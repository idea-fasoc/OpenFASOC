* NGSPICE file created from diff_pair_sample_1502.ext - technology: sky130A

.subckt diff_pair_sample_1502 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t4 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=1.57905 pd=9.9 as=3.7323 ps=19.92 w=9.57 l=3.3
X1 B.t11 B.t9 B.t10 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=0 ps=0 w=9.57 l=3.3
X2 VTAIL.t2 VP.t0 VDD1.t3 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=1.57905 ps=9.9 w=9.57 l=3.3
X3 VDD1.t2 VP.t1 VTAIL.t1 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=1.57905 pd=9.9 as=3.7323 ps=19.92 w=9.57 l=3.3
X4 B.t8 B.t6 B.t7 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=0 ps=0 w=9.57 l=3.3
X5 B.t5 B.t3 B.t4 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=0 ps=0 w=9.57 l=3.3
X6 VTAIL.t0 VP.t2 VDD1.t1 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=1.57905 ps=9.9 w=9.57 l=3.3
X7 VDD2.t2 VN.t1 VTAIL.t5 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=1.57905 pd=9.9 as=3.7323 ps=19.92 w=9.57 l=3.3
X8 VDD1.t0 VP.t3 VTAIL.t7 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=1.57905 pd=9.9 as=3.7323 ps=19.92 w=9.57 l=3.3
X9 B.t2 B.t0 B.t1 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=0 ps=0 w=9.57 l=3.3
X10 VTAIL.t3 VN.t2 VDD2.t1 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=1.57905 ps=9.9 w=9.57 l=3.3
X11 VTAIL.t6 VN.t3 VDD2.t0 w_n3148_n2882# sky130_fd_pr__pfet_01v8 ad=3.7323 pd=19.92 as=1.57905 ps=9.9 w=9.57 l=3.3
R0 VN.n1 VN.t1 104.825
R1 VN.n0 VN.t3 104.825
R2 VN.n0 VN.t0 103.706
R3 VN.n1 VN.t2 103.706
R4 VN VN.n1 49.3386
R5 VN VN.n0 2.48634
R6 VTAIL.n5 VTAIL.t2 63.9563
R7 VTAIL.n4 VTAIL.t5 63.9563
R8 VTAIL.n3 VTAIL.t3 63.9563
R9 VTAIL.n7 VTAIL.t4 63.9562
R10 VTAIL.n0 VTAIL.t6 63.9562
R11 VTAIL.n1 VTAIL.t1 63.9562
R12 VTAIL.n2 VTAIL.t0 63.9562
R13 VTAIL.n6 VTAIL.t7 63.9562
R14 VTAIL.n7 VTAIL.n6 23.7462
R15 VTAIL.n3 VTAIL.n2 23.7462
R16 VTAIL.n4 VTAIL.n3 3.12981
R17 VTAIL.n6 VTAIL.n5 3.12981
R18 VTAIL.n2 VTAIL.n1 3.12981
R19 VTAIL VTAIL.n0 1.62334
R20 VTAIL VTAIL.n7 1.50697
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 118.591
R24 VDD2.n2 VDD2.n1 77.2384
R25 VDD2.n1 VDD2.t1 3.39705
R26 VDD2.n1 VDD2.t2 3.39705
R27 VDD2.n0 VDD2.t0 3.39705
R28 VDD2.n0 VDD2.t3 3.39705
R29 VDD2 VDD2.n2 0.0586897
R30 B.n468 B.n65 585
R31 B.n470 B.n469 585
R32 B.n471 B.n64 585
R33 B.n473 B.n472 585
R34 B.n474 B.n63 585
R35 B.n476 B.n475 585
R36 B.n477 B.n62 585
R37 B.n479 B.n478 585
R38 B.n480 B.n61 585
R39 B.n482 B.n481 585
R40 B.n483 B.n60 585
R41 B.n485 B.n484 585
R42 B.n486 B.n59 585
R43 B.n488 B.n487 585
R44 B.n489 B.n58 585
R45 B.n491 B.n490 585
R46 B.n492 B.n57 585
R47 B.n494 B.n493 585
R48 B.n495 B.n56 585
R49 B.n497 B.n496 585
R50 B.n498 B.n55 585
R51 B.n500 B.n499 585
R52 B.n501 B.n54 585
R53 B.n503 B.n502 585
R54 B.n504 B.n53 585
R55 B.n506 B.n505 585
R56 B.n507 B.n52 585
R57 B.n509 B.n508 585
R58 B.n510 B.n51 585
R59 B.n512 B.n511 585
R60 B.n513 B.n50 585
R61 B.n515 B.n514 585
R62 B.n516 B.n49 585
R63 B.n518 B.n517 585
R64 B.n520 B.n519 585
R65 B.n521 B.n45 585
R66 B.n523 B.n522 585
R67 B.n524 B.n44 585
R68 B.n526 B.n525 585
R69 B.n527 B.n43 585
R70 B.n529 B.n528 585
R71 B.n530 B.n42 585
R72 B.n532 B.n531 585
R73 B.n533 B.n39 585
R74 B.n536 B.n535 585
R75 B.n537 B.n38 585
R76 B.n539 B.n538 585
R77 B.n540 B.n37 585
R78 B.n542 B.n541 585
R79 B.n543 B.n36 585
R80 B.n545 B.n544 585
R81 B.n546 B.n35 585
R82 B.n548 B.n547 585
R83 B.n549 B.n34 585
R84 B.n551 B.n550 585
R85 B.n552 B.n33 585
R86 B.n554 B.n553 585
R87 B.n555 B.n32 585
R88 B.n557 B.n556 585
R89 B.n558 B.n31 585
R90 B.n560 B.n559 585
R91 B.n561 B.n30 585
R92 B.n563 B.n562 585
R93 B.n564 B.n29 585
R94 B.n566 B.n565 585
R95 B.n567 B.n28 585
R96 B.n569 B.n568 585
R97 B.n570 B.n27 585
R98 B.n572 B.n571 585
R99 B.n573 B.n26 585
R100 B.n575 B.n574 585
R101 B.n576 B.n25 585
R102 B.n578 B.n577 585
R103 B.n579 B.n24 585
R104 B.n581 B.n580 585
R105 B.n582 B.n23 585
R106 B.n584 B.n583 585
R107 B.n585 B.n22 585
R108 B.n467 B.n466 585
R109 B.n465 B.n66 585
R110 B.n464 B.n463 585
R111 B.n462 B.n67 585
R112 B.n461 B.n460 585
R113 B.n459 B.n68 585
R114 B.n458 B.n457 585
R115 B.n456 B.n69 585
R116 B.n455 B.n454 585
R117 B.n453 B.n70 585
R118 B.n452 B.n451 585
R119 B.n450 B.n71 585
R120 B.n449 B.n448 585
R121 B.n447 B.n72 585
R122 B.n446 B.n445 585
R123 B.n444 B.n73 585
R124 B.n443 B.n442 585
R125 B.n441 B.n74 585
R126 B.n440 B.n439 585
R127 B.n438 B.n75 585
R128 B.n437 B.n436 585
R129 B.n435 B.n76 585
R130 B.n434 B.n433 585
R131 B.n432 B.n77 585
R132 B.n431 B.n430 585
R133 B.n429 B.n78 585
R134 B.n428 B.n427 585
R135 B.n426 B.n79 585
R136 B.n425 B.n424 585
R137 B.n423 B.n80 585
R138 B.n422 B.n421 585
R139 B.n420 B.n81 585
R140 B.n419 B.n418 585
R141 B.n417 B.n82 585
R142 B.n416 B.n415 585
R143 B.n414 B.n83 585
R144 B.n413 B.n412 585
R145 B.n411 B.n84 585
R146 B.n410 B.n409 585
R147 B.n408 B.n85 585
R148 B.n407 B.n406 585
R149 B.n405 B.n86 585
R150 B.n404 B.n403 585
R151 B.n402 B.n87 585
R152 B.n401 B.n400 585
R153 B.n399 B.n88 585
R154 B.n398 B.n397 585
R155 B.n396 B.n89 585
R156 B.n395 B.n394 585
R157 B.n393 B.n90 585
R158 B.n392 B.n391 585
R159 B.n390 B.n91 585
R160 B.n389 B.n388 585
R161 B.n387 B.n92 585
R162 B.n386 B.n385 585
R163 B.n384 B.n93 585
R164 B.n383 B.n382 585
R165 B.n381 B.n94 585
R166 B.n380 B.n379 585
R167 B.n378 B.n95 585
R168 B.n377 B.n376 585
R169 B.n375 B.n96 585
R170 B.n374 B.n373 585
R171 B.n372 B.n97 585
R172 B.n371 B.n370 585
R173 B.n369 B.n98 585
R174 B.n368 B.n367 585
R175 B.n366 B.n99 585
R176 B.n365 B.n364 585
R177 B.n363 B.n100 585
R178 B.n362 B.n361 585
R179 B.n360 B.n101 585
R180 B.n359 B.n358 585
R181 B.n357 B.n102 585
R182 B.n356 B.n355 585
R183 B.n354 B.n103 585
R184 B.n353 B.n352 585
R185 B.n351 B.n104 585
R186 B.n350 B.n349 585
R187 B.n348 B.n105 585
R188 B.n347 B.n346 585
R189 B.n228 B.n149 585
R190 B.n230 B.n229 585
R191 B.n231 B.n148 585
R192 B.n233 B.n232 585
R193 B.n234 B.n147 585
R194 B.n236 B.n235 585
R195 B.n237 B.n146 585
R196 B.n239 B.n238 585
R197 B.n240 B.n145 585
R198 B.n242 B.n241 585
R199 B.n243 B.n144 585
R200 B.n245 B.n244 585
R201 B.n246 B.n143 585
R202 B.n248 B.n247 585
R203 B.n249 B.n142 585
R204 B.n251 B.n250 585
R205 B.n252 B.n141 585
R206 B.n254 B.n253 585
R207 B.n255 B.n140 585
R208 B.n257 B.n256 585
R209 B.n258 B.n139 585
R210 B.n260 B.n259 585
R211 B.n261 B.n138 585
R212 B.n263 B.n262 585
R213 B.n264 B.n137 585
R214 B.n266 B.n265 585
R215 B.n267 B.n136 585
R216 B.n269 B.n268 585
R217 B.n270 B.n135 585
R218 B.n272 B.n271 585
R219 B.n273 B.n134 585
R220 B.n275 B.n274 585
R221 B.n276 B.n133 585
R222 B.n278 B.n277 585
R223 B.n280 B.n279 585
R224 B.n281 B.n129 585
R225 B.n283 B.n282 585
R226 B.n284 B.n128 585
R227 B.n286 B.n285 585
R228 B.n287 B.n127 585
R229 B.n289 B.n288 585
R230 B.n290 B.n126 585
R231 B.n292 B.n291 585
R232 B.n293 B.n123 585
R233 B.n296 B.n295 585
R234 B.n297 B.n122 585
R235 B.n299 B.n298 585
R236 B.n300 B.n121 585
R237 B.n302 B.n301 585
R238 B.n303 B.n120 585
R239 B.n305 B.n304 585
R240 B.n306 B.n119 585
R241 B.n308 B.n307 585
R242 B.n309 B.n118 585
R243 B.n311 B.n310 585
R244 B.n312 B.n117 585
R245 B.n314 B.n313 585
R246 B.n315 B.n116 585
R247 B.n317 B.n316 585
R248 B.n318 B.n115 585
R249 B.n320 B.n319 585
R250 B.n321 B.n114 585
R251 B.n323 B.n322 585
R252 B.n324 B.n113 585
R253 B.n326 B.n325 585
R254 B.n327 B.n112 585
R255 B.n329 B.n328 585
R256 B.n330 B.n111 585
R257 B.n332 B.n331 585
R258 B.n333 B.n110 585
R259 B.n335 B.n334 585
R260 B.n336 B.n109 585
R261 B.n338 B.n337 585
R262 B.n339 B.n108 585
R263 B.n341 B.n340 585
R264 B.n342 B.n107 585
R265 B.n344 B.n343 585
R266 B.n345 B.n106 585
R267 B.n227 B.n226 585
R268 B.n225 B.n150 585
R269 B.n224 B.n223 585
R270 B.n222 B.n151 585
R271 B.n221 B.n220 585
R272 B.n219 B.n152 585
R273 B.n218 B.n217 585
R274 B.n216 B.n153 585
R275 B.n215 B.n214 585
R276 B.n213 B.n154 585
R277 B.n212 B.n211 585
R278 B.n210 B.n155 585
R279 B.n209 B.n208 585
R280 B.n207 B.n156 585
R281 B.n206 B.n205 585
R282 B.n204 B.n157 585
R283 B.n203 B.n202 585
R284 B.n201 B.n158 585
R285 B.n200 B.n199 585
R286 B.n198 B.n159 585
R287 B.n197 B.n196 585
R288 B.n195 B.n160 585
R289 B.n194 B.n193 585
R290 B.n192 B.n161 585
R291 B.n191 B.n190 585
R292 B.n189 B.n162 585
R293 B.n188 B.n187 585
R294 B.n186 B.n163 585
R295 B.n185 B.n184 585
R296 B.n183 B.n164 585
R297 B.n182 B.n181 585
R298 B.n180 B.n165 585
R299 B.n179 B.n178 585
R300 B.n177 B.n166 585
R301 B.n176 B.n175 585
R302 B.n174 B.n167 585
R303 B.n173 B.n172 585
R304 B.n171 B.n168 585
R305 B.n170 B.n169 585
R306 B.n2 B.n0 585
R307 B.n645 B.n1 585
R308 B.n644 B.n643 585
R309 B.n642 B.n3 585
R310 B.n641 B.n640 585
R311 B.n639 B.n4 585
R312 B.n638 B.n637 585
R313 B.n636 B.n5 585
R314 B.n635 B.n634 585
R315 B.n633 B.n6 585
R316 B.n632 B.n631 585
R317 B.n630 B.n7 585
R318 B.n629 B.n628 585
R319 B.n627 B.n8 585
R320 B.n626 B.n625 585
R321 B.n624 B.n9 585
R322 B.n623 B.n622 585
R323 B.n621 B.n10 585
R324 B.n620 B.n619 585
R325 B.n618 B.n11 585
R326 B.n617 B.n616 585
R327 B.n615 B.n12 585
R328 B.n614 B.n613 585
R329 B.n612 B.n13 585
R330 B.n611 B.n610 585
R331 B.n609 B.n14 585
R332 B.n608 B.n607 585
R333 B.n606 B.n15 585
R334 B.n605 B.n604 585
R335 B.n603 B.n16 585
R336 B.n602 B.n601 585
R337 B.n600 B.n17 585
R338 B.n599 B.n598 585
R339 B.n597 B.n18 585
R340 B.n596 B.n595 585
R341 B.n594 B.n19 585
R342 B.n593 B.n592 585
R343 B.n591 B.n20 585
R344 B.n590 B.n589 585
R345 B.n588 B.n21 585
R346 B.n587 B.n586 585
R347 B.n647 B.n646 585
R348 B.n226 B.n149 564.573
R349 B.n586 B.n585 564.573
R350 B.n346 B.n345 564.573
R351 B.n466 B.n65 564.573
R352 B.n124 B.t6 278.796
R353 B.n130 B.t9 278.796
R354 B.n40 B.t3 278.796
R355 B.n46 B.t0 278.796
R356 B.n124 B.t8 179.206
R357 B.n46 B.t1 179.206
R358 B.n130 B.t11 179.195
R359 B.n40 B.t4 179.195
R360 B.n226 B.n225 163.367
R361 B.n225 B.n224 163.367
R362 B.n224 B.n151 163.367
R363 B.n220 B.n151 163.367
R364 B.n220 B.n219 163.367
R365 B.n219 B.n218 163.367
R366 B.n218 B.n153 163.367
R367 B.n214 B.n153 163.367
R368 B.n214 B.n213 163.367
R369 B.n213 B.n212 163.367
R370 B.n212 B.n155 163.367
R371 B.n208 B.n155 163.367
R372 B.n208 B.n207 163.367
R373 B.n207 B.n206 163.367
R374 B.n206 B.n157 163.367
R375 B.n202 B.n157 163.367
R376 B.n202 B.n201 163.367
R377 B.n201 B.n200 163.367
R378 B.n200 B.n159 163.367
R379 B.n196 B.n159 163.367
R380 B.n196 B.n195 163.367
R381 B.n195 B.n194 163.367
R382 B.n194 B.n161 163.367
R383 B.n190 B.n161 163.367
R384 B.n190 B.n189 163.367
R385 B.n189 B.n188 163.367
R386 B.n188 B.n163 163.367
R387 B.n184 B.n163 163.367
R388 B.n184 B.n183 163.367
R389 B.n183 B.n182 163.367
R390 B.n182 B.n165 163.367
R391 B.n178 B.n165 163.367
R392 B.n178 B.n177 163.367
R393 B.n177 B.n176 163.367
R394 B.n176 B.n167 163.367
R395 B.n172 B.n167 163.367
R396 B.n172 B.n171 163.367
R397 B.n171 B.n170 163.367
R398 B.n170 B.n2 163.367
R399 B.n646 B.n2 163.367
R400 B.n646 B.n645 163.367
R401 B.n645 B.n644 163.367
R402 B.n644 B.n3 163.367
R403 B.n640 B.n3 163.367
R404 B.n640 B.n639 163.367
R405 B.n639 B.n638 163.367
R406 B.n638 B.n5 163.367
R407 B.n634 B.n5 163.367
R408 B.n634 B.n633 163.367
R409 B.n633 B.n632 163.367
R410 B.n632 B.n7 163.367
R411 B.n628 B.n7 163.367
R412 B.n628 B.n627 163.367
R413 B.n627 B.n626 163.367
R414 B.n626 B.n9 163.367
R415 B.n622 B.n9 163.367
R416 B.n622 B.n621 163.367
R417 B.n621 B.n620 163.367
R418 B.n620 B.n11 163.367
R419 B.n616 B.n11 163.367
R420 B.n616 B.n615 163.367
R421 B.n615 B.n614 163.367
R422 B.n614 B.n13 163.367
R423 B.n610 B.n13 163.367
R424 B.n610 B.n609 163.367
R425 B.n609 B.n608 163.367
R426 B.n608 B.n15 163.367
R427 B.n604 B.n15 163.367
R428 B.n604 B.n603 163.367
R429 B.n603 B.n602 163.367
R430 B.n602 B.n17 163.367
R431 B.n598 B.n17 163.367
R432 B.n598 B.n597 163.367
R433 B.n597 B.n596 163.367
R434 B.n596 B.n19 163.367
R435 B.n592 B.n19 163.367
R436 B.n592 B.n591 163.367
R437 B.n591 B.n590 163.367
R438 B.n590 B.n21 163.367
R439 B.n586 B.n21 163.367
R440 B.n230 B.n149 163.367
R441 B.n231 B.n230 163.367
R442 B.n232 B.n231 163.367
R443 B.n232 B.n147 163.367
R444 B.n236 B.n147 163.367
R445 B.n237 B.n236 163.367
R446 B.n238 B.n237 163.367
R447 B.n238 B.n145 163.367
R448 B.n242 B.n145 163.367
R449 B.n243 B.n242 163.367
R450 B.n244 B.n243 163.367
R451 B.n244 B.n143 163.367
R452 B.n248 B.n143 163.367
R453 B.n249 B.n248 163.367
R454 B.n250 B.n249 163.367
R455 B.n250 B.n141 163.367
R456 B.n254 B.n141 163.367
R457 B.n255 B.n254 163.367
R458 B.n256 B.n255 163.367
R459 B.n256 B.n139 163.367
R460 B.n260 B.n139 163.367
R461 B.n261 B.n260 163.367
R462 B.n262 B.n261 163.367
R463 B.n262 B.n137 163.367
R464 B.n266 B.n137 163.367
R465 B.n267 B.n266 163.367
R466 B.n268 B.n267 163.367
R467 B.n268 B.n135 163.367
R468 B.n272 B.n135 163.367
R469 B.n273 B.n272 163.367
R470 B.n274 B.n273 163.367
R471 B.n274 B.n133 163.367
R472 B.n278 B.n133 163.367
R473 B.n279 B.n278 163.367
R474 B.n279 B.n129 163.367
R475 B.n283 B.n129 163.367
R476 B.n284 B.n283 163.367
R477 B.n285 B.n284 163.367
R478 B.n285 B.n127 163.367
R479 B.n289 B.n127 163.367
R480 B.n290 B.n289 163.367
R481 B.n291 B.n290 163.367
R482 B.n291 B.n123 163.367
R483 B.n296 B.n123 163.367
R484 B.n297 B.n296 163.367
R485 B.n298 B.n297 163.367
R486 B.n298 B.n121 163.367
R487 B.n302 B.n121 163.367
R488 B.n303 B.n302 163.367
R489 B.n304 B.n303 163.367
R490 B.n304 B.n119 163.367
R491 B.n308 B.n119 163.367
R492 B.n309 B.n308 163.367
R493 B.n310 B.n309 163.367
R494 B.n310 B.n117 163.367
R495 B.n314 B.n117 163.367
R496 B.n315 B.n314 163.367
R497 B.n316 B.n315 163.367
R498 B.n316 B.n115 163.367
R499 B.n320 B.n115 163.367
R500 B.n321 B.n320 163.367
R501 B.n322 B.n321 163.367
R502 B.n322 B.n113 163.367
R503 B.n326 B.n113 163.367
R504 B.n327 B.n326 163.367
R505 B.n328 B.n327 163.367
R506 B.n328 B.n111 163.367
R507 B.n332 B.n111 163.367
R508 B.n333 B.n332 163.367
R509 B.n334 B.n333 163.367
R510 B.n334 B.n109 163.367
R511 B.n338 B.n109 163.367
R512 B.n339 B.n338 163.367
R513 B.n340 B.n339 163.367
R514 B.n340 B.n107 163.367
R515 B.n344 B.n107 163.367
R516 B.n345 B.n344 163.367
R517 B.n346 B.n105 163.367
R518 B.n350 B.n105 163.367
R519 B.n351 B.n350 163.367
R520 B.n352 B.n351 163.367
R521 B.n352 B.n103 163.367
R522 B.n356 B.n103 163.367
R523 B.n357 B.n356 163.367
R524 B.n358 B.n357 163.367
R525 B.n358 B.n101 163.367
R526 B.n362 B.n101 163.367
R527 B.n363 B.n362 163.367
R528 B.n364 B.n363 163.367
R529 B.n364 B.n99 163.367
R530 B.n368 B.n99 163.367
R531 B.n369 B.n368 163.367
R532 B.n370 B.n369 163.367
R533 B.n370 B.n97 163.367
R534 B.n374 B.n97 163.367
R535 B.n375 B.n374 163.367
R536 B.n376 B.n375 163.367
R537 B.n376 B.n95 163.367
R538 B.n380 B.n95 163.367
R539 B.n381 B.n380 163.367
R540 B.n382 B.n381 163.367
R541 B.n382 B.n93 163.367
R542 B.n386 B.n93 163.367
R543 B.n387 B.n386 163.367
R544 B.n388 B.n387 163.367
R545 B.n388 B.n91 163.367
R546 B.n392 B.n91 163.367
R547 B.n393 B.n392 163.367
R548 B.n394 B.n393 163.367
R549 B.n394 B.n89 163.367
R550 B.n398 B.n89 163.367
R551 B.n399 B.n398 163.367
R552 B.n400 B.n399 163.367
R553 B.n400 B.n87 163.367
R554 B.n404 B.n87 163.367
R555 B.n405 B.n404 163.367
R556 B.n406 B.n405 163.367
R557 B.n406 B.n85 163.367
R558 B.n410 B.n85 163.367
R559 B.n411 B.n410 163.367
R560 B.n412 B.n411 163.367
R561 B.n412 B.n83 163.367
R562 B.n416 B.n83 163.367
R563 B.n417 B.n416 163.367
R564 B.n418 B.n417 163.367
R565 B.n418 B.n81 163.367
R566 B.n422 B.n81 163.367
R567 B.n423 B.n422 163.367
R568 B.n424 B.n423 163.367
R569 B.n424 B.n79 163.367
R570 B.n428 B.n79 163.367
R571 B.n429 B.n428 163.367
R572 B.n430 B.n429 163.367
R573 B.n430 B.n77 163.367
R574 B.n434 B.n77 163.367
R575 B.n435 B.n434 163.367
R576 B.n436 B.n435 163.367
R577 B.n436 B.n75 163.367
R578 B.n440 B.n75 163.367
R579 B.n441 B.n440 163.367
R580 B.n442 B.n441 163.367
R581 B.n442 B.n73 163.367
R582 B.n446 B.n73 163.367
R583 B.n447 B.n446 163.367
R584 B.n448 B.n447 163.367
R585 B.n448 B.n71 163.367
R586 B.n452 B.n71 163.367
R587 B.n453 B.n452 163.367
R588 B.n454 B.n453 163.367
R589 B.n454 B.n69 163.367
R590 B.n458 B.n69 163.367
R591 B.n459 B.n458 163.367
R592 B.n460 B.n459 163.367
R593 B.n460 B.n67 163.367
R594 B.n464 B.n67 163.367
R595 B.n465 B.n464 163.367
R596 B.n466 B.n465 163.367
R597 B.n585 B.n584 163.367
R598 B.n584 B.n23 163.367
R599 B.n580 B.n23 163.367
R600 B.n580 B.n579 163.367
R601 B.n579 B.n578 163.367
R602 B.n578 B.n25 163.367
R603 B.n574 B.n25 163.367
R604 B.n574 B.n573 163.367
R605 B.n573 B.n572 163.367
R606 B.n572 B.n27 163.367
R607 B.n568 B.n27 163.367
R608 B.n568 B.n567 163.367
R609 B.n567 B.n566 163.367
R610 B.n566 B.n29 163.367
R611 B.n562 B.n29 163.367
R612 B.n562 B.n561 163.367
R613 B.n561 B.n560 163.367
R614 B.n560 B.n31 163.367
R615 B.n556 B.n31 163.367
R616 B.n556 B.n555 163.367
R617 B.n555 B.n554 163.367
R618 B.n554 B.n33 163.367
R619 B.n550 B.n33 163.367
R620 B.n550 B.n549 163.367
R621 B.n549 B.n548 163.367
R622 B.n548 B.n35 163.367
R623 B.n544 B.n35 163.367
R624 B.n544 B.n543 163.367
R625 B.n543 B.n542 163.367
R626 B.n542 B.n37 163.367
R627 B.n538 B.n37 163.367
R628 B.n538 B.n537 163.367
R629 B.n537 B.n536 163.367
R630 B.n536 B.n39 163.367
R631 B.n531 B.n39 163.367
R632 B.n531 B.n530 163.367
R633 B.n530 B.n529 163.367
R634 B.n529 B.n43 163.367
R635 B.n525 B.n43 163.367
R636 B.n525 B.n524 163.367
R637 B.n524 B.n523 163.367
R638 B.n523 B.n45 163.367
R639 B.n519 B.n45 163.367
R640 B.n519 B.n518 163.367
R641 B.n518 B.n49 163.367
R642 B.n514 B.n49 163.367
R643 B.n514 B.n513 163.367
R644 B.n513 B.n512 163.367
R645 B.n512 B.n51 163.367
R646 B.n508 B.n51 163.367
R647 B.n508 B.n507 163.367
R648 B.n507 B.n506 163.367
R649 B.n506 B.n53 163.367
R650 B.n502 B.n53 163.367
R651 B.n502 B.n501 163.367
R652 B.n501 B.n500 163.367
R653 B.n500 B.n55 163.367
R654 B.n496 B.n55 163.367
R655 B.n496 B.n495 163.367
R656 B.n495 B.n494 163.367
R657 B.n494 B.n57 163.367
R658 B.n490 B.n57 163.367
R659 B.n490 B.n489 163.367
R660 B.n489 B.n488 163.367
R661 B.n488 B.n59 163.367
R662 B.n484 B.n59 163.367
R663 B.n484 B.n483 163.367
R664 B.n483 B.n482 163.367
R665 B.n482 B.n61 163.367
R666 B.n478 B.n61 163.367
R667 B.n478 B.n477 163.367
R668 B.n477 B.n476 163.367
R669 B.n476 B.n63 163.367
R670 B.n472 B.n63 163.367
R671 B.n472 B.n471 163.367
R672 B.n471 B.n470 163.367
R673 B.n470 B.n65 163.367
R674 B.n125 B.t7 108.805
R675 B.n47 B.t2 108.805
R676 B.n131 B.t10 108.794
R677 B.n41 B.t5 108.794
R678 B.n125 B.n124 70.4005
R679 B.n131 B.n130 70.4005
R680 B.n41 B.n40 70.4005
R681 B.n47 B.n46 70.4005
R682 B.n294 B.n125 59.5399
R683 B.n132 B.n131 59.5399
R684 B.n534 B.n41 59.5399
R685 B.n48 B.n47 59.5399
R686 B.n587 B.n22 36.6834
R687 B.n347 B.n106 36.6834
R688 B.n228 B.n227 36.6834
R689 B.n468 B.n467 36.6834
R690 B B.n647 18.0485
R691 B.n583 B.n22 10.6151
R692 B.n583 B.n582 10.6151
R693 B.n582 B.n581 10.6151
R694 B.n581 B.n24 10.6151
R695 B.n577 B.n24 10.6151
R696 B.n577 B.n576 10.6151
R697 B.n576 B.n575 10.6151
R698 B.n575 B.n26 10.6151
R699 B.n571 B.n26 10.6151
R700 B.n571 B.n570 10.6151
R701 B.n570 B.n569 10.6151
R702 B.n569 B.n28 10.6151
R703 B.n565 B.n28 10.6151
R704 B.n565 B.n564 10.6151
R705 B.n564 B.n563 10.6151
R706 B.n563 B.n30 10.6151
R707 B.n559 B.n30 10.6151
R708 B.n559 B.n558 10.6151
R709 B.n558 B.n557 10.6151
R710 B.n557 B.n32 10.6151
R711 B.n553 B.n32 10.6151
R712 B.n553 B.n552 10.6151
R713 B.n552 B.n551 10.6151
R714 B.n551 B.n34 10.6151
R715 B.n547 B.n34 10.6151
R716 B.n547 B.n546 10.6151
R717 B.n546 B.n545 10.6151
R718 B.n545 B.n36 10.6151
R719 B.n541 B.n36 10.6151
R720 B.n541 B.n540 10.6151
R721 B.n540 B.n539 10.6151
R722 B.n539 B.n38 10.6151
R723 B.n535 B.n38 10.6151
R724 B.n533 B.n532 10.6151
R725 B.n532 B.n42 10.6151
R726 B.n528 B.n42 10.6151
R727 B.n528 B.n527 10.6151
R728 B.n527 B.n526 10.6151
R729 B.n526 B.n44 10.6151
R730 B.n522 B.n44 10.6151
R731 B.n522 B.n521 10.6151
R732 B.n521 B.n520 10.6151
R733 B.n517 B.n516 10.6151
R734 B.n516 B.n515 10.6151
R735 B.n515 B.n50 10.6151
R736 B.n511 B.n50 10.6151
R737 B.n511 B.n510 10.6151
R738 B.n510 B.n509 10.6151
R739 B.n509 B.n52 10.6151
R740 B.n505 B.n52 10.6151
R741 B.n505 B.n504 10.6151
R742 B.n504 B.n503 10.6151
R743 B.n503 B.n54 10.6151
R744 B.n499 B.n54 10.6151
R745 B.n499 B.n498 10.6151
R746 B.n498 B.n497 10.6151
R747 B.n497 B.n56 10.6151
R748 B.n493 B.n56 10.6151
R749 B.n493 B.n492 10.6151
R750 B.n492 B.n491 10.6151
R751 B.n491 B.n58 10.6151
R752 B.n487 B.n58 10.6151
R753 B.n487 B.n486 10.6151
R754 B.n486 B.n485 10.6151
R755 B.n485 B.n60 10.6151
R756 B.n481 B.n60 10.6151
R757 B.n481 B.n480 10.6151
R758 B.n480 B.n479 10.6151
R759 B.n479 B.n62 10.6151
R760 B.n475 B.n62 10.6151
R761 B.n475 B.n474 10.6151
R762 B.n474 B.n473 10.6151
R763 B.n473 B.n64 10.6151
R764 B.n469 B.n64 10.6151
R765 B.n469 B.n468 10.6151
R766 B.n348 B.n347 10.6151
R767 B.n349 B.n348 10.6151
R768 B.n349 B.n104 10.6151
R769 B.n353 B.n104 10.6151
R770 B.n354 B.n353 10.6151
R771 B.n355 B.n354 10.6151
R772 B.n355 B.n102 10.6151
R773 B.n359 B.n102 10.6151
R774 B.n360 B.n359 10.6151
R775 B.n361 B.n360 10.6151
R776 B.n361 B.n100 10.6151
R777 B.n365 B.n100 10.6151
R778 B.n366 B.n365 10.6151
R779 B.n367 B.n366 10.6151
R780 B.n367 B.n98 10.6151
R781 B.n371 B.n98 10.6151
R782 B.n372 B.n371 10.6151
R783 B.n373 B.n372 10.6151
R784 B.n373 B.n96 10.6151
R785 B.n377 B.n96 10.6151
R786 B.n378 B.n377 10.6151
R787 B.n379 B.n378 10.6151
R788 B.n379 B.n94 10.6151
R789 B.n383 B.n94 10.6151
R790 B.n384 B.n383 10.6151
R791 B.n385 B.n384 10.6151
R792 B.n385 B.n92 10.6151
R793 B.n389 B.n92 10.6151
R794 B.n390 B.n389 10.6151
R795 B.n391 B.n390 10.6151
R796 B.n391 B.n90 10.6151
R797 B.n395 B.n90 10.6151
R798 B.n396 B.n395 10.6151
R799 B.n397 B.n396 10.6151
R800 B.n397 B.n88 10.6151
R801 B.n401 B.n88 10.6151
R802 B.n402 B.n401 10.6151
R803 B.n403 B.n402 10.6151
R804 B.n403 B.n86 10.6151
R805 B.n407 B.n86 10.6151
R806 B.n408 B.n407 10.6151
R807 B.n409 B.n408 10.6151
R808 B.n409 B.n84 10.6151
R809 B.n413 B.n84 10.6151
R810 B.n414 B.n413 10.6151
R811 B.n415 B.n414 10.6151
R812 B.n415 B.n82 10.6151
R813 B.n419 B.n82 10.6151
R814 B.n420 B.n419 10.6151
R815 B.n421 B.n420 10.6151
R816 B.n421 B.n80 10.6151
R817 B.n425 B.n80 10.6151
R818 B.n426 B.n425 10.6151
R819 B.n427 B.n426 10.6151
R820 B.n427 B.n78 10.6151
R821 B.n431 B.n78 10.6151
R822 B.n432 B.n431 10.6151
R823 B.n433 B.n432 10.6151
R824 B.n433 B.n76 10.6151
R825 B.n437 B.n76 10.6151
R826 B.n438 B.n437 10.6151
R827 B.n439 B.n438 10.6151
R828 B.n439 B.n74 10.6151
R829 B.n443 B.n74 10.6151
R830 B.n444 B.n443 10.6151
R831 B.n445 B.n444 10.6151
R832 B.n445 B.n72 10.6151
R833 B.n449 B.n72 10.6151
R834 B.n450 B.n449 10.6151
R835 B.n451 B.n450 10.6151
R836 B.n451 B.n70 10.6151
R837 B.n455 B.n70 10.6151
R838 B.n456 B.n455 10.6151
R839 B.n457 B.n456 10.6151
R840 B.n457 B.n68 10.6151
R841 B.n461 B.n68 10.6151
R842 B.n462 B.n461 10.6151
R843 B.n463 B.n462 10.6151
R844 B.n463 B.n66 10.6151
R845 B.n467 B.n66 10.6151
R846 B.n229 B.n228 10.6151
R847 B.n229 B.n148 10.6151
R848 B.n233 B.n148 10.6151
R849 B.n234 B.n233 10.6151
R850 B.n235 B.n234 10.6151
R851 B.n235 B.n146 10.6151
R852 B.n239 B.n146 10.6151
R853 B.n240 B.n239 10.6151
R854 B.n241 B.n240 10.6151
R855 B.n241 B.n144 10.6151
R856 B.n245 B.n144 10.6151
R857 B.n246 B.n245 10.6151
R858 B.n247 B.n246 10.6151
R859 B.n247 B.n142 10.6151
R860 B.n251 B.n142 10.6151
R861 B.n252 B.n251 10.6151
R862 B.n253 B.n252 10.6151
R863 B.n253 B.n140 10.6151
R864 B.n257 B.n140 10.6151
R865 B.n258 B.n257 10.6151
R866 B.n259 B.n258 10.6151
R867 B.n259 B.n138 10.6151
R868 B.n263 B.n138 10.6151
R869 B.n264 B.n263 10.6151
R870 B.n265 B.n264 10.6151
R871 B.n265 B.n136 10.6151
R872 B.n269 B.n136 10.6151
R873 B.n270 B.n269 10.6151
R874 B.n271 B.n270 10.6151
R875 B.n271 B.n134 10.6151
R876 B.n275 B.n134 10.6151
R877 B.n276 B.n275 10.6151
R878 B.n277 B.n276 10.6151
R879 B.n281 B.n280 10.6151
R880 B.n282 B.n281 10.6151
R881 B.n282 B.n128 10.6151
R882 B.n286 B.n128 10.6151
R883 B.n287 B.n286 10.6151
R884 B.n288 B.n287 10.6151
R885 B.n288 B.n126 10.6151
R886 B.n292 B.n126 10.6151
R887 B.n293 B.n292 10.6151
R888 B.n295 B.n122 10.6151
R889 B.n299 B.n122 10.6151
R890 B.n300 B.n299 10.6151
R891 B.n301 B.n300 10.6151
R892 B.n301 B.n120 10.6151
R893 B.n305 B.n120 10.6151
R894 B.n306 B.n305 10.6151
R895 B.n307 B.n306 10.6151
R896 B.n307 B.n118 10.6151
R897 B.n311 B.n118 10.6151
R898 B.n312 B.n311 10.6151
R899 B.n313 B.n312 10.6151
R900 B.n313 B.n116 10.6151
R901 B.n317 B.n116 10.6151
R902 B.n318 B.n317 10.6151
R903 B.n319 B.n318 10.6151
R904 B.n319 B.n114 10.6151
R905 B.n323 B.n114 10.6151
R906 B.n324 B.n323 10.6151
R907 B.n325 B.n324 10.6151
R908 B.n325 B.n112 10.6151
R909 B.n329 B.n112 10.6151
R910 B.n330 B.n329 10.6151
R911 B.n331 B.n330 10.6151
R912 B.n331 B.n110 10.6151
R913 B.n335 B.n110 10.6151
R914 B.n336 B.n335 10.6151
R915 B.n337 B.n336 10.6151
R916 B.n337 B.n108 10.6151
R917 B.n341 B.n108 10.6151
R918 B.n342 B.n341 10.6151
R919 B.n343 B.n342 10.6151
R920 B.n343 B.n106 10.6151
R921 B.n227 B.n150 10.6151
R922 B.n223 B.n150 10.6151
R923 B.n223 B.n222 10.6151
R924 B.n222 B.n221 10.6151
R925 B.n221 B.n152 10.6151
R926 B.n217 B.n152 10.6151
R927 B.n217 B.n216 10.6151
R928 B.n216 B.n215 10.6151
R929 B.n215 B.n154 10.6151
R930 B.n211 B.n154 10.6151
R931 B.n211 B.n210 10.6151
R932 B.n210 B.n209 10.6151
R933 B.n209 B.n156 10.6151
R934 B.n205 B.n156 10.6151
R935 B.n205 B.n204 10.6151
R936 B.n204 B.n203 10.6151
R937 B.n203 B.n158 10.6151
R938 B.n199 B.n158 10.6151
R939 B.n199 B.n198 10.6151
R940 B.n198 B.n197 10.6151
R941 B.n197 B.n160 10.6151
R942 B.n193 B.n160 10.6151
R943 B.n193 B.n192 10.6151
R944 B.n192 B.n191 10.6151
R945 B.n191 B.n162 10.6151
R946 B.n187 B.n162 10.6151
R947 B.n187 B.n186 10.6151
R948 B.n186 B.n185 10.6151
R949 B.n185 B.n164 10.6151
R950 B.n181 B.n164 10.6151
R951 B.n181 B.n180 10.6151
R952 B.n180 B.n179 10.6151
R953 B.n179 B.n166 10.6151
R954 B.n175 B.n166 10.6151
R955 B.n175 B.n174 10.6151
R956 B.n174 B.n173 10.6151
R957 B.n173 B.n168 10.6151
R958 B.n169 B.n168 10.6151
R959 B.n169 B.n0 10.6151
R960 B.n643 B.n1 10.6151
R961 B.n643 B.n642 10.6151
R962 B.n642 B.n641 10.6151
R963 B.n641 B.n4 10.6151
R964 B.n637 B.n4 10.6151
R965 B.n637 B.n636 10.6151
R966 B.n636 B.n635 10.6151
R967 B.n635 B.n6 10.6151
R968 B.n631 B.n6 10.6151
R969 B.n631 B.n630 10.6151
R970 B.n630 B.n629 10.6151
R971 B.n629 B.n8 10.6151
R972 B.n625 B.n8 10.6151
R973 B.n625 B.n624 10.6151
R974 B.n624 B.n623 10.6151
R975 B.n623 B.n10 10.6151
R976 B.n619 B.n10 10.6151
R977 B.n619 B.n618 10.6151
R978 B.n618 B.n617 10.6151
R979 B.n617 B.n12 10.6151
R980 B.n613 B.n12 10.6151
R981 B.n613 B.n612 10.6151
R982 B.n612 B.n611 10.6151
R983 B.n611 B.n14 10.6151
R984 B.n607 B.n14 10.6151
R985 B.n607 B.n606 10.6151
R986 B.n606 B.n605 10.6151
R987 B.n605 B.n16 10.6151
R988 B.n601 B.n16 10.6151
R989 B.n601 B.n600 10.6151
R990 B.n600 B.n599 10.6151
R991 B.n599 B.n18 10.6151
R992 B.n595 B.n18 10.6151
R993 B.n595 B.n594 10.6151
R994 B.n594 B.n593 10.6151
R995 B.n593 B.n20 10.6151
R996 B.n589 B.n20 10.6151
R997 B.n589 B.n588 10.6151
R998 B.n588 B.n587 10.6151
R999 B.n535 B.n534 9.36635
R1000 B.n517 B.n48 9.36635
R1001 B.n277 B.n132 9.36635
R1002 B.n295 B.n294 9.36635
R1003 B.n647 B.n0 2.81026
R1004 B.n647 B.n1 2.81026
R1005 B.n534 B.n533 1.24928
R1006 B.n520 B.n48 1.24928
R1007 B.n280 B.n132 1.24928
R1008 B.n294 B.n293 1.24928
R1009 VP.n17 VP.n16 161.3
R1010 VP.n15 VP.n1 161.3
R1011 VP.n14 VP.n13 161.3
R1012 VP.n12 VP.n2 161.3
R1013 VP.n11 VP.n10 161.3
R1014 VP.n9 VP.n3 161.3
R1015 VP.n8 VP.n7 161.3
R1016 VP.n5 VP.t0 104.825
R1017 VP.n5 VP.t3 103.706
R1018 VP.n6 VP.n4 74.6532
R1019 VP.n18 VP.n0 74.6532
R1020 VP.n4 VP.t2 69.8905
R1021 VP.n0 VP.t1 69.8905
R1022 VP.n6 VP.n5 49.1732
R1023 VP.n10 VP.n2 40.4934
R1024 VP.n14 VP.n2 40.4934
R1025 VP.n9 VP.n8 24.4675
R1026 VP.n10 VP.n9 24.4675
R1027 VP.n15 VP.n14 24.4675
R1028 VP.n16 VP.n15 24.4675
R1029 VP.n8 VP.n4 15.4147
R1030 VP.n16 VP.n0 15.4147
R1031 VP.n7 VP.n6 0.354971
R1032 VP.n18 VP.n17 0.354971
R1033 VP VP.n18 0.26696
R1034 VP.n7 VP.n3 0.189894
R1035 VP.n11 VP.n3 0.189894
R1036 VP.n12 VP.n11 0.189894
R1037 VP.n13 VP.n12 0.189894
R1038 VP.n13 VP.n1 0.189894
R1039 VP.n17 VP.n1 0.189894
R1040 VDD1 VDD1.n1 119.115
R1041 VDD1 VDD1.n0 77.2966
R1042 VDD1.n0 VDD1.t3 3.39705
R1043 VDD1.n0 VDD1.t0 3.39705
R1044 VDD1.n1 VDD1.t1 3.39705
R1045 VDD1.n1 VDD1.t2 3.39705
C0 VP VDD1 4.29483f
C1 B VDD2 1.38369f
C2 VTAIL VDD2 5.10471f
C3 VN VDD2 4.00653f
C4 VP VDD2 0.438694f
C5 B w_n3148_n2882# 9.42482f
C6 VTAIL w_n3148_n2882# 3.46225f
C7 VDD1 VDD2 1.18967f
C8 VN w_n3148_n2882# 5.41757f
C9 VP w_n3148_n2882# 5.82403f
C10 w_n3148_n2882# VDD1 1.51751f
C11 B VTAIL 4.4137f
C12 B VN 1.21312f
C13 VP B 1.89087f
C14 VN VTAIL 4.1295f
C15 VP VTAIL 4.1436f
C16 VP VN 6.24575f
C17 B VDD1 1.31994f
C18 w_n3148_n2882# VDD2 1.5891f
C19 VTAIL VDD1 5.0458f
C20 VN VDD1 0.149479f
C21 VDD2 VSUBS 1.009484f
C22 VDD1 VSUBS 5.83105f
C23 VTAIL VSUBS 1.193881f
C24 VN VSUBS 5.79352f
C25 VP VSUBS 2.573714f
C26 B VSUBS 4.673398f
C27 w_n3148_n2882# VSUBS 0.112157p
C28 VDD1.t3 VSUBS 0.209201f
C29 VDD1.t0 VSUBS 0.209201f
C30 VDD1.n0 VSUBS 1.56471f
C31 VDD1.t1 VSUBS 0.209201f
C32 VDD1.t2 VSUBS 0.209201f
C33 VDD1.n1 VSUBS 2.24226f
C34 VP.t1 VSUBS 2.7557f
C35 VP.n0 VSUBS 1.10987f
C36 VP.n1 VSUBS 0.03226f
C37 VP.n2 VSUBS 0.026079f
C38 VP.n3 VSUBS 0.03226f
C39 VP.t2 VSUBS 2.7557f
C40 VP.n4 VSUBS 1.10987f
C41 VP.t0 VSUBS 3.16411f
C42 VP.t3 VSUBS 3.15156f
C43 VP.n5 VSUBS 3.78057f
C44 VP.n6 VSUBS 1.79009f
C45 VP.n7 VSUBS 0.052067f
C46 VP.n8 VSUBS 0.04914f
C47 VP.n9 VSUBS 0.060124f
C48 VP.n10 VSUBS 0.064116f
C49 VP.n11 VSUBS 0.03226f
C50 VP.n12 VSUBS 0.03226f
C51 VP.n13 VSUBS 0.03226f
C52 VP.n14 VSUBS 0.064116f
C53 VP.n15 VSUBS 0.060124f
C54 VP.n16 VSUBS 0.04914f
C55 VP.n17 VSUBS 0.052067f
C56 VP.n18 VSUBS 0.077094f
C57 B.n0 VSUBS 0.004315f
C58 B.n1 VSUBS 0.004315f
C59 B.n2 VSUBS 0.006824f
C60 B.n3 VSUBS 0.006824f
C61 B.n4 VSUBS 0.006824f
C62 B.n5 VSUBS 0.006824f
C63 B.n6 VSUBS 0.006824f
C64 B.n7 VSUBS 0.006824f
C65 B.n8 VSUBS 0.006824f
C66 B.n9 VSUBS 0.006824f
C67 B.n10 VSUBS 0.006824f
C68 B.n11 VSUBS 0.006824f
C69 B.n12 VSUBS 0.006824f
C70 B.n13 VSUBS 0.006824f
C71 B.n14 VSUBS 0.006824f
C72 B.n15 VSUBS 0.006824f
C73 B.n16 VSUBS 0.006824f
C74 B.n17 VSUBS 0.006824f
C75 B.n18 VSUBS 0.006824f
C76 B.n19 VSUBS 0.006824f
C77 B.n20 VSUBS 0.006824f
C78 B.n21 VSUBS 0.006824f
C79 B.n22 VSUBS 0.017532f
C80 B.n23 VSUBS 0.006824f
C81 B.n24 VSUBS 0.006824f
C82 B.n25 VSUBS 0.006824f
C83 B.n26 VSUBS 0.006824f
C84 B.n27 VSUBS 0.006824f
C85 B.n28 VSUBS 0.006824f
C86 B.n29 VSUBS 0.006824f
C87 B.n30 VSUBS 0.006824f
C88 B.n31 VSUBS 0.006824f
C89 B.n32 VSUBS 0.006824f
C90 B.n33 VSUBS 0.006824f
C91 B.n34 VSUBS 0.006824f
C92 B.n35 VSUBS 0.006824f
C93 B.n36 VSUBS 0.006824f
C94 B.n37 VSUBS 0.006824f
C95 B.n38 VSUBS 0.006824f
C96 B.n39 VSUBS 0.006824f
C97 B.t5 VSUBS 0.295799f
C98 B.t4 VSUBS 0.320502f
C99 B.t3 VSUBS 1.44132f
C100 B.n40 VSUBS 0.177519f
C101 B.n41 VSUBS 0.07261f
C102 B.n42 VSUBS 0.006824f
C103 B.n43 VSUBS 0.006824f
C104 B.n44 VSUBS 0.006824f
C105 B.n45 VSUBS 0.006824f
C106 B.t2 VSUBS 0.295796f
C107 B.t1 VSUBS 0.320498f
C108 B.t0 VSUBS 1.44132f
C109 B.n46 VSUBS 0.177523f
C110 B.n47 VSUBS 0.072614f
C111 B.n48 VSUBS 0.015811f
C112 B.n49 VSUBS 0.006824f
C113 B.n50 VSUBS 0.006824f
C114 B.n51 VSUBS 0.006824f
C115 B.n52 VSUBS 0.006824f
C116 B.n53 VSUBS 0.006824f
C117 B.n54 VSUBS 0.006824f
C118 B.n55 VSUBS 0.006824f
C119 B.n56 VSUBS 0.006824f
C120 B.n57 VSUBS 0.006824f
C121 B.n58 VSUBS 0.006824f
C122 B.n59 VSUBS 0.006824f
C123 B.n60 VSUBS 0.006824f
C124 B.n61 VSUBS 0.006824f
C125 B.n62 VSUBS 0.006824f
C126 B.n63 VSUBS 0.006824f
C127 B.n64 VSUBS 0.006824f
C128 B.n65 VSUBS 0.017532f
C129 B.n66 VSUBS 0.006824f
C130 B.n67 VSUBS 0.006824f
C131 B.n68 VSUBS 0.006824f
C132 B.n69 VSUBS 0.006824f
C133 B.n70 VSUBS 0.006824f
C134 B.n71 VSUBS 0.006824f
C135 B.n72 VSUBS 0.006824f
C136 B.n73 VSUBS 0.006824f
C137 B.n74 VSUBS 0.006824f
C138 B.n75 VSUBS 0.006824f
C139 B.n76 VSUBS 0.006824f
C140 B.n77 VSUBS 0.006824f
C141 B.n78 VSUBS 0.006824f
C142 B.n79 VSUBS 0.006824f
C143 B.n80 VSUBS 0.006824f
C144 B.n81 VSUBS 0.006824f
C145 B.n82 VSUBS 0.006824f
C146 B.n83 VSUBS 0.006824f
C147 B.n84 VSUBS 0.006824f
C148 B.n85 VSUBS 0.006824f
C149 B.n86 VSUBS 0.006824f
C150 B.n87 VSUBS 0.006824f
C151 B.n88 VSUBS 0.006824f
C152 B.n89 VSUBS 0.006824f
C153 B.n90 VSUBS 0.006824f
C154 B.n91 VSUBS 0.006824f
C155 B.n92 VSUBS 0.006824f
C156 B.n93 VSUBS 0.006824f
C157 B.n94 VSUBS 0.006824f
C158 B.n95 VSUBS 0.006824f
C159 B.n96 VSUBS 0.006824f
C160 B.n97 VSUBS 0.006824f
C161 B.n98 VSUBS 0.006824f
C162 B.n99 VSUBS 0.006824f
C163 B.n100 VSUBS 0.006824f
C164 B.n101 VSUBS 0.006824f
C165 B.n102 VSUBS 0.006824f
C166 B.n103 VSUBS 0.006824f
C167 B.n104 VSUBS 0.006824f
C168 B.n105 VSUBS 0.006824f
C169 B.n106 VSUBS 0.017532f
C170 B.n107 VSUBS 0.006824f
C171 B.n108 VSUBS 0.006824f
C172 B.n109 VSUBS 0.006824f
C173 B.n110 VSUBS 0.006824f
C174 B.n111 VSUBS 0.006824f
C175 B.n112 VSUBS 0.006824f
C176 B.n113 VSUBS 0.006824f
C177 B.n114 VSUBS 0.006824f
C178 B.n115 VSUBS 0.006824f
C179 B.n116 VSUBS 0.006824f
C180 B.n117 VSUBS 0.006824f
C181 B.n118 VSUBS 0.006824f
C182 B.n119 VSUBS 0.006824f
C183 B.n120 VSUBS 0.006824f
C184 B.n121 VSUBS 0.006824f
C185 B.n122 VSUBS 0.006824f
C186 B.n123 VSUBS 0.006824f
C187 B.t7 VSUBS 0.295796f
C188 B.t8 VSUBS 0.320498f
C189 B.t6 VSUBS 1.44132f
C190 B.n124 VSUBS 0.177523f
C191 B.n125 VSUBS 0.072614f
C192 B.n126 VSUBS 0.006824f
C193 B.n127 VSUBS 0.006824f
C194 B.n128 VSUBS 0.006824f
C195 B.n129 VSUBS 0.006824f
C196 B.t10 VSUBS 0.295799f
C197 B.t11 VSUBS 0.320502f
C198 B.t9 VSUBS 1.44132f
C199 B.n130 VSUBS 0.177519f
C200 B.n131 VSUBS 0.07261f
C201 B.n132 VSUBS 0.015811f
C202 B.n133 VSUBS 0.006824f
C203 B.n134 VSUBS 0.006824f
C204 B.n135 VSUBS 0.006824f
C205 B.n136 VSUBS 0.006824f
C206 B.n137 VSUBS 0.006824f
C207 B.n138 VSUBS 0.006824f
C208 B.n139 VSUBS 0.006824f
C209 B.n140 VSUBS 0.006824f
C210 B.n141 VSUBS 0.006824f
C211 B.n142 VSUBS 0.006824f
C212 B.n143 VSUBS 0.006824f
C213 B.n144 VSUBS 0.006824f
C214 B.n145 VSUBS 0.006824f
C215 B.n146 VSUBS 0.006824f
C216 B.n147 VSUBS 0.006824f
C217 B.n148 VSUBS 0.006824f
C218 B.n149 VSUBS 0.017532f
C219 B.n150 VSUBS 0.006824f
C220 B.n151 VSUBS 0.006824f
C221 B.n152 VSUBS 0.006824f
C222 B.n153 VSUBS 0.006824f
C223 B.n154 VSUBS 0.006824f
C224 B.n155 VSUBS 0.006824f
C225 B.n156 VSUBS 0.006824f
C226 B.n157 VSUBS 0.006824f
C227 B.n158 VSUBS 0.006824f
C228 B.n159 VSUBS 0.006824f
C229 B.n160 VSUBS 0.006824f
C230 B.n161 VSUBS 0.006824f
C231 B.n162 VSUBS 0.006824f
C232 B.n163 VSUBS 0.006824f
C233 B.n164 VSUBS 0.006824f
C234 B.n165 VSUBS 0.006824f
C235 B.n166 VSUBS 0.006824f
C236 B.n167 VSUBS 0.006824f
C237 B.n168 VSUBS 0.006824f
C238 B.n169 VSUBS 0.006824f
C239 B.n170 VSUBS 0.006824f
C240 B.n171 VSUBS 0.006824f
C241 B.n172 VSUBS 0.006824f
C242 B.n173 VSUBS 0.006824f
C243 B.n174 VSUBS 0.006824f
C244 B.n175 VSUBS 0.006824f
C245 B.n176 VSUBS 0.006824f
C246 B.n177 VSUBS 0.006824f
C247 B.n178 VSUBS 0.006824f
C248 B.n179 VSUBS 0.006824f
C249 B.n180 VSUBS 0.006824f
C250 B.n181 VSUBS 0.006824f
C251 B.n182 VSUBS 0.006824f
C252 B.n183 VSUBS 0.006824f
C253 B.n184 VSUBS 0.006824f
C254 B.n185 VSUBS 0.006824f
C255 B.n186 VSUBS 0.006824f
C256 B.n187 VSUBS 0.006824f
C257 B.n188 VSUBS 0.006824f
C258 B.n189 VSUBS 0.006824f
C259 B.n190 VSUBS 0.006824f
C260 B.n191 VSUBS 0.006824f
C261 B.n192 VSUBS 0.006824f
C262 B.n193 VSUBS 0.006824f
C263 B.n194 VSUBS 0.006824f
C264 B.n195 VSUBS 0.006824f
C265 B.n196 VSUBS 0.006824f
C266 B.n197 VSUBS 0.006824f
C267 B.n198 VSUBS 0.006824f
C268 B.n199 VSUBS 0.006824f
C269 B.n200 VSUBS 0.006824f
C270 B.n201 VSUBS 0.006824f
C271 B.n202 VSUBS 0.006824f
C272 B.n203 VSUBS 0.006824f
C273 B.n204 VSUBS 0.006824f
C274 B.n205 VSUBS 0.006824f
C275 B.n206 VSUBS 0.006824f
C276 B.n207 VSUBS 0.006824f
C277 B.n208 VSUBS 0.006824f
C278 B.n209 VSUBS 0.006824f
C279 B.n210 VSUBS 0.006824f
C280 B.n211 VSUBS 0.006824f
C281 B.n212 VSUBS 0.006824f
C282 B.n213 VSUBS 0.006824f
C283 B.n214 VSUBS 0.006824f
C284 B.n215 VSUBS 0.006824f
C285 B.n216 VSUBS 0.006824f
C286 B.n217 VSUBS 0.006824f
C287 B.n218 VSUBS 0.006824f
C288 B.n219 VSUBS 0.006824f
C289 B.n220 VSUBS 0.006824f
C290 B.n221 VSUBS 0.006824f
C291 B.n222 VSUBS 0.006824f
C292 B.n223 VSUBS 0.006824f
C293 B.n224 VSUBS 0.006824f
C294 B.n225 VSUBS 0.006824f
C295 B.n226 VSUBS 0.01699f
C296 B.n227 VSUBS 0.01699f
C297 B.n228 VSUBS 0.017532f
C298 B.n229 VSUBS 0.006824f
C299 B.n230 VSUBS 0.006824f
C300 B.n231 VSUBS 0.006824f
C301 B.n232 VSUBS 0.006824f
C302 B.n233 VSUBS 0.006824f
C303 B.n234 VSUBS 0.006824f
C304 B.n235 VSUBS 0.006824f
C305 B.n236 VSUBS 0.006824f
C306 B.n237 VSUBS 0.006824f
C307 B.n238 VSUBS 0.006824f
C308 B.n239 VSUBS 0.006824f
C309 B.n240 VSUBS 0.006824f
C310 B.n241 VSUBS 0.006824f
C311 B.n242 VSUBS 0.006824f
C312 B.n243 VSUBS 0.006824f
C313 B.n244 VSUBS 0.006824f
C314 B.n245 VSUBS 0.006824f
C315 B.n246 VSUBS 0.006824f
C316 B.n247 VSUBS 0.006824f
C317 B.n248 VSUBS 0.006824f
C318 B.n249 VSUBS 0.006824f
C319 B.n250 VSUBS 0.006824f
C320 B.n251 VSUBS 0.006824f
C321 B.n252 VSUBS 0.006824f
C322 B.n253 VSUBS 0.006824f
C323 B.n254 VSUBS 0.006824f
C324 B.n255 VSUBS 0.006824f
C325 B.n256 VSUBS 0.006824f
C326 B.n257 VSUBS 0.006824f
C327 B.n258 VSUBS 0.006824f
C328 B.n259 VSUBS 0.006824f
C329 B.n260 VSUBS 0.006824f
C330 B.n261 VSUBS 0.006824f
C331 B.n262 VSUBS 0.006824f
C332 B.n263 VSUBS 0.006824f
C333 B.n264 VSUBS 0.006824f
C334 B.n265 VSUBS 0.006824f
C335 B.n266 VSUBS 0.006824f
C336 B.n267 VSUBS 0.006824f
C337 B.n268 VSUBS 0.006824f
C338 B.n269 VSUBS 0.006824f
C339 B.n270 VSUBS 0.006824f
C340 B.n271 VSUBS 0.006824f
C341 B.n272 VSUBS 0.006824f
C342 B.n273 VSUBS 0.006824f
C343 B.n274 VSUBS 0.006824f
C344 B.n275 VSUBS 0.006824f
C345 B.n276 VSUBS 0.006824f
C346 B.n277 VSUBS 0.006423f
C347 B.n278 VSUBS 0.006824f
C348 B.n279 VSUBS 0.006824f
C349 B.n280 VSUBS 0.003814f
C350 B.n281 VSUBS 0.006824f
C351 B.n282 VSUBS 0.006824f
C352 B.n283 VSUBS 0.006824f
C353 B.n284 VSUBS 0.006824f
C354 B.n285 VSUBS 0.006824f
C355 B.n286 VSUBS 0.006824f
C356 B.n287 VSUBS 0.006824f
C357 B.n288 VSUBS 0.006824f
C358 B.n289 VSUBS 0.006824f
C359 B.n290 VSUBS 0.006824f
C360 B.n291 VSUBS 0.006824f
C361 B.n292 VSUBS 0.006824f
C362 B.n293 VSUBS 0.003814f
C363 B.n294 VSUBS 0.015811f
C364 B.n295 VSUBS 0.006423f
C365 B.n296 VSUBS 0.006824f
C366 B.n297 VSUBS 0.006824f
C367 B.n298 VSUBS 0.006824f
C368 B.n299 VSUBS 0.006824f
C369 B.n300 VSUBS 0.006824f
C370 B.n301 VSUBS 0.006824f
C371 B.n302 VSUBS 0.006824f
C372 B.n303 VSUBS 0.006824f
C373 B.n304 VSUBS 0.006824f
C374 B.n305 VSUBS 0.006824f
C375 B.n306 VSUBS 0.006824f
C376 B.n307 VSUBS 0.006824f
C377 B.n308 VSUBS 0.006824f
C378 B.n309 VSUBS 0.006824f
C379 B.n310 VSUBS 0.006824f
C380 B.n311 VSUBS 0.006824f
C381 B.n312 VSUBS 0.006824f
C382 B.n313 VSUBS 0.006824f
C383 B.n314 VSUBS 0.006824f
C384 B.n315 VSUBS 0.006824f
C385 B.n316 VSUBS 0.006824f
C386 B.n317 VSUBS 0.006824f
C387 B.n318 VSUBS 0.006824f
C388 B.n319 VSUBS 0.006824f
C389 B.n320 VSUBS 0.006824f
C390 B.n321 VSUBS 0.006824f
C391 B.n322 VSUBS 0.006824f
C392 B.n323 VSUBS 0.006824f
C393 B.n324 VSUBS 0.006824f
C394 B.n325 VSUBS 0.006824f
C395 B.n326 VSUBS 0.006824f
C396 B.n327 VSUBS 0.006824f
C397 B.n328 VSUBS 0.006824f
C398 B.n329 VSUBS 0.006824f
C399 B.n330 VSUBS 0.006824f
C400 B.n331 VSUBS 0.006824f
C401 B.n332 VSUBS 0.006824f
C402 B.n333 VSUBS 0.006824f
C403 B.n334 VSUBS 0.006824f
C404 B.n335 VSUBS 0.006824f
C405 B.n336 VSUBS 0.006824f
C406 B.n337 VSUBS 0.006824f
C407 B.n338 VSUBS 0.006824f
C408 B.n339 VSUBS 0.006824f
C409 B.n340 VSUBS 0.006824f
C410 B.n341 VSUBS 0.006824f
C411 B.n342 VSUBS 0.006824f
C412 B.n343 VSUBS 0.006824f
C413 B.n344 VSUBS 0.006824f
C414 B.n345 VSUBS 0.017532f
C415 B.n346 VSUBS 0.01699f
C416 B.n347 VSUBS 0.01699f
C417 B.n348 VSUBS 0.006824f
C418 B.n349 VSUBS 0.006824f
C419 B.n350 VSUBS 0.006824f
C420 B.n351 VSUBS 0.006824f
C421 B.n352 VSUBS 0.006824f
C422 B.n353 VSUBS 0.006824f
C423 B.n354 VSUBS 0.006824f
C424 B.n355 VSUBS 0.006824f
C425 B.n356 VSUBS 0.006824f
C426 B.n357 VSUBS 0.006824f
C427 B.n358 VSUBS 0.006824f
C428 B.n359 VSUBS 0.006824f
C429 B.n360 VSUBS 0.006824f
C430 B.n361 VSUBS 0.006824f
C431 B.n362 VSUBS 0.006824f
C432 B.n363 VSUBS 0.006824f
C433 B.n364 VSUBS 0.006824f
C434 B.n365 VSUBS 0.006824f
C435 B.n366 VSUBS 0.006824f
C436 B.n367 VSUBS 0.006824f
C437 B.n368 VSUBS 0.006824f
C438 B.n369 VSUBS 0.006824f
C439 B.n370 VSUBS 0.006824f
C440 B.n371 VSUBS 0.006824f
C441 B.n372 VSUBS 0.006824f
C442 B.n373 VSUBS 0.006824f
C443 B.n374 VSUBS 0.006824f
C444 B.n375 VSUBS 0.006824f
C445 B.n376 VSUBS 0.006824f
C446 B.n377 VSUBS 0.006824f
C447 B.n378 VSUBS 0.006824f
C448 B.n379 VSUBS 0.006824f
C449 B.n380 VSUBS 0.006824f
C450 B.n381 VSUBS 0.006824f
C451 B.n382 VSUBS 0.006824f
C452 B.n383 VSUBS 0.006824f
C453 B.n384 VSUBS 0.006824f
C454 B.n385 VSUBS 0.006824f
C455 B.n386 VSUBS 0.006824f
C456 B.n387 VSUBS 0.006824f
C457 B.n388 VSUBS 0.006824f
C458 B.n389 VSUBS 0.006824f
C459 B.n390 VSUBS 0.006824f
C460 B.n391 VSUBS 0.006824f
C461 B.n392 VSUBS 0.006824f
C462 B.n393 VSUBS 0.006824f
C463 B.n394 VSUBS 0.006824f
C464 B.n395 VSUBS 0.006824f
C465 B.n396 VSUBS 0.006824f
C466 B.n397 VSUBS 0.006824f
C467 B.n398 VSUBS 0.006824f
C468 B.n399 VSUBS 0.006824f
C469 B.n400 VSUBS 0.006824f
C470 B.n401 VSUBS 0.006824f
C471 B.n402 VSUBS 0.006824f
C472 B.n403 VSUBS 0.006824f
C473 B.n404 VSUBS 0.006824f
C474 B.n405 VSUBS 0.006824f
C475 B.n406 VSUBS 0.006824f
C476 B.n407 VSUBS 0.006824f
C477 B.n408 VSUBS 0.006824f
C478 B.n409 VSUBS 0.006824f
C479 B.n410 VSUBS 0.006824f
C480 B.n411 VSUBS 0.006824f
C481 B.n412 VSUBS 0.006824f
C482 B.n413 VSUBS 0.006824f
C483 B.n414 VSUBS 0.006824f
C484 B.n415 VSUBS 0.006824f
C485 B.n416 VSUBS 0.006824f
C486 B.n417 VSUBS 0.006824f
C487 B.n418 VSUBS 0.006824f
C488 B.n419 VSUBS 0.006824f
C489 B.n420 VSUBS 0.006824f
C490 B.n421 VSUBS 0.006824f
C491 B.n422 VSUBS 0.006824f
C492 B.n423 VSUBS 0.006824f
C493 B.n424 VSUBS 0.006824f
C494 B.n425 VSUBS 0.006824f
C495 B.n426 VSUBS 0.006824f
C496 B.n427 VSUBS 0.006824f
C497 B.n428 VSUBS 0.006824f
C498 B.n429 VSUBS 0.006824f
C499 B.n430 VSUBS 0.006824f
C500 B.n431 VSUBS 0.006824f
C501 B.n432 VSUBS 0.006824f
C502 B.n433 VSUBS 0.006824f
C503 B.n434 VSUBS 0.006824f
C504 B.n435 VSUBS 0.006824f
C505 B.n436 VSUBS 0.006824f
C506 B.n437 VSUBS 0.006824f
C507 B.n438 VSUBS 0.006824f
C508 B.n439 VSUBS 0.006824f
C509 B.n440 VSUBS 0.006824f
C510 B.n441 VSUBS 0.006824f
C511 B.n442 VSUBS 0.006824f
C512 B.n443 VSUBS 0.006824f
C513 B.n444 VSUBS 0.006824f
C514 B.n445 VSUBS 0.006824f
C515 B.n446 VSUBS 0.006824f
C516 B.n447 VSUBS 0.006824f
C517 B.n448 VSUBS 0.006824f
C518 B.n449 VSUBS 0.006824f
C519 B.n450 VSUBS 0.006824f
C520 B.n451 VSUBS 0.006824f
C521 B.n452 VSUBS 0.006824f
C522 B.n453 VSUBS 0.006824f
C523 B.n454 VSUBS 0.006824f
C524 B.n455 VSUBS 0.006824f
C525 B.n456 VSUBS 0.006824f
C526 B.n457 VSUBS 0.006824f
C527 B.n458 VSUBS 0.006824f
C528 B.n459 VSUBS 0.006824f
C529 B.n460 VSUBS 0.006824f
C530 B.n461 VSUBS 0.006824f
C531 B.n462 VSUBS 0.006824f
C532 B.n463 VSUBS 0.006824f
C533 B.n464 VSUBS 0.006824f
C534 B.n465 VSUBS 0.006824f
C535 B.n466 VSUBS 0.01699f
C536 B.n467 VSUBS 0.017708f
C537 B.n468 VSUBS 0.016815f
C538 B.n469 VSUBS 0.006824f
C539 B.n470 VSUBS 0.006824f
C540 B.n471 VSUBS 0.006824f
C541 B.n472 VSUBS 0.006824f
C542 B.n473 VSUBS 0.006824f
C543 B.n474 VSUBS 0.006824f
C544 B.n475 VSUBS 0.006824f
C545 B.n476 VSUBS 0.006824f
C546 B.n477 VSUBS 0.006824f
C547 B.n478 VSUBS 0.006824f
C548 B.n479 VSUBS 0.006824f
C549 B.n480 VSUBS 0.006824f
C550 B.n481 VSUBS 0.006824f
C551 B.n482 VSUBS 0.006824f
C552 B.n483 VSUBS 0.006824f
C553 B.n484 VSUBS 0.006824f
C554 B.n485 VSUBS 0.006824f
C555 B.n486 VSUBS 0.006824f
C556 B.n487 VSUBS 0.006824f
C557 B.n488 VSUBS 0.006824f
C558 B.n489 VSUBS 0.006824f
C559 B.n490 VSUBS 0.006824f
C560 B.n491 VSUBS 0.006824f
C561 B.n492 VSUBS 0.006824f
C562 B.n493 VSUBS 0.006824f
C563 B.n494 VSUBS 0.006824f
C564 B.n495 VSUBS 0.006824f
C565 B.n496 VSUBS 0.006824f
C566 B.n497 VSUBS 0.006824f
C567 B.n498 VSUBS 0.006824f
C568 B.n499 VSUBS 0.006824f
C569 B.n500 VSUBS 0.006824f
C570 B.n501 VSUBS 0.006824f
C571 B.n502 VSUBS 0.006824f
C572 B.n503 VSUBS 0.006824f
C573 B.n504 VSUBS 0.006824f
C574 B.n505 VSUBS 0.006824f
C575 B.n506 VSUBS 0.006824f
C576 B.n507 VSUBS 0.006824f
C577 B.n508 VSUBS 0.006824f
C578 B.n509 VSUBS 0.006824f
C579 B.n510 VSUBS 0.006824f
C580 B.n511 VSUBS 0.006824f
C581 B.n512 VSUBS 0.006824f
C582 B.n513 VSUBS 0.006824f
C583 B.n514 VSUBS 0.006824f
C584 B.n515 VSUBS 0.006824f
C585 B.n516 VSUBS 0.006824f
C586 B.n517 VSUBS 0.006423f
C587 B.n518 VSUBS 0.006824f
C588 B.n519 VSUBS 0.006824f
C589 B.n520 VSUBS 0.003814f
C590 B.n521 VSUBS 0.006824f
C591 B.n522 VSUBS 0.006824f
C592 B.n523 VSUBS 0.006824f
C593 B.n524 VSUBS 0.006824f
C594 B.n525 VSUBS 0.006824f
C595 B.n526 VSUBS 0.006824f
C596 B.n527 VSUBS 0.006824f
C597 B.n528 VSUBS 0.006824f
C598 B.n529 VSUBS 0.006824f
C599 B.n530 VSUBS 0.006824f
C600 B.n531 VSUBS 0.006824f
C601 B.n532 VSUBS 0.006824f
C602 B.n533 VSUBS 0.003814f
C603 B.n534 VSUBS 0.015811f
C604 B.n535 VSUBS 0.006423f
C605 B.n536 VSUBS 0.006824f
C606 B.n537 VSUBS 0.006824f
C607 B.n538 VSUBS 0.006824f
C608 B.n539 VSUBS 0.006824f
C609 B.n540 VSUBS 0.006824f
C610 B.n541 VSUBS 0.006824f
C611 B.n542 VSUBS 0.006824f
C612 B.n543 VSUBS 0.006824f
C613 B.n544 VSUBS 0.006824f
C614 B.n545 VSUBS 0.006824f
C615 B.n546 VSUBS 0.006824f
C616 B.n547 VSUBS 0.006824f
C617 B.n548 VSUBS 0.006824f
C618 B.n549 VSUBS 0.006824f
C619 B.n550 VSUBS 0.006824f
C620 B.n551 VSUBS 0.006824f
C621 B.n552 VSUBS 0.006824f
C622 B.n553 VSUBS 0.006824f
C623 B.n554 VSUBS 0.006824f
C624 B.n555 VSUBS 0.006824f
C625 B.n556 VSUBS 0.006824f
C626 B.n557 VSUBS 0.006824f
C627 B.n558 VSUBS 0.006824f
C628 B.n559 VSUBS 0.006824f
C629 B.n560 VSUBS 0.006824f
C630 B.n561 VSUBS 0.006824f
C631 B.n562 VSUBS 0.006824f
C632 B.n563 VSUBS 0.006824f
C633 B.n564 VSUBS 0.006824f
C634 B.n565 VSUBS 0.006824f
C635 B.n566 VSUBS 0.006824f
C636 B.n567 VSUBS 0.006824f
C637 B.n568 VSUBS 0.006824f
C638 B.n569 VSUBS 0.006824f
C639 B.n570 VSUBS 0.006824f
C640 B.n571 VSUBS 0.006824f
C641 B.n572 VSUBS 0.006824f
C642 B.n573 VSUBS 0.006824f
C643 B.n574 VSUBS 0.006824f
C644 B.n575 VSUBS 0.006824f
C645 B.n576 VSUBS 0.006824f
C646 B.n577 VSUBS 0.006824f
C647 B.n578 VSUBS 0.006824f
C648 B.n579 VSUBS 0.006824f
C649 B.n580 VSUBS 0.006824f
C650 B.n581 VSUBS 0.006824f
C651 B.n582 VSUBS 0.006824f
C652 B.n583 VSUBS 0.006824f
C653 B.n584 VSUBS 0.006824f
C654 B.n585 VSUBS 0.017532f
C655 B.n586 VSUBS 0.01699f
C656 B.n587 VSUBS 0.01699f
C657 B.n588 VSUBS 0.006824f
C658 B.n589 VSUBS 0.006824f
C659 B.n590 VSUBS 0.006824f
C660 B.n591 VSUBS 0.006824f
C661 B.n592 VSUBS 0.006824f
C662 B.n593 VSUBS 0.006824f
C663 B.n594 VSUBS 0.006824f
C664 B.n595 VSUBS 0.006824f
C665 B.n596 VSUBS 0.006824f
C666 B.n597 VSUBS 0.006824f
C667 B.n598 VSUBS 0.006824f
C668 B.n599 VSUBS 0.006824f
C669 B.n600 VSUBS 0.006824f
C670 B.n601 VSUBS 0.006824f
C671 B.n602 VSUBS 0.006824f
C672 B.n603 VSUBS 0.006824f
C673 B.n604 VSUBS 0.006824f
C674 B.n605 VSUBS 0.006824f
C675 B.n606 VSUBS 0.006824f
C676 B.n607 VSUBS 0.006824f
C677 B.n608 VSUBS 0.006824f
C678 B.n609 VSUBS 0.006824f
C679 B.n610 VSUBS 0.006824f
C680 B.n611 VSUBS 0.006824f
C681 B.n612 VSUBS 0.006824f
C682 B.n613 VSUBS 0.006824f
C683 B.n614 VSUBS 0.006824f
C684 B.n615 VSUBS 0.006824f
C685 B.n616 VSUBS 0.006824f
C686 B.n617 VSUBS 0.006824f
C687 B.n618 VSUBS 0.006824f
C688 B.n619 VSUBS 0.006824f
C689 B.n620 VSUBS 0.006824f
C690 B.n621 VSUBS 0.006824f
C691 B.n622 VSUBS 0.006824f
C692 B.n623 VSUBS 0.006824f
C693 B.n624 VSUBS 0.006824f
C694 B.n625 VSUBS 0.006824f
C695 B.n626 VSUBS 0.006824f
C696 B.n627 VSUBS 0.006824f
C697 B.n628 VSUBS 0.006824f
C698 B.n629 VSUBS 0.006824f
C699 B.n630 VSUBS 0.006824f
C700 B.n631 VSUBS 0.006824f
C701 B.n632 VSUBS 0.006824f
C702 B.n633 VSUBS 0.006824f
C703 B.n634 VSUBS 0.006824f
C704 B.n635 VSUBS 0.006824f
C705 B.n636 VSUBS 0.006824f
C706 B.n637 VSUBS 0.006824f
C707 B.n638 VSUBS 0.006824f
C708 B.n639 VSUBS 0.006824f
C709 B.n640 VSUBS 0.006824f
C710 B.n641 VSUBS 0.006824f
C711 B.n642 VSUBS 0.006824f
C712 B.n643 VSUBS 0.006824f
C713 B.n644 VSUBS 0.006824f
C714 B.n645 VSUBS 0.006824f
C715 B.n646 VSUBS 0.006824f
C716 B.n647 VSUBS 0.015452f
C717 VDD2.t0 VSUBS 0.206976f
C718 VDD2.t3 VSUBS 0.206976f
C719 VDD2.n0 VSUBS 2.19398f
C720 VDD2.t1 VSUBS 0.206976f
C721 VDD2.t2 VSUBS 0.206976f
C722 VDD2.n1 VSUBS 1.54748f
C723 VDD2.n2 VSUBS 4.24877f
C724 VTAIL.t6 VSUBS 1.73769f
C725 VTAIL.n0 VSUBS 0.799618f
C726 VTAIL.t1 VSUBS 1.73769f
C727 VTAIL.n1 VSUBS 0.922156f
C728 VTAIL.t0 VSUBS 1.73769f
C729 VTAIL.n2 VSUBS 2.15246f
C730 VTAIL.t3 VSUBS 1.73771f
C731 VTAIL.n3 VSUBS 2.15245f
C732 VTAIL.t5 VSUBS 1.73771f
C733 VTAIL.n4 VSUBS 0.922143f
C734 VTAIL.t2 VSUBS 1.73771f
C735 VTAIL.n5 VSUBS 0.922143f
C736 VTAIL.t7 VSUBS 1.73769f
C737 VTAIL.n6 VSUBS 2.15246f
C738 VTAIL.t4 VSUBS 1.73769f
C739 VTAIL.n7 VSUBS 2.02045f
C740 VN.t0 VSUBS 3.03667f
C741 VN.t3 VSUBS 3.04877f
C742 VN.n0 VSUBS 1.82362f
C743 VN.t2 VSUBS 3.03667f
C744 VN.t1 VSUBS 3.04877f
C745 VN.n1 VSUBS 3.65545f
.ends

