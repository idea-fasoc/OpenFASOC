* NGSPICE file created from diff_pair_sample_0370.ext - technology: sky130A

.subckt diff_pair_sample_0370 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3.14
X1 VTAIL.t2 VN.t0 VDD2.t3 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3.14
X2 VTAIL.t0 VN.t1 VDD2.t2 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3.14
X3 B.t11 B.t9 B.t10 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3.14
X4 VDD2.t1 VN.t2 VTAIL.t1 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3.14
X5 VDD1.t2 VP.t1 VTAIL.t4 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3.14
X6 VDD2.t0 VN.t3 VTAIL.t3 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3.14
X7 VTAIL.t6 VP.t2 VDD1.t1 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3.14
X8 B.t8 B.t6 B.t7 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3.14
X9 VTAIL.t7 VP.t3 VDD1.t0 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3.14
X10 B.t5 B.t3 B.t4 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3.14
X11 B.t2 B.t0 B.t1 w_n3052_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3.14
R0 VP.n15 VP.n14 161.3
R1 VP.n13 VP.n1 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n2 161.3
R4 VP.n9 VP.n8 161.3
R5 VP.n7 VP.n3 161.3
R6 VP.n4 VP.t2 104.742
R7 VP.n4 VP.t0 103.718
R8 VP.n6 VP.t3 70.2282
R9 VP.n0 VP.t1 70.2282
R10 VP.n6 VP.n5 66.3344
R11 VP.n16 VP.n0 66.3344
R12 VP.n12 VP.n2 56.5193
R13 VP.n5 VP.n4 48.7133
R14 VP.n8 VP.n7 24.4675
R15 VP.n8 VP.n2 24.4675
R16 VP.n13 VP.n12 24.4675
R17 VP.n14 VP.n13 24.4675
R18 VP.n7 VP.n6 23.7335
R19 VP.n14 VP.n0 23.7335
R20 VP.n5 VP.n3 0.354971
R21 VP.n16 VP.n15 0.354971
R22 VP VP.n16 0.26696
R23 VP.n9 VP.n3 0.189894
R24 VP.n10 VP.n9 0.189894
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n1 0.189894
R27 VP.n15 VP.n1 0.189894
R28 VTAIL.n6 VTAIL.t5 64.9254
R29 VTAIL.n5 VTAIL.t6 64.9254
R30 VTAIL.n4 VTAIL.t3 64.9254
R31 VTAIL.n3 VTAIL.t0 64.9254
R32 VTAIL.n7 VTAIL.t1 64.9252
R33 VTAIL.n0 VTAIL.t2 64.9252
R34 VTAIL.n1 VTAIL.t4 64.9252
R35 VTAIL.n2 VTAIL.t7 64.9252
R36 VTAIL.n7 VTAIL.n6 23.2462
R37 VTAIL.n3 VTAIL.n2 23.2462
R38 VTAIL.n4 VTAIL.n3 2.99188
R39 VTAIL.n6 VTAIL.n5 2.99188
R40 VTAIL.n2 VTAIL.n1 2.99188
R41 VTAIL VTAIL.n0 1.55438
R42 VTAIL VTAIL.n7 1.438
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 VDD1 VDD1.n1 119.153
R46 VDD1 VDD1.n0 78.1099
R47 VDD1.n0 VDD1.t1 3.55296
R48 VDD1.n0 VDD1.t3 3.55296
R49 VDD1.n1 VDD1.t0 3.55296
R50 VDD1.n1 VDD1.t2 3.55296
R51 VN.n1 VN.t3 104.742
R52 VN.n0 VN.t0 104.742
R53 VN.n0 VN.t2 103.718
R54 VN.n1 VN.t1 103.718
R55 VN VN.n1 48.8787
R56 VN VN.n0 2.76127
R57 VDD2.n2 VDD2.n0 118.629
R58 VDD2.n2 VDD2.n1 78.0517
R59 VDD2.n1 VDD2.t2 3.55296
R60 VDD2.n1 VDD2.t0 3.55296
R61 VDD2.n0 VDD2.t3 3.55296
R62 VDD2.n0 VDD2.t1 3.55296
R63 VDD2 VDD2.n2 0.0586897
R64 B.n334 B.n103 585
R65 B.n333 B.n332 585
R66 B.n331 B.n104 585
R67 B.n330 B.n329 585
R68 B.n328 B.n105 585
R69 B.n327 B.n326 585
R70 B.n325 B.n106 585
R71 B.n324 B.n323 585
R72 B.n322 B.n107 585
R73 B.n321 B.n320 585
R74 B.n319 B.n108 585
R75 B.n318 B.n317 585
R76 B.n316 B.n109 585
R77 B.n315 B.n314 585
R78 B.n313 B.n110 585
R79 B.n312 B.n311 585
R80 B.n310 B.n111 585
R81 B.n309 B.n308 585
R82 B.n307 B.n112 585
R83 B.n306 B.n305 585
R84 B.n304 B.n113 585
R85 B.n303 B.n302 585
R86 B.n301 B.n114 585
R87 B.n300 B.n299 585
R88 B.n298 B.n115 585
R89 B.n297 B.n296 585
R90 B.n295 B.n116 585
R91 B.n294 B.n293 585
R92 B.n292 B.n117 585
R93 B.n291 B.n290 585
R94 B.n289 B.n118 585
R95 B.n288 B.n287 585
R96 B.n286 B.n119 585
R97 B.n285 B.n284 585
R98 B.n280 B.n120 585
R99 B.n279 B.n278 585
R100 B.n277 B.n121 585
R101 B.n276 B.n275 585
R102 B.n274 B.n122 585
R103 B.n273 B.n272 585
R104 B.n271 B.n123 585
R105 B.n270 B.n269 585
R106 B.n268 B.n124 585
R107 B.n266 B.n265 585
R108 B.n264 B.n127 585
R109 B.n263 B.n262 585
R110 B.n261 B.n128 585
R111 B.n260 B.n259 585
R112 B.n258 B.n129 585
R113 B.n257 B.n256 585
R114 B.n255 B.n130 585
R115 B.n254 B.n253 585
R116 B.n252 B.n131 585
R117 B.n251 B.n250 585
R118 B.n249 B.n132 585
R119 B.n248 B.n247 585
R120 B.n246 B.n133 585
R121 B.n245 B.n244 585
R122 B.n243 B.n134 585
R123 B.n242 B.n241 585
R124 B.n240 B.n135 585
R125 B.n239 B.n238 585
R126 B.n237 B.n136 585
R127 B.n236 B.n235 585
R128 B.n234 B.n137 585
R129 B.n233 B.n232 585
R130 B.n231 B.n138 585
R131 B.n230 B.n229 585
R132 B.n228 B.n139 585
R133 B.n227 B.n226 585
R134 B.n225 B.n140 585
R135 B.n224 B.n223 585
R136 B.n222 B.n141 585
R137 B.n221 B.n220 585
R138 B.n219 B.n142 585
R139 B.n218 B.n217 585
R140 B.n336 B.n335 585
R141 B.n337 B.n102 585
R142 B.n339 B.n338 585
R143 B.n340 B.n101 585
R144 B.n342 B.n341 585
R145 B.n343 B.n100 585
R146 B.n345 B.n344 585
R147 B.n346 B.n99 585
R148 B.n348 B.n347 585
R149 B.n349 B.n98 585
R150 B.n351 B.n350 585
R151 B.n352 B.n97 585
R152 B.n354 B.n353 585
R153 B.n355 B.n96 585
R154 B.n357 B.n356 585
R155 B.n358 B.n95 585
R156 B.n360 B.n359 585
R157 B.n361 B.n94 585
R158 B.n363 B.n362 585
R159 B.n364 B.n93 585
R160 B.n366 B.n365 585
R161 B.n367 B.n92 585
R162 B.n369 B.n368 585
R163 B.n370 B.n91 585
R164 B.n372 B.n371 585
R165 B.n373 B.n90 585
R166 B.n375 B.n374 585
R167 B.n376 B.n89 585
R168 B.n378 B.n377 585
R169 B.n379 B.n88 585
R170 B.n381 B.n380 585
R171 B.n382 B.n87 585
R172 B.n384 B.n383 585
R173 B.n385 B.n86 585
R174 B.n387 B.n386 585
R175 B.n388 B.n85 585
R176 B.n390 B.n389 585
R177 B.n391 B.n84 585
R178 B.n393 B.n392 585
R179 B.n394 B.n83 585
R180 B.n396 B.n395 585
R181 B.n397 B.n82 585
R182 B.n399 B.n398 585
R183 B.n400 B.n81 585
R184 B.n402 B.n401 585
R185 B.n403 B.n80 585
R186 B.n405 B.n404 585
R187 B.n406 B.n79 585
R188 B.n408 B.n407 585
R189 B.n409 B.n78 585
R190 B.n411 B.n410 585
R191 B.n412 B.n77 585
R192 B.n414 B.n413 585
R193 B.n415 B.n76 585
R194 B.n417 B.n416 585
R195 B.n418 B.n75 585
R196 B.n420 B.n419 585
R197 B.n421 B.n74 585
R198 B.n423 B.n422 585
R199 B.n424 B.n73 585
R200 B.n426 B.n425 585
R201 B.n427 B.n72 585
R202 B.n429 B.n428 585
R203 B.n430 B.n71 585
R204 B.n432 B.n431 585
R205 B.n433 B.n70 585
R206 B.n435 B.n434 585
R207 B.n436 B.n69 585
R208 B.n438 B.n437 585
R209 B.n439 B.n68 585
R210 B.n441 B.n440 585
R211 B.n442 B.n67 585
R212 B.n444 B.n443 585
R213 B.n445 B.n66 585
R214 B.n447 B.n446 585
R215 B.n448 B.n65 585
R216 B.n450 B.n449 585
R217 B.n451 B.n64 585
R218 B.n566 B.n21 585
R219 B.n565 B.n564 585
R220 B.n563 B.n22 585
R221 B.n562 B.n561 585
R222 B.n560 B.n23 585
R223 B.n559 B.n558 585
R224 B.n557 B.n24 585
R225 B.n556 B.n555 585
R226 B.n554 B.n25 585
R227 B.n553 B.n552 585
R228 B.n551 B.n26 585
R229 B.n550 B.n549 585
R230 B.n548 B.n27 585
R231 B.n547 B.n546 585
R232 B.n545 B.n28 585
R233 B.n544 B.n543 585
R234 B.n542 B.n29 585
R235 B.n541 B.n540 585
R236 B.n539 B.n30 585
R237 B.n538 B.n537 585
R238 B.n536 B.n31 585
R239 B.n535 B.n534 585
R240 B.n533 B.n32 585
R241 B.n532 B.n531 585
R242 B.n530 B.n33 585
R243 B.n529 B.n528 585
R244 B.n527 B.n34 585
R245 B.n526 B.n525 585
R246 B.n524 B.n35 585
R247 B.n523 B.n522 585
R248 B.n521 B.n36 585
R249 B.n520 B.n519 585
R250 B.n518 B.n37 585
R251 B.n516 B.n515 585
R252 B.n514 B.n40 585
R253 B.n513 B.n512 585
R254 B.n511 B.n41 585
R255 B.n510 B.n509 585
R256 B.n508 B.n42 585
R257 B.n507 B.n506 585
R258 B.n505 B.n43 585
R259 B.n504 B.n503 585
R260 B.n502 B.n44 585
R261 B.n501 B.n500 585
R262 B.n499 B.n45 585
R263 B.n498 B.n497 585
R264 B.n496 B.n49 585
R265 B.n495 B.n494 585
R266 B.n493 B.n50 585
R267 B.n492 B.n491 585
R268 B.n490 B.n51 585
R269 B.n489 B.n488 585
R270 B.n487 B.n52 585
R271 B.n486 B.n485 585
R272 B.n484 B.n53 585
R273 B.n483 B.n482 585
R274 B.n481 B.n54 585
R275 B.n480 B.n479 585
R276 B.n478 B.n55 585
R277 B.n477 B.n476 585
R278 B.n475 B.n56 585
R279 B.n474 B.n473 585
R280 B.n472 B.n57 585
R281 B.n471 B.n470 585
R282 B.n469 B.n58 585
R283 B.n468 B.n467 585
R284 B.n466 B.n59 585
R285 B.n465 B.n464 585
R286 B.n463 B.n60 585
R287 B.n462 B.n461 585
R288 B.n460 B.n61 585
R289 B.n459 B.n458 585
R290 B.n457 B.n62 585
R291 B.n456 B.n455 585
R292 B.n454 B.n63 585
R293 B.n453 B.n452 585
R294 B.n568 B.n567 585
R295 B.n569 B.n20 585
R296 B.n571 B.n570 585
R297 B.n572 B.n19 585
R298 B.n574 B.n573 585
R299 B.n575 B.n18 585
R300 B.n577 B.n576 585
R301 B.n578 B.n17 585
R302 B.n580 B.n579 585
R303 B.n581 B.n16 585
R304 B.n583 B.n582 585
R305 B.n584 B.n15 585
R306 B.n586 B.n585 585
R307 B.n587 B.n14 585
R308 B.n589 B.n588 585
R309 B.n590 B.n13 585
R310 B.n592 B.n591 585
R311 B.n593 B.n12 585
R312 B.n595 B.n594 585
R313 B.n596 B.n11 585
R314 B.n598 B.n597 585
R315 B.n599 B.n10 585
R316 B.n601 B.n600 585
R317 B.n602 B.n9 585
R318 B.n604 B.n603 585
R319 B.n605 B.n8 585
R320 B.n607 B.n606 585
R321 B.n608 B.n7 585
R322 B.n610 B.n609 585
R323 B.n611 B.n6 585
R324 B.n613 B.n612 585
R325 B.n614 B.n5 585
R326 B.n616 B.n615 585
R327 B.n617 B.n4 585
R328 B.n619 B.n618 585
R329 B.n620 B.n3 585
R330 B.n622 B.n621 585
R331 B.n623 B.n0 585
R332 B.n2 B.n1 585
R333 B.n162 B.n161 585
R334 B.n164 B.n163 585
R335 B.n165 B.n160 585
R336 B.n167 B.n166 585
R337 B.n168 B.n159 585
R338 B.n170 B.n169 585
R339 B.n171 B.n158 585
R340 B.n173 B.n172 585
R341 B.n174 B.n157 585
R342 B.n176 B.n175 585
R343 B.n177 B.n156 585
R344 B.n179 B.n178 585
R345 B.n180 B.n155 585
R346 B.n182 B.n181 585
R347 B.n183 B.n154 585
R348 B.n185 B.n184 585
R349 B.n186 B.n153 585
R350 B.n188 B.n187 585
R351 B.n189 B.n152 585
R352 B.n191 B.n190 585
R353 B.n192 B.n151 585
R354 B.n194 B.n193 585
R355 B.n195 B.n150 585
R356 B.n197 B.n196 585
R357 B.n198 B.n149 585
R358 B.n200 B.n199 585
R359 B.n201 B.n148 585
R360 B.n203 B.n202 585
R361 B.n204 B.n147 585
R362 B.n206 B.n205 585
R363 B.n207 B.n146 585
R364 B.n209 B.n208 585
R365 B.n210 B.n145 585
R366 B.n212 B.n211 585
R367 B.n213 B.n144 585
R368 B.n215 B.n214 585
R369 B.n216 B.n143 585
R370 B.n217 B.n216 540.549
R371 B.n335 B.n334 540.549
R372 B.n453 B.n64 540.549
R373 B.n568 B.n21 540.549
R374 B.n125 B.t9 278.966
R375 B.n281 B.t6 278.966
R376 B.n46 B.t0 278.966
R377 B.n38 B.t3 278.966
R378 B.n625 B.n624 256.663
R379 B.n624 B.n623 235.042
R380 B.n624 B.n2 235.042
R381 B.n281 B.t7 181.345
R382 B.n46 B.t2 181.345
R383 B.n125 B.t10 181.333
R384 B.n38 B.t5 181.333
R385 B.n217 B.n142 163.367
R386 B.n221 B.n142 163.367
R387 B.n222 B.n221 163.367
R388 B.n223 B.n222 163.367
R389 B.n223 B.n140 163.367
R390 B.n227 B.n140 163.367
R391 B.n228 B.n227 163.367
R392 B.n229 B.n228 163.367
R393 B.n229 B.n138 163.367
R394 B.n233 B.n138 163.367
R395 B.n234 B.n233 163.367
R396 B.n235 B.n234 163.367
R397 B.n235 B.n136 163.367
R398 B.n239 B.n136 163.367
R399 B.n240 B.n239 163.367
R400 B.n241 B.n240 163.367
R401 B.n241 B.n134 163.367
R402 B.n245 B.n134 163.367
R403 B.n246 B.n245 163.367
R404 B.n247 B.n246 163.367
R405 B.n247 B.n132 163.367
R406 B.n251 B.n132 163.367
R407 B.n252 B.n251 163.367
R408 B.n253 B.n252 163.367
R409 B.n253 B.n130 163.367
R410 B.n257 B.n130 163.367
R411 B.n258 B.n257 163.367
R412 B.n259 B.n258 163.367
R413 B.n259 B.n128 163.367
R414 B.n263 B.n128 163.367
R415 B.n264 B.n263 163.367
R416 B.n265 B.n264 163.367
R417 B.n265 B.n124 163.367
R418 B.n270 B.n124 163.367
R419 B.n271 B.n270 163.367
R420 B.n272 B.n271 163.367
R421 B.n272 B.n122 163.367
R422 B.n276 B.n122 163.367
R423 B.n277 B.n276 163.367
R424 B.n278 B.n277 163.367
R425 B.n278 B.n120 163.367
R426 B.n285 B.n120 163.367
R427 B.n286 B.n285 163.367
R428 B.n287 B.n286 163.367
R429 B.n287 B.n118 163.367
R430 B.n291 B.n118 163.367
R431 B.n292 B.n291 163.367
R432 B.n293 B.n292 163.367
R433 B.n293 B.n116 163.367
R434 B.n297 B.n116 163.367
R435 B.n298 B.n297 163.367
R436 B.n299 B.n298 163.367
R437 B.n299 B.n114 163.367
R438 B.n303 B.n114 163.367
R439 B.n304 B.n303 163.367
R440 B.n305 B.n304 163.367
R441 B.n305 B.n112 163.367
R442 B.n309 B.n112 163.367
R443 B.n310 B.n309 163.367
R444 B.n311 B.n310 163.367
R445 B.n311 B.n110 163.367
R446 B.n315 B.n110 163.367
R447 B.n316 B.n315 163.367
R448 B.n317 B.n316 163.367
R449 B.n317 B.n108 163.367
R450 B.n321 B.n108 163.367
R451 B.n322 B.n321 163.367
R452 B.n323 B.n322 163.367
R453 B.n323 B.n106 163.367
R454 B.n327 B.n106 163.367
R455 B.n328 B.n327 163.367
R456 B.n329 B.n328 163.367
R457 B.n329 B.n104 163.367
R458 B.n333 B.n104 163.367
R459 B.n334 B.n333 163.367
R460 B.n449 B.n64 163.367
R461 B.n449 B.n448 163.367
R462 B.n448 B.n447 163.367
R463 B.n447 B.n66 163.367
R464 B.n443 B.n66 163.367
R465 B.n443 B.n442 163.367
R466 B.n442 B.n441 163.367
R467 B.n441 B.n68 163.367
R468 B.n437 B.n68 163.367
R469 B.n437 B.n436 163.367
R470 B.n436 B.n435 163.367
R471 B.n435 B.n70 163.367
R472 B.n431 B.n70 163.367
R473 B.n431 B.n430 163.367
R474 B.n430 B.n429 163.367
R475 B.n429 B.n72 163.367
R476 B.n425 B.n72 163.367
R477 B.n425 B.n424 163.367
R478 B.n424 B.n423 163.367
R479 B.n423 B.n74 163.367
R480 B.n419 B.n74 163.367
R481 B.n419 B.n418 163.367
R482 B.n418 B.n417 163.367
R483 B.n417 B.n76 163.367
R484 B.n413 B.n76 163.367
R485 B.n413 B.n412 163.367
R486 B.n412 B.n411 163.367
R487 B.n411 B.n78 163.367
R488 B.n407 B.n78 163.367
R489 B.n407 B.n406 163.367
R490 B.n406 B.n405 163.367
R491 B.n405 B.n80 163.367
R492 B.n401 B.n80 163.367
R493 B.n401 B.n400 163.367
R494 B.n400 B.n399 163.367
R495 B.n399 B.n82 163.367
R496 B.n395 B.n82 163.367
R497 B.n395 B.n394 163.367
R498 B.n394 B.n393 163.367
R499 B.n393 B.n84 163.367
R500 B.n389 B.n84 163.367
R501 B.n389 B.n388 163.367
R502 B.n388 B.n387 163.367
R503 B.n387 B.n86 163.367
R504 B.n383 B.n86 163.367
R505 B.n383 B.n382 163.367
R506 B.n382 B.n381 163.367
R507 B.n381 B.n88 163.367
R508 B.n377 B.n88 163.367
R509 B.n377 B.n376 163.367
R510 B.n376 B.n375 163.367
R511 B.n375 B.n90 163.367
R512 B.n371 B.n90 163.367
R513 B.n371 B.n370 163.367
R514 B.n370 B.n369 163.367
R515 B.n369 B.n92 163.367
R516 B.n365 B.n92 163.367
R517 B.n365 B.n364 163.367
R518 B.n364 B.n363 163.367
R519 B.n363 B.n94 163.367
R520 B.n359 B.n94 163.367
R521 B.n359 B.n358 163.367
R522 B.n358 B.n357 163.367
R523 B.n357 B.n96 163.367
R524 B.n353 B.n96 163.367
R525 B.n353 B.n352 163.367
R526 B.n352 B.n351 163.367
R527 B.n351 B.n98 163.367
R528 B.n347 B.n98 163.367
R529 B.n347 B.n346 163.367
R530 B.n346 B.n345 163.367
R531 B.n345 B.n100 163.367
R532 B.n341 B.n100 163.367
R533 B.n341 B.n340 163.367
R534 B.n340 B.n339 163.367
R535 B.n339 B.n102 163.367
R536 B.n335 B.n102 163.367
R537 B.n564 B.n21 163.367
R538 B.n564 B.n563 163.367
R539 B.n563 B.n562 163.367
R540 B.n562 B.n23 163.367
R541 B.n558 B.n23 163.367
R542 B.n558 B.n557 163.367
R543 B.n557 B.n556 163.367
R544 B.n556 B.n25 163.367
R545 B.n552 B.n25 163.367
R546 B.n552 B.n551 163.367
R547 B.n551 B.n550 163.367
R548 B.n550 B.n27 163.367
R549 B.n546 B.n27 163.367
R550 B.n546 B.n545 163.367
R551 B.n545 B.n544 163.367
R552 B.n544 B.n29 163.367
R553 B.n540 B.n29 163.367
R554 B.n540 B.n539 163.367
R555 B.n539 B.n538 163.367
R556 B.n538 B.n31 163.367
R557 B.n534 B.n31 163.367
R558 B.n534 B.n533 163.367
R559 B.n533 B.n532 163.367
R560 B.n532 B.n33 163.367
R561 B.n528 B.n33 163.367
R562 B.n528 B.n527 163.367
R563 B.n527 B.n526 163.367
R564 B.n526 B.n35 163.367
R565 B.n522 B.n35 163.367
R566 B.n522 B.n521 163.367
R567 B.n521 B.n520 163.367
R568 B.n520 B.n37 163.367
R569 B.n515 B.n37 163.367
R570 B.n515 B.n514 163.367
R571 B.n514 B.n513 163.367
R572 B.n513 B.n41 163.367
R573 B.n509 B.n41 163.367
R574 B.n509 B.n508 163.367
R575 B.n508 B.n507 163.367
R576 B.n507 B.n43 163.367
R577 B.n503 B.n43 163.367
R578 B.n503 B.n502 163.367
R579 B.n502 B.n501 163.367
R580 B.n501 B.n45 163.367
R581 B.n497 B.n45 163.367
R582 B.n497 B.n496 163.367
R583 B.n496 B.n495 163.367
R584 B.n495 B.n50 163.367
R585 B.n491 B.n50 163.367
R586 B.n491 B.n490 163.367
R587 B.n490 B.n489 163.367
R588 B.n489 B.n52 163.367
R589 B.n485 B.n52 163.367
R590 B.n485 B.n484 163.367
R591 B.n484 B.n483 163.367
R592 B.n483 B.n54 163.367
R593 B.n479 B.n54 163.367
R594 B.n479 B.n478 163.367
R595 B.n478 B.n477 163.367
R596 B.n477 B.n56 163.367
R597 B.n473 B.n56 163.367
R598 B.n473 B.n472 163.367
R599 B.n472 B.n471 163.367
R600 B.n471 B.n58 163.367
R601 B.n467 B.n58 163.367
R602 B.n467 B.n466 163.367
R603 B.n466 B.n465 163.367
R604 B.n465 B.n60 163.367
R605 B.n461 B.n60 163.367
R606 B.n461 B.n460 163.367
R607 B.n460 B.n459 163.367
R608 B.n459 B.n62 163.367
R609 B.n455 B.n62 163.367
R610 B.n455 B.n454 163.367
R611 B.n454 B.n453 163.367
R612 B.n569 B.n568 163.367
R613 B.n570 B.n569 163.367
R614 B.n570 B.n19 163.367
R615 B.n574 B.n19 163.367
R616 B.n575 B.n574 163.367
R617 B.n576 B.n575 163.367
R618 B.n576 B.n17 163.367
R619 B.n580 B.n17 163.367
R620 B.n581 B.n580 163.367
R621 B.n582 B.n581 163.367
R622 B.n582 B.n15 163.367
R623 B.n586 B.n15 163.367
R624 B.n587 B.n586 163.367
R625 B.n588 B.n587 163.367
R626 B.n588 B.n13 163.367
R627 B.n592 B.n13 163.367
R628 B.n593 B.n592 163.367
R629 B.n594 B.n593 163.367
R630 B.n594 B.n11 163.367
R631 B.n598 B.n11 163.367
R632 B.n599 B.n598 163.367
R633 B.n600 B.n599 163.367
R634 B.n600 B.n9 163.367
R635 B.n604 B.n9 163.367
R636 B.n605 B.n604 163.367
R637 B.n606 B.n605 163.367
R638 B.n606 B.n7 163.367
R639 B.n610 B.n7 163.367
R640 B.n611 B.n610 163.367
R641 B.n612 B.n611 163.367
R642 B.n612 B.n5 163.367
R643 B.n616 B.n5 163.367
R644 B.n617 B.n616 163.367
R645 B.n618 B.n617 163.367
R646 B.n618 B.n3 163.367
R647 B.n622 B.n3 163.367
R648 B.n623 B.n622 163.367
R649 B.n162 B.n2 163.367
R650 B.n163 B.n162 163.367
R651 B.n163 B.n160 163.367
R652 B.n167 B.n160 163.367
R653 B.n168 B.n167 163.367
R654 B.n169 B.n168 163.367
R655 B.n169 B.n158 163.367
R656 B.n173 B.n158 163.367
R657 B.n174 B.n173 163.367
R658 B.n175 B.n174 163.367
R659 B.n175 B.n156 163.367
R660 B.n179 B.n156 163.367
R661 B.n180 B.n179 163.367
R662 B.n181 B.n180 163.367
R663 B.n181 B.n154 163.367
R664 B.n185 B.n154 163.367
R665 B.n186 B.n185 163.367
R666 B.n187 B.n186 163.367
R667 B.n187 B.n152 163.367
R668 B.n191 B.n152 163.367
R669 B.n192 B.n191 163.367
R670 B.n193 B.n192 163.367
R671 B.n193 B.n150 163.367
R672 B.n197 B.n150 163.367
R673 B.n198 B.n197 163.367
R674 B.n199 B.n198 163.367
R675 B.n199 B.n148 163.367
R676 B.n203 B.n148 163.367
R677 B.n204 B.n203 163.367
R678 B.n205 B.n204 163.367
R679 B.n205 B.n146 163.367
R680 B.n209 B.n146 163.367
R681 B.n210 B.n209 163.367
R682 B.n211 B.n210 163.367
R683 B.n211 B.n144 163.367
R684 B.n215 B.n144 163.367
R685 B.n216 B.n215 163.367
R686 B.n282 B.t8 114.047
R687 B.n47 B.t1 114.047
R688 B.n126 B.t11 114.037
R689 B.n39 B.t4 114.037
R690 B.n126 B.n125 67.2975
R691 B.n282 B.n281 67.2975
R692 B.n47 B.n46 67.2975
R693 B.n39 B.n38 67.2975
R694 B.n267 B.n126 59.5399
R695 B.n283 B.n282 59.5399
R696 B.n48 B.n47 59.5399
R697 B.n517 B.n39 59.5399
R698 B.n567 B.n566 35.1225
R699 B.n452 B.n451 35.1225
R700 B.n336 B.n103 35.1225
R701 B.n218 B.n143 35.1225
R702 B B.n625 18.0485
R703 B.n567 B.n20 10.6151
R704 B.n571 B.n20 10.6151
R705 B.n572 B.n571 10.6151
R706 B.n573 B.n572 10.6151
R707 B.n573 B.n18 10.6151
R708 B.n577 B.n18 10.6151
R709 B.n578 B.n577 10.6151
R710 B.n579 B.n578 10.6151
R711 B.n579 B.n16 10.6151
R712 B.n583 B.n16 10.6151
R713 B.n584 B.n583 10.6151
R714 B.n585 B.n584 10.6151
R715 B.n585 B.n14 10.6151
R716 B.n589 B.n14 10.6151
R717 B.n590 B.n589 10.6151
R718 B.n591 B.n590 10.6151
R719 B.n591 B.n12 10.6151
R720 B.n595 B.n12 10.6151
R721 B.n596 B.n595 10.6151
R722 B.n597 B.n596 10.6151
R723 B.n597 B.n10 10.6151
R724 B.n601 B.n10 10.6151
R725 B.n602 B.n601 10.6151
R726 B.n603 B.n602 10.6151
R727 B.n603 B.n8 10.6151
R728 B.n607 B.n8 10.6151
R729 B.n608 B.n607 10.6151
R730 B.n609 B.n608 10.6151
R731 B.n609 B.n6 10.6151
R732 B.n613 B.n6 10.6151
R733 B.n614 B.n613 10.6151
R734 B.n615 B.n614 10.6151
R735 B.n615 B.n4 10.6151
R736 B.n619 B.n4 10.6151
R737 B.n620 B.n619 10.6151
R738 B.n621 B.n620 10.6151
R739 B.n621 B.n0 10.6151
R740 B.n566 B.n565 10.6151
R741 B.n565 B.n22 10.6151
R742 B.n561 B.n22 10.6151
R743 B.n561 B.n560 10.6151
R744 B.n560 B.n559 10.6151
R745 B.n559 B.n24 10.6151
R746 B.n555 B.n24 10.6151
R747 B.n555 B.n554 10.6151
R748 B.n554 B.n553 10.6151
R749 B.n553 B.n26 10.6151
R750 B.n549 B.n26 10.6151
R751 B.n549 B.n548 10.6151
R752 B.n548 B.n547 10.6151
R753 B.n547 B.n28 10.6151
R754 B.n543 B.n28 10.6151
R755 B.n543 B.n542 10.6151
R756 B.n542 B.n541 10.6151
R757 B.n541 B.n30 10.6151
R758 B.n537 B.n30 10.6151
R759 B.n537 B.n536 10.6151
R760 B.n536 B.n535 10.6151
R761 B.n535 B.n32 10.6151
R762 B.n531 B.n32 10.6151
R763 B.n531 B.n530 10.6151
R764 B.n530 B.n529 10.6151
R765 B.n529 B.n34 10.6151
R766 B.n525 B.n34 10.6151
R767 B.n525 B.n524 10.6151
R768 B.n524 B.n523 10.6151
R769 B.n523 B.n36 10.6151
R770 B.n519 B.n36 10.6151
R771 B.n519 B.n518 10.6151
R772 B.n516 B.n40 10.6151
R773 B.n512 B.n40 10.6151
R774 B.n512 B.n511 10.6151
R775 B.n511 B.n510 10.6151
R776 B.n510 B.n42 10.6151
R777 B.n506 B.n42 10.6151
R778 B.n506 B.n505 10.6151
R779 B.n505 B.n504 10.6151
R780 B.n504 B.n44 10.6151
R781 B.n500 B.n499 10.6151
R782 B.n499 B.n498 10.6151
R783 B.n498 B.n49 10.6151
R784 B.n494 B.n49 10.6151
R785 B.n494 B.n493 10.6151
R786 B.n493 B.n492 10.6151
R787 B.n492 B.n51 10.6151
R788 B.n488 B.n51 10.6151
R789 B.n488 B.n487 10.6151
R790 B.n487 B.n486 10.6151
R791 B.n486 B.n53 10.6151
R792 B.n482 B.n53 10.6151
R793 B.n482 B.n481 10.6151
R794 B.n481 B.n480 10.6151
R795 B.n480 B.n55 10.6151
R796 B.n476 B.n55 10.6151
R797 B.n476 B.n475 10.6151
R798 B.n475 B.n474 10.6151
R799 B.n474 B.n57 10.6151
R800 B.n470 B.n57 10.6151
R801 B.n470 B.n469 10.6151
R802 B.n469 B.n468 10.6151
R803 B.n468 B.n59 10.6151
R804 B.n464 B.n59 10.6151
R805 B.n464 B.n463 10.6151
R806 B.n463 B.n462 10.6151
R807 B.n462 B.n61 10.6151
R808 B.n458 B.n61 10.6151
R809 B.n458 B.n457 10.6151
R810 B.n457 B.n456 10.6151
R811 B.n456 B.n63 10.6151
R812 B.n452 B.n63 10.6151
R813 B.n451 B.n450 10.6151
R814 B.n450 B.n65 10.6151
R815 B.n446 B.n65 10.6151
R816 B.n446 B.n445 10.6151
R817 B.n445 B.n444 10.6151
R818 B.n444 B.n67 10.6151
R819 B.n440 B.n67 10.6151
R820 B.n440 B.n439 10.6151
R821 B.n439 B.n438 10.6151
R822 B.n438 B.n69 10.6151
R823 B.n434 B.n69 10.6151
R824 B.n434 B.n433 10.6151
R825 B.n433 B.n432 10.6151
R826 B.n432 B.n71 10.6151
R827 B.n428 B.n71 10.6151
R828 B.n428 B.n427 10.6151
R829 B.n427 B.n426 10.6151
R830 B.n426 B.n73 10.6151
R831 B.n422 B.n73 10.6151
R832 B.n422 B.n421 10.6151
R833 B.n421 B.n420 10.6151
R834 B.n420 B.n75 10.6151
R835 B.n416 B.n75 10.6151
R836 B.n416 B.n415 10.6151
R837 B.n415 B.n414 10.6151
R838 B.n414 B.n77 10.6151
R839 B.n410 B.n77 10.6151
R840 B.n410 B.n409 10.6151
R841 B.n409 B.n408 10.6151
R842 B.n408 B.n79 10.6151
R843 B.n404 B.n79 10.6151
R844 B.n404 B.n403 10.6151
R845 B.n403 B.n402 10.6151
R846 B.n402 B.n81 10.6151
R847 B.n398 B.n81 10.6151
R848 B.n398 B.n397 10.6151
R849 B.n397 B.n396 10.6151
R850 B.n396 B.n83 10.6151
R851 B.n392 B.n83 10.6151
R852 B.n392 B.n391 10.6151
R853 B.n391 B.n390 10.6151
R854 B.n390 B.n85 10.6151
R855 B.n386 B.n85 10.6151
R856 B.n386 B.n385 10.6151
R857 B.n385 B.n384 10.6151
R858 B.n384 B.n87 10.6151
R859 B.n380 B.n87 10.6151
R860 B.n380 B.n379 10.6151
R861 B.n379 B.n378 10.6151
R862 B.n378 B.n89 10.6151
R863 B.n374 B.n89 10.6151
R864 B.n374 B.n373 10.6151
R865 B.n373 B.n372 10.6151
R866 B.n372 B.n91 10.6151
R867 B.n368 B.n91 10.6151
R868 B.n368 B.n367 10.6151
R869 B.n367 B.n366 10.6151
R870 B.n366 B.n93 10.6151
R871 B.n362 B.n93 10.6151
R872 B.n362 B.n361 10.6151
R873 B.n361 B.n360 10.6151
R874 B.n360 B.n95 10.6151
R875 B.n356 B.n95 10.6151
R876 B.n356 B.n355 10.6151
R877 B.n355 B.n354 10.6151
R878 B.n354 B.n97 10.6151
R879 B.n350 B.n97 10.6151
R880 B.n350 B.n349 10.6151
R881 B.n349 B.n348 10.6151
R882 B.n348 B.n99 10.6151
R883 B.n344 B.n99 10.6151
R884 B.n344 B.n343 10.6151
R885 B.n343 B.n342 10.6151
R886 B.n342 B.n101 10.6151
R887 B.n338 B.n101 10.6151
R888 B.n338 B.n337 10.6151
R889 B.n337 B.n336 10.6151
R890 B.n161 B.n1 10.6151
R891 B.n164 B.n161 10.6151
R892 B.n165 B.n164 10.6151
R893 B.n166 B.n165 10.6151
R894 B.n166 B.n159 10.6151
R895 B.n170 B.n159 10.6151
R896 B.n171 B.n170 10.6151
R897 B.n172 B.n171 10.6151
R898 B.n172 B.n157 10.6151
R899 B.n176 B.n157 10.6151
R900 B.n177 B.n176 10.6151
R901 B.n178 B.n177 10.6151
R902 B.n178 B.n155 10.6151
R903 B.n182 B.n155 10.6151
R904 B.n183 B.n182 10.6151
R905 B.n184 B.n183 10.6151
R906 B.n184 B.n153 10.6151
R907 B.n188 B.n153 10.6151
R908 B.n189 B.n188 10.6151
R909 B.n190 B.n189 10.6151
R910 B.n190 B.n151 10.6151
R911 B.n194 B.n151 10.6151
R912 B.n195 B.n194 10.6151
R913 B.n196 B.n195 10.6151
R914 B.n196 B.n149 10.6151
R915 B.n200 B.n149 10.6151
R916 B.n201 B.n200 10.6151
R917 B.n202 B.n201 10.6151
R918 B.n202 B.n147 10.6151
R919 B.n206 B.n147 10.6151
R920 B.n207 B.n206 10.6151
R921 B.n208 B.n207 10.6151
R922 B.n208 B.n145 10.6151
R923 B.n212 B.n145 10.6151
R924 B.n213 B.n212 10.6151
R925 B.n214 B.n213 10.6151
R926 B.n214 B.n143 10.6151
R927 B.n219 B.n218 10.6151
R928 B.n220 B.n219 10.6151
R929 B.n220 B.n141 10.6151
R930 B.n224 B.n141 10.6151
R931 B.n225 B.n224 10.6151
R932 B.n226 B.n225 10.6151
R933 B.n226 B.n139 10.6151
R934 B.n230 B.n139 10.6151
R935 B.n231 B.n230 10.6151
R936 B.n232 B.n231 10.6151
R937 B.n232 B.n137 10.6151
R938 B.n236 B.n137 10.6151
R939 B.n237 B.n236 10.6151
R940 B.n238 B.n237 10.6151
R941 B.n238 B.n135 10.6151
R942 B.n242 B.n135 10.6151
R943 B.n243 B.n242 10.6151
R944 B.n244 B.n243 10.6151
R945 B.n244 B.n133 10.6151
R946 B.n248 B.n133 10.6151
R947 B.n249 B.n248 10.6151
R948 B.n250 B.n249 10.6151
R949 B.n250 B.n131 10.6151
R950 B.n254 B.n131 10.6151
R951 B.n255 B.n254 10.6151
R952 B.n256 B.n255 10.6151
R953 B.n256 B.n129 10.6151
R954 B.n260 B.n129 10.6151
R955 B.n261 B.n260 10.6151
R956 B.n262 B.n261 10.6151
R957 B.n262 B.n127 10.6151
R958 B.n266 B.n127 10.6151
R959 B.n269 B.n268 10.6151
R960 B.n269 B.n123 10.6151
R961 B.n273 B.n123 10.6151
R962 B.n274 B.n273 10.6151
R963 B.n275 B.n274 10.6151
R964 B.n275 B.n121 10.6151
R965 B.n279 B.n121 10.6151
R966 B.n280 B.n279 10.6151
R967 B.n284 B.n280 10.6151
R968 B.n288 B.n119 10.6151
R969 B.n289 B.n288 10.6151
R970 B.n290 B.n289 10.6151
R971 B.n290 B.n117 10.6151
R972 B.n294 B.n117 10.6151
R973 B.n295 B.n294 10.6151
R974 B.n296 B.n295 10.6151
R975 B.n296 B.n115 10.6151
R976 B.n300 B.n115 10.6151
R977 B.n301 B.n300 10.6151
R978 B.n302 B.n301 10.6151
R979 B.n302 B.n113 10.6151
R980 B.n306 B.n113 10.6151
R981 B.n307 B.n306 10.6151
R982 B.n308 B.n307 10.6151
R983 B.n308 B.n111 10.6151
R984 B.n312 B.n111 10.6151
R985 B.n313 B.n312 10.6151
R986 B.n314 B.n313 10.6151
R987 B.n314 B.n109 10.6151
R988 B.n318 B.n109 10.6151
R989 B.n319 B.n318 10.6151
R990 B.n320 B.n319 10.6151
R991 B.n320 B.n107 10.6151
R992 B.n324 B.n107 10.6151
R993 B.n325 B.n324 10.6151
R994 B.n326 B.n325 10.6151
R995 B.n326 B.n105 10.6151
R996 B.n330 B.n105 10.6151
R997 B.n331 B.n330 10.6151
R998 B.n332 B.n331 10.6151
R999 B.n332 B.n103 10.6151
R1000 B.n518 B.n517 9.36635
R1001 B.n500 B.n48 9.36635
R1002 B.n267 B.n266 9.36635
R1003 B.n283 B.n119 9.36635
R1004 B.n625 B.n0 8.11757
R1005 B.n625 B.n1 8.11757
R1006 B.n517 B.n516 1.24928
R1007 B.n48 B.n44 1.24928
R1008 B.n268 B.n267 1.24928
R1009 B.n284 B.n283 1.24928
C0 VN VTAIL 3.93481f
C1 w_n3052_n2798# VDD1 1.48133f
C2 VDD2 VDD1 1.15945f
C3 VP VDD1 4.08773f
C4 B VDD1 1.28012f
C5 VDD2 w_n3052_n2798# 1.54941f
C6 B w_n3052_n2798# 9.110519f
C7 w_n3052_n2798# VP 5.59961f
C8 VDD1 VTAIL 4.89573f
C9 B VDD2 1.34123f
C10 VDD2 VP 0.428811f
C11 B VP 1.83366f
C12 w_n3052_n2798# VTAIL 3.36059f
C13 VN VDD1 0.149632f
C14 VDD2 VTAIL 4.95356f
C15 B VTAIL 4.21429f
C16 VP VTAIL 3.94891f
C17 w_n3052_n2798# VN 5.2059f
C18 VDD2 VN 3.80943f
C19 VN VP 6.04957f
C20 B VN 1.1778f
C21 VDD2 VSUBS 0.965778f
C22 VDD1 VSUBS 5.72294f
C23 VTAIL VSUBS 1.154785f
C24 VN VSUBS 5.680901f
C25 VP VSUBS 2.485037f
C26 B VSUBS 4.500538f
C27 w_n3052_n2798# VSUBS 0.10566p
C28 B.n0 VSUBS 0.006175f
C29 B.n1 VSUBS 0.006175f
C30 B.n2 VSUBS 0.009133f
C31 B.n3 VSUBS 0.006999f
C32 B.n4 VSUBS 0.006999f
C33 B.n5 VSUBS 0.006999f
C34 B.n6 VSUBS 0.006999f
C35 B.n7 VSUBS 0.006999f
C36 B.n8 VSUBS 0.006999f
C37 B.n9 VSUBS 0.006999f
C38 B.n10 VSUBS 0.006999f
C39 B.n11 VSUBS 0.006999f
C40 B.n12 VSUBS 0.006999f
C41 B.n13 VSUBS 0.006999f
C42 B.n14 VSUBS 0.006999f
C43 B.n15 VSUBS 0.006999f
C44 B.n16 VSUBS 0.006999f
C45 B.n17 VSUBS 0.006999f
C46 B.n18 VSUBS 0.006999f
C47 B.n19 VSUBS 0.006999f
C48 B.n20 VSUBS 0.006999f
C49 B.n21 VSUBS 0.017685f
C50 B.n22 VSUBS 0.006999f
C51 B.n23 VSUBS 0.006999f
C52 B.n24 VSUBS 0.006999f
C53 B.n25 VSUBS 0.006999f
C54 B.n26 VSUBS 0.006999f
C55 B.n27 VSUBS 0.006999f
C56 B.n28 VSUBS 0.006999f
C57 B.n29 VSUBS 0.006999f
C58 B.n30 VSUBS 0.006999f
C59 B.n31 VSUBS 0.006999f
C60 B.n32 VSUBS 0.006999f
C61 B.n33 VSUBS 0.006999f
C62 B.n34 VSUBS 0.006999f
C63 B.n35 VSUBS 0.006999f
C64 B.n36 VSUBS 0.006999f
C65 B.n37 VSUBS 0.006999f
C66 B.t4 VSUBS 0.288166f
C67 B.t5 VSUBS 0.311855f
C68 B.t3 VSUBS 1.34414f
C69 B.n38 VSUBS 0.17264f
C70 B.n39 VSUBS 0.073812f
C71 B.n40 VSUBS 0.006999f
C72 B.n41 VSUBS 0.006999f
C73 B.n42 VSUBS 0.006999f
C74 B.n43 VSUBS 0.006999f
C75 B.n44 VSUBS 0.003911f
C76 B.n45 VSUBS 0.006999f
C77 B.t1 VSUBS 0.288163f
C78 B.t2 VSUBS 0.311852f
C79 B.t0 VSUBS 1.34414f
C80 B.n46 VSUBS 0.172644f
C81 B.n47 VSUBS 0.073815f
C82 B.n48 VSUBS 0.016215f
C83 B.n49 VSUBS 0.006999f
C84 B.n50 VSUBS 0.006999f
C85 B.n51 VSUBS 0.006999f
C86 B.n52 VSUBS 0.006999f
C87 B.n53 VSUBS 0.006999f
C88 B.n54 VSUBS 0.006999f
C89 B.n55 VSUBS 0.006999f
C90 B.n56 VSUBS 0.006999f
C91 B.n57 VSUBS 0.006999f
C92 B.n58 VSUBS 0.006999f
C93 B.n59 VSUBS 0.006999f
C94 B.n60 VSUBS 0.006999f
C95 B.n61 VSUBS 0.006999f
C96 B.n62 VSUBS 0.006999f
C97 B.n63 VSUBS 0.006999f
C98 B.n64 VSUBS 0.016691f
C99 B.n65 VSUBS 0.006999f
C100 B.n66 VSUBS 0.006999f
C101 B.n67 VSUBS 0.006999f
C102 B.n68 VSUBS 0.006999f
C103 B.n69 VSUBS 0.006999f
C104 B.n70 VSUBS 0.006999f
C105 B.n71 VSUBS 0.006999f
C106 B.n72 VSUBS 0.006999f
C107 B.n73 VSUBS 0.006999f
C108 B.n74 VSUBS 0.006999f
C109 B.n75 VSUBS 0.006999f
C110 B.n76 VSUBS 0.006999f
C111 B.n77 VSUBS 0.006999f
C112 B.n78 VSUBS 0.006999f
C113 B.n79 VSUBS 0.006999f
C114 B.n80 VSUBS 0.006999f
C115 B.n81 VSUBS 0.006999f
C116 B.n82 VSUBS 0.006999f
C117 B.n83 VSUBS 0.006999f
C118 B.n84 VSUBS 0.006999f
C119 B.n85 VSUBS 0.006999f
C120 B.n86 VSUBS 0.006999f
C121 B.n87 VSUBS 0.006999f
C122 B.n88 VSUBS 0.006999f
C123 B.n89 VSUBS 0.006999f
C124 B.n90 VSUBS 0.006999f
C125 B.n91 VSUBS 0.006999f
C126 B.n92 VSUBS 0.006999f
C127 B.n93 VSUBS 0.006999f
C128 B.n94 VSUBS 0.006999f
C129 B.n95 VSUBS 0.006999f
C130 B.n96 VSUBS 0.006999f
C131 B.n97 VSUBS 0.006999f
C132 B.n98 VSUBS 0.006999f
C133 B.n99 VSUBS 0.006999f
C134 B.n100 VSUBS 0.006999f
C135 B.n101 VSUBS 0.006999f
C136 B.n102 VSUBS 0.006999f
C137 B.n103 VSUBS 0.016916f
C138 B.n104 VSUBS 0.006999f
C139 B.n105 VSUBS 0.006999f
C140 B.n106 VSUBS 0.006999f
C141 B.n107 VSUBS 0.006999f
C142 B.n108 VSUBS 0.006999f
C143 B.n109 VSUBS 0.006999f
C144 B.n110 VSUBS 0.006999f
C145 B.n111 VSUBS 0.006999f
C146 B.n112 VSUBS 0.006999f
C147 B.n113 VSUBS 0.006999f
C148 B.n114 VSUBS 0.006999f
C149 B.n115 VSUBS 0.006999f
C150 B.n116 VSUBS 0.006999f
C151 B.n117 VSUBS 0.006999f
C152 B.n118 VSUBS 0.006999f
C153 B.n119 VSUBS 0.006587f
C154 B.n120 VSUBS 0.006999f
C155 B.n121 VSUBS 0.006999f
C156 B.n122 VSUBS 0.006999f
C157 B.n123 VSUBS 0.006999f
C158 B.n124 VSUBS 0.006999f
C159 B.t11 VSUBS 0.288166f
C160 B.t10 VSUBS 0.311855f
C161 B.t9 VSUBS 1.34414f
C162 B.n125 VSUBS 0.17264f
C163 B.n126 VSUBS 0.073812f
C164 B.n127 VSUBS 0.006999f
C165 B.n128 VSUBS 0.006999f
C166 B.n129 VSUBS 0.006999f
C167 B.n130 VSUBS 0.006999f
C168 B.n131 VSUBS 0.006999f
C169 B.n132 VSUBS 0.006999f
C170 B.n133 VSUBS 0.006999f
C171 B.n134 VSUBS 0.006999f
C172 B.n135 VSUBS 0.006999f
C173 B.n136 VSUBS 0.006999f
C174 B.n137 VSUBS 0.006999f
C175 B.n138 VSUBS 0.006999f
C176 B.n139 VSUBS 0.006999f
C177 B.n140 VSUBS 0.006999f
C178 B.n141 VSUBS 0.006999f
C179 B.n142 VSUBS 0.006999f
C180 B.n143 VSUBS 0.016691f
C181 B.n144 VSUBS 0.006999f
C182 B.n145 VSUBS 0.006999f
C183 B.n146 VSUBS 0.006999f
C184 B.n147 VSUBS 0.006999f
C185 B.n148 VSUBS 0.006999f
C186 B.n149 VSUBS 0.006999f
C187 B.n150 VSUBS 0.006999f
C188 B.n151 VSUBS 0.006999f
C189 B.n152 VSUBS 0.006999f
C190 B.n153 VSUBS 0.006999f
C191 B.n154 VSUBS 0.006999f
C192 B.n155 VSUBS 0.006999f
C193 B.n156 VSUBS 0.006999f
C194 B.n157 VSUBS 0.006999f
C195 B.n158 VSUBS 0.006999f
C196 B.n159 VSUBS 0.006999f
C197 B.n160 VSUBS 0.006999f
C198 B.n161 VSUBS 0.006999f
C199 B.n162 VSUBS 0.006999f
C200 B.n163 VSUBS 0.006999f
C201 B.n164 VSUBS 0.006999f
C202 B.n165 VSUBS 0.006999f
C203 B.n166 VSUBS 0.006999f
C204 B.n167 VSUBS 0.006999f
C205 B.n168 VSUBS 0.006999f
C206 B.n169 VSUBS 0.006999f
C207 B.n170 VSUBS 0.006999f
C208 B.n171 VSUBS 0.006999f
C209 B.n172 VSUBS 0.006999f
C210 B.n173 VSUBS 0.006999f
C211 B.n174 VSUBS 0.006999f
C212 B.n175 VSUBS 0.006999f
C213 B.n176 VSUBS 0.006999f
C214 B.n177 VSUBS 0.006999f
C215 B.n178 VSUBS 0.006999f
C216 B.n179 VSUBS 0.006999f
C217 B.n180 VSUBS 0.006999f
C218 B.n181 VSUBS 0.006999f
C219 B.n182 VSUBS 0.006999f
C220 B.n183 VSUBS 0.006999f
C221 B.n184 VSUBS 0.006999f
C222 B.n185 VSUBS 0.006999f
C223 B.n186 VSUBS 0.006999f
C224 B.n187 VSUBS 0.006999f
C225 B.n188 VSUBS 0.006999f
C226 B.n189 VSUBS 0.006999f
C227 B.n190 VSUBS 0.006999f
C228 B.n191 VSUBS 0.006999f
C229 B.n192 VSUBS 0.006999f
C230 B.n193 VSUBS 0.006999f
C231 B.n194 VSUBS 0.006999f
C232 B.n195 VSUBS 0.006999f
C233 B.n196 VSUBS 0.006999f
C234 B.n197 VSUBS 0.006999f
C235 B.n198 VSUBS 0.006999f
C236 B.n199 VSUBS 0.006999f
C237 B.n200 VSUBS 0.006999f
C238 B.n201 VSUBS 0.006999f
C239 B.n202 VSUBS 0.006999f
C240 B.n203 VSUBS 0.006999f
C241 B.n204 VSUBS 0.006999f
C242 B.n205 VSUBS 0.006999f
C243 B.n206 VSUBS 0.006999f
C244 B.n207 VSUBS 0.006999f
C245 B.n208 VSUBS 0.006999f
C246 B.n209 VSUBS 0.006999f
C247 B.n210 VSUBS 0.006999f
C248 B.n211 VSUBS 0.006999f
C249 B.n212 VSUBS 0.006999f
C250 B.n213 VSUBS 0.006999f
C251 B.n214 VSUBS 0.006999f
C252 B.n215 VSUBS 0.006999f
C253 B.n216 VSUBS 0.016691f
C254 B.n217 VSUBS 0.017685f
C255 B.n218 VSUBS 0.017685f
C256 B.n219 VSUBS 0.006999f
C257 B.n220 VSUBS 0.006999f
C258 B.n221 VSUBS 0.006999f
C259 B.n222 VSUBS 0.006999f
C260 B.n223 VSUBS 0.006999f
C261 B.n224 VSUBS 0.006999f
C262 B.n225 VSUBS 0.006999f
C263 B.n226 VSUBS 0.006999f
C264 B.n227 VSUBS 0.006999f
C265 B.n228 VSUBS 0.006999f
C266 B.n229 VSUBS 0.006999f
C267 B.n230 VSUBS 0.006999f
C268 B.n231 VSUBS 0.006999f
C269 B.n232 VSUBS 0.006999f
C270 B.n233 VSUBS 0.006999f
C271 B.n234 VSUBS 0.006999f
C272 B.n235 VSUBS 0.006999f
C273 B.n236 VSUBS 0.006999f
C274 B.n237 VSUBS 0.006999f
C275 B.n238 VSUBS 0.006999f
C276 B.n239 VSUBS 0.006999f
C277 B.n240 VSUBS 0.006999f
C278 B.n241 VSUBS 0.006999f
C279 B.n242 VSUBS 0.006999f
C280 B.n243 VSUBS 0.006999f
C281 B.n244 VSUBS 0.006999f
C282 B.n245 VSUBS 0.006999f
C283 B.n246 VSUBS 0.006999f
C284 B.n247 VSUBS 0.006999f
C285 B.n248 VSUBS 0.006999f
C286 B.n249 VSUBS 0.006999f
C287 B.n250 VSUBS 0.006999f
C288 B.n251 VSUBS 0.006999f
C289 B.n252 VSUBS 0.006999f
C290 B.n253 VSUBS 0.006999f
C291 B.n254 VSUBS 0.006999f
C292 B.n255 VSUBS 0.006999f
C293 B.n256 VSUBS 0.006999f
C294 B.n257 VSUBS 0.006999f
C295 B.n258 VSUBS 0.006999f
C296 B.n259 VSUBS 0.006999f
C297 B.n260 VSUBS 0.006999f
C298 B.n261 VSUBS 0.006999f
C299 B.n262 VSUBS 0.006999f
C300 B.n263 VSUBS 0.006999f
C301 B.n264 VSUBS 0.006999f
C302 B.n265 VSUBS 0.006999f
C303 B.n266 VSUBS 0.006587f
C304 B.n267 VSUBS 0.016215f
C305 B.n268 VSUBS 0.003911f
C306 B.n269 VSUBS 0.006999f
C307 B.n270 VSUBS 0.006999f
C308 B.n271 VSUBS 0.006999f
C309 B.n272 VSUBS 0.006999f
C310 B.n273 VSUBS 0.006999f
C311 B.n274 VSUBS 0.006999f
C312 B.n275 VSUBS 0.006999f
C313 B.n276 VSUBS 0.006999f
C314 B.n277 VSUBS 0.006999f
C315 B.n278 VSUBS 0.006999f
C316 B.n279 VSUBS 0.006999f
C317 B.n280 VSUBS 0.006999f
C318 B.t8 VSUBS 0.288163f
C319 B.t7 VSUBS 0.311852f
C320 B.t6 VSUBS 1.34414f
C321 B.n281 VSUBS 0.172644f
C322 B.n282 VSUBS 0.073815f
C323 B.n283 VSUBS 0.016215f
C324 B.n284 VSUBS 0.003911f
C325 B.n285 VSUBS 0.006999f
C326 B.n286 VSUBS 0.006999f
C327 B.n287 VSUBS 0.006999f
C328 B.n288 VSUBS 0.006999f
C329 B.n289 VSUBS 0.006999f
C330 B.n290 VSUBS 0.006999f
C331 B.n291 VSUBS 0.006999f
C332 B.n292 VSUBS 0.006999f
C333 B.n293 VSUBS 0.006999f
C334 B.n294 VSUBS 0.006999f
C335 B.n295 VSUBS 0.006999f
C336 B.n296 VSUBS 0.006999f
C337 B.n297 VSUBS 0.006999f
C338 B.n298 VSUBS 0.006999f
C339 B.n299 VSUBS 0.006999f
C340 B.n300 VSUBS 0.006999f
C341 B.n301 VSUBS 0.006999f
C342 B.n302 VSUBS 0.006999f
C343 B.n303 VSUBS 0.006999f
C344 B.n304 VSUBS 0.006999f
C345 B.n305 VSUBS 0.006999f
C346 B.n306 VSUBS 0.006999f
C347 B.n307 VSUBS 0.006999f
C348 B.n308 VSUBS 0.006999f
C349 B.n309 VSUBS 0.006999f
C350 B.n310 VSUBS 0.006999f
C351 B.n311 VSUBS 0.006999f
C352 B.n312 VSUBS 0.006999f
C353 B.n313 VSUBS 0.006999f
C354 B.n314 VSUBS 0.006999f
C355 B.n315 VSUBS 0.006999f
C356 B.n316 VSUBS 0.006999f
C357 B.n317 VSUBS 0.006999f
C358 B.n318 VSUBS 0.006999f
C359 B.n319 VSUBS 0.006999f
C360 B.n320 VSUBS 0.006999f
C361 B.n321 VSUBS 0.006999f
C362 B.n322 VSUBS 0.006999f
C363 B.n323 VSUBS 0.006999f
C364 B.n324 VSUBS 0.006999f
C365 B.n325 VSUBS 0.006999f
C366 B.n326 VSUBS 0.006999f
C367 B.n327 VSUBS 0.006999f
C368 B.n328 VSUBS 0.006999f
C369 B.n329 VSUBS 0.006999f
C370 B.n330 VSUBS 0.006999f
C371 B.n331 VSUBS 0.006999f
C372 B.n332 VSUBS 0.006999f
C373 B.n333 VSUBS 0.006999f
C374 B.n334 VSUBS 0.017685f
C375 B.n335 VSUBS 0.016691f
C376 B.n336 VSUBS 0.01746f
C377 B.n337 VSUBS 0.006999f
C378 B.n338 VSUBS 0.006999f
C379 B.n339 VSUBS 0.006999f
C380 B.n340 VSUBS 0.006999f
C381 B.n341 VSUBS 0.006999f
C382 B.n342 VSUBS 0.006999f
C383 B.n343 VSUBS 0.006999f
C384 B.n344 VSUBS 0.006999f
C385 B.n345 VSUBS 0.006999f
C386 B.n346 VSUBS 0.006999f
C387 B.n347 VSUBS 0.006999f
C388 B.n348 VSUBS 0.006999f
C389 B.n349 VSUBS 0.006999f
C390 B.n350 VSUBS 0.006999f
C391 B.n351 VSUBS 0.006999f
C392 B.n352 VSUBS 0.006999f
C393 B.n353 VSUBS 0.006999f
C394 B.n354 VSUBS 0.006999f
C395 B.n355 VSUBS 0.006999f
C396 B.n356 VSUBS 0.006999f
C397 B.n357 VSUBS 0.006999f
C398 B.n358 VSUBS 0.006999f
C399 B.n359 VSUBS 0.006999f
C400 B.n360 VSUBS 0.006999f
C401 B.n361 VSUBS 0.006999f
C402 B.n362 VSUBS 0.006999f
C403 B.n363 VSUBS 0.006999f
C404 B.n364 VSUBS 0.006999f
C405 B.n365 VSUBS 0.006999f
C406 B.n366 VSUBS 0.006999f
C407 B.n367 VSUBS 0.006999f
C408 B.n368 VSUBS 0.006999f
C409 B.n369 VSUBS 0.006999f
C410 B.n370 VSUBS 0.006999f
C411 B.n371 VSUBS 0.006999f
C412 B.n372 VSUBS 0.006999f
C413 B.n373 VSUBS 0.006999f
C414 B.n374 VSUBS 0.006999f
C415 B.n375 VSUBS 0.006999f
C416 B.n376 VSUBS 0.006999f
C417 B.n377 VSUBS 0.006999f
C418 B.n378 VSUBS 0.006999f
C419 B.n379 VSUBS 0.006999f
C420 B.n380 VSUBS 0.006999f
C421 B.n381 VSUBS 0.006999f
C422 B.n382 VSUBS 0.006999f
C423 B.n383 VSUBS 0.006999f
C424 B.n384 VSUBS 0.006999f
C425 B.n385 VSUBS 0.006999f
C426 B.n386 VSUBS 0.006999f
C427 B.n387 VSUBS 0.006999f
C428 B.n388 VSUBS 0.006999f
C429 B.n389 VSUBS 0.006999f
C430 B.n390 VSUBS 0.006999f
C431 B.n391 VSUBS 0.006999f
C432 B.n392 VSUBS 0.006999f
C433 B.n393 VSUBS 0.006999f
C434 B.n394 VSUBS 0.006999f
C435 B.n395 VSUBS 0.006999f
C436 B.n396 VSUBS 0.006999f
C437 B.n397 VSUBS 0.006999f
C438 B.n398 VSUBS 0.006999f
C439 B.n399 VSUBS 0.006999f
C440 B.n400 VSUBS 0.006999f
C441 B.n401 VSUBS 0.006999f
C442 B.n402 VSUBS 0.006999f
C443 B.n403 VSUBS 0.006999f
C444 B.n404 VSUBS 0.006999f
C445 B.n405 VSUBS 0.006999f
C446 B.n406 VSUBS 0.006999f
C447 B.n407 VSUBS 0.006999f
C448 B.n408 VSUBS 0.006999f
C449 B.n409 VSUBS 0.006999f
C450 B.n410 VSUBS 0.006999f
C451 B.n411 VSUBS 0.006999f
C452 B.n412 VSUBS 0.006999f
C453 B.n413 VSUBS 0.006999f
C454 B.n414 VSUBS 0.006999f
C455 B.n415 VSUBS 0.006999f
C456 B.n416 VSUBS 0.006999f
C457 B.n417 VSUBS 0.006999f
C458 B.n418 VSUBS 0.006999f
C459 B.n419 VSUBS 0.006999f
C460 B.n420 VSUBS 0.006999f
C461 B.n421 VSUBS 0.006999f
C462 B.n422 VSUBS 0.006999f
C463 B.n423 VSUBS 0.006999f
C464 B.n424 VSUBS 0.006999f
C465 B.n425 VSUBS 0.006999f
C466 B.n426 VSUBS 0.006999f
C467 B.n427 VSUBS 0.006999f
C468 B.n428 VSUBS 0.006999f
C469 B.n429 VSUBS 0.006999f
C470 B.n430 VSUBS 0.006999f
C471 B.n431 VSUBS 0.006999f
C472 B.n432 VSUBS 0.006999f
C473 B.n433 VSUBS 0.006999f
C474 B.n434 VSUBS 0.006999f
C475 B.n435 VSUBS 0.006999f
C476 B.n436 VSUBS 0.006999f
C477 B.n437 VSUBS 0.006999f
C478 B.n438 VSUBS 0.006999f
C479 B.n439 VSUBS 0.006999f
C480 B.n440 VSUBS 0.006999f
C481 B.n441 VSUBS 0.006999f
C482 B.n442 VSUBS 0.006999f
C483 B.n443 VSUBS 0.006999f
C484 B.n444 VSUBS 0.006999f
C485 B.n445 VSUBS 0.006999f
C486 B.n446 VSUBS 0.006999f
C487 B.n447 VSUBS 0.006999f
C488 B.n448 VSUBS 0.006999f
C489 B.n449 VSUBS 0.006999f
C490 B.n450 VSUBS 0.006999f
C491 B.n451 VSUBS 0.016691f
C492 B.n452 VSUBS 0.017685f
C493 B.n453 VSUBS 0.017685f
C494 B.n454 VSUBS 0.006999f
C495 B.n455 VSUBS 0.006999f
C496 B.n456 VSUBS 0.006999f
C497 B.n457 VSUBS 0.006999f
C498 B.n458 VSUBS 0.006999f
C499 B.n459 VSUBS 0.006999f
C500 B.n460 VSUBS 0.006999f
C501 B.n461 VSUBS 0.006999f
C502 B.n462 VSUBS 0.006999f
C503 B.n463 VSUBS 0.006999f
C504 B.n464 VSUBS 0.006999f
C505 B.n465 VSUBS 0.006999f
C506 B.n466 VSUBS 0.006999f
C507 B.n467 VSUBS 0.006999f
C508 B.n468 VSUBS 0.006999f
C509 B.n469 VSUBS 0.006999f
C510 B.n470 VSUBS 0.006999f
C511 B.n471 VSUBS 0.006999f
C512 B.n472 VSUBS 0.006999f
C513 B.n473 VSUBS 0.006999f
C514 B.n474 VSUBS 0.006999f
C515 B.n475 VSUBS 0.006999f
C516 B.n476 VSUBS 0.006999f
C517 B.n477 VSUBS 0.006999f
C518 B.n478 VSUBS 0.006999f
C519 B.n479 VSUBS 0.006999f
C520 B.n480 VSUBS 0.006999f
C521 B.n481 VSUBS 0.006999f
C522 B.n482 VSUBS 0.006999f
C523 B.n483 VSUBS 0.006999f
C524 B.n484 VSUBS 0.006999f
C525 B.n485 VSUBS 0.006999f
C526 B.n486 VSUBS 0.006999f
C527 B.n487 VSUBS 0.006999f
C528 B.n488 VSUBS 0.006999f
C529 B.n489 VSUBS 0.006999f
C530 B.n490 VSUBS 0.006999f
C531 B.n491 VSUBS 0.006999f
C532 B.n492 VSUBS 0.006999f
C533 B.n493 VSUBS 0.006999f
C534 B.n494 VSUBS 0.006999f
C535 B.n495 VSUBS 0.006999f
C536 B.n496 VSUBS 0.006999f
C537 B.n497 VSUBS 0.006999f
C538 B.n498 VSUBS 0.006999f
C539 B.n499 VSUBS 0.006999f
C540 B.n500 VSUBS 0.006587f
C541 B.n501 VSUBS 0.006999f
C542 B.n502 VSUBS 0.006999f
C543 B.n503 VSUBS 0.006999f
C544 B.n504 VSUBS 0.006999f
C545 B.n505 VSUBS 0.006999f
C546 B.n506 VSUBS 0.006999f
C547 B.n507 VSUBS 0.006999f
C548 B.n508 VSUBS 0.006999f
C549 B.n509 VSUBS 0.006999f
C550 B.n510 VSUBS 0.006999f
C551 B.n511 VSUBS 0.006999f
C552 B.n512 VSUBS 0.006999f
C553 B.n513 VSUBS 0.006999f
C554 B.n514 VSUBS 0.006999f
C555 B.n515 VSUBS 0.006999f
C556 B.n516 VSUBS 0.003911f
C557 B.n517 VSUBS 0.016215f
C558 B.n518 VSUBS 0.006587f
C559 B.n519 VSUBS 0.006999f
C560 B.n520 VSUBS 0.006999f
C561 B.n521 VSUBS 0.006999f
C562 B.n522 VSUBS 0.006999f
C563 B.n523 VSUBS 0.006999f
C564 B.n524 VSUBS 0.006999f
C565 B.n525 VSUBS 0.006999f
C566 B.n526 VSUBS 0.006999f
C567 B.n527 VSUBS 0.006999f
C568 B.n528 VSUBS 0.006999f
C569 B.n529 VSUBS 0.006999f
C570 B.n530 VSUBS 0.006999f
C571 B.n531 VSUBS 0.006999f
C572 B.n532 VSUBS 0.006999f
C573 B.n533 VSUBS 0.006999f
C574 B.n534 VSUBS 0.006999f
C575 B.n535 VSUBS 0.006999f
C576 B.n536 VSUBS 0.006999f
C577 B.n537 VSUBS 0.006999f
C578 B.n538 VSUBS 0.006999f
C579 B.n539 VSUBS 0.006999f
C580 B.n540 VSUBS 0.006999f
C581 B.n541 VSUBS 0.006999f
C582 B.n542 VSUBS 0.006999f
C583 B.n543 VSUBS 0.006999f
C584 B.n544 VSUBS 0.006999f
C585 B.n545 VSUBS 0.006999f
C586 B.n546 VSUBS 0.006999f
C587 B.n547 VSUBS 0.006999f
C588 B.n548 VSUBS 0.006999f
C589 B.n549 VSUBS 0.006999f
C590 B.n550 VSUBS 0.006999f
C591 B.n551 VSUBS 0.006999f
C592 B.n552 VSUBS 0.006999f
C593 B.n553 VSUBS 0.006999f
C594 B.n554 VSUBS 0.006999f
C595 B.n555 VSUBS 0.006999f
C596 B.n556 VSUBS 0.006999f
C597 B.n557 VSUBS 0.006999f
C598 B.n558 VSUBS 0.006999f
C599 B.n559 VSUBS 0.006999f
C600 B.n560 VSUBS 0.006999f
C601 B.n561 VSUBS 0.006999f
C602 B.n562 VSUBS 0.006999f
C603 B.n563 VSUBS 0.006999f
C604 B.n564 VSUBS 0.006999f
C605 B.n565 VSUBS 0.006999f
C606 B.n566 VSUBS 0.017685f
C607 B.n567 VSUBS 0.016691f
C608 B.n568 VSUBS 0.016691f
C609 B.n569 VSUBS 0.006999f
C610 B.n570 VSUBS 0.006999f
C611 B.n571 VSUBS 0.006999f
C612 B.n572 VSUBS 0.006999f
C613 B.n573 VSUBS 0.006999f
C614 B.n574 VSUBS 0.006999f
C615 B.n575 VSUBS 0.006999f
C616 B.n576 VSUBS 0.006999f
C617 B.n577 VSUBS 0.006999f
C618 B.n578 VSUBS 0.006999f
C619 B.n579 VSUBS 0.006999f
C620 B.n580 VSUBS 0.006999f
C621 B.n581 VSUBS 0.006999f
C622 B.n582 VSUBS 0.006999f
C623 B.n583 VSUBS 0.006999f
C624 B.n584 VSUBS 0.006999f
C625 B.n585 VSUBS 0.006999f
C626 B.n586 VSUBS 0.006999f
C627 B.n587 VSUBS 0.006999f
C628 B.n588 VSUBS 0.006999f
C629 B.n589 VSUBS 0.006999f
C630 B.n590 VSUBS 0.006999f
C631 B.n591 VSUBS 0.006999f
C632 B.n592 VSUBS 0.006999f
C633 B.n593 VSUBS 0.006999f
C634 B.n594 VSUBS 0.006999f
C635 B.n595 VSUBS 0.006999f
C636 B.n596 VSUBS 0.006999f
C637 B.n597 VSUBS 0.006999f
C638 B.n598 VSUBS 0.006999f
C639 B.n599 VSUBS 0.006999f
C640 B.n600 VSUBS 0.006999f
C641 B.n601 VSUBS 0.006999f
C642 B.n602 VSUBS 0.006999f
C643 B.n603 VSUBS 0.006999f
C644 B.n604 VSUBS 0.006999f
C645 B.n605 VSUBS 0.006999f
C646 B.n606 VSUBS 0.006999f
C647 B.n607 VSUBS 0.006999f
C648 B.n608 VSUBS 0.006999f
C649 B.n609 VSUBS 0.006999f
C650 B.n610 VSUBS 0.006999f
C651 B.n611 VSUBS 0.006999f
C652 B.n612 VSUBS 0.006999f
C653 B.n613 VSUBS 0.006999f
C654 B.n614 VSUBS 0.006999f
C655 B.n615 VSUBS 0.006999f
C656 B.n616 VSUBS 0.006999f
C657 B.n617 VSUBS 0.006999f
C658 B.n618 VSUBS 0.006999f
C659 B.n619 VSUBS 0.006999f
C660 B.n620 VSUBS 0.006999f
C661 B.n621 VSUBS 0.006999f
C662 B.n622 VSUBS 0.006999f
C663 B.n623 VSUBS 0.009133f
C664 B.n624 VSUBS 0.009729f
C665 B.n625 VSUBS 0.019346f
C666 VDD2.t3 VSUBS 0.198657f
C667 VDD2.t1 VSUBS 0.198657f
C668 VDD2.n0 VSUBS 2.08209f
C669 VDD2.t2 VSUBS 0.198657f
C670 VDD2.t0 VSUBS 0.198657f
C671 VDD2.n1 VSUBS 1.45491f
C672 VDD2.n2 VSUBS 4.19763f
C673 VN.t2 VSUBS 2.87097f
C674 VN.t0 VSUBS 2.88163f
C675 VN.n0 VSUBS 1.74708f
C676 VN.t3 VSUBS 2.88163f
C677 VN.t1 VSUBS 2.87097f
C678 VN.n1 VSUBS 3.57536f
C679 VDD1.t1 VSUBS 0.200856f
C680 VDD1.t3 VSUBS 0.200856f
C681 VDD1.n0 VSUBS 1.4716f
C682 VDD1.t0 VSUBS 0.200856f
C683 VDD1.t2 VSUBS 0.200856f
C684 VDD1.n1 VSUBS 2.12958f
C685 VTAIL.t2 VSUBS 1.63736f
C686 VTAIL.n0 VSUBS 0.808494f
C687 VTAIL.t4 VSUBS 1.63736f
C688 VTAIL.n1 VSUBS 0.926227f
C689 VTAIL.t7 VSUBS 1.63736f
C690 VTAIL.n2 VSUBS 2.12405f
C691 VTAIL.t0 VSUBS 1.63737f
C692 VTAIL.n3 VSUBS 2.12404f
C693 VTAIL.t3 VSUBS 1.63737f
C694 VTAIL.n4 VSUBS 0.926218f
C695 VTAIL.t6 VSUBS 1.63737f
C696 VTAIL.n5 VSUBS 0.926218f
C697 VTAIL.t5 VSUBS 1.63737f
C698 VTAIL.n6 VSUBS 2.12404f
C699 VTAIL.t1 VSUBS 1.63736f
C700 VTAIL.n7 VSUBS 1.99679f
C701 VP.t1 VSUBS 2.60479f
C702 VP.n0 VSUBS 1.07951f
C703 VP.n1 VSUBS 0.033574f
C704 VP.n2 VSUBS 0.049011f
C705 VP.n3 VSUBS 0.054187f
C706 VP.t3 VSUBS 2.60479f
C707 VP.t2 VSUBS 2.99555f
C708 VP.t0 VSUBS 2.98447f
C709 VP.n4 VSUBS 3.70297f
C710 VP.n5 VSUBS 1.81865f
C711 VP.n6 VSUBS 1.07951f
C712 VP.n7 VSUBS 0.061644f
C713 VP.n8 VSUBS 0.062573f
C714 VP.n9 VSUBS 0.033574f
C715 VP.n10 VSUBS 0.033574f
C716 VP.n11 VSUBS 0.033574f
C717 VP.n12 VSUBS 0.049011f
C718 VP.n13 VSUBS 0.062573f
C719 VP.n14 VSUBS 0.061644f
C720 VP.n15 VSUBS 0.054187f
C721 VP.n16 VSUBS 0.064938f
.ends

