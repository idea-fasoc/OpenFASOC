* NGSPICE file created from diff_pair_sample_1303.ext - technology: sky130A

.subckt diff_pair_sample_1303 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=1.88265 ps=11.74 w=11.41 l=1.17
X1 VTAIL.t1 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X2 VDD1.t6 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=4.4499 ps=23.6 w=11.41 l=1.17
X3 VTAIL.t13 VN.t1 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X4 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=0 ps=0 w=11.41 l=1.17
X5 VTAIL.t0 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X6 VDD2.t2 VN.t2 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X7 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=0 ps=0 w=11.41 l=1.17
X8 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=4.4499 ps=23.6 w=11.41 l=1.17
X9 VTAIL.t5 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=1.88265 ps=11.74 w=11.41 l=1.17
X10 VDD2.t6 VN.t3 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=4.4499 ps=23.6 w=11.41 l=1.17
X11 VTAIL.t10 VN.t4 VDD2.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=1.88265 ps=11.74 w=11.41 l=1.17
X12 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=0 ps=0 w=11.41 l=1.17
X13 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=0 ps=0 w=11.41 l=1.17
X14 VTAIL.t9 VN.t5 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X15 VDD2.t1 VN.t6 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=4.4499 ps=23.6 w=11.41 l=1.17
X16 VDD2.t7 VN.t7 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X17 VTAIL.t15 VP.t5 VDD1.t2 B.t21 sky130_fd_pr__nfet_01v8 ad=4.4499 pd=23.6 as=1.88265 ps=11.74 w=11.41 l=1.17
X18 VDD1.t1 VP.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
X19 VDD1.t0 VP.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.88265 pd=11.74 as=1.88265 ps=11.74 w=11.41 l=1.17
R0 VN.n4 VN.t4 265.137
R1 VN.n22 VN.t3 265.137
R2 VN.n3 VN.t2 235.028
R3 VN.n8 VN.t1 235.028
R4 VN.n15 VN.t6 235.028
R5 VN.n21 VN.t5 235.028
R6 VN.n20 VN.t7 235.028
R7 VN.n32 VN.t0 235.028
R8 VN.n16 VN.n15 173.534
R9 VN.n33 VN.n32 173.534
R10 VN.n31 VN.n17 161.3
R11 VN.n30 VN.n29 161.3
R12 VN.n28 VN.n18 161.3
R13 VN.n27 VN.n26 161.3
R14 VN.n25 VN.n19 161.3
R15 VN.n24 VN.n23 161.3
R16 VN.n14 VN.n0 161.3
R17 VN.n13 VN.n12 161.3
R18 VN.n11 VN.n1 161.3
R19 VN.n10 VN.n9 161.3
R20 VN.n7 VN.n2 161.3
R21 VN.n6 VN.n5 161.3
R22 VN.n4 VN.n3 51.4127
R23 VN.n22 VN.n21 51.4127
R24 VN VN.n33 44.0175
R25 VN.n7 VN.n6 40.4934
R26 VN.n9 VN.n7 40.4934
R27 VN.n13 VN.n1 40.4934
R28 VN.n14 VN.n13 40.4934
R29 VN.n25 VN.n24 40.4934
R30 VN.n26 VN.n25 40.4934
R31 VN.n30 VN.n18 40.4934
R32 VN.n31 VN.n30 40.4934
R33 VN.n23 VN.n22 27.0291
R34 VN.n5 VN.n4 27.0291
R35 VN.n6 VN.n3 12.234
R36 VN.n9 VN.n8 12.234
R37 VN.n8 VN.n1 12.234
R38 VN.n15 VN.n14 12.234
R39 VN.n24 VN.n21 12.234
R40 VN.n20 VN.n18 12.234
R41 VN.n26 VN.n20 12.234
R42 VN.n32 VN.n31 12.234
R43 VN.n33 VN.n17 0.189894
R44 VN.n29 VN.n17 0.189894
R45 VN.n29 VN.n28 0.189894
R46 VN.n28 VN.n27 0.189894
R47 VN.n27 VN.n19 0.189894
R48 VN.n23 VN.n19 0.189894
R49 VN.n5 VN.n2 0.189894
R50 VN.n10 VN.n2 0.189894
R51 VN.n11 VN.n10 0.189894
R52 VN.n12 VN.n11 0.189894
R53 VN.n12 VN.n0 0.189894
R54 VN.n16 VN.n0 0.189894
R55 VN VN.n16 0.0516364
R56 VDD2.n2 VDD2.n1 62.8749
R57 VDD2.n2 VDD2.n0 62.8749
R58 VDD2 VDD2.n5 62.872
R59 VDD2.n4 VDD2.n3 62.2838
R60 VDD2.n4 VDD2.n2 39.3705
R61 VDD2.n5 VDD2.t4 1.73582
R62 VDD2.n5 VDD2.t6 1.73582
R63 VDD2.n3 VDD2.t0 1.73582
R64 VDD2.n3 VDD2.t7 1.73582
R65 VDD2.n1 VDD2.t3 1.73582
R66 VDD2.n1 VDD2.t1 1.73582
R67 VDD2.n0 VDD2.t5 1.73582
R68 VDD2.n0 VDD2.t2 1.73582
R69 VDD2 VDD2.n4 0.705241
R70 VTAIL.n498 VTAIL.n442 289.615
R71 VTAIL.n58 VTAIL.n2 289.615
R72 VTAIL.n120 VTAIL.n64 289.615
R73 VTAIL.n184 VTAIL.n128 289.615
R74 VTAIL.n436 VTAIL.n380 289.615
R75 VTAIL.n372 VTAIL.n316 289.615
R76 VTAIL.n310 VTAIL.n254 289.615
R77 VTAIL.n246 VTAIL.n190 289.615
R78 VTAIL.n463 VTAIL.n462 185
R79 VTAIL.n465 VTAIL.n464 185
R80 VTAIL.n458 VTAIL.n457 185
R81 VTAIL.n471 VTAIL.n470 185
R82 VTAIL.n473 VTAIL.n472 185
R83 VTAIL.n454 VTAIL.n453 185
R84 VTAIL.n480 VTAIL.n479 185
R85 VTAIL.n481 VTAIL.n452 185
R86 VTAIL.n483 VTAIL.n482 185
R87 VTAIL.n450 VTAIL.n449 185
R88 VTAIL.n489 VTAIL.n488 185
R89 VTAIL.n491 VTAIL.n490 185
R90 VTAIL.n446 VTAIL.n445 185
R91 VTAIL.n497 VTAIL.n496 185
R92 VTAIL.n499 VTAIL.n498 185
R93 VTAIL.n23 VTAIL.n22 185
R94 VTAIL.n25 VTAIL.n24 185
R95 VTAIL.n18 VTAIL.n17 185
R96 VTAIL.n31 VTAIL.n30 185
R97 VTAIL.n33 VTAIL.n32 185
R98 VTAIL.n14 VTAIL.n13 185
R99 VTAIL.n40 VTAIL.n39 185
R100 VTAIL.n41 VTAIL.n12 185
R101 VTAIL.n43 VTAIL.n42 185
R102 VTAIL.n10 VTAIL.n9 185
R103 VTAIL.n49 VTAIL.n48 185
R104 VTAIL.n51 VTAIL.n50 185
R105 VTAIL.n6 VTAIL.n5 185
R106 VTAIL.n57 VTAIL.n56 185
R107 VTAIL.n59 VTAIL.n58 185
R108 VTAIL.n85 VTAIL.n84 185
R109 VTAIL.n87 VTAIL.n86 185
R110 VTAIL.n80 VTAIL.n79 185
R111 VTAIL.n93 VTAIL.n92 185
R112 VTAIL.n95 VTAIL.n94 185
R113 VTAIL.n76 VTAIL.n75 185
R114 VTAIL.n102 VTAIL.n101 185
R115 VTAIL.n103 VTAIL.n74 185
R116 VTAIL.n105 VTAIL.n104 185
R117 VTAIL.n72 VTAIL.n71 185
R118 VTAIL.n111 VTAIL.n110 185
R119 VTAIL.n113 VTAIL.n112 185
R120 VTAIL.n68 VTAIL.n67 185
R121 VTAIL.n119 VTAIL.n118 185
R122 VTAIL.n121 VTAIL.n120 185
R123 VTAIL.n149 VTAIL.n148 185
R124 VTAIL.n151 VTAIL.n150 185
R125 VTAIL.n144 VTAIL.n143 185
R126 VTAIL.n157 VTAIL.n156 185
R127 VTAIL.n159 VTAIL.n158 185
R128 VTAIL.n140 VTAIL.n139 185
R129 VTAIL.n166 VTAIL.n165 185
R130 VTAIL.n167 VTAIL.n138 185
R131 VTAIL.n169 VTAIL.n168 185
R132 VTAIL.n136 VTAIL.n135 185
R133 VTAIL.n175 VTAIL.n174 185
R134 VTAIL.n177 VTAIL.n176 185
R135 VTAIL.n132 VTAIL.n131 185
R136 VTAIL.n183 VTAIL.n182 185
R137 VTAIL.n185 VTAIL.n184 185
R138 VTAIL.n437 VTAIL.n436 185
R139 VTAIL.n435 VTAIL.n434 185
R140 VTAIL.n384 VTAIL.n383 185
R141 VTAIL.n429 VTAIL.n428 185
R142 VTAIL.n427 VTAIL.n426 185
R143 VTAIL.n388 VTAIL.n387 185
R144 VTAIL.n392 VTAIL.n390 185
R145 VTAIL.n421 VTAIL.n420 185
R146 VTAIL.n419 VTAIL.n418 185
R147 VTAIL.n394 VTAIL.n393 185
R148 VTAIL.n413 VTAIL.n412 185
R149 VTAIL.n411 VTAIL.n410 185
R150 VTAIL.n398 VTAIL.n397 185
R151 VTAIL.n405 VTAIL.n404 185
R152 VTAIL.n403 VTAIL.n402 185
R153 VTAIL.n373 VTAIL.n372 185
R154 VTAIL.n371 VTAIL.n370 185
R155 VTAIL.n320 VTAIL.n319 185
R156 VTAIL.n365 VTAIL.n364 185
R157 VTAIL.n363 VTAIL.n362 185
R158 VTAIL.n324 VTAIL.n323 185
R159 VTAIL.n328 VTAIL.n326 185
R160 VTAIL.n357 VTAIL.n356 185
R161 VTAIL.n355 VTAIL.n354 185
R162 VTAIL.n330 VTAIL.n329 185
R163 VTAIL.n349 VTAIL.n348 185
R164 VTAIL.n347 VTAIL.n346 185
R165 VTAIL.n334 VTAIL.n333 185
R166 VTAIL.n341 VTAIL.n340 185
R167 VTAIL.n339 VTAIL.n338 185
R168 VTAIL.n311 VTAIL.n310 185
R169 VTAIL.n309 VTAIL.n308 185
R170 VTAIL.n258 VTAIL.n257 185
R171 VTAIL.n303 VTAIL.n302 185
R172 VTAIL.n301 VTAIL.n300 185
R173 VTAIL.n262 VTAIL.n261 185
R174 VTAIL.n266 VTAIL.n264 185
R175 VTAIL.n295 VTAIL.n294 185
R176 VTAIL.n293 VTAIL.n292 185
R177 VTAIL.n268 VTAIL.n267 185
R178 VTAIL.n287 VTAIL.n286 185
R179 VTAIL.n285 VTAIL.n284 185
R180 VTAIL.n272 VTAIL.n271 185
R181 VTAIL.n279 VTAIL.n278 185
R182 VTAIL.n277 VTAIL.n276 185
R183 VTAIL.n247 VTAIL.n246 185
R184 VTAIL.n245 VTAIL.n244 185
R185 VTAIL.n194 VTAIL.n193 185
R186 VTAIL.n239 VTAIL.n238 185
R187 VTAIL.n237 VTAIL.n236 185
R188 VTAIL.n198 VTAIL.n197 185
R189 VTAIL.n202 VTAIL.n200 185
R190 VTAIL.n231 VTAIL.n230 185
R191 VTAIL.n229 VTAIL.n228 185
R192 VTAIL.n204 VTAIL.n203 185
R193 VTAIL.n223 VTAIL.n222 185
R194 VTAIL.n221 VTAIL.n220 185
R195 VTAIL.n208 VTAIL.n207 185
R196 VTAIL.n215 VTAIL.n214 185
R197 VTAIL.n213 VTAIL.n212 185
R198 VTAIL.n461 VTAIL.t8 149.524
R199 VTAIL.n21 VTAIL.t10 149.524
R200 VTAIL.n83 VTAIL.t6 149.524
R201 VTAIL.n147 VTAIL.t5 149.524
R202 VTAIL.n401 VTAIL.t3 149.524
R203 VTAIL.n337 VTAIL.t15 149.524
R204 VTAIL.n275 VTAIL.t11 149.524
R205 VTAIL.n211 VTAIL.t14 149.524
R206 VTAIL.n464 VTAIL.n463 104.615
R207 VTAIL.n464 VTAIL.n457 104.615
R208 VTAIL.n471 VTAIL.n457 104.615
R209 VTAIL.n472 VTAIL.n471 104.615
R210 VTAIL.n472 VTAIL.n453 104.615
R211 VTAIL.n480 VTAIL.n453 104.615
R212 VTAIL.n481 VTAIL.n480 104.615
R213 VTAIL.n482 VTAIL.n481 104.615
R214 VTAIL.n482 VTAIL.n449 104.615
R215 VTAIL.n489 VTAIL.n449 104.615
R216 VTAIL.n490 VTAIL.n489 104.615
R217 VTAIL.n490 VTAIL.n445 104.615
R218 VTAIL.n497 VTAIL.n445 104.615
R219 VTAIL.n498 VTAIL.n497 104.615
R220 VTAIL.n24 VTAIL.n23 104.615
R221 VTAIL.n24 VTAIL.n17 104.615
R222 VTAIL.n31 VTAIL.n17 104.615
R223 VTAIL.n32 VTAIL.n31 104.615
R224 VTAIL.n32 VTAIL.n13 104.615
R225 VTAIL.n40 VTAIL.n13 104.615
R226 VTAIL.n41 VTAIL.n40 104.615
R227 VTAIL.n42 VTAIL.n41 104.615
R228 VTAIL.n42 VTAIL.n9 104.615
R229 VTAIL.n49 VTAIL.n9 104.615
R230 VTAIL.n50 VTAIL.n49 104.615
R231 VTAIL.n50 VTAIL.n5 104.615
R232 VTAIL.n57 VTAIL.n5 104.615
R233 VTAIL.n58 VTAIL.n57 104.615
R234 VTAIL.n86 VTAIL.n85 104.615
R235 VTAIL.n86 VTAIL.n79 104.615
R236 VTAIL.n93 VTAIL.n79 104.615
R237 VTAIL.n94 VTAIL.n93 104.615
R238 VTAIL.n94 VTAIL.n75 104.615
R239 VTAIL.n102 VTAIL.n75 104.615
R240 VTAIL.n103 VTAIL.n102 104.615
R241 VTAIL.n104 VTAIL.n103 104.615
R242 VTAIL.n104 VTAIL.n71 104.615
R243 VTAIL.n111 VTAIL.n71 104.615
R244 VTAIL.n112 VTAIL.n111 104.615
R245 VTAIL.n112 VTAIL.n67 104.615
R246 VTAIL.n119 VTAIL.n67 104.615
R247 VTAIL.n120 VTAIL.n119 104.615
R248 VTAIL.n150 VTAIL.n149 104.615
R249 VTAIL.n150 VTAIL.n143 104.615
R250 VTAIL.n157 VTAIL.n143 104.615
R251 VTAIL.n158 VTAIL.n157 104.615
R252 VTAIL.n158 VTAIL.n139 104.615
R253 VTAIL.n166 VTAIL.n139 104.615
R254 VTAIL.n167 VTAIL.n166 104.615
R255 VTAIL.n168 VTAIL.n167 104.615
R256 VTAIL.n168 VTAIL.n135 104.615
R257 VTAIL.n175 VTAIL.n135 104.615
R258 VTAIL.n176 VTAIL.n175 104.615
R259 VTAIL.n176 VTAIL.n131 104.615
R260 VTAIL.n183 VTAIL.n131 104.615
R261 VTAIL.n184 VTAIL.n183 104.615
R262 VTAIL.n436 VTAIL.n435 104.615
R263 VTAIL.n435 VTAIL.n383 104.615
R264 VTAIL.n428 VTAIL.n383 104.615
R265 VTAIL.n428 VTAIL.n427 104.615
R266 VTAIL.n427 VTAIL.n387 104.615
R267 VTAIL.n392 VTAIL.n387 104.615
R268 VTAIL.n420 VTAIL.n392 104.615
R269 VTAIL.n420 VTAIL.n419 104.615
R270 VTAIL.n419 VTAIL.n393 104.615
R271 VTAIL.n412 VTAIL.n393 104.615
R272 VTAIL.n412 VTAIL.n411 104.615
R273 VTAIL.n411 VTAIL.n397 104.615
R274 VTAIL.n404 VTAIL.n397 104.615
R275 VTAIL.n404 VTAIL.n403 104.615
R276 VTAIL.n372 VTAIL.n371 104.615
R277 VTAIL.n371 VTAIL.n319 104.615
R278 VTAIL.n364 VTAIL.n319 104.615
R279 VTAIL.n364 VTAIL.n363 104.615
R280 VTAIL.n363 VTAIL.n323 104.615
R281 VTAIL.n328 VTAIL.n323 104.615
R282 VTAIL.n356 VTAIL.n328 104.615
R283 VTAIL.n356 VTAIL.n355 104.615
R284 VTAIL.n355 VTAIL.n329 104.615
R285 VTAIL.n348 VTAIL.n329 104.615
R286 VTAIL.n348 VTAIL.n347 104.615
R287 VTAIL.n347 VTAIL.n333 104.615
R288 VTAIL.n340 VTAIL.n333 104.615
R289 VTAIL.n340 VTAIL.n339 104.615
R290 VTAIL.n310 VTAIL.n309 104.615
R291 VTAIL.n309 VTAIL.n257 104.615
R292 VTAIL.n302 VTAIL.n257 104.615
R293 VTAIL.n302 VTAIL.n301 104.615
R294 VTAIL.n301 VTAIL.n261 104.615
R295 VTAIL.n266 VTAIL.n261 104.615
R296 VTAIL.n294 VTAIL.n266 104.615
R297 VTAIL.n294 VTAIL.n293 104.615
R298 VTAIL.n293 VTAIL.n267 104.615
R299 VTAIL.n286 VTAIL.n267 104.615
R300 VTAIL.n286 VTAIL.n285 104.615
R301 VTAIL.n285 VTAIL.n271 104.615
R302 VTAIL.n278 VTAIL.n271 104.615
R303 VTAIL.n278 VTAIL.n277 104.615
R304 VTAIL.n246 VTAIL.n245 104.615
R305 VTAIL.n245 VTAIL.n193 104.615
R306 VTAIL.n238 VTAIL.n193 104.615
R307 VTAIL.n238 VTAIL.n237 104.615
R308 VTAIL.n237 VTAIL.n197 104.615
R309 VTAIL.n202 VTAIL.n197 104.615
R310 VTAIL.n230 VTAIL.n202 104.615
R311 VTAIL.n230 VTAIL.n229 104.615
R312 VTAIL.n229 VTAIL.n203 104.615
R313 VTAIL.n222 VTAIL.n203 104.615
R314 VTAIL.n222 VTAIL.n221 104.615
R315 VTAIL.n221 VTAIL.n207 104.615
R316 VTAIL.n214 VTAIL.n207 104.615
R317 VTAIL.n214 VTAIL.n213 104.615
R318 VTAIL.n463 VTAIL.t8 52.3082
R319 VTAIL.n23 VTAIL.t10 52.3082
R320 VTAIL.n85 VTAIL.t6 52.3082
R321 VTAIL.n149 VTAIL.t5 52.3082
R322 VTAIL.n403 VTAIL.t3 52.3082
R323 VTAIL.n339 VTAIL.t15 52.3082
R324 VTAIL.n277 VTAIL.t11 52.3082
R325 VTAIL.n213 VTAIL.t14 52.3082
R326 VTAIL.n379 VTAIL.n378 45.6051
R327 VTAIL.n253 VTAIL.n252 45.6051
R328 VTAIL.n1 VTAIL.n0 45.6049
R329 VTAIL.n127 VTAIL.n126 45.6049
R330 VTAIL.n503 VTAIL.n502 32.3793
R331 VTAIL.n63 VTAIL.n62 32.3793
R332 VTAIL.n125 VTAIL.n124 32.3793
R333 VTAIL.n189 VTAIL.n188 32.3793
R334 VTAIL.n441 VTAIL.n440 32.3793
R335 VTAIL.n377 VTAIL.n376 32.3793
R336 VTAIL.n315 VTAIL.n314 32.3793
R337 VTAIL.n251 VTAIL.n250 32.3793
R338 VTAIL.n503 VTAIL.n441 23.4962
R339 VTAIL.n251 VTAIL.n189 23.4962
R340 VTAIL.n483 VTAIL.n450 13.1884
R341 VTAIL.n43 VTAIL.n10 13.1884
R342 VTAIL.n105 VTAIL.n72 13.1884
R343 VTAIL.n169 VTAIL.n136 13.1884
R344 VTAIL.n390 VTAIL.n388 13.1884
R345 VTAIL.n326 VTAIL.n324 13.1884
R346 VTAIL.n264 VTAIL.n262 13.1884
R347 VTAIL.n200 VTAIL.n198 13.1884
R348 VTAIL.n484 VTAIL.n452 12.8005
R349 VTAIL.n488 VTAIL.n487 12.8005
R350 VTAIL.n44 VTAIL.n12 12.8005
R351 VTAIL.n48 VTAIL.n47 12.8005
R352 VTAIL.n106 VTAIL.n74 12.8005
R353 VTAIL.n110 VTAIL.n109 12.8005
R354 VTAIL.n170 VTAIL.n138 12.8005
R355 VTAIL.n174 VTAIL.n173 12.8005
R356 VTAIL.n426 VTAIL.n425 12.8005
R357 VTAIL.n422 VTAIL.n421 12.8005
R358 VTAIL.n362 VTAIL.n361 12.8005
R359 VTAIL.n358 VTAIL.n357 12.8005
R360 VTAIL.n300 VTAIL.n299 12.8005
R361 VTAIL.n296 VTAIL.n295 12.8005
R362 VTAIL.n236 VTAIL.n235 12.8005
R363 VTAIL.n232 VTAIL.n231 12.8005
R364 VTAIL.n479 VTAIL.n478 12.0247
R365 VTAIL.n491 VTAIL.n448 12.0247
R366 VTAIL.n39 VTAIL.n38 12.0247
R367 VTAIL.n51 VTAIL.n8 12.0247
R368 VTAIL.n101 VTAIL.n100 12.0247
R369 VTAIL.n113 VTAIL.n70 12.0247
R370 VTAIL.n165 VTAIL.n164 12.0247
R371 VTAIL.n177 VTAIL.n134 12.0247
R372 VTAIL.n429 VTAIL.n386 12.0247
R373 VTAIL.n418 VTAIL.n391 12.0247
R374 VTAIL.n365 VTAIL.n322 12.0247
R375 VTAIL.n354 VTAIL.n327 12.0247
R376 VTAIL.n303 VTAIL.n260 12.0247
R377 VTAIL.n292 VTAIL.n265 12.0247
R378 VTAIL.n239 VTAIL.n196 12.0247
R379 VTAIL.n228 VTAIL.n201 12.0247
R380 VTAIL.n477 VTAIL.n454 11.249
R381 VTAIL.n492 VTAIL.n446 11.249
R382 VTAIL.n37 VTAIL.n14 11.249
R383 VTAIL.n52 VTAIL.n6 11.249
R384 VTAIL.n99 VTAIL.n76 11.249
R385 VTAIL.n114 VTAIL.n68 11.249
R386 VTAIL.n163 VTAIL.n140 11.249
R387 VTAIL.n178 VTAIL.n132 11.249
R388 VTAIL.n430 VTAIL.n384 11.249
R389 VTAIL.n417 VTAIL.n394 11.249
R390 VTAIL.n366 VTAIL.n320 11.249
R391 VTAIL.n353 VTAIL.n330 11.249
R392 VTAIL.n304 VTAIL.n258 11.249
R393 VTAIL.n291 VTAIL.n268 11.249
R394 VTAIL.n240 VTAIL.n194 11.249
R395 VTAIL.n227 VTAIL.n204 11.249
R396 VTAIL.n474 VTAIL.n473 10.4732
R397 VTAIL.n496 VTAIL.n495 10.4732
R398 VTAIL.n34 VTAIL.n33 10.4732
R399 VTAIL.n56 VTAIL.n55 10.4732
R400 VTAIL.n96 VTAIL.n95 10.4732
R401 VTAIL.n118 VTAIL.n117 10.4732
R402 VTAIL.n160 VTAIL.n159 10.4732
R403 VTAIL.n182 VTAIL.n181 10.4732
R404 VTAIL.n434 VTAIL.n433 10.4732
R405 VTAIL.n414 VTAIL.n413 10.4732
R406 VTAIL.n370 VTAIL.n369 10.4732
R407 VTAIL.n350 VTAIL.n349 10.4732
R408 VTAIL.n308 VTAIL.n307 10.4732
R409 VTAIL.n288 VTAIL.n287 10.4732
R410 VTAIL.n244 VTAIL.n243 10.4732
R411 VTAIL.n224 VTAIL.n223 10.4732
R412 VTAIL.n462 VTAIL.n461 10.2747
R413 VTAIL.n22 VTAIL.n21 10.2747
R414 VTAIL.n84 VTAIL.n83 10.2747
R415 VTAIL.n148 VTAIL.n147 10.2747
R416 VTAIL.n402 VTAIL.n401 10.2747
R417 VTAIL.n338 VTAIL.n337 10.2747
R418 VTAIL.n276 VTAIL.n275 10.2747
R419 VTAIL.n212 VTAIL.n211 10.2747
R420 VTAIL.n470 VTAIL.n456 9.69747
R421 VTAIL.n499 VTAIL.n444 9.69747
R422 VTAIL.n30 VTAIL.n16 9.69747
R423 VTAIL.n59 VTAIL.n4 9.69747
R424 VTAIL.n92 VTAIL.n78 9.69747
R425 VTAIL.n121 VTAIL.n66 9.69747
R426 VTAIL.n156 VTAIL.n142 9.69747
R427 VTAIL.n185 VTAIL.n130 9.69747
R428 VTAIL.n437 VTAIL.n382 9.69747
R429 VTAIL.n410 VTAIL.n396 9.69747
R430 VTAIL.n373 VTAIL.n318 9.69747
R431 VTAIL.n346 VTAIL.n332 9.69747
R432 VTAIL.n311 VTAIL.n256 9.69747
R433 VTAIL.n284 VTAIL.n270 9.69747
R434 VTAIL.n247 VTAIL.n192 9.69747
R435 VTAIL.n220 VTAIL.n206 9.69747
R436 VTAIL.n502 VTAIL.n501 9.45567
R437 VTAIL.n62 VTAIL.n61 9.45567
R438 VTAIL.n124 VTAIL.n123 9.45567
R439 VTAIL.n188 VTAIL.n187 9.45567
R440 VTAIL.n440 VTAIL.n439 9.45567
R441 VTAIL.n376 VTAIL.n375 9.45567
R442 VTAIL.n314 VTAIL.n313 9.45567
R443 VTAIL.n250 VTAIL.n249 9.45567
R444 VTAIL.n501 VTAIL.n500 9.3005
R445 VTAIL.n444 VTAIL.n443 9.3005
R446 VTAIL.n495 VTAIL.n494 9.3005
R447 VTAIL.n493 VTAIL.n492 9.3005
R448 VTAIL.n448 VTAIL.n447 9.3005
R449 VTAIL.n487 VTAIL.n486 9.3005
R450 VTAIL.n460 VTAIL.n459 9.3005
R451 VTAIL.n467 VTAIL.n466 9.3005
R452 VTAIL.n469 VTAIL.n468 9.3005
R453 VTAIL.n456 VTAIL.n455 9.3005
R454 VTAIL.n475 VTAIL.n474 9.3005
R455 VTAIL.n477 VTAIL.n476 9.3005
R456 VTAIL.n478 VTAIL.n451 9.3005
R457 VTAIL.n485 VTAIL.n484 9.3005
R458 VTAIL.n61 VTAIL.n60 9.3005
R459 VTAIL.n4 VTAIL.n3 9.3005
R460 VTAIL.n55 VTAIL.n54 9.3005
R461 VTAIL.n53 VTAIL.n52 9.3005
R462 VTAIL.n8 VTAIL.n7 9.3005
R463 VTAIL.n47 VTAIL.n46 9.3005
R464 VTAIL.n20 VTAIL.n19 9.3005
R465 VTAIL.n27 VTAIL.n26 9.3005
R466 VTAIL.n29 VTAIL.n28 9.3005
R467 VTAIL.n16 VTAIL.n15 9.3005
R468 VTAIL.n35 VTAIL.n34 9.3005
R469 VTAIL.n37 VTAIL.n36 9.3005
R470 VTAIL.n38 VTAIL.n11 9.3005
R471 VTAIL.n45 VTAIL.n44 9.3005
R472 VTAIL.n123 VTAIL.n122 9.3005
R473 VTAIL.n66 VTAIL.n65 9.3005
R474 VTAIL.n117 VTAIL.n116 9.3005
R475 VTAIL.n115 VTAIL.n114 9.3005
R476 VTAIL.n70 VTAIL.n69 9.3005
R477 VTAIL.n109 VTAIL.n108 9.3005
R478 VTAIL.n82 VTAIL.n81 9.3005
R479 VTAIL.n89 VTAIL.n88 9.3005
R480 VTAIL.n91 VTAIL.n90 9.3005
R481 VTAIL.n78 VTAIL.n77 9.3005
R482 VTAIL.n97 VTAIL.n96 9.3005
R483 VTAIL.n99 VTAIL.n98 9.3005
R484 VTAIL.n100 VTAIL.n73 9.3005
R485 VTAIL.n107 VTAIL.n106 9.3005
R486 VTAIL.n187 VTAIL.n186 9.3005
R487 VTAIL.n130 VTAIL.n129 9.3005
R488 VTAIL.n181 VTAIL.n180 9.3005
R489 VTAIL.n179 VTAIL.n178 9.3005
R490 VTAIL.n134 VTAIL.n133 9.3005
R491 VTAIL.n173 VTAIL.n172 9.3005
R492 VTAIL.n146 VTAIL.n145 9.3005
R493 VTAIL.n153 VTAIL.n152 9.3005
R494 VTAIL.n155 VTAIL.n154 9.3005
R495 VTAIL.n142 VTAIL.n141 9.3005
R496 VTAIL.n161 VTAIL.n160 9.3005
R497 VTAIL.n163 VTAIL.n162 9.3005
R498 VTAIL.n164 VTAIL.n137 9.3005
R499 VTAIL.n171 VTAIL.n170 9.3005
R500 VTAIL.n400 VTAIL.n399 9.3005
R501 VTAIL.n407 VTAIL.n406 9.3005
R502 VTAIL.n409 VTAIL.n408 9.3005
R503 VTAIL.n396 VTAIL.n395 9.3005
R504 VTAIL.n415 VTAIL.n414 9.3005
R505 VTAIL.n417 VTAIL.n416 9.3005
R506 VTAIL.n391 VTAIL.n389 9.3005
R507 VTAIL.n423 VTAIL.n422 9.3005
R508 VTAIL.n439 VTAIL.n438 9.3005
R509 VTAIL.n382 VTAIL.n381 9.3005
R510 VTAIL.n433 VTAIL.n432 9.3005
R511 VTAIL.n431 VTAIL.n430 9.3005
R512 VTAIL.n386 VTAIL.n385 9.3005
R513 VTAIL.n425 VTAIL.n424 9.3005
R514 VTAIL.n336 VTAIL.n335 9.3005
R515 VTAIL.n343 VTAIL.n342 9.3005
R516 VTAIL.n345 VTAIL.n344 9.3005
R517 VTAIL.n332 VTAIL.n331 9.3005
R518 VTAIL.n351 VTAIL.n350 9.3005
R519 VTAIL.n353 VTAIL.n352 9.3005
R520 VTAIL.n327 VTAIL.n325 9.3005
R521 VTAIL.n359 VTAIL.n358 9.3005
R522 VTAIL.n375 VTAIL.n374 9.3005
R523 VTAIL.n318 VTAIL.n317 9.3005
R524 VTAIL.n369 VTAIL.n368 9.3005
R525 VTAIL.n367 VTAIL.n366 9.3005
R526 VTAIL.n322 VTAIL.n321 9.3005
R527 VTAIL.n361 VTAIL.n360 9.3005
R528 VTAIL.n274 VTAIL.n273 9.3005
R529 VTAIL.n281 VTAIL.n280 9.3005
R530 VTAIL.n283 VTAIL.n282 9.3005
R531 VTAIL.n270 VTAIL.n269 9.3005
R532 VTAIL.n289 VTAIL.n288 9.3005
R533 VTAIL.n291 VTAIL.n290 9.3005
R534 VTAIL.n265 VTAIL.n263 9.3005
R535 VTAIL.n297 VTAIL.n296 9.3005
R536 VTAIL.n313 VTAIL.n312 9.3005
R537 VTAIL.n256 VTAIL.n255 9.3005
R538 VTAIL.n307 VTAIL.n306 9.3005
R539 VTAIL.n305 VTAIL.n304 9.3005
R540 VTAIL.n260 VTAIL.n259 9.3005
R541 VTAIL.n299 VTAIL.n298 9.3005
R542 VTAIL.n210 VTAIL.n209 9.3005
R543 VTAIL.n217 VTAIL.n216 9.3005
R544 VTAIL.n219 VTAIL.n218 9.3005
R545 VTAIL.n206 VTAIL.n205 9.3005
R546 VTAIL.n225 VTAIL.n224 9.3005
R547 VTAIL.n227 VTAIL.n226 9.3005
R548 VTAIL.n201 VTAIL.n199 9.3005
R549 VTAIL.n233 VTAIL.n232 9.3005
R550 VTAIL.n249 VTAIL.n248 9.3005
R551 VTAIL.n192 VTAIL.n191 9.3005
R552 VTAIL.n243 VTAIL.n242 9.3005
R553 VTAIL.n241 VTAIL.n240 9.3005
R554 VTAIL.n196 VTAIL.n195 9.3005
R555 VTAIL.n235 VTAIL.n234 9.3005
R556 VTAIL.n469 VTAIL.n458 8.92171
R557 VTAIL.n500 VTAIL.n442 8.92171
R558 VTAIL.n29 VTAIL.n18 8.92171
R559 VTAIL.n60 VTAIL.n2 8.92171
R560 VTAIL.n91 VTAIL.n80 8.92171
R561 VTAIL.n122 VTAIL.n64 8.92171
R562 VTAIL.n155 VTAIL.n144 8.92171
R563 VTAIL.n186 VTAIL.n128 8.92171
R564 VTAIL.n438 VTAIL.n380 8.92171
R565 VTAIL.n409 VTAIL.n398 8.92171
R566 VTAIL.n374 VTAIL.n316 8.92171
R567 VTAIL.n345 VTAIL.n334 8.92171
R568 VTAIL.n312 VTAIL.n254 8.92171
R569 VTAIL.n283 VTAIL.n272 8.92171
R570 VTAIL.n248 VTAIL.n190 8.92171
R571 VTAIL.n219 VTAIL.n208 8.92171
R572 VTAIL.n466 VTAIL.n465 8.14595
R573 VTAIL.n26 VTAIL.n25 8.14595
R574 VTAIL.n88 VTAIL.n87 8.14595
R575 VTAIL.n152 VTAIL.n151 8.14595
R576 VTAIL.n406 VTAIL.n405 8.14595
R577 VTAIL.n342 VTAIL.n341 8.14595
R578 VTAIL.n280 VTAIL.n279 8.14595
R579 VTAIL.n216 VTAIL.n215 8.14595
R580 VTAIL.n462 VTAIL.n460 7.3702
R581 VTAIL.n22 VTAIL.n20 7.3702
R582 VTAIL.n84 VTAIL.n82 7.3702
R583 VTAIL.n148 VTAIL.n146 7.3702
R584 VTAIL.n402 VTAIL.n400 7.3702
R585 VTAIL.n338 VTAIL.n336 7.3702
R586 VTAIL.n276 VTAIL.n274 7.3702
R587 VTAIL.n212 VTAIL.n210 7.3702
R588 VTAIL.n465 VTAIL.n460 5.81868
R589 VTAIL.n25 VTAIL.n20 5.81868
R590 VTAIL.n87 VTAIL.n82 5.81868
R591 VTAIL.n151 VTAIL.n146 5.81868
R592 VTAIL.n405 VTAIL.n400 5.81868
R593 VTAIL.n341 VTAIL.n336 5.81868
R594 VTAIL.n279 VTAIL.n274 5.81868
R595 VTAIL.n215 VTAIL.n210 5.81868
R596 VTAIL.n466 VTAIL.n458 5.04292
R597 VTAIL.n502 VTAIL.n442 5.04292
R598 VTAIL.n26 VTAIL.n18 5.04292
R599 VTAIL.n62 VTAIL.n2 5.04292
R600 VTAIL.n88 VTAIL.n80 5.04292
R601 VTAIL.n124 VTAIL.n64 5.04292
R602 VTAIL.n152 VTAIL.n144 5.04292
R603 VTAIL.n188 VTAIL.n128 5.04292
R604 VTAIL.n440 VTAIL.n380 5.04292
R605 VTAIL.n406 VTAIL.n398 5.04292
R606 VTAIL.n376 VTAIL.n316 5.04292
R607 VTAIL.n342 VTAIL.n334 5.04292
R608 VTAIL.n314 VTAIL.n254 5.04292
R609 VTAIL.n280 VTAIL.n272 5.04292
R610 VTAIL.n250 VTAIL.n190 5.04292
R611 VTAIL.n216 VTAIL.n208 5.04292
R612 VTAIL.n470 VTAIL.n469 4.26717
R613 VTAIL.n500 VTAIL.n499 4.26717
R614 VTAIL.n30 VTAIL.n29 4.26717
R615 VTAIL.n60 VTAIL.n59 4.26717
R616 VTAIL.n92 VTAIL.n91 4.26717
R617 VTAIL.n122 VTAIL.n121 4.26717
R618 VTAIL.n156 VTAIL.n155 4.26717
R619 VTAIL.n186 VTAIL.n185 4.26717
R620 VTAIL.n438 VTAIL.n437 4.26717
R621 VTAIL.n410 VTAIL.n409 4.26717
R622 VTAIL.n374 VTAIL.n373 4.26717
R623 VTAIL.n346 VTAIL.n345 4.26717
R624 VTAIL.n312 VTAIL.n311 4.26717
R625 VTAIL.n284 VTAIL.n283 4.26717
R626 VTAIL.n248 VTAIL.n247 4.26717
R627 VTAIL.n220 VTAIL.n219 4.26717
R628 VTAIL.n473 VTAIL.n456 3.49141
R629 VTAIL.n496 VTAIL.n444 3.49141
R630 VTAIL.n33 VTAIL.n16 3.49141
R631 VTAIL.n56 VTAIL.n4 3.49141
R632 VTAIL.n95 VTAIL.n78 3.49141
R633 VTAIL.n118 VTAIL.n66 3.49141
R634 VTAIL.n159 VTAIL.n142 3.49141
R635 VTAIL.n182 VTAIL.n130 3.49141
R636 VTAIL.n434 VTAIL.n382 3.49141
R637 VTAIL.n413 VTAIL.n396 3.49141
R638 VTAIL.n370 VTAIL.n318 3.49141
R639 VTAIL.n349 VTAIL.n332 3.49141
R640 VTAIL.n308 VTAIL.n256 3.49141
R641 VTAIL.n287 VTAIL.n270 3.49141
R642 VTAIL.n244 VTAIL.n192 3.49141
R643 VTAIL.n223 VTAIL.n206 3.49141
R644 VTAIL.n461 VTAIL.n459 2.84303
R645 VTAIL.n21 VTAIL.n19 2.84303
R646 VTAIL.n83 VTAIL.n81 2.84303
R647 VTAIL.n147 VTAIL.n145 2.84303
R648 VTAIL.n401 VTAIL.n399 2.84303
R649 VTAIL.n337 VTAIL.n335 2.84303
R650 VTAIL.n275 VTAIL.n273 2.84303
R651 VTAIL.n211 VTAIL.n209 2.84303
R652 VTAIL.n474 VTAIL.n454 2.71565
R653 VTAIL.n495 VTAIL.n446 2.71565
R654 VTAIL.n34 VTAIL.n14 2.71565
R655 VTAIL.n55 VTAIL.n6 2.71565
R656 VTAIL.n96 VTAIL.n76 2.71565
R657 VTAIL.n117 VTAIL.n68 2.71565
R658 VTAIL.n160 VTAIL.n140 2.71565
R659 VTAIL.n181 VTAIL.n132 2.71565
R660 VTAIL.n433 VTAIL.n384 2.71565
R661 VTAIL.n414 VTAIL.n394 2.71565
R662 VTAIL.n369 VTAIL.n320 2.71565
R663 VTAIL.n350 VTAIL.n330 2.71565
R664 VTAIL.n307 VTAIL.n258 2.71565
R665 VTAIL.n288 VTAIL.n268 2.71565
R666 VTAIL.n243 VTAIL.n194 2.71565
R667 VTAIL.n224 VTAIL.n204 2.71565
R668 VTAIL.n479 VTAIL.n477 1.93989
R669 VTAIL.n492 VTAIL.n491 1.93989
R670 VTAIL.n39 VTAIL.n37 1.93989
R671 VTAIL.n52 VTAIL.n51 1.93989
R672 VTAIL.n101 VTAIL.n99 1.93989
R673 VTAIL.n114 VTAIL.n113 1.93989
R674 VTAIL.n165 VTAIL.n163 1.93989
R675 VTAIL.n178 VTAIL.n177 1.93989
R676 VTAIL.n430 VTAIL.n429 1.93989
R677 VTAIL.n418 VTAIL.n417 1.93989
R678 VTAIL.n366 VTAIL.n365 1.93989
R679 VTAIL.n354 VTAIL.n353 1.93989
R680 VTAIL.n304 VTAIL.n303 1.93989
R681 VTAIL.n292 VTAIL.n291 1.93989
R682 VTAIL.n240 VTAIL.n239 1.93989
R683 VTAIL.n228 VTAIL.n227 1.93989
R684 VTAIL.n0 VTAIL.t12 1.73582
R685 VTAIL.n0 VTAIL.t13 1.73582
R686 VTAIL.n126 VTAIL.t2 1.73582
R687 VTAIL.n126 VTAIL.t0 1.73582
R688 VTAIL.n378 VTAIL.t4 1.73582
R689 VTAIL.n378 VTAIL.t1 1.73582
R690 VTAIL.n252 VTAIL.t7 1.73582
R691 VTAIL.n252 VTAIL.t9 1.73582
R692 VTAIL.n253 VTAIL.n251 1.2936
R693 VTAIL.n315 VTAIL.n253 1.2936
R694 VTAIL.n379 VTAIL.n377 1.2936
R695 VTAIL.n441 VTAIL.n379 1.2936
R696 VTAIL.n189 VTAIL.n127 1.2936
R697 VTAIL.n127 VTAIL.n125 1.2936
R698 VTAIL.n63 VTAIL.n1 1.2936
R699 VTAIL VTAIL.n503 1.23541
R700 VTAIL.n478 VTAIL.n452 1.16414
R701 VTAIL.n488 VTAIL.n448 1.16414
R702 VTAIL.n38 VTAIL.n12 1.16414
R703 VTAIL.n48 VTAIL.n8 1.16414
R704 VTAIL.n100 VTAIL.n74 1.16414
R705 VTAIL.n110 VTAIL.n70 1.16414
R706 VTAIL.n164 VTAIL.n138 1.16414
R707 VTAIL.n174 VTAIL.n134 1.16414
R708 VTAIL.n426 VTAIL.n386 1.16414
R709 VTAIL.n421 VTAIL.n391 1.16414
R710 VTAIL.n362 VTAIL.n322 1.16414
R711 VTAIL.n357 VTAIL.n327 1.16414
R712 VTAIL.n300 VTAIL.n260 1.16414
R713 VTAIL.n295 VTAIL.n265 1.16414
R714 VTAIL.n236 VTAIL.n196 1.16414
R715 VTAIL.n231 VTAIL.n201 1.16414
R716 VTAIL.n377 VTAIL.n315 0.470328
R717 VTAIL.n125 VTAIL.n63 0.470328
R718 VTAIL.n484 VTAIL.n483 0.388379
R719 VTAIL.n487 VTAIL.n450 0.388379
R720 VTAIL.n44 VTAIL.n43 0.388379
R721 VTAIL.n47 VTAIL.n10 0.388379
R722 VTAIL.n106 VTAIL.n105 0.388379
R723 VTAIL.n109 VTAIL.n72 0.388379
R724 VTAIL.n170 VTAIL.n169 0.388379
R725 VTAIL.n173 VTAIL.n136 0.388379
R726 VTAIL.n425 VTAIL.n388 0.388379
R727 VTAIL.n422 VTAIL.n390 0.388379
R728 VTAIL.n361 VTAIL.n324 0.388379
R729 VTAIL.n358 VTAIL.n326 0.388379
R730 VTAIL.n299 VTAIL.n262 0.388379
R731 VTAIL.n296 VTAIL.n264 0.388379
R732 VTAIL.n235 VTAIL.n198 0.388379
R733 VTAIL.n232 VTAIL.n200 0.388379
R734 VTAIL.n467 VTAIL.n459 0.155672
R735 VTAIL.n468 VTAIL.n467 0.155672
R736 VTAIL.n468 VTAIL.n455 0.155672
R737 VTAIL.n475 VTAIL.n455 0.155672
R738 VTAIL.n476 VTAIL.n475 0.155672
R739 VTAIL.n476 VTAIL.n451 0.155672
R740 VTAIL.n485 VTAIL.n451 0.155672
R741 VTAIL.n486 VTAIL.n485 0.155672
R742 VTAIL.n486 VTAIL.n447 0.155672
R743 VTAIL.n493 VTAIL.n447 0.155672
R744 VTAIL.n494 VTAIL.n493 0.155672
R745 VTAIL.n494 VTAIL.n443 0.155672
R746 VTAIL.n501 VTAIL.n443 0.155672
R747 VTAIL.n27 VTAIL.n19 0.155672
R748 VTAIL.n28 VTAIL.n27 0.155672
R749 VTAIL.n28 VTAIL.n15 0.155672
R750 VTAIL.n35 VTAIL.n15 0.155672
R751 VTAIL.n36 VTAIL.n35 0.155672
R752 VTAIL.n36 VTAIL.n11 0.155672
R753 VTAIL.n45 VTAIL.n11 0.155672
R754 VTAIL.n46 VTAIL.n45 0.155672
R755 VTAIL.n46 VTAIL.n7 0.155672
R756 VTAIL.n53 VTAIL.n7 0.155672
R757 VTAIL.n54 VTAIL.n53 0.155672
R758 VTAIL.n54 VTAIL.n3 0.155672
R759 VTAIL.n61 VTAIL.n3 0.155672
R760 VTAIL.n89 VTAIL.n81 0.155672
R761 VTAIL.n90 VTAIL.n89 0.155672
R762 VTAIL.n90 VTAIL.n77 0.155672
R763 VTAIL.n97 VTAIL.n77 0.155672
R764 VTAIL.n98 VTAIL.n97 0.155672
R765 VTAIL.n98 VTAIL.n73 0.155672
R766 VTAIL.n107 VTAIL.n73 0.155672
R767 VTAIL.n108 VTAIL.n107 0.155672
R768 VTAIL.n108 VTAIL.n69 0.155672
R769 VTAIL.n115 VTAIL.n69 0.155672
R770 VTAIL.n116 VTAIL.n115 0.155672
R771 VTAIL.n116 VTAIL.n65 0.155672
R772 VTAIL.n123 VTAIL.n65 0.155672
R773 VTAIL.n153 VTAIL.n145 0.155672
R774 VTAIL.n154 VTAIL.n153 0.155672
R775 VTAIL.n154 VTAIL.n141 0.155672
R776 VTAIL.n161 VTAIL.n141 0.155672
R777 VTAIL.n162 VTAIL.n161 0.155672
R778 VTAIL.n162 VTAIL.n137 0.155672
R779 VTAIL.n171 VTAIL.n137 0.155672
R780 VTAIL.n172 VTAIL.n171 0.155672
R781 VTAIL.n172 VTAIL.n133 0.155672
R782 VTAIL.n179 VTAIL.n133 0.155672
R783 VTAIL.n180 VTAIL.n179 0.155672
R784 VTAIL.n180 VTAIL.n129 0.155672
R785 VTAIL.n187 VTAIL.n129 0.155672
R786 VTAIL.n439 VTAIL.n381 0.155672
R787 VTAIL.n432 VTAIL.n381 0.155672
R788 VTAIL.n432 VTAIL.n431 0.155672
R789 VTAIL.n431 VTAIL.n385 0.155672
R790 VTAIL.n424 VTAIL.n385 0.155672
R791 VTAIL.n424 VTAIL.n423 0.155672
R792 VTAIL.n423 VTAIL.n389 0.155672
R793 VTAIL.n416 VTAIL.n389 0.155672
R794 VTAIL.n416 VTAIL.n415 0.155672
R795 VTAIL.n415 VTAIL.n395 0.155672
R796 VTAIL.n408 VTAIL.n395 0.155672
R797 VTAIL.n408 VTAIL.n407 0.155672
R798 VTAIL.n407 VTAIL.n399 0.155672
R799 VTAIL.n375 VTAIL.n317 0.155672
R800 VTAIL.n368 VTAIL.n317 0.155672
R801 VTAIL.n368 VTAIL.n367 0.155672
R802 VTAIL.n367 VTAIL.n321 0.155672
R803 VTAIL.n360 VTAIL.n321 0.155672
R804 VTAIL.n360 VTAIL.n359 0.155672
R805 VTAIL.n359 VTAIL.n325 0.155672
R806 VTAIL.n352 VTAIL.n325 0.155672
R807 VTAIL.n352 VTAIL.n351 0.155672
R808 VTAIL.n351 VTAIL.n331 0.155672
R809 VTAIL.n344 VTAIL.n331 0.155672
R810 VTAIL.n344 VTAIL.n343 0.155672
R811 VTAIL.n343 VTAIL.n335 0.155672
R812 VTAIL.n313 VTAIL.n255 0.155672
R813 VTAIL.n306 VTAIL.n255 0.155672
R814 VTAIL.n306 VTAIL.n305 0.155672
R815 VTAIL.n305 VTAIL.n259 0.155672
R816 VTAIL.n298 VTAIL.n259 0.155672
R817 VTAIL.n298 VTAIL.n297 0.155672
R818 VTAIL.n297 VTAIL.n263 0.155672
R819 VTAIL.n290 VTAIL.n263 0.155672
R820 VTAIL.n290 VTAIL.n289 0.155672
R821 VTAIL.n289 VTAIL.n269 0.155672
R822 VTAIL.n282 VTAIL.n269 0.155672
R823 VTAIL.n282 VTAIL.n281 0.155672
R824 VTAIL.n281 VTAIL.n273 0.155672
R825 VTAIL.n249 VTAIL.n191 0.155672
R826 VTAIL.n242 VTAIL.n191 0.155672
R827 VTAIL.n242 VTAIL.n241 0.155672
R828 VTAIL.n241 VTAIL.n195 0.155672
R829 VTAIL.n234 VTAIL.n195 0.155672
R830 VTAIL.n234 VTAIL.n233 0.155672
R831 VTAIL.n233 VTAIL.n199 0.155672
R832 VTAIL.n226 VTAIL.n199 0.155672
R833 VTAIL.n226 VTAIL.n225 0.155672
R834 VTAIL.n225 VTAIL.n205 0.155672
R835 VTAIL.n218 VTAIL.n205 0.155672
R836 VTAIL.n218 VTAIL.n217 0.155672
R837 VTAIL.n217 VTAIL.n209 0.155672
R838 VTAIL VTAIL.n1 0.0586897
R839 B.n521 B.n106 585
R840 B.n106 B.n57 585
R841 B.n523 B.n522 585
R842 B.n525 B.n105 585
R843 B.n528 B.n527 585
R844 B.n529 B.n104 585
R845 B.n531 B.n530 585
R846 B.n533 B.n103 585
R847 B.n536 B.n535 585
R848 B.n537 B.n102 585
R849 B.n539 B.n538 585
R850 B.n541 B.n101 585
R851 B.n544 B.n543 585
R852 B.n545 B.n100 585
R853 B.n547 B.n546 585
R854 B.n549 B.n99 585
R855 B.n552 B.n551 585
R856 B.n553 B.n98 585
R857 B.n555 B.n554 585
R858 B.n557 B.n97 585
R859 B.n560 B.n559 585
R860 B.n561 B.n96 585
R861 B.n563 B.n562 585
R862 B.n565 B.n95 585
R863 B.n568 B.n567 585
R864 B.n569 B.n94 585
R865 B.n571 B.n570 585
R866 B.n573 B.n93 585
R867 B.n576 B.n575 585
R868 B.n577 B.n92 585
R869 B.n579 B.n578 585
R870 B.n581 B.n91 585
R871 B.n584 B.n583 585
R872 B.n585 B.n90 585
R873 B.n587 B.n586 585
R874 B.n589 B.n89 585
R875 B.n592 B.n591 585
R876 B.n593 B.n88 585
R877 B.n595 B.n594 585
R878 B.n597 B.n87 585
R879 B.n600 B.n599 585
R880 B.n602 B.n84 585
R881 B.n604 B.n603 585
R882 B.n606 B.n83 585
R883 B.n609 B.n608 585
R884 B.n610 B.n82 585
R885 B.n612 B.n611 585
R886 B.n614 B.n81 585
R887 B.n617 B.n616 585
R888 B.n618 B.n78 585
R889 B.n621 B.n620 585
R890 B.n623 B.n77 585
R891 B.n626 B.n625 585
R892 B.n627 B.n76 585
R893 B.n629 B.n628 585
R894 B.n631 B.n75 585
R895 B.n634 B.n633 585
R896 B.n635 B.n74 585
R897 B.n637 B.n636 585
R898 B.n639 B.n73 585
R899 B.n642 B.n641 585
R900 B.n643 B.n72 585
R901 B.n645 B.n644 585
R902 B.n647 B.n71 585
R903 B.n650 B.n649 585
R904 B.n651 B.n70 585
R905 B.n653 B.n652 585
R906 B.n655 B.n69 585
R907 B.n658 B.n657 585
R908 B.n659 B.n68 585
R909 B.n661 B.n660 585
R910 B.n663 B.n67 585
R911 B.n666 B.n665 585
R912 B.n667 B.n66 585
R913 B.n669 B.n668 585
R914 B.n671 B.n65 585
R915 B.n674 B.n673 585
R916 B.n675 B.n64 585
R917 B.n677 B.n676 585
R918 B.n679 B.n63 585
R919 B.n682 B.n681 585
R920 B.n683 B.n62 585
R921 B.n685 B.n684 585
R922 B.n687 B.n61 585
R923 B.n690 B.n689 585
R924 B.n691 B.n60 585
R925 B.n693 B.n692 585
R926 B.n695 B.n59 585
R927 B.n698 B.n697 585
R928 B.n699 B.n58 585
R929 B.n520 B.n56 585
R930 B.n702 B.n56 585
R931 B.n519 B.n55 585
R932 B.n703 B.n55 585
R933 B.n518 B.n54 585
R934 B.n704 B.n54 585
R935 B.n517 B.n516 585
R936 B.n516 B.n50 585
R937 B.n515 B.n49 585
R938 B.n710 B.n49 585
R939 B.n514 B.n48 585
R940 B.n711 B.n48 585
R941 B.n513 B.n47 585
R942 B.n712 B.n47 585
R943 B.n512 B.n511 585
R944 B.n511 B.n43 585
R945 B.n510 B.n42 585
R946 B.n718 B.n42 585
R947 B.n509 B.n41 585
R948 B.n719 B.n41 585
R949 B.n508 B.n40 585
R950 B.n720 B.n40 585
R951 B.n507 B.n506 585
R952 B.n506 B.n36 585
R953 B.n505 B.n35 585
R954 B.n726 B.n35 585
R955 B.n504 B.n34 585
R956 B.n727 B.n34 585
R957 B.n503 B.n33 585
R958 B.n728 B.n33 585
R959 B.n502 B.n501 585
R960 B.n501 B.n29 585
R961 B.n500 B.n28 585
R962 B.n734 B.n28 585
R963 B.n499 B.n27 585
R964 B.n735 B.n27 585
R965 B.n498 B.n26 585
R966 B.n736 B.n26 585
R967 B.n497 B.n496 585
R968 B.n496 B.n22 585
R969 B.n495 B.n21 585
R970 B.n742 B.n21 585
R971 B.n494 B.n20 585
R972 B.n743 B.n20 585
R973 B.n493 B.n19 585
R974 B.n744 B.n19 585
R975 B.n492 B.n491 585
R976 B.n491 B.n15 585
R977 B.n490 B.n14 585
R978 B.n750 B.n14 585
R979 B.n489 B.n13 585
R980 B.n751 B.n13 585
R981 B.n488 B.n12 585
R982 B.n752 B.n12 585
R983 B.n487 B.n486 585
R984 B.n486 B.n8 585
R985 B.n485 B.n7 585
R986 B.n758 B.n7 585
R987 B.n484 B.n6 585
R988 B.n759 B.n6 585
R989 B.n483 B.n5 585
R990 B.n760 B.n5 585
R991 B.n482 B.n481 585
R992 B.n481 B.n4 585
R993 B.n480 B.n107 585
R994 B.n480 B.n479 585
R995 B.n470 B.n108 585
R996 B.n109 B.n108 585
R997 B.n472 B.n471 585
R998 B.n473 B.n472 585
R999 B.n469 B.n114 585
R1000 B.n114 B.n113 585
R1001 B.n468 B.n467 585
R1002 B.n467 B.n466 585
R1003 B.n116 B.n115 585
R1004 B.n117 B.n116 585
R1005 B.n459 B.n458 585
R1006 B.n460 B.n459 585
R1007 B.n457 B.n121 585
R1008 B.n125 B.n121 585
R1009 B.n456 B.n455 585
R1010 B.n455 B.n454 585
R1011 B.n123 B.n122 585
R1012 B.n124 B.n123 585
R1013 B.n447 B.n446 585
R1014 B.n448 B.n447 585
R1015 B.n445 B.n129 585
R1016 B.n133 B.n129 585
R1017 B.n444 B.n443 585
R1018 B.n443 B.n442 585
R1019 B.n131 B.n130 585
R1020 B.n132 B.n131 585
R1021 B.n435 B.n434 585
R1022 B.n436 B.n435 585
R1023 B.n433 B.n138 585
R1024 B.n138 B.n137 585
R1025 B.n432 B.n431 585
R1026 B.n431 B.n430 585
R1027 B.n140 B.n139 585
R1028 B.n141 B.n140 585
R1029 B.n423 B.n422 585
R1030 B.n424 B.n423 585
R1031 B.n421 B.n146 585
R1032 B.n146 B.n145 585
R1033 B.n420 B.n419 585
R1034 B.n419 B.n418 585
R1035 B.n148 B.n147 585
R1036 B.n149 B.n148 585
R1037 B.n411 B.n410 585
R1038 B.n412 B.n411 585
R1039 B.n409 B.n153 585
R1040 B.n157 B.n153 585
R1041 B.n408 B.n407 585
R1042 B.n407 B.n406 585
R1043 B.n155 B.n154 585
R1044 B.n156 B.n155 585
R1045 B.n399 B.n398 585
R1046 B.n400 B.n399 585
R1047 B.n397 B.n162 585
R1048 B.n162 B.n161 585
R1049 B.n396 B.n395 585
R1050 B.n395 B.n394 585
R1051 B.n391 B.n166 585
R1052 B.n390 B.n389 585
R1053 B.n387 B.n167 585
R1054 B.n387 B.n165 585
R1055 B.n386 B.n385 585
R1056 B.n384 B.n383 585
R1057 B.n382 B.n169 585
R1058 B.n380 B.n379 585
R1059 B.n378 B.n170 585
R1060 B.n377 B.n376 585
R1061 B.n374 B.n171 585
R1062 B.n372 B.n371 585
R1063 B.n370 B.n172 585
R1064 B.n369 B.n368 585
R1065 B.n366 B.n173 585
R1066 B.n364 B.n363 585
R1067 B.n362 B.n174 585
R1068 B.n361 B.n360 585
R1069 B.n358 B.n175 585
R1070 B.n356 B.n355 585
R1071 B.n354 B.n176 585
R1072 B.n353 B.n352 585
R1073 B.n350 B.n177 585
R1074 B.n348 B.n347 585
R1075 B.n346 B.n178 585
R1076 B.n345 B.n344 585
R1077 B.n342 B.n179 585
R1078 B.n340 B.n339 585
R1079 B.n338 B.n180 585
R1080 B.n337 B.n336 585
R1081 B.n334 B.n181 585
R1082 B.n332 B.n331 585
R1083 B.n330 B.n182 585
R1084 B.n329 B.n328 585
R1085 B.n326 B.n183 585
R1086 B.n324 B.n323 585
R1087 B.n322 B.n184 585
R1088 B.n321 B.n320 585
R1089 B.n318 B.n185 585
R1090 B.n316 B.n315 585
R1091 B.n314 B.n186 585
R1092 B.n312 B.n311 585
R1093 B.n309 B.n189 585
R1094 B.n307 B.n306 585
R1095 B.n305 B.n190 585
R1096 B.n304 B.n303 585
R1097 B.n301 B.n191 585
R1098 B.n299 B.n298 585
R1099 B.n297 B.n192 585
R1100 B.n296 B.n295 585
R1101 B.n293 B.n292 585
R1102 B.n291 B.n290 585
R1103 B.n289 B.n197 585
R1104 B.n287 B.n286 585
R1105 B.n285 B.n198 585
R1106 B.n284 B.n283 585
R1107 B.n281 B.n199 585
R1108 B.n279 B.n278 585
R1109 B.n277 B.n200 585
R1110 B.n276 B.n275 585
R1111 B.n273 B.n201 585
R1112 B.n271 B.n270 585
R1113 B.n269 B.n202 585
R1114 B.n268 B.n267 585
R1115 B.n265 B.n203 585
R1116 B.n263 B.n262 585
R1117 B.n261 B.n204 585
R1118 B.n260 B.n259 585
R1119 B.n257 B.n205 585
R1120 B.n255 B.n254 585
R1121 B.n253 B.n206 585
R1122 B.n252 B.n251 585
R1123 B.n249 B.n207 585
R1124 B.n247 B.n246 585
R1125 B.n245 B.n208 585
R1126 B.n244 B.n243 585
R1127 B.n241 B.n209 585
R1128 B.n239 B.n238 585
R1129 B.n237 B.n210 585
R1130 B.n236 B.n235 585
R1131 B.n233 B.n211 585
R1132 B.n231 B.n230 585
R1133 B.n229 B.n212 585
R1134 B.n228 B.n227 585
R1135 B.n225 B.n213 585
R1136 B.n223 B.n222 585
R1137 B.n221 B.n214 585
R1138 B.n220 B.n219 585
R1139 B.n217 B.n215 585
R1140 B.n164 B.n163 585
R1141 B.n393 B.n392 585
R1142 B.n394 B.n393 585
R1143 B.n160 B.n159 585
R1144 B.n161 B.n160 585
R1145 B.n402 B.n401 585
R1146 B.n401 B.n400 585
R1147 B.n403 B.n158 585
R1148 B.n158 B.n156 585
R1149 B.n405 B.n404 585
R1150 B.n406 B.n405 585
R1151 B.n152 B.n151 585
R1152 B.n157 B.n152 585
R1153 B.n414 B.n413 585
R1154 B.n413 B.n412 585
R1155 B.n415 B.n150 585
R1156 B.n150 B.n149 585
R1157 B.n417 B.n416 585
R1158 B.n418 B.n417 585
R1159 B.n144 B.n143 585
R1160 B.n145 B.n144 585
R1161 B.n426 B.n425 585
R1162 B.n425 B.n424 585
R1163 B.n427 B.n142 585
R1164 B.n142 B.n141 585
R1165 B.n429 B.n428 585
R1166 B.n430 B.n429 585
R1167 B.n136 B.n135 585
R1168 B.n137 B.n136 585
R1169 B.n438 B.n437 585
R1170 B.n437 B.n436 585
R1171 B.n439 B.n134 585
R1172 B.n134 B.n132 585
R1173 B.n441 B.n440 585
R1174 B.n442 B.n441 585
R1175 B.n128 B.n127 585
R1176 B.n133 B.n128 585
R1177 B.n450 B.n449 585
R1178 B.n449 B.n448 585
R1179 B.n451 B.n126 585
R1180 B.n126 B.n124 585
R1181 B.n453 B.n452 585
R1182 B.n454 B.n453 585
R1183 B.n120 B.n119 585
R1184 B.n125 B.n120 585
R1185 B.n462 B.n461 585
R1186 B.n461 B.n460 585
R1187 B.n463 B.n118 585
R1188 B.n118 B.n117 585
R1189 B.n465 B.n464 585
R1190 B.n466 B.n465 585
R1191 B.n112 B.n111 585
R1192 B.n113 B.n112 585
R1193 B.n475 B.n474 585
R1194 B.n474 B.n473 585
R1195 B.n476 B.n110 585
R1196 B.n110 B.n109 585
R1197 B.n478 B.n477 585
R1198 B.n479 B.n478 585
R1199 B.n2 B.n0 585
R1200 B.n4 B.n2 585
R1201 B.n3 B.n1 585
R1202 B.n759 B.n3 585
R1203 B.n757 B.n756 585
R1204 B.n758 B.n757 585
R1205 B.n755 B.n9 585
R1206 B.n9 B.n8 585
R1207 B.n754 B.n753 585
R1208 B.n753 B.n752 585
R1209 B.n11 B.n10 585
R1210 B.n751 B.n11 585
R1211 B.n749 B.n748 585
R1212 B.n750 B.n749 585
R1213 B.n747 B.n16 585
R1214 B.n16 B.n15 585
R1215 B.n746 B.n745 585
R1216 B.n745 B.n744 585
R1217 B.n18 B.n17 585
R1218 B.n743 B.n18 585
R1219 B.n741 B.n740 585
R1220 B.n742 B.n741 585
R1221 B.n739 B.n23 585
R1222 B.n23 B.n22 585
R1223 B.n738 B.n737 585
R1224 B.n737 B.n736 585
R1225 B.n25 B.n24 585
R1226 B.n735 B.n25 585
R1227 B.n733 B.n732 585
R1228 B.n734 B.n733 585
R1229 B.n731 B.n30 585
R1230 B.n30 B.n29 585
R1231 B.n730 B.n729 585
R1232 B.n729 B.n728 585
R1233 B.n32 B.n31 585
R1234 B.n727 B.n32 585
R1235 B.n725 B.n724 585
R1236 B.n726 B.n725 585
R1237 B.n723 B.n37 585
R1238 B.n37 B.n36 585
R1239 B.n722 B.n721 585
R1240 B.n721 B.n720 585
R1241 B.n39 B.n38 585
R1242 B.n719 B.n39 585
R1243 B.n717 B.n716 585
R1244 B.n718 B.n717 585
R1245 B.n715 B.n44 585
R1246 B.n44 B.n43 585
R1247 B.n714 B.n713 585
R1248 B.n713 B.n712 585
R1249 B.n46 B.n45 585
R1250 B.n711 B.n46 585
R1251 B.n709 B.n708 585
R1252 B.n710 B.n709 585
R1253 B.n707 B.n51 585
R1254 B.n51 B.n50 585
R1255 B.n706 B.n705 585
R1256 B.n705 B.n704 585
R1257 B.n53 B.n52 585
R1258 B.n703 B.n53 585
R1259 B.n701 B.n700 585
R1260 B.n702 B.n701 585
R1261 B.n762 B.n761 585
R1262 B.n761 B.n760 585
R1263 B.n393 B.n166 554.963
R1264 B.n701 B.n58 554.963
R1265 B.n395 B.n164 554.963
R1266 B.n106 B.n56 554.963
R1267 B.n193 B.t18 438.985
R1268 B.n187 B.t11 438.985
R1269 B.n79 B.t7 438.985
R1270 B.n85 B.t15 438.985
R1271 B.n193 B.t20 301.132
R1272 B.n85 B.t16 301.132
R1273 B.n187 B.t14 301.132
R1274 B.n79 B.t9 301.132
R1275 B.n194 B.t19 272.041
R1276 B.n86 B.t17 272.041
R1277 B.n188 B.t13 272.041
R1278 B.n80 B.t10 272.041
R1279 B.n524 B.n57 256.663
R1280 B.n526 B.n57 256.663
R1281 B.n532 B.n57 256.663
R1282 B.n534 B.n57 256.663
R1283 B.n540 B.n57 256.663
R1284 B.n542 B.n57 256.663
R1285 B.n548 B.n57 256.663
R1286 B.n550 B.n57 256.663
R1287 B.n556 B.n57 256.663
R1288 B.n558 B.n57 256.663
R1289 B.n564 B.n57 256.663
R1290 B.n566 B.n57 256.663
R1291 B.n572 B.n57 256.663
R1292 B.n574 B.n57 256.663
R1293 B.n580 B.n57 256.663
R1294 B.n582 B.n57 256.663
R1295 B.n588 B.n57 256.663
R1296 B.n590 B.n57 256.663
R1297 B.n596 B.n57 256.663
R1298 B.n598 B.n57 256.663
R1299 B.n605 B.n57 256.663
R1300 B.n607 B.n57 256.663
R1301 B.n613 B.n57 256.663
R1302 B.n615 B.n57 256.663
R1303 B.n622 B.n57 256.663
R1304 B.n624 B.n57 256.663
R1305 B.n630 B.n57 256.663
R1306 B.n632 B.n57 256.663
R1307 B.n638 B.n57 256.663
R1308 B.n640 B.n57 256.663
R1309 B.n646 B.n57 256.663
R1310 B.n648 B.n57 256.663
R1311 B.n654 B.n57 256.663
R1312 B.n656 B.n57 256.663
R1313 B.n662 B.n57 256.663
R1314 B.n664 B.n57 256.663
R1315 B.n670 B.n57 256.663
R1316 B.n672 B.n57 256.663
R1317 B.n678 B.n57 256.663
R1318 B.n680 B.n57 256.663
R1319 B.n686 B.n57 256.663
R1320 B.n688 B.n57 256.663
R1321 B.n694 B.n57 256.663
R1322 B.n696 B.n57 256.663
R1323 B.n388 B.n165 256.663
R1324 B.n168 B.n165 256.663
R1325 B.n381 B.n165 256.663
R1326 B.n375 B.n165 256.663
R1327 B.n373 B.n165 256.663
R1328 B.n367 B.n165 256.663
R1329 B.n365 B.n165 256.663
R1330 B.n359 B.n165 256.663
R1331 B.n357 B.n165 256.663
R1332 B.n351 B.n165 256.663
R1333 B.n349 B.n165 256.663
R1334 B.n343 B.n165 256.663
R1335 B.n341 B.n165 256.663
R1336 B.n335 B.n165 256.663
R1337 B.n333 B.n165 256.663
R1338 B.n327 B.n165 256.663
R1339 B.n325 B.n165 256.663
R1340 B.n319 B.n165 256.663
R1341 B.n317 B.n165 256.663
R1342 B.n310 B.n165 256.663
R1343 B.n308 B.n165 256.663
R1344 B.n302 B.n165 256.663
R1345 B.n300 B.n165 256.663
R1346 B.n294 B.n165 256.663
R1347 B.n196 B.n165 256.663
R1348 B.n288 B.n165 256.663
R1349 B.n282 B.n165 256.663
R1350 B.n280 B.n165 256.663
R1351 B.n274 B.n165 256.663
R1352 B.n272 B.n165 256.663
R1353 B.n266 B.n165 256.663
R1354 B.n264 B.n165 256.663
R1355 B.n258 B.n165 256.663
R1356 B.n256 B.n165 256.663
R1357 B.n250 B.n165 256.663
R1358 B.n248 B.n165 256.663
R1359 B.n242 B.n165 256.663
R1360 B.n240 B.n165 256.663
R1361 B.n234 B.n165 256.663
R1362 B.n232 B.n165 256.663
R1363 B.n226 B.n165 256.663
R1364 B.n224 B.n165 256.663
R1365 B.n218 B.n165 256.663
R1366 B.n216 B.n165 256.663
R1367 B.n393 B.n160 163.367
R1368 B.n401 B.n160 163.367
R1369 B.n401 B.n158 163.367
R1370 B.n405 B.n158 163.367
R1371 B.n405 B.n152 163.367
R1372 B.n413 B.n152 163.367
R1373 B.n413 B.n150 163.367
R1374 B.n417 B.n150 163.367
R1375 B.n417 B.n144 163.367
R1376 B.n425 B.n144 163.367
R1377 B.n425 B.n142 163.367
R1378 B.n429 B.n142 163.367
R1379 B.n429 B.n136 163.367
R1380 B.n437 B.n136 163.367
R1381 B.n437 B.n134 163.367
R1382 B.n441 B.n134 163.367
R1383 B.n441 B.n128 163.367
R1384 B.n449 B.n128 163.367
R1385 B.n449 B.n126 163.367
R1386 B.n453 B.n126 163.367
R1387 B.n453 B.n120 163.367
R1388 B.n461 B.n120 163.367
R1389 B.n461 B.n118 163.367
R1390 B.n465 B.n118 163.367
R1391 B.n465 B.n112 163.367
R1392 B.n474 B.n112 163.367
R1393 B.n474 B.n110 163.367
R1394 B.n478 B.n110 163.367
R1395 B.n478 B.n2 163.367
R1396 B.n761 B.n2 163.367
R1397 B.n761 B.n3 163.367
R1398 B.n757 B.n3 163.367
R1399 B.n757 B.n9 163.367
R1400 B.n753 B.n9 163.367
R1401 B.n753 B.n11 163.367
R1402 B.n749 B.n11 163.367
R1403 B.n749 B.n16 163.367
R1404 B.n745 B.n16 163.367
R1405 B.n745 B.n18 163.367
R1406 B.n741 B.n18 163.367
R1407 B.n741 B.n23 163.367
R1408 B.n737 B.n23 163.367
R1409 B.n737 B.n25 163.367
R1410 B.n733 B.n25 163.367
R1411 B.n733 B.n30 163.367
R1412 B.n729 B.n30 163.367
R1413 B.n729 B.n32 163.367
R1414 B.n725 B.n32 163.367
R1415 B.n725 B.n37 163.367
R1416 B.n721 B.n37 163.367
R1417 B.n721 B.n39 163.367
R1418 B.n717 B.n39 163.367
R1419 B.n717 B.n44 163.367
R1420 B.n713 B.n44 163.367
R1421 B.n713 B.n46 163.367
R1422 B.n709 B.n46 163.367
R1423 B.n709 B.n51 163.367
R1424 B.n705 B.n51 163.367
R1425 B.n705 B.n53 163.367
R1426 B.n701 B.n53 163.367
R1427 B.n389 B.n387 163.367
R1428 B.n387 B.n386 163.367
R1429 B.n383 B.n382 163.367
R1430 B.n380 B.n170 163.367
R1431 B.n376 B.n374 163.367
R1432 B.n372 B.n172 163.367
R1433 B.n368 B.n366 163.367
R1434 B.n364 B.n174 163.367
R1435 B.n360 B.n358 163.367
R1436 B.n356 B.n176 163.367
R1437 B.n352 B.n350 163.367
R1438 B.n348 B.n178 163.367
R1439 B.n344 B.n342 163.367
R1440 B.n340 B.n180 163.367
R1441 B.n336 B.n334 163.367
R1442 B.n332 B.n182 163.367
R1443 B.n328 B.n326 163.367
R1444 B.n324 B.n184 163.367
R1445 B.n320 B.n318 163.367
R1446 B.n316 B.n186 163.367
R1447 B.n311 B.n309 163.367
R1448 B.n307 B.n190 163.367
R1449 B.n303 B.n301 163.367
R1450 B.n299 B.n192 163.367
R1451 B.n295 B.n293 163.367
R1452 B.n290 B.n289 163.367
R1453 B.n287 B.n198 163.367
R1454 B.n283 B.n281 163.367
R1455 B.n279 B.n200 163.367
R1456 B.n275 B.n273 163.367
R1457 B.n271 B.n202 163.367
R1458 B.n267 B.n265 163.367
R1459 B.n263 B.n204 163.367
R1460 B.n259 B.n257 163.367
R1461 B.n255 B.n206 163.367
R1462 B.n251 B.n249 163.367
R1463 B.n247 B.n208 163.367
R1464 B.n243 B.n241 163.367
R1465 B.n239 B.n210 163.367
R1466 B.n235 B.n233 163.367
R1467 B.n231 B.n212 163.367
R1468 B.n227 B.n225 163.367
R1469 B.n223 B.n214 163.367
R1470 B.n219 B.n217 163.367
R1471 B.n395 B.n162 163.367
R1472 B.n399 B.n162 163.367
R1473 B.n399 B.n155 163.367
R1474 B.n407 B.n155 163.367
R1475 B.n407 B.n153 163.367
R1476 B.n411 B.n153 163.367
R1477 B.n411 B.n148 163.367
R1478 B.n419 B.n148 163.367
R1479 B.n419 B.n146 163.367
R1480 B.n423 B.n146 163.367
R1481 B.n423 B.n140 163.367
R1482 B.n431 B.n140 163.367
R1483 B.n431 B.n138 163.367
R1484 B.n435 B.n138 163.367
R1485 B.n435 B.n131 163.367
R1486 B.n443 B.n131 163.367
R1487 B.n443 B.n129 163.367
R1488 B.n447 B.n129 163.367
R1489 B.n447 B.n123 163.367
R1490 B.n455 B.n123 163.367
R1491 B.n455 B.n121 163.367
R1492 B.n459 B.n121 163.367
R1493 B.n459 B.n116 163.367
R1494 B.n467 B.n116 163.367
R1495 B.n467 B.n114 163.367
R1496 B.n472 B.n114 163.367
R1497 B.n472 B.n108 163.367
R1498 B.n480 B.n108 163.367
R1499 B.n481 B.n480 163.367
R1500 B.n481 B.n5 163.367
R1501 B.n6 B.n5 163.367
R1502 B.n7 B.n6 163.367
R1503 B.n486 B.n7 163.367
R1504 B.n486 B.n12 163.367
R1505 B.n13 B.n12 163.367
R1506 B.n14 B.n13 163.367
R1507 B.n491 B.n14 163.367
R1508 B.n491 B.n19 163.367
R1509 B.n20 B.n19 163.367
R1510 B.n21 B.n20 163.367
R1511 B.n496 B.n21 163.367
R1512 B.n496 B.n26 163.367
R1513 B.n27 B.n26 163.367
R1514 B.n28 B.n27 163.367
R1515 B.n501 B.n28 163.367
R1516 B.n501 B.n33 163.367
R1517 B.n34 B.n33 163.367
R1518 B.n35 B.n34 163.367
R1519 B.n506 B.n35 163.367
R1520 B.n506 B.n40 163.367
R1521 B.n41 B.n40 163.367
R1522 B.n42 B.n41 163.367
R1523 B.n511 B.n42 163.367
R1524 B.n511 B.n47 163.367
R1525 B.n48 B.n47 163.367
R1526 B.n49 B.n48 163.367
R1527 B.n516 B.n49 163.367
R1528 B.n516 B.n54 163.367
R1529 B.n55 B.n54 163.367
R1530 B.n56 B.n55 163.367
R1531 B.n697 B.n695 163.367
R1532 B.n693 B.n60 163.367
R1533 B.n689 B.n687 163.367
R1534 B.n685 B.n62 163.367
R1535 B.n681 B.n679 163.367
R1536 B.n677 B.n64 163.367
R1537 B.n673 B.n671 163.367
R1538 B.n669 B.n66 163.367
R1539 B.n665 B.n663 163.367
R1540 B.n661 B.n68 163.367
R1541 B.n657 B.n655 163.367
R1542 B.n653 B.n70 163.367
R1543 B.n649 B.n647 163.367
R1544 B.n645 B.n72 163.367
R1545 B.n641 B.n639 163.367
R1546 B.n637 B.n74 163.367
R1547 B.n633 B.n631 163.367
R1548 B.n629 B.n76 163.367
R1549 B.n625 B.n623 163.367
R1550 B.n621 B.n78 163.367
R1551 B.n616 B.n614 163.367
R1552 B.n612 B.n82 163.367
R1553 B.n608 B.n606 163.367
R1554 B.n604 B.n84 163.367
R1555 B.n599 B.n597 163.367
R1556 B.n595 B.n88 163.367
R1557 B.n591 B.n589 163.367
R1558 B.n587 B.n90 163.367
R1559 B.n583 B.n581 163.367
R1560 B.n579 B.n92 163.367
R1561 B.n575 B.n573 163.367
R1562 B.n571 B.n94 163.367
R1563 B.n567 B.n565 163.367
R1564 B.n563 B.n96 163.367
R1565 B.n559 B.n557 163.367
R1566 B.n555 B.n98 163.367
R1567 B.n551 B.n549 163.367
R1568 B.n547 B.n100 163.367
R1569 B.n543 B.n541 163.367
R1570 B.n539 B.n102 163.367
R1571 B.n535 B.n533 163.367
R1572 B.n531 B.n104 163.367
R1573 B.n527 B.n525 163.367
R1574 B.n523 B.n106 163.367
R1575 B.n394 B.n165 89.0026
R1576 B.n702 B.n57 89.0026
R1577 B.n388 B.n166 71.676
R1578 B.n386 B.n168 71.676
R1579 B.n382 B.n381 71.676
R1580 B.n375 B.n170 71.676
R1581 B.n374 B.n373 71.676
R1582 B.n367 B.n172 71.676
R1583 B.n366 B.n365 71.676
R1584 B.n359 B.n174 71.676
R1585 B.n358 B.n357 71.676
R1586 B.n351 B.n176 71.676
R1587 B.n350 B.n349 71.676
R1588 B.n343 B.n178 71.676
R1589 B.n342 B.n341 71.676
R1590 B.n335 B.n180 71.676
R1591 B.n334 B.n333 71.676
R1592 B.n327 B.n182 71.676
R1593 B.n326 B.n325 71.676
R1594 B.n319 B.n184 71.676
R1595 B.n318 B.n317 71.676
R1596 B.n310 B.n186 71.676
R1597 B.n309 B.n308 71.676
R1598 B.n302 B.n190 71.676
R1599 B.n301 B.n300 71.676
R1600 B.n294 B.n192 71.676
R1601 B.n293 B.n196 71.676
R1602 B.n289 B.n288 71.676
R1603 B.n282 B.n198 71.676
R1604 B.n281 B.n280 71.676
R1605 B.n274 B.n200 71.676
R1606 B.n273 B.n272 71.676
R1607 B.n266 B.n202 71.676
R1608 B.n265 B.n264 71.676
R1609 B.n258 B.n204 71.676
R1610 B.n257 B.n256 71.676
R1611 B.n250 B.n206 71.676
R1612 B.n249 B.n248 71.676
R1613 B.n242 B.n208 71.676
R1614 B.n241 B.n240 71.676
R1615 B.n234 B.n210 71.676
R1616 B.n233 B.n232 71.676
R1617 B.n226 B.n212 71.676
R1618 B.n225 B.n224 71.676
R1619 B.n218 B.n214 71.676
R1620 B.n217 B.n216 71.676
R1621 B.n696 B.n58 71.676
R1622 B.n695 B.n694 71.676
R1623 B.n688 B.n60 71.676
R1624 B.n687 B.n686 71.676
R1625 B.n680 B.n62 71.676
R1626 B.n679 B.n678 71.676
R1627 B.n672 B.n64 71.676
R1628 B.n671 B.n670 71.676
R1629 B.n664 B.n66 71.676
R1630 B.n663 B.n662 71.676
R1631 B.n656 B.n68 71.676
R1632 B.n655 B.n654 71.676
R1633 B.n648 B.n70 71.676
R1634 B.n647 B.n646 71.676
R1635 B.n640 B.n72 71.676
R1636 B.n639 B.n638 71.676
R1637 B.n632 B.n74 71.676
R1638 B.n631 B.n630 71.676
R1639 B.n624 B.n76 71.676
R1640 B.n623 B.n622 71.676
R1641 B.n615 B.n78 71.676
R1642 B.n614 B.n613 71.676
R1643 B.n607 B.n82 71.676
R1644 B.n606 B.n605 71.676
R1645 B.n598 B.n84 71.676
R1646 B.n597 B.n596 71.676
R1647 B.n590 B.n88 71.676
R1648 B.n589 B.n588 71.676
R1649 B.n582 B.n90 71.676
R1650 B.n581 B.n580 71.676
R1651 B.n574 B.n92 71.676
R1652 B.n573 B.n572 71.676
R1653 B.n566 B.n94 71.676
R1654 B.n565 B.n564 71.676
R1655 B.n558 B.n96 71.676
R1656 B.n557 B.n556 71.676
R1657 B.n550 B.n98 71.676
R1658 B.n549 B.n548 71.676
R1659 B.n542 B.n100 71.676
R1660 B.n541 B.n540 71.676
R1661 B.n534 B.n102 71.676
R1662 B.n533 B.n532 71.676
R1663 B.n526 B.n104 71.676
R1664 B.n525 B.n524 71.676
R1665 B.n524 B.n523 71.676
R1666 B.n527 B.n526 71.676
R1667 B.n532 B.n531 71.676
R1668 B.n535 B.n534 71.676
R1669 B.n540 B.n539 71.676
R1670 B.n543 B.n542 71.676
R1671 B.n548 B.n547 71.676
R1672 B.n551 B.n550 71.676
R1673 B.n556 B.n555 71.676
R1674 B.n559 B.n558 71.676
R1675 B.n564 B.n563 71.676
R1676 B.n567 B.n566 71.676
R1677 B.n572 B.n571 71.676
R1678 B.n575 B.n574 71.676
R1679 B.n580 B.n579 71.676
R1680 B.n583 B.n582 71.676
R1681 B.n588 B.n587 71.676
R1682 B.n591 B.n590 71.676
R1683 B.n596 B.n595 71.676
R1684 B.n599 B.n598 71.676
R1685 B.n605 B.n604 71.676
R1686 B.n608 B.n607 71.676
R1687 B.n613 B.n612 71.676
R1688 B.n616 B.n615 71.676
R1689 B.n622 B.n621 71.676
R1690 B.n625 B.n624 71.676
R1691 B.n630 B.n629 71.676
R1692 B.n633 B.n632 71.676
R1693 B.n638 B.n637 71.676
R1694 B.n641 B.n640 71.676
R1695 B.n646 B.n645 71.676
R1696 B.n649 B.n648 71.676
R1697 B.n654 B.n653 71.676
R1698 B.n657 B.n656 71.676
R1699 B.n662 B.n661 71.676
R1700 B.n665 B.n664 71.676
R1701 B.n670 B.n669 71.676
R1702 B.n673 B.n672 71.676
R1703 B.n678 B.n677 71.676
R1704 B.n681 B.n680 71.676
R1705 B.n686 B.n685 71.676
R1706 B.n689 B.n688 71.676
R1707 B.n694 B.n693 71.676
R1708 B.n697 B.n696 71.676
R1709 B.n389 B.n388 71.676
R1710 B.n383 B.n168 71.676
R1711 B.n381 B.n380 71.676
R1712 B.n376 B.n375 71.676
R1713 B.n373 B.n372 71.676
R1714 B.n368 B.n367 71.676
R1715 B.n365 B.n364 71.676
R1716 B.n360 B.n359 71.676
R1717 B.n357 B.n356 71.676
R1718 B.n352 B.n351 71.676
R1719 B.n349 B.n348 71.676
R1720 B.n344 B.n343 71.676
R1721 B.n341 B.n340 71.676
R1722 B.n336 B.n335 71.676
R1723 B.n333 B.n332 71.676
R1724 B.n328 B.n327 71.676
R1725 B.n325 B.n324 71.676
R1726 B.n320 B.n319 71.676
R1727 B.n317 B.n316 71.676
R1728 B.n311 B.n310 71.676
R1729 B.n308 B.n307 71.676
R1730 B.n303 B.n302 71.676
R1731 B.n300 B.n299 71.676
R1732 B.n295 B.n294 71.676
R1733 B.n290 B.n196 71.676
R1734 B.n288 B.n287 71.676
R1735 B.n283 B.n282 71.676
R1736 B.n280 B.n279 71.676
R1737 B.n275 B.n274 71.676
R1738 B.n272 B.n271 71.676
R1739 B.n267 B.n266 71.676
R1740 B.n264 B.n263 71.676
R1741 B.n259 B.n258 71.676
R1742 B.n256 B.n255 71.676
R1743 B.n251 B.n250 71.676
R1744 B.n248 B.n247 71.676
R1745 B.n243 B.n242 71.676
R1746 B.n240 B.n239 71.676
R1747 B.n235 B.n234 71.676
R1748 B.n232 B.n231 71.676
R1749 B.n227 B.n226 71.676
R1750 B.n224 B.n223 71.676
R1751 B.n219 B.n218 71.676
R1752 B.n216 B.n164 71.676
R1753 B.n195 B.n194 59.5399
R1754 B.n313 B.n188 59.5399
R1755 B.n619 B.n80 59.5399
R1756 B.n601 B.n86 59.5399
R1757 B.n394 B.n161 44.8312
R1758 B.n400 B.n161 44.8312
R1759 B.n400 B.n156 44.8312
R1760 B.n406 B.n156 44.8312
R1761 B.n406 B.n157 44.8312
R1762 B.n412 B.n149 44.8312
R1763 B.n418 B.n149 44.8312
R1764 B.n418 B.n145 44.8312
R1765 B.n424 B.n145 44.8312
R1766 B.n424 B.n141 44.8312
R1767 B.n430 B.n141 44.8312
R1768 B.n436 B.n137 44.8312
R1769 B.n436 B.n132 44.8312
R1770 B.n442 B.n132 44.8312
R1771 B.n442 B.n133 44.8312
R1772 B.n448 B.n124 44.8312
R1773 B.n454 B.n124 44.8312
R1774 B.n454 B.n125 44.8312
R1775 B.n460 B.n117 44.8312
R1776 B.n466 B.n117 44.8312
R1777 B.n466 B.n113 44.8312
R1778 B.n473 B.n113 44.8312
R1779 B.n479 B.n109 44.8312
R1780 B.n479 B.n4 44.8312
R1781 B.n760 B.n4 44.8312
R1782 B.n760 B.n759 44.8312
R1783 B.n759 B.n758 44.8312
R1784 B.n758 B.n8 44.8312
R1785 B.n752 B.n751 44.8312
R1786 B.n751 B.n750 44.8312
R1787 B.n750 B.n15 44.8312
R1788 B.n744 B.n15 44.8312
R1789 B.n743 B.n742 44.8312
R1790 B.n742 B.n22 44.8312
R1791 B.n736 B.n22 44.8312
R1792 B.n735 B.n734 44.8312
R1793 B.n734 B.n29 44.8312
R1794 B.n728 B.n29 44.8312
R1795 B.n728 B.n727 44.8312
R1796 B.n726 B.n36 44.8312
R1797 B.n720 B.n36 44.8312
R1798 B.n720 B.n719 44.8312
R1799 B.n719 B.n718 44.8312
R1800 B.n718 B.n43 44.8312
R1801 B.n712 B.n43 44.8312
R1802 B.n711 B.n710 44.8312
R1803 B.n710 B.n50 44.8312
R1804 B.n704 B.n50 44.8312
R1805 B.n704 B.n703 44.8312
R1806 B.n703 B.n702 44.8312
R1807 B.n430 B.t5 42.8534
R1808 B.t3 B.n726 42.8534
R1809 B.t6 B.n109 36.2606
R1810 B.t21 B.n8 36.2606
R1811 B.n700 B.n699 36.059
R1812 B.n521 B.n520 36.059
R1813 B.n396 B.n163 36.059
R1814 B.n392 B.n391 36.059
R1815 B.n125 B.t0 34.9421
R1816 B.t4 B.n743 34.9421
R1817 B.n412 B.t12 29.6679
R1818 B.n712 B.t8 29.6679
R1819 B.n194 B.n193 29.0914
R1820 B.n188 B.n187 29.0914
R1821 B.n80 B.n79 29.0914
R1822 B.n86 B.n85 29.0914
R1823 B.n448 B.t2 28.3493
R1824 B.n736 B.t1 28.3493
R1825 B B.n762 18.0485
R1826 B.n133 B.t2 16.4824
R1827 B.t1 B.n735 16.4824
R1828 B.n157 B.t12 15.1638
R1829 B.t8 B.n711 15.1638
R1830 B.n699 B.n698 10.6151
R1831 B.n698 B.n59 10.6151
R1832 B.n692 B.n59 10.6151
R1833 B.n692 B.n691 10.6151
R1834 B.n691 B.n690 10.6151
R1835 B.n690 B.n61 10.6151
R1836 B.n684 B.n61 10.6151
R1837 B.n684 B.n683 10.6151
R1838 B.n683 B.n682 10.6151
R1839 B.n682 B.n63 10.6151
R1840 B.n676 B.n63 10.6151
R1841 B.n676 B.n675 10.6151
R1842 B.n675 B.n674 10.6151
R1843 B.n674 B.n65 10.6151
R1844 B.n668 B.n65 10.6151
R1845 B.n668 B.n667 10.6151
R1846 B.n667 B.n666 10.6151
R1847 B.n666 B.n67 10.6151
R1848 B.n660 B.n67 10.6151
R1849 B.n660 B.n659 10.6151
R1850 B.n659 B.n658 10.6151
R1851 B.n658 B.n69 10.6151
R1852 B.n652 B.n69 10.6151
R1853 B.n652 B.n651 10.6151
R1854 B.n651 B.n650 10.6151
R1855 B.n650 B.n71 10.6151
R1856 B.n644 B.n71 10.6151
R1857 B.n644 B.n643 10.6151
R1858 B.n643 B.n642 10.6151
R1859 B.n642 B.n73 10.6151
R1860 B.n636 B.n73 10.6151
R1861 B.n636 B.n635 10.6151
R1862 B.n635 B.n634 10.6151
R1863 B.n634 B.n75 10.6151
R1864 B.n628 B.n75 10.6151
R1865 B.n628 B.n627 10.6151
R1866 B.n627 B.n626 10.6151
R1867 B.n626 B.n77 10.6151
R1868 B.n620 B.n77 10.6151
R1869 B.n618 B.n617 10.6151
R1870 B.n617 B.n81 10.6151
R1871 B.n611 B.n81 10.6151
R1872 B.n611 B.n610 10.6151
R1873 B.n610 B.n609 10.6151
R1874 B.n609 B.n83 10.6151
R1875 B.n603 B.n83 10.6151
R1876 B.n603 B.n602 10.6151
R1877 B.n600 B.n87 10.6151
R1878 B.n594 B.n87 10.6151
R1879 B.n594 B.n593 10.6151
R1880 B.n593 B.n592 10.6151
R1881 B.n592 B.n89 10.6151
R1882 B.n586 B.n89 10.6151
R1883 B.n586 B.n585 10.6151
R1884 B.n585 B.n584 10.6151
R1885 B.n584 B.n91 10.6151
R1886 B.n578 B.n91 10.6151
R1887 B.n578 B.n577 10.6151
R1888 B.n577 B.n576 10.6151
R1889 B.n576 B.n93 10.6151
R1890 B.n570 B.n93 10.6151
R1891 B.n570 B.n569 10.6151
R1892 B.n569 B.n568 10.6151
R1893 B.n568 B.n95 10.6151
R1894 B.n562 B.n95 10.6151
R1895 B.n562 B.n561 10.6151
R1896 B.n561 B.n560 10.6151
R1897 B.n560 B.n97 10.6151
R1898 B.n554 B.n97 10.6151
R1899 B.n554 B.n553 10.6151
R1900 B.n553 B.n552 10.6151
R1901 B.n552 B.n99 10.6151
R1902 B.n546 B.n99 10.6151
R1903 B.n546 B.n545 10.6151
R1904 B.n545 B.n544 10.6151
R1905 B.n544 B.n101 10.6151
R1906 B.n538 B.n101 10.6151
R1907 B.n538 B.n537 10.6151
R1908 B.n537 B.n536 10.6151
R1909 B.n536 B.n103 10.6151
R1910 B.n530 B.n103 10.6151
R1911 B.n530 B.n529 10.6151
R1912 B.n529 B.n528 10.6151
R1913 B.n528 B.n105 10.6151
R1914 B.n522 B.n105 10.6151
R1915 B.n522 B.n521 10.6151
R1916 B.n397 B.n396 10.6151
R1917 B.n398 B.n397 10.6151
R1918 B.n398 B.n154 10.6151
R1919 B.n408 B.n154 10.6151
R1920 B.n409 B.n408 10.6151
R1921 B.n410 B.n409 10.6151
R1922 B.n410 B.n147 10.6151
R1923 B.n420 B.n147 10.6151
R1924 B.n421 B.n420 10.6151
R1925 B.n422 B.n421 10.6151
R1926 B.n422 B.n139 10.6151
R1927 B.n432 B.n139 10.6151
R1928 B.n433 B.n432 10.6151
R1929 B.n434 B.n433 10.6151
R1930 B.n434 B.n130 10.6151
R1931 B.n444 B.n130 10.6151
R1932 B.n445 B.n444 10.6151
R1933 B.n446 B.n445 10.6151
R1934 B.n446 B.n122 10.6151
R1935 B.n456 B.n122 10.6151
R1936 B.n457 B.n456 10.6151
R1937 B.n458 B.n457 10.6151
R1938 B.n458 B.n115 10.6151
R1939 B.n468 B.n115 10.6151
R1940 B.n469 B.n468 10.6151
R1941 B.n471 B.n469 10.6151
R1942 B.n471 B.n470 10.6151
R1943 B.n470 B.n107 10.6151
R1944 B.n482 B.n107 10.6151
R1945 B.n483 B.n482 10.6151
R1946 B.n484 B.n483 10.6151
R1947 B.n485 B.n484 10.6151
R1948 B.n487 B.n485 10.6151
R1949 B.n488 B.n487 10.6151
R1950 B.n489 B.n488 10.6151
R1951 B.n490 B.n489 10.6151
R1952 B.n492 B.n490 10.6151
R1953 B.n493 B.n492 10.6151
R1954 B.n494 B.n493 10.6151
R1955 B.n495 B.n494 10.6151
R1956 B.n497 B.n495 10.6151
R1957 B.n498 B.n497 10.6151
R1958 B.n499 B.n498 10.6151
R1959 B.n500 B.n499 10.6151
R1960 B.n502 B.n500 10.6151
R1961 B.n503 B.n502 10.6151
R1962 B.n504 B.n503 10.6151
R1963 B.n505 B.n504 10.6151
R1964 B.n507 B.n505 10.6151
R1965 B.n508 B.n507 10.6151
R1966 B.n509 B.n508 10.6151
R1967 B.n510 B.n509 10.6151
R1968 B.n512 B.n510 10.6151
R1969 B.n513 B.n512 10.6151
R1970 B.n514 B.n513 10.6151
R1971 B.n515 B.n514 10.6151
R1972 B.n517 B.n515 10.6151
R1973 B.n518 B.n517 10.6151
R1974 B.n519 B.n518 10.6151
R1975 B.n520 B.n519 10.6151
R1976 B.n391 B.n390 10.6151
R1977 B.n390 B.n167 10.6151
R1978 B.n385 B.n167 10.6151
R1979 B.n385 B.n384 10.6151
R1980 B.n384 B.n169 10.6151
R1981 B.n379 B.n169 10.6151
R1982 B.n379 B.n378 10.6151
R1983 B.n378 B.n377 10.6151
R1984 B.n377 B.n171 10.6151
R1985 B.n371 B.n171 10.6151
R1986 B.n371 B.n370 10.6151
R1987 B.n370 B.n369 10.6151
R1988 B.n369 B.n173 10.6151
R1989 B.n363 B.n173 10.6151
R1990 B.n363 B.n362 10.6151
R1991 B.n362 B.n361 10.6151
R1992 B.n361 B.n175 10.6151
R1993 B.n355 B.n175 10.6151
R1994 B.n355 B.n354 10.6151
R1995 B.n354 B.n353 10.6151
R1996 B.n353 B.n177 10.6151
R1997 B.n347 B.n177 10.6151
R1998 B.n347 B.n346 10.6151
R1999 B.n346 B.n345 10.6151
R2000 B.n345 B.n179 10.6151
R2001 B.n339 B.n179 10.6151
R2002 B.n339 B.n338 10.6151
R2003 B.n338 B.n337 10.6151
R2004 B.n337 B.n181 10.6151
R2005 B.n331 B.n181 10.6151
R2006 B.n331 B.n330 10.6151
R2007 B.n330 B.n329 10.6151
R2008 B.n329 B.n183 10.6151
R2009 B.n323 B.n183 10.6151
R2010 B.n323 B.n322 10.6151
R2011 B.n322 B.n321 10.6151
R2012 B.n321 B.n185 10.6151
R2013 B.n315 B.n185 10.6151
R2014 B.n315 B.n314 10.6151
R2015 B.n312 B.n189 10.6151
R2016 B.n306 B.n189 10.6151
R2017 B.n306 B.n305 10.6151
R2018 B.n305 B.n304 10.6151
R2019 B.n304 B.n191 10.6151
R2020 B.n298 B.n191 10.6151
R2021 B.n298 B.n297 10.6151
R2022 B.n297 B.n296 10.6151
R2023 B.n292 B.n291 10.6151
R2024 B.n291 B.n197 10.6151
R2025 B.n286 B.n197 10.6151
R2026 B.n286 B.n285 10.6151
R2027 B.n285 B.n284 10.6151
R2028 B.n284 B.n199 10.6151
R2029 B.n278 B.n199 10.6151
R2030 B.n278 B.n277 10.6151
R2031 B.n277 B.n276 10.6151
R2032 B.n276 B.n201 10.6151
R2033 B.n270 B.n201 10.6151
R2034 B.n270 B.n269 10.6151
R2035 B.n269 B.n268 10.6151
R2036 B.n268 B.n203 10.6151
R2037 B.n262 B.n203 10.6151
R2038 B.n262 B.n261 10.6151
R2039 B.n261 B.n260 10.6151
R2040 B.n260 B.n205 10.6151
R2041 B.n254 B.n205 10.6151
R2042 B.n254 B.n253 10.6151
R2043 B.n253 B.n252 10.6151
R2044 B.n252 B.n207 10.6151
R2045 B.n246 B.n207 10.6151
R2046 B.n246 B.n245 10.6151
R2047 B.n245 B.n244 10.6151
R2048 B.n244 B.n209 10.6151
R2049 B.n238 B.n209 10.6151
R2050 B.n238 B.n237 10.6151
R2051 B.n237 B.n236 10.6151
R2052 B.n236 B.n211 10.6151
R2053 B.n230 B.n211 10.6151
R2054 B.n230 B.n229 10.6151
R2055 B.n229 B.n228 10.6151
R2056 B.n228 B.n213 10.6151
R2057 B.n222 B.n213 10.6151
R2058 B.n222 B.n221 10.6151
R2059 B.n221 B.n220 10.6151
R2060 B.n220 B.n215 10.6151
R2061 B.n215 B.n163 10.6151
R2062 B.n392 B.n159 10.6151
R2063 B.n402 B.n159 10.6151
R2064 B.n403 B.n402 10.6151
R2065 B.n404 B.n403 10.6151
R2066 B.n404 B.n151 10.6151
R2067 B.n414 B.n151 10.6151
R2068 B.n415 B.n414 10.6151
R2069 B.n416 B.n415 10.6151
R2070 B.n416 B.n143 10.6151
R2071 B.n426 B.n143 10.6151
R2072 B.n427 B.n426 10.6151
R2073 B.n428 B.n427 10.6151
R2074 B.n428 B.n135 10.6151
R2075 B.n438 B.n135 10.6151
R2076 B.n439 B.n438 10.6151
R2077 B.n440 B.n439 10.6151
R2078 B.n440 B.n127 10.6151
R2079 B.n450 B.n127 10.6151
R2080 B.n451 B.n450 10.6151
R2081 B.n452 B.n451 10.6151
R2082 B.n452 B.n119 10.6151
R2083 B.n462 B.n119 10.6151
R2084 B.n463 B.n462 10.6151
R2085 B.n464 B.n463 10.6151
R2086 B.n464 B.n111 10.6151
R2087 B.n475 B.n111 10.6151
R2088 B.n476 B.n475 10.6151
R2089 B.n477 B.n476 10.6151
R2090 B.n477 B.n0 10.6151
R2091 B.n756 B.n1 10.6151
R2092 B.n756 B.n755 10.6151
R2093 B.n755 B.n754 10.6151
R2094 B.n754 B.n10 10.6151
R2095 B.n748 B.n10 10.6151
R2096 B.n748 B.n747 10.6151
R2097 B.n747 B.n746 10.6151
R2098 B.n746 B.n17 10.6151
R2099 B.n740 B.n17 10.6151
R2100 B.n740 B.n739 10.6151
R2101 B.n739 B.n738 10.6151
R2102 B.n738 B.n24 10.6151
R2103 B.n732 B.n24 10.6151
R2104 B.n732 B.n731 10.6151
R2105 B.n731 B.n730 10.6151
R2106 B.n730 B.n31 10.6151
R2107 B.n724 B.n31 10.6151
R2108 B.n724 B.n723 10.6151
R2109 B.n723 B.n722 10.6151
R2110 B.n722 B.n38 10.6151
R2111 B.n716 B.n38 10.6151
R2112 B.n716 B.n715 10.6151
R2113 B.n715 B.n714 10.6151
R2114 B.n714 B.n45 10.6151
R2115 B.n708 B.n45 10.6151
R2116 B.n708 B.n707 10.6151
R2117 B.n707 B.n706 10.6151
R2118 B.n706 B.n52 10.6151
R2119 B.n700 B.n52 10.6151
R2120 B.n460 B.t0 9.88962
R2121 B.n744 B.t4 9.88962
R2122 B.n473 B.t6 8.57107
R2123 B.n752 B.t21 8.57107
R2124 B.n619 B.n618 6.5566
R2125 B.n602 B.n601 6.5566
R2126 B.n313 B.n312 6.5566
R2127 B.n296 B.n195 6.5566
R2128 B.n620 B.n619 4.05904
R2129 B.n601 B.n600 4.05904
R2130 B.n314 B.n313 4.05904
R2131 B.n292 B.n195 4.05904
R2132 B.n762 B.n0 2.81026
R2133 B.n762 B.n1 2.81026
R2134 B.t5 B.n137 1.97832
R2135 B.n727 B.t3 1.97832
R2136 VP.n10 VP.t5 265.137
R2137 VP.n5 VP.t4 235.028
R2138 VP.n3 VP.t6 235.028
R2139 VP.n32 VP.t2 235.028
R2140 VP.n39 VP.t3 235.028
R2141 VP.n21 VP.t1 235.028
R2142 VP.n14 VP.t0 235.028
R2143 VP.n9 VP.t7 235.028
R2144 VP.n23 VP.n5 173.534
R2145 VP.n40 VP.n39 173.534
R2146 VP.n22 VP.n21 173.534
R2147 VP.n12 VP.n11 161.3
R2148 VP.n13 VP.n8 161.3
R2149 VP.n16 VP.n15 161.3
R2150 VP.n17 VP.n7 161.3
R2151 VP.n19 VP.n18 161.3
R2152 VP.n20 VP.n6 161.3
R2153 VP.n38 VP.n0 161.3
R2154 VP.n37 VP.n36 161.3
R2155 VP.n35 VP.n1 161.3
R2156 VP.n34 VP.n33 161.3
R2157 VP.n31 VP.n2 161.3
R2158 VP.n30 VP.n29 161.3
R2159 VP.n28 VP.n27 161.3
R2160 VP.n26 VP.n4 161.3
R2161 VP.n25 VP.n24 161.3
R2162 VP.n10 VP.n9 51.4127
R2163 VP.n23 VP.n22 43.6369
R2164 VP.n26 VP.n25 40.4934
R2165 VP.n27 VP.n26 40.4934
R2166 VP.n31 VP.n30 40.4934
R2167 VP.n33 VP.n31 40.4934
R2168 VP.n37 VP.n1 40.4934
R2169 VP.n38 VP.n37 40.4934
R2170 VP.n20 VP.n19 40.4934
R2171 VP.n19 VP.n7 40.4934
R2172 VP.n15 VP.n13 40.4934
R2173 VP.n13 VP.n12 40.4934
R2174 VP.n11 VP.n10 27.0291
R2175 VP.n25 VP.n5 12.234
R2176 VP.n27 VP.n3 12.234
R2177 VP.n30 VP.n3 12.234
R2178 VP.n33 VP.n32 12.234
R2179 VP.n32 VP.n1 12.234
R2180 VP.n39 VP.n38 12.234
R2181 VP.n21 VP.n20 12.234
R2182 VP.n15 VP.n14 12.234
R2183 VP.n14 VP.n7 12.234
R2184 VP.n12 VP.n9 12.234
R2185 VP.n11 VP.n8 0.189894
R2186 VP.n16 VP.n8 0.189894
R2187 VP.n17 VP.n16 0.189894
R2188 VP.n18 VP.n17 0.189894
R2189 VP.n18 VP.n6 0.189894
R2190 VP.n22 VP.n6 0.189894
R2191 VP.n24 VP.n23 0.189894
R2192 VP.n24 VP.n4 0.189894
R2193 VP.n28 VP.n4 0.189894
R2194 VP.n29 VP.n28 0.189894
R2195 VP.n29 VP.n2 0.189894
R2196 VP.n34 VP.n2 0.189894
R2197 VP.n35 VP.n34 0.189894
R2198 VP.n36 VP.n35 0.189894
R2199 VP.n36 VP.n0 0.189894
R2200 VP.n40 VP.n0 0.189894
R2201 VP VP.n40 0.0516364
R2202 VDD1 VDD1.n0 62.9886
R2203 VDD1.n3 VDD1.n2 62.8749
R2204 VDD1.n3 VDD1.n1 62.8749
R2205 VDD1.n5 VDD1.n4 62.2837
R2206 VDD1.n5 VDD1.n3 39.9535
R2207 VDD1.n4 VDD1.t7 1.73582
R2208 VDD1.n4 VDD1.t6 1.73582
R2209 VDD1.n0 VDD1.t2 1.73582
R2210 VDD1.n0 VDD1.t0 1.73582
R2211 VDD1.n2 VDD1.t5 1.73582
R2212 VDD1.n2 VDD1.t4 1.73582
R2213 VDD1.n1 VDD1.t3 1.73582
R2214 VDD1.n1 VDD1.t1 1.73582
R2215 VDD1 VDD1.n5 0.588862
C0 VTAIL VN 6.57567f
C1 VN VDD2 6.62615f
C2 VDD1 VP 6.84383f
C3 VDD1 VN 0.148599f
C4 VTAIL VDD2 8.79237f
C5 VP VN 5.80786f
C6 VDD1 VTAIL 8.74754f
C7 VDD1 VDD2 1.05764f
C8 VTAIL VP 6.58977f
C9 VP VDD2 0.36696f
C10 VDD2 B 3.89006f
C11 VDD1 B 4.171769f
C12 VTAIL B 9.028191f
C13 VN B 10.142011f
C14 VP B 8.441841f
C15 VDD1.t2 B 0.229819f
C16 VDD1.t0 B 0.229819f
C17 VDD1.n0 B 2.04586f
C18 VDD1.t3 B 0.229819f
C19 VDD1.t1 B 0.229819f
C20 VDD1.n1 B 2.04508f
C21 VDD1.t5 B 0.229819f
C22 VDD1.t4 B 0.229819f
C23 VDD1.n2 B 2.04508f
C24 VDD1.n3 B 2.5119f
C25 VDD1.t7 B 0.229819f
C26 VDD1.t6 B 0.229819f
C27 VDD1.n4 B 2.04155f
C28 VDD1.n5 B 2.48566f
C29 VP.n0 B 0.035776f
C30 VP.t3 B 1.29935f
C31 VP.n1 B 0.054645f
C32 VP.n2 B 0.035776f
C33 VP.t6 B 1.29935f
C34 VP.n3 B 0.47907f
C35 VP.n4 B 0.035776f
C36 VP.t4 B 1.29935f
C37 VP.n5 B 0.536151f
C38 VP.n6 B 0.035776f
C39 VP.t1 B 1.29935f
C40 VP.n7 B 0.054645f
C41 VP.n8 B 0.035776f
C42 VP.t7 B 1.29935f
C43 VP.n9 B 0.531292f
C44 VP.t5 B 1.36552f
C45 VP.n10 B 0.55774f
C46 VP.n11 B 0.18519f
C47 VP.n12 B 0.054645f
C48 VP.n13 B 0.028921f
C49 VP.t0 B 1.29935f
C50 VP.n14 B 0.47907f
C51 VP.n15 B 0.054645f
C52 VP.n16 B 0.035776f
C53 VP.n17 B 0.035776f
C54 VP.n18 B 0.035776f
C55 VP.n19 B 0.028921f
C56 VP.n20 B 0.054645f
C57 VP.n21 B 0.536151f
C58 VP.n22 B 1.57694f
C59 VP.n23 B 1.60641f
C60 VP.n24 B 0.035776f
C61 VP.n25 B 0.054645f
C62 VP.n26 B 0.028921f
C63 VP.n27 B 0.054645f
C64 VP.n28 B 0.035776f
C65 VP.n29 B 0.035776f
C66 VP.n30 B 0.054645f
C67 VP.n31 B 0.028921f
C68 VP.t2 B 1.29935f
C69 VP.n32 B 0.47907f
C70 VP.n33 B 0.054645f
C71 VP.n34 B 0.035776f
C72 VP.n35 B 0.035776f
C73 VP.n36 B 0.035776f
C74 VP.n37 B 0.028921f
C75 VP.n38 B 0.054645f
C76 VP.n39 B 0.536151f
C77 VP.n40 B 0.032054f
C78 VTAIL.t12 B 0.174851f
C79 VTAIL.t13 B 0.174851f
C80 VTAIL.n0 B 1.49614f
C81 VTAIL.n1 B 0.275012f
C82 VTAIL.n2 B 0.026865f
C83 VTAIL.n3 B 0.019392f
C84 VTAIL.n4 B 0.010421f
C85 VTAIL.n5 B 0.02463f
C86 VTAIL.n6 B 0.011033f
C87 VTAIL.n7 B 0.019392f
C88 VTAIL.n8 B 0.010421f
C89 VTAIL.n9 B 0.02463f
C90 VTAIL.n10 B 0.010727f
C91 VTAIL.n11 B 0.019392f
C92 VTAIL.n12 B 0.011033f
C93 VTAIL.n13 B 0.02463f
C94 VTAIL.n14 B 0.011033f
C95 VTAIL.n15 B 0.019392f
C96 VTAIL.n16 B 0.010421f
C97 VTAIL.n17 B 0.02463f
C98 VTAIL.n18 B 0.011033f
C99 VTAIL.n19 B 0.927415f
C100 VTAIL.n20 B 0.010421f
C101 VTAIL.t10 B 0.041538f
C102 VTAIL.n21 B 0.135424f
C103 VTAIL.n22 B 0.017412f
C104 VTAIL.n23 B 0.018473f
C105 VTAIL.n24 B 0.02463f
C106 VTAIL.n25 B 0.011033f
C107 VTAIL.n26 B 0.010421f
C108 VTAIL.n27 B 0.019392f
C109 VTAIL.n28 B 0.019392f
C110 VTAIL.n29 B 0.010421f
C111 VTAIL.n30 B 0.011033f
C112 VTAIL.n31 B 0.02463f
C113 VTAIL.n32 B 0.02463f
C114 VTAIL.n33 B 0.011033f
C115 VTAIL.n34 B 0.010421f
C116 VTAIL.n35 B 0.019392f
C117 VTAIL.n36 B 0.019392f
C118 VTAIL.n37 B 0.010421f
C119 VTAIL.n38 B 0.010421f
C120 VTAIL.n39 B 0.011033f
C121 VTAIL.n40 B 0.02463f
C122 VTAIL.n41 B 0.02463f
C123 VTAIL.n42 B 0.02463f
C124 VTAIL.n43 B 0.010727f
C125 VTAIL.n44 B 0.010421f
C126 VTAIL.n45 B 0.019392f
C127 VTAIL.n46 B 0.019392f
C128 VTAIL.n47 B 0.010421f
C129 VTAIL.n48 B 0.011033f
C130 VTAIL.n49 B 0.02463f
C131 VTAIL.n50 B 0.02463f
C132 VTAIL.n51 B 0.011033f
C133 VTAIL.n52 B 0.010421f
C134 VTAIL.n53 B 0.019392f
C135 VTAIL.n54 B 0.019392f
C136 VTAIL.n55 B 0.010421f
C137 VTAIL.n56 B 0.011033f
C138 VTAIL.n57 B 0.02463f
C139 VTAIL.n58 B 0.052626f
C140 VTAIL.n59 B 0.011033f
C141 VTAIL.n60 B 0.010421f
C142 VTAIL.n61 B 0.045089f
C143 VTAIL.n62 B 0.029383f
C144 VTAIL.n63 B 0.126871f
C145 VTAIL.n64 B 0.026865f
C146 VTAIL.n65 B 0.019392f
C147 VTAIL.n66 B 0.010421f
C148 VTAIL.n67 B 0.02463f
C149 VTAIL.n68 B 0.011033f
C150 VTAIL.n69 B 0.019392f
C151 VTAIL.n70 B 0.010421f
C152 VTAIL.n71 B 0.02463f
C153 VTAIL.n72 B 0.010727f
C154 VTAIL.n73 B 0.019392f
C155 VTAIL.n74 B 0.011033f
C156 VTAIL.n75 B 0.02463f
C157 VTAIL.n76 B 0.011033f
C158 VTAIL.n77 B 0.019392f
C159 VTAIL.n78 B 0.010421f
C160 VTAIL.n79 B 0.02463f
C161 VTAIL.n80 B 0.011033f
C162 VTAIL.n81 B 0.927415f
C163 VTAIL.n82 B 0.010421f
C164 VTAIL.t6 B 0.041538f
C165 VTAIL.n83 B 0.135424f
C166 VTAIL.n84 B 0.017412f
C167 VTAIL.n85 B 0.018473f
C168 VTAIL.n86 B 0.02463f
C169 VTAIL.n87 B 0.011033f
C170 VTAIL.n88 B 0.010421f
C171 VTAIL.n89 B 0.019392f
C172 VTAIL.n90 B 0.019392f
C173 VTAIL.n91 B 0.010421f
C174 VTAIL.n92 B 0.011033f
C175 VTAIL.n93 B 0.02463f
C176 VTAIL.n94 B 0.02463f
C177 VTAIL.n95 B 0.011033f
C178 VTAIL.n96 B 0.010421f
C179 VTAIL.n97 B 0.019392f
C180 VTAIL.n98 B 0.019392f
C181 VTAIL.n99 B 0.010421f
C182 VTAIL.n100 B 0.010421f
C183 VTAIL.n101 B 0.011033f
C184 VTAIL.n102 B 0.02463f
C185 VTAIL.n103 B 0.02463f
C186 VTAIL.n104 B 0.02463f
C187 VTAIL.n105 B 0.010727f
C188 VTAIL.n106 B 0.010421f
C189 VTAIL.n107 B 0.019392f
C190 VTAIL.n108 B 0.019392f
C191 VTAIL.n109 B 0.010421f
C192 VTAIL.n110 B 0.011033f
C193 VTAIL.n111 B 0.02463f
C194 VTAIL.n112 B 0.02463f
C195 VTAIL.n113 B 0.011033f
C196 VTAIL.n114 B 0.010421f
C197 VTAIL.n115 B 0.019392f
C198 VTAIL.n116 B 0.019392f
C199 VTAIL.n117 B 0.010421f
C200 VTAIL.n118 B 0.011033f
C201 VTAIL.n119 B 0.02463f
C202 VTAIL.n120 B 0.052626f
C203 VTAIL.n121 B 0.011033f
C204 VTAIL.n122 B 0.010421f
C205 VTAIL.n123 B 0.045089f
C206 VTAIL.n124 B 0.029383f
C207 VTAIL.n125 B 0.126871f
C208 VTAIL.t2 B 0.174851f
C209 VTAIL.t0 B 0.174851f
C210 VTAIL.n126 B 1.49614f
C211 VTAIL.n127 B 0.352177f
C212 VTAIL.n128 B 0.026865f
C213 VTAIL.n129 B 0.019392f
C214 VTAIL.n130 B 0.010421f
C215 VTAIL.n131 B 0.02463f
C216 VTAIL.n132 B 0.011033f
C217 VTAIL.n133 B 0.019392f
C218 VTAIL.n134 B 0.010421f
C219 VTAIL.n135 B 0.02463f
C220 VTAIL.n136 B 0.010727f
C221 VTAIL.n137 B 0.019392f
C222 VTAIL.n138 B 0.011033f
C223 VTAIL.n139 B 0.02463f
C224 VTAIL.n140 B 0.011033f
C225 VTAIL.n141 B 0.019392f
C226 VTAIL.n142 B 0.010421f
C227 VTAIL.n143 B 0.02463f
C228 VTAIL.n144 B 0.011033f
C229 VTAIL.n145 B 0.927415f
C230 VTAIL.n146 B 0.010421f
C231 VTAIL.t5 B 0.041538f
C232 VTAIL.n147 B 0.135424f
C233 VTAIL.n148 B 0.017412f
C234 VTAIL.n149 B 0.018473f
C235 VTAIL.n150 B 0.02463f
C236 VTAIL.n151 B 0.011033f
C237 VTAIL.n152 B 0.010421f
C238 VTAIL.n153 B 0.019392f
C239 VTAIL.n154 B 0.019392f
C240 VTAIL.n155 B 0.010421f
C241 VTAIL.n156 B 0.011033f
C242 VTAIL.n157 B 0.02463f
C243 VTAIL.n158 B 0.02463f
C244 VTAIL.n159 B 0.011033f
C245 VTAIL.n160 B 0.010421f
C246 VTAIL.n161 B 0.019392f
C247 VTAIL.n162 B 0.019392f
C248 VTAIL.n163 B 0.010421f
C249 VTAIL.n164 B 0.010421f
C250 VTAIL.n165 B 0.011033f
C251 VTAIL.n166 B 0.02463f
C252 VTAIL.n167 B 0.02463f
C253 VTAIL.n168 B 0.02463f
C254 VTAIL.n169 B 0.010727f
C255 VTAIL.n170 B 0.010421f
C256 VTAIL.n171 B 0.019392f
C257 VTAIL.n172 B 0.019392f
C258 VTAIL.n173 B 0.010421f
C259 VTAIL.n174 B 0.011033f
C260 VTAIL.n175 B 0.02463f
C261 VTAIL.n176 B 0.02463f
C262 VTAIL.n177 B 0.011033f
C263 VTAIL.n178 B 0.010421f
C264 VTAIL.n179 B 0.019392f
C265 VTAIL.n180 B 0.019392f
C266 VTAIL.n181 B 0.010421f
C267 VTAIL.n182 B 0.011033f
C268 VTAIL.n183 B 0.02463f
C269 VTAIL.n184 B 0.052626f
C270 VTAIL.n185 B 0.011033f
C271 VTAIL.n186 B 0.010421f
C272 VTAIL.n187 B 0.045089f
C273 VTAIL.n188 B 0.029383f
C274 VTAIL.n189 B 1.05636f
C275 VTAIL.n190 B 0.026865f
C276 VTAIL.n191 B 0.019392f
C277 VTAIL.n192 B 0.010421f
C278 VTAIL.n193 B 0.02463f
C279 VTAIL.n194 B 0.011033f
C280 VTAIL.n195 B 0.019392f
C281 VTAIL.n196 B 0.010421f
C282 VTAIL.n197 B 0.02463f
C283 VTAIL.n198 B 0.010727f
C284 VTAIL.n199 B 0.019392f
C285 VTAIL.n200 B 0.010727f
C286 VTAIL.n201 B 0.010421f
C287 VTAIL.n202 B 0.02463f
C288 VTAIL.n203 B 0.02463f
C289 VTAIL.n204 B 0.011033f
C290 VTAIL.n205 B 0.019392f
C291 VTAIL.n206 B 0.010421f
C292 VTAIL.n207 B 0.02463f
C293 VTAIL.n208 B 0.011033f
C294 VTAIL.n209 B 0.927415f
C295 VTAIL.n210 B 0.010421f
C296 VTAIL.t14 B 0.041538f
C297 VTAIL.n211 B 0.135424f
C298 VTAIL.n212 B 0.017412f
C299 VTAIL.n213 B 0.018473f
C300 VTAIL.n214 B 0.02463f
C301 VTAIL.n215 B 0.011033f
C302 VTAIL.n216 B 0.010421f
C303 VTAIL.n217 B 0.019392f
C304 VTAIL.n218 B 0.019392f
C305 VTAIL.n219 B 0.010421f
C306 VTAIL.n220 B 0.011033f
C307 VTAIL.n221 B 0.02463f
C308 VTAIL.n222 B 0.02463f
C309 VTAIL.n223 B 0.011033f
C310 VTAIL.n224 B 0.010421f
C311 VTAIL.n225 B 0.019392f
C312 VTAIL.n226 B 0.019392f
C313 VTAIL.n227 B 0.010421f
C314 VTAIL.n228 B 0.011033f
C315 VTAIL.n229 B 0.02463f
C316 VTAIL.n230 B 0.02463f
C317 VTAIL.n231 B 0.011033f
C318 VTAIL.n232 B 0.010421f
C319 VTAIL.n233 B 0.019392f
C320 VTAIL.n234 B 0.019392f
C321 VTAIL.n235 B 0.010421f
C322 VTAIL.n236 B 0.011033f
C323 VTAIL.n237 B 0.02463f
C324 VTAIL.n238 B 0.02463f
C325 VTAIL.n239 B 0.011033f
C326 VTAIL.n240 B 0.010421f
C327 VTAIL.n241 B 0.019392f
C328 VTAIL.n242 B 0.019392f
C329 VTAIL.n243 B 0.010421f
C330 VTAIL.n244 B 0.011033f
C331 VTAIL.n245 B 0.02463f
C332 VTAIL.n246 B 0.052626f
C333 VTAIL.n247 B 0.011033f
C334 VTAIL.n248 B 0.010421f
C335 VTAIL.n249 B 0.045089f
C336 VTAIL.n250 B 0.029383f
C337 VTAIL.n251 B 1.05636f
C338 VTAIL.t7 B 0.174851f
C339 VTAIL.t9 B 0.174851f
C340 VTAIL.n252 B 1.49615f
C341 VTAIL.n253 B 0.352168f
C342 VTAIL.n254 B 0.026865f
C343 VTAIL.n255 B 0.019392f
C344 VTAIL.n256 B 0.010421f
C345 VTAIL.n257 B 0.02463f
C346 VTAIL.n258 B 0.011033f
C347 VTAIL.n259 B 0.019392f
C348 VTAIL.n260 B 0.010421f
C349 VTAIL.n261 B 0.02463f
C350 VTAIL.n262 B 0.010727f
C351 VTAIL.n263 B 0.019392f
C352 VTAIL.n264 B 0.010727f
C353 VTAIL.n265 B 0.010421f
C354 VTAIL.n266 B 0.02463f
C355 VTAIL.n267 B 0.02463f
C356 VTAIL.n268 B 0.011033f
C357 VTAIL.n269 B 0.019392f
C358 VTAIL.n270 B 0.010421f
C359 VTAIL.n271 B 0.02463f
C360 VTAIL.n272 B 0.011033f
C361 VTAIL.n273 B 0.927415f
C362 VTAIL.n274 B 0.010421f
C363 VTAIL.t11 B 0.041538f
C364 VTAIL.n275 B 0.135424f
C365 VTAIL.n276 B 0.017412f
C366 VTAIL.n277 B 0.018473f
C367 VTAIL.n278 B 0.02463f
C368 VTAIL.n279 B 0.011033f
C369 VTAIL.n280 B 0.010421f
C370 VTAIL.n281 B 0.019392f
C371 VTAIL.n282 B 0.019392f
C372 VTAIL.n283 B 0.010421f
C373 VTAIL.n284 B 0.011033f
C374 VTAIL.n285 B 0.02463f
C375 VTAIL.n286 B 0.02463f
C376 VTAIL.n287 B 0.011033f
C377 VTAIL.n288 B 0.010421f
C378 VTAIL.n289 B 0.019392f
C379 VTAIL.n290 B 0.019392f
C380 VTAIL.n291 B 0.010421f
C381 VTAIL.n292 B 0.011033f
C382 VTAIL.n293 B 0.02463f
C383 VTAIL.n294 B 0.02463f
C384 VTAIL.n295 B 0.011033f
C385 VTAIL.n296 B 0.010421f
C386 VTAIL.n297 B 0.019392f
C387 VTAIL.n298 B 0.019392f
C388 VTAIL.n299 B 0.010421f
C389 VTAIL.n300 B 0.011033f
C390 VTAIL.n301 B 0.02463f
C391 VTAIL.n302 B 0.02463f
C392 VTAIL.n303 B 0.011033f
C393 VTAIL.n304 B 0.010421f
C394 VTAIL.n305 B 0.019392f
C395 VTAIL.n306 B 0.019392f
C396 VTAIL.n307 B 0.010421f
C397 VTAIL.n308 B 0.011033f
C398 VTAIL.n309 B 0.02463f
C399 VTAIL.n310 B 0.052626f
C400 VTAIL.n311 B 0.011033f
C401 VTAIL.n312 B 0.010421f
C402 VTAIL.n313 B 0.045089f
C403 VTAIL.n314 B 0.029383f
C404 VTAIL.n315 B 0.126871f
C405 VTAIL.n316 B 0.026865f
C406 VTAIL.n317 B 0.019392f
C407 VTAIL.n318 B 0.010421f
C408 VTAIL.n319 B 0.02463f
C409 VTAIL.n320 B 0.011033f
C410 VTAIL.n321 B 0.019392f
C411 VTAIL.n322 B 0.010421f
C412 VTAIL.n323 B 0.02463f
C413 VTAIL.n324 B 0.010727f
C414 VTAIL.n325 B 0.019392f
C415 VTAIL.n326 B 0.010727f
C416 VTAIL.n327 B 0.010421f
C417 VTAIL.n328 B 0.02463f
C418 VTAIL.n329 B 0.02463f
C419 VTAIL.n330 B 0.011033f
C420 VTAIL.n331 B 0.019392f
C421 VTAIL.n332 B 0.010421f
C422 VTAIL.n333 B 0.02463f
C423 VTAIL.n334 B 0.011033f
C424 VTAIL.n335 B 0.927415f
C425 VTAIL.n336 B 0.010421f
C426 VTAIL.t15 B 0.041538f
C427 VTAIL.n337 B 0.135424f
C428 VTAIL.n338 B 0.017412f
C429 VTAIL.n339 B 0.018473f
C430 VTAIL.n340 B 0.02463f
C431 VTAIL.n341 B 0.011033f
C432 VTAIL.n342 B 0.010421f
C433 VTAIL.n343 B 0.019392f
C434 VTAIL.n344 B 0.019392f
C435 VTAIL.n345 B 0.010421f
C436 VTAIL.n346 B 0.011033f
C437 VTAIL.n347 B 0.02463f
C438 VTAIL.n348 B 0.02463f
C439 VTAIL.n349 B 0.011033f
C440 VTAIL.n350 B 0.010421f
C441 VTAIL.n351 B 0.019392f
C442 VTAIL.n352 B 0.019392f
C443 VTAIL.n353 B 0.010421f
C444 VTAIL.n354 B 0.011033f
C445 VTAIL.n355 B 0.02463f
C446 VTAIL.n356 B 0.02463f
C447 VTAIL.n357 B 0.011033f
C448 VTAIL.n358 B 0.010421f
C449 VTAIL.n359 B 0.019392f
C450 VTAIL.n360 B 0.019392f
C451 VTAIL.n361 B 0.010421f
C452 VTAIL.n362 B 0.011033f
C453 VTAIL.n363 B 0.02463f
C454 VTAIL.n364 B 0.02463f
C455 VTAIL.n365 B 0.011033f
C456 VTAIL.n366 B 0.010421f
C457 VTAIL.n367 B 0.019392f
C458 VTAIL.n368 B 0.019392f
C459 VTAIL.n369 B 0.010421f
C460 VTAIL.n370 B 0.011033f
C461 VTAIL.n371 B 0.02463f
C462 VTAIL.n372 B 0.052626f
C463 VTAIL.n373 B 0.011033f
C464 VTAIL.n374 B 0.010421f
C465 VTAIL.n375 B 0.045089f
C466 VTAIL.n376 B 0.029383f
C467 VTAIL.n377 B 0.126871f
C468 VTAIL.t4 B 0.174851f
C469 VTAIL.t1 B 0.174851f
C470 VTAIL.n378 B 1.49615f
C471 VTAIL.n379 B 0.352168f
C472 VTAIL.n380 B 0.026865f
C473 VTAIL.n381 B 0.019392f
C474 VTAIL.n382 B 0.010421f
C475 VTAIL.n383 B 0.02463f
C476 VTAIL.n384 B 0.011033f
C477 VTAIL.n385 B 0.019392f
C478 VTAIL.n386 B 0.010421f
C479 VTAIL.n387 B 0.02463f
C480 VTAIL.n388 B 0.010727f
C481 VTAIL.n389 B 0.019392f
C482 VTAIL.n390 B 0.010727f
C483 VTAIL.n391 B 0.010421f
C484 VTAIL.n392 B 0.02463f
C485 VTAIL.n393 B 0.02463f
C486 VTAIL.n394 B 0.011033f
C487 VTAIL.n395 B 0.019392f
C488 VTAIL.n396 B 0.010421f
C489 VTAIL.n397 B 0.02463f
C490 VTAIL.n398 B 0.011033f
C491 VTAIL.n399 B 0.927415f
C492 VTAIL.n400 B 0.010421f
C493 VTAIL.t3 B 0.041538f
C494 VTAIL.n401 B 0.135424f
C495 VTAIL.n402 B 0.017412f
C496 VTAIL.n403 B 0.018473f
C497 VTAIL.n404 B 0.02463f
C498 VTAIL.n405 B 0.011033f
C499 VTAIL.n406 B 0.010421f
C500 VTAIL.n407 B 0.019392f
C501 VTAIL.n408 B 0.019392f
C502 VTAIL.n409 B 0.010421f
C503 VTAIL.n410 B 0.011033f
C504 VTAIL.n411 B 0.02463f
C505 VTAIL.n412 B 0.02463f
C506 VTAIL.n413 B 0.011033f
C507 VTAIL.n414 B 0.010421f
C508 VTAIL.n415 B 0.019392f
C509 VTAIL.n416 B 0.019392f
C510 VTAIL.n417 B 0.010421f
C511 VTAIL.n418 B 0.011033f
C512 VTAIL.n419 B 0.02463f
C513 VTAIL.n420 B 0.02463f
C514 VTAIL.n421 B 0.011033f
C515 VTAIL.n422 B 0.010421f
C516 VTAIL.n423 B 0.019392f
C517 VTAIL.n424 B 0.019392f
C518 VTAIL.n425 B 0.010421f
C519 VTAIL.n426 B 0.011033f
C520 VTAIL.n427 B 0.02463f
C521 VTAIL.n428 B 0.02463f
C522 VTAIL.n429 B 0.011033f
C523 VTAIL.n430 B 0.010421f
C524 VTAIL.n431 B 0.019392f
C525 VTAIL.n432 B 0.019392f
C526 VTAIL.n433 B 0.010421f
C527 VTAIL.n434 B 0.011033f
C528 VTAIL.n435 B 0.02463f
C529 VTAIL.n436 B 0.052626f
C530 VTAIL.n437 B 0.011033f
C531 VTAIL.n438 B 0.010421f
C532 VTAIL.n439 B 0.045089f
C533 VTAIL.n440 B 0.029383f
C534 VTAIL.n441 B 1.05636f
C535 VTAIL.n442 B 0.026865f
C536 VTAIL.n443 B 0.019392f
C537 VTAIL.n444 B 0.010421f
C538 VTAIL.n445 B 0.02463f
C539 VTAIL.n446 B 0.011033f
C540 VTAIL.n447 B 0.019392f
C541 VTAIL.n448 B 0.010421f
C542 VTAIL.n449 B 0.02463f
C543 VTAIL.n450 B 0.010727f
C544 VTAIL.n451 B 0.019392f
C545 VTAIL.n452 B 0.011033f
C546 VTAIL.n453 B 0.02463f
C547 VTAIL.n454 B 0.011033f
C548 VTAIL.n455 B 0.019392f
C549 VTAIL.n456 B 0.010421f
C550 VTAIL.n457 B 0.02463f
C551 VTAIL.n458 B 0.011033f
C552 VTAIL.n459 B 0.927415f
C553 VTAIL.n460 B 0.010421f
C554 VTAIL.t8 B 0.041538f
C555 VTAIL.n461 B 0.135424f
C556 VTAIL.n462 B 0.017412f
C557 VTAIL.n463 B 0.018473f
C558 VTAIL.n464 B 0.02463f
C559 VTAIL.n465 B 0.011033f
C560 VTAIL.n466 B 0.010421f
C561 VTAIL.n467 B 0.019392f
C562 VTAIL.n468 B 0.019392f
C563 VTAIL.n469 B 0.010421f
C564 VTAIL.n470 B 0.011033f
C565 VTAIL.n471 B 0.02463f
C566 VTAIL.n472 B 0.02463f
C567 VTAIL.n473 B 0.011033f
C568 VTAIL.n474 B 0.010421f
C569 VTAIL.n475 B 0.019392f
C570 VTAIL.n476 B 0.019392f
C571 VTAIL.n477 B 0.010421f
C572 VTAIL.n478 B 0.010421f
C573 VTAIL.n479 B 0.011033f
C574 VTAIL.n480 B 0.02463f
C575 VTAIL.n481 B 0.02463f
C576 VTAIL.n482 B 0.02463f
C577 VTAIL.n483 B 0.010727f
C578 VTAIL.n484 B 0.010421f
C579 VTAIL.n485 B 0.019392f
C580 VTAIL.n486 B 0.019392f
C581 VTAIL.n487 B 0.010421f
C582 VTAIL.n488 B 0.011033f
C583 VTAIL.n489 B 0.02463f
C584 VTAIL.n490 B 0.02463f
C585 VTAIL.n491 B 0.011033f
C586 VTAIL.n492 B 0.010421f
C587 VTAIL.n493 B 0.019392f
C588 VTAIL.n494 B 0.019392f
C589 VTAIL.n495 B 0.010421f
C590 VTAIL.n496 B 0.011033f
C591 VTAIL.n497 B 0.02463f
C592 VTAIL.n498 B 0.052626f
C593 VTAIL.n499 B 0.011033f
C594 VTAIL.n500 B 0.010421f
C595 VTAIL.n501 B 0.045089f
C596 VTAIL.n502 B 0.029383f
C597 VTAIL.n503 B 1.05273f
C598 VDD2.t5 B 0.229732f
C599 VDD2.t2 B 0.229732f
C600 VDD2.n0 B 2.04431f
C601 VDD2.t3 B 0.229732f
C602 VDD2.t1 B 0.229732f
C603 VDD2.n1 B 2.04431f
C604 VDD2.n2 B 2.45691f
C605 VDD2.t0 B 0.229732f
C606 VDD2.t7 B 0.229732f
C607 VDD2.n3 B 2.04078f
C608 VDD2.n4 B 2.45419f
C609 VDD2.t4 B 0.229732f
C610 VDD2.t6 B 0.229732f
C611 VDD2.n5 B 2.04428f
C612 VN.n0 B 0.035311f
C613 VN.t6 B 1.28246f
C614 VN.n1 B 0.053934f
C615 VN.n2 B 0.035311f
C616 VN.t2 B 1.28246f
C617 VN.n3 B 0.524384f
C618 VN.t4 B 1.34777f
C619 VN.n4 B 0.550488f
C620 VN.n5 B 0.182782f
C621 VN.n6 B 0.053934f
C622 VN.n7 B 0.028546f
C623 VN.t1 B 1.28246f
C624 VN.n8 B 0.472841f
C625 VN.n9 B 0.053934f
C626 VN.n10 B 0.035311f
C627 VN.n11 B 0.035311f
C628 VN.n12 B 0.035311f
C629 VN.n13 B 0.028546f
C630 VN.n14 B 0.053934f
C631 VN.n15 B 0.52918f
C632 VN.n16 B 0.031637f
C633 VN.n17 B 0.035311f
C634 VN.t0 B 1.28246f
C635 VN.n18 B 0.053934f
C636 VN.n19 B 0.035311f
C637 VN.t7 B 1.28246f
C638 VN.n20 B 0.472841f
C639 VN.t5 B 1.28246f
C640 VN.n21 B 0.524384f
C641 VN.t3 B 1.34777f
C642 VN.n22 B 0.550488f
C643 VN.n23 B 0.182782f
C644 VN.n24 B 0.053934f
C645 VN.n25 B 0.028546f
C646 VN.n26 B 0.053934f
C647 VN.n27 B 0.035311f
C648 VN.n28 B 0.035311f
C649 VN.n29 B 0.035311f
C650 VN.n30 B 0.028546f
C651 VN.n31 B 0.053934f
C652 VN.n32 B 0.52918f
C653 VN.n33 B 1.57956f
.ends

