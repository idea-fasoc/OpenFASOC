* NGSPICE file created from diff_pair_sample_0066.ext - technology: sky130A

.subckt diff_pair_sample_0066 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=0 ps=0 w=18.06 l=1.49
X1 VTAIL.t7 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=2.9799 ps=18.39 w=18.06 l=1.49
X2 VTAIL.t6 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=2.9799 ps=18.39 w=18.06 l=1.49
X3 VTAIL.t2 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=2.9799 ps=18.39 w=18.06 l=1.49
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=0 ps=0 w=18.06 l=1.49
X5 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9799 pd=18.39 as=7.0434 ps=36.9 w=18.06 l=1.49
X6 VDD2.t0 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9799 pd=18.39 as=7.0434 ps=36.9 w=18.06 l=1.49
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=0 ps=0 w=18.06 l=1.49
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=0 ps=0 w=18.06 l=1.49
X9 VDD2.t3 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9799 pd=18.39 as=7.0434 ps=36.9 w=18.06 l=1.49
X10 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9799 pd=18.39 as=7.0434 ps=36.9 w=18.06 l=1.49
X11 VTAIL.t3 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0434 pd=36.9 as=2.9799 ps=18.39 w=18.06 l=1.49
R0 B.n844 B.n843 585
R1 B.n368 B.n111 585
R2 B.n367 B.n366 585
R3 B.n365 B.n364 585
R4 B.n363 B.n362 585
R5 B.n361 B.n360 585
R6 B.n359 B.n358 585
R7 B.n357 B.n356 585
R8 B.n355 B.n354 585
R9 B.n353 B.n352 585
R10 B.n351 B.n350 585
R11 B.n349 B.n348 585
R12 B.n347 B.n346 585
R13 B.n345 B.n344 585
R14 B.n343 B.n342 585
R15 B.n341 B.n340 585
R16 B.n339 B.n338 585
R17 B.n337 B.n336 585
R18 B.n335 B.n334 585
R19 B.n333 B.n332 585
R20 B.n331 B.n330 585
R21 B.n329 B.n328 585
R22 B.n327 B.n326 585
R23 B.n325 B.n324 585
R24 B.n323 B.n322 585
R25 B.n321 B.n320 585
R26 B.n319 B.n318 585
R27 B.n317 B.n316 585
R28 B.n315 B.n314 585
R29 B.n313 B.n312 585
R30 B.n311 B.n310 585
R31 B.n309 B.n308 585
R32 B.n307 B.n306 585
R33 B.n305 B.n304 585
R34 B.n303 B.n302 585
R35 B.n301 B.n300 585
R36 B.n299 B.n298 585
R37 B.n297 B.n296 585
R38 B.n295 B.n294 585
R39 B.n293 B.n292 585
R40 B.n291 B.n290 585
R41 B.n289 B.n288 585
R42 B.n287 B.n286 585
R43 B.n285 B.n284 585
R44 B.n283 B.n282 585
R45 B.n281 B.n280 585
R46 B.n279 B.n278 585
R47 B.n277 B.n276 585
R48 B.n275 B.n274 585
R49 B.n273 B.n272 585
R50 B.n271 B.n270 585
R51 B.n269 B.n268 585
R52 B.n267 B.n266 585
R53 B.n265 B.n264 585
R54 B.n263 B.n262 585
R55 B.n261 B.n260 585
R56 B.n259 B.n258 585
R57 B.n257 B.n256 585
R58 B.n255 B.n254 585
R59 B.n252 B.n251 585
R60 B.n250 B.n249 585
R61 B.n248 B.n247 585
R62 B.n246 B.n245 585
R63 B.n244 B.n243 585
R64 B.n242 B.n241 585
R65 B.n240 B.n239 585
R66 B.n238 B.n237 585
R67 B.n236 B.n235 585
R68 B.n234 B.n233 585
R69 B.n231 B.n230 585
R70 B.n229 B.n228 585
R71 B.n227 B.n226 585
R72 B.n225 B.n224 585
R73 B.n223 B.n222 585
R74 B.n221 B.n220 585
R75 B.n219 B.n218 585
R76 B.n217 B.n216 585
R77 B.n215 B.n214 585
R78 B.n213 B.n212 585
R79 B.n211 B.n210 585
R80 B.n209 B.n208 585
R81 B.n207 B.n206 585
R82 B.n205 B.n204 585
R83 B.n203 B.n202 585
R84 B.n201 B.n200 585
R85 B.n199 B.n198 585
R86 B.n197 B.n196 585
R87 B.n195 B.n194 585
R88 B.n193 B.n192 585
R89 B.n191 B.n190 585
R90 B.n189 B.n188 585
R91 B.n187 B.n186 585
R92 B.n185 B.n184 585
R93 B.n183 B.n182 585
R94 B.n181 B.n180 585
R95 B.n179 B.n178 585
R96 B.n177 B.n176 585
R97 B.n175 B.n174 585
R98 B.n173 B.n172 585
R99 B.n171 B.n170 585
R100 B.n169 B.n168 585
R101 B.n167 B.n166 585
R102 B.n165 B.n164 585
R103 B.n163 B.n162 585
R104 B.n161 B.n160 585
R105 B.n159 B.n158 585
R106 B.n157 B.n156 585
R107 B.n155 B.n154 585
R108 B.n153 B.n152 585
R109 B.n151 B.n150 585
R110 B.n149 B.n148 585
R111 B.n147 B.n146 585
R112 B.n145 B.n144 585
R113 B.n143 B.n142 585
R114 B.n141 B.n140 585
R115 B.n139 B.n138 585
R116 B.n137 B.n136 585
R117 B.n135 B.n134 585
R118 B.n133 B.n132 585
R119 B.n131 B.n130 585
R120 B.n129 B.n128 585
R121 B.n127 B.n126 585
R122 B.n125 B.n124 585
R123 B.n123 B.n122 585
R124 B.n121 B.n120 585
R125 B.n119 B.n118 585
R126 B.n117 B.n116 585
R127 B.n46 B.n45 585
R128 B.n842 B.n47 585
R129 B.n847 B.n47 585
R130 B.n841 B.n840 585
R131 B.n840 B.n43 585
R132 B.n839 B.n42 585
R133 B.n853 B.n42 585
R134 B.n838 B.n41 585
R135 B.n854 B.n41 585
R136 B.n837 B.n40 585
R137 B.n855 B.n40 585
R138 B.n836 B.n835 585
R139 B.n835 B.n39 585
R140 B.n834 B.n35 585
R141 B.n861 B.n35 585
R142 B.n833 B.n34 585
R143 B.n862 B.n34 585
R144 B.n832 B.n33 585
R145 B.n863 B.n33 585
R146 B.n831 B.n830 585
R147 B.n830 B.n29 585
R148 B.n829 B.n28 585
R149 B.n869 B.n28 585
R150 B.n828 B.n27 585
R151 B.n870 B.n27 585
R152 B.n827 B.n26 585
R153 B.n871 B.n26 585
R154 B.n826 B.n825 585
R155 B.n825 B.n22 585
R156 B.n824 B.n21 585
R157 B.n877 B.n21 585
R158 B.n823 B.n20 585
R159 B.n878 B.n20 585
R160 B.n822 B.n19 585
R161 B.n879 B.n19 585
R162 B.n821 B.n820 585
R163 B.n820 B.n15 585
R164 B.n819 B.n14 585
R165 B.n885 B.n14 585
R166 B.n818 B.n13 585
R167 B.n886 B.n13 585
R168 B.n817 B.n12 585
R169 B.n887 B.n12 585
R170 B.n816 B.n815 585
R171 B.n815 B.n8 585
R172 B.n814 B.n7 585
R173 B.n893 B.n7 585
R174 B.n813 B.n6 585
R175 B.n894 B.n6 585
R176 B.n812 B.n5 585
R177 B.n895 B.n5 585
R178 B.n811 B.n810 585
R179 B.n810 B.n4 585
R180 B.n809 B.n369 585
R181 B.n809 B.n808 585
R182 B.n799 B.n370 585
R183 B.n371 B.n370 585
R184 B.n801 B.n800 585
R185 B.n802 B.n801 585
R186 B.n798 B.n375 585
R187 B.n379 B.n375 585
R188 B.n797 B.n796 585
R189 B.n796 B.n795 585
R190 B.n377 B.n376 585
R191 B.n378 B.n377 585
R192 B.n788 B.n787 585
R193 B.n789 B.n788 585
R194 B.n786 B.n384 585
R195 B.n384 B.n383 585
R196 B.n785 B.n784 585
R197 B.n784 B.n783 585
R198 B.n386 B.n385 585
R199 B.n387 B.n386 585
R200 B.n776 B.n775 585
R201 B.n777 B.n776 585
R202 B.n774 B.n392 585
R203 B.n392 B.n391 585
R204 B.n773 B.n772 585
R205 B.n772 B.n771 585
R206 B.n394 B.n393 585
R207 B.n395 B.n394 585
R208 B.n764 B.n763 585
R209 B.n765 B.n764 585
R210 B.n762 B.n400 585
R211 B.n400 B.n399 585
R212 B.n761 B.n760 585
R213 B.n760 B.n759 585
R214 B.n402 B.n401 585
R215 B.n752 B.n402 585
R216 B.n751 B.n750 585
R217 B.n753 B.n751 585
R218 B.n749 B.n407 585
R219 B.n407 B.n406 585
R220 B.n748 B.n747 585
R221 B.n747 B.n746 585
R222 B.n409 B.n408 585
R223 B.n410 B.n409 585
R224 B.n739 B.n738 585
R225 B.n740 B.n739 585
R226 B.n413 B.n412 585
R227 B.n486 B.n485 585
R228 B.n487 B.n483 585
R229 B.n483 B.n414 585
R230 B.n489 B.n488 585
R231 B.n491 B.n482 585
R232 B.n494 B.n493 585
R233 B.n495 B.n481 585
R234 B.n497 B.n496 585
R235 B.n499 B.n480 585
R236 B.n502 B.n501 585
R237 B.n503 B.n479 585
R238 B.n505 B.n504 585
R239 B.n507 B.n478 585
R240 B.n510 B.n509 585
R241 B.n511 B.n477 585
R242 B.n513 B.n512 585
R243 B.n515 B.n476 585
R244 B.n518 B.n517 585
R245 B.n519 B.n475 585
R246 B.n521 B.n520 585
R247 B.n523 B.n474 585
R248 B.n526 B.n525 585
R249 B.n527 B.n473 585
R250 B.n529 B.n528 585
R251 B.n531 B.n472 585
R252 B.n534 B.n533 585
R253 B.n535 B.n471 585
R254 B.n537 B.n536 585
R255 B.n539 B.n470 585
R256 B.n542 B.n541 585
R257 B.n543 B.n469 585
R258 B.n545 B.n544 585
R259 B.n547 B.n468 585
R260 B.n550 B.n549 585
R261 B.n551 B.n467 585
R262 B.n553 B.n552 585
R263 B.n555 B.n466 585
R264 B.n558 B.n557 585
R265 B.n559 B.n465 585
R266 B.n561 B.n560 585
R267 B.n563 B.n464 585
R268 B.n566 B.n565 585
R269 B.n567 B.n463 585
R270 B.n569 B.n568 585
R271 B.n571 B.n462 585
R272 B.n574 B.n573 585
R273 B.n575 B.n461 585
R274 B.n577 B.n576 585
R275 B.n579 B.n460 585
R276 B.n582 B.n581 585
R277 B.n583 B.n459 585
R278 B.n585 B.n584 585
R279 B.n587 B.n458 585
R280 B.n590 B.n589 585
R281 B.n591 B.n457 585
R282 B.n593 B.n592 585
R283 B.n595 B.n456 585
R284 B.n598 B.n597 585
R285 B.n599 B.n453 585
R286 B.n602 B.n601 585
R287 B.n604 B.n452 585
R288 B.n607 B.n606 585
R289 B.n608 B.n451 585
R290 B.n610 B.n609 585
R291 B.n612 B.n450 585
R292 B.n615 B.n614 585
R293 B.n616 B.n449 585
R294 B.n618 B.n617 585
R295 B.n620 B.n448 585
R296 B.n623 B.n622 585
R297 B.n624 B.n444 585
R298 B.n626 B.n625 585
R299 B.n628 B.n443 585
R300 B.n631 B.n630 585
R301 B.n632 B.n442 585
R302 B.n634 B.n633 585
R303 B.n636 B.n441 585
R304 B.n639 B.n638 585
R305 B.n640 B.n440 585
R306 B.n642 B.n641 585
R307 B.n644 B.n439 585
R308 B.n647 B.n646 585
R309 B.n648 B.n438 585
R310 B.n650 B.n649 585
R311 B.n652 B.n437 585
R312 B.n655 B.n654 585
R313 B.n656 B.n436 585
R314 B.n658 B.n657 585
R315 B.n660 B.n435 585
R316 B.n663 B.n662 585
R317 B.n664 B.n434 585
R318 B.n666 B.n665 585
R319 B.n668 B.n433 585
R320 B.n671 B.n670 585
R321 B.n672 B.n432 585
R322 B.n674 B.n673 585
R323 B.n676 B.n431 585
R324 B.n679 B.n678 585
R325 B.n680 B.n430 585
R326 B.n682 B.n681 585
R327 B.n684 B.n429 585
R328 B.n687 B.n686 585
R329 B.n688 B.n428 585
R330 B.n690 B.n689 585
R331 B.n692 B.n427 585
R332 B.n695 B.n694 585
R333 B.n696 B.n426 585
R334 B.n698 B.n697 585
R335 B.n700 B.n425 585
R336 B.n703 B.n702 585
R337 B.n704 B.n424 585
R338 B.n706 B.n705 585
R339 B.n708 B.n423 585
R340 B.n711 B.n710 585
R341 B.n712 B.n422 585
R342 B.n714 B.n713 585
R343 B.n716 B.n421 585
R344 B.n719 B.n718 585
R345 B.n720 B.n420 585
R346 B.n722 B.n721 585
R347 B.n724 B.n419 585
R348 B.n727 B.n726 585
R349 B.n728 B.n418 585
R350 B.n730 B.n729 585
R351 B.n732 B.n417 585
R352 B.n733 B.n416 585
R353 B.n736 B.n735 585
R354 B.n737 B.n415 585
R355 B.n415 B.n414 585
R356 B.n742 B.n741 585
R357 B.n741 B.n740 585
R358 B.n743 B.n411 585
R359 B.n411 B.n410 585
R360 B.n745 B.n744 585
R361 B.n746 B.n745 585
R362 B.n405 B.n404 585
R363 B.n406 B.n405 585
R364 B.n755 B.n754 585
R365 B.n754 B.n753 585
R366 B.n756 B.n403 585
R367 B.n752 B.n403 585
R368 B.n758 B.n757 585
R369 B.n759 B.n758 585
R370 B.n398 B.n397 585
R371 B.n399 B.n398 585
R372 B.n767 B.n766 585
R373 B.n766 B.n765 585
R374 B.n768 B.n396 585
R375 B.n396 B.n395 585
R376 B.n770 B.n769 585
R377 B.n771 B.n770 585
R378 B.n390 B.n389 585
R379 B.n391 B.n390 585
R380 B.n779 B.n778 585
R381 B.n778 B.n777 585
R382 B.n780 B.n388 585
R383 B.n388 B.n387 585
R384 B.n782 B.n781 585
R385 B.n783 B.n782 585
R386 B.n382 B.n381 585
R387 B.n383 B.n382 585
R388 B.n791 B.n790 585
R389 B.n790 B.n789 585
R390 B.n792 B.n380 585
R391 B.n380 B.n378 585
R392 B.n794 B.n793 585
R393 B.n795 B.n794 585
R394 B.n374 B.n373 585
R395 B.n379 B.n374 585
R396 B.n804 B.n803 585
R397 B.n803 B.n802 585
R398 B.n805 B.n372 585
R399 B.n372 B.n371 585
R400 B.n807 B.n806 585
R401 B.n808 B.n807 585
R402 B.n2 B.n0 585
R403 B.n4 B.n2 585
R404 B.n3 B.n1 585
R405 B.n894 B.n3 585
R406 B.n892 B.n891 585
R407 B.n893 B.n892 585
R408 B.n890 B.n9 585
R409 B.n9 B.n8 585
R410 B.n889 B.n888 585
R411 B.n888 B.n887 585
R412 B.n11 B.n10 585
R413 B.n886 B.n11 585
R414 B.n884 B.n883 585
R415 B.n885 B.n884 585
R416 B.n882 B.n16 585
R417 B.n16 B.n15 585
R418 B.n881 B.n880 585
R419 B.n880 B.n879 585
R420 B.n18 B.n17 585
R421 B.n878 B.n18 585
R422 B.n876 B.n875 585
R423 B.n877 B.n876 585
R424 B.n874 B.n23 585
R425 B.n23 B.n22 585
R426 B.n873 B.n872 585
R427 B.n872 B.n871 585
R428 B.n25 B.n24 585
R429 B.n870 B.n25 585
R430 B.n868 B.n867 585
R431 B.n869 B.n868 585
R432 B.n866 B.n30 585
R433 B.n30 B.n29 585
R434 B.n865 B.n864 585
R435 B.n864 B.n863 585
R436 B.n32 B.n31 585
R437 B.n862 B.n32 585
R438 B.n860 B.n859 585
R439 B.n861 B.n860 585
R440 B.n858 B.n36 585
R441 B.n39 B.n36 585
R442 B.n857 B.n856 585
R443 B.n856 B.n855 585
R444 B.n38 B.n37 585
R445 B.n854 B.n38 585
R446 B.n852 B.n851 585
R447 B.n853 B.n852 585
R448 B.n850 B.n44 585
R449 B.n44 B.n43 585
R450 B.n849 B.n848 585
R451 B.n848 B.n847 585
R452 B.n897 B.n896 585
R453 B.n896 B.n895 585
R454 B.n741 B.n413 564.573
R455 B.n848 B.n46 564.573
R456 B.n739 B.n415 564.573
R457 B.n844 B.n47 564.573
R458 B.n445 B.t4 497.514
R459 B.n454 B.t15 497.514
R460 B.n114 B.t8 497.514
R461 B.n112 B.t12 497.514
R462 B.n445 B.t7 421.553
R463 B.n112 B.t13 421.553
R464 B.n454 B.t17 421.553
R465 B.n114 B.t10 421.553
R466 B.n446 B.t6 386.257
R467 B.n113 B.t14 386.257
R468 B.n455 B.t16 386.257
R469 B.n115 B.t11 386.257
R470 B.n846 B.n845 256.663
R471 B.n846 B.n110 256.663
R472 B.n846 B.n109 256.663
R473 B.n846 B.n108 256.663
R474 B.n846 B.n107 256.663
R475 B.n846 B.n106 256.663
R476 B.n846 B.n105 256.663
R477 B.n846 B.n104 256.663
R478 B.n846 B.n103 256.663
R479 B.n846 B.n102 256.663
R480 B.n846 B.n101 256.663
R481 B.n846 B.n100 256.663
R482 B.n846 B.n99 256.663
R483 B.n846 B.n98 256.663
R484 B.n846 B.n97 256.663
R485 B.n846 B.n96 256.663
R486 B.n846 B.n95 256.663
R487 B.n846 B.n94 256.663
R488 B.n846 B.n93 256.663
R489 B.n846 B.n92 256.663
R490 B.n846 B.n91 256.663
R491 B.n846 B.n90 256.663
R492 B.n846 B.n89 256.663
R493 B.n846 B.n88 256.663
R494 B.n846 B.n87 256.663
R495 B.n846 B.n86 256.663
R496 B.n846 B.n85 256.663
R497 B.n846 B.n84 256.663
R498 B.n846 B.n83 256.663
R499 B.n846 B.n82 256.663
R500 B.n846 B.n81 256.663
R501 B.n846 B.n80 256.663
R502 B.n846 B.n79 256.663
R503 B.n846 B.n78 256.663
R504 B.n846 B.n77 256.663
R505 B.n846 B.n76 256.663
R506 B.n846 B.n75 256.663
R507 B.n846 B.n74 256.663
R508 B.n846 B.n73 256.663
R509 B.n846 B.n72 256.663
R510 B.n846 B.n71 256.663
R511 B.n846 B.n70 256.663
R512 B.n846 B.n69 256.663
R513 B.n846 B.n68 256.663
R514 B.n846 B.n67 256.663
R515 B.n846 B.n66 256.663
R516 B.n846 B.n65 256.663
R517 B.n846 B.n64 256.663
R518 B.n846 B.n63 256.663
R519 B.n846 B.n62 256.663
R520 B.n846 B.n61 256.663
R521 B.n846 B.n60 256.663
R522 B.n846 B.n59 256.663
R523 B.n846 B.n58 256.663
R524 B.n846 B.n57 256.663
R525 B.n846 B.n56 256.663
R526 B.n846 B.n55 256.663
R527 B.n846 B.n54 256.663
R528 B.n846 B.n53 256.663
R529 B.n846 B.n52 256.663
R530 B.n846 B.n51 256.663
R531 B.n846 B.n50 256.663
R532 B.n846 B.n49 256.663
R533 B.n846 B.n48 256.663
R534 B.n484 B.n414 256.663
R535 B.n490 B.n414 256.663
R536 B.n492 B.n414 256.663
R537 B.n498 B.n414 256.663
R538 B.n500 B.n414 256.663
R539 B.n506 B.n414 256.663
R540 B.n508 B.n414 256.663
R541 B.n514 B.n414 256.663
R542 B.n516 B.n414 256.663
R543 B.n522 B.n414 256.663
R544 B.n524 B.n414 256.663
R545 B.n530 B.n414 256.663
R546 B.n532 B.n414 256.663
R547 B.n538 B.n414 256.663
R548 B.n540 B.n414 256.663
R549 B.n546 B.n414 256.663
R550 B.n548 B.n414 256.663
R551 B.n554 B.n414 256.663
R552 B.n556 B.n414 256.663
R553 B.n562 B.n414 256.663
R554 B.n564 B.n414 256.663
R555 B.n570 B.n414 256.663
R556 B.n572 B.n414 256.663
R557 B.n578 B.n414 256.663
R558 B.n580 B.n414 256.663
R559 B.n586 B.n414 256.663
R560 B.n588 B.n414 256.663
R561 B.n594 B.n414 256.663
R562 B.n596 B.n414 256.663
R563 B.n603 B.n414 256.663
R564 B.n605 B.n414 256.663
R565 B.n611 B.n414 256.663
R566 B.n613 B.n414 256.663
R567 B.n619 B.n414 256.663
R568 B.n621 B.n414 256.663
R569 B.n627 B.n414 256.663
R570 B.n629 B.n414 256.663
R571 B.n635 B.n414 256.663
R572 B.n637 B.n414 256.663
R573 B.n643 B.n414 256.663
R574 B.n645 B.n414 256.663
R575 B.n651 B.n414 256.663
R576 B.n653 B.n414 256.663
R577 B.n659 B.n414 256.663
R578 B.n661 B.n414 256.663
R579 B.n667 B.n414 256.663
R580 B.n669 B.n414 256.663
R581 B.n675 B.n414 256.663
R582 B.n677 B.n414 256.663
R583 B.n683 B.n414 256.663
R584 B.n685 B.n414 256.663
R585 B.n691 B.n414 256.663
R586 B.n693 B.n414 256.663
R587 B.n699 B.n414 256.663
R588 B.n701 B.n414 256.663
R589 B.n707 B.n414 256.663
R590 B.n709 B.n414 256.663
R591 B.n715 B.n414 256.663
R592 B.n717 B.n414 256.663
R593 B.n723 B.n414 256.663
R594 B.n725 B.n414 256.663
R595 B.n731 B.n414 256.663
R596 B.n734 B.n414 256.663
R597 B.n741 B.n411 163.367
R598 B.n745 B.n411 163.367
R599 B.n745 B.n405 163.367
R600 B.n754 B.n405 163.367
R601 B.n754 B.n403 163.367
R602 B.n758 B.n403 163.367
R603 B.n758 B.n398 163.367
R604 B.n766 B.n398 163.367
R605 B.n766 B.n396 163.367
R606 B.n770 B.n396 163.367
R607 B.n770 B.n390 163.367
R608 B.n778 B.n390 163.367
R609 B.n778 B.n388 163.367
R610 B.n782 B.n388 163.367
R611 B.n782 B.n382 163.367
R612 B.n790 B.n382 163.367
R613 B.n790 B.n380 163.367
R614 B.n794 B.n380 163.367
R615 B.n794 B.n374 163.367
R616 B.n803 B.n374 163.367
R617 B.n803 B.n372 163.367
R618 B.n807 B.n372 163.367
R619 B.n807 B.n2 163.367
R620 B.n896 B.n2 163.367
R621 B.n896 B.n3 163.367
R622 B.n892 B.n3 163.367
R623 B.n892 B.n9 163.367
R624 B.n888 B.n9 163.367
R625 B.n888 B.n11 163.367
R626 B.n884 B.n11 163.367
R627 B.n884 B.n16 163.367
R628 B.n880 B.n16 163.367
R629 B.n880 B.n18 163.367
R630 B.n876 B.n18 163.367
R631 B.n876 B.n23 163.367
R632 B.n872 B.n23 163.367
R633 B.n872 B.n25 163.367
R634 B.n868 B.n25 163.367
R635 B.n868 B.n30 163.367
R636 B.n864 B.n30 163.367
R637 B.n864 B.n32 163.367
R638 B.n860 B.n32 163.367
R639 B.n860 B.n36 163.367
R640 B.n856 B.n36 163.367
R641 B.n856 B.n38 163.367
R642 B.n852 B.n38 163.367
R643 B.n852 B.n44 163.367
R644 B.n848 B.n44 163.367
R645 B.n485 B.n483 163.367
R646 B.n489 B.n483 163.367
R647 B.n493 B.n491 163.367
R648 B.n497 B.n481 163.367
R649 B.n501 B.n499 163.367
R650 B.n505 B.n479 163.367
R651 B.n509 B.n507 163.367
R652 B.n513 B.n477 163.367
R653 B.n517 B.n515 163.367
R654 B.n521 B.n475 163.367
R655 B.n525 B.n523 163.367
R656 B.n529 B.n473 163.367
R657 B.n533 B.n531 163.367
R658 B.n537 B.n471 163.367
R659 B.n541 B.n539 163.367
R660 B.n545 B.n469 163.367
R661 B.n549 B.n547 163.367
R662 B.n553 B.n467 163.367
R663 B.n557 B.n555 163.367
R664 B.n561 B.n465 163.367
R665 B.n565 B.n563 163.367
R666 B.n569 B.n463 163.367
R667 B.n573 B.n571 163.367
R668 B.n577 B.n461 163.367
R669 B.n581 B.n579 163.367
R670 B.n585 B.n459 163.367
R671 B.n589 B.n587 163.367
R672 B.n593 B.n457 163.367
R673 B.n597 B.n595 163.367
R674 B.n602 B.n453 163.367
R675 B.n606 B.n604 163.367
R676 B.n610 B.n451 163.367
R677 B.n614 B.n612 163.367
R678 B.n618 B.n449 163.367
R679 B.n622 B.n620 163.367
R680 B.n626 B.n444 163.367
R681 B.n630 B.n628 163.367
R682 B.n634 B.n442 163.367
R683 B.n638 B.n636 163.367
R684 B.n642 B.n440 163.367
R685 B.n646 B.n644 163.367
R686 B.n650 B.n438 163.367
R687 B.n654 B.n652 163.367
R688 B.n658 B.n436 163.367
R689 B.n662 B.n660 163.367
R690 B.n666 B.n434 163.367
R691 B.n670 B.n668 163.367
R692 B.n674 B.n432 163.367
R693 B.n678 B.n676 163.367
R694 B.n682 B.n430 163.367
R695 B.n686 B.n684 163.367
R696 B.n690 B.n428 163.367
R697 B.n694 B.n692 163.367
R698 B.n698 B.n426 163.367
R699 B.n702 B.n700 163.367
R700 B.n706 B.n424 163.367
R701 B.n710 B.n708 163.367
R702 B.n714 B.n422 163.367
R703 B.n718 B.n716 163.367
R704 B.n722 B.n420 163.367
R705 B.n726 B.n724 163.367
R706 B.n730 B.n418 163.367
R707 B.n733 B.n732 163.367
R708 B.n735 B.n415 163.367
R709 B.n739 B.n409 163.367
R710 B.n747 B.n409 163.367
R711 B.n747 B.n407 163.367
R712 B.n751 B.n407 163.367
R713 B.n751 B.n402 163.367
R714 B.n760 B.n402 163.367
R715 B.n760 B.n400 163.367
R716 B.n764 B.n400 163.367
R717 B.n764 B.n394 163.367
R718 B.n772 B.n394 163.367
R719 B.n772 B.n392 163.367
R720 B.n776 B.n392 163.367
R721 B.n776 B.n386 163.367
R722 B.n784 B.n386 163.367
R723 B.n784 B.n384 163.367
R724 B.n788 B.n384 163.367
R725 B.n788 B.n377 163.367
R726 B.n796 B.n377 163.367
R727 B.n796 B.n375 163.367
R728 B.n801 B.n375 163.367
R729 B.n801 B.n370 163.367
R730 B.n809 B.n370 163.367
R731 B.n810 B.n809 163.367
R732 B.n810 B.n5 163.367
R733 B.n6 B.n5 163.367
R734 B.n7 B.n6 163.367
R735 B.n815 B.n7 163.367
R736 B.n815 B.n12 163.367
R737 B.n13 B.n12 163.367
R738 B.n14 B.n13 163.367
R739 B.n820 B.n14 163.367
R740 B.n820 B.n19 163.367
R741 B.n20 B.n19 163.367
R742 B.n21 B.n20 163.367
R743 B.n825 B.n21 163.367
R744 B.n825 B.n26 163.367
R745 B.n27 B.n26 163.367
R746 B.n28 B.n27 163.367
R747 B.n830 B.n28 163.367
R748 B.n830 B.n33 163.367
R749 B.n34 B.n33 163.367
R750 B.n35 B.n34 163.367
R751 B.n835 B.n35 163.367
R752 B.n835 B.n40 163.367
R753 B.n41 B.n40 163.367
R754 B.n42 B.n41 163.367
R755 B.n840 B.n42 163.367
R756 B.n840 B.n47 163.367
R757 B.n118 B.n117 163.367
R758 B.n122 B.n121 163.367
R759 B.n126 B.n125 163.367
R760 B.n130 B.n129 163.367
R761 B.n134 B.n133 163.367
R762 B.n138 B.n137 163.367
R763 B.n142 B.n141 163.367
R764 B.n146 B.n145 163.367
R765 B.n150 B.n149 163.367
R766 B.n154 B.n153 163.367
R767 B.n158 B.n157 163.367
R768 B.n162 B.n161 163.367
R769 B.n166 B.n165 163.367
R770 B.n170 B.n169 163.367
R771 B.n174 B.n173 163.367
R772 B.n178 B.n177 163.367
R773 B.n182 B.n181 163.367
R774 B.n186 B.n185 163.367
R775 B.n190 B.n189 163.367
R776 B.n194 B.n193 163.367
R777 B.n198 B.n197 163.367
R778 B.n202 B.n201 163.367
R779 B.n206 B.n205 163.367
R780 B.n210 B.n209 163.367
R781 B.n214 B.n213 163.367
R782 B.n218 B.n217 163.367
R783 B.n222 B.n221 163.367
R784 B.n226 B.n225 163.367
R785 B.n230 B.n229 163.367
R786 B.n235 B.n234 163.367
R787 B.n239 B.n238 163.367
R788 B.n243 B.n242 163.367
R789 B.n247 B.n246 163.367
R790 B.n251 B.n250 163.367
R791 B.n256 B.n255 163.367
R792 B.n260 B.n259 163.367
R793 B.n264 B.n263 163.367
R794 B.n268 B.n267 163.367
R795 B.n272 B.n271 163.367
R796 B.n276 B.n275 163.367
R797 B.n280 B.n279 163.367
R798 B.n284 B.n283 163.367
R799 B.n288 B.n287 163.367
R800 B.n292 B.n291 163.367
R801 B.n296 B.n295 163.367
R802 B.n300 B.n299 163.367
R803 B.n304 B.n303 163.367
R804 B.n308 B.n307 163.367
R805 B.n312 B.n311 163.367
R806 B.n316 B.n315 163.367
R807 B.n320 B.n319 163.367
R808 B.n324 B.n323 163.367
R809 B.n328 B.n327 163.367
R810 B.n332 B.n331 163.367
R811 B.n336 B.n335 163.367
R812 B.n340 B.n339 163.367
R813 B.n344 B.n343 163.367
R814 B.n348 B.n347 163.367
R815 B.n352 B.n351 163.367
R816 B.n356 B.n355 163.367
R817 B.n360 B.n359 163.367
R818 B.n364 B.n363 163.367
R819 B.n366 B.n111 163.367
R820 B.n484 B.n413 71.676
R821 B.n490 B.n489 71.676
R822 B.n493 B.n492 71.676
R823 B.n498 B.n497 71.676
R824 B.n501 B.n500 71.676
R825 B.n506 B.n505 71.676
R826 B.n509 B.n508 71.676
R827 B.n514 B.n513 71.676
R828 B.n517 B.n516 71.676
R829 B.n522 B.n521 71.676
R830 B.n525 B.n524 71.676
R831 B.n530 B.n529 71.676
R832 B.n533 B.n532 71.676
R833 B.n538 B.n537 71.676
R834 B.n541 B.n540 71.676
R835 B.n546 B.n545 71.676
R836 B.n549 B.n548 71.676
R837 B.n554 B.n553 71.676
R838 B.n557 B.n556 71.676
R839 B.n562 B.n561 71.676
R840 B.n565 B.n564 71.676
R841 B.n570 B.n569 71.676
R842 B.n573 B.n572 71.676
R843 B.n578 B.n577 71.676
R844 B.n581 B.n580 71.676
R845 B.n586 B.n585 71.676
R846 B.n589 B.n588 71.676
R847 B.n594 B.n593 71.676
R848 B.n597 B.n596 71.676
R849 B.n603 B.n602 71.676
R850 B.n606 B.n605 71.676
R851 B.n611 B.n610 71.676
R852 B.n614 B.n613 71.676
R853 B.n619 B.n618 71.676
R854 B.n622 B.n621 71.676
R855 B.n627 B.n626 71.676
R856 B.n630 B.n629 71.676
R857 B.n635 B.n634 71.676
R858 B.n638 B.n637 71.676
R859 B.n643 B.n642 71.676
R860 B.n646 B.n645 71.676
R861 B.n651 B.n650 71.676
R862 B.n654 B.n653 71.676
R863 B.n659 B.n658 71.676
R864 B.n662 B.n661 71.676
R865 B.n667 B.n666 71.676
R866 B.n670 B.n669 71.676
R867 B.n675 B.n674 71.676
R868 B.n678 B.n677 71.676
R869 B.n683 B.n682 71.676
R870 B.n686 B.n685 71.676
R871 B.n691 B.n690 71.676
R872 B.n694 B.n693 71.676
R873 B.n699 B.n698 71.676
R874 B.n702 B.n701 71.676
R875 B.n707 B.n706 71.676
R876 B.n710 B.n709 71.676
R877 B.n715 B.n714 71.676
R878 B.n718 B.n717 71.676
R879 B.n723 B.n722 71.676
R880 B.n726 B.n725 71.676
R881 B.n731 B.n730 71.676
R882 B.n734 B.n733 71.676
R883 B.n48 B.n46 71.676
R884 B.n118 B.n49 71.676
R885 B.n122 B.n50 71.676
R886 B.n126 B.n51 71.676
R887 B.n130 B.n52 71.676
R888 B.n134 B.n53 71.676
R889 B.n138 B.n54 71.676
R890 B.n142 B.n55 71.676
R891 B.n146 B.n56 71.676
R892 B.n150 B.n57 71.676
R893 B.n154 B.n58 71.676
R894 B.n158 B.n59 71.676
R895 B.n162 B.n60 71.676
R896 B.n166 B.n61 71.676
R897 B.n170 B.n62 71.676
R898 B.n174 B.n63 71.676
R899 B.n178 B.n64 71.676
R900 B.n182 B.n65 71.676
R901 B.n186 B.n66 71.676
R902 B.n190 B.n67 71.676
R903 B.n194 B.n68 71.676
R904 B.n198 B.n69 71.676
R905 B.n202 B.n70 71.676
R906 B.n206 B.n71 71.676
R907 B.n210 B.n72 71.676
R908 B.n214 B.n73 71.676
R909 B.n218 B.n74 71.676
R910 B.n222 B.n75 71.676
R911 B.n226 B.n76 71.676
R912 B.n230 B.n77 71.676
R913 B.n235 B.n78 71.676
R914 B.n239 B.n79 71.676
R915 B.n243 B.n80 71.676
R916 B.n247 B.n81 71.676
R917 B.n251 B.n82 71.676
R918 B.n256 B.n83 71.676
R919 B.n260 B.n84 71.676
R920 B.n264 B.n85 71.676
R921 B.n268 B.n86 71.676
R922 B.n272 B.n87 71.676
R923 B.n276 B.n88 71.676
R924 B.n280 B.n89 71.676
R925 B.n284 B.n90 71.676
R926 B.n288 B.n91 71.676
R927 B.n292 B.n92 71.676
R928 B.n296 B.n93 71.676
R929 B.n300 B.n94 71.676
R930 B.n304 B.n95 71.676
R931 B.n308 B.n96 71.676
R932 B.n312 B.n97 71.676
R933 B.n316 B.n98 71.676
R934 B.n320 B.n99 71.676
R935 B.n324 B.n100 71.676
R936 B.n328 B.n101 71.676
R937 B.n332 B.n102 71.676
R938 B.n336 B.n103 71.676
R939 B.n340 B.n104 71.676
R940 B.n344 B.n105 71.676
R941 B.n348 B.n106 71.676
R942 B.n352 B.n107 71.676
R943 B.n356 B.n108 71.676
R944 B.n360 B.n109 71.676
R945 B.n364 B.n110 71.676
R946 B.n845 B.n111 71.676
R947 B.n845 B.n844 71.676
R948 B.n366 B.n110 71.676
R949 B.n363 B.n109 71.676
R950 B.n359 B.n108 71.676
R951 B.n355 B.n107 71.676
R952 B.n351 B.n106 71.676
R953 B.n347 B.n105 71.676
R954 B.n343 B.n104 71.676
R955 B.n339 B.n103 71.676
R956 B.n335 B.n102 71.676
R957 B.n331 B.n101 71.676
R958 B.n327 B.n100 71.676
R959 B.n323 B.n99 71.676
R960 B.n319 B.n98 71.676
R961 B.n315 B.n97 71.676
R962 B.n311 B.n96 71.676
R963 B.n307 B.n95 71.676
R964 B.n303 B.n94 71.676
R965 B.n299 B.n93 71.676
R966 B.n295 B.n92 71.676
R967 B.n291 B.n91 71.676
R968 B.n287 B.n90 71.676
R969 B.n283 B.n89 71.676
R970 B.n279 B.n88 71.676
R971 B.n275 B.n87 71.676
R972 B.n271 B.n86 71.676
R973 B.n267 B.n85 71.676
R974 B.n263 B.n84 71.676
R975 B.n259 B.n83 71.676
R976 B.n255 B.n82 71.676
R977 B.n250 B.n81 71.676
R978 B.n246 B.n80 71.676
R979 B.n242 B.n79 71.676
R980 B.n238 B.n78 71.676
R981 B.n234 B.n77 71.676
R982 B.n229 B.n76 71.676
R983 B.n225 B.n75 71.676
R984 B.n221 B.n74 71.676
R985 B.n217 B.n73 71.676
R986 B.n213 B.n72 71.676
R987 B.n209 B.n71 71.676
R988 B.n205 B.n70 71.676
R989 B.n201 B.n69 71.676
R990 B.n197 B.n68 71.676
R991 B.n193 B.n67 71.676
R992 B.n189 B.n66 71.676
R993 B.n185 B.n65 71.676
R994 B.n181 B.n64 71.676
R995 B.n177 B.n63 71.676
R996 B.n173 B.n62 71.676
R997 B.n169 B.n61 71.676
R998 B.n165 B.n60 71.676
R999 B.n161 B.n59 71.676
R1000 B.n157 B.n58 71.676
R1001 B.n153 B.n57 71.676
R1002 B.n149 B.n56 71.676
R1003 B.n145 B.n55 71.676
R1004 B.n141 B.n54 71.676
R1005 B.n137 B.n53 71.676
R1006 B.n133 B.n52 71.676
R1007 B.n129 B.n51 71.676
R1008 B.n125 B.n50 71.676
R1009 B.n121 B.n49 71.676
R1010 B.n117 B.n48 71.676
R1011 B.n485 B.n484 71.676
R1012 B.n491 B.n490 71.676
R1013 B.n492 B.n481 71.676
R1014 B.n499 B.n498 71.676
R1015 B.n500 B.n479 71.676
R1016 B.n507 B.n506 71.676
R1017 B.n508 B.n477 71.676
R1018 B.n515 B.n514 71.676
R1019 B.n516 B.n475 71.676
R1020 B.n523 B.n522 71.676
R1021 B.n524 B.n473 71.676
R1022 B.n531 B.n530 71.676
R1023 B.n532 B.n471 71.676
R1024 B.n539 B.n538 71.676
R1025 B.n540 B.n469 71.676
R1026 B.n547 B.n546 71.676
R1027 B.n548 B.n467 71.676
R1028 B.n555 B.n554 71.676
R1029 B.n556 B.n465 71.676
R1030 B.n563 B.n562 71.676
R1031 B.n564 B.n463 71.676
R1032 B.n571 B.n570 71.676
R1033 B.n572 B.n461 71.676
R1034 B.n579 B.n578 71.676
R1035 B.n580 B.n459 71.676
R1036 B.n587 B.n586 71.676
R1037 B.n588 B.n457 71.676
R1038 B.n595 B.n594 71.676
R1039 B.n596 B.n453 71.676
R1040 B.n604 B.n603 71.676
R1041 B.n605 B.n451 71.676
R1042 B.n612 B.n611 71.676
R1043 B.n613 B.n449 71.676
R1044 B.n620 B.n619 71.676
R1045 B.n621 B.n444 71.676
R1046 B.n628 B.n627 71.676
R1047 B.n629 B.n442 71.676
R1048 B.n636 B.n635 71.676
R1049 B.n637 B.n440 71.676
R1050 B.n644 B.n643 71.676
R1051 B.n645 B.n438 71.676
R1052 B.n652 B.n651 71.676
R1053 B.n653 B.n436 71.676
R1054 B.n660 B.n659 71.676
R1055 B.n661 B.n434 71.676
R1056 B.n668 B.n667 71.676
R1057 B.n669 B.n432 71.676
R1058 B.n676 B.n675 71.676
R1059 B.n677 B.n430 71.676
R1060 B.n684 B.n683 71.676
R1061 B.n685 B.n428 71.676
R1062 B.n692 B.n691 71.676
R1063 B.n693 B.n426 71.676
R1064 B.n700 B.n699 71.676
R1065 B.n701 B.n424 71.676
R1066 B.n708 B.n707 71.676
R1067 B.n709 B.n422 71.676
R1068 B.n716 B.n715 71.676
R1069 B.n717 B.n420 71.676
R1070 B.n724 B.n723 71.676
R1071 B.n725 B.n418 71.676
R1072 B.n732 B.n731 71.676
R1073 B.n735 B.n734 71.676
R1074 B.n740 B.n414 63.6388
R1075 B.n847 B.n846 63.6388
R1076 B.n447 B.n446 59.5399
R1077 B.n600 B.n455 59.5399
R1078 B.n232 B.n115 59.5399
R1079 B.n253 B.n113 59.5399
R1080 B.n849 B.n45 36.6834
R1081 B.n843 B.n842 36.6834
R1082 B.n738 B.n737 36.6834
R1083 B.n742 B.n412 36.6834
R1084 B.n446 B.n445 35.2975
R1085 B.n455 B.n454 35.2975
R1086 B.n115 B.n114 35.2975
R1087 B.n113 B.n112 35.2975
R1088 B.n740 B.n410 32.0554
R1089 B.n746 B.n410 32.0554
R1090 B.n746 B.n406 32.0554
R1091 B.n753 B.n406 32.0554
R1092 B.n753 B.n752 32.0554
R1093 B.n759 B.n399 32.0554
R1094 B.n765 B.n399 32.0554
R1095 B.n765 B.n395 32.0554
R1096 B.n771 B.n395 32.0554
R1097 B.n771 B.n391 32.0554
R1098 B.n777 B.n391 32.0554
R1099 B.n777 B.n387 32.0554
R1100 B.n783 B.n387 32.0554
R1101 B.n789 B.n383 32.0554
R1102 B.n789 B.n378 32.0554
R1103 B.n795 B.n378 32.0554
R1104 B.n795 B.n379 32.0554
R1105 B.n802 B.n371 32.0554
R1106 B.n808 B.n371 32.0554
R1107 B.n808 B.n4 32.0554
R1108 B.n895 B.n4 32.0554
R1109 B.n895 B.n894 32.0554
R1110 B.n894 B.n893 32.0554
R1111 B.n893 B.n8 32.0554
R1112 B.n887 B.n8 32.0554
R1113 B.n886 B.n885 32.0554
R1114 B.n885 B.n15 32.0554
R1115 B.n879 B.n15 32.0554
R1116 B.n879 B.n878 32.0554
R1117 B.n877 B.n22 32.0554
R1118 B.n871 B.n22 32.0554
R1119 B.n871 B.n870 32.0554
R1120 B.n870 B.n869 32.0554
R1121 B.n869 B.n29 32.0554
R1122 B.n863 B.n29 32.0554
R1123 B.n863 B.n862 32.0554
R1124 B.n862 B.n861 32.0554
R1125 B.n855 B.n39 32.0554
R1126 B.n855 B.n854 32.0554
R1127 B.n854 B.n853 32.0554
R1128 B.n853 B.n43 32.0554
R1129 B.n847 B.n43 32.0554
R1130 B.n752 B.t5 25.9272
R1131 B.n39 B.t9 25.9272
R1132 B.n379 B.t0 23.0989
R1133 B.t2 B.n886 23.0989
R1134 B.t3 B.n383 20.2705
R1135 B.n878 B.t1 20.2705
R1136 B B.n897 18.0485
R1137 B.n783 B.t3 11.7854
R1138 B.t1 B.n877 11.7854
R1139 B.n116 B.n45 10.6151
R1140 B.n119 B.n116 10.6151
R1141 B.n120 B.n119 10.6151
R1142 B.n123 B.n120 10.6151
R1143 B.n124 B.n123 10.6151
R1144 B.n127 B.n124 10.6151
R1145 B.n128 B.n127 10.6151
R1146 B.n131 B.n128 10.6151
R1147 B.n132 B.n131 10.6151
R1148 B.n135 B.n132 10.6151
R1149 B.n136 B.n135 10.6151
R1150 B.n139 B.n136 10.6151
R1151 B.n140 B.n139 10.6151
R1152 B.n143 B.n140 10.6151
R1153 B.n144 B.n143 10.6151
R1154 B.n147 B.n144 10.6151
R1155 B.n148 B.n147 10.6151
R1156 B.n151 B.n148 10.6151
R1157 B.n152 B.n151 10.6151
R1158 B.n155 B.n152 10.6151
R1159 B.n156 B.n155 10.6151
R1160 B.n159 B.n156 10.6151
R1161 B.n160 B.n159 10.6151
R1162 B.n163 B.n160 10.6151
R1163 B.n164 B.n163 10.6151
R1164 B.n167 B.n164 10.6151
R1165 B.n168 B.n167 10.6151
R1166 B.n171 B.n168 10.6151
R1167 B.n172 B.n171 10.6151
R1168 B.n175 B.n172 10.6151
R1169 B.n176 B.n175 10.6151
R1170 B.n179 B.n176 10.6151
R1171 B.n180 B.n179 10.6151
R1172 B.n183 B.n180 10.6151
R1173 B.n184 B.n183 10.6151
R1174 B.n187 B.n184 10.6151
R1175 B.n188 B.n187 10.6151
R1176 B.n191 B.n188 10.6151
R1177 B.n192 B.n191 10.6151
R1178 B.n195 B.n192 10.6151
R1179 B.n196 B.n195 10.6151
R1180 B.n199 B.n196 10.6151
R1181 B.n200 B.n199 10.6151
R1182 B.n203 B.n200 10.6151
R1183 B.n204 B.n203 10.6151
R1184 B.n207 B.n204 10.6151
R1185 B.n208 B.n207 10.6151
R1186 B.n211 B.n208 10.6151
R1187 B.n212 B.n211 10.6151
R1188 B.n215 B.n212 10.6151
R1189 B.n216 B.n215 10.6151
R1190 B.n219 B.n216 10.6151
R1191 B.n220 B.n219 10.6151
R1192 B.n223 B.n220 10.6151
R1193 B.n224 B.n223 10.6151
R1194 B.n227 B.n224 10.6151
R1195 B.n228 B.n227 10.6151
R1196 B.n231 B.n228 10.6151
R1197 B.n236 B.n233 10.6151
R1198 B.n237 B.n236 10.6151
R1199 B.n240 B.n237 10.6151
R1200 B.n241 B.n240 10.6151
R1201 B.n244 B.n241 10.6151
R1202 B.n245 B.n244 10.6151
R1203 B.n248 B.n245 10.6151
R1204 B.n249 B.n248 10.6151
R1205 B.n252 B.n249 10.6151
R1206 B.n257 B.n254 10.6151
R1207 B.n258 B.n257 10.6151
R1208 B.n261 B.n258 10.6151
R1209 B.n262 B.n261 10.6151
R1210 B.n265 B.n262 10.6151
R1211 B.n266 B.n265 10.6151
R1212 B.n269 B.n266 10.6151
R1213 B.n270 B.n269 10.6151
R1214 B.n273 B.n270 10.6151
R1215 B.n274 B.n273 10.6151
R1216 B.n277 B.n274 10.6151
R1217 B.n278 B.n277 10.6151
R1218 B.n281 B.n278 10.6151
R1219 B.n282 B.n281 10.6151
R1220 B.n285 B.n282 10.6151
R1221 B.n286 B.n285 10.6151
R1222 B.n289 B.n286 10.6151
R1223 B.n290 B.n289 10.6151
R1224 B.n293 B.n290 10.6151
R1225 B.n294 B.n293 10.6151
R1226 B.n297 B.n294 10.6151
R1227 B.n298 B.n297 10.6151
R1228 B.n301 B.n298 10.6151
R1229 B.n302 B.n301 10.6151
R1230 B.n305 B.n302 10.6151
R1231 B.n306 B.n305 10.6151
R1232 B.n309 B.n306 10.6151
R1233 B.n310 B.n309 10.6151
R1234 B.n313 B.n310 10.6151
R1235 B.n314 B.n313 10.6151
R1236 B.n317 B.n314 10.6151
R1237 B.n318 B.n317 10.6151
R1238 B.n321 B.n318 10.6151
R1239 B.n322 B.n321 10.6151
R1240 B.n325 B.n322 10.6151
R1241 B.n326 B.n325 10.6151
R1242 B.n329 B.n326 10.6151
R1243 B.n330 B.n329 10.6151
R1244 B.n333 B.n330 10.6151
R1245 B.n334 B.n333 10.6151
R1246 B.n337 B.n334 10.6151
R1247 B.n338 B.n337 10.6151
R1248 B.n341 B.n338 10.6151
R1249 B.n342 B.n341 10.6151
R1250 B.n345 B.n342 10.6151
R1251 B.n346 B.n345 10.6151
R1252 B.n349 B.n346 10.6151
R1253 B.n350 B.n349 10.6151
R1254 B.n353 B.n350 10.6151
R1255 B.n354 B.n353 10.6151
R1256 B.n357 B.n354 10.6151
R1257 B.n358 B.n357 10.6151
R1258 B.n361 B.n358 10.6151
R1259 B.n362 B.n361 10.6151
R1260 B.n365 B.n362 10.6151
R1261 B.n367 B.n365 10.6151
R1262 B.n368 B.n367 10.6151
R1263 B.n843 B.n368 10.6151
R1264 B.n738 B.n408 10.6151
R1265 B.n748 B.n408 10.6151
R1266 B.n749 B.n748 10.6151
R1267 B.n750 B.n749 10.6151
R1268 B.n750 B.n401 10.6151
R1269 B.n761 B.n401 10.6151
R1270 B.n762 B.n761 10.6151
R1271 B.n763 B.n762 10.6151
R1272 B.n763 B.n393 10.6151
R1273 B.n773 B.n393 10.6151
R1274 B.n774 B.n773 10.6151
R1275 B.n775 B.n774 10.6151
R1276 B.n775 B.n385 10.6151
R1277 B.n785 B.n385 10.6151
R1278 B.n786 B.n785 10.6151
R1279 B.n787 B.n786 10.6151
R1280 B.n787 B.n376 10.6151
R1281 B.n797 B.n376 10.6151
R1282 B.n798 B.n797 10.6151
R1283 B.n800 B.n798 10.6151
R1284 B.n800 B.n799 10.6151
R1285 B.n799 B.n369 10.6151
R1286 B.n811 B.n369 10.6151
R1287 B.n812 B.n811 10.6151
R1288 B.n813 B.n812 10.6151
R1289 B.n814 B.n813 10.6151
R1290 B.n816 B.n814 10.6151
R1291 B.n817 B.n816 10.6151
R1292 B.n818 B.n817 10.6151
R1293 B.n819 B.n818 10.6151
R1294 B.n821 B.n819 10.6151
R1295 B.n822 B.n821 10.6151
R1296 B.n823 B.n822 10.6151
R1297 B.n824 B.n823 10.6151
R1298 B.n826 B.n824 10.6151
R1299 B.n827 B.n826 10.6151
R1300 B.n828 B.n827 10.6151
R1301 B.n829 B.n828 10.6151
R1302 B.n831 B.n829 10.6151
R1303 B.n832 B.n831 10.6151
R1304 B.n833 B.n832 10.6151
R1305 B.n834 B.n833 10.6151
R1306 B.n836 B.n834 10.6151
R1307 B.n837 B.n836 10.6151
R1308 B.n838 B.n837 10.6151
R1309 B.n839 B.n838 10.6151
R1310 B.n841 B.n839 10.6151
R1311 B.n842 B.n841 10.6151
R1312 B.n486 B.n412 10.6151
R1313 B.n487 B.n486 10.6151
R1314 B.n488 B.n487 10.6151
R1315 B.n488 B.n482 10.6151
R1316 B.n494 B.n482 10.6151
R1317 B.n495 B.n494 10.6151
R1318 B.n496 B.n495 10.6151
R1319 B.n496 B.n480 10.6151
R1320 B.n502 B.n480 10.6151
R1321 B.n503 B.n502 10.6151
R1322 B.n504 B.n503 10.6151
R1323 B.n504 B.n478 10.6151
R1324 B.n510 B.n478 10.6151
R1325 B.n511 B.n510 10.6151
R1326 B.n512 B.n511 10.6151
R1327 B.n512 B.n476 10.6151
R1328 B.n518 B.n476 10.6151
R1329 B.n519 B.n518 10.6151
R1330 B.n520 B.n519 10.6151
R1331 B.n520 B.n474 10.6151
R1332 B.n526 B.n474 10.6151
R1333 B.n527 B.n526 10.6151
R1334 B.n528 B.n527 10.6151
R1335 B.n528 B.n472 10.6151
R1336 B.n534 B.n472 10.6151
R1337 B.n535 B.n534 10.6151
R1338 B.n536 B.n535 10.6151
R1339 B.n536 B.n470 10.6151
R1340 B.n542 B.n470 10.6151
R1341 B.n543 B.n542 10.6151
R1342 B.n544 B.n543 10.6151
R1343 B.n544 B.n468 10.6151
R1344 B.n550 B.n468 10.6151
R1345 B.n551 B.n550 10.6151
R1346 B.n552 B.n551 10.6151
R1347 B.n552 B.n466 10.6151
R1348 B.n558 B.n466 10.6151
R1349 B.n559 B.n558 10.6151
R1350 B.n560 B.n559 10.6151
R1351 B.n560 B.n464 10.6151
R1352 B.n566 B.n464 10.6151
R1353 B.n567 B.n566 10.6151
R1354 B.n568 B.n567 10.6151
R1355 B.n568 B.n462 10.6151
R1356 B.n574 B.n462 10.6151
R1357 B.n575 B.n574 10.6151
R1358 B.n576 B.n575 10.6151
R1359 B.n576 B.n460 10.6151
R1360 B.n582 B.n460 10.6151
R1361 B.n583 B.n582 10.6151
R1362 B.n584 B.n583 10.6151
R1363 B.n584 B.n458 10.6151
R1364 B.n590 B.n458 10.6151
R1365 B.n591 B.n590 10.6151
R1366 B.n592 B.n591 10.6151
R1367 B.n592 B.n456 10.6151
R1368 B.n598 B.n456 10.6151
R1369 B.n599 B.n598 10.6151
R1370 B.n601 B.n452 10.6151
R1371 B.n607 B.n452 10.6151
R1372 B.n608 B.n607 10.6151
R1373 B.n609 B.n608 10.6151
R1374 B.n609 B.n450 10.6151
R1375 B.n615 B.n450 10.6151
R1376 B.n616 B.n615 10.6151
R1377 B.n617 B.n616 10.6151
R1378 B.n617 B.n448 10.6151
R1379 B.n624 B.n623 10.6151
R1380 B.n625 B.n624 10.6151
R1381 B.n625 B.n443 10.6151
R1382 B.n631 B.n443 10.6151
R1383 B.n632 B.n631 10.6151
R1384 B.n633 B.n632 10.6151
R1385 B.n633 B.n441 10.6151
R1386 B.n639 B.n441 10.6151
R1387 B.n640 B.n639 10.6151
R1388 B.n641 B.n640 10.6151
R1389 B.n641 B.n439 10.6151
R1390 B.n647 B.n439 10.6151
R1391 B.n648 B.n647 10.6151
R1392 B.n649 B.n648 10.6151
R1393 B.n649 B.n437 10.6151
R1394 B.n655 B.n437 10.6151
R1395 B.n656 B.n655 10.6151
R1396 B.n657 B.n656 10.6151
R1397 B.n657 B.n435 10.6151
R1398 B.n663 B.n435 10.6151
R1399 B.n664 B.n663 10.6151
R1400 B.n665 B.n664 10.6151
R1401 B.n665 B.n433 10.6151
R1402 B.n671 B.n433 10.6151
R1403 B.n672 B.n671 10.6151
R1404 B.n673 B.n672 10.6151
R1405 B.n673 B.n431 10.6151
R1406 B.n679 B.n431 10.6151
R1407 B.n680 B.n679 10.6151
R1408 B.n681 B.n680 10.6151
R1409 B.n681 B.n429 10.6151
R1410 B.n687 B.n429 10.6151
R1411 B.n688 B.n687 10.6151
R1412 B.n689 B.n688 10.6151
R1413 B.n689 B.n427 10.6151
R1414 B.n695 B.n427 10.6151
R1415 B.n696 B.n695 10.6151
R1416 B.n697 B.n696 10.6151
R1417 B.n697 B.n425 10.6151
R1418 B.n703 B.n425 10.6151
R1419 B.n704 B.n703 10.6151
R1420 B.n705 B.n704 10.6151
R1421 B.n705 B.n423 10.6151
R1422 B.n711 B.n423 10.6151
R1423 B.n712 B.n711 10.6151
R1424 B.n713 B.n712 10.6151
R1425 B.n713 B.n421 10.6151
R1426 B.n719 B.n421 10.6151
R1427 B.n720 B.n719 10.6151
R1428 B.n721 B.n720 10.6151
R1429 B.n721 B.n419 10.6151
R1430 B.n727 B.n419 10.6151
R1431 B.n728 B.n727 10.6151
R1432 B.n729 B.n728 10.6151
R1433 B.n729 B.n417 10.6151
R1434 B.n417 B.n416 10.6151
R1435 B.n736 B.n416 10.6151
R1436 B.n737 B.n736 10.6151
R1437 B.n743 B.n742 10.6151
R1438 B.n744 B.n743 10.6151
R1439 B.n744 B.n404 10.6151
R1440 B.n755 B.n404 10.6151
R1441 B.n756 B.n755 10.6151
R1442 B.n757 B.n756 10.6151
R1443 B.n757 B.n397 10.6151
R1444 B.n767 B.n397 10.6151
R1445 B.n768 B.n767 10.6151
R1446 B.n769 B.n768 10.6151
R1447 B.n769 B.n389 10.6151
R1448 B.n779 B.n389 10.6151
R1449 B.n780 B.n779 10.6151
R1450 B.n781 B.n780 10.6151
R1451 B.n781 B.n381 10.6151
R1452 B.n791 B.n381 10.6151
R1453 B.n792 B.n791 10.6151
R1454 B.n793 B.n792 10.6151
R1455 B.n793 B.n373 10.6151
R1456 B.n804 B.n373 10.6151
R1457 B.n805 B.n804 10.6151
R1458 B.n806 B.n805 10.6151
R1459 B.n806 B.n0 10.6151
R1460 B.n891 B.n1 10.6151
R1461 B.n891 B.n890 10.6151
R1462 B.n890 B.n889 10.6151
R1463 B.n889 B.n10 10.6151
R1464 B.n883 B.n10 10.6151
R1465 B.n883 B.n882 10.6151
R1466 B.n882 B.n881 10.6151
R1467 B.n881 B.n17 10.6151
R1468 B.n875 B.n17 10.6151
R1469 B.n875 B.n874 10.6151
R1470 B.n874 B.n873 10.6151
R1471 B.n873 B.n24 10.6151
R1472 B.n867 B.n24 10.6151
R1473 B.n867 B.n866 10.6151
R1474 B.n866 B.n865 10.6151
R1475 B.n865 B.n31 10.6151
R1476 B.n859 B.n31 10.6151
R1477 B.n859 B.n858 10.6151
R1478 B.n858 B.n857 10.6151
R1479 B.n857 B.n37 10.6151
R1480 B.n851 B.n37 10.6151
R1481 B.n851 B.n850 10.6151
R1482 B.n850 B.n849 10.6151
R1483 B.n232 B.n231 9.36635
R1484 B.n254 B.n253 9.36635
R1485 B.n600 B.n599 9.36635
R1486 B.n623 B.n447 9.36635
R1487 B.n802 B.t0 8.957
R1488 B.n887 B.t2 8.957
R1489 B.n759 B.t5 6.12863
R1490 B.n861 B.t9 6.12863
R1491 B.n897 B.n0 2.81026
R1492 B.n897 B.n1 2.81026
R1493 B.n233 B.n232 1.24928
R1494 B.n253 B.n252 1.24928
R1495 B.n601 B.n600 1.24928
R1496 B.n448 B.n447 1.24928
R1497 VN.n0 VN.t1 328.408
R1498 VN.n1 VN.t3 328.408
R1499 VN.n0 VN.t2 328.091
R1500 VN.n1 VN.t0 328.091
R1501 VN VN.n1 60.8321
R1502 VN VN.n0 13.0784
R1503 VDD2.n2 VDD2.n0 107.588
R1504 VDD2.n2 VDD2.n1 63.5967
R1505 VDD2.n1 VDD2.t1 1.09685
R1506 VDD2.n1 VDD2.t3 1.09685
R1507 VDD2.n0 VDD2.t2 1.09685
R1508 VDD2.n0 VDD2.t0 1.09685
R1509 VDD2 VDD2.n2 0.0586897
R1510 VTAIL.n798 VTAIL.n797 289.615
R1511 VTAIL.n98 VTAIL.n97 289.615
R1512 VTAIL.n198 VTAIL.n197 289.615
R1513 VTAIL.n298 VTAIL.n297 289.615
R1514 VTAIL.n698 VTAIL.n697 289.615
R1515 VTAIL.n598 VTAIL.n597 289.615
R1516 VTAIL.n498 VTAIL.n497 289.615
R1517 VTAIL.n398 VTAIL.n397 289.615
R1518 VTAIL.n733 VTAIL.n732 185
R1519 VTAIL.n730 VTAIL.n729 185
R1520 VTAIL.n739 VTAIL.n738 185
R1521 VTAIL.n741 VTAIL.n740 185
R1522 VTAIL.n726 VTAIL.n725 185
R1523 VTAIL.n747 VTAIL.n746 185
R1524 VTAIL.n750 VTAIL.n749 185
R1525 VTAIL.n748 VTAIL.n722 185
R1526 VTAIL.n755 VTAIL.n721 185
R1527 VTAIL.n757 VTAIL.n756 185
R1528 VTAIL.n759 VTAIL.n758 185
R1529 VTAIL.n718 VTAIL.n717 185
R1530 VTAIL.n765 VTAIL.n764 185
R1531 VTAIL.n767 VTAIL.n766 185
R1532 VTAIL.n714 VTAIL.n713 185
R1533 VTAIL.n773 VTAIL.n772 185
R1534 VTAIL.n775 VTAIL.n774 185
R1535 VTAIL.n710 VTAIL.n709 185
R1536 VTAIL.n781 VTAIL.n780 185
R1537 VTAIL.n783 VTAIL.n782 185
R1538 VTAIL.n706 VTAIL.n705 185
R1539 VTAIL.n789 VTAIL.n788 185
R1540 VTAIL.n791 VTAIL.n790 185
R1541 VTAIL.n702 VTAIL.n701 185
R1542 VTAIL.n797 VTAIL.n796 185
R1543 VTAIL.n33 VTAIL.n32 185
R1544 VTAIL.n30 VTAIL.n29 185
R1545 VTAIL.n39 VTAIL.n38 185
R1546 VTAIL.n41 VTAIL.n40 185
R1547 VTAIL.n26 VTAIL.n25 185
R1548 VTAIL.n47 VTAIL.n46 185
R1549 VTAIL.n50 VTAIL.n49 185
R1550 VTAIL.n48 VTAIL.n22 185
R1551 VTAIL.n55 VTAIL.n21 185
R1552 VTAIL.n57 VTAIL.n56 185
R1553 VTAIL.n59 VTAIL.n58 185
R1554 VTAIL.n18 VTAIL.n17 185
R1555 VTAIL.n65 VTAIL.n64 185
R1556 VTAIL.n67 VTAIL.n66 185
R1557 VTAIL.n14 VTAIL.n13 185
R1558 VTAIL.n73 VTAIL.n72 185
R1559 VTAIL.n75 VTAIL.n74 185
R1560 VTAIL.n10 VTAIL.n9 185
R1561 VTAIL.n81 VTAIL.n80 185
R1562 VTAIL.n83 VTAIL.n82 185
R1563 VTAIL.n6 VTAIL.n5 185
R1564 VTAIL.n89 VTAIL.n88 185
R1565 VTAIL.n91 VTAIL.n90 185
R1566 VTAIL.n2 VTAIL.n1 185
R1567 VTAIL.n97 VTAIL.n96 185
R1568 VTAIL.n133 VTAIL.n132 185
R1569 VTAIL.n130 VTAIL.n129 185
R1570 VTAIL.n139 VTAIL.n138 185
R1571 VTAIL.n141 VTAIL.n140 185
R1572 VTAIL.n126 VTAIL.n125 185
R1573 VTAIL.n147 VTAIL.n146 185
R1574 VTAIL.n150 VTAIL.n149 185
R1575 VTAIL.n148 VTAIL.n122 185
R1576 VTAIL.n155 VTAIL.n121 185
R1577 VTAIL.n157 VTAIL.n156 185
R1578 VTAIL.n159 VTAIL.n158 185
R1579 VTAIL.n118 VTAIL.n117 185
R1580 VTAIL.n165 VTAIL.n164 185
R1581 VTAIL.n167 VTAIL.n166 185
R1582 VTAIL.n114 VTAIL.n113 185
R1583 VTAIL.n173 VTAIL.n172 185
R1584 VTAIL.n175 VTAIL.n174 185
R1585 VTAIL.n110 VTAIL.n109 185
R1586 VTAIL.n181 VTAIL.n180 185
R1587 VTAIL.n183 VTAIL.n182 185
R1588 VTAIL.n106 VTAIL.n105 185
R1589 VTAIL.n189 VTAIL.n188 185
R1590 VTAIL.n191 VTAIL.n190 185
R1591 VTAIL.n102 VTAIL.n101 185
R1592 VTAIL.n197 VTAIL.n196 185
R1593 VTAIL.n233 VTAIL.n232 185
R1594 VTAIL.n230 VTAIL.n229 185
R1595 VTAIL.n239 VTAIL.n238 185
R1596 VTAIL.n241 VTAIL.n240 185
R1597 VTAIL.n226 VTAIL.n225 185
R1598 VTAIL.n247 VTAIL.n246 185
R1599 VTAIL.n250 VTAIL.n249 185
R1600 VTAIL.n248 VTAIL.n222 185
R1601 VTAIL.n255 VTAIL.n221 185
R1602 VTAIL.n257 VTAIL.n256 185
R1603 VTAIL.n259 VTAIL.n258 185
R1604 VTAIL.n218 VTAIL.n217 185
R1605 VTAIL.n265 VTAIL.n264 185
R1606 VTAIL.n267 VTAIL.n266 185
R1607 VTAIL.n214 VTAIL.n213 185
R1608 VTAIL.n273 VTAIL.n272 185
R1609 VTAIL.n275 VTAIL.n274 185
R1610 VTAIL.n210 VTAIL.n209 185
R1611 VTAIL.n281 VTAIL.n280 185
R1612 VTAIL.n283 VTAIL.n282 185
R1613 VTAIL.n206 VTAIL.n205 185
R1614 VTAIL.n289 VTAIL.n288 185
R1615 VTAIL.n291 VTAIL.n290 185
R1616 VTAIL.n202 VTAIL.n201 185
R1617 VTAIL.n297 VTAIL.n296 185
R1618 VTAIL.n697 VTAIL.n696 185
R1619 VTAIL.n602 VTAIL.n601 185
R1620 VTAIL.n691 VTAIL.n690 185
R1621 VTAIL.n689 VTAIL.n688 185
R1622 VTAIL.n606 VTAIL.n605 185
R1623 VTAIL.n683 VTAIL.n682 185
R1624 VTAIL.n681 VTAIL.n680 185
R1625 VTAIL.n610 VTAIL.n609 185
R1626 VTAIL.n675 VTAIL.n674 185
R1627 VTAIL.n673 VTAIL.n672 185
R1628 VTAIL.n614 VTAIL.n613 185
R1629 VTAIL.n667 VTAIL.n666 185
R1630 VTAIL.n665 VTAIL.n664 185
R1631 VTAIL.n618 VTAIL.n617 185
R1632 VTAIL.n659 VTAIL.n658 185
R1633 VTAIL.n657 VTAIL.n656 185
R1634 VTAIL.n655 VTAIL.n621 185
R1635 VTAIL.n625 VTAIL.n622 185
R1636 VTAIL.n650 VTAIL.n649 185
R1637 VTAIL.n648 VTAIL.n647 185
R1638 VTAIL.n627 VTAIL.n626 185
R1639 VTAIL.n642 VTAIL.n641 185
R1640 VTAIL.n640 VTAIL.n639 185
R1641 VTAIL.n631 VTAIL.n630 185
R1642 VTAIL.n634 VTAIL.n633 185
R1643 VTAIL.n597 VTAIL.n596 185
R1644 VTAIL.n502 VTAIL.n501 185
R1645 VTAIL.n591 VTAIL.n590 185
R1646 VTAIL.n589 VTAIL.n588 185
R1647 VTAIL.n506 VTAIL.n505 185
R1648 VTAIL.n583 VTAIL.n582 185
R1649 VTAIL.n581 VTAIL.n580 185
R1650 VTAIL.n510 VTAIL.n509 185
R1651 VTAIL.n575 VTAIL.n574 185
R1652 VTAIL.n573 VTAIL.n572 185
R1653 VTAIL.n514 VTAIL.n513 185
R1654 VTAIL.n567 VTAIL.n566 185
R1655 VTAIL.n565 VTAIL.n564 185
R1656 VTAIL.n518 VTAIL.n517 185
R1657 VTAIL.n559 VTAIL.n558 185
R1658 VTAIL.n557 VTAIL.n556 185
R1659 VTAIL.n555 VTAIL.n521 185
R1660 VTAIL.n525 VTAIL.n522 185
R1661 VTAIL.n550 VTAIL.n549 185
R1662 VTAIL.n548 VTAIL.n547 185
R1663 VTAIL.n527 VTAIL.n526 185
R1664 VTAIL.n542 VTAIL.n541 185
R1665 VTAIL.n540 VTAIL.n539 185
R1666 VTAIL.n531 VTAIL.n530 185
R1667 VTAIL.n534 VTAIL.n533 185
R1668 VTAIL.n497 VTAIL.n496 185
R1669 VTAIL.n402 VTAIL.n401 185
R1670 VTAIL.n491 VTAIL.n490 185
R1671 VTAIL.n489 VTAIL.n488 185
R1672 VTAIL.n406 VTAIL.n405 185
R1673 VTAIL.n483 VTAIL.n482 185
R1674 VTAIL.n481 VTAIL.n480 185
R1675 VTAIL.n410 VTAIL.n409 185
R1676 VTAIL.n475 VTAIL.n474 185
R1677 VTAIL.n473 VTAIL.n472 185
R1678 VTAIL.n414 VTAIL.n413 185
R1679 VTAIL.n467 VTAIL.n466 185
R1680 VTAIL.n465 VTAIL.n464 185
R1681 VTAIL.n418 VTAIL.n417 185
R1682 VTAIL.n459 VTAIL.n458 185
R1683 VTAIL.n457 VTAIL.n456 185
R1684 VTAIL.n455 VTAIL.n421 185
R1685 VTAIL.n425 VTAIL.n422 185
R1686 VTAIL.n450 VTAIL.n449 185
R1687 VTAIL.n448 VTAIL.n447 185
R1688 VTAIL.n427 VTAIL.n426 185
R1689 VTAIL.n442 VTAIL.n441 185
R1690 VTAIL.n440 VTAIL.n439 185
R1691 VTAIL.n431 VTAIL.n430 185
R1692 VTAIL.n434 VTAIL.n433 185
R1693 VTAIL.n397 VTAIL.n396 185
R1694 VTAIL.n302 VTAIL.n301 185
R1695 VTAIL.n391 VTAIL.n390 185
R1696 VTAIL.n389 VTAIL.n388 185
R1697 VTAIL.n306 VTAIL.n305 185
R1698 VTAIL.n383 VTAIL.n382 185
R1699 VTAIL.n381 VTAIL.n380 185
R1700 VTAIL.n310 VTAIL.n309 185
R1701 VTAIL.n375 VTAIL.n374 185
R1702 VTAIL.n373 VTAIL.n372 185
R1703 VTAIL.n314 VTAIL.n313 185
R1704 VTAIL.n367 VTAIL.n366 185
R1705 VTAIL.n365 VTAIL.n364 185
R1706 VTAIL.n318 VTAIL.n317 185
R1707 VTAIL.n359 VTAIL.n358 185
R1708 VTAIL.n357 VTAIL.n356 185
R1709 VTAIL.n355 VTAIL.n321 185
R1710 VTAIL.n325 VTAIL.n322 185
R1711 VTAIL.n350 VTAIL.n349 185
R1712 VTAIL.n348 VTAIL.n347 185
R1713 VTAIL.n327 VTAIL.n326 185
R1714 VTAIL.n342 VTAIL.n341 185
R1715 VTAIL.n340 VTAIL.n339 185
R1716 VTAIL.n331 VTAIL.n330 185
R1717 VTAIL.n334 VTAIL.n333 185
R1718 VTAIL.t5 VTAIL.n731 149.524
R1719 VTAIL.t6 VTAIL.n31 149.524
R1720 VTAIL.t0 VTAIL.n131 149.524
R1721 VTAIL.t3 VTAIL.n231 149.524
R1722 VTAIL.t1 VTAIL.n632 149.524
R1723 VTAIL.t2 VTAIL.n532 149.524
R1724 VTAIL.t4 VTAIL.n432 149.524
R1725 VTAIL.t7 VTAIL.n332 149.524
R1726 VTAIL.n732 VTAIL.n729 104.615
R1727 VTAIL.n739 VTAIL.n729 104.615
R1728 VTAIL.n740 VTAIL.n739 104.615
R1729 VTAIL.n740 VTAIL.n725 104.615
R1730 VTAIL.n747 VTAIL.n725 104.615
R1731 VTAIL.n749 VTAIL.n747 104.615
R1732 VTAIL.n749 VTAIL.n748 104.615
R1733 VTAIL.n748 VTAIL.n721 104.615
R1734 VTAIL.n757 VTAIL.n721 104.615
R1735 VTAIL.n758 VTAIL.n757 104.615
R1736 VTAIL.n758 VTAIL.n717 104.615
R1737 VTAIL.n765 VTAIL.n717 104.615
R1738 VTAIL.n766 VTAIL.n765 104.615
R1739 VTAIL.n766 VTAIL.n713 104.615
R1740 VTAIL.n773 VTAIL.n713 104.615
R1741 VTAIL.n774 VTAIL.n773 104.615
R1742 VTAIL.n774 VTAIL.n709 104.615
R1743 VTAIL.n781 VTAIL.n709 104.615
R1744 VTAIL.n782 VTAIL.n781 104.615
R1745 VTAIL.n782 VTAIL.n705 104.615
R1746 VTAIL.n789 VTAIL.n705 104.615
R1747 VTAIL.n790 VTAIL.n789 104.615
R1748 VTAIL.n790 VTAIL.n701 104.615
R1749 VTAIL.n797 VTAIL.n701 104.615
R1750 VTAIL.n32 VTAIL.n29 104.615
R1751 VTAIL.n39 VTAIL.n29 104.615
R1752 VTAIL.n40 VTAIL.n39 104.615
R1753 VTAIL.n40 VTAIL.n25 104.615
R1754 VTAIL.n47 VTAIL.n25 104.615
R1755 VTAIL.n49 VTAIL.n47 104.615
R1756 VTAIL.n49 VTAIL.n48 104.615
R1757 VTAIL.n48 VTAIL.n21 104.615
R1758 VTAIL.n57 VTAIL.n21 104.615
R1759 VTAIL.n58 VTAIL.n57 104.615
R1760 VTAIL.n58 VTAIL.n17 104.615
R1761 VTAIL.n65 VTAIL.n17 104.615
R1762 VTAIL.n66 VTAIL.n65 104.615
R1763 VTAIL.n66 VTAIL.n13 104.615
R1764 VTAIL.n73 VTAIL.n13 104.615
R1765 VTAIL.n74 VTAIL.n73 104.615
R1766 VTAIL.n74 VTAIL.n9 104.615
R1767 VTAIL.n81 VTAIL.n9 104.615
R1768 VTAIL.n82 VTAIL.n81 104.615
R1769 VTAIL.n82 VTAIL.n5 104.615
R1770 VTAIL.n89 VTAIL.n5 104.615
R1771 VTAIL.n90 VTAIL.n89 104.615
R1772 VTAIL.n90 VTAIL.n1 104.615
R1773 VTAIL.n97 VTAIL.n1 104.615
R1774 VTAIL.n132 VTAIL.n129 104.615
R1775 VTAIL.n139 VTAIL.n129 104.615
R1776 VTAIL.n140 VTAIL.n139 104.615
R1777 VTAIL.n140 VTAIL.n125 104.615
R1778 VTAIL.n147 VTAIL.n125 104.615
R1779 VTAIL.n149 VTAIL.n147 104.615
R1780 VTAIL.n149 VTAIL.n148 104.615
R1781 VTAIL.n148 VTAIL.n121 104.615
R1782 VTAIL.n157 VTAIL.n121 104.615
R1783 VTAIL.n158 VTAIL.n157 104.615
R1784 VTAIL.n158 VTAIL.n117 104.615
R1785 VTAIL.n165 VTAIL.n117 104.615
R1786 VTAIL.n166 VTAIL.n165 104.615
R1787 VTAIL.n166 VTAIL.n113 104.615
R1788 VTAIL.n173 VTAIL.n113 104.615
R1789 VTAIL.n174 VTAIL.n173 104.615
R1790 VTAIL.n174 VTAIL.n109 104.615
R1791 VTAIL.n181 VTAIL.n109 104.615
R1792 VTAIL.n182 VTAIL.n181 104.615
R1793 VTAIL.n182 VTAIL.n105 104.615
R1794 VTAIL.n189 VTAIL.n105 104.615
R1795 VTAIL.n190 VTAIL.n189 104.615
R1796 VTAIL.n190 VTAIL.n101 104.615
R1797 VTAIL.n197 VTAIL.n101 104.615
R1798 VTAIL.n232 VTAIL.n229 104.615
R1799 VTAIL.n239 VTAIL.n229 104.615
R1800 VTAIL.n240 VTAIL.n239 104.615
R1801 VTAIL.n240 VTAIL.n225 104.615
R1802 VTAIL.n247 VTAIL.n225 104.615
R1803 VTAIL.n249 VTAIL.n247 104.615
R1804 VTAIL.n249 VTAIL.n248 104.615
R1805 VTAIL.n248 VTAIL.n221 104.615
R1806 VTAIL.n257 VTAIL.n221 104.615
R1807 VTAIL.n258 VTAIL.n257 104.615
R1808 VTAIL.n258 VTAIL.n217 104.615
R1809 VTAIL.n265 VTAIL.n217 104.615
R1810 VTAIL.n266 VTAIL.n265 104.615
R1811 VTAIL.n266 VTAIL.n213 104.615
R1812 VTAIL.n273 VTAIL.n213 104.615
R1813 VTAIL.n274 VTAIL.n273 104.615
R1814 VTAIL.n274 VTAIL.n209 104.615
R1815 VTAIL.n281 VTAIL.n209 104.615
R1816 VTAIL.n282 VTAIL.n281 104.615
R1817 VTAIL.n282 VTAIL.n205 104.615
R1818 VTAIL.n289 VTAIL.n205 104.615
R1819 VTAIL.n290 VTAIL.n289 104.615
R1820 VTAIL.n290 VTAIL.n201 104.615
R1821 VTAIL.n297 VTAIL.n201 104.615
R1822 VTAIL.n697 VTAIL.n601 104.615
R1823 VTAIL.n690 VTAIL.n601 104.615
R1824 VTAIL.n690 VTAIL.n689 104.615
R1825 VTAIL.n689 VTAIL.n605 104.615
R1826 VTAIL.n682 VTAIL.n605 104.615
R1827 VTAIL.n682 VTAIL.n681 104.615
R1828 VTAIL.n681 VTAIL.n609 104.615
R1829 VTAIL.n674 VTAIL.n609 104.615
R1830 VTAIL.n674 VTAIL.n673 104.615
R1831 VTAIL.n673 VTAIL.n613 104.615
R1832 VTAIL.n666 VTAIL.n613 104.615
R1833 VTAIL.n666 VTAIL.n665 104.615
R1834 VTAIL.n665 VTAIL.n617 104.615
R1835 VTAIL.n658 VTAIL.n617 104.615
R1836 VTAIL.n658 VTAIL.n657 104.615
R1837 VTAIL.n657 VTAIL.n621 104.615
R1838 VTAIL.n625 VTAIL.n621 104.615
R1839 VTAIL.n649 VTAIL.n625 104.615
R1840 VTAIL.n649 VTAIL.n648 104.615
R1841 VTAIL.n648 VTAIL.n626 104.615
R1842 VTAIL.n641 VTAIL.n626 104.615
R1843 VTAIL.n641 VTAIL.n640 104.615
R1844 VTAIL.n640 VTAIL.n630 104.615
R1845 VTAIL.n633 VTAIL.n630 104.615
R1846 VTAIL.n597 VTAIL.n501 104.615
R1847 VTAIL.n590 VTAIL.n501 104.615
R1848 VTAIL.n590 VTAIL.n589 104.615
R1849 VTAIL.n589 VTAIL.n505 104.615
R1850 VTAIL.n582 VTAIL.n505 104.615
R1851 VTAIL.n582 VTAIL.n581 104.615
R1852 VTAIL.n581 VTAIL.n509 104.615
R1853 VTAIL.n574 VTAIL.n509 104.615
R1854 VTAIL.n574 VTAIL.n573 104.615
R1855 VTAIL.n573 VTAIL.n513 104.615
R1856 VTAIL.n566 VTAIL.n513 104.615
R1857 VTAIL.n566 VTAIL.n565 104.615
R1858 VTAIL.n565 VTAIL.n517 104.615
R1859 VTAIL.n558 VTAIL.n517 104.615
R1860 VTAIL.n558 VTAIL.n557 104.615
R1861 VTAIL.n557 VTAIL.n521 104.615
R1862 VTAIL.n525 VTAIL.n521 104.615
R1863 VTAIL.n549 VTAIL.n525 104.615
R1864 VTAIL.n549 VTAIL.n548 104.615
R1865 VTAIL.n548 VTAIL.n526 104.615
R1866 VTAIL.n541 VTAIL.n526 104.615
R1867 VTAIL.n541 VTAIL.n540 104.615
R1868 VTAIL.n540 VTAIL.n530 104.615
R1869 VTAIL.n533 VTAIL.n530 104.615
R1870 VTAIL.n497 VTAIL.n401 104.615
R1871 VTAIL.n490 VTAIL.n401 104.615
R1872 VTAIL.n490 VTAIL.n489 104.615
R1873 VTAIL.n489 VTAIL.n405 104.615
R1874 VTAIL.n482 VTAIL.n405 104.615
R1875 VTAIL.n482 VTAIL.n481 104.615
R1876 VTAIL.n481 VTAIL.n409 104.615
R1877 VTAIL.n474 VTAIL.n409 104.615
R1878 VTAIL.n474 VTAIL.n473 104.615
R1879 VTAIL.n473 VTAIL.n413 104.615
R1880 VTAIL.n466 VTAIL.n413 104.615
R1881 VTAIL.n466 VTAIL.n465 104.615
R1882 VTAIL.n465 VTAIL.n417 104.615
R1883 VTAIL.n458 VTAIL.n417 104.615
R1884 VTAIL.n458 VTAIL.n457 104.615
R1885 VTAIL.n457 VTAIL.n421 104.615
R1886 VTAIL.n425 VTAIL.n421 104.615
R1887 VTAIL.n449 VTAIL.n425 104.615
R1888 VTAIL.n449 VTAIL.n448 104.615
R1889 VTAIL.n448 VTAIL.n426 104.615
R1890 VTAIL.n441 VTAIL.n426 104.615
R1891 VTAIL.n441 VTAIL.n440 104.615
R1892 VTAIL.n440 VTAIL.n430 104.615
R1893 VTAIL.n433 VTAIL.n430 104.615
R1894 VTAIL.n397 VTAIL.n301 104.615
R1895 VTAIL.n390 VTAIL.n301 104.615
R1896 VTAIL.n390 VTAIL.n389 104.615
R1897 VTAIL.n389 VTAIL.n305 104.615
R1898 VTAIL.n382 VTAIL.n305 104.615
R1899 VTAIL.n382 VTAIL.n381 104.615
R1900 VTAIL.n381 VTAIL.n309 104.615
R1901 VTAIL.n374 VTAIL.n309 104.615
R1902 VTAIL.n374 VTAIL.n373 104.615
R1903 VTAIL.n373 VTAIL.n313 104.615
R1904 VTAIL.n366 VTAIL.n313 104.615
R1905 VTAIL.n366 VTAIL.n365 104.615
R1906 VTAIL.n365 VTAIL.n317 104.615
R1907 VTAIL.n358 VTAIL.n317 104.615
R1908 VTAIL.n358 VTAIL.n357 104.615
R1909 VTAIL.n357 VTAIL.n321 104.615
R1910 VTAIL.n325 VTAIL.n321 104.615
R1911 VTAIL.n349 VTAIL.n325 104.615
R1912 VTAIL.n349 VTAIL.n348 104.615
R1913 VTAIL.n348 VTAIL.n326 104.615
R1914 VTAIL.n341 VTAIL.n326 104.615
R1915 VTAIL.n341 VTAIL.n340 104.615
R1916 VTAIL.n340 VTAIL.n330 104.615
R1917 VTAIL.n333 VTAIL.n330 104.615
R1918 VTAIL.n732 VTAIL.t5 52.3082
R1919 VTAIL.n32 VTAIL.t6 52.3082
R1920 VTAIL.n132 VTAIL.t0 52.3082
R1921 VTAIL.n232 VTAIL.t3 52.3082
R1922 VTAIL.n633 VTAIL.t1 52.3082
R1923 VTAIL.n533 VTAIL.t2 52.3082
R1924 VTAIL.n433 VTAIL.t4 52.3082
R1925 VTAIL.n333 VTAIL.t7 52.3082
R1926 VTAIL.n799 VTAIL.n798 34.5126
R1927 VTAIL.n99 VTAIL.n98 34.5126
R1928 VTAIL.n199 VTAIL.n198 34.5126
R1929 VTAIL.n299 VTAIL.n298 34.5126
R1930 VTAIL.n699 VTAIL.n698 34.5126
R1931 VTAIL.n599 VTAIL.n598 34.5126
R1932 VTAIL.n499 VTAIL.n498 34.5126
R1933 VTAIL.n399 VTAIL.n398 34.5126
R1934 VTAIL.n799 VTAIL.n699 29.5048
R1935 VTAIL.n399 VTAIL.n299 29.5048
R1936 VTAIL.n756 VTAIL.n755 13.1884
R1937 VTAIL.n56 VTAIL.n55 13.1884
R1938 VTAIL.n156 VTAIL.n155 13.1884
R1939 VTAIL.n256 VTAIL.n255 13.1884
R1940 VTAIL.n656 VTAIL.n655 13.1884
R1941 VTAIL.n556 VTAIL.n555 13.1884
R1942 VTAIL.n456 VTAIL.n455 13.1884
R1943 VTAIL.n356 VTAIL.n355 13.1884
R1944 VTAIL.n754 VTAIL.n722 12.8005
R1945 VTAIL.n759 VTAIL.n720 12.8005
R1946 VTAIL.n54 VTAIL.n22 12.8005
R1947 VTAIL.n59 VTAIL.n20 12.8005
R1948 VTAIL.n154 VTAIL.n122 12.8005
R1949 VTAIL.n159 VTAIL.n120 12.8005
R1950 VTAIL.n254 VTAIL.n222 12.8005
R1951 VTAIL.n259 VTAIL.n220 12.8005
R1952 VTAIL.n659 VTAIL.n620 12.8005
R1953 VTAIL.n654 VTAIL.n622 12.8005
R1954 VTAIL.n559 VTAIL.n520 12.8005
R1955 VTAIL.n554 VTAIL.n522 12.8005
R1956 VTAIL.n459 VTAIL.n420 12.8005
R1957 VTAIL.n454 VTAIL.n422 12.8005
R1958 VTAIL.n359 VTAIL.n320 12.8005
R1959 VTAIL.n354 VTAIL.n322 12.8005
R1960 VTAIL.n751 VTAIL.n750 12.0247
R1961 VTAIL.n760 VTAIL.n718 12.0247
R1962 VTAIL.n796 VTAIL.n700 12.0247
R1963 VTAIL.n51 VTAIL.n50 12.0247
R1964 VTAIL.n60 VTAIL.n18 12.0247
R1965 VTAIL.n96 VTAIL.n0 12.0247
R1966 VTAIL.n151 VTAIL.n150 12.0247
R1967 VTAIL.n160 VTAIL.n118 12.0247
R1968 VTAIL.n196 VTAIL.n100 12.0247
R1969 VTAIL.n251 VTAIL.n250 12.0247
R1970 VTAIL.n260 VTAIL.n218 12.0247
R1971 VTAIL.n296 VTAIL.n200 12.0247
R1972 VTAIL.n696 VTAIL.n600 12.0247
R1973 VTAIL.n660 VTAIL.n618 12.0247
R1974 VTAIL.n651 VTAIL.n650 12.0247
R1975 VTAIL.n596 VTAIL.n500 12.0247
R1976 VTAIL.n560 VTAIL.n518 12.0247
R1977 VTAIL.n551 VTAIL.n550 12.0247
R1978 VTAIL.n496 VTAIL.n400 12.0247
R1979 VTAIL.n460 VTAIL.n418 12.0247
R1980 VTAIL.n451 VTAIL.n450 12.0247
R1981 VTAIL.n396 VTAIL.n300 12.0247
R1982 VTAIL.n360 VTAIL.n318 12.0247
R1983 VTAIL.n351 VTAIL.n350 12.0247
R1984 VTAIL.n746 VTAIL.n724 11.249
R1985 VTAIL.n764 VTAIL.n763 11.249
R1986 VTAIL.n795 VTAIL.n702 11.249
R1987 VTAIL.n46 VTAIL.n24 11.249
R1988 VTAIL.n64 VTAIL.n63 11.249
R1989 VTAIL.n95 VTAIL.n2 11.249
R1990 VTAIL.n146 VTAIL.n124 11.249
R1991 VTAIL.n164 VTAIL.n163 11.249
R1992 VTAIL.n195 VTAIL.n102 11.249
R1993 VTAIL.n246 VTAIL.n224 11.249
R1994 VTAIL.n264 VTAIL.n263 11.249
R1995 VTAIL.n295 VTAIL.n202 11.249
R1996 VTAIL.n695 VTAIL.n602 11.249
R1997 VTAIL.n664 VTAIL.n663 11.249
R1998 VTAIL.n647 VTAIL.n624 11.249
R1999 VTAIL.n595 VTAIL.n502 11.249
R2000 VTAIL.n564 VTAIL.n563 11.249
R2001 VTAIL.n547 VTAIL.n524 11.249
R2002 VTAIL.n495 VTAIL.n402 11.249
R2003 VTAIL.n464 VTAIL.n463 11.249
R2004 VTAIL.n447 VTAIL.n424 11.249
R2005 VTAIL.n395 VTAIL.n302 11.249
R2006 VTAIL.n364 VTAIL.n363 11.249
R2007 VTAIL.n347 VTAIL.n324 11.249
R2008 VTAIL.n745 VTAIL.n726 10.4732
R2009 VTAIL.n767 VTAIL.n716 10.4732
R2010 VTAIL.n792 VTAIL.n791 10.4732
R2011 VTAIL.n45 VTAIL.n26 10.4732
R2012 VTAIL.n67 VTAIL.n16 10.4732
R2013 VTAIL.n92 VTAIL.n91 10.4732
R2014 VTAIL.n145 VTAIL.n126 10.4732
R2015 VTAIL.n167 VTAIL.n116 10.4732
R2016 VTAIL.n192 VTAIL.n191 10.4732
R2017 VTAIL.n245 VTAIL.n226 10.4732
R2018 VTAIL.n267 VTAIL.n216 10.4732
R2019 VTAIL.n292 VTAIL.n291 10.4732
R2020 VTAIL.n692 VTAIL.n691 10.4732
R2021 VTAIL.n667 VTAIL.n616 10.4732
R2022 VTAIL.n646 VTAIL.n627 10.4732
R2023 VTAIL.n592 VTAIL.n591 10.4732
R2024 VTAIL.n567 VTAIL.n516 10.4732
R2025 VTAIL.n546 VTAIL.n527 10.4732
R2026 VTAIL.n492 VTAIL.n491 10.4732
R2027 VTAIL.n467 VTAIL.n416 10.4732
R2028 VTAIL.n446 VTAIL.n427 10.4732
R2029 VTAIL.n392 VTAIL.n391 10.4732
R2030 VTAIL.n367 VTAIL.n316 10.4732
R2031 VTAIL.n346 VTAIL.n327 10.4732
R2032 VTAIL.n733 VTAIL.n731 10.2747
R2033 VTAIL.n33 VTAIL.n31 10.2747
R2034 VTAIL.n133 VTAIL.n131 10.2747
R2035 VTAIL.n233 VTAIL.n231 10.2747
R2036 VTAIL.n634 VTAIL.n632 10.2747
R2037 VTAIL.n534 VTAIL.n532 10.2747
R2038 VTAIL.n434 VTAIL.n432 10.2747
R2039 VTAIL.n334 VTAIL.n332 10.2747
R2040 VTAIL.n742 VTAIL.n741 9.69747
R2041 VTAIL.n768 VTAIL.n714 9.69747
R2042 VTAIL.n788 VTAIL.n704 9.69747
R2043 VTAIL.n42 VTAIL.n41 9.69747
R2044 VTAIL.n68 VTAIL.n14 9.69747
R2045 VTAIL.n88 VTAIL.n4 9.69747
R2046 VTAIL.n142 VTAIL.n141 9.69747
R2047 VTAIL.n168 VTAIL.n114 9.69747
R2048 VTAIL.n188 VTAIL.n104 9.69747
R2049 VTAIL.n242 VTAIL.n241 9.69747
R2050 VTAIL.n268 VTAIL.n214 9.69747
R2051 VTAIL.n288 VTAIL.n204 9.69747
R2052 VTAIL.n688 VTAIL.n604 9.69747
R2053 VTAIL.n668 VTAIL.n614 9.69747
R2054 VTAIL.n643 VTAIL.n642 9.69747
R2055 VTAIL.n588 VTAIL.n504 9.69747
R2056 VTAIL.n568 VTAIL.n514 9.69747
R2057 VTAIL.n543 VTAIL.n542 9.69747
R2058 VTAIL.n488 VTAIL.n404 9.69747
R2059 VTAIL.n468 VTAIL.n414 9.69747
R2060 VTAIL.n443 VTAIL.n442 9.69747
R2061 VTAIL.n388 VTAIL.n304 9.69747
R2062 VTAIL.n368 VTAIL.n314 9.69747
R2063 VTAIL.n343 VTAIL.n342 9.69747
R2064 VTAIL.n794 VTAIL.n700 9.45567
R2065 VTAIL.n94 VTAIL.n0 9.45567
R2066 VTAIL.n194 VTAIL.n100 9.45567
R2067 VTAIL.n294 VTAIL.n200 9.45567
R2068 VTAIL.n694 VTAIL.n600 9.45567
R2069 VTAIL.n594 VTAIL.n500 9.45567
R2070 VTAIL.n494 VTAIL.n400 9.45567
R2071 VTAIL.n394 VTAIL.n300 9.45567
R2072 VTAIL.n779 VTAIL.n778 9.3005
R2073 VTAIL.n708 VTAIL.n707 9.3005
R2074 VTAIL.n785 VTAIL.n784 9.3005
R2075 VTAIL.n787 VTAIL.n786 9.3005
R2076 VTAIL.n704 VTAIL.n703 9.3005
R2077 VTAIL.n793 VTAIL.n792 9.3005
R2078 VTAIL.n795 VTAIL.n794 9.3005
R2079 VTAIL.n712 VTAIL.n711 9.3005
R2080 VTAIL.n771 VTAIL.n770 9.3005
R2081 VTAIL.n769 VTAIL.n768 9.3005
R2082 VTAIL.n716 VTAIL.n715 9.3005
R2083 VTAIL.n763 VTAIL.n762 9.3005
R2084 VTAIL.n761 VTAIL.n760 9.3005
R2085 VTAIL.n720 VTAIL.n719 9.3005
R2086 VTAIL.n735 VTAIL.n734 9.3005
R2087 VTAIL.n737 VTAIL.n736 9.3005
R2088 VTAIL.n728 VTAIL.n727 9.3005
R2089 VTAIL.n743 VTAIL.n742 9.3005
R2090 VTAIL.n745 VTAIL.n744 9.3005
R2091 VTAIL.n724 VTAIL.n723 9.3005
R2092 VTAIL.n752 VTAIL.n751 9.3005
R2093 VTAIL.n754 VTAIL.n753 9.3005
R2094 VTAIL.n777 VTAIL.n776 9.3005
R2095 VTAIL.n79 VTAIL.n78 9.3005
R2096 VTAIL.n8 VTAIL.n7 9.3005
R2097 VTAIL.n85 VTAIL.n84 9.3005
R2098 VTAIL.n87 VTAIL.n86 9.3005
R2099 VTAIL.n4 VTAIL.n3 9.3005
R2100 VTAIL.n93 VTAIL.n92 9.3005
R2101 VTAIL.n95 VTAIL.n94 9.3005
R2102 VTAIL.n12 VTAIL.n11 9.3005
R2103 VTAIL.n71 VTAIL.n70 9.3005
R2104 VTAIL.n69 VTAIL.n68 9.3005
R2105 VTAIL.n16 VTAIL.n15 9.3005
R2106 VTAIL.n63 VTAIL.n62 9.3005
R2107 VTAIL.n61 VTAIL.n60 9.3005
R2108 VTAIL.n20 VTAIL.n19 9.3005
R2109 VTAIL.n35 VTAIL.n34 9.3005
R2110 VTAIL.n37 VTAIL.n36 9.3005
R2111 VTAIL.n28 VTAIL.n27 9.3005
R2112 VTAIL.n43 VTAIL.n42 9.3005
R2113 VTAIL.n45 VTAIL.n44 9.3005
R2114 VTAIL.n24 VTAIL.n23 9.3005
R2115 VTAIL.n52 VTAIL.n51 9.3005
R2116 VTAIL.n54 VTAIL.n53 9.3005
R2117 VTAIL.n77 VTAIL.n76 9.3005
R2118 VTAIL.n179 VTAIL.n178 9.3005
R2119 VTAIL.n108 VTAIL.n107 9.3005
R2120 VTAIL.n185 VTAIL.n184 9.3005
R2121 VTAIL.n187 VTAIL.n186 9.3005
R2122 VTAIL.n104 VTAIL.n103 9.3005
R2123 VTAIL.n193 VTAIL.n192 9.3005
R2124 VTAIL.n195 VTAIL.n194 9.3005
R2125 VTAIL.n112 VTAIL.n111 9.3005
R2126 VTAIL.n171 VTAIL.n170 9.3005
R2127 VTAIL.n169 VTAIL.n168 9.3005
R2128 VTAIL.n116 VTAIL.n115 9.3005
R2129 VTAIL.n163 VTAIL.n162 9.3005
R2130 VTAIL.n161 VTAIL.n160 9.3005
R2131 VTAIL.n120 VTAIL.n119 9.3005
R2132 VTAIL.n135 VTAIL.n134 9.3005
R2133 VTAIL.n137 VTAIL.n136 9.3005
R2134 VTAIL.n128 VTAIL.n127 9.3005
R2135 VTAIL.n143 VTAIL.n142 9.3005
R2136 VTAIL.n145 VTAIL.n144 9.3005
R2137 VTAIL.n124 VTAIL.n123 9.3005
R2138 VTAIL.n152 VTAIL.n151 9.3005
R2139 VTAIL.n154 VTAIL.n153 9.3005
R2140 VTAIL.n177 VTAIL.n176 9.3005
R2141 VTAIL.n279 VTAIL.n278 9.3005
R2142 VTAIL.n208 VTAIL.n207 9.3005
R2143 VTAIL.n285 VTAIL.n284 9.3005
R2144 VTAIL.n287 VTAIL.n286 9.3005
R2145 VTAIL.n204 VTAIL.n203 9.3005
R2146 VTAIL.n293 VTAIL.n292 9.3005
R2147 VTAIL.n295 VTAIL.n294 9.3005
R2148 VTAIL.n212 VTAIL.n211 9.3005
R2149 VTAIL.n271 VTAIL.n270 9.3005
R2150 VTAIL.n269 VTAIL.n268 9.3005
R2151 VTAIL.n216 VTAIL.n215 9.3005
R2152 VTAIL.n263 VTAIL.n262 9.3005
R2153 VTAIL.n261 VTAIL.n260 9.3005
R2154 VTAIL.n220 VTAIL.n219 9.3005
R2155 VTAIL.n235 VTAIL.n234 9.3005
R2156 VTAIL.n237 VTAIL.n236 9.3005
R2157 VTAIL.n228 VTAIL.n227 9.3005
R2158 VTAIL.n243 VTAIL.n242 9.3005
R2159 VTAIL.n245 VTAIL.n244 9.3005
R2160 VTAIL.n224 VTAIL.n223 9.3005
R2161 VTAIL.n252 VTAIL.n251 9.3005
R2162 VTAIL.n254 VTAIL.n253 9.3005
R2163 VTAIL.n277 VTAIL.n276 9.3005
R2164 VTAIL.n695 VTAIL.n694 9.3005
R2165 VTAIL.n693 VTAIL.n692 9.3005
R2166 VTAIL.n604 VTAIL.n603 9.3005
R2167 VTAIL.n687 VTAIL.n686 9.3005
R2168 VTAIL.n685 VTAIL.n684 9.3005
R2169 VTAIL.n608 VTAIL.n607 9.3005
R2170 VTAIL.n679 VTAIL.n678 9.3005
R2171 VTAIL.n677 VTAIL.n676 9.3005
R2172 VTAIL.n612 VTAIL.n611 9.3005
R2173 VTAIL.n671 VTAIL.n670 9.3005
R2174 VTAIL.n669 VTAIL.n668 9.3005
R2175 VTAIL.n616 VTAIL.n615 9.3005
R2176 VTAIL.n663 VTAIL.n662 9.3005
R2177 VTAIL.n661 VTAIL.n660 9.3005
R2178 VTAIL.n620 VTAIL.n619 9.3005
R2179 VTAIL.n654 VTAIL.n653 9.3005
R2180 VTAIL.n652 VTAIL.n651 9.3005
R2181 VTAIL.n624 VTAIL.n623 9.3005
R2182 VTAIL.n646 VTAIL.n645 9.3005
R2183 VTAIL.n644 VTAIL.n643 9.3005
R2184 VTAIL.n629 VTAIL.n628 9.3005
R2185 VTAIL.n638 VTAIL.n637 9.3005
R2186 VTAIL.n636 VTAIL.n635 9.3005
R2187 VTAIL.n536 VTAIL.n535 9.3005
R2188 VTAIL.n538 VTAIL.n537 9.3005
R2189 VTAIL.n529 VTAIL.n528 9.3005
R2190 VTAIL.n544 VTAIL.n543 9.3005
R2191 VTAIL.n546 VTAIL.n545 9.3005
R2192 VTAIL.n524 VTAIL.n523 9.3005
R2193 VTAIL.n552 VTAIL.n551 9.3005
R2194 VTAIL.n554 VTAIL.n553 9.3005
R2195 VTAIL.n508 VTAIL.n507 9.3005
R2196 VTAIL.n585 VTAIL.n584 9.3005
R2197 VTAIL.n587 VTAIL.n586 9.3005
R2198 VTAIL.n504 VTAIL.n503 9.3005
R2199 VTAIL.n593 VTAIL.n592 9.3005
R2200 VTAIL.n595 VTAIL.n594 9.3005
R2201 VTAIL.n579 VTAIL.n578 9.3005
R2202 VTAIL.n577 VTAIL.n576 9.3005
R2203 VTAIL.n512 VTAIL.n511 9.3005
R2204 VTAIL.n571 VTAIL.n570 9.3005
R2205 VTAIL.n569 VTAIL.n568 9.3005
R2206 VTAIL.n516 VTAIL.n515 9.3005
R2207 VTAIL.n563 VTAIL.n562 9.3005
R2208 VTAIL.n561 VTAIL.n560 9.3005
R2209 VTAIL.n520 VTAIL.n519 9.3005
R2210 VTAIL.n436 VTAIL.n435 9.3005
R2211 VTAIL.n438 VTAIL.n437 9.3005
R2212 VTAIL.n429 VTAIL.n428 9.3005
R2213 VTAIL.n444 VTAIL.n443 9.3005
R2214 VTAIL.n446 VTAIL.n445 9.3005
R2215 VTAIL.n424 VTAIL.n423 9.3005
R2216 VTAIL.n452 VTAIL.n451 9.3005
R2217 VTAIL.n454 VTAIL.n453 9.3005
R2218 VTAIL.n408 VTAIL.n407 9.3005
R2219 VTAIL.n485 VTAIL.n484 9.3005
R2220 VTAIL.n487 VTAIL.n486 9.3005
R2221 VTAIL.n404 VTAIL.n403 9.3005
R2222 VTAIL.n493 VTAIL.n492 9.3005
R2223 VTAIL.n495 VTAIL.n494 9.3005
R2224 VTAIL.n479 VTAIL.n478 9.3005
R2225 VTAIL.n477 VTAIL.n476 9.3005
R2226 VTAIL.n412 VTAIL.n411 9.3005
R2227 VTAIL.n471 VTAIL.n470 9.3005
R2228 VTAIL.n469 VTAIL.n468 9.3005
R2229 VTAIL.n416 VTAIL.n415 9.3005
R2230 VTAIL.n463 VTAIL.n462 9.3005
R2231 VTAIL.n461 VTAIL.n460 9.3005
R2232 VTAIL.n420 VTAIL.n419 9.3005
R2233 VTAIL.n336 VTAIL.n335 9.3005
R2234 VTAIL.n338 VTAIL.n337 9.3005
R2235 VTAIL.n329 VTAIL.n328 9.3005
R2236 VTAIL.n344 VTAIL.n343 9.3005
R2237 VTAIL.n346 VTAIL.n345 9.3005
R2238 VTAIL.n324 VTAIL.n323 9.3005
R2239 VTAIL.n352 VTAIL.n351 9.3005
R2240 VTAIL.n354 VTAIL.n353 9.3005
R2241 VTAIL.n308 VTAIL.n307 9.3005
R2242 VTAIL.n385 VTAIL.n384 9.3005
R2243 VTAIL.n387 VTAIL.n386 9.3005
R2244 VTAIL.n304 VTAIL.n303 9.3005
R2245 VTAIL.n393 VTAIL.n392 9.3005
R2246 VTAIL.n395 VTAIL.n394 9.3005
R2247 VTAIL.n379 VTAIL.n378 9.3005
R2248 VTAIL.n377 VTAIL.n376 9.3005
R2249 VTAIL.n312 VTAIL.n311 9.3005
R2250 VTAIL.n371 VTAIL.n370 9.3005
R2251 VTAIL.n369 VTAIL.n368 9.3005
R2252 VTAIL.n316 VTAIL.n315 9.3005
R2253 VTAIL.n363 VTAIL.n362 9.3005
R2254 VTAIL.n361 VTAIL.n360 9.3005
R2255 VTAIL.n320 VTAIL.n319 9.3005
R2256 VTAIL.n738 VTAIL.n728 8.92171
R2257 VTAIL.n772 VTAIL.n771 8.92171
R2258 VTAIL.n787 VTAIL.n706 8.92171
R2259 VTAIL.n38 VTAIL.n28 8.92171
R2260 VTAIL.n72 VTAIL.n71 8.92171
R2261 VTAIL.n87 VTAIL.n6 8.92171
R2262 VTAIL.n138 VTAIL.n128 8.92171
R2263 VTAIL.n172 VTAIL.n171 8.92171
R2264 VTAIL.n187 VTAIL.n106 8.92171
R2265 VTAIL.n238 VTAIL.n228 8.92171
R2266 VTAIL.n272 VTAIL.n271 8.92171
R2267 VTAIL.n287 VTAIL.n206 8.92171
R2268 VTAIL.n687 VTAIL.n606 8.92171
R2269 VTAIL.n672 VTAIL.n671 8.92171
R2270 VTAIL.n639 VTAIL.n629 8.92171
R2271 VTAIL.n587 VTAIL.n506 8.92171
R2272 VTAIL.n572 VTAIL.n571 8.92171
R2273 VTAIL.n539 VTAIL.n529 8.92171
R2274 VTAIL.n487 VTAIL.n406 8.92171
R2275 VTAIL.n472 VTAIL.n471 8.92171
R2276 VTAIL.n439 VTAIL.n429 8.92171
R2277 VTAIL.n387 VTAIL.n306 8.92171
R2278 VTAIL.n372 VTAIL.n371 8.92171
R2279 VTAIL.n339 VTAIL.n329 8.92171
R2280 VTAIL.n737 VTAIL.n730 8.14595
R2281 VTAIL.n775 VTAIL.n712 8.14595
R2282 VTAIL.n784 VTAIL.n783 8.14595
R2283 VTAIL.n37 VTAIL.n30 8.14595
R2284 VTAIL.n75 VTAIL.n12 8.14595
R2285 VTAIL.n84 VTAIL.n83 8.14595
R2286 VTAIL.n137 VTAIL.n130 8.14595
R2287 VTAIL.n175 VTAIL.n112 8.14595
R2288 VTAIL.n184 VTAIL.n183 8.14595
R2289 VTAIL.n237 VTAIL.n230 8.14595
R2290 VTAIL.n275 VTAIL.n212 8.14595
R2291 VTAIL.n284 VTAIL.n283 8.14595
R2292 VTAIL.n684 VTAIL.n683 8.14595
R2293 VTAIL.n675 VTAIL.n612 8.14595
R2294 VTAIL.n638 VTAIL.n631 8.14595
R2295 VTAIL.n584 VTAIL.n583 8.14595
R2296 VTAIL.n575 VTAIL.n512 8.14595
R2297 VTAIL.n538 VTAIL.n531 8.14595
R2298 VTAIL.n484 VTAIL.n483 8.14595
R2299 VTAIL.n475 VTAIL.n412 8.14595
R2300 VTAIL.n438 VTAIL.n431 8.14595
R2301 VTAIL.n384 VTAIL.n383 8.14595
R2302 VTAIL.n375 VTAIL.n312 8.14595
R2303 VTAIL.n338 VTAIL.n331 8.14595
R2304 VTAIL.n734 VTAIL.n733 7.3702
R2305 VTAIL.n776 VTAIL.n710 7.3702
R2306 VTAIL.n780 VTAIL.n708 7.3702
R2307 VTAIL.n34 VTAIL.n33 7.3702
R2308 VTAIL.n76 VTAIL.n10 7.3702
R2309 VTAIL.n80 VTAIL.n8 7.3702
R2310 VTAIL.n134 VTAIL.n133 7.3702
R2311 VTAIL.n176 VTAIL.n110 7.3702
R2312 VTAIL.n180 VTAIL.n108 7.3702
R2313 VTAIL.n234 VTAIL.n233 7.3702
R2314 VTAIL.n276 VTAIL.n210 7.3702
R2315 VTAIL.n280 VTAIL.n208 7.3702
R2316 VTAIL.n680 VTAIL.n608 7.3702
R2317 VTAIL.n676 VTAIL.n610 7.3702
R2318 VTAIL.n635 VTAIL.n634 7.3702
R2319 VTAIL.n580 VTAIL.n508 7.3702
R2320 VTAIL.n576 VTAIL.n510 7.3702
R2321 VTAIL.n535 VTAIL.n534 7.3702
R2322 VTAIL.n480 VTAIL.n408 7.3702
R2323 VTAIL.n476 VTAIL.n410 7.3702
R2324 VTAIL.n435 VTAIL.n434 7.3702
R2325 VTAIL.n380 VTAIL.n308 7.3702
R2326 VTAIL.n376 VTAIL.n310 7.3702
R2327 VTAIL.n335 VTAIL.n334 7.3702
R2328 VTAIL.n779 VTAIL.n710 6.59444
R2329 VTAIL.n780 VTAIL.n779 6.59444
R2330 VTAIL.n79 VTAIL.n10 6.59444
R2331 VTAIL.n80 VTAIL.n79 6.59444
R2332 VTAIL.n179 VTAIL.n110 6.59444
R2333 VTAIL.n180 VTAIL.n179 6.59444
R2334 VTAIL.n279 VTAIL.n210 6.59444
R2335 VTAIL.n280 VTAIL.n279 6.59444
R2336 VTAIL.n680 VTAIL.n679 6.59444
R2337 VTAIL.n679 VTAIL.n610 6.59444
R2338 VTAIL.n580 VTAIL.n579 6.59444
R2339 VTAIL.n579 VTAIL.n510 6.59444
R2340 VTAIL.n480 VTAIL.n479 6.59444
R2341 VTAIL.n479 VTAIL.n410 6.59444
R2342 VTAIL.n380 VTAIL.n379 6.59444
R2343 VTAIL.n379 VTAIL.n310 6.59444
R2344 VTAIL.n734 VTAIL.n730 5.81868
R2345 VTAIL.n776 VTAIL.n775 5.81868
R2346 VTAIL.n783 VTAIL.n708 5.81868
R2347 VTAIL.n34 VTAIL.n30 5.81868
R2348 VTAIL.n76 VTAIL.n75 5.81868
R2349 VTAIL.n83 VTAIL.n8 5.81868
R2350 VTAIL.n134 VTAIL.n130 5.81868
R2351 VTAIL.n176 VTAIL.n175 5.81868
R2352 VTAIL.n183 VTAIL.n108 5.81868
R2353 VTAIL.n234 VTAIL.n230 5.81868
R2354 VTAIL.n276 VTAIL.n275 5.81868
R2355 VTAIL.n283 VTAIL.n208 5.81868
R2356 VTAIL.n683 VTAIL.n608 5.81868
R2357 VTAIL.n676 VTAIL.n675 5.81868
R2358 VTAIL.n635 VTAIL.n631 5.81868
R2359 VTAIL.n583 VTAIL.n508 5.81868
R2360 VTAIL.n576 VTAIL.n575 5.81868
R2361 VTAIL.n535 VTAIL.n531 5.81868
R2362 VTAIL.n483 VTAIL.n408 5.81868
R2363 VTAIL.n476 VTAIL.n475 5.81868
R2364 VTAIL.n435 VTAIL.n431 5.81868
R2365 VTAIL.n383 VTAIL.n308 5.81868
R2366 VTAIL.n376 VTAIL.n375 5.81868
R2367 VTAIL.n335 VTAIL.n331 5.81868
R2368 VTAIL.n738 VTAIL.n737 5.04292
R2369 VTAIL.n772 VTAIL.n712 5.04292
R2370 VTAIL.n784 VTAIL.n706 5.04292
R2371 VTAIL.n38 VTAIL.n37 5.04292
R2372 VTAIL.n72 VTAIL.n12 5.04292
R2373 VTAIL.n84 VTAIL.n6 5.04292
R2374 VTAIL.n138 VTAIL.n137 5.04292
R2375 VTAIL.n172 VTAIL.n112 5.04292
R2376 VTAIL.n184 VTAIL.n106 5.04292
R2377 VTAIL.n238 VTAIL.n237 5.04292
R2378 VTAIL.n272 VTAIL.n212 5.04292
R2379 VTAIL.n284 VTAIL.n206 5.04292
R2380 VTAIL.n684 VTAIL.n606 5.04292
R2381 VTAIL.n672 VTAIL.n612 5.04292
R2382 VTAIL.n639 VTAIL.n638 5.04292
R2383 VTAIL.n584 VTAIL.n506 5.04292
R2384 VTAIL.n572 VTAIL.n512 5.04292
R2385 VTAIL.n539 VTAIL.n538 5.04292
R2386 VTAIL.n484 VTAIL.n406 5.04292
R2387 VTAIL.n472 VTAIL.n412 5.04292
R2388 VTAIL.n439 VTAIL.n438 5.04292
R2389 VTAIL.n384 VTAIL.n306 5.04292
R2390 VTAIL.n372 VTAIL.n312 5.04292
R2391 VTAIL.n339 VTAIL.n338 5.04292
R2392 VTAIL.n741 VTAIL.n728 4.26717
R2393 VTAIL.n771 VTAIL.n714 4.26717
R2394 VTAIL.n788 VTAIL.n787 4.26717
R2395 VTAIL.n41 VTAIL.n28 4.26717
R2396 VTAIL.n71 VTAIL.n14 4.26717
R2397 VTAIL.n88 VTAIL.n87 4.26717
R2398 VTAIL.n141 VTAIL.n128 4.26717
R2399 VTAIL.n171 VTAIL.n114 4.26717
R2400 VTAIL.n188 VTAIL.n187 4.26717
R2401 VTAIL.n241 VTAIL.n228 4.26717
R2402 VTAIL.n271 VTAIL.n214 4.26717
R2403 VTAIL.n288 VTAIL.n287 4.26717
R2404 VTAIL.n688 VTAIL.n687 4.26717
R2405 VTAIL.n671 VTAIL.n614 4.26717
R2406 VTAIL.n642 VTAIL.n629 4.26717
R2407 VTAIL.n588 VTAIL.n587 4.26717
R2408 VTAIL.n571 VTAIL.n514 4.26717
R2409 VTAIL.n542 VTAIL.n529 4.26717
R2410 VTAIL.n488 VTAIL.n487 4.26717
R2411 VTAIL.n471 VTAIL.n414 4.26717
R2412 VTAIL.n442 VTAIL.n429 4.26717
R2413 VTAIL.n388 VTAIL.n387 4.26717
R2414 VTAIL.n371 VTAIL.n314 4.26717
R2415 VTAIL.n342 VTAIL.n329 4.26717
R2416 VTAIL.n742 VTAIL.n726 3.49141
R2417 VTAIL.n768 VTAIL.n767 3.49141
R2418 VTAIL.n791 VTAIL.n704 3.49141
R2419 VTAIL.n42 VTAIL.n26 3.49141
R2420 VTAIL.n68 VTAIL.n67 3.49141
R2421 VTAIL.n91 VTAIL.n4 3.49141
R2422 VTAIL.n142 VTAIL.n126 3.49141
R2423 VTAIL.n168 VTAIL.n167 3.49141
R2424 VTAIL.n191 VTAIL.n104 3.49141
R2425 VTAIL.n242 VTAIL.n226 3.49141
R2426 VTAIL.n268 VTAIL.n267 3.49141
R2427 VTAIL.n291 VTAIL.n204 3.49141
R2428 VTAIL.n691 VTAIL.n604 3.49141
R2429 VTAIL.n668 VTAIL.n667 3.49141
R2430 VTAIL.n643 VTAIL.n627 3.49141
R2431 VTAIL.n591 VTAIL.n504 3.49141
R2432 VTAIL.n568 VTAIL.n567 3.49141
R2433 VTAIL.n543 VTAIL.n527 3.49141
R2434 VTAIL.n491 VTAIL.n404 3.49141
R2435 VTAIL.n468 VTAIL.n467 3.49141
R2436 VTAIL.n443 VTAIL.n427 3.49141
R2437 VTAIL.n391 VTAIL.n304 3.49141
R2438 VTAIL.n368 VTAIL.n367 3.49141
R2439 VTAIL.n343 VTAIL.n327 3.49141
R2440 VTAIL.n536 VTAIL.n532 2.84303
R2441 VTAIL.n436 VTAIL.n432 2.84303
R2442 VTAIL.n336 VTAIL.n332 2.84303
R2443 VTAIL.n735 VTAIL.n731 2.84303
R2444 VTAIL.n35 VTAIL.n31 2.84303
R2445 VTAIL.n135 VTAIL.n131 2.84303
R2446 VTAIL.n235 VTAIL.n231 2.84303
R2447 VTAIL.n636 VTAIL.n632 2.84303
R2448 VTAIL.n746 VTAIL.n745 2.71565
R2449 VTAIL.n764 VTAIL.n716 2.71565
R2450 VTAIL.n792 VTAIL.n702 2.71565
R2451 VTAIL.n46 VTAIL.n45 2.71565
R2452 VTAIL.n64 VTAIL.n16 2.71565
R2453 VTAIL.n92 VTAIL.n2 2.71565
R2454 VTAIL.n146 VTAIL.n145 2.71565
R2455 VTAIL.n164 VTAIL.n116 2.71565
R2456 VTAIL.n192 VTAIL.n102 2.71565
R2457 VTAIL.n246 VTAIL.n245 2.71565
R2458 VTAIL.n264 VTAIL.n216 2.71565
R2459 VTAIL.n292 VTAIL.n202 2.71565
R2460 VTAIL.n692 VTAIL.n602 2.71565
R2461 VTAIL.n664 VTAIL.n616 2.71565
R2462 VTAIL.n647 VTAIL.n646 2.71565
R2463 VTAIL.n592 VTAIL.n502 2.71565
R2464 VTAIL.n564 VTAIL.n516 2.71565
R2465 VTAIL.n547 VTAIL.n546 2.71565
R2466 VTAIL.n492 VTAIL.n402 2.71565
R2467 VTAIL.n464 VTAIL.n416 2.71565
R2468 VTAIL.n447 VTAIL.n446 2.71565
R2469 VTAIL.n392 VTAIL.n302 2.71565
R2470 VTAIL.n364 VTAIL.n316 2.71565
R2471 VTAIL.n347 VTAIL.n346 2.71565
R2472 VTAIL.n750 VTAIL.n724 1.93989
R2473 VTAIL.n763 VTAIL.n718 1.93989
R2474 VTAIL.n796 VTAIL.n795 1.93989
R2475 VTAIL.n50 VTAIL.n24 1.93989
R2476 VTAIL.n63 VTAIL.n18 1.93989
R2477 VTAIL.n96 VTAIL.n95 1.93989
R2478 VTAIL.n150 VTAIL.n124 1.93989
R2479 VTAIL.n163 VTAIL.n118 1.93989
R2480 VTAIL.n196 VTAIL.n195 1.93989
R2481 VTAIL.n250 VTAIL.n224 1.93989
R2482 VTAIL.n263 VTAIL.n218 1.93989
R2483 VTAIL.n296 VTAIL.n295 1.93989
R2484 VTAIL.n696 VTAIL.n695 1.93989
R2485 VTAIL.n663 VTAIL.n618 1.93989
R2486 VTAIL.n650 VTAIL.n624 1.93989
R2487 VTAIL.n596 VTAIL.n595 1.93989
R2488 VTAIL.n563 VTAIL.n518 1.93989
R2489 VTAIL.n550 VTAIL.n524 1.93989
R2490 VTAIL.n496 VTAIL.n495 1.93989
R2491 VTAIL.n463 VTAIL.n418 1.93989
R2492 VTAIL.n450 VTAIL.n424 1.93989
R2493 VTAIL.n396 VTAIL.n395 1.93989
R2494 VTAIL.n363 VTAIL.n318 1.93989
R2495 VTAIL.n350 VTAIL.n324 1.93989
R2496 VTAIL.n499 VTAIL.n399 1.56947
R2497 VTAIL.n699 VTAIL.n599 1.56947
R2498 VTAIL.n299 VTAIL.n199 1.56947
R2499 VTAIL.n751 VTAIL.n722 1.16414
R2500 VTAIL.n760 VTAIL.n759 1.16414
R2501 VTAIL.n798 VTAIL.n700 1.16414
R2502 VTAIL.n51 VTAIL.n22 1.16414
R2503 VTAIL.n60 VTAIL.n59 1.16414
R2504 VTAIL.n98 VTAIL.n0 1.16414
R2505 VTAIL.n151 VTAIL.n122 1.16414
R2506 VTAIL.n160 VTAIL.n159 1.16414
R2507 VTAIL.n198 VTAIL.n100 1.16414
R2508 VTAIL.n251 VTAIL.n222 1.16414
R2509 VTAIL.n260 VTAIL.n259 1.16414
R2510 VTAIL.n298 VTAIL.n200 1.16414
R2511 VTAIL.n698 VTAIL.n600 1.16414
R2512 VTAIL.n660 VTAIL.n659 1.16414
R2513 VTAIL.n651 VTAIL.n622 1.16414
R2514 VTAIL.n598 VTAIL.n500 1.16414
R2515 VTAIL.n560 VTAIL.n559 1.16414
R2516 VTAIL.n551 VTAIL.n522 1.16414
R2517 VTAIL.n498 VTAIL.n400 1.16414
R2518 VTAIL.n460 VTAIL.n459 1.16414
R2519 VTAIL.n451 VTAIL.n422 1.16414
R2520 VTAIL.n398 VTAIL.n300 1.16414
R2521 VTAIL.n360 VTAIL.n359 1.16414
R2522 VTAIL.n351 VTAIL.n322 1.16414
R2523 VTAIL VTAIL.n99 0.843172
R2524 VTAIL VTAIL.n799 0.726793
R2525 VTAIL.n599 VTAIL.n499 0.470328
R2526 VTAIL.n199 VTAIL.n99 0.470328
R2527 VTAIL.n755 VTAIL.n754 0.388379
R2528 VTAIL.n756 VTAIL.n720 0.388379
R2529 VTAIL.n55 VTAIL.n54 0.388379
R2530 VTAIL.n56 VTAIL.n20 0.388379
R2531 VTAIL.n155 VTAIL.n154 0.388379
R2532 VTAIL.n156 VTAIL.n120 0.388379
R2533 VTAIL.n255 VTAIL.n254 0.388379
R2534 VTAIL.n256 VTAIL.n220 0.388379
R2535 VTAIL.n656 VTAIL.n620 0.388379
R2536 VTAIL.n655 VTAIL.n654 0.388379
R2537 VTAIL.n556 VTAIL.n520 0.388379
R2538 VTAIL.n555 VTAIL.n554 0.388379
R2539 VTAIL.n456 VTAIL.n420 0.388379
R2540 VTAIL.n455 VTAIL.n454 0.388379
R2541 VTAIL.n356 VTAIL.n320 0.388379
R2542 VTAIL.n355 VTAIL.n354 0.388379
R2543 VTAIL.n736 VTAIL.n735 0.155672
R2544 VTAIL.n736 VTAIL.n727 0.155672
R2545 VTAIL.n743 VTAIL.n727 0.155672
R2546 VTAIL.n744 VTAIL.n743 0.155672
R2547 VTAIL.n744 VTAIL.n723 0.155672
R2548 VTAIL.n752 VTAIL.n723 0.155672
R2549 VTAIL.n753 VTAIL.n752 0.155672
R2550 VTAIL.n753 VTAIL.n719 0.155672
R2551 VTAIL.n761 VTAIL.n719 0.155672
R2552 VTAIL.n762 VTAIL.n761 0.155672
R2553 VTAIL.n762 VTAIL.n715 0.155672
R2554 VTAIL.n769 VTAIL.n715 0.155672
R2555 VTAIL.n770 VTAIL.n769 0.155672
R2556 VTAIL.n770 VTAIL.n711 0.155672
R2557 VTAIL.n777 VTAIL.n711 0.155672
R2558 VTAIL.n778 VTAIL.n777 0.155672
R2559 VTAIL.n778 VTAIL.n707 0.155672
R2560 VTAIL.n785 VTAIL.n707 0.155672
R2561 VTAIL.n786 VTAIL.n785 0.155672
R2562 VTAIL.n786 VTAIL.n703 0.155672
R2563 VTAIL.n793 VTAIL.n703 0.155672
R2564 VTAIL.n794 VTAIL.n793 0.155672
R2565 VTAIL.n36 VTAIL.n35 0.155672
R2566 VTAIL.n36 VTAIL.n27 0.155672
R2567 VTAIL.n43 VTAIL.n27 0.155672
R2568 VTAIL.n44 VTAIL.n43 0.155672
R2569 VTAIL.n44 VTAIL.n23 0.155672
R2570 VTAIL.n52 VTAIL.n23 0.155672
R2571 VTAIL.n53 VTAIL.n52 0.155672
R2572 VTAIL.n53 VTAIL.n19 0.155672
R2573 VTAIL.n61 VTAIL.n19 0.155672
R2574 VTAIL.n62 VTAIL.n61 0.155672
R2575 VTAIL.n62 VTAIL.n15 0.155672
R2576 VTAIL.n69 VTAIL.n15 0.155672
R2577 VTAIL.n70 VTAIL.n69 0.155672
R2578 VTAIL.n70 VTAIL.n11 0.155672
R2579 VTAIL.n77 VTAIL.n11 0.155672
R2580 VTAIL.n78 VTAIL.n77 0.155672
R2581 VTAIL.n78 VTAIL.n7 0.155672
R2582 VTAIL.n85 VTAIL.n7 0.155672
R2583 VTAIL.n86 VTAIL.n85 0.155672
R2584 VTAIL.n86 VTAIL.n3 0.155672
R2585 VTAIL.n93 VTAIL.n3 0.155672
R2586 VTAIL.n94 VTAIL.n93 0.155672
R2587 VTAIL.n136 VTAIL.n135 0.155672
R2588 VTAIL.n136 VTAIL.n127 0.155672
R2589 VTAIL.n143 VTAIL.n127 0.155672
R2590 VTAIL.n144 VTAIL.n143 0.155672
R2591 VTAIL.n144 VTAIL.n123 0.155672
R2592 VTAIL.n152 VTAIL.n123 0.155672
R2593 VTAIL.n153 VTAIL.n152 0.155672
R2594 VTAIL.n153 VTAIL.n119 0.155672
R2595 VTAIL.n161 VTAIL.n119 0.155672
R2596 VTAIL.n162 VTAIL.n161 0.155672
R2597 VTAIL.n162 VTAIL.n115 0.155672
R2598 VTAIL.n169 VTAIL.n115 0.155672
R2599 VTAIL.n170 VTAIL.n169 0.155672
R2600 VTAIL.n170 VTAIL.n111 0.155672
R2601 VTAIL.n177 VTAIL.n111 0.155672
R2602 VTAIL.n178 VTAIL.n177 0.155672
R2603 VTAIL.n178 VTAIL.n107 0.155672
R2604 VTAIL.n185 VTAIL.n107 0.155672
R2605 VTAIL.n186 VTAIL.n185 0.155672
R2606 VTAIL.n186 VTAIL.n103 0.155672
R2607 VTAIL.n193 VTAIL.n103 0.155672
R2608 VTAIL.n194 VTAIL.n193 0.155672
R2609 VTAIL.n236 VTAIL.n235 0.155672
R2610 VTAIL.n236 VTAIL.n227 0.155672
R2611 VTAIL.n243 VTAIL.n227 0.155672
R2612 VTAIL.n244 VTAIL.n243 0.155672
R2613 VTAIL.n244 VTAIL.n223 0.155672
R2614 VTAIL.n252 VTAIL.n223 0.155672
R2615 VTAIL.n253 VTAIL.n252 0.155672
R2616 VTAIL.n253 VTAIL.n219 0.155672
R2617 VTAIL.n261 VTAIL.n219 0.155672
R2618 VTAIL.n262 VTAIL.n261 0.155672
R2619 VTAIL.n262 VTAIL.n215 0.155672
R2620 VTAIL.n269 VTAIL.n215 0.155672
R2621 VTAIL.n270 VTAIL.n269 0.155672
R2622 VTAIL.n270 VTAIL.n211 0.155672
R2623 VTAIL.n277 VTAIL.n211 0.155672
R2624 VTAIL.n278 VTAIL.n277 0.155672
R2625 VTAIL.n278 VTAIL.n207 0.155672
R2626 VTAIL.n285 VTAIL.n207 0.155672
R2627 VTAIL.n286 VTAIL.n285 0.155672
R2628 VTAIL.n286 VTAIL.n203 0.155672
R2629 VTAIL.n293 VTAIL.n203 0.155672
R2630 VTAIL.n294 VTAIL.n293 0.155672
R2631 VTAIL.n694 VTAIL.n693 0.155672
R2632 VTAIL.n693 VTAIL.n603 0.155672
R2633 VTAIL.n686 VTAIL.n603 0.155672
R2634 VTAIL.n686 VTAIL.n685 0.155672
R2635 VTAIL.n685 VTAIL.n607 0.155672
R2636 VTAIL.n678 VTAIL.n607 0.155672
R2637 VTAIL.n678 VTAIL.n677 0.155672
R2638 VTAIL.n677 VTAIL.n611 0.155672
R2639 VTAIL.n670 VTAIL.n611 0.155672
R2640 VTAIL.n670 VTAIL.n669 0.155672
R2641 VTAIL.n669 VTAIL.n615 0.155672
R2642 VTAIL.n662 VTAIL.n615 0.155672
R2643 VTAIL.n662 VTAIL.n661 0.155672
R2644 VTAIL.n661 VTAIL.n619 0.155672
R2645 VTAIL.n653 VTAIL.n619 0.155672
R2646 VTAIL.n653 VTAIL.n652 0.155672
R2647 VTAIL.n652 VTAIL.n623 0.155672
R2648 VTAIL.n645 VTAIL.n623 0.155672
R2649 VTAIL.n645 VTAIL.n644 0.155672
R2650 VTAIL.n644 VTAIL.n628 0.155672
R2651 VTAIL.n637 VTAIL.n628 0.155672
R2652 VTAIL.n637 VTAIL.n636 0.155672
R2653 VTAIL.n594 VTAIL.n593 0.155672
R2654 VTAIL.n593 VTAIL.n503 0.155672
R2655 VTAIL.n586 VTAIL.n503 0.155672
R2656 VTAIL.n586 VTAIL.n585 0.155672
R2657 VTAIL.n585 VTAIL.n507 0.155672
R2658 VTAIL.n578 VTAIL.n507 0.155672
R2659 VTAIL.n578 VTAIL.n577 0.155672
R2660 VTAIL.n577 VTAIL.n511 0.155672
R2661 VTAIL.n570 VTAIL.n511 0.155672
R2662 VTAIL.n570 VTAIL.n569 0.155672
R2663 VTAIL.n569 VTAIL.n515 0.155672
R2664 VTAIL.n562 VTAIL.n515 0.155672
R2665 VTAIL.n562 VTAIL.n561 0.155672
R2666 VTAIL.n561 VTAIL.n519 0.155672
R2667 VTAIL.n553 VTAIL.n519 0.155672
R2668 VTAIL.n553 VTAIL.n552 0.155672
R2669 VTAIL.n552 VTAIL.n523 0.155672
R2670 VTAIL.n545 VTAIL.n523 0.155672
R2671 VTAIL.n545 VTAIL.n544 0.155672
R2672 VTAIL.n544 VTAIL.n528 0.155672
R2673 VTAIL.n537 VTAIL.n528 0.155672
R2674 VTAIL.n537 VTAIL.n536 0.155672
R2675 VTAIL.n494 VTAIL.n493 0.155672
R2676 VTAIL.n493 VTAIL.n403 0.155672
R2677 VTAIL.n486 VTAIL.n403 0.155672
R2678 VTAIL.n486 VTAIL.n485 0.155672
R2679 VTAIL.n485 VTAIL.n407 0.155672
R2680 VTAIL.n478 VTAIL.n407 0.155672
R2681 VTAIL.n478 VTAIL.n477 0.155672
R2682 VTAIL.n477 VTAIL.n411 0.155672
R2683 VTAIL.n470 VTAIL.n411 0.155672
R2684 VTAIL.n470 VTAIL.n469 0.155672
R2685 VTAIL.n469 VTAIL.n415 0.155672
R2686 VTAIL.n462 VTAIL.n415 0.155672
R2687 VTAIL.n462 VTAIL.n461 0.155672
R2688 VTAIL.n461 VTAIL.n419 0.155672
R2689 VTAIL.n453 VTAIL.n419 0.155672
R2690 VTAIL.n453 VTAIL.n452 0.155672
R2691 VTAIL.n452 VTAIL.n423 0.155672
R2692 VTAIL.n445 VTAIL.n423 0.155672
R2693 VTAIL.n445 VTAIL.n444 0.155672
R2694 VTAIL.n444 VTAIL.n428 0.155672
R2695 VTAIL.n437 VTAIL.n428 0.155672
R2696 VTAIL.n437 VTAIL.n436 0.155672
R2697 VTAIL.n394 VTAIL.n393 0.155672
R2698 VTAIL.n393 VTAIL.n303 0.155672
R2699 VTAIL.n386 VTAIL.n303 0.155672
R2700 VTAIL.n386 VTAIL.n385 0.155672
R2701 VTAIL.n385 VTAIL.n307 0.155672
R2702 VTAIL.n378 VTAIL.n307 0.155672
R2703 VTAIL.n378 VTAIL.n377 0.155672
R2704 VTAIL.n377 VTAIL.n311 0.155672
R2705 VTAIL.n370 VTAIL.n311 0.155672
R2706 VTAIL.n370 VTAIL.n369 0.155672
R2707 VTAIL.n369 VTAIL.n315 0.155672
R2708 VTAIL.n362 VTAIL.n315 0.155672
R2709 VTAIL.n362 VTAIL.n361 0.155672
R2710 VTAIL.n361 VTAIL.n319 0.155672
R2711 VTAIL.n353 VTAIL.n319 0.155672
R2712 VTAIL.n353 VTAIL.n352 0.155672
R2713 VTAIL.n352 VTAIL.n323 0.155672
R2714 VTAIL.n345 VTAIL.n323 0.155672
R2715 VTAIL.n345 VTAIL.n344 0.155672
R2716 VTAIL.n344 VTAIL.n328 0.155672
R2717 VTAIL.n337 VTAIL.n328 0.155672
R2718 VTAIL.n337 VTAIL.n336 0.155672
R2719 VP.n2 VP.t0 328.408
R2720 VP.n2 VP.t2 328.091
R2721 VP.n4 VP.t3 292.111
R2722 VP.n11 VP.t1 292.111
R2723 VP.n4 VP.n3 178.023
R2724 VP.n12 VP.n11 178.023
R2725 VP.n10 VP.n0 161.3
R2726 VP.n9 VP.n8 161.3
R2727 VP.n7 VP.n1 161.3
R2728 VP.n6 VP.n5 161.3
R2729 VP.n3 VP.n2 60.4515
R2730 VP.n9 VP.n1 56.5617
R2731 VP.n5 VP.n1 24.5923
R2732 VP.n10 VP.n9 24.5923
R2733 VP.n5 VP.n4 7.86989
R2734 VP.n11 VP.n10 7.86989
R2735 VP.n6 VP.n3 0.189894
R2736 VP.n7 VP.n6 0.189894
R2737 VP.n8 VP.n7 0.189894
R2738 VP.n8 VP.n0 0.189894
R2739 VP.n12 VP.n0 0.189894
R2740 VP VP.n12 0.0516364
R2741 VDD1 VDD1.n1 108.114
R2742 VDD1 VDD1.n0 63.6549
R2743 VDD1.n0 VDD1.t3 1.09685
R2744 VDD1.n0 VDD1.t1 1.09685
R2745 VDD1.n1 VDD1.t0 1.09685
R2746 VDD1.n1 VDD1.t2 1.09685
C0 VDD2 VN 6.13358f
C1 VDD1 VDD2 0.757267f
C2 VP VTAIL 5.6443f
C3 VP VN 6.51152f
C4 VDD1 VP 6.3088f
C5 VDD2 VP 0.324125f
C6 VN VTAIL 5.63019f
C7 VDD1 VTAIL 7.37016f
C8 VDD2 VTAIL 7.416931f
C9 VDD1 VN 0.148448f
C10 VDD2 B 3.617726f
C11 VDD1 B 8.057301f
C12 VTAIL B 12.959926f
C13 VN B 9.44524f
C14 VP B 6.976241f
C15 VDD1.t3 B 0.381333f
C16 VDD1.t1 B 0.381333f
C17 VDD1.n0 B 3.48498f
C18 VDD1.t0 B 0.381333f
C19 VDD1.t2 B 0.381333f
C20 VDD1.n1 B 4.32603f
C21 VP.n0 B 0.034651f
C22 VP.t1 B 2.56492f
C23 VP.n1 B 0.050371f
C24 VP.t0 B 2.67987f
C25 VP.t2 B 2.67885f
C26 VP.n2 B 3.41264f
C27 VP.n3 B 2.18665f
C28 VP.t3 B 2.56492f
C29 VP.n4 B 0.969615f
C30 VP.n5 B 0.042686f
C31 VP.n6 B 0.034651f
C32 VP.n7 B 0.034651f
C33 VP.n8 B 0.034651f
C34 VP.n9 B 0.050371f
C35 VP.n10 B 0.042686f
C36 VP.n11 B 0.969615f
C37 VP.n12 B 0.033783f
C38 VTAIL.n0 B 0.008472f
C39 VTAIL.n1 B 0.0191f
C40 VTAIL.n2 B 0.008556f
C41 VTAIL.n3 B 0.015038f
C42 VTAIL.n4 B 0.008081f
C43 VTAIL.n5 B 0.0191f
C44 VTAIL.n6 B 0.008556f
C45 VTAIL.n7 B 0.015038f
C46 VTAIL.n8 B 0.008081f
C47 VTAIL.n9 B 0.0191f
C48 VTAIL.n10 B 0.008556f
C49 VTAIL.n11 B 0.015038f
C50 VTAIL.n12 B 0.008081f
C51 VTAIL.n13 B 0.0191f
C52 VTAIL.n14 B 0.008556f
C53 VTAIL.n15 B 0.015038f
C54 VTAIL.n16 B 0.008081f
C55 VTAIL.n17 B 0.0191f
C56 VTAIL.n18 B 0.008556f
C57 VTAIL.n19 B 0.015038f
C58 VTAIL.n20 B 0.008081f
C59 VTAIL.n21 B 0.0191f
C60 VTAIL.n22 B 0.008556f
C61 VTAIL.n23 B 0.015038f
C62 VTAIL.n24 B 0.008081f
C63 VTAIL.n25 B 0.0191f
C64 VTAIL.n26 B 0.008556f
C65 VTAIL.n27 B 0.015038f
C66 VTAIL.n28 B 0.008081f
C67 VTAIL.n29 B 0.0191f
C68 VTAIL.n30 B 0.008556f
C69 VTAIL.n31 B 0.143409f
C70 VTAIL.t6 B 0.032749f
C71 VTAIL.n32 B 0.014325f
C72 VTAIL.n33 B 0.013502f
C73 VTAIL.n34 B 0.008081f
C74 VTAIL.n35 B 1.16398f
C75 VTAIL.n36 B 0.015038f
C76 VTAIL.n37 B 0.008081f
C77 VTAIL.n38 B 0.008556f
C78 VTAIL.n39 B 0.0191f
C79 VTAIL.n40 B 0.0191f
C80 VTAIL.n41 B 0.008556f
C81 VTAIL.n42 B 0.008081f
C82 VTAIL.n43 B 0.015038f
C83 VTAIL.n44 B 0.015038f
C84 VTAIL.n45 B 0.008081f
C85 VTAIL.n46 B 0.008556f
C86 VTAIL.n47 B 0.0191f
C87 VTAIL.n48 B 0.0191f
C88 VTAIL.n49 B 0.0191f
C89 VTAIL.n50 B 0.008556f
C90 VTAIL.n51 B 0.008081f
C91 VTAIL.n52 B 0.015038f
C92 VTAIL.n53 B 0.015038f
C93 VTAIL.n54 B 0.008081f
C94 VTAIL.n55 B 0.008318f
C95 VTAIL.n56 B 0.008318f
C96 VTAIL.n57 B 0.0191f
C97 VTAIL.n58 B 0.0191f
C98 VTAIL.n59 B 0.008556f
C99 VTAIL.n60 B 0.008081f
C100 VTAIL.n61 B 0.015038f
C101 VTAIL.n62 B 0.015038f
C102 VTAIL.n63 B 0.008081f
C103 VTAIL.n64 B 0.008556f
C104 VTAIL.n65 B 0.0191f
C105 VTAIL.n66 B 0.0191f
C106 VTAIL.n67 B 0.008556f
C107 VTAIL.n68 B 0.008081f
C108 VTAIL.n69 B 0.015038f
C109 VTAIL.n70 B 0.015038f
C110 VTAIL.n71 B 0.008081f
C111 VTAIL.n72 B 0.008556f
C112 VTAIL.n73 B 0.0191f
C113 VTAIL.n74 B 0.0191f
C114 VTAIL.n75 B 0.008556f
C115 VTAIL.n76 B 0.008081f
C116 VTAIL.n77 B 0.015038f
C117 VTAIL.n78 B 0.015038f
C118 VTAIL.n79 B 0.008081f
C119 VTAIL.n80 B 0.008556f
C120 VTAIL.n81 B 0.0191f
C121 VTAIL.n82 B 0.0191f
C122 VTAIL.n83 B 0.008556f
C123 VTAIL.n84 B 0.008081f
C124 VTAIL.n85 B 0.015038f
C125 VTAIL.n86 B 0.015038f
C126 VTAIL.n87 B 0.008081f
C127 VTAIL.n88 B 0.008556f
C128 VTAIL.n89 B 0.0191f
C129 VTAIL.n90 B 0.0191f
C130 VTAIL.n91 B 0.008556f
C131 VTAIL.n92 B 0.008081f
C132 VTAIL.n93 B 0.015038f
C133 VTAIL.n94 B 0.038457f
C134 VTAIL.n95 B 0.008081f
C135 VTAIL.n96 B 0.008556f
C136 VTAIL.n97 B 0.038119f
C137 VTAIL.n98 B 0.032168f
C138 VTAIL.n99 B 0.077835f
C139 VTAIL.n100 B 0.008472f
C140 VTAIL.n101 B 0.0191f
C141 VTAIL.n102 B 0.008556f
C142 VTAIL.n103 B 0.015038f
C143 VTAIL.n104 B 0.008081f
C144 VTAIL.n105 B 0.0191f
C145 VTAIL.n106 B 0.008556f
C146 VTAIL.n107 B 0.015038f
C147 VTAIL.n108 B 0.008081f
C148 VTAIL.n109 B 0.0191f
C149 VTAIL.n110 B 0.008556f
C150 VTAIL.n111 B 0.015038f
C151 VTAIL.n112 B 0.008081f
C152 VTAIL.n113 B 0.0191f
C153 VTAIL.n114 B 0.008556f
C154 VTAIL.n115 B 0.015038f
C155 VTAIL.n116 B 0.008081f
C156 VTAIL.n117 B 0.0191f
C157 VTAIL.n118 B 0.008556f
C158 VTAIL.n119 B 0.015038f
C159 VTAIL.n120 B 0.008081f
C160 VTAIL.n121 B 0.0191f
C161 VTAIL.n122 B 0.008556f
C162 VTAIL.n123 B 0.015038f
C163 VTAIL.n124 B 0.008081f
C164 VTAIL.n125 B 0.0191f
C165 VTAIL.n126 B 0.008556f
C166 VTAIL.n127 B 0.015038f
C167 VTAIL.n128 B 0.008081f
C168 VTAIL.n129 B 0.0191f
C169 VTAIL.n130 B 0.008556f
C170 VTAIL.n131 B 0.143409f
C171 VTAIL.t0 B 0.032749f
C172 VTAIL.n132 B 0.014325f
C173 VTAIL.n133 B 0.013502f
C174 VTAIL.n134 B 0.008081f
C175 VTAIL.n135 B 1.16398f
C176 VTAIL.n136 B 0.015038f
C177 VTAIL.n137 B 0.008081f
C178 VTAIL.n138 B 0.008556f
C179 VTAIL.n139 B 0.0191f
C180 VTAIL.n140 B 0.0191f
C181 VTAIL.n141 B 0.008556f
C182 VTAIL.n142 B 0.008081f
C183 VTAIL.n143 B 0.015038f
C184 VTAIL.n144 B 0.015038f
C185 VTAIL.n145 B 0.008081f
C186 VTAIL.n146 B 0.008556f
C187 VTAIL.n147 B 0.0191f
C188 VTAIL.n148 B 0.0191f
C189 VTAIL.n149 B 0.0191f
C190 VTAIL.n150 B 0.008556f
C191 VTAIL.n151 B 0.008081f
C192 VTAIL.n152 B 0.015038f
C193 VTAIL.n153 B 0.015038f
C194 VTAIL.n154 B 0.008081f
C195 VTAIL.n155 B 0.008318f
C196 VTAIL.n156 B 0.008318f
C197 VTAIL.n157 B 0.0191f
C198 VTAIL.n158 B 0.0191f
C199 VTAIL.n159 B 0.008556f
C200 VTAIL.n160 B 0.008081f
C201 VTAIL.n161 B 0.015038f
C202 VTAIL.n162 B 0.015038f
C203 VTAIL.n163 B 0.008081f
C204 VTAIL.n164 B 0.008556f
C205 VTAIL.n165 B 0.0191f
C206 VTAIL.n166 B 0.0191f
C207 VTAIL.n167 B 0.008556f
C208 VTAIL.n168 B 0.008081f
C209 VTAIL.n169 B 0.015038f
C210 VTAIL.n170 B 0.015038f
C211 VTAIL.n171 B 0.008081f
C212 VTAIL.n172 B 0.008556f
C213 VTAIL.n173 B 0.0191f
C214 VTAIL.n174 B 0.0191f
C215 VTAIL.n175 B 0.008556f
C216 VTAIL.n176 B 0.008081f
C217 VTAIL.n177 B 0.015038f
C218 VTAIL.n178 B 0.015038f
C219 VTAIL.n179 B 0.008081f
C220 VTAIL.n180 B 0.008556f
C221 VTAIL.n181 B 0.0191f
C222 VTAIL.n182 B 0.0191f
C223 VTAIL.n183 B 0.008556f
C224 VTAIL.n184 B 0.008081f
C225 VTAIL.n185 B 0.015038f
C226 VTAIL.n186 B 0.015038f
C227 VTAIL.n187 B 0.008081f
C228 VTAIL.n188 B 0.008556f
C229 VTAIL.n189 B 0.0191f
C230 VTAIL.n190 B 0.0191f
C231 VTAIL.n191 B 0.008556f
C232 VTAIL.n192 B 0.008081f
C233 VTAIL.n193 B 0.015038f
C234 VTAIL.n194 B 0.038457f
C235 VTAIL.n195 B 0.008081f
C236 VTAIL.n196 B 0.008556f
C237 VTAIL.n197 B 0.038119f
C238 VTAIL.n198 B 0.032168f
C239 VTAIL.n199 B 0.113028f
C240 VTAIL.n200 B 0.008472f
C241 VTAIL.n201 B 0.0191f
C242 VTAIL.n202 B 0.008556f
C243 VTAIL.n203 B 0.015038f
C244 VTAIL.n204 B 0.008081f
C245 VTAIL.n205 B 0.0191f
C246 VTAIL.n206 B 0.008556f
C247 VTAIL.n207 B 0.015038f
C248 VTAIL.n208 B 0.008081f
C249 VTAIL.n209 B 0.0191f
C250 VTAIL.n210 B 0.008556f
C251 VTAIL.n211 B 0.015038f
C252 VTAIL.n212 B 0.008081f
C253 VTAIL.n213 B 0.0191f
C254 VTAIL.n214 B 0.008556f
C255 VTAIL.n215 B 0.015038f
C256 VTAIL.n216 B 0.008081f
C257 VTAIL.n217 B 0.0191f
C258 VTAIL.n218 B 0.008556f
C259 VTAIL.n219 B 0.015038f
C260 VTAIL.n220 B 0.008081f
C261 VTAIL.n221 B 0.0191f
C262 VTAIL.n222 B 0.008556f
C263 VTAIL.n223 B 0.015038f
C264 VTAIL.n224 B 0.008081f
C265 VTAIL.n225 B 0.0191f
C266 VTAIL.n226 B 0.008556f
C267 VTAIL.n227 B 0.015038f
C268 VTAIL.n228 B 0.008081f
C269 VTAIL.n229 B 0.0191f
C270 VTAIL.n230 B 0.008556f
C271 VTAIL.n231 B 0.143409f
C272 VTAIL.t3 B 0.032749f
C273 VTAIL.n232 B 0.014325f
C274 VTAIL.n233 B 0.013502f
C275 VTAIL.n234 B 0.008081f
C276 VTAIL.n235 B 1.16398f
C277 VTAIL.n236 B 0.015038f
C278 VTAIL.n237 B 0.008081f
C279 VTAIL.n238 B 0.008556f
C280 VTAIL.n239 B 0.0191f
C281 VTAIL.n240 B 0.0191f
C282 VTAIL.n241 B 0.008556f
C283 VTAIL.n242 B 0.008081f
C284 VTAIL.n243 B 0.015038f
C285 VTAIL.n244 B 0.015038f
C286 VTAIL.n245 B 0.008081f
C287 VTAIL.n246 B 0.008556f
C288 VTAIL.n247 B 0.0191f
C289 VTAIL.n248 B 0.0191f
C290 VTAIL.n249 B 0.0191f
C291 VTAIL.n250 B 0.008556f
C292 VTAIL.n251 B 0.008081f
C293 VTAIL.n252 B 0.015038f
C294 VTAIL.n253 B 0.015038f
C295 VTAIL.n254 B 0.008081f
C296 VTAIL.n255 B 0.008318f
C297 VTAIL.n256 B 0.008318f
C298 VTAIL.n257 B 0.0191f
C299 VTAIL.n258 B 0.0191f
C300 VTAIL.n259 B 0.008556f
C301 VTAIL.n260 B 0.008081f
C302 VTAIL.n261 B 0.015038f
C303 VTAIL.n262 B 0.015038f
C304 VTAIL.n263 B 0.008081f
C305 VTAIL.n264 B 0.008556f
C306 VTAIL.n265 B 0.0191f
C307 VTAIL.n266 B 0.0191f
C308 VTAIL.n267 B 0.008556f
C309 VTAIL.n268 B 0.008081f
C310 VTAIL.n269 B 0.015038f
C311 VTAIL.n270 B 0.015038f
C312 VTAIL.n271 B 0.008081f
C313 VTAIL.n272 B 0.008556f
C314 VTAIL.n273 B 0.0191f
C315 VTAIL.n274 B 0.0191f
C316 VTAIL.n275 B 0.008556f
C317 VTAIL.n276 B 0.008081f
C318 VTAIL.n277 B 0.015038f
C319 VTAIL.n278 B 0.015038f
C320 VTAIL.n279 B 0.008081f
C321 VTAIL.n280 B 0.008556f
C322 VTAIL.n281 B 0.0191f
C323 VTAIL.n282 B 0.0191f
C324 VTAIL.n283 B 0.008556f
C325 VTAIL.n284 B 0.008081f
C326 VTAIL.n285 B 0.015038f
C327 VTAIL.n286 B 0.015038f
C328 VTAIL.n287 B 0.008081f
C329 VTAIL.n288 B 0.008556f
C330 VTAIL.n289 B 0.0191f
C331 VTAIL.n290 B 0.0191f
C332 VTAIL.n291 B 0.008556f
C333 VTAIL.n292 B 0.008081f
C334 VTAIL.n293 B 0.015038f
C335 VTAIL.n294 B 0.038457f
C336 VTAIL.n295 B 0.008081f
C337 VTAIL.n296 B 0.008556f
C338 VTAIL.n297 B 0.038119f
C339 VTAIL.n298 B 0.032168f
C340 VTAIL.n299 B 1.12497f
C341 VTAIL.n300 B 0.008472f
C342 VTAIL.n301 B 0.0191f
C343 VTAIL.n302 B 0.008556f
C344 VTAIL.n303 B 0.015038f
C345 VTAIL.n304 B 0.008081f
C346 VTAIL.n305 B 0.0191f
C347 VTAIL.n306 B 0.008556f
C348 VTAIL.n307 B 0.015038f
C349 VTAIL.n308 B 0.008081f
C350 VTAIL.n309 B 0.0191f
C351 VTAIL.n310 B 0.008556f
C352 VTAIL.n311 B 0.015038f
C353 VTAIL.n312 B 0.008081f
C354 VTAIL.n313 B 0.0191f
C355 VTAIL.n314 B 0.008556f
C356 VTAIL.n315 B 0.015038f
C357 VTAIL.n316 B 0.008081f
C358 VTAIL.n317 B 0.0191f
C359 VTAIL.n318 B 0.008556f
C360 VTAIL.n319 B 0.015038f
C361 VTAIL.n320 B 0.008081f
C362 VTAIL.n321 B 0.0191f
C363 VTAIL.n322 B 0.008556f
C364 VTAIL.n323 B 0.015038f
C365 VTAIL.n324 B 0.008081f
C366 VTAIL.n325 B 0.0191f
C367 VTAIL.n326 B 0.0191f
C368 VTAIL.n327 B 0.008556f
C369 VTAIL.n328 B 0.015038f
C370 VTAIL.n329 B 0.008081f
C371 VTAIL.n330 B 0.0191f
C372 VTAIL.n331 B 0.008556f
C373 VTAIL.n332 B 0.143409f
C374 VTAIL.t7 B 0.032749f
C375 VTAIL.n333 B 0.014325f
C376 VTAIL.n334 B 0.013502f
C377 VTAIL.n335 B 0.008081f
C378 VTAIL.n336 B 1.16397f
C379 VTAIL.n337 B 0.015038f
C380 VTAIL.n338 B 0.008081f
C381 VTAIL.n339 B 0.008556f
C382 VTAIL.n340 B 0.0191f
C383 VTAIL.n341 B 0.0191f
C384 VTAIL.n342 B 0.008556f
C385 VTAIL.n343 B 0.008081f
C386 VTAIL.n344 B 0.015038f
C387 VTAIL.n345 B 0.015038f
C388 VTAIL.n346 B 0.008081f
C389 VTAIL.n347 B 0.008556f
C390 VTAIL.n348 B 0.0191f
C391 VTAIL.n349 B 0.0191f
C392 VTAIL.n350 B 0.008556f
C393 VTAIL.n351 B 0.008081f
C394 VTAIL.n352 B 0.015038f
C395 VTAIL.n353 B 0.015038f
C396 VTAIL.n354 B 0.008081f
C397 VTAIL.n355 B 0.008318f
C398 VTAIL.n356 B 0.008318f
C399 VTAIL.n357 B 0.0191f
C400 VTAIL.n358 B 0.0191f
C401 VTAIL.n359 B 0.008556f
C402 VTAIL.n360 B 0.008081f
C403 VTAIL.n361 B 0.015038f
C404 VTAIL.n362 B 0.015038f
C405 VTAIL.n363 B 0.008081f
C406 VTAIL.n364 B 0.008556f
C407 VTAIL.n365 B 0.0191f
C408 VTAIL.n366 B 0.0191f
C409 VTAIL.n367 B 0.008556f
C410 VTAIL.n368 B 0.008081f
C411 VTAIL.n369 B 0.015038f
C412 VTAIL.n370 B 0.015038f
C413 VTAIL.n371 B 0.008081f
C414 VTAIL.n372 B 0.008556f
C415 VTAIL.n373 B 0.0191f
C416 VTAIL.n374 B 0.0191f
C417 VTAIL.n375 B 0.008556f
C418 VTAIL.n376 B 0.008081f
C419 VTAIL.n377 B 0.015038f
C420 VTAIL.n378 B 0.015038f
C421 VTAIL.n379 B 0.008081f
C422 VTAIL.n380 B 0.008556f
C423 VTAIL.n381 B 0.0191f
C424 VTAIL.n382 B 0.0191f
C425 VTAIL.n383 B 0.008556f
C426 VTAIL.n384 B 0.008081f
C427 VTAIL.n385 B 0.015038f
C428 VTAIL.n386 B 0.015038f
C429 VTAIL.n387 B 0.008081f
C430 VTAIL.n388 B 0.008556f
C431 VTAIL.n389 B 0.0191f
C432 VTAIL.n390 B 0.0191f
C433 VTAIL.n391 B 0.008556f
C434 VTAIL.n392 B 0.008081f
C435 VTAIL.n393 B 0.015038f
C436 VTAIL.n394 B 0.038457f
C437 VTAIL.n395 B 0.008081f
C438 VTAIL.n396 B 0.008556f
C439 VTAIL.n397 B 0.038119f
C440 VTAIL.n398 B 0.032168f
C441 VTAIL.n399 B 1.12497f
C442 VTAIL.n400 B 0.008472f
C443 VTAIL.n401 B 0.0191f
C444 VTAIL.n402 B 0.008556f
C445 VTAIL.n403 B 0.015038f
C446 VTAIL.n404 B 0.008081f
C447 VTAIL.n405 B 0.0191f
C448 VTAIL.n406 B 0.008556f
C449 VTAIL.n407 B 0.015038f
C450 VTAIL.n408 B 0.008081f
C451 VTAIL.n409 B 0.0191f
C452 VTAIL.n410 B 0.008556f
C453 VTAIL.n411 B 0.015038f
C454 VTAIL.n412 B 0.008081f
C455 VTAIL.n413 B 0.0191f
C456 VTAIL.n414 B 0.008556f
C457 VTAIL.n415 B 0.015038f
C458 VTAIL.n416 B 0.008081f
C459 VTAIL.n417 B 0.0191f
C460 VTAIL.n418 B 0.008556f
C461 VTAIL.n419 B 0.015038f
C462 VTAIL.n420 B 0.008081f
C463 VTAIL.n421 B 0.0191f
C464 VTAIL.n422 B 0.008556f
C465 VTAIL.n423 B 0.015038f
C466 VTAIL.n424 B 0.008081f
C467 VTAIL.n425 B 0.0191f
C468 VTAIL.n426 B 0.0191f
C469 VTAIL.n427 B 0.008556f
C470 VTAIL.n428 B 0.015038f
C471 VTAIL.n429 B 0.008081f
C472 VTAIL.n430 B 0.0191f
C473 VTAIL.n431 B 0.008556f
C474 VTAIL.n432 B 0.143409f
C475 VTAIL.t4 B 0.032749f
C476 VTAIL.n433 B 0.014325f
C477 VTAIL.n434 B 0.013502f
C478 VTAIL.n435 B 0.008081f
C479 VTAIL.n436 B 1.16397f
C480 VTAIL.n437 B 0.015038f
C481 VTAIL.n438 B 0.008081f
C482 VTAIL.n439 B 0.008556f
C483 VTAIL.n440 B 0.0191f
C484 VTAIL.n441 B 0.0191f
C485 VTAIL.n442 B 0.008556f
C486 VTAIL.n443 B 0.008081f
C487 VTAIL.n444 B 0.015038f
C488 VTAIL.n445 B 0.015038f
C489 VTAIL.n446 B 0.008081f
C490 VTAIL.n447 B 0.008556f
C491 VTAIL.n448 B 0.0191f
C492 VTAIL.n449 B 0.0191f
C493 VTAIL.n450 B 0.008556f
C494 VTAIL.n451 B 0.008081f
C495 VTAIL.n452 B 0.015038f
C496 VTAIL.n453 B 0.015038f
C497 VTAIL.n454 B 0.008081f
C498 VTAIL.n455 B 0.008318f
C499 VTAIL.n456 B 0.008318f
C500 VTAIL.n457 B 0.0191f
C501 VTAIL.n458 B 0.0191f
C502 VTAIL.n459 B 0.008556f
C503 VTAIL.n460 B 0.008081f
C504 VTAIL.n461 B 0.015038f
C505 VTAIL.n462 B 0.015038f
C506 VTAIL.n463 B 0.008081f
C507 VTAIL.n464 B 0.008556f
C508 VTAIL.n465 B 0.0191f
C509 VTAIL.n466 B 0.0191f
C510 VTAIL.n467 B 0.008556f
C511 VTAIL.n468 B 0.008081f
C512 VTAIL.n469 B 0.015038f
C513 VTAIL.n470 B 0.015038f
C514 VTAIL.n471 B 0.008081f
C515 VTAIL.n472 B 0.008556f
C516 VTAIL.n473 B 0.0191f
C517 VTAIL.n474 B 0.0191f
C518 VTAIL.n475 B 0.008556f
C519 VTAIL.n476 B 0.008081f
C520 VTAIL.n477 B 0.015038f
C521 VTAIL.n478 B 0.015038f
C522 VTAIL.n479 B 0.008081f
C523 VTAIL.n480 B 0.008556f
C524 VTAIL.n481 B 0.0191f
C525 VTAIL.n482 B 0.0191f
C526 VTAIL.n483 B 0.008556f
C527 VTAIL.n484 B 0.008081f
C528 VTAIL.n485 B 0.015038f
C529 VTAIL.n486 B 0.015038f
C530 VTAIL.n487 B 0.008081f
C531 VTAIL.n488 B 0.008556f
C532 VTAIL.n489 B 0.0191f
C533 VTAIL.n490 B 0.0191f
C534 VTAIL.n491 B 0.008556f
C535 VTAIL.n492 B 0.008081f
C536 VTAIL.n493 B 0.015038f
C537 VTAIL.n494 B 0.038457f
C538 VTAIL.n495 B 0.008081f
C539 VTAIL.n496 B 0.008556f
C540 VTAIL.n497 B 0.038119f
C541 VTAIL.n498 B 0.032168f
C542 VTAIL.n499 B 0.113028f
C543 VTAIL.n500 B 0.008472f
C544 VTAIL.n501 B 0.0191f
C545 VTAIL.n502 B 0.008556f
C546 VTAIL.n503 B 0.015038f
C547 VTAIL.n504 B 0.008081f
C548 VTAIL.n505 B 0.0191f
C549 VTAIL.n506 B 0.008556f
C550 VTAIL.n507 B 0.015038f
C551 VTAIL.n508 B 0.008081f
C552 VTAIL.n509 B 0.0191f
C553 VTAIL.n510 B 0.008556f
C554 VTAIL.n511 B 0.015038f
C555 VTAIL.n512 B 0.008081f
C556 VTAIL.n513 B 0.0191f
C557 VTAIL.n514 B 0.008556f
C558 VTAIL.n515 B 0.015038f
C559 VTAIL.n516 B 0.008081f
C560 VTAIL.n517 B 0.0191f
C561 VTAIL.n518 B 0.008556f
C562 VTAIL.n519 B 0.015038f
C563 VTAIL.n520 B 0.008081f
C564 VTAIL.n521 B 0.0191f
C565 VTAIL.n522 B 0.008556f
C566 VTAIL.n523 B 0.015038f
C567 VTAIL.n524 B 0.008081f
C568 VTAIL.n525 B 0.0191f
C569 VTAIL.n526 B 0.0191f
C570 VTAIL.n527 B 0.008556f
C571 VTAIL.n528 B 0.015038f
C572 VTAIL.n529 B 0.008081f
C573 VTAIL.n530 B 0.0191f
C574 VTAIL.n531 B 0.008556f
C575 VTAIL.n532 B 0.143409f
C576 VTAIL.t2 B 0.032749f
C577 VTAIL.n533 B 0.014325f
C578 VTAIL.n534 B 0.013502f
C579 VTAIL.n535 B 0.008081f
C580 VTAIL.n536 B 1.16397f
C581 VTAIL.n537 B 0.015038f
C582 VTAIL.n538 B 0.008081f
C583 VTAIL.n539 B 0.008556f
C584 VTAIL.n540 B 0.0191f
C585 VTAIL.n541 B 0.0191f
C586 VTAIL.n542 B 0.008556f
C587 VTAIL.n543 B 0.008081f
C588 VTAIL.n544 B 0.015038f
C589 VTAIL.n545 B 0.015038f
C590 VTAIL.n546 B 0.008081f
C591 VTAIL.n547 B 0.008556f
C592 VTAIL.n548 B 0.0191f
C593 VTAIL.n549 B 0.0191f
C594 VTAIL.n550 B 0.008556f
C595 VTAIL.n551 B 0.008081f
C596 VTAIL.n552 B 0.015038f
C597 VTAIL.n553 B 0.015038f
C598 VTAIL.n554 B 0.008081f
C599 VTAIL.n555 B 0.008318f
C600 VTAIL.n556 B 0.008318f
C601 VTAIL.n557 B 0.0191f
C602 VTAIL.n558 B 0.0191f
C603 VTAIL.n559 B 0.008556f
C604 VTAIL.n560 B 0.008081f
C605 VTAIL.n561 B 0.015038f
C606 VTAIL.n562 B 0.015038f
C607 VTAIL.n563 B 0.008081f
C608 VTAIL.n564 B 0.008556f
C609 VTAIL.n565 B 0.0191f
C610 VTAIL.n566 B 0.0191f
C611 VTAIL.n567 B 0.008556f
C612 VTAIL.n568 B 0.008081f
C613 VTAIL.n569 B 0.015038f
C614 VTAIL.n570 B 0.015038f
C615 VTAIL.n571 B 0.008081f
C616 VTAIL.n572 B 0.008556f
C617 VTAIL.n573 B 0.0191f
C618 VTAIL.n574 B 0.0191f
C619 VTAIL.n575 B 0.008556f
C620 VTAIL.n576 B 0.008081f
C621 VTAIL.n577 B 0.015038f
C622 VTAIL.n578 B 0.015038f
C623 VTAIL.n579 B 0.008081f
C624 VTAIL.n580 B 0.008556f
C625 VTAIL.n581 B 0.0191f
C626 VTAIL.n582 B 0.0191f
C627 VTAIL.n583 B 0.008556f
C628 VTAIL.n584 B 0.008081f
C629 VTAIL.n585 B 0.015038f
C630 VTAIL.n586 B 0.015038f
C631 VTAIL.n587 B 0.008081f
C632 VTAIL.n588 B 0.008556f
C633 VTAIL.n589 B 0.0191f
C634 VTAIL.n590 B 0.0191f
C635 VTAIL.n591 B 0.008556f
C636 VTAIL.n592 B 0.008081f
C637 VTAIL.n593 B 0.015038f
C638 VTAIL.n594 B 0.038457f
C639 VTAIL.n595 B 0.008081f
C640 VTAIL.n596 B 0.008556f
C641 VTAIL.n597 B 0.038119f
C642 VTAIL.n598 B 0.032168f
C643 VTAIL.n599 B 0.113028f
C644 VTAIL.n600 B 0.008472f
C645 VTAIL.n601 B 0.0191f
C646 VTAIL.n602 B 0.008556f
C647 VTAIL.n603 B 0.015038f
C648 VTAIL.n604 B 0.008081f
C649 VTAIL.n605 B 0.0191f
C650 VTAIL.n606 B 0.008556f
C651 VTAIL.n607 B 0.015038f
C652 VTAIL.n608 B 0.008081f
C653 VTAIL.n609 B 0.0191f
C654 VTAIL.n610 B 0.008556f
C655 VTAIL.n611 B 0.015038f
C656 VTAIL.n612 B 0.008081f
C657 VTAIL.n613 B 0.0191f
C658 VTAIL.n614 B 0.008556f
C659 VTAIL.n615 B 0.015038f
C660 VTAIL.n616 B 0.008081f
C661 VTAIL.n617 B 0.0191f
C662 VTAIL.n618 B 0.008556f
C663 VTAIL.n619 B 0.015038f
C664 VTAIL.n620 B 0.008081f
C665 VTAIL.n621 B 0.0191f
C666 VTAIL.n622 B 0.008556f
C667 VTAIL.n623 B 0.015038f
C668 VTAIL.n624 B 0.008081f
C669 VTAIL.n625 B 0.0191f
C670 VTAIL.n626 B 0.0191f
C671 VTAIL.n627 B 0.008556f
C672 VTAIL.n628 B 0.015038f
C673 VTAIL.n629 B 0.008081f
C674 VTAIL.n630 B 0.0191f
C675 VTAIL.n631 B 0.008556f
C676 VTAIL.n632 B 0.143409f
C677 VTAIL.t1 B 0.032749f
C678 VTAIL.n633 B 0.014325f
C679 VTAIL.n634 B 0.013502f
C680 VTAIL.n635 B 0.008081f
C681 VTAIL.n636 B 1.16398f
C682 VTAIL.n637 B 0.015038f
C683 VTAIL.n638 B 0.008081f
C684 VTAIL.n639 B 0.008556f
C685 VTAIL.n640 B 0.0191f
C686 VTAIL.n641 B 0.0191f
C687 VTAIL.n642 B 0.008556f
C688 VTAIL.n643 B 0.008081f
C689 VTAIL.n644 B 0.015038f
C690 VTAIL.n645 B 0.015038f
C691 VTAIL.n646 B 0.008081f
C692 VTAIL.n647 B 0.008556f
C693 VTAIL.n648 B 0.0191f
C694 VTAIL.n649 B 0.0191f
C695 VTAIL.n650 B 0.008556f
C696 VTAIL.n651 B 0.008081f
C697 VTAIL.n652 B 0.015038f
C698 VTAIL.n653 B 0.015038f
C699 VTAIL.n654 B 0.008081f
C700 VTAIL.n655 B 0.008318f
C701 VTAIL.n656 B 0.008318f
C702 VTAIL.n657 B 0.0191f
C703 VTAIL.n658 B 0.0191f
C704 VTAIL.n659 B 0.008556f
C705 VTAIL.n660 B 0.008081f
C706 VTAIL.n661 B 0.015038f
C707 VTAIL.n662 B 0.015038f
C708 VTAIL.n663 B 0.008081f
C709 VTAIL.n664 B 0.008556f
C710 VTAIL.n665 B 0.0191f
C711 VTAIL.n666 B 0.0191f
C712 VTAIL.n667 B 0.008556f
C713 VTAIL.n668 B 0.008081f
C714 VTAIL.n669 B 0.015038f
C715 VTAIL.n670 B 0.015038f
C716 VTAIL.n671 B 0.008081f
C717 VTAIL.n672 B 0.008556f
C718 VTAIL.n673 B 0.0191f
C719 VTAIL.n674 B 0.0191f
C720 VTAIL.n675 B 0.008556f
C721 VTAIL.n676 B 0.008081f
C722 VTAIL.n677 B 0.015038f
C723 VTAIL.n678 B 0.015038f
C724 VTAIL.n679 B 0.008081f
C725 VTAIL.n680 B 0.008556f
C726 VTAIL.n681 B 0.0191f
C727 VTAIL.n682 B 0.0191f
C728 VTAIL.n683 B 0.008556f
C729 VTAIL.n684 B 0.008081f
C730 VTAIL.n685 B 0.015038f
C731 VTAIL.n686 B 0.015038f
C732 VTAIL.n687 B 0.008081f
C733 VTAIL.n688 B 0.008556f
C734 VTAIL.n689 B 0.0191f
C735 VTAIL.n690 B 0.0191f
C736 VTAIL.n691 B 0.008556f
C737 VTAIL.n692 B 0.008081f
C738 VTAIL.n693 B 0.015038f
C739 VTAIL.n694 B 0.038457f
C740 VTAIL.n695 B 0.008081f
C741 VTAIL.n696 B 0.008556f
C742 VTAIL.n697 B 0.038119f
C743 VTAIL.n698 B 0.032168f
C744 VTAIL.n699 B 1.12497f
C745 VTAIL.n700 B 0.008472f
C746 VTAIL.n701 B 0.0191f
C747 VTAIL.n702 B 0.008556f
C748 VTAIL.n703 B 0.015038f
C749 VTAIL.n704 B 0.008081f
C750 VTAIL.n705 B 0.0191f
C751 VTAIL.n706 B 0.008556f
C752 VTAIL.n707 B 0.015038f
C753 VTAIL.n708 B 0.008081f
C754 VTAIL.n709 B 0.0191f
C755 VTAIL.n710 B 0.008556f
C756 VTAIL.n711 B 0.015038f
C757 VTAIL.n712 B 0.008081f
C758 VTAIL.n713 B 0.0191f
C759 VTAIL.n714 B 0.008556f
C760 VTAIL.n715 B 0.015038f
C761 VTAIL.n716 B 0.008081f
C762 VTAIL.n717 B 0.0191f
C763 VTAIL.n718 B 0.008556f
C764 VTAIL.n719 B 0.015038f
C765 VTAIL.n720 B 0.008081f
C766 VTAIL.n721 B 0.0191f
C767 VTAIL.n722 B 0.008556f
C768 VTAIL.n723 B 0.015038f
C769 VTAIL.n724 B 0.008081f
C770 VTAIL.n725 B 0.0191f
C771 VTAIL.n726 B 0.008556f
C772 VTAIL.n727 B 0.015038f
C773 VTAIL.n728 B 0.008081f
C774 VTAIL.n729 B 0.0191f
C775 VTAIL.n730 B 0.008556f
C776 VTAIL.n731 B 0.143409f
C777 VTAIL.t5 B 0.032749f
C778 VTAIL.n732 B 0.014325f
C779 VTAIL.n733 B 0.013502f
C780 VTAIL.n734 B 0.008081f
C781 VTAIL.n735 B 1.16398f
C782 VTAIL.n736 B 0.015038f
C783 VTAIL.n737 B 0.008081f
C784 VTAIL.n738 B 0.008556f
C785 VTAIL.n739 B 0.0191f
C786 VTAIL.n740 B 0.0191f
C787 VTAIL.n741 B 0.008556f
C788 VTAIL.n742 B 0.008081f
C789 VTAIL.n743 B 0.015038f
C790 VTAIL.n744 B 0.015038f
C791 VTAIL.n745 B 0.008081f
C792 VTAIL.n746 B 0.008556f
C793 VTAIL.n747 B 0.0191f
C794 VTAIL.n748 B 0.0191f
C795 VTAIL.n749 B 0.0191f
C796 VTAIL.n750 B 0.008556f
C797 VTAIL.n751 B 0.008081f
C798 VTAIL.n752 B 0.015038f
C799 VTAIL.n753 B 0.015038f
C800 VTAIL.n754 B 0.008081f
C801 VTAIL.n755 B 0.008318f
C802 VTAIL.n756 B 0.008318f
C803 VTAIL.n757 B 0.0191f
C804 VTAIL.n758 B 0.0191f
C805 VTAIL.n759 B 0.008556f
C806 VTAIL.n760 B 0.008081f
C807 VTAIL.n761 B 0.015038f
C808 VTAIL.n762 B 0.015038f
C809 VTAIL.n763 B 0.008081f
C810 VTAIL.n764 B 0.008556f
C811 VTAIL.n765 B 0.0191f
C812 VTAIL.n766 B 0.0191f
C813 VTAIL.n767 B 0.008556f
C814 VTAIL.n768 B 0.008081f
C815 VTAIL.n769 B 0.015038f
C816 VTAIL.n770 B 0.015038f
C817 VTAIL.n771 B 0.008081f
C818 VTAIL.n772 B 0.008556f
C819 VTAIL.n773 B 0.0191f
C820 VTAIL.n774 B 0.0191f
C821 VTAIL.n775 B 0.008556f
C822 VTAIL.n776 B 0.008081f
C823 VTAIL.n777 B 0.015038f
C824 VTAIL.n778 B 0.015038f
C825 VTAIL.n779 B 0.008081f
C826 VTAIL.n780 B 0.008556f
C827 VTAIL.n781 B 0.0191f
C828 VTAIL.n782 B 0.0191f
C829 VTAIL.n783 B 0.008556f
C830 VTAIL.n784 B 0.008081f
C831 VTAIL.n785 B 0.015038f
C832 VTAIL.n786 B 0.015038f
C833 VTAIL.n787 B 0.008081f
C834 VTAIL.n788 B 0.008556f
C835 VTAIL.n789 B 0.0191f
C836 VTAIL.n790 B 0.0191f
C837 VTAIL.n791 B 0.008556f
C838 VTAIL.n792 B 0.008081f
C839 VTAIL.n793 B 0.015038f
C840 VTAIL.n794 B 0.038457f
C841 VTAIL.n795 B 0.008081f
C842 VTAIL.n796 B 0.008556f
C843 VTAIL.n797 B 0.038119f
C844 VTAIL.n798 B 0.032168f
C845 VTAIL.n799 B 1.08414f
C846 VDD2.t2 B 0.378492f
C847 VDD2.t0 B 0.378492f
C848 VDD2.n0 B 4.26646f
C849 VDD2.t1 B 0.378492f
C850 VDD2.t3 B 0.378492f
C851 VDD2.n1 B 3.45869f
C852 VDD2.n2 B 4.1211f
C853 VN.t1 B 2.64375f
C854 VN.t2 B 2.64274f
C855 VN.n0 B 1.87533f
C856 VN.t3 B 2.64375f
C857 VN.t0 B 2.64274f
C858 VN.n1 B 3.38671f
.ends

