* NGSPICE file created from tg_sample_0010.ext - technology: sky130A

.subckt tg_sample_0010 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t33 VOUT.t32 VOUT.t33 VCC.t14 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X1 VSS.t18 VSS.t16 VSS.t17 VSS.t13 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=1.63
X2 VCC.t13 VCC.t11 VCC.t12 VCC.t8 sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=3.9
X3 VSS.t15 VSS.t12 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=1.63
X4 VOUT.t11 VGN.t0 VOUT.t10 VSS.t4 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=1.63
X5 VCC.t10 VCC.t7 VCC.t9 VCC.t8 sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=3.9
X6 VOUT.t2 VGN.t1 VOUT.t2 VSS.t2 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X7 VOUT.t31 VOUT.t29 VOUT.t30 VCC.t18 sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=3.9
X8 VOUT.t4 VGN.t2 VOUT.t4 VSS.t2 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X9 VOUT.t1 VGN.t3 VOUT.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X10 VSS.t11 VSS.t9 VSS.t10 VSS.t6 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=1.63
X11 VOUT.t28 VOUT.t27 VOUT.t28 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X12 VOUT.t3 VGN.t4 VOUT.t3 VSS.t3 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X13 VOUT.t26 VOUT.t24 VOUT.t25 VCC.t18 sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=3.9
X14 VOUT.t7 VGN.t5 VOUT.t7 VSS.t3 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X15 VOUT.t23 VOUT.t22 VOUT.t23 VCC.t16 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X16 VOUT.t21 VOUT.t20 VOUT.t21 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X17 VOUT.t19 VOUT.t18 VOUT.t19 VCC.t16 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X18 VOUT.t8 VGN.t6 VOUT.t8 VSS.t1 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X19 VSS.t8 VSS.t5 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=1.63
X20 VOUT.t9 VGN.t7 VOUT.t9 VSS.t0 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X21 VOUT.t17 VOUT.t16 VOUT.t17 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X22 VOUT.t0 VGN.t8 VOUT.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=2.7357 pd=16.91 as=0 ps=0 w=16.58 l=1.63
X23 VCC.t6 VCC.t4 VCC.t5 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=3.9
X24 VOUT.t15 VOUT.t14 VOUT.t15 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X25 VOUT.t13 VOUT.t12 VOUT.t13 VCC.t14 sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=0 ps=0 w=2.99 l=3.9
X26 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=3.9
X27 VOUT.t6 VGN.t9 VOUT.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=1.63
R0 VOUT.n15 VOUT.n12 161.3
R1 VOUT.n17 VOUT.n16 161.3
R2 VOUT.n18 VOUT.n11 161.3
R3 VOUT.n20 VOUT.n19 161.3
R4 VOUT.n21 VOUT.n10 161.3
R5 VOUT.n23 VOUT.n22 161.3
R6 VOUT.n24 VOUT.n9 161.3
R7 VOUT.n26 VOUT.n25 161.3
R8 VOUT.n27 VOUT.n8 161.3
R9 VOUT.n29 VOUT.n28 161.3
R10 VOUT.n30 VOUT.n7 161.3
R11 VOUT.n32 VOUT.n31 161.3
R12 VOUT.n33 VOUT.n6 161.3
R13 VOUT.n35 VOUT.n34 161.3
R14 VOUT.n36 VOUT.n5 161.3
R15 VOUT.n38 VOUT.n37 161.3
R16 VOUT.n39 VOUT.n4 161.3
R17 VOUT.n42 VOUT.n41 161.3
R18 VOUT.n43 VOUT.n3 161.3
R19 VOUT.n45 VOUT.n44 161.3
R20 VOUT.n46 VOUT.n2 161.3
R21 VOUT.n48 VOUT.n47 161.3
R22 VOUT.n49 VOUT.n1 161.3
R23 VOUT.n51 VOUT.n50 161.3
R24 VOUT.n52 VOUT.n0 161.3
R25 VOUT.n114 VOUT.n62 161.3
R26 VOUT.n113 VOUT.n112 161.3
R27 VOUT.n111 VOUT.n63 161.3
R28 VOUT.n110 VOUT.n109 161.3
R29 VOUT.n108 VOUT.n64 161.3
R30 VOUT.n107 VOUT.n106 161.3
R31 VOUT.n105 VOUT.n65 161.3
R32 VOUT.n104 VOUT.n103 161.3
R33 VOUT.n101 VOUT.n66 161.3
R34 VOUT.n100 VOUT.n99 161.3
R35 VOUT.n98 VOUT.n67 161.3
R36 VOUT.n97 VOUT.n96 161.3
R37 VOUT.n95 VOUT.n68 161.3
R38 VOUT.n94 VOUT.n93 161.3
R39 VOUT.n92 VOUT.n69 161.3
R40 VOUT.n91 VOUT.n90 161.3
R41 VOUT.n89 VOUT.n70 161.3
R42 VOUT.n88 VOUT.n87 161.3
R43 VOUT.n86 VOUT.n71 161.3
R44 VOUT.n85 VOUT.n84 161.3
R45 VOUT.n83 VOUT.n72 161.3
R46 VOUT.n82 VOUT.n81 161.3
R47 VOUT.n80 VOUT.n73 161.3
R48 VOUT.n79 VOUT.n78 161.3
R49 VOUT.n77 VOUT.n74 161.3
R50 VOUT.t17 VOUT.n61 157.048
R51 VOUT.n60 VOUT.t15 157.048
R52 VOUT.n125 VOUT.n124 142.53
R53 VOUT.n118 VOUT.n61 142.53
R54 VOUT.n128 VOUT.n127 142.53
R55 VOUT.n60 VOUT.n59 142.53
R56 VOUT.n121 VOUT.t31 136.722
R57 VOUT.n131 VOUT.t26 136.722
R58 VOUT.n130 VOUT.n58 129.499
R59 VOUT.n123 VOUT.n122 125.852
R60 VOUT.n120 VOUT.n119 125.852
R61 VOUT.n130 VOUT.n129 125.852
R62 VOUT.t8 VOUT.n133 66.3487
R63 VOUT.n146 VOUT.t1 66.3487
R64 VOUT.n14 VOUT.n13 63.8768
R65 VOUT.n76 VOUT.n75 63.8768
R66 VOUT.n141 VOUT.n140 63.4648
R67 VOUT.n134 VOUT.n133 63.4648
R68 VOUT.n145 VOUT.n144 63.4648
R69 VOUT.n147 VOUT.n146 63.4648
R70 VOUT.n54 VOUT.n53 59.6721
R71 VOUT.n116 VOUT.n115 59.6721
R72 VOUT.n47 VOUT.n46 55.548
R73 VOUT.n109 VOUT.n108 55.548
R74 VOUT.n34 VOUT.n33 51.663
R75 VOUT.n21 VOUT.n20 51.663
R76 VOUT.n83 VOUT.n82 51.663
R77 VOUT.n96 VOUT.n95 51.663
R78 VOUT.n75 VOUT.t29 50.6168
R79 VOUT.n13 VOUT.t24 50.6164
R80 VOUT.n138 VOUT.n135 48.4757
R81 VOUT.n136 VOUT.t6 47.9802
R82 VOUT.n137 VOUT.t11 47.9802
R83 VOUT.n143 VOUT.n56 46.786
R84 VOUT.n149 VOUT.n148 46.786
R85 VOUT.n139 VOUT.n138 46.786
R86 VOUT.n33 VOUT.n32 29.3238
R87 VOUT.n22 VOUT.n21 29.3238
R88 VOUT.n84 VOUT.n83 29.3238
R89 VOUT.n95 VOUT.n94 29.3238
R90 VOUT.n47 VOUT.n1 25.4388
R91 VOUT.n109 VOUT.n63 25.4388
R92 VOUT.n52 VOUT.n51 24.4675
R93 VOUT.n51 VOUT.n1 24.4675
R94 VOUT.n46 VOUT.n45 24.4675
R95 VOUT.n45 VOUT.n3 24.4675
R96 VOUT.n41 VOUT.n3 24.4675
R97 VOUT.n39 VOUT.n38 24.4675
R98 VOUT.n38 VOUT.n5 24.4675
R99 VOUT.n34 VOUT.n5 24.4675
R100 VOUT.n32 VOUT.n7 24.4675
R101 VOUT.n28 VOUT.n7 24.4675
R102 VOUT.n28 VOUT.n27 24.4675
R103 VOUT.n27 VOUT.n26 24.4675
R104 VOUT.n26 VOUT.n9 24.4675
R105 VOUT.n22 VOUT.n9 24.4675
R106 VOUT.n20 VOUT.n11 24.4675
R107 VOUT.n16 VOUT.n11 24.4675
R108 VOUT.n16 VOUT.n15 24.4675
R109 VOUT.n82 VOUT.n73 24.4675
R110 VOUT.n78 VOUT.n73 24.4675
R111 VOUT.n78 VOUT.n77 24.4675
R112 VOUT.n94 VOUT.n69 24.4675
R113 VOUT.n90 VOUT.n69 24.4675
R114 VOUT.n90 VOUT.n89 24.4675
R115 VOUT.n89 VOUT.n88 24.4675
R116 VOUT.n88 VOUT.n71 24.4675
R117 VOUT.n84 VOUT.n71 24.4675
R118 VOUT.n108 VOUT.n107 24.4675
R119 VOUT.n107 VOUT.n65 24.4675
R120 VOUT.n103 VOUT.n65 24.4675
R121 VOUT.n101 VOUT.n100 24.4675
R122 VOUT.n100 VOUT.n67 24.4675
R123 VOUT.n96 VOUT.n67 24.4675
R124 VOUT.n114 VOUT.n113 24.4675
R125 VOUT.n113 VOUT.n63 24.4675
R126 VOUT.n53 VOUT.n52 22.5101
R127 VOUT.n115 VOUT.n114 22.5101
R128 VIN VOUT.n55 18.841
R129 VOUT.n142 VOUT.n141 18.8065
R130 VOUT.n27 VOUT.t32 18.4772
R131 VOUT.n53 VOUT.t14 18.4772
R132 VOUT.n40 VOUT.t18 18.4772
R133 VOUT.n14 VOUT.t20 18.4772
R134 VOUT.n89 VOUT.t12 18.4772
R135 VOUT.n76 VOUT.t27 18.4772
R136 VOUT.n102 VOUT.t22 18.4772
R137 VOUT.n115 VOUT.t16 18.4772
R138 VOUT.n137 VOUT.n136 17.8281
R139 VOUT.n142 VOUT.n132 15.8865
R140 VOUT.n127 VOUT.n126 14.4315
R141 VOUT.n41 VOUT.n40 13.2127
R142 VOUT.n103 VOUT.n102 13.2127
R143 VOUT.n40 VOUT.n39 11.2553
R144 VOUT.n15 VOUT.n14 11.2553
R145 VOUT.n77 VOUT.n76 11.2553
R146 VOUT.n102 VOUT.n101 11.2553
R147 VOUT.n124 VOUT.t28 10.8717
R148 VOUT.n124 VOUT.t30 10.8717
R149 VOUT.t23 VOUT.n118 10.8717
R150 VOUT.n118 VOUT.t13 10.8717
R151 VOUT.n123 VOUT.t13 10.8717
R152 VOUT.t28 VOUT.n123 10.8717
R153 VOUT.n119 VOUT.t17 10.8717
R154 VOUT.n119 VOUT.t23 10.8717
R155 VOUT.n129 VOUT.t33 10.8717
R156 VOUT.n129 VOUT.t21 10.8717
R157 VOUT.t15 VOUT.n58 10.8717
R158 VOUT.t19 VOUT.n58 10.8717
R159 VOUT.t21 VOUT.n128 10.8717
R160 VOUT.n128 VOUT.t25 10.8717
R161 VOUT.n59 VOUT.t19 10.8717
R162 VOUT.n59 VOUT.t33 10.8717
R163 VOUT.n120 VOUT.n117 6.66429
R164 VOUT.n117 VGP 6.33817
R165 VOUT.n55 VOUT.n54 5.28823
R166 VOUT.n121 VOUT.n57 5.06539
R167 VOUT.n132 VOUT.n131 4.88412
R168 VOUT.n126 VOUT.n57 4.5005
R169 VOUT.n122 VOUT.n120 3.64705
R170 VOUT.n122 VOUT.n121 3.64705
R171 VOUT.n131 VOUT.n130 3.64705
R172 VOUT.n127 VOUT.n60 3.64705
R173 VOUT.n125 VOUT.n61 3.64705
R174 VOUT.n75 VOUT.n74 2.6058
R175 VOUT.n13 VOUT.n12 2.60578
R176 VOUT VOUT.n125 1.94447
R177 VOUT.n145 VOUT.n142 1.74619
R178 VOUT.n138 VOUT.n137 1.69016
R179 VOUT.n149 VOUT.n56 1.69016
R180 VOUT.n136 VOUT.n56 1.69016
R181 VOUT.n141 VOUT.n133 1.69016
R182 VOUT.n146 VOUT.n145 1.69016
R183 VOUT.n132 VOUT.n57 1.48273
R184 VOUT.n143 VOUT.t7 1.19471
R185 VOUT.t9 VOUT.n143 1.19471
R186 VOUT.n148 VOUT.t1 1.19471
R187 VOUT.n148 VOUT.t2 1.19471
R188 VOUT.n139 VOUT.t3 1.19471
R189 VOUT.t0 VOUT.n139 1.19471
R190 VOUT.n135 VOUT.t8 1.19471
R191 VOUT.n135 VOUT.t4 1.19471
R192 VOUT.n140 VOUT.t0 1.19471
R193 VOUT.n140 VOUT.t10 1.19471
R194 VOUT.t4 VOUT.n134 1.19471
R195 VOUT.n134 VOUT.t3 1.19471
R196 VOUT.n144 VOUT.t9 1.19471
R197 VOUT.n144 VOUT.t5 1.19471
R198 VOUT.t2 VOUT.n147 1.19471
R199 VOUT.n147 VOUT.t7 1.19471
R200 VIN VOUT.n149 0.849638
R201 VGP VOUT.n116 0.447322
R202 VOUT.n54 VOUT.n0 0.417535
R203 VOUT.n116 VOUT.n62 0.417535
R204 VOUT.n117 VOUT.n55 0.284154
R205 VOUT.n126 VOUT 0.220328
R206 VOUT.n50 VOUT.n0 0.189894
R207 VOUT.n50 VOUT.n49 0.189894
R208 VOUT.n49 VOUT.n48 0.189894
R209 VOUT.n48 VOUT.n2 0.189894
R210 VOUT.n44 VOUT.n2 0.189894
R211 VOUT.n44 VOUT.n43 0.189894
R212 VOUT.n43 VOUT.n42 0.189894
R213 VOUT.n42 VOUT.n4 0.189894
R214 VOUT.n37 VOUT.n4 0.189894
R215 VOUT.n37 VOUT.n36 0.189894
R216 VOUT.n36 VOUT.n35 0.189894
R217 VOUT.n35 VOUT.n6 0.189894
R218 VOUT.n31 VOUT.n6 0.189894
R219 VOUT.n31 VOUT.n30 0.189894
R220 VOUT.n30 VOUT.n29 0.189894
R221 VOUT.n29 VOUT.n8 0.189894
R222 VOUT.n25 VOUT.n8 0.189894
R223 VOUT.n25 VOUT.n24 0.189894
R224 VOUT.n24 VOUT.n23 0.189894
R225 VOUT.n23 VOUT.n10 0.189894
R226 VOUT.n19 VOUT.n10 0.189894
R227 VOUT.n19 VOUT.n18 0.189894
R228 VOUT.n18 VOUT.n17 0.189894
R229 VOUT.n17 VOUT.n12 0.189894
R230 VOUT.n112 VOUT.n62 0.189894
R231 VOUT.n112 VOUT.n111 0.189894
R232 VOUT.n111 VOUT.n110 0.189894
R233 VOUT.n110 VOUT.n64 0.189894
R234 VOUT.n106 VOUT.n64 0.189894
R235 VOUT.n106 VOUT.n105 0.189894
R236 VOUT.n105 VOUT.n104 0.189894
R237 VOUT.n104 VOUT.n66 0.189894
R238 VOUT.n99 VOUT.n66 0.189894
R239 VOUT.n99 VOUT.n98 0.189894
R240 VOUT.n98 VOUT.n97 0.189894
R241 VOUT.n97 VOUT.n68 0.189894
R242 VOUT.n93 VOUT.n68 0.189894
R243 VOUT.n93 VOUT.n92 0.189894
R244 VOUT.n92 VOUT.n91 0.189894
R245 VOUT.n91 VOUT.n70 0.189894
R246 VOUT.n87 VOUT.n70 0.189894
R247 VOUT.n87 VOUT.n86 0.189894
R248 VOUT.n86 VOUT.n85 0.189894
R249 VOUT.n85 VOUT.n72 0.189894
R250 VOUT.n81 VOUT.n72 0.189894
R251 VOUT.n81 VOUT.n80 0.189894
R252 VOUT.n80 VOUT.n79 0.189894
R253 VOUT.n79 VOUT.n74 0.189894
R254 VCC.n571 VCC.n44 367.317
R255 VCC.n569 VCC.n48 367.317
R256 VCC.n280 VCC.n197 367.317
R257 VCC.n282 VCC.n195 367.317
R258 VCC.n503 VCC.t11 227.897
R259 VCC.n493 VCC.t7 227.897
R260 VCC.n204 VCC.t0 227.897
R261 VCC.n214 VCC.t4 227.897
R262 VCC.n503 VCC.t12 227.101
R263 VCC.n493 VCC.t9 227.101
R264 VCC.n204 VCC.t3 227.101
R265 VCC.n214 VCC.t6 227.101
R266 VCC.n569 VCC.n568 185
R267 VCC.n570 VCC.n569 185
R268 VCC.n49 VCC.n47 185
R269 VCC.n47 VCC.n45 185
R270 VCC.n484 VCC.n483 185
R271 VCC.n483 VCC.n482 185
R272 VCC.n52 VCC.n51 185
R273 VCC.n481 VCC.n52 185
R274 VCC.n479 VCC.n478 185
R275 VCC.n480 VCC.n479 185
R276 VCC.n54 VCC.n53 185
R277 VCC.n471 VCC.n53 185
R278 VCC.n474 VCC.n473 185
R279 VCC.n473 VCC.n472 185
R280 VCC.n57 VCC.n56 185
R281 VCC.n469 VCC.n57 185
R282 VCC.n467 VCC.n466 185
R283 VCC.n468 VCC.n467 185
R284 VCC.n61 VCC.n60 185
R285 VCC.n60 VCC.n59 185
R286 VCC.n462 VCC.n461 185
R287 VCC.n461 VCC.n460 185
R288 VCC.n64 VCC.n63 185
R289 VCC.n459 VCC.n64 185
R290 VCC.n457 VCC.n456 185
R291 VCC.n458 VCC.n457 185
R292 VCC.n68 VCC.n67 185
R293 VCC.n67 VCC.n66 185
R294 VCC.n452 VCC.n451 185
R295 VCC.n451 VCC.n450 185
R296 VCC.n71 VCC.n70 185
R297 VCC.n449 VCC.n71 185
R298 VCC.n447 VCC.n446 185
R299 VCC.n448 VCC.n447 185
R300 VCC.n75 VCC.n74 185
R301 VCC.n74 VCC.n73 185
R302 VCC.n442 VCC.n441 185
R303 VCC.n441 VCC.n440 185
R304 VCC.n78 VCC.n77 185
R305 VCC.n439 VCC.n78 185
R306 VCC.n437 VCC.n436 185
R307 VCC.n438 VCC.n437 185
R308 VCC.n82 VCC.n81 185
R309 VCC.n81 VCC.n80 185
R310 VCC.n432 VCC.n431 185
R311 VCC.n431 VCC.n430 185
R312 VCC.n85 VCC.n84 185
R313 VCC.n429 VCC.n85 185
R314 VCC.n427 VCC.n426 185
R315 VCC.n428 VCC.n427 185
R316 VCC.n89 VCC.n88 185
R317 VCC.n88 VCC.n87 185
R318 VCC.n422 VCC.n421 185
R319 VCC.n421 VCC.n420 185
R320 VCC.n92 VCC.n91 185
R321 VCC.n419 VCC.n92 185
R322 VCC.n417 VCC.n416 185
R323 VCC.n418 VCC.n417 185
R324 VCC.n96 VCC.n95 185
R325 VCC.n95 VCC.n94 185
R326 VCC.n412 VCC.n411 185
R327 VCC.n411 VCC.n410 185
R328 VCC.n99 VCC.n98 185
R329 VCC.n409 VCC.n99 185
R330 VCC.n408 VCC.n407 185
R331 VCC.t14 VCC.n408 185
R332 VCC.n102 VCC.n101 185
R333 VCC.n101 VCC.n100 185
R334 VCC.n403 VCC.n402 185
R335 VCC.n402 VCC.n401 185
R336 VCC.n105 VCC.n104 185
R337 VCC.n106 VCC.n105 185
R338 VCC.n392 VCC.n391 185
R339 VCC.n393 VCC.n392 185
R340 VCC.n115 VCC.n114 185
R341 VCC.n114 VCC.n113 185
R342 VCC.n387 VCC.n386 185
R343 VCC.n386 VCC.n385 185
R344 VCC.n118 VCC.n117 185
R345 VCC.n119 VCC.n118 185
R346 VCC.n376 VCC.n375 185
R347 VCC.n377 VCC.n376 185
R348 VCC.n126 VCC.n125 185
R349 VCC.n131 VCC.n125 185
R350 VCC.n371 VCC.n370 185
R351 VCC.n370 VCC.n369 185
R352 VCC.n129 VCC.n128 185
R353 VCC.n130 VCC.n129 185
R354 VCC.n360 VCC.n359 185
R355 VCC.n361 VCC.n360 185
R356 VCC.n139 VCC.n138 185
R357 VCC.n138 VCC.n137 185
R358 VCC.n355 VCC.n354 185
R359 VCC.n354 VCC.n353 185
R360 VCC.n142 VCC.n141 185
R361 VCC.n143 VCC.n142 185
R362 VCC.n344 VCC.n343 185
R363 VCC.n345 VCC.n344 185
R364 VCC.n150 VCC.n149 185
R365 VCC.n155 VCC.n149 185
R366 VCC.n339 VCC.n338 185
R367 VCC.n338 VCC.n337 185
R368 VCC.n153 VCC.n152 185
R369 VCC.n154 VCC.n153 185
R370 VCC.n328 VCC.n327 185
R371 VCC.n329 VCC.n328 185
R372 VCC.n163 VCC.n162 185
R373 VCC.n162 VCC.n161 185
R374 VCC.n323 VCC.n322 185
R375 VCC.n322 VCC.n321 185
R376 VCC.n166 VCC.n165 185
R377 VCC.n167 VCC.n166 185
R378 VCC.n312 VCC.n311 185
R379 VCC.n313 VCC.n312 185
R380 VCC.n175 VCC.n174 185
R381 VCC.n174 VCC.n173 185
R382 VCC.n307 VCC.n306 185
R383 VCC.n306 VCC.n305 185
R384 VCC.n178 VCC.n177 185
R385 VCC.n179 VCC.n178 185
R386 VCC.n296 VCC.n295 185
R387 VCC.n297 VCC.n296 185
R388 VCC.n187 VCC.n186 185
R389 VCC.n186 VCC.n185 185
R390 VCC.n291 VCC.n290 185
R391 VCC.n290 VCC.n289 185
R392 VCC.n190 VCC.n189 185
R393 VCC.n191 VCC.n190 185
R394 VCC.n280 VCC.n279 185
R395 VCC.n281 VCC.n280 185
R396 VCC.n283 VCC.n282 185
R397 VCC.n282 VCC.n281 185
R398 VCC.n193 VCC.n192 185
R399 VCC.n192 VCC.n191 185
R400 VCC.n288 VCC.n287 185
R401 VCC.n289 VCC.n288 185
R402 VCC.n184 VCC.n183 185
R403 VCC.n185 VCC.n184 185
R404 VCC.n299 VCC.n298 185
R405 VCC.n298 VCC.n297 185
R406 VCC.n181 VCC.n180 185
R407 VCC.n180 VCC.n179 185
R408 VCC.n304 VCC.n303 185
R409 VCC.n305 VCC.n304 185
R410 VCC.n172 VCC.n171 185
R411 VCC.n173 VCC.n172 185
R412 VCC.n315 VCC.n314 185
R413 VCC.n314 VCC.n313 185
R414 VCC.n169 VCC.n168 185
R415 VCC.n168 VCC.n167 185
R416 VCC.n320 VCC.n319 185
R417 VCC.n321 VCC.n320 185
R418 VCC.n160 VCC.n159 185
R419 VCC.n161 VCC.n160 185
R420 VCC.n331 VCC.n330 185
R421 VCC.n330 VCC.n329 185
R422 VCC.n157 VCC.n156 185
R423 VCC.n156 VCC.n154 185
R424 VCC.n336 VCC.n335 185
R425 VCC.n337 VCC.n336 185
R426 VCC.n148 VCC.n147 185
R427 VCC.n155 VCC.n148 185
R428 VCC.n347 VCC.n346 185
R429 VCC.n346 VCC.n345 185
R430 VCC.n145 VCC.n144 185
R431 VCC.n144 VCC.n143 185
R432 VCC.n352 VCC.n351 185
R433 VCC.n353 VCC.n352 185
R434 VCC.n136 VCC.n135 185
R435 VCC.n137 VCC.n136 185
R436 VCC.n363 VCC.n362 185
R437 VCC.n362 VCC.n361 185
R438 VCC.n133 VCC.n132 185
R439 VCC.n132 VCC.n130 185
R440 VCC.n368 VCC.n367 185
R441 VCC.n369 VCC.n368 185
R442 VCC.n124 VCC.n123 185
R443 VCC.n131 VCC.n124 185
R444 VCC.n379 VCC.n378 185
R445 VCC.n378 VCC.n377 185
R446 VCC.n121 VCC.n120 185
R447 VCC.n120 VCC.n119 185
R448 VCC.n384 VCC.n383 185
R449 VCC.n385 VCC.n384 185
R450 VCC.n112 VCC.n111 185
R451 VCC.n113 VCC.n112 185
R452 VCC.n395 VCC.n394 185
R453 VCC.n394 VCC.n393 185
R454 VCC.n109 VCC.n107 185
R455 VCC.n107 VCC.n106 185
R456 VCC.n400 VCC.n399 185
R457 VCC.n401 VCC.n400 185
R458 VCC.n108 VCC.n2 185
R459 VCC.n108 VCC.n100 185
R460 VCC.n620 VCC.n3 185
R461 VCC.t14 VCC.n3 185
R462 VCC.n619 VCC.n4 185
R463 VCC.n409 VCC.n4 185
R464 VCC.n618 VCC.n5 185
R465 VCC.n410 VCC.n5 185
R466 VCC.n93 VCC.n6 185
R467 VCC.n94 VCC.n93 185
R468 VCC.n614 VCC.n8 185
R469 VCC.n418 VCC.n8 185
R470 VCC.n613 VCC.n9 185
R471 VCC.n419 VCC.n9 185
R472 VCC.n612 VCC.n10 185
R473 VCC.n420 VCC.n10 185
R474 VCC.n86 VCC.n11 185
R475 VCC.n87 VCC.n86 185
R476 VCC.n608 VCC.n13 185
R477 VCC.n428 VCC.n13 185
R478 VCC.n607 VCC.n14 185
R479 VCC.n429 VCC.n14 185
R480 VCC.n606 VCC.n15 185
R481 VCC.n430 VCC.n15 185
R482 VCC.n79 VCC.n16 185
R483 VCC.n80 VCC.n79 185
R484 VCC.n602 VCC.n18 185
R485 VCC.n438 VCC.n18 185
R486 VCC.n601 VCC.n19 185
R487 VCC.n439 VCC.n19 185
R488 VCC.n600 VCC.n20 185
R489 VCC.n440 VCC.n20 185
R490 VCC.n72 VCC.n21 185
R491 VCC.n73 VCC.n72 185
R492 VCC.n596 VCC.n23 185
R493 VCC.n448 VCC.n23 185
R494 VCC.n595 VCC.n24 185
R495 VCC.n449 VCC.n24 185
R496 VCC.n594 VCC.n25 185
R497 VCC.n450 VCC.n25 185
R498 VCC.n65 VCC.n26 185
R499 VCC.n66 VCC.n65 185
R500 VCC.n590 VCC.n28 185
R501 VCC.n458 VCC.n28 185
R502 VCC.n589 VCC.n29 185
R503 VCC.n459 VCC.n29 185
R504 VCC.n588 VCC.n30 185
R505 VCC.n460 VCC.n30 185
R506 VCC.n58 VCC.n31 185
R507 VCC.n59 VCC.n58 185
R508 VCC.n584 VCC.n33 185
R509 VCC.n468 VCC.n33 185
R510 VCC.n583 VCC.n34 185
R511 VCC.n469 VCC.n34 185
R512 VCC.n582 VCC.n35 185
R513 VCC.n472 VCC.n35 185
R514 VCC.n470 VCC.n36 185
R515 VCC.n471 VCC.n470 185
R516 VCC.n578 VCC.n38 185
R517 VCC.n480 VCC.n38 185
R518 VCC.n577 VCC.n39 185
R519 VCC.n481 VCC.n39 185
R520 VCC.n576 VCC.n40 185
R521 VCC.n482 VCC.n40 185
R522 VCC.n43 VCC.n41 185
R523 VCC.n45 VCC.n43 185
R524 VCC.n572 VCC.n571 185
R525 VCC.n571 VCC.n570 185
R526 VCC.n566 VCC.n48 185
R527 VCC.n565 VCC.n564 185
R528 VCC.n562 VCC.n487 185
R529 VCC.n560 VCC.n559 185
R530 VCC.n558 VCC.n488 185
R531 VCC.n557 VCC.n556 185
R532 VCC.n554 VCC.n489 185
R533 VCC.n552 VCC.n551 185
R534 VCC.n550 VCC.n490 185
R535 VCC.n549 VCC.n548 185
R536 VCC.n546 VCC.n491 185
R537 VCC.n544 VCC.n543 185
R538 VCC.n542 VCC.n492 185
R539 VCC.n540 VCC.n539 185
R540 VCC.n537 VCC.n495 185
R541 VCC.n535 VCC.n534 185
R542 VCC.n533 VCC.n496 185
R543 VCC.n532 VCC.n531 185
R544 VCC.n529 VCC.n497 185
R545 VCC.n527 VCC.n526 185
R546 VCC.n525 VCC.n498 185
R547 VCC.n524 VCC.n523 185
R548 VCC.n521 VCC.n499 185
R549 VCC.n519 VCC.n518 185
R550 VCC.n517 VCC.n500 185
R551 VCC.n516 VCC.n515 185
R552 VCC.n513 VCC.n501 185
R553 VCC.n511 VCC.n510 185
R554 VCC.n509 VCC.n502 185
R555 VCC.n507 VCC.n506 185
R556 VCC.n44 VCC.n42 185
R557 VCC.n46 VCC.n44 185
R558 VCC.n195 VCC.n194 185
R559 VCC.n218 VCC.n217 185
R560 VCC.n220 VCC.n213 185
R561 VCC.n213 VCC.n196 185
R562 VCC.n222 VCC.n221 185
R563 VCC.n224 VCC.n212 185
R564 VCC.n227 VCC.n226 185
R565 VCC.n228 VCC.n211 185
R566 VCC.n230 VCC.n229 185
R567 VCC.n232 VCC.n210 185
R568 VCC.n235 VCC.n234 185
R569 VCC.n236 VCC.n209 185
R570 VCC.n238 VCC.n237 185
R571 VCC.n240 VCC.n208 185
R572 VCC.n243 VCC.n242 185
R573 VCC.n244 VCC.n207 185
R574 VCC.n246 VCC.n245 185
R575 VCC.n248 VCC.n206 185
R576 VCC.n251 VCC.n250 185
R577 VCC.n253 VCC.n203 185
R578 VCC.n255 VCC.n254 185
R579 VCC.n257 VCC.n202 185
R580 VCC.n260 VCC.n259 185
R581 VCC.n261 VCC.n201 185
R582 VCC.n263 VCC.n262 185
R583 VCC.n265 VCC.n200 185
R584 VCC.n268 VCC.n267 185
R585 VCC.n269 VCC.n199 185
R586 VCC.n271 VCC.n270 185
R587 VCC.n273 VCC.n198 185
R588 VCC.n276 VCC.n275 185
R589 VCC.n277 VCC.n197 185
R590 VCC.n280 VCC.n190 146.341
R591 VCC.n290 VCC.n190 146.341
R592 VCC.n290 VCC.n186 146.341
R593 VCC.n296 VCC.n186 146.341
R594 VCC.n296 VCC.n178 146.341
R595 VCC.n306 VCC.n178 146.341
R596 VCC.n306 VCC.n174 146.341
R597 VCC.n312 VCC.n174 146.341
R598 VCC.n312 VCC.n166 146.341
R599 VCC.n322 VCC.n166 146.341
R600 VCC.n322 VCC.n162 146.341
R601 VCC.n328 VCC.n162 146.341
R602 VCC.n328 VCC.n153 146.341
R603 VCC.n338 VCC.n153 146.341
R604 VCC.n338 VCC.n149 146.341
R605 VCC.n344 VCC.n149 146.341
R606 VCC.n344 VCC.n142 146.341
R607 VCC.n354 VCC.n142 146.341
R608 VCC.n354 VCC.n138 146.341
R609 VCC.n360 VCC.n138 146.341
R610 VCC.n360 VCC.n129 146.341
R611 VCC.n370 VCC.n129 146.341
R612 VCC.n370 VCC.n125 146.341
R613 VCC.n376 VCC.n125 146.341
R614 VCC.n376 VCC.n118 146.341
R615 VCC.n386 VCC.n118 146.341
R616 VCC.n386 VCC.n114 146.341
R617 VCC.n392 VCC.n114 146.341
R618 VCC.n392 VCC.n105 146.341
R619 VCC.n402 VCC.n105 146.341
R620 VCC.n402 VCC.n101 146.341
R621 VCC.n408 VCC.n101 146.341
R622 VCC.n408 VCC.n99 146.341
R623 VCC.n411 VCC.n99 146.341
R624 VCC.n411 VCC.n95 146.341
R625 VCC.n417 VCC.n95 146.341
R626 VCC.n417 VCC.n92 146.341
R627 VCC.n421 VCC.n92 146.341
R628 VCC.n421 VCC.n88 146.341
R629 VCC.n427 VCC.n88 146.341
R630 VCC.n427 VCC.n85 146.341
R631 VCC.n431 VCC.n85 146.341
R632 VCC.n431 VCC.n81 146.341
R633 VCC.n437 VCC.n81 146.341
R634 VCC.n437 VCC.n78 146.341
R635 VCC.n441 VCC.n78 146.341
R636 VCC.n441 VCC.n74 146.341
R637 VCC.n447 VCC.n74 146.341
R638 VCC.n447 VCC.n71 146.341
R639 VCC.n451 VCC.n71 146.341
R640 VCC.n451 VCC.n67 146.341
R641 VCC.n457 VCC.n67 146.341
R642 VCC.n457 VCC.n64 146.341
R643 VCC.n461 VCC.n64 146.341
R644 VCC.n461 VCC.n60 146.341
R645 VCC.n467 VCC.n60 146.341
R646 VCC.n467 VCC.n57 146.341
R647 VCC.n473 VCC.n57 146.341
R648 VCC.n473 VCC.n53 146.341
R649 VCC.n479 VCC.n53 146.341
R650 VCC.n479 VCC.n52 146.341
R651 VCC.n483 VCC.n52 146.341
R652 VCC.n483 VCC.n47 146.341
R653 VCC.n569 VCC.n47 146.341
R654 VCC.n282 VCC.n192 146.341
R655 VCC.n288 VCC.n192 146.341
R656 VCC.n288 VCC.n184 146.341
R657 VCC.n298 VCC.n184 146.341
R658 VCC.n298 VCC.n180 146.341
R659 VCC.n304 VCC.n180 146.341
R660 VCC.n304 VCC.n172 146.341
R661 VCC.n314 VCC.n172 146.341
R662 VCC.n314 VCC.n168 146.341
R663 VCC.n320 VCC.n168 146.341
R664 VCC.n320 VCC.n160 146.341
R665 VCC.n330 VCC.n160 146.341
R666 VCC.n330 VCC.n156 146.341
R667 VCC.n336 VCC.n156 146.341
R668 VCC.n336 VCC.n148 146.341
R669 VCC.n346 VCC.n148 146.341
R670 VCC.n346 VCC.n144 146.341
R671 VCC.n352 VCC.n144 146.341
R672 VCC.n352 VCC.n136 146.341
R673 VCC.n362 VCC.n136 146.341
R674 VCC.n362 VCC.n132 146.341
R675 VCC.n368 VCC.n132 146.341
R676 VCC.n368 VCC.n124 146.341
R677 VCC.n378 VCC.n124 146.341
R678 VCC.n378 VCC.n120 146.341
R679 VCC.n384 VCC.n120 146.341
R680 VCC.n384 VCC.n112 146.341
R681 VCC.n394 VCC.n112 146.341
R682 VCC.n394 VCC.n107 146.341
R683 VCC.n400 VCC.n107 146.341
R684 VCC.n400 VCC.n108 146.341
R685 VCC.n108 VCC.n3 146.341
R686 VCC.n4 VCC.n3 146.341
R687 VCC.n5 VCC.n4 146.341
R688 VCC.n93 VCC.n5 146.341
R689 VCC.n93 VCC.n8 146.341
R690 VCC.n9 VCC.n8 146.341
R691 VCC.n10 VCC.n9 146.341
R692 VCC.n86 VCC.n10 146.341
R693 VCC.n86 VCC.n13 146.341
R694 VCC.n14 VCC.n13 146.341
R695 VCC.n15 VCC.n14 146.341
R696 VCC.n79 VCC.n15 146.341
R697 VCC.n79 VCC.n18 146.341
R698 VCC.n19 VCC.n18 146.341
R699 VCC.n20 VCC.n19 146.341
R700 VCC.n72 VCC.n20 146.341
R701 VCC.n72 VCC.n23 146.341
R702 VCC.n24 VCC.n23 146.341
R703 VCC.n25 VCC.n24 146.341
R704 VCC.n65 VCC.n25 146.341
R705 VCC.n65 VCC.n28 146.341
R706 VCC.n29 VCC.n28 146.341
R707 VCC.n30 VCC.n29 146.341
R708 VCC.n58 VCC.n30 146.341
R709 VCC.n58 VCC.n33 146.341
R710 VCC.n34 VCC.n33 146.341
R711 VCC.n35 VCC.n34 146.341
R712 VCC.n470 VCC.n35 146.341
R713 VCC.n470 VCC.n38 146.341
R714 VCC.n39 VCC.n38 146.341
R715 VCC.n40 VCC.n39 146.341
R716 VCC.n43 VCC.n40 146.341
R717 VCC.n571 VCC.n43 146.341
R718 VCC.n504 VCC.t13 145.065
R719 VCC.n494 VCC.t10 145.065
R720 VCC.n205 VCC.t2 145.065
R721 VCC.n215 VCC.t5 145.065
R722 VCC.n506 VCC.n44 99.5127
R723 VCC.n511 VCC.n502 99.5127
R724 VCC.n515 VCC.n513 99.5127
R725 VCC.n519 VCC.n500 99.5127
R726 VCC.n523 VCC.n521 99.5127
R727 VCC.n527 VCC.n498 99.5127
R728 VCC.n531 VCC.n529 99.5127
R729 VCC.n535 VCC.n496 99.5127
R730 VCC.n539 VCC.n537 99.5127
R731 VCC.n544 VCC.n492 99.5127
R732 VCC.n548 VCC.n546 99.5127
R733 VCC.n552 VCC.n490 99.5127
R734 VCC.n556 VCC.n554 99.5127
R735 VCC.n560 VCC.n488 99.5127
R736 VCC.n564 VCC.n562 99.5127
R737 VCC.n217 VCC.n213 99.5127
R738 VCC.n222 VCC.n213 99.5127
R739 VCC.n226 VCC.n224 99.5127
R740 VCC.n230 VCC.n211 99.5127
R741 VCC.n234 VCC.n232 99.5127
R742 VCC.n238 VCC.n209 99.5127
R743 VCC.n242 VCC.n240 99.5127
R744 VCC.n246 VCC.n207 99.5127
R745 VCC.n250 VCC.n248 99.5127
R746 VCC.n255 VCC.n203 99.5127
R747 VCC.n259 VCC.n257 99.5127
R748 VCC.n263 VCC.n201 99.5127
R749 VCC.n267 VCC.n265 99.5127
R750 VCC.n271 VCC.n199 99.5127
R751 VCC.n275 VCC.n273 99.5127
R752 VCC.n504 VCC.n503 82.0369
R753 VCC.n494 VCC.n493 82.0369
R754 VCC.n205 VCC.n204 82.0369
R755 VCC.n215 VCC.n214 82.0369
R756 VCC.n563 VCC.n46 72.8958
R757 VCC.n561 VCC.n46 72.8958
R758 VCC.n555 VCC.n46 72.8958
R759 VCC.n553 VCC.n46 72.8958
R760 VCC.n547 VCC.n46 72.8958
R761 VCC.n545 VCC.n46 72.8958
R762 VCC.n538 VCC.n46 72.8958
R763 VCC.n536 VCC.n46 72.8958
R764 VCC.n530 VCC.n46 72.8958
R765 VCC.n528 VCC.n46 72.8958
R766 VCC.n522 VCC.n46 72.8958
R767 VCC.n520 VCC.n46 72.8958
R768 VCC.n514 VCC.n46 72.8958
R769 VCC.n512 VCC.n46 72.8958
R770 VCC.n505 VCC.n46 72.8958
R771 VCC.n216 VCC.n196 72.8958
R772 VCC.n223 VCC.n196 72.8958
R773 VCC.n225 VCC.n196 72.8958
R774 VCC.n231 VCC.n196 72.8958
R775 VCC.n233 VCC.n196 72.8958
R776 VCC.n239 VCC.n196 72.8958
R777 VCC.n241 VCC.n196 72.8958
R778 VCC.n247 VCC.n196 72.8958
R779 VCC.n249 VCC.n196 72.8958
R780 VCC.n256 VCC.n196 72.8958
R781 VCC.n258 VCC.n196 72.8958
R782 VCC.n264 VCC.n196 72.8958
R783 VCC.n266 VCC.n196 72.8958
R784 VCC.n272 VCC.n196 72.8958
R785 VCC.n274 VCC.n196 72.8958
R786 VCC.n281 VCC.n196 65.2939
R787 VCC.n570 VCC.n46 65.2939
R788 VCC.n505 VCC.n502 39.2114
R789 VCC.n513 VCC.n512 39.2114
R790 VCC.n514 VCC.n500 39.2114
R791 VCC.n521 VCC.n520 39.2114
R792 VCC.n522 VCC.n498 39.2114
R793 VCC.n529 VCC.n528 39.2114
R794 VCC.n530 VCC.n496 39.2114
R795 VCC.n537 VCC.n536 39.2114
R796 VCC.n538 VCC.n492 39.2114
R797 VCC.n546 VCC.n545 39.2114
R798 VCC.n547 VCC.n490 39.2114
R799 VCC.n554 VCC.n553 39.2114
R800 VCC.n555 VCC.n488 39.2114
R801 VCC.n562 VCC.n561 39.2114
R802 VCC.n563 VCC.n48 39.2114
R803 VCC.n216 VCC.n195 39.2114
R804 VCC.n223 VCC.n222 39.2114
R805 VCC.n226 VCC.n225 39.2114
R806 VCC.n231 VCC.n230 39.2114
R807 VCC.n234 VCC.n233 39.2114
R808 VCC.n239 VCC.n238 39.2114
R809 VCC.n242 VCC.n241 39.2114
R810 VCC.n247 VCC.n246 39.2114
R811 VCC.n250 VCC.n249 39.2114
R812 VCC.n256 VCC.n255 39.2114
R813 VCC.n259 VCC.n258 39.2114
R814 VCC.n264 VCC.n263 39.2114
R815 VCC.n267 VCC.n266 39.2114
R816 VCC.n272 VCC.n271 39.2114
R817 VCC.n275 VCC.n274 39.2114
R818 VCC.n564 VCC.n563 39.2114
R819 VCC.n561 VCC.n560 39.2114
R820 VCC.n556 VCC.n555 39.2114
R821 VCC.n553 VCC.n552 39.2114
R822 VCC.n548 VCC.n547 39.2114
R823 VCC.n545 VCC.n544 39.2114
R824 VCC.n539 VCC.n538 39.2114
R825 VCC.n536 VCC.n535 39.2114
R826 VCC.n531 VCC.n530 39.2114
R827 VCC.n528 VCC.n527 39.2114
R828 VCC.n523 VCC.n522 39.2114
R829 VCC.n520 VCC.n519 39.2114
R830 VCC.n515 VCC.n514 39.2114
R831 VCC.n512 VCC.n511 39.2114
R832 VCC.n506 VCC.n505 39.2114
R833 VCC.n217 VCC.n216 39.2114
R834 VCC.n224 VCC.n223 39.2114
R835 VCC.n225 VCC.n211 39.2114
R836 VCC.n232 VCC.n231 39.2114
R837 VCC.n233 VCC.n209 39.2114
R838 VCC.n240 VCC.n239 39.2114
R839 VCC.n241 VCC.n207 39.2114
R840 VCC.n248 VCC.n247 39.2114
R841 VCC.n249 VCC.n203 39.2114
R842 VCC.n257 VCC.n256 39.2114
R843 VCC.n258 VCC.n201 39.2114
R844 VCC.n265 VCC.n264 39.2114
R845 VCC.n266 VCC.n199 39.2114
R846 VCC.n273 VCC.n272 39.2114
R847 VCC.n274 VCC.n197 39.2114
R848 VCC.n281 VCC.n191 38.1838
R849 VCC.n289 VCC.n191 38.1838
R850 VCC.n289 VCC.n185 38.1838
R851 VCC.n297 VCC.n185 38.1838
R852 VCC.n305 VCC.n179 38.1838
R853 VCC.n305 VCC.n173 38.1838
R854 VCC.n313 VCC.n173 38.1838
R855 VCC.n313 VCC.n167 38.1838
R856 VCC.n321 VCC.n167 38.1838
R857 VCC.n321 VCC.n161 38.1838
R858 VCC.n329 VCC.n161 38.1838
R859 VCC.n329 VCC.n154 38.1838
R860 VCC.n337 VCC.n154 38.1838
R861 VCC.n337 VCC.n155 38.1838
R862 VCC.n345 VCC.n143 38.1838
R863 VCC.n353 VCC.n143 38.1838
R864 VCC.n353 VCC.n137 38.1838
R865 VCC.n361 VCC.n137 38.1838
R866 VCC.n361 VCC.n130 38.1838
R867 VCC.n369 VCC.n130 38.1838
R868 VCC.n369 VCC.n131 38.1838
R869 VCC.n377 VCC.n119 38.1838
R870 VCC.n385 VCC.n119 38.1838
R871 VCC.n385 VCC.n113 38.1838
R872 VCC.n393 VCC.n113 38.1838
R873 VCC.n393 VCC.n106 38.1838
R874 VCC.n401 VCC.n106 38.1838
R875 VCC.n401 VCC.n100 38.1838
R876 VCC.t14 VCC.n100 38.1838
R877 VCC.n409 VCC.t14 38.1838
R878 VCC.n410 VCC.n409 38.1838
R879 VCC.n410 VCC.n94 38.1838
R880 VCC.n418 VCC.n94 38.1838
R881 VCC.n419 VCC.n418 38.1838
R882 VCC.n420 VCC.n419 38.1838
R883 VCC.n420 VCC.n87 38.1838
R884 VCC.n428 VCC.n87 38.1838
R885 VCC.n430 VCC.n429 38.1838
R886 VCC.n430 VCC.n80 38.1838
R887 VCC.n438 VCC.n80 38.1838
R888 VCC.n439 VCC.n438 38.1838
R889 VCC.n440 VCC.n439 38.1838
R890 VCC.n440 VCC.n73 38.1838
R891 VCC.n448 VCC.n73 38.1838
R892 VCC.n450 VCC.n449 38.1838
R893 VCC.n450 VCC.n66 38.1838
R894 VCC.n458 VCC.n66 38.1838
R895 VCC.n459 VCC.n458 38.1838
R896 VCC.n460 VCC.n459 38.1838
R897 VCC.n460 VCC.n59 38.1838
R898 VCC.n468 VCC.n59 38.1838
R899 VCC.n469 VCC.n468 38.1838
R900 VCC.n472 VCC.n469 38.1838
R901 VCC.n472 VCC.n471 38.1838
R902 VCC.n481 VCC.n480 38.1838
R903 VCC.n482 VCC.n481 38.1838
R904 VCC.n482 VCC.n45 38.1838
R905 VCC.n570 VCC.n45 38.1838
R906 VCC.n345 VCC.t15 35.1291
R907 VCC.t18 VCC.n448 35.1291
R908 VCC.n508 VCC.n504 29.2853
R909 VCC.n541 VCC.n494 29.2853
R910 VCC.n252 VCC.n205 29.2853
R911 VCC.n219 VCC.n215 29.2853
R912 VCC.n573 VCC.n42 28.449
R913 VCC.n567 VCC.n566 28.449
R914 VCC.n284 VCC.n194 28.449
R915 VCC.n278 VCC.n277 28.449
R916 VCC.t1 VCC.n179 21.3831
R917 VCC.n471 VCC.t8 21.3831
R918 VCC.n131 VCC.t16 20.6195
R919 VCC.n429 VCC.t17 20.6195
R920 VCC.n279 VCC.n189 19.3944
R921 VCC.n291 VCC.n189 19.3944
R922 VCC.n291 VCC.n187 19.3944
R923 VCC.n295 VCC.n187 19.3944
R924 VCC.n295 VCC.n177 19.3944
R925 VCC.n307 VCC.n177 19.3944
R926 VCC.n307 VCC.n175 19.3944
R927 VCC.n311 VCC.n175 19.3944
R928 VCC.n311 VCC.n165 19.3944
R929 VCC.n323 VCC.n165 19.3944
R930 VCC.n323 VCC.n163 19.3944
R931 VCC.n327 VCC.n163 19.3944
R932 VCC.n327 VCC.n152 19.3944
R933 VCC.n339 VCC.n152 19.3944
R934 VCC.n339 VCC.n150 19.3944
R935 VCC.n343 VCC.n150 19.3944
R936 VCC.n343 VCC.n141 19.3944
R937 VCC.n355 VCC.n141 19.3944
R938 VCC.n355 VCC.n139 19.3944
R939 VCC.n359 VCC.n139 19.3944
R940 VCC.n359 VCC.n128 19.3944
R941 VCC.n371 VCC.n128 19.3944
R942 VCC.n371 VCC.n126 19.3944
R943 VCC.n375 VCC.n126 19.3944
R944 VCC.n375 VCC.n117 19.3944
R945 VCC.n387 VCC.n117 19.3944
R946 VCC.n387 VCC.n115 19.3944
R947 VCC.n391 VCC.n115 19.3944
R948 VCC.n391 VCC.n104 19.3944
R949 VCC.n403 VCC.n104 19.3944
R950 VCC.n403 VCC.n102 19.3944
R951 VCC.n407 VCC.n102 19.3944
R952 VCC.n407 VCC.n98 19.3944
R953 VCC.n412 VCC.n98 19.3944
R954 VCC.n412 VCC.n96 19.3944
R955 VCC.n416 VCC.n96 19.3944
R956 VCC.n416 VCC.n91 19.3944
R957 VCC.n422 VCC.n91 19.3944
R958 VCC.n422 VCC.n89 19.3944
R959 VCC.n426 VCC.n89 19.3944
R960 VCC.n426 VCC.n84 19.3944
R961 VCC.n432 VCC.n84 19.3944
R962 VCC.n432 VCC.n82 19.3944
R963 VCC.n436 VCC.n82 19.3944
R964 VCC.n436 VCC.n77 19.3944
R965 VCC.n442 VCC.n77 19.3944
R966 VCC.n442 VCC.n75 19.3944
R967 VCC.n446 VCC.n75 19.3944
R968 VCC.n446 VCC.n70 19.3944
R969 VCC.n452 VCC.n70 19.3944
R970 VCC.n452 VCC.n68 19.3944
R971 VCC.n456 VCC.n68 19.3944
R972 VCC.n456 VCC.n63 19.3944
R973 VCC.n462 VCC.n63 19.3944
R974 VCC.n462 VCC.n61 19.3944
R975 VCC.n466 VCC.n61 19.3944
R976 VCC.n466 VCC.n56 19.3944
R977 VCC.n474 VCC.n56 19.3944
R978 VCC.n474 VCC.n54 19.3944
R979 VCC.n478 VCC.n54 19.3944
R980 VCC.n478 VCC.n51 19.3944
R981 VCC.n484 VCC.n51 19.3944
R982 VCC.n484 VCC.n49 19.3944
R983 VCC.n568 VCC.n49 19.3944
R984 VCC.n283 VCC.n193 19.3944
R985 VCC.n287 VCC.n193 19.3944
R986 VCC.n287 VCC.n183 19.3944
R987 VCC.n299 VCC.n183 19.3944
R988 VCC.n299 VCC.n181 19.3944
R989 VCC.n303 VCC.n181 19.3944
R990 VCC.n303 VCC.n171 19.3944
R991 VCC.n315 VCC.n171 19.3944
R992 VCC.n315 VCC.n169 19.3944
R993 VCC.n319 VCC.n169 19.3944
R994 VCC.n319 VCC.n159 19.3944
R995 VCC.n331 VCC.n159 19.3944
R996 VCC.n331 VCC.n157 19.3944
R997 VCC.n335 VCC.n157 19.3944
R998 VCC.n335 VCC.n147 19.3944
R999 VCC.n347 VCC.n147 19.3944
R1000 VCC.n347 VCC.n145 19.3944
R1001 VCC.n351 VCC.n145 19.3944
R1002 VCC.n351 VCC.n135 19.3944
R1003 VCC.n363 VCC.n135 19.3944
R1004 VCC.n363 VCC.n133 19.3944
R1005 VCC.n367 VCC.n133 19.3944
R1006 VCC.n367 VCC.n123 19.3944
R1007 VCC.n379 VCC.n123 19.3944
R1008 VCC.n379 VCC.n121 19.3944
R1009 VCC.n383 VCC.n121 19.3944
R1010 VCC.n383 VCC.n111 19.3944
R1011 VCC.n395 VCC.n111 19.3944
R1012 VCC.n395 VCC.n109 19.3944
R1013 VCC.n399 VCC.n109 19.3944
R1014 VCC.n399 VCC.n2 19.3944
R1015 VCC.n620 VCC.n2 19.3944
R1016 VCC.n620 VCC.n619 19.3944
R1017 VCC.n619 VCC.n618 19.3944
R1018 VCC.n618 VCC.n6 19.3944
R1019 VCC.n614 VCC.n6 19.3944
R1020 VCC.n614 VCC.n613 19.3944
R1021 VCC.n613 VCC.n612 19.3944
R1022 VCC.n612 VCC.n11 19.3944
R1023 VCC.n608 VCC.n11 19.3944
R1024 VCC.n608 VCC.n607 19.3944
R1025 VCC.n607 VCC.n606 19.3944
R1026 VCC.n606 VCC.n16 19.3944
R1027 VCC.n602 VCC.n16 19.3944
R1028 VCC.n602 VCC.n601 19.3944
R1029 VCC.n601 VCC.n600 19.3944
R1030 VCC.n600 VCC.n21 19.3944
R1031 VCC.n596 VCC.n21 19.3944
R1032 VCC.n596 VCC.n595 19.3944
R1033 VCC.n595 VCC.n594 19.3944
R1034 VCC.n594 VCC.n26 19.3944
R1035 VCC.n590 VCC.n26 19.3944
R1036 VCC.n590 VCC.n589 19.3944
R1037 VCC.n589 VCC.n588 19.3944
R1038 VCC.n588 VCC.n31 19.3944
R1039 VCC.n584 VCC.n31 19.3944
R1040 VCC.n584 VCC.n583 19.3944
R1041 VCC.n583 VCC.n582 19.3944
R1042 VCC.n582 VCC.n36 19.3944
R1043 VCC.n578 VCC.n36 19.3944
R1044 VCC.n578 VCC.n577 19.3944
R1045 VCC.n577 VCC.n576 19.3944
R1046 VCC.n576 VCC.n41 19.3944
R1047 VCC.n572 VCC.n41 19.3944
R1048 VCC.n377 VCC.t16 17.5648
R1049 VCC.t17 VCC.n428 17.5648
R1050 VCC.n297 VCC.t1 16.8011
R1051 VCC.n480 VCC.t8 16.8011
R1052 VCC.n507 VCC.n42 10.6151
R1053 VCC.n510 VCC.n509 10.6151
R1054 VCC.n510 VCC.n501 10.6151
R1055 VCC.n516 VCC.n501 10.6151
R1056 VCC.n517 VCC.n516 10.6151
R1057 VCC.n518 VCC.n517 10.6151
R1058 VCC.n518 VCC.n499 10.6151
R1059 VCC.n524 VCC.n499 10.6151
R1060 VCC.n525 VCC.n524 10.6151
R1061 VCC.n526 VCC.n525 10.6151
R1062 VCC.n526 VCC.n497 10.6151
R1063 VCC.n532 VCC.n497 10.6151
R1064 VCC.n533 VCC.n532 10.6151
R1065 VCC.n534 VCC.n533 10.6151
R1066 VCC.n534 VCC.n495 10.6151
R1067 VCC.n540 VCC.n495 10.6151
R1068 VCC.n543 VCC.n542 10.6151
R1069 VCC.n543 VCC.n491 10.6151
R1070 VCC.n549 VCC.n491 10.6151
R1071 VCC.n550 VCC.n549 10.6151
R1072 VCC.n551 VCC.n550 10.6151
R1073 VCC.n551 VCC.n489 10.6151
R1074 VCC.n557 VCC.n489 10.6151
R1075 VCC.n558 VCC.n557 10.6151
R1076 VCC.n559 VCC.n558 10.6151
R1077 VCC.n559 VCC.n487 10.6151
R1078 VCC.n565 VCC.n487 10.6151
R1079 VCC.n566 VCC.n565 10.6151
R1080 VCC.n218 VCC.n194 10.6151
R1081 VCC.n221 VCC.n220 10.6151
R1082 VCC.n221 VCC.n212 10.6151
R1083 VCC.n227 VCC.n212 10.6151
R1084 VCC.n228 VCC.n227 10.6151
R1085 VCC.n229 VCC.n228 10.6151
R1086 VCC.n229 VCC.n210 10.6151
R1087 VCC.n235 VCC.n210 10.6151
R1088 VCC.n236 VCC.n235 10.6151
R1089 VCC.n237 VCC.n236 10.6151
R1090 VCC.n237 VCC.n208 10.6151
R1091 VCC.n243 VCC.n208 10.6151
R1092 VCC.n244 VCC.n243 10.6151
R1093 VCC.n245 VCC.n244 10.6151
R1094 VCC.n245 VCC.n206 10.6151
R1095 VCC.n251 VCC.n206 10.6151
R1096 VCC.n254 VCC.n253 10.6151
R1097 VCC.n254 VCC.n202 10.6151
R1098 VCC.n260 VCC.n202 10.6151
R1099 VCC.n261 VCC.n260 10.6151
R1100 VCC.n262 VCC.n261 10.6151
R1101 VCC.n262 VCC.n200 10.6151
R1102 VCC.n268 VCC.n200 10.6151
R1103 VCC.n269 VCC.n268 10.6151
R1104 VCC.n270 VCC.n269 10.6151
R1105 VCC.n270 VCC.n198 10.6151
R1106 VCC.n276 VCC.n198 10.6151
R1107 VCC.n277 VCC.n276 10.6151
R1108 VCC.n508 VCC.n507 10.3029
R1109 VCC.n219 VCC.n218 10.3029
R1110 VCC.n619 VCC.n0 9.3005
R1111 VCC.n618 VCC.n617 9.3005
R1112 VCC.n616 VCC.n6 9.3005
R1113 VCC.n615 VCC.n614 9.3005
R1114 VCC.n613 VCC.n7 9.3005
R1115 VCC.n612 VCC.n611 9.3005
R1116 VCC.n610 VCC.n11 9.3005
R1117 VCC.n609 VCC.n608 9.3005
R1118 VCC.n607 VCC.n12 9.3005
R1119 VCC.n606 VCC.n605 9.3005
R1120 VCC.n604 VCC.n16 9.3005
R1121 VCC.n603 VCC.n602 9.3005
R1122 VCC.n601 VCC.n17 9.3005
R1123 VCC.n600 VCC.n599 9.3005
R1124 VCC.n598 VCC.n21 9.3005
R1125 VCC.n597 VCC.n596 9.3005
R1126 VCC.n595 VCC.n22 9.3005
R1127 VCC.n594 VCC.n593 9.3005
R1128 VCC.n592 VCC.n26 9.3005
R1129 VCC.n591 VCC.n590 9.3005
R1130 VCC.n589 VCC.n27 9.3005
R1131 VCC.n588 VCC.n587 9.3005
R1132 VCC.n586 VCC.n31 9.3005
R1133 VCC.n585 VCC.n584 9.3005
R1134 VCC.n583 VCC.n32 9.3005
R1135 VCC.n582 VCC.n581 9.3005
R1136 VCC.n580 VCC.n36 9.3005
R1137 VCC.n579 VCC.n578 9.3005
R1138 VCC.n577 VCC.n37 9.3005
R1139 VCC.n576 VCC.n575 9.3005
R1140 VCC.n574 VCC.n41 9.3005
R1141 VCC.n573 VCC.n572 9.3005
R1142 VCC.n189 VCC.n188 9.3005
R1143 VCC.n292 VCC.n291 9.3005
R1144 VCC.n293 VCC.n187 9.3005
R1145 VCC.n295 VCC.n294 9.3005
R1146 VCC.n177 VCC.n176 9.3005
R1147 VCC.n308 VCC.n307 9.3005
R1148 VCC.n309 VCC.n175 9.3005
R1149 VCC.n311 VCC.n310 9.3005
R1150 VCC.n165 VCC.n164 9.3005
R1151 VCC.n324 VCC.n323 9.3005
R1152 VCC.n325 VCC.n163 9.3005
R1153 VCC.n327 VCC.n326 9.3005
R1154 VCC.n152 VCC.n151 9.3005
R1155 VCC.n340 VCC.n339 9.3005
R1156 VCC.n341 VCC.n150 9.3005
R1157 VCC.n343 VCC.n342 9.3005
R1158 VCC.n141 VCC.n140 9.3005
R1159 VCC.n356 VCC.n355 9.3005
R1160 VCC.n357 VCC.n139 9.3005
R1161 VCC.n359 VCC.n358 9.3005
R1162 VCC.n128 VCC.n127 9.3005
R1163 VCC.n372 VCC.n371 9.3005
R1164 VCC.n373 VCC.n126 9.3005
R1165 VCC.n375 VCC.n374 9.3005
R1166 VCC.n117 VCC.n116 9.3005
R1167 VCC.n388 VCC.n387 9.3005
R1168 VCC.n389 VCC.n115 9.3005
R1169 VCC.n391 VCC.n390 9.3005
R1170 VCC.n104 VCC.n103 9.3005
R1171 VCC.n404 VCC.n403 9.3005
R1172 VCC.n405 VCC.n102 9.3005
R1173 VCC.n407 VCC.n406 9.3005
R1174 VCC.n98 VCC.n97 9.3005
R1175 VCC.n413 VCC.n412 9.3005
R1176 VCC.n414 VCC.n96 9.3005
R1177 VCC.n416 VCC.n415 9.3005
R1178 VCC.n91 VCC.n90 9.3005
R1179 VCC.n423 VCC.n422 9.3005
R1180 VCC.n424 VCC.n89 9.3005
R1181 VCC.n426 VCC.n425 9.3005
R1182 VCC.n84 VCC.n83 9.3005
R1183 VCC.n433 VCC.n432 9.3005
R1184 VCC.n434 VCC.n82 9.3005
R1185 VCC.n436 VCC.n435 9.3005
R1186 VCC.n77 VCC.n76 9.3005
R1187 VCC.n443 VCC.n442 9.3005
R1188 VCC.n444 VCC.n75 9.3005
R1189 VCC.n446 VCC.n445 9.3005
R1190 VCC.n70 VCC.n69 9.3005
R1191 VCC.n453 VCC.n452 9.3005
R1192 VCC.n454 VCC.n68 9.3005
R1193 VCC.n456 VCC.n455 9.3005
R1194 VCC.n63 VCC.n62 9.3005
R1195 VCC.n463 VCC.n462 9.3005
R1196 VCC.n464 VCC.n61 9.3005
R1197 VCC.n466 VCC.n465 9.3005
R1198 VCC.n56 VCC.n55 9.3005
R1199 VCC.n475 VCC.n474 9.3005
R1200 VCC.n476 VCC.n54 9.3005
R1201 VCC.n478 VCC.n477 9.3005
R1202 VCC.n51 VCC.n50 9.3005
R1203 VCC.n485 VCC.n484 9.3005
R1204 VCC.n486 VCC.n49 9.3005
R1205 VCC.n568 VCC.n567 9.3005
R1206 VCC.n279 VCC.n278 9.3005
R1207 VCC.n284 VCC.n283 9.3005
R1208 VCC.n285 VCC.n193 9.3005
R1209 VCC.n287 VCC.n286 9.3005
R1210 VCC.n183 VCC.n182 9.3005
R1211 VCC.n300 VCC.n299 9.3005
R1212 VCC.n301 VCC.n181 9.3005
R1213 VCC.n303 VCC.n302 9.3005
R1214 VCC.n171 VCC.n170 9.3005
R1215 VCC.n316 VCC.n315 9.3005
R1216 VCC.n317 VCC.n169 9.3005
R1217 VCC.n319 VCC.n318 9.3005
R1218 VCC.n159 VCC.n158 9.3005
R1219 VCC.n332 VCC.n331 9.3005
R1220 VCC.n333 VCC.n157 9.3005
R1221 VCC.n335 VCC.n334 9.3005
R1222 VCC.n147 VCC.n146 9.3005
R1223 VCC.n348 VCC.n347 9.3005
R1224 VCC.n349 VCC.n145 9.3005
R1225 VCC.n351 VCC.n350 9.3005
R1226 VCC.n135 VCC.n134 9.3005
R1227 VCC.n364 VCC.n363 9.3005
R1228 VCC.n365 VCC.n133 9.3005
R1229 VCC.n367 VCC.n366 9.3005
R1230 VCC.n123 VCC.n122 9.3005
R1231 VCC.n380 VCC.n379 9.3005
R1232 VCC.n381 VCC.n121 9.3005
R1233 VCC.n383 VCC.n382 9.3005
R1234 VCC.n111 VCC.n110 9.3005
R1235 VCC.n396 VCC.n395 9.3005
R1236 VCC.n397 VCC.n109 9.3005
R1237 VCC.n399 VCC.n398 9.3005
R1238 VCC.n2 VCC.n1 9.3005
R1239 VCC.n621 VCC.n620 9.3005
R1240 VCC.n542 VCC.n541 5.93221
R1241 VCC.n253 VCC.n252 5.93221
R1242 VCC.n541 VCC.n540 4.68343
R1243 VCC.n252 VCC.n251 4.68343
R1244 VCC.n155 VCC.t15 3.05516
R1245 VCC.n449 VCC.t18 3.05516
R1246 VCC.n509 VCC.n508 0.312695
R1247 VCC.n220 VCC.n219 0.312695
R1248 VCC.n617 VCC.n0 0.152939
R1249 VCC.n617 VCC.n616 0.152939
R1250 VCC.n616 VCC.n615 0.152939
R1251 VCC.n615 VCC.n7 0.152939
R1252 VCC.n611 VCC.n7 0.152939
R1253 VCC.n611 VCC.n610 0.152939
R1254 VCC.n610 VCC.n609 0.152939
R1255 VCC.n609 VCC.n12 0.152939
R1256 VCC.n605 VCC.n12 0.152939
R1257 VCC.n605 VCC.n604 0.152939
R1258 VCC.n604 VCC.n603 0.152939
R1259 VCC.n603 VCC.n17 0.152939
R1260 VCC.n599 VCC.n17 0.152939
R1261 VCC.n599 VCC.n598 0.152939
R1262 VCC.n598 VCC.n597 0.152939
R1263 VCC.n597 VCC.n22 0.152939
R1264 VCC.n593 VCC.n22 0.152939
R1265 VCC.n593 VCC.n592 0.152939
R1266 VCC.n592 VCC.n591 0.152939
R1267 VCC.n591 VCC.n27 0.152939
R1268 VCC.n587 VCC.n27 0.152939
R1269 VCC.n587 VCC.n586 0.152939
R1270 VCC.n586 VCC.n585 0.152939
R1271 VCC.n585 VCC.n32 0.152939
R1272 VCC.n581 VCC.n32 0.152939
R1273 VCC.n581 VCC.n580 0.152939
R1274 VCC.n580 VCC.n579 0.152939
R1275 VCC.n579 VCC.n37 0.152939
R1276 VCC.n575 VCC.n37 0.152939
R1277 VCC.n575 VCC.n574 0.152939
R1278 VCC.n574 VCC.n573 0.152939
R1279 VCC.n278 VCC.n188 0.152939
R1280 VCC.n292 VCC.n188 0.152939
R1281 VCC.n293 VCC.n292 0.152939
R1282 VCC.n294 VCC.n293 0.152939
R1283 VCC.n294 VCC.n176 0.152939
R1284 VCC.n308 VCC.n176 0.152939
R1285 VCC.n309 VCC.n308 0.152939
R1286 VCC.n310 VCC.n309 0.152939
R1287 VCC.n310 VCC.n164 0.152939
R1288 VCC.n324 VCC.n164 0.152939
R1289 VCC.n325 VCC.n324 0.152939
R1290 VCC.n326 VCC.n325 0.152939
R1291 VCC.n326 VCC.n151 0.152939
R1292 VCC.n340 VCC.n151 0.152939
R1293 VCC.n341 VCC.n340 0.152939
R1294 VCC.n342 VCC.n341 0.152939
R1295 VCC.n342 VCC.n140 0.152939
R1296 VCC.n356 VCC.n140 0.152939
R1297 VCC.n357 VCC.n356 0.152939
R1298 VCC.n358 VCC.n357 0.152939
R1299 VCC.n358 VCC.n127 0.152939
R1300 VCC.n372 VCC.n127 0.152939
R1301 VCC.n373 VCC.n372 0.152939
R1302 VCC.n374 VCC.n373 0.152939
R1303 VCC.n374 VCC.n116 0.152939
R1304 VCC.n388 VCC.n116 0.152939
R1305 VCC.n389 VCC.n388 0.152939
R1306 VCC.n390 VCC.n389 0.152939
R1307 VCC.n390 VCC.n103 0.152939
R1308 VCC.n404 VCC.n103 0.152939
R1309 VCC.n405 VCC.n404 0.152939
R1310 VCC.n406 VCC.n405 0.152939
R1311 VCC.n406 VCC.n97 0.152939
R1312 VCC.n413 VCC.n97 0.152939
R1313 VCC.n414 VCC.n413 0.152939
R1314 VCC.n415 VCC.n414 0.152939
R1315 VCC.n415 VCC.n90 0.152939
R1316 VCC.n423 VCC.n90 0.152939
R1317 VCC.n424 VCC.n423 0.152939
R1318 VCC.n425 VCC.n424 0.152939
R1319 VCC.n425 VCC.n83 0.152939
R1320 VCC.n433 VCC.n83 0.152939
R1321 VCC.n434 VCC.n433 0.152939
R1322 VCC.n435 VCC.n434 0.152939
R1323 VCC.n435 VCC.n76 0.152939
R1324 VCC.n443 VCC.n76 0.152939
R1325 VCC.n444 VCC.n443 0.152939
R1326 VCC.n445 VCC.n444 0.152939
R1327 VCC.n445 VCC.n69 0.152939
R1328 VCC.n453 VCC.n69 0.152939
R1329 VCC.n454 VCC.n453 0.152939
R1330 VCC.n455 VCC.n454 0.152939
R1331 VCC.n455 VCC.n62 0.152939
R1332 VCC.n463 VCC.n62 0.152939
R1333 VCC.n464 VCC.n463 0.152939
R1334 VCC.n465 VCC.n464 0.152939
R1335 VCC.n465 VCC.n55 0.152939
R1336 VCC.n475 VCC.n55 0.152939
R1337 VCC.n476 VCC.n475 0.152939
R1338 VCC.n477 VCC.n476 0.152939
R1339 VCC.n477 VCC.n50 0.152939
R1340 VCC.n485 VCC.n50 0.152939
R1341 VCC.n486 VCC.n485 0.152939
R1342 VCC.n567 VCC.n486 0.152939
R1343 VCC.n285 VCC.n284 0.152939
R1344 VCC.n286 VCC.n285 0.152939
R1345 VCC.n286 VCC.n182 0.152939
R1346 VCC.n300 VCC.n182 0.152939
R1347 VCC.n301 VCC.n300 0.152939
R1348 VCC.n302 VCC.n301 0.152939
R1349 VCC.n302 VCC.n170 0.152939
R1350 VCC.n316 VCC.n170 0.152939
R1351 VCC.n317 VCC.n316 0.152939
R1352 VCC.n318 VCC.n317 0.152939
R1353 VCC.n318 VCC.n158 0.152939
R1354 VCC.n332 VCC.n158 0.152939
R1355 VCC.n333 VCC.n332 0.152939
R1356 VCC.n334 VCC.n333 0.152939
R1357 VCC.n334 VCC.n146 0.152939
R1358 VCC.n348 VCC.n146 0.152939
R1359 VCC.n349 VCC.n348 0.152939
R1360 VCC.n350 VCC.n349 0.152939
R1361 VCC.n350 VCC.n134 0.152939
R1362 VCC.n364 VCC.n134 0.152939
R1363 VCC.n365 VCC.n364 0.152939
R1364 VCC.n366 VCC.n365 0.152939
R1365 VCC.n366 VCC.n122 0.152939
R1366 VCC.n380 VCC.n122 0.152939
R1367 VCC.n381 VCC.n380 0.152939
R1368 VCC.n382 VCC.n381 0.152939
R1369 VCC.n382 VCC.n110 0.152939
R1370 VCC.n396 VCC.n110 0.152939
R1371 VCC.n397 VCC.n396 0.152939
R1372 VCC.n398 VCC.n397 0.152939
R1373 VCC.n398 VCC.n1 0.152939
R1374 VCC.n621 VCC.n1 0.13922
R1375 VCC VCC.n0 0.0767195
R1376 VCC VCC.n621 0.063
R1377 VSS.n97 VSS.n96 585
R1378 VSS.n96 VSS.n94 585
R1379 VSS.n387 VSS.n386 585
R1380 VSS.n388 VSS.n387 585
R1381 VSS.n88 VSS.n87 585
R1382 VSS.n95 VSS.n88 585
R1383 VSS.n398 VSS.n397 585
R1384 VSS.n397 VSS.n396 585
R1385 VSS.n85 VSS.n84 585
R1386 VSS.n84 VSS.n83 585
R1387 VSS.n403 VSS.n402 585
R1388 VSS.n404 VSS.n403 585
R1389 VSS.n76 VSS.n75 585
R1390 VSS.n77 VSS.n76 585
R1391 VSS.n415 VSS.n414 585
R1392 VSS.n414 VSS.n413 585
R1393 VSS.n73 VSS.n72 585
R1394 VSS.n412 VSS.n72 585
R1395 VSS.n420 VSS.n419 585
R1396 VSS.n421 VSS.n420 585
R1397 VSS.n65 VSS.n64 585
R1398 VSS.n66 VSS.n65 585
R1399 VSS.n432 VSS.n431 585
R1400 VSS.n431 VSS.n430 585
R1401 VSS.n62 VSS.n61 585
R1402 VSS.n429 VSS.n61 585
R1403 VSS.n437 VSS.n436 585
R1404 VSS.n438 VSS.n437 585
R1405 VSS.n54 VSS.n53 585
R1406 VSS.n55 VSS.n54 585
R1407 VSS.n450 VSS.n449 585
R1408 VSS.n449 VSS.n448 585
R1409 VSS.n51 VSS.n50 585
R1410 VSS.n447 VSS.n50 585
R1411 VSS.n455 VSS.n454 585
R1412 VSS.n456 VSS.n455 585
R1413 VSS.n49 VSS.n48 585
R1414 VSS.n457 VSS.n49 585
R1415 VSS.n462 VSS.n461 585
R1416 VSS.n461 VSS.n460 585
R1417 VSS.n46 VSS.n45 585
R1418 VSS.n459 VSS.n45 585
R1419 VSS.n467 VSS.n466 585
R1420 VSS.n468 VSS.n467 585
R1421 VSS.n44 VSS.n43 585
R1422 VSS.n469 VSS.n44 585
R1423 VSS.n474 VSS.n473 585
R1424 VSS.n473 VSS.n472 585
R1425 VSS.n41 VSS.n40 585
R1426 VSS.n471 VSS.n40 585
R1427 VSS.n479 VSS.n478 585
R1428 VSS.n480 VSS.n479 585
R1429 VSS.n39 VSS.n38 585
R1430 VSS.n481 VSS.n39 585
R1431 VSS.n484 VSS.n483 585
R1432 VSS.n483 VSS.n482 585
R1433 VSS.n36 VSS.n35 585
R1434 VSS.n35 VSS.n34 585
R1435 VSS.n489 VSS.n488 585
R1436 VSS.n490 VSS.n489 585
R1437 VSS.n32 VSS.n31 585
R1438 VSS.n491 VSS.n32 585
R1439 VSS.n494 VSS.n493 585
R1440 VSS.n493 VSS.n492 585
R1441 VSS.n29 VSS.n27 585
R1442 VSS.n27 VSS.n25 585
R1443 VSS.n782 VSS.n781 585
R1444 VSS.n783 VSS.n782 585
R1445 VSS.n785 VSS.n784 585
R1446 VSS.n784 VSS.n783 585
R1447 VSS.n23 VSS.n21 585
R1448 VSS.n25 VSS.n23 585
R1449 VSS.n789 VSS.n20 585
R1450 VSS.n492 VSS.n20 585
R1451 VSS.n790 VSS.n19 585
R1452 VSS.n491 VSS.n19 585
R1453 VSS.n791 VSS.n18 585
R1454 VSS.n490 VSS.n18 585
R1455 VSS.n33 VSS.n16 585
R1456 VSS.n34 VSS.n33 585
R1457 VSS.n795 VSS.n15 585
R1458 VSS.n482 VSS.n15 585
R1459 VSS.n796 VSS.n14 585
R1460 VSS.n481 VSS.n14 585
R1461 VSS.n797 VSS.n13 585
R1462 VSS.n480 VSS.n13 585
R1463 VSS.n470 VSS.n11 585
R1464 VSS.n471 VSS.n470 585
R1465 VSS.n801 VSS.n10 585
R1466 VSS.n472 VSS.n10 585
R1467 VSS.n802 VSS.n9 585
R1468 VSS.n469 VSS.n9 585
R1469 VSS.n803 VSS.n8 585
R1470 VSS.n468 VSS.n8 585
R1471 VSS.n458 VSS.n6 585
R1472 VSS.n459 VSS.n458 585
R1473 VSS.n807 VSS.n5 585
R1474 VSS.n460 VSS.n5 585
R1475 VSS.n808 VSS.n4 585
R1476 VSS.n457 VSS.n4 585
R1477 VSS.n809 VSS.n3 585
R1478 VSS.n456 VSS.n3 585
R1479 VSS.n446 VSS.n2 585
R1480 VSS.n447 VSS.n446 585
R1481 VSS.n445 VSS.n444 585
R1482 VSS.n448 VSS.n445 585
R1483 VSS.n57 VSS.n56 585
R1484 VSS.n56 VSS.n55 585
R1485 VSS.n440 VSS.n439 585
R1486 VSS.n439 VSS.n438 585
R1487 VSS.n60 VSS.n59 585
R1488 VSS.n429 VSS.n60 585
R1489 VSS.n428 VSS.n427 585
R1490 VSS.n430 VSS.n428 585
R1491 VSS.n68 VSS.n67 585
R1492 VSS.n67 VSS.n66 585
R1493 VSS.n423 VSS.n422 585
R1494 VSS.n422 VSS.n421 585
R1495 VSS.n71 VSS.n70 585
R1496 VSS.n412 VSS.n71 585
R1497 VSS.n411 VSS.n410 585
R1498 VSS.n413 VSS.n411 585
R1499 VSS.n79 VSS.n78 585
R1500 VSS.n78 VSS.n77 585
R1501 VSS.n406 VSS.n405 585
R1502 VSS.n405 VSS.n404 585
R1503 VSS.n82 VSS.n81 585
R1504 VSS.n83 VSS.n82 585
R1505 VSS.n395 VSS.n394 585
R1506 VSS.n396 VSS.n395 585
R1507 VSS.n90 VSS.n89 585
R1508 VSS.n95 VSS.n89 585
R1509 VSS.n390 VSS.n389 585
R1510 VSS.n389 VSS.n388 585
R1511 VSS.n93 VSS.n92 585
R1512 VSS.n94 VSS.n93 585
R1513 VSS.n24 VSS.n22 585
R1514 VSS.n586 VSS.n583 585
R1515 VSS.n588 VSS.n587 585
R1516 VSS.n590 VSS.n580 585
R1517 VSS.n592 VSS.n591 585
R1518 VSS.n594 VSS.n578 585
R1519 VSS.n596 VSS.n595 585
R1520 VSS.n597 VSS.n577 585
R1521 VSS.n599 VSS.n598 585
R1522 VSS.n601 VSS.n575 585
R1523 VSS.n603 VSS.n602 585
R1524 VSS.n604 VSS.n574 585
R1525 VSS.n606 VSS.n605 585
R1526 VSS.n608 VSS.n572 585
R1527 VSS.n610 VSS.n609 585
R1528 VSS.n611 VSS.n571 585
R1529 VSS.n613 VSS.n612 585
R1530 VSS.n615 VSS.n569 585
R1531 VSS.n617 VSS.n616 585
R1532 VSS.n618 VSS.n568 585
R1533 VSS.n620 VSS.n619 585
R1534 VSS.n622 VSS.n566 585
R1535 VSS.n624 VSS.n623 585
R1536 VSS.n625 VSS.n565 585
R1537 VSS.n627 VSS.n626 585
R1538 VSS.n629 VSS.n563 585
R1539 VSS.n631 VSS.n630 585
R1540 VSS.n632 VSS.n562 585
R1541 VSS.n634 VSS.n633 585
R1542 VSS.n636 VSS.n560 585
R1543 VSS.n638 VSS.n637 585
R1544 VSS.n639 VSS.n559 585
R1545 VSS.n641 VSS.n640 585
R1546 VSS.n643 VSS.n557 585
R1547 VSS.n645 VSS.n644 585
R1548 VSS.n646 VSS.n556 585
R1549 VSS.n648 VSS.n647 585
R1550 VSS.n650 VSS.n554 585
R1551 VSS.n652 VSS.n651 585
R1552 VSS.n653 VSS.n553 585
R1553 VSS.n655 VSS.n654 585
R1554 VSS.n657 VSS.n551 585
R1555 VSS.n659 VSS.n658 585
R1556 VSS.n660 VSS.n550 585
R1557 VSS.n662 VSS.n661 585
R1558 VSS.n664 VSS.n548 585
R1559 VSS.n666 VSS.n665 585
R1560 VSS.n667 VSS.n547 585
R1561 VSS.n669 VSS.n668 585
R1562 VSS.n671 VSS.n545 585
R1563 VSS.n673 VSS.n672 585
R1564 VSS.n674 VSS.n544 585
R1565 VSS.n676 VSS.n675 585
R1566 VSS.n678 VSS.n542 585
R1567 VSS.n680 VSS.n679 585
R1568 VSS.n681 VSS.n541 585
R1569 VSS.n683 VSS.n682 585
R1570 VSS.n685 VSS.n540 585
R1571 VSS.n687 VSS.n686 585
R1572 VSS.n688 VSS.n535 585
R1573 VSS.n690 VSS.n689 585
R1574 VSS.n692 VSS.n533 585
R1575 VSS.n694 VSS.n693 585
R1576 VSS.n695 VSS.n532 585
R1577 VSS.n697 VSS.n696 585
R1578 VSS.n699 VSS.n530 585
R1579 VSS.n701 VSS.n700 585
R1580 VSS.n702 VSS.n529 585
R1581 VSS.n704 VSS.n703 585
R1582 VSS.n706 VSS.n527 585
R1583 VSS.n708 VSS.n707 585
R1584 VSS.n709 VSS.n526 585
R1585 VSS.n711 VSS.n710 585
R1586 VSS.n713 VSS.n524 585
R1587 VSS.n715 VSS.n714 585
R1588 VSS.n716 VSS.n523 585
R1589 VSS.n718 VSS.n717 585
R1590 VSS.n720 VSS.n521 585
R1591 VSS.n722 VSS.n721 585
R1592 VSS.n723 VSS.n520 585
R1593 VSS.n725 VSS.n724 585
R1594 VSS.n727 VSS.n518 585
R1595 VSS.n729 VSS.n728 585
R1596 VSS.n730 VSS.n517 585
R1597 VSS.n732 VSS.n731 585
R1598 VSS.n734 VSS.n515 585
R1599 VSS.n736 VSS.n735 585
R1600 VSS.n737 VSS.n514 585
R1601 VSS.n739 VSS.n738 585
R1602 VSS.n741 VSS.n512 585
R1603 VSS.n743 VSS.n742 585
R1604 VSS.n744 VSS.n511 585
R1605 VSS.n746 VSS.n745 585
R1606 VSS.n748 VSS.n509 585
R1607 VSS.n750 VSS.n749 585
R1608 VSS.n751 VSS.n508 585
R1609 VSS.n753 VSS.n752 585
R1610 VSS.n755 VSS.n506 585
R1611 VSS.n757 VSS.n756 585
R1612 VSS.n758 VSS.n505 585
R1613 VSS.n760 VSS.n759 585
R1614 VSS.n762 VSS.n503 585
R1615 VSS.n764 VSS.n763 585
R1616 VSS.n765 VSS.n502 585
R1617 VSS.n767 VSS.n766 585
R1618 VSS.n769 VSS.n500 585
R1619 VSS.n771 VSS.n770 585
R1620 VSS.n772 VSS.n499 585
R1621 VSS.n774 VSS.n773 585
R1622 VSS.n776 VSS.n497 585
R1623 VSS.n778 VSS.n777 585
R1624 VSS.n779 VSS.n28 585
R1625 VSS.n383 VSS.n382 585
R1626 VSS.n99 VSS.n98 585
R1627 VSS.n379 VSS.n378 585
R1628 VSS.n380 VSS.n379 585
R1629 VSS.n377 VSS.n155 585
R1630 VSS.n376 VSS.n375 585
R1631 VSS.n374 VSS.n373 585
R1632 VSS.n372 VSS.n371 585
R1633 VSS.n370 VSS.n369 585
R1634 VSS.n368 VSS.n367 585
R1635 VSS.n366 VSS.n365 585
R1636 VSS.n364 VSS.n363 585
R1637 VSS.n362 VSS.n361 585
R1638 VSS.n360 VSS.n359 585
R1639 VSS.n358 VSS.n357 585
R1640 VSS.n356 VSS.n355 585
R1641 VSS.n354 VSS.n353 585
R1642 VSS.n352 VSS.n351 585
R1643 VSS.n350 VSS.n349 585
R1644 VSS.n348 VSS.n347 585
R1645 VSS.n346 VSS.n345 585
R1646 VSS.n344 VSS.n343 585
R1647 VSS.n342 VSS.n341 585
R1648 VSS.n340 VSS.n339 585
R1649 VSS.n338 VSS.n337 585
R1650 VSS.n336 VSS.n335 585
R1651 VSS.n334 VSS.n333 585
R1652 VSS.n332 VSS.n331 585
R1653 VSS.n330 VSS.n329 585
R1654 VSS.n328 VSS.n327 585
R1655 VSS.n326 VSS.n325 585
R1656 VSS.n324 VSS.n323 585
R1657 VSS.n322 VSS.n321 585
R1658 VSS.n320 VSS.n319 585
R1659 VSS.n318 VSS.n317 585
R1660 VSS.n316 VSS.n315 585
R1661 VSS.n314 VSS.n313 585
R1662 VSS.n312 VSS.n311 585
R1663 VSS.n310 VSS.n309 585
R1664 VSS.n308 VSS.n307 585
R1665 VSS.n306 VSS.n305 585
R1666 VSS.n304 VSS.n303 585
R1667 VSS.n302 VSS.n301 585
R1668 VSS.n300 VSS.n299 585
R1669 VSS.n298 VSS.n297 585
R1670 VSS.n296 VSS.n295 585
R1671 VSS.n294 VSS.n293 585
R1672 VSS.n292 VSS.n291 585
R1673 VSS.n290 VSS.n289 585
R1674 VSS.n288 VSS.n287 585
R1675 VSS.n286 VSS.n285 585
R1676 VSS.n284 VSS.n283 585
R1677 VSS.n282 VSS.n281 585
R1678 VSS.n280 VSS.n279 585
R1679 VSS.n278 VSS.n277 585
R1680 VSS.n275 VSS.n274 585
R1681 VSS.n273 VSS.n272 585
R1682 VSS.n271 VSS.n270 585
R1683 VSS.n269 VSS.n268 585
R1684 VSS.n267 VSS.n266 585
R1685 VSS.n265 VSS.n264 585
R1686 VSS.n263 VSS.n262 585
R1687 VSS.n261 VSS.n260 585
R1688 VSS.n259 VSS.n258 585
R1689 VSS.n257 VSS.n256 585
R1690 VSS.n255 VSS.n254 585
R1691 VSS.n253 VSS.n252 585
R1692 VSS.n251 VSS.n250 585
R1693 VSS.n249 VSS.n248 585
R1694 VSS.n247 VSS.n246 585
R1695 VSS.n245 VSS.n244 585
R1696 VSS.n243 VSS.n242 585
R1697 VSS.n241 VSS.n240 585
R1698 VSS.n239 VSS.n238 585
R1699 VSS.n237 VSS.n236 585
R1700 VSS.n235 VSS.n234 585
R1701 VSS.n233 VSS.n232 585
R1702 VSS.n231 VSS.n230 585
R1703 VSS.n229 VSS.n228 585
R1704 VSS.n227 VSS.n226 585
R1705 VSS.n225 VSS.n224 585
R1706 VSS.n223 VSS.n222 585
R1707 VSS.n221 VSS.n220 585
R1708 VSS.n219 VSS.n218 585
R1709 VSS.n217 VSS.n216 585
R1710 VSS.n215 VSS.n214 585
R1711 VSS.n213 VSS.n212 585
R1712 VSS.n211 VSS.n210 585
R1713 VSS.n209 VSS.n208 585
R1714 VSS.n207 VSS.n206 585
R1715 VSS.n205 VSS.n204 585
R1716 VSS.n203 VSS.n202 585
R1717 VSS.n201 VSS.n200 585
R1718 VSS.n199 VSS.n198 585
R1719 VSS.n197 VSS.n196 585
R1720 VSS.n195 VSS.n194 585
R1721 VSS.n193 VSS.n192 585
R1722 VSS.n191 VSS.n190 585
R1723 VSS.n189 VSS.n188 585
R1724 VSS.n187 VSS.n186 585
R1725 VSS.n185 VSS.n184 585
R1726 VSS.n183 VSS.n182 585
R1727 VSS.n181 VSS.n180 585
R1728 VSS.n179 VSS.n178 585
R1729 VSS.n177 VSS.n176 585
R1730 VSS.n175 VSS.n174 585
R1731 VSS.n173 VSS.n172 585
R1732 VSS.n171 VSS.n170 585
R1733 VSS.n169 VSS.n168 585
R1734 VSS.n167 VSS.n166 585
R1735 VSS.n165 VSS.n164 585
R1736 VSS.n163 VSS.n162 585
R1737 VSS.n161 VSS.n154 585
R1738 VSS.n380 VSS.n154 585
R1739 VSS.n382 VSS.n96 545.355
R1740 VSS.n154 VSS.n93 545.355
R1741 VSS.n782 VSS.n28 545.355
R1742 VSS.n784 VSS.n24 545.355
R1743 VSS.n536 VSS.t16 451.034
R1744 VSS.n581 VSS.t12 451.034
R1745 VSS.n158 VSS.t9 451.034
R1746 VSS.n156 VSS.t5 451.034
R1747 VSS.n585 VSS.n26 256.663
R1748 VSS.n584 VSS.n26 256.663
R1749 VSS.n593 VSS.n26 256.663
R1750 VSS.n579 VSS.n26 256.663
R1751 VSS.n600 VSS.n26 256.663
R1752 VSS.n576 VSS.n26 256.663
R1753 VSS.n607 VSS.n26 256.663
R1754 VSS.n573 VSS.n26 256.663
R1755 VSS.n614 VSS.n26 256.663
R1756 VSS.n570 VSS.n26 256.663
R1757 VSS.n621 VSS.n26 256.663
R1758 VSS.n567 VSS.n26 256.663
R1759 VSS.n628 VSS.n26 256.663
R1760 VSS.n564 VSS.n26 256.663
R1761 VSS.n635 VSS.n26 256.663
R1762 VSS.n561 VSS.n26 256.663
R1763 VSS.n642 VSS.n26 256.663
R1764 VSS.n558 VSS.n26 256.663
R1765 VSS.n649 VSS.n26 256.663
R1766 VSS.n555 VSS.n26 256.663
R1767 VSS.n656 VSS.n26 256.663
R1768 VSS.n552 VSS.n26 256.663
R1769 VSS.n663 VSS.n26 256.663
R1770 VSS.n549 VSS.n26 256.663
R1771 VSS.n670 VSS.n26 256.663
R1772 VSS.n546 VSS.n26 256.663
R1773 VSS.n677 VSS.n26 256.663
R1774 VSS.n543 VSS.n26 256.663
R1775 VSS.n684 VSS.n26 256.663
R1776 VSS.n539 VSS.n26 256.663
R1777 VSS.n691 VSS.n26 256.663
R1778 VSS.n534 VSS.n26 256.663
R1779 VSS.n698 VSS.n26 256.663
R1780 VSS.n531 VSS.n26 256.663
R1781 VSS.n705 VSS.n26 256.663
R1782 VSS.n528 VSS.n26 256.663
R1783 VSS.n712 VSS.n26 256.663
R1784 VSS.n525 VSS.n26 256.663
R1785 VSS.n719 VSS.n26 256.663
R1786 VSS.n522 VSS.n26 256.663
R1787 VSS.n726 VSS.n26 256.663
R1788 VSS.n519 VSS.n26 256.663
R1789 VSS.n733 VSS.n26 256.663
R1790 VSS.n516 VSS.n26 256.663
R1791 VSS.n740 VSS.n26 256.663
R1792 VSS.n513 VSS.n26 256.663
R1793 VSS.n747 VSS.n26 256.663
R1794 VSS.n510 VSS.n26 256.663
R1795 VSS.n754 VSS.n26 256.663
R1796 VSS.n507 VSS.n26 256.663
R1797 VSS.n761 VSS.n26 256.663
R1798 VSS.n504 VSS.n26 256.663
R1799 VSS.n768 VSS.n26 256.663
R1800 VSS.n501 VSS.n26 256.663
R1801 VSS.n775 VSS.n26 256.663
R1802 VSS.n498 VSS.n26 256.663
R1803 VSS.n381 VSS.n380 256.663
R1804 VSS.n380 VSS.n100 256.663
R1805 VSS.n380 VSS.n101 256.663
R1806 VSS.n380 VSS.n102 256.663
R1807 VSS.n380 VSS.n103 256.663
R1808 VSS.n380 VSS.n104 256.663
R1809 VSS.n380 VSS.n105 256.663
R1810 VSS.n380 VSS.n106 256.663
R1811 VSS.n380 VSS.n107 256.663
R1812 VSS.n380 VSS.n108 256.663
R1813 VSS.n380 VSS.n109 256.663
R1814 VSS.n380 VSS.n110 256.663
R1815 VSS.n380 VSS.n111 256.663
R1816 VSS.n380 VSS.n112 256.663
R1817 VSS.n380 VSS.n113 256.663
R1818 VSS.n380 VSS.n114 256.663
R1819 VSS.n380 VSS.n115 256.663
R1820 VSS.n380 VSS.n116 256.663
R1821 VSS.n380 VSS.n117 256.663
R1822 VSS.n380 VSS.n118 256.663
R1823 VSS.n380 VSS.n119 256.663
R1824 VSS.n380 VSS.n120 256.663
R1825 VSS.n380 VSS.n121 256.663
R1826 VSS.n380 VSS.n122 256.663
R1827 VSS.n380 VSS.n123 256.663
R1828 VSS.n380 VSS.n124 256.663
R1829 VSS.n380 VSS.n125 256.663
R1830 VSS.n380 VSS.n126 256.663
R1831 VSS.n380 VSS.n127 256.663
R1832 VSS.n380 VSS.n128 256.663
R1833 VSS.n380 VSS.n129 256.663
R1834 VSS.n380 VSS.n130 256.663
R1835 VSS.n380 VSS.n131 256.663
R1836 VSS.n380 VSS.n132 256.663
R1837 VSS.n380 VSS.n133 256.663
R1838 VSS.n380 VSS.n134 256.663
R1839 VSS.n380 VSS.n135 256.663
R1840 VSS.n380 VSS.n136 256.663
R1841 VSS.n380 VSS.n137 256.663
R1842 VSS.n380 VSS.n138 256.663
R1843 VSS.n380 VSS.n139 256.663
R1844 VSS.n380 VSS.n140 256.663
R1845 VSS.n380 VSS.n141 256.663
R1846 VSS.n380 VSS.n142 256.663
R1847 VSS.n380 VSS.n143 256.663
R1848 VSS.n380 VSS.n144 256.663
R1849 VSS.n380 VSS.n145 256.663
R1850 VSS.n380 VSS.n146 256.663
R1851 VSS.n380 VSS.n147 256.663
R1852 VSS.n380 VSS.n148 256.663
R1853 VSS.n380 VSS.n149 256.663
R1854 VSS.n380 VSS.n150 256.663
R1855 VSS.n380 VSS.n151 256.663
R1856 VSS.n380 VSS.n152 256.663
R1857 VSS.n380 VSS.n153 256.663
R1858 VSS.n387 VSS.n96 240.244
R1859 VSS.n387 VSS.n88 240.244
R1860 VSS.n397 VSS.n88 240.244
R1861 VSS.n397 VSS.n84 240.244
R1862 VSS.n403 VSS.n84 240.244
R1863 VSS.n403 VSS.n76 240.244
R1864 VSS.n414 VSS.n76 240.244
R1865 VSS.n414 VSS.n72 240.244
R1866 VSS.n420 VSS.n72 240.244
R1867 VSS.n420 VSS.n65 240.244
R1868 VSS.n431 VSS.n65 240.244
R1869 VSS.n431 VSS.n61 240.244
R1870 VSS.n437 VSS.n61 240.244
R1871 VSS.n437 VSS.n54 240.244
R1872 VSS.n449 VSS.n54 240.244
R1873 VSS.n449 VSS.n50 240.244
R1874 VSS.n455 VSS.n50 240.244
R1875 VSS.n455 VSS.n49 240.244
R1876 VSS.n461 VSS.n49 240.244
R1877 VSS.n461 VSS.n45 240.244
R1878 VSS.n467 VSS.n45 240.244
R1879 VSS.n467 VSS.n44 240.244
R1880 VSS.n473 VSS.n44 240.244
R1881 VSS.n473 VSS.n40 240.244
R1882 VSS.n479 VSS.n40 240.244
R1883 VSS.n479 VSS.n39 240.244
R1884 VSS.n483 VSS.n39 240.244
R1885 VSS.n483 VSS.n35 240.244
R1886 VSS.n489 VSS.n35 240.244
R1887 VSS.n489 VSS.n32 240.244
R1888 VSS.n493 VSS.n32 240.244
R1889 VSS.n493 VSS.n27 240.244
R1890 VSS.n782 VSS.n27 240.244
R1891 VSS.n389 VSS.n93 240.244
R1892 VSS.n389 VSS.n89 240.244
R1893 VSS.n395 VSS.n89 240.244
R1894 VSS.n395 VSS.n82 240.244
R1895 VSS.n405 VSS.n82 240.244
R1896 VSS.n405 VSS.n78 240.244
R1897 VSS.n411 VSS.n78 240.244
R1898 VSS.n411 VSS.n71 240.244
R1899 VSS.n422 VSS.n71 240.244
R1900 VSS.n422 VSS.n67 240.244
R1901 VSS.n428 VSS.n67 240.244
R1902 VSS.n428 VSS.n60 240.244
R1903 VSS.n439 VSS.n60 240.244
R1904 VSS.n439 VSS.n56 240.244
R1905 VSS.n445 VSS.n56 240.244
R1906 VSS.n446 VSS.n445 240.244
R1907 VSS.n446 VSS.n3 240.244
R1908 VSS.n4 VSS.n3 240.244
R1909 VSS.n5 VSS.n4 240.244
R1910 VSS.n458 VSS.n5 240.244
R1911 VSS.n458 VSS.n8 240.244
R1912 VSS.n9 VSS.n8 240.244
R1913 VSS.n10 VSS.n9 240.244
R1914 VSS.n470 VSS.n10 240.244
R1915 VSS.n470 VSS.n13 240.244
R1916 VSS.n14 VSS.n13 240.244
R1917 VSS.n15 VSS.n14 240.244
R1918 VSS.n33 VSS.n15 240.244
R1919 VSS.n33 VSS.n18 240.244
R1920 VSS.n19 VSS.n18 240.244
R1921 VSS.n20 VSS.n19 240.244
R1922 VSS.n23 VSS.n20 240.244
R1923 VSS.n784 VSS.n23 240.244
R1924 VSS.n379 VSS.n99 163.367
R1925 VSS.n379 VSS.n155 163.367
R1926 VSS.n375 VSS.n374 163.367
R1927 VSS.n371 VSS.n370 163.367
R1928 VSS.n367 VSS.n366 163.367
R1929 VSS.n363 VSS.n362 163.367
R1930 VSS.n359 VSS.n358 163.367
R1931 VSS.n355 VSS.n354 163.367
R1932 VSS.n351 VSS.n350 163.367
R1933 VSS.n347 VSS.n346 163.367
R1934 VSS.n343 VSS.n342 163.367
R1935 VSS.n339 VSS.n338 163.367
R1936 VSS.n335 VSS.n334 163.367
R1937 VSS.n331 VSS.n330 163.367
R1938 VSS.n327 VSS.n326 163.367
R1939 VSS.n323 VSS.n322 163.367
R1940 VSS.n319 VSS.n318 163.367
R1941 VSS.n315 VSS.n314 163.367
R1942 VSS.n311 VSS.n310 163.367
R1943 VSS.n307 VSS.n306 163.367
R1944 VSS.n303 VSS.n302 163.367
R1945 VSS.n299 VSS.n298 163.367
R1946 VSS.n295 VSS.n294 163.367
R1947 VSS.n291 VSS.n290 163.367
R1948 VSS.n287 VSS.n286 163.367
R1949 VSS.n283 VSS.n282 163.367
R1950 VSS.n279 VSS.n278 163.367
R1951 VSS.n274 VSS.n273 163.367
R1952 VSS.n270 VSS.n269 163.367
R1953 VSS.n266 VSS.n265 163.367
R1954 VSS.n262 VSS.n261 163.367
R1955 VSS.n258 VSS.n257 163.367
R1956 VSS.n254 VSS.n253 163.367
R1957 VSS.n250 VSS.n249 163.367
R1958 VSS.n246 VSS.n245 163.367
R1959 VSS.n242 VSS.n241 163.367
R1960 VSS.n238 VSS.n237 163.367
R1961 VSS.n234 VSS.n233 163.367
R1962 VSS.n230 VSS.n229 163.367
R1963 VSS.n226 VSS.n225 163.367
R1964 VSS.n222 VSS.n221 163.367
R1965 VSS.n218 VSS.n217 163.367
R1966 VSS.n214 VSS.n213 163.367
R1967 VSS.n210 VSS.n209 163.367
R1968 VSS.n206 VSS.n205 163.367
R1969 VSS.n202 VSS.n201 163.367
R1970 VSS.n198 VSS.n197 163.367
R1971 VSS.n194 VSS.n193 163.367
R1972 VSS.n190 VSS.n189 163.367
R1973 VSS.n186 VSS.n185 163.367
R1974 VSS.n182 VSS.n181 163.367
R1975 VSS.n178 VSS.n177 163.367
R1976 VSS.n174 VSS.n173 163.367
R1977 VSS.n170 VSS.n169 163.367
R1978 VSS.n166 VSS.n165 163.367
R1979 VSS.n162 VSS.n154 163.367
R1980 VSS.n777 VSS.n776 163.367
R1981 VSS.n774 VSS.n499 163.367
R1982 VSS.n770 VSS.n769 163.367
R1983 VSS.n767 VSS.n502 163.367
R1984 VSS.n763 VSS.n762 163.367
R1985 VSS.n760 VSS.n505 163.367
R1986 VSS.n756 VSS.n755 163.367
R1987 VSS.n753 VSS.n508 163.367
R1988 VSS.n749 VSS.n748 163.367
R1989 VSS.n746 VSS.n511 163.367
R1990 VSS.n742 VSS.n741 163.367
R1991 VSS.n739 VSS.n514 163.367
R1992 VSS.n735 VSS.n734 163.367
R1993 VSS.n732 VSS.n517 163.367
R1994 VSS.n728 VSS.n727 163.367
R1995 VSS.n725 VSS.n520 163.367
R1996 VSS.n721 VSS.n720 163.367
R1997 VSS.n718 VSS.n523 163.367
R1998 VSS.n714 VSS.n713 163.367
R1999 VSS.n711 VSS.n526 163.367
R2000 VSS.n707 VSS.n706 163.367
R2001 VSS.n704 VSS.n529 163.367
R2002 VSS.n700 VSS.n699 163.367
R2003 VSS.n697 VSS.n532 163.367
R2004 VSS.n693 VSS.n692 163.367
R2005 VSS.n690 VSS.n535 163.367
R2006 VSS.n686 VSS.n685 163.367
R2007 VSS.n683 VSS.n541 163.367
R2008 VSS.n679 VSS.n678 163.367
R2009 VSS.n676 VSS.n544 163.367
R2010 VSS.n672 VSS.n671 163.367
R2011 VSS.n669 VSS.n547 163.367
R2012 VSS.n665 VSS.n664 163.367
R2013 VSS.n662 VSS.n550 163.367
R2014 VSS.n658 VSS.n657 163.367
R2015 VSS.n655 VSS.n553 163.367
R2016 VSS.n651 VSS.n650 163.367
R2017 VSS.n648 VSS.n556 163.367
R2018 VSS.n644 VSS.n643 163.367
R2019 VSS.n641 VSS.n559 163.367
R2020 VSS.n637 VSS.n636 163.367
R2021 VSS.n634 VSS.n562 163.367
R2022 VSS.n630 VSS.n629 163.367
R2023 VSS.n627 VSS.n565 163.367
R2024 VSS.n623 VSS.n622 163.367
R2025 VSS.n620 VSS.n568 163.367
R2026 VSS.n616 VSS.n615 163.367
R2027 VSS.n613 VSS.n571 163.367
R2028 VSS.n609 VSS.n608 163.367
R2029 VSS.n606 VSS.n574 163.367
R2030 VSS.n602 VSS.n601 163.367
R2031 VSS.n599 VSS.n577 163.367
R2032 VSS.n595 VSS.n594 163.367
R2033 VSS.n592 VSS.n580 163.367
R2034 VSS.n587 VSS.n586 163.367
R2035 VSS.n536 VSS.t17 110.374
R2036 VSS.n581 VSS.t14 110.374
R2037 VSS.n158 VSS.t11 110.374
R2038 VSS.n156 VSS.t8 110.374
R2039 VSS.n380 VSS.n94 86.7054
R2040 VSS.n783 VSS.n26 86.7054
R2041 VSS.n537 VSS.t18 72.3613
R2042 VSS.n582 VSS.t15 72.3613
R2043 VSS.n159 VSS.t10 72.3613
R2044 VSS.n157 VSS.t7 72.3613
R2045 VSS.n382 VSS.n381 71.676
R2046 VSS.n155 VSS.n100 71.676
R2047 VSS.n374 VSS.n101 71.676
R2048 VSS.n370 VSS.n102 71.676
R2049 VSS.n366 VSS.n103 71.676
R2050 VSS.n362 VSS.n104 71.676
R2051 VSS.n358 VSS.n105 71.676
R2052 VSS.n354 VSS.n106 71.676
R2053 VSS.n350 VSS.n107 71.676
R2054 VSS.n346 VSS.n108 71.676
R2055 VSS.n342 VSS.n109 71.676
R2056 VSS.n338 VSS.n110 71.676
R2057 VSS.n334 VSS.n111 71.676
R2058 VSS.n330 VSS.n112 71.676
R2059 VSS.n326 VSS.n113 71.676
R2060 VSS.n322 VSS.n114 71.676
R2061 VSS.n318 VSS.n115 71.676
R2062 VSS.n314 VSS.n116 71.676
R2063 VSS.n310 VSS.n117 71.676
R2064 VSS.n306 VSS.n118 71.676
R2065 VSS.n302 VSS.n119 71.676
R2066 VSS.n298 VSS.n120 71.676
R2067 VSS.n294 VSS.n121 71.676
R2068 VSS.n290 VSS.n122 71.676
R2069 VSS.n286 VSS.n123 71.676
R2070 VSS.n282 VSS.n124 71.676
R2071 VSS.n278 VSS.n125 71.676
R2072 VSS.n273 VSS.n126 71.676
R2073 VSS.n269 VSS.n127 71.676
R2074 VSS.n265 VSS.n128 71.676
R2075 VSS.n261 VSS.n129 71.676
R2076 VSS.n257 VSS.n130 71.676
R2077 VSS.n253 VSS.n131 71.676
R2078 VSS.n249 VSS.n132 71.676
R2079 VSS.n245 VSS.n133 71.676
R2080 VSS.n241 VSS.n134 71.676
R2081 VSS.n237 VSS.n135 71.676
R2082 VSS.n233 VSS.n136 71.676
R2083 VSS.n229 VSS.n137 71.676
R2084 VSS.n225 VSS.n138 71.676
R2085 VSS.n221 VSS.n139 71.676
R2086 VSS.n217 VSS.n140 71.676
R2087 VSS.n213 VSS.n141 71.676
R2088 VSS.n209 VSS.n142 71.676
R2089 VSS.n205 VSS.n143 71.676
R2090 VSS.n201 VSS.n144 71.676
R2091 VSS.n197 VSS.n145 71.676
R2092 VSS.n193 VSS.n146 71.676
R2093 VSS.n189 VSS.n147 71.676
R2094 VSS.n185 VSS.n148 71.676
R2095 VSS.n181 VSS.n149 71.676
R2096 VSS.n177 VSS.n150 71.676
R2097 VSS.n173 VSS.n151 71.676
R2098 VSS.n169 VSS.n152 71.676
R2099 VSS.n165 VSS.n153 71.676
R2100 VSS.n777 VSS.n498 71.676
R2101 VSS.n775 VSS.n774 71.676
R2102 VSS.n770 VSS.n501 71.676
R2103 VSS.n768 VSS.n767 71.676
R2104 VSS.n763 VSS.n504 71.676
R2105 VSS.n761 VSS.n760 71.676
R2106 VSS.n756 VSS.n507 71.676
R2107 VSS.n754 VSS.n753 71.676
R2108 VSS.n749 VSS.n510 71.676
R2109 VSS.n747 VSS.n746 71.676
R2110 VSS.n742 VSS.n513 71.676
R2111 VSS.n740 VSS.n739 71.676
R2112 VSS.n735 VSS.n516 71.676
R2113 VSS.n733 VSS.n732 71.676
R2114 VSS.n728 VSS.n519 71.676
R2115 VSS.n726 VSS.n725 71.676
R2116 VSS.n721 VSS.n522 71.676
R2117 VSS.n719 VSS.n718 71.676
R2118 VSS.n714 VSS.n525 71.676
R2119 VSS.n712 VSS.n711 71.676
R2120 VSS.n707 VSS.n528 71.676
R2121 VSS.n705 VSS.n704 71.676
R2122 VSS.n700 VSS.n531 71.676
R2123 VSS.n698 VSS.n697 71.676
R2124 VSS.n693 VSS.n534 71.676
R2125 VSS.n691 VSS.n690 71.676
R2126 VSS.n686 VSS.n539 71.676
R2127 VSS.n684 VSS.n683 71.676
R2128 VSS.n679 VSS.n543 71.676
R2129 VSS.n677 VSS.n676 71.676
R2130 VSS.n672 VSS.n546 71.676
R2131 VSS.n670 VSS.n669 71.676
R2132 VSS.n665 VSS.n549 71.676
R2133 VSS.n663 VSS.n662 71.676
R2134 VSS.n658 VSS.n552 71.676
R2135 VSS.n656 VSS.n655 71.676
R2136 VSS.n651 VSS.n555 71.676
R2137 VSS.n649 VSS.n648 71.676
R2138 VSS.n644 VSS.n558 71.676
R2139 VSS.n642 VSS.n641 71.676
R2140 VSS.n637 VSS.n561 71.676
R2141 VSS.n635 VSS.n634 71.676
R2142 VSS.n630 VSS.n564 71.676
R2143 VSS.n628 VSS.n627 71.676
R2144 VSS.n623 VSS.n567 71.676
R2145 VSS.n621 VSS.n620 71.676
R2146 VSS.n616 VSS.n570 71.676
R2147 VSS.n614 VSS.n613 71.676
R2148 VSS.n609 VSS.n573 71.676
R2149 VSS.n607 VSS.n606 71.676
R2150 VSS.n602 VSS.n576 71.676
R2151 VSS.n600 VSS.n599 71.676
R2152 VSS.n595 VSS.n579 71.676
R2153 VSS.n593 VSS.n592 71.676
R2154 VSS.n587 VSS.n584 71.676
R2155 VSS.n585 VSS.n24 71.676
R2156 VSS.n586 VSS.n585 71.676
R2157 VSS.n584 VSS.n580 71.676
R2158 VSS.n594 VSS.n593 71.676
R2159 VSS.n579 VSS.n577 71.676
R2160 VSS.n601 VSS.n600 71.676
R2161 VSS.n576 VSS.n574 71.676
R2162 VSS.n608 VSS.n607 71.676
R2163 VSS.n573 VSS.n571 71.676
R2164 VSS.n615 VSS.n614 71.676
R2165 VSS.n570 VSS.n568 71.676
R2166 VSS.n622 VSS.n621 71.676
R2167 VSS.n567 VSS.n565 71.676
R2168 VSS.n629 VSS.n628 71.676
R2169 VSS.n564 VSS.n562 71.676
R2170 VSS.n636 VSS.n635 71.676
R2171 VSS.n561 VSS.n559 71.676
R2172 VSS.n643 VSS.n642 71.676
R2173 VSS.n558 VSS.n556 71.676
R2174 VSS.n650 VSS.n649 71.676
R2175 VSS.n555 VSS.n553 71.676
R2176 VSS.n657 VSS.n656 71.676
R2177 VSS.n552 VSS.n550 71.676
R2178 VSS.n664 VSS.n663 71.676
R2179 VSS.n549 VSS.n547 71.676
R2180 VSS.n671 VSS.n670 71.676
R2181 VSS.n546 VSS.n544 71.676
R2182 VSS.n678 VSS.n677 71.676
R2183 VSS.n543 VSS.n541 71.676
R2184 VSS.n685 VSS.n684 71.676
R2185 VSS.n539 VSS.n535 71.676
R2186 VSS.n692 VSS.n691 71.676
R2187 VSS.n534 VSS.n532 71.676
R2188 VSS.n699 VSS.n698 71.676
R2189 VSS.n531 VSS.n529 71.676
R2190 VSS.n706 VSS.n705 71.676
R2191 VSS.n528 VSS.n526 71.676
R2192 VSS.n713 VSS.n712 71.676
R2193 VSS.n525 VSS.n523 71.676
R2194 VSS.n720 VSS.n719 71.676
R2195 VSS.n522 VSS.n520 71.676
R2196 VSS.n727 VSS.n726 71.676
R2197 VSS.n519 VSS.n517 71.676
R2198 VSS.n734 VSS.n733 71.676
R2199 VSS.n516 VSS.n514 71.676
R2200 VSS.n741 VSS.n740 71.676
R2201 VSS.n513 VSS.n511 71.676
R2202 VSS.n748 VSS.n747 71.676
R2203 VSS.n510 VSS.n508 71.676
R2204 VSS.n755 VSS.n754 71.676
R2205 VSS.n507 VSS.n505 71.676
R2206 VSS.n762 VSS.n761 71.676
R2207 VSS.n504 VSS.n502 71.676
R2208 VSS.n769 VSS.n768 71.676
R2209 VSS.n501 VSS.n499 71.676
R2210 VSS.n776 VSS.n775 71.676
R2211 VSS.n498 VSS.n28 71.676
R2212 VSS.n381 VSS.n99 71.676
R2213 VSS.n375 VSS.n100 71.676
R2214 VSS.n371 VSS.n101 71.676
R2215 VSS.n367 VSS.n102 71.676
R2216 VSS.n363 VSS.n103 71.676
R2217 VSS.n359 VSS.n104 71.676
R2218 VSS.n355 VSS.n105 71.676
R2219 VSS.n351 VSS.n106 71.676
R2220 VSS.n347 VSS.n107 71.676
R2221 VSS.n343 VSS.n108 71.676
R2222 VSS.n339 VSS.n109 71.676
R2223 VSS.n335 VSS.n110 71.676
R2224 VSS.n331 VSS.n111 71.676
R2225 VSS.n327 VSS.n112 71.676
R2226 VSS.n323 VSS.n113 71.676
R2227 VSS.n319 VSS.n114 71.676
R2228 VSS.n315 VSS.n115 71.676
R2229 VSS.n311 VSS.n116 71.676
R2230 VSS.n307 VSS.n117 71.676
R2231 VSS.n303 VSS.n118 71.676
R2232 VSS.n299 VSS.n119 71.676
R2233 VSS.n295 VSS.n120 71.676
R2234 VSS.n291 VSS.n121 71.676
R2235 VSS.n287 VSS.n122 71.676
R2236 VSS.n283 VSS.n123 71.676
R2237 VSS.n279 VSS.n124 71.676
R2238 VSS.n274 VSS.n125 71.676
R2239 VSS.n270 VSS.n126 71.676
R2240 VSS.n266 VSS.n127 71.676
R2241 VSS.n262 VSS.n128 71.676
R2242 VSS.n258 VSS.n129 71.676
R2243 VSS.n254 VSS.n130 71.676
R2244 VSS.n250 VSS.n131 71.676
R2245 VSS.n246 VSS.n132 71.676
R2246 VSS.n242 VSS.n133 71.676
R2247 VSS.n238 VSS.n134 71.676
R2248 VSS.n234 VSS.n135 71.676
R2249 VSS.n230 VSS.n136 71.676
R2250 VSS.n226 VSS.n137 71.676
R2251 VSS.n222 VSS.n138 71.676
R2252 VSS.n218 VSS.n139 71.676
R2253 VSS.n214 VSS.n140 71.676
R2254 VSS.n210 VSS.n141 71.676
R2255 VSS.n206 VSS.n142 71.676
R2256 VSS.n202 VSS.n143 71.676
R2257 VSS.n198 VSS.n144 71.676
R2258 VSS.n194 VSS.n145 71.676
R2259 VSS.n190 VSS.n146 71.676
R2260 VSS.n186 VSS.n147 71.676
R2261 VSS.n182 VSS.n148 71.676
R2262 VSS.n178 VSS.n149 71.676
R2263 VSS.n174 VSS.n150 71.676
R2264 VSS.n170 VSS.n151 71.676
R2265 VSS.n166 VSS.n152 71.676
R2266 VSS.n162 VSS.n153 71.676
R2267 VSS.n388 VSS.n94 54.877
R2268 VSS.n388 VSS.n95 54.877
R2269 VSS.n396 VSS.n83 54.877
R2270 VSS.n404 VSS.n83 54.877
R2271 VSS.n404 VSS.n77 54.877
R2272 VSS.n413 VSS.n77 54.877
R2273 VSS.n413 VSS.n412 54.877
R2274 VSS.n421 VSS.n66 54.877
R2275 VSS.n430 VSS.n66 54.877
R2276 VSS.n430 VSS.n429 54.877
R2277 VSS.n438 VSS.n55 54.877
R2278 VSS.n448 VSS.n55 54.877
R2279 VSS.n448 VSS.n447 54.877
R2280 VSS.n457 VSS.n456 54.877
R2281 VSS.n460 VSS.n457 54.877
R2282 VSS.n460 VSS.n459 54.877
R2283 VSS.n469 VSS.n468 54.877
R2284 VSS.n472 VSS.n469 54.877
R2285 VSS.n472 VSS.n471 54.877
R2286 VSS.n481 VSS.n480 54.877
R2287 VSS.n482 VSS.n481 54.877
R2288 VSS.n482 VSS.n34 54.877
R2289 VSS.n490 VSS.n34 54.877
R2290 VSS.n491 VSS.n490 54.877
R2291 VSS.n492 VSS.n25 54.877
R2292 VSS.n783 VSS.n25 54.877
R2293 VSS.n537 VSS.n536 38.0126
R2294 VSS.n582 VSS.n581 38.0126
R2295 VSS.n159 VSS.n158 38.0126
R2296 VSS.n157 VSS.n156 38.0126
R2297 VSS.n412 VSS.t1 36.219
R2298 VSS.n480 VSS.t4 36.219
R2299 VSS.n538 VSS.n537 34.3278
R2300 VSS.n589 VSS.n582 34.3278
R2301 VSS.n160 VSS.n159 34.3278
R2302 VSS.n276 VSS.n157 34.3278
R2303 VSS.n429 VSS.t2 31.8289
R2304 VSS.n468 VSS.t0 31.8289
R2305 VSS.n95 VSS.t6 30.7314
R2306 VSS.n492 VSS.t13 30.7314
R2307 VSS.n447 VSS.t3 27.4388
R2308 VSS.n456 VSS.t3 27.4388
R2309 VSS.n780 VSS.n779 26.7121
R2310 VSS.n786 VSS.n22 26.7121
R2311 VSS.n384 VSS.n383 26.7121
R2312 VSS.n161 VSS.n91 26.7121
R2313 VSS.n396 VSS.t6 24.1462
R2314 VSS.t13 VSS.n491 24.1462
R2315 VSS.n438 VSS.t2 23.0486
R2316 VSS.n459 VSS.t0 23.0486
R2317 VSS.n386 VSS.n97 19.3944
R2318 VSS.n386 VSS.n87 19.3944
R2319 VSS.n398 VSS.n87 19.3944
R2320 VSS.n398 VSS.n85 19.3944
R2321 VSS.n402 VSS.n85 19.3944
R2322 VSS.n402 VSS.n75 19.3944
R2323 VSS.n415 VSS.n75 19.3944
R2324 VSS.n415 VSS.n73 19.3944
R2325 VSS.n419 VSS.n73 19.3944
R2326 VSS.n419 VSS.n64 19.3944
R2327 VSS.n432 VSS.n64 19.3944
R2328 VSS.n432 VSS.n62 19.3944
R2329 VSS.n436 VSS.n62 19.3944
R2330 VSS.n436 VSS.n53 19.3944
R2331 VSS.n450 VSS.n53 19.3944
R2332 VSS.n450 VSS.n51 19.3944
R2333 VSS.n454 VSS.n51 19.3944
R2334 VSS.n454 VSS.n48 19.3944
R2335 VSS.n462 VSS.n48 19.3944
R2336 VSS.n462 VSS.n46 19.3944
R2337 VSS.n466 VSS.n46 19.3944
R2338 VSS.n466 VSS.n43 19.3944
R2339 VSS.n474 VSS.n43 19.3944
R2340 VSS.n474 VSS.n41 19.3944
R2341 VSS.n478 VSS.n41 19.3944
R2342 VSS.n478 VSS.n38 19.3944
R2343 VSS.n484 VSS.n38 19.3944
R2344 VSS.n484 VSS.n36 19.3944
R2345 VSS.n488 VSS.n36 19.3944
R2346 VSS.n488 VSS.n31 19.3944
R2347 VSS.n494 VSS.n31 19.3944
R2348 VSS.n494 VSS.n29 19.3944
R2349 VSS.n781 VSS.n29 19.3944
R2350 VSS.n390 VSS.n92 19.3944
R2351 VSS.n390 VSS.n90 19.3944
R2352 VSS.n394 VSS.n90 19.3944
R2353 VSS.n394 VSS.n81 19.3944
R2354 VSS.n406 VSS.n81 19.3944
R2355 VSS.n406 VSS.n79 19.3944
R2356 VSS.n410 VSS.n79 19.3944
R2357 VSS.n410 VSS.n70 19.3944
R2358 VSS.n423 VSS.n70 19.3944
R2359 VSS.n423 VSS.n68 19.3944
R2360 VSS.n427 VSS.n68 19.3944
R2361 VSS.n427 VSS.n59 19.3944
R2362 VSS.n440 VSS.n59 19.3944
R2363 VSS.n440 VSS.n57 19.3944
R2364 VSS.n444 VSS.n57 19.3944
R2365 VSS.n444 VSS.n2 19.3944
R2366 VSS.n809 VSS.n2 19.3944
R2367 VSS.n809 VSS.n808 19.3944
R2368 VSS.n808 VSS.n807 19.3944
R2369 VSS.n807 VSS.n6 19.3944
R2370 VSS.n803 VSS.n6 19.3944
R2371 VSS.n803 VSS.n802 19.3944
R2372 VSS.n802 VSS.n801 19.3944
R2373 VSS.n801 VSS.n11 19.3944
R2374 VSS.n797 VSS.n11 19.3944
R2375 VSS.n797 VSS.n796 19.3944
R2376 VSS.n796 VSS.n795 19.3944
R2377 VSS.n795 VSS.n16 19.3944
R2378 VSS.n791 VSS.n16 19.3944
R2379 VSS.n791 VSS.n790 19.3944
R2380 VSS.n790 VSS.n789 19.3944
R2381 VSS.n789 VSS.n21 19.3944
R2382 VSS.n785 VSS.n21 19.3944
R2383 VSS.n421 VSS.t1 18.6585
R2384 VSS.n471 VSS.t4 18.6585
R2385 VSS.n779 VSS.n778 10.6151
R2386 VSS.n778 VSS.n497 10.6151
R2387 VSS.n773 VSS.n497 10.6151
R2388 VSS.n773 VSS.n772 10.6151
R2389 VSS.n772 VSS.n771 10.6151
R2390 VSS.n771 VSS.n500 10.6151
R2391 VSS.n766 VSS.n500 10.6151
R2392 VSS.n766 VSS.n765 10.6151
R2393 VSS.n765 VSS.n764 10.6151
R2394 VSS.n764 VSS.n503 10.6151
R2395 VSS.n759 VSS.n503 10.6151
R2396 VSS.n759 VSS.n758 10.6151
R2397 VSS.n758 VSS.n757 10.6151
R2398 VSS.n757 VSS.n506 10.6151
R2399 VSS.n752 VSS.n506 10.6151
R2400 VSS.n752 VSS.n751 10.6151
R2401 VSS.n751 VSS.n750 10.6151
R2402 VSS.n750 VSS.n509 10.6151
R2403 VSS.n745 VSS.n509 10.6151
R2404 VSS.n745 VSS.n744 10.6151
R2405 VSS.n744 VSS.n743 10.6151
R2406 VSS.n743 VSS.n512 10.6151
R2407 VSS.n738 VSS.n512 10.6151
R2408 VSS.n738 VSS.n737 10.6151
R2409 VSS.n737 VSS.n736 10.6151
R2410 VSS.n736 VSS.n515 10.6151
R2411 VSS.n731 VSS.n515 10.6151
R2412 VSS.n731 VSS.n730 10.6151
R2413 VSS.n730 VSS.n729 10.6151
R2414 VSS.n729 VSS.n518 10.6151
R2415 VSS.n724 VSS.n518 10.6151
R2416 VSS.n724 VSS.n723 10.6151
R2417 VSS.n723 VSS.n722 10.6151
R2418 VSS.n722 VSS.n521 10.6151
R2419 VSS.n717 VSS.n521 10.6151
R2420 VSS.n717 VSS.n716 10.6151
R2421 VSS.n716 VSS.n715 10.6151
R2422 VSS.n715 VSS.n524 10.6151
R2423 VSS.n710 VSS.n524 10.6151
R2424 VSS.n710 VSS.n709 10.6151
R2425 VSS.n709 VSS.n708 10.6151
R2426 VSS.n708 VSS.n527 10.6151
R2427 VSS.n703 VSS.n527 10.6151
R2428 VSS.n703 VSS.n702 10.6151
R2429 VSS.n702 VSS.n701 10.6151
R2430 VSS.n701 VSS.n530 10.6151
R2431 VSS.n696 VSS.n530 10.6151
R2432 VSS.n696 VSS.n695 10.6151
R2433 VSS.n695 VSS.n694 10.6151
R2434 VSS.n694 VSS.n533 10.6151
R2435 VSS.n689 VSS.n533 10.6151
R2436 VSS.n689 VSS.n688 10.6151
R2437 VSS.n688 VSS.n687 10.6151
R2438 VSS.n682 VSS.n540 10.6151
R2439 VSS.n682 VSS.n681 10.6151
R2440 VSS.n681 VSS.n680 10.6151
R2441 VSS.n680 VSS.n542 10.6151
R2442 VSS.n675 VSS.n542 10.6151
R2443 VSS.n675 VSS.n674 10.6151
R2444 VSS.n674 VSS.n673 10.6151
R2445 VSS.n673 VSS.n545 10.6151
R2446 VSS.n668 VSS.n545 10.6151
R2447 VSS.n668 VSS.n667 10.6151
R2448 VSS.n667 VSS.n666 10.6151
R2449 VSS.n666 VSS.n548 10.6151
R2450 VSS.n661 VSS.n548 10.6151
R2451 VSS.n661 VSS.n660 10.6151
R2452 VSS.n660 VSS.n659 10.6151
R2453 VSS.n659 VSS.n551 10.6151
R2454 VSS.n654 VSS.n551 10.6151
R2455 VSS.n654 VSS.n653 10.6151
R2456 VSS.n653 VSS.n652 10.6151
R2457 VSS.n652 VSS.n554 10.6151
R2458 VSS.n647 VSS.n554 10.6151
R2459 VSS.n647 VSS.n646 10.6151
R2460 VSS.n646 VSS.n645 10.6151
R2461 VSS.n645 VSS.n557 10.6151
R2462 VSS.n640 VSS.n557 10.6151
R2463 VSS.n640 VSS.n639 10.6151
R2464 VSS.n639 VSS.n638 10.6151
R2465 VSS.n638 VSS.n560 10.6151
R2466 VSS.n633 VSS.n560 10.6151
R2467 VSS.n633 VSS.n632 10.6151
R2468 VSS.n632 VSS.n631 10.6151
R2469 VSS.n631 VSS.n563 10.6151
R2470 VSS.n626 VSS.n563 10.6151
R2471 VSS.n626 VSS.n625 10.6151
R2472 VSS.n625 VSS.n624 10.6151
R2473 VSS.n624 VSS.n566 10.6151
R2474 VSS.n619 VSS.n566 10.6151
R2475 VSS.n619 VSS.n618 10.6151
R2476 VSS.n618 VSS.n617 10.6151
R2477 VSS.n617 VSS.n569 10.6151
R2478 VSS.n612 VSS.n569 10.6151
R2479 VSS.n612 VSS.n611 10.6151
R2480 VSS.n611 VSS.n610 10.6151
R2481 VSS.n610 VSS.n572 10.6151
R2482 VSS.n605 VSS.n572 10.6151
R2483 VSS.n605 VSS.n604 10.6151
R2484 VSS.n604 VSS.n603 10.6151
R2485 VSS.n603 VSS.n575 10.6151
R2486 VSS.n598 VSS.n575 10.6151
R2487 VSS.n598 VSS.n597 10.6151
R2488 VSS.n597 VSS.n596 10.6151
R2489 VSS.n596 VSS.n578 10.6151
R2490 VSS.n591 VSS.n578 10.6151
R2491 VSS.n591 VSS.n590 10.6151
R2492 VSS.n588 VSS.n583 10.6151
R2493 VSS.n583 VSS.n22 10.6151
R2494 VSS.n383 VSS.n98 10.6151
R2495 VSS.n378 VSS.n98 10.6151
R2496 VSS.n378 VSS.n377 10.6151
R2497 VSS.n377 VSS.n376 10.6151
R2498 VSS.n376 VSS.n373 10.6151
R2499 VSS.n373 VSS.n372 10.6151
R2500 VSS.n372 VSS.n369 10.6151
R2501 VSS.n369 VSS.n368 10.6151
R2502 VSS.n368 VSS.n365 10.6151
R2503 VSS.n365 VSS.n364 10.6151
R2504 VSS.n364 VSS.n361 10.6151
R2505 VSS.n361 VSS.n360 10.6151
R2506 VSS.n360 VSS.n357 10.6151
R2507 VSS.n357 VSS.n356 10.6151
R2508 VSS.n356 VSS.n353 10.6151
R2509 VSS.n353 VSS.n352 10.6151
R2510 VSS.n352 VSS.n349 10.6151
R2511 VSS.n349 VSS.n348 10.6151
R2512 VSS.n348 VSS.n345 10.6151
R2513 VSS.n345 VSS.n344 10.6151
R2514 VSS.n344 VSS.n341 10.6151
R2515 VSS.n341 VSS.n340 10.6151
R2516 VSS.n340 VSS.n337 10.6151
R2517 VSS.n337 VSS.n336 10.6151
R2518 VSS.n336 VSS.n333 10.6151
R2519 VSS.n333 VSS.n332 10.6151
R2520 VSS.n332 VSS.n329 10.6151
R2521 VSS.n329 VSS.n328 10.6151
R2522 VSS.n328 VSS.n325 10.6151
R2523 VSS.n325 VSS.n324 10.6151
R2524 VSS.n324 VSS.n321 10.6151
R2525 VSS.n321 VSS.n320 10.6151
R2526 VSS.n320 VSS.n317 10.6151
R2527 VSS.n317 VSS.n316 10.6151
R2528 VSS.n316 VSS.n313 10.6151
R2529 VSS.n313 VSS.n312 10.6151
R2530 VSS.n312 VSS.n309 10.6151
R2531 VSS.n309 VSS.n308 10.6151
R2532 VSS.n308 VSS.n305 10.6151
R2533 VSS.n305 VSS.n304 10.6151
R2534 VSS.n304 VSS.n301 10.6151
R2535 VSS.n301 VSS.n300 10.6151
R2536 VSS.n300 VSS.n297 10.6151
R2537 VSS.n297 VSS.n296 10.6151
R2538 VSS.n296 VSS.n293 10.6151
R2539 VSS.n293 VSS.n292 10.6151
R2540 VSS.n292 VSS.n289 10.6151
R2541 VSS.n289 VSS.n288 10.6151
R2542 VSS.n288 VSS.n285 10.6151
R2543 VSS.n285 VSS.n284 10.6151
R2544 VSS.n284 VSS.n281 10.6151
R2545 VSS.n281 VSS.n280 10.6151
R2546 VSS.n280 VSS.n277 10.6151
R2547 VSS.n275 VSS.n272 10.6151
R2548 VSS.n272 VSS.n271 10.6151
R2549 VSS.n271 VSS.n268 10.6151
R2550 VSS.n268 VSS.n267 10.6151
R2551 VSS.n267 VSS.n264 10.6151
R2552 VSS.n264 VSS.n263 10.6151
R2553 VSS.n263 VSS.n260 10.6151
R2554 VSS.n260 VSS.n259 10.6151
R2555 VSS.n259 VSS.n256 10.6151
R2556 VSS.n256 VSS.n255 10.6151
R2557 VSS.n255 VSS.n252 10.6151
R2558 VSS.n252 VSS.n251 10.6151
R2559 VSS.n251 VSS.n248 10.6151
R2560 VSS.n248 VSS.n247 10.6151
R2561 VSS.n247 VSS.n244 10.6151
R2562 VSS.n244 VSS.n243 10.6151
R2563 VSS.n243 VSS.n240 10.6151
R2564 VSS.n240 VSS.n239 10.6151
R2565 VSS.n239 VSS.n236 10.6151
R2566 VSS.n236 VSS.n235 10.6151
R2567 VSS.n235 VSS.n232 10.6151
R2568 VSS.n232 VSS.n231 10.6151
R2569 VSS.n231 VSS.n228 10.6151
R2570 VSS.n228 VSS.n227 10.6151
R2571 VSS.n227 VSS.n224 10.6151
R2572 VSS.n224 VSS.n223 10.6151
R2573 VSS.n223 VSS.n220 10.6151
R2574 VSS.n220 VSS.n219 10.6151
R2575 VSS.n219 VSS.n216 10.6151
R2576 VSS.n216 VSS.n215 10.6151
R2577 VSS.n215 VSS.n212 10.6151
R2578 VSS.n212 VSS.n211 10.6151
R2579 VSS.n211 VSS.n208 10.6151
R2580 VSS.n208 VSS.n207 10.6151
R2581 VSS.n207 VSS.n204 10.6151
R2582 VSS.n204 VSS.n203 10.6151
R2583 VSS.n203 VSS.n200 10.6151
R2584 VSS.n200 VSS.n199 10.6151
R2585 VSS.n199 VSS.n196 10.6151
R2586 VSS.n196 VSS.n195 10.6151
R2587 VSS.n195 VSS.n192 10.6151
R2588 VSS.n192 VSS.n191 10.6151
R2589 VSS.n191 VSS.n188 10.6151
R2590 VSS.n188 VSS.n187 10.6151
R2591 VSS.n187 VSS.n184 10.6151
R2592 VSS.n184 VSS.n183 10.6151
R2593 VSS.n183 VSS.n180 10.6151
R2594 VSS.n180 VSS.n179 10.6151
R2595 VSS.n179 VSS.n176 10.6151
R2596 VSS.n176 VSS.n175 10.6151
R2597 VSS.n175 VSS.n172 10.6151
R2598 VSS.n172 VSS.n171 10.6151
R2599 VSS.n171 VSS.n168 10.6151
R2600 VSS.n168 VSS.n167 10.6151
R2601 VSS.n164 VSS.n163 10.6151
R2602 VSS.n163 VSS.n161 10.6151
R2603 VSS.n540 VSS.n538 9.83465
R2604 VSS.n276 VSS.n275 9.83465
R2605 VSS.n808 VSS.n0 9.3005
R2606 VSS.n807 VSS.n806 9.3005
R2607 VSS.n805 VSS.n6 9.3005
R2608 VSS.n804 VSS.n803 9.3005
R2609 VSS.n802 VSS.n7 9.3005
R2610 VSS.n801 VSS.n800 9.3005
R2611 VSS.n799 VSS.n11 9.3005
R2612 VSS.n798 VSS.n797 9.3005
R2613 VSS.n796 VSS.n12 9.3005
R2614 VSS.n795 VSS.n794 9.3005
R2615 VSS.n793 VSS.n16 9.3005
R2616 VSS.n792 VSS.n791 9.3005
R2617 VSS.n790 VSS.n17 9.3005
R2618 VSS.n789 VSS.n788 9.3005
R2619 VSS.n787 VSS.n21 9.3005
R2620 VSS.n786 VSS.n785 9.3005
R2621 VSS.n384 VSS.n97 9.3005
R2622 VSS.n386 VSS.n385 9.3005
R2623 VSS.n87 VSS.n86 9.3005
R2624 VSS.n399 VSS.n398 9.3005
R2625 VSS.n400 VSS.n85 9.3005
R2626 VSS.n402 VSS.n401 9.3005
R2627 VSS.n75 VSS.n74 9.3005
R2628 VSS.n416 VSS.n415 9.3005
R2629 VSS.n417 VSS.n73 9.3005
R2630 VSS.n419 VSS.n418 9.3005
R2631 VSS.n64 VSS.n63 9.3005
R2632 VSS.n433 VSS.n432 9.3005
R2633 VSS.n434 VSS.n62 9.3005
R2634 VSS.n436 VSS.n435 9.3005
R2635 VSS.n53 VSS.n52 9.3005
R2636 VSS.n451 VSS.n450 9.3005
R2637 VSS.n452 VSS.n51 9.3005
R2638 VSS.n454 VSS.n453 9.3005
R2639 VSS.n48 VSS.n47 9.3005
R2640 VSS.n463 VSS.n462 9.3005
R2641 VSS.n464 VSS.n46 9.3005
R2642 VSS.n466 VSS.n465 9.3005
R2643 VSS.n43 VSS.n42 9.3005
R2644 VSS.n475 VSS.n474 9.3005
R2645 VSS.n476 VSS.n41 9.3005
R2646 VSS.n478 VSS.n477 9.3005
R2647 VSS.n38 VSS.n37 9.3005
R2648 VSS.n485 VSS.n484 9.3005
R2649 VSS.n486 VSS.n36 9.3005
R2650 VSS.n488 VSS.n487 9.3005
R2651 VSS.n31 VSS.n30 9.3005
R2652 VSS.n495 VSS.n494 9.3005
R2653 VSS.n496 VSS.n29 9.3005
R2654 VSS.n781 VSS.n780 9.3005
R2655 VSS.n391 VSS.n390 9.3005
R2656 VSS.n392 VSS.n90 9.3005
R2657 VSS.n394 VSS.n393 9.3005
R2658 VSS.n81 VSS.n80 9.3005
R2659 VSS.n407 VSS.n406 9.3005
R2660 VSS.n408 VSS.n79 9.3005
R2661 VSS.n410 VSS.n409 9.3005
R2662 VSS.n70 VSS.n69 9.3005
R2663 VSS.n424 VSS.n423 9.3005
R2664 VSS.n425 VSS.n68 9.3005
R2665 VSS.n427 VSS.n426 9.3005
R2666 VSS.n59 VSS.n58 9.3005
R2667 VSS.n441 VSS.n440 9.3005
R2668 VSS.n442 VSS.n57 9.3005
R2669 VSS.n444 VSS.n443 9.3005
R2670 VSS.n2 VSS.n1 9.3005
R2671 VSS.n92 VSS.n91 9.3005
R2672 VSS VSS.n809 9.3005
R2673 VSS.n589 VSS.n588 5.46391
R2674 VSS.n164 VSS.n160 5.46391
R2675 VSS.n590 VSS.n589 5.15172
R2676 VSS.n167 VSS.n160 5.15172
R2677 VSS.n687 VSS.n538 0.780988
R2678 VSS.n277 VSS.n276 0.780988
R2679 VSS VSS.n0 0.152939
R2680 VSS.n806 VSS.n0 0.152939
R2681 VSS.n806 VSS.n805 0.152939
R2682 VSS.n805 VSS.n804 0.152939
R2683 VSS.n804 VSS.n7 0.152939
R2684 VSS.n800 VSS.n7 0.152939
R2685 VSS.n800 VSS.n799 0.152939
R2686 VSS.n799 VSS.n798 0.152939
R2687 VSS.n798 VSS.n12 0.152939
R2688 VSS.n794 VSS.n12 0.152939
R2689 VSS.n794 VSS.n793 0.152939
R2690 VSS.n793 VSS.n792 0.152939
R2691 VSS.n792 VSS.n17 0.152939
R2692 VSS.n788 VSS.n17 0.152939
R2693 VSS.n788 VSS.n787 0.152939
R2694 VSS.n787 VSS.n786 0.152939
R2695 VSS.n385 VSS.n384 0.152939
R2696 VSS.n385 VSS.n86 0.152939
R2697 VSS.n399 VSS.n86 0.152939
R2698 VSS.n400 VSS.n399 0.152939
R2699 VSS.n401 VSS.n400 0.152939
R2700 VSS.n401 VSS.n74 0.152939
R2701 VSS.n416 VSS.n74 0.152939
R2702 VSS.n417 VSS.n416 0.152939
R2703 VSS.n418 VSS.n417 0.152939
R2704 VSS.n418 VSS.n63 0.152939
R2705 VSS.n433 VSS.n63 0.152939
R2706 VSS.n434 VSS.n433 0.152939
R2707 VSS.n435 VSS.n434 0.152939
R2708 VSS.n435 VSS.n52 0.152939
R2709 VSS.n451 VSS.n52 0.152939
R2710 VSS.n452 VSS.n451 0.152939
R2711 VSS.n453 VSS.n452 0.152939
R2712 VSS.n453 VSS.n47 0.152939
R2713 VSS.n463 VSS.n47 0.152939
R2714 VSS.n464 VSS.n463 0.152939
R2715 VSS.n465 VSS.n464 0.152939
R2716 VSS.n465 VSS.n42 0.152939
R2717 VSS.n475 VSS.n42 0.152939
R2718 VSS.n476 VSS.n475 0.152939
R2719 VSS.n477 VSS.n476 0.152939
R2720 VSS.n477 VSS.n37 0.152939
R2721 VSS.n485 VSS.n37 0.152939
R2722 VSS.n486 VSS.n485 0.152939
R2723 VSS.n487 VSS.n486 0.152939
R2724 VSS.n487 VSS.n30 0.152939
R2725 VSS.n495 VSS.n30 0.152939
R2726 VSS.n496 VSS.n495 0.152939
R2727 VSS.n780 VSS.n496 0.152939
R2728 VSS.n391 VSS.n91 0.152939
R2729 VSS.n392 VSS.n391 0.152939
R2730 VSS.n393 VSS.n392 0.152939
R2731 VSS.n393 VSS.n80 0.152939
R2732 VSS.n407 VSS.n80 0.152939
R2733 VSS.n408 VSS.n407 0.152939
R2734 VSS.n409 VSS.n408 0.152939
R2735 VSS.n409 VSS.n69 0.152939
R2736 VSS.n424 VSS.n69 0.152939
R2737 VSS.n425 VSS.n424 0.152939
R2738 VSS.n426 VSS.n425 0.152939
R2739 VSS.n426 VSS.n58 0.152939
R2740 VSS.n441 VSS.n58 0.152939
R2741 VSS.n442 VSS.n441 0.152939
R2742 VSS.n443 VSS.n442 0.152939
R2743 VSS.n443 VSS.n1 0.152939
R2744 VSS VSS.n1 0.1255
R2745 VGN.n36 VGN.t9 278.067
R2746 VGN.n6 VGN.t0 278.067
R2747 VGN.n58 VGN.t3 245.141
R2748 VGN.n51 VGN.t1 245.141
R2749 VGN.n44 VGN.t5 245.141
R2750 VGN.n37 VGN.t7 245.141
R2751 VGN.n7 VGN.t8 245.141
R2752 VGN.n14 VGN.t4 245.141
R2753 VGN.n21 VGN.t2 245.141
R2754 VGN.n28 VGN.t6 245.141
R2755 VGN.n59 VGN.n58 177.531
R2756 VGN.n29 VGN.n28 177.531
R2757 VGN.n27 VGN.n0 161.3
R2758 VGN.n26 VGN.n25 161.3
R2759 VGN.n24 VGN.n1 161.3
R2760 VGN.n23 VGN.n22 161.3
R2761 VGN.n20 VGN.n2 161.3
R2762 VGN.n19 VGN.n18 161.3
R2763 VGN.n17 VGN.n3 161.3
R2764 VGN.n16 VGN.n15 161.3
R2765 VGN.n13 VGN.n4 161.3
R2766 VGN.n12 VGN.n11 161.3
R2767 VGN.n10 VGN.n5 161.3
R2768 VGN.n9 VGN.n8 161.3
R2769 VGN.n39 VGN.n38 161.3
R2770 VGN.n40 VGN.n35 161.3
R2771 VGN.n42 VGN.n41 161.3
R2772 VGN.n43 VGN.n34 161.3
R2773 VGN.n46 VGN.n45 161.3
R2774 VGN.n47 VGN.n33 161.3
R2775 VGN.n49 VGN.n48 161.3
R2776 VGN.n50 VGN.n32 161.3
R2777 VGN.n53 VGN.n52 161.3
R2778 VGN.n54 VGN.n31 161.3
R2779 VGN.n56 VGN.n55 161.3
R2780 VGN.n57 VGN.n30 161.3
R2781 VGN.n56 VGN.n31 56.5617
R2782 VGN.n26 VGN.n1 56.5617
R2783 VGN.n49 VGN.n33 56.5617
R2784 VGN.n42 VGN.n35 56.5617
R2785 VGN.n12 VGN.n5 56.5617
R2786 VGN.n19 VGN.n3 56.5617
R2787 VGN.n37 VGN.n36 56.0889
R2788 VGN.n7 VGN.n6 56.0889
R2789 VGN.n57 VGN.n56 24.5923
R2790 VGN.n52 VGN.n31 24.5923
R2791 VGN.n50 VGN.n49 24.5923
R2792 VGN.n45 VGN.n33 24.5923
R2793 VGN.n43 VGN.n42 24.5923
R2794 VGN.n38 VGN.n35 24.5923
R2795 VGN.n8 VGN.n5 24.5923
R2796 VGN.n15 VGN.n3 24.5923
R2797 VGN.n13 VGN.n12 24.5923
R2798 VGN.n22 VGN.n1 24.5923
R2799 VGN.n20 VGN.n19 24.5923
R2800 VGN.n27 VGN.n26 24.5923
R2801 VGN.n9 VGN.n6 17.9261
R2802 VGN.n39 VGN.n36 17.9261
R2803 VGN VGN.n29 16.9134
R2804 VGN.n52 VGN.n51 14.2638
R2805 VGN.n22 VGN.n21 14.2638
R2806 VGN.n45 VGN.n44 12.2964
R2807 VGN.n44 VGN.n43 12.2964
R2808 VGN.n15 VGN.n14 12.2964
R2809 VGN.n14 VGN.n13 12.2964
R2810 VGN.n51 VGN.n50 10.3291
R2811 VGN.n38 VGN.n37 10.3291
R2812 VGN.n8 VGN.n7 10.3291
R2813 VGN.n21 VGN.n20 10.3291
R2814 VGN.n58 VGN.n57 8.36172
R2815 VGN.n28 VGN.n27 8.36172
R2816 VGN.n29 VGN.n0 0.189894
R2817 VGN.n25 VGN.n0 0.189894
R2818 VGN.n25 VGN.n24 0.189894
R2819 VGN.n24 VGN.n23 0.189894
R2820 VGN.n23 VGN.n2 0.189894
R2821 VGN.n18 VGN.n2 0.189894
R2822 VGN.n18 VGN.n17 0.189894
R2823 VGN.n17 VGN.n16 0.189894
R2824 VGN.n16 VGN.n4 0.189894
R2825 VGN.n11 VGN.n4 0.189894
R2826 VGN.n11 VGN.n10 0.189894
R2827 VGN.n10 VGN.n9 0.189894
R2828 VGN.n59 VGN.n30 0.189894
R2829 VGN.n55 VGN.n30 0.189894
R2830 VGN.n55 VGN.n54 0.189894
R2831 VGN.n54 VGN.n53 0.189894
R2832 VGN.n53 VGN.n32 0.189894
R2833 VGN.n48 VGN.n32 0.189894
R2834 VGN.n48 VGN.n47 0.189894
R2835 VGN.n47 VGN.n46 0.189894
R2836 VGN.n46 VGN.n34 0.189894
R2837 VGN.n41 VGN.n34 0.189894
R2838 VGN.n41 VGN.n40 0.189894
R2839 VGN.n40 VGN.n39 0.189894
R2840 VGN VGN.n59 0.133076
C0 VGN VCC 0.030258f
C1 VGN VOUT 26.322401f
C2 VCC VOUT 18.7081f
C3 VGN VSS 9.645183f
C4 VOUT VSS 18.778307f
C5 VGP VSS 0.119239f
C6 VIN VSS 0.433798f
C7 VCC VSS 57.062347f
C8 VGN.n0 VSS 0.02343f
C9 VGN.t6 VSS 1.73884f
C10 VGN.n1 VSS 0.030169f
C11 VGN.n2 VSS 0.02343f
C12 VGN.t2 VSS 1.73884f
C13 VGN.n3 VSS 0.032762f
C14 VGN.n4 VSS 0.02343f
C15 VGN.t4 VSS 1.73884f
C16 VGN.n5 VSS 0.035355f
C17 VGN.t0 VSS 1.82286f
C18 VGN.n6 VSS 0.670151f
C19 VGN.t8 VSS 1.73884f
C20 VGN.n7 VSS 0.657309f
C21 VGN.n8 VSS 0.031008f
C22 VGN.n9 VSS 0.149969f
C23 VGN.n10 VSS 0.02343f
C24 VGN.n11 VSS 0.02343f
C25 VGN.n12 VSS 0.032762f
C26 VGN.n13 VSS 0.032724f
C27 VGN.n14 VSS 0.612956f
C28 VGN.n15 VSS 0.032724f
C29 VGN.n16 VSS 0.02343f
C30 VGN.n17 VSS 0.02343f
C31 VGN.n18 VSS 0.02343f
C32 VGN.n19 VSS 0.035355f
C33 VGN.n20 VSS 0.031008f
C34 VGN.n21 VSS 0.612956f
C35 VGN.n22 VSS 0.03444f
C36 VGN.n23 VSS 0.02343f
C37 VGN.n24 VSS 0.02343f
C38 VGN.n25 VSS 0.02343f
C39 VGN.n26 VSS 0.037948f
C40 VGN.n27 VSS 0.029292f
C41 VGN.n28 VSS 0.664125f
C42 VGN.n29 VSS 0.348474f
C43 VGN.n30 VSS 0.02343f
C44 VGN.t3 VSS 1.73884f
C45 VGN.n31 VSS 0.030169f
C46 VGN.n32 VSS 0.02343f
C47 VGN.t1 VSS 1.73884f
C48 VGN.n33 VSS 0.032762f
C49 VGN.n34 VSS 0.02343f
C50 VGN.t5 VSS 1.73884f
C51 VGN.n35 VSS 0.035355f
C52 VGN.t9 VSS 1.82286f
C53 VGN.n36 VSS 0.670152f
C54 VGN.t7 VSS 1.73884f
C55 VGN.n37 VSS 0.657309f
C56 VGN.n38 VSS 0.031008f
C57 VGN.n39 VSS 0.149969f
C58 VGN.n40 VSS 0.02343f
C59 VGN.n41 VSS 0.02343f
C60 VGN.n42 VSS 0.032762f
C61 VGN.n43 VSS 0.032724f
C62 VGN.n44 VSS 0.612956f
C63 VGN.n45 VSS 0.032724f
C64 VGN.n46 VSS 0.02343f
C65 VGN.n47 VSS 0.02343f
C66 VGN.n48 VSS 0.02343f
C67 VGN.n49 VSS 0.035355f
C68 VGN.n50 VSS 0.031008f
C69 VGN.n51 VSS 0.612956f
C70 VGN.n52 VSS 0.03444f
C71 VGN.n53 VSS 0.02343f
C72 VGN.n54 VSS 0.02343f
C73 VGN.n55 VSS 0.02343f
C74 VGN.n56 VSS 0.037948f
C75 VGN.n57 VSS 0.029292f
C76 VGN.n58 VSS 0.664125f
C77 VGN.n59 VSS 0.026412f
C78 VCC.n0 VSS 0.004792f
C79 VCC.n1 VSS 0.006389f
C80 VCC.n2 VSS 0.005143f
C81 VCC.n3 VSS 0.006389f
C82 VCC.n4 VSS 0.006389f
C83 VCC.n5 VSS 0.006389f
C84 VCC.n6 VSS 0.005143f
C85 VCC.n7 VSS 0.006389f
C86 VCC.n8 VSS 0.006389f
C87 VCC.n9 VSS 0.006389f
C88 VCC.n10 VSS 0.006389f
C89 VCC.n11 VSS 0.005143f
C90 VCC.n12 VSS 0.006389f
C91 VCC.n13 VSS 0.006389f
C92 VCC.n14 VSS 0.006389f
C93 VCC.n15 VSS 0.006389f
C94 VCC.n16 VSS 0.005143f
C95 VCC.n17 VSS 0.006389f
C96 VCC.n18 VSS 0.006389f
C97 VCC.n19 VSS 0.006389f
C98 VCC.n20 VSS 0.006389f
C99 VCC.n21 VSS 0.005143f
C100 VCC.n22 VSS 0.006389f
C101 VCC.n23 VSS 0.006389f
C102 VCC.n24 VSS 0.006389f
C103 VCC.n25 VSS 0.006389f
C104 VCC.n26 VSS 0.005143f
C105 VCC.n27 VSS 0.006389f
C106 VCC.n28 VSS 0.006389f
C107 VCC.n29 VSS 0.006389f
C108 VCC.n30 VSS 0.006389f
C109 VCC.n31 VSS 0.005143f
C110 VCC.n32 VSS 0.006389f
C111 VCC.n33 VSS 0.006389f
C112 VCC.n34 VSS 0.006389f
C113 VCC.n35 VSS 0.006389f
C114 VCC.n36 VSS 0.005143f
C115 VCC.n37 VSS 0.006389f
C116 VCC.n38 VSS 0.006389f
C117 VCC.n39 VSS 0.006389f
C118 VCC.n40 VSS 0.006389f
C119 VCC.n41 VSS 0.005143f
C120 VCC.n42 VSS 0.008292f
C121 VCC.n43 VSS 0.006389f
C122 VCC.n44 VSS 0.011976f
C123 VCC.n45 VSS 0.193864f
C124 VCC.n46 VSS 0.365434f
C125 VCC.n47 VSS 0.006389f
C126 VCC.n48 VSS 0.011976f
C127 VCC.n49 VSS 0.005143f
C128 VCC.n50 VSS 0.006389f
C129 VCC.n51 VSS 0.005143f
C130 VCC.n52 VSS 0.006389f
C131 VCC.t8 VSS 0.096932f
C132 VCC.n53 VSS 0.006389f
C133 VCC.n54 VSS 0.005143f
C134 VCC.n55 VSS 0.006389f
C135 VCC.n56 VSS 0.005143f
C136 VCC.n57 VSS 0.006389f
C137 VCC.n58 VSS 0.006389f
C138 VCC.n59 VSS 0.193864f
C139 VCC.n60 VSS 0.006389f
C140 VCC.n61 VSS 0.005143f
C141 VCC.n62 VSS 0.006389f
C142 VCC.n63 VSS 0.005143f
C143 VCC.n64 VSS 0.006389f
C144 VCC.n65 VSS 0.006389f
C145 VCC.n66 VSS 0.193864f
C146 VCC.n67 VSS 0.006389f
C147 VCC.n68 VSS 0.005143f
C148 VCC.n69 VSS 0.006389f
C149 VCC.n70 VSS 0.005143f
C150 VCC.n71 VSS 0.006389f
C151 VCC.n72 VSS 0.006389f
C152 VCC.n73 VSS 0.193864f
C153 VCC.n74 VSS 0.006389f
C154 VCC.n75 VSS 0.005143f
C155 VCC.n76 VSS 0.006389f
C156 VCC.n77 VSS 0.005143f
C157 VCC.n78 VSS 0.006389f
C158 VCC.n79 VSS 0.006389f
C159 VCC.n80 VSS 0.193864f
C160 VCC.n81 VSS 0.006389f
C161 VCC.n82 VSS 0.005143f
C162 VCC.n83 VSS 0.006389f
C163 VCC.n84 VSS 0.005143f
C164 VCC.n85 VSS 0.006389f
C165 VCC.n86 VSS 0.006389f
C166 VCC.n87 VSS 0.193864f
C167 VCC.n88 VSS 0.006389f
C168 VCC.n89 VSS 0.005143f
C169 VCC.n90 VSS 0.006389f
C170 VCC.n91 VSS 0.005143f
C171 VCC.n92 VSS 0.006389f
C172 VCC.n93 VSS 0.006389f
C173 VCC.n94 VSS 0.193864f
C174 VCC.n95 VSS 0.006389f
C175 VCC.n96 VSS 0.005143f
C176 VCC.n97 VSS 0.006389f
C177 VCC.n98 VSS 0.005143f
C178 VCC.n99 VSS 0.006389f
C179 VCC.n100 VSS 0.193864f
C180 VCC.n101 VSS 0.006389f
C181 VCC.n102 VSS 0.005143f
C182 VCC.n103 VSS 0.006389f
C183 VCC.n104 VSS 0.005143f
C184 VCC.n105 VSS 0.006389f
C185 VCC.n106 VSS 0.193864f
C186 VCC.n107 VSS 0.006389f
C187 VCC.n108 VSS 0.006389f
C188 VCC.n109 VSS 0.005143f
C189 VCC.n110 VSS 0.006389f
C190 VCC.n111 VSS 0.005143f
C191 VCC.n112 VSS 0.006389f
C192 VCC.n113 VSS 0.193864f
C193 VCC.n114 VSS 0.006389f
C194 VCC.n115 VSS 0.005143f
C195 VCC.n116 VSS 0.006389f
C196 VCC.n117 VSS 0.005143f
C197 VCC.n118 VSS 0.006389f
C198 VCC.n119 VSS 0.193864f
C199 VCC.n120 VSS 0.006389f
C200 VCC.n121 VSS 0.005143f
C201 VCC.n122 VSS 0.006389f
C202 VCC.n123 VSS 0.005143f
C203 VCC.n124 VSS 0.006389f
C204 VCC.t16 VSS 0.096932f
C205 VCC.n125 VSS 0.006389f
C206 VCC.n126 VSS 0.005143f
C207 VCC.n127 VSS 0.006389f
C208 VCC.n128 VSS 0.005143f
C209 VCC.n129 VSS 0.006389f
C210 VCC.n130 VSS 0.193864f
C211 VCC.n131 VSS 0.149275f
C212 VCC.n132 VSS 0.006389f
C213 VCC.n133 VSS 0.005143f
C214 VCC.n134 VSS 0.006389f
C215 VCC.n135 VSS 0.005143f
C216 VCC.n136 VSS 0.006389f
C217 VCC.n137 VSS 0.193864f
C218 VCC.n138 VSS 0.006389f
C219 VCC.n139 VSS 0.005143f
C220 VCC.n140 VSS 0.006389f
C221 VCC.n141 VSS 0.005143f
C222 VCC.n142 VSS 0.006389f
C223 VCC.n143 VSS 0.193864f
C224 VCC.n144 VSS 0.006389f
C225 VCC.n145 VSS 0.005143f
C226 VCC.n146 VSS 0.006389f
C227 VCC.n147 VSS 0.005143f
C228 VCC.n148 VSS 0.006389f
C229 VCC.t15 VSS 0.096932f
C230 VCC.n149 VSS 0.006389f
C231 VCC.n150 VSS 0.005143f
C232 VCC.n151 VSS 0.006389f
C233 VCC.n152 VSS 0.005143f
C234 VCC.n153 VSS 0.006389f
C235 VCC.n154 VSS 0.193864f
C236 VCC.n155 VSS 0.104687f
C237 VCC.n156 VSS 0.006389f
C238 VCC.n157 VSS 0.005143f
C239 VCC.n158 VSS 0.006389f
C240 VCC.n159 VSS 0.005143f
C241 VCC.n160 VSS 0.006389f
C242 VCC.n161 VSS 0.193864f
C243 VCC.n162 VSS 0.006389f
C244 VCC.n163 VSS 0.005143f
C245 VCC.n164 VSS 0.006389f
C246 VCC.n165 VSS 0.005143f
C247 VCC.n166 VSS 0.006389f
C248 VCC.n167 VSS 0.193864f
C249 VCC.n168 VSS 0.006389f
C250 VCC.n169 VSS 0.005143f
C251 VCC.n170 VSS 0.006389f
C252 VCC.n171 VSS 0.005143f
C253 VCC.n172 VSS 0.006389f
C254 VCC.n173 VSS 0.193864f
C255 VCC.n174 VSS 0.006389f
C256 VCC.n175 VSS 0.005143f
C257 VCC.n176 VSS 0.006389f
C258 VCC.n177 VSS 0.005143f
C259 VCC.n178 VSS 0.006389f
C260 VCC.n179 VSS 0.151214f
C261 VCC.n180 VSS 0.006389f
C262 VCC.n181 VSS 0.005143f
C263 VCC.n182 VSS 0.006389f
C264 VCC.n183 VSS 0.005143f
C265 VCC.n184 VSS 0.006389f
C266 VCC.n185 VSS 0.193864f
C267 VCC.n186 VSS 0.006389f
C268 VCC.n187 VSS 0.005143f
C269 VCC.n188 VSS 0.006389f
C270 VCC.n189 VSS 0.005143f
C271 VCC.n190 VSS 0.006389f
C272 VCC.n191 VSS 0.193864f
C273 VCC.n192 VSS 0.006389f
C274 VCC.n193 VSS 0.005143f
C275 VCC.n194 VSS 0.008292f
C276 VCC.n195 VSS 0.011976f
C277 VCC.n196 VSS 0.365434f
C278 VCC.n197 VSS 0.011976f
C279 VCC.n198 VSS 0.004345f
C280 VCC.n199 VSS 0.004345f
C281 VCC.n200 VSS 0.004345f
C282 VCC.n201 VSS 0.004345f
C283 VCC.n202 VSS 0.004345f
C284 VCC.n203 VSS 0.004345f
C285 VCC.t2 VSS 0.044506f
C286 VCC.t3 VSS 0.058138f
C287 VCC.t0 VSS 0.355333f
C288 VCC.n204 VSS 0.057369f
C289 VCC.n205 VSS 0.039923f
C290 VCC.n206 VSS 0.004345f
C291 VCC.n207 VSS 0.004345f
C292 VCC.n208 VSS 0.004345f
C293 VCC.n209 VSS 0.004345f
C294 VCC.n210 VSS 0.004345f
C295 VCC.n211 VSS 0.004345f
C296 VCC.n212 VSS 0.004345f
C297 VCC.n213 VSS 0.004345f
C298 VCC.t5 VSS 0.044506f
C299 VCC.t6 VSS 0.058138f
C300 VCC.t4 VSS 0.355333f
C301 VCC.n214 VSS 0.057369f
C302 VCC.n215 VSS 0.039923f
C303 VCC.n217 VSS 0.004345f
C304 VCC.n218 VSS 0.004281f
C305 VCC.n219 VSS 0.006055f
C306 VCC.n220 VSS 0.002236f
C307 VCC.n221 VSS 0.004345f
C308 VCC.n222 VSS 0.004345f
C309 VCC.n224 VSS 0.004345f
C310 VCC.n226 VSS 0.004345f
C311 VCC.n227 VSS 0.004345f
C312 VCC.n228 VSS 0.004345f
C313 VCC.n229 VSS 0.004345f
C314 VCC.n230 VSS 0.004345f
C315 VCC.n232 VSS 0.004345f
C316 VCC.n234 VSS 0.004345f
C317 VCC.n235 VSS 0.004345f
C318 VCC.n236 VSS 0.004345f
C319 VCC.n237 VSS 0.004345f
C320 VCC.n238 VSS 0.004345f
C321 VCC.n240 VSS 0.004345f
C322 VCC.n242 VSS 0.004345f
C323 VCC.n243 VSS 0.004345f
C324 VCC.n244 VSS 0.004345f
C325 VCC.n245 VSS 0.004345f
C326 VCC.n246 VSS 0.004345f
C327 VCC.n248 VSS 0.004345f
C328 VCC.n250 VSS 0.004345f
C329 VCC.n251 VSS 0.003131f
C330 VCC.n252 VSS 0.006055f
C331 VCC.n253 VSS 0.003386f
C332 VCC.n254 VSS 0.004345f
C333 VCC.n255 VSS 0.004345f
C334 VCC.n257 VSS 0.004345f
C335 VCC.n259 VSS 0.004345f
C336 VCC.n260 VSS 0.004345f
C337 VCC.n261 VSS 0.004345f
C338 VCC.n262 VSS 0.004345f
C339 VCC.n263 VSS 0.004345f
C340 VCC.n265 VSS 0.004345f
C341 VCC.n267 VSS 0.004345f
C342 VCC.n268 VSS 0.004345f
C343 VCC.n269 VSS 0.004345f
C344 VCC.n270 VSS 0.004345f
C345 VCC.n271 VSS 0.004345f
C346 VCC.n273 VSS 0.004345f
C347 VCC.n275 VSS 0.004345f
C348 VCC.n276 VSS 0.004345f
C349 VCC.n277 VSS 0.008292f
C350 VCC.n278 VSS 0.020972f
C351 VCC.n279 VSS 0.004268f
C352 VCC.n280 VSS 0.012048f
C353 VCC.n281 VSS 0.262686f
C354 VCC.n282 VSS 0.012048f
C355 VCC.n283 VSS 0.004268f
C356 VCC.n284 VSS 0.020972f
C357 VCC.n285 VSS 0.006389f
C358 VCC.n286 VSS 0.006389f
C359 VCC.n287 VSS 0.005143f
C360 VCC.n288 VSS 0.006389f
C361 VCC.n289 VSS 0.193864f
C362 VCC.n290 VSS 0.006389f
C363 VCC.n291 VSS 0.005143f
C364 VCC.n292 VSS 0.006389f
C365 VCC.n293 VSS 0.006389f
C366 VCC.n294 VSS 0.006389f
C367 VCC.n295 VSS 0.005143f
C368 VCC.n296 VSS 0.006389f
C369 VCC.t1 VSS 0.096932f
C370 VCC.n297 VSS 0.139582f
C371 VCC.n298 VSS 0.006389f
C372 VCC.n299 VSS 0.005143f
C373 VCC.n300 VSS 0.006389f
C374 VCC.n301 VSS 0.006389f
C375 VCC.n302 VSS 0.006389f
C376 VCC.n303 VSS 0.005143f
C377 VCC.n304 VSS 0.006389f
C378 VCC.n305 VSS 0.193864f
C379 VCC.n306 VSS 0.006389f
C380 VCC.n307 VSS 0.005143f
C381 VCC.n308 VSS 0.006389f
C382 VCC.n309 VSS 0.006389f
C383 VCC.n310 VSS 0.006389f
C384 VCC.n311 VSS 0.005143f
C385 VCC.n312 VSS 0.006389f
C386 VCC.n313 VSS 0.193864f
C387 VCC.n314 VSS 0.006389f
C388 VCC.n315 VSS 0.005143f
C389 VCC.n316 VSS 0.006389f
C390 VCC.n317 VSS 0.006389f
C391 VCC.n318 VSS 0.006389f
C392 VCC.n319 VSS 0.005143f
C393 VCC.n320 VSS 0.006389f
C394 VCC.n321 VSS 0.193864f
C395 VCC.n322 VSS 0.006389f
C396 VCC.n323 VSS 0.005143f
C397 VCC.n324 VSS 0.006389f
C398 VCC.n325 VSS 0.006389f
C399 VCC.n326 VSS 0.006389f
C400 VCC.n327 VSS 0.005143f
C401 VCC.n328 VSS 0.006389f
C402 VCC.n329 VSS 0.193864f
C403 VCC.n330 VSS 0.006389f
C404 VCC.n331 VSS 0.005143f
C405 VCC.n332 VSS 0.006389f
C406 VCC.n333 VSS 0.006389f
C407 VCC.n334 VSS 0.006389f
C408 VCC.n335 VSS 0.005143f
C409 VCC.n336 VSS 0.006389f
C410 VCC.n337 VSS 0.193864f
C411 VCC.n338 VSS 0.006389f
C412 VCC.n339 VSS 0.005143f
C413 VCC.n340 VSS 0.006389f
C414 VCC.n341 VSS 0.006389f
C415 VCC.n342 VSS 0.006389f
C416 VCC.n343 VSS 0.005143f
C417 VCC.n344 VSS 0.006389f
C418 VCC.n345 VSS 0.186109f
C419 VCC.n346 VSS 0.006389f
C420 VCC.n347 VSS 0.005143f
C421 VCC.n348 VSS 0.006389f
C422 VCC.n349 VSS 0.006389f
C423 VCC.n350 VSS 0.006389f
C424 VCC.n351 VSS 0.005143f
C425 VCC.n352 VSS 0.006389f
C426 VCC.n353 VSS 0.193864f
C427 VCC.n354 VSS 0.006389f
C428 VCC.n355 VSS 0.005143f
C429 VCC.n356 VSS 0.006389f
C430 VCC.n357 VSS 0.006389f
C431 VCC.n358 VSS 0.006389f
C432 VCC.n359 VSS 0.005143f
C433 VCC.n360 VSS 0.006389f
C434 VCC.n361 VSS 0.193864f
C435 VCC.n362 VSS 0.006389f
C436 VCC.n363 VSS 0.005143f
C437 VCC.n364 VSS 0.006389f
C438 VCC.n365 VSS 0.006389f
C439 VCC.n366 VSS 0.006389f
C440 VCC.n367 VSS 0.005143f
C441 VCC.n368 VSS 0.006389f
C442 VCC.n369 VSS 0.193864f
C443 VCC.n370 VSS 0.006389f
C444 VCC.n371 VSS 0.005143f
C445 VCC.n372 VSS 0.006389f
C446 VCC.n373 VSS 0.006389f
C447 VCC.n374 VSS 0.006389f
C448 VCC.n375 VSS 0.005143f
C449 VCC.n376 VSS 0.006389f
C450 VCC.n377 VSS 0.141521f
C451 VCC.n378 VSS 0.006389f
C452 VCC.n379 VSS 0.005143f
C453 VCC.n380 VSS 0.006389f
C454 VCC.n381 VSS 0.006389f
C455 VCC.n382 VSS 0.006389f
C456 VCC.n383 VSS 0.005143f
C457 VCC.n384 VSS 0.006389f
C458 VCC.n385 VSS 0.193864f
C459 VCC.n386 VSS 0.006389f
C460 VCC.n387 VSS 0.005143f
C461 VCC.n388 VSS 0.006389f
C462 VCC.n389 VSS 0.006389f
C463 VCC.n390 VSS 0.006389f
C464 VCC.n391 VSS 0.005143f
C465 VCC.n392 VSS 0.006389f
C466 VCC.n393 VSS 0.193864f
C467 VCC.n394 VSS 0.006389f
C468 VCC.n395 VSS 0.005143f
C469 VCC.n396 VSS 0.006389f
C470 VCC.n397 VSS 0.006389f
C471 VCC.n398 VSS 0.006389f
C472 VCC.n399 VSS 0.005143f
C473 VCC.n400 VSS 0.006389f
C474 VCC.n401 VSS 0.193864f
C475 VCC.n402 VSS 0.006389f
C476 VCC.n403 VSS 0.005143f
C477 VCC.n404 VSS 0.006389f
C478 VCC.n405 VSS 0.006389f
C479 VCC.n406 VSS 0.006389f
C480 VCC.n407 VSS 0.005143f
C481 VCC.n408 VSS 0.006389f
C482 VCC.t14 VSS 0.193864f
C483 VCC.n409 VSS 0.193864f
C484 VCC.n410 VSS 0.193864f
C485 VCC.n411 VSS 0.006389f
C486 VCC.n412 VSS 0.005143f
C487 VCC.n413 VSS 0.006389f
C488 VCC.n414 VSS 0.006389f
C489 VCC.n415 VSS 0.006389f
C490 VCC.n416 VSS 0.005143f
C491 VCC.n417 VSS 0.006389f
C492 VCC.n418 VSS 0.193864f
C493 VCC.n419 VSS 0.193864f
C494 VCC.n420 VSS 0.193864f
C495 VCC.n421 VSS 0.006389f
C496 VCC.n422 VSS 0.005143f
C497 VCC.n423 VSS 0.006389f
C498 VCC.n424 VSS 0.006389f
C499 VCC.n425 VSS 0.006389f
C500 VCC.n426 VSS 0.005143f
C501 VCC.n427 VSS 0.006389f
C502 VCC.n428 VSS 0.141521f
C503 VCC.t17 VSS 0.096932f
C504 VCC.n429 VSS 0.149275f
C505 VCC.n430 VSS 0.193864f
C506 VCC.n431 VSS 0.006389f
C507 VCC.n432 VSS 0.005143f
C508 VCC.n433 VSS 0.006389f
C509 VCC.n434 VSS 0.006389f
C510 VCC.n435 VSS 0.006389f
C511 VCC.n436 VSS 0.005143f
C512 VCC.n437 VSS 0.006389f
C513 VCC.n438 VSS 0.193864f
C514 VCC.n439 VSS 0.193864f
C515 VCC.n440 VSS 0.193864f
C516 VCC.n441 VSS 0.006389f
C517 VCC.n442 VSS 0.005143f
C518 VCC.n443 VSS 0.006389f
C519 VCC.n444 VSS 0.006389f
C520 VCC.n445 VSS 0.006389f
C521 VCC.n446 VSS 0.005143f
C522 VCC.n447 VSS 0.006389f
C523 VCC.n448 VSS 0.186109f
C524 VCC.t18 VSS 0.096932f
C525 VCC.n449 VSS 0.104687f
C526 VCC.n450 VSS 0.193864f
C527 VCC.n451 VSS 0.006389f
C528 VCC.n452 VSS 0.005143f
C529 VCC.n453 VSS 0.006389f
C530 VCC.n454 VSS 0.006389f
C531 VCC.n455 VSS 0.006389f
C532 VCC.n456 VSS 0.005143f
C533 VCC.n457 VSS 0.006389f
C534 VCC.n458 VSS 0.193864f
C535 VCC.n459 VSS 0.193864f
C536 VCC.n460 VSS 0.193864f
C537 VCC.n461 VSS 0.006389f
C538 VCC.n462 VSS 0.005143f
C539 VCC.n463 VSS 0.006389f
C540 VCC.n464 VSS 0.006389f
C541 VCC.n465 VSS 0.006389f
C542 VCC.n466 VSS 0.005143f
C543 VCC.n467 VSS 0.006389f
C544 VCC.n468 VSS 0.193864f
C545 VCC.n469 VSS 0.193864f
C546 VCC.n470 VSS 0.006389f
C547 VCC.n471 VSS 0.151214f
C548 VCC.n472 VSS 0.193864f
C549 VCC.n473 VSS 0.006389f
C550 VCC.n474 VSS 0.005143f
C551 VCC.n475 VSS 0.006389f
C552 VCC.n476 VSS 0.006389f
C553 VCC.n477 VSS 0.006389f
C554 VCC.n478 VSS 0.005143f
C555 VCC.n479 VSS 0.006389f
C556 VCC.n480 VSS 0.139582f
C557 VCC.n481 VSS 0.193864f
C558 VCC.n482 VSS 0.193864f
C559 VCC.n483 VSS 0.006389f
C560 VCC.n484 VSS 0.005143f
C561 VCC.n485 VSS 0.006389f
C562 VCC.n486 VSS 0.006389f
C563 VCC.n487 VSS 0.004345f
C564 VCC.n488 VSS 0.004345f
C565 VCC.n489 VSS 0.004345f
C566 VCC.n490 VSS 0.004345f
C567 VCC.n491 VSS 0.004345f
C568 VCC.n492 VSS 0.004345f
C569 VCC.t10 VSS 0.044506f
C570 VCC.t9 VSS 0.058138f
C571 VCC.t7 VSS 0.355333f
C572 VCC.n493 VSS 0.057369f
C573 VCC.n494 VSS 0.039923f
C574 VCC.n495 VSS 0.004345f
C575 VCC.n496 VSS 0.004345f
C576 VCC.n497 VSS 0.004345f
C577 VCC.n498 VSS 0.004345f
C578 VCC.n499 VSS 0.004345f
C579 VCC.n500 VSS 0.004345f
C580 VCC.n501 VSS 0.004345f
C581 VCC.n502 VSS 0.004345f
C582 VCC.t13 VSS 0.044506f
C583 VCC.t12 VSS 0.058138f
C584 VCC.t11 VSS 0.355333f
C585 VCC.n503 VSS 0.057369f
C586 VCC.n504 VSS 0.039923f
C587 VCC.n506 VSS 0.004345f
C588 VCC.n507 VSS 0.004281f
C589 VCC.n508 VSS 0.006055f
C590 VCC.n509 VSS 0.002236f
C591 VCC.n510 VSS 0.004345f
C592 VCC.n511 VSS 0.004345f
C593 VCC.n513 VSS 0.004345f
C594 VCC.n515 VSS 0.004345f
C595 VCC.n516 VSS 0.004345f
C596 VCC.n517 VSS 0.004345f
C597 VCC.n518 VSS 0.004345f
C598 VCC.n519 VSS 0.004345f
C599 VCC.n521 VSS 0.004345f
C600 VCC.n523 VSS 0.004345f
C601 VCC.n524 VSS 0.004345f
C602 VCC.n525 VSS 0.004345f
C603 VCC.n526 VSS 0.004345f
C604 VCC.n527 VSS 0.004345f
C605 VCC.n529 VSS 0.004345f
C606 VCC.n531 VSS 0.004345f
C607 VCC.n532 VSS 0.004345f
C608 VCC.n533 VSS 0.004345f
C609 VCC.n534 VSS 0.004345f
C610 VCC.n535 VSS 0.004345f
C611 VCC.n537 VSS 0.004345f
C612 VCC.n539 VSS 0.004345f
C613 VCC.n540 VSS 0.003131f
C614 VCC.n541 VSS 0.006055f
C615 VCC.n542 VSS 0.003386f
C616 VCC.n543 VSS 0.004345f
C617 VCC.n544 VSS 0.004345f
C618 VCC.n546 VSS 0.004345f
C619 VCC.n548 VSS 0.004345f
C620 VCC.n549 VSS 0.004345f
C621 VCC.n550 VSS 0.004345f
C622 VCC.n551 VSS 0.004345f
C623 VCC.n552 VSS 0.004345f
C624 VCC.n554 VSS 0.004345f
C625 VCC.n556 VSS 0.004345f
C626 VCC.n557 VSS 0.004345f
C627 VCC.n558 VSS 0.004345f
C628 VCC.n559 VSS 0.004345f
C629 VCC.n560 VSS 0.004345f
C630 VCC.n562 VSS 0.004345f
C631 VCC.n564 VSS 0.004345f
C632 VCC.n565 VSS 0.004345f
C633 VCC.n566 VSS 0.008292f
C634 VCC.n567 VSS 0.020972f
C635 VCC.n568 VSS 0.004268f
C636 VCC.n569 VSS 0.012048f
C637 VCC.n570 VSS 0.262686f
C638 VCC.n571 VSS 0.012048f
C639 VCC.n572 VSS 0.004268f
C640 VCC.n573 VSS 0.020972f
C641 VCC.n574 VSS 0.006389f
C642 VCC.n575 VSS 0.006389f
C643 VCC.n576 VSS 0.005143f
C644 VCC.n577 VSS 0.005143f
C645 VCC.n578 VSS 0.005143f
C646 VCC.n579 VSS 0.006389f
C647 VCC.n580 VSS 0.006389f
C648 VCC.n581 VSS 0.006389f
C649 VCC.n582 VSS 0.005143f
C650 VCC.n583 VSS 0.005143f
C651 VCC.n584 VSS 0.005143f
C652 VCC.n585 VSS 0.006389f
C653 VCC.n586 VSS 0.006389f
C654 VCC.n587 VSS 0.006389f
C655 VCC.n588 VSS 0.005143f
C656 VCC.n589 VSS 0.005143f
C657 VCC.n590 VSS 0.005143f
C658 VCC.n591 VSS 0.006389f
C659 VCC.n592 VSS 0.006389f
C660 VCC.n593 VSS 0.006389f
C661 VCC.n594 VSS 0.005143f
C662 VCC.n595 VSS 0.005143f
C663 VCC.n596 VSS 0.005143f
C664 VCC.n597 VSS 0.006389f
C665 VCC.n598 VSS 0.006389f
C666 VCC.n599 VSS 0.006389f
C667 VCC.n600 VSS 0.005143f
C668 VCC.n601 VSS 0.005143f
C669 VCC.n602 VSS 0.005143f
C670 VCC.n603 VSS 0.006389f
C671 VCC.n604 VSS 0.006389f
C672 VCC.n605 VSS 0.006389f
C673 VCC.n606 VSS 0.005143f
C674 VCC.n607 VSS 0.005143f
C675 VCC.n608 VSS 0.005143f
C676 VCC.n609 VSS 0.006389f
C677 VCC.n610 VSS 0.006389f
C678 VCC.n611 VSS 0.006389f
C679 VCC.n612 VSS 0.005143f
C680 VCC.n613 VSS 0.005143f
C681 VCC.n614 VSS 0.005143f
C682 VCC.n615 VSS 0.006389f
C683 VCC.n616 VSS 0.006389f
C684 VCC.n617 VSS 0.006389f
C685 VCC.n618 VSS 0.005143f
C686 VCC.n619 VSS 0.005143f
C687 VCC.n620 VSS 0.005143f
C688 VCC.n621 VSS 0.005844f
C689 VOUT.n0 VSS 0.047327f
C690 VOUT.t14 VSS 0.730564f
C691 VOUT.n1 VSS 0.047741f
C692 VOUT.n2 VSS 0.02516f
C693 VOUT.n3 VSS 0.046893f
C694 VOUT.n4 VSS 0.02516f
C695 VOUT.t18 VSS 0.730564f
C696 VOUT.n5 VSS 0.046893f
C697 VOUT.n6 VSS 0.02516f
C698 VOUT.n7 VSS 0.046893f
C699 VOUT.n8 VSS 0.02516f
C700 VOUT.t32 VSS 0.730564f
C701 VOUT.n9 VSS 0.046893f
C702 VOUT.n10 VSS 0.02516f
C703 VOUT.n11 VSS 0.046893f
C704 VOUT.n12 VSS 0.330792f
C705 VOUT.t20 VSS 0.730564f
C706 VOUT.t24 VSS 1.04602f
C707 VOUT.n13 VSS 0.416119f
C708 VOUT.n14 VSS 0.387538f
C709 VOUT.n15 VSS 0.034391f
C710 VOUT.n16 VSS 0.046893f
C711 VOUT.n17 VSS 0.02516f
C712 VOUT.n18 VSS 0.02516f
C713 VOUT.n19 VSS 0.02516f
C714 VOUT.n20 VSS 0.04543f
C715 VOUT.n21 VSS 0.024966f
C716 VOUT.n22 VSS 0.04996f
C717 VOUT.n23 VSS 0.02516f
C718 VOUT.n24 VSS 0.02516f
C719 VOUT.n25 VSS 0.02516f
C720 VOUT.n26 VSS 0.046893f
C721 VOUT.n27 VSS 0.320969f
C722 VOUT.n28 VSS 0.046893f
C723 VOUT.n29 VSS 0.02516f
C724 VOUT.n30 VSS 0.02516f
C725 VOUT.n31 VSS 0.02516f
C726 VOUT.n32 VSS 0.04996f
C727 VOUT.n33 VSS 0.024966f
C728 VOUT.n34 VSS 0.04543f
C729 VOUT.n35 VSS 0.02516f
C730 VOUT.n36 VSS 0.02516f
C731 VOUT.n37 VSS 0.02516f
C732 VOUT.n38 VSS 0.046893f
C733 VOUT.n39 VSS 0.034391f
C734 VOUT.n40 VSS 0.297227f
C735 VOUT.n41 VSS 0.036243f
C736 VOUT.n42 VSS 0.02516f
C737 VOUT.n43 VSS 0.02516f
C738 VOUT.n44 VSS 0.02516f
C739 VOUT.n45 VSS 0.046893f
C740 VOUT.n46 VSS 0.043265f
C741 VOUT.n47 VSS 0.02935f
C742 VOUT.n48 VSS 0.02516f
C743 VOUT.n49 VSS 0.02516f
C744 VOUT.n50 VSS 0.02516f
C745 VOUT.n51 VSS 0.046893f
C746 VOUT.n52 VSS 0.04504f
C747 VOUT.n53 VSS 0.410158f
C748 VOUT.n54 VSS 0.177199f
C749 VOUT.n55 VSS 0.571454f
C750 VOUT.n56 VSS 0.201193f
C751 VOUT.t1 VSS 1.62653f
C752 VOUT.t7 VSS 0.257196f
C753 VOUT.n57 VSS 0.119112f
C754 VOUT.n58 VSS 0.11496f
C755 VOUT.t33 VSS 0.046382f
C756 VOUT.t15 VSS 0.20198f
C757 VOUT.t19 VSS 0.046382f
C758 VOUT.n59 VSS 0.121029f
C759 VOUT.n60 VSS 0.604649f
C760 VOUT.n61 VSS 0.604649f
C761 VOUT.t13 VSS 0.046382f
C762 VOUT.n62 VSS 0.047327f
C763 VOUT.t16 VSS 0.730564f
C764 VOUT.n63 VSS 0.047741f
C765 VOUT.n64 VSS 0.02516f
C766 VOUT.n65 VSS 0.046893f
C767 VOUT.n66 VSS 0.02516f
C768 VOUT.t22 VSS 0.730564f
C769 VOUT.n67 VSS 0.046893f
C770 VOUT.n68 VSS 0.02516f
C771 VOUT.n69 VSS 0.046893f
C772 VOUT.n70 VSS 0.02516f
C773 VOUT.t12 VSS 0.730564f
C774 VOUT.n71 VSS 0.046893f
C775 VOUT.n72 VSS 0.02516f
C776 VOUT.n73 VSS 0.046893f
C777 VOUT.n74 VSS 0.330791f
C778 VOUT.t27 VSS 0.730564f
C779 VOUT.t29 VSS 1.04602f
C780 VOUT.n75 VSS 0.416118f
C781 VOUT.n76 VSS 0.387538f
C782 VOUT.n77 VSS 0.034391f
C783 VOUT.n78 VSS 0.046893f
C784 VOUT.n79 VSS 0.02516f
C785 VOUT.n80 VSS 0.02516f
C786 VOUT.n81 VSS 0.02516f
C787 VOUT.n82 VSS 0.04543f
C788 VOUT.n83 VSS 0.024966f
C789 VOUT.n84 VSS 0.04996f
C790 VOUT.n85 VSS 0.02516f
C791 VOUT.n86 VSS 0.02516f
C792 VOUT.n87 VSS 0.02516f
C793 VOUT.n88 VSS 0.046893f
C794 VOUT.n89 VSS 0.320969f
C795 VOUT.n90 VSS 0.046893f
C796 VOUT.n91 VSS 0.02516f
C797 VOUT.n92 VSS 0.02516f
C798 VOUT.n93 VSS 0.02516f
C799 VOUT.n94 VSS 0.04996f
C800 VOUT.n95 VSS 0.024966f
C801 VOUT.n96 VSS 0.04543f
C802 VOUT.n97 VSS 0.02516f
C803 VOUT.n98 VSS 0.02516f
C804 VOUT.n99 VSS 0.02516f
C805 VOUT.n100 VSS 0.046893f
C806 VOUT.n101 VSS 0.034391f
C807 VOUT.n102 VSS 0.297227f
C808 VOUT.n103 VSS 0.036243f
C809 VOUT.n104 VSS 0.02516f
C810 VOUT.n105 VSS 0.02516f
C811 VOUT.n106 VSS 0.02516f
C812 VOUT.n107 VSS 0.046893f
C813 VOUT.n108 VSS 0.043265f
C814 VOUT.n109 VSS 0.02935f
C815 VOUT.n110 VSS 0.02516f
C816 VOUT.n111 VSS 0.02516f
C817 VOUT.n112 VSS 0.02516f
C818 VOUT.n113 VSS 0.046893f
C819 VOUT.n114 VSS 0.04504f
C820 VOUT.n115 VSS 0.410158f
C821 VOUT.n116 VSS 0.084343f
C822 VOUT.n117 VSS 0.17772f
C823 VOUT.t17 VSS 0.20198f
C824 VOUT.n118 VSS 0.121029f
C825 VOUT.t23 VSS 0.046382f
C826 VOUT.n119 VSS 0.104762f
C827 VOUT.n120 VSS 0.366603f
C828 VOUT.t31 VSS 0.156495f
C829 VOUT.n121 VSS 0.290859f
C830 VOUT.n122 VSS 0.358194f
C831 VOUT.n123 VSS 0.104762f
C832 VOUT.t28 VSS 0.046382f
C833 VOUT.t30 VSS 0.023191f
C834 VOUT.n124 VSS 0.121029f
C835 VOUT.n125 VSS 0.301421f
C836 VOUT.n126 VSS 0.174641f
C837 VOUT.n127 VSS 0.478304f
C838 VOUT.t25 VSS 0.023191f
C839 VOUT.n128 VSS 0.121029f
C840 VOUT.t21 VSS 0.046382f
C841 VOUT.n129 VSS 0.104762f
C842 VOUT.n130 VSS 0.710144f
C843 VOUT.t26 VSS 0.156495f
C844 VOUT.n131 VSS 0.290099f
C845 VOUT.n132 VSS 0.531263f
C846 VOUT.n133 VSS 0.345517f
C847 VOUT.t3 VSS 0.257196f
C848 VOUT.t8 VSS 1.62653f
C849 VOUT.n134 VSS 1.16875f
C850 VOUT.t4 VSS 0.257196f
C851 VOUT.n135 VSS 1.1481f
C852 VOUT.t6 VSS 1.45774f
C853 VOUT.n136 VSS 0.487727f
C854 VOUT.t11 VSS 1.45774f
C855 VOUT.n137 VSS 0.487727f
C856 VOUT.n138 VSS 0.399188f
C857 VOUT.n139 VSS 1.14095f
C858 VOUT.t0 VSS 0.257196f
C859 VOUT.t10 VSS 0.128598f
C860 VOUT.n140 VSS 1.16875f
C861 VOUT.n141 VSS 0.49422f
C862 VOUT.n142 VSS 0.674999f
C863 VOUT.n143 VSS 1.14095f
C864 VOUT.t9 VSS 0.257196f
C865 VOUT.t5 VSS 0.128598f
C866 VOUT.n144 VSS 1.16875f
C867 VOUT.n145 VSS 0.188588f
C868 VOUT.n146 VSS 0.345517f
C869 VOUT.n147 VSS 1.16875f
C870 VOUT.t2 VSS 0.257196f
C871 VOUT.n148 VSS 1.14095f
C872 VOUT.n149 VSS 0.17461f
.ends

