* NGSPICE file created from diff_pair_sample_1105.ext - technology: sky130A

.subckt diff_pair_sample_1105 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.65155 pd=16.4 as=6.2673 ps=32.92 w=16.07 l=3.6
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=0 ps=0 w=16.07 l=3.6
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=0 ps=0 w=16.07 l=3.6
X3 VTAIL.t4 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=2.65155 ps=16.4 w=16.07 l=3.6
X4 VDD1.t1 VP.t2 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.65155 pd=16.4 as=6.2673 ps=32.92 w=16.07 l=3.6
X5 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=0 ps=0 w=16.07 l=3.6
X6 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.65155 pd=16.4 as=6.2673 ps=32.92 w=16.07 l=3.6
X7 VDD2.t2 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.65155 pd=16.4 as=6.2673 ps=32.92 w=16.07 l=3.6
X8 VTAIL.t1 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=2.65155 ps=16.4 w=16.07 l=3.6
X9 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=2.65155 ps=16.4 w=16.07 l=3.6
X10 VTAIL.t7 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=2.65155 ps=16.4 w=16.07 l=3.6
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.2673 pd=32.92 as=0 ps=0 w=16.07 l=3.6
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n5 VP.t3 142.452
R9 VP.n5 VP.t0 141.208
R10 VP.n6 VP.t1 107.581
R11 VP.n0 VP.t2 107.581
R12 VP.n7 VP.n6 79.5466
R13 VP.n20 VP.n0 79.5466
R14 VP.n12 VP.n2 56.5193
R15 VP.n7 VP.n5 54.6571
R16 VP.n10 VP.n4 24.4675
R17 VP.n11 VP.n10 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n16 VP.n2 24.4675
R20 VP.n17 VP.n16 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n6 VP.n4 10.5213
R23 VP.n18 VP.n0 10.5213
R24 VP.n8 VP.n7 0.354971
R25 VP.n20 VP.n19 0.354971
R26 VP VP.n20 0.26696
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VTAIL.n714 VTAIL.n630 289.615
R35 VTAIL.n84 VTAIL.n0 289.615
R36 VTAIL.n174 VTAIL.n90 289.615
R37 VTAIL.n264 VTAIL.n180 289.615
R38 VTAIL.n624 VTAIL.n540 289.615
R39 VTAIL.n534 VTAIL.n450 289.615
R40 VTAIL.n444 VTAIL.n360 289.615
R41 VTAIL.n354 VTAIL.n270 289.615
R42 VTAIL.n658 VTAIL.n657 185
R43 VTAIL.n663 VTAIL.n662 185
R44 VTAIL.n665 VTAIL.n664 185
R45 VTAIL.n654 VTAIL.n653 185
R46 VTAIL.n671 VTAIL.n670 185
R47 VTAIL.n673 VTAIL.n672 185
R48 VTAIL.n650 VTAIL.n649 185
R49 VTAIL.n679 VTAIL.n678 185
R50 VTAIL.n681 VTAIL.n680 185
R51 VTAIL.n646 VTAIL.n645 185
R52 VTAIL.n687 VTAIL.n686 185
R53 VTAIL.n689 VTAIL.n688 185
R54 VTAIL.n642 VTAIL.n641 185
R55 VTAIL.n695 VTAIL.n694 185
R56 VTAIL.n697 VTAIL.n696 185
R57 VTAIL.n638 VTAIL.n637 185
R58 VTAIL.n704 VTAIL.n703 185
R59 VTAIL.n705 VTAIL.n636 185
R60 VTAIL.n707 VTAIL.n706 185
R61 VTAIL.n634 VTAIL.n633 185
R62 VTAIL.n713 VTAIL.n712 185
R63 VTAIL.n715 VTAIL.n714 185
R64 VTAIL.n28 VTAIL.n27 185
R65 VTAIL.n33 VTAIL.n32 185
R66 VTAIL.n35 VTAIL.n34 185
R67 VTAIL.n24 VTAIL.n23 185
R68 VTAIL.n41 VTAIL.n40 185
R69 VTAIL.n43 VTAIL.n42 185
R70 VTAIL.n20 VTAIL.n19 185
R71 VTAIL.n49 VTAIL.n48 185
R72 VTAIL.n51 VTAIL.n50 185
R73 VTAIL.n16 VTAIL.n15 185
R74 VTAIL.n57 VTAIL.n56 185
R75 VTAIL.n59 VTAIL.n58 185
R76 VTAIL.n12 VTAIL.n11 185
R77 VTAIL.n65 VTAIL.n64 185
R78 VTAIL.n67 VTAIL.n66 185
R79 VTAIL.n8 VTAIL.n7 185
R80 VTAIL.n74 VTAIL.n73 185
R81 VTAIL.n75 VTAIL.n6 185
R82 VTAIL.n77 VTAIL.n76 185
R83 VTAIL.n4 VTAIL.n3 185
R84 VTAIL.n83 VTAIL.n82 185
R85 VTAIL.n85 VTAIL.n84 185
R86 VTAIL.n118 VTAIL.n117 185
R87 VTAIL.n123 VTAIL.n122 185
R88 VTAIL.n125 VTAIL.n124 185
R89 VTAIL.n114 VTAIL.n113 185
R90 VTAIL.n131 VTAIL.n130 185
R91 VTAIL.n133 VTAIL.n132 185
R92 VTAIL.n110 VTAIL.n109 185
R93 VTAIL.n139 VTAIL.n138 185
R94 VTAIL.n141 VTAIL.n140 185
R95 VTAIL.n106 VTAIL.n105 185
R96 VTAIL.n147 VTAIL.n146 185
R97 VTAIL.n149 VTAIL.n148 185
R98 VTAIL.n102 VTAIL.n101 185
R99 VTAIL.n155 VTAIL.n154 185
R100 VTAIL.n157 VTAIL.n156 185
R101 VTAIL.n98 VTAIL.n97 185
R102 VTAIL.n164 VTAIL.n163 185
R103 VTAIL.n165 VTAIL.n96 185
R104 VTAIL.n167 VTAIL.n166 185
R105 VTAIL.n94 VTAIL.n93 185
R106 VTAIL.n173 VTAIL.n172 185
R107 VTAIL.n175 VTAIL.n174 185
R108 VTAIL.n208 VTAIL.n207 185
R109 VTAIL.n213 VTAIL.n212 185
R110 VTAIL.n215 VTAIL.n214 185
R111 VTAIL.n204 VTAIL.n203 185
R112 VTAIL.n221 VTAIL.n220 185
R113 VTAIL.n223 VTAIL.n222 185
R114 VTAIL.n200 VTAIL.n199 185
R115 VTAIL.n229 VTAIL.n228 185
R116 VTAIL.n231 VTAIL.n230 185
R117 VTAIL.n196 VTAIL.n195 185
R118 VTAIL.n237 VTAIL.n236 185
R119 VTAIL.n239 VTAIL.n238 185
R120 VTAIL.n192 VTAIL.n191 185
R121 VTAIL.n245 VTAIL.n244 185
R122 VTAIL.n247 VTAIL.n246 185
R123 VTAIL.n188 VTAIL.n187 185
R124 VTAIL.n254 VTAIL.n253 185
R125 VTAIL.n255 VTAIL.n186 185
R126 VTAIL.n257 VTAIL.n256 185
R127 VTAIL.n184 VTAIL.n183 185
R128 VTAIL.n263 VTAIL.n262 185
R129 VTAIL.n265 VTAIL.n264 185
R130 VTAIL.n625 VTAIL.n624 185
R131 VTAIL.n623 VTAIL.n622 185
R132 VTAIL.n544 VTAIL.n543 185
R133 VTAIL.n617 VTAIL.n616 185
R134 VTAIL.n615 VTAIL.n546 185
R135 VTAIL.n614 VTAIL.n613 185
R136 VTAIL.n549 VTAIL.n547 185
R137 VTAIL.n608 VTAIL.n607 185
R138 VTAIL.n606 VTAIL.n605 185
R139 VTAIL.n553 VTAIL.n552 185
R140 VTAIL.n600 VTAIL.n599 185
R141 VTAIL.n598 VTAIL.n597 185
R142 VTAIL.n557 VTAIL.n556 185
R143 VTAIL.n592 VTAIL.n591 185
R144 VTAIL.n590 VTAIL.n589 185
R145 VTAIL.n561 VTAIL.n560 185
R146 VTAIL.n584 VTAIL.n583 185
R147 VTAIL.n582 VTAIL.n581 185
R148 VTAIL.n565 VTAIL.n564 185
R149 VTAIL.n576 VTAIL.n575 185
R150 VTAIL.n574 VTAIL.n573 185
R151 VTAIL.n569 VTAIL.n568 185
R152 VTAIL.n535 VTAIL.n534 185
R153 VTAIL.n533 VTAIL.n532 185
R154 VTAIL.n454 VTAIL.n453 185
R155 VTAIL.n527 VTAIL.n526 185
R156 VTAIL.n525 VTAIL.n456 185
R157 VTAIL.n524 VTAIL.n523 185
R158 VTAIL.n459 VTAIL.n457 185
R159 VTAIL.n518 VTAIL.n517 185
R160 VTAIL.n516 VTAIL.n515 185
R161 VTAIL.n463 VTAIL.n462 185
R162 VTAIL.n510 VTAIL.n509 185
R163 VTAIL.n508 VTAIL.n507 185
R164 VTAIL.n467 VTAIL.n466 185
R165 VTAIL.n502 VTAIL.n501 185
R166 VTAIL.n500 VTAIL.n499 185
R167 VTAIL.n471 VTAIL.n470 185
R168 VTAIL.n494 VTAIL.n493 185
R169 VTAIL.n492 VTAIL.n491 185
R170 VTAIL.n475 VTAIL.n474 185
R171 VTAIL.n486 VTAIL.n485 185
R172 VTAIL.n484 VTAIL.n483 185
R173 VTAIL.n479 VTAIL.n478 185
R174 VTAIL.n445 VTAIL.n444 185
R175 VTAIL.n443 VTAIL.n442 185
R176 VTAIL.n364 VTAIL.n363 185
R177 VTAIL.n437 VTAIL.n436 185
R178 VTAIL.n435 VTAIL.n366 185
R179 VTAIL.n434 VTAIL.n433 185
R180 VTAIL.n369 VTAIL.n367 185
R181 VTAIL.n428 VTAIL.n427 185
R182 VTAIL.n426 VTAIL.n425 185
R183 VTAIL.n373 VTAIL.n372 185
R184 VTAIL.n420 VTAIL.n419 185
R185 VTAIL.n418 VTAIL.n417 185
R186 VTAIL.n377 VTAIL.n376 185
R187 VTAIL.n412 VTAIL.n411 185
R188 VTAIL.n410 VTAIL.n409 185
R189 VTAIL.n381 VTAIL.n380 185
R190 VTAIL.n404 VTAIL.n403 185
R191 VTAIL.n402 VTAIL.n401 185
R192 VTAIL.n385 VTAIL.n384 185
R193 VTAIL.n396 VTAIL.n395 185
R194 VTAIL.n394 VTAIL.n393 185
R195 VTAIL.n389 VTAIL.n388 185
R196 VTAIL.n355 VTAIL.n354 185
R197 VTAIL.n353 VTAIL.n352 185
R198 VTAIL.n274 VTAIL.n273 185
R199 VTAIL.n347 VTAIL.n346 185
R200 VTAIL.n345 VTAIL.n276 185
R201 VTAIL.n344 VTAIL.n343 185
R202 VTAIL.n279 VTAIL.n277 185
R203 VTAIL.n338 VTAIL.n337 185
R204 VTAIL.n336 VTAIL.n335 185
R205 VTAIL.n283 VTAIL.n282 185
R206 VTAIL.n330 VTAIL.n329 185
R207 VTAIL.n328 VTAIL.n327 185
R208 VTAIL.n287 VTAIL.n286 185
R209 VTAIL.n322 VTAIL.n321 185
R210 VTAIL.n320 VTAIL.n319 185
R211 VTAIL.n291 VTAIL.n290 185
R212 VTAIL.n314 VTAIL.n313 185
R213 VTAIL.n312 VTAIL.n311 185
R214 VTAIL.n295 VTAIL.n294 185
R215 VTAIL.n306 VTAIL.n305 185
R216 VTAIL.n304 VTAIL.n303 185
R217 VTAIL.n299 VTAIL.n298 185
R218 VTAIL.n659 VTAIL.t3 147.659
R219 VTAIL.n29 VTAIL.t1 147.659
R220 VTAIL.n119 VTAIL.t6 147.659
R221 VTAIL.n209 VTAIL.t4 147.659
R222 VTAIL.n570 VTAIL.t5 147.659
R223 VTAIL.n480 VTAIL.t7 147.659
R224 VTAIL.n390 VTAIL.t0 147.659
R225 VTAIL.n300 VTAIL.t2 147.659
R226 VTAIL.n663 VTAIL.n657 104.615
R227 VTAIL.n664 VTAIL.n663 104.615
R228 VTAIL.n664 VTAIL.n653 104.615
R229 VTAIL.n671 VTAIL.n653 104.615
R230 VTAIL.n672 VTAIL.n671 104.615
R231 VTAIL.n672 VTAIL.n649 104.615
R232 VTAIL.n679 VTAIL.n649 104.615
R233 VTAIL.n680 VTAIL.n679 104.615
R234 VTAIL.n680 VTAIL.n645 104.615
R235 VTAIL.n687 VTAIL.n645 104.615
R236 VTAIL.n688 VTAIL.n687 104.615
R237 VTAIL.n688 VTAIL.n641 104.615
R238 VTAIL.n695 VTAIL.n641 104.615
R239 VTAIL.n696 VTAIL.n695 104.615
R240 VTAIL.n696 VTAIL.n637 104.615
R241 VTAIL.n704 VTAIL.n637 104.615
R242 VTAIL.n705 VTAIL.n704 104.615
R243 VTAIL.n706 VTAIL.n705 104.615
R244 VTAIL.n706 VTAIL.n633 104.615
R245 VTAIL.n713 VTAIL.n633 104.615
R246 VTAIL.n714 VTAIL.n713 104.615
R247 VTAIL.n33 VTAIL.n27 104.615
R248 VTAIL.n34 VTAIL.n33 104.615
R249 VTAIL.n34 VTAIL.n23 104.615
R250 VTAIL.n41 VTAIL.n23 104.615
R251 VTAIL.n42 VTAIL.n41 104.615
R252 VTAIL.n42 VTAIL.n19 104.615
R253 VTAIL.n49 VTAIL.n19 104.615
R254 VTAIL.n50 VTAIL.n49 104.615
R255 VTAIL.n50 VTAIL.n15 104.615
R256 VTAIL.n57 VTAIL.n15 104.615
R257 VTAIL.n58 VTAIL.n57 104.615
R258 VTAIL.n58 VTAIL.n11 104.615
R259 VTAIL.n65 VTAIL.n11 104.615
R260 VTAIL.n66 VTAIL.n65 104.615
R261 VTAIL.n66 VTAIL.n7 104.615
R262 VTAIL.n74 VTAIL.n7 104.615
R263 VTAIL.n75 VTAIL.n74 104.615
R264 VTAIL.n76 VTAIL.n75 104.615
R265 VTAIL.n76 VTAIL.n3 104.615
R266 VTAIL.n83 VTAIL.n3 104.615
R267 VTAIL.n84 VTAIL.n83 104.615
R268 VTAIL.n123 VTAIL.n117 104.615
R269 VTAIL.n124 VTAIL.n123 104.615
R270 VTAIL.n124 VTAIL.n113 104.615
R271 VTAIL.n131 VTAIL.n113 104.615
R272 VTAIL.n132 VTAIL.n131 104.615
R273 VTAIL.n132 VTAIL.n109 104.615
R274 VTAIL.n139 VTAIL.n109 104.615
R275 VTAIL.n140 VTAIL.n139 104.615
R276 VTAIL.n140 VTAIL.n105 104.615
R277 VTAIL.n147 VTAIL.n105 104.615
R278 VTAIL.n148 VTAIL.n147 104.615
R279 VTAIL.n148 VTAIL.n101 104.615
R280 VTAIL.n155 VTAIL.n101 104.615
R281 VTAIL.n156 VTAIL.n155 104.615
R282 VTAIL.n156 VTAIL.n97 104.615
R283 VTAIL.n164 VTAIL.n97 104.615
R284 VTAIL.n165 VTAIL.n164 104.615
R285 VTAIL.n166 VTAIL.n165 104.615
R286 VTAIL.n166 VTAIL.n93 104.615
R287 VTAIL.n173 VTAIL.n93 104.615
R288 VTAIL.n174 VTAIL.n173 104.615
R289 VTAIL.n213 VTAIL.n207 104.615
R290 VTAIL.n214 VTAIL.n213 104.615
R291 VTAIL.n214 VTAIL.n203 104.615
R292 VTAIL.n221 VTAIL.n203 104.615
R293 VTAIL.n222 VTAIL.n221 104.615
R294 VTAIL.n222 VTAIL.n199 104.615
R295 VTAIL.n229 VTAIL.n199 104.615
R296 VTAIL.n230 VTAIL.n229 104.615
R297 VTAIL.n230 VTAIL.n195 104.615
R298 VTAIL.n237 VTAIL.n195 104.615
R299 VTAIL.n238 VTAIL.n237 104.615
R300 VTAIL.n238 VTAIL.n191 104.615
R301 VTAIL.n245 VTAIL.n191 104.615
R302 VTAIL.n246 VTAIL.n245 104.615
R303 VTAIL.n246 VTAIL.n187 104.615
R304 VTAIL.n254 VTAIL.n187 104.615
R305 VTAIL.n255 VTAIL.n254 104.615
R306 VTAIL.n256 VTAIL.n255 104.615
R307 VTAIL.n256 VTAIL.n183 104.615
R308 VTAIL.n263 VTAIL.n183 104.615
R309 VTAIL.n264 VTAIL.n263 104.615
R310 VTAIL.n624 VTAIL.n623 104.615
R311 VTAIL.n623 VTAIL.n543 104.615
R312 VTAIL.n616 VTAIL.n543 104.615
R313 VTAIL.n616 VTAIL.n615 104.615
R314 VTAIL.n615 VTAIL.n614 104.615
R315 VTAIL.n614 VTAIL.n547 104.615
R316 VTAIL.n607 VTAIL.n547 104.615
R317 VTAIL.n607 VTAIL.n606 104.615
R318 VTAIL.n606 VTAIL.n552 104.615
R319 VTAIL.n599 VTAIL.n552 104.615
R320 VTAIL.n599 VTAIL.n598 104.615
R321 VTAIL.n598 VTAIL.n556 104.615
R322 VTAIL.n591 VTAIL.n556 104.615
R323 VTAIL.n591 VTAIL.n590 104.615
R324 VTAIL.n590 VTAIL.n560 104.615
R325 VTAIL.n583 VTAIL.n560 104.615
R326 VTAIL.n583 VTAIL.n582 104.615
R327 VTAIL.n582 VTAIL.n564 104.615
R328 VTAIL.n575 VTAIL.n564 104.615
R329 VTAIL.n575 VTAIL.n574 104.615
R330 VTAIL.n574 VTAIL.n568 104.615
R331 VTAIL.n534 VTAIL.n533 104.615
R332 VTAIL.n533 VTAIL.n453 104.615
R333 VTAIL.n526 VTAIL.n453 104.615
R334 VTAIL.n526 VTAIL.n525 104.615
R335 VTAIL.n525 VTAIL.n524 104.615
R336 VTAIL.n524 VTAIL.n457 104.615
R337 VTAIL.n517 VTAIL.n457 104.615
R338 VTAIL.n517 VTAIL.n516 104.615
R339 VTAIL.n516 VTAIL.n462 104.615
R340 VTAIL.n509 VTAIL.n462 104.615
R341 VTAIL.n509 VTAIL.n508 104.615
R342 VTAIL.n508 VTAIL.n466 104.615
R343 VTAIL.n501 VTAIL.n466 104.615
R344 VTAIL.n501 VTAIL.n500 104.615
R345 VTAIL.n500 VTAIL.n470 104.615
R346 VTAIL.n493 VTAIL.n470 104.615
R347 VTAIL.n493 VTAIL.n492 104.615
R348 VTAIL.n492 VTAIL.n474 104.615
R349 VTAIL.n485 VTAIL.n474 104.615
R350 VTAIL.n485 VTAIL.n484 104.615
R351 VTAIL.n484 VTAIL.n478 104.615
R352 VTAIL.n444 VTAIL.n443 104.615
R353 VTAIL.n443 VTAIL.n363 104.615
R354 VTAIL.n436 VTAIL.n363 104.615
R355 VTAIL.n436 VTAIL.n435 104.615
R356 VTAIL.n435 VTAIL.n434 104.615
R357 VTAIL.n434 VTAIL.n367 104.615
R358 VTAIL.n427 VTAIL.n367 104.615
R359 VTAIL.n427 VTAIL.n426 104.615
R360 VTAIL.n426 VTAIL.n372 104.615
R361 VTAIL.n419 VTAIL.n372 104.615
R362 VTAIL.n419 VTAIL.n418 104.615
R363 VTAIL.n418 VTAIL.n376 104.615
R364 VTAIL.n411 VTAIL.n376 104.615
R365 VTAIL.n411 VTAIL.n410 104.615
R366 VTAIL.n410 VTAIL.n380 104.615
R367 VTAIL.n403 VTAIL.n380 104.615
R368 VTAIL.n403 VTAIL.n402 104.615
R369 VTAIL.n402 VTAIL.n384 104.615
R370 VTAIL.n395 VTAIL.n384 104.615
R371 VTAIL.n395 VTAIL.n394 104.615
R372 VTAIL.n394 VTAIL.n388 104.615
R373 VTAIL.n354 VTAIL.n353 104.615
R374 VTAIL.n353 VTAIL.n273 104.615
R375 VTAIL.n346 VTAIL.n273 104.615
R376 VTAIL.n346 VTAIL.n345 104.615
R377 VTAIL.n345 VTAIL.n344 104.615
R378 VTAIL.n344 VTAIL.n277 104.615
R379 VTAIL.n337 VTAIL.n277 104.615
R380 VTAIL.n337 VTAIL.n336 104.615
R381 VTAIL.n336 VTAIL.n282 104.615
R382 VTAIL.n329 VTAIL.n282 104.615
R383 VTAIL.n329 VTAIL.n328 104.615
R384 VTAIL.n328 VTAIL.n286 104.615
R385 VTAIL.n321 VTAIL.n286 104.615
R386 VTAIL.n321 VTAIL.n320 104.615
R387 VTAIL.n320 VTAIL.n290 104.615
R388 VTAIL.n313 VTAIL.n290 104.615
R389 VTAIL.n313 VTAIL.n312 104.615
R390 VTAIL.n312 VTAIL.n294 104.615
R391 VTAIL.n305 VTAIL.n294 104.615
R392 VTAIL.n305 VTAIL.n304 104.615
R393 VTAIL.n304 VTAIL.n298 104.615
R394 VTAIL.t3 VTAIL.n657 52.3082
R395 VTAIL.t1 VTAIL.n27 52.3082
R396 VTAIL.t6 VTAIL.n117 52.3082
R397 VTAIL.t4 VTAIL.n207 52.3082
R398 VTAIL.t5 VTAIL.n568 52.3082
R399 VTAIL.t7 VTAIL.n478 52.3082
R400 VTAIL.t0 VTAIL.n388 52.3082
R401 VTAIL.t2 VTAIL.n298 52.3082
R402 VTAIL.n719 VTAIL.n718 31.9914
R403 VTAIL.n89 VTAIL.n88 31.9914
R404 VTAIL.n179 VTAIL.n178 31.9914
R405 VTAIL.n269 VTAIL.n268 31.9914
R406 VTAIL.n629 VTAIL.n628 31.9914
R407 VTAIL.n539 VTAIL.n538 31.9914
R408 VTAIL.n449 VTAIL.n448 31.9914
R409 VTAIL.n359 VTAIL.n358 31.9914
R410 VTAIL.n719 VTAIL.n629 29.6083
R411 VTAIL.n359 VTAIL.n269 29.6083
R412 VTAIL.n659 VTAIL.n658 15.6677
R413 VTAIL.n29 VTAIL.n28 15.6677
R414 VTAIL.n119 VTAIL.n118 15.6677
R415 VTAIL.n209 VTAIL.n208 15.6677
R416 VTAIL.n570 VTAIL.n569 15.6677
R417 VTAIL.n480 VTAIL.n479 15.6677
R418 VTAIL.n390 VTAIL.n389 15.6677
R419 VTAIL.n300 VTAIL.n299 15.6677
R420 VTAIL.n707 VTAIL.n636 13.1884
R421 VTAIL.n77 VTAIL.n6 13.1884
R422 VTAIL.n167 VTAIL.n96 13.1884
R423 VTAIL.n257 VTAIL.n186 13.1884
R424 VTAIL.n617 VTAIL.n546 13.1884
R425 VTAIL.n527 VTAIL.n456 13.1884
R426 VTAIL.n437 VTAIL.n366 13.1884
R427 VTAIL.n347 VTAIL.n276 13.1884
R428 VTAIL.n662 VTAIL.n661 12.8005
R429 VTAIL.n703 VTAIL.n702 12.8005
R430 VTAIL.n708 VTAIL.n634 12.8005
R431 VTAIL.n32 VTAIL.n31 12.8005
R432 VTAIL.n73 VTAIL.n72 12.8005
R433 VTAIL.n78 VTAIL.n4 12.8005
R434 VTAIL.n122 VTAIL.n121 12.8005
R435 VTAIL.n163 VTAIL.n162 12.8005
R436 VTAIL.n168 VTAIL.n94 12.8005
R437 VTAIL.n212 VTAIL.n211 12.8005
R438 VTAIL.n253 VTAIL.n252 12.8005
R439 VTAIL.n258 VTAIL.n184 12.8005
R440 VTAIL.n618 VTAIL.n544 12.8005
R441 VTAIL.n613 VTAIL.n548 12.8005
R442 VTAIL.n573 VTAIL.n572 12.8005
R443 VTAIL.n528 VTAIL.n454 12.8005
R444 VTAIL.n523 VTAIL.n458 12.8005
R445 VTAIL.n483 VTAIL.n482 12.8005
R446 VTAIL.n438 VTAIL.n364 12.8005
R447 VTAIL.n433 VTAIL.n368 12.8005
R448 VTAIL.n393 VTAIL.n392 12.8005
R449 VTAIL.n348 VTAIL.n274 12.8005
R450 VTAIL.n343 VTAIL.n278 12.8005
R451 VTAIL.n303 VTAIL.n302 12.8005
R452 VTAIL.n665 VTAIL.n656 12.0247
R453 VTAIL.n701 VTAIL.n638 12.0247
R454 VTAIL.n712 VTAIL.n711 12.0247
R455 VTAIL.n35 VTAIL.n26 12.0247
R456 VTAIL.n71 VTAIL.n8 12.0247
R457 VTAIL.n82 VTAIL.n81 12.0247
R458 VTAIL.n125 VTAIL.n116 12.0247
R459 VTAIL.n161 VTAIL.n98 12.0247
R460 VTAIL.n172 VTAIL.n171 12.0247
R461 VTAIL.n215 VTAIL.n206 12.0247
R462 VTAIL.n251 VTAIL.n188 12.0247
R463 VTAIL.n262 VTAIL.n261 12.0247
R464 VTAIL.n622 VTAIL.n621 12.0247
R465 VTAIL.n612 VTAIL.n549 12.0247
R466 VTAIL.n576 VTAIL.n567 12.0247
R467 VTAIL.n532 VTAIL.n531 12.0247
R468 VTAIL.n522 VTAIL.n459 12.0247
R469 VTAIL.n486 VTAIL.n477 12.0247
R470 VTAIL.n442 VTAIL.n441 12.0247
R471 VTAIL.n432 VTAIL.n369 12.0247
R472 VTAIL.n396 VTAIL.n387 12.0247
R473 VTAIL.n352 VTAIL.n351 12.0247
R474 VTAIL.n342 VTAIL.n279 12.0247
R475 VTAIL.n306 VTAIL.n297 12.0247
R476 VTAIL.n666 VTAIL.n654 11.249
R477 VTAIL.n698 VTAIL.n697 11.249
R478 VTAIL.n715 VTAIL.n632 11.249
R479 VTAIL.n36 VTAIL.n24 11.249
R480 VTAIL.n68 VTAIL.n67 11.249
R481 VTAIL.n85 VTAIL.n2 11.249
R482 VTAIL.n126 VTAIL.n114 11.249
R483 VTAIL.n158 VTAIL.n157 11.249
R484 VTAIL.n175 VTAIL.n92 11.249
R485 VTAIL.n216 VTAIL.n204 11.249
R486 VTAIL.n248 VTAIL.n247 11.249
R487 VTAIL.n265 VTAIL.n182 11.249
R488 VTAIL.n625 VTAIL.n542 11.249
R489 VTAIL.n609 VTAIL.n608 11.249
R490 VTAIL.n577 VTAIL.n565 11.249
R491 VTAIL.n535 VTAIL.n452 11.249
R492 VTAIL.n519 VTAIL.n518 11.249
R493 VTAIL.n487 VTAIL.n475 11.249
R494 VTAIL.n445 VTAIL.n362 11.249
R495 VTAIL.n429 VTAIL.n428 11.249
R496 VTAIL.n397 VTAIL.n385 11.249
R497 VTAIL.n355 VTAIL.n272 11.249
R498 VTAIL.n339 VTAIL.n338 11.249
R499 VTAIL.n307 VTAIL.n295 11.249
R500 VTAIL.n670 VTAIL.n669 10.4732
R501 VTAIL.n694 VTAIL.n640 10.4732
R502 VTAIL.n716 VTAIL.n630 10.4732
R503 VTAIL.n40 VTAIL.n39 10.4732
R504 VTAIL.n64 VTAIL.n10 10.4732
R505 VTAIL.n86 VTAIL.n0 10.4732
R506 VTAIL.n130 VTAIL.n129 10.4732
R507 VTAIL.n154 VTAIL.n100 10.4732
R508 VTAIL.n176 VTAIL.n90 10.4732
R509 VTAIL.n220 VTAIL.n219 10.4732
R510 VTAIL.n244 VTAIL.n190 10.4732
R511 VTAIL.n266 VTAIL.n180 10.4732
R512 VTAIL.n626 VTAIL.n540 10.4732
R513 VTAIL.n605 VTAIL.n551 10.4732
R514 VTAIL.n581 VTAIL.n580 10.4732
R515 VTAIL.n536 VTAIL.n450 10.4732
R516 VTAIL.n515 VTAIL.n461 10.4732
R517 VTAIL.n491 VTAIL.n490 10.4732
R518 VTAIL.n446 VTAIL.n360 10.4732
R519 VTAIL.n425 VTAIL.n371 10.4732
R520 VTAIL.n401 VTAIL.n400 10.4732
R521 VTAIL.n356 VTAIL.n270 10.4732
R522 VTAIL.n335 VTAIL.n281 10.4732
R523 VTAIL.n311 VTAIL.n310 10.4732
R524 VTAIL.n673 VTAIL.n652 9.69747
R525 VTAIL.n693 VTAIL.n642 9.69747
R526 VTAIL.n43 VTAIL.n22 9.69747
R527 VTAIL.n63 VTAIL.n12 9.69747
R528 VTAIL.n133 VTAIL.n112 9.69747
R529 VTAIL.n153 VTAIL.n102 9.69747
R530 VTAIL.n223 VTAIL.n202 9.69747
R531 VTAIL.n243 VTAIL.n192 9.69747
R532 VTAIL.n604 VTAIL.n553 9.69747
R533 VTAIL.n584 VTAIL.n563 9.69747
R534 VTAIL.n514 VTAIL.n463 9.69747
R535 VTAIL.n494 VTAIL.n473 9.69747
R536 VTAIL.n424 VTAIL.n373 9.69747
R537 VTAIL.n404 VTAIL.n383 9.69747
R538 VTAIL.n334 VTAIL.n283 9.69747
R539 VTAIL.n314 VTAIL.n293 9.69747
R540 VTAIL.n718 VTAIL.n717 9.45567
R541 VTAIL.n88 VTAIL.n87 9.45567
R542 VTAIL.n178 VTAIL.n177 9.45567
R543 VTAIL.n268 VTAIL.n267 9.45567
R544 VTAIL.n628 VTAIL.n627 9.45567
R545 VTAIL.n538 VTAIL.n537 9.45567
R546 VTAIL.n448 VTAIL.n447 9.45567
R547 VTAIL.n358 VTAIL.n357 9.45567
R548 VTAIL.n717 VTAIL.n716 9.3005
R549 VTAIL.n632 VTAIL.n631 9.3005
R550 VTAIL.n711 VTAIL.n710 9.3005
R551 VTAIL.n709 VTAIL.n708 9.3005
R552 VTAIL.n648 VTAIL.n647 9.3005
R553 VTAIL.n677 VTAIL.n676 9.3005
R554 VTAIL.n675 VTAIL.n674 9.3005
R555 VTAIL.n652 VTAIL.n651 9.3005
R556 VTAIL.n669 VTAIL.n668 9.3005
R557 VTAIL.n667 VTAIL.n666 9.3005
R558 VTAIL.n656 VTAIL.n655 9.3005
R559 VTAIL.n661 VTAIL.n660 9.3005
R560 VTAIL.n683 VTAIL.n682 9.3005
R561 VTAIL.n685 VTAIL.n684 9.3005
R562 VTAIL.n644 VTAIL.n643 9.3005
R563 VTAIL.n691 VTAIL.n690 9.3005
R564 VTAIL.n693 VTAIL.n692 9.3005
R565 VTAIL.n640 VTAIL.n639 9.3005
R566 VTAIL.n699 VTAIL.n698 9.3005
R567 VTAIL.n701 VTAIL.n700 9.3005
R568 VTAIL.n702 VTAIL.n635 9.3005
R569 VTAIL.n87 VTAIL.n86 9.3005
R570 VTAIL.n2 VTAIL.n1 9.3005
R571 VTAIL.n81 VTAIL.n80 9.3005
R572 VTAIL.n79 VTAIL.n78 9.3005
R573 VTAIL.n18 VTAIL.n17 9.3005
R574 VTAIL.n47 VTAIL.n46 9.3005
R575 VTAIL.n45 VTAIL.n44 9.3005
R576 VTAIL.n22 VTAIL.n21 9.3005
R577 VTAIL.n39 VTAIL.n38 9.3005
R578 VTAIL.n37 VTAIL.n36 9.3005
R579 VTAIL.n26 VTAIL.n25 9.3005
R580 VTAIL.n31 VTAIL.n30 9.3005
R581 VTAIL.n53 VTAIL.n52 9.3005
R582 VTAIL.n55 VTAIL.n54 9.3005
R583 VTAIL.n14 VTAIL.n13 9.3005
R584 VTAIL.n61 VTAIL.n60 9.3005
R585 VTAIL.n63 VTAIL.n62 9.3005
R586 VTAIL.n10 VTAIL.n9 9.3005
R587 VTAIL.n69 VTAIL.n68 9.3005
R588 VTAIL.n71 VTAIL.n70 9.3005
R589 VTAIL.n72 VTAIL.n5 9.3005
R590 VTAIL.n177 VTAIL.n176 9.3005
R591 VTAIL.n92 VTAIL.n91 9.3005
R592 VTAIL.n171 VTAIL.n170 9.3005
R593 VTAIL.n169 VTAIL.n168 9.3005
R594 VTAIL.n108 VTAIL.n107 9.3005
R595 VTAIL.n137 VTAIL.n136 9.3005
R596 VTAIL.n135 VTAIL.n134 9.3005
R597 VTAIL.n112 VTAIL.n111 9.3005
R598 VTAIL.n129 VTAIL.n128 9.3005
R599 VTAIL.n127 VTAIL.n126 9.3005
R600 VTAIL.n116 VTAIL.n115 9.3005
R601 VTAIL.n121 VTAIL.n120 9.3005
R602 VTAIL.n143 VTAIL.n142 9.3005
R603 VTAIL.n145 VTAIL.n144 9.3005
R604 VTAIL.n104 VTAIL.n103 9.3005
R605 VTAIL.n151 VTAIL.n150 9.3005
R606 VTAIL.n153 VTAIL.n152 9.3005
R607 VTAIL.n100 VTAIL.n99 9.3005
R608 VTAIL.n159 VTAIL.n158 9.3005
R609 VTAIL.n161 VTAIL.n160 9.3005
R610 VTAIL.n162 VTAIL.n95 9.3005
R611 VTAIL.n267 VTAIL.n266 9.3005
R612 VTAIL.n182 VTAIL.n181 9.3005
R613 VTAIL.n261 VTAIL.n260 9.3005
R614 VTAIL.n259 VTAIL.n258 9.3005
R615 VTAIL.n198 VTAIL.n197 9.3005
R616 VTAIL.n227 VTAIL.n226 9.3005
R617 VTAIL.n225 VTAIL.n224 9.3005
R618 VTAIL.n202 VTAIL.n201 9.3005
R619 VTAIL.n219 VTAIL.n218 9.3005
R620 VTAIL.n217 VTAIL.n216 9.3005
R621 VTAIL.n206 VTAIL.n205 9.3005
R622 VTAIL.n211 VTAIL.n210 9.3005
R623 VTAIL.n233 VTAIL.n232 9.3005
R624 VTAIL.n235 VTAIL.n234 9.3005
R625 VTAIL.n194 VTAIL.n193 9.3005
R626 VTAIL.n241 VTAIL.n240 9.3005
R627 VTAIL.n243 VTAIL.n242 9.3005
R628 VTAIL.n190 VTAIL.n189 9.3005
R629 VTAIL.n249 VTAIL.n248 9.3005
R630 VTAIL.n251 VTAIL.n250 9.3005
R631 VTAIL.n252 VTAIL.n185 9.3005
R632 VTAIL.n596 VTAIL.n595 9.3005
R633 VTAIL.n555 VTAIL.n554 9.3005
R634 VTAIL.n602 VTAIL.n601 9.3005
R635 VTAIL.n604 VTAIL.n603 9.3005
R636 VTAIL.n551 VTAIL.n550 9.3005
R637 VTAIL.n610 VTAIL.n609 9.3005
R638 VTAIL.n612 VTAIL.n611 9.3005
R639 VTAIL.n548 VTAIL.n545 9.3005
R640 VTAIL.n627 VTAIL.n626 9.3005
R641 VTAIL.n542 VTAIL.n541 9.3005
R642 VTAIL.n621 VTAIL.n620 9.3005
R643 VTAIL.n619 VTAIL.n618 9.3005
R644 VTAIL.n594 VTAIL.n593 9.3005
R645 VTAIL.n559 VTAIL.n558 9.3005
R646 VTAIL.n588 VTAIL.n587 9.3005
R647 VTAIL.n586 VTAIL.n585 9.3005
R648 VTAIL.n563 VTAIL.n562 9.3005
R649 VTAIL.n580 VTAIL.n579 9.3005
R650 VTAIL.n578 VTAIL.n577 9.3005
R651 VTAIL.n567 VTAIL.n566 9.3005
R652 VTAIL.n572 VTAIL.n571 9.3005
R653 VTAIL.n506 VTAIL.n505 9.3005
R654 VTAIL.n465 VTAIL.n464 9.3005
R655 VTAIL.n512 VTAIL.n511 9.3005
R656 VTAIL.n514 VTAIL.n513 9.3005
R657 VTAIL.n461 VTAIL.n460 9.3005
R658 VTAIL.n520 VTAIL.n519 9.3005
R659 VTAIL.n522 VTAIL.n521 9.3005
R660 VTAIL.n458 VTAIL.n455 9.3005
R661 VTAIL.n537 VTAIL.n536 9.3005
R662 VTAIL.n452 VTAIL.n451 9.3005
R663 VTAIL.n531 VTAIL.n530 9.3005
R664 VTAIL.n529 VTAIL.n528 9.3005
R665 VTAIL.n504 VTAIL.n503 9.3005
R666 VTAIL.n469 VTAIL.n468 9.3005
R667 VTAIL.n498 VTAIL.n497 9.3005
R668 VTAIL.n496 VTAIL.n495 9.3005
R669 VTAIL.n473 VTAIL.n472 9.3005
R670 VTAIL.n490 VTAIL.n489 9.3005
R671 VTAIL.n488 VTAIL.n487 9.3005
R672 VTAIL.n477 VTAIL.n476 9.3005
R673 VTAIL.n482 VTAIL.n481 9.3005
R674 VTAIL.n416 VTAIL.n415 9.3005
R675 VTAIL.n375 VTAIL.n374 9.3005
R676 VTAIL.n422 VTAIL.n421 9.3005
R677 VTAIL.n424 VTAIL.n423 9.3005
R678 VTAIL.n371 VTAIL.n370 9.3005
R679 VTAIL.n430 VTAIL.n429 9.3005
R680 VTAIL.n432 VTAIL.n431 9.3005
R681 VTAIL.n368 VTAIL.n365 9.3005
R682 VTAIL.n447 VTAIL.n446 9.3005
R683 VTAIL.n362 VTAIL.n361 9.3005
R684 VTAIL.n441 VTAIL.n440 9.3005
R685 VTAIL.n439 VTAIL.n438 9.3005
R686 VTAIL.n414 VTAIL.n413 9.3005
R687 VTAIL.n379 VTAIL.n378 9.3005
R688 VTAIL.n408 VTAIL.n407 9.3005
R689 VTAIL.n406 VTAIL.n405 9.3005
R690 VTAIL.n383 VTAIL.n382 9.3005
R691 VTAIL.n400 VTAIL.n399 9.3005
R692 VTAIL.n398 VTAIL.n397 9.3005
R693 VTAIL.n387 VTAIL.n386 9.3005
R694 VTAIL.n392 VTAIL.n391 9.3005
R695 VTAIL.n326 VTAIL.n325 9.3005
R696 VTAIL.n285 VTAIL.n284 9.3005
R697 VTAIL.n332 VTAIL.n331 9.3005
R698 VTAIL.n334 VTAIL.n333 9.3005
R699 VTAIL.n281 VTAIL.n280 9.3005
R700 VTAIL.n340 VTAIL.n339 9.3005
R701 VTAIL.n342 VTAIL.n341 9.3005
R702 VTAIL.n278 VTAIL.n275 9.3005
R703 VTAIL.n357 VTAIL.n356 9.3005
R704 VTAIL.n272 VTAIL.n271 9.3005
R705 VTAIL.n351 VTAIL.n350 9.3005
R706 VTAIL.n349 VTAIL.n348 9.3005
R707 VTAIL.n324 VTAIL.n323 9.3005
R708 VTAIL.n289 VTAIL.n288 9.3005
R709 VTAIL.n318 VTAIL.n317 9.3005
R710 VTAIL.n316 VTAIL.n315 9.3005
R711 VTAIL.n293 VTAIL.n292 9.3005
R712 VTAIL.n310 VTAIL.n309 9.3005
R713 VTAIL.n308 VTAIL.n307 9.3005
R714 VTAIL.n297 VTAIL.n296 9.3005
R715 VTAIL.n302 VTAIL.n301 9.3005
R716 VTAIL.n674 VTAIL.n650 8.92171
R717 VTAIL.n690 VTAIL.n689 8.92171
R718 VTAIL.n44 VTAIL.n20 8.92171
R719 VTAIL.n60 VTAIL.n59 8.92171
R720 VTAIL.n134 VTAIL.n110 8.92171
R721 VTAIL.n150 VTAIL.n149 8.92171
R722 VTAIL.n224 VTAIL.n200 8.92171
R723 VTAIL.n240 VTAIL.n239 8.92171
R724 VTAIL.n601 VTAIL.n600 8.92171
R725 VTAIL.n585 VTAIL.n561 8.92171
R726 VTAIL.n511 VTAIL.n510 8.92171
R727 VTAIL.n495 VTAIL.n471 8.92171
R728 VTAIL.n421 VTAIL.n420 8.92171
R729 VTAIL.n405 VTAIL.n381 8.92171
R730 VTAIL.n331 VTAIL.n330 8.92171
R731 VTAIL.n315 VTAIL.n291 8.92171
R732 VTAIL.n678 VTAIL.n677 8.14595
R733 VTAIL.n686 VTAIL.n644 8.14595
R734 VTAIL.n48 VTAIL.n47 8.14595
R735 VTAIL.n56 VTAIL.n14 8.14595
R736 VTAIL.n138 VTAIL.n137 8.14595
R737 VTAIL.n146 VTAIL.n104 8.14595
R738 VTAIL.n228 VTAIL.n227 8.14595
R739 VTAIL.n236 VTAIL.n194 8.14595
R740 VTAIL.n597 VTAIL.n555 8.14595
R741 VTAIL.n589 VTAIL.n588 8.14595
R742 VTAIL.n507 VTAIL.n465 8.14595
R743 VTAIL.n499 VTAIL.n498 8.14595
R744 VTAIL.n417 VTAIL.n375 8.14595
R745 VTAIL.n409 VTAIL.n408 8.14595
R746 VTAIL.n327 VTAIL.n285 8.14595
R747 VTAIL.n319 VTAIL.n318 8.14595
R748 VTAIL.n681 VTAIL.n648 7.3702
R749 VTAIL.n685 VTAIL.n646 7.3702
R750 VTAIL.n51 VTAIL.n18 7.3702
R751 VTAIL.n55 VTAIL.n16 7.3702
R752 VTAIL.n141 VTAIL.n108 7.3702
R753 VTAIL.n145 VTAIL.n106 7.3702
R754 VTAIL.n231 VTAIL.n198 7.3702
R755 VTAIL.n235 VTAIL.n196 7.3702
R756 VTAIL.n596 VTAIL.n557 7.3702
R757 VTAIL.n592 VTAIL.n559 7.3702
R758 VTAIL.n506 VTAIL.n467 7.3702
R759 VTAIL.n502 VTAIL.n469 7.3702
R760 VTAIL.n416 VTAIL.n377 7.3702
R761 VTAIL.n412 VTAIL.n379 7.3702
R762 VTAIL.n326 VTAIL.n287 7.3702
R763 VTAIL.n322 VTAIL.n289 7.3702
R764 VTAIL.n682 VTAIL.n681 6.59444
R765 VTAIL.n682 VTAIL.n646 6.59444
R766 VTAIL.n52 VTAIL.n51 6.59444
R767 VTAIL.n52 VTAIL.n16 6.59444
R768 VTAIL.n142 VTAIL.n141 6.59444
R769 VTAIL.n142 VTAIL.n106 6.59444
R770 VTAIL.n232 VTAIL.n231 6.59444
R771 VTAIL.n232 VTAIL.n196 6.59444
R772 VTAIL.n593 VTAIL.n557 6.59444
R773 VTAIL.n593 VTAIL.n592 6.59444
R774 VTAIL.n503 VTAIL.n467 6.59444
R775 VTAIL.n503 VTAIL.n502 6.59444
R776 VTAIL.n413 VTAIL.n377 6.59444
R777 VTAIL.n413 VTAIL.n412 6.59444
R778 VTAIL.n323 VTAIL.n287 6.59444
R779 VTAIL.n323 VTAIL.n322 6.59444
R780 VTAIL.n678 VTAIL.n648 5.81868
R781 VTAIL.n686 VTAIL.n685 5.81868
R782 VTAIL.n48 VTAIL.n18 5.81868
R783 VTAIL.n56 VTAIL.n55 5.81868
R784 VTAIL.n138 VTAIL.n108 5.81868
R785 VTAIL.n146 VTAIL.n145 5.81868
R786 VTAIL.n228 VTAIL.n198 5.81868
R787 VTAIL.n236 VTAIL.n235 5.81868
R788 VTAIL.n597 VTAIL.n596 5.81868
R789 VTAIL.n589 VTAIL.n559 5.81868
R790 VTAIL.n507 VTAIL.n506 5.81868
R791 VTAIL.n499 VTAIL.n469 5.81868
R792 VTAIL.n417 VTAIL.n416 5.81868
R793 VTAIL.n409 VTAIL.n379 5.81868
R794 VTAIL.n327 VTAIL.n326 5.81868
R795 VTAIL.n319 VTAIL.n289 5.81868
R796 VTAIL.n677 VTAIL.n650 5.04292
R797 VTAIL.n689 VTAIL.n644 5.04292
R798 VTAIL.n47 VTAIL.n20 5.04292
R799 VTAIL.n59 VTAIL.n14 5.04292
R800 VTAIL.n137 VTAIL.n110 5.04292
R801 VTAIL.n149 VTAIL.n104 5.04292
R802 VTAIL.n227 VTAIL.n200 5.04292
R803 VTAIL.n239 VTAIL.n194 5.04292
R804 VTAIL.n600 VTAIL.n555 5.04292
R805 VTAIL.n588 VTAIL.n561 5.04292
R806 VTAIL.n510 VTAIL.n465 5.04292
R807 VTAIL.n498 VTAIL.n471 5.04292
R808 VTAIL.n420 VTAIL.n375 5.04292
R809 VTAIL.n408 VTAIL.n381 5.04292
R810 VTAIL.n330 VTAIL.n285 5.04292
R811 VTAIL.n318 VTAIL.n291 5.04292
R812 VTAIL.n660 VTAIL.n659 4.38563
R813 VTAIL.n30 VTAIL.n29 4.38563
R814 VTAIL.n120 VTAIL.n119 4.38563
R815 VTAIL.n210 VTAIL.n209 4.38563
R816 VTAIL.n571 VTAIL.n570 4.38563
R817 VTAIL.n481 VTAIL.n480 4.38563
R818 VTAIL.n391 VTAIL.n390 4.38563
R819 VTAIL.n301 VTAIL.n300 4.38563
R820 VTAIL.n674 VTAIL.n673 4.26717
R821 VTAIL.n690 VTAIL.n642 4.26717
R822 VTAIL.n44 VTAIL.n43 4.26717
R823 VTAIL.n60 VTAIL.n12 4.26717
R824 VTAIL.n134 VTAIL.n133 4.26717
R825 VTAIL.n150 VTAIL.n102 4.26717
R826 VTAIL.n224 VTAIL.n223 4.26717
R827 VTAIL.n240 VTAIL.n192 4.26717
R828 VTAIL.n601 VTAIL.n553 4.26717
R829 VTAIL.n585 VTAIL.n584 4.26717
R830 VTAIL.n511 VTAIL.n463 4.26717
R831 VTAIL.n495 VTAIL.n494 4.26717
R832 VTAIL.n421 VTAIL.n373 4.26717
R833 VTAIL.n405 VTAIL.n404 4.26717
R834 VTAIL.n331 VTAIL.n283 4.26717
R835 VTAIL.n315 VTAIL.n314 4.26717
R836 VTAIL.n670 VTAIL.n652 3.49141
R837 VTAIL.n694 VTAIL.n693 3.49141
R838 VTAIL.n718 VTAIL.n630 3.49141
R839 VTAIL.n40 VTAIL.n22 3.49141
R840 VTAIL.n64 VTAIL.n63 3.49141
R841 VTAIL.n88 VTAIL.n0 3.49141
R842 VTAIL.n130 VTAIL.n112 3.49141
R843 VTAIL.n154 VTAIL.n153 3.49141
R844 VTAIL.n178 VTAIL.n90 3.49141
R845 VTAIL.n220 VTAIL.n202 3.49141
R846 VTAIL.n244 VTAIL.n243 3.49141
R847 VTAIL.n268 VTAIL.n180 3.49141
R848 VTAIL.n628 VTAIL.n540 3.49141
R849 VTAIL.n605 VTAIL.n604 3.49141
R850 VTAIL.n581 VTAIL.n563 3.49141
R851 VTAIL.n538 VTAIL.n450 3.49141
R852 VTAIL.n515 VTAIL.n514 3.49141
R853 VTAIL.n491 VTAIL.n473 3.49141
R854 VTAIL.n448 VTAIL.n360 3.49141
R855 VTAIL.n425 VTAIL.n424 3.49141
R856 VTAIL.n401 VTAIL.n383 3.49141
R857 VTAIL.n358 VTAIL.n270 3.49141
R858 VTAIL.n335 VTAIL.n334 3.49141
R859 VTAIL.n311 VTAIL.n293 3.49141
R860 VTAIL.n449 VTAIL.n359 3.38843
R861 VTAIL.n629 VTAIL.n539 3.38843
R862 VTAIL.n269 VTAIL.n179 3.38843
R863 VTAIL.n669 VTAIL.n654 2.71565
R864 VTAIL.n697 VTAIL.n640 2.71565
R865 VTAIL.n716 VTAIL.n715 2.71565
R866 VTAIL.n39 VTAIL.n24 2.71565
R867 VTAIL.n67 VTAIL.n10 2.71565
R868 VTAIL.n86 VTAIL.n85 2.71565
R869 VTAIL.n129 VTAIL.n114 2.71565
R870 VTAIL.n157 VTAIL.n100 2.71565
R871 VTAIL.n176 VTAIL.n175 2.71565
R872 VTAIL.n219 VTAIL.n204 2.71565
R873 VTAIL.n247 VTAIL.n190 2.71565
R874 VTAIL.n266 VTAIL.n265 2.71565
R875 VTAIL.n626 VTAIL.n625 2.71565
R876 VTAIL.n608 VTAIL.n551 2.71565
R877 VTAIL.n580 VTAIL.n565 2.71565
R878 VTAIL.n536 VTAIL.n535 2.71565
R879 VTAIL.n518 VTAIL.n461 2.71565
R880 VTAIL.n490 VTAIL.n475 2.71565
R881 VTAIL.n446 VTAIL.n445 2.71565
R882 VTAIL.n428 VTAIL.n371 2.71565
R883 VTAIL.n400 VTAIL.n385 2.71565
R884 VTAIL.n356 VTAIL.n355 2.71565
R885 VTAIL.n338 VTAIL.n281 2.71565
R886 VTAIL.n310 VTAIL.n295 2.71565
R887 VTAIL.n666 VTAIL.n665 1.93989
R888 VTAIL.n698 VTAIL.n638 1.93989
R889 VTAIL.n712 VTAIL.n632 1.93989
R890 VTAIL.n36 VTAIL.n35 1.93989
R891 VTAIL.n68 VTAIL.n8 1.93989
R892 VTAIL.n82 VTAIL.n2 1.93989
R893 VTAIL.n126 VTAIL.n125 1.93989
R894 VTAIL.n158 VTAIL.n98 1.93989
R895 VTAIL.n172 VTAIL.n92 1.93989
R896 VTAIL.n216 VTAIL.n215 1.93989
R897 VTAIL.n248 VTAIL.n188 1.93989
R898 VTAIL.n262 VTAIL.n182 1.93989
R899 VTAIL.n622 VTAIL.n542 1.93989
R900 VTAIL.n609 VTAIL.n549 1.93989
R901 VTAIL.n577 VTAIL.n576 1.93989
R902 VTAIL.n532 VTAIL.n452 1.93989
R903 VTAIL.n519 VTAIL.n459 1.93989
R904 VTAIL.n487 VTAIL.n486 1.93989
R905 VTAIL.n442 VTAIL.n362 1.93989
R906 VTAIL.n429 VTAIL.n369 1.93989
R907 VTAIL.n397 VTAIL.n396 1.93989
R908 VTAIL.n352 VTAIL.n272 1.93989
R909 VTAIL.n339 VTAIL.n279 1.93989
R910 VTAIL.n307 VTAIL.n306 1.93989
R911 VTAIL VTAIL.n89 1.75266
R912 VTAIL VTAIL.n719 1.63628
R913 VTAIL.n662 VTAIL.n656 1.16414
R914 VTAIL.n703 VTAIL.n701 1.16414
R915 VTAIL.n711 VTAIL.n634 1.16414
R916 VTAIL.n32 VTAIL.n26 1.16414
R917 VTAIL.n73 VTAIL.n71 1.16414
R918 VTAIL.n81 VTAIL.n4 1.16414
R919 VTAIL.n122 VTAIL.n116 1.16414
R920 VTAIL.n163 VTAIL.n161 1.16414
R921 VTAIL.n171 VTAIL.n94 1.16414
R922 VTAIL.n212 VTAIL.n206 1.16414
R923 VTAIL.n253 VTAIL.n251 1.16414
R924 VTAIL.n261 VTAIL.n184 1.16414
R925 VTAIL.n621 VTAIL.n544 1.16414
R926 VTAIL.n613 VTAIL.n612 1.16414
R927 VTAIL.n573 VTAIL.n567 1.16414
R928 VTAIL.n531 VTAIL.n454 1.16414
R929 VTAIL.n523 VTAIL.n522 1.16414
R930 VTAIL.n483 VTAIL.n477 1.16414
R931 VTAIL.n441 VTAIL.n364 1.16414
R932 VTAIL.n433 VTAIL.n432 1.16414
R933 VTAIL.n393 VTAIL.n387 1.16414
R934 VTAIL.n351 VTAIL.n274 1.16414
R935 VTAIL.n343 VTAIL.n342 1.16414
R936 VTAIL.n303 VTAIL.n297 1.16414
R937 VTAIL.n539 VTAIL.n449 0.470328
R938 VTAIL.n179 VTAIL.n89 0.470328
R939 VTAIL.n661 VTAIL.n658 0.388379
R940 VTAIL.n702 VTAIL.n636 0.388379
R941 VTAIL.n708 VTAIL.n707 0.388379
R942 VTAIL.n31 VTAIL.n28 0.388379
R943 VTAIL.n72 VTAIL.n6 0.388379
R944 VTAIL.n78 VTAIL.n77 0.388379
R945 VTAIL.n121 VTAIL.n118 0.388379
R946 VTAIL.n162 VTAIL.n96 0.388379
R947 VTAIL.n168 VTAIL.n167 0.388379
R948 VTAIL.n211 VTAIL.n208 0.388379
R949 VTAIL.n252 VTAIL.n186 0.388379
R950 VTAIL.n258 VTAIL.n257 0.388379
R951 VTAIL.n618 VTAIL.n617 0.388379
R952 VTAIL.n548 VTAIL.n546 0.388379
R953 VTAIL.n572 VTAIL.n569 0.388379
R954 VTAIL.n528 VTAIL.n527 0.388379
R955 VTAIL.n458 VTAIL.n456 0.388379
R956 VTAIL.n482 VTAIL.n479 0.388379
R957 VTAIL.n438 VTAIL.n437 0.388379
R958 VTAIL.n368 VTAIL.n366 0.388379
R959 VTAIL.n392 VTAIL.n389 0.388379
R960 VTAIL.n348 VTAIL.n347 0.388379
R961 VTAIL.n278 VTAIL.n276 0.388379
R962 VTAIL.n302 VTAIL.n299 0.388379
R963 VTAIL.n660 VTAIL.n655 0.155672
R964 VTAIL.n667 VTAIL.n655 0.155672
R965 VTAIL.n668 VTAIL.n667 0.155672
R966 VTAIL.n668 VTAIL.n651 0.155672
R967 VTAIL.n675 VTAIL.n651 0.155672
R968 VTAIL.n676 VTAIL.n675 0.155672
R969 VTAIL.n676 VTAIL.n647 0.155672
R970 VTAIL.n683 VTAIL.n647 0.155672
R971 VTAIL.n684 VTAIL.n683 0.155672
R972 VTAIL.n684 VTAIL.n643 0.155672
R973 VTAIL.n691 VTAIL.n643 0.155672
R974 VTAIL.n692 VTAIL.n691 0.155672
R975 VTAIL.n692 VTAIL.n639 0.155672
R976 VTAIL.n699 VTAIL.n639 0.155672
R977 VTAIL.n700 VTAIL.n699 0.155672
R978 VTAIL.n700 VTAIL.n635 0.155672
R979 VTAIL.n709 VTAIL.n635 0.155672
R980 VTAIL.n710 VTAIL.n709 0.155672
R981 VTAIL.n710 VTAIL.n631 0.155672
R982 VTAIL.n717 VTAIL.n631 0.155672
R983 VTAIL.n30 VTAIL.n25 0.155672
R984 VTAIL.n37 VTAIL.n25 0.155672
R985 VTAIL.n38 VTAIL.n37 0.155672
R986 VTAIL.n38 VTAIL.n21 0.155672
R987 VTAIL.n45 VTAIL.n21 0.155672
R988 VTAIL.n46 VTAIL.n45 0.155672
R989 VTAIL.n46 VTAIL.n17 0.155672
R990 VTAIL.n53 VTAIL.n17 0.155672
R991 VTAIL.n54 VTAIL.n53 0.155672
R992 VTAIL.n54 VTAIL.n13 0.155672
R993 VTAIL.n61 VTAIL.n13 0.155672
R994 VTAIL.n62 VTAIL.n61 0.155672
R995 VTAIL.n62 VTAIL.n9 0.155672
R996 VTAIL.n69 VTAIL.n9 0.155672
R997 VTAIL.n70 VTAIL.n69 0.155672
R998 VTAIL.n70 VTAIL.n5 0.155672
R999 VTAIL.n79 VTAIL.n5 0.155672
R1000 VTAIL.n80 VTAIL.n79 0.155672
R1001 VTAIL.n80 VTAIL.n1 0.155672
R1002 VTAIL.n87 VTAIL.n1 0.155672
R1003 VTAIL.n120 VTAIL.n115 0.155672
R1004 VTAIL.n127 VTAIL.n115 0.155672
R1005 VTAIL.n128 VTAIL.n127 0.155672
R1006 VTAIL.n128 VTAIL.n111 0.155672
R1007 VTAIL.n135 VTAIL.n111 0.155672
R1008 VTAIL.n136 VTAIL.n135 0.155672
R1009 VTAIL.n136 VTAIL.n107 0.155672
R1010 VTAIL.n143 VTAIL.n107 0.155672
R1011 VTAIL.n144 VTAIL.n143 0.155672
R1012 VTAIL.n144 VTAIL.n103 0.155672
R1013 VTAIL.n151 VTAIL.n103 0.155672
R1014 VTAIL.n152 VTAIL.n151 0.155672
R1015 VTAIL.n152 VTAIL.n99 0.155672
R1016 VTAIL.n159 VTAIL.n99 0.155672
R1017 VTAIL.n160 VTAIL.n159 0.155672
R1018 VTAIL.n160 VTAIL.n95 0.155672
R1019 VTAIL.n169 VTAIL.n95 0.155672
R1020 VTAIL.n170 VTAIL.n169 0.155672
R1021 VTAIL.n170 VTAIL.n91 0.155672
R1022 VTAIL.n177 VTAIL.n91 0.155672
R1023 VTAIL.n210 VTAIL.n205 0.155672
R1024 VTAIL.n217 VTAIL.n205 0.155672
R1025 VTAIL.n218 VTAIL.n217 0.155672
R1026 VTAIL.n218 VTAIL.n201 0.155672
R1027 VTAIL.n225 VTAIL.n201 0.155672
R1028 VTAIL.n226 VTAIL.n225 0.155672
R1029 VTAIL.n226 VTAIL.n197 0.155672
R1030 VTAIL.n233 VTAIL.n197 0.155672
R1031 VTAIL.n234 VTAIL.n233 0.155672
R1032 VTAIL.n234 VTAIL.n193 0.155672
R1033 VTAIL.n241 VTAIL.n193 0.155672
R1034 VTAIL.n242 VTAIL.n241 0.155672
R1035 VTAIL.n242 VTAIL.n189 0.155672
R1036 VTAIL.n249 VTAIL.n189 0.155672
R1037 VTAIL.n250 VTAIL.n249 0.155672
R1038 VTAIL.n250 VTAIL.n185 0.155672
R1039 VTAIL.n259 VTAIL.n185 0.155672
R1040 VTAIL.n260 VTAIL.n259 0.155672
R1041 VTAIL.n260 VTAIL.n181 0.155672
R1042 VTAIL.n267 VTAIL.n181 0.155672
R1043 VTAIL.n627 VTAIL.n541 0.155672
R1044 VTAIL.n620 VTAIL.n541 0.155672
R1045 VTAIL.n620 VTAIL.n619 0.155672
R1046 VTAIL.n619 VTAIL.n545 0.155672
R1047 VTAIL.n611 VTAIL.n545 0.155672
R1048 VTAIL.n611 VTAIL.n610 0.155672
R1049 VTAIL.n610 VTAIL.n550 0.155672
R1050 VTAIL.n603 VTAIL.n550 0.155672
R1051 VTAIL.n603 VTAIL.n602 0.155672
R1052 VTAIL.n602 VTAIL.n554 0.155672
R1053 VTAIL.n595 VTAIL.n554 0.155672
R1054 VTAIL.n595 VTAIL.n594 0.155672
R1055 VTAIL.n594 VTAIL.n558 0.155672
R1056 VTAIL.n587 VTAIL.n558 0.155672
R1057 VTAIL.n587 VTAIL.n586 0.155672
R1058 VTAIL.n586 VTAIL.n562 0.155672
R1059 VTAIL.n579 VTAIL.n562 0.155672
R1060 VTAIL.n579 VTAIL.n578 0.155672
R1061 VTAIL.n578 VTAIL.n566 0.155672
R1062 VTAIL.n571 VTAIL.n566 0.155672
R1063 VTAIL.n537 VTAIL.n451 0.155672
R1064 VTAIL.n530 VTAIL.n451 0.155672
R1065 VTAIL.n530 VTAIL.n529 0.155672
R1066 VTAIL.n529 VTAIL.n455 0.155672
R1067 VTAIL.n521 VTAIL.n455 0.155672
R1068 VTAIL.n521 VTAIL.n520 0.155672
R1069 VTAIL.n520 VTAIL.n460 0.155672
R1070 VTAIL.n513 VTAIL.n460 0.155672
R1071 VTAIL.n513 VTAIL.n512 0.155672
R1072 VTAIL.n512 VTAIL.n464 0.155672
R1073 VTAIL.n505 VTAIL.n464 0.155672
R1074 VTAIL.n505 VTAIL.n504 0.155672
R1075 VTAIL.n504 VTAIL.n468 0.155672
R1076 VTAIL.n497 VTAIL.n468 0.155672
R1077 VTAIL.n497 VTAIL.n496 0.155672
R1078 VTAIL.n496 VTAIL.n472 0.155672
R1079 VTAIL.n489 VTAIL.n472 0.155672
R1080 VTAIL.n489 VTAIL.n488 0.155672
R1081 VTAIL.n488 VTAIL.n476 0.155672
R1082 VTAIL.n481 VTAIL.n476 0.155672
R1083 VTAIL.n447 VTAIL.n361 0.155672
R1084 VTAIL.n440 VTAIL.n361 0.155672
R1085 VTAIL.n440 VTAIL.n439 0.155672
R1086 VTAIL.n439 VTAIL.n365 0.155672
R1087 VTAIL.n431 VTAIL.n365 0.155672
R1088 VTAIL.n431 VTAIL.n430 0.155672
R1089 VTAIL.n430 VTAIL.n370 0.155672
R1090 VTAIL.n423 VTAIL.n370 0.155672
R1091 VTAIL.n423 VTAIL.n422 0.155672
R1092 VTAIL.n422 VTAIL.n374 0.155672
R1093 VTAIL.n415 VTAIL.n374 0.155672
R1094 VTAIL.n415 VTAIL.n414 0.155672
R1095 VTAIL.n414 VTAIL.n378 0.155672
R1096 VTAIL.n407 VTAIL.n378 0.155672
R1097 VTAIL.n407 VTAIL.n406 0.155672
R1098 VTAIL.n406 VTAIL.n382 0.155672
R1099 VTAIL.n399 VTAIL.n382 0.155672
R1100 VTAIL.n399 VTAIL.n398 0.155672
R1101 VTAIL.n398 VTAIL.n386 0.155672
R1102 VTAIL.n391 VTAIL.n386 0.155672
R1103 VTAIL.n357 VTAIL.n271 0.155672
R1104 VTAIL.n350 VTAIL.n271 0.155672
R1105 VTAIL.n350 VTAIL.n349 0.155672
R1106 VTAIL.n349 VTAIL.n275 0.155672
R1107 VTAIL.n341 VTAIL.n275 0.155672
R1108 VTAIL.n341 VTAIL.n340 0.155672
R1109 VTAIL.n340 VTAIL.n280 0.155672
R1110 VTAIL.n333 VTAIL.n280 0.155672
R1111 VTAIL.n333 VTAIL.n332 0.155672
R1112 VTAIL.n332 VTAIL.n284 0.155672
R1113 VTAIL.n325 VTAIL.n284 0.155672
R1114 VTAIL.n325 VTAIL.n324 0.155672
R1115 VTAIL.n324 VTAIL.n288 0.155672
R1116 VTAIL.n317 VTAIL.n288 0.155672
R1117 VTAIL.n317 VTAIL.n316 0.155672
R1118 VTAIL.n316 VTAIL.n292 0.155672
R1119 VTAIL.n309 VTAIL.n292 0.155672
R1120 VTAIL.n309 VTAIL.n308 0.155672
R1121 VTAIL.n308 VTAIL.n296 0.155672
R1122 VTAIL.n301 VTAIL.n296 0.155672
R1123 VDD1 VDD1.n1 108.841
R1124 VDD1 VDD1.n0 60.6418
R1125 VDD1.n0 VDD1.t0 1.23261
R1126 VDD1.n0 VDD1.t3 1.23261
R1127 VDD1.n1 VDD1.t2 1.23261
R1128 VDD1.n1 VDD1.t1 1.23261
R1129 B.n940 B.n939 585
R1130 B.n941 B.n940 585
R1131 B.n373 B.n139 585
R1132 B.n372 B.n371 585
R1133 B.n370 B.n369 585
R1134 B.n368 B.n367 585
R1135 B.n366 B.n365 585
R1136 B.n364 B.n363 585
R1137 B.n362 B.n361 585
R1138 B.n360 B.n359 585
R1139 B.n358 B.n357 585
R1140 B.n356 B.n355 585
R1141 B.n354 B.n353 585
R1142 B.n352 B.n351 585
R1143 B.n350 B.n349 585
R1144 B.n348 B.n347 585
R1145 B.n346 B.n345 585
R1146 B.n344 B.n343 585
R1147 B.n342 B.n341 585
R1148 B.n340 B.n339 585
R1149 B.n338 B.n337 585
R1150 B.n336 B.n335 585
R1151 B.n334 B.n333 585
R1152 B.n332 B.n331 585
R1153 B.n330 B.n329 585
R1154 B.n328 B.n327 585
R1155 B.n326 B.n325 585
R1156 B.n324 B.n323 585
R1157 B.n322 B.n321 585
R1158 B.n320 B.n319 585
R1159 B.n318 B.n317 585
R1160 B.n316 B.n315 585
R1161 B.n314 B.n313 585
R1162 B.n312 B.n311 585
R1163 B.n310 B.n309 585
R1164 B.n308 B.n307 585
R1165 B.n306 B.n305 585
R1166 B.n304 B.n303 585
R1167 B.n302 B.n301 585
R1168 B.n300 B.n299 585
R1169 B.n298 B.n297 585
R1170 B.n296 B.n295 585
R1171 B.n294 B.n293 585
R1172 B.n292 B.n291 585
R1173 B.n290 B.n289 585
R1174 B.n288 B.n287 585
R1175 B.n286 B.n285 585
R1176 B.n284 B.n283 585
R1177 B.n282 B.n281 585
R1178 B.n280 B.n279 585
R1179 B.n278 B.n277 585
R1180 B.n276 B.n275 585
R1181 B.n274 B.n273 585
R1182 B.n272 B.n271 585
R1183 B.n270 B.n269 585
R1184 B.n267 B.n266 585
R1185 B.n265 B.n264 585
R1186 B.n263 B.n262 585
R1187 B.n261 B.n260 585
R1188 B.n259 B.n258 585
R1189 B.n257 B.n256 585
R1190 B.n255 B.n254 585
R1191 B.n253 B.n252 585
R1192 B.n251 B.n250 585
R1193 B.n249 B.n248 585
R1194 B.n247 B.n246 585
R1195 B.n245 B.n244 585
R1196 B.n243 B.n242 585
R1197 B.n241 B.n240 585
R1198 B.n239 B.n238 585
R1199 B.n237 B.n236 585
R1200 B.n235 B.n234 585
R1201 B.n233 B.n232 585
R1202 B.n231 B.n230 585
R1203 B.n229 B.n228 585
R1204 B.n227 B.n226 585
R1205 B.n225 B.n224 585
R1206 B.n223 B.n222 585
R1207 B.n221 B.n220 585
R1208 B.n219 B.n218 585
R1209 B.n217 B.n216 585
R1210 B.n215 B.n214 585
R1211 B.n213 B.n212 585
R1212 B.n211 B.n210 585
R1213 B.n209 B.n208 585
R1214 B.n207 B.n206 585
R1215 B.n205 B.n204 585
R1216 B.n203 B.n202 585
R1217 B.n201 B.n200 585
R1218 B.n199 B.n198 585
R1219 B.n197 B.n196 585
R1220 B.n195 B.n194 585
R1221 B.n193 B.n192 585
R1222 B.n191 B.n190 585
R1223 B.n189 B.n188 585
R1224 B.n187 B.n186 585
R1225 B.n185 B.n184 585
R1226 B.n183 B.n182 585
R1227 B.n181 B.n180 585
R1228 B.n179 B.n178 585
R1229 B.n177 B.n176 585
R1230 B.n175 B.n174 585
R1231 B.n173 B.n172 585
R1232 B.n171 B.n170 585
R1233 B.n169 B.n168 585
R1234 B.n167 B.n166 585
R1235 B.n165 B.n164 585
R1236 B.n163 B.n162 585
R1237 B.n161 B.n160 585
R1238 B.n159 B.n158 585
R1239 B.n157 B.n156 585
R1240 B.n155 B.n154 585
R1241 B.n153 B.n152 585
R1242 B.n151 B.n150 585
R1243 B.n149 B.n148 585
R1244 B.n147 B.n146 585
R1245 B.n81 B.n80 585
R1246 B.n944 B.n943 585
R1247 B.n938 B.n140 585
R1248 B.n140 B.n78 585
R1249 B.n937 B.n77 585
R1250 B.n948 B.n77 585
R1251 B.n936 B.n76 585
R1252 B.n949 B.n76 585
R1253 B.n935 B.n75 585
R1254 B.n950 B.n75 585
R1255 B.n934 B.n933 585
R1256 B.n933 B.n71 585
R1257 B.n932 B.n70 585
R1258 B.n956 B.n70 585
R1259 B.n931 B.n69 585
R1260 B.n957 B.n69 585
R1261 B.n930 B.n68 585
R1262 B.n958 B.n68 585
R1263 B.n929 B.n928 585
R1264 B.n928 B.n64 585
R1265 B.n927 B.n63 585
R1266 B.n964 B.n63 585
R1267 B.n926 B.n62 585
R1268 B.n965 B.n62 585
R1269 B.n925 B.n61 585
R1270 B.n966 B.n61 585
R1271 B.n924 B.n923 585
R1272 B.n923 B.n57 585
R1273 B.n922 B.n56 585
R1274 B.n972 B.n56 585
R1275 B.n921 B.n55 585
R1276 B.n973 B.n55 585
R1277 B.n920 B.n54 585
R1278 B.n974 B.n54 585
R1279 B.n919 B.n918 585
R1280 B.n918 B.n50 585
R1281 B.n917 B.n49 585
R1282 B.n980 B.n49 585
R1283 B.n916 B.n48 585
R1284 B.n981 B.n48 585
R1285 B.n915 B.n47 585
R1286 B.n982 B.n47 585
R1287 B.n914 B.n913 585
R1288 B.n913 B.n43 585
R1289 B.n912 B.n42 585
R1290 B.n988 B.n42 585
R1291 B.n911 B.n41 585
R1292 B.n989 B.n41 585
R1293 B.n910 B.n40 585
R1294 B.n990 B.n40 585
R1295 B.n909 B.n908 585
R1296 B.n908 B.n39 585
R1297 B.n907 B.n35 585
R1298 B.n996 B.n35 585
R1299 B.n906 B.n34 585
R1300 B.n997 B.n34 585
R1301 B.n905 B.n33 585
R1302 B.n998 B.n33 585
R1303 B.n904 B.n903 585
R1304 B.n903 B.n29 585
R1305 B.n902 B.n28 585
R1306 B.n1004 B.n28 585
R1307 B.n901 B.n27 585
R1308 B.n1005 B.n27 585
R1309 B.n900 B.n26 585
R1310 B.n1006 B.n26 585
R1311 B.n899 B.n898 585
R1312 B.n898 B.n22 585
R1313 B.n897 B.n21 585
R1314 B.n1012 B.n21 585
R1315 B.n896 B.n20 585
R1316 B.n1013 B.n20 585
R1317 B.n895 B.n19 585
R1318 B.n1014 B.n19 585
R1319 B.n894 B.n893 585
R1320 B.n893 B.n15 585
R1321 B.n892 B.n14 585
R1322 B.n1020 B.n14 585
R1323 B.n891 B.n13 585
R1324 B.n1021 B.n13 585
R1325 B.n890 B.n12 585
R1326 B.n1022 B.n12 585
R1327 B.n889 B.n888 585
R1328 B.n888 B.n8 585
R1329 B.n887 B.n7 585
R1330 B.n1028 B.n7 585
R1331 B.n886 B.n6 585
R1332 B.n1029 B.n6 585
R1333 B.n885 B.n5 585
R1334 B.n1030 B.n5 585
R1335 B.n884 B.n883 585
R1336 B.n883 B.n4 585
R1337 B.n882 B.n374 585
R1338 B.n882 B.n881 585
R1339 B.n872 B.n375 585
R1340 B.n376 B.n375 585
R1341 B.n874 B.n873 585
R1342 B.n875 B.n874 585
R1343 B.n871 B.n381 585
R1344 B.n381 B.n380 585
R1345 B.n870 B.n869 585
R1346 B.n869 B.n868 585
R1347 B.n383 B.n382 585
R1348 B.n384 B.n383 585
R1349 B.n861 B.n860 585
R1350 B.n862 B.n861 585
R1351 B.n859 B.n389 585
R1352 B.n389 B.n388 585
R1353 B.n858 B.n857 585
R1354 B.n857 B.n856 585
R1355 B.n391 B.n390 585
R1356 B.n392 B.n391 585
R1357 B.n849 B.n848 585
R1358 B.n850 B.n849 585
R1359 B.n847 B.n397 585
R1360 B.n397 B.n396 585
R1361 B.n846 B.n845 585
R1362 B.n845 B.n844 585
R1363 B.n399 B.n398 585
R1364 B.n400 B.n399 585
R1365 B.n837 B.n836 585
R1366 B.n838 B.n837 585
R1367 B.n835 B.n405 585
R1368 B.n405 B.n404 585
R1369 B.n834 B.n833 585
R1370 B.n833 B.n832 585
R1371 B.n407 B.n406 585
R1372 B.n825 B.n407 585
R1373 B.n824 B.n823 585
R1374 B.n826 B.n824 585
R1375 B.n822 B.n412 585
R1376 B.n412 B.n411 585
R1377 B.n821 B.n820 585
R1378 B.n820 B.n819 585
R1379 B.n414 B.n413 585
R1380 B.n415 B.n414 585
R1381 B.n812 B.n811 585
R1382 B.n813 B.n812 585
R1383 B.n810 B.n420 585
R1384 B.n420 B.n419 585
R1385 B.n809 B.n808 585
R1386 B.n808 B.n807 585
R1387 B.n422 B.n421 585
R1388 B.n423 B.n422 585
R1389 B.n800 B.n799 585
R1390 B.n801 B.n800 585
R1391 B.n798 B.n428 585
R1392 B.n428 B.n427 585
R1393 B.n797 B.n796 585
R1394 B.n796 B.n795 585
R1395 B.n430 B.n429 585
R1396 B.n431 B.n430 585
R1397 B.n788 B.n787 585
R1398 B.n789 B.n788 585
R1399 B.n786 B.n436 585
R1400 B.n436 B.n435 585
R1401 B.n785 B.n784 585
R1402 B.n784 B.n783 585
R1403 B.n438 B.n437 585
R1404 B.n439 B.n438 585
R1405 B.n776 B.n775 585
R1406 B.n777 B.n776 585
R1407 B.n774 B.n444 585
R1408 B.n444 B.n443 585
R1409 B.n773 B.n772 585
R1410 B.n772 B.n771 585
R1411 B.n446 B.n445 585
R1412 B.n447 B.n446 585
R1413 B.n764 B.n763 585
R1414 B.n765 B.n764 585
R1415 B.n762 B.n452 585
R1416 B.n452 B.n451 585
R1417 B.n761 B.n760 585
R1418 B.n760 B.n759 585
R1419 B.n454 B.n453 585
R1420 B.n455 B.n454 585
R1421 B.n755 B.n754 585
R1422 B.n458 B.n457 585
R1423 B.n751 B.n750 585
R1424 B.n752 B.n751 585
R1425 B.n749 B.n516 585
R1426 B.n748 B.n747 585
R1427 B.n746 B.n745 585
R1428 B.n744 B.n743 585
R1429 B.n742 B.n741 585
R1430 B.n740 B.n739 585
R1431 B.n738 B.n737 585
R1432 B.n736 B.n735 585
R1433 B.n734 B.n733 585
R1434 B.n732 B.n731 585
R1435 B.n730 B.n729 585
R1436 B.n728 B.n727 585
R1437 B.n726 B.n725 585
R1438 B.n724 B.n723 585
R1439 B.n722 B.n721 585
R1440 B.n720 B.n719 585
R1441 B.n718 B.n717 585
R1442 B.n716 B.n715 585
R1443 B.n714 B.n713 585
R1444 B.n712 B.n711 585
R1445 B.n710 B.n709 585
R1446 B.n708 B.n707 585
R1447 B.n706 B.n705 585
R1448 B.n704 B.n703 585
R1449 B.n702 B.n701 585
R1450 B.n700 B.n699 585
R1451 B.n698 B.n697 585
R1452 B.n696 B.n695 585
R1453 B.n694 B.n693 585
R1454 B.n692 B.n691 585
R1455 B.n690 B.n689 585
R1456 B.n688 B.n687 585
R1457 B.n686 B.n685 585
R1458 B.n684 B.n683 585
R1459 B.n682 B.n681 585
R1460 B.n680 B.n679 585
R1461 B.n678 B.n677 585
R1462 B.n676 B.n675 585
R1463 B.n674 B.n673 585
R1464 B.n672 B.n671 585
R1465 B.n670 B.n669 585
R1466 B.n668 B.n667 585
R1467 B.n666 B.n665 585
R1468 B.n664 B.n663 585
R1469 B.n662 B.n661 585
R1470 B.n660 B.n659 585
R1471 B.n658 B.n657 585
R1472 B.n656 B.n655 585
R1473 B.n654 B.n653 585
R1474 B.n652 B.n651 585
R1475 B.n650 B.n649 585
R1476 B.n647 B.n646 585
R1477 B.n645 B.n644 585
R1478 B.n643 B.n642 585
R1479 B.n641 B.n640 585
R1480 B.n639 B.n638 585
R1481 B.n637 B.n636 585
R1482 B.n635 B.n634 585
R1483 B.n633 B.n632 585
R1484 B.n631 B.n630 585
R1485 B.n629 B.n628 585
R1486 B.n627 B.n626 585
R1487 B.n625 B.n624 585
R1488 B.n623 B.n622 585
R1489 B.n621 B.n620 585
R1490 B.n619 B.n618 585
R1491 B.n617 B.n616 585
R1492 B.n615 B.n614 585
R1493 B.n613 B.n612 585
R1494 B.n611 B.n610 585
R1495 B.n609 B.n608 585
R1496 B.n607 B.n606 585
R1497 B.n605 B.n604 585
R1498 B.n603 B.n602 585
R1499 B.n601 B.n600 585
R1500 B.n599 B.n598 585
R1501 B.n597 B.n596 585
R1502 B.n595 B.n594 585
R1503 B.n593 B.n592 585
R1504 B.n591 B.n590 585
R1505 B.n589 B.n588 585
R1506 B.n587 B.n586 585
R1507 B.n585 B.n584 585
R1508 B.n583 B.n582 585
R1509 B.n581 B.n580 585
R1510 B.n579 B.n578 585
R1511 B.n577 B.n576 585
R1512 B.n575 B.n574 585
R1513 B.n573 B.n572 585
R1514 B.n571 B.n570 585
R1515 B.n569 B.n568 585
R1516 B.n567 B.n566 585
R1517 B.n565 B.n564 585
R1518 B.n563 B.n562 585
R1519 B.n561 B.n560 585
R1520 B.n559 B.n558 585
R1521 B.n557 B.n556 585
R1522 B.n555 B.n554 585
R1523 B.n553 B.n552 585
R1524 B.n551 B.n550 585
R1525 B.n549 B.n548 585
R1526 B.n547 B.n546 585
R1527 B.n545 B.n544 585
R1528 B.n543 B.n542 585
R1529 B.n541 B.n540 585
R1530 B.n539 B.n538 585
R1531 B.n537 B.n536 585
R1532 B.n535 B.n534 585
R1533 B.n533 B.n532 585
R1534 B.n531 B.n530 585
R1535 B.n529 B.n528 585
R1536 B.n527 B.n526 585
R1537 B.n525 B.n524 585
R1538 B.n523 B.n522 585
R1539 B.n756 B.n456 585
R1540 B.n456 B.n455 585
R1541 B.n758 B.n757 585
R1542 B.n759 B.n758 585
R1543 B.n450 B.n449 585
R1544 B.n451 B.n450 585
R1545 B.n767 B.n766 585
R1546 B.n766 B.n765 585
R1547 B.n768 B.n448 585
R1548 B.n448 B.n447 585
R1549 B.n770 B.n769 585
R1550 B.n771 B.n770 585
R1551 B.n442 B.n441 585
R1552 B.n443 B.n442 585
R1553 B.n779 B.n778 585
R1554 B.n778 B.n777 585
R1555 B.n780 B.n440 585
R1556 B.n440 B.n439 585
R1557 B.n782 B.n781 585
R1558 B.n783 B.n782 585
R1559 B.n434 B.n433 585
R1560 B.n435 B.n434 585
R1561 B.n791 B.n790 585
R1562 B.n790 B.n789 585
R1563 B.n792 B.n432 585
R1564 B.n432 B.n431 585
R1565 B.n794 B.n793 585
R1566 B.n795 B.n794 585
R1567 B.n426 B.n425 585
R1568 B.n427 B.n426 585
R1569 B.n803 B.n802 585
R1570 B.n802 B.n801 585
R1571 B.n804 B.n424 585
R1572 B.n424 B.n423 585
R1573 B.n806 B.n805 585
R1574 B.n807 B.n806 585
R1575 B.n418 B.n417 585
R1576 B.n419 B.n418 585
R1577 B.n815 B.n814 585
R1578 B.n814 B.n813 585
R1579 B.n816 B.n416 585
R1580 B.n416 B.n415 585
R1581 B.n818 B.n817 585
R1582 B.n819 B.n818 585
R1583 B.n410 B.n409 585
R1584 B.n411 B.n410 585
R1585 B.n828 B.n827 585
R1586 B.n827 B.n826 585
R1587 B.n829 B.n408 585
R1588 B.n825 B.n408 585
R1589 B.n831 B.n830 585
R1590 B.n832 B.n831 585
R1591 B.n403 B.n402 585
R1592 B.n404 B.n403 585
R1593 B.n840 B.n839 585
R1594 B.n839 B.n838 585
R1595 B.n841 B.n401 585
R1596 B.n401 B.n400 585
R1597 B.n843 B.n842 585
R1598 B.n844 B.n843 585
R1599 B.n395 B.n394 585
R1600 B.n396 B.n395 585
R1601 B.n852 B.n851 585
R1602 B.n851 B.n850 585
R1603 B.n853 B.n393 585
R1604 B.n393 B.n392 585
R1605 B.n855 B.n854 585
R1606 B.n856 B.n855 585
R1607 B.n387 B.n386 585
R1608 B.n388 B.n387 585
R1609 B.n864 B.n863 585
R1610 B.n863 B.n862 585
R1611 B.n865 B.n385 585
R1612 B.n385 B.n384 585
R1613 B.n867 B.n866 585
R1614 B.n868 B.n867 585
R1615 B.n379 B.n378 585
R1616 B.n380 B.n379 585
R1617 B.n877 B.n876 585
R1618 B.n876 B.n875 585
R1619 B.n878 B.n377 585
R1620 B.n377 B.n376 585
R1621 B.n880 B.n879 585
R1622 B.n881 B.n880 585
R1623 B.n2 B.n0 585
R1624 B.n4 B.n2 585
R1625 B.n3 B.n1 585
R1626 B.n1029 B.n3 585
R1627 B.n1027 B.n1026 585
R1628 B.n1028 B.n1027 585
R1629 B.n1025 B.n9 585
R1630 B.n9 B.n8 585
R1631 B.n1024 B.n1023 585
R1632 B.n1023 B.n1022 585
R1633 B.n11 B.n10 585
R1634 B.n1021 B.n11 585
R1635 B.n1019 B.n1018 585
R1636 B.n1020 B.n1019 585
R1637 B.n1017 B.n16 585
R1638 B.n16 B.n15 585
R1639 B.n1016 B.n1015 585
R1640 B.n1015 B.n1014 585
R1641 B.n18 B.n17 585
R1642 B.n1013 B.n18 585
R1643 B.n1011 B.n1010 585
R1644 B.n1012 B.n1011 585
R1645 B.n1009 B.n23 585
R1646 B.n23 B.n22 585
R1647 B.n1008 B.n1007 585
R1648 B.n1007 B.n1006 585
R1649 B.n25 B.n24 585
R1650 B.n1005 B.n25 585
R1651 B.n1003 B.n1002 585
R1652 B.n1004 B.n1003 585
R1653 B.n1001 B.n30 585
R1654 B.n30 B.n29 585
R1655 B.n1000 B.n999 585
R1656 B.n999 B.n998 585
R1657 B.n32 B.n31 585
R1658 B.n997 B.n32 585
R1659 B.n995 B.n994 585
R1660 B.n996 B.n995 585
R1661 B.n993 B.n36 585
R1662 B.n39 B.n36 585
R1663 B.n992 B.n991 585
R1664 B.n991 B.n990 585
R1665 B.n38 B.n37 585
R1666 B.n989 B.n38 585
R1667 B.n987 B.n986 585
R1668 B.n988 B.n987 585
R1669 B.n985 B.n44 585
R1670 B.n44 B.n43 585
R1671 B.n984 B.n983 585
R1672 B.n983 B.n982 585
R1673 B.n46 B.n45 585
R1674 B.n981 B.n46 585
R1675 B.n979 B.n978 585
R1676 B.n980 B.n979 585
R1677 B.n977 B.n51 585
R1678 B.n51 B.n50 585
R1679 B.n976 B.n975 585
R1680 B.n975 B.n974 585
R1681 B.n53 B.n52 585
R1682 B.n973 B.n53 585
R1683 B.n971 B.n970 585
R1684 B.n972 B.n971 585
R1685 B.n969 B.n58 585
R1686 B.n58 B.n57 585
R1687 B.n968 B.n967 585
R1688 B.n967 B.n966 585
R1689 B.n60 B.n59 585
R1690 B.n965 B.n60 585
R1691 B.n963 B.n962 585
R1692 B.n964 B.n963 585
R1693 B.n961 B.n65 585
R1694 B.n65 B.n64 585
R1695 B.n960 B.n959 585
R1696 B.n959 B.n958 585
R1697 B.n67 B.n66 585
R1698 B.n957 B.n67 585
R1699 B.n955 B.n954 585
R1700 B.n956 B.n955 585
R1701 B.n953 B.n72 585
R1702 B.n72 B.n71 585
R1703 B.n952 B.n951 585
R1704 B.n951 B.n950 585
R1705 B.n74 B.n73 585
R1706 B.n949 B.n74 585
R1707 B.n947 B.n946 585
R1708 B.n948 B.n947 585
R1709 B.n945 B.n79 585
R1710 B.n79 B.n78 585
R1711 B.n1032 B.n1031 585
R1712 B.n1031 B.n1030 585
R1713 B.n754 B.n456 444.452
R1714 B.n943 B.n79 444.452
R1715 B.n522 B.n454 444.452
R1716 B.n940 B.n140 444.452
R1717 B.n519 B.t7 428.307
R1718 B.n141 B.t16 428.307
R1719 B.n517 B.t10 428.307
R1720 B.n143 B.t13 428.307
R1721 B.n520 B.t6 352.089
R1722 B.n142 B.t17 352.089
R1723 B.n518 B.t9 352.089
R1724 B.n144 B.t14 352.089
R1725 B.n519 B.t4 316.762
R1726 B.n517 B.t8 316.762
R1727 B.n143 B.t11 316.762
R1728 B.n141 B.t15 316.762
R1729 B.n941 B.n138 256.663
R1730 B.n941 B.n137 256.663
R1731 B.n941 B.n136 256.663
R1732 B.n941 B.n135 256.663
R1733 B.n941 B.n134 256.663
R1734 B.n941 B.n133 256.663
R1735 B.n941 B.n132 256.663
R1736 B.n941 B.n131 256.663
R1737 B.n941 B.n130 256.663
R1738 B.n941 B.n129 256.663
R1739 B.n941 B.n128 256.663
R1740 B.n941 B.n127 256.663
R1741 B.n941 B.n126 256.663
R1742 B.n941 B.n125 256.663
R1743 B.n941 B.n124 256.663
R1744 B.n941 B.n123 256.663
R1745 B.n941 B.n122 256.663
R1746 B.n941 B.n121 256.663
R1747 B.n941 B.n120 256.663
R1748 B.n941 B.n119 256.663
R1749 B.n941 B.n118 256.663
R1750 B.n941 B.n117 256.663
R1751 B.n941 B.n116 256.663
R1752 B.n941 B.n115 256.663
R1753 B.n941 B.n114 256.663
R1754 B.n941 B.n113 256.663
R1755 B.n941 B.n112 256.663
R1756 B.n941 B.n111 256.663
R1757 B.n941 B.n110 256.663
R1758 B.n941 B.n109 256.663
R1759 B.n941 B.n108 256.663
R1760 B.n941 B.n107 256.663
R1761 B.n941 B.n106 256.663
R1762 B.n941 B.n105 256.663
R1763 B.n941 B.n104 256.663
R1764 B.n941 B.n103 256.663
R1765 B.n941 B.n102 256.663
R1766 B.n941 B.n101 256.663
R1767 B.n941 B.n100 256.663
R1768 B.n941 B.n99 256.663
R1769 B.n941 B.n98 256.663
R1770 B.n941 B.n97 256.663
R1771 B.n941 B.n96 256.663
R1772 B.n941 B.n95 256.663
R1773 B.n941 B.n94 256.663
R1774 B.n941 B.n93 256.663
R1775 B.n941 B.n92 256.663
R1776 B.n941 B.n91 256.663
R1777 B.n941 B.n90 256.663
R1778 B.n941 B.n89 256.663
R1779 B.n941 B.n88 256.663
R1780 B.n941 B.n87 256.663
R1781 B.n941 B.n86 256.663
R1782 B.n941 B.n85 256.663
R1783 B.n941 B.n84 256.663
R1784 B.n941 B.n83 256.663
R1785 B.n941 B.n82 256.663
R1786 B.n942 B.n941 256.663
R1787 B.n753 B.n752 256.663
R1788 B.n752 B.n459 256.663
R1789 B.n752 B.n460 256.663
R1790 B.n752 B.n461 256.663
R1791 B.n752 B.n462 256.663
R1792 B.n752 B.n463 256.663
R1793 B.n752 B.n464 256.663
R1794 B.n752 B.n465 256.663
R1795 B.n752 B.n466 256.663
R1796 B.n752 B.n467 256.663
R1797 B.n752 B.n468 256.663
R1798 B.n752 B.n469 256.663
R1799 B.n752 B.n470 256.663
R1800 B.n752 B.n471 256.663
R1801 B.n752 B.n472 256.663
R1802 B.n752 B.n473 256.663
R1803 B.n752 B.n474 256.663
R1804 B.n752 B.n475 256.663
R1805 B.n752 B.n476 256.663
R1806 B.n752 B.n477 256.663
R1807 B.n752 B.n478 256.663
R1808 B.n752 B.n479 256.663
R1809 B.n752 B.n480 256.663
R1810 B.n752 B.n481 256.663
R1811 B.n752 B.n482 256.663
R1812 B.n752 B.n483 256.663
R1813 B.n752 B.n484 256.663
R1814 B.n752 B.n485 256.663
R1815 B.n752 B.n486 256.663
R1816 B.n752 B.n487 256.663
R1817 B.n752 B.n488 256.663
R1818 B.n752 B.n489 256.663
R1819 B.n752 B.n490 256.663
R1820 B.n752 B.n491 256.663
R1821 B.n752 B.n492 256.663
R1822 B.n752 B.n493 256.663
R1823 B.n752 B.n494 256.663
R1824 B.n752 B.n495 256.663
R1825 B.n752 B.n496 256.663
R1826 B.n752 B.n497 256.663
R1827 B.n752 B.n498 256.663
R1828 B.n752 B.n499 256.663
R1829 B.n752 B.n500 256.663
R1830 B.n752 B.n501 256.663
R1831 B.n752 B.n502 256.663
R1832 B.n752 B.n503 256.663
R1833 B.n752 B.n504 256.663
R1834 B.n752 B.n505 256.663
R1835 B.n752 B.n506 256.663
R1836 B.n752 B.n507 256.663
R1837 B.n752 B.n508 256.663
R1838 B.n752 B.n509 256.663
R1839 B.n752 B.n510 256.663
R1840 B.n752 B.n511 256.663
R1841 B.n752 B.n512 256.663
R1842 B.n752 B.n513 256.663
R1843 B.n752 B.n514 256.663
R1844 B.n752 B.n515 256.663
R1845 B.n758 B.n456 163.367
R1846 B.n758 B.n450 163.367
R1847 B.n766 B.n450 163.367
R1848 B.n766 B.n448 163.367
R1849 B.n770 B.n448 163.367
R1850 B.n770 B.n442 163.367
R1851 B.n778 B.n442 163.367
R1852 B.n778 B.n440 163.367
R1853 B.n782 B.n440 163.367
R1854 B.n782 B.n434 163.367
R1855 B.n790 B.n434 163.367
R1856 B.n790 B.n432 163.367
R1857 B.n794 B.n432 163.367
R1858 B.n794 B.n426 163.367
R1859 B.n802 B.n426 163.367
R1860 B.n802 B.n424 163.367
R1861 B.n806 B.n424 163.367
R1862 B.n806 B.n418 163.367
R1863 B.n814 B.n418 163.367
R1864 B.n814 B.n416 163.367
R1865 B.n818 B.n416 163.367
R1866 B.n818 B.n410 163.367
R1867 B.n827 B.n410 163.367
R1868 B.n827 B.n408 163.367
R1869 B.n831 B.n408 163.367
R1870 B.n831 B.n403 163.367
R1871 B.n839 B.n403 163.367
R1872 B.n839 B.n401 163.367
R1873 B.n843 B.n401 163.367
R1874 B.n843 B.n395 163.367
R1875 B.n851 B.n395 163.367
R1876 B.n851 B.n393 163.367
R1877 B.n855 B.n393 163.367
R1878 B.n855 B.n387 163.367
R1879 B.n863 B.n387 163.367
R1880 B.n863 B.n385 163.367
R1881 B.n867 B.n385 163.367
R1882 B.n867 B.n379 163.367
R1883 B.n876 B.n379 163.367
R1884 B.n876 B.n377 163.367
R1885 B.n880 B.n377 163.367
R1886 B.n880 B.n2 163.367
R1887 B.n1031 B.n2 163.367
R1888 B.n1031 B.n3 163.367
R1889 B.n1027 B.n3 163.367
R1890 B.n1027 B.n9 163.367
R1891 B.n1023 B.n9 163.367
R1892 B.n1023 B.n11 163.367
R1893 B.n1019 B.n11 163.367
R1894 B.n1019 B.n16 163.367
R1895 B.n1015 B.n16 163.367
R1896 B.n1015 B.n18 163.367
R1897 B.n1011 B.n18 163.367
R1898 B.n1011 B.n23 163.367
R1899 B.n1007 B.n23 163.367
R1900 B.n1007 B.n25 163.367
R1901 B.n1003 B.n25 163.367
R1902 B.n1003 B.n30 163.367
R1903 B.n999 B.n30 163.367
R1904 B.n999 B.n32 163.367
R1905 B.n995 B.n32 163.367
R1906 B.n995 B.n36 163.367
R1907 B.n991 B.n36 163.367
R1908 B.n991 B.n38 163.367
R1909 B.n987 B.n38 163.367
R1910 B.n987 B.n44 163.367
R1911 B.n983 B.n44 163.367
R1912 B.n983 B.n46 163.367
R1913 B.n979 B.n46 163.367
R1914 B.n979 B.n51 163.367
R1915 B.n975 B.n51 163.367
R1916 B.n975 B.n53 163.367
R1917 B.n971 B.n53 163.367
R1918 B.n971 B.n58 163.367
R1919 B.n967 B.n58 163.367
R1920 B.n967 B.n60 163.367
R1921 B.n963 B.n60 163.367
R1922 B.n963 B.n65 163.367
R1923 B.n959 B.n65 163.367
R1924 B.n959 B.n67 163.367
R1925 B.n955 B.n67 163.367
R1926 B.n955 B.n72 163.367
R1927 B.n951 B.n72 163.367
R1928 B.n951 B.n74 163.367
R1929 B.n947 B.n74 163.367
R1930 B.n947 B.n79 163.367
R1931 B.n751 B.n458 163.367
R1932 B.n751 B.n516 163.367
R1933 B.n747 B.n746 163.367
R1934 B.n743 B.n742 163.367
R1935 B.n739 B.n738 163.367
R1936 B.n735 B.n734 163.367
R1937 B.n731 B.n730 163.367
R1938 B.n727 B.n726 163.367
R1939 B.n723 B.n722 163.367
R1940 B.n719 B.n718 163.367
R1941 B.n715 B.n714 163.367
R1942 B.n711 B.n710 163.367
R1943 B.n707 B.n706 163.367
R1944 B.n703 B.n702 163.367
R1945 B.n699 B.n698 163.367
R1946 B.n695 B.n694 163.367
R1947 B.n691 B.n690 163.367
R1948 B.n687 B.n686 163.367
R1949 B.n683 B.n682 163.367
R1950 B.n679 B.n678 163.367
R1951 B.n675 B.n674 163.367
R1952 B.n671 B.n670 163.367
R1953 B.n667 B.n666 163.367
R1954 B.n663 B.n662 163.367
R1955 B.n659 B.n658 163.367
R1956 B.n655 B.n654 163.367
R1957 B.n651 B.n650 163.367
R1958 B.n646 B.n645 163.367
R1959 B.n642 B.n641 163.367
R1960 B.n638 B.n637 163.367
R1961 B.n634 B.n633 163.367
R1962 B.n630 B.n629 163.367
R1963 B.n626 B.n625 163.367
R1964 B.n622 B.n621 163.367
R1965 B.n618 B.n617 163.367
R1966 B.n614 B.n613 163.367
R1967 B.n610 B.n609 163.367
R1968 B.n606 B.n605 163.367
R1969 B.n602 B.n601 163.367
R1970 B.n598 B.n597 163.367
R1971 B.n594 B.n593 163.367
R1972 B.n590 B.n589 163.367
R1973 B.n586 B.n585 163.367
R1974 B.n582 B.n581 163.367
R1975 B.n578 B.n577 163.367
R1976 B.n574 B.n573 163.367
R1977 B.n570 B.n569 163.367
R1978 B.n566 B.n565 163.367
R1979 B.n562 B.n561 163.367
R1980 B.n558 B.n557 163.367
R1981 B.n554 B.n553 163.367
R1982 B.n550 B.n549 163.367
R1983 B.n546 B.n545 163.367
R1984 B.n542 B.n541 163.367
R1985 B.n538 B.n537 163.367
R1986 B.n534 B.n533 163.367
R1987 B.n530 B.n529 163.367
R1988 B.n526 B.n525 163.367
R1989 B.n760 B.n454 163.367
R1990 B.n760 B.n452 163.367
R1991 B.n764 B.n452 163.367
R1992 B.n764 B.n446 163.367
R1993 B.n772 B.n446 163.367
R1994 B.n772 B.n444 163.367
R1995 B.n776 B.n444 163.367
R1996 B.n776 B.n438 163.367
R1997 B.n784 B.n438 163.367
R1998 B.n784 B.n436 163.367
R1999 B.n788 B.n436 163.367
R2000 B.n788 B.n430 163.367
R2001 B.n796 B.n430 163.367
R2002 B.n796 B.n428 163.367
R2003 B.n800 B.n428 163.367
R2004 B.n800 B.n422 163.367
R2005 B.n808 B.n422 163.367
R2006 B.n808 B.n420 163.367
R2007 B.n812 B.n420 163.367
R2008 B.n812 B.n414 163.367
R2009 B.n820 B.n414 163.367
R2010 B.n820 B.n412 163.367
R2011 B.n824 B.n412 163.367
R2012 B.n824 B.n407 163.367
R2013 B.n833 B.n407 163.367
R2014 B.n833 B.n405 163.367
R2015 B.n837 B.n405 163.367
R2016 B.n837 B.n399 163.367
R2017 B.n845 B.n399 163.367
R2018 B.n845 B.n397 163.367
R2019 B.n849 B.n397 163.367
R2020 B.n849 B.n391 163.367
R2021 B.n857 B.n391 163.367
R2022 B.n857 B.n389 163.367
R2023 B.n861 B.n389 163.367
R2024 B.n861 B.n383 163.367
R2025 B.n869 B.n383 163.367
R2026 B.n869 B.n381 163.367
R2027 B.n874 B.n381 163.367
R2028 B.n874 B.n375 163.367
R2029 B.n882 B.n375 163.367
R2030 B.n883 B.n882 163.367
R2031 B.n883 B.n5 163.367
R2032 B.n6 B.n5 163.367
R2033 B.n7 B.n6 163.367
R2034 B.n888 B.n7 163.367
R2035 B.n888 B.n12 163.367
R2036 B.n13 B.n12 163.367
R2037 B.n14 B.n13 163.367
R2038 B.n893 B.n14 163.367
R2039 B.n893 B.n19 163.367
R2040 B.n20 B.n19 163.367
R2041 B.n21 B.n20 163.367
R2042 B.n898 B.n21 163.367
R2043 B.n898 B.n26 163.367
R2044 B.n27 B.n26 163.367
R2045 B.n28 B.n27 163.367
R2046 B.n903 B.n28 163.367
R2047 B.n903 B.n33 163.367
R2048 B.n34 B.n33 163.367
R2049 B.n35 B.n34 163.367
R2050 B.n908 B.n35 163.367
R2051 B.n908 B.n40 163.367
R2052 B.n41 B.n40 163.367
R2053 B.n42 B.n41 163.367
R2054 B.n913 B.n42 163.367
R2055 B.n913 B.n47 163.367
R2056 B.n48 B.n47 163.367
R2057 B.n49 B.n48 163.367
R2058 B.n918 B.n49 163.367
R2059 B.n918 B.n54 163.367
R2060 B.n55 B.n54 163.367
R2061 B.n56 B.n55 163.367
R2062 B.n923 B.n56 163.367
R2063 B.n923 B.n61 163.367
R2064 B.n62 B.n61 163.367
R2065 B.n63 B.n62 163.367
R2066 B.n928 B.n63 163.367
R2067 B.n928 B.n68 163.367
R2068 B.n69 B.n68 163.367
R2069 B.n70 B.n69 163.367
R2070 B.n933 B.n70 163.367
R2071 B.n933 B.n75 163.367
R2072 B.n76 B.n75 163.367
R2073 B.n77 B.n76 163.367
R2074 B.n140 B.n77 163.367
R2075 B.n146 B.n81 163.367
R2076 B.n150 B.n149 163.367
R2077 B.n154 B.n153 163.367
R2078 B.n158 B.n157 163.367
R2079 B.n162 B.n161 163.367
R2080 B.n166 B.n165 163.367
R2081 B.n170 B.n169 163.367
R2082 B.n174 B.n173 163.367
R2083 B.n178 B.n177 163.367
R2084 B.n182 B.n181 163.367
R2085 B.n186 B.n185 163.367
R2086 B.n190 B.n189 163.367
R2087 B.n194 B.n193 163.367
R2088 B.n198 B.n197 163.367
R2089 B.n202 B.n201 163.367
R2090 B.n206 B.n205 163.367
R2091 B.n210 B.n209 163.367
R2092 B.n214 B.n213 163.367
R2093 B.n218 B.n217 163.367
R2094 B.n222 B.n221 163.367
R2095 B.n226 B.n225 163.367
R2096 B.n230 B.n229 163.367
R2097 B.n234 B.n233 163.367
R2098 B.n238 B.n237 163.367
R2099 B.n242 B.n241 163.367
R2100 B.n246 B.n245 163.367
R2101 B.n250 B.n249 163.367
R2102 B.n254 B.n253 163.367
R2103 B.n258 B.n257 163.367
R2104 B.n262 B.n261 163.367
R2105 B.n266 B.n265 163.367
R2106 B.n271 B.n270 163.367
R2107 B.n275 B.n274 163.367
R2108 B.n279 B.n278 163.367
R2109 B.n283 B.n282 163.367
R2110 B.n287 B.n286 163.367
R2111 B.n291 B.n290 163.367
R2112 B.n295 B.n294 163.367
R2113 B.n299 B.n298 163.367
R2114 B.n303 B.n302 163.367
R2115 B.n307 B.n306 163.367
R2116 B.n311 B.n310 163.367
R2117 B.n315 B.n314 163.367
R2118 B.n319 B.n318 163.367
R2119 B.n323 B.n322 163.367
R2120 B.n327 B.n326 163.367
R2121 B.n331 B.n330 163.367
R2122 B.n335 B.n334 163.367
R2123 B.n339 B.n338 163.367
R2124 B.n343 B.n342 163.367
R2125 B.n347 B.n346 163.367
R2126 B.n351 B.n350 163.367
R2127 B.n355 B.n354 163.367
R2128 B.n359 B.n358 163.367
R2129 B.n363 B.n362 163.367
R2130 B.n367 B.n366 163.367
R2131 B.n371 B.n370 163.367
R2132 B.n940 B.n139 163.367
R2133 B.n520 B.n519 76.2187
R2134 B.n518 B.n517 76.2187
R2135 B.n144 B.n143 76.2187
R2136 B.n142 B.n141 76.2187
R2137 B.n754 B.n753 71.676
R2138 B.n516 B.n459 71.676
R2139 B.n746 B.n460 71.676
R2140 B.n742 B.n461 71.676
R2141 B.n738 B.n462 71.676
R2142 B.n734 B.n463 71.676
R2143 B.n730 B.n464 71.676
R2144 B.n726 B.n465 71.676
R2145 B.n722 B.n466 71.676
R2146 B.n718 B.n467 71.676
R2147 B.n714 B.n468 71.676
R2148 B.n710 B.n469 71.676
R2149 B.n706 B.n470 71.676
R2150 B.n702 B.n471 71.676
R2151 B.n698 B.n472 71.676
R2152 B.n694 B.n473 71.676
R2153 B.n690 B.n474 71.676
R2154 B.n686 B.n475 71.676
R2155 B.n682 B.n476 71.676
R2156 B.n678 B.n477 71.676
R2157 B.n674 B.n478 71.676
R2158 B.n670 B.n479 71.676
R2159 B.n666 B.n480 71.676
R2160 B.n662 B.n481 71.676
R2161 B.n658 B.n482 71.676
R2162 B.n654 B.n483 71.676
R2163 B.n650 B.n484 71.676
R2164 B.n645 B.n485 71.676
R2165 B.n641 B.n486 71.676
R2166 B.n637 B.n487 71.676
R2167 B.n633 B.n488 71.676
R2168 B.n629 B.n489 71.676
R2169 B.n625 B.n490 71.676
R2170 B.n621 B.n491 71.676
R2171 B.n617 B.n492 71.676
R2172 B.n613 B.n493 71.676
R2173 B.n609 B.n494 71.676
R2174 B.n605 B.n495 71.676
R2175 B.n601 B.n496 71.676
R2176 B.n597 B.n497 71.676
R2177 B.n593 B.n498 71.676
R2178 B.n589 B.n499 71.676
R2179 B.n585 B.n500 71.676
R2180 B.n581 B.n501 71.676
R2181 B.n577 B.n502 71.676
R2182 B.n573 B.n503 71.676
R2183 B.n569 B.n504 71.676
R2184 B.n565 B.n505 71.676
R2185 B.n561 B.n506 71.676
R2186 B.n557 B.n507 71.676
R2187 B.n553 B.n508 71.676
R2188 B.n549 B.n509 71.676
R2189 B.n545 B.n510 71.676
R2190 B.n541 B.n511 71.676
R2191 B.n537 B.n512 71.676
R2192 B.n533 B.n513 71.676
R2193 B.n529 B.n514 71.676
R2194 B.n525 B.n515 71.676
R2195 B.n943 B.n942 71.676
R2196 B.n146 B.n82 71.676
R2197 B.n150 B.n83 71.676
R2198 B.n154 B.n84 71.676
R2199 B.n158 B.n85 71.676
R2200 B.n162 B.n86 71.676
R2201 B.n166 B.n87 71.676
R2202 B.n170 B.n88 71.676
R2203 B.n174 B.n89 71.676
R2204 B.n178 B.n90 71.676
R2205 B.n182 B.n91 71.676
R2206 B.n186 B.n92 71.676
R2207 B.n190 B.n93 71.676
R2208 B.n194 B.n94 71.676
R2209 B.n198 B.n95 71.676
R2210 B.n202 B.n96 71.676
R2211 B.n206 B.n97 71.676
R2212 B.n210 B.n98 71.676
R2213 B.n214 B.n99 71.676
R2214 B.n218 B.n100 71.676
R2215 B.n222 B.n101 71.676
R2216 B.n226 B.n102 71.676
R2217 B.n230 B.n103 71.676
R2218 B.n234 B.n104 71.676
R2219 B.n238 B.n105 71.676
R2220 B.n242 B.n106 71.676
R2221 B.n246 B.n107 71.676
R2222 B.n250 B.n108 71.676
R2223 B.n254 B.n109 71.676
R2224 B.n258 B.n110 71.676
R2225 B.n262 B.n111 71.676
R2226 B.n266 B.n112 71.676
R2227 B.n271 B.n113 71.676
R2228 B.n275 B.n114 71.676
R2229 B.n279 B.n115 71.676
R2230 B.n283 B.n116 71.676
R2231 B.n287 B.n117 71.676
R2232 B.n291 B.n118 71.676
R2233 B.n295 B.n119 71.676
R2234 B.n299 B.n120 71.676
R2235 B.n303 B.n121 71.676
R2236 B.n307 B.n122 71.676
R2237 B.n311 B.n123 71.676
R2238 B.n315 B.n124 71.676
R2239 B.n319 B.n125 71.676
R2240 B.n323 B.n126 71.676
R2241 B.n327 B.n127 71.676
R2242 B.n331 B.n128 71.676
R2243 B.n335 B.n129 71.676
R2244 B.n339 B.n130 71.676
R2245 B.n343 B.n131 71.676
R2246 B.n347 B.n132 71.676
R2247 B.n351 B.n133 71.676
R2248 B.n355 B.n134 71.676
R2249 B.n359 B.n135 71.676
R2250 B.n363 B.n136 71.676
R2251 B.n367 B.n137 71.676
R2252 B.n371 B.n138 71.676
R2253 B.n139 B.n138 71.676
R2254 B.n370 B.n137 71.676
R2255 B.n366 B.n136 71.676
R2256 B.n362 B.n135 71.676
R2257 B.n358 B.n134 71.676
R2258 B.n354 B.n133 71.676
R2259 B.n350 B.n132 71.676
R2260 B.n346 B.n131 71.676
R2261 B.n342 B.n130 71.676
R2262 B.n338 B.n129 71.676
R2263 B.n334 B.n128 71.676
R2264 B.n330 B.n127 71.676
R2265 B.n326 B.n126 71.676
R2266 B.n322 B.n125 71.676
R2267 B.n318 B.n124 71.676
R2268 B.n314 B.n123 71.676
R2269 B.n310 B.n122 71.676
R2270 B.n306 B.n121 71.676
R2271 B.n302 B.n120 71.676
R2272 B.n298 B.n119 71.676
R2273 B.n294 B.n118 71.676
R2274 B.n290 B.n117 71.676
R2275 B.n286 B.n116 71.676
R2276 B.n282 B.n115 71.676
R2277 B.n278 B.n114 71.676
R2278 B.n274 B.n113 71.676
R2279 B.n270 B.n112 71.676
R2280 B.n265 B.n111 71.676
R2281 B.n261 B.n110 71.676
R2282 B.n257 B.n109 71.676
R2283 B.n253 B.n108 71.676
R2284 B.n249 B.n107 71.676
R2285 B.n245 B.n106 71.676
R2286 B.n241 B.n105 71.676
R2287 B.n237 B.n104 71.676
R2288 B.n233 B.n103 71.676
R2289 B.n229 B.n102 71.676
R2290 B.n225 B.n101 71.676
R2291 B.n221 B.n100 71.676
R2292 B.n217 B.n99 71.676
R2293 B.n213 B.n98 71.676
R2294 B.n209 B.n97 71.676
R2295 B.n205 B.n96 71.676
R2296 B.n201 B.n95 71.676
R2297 B.n197 B.n94 71.676
R2298 B.n193 B.n93 71.676
R2299 B.n189 B.n92 71.676
R2300 B.n185 B.n91 71.676
R2301 B.n181 B.n90 71.676
R2302 B.n177 B.n89 71.676
R2303 B.n173 B.n88 71.676
R2304 B.n169 B.n87 71.676
R2305 B.n165 B.n86 71.676
R2306 B.n161 B.n85 71.676
R2307 B.n157 B.n84 71.676
R2308 B.n153 B.n83 71.676
R2309 B.n149 B.n82 71.676
R2310 B.n942 B.n81 71.676
R2311 B.n753 B.n458 71.676
R2312 B.n747 B.n459 71.676
R2313 B.n743 B.n460 71.676
R2314 B.n739 B.n461 71.676
R2315 B.n735 B.n462 71.676
R2316 B.n731 B.n463 71.676
R2317 B.n727 B.n464 71.676
R2318 B.n723 B.n465 71.676
R2319 B.n719 B.n466 71.676
R2320 B.n715 B.n467 71.676
R2321 B.n711 B.n468 71.676
R2322 B.n707 B.n469 71.676
R2323 B.n703 B.n470 71.676
R2324 B.n699 B.n471 71.676
R2325 B.n695 B.n472 71.676
R2326 B.n691 B.n473 71.676
R2327 B.n687 B.n474 71.676
R2328 B.n683 B.n475 71.676
R2329 B.n679 B.n476 71.676
R2330 B.n675 B.n477 71.676
R2331 B.n671 B.n478 71.676
R2332 B.n667 B.n479 71.676
R2333 B.n663 B.n480 71.676
R2334 B.n659 B.n481 71.676
R2335 B.n655 B.n482 71.676
R2336 B.n651 B.n483 71.676
R2337 B.n646 B.n484 71.676
R2338 B.n642 B.n485 71.676
R2339 B.n638 B.n486 71.676
R2340 B.n634 B.n487 71.676
R2341 B.n630 B.n488 71.676
R2342 B.n626 B.n489 71.676
R2343 B.n622 B.n490 71.676
R2344 B.n618 B.n491 71.676
R2345 B.n614 B.n492 71.676
R2346 B.n610 B.n493 71.676
R2347 B.n606 B.n494 71.676
R2348 B.n602 B.n495 71.676
R2349 B.n598 B.n496 71.676
R2350 B.n594 B.n497 71.676
R2351 B.n590 B.n498 71.676
R2352 B.n586 B.n499 71.676
R2353 B.n582 B.n500 71.676
R2354 B.n578 B.n501 71.676
R2355 B.n574 B.n502 71.676
R2356 B.n570 B.n503 71.676
R2357 B.n566 B.n504 71.676
R2358 B.n562 B.n505 71.676
R2359 B.n558 B.n506 71.676
R2360 B.n554 B.n507 71.676
R2361 B.n550 B.n508 71.676
R2362 B.n546 B.n509 71.676
R2363 B.n542 B.n510 71.676
R2364 B.n538 B.n511 71.676
R2365 B.n534 B.n512 71.676
R2366 B.n530 B.n513 71.676
R2367 B.n526 B.n514 71.676
R2368 B.n522 B.n515 71.676
R2369 B.n521 B.n520 59.5399
R2370 B.n648 B.n518 59.5399
R2371 B.n145 B.n144 59.5399
R2372 B.n268 B.n142 59.5399
R2373 B.n752 B.n455 56.1729
R2374 B.n941 B.n78 56.1729
R2375 B.n759 B.n455 35.0438
R2376 B.n759 B.n451 35.0438
R2377 B.n765 B.n451 35.0438
R2378 B.n765 B.n447 35.0438
R2379 B.n771 B.n447 35.0438
R2380 B.n771 B.n443 35.0438
R2381 B.n777 B.n443 35.0438
R2382 B.n777 B.n439 35.0438
R2383 B.n783 B.n439 35.0438
R2384 B.n789 B.n435 35.0438
R2385 B.n789 B.n431 35.0438
R2386 B.n795 B.n431 35.0438
R2387 B.n795 B.n427 35.0438
R2388 B.n801 B.n427 35.0438
R2389 B.n801 B.n423 35.0438
R2390 B.n807 B.n423 35.0438
R2391 B.n807 B.n419 35.0438
R2392 B.n813 B.n419 35.0438
R2393 B.n813 B.n415 35.0438
R2394 B.n819 B.n415 35.0438
R2395 B.n819 B.n411 35.0438
R2396 B.n826 B.n411 35.0438
R2397 B.n826 B.n825 35.0438
R2398 B.n832 B.n404 35.0438
R2399 B.n838 B.n404 35.0438
R2400 B.n838 B.n400 35.0438
R2401 B.n844 B.n400 35.0438
R2402 B.n844 B.n396 35.0438
R2403 B.n850 B.n396 35.0438
R2404 B.n850 B.n392 35.0438
R2405 B.n856 B.n392 35.0438
R2406 B.n856 B.n388 35.0438
R2407 B.n862 B.n388 35.0438
R2408 B.n868 B.n384 35.0438
R2409 B.n868 B.n380 35.0438
R2410 B.n875 B.n380 35.0438
R2411 B.n875 B.n376 35.0438
R2412 B.n881 B.n376 35.0438
R2413 B.n881 B.n4 35.0438
R2414 B.n1030 B.n4 35.0438
R2415 B.n1030 B.n1029 35.0438
R2416 B.n1029 B.n1028 35.0438
R2417 B.n1028 B.n8 35.0438
R2418 B.n1022 B.n8 35.0438
R2419 B.n1022 B.n1021 35.0438
R2420 B.n1021 B.n1020 35.0438
R2421 B.n1020 B.n15 35.0438
R2422 B.n1014 B.n1013 35.0438
R2423 B.n1013 B.n1012 35.0438
R2424 B.n1012 B.n22 35.0438
R2425 B.n1006 B.n22 35.0438
R2426 B.n1006 B.n1005 35.0438
R2427 B.n1005 B.n1004 35.0438
R2428 B.n1004 B.n29 35.0438
R2429 B.n998 B.n29 35.0438
R2430 B.n998 B.n997 35.0438
R2431 B.n997 B.n996 35.0438
R2432 B.n990 B.n39 35.0438
R2433 B.n990 B.n989 35.0438
R2434 B.n989 B.n988 35.0438
R2435 B.n988 B.n43 35.0438
R2436 B.n982 B.n43 35.0438
R2437 B.n982 B.n981 35.0438
R2438 B.n981 B.n980 35.0438
R2439 B.n980 B.n50 35.0438
R2440 B.n974 B.n50 35.0438
R2441 B.n974 B.n973 35.0438
R2442 B.n973 B.n972 35.0438
R2443 B.n972 B.n57 35.0438
R2444 B.n966 B.n57 35.0438
R2445 B.n966 B.n965 35.0438
R2446 B.n964 B.n64 35.0438
R2447 B.n958 B.n64 35.0438
R2448 B.n958 B.n957 35.0438
R2449 B.n957 B.n956 35.0438
R2450 B.n956 B.n71 35.0438
R2451 B.n950 B.n71 35.0438
R2452 B.n950 B.n949 35.0438
R2453 B.n949 B.n948 35.0438
R2454 B.n948 B.n78 35.0438
R2455 B.n832 B.t2 32.9825
R2456 B.n996 B.t3 32.9825
R2457 B.n945 B.n944 28.8785
R2458 B.n523 B.n453 28.8785
R2459 B.n756 B.n755 28.8785
R2460 B.n939 B.n938 28.8785
R2461 B.t5 B.n435 24.737
R2462 B.n965 B.t12 24.737
R2463 B.n862 B.t0 21.6449
R2464 B.n1014 B.t1 21.6449
R2465 B B.n1032 18.0485
R2466 B.t0 B.n384 13.3994
R2467 B.t1 B.n15 13.3994
R2468 B.n944 B.n80 10.6151
R2469 B.n147 B.n80 10.6151
R2470 B.n148 B.n147 10.6151
R2471 B.n151 B.n148 10.6151
R2472 B.n152 B.n151 10.6151
R2473 B.n155 B.n152 10.6151
R2474 B.n156 B.n155 10.6151
R2475 B.n159 B.n156 10.6151
R2476 B.n160 B.n159 10.6151
R2477 B.n163 B.n160 10.6151
R2478 B.n164 B.n163 10.6151
R2479 B.n167 B.n164 10.6151
R2480 B.n168 B.n167 10.6151
R2481 B.n171 B.n168 10.6151
R2482 B.n172 B.n171 10.6151
R2483 B.n175 B.n172 10.6151
R2484 B.n176 B.n175 10.6151
R2485 B.n179 B.n176 10.6151
R2486 B.n180 B.n179 10.6151
R2487 B.n183 B.n180 10.6151
R2488 B.n184 B.n183 10.6151
R2489 B.n187 B.n184 10.6151
R2490 B.n188 B.n187 10.6151
R2491 B.n191 B.n188 10.6151
R2492 B.n192 B.n191 10.6151
R2493 B.n195 B.n192 10.6151
R2494 B.n196 B.n195 10.6151
R2495 B.n199 B.n196 10.6151
R2496 B.n200 B.n199 10.6151
R2497 B.n203 B.n200 10.6151
R2498 B.n204 B.n203 10.6151
R2499 B.n207 B.n204 10.6151
R2500 B.n208 B.n207 10.6151
R2501 B.n211 B.n208 10.6151
R2502 B.n212 B.n211 10.6151
R2503 B.n215 B.n212 10.6151
R2504 B.n216 B.n215 10.6151
R2505 B.n219 B.n216 10.6151
R2506 B.n220 B.n219 10.6151
R2507 B.n223 B.n220 10.6151
R2508 B.n224 B.n223 10.6151
R2509 B.n227 B.n224 10.6151
R2510 B.n228 B.n227 10.6151
R2511 B.n231 B.n228 10.6151
R2512 B.n232 B.n231 10.6151
R2513 B.n235 B.n232 10.6151
R2514 B.n236 B.n235 10.6151
R2515 B.n239 B.n236 10.6151
R2516 B.n240 B.n239 10.6151
R2517 B.n243 B.n240 10.6151
R2518 B.n244 B.n243 10.6151
R2519 B.n247 B.n244 10.6151
R2520 B.n248 B.n247 10.6151
R2521 B.n252 B.n251 10.6151
R2522 B.n255 B.n252 10.6151
R2523 B.n256 B.n255 10.6151
R2524 B.n259 B.n256 10.6151
R2525 B.n260 B.n259 10.6151
R2526 B.n263 B.n260 10.6151
R2527 B.n264 B.n263 10.6151
R2528 B.n267 B.n264 10.6151
R2529 B.n272 B.n269 10.6151
R2530 B.n273 B.n272 10.6151
R2531 B.n276 B.n273 10.6151
R2532 B.n277 B.n276 10.6151
R2533 B.n280 B.n277 10.6151
R2534 B.n281 B.n280 10.6151
R2535 B.n284 B.n281 10.6151
R2536 B.n285 B.n284 10.6151
R2537 B.n288 B.n285 10.6151
R2538 B.n289 B.n288 10.6151
R2539 B.n292 B.n289 10.6151
R2540 B.n293 B.n292 10.6151
R2541 B.n296 B.n293 10.6151
R2542 B.n297 B.n296 10.6151
R2543 B.n300 B.n297 10.6151
R2544 B.n301 B.n300 10.6151
R2545 B.n304 B.n301 10.6151
R2546 B.n305 B.n304 10.6151
R2547 B.n308 B.n305 10.6151
R2548 B.n309 B.n308 10.6151
R2549 B.n312 B.n309 10.6151
R2550 B.n313 B.n312 10.6151
R2551 B.n316 B.n313 10.6151
R2552 B.n317 B.n316 10.6151
R2553 B.n320 B.n317 10.6151
R2554 B.n321 B.n320 10.6151
R2555 B.n324 B.n321 10.6151
R2556 B.n325 B.n324 10.6151
R2557 B.n328 B.n325 10.6151
R2558 B.n329 B.n328 10.6151
R2559 B.n332 B.n329 10.6151
R2560 B.n333 B.n332 10.6151
R2561 B.n336 B.n333 10.6151
R2562 B.n337 B.n336 10.6151
R2563 B.n340 B.n337 10.6151
R2564 B.n341 B.n340 10.6151
R2565 B.n344 B.n341 10.6151
R2566 B.n345 B.n344 10.6151
R2567 B.n348 B.n345 10.6151
R2568 B.n349 B.n348 10.6151
R2569 B.n352 B.n349 10.6151
R2570 B.n353 B.n352 10.6151
R2571 B.n356 B.n353 10.6151
R2572 B.n357 B.n356 10.6151
R2573 B.n360 B.n357 10.6151
R2574 B.n361 B.n360 10.6151
R2575 B.n364 B.n361 10.6151
R2576 B.n365 B.n364 10.6151
R2577 B.n368 B.n365 10.6151
R2578 B.n369 B.n368 10.6151
R2579 B.n372 B.n369 10.6151
R2580 B.n373 B.n372 10.6151
R2581 B.n939 B.n373 10.6151
R2582 B.n761 B.n453 10.6151
R2583 B.n762 B.n761 10.6151
R2584 B.n763 B.n762 10.6151
R2585 B.n763 B.n445 10.6151
R2586 B.n773 B.n445 10.6151
R2587 B.n774 B.n773 10.6151
R2588 B.n775 B.n774 10.6151
R2589 B.n775 B.n437 10.6151
R2590 B.n785 B.n437 10.6151
R2591 B.n786 B.n785 10.6151
R2592 B.n787 B.n786 10.6151
R2593 B.n787 B.n429 10.6151
R2594 B.n797 B.n429 10.6151
R2595 B.n798 B.n797 10.6151
R2596 B.n799 B.n798 10.6151
R2597 B.n799 B.n421 10.6151
R2598 B.n809 B.n421 10.6151
R2599 B.n810 B.n809 10.6151
R2600 B.n811 B.n810 10.6151
R2601 B.n811 B.n413 10.6151
R2602 B.n821 B.n413 10.6151
R2603 B.n822 B.n821 10.6151
R2604 B.n823 B.n822 10.6151
R2605 B.n823 B.n406 10.6151
R2606 B.n834 B.n406 10.6151
R2607 B.n835 B.n834 10.6151
R2608 B.n836 B.n835 10.6151
R2609 B.n836 B.n398 10.6151
R2610 B.n846 B.n398 10.6151
R2611 B.n847 B.n846 10.6151
R2612 B.n848 B.n847 10.6151
R2613 B.n848 B.n390 10.6151
R2614 B.n858 B.n390 10.6151
R2615 B.n859 B.n858 10.6151
R2616 B.n860 B.n859 10.6151
R2617 B.n860 B.n382 10.6151
R2618 B.n870 B.n382 10.6151
R2619 B.n871 B.n870 10.6151
R2620 B.n873 B.n871 10.6151
R2621 B.n873 B.n872 10.6151
R2622 B.n872 B.n374 10.6151
R2623 B.n884 B.n374 10.6151
R2624 B.n885 B.n884 10.6151
R2625 B.n886 B.n885 10.6151
R2626 B.n887 B.n886 10.6151
R2627 B.n889 B.n887 10.6151
R2628 B.n890 B.n889 10.6151
R2629 B.n891 B.n890 10.6151
R2630 B.n892 B.n891 10.6151
R2631 B.n894 B.n892 10.6151
R2632 B.n895 B.n894 10.6151
R2633 B.n896 B.n895 10.6151
R2634 B.n897 B.n896 10.6151
R2635 B.n899 B.n897 10.6151
R2636 B.n900 B.n899 10.6151
R2637 B.n901 B.n900 10.6151
R2638 B.n902 B.n901 10.6151
R2639 B.n904 B.n902 10.6151
R2640 B.n905 B.n904 10.6151
R2641 B.n906 B.n905 10.6151
R2642 B.n907 B.n906 10.6151
R2643 B.n909 B.n907 10.6151
R2644 B.n910 B.n909 10.6151
R2645 B.n911 B.n910 10.6151
R2646 B.n912 B.n911 10.6151
R2647 B.n914 B.n912 10.6151
R2648 B.n915 B.n914 10.6151
R2649 B.n916 B.n915 10.6151
R2650 B.n917 B.n916 10.6151
R2651 B.n919 B.n917 10.6151
R2652 B.n920 B.n919 10.6151
R2653 B.n921 B.n920 10.6151
R2654 B.n922 B.n921 10.6151
R2655 B.n924 B.n922 10.6151
R2656 B.n925 B.n924 10.6151
R2657 B.n926 B.n925 10.6151
R2658 B.n927 B.n926 10.6151
R2659 B.n929 B.n927 10.6151
R2660 B.n930 B.n929 10.6151
R2661 B.n931 B.n930 10.6151
R2662 B.n932 B.n931 10.6151
R2663 B.n934 B.n932 10.6151
R2664 B.n935 B.n934 10.6151
R2665 B.n936 B.n935 10.6151
R2666 B.n937 B.n936 10.6151
R2667 B.n938 B.n937 10.6151
R2668 B.n755 B.n457 10.6151
R2669 B.n750 B.n457 10.6151
R2670 B.n750 B.n749 10.6151
R2671 B.n749 B.n748 10.6151
R2672 B.n748 B.n745 10.6151
R2673 B.n745 B.n744 10.6151
R2674 B.n744 B.n741 10.6151
R2675 B.n741 B.n740 10.6151
R2676 B.n740 B.n737 10.6151
R2677 B.n737 B.n736 10.6151
R2678 B.n736 B.n733 10.6151
R2679 B.n733 B.n732 10.6151
R2680 B.n732 B.n729 10.6151
R2681 B.n729 B.n728 10.6151
R2682 B.n728 B.n725 10.6151
R2683 B.n725 B.n724 10.6151
R2684 B.n724 B.n721 10.6151
R2685 B.n721 B.n720 10.6151
R2686 B.n720 B.n717 10.6151
R2687 B.n717 B.n716 10.6151
R2688 B.n716 B.n713 10.6151
R2689 B.n713 B.n712 10.6151
R2690 B.n712 B.n709 10.6151
R2691 B.n709 B.n708 10.6151
R2692 B.n708 B.n705 10.6151
R2693 B.n705 B.n704 10.6151
R2694 B.n704 B.n701 10.6151
R2695 B.n701 B.n700 10.6151
R2696 B.n700 B.n697 10.6151
R2697 B.n697 B.n696 10.6151
R2698 B.n696 B.n693 10.6151
R2699 B.n693 B.n692 10.6151
R2700 B.n692 B.n689 10.6151
R2701 B.n689 B.n688 10.6151
R2702 B.n688 B.n685 10.6151
R2703 B.n685 B.n684 10.6151
R2704 B.n684 B.n681 10.6151
R2705 B.n681 B.n680 10.6151
R2706 B.n680 B.n677 10.6151
R2707 B.n677 B.n676 10.6151
R2708 B.n676 B.n673 10.6151
R2709 B.n673 B.n672 10.6151
R2710 B.n672 B.n669 10.6151
R2711 B.n669 B.n668 10.6151
R2712 B.n668 B.n665 10.6151
R2713 B.n665 B.n664 10.6151
R2714 B.n664 B.n661 10.6151
R2715 B.n661 B.n660 10.6151
R2716 B.n660 B.n657 10.6151
R2717 B.n657 B.n656 10.6151
R2718 B.n656 B.n653 10.6151
R2719 B.n653 B.n652 10.6151
R2720 B.n652 B.n649 10.6151
R2721 B.n647 B.n644 10.6151
R2722 B.n644 B.n643 10.6151
R2723 B.n643 B.n640 10.6151
R2724 B.n640 B.n639 10.6151
R2725 B.n639 B.n636 10.6151
R2726 B.n636 B.n635 10.6151
R2727 B.n635 B.n632 10.6151
R2728 B.n632 B.n631 10.6151
R2729 B.n628 B.n627 10.6151
R2730 B.n627 B.n624 10.6151
R2731 B.n624 B.n623 10.6151
R2732 B.n623 B.n620 10.6151
R2733 B.n620 B.n619 10.6151
R2734 B.n619 B.n616 10.6151
R2735 B.n616 B.n615 10.6151
R2736 B.n615 B.n612 10.6151
R2737 B.n612 B.n611 10.6151
R2738 B.n611 B.n608 10.6151
R2739 B.n608 B.n607 10.6151
R2740 B.n607 B.n604 10.6151
R2741 B.n604 B.n603 10.6151
R2742 B.n603 B.n600 10.6151
R2743 B.n600 B.n599 10.6151
R2744 B.n599 B.n596 10.6151
R2745 B.n596 B.n595 10.6151
R2746 B.n595 B.n592 10.6151
R2747 B.n592 B.n591 10.6151
R2748 B.n591 B.n588 10.6151
R2749 B.n588 B.n587 10.6151
R2750 B.n587 B.n584 10.6151
R2751 B.n584 B.n583 10.6151
R2752 B.n583 B.n580 10.6151
R2753 B.n580 B.n579 10.6151
R2754 B.n579 B.n576 10.6151
R2755 B.n576 B.n575 10.6151
R2756 B.n575 B.n572 10.6151
R2757 B.n572 B.n571 10.6151
R2758 B.n571 B.n568 10.6151
R2759 B.n568 B.n567 10.6151
R2760 B.n567 B.n564 10.6151
R2761 B.n564 B.n563 10.6151
R2762 B.n563 B.n560 10.6151
R2763 B.n560 B.n559 10.6151
R2764 B.n559 B.n556 10.6151
R2765 B.n556 B.n555 10.6151
R2766 B.n555 B.n552 10.6151
R2767 B.n552 B.n551 10.6151
R2768 B.n551 B.n548 10.6151
R2769 B.n548 B.n547 10.6151
R2770 B.n547 B.n544 10.6151
R2771 B.n544 B.n543 10.6151
R2772 B.n543 B.n540 10.6151
R2773 B.n540 B.n539 10.6151
R2774 B.n539 B.n536 10.6151
R2775 B.n536 B.n535 10.6151
R2776 B.n535 B.n532 10.6151
R2777 B.n532 B.n531 10.6151
R2778 B.n531 B.n528 10.6151
R2779 B.n528 B.n527 10.6151
R2780 B.n527 B.n524 10.6151
R2781 B.n524 B.n523 10.6151
R2782 B.n757 B.n756 10.6151
R2783 B.n757 B.n449 10.6151
R2784 B.n767 B.n449 10.6151
R2785 B.n768 B.n767 10.6151
R2786 B.n769 B.n768 10.6151
R2787 B.n769 B.n441 10.6151
R2788 B.n779 B.n441 10.6151
R2789 B.n780 B.n779 10.6151
R2790 B.n781 B.n780 10.6151
R2791 B.n781 B.n433 10.6151
R2792 B.n791 B.n433 10.6151
R2793 B.n792 B.n791 10.6151
R2794 B.n793 B.n792 10.6151
R2795 B.n793 B.n425 10.6151
R2796 B.n803 B.n425 10.6151
R2797 B.n804 B.n803 10.6151
R2798 B.n805 B.n804 10.6151
R2799 B.n805 B.n417 10.6151
R2800 B.n815 B.n417 10.6151
R2801 B.n816 B.n815 10.6151
R2802 B.n817 B.n816 10.6151
R2803 B.n817 B.n409 10.6151
R2804 B.n828 B.n409 10.6151
R2805 B.n829 B.n828 10.6151
R2806 B.n830 B.n829 10.6151
R2807 B.n830 B.n402 10.6151
R2808 B.n840 B.n402 10.6151
R2809 B.n841 B.n840 10.6151
R2810 B.n842 B.n841 10.6151
R2811 B.n842 B.n394 10.6151
R2812 B.n852 B.n394 10.6151
R2813 B.n853 B.n852 10.6151
R2814 B.n854 B.n853 10.6151
R2815 B.n854 B.n386 10.6151
R2816 B.n864 B.n386 10.6151
R2817 B.n865 B.n864 10.6151
R2818 B.n866 B.n865 10.6151
R2819 B.n866 B.n378 10.6151
R2820 B.n877 B.n378 10.6151
R2821 B.n878 B.n877 10.6151
R2822 B.n879 B.n878 10.6151
R2823 B.n879 B.n0 10.6151
R2824 B.n1026 B.n1 10.6151
R2825 B.n1026 B.n1025 10.6151
R2826 B.n1025 B.n1024 10.6151
R2827 B.n1024 B.n10 10.6151
R2828 B.n1018 B.n10 10.6151
R2829 B.n1018 B.n1017 10.6151
R2830 B.n1017 B.n1016 10.6151
R2831 B.n1016 B.n17 10.6151
R2832 B.n1010 B.n17 10.6151
R2833 B.n1010 B.n1009 10.6151
R2834 B.n1009 B.n1008 10.6151
R2835 B.n1008 B.n24 10.6151
R2836 B.n1002 B.n24 10.6151
R2837 B.n1002 B.n1001 10.6151
R2838 B.n1001 B.n1000 10.6151
R2839 B.n1000 B.n31 10.6151
R2840 B.n994 B.n31 10.6151
R2841 B.n994 B.n993 10.6151
R2842 B.n993 B.n992 10.6151
R2843 B.n992 B.n37 10.6151
R2844 B.n986 B.n37 10.6151
R2845 B.n986 B.n985 10.6151
R2846 B.n985 B.n984 10.6151
R2847 B.n984 B.n45 10.6151
R2848 B.n978 B.n45 10.6151
R2849 B.n978 B.n977 10.6151
R2850 B.n977 B.n976 10.6151
R2851 B.n976 B.n52 10.6151
R2852 B.n970 B.n52 10.6151
R2853 B.n970 B.n969 10.6151
R2854 B.n969 B.n968 10.6151
R2855 B.n968 B.n59 10.6151
R2856 B.n962 B.n59 10.6151
R2857 B.n962 B.n961 10.6151
R2858 B.n961 B.n960 10.6151
R2859 B.n960 B.n66 10.6151
R2860 B.n954 B.n66 10.6151
R2861 B.n954 B.n953 10.6151
R2862 B.n953 B.n952 10.6151
R2863 B.n952 B.n73 10.6151
R2864 B.n946 B.n73 10.6151
R2865 B.n946 B.n945 10.6151
R2866 B.n783 B.t5 10.3074
R2867 B.t12 B.n964 10.3074
R2868 B.n251 B.n145 6.5566
R2869 B.n268 B.n267 6.5566
R2870 B.n648 B.n647 6.5566
R2871 B.n631 B.n521 6.5566
R2872 B.n248 B.n145 4.05904
R2873 B.n269 B.n268 4.05904
R2874 B.n649 B.n648 4.05904
R2875 B.n628 B.n521 4.05904
R2876 B.n1032 B.n0 2.81026
R2877 B.n1032 B.n1 2.81026
R2878 B.n825 B.t2 2.06187
R2879 B.n39 B.t3 2.06187
R2880 VN.n1 VN.t0 142.452
R2881 VN.n0 VN.t2 142.452
R2882 VN.n0 VN.t1 141.208
R2883 VN.n1 VN.t3 141.208
R2884 VN VN.n1 54.8225
R2885 VN VN.n0 2.09897
R2886 VDD2.n2 VDD2.n0 108.316
R2887 VDD2.n2 VDD2.n1 60.5836
R2888 VDD2.n1 VDD2.t0 1.23261
R2889 VDD2.n1 VDD2.t3 1.23261
R2890 VDD2.n0 VDD2.t1 1.23261
R2891 VDD2.n0 VDD2.t2 1.23261
R2892 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.150056f
C1 VN VTAIL 6.44773f
C2 VDD1 VTAIL 6.5373f
C3 VDD2 VP 0.458089f
C4 VP VN 7.66409f
C5 VDD1 VP 6.88526f
C6 VP VTAIL 6.46183f
C7 VDD2 VN 6.57821f
C8 VDD1 VDD2 1.26764f
C9 VDD2 VTAIL 6.59821f
C10 VDD2 B 4.654099f
C11 VDD1 B 9.54391f
C12 VTAIL B 13.097765f
C13 VN B 12.93845f
C14 VP B 11.334183f
C15 VDD2.t1 B 0.341351f
C16 VDD2.t2 B 0.341351f
C17 VDD2.n0 B 3.98531f
C18 VDD2.t0 B 0.341351f
C19 VDD2.t3 B 0.341351f
C20 VDD2.n1 B 3.09466f
C21 VDD2.n2 B 4.45541f
C22 VN.t1 B 3.42008f
C23 VN.t2 B 3.43041f
C24 VN.n0 B 2.0709f
C25 VN.t0 B 3.43041f
C26 VN.t3 B 3.42008f
C27 VN.n1 B 3.43837f
C28 VDD1.t0 B 0.343936f
C29 VDD1.t3 B 0.343936f
C30 VDD1.n0 B 3.11861f
C31 VDD1.t2 B 0.343936f
C32 VDD1.t1 B 0.343936f
C33 VDD1.n1 B 4.04448f
C34 VTAIL.n0 B 0.02111f
C35 VTAIL.n1 B 0.016018f
C36 VTAIL.n2 B 0.008607f
C37 VTAIL.n3 B 0.020345f
C38 VTAIL.n4 B 0.009114f
C39 VTAIL.n5 B 0.016018f
C40 VTAIL.n6 B 0.008861f
C41 VTAIL.n7 B 0.020345f
C42 VTAIL.n8 B 0.009114f
C43 VTAIL.n9 B 0.016018f
C44 VTAIL.n10 B 0.008607f
C45 VTAIL.n11 B 0.020345f
C46 VTAIL.n12 B 0.009114f
C47 VTAIL.n13 B 0.016018f
C48 VTAIL.n14 B 0.008607f
C49 VTAIL.n15 B 0.020345f
C50 VTAIL.n16 B 0.009114f
C51 VTAIL.n17 B 0.016018f
C52 VTAIL.n18 B 0.008607f
C53 VTAIL.n19 B 0.020345f
C54 VTAIL.n20 B 0.009114f
C55 VTAIL.n21 B 0.016018f
C56 VTAIL.n22 B 0.008607f
C57 VTAIL.n23 B 0.020345f
C58 VTAIL.n24 B 0.009114f
C59 VTAIL.n25 B 0.016018f
C60 VTAIL.n26 B 0.008607f
C61 VTAIL.n27 B 0.015259f
C62 VTAIL.n28 B 0.012018f
C63 VTAIL.t1 B 0.033605f
C64 VTAIL.n29 B 0.108771f
C65 VTAIL.n30 B 1.12071f
C66 VTAIL.n31 B 0.008607f
C67 VTAIL.n32 B 0.009114f
C68 VTAIL.n33 B 0.020345f
C69 VTAIL.n34 B 0.020345f
C70 VTAIL.n35 B 0.009114f
C71 VTAIL.n36 B 0.008607f
C72 VTAIL.n37 B 0.016018f
C73 VTAIL.n38 B 0.016018f
C74 VTAIL.n39 B 0.008607f
C75 VTAIL.n40 B 0.009114f
C76 VTAIL.n41 B 0.020345f
C77 VTAIL.n42 B 0.020345f
C78 VTAIL.n43 B 0.009114f
C79 VTAIL.n44 B 0.008607f
C80 VTAIL.n45 B 0.016018f
C81 VTAIL.n46 B 0.016018f
C82 VTAIL.n47 B 0.008607f
C83 VTAIL.n48 B 0.009114f
C84 VTAIL.n49 B 0.020345f
C85 VTAIL.n50 B 0.020345f
C86 VTAIL.n51 B 0.009114f
C87 VTAIL.n52 B 0.008607f
C88 VTAIL.n53 B 0.016018f
C89 VTAIL.n54 B 0.016018f
C90 VTAIL.n55 B 0.008607f
C91 VTAIL.n56 B 0.009114f
C92 VTAIL.n57 B 0.020345f
C93 VTAIL.n58 B 0.020345f
C94 VTAIL.n59 B 0.009114f
C95 VTAIL.n60 B 0.008607f
C96 VTAIL.n61 B 0.016018f
C97 VTAIL.n62 B 0.016018f
C98 VTAIL.n63 B 0.008607f
C99 VTAIL.n64 B 0.009114f
C100 VTAIL.n65 B 0.020345f
C101 VTAIL.n66 B 0.020345f
C102 VTAIL.n67 B 0.009114f
C103 VTAIL.n68 B 0.008607f
C104 VTAIL.n69 B 0.016018f
C105 VTAIL.n70 B 0.016018f
C106 VTAIL.n71 B 0.008607f
C107 VTAIL.n72 B 0.008607f
C108 VTAIL.n73 B 0.009114f
C109 VTAIL.n74 B 0.020345f
C110 VTAIL.n75 B 0.020345f
C111 VTAIL.n76 B 0.020345f
C112 VTAIL.n77 B 0.008861f
C113 VTAIL.n78 B 0.008607f
C114 VTAIL.n79 B 0.016018f
C115 VTAIL.n80 B 0.016018f
C116 VTAIL.n81 B 0.008607f
C117 VTAIL.n82 B 0.009114f
C118 VTAIL.n83 B 0.020345f
C119 VTAIL.n84 B 0.041559f
C120 VTAIL.n85 B 0.009114f
C121 VTAIL.n86 B 0.008607f
C122 VTAIL.n87 B 0.036806f
C123 VTAIL.n88 B 0.022992f
C124 VTAIL.n89 B 0.128242f
C125 VTAIL.n90 B 0.02111f
C126 VTAIL.n91 B 0.016018f
C127 VTAIL.n92 B 0.008607f
C128 VTAIL.n93 B 0.020345f
C129 VTAIL.n94 B 0.009114f
C130 VTAIL.n95 B 0.016018f
C131 VTAIL.n96 B 0.008861f
C132 VTAIL.n97 B 0.020345f
C133 VTAIL.n98 B 0.009114f
C134 VTAIL.n99 B 0.016018f
C135 VTAIL.n100 B 0.008607f
C136 VTAIL.n101 B 0.020345f
C137 VTAIL.n102 B 0.009114f
C138 VTAIL.n103 B 0.016018f
C139 VTAIL.n104 B 0.008607f
C140 VTAIL.n105 B 0.020345f
C141 VTAIL.n106 B 0.009114f
C142 VTAIL.n107 B 0.016018f
C143 VTAIL.n108 B 0.008607f
C144 VTAIL.n109 B 0.020345f
C145 VTAIL.n110 B 0.009114f
C146 VTAIL.n111 B 0.016018f
C147 VTAIL.n112 B 0.008607f
C148 VTAIL.n113 B 0.020345f
C149 VTAIL.n114 B 0.009114f
C150 VTAIL.n115 B 0.016018f
C151 VTAIL.n116 B 0.008607f
C152 VTAIL.n117 B 0.015259f
C153 VTAIL.n118 B 0.012018f
C154 VTAIL.t6 B 0.033605f
C155 VTAIL.n119 B 0.108771f
C156 VTAIL.n120 B 1.12071f
C157 VTAIL.n121 B 0.008607f
C158 VTAIL.n122 B 0.009114f
C159 VTAIL.n123 B 0.020345f
C160 VTAIL.n124 B 0.020345f
C161 VTAIL.n125 B 0.009114f
C162 VTAIL.n126 B 0.008607f
C163 VTAIL.n127 B 0.016018f
C164 VTAIL.n128 B 0.016018f
C165 VTAIL.n129 B 0.008607f
C166 VTAIL.n130 B 0.009114f
C167 VTAIL.n131 B 0.020345f
C168 VTAIL.n132 B 0.020345f
C169 VTAIL.n133 B 0.009114f
C170 VTAIL.n134 B 0.008607f
C171 VTAIL.n135 B 0.016018f
C172 VTAIL.n136 B 0.016018f
C173 VTAIL.n137 B 0.008607f
C174 VTAIL.n138 B 0.009114f
C175 VTAIL.n139 B 0.020345f
C176 VTAIL.n140 B 0.020345f
C177 VTAIL.n141 B 0.009114f
C178 VTAIL.n142 B 0.008607f
C179 VTAIL.n143 B 0.016018f
C180 VTAIL.n144 B 0.016018f
C181 VTAIL.n145 B 0.008607f
C182 VTAIL.n146 B 0.009114f
C183 VTAIL.n147 B 0.020345f
C184 VTAIL.n148 B 0.020345f
C185 VTAIL.n149 B 0.009114f
C186 VTAIL.n150 B 0.008607f
C187 VTAIL.n151 B 0.016018f
C188 VTAIL.n152 B 0.016018f
C189 VTAIL.n153 B 0.008607f
C190 VTAIL.n154 B 0.009114f
C191 VTAIL.n155 B 0.020345f
C192 VTAIL.n156 B 0.020345f
C193 VTAIL.n157 B 0.009114f
C194 VTAIL.n158 B 0.008607f
C195 VTAIL.n159 B 0.016018f
C196 VTAIL.n160 B 0.016018f
C197 VTAIL.n161 B 0.008607f
C198 VTAIL.n162 B 0.008607f
C199 VTAIL.n163 B 0.009114f
C200 VTAIL.n164 B 0.020345f
C201 VTAIL.n165 B 0.020345f
C202 VTAIL.n166 B 0.020345f
C203 VTAIL.n167 B 0.008861f
C204 VTAIL.n168 B 0.008607f
C205 VTAIL.n169 B 0.016018f
C206 VTAIL.n170 B 0.016018f
C207 VTAIL.n171 B 0.008607f
C208 VTAIL.n172 B 0.009114f
C209 VTAIL.n173 B 0.020345f
C210 VTAIL.n174 B 0.041559f
C211 VTAIL.n175 B 0.009114f
C212 VTAIL.n176 B 0.008607f
C213 VTAIL.n177 B 0.036806f
C214 VTAIL.n178 B 0.022992f
C215 VTAIL.n179 B 0.212671f
C216 VTAIL.n180 B 0.02111f
C217 VTAIL.n181 B 0.016018f
C218 VTAIL.n182 B 0.008607f
C219 VTAIL.n183 B 0.020345f
C220 VTAIL.n184 B 0.009114f
C221 VTAIL.n185 B 0.016018f
C222 VTAIL.n186 B 0.008861f
C223 VTAIL.n187 B 0.020345f
C224 VTAIL.n188 B 0.009114f
C225 VTAIL.n189 B 0.016018f
C226 VTAIL.n190 B 0.008607f
C227 VTAIL.n191 B 0.020345f
C228 VTAIL.n192 B 0.009114f
C229 VTAIL.n193 B 0.016018f
C230 VTAIL.n194 B 0.008607f
C231 VTAIL.n195 B 0.020345f
C232 VTAIL.n196 B 0.009114f
C233 VTAIL.n197 B 0.016018f
C234 VTAIL.n198 B 0.008607f
C235 VTAIL.n199 B 0.020345f
C236 VTAIL.n200 B 0.009114f
C237 VTAIL.n201 B 0.016018f
C238 VTAIL.n202 B 0.008607f
C239 VTAIL.n203 B 0.020345f
C240 VTAIL.n204 B 0.009114f
C241 VTAIL.n205 B 0.016018f
C242 VTAIL.n206 B 0.008607f
C243 VTAIL.n207 B 0.015259f
C244 VTAIL.n208 B 0.012018f
C245 VTAIL.t4 B 0.033605f
C246 VTAIL.n209 B 0.108771f
C247 VTAIL.n210 B 1.12071f
C248 VTAIL.n211 B 0.008607f
C249 VTAIL.n212 B 0.009114f
C250 VTAIL.n213 B 0.020345f
C251 VTAIL.n214 B 0.020345f
C252 VTAIL.n215 B 0.009114f
C253 VTAIL.n216 B 0.008607f
C254 VTAIL.n217 B 0.016018f
C255 VTAIL.n218 B 0.016018f
C256 VTAIL.n219 B 0.008607f
C257 VTAIL.n220 B 0.009114f
C258 VTAIL.n221 B 0.020345f
C259 VTAIL.n222 B 0.020345f
C260 VTAIL.n223 B 0.009114f
C261 VTAIL.n224 B 0.008607f
C262 VTAIL.n225 B 0.016018f
C263 VTAIL.n226 B 0.016018f
C264 VTAIL.n227 B 0.008607f
C265 VTAIL.n228 B 0.009114f
C266 VTAIL.n229 B 0.020345f
C267 VTAIL.n230 B 0.020345f
C268 VTAIL.n231 B 0.009114f
C269 VTAIL.n232 B 0.008607f
C270 VTAIL.n233 B 0.016018f
C271 VTAIL.n234 B 0.016018f
C272 VTAIL.n235 B 0.008607f
C273 VTAIL.n236 B 0.009114f
C274 VTAIL.n237 B 0.020345f
C275 VTAIL.n238 B 0.020345f
C276 VTAIL.n239 B 0.009114f
C277 VTAIL.n240 B 0.008607f
C278 VTAIL.n241 B 0.016018f
C279 VTAIL.n242 B 0.016018f
C280 VTAIL.n243 B 0.008607f
C281 VTAIL.n244 B 0.009114f
C282 VTAIL.n245 B 0.020345f
C283 VTAIL.n246 B 0.020345f
C284 VTAIL.n247 B 0.009114f
C285 VTAIL.n248 B 0.008607f
C286 VTAIL.n249 B 0.016018f
C287 VTAIL.n250 B 0.016018f
C288 VTAIL.n251 B 0.008607f
C289 VTAIL.n252 B 0.008607f
C290 VTAIL.n253 B 0.009114f
C291 VTAIL.n254 B 0.020345f
C292 VTAIL.n255 B 0.020345f
C293 VTAIL.n256 B 0.020345f
C294 VTAIL.n257 B 0.008861f
C295 VTAIL.n258 B 0.008607f
C296 VTAIL.n259 B 0.016018f
C297 VTAIL.n260 B 0.016018f
C298 VTAIL.n261 B 0.008607f
C299 VTAIL.n262 B 0.009114f
C300 VTAIL.n263 B 0.020345f
C301 VTAIL.n264 B 0.041559f
C302 VTAIL.n265 B 0.009114f
C303 VTAIL.n266 B 0.008607f
C304 VTAIL.n267 B 0.036806f
C305 VTAIL.n268 B 0.022992f
C306 VTAIL.n269 B 1.2959f
C307 VTAIL.n270 B 0.02111f
C308 VTAIL.n271 B 0.016018f
C309 VTAIL.n272 B 0.008607f
C310 VTAIL.n273 B 0.020345f
C311 VTAIL.n274 B 0.009114f
C312 VTAIL.n275 B 0.016018f
C313 VTAIL.n276 B 0.008861f
C314 VTAIL.n277 B 0.020345f
C315 VTAIL.n278 B 0.008607f
C316 VTAIL.n279 B 0.009114f
C317 VTAIL.n280 B 0.016018f
C318 VTAIL.n281 B 0.008607f
C319 VTAIL.n282 B 0.020345f
C320 VTAIL.n283 B 0.009114f
C321 VTAIL.n284 B 0.016018f
C322 VTAIL.n285 B 0.008607f
C323 VTAIL.n286 B 0.020345f
C324 VTAIL.n287 B 0.009114f
C325 VTAIL.n288 B 0.016018f
C326 VTAIL.n289 B 0.008607f
C327 VTAIL.n290 B 0.020345f
C328 VTAIL.n291 B 0.009114f
C329 VTAIL.n292 B 0.016018f
C330 VTAIL.n293 B 0.008607f
C331 VTAIL.n294 B 0.020345f
C332 VTAIL.n295 B 0.009114f
C333 VTAIL.n296 B 0.016018f
C334 VTAIL.n297 B 0.008607f
C335 VTAIL.n298 B 0.015259f
C336 VTAIL.n299 B 0.012018f
C337 VTAIL.t2 B 0.033605f
C338 VTAIL.n300 B 0.108771f
C339 VTAIL.n301 B 1.12071f
C340 VTAIL.n302 B 0.008607f
C341 VTAIL.n303 B 0.009114f
C342 VTAIL.n304 B 0.020345f
C343 VTAIL.n305 B 0.020345f
C344 VTAIL.n306 B 0.009114f
C345 VTAIL.n307 B 0.008607f
C346 VTAIL.n308 B 0.016018f
C347 VTAIL.n309 B 0.016018f
C348 VTAIL.n310 B 0.008607f
C349 VTAIL.n311 B 0.009114f
C350 VTAIL.n312 B 0.020345f
C351 VTAIL.n313 B 0.020345f
C352 VTAIL.n314 B 0.009114f
C353 VTAIL.n315 B 0.008607f
C354 VTAIL.n316 B 0.016018f
C355 VTAIL.n317 B 0.016018f
C356 VTAIL.n318 B 0.008607f
C357 VTAIL.n319 B 0.009114f
C358 VTAIL.n320 B 0.020345f
C359 VTAIL.n321 B 0.020345f
C360 VTAIL.n322 B 0.009114f
C361 VTAIL.n323 B 0.008607f
C362 VTAIL.n324 B 0.016018f
C363 VTAIL.n325 B 0.016018f
C364 VTAIL.n326 B 0.008607f
C365 VTAIL.n327 B 0.009114f
C366 VTAIL.n328 B 0.020345f
C367 VTAIL.n329 B 0.020345f
C368 VTAIL.n330 B 0.009114f
C369 VTAIL.n331 B 0.008607f
C370 VTAIL.n332 B 0.016018f
C371 VTAIL.n333 B 0.016018f
C372 VTAIL.n334 B 0.008607f
C373 VTAIL.n335 B 0.009114f
C374 VTAIL.n336 B 0.020345f
C375 VTAIL.n337 B 0.020345f
C376 VTAIL.n338 B 0.009114f
C377 VTAIL.n339 B 0.008607f
C378 VTAIL.n340 B 0.016018f
C379 VTAIL.n341 B 0.016018f
C380 VTAIL.n342 B 0.008607f
C381 VTAIL.n343 B 0.009114f
C382 VTAIL.n344 B 0.020345f
C383 VTAIL.n345 B 0.020345f
C384 VTAIL.n346 B 0.020345f
C385 VTAIL.n347 B 0.008861f
C386 VTAIL.n348 B 0.008607f
C387 VTAIL.n349 B 0.016018f
C388 VTAIL.n350 B 0.016018f
C389 VTAIL.n351 B 0.008607f
C390 VTAIL.n352 B 0.009114f
C391 VTAIL.n353 B 0.020345f
C392 VTAIL.n354 B 0.041559f
C393 VTAIL.n355 B 0.009114f
C394 VTAIL.n356 B 0.008607f
C395 VTAIL.n357 B 0.036806f
C396 VTAIL.n358 B 0.022992f
C397 VTAIL.n359 B 1.2959f
C398 VTAIL.n360 B 0.02111f
C399 VTAIL.n361 B 0.016018f
C400 VTAIL.n362 B 0.008607f
C401 VTAIL.n363 B 0.020345f
C402 VTAIL.n364 B 0.009114f
C403 VTAIL.n365 B 0.016018f
C404 VTAIL.n366 B 0.008861f
C405 VTAIL.n367 B 0.020345f
C406 VTAIL.n368 B 0.008607f
C407 VTAIL.n369 B 0.009114f
C408 VTAIL.n370 B 0.016018f
C409 VTAIL.n371 B 0.008607f
C410 VTAIL.n372 B 0.020345f
C411 VTAIL.n373 B 0.009114f
C412 VTAIL.n374 B 0.016018f
C413 VTAIL.n375 B 0.008607f
C414 VTAIL.n376 B 0.020345f
C415 VTAIL.n377 B 0.009114f
C416 VTAIL.n378 B 0.016018f
C417 VTAIL.n379 B 0.008607f
C418 VTAIL.n380 B 0.020345f
C419 VTAIL.n381 B 0.009114f
C420 VTAIL.n382 B 0.016018f
C421 VTAIL.n383 B 0.008607f
C422 VTAIL.n384 B 0.020345f
C423 VTAIL.n385 B 0.009114f
C424 VTAIL.n386 B 0.016018f
C425 VTAIL.n387 B 0.008607f
C426 VTAIL.n388 B 0.015259f
C427 VTAIL.n389 B 0.012018f
C428 VTAIL.t0 B 0.033605f
C429 VTAIL.n390 B 0.108771f
C430 VTAIL.n391 B 1.12071f
C431 VTAIL.n392 B 0.008607f
C432 VTAIL.n393 B 0.009114f
C433 VTAIL.n394 B 0.020345f
C434 VTAIL.n395 B 0.020345f
C435 VTAIL.n396 B 0.009114f
C436 VTAIL.n397 B 0.008607f
C437 VTAIL.n398 B 0.016018f
C438 VTAIL.n399 B 0.016018f
C439 VTAIL.n400 B 0.008607f
C440 VTAIL.n401 B 0.009114f
C441 VTAIL.n402 B 0.020345f
C442 VTAIL.n403 B 0.020345f
C443 VTAIL.n404 B 0.009114f
C444 VTAIL.n405 B 0.008607f
C445 VTAIL.n406 B 0.016018f
C446 VTAIL.n407 B 0.016018f
C447 VTAIL.n408 B 0.008607f
C448 VTAIL.n409 B 0.009114f
C449 VTAIL.n410 B 0.020345f
C450 VTAIL.n411 B 0.020345f
C451 VTAIL.n412 B 0.009114f
C452 VTAIL.n413 B 0.008607f
C453 VTAIL.n414 B 0.016018f
C454 VTAIL.n415 B 0.016018f
C455 VTAIL.n416 B 0.008607f
C456 VTAIL.n417 B 0.009114f
C457 VTAIL.n418 B 0.020345f
C458 VTAIL.n419 B 0.020345f
C459 VTAIL.n420 B 0.009114f
C460 VTAIL.n421 B 0.008607f
C461 VTAIL.n422 B 0.016018f
C462 VTAIL.n423 B 0.016018f
C463 VTAIL.n424 B 0.008607f
C464 VTAIL.n425 B 0.009114f
C465 VTAIL.n426 B 0.020345f
C466 VTAIL.n427 B 0.020345f
C467 VTAIL.n428 B 0.009114f
C468 VTAIL.n429 B 0.008607f
C469 VTAIL.n430 B 0.016018f
C470 VTAIL.n431 B 0.016018f
C471 VTAIL.n432 B 0.008607f
C472 VTAIL.n433 B 0.009114f
C473 VTAIL.n434 B 0.020345f
C474 VTAIL.n435 B 0.020345f
C475 VTAIL.n436 B 0.020345f
C476 VTAIL.n437 B 0.008861f
C477 VTAIL.n438 B 0.008607f
C478 VTAIL.n439 B 0.016018f
C479 VTAIL.n440 B 0.016018f
C480 VTAIL.n441 B 0.008607f
C481 VTAIL.n442 B 0.009114f
C482 VTAIL.n443 B 0.020345f
C483 VTAIL.n444 B 0.041559f
C484 VTAIL.n445 B 0.009114f
C485 VTAIL.n446 B 0.008607f
C486 VTAIL.n447 B 0.036806f
C487 VTAIL.n448 B 0.022992f
C488 VTAIL.n449 B 0.212671f
C489 VTAIL.n450 B 0.02111f
C490 VTAIL.n451 B 0.016018f
C491 VTAIL.n452 B 0.008607f
C492 VTAIL.n453 B 0.020345f
C493 VTAIL.n454 B 0.009114f
C494 VTAIL.n455 B 0.016018f
C495 VTAIL.n456 B 0.008861f
C496 VTAIL.n457 B 0.020345f
C497 VTAIL.n458 B 0.008607f
C498 VTAIL.n459 B 0.009114f
C499 VTAIL.n460 B 0.016018f
C500 VTAIL.n461 B 0.008607f
C501 VTAIL.n462 B 0.020345f
C502 VTAIL.n463 B 0.009114f
C503 VTAIL.n464 B 0.016018f
C504 VTAIL.n465 B 0.008607f
C505 VTAIL.n466 B 0.020345f
C506 VTAIL.n467 B 0.009114f
C507 VTAIL.n468 B 0.016018f
C508 VTAIL.n469 B 0.008607f
C509 VTAIL.n470 B 0.020345f
C510 VTAIL.n471 B 0.009114f
C511 VTAIL.n472 B 0.016018f
C512 VTAIL.n473 B 0.008607f
C513 VTAIL.n474 B 0.020345f
C514 VTAIL.n475 B 0.009114f
C515 VTAIL.n476 B 0.016018f
C516 VTAIL.n477 B 0.008607f
C517 VTAIL.n478 B 0.015259f
C518 VTAIL.n479 B 0.012018f
C519 VTAIL.t7 B 0.033605f
C520 VTAIL.n480 B 0.108771f
C521 VTAIL.n481 B 1.12071f
C522 VTAIL.n482 B 0.008607f
C523 VTAIL.n483 B 0.009114f
C524 VTAIL.n484 B 0.020345f
C525 VTAIL.n485 B 0.020345f
C526 VTAIL.n486 B 0.009114f
C527 VTAIL.n487 B 0.008607f
C528 VTAIL.n488 B 0.016018f
C529 VTAIL.n489 B 0.016018f
C530 VTAIL.n490 B 0.008607f
C531 VTAIL.n491 B 0.009114f
C532 VTAIL.n492 B 0.020345f
C533 VTAIL.n493 B 0.020345f
C534 VTAIL.n494 B 0.009114f
C535 VTAIL.n495 B 0.008607f
C536 VTAIL.n496 B 0.016018f
C537 VTAIL.n497 B 0.016018f
C538 VTAIL.n498 B 0.008607f
C539 VTAIL.n499 B 0.009114f
C540 VTAIL.n500 B 0.020345f
C541 VTAIL.n501 B 0.020345f
C542 VTAIL.n502 B 0.009114f
C543 VTAIL.n503 B 0.008607f
C544 VTAIL.n504 B 0.016018f
C545 VTAIL.n505 B 0.016018f
C546 VTAIL.n506 B 0.008607f
C547 VTAIL.n507 B 0.009114f
C548 VTAIL.n508 B 0.020345f
C549 VTAIL.n509 B 0.020345f
C550 VTAIL.n510 B 0.009114f
C551 VTAIL.n511 B 0.008607f
C552 VTAIL.n512 B 0.016018f
C553 VTAIL.n513 B 0.016018f
C554 VTAIL.n514 B 0.008607f
C555 VTAIL.n515 B 0.009114f
C556 VTAIL.n516 B 0.020345f
C557 VTAIL.n517 B 0.020345f
C558 VTAIL.n518 B 0.009114f
C559 VTAIL.n519 B 0.008607f
C560 VTAIL.n520 B 0.016018f
C561 VTAIL.n521 B 0.016018f
C562 VTAIL.n522 B 0.008607f
C563 VTAIL.n523 B 0.009114f
C564 VTAIL.n524 B 0.020345f
C565 VTAIL.n525 B 0.020345f
C566 VTAIL.n526 B 0.020345f
C567 VTAIL.n527 B 0.008861f
C568 VTAIL.n528 B 0.008607f
C569 VTAIL.n529 B 0.016018f
C570 VTAIL.n530 B 0.016018f
C571 VTAIL.n531 B 0.008607f
C572 VTAIL.n532 B 0.009114f
C573 VTAIL.n533 B 0.020345f
C574 VTAIL.n534 B 0.041559f
C575 VTAIL.n535 B 0.009114f
C576 VTAIL.n536 B 0.008607f
C577 VTAIL.n537 B 0.036806f
C578 VTAIL.n538 B 0.022992f
C579 VTAIL.n539 B 0.212671f
C580 VTAIL.n540 B 0.02111f
C581 VTAIL.n541 B 0.016018f
C582 VTAIL.n542 B 0.008607f
C583 VTAIL.n543 B 0.020345f
C584 VTAIL.n544 B 0.009114f
C585 VTAIL.n545 B 0.016018f
C586 VTAIL.n546 B 0.008861f
C587 VTAIL.n547 B 0.020345f
C588 VTAIL.n548 B 0.008607f
C589 VTAIL.n549 B 0.009114f
C590 VTAIL.n550 B 0.016018f
C591 VTAIL.n551 B 0.008607f
C592 VTAIL.n552 B 0.020345f
C593 VTAIL.n553 B 0.009114f
C594 VTAIL.n554 B 0.016018f
C595 VTAIL.n555 B 0.008607f
C596 VTAIL.n556 B 0.020345f
C597 VTAIL.n557 B 0.009114f
C598 VTAIL.n558 B 0.016018f
C599 VTAIL.n559 B 0.008607f
C600 VTAIL.n560 B 0.020345f
C601 VTAIL.n561 B 0.009114f
C602 VTAIL.n562 B 0.016018f
C603 VTAIL.n563 B 0.008607f
C604 VTAIL.n564 B 0.020345f
C605 VTAIL.n565 B 0.009114f
C606 VTAIL.n566 B 0.016018f
C607 VTAIL.n567 B 0.008607f
C608 VTAIL.n568 B 0.015259f
C609 VTAIL.n569 B 0.012018f
C610 VTAIL.t5 B 0.033605f
C611 VTAIL.n570 B 0.108771f
C612 VTAIL.n571 B 1.12071f
C613 VTAIL.n572 B 0.008607f
C614 VTAIL.n573 B 0.009114f
C615 VTAIL.n574 B 0.020345f
C616 VTAIL.n575 B 0.020345f
C617 VTAIL.n576 B 0.009114f
C618 VTAIL.n577 B 0.008607f
C619 VTAIL.n578 B 0.016018f
C620 VTAIL.n579 B 0.016018f
C621 VTAIL.n580 B 0.008607f
C622 VTAIL.n581 B 0.009114f
C623 VTAIL.n582 B 0.020345f
C624 VTAIL.n583 B 0.020345f
C625 VTAIL.n584 B 0.009114f
C626 VTAIL.n585 B 0.008607f
C627 VTAIL.n586 B 0.016018f
C628 VTAIL.n587 B 0.016018f
C629 VTAIL.n588 B 0.008607f
C630 VTAIL.n589 B 0.009114f
C631 VTAIL.n590 B 0.020345f
C632 VTAIL.n591 B 0.020345f
C633 VTAIL.n592 B 0.009114f
C634 VTAIL.n593 B 0.008607f
C635 VTAIL.n594 B 0.016018f
C636 VTAIL.n595 B 0.016018f
C637 VTAIL.n596 B 0.008607f
C638 VTAIL.n597 B 0.009114f
C639 VTAIL.n598 B 0.020345f
C640 VTAIL.n599 B 0.020345f
C641 VTAIL.n600 B 0.009114f
C642 VTAIL.n601 B 0.008607f
C643 VTAIL.n602 B 0.016018f
C644 VTAIL.n603 B 0.016018f
C645 VTAIL.n604 B 0.008607f
C646 VTAIL.n605 B 0.009114f
C647 VTAIL.n606 B 0.020345f
C648 VTAIL.n607 B 0.020345f
C649 VTAIL.n608 B 0.009114f
C650 VTAIL.n609 B 0.008607f
C651 VTAIL.n610 B 0.016018f
C652 VTAIL.n611 B 0.016018f
C653 VTAIL.n612 B 0.008607f
C654 VTAIL.n613 B 0.009114f
C655 VTAIL.n614 B 0.020345f
C656 VTAIL.n615 B 0.020345f
C657 VTAIL.n616 B 0.020345f
C658 VTAIL.n617 B 0.008861f
C659 VTAIL.n618 B 0.008607f
C660 VTAIL.n619 B 0.016018f
C661 VTAIL.n620 B 0.016018f
C662 VTAIL.n621 B 0.008607f
C663 VTAIL.n622 B 0.009114f
C664 VTAIL.n623 B 0.020345f
C665 VTAIL.n624 B 0.041559f
C666 VTAIL.n625 B 0.009114f
C667 VTAIL.n626 B 0.008607f
C668 VTAIL.n627 B 0.036806f
C669 VTAIL.n628 B 0.022992f
C670 VTAIL.n629 B 1.2959f
C671 VTAIL.n630 B 0.02111f
C672 VTAIL.n631 B 0.016018f
C673 VTAIL.n632 B 0.008607f
C674 VTAIL.n633 B 0.020345f
C675 VTAIL.n634 B 0.009114f
C676 VTAIL.n635 B 0.016018f
C677 VTAIL.n636 B 0.008861f
C678 VTAIL.n637 B 0.020345f
C679 VTAIL.n638 B 0.009114f
C680 VTAIL.n639 B 0.016018f
C681 VTAIL.n640 B 0.008607f
C682 VTAIL.n641 B 0.020345f
C683 VTAIL.n642 B 0.009114f
C684 VTAIL.n643 B 0.016018f
C685 VTAIL.n644 B 0.008607f
C686 VTAIL.n645 B 0.020345f
C687 VTAIL.n646 B 0.009114f
C688 VTAIL.n647 B 0.016018f
C689 VTAIL.n648 B 0.008607f
C690 VTAIL.n649 B 0.020345f
C691 VTAIL.n650 B 0.009114f
C692 VTAIL.n651 B 0.016018f
C693 VTAIL.n652 B 0.008607f
C694 VTAIL.n653 B 0.020345f
C695 VTAIL.n654 B 0.009114f
C696 VTAIL.n655 B 0.016018f
C697 VTAIL.n656 B 0.008607f
C698 VTAIL.n657 B 0.015259f
C699 VTAIL.n658 B 0.012018f
C700 VTAIL.t3 B 0.033605f
C701 VTAIL.n659 B 0.108771f
C702 VTAIL.n660 B 1.12071f
C703 VTAIL.n661 B 0.008607f
C704 VTAIL.n662 B 0.009114f
C705 VTAIL.n663 B 0.020345f
C706 VTAIL.n664 B 0.020345f
C707 VTAIL.n665 B 0.009114f
C708 VTAIL.n666 B 0.008607f
C709 VTAIL.n667 B 0.016018f
C710 VTAIL.n668 B 0.016018f
C711 VTAIL.n669 B 0.008607f
C712 VTAIL.n670 B 0.009114f
C713 VTAIL.n671 B 0.020345f
C714 VTAIL.n672 B 0.020345f
C715 VTAIL.n673 B 0.009114f
C716 VTAIL.n674 B 0.008607f
C717 VTAIL.n675 B 0.016018f
C718 VTAIL.n676 B 0.016018f
C719 VTAIL.n677 B 0.008607f
C720 VTAIL.n678 B 0.009114f
C721 VTAIL.n679 B 0.020345f
C722 VTAIL.n680 B 0.020345f
C723 VTAIL.n681 B 0.009114f
C724 VTAIL.n682 B 0.008607f
C725 VTAIL.n683 B 0.016018f
C726 VTAIL.n684 B 0.016018f
C727 VTAIL.n685 B 0.008607f
C728 VTAIL.n686 B 0.009114f
C729 VTAIL.n687 B 0.020345f
C730 VTAIL.n688 B 0.020345f
C731 VTAIL.n689 B 0.009114f
C732 VTAIL.n690 B 0.008607f
C733 VTAIL.n691 B 0.016018f
C734 VTAIL.n692 B 0.016018f
C735 VTAIL.n693 B 0.008607f
C736 VTAIL.n694 B 0.009114f
C737 VTAIL.n695 B 0.020345f
C738 VTAIL.n696 B 0.020345f
C739 VTAIL.n697 B 0.009114f
C740 VTAIL.n698 B 0.008607f
C741 VTAIL.n699 B 0.016018f
C742 VTAIL.n700 B 0.016018f
C743 VTAIL.n701 B 0.008607f
C744 VTAIL.n702 B 0.008607f
C745 VTAIL.n703 B 0.009114f
C746 VTAIL.n704 B 0.020345f
C747 VTAIL.n705 B 0.020345f
C748 VTAIL.n706 B 0.020345f
C749 VTAIL.n707 B 0.008861f
C750 VTAIL.n708 B 0.008607f
C751 VTAIL.n709 B 0.016018f
C752 VTAIL.n710 B 0.016018f
C753 VTAIL.n711 B 0.008607f
C754 VTAIL.n712 B 0.009114f
C755 VTAIL.n713 B 0.020345f
C756 VTAIL.n714 B 0.041559f
C757 VTAIL.n715 B 0.009114f
C758 VTAIL.n716 B 0.008607f
C759 VTAIL.n717 B 0.036806f
C760 VTAIL.n718 B 0.022992f
C761 VTAIL.n719 B 1.20547f
C762 VP.t2 B 3.19163f
C763 VP.n0 B 1.18516f
C764 VP.n1 B 0.020103f
C765 VP.n2 B 0.029347f
C766 VP.n3 B 0.020103f
C767 VP.n4 B 0.026922f
C768 VP.t3 B 3.50138f
C769 VP.t0 B 3.49084f
C770 VP.n5 B 3.50156f
C771 VP.t1 B 3.19163f
C772 VP.n6 B 1.18516f
C773 VP.n7 B 1.30639f
C774 VP.n8 B 0.032445f
C775 VP.n9 B 0.020103f
C776 VP.n10 B 0.037467f
C777 VP.n11 B 0.037467f
C778 VP.n12 B 0.029347f
C779 VP.n13 B 0.020103f
C780 VP.n14 B 0.020103f
C781 VP.n15 B 0.020103f
C782 VP.n16 B 0.037467f
C783 VP.n17 B 0.037467f
C784 VP.n18 B 0.026922f
C785 VP.n19 B 0.032445f
C786 VP.n20 B 0.054554f
.ends

