* NGSPICE file created from diff_pair_sample_0993.ext - technology: sky130A

.subckt diff_pair_sample_0993 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X1 VTAIL.t14 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X2 VDD1.t9 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=5.0271 ps=26.56 w=12.89 l=0.39
X3 VDD1.t8 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=5.0271 ps=26.56 w=12.89 l=0.39
X4 VTAIL.t13 VN.t2 VDD2.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X5 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=0 ps=0 w=12.89 l=0.39
X6 VDD2.t4 VN.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X7 VDD1.t7 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X8 VDD1.t6 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=2.12685 ps=13.22 w=12.89 l=0.39
X9 VTAIL.t3 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X10 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=0 ps=0 w=12.89 l=0.39
X11 VDD2.t7 VN.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=5.0271 ps=26.56 w=12.89 l=0.39
X12 VDD1.t4 VP.t5 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=2.12685 ps=13.22 w=12.89 l=0.39
X13 VDD2.t1 VN.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=5.0271 ps=26.56 w=12.89 l=0.39
X14 VDD2.t6 VN.t6 VTAIL.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=0 ps=0 w=12.89 l=0.39
X16 VDD2.t9 VN.t7 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=2.12685 ps=13.22 w=12.89 l=0.39
X17 VDD2.t3 VN.t8 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=2.12685 ps=13.22 w=12.89 l=0.39
X18 VTAIL.t17 VP.t6 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X19 VTAIL.t18 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X20 VTAIL.t6 VN.t9 VDD2.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X21 VDD1.t1 VP.t8 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0271 pd=26.56 as=0 ps=0 w=12.89 l=0.39
X23 VTAIL.t2 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.12685 pd=13.22 as=2.12685 ps=13.22 w=12.89 l=0.39
R0 VN.n2 VN.t8 918.861
R1 VN.n13 VN.t5 918.861
R2 VN.n3 VN.t2 897.88
R3 VN.n1 VN.t3 897.88
R4 VN.n8 VN.t9 897.88
R5 VN.n9 VN.t4 897.88
R6 VN.n14 VN.t0 897.88
R7 VN.n12 VN.t6 897.88
R8 VN.n19 VN.t1 897.88
R9 VN.n20 VN.t7 897.88
R10 VN.n10 VN.n9 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n11 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n8 VN.n0 161.3
R16 VN.n7 VN.n6 161.3
R17 VN.n5 VN.n4 161.3
R18 VN.n16 VN.n13 70.4033
R19 VN.n5 VN.n2 70.4033
R20 VN.n9 VN.n8 48.2005
R21 VN.n20 VN.n19 48.2005
R22 VN VN.n21 42.1766
R23 VN.n4 VN.n3 40.1672
R24 VN.n8 VN.n7 40.1672
R25 VN.n15 VN.n14 40.1672
R26 VN.n19 VN.n18 40.1672
R27 VN.n14 VN.n13 20.9576
R28 VN.n3 VN.n2 20.9576
R29 VN.n4 VN.n1 8.03383
R30 VN.n7 VN.n1 8.03383
R31 VN.n15 VN.n12 8.03383
R32 VN.n18 VN.n12 8.03383
R33 VN.n21 VN.n11 0.189894
R34 VN.n17 VN.n11 0.189894
R35 VN.n17 VN.n16 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n6 VN.n0 0.189894
R38 VN.n10 VN.n0 0.189894
R39 VN VN.n10 0.0516364
R40 VDD2.n137 VDD2.n73 289.615
R41 VDD2.n64 VDD2.n0 289.615
R42 VDD2.n138 VDD2.n137 185
R43 VDD2.n136 VDD2.n135 185
R44 VDD2.n77 VDD2.n76 185
R45 VDD2.n130 VDD2.n129 185
R46 VDD2.n128 VDD2.n127 185
R47 VDD2.n81 VDD2.n80 185
R48 VDD2.n122 VDD2.n121 185
R49 VDD2.n120 VDD2.n119 185
R50 VDD2.n118 VDD2.n84 185
R51 VDD2.n88 VDD2.n85 185
R52 VDD2.n113 VDD2.n112 185
R53 VDD2.n111 VDD2.n110 185
R54 VDD2.n90 VDD2.n89 185
R55 VDD2.n105 VDD2.n104 185
R56 VDD2.n103 VDD2.n102 185
R57 VDD2.n94 VDD2.n93 185
R58 VDD2.n97 VDD2.n96 185
R59 VDD2.n23 VDD2.n22 185
R60 VDD2.n20 VDD2.n19 185
R61 VDD2.n29 VDD2.n28 185
R62 VDD2.n31 VDD2.n30 185
R63 VDD2.n16 VDD2.n15 185
R64 VDD2.n37 VDD2.n36 185
R65 VDD2.n40 VDD2.n39 185
R66 VDD2.n38 VDD2.n12 185
R67 VDD2.n45 VDD2.n11 185
R68 VDD2.n47 VDD2.n46 185
R69 VDD2.n49 VDD2.n48 185
R70 VDD2.n8 VDD2.n7 185
R71 VDD2.n55 VDD2.n54 185
R72 VDD2.n57 VDD2.n56 185
R73 VDD2.n4 VDD2.n3 185
R74 VDD2.n63 VDD2.n62 185
R75 VDD2.n65 VDD2.n64 185
R76 VDD2.t9 VDD2.n95 149.524
R77 VDD2.t3 VDD2.n21 149.524
R78 VDD2.n137 VDD2.n136 104.615
R79 VDD2.n136 VDD2.n76 104.615
R80 VDD2.n129 VDD2.n76 104.615
R81 VDD2.n129 VDD2.n128 104.615
R82 VDD2.n128 VDD2.n80 104.615
R83 VDD2.n121 VDD2.n80 104.615
R84 VDD2.n121 VDD2.n120 104.615
R85 VDD2.n120 VDD2.n84 104.615
R86 VDD2.n88 VDD2.n84 104.615
R87 VDD2.n112 VDD2.n88 104.615
R88 VDD2.n112 VDD2.n111 104.615
R89 VDD2.n111 VDD2.n89 104.615
R90 VDD2.n104 VDD2.n89 104.615
R91 VDD2.n104 VDD2.n103 104.615
R92 VDD2.n103 VDD2.n93 104.615
R93 VDD2.n96 VDD2.n93 104.615
R94 VDD2.n22 VDD2.n19 104.615
R95 VDD2.n29 VDD2.n19 104.615
R96 VDD2.n30 VDD2.n29 104.615
R97 VDD2.n30 VDD2.n15 104.615
R98 VDD2.n37 VDD2.n15 104.615
R99 VDD2.n39 VDD2.n37 104.615
R100 VDD2.n39 VDD2.n38 104.615
R101 VDD2.n38 VDD2.n11 104.615
R102 VDD2.n47 VDD2.n11 104.615
R103 VDD2.n48 VDD2.n47 104.615
R104 VDD2.n48 VDD2.n7 104.615
R105 VDD2.n55 VDD2.n7 104.615
R106 VDD2.n56 VDD2.n55 104.615
R107 VDD2.n56 VDD2.n3 104.615
R108 VDD2.n63 VDD2.n3 104.615
R109 VDD2.n64 VDD2.n63 104.615
R110 VDD2.n72 VDD2.n71 63.0831
R111 VDD2 VDD2.n145 63.0801
R112 VDD2.n144 VDD2.n143 62.673
R113 VDD2.n70 VDD2.n69 62.673
R114 VDD2.n96 VDD2.t9 52.3082
R115 VDD2.n22 VDD2.t3 52.3082
R116 VDD2.n70 VDD2.n68 50.4545
R117 VDD2.n142 VDD2.n141 49.8338
R118 VDD2.n142 VDD2.n72 37.7756
R119 VDD2.n119 VDD2.n118 13.1884
R120 VDD2.n46 VDD2.n45 13.1884
R121 VDD2.n122 VDD2.n83 12.8005
R122 VDD2.n117 VDD2.n85 12.8005
R123 VDD2.n44 VDD2.n12 12.8005
R124 VDD2.n49 VDD2.n10 12.8005
R125 VDD2.n123 VDD2.n81 12.0247
R126 VDD2.n114 VDD2.n113 12.0247
R127 VDD2.n41 VDD2.n40 12.0247
R128 VDD2.n50 VDD2.n8 12.0247
R129 VDD2.n127 VDD2.n126 11.249
R130 VDD2.n110 VDD2.n87 11.249
R131 VDD2.n36 VDD2.n14 11.249
R132 VDD2.n54 VDD2.n53 11.249
R133 VDD2.n130 VDD2.n79 10.4732
R134 VDD2.n109 VDD2.n90 10.4732
R135 VDD2.n35 VDD2.n16 10.4732
R136 VDD2.n57 VDD2.n6 10.4732
R137 VDD2.n97 VDD2.n95 10.2747
R138 VDD2.n23 VDD2.n21 10.2747
R139 VDD2.n131 VDD2.n77 9.69747
R140 VDD2.n106 VDD2.n105 9.69747
R141 VDD2.n32 VDD2.n31 9.69747
R142 VDD2.n58 VDD2.n4 9.69747
R143 VDD2.n141 VDD2.n140 9.45567
R144 VDD2.n68 VDD2.n67 9.45567
R145 VDD2.n99 VDD2.n98 9.3005
R146 VDD2.n101 VDD2.n100 9.3005
R147 VDD2.n92 VDD2.n91 9.3005
R148 VDD2.n107 VDD2.n106 9.3005
R149 VDD2.n109 VDD2.n108 9.3005
R150 VDD2.n87 VDD2.n86 9.3005
R151 VDD2.n115 VDD2.n114 9.3005
R152 VDD2.n117 VDD2.n116 9.3005
R153 VDD2.n140 VDD2.n139 9.3005
R154 VDD2.n75 VDD2.n74 9.3005
R155 VDD2.n134 VDD2.n133 9.3005
R156 VDD2.n132 VDD2.n131 9.3005
R157 VDD2.n79 VDD2.n78 9.3005
R158 VDD2.n126 VDD2.n125 9.3005
R159 VDD2.n124 VDD2.n123 9.3005
R160 VDD2.n83 VDD2.n82 9.3005
R161 VDD2.n2 VDD2.n1 9.3005
R162 VDD2.n61 VDD2.n60 9.3005
R163 VDD2.n59 VDD2.n58 9.3005
R164 VDD2.n6 VDD2.n5 9.3005
R165 VDD2.n53 VDD2.n52 9.3005
R166 VDD2.n51 VDD2.n50 9.3005
R167 VDD2.n10 VDD2.n9 9.3005
R168 VDD2.n25 VDD2.n24 9.3005
R169 VDD2.n27 VDD2.n26 9.3005
R170 VDD2.n18 VDD2.n17 9.3005
R171 VDD2.n33 VDD2.n32 9.3005
R172 VDD2.n35 VDD2.n34 9.3005
R173 VDD2.n14 VDD2.n13 9.3005
R174 VDD2.n42 VDD2.n41 9.3005
R175 VDD2.n44 VDD2.n43 9.3005
R176 VDD2.n67 VDD2.n66 9.3005
R177 VDD2.n135 VDD2.n134 8.92171
R178 VDD2.n102 VDD2.n92 8.92171
R179 VDD2.n28 VDD2.n18 8.92171
R180 VDD2.n62 VDD2.n61 8.92171
R181 VDD2.n138 VDD2.n75 8.14595
R182 VDD2.n101 VDD2.n94 8.14595
R183 VDD2.n27 VDD2.n20 8.14595
R184 VDD2.n65 VDD2.n2 8.14595
R185 VDD2.n139 VDD2.n73 7.3702
R186 VDD2.n98 VDD2.n97 7.3702
R187 VDD2.n24 VDD2.n23 7.3702
R188 VDD2.n66 VDD2.n0 7.3702
R189 VDD2.n141 VDD2.n73 6.59444
R190 VDD2.n68 VDD2.n0 6.59444
R191 VDD2.n139 VDD2.n138 5.81868
R192 VDD2.n98 VDD2.n94 5.81868
R193 VDD2.n24 VDD2.n20 5.81868
R194 VDD2.n66 VDD2.n65 5.81868
R195 VDD2.n135 VDD2.n75 5.04292
R196 VDD2.n102 VDD2.n101 5.04292
R197 VDD2.n28 VDD2.n27 5.04292
R198 VDD2.n62 VDD2.n2 5.04292
R199 VDD2.n134 VDD2.n77 4.26717
R200 VDD2.n105 VDD2.n92 4.26717
R201 VDD2.n31 VDD2.n18 4.26717
R202 VDD2.n61 VDD2.n4 4.26717
R203 VDD2.n131 VDD2.n130 3.49141
R204 VDD2.n106 VDD2.n90 3.49141
R205 VDD2.n32 VDD2.n16 3.49141
R206 VDD2.n58 VDD2.n57 3.49141
R207 VDD2.n99 VDD2.n95 2.84303
R208 VDD2.n25 VDD2.n21 2.84303
R209 VDD2.n127 VDD2.n79 2.71565
R210 VDD2.n110 VDD2.n109 2.71565
R211 VDD2.n36 VDD2.n35 2.71565
R212 VDD2.n54 VDD2.n6 2.71565
R213 VDD2.n126 VDD2.n81 1.93989
R214 VDD2.n113 VDD2.n87 1.93989
R215 VDD2.n40 VDD2.n14 1.93989
R216 VDD2.n53 VDD2.n8 1.93989
R217 VDD2.n145 VDD2.t5 1.53657
R218 VDD2.n145 VDD2.t1 1.53657
R219 VDD2.n143 VDD2.t2 1.53657
R220 VDD2.n143 VDD2.t6 1.53657
R221 VDD2.n71 VDD2.t8 1.53657
R222 VDD2.n71 VDD2.t7 1.53657
R223 VDD2.n69 VDD2.t0 1.53657
R224 VDD2.n69 VDD2.t4 1.53657
R225 VDD2.n123 VDD2.n122 1.16414
R226 VDD2.n114 VDD2.n85 1.16414
R227 VDD2.n41 VDD2.n12 1.16414
R228 VDD2.n50 VDD2.n49 1.16414
R229 VDD2.n144 VDD2.n142 0.62119
R230 VDD2.n119 VDD2.n83 0.388379
R231 VDD2.n118 VDD2.n117 0.388379
R232 VDD2.n45 VDD2.n44 0.388379
R233 VDD2.n46 VDD2.n10 0.388379
R234 VDD2 VDD2.n144 0.213862
R235 VDD2.n140 VDD2.n74 0.155672
R236 VDD2.n133 VDD2.n74 0.155672
R237 VDD2.n133 VDD2.n132 0.155672
R238 VDD2.n132 VDD2.n78 0.155672
R239 VDD2.n125 VDD2.n78 0.155672
R240 VDD2.n125 VDD2.n124 0.155672
R241 VDD2.n124 VDD2.n82 0.155672
R242 VDD2.n116 VDD2.n82 0.155672
R243 VDD2.n116 VDD2.n115 0.155672
R244 VDD2.n115 VDD2.n86 0.155672
R245 VDD2.n108 VDD2.n86 0.155672
R246 VDD2.n108 VDD2.n107 0.155672
R247 VDD2.n107 VDD2.n91 0.155672
R248 VDD2.n100 VDD2.n91 0.155672
R249 VDD2.n100 VDD2.n99 0.155672
R250 VDD2.n26 VDD2.n25 0.155672
R251 VDD2.n26 VDD2.n17 0.155672
R252 VDD2.n33 VDD2.n17 0.155672
R253 VDD2.n34 VDD2.n33 0.155672
R254 VDD2.n34 VDD2.n13 0.155672
R255 VDD2.n42 VDD2.n13 0.155672
R256 VDD2.n43 VDD2.n42 0.155672
R257 VDD2.n43 VDD2.n9 0.155672
R258 VDD2.n51 VDD2.n9 0.155672
R259 VDD2.n52 VDD2.n51 0.155672
R260 VDD2.n52 VDD2.n5 0.155672
R261 VDD2.n59 VDD2.n5 0.155672
R262 VDD2.n60 VDD2.n59 0.155672
R263 VDD2.n60 VDD2.n1 0.155672
R264 VDD2.n67 VDD2.n1 0.155672
R265 VDD2.n72 VDD2.n70 0.100326
R266 VTAIL.n288 VTAIL.n224 289.615
R267 VTAIL.n66 VTAIL.n2 289.615
R268 VTAIL.n218 VTAIL.n154 289.615
R269 VTAIL.n144 VTAIL.n80 289.615
R270 VTAIL.n247 VTAIL.n246 185
R271 VTAIL.n244 VTAIL.n243 185
R272 VTAIL.n253 VTAIL.n252 185
R273 VTAIL.n255 VTAIL.n254 185
R274 VTAIL.n240 VTAIL.n239 185
R275 VTAIL.n261 VTAIL.n260 185
R276 VTAIL.n264 VTAIL.n263 185
R277 VTAIL.n262 VTAIL.n236 185
R278 VTAIL.n269 VTAIL.n235 185
R279 VTAIL.n271 VTAIL.n270 185
R280 VTAIL.n273 VTAIL.n272 185
R281 VTAIL.n232 VTAIL.n231 185
R282 VTAIL.n279 VTAIL.n278 185
R283 VTAIL.n281 VTAIL.n280 185
R284 VTAIL.n228 VTAIL.n227 185
R285 VTAIL.n287 VTAIL.n286 185
R286 VTAIL.n289 VTAIL.n288 185
R287 VTAIL.n25 VTAIL.n24 185
R288 VTAIL.n22 VTAIL.n21 185
R289 VTAIL.n31 VTAIL.n30 185
R290 VTAIL.n33 VTAIL.n32 185
R291 VTAIL.n18 VTAIL.n17 185
R292 VTAIL.n39 VTAIL.n38 185
R293 VTAIL.n42 VTAIL.n41 185
R294 VTAIL.n40 VTAIL.n14 185
R295 VTAIL.n47 VTAIL.n13 185
R296 VTAIL.n49 VTAIL.n48 185
R297 VTAIL.n51 VTAIL.n50 185
R298 VTAIL.n10 VTAIL.n9 185
R299 VTAIL.n57 VTAIL.n56 185
R300 VTAIL.n59 VTAIL.n58 185
R301 VTAIL.n6 VTAIL.n5 185
R302 VTAIL.n65 VTAIL.n64 185
R303 VTAIL.n67 VTAIL.n66 185
R304 VTAIL.n219 VTAIL.n218 185
R305 VTAIL.n217 VTAIL.n216 185
R306 VTAIL.n158 VTAIL.n157 185
R307 VTAIL.n211 VTAIL.n210 185
R308 VTAIL.n209 VTAIL.n208 185
R309 VTAIL.n162 VTAIL.n161 185
R310 VTAIL.n203 VTAIL.n202 185
R311 VTAIL.n201 VTAIL.n200 185
R312 VTAIL.n199 VTAIL.n165 185
R313 VTAIL.n169 VTAIL.n166 185
R314 VTAIL.n194 VTAIL.n193 185
R315 VTAIL.n192 VTAIL.n191 185
R316 VTAIL.n171 VTAIL.n170 185
R317 VTAIL.n186 VTAIL.n185 185
R318 VTAIL.n184 VTAIL.n183 185
R319 VTAIL.n175 VTAIL.n174 185
R320 VTAIL.n178 VTAIL.n177 185
R321 VTAIL.n145 VTAIL.n144 185
R322 VTAIL.n143 VTAIL.n142 185
R323 VTAIL.n84 VTAIL.n83 185
R324 VTAIL.n137 VTAIL.n136 185
R325 VTAIL.n135 VTAIL.n134 185
R326 VTAIL.n88 VTAIL.n87 185
R327 VTAIL.n129 VTAIL.n128 185
R328 VTAIL.n127 VTAIL.n126 185
R329 VTAIL.n125 VTAIL.n91 185
R330 VTAIL.n95 VTAIL.n92 185
R331 VTAIL.n120 VTAIL.n119 185
R332 VTAIL.n118 VTAIL.n117 185
R333 VTAIL.n97 VTAIL.n96 185
R334 VTAIL.n112 VTAIL.n111 185
R335 VTAIL.n110 VTAIL.n109 185
R336 VTAIL.n101 VTAIL.n100 185
R337 VTAIL.n104 VTAIL.n103 185
R338 VTAIL.t11 VTAIL.n245 149.524
R339 VTAIL.t5 VTAIL.n23 149.524
R340 VTAIL.t0 VTAIL.n176 149.524
R341 VTAIL.t10 VTAIL.n102 149.524
R342 VTAIL.n246 VTAIL.n243 104.615
R343 VTAIL.n253 VTAIL.n243 104.615
R344 VTAIL.n254 VTAIL.n253 104.615
R345 VTAIL.n254 VTAIL.n239 104.615
R346 VTAIL.n261 VTAIL.n239 104.615
R347 VTAIL.n263 VTAIL.n261 104.615
R348 VTAIL.n263 VTAIL.n262 104.615
R349 VTAIL.n262 VTAIL.n235 104.615
R350 VTAIL.n271 VTAIL.n235 104.615
R351 VTAIL.n272 VTAIL.n271 104.615
R352 VTAIL.n272 VTAIL.n231 104.615
R353 VTAIL.n279 VTAIL.n231 104.615
R354 VTAIL.n280 VTAIL.n279 104.615
R355 VTAIL.n280 VTAIL.n227 104.615
R356 VTAIL.n287 VTAIL.n227 104.615
R357 VTAIL.n288 VTAIL.n287 104.615
R358 VTAIL.n24 VTAIL.n21 104.615
R359 VTAIL.n31 VTAIL.n21 104.615
R360 VTAIL.n32 VTAIL.n31 104.615
R361 VTAIL.n32 VTAIL.n17 104.615
R362 VTAIL.n39 VTAIL.n17 104.615
R363 VTAIL.n41 VTAIL.n39 104.615
R364 VTAIL.n41 VTAIL.n40 104.615
R365 VTAIL.n40 VTAIL.n13 104.615
R366 VTAIL.n49 VTAIL.n13 104.615
R367 VTAIL.n50 VTAIL.n49 104.615
R368 VTAIL.n50 VTAIL.n9 104.615
R369 VTAIL.n57 VTAIL.n9 104.615
R370 VTAIL.n58 VTAIL.n57 104.615
R371 VTAIL.n58 VTAIL.n5 104.615
R372 VTAIL.n65 VTAIL.n5 104.615
R373 VTAIL.n66 VTAIL.n65 104.615
R374 VTAIL.n218 VTAIL.n217 104.615
R375 VTAIL.n217 VTAIL.n157 104.615
R376 VTAIL.n210 VTAIL.n157 104.615
R377 VTAIL.n210 VTAIL.n209 104.615
R378 VTAIL.n209 VTAIL.n161 104.615
R379 VTAIL.n202 VTAIL.n161 104.615
R380 VTAIL.n202 VTAIL.n201 104.615
R381 VTAIL.n201 VTAIL.n165 104.615
R382 VTAIL.n169 VTAIL.n165 104.615
R383 VTAIL.n193 VTAIL.n169 104.615
R384 VTAIL.n193 VTAIL.n192 104.615
R385 VTAIL.n192 VTAIL.n170 104.615
R386 VTAIL.n185 VTAIL.n170 104.615
R387 VTAIL.n185 VTAIL.n184 104.615
R388 VTAIL.n184 VTAIL.n174 104.615
R389 VTAIL.n177 VTAIL.n174 104.615
R390 VTAIL.n144 VTAIL.n143 104.615
R391 VTAIL.n143 VTAIL.n83 104.615
R392 VTAIL.n136 VTAIL.n83 104.615
R393 VTAIL.n136 VTAIL.n135 104.615
R394 VTAIL.n135 VTAIL.n87 104.615
R395 VTAIL.n128 VTAIL.n87 104.615
R396 VTAIL.n128 VTAIL.n127 104.615
R397 VTAIL.n127 VTAIL.n91 104.615
R398 VTAIL.n95 VTAIL.n91 104.615
R399 VTAIL.n119 VTAIL.n95 104.615
R400 VTAIL.n119 VTAIL.n118 104.615
R401 VTAIL.n118 VTAIL.n96 104.615
R402 VTAIL.n111 VTAIL.n96 104.615
R403 VTAIL.n111 VTAIL.n110 104.615
R404 VTAIL.n110 VTAIL.n100 104.615
R405 VTAIL.n103 VTAIL.n100 104.615
R406 VTAIL.n246 VTAIL.t11 52.3082
R407 VTAIL.n24 VTAIL.t5 52.3082
R408 VTAIL.n177 VTAIL.t0 52.3082
R409 VTAIL.n103 VTAIL.t10 52.3082
R410 VTAIL.n295 VTAIL.n294 45.9942
R411 VTAIL.n1 VTAIL.n0 45.9942
R412 VTAIL.n73 VTAIL.n72 45.9942
R413 VTAIL.n75 VTAIL.n74 45.9942
R414 VTAIL.n153 VTAIL.n152 45.9942
R415 VTAIL.n151 VTAIL.n150 45.9942
R416 VTAIL.n79 VTAIL.n78 45.9942
R417 VTAIL.n77 VTAIL.n76 45.9942
R418 VTAIL.n293 VTAIL.n292 33.155
R419 VTAIL.n71 VTAIL.n70 33.155
R420 VTAIL.n223 VTAIL.n222 33.155
R421 VTAIL.n149 VTAIL.n148 33.155
R422 VTAIL.n77 VTAIL.n75 24.7203
R423 VTAIL.n293 VTAIL.n223 24.0996
R424 VTAIL.n270 VTAIL.n269 13.1884
R425 VTAIL.n48 VTAIL.n47 13.1884
R426 VTAIL.n200 VTAIL.n199 13.1884
R427 VTAIL.n126 VTAIL.n125 13.1884
R428 VTAIL.n268 VTAIL.n236 12.8005
R429 VTAIL.n273 VTAIL.n234 12.8005
R430 VTAIL.n46 VTAIL.n14 12.8005
R431 VTAIL.n51 VTAIL.n12 12.8005
R432 VTAIL.n203 VTAIL.n164 12.8005
R433 VTAIL.n198 VTAIL.n166 12.8005
R434 VTAIL.n129 VTAIL.n90 12.8005
R435 VTAIL.n124 VTAIL.n92 12.8005
R436 VTAIL.n265 VTAIL.n264 12.0247
R437 VTAIL.n274 VTAIL.n232 12.0247
R438 VTAIL.n43 VTAIL.n42 12.0247
R439 VTAIL.n52 VTAIL.n10 12.0247
R440 VTAIL.n204 VTAIL.n162 12.0247
R441 VTAIL.n195 VTAIL.n194 12.0247
R442 VTAIL.n130 VTAIL.n88 12.0247
R443 VTAIL.n121 VTAIL.n120 12.0247
R444 VTAIL.n260 VTAIL.n238 11.249
R445 VTAIL.n278 VTAIL.n277 11.249
R446 VTAIL.n38 VTAIL.n16 11.249
R447 VTAIL.n56 VTAIL.n55 11.249
R448 VTAIL.n208 VTAIL.n207 11.249
R449 VTAIL.n191 VTAIL.n168 11.249
R450 VTAIL.n134 VTAIL.n133 11.249
R451 VTAIL.n117 VTAIL.n94 11.249
R452 VTAIL.n259 VTAIL.n240 10.4732
R453 VTAIL.n281 VTAIL.n230 10.4732
R454 VTAIL.n37 VTAIL.n18 10.4732
R455 VTAIL.n59 VTAIL.n8 10.4732
R456 VTAIL.n211 VTAIL.n160 10.4732
R457 VTAIL.n190 VTAIL.n171 10.4732
R458 VTAIL.n137 VTAIL.n86 10.4732
R459 VTAIL.n116 VTAIL.n97 10.4732
R460 VTAIL.n247 VTAIL.n245 10.2747
R461 VTAIL.n25 VTAIL.n23 10.2747
R462 VTAIL.n178 VTAIL.n176 10.2747
R463 VTAIL.n104 VTAIL.n102 10.2747
R464 VTAIL.n256 VTAIL.n255 9.69747
R465 VTAIL.n282 VTAIL.n228 9.69747
R466 VTAIL.n34 VTAIL.n33 9.69747
R467 VTAIL.n60 VTAIL.n6 9.69747
R468 VTAIL.n212 VTAIL.n158 9.69747
R469 VTAIL.n187 VTAIL.n186 9.69747
R470 VTAIL.n138 VTAIL.n84 9.69747
R471 VTAIL.n113 VTAIL.n112 9.69747
R472 VTAIL.n292 VTAIL.n291 9.45567
R473 VTAIL.n70 VTAIL.n69 9.45567
R474 VTAIL.n222 VTAIL.n221 9.45567
R475 VTAIL.n148 VTAIL.n147 9.45567
R476 VTAIL.n226 VTAIL.n225 9.3005
R477 VTAIL.n285 VTAIL.n284 9.3005
R478 VTAIL.n283 VTAIL.n282 9.3005
R479 VTAIL.n230 VTAIL.n229 9.3005
R480 VTAIL.n277 VTAIL.n276 9.3005
R481 VTAIL.n275 VTAIL.n274 9.3005
R482 VTAIL.n234 VTAIL.n233 9.3005
R483 VTAIL.n249 VTAIL.n248 9.3005
R484 VTAIL.n251 VTAIL.n250 9.3005
R485 VTAIL.n242 VTAIL.n241 9.3005
R486 VTAIL.n257 VTAIL.n256 9.3005
R487 VTAIL.n259 VTAIL.n258 9.3005
R488 VTAIL.n238 VTAIL.n237 9.3005
R489 VTAIL.n266 VTAIL.n265 9.3005
R490 VTAIL.n268 VTAIL.n267 9.3005
R491 VTAIL.n291 VTAIL.n290 9.3005
R492 VTAIL.n4 VTAIL.n3 9.3005
R493 VTAIL.n63 VTAIL.n62 9.3005
R494 VTAIL.n61 VTAIL.n60 9.3005
R495 VTAIL.n8 VTAIL.n7 9.3005
R496 VTAIL.n55 VTAIL.n54 9.3005
R497 VTAIL.n53 VTAIL.n52 9.3005
R498 VTAIL.n12 VTAIL.n11 9.3005
R499 VTAIL.n27 VTAIL.n26 9.3005
R500 VTAIL.n29 VTAIL.n28 9.3005
R501 VTAIL.n20 VTAIL.n19 9.3005
R502 VTAIL.n35 VTAIL.n34 9.3005
R503 VTAIL.n37 VTAIL.n36 9.3005
R504 VTAIL.n16 VTAIL.n15 9.3005
R505 VTAIL.n44 VTAIL.n43 9.3005
R506 VTAIL.n46 VTAIL.n45 9.3005
R507 VTAIL.n69 VTAIL.n68 9.3005
R508 VTAIL.n180 VTAIL.n179 9.3005
R509 VTAIL.n182 VTAIL.n181 9.3005
R510 VTAIL.n173 VTAIL.n172 9.3005
R511 VTAIL.n188 VTAIL.n187 9.3005
R512 VTAIL.n190 VTAIL.n189 9.3005
R513 VTAIL.n168 VTAIL.n167 9.3005
R514 VTAIL.n196 VTAIL.n195 9.3005
R515 VTAIL.n198 VTAIL.n197 9.3005
R516 VTAIL.n221 VTAIL.n220 9.3005
R517 VTAIL.n156 VTAIL.n155 9.3005
R518 VTAIL.n215 VTAIL.n214 9.3005
R519 VTAIL.n213 VTAIL.n212 9.3005
R520 VTAIL.n160 VTAIL.n159 9.3005
R521 VTAIL.n207 VTAIL.n206 9.3005
R522 VTAIL.n205 VTAIL.n204 9.3005
R523 VTAIL.n164 VTAIL.n163 9.3005
R524 VTAIL.n106 VTAIL.n105 9.3005
R525 VTAIL.n108 VTAIL.n107 9.3005
R526 VTAIL.n99 VTAIL.n98 9.3005
R527 VTAIL.n114 VTAIL.n113 9.3005
R528 VTAIL.n116 VTAIL.n115 9.3005
R529 VTAIL.n94 VTAIL.n93 9.3005
R530 VTAIL.n122 VTAIL.n121 9.3005
R531 VTAIL.n124 VTAIL.n123 9.3005
R532 VTAIL.n147 VTAIL.n146 9.3005
R533 VTAIL.n82 VTAIL.n81 9.3005
R534 VTAIL.n141 VTAIL.n140 9.3005
R535 VTAIL.n139 VTAIL.n138 9.3005
R536 VTAIL.n86 VTAIL.n85 9.3005
R537 VTAIL.n133 VTAIL.n132 9.3005
R538 VTAIL.n131 VTAIL.n130 9.3005
R539 VTAIL.n90 VTAIL.n89 9.3005
R540 VTAIL.n252 VTAIL.n242 8.92171
R541 VTAIL.n286 VTAIL.n285 8.92171
R542 VTAIL.n30 VTAIL.n20 8.92171
R543 VTAIL.n64 VTAIL.n63 8.92171
R544 VTAIL.n216 VTAIL.n215 8.92171
R545 VTAIL.n183 VTAIL.n173 8.92171
R546 VTAIL.n142 VTAIL.n141 8.92171
R547 VTAIL.n109 VTAIL.n99 8.92171
R548 VTAIL.n251 VTAIL.n244 8.14595
R549 VTAIL.n289 VTAIL.n226 8.14595
R550 VTAIL.n29 VTAIL.n22 8.14595
R551 VTAIL.n67 VTAIL.n4 8.14595
R552 VTAIL.n219 VTAIL.n156 8.14595
R553 VTAIL.n182 VTAIL.n175 8.14595
R554 VTAIL.n145 VTAIL.n82 8.14595
R555 VTAIL.n108 VTAIL.n101 8.14595
R556 VTAIL.n248 VTAIL.n247 7.3702
R557 VTAIL.n290 VTAIL.n224 7.3702
R558 VTAIL.n26 VTAIL.n25 7.3702
R559 VTAIL.n68 VTAIL.n2 7.3702
R560 VTAIL.n220 VTAIL.n154 7.3702
R561 VTAIL.n179 VTAIL.n178 7.3702
R562 VTAIL.n146 VTAIL.n80 7.3702
R563 VTAIL.n105 VTAIL.n104 7.3702
R564 VTAIL.n292 VTAIL.n224 6.59444
R565 VTAIL.n70 VTAIL.n2 6.59444
R566 VTAIL.n222 VTAIL.n154 6.59444
R567 VTAIL.n148 VTAIL.n80 6.59444
R568 VTAIL.n248 VTAIL.n244 5.81868
R569 VTAIL.n290 VTAIL.n289 5.81868
R570 VTAIL.n26 VTAIL.n22 5.81868
R571 VTAIL.n68 VTAIL.n67 5.81868
R572 VTAIL.n220 VTAIL.n219 5.81868
R573 VTAIL.n179 VTAIL.n175 5.81868
R574 VTAIL.n146 VTAIL.n145 5.81868
R575 VTAIL.n105 VTAIL.n101 5.81868
R576 VTAIL.n252 VTAIL.n251 5.04292
R577 VTAIL.n286 VTAIL.n226 5.04292
R578 VTAIL.n30 VTAIL.n29 5.04292
R579 VTAIL.n64 VTAIL.n4 5.04292
R580 VTAIL.n216 VTAIL.n156 5.04292
R581 VTAIL.n183 VTAIL.n182 5.04292
R582 VTAIL.n142 VTAIL.n82 5.04292
R583 VTAIL.n109 VTAIL.n108 5.04292
R584 VTAIL.n255 VTAIL.n242 4.26717
R585 VTAIL.n285 VTAIL.n228 4.26717
R586 VTAIL.n33 VTAIL.n20 4.26717
R587 VTAIL.n63 VTAIL.n6 4.26717
R588 VTAIL.n215 VTAIL.n158 4.26717
R589 VTAIL.n186 VTAIL.n173 4.26717
R590 VTAIL.n141 VTAIL.n84 4.26717
R591 VTAIL.n112 VTAIL.n99 4.26717
R592 VTAIL.n256 VTAIL.n240 3.49141
R593 VTAIL.n282 VTAIL.n281 3.49141
R594 VTAIL.n34 VTAIL.n18 3.49141
R595 VTAIL.n60 VTAIL.n59 3.49141
R596 VTAIL.n212 VTAIL.n211 3.49141
R597 VTAIL.n187 VTAIL.n171 3.49141
R598 VTAIL.n138 VTAIL.n137 3.49141
R599 VTAIL.n113 VTAIL.n97 3.49141
R600 VTAIL.n249 VTAIL.n245 2.84303
R601 VTAIL.n27 VTAIL.n23 2.84303
R602 VTAIL.n180 VTAIL.n176 2.84303
R603 VTAIL.n106 VTAIL.n102 2.84303
R604 VTAIL.n260 VTAIL.n259 2.71565
R605 VTAIL.n278 VTAIL.n230 2.71565
R606 VTAIL.n38 VTAIL.n37 2.71565
R607 VTAIL.n56 VTAIL.n8 2.71565
R608 VTAIL.n208 VTAIL.n160 2.71565
R609 VTAIL.n191 VTAIL.n190 2.71565
R610 VTAIL.n134 VTAIL.n86 2.71565
R611 VTAIL.n117 VTAIL.n116 2.71565
R612 VTAIL.n264 VTAIL.n238 1.93989
R613 VTAIL.n277 VTAIL.n232 1.93989
R614 VTAIL.n42 VTAIL.n16 1.93989
R615 VTAIL.n55 VTAIL.n10 1.93989
R616 VTAIL.n207 VTAIL.n162 1.93989
R617 VTAIL.n194 VTAIL.n168 1.93989
R618 VTAIL.n133 VTAIL.n88 1.93989
R619 VTAIL.n120 VTAIL.n94 1.93989
R620 VTAIL.n294 VTAIL.t12 1.53657
R621 VTAIL.n294 VTAIL.t6 1.53657
R622 VTAIL.n0 VTAIL.t7 1.53657
R623 VTAIL.n0 VTAIL.t13 1.53657
R624 VTAIL.n72 VTAIL.t19 1.53657
R625 VTAIL.n72 VTAIL.t2 1.53657
R626 VTAIL.n74 VTAIL.t16 1.53657
R627 VTAIL.n74 VTAIL.t3 1.53657
R628 VTAIL.n152 VTAIL.t1 1.53657
R629 VTAIL.n152 VTAIL.t17 1.53657
R630 VTAIL.n150 VTAIL.t4 1.53657
R631 VTAIL.n150 VTAIL.t18 1.53657
R632 VTAIL.n78 VTAIL.t9 1.53657
R633 VTAIL.n78 VTAIL.t15 1.53657
R634 VTAIL.n76 VTAIL.t8 1.53657
R635 VTAIL.n76 VTAIL.t14 1.53657
R636 VTAIL.n265 VTAIL.n236 1.16414
R637 VTAIL.n274 VTAIL.n273 1.16414
R638 VTAIL.n43 VTAIL.n14 1.16414
R639 VTAIL.n52 VTAIL.n51 1.16414
R640 VTAIL.n204 VTAIL.n203 1.16414
R641 VTAIL.n195 VTAIL.n166 1.16414
R642 VTAIL.n130 VTAIL.n129 1.16414
R643 VTAIL.n121 VTAIL.n92 1.16414
R644 VTAIL.n151 VTAIL.n149 0.780672
R645 VTAIL.n71 VTAIL.n1 0.780672
R646 VTAIL.n79 VTAIL.n77 0.62119
R647 VTAIL.n149 VTAIL.n79 0.62119
R648 VTAIL.n153 VTAIL.n151 0.62119
R649 VTAIL.n223 VTAIL.n153 0.62119
R650 VTAIL.n75 VTAIL.n73 0.62119
R651 VTAIL.n73 VTAIL.n71 0.62119
R652 VTAIL.n295 VTAIL.n293 0.62119
R653 VTAIL VTAIL.n1 0.524207
R654 VTAIL.n269 VTAIL.n268 0.388379
R655 VTAIL.n270 VTAIL.n234 0.388379
R656 VTAIL.n47 VTAIL.n46 0.388379
R657 VTAIL.n48 VTAIL.n12 0.388379
R658 VTAIL.n200 VTAIL.n164 0.388379
R659 VTAIL.n199 VTAIL.n198 0.388379
R660 VTAIL.n126 VTAIL.n90 0.388379
R661 VTAIL.n125 VTAIL.n124 0.388379
R662 VTAIL.n250 VTAIL.n249 0.155672
R663 VTAIL.n250 VTAIL.n241 0.155672
R664 VTAIL.n257 VTAIL.n241 0.155672
R665 VTAIL.n258 VTAIL.n257 0.155672
R666 VTAIL.n258 VTAIL.n237 0.155672
R667 VTAIL.n266 VTAIL.n237 0.155672
R668 VTAIL.n267 VTAIL.n266 0.155672
R669 VTAIL.n267 VTAIL.n233 0.155672
R670 VTAIL.n275 VTAIL.n233 0.155672
R671 VTAIL.n276 VTAIL.n275 0.155672
R672 VTAIL.n276 VTAIL.n229 0.155672
R673 VTAIL.n283 VTAIL.n229 0.155672
R674 VTAIL.n284 VTAIL.n283 0.155672
R675 VTAIL.n284 VTAIL.n225 0.155672
R676 VTAIL.n291 VTAIL.n225 0.155672
R677 VTAIL.n28 VTAIL.n27 0.155672
R678 VTAIL.n28 VTAIL.n19 0.155672
R679 VTAIL.n35 VTAIL.n19 0.155672
R680 VTAIL.n36 VTAIL.n35 0.155672
R681 VTAIL.n36 VTAIL.n15 0.155672
R682 VTAIL.n44 VTAIL.n15 0.155672
R683 VTAIL.n45 VTAIL.n44 0.155672
R684 VTAIL.n45 VTAIL.n11 0.155672
R685 VTAIL.n53 VTAIL.n11 0.155672
R686 VTAIL.n54 VTAIL.n53 0.155672
R687 VTAIL.n54 VTAIL.n7 0.155672
R688 VTAIL.n61 VTAIL.n7 0.155672
R689 VTAIL.n62 VTAIL.n61 0.155672
R690 VTAIL.n62 VTAIL.n3 0.155672
R691 VTAIL.n69 VTAIL.n3 0.155672
R692 VTAIL.n221 VTAIL.n155 0.155672
R693 VTAIL.n214 VTAIL.n155 0.155672
R694 VTAIL.n214 VTAIL.n213 0.155672
R695 VTAIL.n213 VTAIL.n159 0.155672
R696 VTAIL.n206 VTAIL.n159 0.155672
R697 VTAIL.n206 VTAIL.n205 0.155672
R698 VTAIL.n205 VTAIL.n163 0.155672
R699 VTAIL.n197 VTAIL.n163 0.155672
R700 VTAIL.n197 VTAIL.n196 0.155672
R701 VTAIL.n196 VTAIL.n167 0.155672
R702 VTAIL.n189 VTAIL.n167 0.155672
R703 VTAIL.n189 VTAIL.n188 0.155672
R704 VTAIL.n188 VTAIL.n172 0.155672
R705 VTAIL.n181 VTAIL.n172 0.155672
R706 VTAIL.n181 VTAIL.n180 0.155672
R707 VTAIL.n147 VTAIL.n81 0.155672
R708 VTAIL.n140 VTAIL.n81 0.155672
R709 VTAIL.n140 VTAIL.n139 0.155672
R710 VTAIL.n139 VTAIL.n85 0.155672
R711 VTAIL.n132 VTAIL.n85 0.155672
R712 VTAIL.n132 VTAIL.n131 0.155672
R713 VTAIL.n131 VTAIL.n89 0.155672
R714 VTAIL.n123 VTAIL.n89 0.155672
R715 VTAIL.n123 VTAIL.n122 0.155672
R716 VTAIL.n122 VTAIL.n93 0.155672
R717 VTAIL.n115 VTAIL.n93 0.155672
R718 VTAIL.n115 VTAIL.n114 0.155672
R719 VTAIL.n114 VTAIL.n98 0.155672
R720 VTAIL.n107 VTAIL.n98 0.155672
R721 VTAIL.n107 VTAIL.n106 0.155672
R722 VTAIL VTAIL.n295 0.0974828
R723 B.n381 B.t10 1006.34
R724 B.n379 B.t14 1006.34
R725 B.n94 B.t21 1006.34
R726 B.n91 B.t17 1006.34
R727 B.n671 B.n670 585
R728 B.n289 B.n90 585
R729 B.n288 B.n287 585
R730 B.n286 B.n285 585
R731 B.n284 B.n283 585
R732 B.n282 B.n281 585
R733 B.n280 B.n279 585
R734 B.n278 B.n277 585
R735 B.n276 B.n275 585
R736 B.n274 B.n273 585
R737 B.n272 B.n271 585
R738 B.n270 B.n269 585
R739 B.n268 B.n267 585
R740 B.n266 B.n265 585
R741 B.n264 B.n263 585
R742 B.n262 B.n261 585
R743 B.n260 B.n259 585
R744 B.n258 B.n257 585
R745 B.n256 B.n255 585
R746 B.n254 B.n253 585
R747 B.n252 B.n251 585
R748 B.n250 B.n249 585
R749 B.n248 B.n247 585
R750 B.n246 B.n245 585
R751 B.n244 B.n243 585
R752 B.n242 B.n241 585
R753 B.n240 B.n239 585
R754 B.n238 B.n237 585
R755 B.n236 B.n235 585
R756 B.n234 B.n233 585
R757 B.n232 B.n231 585
R758 B.n230 B.n229 585
R759 B.n228 B.n227 585
R760 B.n226 B.n225 585
R761 B.n224 B.n223 585
R762 B.n222 B.n221 585
R763 B.n220 B.n219 585
R764 B.n218 B.n217 585
R765 B.n216 B.n215 585
R766 B.n214 B.n213 585
R767 B.n212 B.n211 585
R768 B.n210 B.n209 585
R769 B.n208 B.n207 585
R770 B.n206 B.n205 585
R771 B.n204 B.n203 585
R772 B.n202 B.n201 585
R773 B.n200 B.n199 585
R774 B.n198 B.n197 585
R775 B.n196 B.n195 585
R776 B.n194 B.n193 585
R777 B.n192 B.n191 585
R778 B.n190 B.n189 585
R779 B.n188 B.n187 585
R780 B.n186 B.n185 585
R781 B.n184 B.n183 585
R782 B.n182 B.n181 585
R783 B.n180 B.n179 585
R784 B.n178 B.n177 585
R785 B.n176 B.n175 585
R786 B.n174 B.n173 585
R787 B.n172 B.n171 585
R788 B.n170 B.n169 585
R789 B.n168 B.n167 585
R790 B.n166 B.n165 585
R791 B.n164 B.n163 585
R792 B.n162 B.n161 585
R793 B.n160 B.n159 585
R794 B.n158 B.n157 585
R795 B.n156 B.n155 585
R796 B.n154 B.n153 585
R797 B.n152 B.n151 585
R798 B.n150 B.n149 585
R799 B.n148 B.n147 585
R800 B.n146 B.n145 585
R801 B.n144 B.n143 585
R802 B.n142 B.n141 585
R803 B.n140 B.n139 585
R804 B.n138 B.n137 585
R805 B.n136 B.n135 585
R806 B.n134 B.n133 585
R807 B.n132 B.n131 585
R808 B.n130 B.n129 585
R809 B.n128 B.n127 585
R810 B.n126 B.n125 585
R811 B.n124 B.n123 585
R812 B.n122 B.n121 585
R813 B.n120 B.n119 585
R814 B.n118 B.n117 585
R815 B.n116 B.n115 585
R816 B.n114 B.n113 585
R817 B.n112 B.n111 585
R818 B.n110 B.n109 585
R819 B.n108 B.n107 585
R820 B.n106 B.n105 585
R821 B.n104 B.n103 585
R822 B.n102 B.n101 585
R823 B.n100 B.n99 585
R824 B.n98 B.n97 585
R825 B.n669 B.n41 585
R826 B.n674 B.n41 585
R827 B.n668 B.n40 585
R828 B.n675 B.n40 585
R829 B.n667 B.n666 585
R830 B.n666 B.n36 585
R831 B.n665 B.n35 585
R832 B.n681 B.n35 585
R833 B.n664 B.n34 585
R834 B.n682 B.n34 585
R835 B.n663 B.n33 585
R836 B.n683 B.n33 585
R837 B.n662 B.n661 585
R838 B.n661 B.n29 585
R839 B.n660 B.n28 585
R840 B.n689 B.n28 585
R841 B.n659 B.n27 585
R842 B.n690 B.n27 585
R843 B.n658 B.n26 585
R844 B.n691 B.n26 585
R845 B.n657 B.n656 585
R846 B.n656 B.n22 585
R847 B.n655 B.n21 585
R848 B.n697 B.n21 585
R849 B.n654 B.n20 585
R850 B.n698 B.n20 585
R851 B.n653 B.n19 585
R852 B.n699 B.n19 585
R853 B.n652 B.n651 585
R854 B.n651 B.n18 585
R855 B.n650 B.n14 585
R856 B.n705 B.n14 585
R857 B.n649 B.n13 585
R858 B.n706 B.n13 585
R859 B.n648 B.n12 585
R860 B.n707 B.n12 585
R861 B.n647 B.n646 585
R862 B.n646 B.n11 585
R863 B.n645 B.n7 585
R864 B.n713 B.n7 585
R865 B.n644 B.n6 585
R866 B.n714 B.n6 585
R867 B.n643 B.n5 585
R868 B.n715 B.n5 585
R869 B.n642 B.n641 585
R870 B.n641 B.n4 585
R871 B.n640 B.n290 585
R872 B.n640 B.n639 585
R873 B.n629 B.n291 585
R874 B.n632 B.n291 585
R875 B.n631 B.n630 585
R876 B.n633 B.n631 585
R877 B.n628 B.n295 585
R878 B.n298 B.n295 585
R879 B.n627 B.n626 585
R880 B.n626 B.n625 585
R881 B.n297 B.n296 585
R882 B.n618 B.n297 585
R883 B.n617 B.n616 585
R884 B.n619 B.n617 585
R885 B.n615 B.n303 585
R886 B.n303 B.n302 585
R887 B.n614 B.n613 585
R888 B.n613 B.n612 585
R889 B.n305 B.n304 585
R890 B.n306 B.n305 585
R891 B.n605 B.n604 585
R892 B.n606 B.n605 585
R893 B.n603 B.n311 585
R894 B.n311 B.n310 585
R895 B.n602 B.n601 585
R896 B.n601 B.n600 585
R897 B.n313 B.n312 585
R898 B.n314 B.n313 585
R899 B.n593 B.n592 585
R900 B.n594 B.n593 585
R901 B.n591 B.n318 585
R902 B.n322 B.n318 585
R903 B.n590 B.n589 585
R904 B.n589 B.n588 585
R905 B.n320 B.n319 585
R906 B.n321 B.n320 585
R907 B.n581 B.n580 585
R908 B.n582 B.n581 585
R909 B.n579 B.n327 585
R910 B.n327 B.n326 585
R911 B.n574 B.n573 585
R912 B.n572 B.n378 585
R913 B.n571 B.n377 585
R914 B.n576 B.n377 585
R915 B.n570 B.n569 585
R916 B.n568 B.n567 585
R917 B.n566 B.n565 585
R918 B.n564 B.n563 585
R919 B.n562 B.n561 585
R920 B.n560 B.n559 585
R921 B.n558 B.n557 585
R922 B.n556 B.n555 585
R923 B.n554 B.n553 585
R924 B.n552 B.n551 585
R925 B.n550 B.n549 585
R926 B.n548 B.n547 585
R927 B.n546 B.n545 585
R928 B.n544 B.n543 585
R929 B.n542 B.n541 585
R930 B.n540 B.n539 585
R931 B.n538 B.n537 585
R932 B.n536 B.n535 585
R933 B.n534 B.n533 585
R934 B.n532 B.n531 585
R935 B.n530 B.n529 585
R936 B.n528 B.n527 585
R937 B.n526 B.n525 585
R938 B.n524 B.n523 585
R939 B.n522 B.n521 585
R940 B.n520 B.n519 585
R941 B.n518 B.n517 585
R942 B.n516 B.n515 585
R943 B.n514 B.n513 585
R944 B.n512 B.n511 585
R945 B.n510 B.n509 585
R946 B.n508 B.n507 585
R947 B.n506 B.n505 585
R948 B.n504 B.n503 585
R949 B.n502 B.n501 585
R950 B.n500 B.n499 585
R951 B.n498 B.n497 585
R952 B.n496 B.n495 585
R953 B.n494 B.n493 585
R954 B.n492 B.n491 585
R955 B.n490 B.n489 585
R956 B.n487 B.n486 585
R957 B.n485 B.n484 585
R958 B.n483 B.n482 585
R959 B.n481 B.n480 585
R960 B.n479 B.n478 585
R961 B.n477 B.n476 585
R962 B.n475 B.n474 585
R963 B.n473 B.n472 585
R964 B.n471 B.n470 585
R965 B.n469 B.n468 585
R966 B.n466 B.n465 585
R967 B.n464 B.n463 585
R968 B.n462 B.n461 585
R969 B.n460 B.n459 585
R970 B.n458 B.n457 585
R971 B.n456 B.n455 585
R972 B.n454 B.n453 585
R973 B.n452 B.n451 585
R974 B.n450 B.n449 585
R975 B.n448 B.n447 585
R976 B.n446 B.n445 585
R977 B.n444 B.n443 585
R978 B.n442 B.n441 585
R979 B.n440 B.n439 585
R980 B.n438 B.n437 585
R981 B.n436 B.n435 585
R982 B.n434 B.n433 585
R983 B.n432 B.n431 585
R984 B.n430 B.n429 585
R985 B.n428 B.n427 585
R986 B.n426 B.n425 585
R987 B.n424 B.n423 585
R988 B.n422 B.n421 585
R989 B.n420 B.n419 585
R990 B.n418 B.n417 585
R991 B.n416 B.n415 585
R992 B.n414 B.n413 585
R993 B.n412 B.n411 585
R994 B.n410 B.n409 585
R995 B.n408 B.n407 585
R996 B.n406 B.n405 585
R997 B.n404 B.n403 585
R998 B.n402 B.n401 585
R999 B.n400 B.n399 585
R1000 B.n398 B.n397 585
R1001 B.n396 B.n395 585
R1002 B.n394 B.n393 585
R1003 B.n392 B.n391 585
R1004 B.n390 B.n389 585
R1005 B.n388 B.n387 585
R1006 B.n386 B.n385 585
R1007 B.n384 B.n383 585
R1008 B.n329 B.n328 585
R1009 B.n578 B.n577 585
R1010 B.n577 B.n576 585
R1011 B.n325 B.n324 585
R1012 B.n326 B.n325 585
R1013 B.n584 B.n583 585
R1014 B.n583 B.n582 585
R1015 B.n585 B.n323 585
R1016 B.n323 B.n321 585
R1017 B.n587 B.n586 585
R1018 B.n588 B.n587 585
R1019 B.n317 B.n316 585
R1020 B.n322 B.n317 585
R1021 B.n596 B.n595 585
R1022 B.n595 B.n594 585
R1023 B.n597 B.n315 585
R1024 B.n315 B.n314 585
R1025 B.n599 B.n598 585
R1026 B.n600 B.n599 585
R1027 B.n309 B.n308 585
R1028 B.n310 B.n309 585
R1029 B.n608 B.n607 585
R1030 B.n607 B.n606 585
R1031 B.n609 B.n307 585
R1032 B.n307 B.n306 585
R1033 B.n611 B.n610 585
R1034 B.n612 B.n611 585
R1035 B.n301 B.n300 585
R1036 B.n302 B.n301 585
R1037 B.n621 B.n620 585
R1038 B.n620 B.n619 585
R1039 B.n622 B.n299 585
R1040 B.n618 B.n299 585
R1041 B.n624 B.n623 585
R1042 B.n625 B.n624 585
R1043 B.n294 B.n293 585
R1044 B.n298 B.n294 585
R1045 B.n635 B.n634 585
R1046 B.n634 B.n633 585
R1047 B.n636 B.n292 585
R1048 B.n632 B.n292 585
R1049 B.n638 B.n637 585
R1050 B.n639 B.n638 585
R1051 B.n2 B.n0 585
R1052 B.n4 B.n2 585
R1053 B.n3 B.n1 585
R1054 B.n714 B.n3 585
R1055 B.n712 B.n711 585
R1056 B.n713 B.n712 585
R1057 B.n710 B.n8 585
R1058 B.n11 B.n8 585
R1059 B.n709 B.n708 585
R1060 B.n708 B.n707 585
R1061 B.n10 B.n9 585
R1062 B.n706 B.n10 585
R1063 B.n704 B.n703 585
R1064 B.n705 B.n704 585
R1065 B.n702 B.n15 585
R1066 B.n18 B.n15 585
R1067 B.n701 B.n700 585
R1068 B.n700 B.n699 585
R1069 B.n17 B.n16 585
R1070 B.n698 B.n17 585
R1071 B.n696 B.n695 585
R1072 B.n697 B.n696 585
R1073 B.n694 B.n23 585
R1074 B.n23 B.n22 585
R1075 B.n693 B.n692 585
R1076 B.n692 B.n691 585
R1077 B.n25 B.n24 585
R1078 B.n690 B.n25 585
R1079 B.n688 B.n687 585
R1080 B.n689 B.n688 585
R1081 B.n686 B.n30 585
R1082 B.n30 B.n29 585
R1083 B.n685 B.n684 585
R1084 B.n684 B.n683 585
R1085 B.n32 B.n31 585
R1086 B.n682 B.n32 585
R1087 B.n680 B.n679 585
R1088 B.n681 B.n680 585
R1089 B.n678 B.n37 585
R1090 B.n37 B.n36 585
R1091 B.n677 B.n676 585
R1092 B.n676 B.n675 585
R1093 B.n39 B.n38 585
R1094 B.n674 B.n39 585
R1095 B.n717 B.n716 585
R1096 B.n716 B.n715 585
R1097 B.n574 B.n325 473.281
R1098 B.n97 B.n39 473.281
R1099 B.n577 B.n327 473.281
R1100 B.n671 B.n41 473.281
R1101 B.n381 B.t13 311.757
R1102 B.n91 B.t19 311.757
R1103 B.n379 B.t16 311.757
R1104 B.n94 B.t22 311.757
R1105 B.n382 B.t12 297.793
R1106 B.n92 B.t20 297.793
R1107 B.n380 B.t15 297.793
R1108 B.n95 B.t23 297.793
R1109 B.n673 B.n672 256.663
R1110 B.n673 B.n89 256.663
R1111 B.n673 B.n88 256.663
R1112 B.n673 B.n87 256.663
R1113 B.n673 B.n86 256.663
R1114 B.n673 B.n85 256.663
R1115 B.n673 B.n84 256.663
R1116 B.n673 B.n83 256.663
R1117 B.n673 B.n82 256.663
R1118 B.n673 B.n81 256.663
R1119 B.n673 B.n80 256.663
R1120 B.n673 B.n79 256.663
R1121 B.n673 B.n78 256.663
R1122 B.n673 B.n77 256.663
R1123 B.n673 B.n76 256.663
R1124 B.n673 B.n75 256.663
R1125 B.n673 B.n74 256.663
R1126 B.n673 B.n73 256.663
R1127 B.n673 B.n72 256.663
R1128 B.n673 B.n71 256.663
R1129 B.n673 B.n70 256.663
R1130 B.n673 B.n69 256.663
R1131 B.n673 B.n68 256.663
R1132 B.n673 B.n67 256.663
R1133 B.n673 B.n66 256.663
R1134 B.n673 B.n65 256.663
R1135 B.n673 B.n64 256.663
R1136 B.n673 B.n63 256.663
R1137 B.n673 B.n62 256.663
R1138 B.n673 B.n61 256.663
R1139 B.n673 B.n60 256.663
R1140 B.n673 B.n59 256.663
R1141 B.n673 B.n58 256.663
R1142 B.n673 B.n57 256.663
R1143 B.n673 B.n56 256.663
R1144 B.n673 B.n55 256.663
R1145 B.n673 B.n54 256.663
R1146 B.n673 B.n53 256.663
R1147 B.n673 B.n52 256.663
R1148 B.n673 B.n51 256.663
R1149 B.n673 B.n50 256.663
R1150 B.n673 B.n49 256.663
R1151 B.n673 B.n48 256.663
R1152 B.n673 B.n47 256.663
R1153 B.n673 B.n46 256.663
R1154 B.n673 B.n45 256.663
R1155 B.n673 B.n44 256.663
R1156 B.n673 B.n43 256.663
R1157 B.n673 B.n42 256.663
R1158 B.n576 B.n575 256.663
R1159 B.n576 B.n330 256.663
R1160 B.n576 B.n331 256.663
R1161 B.n576 B.n332 256.663
R1162 B.n576 B.n333 256.663
R1163 B.n576 B.n334 256.663
R1164 B.n576 B.n335 256.663
R1165 B.n576 B.n336 256.663
R1166 B.n576 B.n337 256.663
R1167 B.n576 B.n338 256.663
R1168 B.n576 B.n339 256.663
R1169 B.n576 B.n340 256.663
R1170 B.n576 B.n341 256.663
R1171 B.n576 B.n342 256.663
R1172 B.n576 B.n343 256.663
R1173 B.n576 B.n344 256.663
R1174 B.n576 B.n345 256.663
R1175 B.n576 B.n346 256.663
R1176 B.n576 B.n347 256.663
R1177 B.n576 B.n348 256.663
R1178 B.n576 B.n349 256.663
R1179 B.n576 B.n350 256.663
R1180 B.n576 B.n351 256.663
R1181 B.n576 B.n352 256.663
R1182 B.n576 B.n353 256.663
R1183 B.n576 B.n354 256.663
R1184 B.n576 B.n355 256.663
R1185 B.n576 B.n356 256.663
R1186 B.n576 B.n357 256.663
R1187 B.n576 B.n358 256.663
R1188 B.n576 B.n359 256.663
R1189 B.n576 B.n360 256.663
R1190 B.n576 B.n361 256.663
R1191 B.n576 B.n362 256.663
R1192 B.n576 B.n363 256.663
R1193 B.n576 B.n364 256.663
R1194 B.n576 B.n365 256.663
R1195 B.n576 B.n366 256.663
R1196 B.n576 B.n367 256.663
R1197 B.n576 B.n368 256.663
R1198 B.n576 B.n369 256.663
R1199 B.n576 B.n370 256.663
R1200 B.n576 B.n371 256.663
R1201 B.n576 B.n372 256.663
R1202 B.n576 B.n373 256.663
R1203 B.n576 B.n374 256.663
R1204 B.n576 B.n375 256.663
R1205 B.n576 B.n376 256.663
R1206 B.n583 B.n325 163.367
R1207 B.n583 B.n323 163.367
R1208 B.n587 B.n323 163.367
R1209 B.n587 B.n317 163.367
R1210 B.n595 B.n317 163.367
R1211 B.n595 B.n315 163.367
R1212 B.n599 B.n315 163.367
R1213 B.n599 B.n309 163.367
R1214 B.n607 B.n309 163.367
R1215 B.n607 B.n307 163.367
R1216 B.n611 B.n307 163.367
R1217 B.n611 B.n301 163.367
R1218 B.n620 B.n301 163.367
R1219 B.n620 B.n299 163.367
R1220 B.n624 B.n299 163.367
R1221 B.n624 B.n294 163.367
R1222 B.n634 B.n294 163.367
R1223 B.n634 B.n292 163.367
R1224 B.n638 B.n292 163.367
R1225 B.n638 B.n2 163.367
R1226 B.n716 B.n2 163.367
R1227 B.n716 B.n3 163.367
R1228 B.n712 B.n3 163.367
R1229 B.n712 B.n8 163.367
R1230 B.n708 B.n8 163.367
R1231 B.n708 B.n10 163.367
R1232 B.n704 B.n10 163.367
R1233 B.n704 B.n15 163.367
R1234 B.n700 B.n15 163.367
R1235 B.n700 B.n17 163.367
R1236 B.n696 B.n17 163.367
R1237 B.n696 B.n23 163.367
R1238 B.n692 B.n23 163.367
R1239 B.n692 B.n25 163.367
R1240 B.n688 B.n25 163.367
R1241 B.n688 B.n30 163.367
R1242 B.n684 B.n30 163.367
R1243 B.n684 B.n32 163.367
R1244 B.n680 B.n32 163.367
R1245 B.n680 B.n37 163.367
R1246 B.n676 B.n37 163.367
R1247 B.n676 B.n39 163.367
R1248 B.n378 B.n377 163.367
R1249 B.n569 B.n377 163.367
R1250 B.n567 B.n566 163.367
R1251 B.n563 B.n562 163.367
R1252 B.n559 B.n558 163.367
R1253 B.n555 B.n554 163.367
R1254 B.n551 B.n550 163.367
R1255 B.n547 B.n546 163.367
R1256 B.n543 B.n542 163.367
R1257 B.n539 B.n538 163.367
R1258 B.n535 B.n534 163.367
R1259 B.n531 B.n530 163.367
R1260 B.n527 B.n526 163.367
R1261 B.n523 B.n522 163.367
R1262 B.n519 B.n518 163.367
R1263 B.n515 B.n514 163.367
R1264 B.n511 B.n510 163.367
R1265 B.n507 B.n506 163.367
R1266 B.n503 B.n502 163.367
R1267 B.n499 B.n498 163.367
R1268 B.n495 B.n494 163.367
R1269 B.n491 B.n490 163.367
R1270 B.n486 B.n485 163.367
R1271 B.n482 B.n481 163.367
R1272 B.n478 B.n477 163.367
R1273 B.n474 B.n473 163.367
R1274 B.n470 B.n469 163.367
R1275 B.n465 B.n464 163.367
R1276 B.n461 B.n460 163.367
R1277 B.n457 B.n456 163.367
R1278 B.n453 B.n452 163.367
R1279 B.n449 B.n448 163.367
R1280 B.n445 B.n444 163.367
R1281 B.n441 B.n440 163.367
R1282 B.n437 B.n436 163.367
R1283 B.n433 B.n432 163.367
R1284 B.n429 B.n428 163.367
R1285 B.n425 B.n424 163.367
R1286 B.n421 B.n420 163.367
R1287 B.n417 B.n416 163.367
R1288 B.n413 B.n412 163.367
R1289 B.n409 B.n408 163.367
R1290 B.n405 B.n404 163.367
R1291 B.n401 B.n400 163.367
R1292 B.n397 B.n396 163.367
R1293 B.n393 B.n392 163.367
R1294 B.n389 B.n388 163.367
R1295 B.n385 B.n384 163.367
R1296 B.n577 B.n329 163.367
R1297 B.n581 B.n327 163.367
R1298 B.n581 B.n320 163.367
R1299 B.n589 B.n320 163.367
R1300 B.n589 B.n318 163.367
R1301 B.n593 B.n318 163.367
R1302 B.n593 B.n313 163.367
R1303 B.n601 B.n313 163.367
R1304 B.n601 B.n311 163.367
R1305 B.n605 B.n311 163.367
R1306 B.n605 B.n305 163.367
R1307 B.n613 B.n305 163.367
R1308 B.n613 B.n303 163.367
R1309 B.n617 B.n303 163.367
R1310 B.n617 B.n297 163.367
R1311 B.n626 B.n297 163.367
R1312 B.n626 B.n295 163.367
R1313 B.n631 B.n295 163.367
R1314 B.n631 B.n291 163.367
R1315 B.n640 B.n291 163.367
R1316 B.n641 B.n640 163.367
R1317 B.n641 B.n5 163.367
R1318 B.n6 B.n5 163.367
R1319 B.n7 B.n6 163.367
R1320 B.n646 B.n7 163.367
R1321 B.n646 B.n12 163.367
R1322 B.n13 B.n12 163.367
R1323 B.n14 B.n13 163.367
R1324 B.n651 B.n14 163.367
R1325 B.n651 B.n19 163.367
R1326 B.n20 B.n19 163.367
R1327 B.n21 B.n20 163.367
R1328 B.n656 B.n21 163.367
R1329 B.n656 B.n26 163.367
R1330 B.n27 B.n26 163.367
R1331 B.n28 B.n27 163.367
R1332 B.n661 B.n28 163.367
R1333 B.n661 B.n33 163.367
R1334 B.n34 B.n33 163.367
R1335 B.n35 B.n34 163.367
R1336 B.n666 B.n35 163.367
R1337 B.n666 B.n40 163.367
R1338 B.n41 B.n40 163.367
R1339 B.n101 B.n100 163.367
R1340 B.n105 B.n104 163.367
R1341 B.n109 B.n108 163.367
R1342 B.n113 B.n112 163.367
R1343 B.n117 B.n116 163.367
R1344 B.n121 B.n120 163.367
R1345 B.n125 B.n124 163.367
R1346 B.n129 B.n128 163.367
R1347 B.n133 B.n132 163.367
R1348 B.n137 B.n136 163.367
R1349 B.n141 B.n140 163.367
R1350 B.n145 B.n144 163.367
R1351 B.n149 B.n148 163.367
R1352 B.n153 B.n152 163.367
R1353 B.n157 B.n156 163.367
R1354 B.n161 B.n160 163.367
R1355 B.n165 B.n164 163.367
R1356 B.n169 B.n168 163.367
R1357 B.n173 B.n172 163.367
R1358 B.n177 B.n176 163.367
R1359 B.n181 B.n180 163.367
R1360 B.n185 B.n184 163.367
R1361 B.n189 B.n188 163.367
R1362 B.n193 B.n192 163.367
R1363 B.n197 B.n196 163.367
R1364 B.n201 B.n200 163.367
R1365 B.n205 B.n204 163.367
R1366 B.n209 B.n208 163.367
R1367 B.n213 B.n212 163.367
R1368 B.n217 B.n216 163.367
R1369 B.n221 B.n220 163.367
R1370 B.n225 B.n224 163.367
R1371 B.n229 B.n228 163.367
R1372 B.n233 B.n232 163.367
R1373 B.n237 B.n236 163.367
R1374 B.n241 B.n240 163.367
R1375 B.n245 B.n244 163.367
R1376 B.n249 B.n248 163.367
R1377 B.n253 B.n252 163.367
R1378 B.n257 B.n256 163.367
R1379 B.n261 B.n260 163.367
R1380 B.n265 B.n264 163.367
R1381 B.n269 B.n268 163.367
R1382 B.n273 B.n272 163.367
R1383 B.n277 B.n276 163.367
R1384 B.n281 B.n280 163.367
R1385 B.n285 B.n284 163.367
R1386 B.n287 B.n90 163.367
R1387 B.n575 B.n574 71.676
R1388 B.n569 B.n330 71.676
R1389 B.n566 B.n331 71.676
R1390 B.n562 B.n332 71.676
R1391 B.n558 B.n333 71.676
R1392 B.n554 B.n334 71.676
R1393 B.n550 B.n335 71.676
R1394 B.n546 B.n336 71.676
R1395 B.n542 B.n337 71.676
R1396 B.n538 B.n338 71.676
R1397 B.n534 B.n339 71.676
R1398 B.n530 B.n340 71.676
R1399 B.n526 B.n341 71.676
R1400 B.n522 B.n342 71.676
R1401 B.n518 B.n343 71.676
R1402 B.n514 B.n344 71.676
R1403 B.n510 B.n345 71.676
R1404 B.n506 B.n346 71.676
R1405 B.n502 B.n347 71.676
R1406 B.n498 B.n348 71.676
R1407 B.n494 B.n349 71.676
R1408 B.n490 B.n350 71.676
R1409 B.n485 B.n351 71.676
R1410 B.n481 B.n352 71.676
R1411 B.n477 B.n353 71.676
R1412 B.n473 B.n354 71.676
R1413 B.n469 B.n355 71.676
R1414 B.n464 B.n356 71.676
R1415 B.n460 B.n357 71.676
R1416 B.n456 B.n358 71.676
R1417 B.n452 B.n359 71.676
R1418 B.n448 B.n360 71.676
R1419 B.n444 B.n361 71.676
R1420 B.n440 B.n362 71.676
R1421 B.n436 B.n363 71.676
R1422 B.n432 B.n364 71.676
R1423 B.n428 B.n365 71.676
R1424 B.n424 B.n366 71.676
R1425 B.n420 B.n367 71.676
R1426 B.n416 B.n368 71.676
R1427 B.n412 B.n369 71.676
R1428 B.n408 B.n370 71.676
R1429 B.n404 B.n371 71.676
R1430 B.n400 B.n372 71.676
R1431 B.n396 B.n373 71.676
R1432 B.n392 B.n374 71.676
R1433 B.n388 B.n375 71.676
R1434 B.n384 B.n376 71.676
R1435 B.n97 B.n42 71.676
R1436 B.n101 B.n43 71.676
R1437 B.n105 B.n44 71.676
R1438 B.n109 B.n45 71.676
R1439 B.n113 B.n46 71.676
R1440 B.n117 B.n47 71.676
R1441 B.n121 B.n48 71.676
R1442 B.n125 B.n49 71.676
R1443 B.n129 B.n50 71.676
R1444 B.n133 B.n51 71.676
R1445 B.n137 B.n52 71.676
R1446 B.n141 B.n53 71.676
R1447 B.n145 B.n54 71.676
R1448 B.n149 B.n55 71.676
R1449 B.n153 B.n56 71.676
R1450 B.n157 B.n57 71.676
R1451 B.n161 B.n58 71.676
R1452 B.n165 B.n59 71.676
R1453 B.n169 B.n60 71.676
R1454 B.n173 B.n61 71.676
R1455 B.n177 B.n62 71.676
R1456 B.n181 B.n63 71.676
R1457 B.n185 B.n64 71.676
R1458 B.n189 B.n65 71.676
R1459 B.n193 B.n66 71.676
R1460 B.n197 B.n67 71.676
R1461 B.n201 B.n68 71.676
R1462 B.n205 B.n69 71.676
R1463 B.n209 B.n70 71.676
R1464 B.n213 B.n71 71.676
R1465 B.n217 B.n72 71.676
R1466 B.n221 B.n73 71.676
R1467 B.n225 B.n74 71.676
R1468 B.n229 B.n75 71.676
R1469 B.n233 B.n76 71.676
R1470 B.n237 B.n77 71.676
R1471 B.n241 B.n78 71.676
R1472 B.n245 B.n79 71.676
R1473 B.n249 B.n80 71.676
R1474 B.n253 B.n81 71.676
R1475 B.n257 B.n82 71.676
R1476 B.n261 B.n83 71.676
R1477 B.n265 B.n84 71.676
R1478 B.n269 B.n85 71.676
R1479 B.n273 B.n86 71.676
R1480 B.n277 B.n87 71.676
R1481 B.n281 B.n88 71.676
R1482 B.n285 B.n89 71.676
R1483 B.n672 B.n90 71.676
R1484 B.n672 B.n671 71.676
R1485 B.n287 B.n89 71.676
R1486 B.n284 B.n88 71.676
R1487 B.n280 B.n87 71.676
R1488 B.n276 B.n86 71.676
R1489 B.n272 B.n85 71.676
R1490 B.n268 B.n84 71.676
R1491 B.n264 B.n83 71.676
R1492 B.n260 B.n82 71.676
R1493 B.n256 B.n81 71.676
R1494 B.n252 B.n80 71.676
R1495 B.n248 B.n79 71.676
R1496 B.n244 B.n78 71.676
R1497 B.n240 B.n77 71.676
R1498 B.n236 B.n76 71.676
R1499 B.n232 B.n75 71.676
R1500 B.n228 B.n74 71.676
R1501 B.n224 B.n73 71.676
R1502 B.n220 B.n72 71.676
R1503 B.n216 B.n71 71.676
R1504 B.n212 B.n70 71.676
R1505 B.n208 B.n69 71.676
R1506 B.n204 B.n68 71.676
R1507 B.n200 B.n67 71.676
R1508 B.n196 B.n66 71.676
R1509 B.n192 B.n65 71.676
R1510 B.n188 B.n64 71.676
R1511 B.n184 B.n63 71.676
R1512 B.n180 B.n62 71.676
R1513 B.n176 B.n61 71.676
R1514 B.n172 B.n60 71.676
R1515 B.n168 B.n59 71.676
R1516 B.n164 B.n58 71.676
R1517 B.n160 B.n57 71.676
R1518 B.n156 B.n56 71.676
R1519 B.n152 B.n55 71.676
R1520 B.n148 B.n54 71.676
R1521 B.n144 B.n53 71.676
R1522 B.n140 B.n52 71.676
R1523 B.n136 B.n51 71.676
R1524 B.n132 B.n50 71.676
R1525 B.n128 B.n49 71.676
R1526 B.n124 B.n48 71.676
R1527 B.n120 B.n47 71.676
R1528 B.n116 B.n46 71.676
R1529 B.n112 B.n45 71.676
R1530 B.n108 B.n44 71.676
R1531 B.n104 B.n43 71.676
R1532 B.n100 B.n42 71.676
R1533 B.n575 B.n378 71.676
R1534 B.n567 B.n330 71.676
R1535 B.n563 B.n331 71.676
R1536 B.n559 B.n332 71.676
R1537 B.n555 B.n333 71.676
R1538 B.n551 B.n334 71.676
R1539 B.n547 B.n335 71.676
R1540 B.n543 B.n336 71.676
R1541 B.n539 B.n337 71.676
R1542 B.n535 B.n338 71.676
R1543 B.n531 B.n339 71.676
R1544 B.n527 B.n340 71.676
R1545 B.n523 B.n341 71.676
R1546 B.n519 B.n342 71.676
R1547 B.n515 B.n343 71.676
R1548 B.n511 B.n344 71.676
R1549 B.n507 B.n345 71.676
R1550 B.n503 B.n346 71.676
R1551 B.n499 B.n347 71.676
R1552 B.n495 B.n348 71.676
R1553 B.n491 B.n349 71.676
R1554 B.n486 B.n350 71.676
R1555 B.n482 B.n351 71.676
R1556 B.n478 B.n352 71.676
R1557 B.n474 B.n353 71.676
R1558 B.n470 B.n354 71.676
R1559 B.n465 B.n355 71.676
R1560 B.n461 B.n356 71.676
R1561 B.n457 B.n357 71.676
R1562 B.n453 B.n358 71.676
R1563 B.n449 B.n359 71.676
R1564 B.n445 B.n360 71.676
R1565 B.n441 B.n361 71.676
R1566 B.n437 B.n362 71.676
R1567 B.n433 B.n363 71.676
R1568 B.n429 B.n364 71.676
R1569 B.n425 B.n365 71.676
R1570 B.n421 B.n366 71.676
R1571 B.n417 B.n367 71.676
R1572 B.n413 B.n368 71.676
R1573 B.n409 B.n369 71.676
R1574 B.n405 B.n370 71.676
R1575 B.n401 B.n371 71.676
R1576 B.n397 B.n372 71.676
R1577 B.n393 B.n373 71.676
R1578 B.n389 B.n374 71.676
R1579 B.n385 B.n375 71.676
R1580 B.n376 B.n329 71.676
R1581 B.n576 B.n326 67.2177
R1582 B.n674 B.n673 67.2177
R1583 B.n467 B.n382 59.5399
R1584 B.n488 B.n380 59.5399
R1585 B.n96 B.n95 59.5399
R1586 B.n93 B.n92 59.5399
R1587 B.n582 B.n326 41.1786
R1588 B.n582 B.n321 41.1786
R1589 B.n588 B.n321 41.1786
R1590 B.n588 B.n322 41.1786
R1591 B.n594 B.n314 41.1786
R1592 B.n600 B.n314 41.1786
R1593 B.n600 B.n310 41.1786
R1594 B.n606 B.n310 41.1786
R1595 B.n612 B.n306 41.1786
R1596 B.n619 B.n302 41.1786
R1597 B.n619 B.n618 41.1786
R1598 B.n625 B.n298 41.1786
R1599 B.n633 B.n632 41.1786
R1600 B.n639 B.n4 41.1786
R1601 B.n715 B.n4 41.1786
R1602 B.n715 B.n714 41.1786
R1603 B.n714 B.n713 41.1786
R1604 B.n707 B.n11 41.1786
R1605 B.n706 B.n705 41.1786
R1606 B.n699 B.n18 41.1786
R1607 B.n699 B.n698 41.1786
R1608 B.n697 B.n22 41.1786
R1609 B.n691 B.n690 41.1786
R1610 B.n690 B.n689 41.1786
R1611 B.n689 B.n29 41.1786
R1612 B.n683 B.n29 41.1786
R1613 B.n682 B.n681 41.1786
R1614 B.n681 B.n36 41.1786
R1615 B.n675 B.n36 41.1786
R1616 B.n675 B.n674 41.1786
R1617 B.n612 B.t3 40.573
R1618 B.t6 B.n697 40.573
R1619 B.n625 B.t8 36.9397
R1620 B.n705 B.t1 36.9397
R1621 B.n606 B.t7 35.7285
R1622 B.n691 B.t0 35.7285
R1623 B.n633 B.t2 32.0952
R1624 B.n707 B.t9 32.0952
R1625 B.n98 B.n38 30.7517
R1626 B.n579 B.n578 30.7517
R1627 B.n573 B.n324 30.7517
R1628 B.n670 B.n669 30.7517
R1629 B.n639 B.t5 27.2507
R1630 B.n713 B.t4 27.2507
R1631 B.n322 B.t11 22.4062
R1632 B.t18 B.n682 22.4062
R1633 B.n594 B.t11 18.7729
R1634 B.n683 B.t18 18.7729
R1635 B B.n717 18.0485
R1636 B.n382 B.n381 13.9641
R1637 B.n380 B.n379 13.9641
R1638 B.n95 B.n94 13.9641
R1639 B.n92 B.n91 13.9641
R1640 B.n632 B.t5 13.9284
R1641 B.n11 B.t4 13.9284
R1642 B.n99 B.n98 10.6151
R1643 B.n102 B.n99 10.6151
R1644 B.n103 B.n102 10.6151
R1645 B.n106 B.n103 10.6151
R1646 B.n107 B.n106 10.6151
R1647 B.n110 B.n107 10.6151
R1648 B.n111 B.n110 10.6151
R1649 B.n114 B.n111 10.6151
R1650 B.n115 B.n114 10.6151
R1651 B.n118 B.n115 10.6151
R1652 B.n119 B.n118 10.6151
R1653 B.n122 B.n119 10.6151
R1654 B.n123 B.n122 10.6151
R1655 B.n126 B.n123 10.6151
R1656 B.n127 B.n126 10.6151
R1657 B.n130 B.n127 10.6151
R1658 B.n131 B.n130 10.6151
R1659 B.n134 B.n131 10.6151
R1660 B.n135 B.n134 10.6151
R1661 B.n138 B.n135 10.6151
R1662 B.n139 B.n138 10.6151
R1663 B.n142 B.n139 10.6151
R1664 B.n143 B.n142 10.6151
R1665 B.n146 B.n143 10.6151
R1666 B.n147 B.n146 10.6151
R1667 B.n150 B.n147 10.6151
R1668 B.n151 B.n150 10.6151
R1669 B.n154 B.n151 10.6151
R1670 B.n155 B.n154 10.6151
R1671 B.n158 B.n155 10.6151
R1672 B.n159 B.n158 10.6151
R1673 B.n162 B.n159 10.6151
R1674 B.n163 B.n162 10.6151
R1675 B.n166 B.n163 10.6151
R1676 B.n167 B.n166 10.6151
R1677 B.n170 B.n167 10.6151
R1678 B.n171 B.n170 10.6151
R1679 B.n174 B.n171 10.6151
R1680 B.n175 B.n174 10.6151
R1681 B.n178 B.n175 10.6151
R1682 B.n179 B.n178 10.6151
R1683 B.n182 B.n179 10.6151
R1684 B.n183 B.n182 10.6151
R1685 B.n187 B.n186 10.6151
R1686 B.n190 B.n187 10.6151
R1687 B.n191 B.n190 10.6151
R1688 B.n194 B.n191 10.6151
R1689 B.n195 B.n194 10.6151
R1690 B.n198 B.n195 10.6151
R1691 B.n199 B.n198 10.6151
R1692 B.n202 B.n199 10.6151
R1693 B.n203 B.n202 10.6151
R1694 B.n207 B.n206 10.6151
R1695 B.n210 B.n207 10.6151
R1696 B.n211 B.n210 10.6151
R1697 B.n214 B.n211 10.6151
R1698 B.n215 B.n214 10.6151
R1699 B.n218 B.n215 10.6151
R1700 B.n219 B.n218 10.6151
R1701 B.n222 B.n219 10.6151
R1702 B.n223 B.n222 10.6151
R1703 B.n226 B.n223 10.6151
R1704 B.n227 B.n226 10.6151
R1705 B.n230 B.n227 10.6151
R1706 B.n231 B.n230 10.6151
R1707 B.n234 B.n231 10.6151
R1708 B.n235 B.n234 10.6151
R1709 B.n238 B.n235 10.6151
R1710 B.n239 B.n238 10.6151
R1711 B.n242 B.n239 10.6151
R1712 B.n243 B.n242 10.6151
R1713 B.n246 B.n243 10.6151
R1714 B.n247 B.n246 10.6151
R1715 B.n250 B.n247 10.6151
R1716 B.n251 B.n250 10.6151
R1717 B.n254 B.n251 10.6151
R1718 B.n255 B.n254 10.6151
R1719 B.n258 B.n255 10.6151
R1720 B.n259 B.n258 10.6151
R1721 B.n262 B.n259 10.6151
R1722 B.n263 B.n262 10.6151
R1723 B.n266 B.n263 10.6151
R1724 B.n267 B.n266 10.6151
R1725 B.n270 B.n267 10.6151
R1726 B.n271 B.n270 10.6151
R1727 B.n274 B.n271 10.6151
R1728 B.n275 B.n274 10.6151
R1729 B.n278 B.n275 10.6151
R1730 B.n279 B.n278 10.6151
R1731 B.n282 B.n279 10.6151
R1732 B.n283 B.n282 10.6151
R1733 B.n286 B.n283 10.6151
R1734 B.n288 B.n286 10.6151
R1735 B.n289 B.n288 10.6151
R1736 B.n670 B.n289 10.6151
R1737 B.n580 B.n579 10.6151
R1738 B.n580 B.n319 10.6151
R1739 B.n590 B.n319 10.6151
R1740 B.n591 B.n590 10.6151
R1741 B.n592 B.n591 10.6151
R1742 B.n592 B.n312 10.6151
R1743 B.n602 B.n312 10.6151
R1744 B.n603 B.n602 10.6151
R1745 B.n604 B.n603 10.6151
R1746 B.n604 B.n304 10.6151
R1747 B.n614 B.n304 10.6151
R1748 B.n615 B.n614 10.6151
R1749 B.n616 B.n615 10.6151
R1750 B.n616 B.n296 10.6151
R1751 B.n627 B.n296 10.6151
R1752 B.n628 B.n627 10.6151
R1753 B.n630 B.n628 10.6151
R1754 B.n630 B.n629 10.6151
R1755 B.n629 B.n290 10.6151
R1756 B.n642 B.n290 10.6151
R1757 B.n643 B.n642 10.6151
R1758 B.n644 B.n643 10.6151
R1759 B.n645 B.n644 10.6151
R1760 B.n647 B.n645 10.6151
R1761 B.n648 B.n647 10.6151
R1762 B.n649 B.n648 10.6151
R1763 B.n650 B.n649 10.6151
R1764 B.n652 B.n650 10.6151
R1765 B.n653 B.n652 10.6151
R1766 B.n654 B.n653 10.6151
R1767 B.n655 B.n654 10.6151
R1768 B.n657 B.n655 10.6151
R1769 B.n658 B.n657 10.6151
R1770 B.n659 B.n658 10.6151
R1771 B.n660 B.n659 10.6151
R1772 B.n662 B.n660 10.6151
R1773 B.n663 B.n662 10.6151
R1774 B.n664 B.n663 10.6151
R1775 B.n665 B.n664 10.6151
R1776 B.n667 B.n665 10.6151
R1777 B.n668 B.n667 10.6151
R1778 B.n669 B.n668 10.6151
R1779 B.n573 B.n572 10.6151
R1780 B.n572 B.n571 10.6151
R1781 B.n571 B.n570 10.6151
R1782 B.n570 B.n568 10.6151
R1783 B.n568 B.n565 10.6151
R1784 B.n565 B.n564 10.6151
R1785 B.n564 B.n561 10.6151
R1786 B.n561 B.n560 10.6151
R1787 B.n560 B.n557 10.6151
R1788 B.n557 B.n556 10.6151
R1789 B.n556 B.n553 10.6151
R1790 B.n553 B.n552 10.6151
R1791 B.n552 B.n549 10.6151
R1792 B.n549 B.n548 10.6151
R1793 B.n548 B.n545 10.6151
R1794 B.n545 B.n544 10.6151
R1795 B.n544 B.n541 10.6151
R1796 B.n541 B.n540 10.6151
R1797 B.n540 B.n537 10.6151
R1798 B.n537 B.n536 10.6151
R1799 B.n536 B.n533 10.6151
R1800 B.n533 B.n532 10.6151
R1801 B.n532 B.n529 10.6151
R1802 B.n529 B.n528 10.6151
R1803 B.n528 B.n525 10.6151
R1804 B.n525 B.n524 10.6151
R1805 B.n524 B.n521 10.6151
R1806 B.n521 B.n520 10.6151
R1807 B.n520 B.n517 10.6151
R1808 B.n517 B.n516 10.6151
R1809 B.n516 B.n513 10.6151
R1810 B.n513 B.n512 10.6151
R1811 B.n512 B.n509 10.6151
R1812 B.n509 B.n508 10.6151
R1813 B.n508 B.n505 10.6151
R1814 B.n505 B.n504 10.6151
R1815 B.n504 B.n501 10.6151
R1816 B.n501 B.n500 10.6151
R1817 B.n500 B.n497 10.6151
R1818 B.n497 B.n496 10.6151
R1819 B.n496 B.n493 10.6151
R1820 B.n493 B.n492 10.6151
R1821 B.n492 B.n489 10.6151
R1822 B.n487 B.n484 10.6151
R1823 B.n484 B.n483 10.6151
R1824 B.n483 B.n480 10.6151
R1825 B.n480 B.n479 10.6151
R1826 B.n479 B.n476 10.6151
R1827 B.n476 B.n475 10.6151
R1828 B.n475 B.n472 10.6151
R1829 B.n472 B.n471 10.6151
R1830 B.n471 B.n468 10.6151
R1831 B.n466 B.n463 10.6151
R1832 B.n463 B.n462 10.6151
R1833 B.n462 B.n459 10.6151
R1834 B.n459 B.n458 10.6151
R1835 B.n458 B.n455 10.6151
R1836 B.n455 B.n454 10.6151
R1837 B.n454 B.n451 10.6151
R1838 B.n451 B.n450 10.6151
R1839 B.n450 B.n447 10.6151
R1840 B.n447 B.n446 10.6151
R1841 B.n446 B.n443 10.6151
R1842 B.n443 B.n442 10.6151
R1843 B.n442 B.n439 10.6151
R1844 B.n439 B.n438 10.6151
R1845 B.n438 B.n435 10.6151
R1846 B.n435 B.n434 10.6151
R1847 B.n434 B.n431 10.6151
R1848 B.n431 B.n430 10.6151
R1849 B.n430 B.n427 10.6151
R1850 B.n427 B.n426 10.6151
R1851 B.n426 B.n423 10.6151
R1852 B.n423 B.n422 10.6151
R1853 B.n422 B.n419 10.6151
R1854 B.n419 B.n418 10.6151
R1855 B.n418 B.n415 10.6151
R1856 B.n415 B.n414 10.6151
R1857 B.n414 B.n411 10.6151
R1858 B.n411 B.n410 10.6151
R1859 B.n410 B.n407 10.6151
R1860 B.n407 B.n406 10.6151
R1861 B.n406 B.n403 10.6151
R1862 B.n403 B.n402 10.6151
R1863 B.n402 B.n399 10.6151
R1864 B.n399 B.n398 10.6151
R1865 B.n398 B.n395 10.6151
R1866 B.n395 B.n394 10.6151
R1867 B.n394 B.n391 10.6151
R1868 B.n391 B.n390 10.6151
R1869 B.n390 B.n387 10.6151
R1870 B.n387 B.n386 10.6151
R1871 B.n386 B.n383 10.6151
R1872 B.n383 B.n328 10.6151
R1873 B.n578 B.n328 10.6151
R1874 B.n584 B.n324 10.6151
R1875 B.n585 B.n584 10.6151
R1876 B.n586 B.n585 10.6151
R1877 B.n586 B.n316 10.6151
R1878 B.n596 B.n316 10.6151
R1879 B.n597 B.n596 10.6151
R1880 B.n598 B.n597 10.6151
R1881 B.n598 B.n308 10.6151
R1882 B.n608 B.n308 10.6151
R1883 B.n609 B.n608 10.6151
R1884 B.n610 B.n609 10.6151
R1885 B.n610 B.n300 10.6151
R1886 B.n621 B.n300 10.6151
R1887 B.n622 B.n621 10.6151
R1888 B.n623 B.n622 10.6151
R1889 B.n623 B.n293 10.6151
R1890 B.n635 B.n293 10.6151
R1891 B.n636 B.n635 10.6151
R1892 B.n637 B.n636 10.6151
R1893 B.n637 B.n0 10.6151
R1894 B.n711 B.n1 10.6151
R1895 B.n711 B.n710 10.6151
R1896 B.n710 B.n709 10.6151
R1897 B.n709 B.n9 10.6151
R1898 B.n703 B.n9 10.6151
R1899 B.n703 B.n702 10.6151
R1900 B.n702 B.n701 10.6151
R1901 B.n701 B.n16 10.6151
R1902 B.n695 B.n16 10.6151
R1903 B.n695 B.n694 10.6151
R1904 B.n694 B.n693 10.6151
R1905 B.n693 B.n24 10.6151
R1906 B.n687 B.n24 10.6151
R1907 B.n687 B.n686 10.6151
R1908 B.n686 B.n685 10.6151
R1909 B.n685 B.n31 10.6151
R1910 B.n679 B.n31 10.6151
R1911 B.n679 B.n678 10.6151
R1912 B.n678 B.n677 10.6151
R1913 B.n677 B.n38 10.6151
R1914 B.n183 B.n96 9.36635
R1915 B.n206 B.n93 9.36635
R1916 B.n489 B.n488 9.36635
R1917 B.n467 B.n466 9.36635
R1918 B.n298 B.t2 9.0839
R1919 B.t9 B.n706 9.0839
R1920 B.t7 B.n306 5.45054
R1921 B.t0 B.n22 5.45054
R1922 B.n618 B.t8 4.23942
R1923 B.n18 B.t1 4.23942
R1924 B.n717 B.n0 2.81026
R1925 B.n717 B.n1 2.81026
R1926 B.n186 B.n96 1.24928
R1927 B.n203 B.n93 1.24928
R1928 B.n488 B.n487 1.24928
R1929 B.n468 B.n467 1.24928
R1930 B.t3 B.n302 0.60606
R1931 B.n698 B.t6 0.60606
R1932 VP.n5 VP.t3 918.861
R1933 VP.n15 VP.t5 897.88
R1934 VP.n16 VP.t4 897.88
R1935 VP.n1 VP.t8 897.88
R1936 VP.n21 VP.t9 897.88
R1937 VP.n22 VP.t1 897.88
R1938 VP.n12 VP.t0 897.88
R1939 VP.n11 VP.t6 897.88
R1940 VP.n4 VP.t2 897.88
R1941 VP.n6 VP.t7 897.88
R1942 VP.n23 VP.n22 161.3
R1943 VP.n8 VP.n7 161.3
R1944 VP.n10 VP.n9 161.3
R1945 VP.n11 VP.n3 161.3
R1946 VP.n13 VP.n12 161.3
R1947 VP.n21 VP.n0 161.3
R1948 VP.n20 VP.n19 161.3
R1949 VP.n18 VP.n17 161.3
R1950 VP.n16 VP.n2 161.3
R1951 VP.n15 VP.n14 161.3
R1952 VP.n8 VP.n5 70.4033
R1953 VP.n16 VP.n15 48.2005
R1954 VP.n22 VP.n21 48.2005
R1955 VP.n12 VP.n11 48.2005
R1956 VP.n14 VP.n13 41.796
R1957 VP.n17 VP.n16 40.1672
R1958 VP.n21 VP.n20 40.1672
R1959 VP.n11 VP.n10 40.1672
R1960 VP.n7 VP.n6 40.1672
R1961 VP.n6 VP.n5 20.9576
R1962 VP.n17 VP.n1 8.03383
R1963 VP.n20 VP.n1 8.03383
R1964 VP.n10 VP.n4 8.03383
R1965 VP.n7 VP.n4 8.03383
R1966 VP.n9 VP.n8 0.189894
R1967 VP.n9 VP.n3 0.189894
R1968 VP.n13 VP.n3 0.189894
R1969 VP.n14 VP.n2 0.189894
R1970 VP.n18 VP.n2 0.189894
R1971 VP.n19 VP.n18 0.189894
R1972 VP.n19 VP.n0 0.189894
R1973 VP.n23 VP.n0 0.189894
R1974 VP VP.n23 0.0516364
R1975 VDD1.n64 VDD1.n0 289.615
R1976 VDD1.n135 VDD1.n71 289.615
R1977 VDD1.n65 VDD1.n64 185
R1978 VDD1.n63 VDD1.n62 185
R1979 VDD1.n4 VDD1.n3 185
R1980 VDD1.n57 VDD1.n56 185
R1981 VDD1.n55 VDD1.n54 185
R1982 VDD1.n8 VDD1.n7 185
R1983 VDD1.n49 VDD1.n48 185
R1984 VDD1.n47 VDD1.n46 185
R1985 VDD1.n45 VDD1.n11 185
R1986 VDD1.n15 VDD1.n12 185
R1987 VDD1.n40 VDD1.n39 185
R1988 VDD1.n38 VDD1.n37 185
R1989 VDD1.n17 VDD1.n16 185
R1990 VDD1.n32 VDD1.n31 185
R1991 VDD1.n30 VDD1.n29 185
R1992 VDD1.n21 VDD1.n20 185
R1993 VDD1.n24 VDD1.n23 185
R1994 VDD1.n94 VDD1.n93 185
R1995 VDD1.n91 VDD1.n90 185
R1996 VDD1.n100 VDD1.n99 185
R1997 VDD1.n102 VDD1.n101 185
R1998 VDD1.n87 VDD1.n86 185
R1999 VDD1.n108 VDD1.n107 185
R2000 VDD1.n111 VDD1.n110 185
R2001 VDD1.n109 VDD1.n83 185
R2002 VDD1.n116 VDD1.n82 185
R2003 VDD1.n118 VDD1.n117 185
R2004 VDD1.n120 VDD1.n119 185
R2005 VDD1.n79 VDD1.n78 185
R2006 VDD1.n126 VDD1.n125 185
R2007 VDD1.n128 VDD1.n127 185
R2008 VDD1.n75 VDD1.n74 185
R2009 VDD1.n134 VDD1.n133 185
R2010 VDD1.n136 VDD1.n135 185
R2011 VDD1.t6 VDD1.n22 149.524
R2012 VDD1.t4 VDD1.n92 149.524
R2013 VDD1.n64 VDD1.n63 104.615
R2014 VDD1.n63 VDD1.n3 104.615
R2015 VDD1.n56 VDD1.n3 104.615
R2016 VDD1.n56 VDD1.n55 104.615
R2017 VDD1.n55 VDD1.n7 104.615
R2018 VDD1.n48 VDD1.n7 104.615
R2019 VDD1.n48 VDD1.n47 104.615
R2020 VDD1.n47 VDD1.n11 104.615
R2021 VDD1.n15 VDD1.n11 104.615
R2022 VDD1.n39 VDD1.n15 104.615
R2023 VDD1.n39 VDD1.n38 104.615
R2024 VDD1.n38 VDD1.n16 104.615
R2025 VDD1.n31 VDD1.n16 104.615
R2026 VDD1.n31 VDD1.n30 104.615
R2027 VDD1.n30 VDD1.n20 104.615
R2028 VDD1.n23 VDD1.n20 104.615
R2029 VDD1.n93 VDD1.n90 104.615
R2030 VDD1.n100 VDD1.n90 104.615
R2031 VDD1.n101 VDD1.n100 104.615
R2032 VDD1.n101 VDD1.n86 104.615
R2033 VDD1.n108 VDD1.n86 104.615
R2034 VDD1.n110 VDD1.n108 104.615
R2035 VDD1.n110 VDD1.n109 104.615
R2036 VDD1.n109 VDD1.n82 104.615
R2037 VDD1.n118 VDD1.n82 104.615
R2038 VDD1.n119 VDD1.n118 104.615
R2039 VDD1.n119 VDD1.n78 104.615
R2040 VDD1.n126 VDD1.n78 104.615
R2041 VDD1.n127 VDD1.n126 104.615
R2042 VDD1.n127 VDD1.n74 104.615
R2043 VDD1.n134 VDD1.n74 104.615
R2044 VDD1.n135 VDD1.n134 104.615
R2045 VDD1.n143 VDD1.n142 63.0831
R2046 VDD1.n70 VDD1.n69 62.673
R2047 VDD1.n141 VDD1.n140 62.673
R2048 VDD1.n145 VDD1.n144 62.6728
R2049 VDD1.n23 VDD1.t6 52.3082
R2050 VDD1.n93 VDD1.t4 52.3082
R2051 VDD1.n70 VDD1.n68 50.4545
R2052 VDD1.n141 VDD1.n139 50.4545
R2053 VDD1.n145 VDD1.n143 38.669
R2054 VDD1.n46 VDD1.n45 13.1884
R2055 VDD1.n117 VDD1.n116 13.1884
R2056 VDD1.n49 VDD1.n10 12.8005
R2057 VDD1.n44 VDD1.n12 12.8005
R2058 VDD1.n115 VDD1.n83 12.8005
R2059 VDD1.n120 VDD1.n81 12.8005
R2060 VDD1.n50 VDD1.n8 12.0247
R2061 VDD1.n41 VDD1.n40 12.0247
R2062 VDD1.n112 VDD1.n111 12.0247
R2063 VDD1.n121 VDD1.n79 12.0247
R2064 VDD1.n54 VDD1.n53 11.249
R2065 VDD1.n37 VDD1.n14 11.249
R2066 VDD1.n107 VDD1.n85 11.249
R2067 VDD1.n125 VDD1.n124 11.249
R2068 VDD1.n57 VDD1.n6 10.4732
R2069 VDD1.n36 VDD1.n17 10.4732
R2070 VDD1.n106 VDD1.n87 10.4732
R2071 VDD1.n128 VDD1.n77 10.4732
R2072 VDD1.n24 VDD1.n22 10.2747
R2073 VDD1.n94 VDD1.n92 10.2747
R2074 VDD1.n58 VDD1.n4 9.69747
R2075 VDD1.n33 VDD1.n32 9.69747
R2076 VDD1.n103 VDD1.n102 9.69747
R2077 VDD1.n129 VDD1.n75 9.69747
R2078 VDD1.n68 VDD1.n67 9.45567
R2079 VDD1.n139 VDD1.n138 9.45567
R2080 VDD1.n26 VDD1.n25 9.3005
R2081 VDD1.n28 VDD1.n27 9.3005
R2082 VDD1.n19 VDD1.n18 9.3005
R2083 VDD1.n34 VDD1.n33 9.3005
R2084 VDD1.n36 VDD1.n35 9.3005
R2085 VDD1.n14 VDD1.n13 9.3005
R2086 VDD1.n42 VDD1.n41 9.3005
R2087 VDD1.n44 VDD1.n43 9.3005
R2088 VDD1.n67 VDD1.n66 9.3005
R2089 VDD1.n2 VDD1.n1 9.3005
R2090 VDD1.n61 VDD1.n60 9.3005
R2091 VDD1.n59 VDD1.n58 9.3005
R2092 VDD1.n6 VDD1.n5 9.3005
R2093 VDD1.n53 VDD1.n52 9.3005
R2094 VDD1.n51 VDD1.n50 9.3005
R2095 VDD1.n10 VDD1.n9 9.3005
R2096 VDD1.n73 VDD1.n72 9.3005
R2097 VDD1.n132 VDD1.n131 9.3005
R2098 VDD1.n130 VDD1.n129 9.3005
R2099 VDD1.n77 VDD1.n76 9.3005
R2100 VDD1.n124 VDD1.n123 9.3005
R2101 VDD1.n122 VDD1.n121 9.3005
R2102 VDD1.n81 VDD1.n80 9.3005
R2103 VDD1.n96 VDD1.n95 9.3005
R2104 VDD1.n98 VDD1.n97 9.3005
R2105 VDD1.n89 VDD1.n88 9.3005
R2106 VDD1.n104 VDD1.n103 9.3005
R2107 VDD1.n106 VDD1.n105 9.3005
R2108 VDD1.n85 VDD1.n84 9.3005
R2109 VDD1.n113 VDD1.n112 9.3005
R2110 VDD1.n115 VDD1.n114 9.3005
R2111 VDD1.n138 VDD1.n137 9.3005
R2112 VDD1.n62 VDD1.n61 8.92171
R2113 VDD1.n29 VDD1.n19 8.92171
R2114 VDD1.n99 VDD1.n89 8.92171
R2115 VDD1.n133 VDD1.n132 8.92171
R2116 VDD1.n65 VDD1.n2 8.14595
R2117 VDD1.n28 VDD1.n21 8.14595
R2118 VDD1.n98 VDD1.n91 8.14595
R2119 VDD1.n136 VDD1.n73 8.14595
R2120 VDD1.n66 VDD1.n0 7.3702
R2121 VDD1.n25 VDD1.n24 7.3702
R2122 VDD1.n95 VDD1.n94 7.3702
R2123 VDD1.n137 VDD1.n71 7.3702
R2124 VDD1.n68 VDD1.n0 6.59444
R2125 VDD1.n139 VDD1.n71 6.59444
R2126 VDD1.n66 VDD1.n65 5.81868
R2127 VDD1.n25 VDD1.n21 5.81868
R2128 VDD1.n95 VDD1.n91 5.81868
R2129 VDD1.n137 VDD1.n136 5.81868
R2130 VDD1.n62 VDD1.n2 5.04292
R2131 VDD1.n29 VDD1.n28 5.04292
R2132 VDD1.n99 VDD1.n98 5.04292
R2133 VDD1.n133 VDD1.n73 5.04292
R2134 VDD1.n61 VDD1.n4 4.26717
R2135 VDD1.n32 VDD1.n19 4.26717
R2136 VDD1.n102 VDD1.n89 4.26717
R2137 VDD1.n132 VDD1.n75 4.26717
R2138 VDD1.n58 VDD1.n57 3.49141
R2139 VDD1.n33 VDD1.n17 3.49141
R2140 VDD1.n103 VDD1.n87 3.49141
R2141 VDD1.n129 VDD1.n128 3.49141
R2142 VDD1.n26 VDD1.n22 2.84303
R2143 VDD1.n96 VDD1.n92 2.84303
R2144 VDD1.n54 VDD1.n6 2.71565
R2145 VDD1.n37 VDD1.n36 2.71565
R2146 VDD1.n107 VDD1.n106 2.71565
R2147 VDD1.n125 VDD1.n77 2.71565
R2148 VDD1.n53 VDD1.n8 1.93989
R2149 VDD1.n40 VDD1.n14 1.93989
R2150 VDD1.n111 VDD1.n85 1.93989
R2151 VDD1.n124 VDD1.n79 1.93989
R2152 VDD1.n144 VDD1.t3 1.53657
R2153 VDD1.n144 VDD1.t9 1.53657
R2154 VDD1.n69 VDD1.t2 1.53657
R2155 VDD1.n69 VDD1.t7 1.53657
R2156 VDD1.n142 VDD1.t0 1.53657
R2157 VDD1.n142 VDD1.t8 1.53657
R2158 VDD1.n140 VDD1.t5 1.53657
R2159 VDD1.n140 VDD1.t1 1.53657
R2160 VDD1.n50 VDD1.n49 1.16414
R2161 VDD1.n41 VDD1.n12 1.16414
R2162 VDD1.n112 VDD1.n83 1.16414
R2163 VDD1.n121 VDD1.n120 1.16414
R2164 VDD1 VDD1.n145 0.407828
R2165 VDD1.n46 VDD1.n10 0.388379
R2166 VDD1.n45 VDD1.n44 0.388379
R2167 VDD1.n116 VDD1.n115 0.388379
R2168 VDD1.n117 VDD1.n81 0.388379
R2169 VDD1 VDD1.n70 0.213862
R2170 VDD1.n67 VDD1.n1 0.155672
R2171 VDD1.n60 VDD1.n1 0.155672
R2172 VDD1.n60 VDD1.n59 0.155672
R2173 VDD1.n59 VDD1.n5 0.155672
R2174 VDD1.n52 VDD1.n5 0.155672
R2175 VDD1.n52 VDD1.n51 0.155672
R2176 VDD1.n51 VDD1.n9 0.155672
R2177 VDD1.n43 VDD1.n9 0.155672
R2178 VDD1.n43 VDD1.n42 0.155672
R2179 VDD1.n42 VDD1.n13 0.155672
R2180 VDD1.n35 VDD1.n13 0.155672
R2181 VDD1.n35 VDD1.n34 0.155672
R2182 VDD1.n34 VDD1.n18 0.155672
R2183 VDD1.n27 VDD1.n18 0.155672
R2184 VDD1.n27 VDD1.n26 0.155672
R2185 VDD1.n97 VDD1.n96 0.155672
R2186 VDD1.n97 VDD1.n88 0.155672
R2187 VDD1.n104 VDD1.n88 0.155672
R2188 VDD1.n105 VDD1.n104 0.155672
R2189 VDD1.n105 VDD1.n84 0.155672
R2190 VDD1.n113 VDD1.n84 0.155672
R2191 VDD1.n114 VDD1.n113 0.155672
R2192 VDD1.n114 VDD1.n80 0.155672
R2193 VDD1.n122 VDD1.n80 0.155672
R2194 VDD1.n123 VDD1.n122 0.155672
R2195 VDD1.n123 VDD1.n76 0.155672
R2196 VDD1.n130 VDD1.n76 0.155672
R2197 VDD1.n131 VDD1.n130 0.155672
R2198 VDD1.n131 VDD1.n72 0.155672
R2199 VDD1.n138 VDD1.n72 0.155672
R2200 VDD1.n143 VDD1.n141 0.100326
C0 VN VP 5.30648f
C1 VP VDD2 0.302372f
C2 VDD1 VTAIL 19.773802f
C3 VP VTAIL 4.68502f
C4 VN VDD2 5.04536f
C5 VN VTAIL 4.67026f
C6 VDD2 VTAIL 19.8039f
C7 VDD1 VP 5.19397f
C8 VDD1 VN 0.148326f
C9 VDD1 VDD2 0.781156f
C10 VDD2 B 4.792572f
C11 VDD1 B 4.672749f
C12 VTAIL B 6.483735f
C13 VN B 8.270651f
C14 VP B 6.066381f
C15 VDD1.n0 B 0.040866f
C16 VDD1.n1 B 0.02787f
C17 VDD1.n2 B 0.014976f
C18 VDD1.n3 B 0.035398f
C19 VDD1.n4 B 0.015857f
C20 VDD1.n5 B 0.02787f
C21 VDD1.n6 B 0.014976f
C22 VDD1.n7 B 0.035398f
C23 VDD1.n8 B 0.015857f
C24 VDD1.n9 B 0.02787f
C25 VDD1.n10 B 0.014976f
C26 VDD1.n11 B 0.035398f
C27 VDD1.n12 B 0.015857f
C28 VDD1.n13 B 0.02787f
C29 VDD1.n14 B 0.014976f
C30 VDD1.n15 B 0.035398f
C31 VDD1.n16 B 0.035398f
C32 VDD1.n17 B 0.015857f
C33 VDD1.n18 B 0.02787f
C34 VDD1.n19 B 0.014976f
C35 VDD1.n20 B 0.035398f
C36 VDD1.n21 B 0.015857f
C37 VDD1.n22 B 0.21046f
C38 VDD1.t6 B 0.059918f
C39 VDD1.n23 B 0.026548f
C40 VDD1.n24 B 0.025024f
C41 VDD1.n25 B 0.014976f
C42 VDD1.n26 B 1.5163f
C43 VDD1.n27 B 0.02787f
C44 VDD1.n28 B 0.014976f
C45 VDD1.n29 B 0.015857f
C46 VDD1.n30 B 0.035398f
C47 VDD1.n31 B 0.035398f
C48 VDD1.n32 B 0.015857f
C49 VDD1.n33 B 0.014976f
C50 VDD1.n34 B 0.02787f
C51 VDD1.n35 B 0.02787f
C52 VDD1.n36 B 0.014976f
C53 VDD1.n37 B 0.015857f
C54 VDD1.n38 B 0.035398f
C55 VDD1.n39 B 0.035398f
C56 VDD1.n40 B 0.015857f
C57 VDD1.n41 B 0.014976f
C58 VDD1.n42 B 0.02787f
C59 VDD1.n43 B 0.02787f
C60 VDD1.n44 B 0.014976f
C61 VDD1.n45 B 0.015416f
C62 VDD1.n46 B 0.015416f
C63 VDD1.n47 B 0.035398f
C64 VDD1.n48 B 0.035398f
C65 VDD1.n49 B 0.015857f
C66 VDD1.n50 B 0.014976f
C67 VDD1.n51 B 0.02787f
C68 VDD1.n52 B 0.02787f
C69 VDD1.n53 B 0.014976f
C70 VDD1.n54 B 0.015857f
C71 VDD1.n55 B 0.035398f
C72 VDD1.n56 B 0.035398f
C73 VDD1.n57 B 0.015857f
C74 VDD1.n58 B 0.014976f
C75 VDD1.n59 B 0.02787f
C76 VDD1.n60 B 0.02787f
C77 VDD1.n61 B 0.014976f
C78 VDD1.n62 B 0.015857f
C79 VDD1.n63 B 0.035398f
C80 VDD1.n64 B 0.079623f
C81 VDD1.n65 B 0.015857f
C82 VDD1.n66 B 0.014976f
C83 VDD1.n67 B 0.066323f
C84 VDD1.n68 B 0.065505f
C85 VDD1.t2 B 0.283883f
C86 VDD1.t7 B 0.283883f
C87 VDD1.n69 B 2.54107f
C88 VDD1.n70 B 0.415068f
C89 VDD1.n71 B 0.040866f
C90 VDD1.n72 B 0.02787f
C91 VDD1.n73 B 0.014976f
C92 VDD1.n74 B 0.035398f
C93 VDD1.n75 B 0.015857f
C94 VDD1.n76 B 0.02787f
C95 VDD1.n77 B 0.014976f
C96 VDD1.n78 B 0.035398f
C97 VDD1.n79 B 0.015857f
C98 VDD1.n80 B 0.02787f
C99 VDD1.n81 B 0.014976f
C100 VDD1.n82 B 0.035398f
C101 VDD1.n83 B 0.015857f
C102 VDD1.n84 B 0.02787f
C103 VDD1.n85 B 0.014976f
C104 VDD1.n86 B 0.035398f
C105 VDD1.n87 B 0.015857f
C106 VDD1.n88 B 0.02787f
C107 VDD1.n89 B 0.014976f
C108 VDD1.n90 B 0.035398f
C109 VDD1.n91 B 0.015857f
C110 VDD1.n92 B 0.21046f
C111 VDD1.t4 B 0.059918f
C112 VDD1.n93 B 0.026548f
C113 VDD1.n94 B 0.025024f
C114 VDD1.n95 B 0.014976f
C115 VDD1.n96 B 1.5163f
C116 VDD1.n97 B 0.02787f
C117 VDD1.n98 B 0.014976f
C118 VDD1.n99 B 0.015857f
C119 VDD1.n100 B 0.035398f
C120 VDD1.n101 B 0.035398f
C121 VDD1.n102 B 0.015857f
C122 VDD1.n103 B 0.014976f
C123 VDD1.n104 B 0.02787f
C124 VDD1.n105 B 0.02787f
C125 VDD1.n106 B 0.014976f
C126 VDD1.n107 B 0.015857f
C127 VDD1.n108 B 0.035398f
C128 VDD1.n109 B 0.035398f
C129 VDD1.n110 B 0.035398f
C130 VDD1.n111 B 0.015857f
C131 VDD1.n112 B 0.014976f
C132 VDD1.n113 B 0.02787f
C133 VDD1.n114 B 0.02787f
C134 VDD1.n115 B 0.014976f
C135 VDD1.n116 B 0.015416f
C136 VDD1.n117 B 0.015416f
C137 VDD1.n118 B 0.035398f
C138 VDD1.n119 B 0.035398f
C139 VDD1.n120 B 0.015857f
C140 VDD1.n121 B 0.014976f
C141 VDD1.n122 B 0.02787f
C142 VDD1.n123 B 0.02787f
C143 VDD1.n124 B 0.014976f
C144 VDD1.n125 B 0.015857f
C145 VDD1.n126 B 0.035398f
C146 VDD1.n127 B 0.035398f
C147 VDD1.n128 B 0.015857f
C148 VDD1.n129 B 0.014976f
C149 VDD1.n130 B 0.02787f
C150 VDD1.n131 B 0.02787f
C151 VDD1.n132 B 0.014976f
C152 VDD1.n133 B 0.015857f
C153 VDD1.n134 B 0.035398f
C154 VDD1.n135 B 0.079623f
C155 VDD1.n136 B 0.015857f
C156 VDD1.n137 B 0.014976f
C157 VDD1.n138 B 0.066323f
C158 VDD1.n139 B 0.065505f
C159 VDD1.t5 B 0.283883f
C160 VDD1.t1 B 0.283883f
C161 VDD1.n140 B 2.54107f
C162 VDD1.n141 B 0.411347f
C163 VDD1.t0 B 0.283883f
C164 VDD1.t8 B 0.283883f
C165 VDD1.n142 B 2.54325f
C166 VDD1.n143 B 2.0754f
C167 VDD1.t3 B 0.283883f
C168 VDD1.t9 B 0.283883f
C169 VDD1.n144 B 2.54106f
C170 VDD1.n145 B 2.59663f
C171 VP.n0 B 0.051496f
C172 VP.t8 B 0.737494f
C173 VP.n1 B 0.288471f
C174 VP.n2 B 0.051496f
C175 VP.n3 B 0.051496f
C176 VP.t0 B 0.737494f
C177 VP.t6 B 0.737494f
C178 VP.t2 B 0.737494f
C179 VP.n4 B 0.288471f
C180 VP.t3 B 0.744269f
C181 VP.n5 B 0.290259f
C182 VP.t7 B 0.737494f
C183 VP.n6 B 0.305396f
C184 VP.n7 B 0.011685f
C185 VP.n8 B 0.162689f
C186 VP.n9 B 0.051496f
C187 VP.n10 B 0.011685f
C188 VP.n11 B 0.305396f
C189 VP.n12 B 0.296664f
C190 VP.n13 B 2.10837f
C191 VP.n14 B 2.15266f
C192 VP.t5 B 0.737494f
C193 VP.n15 B 0.296664f
C194 VP.t4 B 0.737494f
C195 VP.n16 B 0.305396f
C196 VP.n17 B 0.011685f
C197 VP.n18 B 0.051496f
C198 VP.n19 B 0.051496f
C199 VP.n20 B 0.011685f
C200 VP.t9 B 0.737494f
C201 VP.n21 B 0.305396f
C202 VP.t1 B 0.737494f
C203 VP.n22 B 0.296664f
C204 VP.n23 B 0.039907f
C205 VTAIL.t7 B 0.293081f
C206 VTAIL.t13 B 0.293081f
C207 VTAIL.n0 B 2.5389f
C208 VTAIL.n1 B 0.404809f
C209 VTAIL.n2 B 0.04219f
C210 VTAIL.n3 B 0.028773f
C211 VTAIL.n4 B 0.015461f
C212 VTAIL.n5 B 0.036545f
C213 VTAIL.n6 B 0.016371f
C214 VTAIL.n7 B 0.028773f
C215 VTAIL.n8 B 0.015461f
C216 VTAIL.n9 B 0.036545f
C217 VTAIL.n10 B 0.016371f
C218 VTAIL.n11 B 0.028773f
C219 VTAIL.n12 B 0.015461f
C220 VTAIL.n13 B 0.036545f
C221 VTAIL.n14 B 0.016371f
C222 VTAIL.n15 B 0.028773f
C223 VTAIL.n16 B 0.015461f
C224 VTAIL.n17 B 0.036545f
C225 VTAIL.n18 B 0.016371f
C226 VTAIL.n19 B 0.028773f
C227 VTAIL.n20 B 0.015461f
C228 VTAIL.n21 B 0.036545f
C229 VTAIL.n22 B 0.016371f
C230 VTAIL.n23 B 0.21728f
C231 VTAIL.t5 B 0.061859f
C232 VTAIL.n24 B 0.027409f
C233 VTAIL.n25 B 0.025834f
C234 VTAIL.n26 B 0.015461f
C235 VTAIL.n27 B 1.56544f
C236 VTAIL.n28 B 0.028773f
C237 VTAIL.n29 B 0.015461f
C238 VTAIL.n30 B 0.016371f
C239 VTAIL.n31 B 0.036545f
C240 VTAIL.n32 B 0.036545f
C241 VTAIL.n33 B 0.016371f
C242 VTAIL.n34 B 0.015461f
C243 VTAIL.n35 B 0.028773f
C244 VTAIL.n36 B 0.028773f
C245 VTAIL.n37 B 0.015461f
C246 VTAIL.n38 B 0.016371f
C247 VTAIL.n39 B 0.036545f
C248 VTAIL.n40 B 0.036545f
C249 VTAIL.n41 B 0.036545f
C250 VTAIL.n42 B 0.016371f
C251 VTAIL.n43 B 0.015461f
C252 VTAIL.n44 B 0.028773f
C253 VTAIL.n45 B 0.028773f
C254 VTAIL.n46 B 0.015461f
C255 VTAIL.n47 B 0.015916f
C256 VTAIL.n48 B 0.015916f
C257 VTAIL.n49 B 0.036545f
C258 VTAIL.n50 B 0.036545f
C259 VTAIL.n51 B 0.016371f
C260 VTAIL.n52 B 0.015461f
C261 VTAIL.n53 B 0.028773f
C262 VTAIL.n54 B 0.028773f
C263 VTAIL.n55 B 0.015461f
C264 VTAIL.n56 B 0.016371f
C265 VTAIL.n57 B 0.036545f
C266 VTAIL.n58 B 0.036545f
C267 VTAIL.n59 B 0.016371f
C268 VTAIL.n60 B 0.015461f
C269 VTAIL.n61 B 0.028773f
C270 VTAIL.n62 B 0.028773f
C271 VTAIL.n63 B 0.015461f
C272 VTAIL.n64 B 0.016371f
C273 VTAIL.n65 B 0.036545f
C274 VTAIL.n66 B 0.082203f
C275 VTAIL.n67 B 0.016371f
C276 VTAIL.n68 B 0.015461f
C277 VTAIL.n69 B 0.068472f
C278 VTAIL.n70 B 0.046373f
C279 VTAIL.n71 B 0.155561f
C280 VTAIL.t19 B 0.293081f
C281 VTAIL.t2 B 0.293081f
C282 VTAIL.n72 B 2.5389f
C283 VTAIL.n73 B 0.399014f
C284 VTAIL.t16 B 0.293081f
C285 VTAIL.t3 B 0.293081f
C286 VTAIL.n74 B 2.5389f
C287 VTAIL.n75 B 1.87763f
C288 VTAIL.t8 B 0.293081f
C289 VTAIL.t14 B 0.293081f
C290 VTAIL.n76 B 2.5389f
C291 VTAIL.n77 B 1.87763f
C292 VTAIL.t9 B 0.293081f
C293 VTAIL.t15 B 0.293081f
C294 VTAIL.n78 B 2.5389f
C295 VTAIL.n79 B 0.399011f
C296 VTAIL.n80 B 0.04219f
C297 VTAIL.n81 B 0.028773f
C298 VTAIL.n82 B 0.015461f
C299 VTAIL.n83 B 0.036545f
C300 VTAIL.n84 B 0.016371f
C301 VTAIL.n85 B 0.028773f
C302 VTAIL.n86 B 0.015461f
C303 VTAIL.n87 B 0.036545f
C304 VTAIL.n88 B 0.016371f
C305 VTAIL.n89 B 0.028773f
C306 VTAIL.n90 B 0.015461f
C307 VTAIL.n91 B 0.036545f
C308 VTAIL.n92 B 0.016371f
C309 VTAIL.n93 B 0.028773f
C310 VTAIL.n94 B 0.015461f
C311 VTAIL.n95 B 0.036545f
C312 VTAIL.n96 B 0.036545f
C313 VTAIL.n97 B 0.016371f
C314 VTAIL.n98 B 0.028773f
C315 VTAIL.n99 B 0.015461f
C316 VTAIL.n100 B 0.036545f
C317 VTAIL.n101 B 0.016371f
C318 VTAIL.n102 B 0.21728f
C319 VTAIL.t10 B 0.061859f
C320 VTAIL.n103 B 0.027409f
C321 VTAIL.n104 B 0.025834f
C322 VTAIL.n105 B 0.015461f
C323 VTAIL.n106 B 1.56544f
C324 VTAIL.n107 B 0.028773f
C325 VTAIL.n108 B 0.015461f
C326 VTAIL.n109 B 0.016371f
C327 VTAIL.n110 B 0.036545f
C328 VTAIL.n111 B 0.036545f
C329 VTAIL.n112 B 0.016371f
C330 VTAIL.n113 B 0.015461f
C331 VTAIL.n114 B 0.028773f
C332 VTAIL.n115 B 0.028773f
C333 VTAIL.n116 B 0.015461f
C334 VTAIL.n117 B 0.016371f
C335 VTAIL.n118 B 0.036545f
C336 VTAIL.n119 B 0.036545f
C337 VTAIL.n120 B 0.016371f
C338 VTAIL.n121 B 0.015461f
C339 VTAIL.n122 B 0.028773f
C340 VTAIL.n123 B 0.028773f
C341 VTAIL.n124 B 0.015461f
C342 VTAIL.n125 B 0.015916f
C343 VTAIL.n126 B 0.015916f
C344 VTAIL.n127 B 0.036545f
C345 VTAIL.n128 B 0.036545f
C346 VTAIL.n129 B 0.016371f
C347 VTAIL.n130 B 0.015461f
C348 VTAIL.n131 B 0.028773f
C349 VTAIL.n132 B 0.028773f
C350 VTAIL.n133 B 0.015461f
C351 VTAIL.n134 B 0.016371f
C352 VTAIL.n135 B 0.036545f
C353 VTAIL.n136 B 0.036545f
C354 VTAIL.n137 B 0.016371f
C355 VTAIL.n138 B 0.015461f
C356 VTAIL.n139 B 0.028773f
C357 VTAIL.n140 B 0.028773f
C358 VTAIL.n141 B 0.015461f
C359 VTAIL.n142 B 0.016371f
C360 VTAIL.n143 B 0.036545f
C361 VTAIL.n144 B 0.082203f
C362 VTAIL.n145 B 0.016371f
C363 VTAIL.n146 B 0.015461f
C364 VTAIL.n147 B 0.068472f
C365 VTAIL.n148 B 0.046373f
C366 VTAIL.n149 B 0.155561f
C367 VTAIL.t4 B 0.293081f
C368 VTAIL.t18 B 0.293081f
C369 VTAIL.n150 B 2.5389f
C370 VTAIL.n151 B 0.413797f
C371 VTAIL.t1 B 0.293081f
C372 VTAIL.t17 B 0.293081f
C373 VTAIL.n152 B 2.5389f
C374 VTAIL.n153 B 0.399011f
C375 VTAIL.n154 B 0.04219f
C376 VTAIL.n155 B 0.028773f
C377 VTAIL.n156 B 0.015461f
C378 VTAIL.n157 B 0.036545f
C379 VTAIL.n158 B 0.016371f
C380 VTAIL.n159 B 0.028773f
C381 VTAIL.n160 B 0.015461f
C382 VTAIL.n161 B 0.036545f
C383 VTAIL.n162 B 0.016371f
C384 VTAIL.n163 B 0.028773f
C385 VTAIL.n164 B 0.015461f
C386 VTAIL.n165 B 0.036545f
C387 VTAIL.n166 B 0.016371f
C388 VTAIL.n167 B 0.028773f
C389 VTAIL.n168 B 0.015461f
C390 VTAIL.n169 B 0.036545f
C391 VTAIL.n170 B 0.036545f
C392 VTAIL.n171 B 0.016371f
C393 VTAIL.n172 B 0.028773f
C394 VTAIL.n173 B 0.015461f
C395 VTAIL.n174 B 0.036545f
C396 VTAIL.n175 B 0.016371f
C397 VTAIL.n176 B 0.21728f
C398 VTAIL.t0 B 0.061859f
C399 VTAIL.n177 B 0.027409f
C400 VTAIL.n178 B 0.025834f
C401 VTAIL.n179 B 0.015461f
C402 VTAIL.n180 B 1.56544f
C403 VTAIL.n181 B 0.028773f
C404 VTAIL.n182 B 0.015461f
C405 VTAIL.n183 B 0.016371f
C406 VTAIL.n184 B 0.036545f
C407 VTAIL.n185 B 0.036545f
C408 VTAIL.n186 B 0.016371f
C409 VTAIL.n187 B 0.015461f
C410 VTAIL.n188 B 0.028773f
C411 VTAIL.n189 B 0.028773f
C412 VTAIL.n190 B 0.015461f
C413 VTAIL.n191 B 0.016371f
C414 VTAIL.n192 B 0.036545f
C415 VTAIL.n193 B 0.036545f
C416 VTAIL.n194 B 0.016371f
C417 VTAIL.n195 B 0.015461f
C418 VTAIL.n196 B 0.028773f
C419 VTAIL.n197 B 0.028773f
C420 VTAIL.n198 B 0.015461f
C421 VTAIL.n199 B 0.015916f
C422 VTAIL.n200 B 0.015916f
C423 VTAIL.n201 B 0.036545f
C424 VTAIL.n202 B 0.036545f
C425 VTAIL.n203 B 0.016371f
C426 VTAIL.n204 B 0.015461f
C427 VTAIL.n205 B 0.028773f
C428 VTAIL.n206 B 0.028773f
C429 VTAIL.n207 B 0.015461f
C430 VTAIL.n208 B 0.016371f
C431 VTAIL.n209 B 0.036545f
C432 VTAIL.n210 B 0.036545f
C433 VTAIL.n211 B 0.016371f
C434 VTAIL.n212 B 0.015461f
C435 VTAIL.n213 B 0.028773f
C436 VTAIL.n214 B 0.028773f
C437 VTAIL.n215 B 0.015461f
C438 VTAIL.n216 B 0.016371f
C439 VTAIL.n217 B 0.036545f
C440 VTAIL.n218 B 0.082203f
C441 VTAIL.n219 B 0.016371f
C442 VTAIL.n220 B 0.015461f
C443 VTAIL.n221 B 0.068472f
C444 VTAIL.n222 B 0.046373f
C445 VTAIL.n223 B 1.56185f
C446 VTAIL.n224 B 0.04219f
C447 VTAIL.n225 B 0.028773f
C448 VTAIL.n226 B 0.015461f
C449 VTAIL.n227 B 0.036545f
C450 VTAIL.n228 B 0.016371f
C451 VTAIL.n229 B 0.028773f
C452 VTAIL.n230 B 0.015461f
C453 VTAIL.n231 B 0.036545f
C454 VTAIL.n232 B 0.016371f
C455 VTAIL.n233 B 0.028773f
C456 VTAIL.n234 B 0.015461f
C457 VTAIL.n235 B 0.036545f
C458 VTAIL.n236 B 0.016371f
C459 VTAIL.n237 B 0.028773f
C460 VTAIL.n238 B 0.015461f
C461 VTAIL.n239 B 0.036545f
C462 VTAIL.n240 B 0.016371f
C463 VTAIL.n241 B 0.028773f
C464 VTAIL.n242 B 0.015461f
C465 VTAIL.n243 B 0.036545f
C466 VTAIL.n244 B 0.016371f
C467 VTAIL.n245 B 0.21728f
C468 VTAIL.t11 B 0.061859f
C469 VTAIL.n246 B 0.027409f
C470 VTAIL.n247 B 0.025834f
C471 VTAIL.n248 B 0.015461f
C472 VTAIL.n249 B 1.56544f
C473 VTAIL.n250 B 0.028773f
C474 VTAIL.n251 B 0.015461f
C475 VTAIL.n252 B 0.016371f
C476 VTAIL.n253 B 0.036545f
C477 VTAIL.n254 B 0.036545f
C478 VTAIL.n255 B 0.016371f
C479 VTAIL.n256 B 0.015461f
C480 VTAIL.n257 B 0.028773f
C481 VTAIL.n258 B 0.028773f
C482 VTAIL.n259 B 0.015461f
C483 VTAIL.n260 B 0.016371f
C484 VTAIL.n261 B 0.036545f
C485 VTAIL.n262 B 0.036545f
C486 VTAIL.n263 B 0.036545f
C487 VTAIL.n264 B 0.016371f
C488 VTAIL.n265 B 0.015461f
C489 VTAIL.n266 B 0.028773f
C490 VTAIL.n267 B 0.028773f
C491 VTAIL.n268 B 0.015461f
C492 VTAIL.n269 B 0.015916f
C493 VTAIL.n270 B 0.015916f
C494 VTAIL.n271 B 0.036545f
C495 VTAIL.n272 B 0.036545f
C496 VTAIL.n273 B 0.016371f
C497 VTAIL.n274 B 0.015461f
C498 VTAIL.n275 B 0.028773f
C499 VTAIL.n276 B 0.028773f
C500 VTAIL.n277 B 0.015461f
C501 VTAIL.n278 B 0.016371f
C502 VTAIL.n279 B 0.036545f
C503 VTAIL.n280 B 0.036545f
C504 VTAIL.n281 B 0.016371f
C505 VTAIL.n282 B 0.015461f
C506 VTAIL.n283 B 0.028773f
C507 VTAIL.n284 B 0.028773f
C508 VTAIL.n285 B 0.015461f
C509 VTAIL.n286 B 0.016371f
C510 VTAIL.n287 B 0.036545f
C511 VTAIL.n288 B 0.082203f
C512 VTAIL.n289 B 0.016371f
C513 VTAIL.n290 B 0.015461f
C514 VTAIL.n291 B 0.068472f
C515 VTAIL.n292 B 0.046373f
C516 VTAIL.n293 B 1.56184f
C517 VTAIL.t12 B 0.293081f
C518 VTAIL.t6 B 0.293081f
C519 VTAIL.n294 B 2.5389f
C520 VTAIL.n295 B 0.35046f
C521 VDD2.n0 B 0.040706f
C522 VDD2.n1 B 0.027761f
C523 VDD2.n2 B 0.014918f
C524 VDD2.n3 B 0.03526f
C525 VDD2.n4 B 0.015795f
C526 VDD2.n5 B 0.027761f
C527 VDD2.n6 B 0.014918f
C528 VDD2.n7 B 0.03526f
C529 VDD2.n8 B 0.015795f
C530 VDD2.n9 B 0.027761f
C531 VDD2.n10 B 0.014918f
C532 VDD2.n11 B 0.03526f
C533 VDD2.n12 B 0.015795f
C534 VDD2.n13 B 0.027761f
C535 VDD2.n14 B 0.014918f
C536 VDD2.n15 B 0.03526f
C537 VDD2.n16 B 0.015795f
C538 VDD2.n17 B 0.027761f
C539 VDD2.n18 B 0.014918f
C540 VDD2.n19 B 0.03526f
C541 VDD2.n20 B 0.015795f
C542 VDD2.n21 B 0.209639f
C543 VDD2.t3 B 0.059684f
C544 VDD2.n22 B 0.026445f
C545 VDD2.n23 B 0.024926f
C546 VDD2.n24 B 0.014918f
C547 VDD2.n25 B 1.51039f
C548 VDD2.n26 B 0.027761f
C549 VDD2.n27 B 0.014918f
C550 VDD2.n28 B 0.015795f
C551 VDD2.n29 B 0.03526f
C552 VDD2.n30 B 0.03526f
C553 VDD2.n31 B 0.015795f
C554 VDD2.n32 B 0.014918f
C555 VDD2.n33 B 0.027761f
C556 VDD2.n34 B 0.027761f
C557 VDD2.n35 B 0.014918f
C558 VDD2.n36 B 0.015795f
C559 VDD2.n37 B 0.03526f
C560 VDD2.n38 B 0.03526f
C561 VDD2.n39 B 0.03526f
C562 VDD2.n40 B 0.015795f
C563 VDD2.n41 B 0.014918f
C564 VDD2.n42 B 0.027761f
C565 VDD2.n43 B 0.027761f
C566 VDD2.n44 B 0.014918f
C567 VDD2.n45 B 0.015356f
C568 VDD2.n46 B 0.015356f
C569 VDD2.n47 B 0.03526f
C570 VDD2.n48 B 0.03526f
C571 VDD2.n49 B 0.015795f
C572 VDD2.n50 B 0.014918f
C573 VDD2.n51 B 0.027761f
C574 VDD2.n52 B 0.027761f
C575 VDD2.n53 B 0.014918f
C576 VDD2.n54 B 0.015795f
C577 VDD2.n55 B 0.03526f
C578 VDD2.n56 B 0.03526f
C579 VDD2.n57 B 0.015795f
C580 VDD2.n58 B 0.014918f
C581 VDD2.n59 B 0.027761f
C582 VDD2.n60 B 0.027761f
C583 VDD2.n61 B 0.014918f
C584 VDD2.n62 B 0.015795f
C585 VDD2.n63 B 0.03526f
C586 VDD2.n64 B 0.079312f
C587 VDD2.n65 B 0.015795f
C588 VDD2.n66 B 0.014918f
C589 VDD2.n67 B 0.066064f
C590 VDD2.n68 B 0.06525f
C591 VDD2.t0 B 0.282776f
C592 VDD2.t4 B 0.282776f
C593 VDD2.n69 B 2.53116f
C594 VDD2.n70 B 0.409743f
C595 VDD2.t8 B 0.282776f
C596 VDD2.t7 B 0.282776f
C597 VDD2.n71 B 2.53334f
C598 VDD2.n72 B 1.98954f
C599 VDD2.n73 B 0.040706f
C600 VDD2.n74 B 0.027761f
C601 VDD2.n75 B 0.014918f
C602 VDD2.n76 B 0.03526f
C603 VDD2.n77 B 0.015795f
C604 VDD2.n78 B 0.027761f
C605 VDD2.n79 B 0.014918f
C606 VDD2.n80 B 0.03526f
C607 VDD2.n81 B 0.015795f
C608 VDD2.n82 B 0.027761f
C609 VDD2.n83 B 0.014918f
C610 VDD2.n84 B 0.03526f
C611 VDD2.n85 B 0.015795f
C612 VDD2.n86 B 0.027761f
C613 VDD2.n87 B 0.014918f
C614 VDD2.n88 B 0.03526f
C615 VDD2.n89 B 0.03526f
C616 VDD2.n90 B 0.015795f
C617 VDD2.n91 B 0.027761f
C618 VDD2.n92 B 0.014918f
C619 VDD2.n93 B 0.03526f
C620 VDD2.n94 B 0.015795f
C621 VDD2.n95 B 0.209639f
C622 VDD2.t9 B 0.059684f
C623 VDD2.n96 B 0.026445f
C624 VDD2.n97 B 0.024926f
C625 VDD2.n98 B 0.014918f
C626 VDD2.n99 B 1.51039f
C627 VDD2.n100 B 0.027761f
C628 VDD2.n101 B 0.014918f
C629 VDD2.n102 B 0.015795f
C630 VDD2.n103 B 0.03526f
C631 VDD2.n104 B 0.03526f
C632 VDD2.n105 B 0.015795f
C633 VDD2.n106 B 0.014918f
C634 VDD2.n107 B 0.027761f
C635 VDD2.n108 B 0.027761f
C636 VDD2.n109 B 0.014918f
C637 VDD2.n110 B 0.015795f
C638 VDD2.n111 B 0.03526f
C639 VDD2.n112 B 0.03526f
C640 VDD2.n113 B 0.015795f
C641 VDD2.n114 B 0.014918f
C642 VDD2.n115 B 0.027761f
C643 VDD2.n116 B 0.027761f
C644 VDD2.n117 B 0.014918f
C645 VDD2.n118 B 0.015356f
C646 VDD2.n119 B 0.015356f
C647 VDD2.n120 B 0.03526f
C648 VDD2.n121 B 0.03526f
C649 VDD2.n122 B 0.015795f
C650 VDD2.n123 B 0.014918f
C651 VDD2.n124 B 0.027761f
C652 VDD2.n125 B 0.027761f
C653 VDD2.n126 B 0.014918f
C654 VDD2.n127 B 0.015795f
C655 VDD2.n128 B 0.03526f
C656 VDD2.n129 B 0.03526f
C657 VDD2.n130 B 0.015795f
C658 VDD2.n131 B 0.014918f
C659 VDD2.n132 B 0.027761f
C660 VDD2.n133 B 0.027761f
C661 VDD2.n134 B 0.014918f
C662 VDD2.n135 B 0.015795f
C663 VDD2.n136 B 0.03526f
C664 VDD2.n137 B 0.079312f
C665 VDD2.n138 B 0.015795f
C666 VDD2.n139 B 0.014918f
C667 VDD2.n140 B 0.066064f
C668 VDD2.n141 B 0.063896f
C669 VDD2.n142 B 2.33853f
C670 VDD2.t2 B 0.282776f
C671 VDD2.t6 B 0.282776f
C672 VDD2.n143 B 2.53116f
C673 VDD2.n144 B 0.30474f
C674 VDD2.t5 B 0.282776f
C675 VDD2.t1 B 0.282776f
C676 VDD2.n145 B 2.5333f
C677 VN.n0 B 0.050577f
C678 VN.t3 B 0.72434f
C679 VN.n1 B 0.283327f
C680 VN.t8 B 0.730995f
C681 VN.n2 B 0.285082f
C682 VN.t2 B 0.72434f
C683 VN.n3 B 0.299949f
C684 VN.n4 B 0.011477f
C685 VN.n5 B 0.159787f
C686 VN.n6 B 0.050577f
C687 VN.n7 B 0.011477f
C688 VN.t9 B 0.72434f
C689 VN.n8 B 0.299949f
C690 VN.t4 B 0.72434f
C691 VN.n9 B 0.291373f
C692 VN.n10 B 0.039195f
C693 VN.n11 B 0.050577f
C694 VN.t6 B 0.72434f
C695 VN.n12 B 0.283327f
C696 VN.t5 B 0.730995f
C697 VN.n13 B 0.285082f
C698 VN.t0 B 0.72434f
C699 VN.n14 B 0.299949f
C700 VN.n15 B 0.011477f
C701 VN.n16 B 0.159787f
C702 VN.n17 B 0.050577f
C703 VN.n18 B 0.011477f
C704 VN.t1 B 0.72434f
C705 VN.n19 B 0.299949f
C706 VN.t7 B 0.72434f
C707 VN.n20 B 0.291373f
C708 VN.n21 B 2.10398f
.ends

