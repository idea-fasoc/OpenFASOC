* NGSPICE file created from diff_pair_sample_1683.ext - technology: sky130A

.subckt diff_pair_sample_1683 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=4.7931 ps=25.36 w=12.29 l=2.38
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=0 ps=0 w=12.29 l=2.38
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=0 ps=0 w=12.29 l=2.38
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=0 ps=0 w=12.29 l=2.38
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=4.7931 ps=25.36 w=12.29 l=2.38
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=0 ps=0 w=12.29 l=2.38
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=4.7931 ps=25.36 w=12.29 l=2.38
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7931 pd=25.36 as=4.7931 ps=25.36 w=12.29 l=2.38
R0 VP.n0 VP.t1 217.912
R1 VP.n0 VP.t0 173.619
R2 VP VP.n0 0.336784
R3 VTAIL.n1 VTAIL.t1 49.473
R4 VTAIL.n3 VTAIL.t0 49.4719
R5 VTAIL.n0 VTAIL.t3 49.4719
R6 VTAIL.n2 VTAIL.t2 49.4718
R7 VTAIL.n1 VTAIL.n0 27.6341
R8 VTAIL.n3 VTAIL.n2 25.2979
R9 VTAIL.n2 VTAIL.n1 1.63843
R10 VTAIL VTAIL.n0 1.11257
R11 VTAIL VTAIL.n3 0.526362
R12 VDD1 VDD1.t1 106.186
R13 VDD1 VDD1.t0 66.7928
R14 B.n680 B.n679 585
R15 B.n681 B.n680 585
R16 B.n286 B.n95 585
R17 B.n285 B.n284 585
R18 B.n283 B.n282 585
R19 B.n281 B.n280 585
R20 B.n279 B.n278 585
R21 B.n277 B.n276 585
R22 B.n275 B.n274 585
R23 B.n273 B.n272 585
R24 B.n271 B.n270 585
R25 B.n269 B.n268 585
R26 B.n267 B.n266 585
R27 B.n265 B.n264 585
R28 B.n263 B.n262 585
R29 B.n261 B.n260 585
R30 B.n259 B.n258 585
R31 B.n257 B.n256 585
R32 B.n255 B.n254 585
R33 B.n253 B.n252 585
R34 B.n251 B.n250 585
R35 B.n249 B.n248 585
R36 B.n247 B.n246 585
R37 B.n245 B.n244 585
R38 B.n243 B.n242 585
R39 B.n241 B.n240 585
R40 B.n239 B.n238 585
R41 B.n237 B.n236 585
R42 B.n235 B.n234 585
R43 B.n233 B.n232 585
R44 B.n231 B.n230 585
R45 B.n229 B.n228 585
R46 B.n227 B.n226 585
R47 B.n225 B.n224 585
R48 B.n223 B.n222 585
R49 B.n221 B.n220 585
R50 B.n219 B.n218 585
R51 B.n217 B.n216 585
R52 B.n215 B.n214 585
R53 B.n213 B.n212 585
R54 B.n211 B.n210 585
R55 B.n209 B.n208 585
R56 B.n207 B.n206 585
R57 B.n205 B.n204 585
R58 B.n203 B.n202 585
R59 B.n201 B.n200 585
R60 B.n199 B.n198 585
R61 B.n197 B.n196 585
R62 B.n195 B.n194 585
R63 B.n193 B.n192 585
R64 B.n191 B.n190 585
R65 B.n189 B.n188 585
R66 B.n187 B.n186 585
R67 B.n184 B.n183 585
R68 B.n182 B.n181 585
R69 B.n180 B.n179 585
R70 B.n178 B.n177 585
R71 B.n176 B.n175 585
R72 B.n174 B.n173 585
R73 B.n172 B.n171 585
R74 B.n170 B.n169 585
R75 B.n168 B.n167 585
R76 B.n166 B.n165 585
R77 B.n164 B.n163 585
R78 B.n162 B.n161 585
R79 B.n160 B.n159 585
R80 B.n158 B.n157 585
R81 B.n156 B.n155 585
R82 B.n154 B.n153 585
R83 B.n152 B.n151 585
R84 B.n150 B.n149 585
R85 B.n148 B.n147 585
R86 B.n146 B.n145 585
R87 B.n144 B.n143 585
R88 B.n142 B.n141 585
R89 B.n140 B.n139 585
R90 B.n138 B.n137 585
R91 B.n136 B.n135 585
R92 B.n134 B.n133 585
R93 B.n132 B.n131 585
R94 B.n130 B.n129 585
R95 B.n128 B.n127 585
R96 B.n126 B.n125 585
R97 B.n124 B.n123 585
R98 B.n122 B.n121 585
R99 B.n120 B.n119 585
R100 B.n118 B.n117 585
R101 B.n116 B.n115 585
R102 B.n114 B.n113 585
R103 B.n112 B.n111 585
R104 B.n110 B.n109 585
R105 B.n108 B.n107 585
R106 B.n106 B.n105 585
R107 B.n104 B.n103 585
R108 B.n102 B.n101 585
R109 B.n46 B.n45 585
R110 B.n678 B.n47 585
R111 B.n682 B.n47 585
R112 B.n677 B.n676 585
R113 B.n676 B.n43 585
R114 B.n675 B.n42 585
R115 B.n688 B.n42 585
R116 B.n674 B.n41 585
R117 B.n689 B.n41 585
R118 B.n673 B.n40 585
R119 B.n690 B.n40 585
R120 B.n672 B.n671 585
R121 B.n671 B.n36 585
R122 B.n670 B.n35 585
R123 B.n696 B.n35 585
R124 B.n669 B.n34 585
R125 B.n697 B.n34 585
R126 B.n668 B.n33 585
R127 B.n698 B.n33 585
R128 B.n667 B.n666 585
R129 B.n666 B.n29 585
R130 B.n665 B.n28 585
R131 B.n704 B.n28 585
R132 B.n664 B.n27 585
R133 B.n705 B.n27 585
R134 B.n663 B.n26 585
R135 B.n706 B.n26 585
R136 B.n662 B.n661 585
R137 B.n661 B.n22 585
R138 B.n660 B.n21 585
R139 B.n712 B.n21 585
R140 B.n659 B.n20 585
R141 B.n713 B.n20 585
R142 B.n658 B.n19 585
R143 B.n714 B.n19 585
R144 B.n657 B.n656 585
R145 B.n656 B.n15 585
R146 B.n655 B.n14 585
R147 B.n720 B.n14 585
R148 B.n654 B.n13 585
R149 B.n721 B.n13 585
R150 B.n653 B.n12 585
R151 B.n722 B.n12 585
R152 B.n652 B.n651 585
R153 B.n651 B.n8 585
R154 B.n650 B.n7 585
R155 B.n728 B.n7 585
R156 B.n649 B.n6 585
R157 B.n729 B.n6 585
R158 B.n648 B.n5 585
R159 B.n730 B.n5 585
R160 B.n647 B.n646 585
R161 B.n646 B.n4 585
R162 B.n645 B.n287 585
R163 B.n645 B.n644 585
R164 B.n635 B.n288 585
R165 B.n289 B.n288 585
R166 B.n637 B.n636 585
R167 B.n638 B.n637 585
R168 B.n634 B.n294 585
R169 B.n294 B.n293 585
R170 B.n633 B.n632 585
R171 B.n632 B.n631 585
R172 B.n296 B.n295 585
R173 B.n297 B.n296 585
R174 B.n624 B.n623 585
R175 B.n625 B.n624 585
R176 B.n622 B.n302 585
R177 B.n302 B.n301 585
R178 B.n621 B.n620 585
R179 B.n620 B.n619 585
R180 B.n304 B.n303 585
R181 B.n305 B.n304 585
R182 B.n612 B.n611 585
R183 B.n613 B.n612 585
R184 B.n610 B.n310 585
R185 B.n310 B.n309 585
R186 B.n609 B.n608 585
R187 B.n608 B.n607 585
R188 B.n312 B.n311 585
R189 B.n313 B.n312 585
R190 B.n600 B.n599 585
R191 B.n601 B.n600 585
R192 B.n598 B.n317 585
R193 B.n321 B.n317 585
R194 B.n597 B.n596 585
R195 B.n596 B.n595 585
R196 B.n319 B.n318 585
R197 B.n320 B.n319 585
R198 B.n588 B.n587 585
R199 B.n589 B.n588 585
R200 B.n586 B.n326 585
R201 B.n326 B.n325 585
R202 B.n585 B.n584 585
R203 B.n584 B.n583 585
R204 B.n328 B.n327 585
R205 B.n329 B.n328 585
R206 B.n576 B.n575 585
R207 B.n577 B.n576 585
R208 B.n332 B.n331 585
R209 B.n385 B.n384 585
R210 B.n386 B.n382 585
R211 B.n382 B.n333 585
R212 B.n388 B.n387 585
R213 B.n390 B.n381 585
R214 B.n393 B.n392 585
R215 B.n394 B.n380 585
R216 B.n396 B.n395 585
R217 B.n398 B.n379 585
R218 B.n401 B.n400 585
R219 B.n402 B.n378 585
R220 B.n404 B.n403 585
R221 B.n406 B.n377 585
R222 B.n409 B.n408 585
R223 B.n410 B.n376 585
R224 B.n412 B.n411 585
R225 B.n414 B.n375 585
R226 B.n417 B.n416 585
R227 B.n418 B.n374 585
R228 B.n420 B.n419 585
R229 B.n422 B.n373 585
R230 B.n425 B.n424 585
R231 B.n426 B.n372 585
R232 B.n428 B.n427 585
R233 B.n430 B.n371 585
R234 B.n433 B.n432 585
R235 B.n434 B.n370 585
R236 B.n436 B.n435 585
R237 B.n438 B.n369 585
R238 B.n441 B.n440 585
R239 B.n442 B.n368 585
R240 B.n444 B.n443 585
R241 B.n446 B.n367 585
R242 B.n449 B.n448 585
R243 B.n450 B.n366 585
R244 B.n452 B.n451 585
R245 B.n454 B.n365 585
R246 B.n457 B.n456 585
R247 B.n458 B.n364 585
R248 B.n460 B.n459 585
R249 B.n462 B.n363 585
R250 B.n465 B.n464 585
R251 B.n466 B.n360 585
R252 B.n469 B.n468 585
R253 B.n471 B.n359 585
R254 B.n474 B.n473 585
R255 B.n475 B.n358 585
R256 B.n477 B.n476 585
R257 B.n479 B.n357 585
R258 B.n482 B.n481 585
R259 B.n483 B.n356 585
R260 B.n488 B.n487 585
R261 B.n490 B.n355 585
R262 B.n493 B.n492 585
R263 B.n494 B.n354 585
R264 B.n496 B.n495 585
R265 B.n498 B.n353 585
R266 B.n501 B.n500 585
R267 B.n502 B.n352 585
R268 B.n504 B.n503 585
R269 B.n506 B.n351 585
R270 B.n509 B.n508 585
R271 B.n510 B.n350 585
R272 B.n512 B.n511 585
R273 B.n514 B.n349 585
R274 B.n517 B.n516 585
R275 B.n518 B.n348 585
R276 B.n520 B.n519 585
R277 B.n522 B.n347 585
R278 B.n525 B.n524 585
R279 B.n526 B.n346 585
R280 B.n528 B.n527 585
R281 B.n530 B.n345 585
R282 B.n533 B.n532 585
R283 B.n534 B.n344 585
R284 B.n536 B.n535 585
R285 B.n538 B.n343 585
R286 B.n541 B.n540 585
R287 B.n542 B.n342 585
R288 B.n544 B.n543 585
R289 B.n546 B.n341 585
R290 B.n549 B.n548 585
R291 B.n550 B.n340 585
R292 B.n552 B.n551 585
R293 B.n554 B.n339 585
R294 B.n557 B.n556 585
R295 B.n558 B.n338 585
R296 B.n560 B.n559 585
R297 B.n562 B.n337 585
R298 B.n565 B.n564 585
R299 B.n566 B.n336 585
R300 B.n568 B.n567 585
R301 B.n570 B.n335 585
R302 B.n573 B.n572 585
R303 B.n574 B.n334 585
R304 B.n579 B.n578 585
R305 B.n578 B.n577 585
R306 B.n580 B.n330 585
R307 B.n330 B.n329 585
R308 B.n582 B.n581 585
R309 B.n583 B.n582 585
R310 B.n324 B.n323 585
R311 B.n325 B.n324 585
R312 B.n591 B.n590 585
R313 B.n590 B.n589 585
R314 B.n592 B.n322 585
R315 B.n322 B.n320 585
R316 B.n594 B.n593 585
R317 B.n595 B.n594 585
R318 B.n316 B.n315 585
R319 B.n321 B.n316 585
R320 B.n603 B.n602 585
R321 B.n602 B.n601 585
R322 B.n604 B.n314 585
R323 B.n314 B.n313 585
R324 B.n606 B.n605 585
R325 B.n607 B.n606 585
R326 B.n308 B.n307 585
R327 B.n309 B.n308 585
R328 B.n615 B.n614 585
R329 B.n614 B.n613 585
R330 B.n616 B.n306 585
R331 B.n306 B.n305 585
R332 B.n618 B.n617 585
R333 B.n619 B.n618 585
R334 B.n300 B.n299 585
R335 B.n301 B.n300 585
R336 B.n627 B.n626 585
R337 B.n626 B.n625 585
R338 B.n628 B.n298 585
R339 B.n298 B.n297 585
R340 B.n630 B.n629 585
R341 B.n631 B.n630 585
R342 B.n292 B.n291 585
R343 B.n293 B.n292 585
R344 B.n640 B.n639 585
R345 B.n639 B.n638 585
R346 B.n641 B.n290 585
R347 B.n290 B.n289 585
R348 B.n643 B.n642 585
R349 B.n644 B.n643 585
R350 B.n2 B.n0 585
R351 B.n4 B.n2 585
R352 B.n3 B.n1 585
R353 B.n729 B.n3 585
R354 B.n727 B.n726 585
R355 B.n728 B.n727 585
R356 B.n725 B.n9 585
R357 B.n9 B.n8 585
R358 B.n724 B.n723 585
R359 B.n723 B.n722 585
R360 B.n11 B.n10 585
R361 B.n721 B.n11 585
R362 B.n719 B.n718 585
R363 B.n720 B.n719 585
R364 B.n717 B.n16 585
R365 B.n16 B.n15 585
R366 B.n716 B.n715 585
R367 B.n715 B.n714 585
R368 B.n18 B.n17 585
R369 B.n713 B.n18 585
R370 B.n711 B.n710 585
R371 B.n712 B.n711 585
R372 B.n709 B.n23 585
R373 B.n23 B.n22 585
R374 B.n708 B.n707 585
R375 B.n707 B.n706 585
R376 B.n25 B.n24 585
R377 B.n705 B.n25 585
R378 B.n703 B.n702 585
R379 B.n704 B.n703 585
R380 B.n701 B.n30 585
R381 B.n30 B.n29 585
R382 B.n700 B.n699 585
R383 B.n699 B.n698 585
R384 B.n32 B.n31 585
R385 B.n697 B.n32 585
R386 B.n695 B.n694 585
R387 B.n696 B.n695 585
R388 B.n693 B.n37 585
R389 B.n37 B.n36 585
R390 B.n692 B.n691 585
R391 B.n691 B.n690 585
R392 B.n39 B.n38 585
R393 B.n689 B.n39 585
R394 B.n687 B.n686 585
R395 B.n688 B.n687 585
R396 B.n685 B.n44 585
R397 B.n44 B.n43 585
R398 B.n684 B.n683 585
R399 B.n683 B.n682 585
R400 B.n732 B.n731 585
R401 B.n731 B.n730 585
R402 B.n578 B.n332 468.476
R403 B.n683 B.n46 468.476
R404 B.n576 B.n334 468.476
R405 B.n680 B.n47 468.476
R406 B.n484 B.t6 332.139
R407 B.n361 B.t10 332.139
R408 B.n99 B.t13 332.139
R409 B.n96 B.t2 332.139
R410 B.n681 B.n94 256.663
R411 B.n681 B.n93 256.663
R412 B.n681 B.n92 256.663
R413 B.n681 B.n91 256.663
R414 B.n681 B.n90 256.663
R415 B.n681 B.n89 256.663
R416 B.n681 B.n88 256.663
R417 B.n681 B.n87 256.663
R418 B.n681 B.n86 256.663
R419 B.n681 B.n85 256.663
R420 B.n681 B.n84 256.663
R421 B.n681 B.n83 256.663
R422 B.n681 B.n82 256.663
R423 B.n681 B.n81 256.663
R424 B.n681 B.n80 256.663
R425 B.n681 B.n79 256.663
R426 B.n681 B.n78 256.663
R427 B.n681 B.n77 256.663
R428 B.n681 B.n76 256.663
R429 B.n681 B.n75 256.663
R430 B.n681 B.n74 256.663
R431 B.n681 B.n73 256.663
R432 B.n681 B.n72 256.663
R433 B.n681 B.n71 256.663
R434 B.n681 B.n70 256.663
R435 B.n681 B.n69 256.663
R436 B.n681 B.n68 256.663
R437 B.n681 B.n67 256.663
R438 B.n681 B.n66 256.663
R439 B.n681 B.n65 256.663
R440 B.n681 B.n64 256.663
R441 B.n681 B.n63 256.663
R442 B.n681 B.n62 256.663
R443 B.n681 B.n61 256.663
R444 B.n681 B.n60 256.663
R445 B.n681 B.n59 256.663
R446 B.n681 B.n58 256.663
R447 B.n681 B.n57 256.663
R448 B.n681 B.n56 256.663
R449 B.n681 B.n55 256.663
R450 B.n681 B.n54 256.663
R451 B.n681 B.n53 256.663
R452 B.n681 B.n52 256.663
R453 B.n681 B.n51 256.663
R454 B.n681 B.n50 256.663
R455 B.n681 B.n49 256.663
R456 B.n681 B.n48 256.663
R457 B.n383 B.n333 256.663
R458 B.n389 B.n333 256.663
R459 B.n391 B.n333 256.663
R460 B.n397 B.n333 256.663
R461 B.n399 B.n333 256.663
R462 B.n405 B.n333 256.663
R463 B.n407 B.n333 256.663
R464 B.n413 B.n333 256.663
R465 B.n415 B.n333 256.663
R466 B.n421 B.n333 256.663
R467 B.n423 B.n333 256.663
R468 B.n429 B.n333 256.663
R469 B.n431 B.n333 256.663
R470 B.n437 B.n333 256.663
R471 B.n439 B.n333 256.663
R472 B.n445 B.n333 256.663
R473 B.n447 B.n333 256.663
R474 B.n453 B.n333 256.663
R475 B.n455 B.n333 256.663
R476 B.n461 B.n333 256.663
R477 B.n463 B.n333 256.663
R478 B.n470 B.n333 256.663
R479 B.n472 B.n333 256.663
R480 B.n478 B.n333 256.663
R481 B.n480 B.n333 256.663
R482 B.n489 B.n333 256.663
R483 B.n491 B.n333 256.663
R484 B.n497 B.n333 256.663
R485 B.n499 B.n333 256.663
R486 B.n505 B.n333 256.663
R487 B.n507 B.n333 256.663
R488 B.n513 B.n333 256.663
R489 B.n515 B.n333 256.663
R490 B.n521 B.n333 256.663
R491 B.n523 B.n333 256.663
R492 B.n529 B.n333 256.663
R493 B.n531 B.n333 256.663
R494 B.n537 B.n333 256.663
R495 B.n539 B.n333 256.663
R496 B.n545 B.n333 256.663
R497 B.n547 B.n333 256.663
R498 B.n553 B.n333 256.663
R499 B.n555 B.n333 256.663
R500 B.n561 B.n333 256.663
R501 B.n563 B.n333 256.663
R502 B.n569 B.n333 256.663
R503 B.n571 B.n333 256.663
R504 B.n578 B.n330 163.367
R505 B.n582 B.n330 163.367
R506 B.n582 B.n324 163.367
R507 B.n590 B.n324 163.367
R508 B.n590 B.n322 163.367
R509 B.n594 B.n322 163.367
R510 B.n594 B.n316 163.367
R511 B.n602 B.n316 163.367
R512 B.n602 B.n314 163.367
R513 B.n606 B.n314 163.367
R514 B.n606 B.n308 163.367
R515 B.n614 B.n308 163.367
R516 B.n614 B.n306 163.367
R517 B.n618 B.n306 163.367
R518 B.n618 B.n300 163.367
R519 B.n626 B.n300 163.367
R520 B.n626 B.n298 163.367
R521 B.n630 B.n298 163.367
R522 B.n630 B.n292 163.367
R523 B.n639 B.n292 163.367
R524 B.n639 B.n290 163.367
R525 B.n643 B.n290 163.367
R526 B.n643 B.n2 163.367
R527 B.n731 B.n2 163.367
R528 B.n731 B.n3 163.367
R529 B.n727 B.n3 163.367
R530 B.n727 B.n9 163.367
R531 B.n723 B.n9 163.367
R532 B.n723 B.n11 163.367
R533 B.n719 B.n11 163.367
R534 B.n719 B.n16 163.367
R535 B.n715 B.n16 163.367
R536 B.n715 B.n18 163.367
R537 B.n711 B.n18 163.367
R538 B.n711 B.n23 163.367
R539 B.n707 B.n23 163.367
R540 B.n707 B.n25 163.367
R541 B.n703 B.n25 163.367
R542 B.n703 B.n30 163.367
R543 B.n699 B.n30 163.367
R544 B.n699 B.n32 163.367
R545 B.n695 B.n32 163.367
R546 B.n695 B.n37 163.367
R547 B.n691 B.n37 163.367
R548 B.n691 B.n39 163.367
R549 B.n687 B.n39 163.367
R550 B.n687 B.n44 163.367
R551 B.n683 B.n44 163.367
R552 B.n384 B.n382 163.367
R553 B.n388 B.n382 163.367
R554 B.n392 B.n390 163.367
R555 B.n396 B.n380 163.367
R556 B.n400 B.n398 163.367
R557 B.n404 B.n378 163.367
R558 B.n408 B.n406 163.367
R559 B.n412 B.n376 163.367
R560 B.n416 B.n414 163.367
R561 B.n420 B.n374 163.367
R562 B.n424 B.n422 163.367
R563 B.n428 B.n372 163.367
R564 B.n432 B.n430 163.367
R565 B.n436 B.n370 163.367
R566 B.n440 B.n438 163.367
R567 B.n444 B.n368 163.367
R568 B.n448 B.n446 163.367
R569 B.n452 B.n366 163.367
R570 B.n456 B.n454 163.367
R571 B.n460 B.n364 163.367
R572 B.n464 B.n462 163.367
R573 B.n469 B.n360 163.367
R574 B.n473 B.n471 163.367
R575 B.n477 B.n358 163.367
R576 B.n481 B.n479 163.367
R577 B.n488 B.n356 163.367
R578 B.n492 B.n490 163.367
R579 B.n496 B.n354 163.367
R580 B.n500 B.n498 163.367
R581 B.n504 B.n352 163.367
R582 B.n508 B.n506 163.367
R583 B.n512 B.n350 163.367
R584 B.n516 B.n514 163.367
R585 B.n520 B.n348 163.367
R586 B.n524 B.n522 163.367
R587 B.n528 B.n346 163.367
R588 B.n532 B.n530 163.367
R589 B.n536 B.n344 163.367
R590 B.n540 B.n538 163.367
R591 B.n544 B.n342 163.367
R592 B.n548 B.n546 163.367
R593 B.n552 B.n340 163.367
R594 B.n556 B.n554 163.367
R595 B.n560 B.n338 163.367
R596 B.n564 B.n562 163.367
R597 B.n568 B.n336 163.367
R598 B.n572 B.n570 163.367
R599 B.n576 B.n328 163.367
R600 B.n584 B.n328 163.367
R601 B.n584 B.n326 163.367
R602 B.n588 B.n326 163.367
R603 B.n588 B.n319 163.367
R604 B.n596 B.n319 163.367
R605 B.n596 B.n317 163.367
R606 B.n600 B.n317 163.367
R607 B.n600 B.n312 163.367
R608 B.n608 B.n312 163.367
R609 B.n608 B.n310 163.367
R610 B.n612 B.n310 163.367
R611 B.n612 B.n304 163.367
R612 B.n620 B.n304 163.367
R613 B.n620 B.n302 163.367
R614 B.n624 B.n302 163.367
R615 B.n624 B.n296 163.367
R616 B.n632 B.n296 163.367
R617 B.n632 B.n294 163.367
R618 B.n637 B.n294 163.367
R619 B.n637 B.n288 163.367
R620 B.n645 B.n288 163.367
R621 B.n646 B.n645 163.367
R622 B.n646 B.n5 163.367
R623 B.n6 B.n5 163.367
R624 B.n7 B.n6 163.367
R625 B.n651 B.n7 163.367
R626 B.n651 B.n12 163.367
R627 B.n13 B.n12 163.367
R628 B.n14 B.n13 163.367
R629 B.n656 B.n14 163.367
R630 B.n656 B.n19 163.367
R631 B.n20 B.n19 163.367
R632 B.n21 B.n20 163.367
R633 B.n661 B.n21 163.367
R634 B.n661 B.n26 163.367
R635 B.n27 B.n26 163.367
R636 B.n28 B.n27 163.367
R637 B.n666 B.n28 163.367
R638 B.n666 B.n33 163.367
R639 B.n34 B.n33 163.367
R640 B.n35 B.n34 163.367
R641 B.n671 B.n35 163.367
R642 B.n671 B.n40 163.367
R643 B.n41 B.n40 163.367
R644 B.n42 B.n41 163.367
R645 B.n676 B.n42 163.367
R646 B.n676 B.n47 163.367
R647 B.n103 B.n102 163.367
R648 B.n107 B.n106 163.367
R649 B.n111 B.n110 163.367
R650 B.n115 B.n114 163.367
R651 B.n119 B.n118 163.367
R652 B.n123 B.n122 163.367
R653 B.n127 B.n126 163.367
R654 B.n131 B.n130 163.367
R655 B.n135 B.n134 163.367
R656 B.n139 B.n138 163.367
R657 B.n143 B.n142 163.367
R658 B.n147 B.n146 163.367
R659 B.n151 B.n150 163.367
R660 B.n155 B.n154 163.367
R661 B.n159 B.n158 163.367
R662 B.n163 B.n162 163.367
R663 B.n167 B.n166 163.367
R664 B.n171 B.n170 163.367
R665 B.n175 B.n174 163.367
R666 B.n179 B.n178 163.367
R667 B.n183 B.n182 163.367
R668 B.n188 B.n187 163.367
R669 B.n192 B.n191 163.367
R670 B.n196 B.n195 163.367
R671 B.n200 B.n199 163.367
R672 B.n204 B.n203 163.367
R673 B.n208 B.n207 163.367
R674 B.n212 B.n211 163.367
R675 B.n216 B.n215 163.367
R676 B.n220 B.n219 163.367
R677 B.n224 B.n223 163.367
R678 B.n228 B.n227 163.367
R679 B.n232 B.n231 163.367
R680 B.n236 B.n235 163.367
R681 B.n240 B.n239 163.367
R682 B.n244 B.n243 163.367
R683 B.n248 B.n247 163.367
R684 B.n252 B.n251 163.367
R685 B.n256 B.n255 163.367
R686 B.n260 B.n259 163.367
R687 B.n264 B.n263 163.367
R688 B.n268 B.n267 163.367
R689 B.n272 B.n271 163.367
R690 B.n276 B.n275 163.367
R691 B.n280 B.n279 163.367
R692 B.n284 B.n283 163.367
R693 B.n680 B.n95 163.367
R694 B.n484 B.t9 121.278
R695 B.n96 B.t4 121.278
R696 B.n361 B.t12 121.263
R697 B.n99 B.t14 121.263
R698 B.n577 B.n333 79.5337
R699 B.n682 B.n681 79.5337
R700 B.n383 B.n332 71.676
R701 B.n389 B.n388 71.676
R702 B.n392 B.n391 71.676
R703 B.n397 B.n396 71.676
R704 B.n400 B.n399 71.676
R705 B.n405 B.n404 71.676
R706 B.n408 B.n407 71.676
R707 B.n413 B.n412 71.676
R708 B.n416 B.n415 71.676
R709 B.n421 B.n420 71.676
R710 B.n424 B.n423 71.676
R711 B.n429 B.n428 71.676
R712 B.n432 B.n431 71.676
R713 B.n437 B.n436 71.676
R714 B.n440 B.n439 71.676
R715 B.n445 B.n444 71.676
R716 B.n448 B.n447 71.676
R717 B.n453 B.n452 71.676
R718 B.n456 B.n455 71.676
R719 B.n461 B.n460 71.676
R720 B.n464 B.n463 71.676
R721 B.n470 B.n469 71.676
R722 B.n473 B.n472 71.676
R723 B.n478 B.n477 71.676
R724 B.n481 B.n480 71.676
R725 B.n489 B.n488 71.676
R726 B.n492 B.n491 71.676
R727 B.n497 B.n496 71.676
R728 B.n500 B.n499 71.676
R729 B.n505 B.n504 71.676
R730 B.n508 B.n507 71.676
R731 B.n513 B.n512 71.676
R732 B.n516 B.n515 71.676
R733 B.n521 B.n520 71.676
R734 B.n524 B.n523 71.676
R735 B.n529 B.n528 71.676
R736 B.n532 B.n531 71.676
R737 B.n537 B.n536 71.676
R738 B.n540 B.n539 71.676
R739 B.n545 B.n544 71.676
R740 B.n548 B.n547 71.676
R741 B.n553 B.n552 71.676
R742 B.n556 B.n555 71.676
R743 B.n561 B.n560 71.676
R744 B.n564 B.n563 71.676
R745 B.n569 B.n568 71.676
R746 B.n572 B.n571 71.676
R747 B.n48 B.n46 71.676
R748 B.n103 B.n49 71.676
R749 B.n107 B.n50 71.676
R750 B.n111 B.n51 71.676
R751 B.n115 B.n52 71.676
R752 B.n119 B.n53 71.676
R753 B.n123 B.n54 71.676
R754 B.n127 B.n55 71.676
R755 B.n131 B.n56 71.676
R756 B.n135 B.n57 71.676
R757 B.n139 B.n58 71.676
R758 B.n143 B.n59 71.676
R759 B.n147 B.n60 71.676
R760 B.n151 B.n61 71.676
R761 B.n155 B.n62 71.676
R762 B.n159 B.n63 71.676
R763 B.n163 B.n64 71.676
R764 B.n167 B.n65 71.676
R765 B.n171 B.n66 71.676
R766 B.n175 B.n67 71.676
R767 B.n179 B.n68 71.676
R768 B.n183 B.n69 71.676
R769 B.n188 B.n70 71.676
R770 B.n192 B.n71 71.676
R771 B.n196 B.n72 71.676
R772 B.n200 B.n73 71.676
R773 B.n204 B.n74 71.676
R774 B.n208 B.n75 71.676
R775 B.n212 B.n76 71.676
R776 B.n216 B.n77 71.676
R777 B.n220 B.n78 71.676
R778 B.n224 B.n79 71.676
R779 B.n228 B.n80 71.676
R780 B.n232 B.n81 71.676
R781 B.n236 B.n82 71.676
R782 B.n240 B.n83 71.676
R783 B.n244 B.n84 71.676
R784 B.n248 B.n85 71.676
R785 B.n252 B.n86 71.676
R786 B.n256 B.n87 71.676
R787 B.n260 B.n88 71.676
R788 B.n264 B.n89 71.676
R789 B.n268 B.n90 71.676
R790 B.n272 B.n91 71.676
R791 B.n276 B.n92 71.676
R792 B.n280 B.n93 71.676
R793 B.n284 B.n94 71.676
R794 B.n95 B.n94 71.676
R795 B.n283 B.n93 71.676
R796 B.n279 B.n92 71.676
R797 B.n275 B.n91 71.676
R798 B.n271 B.n90 71.676
R799 B.n267 B.n89 71.676
R800 B.n263 B.n88 71.676
R801 B.n259 B.n87 71.676
R802 B.n255 B.n86 71.676
R803 B.n251 B.n85 71.676
R804 B.n247 B.n84 71.676
R805 B.n243 B.n83 71.676
R806 B.n239 B.n82 71.676
R807 B.n235 B.n81 71.676
R808 B.n231 B.n80 71.676
R809 B.n227 B.n79 71.676
R810 B.n223 B.n78 71.676
R811 B.n219 B.n77 71.676
R812 B.n215 B.n76 71.676
R813 B.n211 B.n75 71.676
R814 B.n207 B.n74 71.676
R815 B.n203 B.n73 71.676
R816 B.n199 B.n72 71.676
R817 B.n195 B.n71 71.676
R818 B.n191 B.n70 71.676
R819 B.n187 B.n69 71.676
R820 B.n182 B.n68 71.676
R821 B.n178 B.n67 71.676
R822 B.n174 B.n66 71.676
R823 B.n170 B.n65 71.676
R824 B.n166 B.n64 71.676
R825 B.n162 B.n63 71.676
R826 B.n158 B.n62 71.676
R827 B.n154 B.n61 71.676
R828 B.n150 B.n60 71.676
R829 B.n146 B.n59 71.676
R830 B.n142 B.n58 71.676
R831 B.n138 B.n57 71.676
R832 B.n134 B.n56 71.676
R833 B.n130 B.n55 71.676
R834 B.n126 B.n54 71.676
R835 B.n122 B.n53 71.676
R836 B.n118 B.n52 71.676
R837 B.n114 B.n51 71.676
R838 B.n110 B.n50 71.676
R839 B.n106 B.n49 71.676
R840 B.n102 B.n48 71.676
R841 B.n384 B.n383 71.676
R842 B.n390 B.n389 71.676
R843 B.n391 B.n380 71.676
R844 B.n398 B.n397 71.676
R845 B.n399 B.n378 71.676
R846 B.n406 B.n405 71.676
R847 B.n407 B.n376 71.676
R848 B.n414 B.n413 71.676
R849 B.n415 B.n374 71.676
R850 B.n422 B.n421 71.676
R851 B.n423 B.n372 71.676
R852 B.n430 B.n429 71.676
R853 B.n431 B.n370 71.676
R854 B.n438 B.n437 71.676
R855 B.n439 B.n368 71.676
R856 B.n446 B.n445 71.676
R857 B.n447 B.n366 71.676
R858 B.n454 B.n453 71.676
R859 B.n455 B.n364 71.676
R860 B.n462 B.n461 71.676
R861 B.n463 B.n360 71.676
R862 B.n471 B.n470 71.676
R863 B.n472 B.n358 71.676
R864 B.n479 B.n478 71.676
R865 B.n480 B.n356 71.676
R866 B.n490 B.n489 71.676
R867 B.n491 B.n354 71.676
R868 B.n498 B.n497 71.676
R869 B.n499 B.n352 71.676
R870 B.n506 B.n505 71.676
R871 B.n507 B.n350 71.676
R872 B.n514 B.n513 71.676
R873 B.n515 B.n348 71.676
R874 B.n522 B.n521 71.676
R875 B.n523 B.n346 71.676
R876 B.n530 B.n529 71.676
R877 B.n531 B.n344 71.676
R878 B.n538 B.n537 71.676
R879 B.n539 B.n342 71.676
R880 B.n546 B.n545 71.676
R881 B.n547 B.n340 71.676
R882 B.n554 B.n553 71.676
R883 B.n555 B.n338 71.676
R884 B.n562 B.n561 71.676
R885 B.n563 B.n336 71.676
R886 B.n570 B.n569 71.676
R887 B.n571 B.n334 71.676
R888 B.n485 B.t8 68.7211
R889 B.n97 B.t5 68.7211
R890 B.n362 B.t11 68.7054
R891 B.n100 B.t15 68.7054
R892 B.n486 B.n485 59.5399
R893 B.n467 B.n362 59.5399
R894 B.n185 B.n100 59.5399
R895 B.n98 B.n97 59.5399
R896 B.n485 B.n484 52.5581
R897 B.n362 B.n361 52.5581
R898 B.n100 B.n99 52.5581
R899 B.n97 B.n96 52.5581
R900 B.n577 B.n329 42.5852
R901 B.n583 B.n329 42.5852
R902 B.n583 B.n325 42.5852
R903 B.n589 B.n325 42.5852
R904 B.n589 B.n320 42.5852
R905 B.n595 B.n320 42.5852
R906 B.n595 B.n321 42.5852
R907 B.n601 B.n313 42.5852
R908 B.n607 B.n313 42.5852
R909 B.n607 B.n309 42.5852
R910 B.n613 B.n309 42.5852
R911 B.n613 B.n305 42.5852
R912 B.n619 B.n305 42.5852
R913 B.n619 B.n301 42.5852
R914 B.n625 B.n301 42.5852
R915 B.n625 B.n297 42.5852
R916 B.n631 B.n297 42.5852
R917 B.n638 B.n293 42.5852
R918 B.n638 B.n289 42.5852
R919 B.n644 B.n289 42.5852
R920 B.n644 B.n4 42.5852
R921 B.n730 B.n4 42.5852
R922 B.n730 B.n729 42.5852
R923 B.n729 B.n728 42.5852
R924 B.n728 B.n8 42.5852
R925 B.n722 B.n8 42.5852
R926 B.n722 B.n721 42.5852
R927 B.n720 B.n15 42.5852
R928 B.n714 B.n15 42.5852
R929 B.n714 B.n713 42.5852
R930 B.n713 B.n712 42.5852
R931 B.n712 B.n22 42.5852
R932 B.n706 B.n22 42.5852
R933 B.n706 B.n705 42.5852
R934 B.n705 B.n704 42.5852
R935 B.n704 B.n29 42.5852
R936 B.n698 B.n29 42.5852
R937 B.n697 B.n696 42.5852
R938 B.n696 B.n36 42.5852
R939 B.n690 B.n36 42.5852
R940 B.n690 B.n689 42.5852
R941 B.n689 B.n688 42.5852
R942 B.n688 B.n43 42.5852
R943 B.n682 B.n43 42.5852
R944 B.n601 B.t7 32.5653
R945 B.n698 B.t3 32.5653
R946 B.n679 B.n678 30.4395
R947 B.n684 B.n45 30.4395
R948 B.n575 B.n574 30.4395
R949 B.n579 B.n331 30.4395
R950 B.t1 B.n293 25.0503
R951 B.n721 B.t0 25.0503
R952 B B.n732 18.0485
R953 B.n631 B.t1 17.5354
R954 B.t0 B.n720 17.5354
R955 B.n101 B.n45 10.6151
R956 B.n104 B.n101 10.6151
R957 B.n105 B.n104 10.6151
R958 B.n108 B.n105 10.6151
R959 B.n109 B.n108 10.6151
R960 B.n112 B.n109 10.6151
R961 B.n113 B.n112 10.6151
R962 B.n116 B.n113 10.6151
R963 B.n117 B.n116 10.6151
R964 B.n120 B.n117 10.6151
R965 B.n121 B.n120 10.6151
R966 B.n124 B.n121 10.6151
R967 B.n125 B.n124 10.6151
R968 B.n128 B.n125 10.6151
R969 B.n129 B.n128 10.6151
R970 B.n132 B.n129 10.6151
R971 B.n133 B.n132 10.6151
R972 B.n136 B.n133 10.6151
R973 B.n137 B.n136 10.6151
R974 B.n140 B.n137 10.6151
R975 B.n141 B.n140 10.6151
R976 B.n144 B.n141 10.6151
R977 B.n145 B.n144 10.6151
R978 B.n148 B.n145 10.6151
R979 B.n149 B.n148 10.6151
R980 B.n152 B.n149 10.6151
R981 B.n153 B.n152 10.6151
R982 B.n156 B.n153 10.6151
R983 B.n157 B.n156 10.6151
R984 B.n160 B.n157 10.6151
R985 B.n161 B.n160 10.6151
R986 B.n164 B.n161 10.6151
R987 B.n165 B.n164 10.6151
R988 B.n168 B.n165 10.6151
R989 B.n169 B.n168 10.6151
R990 B.n172 B.n169 10.6151
R991 B.n173 B.n172 10.6151
R992 B.n176 B.n173 10.6151
R993 B.n177 B.n176 10.6151
R994 B.n180 B.n177 10.6151
R995 B.n181 B.n180 10.6151
R996 B.n184 B.n181 10.6151
R997 B.n189 B.n186 10.6151
R998 B.n190 B.n189 10.6151
R999 B.n193 B.n190 10.6151
R1000 B.n194 B.n193 10.6151
R1001 B.n197 B.n194 10.6151
R1002 B.n198 B.n197 10.6151
R1003 B.n201 B.n198 10.6151
R1004 B.n202 B.n201 10.6151
R1005 B.n206 B.n205 10.6151
R1006 B.n209 B.n206 10.6151
R1007 B.n210 B.n209 10.6151
R1008 B.n213 B.n210 10.6151
R1009 B.n214 B.n213 10.6151
R1010 B.n217 B.n214 10.6151
R1011 B.n218 B.n217 10.6151
R1012 B.n221 B.n218 10.6151
R1013 B.n222 B.n221 10.6151
R1014 B.n225 B.n222 10.6151
R1015 B.n226 B.n225 10.6151
R1016 B.n229 B.n226 10.6151
R1017 B.n230 B.n229 10.6151
R1018 B.n233 B.n230 10.6151
R1019 B.n234 B.n233 10.6151
R1020 B.n237 B.n234 10.6151
R1021 B.n238 B.n237 10.6151
R1022 B.n241 B.n238 10.6151
R1023 B.n242 B.n241 10.6151
R1024 B.n245 B.n242 10.6151
R1025 B.n246 B.n245 10.6151
R1026 B.n249 B.n246 10.6151
R1027 B.n250 B.n249 10.6151
R1028 B.n253 B.n250 10.6151
R1029 B.n254 B.n253 10.6151
R1030 B.n257 B.n254 10.6151
R1031 B.n258 B.n257 10.6151
R1032 B.n261 B.n258 10.6151
R1033 B.n262 B.n261 10.6151
R1034 B.n265 B.n262 10.6151
R1035 B.n266 B.n265 10.6151
R1036 B.n269 B.n266 10.6151
R1037 B.n270 B.n269 10.6151
R1038 B.n273 B.n270 10.6151
R1039 B.n274 B.n273 10.6151
R1040 B.n277 B.n274 10.6151
R1041 B.n278 B.n277 10.6151
R1042 B.n281 B.n278 10.6151
R1043 B.n282 B.n281 10.6151
R1044 B.n285 B.n282 10.6151
R1045 B.n286 B.n285 10.6151
R1046 B.n679 B.n286 10.6151
R1047 B.n575 B.n327 10.6151
R1048 B.n585 B.n327 10.6151
R1049 B.n586 B.n585 10.6151
R1050 B.n587 B.n586 10.6151
R1051 B.n587 B.n318 10.6151
R1052 B.n597 B.n318 10.6151
R1053 B.n598 B.n597 10.6151
R1054 B.n599 B.n598 10.6151
R1055 B.n599 B.n311 10.6151
R1056 B.n609 B.n311 10.6151
R1057 B.n610 B.n609 10.6151
R1058 B.n611 B.n610 10.6151
R1059 B.n611 B.n303 10.6151
R1060 B.n621 B.n303 10.6151
R1061 B.n622 B.n621 10.6151
R1062 B.n623 B.n622 10.6151
R1063 B.n623 B.n295 10.6151
R1064 B.n633 B.n295 10.6151
R1065 B.n634 B.n633 10.6151
R1066 B.n636 B.n634 10.6151
R1067 B.n636 B.n635 10.6151
R1068 B.n635 B.n287 10.6151
R1069 B.n647 B.n287 10.6151
R1070 B.n648 B.n647 10.6151
R1071 B.n649 B.n648 10.6151
R1072 B.n650 B.n649 10.6151
R1073 B.n652 B.n650 10.6151
R1074 B.n653 B.n652 10.6151
R1075 B.n654 B.n653 10.6151
R1076 B.n655 B.n654 10.6151
R1077 B.n657 B.n655 10.6151
R1078 B.n658 B.n657 10.6151
R1079 B.n659 B.n658 10.6151
R1080 B.n660 B.n659 10.6151
R1081 B.n662 B.n660 10.6151
R1082 B.n663 B.n662 10.6151
R1083 B.n664 B.n663 10.6151
R1084 B.n665 B.n664 10.6151
R1085 B.n667 B.n665 10.6151
R1086 B.n668 B.n667 10.6151
R1087 B.n669 B.n668 10.6151
R1088 B.n670 B.n669 10.6151
R1089 B.n672 B.n670 10.6151
R1090 B.n673 B.n672 10.6151
R1091 B.n674 B.n673 10.6151
R1092 B.n675 B.n674 10.6151
R1093 B.n677 B.n675 10.6151
R1094 B.n678 B.n677 10.6151
R1095 B.n385 B.n331 10.6151
R1096 B.n386 B.n385 10.6151
R1097 B.n387 B.n386 10.6151
R1098 B.n387 B.n381 10.6151
R1099 B.n393 B.n381 10.6151
R1100 B.n394 B.n393 10.6151
R1101 B.n395 B.n394 10.6151
R1102 B.n395 B.n379 10.6151
R1103 B.n401 B.n379 10.6151
R1104 B.n402 B.n401 10.6151
R1105 B.n403 B.n402 10.6151
R1106 B.n403 B.n377 10.6151
R1107 B.n409 B.n377 10.6151
R1108 B.n410 B.n409 10.6151
R1109 B.n411 B.n410 10.6151
R1110 B.n411 B.n375 10.6151
R1111 B.n417 B.n375 10.6151
R1112 B.n418 B.n417 10.6151
R1113 B.n419 B.n418 10.6151
R1114 B.n419 B.n373 10.6151
R1115 B.n425 B.n373 10.6151
R1116 B.n426 B.n425 10.6151
R1117 B.n427 B.n426 10.6151
R1118 B.n427 B.n371 10.6151
R1119 B.n433 B.n371 10.6151
R1120 B.n434 B.n433 10.6151
R1121 B.n435 B.n434 10.6151
R1122 B.n435 B.n369 10.6151
R1123 B.n441 B.n369 10.6151
R1124 B.n442 B.n441 10.6151
R1125 B.n443 B.n442 10.6151
R1126 B.n443 B.n367 10.6151
R1127 B.n449 B.n367 10.6151
R1128 B.n450 B.n449 10.6151
R1129 B.n451 B.n450 10.6151
R1130 B.n451 B.n365 10.6151
R1131 B.n457 B.n365 10.6151
R1132 B.n458 B.n457 10.6151
R1133 B.n459 B.n458 10.6151
R1134 B.n459 B.n363 10.6151
R1135 B.n465 B.n363 10.6151
R1136 B.n466 B.n465 10.6151
R1137 B.n468 B.n359 10.6151
R1138 B.n474 B.n359 10.6151
R1139 B.n475 B.n474 10.6151
R1140 B.n476 B.n475 10.6151
R1141 B.n476 B.n357 10.6151
R1142 B.n482 B.n357 10.6151
R1143 B.n483 B.n482 10.6151
R1144 B.n487 B.n483 10.6151
R1145 B.n493 B.n355 10.6151
R1146 B.n494 B.n493 10.6151
R1147 B.n495 B.n494 10.6151
R1148 B.n495 B.n353 10.6151
R1149 B.n501 B.n353 10.6151
R1150 B.n502 B.n501 10.6151
R1151 B.n503 B.n502 10.6151
R1152 B.n503 B.n351 10.6151
R1153 B.n509 B.n351 10.6151
R1154 B.n510 B.n509 10.6151
R1155 B.n511 B.n510 10.6151
R1156 B.n511 B.n349 10.6151
R1157 B.n517 B.n349 10.6151
R1158 B.n518 B.n517 10.6151
R1159 B.n519 B.n518 10.6151
R1160 B.n519 B.n347 10.6151
R1161 B.n525 B.n347 10.6151
R1162 B.n526 B.n525 10.6151
R1163 B.n527 B.n526 10.6151
R1164 B.n527 B.n345 10.6151
R1165 B.n533 B.n345 10.6151
R1166 B.n534 B.n533 10.6151
R1167 B.n535 B.n534 10.6151
R1168 B.n535 B.n343 10.6151
R1169 B.n541 B.n343 10.6151
R1170 B.n542 B.n541 10.6151
R1171 B.n543 B.n542 10.6151
R1172 B.n543 B.n341 10.6151
R1173 B.n549 B.n341 10.6151
R1174 B.n550 B.n549 10.6151
R1175 B.n551 B.n550 10.6151
R1176 B.n551 B.n339 10.6151
R1177 B.n557 B.n339 10.6151
R1178 B.n558 B.n557 10.6151
R1179 B.n559 B.n558 10.6151
R1180 B.n559 B.n337 10.6151
R1181 B.n565 B.n337 10.6151
R1182 B.n566 B.n565 10.6151
R1183 B.n567 B.n566 10.6151
R1184 B.n567 B.n335 10.6151
R1185 B.n573 B.n335 10.6151
R1186 B.n574 B.n573 10.6151
R1187 B.n580 B.n579 10.6151
R1188 B.n581 B.n580 10.6151
R1189 B.n581 B.n323 10.6151
R1190 B.n591 B.n323 10.6151
R1191 B.n592 B.n591 10.6151
R1192 B.n593 B.n592 10.6151
R1193 B.n593 B.n315 10.6151
R1194 B.n603 B.n315 10.6151
R1195 B.n604 B.n603 10.6151
R1196 B.n605 B.n604 10.6151
R1197 B.n605 B.n307 10.6151
R1198 B.n615 B.n307 10.6151
R1199 B.n616 B.n615 10.6151
R1200 B.n617 B.n616 10.6151
R1201 B.n617 B.n299 10.6151
R1202 B.n627 B.n299 10.6151
R1203 B.n628 B.n627 10.6151
R1204 B.n629 B.n628 10.6151
R1205 B.n629 B.n291 10.6151
R1206 B.n640 B.n291 10.6151
R1207 B.n641 B.n640 10.6151
R1208 B.n642 B.n641 10.6151
R1209 B.n642 B.n0 10.6151
R1210 B.n726 B.n1 10.6151
R1211 B.n726 B.n725 10.6151
R1212 B.n725 B.n724 10.6151
R1213 B.n724 B.n10 10.6151
R1214 B.n718 B.n10 10.6151
R1215 B.n718 B.n717 10.6151
R1216 B.n717 B.n716 10.6151
R1217 B.n716 B.n17 10.6151
R1218 B.n710 B.n17 10.6151
R1219 B.n710 B.n709 10.6151
R1220 B.n709 B.n708 10.6151
R1221 B.n708 B.n24 10.6151
R1222 B.n702 B.n24 10.6151
R1223 B.n702 B.n701 10.6151
R1224 B.n701 B.n700 10.6151
R1225 B.n700 B.n31 10.6151
R1226 B.n694 B.n31 10.6151
R1227 B.n694 B.n693 10.6151
R1228 B.n693 B.n692 10.6151
R1229 B.n692 B.n38 10.6151
R1230 B.n686 B.n38 10.6151
R1231 B.n686 B.n685 10.6151
R1232 B.n685 B.n684 10.6151
R1233 B.n321 B.t7 10.0204
R1234 B.t3 B.n697 10.0204
R1235 B.n186 B.n185 6.5566
R1236 B.n202 B.n98 6.5566
R1237 B.n468 B.n467 6.5566
R1238 B.n487 B.n486 6.5566
R1239 B.n185 B.n184 4.05904
R1240 B.n205 B.n98 4.05904
R1241 B.n467 B.n466 4.05904
R1242 B.n486 B.n355 4.05904
R1243 B.n732 B.n0 2.81026
R1244 B.n732 B.n1 2.81026
R1245 VN VN.t0 218.01
R1246 VN VN.t1 173.957
R1247 VDD2.n0 VDD2.t0 105.078
R1248 VDD2.n0 VDD2.t1 66.1506
R1249 VDD2 VDD2.n0 0.642741
C0 VTAIL VDD1 5.11782f
C1 VP VDD2 0.32386f
C2 VN VDD2 2.80134f
C3 VP VTAIL 2.44848f
C4 VN VTAIL 2.43417f
C5 VP VDD1 2.97447f
C6 VDD2 VTAIL 5.16664f
C7 VN VDD1 0.148021f
C8 VDD2 VDD1 0.648332f
C9 VP VN 5.40619f
C10 VDD2 B 4.406115f
C11 VDD1 B 7.50216f
C12 VTAIL B 7.39113f
C13 VN B 10.528509f
C14 VP B 6.14569f
C15 VDD2.t0 B 2.77701f
C16 VDD2.t1 B 2.25223f
C17 VDD2.n0 B 2.85184f
C18 VN.t1 B 2.88913f
C19 VN.t0 B 3.37364f
C20 VDD1.t0 B 2.26175f
C21 VDD1.t1 B 2.82006f
C22 VTAIL.t3 B 2.20215f
C23 VTAIL.n0 B 1.61522f
C24 VTAIL.t1 B 2.20214f
C25 VTAIL.n1 B 1.64992f
C26 VTAIL.t2 B 2.20214f
C27 VTAIL.n2 B 1.4958f
C28 VTAIL.t0 B 2.20215f
C29 VTAIL.n3 B 1.42242f
C30 VP.t1 B 3.44882f
C31 VP.t0 B 2.95446f
C32 VP.n0 B 4.32435f
.ends

