* NGSPICE file created from diff_pair_sample_0619.ext - technology: sky130A

.subckt diff_pair_sample_0619 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X1 VTAIL.t5 VN.t0 VDD2.t9 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X2 VDD1.t8 VP.t1 VTAIL.t17 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.54
X3 VTAIL.t10 VP.t2 VDD1.t7 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X4 B.t11 B.t9 B.t10 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.54
X5 VTAIL.t19 VP.t3 VDD1.t6 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X6 VTAIL.t12 VP.t4 VDD1.t5 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X7 VTAIL.t7 VN.t1 VDD2.t8 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X8 VDD2.t7 VN.t2 VTAIL.t1 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.54
X9 VDD2.t6 VN.t3 VTAIL.t4 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.54
X10 VDD2.t5 VN.t4 VTAIL.t6 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X11 B.t8 B.t6 B.t7 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.54
X12 VDD2.t4 VN.t5 VTAIL.t0 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.54
X13 VDD1.t4 VP.t5 VTAIL.t13 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.54
X14 VTAIL.t2 VN.t6 VDD2.t3 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X15 VDD2.t2 VN.t7 VTAIL.t9 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X16 VDD2.t1 VN.t8 VTAIL.t8 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.54
X17 B.t5 B.t3 B.t4 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.54
X18 VTAIL.t3 VN.t9 VDD2.t0 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X19 VTAIL.t14 VP.t6 VDD1.t3 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X20 VDD1.t2 VP.t7 VTAIL.t11 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.54
X21 VDD1.t1 VP.t8 VTAIL.t15 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.54
X22 B.t2 B.t0 B.t1 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.54
X23 VDD1.t0 VP.t9 VTAIL.t16 w_n3214_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.54
R0 VP.n15 VP.t8 208.109
R1 VP.n36 VP.n35 174.089
R2 VP.n62 VP.n61 174.089
R3 VP.n34 VP.n33 174.089
R4 VP.n48 VP.t7 173.395
R5 VP.n35 VP.t9 173.395
R6 VP.n41 VP.t6 173.395
R7 VP.n54 VP.t3 173.395
R8 VP.n61 VP.t1 173.395
R9 VP.n20 VP.t0 173.395
R10 VP.n33 VP.t5 173.395
R11 VP.n26 VP.t4 173.395
R12 VP.n14 VP.t2 173.395
R13 VP.n16 VP.n13 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n12 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n11 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n25 VP.n10 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n29 VP.n9 161.3
R22 VP.n31 VP.n30 161.3
R23 VP.n32 VP.n8 161.3
R24 VP.n60 VP.n0 161.3
R25 VP.n59 VP.n58 161.3
R26 VP.n57 VP.n1 161.3
R27 VP.n56 VP.n55 161.3
R28 VP.n53 VP.n2 161.3
R29 VP.n52 VP.n51 161.3
R30 VP.n50 VP.n3 161.3
R31 VP.n49 VP.n48 161.3
R32 VP.n47 VP.n4 161.3
R33 VP.n46 VP.n45 161.3
R34 VP.n44 VP.n5 161.3
R35 VP.n43 VP.n42 161.3
R36 VP.n40 VP.n6 161.3
R37 VP.n39 VP.n38 161.3
R38 VP.n37 VP.n7 161.3
R39 VP.n40 VP.n39 56.5617
R40 VP.n59 VP.n1 56.5617
R41 VP.n31 VP.n9 56.5617
R42 VP.n15 VP.n14 48.5587
R43 VP.n47 VP.n46 46.874
R44 VP.n52 VP.n3 46.874
R45 VP.n24 VP.n11 46.874
R46 VP.n19 VP.n18 46.874
R47 VP.n36 VP.n34 46.6179
R48 VP.n46 VP.n5 34.28
R49 VP.n53 VP.n52 34.28
R50 VP.n25 VP.n24 34.28
R51 VP.n18 VP.n13 34.28
R52 VP.n39 VP.n7 24.5923
R53 VP.n42 VP.n40 24.5923
R54 VP.n48 VP.n47 24.5923
R55 VP.n48 VP.n3 24.5923
R56 VP.n55 VP.n1 24.5923
R57 VP.n60 VP.n59 24.5923
R58 VP.n32 VP.n31 24.5923
R59 VP.n27 VP.n9 24.5923
R60 VP.n20 VP.n19 24.5923
R61 VP.n20 VP.n11 24.5923
R62 VP.n41 VP.n5 18.1985
R63 VP.n54 VP.n53 18.1985
R64 VP.n26 VP.n25 18.1985
R65 VP.n14 VP.n13 18.1985
R66 VP.n16 VP.n15 17.587
R67 VP.n35 VP.n7 11.8046
R68 VP.n61 VP.n60 11.8046
R69 VP.n33 VP.n32 11.8046
R70 VP.n42 VP.n41 6.39438
R71 VP.n55 VP.n54 6.39438
R72 VP.n27 VP.n26 6.39438
R73 VP.n17 VP.n16 0.189894
R74 VP.n17 VP.n12 0.189894
R75 VP.n21 VP.n12 0.189894
R76 VP.n22 VP.n21 0.189894
R77 VP.n23 VP.n22 0.189894
R78 VP.n23 VP.n10 0.189894
R79 VP.n28 VP.n10 0.189894
R80 VP.n29 VP.n28 0.189894
R81 VP.n30 VP.n29 0.189894
R82 VP.n30 VP.n8 0.189894
R83 VP.n34 VP.n8 0.189894
R84 VP.n37 VP.n36 0.189894
R85 VP.n38 VP.n37 0.189894
R86 VP.n38 VP.n6 0.189894
R87 VP.n43 VP.n6 0.189894
R88 VP.n44 VP.n43 0.189894
R89 VP.n45 VP.n44 0.189894
R90 VP.n45 VP.n4 0.189894
R91 VP.n49 VP.n4 0.189894
R92 VP.n50 VP.n49 0.189894
R93 VP.n51 VP.n50 0.189894
R94 VP.n51 VP.n2 0.189894
R95 VP.n56 VP.n2 0.189894
R96 VP.n57 VP.n56 0.189894
R97 VP.n58 VP.n57 0.189894
R98 VP.n58 VP.n0 0.189894
R99 VP.n62 VP.n0 0.189894
R100 VP VP.n62 0.0516364
R101 VTAIL.n11 VTAIL.t4 62.3356
R102 VTAIL.n17 VTAIL.t0 62.3355
R103 VTAIL.n2 VTAIL.t17 62.3355
R104 VTAIL.n16 VTAIL.t13 62.3355
R105 VTAIL.n15 VTAIL.n14 59.402
R106 VTAIL.n13 VTAIL.n12 59.402
R107 VTAIL.n10 VTAIL.n9 59.402
R108 VTAIL.n8 VTAIL.n7 59.402
R109 VTAIL.n19 VTAIL.n18 59.4018
R110 VTAIL.n1 VTAIL.n0 59.4018
R111 VTAIL.n4 VTAIL.n3 59.4018
R112 VTAIL.n6 VTAIL.n5 59.4018
R113 VTAIL.n8 VTAIL.n6 25.1427
R114 VTAIL.n17 VTAIL.n16 23.5307
R115 VTAIL.n18 VTAIL.t6 2.93416
R116 VTAIL.n18 VTAIL.t7 2.93416
R117 VTAIL.n0 VTAIL.t8 2.93416
R118 VTAIL.n0 VTAIL.t2 2.93416
R119 VTAIL.n3 VTAIL.t11 2.93416
R120 VTAIL.n3 VTAIL.t19 2.93416
R121 VTAIL.n5 VTAIL.t16 2.93416
R122 VTAIL.n5 VTAIL.t14 2.93416
R123 VTAIL.n14 VTAIL.t18 2.93416
R124 VTAIL.n14 VTAIL.t12 2.93416
R125 VTAIL.n12 VTAIL.t15 2.93416
R126 VTAIL.n12 VTAIL.t10 2.93416
R127 VTAIL.n9 VTAIL.t9 2.93416
R128 VTAIL.n9 VTAIL.t3 2.93416
R129 VTAIL.n7 VTAIL.t1 2.93416
R130 VTAIL.n7 VTAIL.t5 2.93416
R131 VTAIL.n10 VTAIL.n8 1.61257
R132 VTAIL.n11 VTAIL.n10 1.61257
R133 VTAIL.n15 VTAIL.n13 1.61257
R134 VTAIL.n16 VTAIL.n15 1.61257
R135 VTAIL.n6 VTAIL.n4 1.61257
R136 VTAIL.n4 VTAIL.n2 1.61257
R137 VTAIL.n19 VTAIL.n17 1.61257
R138 VTAIL.n13 VTAIL.n11 1.27636
R139 VTAIL.n2 VTAIL.n1 1.27636
R140 VTAIL VTAIL.n1 1.26774
R141 VTAIL VTAIL.n19 0.345328
R142 VDD1.n1 VDD1.t1 80.6265
R143 VDD1.n3 VDD1.t0 80.6264
R144 VDD1.n5 VDD1.n4 77.2343
R145 VDD1.n1 VDD1.n0 76.0808
R146 VDD1.n7 VDD1.n6 76.0806
R147 VDD1.n3 VDD1.n2 76.0806
R148 VDD1.n7 VDD1.n5 42.3134
R149 VDD1.n6 VDD1.t5 2.93416
R150 VDD1.n6 VDD1.t4 2.93416
R151 VDD1.n0 VDD1.t7 2.93416
R152 VDD1.n0 VDD1.t9 2.93416
R153 VDD1.n4 VDD1.t6 2.93416
R154 VDD1.n4 VDD1.t8 2.93416
R155 VDD1.n2 VDD1.t3 2.93416
R156 VDD1.n2 VDD1.t2 2.93416
R157 VDD1 VDD1.n7 1.15136
R158 VDD1 VDD1.n1 0.461707
R159 VDD1.n5 VDD1.n3 0.348171
R160 VN.n7 VN.t8 208.109
R161 VN.n34 VN.t3 208.109
R162 VN.n26 VN.n25 174.089
R163 VN.n53 VN.n52 174.089
R164 VN.n12 VN.t4 173.395
R165 VN.n6 VN.t6 173.395
R166 VN.n18 VN.t1 173.395
R167 VN.n25 VN.t5 173.395
R168 VN.n39 VN.t7 173.395
R169 VN.n33 VN.t9 173.395
R170 VN.n45 VN.t0 173.395
R171 VN.n52 VN.t2 173.395
R172 VN.n51 VN.n27 161.3
R173 VN.n50 VN.n49 161.3
R174 VN.n48 VN.n28 161.3
R175 VN.n47 VN.n46 161.3
R176 VN.n44 VN.n29 161.3
R177 VN.n43 VN.n42 161.3
R178 VN.n41 VN.n30 161.3
R179 VN.n40 VN.n39 161.3
R180 VN.n38 VN.n31 161.3
R181 VN.n37 VN.n36 161.3
R182 VN.n35 VN.n32 161.3
R183 VN.n24 VN.n0 161.3
R184 VN.n23 VN.n22 161.3
R185 VN.n21 VN.n1 161.3
R186 VN.n20 VN.n19 161.3
R187 VN.n17 VN.n2 161.3
R188 VN.n16 VN.n15 161.3
R189 VN.n14 VN.n3 161.3
R190 VN.n13 VN.n12 161.3
R191 VN.n11 VN.n4 161.3
R192 VN.n10 VN.n9 161.3
R193 VN.n8 VN.n5 161.3
R194 VN.n23 VN.n1 56.5617
R195 VN.n50 VN.n28 56.5617
R196 VN.n7 VN.n6 48.5587
R197 VN.n34 VN.n33 48.5587
R198 VN VN.n53 46.9986
R199 VN.n11 VN.n10 46.874
R200 VN.n16 VN.n3 46.874
R201 VN.n38 VN.n37 46.874
R202 VN.n43 VN.n30 46.874
R203 VN.n10 VN.n5 34.28
R204 VN.n17 VN.n16 34.28
R205 VN.n37 VN.n32 34.28
R206 VN.n44 VN.n43 34.28
R207 VN.n12 VN.n11 24.5923
R208 VN.n12 VN.n3 24.5923
R209 VN.n19 VN.n1 24.5923
R210 VN.n24 VN.n23 24.5923
R211 VN.n39 VN.n30 24.5923
R212 VN.n39 VN.n38 24.5923
R213 VN.n46 VN.n28 24.5923
R214 VN.n51 VN.n50 24.5923
R215 VN.n6 VN.n5 18.1985
R216 VN.n18 VN.n17 18.1985
R217 VN.n33 VN.n32 18.1985
R218 VN.n45 VN.n44 18.1985
R219 VN.n35 VN.n34 17.587
R220 VN.n8 VN.n7 17.587
R221 VN.n25 VN.n24 11.8046
R222 VN.n52 VN.n51 11.8046
R223 VN.n19 VN.n18 6.39438
R224 VN.n46 VN.n45 6.39438
R225 VN.n53 VN.n27 0.189894
R226 VN.n49 VN.n27 0.189894
R227 VN.n49 VN.n48 0.189894
R228 VN.n48 VN.n47 0.189894
R229 VN.n47 VN.n29 0.189894
R230 VN.n42 VN.n29 0.189894
R231 VN.n42 VN.n41 0.189894
R232 VN.n41 VN.n40 0.189894
R233 VN.n40 VN.n31 0.189894
R234 VN.n36 VN.n31 0.189894
R235 VN.n36 VN.n35 0.189894
R236 VN.n9 VN.n8 0.189894
R237 VN.n9 VN.n4 0.189894
R238 VN.n13 VN.n4 0.189894
R239 VN.n14 VN.n13 0.189894
R240 VN.n15 VN.n14 0.189894
R241 VN.n15 VN.n2 0.189894
R242 VN.n20 VN.n2 0.189894
R243 VN.n21 VN.n20 0.189894
R244 VN.n22 VN.n21 0.189894
R245 VN.n22 VN.n0 0.189894
R246 VN.n26 VN.n0 0.189894
R247 VN VN.n26 0.0516364
R248 VDD2.n1 VDD2.t1 80.6264
R249 VDD2.n4 VDD2.t7 79.0144
R250 VDD2.n3 VDD2.n2 77.2343
R251 VDD2 VDD2.n7 77.2315
R252 VDD2.n6 VDD2.n5 76.0808
R253 VDD2.n1 VDD2.n0 76.0806
R254 VDD2.n4 VDD2.n3 40.9243
R255 VDD2.n7 VDD2.t0 2.93416
R256 VDD2.n7 VDD2.t6 2.93416
R257 VDD2.n5 VDD2.t9 2.93416
R258 VDD2.n5 VDD2.t2 2.93416
R259 VDD2.n2 VDD2.t8 2.93416
R260 VDD2.n2 VDD2.t4 2.93416
R261 VDD2.n0 VDD2.t3 2.93416
R262 VDD2.n0 VDD2.t5 2.93416
R263 VDD2.n6 VDD2.n4 1.61257
R264 VDD2 VDD2.n6 0.461707
R265 VDD2.n3 VDD2.n1 0.348171
R266 B.n497 B.n70 585
R267 B.n499 B.n498 585
R268 B.n500 B.n69 585
R269 B.n502 B.n501 585
R270 B.n503 B.n68 585
R271 B.n505 B.n504 585
R272 B.n506 B.n67 585
R273 B.n508 B.n507 585
R274 B.n509 B.n66 585
R275 B.n511 B.n510 585
R276 B.n512 B.n65 585
R277 B.n514 B.n513 585
R278 B.n515 B.n64 585
R279 B.n517 B.n516 585
R280 B.n518 B.n63 585
R281 B.n520 B.n519 585
R282 B.n521 B.n62 585
R283 B.n523 B.n522 585
R284 B.n524 B.n61 585
R285 B.n526 B.n525 585
R286 B.n527 B.n60 585
R287 B.n529 B.n528 585
R288 B.n530 B.n59 585
R289 B.n532 B.n531 585
R290 B.n533 B.n58 585
R291 B.n535 B.n534 585
R292 B.n536 B.n57 585
R293 B.n538 B.n537 585
R294 B.n539 B.n56 585
R295 B.n541 B.n540 585
R296 B.n542 B.n55 585
R297 B.n544 B.n543 585
R298 B.n545 B.n54 585
R299 B.n547 B.n546 585
R300 B.n548 B.n53 585
R301 B.n550 B.n549 585
R302 B.n551 B.n52 585
R303 B.n553 B.n552 585
R304 B.n554 B.n49 585
R305 B.n557 B.n556 585
R306 B.n558 B.n48 585
R307 B.n560 B.n559 585
R308 B.n561 B.n47 585
R309 B.n563 B.n562 585
R310 B.n564 B.n46 585
R311 B.n566 B.n565 585
R312 B.n567 B.n45 585
R313 B.n569 B.n568 585
R314 B.n571 B.n570 585
R315 B.n572 B.n41 585
R316 B.n574 B.n573 585
R317 B.n575 B.n40 585
R318 B.n577 B.n576 585
R319 B.n578 B.n39 585
R320 B.n580 B.n579 585
R321 B.n581 B.n38 585
R322 B.n583 B.n582 585
R323 B.n584 B.n37 585
R324 B.n586 B.n585 585
R325 B.n587 B.n36 585
R326 B.n589 B.n588 585
R327 B.n590 B.n35 585
R328 B.n592 B.n591 585
R329 B.n593 B.n34 585
R330 B.n595 B.n594 585
R331 B.n596 B.n33 585
R332 B.n598 B.n597 585
R333 B.n599 B.n32 585
R334 B.n601 B.n600 585
R335 B.n602 B.n31 585
R336 B.n604 B.n603 585
R337 B.n605 B.n30 585
R338 B.n607 B.n606 585
R339 B.n608 B.n29 585
R340 B.n610 B.n609 585
R341 B.n611 B.n28 585
R342 B.n613 B.n612 585
R343 B.n614 B.n27 585
R344 B.n616 B.n615 585
R345 B.n617 B.n26 585
R346 B.n619 B.n618 585
R347 B.n620 B.n25 585
R348 B.n622 B.n621 585
R349 B.n623 B.n24 585
R350 B.n625 B.n624 585
R351 B.n626 B.n23 585
R352 B.n628 B.n627 585
R353 B.n496 B.n495 585
R354 B.n494 B.n71 585
R355 B.n493 B.n492 585
R356 B.n491 B.n72 585
R357 B.n490 B.n489 585
R358 B.n488 B.n73 585
R359 B.n487 B.n486 585
R360 B.n485 B.n74 585
R361 B.n484 B.n483 585
R362 B.n482 B.n75 585
R363 B.n481 B.n480 585
R364 B.n479 B.n76 585
R365 B.n478 B.n477 585
R366 B.n476 B.n77 585
R367 B.n475 B.n474 585
R368 B.n473 B.n78 585
R369 B.n472 B.n471 585
R370 B.n470 B.n79 585
R371 B.n469 B.n468 585
R372 B.n467 B.n80 585
R373 B.n466 B.n465 585
R374 B.n464 B.n81 585
R375 B.n463 B.n462 585
R376 B.n461 B.n82 585
R377 B.n460 B.n459 585
R378 B.n458 B.n83 585
R379 B.n457 B.n456 585
R380 B.n455 B.n84 585
R381 B.n454 B.n453 585
R382 B.n452 B.n85 585
R383 B.n451 B.n450 585
R384 B.n449 B.n86 585
R385 B.n448 B.n447 585
R386 B.n446 B.n87 585
R387 B.n445 B.n444 585
R388 B.n443 B.n88 585
R389 B.n442 B.n441 585
R390 B.n440 B.n89 585
R391 B.n439 B.n438 585
R392 B.n437 B.n90 585
R393 B.n436 B.n435 585
R394 B.n434 B.n91 585
R395 B.n433 B.n432 585
R396 B.n431 B.n92 585
R397 B.n430 B.n429 585
R398 B.n428 B.n93 585
R399 B.n427 B.n426 585
R400 B.n425 B.n94 585
R401 B.n424 B.n423 585
R402 B.n422 B.n95 585
R403 B.n421 B.n420 585
R404 B.n419 B.n96 585
R405 B.n418 B.n417 585
R406 B.n416 B.n97 585
R407 B.n415 B.n414 585
R408 B.n413 B.n98 585
R409 B.n412 B.n411 585
R410 B.n410 B.n99 585
R411 B.n409 B.n408 585
R412 B.n407 B.n100 585
R413 B.n406 B.n405 585
R414 B.n404 B.n101 585
R415 B.n403 B.n402 585
R416 B.n401 B.n102 585
R417 B.n400 B.n399 585
R418 B.n398 B.n103 585
R419 B.n397 B.n396 585
R420 B.n395 B.n104 585
R421 B.n394 B.n393 585
R422 B.n392 B.n105 585
R423 B.n391 B.n390 585
R424 B.n389 B.n106 585
R425 B.n388 B.n387 585
R426 B.n386 B.n107 585
R427 B.n385 B.n384 585
R428 B.n383 B.n108 585
R429 B.n382 B.n381 585
R430 B.n380 B.n109 585
R431 B.n379 B.n378 585
R432 B.n377 B.n110 585
R433 B.n376 B.n375 585
R434 B.n374 B.n111 585
R435 B.n373 B.n372 585
R436 B.n241 B.n240 585
R437 B.n242 B.n159 585
R438 B.n244 B.n243 585
R439 B.n245 B.n158 585
R440 B.n247 B.n246 585
R441 B.n248 B.n157 585
R442 B.n250 B.n249 585
R443 B.n251 B.n156 585
R444 B.n253 B.n252 585
R445 B.n254 B.n155 585
R446 B.n256 B.n255 585
R447 B.n257 B.n154 585
R448 B.n259 B.n258 585
R449 B.n260 B.n153 585
R450 B.n262 B.n261 585
R451 B.n263 B.n152 585
R452 B.n265 B.n264 585
R453 B.n266 B.n151 585
R454 B.n268 B.n267 585
R455 B.n269 B.n150 585
R456 B.n271 B.n270 585
R457 B.n272 B.n149 585
R458 B.n274 B.n273 585
R459 B.n275 B.n148 585
R460 B.n277 B.n276 585
R461 B.n278 B.n147 585
R462 B.n280 B.n279 585
R463 B.n281 B.n146 585
R464 B.n283 B.n282 585
R465 B.n284 B.n145 585
R466 B.n286 B.n285 585
R467 B.n287 B.n144 585
R468 B.n289 B.n288 585
R469 B.n290 B.n143 585
R470 B.n292 B.n291 585
R471 B.n293 B.n142 585
R472 B.n295 B.n294 585
R473 B.n296 B.n141 585
R474 B.n298 B.n297 585
R475 B.n300 B.n299 585
R476 B.n301 B.n137 585
R477 B.n303 B.n302 585
R478 B.n304 B.n136 585
R479 B.n306 B.n305 585
R480 B.n307 B.n135 585
R481 B.n309 B.n308 585
R482 B.n310 B.n134 585
R483 B.n312 B.n311 585
R484 B.n314 B.n131 585
R485 B.n316 B.n315 585
R486 B.n317 B.n130 585
R487 B.n319 B.n318 585
R488 B.n320 B.n129 585
R489 B.n322 B.n321 585
R490 B.n323 B.n128 585
R491 B.n325 B.n324 585
R492 B.n326 B.n127 585
R493 B.n328 B.n327 585
R494 B.n329 B.n126 585
R495 B.n331 B.n330 585
R496 B.n332 B.n125 585
R497 B.n334 B.n333 585
R498 B.n335 B.n124 585
R499 B.n337 B.n336 585
R500 B.n338 B.n123 585
R501 B.n340 B.n339 585
R502 B.n341 B.n122 585
R503 B.n343 B.n342 585
R504 B.n344 B.n121 585
R505 B.n346 B.n345 585
R506 B.n347 B.n120 585
R507 B.n349 B.n348 585
R508 B.n350 B.n119 585
R509 B.n352 B.n351 585
R510 B.n353 B.n118 585
R511 B.n355 B.n354 585
R512 B.n356 B.n117 585
R513 B.n358 B.n357 585
R514 B.n359 B.n116 585
R515 B.n361 B.n360 585
R516 B.n362 B.n115 585
R517 B.n364 B.n363 585
R518 B.n365 B.n114 585
R519 B.n367 B.n366 585
R520 B.n368 B.n113 585
R521 B.n370 B.n369 585
R522 B.n371 B.n112 585
R523 B.n239 B.n160 585
R524 B.n238 B.n237 585
R525 B.n236 B.n161 585
R526 B.n235 B.n234 585
R527 B.n233 B.n162 585
R528 B.n232 B.n231 585
R529 B.n230 B.n163 585
R530 B.n229 B.n228 585
R531 B.n227 B.n164 585
R532 B.n226 B.n225 585
R533 B.n224 B.n165 585
R534 B.n223 B.n222 585
R535 B.n221 B.n166 585
R536 B.n220 B.n219 585
R537 B.n218 B.n167 585
R538 B.n217 B.n216 585
R539 B.n215 B.n168 585
R540 B.n214 B.n213 585
R541 B.n212 B.n169 585
R542 B.n211 B.n210 585
R543 B.n209 B.n170 585
R544 B.n208 B.n207 585
R545 B.n206 B.n171 585
R546 B.n205 B.n204 585
R547 B.n203 B.n172 585
R548 B.n202 B.n201 585
R549 B.n200 B.n173 585
R550 B.n199 B.n198 585
R551 B.n197 B.n174 585
R552 B.n196 B.n195 585
R553 B.n194 B.n175 585
R554 B.n193 B.n192 585
R555 B.n191 B.n176 585
R556 B.n190 B.n189 585
R557 B.n188 B.n177 585
R558 B.n187 B.n186 585
R559 B.n185 B.n178 585
R560 B.n184 B.n183 585
R561 B.n182 B.n179 585
R562 B.n181 B.n180 585
R563 B.n2 B.n0 585
R564 B.n689 B.n1 585
R565 B.n688 B.n687 585
R566 B.n686 B.n3 585
R567 B.n685 B.n684 585
R568 B.n683 B.n4 585
R569 B.n682 B.n681 585
R570 B.n680 B.n5 585
R571 B.n679 B.n678 585
R572 B.n677 B.n6 585
R573 B.n676 B.n675 585
R574 B.n674 B.n7 585
R575 B.n673 B.n672 585
R576 B.n671 B.n8 585
R577 B.n670 B.n669 585
R578 B.n668 B.n9 585
R579 B.n667 B.n666 585
R580 B.n665 B.n10 585
R581 B.n664 B.n663 585
R582 B.n662 B.n11 585
R583 B.n661 B.n660 585
R584 B.n659 B.n12 585
R585 B.n658 B.n657 585
R586 B.n656 B.n13 585
R587 B.n655 B.n654 585
R588 B.n653 B.n14 585
R589 B.n652 B.n651 585
R590 B.n650 B.n15 585
R591 B.n649 B.n648 585
R592 B.n647 B.n16 585
R593 B.n646 B.n645 585
R594 B.n644 B.n17 585
R595 B.n643 B.n642 585
R596 B.n641 B.n18 585
R597 B.n640 B.n639 585
R598 B.n638 B.n19 585
R599 B.n637 B.n636 585
R600 B.n635 B.n20 585
R601 B.n634 B.n633 585
R602 B.n632 B.n21 585
R603 B.n631 B.n630 585
R604 B.n629 B.n22 585
R605 B.n691 B.n690 585
R606 B.n240 B.n239 550.159
R607 B.n629 B.n628 550.159
R608 B.n372 B.n371 550.159
R609 B.n497 B.n496 550.159
R610 B.n132 B.t3 378.981
R611 B.n138 B.t0 378.981
R612 B.n42 B.t9 378.981
R613 B.n50 B.t6 378.981
R614 B.n239 B.n238 163.367
R615 B.n238 B.n161 163.367
R616 B.n234 B.n161 163.367
R617 B.n234 B.n233 163.367
R618 B.n233 B.n232 163.367
R619 B.n232 B.n163 163.367
R620 B.n228 B.n163 163.367
R621 B.n228 B.n227 163.367
R622 B.n227 B.n226 163.367
R623 B.n226 B.n165 163.367
R624 B.n222 B.n165 163.367
R625 B.n222 B.n221 163.367
R626 B.n221 B.n220 163.367
R627 B.n220 B.n167 163.367
R628 B.n216 B.n167 163.367
R629 B.n216 B.n215 163.367
R630 B.n215 B.n214 163.367
R631 B.n214 B.n169 163.367
R632 B.n210 B.n169 163.367
R633 B.n210 B.n209 163.367
R634 B.n209 B.n208 163.367
R635 B.n208 B.n171 163.367
R636 B.n204 B.n171 163.367
R637 B.n204 B.n203 163.367
R638 B.n203 B.n202 163.367
R639 B.n202 B.n173 163.367
R640 B.n198 B.n173 163.367
R641 B.n198 B.n197 163.367
R642 B.n197 B.n196 163.367
R643 B.n196 B.n175 163.367
R644 B.n192 B.n175 163.367
R645 B.n192 B.n191 163.367
R646 B.n191 B.n190 163.367
R647 B.n190 B.n177 163.367
R648 B.n186 B.n177 163.367
R649 B.n186 B.n185 163.367
R650 B.n185 B.n184 163.367
R651 B.n184 B.n179 163.367
R652 B.n180 B.n179 163.367
R653 B.n180 B.n2 163.367
R654 B.n690 B.n2 163.367
R655 B.n690 B.n689 163.367
R656 B.n689 B.n688 163.367
R657 B.n688 B.n3 163.367
R658 B.n684 B.n3 163.367
R659 B.n684 B.n683 163.367
R660 B.n683 B.n682 163.367
R661 B.n682 B.n5 163.367
R662 B.n678 B.n5 163.367
R663 B.n678 B.n677 163.367
R664 B.n677 B.n676 163.367
R665 B.n676 B.n7 163.367
R666 B.n672 B.n7 163.367
R667 B.n672 B.n671 163.367
R668 B.n671 B.n670 163.367
R669 B.n670 B.n9 163.367
R670 B.n666 B.n9 163.367
R671 B.n666 B.n665 163.367
R672 B.n665 B.n664 163.367
R673 B.n664 B.n11 163.367
R674 B.n660 B.n11 163.367
R675 B.n660 B.n659 163.367
R676 B.n659 B.n658 163.367
R677 B.n658 B.n13 163.367
R678 B.n654 B.n13 163.367
R679 B.n654 B.n653 163.367
R680 B.n653 B.n652 163.367
R681 B.n652 B.n15 163.367
R682 B.n648 B.n15 163.367
R683 B.n648 B.n647 163.367
R684 B.n647 B.n646 163.367
R685 B.n646 B.n17 163.367
R686 B.n642 B.n17 163.367
R687 B.n642 B.n641 163.367
R688 B.n641 B.n640 163.367
R689 B.n640 B.n19 163.367
R690 B.n636 B.n19 163.367
R691 B.n636 B.n635 163.367
R692 B.n635 B.n634 163.367
R693 B.n634 B.n21 163.367
R694 B.n630 B.n21 163.367
R695 B.n630 B.n629 163.367
R696 B.n240 B.n159 163.367
R697 B.n244 B.n159 163.367
R698 B.n245 B.n244 163.367
R699 B.n246 B.n245 163.367
R700 B.n246 B.n157 163.367
R701 B.n250 B.n157 163.367
R702 B.n251 B.n250 163.367
R703 B.n252 B.n251 163.367
R704 B.n252 B.n155 163.367
R705 B.n256 B.n155 163.367
R706 B.n257 B.n256 163.367
R707 B.n258 B.n257 163.367
R708 B.n258 B.n153 163.367
R709 B.n262 B.n153 163.367
R710 B.n263 B.n262 163.367
R711 B.n264 B.n263 163.367
R712 B.n264 B.n151 163.367
R713 B.n268 B.n151 163.367
R714 B.n269 B.n268 163.367
R715 B.n270 B.n269 163.367
R716 B.n270 B.n149 163.367
R717 B.n274 B.n149 163.367
R718 B.n275 B.n274 163.367
R719 B.n276 B.n275 163.367
R720 B.n276 B.n147 163.367
R721 B.n280 B.n147 163.367
R722 B.n281 B.n280 163.367
R723 B.n282 B.n281 163.367
R724 B.n282 B.n145 163.367
R725 B.n286 B.n145 163.367
R726 B.n287 B.n286 163.367
R727 B.n288 B.n287 163.367
R728 B.n288 B.n143 163.367
R729 B.n292 B.n143 163.367
R730 B.n293 B.n292 163.367
R731 B.n294 B.n293 163.367
R732 B.n294 B.n141 163.367
R733 B.n298 B.n141 163.367
R734 B.n299 B.n298 163.367
R735 B.n299 B.n137 163.367
R736 B.n303 B.n137 163.367
R737 B.n304 B.n303 163.367
R738 B.n305 B.n304 163.367
R739 B.n305 B.n135 163.367
R740 B.n309 B.n135 163.367
R741 B.n310 B.n309 163.367
R742 B.n311 B.n310 163.367
R743 B.n311 B.n131 163.367
R744 B.n316 B.n131 163.367
R745 B.n317 B.n316 163.367
R746 B.n318 B.n317 163.367
R747 B.n318 B.n129 163.367
R748 B.n322 B.n129 163.367
R749 B.n323 B.n322 163.367
R750 B.n324 B.n323 163.367
R751 B.n324 B.n127 163.367
R752 B.n328 B.n127 163.367
R753 B.n329 B.n328 163.367
R754 B.n330 B.n329 163.367
R755 B.n330 B.n125 163.367
R756 B.n334 B.n125 163.367
R757 B.n335 B.n334 163.367
R758 B.n336 B.n335 163.367
R759 B.n336 B.n123 163.367
R760 B.n340 B.n123 163.367
R761 B.n341 B.n340 163.367
R762 B.n342 B.n341 163.367
R763 B.n342 B.n121 163.367
R764 B.n346 B.n121 163.367
R765 B.n347 B.n346 163.367
R766 B.n348 B.n347 163.367
R767 B.n348 B.n119 163.367
R768 B.n352 B.n119 163.367
R769 B.n353 B.n352 163.367
R770 B.n354 B.n353 163.367
R771 B.n354 B.n117 163.367
R772 B.n358 B.n117 163.367
R773 B.n359 B.n358 163.367
R774 B.n360 B.n359 163.367
R775 B.n360 B.n115 163.367
R776 B.n364 B.n115 163.367
R777 B.n365 B.n364 163.367
R778 B.n366 B.n365 163.367
R779 B.n366 B.n113 163.367
R780 B.n370 B.n113 163.367
R781 B.n371 B.n370 163.367
R782 B.n372 B.n111 163.367
R783 B.n376 B.n111 163.367
R784 B.n377 B.n376 163.367
R785 B.n378 B.n377 163.367
R786 B.n378 B.n109 163.367
R787 B.n382 B.n109 163.367
R788 B.n383 B.n382 163.367
R789 B.n384 B.n383 163.367
R790 B.n384 B.n107 163.367
R791 B.n388 B.n107 163.367
R792 B.n389 B.n388 163.367
R793 B.n390 B.n389 163.367
R794 B.n390 B.n105 163.367
R795 B.n394 B.n105 163.367
R796 B.n395 B.n394 163.367
R797 B.n396 B.n395 163.367
R798 B.n396 B.n103 163.367
R799 B.n400 B.n103 163.367
R800 B.n401 B.n400 163.367
R801 B.n402 B.n401 163.367
R802 B.n402 B.n101 163.367
R803 B.n406 B.n101 163.367
R804 B.n407 B.n406 163.367
R805 B.n408 B.n407 163.367
R806 B.n408 B.n99 163.367
R807 B.n412 B.n99 163.367
R808 B.n413 B.n412 163.367
R809 B.n414 B.n413 163.367
R810 B.n414 B.n97 163.367
R811 B.n418 B.n97 163.367
R812 B.n419 B.n418 163.367
R813 B.n420 B.n419 163.367
R814 B.n420 B.n95 163.367
R815 B.n424 B.n95 163.367
R816 B.n425 B.n424 163.367
R817 B.n426 B.n425 163.367
R818 B.n426 B.n93 163.367
R819 B.n430 B.n93 163.367
R820 B.n431 B.n430 163.367
R821 B.n432 B.n431 163.367
R822 B.n432 B.n91 163.367
R823 B.n436 B.n91 163.367
R824 B.n437 B.n436 163.367
R825 B.n438 B.n437 163.367
R826 B.n438 B.n89 163.367
R827 B.n442 B.n89 163.367
R828 B.n443 B.n442 163.367
R829 B.n444 B.n443 163.367
R830 B.n444 B.n87 163.367
R831 B.n448 B.n87 163.367
R832 B.n449 B.n448 163.367
R833 B.n450 B.n449 163.367
R834 B.n450 B.n85 163.367
R835 B.n454 B.n85 163.367
R836 B.n455 B.n454 163.367
R837 B.n456 B.n455 163.367
R838 B.n456 B.n83 163.367
R839 B.n460 B.n83 163.367
R840 B.n461 B.n460 163.367
R841 B.n462 B.n461 163.367
R842 B.n462 B.n81 163.367
R843 B.n466 B.n81 163.367
R844 B.n467 B.n466 163.367
R845 B.n468 B.n467 163.367
R846 B.n468 B.n79 163.367
R847 B.n472 B.n79 163.367
R848 B.n473 B.n472 163.367
R849 B.n474 B.n473 163.367
R850 B.n474 B.n77 163.367
R851 B.n478 B.n77 163.367
R852 B.n479 B.n478 163.367
R853 B.n480 B.n479 163.367
R854 B.n480 B.n75 163.367
R855 B.n484 B.n75 163.367
R856 B.n485 B.n484 163.367
R857 B.n486 B.n485 163.367
R858 B.n486 B.n73 163.367
R859 B.n490 B.n73 163.367
R860 B.n491 B.n490 163.367
R861 B.n492 B.n491 163.367
R862 B.n492 B.n71 163.367
R863 B.n496 B.n71 163.367
R864 B.n628 B.n23 163.367
R865 B.n624 B.n23 163.367
R866 B.n624 B.n623 163.367
R867 B.n623 B.n622 163.367
R868 B.n622 B.n25 163.367
R869 B.n618 B.n25 163.367
R870 B.n618 B.n617 163.367
R871 B.n617 B.n616 163.367
R872 B.n616 B.n27 163.367
R873 B.n612 B.n27 163.367
R874 B.n612 B.n611 163.367
R875 B.n611 B.n610 163.367
R876 B.n610 B.n29 163.367
R877 B.n606 B.n29 163.367
R878 B.n606 B.n605 163.367
R879 B.n605 B.n604 163.367
R880 B.n604 B.n31 163.367
R881 B.n600 B.n31 163.367
R882 B.n600 B.n599 163.367
R883 B.n599 B.n598 163.367
R884 B.n598 B.n33 163.367
R885 B.n594 B.n33 163.367
R886 B.n594 B.n593 163.367
R887 B.n593 B.n592 163.367
R888 B.n592 B.n35 163.367
R889 B.n588 B.n35 163.367
R890 B.n588 B.n587 163.367
R891 B.n587 B.n586 163.367
R892 B.n586 B.n37 163.367
R893 B.n582 B.n37 163.367
R894 B.n582 B.n581 163.367
R895 B.n581 B.n580 163.367
R896 B.n580 B.n39 163.367
R897 B.n576 B.n39 163.367
R898 B.n576 B.n575 163.367
R899 B.n575 B.n574 163.367
R900 B.n574 B.n41 163.367
R901 B.n570 B.n41 163.367
R902 B.n570 B.n569 163.367
R903 B.n569 B.n45 163.367
R904 B.n565 B.n45 163.367
R905 B.n565 B.n564 163.367
R906 B.n564 B.n563 163.367
R907 B.n563 B.n47 163.367
R908 B.n559 B.n47 163.367
R909 B.n559 B.n558 163.367
R910 B.n558 B.n557 163.367
R911 B.n557 B.n49 163.367
R912 B.n552 B.n49 163.367
R913 B.n552 B.n551 163.367
R914 B.n551 B.n550 163.367
R915 B.n550 B.n53 163.367
R916 B.n546 B.n53 163.367
R917 B.n546 B.n545 163.367
R918 B.n545 B.n544 163.367
R919 B.n544 B.n55 163.367
R920 B.n540 B.n55 163.367
R921 B.n540 B.n539 163.367
R922 B.n539 B.n538 163.367
R923 B.n538 B.n57 163.367
R924 B.n534 B.n57 163.367
R925 B.n534 B.n533 163.367
R926 B.n533 B.n532 163.367
R927 B.n532 B.n59 163.367
R928 B.n528 B.n59 163.367
R929 B.n528 B.n527 163.367
R930 B.n527 B.n526 163.367
R931 B.n526 B.n61 163.367
R932 B.n522 B.n61 163.367
R933 B.n522 B.n521 163.367
R934 B.n521 B.n520 163.367
R935 B.n520 B.n63 163.367
R936 B.n516 B.n63 163.367
R937 B.n516 B.n515 163.367
R938 B.n515 B.n514 163.367
R939 B.n514 B.n65 163.367
R940 B.n510 B.n65 163.367
R941 B.n510 B.n509 163.367
R942 B.n509 B.n508 163.367
R943 B.n508 B.n67 163.367
R944 B.n504 B.n67 163.367
R945 B.n504 B.n503 163.367
R946 B.n503 B.n502 163.367
R947 B.n502 B.n69 163.367
R948 B.n498 B.n69 163.367
R949 B.n498 B.n497 163.367
R950 B.n132 B.t5 147.483
R951 B.n50 B.t7 147.483
R952 B.n138 B.t2 147.47
R953 B.n42 B.t10 147.47
R954 B.n133 B.t4 111.216
R955 B.n51 B.t8 111.216
R956 B.n139 B.t1 111.204
R957 B.n43 B.t11 111.204
R958 B.n313 B.n133 59.5399
R959 B.n140 B.n139 59.5399
R960 B.n44 B.n43 59.5399
R961 B.n555 B.n51 59.5399
R962 B.n133 B.n132 36.2672
R963 B.n139 B.n138 36.2672
R964 B.n43 B.n42 36.2672
R965 B.n51 B.n50 36.2672
R966 B.n627 B.n22 35.7468
R967 B.n373 B.n112 35.7468
R968 B.n241 B.n160 35.7468
R969 B.n495 B.n70 35.7468
R970 B B.n691 18.0485
R971 B.n627 B.n626 10.6151
R972 B.n626 B.n625 10.6151
R973 B.n625 B.n24 10.6151
R974 B.n621 B.n24 10.6151
R975 B.n621 B.n620 10.6151
R976 B.n620 B.n619 10.6151
R977 B.n619 B.n26 10.6151
R978 B.n615 B.n26 10.6151
R979 B.n615 B.n614 10.6151
R980 B.n614 B.n613 10.6151
R981 B.n613 B.n28 10.6151
R982 B.n609 B.n28 10.6151
R983 B.n609 B.n608 10.6151
R984 B.n608 B.n607 10.6151
R985 B.n607 B.n30 10.6151
R986 B.n603 B.n30 10.6151
R987 B.n603 B.n602 10.6151
R988 B.n602 B.n601 10.6151
R989 B.n601 B.n32 10.6151
R990 B.n597 B.n32 10.6151
R991 B.n597 B.n596 10.6151
R992 B.n596 B.n595 10.6151
R993 B.n595 B.n34 10.6151
R994 B.n591 B.n34 10.6151
R995 B.n591 B.n590 10.6151
R996 B.n590 B.n589 10.6151
R997 B.n589 B.n36 10.6151
R998 B.n585 B.n36 10.6151
R999 B.n585 B.n584 10.6151
R1000 B.n584 B.n583 10.6151
R1001 B.n583 B.n38 10.6151
R1002 B.n579 B.n38 10.6151
R1003 B.n579 B.n578 10.6151
R1004 B.n578 B.n577 10.6151
R1005 B.n577 B.n40 10.6151
R1006 B.n573 B.n40 10.6151
R1007 B.n573 B.n572 10.6151
R1008 B.n572 B.n571 10.6151
R1009 B.n568 B.n567 10.6151
R1010 B.n567 B.n566 10.6151
R1011 B.n566 B.n46 10.6151
R1012 B.n562 B.n46 10.6151
R1013 B.n562 B.n561 10.6151
R1014 B.n561 B.n560 10.6151
R1015 B.n560 B.n48 10.6151
R1016 B.n556 B.n48 10.6151
R1017 B.n554 B.n553 10.6151
R1018 B.n553 B.n52 10.6151
R1019 B.n549 B.n52 10.6151
R1020 B.n549 B.n548 10.6151
R1021 B.n548 B.n547 10.6151
R1022 B.n547 B.n54 10.6151
R1023 B.n543 B.n54 10.6151
R1024 B.n543 B.n542 10.6151
R1025 B.n542 B.n541 10.6151
R1026 B.n541 B.n56 10.6151
R1027 B.n537 B.n56 10.6151
R1028 B.n537 B.n536 10.6151
R1029 B.n536 B.n535 10.6151
R1030 B.n535 B.n58 10.6151
R1031 B.n531 B.n58 10.6151
R1032 B.n531 B.n530 10.6151
R1033 B.n530 B.n529 10.6151
R1034 B.n529 B.n60 10.6151
R1035 B.n525 B.n60 10.6151
R1036 B.n525 B.n524 10.6151
R1037 B.n524 B.n523 10.6151
R1038 B.n523 B.n62 10.6151
R1039 B.n519 B.n62 10.6151
R1040 B.n519 B.n518 10.6151
R1041 B.n518 B.n517 10.6151
R1042 B.n517 B.n64 10.6151
R1043 B.n513 B.n64 10.6151
R1044 B.n513 B.n512 10.6151
R1045 B.n512 B.n511 10.6151
R1046 B.n511 B.n66 10.6151
R1047 B.n507 B.n66 10.6151
R1048 B.n507 B.n506 10.6151
R1049 B.n506 B.n505 10.6151
R1050 B.n505 B.n68 10.6151
R1051 B.n501 B.n68 10.6151
R1052 B.n501 B.n500 10.6151
R1053 B.n500 B.n499 10.6151
R1054 B.n499 B.n70 10.6151
R1055 B.n374 B.n373 10.6151
R1056 B.n375 B.n374 10.6151
R1057 B.n375 B.n110 10.6151
R1058 B.n379 B.n110 10.6151
R1059 B.n380 B.n379 10.6151
R1060 B.n381 B.n380 10.6151
R1061 B.n381 B.n108 10.6151
R1062 B.n385 B.n108 10.6151
R1063 B.n386 B.n385 10.6151
R1064 B.n387 B.n386 10.6151
R1065 B.n387 B.n106 10.6151
R1066 B.n391 B.n106 10.6151
R1067 B.n392 B.n391 10.6151
R1068 B.n393 B.n392 10.6151
R1069 B.n393 B.n104 10.6151
R1070 B.n397 B.n104 10.6151
R1071 B.n398 B.n397 10.6151
R1072 B.n399 B.n398 10.6151
R1073 B.n399 B.n102 10.6151
R1074 B.n403 B.n102 10.6151
R1075 B.n404 B.n403 10.6151
R1076 B.n405 B.n404 10.6151
R1077 B.n405 B.n100 10.6151
R1078 B.n409 B.n100 10.6151
R1079 B.n410 B.n409 10.6151
R1080 B.n411 B.n410 10.6151
R1081 B.n411 B.n98 10.6151
R1082 B.n415 B.n98 10.6151
R1083 B.n416 B.n415 10.6151
R1084 B.n417 B.n416 10.6151
R1085 B.n417 B.n96 10.6151
R1086 B.n421 B.n96 10.6151
R1087 B.n422 B.n421 10.6151
R1088 B.n423 B.n422 10.6151
R1089 B.n423 B.n94 10.6151
R1090 B.n427 B.n94 10.6151
R1091 B.n428 B.n427 10.6151
R1092 B.n429 B.n428 10.6151
R1093 B.n429 B.n92 10.6151
R1094 B.n433 B.n92 10.6151
R1095 B.n434 B.n433 10.6151
R1096 B.n435 B.n434 10.6151
R1097 B.n435 B.n90 10.6151
R1098 B.n439 B.n90 10.6151
R1099 B.n440 B.n439 10.6151
R1100 B.n441 B.n440 10.6151
R1101 B.n441 B.n88 10.6151
R1102 B.n445 B.n88 10.6151
R1103 B.n446 B.n445 10.6151
R1104 B.n447 B.n446 10.6151
R1105 B.n447 B.n86 10.6151
R1106 B.n451 B.n86 10.6151
R1107 B.n452 B.n451 10.6151
R1108 B.n453 B.n452 10.6151
R1109 B.n453 B.n84 10.6151
R1110 B.n457 B.n84 10.6151
R1111 B.n458 B.n457 10.6151
R1112 B.n459 B.n458 10.6151
R1113 B.n459 B.n82 10.6151
R1114 B.n463 B.n82 10.6151
R1115 B.n464 B.n463 10.6151
R1116 B.n465 B.n464 10.6151
R1117 B.n465 B.n80 10.6151
R1118 B.n469 B.n80 10.6151
R1119 B.n470 B.n469 10.6151
R1120 B.n471 B.n470 10.6151
R1121 B.n471 B.n78 10.6151
R1122 B.n475 B.n78 10.6151
R1123 B.n476 B.n475 10.6151
R1124 B.n477 B.n476 10.6151
R1125 B.n477 B.n76 10.6151
R1126 B.n481 B.n76 10.6151
R1127 B.n482 B.n481 10.6151
R1128 B.n483 B.n482 10.6151
R1129 B.n483 B.n74 10.6151
R1130 B.n487 B.n74 10.6151
R1131 B.n488 B.n487 10.6151
R1132 B.n489 B.n488 10.6151
R1133 B.n489 B.n72 10.6151
R1134 B.n493 B.n72 10.6151
R1135 B.n494 B.n493 10.6151
R1136 B.n495 B.n494 10.6151
R1137 B.n242 B.n241 10.6151
R1138 B.n243 B.n242 10.6151
R1139 B.n243 B.n158 10.6151
R1140 B.n247 B.n158 10.6151
R1141 B.n248 B.n247 10.6151
R1142 B.n249 B.n248 10.6151
R1143 B.n249 B.n156 10.6151
R1144 B.n253 B.n156 10.6151
R1145 B.n254 B.n253 10.6151
R1146 B.n255 B.n254 10.6151
R1147 B.n255 B.n154 10.6151
R1148 B.n259 B.n154 10.6151
R1149 B.n260 B.n259 10.6151
R1150 B.n261 B.n260 10.6151
R1151 B.n261 B.n152 10.6151
R1152 B.n265 B.n152 10.6151
R1153 B.n266 B.n265 10.6151
R1154 B.n267 B.n266 10.6151
R1155 B.n267 B.n150 10.6151
R1156 B.n271 B.n150 10.6151
R1157 B.n272 B.n271 10.6151
R1158 B.n273 B.n272 10.6151
R1159 B.n273 B.n148 10.6151
R1160 B.n277 B.n148 10.6151
R1161 B.n278 B.n277 10.6151
R1162 B.n279 B.n278 10.6151
R1163 B.n279 B.n146 10.6151
R1164 B.n283 B.n146 10.6151
R1165 B.n284 B.n283 10.6151
R1166 B.n285 B.n284 10.6151
R1167 B.n285 B.n144 10.6151
R1168 B.n289 B.n144 10.6151
R1169 B.n290 B.n289 10.6151
R1170 B.n291 B.n290 10.6151
R1171 B.n291 B.n142 10.6151
R1172 B.n295 B.n142 10.6151
R1173 B.n296 B.n295 10.6151
R1174 B.n297 B.n296 10.6151
R1175 B.n301 B.n300 10.6151
R1176 B.n302 B.n301 10.6151
R1177 B.n302 B.n136 10.6151
R1178 B.n306 B.n136 10.6151
R1179 B.n307 B.n306 10.6151
R1180 B.n308 B.n307 10.6151
R1181 B.n308 B.n134 10.6151
R1182 B.n312 B.n134 10.6151
R1183 B.n315 B.n314 10.6151
R1184 B.n315 B.n130 10.6151
R1185 B.n319 B.n130 10.6151
R1186 B.n320 B.n319 10.6151
R1187 B.n321 B.n320 10.6151
R1188 B.n321 B.n128 10.6151
R1189 B.n325 B.n128 10.6151
R1190 B.n326 B.n325 10.6151
R1191 B.n327 B.n326 10.6151
R1192 B.n327 B.n126 10.6151
R1193 B.n331 B.n126 10.6151
R1194 B.n332 B.n331 10.6151
R1195 B.n333 B.n332 10.6151
R1196 B.n333 B.n124 10.6151
R1197 B.n337 B.n124 10.6151
R1198 B.n338 B.n337 10.6151
R1199 B.n339 B.n338 10.6151
R1200 B.n339 B.n122 10.6151
R1201 B.n343 B.n122 10.6151
R1202 B.n344 B.n343 10.6151
R1203 B.n345 B.n344 10.6151
R1204 B.n345 B.n120 10.6151
R1205 B.n349 B.n120 10.6151
R1206 B.n350 B.n349 10.6151
R1207 B.n351 B.n350 10.6151
R1208 B.n351 B.n118 10.6151
R1209 B.n355 B.n118 10.6151
R1210 B.n356 B.n355 10.6151
R1211 B.n357 B.n356 10.6151
R1212 B.n357 B.n116 10.6151
R1213 B.n361 B.n116 10.6151
R1214 B.n362 B.n361 10.6151
R1215 B.n363 B.n362 10.6151
R1216 B.n363 B.n114 10.6151
R1217 B.n367 B.n114 10.6151
R1218 B.n368 B.n367 10.6151
R1219 B.n369 B.n368 10.6151
R1220 B.n369 B.n112 10.6151
R1221 B.n237 B.n160 10.6151
R1222 B.n237 B.n236 10.6151
R1223 B.n236 B.n235 10.6151
R1224 B.n235 B.n162 10.6151
R1225 B.n231 B.n162 10.6151
R1226 B.n231 B.n230 10.6151
R1227 B.n230 B.n229 10.6151
R1228 B.n229 B.n164 10.6151
R1229 B.n225 B.n164 10.6151
R1230 B.n225 B.n224 10.6151
R1231 B.n224 B.n223 10.6151
R1232 B.n223 B.n166 10.6151
R1233 B.n219 B.n166 10.6151
R1234 B.n219 B.n218 10.6151
R1235 B.n218 B.n217 10.6151
R1236 B.n217 B.n168 10.6151
R1237 B.n213 B.n168 10.6151
R1238 B.n213 B.n212 10.6151
R1239 B.n212 B.n211 10.6151
R1240 B.n211 B.n170 10.6151
R1241 B.n207 B.n170 10.6151
R1242 B.n207 B.n206 10.6151
R1243 B.n206 B.n205 10.6151
R1244 B.n205 B.n172 10.6151
R1245 B.n201 B.n172 10.6151
R1246 B.n201 B.n200 10.6151
R1247 B.n200 B.n199 10.6151
R1248 B.n199 B.n174 10.6151
R1249 B.n195 B.n174 10.6151
R1250 B.n195 B.n194 10.6151
R1251 B.n194 B.n193 10.6151
R1252 B.n193 B.n176 10.6151
R1253 B.n189 B.n176 10.6151
R1254 B.n189 B.n188 10.6151
R1255 B.n188 B.n187 10.6151
R1256 B.n187 B.n178 10.6151
R1257 B.n183 B.n178 10.6151
R1258 B.n183 B.n182 10.6151
R1259 B.n182 B.n181 10.6151
R1260 B.n181 B.n0 10.6151
R1261 B.n687 B.n1 10.6151
R1262 B.n687 B.n686 10.6151
R1263 B.n686 B.n685 10.6151
R1264 B.n685 B.n4 10.6151
R1265 B.n681 B.n4 10.6151
R1266 B.n681 B.n680 10.6151
R1267 B.n680 B.n679 10.6151
R1268 B.n679 B.n6 10.6151
R1269 B.n675 B.n6 10.6151
R1270 B.n675 B.n674 10.6151
R1271 B.n674 B.n673 10.6151
R1272 B.n673 B.n8 10.6151
R1273 B.n669 B.n8 10.6151
R1274 B.n669 B.n668 10.6151
R1275 B.n668 B.n667 10.6151
R1276 B.n667 B.n10 10.6151
R1277 B.n663 B.n10 10.6151
R1278 B.n663 B.n662 10.6151
R1279 B.n662 B.n661 10.6151
R1280 B.n661 B.n12 10.6151
R1281 B.n657 B.n12 10.6151
R1282 B.n657 B.n656 10.6151
R1283 B.n656 B.n655 10.6151
R1284 B.n655 B.n14 10.6151
R1285 B.n651 B.n14 10.6151
R1286 B.n651 B.n650 10.6151
R1287 B.n650 B.n649 10.6151
R1288 B.n649 B.n16 10.6151
R1289 B.n645 B.n16 10.6151
R1290 B.n645 B.n644 10.6151
R1291 B.n644 B.n643 10.6151
R1292 B.n643 B.n18 10.6151
R1293 B.n639 B.n18 10.6151
R1294 B.n639 B.n638 10.6151
R1295 B.n638 B.n637 10.6151
R1296 B.n637 B.n20 10.6151
R1297 B.n633 B.n20 10.6151
R1298 B.n633 B.n632 10.6151
R1299 B.n632 B.n631 10.6151
R1300 B.n631 B.n22 10.6151
R1301 B.n568 B.n44 6.5566
R1302 B.n556 B.n555 6.5566
R1303 B.n300 B.n140 6.5566
R1304 B.n313 B.n312 6.5566
R1305 B.n571 B.n44 4.05904
R1306 B.n555 B.n554 4.05904
R1307 B.n297 B.n140 4.05904
R1308 B.n314 B.n313 4.05904
R1309 B.n691 B.n0 2.81026
R1310 B.n691 B.n1 2.81026
C0 VN B 1.00571f
C1 VTAIL B 3.04856f
C2 VN VDD1 0.151225f
C3 VN VP 6.65835f
C4 VTAIL VDD1 10.301201f
C5 VTAIL VP 8.90726f
C6 VN w_n3214_n3184# 6.52073f
C7 VTAIL w_n3214_n3184# 2.94708f
C8 VDD2 B 2.06397f
C9 VDD2 VDD1 1.48473f
C10 VDD2 VP 0.448649f
C11 VTAIL VN 8.89287f
C12 w_n3214_n3184# VDD2 2.40603f
C13 VDD1 B 1.98733f
C14 B VP 1.69801f
C15 w_n3214_n3184# B 8.50603f
C16 VDD1 VP 8.94953f
C17 VN VDD2 8.655941f
C18 w_n3214_n3184# VDD1 2.31751f
C19 VTAIL VDD2 10.3438f
C20 w_n3214_n3184# VP 6.93591f
C21 VDD2 VSUBS 1.731337f
C22 VDD1 VSUBS 1.482542f
C23 VTAIL VSUBS 1.005174f
C24 VN VSUBS 5.95739f
C25 VP VSUBS 2.844309f
C26 B VSUBS 3.973086f
C27 w_n3214_n3184# VSUBS 0.126156p
C28 B.n0 VSUBS 0.005075f
C29 B.n1 VSUBS 0.005075f
C30 B.n2 VSUBS 0.008025f
C31 B.n3 VSUBS 0.008025f
C32 B.n4 VSUBS 0.008025f
C33 B.n5 VSUBS 0.008025f
C34 B.n6 VSUBS 0.008025f
C35 B.n7 VSUBS 0.008025f
C36 B.n8 VSUBS 0.008025f
C37 B.n9 VSUBS 0.008025f
C38 B.n10 VSUBS 0.008025f
C39 B.n11 VSUBS 0.008025f
C40 B.n12 VSUBS 0.008025f
C41 B.n13 VSUBS 0.008025f
C42 B.n14 VSUBS 0.008025f
C43 B.n15 VSUBS 0.008025f
C44 B.n16 VSUBS 0.008025f
C45 B.n17 VSUBS 0.008025f
C46 B.n18 VSUBS 0.008025f
C47 B.n19 VSUBS 0.008025f
C48 B.n20 VSUBS 0.008025f
C49 B.n21 VSUBS 0.008025f
C50 B.n22 VSUBS 0.019596f
C51 B.n23 VSUBS 0.008025f
C52 B.n24 VSUBS 0.008025f
C53 B.n25 VSUBS 0.008025f
C54 B.n26 VSUBS 0.008025f
C55 B.n27 VSUBS 0.008025f
C56 B.n28 VSUBS 0.008025f
C57 B.n29 VSUBS 0.008025f
C58 B.n30 VSUBS 0.008025f
C59 B.n31 VSUBS 0.008025f
C60 B.n32 VSUBS 0.008025f
C61 B.n33 VSUBS 0.008025f
C62 B.n34 VSUBS 0.008025f
C63 B.n35 VSUBS 0.008025f
C64 B.n36 VSUBS 0.008025f
C65 B.n37 VSUBS 0.008025f
C66 B.n38 VSUBS 0.008025f
C67 B.n39 VSUBS 0.008025f
C68 B.n40 VSUBS 0.008025f
C69 B.n41 VSUBS 0.008025f
C70 B.t11 VSUBS 0.410286f
C71 B.t10 VSUBS 0.426455f
C72 B.t9 VSUBS 0.862141f
C73 B.n42 VSUBS 0.193788f
C74 B.n43 VSUBS 0.077191f
C75 B.n44 VSUBS 0.018593f
C76 B.n45 VSUBS 0.008025f
C77 B.n46 VSUBS 0.008025f
C78 B.n47 VSUBS 0.008025f
C79 B.n48 VSUBS 0.008025f
C80 B.n49 VSUBS 0.008025f
C81 B.t8 VSUBS 0.41028f
C82 B.t7 VSUBS 0.426448f
C83 B.t6 VSUBS 0.862141f
C84 B.n50 VSUBS 0.193794f
C85 B.n51 VSUBS 0.077198f
C86 B.n52 VSUBS 0.008025f
C87 B.n53 VSUBS 0.008025f
C88 B.n54 VSUBS 0.008025f
C89 B.n55 VSUBS 0.008025f
C90 B.n56 VSUBS 0.008025f
C91 B.n57 VSUBS 0.008025f
C92 B.n58 VSUBS 0.008025f
C93 B.n59 VSUBS 0.008025f
C94 B.n60 VSUBS 0.008025f
C95 B.n61 VSUBS 0.008025f
C96 B.n62 VSUBS 0.008025f
C97 B.n63 VSUBS 0.008025f
C98 B.n64 VSUBS 0.008025f
C99 B.n65 VSUBS 0.008025f
C100 B.n66 VSUBS 0.008025f
C101 B.n67 VSUBS 0.008025f
C102 B.n68 VSUBS 0.008025f
C103 B.n69 VSUBS 0.008025f
C104 B.n70 VSUBS 0.019427f
C105 B.n71 VSUBS 0.008025f
C106 B.n72 VSUBS 0.008025f
C107 B.n73 VSUBS 0.008025f
C108 B.n74 VSUBS 0.008025f
C109 B.n75 VSUBS 0.008025f
C110 B.n76 VSUBS 0.008025f
C111 B.n77 VSUBS 0.008025f
C112 B.n78 VSUBS 0.008025f
C113 B.n79 VSUBS 0.008025f
C114 B.n80 VSUBS 0.008025f
C115 B.n81 VSUBS 0.008025f
C116 B.n82 VSUBS 0.008025f
C117 B.n83 VSUBS 0.008025f
C118 B.n84 VSUBS 0.008025f
C119 B.n85 VSUBS 0.008025f
C120 B.n86 VSUBS 0.008025f
C121 B.n87 VSUBS 0.008025f
C122 B.n88 VSUBS 0.008025f
C123 B.n89 VSUBS 0.008025f
C124 B.n90 VSUBS 0.008025f
C125 B.n91 VSUBS 0.008025f
C126 B.n92 VSUBS 0.008025f
C127 B.n93 VSUBS 0.008025f
C128 B.n94 VSUBS 0.008025f
C129 B.n95 VSUBS 0.008025f
C130 B.n96 VSUBS 0.008025f
C131 B.n97 VSUBS 0.008025f
C132 B.n98 VSUBS 0.008025f
C133 B.n99 VSUBS 0.008025f
C134 B.n100 VSUBS 0.008025f
C135 B.n101 VSUBS 0.008025f
C136 B.n102 VSUBS 0.008025f
C137 B.n103 VSUBS 0.008025f
C138 B.n104 VSUBS 0.008025f
C139 B.n105 VSUBS 0.008025f
C140 B.n106 VSUBS 0.008025f
C141 B.n107 VSUBS 0.008025f
C142 B.n108 VSUBS 0.008025f
C143 B.n109 VSUBS 0.008025f
C144 B.n110 VSUBS 0.008025f
C145 B.n111 VSUBS 0.008025f
C146 B.n112 VSUBS 0.020294f
C147 B.n113 VSUBS 0.008025f
C148 B.n114 VSUBS 0.008025f
C149 B.n115 VSUBS 0.008025f
C150 B.n116 VSUBS 0.008025f
C151 B.n117 VSUBS 0.008025f
C152 B.n118 VSUBS 0.008025f
C153 B.n119 VSUBS 0.008025f
C154 B.n120 VSUBS 0.008025f
C155 B.n121 VSUBS 0.008025f
C156 B.n122 VSUBS 0.008025f
C157 B.n123 VSUBS 0.008025f
C158 B.n124 VSUBS 0.008025f
C159 B.n125 VSUBS 0.008025f
C160 B.n126 VSUBS 0.008025f
C161 B.n127 VSUBS 0.008025f
C162 B.n128 VSUBS 0.008025f
C163 B.n129 VSUBS 0.008025f
C164 B.n130 VSUBS 0.008025f
C165 B.n131 VSUBS 0.008025f
C166 B.t4 VSUBS 0.41028f
C167 B.t5 VSUBS 0.426448f
C168 B.t3 VSUBS 0.862141f
C169 B.n132 VSUBS 0.193794f
C170 B.n133 VSUBS 0.077198f
C171 B.n134 VSUBS 0.008025f
C172 B.n135 VSUBS 0.008025f
C173 B.n136 VSUBS 0.008025f
C174 B.n137 VSUBS 0.008025f
C175 B.t1 VSUBS 0.410286f
C176 B.t2 VSUBS 0.426455f
C177 B.t0 VSUBS 0.862141f
C178 B.n138 VSUBS 0.193788f
C179 B.n139 VSUBS 0.077191f
C180 B.n140 VSUBS 0.018593f
C181 B.n141 VSUBS 0.008025f
C182 B.n142 VSUBS 0.008025f
C183 B.n143 VSUBS 0.008025f
C184 B.n144 VSUBS 0.008025f
C185 B.n145 VSUBS 0.008025f
C186 B.n146 VSUBS 0.008025f
C187 B.n147 VSUBS 0.008025f
C188 B.n148 VSUBS 0.008025f
C189 B.n149 VSUBS 0.008025f
C190 B.n150 VSUBS 0.008025f
C191 B.n151 VSUBS 0.008025f
C192 B.n152 VSUBS 0.008025f
C193 B.n153 VSUBS 0.008025f
C194 B.n154 VSUBS 0.008025f
C195 B.n155 VSUBS 0.008025f
C196 B.n156 VSUBS 0.008025f
C197 B.n157 VSUBS 0.008025f
C198 B.n158 VSUBS 0.008025f
C199 B.n159 VSUBS 0.008025f
C200 B.n160 VSUBS 0.019596f
C201 B.n161 VSUBS 0.008025f
C202 B.n162 VSUBS 0.008025f
C203 B.n163 VSUBS 0.008025f
C204 B.n164 VSUBS 0.008025f
C205 B.n165 VSUBS 0.008025f
C206 B.n166 VSUBS 0.008025f
C207 B.n167 VSUBS 0.008025f
C208 B.n168 VSUBS 0.008025f
C209 B.n169 VSUBS 0.008025f
C210 B.n170 VSUBS 0.008025f
C211 B.n171 VSUBS 0.008025f
C212 B.n172 VSUBS 0.008025f
C213 B.n173 VSUBS 0.008025f
C214 B.n174 VSUBS 0.008025f
C215 B.n175 VSUBS 0.008025f
C216 B.n176 VSUBS 0.008025f
C217 B.n177 VSUBS 0.008025f
C218 B.n178 VSUBS 0.008025f
C219 B.n179 VSUBS 0.008025f
C220 B.n180 VSUBS 0.008025f
C221 B.n181 VSUBS 0.008025f
C222 B.n182 VSUBS 0.008025f
C223 B.n183 VSUBS 0.008025f
C224 B.n184 VSUBS 0.008025f
C225 B.n185 VSUBS 0.008025f
C226 B.n186 VSUBS 0.008025f
C227 B.n187 VSUBS 0.008025f
C228 B.n188 VSUBS 0.008025f
C229 B.n189 VSUBS 0.008025f
C230 B.n190 VSUBS 0.008025f
C231 B.n191 VSUBS 0.008025f
C232 B.n192 VSUBS 0.008025f
C233 B.n193 VSUBS 0.008025f
C234 B.n194 VSUBS 0.008025f
C235 B.n195 VSUBS 0.008025f
C236 B.n196 VSUBS 0.008025f
C237 B.n197 VSUBS 0.008025f
C238 B.n198 VSUBS 0.008025f
C239 B.n199 VSUBS 0.008025f
C240 B.n200 VSUBS 0.008025f
C241 B.n201 VSUBS 0.008025f
C242 B.n202 VSUBS 0.008025f
C243 B.n203 VSUBS 0.008025f
C244 B.n204 VSUBS 0.008025f
C245 B.n205 VSUBS 0.008025f
C246 B.n206 VSUBS 0.008025f
C247 B.n207 VSUBS 0.008025f
C248 B.n208 VSUBS 0.008025f
C249 B.n209 VSUBS 0.008025f
C250 B.n210 VSUBS 0.008025f
C251 B.n211 VSUBS 0.008025f
C252 B.n212 VSUBS 0.008025f
C253 B.n213 VSUBS 0.008025f
C254 B.n214 VSUBS 0.008025f
C255 B.n215 VSUBS 0.008025f
C256 B.n216 VSUBS 0.008025f
C257 B.n217 VSUBS 0.008025f
C258 B.n218 VSUBS 0.008025f
C259 B.n219 VSUBS 0.008025f
C260 B.n220 VSUBS 0.008025f
C261 B.n221 VSUBS 0.008025f
C262 B.n222 VSUBS 0.008025f
C263 B.n223 VSUBS 0.008025f
C264 B.n224 VSUBS 0.008025f
C265 B.n225 VSUBS 0.008025f
C266 B.n226 VSUBS 0.008025f
C267 B.n227 VSUBS 0.008025f
C268 B.n228 VSUBS 0.008025f
C269 B.n229 VSUBS 0.008025f
C270 B.n230 VSUBS 0.008025f
C271 B.n231 VSUBS 0.008025f
C272 B.n232 VSUBS 0.008025f
C273 B.n233 VSUBS 0.008025f
C274 B.n234 VSUBS 0.008025f
C275 B.n235 VSUBS 0.008025f
C276 B.n236 VSUBS 0.008025f
C277 B.n237 VSUBS 0.008025f
C278 B.n238 VSUBS 0.008025f
C279 B.n239 VSUBS 0.019596f
C280 B.n240 VSUBS 0.020294f
C281 B.n241 VSUBS 0.020294f
C282 B.n242 VSUBS 0.008025f
C283 B.n243 VSUBS 0.008025f
C284 B.n244 VSUBS 0.008025f
C285 B.n245 VSUBS 0.008025f
C286 B.n246 VSUBS 0.008025f
C287 B.n247 VSUBS 0.008025f
C288 B.n248 VSUBS 0.008025f
C289 B.n249 VSUBS 0.008025f
C290 B.n250 VSUBS 0.008025f
C291 B.n251 VSUBS 0.008025f
C292 B.n252 VSUBS 0.008025f
C293 B.n253 VSUBS 0.008025f
C294 B.n254 VSUBS 0.008025f
C295 B.n255 VSUBS 0.008025f
C296 B.n256 VSUBS 0.008025f
C297 B.n257 VSUBS 0.008025f
C298 B.n258 VSUBS 0.008025f
C299 B.n259 VSUBS 0.008025f
C300 B.n260 VSUBS 0.008025f
C301 B.n261 VSUBS 0.008025f
C302 B.n262 VSUBS 0.008025f
C303 B.n263 VSUBS 0.008025f
C304 B.n264 VSUBS 0.008025f
C305 B.n265 VSUBS 0.008025f
C306 B.n266 VSUBS 0.008025f
C307 B.n267 VSUBS 0.008025f
C308 B.n268 VSUBS 0.008025f
C309 B.n269 VSUBS 0.008025f
C310 B.n270 VSUBS 0.008025f
C311 B.n271 VSUBS 0.008025f
C312 B.n272 VSUBS 0.008025f
C313 B.n273 VSUBS 0.008025f
C314 B.n274 VSUBS 0.008025f
C315 B.n275 VSUBS 0.008025f
C316 B.n276 VSUBS 0.008025f
C317 B.n277 VSUBS 0.008025f
C318 B.n278 VSUBS 0.008025f
C319 B.n279 VSUBS 0.008025f
C320 B.n280 VSUBS 0.008025f
C321 B.n281 VSUBS 0.008025f
C322 B.n282 VSUBS 0.008025f
C323 B.n283 VSUBS 0.008025f
C324 B.n284 VSUBS 0.008025f
C325 B.n285 VSUBS 0.008025f
C326 B.n286 VSUBS 0.008025f
C327 B.n287 VSUBS 0.008025f
C328 B.n288 VSUBS 0.008025f
C329 B.n289 VSUBS 0.008025f
C330 B.n290 VSUBS 0.008025f
C331 B.n291 VSUBS 0.008025f
C332 B.n292 VSUBS 0.008025f
C333 B.n293 VSUBS 0.008025f
C334 B.n294 VSUBS 0.008025f
C335 B.n295 VSUBS 0.008025f
C336 B.n296 VSUBS 0.008025f
C337 B.n297 VSUBS 0.005547f
C338 B.n298 VSUBS 0.008025f
C339 B.n299 VSUBS 0.008025f
C340 B.n300 VSUBS 0.006491f
C341 B.n301 VSUBS 0.008025f
C342 B.n302 VSUBS 0.008025f
C343 B.n303 VSUBS 0.008025f
C344 B.n304 VSUBS 0.008025f
C345 B.n305 VSUBS 0.008025f
C346 B.n306 VSUBS 0.008025f
C347 B.n307 VSUBS 0.008025f
C348 B.n308 VSUBS 0.008025f
C349 B.n309 VSUBS 0.008025f
C350 B.n310 VSUBS 0.008025f
C351 B.n311 VSUBS 0.008025f
C352 B.n312 VSUBS 0.006491f
C353 B.n313 VSUBS 0.018593f
C354 B.n314 VSUBS 0.005547f
C355 B.n315 VSUBS 0.008025f
C356 B.n316 VSUBS 0.008025f
C357 B.n317 VSUBS 0.008025f
C358 B.n318 VSUBS 0.008025f
C359 B.n319 VSUBS 0.008025f
C360 B.n320 VSUBS 0.008025f
C361 B.n321 VSUBS 0.008025f
C362 B.n322 VSUBS 0.008025f
C363 B.n323 VSUBS 0.008025f
C364 B.n324 VSUBS 0.008025f
C365 B.n325 VSUBS 0.008025f
C366 B.n326 VSUBS 0.008025f
C367 B.n327 VSUBS 0.008025f
C368 B.n328 VSUBS 0.008025f
C369 B.n329 VSUBS 0.008025f
C370 B.n330 VSUBS 0.008025f
C371 B.n331 VSUBS 0.008025f
C372 B.n332 VSUBS 0.008025f
C373 B.n333 VSUBS 0.008025f
C374 B.n334 VSUBS 0.008025f
C375 B.n335 VSUBS 0.008025f
C376 B.n336 VSUBS 0.008025f
C377 B.n337 VSUBS 0.008025f
C378 B.n338 VSUBS 0.008025f
C379 B.n339 VSUBS 0.008025f
C380 B.n340 VSUBS 0.008025f
C381 B.n341 VSUBS 0.008025f
C382 B.n342 VSUBS 0.008025f
C383 B.n343 VSUBS 0.008025f
C384 B.n344 VSUBS 0.008025f
C385 B.n345 VSUBS 0.008025f
C386 B.n346 VSUBS 0.008025f
C387 B.n347 VSUBS 0.008025f
C388 B.n348 VSUBS 0.008025f
C389 B.n349 VSUBS 0.008025f
C390 B.n350 VSUBS 0.008025f
C391 B.n351 VSUBS 0.008025f
C392 B.n352 VSUBS 0.008025f
C393 B.n353 VSUBS 0.008025f
C394 B.n354 VSUBS 0.008025f
C395 B.n355 VSUBS 0.008025f
C396 B.n356 VSUBS 0.008025f
C397 B.n357 VSUBS 0.008025f
C398 B.n358 VSUBS 0.008025f
C399 B.n359 VSUBS 0.008025f
C400 B.n360 VSUBS 0.008025f
C401 B.n361 VSUBS 0.008025f
C402 B.n362 VSUBS 0.008025f
C403 B.n363 VSUBS 0.008025f
C404 B.n364 VSUBS 0.008025f
C405 B.n365 VSUBS 0.008025f
C406 B.n366 VSUBS 0.008025f
C407 B.n367 VSUBS 0.008025f
C408 B.n368 VSUBS 0.008025f
C409 B.n369 VSUBS 0.008025f
C410 B.n370 VSUBS 0.008025f
C411 B.n371 VSUBS 0.020294f
C412 B.n372 VSUBS 0.019596f
C413 B.n373 VSUBS 0.019596f
C414 B.n374 VSUBS 0.008025f
C415 B.n375 VSUBS 0.008025f
C416 B.n376 VSUBS 0.008025f
C417 B.n377 VSUBS 0.008025f
C418 B.n378 VSUBS 0.008025f
C419 B.n379 VSUBS 0.008025f
C420 B.n380 VSUBS 0.008025f
C421 B.n381 VSUBS 0.008025f
C422 B.n382 VSUBS 0.008025f
C423 B.n383 VSUBS 0.008025f
C424 B.n384 VSUBS 0.008025f
C425 B.n385 VSUBS 0.008025f
C426 B.n386 VSUBS 0.008025f
C427 B.n387 VSUBS 0.008025f
C428 B.n388 VSUBS 0.008025f
C429 B.n389 VSUBS 0.008025f
C430 B.n390 VSUBS 0.008025f
C431 B.n391 VSUBS 0.008025f
C432 B.n392 VSUBS 0.008025f
C433 B.n393 VSUBS 0.008025f
C434 B.n394 VSUBS 0.008025f
C435 B.n395 VSUBS 0.008025f
C436 B.n396 VSUBS 0.008025f
C437 B.n397 VSUBS 0.008025f
C438 B.n398 VSUBS 0.008025f
C439 B.n399 VSUBS 0.008025f
C440 B.n400 VSUBS 0.008025f
C441 B.n401 VSUBS 0.008025f
C442 B.n402 VSUBS 0.008025f
C443 B.n403 VSUBS 0.008025f
C444 B.n404 VSUBS 0.008025f
C445 B.n405 VSUBS 0.008025f
C446 B.n406 VSUBS 0.008025f
C447 B.n407 VSUBS 0.008025f
C448 B.n408 VSUBS 0.008025f
C449 B.n409 VSUBS 0.008025f
C450 B.n410 VSUBS 0.008025f
C451 B.n411 VSUBS 0.008025f
C452 B.n412 VSUBS 0.008025f
C453 B.n413 VSUBS 0.008025f
C454 B.n414 VSUBS 0.008025f
C455 B.n415 VSUBS 0.008025f
C456 B.n416 VSUBS 0.008025f
C457 B.n417 VSUBS 0.008025f
C458 B.n418 VSUBS 0.008025f
C459 B.n419 VSUBS 0.008025f
C460 B.n420 VSUBS 0.008025f
C461 B.n421 VSUBS 0.008025f
C462 B.n422 VSUBS 0.008025f
C463 B.n423 VSUBS 0.008025f
C464 B.n424 VSUBS 0.008025f
C465 B.n425 VSUBS 0.008025f
C466 B.n426 VSUBS 0.008025f
C467 B.n427 VSUBS 0.008025f
C468 B.n428 VSUBS 0.008025f
C469 B.n429 VSUBS 0.008025f
C470 B.n430 VSUBS 0.008025f
C471 B.n431 VSUBS 0.008025f
C472 B.n432 VSUBS 0.008025f
C473 B.n433 VSUBS 0.008025f
C474 B.n434 VSUBS 0.008025f
C475 B.n435 VSUBS 0.008025f
C476 B.n436 VSUBS 0.008025f
C477 B.n437 VSUBS 0.008025f
C478 B.n438 VSUBS 0.008025f
C479 B.n439 VSUBS 0.008025f
C480 B.n440 VSUBS 0.008025f
C481 B.n441 VSUBS 0.008025f
C482 B.n442 VSUBS 0.008025f
C483 B.n443 VSUBS 0.008025f
C484 B.n444 VSUBS 0.008025f
C485 B.n445 VSUBS 0.008025f
C486 B.n446 VSUBS 0.008025f
C487 B.n447 VSUBS 0.008025f
C488 B.n448 VSUBS 0.008025f
C489 B.n449 VSUBS 0.008025f
C490 B.n450 VSUBS 0.008025f
C491 B.n451 VSUBS 0.008025f
C492 B.n452 VSUBS 0.008025f
C493 B.n453 VSUBS 0.008025f
C494 B.n454 VSUBS 0.008025f
C495 B.n455 VSUBS 0.008025f
C496 B.n456 VSUBS 0.008025f
C497 B.n457 VSUBS 0.008025f
C498 B.n458 VSUBS 0.008025f
C499 B.n459 VSUBS 0.008025f
C500 B.n460 VSUBS 0.008025f
C501 B.n461 VSUBS 0.008025f
C502 B.n462 VSUBS 0.008025f
C503 B.n463 VSUBS 0.008025f
C504 B.n464 VSUBS 0.008025f
C505 B.n465 VSUBS 0.008025f
C506 B.n466 VSUBS 0.008025f
C507 B.n467 VSUBS 0.008025f
C508 B.n468 VSUBS 0.008025f
C509 B.n469 VSUBS 0.008025f
C510 B.n470 VSUBS 0.008025f
C511 B.n471 VSUBS 0.008025f
C512 B.n472 VSUBS 0.008025f
C513 B.n473 VSUBS 0.008025f
C514 B.n474 VSUBS 0.008025f
C515 B.n475 VSUBS 0.008025f
C516 B.n476 VSUBS 0.008025f
C517 B.n477 VSUBS 0.008025f
C518 B.n478 VSUBS 0.008025f
C519 B.n479 VSUBS 0.008025f
C520 B.n480 VSUBS 0.008025f
C521 B.n481 VSUBS 0.008025f
C522 B.n482 VSUBS 0.008025f
C523 B.n483 VSUBS 0.008025f
C524 B.n484 VSUBS 0.008025f
C525 B.n485 VSUBS 0.008025f
C526 B.n486 VSUBS 0.008025f
C527 B.n487 VSUBS 0.008025f
C528 B.n488 VSUBS 0.008025f
C529 B.n489 VSUBS 0.008025f
C530 B.n490 VSUBS 0.008025f
C531 B.n491 VSUBS 0.008025f
C532 B.n492 VSUBS 0.008025f
C533 B.n493 VSUBS 0.008025f
C534 B.n494 VSUBS 0.008025f
C535 B.n495 VSUBS 0.020463f
C536 B.n496 VSUBS 0.019596f
C537 B.n497 VSUBS 0.020294f
C538 B.n498 VSUBS 0.008025f
C539 B.n499 VSUBS 0.008025f
C540 B.n500 VSUBS 0.008025f
C541 B.n501 VSUBS 0.008025f
C542 B.n502 VSUBS 0.008025f
C543 B.n503 VSUBS 0.008025f
C544 B.n504 VSUBS 0.008025f
C545 B.n505 VSUBS 0.008025f
C546 B.n506 VSUBS 0.008025f
C547 B.n507 VSUBS 0.008025f
C548 B.n508 VSUBS 0.008025f
C549 B.n509 VSUBS 0.008025f
C550 B.n510 VSUBS 0.008025f
C551 B.n511 VSUBS 0.008025f
C552 B.n512 VSUBS 0.008025f
C553 B.n513 VSUBS 0.008025f
C554 B.n514 VSUBS 0.008025f
C555 B.n515 VSUBS 0.008025f
C556 B.n516 VSUBS 0.008025f
C557 B.n517 VSUBS 0.008025f
C558 B.n518 VSUBS 0.008025f
C559 B.n519 VSUBS 0.008025f
C560 B.n520 VSUBS 0.008025f
C561 B.n521 VSUBS 0.008025f
C562 B.n522 VSUBS 0.008025f
C563 B.n523 VSUBS 0.008025f
C564 B.n524 VSUBS 0.008025f
C565 B.n525 VSUBS 0.008025f
C566 B.n526 VSUBS 0.008025f
C567 B.n527 VSUBS 0.008025f
C568 B.n528 VSUBS 0.008025f
C569 B.n529 VSUBS 0.008025f
C570 B.n530 VSUBS 0.008025f
C571 B.n531 VSUBS 0.008025f
C572 B.n532 VSUBS 0.008025f
C573 B.n533 VSUBS 0.008025f
C574 B.n534 VSUBS 0.008025f
C575 B.n535 VSUBS 0.008025f
C576 B.n536 VSUBS 0.008025f
C577 B.n537 VSUBS 0.008025f
C578 B.n538 VSUBS 0.008025f
C579 B.n539 VSUBS 0.008025f
C580 B.n540 VSUBS 0.008025f
C581 B.n541 VSUBS 0.008025f
C582 B.n542 VSUBS 0.008025f
C583 B.n543 VSUBS 0.008025f
C584 B.n544 VSUBS 0.008025f
C585 B.n545 VSUBS 0.008025f
C586 B.n546 VSUBS 0.008025f
C587 B.n547 VSUBS 0.008025f
C588 B.n548 VSUBS 0.008025f
C589 B.n549 VSUBS 0.008025f
C590 B.n550 VSUBS 0.008025f
C591 B.n551 VSUBS 0.008025f
C592 B.n552 VSUBS 0.008025f
C593 B.n553 VSUBS 0.008025f
C594 B.n554 VSUBS 0.005547f
C595 B.n555 VSUBS 0.018593f
C596 B.n556 VSUBS 0.006491f
C597 B.n557 VSUBS 0.008025f
C598 B.n558 VSUBS 0.008025f
C599 B.n559 VSUBS 0.008025f
C600 B.n560 VSUBS 0.008025f
C601 B.n561 VSUBS 0.008025f
C602 B.n562 VSUBS 0.008025f
C603 B.n563 VSUBS 0.008025f
C604 B.n564 VSUBS 0.008025f
C605 B.n565 VSUBS 0.008025f
C606 B.n566 VSUBS 0.008025f
C607 B.n567 VSUBS 0.008025f
C608 B.n568 VSUBS 0.006491f
C609 B.n569 VSUBS 0.008025f
C610 B.n570 VSUBS 0.008025f
C611 B.n571 VSUBS 0.005547f
C612 B.n572 VSUBS 0.008025f
C613 B.n573 VSUBS 0.008025f
C614 B.n574 VSUBS 0.008025f
C615 B.n575 VSUBS 0.008025f
C616 B.n576 VSUBS 0.008025f
C617 B.n577 VSUBS 0.008025f
C618 B.n578 VSUBS 0.008025f
C619 B.n579 VSUBS 0.008025f
C620 B.n580 VSUBS 0.008025f
C621 B.n581 VSUBS 0.008025f
C622 B.n582 VSUBS 0.008025f
C623 B.n583 VSUBS 0.008025f
C624 B.n584 VSUBS 0.008025f
C625 B.n585 VSUBS 0.008025f
C626 B.n586 VSUBS 0.008025f
C627 B.n587 VSUBS 0.008025f
C628 B.n588 VSUBS 0.008025f
C629 B.n589 VSUBS 0.008025f
C630 B.n590 VSUBS 0.008025f
C631 B.n591 VSUBS 0.008025f
C632 B.n592 VSUBS 0.008025f
C633 B.n593 VSUBS 0.008025f
C634 B.n594 VSUBS 0.008025f
C635 B.n595 VSUBS 0.008025f
C636 B.n596 VSUBS 0.008025f
C637 B.n597 VSUBS 0.008025f
C638 B.n598 VSUBS 0.008025f
C639 B.n599 VSUBS 0.008025f
C640 B.n600 VSUBS 0.008025f
C641 B.n601 VSUBS 0.008025f
C642 B.n602 VSUBS 0.008025f
C643 B.n603 VSUBS 0.008025f
C644 B.n604 VSUBS 0.008025f
C645 B.n605 VSUBS 0.008025f
C646 B.n606 VSUBS 0.008025f
C647 B.n607 VSUBS 0.008025f
C648 B.n608 VSUBS 0.008025f
C649 B.n609 VSUBS 0.008025f
C650 B.n610 VSUBS 0.008025f
C651 B.n611 VSUBS 0.008025f
C652 B.n612 VSUBS 0.008025f
C653 B.n613 VSUBS 0.008025f
C654 B.n614 VSUBS 0.008025f
C655 B.n615 VSUBS 0.008025f
C656 B.n616 VSUBS 0.008025f
C657 B.n617 VSUBS 0.008025f
C658 B.n618 VSUBS 0.008025f
C659 B.n619 VSUBS 0.008025f
C660 B.n620 VSUBS 0.008025f
C661 B.n621 VSUBS 0.008025f
C662 B.n622 VSUBS 0.008025f
C663 B.n623 VSUBS 0.008025f
C664 B.n624 VSUBS 0.008025f
C665 B.n625 VSUBS 0.008025f
C666 B.n626 VSUBS 0.008025f
C667 B.n627 VSUBS 0.020294f
C668 B.n628 VSUBS 0.020294f
C669 B.n629 VSUBS 0.019596f
C670 B.n630 VSUBS 0.008025f
C671 B.n631 VSUBS 0.008025f
C672 B.n632 VSUBS 0.008025f
C673 B.n633 VSUBS 0.008025f
C674 B.n634 VSUBS 0.008025f
C675 B.n635 VSUBS 0.008025f
C676 B.n636 VSUBS 0.008025f
C677 B.n637 VSUBS 0.008025f
C678 B.n638 VSUBS 0.008025f
C679 B.n639 VSUBS 0.008025f
C680 B.n640 VSUBS 0.008025f
C681 B.n641 VSUBS 0.008025f
C682 B.n642 VSUBS 0.008025f
C683 B.n643 VSUBS 0.008025f
C684 B.n644 VSUBS 0.008025f
C685 B.n645 VSUBS 0.008025f
C686 B.n646 VSUBS 0.008025f
C687 B.n647 VSUBS 0.008025f
C688 B.n648 VSUBS 0.008025f
C689 B.n649 VSUBS 0.008025f
C690 B.n650 VSUBS 0.008025f
C691 B.n651 VSUBS 0.008025f
C692 B.n652 VSUBS 0.008025f
C693 B.n653 VSUBS 0.008025f
C694 B.n654 VSUBS 0.008025f
C695 B.n655 VSUBS 0.008025f
C696 B.n656 VSUBS 0.008025f
C697 B.n657 VSUBS 0.008025f
C698 B.n658 VSUBS 0.008025f
C699 B.n659 VSUBS 0.008025f
C700 B.n660 VSUBS 0.008025f
C701 B.n661 VSUBS 0.008025f
C702 B.n662 VSUBS 0.008025f
C703 B.n663 VSUBS 0.008025f
C704 B.n664 VSUBS 0.008025f
C705 B.n665 VSUBS 0.008025f
C706 B.n666 VSUBS 0.008025f
C707 B.n667 VSUBS 0.008025f
C708 B.n668 VSUBS 0.008025f
C709 B.n669 VSUBS 0.008025f
C710 B.n670 VSUBS 0.008025f
C711 B.n671 VSUBS 0.008025f
C712 B.n672 VSUBS 0.008025f
C713 B.n673 VSUBS 0.008025f
C714 B.n674 VSUBS 0.008025f
C715 B.n675 VSUBS 0.008025f
C716 B.n676 VSUBS 0.008025f
C717 B.n677 VSUBS 0.008025f
C718 B.n678 VSUBS 0.008025f
C719 B.n679 VSUBS 0.008025f
C720 B.n680 VSUBS 0.008025f
C721 B.n681 VSUBS 0.008025f
C722 B.n682 VSUBS 0.008025f
C723 B.n683 VSUBS 0.008025f
C724 B.n684 VSUBS 0.008025f
C725 B.n685 VSUBS 0.008025f
C726 B.n686 VSUBS 0.008025f
C727 B.n687 VSUBS 0.008025f
C728 B.n688 VSUBS 0.008025f
C729 B.n689 VSUBS 0.008025f
C730 B.n690 VSUBS 0.008025f
C731 B.n691 VSUBS 0.018172f
C732 VDD2.t1 VSUBS 2.47115f
C733 VDD2.t3 VSUBS 0.243598f
C734 VDD2.t5 VSUBS 0.243598f
C735 VDD2.n0 VSUBS 1.87706f
C736 VDD2.n1 VSUBS 1.42673f
C737 VDD2.t8 VSUBS 0.243598f
C738 VDD2.t4 VSUBS 0.243598f
C739 VDD2.n2 VSUBS 1.88858f
C740 VDD2.n3 VSUBS 2.83151f
C741 VDD2.t7 VSUBS 2.45611f
C742 VDD2.n4 VSUBS 3.23348f
C743 VDD2.t9 VSUBS 0.243598f
C744 VDD2.t2 VSUBS 0.243598f
C745 VDD2.n5 VSUBS 1.87707f
C746 VDD2.n6 VSUBS 0.697458f
C747 VDD2.t0 VSUBS 0.243598f
C748 VDD2.t6 VSUBS 0.243598f
C749 VDD2.n7 VSUBS 1.88854f
C750 VN.n0 VSUBS 0.037739f
C751 VN.t5 VSUBS 1.75034f
C752 VN.n1 VSUBS 0.060602f
C753 VN.n2 VSUBS 0.037739f
C754 VN.t1 VSUBS 1.75034f
C755 VN.n3 VSUBS 0.071297f
C756 VN.n4 VSUBS 0.037739f
C757 VN.t4 VSUBS 1.75034f
C758 VN.n5 VSUBS 0.066859f
C759 VN.t8 VSUBS 1.88147f
C760 VN.t6 VSUBS 1.75034f
C761 VN.n6 VSUBS 0.715624f
C762 VN.n7 VSUBS 0.718526f
C763 VN.n8 VSUBS 0.240924f
C764 VN.n9 VSUBS 0.037739f
C765 VN.n10 VSUBS 0.032563f
C766 VN.n11 VSUBS 0.071297f
C767 VN.n12 VSUBS 0.671527f
C768 VN.n13 VSUBS 0.037739f
C769 VN.n14 VSUBS 0.037739f
C770 VN.n15 VSUBS 0.037739f
C771 VN.n16 VSUBS 0.032563f
C772 VN.n17 VSUBS 0.066859f
C773 VN.n18 VSUBS 0.636093f
C774 VN.n19 VSUBS 0.044417f
C775 VN.n20 VSUBS 0.037739f
C776 VN.n21 VSUBS 0.037739f
C777 VN.n22 VSUBS 0.037739f
C778 VN.n23 VSUBS 0.049116f
C779 VN.n24 VSUBS 0.052018f
C780 VN.n25 VSUBS 0.718861f
C781 VN.n26 VSUBS 0.035808f
C782 VN.n27 VSUBS 0.037739f
C783 VN.t2 VSUBS 1.75034f
C784 VN.n28 VSUBS 0.060602f
C785 VN.n29 VSUBS 0.037739f
C786 VN.t0 VSUBS 1.75034f
C787 VN.n30 VSUBS 0.071297f
C788 VN.n31 VSUBS 0.037739f
C789 VN.t7 VSUBS 1.75034f
C790 VN.n32 VSUBS 0.066859f
C791 VN.t3 VSUBS 1.88147f
C792 VN.t9 VSUBS 1.75034f
C793 VN.n33 VSUBS 0.715624f
C794 VN.n34 VSUBS 0.718526f
C795 VN.n35 VSUBS 0.240924f
C796 VN.n36 VSUBS 0.037739f
C797 VN.n37 VSUBS 0.032563f
C798 VN.n38 VSUBS 0.071297f
C799 VN.n39 VSUBS 0.671527f
C800 VN.n40 VSUBS 0.037739f
C801 VN.n41 VSUBS 0.037739f
C802 VN.n42 VSUBS 0.037739f
C803 VN.n43 VSUBS 0.032563f
C804 VN.n44 VSUBS 0.066859f
C805 VN.n45 VSUBS 0.636093f
C806 VN.n46 VSUBS 0.044417f
C807 VN.n47 VSUBS 0.037739f
C808 VN.n48 VSUBS 0.037739f
C809 VN.n49 VSUBS 0.037739f
C810 VN.n50 VSUBS 0.049116f
C811 VN.n51 VSUBS 0.052018f
C812 VN.n52 VSUBS 0.718861f
C813 VN.n53 VSUBS 1.87415f
C814 VDD1.t1 VSUBS 2.25101f
C815 VDD1.t7 VSUBS 0.221896f
C816 VDD1.t9 VSUBS 0.221896f
C817 VDD1.n0 VSUBS 1.70984f
C818 VDD1.n1 VSUBS 1.30719f
C819 VDD1.t0 VSUBS 2.25099f
C820 VDD1.t3 VSUBS 0.221896f
C821 VDD1.t2 VSUBS 0.221896f
C822 VDD1.n2 VSUBS 1.70983f
C823 VDD1.n3 VSUBS 1.29963f
C824 VDD1.t6 VSUBS 0.221896f
C825 VDD1.t8 VSUBS 0.221896f
C826 VDD1.n4 VSUBS 1.72033f
C827 VDD1.n5 VSUBS 2.67754f
C828 VDD1.t5 VSUBS 0.221896f
C829 VDD1.t4 VSUBS 0.221896f
C830 VDD1.n6 VSUBS 1.70983f
C831 VDD1.n7 VSUBS 2.95701f
C832 VTAIL.t8 VSUBS 0.249f
C833 VTAIL.t2 VSUBS 0.249f
C834 VTAIL.n0 VSUBS 1.77338f
C835 VTAIL.n1 VSUBS 0.862645f
C836 VTAIL.t17 VSUBS 2.34876f
C837 VTAIL.n2 VSUBS 0.997949f
C838 VTAIL.t11 VSUBS 0.249f
C839 VTAIL.t19 VSUBS 0.249f
C840 VTAIL.n3 VSUBS 1.77338f
C841 VTAIL.n4 VSUBS 0.925051f
C842 VTAIL.t16 VSUBS 0.249f
C843 VTAIL.t14 VSUBS 0.249f
C844 VTAIL.n5 VSUBS 1.77338f
C845 VTAIL.n6 VSUBS 2.33435f
C846 VTAIL.t1 VSUBS 0.249f
C847 VTAIL.t5 VSUBS 0.249f
C848 VTAIL.n7 VSUBS 1.77338f
C849 VTAIL.n8 VSUBS 2.33434f
C850 VTAIL.t9 VSUBS 0.249f
C851 VTAIL.t3 VSUBS 0.249f
C852 VTAIL.n9 VSUBS 1.77338f
C853 VTAIL.n10 VSUBS 0.925044f
C854 VTAIL.t4 VSUBS 2.34878f
C855 VTAIL.n11 VSUBS 0.997933f
C856 VTAIL.t15 VSUBS 0.249f
C857 VTAIL.t10 VSUBS 0.249f
C858 VTAIL.n12 VSUBS 1.77338f
C859 VTAIL.n13 VSUBS 0.894236f
C860 VTAIL.t18 VSUBS 0.249f
C861 VTAIL.t12 VSUBS 0.249f
C862 VTAIL.n14 VSUBS 1.77338f
C863 VTAIL.n15 VSUBS 0.925044f
C864 VTAIL.t13 VSUBS 2.34876f
C865 VTAIL.n16 VSUBS 2.29033f
C866 VTAIL.t0 VSUBS 2.34876f
C867 VTAIL.n17 VSUBS 2.29033f
C868 VTAIL.t6 VSUBS 0.249f
C869 VTAIL.t7 VSUBS 0.249f
C870 VTAIL.n18 VSUBS 1.77338f
C871 VTAIL.n19 VSUBS 0.808928f
C872 VP.n0 VSUBS 0.03854f
C873 VP.t1 VSUBS 1.78752f
C874 VP.n1 VSUBS 0.061889f
C875 VP.n2 VSUBS 0.03854f
C876 VP.t3 VSUBS 1.78752f
C877 VP.n3 VSUBS 0.072811f
C878 VP.n4 VSUBS 0.03854f
C879 VP.t7 VSUBS 1.78752f
C880 VP.n5 VSUBS 0.068279f
C881 VP.n6 VSUBS 0.03854f
C882 VP.n7 VSUBS 0.053122f
C883 VP.n8 VSUBS 0.03854f
C884 VP.t5 VSUBS 1.78752f
C885 VP.n9 VSUBS 0.061889f
C886 VP.n10 VSUBS 0.03854f
C887 VP.t4 VSUBS 1.78752f
C888 VP.n11 VSUBS 0.072811f
C889 VP.n12 VSUBS 0.03854f
C890 VP.t0 VSUBS 1.78752f
C891 VP.n13 VSUBS 0.068279f
C892 VP.t8 VSUBS 1.92143f
C893 VP.t2 VSUBS 1.78752f
C894 VP.n14 VSUBS 0.730824f
C895 VP.n15 VSUBS 0.733787f
C896 VP.n16 VSUBS 0.246041f
C897 VP.n17 VSUBS 0.03854f
C898 VP.n18 VSUBS 0.033255f
C899 VP.n19 VSUBS 0.072811f
C900 VP.n20 VSUBS 0.68579f
C901 VP.n21 VSUBS 0.03854f
C902 VP.n22 VSUBS 0.03854f
C903 VP.n23 VSUBS 0.03854f
C904 VP.n24 VSUBS 0.033255f
C905 VP.n25 VSUBS 0.068279f
C906 VP.n26 VSUBS 0.649603f
C907 VP.n27 VSUBS 0.04536f
C908 VP.n28 VSUBS 0.03854f
C909 VP.n29 VSUBS 0.03854f
C910 VP.n30 VSUBS 0.03854f
C911 VP.n31 VSUBS 0.05016f
C912 VP.n32 VSUBS 0.053122f
C913 VP.n33 VSUBS 0.734129f
C914 VP.n34 VSUBS 1.8888f
C915 VP.t9 VSUBS 1.78752f
C916 VP.n35 VSUBS 0.734129f
C917 VP.n36 VSUBS 1.91861f
C918 VP.n37 VSUBS 0.03854f
C919 VP.n38 VSUBS 0.03854f
C920 VP.n39 VSUBS 0.05016f
C921 VP.n40 VSUBS 0.061889f
C922 VP.t6 VSUBS 1.78752f
C923 VP.n41 VSUBS 0.649603f
C924 VP.n42 VSUBS 0.04536f
C925 VP.n43 VSUBS 0.03854f
C926 VP.n44 VSUBS 0.03854f
C927 VP.n45 VSUBS 0.03854f
C928 VP.n46 VSUBS 0.033255f
C929 VP.n47 VSUBS 0.072811f
C930 VP.n48 VSUBS 0.68579f
C931 VP.n49 VSUBS 0.03854f
C932 VP.n50 VSUBS 0.03854f
C933 VP.n51 VSUBS 0.03854f
C934 VP.n52 VSUBS 0.033255f
C935 VP.n53 VSUBS 0.068279f
C936 VP.n54 VSUBS 0.649603f
C937 VP.n55 VSUBS 0.04536f
C938 VP.n56 VSUBS 0.03854f
C939 VP.n57 VSUBS 0.03854f
C940 VP.n58 VSUBS 0.03854f
C941 VP.n59 VSUBS 0.05016f
C942 VP.n60 VSUBS 0.053122f
C943 VP.n61 VSUBS 0.734129f
C944 VP.n62 VSUBS 0.036568f
.ends

