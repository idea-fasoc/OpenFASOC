* NGSPICE file created from diff_pair_sample_1318.ext - technology: sky130A

.subckt diff_pair_sample_1318 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=2.58
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=2.58
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=2.58
X3 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=2.58
X4 VTAIL.t7 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=2.58
X5 VDD2.t3 VN.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=2.58
X6 VDD2.t2 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=2.58
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=2.58
X8 VTAIL.t5 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=2.58
X9 VTAIL.t9 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=2.58
X10 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=2.58
X11 VTAIL.t0 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=2.58
X12 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=2.58
X13 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=2.58
X14 VDD2.t0 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=2.58
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=2.58
R0 VN.n29 VN.n16 161.3
R1 VN.n28 VN.n27 161.3
R2 VN.n26 VN.n17 161.3
R3 VN.n25 VN.n24 161.3
R4 VN.n23 VN.n18 161.3
R5 VN.n22 VN.n21 161.3
R6 VN.n13 VN.n0 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n10 VN.n1 161.3
R9 VN.n9 VN.n8 161.3
R10 VN.n7 VN.n2 161.3
R11 VN.n6 VN.n5 161.3
R12 VN.n4 VN.t0 107.779
R13 VN.n20 VN.t3 107.779
R14 VN.n15 VN.n14 103.038
R15 VN.n31 VN.n30 103.038
R16 VN.n3 VN.t1 74.7292
R17 VN.n14 VN.t2 74.7292
R18 VN.n19 VN.t4 74.7292
R19 VN.n30 VN.t5 74.7292
R20 VN.n4 VN.n3 60.2499
R21 VN.n20 VN.n19 60.2499
R22 VN.n8 VN.n1 56.5617
R23 VN.n24 VN.n17 56.5617
R24 VN VN.n31 45.8277
R25 VN.n7 VN.n6 24.5923
R26 VN.n8 VN.n7 24.5923
R27 VN.n12 VN.n1 24.5923
R28 VN.n13 VN.n12 24.5923
R29 VN.n24 VN.n23 24.5923
R30 VN.n23 VN.n22 24.5923
R31 VN.n29 VN.n28 24.5923
R32 VN.n28 VN.n17 24.5923
R33 VN.n6 VN.n3 12.2964
R34 VN.n22 VN.n19 12.2964
R35 VN.n14 VN.n13 7.86989
R36 VN.n30 VN.n29 7.86989
R37 VN.n21 VN.n20 6.96699
R38 VN.n5 VN.n4 6.96699
R39 VN.n31 VN.n16 0.278335
R40 VN.n15 VN.n0 0.278335
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153485
R52 VTAIL.n170 VTAIL.n134 289.615
R53 VTAIL.n38 VTAIL.n2 289.615
R54 VTAIL.n128 VTAIL.n92 289.615
R55 VTAIL.n84 VTAIL.n48 289.615
R56 VTAIL.n146 VTAIL.n145 185
R57 VTAIL.n151 VTAIL.n150 185
R58 VTAIL.n153 VTAIL.n152 185
R59 VTAIL.n142 VTAIL.n141 185
R60 VTAIL.n159 VTAIL.n158 185
R61 VTAIL.n161 VTAIL.n160 185
R62 VTAIL.n138 VTAIL.n137 185
R63 VTAIL.n168 VTAIL.n167 185
R64 VTAIL.n169 VTAIL.n136 185
R65 VTAIL.n171 VTAIL.n170 185
R66 VTAIL.n14 VTAIL.n13 185
R67 VTAIL.n19 VTAIL.n18 185
R68 VTAIL.n21 VTAIL.n20 185
R69 VTAIL.n10 VTAIL.n9 185
R70 VTAIL.n27 VTAIL.n26 185
R71 VTAIL.n29 VTAIL.n28 185
R72 VTAIL.n6 VTAIL.n5 185
R73 VTAIL.n36 VTAIL.n35 185
R74 VTAIL.n37 VTAIL.n4 185
R75 VTAIL.n39 VTAIL.n38 185
R76 VTAIL.n129 VTAIL.n128 185
R77 VTAIL.n127 VTAIL.n94 185
R78 VTAIL.n126 VTAIL.n125 185
R79 VTAIL.n97 VTAIL.n95 185
R80 VTAIL.n120 VTAIL.n119 185
R81 VTAIL.n118 VTAIL.n117 185
R82 VTAIL.n101 VTAIL.n100 185
R83 VTAIL.n112 VTAIL.n111 185
R84 VTAIL.n110 VTAIL.n109 185
R85 VTAIL.n105 VTAIL.n104 185
R86 VTAIL.n85 VTAIL.n84 185
R87 VTAIL.n83 VTAIL.n50 185
R88 VTAIL.n82 VTAIL.n81 185
R89 VTAIL.n53 VTAIL.n51 185
R90 VTAIL.n76 VTAIL.n75 185
R91 VTAIL.n74 VTAIL.n73 185
R92 VTAIL.n57 VTAIL.n56 185
R93 VTAIL.n68 VTAIL.n67 185
R94 VTAIL.n66 VTAIL.n65 185
R95 VTAIL.n61 VTAIL.n60 185
R96 VTAIL.n147 VTAIL.t11 149.524
R97 VTAIL.n15 VTAIL.t2 149.524
R98 VTAIL.n106 VTAIL.t3 149.524
R99 VTAIL.n62 VTAIL.t8 149.524
R100 VTAIL.n151 VTAIL.n145 104.615
R101 VTAIL.n152 VTAIL.n151 104.615
R102 VTAIL.n152 VTAIL.n141 104.615
R103 VTAIL.n159 VTAIL.n141 104.615
R104 VTAIL.n160 VTAIL.n159 104.615
R105 VTAIL.n160 VTAIL.n137 104.615
R106 VTAIL.n168 VTAIL.n137 104.615
R107 VTAIL.n169 VTAIL.n168 104.615
R108 VTAIL.n170 VTAIL.n169 104.615
R109 VTAIL.n19 VTAIL.n13 104.615
R110 VTAIL.n20 VTAIL.n19 104.615
R111 VTAIL.n20 VTAIL.n9 104.615
R112 VTAIL.n27 VTAIL.n9 104.615
R113 VTAIL.n28 VTAIL.n27 104.615
R114 VTAIL.n28 VTAIL.n5 104.615
R115 VTAIL.n36 VTAIL.n5 104.615
R116 VTAIL.n37 VTAIL.n36 104.615
R117 VTAIL.n38 VTAIL.n37 104.615
R118 VTAIL.n128 VTAIL.n127 104.615
R119 VTAIL.n127 VTAIL.n126 104.615
R120 VTAIL.n126 VTAIL.n95 104.615
R121 VTAIL.n119 VTAIL.n95 104.615
R122 VTAIL.n119 VTAIL.n118 104.615
R123 VTAIL.n118 VTAIL.n100 104.615
R124 VTAIL.n111 VTAIL.n100 104.615
R125 VTAIL.n111 VTAIL.n110 104.615
R126 VTAIL.n110 VTAIL.n104 104.615
R127 VTAIL.n84 VTAIL.n83 104.615
R128 VTAIL.n83 VTAIL.n82 104.615
R129 VTAIL.n82 VTAIL.n51 104.615
R130 VTAIL.n75 VTAIL.n51 104.615
R131 VTAIL.n75 VTAIL.n74 104.615
R132 VTAIL.n74 VTAIL.n56 104.615
R133 VTAIL.n67 VTAIL.n56 104.615
R134 VTAIL.n67 VTAIL.n66 104.615
R135 VTAIL.n66 VTAIL.n60 104.615
R136 VTAIL.t11 VTAIL.n145 52.3082
R137 VTAIL.t2 VTAIL.n13 52.3082
R138 VTAIL.t3 VTAIL.n104 52.3082
R139 VTAIL.t8 VTAIL.n60 52.3082
R140 VTAIL.n91 VTAIL.n90 51.178
R141 VTAIL.n47 VTAIL.n46 51.178
R142 VTAIL.n1 VTAIL.n0 51.1778
R143 VTAIL.n45 VTAIL.n44 51.1778
R144 VTAIL.n175 VTAIL.n174 36.0641
R145 VTAIL.n43 VTAIL.n42 36.0641
R146 VTAIL.n133 VTAIL.n132 36.0641
R147 VTAIL.n89 VTAIL.n88 36.0641
R148 VTAIL.n47 VTAIL.n45 24.2807
R149 VTAIL.n175 VTAIL.n133 21.7721
R150 VTAIL.n171 VTAIL.n136 13.1884
R151 VTAIL.n39 VTAIL.n4 13.1884
R152 VTAIL.n129 VTAIL.n94 13.1884
R153 VTAIL.n85 VTAIL.n50 13.1884
R154 VTAIL.n167 VTAIL.n166 12.8005
R155 VTAIL.n172 VTAIL.n134 12.8005
R156 VTAIL.n35 VTAIL.n34 12.8005
R157 VTAIL.n40 VTAIL.n2 12.8005
R158 VTAIL.n130 VTAIL.n92 12.8005
R159 VTAIL.n125 VTAIL.n96 12.8005
R160 VTAIL.n86 VTAIL.n48 12.8005
R161 VTAIL.n81 VTAIL.n52 12.8005
R162 VTAIL.n165 VTAIL.n138 12.0247
R163 VTAIL.n33 VTAIL.n6 12.0247
R164 VTAIL.n124 VTAIL.n97 12.0247
R165 VTAIL.n80 VTAIL.n53 12.0247
R166 VTAIL.n162 VTAIL.n161 11.249
R167 VTAIL.n30 VTAIL.n29 11.249
R168 VTAIL.n121 VTAIL.n120 11.249
R169 VTAIL.n77 VTAIL.n76 11.249
R170 VTAIL.n158 VTAIL.n140 10.4732
R171 VTAIL.n26 VTAIL.n8 10.4732
R172 VTAIL.n117 VTAIL.n99 10.4732
R173 VTAIL.n73 VTAIL.n55 10.4732
R174 VTAIL.n147 VTAIL.n146 10.2747
R175 VTAIL.n15 VTAIL.n14 10.2747
R176 VTAIL.n106 VTAIL.n105 10.2747
R177 VTAIL.n62 VTAIL.n61 10.2747
R178 VTAIL.n157 VTAIL.n142 9.69747
R179 VTAIL.n25 VTAIL.n10 9.69747
R180 VTAIL.n116 VTAIL.n101 9.69747
R181 VTAIL.n72 VTAIL.n57 9.69747
R182 VTAIL.n174 VTAIL.n173 9.45567
R183 VTAIL.n42 VTAIL.n41 9.45567
R184 VTAIL.n132 VTAIL.n131 9.45567
R185 VTAIL.n88 VTAIL.n87 9.45567
R186 VTAIL.n173 VTAIL.n172 9.3005
R187 VTAIL.n149 VTAIL.n148 9.3005
R188 VTAIL.n144 VTAIL.n143 9.3005
R189 VTAIL.n155 VTAIL.n154 9.3005
R190 VTAIL.n157 VTAIL.n156 9.3005
R191 VTAIL.n140 VTAIL.n139 9.3005
R192 VTAIL.n163 VTAIL.n162 9.3005
R193 VTAIL.n165 VTAIL.n164 9.3005
R194 VTAIL.n166 VTAIL.n135 9.3005
R195 VTAIL.n41 VTAIL.n40 9.3005
R196 VTAIL.n17 VTAIL.n16 9.3005
R197 VTAIL.n12 VTAIL.n11 9.3005
R198 VTAIL.n23 VTAIL.n22 9.3005
R199 VTAIL.n25 VTAIL.n24 9.3005
R200 VTAIL.n8 VTAIL.n7 9.3005
R201 VTAIL.n31 VTAIL.n30 9.3005
R202 VTAIL.n33 VTAIL.n32 9.3005
R203 VTAIL.n34 VTAIL.n3 9.3005
R204 VTAIL.n108 VTAIL.n107 9.3005
R205 VTAIL.n103 VTAIL.n102 9.3005
R206 VTAIL.n114 VTAIL.n113 9.3005
R207 VTAIL.n116 VTAIL.n115 9.3005
R208 VTAIL.n99 VTAIL.n98 9.3005
R209 VTAIL.n122 VTAIL.n121 9.3005
R210 VTAIL.n124 VTAIL.n123 9.3005
R211 VTAIL.n96 VTAIL.n93 9.3005
R212 VTAIL.n131 VTAIL.n130 9.3005
R213 VTAIL.n64 VTAIL.n63 9.3005
R214 VTAIL.n59 VTAIL.n58 9.3005
R215 VTAIL.n70 VTAIL.n69 9.3005
R216 VTAIL.n72 VTAIL.n71 9.3005
R217 VTAIL.n55 VTAIL.n54 9.3005
R218 VTAIL.n78 VTAIL.n77 9.3005
R219 VTAIL.n80 VTAIL.n79 9.3005
R220 VTAIL.n52 VTAIL.n49 9.3005
R221 VTAIL.n87 VTAIL.n86 9.3005
R222 VTAIL.n154 VTAIL.n153 8.92171
R223 VTAIL.n22 VTAIL.n21 8.92171
R224 VTAIL.n113 VTAIL.n112 8.92171
R225 VTAIL.n69 VTAIL.n68 8.92171
R226 VTAIL.n150 VTAIL.n144 8.14595
R227 VTAIL.n18 VTAIL.n12 8.14595
R228 VTAIL.n109 VTAIL.n103 8.14595
R229 VTAIL.n65 VTAIL.n59 8.14595
R230 VTAIL.n149 VTAIL.n146 7.3702
R231 VTAIL.n17 VTAIL.n14 7.3702
R232 VTAIL.n108 VTAIL.n105 7.3702
R233 VTAIL.n64 VTAIL.n61 7.3702
R234 VTAIL.n150 VTAIL.n149 5.81868
R235 VTAIL.n18 VTAIL.n17 5.81868
R236 VTAIL.n109 VTAIL.n108 5.81868
R237 VTAIL.n65 VTAIL.n64 5.81868
R238 VTAIL.n153 VTAIL.n144 5.04292
R239 VTAIL.n21 VTAIL.n12 5.04292
R240 VTAIL.n112 VTAIL.n103 5.04292
R241 VTAIL.n68 VTAIL.n59 5.04292
R242 VTAIL.n154 VTAIL.n142 4.26717
R243 VTAIL.n22 VTAIL.n10 4.26717
R244 VTAIL.n113 VTAIL.n101 4.26717
R245 VTAIL.n69 VTAIL.n57 4.26717
R246 VTAIL.n158 VTAIL.n157 3.49141
R247 VTAIL.n26 VTAIL.n25 3.49141
R248 VTAIL.n117 VTAIL.n116 3.49141
R249 VTAIL.n73 VTAIL.n72 3.49141
R250 VTAIL.n148 VTAIL.n147 2.84304
R251 VTAIL.n16 VTAIL.n15 2.84304
R252 VTAIL.n107 VTAIL.n106 2.84304
R253 VTAIL.n63 VTAIL.n62 2.84304
R254 VTAIL.n161 VTAIL.n140 2.71565
R255 VTAIL.n29 VTAIL.n8 2.71565
R256 VTAIL.n120 VTAIL.n99 2.71565
R257 VTAIL.n76 VTAIL.n55 2.71565
R258 VTAIL.n89 VTAIL.n47 2.50912
R259 VTAIL.n133 VTAIL.n91 2.50912
R260 VTAIL.n45 VTAIL.n43 2.50912
R261 VTAIL.n0 VTAIL.t6 2.4755
R262 VTAIL.n0 VTAIL.t7 2.4755
R263 VTAIL.n44 VTAIL.t4 2.4755
R264 VTAIL.n44 VTAIL.t5 2.4755
R265 VTAIL.n90 VTAIL.t1 2.4755
R266 VTAIL.n90 VTAIL.t0 2.4755
R267 VTAIL.n46 VTAIL.t10 2.4755
R268 VTAIL.n46 VTAIL.t9 2.4755
R269 VTAIL.n162 VTAIL.n138 1.93989
R270 VTAIL.n30 VTAIL.n6 1.93989
R271 VTAIL.n121 VTAIL.n97 1.93989
R272 VTAIL.n77 VTAIL.n53 1.93989
R273 VTAIL VTAIL.n175 1.82378
R274 VTAIL.n91 VTAIL.n89 1.72464
R275 VTAIL.n43 VTAIL.n1 1.72464
R276 VTAIL.n167 VTAIL.n165 1.16414
R277 VTAIL.n174 VTAIL.n134 1.16414
R278 VTAIL.n35 VTAIL.n33 1.16414
R279 VTAIL.n42 VTAIL.n2 1.16414
R280 VTAIL.n132 VTAIL.n92 1.16414
R281 VTAIL.n125 VTAIL.n124 1.16414
R282 VTAIL.n88 VTAIL.n48 1.16414
R283 VTAIL.n81 VTAIL.n80 1.16414
R284 VTAIL VTAIL.n1 0.685845
R285 VTAIL.n166 VTAIL.n136 0.388379
R286 VTAIL.n172 VTAIL.n171 0.388379
R287 VTAIL.n34 VTAIL.n4 0.388379
R288 VTAIL.n40 VTAIL.n39 0.388379
R289 VTAIL.n130 VTAIL.n129 0.388379
R290 VTAIL.n96 VTAIL.n94 0.388379
R291 VTAIL.n86 VTAIL.n85 0.388379
R292 VTAIL.n52 VTAIL.n50 0.388379
R293 VTAIL.n148 VTAIL.n143 0.155672
R294 VTAIL.n155 VTAIL.n143 0.155672
R295 VTAIL.n156 VTAIL.n155 0.155672
R296 VTAIL.n156 VTAIL.n139 0.155672
R297 VTAIL.n163 VTAIL.n139 0.155672
R298 VTAIL.n164 VTAIL.n163 0.155672
R299 VTAIL.n164 VTAIL.n135 0.155672
R300 VTAIL.n173 VTAIL.n135 0.155672
R301 VTAIL.n16 VTAIL.n11 0.155672
R302 VTAIL.n23 VTAIL.n11 0.155672
R303 VTAIL.n24 VTAIL.n23 0.155672
R304 VTAIL.n24 VTAIL.n7 0.155672
R305 VTAIL.n31 VTAIL.n7 0.155672
R306 VTAIL.n32 VTAIL.n31 0.155672
R307 VTAIL.n32 VTAIL.n3 0.155672
R308 VTAIL.n41 VTAIL.n3 0.155672
R309 VTAIL.n131 VTAIL.n93 0.155672
R310 VTAIL.n123 VTAIL.n93 0.155672
R311 VTAIL.n123 VTAIL.n122 0.155672
R312 VTAIL.n122 VTAIL.n98 0.155672
R313 VTAIL.n115 VTAIL.n98 0.155672
R314 VTAIL.n115 VTAIL.n114 0.155672
R315 VTAIL.n114 VTAIL.n102 0.155672
R316 VTAIL.n107 VTAIL.n102 0.155672
R317 VTAIL.n87 VTAIL.n49 0.155672
R318 VTAIL.n79 VTAIL.n49 0.155672
R319 VTAIL.n79 VTAIL.n78 0.155672
R320 VTAIL.n78 VTAIL.n54 0.155672
R321 VTAIL.n71 VTAIL.n54 0.155672
R322 VTAIL.n71 VTAIL.n70 0.155672
R323 VTAIL.n70 VTAIL.n58 0.155672
R324 VTAIL.n63 VTAIL.n58 0.155672
R325 VDD2.n79 VDD2.n43 289.615
R326 VDD2.n36 VDD2.n0 289.615
R327 VDD2.n80 VDD2.n79 185
R328 VDD2.n78 VDD2.n45 185
R329 VDD2.n77 VDD2.n76 185
R330 VDD2.n48 VDD2.n46 185
R331 VDD2.n71 VDD2.n70 185
R332 VDD2.n69 VDD2.n68 185
R333 VDD2.n52 VDD2.n51 185
R334 VDD2.n63 VDD2.n62 185
R335 VDD2.n61 VDD2.n60 185
R336 VDD2.n56 VDD2.n55 185
R337 VDD2.n12 VDD2.n11 185
R338 VDD2.n17 VDD2.n16 185
R339 VDD2.n19 VDD2.n18 185
R340 VDD2.n8 VDD2.n7 185
R341 VDD2.n25 VDD2.n24 185
R342 VDD2.n27 VDD2.n26 185
R343 VDD2.n4 VDD2.n3 185
R344 VDD2.n34 VDD2.n33 185
R345 VDD2.n35 VDD2.n2 185
R346 VDD2.n37 VDD2.n36 185
R347 VDD2.n57 VDD2.t0 149.524
R348 VDD2.n13 VDD2.t5 149.524
R349 VDD2.n79 VDD2.n78 104.615
R350 VDD2.n78 VDD2.n77 104.615
R351 VDD2.n77 VDD2.n46 104.615
R352 VDD2.n70 VDD2.n46 104.615
R353 VDD2.n70 VDD2.n69 104.615
R354 VDD2.n69 VDD2.n51 104.615
R355 VDD2.n62 VDD2.n51 104.615
R356 VDD2.n62 VDD2.n61 104.615
R357 VDD2.n61 VDD2.n55 104.615
R358 VDD2.n17 VDD2.n11 104.615
R359 VDD2.n18 VDD2.n17 104.615
R360 VDD2.n18 VDD2.n7 104.615
R361 VDD2.n25 VDD2.n7 104.615
R362 VDD2.n26 VDD2.n25 104.615
R363 VDD2.n26 VDD2.n3 104.615
R364 VDD2.n34 VDD2.n3 104.615
R365 VDD2.n35 VDD2.n34 104.615
R366 VDD2.n36 VDD2.n35 104.615
R367 VDD2.n42 VDD2.n41 68.4284
R368 VDD2 VDD2.n85 68.4256
R369 VDD2.n42 VDD2.n40 54.569
R370 VDD2.n84 VDD2.n83 52.7429
R371 VDD2.t0 VDD2.n55 52.3082
R372 VDD2.t5 VDD2.n11 52.3082
R373 VDD2.n84 VDD2.n42 38.7649
R374 VDD2.n80 VDD2.n45 13.1884
R375 VDD2.n37 VDD2.n2 13.1884
R376 VDD2.n81 VDD2.n43 12.8005
R377 VDD2.n76 VDD2.n47 12.8005
R378 VDD2.n33 VDD2.n32 12.8005
R379 VDD2.n38 VDD2.n0 12.8005
R380 VDD2.n75 VDD2.n48 12.0247
R381 VDD2.n31 VDD2.n4 12.0247
R382 VDD2.n72 VDD2.n71 11.249
R383 VDD2.n28 VDD2.n27 11.249
R384 VDD2.n68 VDD2.n50 10.4732
R385 VDD2.n24 VDD2.n6 10.4732
R386 VDD2.n57 VDD2.n56 10.2747
R387 VDD2.n13 VDD2.n12 10.2747
R388 VDD2.n67 VDD2.n52 9.69747
R389 VDD2.n23 VDD2.n8 9.69747
R390 VDD2.n83 VDD2.n82 9.45567
R391 VDD2.n40 VDD2.n39 9.45567
R392 VDD2.n59 VDD2.n58 9.3005
R393 VDD2.n54 VDD2.n53 9.3005
R394 VDD2.n65 VDD2.n64 9.3005
R395 VDD2.n67 VDD2.n66 9.3005
R396 VDD2.n50 VDD2.n49 9.3005
R397 VDD2.n73 VDD2.n72 9.3005
R398 VDD2.n75 VDD2.n74 9.3005
R399 VDD2.n47 VDD2.n44 9.3005
R400 VDD2.n82 VDD2.n81 9.3005
R401 VDD2.n39 VDD2.n38 9.3005
R402 VDD2.n15 VDD2.n14 9.3005
R403 VDD2.n10 VDD2.n9 9.3005
R404 VDD2.n21 VDD2.n20 9.3005
R405 VDD2.n23 VDD2.n22 9.3005
R406 VDD2.n6 VDD2.n5 9.3005
R407 VDD2.n29 VDD2.n28 9.3005
R408 VDD2.n31 VDD2.n30 9.3005
R409 VDD2.n32 VDD2.n1 9.3005
R410 VDD2.n64 VDD2.n63 8.92171
R411 VDD2.n20 VDD2.n19 8.92171
R412 VDD2.n60 VDD2.n54 8.14595
R413 VDD2.n16 VDD2.n10 8.14595
R414 VDD2.n59 VDD2.n56 7.3702
R415 VDD2.n15 VDD2.n12 7.3702
R416 VDD2.n60 VDD2.n59 5.81868
R417 VDD2.n16 VDD2.n15 5.81868
R418 VDD2.n63 VDD2.n54 5.04292
R419 VDD2.n19 VDD2.n10 5.04292
R420 VDD2.n64 VDD2.n52 4.26717
R421 VDD2.n20 VDD2.n8 4.26717
R422 VDD2.n68 VDD2.n67 3.49141
R423 VDD2.n24 VDD2.n23 3.49141
R424 VDD2.n58 VDD2.n57 2.84304
R425 VDD2.n14 VDD2.n13 2.84304
R426 VDD2.n71 VDD2.n50 2.71565
R427 VDD2.n27 VDD2.n6 2.71565
R428 VDD2.n85 VDD2.t1 2.4755
R429 VDD2.n85 VDD2.t2 2.4755
R430 VDD2.n41 VDD2.t4 2.4755
R431 VDD2.n41 VDD2.t3 2.4755
R432 VDD2 VDD2.n84 1.94016
R433 VDD2.n72 VDD2.n48 1.93989
R434 VDD2.n28 VDD2.n4 1.93989
R435 VDD2.n83 VDD2.n43 1.16414
R436 VDD2.n76 VDD2.n75 1.16414
R437 VDD2.n33 VDD2.n31 1.16414
R438 VDD2.n40 VDD2.n0 1.16414
R439 VDD2.n81 VDD2.n80 0.388379
R440 VDD2.n47 VDD2.n45 0.388379
R441 VDD2.n32 VDD2.n2 0.388379
R442 VDD2.n38 VDD2.n37 0.388379
R443 VDD2.n82 VDD2.n44 0.155672
R444 VDD2.n74 VDD2.n44 0.155672
R445 VDD2.n74 VDD2.n73 0.155672
R446 VDD2.n73 VDD2.n49 0.155672
R447 VDD2.n66 VDD2.n49 0.155672
R448 VDD2.n66 VDD2.n65 0.155672
R449 VDD2.n65 VDD2.n53 0.155672
R450 VDD2.n58 VDD2.n53 0.155672
R451 VDD2.n14 VDD2.n9 0.155672
R452 VDD2.n21 VDD2.n9 0.155672
R453 VDD2.n22 VDD2.n21 0.155672
R454 VDD2.n22 VDD2.n5 0.155672
R455 VDD2.n29 VDD2.n5 0.155672
R456 VDD2.n30 VDD2.n29 0.155672
R457 VDD2.n30 VDD2.n1 0.155672
R458 VDD2.n39 VDD2.n1 0.155672
R459 B.n561 B.n560 585
R460 B.n561 B.n79 585
R461 B.n564 B.n563 585
R462 B.n565 B.n118 585
R463 B.n567 B.n566 585
R464 B.n569 B.n117 585
R465 B.n572 B.n571 585
R466 B.n573 B.n116 585
R467 B.n575 B.n574 585
R468 B.n577 B.n115 585
R469 B.n580 B.n579 585
R470 B.n581 B.n114 585
R471 B.n583 B.n582 585
R472 B.n585 B.n113 585
R473 B.n588 B.n587 585
R474 B.n589 B.n112 585
R475 B.n591 B.n590 585
R476 B.n593 B.n111 585
R477 B.n596 B.n595 585
R478 B.n597 B.n110 585
R479 B.n599 B.n598 585
R480 B.n601 B.n109 585
R481 B.n604 B.n603 585
R482 B.n605 B.n108 585
R483 B.n607 B.n606 585
R484 B.n609 B.n107 585
R485 B.n612 B.n611 585
R486 B.n613 B.n106 585
R487 B.n615 B.n614 585
R488 B.n617 B.n105 585
R489 B.n620 B.n619 585
R490 B.n622 B.n102 585
R491 B.n624 B.n623 585
R492 B.n626 B.n101 585
R493 B.n629 B.n628 585
R494 B.n630 B.n100 585
R495 B.n632 B.n631 585
R496 B.n634 B.n99 585
R497 B.n636 B.n635 585
R498 B.n638 B.n637 585
R499 B.n641 B.n640 585
R500 B.n642 B.n94 585
R501 B.n644 B.n643 585
R502 B.n646 B.n93 585
R503 B.n649 B.n648 585
R504 B.n650 B.n92 585
R505 B.n652 B.n651 585
R506 B.n654 B.n91 585
R507 B.n657 B.n656 585
R508 B.n658 B.n90 585
R509 B.n660 B.n659 585
R510 B.n662 B.n89 585
R511 B.n665 B.n664 585
R512 B.n666 B.n88 585
R513 B.n668 B.n667 585
R514 B.n670 B.n87 585
R515 B.n673 B.n672 585
R516 B.n674 B.n86 585
R517 B.n676 B.n675 585
R518 B.n678 B.n85 585
R519 B.n681 B.n680 585
R520 B.n682 B.n84 585
R521 B.n684 B.n683 585
R522 B.n686 B.n83 585
R523 B.n689 B.n688 585
R524 B.n690 B.n82 585
R525 B.n692 B.n691 585
R526 B.n694 B.n81 585
R527 B.n697 B.n696 585
R528 B.n698 B.n80 585
R529 B.n559 B.n78 585
R530 B.n701 B.n78 585
R531 B.n558 B.n77 585
R532 B.n702 B.n77 585
R533 B.n557 B.n76 585
R534 B.n703 B.n76 585
R535 B.n556 B.n555 585
R536 B.n555 B.n72 585
R537 B.n554 B.n71 585
R538 B.n709 B.n71 585
R539 B.n553 B.n70 585
R540 B.n710 B.n70 585
R541 B.n552 B.n69 585
R542 B.n711 B.n69 585
R543 B.n551 B.n550 585
R544 B.n550 B.n68 585
R545 B.n549 B.n64 585
R546 B.n717 B.n64 585
R547 B.n548 B.n63 585
R548 B.n718 B.n63 585
R549 B.n547 B.n62 585
R550 B.n719 B.n62 585
R551 B.n546 B.n545 585
R552 B.n545 B.n58 585
R553 B.n544 B.n57 585
R554 B.n725 B.n57 585
R555 B.n543 B.n56 585
R556 B.n726 B.n56 585
R557 B.n542 B.n55 585
R558 B.n727 B.n55 585
R559 B.n541 B.n540 585
R560 B.n540 B.n51 585
R561 B.n539 B.n50 585
R562 B.n733 B.n50 585
R563 B.n538 B.n49 585
R564 B.n734 B.n49 585
R565 B.n537 B.n48 585
R566 B.n735 B.n48 585
R567 B.n536 B.n535 585
R568 B.n535 B.n47 585
R569 B.n534 B.n43 585
R570 B.n741 B.n43 585
R571 B.n533 B.n42 585
R572 B.n742 B.n42 585
R573 B.n532 B.n41 585
R574 B.n743 B.n41 585
R575 B.n531 B.n530 585
R576 B.n530 B.n37 585
R577 B.n529 B.n36 585
R578 B.n749 B.n36 585
R579 B.n528 B.n35 585
R580 B.n750 B.n35 585
R581 B.n527 B.n34 585
R582 B.n751 B.n34 585
R583 B.n526 B.n525 585
R584 B.n525 B.n30 585
R585 B.n524 B.n29 585
R586 B.n757 B.n29 585
R587 B.n523 B.n28 585
R588 B.n758 B.n28 585
R589 B.n522 B.n27 585
R590 B.n759 B.n27 585
R591 B.n521 B.n520 585
R592 B.n520 B.n23 585
R593 B.n519 B.n22 585
R594 B.n765 B.n22 585
R595 B.n518 B.n21 585
R596 B.n766 B.n21 585
R597 B.n517 B.n20 585
R598 B.n767 B.n20 585
R599 B.n516 B.n515 585
R600 B.n515 B.n16 585
R601 B.n514 B.n15 585
R602 B.n773 B.n15 585
R603 B.n513 B.n14 585
R604 B.n774 B.n14 585
R605 B.n512 B.n13 585
R606 B.n775 B.n13 585
R607 B.n511 B.n510 585
R608 B.n510 B.n12 585
R609 B.n509 B.n508 585
R610 B.n509 B.n8 585
R611 B.n507 B.n7 585
R612 B.n782 B.n7 585
R613 B.n506 B.n6 585
R614 B.n783 B.n6 585
R615 B.n505 B.n5 585
R616 B.n784 B.n5 585
R617 B.n504 B.n503 585
R618 B.n503 B.n4 585
R619 B.n502 B.n119 585
R620 B.n502 B.n501 585
R621 B.n492 B.n120 585
R622 B.n121 B.n120 585
R623 B.n494 B.n493 585
R624 B.n495 B.n494 585
R625 B.n491 B.n126 585
R626 B.n126 B.n125 585
R627 B.n490 B.n489 585
R628 B.n489 B.n488 585
R629 B.n128 B.n127 585
R630 B.n129 B.n128 585
R631 B.n481 B.n480 585
R632 B.n482 B.n481 585
R633 B.n479 B.n134 585
R634 B.n134 B.n133 585
R635 B.n478 B.n477 585
R636 B.n477 B.n476 585
R637 B.n136 B.n135 585
R638 B.n137 B.n136 585
R639 B.n469 B.n468 585
R640 B.n470 B.n469 585
R641 B.n467 B.n142 585
R642 B.n142 B.n141 585
R643 B.n466 B.n465 585
R644 B.n465 B.n464 585
R645 B.n144 B.n143 585
R646 B.n145 B.n144 585
R647 B.n457 B.n456 585
R648 B.n458 B.n457 585
R649 B.n455 B.n150 585
R650 B.n150 B.n149 585
R651 B.n454 B.n453 585
R652 B.n453 B.n452 585
R653 B.n152 B.n151 585
R654 B.n153 B.n152 585
R655 B.n445 B.n444 585
R656 B.n446 B.n445 585
R657 B.n443 B.n158 585
R658 B.n158 B.n157 585
R659 B.n442 B.n441 585
R660 B.n441 B.n440 585
R661 B.n160 B.n159 585
R662 B.n433 B.n160 585
R663 B.n432 B.n431 585
R664 B.n434 B.n432 585
R665 B.n430 B.n165 585
R666 B.n165 B.n164 585
R667 B.n429 B.n428 585
R668 B.n428 B.n427 585
R669 B.n167 B.n166 585
R670 B.n168 B.n167 585
R671 B.n420 B.n419 585
R672 B.n421 B.n420 585
R673 B.n418 B.n173 585
R674 B.n173 B.n172 585
R675 B.n417 B.n416 585
R676 B.n416 B.n415 585
R677 B.n175 B.n174 585
R678 B.n176 B.n175 585
R679 B.n408 B.n407 585
R680 B.n409 B.n408 585
R681 B.n406 B.n181 585
R682 B.n181 B.n180 585
R683 B.n405 B.n404 585
R684 B.n404 B.n403 585
R685 B.n183 B.n182 585
R686 B.n396 B.n183 585
R687 B.n395 B.n394 585
R688 B.n397 B.n395 585
R689 B.n393 B.n188 585
R690 B.n188 B.n187 585
R691 B.n392 B.n391 585
R692 B.n391 B.n390 585
R693 B.n190 B.n189 585
R694 B.n191 B.n190 585
R695 B.n383 B.n382 585
R696 B.n384 B.n383 585
R697 B.n381 B.n196 585
R698 B.n196 B.n195 585
R699 B.n380 B.n379 585
R700 B.n379 B.n378 585
R701 B.n375 B.n200 585
R702 B.n374 B.n373 585
R703 B.n371 B.n201 585
R704 B.n371 B.n199 585
R705 B.n370 B.n369 585
R706 B.n368 B.n367 585
R707 B.n366 B.n203 585
R708 B.n364 B.n363 585
R709 B.n362 B.n204 585
R710 B.n361 B.n360 585
R711 B.n358 B.n205 585
R712 B.n356 B.n355 585
R713 B.n354 B.n206 585
R714 B.n353 B.n352 585
R715 B.n350 B.n207 585
R716 B.n348 B.n347 585
R717 B.n346 B.n208 585
R718 B.n345 B.n344 585
R719 B.n342 B.n209 585
R720 B.n340 B.n339 585
R721 B.n338 B.n210 585
R722 B.n337 B.n336 585
R723 B.n334 B.n211 585
R724 B.n332 B.n331 585
R725 B.n330 B.n212 585
R726 B.n329 B.n328 585
R727 B.n326 B.n213 585
R728 B.n324 B.n323 585
R729 B.n322 B.n214 585
R730 B.n321 B.n320 585
R731 B.n318 B.n215 585
R732 B.n316 B.n315 585
R733 B.n314 B.n216 585
R734 B.n313 B.n312 585
R735 B.n310 B.n220 585
R736 B.n308 B.n307 585
R737 B.n306 B.n221 585
R738 B.n305 B.n304 585
R739 B.n302 B.n222 585
R740 B.n300 B.n299 585
R741 B.n297 B.n223 585
R742 B.n296 B.n295 585
R743 B.n293 B.n226 585
R744 B.n291 B.n290 585
R745 B.n289 B.n227 585
R746 B.n288 B.n287 585
R747 B.n285 B.n228 585
R748 B.n283 B.n282 585
R749 B.n281 B.n229 585
R750 B.n280 B.n279 585
R751 B.n277 B.n230 585
R752 B.n275 B.n274 585
R753 B.n273 B.n231 585
R754 B.n272 B.n271 585
R755 B.n269 B.n232 585
R756 B.n267 B.n266 585
R757 B.n265 B.n233 585
R758 B.n264 B.n263 585
R759 B.n261 B.n234 585
R760 B.n259 B.n258 585
R761 B.n257 B.n235 585
R762 B.n256 B.n255 585
R763 B.n253 B.n236 585
R764 B.n251 B.n250 585
R765 B.n249 B.n237 585
R766 B.n248 B.n247 585
R767 B.n245 B.n238 585
R768 B.n243 B.n242 585
R769 B.n241 B.n240 585
R770 B.n198 B.n197 585
R771 B.n377 B.n376 585
R772 B.n378 B.n377 585
R773 B.n194 B.n193 585
R774 B.n195 B.n194 585
R775 B.n386 B.n385 585
R776 B.n385 B.n384 585
R777 B.n387 B.n192 585
R778 B.n192 B.n191 585
R779 B.n389 B.n388 585
R780 B.n390 B.n389 585
R781 B.n186 B.n185 585
R782 B.n187 B.n186 585
R783 B.n399 B.n398 585
R784 B.n398 B.n397 585
R785 B.n400 B.n184 585
R786 B.n396 B.n184 585
R787 B.n402 B.n401 585
R788 B.n403 B.n402 585
R789 B.n179 B.n178 585
R790 B.n180 B.n179 585
R791 B.n411 B.n410 585
R792 B.n410 B.n409 585
R793 B.n412 B.n177 585
R794 B.n177 B.n176 585
R795 B.n414 B.n413 585
R796 B.n415 B.n414 585
R797 B.n171 B.n170 585
R798 B.n172 B.n171 585
R799 B.n423 B.n422 585
R800 B.n422 B.n421 585
R801 B.n424 B.n169 585
R802 B.n169 B.n168 585
R803 B.n426 B.n425 585
R804 B.n427 B.n426 585
R805 B.n163 B.n162 585
R806 B.n164 B.n163 585
R807 B.n436 B.n435 585
R808 B.n435 B.n434 585
R809 B.n437 B.n161 585
R810 B.n433 B.n161 585
R811 B.n439 B.n438 585
R812 B.n440 B.n439 585
R813 B.n156 B.n155 585
R814 B.n157 B.n156 585
R815 B.n448 B.n447 585
R816 B.n447 B.n446 585
R817 B.n449 B.n154 585
R818 B.n154 B.n153 585
R819 B.n451 B.n450 585
R820 B.n452 B.n451 585
R821 B.n148 B.n147 585
R822 B.n149 B.n148 585
R823 B.n460 B.n459 585
R824 B.n459 B.n458 585
R825 B.n461 B.n146 585
R826 B.n146 B.n145 585
R827 B.n463 B.n462 585
R828 B.n464 B.n463 585
R829 B.n140 B.n139 585
R830 B.n141 B.n140 585
R831 B.n472 B.n471 585
R832 B.n471 B.n470 585
R833 B.n473 B.n138 585
R834 B.n138 B.n137 585
R835 B.n475 B.n474 585
R836 B.n476 B.n475 585
R837 B.n132 B.n131 585
R838 B.n133 B.n132 585
R839 B.n484 B.n483 585
R840 B.n483 B.n482 585
R841 B.n485 B.n130 585
R842 B.n130 B.n129 585
R843 B.n487 B.n486 585
R844 B.n488 B.n487 585
R845 B.n124 B.n123 585
R846 B.n125 B.n124 585
R847 B.n497 B.n496 585
R848 B.n496 B.n495 585
R849 B.n498 B.n122 585
R850 B.n122 B.n121 585
R851 B.n500 B.n499 585
R852 B.n501 B.n500 585
R853 B.n3 B.n0 585
R854 B.n4 B.n3 585
R855 B.n781 B.n1 585
R856 B.n782 B.n781 585
R857 B.n780 B.n779 585
R858 B.n780 B.n8 585
R859 B.n778 B.n9 585
R860 B.n12 B.n9 585
R861 B.n777 B.n776 585
R862 B.n776 B.n775 585
R863 B.n11 B.n10 585
R864 B.n774 B.n11 585
R865 B.n772 B.n771 585
R866 B.n773 B.n772 585
R867 B.n770 B.n17 585
R868 B.n17 B.n16 585
R869 B.n769 B.n768 585
R870 B.n768 B.n767 585
R871 B.n19 B.n18 585
R872 B.n766 B.n19 585
R873 B.n764 B.n763 585
R874 B.n765 B.n764 585
R875 B.n762 B.n24 585
R876 B.n24 B.n23 585
R877 B.n761 B.n760 585
R878 B.n760 B.n759 585
R879 B.n26 B.n25 585
R880 B.n758 B.n26 585
R881 B.n756 B.n755 585
R882 B.n757 B.n756 585
R883 B.n754 B.n31 585
R884 B.n31 B.n30 585
R885 B.n753 B.n752 585
R886 B.n752 B.n751 585
R887 B.n33 B.n32 585
R888 B.n750 B.n33 585
R889 B.n748 B.n747 585
R890 B.n749 B.n748 585
R891 B.n746 B.n38 585
R892 B.n38 B.n37 585
R893 B.n745 B.n744 585
R894 B.n744 B.n743 585
R895 B.n40 B.n39 585
R896 B.n742 B.n40 585
R897 B.n740 B.n739 585
R898 B.n741 B.n740 585
R899 B.n738 B.n44 585
R900 B.n47 B.n44 585
R901 B.n737 B.n736 585
R902 B.n736 B.n735 585
R903 B.n46 B.n45 585
R904 B.n734 B.n46 585
R905 B.n732 B.n731 585
R906 B.n733 B.n732 585
R907 B.n730 B.n52 585
R908 B.n52 B.n51 585
R909 B.n729 B.n728 585
R910 B.n728 B.n727 585
R911 B.n54 B.n53 585
R912 B.n726 B.n54 585
R913 B.n724 B.n723 585
R914 B.n725 B.n724 585
R915 B.n722 B.n59 585
R916 B.n59 B.n58 585
R917 B.n721 B.n720 585
R918 B.n720 B.n719 585
R919 B.n61 B.n60 585
R920 B.n718 B.n61 585
R921 B.n716 B.n715 585
R922 B.n717 B.n716 585
R923 B.n714 B.n65 585
R924 B.n68 B.n65 585
R925 B.n713 B.n712 585
R926 B.n712 B.n711 585
R927 B.n67 B.n66 585
R928 B.n710 B.n67 585
R929 B.n708 B.n707 585
R930 B.n709 B.n708 585
R931 B.n706 B.n73 585
R932 B.n73 B.n72 585
R933 B.n705 B.n704 585
R934 B.n704 B.n703 585
R935 B.n75 B.n74 585
R936 B.n702 B.n75 585
R937 B.n700 B.n699 585
R938 B.n701 B.n700 585
R939 B.n785 B.n784 585
R940 B.n783 B.n2 585
R941 B.n700 B.n80 497.305
R942 B.n561 B.n78 497.305
R943 B.n379 B.n198 497.305
R944 B.n377 B.n200 497.305
R945 B.n95 B.t14 282.745
R946 B.n103 B.t10 282.745
R947 B.n224 B.t6 282.745
R948 B.n217 B.t17 282.745
R949 B.n103 B.t12 269.728
R950 B.n224 B.t9 269.728
R951 B.n95 B.t15 269.728
R952 B.n217 B.t19 269.728
R953 B.n562 B.n79 256.663
R954 B.n568 B.n79 256.663
R955 B.n570 B.n79 256.663
R956 B.n576 B.n79 256.663
R957 B.n578 B.n79 256.663
R958 B.n584 B.n79 256.663
R959 B.n586 B.n79 256.663
R960 B.n592 B.n79 256.663
R961 B.n594 B.n79 256.663
R962 B.n600 B.n79 256.663
R963 B.n602 B.n79 256.663
R964 B.n608 B.n79 256.663
R965 B.n610 B.n79 256.663
R966 B.n616 B.n79 256.663
R967 B.n618 B.n79 256.663
R968 B.n625 B.n79 256.663
R969 B.n627 B.n79 256.663
R970 B.n633 B.n79 256.663
R971 B.n98 B.n79 256.663
R972 B.n639 B.n79 256.663
R973 B.n645 B.n79 256.663
R974 B.n647 B.n79 256.663
R975 B.n653 B.n79 256.663
R976 B.n655 B.n79 256.663
R977 B.n661 B.n79 256.663
R978 B.n663 B.n79 256.663
R979 B.n669 B.n79 256.663
R980 B.n671 B.n79 256.663
R981 B.n677 B.n79 256.663
R982 B.n679 B.n79 256.663
R983 B.n685 B.n79 256.663
R984 B.n687 B.n79 256.663
R985 B.n693 B.n79 256.663
R986 B.n695 B.n79 256.663
R987 B.n372 B.n199 256.663
R988 B.n202 B.n199 256.663
R989 B.n365 B.n199 256.663
R990 B.n359 B.n199 256.663
R991 B.n357 B.n199 256.663
R992 B.n351 B.n199 256.663
R993 B.n349 B.n199 256.663
R994 B.n343 B.n199 256.663
R995 B.n341 B.n199 256.663
R996 B.n335 B.n199 256.663
R997 B.n333 B.n199 256.663
R998 B.n327 B.n199 256.663
R999 B.n325 B.n199 256.663
R1000 B.n319 B.n199 256.663
R1001 B.n317 B.n199 256.663
R1002 B.n311 B.n199 256.663
R1003 B.n309 B.n199 256.663
R1004 B.n303 B.n199 256.663
R1005 B.n301 B.n199 256.663
R1006 B.n294 B.n199 256.663
R1007 B.n292 B.n199 256.663
R1008 B.n286 B.n199 256.663
R1009 B.n284 B.n199 256.663
R1010 B.n278 B.n199 256.663
R1011 B.n276 B.n199 256.663
R1012 B.n270 B.n199 256.663
R1013 B.n268 B.n199 256.663
R1014 B.n262 B.n199 256.663
R1015 B.n260 B.n199 256.663
R1016 B.n254 B.n199 256.663
R1017 B.n252 B.n199 256.663
R1018 B.n246 B.n199 256.663
R1019 B.n244 B.n199 256.663
R1020 B.n239 B.n199 256.663
R1021 B.n787 B.n786 256.663
R1022 B.n104 B.t13 213.292
R1023 B.n225 B.t8 213.292
R1024 B.n96 B.t16 213.292
R1025 B.n218 B.t18 213.292
R1026 B.n696 B.n694 163.367
R1027 B.n692 B.n82 163.367
R1028 B.n688 B.n686 163.367
R1029 B.n684 B.n84 163.367
R1030 B.n680 B.n678 163.367
R1031 B.n676 B.n86 163.367
R1032 B.n672 B.n670 163.367
R1033 B.n668 B.n88 163.367
R1034 B.n664 B.n662 163.367
R1035 B.n660 B.n90 163.367
R1036 B.n656 B.n654 163.367
R1037 B.n652 B.n92 163.367
R1038 B.n648 B.n646 163.367
R1039 B.n644 B.n94 163.367
R1040 B.n640 B.n638 163.367
R1041 B.n635 B.n634 163.367
R1042 B.n632 B.n100 163.367
R1043 B.n628 B.n626 163.367
R1044 B.n624 B.n102 163.367
R1045 B.n619 B.n617 163.367
R1046 B.n615 B.n106 163.367
R1047 B.n611 B.n609 163.367
R1048 B.n607 B.n108 163.367
R1049 B.n603 B.n601 163.367
R1050 B.n599 B.n110 163.367
R1051 B.n595 B.n593 163.367
R1052 B.n591 B.n112 163.367
R1053 B.n587 B.n585 163.367
R1054 B.n583 B.n114 163.367
R1055 B.n579 B.n577 163.367
R1056 B.n575 B.n116 163.367
R1057 B.n571 B.n569 163.367
R1058 B.n567 B.n118 163.367
R1059 B.n563 B.n561 163.367
R1060 B.n379 B.n196 163.367
R1061 B.n383 B.n196 163.367
R1062 B.n383 B.n190 163.367
R1063 B.n391 B.n190 163.367
R1064 B.n391 B.n188 163.367
R1065 B.n395 B.n188 163.367
R1066 B.n395 B.n183 163.367
R1067 B.n404 B.n183 163.367
R1068 B.n404 B.n181 163.367
R1069 B.n408 B.n181 163.367
R1070 B.n408 B.n175 163.367
R1071 B.n416 B.n175 163.367
R1072 B.n416 B.n173 163.367
R1073 B.n420 B.n173 163.367
R1074 B.n420 B.n167 163.367
R1075 B.n428 B.n167 163.367
R1076 B.n428 B.n165 163.367
R1077 B.n432 B.n165 163.367
R1078 B.n432 B.n160 163.367
R1079 B.n441 B.n160 163.367
R1080 B.n441 B.n158 163.367
R1081 B.n445 B.n158 163.367
R1082 B.n445 B.n152 163.367
R1083 B.n453 B.n152 163.367
R1084 B.n453 B.n150 163.367
R1085 B.n457 B.n150 163.367
R1086 B.n457 B.n144 163.367
R1087 B.n465 B.n144 163.367
R1088 B.n465 B.n142 163.367
R1089 B.n469 B.n142 163.367
R1090 B.n469 B.n136 163.367
R1091 B.n477 B.n136 163.367
R1092 B.n477 B.n134 163.367
R1093 B.n481 B.n134 163.367
R1094 B.n481 B.n128 163.367
R1095 B.n489 B.n128 163.367
R1096 B.n489 B.n126 163.367
R1097 B.n494 B.n126 163.367
R1098 B.n494 B.n120 163.367
R1099 B.n502 B.n120 163.367
R1100 B.n503 B.n502 163.367
R1101 B.n503 B.n5 163.367
R1102 B.n6 B.n5 163.367
R1103 B.n7 B.n6 163.367
R1104 B.n509 B.n7 163.367
R1105 B.n510 B.n509 163.367
R1106 B.n510 B.n13 163.367
R1107 B.n14 B.n13 163.367
R1108 B.n15 B.n14 163.367
R1109 B.n515 B.n15 163.367
R1110 B.n515 B.n20 163.367
R1111 B.n21 B.n20 163.367
R1112 B.n22 B.n21 163.367
R1113 B.n520 B.n22 163.367
R1114 B.n520 B.n27 163.367
R1115 B.n28 B.n27 163.367
R1116 B.n29 B.n28 163.367
R1117 B.n525 B.n29 163.367
R1118 B.n525 B.n34 163.367
R1119 B.n35 B.n34 163.367
R1120 B.n36 B.n35 163.367
R1121 B.n530 B.n36 163.367
R1122 B.n530 B.n41 163.367
R1123 B.n42 B.n41 163.367
R1124 B.n43 B.n42 163.367
R1125 B.n535 B.n43 163.367
R1126 B.n535 B.n48 163.367
R1127 B.n49 B.n48 163.367
R1128 B.n50 B.n49 163.367
R1129 B.n540 B.n50 163.367
R1130 B.n540 B.n55 163.367
R1131 B.n56 B.n55 163.367
R1132 B.n57 B.n56 163.367
R1133 B.n545 B.n57 163.367
R1134 B.n545 B.n62 163.367
R1135 B.n63 B.n62 163.367
R1136 B.n64 B.n63 163.367
R1137 B.n550 B.n64 163.367
R1138 B.n550 B.n69 163.367
R1139 B.n70 B.n69 163.367
R1140 B.n71 B.n70 163.367
R1141 B.n555 B.n71 163.367
R1142 B.n555 B.n76 163.367
R1143 B.n77 B.n76 163.367
R1144 B.n78 B.n77 163.367
R1145 B.n373 B.n371 163.367
R1146 B.n371 B.n370 163.367
R1147 B.n367 B.n366 163.367
R1148 B.n364 B.n204 163.367
R1149 B.n360 B.n358 163.367
R1150 B.n356 B.n206 163.367
R1151 B.n352 B.n350 163.367
R1152 B.n348 B.n208 163.367
R1153 B.n344 B.n342 163.367
R1154 B.n340 B.n210 163.367
R1155 B.n336 B.n334 163.367
R1156 B.n332 B.n212 163.367
R1157 B.n328 B.n326 163.367
R1158 B.n324 B.n214 163.367
R1159 B.n320 B.n318 163.367
R1160 B.n316 B.n216 163.367
R1161 B.n312 B.n310 163.367
R1162 B.n308 B.n221 163.367
R1163 B.n304 B.n302 163.367
R1164 B.n300 B.n223 163.367
R1165 B.n295 B.n293 163.367
R1166 B.n291 B.n227 163.367
R1167 B.n287 B.n285 163.367
R1168 B.n283 B.n229 163.367
R1169 B.n279 B.n277 163.367
R1170 B.n275 B.n231 163.367
R1171 B.n271 B.n269 163.367
R1172 B.n267 B.n233 163.367
R1173 B.n263 B.n261 163.367
R1174 B.n259 B.n235 163.367
R1175 B.n255 B.n253 163.367
R1176 B.n251 B.n237 163.367
R1177 B.n247 B.n245 163.367
R1178 B.n243 B.n240 163.367
R1179 B.n377 B.n194 163.367
R1180 B.n385 B.n194 163.367
R1181 B.n385 B.n192 163.367
R1182 B.n389 B.n192 163.367
R1183 B.n389 B.n186 163.367
R1184 B.n398 B.n186 163.367
R1185 B.n398 B.n184 163.367
R1186 B.n402 B.n184 163.367
R1187 B.n402 B.n179 163.367
R1188 B.n410 B.n179 163.367
R1189 B.n410 B.n177 163.367
R1190 B.n414 B.n177 163.367
R1191 B.n414 B.n171 163.367
R1192 B.n422 B.n171 163.367
R1193 B.n422 B.n169 163.367
R1194 B.n426 B.n169 163.367
R1195 B.n426 B.n163 163.367
R1196 B.n435 B.n163 163.367
R1197 B.n435 B.n161 163.367
R1198 B.n439 B.n161 163.367
R1199 B.n439 B.n156 163.367
R1200 B.n447 B.n156 163.367
R1201 B.n447 B.n154 163.367
R1202 B.n451 B.n154 163.367
R1203 B.n451 B.n148 163.367
R1204 B.n459 B.n148 163.367
R1205 B.n459 B.n146 163.367
R1206 B.n463 B.n146 163.367
R1207 B.n463 B.n140 163.367
R1208 B.n471 B.n140 163.367
R1209 B.n471 B.n138 163.367
R1210 B.n475 B.n138 163.367
R1211 B.n475 B.n132 163.367
R1212 B.n483 B.n132 163.367
R1213 B.n483 B.n130 163.367
R1214 B.n487 B.n130 163.367
R1215 B.n487 B.n124 163.367
R1216 B.n496 B.n124 163.367
R1217 B.n496 B.n122 163.367
R1218 B.n500 B.n122 163.367
R1219 B.n500 B.n3 163.367
R1220 B.n785 B.n3 163.367
R1221 B.n781 B.n2 163.367
R1222 B.n781 B.n780 163.367
R1223 B.n780 B.n9 163.367
R1224 B.n776 B.n9 163.367
R1225 B.n776 B.n11 163.367
R1226 B.n772 B.n11 163.367
R1227 B.n772 B.n17 163.367
R1228 B.n768 B.n17 163.367
R1229 B.n768 B.n19 163.367
R1230 B.n764 B.n19 163.367
R1231 B.n764 B.n24 163.367
R1232 B.n760 B.n24 163.367
R1233 B.n760 B.n26 163.367
R1234 B.n756 B.n26 163.367
R1235 B.n756 B.n31 163.367
R1236 B.n752 B.n31 163.367
R1237 B.n752 B.n33 163.367
R1238 B.n748 B.n33 163.367
R1239 B.n748 B.n38 163.367
R1240 B.n744 B.n38 163.367
R1241 B.n744 B.n40 163.367
R1242 B.n740 B.n40 163.367
R1243 B.n740 B.n44 163.367
R1244 B.n736 B.n44 163.367
R1245 B.n736 B.n46 163.367
R1246 B.n732 B.n46 163.367
R1247 B.n732 B.n52 163.367
R1248 B.n728 B.n52 163.367
R1249 B.n728 B.n54 163.367
R1250 B.n724 B.n54 163.367
R1251 B.n724 B.n59 163.367
R1252 B.n720 B.n59 163.367
R1253 B.n720 B.n61 163.367
R1254 B.n716 B.n61 163.367
R1255 B.n716 B.n65 163.367
R1256 B.n712 B.n65 163.367
R1257 B.n712 B.n67 163.367
R1258 B.n708 B.n67 163.367
R1259 B.n708 B.n73 163.367
R1260 B.n704 B.n73 163.367
R1261 B.n704 B.n75 163.367
R1262 B.n700 B.n75 163.367
R1263 B.n378 B.n199 93.6352
R1264 B.n701 B.n79 93.6352
R1265 B.n695 B.n80 71.676
R1266 B.n694 B.n693 71.676
R1267 B.n687 B.n82 71.676
R1268 B.n686 B.n685 71.676
R1269 B.n679 B.n84 71.676
R1270 B.n678 B.n677 71.676
R1271 B.n671 B.n86 71.676
R1272 B.n670 B.n669 71.676
R1273 B.n663 B.n88 71.676
R1274 B.n662 B.n661 71.676
R1275 B.n655 B.n90 71.676
R1276 B.n654 B.n653 71.676
R1277 B.n647 B.n92 71.676
R1278 B.n646 B.n645 71.676
R1279 B.n639 B.n94 71.676
R1280 B.n638 B.n98 71.676
R1281 B.n634 B.n633 71.676
R1282 B.n627 B.n100 71.676
R1283 B.n626 B.n625 71.676
R1284 B.n618 B.n102 71.676
R1285 B.n617 B.n616 71.676
R1286 B.n610 B.n106 71.676
R1287 B.n609 B.n608 71.676
R1288 B.n602 B.n108 71.676
R1289 B.n601 B.n600 71.676
R1290 B.n594 B.n110 71.676
R1291 B.n593 B.n592 71.676
R1292 B.n586 B.n112 71.676
R1293 B.n585 B.n584 71.676
R1294 B.n578 B.n114 71.676
R1295 B.n577 B.n576 71.676
R1296 B.n570 B.n116 71.676
R1297 B.n569 B.n568 71.676
R1298 B.n562 B.n118 71.676
R1299 B.n563 B.n562 71.676
R1300 B.n568 B.n567 71.676
R1301 B.n571 B.n570 71.676
R1302 B.n576 B.n575 71.676
R1303 B.n579 B.n578 71.676
R1304 B.n584 B.n583 71.676
R1305 B.n587 B.n586 71.676
R1306 B.n592 B.n591 71.676
R1307 B.n595 B.n594 71.676
R1308 B.n600 B.n599 71.676
R1309 B.n603 B.n602 71.676
R1310 B.n608 B.n607 71.676
R1311 B.n611 B.n610 71.676
R1312 B.n616 B.n615 71.676
R1313 B.n619 B.n618 71.676
R1314 B.n625 B.n624 71.676
R1315 B.n628 B.n627 71.676
R1316 B.n633 B.n632 71.676
R1317 B.n635 B.n98 71.676
R1318 B.n640 B.n639 71.676
R1319 B.n645 B.n644 71.676
R1320 B.n648 B.n647 71.676
R1321 B.n653 B.n652 71.676
R1322 B.n656 B.n655 71.676
R1323 B.n661 B.n660 71.676
R1324 B.n664 B.n663 71.676
R1325 B.n669 B.n668 71.676
R1326 B.n672 B.n671 71.676
R1327 B.n677 B.n676 71.676
R1328 B.n680 B.n679 71.676
R1329 B.n685 B.n684 71.676
R1330 B.n688 B.n687 71.676
R1331 B.n693 B.n692 71.676
R1332 B.n696 B.n695 71.676
R1333 B.n372 B.n200 71.676
R1334 B.n370 B.n202 71.676
R1335 B.n366 B.n365 71.676
R1336 B.n359 B.n204 71.676
R1337 B.n358 B.n357 71.676
R1338 B.n351 B.n206 71.676
R1339 B.n350 B.n349 71.676
R1340 B.n343 B.n208 71.676
R1341 B.n342 B.n341 71.676
R1342 B.n335 B.n210 71.676
R1343 B.n334 B.n333 71.676
R1344 B.n327 B.n212 71.676
R1345 B.n326 B.n325 71.676
R1346 B.n319 B.n214 71.676
R1347 B.n318 B.n317 71.676
R1348 B.n311 B.n216 71.676
R1349 B.n310 B.n309 71.676
R1350 B.n303 B.n221 71.676
R1351 B.n302 B.n301 71.676
R1352 B.n294 B.n223 71.676
R1353 B.n293 B.n292 71.676
R1354 B.n286 B.n227 71.676
R1355 B.n285 B.n284 71.676
R1356 B.n278 B.n229 71.676
R1357 B.n277 B.n276 71.676
R1358 B.n270 B.n231 71.676
R1359 B.n269 B.n268 71.676
R1360 B.n262 B.n233 71.676
R1361 B.n261 B.n260 71.676
R1362 B.n254 B.n235 71.676
R1363 B.n253 B.n252 71.676
R1364 B.n246 B.n237 71.676
R1365 B.n245 B.n244 71.676
R1366 B.n240 B.n239 71.676
R1367 B.n373 B.n372 71.676
R1368 B.n367 B.n202 71.676
R1369 B.n365 B.n364 71.676
R1370 B.n360 B.n359 71.676
R1371 B.n357 B.n356 71.676
R1372 B.n352 B.n351 71.676
R1373 B.n349 B.n348 71.676
R1374 B.n344 B.n343 71.676
R1375 B.n341 B.n340 71.676
R1376 B.n336 B.n335 71.676
R1377 B.n333 B.n332 71.676
R1378 B.n328 B.n327 71.676
R1379 B.n325 B.n324 71.676
R1380 B.n320 B.n319 71.676
R1381 B.n317 B.n316 71.676
R1382 B.n312 B.n311 71.676
R1383 B.n309 B.n308 71.676
R1384 B.n304 B.n303 71.676
R1385 B.n301 B.n300 71.676
R1386 B.n295 B.n294 71.676
R1387 B.n292 B.n291 71.676
R1388 B.n287 B.n286 71.676
R1389 B.n284 B.n283 71.676
R1390 B.n279 B.n278 71.676
R1391 B.n276 B.n275 71.676
R1392 B.n271 B.n270 71.676
R1393 B.n268 B.n267 71.676
R1394 B.n263 B.n262 71.676
R1395 B.n260 B.n259 71.676
R1396 B.n255 B.n254 71.676
R1397 B.n252 B.n251 71.676
R1398 B.n247 B.n246 71.676
R1399 B.n244 B.n243 71.676
R1400 B.n239 B.n198 71.676
R1401 B.n786 B.n785 71.676
R1402 B.n786 B.n2 71.676
R1403 B.n97 B.n96 59.5399
R1404 B.n621 B.n104 59.5399
R1405 B.n298 B.n225 59.5399
R1406 B.n219 B.n218 59.5399
R1407 B.n96 B.n95 56.4369
R1408 B.n104 B.n103 56.4369
R1409 B.n225 B.n224 56.4369
R1410 B.n218 B.n217 56.4369
R1411 B.n378 B.n195 56.347
R1412 B.n384 B.n195 56.347
R1413 B.n384 B.n191 56.347
R1414 B.n390 B.n191 56.347
R1415 B.n390 B.n187 56.347
R1416 B.n397 B.n187 56.347
R1417 B.n397 B.n396 56.347
R1418 B.n403 B.n180 56.347
R1419 B.n409 B.n180 56.347
R1420 B.n409 B.n176 56.347
R1421 B.n415 B.n176 56.347
R1422 B.n415 B.n172 56.347
R1423 B.n421 B.n172 56.347
R1424 B.n421 B.n168 56.347
R1425 B.n427 B.n168 56.347
R1426 B.n427 B.n164 56.347
R1427 B.n434 B.n164 56.347
R1428 B.n434 B.n433 56.347
R1429 B.n440 B.n157 56.347
R1430 B.n446 B.n157 56.347
R1431 B.n446 B.n153 56.347
R1432 B.n452 B.n153 56.347
R1433 B.n452 B.n149 56.347
R1434 B.n458 B.n149 56.347
R1435 B.n458 B.n145 56.347
R1436 B.n464 B.n145 56.347
R1437 B.n470 B.n141 56.347
R1438 B.n470 B.n137 56.347
R1439 B.n476 B.n137 56.347
R1440 B.n476 B.n133 56.347
R1441 B.n482 B.n133 56.347
R1442 B.n482 B.n129 56.347
R1443 B.n488 B.n129 56.347
R1444 B.n495 B.n125 56.347
R1445 B.n495 B.n121 56.347
R1446 B.n501 B.n121 56.347
R1447 B.n501 B.n4 56.347
R1448 B.n784 B.n4 56.347
R1449 B.n784 B.n783 56.347
R1450 B.n783 B.n782 56.347
R1451 B.n782 B.n8 56.347
R1452 B.n12 B.n8 56.347
R1453 B.n775 B.n12 56.347
R1454 B.n775 B.n774 56.347
R1455 B.n773 B.n16 56.347
R1456 B.n767 B.n16 56.347
R1457 B.n767 B.n766 56.347
R1458 B.n766 B.n765 56.347
R1459 B.n765 B.n23 56.347
R1460 B.n759 B.n23 56.347
R1461 B.n759 B.n758 56.347
R1462 B.n757 B.n30 56.347
R1463 B.n751 B.n30 56.347
R1464 B.n751 B.n750 56.347
R1465 B.n750 B.n749 56.347
R1466 B.n749 B.n37 56.347
R1467 B.n743 B.n37 56.347
R1468 B.n743 B.n742 56.347
R1469 B.n742 B.n741 56.347
R1470 B.n735 B.n47 56.347
R1471 B.n735 B.n734 56.347
R1472 B.n734 B.n733 56.347
R1473 B.n733 B.n51 56.347
R1474 B.n727 B.n51 56.347
R1475 B.n727 B.n726 56.347
R1476 B.n726 B.n725 56.347
R1477 B.n725 B.n58 56.347
R1478 B.n719 B.n58 56.347
R1479 B.n719 B.n718 56.347
R1480 B.n718 B.n717 56.347
R1481 B.n711 B.n68 56.347
R1482 B.n711 B.n710 56.347
R1483 B.n710 B.n709 56.347
R1484 B.n709 B.n72 56.347
R1485 B.n703 B.n72 56.347
R1486 B.n703 B.n702 56.347
R1487 B.n702 B.n701 56.347
R1488 B.t5 B.n141 53.0325
R1489 B.n758 B.t0 53.0325
R1490 B.n396 B.t7 41.4318
R1491 B.n68 B.t11 41.4318
R1492 B.n488 B.t2 34.8028
R1493 B.t1 B.n773 34.8028
R1494 B.n376 B.n375 32.3127
R1495 B.n380 B.n197 32.3127
R1496 B.n560 B.n559 32.3127
R1497 B.n699 B.n698 32.3127
R1498 B.n433 B.t4 28.1738
R1499 B.n440 B.t4 28.1738
R1500 B.n741 B.t3 28.1738
R1501 B.n47 B.t3 28.1738
R1502 B.t2 B.n125 21.5448
R1503 B.n774 B.t1 21.5448
R1504 B B.n787 18.0485
R1505 B.n403 B.t7 14.9158
R1506 B.n717 B.t11 14.9158
R1507 B.n376 B.n193 10.6151
R1508 B.n386 B.n193 10.6151
R1509 B.n387 B.n386 10.6151
R1510 B.n388 B.n387 10.6151
R1511 B.n388 B.n185 10.6151
R1512 B.n399 B.n185 10.6151
R1513 B.n400 B.n399 10.6151
R1514 B.n401 B.n400 10.6151
R1515 B.n401 B.n178 10.6151
R1516 B.n411 B.n178 10.6151
R1517 B.n412 B.n411 10.6151
R1518 B.n413 B.n412 10.6151
R1519 B.n413 B.n170 10.6151
R1520 B.n423 B.n170 10.6151
R1521 B.n424 B.n423 10.6151
R1522 B.n425 B.n424 10.6151
R1523 B.n425 B.n162 10.6151
R1524 B.n436 B.n162 10.6151
R1525 B.n437 B.n436 10.6151
R1526 B.n438 B.n437 10.6151
R1527 B.n438 B.n155 10.6151
R1528 B.n448 B.n155 10.6151
R1529 B.n449 B.n448 10.6151
R1530 B.n450 B.n449 10.6151
R1531 B.n450 B.n147 10.6151
R1532 B.n460 B.n147 10.6151
R1533 B.n461 B.n460 10.6151
R1534 B.n462 B.n461 10.6151
R1535 B.n462 B.n139 10.6151
R1536 B.n472 B.n139 10.6151
R1537 B.n473 B.n472 10.6151
R1538 B.n474 B.n473 10.6151
R1539 B.n474 B.n131 10.6151
R1540 B.n484 B.n131 10.6151
R1541 B.n485 B.n484 10.6151
R1542 B.n486 B.n485 10.6151
R1543 B.n486 B.n123 10.6151
R1544 B.n497 B.n123 10.6151
R1545 B.n498 B.n497 10.6151
R1546 B.n499 B.n498 10.6151
R1547 B.n499 B.n0 10.6151
R1548 B.n375 B.n374 10.6151
R1549 B.n374 B.n201 10.6151
R1550 B.n369 B.n201 10.6151
R1551 B.n369 B.n368 10.6151
R1552 B.n368 B.n203 10.6151
R1553 B.n363 B.n203 10.6151
R1554 B.n363 B.n362 10.6151
R1555 B.n362 B.n361 10.6151
R1556 B.n361 B.n205 10.6151
R1557 B.n355 B.n205 10.6151
R1558 B.n355 B.n354 10.6151
R1559 B.n354 B.n353 10.6151
R1560 B.n353 B.n207 10.6151
R1561 B.n347 B.n207 10.6151
R1562 B.n347 B.n346 10.6151
R1563 B.n346 B.n345 10.6151
R1564 B.n345 B.n209 10.6151
R1565 B.n339 B.n209 10.6151
R1566 B.n339 B.n338 10.6151
R1567 B.n338 B.n337 10.6151
R1568 B.n337 B.n211 10.6151
R1569 B.n331 B.n211 10.6151
R1570 B.n331 B.n330 10.6151
R1571 B.n330 B.n329 10.6151
R1572 B.n329 B.n213 10.6151
R1573 B.n323 B.n213 10.6151
R1574 B.n323 B.n322 10.6151
R1575 B.n322 B.n321 10.6151
R1576 B.n321 B.n215 10.6151
R1577 B.n315 B.n314 10.6151
R1578 B.n314 B.n313 10.6151
R1579 B.n313 B.n220 10.6151
R1580 B.n307 B.n220 10.6151
R1581 B.n307 B.n306 10.6151
R1582 B.n306 B.n305 10.6151
R1583 B.n305 B.n222 10.6151
R1584 B.n299 B.n222 10.6151
R1585 B.n297 B.n296 10.6151
R1586 B.n296 B.n226 10.6151
R1587 B.n290 B.n226 10.6151
R1588 B.n290 B.n289 10.6151
R1589 B.n289 B.n288 10.6151
R1590 B.n288 B.n228 10.6151
R1591 B.n282 B.n228 10.6151
R1592 B.n282 B.n281 10.6151
R1593 B.n281 B.n280 10.6151
R1594 B.n280 B.n230 10.6151
R1595 B.n274 B.n230 10.6151
R1596 B.n274 B.n273 10.6151
R1597 B.n273 B.n272 10.6151
R1598 B.n272 B.n232 10.6151
R1599 B.n266 B.n232 10.6151
R1600 B.n266 B.n265 10.6151
R1601 B.n265 B.n264 10.6151
R1602 B.n264 B.n234 10.6151
R1603 B.n258 B.n234 10.6151
R1604 B.n258 B.n257 10.6151
R1605 B.n257 B.n256 10.6151
R1606 B.n256 B.n236 10.6151
R1607 B.n250 B.n236 10.6151
R1608 B.n250 B.n249 10.6151
R1609 B.n249 B.n248 10.6151
R1610 B.n248 B.n238 10.6151
R1611 B.n242 B.n238 10.6151
R1612 B.n242 B.n241 10.6151
R1613 B.n241 B.n197 10.6151
R1614 B.n381 B.n380 10.6151
R1615 B.n382 B.n381 10.6151
R1616 B.n382 B.n189 10.6151
R1617 B.n392 B.n189 10.6151
R1618 B.n393 B.n392 10.6151
R1619 B.n394 B.n393 10.6151
R1620 B.n394 B.n182 10.6151
R1621 B.n405 B.n182 10.6151
R1622 B.n406 B.n405 10.6151
R1623 B.n407 B.n406 10.6151
R1624 B.n407 B.n174 10.6151
R1625 B.n417 B.n174 10.6151
R1626 B.n418 B.n417 10.6151
R1627 B.n419 B.n418 10.6151
R1628 B.n419 B.n166 10.6151
R1629 B.n429 B.n166 10.6151
R1630 B.n430 B.n429 10.6151
R1631 B.n431 B.n430 10.6151
R1632 B.n431 B.n159 10.6151
R1633 B.n442 B.n159 10.6151
R1634 B.n443 B.n442 10.6151
R1635 B.n444 B.n443 10.6151
R1636 B.n444 B.n151 10.6151
R1637 B.n454 B.n151 10.6151
R1638 B.n455 B.n454 10.6151
R1639 B.n456 B.n455 10.6151
R1640 B.n456 B.n143 10.6151
R1641 B.n466 B.n143 10.6151
R1642 B.n467 B.n466 10.6151
R1643 B.n468 B.n467 10.6151
R1644 B.n468 B.n135 10.6151
R1645 B.n478 B.n135 10.6151
R1646 B.n479 B.n478 10.6151
R1647 B.n480 B.n479 10.6151
R1648 B.n480 B.n127 10.6151
R1649 B.n490 B.n127 10.6151
R1650 B.n491 B.n490 10.6151
R1651 B.n493 B.n491 10.6151
R1652 B.n493 B.n492 10.6151
R1653 B.n492 B.n119 10.6151
R1654 B.n504 B.n119 10.6151
R1655 B.n505 B.n504 10.6151
R1656 B.n506 B.n505 10.6151
R1657 B.n507 B.n506 10.6151
R1658 B.n508 B.n507 10.6151
R1659 B.n511 B.n508 10.6151
R1660 B.n512 B.n511 10.6151
R1661 B.n513 B.n512 10.6151
R1662 B.n514 B.n513 10.6151
R1663 B.n516 B.n514 10.6151
R1664 B.n517 B.n516 10.6151
R1665 B.n518 B.n517 10.6151
R1666 B.n519 B.n518 10.6151
R1667 B.n521 B.n519 10.6151
R1668 B.n522 B.n521 10.6151
R1669 B.n523 B.n522 10.6151
R1670 B.n524 B.n523 10.6151
R1671 B.n526 B.n524 10.6151
R1672 B.n527 B.n526 10.6151
R1673 B.n528 B.n527 10.6151
R1674 B.n529 B.n528 10.6151
R1675 B.n531 B.n529 10.6151
R1676 B.n532 B.n531 10.6151
R1677 B.n533 B.n532 10.6151
R1678 B.n534 B.n533 10.6151
R1679 B.n536 B.n534 10.6151
R1680 B.n537 B.n536 10.6151
R1681 B.n538 B.n537 10.6151
R1682 B.n539 B.n538 10.6151
R1683 B.n541 B.n539 10.6151
R1684 B.n542 B.n541 10.6151
R1685 B.n543 B.n542 10.6151
R1686 B.n544 B.n543 10.6151
R1687 B.n546 B.n544 10.6151
R1688 B.n547 B.n546 10.6151
R1689 B.n548 B.n547 10.6151
R1690 B.n549 B.n548 10.6151
R1691 B.n551 B.n549 10.6151
R1692 B.n552 B.n551 10.6151
R1693 B.n553 B.n552 10.6151
R1694 B.n554 B.n553 10.6151
R1695 B.n556 B.n554 10.6151
R1696 B.n557 B.n556 10.6151
R1697 B.n558 B.n557 10.6151
R1698 B.n559 B.n558 10.6151
R1699 B.n779 B.n1 10.6151
R1700 B.n779 B.n778 10.6151
R1701 B.n778 B.n777 10.6151
R1702 B.n777 B.n10 10.6151
R1703 B.n771 B.n10 10.6151
R1704 B.n771 B.n770 10.6151
R1705 B.n770 B.n769 10.6151
R1706 B.n769 B.n18 10.6151
R1707 B.n763 B.n18 10.6151
R1708 B.n763 B.n762 10.6151
R1709 B.n762 B.n761 10.6151
R1710 B.n761 B.n25 10.6151
R1711 B.n755 B.n25 10.6151
R1712 B.n755 B.n754 10.6151
R1713 B.n754 B.n753 10.6151
R1714 B.n753 B.n32 10.6151
R1715 B.n747 B.n32 10.6151
R1716 B.n747 B.n746 10.6151
R1717 B.n746 B.n745 10.6151
R1718 B.n745 B.n39 10.6151
R1719 B.n739 B.n39 10.6151
R1720 B.n739 B.n738 10.6151
R1721 B.n738 B.n737 10.6151
R1722 B.n737 B.n45 10.6151
R1723 B.n731 B.n45 10.6151
R1724 B.n731 B.n730 10.6151
R1725 B.n730 B.n729 10.6151
R1726 B.n729 B.n53 10.6151
R1727 B.n723 B.n53 10.6151
R1728 B.n723 B.n722 10.6151
R1729 B.n722 B.n721 10.6151
R1730 B.n721 B.n60 10.6151
R1731 B.n715 B.n60 10.6151
R1732 B.n715 B.n714 10.6151
R1733 B.n714 B.n713 10.6151
R1734 B.n713 B.n66 10.6151
R1735 B.n707 B.n66 10.6151
R1736 B.n707 B.n706 10.6151
R1737 B.n706 B.n705 10.6151
R1738 B.n705 B.n74 10.6151
R1739 B.n699 B.n74 10.6151
R1740 B.n698 B.n697 10.6151
R1741 B.n697 B.n81 10.6151
R1742 B.n691 B.n81 10.6151
R1743 B.n691 B.n690 10.6151
R1744 B.n690 B.n689 10.6151
R1745 B.n689 B.n83 10.6151
R1746 B.n683 B.n83 10.6151
R1747 B.n683 B.n682 10.6151
R1748 B.n682 B.n681 10.6151
R1749 B.n681 B.n85 10.6151
R1750 B.n675 B.n85 10.6151
R1751 B.n675 B.n674 10.6151
R1752 B.n674 B.n673 10.6151
R1753 B.n673 B.n87 10.6151
R1754 B.n667 B.n87 10.6151
R1755 B.n667 B.n666 10.6151
R1756 B.n666 B.n665 10.6151
R1757 B.n665 B.n89 10.6151
R1758 B.n659 B.n89 10.6151
R1759 B.n659 B.n658 10.6151
R1760 B.n658 B.n657 10.6151
R1761 B.n657 B.n91 10.6151
R1762 B.n651 B.n91 10.6151
R1763 B.n651 B.n650 10.6151
R1764 B.n650 B.n649 10.6151
R1765 B.n649 B.n93 10.6151
R1766 B.n643 B.n93 10.6151
R1767 B.n643 B.n642 10.6151
R1768 B.n642 B.n641 10.6151
R1769 B.n637 B.n636 10.6151
R1770 B.n636 B.n99 10.6151
R1771 B.n631 B.n99 10.6151
R1772 B.n631 B.n630 10.6151
R1773 B.n630 B.n629 10.6151
R1774 B.n629 B.n101 10.6151
R1775 B.n623 B.n101 10.6151
R1776 B.n623 B.n622 10.6151
R1777 B.n620 B.n105 10.6151
R1778 B.n614 B.n105 10.6151
R1779 B.n614 B.n613 10.6151
R1780 B.n613 B.n612 10.6151
R1781 B.n612 B.n107 10.6151
R1782 B.n606 B.n107 10.6151
R1783 B.n606 B.n605 10.6151
R1784 B.n605 B.n604 10.6151
R1785 B.n604 B.n109 10.6151
R1786 B.n598 B.n109 10.6151
R1787 B.n598 B.n597 10.6151
R1788 B.n597 B.n596 10.6151
R1789 B.n596 B.n111 10.6151
R1790 B.n590 B.n111 10.6151
R1791 B.n590 B.n589 10.6151
R1792 B.n589 B.n588 10.6151
R1793 B.n588 B.n113 10.6151
R1794 B.n582 B.n113 10.6151
R1795 B.n582 B.n581 10.6151
R1796 B.n581 B.n580 10.6151
R1797 B.n580 B.n115 10.6151
R1798 B.n574 B.n115 10.6151
R1799 B.n574 B.n573 10.6151
R1800 B.n573 B.n572 10.6151
R1801 B.n572 B.n117 10.6151
R1802 B.n566 B.n117 10.6151
R1803 B.n566 B.n565 10.6151
R1804 B.n565 B.n564 10.6151
R1805 B.n564 B.n560 10.6151
R1806 B.n787 B.n0 8.11757
R1807 B.n787 B.n1 8.11757
R1808 B.n315 B.n219 6.5566
R1809 B.n299 B.n298 6.5566
R1810 B.n637 B.n97 6.5566
R1811 B.n622 B.n621 6.5566
R1812 B.n219 B.n215 4.05904
R1813 B.n298 B.n297 4.05904
R1814 B.n641 B.n97 4.05904
R1815 B.n621 B.n620 4.05904
R1816 B.n464 B.t5 3.315
R1817 B.t0 B.n757 3.315
R1818 VP.n13 VP.n12 161.3
R1819 VP.n14 VP.n9 161.3
R1820 VP.n16 VP.n15 161.3
R1821 VP.n17 VP.n8 161.3
R1822 VP.n19 VP.n18 161.3
R1823 VP.n20 VP.n7 161.3
R1824 VP.n42 VP.n0 161.3
R1825 VP.n41 VP.n40 161.3
R1826 VP.n39 VP.n1 161.3
R1827 VP.n38 VP.n37 161.3
R1828 VP.n36 VP.n2 161.3
R1829 VP.n35 VP.n34 161.3
R1830 VP.n33 VP.n32 161.3
R1831 VP.n31 VP.n4 161.3
R1832 VP.n30 VP.n29 161.3
R1833 VP.n28 VP.n5 161.3
R1834 VP.n27 VP.n26 161.3
R1835 VP.n25 VP.n6 161.3
R1836 VP.n11 VP.t4 107.779
R1837 VP.n24 VP.n23 103.038
R1838 VP.n44 VP.n43 103.038
R1839 VP.n22 VP.n21 103.038
R1840 VP.n24 VP.t2 74.7292
R1841 VP.n3 VP.t1 74.7292
R1842 VP.n43 VP.t0 74.7292
R1843 VP.n21 VP.t5 74.7292
R1844 VP.n10 VP.t3 74.7292
R1845 VP.n11 VP.n10 60.2499
R1846 VP.n30 VP.n5 56.5617
R1847 VP.n37 VP.n1 56.5617
R1848 VP.n15 VP.n8 56.5617
R1849 VP.n23 VP.n22 45.5489
R1850 VP.n26 VP.n25 24.5923
R1851 VP.n26 VP.n5 24.5923
R1852 VP.n31 VP.n30 24.5923
R1853 VP.n32 VP.n31 24.5923
R1854 VP.n36 VP.n35 24.5923
R1855 VP.n37 VP.n36 24.5923
R1856 VP.n41 VP.n1 24.5923
R1857 VP.n42 VP.n41 24.5923
R1858 VP.n19 VP.n8 24.5923
R1859 VP.n20 VP.n19 24.5923
R1860 VP.n14 VP.n13 24.5923
R1861 VP.n15 VP.n14 24.5923
R1862 VP.n32 VP.n3 12.2964
R1863 VP.n35 VP.n3 12.2964
R1864 VP.n13 VP.n10 12.2964
R1865 VP.n25 VP.n24 7.86989
R1866 VP.n43 VP.n42 7.86989
R1867 VP.n21 VP.n20 7.86989
R1868 VP.n12 VP.n11 6.96699
R1869 VP.n22 VP.n7 0.278335
R1870 VP.n23 VP.n6 0.278335
R1871 VP.n44 VP.n0 0.278335
R1872 VP.n12 VP.n9 0.189894
R1873 VP.n16 VP.n9 0.189894
R1874 VP.n17 VP.n16 0.189894
R1875 VP.n18 VP.n17 0.189894
R1876 VP.n18 VP.n7 0.189894
R1877 VP.n27 VP.n6 0.189894
R1878 VP.n28 VP.n27 0.189894
R1879 VP.n29 VP.n28 0.189894
R1880 VP.n29 VP.n4 0.189894
R1881 VP.n33 VP.n4 0.189894
R1882 VP.n34 VP.n33 0.189894
R1883 VP.n34 VP.n2 0.189894
R1884 VP.n38 VP.n2 0.189894
R1885 VP.n39 VP.n38 0.189894
R1886 VP.n40 VP.n39 0.189894
R1887 VP.n40 VP.n0 0.189894
R1888 VP VP.n44 0.153485
R1889 VDD1.n36 VDD1.n0 289.615
R1890 VDD1.n77 VDD1.n41 289.615
R1891 VDD1.n37 VDD1.n36 185
R1892 VDD1.n35 VDD1.n2 185
R1893 VDD1.n34 VDD1.n33 185
R1894 VDD1.n5 VDD1.n3 185
R1895 VDD1.n28 VDD1.n27 185
R1896 VDD1.n26 VDD1.n25 185
R1897 VDD1.n9 VDD1.n8 185
R1898 VDD1.n20 VDD1.n19 185
R1899 VDD1.n18 VDD1.n17 185
R1900 VDD1.n13 VDD1.n12 185
R1901 VDD1.n53 VDD1.n52 185
R1902 VDD1.n58 VDD1.n57 185
R1903 VDD1.n60 VDD1.n59 185
R1904 VDD1.n49 VDD1.n48 185
R1905 VDD1.n66 VDD1.n65 185
R1906 VDD1.n68 VDD1.n67 185
R1907 VDD1.n45 VDD1.n44 185
R1908 VDD1.n75 VDD1.n74 185
R1909 VDD1.n76 VDD1.n43 185
R1910 VDD1.n78 VDD1.n77 185
R1911 VDD1.n14 VDD1.t1 149.524
R1912 VDD1.n54 VDD1.t3 149.524
R1913 VDD1.n36 VDD1.n35 104.615
R1914 VDD1.n35 VDD1.n34 104.615
R1915 VDD1.n34 VDD1.n3 104.615
R1916 VDD1.n27 VDD1.n3 104.615
R1917 VDD1.n27 VDD1.n26 104.615
R1918 VDD1.n26 VDD1.n8 104.615
R1919 VDD1.n19 VDD1.n8 104.615
R1920 VDD1.n19 VDD1.n18 104.615
R1921 VDD1.n18 VDD1.n12 104.615
R1922 VDD1.n58 VDD1.n52 104.615
R1923 VDD1.n59 VDD1.n58 104.615
R1924 VDD1.n59 VDD1.n48 104.615
R1925 VDD1.n66 VDD1.n48 104.615
R1926 VDD1.n67 VDD1.n66 104.615
R1927 VDD1.n67 VDD1.n44 104.615
R1928 VDD1.n75 VDD1.n44 104.615
R1929 VDD1.n76 VDD1.n75 104.615
R1930 VDD1.n77 VDD1.n76 104.615
R1931 VDD1.n83 VDD1.n82 68.4284
R1932 VDD1.n85 VDD1.n84 67.8566
R1933 VDD1 VDD1.n40 54.6826
R1934 VDD1.n83 VDD1.n81 54.569
R1935 VDD1.t1 VDD1.n12 52.3082
R1936 VDD1.t3 VDD1.n52 52.3082
R1937 VDD1.n85 VDD1.n83 40.6022
R1938 VDD1.n37 VDD1.n2 13.1884
R1939 VDD1.n78 VDD1.n43 13.1884
R1940 VDD1.n38 VDD1.n0 12.8005
R1941 VDD1.n33 VDD1.n4 12.8005
R1942 VDD1.n74 VDD1.n73 12.8005
R1943 VDD1.n79 VDD1.n41 12.8005
R1944 VDD1.n32 VDD1.n5 12.0247
R1945 VDD1.n72 VDD1.n45 12.0247
R1946 VDD1.n29 VDD1.n28 11.249
R1947 VDD1.n69 VDD1.n68 11.249
R1948 VDD1.n25 VDD1.n7 10.4732
R1949 VDD1.n65 VDD1.n47 10.4732
R1950 VDD1.n14 VDD1.n13 10.2747
R1951 VDD1.n54 VDD1.n53 10.2747
R1952 VDD1.n24 VDD1.n9 9.69747
R1953 VDD1.n64 VDD1.n49 9.69747
R1954 VDD1.n40 VDD1.n39 9.45567
R1955 VDD1.n81 VDD1.n80 9.45567
R1956 VDD1.n16 VDD1.n15 9.3005
R1957 VDD1.n11 VDD1.n10 9.3005
R1958 VDD1.n22 VDD1.n21 9.3005
R1959 VDD1.n24 VDD1.n23 9.3005
R1960 VDD1.n7 VDD1.n6 9.3005
R1961 VDD1.n30 VDD1.n29 9.3005
R1962 VDD1.n32 VDD1.n31 9.3005
R1963 VDD1.n4 VDD1.n1 9.3005
R1964 VDD1.n39 VDD1.n38 9.3005
R1965 VDD1.n80 VDD1.n79 9.3005
R1966 VDD1.n56 VDD1.n55 9.3005
R1967 VDD1.n51 VDD1.n50 9.3005
R1968 VDD1.n62 VDD1.n61 9.3005
R1969 VDD1.n64 VDD1.n63 9.3005
R1970 VDD1.n47 VDD1.n46 9.3005
R1971 VDD1.n70 VDD1.n69 9.3005
R1972 VDD1.n72 VDD1.n71 9.3005
R1973 VDD1.n73 VDD1.n42 9.3005
R1974 VDD1.n21 VDD1.n20 8.92171
R1975 VDD1.n61 VDD1.n60 8.92171
R1976 VDD1.n17 VDD1.n11 8.14595
R1977 VDD1.n57 VDD1.n51 8.14595
R1978 VDD1.n16 VDD1.n13 7.3702
R1979 VDD1.n56 VDD1.n53 7.3702
R1980 VDD1.n17 VDD1.n16 5.81868
R1981 VDD1.n57 VDD1.n56 5.81868
R1982 VDD1.n20 VDD1.n11 5.04292
R1983 VDD1.n60 VDD1.n51 5.04292
R1984 VDD1.n21 VDD1.n9 4.26717
R1985 VDD1.n61 VDD1.n49 4.26717
R1986 VDD1.n25 VDD1.n24 3.49141
R1987 VDD1.n65 VDD1.n64 3.49141
R1988 VDD1.n15 VDD1.n14 2.84304
R1989 VDD1.n55 VDD1.n54 2.84304
R1990 VDD1.n28 VDD1.n7 2.71565
R1991 VDD1.n68 VDD1.n47 2.71565
R1992 VDD1.n84 VDD1.t2 2.4755
R1993 VDD1.n84 VDD1.t0 2.4755
R1994 VDD1.n82 VDD1.t4 2.4755
R1995 VDD1.n82 VDD1.t5 2.4755
R1996 VDD1.n29 VDD1.n5 1.93989
R1997 VDD1.n69 VDD1.n45 1.93989
R1998 VDD1.n40 VDD1.n0 1.16414
R1999 VDD1.n33 VDD1.n32 1.16414
R2000 VDD1.n74 VDD1.n72 1.16414
R2001 VDD1.n81 VDD1.n41 1.16414
R2002 VDD1 VDD1.n85 0.569465
R2003 VDD1.n38 VDD1.n37 0.388379
R2004 VDD1.n4 VDD1.n2 0.388379
R2005 VDD1.n73 VDD1.n43 0.388379
R2006 VDD1.n79 VDD1.n78 0.388379
R2007 VDD1.n39 VDD1.n1 0.155672
R2008 VDD1.n31 VDD1.n1 0.155672
R2009 VDD1.n31 VDD1.n30 0.155672
R2010 VDD1.n30 VDD1.n6 0.155672
R2011 VDD1.n23 VDD1.n6 0.155672
R2012 VDD1.n23 VDD1.n22 0.155672
R2013 VDD1.n22 VDD1.n10 0.155672
R2014 VDD1.n15 VDD1.n10 0.155672
R2015 VDD1.n55 VDD1.n50 0.155672
R2016 VDD1.n62 VDD1.n50 0.155672
R2017 VDD1.n63 VDD1.n62 0.155672
R2018 VDD1.n63 VDD1.n46 0.155672
R2019 VDD1.n70 VDD1.n46 0.155672
R2020 VDD1.n71 VDD1.n70 0.155672
R2021 VDD1.n71 VDD1.n42 0.155672
R2022 VDD1.n80 VDD1.n42 0.155672
C0 VDD1 VDD2 1.39929f
C1 VN VP 6.16218f
C2 VTAIL VDD2 6.32315f
C3 VN VDD2 4.60026f
C4 VDD2 VP 0.456719f
C5 VTAIL VDD1 6.27154f
C6 VN VDD1 0.151126f
C7 VDD1 VP 4.90336f
C8 VN VTAIL 4.93054f
C9 VTAIL VP 4.94477f
C10 VDD2 B 5.257894f
C11 VDD1 B 5.394695f
C12 VTAIL B 6.207696f
C13 VN B 12.501869f
C14 VP B 11.176163f
C15 VDD1.n0 B 0.030357f
C16 VDD1.n1 B 0.02202f
C17 VDD1.n2 B 0.012181f
C18 VDD1.n3 B 0.027968f
C19 VDD1.n4 B 0.011833f
C20 VDD1.n5 B 0.012529f
C21 VDD1.n6 B 0.02202f
C22 VDD1.n7 B 0.011833f
C23 VDD1.n8 B 0.027968f
C24 VDD1.n9 B 0.012529f
C25 VDD1.n10 B 0.02202f
C26 VDD1.n11 B 0.011833f
C27 VDD1.n12 B 0.020976f
C28 VDD1.n13 B 0.019771f
C29 VDD1.t1 B 0.04678f
C30 VDD1.n14 B 0.124979f
C31 VDD1.n15 B 0.719066f
C32 VDD1.n16 B 0.011833f
C33 VDD1.n17 B 0.012529f
C34 VDD1.n18 B 0.027968f
C35 VDD1.n19 B 0.027968f
C36 VDD1.n20 B 0.012529f
C37 VDD1.n21 B 0.011833f
C38 VDD1.n22 B 0.02202f
C39 VDD1.n23 B 0.02202f
C40 VDD1.n24 B 0.011833f
C41 VDD1.n25 B 0.012529f
C42 VDD1.n26 B 0.027968f
C43 VDD1.n27 B 0.027968f
C44 VDD1.n28 B 0.012529f
C45 VDD1.n29 B 0.011833f
C46 VDD1.n30 B 0.02202f
C47 VDD1.n31 B 0.02202f
C48 VDD1.n32 B 0.011833f
C49 VDD1.n33 B 0.012529f
C50 VDD1.n34 B 0.027968f
C51 VDD1.n35 B 0.027968f
C52 VDD1.n36 B 0.059496f
C53 VDD1.n37 B 0.012181f
C54 VDD1.n38 B 0.011833f
C55 VDD1.n39 B 0.056915f
C56 VDD1.n40 B 0.055029f
C57 VDD1.n41 B 0.030357f
C58 VDD1.n42 B 0.02202f
C59 VDD1.n43 B 0.012181f
C60 VDD1.n44 B 0.027968f
C61 VDD1.n45 B 0.012529f
C62 VDD1.n46 B 0.02202f
C63 VDD1.n47 B 0.011833f
C64 VDD1.n48 B 0.027968f
C65 VDD1.n49 B 0.012529f
C66 VDD1.n50 B 0.02202f
C67 VDD1.n51 B 0.011833f
C68 VDD1.n52 B 0.020976f
C69 VDD1.n53 B 0.019771f
C70 VDD1.t3 B 0.04678f
C71 VDD1.n54 B 0.124979f
C72 VDD1.n55 B 0.719066f
C73 VDD1.n56 B 0.011833f
C74 VDD1.n57 B 0.012529f
C75 VDD1.n58 B 0.027968f
C76 VDD1.n59 B 0.027968f
C77 VDD1.n60 B 0.012529f
C78 VDD1.n61 B 0.011833f
C79 VDD1.n62 B 0.02202f
C80 VDD1.n63 B 0.02202f
C81 VDD1.n64 B 0.011833f
C82 VDD1.n65 B 0.012529f
C83 VDD1.n66 B 0.027968f
C84 VDD1.n67 B 0.027968f
C85 VDD1.n68 B 0.012529f
C86 VDD1.n69 B 0.011833f
C87 VDD1.n70 B 0.02202f
C88 VDD1.n71 B 0.02202f
C89 VDD1.n72 B 0.011833f
C90 VDD1.n73 B 0.011833f
C91 VDD1.n74 B 0.012529f
C92 VDD1.n75 B 0.027968f
C93 VDD1.n76 B 0.027968f
C94 VDD1.n77 B 0.059496f
C95 VDD1.n78 B 0.012181f
C96 VDD1.n79 B 0.011833f
C97 VDD1.n80 B 0.056915f
C98 VDD1.n81 B 0.054401f
C99 VDD1.t4 B 0.139209f
C100 VDD1.t5 B 0.139209f
C101 VDD1.n82 B 1.21005f
C102 VDD1.n83 B 2.23909f
C103 VDD1.t2 B 0.139209f
C104 VDD1.t0 B 0.139209f
C105 VDD1.n84 B 1.20669f
C106 VDD1.n85 B 2.17336f
C107 VP.n0 B 0.033368f
C108 VP.t0 B 1.40305f
C109 VP.n1 B 0.039944f
C110 VP.n2 B 0.025311f
C111 VP.t1 B 1.40305f
C112 VP.n3 B 0.511189f
C113 VP.n4 B 0.025311f
C114 VP.n5 B 0.039944f
C115 VP.n6 B 0.033368f
C116 VP.t2 B 1.40305f
C117 VP.n7 B 0.033368f
C118 VP.t5 B 1.40305f
C119 VP.n8 B 0.039944f
C120 VP.n9 B 0.025311f
C121 VP.t3 B 1.40305f
C122 VP.n10 B 0.583336f
C123 VP.t4 B 1.60706f
C124 VP.n11 B 0.564035f
C125 VP.n12 B 0.244023f
C126 VP.n13 B 0.035351f
C127 VP.n14 B 0.046937f
C128 VP.n15 B 0.033642f
C129 VP.n16 B 0.025311f
C130 VP.n17 B 0.025311f
C131 VP.n18 B 0.025311f
C132 VP.n19 B 0.046937f
C133 VP.n20 B 0.03118f
C134 VP.n21 B 0.591889f
C135 VP.n22 B 1.22493f
C136 VP.n23 B 1.24497f
C137 VP.n24 B 0.591889f
C138 VP.n25 B 0.03118f
C139 VP.n26 B 0.046937f
C140 VP.n27 B 0.025311f
C141 VP.n28 B 0.025311f
C142 VP.n29 B 0.025311f
C143 VP.n30 B 0.033642f
C144 VP.n31 B 0.046937f
C145 VP.n32 B 0.035351f
C146 VP.n33 B 0.025311f
C147 VP.n34 B 0.025311f
C148 VP.n35 B 0.035351f
C149 VP.n36 B 0.046937f
C150 VP.n37 B 0.033642f
C151 VP.n38 B 0.025311f
C152 VP.n39 B 0.025311f
C153 VP.n40 B 0.025311f
C154 VP.n41 B 0.046937f
C155 VP.n42 B 0.03118f
C156 VP.n43 B 0.591889f
C157 VP.n44 B 0.04234f
C158 VDD2.n0 B 0.02976f
C159 VDD2.n1 B 0.021587f
C160 VDD2.n2 B 0.011941f
C161 VDD2.n3 B 0.027418f
C162 VDD2.n4 B 0.012282f
C163 VDD2.n5 B 0.021587f
C164 VDD2.n6 B 0.0116f
C165 VDD2.n7 B 0.027418f
C166 VDD2.n8 B 0.012282f
C167 VDD2.n9 B 0.021587f
C168 VDD2.n10 B 0.0116f
C169 VDD2.n11 B 0.020564f
C170 VDD2.n12 B 0.019383f
C171 VDD2.t5 B 0.04586f
C172 VDD2.n13 B 0.122521f
C173 VDD2.n14 B 0.704925f
C174 VDD2.n15 B 0.0116f
C175 VDD2.n16 B 0.012282f
C176 VDD2.n17 B 0.027418f
C177 VDD2.n18 B 0.027418f
C178 VDD2.n19 B 0.012282f
C179 VDD2.n20 B 0.0116f
C180 VDD2.n21 B 0.021587f
C181 VDD2.n22 B 0.021587f
C182 VDD2.n23 B 0.0116f
C183 VDD2.n24 B 0.012282f
C184 VDD2.n25 B 0.027418f
C185 VDD2.n26 B 0.027418f
C186 VDD2.n27 B 0.012282f
C187 VDD2.n28 B 0.0116f
C188 VDD2.n29 B 0.021587f
C189 VDD2.n30 B 0.021587f
C190 VDD2.n31 B 0.0116f
C191 VDD2.n32 B 0.0116f
C192 VDD2.n33 B 0.012282f
C193 VDD2.n34 B 0.027418f
C194 VDD2.n35 B 0.027418f
C195 VDD2.n36 B 0.058326f
C196 VDD2.n37 B 0.011941f
C197 VDD2.n38 B 0.0116f
C198 VDD2.n39 B 0.055796f
C199 VDD2.n40 B 0.053331f
C200 VDD2.t4 B 0.136471f
C201 VDD2.t3 B 0.136471f
C202 VDD2.n41 B 1.18625f
C203 VDD2.n42 B 2.09133f
C204 VDD2.n43 B 0.02976f
C205 VDD2.n44 B 0.021587f
C206 VDD2.n45 B 0.011941f
C207 VDD2.n46 B 0.027418f
C208 VDD2.n47 B 0.0116f
C209 VDD2.n48 B 0.012282f
C210 VDD2.n49 B 0.021587f
C211 VDD2.n50 B 0.0116f
C212 VDD2.n51 B 0.027418f
C213 VDD2.n52 B 0.012282f
C214 VDD2.n53 B 0.021587f
C215 VDD2.n54 B 0.0116f
C216 VDD2.n55 B 0.020564f
C217 VDD2.n56 B 0.019383f
C218 VDD2.t0 B 0.04586f
C219 VDD2.n57 B 0.122521f
C220 VDD2.n58 B 0.704925f
C221 VDD2.n59 B 0.0116f
C222 VDD2.n60 B 0.012282f
C223 VDD2.n61 B 0.027418f
C224 VDD2.n62 B 0.027418f
C225 VDD2.n63 B 0.012282f
C226 VDD2.n64 B 0.0116f
C227 VDD2.n65 B 0.021587f
C228 VDD2.n66 B 0.021587f
C229 VDD2.n67 B 0.0116f
C230 VDD2.n68 B 0.012282f
C231 VDD2.n69 B 0.027418f
C232 VDD2.n70 B 0.027418f
C233 VDD2.n71 B 0.012282f
C234 VDD2.n72 B 0.0116f
C235 VDD2.n73 B 0.021587f
C236 VDD2.n74 B 0.021587f
C237 VDD2.n75 B 0.0116f
C238 VDD2.n76 B 0.012282f
C239 VDD2.n77 B 0.027418f
C240 VDD2.n78 B 0.027418f
C241 VDD2.n79 B 0.058326f
C242 VDD2.n80 B 0.011941f
C243 VDD2.n81 B 0.0116f
C244 VDD2.n82 B 0.055796f
C245 VDD2.n83 B 0.047567f
C246 VDD2.n84 B 1.94119f
C247 VDD2.t1 B 0.136471f
C248 VDD2.t2 B 0.136471f
C249 VDD2.n85 B 1.18623f
C250 VTAIL.t6 B 0.159315f
C251 VTAIL.t7 B 0.159315f
C252 VTAIL.n0 B 1.31766f
C253 VTAIL.n1 B 0.423775f
C254 VTAIL.n2 B 0.034742f
C255 VTAIL.n3 B 0.025201f
C256 VTAIL.n4 B 0.01394f
C257 VTAIL.n5 B 0.032008f
C258 VTAIL.n6 B 0.014338f
C259 VTAIL.n7 B 0.025201f
C260 VTAIL.n8 B 0.013542f
C261 VTAIL.n9 B 0.032008f
C262 VTAIL.n10 B 0.014338f
C263 VTAIL.n11 B 0.025201f
C264 VTAIL.n12 B 0.013542f
C265 VTAIL.n13 B 0.024006f
C266 VTAIL.n14 B 0.022627f
C267 VTAIL.t2 B 0.053536f
C268 VTAIL.n15 B 0.14303f
C269 VTAIL.n16 B 0.822921f
C270 VTAIL.n17 B 0.013542f
C271 VTAIL.n18 B 0.014338f
C272 VTAIL.n19 B 0.032008f
C273 VTAIL.n20 B 0.032008f
C274 VTAIL.n21 B 0.014338f
C275 VTAIL.n22 B 0.013542f
C276 VTAIL.n23 B 0.025201f
C277 VTAIL.n24 B 0.025201f
C278 VTAIL.n25 B 0.013542f
C279 VTAIL.n26 B 0.014338f
C280 VTAIL.n27 B 0.032008f
C281 VTAIL.n28 B 0.032008f
C282 VTAIL.n29 B 0.014338f
C283 VTAIL.n30 B 0.013542f
C284 VTAIL.n31 B 0.025201f
C285 VTAIL.n32 B 0.025201f
C286 VTAIL.n33 B 0.013542f
C287 VTAIL.n34 B 0.013542f
C288 VTAIL.n35 B 0.014338f
C289 VTAIL.n36 B 0.032008f
C290 VTAIL.n37 B 0.032008f
C291 VTAIL.n38 B 0.068089f
C292 VTAIL.n39 B 0.01394f
C293 VTAIL.n40 B 0.013542f
C294 VTAIL.n41 B 0.065136f
C295 VTAIL.n42 B 0.038176f
C296 VTAIL.n43 B 0.36913f
C297 VTAIL.t4 B 0.159315f
C298 VTAIL.t5 B 0.159315f
C299 VTAIL.n44 B 1.31766f
C300 VTAIL.n45 B 1.74158f
C301 VTAIL.t10 B 0.159315f
C302 VTAIL.t9 B 0.159315f
C303 VTAIL.n46 B 1.31767f
C304 VTAIL.n47 B 1.74157f
C305 VTAIL.n48 B 0.034742f
C306 VTAIL.n49 B 0.025201f
C307 VTAIL.n50 B 0.01394f
C308 VTAIL.n51 B 0.032008f
C309 VTAIL.n52 B 0.013542f
C310 VTAIL.n53 B 0.014338f
C311 VTAIL.n54 B 0.025201f
C312 VTAIL.n55 B 0.013542f
C313 VTAIL.n56 B 0.032008f
C314 VTAIL.n57 B 0.014338f
C315 VTAIL.n58 B 0.025201f
C316 VTAIL.n59 B 0.013542f
C317 VTAIL.n60 B 0.024006f
C318 VTAIL.n61 B 0.022627f
C319 VTAIL.t8 B 0.053536f
C320 VTAIL.n62 B 0.14303f
C321 VTAIL.n63 B 0.822921f
C322 VTAIL.n64 B 0.013542f
C323 VTAIL.n65 B 0.014338f
C324 VTAIL.n66 B 0.032008f
C325 VTAIL.n67 B 0.032008f
C326 VTAIL.n68 B 0.014338f
C327 VTAIL.n69 B 0.013542f
C328 VTAIL.n70 B 0.025201f
C329 VTAIL.n71 B 0.025201f
C330 VTAIL.n72 B 0.013542f
C331 VTAIL.n73 B 0.014338f
C332 VTAIL.n74 B 0.032008f
C333 VTAIL.n75 B 0.032008f
C334 VTAIL.n76 B 0.014338f
C335 VTAIL.n77 B 0.013542f
C336 VTAIL.n78 B 0.025201f
C337 VTAIL.n79 B 0.025201f
C338 VTAIL.n80 B 0.013542f
C339 VTAIL.n81 B 0.014338f
C340 VTAIL.n82 B 0.032008f
C341 VTAIL.n83 B 0.032008f
C342 VTAIL.n84 B 0.068089f
C343 VTAIL.n85 B 0.01394f
C344 VTAIL.n86 B 0.013542f
C345 VTAIL.n87 B 0.065136f
C346 VTAIL.n88 B 0.038176f
C347 VTAIL.n89 B 0.36913f
C348 VTAIL.t1 B 0.159315f
C349 VTAIL.t0 B 0.159315f
C350 VTAIL.n90 B 1.31767f
C351 VTAIL.n91 B 0.571821f
C352 VTAIL.n92 B 0.034742f
C353 VTAIL.n93 B 0.025201f
C354 VTAIL.n94 B 0.01394f
C355 VTAIL.n95 B 0.032008f
C356 VTAIL.n96 B 0.013542f
C357 VTAIL.n97 B 0.014338f
C358 VTAIL.n98 B 0.025201f
C359 VTAIL.n99 B 0.013542f
C360 VTAIL.n100 B 0.032008f
C361 VTAIL.n101 B 0.014338f
C362 VTAIL.n102 B 0.025201f
C363 VTAIL.n103 B 0.013542f
C364 VTAIL.n104 B 0.024006f
C365 VTAIL.n105 B 0.022627f
C366 VTAIL.t3 B 0.053536f
C367 VTAIL.n106 B 0.14303f
C368 VTAIL.n107 B 0.822921f
C369 VTAIL.n108 B 0.013542f
C370 VTAIL.n109 B 0.014338f
C371 VTAIL.n110 B 0.032008f
C372 VTAIL.n111 B 0.032008f
C373 VTAIL.n112 B 0.014338f
C374 VTAIL.n113 B 0.013542f
C375 VTAIL.n114 B 0.025201f
C376 VTAIL.n115 B 0.025201f
C377 VTAIL.n116 B 0.013542f
C378 VTAIL.n117 B 0.014338f
C379 VTAIL.n118 B 0.032008f
C380 VTAIL.n119 B 0.032008f
C381 VTAIL.n120 B 0.014338f
C382 VTAIL.n121 B 0.013542f
C383 VTAIL.n122 B 0.025201f
C384 VTAIL.n123 B 0.025201f
C385 VTAIL.n124 B 0.013542f
C386 VTAIL.n125 B 0.014338f
C387 VTAIL.n126 B 0.032008f
C388 VTAIL.n127 B 0.032008f
C389 VTAIL.n128 B 0.068089f
C390 VTAIL.n129 B 0.01394f
C391 VTAIL.n130 B 0.013542f
C392 VTAIL.n131 B 0.065136f
C393 VTAIL.n132 B 0.038176f
C394 VTAIL.n133 B 1.33517f
C395 VTAIL.n134 B 0.034742f
C396 VTAIL.n135 B 0.025201f
C397 VTAIL.n136 B 0.01394f
C398 VTAIL.n137 B 0.032008f
C399 VTAIL.n138 B 0.014338f
C400 VTAIL.n139 B 0.025201f
C401 VTAIL.n140 B 0.013542f
C402 VTAIL.n141 B 0.032008f
C403 VTAIL.n142 B 0.014338f
C404 VTAIL.n143 B 0.025201f
C405 VTAIL.n144 B 0.013542f
C406 VTAIL.n145 B 0.024006f
C407 VTAIL.n146 B 0.022627f
C408 VTAIL.t11 B 0.053536f
C409 VTAIL.n147 B 0.14303f
C410 VTAIL.n148 B 0.822921f
C411 VTAIL.n149 B 0.013542f
C412 VTAIL.n150 B 0.014338f
C413 VTAIL.n151 B 0.032008f
C414 VTAIL.n152 B 0.032008f
C415 VTAIL.n153 B 0.014338f
C416 VTAIL.n154 B 0.013542f
C417 VTAIL.n155 B 0.025201f
C418 VTAIL.n156 B 0.025201f
C419 VTAIL.n157 B 0.013542f
C420 VTAIL.n158 B 0.014338f
C421 VTAIL.n159 B 0.032008f
C422 VTAIL.n160 B 0.032008f
C423 VTAIL.n161 B 0.014338f
C424 VTAIL.n162 B 0.013542f
C425 VTAIL.n163 B 0.025201f
C426 VTAIL.n164 B 0.025201f
C427 VTAIL.n165 B 0.013542f
C428 VTAIL.n166 B 0.013542f
C429 VTAIL.n167 B 0.014338f
C430 VTAIL.n168 B 0.032008f
C431 VTAIL.n169 B 0.032008f
C432 VTAIL.n170 B 0.068089f
C433 VTAIL.n171 B 0.01394f
C434 VTAIL.n172 B 0.013542f
C435 VTAIL.n173 B 0.065136f
C436 VTAIL.n174 B 0.038176f
C437 VTAIL.n175 B 1.27952f
C438 VN.n0 B 0.03267f
C439 VN.t2 B 1.37369f
C440 VN.n1 B 0.039109f
C441 VN.n2 B 0.024781f
C442 VN.t1 B 1.37369f
C443 VN.n3 B 0.571128f
C444 VN.t0 B 1.57343f
C445 VN.n4 B 0.552232f
C446 VN.n5 B 0.238916f
C447 VN.n6 B 0.034611f
C448 VN.n7 B 0.045954f
C449 VN.n8 B 0.032938f
C450 VN.n9 B 0.024781f
C451 VN.n10 B 0.024781f
C452 VN.n11 B 0.024781f
C453 VN.n12 B 0.045954f
C454 VN.n13 B 0.030528f
C455 VN.n14 B 0.579502f
C456 VN.n15 B 0.041454f
C457 VN.n16 B 0.03267f
C458 VN.t5 B 1.37369f
C459 VN.n17 B 0.039109f
C460 VN.n18 B 0.024781f
C461 VN.t4 B 1.37369f
C462 VN.n19 B 0.571128f
C463 VN.t3 B 1.57343f
C464 VN.n20 B 0.552232f
C465 VN.n21 B 0.238916f
C466 VN.n22 B 0.034611f
C467 VN.n23 B 0.045954f
C468 VN.n24 B 0.032938f
C469 VN.n25 B 0.024781f
C470 VN.n26 B 0.024781f
C471 VN.n27 B 0.024781f
C472 VN.n28 B 0.045954f
C473 VN.n29 B 0.030528f
C474 VN.n30 B 0.579502f
C475 VN.n31 B 1.21282f
.ends

