* NGSPICE file created from diff_pair_sample_0318.ext - technology: sky130A

.subckt diff_pair_sample_0318 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.14675 pd=7.28 as=2.7105 ps=14.68 w=6.95 l=3.5
X1 VDD1.t2 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.14675 pd=7.28 as=2.7105 ps=14.68 w=6.95 l=3.5
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=0 ps=0 w=6.95 l=3.5
X3 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.14675 pd=7.28 as=2.7105 ps=14.68 w=6.95 l=3.5
X4 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=1.14675 ps=7.28 w=6.95 l=3.5
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=0 ps=0 w=6.95 l=3.5
X6 VTAIL.t7 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=1.14675 ps=7.28 w=6.95 l=3.5
X7 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.14675 pd=7.28 as=2.7105 ps=14.68 w=6.95 l=3.5
X8 VTAIL.t5 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=1.14675 ps=7.28 w=6.95 l=3.5
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=0 ps=0 w=6.95 l=3.5
X10 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=1.14675 ps=7.28 w=6.95 l=3.5
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7105 pd=14.68 as=0 ps=0 w=6.95 l=3.5
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n5 VP.t2 82.2952
R9 VP.n7 VP.n6 81.9933
R10 VP.n20 VP.n0 81.9933
R11 VP.n5 VP.t0 81.0755
R12 VP.n12 VP.n2 56.5193
R13 VP.n6 VP.t3 47.8562
R14 VP.n0 VP.t1 47.8562
R15 VP.n7 VP.n5 47.4711
R16 VP.n10 VP.n4 24.4675
R17 VP.n11 VP.n10 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n16 VP.n2 24.4675
R20 VP.n17 VP.n16 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n6 VP.n4 8.07461
R23 VP.n18 VP.n0 8.07461
R24 VP.n8 VP.n7 0.354971
R25 VP.n20 VP.n19 0.354971
R26 VP VP.n20 0.26696
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VTAIL.n5 VTAIL.t7 55.6507
R35 VTAIL.n4 VTAIL.t2 55.6507
R36 VTAIL.n3 VTAIL.t1 55.6507
R37 VTAIL.n7 VTAIL.t0 55.6505
R38 VTAIL.n0 VTAIL.t3 55.6505
R39 VTAIL.n1 VTAIL.t6 55.6505
R40 VTAIL.n2 VTAIL.t5 55.6505
R41 VTAIL.n6 VTAIL.t4 55.6505
R42 VTAIL.n7 VTAIL.n6 21.66
R43 VTAIL.n3 VTAIL.n2 21.66
R44 VTAIL.n4 VTAIL.n3 3.30222
R45 VTAIL.n6 VTAIL.n5 3.30222
R46 VTAIL.n2 VTAIL.n1 3.30222
R47 VTAIL VTAIL.n0 1.70955
R48 VTAIL VTAIL.n7 1.59317
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 VDD1 VDD1.n1 109.615
R52 VDD1 VDD1.n0 69.5386
R53 VDD1.n0 VDD1.t1 2.84942
R54 VDD1.n0 VDD1.t3 2.84942
R55 VDD1.n1 VDD1.t0 2.84942
R56 VDD1.n1 VDD1.t2 2.84942
R57 B.n540 B.n539 585
R58 B.n540 B.n78 585
R59 B.n543 B.n542 585
R60 B.n544 B.n114 585
R61 B.n546 B.n545 585
R62 B.n548 B.n113 585
R63 B.n551 B.n550 585
R64 B.n552 B.n112 585
R65 B.n554 B.n553 585
R66 B.n556 B.n111 585
R67 B.n559 B.n558 585
R68 B.n560 B.n110 585
R69 B.n562 B.n561 585
R70 B.n564 B.n109 585
R71 B.n567 B.n566 585
R72 B.n568 B.n108 585
R73 B.n570 B.n569 585
R74 B.n572 B.n107 585
R75 B.n575 B.n574 585
R76 B.n576 B.n106 585
R77 B.n578 B.n577 585
R78 B.n580 B.n105 585
R79 B.n583 B.n582 585
R80 B.n584 B.n104 585
R81 B.n586 B.n585 585
R82 B.n588 B.n103 585
R83 B.n591 B.n590 585
R84 B.n592 B.n100 585
R85 B.n595 B.n594 585
R86 B.n597 B.n99 585
R87 B.n600 B.n599 585
R88 B.n601 B.n98 585
R89 B.n603 B.n602 585
R90 B.n605 B.n97 585
R91 B.n608 B.n607 585
R92 B.n609 B.n93 585
R93 B.n611 B.n610 585
R94 B.n613 B.n92 585
R95 B.n616 B.n615 585
R96 B.n617 B.n91 585
R97 B.n619 B.n618 585
R98 B.n621 B.n90 585
R99 B.n624 B.n623 585
R100 B.n625 B.n89 585
R101 B.n627 B.n626 585
R102 B.n629 B.n88 585
R103 B.n632 B.n631 585
R104 B.n633 B.n87 585
R105 B.n635 B.n634 585
R106 B.n637 B.n86 585
R107 B.n640 B.n639 585
R108 B.n641 B.n85 585
R109 B.n643 B.n642 585
R110 B.n645 B.n84 585
R111 B.n648 B.n647 585
R112 B.n649 B.n83 585
R113 B.n651 B.n650 585
R114 B.n653 B.n82 585
R115 B.n656 B.n655 585
R116 B.n657 B.n81 585
R117 B.n659 B.n658 585
R118 B.n661 B.n80 585
R119 B.n664 B.n663 585
R120 B.n665 B.n79 585
R121 B.n538 B.n77 585
R122 B.n668 B.n77 585
R123 B.n537 B.n76 585
R124 B.n669 B.n76 585
R125 B.n536 B.n75 585
R126 B.n670 B.n75 585
R127 B.n535 B.n534 585
R128 B.n534 B.n71 585
R129 B.n533 B.n70 585
R130 B.n676 B.n70 585
R131 B.n532 B.n69 585
R132 B.n677 B.n69 585
R133 B.n531 B.n68 585
R134 B.n678 B.n68 585
R135 B.n530 B.n529 585
R136 B.n529 B.n64 585
R137 B.n528 B.n63 585
R138 B.n684 B.n63 585
R139 B.n527 B.n62 585
R140 B.n685 B.n62 585
R141 B.n526 B.n61 585
R142 B.n686 B.n61 585
R143 B.n525 B.n524 585
R144 B.n524 B.n57 585
R145 B.n523 B.n56 585
R146 B.n692 B.n56 585
R147 B.n522 B.n55 585
R148 B.n693 B.n55 585
R149 B.n521 B.n54 585
R150 B.n694 B.n54 585
R151 B.n520 B.n519 585
R152 B.n519 B.n50 585
R153 B.n518 B.n49 585
R154 B.n700 B.n49 585
R155 B.n517 B.n48 585
R156 B.n701 B.n48 585
R157 B.n516 B.n47 585
R158 B.n702 B.n47 585
R159 B.n515 B.n514 585
R160 B.n514 B.n43 585
R161 B.n513 B.n42 585
R162 B.n708 B.n42 585
R163 B.n512 B.n41 585
R164 B.n709 B.n41 585
R165 B.n511 B.n40 585
R166 B.n710 B.n40 585
R167 B.n510 B.n509 585
R168 B.n509 B.n39 585
R169 B.n508 B.n35 585
R170 B.n716 B.n35 585
R171 B.n507 B.n34 585
R172 B.n717 B.n34 585
R173 B.n506 B.n33 585
R174 B.n718 B.n33 585
R175 B.n505 B.n504 585
R176 B.n504 B.n29 585
R177 B.n503 B.n28 585
R178 B.n724 B.n28 585
R179 B.n502 B.n27 585
R180 B.n725 B.n27 585
R181 B.n501 B.n26 585
R182 B.n726 B.n26 585
R183 B.n500 B.n499 585
R184 B.n499 B.n22 585
R185 B.n498 B.n21 585
R186 B.n732 B.n21 585
R187 B.n497 B.n20 585
R188 B.n733 B.n20 585
R189 B.n496 B.n19 585
R190 B.n734 B.n19 585
R191 B.n495 B.n494 585
R192 B.n494 B.n15 585
R193 B.n493 B.n14 585
R194 B.n740 B.n14 585
R195 B.n492 B.n13 585
R196 B.n741 B.n13 585
R197 B.n491 B.n12 585
R198 B.n742 B.n12 585
R199 B.n490 B.n489 585
R200 B.n489 B.n8 585
R201 B.n488 B.n7 585
R202 B.n748 B.n7 585
R203 B.n487 B.n6 585
R204 B.n749 B.n6 585
R205 B.n486 B.n5 585
R206 B.n750 B.n5 585
R207 B.n485 B.n484 585
R208 B.n484 B.n4 585
R209 B.n483 B.n115 585
R210 B.n483 B.n482 585
R211 B.n473 B.n116 585
R212 B.n117 B.n116 585
R213 B.n475 B.n474 585
R214 B.n476 B.n475 585
R215 B.n472 B.n122 585
R216 B.n122 B.n121 585
R217 B.n471 B.n470 585
R218 B.n470 B.n469 585
R219 B.n124 B.n123 585
R220 B.n125 B.n124 585
R221 B.n462 B.n461 585
R222 B.n463 B.n462 585
R223 B.n460 B.n130 585
R224 B.n130 B.n129 585
R225 B.n459 B.n458 585
R226 B.n458 B.n457 585
R227 B.n132 B.n131 585
R228 B.n133 B.n132 585
R229 B.n450 B.n449 585
R230 B.n451 B.n450 585
R231 B.n448 B.n138 585
R232 B.n138 B.n137 585
R233 B.n447 B.n446 585
R234 B.n446 B.n445 585
R235 B.n140 B.n139 585
R236 B.n141 B.n140 585
R237 B.n438 B.n437 585
R238 B.n439 B.n438 585
R239 B.n436 B.n146 585
R240 B.n146 B.n145 585
R241 B.n435 B.n434 585
R242 B.n434 B.n433 585
R243 B.n148 B.n147 585
R244 B.n426 B.n148 585
R245 B.n425 B.n424 585
R246 B.n427 B.n425 585
R247 B.n423 B.n153 585
R248 B.n153 B.n152 585
R249 B.n422 B.n421 585
R250 B.n421 B.n420 585
R251 B.n155 B.n154 585
R252 B.n156 B.n155 585
R253 B.n413 B.n412 585
R254 B.n414 B.n413 585
R255 B.n411 B.n161 585
R256 B.n161 B.n160 585
R257 B.n410 B.n409 585
R258 B.n409 B.n408 585
R259 B.n163 B.n162 585
R260 B.n164 B.n163 585
R261 B.n401 B.n400 585
R262 B.n402 B.n401 585
R263 B.n399 B.n169 585
R264 B.n169 B.n168 585
R265 B.n398 B.n397 585
R266 B.n397 B.n396 585
R267 B.n171 B.n170 585
R268 B.n172 B.n171 585
R269 B.n389 B.n388 585
R270 B.n390 B.n389 585
R271 B.n387 B.n176 585
R272 B.n180 B.n176 585
R273 B.n386 B.n385 585
R274 B.n385 B.n384 585
R275 B.n178 B.n177 585
R276 B.n179 B.n178 585
R277 B.n377 B.n376 585
R278 B.n378 B.n377 585
R279 B.n375 B.n185 585
R280 B.n185 B.n184 585
R281 B.n374 B.n373 585
R282 B.n373 B.n372 585
R283 B.n187 B.n186 585
R284 B.n188 B.n187 585
R285 B.n365 B.n364 585
R286 B.n366 B.n365 585
R287 B.n363 B.n193 585
R288 B.n193 B.n192 585
R289 B.n362 B.n361 585
R290 B.n361 B.n360 585
R291 B.n357 B.n197 585
R292 B.n356 B.n355 585
R293 B.n353 B.n198 585
R294 B.n353 B.n196 585
R295 B.n352 B.n351 585
R296 B.n350 B.n349 585
R297 B.n348 B.n200 585
R298 B.n346 B.n345 585
R299 B.n344 B.n201 585
R300 B.n343 B.n342 585
R301 B.n340 B.n202 585
R302 B.n338 B.n337 585
R303 B.n336 B.n203 585
R304 B.n335 B.n334 585
R305 B.n332 B.n204 585
R306 B.n330 B.n329 585
R307 B.n328 B.n205 585
R308 B.n327 B.n326 585
R309 B.n324 B.n206 585
R310 B.n322 B.n321 585
R311 B.n320 B.n207 585
R312 B.n319 B.n318 585
R313 B.n316 B.n208 585
R314 B.n314 B.n313 585
R315 B.n312 B.n209 585
R316 B.n311 B.n310 585
R317 B.n308 B.n210 585
R318 B.n306 B.n305 585
R319 B.n303 B.n211 585
R320 B.n302 B.n301 585
R321 B.n299 B.n214 585
R322 B.n297 B.n296 585
R323 B.n295 B.n215 585
R324 B.n294 B.n293 585
R325 B.n291 B.n216 585
R326 B.n289 B.n288 585
R327 B.n287 B.n217 585
R328 B.n285 B.n284 585
R329 B.n282 B.n220 585
R330 B.n280 B.n279 585
R331 B.n278 B.n221 585
R332 B.n277 B.n276 585
R333 B.n274 B.n222 585
R334 B.n272 B.n271 585
R335 B.n270 B.n223 585
R336 B.n269 B.n268 585
R337 B.n266 B.n224 585
R338 B.n264 B.n263 585
R339 B.n262 B.n225 585
R340 B.n261 B.n260 585
R341 B.n258 B.n226 585
R342 B.n256 B.n255 585
R343 B.n254 B.n227 585
R344 B.n253 B.n252 585
R345 B.n250 B.n228 585
R346 B.n248 B.n247 585
R347 B.n246 B.n229 585
R348 B.n245 B.n244 585
R349 B.n242 B.n230 585
R350 B.n240 B.n239 585
R351 B.n238 B.n231 585
R352 B.n237 B.n236 585
R353 B.n234 B.n232 585
R354 B.n195 B.n194 585
R355 B.n359 B.n358 585
R356 B.n360 B.n359 585
R357 B.n191 B.n190 585
R358 B.n192 B.n191 585
R359 B.n368 B.n367 585
R360 B.n367 B.n366 585
R361 B.n369 B.n189 585
R362 B.n189 B.n188 585
R363 B.n371 B.n370 585
R364 B.n372 B.n371 585
R365 B.n183 B.n182 585
R366 B.n184 B.n183 585
R367 B.n380 B.n379 585
R368 B.n379 B.n378 585
R369 B.n381 B.n181 585
R370 B.n181 B.n179 585
R371 B.n383 B.n382 585
R372 B.n384 B.n383 585
R373 B.n175 B.n174 585
R374 B.n180 B.n175 585
R375 B.n392 B.n391 585
R376 B.n391 B.n390 585
R377 B.n393 B.n173 585
R378 B.n173 B.n172 585
R379 B.n395 B.n394 585
R380 B.n396 B.n395 585
R381 B.n167 B.n166 585
R382 B.n168 B.n167 585
R383 B.n404 B.n403 585
R384 B.n403 B.n402 585
R385 B.n405 B.n165 585
R386 B.n165 B.n164 585
R387 B.n407 B.n406 585
R388 B.n408 B.n407 585
R389 B.n159 B.n158 585
R390 B.n160 B.n159 585
R391 B.n416 B.n415 585
R392 B.n415 B.n414 585
R393 B.n417 B.n157 585
R394 B.n157 B.n156 585
R395 B.n419 B.n418 585
R396 B.n420 B.n419 585
R397 B.n151 B.n150 585
R398 B.n152 B.n151 585
R399 B.n429 B.n428 585
R400 B.n428 B.n427 585
R401 B.n430 B.n149 585
R402 B.n426 B.n149 585
R403 B.n432 B.n431 585
R404 B.n433 B.n432 585
R405 B.n144 B.n143 585
R406 B.n145 B.n144 585
R407 B.n441 B.n440 585
R408 B.n440 B.n439 585
R409 B.n442 B.n142 585
R410 B.n142 B.n141 585
R411 B.n444 B.n443 585
R412 B.n445 B.n444 585
R413 B.n136 B.n135 585
R414 B.n137 B.n136 585
R415 B.n453 B.n452 585
R416 B.n452 B.n451 585
R417 B.n454 B.n134 585
R418 B.n134 B.n133 585
R419 B.n456 B.n455 585
R420 B.n457 B.n456 585
R421 B.n128 B.n127 585
R422 B.n129 B.n128 585
R423 B.n465 B.n464 585
R424 B.n464 B.n463 585
R425 B.n466 B.n126 585
R426 B.n126 B.n125 585
R427 B.n468 B.n467 585
R428 B.n469 B.n468 585
R429 B.n120 B.n119 585
R430 B.n121 B.n120 585
R431 B.n478 B.n477 585
R432 B.n477 B.n476 585
R433 B.n479 B.n118 585
R434 B.n118 B.n117 585
R435 B.n481 B.n480 585
R436 B.n482 B.n481 585
R437 B.n2 B.n0 585
R438 B.n4 B.n2 585
R439 B.n3 B.n1 585
R440 B.n749 B.n3 585
R441 B.n747 B.n746 585
R442 B.n748 B.n747 585
R443 B.n745 B.n9 585
R444 B.n9 B.n8 585
R445 B.n744 B.n743 585
R446 B.n743 B.n742 585
R447 B.n11 B.n10 585
R448 B.n741 B.n11 585
R449 B.n739 B.n738 585
R450 B.n740 B.n739 585
R451 B.n737 B.n16 585
R452 B.n16 B.n15 585
R453 B.n736 B.n735 585
R454 B.n735 B.n734 585
R455 B.n18 B.n17 585
R456 B.n733 B.n18 585
R457 B.n731 B.n730 585
R458 B.n732 B.n731 585
R459 B.n729 B.n23 585
R460 B.n23 B.n22 585
R461 B.n728 B.n727 585
R462 B.n727 B.n726 585
R463 B.n25 B.n24 585
R464 B.n725 B.n25 585
R465 B.n723 B.n722 585
R466 B.n724 B.n723 585
R467 B.n721 B.n30 585
R468 B.n30 B.n29 585
R469 B.n720 B.n719 585
R470 B.n719 B.n718 585
R471 B.n32 B.n31 585
R472 B.n717 B.n32 585
R473 B.n715 B.n714 585
R474 B.n716 B.n715 585
R475 B.n713 B.n36 585
R476 B.n39 B.n36 585
R477 B.n712 B.n711 585
R478 B.n711 B.n710 585
R479 B.n38 B.n37 585
R480 B.n709 B.n38 585
R481 B.n707 B.n706 585
R482 B.n708 B.n707 585
R483 B.n705 B.n44 585
R484 B.n44 B.n43 585
R485 B.n704 B.n703 585
R486 B.n703 B.n702 585
R487 B.n46 B.n45 585
R488 B.n701 B.n46 585
R489 B.n699 B.n698 585
R490 B.n700 B.n699 585
R491 B.n697 B.n51 585
R492 B.n51 B.n50 585
R493 B.n696 B.n695 585
R494 B.n695 B.n694 585
R495 B.n53 B.n52 585
R496 B.n693 B.n53 585
R497 B.n691 B.n690 585
R498 B.n692 B.n691 585
R499 B.n689 B.n58 585
R500 B.n58 B.n57 585
R501 B.n688 B.n687 585
R502 B.n687 B.n686 585
R503 B.n60 B.n59 585
R504 B.n685 B.n60 585
R505 B.n683 B.n682 585
R506 B.n684 B.n683 585
R507 B.n681 B.n65 585
R508 B.n65 B.n64 585
R509 B.n680 B.n679 585
R510 B.n679 B.n678 585
R511 B.n67 B.n66 585
R512 B.n677 B.n67 585
R513 B.n675 B.n674 585
R514 B.n676 B.n675 585
R515 B.n673 B.n72 585
R516 B.n72 B.n71 585
R517 B.n672 B.n671 585
R518 B.n671 B.n670 585
R519 B.n74 B.n73 585
R520 B.n669 B.n74 585
R521 B.n667 B.n666 585
R522 B.n668 B.n667 585
R523 B.n752 B.n751 585
R524 B.n751 B.n750 585
R525 B.n359 B.n197 492.5
R526 B.n667 B.n79 492.5
R527 B.n361 B.n195 492.5
R528 B.n540 B.n77 492.5
R529 B.n218 B.t15 256.95
R530 B.n212 B.t11 256.95
R531 B.n94 B.t8 256.95
R532 B.n101 B.t4 256.95
R533 B.n541 B.n78 256.663
R534 B.n547 B.n78 256.663
R535 B.n549 B.n78 256.663
R536 B.n555 B.n78 256.663
R537 B.n557 B.n78 256.663
R538 B.n563 B.n78 256.663
R539 B.n565 B.n78 256.663
R540 B.n571 B.n78 256.663
R541 B.n573 B.n78 256.663
R542 B.n579 B.n78 256.663
R543 B.n581 B.n78 256.663
R544 B.n587 B.n78 256.663
R545 B.n589 B.n78 256.663
R546 B.n596 B.n78 256.663
R547 B.n598 B.n78 256.663
R548 B.n604 B.n78 256.663
R549 B.n606 B.n78 256.663
R550 B.n612 B.n78 256.663
R551 B.n614 B.n78 256.663
R552 B.n620 B.n78 256.663
R553 B.n622 B.n78 256.663
R554 B.n628 B.n78 256.663
R555 B.n630 B.n78 256.663
R556 B.n636 B.n78 256.663
R557 B.n638 B.n78 256.663
R558 B.n644 B.n78 256.663
R559 B.n646 B.n78 256.663
R560 B.n652 B.n78 256.663
R561 B.n654 B.n78 256.663
R562 B.n660 B.n78 256.663
R563 B.n662 B.n78 256.663
R564 B.n354 B.n196 256.663
R565 B.n199 B.n196 256.663
R566 B.n347 B.n196 256.663
R567 B.n341 B.n196 256.663
R568 B.n339 B.n196 256.663
R569 B.n333 B.n196 256.663
R570 B.n331 B.n196 256.663
R571 B.n325 B.n196 256.663
R572 B.n323 B.n196 256.663
R573 B.n317 B.n196 256.663
R574 B.n315 B.n196 256.663
R575 B.n309 B.n196 256.663
R576 B.n307 B.n196 256.663
R577 B.n300 B.n196 256.663
R578 B.n298 B.n196 256.663
R579 B.n292 B.n196 256.663
R580 B.n290 B.n196 256.663
R581 B.n283 B.n196 256.663
R582 B.n281 B.n196 256.663
R583 B.n275 B.n196 256.663
R584 B.n273 B.n196 256.663
R585 B.n267 B.n196 256.663
R586 B.n265 B.n196 256.663
R587 B.n259 B.n196 256.663
R588 B.n257 B.n196 256.663
R589 B.n251 B.n196 256.663
R590 B.n249 B.n196 256.663
R591 B.n243 B.n196 256.663
R592 B.n241 B.n196 256.663
R593 B.n235 B.n196 256.663
R594 B.n233 B.n196 256.663
R595 B.n359 B.n191 163.367
R596 B.n367 B.n191 163.367
R597 B.n367 B.n189 163.367
R598 B.n371 B.n189 163.367
R599 B.n371 B.n183 163.367
R600 B.n379 B.n183 163.367
R601 B.n379 B.n181 163.367
R602 B.n383 B.n181 163.367
R603 B.n383 B.n175 163.367
R604 B.n391 B.n175 163.367
R605 B.n391 B.n173 163.367
R606 B.n395 B.n173 163.367
R607 B.n395 B.n167 163.367
R608 B.n403 B.n167 163.367
R609 B.n403 B.n165 163.367
R610 B.n407 B.n165 163.367
R611 B.n407 B.n159 163.367
R612 B.n415 B.n159 163.367
R613 B.n415 B.n157 163.367
R614 B.n419 B.n157 163.367
R615 B.n419 B.n151 163.367
R616 B.n428 B.n151 163.367
R617 B.n428 B.n149 163.367
R618 B.n432 B.n149 163.367
R619 B.n432 B.n144 163.367
R620 B.n440 B.n144 163.367
R621 B.n440 B.n142 163.367
R622 B.n444 B.n142 163.367
R623 B.n444 B.n136 163.367
R624 B.n452 B.n136 163.367
R625 B.n452 B.n134 163.367
R626 B.n456 B.n134 163.367
R627 B.n456 B.n128 163.367
R628 B.n464 B.n128 163.367
R629 B.n464 B.n126 163.367
R630 B.n468 B.n126 163.367
R631 B.n468 B.n120 163.367
R632 B.n477 B.n120 163.367
R633 B.n477 B.n118 163.367
R634 B.n481 B.n118 163.367
R635 B.n481 B.n2 163.367
R636 B.n751 B.n2 163.367
R637 B.n751 B.n3 163.367
R638 B.n747 B.n3 163.367
R639 B.n747 B.n9 163.367
R640 B.n743 B.n9 163.367
R641 B.n743 B.n11 163.367
R642 B.n739 B.n11 163.367
R643 B.n739 B.n16 163.367
R644 B.n735 B.n16 163.367
R645 B.n735 B.n18 163.367
R646 B.n731 B.n18 163.367
R647 B.n731 B.n23 163.367
R648 B.n727 B.n23 163.367
R649 B.n727 B.n25 163.367
R650 B.n723 B.n25 163.367
R651 B.n723 B.n30 163.367
R652 B.n719 B.n30 163.367
R653 B.n719 B.n32 163.367
R654 B.n715 B.n32 163.367
R655 B.n715 B.n36 163.367
R656 B.n711 B.n36 163.367
R657 B.n711 B.n38 163.367
R658 B.n707 B.n38 163.367
R659 B.n707 B.n44 163.367
R660 B.n703 B.n44 163.367
R661 B.n703 B.n46 163.367
R662 B.n699 B.n46 163.367
R663 B.n699 B.n51 163.367
R664 B.n695 B.n51 163.367
R665 B.n695 B.n53 163.367
R666 B.n691 B.n53 163.367
R667 B.n691 B.n58 163.367
R668 B.n687 B.n58 163.367
R669 B.n687 B.n60 163.367
R670 B.n683 B.n60 163.367
R671 B.n683 B.n65 163.367
R672 B.n679 B.n65 163.367
R673 B.n679 B.n67 163.367
R674 B.n675 B.n67 163.367
R675 B.n675 B.n72 163.367
R676 B.n671 B.n72 163.367
R677 B.n671 B.n74 163.367
R678 B.n667 B.n74 163.367
R679 B.n355 B.n353 163.367
R680 B.n353 B.n352 163.367
R681 B.n349 B.n348 163.367
R682 B.n346 B.n201 163.367
R683 B.n342 B.n340 163.367
R684 B.n338 B.n203 163.367
R685 B.n334 B.n332 163.367
R686 B.n330 B.n205 163.367
R687 B.n326 B.n324 163.367
R688 B.n322 B.n207 163.367
R689 B.n318 B.n316 163.367
R690 B.n314 B.n209 163.367
R691 B.n310 B.n308 163.367
R692 B.n306 B.n211 163.367
R693 B.n301 B.n299 163.367
R694 B.n297 B.n215 163.367
R695 B.n293 B.n291 163.367
R696 B.n289 B.n217 163.367
R697 B.n284 B.n282 163.367
R698 B.n280 B.n221 163.367
R699 B.n276 B.n274 163.367
R700 B.n272 B.n223 163.367
R701 B.n268 B.n266 163.367
R702 B.n264 B.n225 163.367
R703 B.n260 B.n258 163.367
R704 B.n256 B.n227 163.367
R705 B.n252 B.n250 163.367
R706 B.n248 B.n229 163.367
R707 B.n244 B.n242 163.367
R708 B.n240 B.n231 163.367
R709 B.n236 B.n234 163.367
R710 B.n361 B.n193 163.367
R711 B.n365 B.n193 163.367
R712 B.n365 B.n187 163.367
R713 B.n373 B.n187 163.367
R714 B.n373 B.n185 163.367
R715 B.n377 B.n185 163.367
R716 B.n377 B.n178 163.367
R717 B.n385 B.n178 163.367
R718 B.n385 B.n176 163.367
R719 B.n389 B.n176 163.367
R720 B.n389 B.n171 163.367
R721 B.n397 B.n171 163.367
R722 B.n397 B.n169 163.367
R723 B.n401 B.n169 163.367
R724 B.n401 B.n163 163.367
R725 B.n409 B.n163 163.367
R726 B.n409 B.n161 163.367
R727 B.n413 B.n161 163.367
R728 B.n413 B.n155 163.367
R729 B.n421 B.n155 163.367
R730 B.n421 B.n153 163.367
R731 B.n425 B.n153 163.367
R732 B.n425 B.n148 163.367
R733 B.n434 B.n148 163.367
R734 B.n434 B.n146 163.367
R735 B.n438 B.n146 163.367
R736 B.n438 B.n140 163.367
R737 B.n446 B.n140 163.367
R738 B.n446 B.n138 163.367
R739 B.n450 B.n138 163.367
R740 B.n450 B.n132 163.367
R741 B.n458 B.n132 163.367
R742 B.n458 B.n130 163.367
R743 B.n462 B.n130 163.367
R744 B.n462 B.n124 163.367
R745 B.n470 B.n124 163.367
R746 B.n470 B.n122 163.367
R747 B.n475 B.n122 163.367
R748 B.n475 B.n116 163.367
R749 B.n483 B.n116 163.367
R750 B.n484 B.n483 163.367
R751 B.n484 B.n5 163.367
R752 B.n6 B.n5 163.367
R753 B.n7 B.n6 163.367
R754 B.n489 B.n7 163.367
R755 B.n489 B.n12 163.367
R756 B.n13 B.n12 163.367
R757 B.n14 B.n13 163.367
R758 B.n494 B.n14 163.367
R759 B.n494 B.n19 163.367
R760 B.n20 B.n19 163.367
R761 B.n21 B.n20 163.367
R762 B.n499 B.n21 163.367
R763 B.n499 B.n26 163.367
R764 B.n27 B.n26 163.367
R765 B.n28 B.n27 163.367
R766 B.n504 B.n28 163.367
R767 B.n504 B.n33 163.367
R768 B.n34 B.n33 163.367
R769 B.n35 B.n34 163.367
R770 B.n509 B.n35 163.367
R771 B.n509 B.n40 163.367
R772 B.n41 B.n40 163.367
R773 B.n42 B.n41 163.367
R774 B.n514 B.n42 163.367
R775 B.n514 B.n47 163.367
R776 B.n48 B.n47 163.367
R777 B.n49 B.n48 163.367
R778 B.n519 B.n49 163.367
R779 B.n519 B.n54 163.367
R780 B.n55 B.n54 163.367
R781 B.n56 B.n55 163.367
R782 B.n524 B.n56 163.367
R783 B.n524 B.n61 163.367
R784 B.n62 B.n61 163.367
R785 B.n63 B.n62 163.367
R786 B.n529 B.n63 163.367
R787 B.n529 B.n68 163.367
R788 B.n69 B.n68 163.367
R789 B.n70 B.n69 163.367
R790 B.n534 B.n70 163.367
R791 B.n534 B.n75 163.367
R792 B.n76 B.n75 163.367
R793 B.n77 B.n76 163.367
R794 B.n663 B.n661 163.367
R795 B.n659 B.n81 163.367
R796 B.n655 B.n653 163.367
R797 B.n651 B.n83 163.367
R798 B.n647 B.n645 163.367
R799 B.n643 B.n85 163.367
R800 B.n639 B.n637 163.367
R801 B.n635 B.n87 163.367
R802 B.n631 B.n629 163.367
R803 B.n627 B.n89 163.367
R804 B.n623 B.n621 163.367
R805 B.n619 B.n91 163.367
R806 B.n615 B.n613 163.367
R807 B.n611 B.n93 163.367
R808 B.n607 B.n605 163.367
R809 B.n603 B.n98 163.367
R810 B.n599 B.n597 163.367
R811 B.n595 B.n100 163.367
R812 B.n590 B.n588 163.367
R813 B.n586 B.n104 163.367
R814 B.n582 B.n580 163.367
R815 B.n578 B.n106 163.367
R816 B.n574 B.n572 163.367
R817 B.n570 B.n108 163.367
R818 B.n566 B.n564 163.367
R819 B.n562 B.n110 163.367
R820 B.n558 B.n556 163.367
R821 B.n554 B.n112 163.367
R822 B.n550 B.n548 163.367
R823 B.n546 B.n114 163.367
R824 B.n542 B.n540 163.367
R825 B.n218 B.t17 146.173
R826 B.n101 B.t6 146.173
R827 B.n212 B.t14 146.166
R828 B.n94 B.t9 146.166
R829 B.n360 B.n196 105.276
R830 B.n668 B.n78 105.276
R831 B.n219 B.n218 74.2793
R832 B.n213 B.n212 74.2793
R833 B.n95 B.n94 74.2793
R834 B.n102 B.n101 74.2793
R835 B.n219 B.t16 71.8945
R836 B.n102 B.t7 71.8945
R837 B.n213 B.t13 71.8867
R838 B.n95 B.t10 71.8867
R839 B.n354 B.n197 71.676
R840 B.n352 B.n199 71.676
R841 B.n348 B.n347 71.676
R842 B.n341 B.n201 71.676
R843 B.n340 B.n339 71.676
R844 B.n333 B.n203 71.676
R845 B.n332 B.n331 71.676
R846 B.n325 B.n205 71.676
R847 B.n324 B.n323 71.676
R848 B.n317 B.n207 71.676
R849 B.n316 B.n315 71.676
R850 B.n309 B.n209 71.676
R851 B.n308 B.n307 71.676
R852 B.n300 B.n211 71.676
R853 B.n299 B.n298 71.676
R854 B.n292 B.n215 71.676
R855 B.n291 B.n290 71.676
R856 B.n283 B.n217 71.676
R857 B.n282 B.n281 71.676
R858 B.n275 B.n221 71.676
R859 B.n274 B.n273 71.676
R860 B.n267 B.n223 71.676
R861 B.n266 B.n265 71.676
R862 B.n259 B.n225 71.676
R863 B.n258 B.n257 71.676
R864 B.n251 B.n227 71.676
R865 B.n250 B.n249 71.676
R866 B.n243 B.n229 71.676
R867 B.n242 B.n241 71.676
R868 B.n235 B.n231 71.676
R869 B.n234 B.n233 71.676
R870 B.n662 B.n79 71.676
R871 B.n661 B.n660 71.676
R872 B.n654 B.n81 71.676
R873 B.n653 B.n652 71.676
R874 B.n646 B.n83 71.676
R875 B.n645 B.n644 71.676
R876 B.n638 B.n85 71.676
R877 B.n637 B.n636 71.676
R878 B.n630 B.n87 71.676
R879 B.n629 B.n628 71.676
R880 B.n622 B.n89 71.676
R881 B.n621 B.n620 71.676
R882 B.n614 B.n91 71.676
R883 B.n613 B.n612 71.676
R884 B.n606 B.n93 71.676
R885 B.n605 B.n604 71.676
R886 B.n598 B.n98 71.676
R887 B.n597 B.n596 71.676
R888 B.n589 B.n100 71.676
R889 B.n588 B.n587 71.676
R890 B.n581 B.n104 71.676
R891 B.n580 B.n579 71.676
R892 B.n573 B.n106 71.676
R893 B.n572 B.n571 71.676
R894 B.n565 B.n108 71.676
R895 B.n564 B.n563 71.676
R896 B.n557 B.n110 71.676
R897 B.n556 B.n555 71.676
R898 B.n549 B.n112 71.676
R899 B.n548 B.n547 71.676
R900 B.n541 B.n114 71.676
R901 B.n542 B.n541 71.676
R902 B.n547 B.n546 71.676
R903 B.n550 B.n549 71.676
R904 B.n555 B.n554 71.676
R905 B.n558 B.n557 71.676
R906 B.n563 B.n562 71.676
R907 B.n566 B.n565 71.676
R908 B.n571 B.n570 71.676
R909 B.n574 B.n573 71.676
R910 B.n579 B.n578 71.676
R911 B.n582 B.n581 71.676
R912 B.n587 B.n586 71.676
R913 B.n590 B.n589 71.676
R914 B.n596 B.n595 71.676
R915 B.n599 B.n598 71.676
R916 B.n604 B.n603 71.676
R917 B.n607 B.n606 71.676
R918 B.n612 B.n611 71.676
R919 B.n615 B.n614 71.676
R920 B.n620 B.n619 71.676
R921 B.n623 B.n622 71.676
R922 B.n628 B.n627 71.676
R923 B.n631 B.n630 71.676
R924 B.n636 B.n635 71.676
R925 B.n639 B.n638 71.676
R926 B.n644 B.n643 71.676
R927 B.n647 B.n646 71.676
R928 B.n652 B.n651 71.676
R929 B.n655 B.n654 71.676
R930 B.n660 B.n659 71.676
R931 B.n663 B.n662 71.676
R932 B.n355 B.n354 71.676
R933 B.n349 B.n199 71.676
R934 B.n347 B.n346 71.676
R935 B.n342 B.n341 71.676
R936 B.n339 B.n338 71.676
R937 B.n334 B.n333 71.676
R938 B.n331 B.n330 71.676
R939 B.n326 B.n325 71.676
R940 B.n323 B.n322 71.676
R941 B.n318 B.n317 71.676
R942 B.n315 B.n314 71.676
R943 B.n310 B.n309 71.676
R944 B.n307 B.n306 71.676
R945 B.n301 B.n300 71.676
R946 B.n298 B.n297 71.676
R947 B.n293 B.n292 71.676
R948 B.n290 B.n289 71.676
R949 B.n284 B.n283 71.676
R950 B.n281 B.n280 71.676
R951 B.n276 B.n275 71.676
R952 B.n273 B.n272 71.676
R953 B.n268 B.n267 71.676
R954 B.n265 B.n264 71.676
R955 B.n260 B.n259 71.676
R956 B.n257 B.n256 71.676
R957 B.n252 B.n251 71.676
R958 B.n249 B.n248 71.676
R959 B.n244 B.n243 71.676
R960 B.n241 B.n240 71.676
R961 B.n236 B.n235 71.676
R962 B.n233 B.n195 71.676
R963 B.n360 B.n192 61.1866
R964 B.n366 B.n192 61.1866
R965 B.n366 B.n188 61.1866
R966 B.n372 B.n188 61.1866
R967 B.n372 B.n184 61.1866
R968 B.n378 B.n184 61.1866
R969 B.n378 B.n179 61.1866
R970 B.n384 B.n179 61.1866
R971 B.n384 B.n180 61.1866
R972 B.n390 B.n172 61.1866
R973 B.n396 B.n172 61.1866
R974 B.n396 B.n168 61.1866
R975 B.n402 B.n168 61.1866
R976 B.n402 B.n164 61.1866
R977 B.n408 B.n164 61.1866
R978 B.n408 B.n160 61.1866
R979 B.n414 B.n160 61.1866
R980 B.n414 B.n156 61.1866
R981 B.n420 B.n156 61.1866
R982 B.n420 B.n152 61.1866
R983 B.n427 B.n152 61.1866
R984 B.n427 B.n426 61.1866
R985 B.n433 B.n145 61.1866
R986 B.n439 B.n145 61.1866
R987 B.n439 B.n141 61.1866
R988 B.n445 B.n141 61.1866
R989 B.n445 B.n137 61.1866
R990 B.n451 B.n137 61.1866
R991 B.n451 B.n133 61.1866
R992 B.n457 B.n133 61.1866
R993 B.n457 B.n129 61.1866
R994 B.n463 B.n129 61.1866
R995 B.n469 B.n125 61.1866
R996 B.n469 B.n121 61.1866
R997 B.n476 B.n121 61.1866
R998 B.n476 B.n117 61.1866
R999 B.n482 B.n117 61.1866
R1000 B.n482 B.n4 61.1866
R1001 B.n750 B.n4 61.1866
R1002 B.n750 B.n749 61.1866
R1003 B.n749 B.n748 61.1866
R1004 B.n748 B.n8 61.1866
R1005 B.n742 B.n8 61.1866
R1006 B.n742 B.n741 61.1866
R1007 B.n741 B.n740 61.1866
R1008 B.n740 B.n15 61.1866
R1009 B.n734 B.n733 61.1866
R1010 B.n733 B.n732 61.1866
R1011 B.n732 B.n22 61.1866
R1012 B.n726 B.n22 61.1866
R1013 B.n726 B.n725 61.1866
R1014 B.n725 B.n724 61.1866
R1015 B.n724 B.n29 61.1866
R1016 B.n718 B.n29 61.1866
R1017 B.n718 B.n717 61.1866
R1018 B.n717 B.n716 61.1866
R1019 B.n710 B.n39 61.1866
R1020 B.n710 B.n709 61.1866
R1021 B.n709 B.n708 61.1866
R1022 B.n708 B.n43 61.1866
R1023 B.n702 B.n43 61.1866
R1024 B.n702 B.n701 61.1866
R1025 B.n701 B.n700 61.1866
R1026 B.n700 B.n50 61.1866
R1027 B.n694 B.n50 61.1866
R1028 B.n694 B.n693 61.1866
R1029 B.n693 B.n692 61.1866
R1030 B.n692 B.n57 61.1866
R1031 B.n686 B.n57 61.1866
R1032 B.n685 B.n684 61.1866
R1033 B.n684 B.n64 61.1866
R1034 B.n678 B.n64 61.1866
R1035 B.n678 B.n677 61.1866
R1036 B.n677 B.n676 61.1866
R1037 B.n676 B.n71 61.1866
R1038 B.n670 B.n71 61.1866
R1039 B.n670 B.n669 61.1866
R1040 B.n669 B.n668 61.1866
R1041 B.n286 B.n219 59.5399
R1042 B.n304 B.n213 59.5399
R1043 B.n96 B.n95 59.5399
R1044 B.n593 B.n102 59.5399
R1045 B.n390 B.t12 59.387
R1046 B.n686 B.t5 59.387
R1047 B.n463 B.t2 46.7899
R1048 B.n734 B.t3 46.7899
R1049 B.n666 B.n665 32.0005
R1050 B.n539 B.n538 32.0005
R1051 B.n362 B.n194 32.0005
R1052 B.n358 B.n357 32.0005
R1053 B.n426 B.t1 30.5935
R1054 B.n433 B.t1 30.5935
R1055 B.n716 B.t0 30.5935
R1056 B.n39 B.t0 30.5935
R1057 B B.n752 18.0485
R1058 B.t2 B.n125 14.3972
R1059 B.t3 B.n15 14.3972
R1060 B.n665 B.n664 10.6151
R1061 B.n664 B.n80 10.6151
R1062 B.n658 B.n80 10.6151
R1063 B.n658 B.n657 10.6151
R1064 B.n657 B.n656 10.6151
R1065 B.n656 B.n82 10.6151
R1066 B.n650 B.n82 10.6151
R1067 B.n650 B.n649 10.6151
R1068 B.n649 B.n648 10.6151
R1069 B.n648 B.n84 10.6151
R1070 B.n642 B.n84 10.6151
R1071 B.n642 B.n641 10.6151
R1072 B.n641 B.n640 10.6151
R1073 B.n640 B.n86 10.6151
R1074 B.n634 B.n86 10.6151
R1075 B.n634 B.n633 10.6151
R1076 B.n633 B.n632 10.6151
R1077 B.n632 B.n88 10.6151
R1078 B.n626 B.n88 10.6151
R1079 B.n626 B.n625 10.6151
R1080 B.n625 B.n624 10.6151
R1081 B.n624 B.n90 10.6151
R1082 B.n618 B.n90 10.6151
R1083 B.n618 B.n617 10.6151
R1084 B.n617 B.n616 10.6151
R1085 B.n616 B.n92 10.6151
R1086 B.n610 B.n609 10.6151
R1087 B.n609 B.n608 10.6151
R1088 B.n608 B.n97 10.6151
R1089 B.n602 B.n97 10.6151
R1090 B.n602 B.n601 10.6151
R1091 B.n601 B.n600 10.6151
R1092 B.n600 B.n99 10.6151
R1093 B.n594 B.n99 10.6151
R1094 B.n592 B.n591 10.6151
R1095 B.n591 B.n103 10.6151
R1096 B.n585 B.n103 10.6151
R1097 B.n585 B.n584 10.6151
R1098 B.n584 B.n583 10.6151
R1099 B.n583 B.n105 10.6151
R1100 B.n577 B.n105 10.6151
R1101 B.n577 B.n576 10.6151
R1102 B.n576 B.n575 10.6151
R1103 B.n575 B.n107 10.6151
R1104 B.n569 B.n107 10.6151
R1105 B.n569 B.n568 10.6151
R1106 B.n568 B.n567 10.6151
R1107 B.n567 B.n109 10.6151
R1108 B.n561 B.n109 10.6151
R1109 B.n561 B.n560 10.6151
R1110 B.n560 B.n559 10.6151
R1111 B.n559 B.n111 10.6151
R1112 B.n553 B.n111 10.6151
R1113 B.n553 B.n552 10.6151
R1114 B.n552 B.n551 10.6151
R1115 B.n551 B.n113 10.6151
R1116 B.n545 B.n113 10.6151
R1117 B.n545 B.n544 10.6151
R1118 B.n544 B.n543 10.6151
R1119 B.n543 B.n539 10.6151
R1120 B.n363 B.n362 10.6151
R1121 B.n364 B.n363 10.6151
R1122 B.n364 B.n186 10.6151
R1123 B.n374 B.n186 10.6151
R1124 B.n375 B.n374 10.6151
R1125 B.n376 B.n375 10.6151
R1126 B.n376 B.n177 10.6151
R1127 B.n386 B.n177 10.6151
R1128 B.n387 B.n386 10.6151
R1129 B.n388 B.n387 10.6151
R1130 B.n388 B.n170 10.6151
R1131 B.n398 B.n170 10.6151
R1132 B.n399 B.n398 10.6151
R1133 B.n400 B.n399 10.6151
R1134 B.n400 B.n162 10.6151
R1135 B.n410 B.n162 10.6151
R1136 B.n411 B.n410 10.6151
R1137 B.n412 B.n411 10.6151
R1138 B.n412 B.n154 10.6151
R1139 B.n422 B.n154 10.6151
R1140 B.n423 B.n422 10.6151
R1141 B.n424 B.n423 10.6151
R1142 B.n424 B.n147 10.6151
R1143 B.n435 B.n147 10.6151
R1144 B.n436 B.n435 10.6151
R1145 B.n437 B.n436 10.6151
R1146 B.n437 B.n139 10.6151
R1147 B.n447 B.n139 10.6151
R1148 B.n448 B.n447 10.6151
R1149 B.n449 B.n448 10.6151
R1150 B.n449 B.n131 10.6151
R1151 B.n459 B.n131 10.6151
R1152 B.n460 B.n459 10.6151
R1153 B.n461 B.n460 10.6151
R1154 B.n461 B.n123 10.6151
R1155 B.n471 B.n123 10.6151
R1156 B.n472 B.n471 10.6151
R1157 B.n474 B.n472 10.6151
R1158 B.n474 B.n473 10.6151
R1159 B.n473 B.n115 10.6151
R1160 B.n485 B.n115 10.6151
R1161 B.n486 B.n485 10.6151
R1162 B.n487 B.n486 10.6151
R1163 B.n488 B.n487 10.6151
R1164 B.n490 B.n488 10.6151
R1165 B.n491 B.n490 10.6151
R1166 B.n492 B.n491 10.6151
R1167 B.n493 B.n492 10.6151
R1168 B.n495 B.n493 10.6151
R1169 B.n496 B.n495 10.6151
R1170 B.n497 B.n496 10.6151
R1171 B.n498 B.n497 10.6151
R1172 B.n500 B.n498 10.6151
R1173 B.n501 B.n500 10.6151
R1174 B.n502 B.n501 10.6151
R1175 B.n503 B.n502 10.6151
R1176 B.n505 B.n503 10.6151
R1177 B.n506 B.n505 10.6151
R1178 B.n507 B.n506 10.6151
R1179 B.n508 B.n507 10.6151
R1180 B.n510 B.n508 10.6151
R1181 B.n511 B.n510 10.6151
R1182 B.n512 B.n511 10.6151
R1183 B.n513 B.n512 10.6151
R1184 B.n515 B.n513 10.6151
R1185 B.n516 B.n515 10.6151
R1186 B.n517 B.n516 10.6151
R1187 B.n518 B.n517 10.6151
R1188 B.n520 B.n518 10.6151
R1189 B.n521 B.n520 10.6151
R1190 B.n522 B.n521 10.6151
R1191 B.n523 B.n522 10.6151
R1192 B.n525 B.n523 10.6151
R1193 B.n526 B.n525 10.6151
R1194 B.n527 B.n526 10.6151
R1195 B.n528 B.n527 10.6151
R1196 B.n530 B.n528 10.6151
R1197 B.n531 B.n530 10.6151
R1198 B.n532 B.n531 10.6151
R1199 B.n533 B.n532 10.6151
R1200 B.n535 B.n533 10.6151
R1201 B.n536 B.n535 10.6151
R1202 B.n537 B.n536 10.6151
R1203 B.n538 B.n537 10.6151
R1204 B.n357 B.n356 10.6151
R1205 B.n356 B.n198 10.6151
R1206 B.n351 B.n198 10.6151
R1207 B.n351 B.n350 10.6151
R1208 B.n350 B.n200 10.6151
R1209 B.n345 B.n200 10.6151
R1210 B.n345 B.n344 10.6151
R1211 B.n344 B.n343 10.6151
R1212 B.n343 B.n202 10.6151
R1213 B.n337 B.n202 10.6151
R1214 B.n337 B.n336 10.6151
R1215 B.n336 B.n335 10.6151
R1216 B.n335 B.n204 10.6151
R1217 B.n329 B.n204 10.6151
R1218 B.n329 B.n328 10.6151
R1219 B.n328 B.n327 10.6151
R1220 B.n327 B.n206 10.6151
R1221 B.n321 B.n206 10.6151
R1222 B.n321 B.n320 10.6151
R1223 B.n320 B.n319 10.6151
R1224 B.n319 B.n208 10.6151
R1225 B.n313 B.n208 10.6151
R1226 B.n313 B.n312 10.6151
R1227 B.n312 B.n311 10.6151
R1228 B.n311 B.n210 10.6151
R1229 B.n305 B.n210 10.6151
R1230 B.n303 B.n302 10.6151
R1231 B.n302 B.n214 10.6151
R1232 B.n296 B.n214 10.6151
R1233 B.n296 B.n295 10.6151
R1234 B.n295 B.n294 10.6151
R1235 B.n294 B.n216 10.6151
R1236 B.n288 B.n216 10.6151
R1237 B.n288 B.n287 10.6151
R1238 B.n285 B.n220 10.6151
R1239 B.n279 B.n220 10.6151
R1240 B.n279 B.n278 10.6151
R1241 B.n278 B.n277 10.6151
R1242 B.n277 B.n222 10.6151
R1243 B.n271 B.n222 10.6151
R1244 B.n271 B.n270 10.6151
R1245 B.n270 B.n269 10.6151
R1246 B.n269 B.n224 10.6151
R1247 B.n263 B.n224 10.6151
R1248 B.n263 B.n262 10.6151
R1249 B.n262 B.n261 10.6151
R1250 B.n261 B.n226 10.6151
R1251 B.n255 B.n226 10.6151
R1252 B.n255 B.n254 10.6151
R1253 B.n254 B.n253 10.6151
R1254 B.n253 B.n228 10.6151
R1255 B.n247 B.n228 10.6151
R1256 B.n247 B.n246 10.6151
R1257 B.n246 B.n245 10.6151
R1258 B.n245 B.n230 10.6151
R1259 B.n239 B.n230 10.6151
R1260 B.n239 B.n238 10.6151
R1261 B.n238 B.n237 10.6151
R1262 B.n237 B.n232 10.6151
R1263 B.n232 B.n194 10.6151
R1264 B.n358 B.n190 10.6151
R1265 B.n368 B.n190 10.6151
R1266 B.n369 B.n368 10.6151
R1267 B.n370 B.n369 10.6151
R1268 B.n370 B.n182 10.6151
R1269 B.n380 B.n182 10.6151
R1270 B.n381 B.n380 10.6151
R1271 B.n382 B.n381 10.6151
R1272 B.n382 B.n174 10.6151
R1273 B.n392 B.n174 10.6151
R1274 B.n393 B.n392 10.6151
R1275 B.n394 B.n393 10.6151
R1276 B.n394 B.n166 10.6151
R1277 B.n404 B.n166 10.6151
R1278 B.n405 B.n404 10.6151
R1279 B.n406 B.n405 10.6151
R1280 B.n406 B.n158 10.6151
R1281 B.n416 B.n158 10.6151
R1282 B.n417 B.n416 10.6151
R1283 B.n418 B.n417 10.6151
R1284 B.n418 B.n150 10.6151
R1285 B.n429 B.n150 10.6151
R1286 B.n430 B.n429 10.6151
R1287 B.n431 B.n430 10.6151
R1288 B.n431 B.n143 10.6151
R1289 B.n441 B.n143 10.6151
R1290 B.n442 B.n441 10.6151
R1291 B.n443 B.n442 10.6151
R1292 B.n443 B.n135 10.6151
R1293 B.n453 B.n135 10.6151
R1294 B.n454 B.n453 10.6151
R1295 B.n455 B.n454 10.6151
R1296 B.n455 B.n127 10.6151
R1297 B.n465 B.n127 10.6151
R1298 B.n466 B.n465 10.6151
R1299 B.n467 B.n466 10.6151
R1300 B.n467 B.n119 10.6151
R1301 B.n478 B.n119 10.6151
R1302 B.n479 B.n478 10.6151
R1303 B.n480 B.n479 10.6151
R1304 B.n480 B.n0 10.6151
R1305 B.n746 B.n1 10.6151
R1306 B.n746 B.n745 10.6151
R1307 B.n745 B.n744 10.6151
R1308 B.n744 B.n10 10.6151
R1309 B.n738 B.n10 10.6151
R1310 B.n738 B.n737 10.6151
R1311 B.n737 B.n736 10.6151
R1312 B.n736 B.n17 10.6151
R1313 B.n730 B.n17 10.6151
R1314 B.n730 B.n729 10.6151
R1315 B.n729 B.n728 10.6151
R1316 B.n728 B.n24 10.6151
R1317 B.n722 B.n24 10.6151
R1318 B.n722 B.n721 10.6151
R1319 B.n721 B.n720 10.6151
R1320 B.n720 B.n31 10.6151
R1321 B.n714 B.n31 10.6151
R1322 B.n714 B.n713 10.6151
R1323 B.n713 B.n712 10.6151
R1324 B.n712 B.n37 10.6151
R1325 B.n706 B.n37 10.6151
R1326 B.n706 B.n705 10.6151
R1327 B.n705 B.n704 10.6151
R1328 B.n704 B.n45 10.6151
R1329 B.n698 B.n45 10.6151
R1330 B.n698 B.n697 10.6151
R1331 B.n697 B.n696 10.6151
R1332 B.n696 B.n52 10.6151
R1333 B.n690 B.n52 10.6151
R1334 B.n690 B.n689 10.6151
R1335 B.n689 B.n688 10.6151
R1336 B.n688 B.n59 10.6151
R1337 B.n682 B.n59 10.6151
R1338 B.n682 B.n681 10.6151
R1339 B.n681 B.n680 10.6151
R1340 B.n680 B.n66 10.6151
R1341 B.n674 B.n66 10.6151
R1342 B.n674 B.n673 10.6151
R1343 B.n673 B.n672 10.6151
R1344 B.n672 B.n73 10.6151
R1345 B.n666 B.n73 10.6151
R1346 B.n610 B.n96 6.5566
R1347 B.n594 B.n593 6.5566
R1348 B.n304 B.n303 6.5566
R1349 B.n287 B.n286 6.5566
R1350 B.n96 B.n92 4.05904
R1351 B.n593 B.n592 4.05904
R1352 B.n305 B.n304 4.05904
R1353 B.n286 B.n285 4.05904
R1354 B.n752 B.n0 2.81026
R1355 B.n752 B.n1 2.81026
R1356 B.n180 B.t12 1.80009
R1357 B.t5 B.n685 1.80009
R1358 VN.n0 VN.t3 82.2953
R1359 VN.n1 VN.t2 82.2953
R1360 VN.n1 VN.t1 81.0755
R1361 VN.n0 VN.t0 81.0755
R1362 VN VN.n1 47.6365
R1363 VN VN.n0 2.20088
R1364 VDD2.n2 VDD2.n0 109.091
R1365 VDD2.n2 VDD2.n1 69.4804
R1366 VDD2.n1 VDD2.t2 2.84942
R1367 VDD2.n1 VDD2.t1 2.84942
R1368 VDD2.n0 VDD2.t0 2.84942
R1369 VDD2.n0 VDD2.t3 2.84942
R1370 VDD2 VDD2.n2 0.0586897
C0 VN VDD2 3.01617f
C1 VDD2 VP 0.451724f
C2 VN VTAIL 3.43996f
C3 VP VTAIL 3.45407f
C4 VDD1 VDD2 1.24157f
C5 VDD1 VTAIL 4.5614f
C6 VN VP 5.90642f
C7 VDD2 VTAIL 4.62164f
C8 VN VDD1 0.149964f
C9 VDD1 VP 3.31697f
C10 VDD2 B 3.898477f
C11 VDD1 B 7.94742f
C12 VTAIL B 7.203583f
C13 VN B 11.964861f
C14 VP B 10.360171f
C15 VDD2.t0 B 0.152873f
C16 VDD2.t3 B 0.152873f
C17 VDD2.n0 B 1.8298f
C18 VDD2.t2 B 0.152873f
C19 VDD2.t1 B 0.152873f
C20 VDD2.n1 B 1.30842f
C21 VDD2.n2 B 3.54816f
C22 VN.t0 B 1.81861f
C23 VN.t3 B 1.82917f
C24 VN.n0 B 1.08037f
C25 VN.t2 B 1.82917f
C26 VN.t1 B 1.81861f
C27 VN.n1 B 2.4277f
C28 VDD1.t1 B 0.156787f
C29 VDD1.t3 B 0.156787f
C30 VDD1.n0 B 1.34237f
C31 VDD1.t0 B 0.156787f
C32 VDD1.t2 B 0.156787f
C33 VDD1.n1 B 1.90196f
C34 VTAIL.t3 B 1.12555f
C35 VTAIL.n0 B 0.369093f
C36 VTAIL.t6 B 1.12555f
C37 VTAIL.n1 B 0.470765f
C38 VTAIL.t5 B 1.12555f
C39 VTAIL.n2 B 1.30314f
C40 VTAIL.t1 B 1.12556f
C41 VTAIL.n3 B 1.30313f
C42 VTAIL.t2 B 1.12556f
C43 VTAIL.n4 B 0.470755f
C44 VTAIL.t7 B 1.12556f
C45 VTAIL.n5 B 0.470755f
C46 VTAIL.t4 B 1.12555f
C47 VTAIL.n6 B 1.30314f
C48 VTAIL.t0 B 1.12555f
C49 VTAIL.n7 B 1.19404f
C50 VP.t1 B 1.57471f
C51 VP.n0 B 0.66459f
C52 VP.n1 B 0.024263f
C53 VP.n2 B 0.03542f
C54 VP.n3 B 0.024263f
C55 VP.n4 B 0.030261f
C56 VP.t2 B 1.89373f
C57 VP.t0 B 1.88279f
C58 VP.n5 B 2.50332f
C59 VP.t3 B 1.57471f
C60 VP.n6 B 0.66459f
C61 VP.n7 B 1.29048f
C62 VP.n8 B 0.039161f
C63 VP.n9 B 0.024263f
C64 VP.n10 B 0.045221f
C65 VP.n11 B 0.045221f
C66 VP.n12 B 0.03542f
C67 VP.n13 B 0.024263f
C68 VP.n14 B 0.024263f
C69 VP.n15 B 0.024263f
C70 VP.n16 B 0.045221f
C71 VP.n17 B 0.045221f
C72 VP.n18 B 0.030261f
C73 VP.n19 B 0.039161f
C74 VP.n20 B 0.066765f
.ends

