* NGSPICE file created from diff_pair_sample_1749.ext - technology: sky130A

.subckt diff_pair_sample_1749 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=0.69465 ps=4.54 w=4.21 l=0.71
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=1.6419 ps=9.2 w=4.21 l=0.71
X2 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=1.6419 ps=9.2 w=4.21 l=0.71
X3 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0.69465 ps=4.54 w=4.21 l=0.71
X4 VTAIL.t9 VP.t2 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=0.69465 ps=4.54 w=4.21 l=0.71
X5 VTAIL.t5 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=0.69465 ps=4.54 w=4.21 l=0.71
X6 VDD1.t0 VP.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0.69465 ps=4.54 w=4.21 l=0.71
X7 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0 ps=0 w=4.21 l=0.71
X8 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0.69465 ps=4.54 w=4.21 l=0.71
X9 VDD1.t5 VP.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0.69465 ps=4.54 w=4.21 l=0.71
X10 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0 ps=0 w=4.21 l=0.71
X11 VDD2.t1 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=1.6419 ps=9.2 w=4.21 l=0.71
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0 ps=0 w=4.21 l=0.71
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6419 pd=9.2 as=0 ps=0 w=4.21 l=0.71
X14 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=0.69465 ps=4.54 w=4.21 l=0.71
X15 VDD1.t3 VP.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.69465 pd=4.54 as=1.6419 ps=9.2 w=4.21 l=0.71
R0 VP.n3 VP.t3 220.362
R1 VP.n8 VP.t4 198.571
R2 VP.n12 VP.t0 198.571
R3 VP.n14 VP.t5 198.571
R4 VP.n6 VP.t1 198.571
R5 VP.n4 VP.t2 198.571
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.8565
R14 VP.n9 VP.n7 35.349
R15 VP.n8 VP.n1 27.0217
R16 VP.n14 VP.n13 27.0217
R17 VP.n6 VP.n5 27.0217
R18 VP.n12 VP.n1 21.1793
R19 VP.n13 VP.n12 21.1793
R20 VP.n5 VP.n4 21.1793
R21 VP.n4 VP.n3 20.1275
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VDD1 VDD1.t0 77.5461
R29 VDD1.n1 VDD1.t5 77.4323
R30 VDD1.n1 VDD1.n0 72.281
R31 VDD1.n3 VDD1.n2 72.1122
R32 VDD1.n3 VDD1.n1 31.2897
R33 VDD1.n2 VDD1.t2 4.70359
R34 VDD1.n2 VDD1.t4 4.70359
R35 VDD1.n0 VDD1.t1 4.70359
R36 VDD1.n0 VDD1.t3 4.70359
R37 VDD1 VDD1.n3 0.166448
R38 VTAIL.n7 VTAIL.t2 60.1367
R39 VTAIL.n10 VTAIL.t10 60.1365
R40 VTAIL.n11 VTAIL.t1 60.1365
R41 VTAIL.n2 VTAIL.t6 60.1365
R42 VTAIL.n9 VTAIL.n8 55.4336
R43 VTAIL.n6 VTAIL.n5 55.4336
R44 VTAIL.n1 VTAIL.n0 55.4334
R45 VTAIL.n4 VTAIL.n3 55.4334
R46 VTAIL.n6 VTAIL.n4 17.7893
R47 VTAIL.n11 VTAIL.n10 16.8927
R48 VTAIL.n0 VTAIL.t4 4.70359
R49 VTAIL.n0 VTAIL.t0 4.70359
R50 VTAIL.n3 VTAIL.t7 4.70359
R51 VTAIL.n3 VTAIL.t11 4.70359
R52 VTAIL.n8 VTAIL.t8 4.70359
R53 VTAIL.n8 VTAIL.t9 4.70359
R54 VTAIL.n5 VTAIL.t3 4.70359
R55 VTAIL.n5 VTAIL.t5 4.70359
R56 VTAIL.n9 VTAIL.n7 0.918603
R57 VTAIL.n2 VTAIL.n1 0.918603
R58 VTAIL.n7 VTAIL.n6 0.897052
R59 VTAIL.n10 VTAIL.n9 0.897052
R60 VTAIL.n4 VTAIL.n2 0.897052
R61 VTAIL VTAIL.n11 0.614724
R62 VTAIL VTAIL.n1 0.282828
R63 B.n411 B.n410 585
R64 B.n412 B.n411 585
R65 B.n160 B.n65 585
R66 B.n159 B.n158 585
R67 B.n157 B.n156 585
R68 B.n155 B.n154 585
R69 B.n153 B.n152 585
R70 B.n151 B.n150 585
R71 B.n149 B.n148 585
R72 B.n147 B.n146 585
R73 B.n145 B.n144 585
R74 B.n143 B.n142 585
R75 B.n141 B.n140 585
R76 B.n139 B.n138 585
R77 B.n137 B.n136 585
R78 B.n135 B.n134 585
R79 B.n133 B.n132 585
R80 B.n131 B.n130 585
R81 B.n129 B.n128 585
R82 B.n127 B.n126 585
R83 B.n125 B.n124 585
R84 B.n123 B.n122 585
R85 B.n121 B.n120 585
R86 B.n119 B.n118 585
R87 B.n117 B.n116 585
R88 B.n115 B.n114 585
R89 B.n113 B.n112 585
R90 B.n111 B.n110 585
R91 B.n109 B.n108 585
R92 B.n106 B.n105 585
R93 B.n104 B.n103 585
R94 B.n102 B.n101 585
R95 B.n100 B.n99 585
R96 B.n98 B.n97 585
R97 B.n96 B.n95 585
R98 B.n94 B.n93 585
R99 B.n92 B.n91 585
R100 B.n90 B.n89 585
R101 B.n88 B.n87 585
R102 B.n86 B.n85 585
R103 B.n84 B.n83 585
R104 B.n82 B.n81 585
R105 B.n80 B.n79 585
R106 B.n78 B.n77 585
R107 B.n76 B.n75 585
R108 B.n74 B.n73 585
R109 B.n72 B.n71 585
R110 B.n40 B.n39 585
R111 B.n409 B.n41 585
R112 B.n413 B.n41 585
R113 B.n408 B.n407 585
R114 B.n407 B.n37 585
R115 B.n406 B.n36 585
R116 B.n419 B.n36 585
R117 B.n405 B.n35 585
R118 B.n420 B.n35 585
R119 B.n404 B.n34 585
R120 B.n421 B.n34 585
R121 B.n403 B.n402 585
R122 B.n402 B.n30 585
R123 B.n401 B.n29 585
R124 B.n427 B.n29 585
R125 B.n400 B.n28 585
R126 B.n428 B.n28 585
R127 B.n399 B.n27 585
R128 B.n429 B.n27 585
R129 B.n398 B.n397 585
R130 B.n397 B.n23 585
R131 B.n396 B.n22 585
R132 B.n435 B.n22 585
R133 B.n395 B.n21 585
R134 B.n436 B.n21 585
R135 B.n394 B.n20 585
R136 B.n437 B.n20 585
R137 B.n393 B.n392 585
R138 B.n392 B.n16 585
R139 B.n391 B.n15 585
R140 B.n443 B.n15 585
R141 B.n390 B.n14 585
R142 B.n444 B.n14 585
R143 B.n389 B.n13 585
R144 B.n445 B.n13 585
R145 B.n388 B.n387 585
R146 B.n387 B.n12 585
R147 B.n386 B.n385 585
R148 B.n386 B.n8 585
R149 B.n384 B.n7 585
R150 B.n452 B.n7 585
R151 B.n383 B.n6 585
R152 B.n453 B.n6 585
R153 B.n382 B.n5 585
R154 B.n454 B.n5 585
R155 B.n381 B.n380 585
R156 B.n380 B.n4 585
R157 B.n379 B.n161 585
R158 B.n379 B.n378 585
R159 B.n368 B.n162 585
R160 B.n371 B.n162 585
R161 B.n370 B.n369 585
R162 B.n372 B.n370 585
R163 B.n367 B.n167 585
R164 B.n167 B.n166 585
R165 B.n366 B.n365 585
R166 B.n365 B.n364 585
R167 B.n169 B.n168 585
R168 B.n170 B.n169 585
R169 B.n357 B.n356 585
R170 B.n358 B.n357 585
R171 B.n355 B.n174 585
R172 B.n178 B.n174 585
R173 B.n354 B.n353 585
R174 B.n353 B.n352 585
R175 B.n176 B.n175 585
R176 B.n177 B.n176 585
R177 B.n345 B.n344 585
R178 B.n346 B.n345 585
R179 B.n343 B.n183 585
R180 B.n183 B.n182 585
R181 B.n342 B.n341 585
R182 B.n341 B.n340 585
R183 B.n185 B.n184 585
R184 B.n186 B.n185 585
R185 B.n333 B.n332 585
R186 B.n334 B.n333 585
R187 B.n331 B.n191 585
R188 B.n191 B.n190 585
R189 B.n330 B.n329 585
R190 B.n329 B.n328 585
R191 B.n193 B.n192 585
R192 B.n194 B.n193 585
R193 B.n321 B.n320 585
R194 B.n322 B.n321 585
R195 B.n197 B.n196 585
R196 B.n226 B.n225 585
R197 B.n227 B.n223 585
R198 B.n223 B.n198 585
R199 B.n229 B.n228 585
R200 B.n231 B.n222 585
R201 B.n234 B.n233 585
R202 B.n235 B.n221 585
R203 B.n237 B.n236 585
R204 B.n239 B.n220 585
R205 B.n242 B.n241 585
R206 B.n243 B.n219 585
R207 B.n245 B.n244 585
R208 B.n247 B.n218 585
R209 B.n250 B.n249 585
R210 B.n251 B.n217 585
R211 B.n253 B.n252 585
R212 B.n255 B.n216 585
R213 B.n258 B.n257 585
R214 B.n259 B.n213 585
R215 B.n262 B.n261 585
R216 B.n264 B.n212 585
R217 B.n267 B.n266 585
R218 B.n268 B.n211 585
R219 B.n270 B.n269 585
R220 B.n272 B.n210 585
R221 B.n275 B.n274 585
R222 B.n276 B.n209 585
R223 B.n281 B.n280 585
R224 B.n283 B.n208 585
R225 B.n286 B.n285 585
R226 B.n287 B.n207 585
R227 B.n289 B.n288 585
R228 B.n291 B.n206 585
R229 B.n294 B.n293 585
R230 B.n295 B.n205 585
R231 B.n297 B.n296 585
R232 B.n299 B.n204 585
R233 B.n302 B.n301 585
R234 B.n303 B.n203 585
R235 B.n305 B.n304 585
R236 B.n307 B.n202 585
R237 B.n310 B.n309 585
R238 B.n311 B.n201 585
R239 B.n313 B.n312 585
R240 B.n315 B.n200 585
R241 B.n318 B.n317 585
R242 B.n319 B.n199 585
R243 B.n324 B.n323 585
R244 B.n323 B.n322 585
R245 B.n325 B.n195 585
R246 B.n195 B.n194 585
R247 B.n327 B.n326 585
R248 B.n328 B.n327 585
R249 B.n189 B.n188 585
R250 B.n190 B.n189 585
R251 B.n336 B.n335 585
R252 B.n335 B.n334 585
R253 B.n337 B.n187 585
R254 B.n187 B.n186 585
R255 B.n339 B.n338 585
R256 B.n340 B.n339 585
R257 B.n181 B.n180 585
R258 B.n182 B.n181 585
R259 B.n348 B.n347 585
R260 B.n347 B.n346 585
R261 B.n349 B.n179 585
R262 B.n179 B.n177 585
R263 B.n351 B.n350 585
R264 B.n352 B.n351 585
R265 B.n173 B.n172 585
R266 B.n178 B.n173 585
R267 B.n360 B.n359 585
R268 B.n359 B.n358 585
R269 B.n361 B.n171 585
R270 B.n171 B.n170 585
R271 B.n363 B.n362 585
R272 B.n364 B.n363 585
R273 B.n165 B.n164 585
R274 B.n166 B.n165 585
R275 B.n374 B.n373 585
R276 B.n373 B.n372 585
R277 B.n375 B.n163 585
R278 B.n371 B.n163 585
R279 B.n377 B.n376 585
R280 B.n378 B.n377 585
R281 B.n3 B.n0 585
R282 B.n4 B.n3 585
R283 B.n451 B.n1 585
R284 B.n452 B.n451 585
R285 B.n450 B.n449 585
R286 B.n450 B.n8 585
R287 B.n448 B.n9 585
R288 B.n12 B.n9 585
R289 B.n447 B.n446 585
R290 B.n446 B.n445 585
R291 B.n11 B.n10 585
R292 B.n444 B.n11 585
R293 B.n442 B.n441 585
R294 B.n443 B.n442 585
R295 B.n440 B.n17 585
R296 B.n17 B.n16 585
R297 B.n439 B.n438 585
R298 B.n438 B.n437 585
R299 B.n19 B.n18 585
R300 B.n436 B.n19 585
R301 B.n434 B.n433 585
R302 B.n435 B.n434 585
R303 B.n432 B.n24 585
R304 B.n24 B.n23 585
R305 B.n431 B.n430 585
R306 B.n430 B.n429 585
R307 B.n26 B.n25 585
R308 B.n428 B.n26 585
R309 B.n426 B.n425 585
R310 B.n427 B.n426 585
R311 B.n424 B.n31 585
R312 B.n31 B.n30 585
R313 B.n423 B.n422 585
R314 B.n422 B.n421 585
R315 B.n33 B.n32 585
R316 B.n420 B.n33 585
R317 B.n418 B.n417 585
R318 B.n419 B.n418 585
R319 B.n416 B.n38 585
R320 B.n38 B.n37 585
R321 B.n415 B.n414 585
R322 B.n414 B.n413 585
R323 B.n455 B.n454 585
R324 B.n453 B.n2 585
R325 B.n414 B.n40 473.281
R326 B.n411 B.n41 473.281
R327 B.n321 B.n199 473.281
R328 B.n323 B.n197 473.281
R329 B.n69 B.t10 345.747
R330 B.n66 B.t14 345.747
R331 B.n277 B.t6 345.747
R332 B.n214 B.t17 345.747
R333 B.n412 B.n64 256.663
R334 B.n412 B.n63 256.663
R335 B.n412 B.n62 256.663
R336 B.n412 B.n61 256.663
R337 B.n412 B.n60 256.663
R338 B.n412 B.n59 256.663
R339 B.n412 B.n58 256.663
R340 B.n412 B.n57 256.663
R341 B.n412 B.n56 256.663
R342 B.n412 B.n55 256.663
R343 B.n412 B.n54 256.663
R344 B.n412 B.n53 256.663
R345 B.n412 B.n52 256.663
R346 B.n412 B.n51 256.663
R347 B.n412 B.n50 256.663
R348 B.n412 B.n49 256.663
R349 B.n412 B.n48 256.663
R350 B.n412 B.n47 256.663
R351 B.n412 B.n46 256.663
R352 B.n412 B.n45 256.663
R353 B.n412 B.n44 256.663
R354 B.n412 B.n43 256.663
R355 B.n412 B.n42 256.663
R356 B.n224 B.n198 256.663
R357 B.n230 B.n198 256.663
R358 B.n232 B.n198 256.663
R359 B.n238 B.n198 256.663
R360 B.n240 B.n198 256.663
R361 B.n246 B.n198 256.663
R362 B.n248 B.n198 256.663
R363 B.n254 B.n198 256.663
R364 B.n256 B.n198 256.663
R365 B.n263 B.n198 256.663
R366 B.n265 B.n198 256.663
R367 B.n271 B.n198 256.663
R368 B.n273 B.n198 256.663
R369 B.n282 B.n198 256.663
R370 B.n284 B.n198 256.663
R371 B.n290 B.n198 256.663
R372 B.n292 B.n198 256.663
R373 B.n298 B.n198 256.663
R374 B.n300 B.n198 256.663
R375 B.n306 B.n198 256.663
R376 B.n308 B.n198 256.663
R377 B.n314 B.n198 256.663
R378 B.n316 B.n198 256.663
R379 B.n457 B.n456 256.663
R380 B.n73 B.n72 163.367
R381 B.n77 B.n76 163.367
R382 B.n81 B.n80 163.367
R383 B.n85 B.n84 163.367
R384 B.n89 B.n88 163.367
R385 B.n93 B.n92 163.367
R386 B.n97 B.n96 163.367
R387 B.n101 B.n100 163.367
R388 B.n105 B.n104 163.367
R389 B.n110 B.n109 163.367
R390 B.n114 B.n113 163.367
R391 B.n118 B.n117 163.367
R392 B.n122 B.n121 163.367
R393 B.n126 B.n125 163.367
R394 B.n130 B.n129 163.367
R395 B.n134 B.n133 163.367
R396 B.n138 B.n137 163.367
R397 B.n142 B.n141 163.367
R398 B.n146 B.n145 163.367
R399 B.n150 B.n149 163.367
R400 B.n154 B.n153 163.367
R401 B.n158 B.n157 163.367
R402 B.n411 B.n65 163.367
R403 B.n321 B.n193 163.367
R404 B.n329 B.n193 163.367
R405 B.n329 B.n191 163.367
R406 B.n333 B.n191 163.367
R407 B.n333 B.n185 163.367
R408 B.n341 B.n185 163.367
R409 B.n341 B.n183 163.367
R410 B.n345 B.n183 163.367
R411 B.n345 B.n176 163.367
R412 B.n353 B.n176 163.367
R413 B.n353 B.n174 163.367
R414 B.n357 B.n174 163.367
R415 B.n357 B.n169 163.367
R416 B.n365 B.n169 163.367
R417 B.n365 B.n167 163.367
R418 B.n370 B.n167 163.367
R419 B.n370 B.n162 163.367
R420 B.n379 B.n162 163.367
R421 B.n380 B.n379 163.367
R422 B.n380 B.n5 163.367
R423 B.n6 B.n5 163.367
R424 B.n7 B.n6 163.367
R425 B.n386 B.n7 163.367
R426 B.n387 B.n386 163.367
R427 B.n387 B.n13 163.367
R428 B.n14 B.n13 163.367
R429 B.n15 B.n14 163.367
R430 B.n392 B.n15 163.367
R431 B.n392 B.n20 163.367
R432 B.n21 B.n20 163.367
R433 B.n22 B.n21 163.367
R434 B.n397 B.n22 163.367
R435 B.n397 B.n27 163.367
R436 B.n28 B.n27 163.367
R437 B.n29 B.n28 163.367
R438 B.n402 B.n29 163.367
R439 B.n402 B.n34 163.367
R440 B.n35 B.n34 163.367
R441 B.n36 B.n35 163.367
R442 B.n407 B.n36 163.367
R443 B.n407 B.n41 163.367
R444 B.n225 B.n223 163.367
R445 B.n229 B.n223 163.367
R446 B.n233 B.n231 163.367
R447 B.n237 B.n221 163.367
R448 B.n241 B.n239 163.367
R449 B.n245 B.n219 163.367
R450 B.n249 B.n247 163.367
R451 B.n253 B.n217 163.367
R452 B.n257 B.n255 163.367
R453 B.n262 B.n213 163.367
R454 B.n266 B.n264 163.367
R455 B.n270 B.n211 163.367
R456 B.n274 B.n272 163.367
R457 B.n281 B.n209 163.367
R458 B.n285 B.n283 163.367
R459 B.n289 B.n207 163.367
R460 B.n293 B.n291 163.367
R461 B.n297 B.n205 163.367
R462 B.n301 B.n299 163.367
R463 B.n305 B.n203 163.367
R464 B.n309 B.n307 163.367
R465 B.n313 B.n201 163.367
R466 B.n317 B.n315 163.367
R467 B.n323 B.n195 163.367
R468 B.n327 B.n195 163.367
R469 B.n327 B.n189 163.367
R470 B.n335 B.n189 163.367
R471 B.n335 B.n187 163.367
R472 B.n339 B.n187 163.367
R473 B.n339 B.n181 163.367
R474 B.n347 B.n181 163.367
R475 B.n347 B.n179 163.367
R476 B.n351 B.n179 163.367
R477 B.n351 B.n173 163.367
R478 B.n359 B.n173 163.367
R479 B.n359 B.n171 163.367
R480 B.n363 B.n171 163.367
R481 B.n363 B.n165 163.367
R482 B.n373 B.n165 163.367
R483 B.n373 B.n163 163.367
R484 B.n377 B.n163 163.367
R485 B.n377 B.n3 163.367
R486 B.n455 B.n3 163.367
R487 B.n451 B.n2 163.367
R488 B.n451 B.n450 163.367
R489 B.n450 B.n9 163.367
R490 B.n446 B.n9 163.367
R491 B.n446 B.n11 163.367
R492 B.n442 B.n11 163.367
R493 B.n442 B.n17 163.367
R494 B.n438 B.n17 163.367
R495 B.n438 B.n19 163.367
R496 B.n434 B.n19 163.367
R497 B.n434 B.n24 163.367
R498 B.n430 B.n24 163.367
R499 B.n430 B.n26 163.367
R500 B.n426 B.n26 163.367
R501 B.n426 B.n31 163.367
R502 B.n422 B.n31 163.367
R503 B.n422 B.n33 163.367
R504 B.n418 B.n33 163.367
R505 B.n418 B.n38 163.367
R506 B.n414 B.n38 163.367
R507 B.n322 B.n198 131.049
R508 B.n413 B.n412 131.049
R509 B.n66 B.t15 93.8085
R510 B.n277 B.t9 93.8085
R511 B.n69 B.t12 93.8046
R512 B.n214 B.t19 93.8046
R513 B.n322 B.n194 78.8619
R514 B.n328 B.n194 78.8619
R515 B.n328 B.n190 78.8619
R516 B.n334 B.n190 78.8619
R517 B.n340 B.n186 78.8619
R518 B.n340 B.n182 78.8619
R519 B.n346 B.n182 78.8619
R520 B.n346 B.n177 78.8619
R521 B.n352 B.n177 78.8619
R522 B.n352 B.n178 78.8619
R523 B.n358 B.n170 78.8619
R524 B.n364 B.n170 78.8619
R525 B.n372 B.n166 78.8619
R526 B.n372 B.n371 78.8619
R527 B.n378 B.n4 78.8619
R528 B.n454 B.n4 78.8619
R529 B.n454 B.n453 78.8619
R530 B.n453 B.n452 78.8619
R531 B.n452 B.n8 78.8619
R532 B.n445 B.n12 78.8619
R533 B.n445 B.n444 78.8619
R534 B.n443 B.n16 78.8619
R535 B.n437 B.n16 78.8619
R536 B.n436 B.n435 78.8619
R537 B.n435 B.n23 78.8619
R538 B.n429 B.n23 78.8619
R539 B.n429 B.n428 78.8619
R540 B.n428 B.n427 78.8619
R541 B.n427 B.n30 78.8619
R542 B.n421 B.n420 78.8619
R543 B.n420 B.n419 78.8619
R544 B.n419 B.n37 78.8619
R545 B.n413 B.n37 78.8619
R546 B.n334 B.t7 77.7021
R547 B.n421 B.t11 77.7021
R548 B.n67 B.t16 73.6388
R549 B.n278 B.t8 73.6388
R550 B.n70 B.t13 73.6349
R551 B.n215 B.t18 73.6349
R552 B.n42 B.n40 71.676
R553 B.n73 B.n43 71.676
R554 B.n77 B.n44 71.676
R555 B.n81 B.n45 71.676
R556 B.n85 B.n46 71.676
R557 B.n89 B.n47 71.676
R558 B.n93 B.n48 71.676
R559 B.n97 B.n49 71.676
R560 B.n101 B.n50 71.676
R561 B.n105 B.n51 71.676
R562 B.n110 B.n52 71.676
R563 B.n114 B.n53 71.676
R564 B.n118 B.n54 71.676
R565 B.n122 B.n55 71.676
R566 B.n126 B.n56 71.676
R567 B.n130 B.n57 71.676
R568 B.n134 B.n58 71.676
R569 B.n138 B.n59 71.676
R570 B.n142 B.n60 71.676
R571 B.n146 B.n61 71.676
R572 B.n150 B.n62 71.676
R573 B.n154 B.n63 71.676
R574 B.n158 B.n64 71.676
R575 B.n65 B.n64 71.676
R576 B.n157 B.n63 71.676
R577 B.n153 B.n62 71.676
R578 B.n149 B.n61 71.676
R579 B.n145 B.n60 71.676
R580 B.n141 B.n59 71.676
R581 B.n137 B.n58 71.676
R582 B.n133 B.n57 71.676
R583 B.n129 B.n56 71.676
R584 B.n125 B.n55 71.676
R585 B.n121 B.n54 71.676
R586 B.n117 B.n53 71.676
R587 B.n113 B.n52 71.676
R588 B.n109 B.n51 71.676
R589 B.n104 B.n50 71.676
R590 B.n100 B.n49 71.676
R591 B.n96 B.n48 71.676
R592 B.n92 B.n47 71.676
R593 B.n88 B.n46 71.676
R594 B.n84 B.n45 71.676
R595 B.n80 B.n44 71.676
R596 B.n76 B.n43 71.676
R597 B.n72 B.n42 71.676
R598 B.n224 B.n197 71.676
R599 B.n230 B.n229 71.676
R600 B.n233 B.n232 71.676
R601 B.n238 B.n237 71.676
R602 B.n241 B.n240 71.676
R603 B.n246 B.n245 71.676
R604 B.n249 B.n248 71.676
R605 B.n254 B.n253 71.676
R606 B.n257 B.n256 71.676
R607 B.n263 B.n262 71.676
R608 B.n266 B.n265 71.676
R609 B.n271 B.n270 71.676
R610 B.n274 B.n273 71.676
R611 B.n282 B.n281 71.676
R612 B.n285 B.n284 71.676
R613 B.n290 B.n289 71.676
R614 B.n293 B.n292 71.676
R615 B.n298 B.n297 71.676
R616 B.n301 B.n300 71.676
R617 B.n306 B.n305 71.676
R618 B.n309 B.n308 71.676
R619 B.n314 B.n313 71.676
R620 B.n317 B.n316 71.676
R621 B.n225 B.n224 71.676
R622 B.n231 B.n230 71.676
R623 B.n232 B.n221 71.676
R624 B.n239 B.n238 71.676
R625 B.n240 B.n219 71.676
R626 B.n247 B.n246 71.676
R627 B.n248 B.n217 71.676
R628 B.n255 B.n254 71.676
R629 B.n256 B.n213 71.676
R630 B.n264 B.n263 71.676
R631 B.n265 B.n211 71.676
R632 B.n272 B.n271 71.676
R633 B.n273 B.n209 71.676
R634 B.n283 B.n282 71.676
R635 B.n284 B.n207 71.676
R636 B.n291 B.n290 71.676
R637 B.n292 B.n205 71.676
R638 B.n299 B.n298 71.676
R639 B.n300 B.n203 71.676
R640 B.n307 B.n306 71.676
R641 B.n308 B.n201 71.676
R642 B.n315 B.n314 71.676
R643 B.n316 B.n199 71.676
R644 B.n456 B.n455 71.676
R645 B.n456 B.n2 71.676
R646 B.n107 B.n70 59.5399
R647 B.n68 B.n67 59.5399
R648 B.n279 B.n278 59.5399
R649 B.n260 B.n215 59.5399
R650 B.n358 B.t3 59.1465
R651 B.n437 B.t1 59.1465
R652 B.t5 B.n166 54.5076
R653 B.n444 B.t0 54.5076
R654 B.n378 B.t2 49.8687
R655 B.t4 B.n8 49.8687
R656 B.n324 B.n196 30.7517
R657 B.n320 B.n319 30.7517
R658 B.n410 B.n409 30.7517
R659 B.n415 B.n39 30.7517
R660 B.n371 B.t2 28.9936
R661 B.n12 B.t4 28.9936
R662 B.n364 B.t5 24.3547
R663 B.t0 B.n443 24.3547
R664 B.n70 B.n69 20.1702
R665 B.n67 B.n66 20.1702
R666 B.n278 B.n277 20.1702
R667 B.n215 B.n214 20.1702
R668 B.n178 B.t3 19.7158
R669 B.t1 B.n436 19.7158
R670 B B.n457 18.0485
R671 B.n325 B.n324 10.6151
R672 B.n326 B.n325 10.6151
R673 B.n326 B.n188 10.6151
R674 B.n336 B.n188 10.6151
R675 B.n337 B.n336 10.6151
R676 B.n338 B.n337 10.6151
R677 B.n338 B.n180 10.6151
R678 B.n348 B.n180 10.6151
R679 B.n349 B.n348 10.6151
R680 B.n350 B.n349 10.6151
R681 B.n350 B.n172 10.6151
R682 B.n360 B.n172 10.6151
R683 B.n361 B.n360 10.6151
R684 B.n362 B.n361 10.6151
R685 B.n362 B.n164 10.6151
R686 B.n374 B.n164 10.6151
R687 B.n375 B.n374 10.6151
R688 B.n376 B.n375 10.6151
R689 B.n376 B.n0 10.6151
R690 B.n226 B.n196 10.6151
R691 B.n227 B.n226 10.6151
R692 B.n228 B.n227 10.6151
R693 B.n228 B.n222 10.6151
R694 B.n234 B.n222 10.6151
R695 B.n235 B.n234 10.6151
R696 B.n236 B.n235 10.6151
R697 B.n236 B.n220 10.6151
R698 B.n242 B.n220 10.6151
R699 B.n243 B.n242 10.6151
R700 B.n244 B.n243 10.6151
R701 B.n244 B.n218 10.6151
R702 B.n250 B.n218 10.6151
R703 B.n251 B.n250 10.6151
R704 B.n252 B.n251 10.6151
R705 B.n252 B.n216 10.6151
R706 B.n258 B.n216 10.6151
R707 B.n259 B.n258 10.6151
R708 B.n261 B.n212 10.6151
R709 B.n267 B.n212 10.6151
R710 B.n268 B.n267 10.6151
R711 B.n269 B.n268 10.6151
R712 B.n269 B.n210 10.6151
R713 B.n275 B.n210 10.6151
R714 B.n276 B.n275 10.6151
R715 B.n280 B.n276 10.6151
R716 B.n286 B.n208 10.6151
R717 B.n287 B.n286 10.6151
R718 B.n288 B.n287 10.6151
R719 B.n288 B.n206 10.6151
R720 B.n294 B.n206 10.6151
R721 B.n295 B.n294 10.6151
R722 B.n296 B.n295 10.6151
R723 B.n296 B.n204 10.6151
R724 B.n302 B.n204 10.6151
R725 B.n303 B.n302 10.6151
R726 B.n304 B.n303 10.6151
R727 B.n304 B.n202 10.6151
R728 B.n310 B.n202 10.6151
R729 B.n311 B.n310 10.6151
R730 B.n312 B.n311 10.6151
R731 B.n312 B.n200 10.6151
R732 B.n318 B.n200 10.6151
R733 B.n319 B.n318 10.6151
R734 B.n320 B.n192 10.6151
R735 B.n330 B.n192 10.6151
R736 B.n331 B.n330 10.6151
R737 B.n332 B.n331 10.6151
R738 B.n332 B.n184 10.6151
R739 B.n342 B.n184 10.6151
R740 B.n343 B.n342 10.6151
R741 B.n344 B.n343 10.6151
R742 B.n344 B.n175 10.6151
R743 B.n354 B.n175 10.6151
R744 B.n355 B.n354 10.6151
R745 B.n356 B.n355 10.6151
R746 B.n356 B.n168 10.6151
R747 B.n366 B.n168 10.6151
R748 B.n367 B.n366 10.6151
R749 B.n369 B.n367 10.6151
R750 B.n369 B.n368 10.6151
R751 B.n368 B.n161 10.6151
R752 B.n381 B.n161 10.6151
R753 B.n382 B.n381 10.6151
R754 B.n383 B.n382 10.6151
R755 B.n384 B.n383 10.6151
R756 B.n385 B.n384 10.6151
R757 B.n388 B.n385 10.6151
R758 B.n389 B.n388 10.6151
R759 B.n390 B.n389 10.6151
R760 B.n391 B.n390 10.6151
R761 B.n393 B.n391 10.6151
R762 B.n394 B.n393 10.6151
R763 B.n395 B.n394 10.6151
R764 B.n396 B.n395 10.6151
R765 B.n398 B.n396 10.6151
R766 B.n399 B.n398 10.6151
R767 B.n400 B.n399 10.6151
R768 B.n401 B.n400 10.6151
R769 B.n403 B.n401 10.6151
R770 B.n404 B.n403 10.6151
R771 B.n405 B.n404 10.6151
R772 B.n406 B.n405 10.6151
R773 B.n408 B.n406 10.6151
R774 B.n409 B.n408 10.6151
R775 B.n449 B.n1 10.6151
R776 B.n449 B.n448 10.6151
R777 B.n448 B.n447 10.6151
R778 B.n447 B.n10 10.6151
R779 B.n441 B.n10 10.6151
R780 B.n441 B.n440 10.6151
R781 B.n440 B.n439 10.6151
R782 B.n439 B.n18 10.6151
R783 B.n433 B.n18 10.6151
R784 B.n433 B.n432 10.6151
R785 B.n432 B.n431 10.6151
R786 B.n431 B.n25 10.6151
R787 B.n425 B.n25 10.6151
R788 B.n425 B.n424 10.6151
R789 B.n424 B.n423 10.6151
R790 B.n423 B.n32 10.6151
R791 B.n417 B.n32 10.6151
R792 B.n417 B.n416 10.6151
R793 B.n416 B.n415 10.6151
R794 B.n71 B.n39 10.6151
R795 B.n74 B.n71 10.6151
R796 B.n75 B.n74 10.6151
R797 B.n78 B.n75 10.6151
R798 B.n79 B.n78 10.6151
R799 B.n82 B.n79 10.6151
R800 B.n83 B.n82 10.6151
R801 B.n86 B.n83 10.6151
R802 B.n87 B.n86 10.6151
R803 B.n90 B.n87 10.6151
R804 B.n91 B.n90 10.6151
R805 B.n94 B.n91 10.6151
R806 B.n95 B.n94 10.6151
R807 B.n98 B.n95 10.6151
R808 B.n99 B.n98 10.6151
R809 B.n102 B.n99 10.6151
R810 B.n103 B.n102 10.6151
R811 B.n106 B.n103 10.6151
R812 B.n111 B.n108 10.6151
R813 B.n112 B.n111 10.6151
R814 B.n115 B.n112 10.6151
R815 B.n116 B.n115 10.6151
R816 B.n119 B.n116 10.6151
R817 B.n120 B.n119 10.6151
R818 B.n123 B.n120 10.6151
R819 B.n124 B.n123 10.6151
R820 B.n128 B.n127 10.6151
R821 B.n131 B.n128 10.6151
R822 B.n132 B.n131 10.6151
R823 B.n135 B.n132 10.6151
R824 B.n136 B.n135 10.6151
R825 B.n139 B.n136 10.6151
R826 B.n140 B.n139 10.6151
R827 B.n143 B.n140 10.6151
R828 B.n144 B.n143 10.6151
R829 B.n147 B.n144 10.6151
R830 B.n148 B.n147 10.6151
R831 B.n151 B.n148 10.6151
R832 B.n152 B.n151 10.6151
R833 B.n155 B.n152 10.6151
R834 B.n156 B.n155 10.6151
R835 B.n159 B.n156 10.6151
R836 B.n160 B.n159 10.6151
R837 B.n410 B.n160 10.6151
R838 B.n457 B.n0 8.11757
R839 B.n457 B.n1 8.11757
R840 B.n261 B.n260 6.5566
R841 B.n280 B.n279 6.5566
R842 B.n108 B.n107 6.5566
R843 B.n124 B.n68 6.5566
R844 B.n260 B.n259 4.05904
R845 B.n279 B.n208 4.05904
R846 B.n107 B.n106 4.05904
R847 B.n127 B.n68 4.05904
R848 B.t7 B.n186 1.16023
R849 B.t11 B.n30 1.16023
R850 VN.n1 VN.t3 220.362
R851 VN.n7 VN.t4 220.362
R852 VN.n2 VN.t5 198.571
R853 VN.n4 VN.t0 198.571
R854 VN.n8 VN.t2 198.571
R855 VN.n10 VN.t1 198.571
R856 VN.n5 VN.n4 161.3
R857 VN.n11 VN.n10 161.3
R858 VN.n9 VN.n6 161.3
R859 VN.n3 VN.n0 161.3
R860 VN.n7 VN.n6 44.8565
R861 VN.n1 VN.n0 44.8565
R862 VN VN.n11 35.7297
R863 VN.n4 VN.n3 27.0217
R864 VN.n10 VN.n9 27.0217
R865 VN.n3 VN.n2 21.1793
R866 VN.n9 VN.n8 21.1793
R867 VN.n2 VN.n1 20.1275
R868 VN.n8 VN.n7 20.1275
R869 VN.n11 VN.n6 0.189894
R870 VN.n5 VN.n0 0.189894
R871 VN VN.n5 0.0516364
R872 VDD2.n1 VDD2.t2 77.4323
R873 VDD2.n2 VDD2.t4 76.8155
R874 VDD2.n1 VDD2.n0 72.281
R875 VDD2 VDD2.n3 72.2782
R876 VDD2.n2 VDD2.n1 30.2584
R877 VDD2.n3 VDD2.t3 4.70359
R878 VDD2.n3 VDD2.t1 4.70359
R879 VDD2.n0 VDD2.t0 4.70359
R880 VDD2.n0 VDD2.t5 4.70359
R881 VDD2 VDD2.n2 0.731103
C0 VTAIL VDD1 4.68791f
C1 VDD2 VN 1.75503f
C2 VDD1 VP 1.90233f
C3 VTAIL VN 1.82593f
C4 VDD2 VTAIL 4.7264f
C5 VP VN 3.65413f
C6 VDD1 VN 0.152107f
C7 VDD2 VP 0.30158f
C8 VDD2 VDD1 0.710838f
C9 VTAIL VP 1.84021f
C10 VDD2 B 2.990646f
C11 VDD1 B 3.201733f
C12 VTAIL B 3.358459f
C13 VN B 6.029113f
C14 VP B 5.151605f
C15 VDD2.t2 B 0.570732f
C16 VDD2.t0 B 0.056523f
C17 VDD2.t5 B 0.056523f
C18 VDD2.n0 B 0.44882f
C19 VDD2.n1 B 1.08266f
C20 VDD2.t4 B 0.56908f
C21 VDD2.n2 B 1.10746f
C22 VDD2.t3 B 0.056523f
C23 VDD2.t1 B 0.056523f
C24 VDD2.n3 B 0.448806f
C25 VN.n0 B 0.101161f
C26 VN.t3 B 0.224977f
C27 VN.n1 B 0.101477f
C28 VN.t5 B 0.214104f
C29 VN.n2 B 0.112f
C30 VN.n3 B 0.00552f
C31 VN.t0 B 0.214104f
C32 VN.n4 B 0.108381f
C33 VN.n5 B 0.018852f
C34 VN.n6 B 0.101161f
C35 VN.t4 B 0.224977f
C36 VN.n7 B 0.101477f
C37 VN.t2 B 0.214104f
C38 VN.n8 B 0.112f
C39 VN.n9 B 0.00552f
C40 VN.t1 B 0.214104f
C41 VN.n10 B 0.108381f
C42 VN.n11 B 0.754965f
C43 VTAIL.t4 B 0.065283f
C44 VTAIL.t0 B 0.065283f
C45 VTAIL.n0 B 0.472847f
C46 VTAIL.n1 B 0.247499f
C47 VTAIL.t6 B 0.605094f
C48 VTAIL.n2 B 0.332136f
C49 VTAIL.t7 B 0.065283f
C50 VTAIL.t11 B 0.065283f
C51 VTAIL.n3 B 0.472847f
C52 VTAIL.n4 B 0.837701f
C53 VTAIL.t3 B 0.065283f
C54 VTAIL.t5 B 0.065283f
C55 VTAIL.n5 B 0.472849f
C56 VTAIL.n6 B 0.837699f
C57 VTAIL.t2 B 0.605096f
C58 VTAIL.n7 B 0.332133f
C59 VTAIL.t8 B 0.065283f
C60 VTAIL.t9 B 0.065283f
C61 VTAIL.n8 B 0.472849f
C62 VTAIL.n9 B 0.286334f
C63 VTAIL.t10 B 0.605094f
C64 VTAIL.n10 B 0.826811f
C65 VTAIL.t1 B 0.605094f
C66 VTAIL.n11 B 0.80896f
C67 VDD1.t0 B 0.563562f
C68 VDD1.t5 B 0.563212f
C69 VDD1.t1 B 0.055779f
C70 VDD1.t3 B 0.055779f
C71 VDD1.n0 B 0.442907f
C72 VDD1.n1 B 1.11785f
C73 VDD1.t2 B 0.055779f
C74 VDD1.t4 B 0.055779f
C75 VDD1.n2 B 0.442445f
C76 VDD1.n3 B 1.09029f
C77 VP.n0 B 0.024553f
C78 VP.n1 B 0.005572f
C79 VP.n2 B 0.102105f
C80 VP.t1 B 0.216102f
C81 VP.t2 B 0.216102f
C82 VP.t3 B 0.227076f
C83 VP.n3 B 0.102423f
C84 VP.n4 B 0.113045f
C85 VP.n5 B 0.005572f
C86 VP.n6 B 0.109392f
C87 VP.n7 B 0.7457f
C88 VP.t4 B 0.216102f
C89 VP.n8 B 0.109392f
C90 VP.n9 B 0.770669f
C91 VP.n10 B 0.024553f
C92 VP.n11 B 0.024553f
C93 VP.t0 B 0.216102f
C94 VP.n12 B 0.110981f
C95 VP.n13 B 0.005572f
C96 VP.t5 B 0.216102f
C97 VP.n14 B 0.109392f
C98 VP.n15 B 0.019028f
.ends

