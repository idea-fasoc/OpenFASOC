* NGSPICE file created from diff_pair_sample_1540.ext - technology: sky130A

.subckt diff_pair_sample_1540 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=1.6263 ps=9.12 w=4.17 l=3.79
X1 VDD1.t8 VP.t1 VTAIL.t18 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0.68805 ps=4.5 w=4.17 l=3.79
X2 VDD2.t9 VN.t0 VTAIL.t19 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X3 VDD2.t8 VN.t1 VTAIL.t3 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0.68805 ps=4.5 w=4.17 l=3.79
X4 VTAIL.t0 VN.t2 VDD2.t7 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X5 VDD2.t6 VN.t3 VTAIL.t1 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X6 B.t11 B.t9 B.t10 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=3.79
X7 B.t8 B.t6 B.t7 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=3.79
X8 VTAIL.t12 VP.t2 VDD1.t7 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X9 VTAIL.t16 VP.t3 VDD1.t6 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X10 VDD1.t5 VP.t4 VTAIL.t10 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0.68805 ps=4.5 w=4.17 l=3.79
X11 VDD2.t5 VN.t4 VTAIL.t5 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=1.6263 ps=9.12 w=4.17 l=3.79
X12 VTAIL.t4 VN.t5 VDD2.t4 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X13 VDD2.t3 VN.t6 VTAIL.t2 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0.68805 ps=4.5 w=4.17 l=3.79
X14 B.t5 B.t3 B.t4 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=3.79
X15 VTAIL.t17 VP.t5 VDD1.t4 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X16 VTAIL.t14 VP.t6 VDD1.t3 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X17 B.t2 B.t0 B.t1 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=3.79
X18 VTAIL.t8 VN.t7 VDD2.t2 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X19 VDD1.t2 VP.t7 VTAIL.t11 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X20 VDD1.t1 VP.t8 VTAIL.t13 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X21 VTAIL.t7 VN.t8 VDD2.t1 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=0.68805 ps=4.5 w=4.17 l=3.79
X22 VDD2.t0 VN.t9 VTAIL.t6 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=1.6263 ps=9.12 w=4.17 l=3.79
X23 VDD1.t0 VP.t9 VTAIL.t9 w_n5914_n1802# sky130_fd_pr__pfet_01v8 ad=0.68805 pd=4.5 as=1.6263 ps=9.12 w=4.17 l=3.79
R0 VP.n31 VP.n30 161.3
R1 VP.n32 VP.n27 161.3
R2 VP.n34 VP.n33 161.3
R3 VP.n35 VP.n26 161.3
R4 VP.n37 VP.n36 161.3
R5 VP.n38 VP.n25 161.3
R6 VP.n40 VP.n39 161.3
R7 VP.n41 VP.n24 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n23 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n22 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n21 161.3
R14 VP.n53 VP.n52 161.3
R15 VP.n54 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n17 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n67 VP.n16 161.3
R24 VP.n122 VP.n0 161.3
R25 VP.n121 VP.n120 161.3
R26 VP.n119 VP.n1 161.3
R27 VP.n118 VP.n117 161.3
R28 VP.n116 VP.n2 161.3
R29 VP.n115 VP.n114 161.3
R30 VP.n113 VP.n3 161.3
R31 VP.n112 VP.n111 161.3
R32 VP.n109 VP.n4 161.3
R33 VP.n108 VP.n107 161.3
R34 VP.n106 VP.n5 161.3
R35 VP.n105 VP.n104 161.3
R36 VP.n103 VP.n6 161.3
R37 VP.n102 VP.n101 161.3
R38 VP.n100 VP.n7 161.3
R39 VP.n99 VP.n98 161.3
R40 VP.n96 VP.n8 161.3
R41 VP.n95 VP.n94 161.3
R42 VP.n93 VP.n9 161.3
R43 VP.n92 VP.n91 161.3
R44 VP.n90 VP.n10 161.3
R45 VP.n89 VP.n88 161.3
R46 VP.n87 VP.n11 161.3
R47 VP.n86 VP.n85 161.3
R48 VP.n83 VP.n12 161.3
R49 VP.n82 VP.n81 161.3
R50 VP.n80 VP.n13 161.3
R51 VP.n79 VP.n78 161.3
R52 VP.n77 VP.n14 161.3
R53 VP.n76 VP.n75 161.3
R54 VP.n74 VP.n15 161.3
R55 VP.n73 VP.n72 161.3
R56 VP.n28 VP.t4 58.6168
R57 VP.n71 VP.n70 58.2041
R58 VP.n124 VP.n123 58.2041
R59 VP.n69 VP.n68 58.2041
R60 VP.n29 VP.n28 56.9469
R61 VP.n91 VP.n90 56.5193
R62 VP.n104 VP.n103 56.5193
R63 VP.n49 VP.n48 56.5193
R64 VP.n36 VP.n35 56.5193
R65 VP.n70 VP.n69 53.9055
R66 VP.n78 VP.n77 47.2923
R67 VP.n117 VP.n116 47.2923
R68 VP.n62 VP.n61 47.2923
R69 VP.n77 VP.n76 33.6945
R70 VP.n117 VP.n1 33.6945
R71 VP.n62 VP.n17 33.6945
R72 VP.n71 VP.t1 26.5169
R73 VP.n84 VP.t5 26.5169
R74 VP.n97 VP.t7 26.5169
R75 VP.n110 VP.t6 26.5169
R76 VP.n123 VP.t0 26.5169
R77 VP.n68 VP.t9 26.5169
R78 VP.n55 VP.t3 26.5169
R79 VP.n42 VP.t8 26.5169
R80 VP.n29 VP.t2 26.5169
R81 VP.n72 VP.n15 24.4675
R82 VP.n76 VP.n15 24.4675
R83 VP.n78 VP.n13 24.4675
R84 VP.n82 VP.n13 24.4675
R85 VP.n83 VP.n82 24.4675
R86 VP.n85 VP.n11 24.4675
R87 VP.n89 VP.n11 24.4675
R88 VP.n90 VP.n89 24.4675
R89 VP.n91 VP.n9 24.4675
R90 VP.n95 VP.n9 24.4675
R91 VP.n96 VP.n95 24.4675
R92 VP.n98 VP.n7 24.4675
R93 VP.n102 VP.n7 24.4675
R94 VP.n103 VP.n102 24.4675
R95 VP.n104 VP.n5 24.4675
R96 VP.n108 VP.n5 24.4675
R97 VP.n109 VP.n108 24.4675
R98 VP.n111 VP.n3 24.4675
R99 VP.n115 VP.n3 24.4675
R100 VP.n116 VP.n115 24.4675
R101 VP.n121 VP.n1 24.4675
R102 VP.n122 VP.n121 24.4675
R103 VP.n66 VP.n17 24.4675
R104 VP.n67 VP.n66 24.4675
R105 VP.n49 VP.n21 24.4675
R106 VP.n53 VP.n21 24.4675
R107 VP.n54 VP.n53 24.4675
R108 VP.n56 VP.n19 24.4675
R109 VP.n60 VP.n19 24.4675
R110 VP.n61 VP.n60 24.4675
R111 VP.n36 VP.n25 24.4675
R112 VP.n40 VP.n25 24.4675
R113 VP.n41 VP.n40 24.4675
R114 VP.n43 VP.n23 24.4675
R115 VP.n47 VP.n23 24.4675
R116 VP.n48 VP.n47 24.4675
R117 VP.n30 VP.n27 24.4675
R118 VP.n34 VP.n27 24.4675
R119 VP.n35 VP.n34 24.4675
R120 VP.n72 VP.n71 23.9782
R121 VP.n123 VP.n122 23.9782
R122 VP.n68 VP.n67 23.9782
R123 VP.n85 VP.n84 18.1061
R124 VP.n110 VP.n109 18.1061
R125 VP.n55 VP.n54 18.1061
R126 VP.n30 VP.n29 18.1061
R127 VP.n97 VP.n96 12.234
R128 VP.n98 VP.n97 12.234
R129 VP.n42 VP.n41 12.234
R130 VP.n43 VP.n42 12.234
R131 VP.n84 VP.n83 6.36192
R132 VP.n111 VP.n110 6.36192
R133 VP.n56 VP.n55 6.36192
R134 VP.n31 VP.n28 2.54561
R135 VP.n69 VP.n16 0.417535
R136 VP.n73 VP.n70 0.417535
R137 VP.n124 VP.n0 0.417535
R138 VP VP.n124 0.394291
R139 VP.n32 VP.n31 0.189894
R140 VP.n33 VP.n32 0.189894
R141 VP.n33 VP.n26 0.189894
R142 VP.n37 VP.n26 0.189894
R143 VP.n38 VP.n37 0.189894
R144 VP.n39 VP.n38 0.189894
R145 VP.n39 VP.n24 0.189894
R146 VP.n44 VP.n24 0.189894
R147 VP.n45 VP.n44 0.189894
R148 VP.n46 VP.n45 0.189894
R149 VP.n46 VP.n22 0.189894
R150 VP.n50 VP.n22 0.189894
R151 VP.n51 VP.n50 0.189894
R152 VP.n52 VP.n51 0.189894
R153 VP.n52 VP.n20 0.189894
R154 VP.n57 VP.n20 0.189894
R155 VP.n58 VP.n57 0.189894
R156 VP.n59 VP.n58 0.189894
R157 VP.n59 VP.n18 0.189894
R158 VP.n63 VP.n18 0.189894
R159 VP.n64 VP.n63 0.189894
R160 VP.n65 VP.n64 0.189894
R161 VP.n65 VP.n16 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n75 VP.n74 0.189894
R164 VP.n75 VP.n14 0.189894
R165 VP.n79 VP.n14 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n81 VP.n80 0.189894
R168 VP.n81 VP.n12 0.189894
R169 VP.n86 VP.n12 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n88 VP.n87 0.189894
R172 VP.n88 VP.n10 0.189894
R173 VP.n92 VP.n10 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n94 VP.n93 0.189894
R176 VP.n94 VP.n8 0.189894
R177 VP.n99 VP.n8 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n101 VP.n100 0.189894
R180 VP.n101 VP.n6 0.189894
R181 VP.n105 VP.n6 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n107 VP.n106 0.189894
R184 VP.n107 VP.n4 0.189894
R185 VP.n112 VP.n4 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n114 VP.n113 0.189894
R188 VP.n114 VP.n2 0.189894
R189 VP.n118 VP.n2 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n120 VP.n119 0.189894
R192 VP.n120 VP.n0 0.189894
R193 VTAIL.n11 VTAIL.t5 98.921
R194 VTAIL.n17 VTAIL.t6 98.9207
R195 VTAIL.n2 VTAIL.t15 98.9207
R196 VTAIL.n16 VTAIL.t9 98.9207
R197 VTAIL.n15 VTAIL.n14 91.126
R198 VTAIL.n13 VTAIL.n12 91.126
R199 VTAIL.n10 VTAIL.n9 91.126
R200 VTAIL.n8 VTAIL.n7 91.126
R201 VTAIL.n19 VTAIL.n18 91.1258
R202 VTAIL.n1 VTAIL.n0 91.1258
R203 VTAIL.n4 VTAIL.n3 91.1258
R204 VTAIL.n6 VTAIL.n5 91.1258
R205 VTAIL.n8 VTAIL.n6 23.0652
R206 VTAIL.n17 VTAIL.n16 19.5134
R207 VTAIL.n18 VTAIL.t1 7.79546
R208 VTAIL.n18 VTAIL.t4 7.79546
R209 VTAIL.n0 VTAIL.t3 7.79546
R210 VTAIL.n0 VTAIL.t8 7.79546
R211 VTAIL.n3 VTAIL.t11 7.79546
R212 VTAIL.n3 VTAIL.t14 7.79546
R213 VTAIL.n5 VTAIL.t18 7.79546
R214 VTAIL.n5 VTAIL.t17 7.79546
R215 VTAIL.n14 VTAIL.t13 7.79546
R216 VTAIL.n14 VTAIL.t16 7.79546
R217 VTAIL.n12 VTAIL.t10 7.79546
R218 VTAIL.n12 VTAIL.t12 7.79546
R219 VTAIL.n9 VTAIL.t19 7.79546
R220 VTAIL.n9 VTAIL.t0 7.79546
R221 VTAIL.n7 VTAIL.t2 7.79546
R222 VTAIL.n7 VTAIL.t7 7.79546
R223 VTAIL.n10 VTAIL.n8 3.55222
R224 VTAIL.n11 VTAIL.n10 3.55222
R225 VTAIL.n15 VTAIL.n13 3.55222
R226 VTAIL.n16 VTAIL.n15 3.55222
R227 VTAIL.n6 VTAIL.n4 3.55222
R228 VTAIL.n4 VTAIL.n2 3.55222
R229 VTAIL.n19 VTAIL.n17 3.55222
R230 VTAIL VTAIL.n1 2.72248
R231 VTAIL.n13 VTAIL.n11 2.24619
R232 VTAIL.n2 VTAIL.n1 2.24619
R233 VTAIL VTAIL.n19 0.830241
R234 VDD1.n1 VDD1.t5 119.151
R235 VDD1.n3 VDD1.t8 119.151
R236 VDD1.n5 VDD1.n4 110.413
R237 VDD1.n1 VDD1.n0 107.805
R238 VDD1.n7 VDD1.n6 107.805
R239 VDD1.n3 VDD1.n2 107.805
R240 VDD1.n7 VDD1.n5 46.5397
R241 VDD1.n6 VDD1.t6 7.79546
R242 VDD1.n6 VDD1.t0 7.79546
R243 VDD1.n0 VDD1.t7 7.79546
R244 VDD1.n0 VDD1.t1 7.79546
R245 VDD1.n4 VDD1.t3 7.79546
R246 VDD1.n4 VDD1.t9 7.79546
R247 VDD1.n2 VDD1.t4 7.79546
R248 VDD1.n2 VDD1.t2 7.79546
R249 VDD1 VDD1.n7 2.6061
R250 VDD1 VDD1.n1 0.946621
R251 VDD1.n5 VDD1.n3 0.833085
R252 VN.n105 VN.n54 161.3
R253 VN.n104 VN.n103 161.3
R254 VN.n102 VN.n55 161.3
R255 VN.n101 VN.n100 161.3
R256 VN.n99 VN.n56 161.3
R257 VN.n98 VN.n97 161.3
R258 VN.n96 VN.n57 161.3
R259 VN.n95 VN.n94 161.3
R260 VN.n92 VN.n58 161.3
R261 VN.n91 VN.n90 161.3
R262 VN.n89 VN.n59 161.3
R263 VN.n88 VN.n87 161.3
R264 VN.n86 VN.n60 161.3
R265 VN.n85 VN.n84 161.3
R266 VN.n83 VN.n61 161.3
R267 VN.n82 VN.n81 161.3
R268 VN.n79 VN.n62 161.3
R269 VN.n78 VN.n77 161.3
R270 VN.n76 VN.n63 161.3
R271 VN.n75 VN.n74 161.3
R272 VN.n73 VN.n64 161.3
R273 VN.n72 VN.n71 161.3
R274 VN.n70 VN.n65 161.3
R275 VN.n69 VN.n68 161.3
R276 VN.n51 VN.n0 161.3
R277 VN.n50 VN.n49 161.3
R278 VN.n48 VN.n1 161.3
R279 VN.n47 VN.n46 161.3
R280 VN.n45 VN.n2 161.3
R281 VN.n44 VN.n43 161.3
R282 VN.n42 VN.n3 161.3
R283 VN.n41 VN.n40 161.3
R284 VN.n38 VN.n4 161.3
R285 VN.n37 VN.n36 161.3
R286 VN.n35 VN.n5 161.3
R287 VN.n34 VN.n33 161.3
R288 VN.n32 VN.n6 161.3
R289 VN.n31 VN.n30 161.3
R290 VN.n29 VN.n7 161.3
R291 VN.n28 VN.n27 161.3
R292 VN.n25 VN.n8 161.3
R293 VN.n24 VN.n23 161.3
R294 VN.n22 VN.n9 161.3
R295 VN.n21 VN.n20 161.3
R296 VN.n19 VN.n10 161.3
R297 VN.n18 VN.n17 161.3
R298 VN.n16 VN.n11 161.3
R299 VN.n15 VN.n14 161.3
R300 VN.n12 VN.t1 58.6172
R301 VN.n66 VN.t4 58.6172
R302 VN.n53 VN.n52 58.2041
R303 VN.n107 VN.n106 58.2041
R304 VN.n13 VN.n12 56.9468
R305 VN.n67 VN.n66 56.9468
R306 VN.n20 VN.n19 56.5193
R307 VN.n33 VN.n32 56.5193
R308 VN.n74 VN.n73 56.5193
R309 VN.n87 VN.n86 56.5193
R310 VN VN.n107 53.9435
R311 VN.n46 VN.n45 47.2923
R312 VN.n100 VN.n99 47.2923
R313 VN.n46 VN.n1 33.6945
R314 VN.n100 VN.n55 33.6945
R315 VN.n13 VN.t7 26.5169
R316 VN.n26 VN.t3 26.5169
R317 VN.n39 VN.t5 26.5169
R318 VN.n52 VN.t9 26.5169
R319 VN.n67 VN.t2 26.5169
R320 VN.n80 VN.t0 26.5169
R321 VN.n93 VN.t8 26.5169
R322 VN.n106 VN.t6 26.5169
R323 VN.n14 VN.n11 24.4675
R324 VN.n18 VN.n11 24.4675
R325 VN.n19 VN.n18 24.4675
R326 VN.n20 VN.n9 24.4675
R327 VN.n24 VN.n9 24.4675
R328 VN.n25 VN.n24 24.4675
R329 VN.n27 VN.n7 24.4675
R330 VN.n31 VN.n7 24.4675
R331 VN.n32 VN.n31 24.4675
R332 VN.n33 VN.n5 24.4675
R333 VN.n37 VN.n5 24.4675
R334 VN.n38 VN.n37 24.4675
R335 VN.n40 VN.n3 24.4675
R336 VN.n44 VN.n3 24.4675
R337 VN.n45 VN.n44 24.4675
R338 VN.n50 VN.n1 24.4675
R339 VN.n51 VN.n50 24.4675
R340 VN.n73 VN.n72 24.4675
R341 VN.n72 VN.n65 24.4675
R342 VN.n68 VN.n65 24.4675
R343 VN.n86 VN.n85 24.4675
R344 VN.n85 VN.n61 24.4675
R345 VN.n81 VN.n61 24.4675
R346 VN.n79 VN.n78 24.4675
R347 VN.n78 VN.n63 24.4675
R348 VN.n74 VN.n63 24.4675
R349 VN.n99 VN.n98 24.4675
R350 VN.n98 VN.n57 24.4675
R351 VN.n94 VN.n57 24.4675
R352 VN.n92 VN.n91 24.4675
R353 VN.n91 VN.n59 24.4675
R354 VN.n87 VN.n59 24.4675
R355 VN.n105 VN.n104 24.4675
R356 VN.n104 VN.n55 24.4675
R357 VN.n52 VN.n51 23.9782
R358 VN.n106 VN.n105 23.9782
R359 VN.n14 VN.n13 18.1061
R360 VN.n39 VN.n38 18.1061
R361 VN.n68 VN.n67 18.1061
R362 VN.n93 VN.n92 18.1061
R363 VN.n26 VN.n25 12.234
R364 VN.n27 VN.n26 12.234
R365 VN.n81 VN.n80 12.234
R366 VN.n80 VN.n79 12.234
R367 VN.n40 VN.n39 6.36192
R368 VN.n94 VN.n93 6.36192
R369 VN.n69 VN.n66 2.54564
R370 VN.n15 VN.n12 2.54564
R371 VN.n107 VN.n54 0.417535
R372 VN.n53 VN.n0 0.417535
R373 VN VN.n53 0.394291
R374 VN.n103 VN.n54 0.189894
R375 VN.n103 VN.n102 0.189894
R376 VN.n102 VN.n101 0.189894
R377 VN.n101 VN.n56 0.189894
R378 VN.n97 VN.n56 0.189894
R379 VN.n97 VN.n96 0.189894
R380 VN.n96 VN.n95 0.189894
R381 VN.n95 VN.n58 0.189894
R382 VN.n90 VN.n58 0.189894
R383 VN.n90 VN.n89 0.189894
R384 VN.n89 VN.n88 0.189894
R385 VN.n88 VN.n60 0.189894
R386 VN.n84 VN.n60 0.189894
R387 VN.n84 VN.n83 0.189894
R388 VN.n83 VN.n82 0.189894
R389 VN.n82 VN.n62 0.189894
R390 VN.n77 VN.n62 0.189894
R391 VN.n77 VN.n76 0.189894
R392 VN.n76 VN.n75 0.189894
R393 VN.n75 VN.n64 0.189894
R394 VN.n71 VN.n64 0.189894
R395 VN.n71 VN.n70 0.189894
R396 VN.n70 VN.n69 0.189894
R397 VN.n16 VN.n15 0.189894
R398 VN.n17 VN.n16 0.189894
R399 VN.n17 VN.n10 0.189894
R400 VN.n21 VN.n10 0.189894
R401 VN.n22 VN.n21 0.189894
R402 VN.n23 VN.n22 0.189894
R403 VN.n23 VN.n8 0.189894
R404 VN.n28 VN.n8 0.189894
R405 VN.n29 VN.n28 0.189894
R406 VN.n30 VN.n29 0.189894
R407 VN.n30 VN.n6 0.189894
R408 VN.n34 VN.n6 0.189894
R409 VN.n35 VN.n34 0.189894
R410 VN.n36 VN.n35 0.189894
R411 VN.n36 VN.n4 0.189894
R412 VN.n41 VN.n4 0.189894
R413 VN.n42 VN.n41 0.189894
R414 VN.n43 VN.n42 0.189894
R415 VN.n43 VN.n2 0.189894
R416 VN.n47 VN.n2 0.189894
R417 VN.n48 VN.n47 0.189894
R418 VN.n49 VN.n48 0.189894
R419 VN.n49 VN.n0 0.189894
R420 VDD2.n1 VDD2.t8 119.151
R421 VDD2.n4 VDD2.t3 115.6
R422 VDD2.n3 VDD2.n2 110.413
R423 VDD2 VDD2.n7 110.41
R424 VDD2.n6 VDD2.n5 107.805
R425 VDD2.n1 VDD2.n0 107.805
R426 VDD2.n4 VDD2.n3 44.1808
R427 VDD2.n7 VDD2.t7 7.79546
R428 VDD2.n7 VDD2.t5 7.79546
R429 VDD2.n5 VDD2.t1 7.79546
R430 VDD2.n5 VDD2.t9 7.79546
R431 VDD2.n2 VDD2.t4 7.79546
R432 VDD2.n2 VDD2.t0 7.79546
R433 VDD2.n0 VDD2.t2 7.79546
R434 VDD2.n0 VDD2.t6 7.79546
R435 VDD2.n6 VDD2.n4 3.55222
R436 VDD2 VDD2.n6 0.946621
R437 VDD2.n3 VDD2.n1 0.833085
R438 B.n657 B.n70 585
R439 B.n659 B.n658 585
R440 B.n660 B.n69 585
R441 B.n662 B.n661 585
R442 B.n663 B.n68 585
R443 B.n665 B.n664 585
R444 B.n666 B.n67 585
R445 B.n668 B.n667 585
R446 B.n669 B.n66 585
R447 B.n671 B.n670 585
R448 B.n672 B.n65 585
R449 B.n674 B.n673 585
R450 B.n675 B.n64 585
R451 B.n677 B.n676 585
R452 B.n678 B.n63 585
R453 B.n680 B.n679 585
R454 B.n681 B.n62 585
R455 B.n683 B.n682 585
R456 B.n684 B.n59 585
R457 B.n687 B.n686 585
R458 B.n688 B.n58 585
R459 B.n690 B.n689 585
R460 B.n691 B.n57 585
R461 B.n693 B.n692 585
R462 B.n694 B.n56 585
R463 B.n696 B.n695 585
R464 B.n697 B.n55 585
R465 B.n699 B.n698 585
R466 B.n701 B.n700 585
R467 B.n702 B.n51 585
R468 B.n704 B.n703 585
R469 B.n705 B.n50 585
R470 B.n707 B.n706 585
R471 B.n708 B.n49 585
R472 B.n710 B.n709 585
R473 B.n711 B.n48 585
R474 B.n713 B.n712 585
R475 B.n714 B.n47 585
R476 B.n716 B.n715 585
R477 B.n717 B.n46 585
R478 B.n719 B.n718 585
R479 B.n720 B.n45 585
R480 B.n722 B.n721 585
R481 B.n723 B.n44 585
R482 B.n725 B.n724 585
R483 B.n726 B.n43 585
R484 B.n728 B.n727 585
R485 B.n656 B.n655 585
R486 B.n654 B.n71 585
R487 B.n653 B.n652 585
R488 B.n651 B.n72 585
R489 B.n650 B.n649 585
R490 B.n648 B.n73 585
R491 B.n647 B.n646 585
R492 B.n645 B.n74 585
R493 B.n644 B.n643 585
R494 B.n642 B.n75 585
R495 B.n641 B.n640 585
R496 B.n639 B.n76 585
R497 B.n638 B.n637 585
R498 B.n636 B.n77 585
R499 B.n635 B.n634 585
R500 B.n633 B.n78 585
R501 B.n632 B.n631 585
R502 B.n630 B.n79 585
R503 B.n629 B.n628 585
R504 B.n627 B.n80 585
R505 B.n626 B.n625 585
R506 B.n624 B.n81 585
R507 B.n623 B.n622 585
R508 B.n621 B.n82 585
R509 B.n620 B.n619 585
R510 B.n618 B.n83 585
R511 B.n617 B.n616 585
R512 B.n615 B.n84 585
R513 B.n614 B.n613 585
R514 B.n612 B.n85 585
R515 B.n611 B.n610 585
R516 B.n609 B.n86 585
R517 B.n608 B.n607 585
R518 B.n606 B.n87 585
R519 B.n605 B.n604 585
R520 B.n603 B.n88 585
R521 B.n602 B.n601 585
R522 B.n600 B.n89 585
R523 B.n599 B.n598 585
R524 B.n597 B.n90 585
R525 B.n596 B.n595 585
R526 B.n594 B.n91 585
R527 B.n593 B.n592 585
R528 B.n591 B.n92 585
R529 B.n590 B.n589 585
R530 B.n588 B.n93 585
R531 B.n587 B.n586 585
R532 B.n585 B.n94 585
R533 B.n584 B.n583 585
R534 B.n582 B.n95 585
R535 B.n581 B.n580 585
R536 B.n579 B.n96 585
R537 B.n578 B.n577 585
R538 B.n576 B.n97 585
R539 B.n575 B.n574 585
R540 B.n573 B.n98 585
R541 B.n572 B.n571 585
R542 B.n570 B.n99 585
R543 B.n569 B.n568 585
R544 B.n567 B.n100 585
R545 B.n566 B.n565 585
R546 B.n564 B.n101 585
R547 B.n563 B.n562 585
R548 B.n561 B.n102 585
R549 B.n560 B.n559 585
R550 B.n558 B.n103 585
R551 B.n557 B.n556 585
R552 B.n555 B.n104 585
R553 B.n554 B.n553 585
R554 B.n552 B.n105 585
R555 B.n551 B.n550 585
R556 B.n549 B.n106 585
R557 B.n548 B.n547 585
R558 B.n546 B.n107 585
R559 B.n545 B.n544 585
R560 B.n543 B.n108 585
R561 B.n542 B.n541 585
R562 B.n540 B.n109 585
R563 B.n539 B.n538 585
R564 B.n537 B.n110 585
R565 B.n536 B.n535 585
R566 B.n534 B.n111 585
R567 B.n533 B.n532 585
R568 B.n531 B.n112 585
R569 B.n530 B.n529 585
R570 B.n528 B.n113 585
R571 B.n527 B.n526 585
R572 B.n525 B.n114 585
R573 B.n524 B.n523 585
R574 B.n522 B.n115 585
R575 B.n521 B.n520 585
R576 B.n519 B.n116 585
R577 B.n518 B.n517 585
R578 B.n516 B.n117 585
R579 B.n515 B.n514 585
R580 B.n513 B.n118 585
R581 B.n512 B.n511 585
R582 B.n510 B.n119 585
R583 B.n509 B.n508 585
R584 B.n507 B.n120 585
R585 B.n506 B.n505 585
R586 B.n504 B.n121 585
R587 B.n503 B.n502 585
R588 B.n501 B.n122 585
R589 B.n500 B.n499 585
R590 B.n498 B.n123 585
R591 B.n497 B.n496 585
R592 B.n495 B.n124 585
R593 B.n494 B.n493 585
R594 B.n492 B.n125 585
R595 B.n491 B.n490 585
R596 B.n489 B.n126 585
R597 B.n488 B.n487 585
R598 B.n486 B.n127 585
R599 B.n485 B.n484 585
R600 B.n483 B.n128 585
R601 B.n482 B.n481 585
R602 B.n480 B.n129 585
R603 B.n479 B.n478 585
R604 B.n477 B.n130 585
R605 B.n476 B.n475 585
R606 B.n474 B.n131 585
R607 B.n473 B.n472 585
R608 B.n471 B.n132 585
R609 B.n470 B.n469 585
R610 B.n468 B.n133 585
R611 B.n467 B.n466 585
R612 B.n465 B.n134 585
R613 B.n464 B.n463 585
R614 B.n462 B.n135 585
R615 B.n461 B.n460 585
R616 B.n459 B.n136 585
R617 B.n458 B.n457 585
R618 B.n456 B.n137 585
R619 B.n455 B.n454 585
R620 B.n453 B.n138 585
R621 B.n452 B.n451 585
R622 B.n450 B.n139 585
R623 B.n449 B.n448 585
R624 B.n447 B.n140 585
R625 B.n446 B.n445 585
R626 B.n444 B.n141 585
R627 B.n443 B.n442 585
R628 B.n441 B.n142 585
R629 B.n440 B.n439 585
R630 B.n438 B.n143 585
R631 B.n437 B.n436 585
R632 B.n435 B.n144 585
R633 B.n434 B.n433 585
R634 B.n432 B.n145 585
R635 B.n431 B.n430 585
R636 B.n429 B.n146 585
R637 B.n428 B.n427 585
R638 B.n426 B.n147 585
R639 B.n425 B.n424 585
R640 B.n423 B.n148 585
R641 B.n422 B.n421 585
R642 B.n420 B.n149 585
R643 B.n419 B.n418 585
R644 B.n417 B.n150 585
R645 B.n416 B.n415 585
R646 B.n414 B.n151 585
R647 B.n413 B.n412 585
R648 B.n341 B.n340 585
R649 B.n342 B.n179 585
R650 B.n344 B.n343 585
R651 B.n345 B.n178 585
R652 B.n347 B.n346 585
R653 B.n348 B.n177 585
R654 B.n350 B.n349 585
R655 B.n351 B.n176 585
R656 B.n353 B.n352 585
R657 B.n354 B.n175 585
R658 B.n356 B.n355 585
R659 B.n357 B.n174 585
R660 B.n359 B.n358 585
R661 B.n360 B.n173 585
R662 B.n362 B.n361 585
R663 B.n363 B.n172 585
R664 B.n365 B.n364 585
R665 B.n366 B.n171 585
R666 B.n368 B.n367 585
R667 B.n370 B.n369 585
R668 B.n371 B.n167 585
R669 B.n373 B.n372 585
R670 B.n374 B.n166 585
R671 B.n376 B.n375 585
R672 B.n377 B.n165 585
R673 B.n379 B.n378 585
R674 B.n380 B.n164 585
R675 B.n382 B.n381 585
R676 B.n384 B.n161 585
R677 B.n386 B.n385 585
R678 B.n387 B.n160 585
R679 B.n389 B.n388 585
R680 B.n390 B.n159 585
R681 B.n392 B.n391 585
R682 B.n393 B.n158 585
R683 B.n395 B.n394 585
R684 B.n396 B.n157 585
R685 B.n398 B.n397 585
R686 B.n399 B.n156 585
R687 B.n401 B.n400 585
R688 B.n402 B.n155 585
R689 B.n404 B.n403 585
R690 B.n405 B.n154 585
R691 B.n407 B.n406 585
R692 B.n408 B.n153 585
R693 B.n410 B.n409 585
R694 B.n411 B.n152 585
R695 B.n339 B.n180 585
R696 B.n338 B.n337 585
R697 B.n336 B.n181 585
R698 B.n335 B.n334 585
R699 B.n333 B.n182 585
R700 B.n332 B.n331 585
R701 B.n330 B.n183 585
R702 B.n329 B.n328 585
R703 B.n327 B.n184 585
R704 B.n326 B.n325 585
R705 B.n324 B.n185 585
R706 B.n323 B.n322 585
R707 B.n321 B.n186 585
R708 B.n320 B.n319 585
R709 B.n318 B.n187 585
R710 B.n317 B.n316 585
R711 B.n315 B.n188 585
R712 B.n314 B.n313 585
R713 B.n312 B.n189 585
R714 B.n311 B.n310 585
R715 B.n309 B.n190 585
R716 B.n308 B.n307 585
R717 B.n306 B.n191 585
R718 B.n305 B.n304 585
R719 B.n303 B.n192 585
R720 B.n302 B.n301 585
R721 B.n300 B.n193 585
R722 B.n299 B.n298 585
R723 B.n297 B.n194 585
R724 B.n296 B.n295 585
R725 B.n294 B.n195 585
R726 B.n293 B.n292 585
R727 B.n291 B.n196 585
R728 B.n290 B.n289 585
R729 B.n288 B.n197 585
R730 B.n287 B.n286 585
R731 B.n285 B.n198 585
R732 B.n284 B.n283 585
R733 B.n282 B.n199 585
R734 B.n281 B.n280 585
R735 B.n279 B.n200 585
R736 B.n278 B.n277 585
R737 B.n276 B.n201 585
R738 B.n275 B.n274 585
R739 B.n273 B.n202 585
R740 B.n272 B.n271 585
R741 B.n270 B.n203 585
R742 B.n269 B.n268 585
R743 B.n267 B.n204 585
R744 B.n266 B.n265 585
R745 B.n264 B.n205 585
R746 B.n263 B.n262 585
R747 B.n261 B.n206 585
R748 B.n260 B.n259 585
R749 B.n258 B.n207 585
R750 B.n257 B.n256 585
R751 B.n255 B.n208 585
R752 B.n254 B.n253 585
R753 B.n252 B.n209 585
R754 B.n251 B.n250 585
R755 B.n249 B.n210 585
R756 B.n248 B.n247 585
R757 B.n246 B.n211 585
R758 B.n245 B.n244 585
R759 B.n243 B.n212 585
R760 B.n242 B.n241 585
R761 B.n240 B.n213 585
R762 B.n239 B.n238 585
R763 B.n237 B.n214 585
R764 B.n236 B.n235 585
R765 B.n234 B.n215 585
R766 B.n233 B.n232 585
R767 B.n231 B.n216 585
R768 B.n230 B.n229 585
R769 B.n228 B.n217 585
R770 B.n227 B.n226 585
R771 B.n225 B.n218 585
R772 B.n224 B.n223 585
R773 B.n222 B.n219 585
R774 B.n221 B.n220 585
R775 B.n2 B.n0 585
R776 B.n849 B.n1 585
R777 B.n848 B.n847 585
R778 B.n846 B.n3 585
R779 B.n845 B.n844 585
R780 B.n843 B.n4 585
R781 B.n842 B.n841 585
R782 B.n840 B.n5 585
R783 B.n839 B.n838 585
R784 B.n837 B.n6 585
R785 B.n836 B.n835 585
R786 B.n834 B.n7 585
R787 B.n833 B.n832 585
R788 B.n831 B.n8 585
R789 B.n830 B.n829 585
R790 B.n828 B.n9 585
R791 B.n827 B.n826 585
R792 B.n825 B.n10 585
R793 B.n824 B.n823 585
R794 B.n822 B.n11 585
R795 B.n821 B.n820 585
R796 B.n819 B.n12 585
R797 B.n818 B.n817 585
R798 B.n816 B.n13 585
R799 B.n815 B.n814 585
R800 B.n813 B.n14 585
R801 B.n812 B.n811 585
R802 B.n810 B.n15 585
R803 B.n809 B.n808 585
R804 B.n807 B.n16 585
R805 B.n806 B.n805 585
R806 B.n804 B.n17 585
R807 B.n803 B.n802 585
R808 B.n801 B.n18 585
R809 B.n800 B.n799 585
R810 B.n798 B.n19 585
R811 B.n797 B.n796 585
R812 B.n795 B.n20 585
R813 B.n794 B.n793 585
R814 B.n792 B.n21 585
R815 B.n791 B.n790 585
R816 B.n789 B.n22 585
R817 B.n788 B.n787 585
R818 B.n786 B.n23 585
R819 B.n785 B.n784 585
R820 B.n783 B.n24 585
R821 B.n782 B.n781 585
R822 B.n780 B.n25 585
R823 B.n779 B.n778 585
R824 B.n777 B.n26 585
R825 B.n776 B.n775 585
R826 B.n774 B.n27 585
R827 B.n773 B.n772 585
R828 B.n771 B.n28 585
R829 B.n770 B.n769 585
R830 B.n768 B.n29 585
R831 B.n767 B.n766 585
R832 B.n765 B.n30 585
R833 B.n764 B.n763 585
R834 B.n762 B.n31 585
R835 B.n761 B.n760 585
R836 B.n759 B.n32 585
R837 B.n758 B.n757 585
R838 B.n756 B.n33 585
R839 B.n755 B.n754 585
R840 B.n753 B.n34 585
R841 B.n752 B.n751 585
R842 B.n750 B.n35 585
R843 B.n749 B.n748 585
R844 B.n747 B.n36 585
R845 B.n746 B.n745 585
R846 B.n744 B.n37 585
R847 B.n743 B.n742 585
R848 B.n741 B.n38 585
R849 B.n740 B.n739 585
R850 B.n738 B.n39 585
R851 B.n737 B.n736 585
R852 B.n735 B.n40 585
R853 B.n734 B.n733 585
R854 B.n732 B.n41 585
R855 B.n731 B.n730 585
R856 B.n729 B.n42 585
R857 B.n851 B.n850 585
R858 B.n340 B.n339 449.257
R859 B.n729 B.n728 449.257
R860 B.n412 B.n411 449.257
R861 B.n657 B.n656 449.257
R862 B.n162 B.t9 235.852
R863 B.n168 B.t3 235.852
R864 B.n52 B.t6 235.852
R865 B.n60 B.t0 235.852
R866 B.n162 B.t11 200.567
R867 B.n60 B.t1 200.567
R868 B.n168 B.t5 200.564
R869 B.n52 B.t7 200.564
R870 B.n339 B.n338 163.367
R871 B.n338 B.n181 163.367
R872 B.n334 B.n181 163.367
R873 B.n334 B.n333 163.367
R874 B.n333 B.n332 163.367
R875 B.n332 B.n183 163.367
R876 B.n328 B.n183 163.367
R877 B.n328 B.n327 163.367
R878 B.n327 B.n326 163.367
R879 B.n326 B.n185 163.367
R880 B.n322 B.n185 163.367
R881 B.n322 B.n321 163.367
R882 B.n321 B.n320 163.367
R883 B.n320 B.n187 163.367
R884 B.n316 B.n187 163.367
R885 B.n316 B.n315 163.367
R886 B.n315 B.n314 163.367
R887 B.n314 B.n189 163.367
R888 B.n310 B.n189 163.367
R889 B.n310 B.n309 163.367
R890 B.n309 B.n308 163.367
R891 B.n308 B.n191 163.367
R892 B.n304 B.n191 163.367
R893 B.n304 B.n303 163.367
R894 B.n303 B.n302 163.367
R895 B.n302 B.n193 163.367
R896 B.n298 B.n193 163.367
R897 B.n298 B.n297 163.367
R898 B.n297 B.n296 163.367
R899 B.n296 B.n195 163.367
R900 B.n292 B.n195 163.367
R901 B.n292 B.n291 163.367
R902 B.n291 B.n290 163.367
R903 B.n290 B.n197 163.367
R904 B.n286 B.n197 163.367
R905 B.n286 B.n285 163.367
R906 B.n285 B.n284 163.367
R907 B.n284 B.n199 163.367
R908 B.n280 B.n199 163.367
R909 B.n280 B.n279 163.367
R910 B.n279 B.n278 163.367
R911 B.n278 B.n201 163.367
R912 B.n274 B.n201 163.367
R913 B.n274 B.n273 163.367
R914 B.n273 B.n272 163.367
R915 B.n272 B.n203 163.367
R916 B.n268 B.n203 163.367
R917 B.n268 B.n267 163.367
R918 B.n267 B.n266 163.367
R919 B.n266 B.n205 163.367
R920 B.n262 B.n205 163.367
R921 B.n262 B.n261 163.367
R922 B.n261 B.n260 163.367
R923 B.n260 B.n207 163.367
R924 B.n256 B.n207 163.367
R925 B.n256 B.n255 163.367
R926 B.n255 B.n254 163.367
R927 B.n254 B.n209 163.367
R928 B.n250 B.n209 163.367
R929 B.n250 B.n249 163.367
R930 B.n249 B.n248 163.367
R931 B.n248 B.n211 163.367
R932 B.n244 B.n211 163.367
R933 B.n244 B.n243 163.367
R934 B.n243 B.n242 163.367
R935 B.n242 B.n213 163.367
R936 B.n238 B.n213 163.367
R937 B.n238 B.n237 163.367
R938 B.n237 B.n236 163.367
R939 B.n236 B.n215 163.367
R940 B.n232 B.n215 163.367
R941 B.n232 B.n231 163.367
R942 B.n231 B.n230 163.367
R943 B.n230 B.n217 163.367
R944 B.n226 B.n217 163.367
R945 B.n226 B.n225 163.367
R946 B.n225 B.n224 163.367
R947 B.n224 B.n219 163.367
R948 B.n220 B.n219 163.367
R949 B.n220 B.n2 163.367
R950 B.n850 B.n2 163.367
R951 B.n850 B.n849 163.367
R952 B.n849 B.n848 163.367
R953 B.n848 B.n3 163.367
R954 B.n844 B.n3 163.367
R955 B.n844 B.n843 163.367
R956 B.n843 B.n842 163.367
R957 B.n842 B.n5 163.367
R958 B.n838 B.n5 163.367
R959 B.n838 B.n837 163.367
R960 B.n837 B.n836 163.367
R961 B.n836 B.n7 163.367
R962 B.n832 B.n7 163.367
R963 B.n832 B.n831 163.367
R964 B.n831 B.n830 163.367
R965 B.n830 B.n9 163.367
R966 B.n826 B.n9 163.367
R967 B.n826 B.n825 163.367
R968 B.n825 B.n824 163.367
R969 B.n824 B.n11 163.367
R970 B.n820 B.n11 163.367
R971 B.n820 B.n819 163.367
R972 B.n819 B.n818 163.367
R973 B.n818 B.n13 163.367
R974 B.n814 B.n13 163.367
R975 B.n814 B.n813 163.367
R976 B.n813 B.n812 163.367
R977 B.n812 B.n15 163.367
R978 B.n808 B.n15 163.367
R979 B.n808 B.n807 163.367
R980 B.n807 B.n806 163.367
R981 B.n806 B.n17 163.367
R982 B.n802 B.n17 163.367
R983 B.n802 B.n801 163.367
R984 B.n801 B.n800 163.367
R985 B.n800 B.n19 163.367
R986 B.n796 B.n19 163.367
R987 B.n796 B.n795 163.367
R988 B.n795 B.n794 163.367
R989 B.n794 B.n21 163.367
R990 B.n790 B.n21 163.367
R991 B.n790 B.n789 163.367
R992 B.n789 B.n788 163.367
R993 B.n788 B.n23 163.367
R994 B.n784 B.n23 163.367
R995 B.n784 B.n783 163.367
R996 B.n783 B.n782 163.367
R997 B.n782 B.n25 163.367
R998 B.n778 B.n25 163.367
R999 B.n778 B.n777 163.367
R1000 B.n777 B.n776 163.367
R1001 B.n776 B.n27 163.367
R1002 B.n772 B.n27 163.367
R1003 B.n772 B.n771 163.367
R1004 B.n771 B.n770 163.367
R1005 B.n770 B.n29 163.367
R1006 B.n766 B.n29 163.367
R1007 B.n766 B.n765 163.367
R1008 B.n765 B.n764 163.367
R1009 B.n764 B.n31 163.367
R1010 B.n760 B.n31 163.367
R1011 B.n760 B.n759 163.367
R1012 B.n759 B.n758 163.367
R1013 B.n758 B.n33 163.367
R1014 B.n754 B.n33 163.367
R1015 B.n754 B.n753 163.367
R1016 B.n753 B.n752 163.367
R1017 B.n752 B.n35 163.367
R1018 B.n748 B.n35 163.367
R1019 B.n748 B.n747 163.367
R1020 B.n747 B.n746 163.367
R1021 B.n746 B.n37 163.367
R1022 B.n742 B.n37 163.367
R1023 B.n742 B.n741 163.367
R1024 B.n741 B.n740 163.367
R1025 B.n740 B.n39 163.367
R1026 B.n736 B.n39 163.367
R1027 B.n736 B.n735 163.367
R1028 B.n735 B.n734 163.367
R1029 B.n734 B.n41 163.367
R1030 B.n730 B.n41 163.367
R1031 B.n730 B.n729 163.367
R1032 B.n340 B.n179 163.367
R1033 B.n344 B.n179 163.367
R1034 B.n345 B.n344 163.367
R1035 B.n346 B.n345 163.367
R1036 B.n346 B.n177 163.367
R1037 B.n350 B.n177 163.367
R1038 B.n351 B.n350 163.367
R1039 B.n352 B.n351 163.367
R1040 B.n352 B.n175 163.367
R1041 B.n356 B.n175 163.367
R1042 B.n357 B.n356 163.367
R1043 B.n358 B.n357 163.367
R1044 B.n358 B.n173 163.367
R1045 B.n362 B.n173 163.367
R1046 B.n363 B.n362 163.367
R1047 B.n364 B.n363 163.367
R1048 B.n364 B.n171 163.367
R1049 B.n368 B.n171 163.367
R1050 B.n369 B.n368 163.367
R1051 B.n369 B.n167 163.367
R1052 B.n373 B.n167 163.367
R1053 B.n374 B.n373 163.367
R1054 B.n375 B.n374 163.367
R1055 B.n375 B.n165 163.367
R1056 B.n379 B.n165 163.367
R1057 B.n380 B.n379 163.367
R1058 B.n381 B.n380 163.367
R1059 B.n381 B.n161 163.367
R1060 B.n386 B.n161 163.367
R1061 B.n387 B.n386 163.367
R1062 B.n388 B.n387 163.367
R1063 B.n388 B.n159 163.367
R1064 B.n392 B.n159 163.367
R1065 B.n393 B.n392 163.367
R1066 B.n394 B.n393 163.367
R1067 B.n394 B.n157 163.367
R1068 B.n398 B.n157 163.367
R1069 B.n399 B.n398 163.367
R1070 B.n400 B.n399 163.367
R1071 B.n400 B.n155 163.367
R1072 B.n404 B.n155 163.367
R1073 B.n405 B.n404 163.367
R1074 B.n406 B.n405 163.367
R1075 B.n406 B.n153 163.367
R1076 B.n410 B.n153 163.367
R1077 B.n411 B.n410 163.367
R1078 B.n412 B.n151 163.367
R1079 B.n416 B.n151 163.367
R1080 B.n417 B.n416 163.367
R1081 B.n418 B.n417 163.367
R1082 B.n418 B.n149 163.367
R1083 B.n422 B.n149 163.367
R1084 B.n423 B.n422 163.367
R1085 B.n424 B.n423 163.367
R1086 B.n424 B.n147 163.367
R1087 B.n428 B.n147 163.367
R1088 B.n429 B.n428 163.367
R1089 B.n430 B.n429 163.367
R1090 B.n430 B.n145 163.367
R1091 B.n434 B.n145 163.367
R1092 B.n435 B.n434 163.367
R1093 B.n436 B.n435 163.367
R1094 B.n436 B.n143 163.367
R1095 B.n440 B.n143 163.367
R1096 B.n441 B.n440 163.367
R1097 B.n442 B.n441 163.367
R1098 B.n442 B.n141 163.367
R1099 B.n446 B.n141 163.367
R1100 B.n447 B.n446 163.367
R1101 B.n448 B.n447 163.367
R1102 B.n448 B.n139 163.367
R1103 B.n452 B.n139 163.367
R1104 B.n453 B.n452 163.367
R1105 B.n454 B.n453 163.367
R1106 B.n454 B.n137 163.367
R1107 B.n458 B.n137 163.367
R1108 B.n459 B.n458 163.367
R1109 B.n460 B.n459 163.367
R1110 B.n460 B.n135 163.367
R1111 B.n464 B.n135 163.367
R1112 B.n465 B.n464 163.367
R1113 B.n466 B.n465 163.367
R1114 B.n466 B.n133 163.367
R1115 B.n470 B.n133 163.367
R1116 B.n471 B.n470 163.367
R1117 B.n472 B.n471 163.367
R1118 B.n472 B.n131 163.367
R1119 B.n476 B.n131 163.367
R1120 B.n477 B.n476 163.367
R1121 B.n478 B.n477 163.367
R1122 B.n478 B.n129 163.367
R1123 B.n482 B.n129 163.367
R1124 B.n483 B.n482 163.367
R1125 B.n484 B.n483 163.367
R1126 B.n484 B.n127 163.367
R1127 B.n488 B.n127 163.367
R1128 B.n489 B.n488 163.367
R1129 B.n490 B.n489 163.367
R1130 B.n490 B.n125 163.367
R1131 B.n494 B.n125 163.367
R1132 B.n495 B.n494 163.367
R1133 B.n496 B.n495 163.367
R1134 B.n496 B.n123 163.367
R1135 B.n500 B.n123 163.367
R1136 B.n501 B.n500 163.367
R1137 B.n502 B.n501 163.367
R1138 B.n502 B.n121 163.367
R1139 B.n506 B.n121 163.367
R1140 B.n507 B.n506 163.367
R1141 B.n508 B.n507 163.367
R1142 B.n508 B.n119 163.367
R1143 B.n512 B.n119 163.367
R1144 B.n513 B.n512 163.367
R1145 B.n514 B.n513 163.367
R1146 B.n514 B.n117 163.367
R1147 B.n518 B.n117 163.367
R1148 B.n519 B.n518 163.367
R1149 B.n520 B.n519 163.367
R1150 B.n520 B.n115 163.367
R1151 B.n524 B.n115 163.367
R1152 B.n525 B.n524 163.367
R1153 B.n526 B.n525 163.367
R1154 B.n526 B.n113 163.367
R1155 B.n530 B.n113 163.367
R1156 B.n531 B.n530 163.367
R1157 B.n532 B.n531 163.367
R1158 B.n532 B.n111 163.367
R1159 B.n536 B.n111 163.367
R1160 B.n537 B.n536 163.367
R1161 B.n538 B.n537 163.367
R1162 B.n538 B.n109 163.367
R1163 B.n542 B.n109 163.367
R1164 B.n543 B.n542 163.367
R1165 B.n544 B.n543 163.367
R1166 B.n544 B.n107 163.367
R1167 B.n548 B.n107 163.367
R1168 B.n549 B.n548 163.367
R1169 B.n550 B.n549 163.367
R1170 B.n550 B.n105 163.367
R1171 B.n554 B.n105 163.367
R1172 B.n555 B.n554 163.367
R1173 B.n556 B.n555 163.367
R1174 B.n556 B.n103 163.367
R1175 B.n560 B.n103 163.367
R1176 B.n561 B.n560 163.367
R1177 B.n562 B.n561 163.367
R1178 B.n562 B.n101 163.367
R1179 B.n566 B.n101 163.367
R1180 B.n567 B.n566 163.367
R1181 B.n568 B.n567 163.367
R1182 B.n568 B.n99 163.367
R1183 B.n572 B.n99 163.367
R1184 B.n573 B.n572 163.367
R1185 B.n574 B.n573 163.367
R1186 B.n574 B.n97 163.367
R1187 B.n578 B.n97 163.367
R1188 B.n579 B.n578 163.367
R1189 B.n580 B.n579 163.367
R1190 B.n580 B.n95 163.367
R1191 B.n584 B.n95 163.367
R1192 B.n585 B.n584 163.367
R1193 B.n586 B.n585 163.367
R1194 B.n586 B.n93 163.367
R1195 B.n590 B.n93 163.367
R1196 B.n591 B.n590 163.367
R1197 B.n592 B.n591 163.367
R1198 B.n592 B.n91 163.367
R1199 B.n596 B.n91 163.367
R1200 B.n597 B.n596 163.367
R1201 B.n598 B.n597 163.367
R1202 B.n598 B.n89 163.367
R1203 B.n602 B.n89 163.367
R1204 B.n603 B.n602 163.367
R1205 B.n604 B.n603 163.367
R1206 B.n604 B.n87 163.367
R1207 B.n608 B.n87 163.367
R1208 B.n609 B.n608 163.367
R1209 B.n610 B.n609 163.367
R1210 B.n610 B.n85 163.367
R1211 B.n614 B.n85 163.367
R1212 B.n615 B.n614 163.367
R1213 B.n616 B.n615 163.367
R1214 B.n616 B.n83 163.367
R1215 B.n620 B.n83 163.367
R1216 B.n621 B.n620 163.367
R1217 B.n622 B.n621 163.367
R1218 B.n622 B.n81 163.367
R1219 B.n626 B.n81 163.367
R1220 B.n627 B.n626 163.367
R1221 B.n628 B.n627 163.367
R1222 B.n628 B.n79 163.367
R1223 B.n632 B.n79 163.367
R1224 B.n633 B.n632 163.367
R1225 B.n634 B.n633 163.367
R1226 B.n634 B.n77 163.367
R1227 B.n638 B.n77 163.367
R1228 B.n639 B.n638 163.367
R1229 B.n640 B.n639 163.367
R1230 B.n640 B.n75 163.367
R1231 B.n644 B.n75 163.367
R1232 B.n645 B.n644 163.367
R1233 B.n646 B.n645 163.367
R1234 B.n646 B.n73 163.367
R1235 B.n650 B.n73 163.367
R1236 B.n651 B.n650 163.367
R1237 B.n652 B.n651 163.367
R1238 B.n652 B.n71 163.367
R1239 B.n656 B.n71 163.367
R1240 B.n728 B.n43 163.367
R1241 B.n724 B.n43 163.367
R1242 B.n724 B.n723 163.367
R1243 B.n723 B.n722 163.367
R1244 B.n722 B.n45 163.367
R1245 B.n718 B.n45 163.367
R1246 B.n718 B.n717 163.367
R1247 B.n717 B.n716 163.367
R1248 B.n716 B.n47 163.367
R1249 B.n712 B.n47 163.367
R1250 B.n712 B.n711 163.367
R1251 B.n711 B.n710 163.367
R1252 B.n710 B.n49 163.367
R1253 B.n706 B.n49 163.367
R1254 B.n706 B.n705 163.367
R1255 B.n705 B.n704 163.367
R1256 B.n704 B.n51 163.367
R1257 B.n700 B.n51 163.367
R1258 B.n700 B.n699 163.367
R1259 B.n699 B.n55 163.367
R1260 B.n695 B.n55 163.367
R1261 B.n695 B.n694 163.367
R1262 B.n694 B.n693 163.367
R1263 B.n693 B.n57 163.367
R1264 B.n689 B.n57 163.367
R1265 B.n689 B.n688 163.367
R1266 B.n688 B.n687 163.367
R1267 B.n687 B.n59 163.367
R1268 B.n682 B.n59 163.367
R1269 B.n682 B.n681 163.367
R1270 B.n681 B.n680 163.367
R1271 B.n680 B.n63 163.367
R1272 B.n676 B.n63 163.367
R1273 B.n676 B.n675 163.367
R1274 B.n675 B.n674 163.367
R1275 B.n674 B.n65 163.367
R1276 B.n670 B.n65 163.367
R1277 B.n670 B.n669 163.367
R1278 B.n669 B.n668 163.367
R1279 B.n668 B.n67 163.367
R1280 B.n664 B.n67 163.367
R1281 B.n664 B.n663 163.367
R1282 B.n663 B.n662 163.367
R1283 B.n662 B.n69 163.367
R1284 B.n658 B.n69 163.367
R1285 B.n658 B.n657 163.367
R1286 B.n163 B.t10 120.665
R1287 B.n61 B.t2 120.665
R1288 B.n169 B.t4 120.66
R1289 B.n53 B.t8 120.66
R1290 B.n163 B.n162 79.9035
R1291 B.n169 B.n168 79.9035
R1292 B.n53 B.n52 79.9035
R1293 B.n61 B.n60 79.9035
R1294 B.n383 B.n163 59.5399
R1295 B.n170 B.n169 59.5399
R1296 B.n54 B.n53 59.5399
R1297 B.n685 B.n61 59.5399
R1298 B.n727 B.n42 29.1907
R1299 B.n413 B.n152 29.1907
R1300 B.n341 B.n180 29.1907
R1301 B.n655 B.n70 29.1907
R1302 B B.n851 18.0485
R1303 B.n727 B.n726 10.6151
R1304 B.n726 B.n725 10.6151
R1305 B.n725 B.n44 10.6151
R1306 B.n721 B.n44 10.6151
R1307 B.n721 B.n720 10.6151
R1308 B.n720 B.n719 10.6151
R1309 B.n719 B.n46 10.6151
R1310 B.n715 B.n46 10.6151
R1311 B.n715 B.n714 10.6151
R1312 B.n714 B.n713 10.6151
R1313 B.n713 B.n48 10.6151
R1314 B.n709 B.n48 10.6151
R1315 B.n709 B.n708 10.6151
R1316 B.n708 B.n707 10.6151
R1317 B.n707 B.n50 10.6151
R1318 B.n703 B.n50 10.6151
R1319 B.n703 B.n702 10.6151
R1320 B.n702 B.n701 10.6151
R1321 B.n698 B.n697 10.6151
R1322 B.n697 B.n696 10.6151
R1323 B.n696 B.n56 10.6151
R1324 B.n692 B.n56 10.6151
R1325 B.n692 B.n691 10.6151
R1326 B.n691 B.n690 10.6151
R1327 B.n690 B.n58 10.6151
R1328 B.n686 B.n58 10.6151
R1329 B.n684 B.n683 10.6151
R1330 B.n683 B.n62 10.6151
R1331 B.n679 B.n62 10.6151
R1332 B.n679 B.n678 10.6151
R1333 B.n678 B.n677 10.6151
R1334 B.n677 B.n64 10.6151
R1335 B.n673 B.n64 10.6151
R1336 B.n673 B.n672 10.6151
R1337 B.n672 B.n671 10.6151
R1338 B.n671 B.n66 10.6151
R1339 B.n667 B.n66 10.6151
R1340 B.n667 B.n666 10.6151
R1341 B.n666 B.n665 10.6151
R1342 B.n665 B.n68 10.6151
R1343 B.n661 B.n68 10.6151
R1344 B.n661 B.n660 10.6151
R1345 B.n660 B.n659 10.6151
R1346 B.n659 B.n70 10.6151
R1347 B.n414 B.n413 10.6151
R1348 B.n415 B.n414 10.6151
R1349 B.n415 B.n150 10.6151
R1350 B.n419 B.n150 10.6151
R1351 B.n420 B.n419 10.6151
R1352 B.n421 B.n420 10.6151
R1353 B.n421 B.n148 10.6151
R1354 B.n425 B.n148 10.6151
R1355 B.n426 B.n425 10.6151
R1356 B.n427 B.n426 10.6151
R1357 B.n427 B.n146 10.6151
R1358 B.n431 B.n146 10.6151
R1359 B.n432 B.n431 10.6151
R1360 B.n433 B.n432 10.6151
R1361 B.n433 B.n144 10.6151
R1362 B.n437 B.n144 10.6151
R1363 B.n438 B.n437 10.6151
R1364 B.n439 B.n438 10.6151
R1365 B.n439 B.n142 10.6151
R1366 B.n443 B.n142 10.6151
R1367 B.n444 B.n443 10.6151
R1368 B.n445 B.n444 10.6151
R1369 B.n445 B.n140 10.6151
R1370 B.n449 B.n140 10.6151
R1371 B.n450 B.n449 10.6151
R1372 B.n451 B.n450 10.6151
R1373 B.n451 B.n138 10.6151
R1374 B.n455 B.n138 10.6151
R1375 B.n456 B.n455 10.6151
R1376 B.n457 B.n456 10.6151
R1377 B.n457 B.n136 10.6151
R1378 B.n461 B.n136 10.6151
R1379 B.n462 B.n461 10.6151
R1380 B.n463 B.n462 10.6151
R1381 B.n463 B.n134 10.6151
R1382 B.n467 B.n134 10.6151
R1383 B.n468 B.n467 10.6151
R1384 B.n469 B.n468 10.6151
R1385 B.n469 B.n132 10.6151
R1386 B.n473 B.n132 10.6151
R1387 B.n474 B.n473 10.6151
R1388 B.n475 B.n474 10.6151
R1389 B.n475 B.n130 10.6151
R1390 B.n479 B.n130 10.6151
R1391 B.n480 B.n479 10.6151
R1392 B.n481 B.n480 10.6151
R1393 B.n481 B.n128 10.6151
R1394 B.n485 B.n128 10.6151
R1395 B.n486 B.n485 10.6151
R1396 B.n487 B.n486 10.6151
R1397 B.n487 B.n126 10.6151
R1398 B.n491 B.n126 10.6151
R1399 B.n492 B.n491 10.6151
R1400 B.n493 B.n492 10.6151
R1401 B.n493 B.n124 10.6151
R1402 B.n497 B.n124 10.6151
R1403 B.n498 B.n497 10.6151
R1404 B.n499 B.n498 10.6151
R1405 B.n499 B.n122 10.6151
R1406 B.n503 B.n122 10.6151
R1407 B.n504 B.n503 10.6151
R1408 B.n505 B.n504 10.6151
R1409 B.n505 B.n120 10.6151
R1410 B.n509 B.n120 10.6151
R1411 B.n510 B.n509 10.6151
R1412 B.n511 B.n510 10.6151
R1413 B.n511 B.n118 10.6151
R1414 B.n515 B.n118 10.6151
R1415 B.n516 B.n515 10.6151
R1416 B.n517 B.n516 10.6151
R1417 B.n517 B.n116 10.6151
R1418 B.n521 B.n116 10.6151
R1419 B.n522 B.n521 10.6151
R1420 B.n523 B.n522 10.6151
R1421 B.n523 B.n114 10.6151
R1422 B.n527 B.n114 10.6151
R1423 B.n528 B.n527 10.6151
R1424 B.n529 B.n528 10.6151
R1425 B.n529 B.n112 10.6151
R1426 B.n533 B.n112 10.6151
R1427 B.n534 B.n533 10.6151
R1428 B.n535 B.n534 10.6151
R1429 B.n535 B.n110 10.6151
R1430 B.n539 B.n110 10.6151
R1431 B.n540 B.n539 10.6151
R1432 B.n541 B.n540 10.6151
R1433 B.n541 B.n108 10.6151
R1434 B.n545 B.n108 10.6151
R1435 B.n546 B.n545 10.6151
R1436 B.n547 B.n546 10.6151
R1437 B.n547 B.n106 10.6151
R1438 B.n551 B.n106 10.6151
R1439 B.n552 B.n551 10.6151
R1440 B.n553 B.n552 10.6151
R1441 B.n553 B.n104 10.6151
R1442 B.n557 B.n104 10.6151
R1443 B.n558 B.n557 10.6151
R1444 B.n559 B.n558 10.6151
R1445 B.n559 B.n102 10.6151
R1446 B.n563 B.n102 10.6151
R1447 B.n564 B.n563 10.6151
R1448 B.n565 B.n564 10.6151
R1449 B.n565 B.n100 10.6151
R1450 B.n569 B.n100 10.6151
R1451 B.n570 B.n569 10.6151
R1452 B.n571 B.n570 10.6151
R1453 B.n571 B.n98 10.6151
R1454 B.n575 B.n98 10.6151
R1455 B.n576 B.n575 10.6151
R1456 B.n577 B.n576 10.6151
R1457 B.n577 B.n96 10.6151
R1458 B.n581 B.n96 10.6151
R1459 B.n582 B.n581 10.6151
R1460 B.n583 B.n582 10.6151
R1461 B.n583 B.n94 10.6151
R1462 B.n587 B.n94 10.6151
R1463 B.n588 B.n587 10.6151
R1464 B.n589 B.n588 10.6151
R1465 B.n589 B.n92 10.6151
R1466 B.n593 B.n92 10.6151
R1467 B.n594 B.n593 10.6151
R1468 B.n595 B.n594 10.6151
R1469 B.n595 B.n90 10.6151
R1470 B.n599 B.n90 10.6151
R1471 B.n600 B.n599 10.6151
R1472 B.n601 B.n600 10.6151
R1473 B.n601 B.n88 10.6151
R1474 B.n605 B.n88 10.6151
R1475 B.n606 B.n605 10.6151
R1476 B.n607 B.n606 10.6151
R1477 B.n607 B.n86 10.6151
R1478 B.n611 B.n86 10.6151
R1479 B.n612 B.n611 10.6151
R1480 B.n613 B.n612 10.6151
R1481 B.n613 B.n84 10.6151
R1482 B.n617 B.n84 10.6151
R1483 B.n618 B.n617 10.6151
R1484 B.n619 B.n618 10.6151
R1485 B.n619 B.n82 10.6151
R1486 B.n623 B.n82 10.6151
R1487 B.n624 B.n623 10.6151
R1488 B.n625 B.n624 10.6151
R1489 B.n625 B.n80 10.6151
R1490 B.n629 B.n80 10.6151
R1491 B.n630 B.n629 10.6151
R1492 B.n631 B.n630 10.6151
R1493 B.n631 B.n78 10.6151
R1494 B.n635 B.n78 10.6151
R1495 B.n636 B.n635 10.6151
R1496 B.n637 B.n636 10.6151
R1497 B.n637 B.n76 10.6151
R1498 B.n641 B.n76 10.6151
R1499 B.n642 B.n641 10.6151
R1500 B.n643 B.n642 10.6151
R1501 B.n643 B.n74 10.6151
R1502 B.n647 B.n74 10.6151
R1503 B.n648 B.n647 10.6151
R1504 B.n649 B.n648 10.6151
R1505 B.n649 B.n72 10.6151
R1506 B.n653 B.n72 10.6151
R1507 B.n654 B.n653 10.6151
R1508 B.n655 B.n654 10.6151
R1509 B.n342 B.n341 10.6151
R1510 B.n343 B.n342 10.6151
R1511 B.n343 B.n178 10.6151
R1512 B.n347 B.n178 10.6151
R1513 B.n348 B.n347 10.6151
R1514 B.n349 B.n348 10.6151
R1515 B.n349 B.n176 10.6151
R1516 B.n353 B.n176 10.6151
R1517 B.n354 B.n353 10.6151
R1518 B.n355 B.n354 10.6151
R1519 B.n355 B.n174 10.6151
R1520 B.n359 B.n174 10.6151
R1521 B.n360 B.n359 10.6151
R1522 B.n361 B.n360 10.6151
R1523 B.n361 B.n172 10.6151
R1524 B.n365 B.n172 10.6151
R1525 B.n366 B.n365 10.6151
R1526 B.n367 B.n366 10.6151
R1527 B.n371 B.n370 10.6151
R1528 B.n372 B.n371 10.6151
R1529 B.n372 B.n166 10.6151
R1530 B.n376 B.n166 10.6151
R1531 B.n377 B.n376 10.6151
R1532 B.n378 B.n377 10.6151
R1533 B.n378 B.n164 10.6151
R1534 B.n382 B.n164 10.6151
R1535 B.n385 B.n384 10.6151
R1536 B.n385 B.n160 10.6151
R1537 B.n389 B.n160 10.6151
R1538 B.n390 B.n389 10.6151
R1539 B.n391 B.n390 10.6151
R1540 B.n391 B.n158 10.6151
R1541 B.n395 B.n158 10.6151
R1542 B.n396 B.n395 10.6151
R1543 B.n397 B.n396 10.6151
R1544 B.n397 B.n156 10.6151
R1545 B.n401 B.n156 10.6151
R1546 B.n402 B.n401 10.6151
R1547 B.n403 B.n402 10.6151
R1548 B.n403 B.n154 10.6151
R1549 B.n407 B.n154 10.6151
R1550 B.n408 B.n407 10.6151
R1551 B.n409 B.n408 10.6151
R1552 B.n409 B.n152 10.6151
R1553 B.n337 B.n180 10.6151
R1554 B.n337 B.n336 10.6151
R1555 B.n336 B.n335 10.6151
R1556 B.n335 B.n182 10.6151
R1557 B.n331 B.n182 10.6151
R1558 B.n331 B.n330 10.6151
R1559 B.n330 B.n329 10.6151
R1560 B.n329 B.n184 10.6151
R1561 B.n325 B.n184 10.6151
R1562 B.n325 B.n324 10.6151
R1563 B.n324 B.n323 10.6151
R1564 B.n323 B.n186 10.6151
R1565 B.n319 B.n186 10.6151
R1566 B.n319 B.n318 10.6151
R1567 B.n318 B.n317 10.6151
R1568 B.n317 B.n188 10.6151
R1569 B.n313 B.n188 10.6151
R1570 B.n313 B.n312 10.6151
R1571 B.n312 B.n311 10.6151
R1572 B.n311 B.n190 10.6151
R1573 B.n307 B.n190 10.6151
R1574 B.n307 B.n306 10.6151
R1575 B.n306 B.n305 10.6151
R1576 B.n305 B.n192 10.6151
R1577 B.n301 B.n192 10.6151
R1578 B.n301 B.n300 10.6151
R1579 B.n300 B.n299 10.6151
R1580 B.n299 B.n194 10.6151
R1581 B.n295 B.n194 10.6151
R1582 B.n295 B.n294 10.6151
R1583 B.n294 B.n293 10.6151
R1584 B.n293 B.n196 10.6151
R1585 B.n289 B.n196 10.6151
R1586 B.n289 B.n288 10.6151
R1587 B.n288 B.n287 10.6151
R1588 B.n287 B.n198 10.6151
R1589 B.n283 B.n198 10.6151
R1590 B.n283 B.n282 10.6151
R1591 B.n282 B.n281 10.6151
R1592 B.n281 B.n200 10.6151
R1593 B.n277 B.n200 10.6151
R1594 B.n277 B.n276 10.6151
R1595 B.n276 B.n275 10.6151
R1596 B.n275 B.n202 10.6151
R1597 B.n271 B.n202 10.6151
R1598 B.n271 B.n270 10.6151
R1599 B.n270 B.n269 10.6151
R1600 B.n269 B.n204 10.6151
R1601 B.n265 B.n204 10.6151
R1602 B.n265 B.n264 10.6151
R1603 B.n264 B.n263 10.6151
R1604 B.n263 B.n206 10.6151
R1605 B.n259 B.n206 10.6151
R1606 B.n259 B.n258 10.6151
R1607 B.n258 B.n257 10.6151
R1608 B.n257 B.n208 10.6151
R1609 B.n253 B.n208 10.6151
R1610 B.n253 B.n252 10.6151
R1611 B.n252 B.n251 10.6151
R1612 B.n251 B.n210 10.6151
R1613 B.n247 B.n210 10.6151
R1614 B.n247 B.n246 10.6151
R1615 B.n246 B.n245 10.6151
R1616 B.n245 B.n212 10.6151
R1617 B.n241 B.n212 10.6151
R1618 B.n241 B.n240 10.6151
R1619 B.n240 B.n239 10.6151
R1620 B.n239 B.n214 10.6151
R1621 B.n235 B.n214 10.6151
R1622 B.n235 B.n234 10.6151
R1623 B.n234 B.n233 10.6151
R1624 B.n233 B.n216 10.6151
R1625 B.n229 B.n216 10.6151
R1626 B.n229 B.n228 10.6151
R1627 B.n228 B.n227 10.6151
R1628 B.n227 B.n218 10.6151
R1629 B.n223 B.n218 10.6151
R1630 B.n223 B.n222 10.6151
R1631 B.n222 B.n221 10.6151
R1632 B.n221 B.n0 10.6151
R1633 B.n847 B.n1 10.6151
R1634 B.n847 B.n846 10.6151
R1635 B.n846 B.n845 10.6151
R1636 B.n845 B.n4 10.6151
R1637 B.n841 B.n4 10.6151
R1638 B.n841 B.n840 10.6151
R1639 B.n840 B.n839 10.6151
R1640 B.n839 B.n6 10.6151
R1641 B.n835 B.n6 10.6151
R1642 B.n835 B.n834 10.6151
R1643 B.n834 B.n833 10.6151
R1644 B.n833 B.n8 10.6151
R1645 B.n829 B.n8 10.6151
R1646 B.n829 B.n828 10.6151
R1647 B.n828 B.n827 10.6151
R1648 B.n827 B.n10 10.6151
R1649 B.n823 B.n10 10.6151
R1650 B.n823 B.n822 10.6151
R1651 B.n822 B.n821 10.6151
R1652 B.n821 B.n12 10.6151
R1653 B.n817 B.n12 10.6151
R1654 B.n817 B.n816 10.6151
R1655 B.n816 B.n815 10.6151
R1656 B.n815 B.n14 10.6151
R1657 B.n811 B.n14 10.6151
R1658 B.n811 B.n810 10.6151
R1659 B.n810 B.n809 10.6151
R1660 B.n809 B.n16 10.6151
R1661 B.n805 B.n16 10.6151
R1662 B.n805 B.n804 10.6151
R1663 B.n804 B.n803 10.6151
R1664 B.n803 B.n18 10.6151
R1665 B.n799 B.n18 10.6151
R1666 B.n799 B.n798 10.6151
R1667 B.n798 B.n797 10.6151
R1668 B.n797 B.n20 10.6151
R1669 B.n793 B.n20 10.6151
R1670 B.n793 B.n792 10.6151
R1671 B.n792 B.n791 10.6151
R1672 B.n791 B.n22 10.6151
R1673 B.n787 B.n22 10.6151
R1674 B.n787 B.n786 10.6151
R1675 B.n786 B.n785 10.6151
R1676 B.n785 B.n24 10.6151
R1677 B.n781 B.n24 10.6151
R1678 B.n781 B.n780 10.6151
R1679 B.n780 B.n779 10.6151
R1680 B.n779 B.n26 10.6151
R1681 B.n775 B.n26 10.6151
R1682 B.n775 B.n774 10.6151
R1683 B.n774 B.n773 10.6151
R1684 B.n773 B.n28 10.6151
R1685 B.n769 B.n28 10.6151
R1686 B.n769 B.n768 10.6151
R1687 B.n768 B.n767 10.6151
R1688 B.n767 B.n30 10.6151
R1689 B.n763 B.n30 10.6151
R1690 B.n763 B.n762 10.6151
R1691 B.n762 B.n761 10.6151
R1692 B.n761 B.n32 10.6151
R1693 B.n757 B.n32 10.6151
R1694 B.n757 B.n756 10.6151
R1695 B.n756 B.n755 10.6151
R1696 B.n755 B.n34 10.6151
R1697 B.n751 B.n34 10.6151
R1698 B.n751 B.n750 10.6151
R1699 B.n750 B.n749 10.6151
R1700 B.n749 B.n36 10.6151
R1701 B.n745 B.n36 10.6151
R1702 B.n745 B.n744 10.6151
R1703 B.n744 B.n743 10.6151
R1704 B.n743 B.n38 10.6151
R1705 B.n739 B.n38 10.6151
R1706 B.n739 B.n738 10.6151
R1707 B.n738 B.n737 10.6151
R1708 B.n737 B.n40 10.6151
R1709 B.n733 B.n40 10.6151
R1710 B.n733 B.n732 10.6151
R1711 B.n732 B.n731 10.6151
R1712 B.n731 B.n42 10.6151
R1713 B.n698 B.n54 6.5566
R1714 B.n686 B.n685 6.5566
R1715 B.n370 B.n170 6.5566
R1716 B.n383 B.n382 6.5566
R1717 B.n701 B.n54 4.05904
R1718 B.n685 B.n684 4.05904
R1719 B.n367 B.n170 4.05904
R1720 B.n384 B.n383 4.05904
R1721 B.n851 B.n0 2.81026
R1722 B.n851 B.n1 2.81026
C0 B VDD1 2.30947f
C1 VTAIL w_n5914_n1802# 2.3127f
C2 VDD2 w_n5914_n1802# 2.90862f
C3 VTAIL VP 6.18186f
C4 VDD2 VP 0.739821f
C5 VDD1 VN 0.160302f
C6 VDD2 VTAIL 8.02878f
C7 B w_n5914_n1802# 10.3852f
C8 B VP 2.85914f
C9 B VTAIL 2.26179f
C10 VN w_n5914_n1802# 12.9015f
C11 B VDD2 2.47392f
C12 VDD1 w_n5914_n1802# 2.70358f
C13 VN VP 8.711889f
C14 VDD1 VP 4.88913f
C15 VTAIL VN 6.16754f
C16 VDD1 VTAIL 7.96768f
C17 VDD2 VN 4.31351f
C18 VDD2 VDD1 2.94914f
C19 B VN 1.55182f
C20 VP w_n5914_n1802# 13.6744f
C21 VDD2 VSUBS 2.568357f
C22 VDD1 VSUBS 2.302459f
C23 VTAIL VSUBS 0.77925f
C24 VN VSUBS 9.55648f
C25 VP VSUBS 5.083108f
C26 B VSUBS 5.790497f
C27 w_n5914_n1802# VSUBS 0.134059p
C28 B.n0 VSUBS 0.008326f
C29 B.n1 VSUBS 0.008326f
C30 B.n2 VSUBS 0.013167f
C31 B.n3 VSUBS 0.013167f
C32 B.n4 VSUBS 0.013167f
C33 B.n5 VSUBS 0.013167f
C34 B.n6 VSUBS 0.013167f
C35 B.n7 VSUBS 0.013167f
C36 B.n8 VSUBS 0.013167f
C37 B.n9 VSUBS 0.013167f
C38 B.n10 VSUBS 0.013167f
C39 B.n11 VSUBS 0.013167f
C40 B.n12 VSUBS 0.013167f
C41 B.n13 VSUBS 0.013167f
C42 B.n14 VSUBS 0.013167f
C43 B.n15 VSUBS 0.013167f
C44 B.n16 VSUBS 0.013167f
C45 B.n17 VSUBS 0.013167f
C46 B.n18 VSUBS 0.013167f
C47 B.n19 VSUBS 0.013167f
C48 B.n20 VSUBS 0.013167f
C49 B.n21 VSUBS 0.013167f
C50 B.n22 VSUBS 0.013167f
C51 B.n23 VSUBS 0.013167f
C52 B.n24 VSUBS 0.013167f
C53 B.n25 VSUBS 0.013167f
C54 B.n26 VSUBS 0.013167f
C55 B.n27 VSUBS 0.013167f
C56 B.n28 VSUBS 0.013167f
C57 B.n29 VSUBS 0.013167f
C58 B.n30 VSUBS 0.013167f
C59 B.n31 VSUBS 0.013167f
C60 B.n32 VSUBS 0.013167f
C61 B.n33 VSUBS 0.013167f
C62 B.n34 VSUBS 0.013167f
C63 B.n35 VSUBS 0.013167f
C64 B.n36 VSUBS 0.013167f
C65 B.n37 VSUBS 0.013167f
C66 B.n38 VSUBS 0.013167f
C67 B.n39 VSUBS 0.013167f
C68 B.n40 VSUBS 0.013167f
C69 B.n41 VSUBS 0.013167f
C70 B.n42 VSUBS 0.027914f
C71 B.n43 VSUBS 0.013167f
C72 B.n44 VSUBS 0.013167f
C73 B.n45 VSUBS 0.013167f
C74 B.n46 VSUBS 0.013167f
C75 B.n47 VSUBS 0.013167f
C76 B.n48 VSUBS 0.013167f
C77 B.n49 VSUBS 0.013167f
C78 B.n50 VSUBS 0.013167f
C79 B.n51 VSUBS 0.013167f
C80 B.t8 VSUBS 0.208699f
C81 B.t7 VSUBS 0.256474f
C82 B.t6 VSUBS 1.44579f
C83 B.n52 VSUBS 0.193584f
C84 B.n53 VSUBS 0.1387f
C85 B.n54 VSUBS 0.030505f
C86 B.n55 VSUBS 0.013167f
C87 B.n56 VSUBS 0.013167f
C88 B.n57 VSUBS 0.013167f
C89 B.n58 VSUBS 0.013167f
C90 B.n59 VSUBS 0.013167f
C91 B.t2 VSUBS 0.208699f
C92 B.t1 VSUBS 0.256474f
C93 B.t0 VSUBS 1.44579f
C94 B.n60 VSUBS 0.193585f
C95 B.n61 VSUBS 0.1387f
C96 B.n62 VSUBS 0.013167f
C97 B.n63 VSUBS 0.013167f
C98 B.n64 VSUBS 0.013167f
C99 B.n65 VSUBS 0.013167f
C100 B.n66 VSUBS 0.013167f
C101 B.n67 VSUBS 0.013167f
C102 B.n68 VSUBS 0.013167f
C103 B.n69 VSUBS 0.013167f
C104 B.n70 VSUBS 0.027659f
C105 B.n71 VSUBS 0.013167f
C106 B.n72 VSUBS 0.013167f
C107 B.n73 VSUBS 0.013167f
C108 B.n74 VSUBS 0.013167f
C109 B.n75 VSUBS 0.013167f
C110 B.n76 VSUBS 0.013167f
C111 B.n77 VSUBS 0.013167f
C112 B.n78 VSUBS 0.013167f
C113 B.n79 VSUBS 0.013167f
C114 B.n80 VSUBS 0.013167f
C115 B.n81 VSUBS 0.013167f
C116 B.n82 VSUBS 0.013167f
C117 B.n83 VSUBS 0.013167f
C118 B.n84 VSUBS 0.013167f
C119 B.n85 VSUBS 0.013167f
C120 B.n86 VSUBS 0.013167f
C121 B.n87 VSUBS 0.013167f
C122 B.n88 VSUBS 0.013167f
C123 B.n89 VSUBS 0.013167f
C124 B.n90 VSUBS 0.013167f
C125 B.n91 VSUBS 0.013167f
C126 B.n92 VSUBS 0.013167f
C127 B.n93 VSUBS 0.013167f
C128 B.n94 VSUBS 0.013167f
C129 B.n95 VSUBS 0.013167f
C130 B.n96 VSUBS 0.013167f
C131 B.n97 VSUBS 0.013167f
C132 B.n98 VSUBS 0.013167f
C133 B.n99 VSUBS 0.013167f
C134 B.n100 VSUBS 0.013167f
C135 B.n101 VSUBS 0.013167f
C136 B.n102 VSUBS 0.013167f
C137 B.n103 VSUBS 0.013167f
C138 B.n104 VSUBS 0.013167f
C139 B.n105 VSUBS 0.013167f
C140 B.n106 VSUBS 0.013167f
C141 B.n107 VSUBS 0.013167f
C142 B.n108 VSUBS 0.013167f
C143 B.n109 VSUBS 0.013167f
C144 B.n110 VSUBS 0.013167f
C145 B.n111 VSUBS 0.013167f
C146 B.n112 VSUBS 0.013167f
C147 B.n113 VSUBS 0.013167f
C148 B.n114 VSUBS 0.013167f
C149 B.n115 VSUBS 0.013167f
C150 B.n116 VSUBS 0.013167f
C151 B.n117 VSUBS 0.013167f
C152 B.n118 VSUBS 0.013167f
C153 B.n119 VSUBS 0.013167f
C154 B.n120 VSUBS 0.013167f
C155 B.n121 VSUBS 0.013167f
C156 B.n122 VSUBS 0.013167f
C157 B.n123 VSUBS 0.013167f
C158 B.n124 VSUBS 0.013167f
C159 B.n125 VSUBS 0.013167f
C160 B.n126 VSUBS 0.013167f
C161 B.n127 VSUBS 0.013167f
C162 B.n128 VSUBS 0.013167f
C163 B.n129 VSUBS 0.013167f
C164 B.n130 VSUBS 0.013167f
C165 B.n131 VSUBS 0.013167f
C166 B.n132 VSUBS 0.013167f
C167 B.n133 VSUBS 0.013167f
C168 B.n134 VSUBS 0.013167f
C169 B.n135 VSUBS 0.013167f
C170 B.n136 VSUBS 0.013167f
C171 B.n137 VSUBS 0.013167f
C172 B.n138 VSUBS 0.013167f
C173 B.n139 VSUBS 0.013167f
C174 B.n140 VSUBS 0.013167f
C175 B.n141 VSUBS 0.013167f
C176 B.n142 VSUBS 0.013167f
C177 B.n143 VSUBS 0.013167f
C178 B.n144 VSUBS 0.013167f
C179 B.n145 VSUBS 0.013167f
C180 B.n146 VSUBS 0.013167f
C181 B.n147 VSUBS 0.013167f
C182 B.n148 VSUBS 0.013167f
C183 B.n149 VSUBS 0.013167f
C184 B.n150 VSUBS 0.013167f
C185 B.n151 VSUBS 0.013167f
C186 B.n152 VSUBS 0.029399f
C187 B.n153 VSUBS 0.013167f
C188 B.n154 VSUBS 0.013167f
C189 B.n155 VSUBS 0.013167f
C190 B.n156 VSUBS 0.013167f
C191 B.n157 VSUBS 0.013167f
C192 B.n158 VSUBS 0.013167f
C193 B.n159 VSUBS 0.013167f
C194 B.n160 VSUBS 0.013167f
C195 B.n161 VSUBS 0.013167f
C196 B.t10 VSUBS 0.208699f
C197 B.t11 VSUBS 0.256474f
C198 B.t9 VSUBS 1.44579f
C199 B.n162 VSUBS 0.193585f
C200 B.n163 VSUBS 0.1387f
C201 B.n164 VSUBS 0.013167f
C202 B.n165 VSUBS 0.013167f
C203 B.n166 VSUBS 0.013167f
C204 B.n167 VSUBS 0.013167f
C205 B.t4 VSUBS 0.208699f
C206 B.t5 VSUBS 0.256474f
C207 B.t3 VSUBS 1.44579f
C208 B.n168 VSUBS 0.193584f
C209 B.n169 VSUBS 0.1387f
C210 B.n170 VSUBS 0.030505f
C211 B.n171 VSUBS 0.013167f
C212 B.n172 VSUBS 0.013167f
C213 B.n173 VSUBS 0.013167f
C214 B.n174 VSUBS 0.013167f
C215 B.n175 VSUBS 0.013167f
C216 B.n176 VSUBS 0.013167f
C217 B.n177 VSUBS 0.013167f
C218 B.n178 VSUBS 0.013167f
C219 B.n179 VSUBS 0.013167f
C220 B.n180 VSUBS 0.027914f
C221 B.n181 VSUBS 0.013167f
C222 B.n182 VSUBS 0.013167f
C223 B.n183 VSUBS 0.013167f
C224 B.n184 VSUBS 0.013167f
C225 B.n185 VSUBS 0.013167f
C226 B.n186 VSUBS 0.013167f
C227 B.n187 VSUBS 0.013167f
C228 B.n188 VSUBS 0.013167f
C229 B.n189 VSUBS 0.013167f
C230 B.n190 VSUBS 0.013167f
C231 B.n191 VSUBS 0.013167f
C232 B.n192 VSUBS 0.013167f
C233 B.n193 VSUBS 0.013167f
C234 B.n194 VSUBS 0.013167f
C235 B.n195 VSUBS 0.013167f
C236 B.n196 VSUBS 0.013167f
C237 B.n197 VSUBS 0.013167f
C238 B.n198 VSUBS 0.013167f
C239 B.n199 VSUBS 0.013167f
C240 B.n200 VSUBS 0.013167f
C241 B.n201 VSUBS 0.013167f
C242 B.n202 VSUBS 0.013167f
C243 B.n203 VSUBS 0.013167f
C244 B.n204 VSUBS 0.013167f
C245 B.n205 VSUBS 0.013167f
C246 B.n206 VSUBS 0.013167f
C247 B.n207 VSUBS 0.013167f
C248 B.n208 VSUBS 0.013167f
C249 B.n209 VSUBS 0.013167f
C250 B.n210 VSUBS 0.013167f
C251 B.n211 VSUBS 0.013167f
C252 B.n212 VSUBS 0.013167f
C253 B.n213 VSUBS 0.013167f
C254 B.n214 VSUBS 0.013167f
C255 B.n215 VSUBS 0.013167f
C256 B.n216 VSUBS 0.013167f
C257 B.n217 VSUBS 0.013167f
C258 B.n218 VSUBS 0.013167f
C259 B.n219 VSUBS 0.013167f
C260 B.n220 VSUBS 0.013167f
C261 B.n221 VSUBS 0.013167f
C262 B.n222 VSUBS 0.013167f
C263 B.n223 VSUBS 0.013167f
C264 B.n224 VSUBS 0.013167f
C265 B.n225 VSUBS 0.013167f
C266 B.n226 VSUBS 0.013167f
C267 B.n227 VSUBS 0.013167f
C268 B.n228 VSUBS 0.013167f
C269 B.n229 VSUBS 0.013167f
C270 B.n230 VSUBS 0.013167f
C271 B.n231 VSUBS 0.013167f
C272 B.n232 VSUBS 0.013167f
C273 B.n233 VSUBS 0.013167f
C274 B.n234 VSUBS 0.013167f
C275 B.n235 VSUBS 0.013167f
C276 B.n236 VSUBS 0.013167f
C277 B.n237 VSUBS 0.013167f
C278 B.n238 VSUBS 0.013167f
C279 B.n239 VSUBS 0.013167f
C280 B.n240 VSUBS 0.013167f
C281 B.n241 VSUBS 0.013167f
C282 B.n242 VSUBS 0.013167f
C283 B.n243 VSUBS 0.013167f
C284 B.n244 VSUBS 0.013167f
C285 B.n245 VSUBS 0.013167f
C286 B.n246 VSUBS 0.013167f
C287 B.n247 VSUBS 0.013167f
C288 B.n248 VSUBS 0.013167f
C289 B.n249 VSUBS 0.013167f
C290 B.n250 VSUBS 0.013167f
C291 B.n251 VSUBS 0.013167f
C292 B.n252 VSUBS 0.013167f
C293 B.n253 VSUBS 0.013167f
C294 B.n254 VSUBS 0.013167f
C295 B.n255 VSUBS 0.013167f
C296 B.n256 VSUBS 0.013167f
C297 B.n257 VSUBS 0.013167f
C298 B.n258 VSUBS 0.013167f
C299 B.n259 VSUBS 0.013167f
C300 B.n260 VSUBS 0.013167f
C301 B.n261 VSUBS 0.013167f
C302 B.n262 VSUBS 0.013167f
C303 B.n263 VSUBS 0.013167f
C304 B.n264 VSUBS 0.013167f
C305 B.n265 VSUBS 0.013167f
C306 B.n266 VSUBS 0.013167f
C307 B.n267 VSUBS 0.013167f
C308 B.n268 VSUBS 0.013167f
C309 B.n269 VSUBS 0.013167f
C310 B.n270 VSUBS 0.013167f
C311 B.n271 VSUBS 0.013167f
C312 B.n272 VSUBS 0.013167f
C313 B.n273 VSUBS 0.013167f
C314 B.n274 VSUBS 0.013167f
C315 B.n275 VSUBS 0.013167f
C316 B.n276 VSUBS 0.013167f
C317 B.n277 VSUBS 0.013167f
C318 B.n278 VSUBS 0.013167f
C319 B.n279 VSUBS 0.013167f
C320 B.n280 VSUBS 0.013167f
C321 B.n281 VSUBS 0.013167f
C322 B.n282 VSUBS 0.013167f
C323 B.n283 VSUBS 0.013167f
C324 B.n284 VSUBS 0.013167f
C325 B.n285 VSUBS 0.013167f
C326 B.n286 VSUBS 0.013167f
C327 B.n287 VSUBS 0.013167f
C328 B.n288 VSUBS 0.013167f
C329 B.n289 VSUBS 0.013167f
C330 B.n290 VSUBS 0.013167f
C331 B.n291 VSUBS 0.013167f
C332 B.n292 VSUBS 0.013167f
C333 B.n293 VSUBS 0.013167f
C334 B.n294 VSUBS 0.013167f
C335 B.n295 VSUBS 0.013167f
C336 B.n296 VSUBS 0.013167f
C337 B.n297 VSUBS 0.013167f
C338 B.n298 VSUBS 0.013167f
C339 B.n299 VSUBS 0.013167f
C340 B.n300 VSUBS 0.013167f
C341 B.n301 VSUBS 0.013167f
C342 B.n302 VSUBS 0.013167f
C343 B.n303 VSUBS 0.013167f
C344 B.n304 VSUBS 0.013167f
C345 B.n305 VSUBS 0.013167f
C346 B.n306 VSUBS 0.013167f
C347 B.n307 VSUBS 0.013167f
C348 B.n308 VSUBS 0.013167f
C349 B.n309 VSUBS 0.013167f
C350 B.n310 VSUBS 0.013167f
C351 B.n311 VSUBS 0.013167f
C352 B.n312 VSUBS 0.013167f
C353 B.n313 VSUBS 0.013167f
C354 B.n314 VSUBS 0.013167f
C355 B.n315 VSUBS 0.013167f
C356 B.n316 VSUBS 0.013167f
C357 B.n317 VSUBS 0.013167f
C358 B.n318 VSUBS 0.013167f
C359 B.n319 VSUBS 0.013167f
C360 B.n320 VSUBS 0.013167f
C361 B.n321 VSUBS 0.013167f
C362 B.n322 VSUBS 0.013167f
C363 B.n323 VSUBS 0.013167f
C364 B.n324 VSUBS 0.013167f
C365 B.n325 VSUBS 0.013167f
C366 B.n326 VSUBS 0.013167f
C367 B.n327 VSUBS 0.013167f
C368 B.n328 VSUBS 0.013167f
C369 B.n329 VSUBS 0.013167f
C370 B.n330 VSUBS 0.013167f
C371 B.n331 VSUBS 0.013167f
C372 B.n332 VSUBS 0.013167f
C373 B.n333 VSUBS 0.013167f
C374 B.n334 VSUBS 0.013167f
C375 B.n335 VSUBS 0.013167f
C376 B.n336 VSUBS 0.013167f
C377 B.n337 VSUBS 0.013167f
C378 B.n338 VSUBS 0.013167f
C379 B.n339 VSUBS 0.027914f
C380 B.n340 VSUBS 0.029399f
C381 B.n341 VSUBS 0.029399f
C382 B.n342 VSUBS 0.013167f
C383 B.n343 VSUBS 0.013167f
C384 B.n344 VSUBS 0.013167f
C385 B.n345 VSUBS 0.013167f
C386 B.n346 VSUBS 0.013167f
C387 B.n347 VSUBS 0.013167f
C388 B.n348 VSUBS 0.013167f
C389 B.n349 VSUBS 0.013167f
C390 B.n350 VSUBS 0.013167f
C391 B.n351 VSUBS 0.013167f
C392 B.n352 VSUBS 0.013167f
C393 B.n353 VSUBS 0.013167f
C394 B.n354 VSUBS 0.013167f
C395 B.n355 VSUBS 0.013167f
C396 B.n356 VSUBS 0.013167f
C397 B.n357 VSUBS 0.013167f
C398 B.n358 VSUBS 0.013167f
C399 B.n359 VSUBS 0.013167f
C400 B.n360 VSUBS 0.013167f
C401 B.n361 VSUBS 0.013167f
C402 B.n362 VSUBS 0.013167f
C403 B.n363 VSUBS 0.013167f
C404 B.n364 VSUBS 0.013167f
C405 B.n365 VSUBS 0.013167f
C406 B.n366 VSUBS 0.013167f
C407 B.n367 VSUBS 0.0091f
C408 B.n368 VSUBS 0.013167f
C409 B.n369 VSUBS 0.013167f
C410 B.n370 VSUBS 0.010649f
C411 B.n371 VSUBS 0.013167f
C412 B.n372 VSUBS 0.013167f
C413 B.n373 VSUBS 0.013167f
C414 B.n374 VSUBS 0.013167f
C415 B.n375 VSUBS 0.013167f
C416 B.n376 VSUBS 0.013167f
C417 B.n377 VSUBS 0.013167f
C418 B.n378 VSUBS 0.013167f
C419 B.n379 VSUBS 0.013167f
C420 B.n380 VSUBS 0.013167f
C421 B.n381 VSUBS 0.013167f
C422 B.n382 VSUBS 0.010649f
C423 B.n383 VSUBS 0.030505f
C424 B.n384 VSUBS 0.0091f
C425 B.n385 VSUBS 0.013167f
C426 B.n386 VSUBS 0.013167f
C427 B.n387 VSUBS 0.013167f
C428 B.n388 VSUBS 0.013167f
C429 B.n389 VSUBS 0.013167f
C430 B.n390 VSUBS 0.013167f
C431 B.n391 VSUBS 0.013167f
C432 B.n392 VSUBS 0.013167f
C433 B.n393 VSUBS 0.013167f
C434 B.n394 VSUBS 0.013167f
C435 B.n395 VSUBS 0.013167f
C436 B.n396 VSUBS 0.013167f
C437 B.n397 VSUBS 0.013167f
C438 B.n398 VSUBS 0.013167f
C439 B.n399 VSUBS 0.013167f
C440 B.n400 VSUBS 0.013167f
C441 B.n401 VSUBS 0.013167f
C442 B.n402 VSUBS 0.013167f
C443 B.n403 VSUBS 0.013167f
C444 B.n404 VSUBS 0.013167f
C445 B.n405 VSUBS 0.013167f
C446 B.n406 VSUBS 0.013167f
C447 B.n407 VSUBS 0.013167f
C448 B.n408 VSUBS 0.013167f
C449 B.n409 VSUBS 0.013167f
C450 B.n410 VSUBS 0.013167f
C451 B.n411 VSUBS 0.029399f
C452 B.n412 VSUBS 0.027914f
C453 B.n413 VSUBS 0.027914f
C454 B.n414 VSUBS 0.013167f
C455 B.n415 VSUBS 0.013167f
C456 B.n416 VSUBS 0.013167f
C457 B.n417 VSUBS 0.013167f
C458 B.n418 VSUBS 0.013167f
C459 B.n419 VSUBS 0.013167f
C460 B.n420 VSUBS 0.013167f
C461 B.n421 VSUBS 0.013167f
C462 B.n422 VSUBS 0.013167f
C463 B.n423 VSUBS 0.013167f
C464 B.n424 VSUBS 0.013167f
C465 B.n425 VSUBS 0.013167f
C466 B.n426 VSUBS 0.013167f
C467 B.n427 VSUBS 0.013167f
C468 B.n428 VSUBS 0.013167f
C469 B.n429 VSUBS 0.013167f
C470 B.n430 VSUBS 0.013167f
C471 B.n431 VSUBS 0.013167f
C472 B.n432 VSUBS 0.013167f
C473 B.n433 VSUBS 0.013167f
C474 B.n434 VSUBS 0.013167f
C475 B.n435 VSUBS 0.013167f
C476 B.n436 VSUBS 0.013167f
C477 B.n437 VSUBS 0.013167f
C478 B.n438 VSUBS 0.013167f
C479 B.n439 VSUBS 0.013167f
C480 B.n440 VSUBS 0.013167f
C481 B.n441 VSUBS 0.013167f
C482 B.n442 VSUBS 0.013167f
C483 B.n443 VSUBS 0.013167f
C484 B.n444 VSUBS 0.013167f
C485 B.n445 VSUBS 0.013167f
C486 B.n446 VSUBS 0.013167f
C487 B.n447 VSUBS 0.013167f
C488 B.n448 VSUBS 0.013167f
C489 B.n449 VSUBS 0.013167f
C490 B.n450 VSUBS 0.013167f
C491 B.n451 VSUBS 0.013167f
C492 B.n452 VSUBS 0.013167f
C493 B.n453 VSUBS 0.013167f
C494 B.n454 VSUBS 0.013167f
C495 B.n455 VSUBS 0.013167f
C496 B.n456 VSUBS 0.013167f
C497 B.n457 VSUBS 0.013167f
C498 B.n458 VSUBS 0.013167f
C499 B.n459 VSUBS 0.013167f
C500 B.n460 VSUBS 0.013167f
C501 B.n461 VSUBS 0.013167f
C502 B.n462 VSUBS 0.013167f
C503 B.n463 VSUBS 0.013167f
C504 B.n464 VSUBS 0.013167f
C505 B.n465 VSUBS 0.013167f
C506 B.n466 VSUBS 0.013167f
C507 B.n467 VSUBS 0.013167f
C508 B.n468 VSUBS 0.013167f
C509 B.n469 VSUBS 0.013167f
C510 B.n470 VSUBS 0.013167f
C511 B.n471 VSUBS 0.013167f
C512 B.n472 VSUBS 0.013167f
C513 B.n473 VSUBS 0.013167f
C514 B.n474 VSUBS 0.013167f
C515 B.n475 VSUBS 0.013167f
C516 B.n476 VSUBS 0.013167f
C517 B.n477 VSUBS 0.013167f
C518 B.n478 VSUBS 0.013167f
C519 B.n479 VSUBS 0.013167f
C520 B.n480 VSUBS 0.013167f
C521 B.n481 VSUBS 0.013167f
C522 B.n482 VSUBS 0.013167f
C523 B.n483 VSUBS 0.013167f
C524 B.n484 VSUBS 0.013167f
C525 B.n485 VSUBS 0.013167f
C526 B.n486 VSUBS 0.013167f
C527 B.n487 VSUBS 0.013167f
C528 B.n488 VSUBS 0.013167f
C529 B.n489 VSUBS 0.013167f
C530 B.n490 VSUBS 0.013167f
C531 B.n491 VSUBS 0.013167f
C532 B.n492 VSUBS 0.013167f
C533 B.n493 VSUBS 0.013167f
C534 B.n494 VSUBS 0.013167f
C535 B.n495 VSUBS 0.013167f
C536 B.n496 VSUBS 0.013167f
C537 B.n497 VSUBS 0.013167f
C538 B.n498 VSUBS 0.013167f
C539 B.n499 VSUBS 0.013167f
C540 B.n500 VSUBS 0.013167f
C541 B.n501 VSUBS 0.013167f
C542 B.n502 VSUBS 0.013167f
C543 B.n503 VSUBS 0.013167f
C544 B.n504 VSUBS 0.013167f
C545 B.n505 VSUBS 0.013167f
C546 B.n506 VSUBS 0.013167f
C547 B.n507 VSUBS 0.013167f
C548 B.n508 VSUBS 0.013167f
C549 B.n509 VSUBS 0.013167f
C550 B.n510 VSUBS 0.013167f
C551 B.n511 VSUBS 0.013167f
C552 B.n512 VSUBS 0.013167f
C553 B.n513 VSUBS 0.013167f
C554 B.n514 VSUBS 0.013167f
C555 B.n515 VSUBS 0.013167f
C556 B.n516 VSUBS 0.013167f
C557 B.n517 VSUBS 0.013167f
C558 B.n518 VSUBS 0.013167f
C559 B.n519 VSUBS 0.013167f
C560 B.n520 VSUBS 0.013167f
C561 B.n521 VSUBS 0.013167f
C562 B.n522 VSUBS 0.013167f
C563 B.n523 VSUBS 0.013167f
C564 B.n524 VSUBS 0.013167f
C565 B.n525 VSUBS 0.013167f
C566 B.n526 VSUBS 0.013167f
C567 B.n527 VSUBS 0.013167f
C568 B.n528 VSUBS 0.013167f
C569 B.n529 VSUBS 0.013167f
C570 B.n530 VSUBS 0.013167f
C571 B.n531 VSUBS 0.013167f
C572 B.n532 VSUBS 0.013167f
C573 B.n533 VSUBS 0.013167f
C574 B.n534 VSUBS 0.013167f
C575 B.n535 VSUBS 0.013167f
C576 B.n536 VSUBS 0.013167f
C577 B.n537 VSUBS 0.013167f
C578 B.n538 VSUBS 0.013167f
C579 B.n539 VSUBS 0.013167f
C580 B.n540 VSUBS 0.013167f
C581 B.n541 VSUBS 0.013167f
C582 B.n542 VSUBS 0.013167f
C583 B.n543 VSUBS 0.013167f
C584 B.n544 VSUBS 0.013167f
C585 B.n545 VSUBS 0.013167f
C586 B.n546 VSUBS 0.013167f
C587 B.n547 VSUBS 0.013167f
C588 B.n548 VSUBS 0.013167f
C589 B.n549 VSUBS 0.013167f
C590 B.n550 VSUBS 0.013167f
C591 B.n551 VSUBS 0.013167f
C592 B.n552 VSUBS 0.013167f
C593 B.n553 VSUBS 0.013167f
C594 B.n554 VSUBS 0.013167f
C595 B.n555 VSUBS 0.013167f
C596 B.n556 VSUBS 0.013167f
C597 B.n557 VSUBS 0.013167f
C598 B.n558 VSUBS 0.013167f
C599 B.n559 VSUBS 0.013167f
C600 B.n560 VSUBS 0.013167f
C601 B.n561 VSUBS 0.013167f
C602 B.n562 VSUBS 0.013167f
C603 B.n563 VSUBS 0.013167f
C604 B.n564 VSUBS 0.013167f
C605 B.n565 VSUBS 0.013167f
C606 B.n566 VSUBS 0.013167f
C607 B.n567 VSUBS 0.013167f
C608 B.n568 VSUBS 0.013167f
C609 B.n569 VSUBS 0.013167f
C610 B.n570 VSUBS 0.013167f
C611 B.n571 VSUBS 0.013167f
C612 B.n572 VSUBS 0.013167f
C613 B.n573 VSUBS 0.013167f
C614 B.n574 VSUBS 0.013167f
C615 B.n575 VSUBS 0.013167f
C616 B.n576 VSUBS 0.013167f
C617 B.n577 VSUBS 0.013167f
C618 B.n578 VSUBS 0.013167f
C619 B.n579 VSUBS 0.013167f
C620 B.n580 VSUBS 0.013167f
C621 B.n581 VSUBS 0.013167f
C622 B.n582 VSUBS 0.013167f
C623 B.n583 VSUBS 0.013167f
C624 B.n584 VSUBS 0.013167f
C625 B.n585 VSUBS 0.013167f
C626 B.n586 VSUBS 0.013167f
C627 B.n587 VSUBS 0.013167f
C628 B.n588 VSUBS 0.013167f
C629 B.n589 VSUBS 0.013167f
C630 B.n590 VSUBS 0.013167f
C631 B.n591 VSUBS 0.013167f
C632 B.n592 VSUBS 0.013167f
C633 B.n593 VSUBS 0.013167f
C634 B.n594 VSUBS 0.013167f
C635 B.n595 VSUBS 0.013167f
C636 B.n596 VSUBS 0.013167f
C637 B.n597 VSUBS 0.013167f
C638 B.n598 VSUBS 0.013167f
C639 B.n599 VSUBS 0.013167f
C640 B.n600 VSUBS 0.013167f
C641 B.n601 VSUBS 0.013167f
C642 B.n602 VSUBS 0.013167f
C643 B.n603 VSUBS 0.013167f
C644 B.n604 VSUBS 0.013167f
C645 B.n605 VSUBS 0.013167f
C646 B.n606 VSUBS 0.013167f
C647 B.n607 VSUBS 0.013167f
C648 B.n608 VSUBS 0.013167f
C649 B.n609 VSUBS 0.013167f
C650 B.n610 VSUBS 0.013167f
C651 B.n611 VSUBS 0.013167f
C652 B.n612 VSUBS 0.013167f
C653 B.n613 VSUBS 0.013167f
C654 B.n614 VSUBS 0.013167f
C655 B.n615 VSUBS 0.013167f
C656 B.n616 VSUBS 0.013167f
C657 B.n617 VSUBS 0.013167f
C658 B.n618 VSUBS 0.013167f
C659 B.n619 VSUBS 0.013167f
C660 B.n620 VSUBS 0.013167f
C661 B.n621 VSUBS 0.013167f
C662 B.n622 VSUBS 0.013167f
C663 B.n623 VSUBS 0.013167f
C664 B.n624 VSUBS 0.013167f
C665 B.n625 VSUBS 0.013167f
C666 B.n626 VSUBS 0.013167f
C667 B.n627 VSUBS 0.013167f
C668 B.n628 VSUBS 0.013167f
C669 B.n629 VSUBS 0.013167f
C670 B.n630 VSUBS 0.013167f
C671 B.n631 VSUBS 0.013167f
C672 B.n632 VSUBS 0.013167f
C673 B.n633 VSUBS 0.013167f
C674 B.n634 VSUBS 0.013167f
C675 B.n635 VSUBS 0.013167f
C676 B.n636 VSUBS 0.013167f
C677 B.n637 VSUBS 0.013167f
C678 B.n638 VSUBS 0.013167f
C679 B.n639 VSUBS 0.013167f
C680 B.n640 VSUBS 0.013167f
C681 B.n641 VSUBS 0.013167f
C682 B.n642 VSUBS 0.013167f
C683 B.n643 VSUBS 0.013167f
C684 B.n644 VSUBS 0.013167f
C685 B.n645 VSUBS 0.013167f
C686 B.n646 VSUBS 0.013167f
C687 B.n647 VSUBS 0.013167f
C688 B.n648 VSUBS 0.013167f
C689 B.n649 VSUBS 0.013167f
C690 B.n650 VSUBS 0.013167f
C691 B.n651 VSUBS 0.013167f
C692 B.n652 VSUBS 0.013167f
C693 B.n653 VSUBS 0.013167f
C694 B.n654 VSUBS 0.013167f
C695 B.n655 VSUBS 0.029654f
C696 B.n656 VSUBS 0.027914f
C697 B.n657 VSUBS 0.029399f
C698 B.n658 VSUBS 0.013167f
C699 B.n659 VSUBS 0.013167f
C700 B.n660 VSUBS 0.013167f
C701 B.n661 VSUBS 0.013167f
C702 B.n662 VSUBS 0.013167f
C703 B.n663 VSUBS 0.013167f
C704 B.n664 VSUBS 0.013167f
C705 B.n665 VSUBS 0.013167f
C706 B.n666 VSUBS 0.013167f
C707 B.n667 VSUBS 0.013167f
C708 B.n668 VSUBS 0.013167f
C709 B.n669 VSUBS 0.013167f
C710 B.n670 VSUBS 0.013167f
C711 B.n671 VSUBS 0.013167f
C712 B.n672 VSUBS 0.013167f
C713 B.n673 VSUBS 0.013167f
C714 B.n674 VSUBS 0.013167f
C715 B.n675 VSUBS 0.013167f
C716 B.n676 VSUBS 0.013167f
C717 B.n677 VSUBS 0.013167f
C718 B.n678 VSUBS 0.013167f
C719 B.n679 VSUBS 0.013167f
C720 B.n680 VSUBS 0.013167f
C721 B.n681 VSUBS 0.013167f
C722 B.n682 VSUBS 0.013167f
C723 B.n683 VSUBS 0.013167f
C724 B.n684 VSUBS 0.0091f
C725 B.n685 VSUBS 0.030505f
C726 B.n686 VSUBS 0.010649f
C727 B.n687 VSUBS 0.013167f
C728 B.n688 VSUBS 0.013167f
C729 B.n689 VSUBS 0.013167f
C730 B.n690 VSUBS 0.013167f
C731 B.n691 VSUBS 0.013167f
C732 B.n692 VSUBS 0.013167f
C733 B.n693 VSUBS 0.013167f
C734 B.n694 VSUBS 0.013167f
C735 B.n695 VSUBS 0.013167f
C736 B.n696 VSUBS 0.013167f
C737 B.n697 VSUBS 0.013167f
C738 B.n698 VSUBS 0.010649f
C739 B.n699 VSUBS 0.013167f
C740 B.n700 VSUBS 0.013167f
C741 B.n701 VSUBS 0.0091f
C742 B.n702 VSUBS 0.013167f
C743 B.n703 VSUBS 0.013167f
C744 B.n704 VSUBS 0.013167f
C745 B.n705 VSUBS 0.013167f
C746 B.n706 VSUBS 0.013167f
C747 B.n707 VSUBS 0.013167f
C748 B.n708 VSUBS 0.013167f
C749 B.n709 VSUBS 0.013167f
C750 B.n710 VSUBS 0.013167f
C751 B.n711 VSUBS 0.013167f
C752 B.n712 VSUBS 0.013167f
C753 B.n713 VSUBS 0.013167f
C754 B.n714 VSUBS 0.013167f
C755 B.n715 VSUBS 0.013167f
C756 B.n716 VSUBS 0.013167f
C757 B.n717 VSUBS 0.013167f
C758 B.n718 VSUBS 0.013167f
C759 B.n719 VSUBS 0.013167f
C760 B.n720 VSUBS 0.013167f
C761 B.n721 VSUBS 0.013167f
C762 B.n722 VSUBS 0.013167f
C763 B.n723 VSUBS 0.013167f
C764 B.n724 VSUBS 0.013167f
C765 B.n725 VSUBS 0.013167f
C766 B.n726 VSUBS 0.013167f
C767 B.n727 VSUBS 0.029399f
C768 B.n728 VSUBS 0.029399f
C769 B.n729 VSUBS 0.027914f
C770 B.n730 VSUBS 0.013167f
C771 B.n731 VSUBS 0.013167f
C772 B.n732 VSUBS 0.013167f
C773 B.n733 VSUBS 0.013167f
C774 B.n734 VSUBS 0.013167f
C775 B.n735 VSUBS 0.013167f
C776 B.n736 VSUBS 0.013167f
C777 B.n737 VSUBS 0.013167f
C778 B.n738 VSUBS 0.013167f
C779 B.n739 VSUBS 0.013167f
C780 B.n740 VSUBS 0.013167f
C781 B.n741 VSUBS 0.013167f
C782 B.n742 VSUBS 0.013167f
C783 B.n743 VSUBS 0.013167f
C784 B.n744 VSUBS 0.013167f
C785 B.n745 VSUBS 0.013167f
C786 B.n746 VSUBS 0.013167f
C787 B.n747 VSUBS 0.013167f
C788 B.n748 VSUBS 0.013167f
C789 B.n749 VSUBS 0.013167f
C790 B.n750 VSUBS 0.013167f
C791 B.n751 VSUBS 0.013167f
C792 B.n752 VSUBS 0.013167f
C793 B.n753 VSUBS 0.013167f
C794 B.n754 VSUBS 0.013167f
C795 B.n755 VSUBS 0.013167f
C796 B.n756 VSUBS 0.013167f
C797 B.n757 VSUBS 0.013167f
C798 B.n758 VSUBS 0.013167f
C799 B.n759 VSUBS 0.013167f
C800 B.n760 VSUBS 0.013167f
C801 B.n761 VSUBS 0.013167f
C802 B.n762 VSUBS 0.013167f
C803 B.n763 VSUBS 0.013167f
C804 B.n764 VSUBS 0.013167f
C805 B.n765 VSUBS 0.013167f
C806 B.n766 VSUBS 0.013167f
C807 B.n767 VSUBS 0.013167f
C808 B.n768 VSUBS 0.013167f
C809 B.n769 VSUBS 0.013167f
C810 B.n770 VSUBS 0.013167f
C811 B.n771 VSUBS 0.013167f
C812 B.n772 VSUBS 0.013167f
C813 B.n773 VSUBS 0.013167f
C814 B.n774 VSUBS 0.013167f
C815 B.n775 VSUBS 0.013167f
C816 B.n776 VSUBS 0.013167f
C817 B.n777 VSUBS 0.013167f
C818 B.n778 VSUBS 0.013167f
C819 B.n779 VSUBS 0.013167f
C820 B.n780 VSUBS 0.013167f
C821 B.n781 VSUBS 0.013167f
C822 B.n782 VSUBS 0.013167f
C823 B.n783 VSUBS 0.013167f
C824 B.n784 VSUBS 0.013167f
C825 B.n785 VSUBS 0.013167f
C826 B.n786 VSUBS 0.013167f
C827 B.n787 VSUBS 0.013167f
C828 B.n788 VSUBS 0.013167f
C829 B.n789 VSUBS 0.013167f
C830 B.n790 VSUBS 0.013167f
C831 B.n791 VSUBS 0.013167f
C832 B.n792 VSUBS 0.013167f
C833 B.n793 VSUBS 0.013167f
C834 B.n794 VSUBS 0.013167f
C835 B.n795 VSUBS 0.013167f
C836 B.n796 VSUBS 0.013167f
C837 B.n797 VSUBS 0.013167f
C838 B.n798 VSUBS 0.013167f
C839 B.n799 VSUBS 0.013167f
C840 B.n800 VSUBS 0.013167f
C841 B.n801 VSUBS 0.013167f
C842 B.n802 VSUBS 0.013167f
C843 B.n803 VSUBS 0.013167f
C844 B.n804 VSUBS 0.013167f
C845 B.n805 VSUBS 0.013167f
C846 B.n806 VSUBS 0.013167f
C847 B.n807 VSUBS 0.013167f
C848 B.n808 VSUBS 0.013167f
C849 B.n809 VSUBS 0.013167f
C850 B.n810 VSUBS 0.013167f
C851 B.n811 VSUBS 0.013167f
C852 B.n812 VSUBS 0.013167f
C853 B.n813 VSUBS 0.013167f
C854 B.n814 VSUBS 0.013167f
C855 B.n815 VSUBS 0.013167f
C856 B.n816 VSUBS 0.013167f
C857 B.n817 VSUBS 0.013167f
C858 B.n818 VSUBS 0.013167f
C859 B.n819 VSUBS 0.013167f
C860 B.n820 VSUBS 0.013167f
C861 B.n821 VSUBS 0.013167f
C862 B.n822 VSUBS 0.013167f
C863 B.n823 VSUBS 0.013167f
C864 B.n824 VSUBS 0.013167f
C865 B.n825 VSUBS 0.013167f
C866 B.n826 VSUBS 0.013167f
C867 B.n827 VSUBS 0.013167f
C868 B.n828 VSUBS 0.013167f
C869 B.n829 VSUBS 0.013167f
C870 B.n830 VSUBS 0.013167f
C871 B.n831 VSUBS 0.013167f
C872 B.n832 VSUBS 0.013167f
C873 B.n833 VSUBS 0.013167f
C874 B.n834 VSUBS 0.013167f
C875 B.n835 VSUBS 0.013167f
C876 B.n836 VSUBS 0.013167f
C877 B.n837 VSUBS 0.013167f
C878 B.n838 VSUBS 0.013167f
C879 B.n839 VSUBS 0.013167f
C880 B.n840 VSUBS 0.013167f
C881 B.n841 VSUBS 0.013167f
C882 B.n842 VSUBS 0.013167f
C883 B.n843 VSUBS 0.013167f
C884 B.n844 VSUBS 0.013167f
C885 B.n845 VSUBS 0.013167f
C886 B.n846 VSUBS 0.013167f
C887 B.n847 VSUBS 0.013167f
C888 B.n848 VSUBS 0.013167f
C889 B.n849 VSUBS 0.013167f
C890 B.n850 VSUBS 0.013167f
C891 B.n851 VSUBS 0.029813f
C892 VDD2.t8 VSUBS 1.04888f
C893 VDD2.t2 VSUBS 0.125026f
C894 VDD2.t6 VSUBS 0.125026f
C895 VDD2.n0 VSUBS 0.740835f
C896 VDD2.n1 VSUBS 2.1102f
C897 VDD2.t4 VSUBS 0.125026f
C898 VDD2.t0 VSUBS 0.125026f
C899 VDD2.n2 VSUBS 0.77188f
C900 VDD2.n3 VSUBS 4.86471f
C901 VDD2.t3 VSUBS 1.0173f
C902 VDD2.n4 VSUBS 4.72148f
C903 VDD2.t1 VSUBS 0.125026f
C904 VDD2.t9 VSUBS 0.125026f
C905 VDD2.n5 VSUBS 0.740838f
C906 VDD2.n6 VSUBS 1.09523f
C907 VDD2.t7 VSUBS 0.125026f
C908 VDD2.t5 VSUBS 0.125026f
C909 VDD2.n7 VSUBS 0.77183f
C910 VN.n0 VSUBS 0.067131f
C911 VN.t9 VSUBS 1.45434f
C912 VN.n1 VSUBS 0.072088f
C913 VN.n2 VSUBS 0.035689f
C914 VN.n3 VSUBS 0.066515f
C915 VN.n4 VSUBS 0.035689f
C916 VN.t5 VSUBS 1.45434f
C917 VN.n5 VSUBS 0.066515f
C918 VN.n6 VSUBS 0.035689f
C919 VN.n7 VSUBS 0.066515f
C920 VN.n8 VSUBS 0.035689f
C921 VN.t3 VSUBS 1.45434f
C922 VN.n9 VSUBS 0.066515f
C923 VN.n10 VSUBS 0.035689f
C924 VN.n11 VSUBS 0.066515f
C925 VN.t1 VSUBS 1.91554f
C926 VN.n12 VSUBS 0.700772f
C927 VN.t7 VSUBS 1.45434f
C928 VN.n13 VSUBS 0.696113f
C929 VN.n14 VSUBS 0.057977f
C930 VN.n15 VSUBS 0.461229f
C931 VN.n16 VSUBS 0.035689f
C932 VN.n17 VSUBS 0.035689f
C933 VN.n18 VSUBS 0.066515f
C934 VN.n19 VSUBS 0.046132f
C935 VN.n20 VSUBS 0.058066f
C936 VN.n21 VSUBS 0.035689f
C937 VN.n22 VSUBS 0.035689f
C938 VN.n23 VSUBS 0.035689f
C939 VN.n24 VSUBS 0.066515f
C940 VN.n25 VSUBS 0.050096f
C941 VN.n26 VSUBS 0.559737f
C942 VN.n27 VSUBS 0.050096f
C943 VN.n28 VSUBS 0.035689f
C944 VN.n29 VSUBS 0.035689f
C945 VN.n30 VSUBS 0.035689f
C946 VN.n31 VSUBS 0.066515f
C947 VN.n32 VSUBS 0.058066f
C948 VN.n33 VSUBS 0.046132f
C949 VN.n34 VSUBS 0.035689f
C950 VN.n35 VSUBS 0.035689f
C951 VN.n36 VSUBS 0.035689f
C952 VN.n37 VSUBS 0.066515f
C953 VN.n38 VSUBS 0.057977f
C954 VN.n39 VSUBS 0.559737f
C955 VN.n40 VSUBS 0.042214f
C956 VN.n41 VSUBS 0.035689f
C957 VN.n42 VSUBS 0.035689f
C958 VN.n43 VSUBS 0.035689f
C959 VN.n44 VSUBS 0.066515f
C960 VN.n45 VSUBS 0.067463f
C961 VN.n46 VSUBS 0.031162f
C962 VN.n47 VSUBS 0.035689f
C963 VN.n48 VSUBS 0.035689f
C964 VN.n49 VSUBS 0.035689f
C965 VN.n50 VSUBS 0.066515f
C966 VN.n51 VSUBS 0.065858f
C967 VN.n52 VSUBS 0.720407f
C968 VN.n53 VSUBS 0.103225f
C969 VN.n54 VSUBS 0.067131f
C970 VN.t6 VSUBS 1.45434f
C971 VN.n55 VSUBS 0.072088f
C972 VN.n56 VSUBS 0.035689f
C973 VN.n57 VSUBS 0.066515f
C974 VN.n58 VSUBS 0.035689f
C975 VN.t8 VSUBS 1.45434f
C976 VN.n59 VSUBS 0.066515f
C977 VN.n60 VSUBS 0.035689f
C978 VN.n61 VSUBS 0.066515f
C979 VN.n62 VSUBS 0.035689f
C980 VN.t0 VSUBS 1.45434f
C981 VN.n63 VSUBS 0.066515f
C982 VN.n64 VSUBS 0.035689f
C983 VN.n65 VSUBS 0.066515f
C984 VN.t4 VSUBS 1.91554f
C985 VN.n66 VSUBS 0.700772f
C986 VN.t2 VSUBS 1.45434f
C987 VN.n67 VSUBS 0.696113f
C988 VN.n68 VSUBS 0.057977f
C989 VN.n69 VSUBS 0.461229f
C990 VN.n70 VSUBS 0.035689f
C991 VN.n71 VSUBS 0.035689f
C992 VN.n72 VSUBS 0.066515f
C993 VN.n73 VSUBS 0.046132f
C994 VN.n74 VSUBS 0.058066f
C995 VN.n75 VSUBS 0.035689f
C996 VN.n76 VSUBS 0.035689f
C997 VN.n77 VSUBS 0.035689f
C998 VN.n78 VSUBS 0.066515f
C999 VN.n79 VSUBS 0.050096f
C1000 VN.n80 VSUBS 0.559737f
C1001 VN.n81 VSUBS 0.050096f
C1002 VN.n82 VSUBS 0.035689f
C1003 VN.n83 VSUBS 0.035689f
C1004 VN.n84 VSUBS 0.035689f
C1005 VN.n85 VSUBS 0.066515f
C1006 VN.n86 VSUBS 0.058066f
C1007 VN.n87 VSUBS 0.046132f
C1008 VN.n88 VSUBS 0.035689f
C1009 VN.n89 VSUBS 0.035689f
C1010 VN.n90 VSUBS 0.035689f
C1011 VN.n91 VSUBS 0.066515f
C1012 VN.n92 VSUBS 0.057977f
C1013 VN.n93 VSUBS 0.559737f
C1014 VN.n94 VSUBS 0.042214f
C1015 VN.n95 VSUBS 0.035689f
C1016 VN.n96 VSUBS 0.035689f
C1017 VN.n97 VSUBS 0.035689f
C1018 VN.n98 VSUBS 0.066515f
C1019 VN.n99 VSUBS 0.067463f
C1020 VN.n100 VSUBS 0.031162f
C1021 VN.n101 VSUBS 0.035689f
C1022 VN.n102 VSUBS 0.035689f
C1023 VN.n103 VSUBS 0.035689f
C1024 VN.n104 VSUBS 0.066515f
C1025 VN.n105 VSUBS 0.065858f
C1026 VN.n106 VSUBS 0.720407f
C1027 VN.n107 VSUBS 2.30366f
C1028 VDD1.t5 VSUBS 1.05191f
C1029 VDD1.t7 VSUBS 0.125387f
C1030 VDD1.t1 VSUBS 0.125387f
C1031 VDD1.n0 VSUBS 0.742977f
C1032 VDD1.n1 VSUBS 2.12914f
C1033 VDD1.t8 VSUBS 1.0519f
C1034 VDD1.t4 VSUBS 0.125387f
C1035 VDD1.t2 VSUBS 0.125387f
C1036 VDD1.n2 VSUBS 0.742974f
C1037 VDD1.n3 VSUBS 2.11629f
C1038 VDD1.t3 VSUBS 0.125387f
C1039 VDD1.t9 VSUBS 0.125387f
C1040 VDD1.n4 VSUBS 0.774108f
C1041 VDD1.n5 VSUBS 5.10747f
C1042 VDD1.t6 VSUBS 0.125387f
C1043 VDD1.t0 VSUBS 0.125387f
C1044 VDD1.n6 VSUBS 0.742973f
C1045 VDD1.n7 VSUBS 4.9017f
C1046 VTAIL.t3 VSUBS 0.126366f
C1047 VTAIL.t8 VSUBS 0.126366f
C1048 VTAIL.n0 VSUBS 0.649224f
C1049 VTAIL.n1 VSUBS 1.21245f
C1050 VTAIL.t15 VSUBS 0.925499f
C1051 VTAIL.n2 VSUBS 1.38334f
C1052 VTAIL.t11 VSUBS 0.126366f
C1053 VTAIL.t14 VSUBS 0.126366f
C1054 VTAIL.n3 VSUBS 0.649224f
C1055 VTAIL.n4 VSUBS 1.47636f
C1056 VTAIL.t18 VSUBS 0.126366f
C1057 VTAIL.t17 VSUBS 0.126366f
C1058 VTAIL.n5 VSUBS 0.649224f
C1059 VTAIL.n6 VSUBS 2.88033f
C1060 VTAIL.t2 VSUBS 0.126366f
C1061 VTAIL.t7 VSUBS 0.126366f
C1062 VTAIL.n7 VSUBS 0.649228f
C1063 VTAIL.n8 VSUBS 2.88033f
C1064 VTAIL.t19 VSUBS 0.126366f
C1065 VTAIL.t0 VSUBS 0.126366f
C1066 VTAIL.n9 VSUBS 0.649228f
C1067 VTAIL.n10 VSUBS 1.47635f
C1068 VTAIL.t5 VSUBS 0.925503f
C1069 VTAIL.n11 VSUBS 1.38333f
C1070 VTAIL.t10 VSUBS 0.126366f
C1071 VTAIL.t12 VSUBS 0.126366f
C1072 VTAIL.n12 VSUBS 0.649228f
C1073 VTAIL.n13 VSUBS 1.31497f
C1074 VTAIL.t13 VSUBS 0.126366f
C1075 VTAIL.t16 VSUBS 0.126366f
C1076 VTAIL.n14 VSUBS 0.649228f
C1077 VTAIL.n15 VSUBS 1.47635f
C1078 VTAIL.t9 VSUBS 0.925499f
C1079 VTAIL.n16 VSUBS 2.50982f
C1080 VTAIL.t6 VSUBS 0.925499f
C1081 VTAIL.n17 VSUBS 2.50982f
C1082 VTAIL.t1 VSUBS 0.126366f
C1083 VTAIL.t4 VSUBS 0.126366f
C1084 VTAIL.n18 VSUBS 0.649224f
C1085 VTAIL.n19 VSUBS 1.14002f
C1086 VP.n0 VSUBS 0.076242f
C1087 VP.t0 VSUBS 1.65174f
C1088 VP.n1 VSUBS 0.081873f
C1089 VP.n2 VSUBS 0.040533f
C1090 VP.n3 VSUBS 0.075543f
C1091 VP.n4 VSUBS 0.040533f
C1092 VP.t6 VSUBS 1.65174f
C1093 VP.n5 VSUBS 0.075543f
C1094 VP.n6 VSUBS 0.040533f
C1095 VP.n7 VSUBS 0.075543f
C1096 VP.n8 VSUBS 0.040533f
C1097 VP.t7 VSUBS 1.65174f
C1098 VP.n9 VSUBS 0.075543f
C1099 VP.n10 VSUBS 0.040533f
C1100 VP.n11 VSUBS 0.075543f
C1101 VP.n12 VSUBS 0.040533f
C1102 VP.t5 VSUBS 1.65174f
C1103 VP.n13 VSUBS 0.075543f
C1104 VP.n14 VSUBS 0.040533f
C1105 VP.n15 VSUBS 0.075543f
C1106 VP.n16 VSUBS 0.076242f
C1107 VP.t9 VSUBS 1.65174f
C1108 VP.n17 VSUBS 0.081873f
C1109 VP.n18 VSUBS 0.040533f
C1110 VP.n19 VSUBS 0.075543f
C1111 VP.n20 VSUBS 0.040533f
C1112 VP.t3 VSUBS 1.65174f
C1113 VP.n21 VSUBS 0.075543f
C1114 VP.n22 VSUBS 0.040533f
C1115 VP.n23 VSUBS 0.075543f
C1116 VP.n24 VSUBS 0.040533f
C1117 VP.t8 VSUBS 1.65174f
C1118 VP.n25 VSUBS 0.075543f
C1119 VP.n26 VSUBS 0.040533f
C1120 VP.n27 VSUBS 0.075543f
C1121 VP.t4 VSUBS 2.17553f
C1122 VP.n28 VSUBS 0.795891f
C1123 VP.t2 VSUBS 1.65174f
C1124 VP.n29 VSUBS 0.790597f
C1125 VP.n30 VSUBS 0.065846f
C1126 VP.n31 VSUBS 0.523833f
C1127 VP.n32 VSUBS 0.040533f
C1128 VP.n33 VSUBS 0.040533f
C1129 VP.n34 VSUBS 0.075543f
C1130 VP.n35 VSUBS 0.052394f
C1131 VP.n36 VSUBS 0.065948f
C1132 VP.n37 VSUBS 0.040533f
C1133 VP.n38 VSUBS 0.040533f
C1134 VP.n39 VSUBS 0.040533f
C1135 VP.n40 VSUBS 0.075543f
C1136 VP.n41 VSUBS 0.056895f
C1137 VP.n42 VSUBS 0.635711f
C1138 VP.n43 VSUBS 0.056895f
C1139 VP.n44 VSUBS 0.040533f
C1140 VP.n45 VSUBS 0.040533f
C1141 VP.n46 VSUBS 0.040533f
C1142 VP.n47 VSUBS 0.075543f
C1143 VP.n48 VSUBS 0.065948f
C1144 VP.n49 VSUBS 0.052394f
C1145 VP.n50 VSUBS 0.040533f
C1146 VP.n51 VSUBS 0.040533f
C1147 VP.n52 VSUBS 0.040533f
C1148 VP.n53 VSUBS 0.075543f
C1149 VP.n54 VSUBS 0.065846f
C1150 VP.n55 VSUBS 0.635711f
C1151 VP.n56 VSUBS 0.047944f
C1152 VP.n57 VSUBS 0.040533f
C1153 VP.n58 VSUBS 0.040533f
C1154 VP.n59 VSUBS 0.040533f
C1155 VP.n60 VSUBS 0.075543f
C1156 VP.n61 VSUBS 0.07662f
C1157 VP.n62 VSUBS 0.035392f
C1158 VP.n63 VSUBS 0.040533f
C1159 VP.n64 VSUBS 0.040533f
C1160 VP.n65 VSUBS 0.040533f
C1161 VP.n66 VSUBS 0.075543f
C1162 VP.n67 VSUBS 0.074797f
C1163 VP.n68 VSUBS 0.818189f
C1164 VP.n69 VSUBS 2.60632f
C1165 VP.n70 VSUBS 2.63335f
C1166 VP.t1 VSUBS 1.65174f
C1167 VP.n71 VSUBS 0.818189f
C1168 VP.n72 VSUBS 0.074797f
C1169 VP.n73 VSUBS 0.076242f
C1170 VP.n74 VSUBS 0.040533f
C1171 VP.n75 VSUBS 0.040533f
C1172 VP.n76 VSUBS 0.081873f
C1173 VP.n77 VSUBS 0.035392f
C1174 VP.n78 VSUBS 0.07662f
C1175 VP.n79 VSUBS 0.040533f
C1176 VP.n80 VSUBS 0.040533f
C1177 VP.n81 VSUBS 0.040533f
C1178 VP.n82 VSUBS 0.075543f
C1179 VP.n83 VSUBS 0.047944f
C1180 VP.n84 VSUBS 0.635711f
C1181 VP.n85 VSUBS 0.065846f
C1182 VP.n86 VSUBS 0.040533f
C1183 VP.n87 VSUBS 0.040533f
C1184 VP.n88 VSUBS 0.040533f
C1185 VP.n89 VSUBS 0.075543f
C1186 VP.n90 VSUBS 0.052394f
C1187 VP.n91 VSUBS 0.065948f
C1188 VP.n92 VSUBS 0.040533f
C1189 VP.n93 VSUBS 0.040533f
C1190 VP.n94 VSUBS 0.040533f
C1191 VP.n95 VSUBS 0.075543f
C1192 VP.n96 VSUBS 0.056895f
C1193 VP.n97 VSUBS 0.635711f
C1194 VP.n98 VSUBS 0.056895f
C1195 VP.n99 VSUBS 0.040533f
C1196 VP.n100 VSUBS 0.040533f
C1197 VP.n101 VSUBS 0.040533f
C1198 VP.n102 VSUBS 0.075543f
C1199 VP.n103 VSUBS 0.065948f
C1200 VP.n104 VSUBS 0.052394f
C1201 VP.n105 VSUBS 0.040533f
C1202 VP.n106 VSUBS 0.040533f
C1203 VP.n107 VSUBS 0.040533f
C1204 VP.n108 VSUBS 0.075543f
C1205 VP.n109 VSUBS 0.065846f
C1206 VP.n110 VSUBS 0.635711f
C1207 VP.n111 VSUBS 0.047944f
C1208 VP.n112 VSUBS 0.040533f
C1209 VP.n113 VSUBS 0.040533f
C1210 VP.n114 VSUBS 0.040533f
C1211 VP.n115 VSUBS 0.075543f
C1212 VP.n116 VSUBS 0.07662f
C1213 VP.n117 VSUBS 0.035392f
C1214 VP.n118 VSUBS 0.040533f
C1215 VP.n119 VSUBS 0.040533f
C1216 VP.n120 VSUBS 0.040533f
C1217 VP.n121 VSUBS 0.075543f
C1218 VP.n122 VSUBS 0.074797f
C1219 VP.n123 VSUBS 0.818189f
C1220 VP.n124 VSUBS 0.117236f
.ends

