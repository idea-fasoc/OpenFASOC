* NGSPICE file created from diff_pair_sample_0229.ext - technology: sky130A

.subckt diff_pair_sample_0229 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=0 ps=0 w=8.18 l=1.83
X1 VTAIL.t11 VN.t0 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=1.3497 ps=8.51 w=8.18 l=1.83
X2 VDD1.t5 VP.t0 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=3.1902 ps=17.14 w=8.18 l=1.83
X3 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=1.3497 ps=8.51 w=8.18 l=1.83
X4 VDD1.t3 VP.t2 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=1.3497 ps=8.51 w=8.18 l=1.83
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=0 ps=0 w=8.18 l=1.83
X6 VDD1.t2 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=3.1902 ps=17.14 w=8.18 l=1.83
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=0 ps=0 w=8.18 l=1.83
X8 VDD2.t5 VN.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=1.3497 ps=8.51 w=8.18 l=1.83
X9 VDD2.t4 VN.t2 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=3.1902 ps=17.14 w=8.18 l=1.83
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=0 ps=0 w=8.18 l=1.83
X11 VDD2.t3 VN.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1902 pd=17.14 as=1.3497 ps=8.51 w=8.18 l=1.83
X12 VTAIL.t2 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=1.3497 ps=8.51 w=8.18 l=1.83
X13 VTAIL.t3 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=1.3497 ps=8.51 w=8.18 l=1.83
X14 VTAIL.t7 VN.t4 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=1.3497 ps=8.51 w=8.18 l=1.83
X15 VDD2.t1 VN.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3497 pd=8.51 as=3.1902 ps=17.14 w=8.18 l=1.83
R0 B.n630 B.n629 585
R1 B.n241 B.n98 585
R2 B.n240 B.n239 585
R3 B.n238 B.n237 585
R4 B.n236 B.n235 585
R5 B.n234 B.n233 585
R6 B.n232 B.n231 585
R7 B.n230 B.n229 585
R8 B.n228 B.n227 585
R9 B.n226 B.n225 585
R10 B.n224 B.n223 585
R11 B.n222 B.n221 585
R12 B.n220 B.n219 585
R13 B.n218 B.n217 585
R14 B.n216 B.n215 585
R15 B.n214 B.n213 585
R16 B.n212 B.n211 585
R17 B.n210 B.n209 585
R18 B.n208 B.n207 585
R19 B.n206 B.n205 585
R20 B.n204 B.n203 585
R21 B.n202 B.n201 585
R22 B.n200 B.n199 585
R23 B.n198 B.n197 585
R24 B.n196 B.n195 585
R25 B.n194 B.n193 585
R26 B.n192 B.n191 585
R27 B.n190 B.n189 585
R28 B.n188 B.n187 585
R29 B.n186 B.n185 585
R30 B.n184 B.n183 585
R31 B.n182 B.n181 585
R32 B.n180 B.n179 585
R33 B.n178 B.n177 585
R34 B.n176 B.n175 585
R35 B.n174 B.n173 585
R36 B.n172 B.n171 585
R37 B.n170 B.n169 585
R38 B.n168 B.n167 585
R39 B.n166 B.n165 585
R40 B.n164 B.n163 585
R41 B.n162 B.n161 585
R42 B.n160 B.n159 585
R43 B.n158 B.n157 585
R44 B.n156 B.n155 585
R45 B.n154 B.n153 585
R46 B.n152 B.n151 585
R47 B.n150 B.n149 585
R48 B.n148 B.n147 585
R49 B.n146 B.n145 585
R50 B.n144 B.n143 585
R51 B.n142 B.n141 585
R52 B.n140 B.n139 585
R53 B.n138 B.n137 585
R54 B.n136 B.n135 585
R55 B.n134 B.n133 585
R56 B.n132 B.n131 585
R57 B.n130 B.n129 585
R58 B.n128 B.n127 585
R59 B.n126 B.n125 585
R60 B.n124 B.n123 585
R61 B.n122 B.n121 585
R62 B.n120 B.n119 585
R63 B.n118 B.n117 585
R64 B.n116 B.n115 585
R65 B.n114 B.n113 585
R66 B.n112 B.n111 585
R67 B.n110 B.n109 585
R68 B.n108 B.n107 585
R69 B.n106 B.n105 585
R70 B.n628 B.n63 585
R71 B.n633 B.n63 585
R72 B.n627 B.n62 585
R73 B.n634 B.n62 585
R74 B.n626 B.n625 585
R75 B.n625 B.n58 585
R76 B.n624 B.n57 585
R77 B.n640 B.n57 585
R78 B.n623 B.n56 585
R79 B.n641 B.n56 585
R80 B.n622 B.n55 585
R81 B.n642 B.n55 585
R82 B.n621 B.n620 585
R83 B.n620 B.n54 585
R84 B.n619 B.n50 585
R85 B.n648 B.n50 585
R86 B.n618 B.n49 585
R87 B.n649 B.n49 585
R88 B.n617 B.n48 585
R89 B.n650 B.n48 585
R90 B.n616 B.n615 585
R91 B.n615 B.n44 585
R92 B.n614 B.n43 585
R93 B.n656 B.n43 585
R94 B.n613 B.n42 585
R95 B.n657 B.n42 585
R96 B.n612 B.n41 585
R97 B.n658 B.n41 585
R98 B.n611 B.n610 585
R99 B.n610 B.n37 585
R100 B.n609 B.n36 585
R101 B.n664 B.n36 585
R102 B.n608 B.n35 585
R103 B.n665 B.n35 585
R104 B.n607 B.n34 585
R105 B.n666 B.n34 585
R106 B.n606 B.n605 585
R107 B.n605 B.n30 585
R108 B.n604 B.n29 585
R109 B.n672 B.n29 585
R110 B.n603 B.n28 585
R111 B.n673 B.n28 585
R112 B.n602 B.n27 585
R113 B.n674 B.n27 585
R114 B.n601 B.n600 585
R115 B.n600 B.n26 585
R116 B.n599 B.n22 585
R117 B.n680 B.n22 585
R118 B.n598 B.n21 585
R119 B.n681 B.n21 585
R120 B.n597 B.n20 585
R121 B.n682 B.n20 585
R122 B.n596 B.n595 585
R123 B.n595 B.n16 585
R124 B.n594 B.n15 585
R125 B.n688 B.n15 585
R126 B.n593 B.n14 585
R127 B.n689 B.n14 585
R128 B.n592 B.n13 585
R129 B.n690 B.n13 585
R130 B.n591 B.n590 585
R131 B.n590 B.n12 585
R132 B.n589 B.n588 585
R133 B.n589 B.n8 585
R134 B.n587 B.n7 585
R135 B.n697 B.n7 585
R136 B.n586 B.n6 585
R137 B.n698 B.n6 585
R138 B.n585 B.n5 585
R139 B.n699 B.n5 585
R140 B.n584 B.n583 585
R141 B.n583 B.n4 585
R142 B.n582 B.n242 585
R143 B.n582 B.n581 585
R144 B.n572 B.n243 585
R145 B.n244 B.n243 585
R146 B.n574 B.n573 585
R147 B.n575 B.n574 585
R148 B.n571 B.n248 585
R149 B.n252 B.n248 585
R150 B.n570 B.n569 585
R151 B.n569 B.n568 585
R152 B.n250 B.n249 585
R153 B.n251 B.n250 585
R154 B.n561 B.n560 585
R155 B.n562 B.n561 585
R156 B.n559 B.n257 585
R157 B.n257 B.n256 585
R158 B.n558 B.n557 585
R159 B.n557 B.n556 585
R160 B.n259 B.n258 585
R161 B.n549 B.n259 585
R162 B.n548 B.n547 585
R163 B.n550 B.n548 585
R164 B.n546 B.n264 585
R165 B.n264 B.n263 585
R166 B.n545 B.n544 585
R167 B.n544 B.n543 585
R168 B.n266 B.n265 585
R169 B.n267 B.n266 585
R170 B.n536 B.n535 585
R171 B.n537 B.n536 585
R172 B.n534 B.n271 585
R173 B.n275 B.n271 585
R174 B.n533 B.n532 585
R175 B.n532 B.n531 585
R176 B.n273 B.n272 585
R177 B.n274 B.n273 585
R178 B.n524 B.n523 585
R179 B.n525 B.n524 585
R180 B.n522 B.n280 585
R181 B.n280 B.n279 585
R182 B.n521 B.n520 585
R183 B.n520 B.n519 585
R184 B.n282 B.n281 585
R185 B.n283 B.n282 585
R186 B.n512 B.n511 585
R187 B.n513 B.n512 585
R188 B.n510 B.n288 585
R189 B.n288 B.n287 585
R190 B.n509 B.n508 585
R191 B.n508 B.n507 585
R192 B.n290 B.n289 585
R193 B.n500 B.n290 585
R194 B.n499 B.n498 585
R195 B.n501 B.n499 585
R196 B.n497 B.n295 585
R197 B.n295 B.n294 585
R198 B.n496 B.n495 585
R199 B.n495 B.n494 585
R200 B.n297 B.n296 585
R201 B.n298 B.n297 585
R202 B.n487 B.n486 585
R203 B.n488 B.n487 585
R204 B.n485 B.n303 585
R205 B.n303 B.n302 585
R206 B.n480 B.n479 585
R207 B.n478 B.n340 585
R208 B.n477 B.n339 585
R209 B.n482 B.n339 585
R210 B.n476 B.n475 585
R211 B.n474 B.n473 585
R212 B.n472 B.n471 585
R213 B.n470 B.n469 585
R214 B.n468 B.n467 585
R215 B.n466 B.n465 585
R216 B.n464 B.n463 585
R217 B.n462 B.n461 585
R218 B.n460 B.n459 585
R219 B.n458 B.n457 585
R220 B.n456 B.n455 585
R221 B.n454 B.n453 585
R222 B.n452 B.n451 585
R223 B.n450 B.n449 585
R224 B.n448 B.n447 585
R225 B.n446 B.n445 585
R226 B.n444 B.n443 585
R227 B.n442 B.n441 585
R228 B.n440 B.n439 585
R229 B.n438 B.n437 585
R230 B.n436 B.n435 585
R231 B.n434 B.n433 585
R232 B.n432 B.n431 585
R233 B.n430 B.n429 585
R234 B.n428 B.n427 585
R235 B.n426 B.n425 585
R236 B.n424 B.n423 585
R237 B.n421 B.n420 585
R238 B.n419 B.n418 585
R239 B.n417 B.n416 585
R240 B.n415 B.n414 585
R241 B.n413 B.n412 585
R242 B.n411 B.n410 585
R243 B.n409 B.n408 585
R244 B.n407 B.n406 585
R245 B.n405 B.n404 585
R246 B.n403 B.n402 585
R247 B.n400 B.n399 585
R248 B.n398 B.n397 585
R249 B.n396 B.n395 585
R250 B.n394 B.n393 585
R251 B.n392 B.n391 585
R252 B.n390 B.n389 585
R253 B.n388 B.n387 585
R254 B.n386 B.n385 585
R255 B.n384 B.n383 585
R256 B.n382 B.n381 585
R257 B.n380 B.n379 585
R258 B.n378 B.n377 585
R259 B.n376 B.n375 585
R260 B.n374 B.n373 585
R261 B.n372 B.n371 585
R262 B.n370 B.n369 585
R263 B.n368 B.n367 585
R264 B.n366 B.n365 585
R265 B.n364 B.n363 585
R266 B.n362 B.n361 585
R267 B.n360 B.n359 585
R268 B.n358 B.n357 585
R269 B.n356 B.n355 585
R270 B.n354 B.n353 585
R271 B.n352 B.n351 585
R272 B.n350 B.n349 585
R273 B.n348 B.n347 585
R274 B.n346 B.n345 585
R275 B.n305 B.n304 585
R276 B.n484 B.n483 585
R277 B.n483 B.n482 585
R278 B.n301 B.n300 585
R279 B.n302 B.n301 585
R280 B.n490 B.n489 585
R281 B.n489 B.n488 585
R282 B.n491 B.n299 585
R283 B.n299 B.n298 585
R284 B.n493 B.n492 585
R285 B.n494 B.n493 585
R286 B.n293 B.n292 585
R287 B.n294 B.n293 585
R288 B.n503 B.n502 585
R289 B.n502 B.n501 585
R290 B.n504 B.n291 585
R291 B.n500 B.n291 585
R292 B.n506 B.n505 585
R293 B.n507 B.n506 585
R294 B.n286 B.n285 585
R295 B.n287 B.n286 585
R296 B.n515 B.n514 585
R297 B.n514 B.n513 585
R298 B.n516 B.n284 585
R299 B.n284 B.n283 585
R300 B.n518 B.n517 585
R301 B.n519 B.n518 585
R302 B.n278 B.n277 585
R303 B.n279 B.n278 585
R304 B.n527 B.n526 585
R305 B.n526 B.n525 585
R306 B.n528 B.n276 585
R307 B.n276 B.n274 585
R308 B.n530 B.n529 585
R309 B.n531 B.n530 585
R310 B.n270 B.n269 585
R311 B.n275 B.n270 585
R312 B.n539 B.n538 585
R313 B.n538 B.n537 585
R314 B.n540 B.n268 585
R315 B.n268 B.n267 585
R316 B.n542 B.n541 585
R317 B.n543 B.n542 585
R318 B.n262 B.n261 585
R319 B.n263 B.n262 585
R320 B.n552 B.n551 585
R321 B.n551 B.n550 585
R322 B.n553 B.n260 585
R323 B.n549 B.n260 585
R324 B.n555 B.n554 585
R325 B.n556 B.n555 585
R326 B.n255 B.n254 585
R327 B.n256 B.n255 585
R328 B.n564 B.n563 585
R329 B.n563 B.n562 585
R330 B.n565 B.n253 585
R331 B.n253 B.n251 585
R332 B.n567 B.n566 585
R333 B.n568 B.n567 585
R334 B.n247 B.n246 585
R335 B.n252 B.n247 585
R336 B.n577 B.n576 585
R337 B.n576 B.n575 585
R338 B.n578 B.n245 585
R339 B.n245 B.n244 585
R340 B.n580 B.n579 585
R341 B.n581 B.n580 585
R342 B.n3 B.n0 585
R343 B.n4 B.n3 585
R344 B.n696 B.n1 585
R345 B.n697 B.n696 585
R346 B.n695 B.n694 585
R347 B.n695 B.n8 585
R348 B.n693 B.n9 585
R349 B.n12 B.n9 585
R350 B.n692 B.n691 585
R351 B.n691 B.n690 585
R352 B.n11 B.n10 585
R353 B.n689 B.n11 585
R354 B.n687 B.n686 585
R355 B.n688 B.n687 585
R356 B.n685 B.n17 585
R357 B.n17 B.n16 585
R358 B.n684 B.n683 585
R359 B.n683 B.n682 585
R360 B.n19 B.n18 585
R361 B.n681 B.n19 585
R362 B.n679 B.n678 585
R363 B.n680 B.n679 585
R364 B.n677 B.n23 585
R365 B.n26 B.n23 585
R366 B.n676 B.n675 585
R367 B.n675 B.n674 585
R368 B.n25 B.n24 585
R369 B.n673 B.n25 585
R370 B.n671 B.n670 585
R371 B.n672 B.n671 585
R372 B.n669 B.n31 585
R373 B.n31 B.n30 585
R374 B.n668 B.n667 585
R375 B.n667 B.n666 585
R376 B.n33 B.n32 585
R377 B.n665 B.n33 585
R378 B.n663 B.n662 585
R379 B.n664 B.n663 585
R380 B.n661 B.n38 585
R381 B.n38 B.n37 585
R382 B.n660 B.n659 585
R383 B.n659 B.n658 585
R384 B.n40 B.n39 585
R385 B.n657 B.n40 585
R386 B.n655 B.n654 585
R387 B.n656 B.n655 585
R388 B.n653 B.n45 585
R389 B.n45 B.n44 585
R390 B.n652 B.n651 585
R391 B.n651 B.n650 585
R392 B.n47 B.n46 585
R393 B.n649 B.n47 585
R394 B.n647 B.n646 585
R395 B.n648 B.n647 585
R396 B.n645 B.n51 585
R397 B.n54 B.n51 585
R398 B.n644 B.n643 585
R399 B.n643 B.n642 585
R400 B.n53 B.n52 585
R401 B.n641 B.n53 585
R402 B.n639 B.n638 585
R403 B.n640 B.n639 585
R404 B.n637 B.n59 585
R405 B.n59 B.n58 585
R406 B.n636 B.n635 585
R407 B.n635 B.n634 585
R408 B.n61 B.n60 585
R409 B.n633 B.n61 585
R410 B.n700 B.n699 585
R411 B.n698 B.n2 585
R412 B.n105 B.n61 530.939
R413 B.n630 B.n63 530.939
R414 B.n483 B.n303 530.939
R415 B.n480 B.n301 530.939
R416 B.n102 B.t17 314.214
R417 B.n99 B.t13 314.214
R418 B.n343 B.t10 314.214
R419 B.n341 B.t6 314.214
R420 B.n632 B.n631 256.663
R421 B.n632 B.n97 256.663
R422 B.n632 B.n96 256.663
R423 B.n632 B.n95 256.663
R424 B.n632 B.n94 256.663
R425 B.n632 B.n93 256.663
R426 B.n632 B.n92 256.663
R427 B.n632 B.n91 256.663
R428 B.n632 B.n90 256.663
R429 B.n632 B.n89 256.663
R430 B.n632 B.n88 256.663
R431 B.n632 B.n87 256.663
R432 B.n632 B.n86 256.663
R433 B.n632 B.n85 256.663
R434 B.n632 B.n84 256.663
R435 B.n632 B.n83 256.663
R436 B.n632 B.n82 256.663
R437 B.n632 B.n81 256.663
R438 B.n632 B.n80 256.663
R439 B.n632 B.n79 256.663
R440 B.n632 B.n78 256.663
R441 B.n632 B.n77 256.663
R442 B.n632 B.n76 256.663
R443 B.n632 B.n75 256.663
R444 B.n632 B.n74 256.663
R445 B.n632 B.n73 256.663
R446 B.n632 B.n72 256.663
R447 B.n632 B.n71 256.663
R448 B.n632 B.n70 256.663
R449 B.n632 B.n69 256.663
R450 B.n632 B.n68 256.663
R451 B.n632 B.n67 256.663
R452 B.n632 B.n66 256.663
R453 B.n632 B.n65 256.663
R454 B.n632 B.n64 256.663
R455 B.n482 B.n481 256.663
R456 B.n482 B.n306 256.663
R457 B.n482 B.n307 256.663
R458 B.n482 B.n308 256.663
R459 B.n482 B.n309 256.663
R460 B.n482 B.n310 256.663
R461 B.n482 B.n311 256.663
R462 B.n482 B.n312 256.663
R463 B.n482 B.n313 256.663
R464 B.n482 B.n314 256.663
R465 B.n482 B.n315 256.663
R466 B.n482 B.n316 256.663
R467 B.n482 B.n317 256.663
R468 B.n482 B.n318 256.663
R469 B.n482 B.n319 256.663
R470 B.n482 B.n320 256.663
R471 B.n482 B.n321 256.663
R472 B.n482 B.n322 256.663
R473 B.n482 B.n323 256.663
R474 B.n482 B.n324 256.663
R475 B.n482 B.n325 256.663
R476 B.n482 B.n326 256.663
R477 B.n482 B.n327 256.663
R478 B.n482 B.n328 256.663
R479 B.n482 B.n329 256.663
R480 B.n482 B.n330 256.663
R481 B.n482 B.n331 256.663
R482 B.n482 B.n332 256.663
R483 B.n482 B.n333 256.663
R484 B.n482 B.n334 256.663
R485 B.n482 B.n335 256.663
R486 B.n482 B.n336 256.663
R487 B.n482 B.n337 256.663
R488 B.n482 B.n338 256.663
R489 B.n702 B.n701 256.663
R490 B.n109 B.n108 163.367
R491 B.n113 B.n112 163.367
R492 B.n117 B.n116 163.367
R493 B.n121 B.n120 163.367
R494 B.n125 B.n124 163.367
R495 B.n129 B.n128 163.367
R496 B.n133 B.n132 163.367
R497 B.n137 B.n136 163.367
R498 B.n141 B.n140 163.367
R499 B.n145 B.n144 163.367
R500 B.n149 B.n148 163.367
R501 B.n153 B.n152 163.367
R502 B.n157 B.n156 163.367
R503 B.n161 B.n160 163.367
R504 B.n165 B.n164 163.367
R505 B.n169 B.n168 163.367
R506 B.n173 B.n172 163.367
R507 B.n177 B.n176 163.367
R508 B.n181 B.n180 163.367
R509 B.n185 B.n184 163.367
R510 B.n189 B.n188 163.367
R511 B.n193 B.n192 163.367
R512 B.n197 B.n196 163.367
R513 B.n201 B.n200 163.367
R514 B.n205 B.n204 163.367
R515 B.n209 B.n208 163.367
R516 B.n213 B.n212 163.367
R517 B.n217 B.n216 163.367
R518 B.n221 B.n220 163.367
R519 B.n225 B.n224 163.367
R520 B.n229 B.n228 163.367
R521 B.n233 B.n232 163.367
R522 B.n237 B.n236 163.367
R523 B.n239 B.n98 163.367
R524 B.n487 B.n303 163.367
R525 B.n487 B.n297 163.367
R526 B.n495 B.n297 163.367
R527 B.n495 B.n295 163.367
R528 B.n499 B.n295 163.367
R529 B.n499 B.n290 163.367
R530 B.n508 B.n290 163.367
R531 B.n508 B.n288 163.367
R532 B.n512 B.n288 163.367
R533 B.n512 B.n282 163.367
R534 B.n520 B.n282 163.367
R535 B.n520 B.n280 163.367
R536 B.n524 B.n280 163.367
R537 B.n524 B.n273 163.367
R538 B.n532 B.n273 163.367
R539 B.n532 B.n271 163.367
R540 B.n536 B.n271 163.367
R541 B.n536 B.n266 163.367
R542 B.n544 B.n266 163.367
R543 B.n544 B.n264 163.367
R544 B.n548 B.n264 163.367
R545 B.n548 B.n259 163.367
R546 B.n557 B.n259 163.367
R547 B.n557 B.n257 163.367
R548 B.n561 B.n257 163.367
R549 B.n561 B.n250 163.367
R550 B.n569 B.n250 163.367
R551 B.n569 B.n248 163.367
R552 B.n574 B.n248 163.367
R553 B.n574 B.n243 163.367
R554 B.n582 B.n243 163.367
R555 B.n583 B.n582 163.367
R556 B.n583 B.n5 163.367
R557 B.n6 B.n5 163.367
R558 B.n7 B.n6 163.367
R559 B.n589 B.n7 163.367
R560 B.n590 B.n589 163.367
R561 B.n590 B.n13 163.367
R562 B.n14 B.n13 163.367
R563 B.n15 B.n14 163.367
R564 B.n595 B.n15 163.367
R565 B.n595 B.n20 163.367
R566 B.n21 B.n20 163.367
R567 B.n22 B.n21 163.367
R568 B.n600 B.n22 163.367
R569 B.n600 B.n27 163.367
R570 B.n28 B.n27 163.367
R571 B.n29 B.n28 163.367
R572 B.n605 B.n29 163.367
R573 B.n605 B.n34 163.367
R574 B.n35 B.n34 163.367
R575 B.n36 B.n35 163.367
R576 B.n610 B.n36 163.367
R577 B.n610 B.n41 163.367
R578 B.n42 B.n41 163.367
R579 B.n43 B.n42 163.367
R580 B.n615 B.n43 163.367
R581 B.n615 B.n48 163.367
R582 B.n49 B.n48 163.367
R583 B.n50 B.n49 163.367
R584 B.n620 B.n50 163.367
R585 B.n620 B.n55 163.367
R586 B.n56 B.n55 163.367
R587 B.n57 B.n56 163.367
R588 B.n625 B.n57 163.367
R589 B.n625 B.n62 163.367
R590 B.n63 B.n62 163.367
R591 B.n340 B.n339 163.367
R592 B.n475 B.n339 163.367
R593 B.n473 B.n472 163.367
R594 B.n469 B.n468 163.367
R595 B.n465 B.n464 163.367
R596 B.n461 B.n460 163.367
R597 B.n457 B.n456 163.367
R598 B.n453 B.n452 163.367
R599 B.n449 B.n448 163.367
R600 B.n445 B.n444 163.367
R601 B.n441 B.n440 163.367
R602 B.n437 B.n436 163.367
R603 B.n433 B.n432 163.367
R604 B.n429 B.n428 163.367
R605 B.n425 B.n424 163.367
R606 B.n420 B.n419 163.367
R607 B.n416 B.n415 163.367
R608 B.n412 B.n411 163.367
R609 B.n408 B.n407 163.367
R610 B.n404 B.n403 163.367
R611 B.n399 B.n398 163.367
R612 B.n395 B.n394 163.367
R613 B.n391 B.n390 163.367
R614 B.n387 B.n386 163.367
R615 B.n383 B.n382 163.367
R616 B.n379 B.n378 163.367
R617 B.n375 B.n374 163.367
R618 B.n371 B.n370 163.367
R619 B.n367 B.n366 163.367
R620 B.n363 B.n362 163.367
R621 B.n359 B.n358 163.367
R622 B.n355 B.n354 163.367
R623 B.n351 B.n350 163.367
R624 B.n347 B.n346 163.367
R625 B.n483 B.n305 163.367
R626 B.n489 B.n301 163.367
R627 B.n489 B.n299 163.367
R628 B.n493 B.n299 163.367
R629 B.n493 B.n293 163.367
R630 B.n502 B.n293 163.367
R631 B.n502 B.n291 163.367
R632 B.n506 B.n291 163.367
R633 B.n506 B.n286 163.367
R634 B.n514 B.n286 163.367
R635 B.n514 B.n284 163.367
R636 B.n518 B.n284 163.367
R637 B.n518 B.n278 163.367
R638 B.n526 B.n278 163.367
R639 B.n526 B.n276 163.367
R640 B.n530 B.n276 163.367
R641 B.n530 B.n270 163.367
R642 B.n538 B.n270 163.367
R643 B.n538 B.n268 163.367
R644 B.n542 B.n268 163.367
R645 B.n542 B.n262 163.367
R646 B.n551 B.n262 163.367
R647 B.n551 B.n260 163.367
R648 B.n555 B.n260 163.367
R649 B.n555 B.n255 163.367
R650 B.n563 B.n255 163.367
R651 B.n563 B.n253 163.367
R652 B.n567 B.n253 163.367
R653 B.n567 B.n247 163.367
R654 B.n576 B.n247 163.367
R655 B.n576 B.n245 163.367
R656 B.n580 B.n245 163.367
R657 B.n580 B.n3 163.367
R658 B.n700 B.n3 163.367
R659 B.n696 B.n2 163.367
R660 B.n696 B.n695 163.367
R661 B.n695 B.n9 163.367
R662 B.n691 B.n9 163.367
R663 B.n691 B.n11 163.367
R664 B.n687 B.n11 163.367
R665 B.n687 B.n17 163.367
R666 B.n683 B.n17 163.367
R667 B.n683 B.n19 163.367
R668 B.n679 B.n19 163.367
R669 B.n679 B.n23 163.367
R670 B.n675 B.n23 163.367
R671 B.n675 B.n25 163.367
R672 B.n671 B.n25 163.367
R673 B.n671 B.n31 163.367
R674 B.n667 B.n31 163.367
R675 B.n667 B.n33 163.367
R676 B.n663 B.n33 163.367
R677 B.n663 B.n38 163.367
R678 B.n659 B.n38 163.367
R679 B.n659 B.n40 163.367
R680 B.n655 B.n40 163.367
R681 B.n655 B.n45 163.367
R682 B.n651 B.n45 163.367
R683 B.n651 B.n47 163.367
R684 B.n647 B.n47 163.367
R685 B.n647 B.n51 163.367
R686 B.n643 B.n51 163.367
R687 B.n643 B.n53 163.367
R688 B.n639 B.n53 163.367
R689 B.n639 B.n59 163.367
R690 B.n635 B.n59 163.367
R691 B.n635 B.n61 163.367
R692 B.n99 B.t15 110.835
R693 B.n343 B.t12 110.835
R694 B.n102 B.t18 110.825
R695 B.n341 B.t9 110.825
R696 B.n482 B.n302 102.192
R697 B.n633 B.n632 102.192
R698 B.n105 B.n64 71.676
R699 B.n109 B.n65 71.676
R700 B.n113 B.n66 71.676
R701 B.n117 B.n67 71.676
R702 B.n121 B.n68 71.676
R703 B.n125 B.n69 71.676
R704 B.n129 B.n70 71.676
R705 B.n133 B.n71 71.676
R706 B.n137 B.n72 71.676
R707 B.n141 B.n73 71.676
R708 B.n145 B.n74 71.676
R709 B.n149 B.n75 71.676
R710 B.n153 B.n76 71.676
R711 B.n157 B.n77 71.676
R712 B.n161 B.n78 71.676
R713 B.n165 B.n79 71.676
R714 B.n169 B.n80 71.676
R715 B.n173 B.n81 71.676
R716 B.n177 B.n82 71.676
R717 B.n181 B.n83 71.676
R718 B.n185 B.n84 71.676
R719 B.n189 B.n85 71.676
R720 B.n193 B.n86 71.676
R721 B.n197 B.n87 71.676
R722 B.n201 B.n88 71.676
R723 B.n205 B.n89 71.676
R724 B.n209 B.n90 71.676
R725 B.n213 B.n91 71.676
R726 B.n217 B.n92 71.676
R727 B.n221 B.n93 71.676
R728 B.n225 B.n94 71.676
R729 B.n229 B.n95 71.676
R730 B.n233 B.n96 71.676
R731 B.n237 B.n97 71.676
R732 B.n631 B.n98 71.676
R733 B.n631 B.n630 71.676
R734 B.n239 B.n97 71.676
R735 B.n236 B.n96 71.676
R736 B.n232 B.n95 71.676
R737 B.n228 B.n94 71.676
R738 B.n224 B.n93 71.676
R739 B.n220 B.n92 71.676
R740 B.n216 B.n91 71.676
R741 B.n212 B.n90 71.676
R742 B.n208 B.n89 71.676
R743 B.n204 B.n88 71.676
R744 B.n200 B.n87 71.676
R745 B.n196 B.n86 71.676
R746 B.n192 B.n85 71.676
R747 B.n188 B.n84 71.676
R748 B.n184 B.n83 71.676
R749 B.n180 B.n82 71.676
R750 B.n176 B.n81 71.676
R751 B.n172 B.n80 71.676
R752 B.n168 B.n79 71.676
R753 B.n164 B.n78 71.676
R754 B.n160 B.n77 71.676
R755 B.n156 B.n76 71.676
R756 B.n152 B.n75 71.676
R757 B.n148 B.n74 71.676
R758 B.n144 B.n73 71.676
R759 B.n140 B.n72 71.676
R760 B.n136 B.n71 71.676
R761 B.n132 B.n70 71.676
R762 B.n128 B.n69 71.676
R763 B.n124 B.n68 71.676
R764 B.n120 B.n67 71.676
R765 B.n116 B.n66 71.676
R766 B.n112 B.n65 71.676
R767 B.n108 B.n64 71.676
R768 B.n481 B.n480 71.676
R769 B.n475 B.n306 71.676
R770 B.n472 B.n307 71.676
R771 B.n468 B.n308 71.676
R772 B.n464 B.n309 71.676
R773 B.n460 B.n310 71.676
R774 B.n456 B.n311 71.676
R775 B.n452 B.n312 71.676
R776 B.n448 B.n313 71.676
R777 B.n444 B.n314 71.676
R778 B.n440 B.n315 71.676
R779 B.n436 B.n316 71.676
R780 B.n432 B.n317 71.676
R781 B.n428 B.n318 71.676
R782 B.n424 B.n319 71.676
R783 B.n419 B.n320 71.676
R784 B.n415 B.n321 71.676
R785 B.n411 B.n322 71.676
R786 B.n407 B.n323 71.676
R787 B.n403 B.n324 71.676
R788 B.n398 B.n325 71.676
R789 B.n394 B.n326 71.676
R790 B.n390 B.n327 71.676
R791 B.n386 B.n328 71.676
R792 B.n382 B.n329 71.676
R793 B.n378 B.n330 71.676
R794 B.n374 B.n331 71.676
R795 B.n370 B.n332 71.676
R796 B.n366 B.n333 71.676
R797 B.n362 B.n334 71.676
R798 B.n358 B.n335 71.676
R799 B.n354 B.n336 71.676
R800 B.n350 B.n337 71.676
R801 B.n346 B.n338 71.676
R802 B.n481 B.n340 71.676
R803 B.n473 B.n306 71.676
R804 B.n469 B.n307 71.676
R805 B.n465 B.n308 71.676
R806 B.n461 B.n309 71.676
R807 B.n457 B.n310 71.676
R808 B.n453 B.n311 71.676
R809 B.n449 B.n312 71.676
R810 B.n445 B.n313 71.676
R811 B.n441 B.n314 71.676
R812 B.n437 B.n315 71.676
R813 B.n433 B.n316 71.676
R814 B.n429 B.n317 71.676
R815 B.n425 B.n318 71.676
R816 B.n420 B.n319 71.676
R817 B.n416 B.n320 71.676
R818 B.n412 B.n321 71.676
R819 B.n408 B.n322 71.676
R820 B.n404 B.n323 71.676
R821 B.n399 B.n324 71.676
R822 B.n395 B.n325 71.676
R823 B.n391 B.n326 71.676
R824 B.n387 B.n327 71.676
R825 B.n383 B.n328 71.676
R826 B.n379 B.n329 71.676
R827 B.n375 B.n330 71.676
R828 B.n371 B.n331 71.676
R829 B.n367 B.n332 71.676
R830 B.n363 B.n333 71.676
R831 B.n359 B.n334 71.676
R832 B.n355 B.n335 71.676
R833 B.n351 B.n336 71.676
R834 B.n347 B.n337 71.676
R835 B.n338 B.n305 71.676
R836 B.n701 B.n700 71.676
R837 B.n701 B.n2 71.676
R838 B.n100 B.t16 68.9433
R839 B.n344 B.t11 68.9433
R840 B.n103 B.t19 68.9336
R841 B.n342 B.t8 68.9336
R842 B.n104 B.n103 59.5399
R843 B.n101 B.n100 59.5399
R844 B.n401 B.n344 59.5399
R845 B.n422 B.n342 59.5399
R846 B.n488 B.n302 55.5932
R847 B.n488 B.n298 55.5932
R848 B.n494 B.n298 55.5932
R849 B.n494 B.n294 55.5932
R850 B.n501 B.n294 55.5932
R851 B.n501 B.n500 55.5932
R852 B.n507 B.n287 55.5932
R853 B.n513 B.n287 55.5932
R854 B.n513 B.n283 55.5932
R855 B.n519 B.n283 55.5932
R856 B.n519 B.n279 55.5932
R857 B.n525 B.n279 55.5932
R858 B.n525 B.n274 55.5932
R859 B.n531 B.n274 55.5932
R860 B.n531 B.n275 55.5932
R861 B.n537 B.n267 55.5932
R862 B.n543 B.n267 55.5932
R863 B.n543 B.n263 55.5932
R864 B.n550 B.n263 55.5932
R865 B.n550 B.n549 55.5932
R866 B.n556 B.n256 55.5932
R867 B.n562 B.n256 55.5932
R868 B.n562 B.n251 55.5932
R869 B.n568 B.n251 55.5932
R870 B.n568 B.n252 55.5932
R871 B.n575 B.n244 55.5932
R872 B.n581 B.n244 55.5932
R873 B.n581 B.n4 55.5932
R874 B.n699 B.n4 55.5932
R875 B.n699 B.n698 55.5932
R876 B.n698 B.n697 55.5932
R877 B.n697 B.n8 55.5932
R878 B.n12 B.n8 55.5932
R879 B.n690 B.n12 55.5932
R880 B.n689 B.n688 55.5932
R881 B.n688 B.n16 55.5932
R882 B.n682 B.n16 55.5932
R883 B.n682 B.n681 55.5932
R884 B.n681 B.n680 55.5932
R885 B.n674 B.n26 55.5932
R886 B.n674 B.n673 55.5932
R887 B.n673 B.n672 55.5932
R888 B.n672 B.n30 55.5932
R889 B.n666 B.n30 55.5932
R890 B.n665 B.n664 55.5932
R891 B.n664 B.n37 55.5932
R892 B.n658 B.n37 55.5932
R893 B.n658 B.n657 55.5932
R894 B.n657 B.n656 55.5932
R895 B.n656 B.n44 55.5932
R896 B.n650 B.n44 55.5932
R897 B.n650 B.n649 55.5932
R898 B.n649 B.n648 55.5932
R899 B.n642 B.n54 55.5932
R900 B.n642 B.n641 55.5932
R901 B.n641 B.n640 55.5932
R902 B.n640 B.n58 55.5932
R903 B.n634 B.n58 55.5932
R904 B.n634 B.n633 55.5932
R905 B.n537 B.t0 54.7757
R906 B.n666 B.t3 54.7757
R907 B.n103 B.n102 41.8914
R908 B.n100 B.n99 41.8914
R909 B.n344 B.n343 41.8914
R910 B.n342 B.n341 41.8914
R911 B.n252 B.t1 40.06
R912 B.t5 B.n689 40.06
R913 B.n556 B.t4 35.1547
R914 B.n680 B.t2 35.1547
R915 B.n479 B.n300 34.4981
R916 B.n485 B.n484 34.4981
R917 B.n629 B.n628 34.4981
R918 B.n106 B.n60 34.4981
R919 B.n507 B.t7 30.2495
R920 B.n648 B.t14 30.2495
R921 B.n500 B.t7 25.3442
R922 B.n54 B.t14 25.3442
R923 B.n549 B.t4 20.439
R924 B.n26 B.t2 20.439
R925 B B.n702 18.0485
R926 B.n575 B.t1 15.5338
R927 B.n690 B.t5 15.5338
R928 B.n490 B.n300 10.6151
R929 B.n491 B.n490 10.6151
R930 B.n492 B.n491 10.6151
R931 B.n492 B.n292 10.6151
R932 B.n503 B.n292 10.6151
R933 B.n504 B.n503 10.6151
R934 B.n505 B.n504 10.6151
R935 B.n505 B.n285 10.6151
R936 B.n515 B.n285 10.6151
R937 B.n516 B.n515 10.6151
R938 B.n517 B.n516 10.6151
R939 B.n517 B.n277 10.6151
R940 B.n527 B.n277 10.6151
R941 B.n528 B.n527 10.6151
R942 B.n529 B.n528 10.6151
R943 B.n529 B.n269 10.6151
R944 B.n539 B.n269 10.6151
R945 B.n540 B.n539 10.6151
R946 B.n541 B.n540 10.6151
R947 B.n541 B.n261 10.6151
R948 B.n552 B.n261 10.6151
R949 B.n553 B.n552 10.6151
R950 B.n554 B.n553 10.6151
R951 B.n554 B.n254 10.6151
R952 B.n564 B.n254 10.6151
R953 B.n565 B.n564 10.6151
R954 B.n566 B.n565 10.6151
R955 B.n566 B.n246 10.6151
R956 B.n577 B.n246 10.6151
R957 B.n578 B.n577 10.6151
R958 B.n579 B.n578 10.6151
R959 B.n579 B.n0 10.6151
R960 B.n479 B.n478 10.6151
R961 B.n478 B.n477 10.6151
R962 B.n477 B.n476 10.6151
R963 B.n476 B.n474 10.6151
R964 B.n474 B.n471 10.6151
R965 B.n471 B.n470 10.6151
R966 B.n470 B.n467 10.6151
R967 B.n467 B.n466 10.6151
R968 B.n466 B.n463 10.6151
R969 B.n463 B.n462 10.6151
R970 B.n462 B.n459 10.6151
R971 B.n459 B.n458 10.6151
R972 B.n458 B.n455 10.6151
R973 B.n455 B.n454 10.6151
R974 B.n454 B.n451 10.6151
R975 B.n451 B.n450 10.6151
R976 B.n450 B.n447 10.6151
R977 B.n447 B.n446 10.6151
R978 B.n446 B.n443 10.6151
R979 B.n443 B.n442 10.6151
R980 B.n442 B.n439 10.6151
R981 B.n439 B.n438 10.6151
R982 B.n438 B.n435 10.6151
R983 B.n435 B.n434 10.6151
R984 B.n434 B.n431 10.6151
R985 B.n431 B.n430 10.6151
R986 B.n430 B.n427 10.6151
R987 B.n427 B.n426 10.6151
R988 B.n426 B.n423 10.6151
R989 B.n421 B.n418 10.6151
R990 B.n418 B.n417 10.6151
R991 B.n417 B.n414 10.6151
R992 B.n414 B.n413 10.6151
R993 B.n413 B.n410 10.6151
R994 B.n410 B.n409 10.6151
R995 B.n409 B.n406 10.6151
R996 B.n406 B.n405 10.6151
R997 B.n405 B.n402 10.6151
R998 B.n400 B.n397 10.6151
R999 B.n397 B.n396 10.6151
R1000 B.n396 B.n393 10.6151
R1001 B.n393 B.n392 10.6151
R1002 B.n392 B.n389 10.6151
R1003 B.n389 B.n388 10.6151
R1004 B.n388 B.n385 10.6151
R1005 B.n385 B.n384 10.6151
R1006 B.n384 B.n381 10.6151
R1007 B.n381 B.n380 10.6151
R1008 B.n380 B.n377 10.6151
R1009 B.n377 B.n376 10.6151
R1010 B.n376 B.n373 10.6151
R1011 B.n373 B.n372 10.6151
R1012 B.n372 B.n369 10.6151
R1013 B.n369 B.n368 10.6151
R1014 B.n368 B.n365 10.6151
R1015 B.n365 B.n364 10.6151
R1016 B.n364 B.n361 10.6151
R1017 B.n361 B.n360 10.6151
R1018 B.n360 B.n357 10.6151
R1019 B.n357 B.n356 10.6151
R1020 B.n356 B.n353 10.6151
R1021 B.n353 B.n352 10.6151
R1022 B.n352 B.n349 10.6151
R1023 B.n349 B.n348 10.6151
R1024 B.n348 B.n345 10.6151
R1025 B.n345 B.n304 10.6151
R1026 B.n484 B.n304 10.6151
R1027 B.n486 B.n485 10.6151
R1028 B.n486 B.n296 10.6151
R1029 B.n496 B.n296 10.6151
R1030 B.n497 B.n496 10.6151
R1031 B.n498 B.n497 10.6151
R1032 B.n498 B.n289 10.6151
R1033 B.n509 B.n289 10.6151
R1034 B.n510 B.n509 10.6151
R1035 B.n511 B.n510 10.6151
R1036 B.n511 B.n281 10.6151
R1037 B.n521 B.n281 10.6151
R1038 B.n522 B.n521 10.6151
R1039 B.n523 B.n522 10.6151
R1040 B.n523 B.n272 10.6151
R1041 B.n533 B.n272 10.6151
R1042 B.n534 B.n533 10.6151
R1043 B.n535 B.n534 10.6151
R1044 B.n535 B.n265 10.6151
R1045 B.n545 B.n265 10.6151
R1046 B.n546 B.n545 10.6151
R1047 B.n547 B.n546 10.6151
R1048 B.n547 B.n258 10.6151
R1049 B.n558 B.n258 10.6151
R1050 B.n559 B.n558 10.6151
R1051 B.n560 B.n559 10.6151
R1052 B.n560 B.n249 10.6151
R1053 B.n570 B.n249 10.6151
R1054 B.n571 B.n570 10.6151
R1055 B.n573 B.n571 10.6151
R1056 B.n573 B.n572 10.6151
R1057 B.n572 B.n242 10.6151
R1058 B.n584 B.n242 10.6151
R1059 B.n585 B.n584 10.6151
R1060 B.n586 B.n585 10.6151
R1061 B.n587 B.n586 10.6151
R1062 B.n588 B.n587 10.6151
R1063 B.n591 B.n588 10.6151
R1064 B.n592 B.n591 10.6151
R1065 B.n593 B.n592 10.6151
R1066 B.n594 B.n593 10.6151
R1067 B.n596 B.n594 10.6151
R1068 B.n597 B.n596 10.6151
R1069 B.n598 B.n597 10.6151
R1070 B.n599 B.n598 10.6151
R1071 B.n601 B.n599 10.6151
R1072 B.n602 B.n601 10.6151
R1073 B.n603 B.n602 10.6151
R1074 B.n604 B.n603 10.6151
R1075 B.n606 B.n604 10.6151
R1076 B.n607 B.n606 10.6151
R1077 B.n608 B.n607 10.6151
R1078 B.n609 B.n608 10.6151
R1079 B.n611 B.n609 10.6151
R1080 B.n612 B.n611 10.6151
R1081 B.n613 B.n612 10.6151
R1082 B.n614 B.n613 10.6151
R1083 B.n616 B.n614 10.6151
R1084 B.n617 B.n616 10.6151
R1085 B.n618 B.n617 10.6151
R1086 B.n619 B.n618 10.6151
R1087 B.n621 B.n619 10.6151
R1088 B.n622 B.n621 10.6151
R1089 B.n623 B.n622 10.6151
R1090 B.n624 B.n623 10.6151
R1091 B.n626 B.n624 10.6151
R1092 B.n627 B.n626 10.6151
R1093 B.n628 B.n627 10.6151
R1094 B.n694 B.n1 10.6151
R1095 B.n694 B.n693 10.6151
R1096 B.n693 B.n692 10.6151
R1097 B.n692 B.n10 10.6151
R1098 B.n686 B.n10 10.6151
R1099 B.n686 B.n685 10.6151
R1100 B.n685 B.n684 10.6151
R1101 B.n684 B.n18 10.6151
R1102 B.n678 B.n18 10.6151
R1103 B.n678 B.n677 10.6151
R1104 B.n677 B.n676 10.6151
R1105 B.n676 B.n24 10.6151
R1106 B.n670 B.n24 10.6151
R1107 B.n670 B.n669 10.6151
R1108 B.n669 B.n668 10.6151
R1109 B.n668 B.n32 10.6151
R1110 B.n662 B.n32 10.6151
R1111 B.n662 B.n661 10.6151
R1112 B.n661 B.n660 10.6151
R1113 B.n660 B.n39 10.6151
R1114 B.n654 B.n39 10.6151
R1115 B.n654 B.n653 10.6151
R1116 B.n653 B.n652 10.6151
R1117 B.n652 B.n46 10.6151
R1118 B.n646 B.n46 10.6151
R1119 B.n646 B.n645 10.6151
R1120 B.n645 B.n644 10.6151
R1121 B.n644 B.n52 10.6151
R1122 B.n638 B.n52 10.6151
R1123 B.n638 B.n637 10.6151
R1124 B.n637 B.n636 10.6151
R1125 B.n636 B.n60 10.6151
R1126 B.n107 B.n106 10.6151
R1127 B.n110 B.n107 10.6151
R1128 B.n111 B.n110 10.6151
R1129 B.n114 B.n111 10.6151
R1130 B.n115 B.n114 10.6151
R1131 B.n118 B.n115 10.6151
R1132 B.n119 B.n118 10.6151
R1133 B.n122 B.n119 10.6151
R1134 B.n123 B.n122 10.6151
R1135 B.n126 B.n123 10.6151
R1136 B.n127 B.n126 10.6151
R1137 B.n130 B.n127 10.6151
R1138 B.n131 B.n130 10.6151
R1139 B.n134 B.n131 10.6151
R1140 B.n135 B.n134 10.6151
R1141 B.n138 B.n135 10.6151
R1142 B.n139 B.n138 10.6151
R1143 B.n142 B.n139 10.6151
R1144 B.n143 B.n142 10.6151
R1145 B.n146 B.n143 10.6151
R1146 B.n147 B.n146 10.6151
R1147 B.n150 B.n147 10.6151
R1148 B.n151 B.n150 10.6151
R1149 B.n154 B.n151 10.6151
R1150 B.n155 B.n154 10.6151
R1151 B.n158 B.n155 10.6151
R1152 B.n159 B.n158 10.6151
R1153 B.n162 B.n159 10.6151
R1154 B.n163 B.n162 10.6151
R1155 B.n167 B.n166 10.6151
R1156 B.n170 B.n167 10.6151
R1157 B.n171 B.n170 10.6151
R1158 B.n174 B.n171 10.6151
R1159 B.n175 B.n174 10.6151
R1160 B.n178 B.n175 10.6151
R1161 B.n179 B.n178 10.6151
R1162 B.n182 B.n179 10.6151
R1163 B.n183 B.n182 10.6151
R1164 B.n187 B.n186 10.6151
R1165 B.n190 B.n187 10.6151
R1166 B.n191 B.n190 10.6151
R1167 B.n194 B.n191 10.6151
R1168 B.n195 B.n194 10.6151
R1169 B.n198 B.n195 10.6151
R1170 B.n199 B.n198 10.6151
R1171 B.n202 B.n199 10.6151
R1172 B.n203 B.n202 10.6151
R1173 B.n206 B.n203 10.6151
R1174 B.n207 B.n206 10.6151
R1175 B.n210 B.n207 10.6151
R1176 B.n211 B.n210 10.6151
R1177 B.n214 B.n211 10.6151
R1178 B.n215 B.n214 10.6151
R1179 B.n218 B.n215 10.6151
R1180 B.n219 B.n218 10.6151
R1181 B.n222 B.n219 10.6151
R1182 B.n223 B.n222 10.6151
R1183 B.n226 B.n223 10.6151
R1184 B.n227 B.n226 10.6151
R1185 B.n230 B.n227 10.6151
R1186 B.n231 B.n230 10.6151
R1187 B.n234 B.n231 10.6151
R1188 B.n235 B.n234 10.6151
R1189 B.n238 B.n235 10.6151
R1190 B.n240 B.n238 10.6151
R1191 B.n241 B.n240 10.6151
R1192 B.n629 B.n241 10.6151
R1193 B.n423 B.n422 9.36635
R1194 B.n401 B.n400 9.36635
R1195 B.n163 B.n104 9.36635
R1196 B.n186 B.n101 9.36635
R1197 B.n702 B.n0 8.11757
R1198 B.n702 B.n1 8.11757
R1199 B.n422 B.n421 1.24928
R1200 B.n402 B.n401 1.24928
R1201 B.n166 B.n104 1.24928
R1202 B.n183 B.n101 1.24928
R1203 B.n275 B.t0 0.81804
R1204 B.t3 B.n665 0.81804
R1205 VN.n21 VN.n12 161.3
R1206 VN.n20 VN.n19 161.3
R1207 VN.n18 VN.n13 161.3
R1208 VN.n17 VN.n16 161.3
R1209 VN.n9 VN.n0 161.3
R1210 VN.n8 VN.n7 161.3
R1211 VN.n6 VN.n1 161.3
R1212 VN.n5 VN.n4 161.3
R1213 VN.n2 VN.t1 138.171
R1214 VN.n14 VN.t2 138.171
R1215 VN.n3 VN.t4 107.727
R1216 VN.n10 VN.t5 107.727
R1217 VN.n15 VN.t0 107.727
R1218 VN.n22 VN.t3 107.727
R1219 VN.n11 VN.n10 90.7429
R1220 VN.n23 VN.n22 90.7429
R1221 VN.n3 VN.n2 57.7341
R1222 VN.n15 VN.n14 57.7341
R1223 VN.n8 VN.n1 56.5617
R1224 VN.n20 VN.n13 56.5617
R1225 VN VN.n23 43.0285
R1226 VN.n4 VN.n1 24.5923
R1227 VN.n9 VN.n8 24.5923
R1228 VN.n16 VN.n13 24.5923
R1229 VN.n21 VN.n20 24.5923
R1230 VN.n10 VN.n9 20.1658
R1231 VN.n22 VN.n21 20.1658
R1232 VN.n17 VN.n14 13.2724
R1233 VN.n5 VN.n2 13.2724
R1234 VN.n4 VN.n3 12.2964
R1235 VN.n16 VN.n15 12.2964
R1236 VN.n23 VN.n12 0.278335
R1237 VN.n11 VN.n0 0.278335
R1238 VN.n19 VN.n12 0.189894
R1239 VN.n19 VN.n18 0.189894
R1240 VN.n18 VN.n17 0.189894
R1241 VN.n6 VN.n5 0.189894
R1242 VN.n7 VN.n6 0.189894
R1243 VN.n7 VN.n0 0.189894
R1244 VN VN.n11 0.153485
R1245 VDD2.n1 VDD2.t5 67.8452
R1246 VDD2.n2 VDD2.t3 66.5041
R1247 VDD2.n1 VDD2.n0 64.4935
R1248 VDD2 VDD2.n3 64.4908
R1249 VDD2.n2 VDD2.n1 36.8187
R1250 VDD2.n3 VDD2.t0 2.42104
R1251 VDD2.n3 VDD2.t4 2.42104
R1252 VDD2.n0 VDD2.t2 2.42104
R1253 VDD2.n0 VDD2.t1 2.42104
R1254 VDD2 VDD2.n2 1.45524
R1255 VTAIL.n7 VTAIL.t9 49.8253
R1256 VTAIL.n10 VTAIL.t5 49.8252
R1257 VTAIL.n11 VTAIL.t6 49.8252
R1258 VTAIL.n2 VTAIL.t1 49.8252
R1259 VTAIL.n9 VTAIL.n8 47.4048
R1260 VTAIL.n6 VTAIL.n5 47.4048
R1261 VTAIL.n1 VTAIL.n0 47.4046
R1262 VTAIL.n4 VTAIL.n3 47.4046
R1263 VTAIL.n6 VTAIL.n4 23.1427
R1264 VTAIL.n11 VTAIL.n10 21.2807
R1265 VTAIL.n0 VTAIL.t10 2.42104
R1266 VTAIL.n0 VTAIL.t7 2.42104
R1267 VTAIL.n3 VTAIL.t0 2.42104
R1268 VTAIL.n3 VTAIL.t3 2.42104
R1269 VTAIL.n8 VTAIL.t4 2.42104
R1270 VTAIL.n8 VTAIL.t2 2.42104
R1271 VTAIL.n5 VTAIL.t8 2.42104
R1272 VTAIL.n5 VTAIL.t11 2.42104
R1273 VTAIL.n7 VTAIL.n6 1.86257
R1274 VTAIL.n10 VTAIL.n9 1.86257
R1275 VTAIL.n4 VTAIL.n2 1.86257
R1276 VTAIL.n9 VTAIL.n7 1.40136
R1277 VTAIL.n2 VTAIL.n1 1.40136
R1278 VTAIL VTAIL.n11 1.33886
R1279 VTAIL VTAIL.n1 0.524207
R1280 VP.n9 VP.n8 161.3
R1281 VP.n10 VP.n5 161.3
R1282 VP.n12 VP.n11 161.3
R1283 VP.n13 VP.n4 161.3
R1284 VP.n30 VP.n0 161.3
R1285 VP.n29 VP.n28 161.3
R1286 VP.n27 VP.n1 161.3
R1287 VP.n26 VP.n25 161.3
R1288 VP.n23 VP.n2 161.3
R1289 VP.n22 VP.n21 161.3
R1290 VP.n20 VP.n3 161.3
R1291 VP.n19 VP.n18 161.3
R1292 VP.n6 VP.t2 138.171
R1293 VP.n17 VP.t1 107.727
R1294 VP.n24 VP.t5 107.727
R1295 VP.n31 VP.t3 107.727
R1296 VP.n14 VP.t0 107.727
R1297 VP.n7 VP.t4 107.727
R1298 VP.n17 VP.n16 90.7429
R1299 VP.n32 VP.n31 90.7429
R1300 VP.n15 VP.n14 90.7429
R1301 VP.n7 VP.n6 57.7341
R1302 VP.n22 VP.n3 56.5617
R1303 VP.n29 VP.n1 56.5617
R1304 VP.n12 VP.n5 56.5617
R1305 VP.n16 VP.n15 42.7497
R1306 VP.n18 VP.n3 24.5923
R1307 VP.n23 VP.n22 24.5923
R1308 VP.n25 VP.n1 24.5923
R1309 VP.n30 VP.n29 24.5923
R1310 VP.n13 VP.n12 24.5923
R1311 VP.n8 VP.n5 24.5923
R1312 VP.n18 VP.n17 20.1658
R1313 VP.n31 VP.n30 20.1658
R1314 VP.n14 VP.n13 20.1658
R1315 VP.n9 VP.n6 13.2724
R1316 VP.n24 VP.n23 12.2964
R1317 VP.n25 VP.n24 12.2964
R1318 VP.n8 VP.n7 12.2964
R1319 VP.n15 VP.n4 0.278335
R1320 VP.n19 VP.n16 0.278335
R1321 VP.n32 VP.n0 0.278335
R1322 VP.n10 VP.n9 0.189894
R1323 VP.n11 VP.n10 0.189894
R1324 VP.n11 VP.n4 0.189894
R1325 VP.n20 VP.n19 0.189894
R1326 VP.n21 VP.n20 0.189894
R1327 VP.n21 VP.n2 0.189894
R1328 VP.n26 VP.n2 0.189894
R1329 VP.n27 VP.n26 0.189894
R1330 VP.n28 VP.n27 0.189894
R1331 VP.n28 VP.n0 0.189894
R1332 VP VP.n32 0.153485
R1333 VDD1 VDD1.t3 67.9588
R1334 VDD1.n1 VDD1.t4 67.8452
R1335 VDD1.n1 VDD1.n0 64.4935
R1336 VDD1.n3 VDD1.n2 64.0834
R1337 VDD1.n3 VDD1.n1 38.3328
R1338 VDD1.n2 VDD1.t1 2.42104
R1339 VDD1.n2 VDD1.t5 2.42104
R1340 VDD1.n0 VDD1.t0 2.42104
R1341 VDD1.n0 VDD1.t2 2.42104
R1342 VDD1 VDD1.n3 0.407828
C0 VP VN 5.47113f
C1 VTAIL VDD1 6.18441f
C2 VTAIL VDD2 6.23024f
C3 VDD2 VDD1 1.13199f
C4 VN VTAIL 4.49243f
C5 VP VTAIL 4.50671f
C6 VN VDD1 0.15009f
C7 VN VDD2 4.35126f
C8 VP VDD1 4.59166f
C9 VP VDD2 0.39312f
C10 VDD2 B 4.686835f
C11 VDD1 B 4.970611f
C12 VTAIL B 5.801569f
C13 VN B 10.36742f
C14 VP B 8.936573f
C15 VDD1.t3 B 1.57642f
C16 VDD1.t4 B 1.5757f
C17 VDD1.t0 B 0.142376f
C18 VDD1.t2 B 0.142376f
C19 VDD1.n0 B 1.23689f
C20 VDD1.n1 B 2.1397f
C21 VDD1.t1 B 0.142376f
C22 VDD1.t5 B 0.142376f
C23 VDD1.n2 B 1.23468f
C24 VDD1.n3 B 2.00019f
C25 VP.n0 B 0.040511f
C26 VP.t3 B 1.23658f
C27 VP.n1 B 0.051471f
C28 VP.n2 B 0.030729f
C29 VP.t5 B 1.23658f
C30 VP.n3 B 0.037868f
C31 VP.n4 B 0.040511f
C32 VP.t0 B 1.23658f
C33 VP.n5 B 0.051471f
C34 VP.t2 B 1.36816f
C35 VP.n6 B 0.533816f
C36 VP.t4 B 1.23658f
C37 VP.n7 B 0.526424f
C38 VP.n8 B 0.042918f
C39 VP.n9 B 0.225317f
C40 VP.n10 B 0.030729f
C41 VP.n11 B 0.030729f
C42 VP.n12 B 0.037868f
C43 VP.n13 B 0.05192f
C44 VP.n14 B 0.544097f
C45 VP.n15 B 1.32992f
C46 VP.n16 B 1.35583f
C47 VP.t1 B 1.23658f
C48 VP.n17 B 0.544097f
C49 VP.n18 B 0.05192f
C50 VP.n19 B 0.040511f
C51 VP.n20 B 0.030729f
C52 VP.n21 B 0.030729f
C53 VP.n22 B 0.051471f
C54 VP.n23 B 0.042918f
C55 VP.n24 B 0.457836f
C56 VP.n25 B 0.042918f
C57 VP.n26 B 0.030729f
C58 VP.n27 B 0.030729f
C59 VP.n28 B 0.030729f
C60 VP.n29 B 0.037868f
C61 VP.n30 B 0.05192f
C62 VP.n31 B 0.544097f
C63 VP.n32 B 0.036224f
C64 VTAIL.t10 B 0.158811f
C65 VTAIL.t7 B 0.158811f
C66 VTAIL.n0 B 1.30974f
C67 VTAIL.n1 B 0.382841f
C68 VTAIL.t1 B 1.66591f
C69 VTAIL.n2 B 0.56575f
C70 VTAIL.t0 B 0.158811f
C71 VTAIL.t3 B 0.158811f
C72 VTAIL.n3 B 1.30974f
C73 VTAIL.n4 B 1.56468f
C74 VTAIL.t8 B 0.158811f
C75 VTAIL.t11 B 0.158811f
C76 VTAIL.n5 B 1.30975f
C77 VTAIL.n6 B 1.56468f
C78 VTAIL.t9 B 1.66592f
C79 VTAIL.n7 B 0.565738f
C80 VTAIL.t4 B 0.158811f
C81 VTAIL.t2 B 0.158811f
C82 VTAIL.n8 B 1.30975f
C83 VTAIL.n9 B 0.488787f
C84 VTAIL.t5 B 1.6659f
C85 VTAIL.n10 B 1.49423f
C86 VTAIL.t6 B 1.66591f
C87 VTAIL.n11 B 1.45278f
C88 VDD2.t5 B 1.55826f
C89 VDD2.t2 B 0.1408f
C90 VDD2.t1 B 0.1408f
C91 VDD2.n0 B 1.2232f
C92 VDD2.n1 B 2.02738f
C93 VDD2.t3 B 1.55173f
C94 VDD2.n2 B 1.98234f
C95 VDD2.t0 B 0.1408f
C96 VDD2.t4 B 0.1408f
C97 VDD2.n3 B 1.22317f
C98 VN.n0 B 0.039838f
C99 VN.t5 B 1.21605f
C100 VN.n1 B 0.050616f
C101 VN.t1 B 1.34544f
C102 VN.n2 B 0.52495f
C103 VN.t4 B 1.21605f
C104 VN.n3 B 0.517681f
C105 VN.n4 B 0.042205f
C106 VN.n5 B 0.221575f
C107 VN.n6 B 0.030218f
C108 VN.n7 B 0.030218f
C109 VN.n8 B 0.037239f
C110 VN.n9 B 0.051058f
C111 VN.n10 B 0.535061f
C112 VN.n11 B 0.035622f
C113 VN.n12 B 0.039838f
C114 VN.t3 B 1.21605f
C115 VN.n13 B 0.050616f
C116 VN.t2 B 1.34544f
C117 VN.n14 B 0.52495f
C118 VN.t0 B 1.21605f
C119 VN.n15 B 0.517681f
C120 VN.n16 B 0.042205f
C121 VN.n17 B 0.221575f
C122 VN.n18 B 0.030218f
C123 VN.n19 B 0.030218f
C124 VN.n20 B 0.037239f
C125 VN.n21 B 0.051058f
C126 VN.n22 B 0.535061f
C127 VN.n23 B 1.32451f
.ends

