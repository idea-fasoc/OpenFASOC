* NGSPICE file created from diff_pair_sample_0433.ext - technology: sky130A

.subckt diff_pair_sample_0433 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=0 ps=0 w=14.72 l=2.19
X1 VDD1.t3 VP.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4288 pd=15.05 as=5.7408 ps=30.22 w=14.72 l=2.19
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=0 ps=0 w=14.72 l=2.19
X3 VTAIL.t0 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=2.4288 ps=15.05 w=14.72 l=2.19
X4 VDD2.t2 VN.t1 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4288 pd=15.05 as=5.7408 ps=30.22 w=14.72 l=2.19
X5 VDD1.t2 VP.t1 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4288 pd=15.05 as=5.7408 ps=30.22 w=14.72 l=2.19
X6 VDD2.t1 VN.t2 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4288 pd=15.05 as=5.7408 ps=30.22 w=14.72 l=2.19
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=0 ps=0 w=14.72 l=2.19
X8 VTAIL.t2 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=2.4288 ps=15.05 w=14.72 l=2.19
X9 VTAIL.t4 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=2.4288 ps=15.05 w=14.72 l=2.19
X10 VTAIL.t6 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=2.4288 ps=15.05 w=14.72 l=2.19
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7408 pd=30.22 as=0 ps=0 w=14.72 l=2.19
R0 B.n585 B.n584 585
R1 B.n585 B.n58 585
R2 B.n588 B.n587 585
R3 B.n589 B.n117 585
R4 B.n591 B.n590 585
R5 B.n593 B.n116 585
R6 B.n596 B.n595 585
R7 B.n597 B.n115 585
R8 B.n599 B.n598 585
R9 B.n601 B.n114 585
R10 B.n604 B.n603 585
R11 B.n605 B.n113 585
R12 B.n607 B.n606 585
R13 B.n609 B.n112 585
R14 B.n612 B.n611 585
R15 B.n613 B.n111 585
R16 B.n615 B.n614 585
R17 B.n617 B.n110 585
R18 B.n620 B.n619 585
R19 B.n621 B.n109 585
R20 B.n623 B.n622 585
R21 B.n625 B.n108 585
R22 B.n628 B.n627 585
R23 B.n629 B.n107 585
R24 B.n631 B.n630 585
R25 B.n633 B.n106 585
R26 B.n636 B.n635 585
R27 B.n637 B.n105 585
R28 B.n639 B.n638 585
R29 B.n641 B.n104 585
R30 B.n644 B.n643 585
R31 B.n645 B.n103 585
R32 B.n647 B.n646 585
R33 B.n649 B.n102 585
R34 B.n652 B.n651 585
R35 B.n653 B.n101 585
R36 B.n655 B.n654 585
R37 B.n657 B.n100 585
R38 B.n660 B.n659 585
R39 B.n661 B.n99 585
R40 B.n663 B.n662 585
R41 B.n665 B.n98 585
R42 B.n668 B.n667 585
R43 B.n669 B.n97 585
R44 B.n671 B.n670 585
R45 B.n673 B.n96 585
R46 B.n676 B.n675 585
R47 B.n677 B.n95 585
R48 B.n679 B.n678 585
R49 B.n681 B.n94 585
R50 B.n684 B.n683 585
R51 B.n686 B.n91 585
R52 B.n688 B.n687 585
R53 B.n690 B.n90 585
R54 B.n693 B.n692 585
R55 B.n694 B.n89 585
R56 B.n696 B.n695 585
R57 B.n698 B.n88 585
R58 B.n700 B.n699 585
R59 B.n702 B.n701 585
R60 B.n705 B.n704 585
R61 B.n706 B.n83 585
R62 B.n708 B.n707 585
R63 B.n710 B.n82 585
R64 B.n713 B.n712 585
R65 B.n714 B.n81 585
R66 B.n716 B.n715 585
R67 B.n718 B.n80 585
R68 B.n721 B.n720 585
R69 B.n722 B.n79 585
R70 B.n724 B.n723 585
R71 B.n726 B.n78 585
R72 B.n729 B.n728 585
R73 B.n730 B.n77 585
R74 B.n732 B.n731 585
R75 B.n734 B.n76 585
R76 B.n737 B.n736 585
R77 B.n738 B.n75 585
R78 B.n740 B.n739 585
R79 B.n742 B.n74 585
R80 B.n745 B.n744 585
R81 B.n746 B.n73 585
R82 B.n748 B.n747 585
R83 B.n750 B.n72 585
R84 B.n753 B.n752 585
R85 B.n754 B.n71 585
R86 B.n756 B.n755 585
R87 B.n758 B.n70 585
R88 B.n761 B.n760 585
R89 B.n762 B.n69 585
R90 B.n764 B.n763 585
R91 B.n766 B.n68 585
R92 B.n769 B.n768 585
R93 B.n770 B.n67 585
R94 B.n772 B.n771 585
R95 B.n774 B.n66 585
R96 B.n777 B.n776 585
R97 B.n778 B.n65 585
R98 B.n780 B.n779 585
R99 B.n782 B.n64 585
R100 B.n785 B.n784 585
R101 B.n786 B.n63 585
R102 B.n788 B.n787 585
R103 B.n790 B.n62 585
R104 B.n793 B.n792 585
R105 B.n794 B.n61 585
R106 B.n796 B.n795 585
R107 B.n798 B.n60 585
R108 B.n801 B.n800 585
R109 B.n802 B.n59 585
R110 B.n583 B.n57 585
R111 B.n805 B.n57 585
R112 B.n582 B.n56 585
R113 B.n806 B.n56 585
R114 B.n581 B.n55 585
R115 B.n807 B.n55 585
R116 B.n580 B.n579 585
R117 B.n579 B.n51 585
R118 B.n578 B.n50 585
R119 B.n813 B.n50 585
R120 B.n577 B.n49 585
R121 B.n814 B.n49 585
R122 B.n576 B.n48 585
R123 B.n815 B.n48 585
R124 B.n575 B.n574 585
R125 B.n574 B.n47 585
R126 B.n573 B.n43 585
R127 B.n821 B.n43 585
R128 B.n572 B.n42 585
R129 B.n822 B.n42 585
R130 B.n571 B.n41 585
R131 B.n823 B.n41 585
R132 B.n570 B.n569 585
R133 B.n569 B.n37 585
R134 B.n568 B.n36 585
R135 B.n829 B.n36 585
R136 B.n567 B.n35 585
R137 B.n830 B.n35 585
R138 B.n566 B.n34 585
R139 B.n831 B.n34 585
R140 B.n565 B.n564 585
R141 B.n564 B.n30 585
R142 B.n563 B.n29 585
R143 B.n837 B.n29 585
R144 B.n562 B.n28 585
R145 B.n838 B.n28 585
R146 B.n561 B.n27 585
R147 B.n839 B.n27 585
R148 B.n560 B.n559 585
R149 B.n559 B.n23 585
R150 B.n558 B.n22 585
R151 B.n845 B.n22 585
R152 B.n557 B.n21 585
R153 B.n846 B.n21 585
R154 B.n556 B.n20 585
R155 B.n847 B.n20 585
R156 B.n555 B.n554 585
R157 B.n554 B.n16 585
R158 B.n553 B.n15 585
R159 B.n853 B.n15 585
R160 B.n552 B.n14 585
R161 B.n854 B.n14 585
R162 B.n551 B.n13 585
R163 B.n855 B.n13 585
R164 B.n550 B.n549 585
R165 B.n549 B.n12 585
R166 B.n548 B.n547 585
R167 B.n548 B.n8 585
R168 B.n546 B.n7 585
R169 B.n862 B.n7 585
R170 B.n545 B.n6 585
R171 B.n863 B.n6 585
R172 B.n544 B.n5 585
R173 B.n864 B.n5 585
R174 B.n543 B.n542 585
R175 B.n542 B.n4 585
R176 B.n541 B.n118 585
R177 B.n541 B.n540 585
R178 B.n531 B.n119 585
R179 B.n120 B.n119 585
R180 B.n533 B.n532 585
R181 B.n534 B.n533 585
R182 B.n530 B.n124 585
R183 B.n128 B.n124 585
R184 B.n529 B.n528 585
R185 B.n528 B.n527 585
R186 B.n126 B.n125 585
R187 B.n127 B.n126 585
R188 B.n520 B.n519 585
R189 B.n521 B.n520 585
R190 B.n518 B.n133 585
R191 B.n133 B.n132 585
R192 B.n517 B.n516 585
R193 B.n516 B.n515 585
R194 B.n135 B.n134 585
R195 B.n136 B.n135 585
R196 B.n508 B.n507 585
R197 B.n509 B.n508 585
R198 B.n506 B.n140 585
R199 B.n144 B.n140 585
R200 B.n505 B.n504 585
R201 B.n504 B.n503 585
R202 B.n142 B.n141 585
R203 B.n143 B.n142 585
R204 B.n496 B.n495 585
R205 B.n497 B.n496 585
R206 B.n494 B.n149 585
R207 B.n149 B.n148 585
R208 B.n493 B.n492 585
R209 B.n492 B.n491 585
R210 B.n151 B.n150 585
R211 B.n152 B.n151 585
R212 B.n484 B.n483 585
R213 B.n485 B.n484 585
R214 B.n482 B.n157 585
R215 B.n157 B.n156 585
R216 B.n481 B.n480 585
R217 B.n480 B.n479 585
R218 B.n159 B.n158 585
R219 B.n472 B.n159 585
R220 B.n471 B.n470 585
R221 B.n473 B.n471 585
R222 B.n469 B.n164 585
R223 B.n164 B.n163 585
R224 B.n468 B.n467 585
R225 B.n467 B.n466 585
R226 B.n166 B.n165 585
R227 B.n167 B.n166 585
R228 B.n459 B.n458 585
R229 B.n460 B.n459 585
R230 B.n457 B.n172 585
R231 B.n172 B.n171 585
R232 B.n456 B.n455 585
R233 B.n455 B.n454 585
R234 B.n451 B.n176 585
R235 B.n450 B.n449 585
R236 B.n447 B.n177 585
R237 B.n447 B.n175 585
R238 B.n446 B.n445 585
R239 B.n444 B.n443 585
R240 B.n442 B.n179 585
R241 B.n440 B.n439 585
R242 B.n438 B.n180 585
R243 B.n437 B.n436 585
R244 B.n434 B.n181 585
R245 B.n432 B.n431 585
R246 B.n430 B.n182 585
R247 B.n429 B.n428 585
R248 B.n426 B.n183 585
R249 B.n424 B.n423 585
R250 B.n422 B.n184 585
R251 B.n421 B.n420 585
R252 B.n418 B.n185 585
R253 B.n416 B.n415 585
R254 B.n414 B.n186 585
R255 B.n413 B.n412 585
R256 B.n410 B.n187 585
R257 B.n408 B.n407 585
R258 B.n406 B.n188 585
R259 B.n405 B.n404 585
R260 B.n402 B.n189 585
R261 B.n400 B.n399 585
R262 B.n398 B.n190 585
R263 B.n397 B.n396 585
R264 B.n394 B.n191 585
R265 B.n392 B.n391 585
R266 B.n390 B.n192 585
R267 B.n389 B.n388 585
R268 B.n386 B.n193 585
R269 B.n384 B.n383 585
R270 B.n382 B.n194 585
R271 B.n381 B.n380 585
R272 B.n378 B.n195 585
R273 B.n376 B.n375 585
R274 B.n374 B.n196 585
R275 B.n373 B.n372 585
R276 B.n370 B.n197 585
R277 B.n368 B.n367 585
R278 B.n366 B.n198 585
R279 B.n365 B.n364 585
R280 B.n362 B.n199 585
R281 B.n360 B.n359 585
R282 B.n358 B.n200 585
R283 B.n357 B.n356 585
R284 B.n354 B.n201 585
R285 B.n352 B.n351 585
R286 B.n350 B.n202 585
R287 B.n349 B.n348 585
R288 B.n346 B.n206 585
R289 B.n344 B.n343 585
R290 B.n342 B.n207 585
R291 B.n341 B.n340 585
R292 B.n338 B.n208 585
R293 B.n336 B.n335 585
R294 B.n333 B.n209 585
R295 B.n332 B.n331 585
R296 B.n329 B.n212 585
R297 B.n327 B.n326 585
R298 B.n325 B.n213 585
R299 B.n324 B.n323 585
R300 B.n321 B.n214 585
R301 B.n319 B.n318 585
R302 B.n317 B.n215 585
R303 B.n316 B.n315 585
R304 B.n313 B.n216 585
R305 B.n311 B.n310 585
R306 B.n309 B.n217 585
R307 B.n308 B.n307 585
R308 B.n305 B.n218 585
R309 B.n303 B.n302 585
R310 B.n301 B.n219 585
R311 B.n300 B.n299 585
R312 B.n297 B.n220 585
R313 B.n295 B.n294 585
R314 B.n293 B.n221 585
R315 B.n292 B.n291 585
R316 B.n289 B.n222 585
R317 B.n287 B.n286 585
R318 B.n285 B.n223 585
R319 B.n284 B.n283 585
R320 B.n281 B.n224 585
R321 B.n279 B.n278 585
R322 B.n277 B.n225 585
R323 B.n276 B.n275 585
R324 B.n273 B.n226 585
R325 B.n271 B.n270 585
R326 B.n269 B.n227 585
R327 B.n268 B.n267 585
R328 B.n265 B.n228 585
R329 B.n263 B.n262 585
R330 B.n261 B.n229 585
R331 B.n260 B.n259 585
R332 B.n257 B.n230 585
R333 B.n255 B.n254 585
R334 B.n253 B.n231 585
R335 B.n252 B.n251 585
R336 B.n249 B.n232 585
R337 B.n247 B.n246 585
R338 B.n245 B.n233 585
R339 B.n244 B.n243 585
R340 B.n241 B.n234 585
R341 B.n239 B.n238 585
R342 B.n237 B.n236 585
R343 B.n174 B.n173 585
R344 B.n453 B.n452 585
R345 B.n454 B.n453 585
R346 B.n170 B.n169 585
R347 B.n171 B.n170 585
R348 B.n462 B.n461 585
R349 B.n461 B.n460 585
R350 B.n463 B.n168 585
R351 B.n168 B.n167 585
R352 B.n465 B.n464 585
R353 B.n466 B.n465 585
R354 B.n162 B.n161 585
R355 B.n163 B.n162 585
R356 B.n475 B.n474 585
R357 B.n474 B.n473 585
R358 B.n476 B.n160 585
R359 B.n472 B.n160 585
R360 B.n478 B.n477 585
R361 B.n479 B.n478 585
R362 B.n155 B.n154 585
R363 B.n156 B.n155 585
R364 B.n487 B.n486 585
R365 B.n486 B.n485 585
R366 B.n488 B.n153 585
R367 B.n153 B.n152 585
R368 B.n490 B.n489 585
R369 B.n491 B.n490 585
R370 B.n147 B.n146 585
R371 B.n148 B.n147 585
R372 B.n499 B.n498 585
R373 B.n498 B.n497 585
R374 B.n500 B.n145 585
R375 B.n145 B.n143 585
R376 B.n502 B.n501 585
R377 B.n503 B.n502 585
R378 B.n139 B.n138 585
R379 B.n144 B.n139 585
R380 B.n511 B.n510 585
R381 B.n510 B.n509 585
R382 B.n512 B.n137 585
R383 B.n137 B.n136 585
R384 B.n514 B.n513 585
R385 B.n515 B.n514 585
R386 B.n131 B.n130 585
R387 B.n132 B.n131 585
R388 B.n523 B.n522 585
R389 B.n522 B.n521 585
R390 B.n524 B.n129 585
R391 B.n129 B.n127 585
R392 B.n526 B.n525 585
R393 B.n527 B.n526 585
R394 B.n123 B.n122 585
R395 B.n128 B.n123 585
R396 B.n536 B.n535 585
R397 B.n535 B.n534 585
R398 B.n537 B.n121 585
R399 B.n121 B.n120 585
R400 B.n539 B.n538 585
R401 B.n540 B.n539 585
R402 B.n3 B.n0 585
R403 B.n4 B.n3 585
R404 B.n861 B.n1 585
R405 B.n862 B.n861 585
R406 B.n860 B.n859 585
R407 B.n860 B.n8 585
R408 B.n858 B.n9 585
R409 B.n12 B.n9 585
R410 B.n857 B.n856 585
R411 B.n856 B.n855 585
R412 B.n11 B.n10 585
R413 B.n854 B.n11 585
R414 B.n852 B.n851 585
R415 B.n853 B.n852 585
R416 B.n850 B.n17 585
R417 B.n17 B.n16 585
R418 B.n849 B.n848 585
R419 B.n848 B.n847 585
R420 B.n19 B.n18 585
R421 B.n846 B.n19 585
R422 B.n844 B.n843 585
R423 B.n845 B.n844 585
R424 B.n842 B.n24 585
R425 B.n24 B.n23 585
R426 B.n841 B.n840 585
R427 B.n840 B.n839 585
R428 B.n26 B.n25 585
R429 B.n838 B.n26 585
R430 B.n836 B.n835 585
R431 B.n837 B.n836 585
R432 B.n834 B.n31 585
R433 B.n31 B.n30 585
R434 B.n833 B.n832 585
R435 B.n832 B.n831 585
R436 B.n33 B.n32 585
R437 B.n830 B.n33 585
R438 B.n828 B.n827 585
R439 B.n829 B.n828 585
R440 B.n826 B.n38 585
R441 B.n38 B.n37 585
R442 B.n825 B.n824 585
R443 B.n824 B.n823 585
R444 B.n40 B.n39 585
R445 B.n822 B.n40 585
R446 B.n820 B.n819 585
R447 B.n821 B.n820 585
R448 B.n818 B.n44 585
R449 B.n47 B.n44 585
R450 B.n817 B.n816 585
R451 B.n816 B.n815 585
R452 B.n46 B.n45 585
R453 B.n814 B.n46 585
R454 B.n812 B.n811 585
R455 B.n813 B.n812 585
R456 B.n810 B.n52 585
R457 B.n52 B.n51 585
R458 B.n809 B.n808 585
R459 B.n808 B.n807 585
R460 B.n54 B.n53 585
R461 B.n806 B.n54 585
R462 B.n804 B.n803 585
R463 B.n805 B.n804 585
R464 B.n865 B.n864 585
R465 B.n863 B.n2 585
R466 B.n804 B.n59 458.866
R467 B.n585 B.n57 458.866
R468 B.n455 B.n174 458.866
R469 B.n453 B.n176 458.866
R470 B.n92 B.t16 377.731
R471 B.n210 B.t7 377.731
R472 B.n84 B.t13 377.731
R473 B.n203 B.t10 377.731
R474 B.n84 B.t11 369.318
R475 B.n92 B.t15 369.318
R476 B.n210 B.t4 369.318
R477 B.n203 B.t8 369.318
R478 B.n93 B.t17 328.858
R479 B.n211 B.t6 328.858
R480 B.n85 B.t14 328.858
R481 B.n204 B.t9 328.858
R482 B.n586 B.n58 256.663
R483 B.n592 B.n58 256.663
R484 B.n594 B.n58 256.663
R485 B.n600 B.n58 256.663
R486 B.n602 B.n58 256.663
R487 B.n608 B.n58 256.663
R488 B.n610 B.n58 256.663
R489 B.n616 B.n58 256.663
R490 B.n618 B.n58 256.663
R491 B.n624 B.n58 256.663
R492 B.n626 B.n58 256.663
R493 B.n632 B.n58 256.663
R494 B.n634 B.n58 256.663
R495 B.n640 B.n58 256.663
R496 B.n642 B.n58 256.663
R497 B.n648 B.n58 256.663
R498 B.n650 B.n58 256.663
R499 B.n656 B.n58 256.663
R500 B.n658 B.n58 256.663
R501 B.n664 B.n58 256.663
R502 B.n666 B.n58 256.663
R503 B.n672 B.n58 256.663
R504 B.n674 B.n58 256.663
R505 B.n680 B.n58 256.663
R506 B.n682 B.n58 256.663
R507 B.n689 B.n58 256.663
R508 B.n691 B.n58 256.663
R509 B.n697 B.n58 256.663
R510 B.n87 B.n58 256.663
R511 B.n703 B.n58 256.663
R512 B.n709 B.n58 256.663
R513 B.n711 B.n58 256.663
R514 B.n717 B.n58 256.663
R515 B.n719 B.n58 256.663
R516 B.n725 B.n58 256.663
R517 B.n727 B.n58 256.663
R518 B.n733 B.n58 256.663
R519 B.n735 B.n58 256.663
R520 B.n741 B.n58 256.663
R521 B.n743 B.n58 256.663
R522 B.n749 B.n58 256.663
R523 B.n751 B.n58 256.663
R524 B.n757 B.n58 256.663
R525 B.n759 B.n58 256.663
R526 B.n765 B.n58 256.663
R527 B.n767 B.n58 256.663
R528 B.n773 B.n58 256.663
R529 B.n775 B.n58 256.663
R530 B.n781 B.n58 256.663
R531 B.n783 B.n58 256.663
R532 B.n789 B.n58 256.663
R533 B.n791 B.n58 256.663
R534 B.n797 B.n58 256.663
R535 B.n799 B.n58 256.663
R536 B.n448 B.n175 256.663
R537 B.n178 B.n175 256.663
R538 B.n441 B.n175 256.663
R539 B.n435 B.n175 256.663
R540 B.n433 B.n175 256.663
R541 B.n427 B.n175 256.663
R542 B.n425 B.n175 256.663
R543 B.n419 B.n175 256.663
R544 B.n417 B.n175 256.663
R545 B.n411 B.n175 256.663
R546 B.n409 B.n175 256.663
R547 B.n403 B.n175 256.663
R548 B.n401 B.n175 256.663
R549 B.n395 B.n175 256.663
R550 B.n393 B.n175 256.663
R551 B.n387 B.n175 256.663
R552 B.n385 B.n175 256.663
R553 B.n379 B.n175 256.663
R554 B.n377 B.n175 256.663
R555 B.n371 B.n175 256.663
R556 B.n369 B.n175 256.663
R557 B.n363 B.n175 256.663
R558 B.n361 B.n175 256.663
R559 B.n355 B.n175 256.663
R560 B.n353 B.n175 256.663
R561 B.n347 B.n175 256.663
R562 B.n345 B.n175 256.663
R563 B.n339 B.n175 256.663
R564 B.n337 B.n175 256.663
R565 B.n330 B.n175 256.663
R566 B.n328 B.n175 256.663
R567 B.n322 B.n175 256.663
R568 B.n320 B.n175 256.663
R569 B.n314 B.n175 256.663
R570 B.n312 B.n175 256.663
R571 B.n306 B.n175 256.663
R572 B.n304 B.n175 256.663
R573 B.n298 B.n175 256.663
R574 B.n296 B.n175 256.663
R575 B.n290 B.n175 256.663
R576 B.n288 B.n175 256.663
R577 B.n282 B.n175 256.663
R578 B.n280 B.n175 256.663
R579 B.n274 B.n175 256.663
R580 B.n272 B.n175 256.663
R581 B.n266 B.n175 256.663
R582 B.n264 B.n175 256.663
R583 B.n258 B.n175 256.663
R584 B.n256 B.n175 256.663
R585 B.n250 B.n175 256.663
R586 B.n248 B.n175 256.663
R587 B.n242 B.n175 256.663
R588 B.n240 B.n175 256.663
R589 B.n235 B.n175 256.663
R590 B.n867 B.n866 256.663
R591 B.n800 B.n798 163.367
R592 B.n796 B.n61 163.367
R593 B.n792 B.n790 163.367
R594 B.n788 B.n63 163.367
R595 B.n784 B.n782 163.367
R596 B.n780 B.n65 163.367
R597 B.n776 B.n774 163.367
R598 B.n772 B.n67 163.367
R599 B.n768 B.n766 163.367
R600 B.n764 B.n69 163.367
R601 B.n760 B.n758 163.367
R602 B.n756 B.n71 163.367
R603 B.n752 B.n750 163.367
R604 B.n748 B.n73 163.367
R605 B.n744 B.n742 163.367
R606 B.n740 B.n75 163.367
R607 B.n736 B.n734 163.367
R608 B.n732 B.n77 163.367
R609 B.n728 B.n726 163.367
R610 B.n724 B.n79 163.367
R611 B.n720 B.n718 163.367
R612 B.n716 B.n81 163.367
R613 B.n712 B.n710 163.367
R614 B.n708 B.n83 163.367
R615 B.n704 B.n702 163.367
R616 B.n699 B.n698 163.367
R617 B.n696 B.n89 163.367
R618 B.n692 B.n690 163.367
R619 B.n688 B.n91 163.367
R620 B.n683 B.n681 163.367
R621 B.n679 B.n95 163.367
R622 B.n675 B.n673 163.367
R623 B.n671 B.n97 163.367
R624 B.n667 B.n665 163.367
R625 B.n663 B.n99 163.367
R626 B.n659 B.n657 163.367
R627 B.n655 B.n101 163.367
R628 B.n651 B.n649 163.367
R629 B.n647 B.n103 163.367
R630 B.n643 B.n641 163.367
R631 B.n639 B.n105 163.367
R632 B.n635 B.n633 163.367
R633 B.n631 B.n107 163.367
R634 B.n627 B.n625 163.367
R635 B.n623 B.n109 163.367
R636 B.n619 B.n617 163.367
R637 B.n615 B.n111 163.367
R638 B.n611 B.n609 163.367
R639 B.n607 B.n113 163.367
R640 B.n603 B.n601 163.367
R641 B.n599 B.n115 163.367
R642 B.n595 B.n593 163.367
R643 B.n591 B.n117 163.367
R644 B.n587 B.n585 163.367
R645 B.n455 B.n172 163.367
R646 B.n459 B.n172 163.367
R647 B.n459 B.n166 163.367
R648 B.n467 B.n166 163.367
R649 B.n467 B.n164 163.367
R650 B.n471 B.n164 163.367
R651 B.n471 B.n159 163.367
R652 B.n480 B.n159 163.367
R653 B.n480 B.n157 163.367
R654 B.n484 B.n157 163.367
R655 B.n484 B.n151 163.367
R656 B.n492 B.n151 163.367
R657 B.n492 B.n149 163.367
R658 B.n496 B.n149 163.367
R659 B.n496 B.n142 163.367
R660 B.n504 B.n142 163.367
R661 B.n504 B.n140 163.367
R662 B.n508 B.n140 163.367
R663 B.n508 B.n135 163.367
R664 B.n516 B.n135 163.367
R665 B.n516 B.n133 163.367
R666 B.n520 B.n133 163.367
R667 B.n520 B.n126 163.367
R668 B.n528 B.n126 163.367
R669 B.n528 B.n124 163.367
R670 B.n533 B.n124 163.367
R671 B.n533 B.n119 163.367
R672 B.n541 B.n119 163.367
R673 B.n542 B.n541 163.367
R674 B.n542 B.n5 163.367
R675 B.n6 B.n5 163.367
R676 B.n7 B.n6 163.367
R677 B.n548 B.n7 163.367
R678 B.n549 B.n548 163.367
R679 B.n549 B.n13 163.367
R680 B.n14 B.n13 163.367
R681 B.n15 B.n14 163.367
R682 B.n554 B.n15 163.367
R683 B.n554 B.n20 163.367
R684 B.n21 B.n20 163.367
R685 B.n22 B.n21 163.367
R686 B.n559 B.n22 163.367
R687 B.n559 B.n27 163.367
R688 B.n28 B.n27 163.367
R689 B.n29 B.n28 163.367
R690 B.n564 B.n29 163.367
R691 B.n564 B.n34 163.367
R692 B.n35 B.n34 163.367
R693 B.n36 B.n35 163.367
R694 B.n569 B.n36 163.367
R695 B.n569 B.n41 163.367
R696 B.n42 B.n41 163.367
R697 B.n43 B.n42 163.367
R698 B.n574 B.n43 163.367
R699 B.n574 B.n48 163.367
R700 B.n49 B.n48 163.367
R701 B.n50 B.n49 163.367
R702 B.n579 B.n50 163.367
R703 B.n579 B.n55 163.367
R704 B.n56 B.n55 163.367
R705 B.n57 B.n56 163.367
R706 B.n449 B.n447 163.367
R707 B.n447 B.n446 163.367
R708 B.n443 B.n442 163.367
R709 B.n440 B.n180 163.367
R710 B.n436 B.n434 163.367
R711 B.n432 B.n182 163.367
R712 B.n428 B.n426 163.367
R713 B.n424 B.n184 163.367
R714 B.n420 B.n418 163.367
R715 B.n416 B.n186 163.367
R716 B.n412 B.n410 163.367
R717 B.n408 B.n188 163.367
R718 B.n404 B.n402 163.367
R719 B.n400 B.n190 163.367
R720 B.n396 B.n394 163.367
R721 B.n392 B.n192 163.367
R722 B.n388 B.n386 163.367
R723 B.n384 B.n194 163.367
R724 B.n380 B.n378 163.367
R725 B.n376 B.n196 163.367
R726 B.n372 B.n370 163.367
R727 B.n368 B.n198 163.367
R728 B.n364 B.n362 163.367
R729 B.n360 B.n200 163.367
R730 B.n356 B.n354 163.367
R731 B.n352 B.n202 163.367
R732 B.n348 B.n346 163.367
R733 B.n344 B.n207 163.367
R734 B.n340 B.n338 163.367
R735 B.n336 B.n209 163.367
R736 B.n331 B.n329 163.367
R737 B.n327 B.n213 163.367
R738 B.n323 B.n321 163.367
R739 B.n319 B.n215 163.367
R740 B.n315 B.n313 163.367
R741 B.n311 B.n217 163.367
R742 B.n307 B.n305 163.367
R743 B.n303 B.n219 163.367
R744 B.n299 B.n297 163.367
R745 B.n295 B.n221 163.367
R746 B.n291 B.n289 163.367
R747 B.n287 B.n223 163.367
R748 B.n283 B.n281 163.367
R749 B.n279 B.n225 163.367
R750 B.n275 B.n273 163.367
R751 B.n271 B.n227 163.367
R752 B.n267 B.n265 163.367
R753 B.n263 B.n229 163.367
R754 B.n259 B.n257 163.367
R755 B.n255 B.n231 163.367
R756 B.n251 B.n249 163.367
R757 B.n247 B.n233 163.367
R758 B.n243 B.n241 163.367
R759 B.n239 B.n236 163.367
R760 B.n453 B.n170 163.367
R761 B.n461 B.n170 163.367
R762 B.n461 B.n168 163.367
R763 B.n465 B.n168 163.367
R764 B.n465 B.n162 163.367
R765 B.n474 B.n162 163.367
R766 B.n474 B.n160 163.367
R767 B.n478 B.n160 163.367
R768 B.n478 B.n155 163.367
R769 B.n486 B.n155 163.367
R770 B.n486 B.n153 163.367
R771 B.n490 B.n153 163.367
R772 B.n490 B.n147 163.367
R773 B.n498 B.n147 163.367
R774 B.n498 B.n145 163.367
R775 B.n502 B.n145 163.367
R776 B.n502 B.n139 163.367
R777 B.n510 B.n139 163.367
R778 B.n510 B.n137 163.367
R779 B.n514 B.n137 163.367
R780 B.n514 B.n131 163.367
R781 B.n522 B.n131 163.367
R782 B.n522 B.n129 163.367
R783 B.n526 B.n129 163.367
R784 B.n526 B.n123 163.367
R785 B.n535 B.n123 163.367
R786 B.n535 B.n121 163.367
R787 B.n539 B.n121 163.367
R788 B.n539 B.n3 163.367
R789 B.n865 B.n3 163.367
R790 B.n861 B.n2 163.367
R791 B.n861 B.n860 163.367
R792 B.n860 B.n9 163.367
R793 B.n856 B.n9 163.367
R794 B.n856 B.n11 163.367
R795 B.n852 B.n11 163.367
R796 B.n852 B.n17 163.367
R797 B.n848 B.n17 163.367
R798 B.n848 B.n19 163.367
R799 B.n844 B.n19 163.367
R800 B.n844 B.n24 163.367
R801 B.n840 B.n24 163.367
R802 B.n840 B.n26 163.367
R803 B.n836 B.n26 163.367
R804 B.n836 B.n31 163.367
R805 B.n832 B.n31 163.367
R806 B.n832 B.n33 163.367
R807 B.n828 B.n33 163.367
R808 B.n828 B.n38 163.367
R809 B.n824 B.n38 163.367
R810 B.n824 B.n40 163.367
R811 B.n820 B.n40 163.367
R812 B.n820 B.n44 163.367
R813 B.n816 B.n44 163.367
R814 B.n816 B.n46 163.367
R815 B.n812 B.n46 163.367
R816 B.n812 B.n52 163.367
R817 B.n808 B.n52 163.367
R818 B.n808 B.n54 163.367
R819 B.n804 B.n54 163.367
R820 B.n799 B.n59 71.676
R821 B.n798 B.n797 71.676
R822 B.n791 B.n61 71.676
R823 B.n790 B.n789 71.676
R824 B.n783 B.n63 71.676
R825 B.n782 B.n781 71.676
R826 B.n775 B.n65 71.676
R827 B.n774 B.n773 71.676
R828 B.n767 B.n67 71.676
R829 B.n766 B.n765 71.676
R830 B.n759 B.n69 71.676
R831 B.n758 B.n757 71.676
R832 B.n751 B.n71 71.676
R833 B.n750 B.n749 71.676
R834 B.n743 B.n73 71.676
R835 B.n742 B.n741 71.676
R836 B.n735 B.n75 71.676
R837 B.n734 B.n733 71.676
R838 B.n727 B.n77 71.676
R839 B.n726 B.n725 71.676
R840 B.n719 B.n79 71.676
R841 B.n718 B.n717 71.676
R842 B.n711 B.n81 71.676
R843 B.n710 B.n709 71.676
R844 B.n703 B.n83 71.676
R845 B.n702 B.n87 71.676
R846 B.n698 B.n697 71.676
R847 B.n691 B.n89 71.676
R848 B.n690 B.n689 71.676
R849 B.n682 B.n91 71.676
R850 B.n681 B.n680 71.676
R851 B.n674 B.n95 71.676
R852 B.n673 B.n672 71.676
R853 B.n666 B.n97 71.676
R854 B.n665 B.n664 71.676
R855 B.n658 B.n99 71.676
R856 B.n657 B.n656 71.676
R857 B.n650 B.n101 71.676
R858 B.n649 B.n648 71.676
R859 B.n642 B.n103 71.676
R860 B.n641 B.n640 71.676
R861 B.n634 B.n105 71.676
R862 B.n633 B.n632 71.676
R863 B.n626 B.n107 71.676
R864 B.n625 B.n624 71.676
R865 B.n618 B.n109 71.676
R866 B.n617 B.n616 71.676
R867 B.n610 B.n111 71.676
R868 B.n609 B.n608 71.676
R869 B.n602 B.n113 71.676
R870 B.n601 B.n600 71.676
R871 B.n594 B.n115 71.676
R872 B.n593 B.n592 71.676
R873 B.n586 B.n117 71.676
R874 B.n587 B.n586 71.676
R875 B.n592 B.n591 71.676
R876 B.n595 B.n594 71.676
R877 B.n600 B.n599 71.676
R878 B.n603 B.n602 71.676
R879 B.n608 B.n607 71.676
R880 B.n611 B.n610 71.676
R881 B.n616 B.n615 71.676
R882 B.n619 B.n618 71.676
R883 B.n624 B.n623 71.676
R884 B.n627 B.n626 71.676
R885 B.n632 B.n631 71.676
R886 B.n635 B.n634 71.676
R887 B.n640 B.n639 71.676
R888 B.n643 B.n642 71.676
R889 B.n648 B.n647 71.676
R890 B.n651 B.n650 71.676
R891 B.n656 B.n655 71.676
R892 B.n659 B.n658 71.676
R893 B.n664 B.n663 71.676
R894 B.n667 B.n666 71.676
R895 B.n672 B.n671 71.676
R896 B.n675 B.n674 71.676
R897 B.n680 B.n679 71.676
R898 B.n683 B.n682 71.676
R899 B.n689 B.n688 71.676
R900 B.n692 B.n691 71.676
R901 B.n697 B.n696 71.676
R902 B.n699 B.n87 71.676
R903 B.n704 B.n703 71.676
R904 B.n709 B.n708 71.676
R905 B.n712 B.n711 71.676
R906 B.n717 B.n716 71.676
R907 B.n720 B.n719 71.676
R908 B.n725 B.n724 71.676
R909 B.n728 B.n727 71.676
R910 B.n733 B.n732 71.676
R911 B.n736 B.n735 71.676
R912 B.n741 B.n740 71.676
R913 B.n744 B.n743 71.676
R914 B.n749 B.n748 71.676
R915 B.n752 B.n751 71.676
R916 B.n757 B.n756 71.676
R917 B.n760 B.n759 71.676
R918 B.n765 B.n764 71.676
R919 B.n768 B.n767 71.676
R920 B.n773 B.n772 71.676
R921 B.n776 B.n775 71.676
R922 B.n781 B.n780 71.676
R923 B.n784 B.n783 71.676
R924 B.n789 B.n788 71.676
R925 B.n792 B.n791 71.676
R926 B.n797 B.n796 71.676
R927 B.n800 B.n799 71.676
R928 B.n448 B.n176 71.676
R929 B.n446 B.n178 71.676
R930 B.n442 B.n441 71.676
R931 B.n435 B.n180 71.676
R932 B.n434 B.n433 71.676
R933 B.n427 B.n182 71.676
R934 B.n426 B.n425 71.676
R935 B.n419 B.n184 71.676
R936 B.n418 B.n417 71.676
R937 B.n411 B.n186 71.676
R938 B.n410 B.n409 71.676
R939 B.n403 B.n188 71.676
R940 B.n402 B.n401 71.676
R941 B.n395 B.n190 71.676
R942 B.n394 B.n393 71.676
R943 B.n387 B.n192 71.676
R944 B.n386 B.n385 71.676
R945 B.n379 B.n194 71.676
R946 B.n378 B.n377 71.676
R947 B.n371 B.n196 71.676
R948 B.n370 B.n369 71.676
R949 B.n363 B.n198 71.676
R950 B.n362 B.n361 71.676
R951 B.n355 B.n200 71.676
R952 B.n354 B.n353 71.676
R953 B.n347 B.n202 71.676
R954 B.n346 B.n345 71.676
R955 B.n339 B.n207 71.676
R956 B.n338 B.n337 71.676
R957 B.n330 B.n209 71.676
R958 B.n329 B.n328 71.676
R959 B.n322 B.n213 71.676
R960 B.n321 B.n320 71.676
R961 B.n314 B.n215 71.676
R962 B.n313 B.n312 71.676
R963 B.n306 B.n217 71.676
R964 B.n305 B.n304 71.676
R965 B.n298 B.n219 71.676
R966 B.n297 B.n296 71.676
R967 B.n290 B.n221 71.676
R968 B.n289 B.n288 71.676
R969 B.n282 B.n223 71.676
R970 B.n281 B.n280 71.676
R971 B.n274 B.n225 71.676
R972 B.n273 B.n272 71.676
R973 B.n266 B.n227 71.676
R974 B.n265 B.n264 71.676
R975 B.n258 B.n229 71.676
R976 B.n257 B.n256 71.676
R977 B.n250 B.n231 71.676
R978 B.n249 B.n248 71.676
R979 B.n242 B.n233 71.676
R980 B.n241 B.n240 71.676
R981 B.n236 B.n235 71.676
R982 B.n449 B.n448 71.676
R983 B.n443 B.n178 71.676
R984 B.n441 B.n440 71.676
R985 B.n436 B.n435 71.676
R986 B.n433 B.n432 71.676
R987 B.n428 B.n427 71.676
R988 B.n425 B.n424 71.676
R989 B.n420 B.n419 71.676
R990 B.n417 B.n416 71.676
R991 B.n412 B.n411 71.676
R992 B.n409 B.n408 71.676
R993 B.n404 B.n403 71.676
R994 B.n401 B.n400 71.676
R995 B.n396 B.n395 71.676
R996 B.n393 B.n392 71.676
R997 B.n388 B.n387 71.676
R998 B.n385 B.n384 71.676
R999 B.n380 B.n379 71.676
R1000 B.n377 B.n376 71.676
R1001 B.n372 B.n371 71.676
R1002 B.n369 B.n368 71.676
R1003 B.n364 B.n363 71.676
R1004 B.n361 B.n360 71.676
R1005 B.n356 B.n355 71.676
R1006 B.n353 B.n352 71.676
R1007 B.n348 B.n347 71.676
R1008 B.n345 B.n344 71.676
R1009 B.n340 B.n339 71.676
R1010 B.n337 B.n336 71.676
R1011 B.n331 B.n330 71.676
R1012 B.n328 B.n327 71.676
R1013 B.n323 B.n322 71.676
R1014 B.n320 B.n319 71.676
R1015 B.n315 B.n314 71.676
R1016 B.n312 B.n311 71.676
R1017 B.n307 B.n306 71.676
R1018 B.n304 B.n303 71.676
R1019 B.n299 B.n298 71.676
R1020 B.n296 B.n295 71.676
R1021 B.n291 B.n290 71.676
R1022 B.n288 B.n287 71.676
R1023 B.n283 B.n282 71.676
R1024 B.n280 B.n279 71.676
R1025 B.n275 B.n274 71.676
R1026 B.n272 B.n271 71.676
R1027 B.n267 B.n266 71.676
R1028 B.n264 B.n263 71.676
R1029 B.n259 B.n258 71.676
R1030 B.n256 B.n255 71.676
R1031 B.n251 B.n250 71.676
R1032 B.n248 B.n247 71.676
R1033 B.n243 B.n242 71.676
R1034 B.n240 B.n239 71.676
R1035 B.n235 B.n174 71.676
R1036 B.n866 B.n865 71.676
R1037 B.n866 B.n2 71.676
R1038 B.n454 B.n175 62.166
R1039 B.n805 B.n58 62.166
R1040 B.n86 B.n85 59.5399
R1041 B.n685 B.n93 59.5399
R1042 B.n334 B.n211 59.5399
R1043 B.n205 B.n204 59.5399
R1044 B.n85 B.n84 48.8732
R1045 B.n93 B.n92 48.8732
R1046 B.n211 B.n210 48.8732
R1047 B.n204 B.n203 48.8732
R1048 B.n454 B.n171 37.4099
R1049 B.n460 B.n171 37.4099
R1050 B.n460 B.n167 37.4099
R1051 B.n466 B.n167 37.4099
R1052 B.n466 B.n163 37.4099
R1053 B.n473 B.n163 37.4099
R1054 B.n473 B.n472 37.4099
R1055 B.n479 B.n156 37.4099
R1056 B.n485 B.n156 37.4099
R1057 B.n485 B.n152 37.4099
R1058 B.n491 B.n152 37.4099
R1059 B.n491 B.n148 37.4099
R1060 B.n497 B.n148 37.4099
R1061 B.n497 B.n143 37.4099
R1062 B.n503 B.n143 37.4099
R1063 B.n503 B.n144 37.4099
R1064 B.n509 B.n136 37.4099
R1065 B.n515 B.n136 37.4099
R1066 B.n515 B.n132 37.4099
R1067 B.n521 B.n132 37.4099
R1068 B.n521 B.n127 37.4099
R1069 B.n527 B.n127 37.4099
R1070 B.n527 B.n128 37.4099
R1071 B.n534 B.n120 37.4099
R1072 B.n540 B.n120 37.4099
R1073 B.n540 B.n4 37.4099
R1074 B.n864 B.n4 37.4099
R1075 B.n864 B.n863 37.4099
R1076 B.n863 B.n862 37.4099
R1077 B.n862 B.n8 37.4099
R1078 B.n12 B.n8 37.4099
R1079 B.n855 B.n12 37.4099
R1080 B.n854 B.n853 37.4099
R1081 B.n853 B.n16 37.4099
R1082 B.n847 B.n16 37.4099
R1083 B.n847 B.n846 37.4099
R1084 B.n846 B.n845 37.4099
R1085 B.n845 B.n23 37.4099
R1086 B.n839 B.n23 37.4099
R1087 B.n838 B.n837 37.4099
R1088 B.n837 B.n30 37.4099
R1089 B.n831 B.n30 37.4099
R1090 B.n831 B.n830 37.4099
R1091 B.n830 B.n829 37.4099
R1092 B.n829 B.n37 37.4099
R1093 B.n823 B.n37 37.4099
R1094 B.n823 B.n822 37.4099
R1095 B.n822 B.n821 37.4099
R1096 B.n815 B.n47 37.4099
R1097 B.n815 B.n814 37.4099
R1098 B.n814 B.n813 37.4099
R1099 B.n813 B.n51 37.4099
R1100 B.n807 B.n51 37.4099
R1101 B.n807 B.n806 37.4099
R1102 B.n806 B.n805 37.4099
R1103 B.n479 B.t5 31.3583
R1104 B.n821 B.t12 31.3583
R1105 B.n534 B.t1 30.2581
R1106 B.n855 B.t3 30.2581
R1107 B.n452 B.n451 29.8151
R1108 B.n456 B.n173 29.8151
R1109 B.n584 B.n583 29.8151
R1110 B.n803 B.n802 29.8151
R1111 B.n144 B.t0 29.1578
R1112 B.t2 B.n838 29.1578
R1113 B B.n867 18.0485
R1114 B.n452 B.n169 10.6151
R1115 B.n462 B.n169 10.6151
R1116 B.n463 B.n462 10.6151
R1117 B.n464 B.n463 10.6151
R1118 B.n464 B.n161 10.6151
R1119 B.n475 B.n161 10.6151
R1120 B.n476 B.n475 10.6151
R1121 B.n477 B.n476 10.6151
R1122 B.n477 B.n154 10.6151
R1123 B.n487 B.n154 10.6151
R1124 B.n488 B.n487 10.6151
R1125 B.n489 B.n488 10.6151
R1126 B.n489 B.n146 10.6151
R1127 B.n499 B.n146 10.6151
R1128 B.n500 B.n499 10.6151
R1129 B.n501 B.n500 10.6151
R1130 B.n501 B.n138 10.6151
R1131 B.n511 B.n138 10.6151
R1132 B.n512 B.n511 10.6151
R1133 B.n513 B.n512 10.6151
R1134 B.n513 B.n130 10.6151
R1135 B.n523 B.n130 10.6151
R1136 B.n524 B.n523 10.6151
R1137 B.n525 B.n524 10.6151
R1138 B.n525 B.n122 10.6151
R1139 B.n536 B.n122 10.6151
R1140 B.n537 B.n536 10.6151
R1141 B.n538 B.n537 10.6151
R1142 B.n538 B.n0 10.6151
R1143 B.n451 B.n450 10.6151
R1144 B.n450 B.n177 10.6151
R1145 B.n445 B.n177 10.6151
R1146 B.n445 B.n444 10.6151
R1147 B.n444 B.n179 10.6151
R1148 B.n439 B.n179 10.6151
R1149 B.n439 B.n438 10.6151
R1150 B.n438 B.n437 10.6151
R1151 B.n437 B.n181 10.6151
R1152 B.n431 B.n181 10.6151
R1153 B.n431 B.n430 10.6151
R1154 B.n430 B.n429 10.6151
R1155 B.n429 B.n183 10.6151
R1156 B.n423 B.n183 10.6151
R1157 B.n423 B.n422 10.6151
R1158 B.n422 B.n421 10.6151
R1159 B.n421 B.n185 10.6151
R1160 B.n415 B.n185 10.6151
R1161 B.n415 B.n414 10.6151
R1162 B.n414 B.n413 10.6151
R1163 B.n413 B.n187 10.6151
R1164 B.n407 B.n187 10.6151
R1165 B.n407 B.n406 10.6151
R1166 B.n406 B.n405 10.6151
R1167 B.n405 B.n189 10.6151
R1168 B.n399 B.n189 10.6151
R1169 B.n399 B.n398 10.6151
R1170 B.n398 B.n397 10.6151
R1171 B.n397 B.n191 10.6151
R1172 B.n391 B.n191 10.6151
R1173 B.n391 B.n390 10.6151
R1174 B.n390 B.n389 10.6151
R1175 B.n389 B.n193 10.6151
R1176 B.n383 B.n193 10.6151
R1177 B.n383 B.n382 10.6151
R1178 B.n382 B.n381 10.6151
R1179 B.n381 B.n195 10.6151
R1180 B.n375 B.n195 10.6151
R1181 B.n375 B.n374 10.6151
R1182 B.n374 B.n373 10.6151
R1183 B.n373 B.n197 10.6151
R1184 B.n367 B.n197 10.6151
R1185 B.n367 B.n366 10.6151
R1186 B.n366 B.n365 10.6151
R1187 B.n365 B.n199 10.6151
R1188 B.n359 B.n199 10.6151
R1189 B.n359 B.n358 10.6151
R1190 B.n358 B.n357 10.6151
R1191 B.n357 B.n201 10.6151
R1192 B.n351 B.n350 10.6151
R1193 B.n350 B.n349 10.6151
R1194 B.n349 B.n206 10.6151
R1195 B.n343 B.n206 10.6151
R1196 B.n343 B.n342 10.6151
R1197 B.n342 B.n341 10.6151
R1198 B.n341 B.n208 10.6151
R1199 B.n335 B.n208 10.6151
R1200 B.n333 B.n332 10.6151
R1201 B.n332 B.n212 10.6151
R1202 B.n326 B.n212 10.6151
R1203 B.n326 B.n325 10.6151
R1204 B.n325 B.n324 10.6151
R1205 B.n324 B.n214 10.6151
R1206 B.n318 B.n214 10.6151
R1207 B.n318 B.n317 10.6151
R1208 B.n317 B.n316 10.6151
R1209 B.n316 B.n216 10.6151
R1210 B.n310 B.n216 10.6151
R1211 B.n310 B.n309 10.6151
R1212 B.n309 B.n308 10.6151
R1213 B.n308 B.n218 10.6151
R1214 B.n302 B.n218 10.6151
R1215 B.n302 B.n301 10.6151
R1216 B.n301 B.n300 10.6151
R1217 B.n300 B.n220 10.6151
R1218 B.n294 B.n220 10.6151
R1219 B.n294 B.n293 10.6151
R1220 B.n293 B.n292 10.6151
R1221 B.n292 B.n222 10.6151
R1222 B.n286 B.n222 10.6151
R1223 B.n286 B.n285 10.6151
R1224 B.n285 B.n284 10.6151
R1225 B.n284 B.n224 10.6151
R1226 B.n278 B.n224 10.6151
R1227 B.n278 B.n277 10.6151
R1228 B.n277 B.n276 10.6151
R1229 B.n276 B.n226 10.6151
R1230 B.n270 B.n226 10.6151
R1231 B.n270 B.n269 10.6151
R1232 B.n269 B.n268 10.6151
R1233 B.n268 B.n228 10.6151
R1234 B.n262 B.n228 10.6151
R1235 B.n262 B.n261 10.6151
R1236 B.n261 B.n260 10.6151
R1237 B.n260 B.n230 10.6151
R1238 B.n254 B.n230 10.6151
R1239 B.n254 B.n253 10.6151
R1240 B.n253 B.n252 10.6151
R1241 B.n252 B.n232 10.6151
R1242 B.n246 B.n232 10.6151
R1243 B.n246 B.n245 10.6151
R1244 B.n245 B.n244 10.6151
R1245 B.n244 B.n234 10.6151
R1246 B.n238 B.n234 10.6151
R1247 B.n238 B.n237 10.6151
R1248 B.n237 B.n173 10.6151
R1249 B.n457 B.n456 10.6151
R1250 B.n458 B.n457 10.6151
R1251 B.n458 B.n165 10.6151
R1252 B.n468 B.n165 10.6151
R1253 B.n469 B.n468 10.6151
R1254 B.n470 B.n469 10.6151
R1255 B.n470 B.n158 10.6151
R1256 B.n481 B.n158 10.6151
R1257 B.n482 B.n481 10.6151
R1258 B.n483 B.n482 10.6151
R1259 B.n483 B.n150 10.6151
R1260 B.n493 B.n150 10.6151
R1261 B.n494 B.n493 10.6151
R1262 B.n495 B.n494 10.6151
R1263 B.n495 B.n141 10.6151
R1264 B.n505 B.n141 10.6151
R1265 B.n506 B.n505 10.6151
R1266 B.n507 B.n506 10.6151
R1267 B.n507 B.n134 10.6151
R1268 B.n517 B.n134 10.6151
R1269 B.n518 B.n517 10.6151
R1270 B.n519 B.n518 10.6151
R1271 B.n519 B.n125 10.6151
R1272 B.n529 B.n125 10.6151
R1273 B.n530 B.n529 10.6151
R1274 B.n532 B.n530 10.6151
R1275 B.n532 B.n531 10.6151
R1276 B.n531 B.n118 10.6151
R1277 B.n543 B.n118 10.6151
R1278 B.n544 B.n543 10.6151
R1279 B.n545 B.n544 10.6151
R1280 B.n546 B.n545 10.6151
R1281 B.n547 B.n546 10.6151
R1282 B.n550 B.n547 10.6151
R1283 B.n551 B.n550 10.6151
R1284 B.n552 B.n551 10.6151
R1285 B.n553 B.n552 10.6151
R1286 B.n555 B.n553 10.6151
R1287 B.n556 B.n555 10.6151
R1288 B.n557 B.n556 10.6151
R1289 B.n558 B.n557 10.6151
R1290 B.n560 B.n558 10.6151
R1291 B.n561 B.n560 10.6151
R1292 B.n562 B.n561 10.6151
R1293 B.n563 B.n562 10.6151
R1294 B.n565 B.n563 10.6151
R1295 B.n566 B.n565 10.6151
R1296 B.n567 B.n566 10.6151
R1297 B.n568 B.n567 10.6151
R1298 B.n570 B.n568 10.6151
R1299 B.n571 B.n570 10.6151
R1300 B.n572 B.n571 10.6151
R1301 B.n573 B.n572 10.6151
R1302 B.n575 B.n573 10.6151
R1303 B.n576 B.n575 10.6151
R1304 B.n577 B.n576 10.6151
R1305 B.n578 B.n577 10.6151
R1306 B.n580 B.n578 10.6151
R1307 B.n581 B.n580 10.6151
R1308 B.n582 B.n581 10.6151
R1309 B.n583 B.n582 10.6151
R1310 B.n859 B.n1 10.6151
R1311 B.n859 B.n858 10.6151
R1312 B.n858 B.n857 10.6151
R1313 B.n857 B.n10 10.6151
R1314 B.n851 B.n10 10.6151
R1315 B.n851 B.n850 10.6151
R1316 B.n850 B.n849 10.6151
R1317 B.n849 B.n18 10.6151
R1318 B.n843 B.n18 10.6151
R1319 B.n843 B.n842 10.6151
R1320 B.n842 B.n841 10.6151
R1321 B.n841 B.n25 10.6151
R1322 B.n835 B.n25 10.6151
R1323 B.n835 B.n834 10.6151
R1324 B.n834 B.n833 10.6151
R1325 B.n833 B.n32 10.6151
R1326 B.n827 B.n32 10.6151
R1327 B.n827 B.n826 10.6151
R1328 B.n826 B.n825 10.6151
R1329 B.n825 B.n39 10.6151
R1330 B.n819 B.n39 10.6151
R1331 B.n819 B.n818 10.6151
R1332 B.n818 B.n817 10.6151
R1333 B.n817 B.n45 10.6151
R1334 B.n811 B.n45 10.6151
R1335 B.n811 B.n810 10.6151
R1336 B.n810 B.n809 10.6151
R1337 B.n809 B.n53 10.6151
R1338 B.n803 B.n53 10.6151
R1339 B.n802 B.n801 10.6151
R1340 B.n801 B.n60 10.6151
R1341 B.n795 B.n60 10.6151
R1342 B.n795 B.n794 10.6151
R1343 B.n794 B.n793 10.6151
R1344 B.n793 B.n62 10.6151
R1345 B.n787 B.n62 10.6151
R1346 B.n787 B.n786 10.6151
R1347 B.n786 B.n785 10.6151
R1348 B.n785 B.n64 10.6151
R1349 B.n779 B.n64 10.6151
R1350 B.n779 B.n778 10.6151
R1351 B.n778 B.n777 10.6151
R1352 B.n777 B.n66 10.6151
R1353 B.n771 B.n66 10.6151
R1354 B.n771 B.n770 10.6151
R1355 B.n770 B.n769 10.6151
R1356 B.n769 B.n68 10.6151
R1357 B.n763 B.n68 10.6151
R1358 B.n763 B.n762 10.6151
R1359 B.n762 B.n761 10.6151
R1360 B.n761 B.n70 10.6151
R1361 B.n755 B.n70 10.6151
R1362 B.n755 B.n754 10.6151
R1363 B.n754 B.n753 10.6151
R1364 B.n753 B.n72 10.6151
R1365 B.n747 B.n72 10.6151
R1366 B.n747 B.n746 10.6151
R1367 B.n746 B.n745 10.6151
R1368 B.n745 B.n74 10.6151
R1369 B.n739 B.n74 10.6151
R1370 B.n739 B.n738 10.6151
R1371 B.n738 B.n737 10.6151
R1372 B.n737 B.n76 10.6151
R1373 B.n731 B.n76 10.6151
R1374 B.n731 B.n730 10.6151
R1375 B.n730 B.n729 10.6151
R1376 B.n729 B.n78 10.6151
R1377 B.n723 B.n78 10.6151
R1378 B.n723 B.n722 10.6151
R1379 B.n722 B.n721 10.6151
R1380 B.n721 B.n80 10.6151
R1381 B.n715 B.n80 10.6151
R1382 B.n715 B.n714 10.6151
R1383 B.n714 B.n713 10.6151
R1384 B.n713 B.n82 10.6151
R1385 B.n707 B.n82 10.6151
R1386 B.n707 B.n706 10.6151
R1387 B.n706 B.n705 10.6151
R1388 B.n701 B.n700 10.6151
R1389 B.n700 B.n88 10.6151
R1390 B.n695 B.n88 10.6151
R1391 B.n695 B.n694 10.6151
R1392 B.n694 B.n693 10.6151
R1393 B.n693 B.n90 10.6151
R1394 B.n687 B.n90 10.6151
R1395 B.n687 B.n686 10.6151
R1396 B.n684 B.n94 10.6151
R1397 B.n678 B.n94 10.6151
R1398 B.n678 B.n677 10.6151
R1399 B.n677 B.n676 10.6151
R1400 B.n676 B.n96 10.6151
R1401 B.n670 B.n96 10.6151
R1402 B.n670 B.n669 10.6151
R1403 B.n669 B.n668 10.6151
R1404 B.n668 B.n98 10.6151
R1405 B.n662 B.n98 10.6151
R1406 B.n662 B.n661 10.6151
R1407 B.n661 B.n660 10.6151
R1408 B.n660 B.n100 10.6151
R1409 B.n654 B.n100 10.6151
R1410 B.n654 B.n653 10.6151
R1411 B.n653 B.n652 10.6151
R1412 B.n652 B.n102 10.6151
R1413 B.n646 B.n102 10.6151
R1414 B.n646 B.n645 10.6151
R1415 B.n645 B.n644 10.6151
R1416 B.n644 B.n104 10.6151
R1417 B.n638 B.n104 10.6151
R1418 B.n638 B.n637 10.6151
R1419 B.n637 B.n636 10.6151
R1420 B.n636 B.n106 10.6151
R1421 B.n630 B.n106 10.6151
R1422 B.n630 B.n629 10.6151
R1423 B.n629 B.n628 10.6151
R1424 B.n628 B.n108 10.6151
R1425 B.n622 B.n108 10.6151
R1426 B.n622 B.n621 10.6151
R1427 B.n621 B.n620 10.6151
R1428 B.n620 B.n110 10.6151
R1429 B.n614 B.n110 10.6151
R1430 B.n614 B.n613 10.6151
R1431 B.n613 B.n612 10.6151
R1432 B.n612 B.n112 10.6151
R1433 B.n606 B.n112 10.6151
R1434 B.n606 B.n605 10.6151
R1435 B.n605 B.n604 10.6151
R1436 B.n604 B.n114 10.6151
R1437 B.n598 B.n114 10.6151
R1438 B.n598 B.n597 10.6151
R1439 B.n597 B.n596 10.6151
R1440 B.n596 B.n116 10.6151
R1441 B.n590 B.n116 10.6151
R1442 B.n590 B.n589 10.6151
R1443 B.n589 B.n588 10.6151
R1444 B.n588 B.n584 10.6151
R1445 B.n509 B.t0 8.25256
R1446 B.n839 B.t2 8.25256
R1447 B.n867 B.n0 8.11757
R1448 B.n867 B.n1 8.11757
R1449 B.n128 B.t1 7.15229
R1450 B.t3 B.n854 7.15229
R1451 B.n351 B.n205 6.5566
R1452 B.n335 B.n334 6.5566
R1453 B.n701 B.n86 6.5566
R1454 B.n686 B.n685 6.5566
R1455 B.n472 B.t5 6.05201
R1456 B.n47 B.t12 6.05201
R1457 B.n205 B.n201 4.05904
R1458 B.n334 B.n333 4.05904
R1459 B.n705 B.n86 4.05904
R1460 B.n685 B.n684 4.05904
R1461 VP.n3 VP.t3 197.677
R1462 VP.n3 VP.t0 197.042
R1463 VP.n5 VP.t2 161.988
R1464 VP.n13 VP.t1 161.988
R1465 VP.n12 VP.n0 161.3
R1466 VP.n11 VP.n10 161.3
R1467 VP.n9 VP.n1 161.3
R1468 VP.n8 VP.n7 161.3
R1469 VP.n6 VP.n2 161.3
R1470 VP.n5 VP.n4 98.1205
R1471 VP.n14 VP.n13 98.1205
R1472 VP.n4 VP.n3 52.8813
R1473 VP.n7 VP.n1 40.577
R1474 VP.n11 VP.n1 40.577
R1475 VP.n7 VP.n6 24.5923
R1476 VP.n12 VP.n11 24.5923
R1477 VP.n6 VP.n5 12.7883
R1478 VP.n13 VP.n12 12.7883
R1479 VP.n4 VP.n2 0.278335
R1480 VP.n14 VP.n0 0.278335
R1481 VP.n8 VP.n2 0.189894
R1482 VP.n9 VP.n8 0.189894
R1483 VP.n10 VP.n9 0.189894
R1484 VP.n10 VP.n0 0.189894
R1485 VP VP.n14 0.153485
R1486 VTAIL.n650 VTAIL.n574 289.615
R1487 VTAIL.n76 VTAIL.n0 289.615
R1488 VTAIL.n158 VTAIL.n82 289.615
R1489 VTAIL.n240 VTAIL.n164 289.615
R1490 VTAIL.n568 VTAIL.n492 289.615
R1491 VTAIL.n486 VTAIL.n410 289.615
R1492 VTAIL.n404 VTAIL.n328 289.615
R1493 VTAIL.n322 VTAIL.n246 289.615
R1494 VTAIL.n601 VTAIL.n600 185
R1495 VTAIL.n598 VTAIL.n597 185
R1496 VTAIL.n607 VTAIL.n606 185
R1497 VTAIL.n609 VTAIL.n608 185
R1498 VTAIL.n594 VTAIL.n593 185
R1499 VTAIL.n615 VTAIL.n614 185
R1500 VTAIL.n617 VTAIL.n616 185
R1501 VTAIL.n590 VTAIL.n589 185
R1502 VTAIL.n623 VTAIL.n622 185
R1503 VTAIL.n625 VTAIL.n624 185
R1504 VTAIL.n586 VTAIL.n585 185
R1505 VTAIL.n631 VTAIL.n630 185
R1506 VTAIL.n633 VTAIL.n632 185
R1507 VTAIL.n582 VTAIL.n581 185
R1508 VTAIL.n639 VTAIL.n638 185
R1509 VTAIL.n642 VTAIL.n641 185
R1510 VTAIL.n640 VTAIL.n578 185
R1511 VTAIL.n647 VTAIL.n577 185
R1512 VTAIL.n649 VTAIL.n648 185
R1513 VTAIL.n651 VTAIL.n650 185
R1514 VTAIL.n27 VTAIL.n26 185
R1515 VTAIL.n24 VTAIL.n23 185
R1516 VTAIL.n33 VTAIL.n32 185
R1517 VTAIL.n35 VTAIL.n34 185
R1518 VTAIL.n20 VTAIL.n19 185
R1519 VTAIL.n41 VTAIL.n40 185
R1520 VTAIL.n43 VTAIL.n42 185
R1521 VTAIL.n16 VTAIL.n15 185
R1522 VTAIL.n49 VTAIL.n48 185
R1523 VTAIL.n51 VTAIL.n50 185
R1524 VTAIL.n12 VTAIL.n11 185
R1525 VTAIL.n57 VTAIL.n56 185
R1526 VTAIL.n59 VTAIL.n58 185
R1527 VTAIL.n8 VTAIL.n7 185
R1528 VTAIL.n65 VTAIL.n64 185
R1529 VTAIL.n68 VTAIL.n67 185
R1530 VTAIL.n66 VTAIL.n4 185
R1531 VTAIL.n73 VTAIL.n3 185
R1532 VTAIL.n75 VTAIL.n74 185
R1533 VTAIL.n77 VTAIL.n76 185
R1534 VTAIL.n109 VTAIL.n108 185
R1535 VTAIL.n106 VTAIL.n105 185
R1536 VTAIL.n115 VTAIL.n114 185
R1537 VTAIL.n117 VTAIL.n116 185
R1538 VTAIL.n102 VTAIL.n101 185
R1539 VTAIL.n123 VTAIL.n122 185
R1540 VTAIL.n125 VTAIL.n124 185
R1541 VTAIL.n98 VTAIL.n97 185
R1542 VTAIL.n131 VTAIL.n130 185
R1543 VTAIL.n133 VTAIL.n132 185
R1544 VTAIL.n94 VTAIL.n93 185
R1545 VTAIL.n139 VTAIL.n138 185
R1546 VTAIL.n141 VTAIL.n140 185
R1547 VTAIL.n90 VTAIL.n89 185
R1548 VTAIL.n147 VTAIL.n146 185
R1549 VTAIL.n150 VTAIL.n149 185
R1550 VTAIL.n148 VTAIL.n86 185
R1551 VTAIL.n155 VTAIL.n85 185
R1552 VTAIL.n157 VTAIL.n156 185
R1553 VTAIL.n159 VTAIL.n158 185
R1554 VTAIL.n191 VTAIL.n190 185
R1555 VTAIL.n188 VTAIL.n187 185
R1556 VTAIL.n197 VTAIL.n196 185
R1557 VTAIL.n199 VTAIL.n198 185
R1558 VTAIL.n184 VTAIL.n183 185
R1559 VTAIL.n205 VTAIL.n204 185
R1560 VTAIL.n207 VTAIL.n206 185
R1561 VTAIL.n180 VTAIL.n179 185
R1562 VTAIL.n213 VTAIL.n212 185
R1563 VTAIL.n215 VTAIL.n214 185
R1564 VTAIL.n176 VTAIL.n175 185
R1565 VTAIL.n221 VTAIL.n220 185
R1566 VTAIL.n223 VTAIL.n222 185
R1567 VTAIL.n172 VTAIL.n171 185
R1568 VTAIL.n229 VTAIL.n228 185
R1569 VTAIL.n232 VTAIL.n231 185
R1570 VTAIL.n230 VTAIL.n168 185
R1571 VTAIL.n237 VTAIL.n167 185
R1572 VTAIL.n239 VTAIL.n238 185
R1573 VTAIL.n241 VTAIL.n240 185
R1574 VTAIL.n569 VTAIL.n568 185
R1575 VTAIL.n567 VTAIL.n566 185
R1576 VTAIL.n565 VTAIL.n495 185
R1577 VTAIL.n499 VTAIL.n496 185
R1578 VTAIL.n560 VTAIL.n559 185
R1579 VTAIL.n558 VTAIL.n557 185
R1580 VTAIL.n501 VTAIL.n500 185
R1581 VTAIL.n552 VTAIL.n551 185
R1582 VTAIL.n550 VTAIL.n549 185
R1583 VTAIL.n505 VTAIL.n504 185
R1584 VTAIL.n544 VTAIL.n543 185
R1585 VTAIL.n542 VTAIL.n541 185
R1586 VTAIL.n509 VTAIL.n508 185
R1587 VTAIL.n536 VTAIL.n535 185
R1588 VTAIL.n534 VTAIL.n533 185
R1589 VTAIL.n513 VTAIL.n512 185
R1590 VTAIL.n528 VTAIL.n527 185
R1591 VTAIL.n526 VTAIL.n525 185
R1592 VTAIL.n517 VTAIL.n516 185
R1593 VTAIL.n520 VTAIL.n519 185
R1594 VTAIL.n487 VTAIL.n486 185
R1595 VTAIL.n485 VTAIL.n484 185
R1596 VTAIL.n483 VTAIL.n413 185
R1597 VTAIL.n417 VTAIL.n414 185
R1598 VTAIL.n478 VTAIL.n477 185
R1599 VTAIL.n476 VTAIL.n475 185
R1600 VTAIL.n419 VTAIL.n418 185
R1601 VTAIL.n470 VTAIL.n469 185
R1602 VTAIL.n468 VTAIL.n467 185
R1603 VTAIL.n423 VTAIL.n422 185
R1604 VTAIL.n462 VTAIL.n461 185
R1605 VTAIL.n460 VTAIL.n459 185
R1606 VTAIL.n427 VTAIL.n426 185
R1607 VTAIL.n454 VTAIL.n453 185
R1608 VTAIL.n452 VTAIL.n451 185
R1609 VTAIL.n431 VTAIL.n430 185
R1610 VTAIL.n446 VTAIL.n445 185
R1611 VTAIL.n444 VTAIL.n443 185
R1612 VTAIL.n435 VTAIL.n434 185
R1613 VTAIL.n438 VTAIL.n437 185
R1614 VTAIL.n405 VTAIL.n404 185
R1615 VTAIL.n403 VTAIL.n402 185
R1616 VTAIL.n401 VTAIL.n331 185
R1617 VTAIL.n335 VTAIL.n332 185
R1618 VTAIL.n396 VTAIL.n395 185
R1619 VTAIL.n394 VTAIL.n393 185
R1620 VTAIL.n337 VTAIL.n336 185
R1621 VTAIL.n388 VTAIL.n387 185
R1622 VTAIL.n386 VTAIL.n385 185
R1623 VTAIL.n341 VTAIL.n340 185
R1624 VTAIL.n380 VTAIL.n379 185
R1625 VTAIL.n378 VTAIL.n377 185
R1626 VTAIL.n345 VTAIL.n344 185
R1627 VTAIL.n372 VTAIL.n371 185
R1628 VTAIL.n370 VTAIL.n369 185
R1629 VTAIL.n349 VTAIL.n348 185
R1630 VTAIL.n364 VTAIL.n363 185
R1631 VTAIL.n362 VTAIL.n361 185
R1632 VTAIL.n353 VTAIL.n352 185
R1633 VTAIL.n356 VTAIL.n355 185
R1634 VTAIL.n323 VTAIL.n322 185
R1635 VTAIL.n321 VTAIL.n320 185
R1636 VTAIL.n319 VTAIL.n249 185
R1637 VTAIL.n253 VTAIL.n250 185
R1638 VTAIL.n314 VTAIL.n313 185
R1639 VTAIL.n312 VTAIL.n311 185
R1640 VTAIL.n255 VTAIL.n254 185
R1641 VTAIL.n306 VTAIL.n305 185
R1642 VTAIL.n304 VTAIL.n303 185
R1643 VTAIL.n259 VTAIL.n258 185
R1644 VTAIL.n298 VTAIL.n297 185
R1645 VTAIL.n296 VTAIL.n295 185
R1646 VTAIL.n263 VTAIL.n262 185
R1647 VTAIL.n290 VTAIL.n289 185
R1648 VTAIL.n288 VTAIL.n287 185
R1649 VTAIL.n267 VTAIL.n266 185
R1650 VTAIL.n282 VTAIL.n281 185
R1651 VTAIL.n280 VTAIL.n279 185
R1652 VTAIL.n271 VTAIL.n270 185
R1653 VTAIL.n274 VTAIL.n273 185
R1654 VTAIL.t7 VTAIL.n518 147.659
R1655 VTAIL.t6 VTAIL.n436 147.659
R1656 VTAIL.t3 VTAIL.n354 147.659
R1657 VTAIL.t2 VTAIL.n272 147.659
R1658 VTAIL.t1 VTAIL.n599 147.659
R1659 VTAIL.t0 VTAIL.n25 147.659
R1660 VTAIL.t5 VTAIL.n107 147.659
R1661 VTAIL.t4 VTAIL.n189 147.659
R1662 VTAIL.n600 VTAIL.n597 104.615
R1663 VTAIL.n607 VTAIL.n597 104.615
R1664 VTAIL.n608 VTAIL.n607 104.615
R1665 VTAIL.n608 VTAIL.n593 104.615
R1666 VTAIL.n615 VTAIL.n593 104.615
R1667 VTAIL.n616 VTAIL.n615 104.615
R1668 VTAIL.n616 VTAIL.n589 104.615
R1669 VTAIL.n623 VTAIL.n589 104.615
R1670 VTAIL.n624 VTAIL.n623 104.615
R1671 VTAIL.n624 VTAIL.n585 104.615
R1672 VTAIL.n631 VTAIL.n585 104.615
R1673 VTAIL.n632 VTAIL.n631 104.615
R1674 VTAIL.n632 VTAIL.n581 104.615
R1675 VTAIL.n639 VTAIL.n581 104.615
R1676 VTAIL.n641 VTAIL.n639 104.615
R1677 VTAIL.n641 VTAIL.n640 104.615
R1678 VTAIL.n640 VTAIL.n577 104.615
R1679 VTAIL.n649 VTAIL.n577 104.615
R1680 VTAIL.n650 VTAIL.n649 104.615
R1681 VTAIL.n26 VTAIL.n23 104.615
R1682 VTAIL.n33 VTAIL.n23 104.615
R1683 VTAIL.n34 VTAIL.n33 104.615
R1684 VTAIL.n34 VTAIL.n19 104.615
R1685 VTAIL.n41 VTAIL.n19 104.615
R1686 VTAIL.n42 VTAIL.n41 104.615
R1687 VTAIL.n42 VTAIL.n15 104.615
R1688 VTAIL.n49 VTAIL.n15 104.615
R1689 VTAIL.n50 VTAIL.n49 104.615
R1690 VTAIL.n50 VTAIL.n11 104.615
R1691 VTAIL.n57 VTAIL.n11 104.615
R1692 VTAIL.n58 VTAIL.n57 104.615
R1693 VTAIL.n58 VTAIL.n7 104.615
R1694 VTAIL.n65 VTAIL.n7 104.615
R1695 VTAIL.n67 VTAIL.n65 104.615
R1696 VTAIL.n67 VTAIL.n66 104.615
R1697 VTAIL.n66 VTAIL.n3 104.615
R1698 VTAIL.n75 VTAIL.n3 104.615
R1699 VTAIL.n76 VTAIL.n75 104.615
R1700 VTAIL.n108 VTAIL.n105 104.615
R1701 VTAIL.n115 VTAIL.n105 104.615
R1702 VTAIL.n116 VTAIL.n115 104.615
R1703 VTAIL.n116 VTAIL.n101 104.615
R1704 VTAIL.n123 VTAIL.n101 104.615
R1705 VTAIL.n124 VTAIL.n123 104.615
R1706 VTAIL.n124 VTAIL.n97 104.615
R1707 VTAIL.n131 VTAIL.n97 104.615
R1708 VTAIL.n132 VTAIL.n131 104.615
R1709 VTAIL.n132 VTAIL.n93 104.615
R1710 VTAIL.n139 VTAIL.n93 104.615
R1711 VTAIL.n140 VTAIL.n139 104.615
R1712 VTAIL.n140 VTAIL.n89 104.615
R1713 VTAIL.n147 VTAIL.n89 104.615
R1714 VTAIL.n149 VTAIL.n147 104.615
R1715 VTAIL.n149 VTAIL.n148 104.615
R1716 VTAIL.n148 VTAIL.n85 104.615
R1717 VTAIL.n157 VTAIL.n85 104.615
R1718 VTAIL.n158 VTAIL.n157 104.615
R1719 VTAIL.n190 VTAIL.n187 104.615
R1720 VTAIL.n197 VTAIL.n187 104.615
R1721 VTAIL.n198 VTAIL.n197 104.615
R1722 VTAIL.n198 VTAIL.n183 104.615
R1723 VTAIL.n205 VTAIL.n183 104.615
R1724 VTAIL.n206 VTAIL.n205 104.615
R1725 VTAIL.n206 VTAIL.n179 104.615
R1726 VTAIL.n213 VTAIL.n179 104.615
R1727 VTAIL.n214 VTAIL.n213 104.615
R1728 VTAIL.n214 VTAIL.n175 104.615
R1729 VTAIL.n221 VTAIL.n175 104.615
R1730 VTAIL.n222 VTAIL.n221 104.615
R1731 VTAIL.n222 VTAIL.n171 104.615
R1732 VTAIL.n229 VTAIL.n171 104.615
R1733 VTAIL.n231 VTAIL.n229 104.615
R1734 VTAIL.n231 VTAIL.n230 104.615
R1735 VTAIL.n230 VTAIL.n167 104.615
R1736 VTAIL.n239 VTAIL.n167 104.615
R1737 VTAIL.n240 VTAIL.n239 104.615
R1738 VTAIL.n568 VTAIL.n567 104.615
R1739 VTAIL.n567 VTAIL.n495 104.615
R1740 VTAIL.n499 VTAIL.n495 104.615
R1741 VTAIL.n559 VTAIL.n499 104.615
R1742 VTAIL.n559 VTAIL.n558 104.615
R1743 VTAIL.n558 VTAIL.n500 104.615
R1744 VTAIL.n551 VTAIL.n500 104.615
R1745 VTAIL.n551 VTAIL.n550 104.615
R1746 VTAIL.n550 VTAIL.n504 104.615
R1747 VTAIL.n543 VTAIL.n504 104.615
R1748 VTAIL.n543 VTAIL.n542 104.615
R1749 VTAIL.n542 VTAIL.n508 104.615
R1750 VTAIL.n535 VTAIL.n508 104.615
R1751 VTAIL.n535 VTAIL.n534 104.615
R1752 VTAIL.n534 VTAIL.n512 104.615
R1753 VTAIL.n527 VTAIL.n512 104.615
R1754 VTAIL.n527 VTAIL.n526 104.615
R1755 VTAIL.n526 VTAIL.n516 104.615
R1756 VTAIL.n519 VTAIL.n516 104.615
R1757 VTAIL.n486 VTAIL.n485 104.615
R1758 VTAIL.n485 VTAIL.n413 104.615
R1759 VTAIL.n417 VTAIL.n413 104.615
R1760 VTAIL.n477 VTAIL.n417 104.615
R1761 VTAIL.n477 VTAIL.n476 104.615
R1762 VTAIL.n476 VTAIL.n418 104.615
R1763 VTAIL.n469 VTAIL.n418 104.615
R1764 VTAIL.n469 VTAIL.n468 104.615
R1765 VTAIL.n468 VTAIL.n422 104.615
R1766 VTAIL.n461 VTAIL.n422 104.615
R1767 VTAIL.n461 VTAIL.n460 104.615
R1768 VTAIL.n460 VTAIL.n426 104.615
R1769 VTAIL.n453 VTAIL.n426 104.615
R1770 VTAIL.n453 VTAIL.n452 104.615
R1771 VTAIL.n452 VTAIL.n430 104.615
R1772 VTAIL.n445 VTAIL.n430 104.615
R1773 VTAIL.n445 VTAIL.n444 104.615
R1774 VTAIL.n444 VTAIL.n434 104.615
R1775 VTAIL.n437 VTAIL.n434 104.615
R1776 VTAIL.n404 VTAIL.n403 104.615
R1777 VTAIL.n403 VTAIL.n331 104.615
R1778 VTAIL.n335 VTAIL.n331 104.615
R1779 VTAIL.n395 VTAIL.n335 104.615
R1780 VTAIL.n395 VTAIL.n394 104.615
R1781 VTAIL.n394 VTAIL.n336 104.615
R1782 VTAIL.n387 VTAIL.n336 104.615
R1783 VTAIL.n387 VTAIL.n386 104.615
R1784 VTAIL.n386 VTAIL.n340 104.615
R1785 VTAIL.n379 VTAIL.n340 104.615
R1786 VTAIL.n379 VTAIL.n378 104.615
R1787 VTAIL.n378 VTAIL.n344 104.615
R1788 VTAIL.n371 VTAIL.n344 104.615
R1789 VTAIL.n371 VTAIL.n370 104.615
R1790 VTAIL.n370 VTAIL.n348 104.615
R1791 VTAIL.n363 VTAIL.n348 104.615
R1792 VTAIL.n363 VTAIL.n362 104.615
R1793 VTAIL.n362 VTAIL.n352 104.615
R1794 VTAIL.n355 VTAIL.n352 104.615
R1795 VTAIL.n322 VTAIL.n321 104.615
R1796 VTAIL.n321 VTAIL.n249 104.615
R1797 VTAIL.n253 VTAIL.n249 104.615
R1798 VTAIL.n313 VTAIL.n253 104.615
R1799 VTAIL.n313 VTAIL.n312 104.615
R1800 VTAIL.n312 VTAIL.n254 104.615
R1801 VTAIL.n305 VTAIL.n254 104.615
R1802 VTAIL.n305 VTAIL.n304 104.615
R1803 VTAIL.n304 VTAIL.n258 104.615
R1804 VTAIL.n297 VTAIL.n258 104.615
R1805 VTAIL.n297 VTAIL.n296 104.615
R1806 VTAIL.n296 VTAIL.n262 104.615
R1807 VTAIL.n289 VTAIL.n262 104.615
R1808 VTAIL.n289 VTAIL.n288 104.615
R1809 VTAIL.n288 VTAIL.n266 104.615
R1810 VTAIL.n281 VTAIL.n266 104.615
R1811 VTAIL.n281 VTAIL.n280 104.615
R1812 VTAIL.n280 VTAIL.n270 104.615
R1813 VTAIL.n273 VTAIL.n270 104.615
R1814 VTAIL.n600 VTAIL.t1 52.3082
R1815 VTAIL.n26 VTAIL.t0 52.3082
R1816 VTAIL.n108 VTAIL.t5 52.3082
R1817 VTAIL.n190 VTAIL.t4 52.3082
R1818 VTAIL.n519 VTAIL.t7 52.3082
R1819 VTAIL.n437 VTAIL.t6 52.3082
R1820 VTAIL.n355 VTAIL.t3 52.3082
R1821 VTAIL.n273 VTAIL.t2 52.3082
R1822 VTAIL.n655 VTAIL.n654 33.7369
R1823 VTAIL.n81 VTAIL.n80 33.7369
R1824 VTAIL.n163 VTAIL.n162 33.7369
R1825 VTAIL.n245 VTAIL.n244 33.7369
R1826 VTAIL.n573 VTAIL.n572 33.7369
R1827 VTAIL.n491 VTAIL.n490 33.7369
R1828 VTAIL.n409 VTAIL.n408 33.7369
R1829 VTAIL.n327 VTAIL.n326 33.7369
R1830 VTAIL.n655 VTAIL.n573 27.2289
R1831 VTAIL.n327 VTAIL.n245 27.2289
R1832 VTAIL.n601 VTAIL.n599 15.6677
R1833 VTAIL.n27 VTAIL.n25 15.6677
R1834 VTAIL.n109 VTAIL.n107 15.6677
R1835 VTAIL.n191 VTAIL.n189 15.6677
R1836 VTAIL.n520 VTAIL.n518 15.6677
R1837 VTAIL.n438 VTAIL.n436 15.6677
R1838 VTAIL.n356 VTAIL.n354 15.6677
R1839 VTAIL.n274 VTAIL.n272 15.6677
R1840 VTAIL.n648 VTAIL.n647 13.1884
R1841 VTAIL.n74 VTAIL.n73 13.1884
R1842 VTAIL.n156 VTAIL.n155 13.1884
R1843 VTAIL.n238 VTAIL.n237 13.1884
R1844 VTAIL.n566 VTAIL.n565 13.1884
R1845 VTAIL.n484 VTAIL.n483 13.1884
R1846 VTAIL.n402 VTAIL.n401 13.1884
R1847 VTAIL.n320 VTAIL.n319 13.1884
R1848 VTAIL.n602 VTAIL.n598 12.8005
R1849 VTAIL.n646 VTAIL.n578 12.8005
R1850 VTAIL.n651 VTAIL.n576 12.8005
R1851 VTAIL.n28 VTAIL.n24 12.8005
R1852 VTAIL.n72 VTAIL.n4 12.8005
R1853 VTAIL.n77 VTAIL.n2 12.8005
R1854 VTAIL.n110 VTAIL.n106 12.8005
R1855 VTAIL.n154 VTAIL.n86 12.8005
R1856 VTAIL.n159 VTAIL.n84 12.8005
R1857 VTAIL.n192 VTAIL.n188 12.8005
R1858 VTAIL.n236 VTAIL.n168 12.8005
R1859 VTAIL.n241 VTAIL.n166 12.8005
R1860 VTAIL.n569 VTAIL.n494 12.8005
R1861 VTAIL.n564 VTAIL.n496 12.8005
R1862 VTAIL.n521 VTAIL.n517 12.8005
R1863 VTAIL.n487 VTAIL.n412 12.8005
R1864 VTAIL.n482 VTAIL.n414 12.8005
R1865 VTAIL.n439 VTAIL.n435 12.8005
R1866 VTAIL.n405 VTAIL.n330 12.8005
R1867 VTAIL.n400 VTAIL.n332 12.8005
R1868 VTAIL.n357 VTAIL.n353 12.8005
R1869 VTAIL.n323 VTAIL.n248 12.8005
R1870 VTAIL.n318 VTAIL.n250 12.8005
R1871 VTAIL.n275 VTAIL.n271 12.8005
R1872 VTAIL.n606 VTAIL.n605 12.0247
R1873 VTAIL.n643 VTAIL.n642 12.0247
R1874 VTAIL.n652 VTAIL.n574 12.0247
R1875 VTAIL.n32 VTAIL.n31 12.0247
R1876 VTAIL.n69 VTAIL.n68 12.0247
R1877 VTAIL.n78 VTAIL.n0 12.0247
R1878 VTAIL.n114 VTAIL.n113 12.0247
R1879 VTAIL.n151 VTAIL.n150 12.0247
R1880 VTAIL.n160 VTAIL.n82 12.0247
R1881 VTAIL.n196 VTAIL.n195 12.0247
R1882 VTAIL.n233 VTAIL.n232 12.0247
R1883 VTAIL.n242 VTAIL.n164 12.0247
R1884 VTAIL.n570 VTAIL.n492 12.0247
R1885 VTAIL.n561 VTAIL.n560 12.0247
R1886 VTAIL.n525 VTAIL.n524 12.0247
R1887 VTAIL.n488 VTAIL.n410 12.0247
R1888 VTAIL.n479 VTAIL.n478 12.0247
R1889 VTAIL.n443 VTAIL.n442 12.0247
R1890 VTAIL.n406 VTAIL.n328 12.0247
R1891 VTAIL.n397 VTAIL.n396 12.0247
R1892 VTAIL.n361 VTAIL.n360 12.0247
R1893 VTAIL.n324 VTAIL.n246 12.0247
R1894 VTAIL.n315 VTAIL.n314 12.0247
R1895 VTAIL.n279 VTAIL.n278 12.0247
R1896 VTAIL.n609 VTAIL.n596 11.249
R1897 VTAIL.n638 VTAIL.n580 11.249
R1898 VTAIL.n35 VTAIL.n22 11.249
R1899 VTAIL.n64 VTAIL.n6 11.249
R1900 VTAIL.n117 VTAIL.n104 11.249
R1901 VTAIL.n146 VTAIL.n88 11.249
R1902 VTAIL.n199 VTAIL.n186 11.249
R1903 VTAIL.n228 VTAIL.n170 11.249
R1904 VTAIL.n557 VTAIL.n498 11.249
R1905 VTAIL.n528 VTAIL.n515 11.249
R1906 VTAIL.n475 VTAIL.n416 11.249
R1907 VTAIL.n446 VTAIL.n433 11.249
R1908 VTAIL.n393 VTAIL.n334 11.249
R1909 VTAIL.n364 VTAIL.n351 11.249
R1910 VTAIL.n311 VTAIL.n252 11.249
R1911 VTAIL.n282 VTAIL.n269 11.249
R1912 VTAIL.n610 VTAIL.n594 10.4732
R1913 VTAIL.n637 VTAIL.n582 10.4732
R1914 VTAIL.n36 VTAIL.n20 10.4732
R1915 VTAIL.n63 VTAIL.n8 10.4732
R1916 VTAIL.n118 VTAIL.n102 10.4732
R1917 VTAIL.n145 VTAIL.n90 10.4732
R1918 VTAIL.n200 VTAIL.n184 10.4732
R1919 VTAIL.n227 VTAIL.n172 10.4732
R1920 VTAIL.n556 VTAIL.n501 10.4732
R1921 VTAIL.n529 VTAIL.n513 10.4732
R1922 VTAIL.n474 VTAIL.n419 10.4732
R1923 VTAIL.n447 VTAIL.n431 10.4732
R1924 VTAIL.n392 VTAIL.n337 10.4732
R1925 VTAIL.n365 VTAIL.n349 10.4732
R1926 VTAIL.n310 VTAIL.n255 10.4732
R1927 VTAIL.n283 VTAIL.n267 10.4732
R1928 VTAIL.n614 VTAIL.n613 9.69747
R1929 VTAIL.n634 VTAIL.n633 9.69747
R1930 VTAIL.n40 VTAIL.n39 9.69747
R1931 VTAIL.n60 VTAIL.n59 9.69747
R1932 VTAIL.n122 VTAIL.n121 9.69747
R1933 VTAIL.n142 VTAIL.n141 9.69747
R1934 VTAIL.n204 VTAIL.n203 9.69747
R1935 VTAIL.n224 VTAIL.n223 9.69747
R1936 VTAIL.n553 VTAIL.n552 9.69747
R1937 VTAIL.n533 VTAIL.n532 9.69747
R1938 VTAIL.n471 VTAIL.n470 9.69747
R1939 VTAIL.n451 VTAIL.n450 9.69747
R1940 VTAIL.n389 VTAIL.n388 9.69747
R1941 VTAIL.n369 VTAIL.n368 9.69747
R1942 VTAIL.n307 VTAIL.n306 9.69747
R1943 VTAIL.n287 VTAIL.n286 9.69747
R1944 VTAIL.n654 VTAIL.n653 9.45567
R1945 VTAIL.n80 VTAIL.n79 9.45567
R1946 VTAIL.n162 VTAIL.n161 9.45567
R1947 VTAIL.n244 VTAIL.n243 9.45567
R1948 VTAIL.n572 VTAIL.n571 9.45567
R1949 VTAIL.n490 VTAIL.n489 9.45567
R1950 VTAIL.n408 VTAIL.n407 9.45567
R1951 VTAIL.n326 VTAIL.n325 9.45567
R1952 VTAIL.n653 VTAIL.n652 9.3005
R1953 VTAIL.n576 VTAIL.n575 9.3005
R1954 VTAIL.n621 VTAIL.n620 9.3005
R1955 VTAIL.n619 VTAIL.n618 9.3005
R1956 VTAIL.n592 VTAIL.n591 9.3005
R1957 VTAIL.n613 VTAIL.n612 9.3005
R1958 VTAIL.n611 VTAIL.n610 9.3005
R1959 VTAIL.n596 VTAIL.n595 9.3005
R1960 VTAIL.n605 VTAIL.n604 9.3005
R1961 VTAIL.n603 VTAIL.n602 9.3005
R1962 VTAIL.n588 VTAIL.n587 9.3005
R1963 VTAIL.n627 VTAIL.n626 9.3005
R1964 VTAIL.n629 VTAIL.n628 9.3005
R1965 VTAIL.n584 VTAIL.n583 9.3005
R1966 VTAIL.n635 VTAIL.n634 9.3005
R1967 VTAIL.n637 VTAIL.n636 9.3005
R1968 VTAIL.n580 VTAIL.n579 9.3005
R1969 VTAIL.n644 VTAIL.n643 9.3005
R1970 VTAIL.n646 VTAIL.n645 9.3005
R1971 VTAIL.n79 VTAIL.n78 9.3005
R1972 VTAIL.n2 VTAIL.n1 9.3005
R1973 VTAIL.n47 VTAIL.n46 9.3005
R1974 VTAIL.n45 VTAIL.n44 9.3005
R1975 VTAIL.n18 VTAIL.n17 9.3005
R1976 VTAIL.n39 VTAIL.n38 9.3005
R1977 VTAIL.n37 VTAIL.n36 9.3005
R1978 VTAIL.n22 VTAIL.n21 9.3005
R1979 VTAIL.n31 VTAIL.n30 9.3005
R1980 VTAIL.n29 VTAIL.n28 9.3005
R1981 VTAIL.n14 VTAIL.n13 9.3005
R1982 VTAIL.n53 VTAIL.n52 9.3005
R1983 VTAIL.n55 VTAIL.n54 9.3005
R1984 VTAIL.n10 VTAIL.n9 9.3005
R1985 VTAIL.n61 VTAIL.n60 9.3005
R1986 VTAIL.n63 VTAIL.n62 9.3005
R1987 VTAIL.n6 VTAIL.n5 9.3005
R1988 VTAIL.n70 VTAIL.n69 9.3005
R1989 VTAIL.n72 VTAIL.n71 9.3005
R1990 VTAIL.n161 VTAIL.n160 9.3005
R1991 VTAIL.n84 VTAIL.n83 9.3005
R1992 VTAIL.n129 VTAIL.n128 9.3005
R1993 VTAIL.n127 VTAIL.n126 9.3005
R1994 VTAIL.n100 VTAIL.n99 9.3005
R1995 VTAIL.n121 VTAIL.n120 9.3005
R1996 VTAIL.n119 VTAIL.n118 9.3005
R1997 VTAIL.n104 VTAIL.n103 9.3005
R1998 VTAIL.n113 VTAIL.n112 9.3005
R1999 VTAIL.n111 VTAIL.n110 9.3005
R2000 VTAIL.n96 VTAIL.n95 9.3005
R2001 VTAIL.n135 VTAIL.n134 9.3005
R2002 VTAIL.n137 VTAIL.n136 9.3005
R2003 VTAIL.n92 VTAIL.n91 9.3005
R2004 VTAIL.n143 VTAIL.n142 9.3005
R2005 VTAIL.n145 VTAIL.n144 9.3005
R2006 VTAIL.n88 VTAIL.n87 9.3005
R2007 VTAIL.n152 VTAIL.n151 9.3005
R2008 VTAIL.n154 VTAIL.n153 9.3005
R2009 VTAIL.n243 VTAIL.n242 9.3005
R2010 VTAIL.n166 VTAIL.n165 9.3005
R2011 VTAIL.n211 VTAIL.n210 9.3005
R2012 VTAIL.n209 VTAIL.n208 9.3005
R2013 VTAIL.n182 VTAIL.n181 9.3005
R2014 VTAIL.n203 VTAIL.n202 9.3005
R2015 VTAIL.n201 VTAIL.n200 9.3005
R2016 VTAIL.n186 VTAIL.n185 9.3005
R2017 VTAIL.n195 VTAIL.n194 9.3005
R2018 VTAIL.n193 VTAIL.n192 9.3005
R2019 VTAIL.n178 VTAIL.n177 9.3005
R2020 VTAIL.n217 VTAIL.n216 9.3005
R2021 VTAIL.n219 VTAIL.n218 9.3005
R2022 VTAIL.n174 VTAIL.n173 9.3005
R2023 VTAIL.n225 VTAIL.n224 9.3005
R2024 VTAIL.n227 VTAIL.n226 9.3005
R2025 VTAIL.n170 VTAIL.n169 9.3005
R2026 VTAIL.n234 VTAIL.n233 9.3005
R2027 VTAIL.n236 VTAIL.n235 9.3005
R2028 VTAIL.n546 VTAIL.n545 9.3005
R2029 VTAIL.n548 VTAIL.n547 9.3005
R2030 VTAIL.n503 VTAIL.n502 9.3005
R2031 VTAIL.n554 VTAIL.n553 9.3005
R2032 VTAIL.n556 VTAIL.n555 9.3005
R2033 VTAIL.n498 VTAIL.n497 9.3005
R2034 VTAIL.n562 VTAIL.n561 9.3005
R2035 VTAIL.n564 VTAIL.n563 9.3005
R2036 VTAIL.n571 VTAIL.n570 9.3005
R2037 VTAIL.n494 VTAIL.n493 9.3005
R2038 VTAIL.n507 VTAIL.n506 9.3005
R2039 VTAIL.n540 VTAIL.n539 9.3005
R2040 VTAIL.n538 VTAIL.n537 9.3005
R2041 VTAIL.n511 VTAIL.n510 9.3005
R2042 VTAIL.n532 VTAIL.n531 9.3005
R2043 VTAIL.n530 VTAIL.n529 9.3005
R2044 VTAIL.n515 VTAIL.n514 9.3005
R2045 VTAIL.n524 VTAIL.n523 9.3005
R2046 VTAIL.n522 VTAIL.n521 9.3005
R2047 VTAIL.n464 VTAIL.n463 9.3005
R2048 VTAIL.n466 VTAIL.n465 9.3005
R2049 VTAIL.n421 VTAIL.n420 9.3005
R2050 VTAIL.n472 VTAIL.n471 9.3005
R2051 VTAIL.n474 VTAIL.n473 9.3005
R2052 VTAIL.n416 VTAIL.n415 9.3005
R2053 VTAIL.n480 VTAIL.n479 9.3005
R2054 VTAIL.n482 VTAIL.n481 9.3005
R2055 VTAIL.n489 VTAIL.n488 9.3005
R2056 VTAIL.n412 VTAIL.n411 9.3005
R2057 VTAIL.n425 VTAIL.n424 9.3005
R2058 VTAIL.n458 VTAIL.n457 9.3005
R2059 VTAIL.n456 VTAIL.n455 9.3005
R2060 VTAIL.n429 VTAIL.n428 9.3005
R2061 VTAIL.n450 VTAIL.n449 9.3005
R2062 VTAIL.n448 VTAIL.n447 9.3005
R2063 VTAIL.n433 VTAIL.n432 9.3005
R2064 VTAIL.n442 VTAIL.n441 9.3005
R2065 VTAIL.n440 VTAIL.n439 9.3005
R2066 VTAIL.n382 VTAIL.n381 9.3005
R2067 VTAIL.n384 VTAIL.n383 9.3005
R2068 VTAIL.n339 VTAIL.n338 9.3005
R2069 VTAIL.n390 VTAIL.n389 9.3005
R2070 VTAIL.n392 VTAIL.n391 9.3005
R2071 VTAIL.n334 VTAIL.n333 9.3005
R2072 VTAIL.n398 VTAIL.n397 9.3005
R2073 VTAIL.n400 VTAIL.n399 9.3005
R2074 VTAIL.n407 VTAIL.n406 9.3005
R2075 VTAIL.n330 VTAIL.n329 9.3005
R2076 VTAIL.n343 VTAIL.n342 9.3005
R2077 VTAIL.n376 VTAIL.n375 9.3005
R2078 VTAIL.n374 VTAIL.n373 9.3005
R2079 VTAIL.n347 VTAIL.n346 9.3005
R2080 VTAIL.n368 VTAIL.n367 9.3005
R2081 VTAIL.n366 VTAIL.n365 9.3005
R2082 VTAIL.n351 VTAIL.n350 9.3005
R2083 VTAIL.n360 VTAIL.n359 9.3005
R2084 VTAIL.n358 VTAIL.n357 9.3005
R2085 VTAIL.n300 VTAIL.n299 9.3005
R2086 VTAIL.n302 VTAIL.n301 9.3005
R2087 VTAIL.n257 VTAIL.n256 9.3005
R2088 VTAIL.n308 VTAIL.n307 9.3005
R2089 VTAIL.n310 VTAIL.n309 9.3005
R2090 VTAIL.n252 VTAIL.n251 9.3005
R2091 VTAIL.n316 VTAIL.n315 9.3005
R2092 VTAIL.n318 VTAIL.n317 9.3005
R2093 VTAIL.n325 VTAIL.n324 9.3005
R2094 VTAIL.n248 VTAIL.n247 9.3005
R2095 VTAIL.n261 VTAIL.n260 9.3005
R2096 VTAIL.n294 VTAIL.n293 9.3005
R2097 VTAIL.n292 VTAIL.n291 9.3005
R2098 VTAIL.n265 VTAIL.n264 9.3005
R2099 VTAIL.n286 VTAIL.n285 9.3005
R2100 VTAIL.n284 VTAIL.n283 9.3005
R2101 VTAIL.n269 VTAIL.n268 9.3005
R2102 VTAIL.n278 VTAIL.n277 9.3005
R2103 VTAIL.n276 VTAIL.n275 9.3005
R2104 VTAIL.n617 VTAIL.n592 8.92171
R2105 VTAIL.n630 VTAIL.n584 8.92171
R2106 VTAIL.n43 VTAIL.n18 8.92171
R2107 VTAIL.n56 VTAIL.n10 8.92171
R2108 VTAIL.n125 VTAIL.n100 8.92171
R2109 VTAIL.n138 VTAIL.n92 8.92171
R2110 VTAIL.n207 VTAIL.n182 8.92171
R2111 VTAIL.n220 VTAIL.n174 8.92171
R2112 VTAIL.n549 VTAIL.n503 8.92171
R2113 VTAIL.n536 VTAIL.n511 8.92171
R2114 VTAIL.n467 VTAIL.n421 8.92171
R2115 VTAIL.n454 VTAIL.n429 8.92171
R2116 VTAIL.n385 VTAIL.n339 8.92171
R2117 VTAIL.n372 VTAIL.n347 8.92171
R2118 VTAIL.n303 VTAIL.n257 8.92171
R2119 VTAIL.n290 VTAIL.n265 8.92171
R2120 VTAIL.n618 VTAIL.n590 8.14595
R2121 VTAIL.n629 VTAIL.n586 8.14595
R2122 VTAIL.n44 VTAIL.n16 8.14595
R2123 VTAIL.n55 VTAIL.n12 8.14595
R2124 VTAIL.n126 VTAIL.n98 8.14595
R2125 VTAIL.n137 VTAIL.n94 8.14595
R2126 VTAIL.n208 VTAIL.n180 8.14595
R2127 VTAIL.n219 VTAIL.n176 8.14595
R2128 VTAIL.n548 VTAIL.n505 8.14595
R2129 VTAIL.n537 VTAIL.n509 8.14595
R2130 VTAIL.n466 VTAIL.n423 8.14595
R2131 VTAIL.n455 VTAIL.n427 8.14595
R2132 VTAIL.n384 VTAIL.n341 8.14595
R2133 VTAIL.n373 VTAIL.n345 8.14595
R2134 VTAIL.n302 VTAIL.n259 8.14595
R2135 VTAIL.n291 VTAIL.n263 8.14595
R2136 VTAIL.n622 VTAIL.n621 7.3702
R2137 VTAIL.n626 VTAIL.n625 7.3702
R2138 VTAIL.n48 VTAIL.n47 7.3702
R2139 VTAIL.n52 VTAIL.n51 7.3702
R2140 VTAIL.n130 VTAIL.n129 7.3702
R2141 VTAIL.n134 VTAIL.n133 7.3702
R2142 VTAIL.n212 VTAIL.n211 7.3702
R2143 VTAIL.n216 VTAIL.n215 7.3702
R2144 VTAIL.n545 VTAIL.n544 7.3702
R2145 VTAIL.n541 VTAIL.n540 7.3702
R2146 VTAIL.n463 VTAIL.n462 7.3702
R2147 VTAIL.n459 VTAIL.n458 7.3702
R2148 VTAIL.n381 VTAIL.n380 7.3702
R2149 VTAIL.n377 VTAIL.n376 7.3702
R2150 VTAIL.n299 VTAIL.n298 7.3702
R2151 VTAIL.n295 VTAIL.n294 7.3702
R2152 VTAIL.n622 VTAIL.n588 6.59444
R2153 VTAIL.n625 VTAIL.n588 6.59444
R2154 VTAIL.n48 VTAIL.n14 6.59444
R2155 VTAIL.n51 VTAIL.n14 6.59444
R2156 VTAIL.n130 VTAIL.n96 6.59444
R2157 VTAIL.n133 VTAIL.n96 6.59444
R2158 VTAIL.n212 VTAIL.n178 6.59444
R2159 VTAIL.n215 VTAIL.n178 6.59444
R2160 VTAIL.n544 VTAIL.n507 6.59444
R2161 VTAIL.n541 VTAIL.n507 6.59444
R2162 VTAIL.n462 VTAIL.n425 6.59444
R2163 VTAIL.n459 VTAIL.n425 6.59444
R2164 VTAIL.n380 VTAIL.n343 6.59444
R2165 VTAIL.n377 VTAIL.n343 6.59444
R2166 VTAIL.n298 VTAIL.n261 6.59444
R2167 VTAIL.n295 VTAIL.n261 6.59444
R2168 VTAIL.n621 VTAIL.n590 5.81868
R2169 VTAIL.n626 VTAIL.n586 5.81868
R2170 VTAIL.n47 VTAIL.n16 5.81868
R2171 VTAIL.n52 VTAIL.n12 5.81868
R2172 VTAIL.n129 VTAIL.n98 5.81868
R2173 VTAIL.n134 VTAIL.n94 5.81868
R2174 VTAIL.n211 VTAIL.n180 5.81868
R2175 VTAIL.n216 VTAIL.n176 5.81868
R2176 VTAIL.n545 VTAIL.n505 5.81868
R2177 VTAIL.n540 VTAIL.n509 5.81868
R2178 VTAIL.n463 VTAIL.n423 5.81868
R2179 VTAIL.n458 VTAIL.n427 5.81868
R2180 VTAIL.n381 VTAIL.n341 5.81868
R2181 VTAIL.n376 VTAIL.n345 5.81868
R2182 VTAIL.n299 VTAIL.n259 5.81868
R2183 VTAIL.n294 VTAIL.n263 5.81868
R2184 VTAIL.n618 VTAIL.n617 5.04292
R2185 VTAIL.n630 VTAIL.n629 5.04292
R2186 VTAIL.n44 VTAIL.n43 5.04292
R2187 VTAIL.n56 VTAIL.n55 5.04292
R2188 VTAIL.n126 VTAIL.n125 5.04292
R2189 VTAIL.n138 VTAIL.n137 5.04292
R2190 VTAIL.n208 VTAIL.n207 5.04292
R2191 VTAIL.n220 VTAIL.n219 5.04292
R2192 VTAIL.n549 VTAIL.n548 5.04292
R2193 VTAIL.n537 VTAIL.n536 5.04292
R2194 VTAIL.n467 VTAIL.n466 5.04292
R2195 VTAIL.n455 VTAIL.n454 5.04292
R2196 VTAIL.n385 VTAIL.n384 5.04292
R2197 VTAIL.n373 VTAIL.n372 5.04292
R2198 VTAIL.n303 VTAIL.n302 5.04292
R2199 VTAIL.n291 VTAIL.n290 5.04292
R2200 VTAIL.n522 VTAIL.n518 4.38563
R2201 VTAIL.n440 VTAIL.n436 4.38563
R2202 VTAIL.n358 VTAIL.n354 4.38563
R2203 VTAIL.n276 VTAIL.n272 4.38563
R2204 VTAIL.n603 VTAIL.n599 4.38563
R2205 VTAIL.n29 VTAIL.n25 4.38563
R2206 VTAIL.n111 VTAIL.n107 4.38563
R2207 VTAIL.n193 VTAIL.n189 4.38563
R2208 VTAIL.n614 VTAIL.n592 4.26717
R2209 VTAIL.n633 VTAIL.n584 4.26717
R2210 VTAIL.n40 VTAIL.n18 4.26717
R2211 VTAIL.n59 VTAIL.n10 4.26717
R2212 VTAIL.n122 VTAIL.n100 4.26717
R2213 VTAIL.n141 VTAIL.n92 4.26717
R2214 VTAIL.n204 VTAIL.n182 4.26717
R2215 VTAIL.n223 VTAIL.n174 4.26717
R2216 VTAIL.n552 VTAIL.n503 4.26717
R2217 VTAIL.n533 VTAIL.n511 4.26717
R2218 VTAIL.n470 VTAIL.n421 4.26717
R2219 VTAIL.n451 VTAIL.n429 4.26717
R2220 VTAIL.n388 VTAIL.n339 4.26717
R2221 VTAIL.n369 VTAIL.n347 4.26717
R2222 VTAIL.n306 VTAIL.n257 4.26717
R2223 VTAIL.n287 VTAIL.n265 4.26717
R2224 VTAIL.n613 VTAIL.n594 3.49141
R2225 VTAIL.n634 VTAIL.n582 3.49141
R2226 VTAIL.n39 VTAIL.n20 3.49141
R2227 VTAIL.n60 VTAIL.n8 3.49141
R2228 VTAIL.n121 VTAIL.n102 3.49141
R2229 VTAIL.n142 VTAIL.n90 3.49141
R2230 VTAIL.n203 VTAIL.n184 3.49141
R2231 VTAIL.n224 VTAIL.n172 3.49141
R2232 VTAIL.n553 VTAIL.n501 3.49141
R2233 VTAIL.n532 VTAIL.n513 3.49141
R2234 VTAIL.n471 VTAIL.n419 3.49141
R2235 VTAIL.n450 VTAIL.n431 3.49141
R2236 VTAIL.n389 VTAIL.n337 3.49141
R2237 VTAIL.n368 VTAIL.n349 3.49141
R2238 VTAIL.n307 VTAIL.n255 3.49141
R2239 VTAIL.n286 VTAIL.n267 3.49141
R2240 VTAIL.n610 VTAIL.n609 2.71565
R2241 VTAIL.n638 VTAIL.n637 2.71565
R2242 VTAIL.n36 VTAIL.n35 2.71565
R2243 VTAIL.n64 VTAIL.n63 2.71565
R2244 VTAIL.n118 VTAIL.n117 2.71565
R2245 VTAIL.n146 VTAIL.n145 2.71565
R2246 VTAIL.n200 VTAIL.n199 2.71565
R2247 VTAIL.n228 VTAIL.n227 2.71565
R2248 VTAIL.n557 VTAIL.n556 2.71565
R2249 VTAIL.n529 VTAIL.n528 2.71565
R2250 VTAIL.n475 VTAIL.n474 2.71565
R2251 VTAIL.n447 VTAIL.n446 2.71565
R2252 VTAIL.n393 VTAIL.n392 2.71565
R2253 VTAIL.n365 VTAIL.n364 2.71565
R2254 VTAIL.n311 VTAIL.n310 2.71565
R2255 VTAIL.n283 VTAIL.n282 2.71565
R2256 VTAIL.n409 VTAIL.n327 2.17291
R2257 VTAIL.n573 VTAIL.n491 2.17291
R2258 VTAIL.n245 VTAIL.n163 2.17291
R2259 VTAIL.n606 VTAIL.n596 1.93989
R2260 VTAIL.n642 VTAIL.n580 1.93989
R2261 VTAIL.n654 VTAIL.n574 1.93989
R2262 VTAIL.n32 VTAIL.n22 1.93989
R2263 VTAIL.n68 VTAIL.n6 1.93989
R2264 VTAIL.n80 VTAIL.n0 1.93989
R2265 VTAIL.n114 VTAIL.n104 1.93989
R2266 VTAIL.n150 VTAIL.n88 1.93989
R2267 VTAIL.n162 VTAIL.n82 1.93989
R2268 VTAIL.n196 VTAIL.n186 1.93989
R2269 VTAIL.n232 VTAIL.n170 1.93989
R2270 VTAIL.n244 VTAIL.n164 1.93989
R2271 VTAIL.n572 VTAIL.n492 1.93989
R2272 VTAIL.n560 VTAIL.n498 1.93989
R2273 VTAIL.n525 VTAIL.n515 1.93989
R2274 VTAIL.n490 VTAIL.n410 1.93989
R2275 VTAIL.n478 VTAIL.n416 1.93989
R2276 VTAIL.n443 VTAIL.n433 1.93989
R2277 VTAIL.n408 VTAIL.n328 1.93989
R2278 VTAIL.n396 VTAIL.n334 1.93989
R2279 VTAIL.n361 VTAIL.n351 1.93989
R2280 VTAIL.n326 VTAIL.n246 1.93989
R2281 VTAIL.n314 VTAIL.n252 1.93989
R2282 VTAIL.n279 VTAIL.n269 1.93989
R2283 VTAIL.n605 VTAIL.n598 1.16414
R2284 VTAIL.n643 VTAIL.n578 1.16414
R2285 VTAIL.n652 VTAIL.n651 1.16414
R2286 VTAIL.n31 VTAIL.n24 1.16414
R2287 VTAIL.n69 VTAIL.n4 1.16414
R2288 VTAIL.n78 VTAIL.n77 1.16414
R2289 VTAIL.n113 VTAIL.n106 1.16414
R2290 VTAIL.n151 VTAIL.n86 1.16414
R2291 VTAIL.n160 VTAIL.n159 1.16414
R2292 VTAIL.n195 VTAIL.n188 1.16414
R2293 VTAIL.n233 VTAIL.n168 1.16414
R2294 VTAIL.n242 VTAIL.n241 1.16414
R2295 VTAIL.n570 VTAIL.n569 1.16414
R2296 VTAIL.n561 VTAIL.n496 1.16414
R2297 VTAIL.n524 VTAIL.n517 1.16414
R2298 VTAIL.n488 VTAIL.n487 1.16414
R2299 VTAIL.n479 VTAIL.n414 1.16414
R2300 VTAIL.n442 VTAIL.n435 1.16414
R2301 VTAIL.n406 VTAIL.n405 1.16414
R2302 VTAIL.n397 VTAIL.n332 1.16414
R2303 VTAIL.n360 VTAIL.n353 1.16414
R2304 VTAIL.n324 VTAIL.n323 1.16414
R2305 VTAIL.n315 VTAIL.n250 1.16414
R2306 VTAIL.n278 VTAIL.n271 1.16414
R2307 VTAIL VTAIL.n81 1.1449
R2308 VTAIL VTAIL.n655 1.02852
R2309 VTAIL.n491 VTAIL.n409 0.470328
R2310 VTAIL.n163 VTAIL.n81 0.470328
R2311 VTAIL.n602 VTAIL.n601 0.388379
R2312 VTAIL.n647 VTAIL.n646 0.388379
R2313 VTAIL.n648 VTAIL.n576 0.388379
R2314 VTAIL.n28 VTAIL.n27 0.388379
R2315 VTAIL.n73 VTAIL.n72 0.388379
R2316 VTAIL.n74 VTAIL.n2 0.388379
R2317 VTAIL.n110 VTAIL.n109 0.388379
R2318 VTAIL.n155 VTAIL.n154 0.388379
R2319 VTAIL.n156 VTAIL.n84 0.388379
R2320 VTAIL.n192 VTAIL.n191 0.388379
R2321 VTAIL.n237 VTAIL.n236 0.388379
R2322 VTAIL.n238 VTAIL.n166 0.388379
R2323 VTAIL.n566 VTAIL.n494 0.388379
R2324 VTAIL.n565 VTAIL.n564 0.388379
R2325 VTAIL.n521 VTAIL.n520 0.388379
R2326 VTAIL.n484 VTAIL.n412 0.388379
R2327 VTAIL.n483 VTAIL.n482 0.388379
R2328 VTAIL.n439 VTAIL.n438 0.388379
R2329 VTAIL.n402 VTAIL.n330 0.388379
R2330 VTAIL.n401 VTAIL.n400 0.388379
R2331 VTAIL.n357 VTAIL.n356 0.388379
R2332 VTAIL.n320 VTAIL.n248 0.388379
R2333 VTAIL.n319 VTAIL.n318 0.388379
R2334 VTAIL.n275 VTAIL.n274 0.388379
R2335 VTAIL.n604 VTAIL.n603 0.155672
R2336 VTAIL.n604 VTAIL.n595 0.155672
R2337 VTAIL.n611 VTAIL.n595 0.155672
R2338 VTAIL.n612 VTAIL.n611 0.155672
R2339 VTAIL.n612 VTAIL.n591 0.155672
R2340 VTAIL.n619 VTAIL.n591 0.155672
R2341 VTAIL.n620 VTAIL.n619 0.155672
R2342 VTAIL.n620 VTAIL.n587 0.155672
R2343 VTAIL.n627 VTAIL.n587 0.155672
R2344 VTAIL.n628 VTAIL.n627 0.155672
R2345 VTAIL.n628 VTAIL.n583 0.155672
R2346 VTAIL.n635 VTAIL.n583 0.155672
R2347 VTAIL.n636 VTAIL.n635 0.155672
R2348 VTAIL.n636 VTAIL.n579 0.155672
R2349 VTAIL.n644 VTAIL.n579 0.155672
R2350 VTAIL.n645 VTAIL.n644 0.155672
R2351 VTAIL.n645 VTAIL.n575 0.155672
R2352 VTAIL.n653 VTAIL.n575 0.155672
R2353 VTAIL.n30 VTAIL.n29 0.155672
R2354 VTAIL.n30 VTAIL.n21 0.155672
R2355 VTAIL.n37 VTAIL.n21 0.155672
R2356 VTAIL.n38 VTAIL.n37 0.155672
R2357 VTAIL.n38 VTAIL.n17 0.155672
R2358 VTAIL.n45 VTAIL.n17 0.155672
R2359 VTAIL.n46 VTAIL.n45 0.155672
R2360 VTAIL.n46 VTAIL.n13 0.155672
R2361 VTAIL.n53 VTAIL.n13 0.155672
R2362 VTAIL.n54 VTAIL.n53 0.155672
R2363 VTAIL.n54 VTAIL.n9 0.155672
R2364 VTAIL.n61 VTAIL.n9 0.155672
R2365 VTAIL.n62 VTAIL.n61 0.155672
R2366 VTAIL.n62 VTAIL.n5 0.155672
R2367 VTAIL.n70 VTAIL.n5 0.155672
R2368 VTAIL.n71 VTAIL.n70 0.155672
R2369 VTAIL.n71 VTAIL.n1 0.155672
R2370 VTAIL.n79 VTAIL.n1 0.155672
R2371 VTAIL.n112 VTAIL.n111 0.155672
R2372 VTAIL.n112 VTAIL.n103 0.155672
R2373 VTAIL.n119 VTAIL.n103 0.155672
R2374 VTAIL.n120 VTAIL.n119 0.155672
R2375 VTAIL.n120 VTAIL.n99 0.155672
R2376 VTAIL.n127 VTAIL.n99 0.155672
R2377 VTAIL.n128 VTAIL.n127 0.155672
R2378 VTAIL.n128 VTAIL.n95 0.155672
R2379 VTAIL.n135 VTAIL.n95 0.155672
R2380 VTAIL.n136 VTAIL.n135 0.155672
R2381 VTAIL.n136 VTAIL.n91 0.155672
R2382 VTAIL.n143 VTAIL.n91 0.155672
R2383 VTAIL.n144 VTAIL.n143 0.155672
R2384 VTAIL.n144 VTAIL.n87 0.155672
R2385 VTAIL.n152 VTAIL.n87 0.155672
R2386 VTAIL.n153 VTAIL.n152 0.155672
R2387 VTAIL.n153 VTAIL.n83 0.155672
R2388 VTAIL.n161 VTAIL.n83 0.155672
R2389 VTAIL.n194 VTAIL.n193 0.155672
R2390 VTAIL.n194 VTAIL.n185 0.155672
R2391 VTAIL.n201 VTAIL.n185 0.155672
R2392 VTAIL.n202 VTAIL.n201 0.155672
R2393 VTAIL.n202 VTAIL.n181 0.155672
R2394 VTAIL.n209 VTAIL.n181 0.155672
R2395 VTAIL.n210 VTAIL.n209 0.155672
R2396 VTAIL.n210 VTAIL.n177 0.155672
R2397 VTAIL.n217 VTAIL.n177 0.155672
R2398 VTAIL.n218 VTAIL.n217 0.155672
R2399 VTAIL.n218 VTAIL.n173 0.155672
R2400 VTAIL.n225 VTAIL.n173 0.155672
R2401 VTAIL.n226 VTAIL.n225 0.155672
R2402 VTAIL.n226 VTAIL.n169 0.155672
R2403 VTAIL.n234 VTAIL.n169 0.155672
R2404 VTAIL.n235 VTAIL.n234 0.155672
R2405 VTAIL.n235 VTAIL.n165 0.155672
R2406 VTAIL.n243 VTAIL.n165 0.155672
R2407 VTAIL.n571 VTAIL.n493 0.155672
R2408 VTAIL.n563 VTAIL.n493 0.155672
R2409 VTAIL.n563 VTAIL.n562 0.155672
R2410 VTAIL.n562 VTAIL.n497 0.155672
R2411 VTAIL.n555 VTAIL.n497 0.155672
R2412 VTAIL.n555 VTAIL.n554 0.155672
R2413 VTAIL.n554 VTAIL.n502 0.155672
R2414 VTAIL.n547 VTAIL.n502 0.155672
R2415 VTAIL.n547 VTAIL.n546 0.155672
R2416 VTAIL.n546 VTAIL.n506 0.155672
R2417 VTAIL.n539 VTAIL.n506 0.155672
R2418 VTAIL.n539 VTAIL.n538 0.155672
R2419 VTAIL.n538 VTAIL.n510 0.155672
R2420 VTAIL.n531 VTAIL.n510 0.155672
R2421 VTAIL.n531 VTAIL.n530 0.155672
R2422 VTAIL.n530 VTAIL.n514 0.155672
R2423 VTAIL.n523 VTAIL.n514 0.155672
R2424 VTAIL.n523 VTAIL.n522 0.155672
R2425 VTAIL.n489 VTAIL.n411 0.155672
R2426 VTAIL.n481 VTAIL.n411 0.155672
R2427 VTAIL.n481 VTAIL.n480 0.155672
R2428 VTAIL.n480 VTAIL.n415 0.155672
R2429 VTAIL.n473 VTAIL.n415 0.155672
R2430 VTAIL.n473 VTAIL.n472 0.155672
R2431 VTAIL.n472 VTAIL.n420 0.155672
R2432 VTAIL.n465 VTAIL.n420 0.155672
R2433 VTAIL.n465 VTAIL.n464 0.155672
R2434 VTAIL.n464 VTAIL.n424 0.155672
R2435 VTAIL.n457 VTAIL.n424 0.155672
R2436 VTAIL.n457 VTAIL.n456 0.155672
R2437 VTAIL.n456 VTAIL.n428 0.155672
R2438 VTAIL.n449 VTAIL.n428 0.155672
R2439 VTAIL.n449 VTAIL.n448 0.155672
R2440 VTAIL.n448 VTAIL.n432 0.155672
R2441 VTAIL.n441 VTAIL.n432 0.155672
R2442 VTAIL.n441 VTAIL.n440 0.155672
R2443 VTAIL.n407 VTAIL.n329 0.155672
R2444 VTAIL.n399 VTAIL.n329 0.155672
R2445 VTAIL.n399 VTAIL.n398 0.155672
R2446 VTAIL.n398 VTAIL.n333 0.155672
R2447 VTAIL.n391 VTAIL.n333 0.155672
R2448 VTAIL.n391 VTAIL.n390 0.155672
R2449 VTAIL.n390 VTAIL.n338 0.155672
R2450 VTAIL.n383 VTAIL.n338 0.155672
R2451 VTAIL.n383 VTAIL.n382 0.155672
R2452 VTAIL.n382 VTAIL.n342 0.155672
R2453 VTAIL.n375 VTAIL.n342 0.155672
R2454 VTAIL.n375 VTAIL.n374 0.155672
R2455 VTAIL.n374 VTAIL.n346 0.155672
R2456 VTAIL.n367 VTAIL.n346 0.155672
R2457 VTAIL.n367 VTAIL.n366 0.155672
R2458 VTAIL.n366 VTAIL.n350 0.155672
R2459 VTAIL.n359 VTAIL.n350 0.155672
R2460 VTAIL.n359 VTAIL.n358 0.155672
R2461 VTAIL.n325 VTAIL.n247 0.155672
R2462 VTAIL.n317 VTAIL.n247 0.155672
R2463 VTAIL.n317 VTAIL.n316 0.155672
R2464 VTAIL.n316 VTAIL.n251 0.155672
R2465 VTAIL.n309 VTAIL.n251 0.155672
R2466 VTAIL.n309 VTAIL.n308 0.155672
R2467 VTAIL.n308 VTAIL.n256 0.155672
R2468 VTAIL.n301 VTAIL.n256 0.155672
R2469 VTAIL.n301 VTAIL.n300 0.155672
R2470 VTAIL.n300 VTAIL.n260 0.155672
R2471 VTAIL.n293 VTAIL.n260 0.155672
R2472 VTAIL.n293 VTAIL.n292 0.155672
R2473 VTAIL.n292 VTAIL.n264 0.155672
R2474 VTAIL.n285 VTAIL.n264 0.155672
R2475 VTAIL.n285 VTAIL.n284 0.155672
R2476 VTAIL.n284 VTAIL.n268 0.155672
R2477 VTAIL.n277 VTAIL.n268 0.155672
R2478 VTAIL.n277 VTAIL.n276 0.155672
R2479 VDD1 VDD1.n1 105.918
R2480 VDD1 VDD1.n0 62.5306
R2481 VDD1.n0 VDD1.t0 1.34561
R2482 VDD1.n0 VDD1.t3 1.34561
R2483 VDD1.n1 VDD1.t1 1.34561
R2484 VDD1.n1 VDD1.t2 1.34561
R2485 VN.n0 VN.t0 197.677
R2486 VN.n1 VN.t2 197.677
R2487 VN.n0 VN.t1 197.042
R2488 VN.n1 VN.t3 197.042
R2489 VN VN.n1 53.1602
R2490 VN VN.n0 5.85334
R2491 VDD2.n2 VDD2.n0 105.394
R2492 VDD2.n2 VDD2.n1 62.4724
R2493 VDD2.n1 VDD2.t0 1.34561
R2494 VDD2.n1 VDD2.t1 1.34561
R2495 VDD2.n0 VDD2.t3 1.34561
R2496 VDD2.n0 VDD2.t2 1.34561
R2497 VDD2 VDD2.n2 0.0586897
C0 VP VN 6.39888f
C1 VDD2 VTAIL 6.11636f
C2 VDD1 VN 0.148792f
C3 VDD1 VP 5.78934f
C4 VDD2 VN 5.57039f
C5 VDD2 VP 0.368378f
C6 VDD1 VDD2 0.92934f
C7 VN VTAIL 5.30323f
C8 VP VTAIL 5.31734f
C9 VDD1 VTAIL 6.0649f
C10 VDD2 B 3.739515f
C11 VDD1 B 8.033219f
C12 VTAIL B 11.460465f
C13 VN B 10.19492f
C14 VP B 8.256827f
C15 VDD2.t3 B 0.309721f
C16 VDD2.t2 B 0.309721f
C17 VDD2.n0 B 3.53642f
C18 VDD2.t0 B 0.309721f
C19 VDD2.t1 B 0.309721f
C20 VDD2.n1 B 2.79891f
C21 VDD2.n2 B 3.93368f
C22 VN.t0 B 2.63021f
C23 VN.t1 B 2.62696f
C24 VN.n0 B 1.74701f
C25 VN.t2 B 2.63021f
C26 VN.t3 B 2.62696f
C27 VN.n1 B 3.20223f
C28 VDD1.t0 B 0.31239f
C29 VDD1.t3 B 0.31239f
C30 VDD1.n0 B 2.82341f
C31 VDD1.t1 B 0.31239f
C32 VDD1.t2 B 0.31239f
C33 VDD1.n1 B 3.59413f
C34 VTAIL.n0 B 0.020733f
C35 VTAIL.n1 B 0.015652f
C36 VTAIL.n2 B 0.008411f
C37 VTAIL.n3 B 0.01988f
C38 VTAIL.n4 B 0.008905f
C39 VTAIL.n5 B 0.015652f
C40 VTAIL.n6 B 0.008411f
C41 VTAIL.n7 B 0.01988f
C42 VTAIL.n8 B 0.008905f
C43 VTAIL.n9 B 0.015652f
C44 VTAIL.n10 B 0.008411f
C45 VTAIL.n11 B 0.01988f
C46 VTAIL.n12 B 0.008905f
C47 VTAIL.n13 B 0.015652f
C48 VTAIL.n14 B 0.008411f
C49 VTAIL.n15 B 0.01988f
C50 VTAIL.n16 B 0.008905f
C51 VTAIL.n17 B 0.015652f
C52 VTAIL.n18 B 0.008411f
C53 VTAIL.n19 B 0.01988f
C54 VTAIL.n20 B 0.008905f
C55 VTAIL.n21 B 0.015652f
C56 VTAIL.n22 B 0.008411f
C57 VTAIL.n23 B 0.01988f
C58 VTAIL.n24 B 0.008905f
C59 VTAIL.n25 B 0.100987f
C60 VTAIL.t0 B 0.032764f
C61 VTAIL.n26 B 0.01491f
C62 VTAIL.n27 B 0.011744f
C63 VTAIL.n28 B 0.008411f
C64 VTAIL.n29 B 0.998259f
C65 VTAIL.n30 B 0.015652f
C66 VTAIL.n31 B 0.008411f
C67 VTAIL.n32 B 0.008905f
C68 VTAIL.n33 B 0.01988f
C69 VTAIL.n34 B 0.01988f
C70 VTAIL.n35 B 0.008905f
C71 VTAIL.n36 B 0.008411f
C72 VTAIL.n37 B 0.015652f
C73 VTAIL.n38 B 0.015652f
C74 VTAIL.n39 B 0.008411f
C75 VTAIL.n40 B 0.008905f
C76 VTAIL.n41 B 0.01988f
C77 VTAIL.n42 B 0.01988f
C78 VTAIL.n43 B 0.008905f
C79 VTAIL.n44 B 0.008411f
C80 VTAIL.n45 B 0.015652f
C81 VTAIL.n46 B 0.015652f
C82 VTAIL.n47 B 0.008411f
C83 VTAIL.n48 B 0.008905f
C84 VTAIL.n49 B 0.01988f
C85 VTAIL.n50 B 0.01988f
C86 VTAIL.n51 B 0.008905f
C87 VTAIL.n52 B 0.008411f
C88 VTAIL.n53 B 0.015652f
C89 VTAIL.n54 B 0.015652f
C90 VTAIL.n55 B 0.008411f
C91 VTAIL.n56 B 0.008905f
C92 VTAIL.n57 B 0.01988f
C93 VTAIL.n58 B 0.01988f
C94 VTAIL.n59 B 0.008905f
C95 VTAIL.n60 B 0.008411f
C96 VTAIL.n61 B 0.015652f
C97 VTAIL.n62 B 0.015652f
C98 VTAIL.n63 B 0.008411f
C99 VTAIL.n64 B 0.008905f
C100 VTAIL.n65 B 0.01988f
C101 VTAIL.n66 B 0.01988f
C102 VTAIL.n67 B 0.01988f
C103 VTAIL.n68 B 0.008905f
C104 VTAIL.n69 B 0.008411f
C105 VTAIL.n70 B 0.015652f
C106 VTAIL.n71 B 0.015652f
C107 VTAIL.n72 B 0.008411f
C108 VTAIL.n73 B 0.008658f
C109 VTAIL.n74 B 0.008658f
C110 VTAIL.n75 B 0.01988f
C111 VTAIL.n76 B 0.040796f
C112 VTAIL.n77 B 0.008905f
C113 VTAIL.n78 B 0.008411f
C114 VTAIL.n79 B 0.037889f
C115 VTAIL.n80 B 0.022648f
C116 VTAIL.n81 B 0.095747f
C117 VTAIL.n82 B 0.020733f
C118 VTAIL.n83 B 0.015652f
C119 VTAIL.n84 B 0.008411f
C120 VTAIL.n85 B 0.01988f
C121 VTAIL.n86 B 0.008905f
C122 VTAIL.n87 B 0.015652f
C123 VTAIL.n88 B 0.008411f
C124 VTAIL.n89 B 0.01988f
C125 VTAIL.n90 B 0.008905f
C126 VTAIL.n91 B 0.015652f
C127 VTAIL.n92 B 0.008411f
C128 VTAIL.n93 B 0.01988f
C129 VTAIL.n94 B 0.008905f
C130 VTAIL.n95 B 0.015652f
C131 VTAIL.n96 B 0.008411f
C132 VTAIL.n97 B 0.01988f
C133 VTAIL.n98 B 0.008905f
C134 VTAIL.n99 B 0.015652f
C135 VTAIL.n100 B 0.008411f
C136 VTAIL.n101 B 0.01988f
C137 VTAIL.n102 B 0.008905f
C138 VTAIL.n103 B 0.015652f
C139 VTAIL.n104 B 0.008411f
C140 VTAIL.n105 B 0.01988f
C141 VTAIL.n106 B 0.008905f
C142 VTAIL.n107 B 0.100987f
C143 VTAIL.t5 B 0.032764f
C144 VTAIL.n108 B 0.01491f
C145 VTAIL.n109 B 0.011744f
C146 VTAIL.n110 B 0.008411f
C147 VTAIL.n111 B 0.998259f
C148 VTAIL.n112 B 0.015652f
C149 VTAIL.n113 B 0.008411f
C150 VTAIL.n114 B 0.008905f
C151 VTAIL.n115 B 0.01988f
C152 VTAIL.n116 B 0.01988f
C153 VTAIL.n117 B 0.008905f
C154 VTAIL.n118 B 0.008411f
C155 VTAIL.n119 B 0.015652f
C156 VTAIL.n120 B 0.015652f
C157 VTAIL.n121 B 0.008411f
C158 VTAIL.n122 B 0.008905f
C159 VTAIL.n123 B 0.01988f
C160 VTAIL.n124 B 0.01988f
C161 VTAIL.n125 B 0.008905f
C162 VTAIL.n126 B 0.008411f
C163 VTAIL.n127 B 0.015652f
C164 VTAIL.n128 B 0.015652f
C165 VTAIL.n129 B 0.008411f
C166 VTAIL.n130 B 0.008905f
C167 VTAIL.n131 B 0.01988f
C168 VTAIL.n132 B 0.01988f
C169 VTAIL.n133 B 0.008905f
C170 VTAIL.n134 B 0.008411f
C171 VTAIL.n135 B 0.015652f
C172 VTAIL.n136 B 0.015652f
C173 VTAIL.n137 B 0.008411f
C174 VTAIL.n138 B 0.008905f
C175 VTAIL.n139 B 0.01988f
C176 VTAIL.n140 B 0.01988f
C177 VTAIL.n141 B 0.008905f
C178 VTAIL.n142 B 0.008411f
C179 VTAIL.n143 B 0.015652f
C180 VTAIL.n144 B 0.015652f
C181 VTAIL.n145 B 0.008411f
C182 VTAIL.n146 B 0.008905f
C183 VTAIL.n147 B 0.01988f
C184 VTAIL.n148 B 0.01988f
C185 VTAIL.n149 B 0.01988f
C186 VTAIL.n150 B 0.008905f
C187 VTAIL.n151 B 0.008411f
C188 VTAIL.n152 B 0.015652f
C189 VTAIL.n153 B 0.015652f
C190 VTAIL.n154 B 0.008411f
C191 VTAIL.n155 B 0.008658f
C192 VTAIL.n156 B 0.008658f
C193 VTAIL.n157 B 0.01988f
C194 VTAIL.n158 B 0.040796f
C195 VTAIL.n159 B 0.008905f
C196 VTAIL.n160 B 0.008411f
C197 VTAIL.n161 B 0.037889f
C198 VTAIL.n162 B 0.022648f
C199 VTAIL.n163 B 0.147594f
C200 VTAIL.n164 B 0.020733f
C201 VTAIL.n165 B 0.015652f
C202 VTAIL.n166 B 0.008411f
C203 VTAIL.n167 B 0.01988f
C204 VTAIL.n168 B 0.008905f
C205 VTAIL.n169 B 0.015652f
C206 VTAIL.n170 B 0.008411f
C207 VTAIL.n171 B 0.01988f
C208 VTAIL.n172 B 0.008905f
C209 VTAIL.n173 B 0.015652f
C210 VTAIL.n174 B 0.008411f
C211 VTAIL.n175 B 0.01988f
C212 VTAIL.n176 B 0.008905f
C213 VTAIL.n177 B 0.015652f
C214 VTAIL.n178 B 0.008411f
C215 VTAIL.n179 B 0.01988f
C216 VTAIL.n180 B 0.008905f
C217 VTAIL.n181 B 0.015652f
C218 VTAIL.n182 B 0.008411f
C219 VTAIL.n183 B 0.01988f
C220 VTAIL.n184 B 0.008905f
C221 VTAIL.n185 B 0.015652f
C222 VTAIL.n186 B 0.008411f
C223 VTAIL.n187 B 0.01988f
C224 VTAIL.n188 B 0.008905f
C225 VTAIL.n189 B 0.100987f
C226 VTAIL.t4 B 0.032764f
C227 VTAIL.n190 B 0.01491f
C228 VTAIL.n191 B 0.011744f
C229 VTAIL.n192 B 0.008411f
C230 VTAIL.n193 B 0.998259f
C231 VTAIL.n194 B 0.015652f
C232 VTAIL.n195 B 0.008411f
C233 VTAIL.n196 B 0.008905f
C234 VTAIL.n197 B 0.01988f
C235 VTAIL.n198 B 0.01988f
C236 VTAIL.n199 B 0.008905f
C237 VTAIL.n200 B 0.008411f
C238 VTAIL.n201 B 0.015652f
C239 VTAIL.n202 B 0.015652f
C240 VTAIL.n203 B 0.008411f
C241 VTAIL.n204 B 0.008905f
C242 VTAIL.n205 B 0.01988f
C243 VTAIL.n206 B 0.01988f
C244 VTAIL.n207 B 0.008905f
C245 VTAIL.n208 B 0.008411f
C246 VTAIL.n209 B 0.015652f
C247 VTAIL.n210 B 0.015652f
C248 VTAIL.n211 B 0.008411f
C249 VTAIL.n212 B 0.008905f
C250 VTAIL.n213 B 0.01988f
C251 VTAIL.n214 B 0.01988f
C252 VTAIL.n215 B 0.008905f
C253 VTAIL.n216 B 0.008411f
C254 VTAIL.n217 B 0.015652f
C255 VTAIL.n218 B 0.015652f
C256 VTAIL.n219 B 0.008411f
C257 VTAIL.n220 B 0.008905f
C258 VTAIL.n221 B 0.01988f
C259 VTAIL.n222 B 0.01988f
C260 VTAIL.n223 B 0.008905f
C261 VTAIL.n224 B 0.008411f
C262 VTAIL.n225 B 0.015652f
C263 VTAIL.n226 B 0.015652f
C264 VTAIL.n227 B 0.008411f
C265 VTAIL.n228 B 0.008905f
C266 VTAIL.n229 B 0.01988f
C267 VTAIL.n230 B 0.01988f
C268 VTAIL.n231 B 0.01988f
C269 VTAIL.n232 B 0.008905f
C270 VTAIL.n233 B 0.008411f
C271 VTAIL.n234 B 0.015652f
C272 VTAIL.n235 B 0.015652f
C273 VTAIL.n236 B 0.008411f
C274 VTAIL.n237 B 0.008658f
C275 VTAIL.n238 B 0.008658f
C276 VTAIL.n239 B 0.01988f
C277 VTAIL.n240 B 0.040796f
C278 VTAIL.n241 B 0.008905f
C279 VTAIL.n242 B 0.008411f
C280 VTAIL.n243 B 0.037889f
C281 VTAIL.n244 B 0.022648f
C282 VTAIL.n245 B 1.08607f
C283 VTAIL.n246 B 0.020733f
C284 VTAIL.n247 B 0.015652f
C285 VTAIL.n248 B 0.008411f
C286 VTAIL.n249 B 0.01988f
C287 VTAIL.n250 B 0.008905f
C288 VTAIL.n251 B 0.015652f
C289 VTAIL.n252 B 0.008411f
C290 VTAIL.n253 B 0.01988f
C291 VTAIL.n254 B 0.01988f
C292 VTAIL.n255 B 0.008905f
C293 VTAIL.n256 B 0.015652f
C294 VTAIL.n257 B 0.008411f
C295 VTAIL.n258 B 0.01988f
C296 VTAIL.n259 B 0.008905f
C297 VTAIL.n260 B 0.015652f
C298 VTAIL.n261 B 0.008411f
C299 VTAIL.n262 B 0.01988f
C300 VTAIL.n263 B 0.008905f
C301 VTAIL.n264 B 0.015652f
C302 VTAIL.n265 B 0.008411f
C303 VTAIL.n266 B 0.01988f
C304 VTAIL.n267 B 0.008905f
C305 VTAIL.n268 B 0.015652f
C306 VTAIL.n269 B 0.008411f
C307 VTAIL.n270 B 0.01988f
C308 VTAIL.n271 B 0.008905f
C309 VTAIL.n272 B 0.100987f
C310 VTAIL.t2 B 0.032764f
C311 VTAIL.n273 B 0.01491f
C312 VTAIL.n274 B 0.011744f
C313 VTAIL.n275 B 0.008411f
C314 VTAIL.n276 B 0.998259f
C315 VTAIL.n277 B 0.015652f
C316 VTAIL.n278 B 0.008411f
C317 VTAIL.n279 B 0.008905f
C318 VTAIL.n280 B 0.01988f
C319 VTAIL.n281 B 0.01988f
C320 VTAIL.n282 B 0.008905f
C321 VTAIL.n283 B 0.008411f
C322 VTAIL.n284 B 0.015652f
C323 VTAIL.n285 B 0.015652f
C324 VTAIL.n286 B 0.008411f
C325 VTAIL.n287 B 0.008905f
C326 VTAIL.n288 B 0.01988f
C327 VTAIL.n289 B 0.01988f
C328 VTAIL.n290 B 0.008905f
C329 VTAIL.n291 B 0.008411f
C330 VTAIL.n292 B 0.015652f
C331 VTAIL.n293 B 0.015652f
C332 VTAIL.n294 B 0.008411f
C333 VTAIL.n295 B 0.008905f
C334 VTAIL.n296 B 0.01988f
C335 VTAIL.n297 B 0.01988f
C336 VTAIL.n298 B 0.008905f
C337 VTAIL.n299 B 0.008411f
C338 VTAIL.n300 B 0.015652f
C339 VTAIL.n301 B 0.015652f
C340 VTAIL.n302 B 0.008411f
C341 VTAIL.n303 B 0.008905f
C342 VTAIL.n304 B 0.01988f
C343 VTAIL.n305 B 0.01988f
C344 VTAIL.n306 B 0.008905f
C345 VTAIL.n307 B 0.008411f
C346 VTAIL.n308 B 0.015652f
C347 VTAIL.n309 B 0.015652f
C348 VTAIL.n310 B 0.008411f
C349 VTAIL.n311 B 0.008905f
C350 VTAIL.n312 B 0.01988f
C351 VTAIL.n313 B 0.01988f
C352 VTAIL.n314 B 0.008905f
C353 VTAIL.n315 B 0.008411f
C354 VTAIL.n316 B 0.015652f
C355 VTAIL.n317 B 0.015652f
C356 VTAIL.n318 B 0.008411f
C357 VTAIL.n319 B 0.008658f
C358 VTAIL.n320 B 0.008658f
C359 VTAIL.n321 B 0.01988f
C360 VTAIL.n322 B 0.040796f
C361 VTAIL.n323 B 0.008905f
C362 VTAIL.n324 B 0.008411f
C363 VTAIL.n325 B 0.037889f
C364 VTAIL.n326 B 0.022648f
C365 VTAIL.n327 B 1.08607f
C366 VTAIL.n328 B 0.020733f
C367 VTAIL.n329 B 0.015652f
C368 VTAIL.n330 B 0.008411f
C369 VTAIL.n331 B 0.01988f
C370 VTAIL.n332 B 0.008905f
C371 VTAIL.n333 B 0.015652f
C372 VTAIL.n334 B 0.008411f
C373 VTAIL.n335 B 0.01988f
C374 VTAIL.n336 B 0.01988f
C375 VTAIL.n337 B 0.008905f
C376 VTAIL.n338 B 0.015652f
C377 VTAIL.n339 B 0.008411f
C378 VTAIL.n340 B 0.01988f
C379 VTAIL.n341 B 0.008905f
C380 VTAIL.n342 B 0.015652f
C381 VTAIL.n343 B 0.008411f
C382 VTAIL.n344 B 0.01988f
C383 VTAIL.n345 B 0.008905f
C384 VTAIL.n346 B 0.015652f
C385 VTAIL.n347 B 0.008411f
C386 VTAIL.n348 B 0.01988f
C387 VTAIL.n349 B 0.008905f
C388 VTAIL.n350 B 0.015652f
C389 VTAIL.n351 B 0.008411f
C390 VTAIL.n352 B 0.01988f
C391 VTAIL.n353 B 0.008905f
C392 VTAIL.n354 B 0.100987f
C393 VTAIL.t3 B 0.032764f
C394 VTAIL.n355 B 0.01491f
C395 VTAIL.n356 B 0.011744f
C396 VTAIL.n357 B 0.008411f
C397 VTAIL.n358 B 0.998259f
C398 VTAIL.n359 B 0.015652f
C399 VTAIL.n360 B 0.008411f
C400 VTAIL.n361 B 0.008905f
C401 VTAIL.n362 B 0.01988f
C402 VTAIL.n363 B 0.01988f
C403 VTAIL.n364 B 0.008905f
C404 VTAIL.n365 B 0.008411f
C405 VTAIL.n366 B 0.015652f
C406 VTAIL.n367 B 0.015652f
C407 VTAIL.n368 B 0.008411f
C408 VTAIL.n369 B 0.008905f
C409 VTAIL.n370 B 0.01988f
C410 VTAIL.n371 B 0.01988f
C411 VTAIL.n372 B 0.008905f
C412 VTAIL.n373 B 0.008411f
C413 VTAIL.n374 B 0.015652f
C414 VTAIL.n375 B 0.015652f
C415 VTAIL.n376 B 0.008411f
C416 VTAIL.n377 B 0.008905f
C417 VTAIL.n378 B 0.01988f
C418 VTAIL.n379 B 0.01988f
C419 VTAIL.n380 B 0.008905f
C420 VTAIL.n381 B 0.008411f
C421 VTAIL.n382 B 0.015652f
C422 VTAIL.n383 B 0.015652f
C423 VTAIL.n384 B 0.008411f
C424 VTAIL.n385 B 0.008905f
C425 VTAIL.n386 B 0.01988f
C426 VTAIL.n387 B 0.01988f
C427 VTAIL.n388 B 0.008905f
C428 VTAIL.n389 B 0.008411f
C429 VTAIL.n390 B 0.015652f
C430 VTAIL.n391 B 0.015652f
C431 VTAIL.n392 B 0.008411f
C432 VTAIL.n393 B 0.008905f
C433 VTAIL.n394 B 0.01988f
C434 VTAIL.n395 B 0.01988f
C435 VTAIL.n396 B 0.008905f
C436 VTAIL.n397 B 0.008411f
C437 VTAIL.n398 B 0.015652f
C438 VTAIL.n399 B 0.015652f
C439 VTAIL.n400 B 0.008411f
C440 VTAIL.n401 B 0.008658f
C441 VTAIL.n402 B 0.008658f
C442 VTAIL.n403 B 0.01988f
C443 VTAIL.n404 B 0.040796f
C444 VTAIL.n405 B 0.008905f
C445 VTAIL.n406 B 0.008411f
C446 VTAIL.n407 B 0.037889f
C447 VTAIL.n408 B 0.022648f
C448 VTAIL.n409 B 0.147594f
C449 VTAIL.n410 B 0.020733f
C450 VTAIL.n411 B 0.015652f
C451 VTAIL.n412 B 0.008411f
C452 VTAIL.n413 B 0.01988f
C453 VTAIL.n414 B 0.008905f
C454 VTAIL.n415 B 0.015652f
C455 VTAIL.n416 B 0.008411f
C456 VTAIL.n417 B 0.01988f
C457 VTAIL.n418 B 0.01988f
C458 VTAIL.n419 B 0.008905f
C459 VTAIL.n420 B 0.015652f
C460 VTAIL.n421 B 0.008411f
C461 VTAIL.n422 B 0.01988f
C462 VTAIL.n423 B 0.008905f
C463 VTAIL.n424 B 0.015652f
C464 VTAIL.n425 B 0.008411f
C465 VTAIL.n426 B 0.01988f
C466 VTAIL.n427 B 0.008905f
C467 VTAIL.n428 B 0.015652f
C468 VTAIL.n429 B 0.008411f
C469 VTAIL.n430 B 0.01988f
C470 VTAIL.n431 B 0.008905f
C471 VTAIL.n432 B 0.015652f
C472 VTAIL.n433 B 0.008411f
C473 VTAIL.n434 B 0.01988f
C474 VTAIL.n435 B 0.008905f
C475 VTAIL.n436 B 0.100987f
C476 VTAIL.t6 B 0.032764f
C477 VTAIL.n437 B 0.01491f
C478 VTAIL.n438 B 0.011744f
C479 VTAIL.n439 B 0.008411f
C480 VTAIL.n440 B 0.998259f
C481 VTAIL.n441 B 0.015652f
C482 VTAIL.n442 B 0.008411f
C483 VTAIL.n443 B 0.008905f
C484 VTAIL.n444 B 0.01988f
C485 VTAIL.n445 B 0.01988f
C486 VTAIL.n446 B 0.008905f
C487 VTAIL.n447 B 0.008411f
C488 VTAIL.n448 B 0.015652f
C489 VTAIL.n449 B 0.015652f
C490 VTAIL.n450 B 0.008411f
C491 VTAIL.n451 B 0.008905f
C492 VTAIL.n452 B 0.01988f
C493 VTAIL.n453 B 0.01988f
C494 VTAIL.n454 B 0.008905f
C495 VTAIL.n455 B 0.008411f
C496 VTAIL.n456 B 0.015652f
C497 VTAIL.n457 B 0.015652f
C498 VTAIL.n458 B 0.008411f
C499 VTAIL.n459 B 0.008905f
C500 VTAIL.n460 B 0.01988f
C501 VTAIL.n461 B 0.01988f
C502 VTAIL.n462 B 0.008905f
C503 VTAIL.n463 B 0.008411f
C504 VTAIL.n464 B 0.015652f
C505 VTAIL.n465 B 0.015652f
C506 VTAIL.n466 B 0.008411f
C507 VTAIL.n467 B 0.008905f
C508 VTAIL.n468 B 0.01988f
C509 VTAIL.n469 B 0.01988f
C510 VTAIL.n470 B 0.008905f
C511 VTAIL.n471 B 0.008411f
C512 VTAIL.n472 B 0.015652f
C513 VTAIL.n473 B 0.015652f
C514 VTAIL.n474 B 0.008411f
C515 VTAIL.n475 B 0.008905f
C516 VTAIL.n476 B 0.01988f
C517 VTAIL.n477 B 0.01988f
C518 VTAIL.n478 B 0.008905f
C519 VTAIL.n479 B 0.008411f
C520 VTAIL.n480 B 0.015652f
C521 VTAIL.n481 B 0.015652f
C522 VTAIL.n482 B 0.008411f
C523 VTAIL.n483 B 0.008658f
C524 VTAIL.n484 B 0.008658f
C525 VTAIL.n485 B 0.01988f
C526 VTAIL.n486 B 0.040796f
C527 VTAIL.n487 B 0.008905f
C528 VTAIL.n488 B 0.008411f
C529 VTAIL.n489 B 0.037889f
C530 VTAIL.n490 B 0.022648f
C531 VTAIL.n491 B 0.147594f
C532 VTAIL.n492 B 0.020733f
C533 VTAIL.n493 B 0.015652f
C534 VTAIL.n494 B 0.008411f
C535 VTAIL.n495 B 0.01988f
C536 VTAIL.n496 B 0.008905f
C537 VTAIL.n497 B 0.015652f
C538 VTAIL.n498 B 0.008411f
C539 VTAIL.n499 B 0.01988f
C540 VTAIL.n500 B 0.01988f
C541 VTAIL.n501 B 0.008905f
C542 VTAIL.n502 B 0.015652f
C543 VTAIL.n503 B 0.008411f
C544 VTAIL.n504 B 0.01988f
C545 VTAIL.n505 B 0.008905f
C546 VTAIL.n506 B 0.015652f
C547 VTAIL.n507 B 0.008411f
C548 VTAIL.n508 B 0.01988f
C549 VTAIL.n509 B 0.008905f
C550 VTAIL.n510 B 0.015652f
C551 VTAIL.n511 B 0.008411f
C552 VTAIL.n512 B 0.01988f
C553 VTAIL.n513 B 0.008905f
C554 VTAIL.n514 B 0.015652f
C555 VTAIL.n515 B 0.008411f
C556 VTAIL.n516 B 0.01988f
C557 VTAIL.n517 B 0.008905f
C558 VTAIL.n518 B 0.100987f
C559 VTAIL.t7 B 0.032764f
C560 VTAIL.n519 B 0.01491f
C561 VTAIL.n520 B 0.011744f
C562 VTAIL.n521 B 0.008411f
C563 VTAIL.n522 B 0.998259f
C564 VTAIL.n523 B 0.015652f
C565 VTAIL.n524 B 0.008411f
C566 VTAIL.n525 B 0.008905f
C567 VTAIL.n526 B 0.01988f
C568 VTAIL.n527 B 0.01988f
C569 VTAIL.n528 B 0.008905f
C570 VTAIL.n529 B 0.008411f
C571 VTAIL.n530 B 0.015652f
C572 VTAIL.n531 B 0.015652f
C573 VTAIL.n532 B 0.008411f
C574 VTAIL.n533 B 0.008905f
C575 VTAIL.n534 B 0.01988f
C576 VTAIL.n535 B 0.01988f
C577 VTAIL.n536 B 0.008905f
C578 VTAIL.n537 B 0.008411f
C579 VTAIL.n538 B 0.015652f
C580 VTAIL.n539 B 0.015652f
C581 VTAIL.n540 B 0.008411f
C582 VTAIL.n541 B 0.008905f
C583 VTAIL.n542 B 0.01988f
C584 VTAIL.n543 B 0.01988f
C585 VTAIL.n544 B 0.008905f
C586 VTAIL.n545 B 0.008411f
C587 VTAIL.n546 B 0.015652f
C588 VTAIL.n547 B 0.015652f
C589 VTAIL.n548 B 0.008411f
C590 VTAIL.n549 B 0.008905f
C591 VTAIL.n550 B 0.01988f
C592 VTAIL.n551 B 0.01988f
C593 VTAIL.n552 B 0.008905f
C594 VTAIL.n553 B 0.008411f
C595 VTAIL.n554 B 0.015652f
C596 VTAIL.n555 B 0.015652f
C597 VTAIL.n556 B 0.008411f
C598 VTAIL.n557 B 0.008905f
C599 VTAIL.n558 B 0.01988f
C600 VTAIL.n559 B 0.01988f
C601 VTAIL.n560 B 0.008905f
C602 VTAIL.n561 B 0.008411f
C603 VTAIL.n562 B 0.015652f
C604 VTAIL.n563 B 0.015652f
C605 VTAIL.n564 B 0.008411f
C606 VTAIL.n565 B 0.008658f
C607 VTAIL.n566 B 0.008658f
C608 VTAIL.n567 B 0.01988f
C609 VTAIL.n568 B 0.040796f
C610 VTAIL.n569 B 0.008905f
C611 VTAIL.n570 B 0.008411f
C612 VTAIL.n571 B 0.037889f
C613 VTAIL.n572 B 0.022648f
C614 VTAIL.n573 B 1.08607f
C615 VTAIL.n574 B 0.020733f
C616 VTAIL.n575 B 0.015652f
C617 VTAIL.n576 B 0.008411f
C618 VTAIL.n577 B 0.01988f
C619 VTAIL.n578 B 0.008905f
C620 VTAIL.n579 B 0.015652f
C621 VTAIL.n580 B 0.008411f
C622 VTAIL.n581 B 0.01988f
C623 VTAIL.n582 B 0.008905f
C624 VTAIL.n583 B 0.015652f
C625 VTAIL.n584 B 0.008411f
C626 VTAIL.n585 B 0.01988f
C627 VTAIL.n586 B 0.008905f
C628 VTAIL.n587 B 0.015652f
C629 VTAIL.n588 B 0.008411f
C630 VTAIL.n589 B 0.01988f
C631 VTAIL.n590 B 0.008905f
C632 VTAIL.n591 B 0.015652f
C633 VTAIL.n592 B 0.008411f
C634 VTAIL.n593 B 0.01988f
C635 VTAIL.n594 B 0.008905f
C636 VTAIL.n595 B 0.015652f
C637 VTAIL.n596 B 0.008411f
C638 VTAIL.n597 B 0.01988f
C639 VTAIL.n598 B 0.008905f
C640 VTAIL.n599 B 0.100987f
C641 VTAIL.t1 B 0.032764f
C642 VTAIL.n600 B 0.01491f
C643 VTAIL.n601 B 0.011744f
C644 VTAIL.n602 B 0.008411f
C645 VTAIL.n603 B 0.998259f
C646 VTAIL.n604 B 0.015652f
C647 VTAIL.n605 B 0.008411f
C648 VTAIL.n606 B 0.008905f
C649 VTAIL.n607 B 0.01988f
C650 VTAIL.n608 B 0.01988f
C651 VTAIL.n609 B 0.008905f
C652 VTAIL.n610 B 0.008411f
C653 VTAIL.n611 B 0.015652f
C654 VTAIL.n612 B 0.015652f
C655 VTAIL.n613 B 0.008411f
C656 VTAIL.n614 B 0.008905f
C657 VTAIL.n615 B 0.01988f
C658 VTAIL.n616 B 0.01988f
C659 VTAIL.n617 B 0.008905f
C660 VTAIL.n618 B 0.008411f
C661 VTAIL.n619 B 0.015652f
C662 VTAIL.n620 B 0.015652f
C663 VTAIL.n621 B 0.008411f
C664 VTAIL.n622 B 0.008905f
C665 VTAIL.n623 B 0.01988f
C666 VTAIL.n624 B 0.01988f
C667 VTAIL.n625 B 0.008905f
C668 VTAIL.n626 B 0.008411f
C669 VTAIL.n627 B 0.015652f
C670 VTAIL.n628 B 0.015652f
C671 VTAIL.n629 B 0.008411f
C672 VTAIL.n630 B 0.008905f
C673 VTAIL.n631 B 0.01988f
C674 VTAIL.n632 B 0.01988f
C675 VTAIL.n633 B 0.008905f
C676 VTAIL.n634 B 0.008411f
C677 VTAIL.n635 B 0.015652f
C678 VTAIL.n636 B 0.015652f
C679 VTAIL.n637 B 0.008411f
C680 VTAIL.n638 B 0.008905f
C681 VTAIL.n639 B 0.01988f
C682 VTAIL.n640 B 0.01988f
C683 VTAIL.n641 B 0.01988f
C684 VTAIL.n642 B 0.008905f
C685 VTAIL.n643 B 0.008411f
C686 VTAIL.n644 B 0.015652f
C687 VTAIL.n645 B 0.015652f
C688 VTAIL.n646 B 0.008411f
C689 VTAIL.n647 B 0.008658f
C690 VTAIL.n648 B 0.008658f
C691 VTAIL.n649 B 0.01988f
C692 VTAIL.n650 B 0.040796f
C693 VTAIL.n651 B 0.008905f
C694 VTAIL.n652 B 0.008411f
C695 VTAIL.n653 B 0.037889f
C696 VTAIL.n654 B 0.022648f
C697 VTAIL.n655 B 1.02836f
C698 VP.n0 B 0.037042f
C699 VP.t1 B 2.48092f
C700 VP.n1 B 0.022693f
C701 VP.n2 B 0.037042f
C702 VP.t2 B 2.48092f
C703 VP.t0 B 2.66333f
C704 VP.t3 B 2.66663f
C705 VP.n3 B 3.23202f
C706 VP.n4 B 1.62618f
C707 VP.n5 B 0.953944f
C708 VP.n6 B 0.039757f
C709 VP.n7 B 0.055549f
C710 VP.n8 B 0.028097f
C711 VP.n9 B 0.028097f
C712 VP.n10 B 0.028097f
C713 VP.n11 B 0.055549f
C714 VP.n12 B 0.039757f
C715 VP.n13 B 0.953944f
C716 VP.n14 B 0.040439f
.ends

