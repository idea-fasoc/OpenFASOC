* NGSPICE file created from diff_pair_sample_1195.ext - technology: sky130A

.subckt diff_pair_sample_1195 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=0 ps=0 w=11.46 l=3.23
X1 B.t8 B.t6 B.t7 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=0 ps=0 w=11.46 l=3.23
X2 VDD2.t5 VN.t0 VTAIL.t11 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=4.4694 ps=23.7 w=11.46 l=3.23
X3 VTAIL.t7 VN.t1 VDD2.t4 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=1.8909 ps=11.79 w=11.46 l=3.23
X4 VTAIL.t8 VN.t2 VDD2.t3 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=1.8909 ps=11.79 w=11.46 l=3.23
X5 VDD1.t5 VP.t0 VTAIL.t3 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=4.4694 ps=23.7 w=11.46 l=3.23
X6 VTAIL.t2 VP.t1 VDD1.t4 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=1.8909 ps=11.79 w=11.46 l=3.23
X7 VTAIL.t4 VP.t2 VDD1.t3 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=1.8909 ps=11.79 w=11.46 l=3.23
X8 VDD2.t2 VN.t3 VTAIL.t6 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=1.8909 ps=11.79 w=11.46 l=3.23
X9 VDD1.t2 VP.t3 VTAIL.t1 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=1.8909 ps=11.79 w=11.46 l=3.23
X10 B.t5 B.t3 B.t4 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=0 ps=0 w=11.46 l=3.23
X11 B.t2 B.t0 B.t1 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=0 ps=0 w=11.46 l=3.23
X12 VDD1.t1 VP.t4 VTAIL.t5 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=1.8909 ps=11.79 w=11.46 l=3.23
X13 VDD2.t1 VN.t4 VTAIL.t9 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=4.4694 ps=23.7 w=11.46 l=3.23
X14 VDD2.t0 VN.t5 VTAIL.t10 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=4.4694 pd=23.7 as=1.8909 ps=11.79 w=11.46 l=3.23
X15 VDD1.t0 VP.t5 VTAIL.t0 w_n3818_n3260# sky130_fd_pr__pfet_01v8 ad=1.8909 pd=11.79 as=4.4694 ps=23.7 w=11.46 l=3.23
R0 B.n563 B.n76 585
R1 B.n565 B.n564 585
R2 B.n566 B.n75 585
R3 B.n568 B.n567 585
R4 B.n569 B.n74 585
R5 B.n571 B.n570 585
R6 B.n572 B.n73 585
R7 B.n574 B.n573 585
R8 B.n575 B.n72 585
R9 B.n577 B.n576 585
R10 B.n578 B.n71 585
R11 B.n580 B.n579 585
R12 B.n581 B.n70 585
R13 B.n583 B.n582 585
R14 B.n584 B.n69 585
R15 B.n586 B.n585 585
R16 B.n587 B.n68 585
R17 B.n589 B.n588 585
R18 B.n590 B.n67 585
R19 B.n592 B.n591 585
R20 B.n593 B.n66 585
R21 B.n595 B.n594 585
R22 B.n596 B.n65 585
R23 B.n598 B.n597 585
R24 B.n599 B.n64 585
R25 B.n601 B.n600 585
R26 B.n602 B.n63 585
R27 B.n604 B.n603 585
R28 B.n605 B.n62 585
R29 B.n607 B.n606 585
R30 B.n608 B.n61 585
R31 B.n610 B.n609 585
R32 B.n611 B.n60 585
R33 B.n613 B.n612 585
R34 B.n614 B.n59 585
R35 B.n616 B.n615 585
R36 B.n617 B.n58 585
R37 B.n619 B.n618 585
R38 B.n620 B.n57 585
R39 B.n622 B.n621 585
R40 B.n624 B.n623 585
R41 B.n625 B.n53 585
R42 B.n627 B.n626 585
R43 B.n628 B.n52 585
R44 B.n630 B.n629 585
R45 B.n631 B.n51 585
R46 B.n633 B.n632 585
R47 B.n634 B.n50 585
R48 B.n636 B.n635 585
R49 B.n637 B.n47 585
R50 B.n640 B.n639 585
R51 B.n641 B.n46 585
R52 B.n643 B.n642 585
R53 B.n644 B.n45 585
R54 B.n646 B.n645 585
R55 B.n647 B.n44 585
R56 B.n649 B.n648 585
R57 B.n650 B.n43 585
R58 B.n652 B.n651 585
R59 B.n653 B.n42 585
R60 B.n655 B.n654 585
R61 B.n656 B.n41 585
R62 B.n658 B.n657 585
R63 B.n659 B.n40 585
R64 B.n661 B.n660 585
R65 B.n662 B.n39 585
R66 B.n664 B.n663 585
R67 B.n665 B.n38 585
R68 B.n667 B.n666 585
R69 B.n668 B.n37 585
R70 B.n670 B.n669 585
R71 B.n671 B.n36 585
R72 B.n673 B.n672 585
R73 B.n674 B.n35 585
R74 B.n676 B.n675 585
R75 B.n677 B.n34 585
R76 B.n679 B.n678 585
R77 B.n680 B.n33 585
R78 B.n682 B.n681 585
R79 B.n683 B.n32 585
R80 B.n685 B.n684 585
R81 B.n686 B.n31 585
R82 B.n688 B.n687 585
R83 B.n689 B.n30 585
R84 B.n691 B.n690 585
R85 B.n692 B.n29 585
R86 B.n694 B.n693 585
R87 B.n695 B.n28 585
R88 B.n697 B.n696 585
R89 B.n698 B.n27 585
R90 B.n562 B.n561 585
R91 B.n560 B.n77 585
R92 B.n559 B.n558 585
R93 B.n557 B.n78 585
R94 B.n556 B.n555 585
R95 B.n554 B.n79 585
R96 B.n553 B.n552 585
R97 B.n551 B.n80 585
R98 B.n550 B.n549 585
R99 B.n548 B.n81 585
R100 B.n547 B.n546 585
R101 B.n545 B.n82 585
R102 B.n544 B.n543 585
R103 B.n542 B.n83 585
R104 B.n541 B.n540 585
R105 B.n539 B.n84 585
R106 B.n538 B.n537 585
R107 B.n536 B.n85 585
R108 B.n535 B.n534 585
R109 B.n533 B.n86 585
R110 B.n532 B.n531 585
R111 B.n530 B.n87 585
R112 B.n529 B.n528 585
R113 B.n527 B.n88 585
R114 B.n526 B.n525 585
R115 B.n524 B.n89 585
R116 B.n523 B.n522 585
R117 B.n521 B.n90 585
R118 B.n520 B.n519 585
R119 B.n518 B.n91 585
R120 B.n517 B.n516 585
R121 B.n515 B.n92 585
R122 B.n514 B.n513 585
R123 B.n512 B.n93 585
R124 B.n511 B.n510 585
R125 B.n509 B.n94 585
R126 B.n508 B.n507 585
R127 B.n506 B.n95 585
R128 B.n505 B.n504 585
R129 B.n503 B.n96 585
R130 B.n502 B.n501 585
R131 B.n500 B.n97 585
R132 B.n499 B.n498 585
R133 B.n497 B.n98 585
R134 B.n496 B.n495 585
R135 B.n494 B.n99 585
R136 B.n493 B.n492 585
R137 B.n491 B.n100 585
R138 B.n490 B.n489 585
R139 B.n488 B.n101 585
R140 B.n487 B.n486 585
R141 B.n485 B.n102 585
R142 B.n484 B.n483 585
R143 B.n482 B.n103 585
R144 B.n481 B.n480 585
R145 B.n479 B.n104 585
R146 B.n478 B.n477 585
R147 B.n476 B.n105 585
R148 B.n475 B.n474 585
R149 B.n473 B.n106 585
R150 B.n472 B.n471 585
R151 B.n470 B.n107 585
R152 B.n469 B.n468 585
R153 B.n467 B.n108 585
R154 B.n466 B.n465 585
R155 B.n464 B.n109 585
R156 B.n463 B.n462 585
R157 B.n461 B.n110 585
R158 B.n460 B.n459 585
R159 B.n458 B.n111 585
R160 B.n457 B.n456 585
R161 B.n455 B.n112 585
R162 B.n454 B.n453 585
R163 B.n452 B.n113 585
R164 B.n451 B.n450 585
R165 B.n449 B.n114 585
R166 B.n448 B.n447 585
R167 B.n446 B.n115 585
R168 B.n445 B.n444 585
R169 B.n443 B.n116 585
R170 B.n442 B.n441 585
R171 B.n440 B.n117 585
R172 B.n439 B.n438 585
R173 B.n437 B.n118 585
R174 B.n436 B.n435 585
R175 B.n434 B.n119 585
R176 B.n433 B.n432 585
R177 B.n431 B.n120 585
R178 B.n430 B.n429 585
R179 B.n428 B.n121 585
R180 B.n427 B.n426 585
R181 B.n425 B.n122 585
R182 B.n424 B.n423 585
R183 B.n422 B.n123 585
R184 B.n421 B.n420 585
R185 B.n419 B.n124 585
R186 B.n418 B.n417 585
R187 B.n416 B.n125 585
R188 B.n415 B.n414 585
R189 B.n413 B.n126 585
R190 B.n412 B.n411 585
R191 B.n275 B.n176 585
R192 B.n277 B.n276 585
R193 B.n278 B.n175 585
R194 B.n280 B.n279 585
R195 B.n281 B.n174 585
R196 B.n283 B.n282 585
R197 B.n284 B.n173 585
R198 B.n286 B.n285 585
R199 B.n287 B.n172 585
R200 B.n289 B.n288 585
R201 B.n290 B.n171 585
R202 B.n292 B.n291 585
R203 B.n293 B.n170 585
R204 B.n295 B.n294 585
R205 B.n296 B.n169 585
R206 B.n298 B.n297 585
R207 B.n299 B.n168 585
R208 B.n301 B.n300 585
R209 B.n302 B.n167 585
R210 B.n304 B.n303 585
R211 B.n305 B.n166 585
R212 B.n307 B.n306 585
R213 B.n308 B.n165 585
R214 B.n310 B.n309 585
R215 B.n311 B.n164 585
R216 B.n313 B.n312 585
R217 B.n314 B.n163 585
R218 B.n316 B.n315 585
R219 B.n317 B.n162 585
R220 B.n319 B.n318 585
R221 B.n320 B.n161 585
R222 B.n322 B.n321 585
R223 B.n323 B.n160 585
R224 B.n325 B.n324 585
R225 B.n326 B.n159 585
R226 B.n328 B.n327 585
R227 B.n329 B.n158 585
R228 B.n331 B.n330 585
R229 B.n332 B.n157 585
R230 B.n334 B.n333 585
R231 B.n336 B.n335 585
R232 B.n337 B.n153 585
R233 B.n339 B.n338 585
R234 B.n340 B.n152 585
R235 B.n342 B.n341 585
R236 B.n343 B.n151 585
R237 B.n345 B.n344 585
R238 B.n346 B.n150 585
R239 B.n348 B.n347 585
R240 B.n349 B.n147 585
R241 B.n352 B.n351 585
R242 B.n353 B.n146 585
R243 B.n355 B.n354 585
R244 B.n356 B.n145 585
R245 B.n358 B.n357 585
R246 B.n359 B.n144 585
R247 B.n361 B.n360 585
R248 B.n362 B.n143 585
R249 B.n364 B.n363 585
R250 B.n365 B.n142 585
R251 B.n367 B.n366 585
R252 B.n368 B.n141 585
R253 B.n370 B.n369 585
R254 B.n371 B.n140 585
R255 B.n373 B.n372 585
R256 B.n374 B.n139 585
R257 B.n376 B.n375 585
R258 B.n377 B.n138 585
R259 B.n379 B.n378 585
R260 B.n380 B.n137 585
R261 B.n382 B.n381 585
R262 B.n383 B.n136 585
R263 B.n385 B.n384 585
R264 B.n386 B.n135 585
R265 B.n388 B.n387 585
R266 B.n389 B.n134 585
R267 B.n391 B.n390 585
R268 B.n392 B.n133 585
R269 B.n394 B.n393 585
R270 B.n395 B.n132 585
R271 B.n397 B.n396 585
R272 B.n398 B.n131 585
R273 B.n400 B.n399 585
R274 B.n401 B.n130 585
R275 B.n403 B.n402 585
R276 B.n404 B.n129 585
R277 B.n406 B.n405 585
R278 B.n407 B.n128 585
R279 B.n409 B.n408 585
R280 B.n410 B.n127 585
R281 B.n274 B.n273 585
R282 B.n272 B.n177 585
R283 B.n271 B.n270 585
R284 B.n269 B.n178 585
R285 B.n268 B.n267 585
R286 B.n266 B.n179 585
R287 B.n265 B.n264 585
R288 B.n263 B.n180 585
R289 B.n262 B.n261 585
R290 B.n260 B.n181 585
R291 B.n259 B.n258 585
R292 B.n257 B.n182 585
R293 B.n256 B.n255 585
R294 B.n254 B.n183 585
R295 B.n253 B.n252 585
R296 B.n251 B.n184 585
R297 B.n250 B.n249 585
R298 B.n248 B.n185 585
R299 B.n247 B.n246 585
R300 B.n245 B.n186 585
R301 B.n244 B.n243 585
R302 B.n242 B.n187 585
R303 B.n241 B.n240 585
R304 B.n239 B.n188 585
R305 B.n238 B.n237 585
R306 B.n236 B.n189 585
R307 B.n235 B.n234 585
R308 B.n233 B.n190 585
R309 B.n232 B.n231 585
R310 B.n230 B.n191 585
R311 B.n229 B.n228 585
R312 B.n227 B.n192 585
R313 B.n226 B.n225 585
R314 B.n224 B.n193 585
R315 B.n223 B.n222 585
R316 B.n221 B.n194 585
R317 B.n220 B.n219 585
R318 B.n218 B.n195 585
R319 B.n217 B.n216 585
R320 B.n215 B.n196 585
R321 B.n214 B.n213 585
R322 B.n212 B.n197 585
R323 B.n211 B.n210 585
R324 B.n209 B.n198 585
R325 B.n208 B.n207 585
R326 B.n206 B.n199 585
R327 B.n205 B.n204 585
R328 B.n203 B.n200 585
R329 B.n202 B.n201 585
R330 B.n2 B.n0 585
R331 B.n773 B.n1 585
R332 B.n772 B.n771 585
R333 B.n770 B.n3 585
R334 B.n769 B.n768 585
R335 B.n767 B.n4 585
R336 B.n766 B.n765 585
R337 B.n764 B.n5 585
R338 B.n763 B.n762 585
R339 B.n761 B.n6 585
R340 B.n760 B.n759 585
R341 B.n758 B.n7 585
R342 B.n757 B.n756 585
R343 B.n755 B.n8 585
R344 B.n754 B.n753 585
R345 B.n752 B.n9 585
R346 B.n751 B.n750 585
R347 B.n749 B.n10 585
R348 B.n748 B.n747 585
R349 B.n746 B.n11 585
R350 B.n745 B.n744 585
R351 B.n743 B.n12 585
R352 B.n742 B.n741 585
R353 B.n740 B.n13 585
R354 B.n739 B.n738 585
R355 B.n737 B.n14 585
R356 B.n736 B.n735 585
R357 B.n734 B.n15 585
R358 B.n733 B.n732 585
R359 B.n731 B.n16 585
R360 B.n730 B.n729 585
R361 B.n728 B.n17 585
R362 B.n727 B.n726 585
R363 B.n725 B.n18 585
R364 B.n724 B.n723 585
R365 B.n722 B.n19 585
R366 B.n721 B.n720 585
R367 B.n719 B.n20 585
R368 B.n718 B.n717 585
R369 B.n716 B.n21 585
R370 B.n715 B.n714 585
R371 B.n713 B.n22 585
R372 B.n712 B.n711 585
R373 B.n710 B.n23 585
R374 B.n709 B.n708 585
R375 B.n707 B.n24 585
R376 B.n706 B.n705 585
R377 B.n704 B.n25 585
R378 B.n703 B.n702 585
R379 B.n701 B.n26 585
R380 B.n700 B.n699 585
R381 B.n775 B.n774 585
R382 B.n275 B.n274 468.476
R383 B.n700 B.n27 468.476
R384 B.n412 B.n127 468.476
R385 B.n563 B.n562 468.476
R386 B.n148 B.t11 435.041
R387 B.n54 B.t7 435.041
R388 B.n154 B.t2 435.041
R389 B.n48 B.t4 435.041
R390 B.n149 B.t10 366
R391 B.n55 B.t8 366
R392 B.n155 B.t1 366
R393 B.n49 B.t5 366
R394 B.n148 B.t9 294.341
R395 B.n154 B.t0 294.341
R396 B.n48 B.t3 294.341
R397 B.n54 B.t6 294.341
R398 B.n274 B.n177 163.367
R399 B.n270 B.n177 163.367
R400 B.n270 B.n269 163.367
R401 B.n269 B.n268 163.367
R402 B.n268 B.n179 163.367
R403 B.n264 B.n179 163.367
R404 B.n264 B.n263 163.367
R405 B.n263 B.n262 163.367
R406 B.n262 B.n181 163.367
R407 B.n258 B.n181 163.367
R408 B.n258 B.n257 163.367
R409 B.n257 B.n256 163.367
R410 B.n256 B.n183 163.367
R411 B.n252 B.n183 163.367
R412 B.n252 B.n251 163.367
R413 B.n251 B.n250 163.367
R414 B.n250 B.n185 163.367
R415 B.n246 B.n185 163.367
R416 B.n246 B.n245 163.367
R417 B.n245 B.n244 163.367
R418 B.n244 B.n187 163.367
R419 B.n240 B.n187 163.367
R420 B.n240 B.n239 163.367
R421 B.n239 B.n238 163.367
R422 B.n238 B.n189 163.367
R423 B.n234 B.n189 163.367
R424 B.n234 B.n233 163.367
R425 B.n233 B.n232 163.367
R426 B.n232 B.n191 163.367
R427 B.n228 B.n191 163.367
R428 B.n228 B.n227 163.367
R429 B.n227 B.n226 163.367
R430 B.n226 B.n193 163.367
R431 B.n222 B.n193 163.367
R432 B.n222 B.n221 163.367
R433 B.n221 B.n220 163.367
R434 B.n220 B.n195 163.367
R435 B.n216 B.n195 163.367
R436 B.n216 B.n215 163.367
R437 B.n215 B.n214 163.367
R438 B.n214 B.n197 163.367
R439 B.n210 B.n197 163.367
R440 B.n210 B.n209 163.367
R441 B.n209 B.n208 163.367
R442 B.n208 B.n199 163.367
R443 B.n204 B.n199 163.367
R444 B.n204 B.n203 163.367
R445 B.n203 B.n202 163.367
R446 B.n202 B.n2 163.367
R447 B.n774 B.n2 163.367
R448 B.n774 B.n773 163.367
R449 B.n773 B.n772 163.367
R450 B.n772 B.n3 163.367
R451 B.n768 B.n3 163.367
R452 B.n768 B.n767 163.367
R453 B.n767 B.n766 163.367
R454 B.n766 B.n5 163.367
R455 B.n762 B.n5 163.367
R456 B.n762 B.n761 163.367
R457 B.n761 B.n760 163.367
R458 B.n760 B.n7 163.367
R459 B.n756 B.n7 163.367
R460 B.n756 B.n755 163.367
R461 B.n755 B.n754 163.367
R462 B.n754 B.n9 163.367
R463 B.n750 B.n9 163.367
R464 B.n750 B.n749 163.367
R465 B.n749 B.n748 163.367
R466 B.n748 B.n11 163.367
R467 B.n744 B.n11 163.367
R468 B.n744 B.n743 163.367
R469 B.n743 B.n742 163.367
R470 B.n742 B.n13 163.367
R471 B.n738 B.n13 163.367
R472 B.n738 B.n737 163.367
R473 B.n737 B.n736 163.367
R474 B.n736 B.n15 163.367
R475 B.n732 B.n15 163.367
R476 B.n732 B.n731 163.367
R477 B.n731 B.n730 163.367
R478 B.n730 B.n17 163.367
R479 B.n726 B.n17 163.367
R480 B.n726 B.n725 163.367
R481 B.n725 B.n724 163.367
R482 B.n724 B.n19 163.367
R483 B.n720 B.n19 163.367
R484 B.n720 B.n719 163.367
R485 B.n719 B.n718 163.367
R486 B.n718 B.n21 163.367
R487 B.n714 B.n21 163.367
R488 B.n714 B.n713 163.367
R489 B.n713 B.n712 163.367
R490 B.n712 B.n23 163.367
R491 B.n708 B.n23 163.367
R492 B.n708 B.n707 163.367
R493 B.n707 B.n706 163.367
R494 B.n706 B.n25 163.367
R495 B.n702 B.n25 163.367
R496 B.n702 B.n701 163.367
R497 B.n701 B.n700 163.367
R498 B.n276 B.n275 163.367
R499 B.n276 B.n175 163.367
R500 B.n280 B.n175 163.367
R501 B.n281 B.n280 163.367
R502 B.n282 B.n281 163.367
R503 B.n282 B.n173 163.367
R504 B.n286 B.n173 163.367
R505 B.n287 B.n286 163.367
R506 B.n288 B.n287 163.367
R507 B.n288 B.n171 163.367
R508 B.n292 B.n171 163.367
R509 B.n293 B.n292 163.367
R510 B.n294 B.n293 163.367
R511 B.n294 B.n169 163.367
R512 B.n298 B.n169 163.367
R513 B.n299 B.n298 163.367
R514 B.n300 B.n299 163.367
R515 B.n300 B.n167 163.367
R516 B.n304 B.n167 163.367
R517 B.n305 B.n304 163.367
R518 B.n306 B.n305 163.367
R519 B.n306 B.n165 163.367
R520 B.n310 B.n165 163.367
R521 B.n311 B.n310 163.367
R522 B.n312 B.n311 163.367
R523 B.n312 B.n163 163.367
R524 B.n316 B.n163 163.367
R525 B.n317 B.n316 163.367
R526 B.n318 B.n317 163.367
R527 B.n318 B.n161 163.367
R528 B.n322 B.n161 163.367
R529 B.n323 B.n322 163.367
R530 B.n324 B.n323 163.367
R531 B.n324 B.n159 163.367
R532 B.n328 B.n159 163.367
R533 B.n329 B.n328 163.367
R534 B.n330 B.n329 163.367
R535 B.n330 B.n157 163.367
R536 B.n334 B.n157 163.367
R537 B.n335 B.n334 163.367
R538 B.n335 B.n153 163.367
R539 B.n339 B.n153 163.367
R540 B.n340 B.n339 163.367
R541 B.n341 B.n340 163.367
R542 B.n341 B.n151 163.367
R543 B.n345 B.n151 163.367
R544 B.n346 B.n345 163.367
R545 B.n347 B.n346 163.367
R546 B.n347 B.n147 163.367
R547 B.n352 B.n147 163.367
R548 B.n353 B.n352 163.367
R549 B.n354 B.n353 163.367
R550 B.n354 B.n145 163.367
R551 B.n358 B.n145 163.367
R552 B.n359 B.n358 163.367
R553 B.n360 B.n359 163.367
R554 B.n360 B.n143 163.367
R555 B.n364 B.n143 163.367
R556 B.n365 B.n364 163.367
R557 B.n366 B.n365 163.367
R558 B.n366 B.n141 163.367
R559 B.n370 B.n141 163.367
R560 B.n371 B.n370 163.367
R561 B.n372 B.n371 163.367
R562 B.n372 B.n139 163.367
R563 B.n376 B.n139 163.367
R564 B.n377 B.n376 163.367
R565 B.n378 B.n377 163.367
R566 B.n378 B.n137 163.367
R567 B.n382 B.n137 163.367
R568 B.n383 B.n382 163.367
R569 B.n384 B.n383 163.367
R570 B.n384 B.n135 163.367
R571 B.n388 B.n135 163.367
R572 B.n389 B.n388 163.367
R573 B.n390 B.n389 163.367
R574 B.n390 B.n133 163.367
R575 B.n394 B.n133 163.367
R576 B.n395 B.n394 163.367
R577 B.n396 B.n395 163.367
R578 B.n396 B.n131 163.367
R579 B.n400 B.n131 163.367
R580 B.n401 B.n400 163.367
R581 B.n402 B.n401 163.367
R582 B.n402 B.n129 163.367
R583 B.n406 B.n129 163.367
R584 B.n407 B.n406 163.367
R585 B.n408 B.n407 163.367
R586 B.n408 B.n127 163.367
R587 B.n413 B.n412 163.367
R588 B.n414 B.n413 163.367
R589 B.n414 B.n125 163.367
R590 B.n418 B.n125 163.367
R591 B.n419 B.n418 163.367
R592 B.n420 B.n419 163.367
R593 B.n420 B.n123 163.367
R594 B.n424 B.n123 163.367
R595 B.n425 B.n424 163.367
R596 B.n426 B.n425 163.367
R597 B.n426 B.n121 163.367
R598 B.n430 B.n121 163.367
R599 B.n431 B.n430 163.367
R600 B.n432 B.n431 163.367
R601 B.n432 B.n119 163.367
R602 B.n436 B.n119 163.367
R603 B.n437 B.n436 163.367
R604 B.n438 B.n437 163.367
R605 B.n438 B.n117 163.367
R606 B.n442 B.n117 163.367
R607 B.n443 B.n442 163.367
R608 B.n444 B.n443 163.367
R609 B.n444 B.n115 163.367
R610 B.n448 B.n115 163.367
R611 B.n449 B.n448 163.367
R612 B.n450 B.n449 163.367
R613 B.n450 B.n113 163.367
R614 B.n454 B.n113 163.367
R615 B.n455 B.n454 163.367
R616 B.n456 B.n455 163.367
R617 B.n456 B.n111 163.367
R618 B.n460 B.n111 163.367
R619 B.n461 B.n460 163.367
R620 B.n462 B.n461 163.367
R621 B.n462 B.n109 163.367
R622 B.n466 B.n109 163.367
R623 B.n467 B.n466 163.367
R624 B.n468 B.n467 163.367
R625 B.n468 B.n107 163.367
R626 B.n472 B.n107 163.367
R627 B.n473 B.n472 163.367
R628 B.n474 B.n473 163.367
R629 B.n474 B.n105 163.367
R630 B.n478 B.n105 163.367
R631 B.n479 B.n478 163.367
R632 B.n480 B.n479 163.367
R633 B.n480 B.n103 163.367
R634 B.n484 B.n103 163.367
R635 B.n485 B.n484 163.367
R636 B.n486 B.n485 163.367
R637 B.n486 B.n101 163.367
R638 B.n490 B.n101 163.367
R639 B.n491 B.n490 163.367
R640 B.n492 B.n491 163.367
R641 B.n492 B.n99 163.367
R642 B.n496 B.n99 163.367
R643 B.n497 B.n496 163.367
R644 B.n498 B.n497 163.367
R645 B.n498 B.n97 163.367
R646 B.n502 B.n97 163.367
R647 B.n503 B.n502 163.367
R648 B.n504 B.n503 163.367
R649 B.n504 B.n95 163.367
R650 B.n508 B.n95 163.367
R651 B.n509 B.n508 163.367
R652 B.n510 B.n509 163.367
R653 B.n510 B.n93 163.367
R654 B.n514 B.n93 163.367
R655 B.n515 B.n514 163.367
R656 B.n516 B.n515 163.367
R657 B.n516 B.n91 163.367
R658 B.n520 B.n91 163.367
R659 B.n521 B.n520 163.367
R660 B.n522 B.n521 163.367
R661 B.n522 B.n89 163.367
R662 B.n526 B.n89 163.367
R663 B.n527 B.n526 163.367
R664 B.n528 B.n527 163.367
R665 B.n528 B.n87 163.367
R666 B.n532 B.n87 163.367
R667 B.n533 B.n532 163.367
R668 B.n534 B.n533 163.367
R669 B.n534 B.n85 163.367
R670 B.n538 B.n85 163.367
R671 B.n539 B.n538 163.367
R672 B.n540 B.n539 163.367
R673 B.n540 B.n83 163.367
R674 B.n544 B.n83 163.367
R675 B.n545 B.n544 163.367
R676 B.n546 B.n545 163.367
R677 B.n546 B.n81 163.367
R678 B.n550 B.n81 163.367
R679 B.n551 B.n550 163.367
R680 B.n552 B.n551 163.367
R681 B.n552 B.n79 163.367
R682 B.n556 B.n79 163.367
R683 B.n557 B.n556 163.367
R684 B.n558 B.n557 163.367
R685 B.n558 B.n77 163.367
R686 B.n562 B.n77 163.367
R687 B.n696 B.n27 163.367
R688 B.n696 B.n695 163.367
R689 B.n695 B.n694 163.367
R690 B.n694 B.n29 163.367
R691 B.n690 B.n29 163.367
R692 B.n690 B.n689 163.367
R693 B.n689 B.n688 163.367
R694 B.n688 B.n31 163.367
R695 B.n684 B.n31 163.367
R696 B.n684 B.n683 163.367
R697 B.n683 B.n682 163.367
R698 B.n682 B.n33 163.367
R699 B.n678 B.n33 163.367
R700 B.n678 B.n677 163.367
R701 B.n677 B.n676 163.367
R702 B.n676 B.n35 163.367
R703 B.n672 B.n35 163.367
R704 B.n672 B.n671 163.367
R705 B.n671 B.n670 163.367
R706 B.n670 B.n37 163.367
R707 B.n666 B.n37 163.367
R708 B.n666 B.n665 163.367
R709 B.n665 B.n664 163.367
R710 B.n664 B.n39 163.367
R711 B.n660 B.n39 163.367
R712 B.n660 B.n659 163.367
R713 B.n659 B.n658 163.367
R714 B.n658 B.n41 163.367
R715 B.n654 B.n41 163.367
R716 B.n654 B.n653 163.367
R717 B.n653 B.n652 163.367
R718 B.n652 B.n43 163.367
R719 B.n648 B.n43 163.367
R720 B.n648 B.n647 163.367
R721 B.n647 B.n646 163.367
R722 B.n646 B.n45 163.367
R723 B.n642 B.n45 163.367
R724 B.n642 B.n641 163.367
R725 B.n641 B.n640 163.367
R726 B.n640 B.n47 163.367
R727 B.n635 B.n47 163.367
R728 B.n635 B.n634 163.367
R729 B.n634 B.n633 163.367
R730 B.n633 B.n51 163.367
R731 B.n629 B.n51 163.367
R732 B.n629 B.n628 163.367
R733 B.n628 B.n627 163.367
R734 B.n627 B.n53 163.367
R735 B.n623 B.n53 163.367
R736 B.n623 B.n622 163.367
R737 B.n622 B.n57 163.367
R738 B.n618 B.n57 163.367
R739 B.n618 B.n617 163.367
R740 B.n617 B.n616 163.367
R741 B.n616 B.n59 163.367
R742 B.n612 B.n59 163.367
R743 B.n612 B.n611 163.367
R744 B.n611 B.n610 163.367
R745 B.n610 B.n61 163.367
R746 B.n606 B.n61 163.367
R747 B.n606 B.n605 163.367
R748 B.n605 B.n604 163.367
R749 B.n604 B.n63 163.367
R750 B.n600 B.n63 163.367
R751 B.n600 B.n599 163.367
R752 B.n599 B.n598 163.367
R753 B.n598 B.n65 163.367
R754 B.n594 B.n65 163.367
R755 B.n594 B.n593 163.367
R756 B.n593 B.n592 163.367
R757 B.n592 B.n67 163.367
R758 B.n588 B.n67 163.367
R759 B.n588 B.n587 163.367
R760 B.n587 B.n586 163.367
R761 B.n586 B.n69 163.367
R762 B.n582 B.n69 163.367
R763 B.n582 B.n581 163.367
R764 B.n581 B.n580 163.367
R765 B.n580 B.n71 163.367
R766 B.n576 B.n71 163.367
R767 B.n576 B.n575 163.367
R768 B.n575 B.n574 163.367
R769 B.n574 B.n73 163.367
R770 B.n570 B.n73 163.367
R771 B.n570 B.n569 163.367
R772 B.n569 B.n568 163.367
R773 B.n568 B.n75 163.367
R774 B.n564 B.n75 163.367
R775 B.n564 B.n563 163.367
R776 B.n149 B.n148 69.0429
R777 B.n155 B.n154 69.0429
R778 B.n49 B.n48 69.0429
R779 B.n55 B.n54 69.0429
R780 B.n350 B.n149 59.5399
R781 B.n156 B.n155 59.5399
R782 B.n638 B.n49 59.5399
R783 B.n56 B.n55 59.5399
R784 B.n699 B.n698 30.4395
R785 B.n561 B.n76 30.4395
R786 B.n411 B.n410 30.4395
R787 B.n273 B.n176 30.4395
R788 B B.n775 18.0485
R789 B.n698 B.n697 10.6151
R790 B.n697 B.n28 10.6151
R791 B.n693 B.n28 10.6151
R792 B.n693 B.n692 10.6151
R793 B.n692 B.n691 10.6151
R794 B.n691 B.n30 10.6151
R795 B.n687 B.n30 10.6151
R796 B.n687 B.n686 10.6151
R797 B.n686 B.n685 10.6151
R798 B.n685 B.n32 10.6151
R799 B.n681 B.n32 10.6151
R800 B.n681 B.n680 10.6151
R801 B.n680 B.n679 10.6151
R802 B.n679 B.n34 10.6151
R803 B.n675 B.n34 10.6151
R804 B.n675 B.n674 10.6151
R805 B.n674 B.n673 10.6151
R806 B.n673 B.n36 10.6151
R807 B.n669 B.n36 10.6151
R808 B.n669 B.n668 10.6151
R809 B.n668 B.n667 10.6151
R810 B.n667 B.n38 10.6151
R811 B.n663 B.n38 10.6151
R812 B.n663 B.n662 10.6151
R813 B.n662 B.n661 10.6151
R814 B.n661 B.n40 10.6151
R815 B.n657 B.n40 10.6151
R816 B.n657 B.n656 10.6151
R817 B.n656 B.n655 10.6151
R818 B.n655 B.n42 10.6151
R819 B.n651 B.n42 10.6151
R820 B.n651 B.n650 10.6151
R821 B.n650 B.n649 10.6151
R822 B.n649 B.n44 10.6151
R823 B.n645 B.n44 10.6151
R824 B.n645 B.n644 10.6151
R825 B.n644 B.n643 10.6151
R826 B.n643 B.n46 10.6151
R827 B.n639 B.n46 10.6151
R828 B.n637 B.n636 10.6151
R829 B.n636 B.n50 10.6151
R830 B.n632 B.n50 10.6151
R831 B.n632 B.n631 10.6151
R832 B.n631 B.n630 10.6151
R833 B.n630 B.n52 10.6151
R834 B.n626 B.n52 10.6151
R835 B.n626 B.n625 10.6151
R836 B.n625 B.n624 10.6151
R837 B.n621 B.n620 10.6151
R838 B.n620 B.n619 10.6151
R839 B.n619 B.n58 10.6151
R840 B.n615 B.n58 10.6151
R841 B.n615 B.n614 10.6151
R842 B.n614 B.n613 10.6151
R843 B.n613 B.n60 10.6151
R844 B.n609 B.n60 10.6151
R845 B.n609 B.n608 10.6151
R846 B.n608 B.n607 10.6151
R847 B.n607 B.n62 10.6151
R848 B.n603 B.n62 10.6151
R849 B.n603 B.n602 10.6151
R850 B.n602 B.n601 10.6151
R851 B.n601 B.n64 10.6151
R852 B.n597 B.n64 10.6151
R853 B.n597 B.n596 10.6151
R854 B.n596 B.n595 10.6151
R855 B.n595 B.n66 10.6151
R856 B.n591 B.n66 10.6151
R857 B.n591 B.n590 10.6151
R858 B.n590 B.n589 10.6151
R859 B.n589 B.n68 10.6151
R860 B.n585 B.n68 10.6151
R861 B.n585 B.n584 10.6151
R862 B.n584 B.n583 10.6151
R863 B.n583 B.n70 10.6151
R864 B.n579 B.n70 10.6151
R865 B.n579 B.n578 10.6151
R866 B.n578 B.n577 10.6151
R867 B.n577 B.n72 10.6151
R868 B.n573 B.n72 10.6151
R869 B.n573 B.n572 10.6151
R870 B.n572 B.n571 10.6151
R871 B.n571 B.n74 10.6151
R872 B.n567 B.n74 10.6151
R873 B.n567 B.n566 10.6151
R874 B.n566 B.n565 10.6151
R875 B.n565 B.n76 10.6151
R876 B.n411 B.n126 10.6151
R877 B.n415 B.n126 10.6151
R878 B.n416 B.n415 10.6151
R879 B.n417 B.n416 10.6151
R880 B.n417 B.n124 10.6151
R881 B.n421 B.n124 10.6151
R882 B.n422 B.n421 10.6151
R883 B.n423 B.n422 10.6151
R884 B.n423 B.n122 10.6151
R885 B.n427 B.n122 10.6151
R886 B.n428 B.n427 10.6151
R887 B.n429 B.n428 10.6151
R888 B.n429 B.n120 10.6151
R889 B.n433 B.n120 10.6151
R890 B.n434 B.n433 10.6151
R891 B.n435 B.n434 10.6151
R892 B.n435 B.n118 10.6151
R893 B.n439 B.n118 10.6151
R894 B.n440 B.n439 10.6151
R895 B.n441 B.n440 10.6151
R896 B.n441 B.n116 10.6151
R897 B.n445 B.n116 10.6151
R898 B.n446 B.n445 10.6151
R899 B.n447 B.n446 10.6151
R900 B.n447 B.n114 10.6151
R901 B.n451 B.n114 10.6151
R902 B.n452 B.n451 10.6151
R903 B.n453 B.n452 10.6151
R904 B.n453 B.n112 10.6151
R905 B.n457 B.n112 10.6151
R906 B.n458 B.n457 10.6151
R907 B.n459 B.n458 10.6151
R908 B.n459 B.n110 10.6151
R909 B.n463 B.n110 10.6151
R910 B.n464 B.n463 10.6151
R911 B.n465 B.n464 10.6151
R912 B.n465 B.n108 10.6151
R913 B.n469 B.n108 10.6151
R914 B.n470 B.n469 10.6151
R915 B.n471 B.n470 10.6151
R916 B.n471 B.n106 10.6151
R917 B.n475 B.n106 10.6151
R918 B.n476 B.n475 10.6151
R919 B.n477 B.n476 10.6151
R920 B.n477 B.n104 10.6151
R921 B.n481 B.n104 10.6151
R922 B.n482 B.n481 10.6151
R923 B.n483 B.n482 10.6151
R924 B.n483 B.n102 10.6151
R925 B.n487 B.n102 10.6151
R926 B.n488 B.n487 10.6151
R927 B.n489 B.n488 10.6151
R928 B.n489 B.n100 10.6151
R929 B.n493 B.n100 10.6151
R930 B.n494 B.n493 10.6151
R931 B.n495 B.n494 10.6151
R932 B.n495 B.n98 10.6151
R933 B.n499 B.n98 10.6151
R934 B.n500 B.n499 10.6151
R935 B.n501 B.n500 10.6151
R936 B.n501 B.n96 10.6151
R937 B.n505 B.n96 10.6151
R938 B.n506 B.n505 10.6151
R939 B.n507 B.n506 10.6151
R940 B.n507 B.n94 10.6151
R941 B.n511 B.n94 10.6151
R942 B.n512 B.n511 10.6151
R943 B.n513 B.n512 10.6151
R944 B.n513 B.n92 10.6151
R945 B.n517 B.n92 10.6151
R946 B.n518 B.n517 10.6151
R947 B.n519 B.n518 10.6151
R948 B.n519 B.n90 10.6151
R949 B.n523 B.n90 10.6151
R950 B.n524 B.n523 10.6151
R951 B.n525 B.n524 10.6151
R952 B.n525 B.n88 10.6151
R953 B.n529 B.n88 10.6151
R954 B.n530 B.n529 10.6151
R955 B.n531 B.n530 10.6151
R956 B.n531 B.n86 10.6151
R957 B.n535 B.n86 10.6151
R958 B.n536 B.n535 10.6151
R959 B.n537 B.n536 10.6151
R960 B.n537 B.n84 10.6151
R961 B.n541 B.n84 10.6151
R962 B.n542 B.n541 10.6151
R963 B.n543 B.n542 10.6151
R964 B.n543 B.n82 10.6151
R965 B.n547 B.n82 10.6151
R966 B.n548 B.n547 10.6151
R967 B.n549 B.n548 10.6151
R968 B.n549 B.n80 10.6151
R969 B.n553 B.n80 10.6151
R970 B.n554 B.n553 10.6151
R971 B.n555 B.n554 10.6151
R972 B.n555 B.n78 10.6151
R973 B.n559 B.n78 10.6151
R974 B.n560 B.n559 10.6151
R975 B.n561 B.n560 10.6151
R976 B.n277 B.n176 10.6151
R977 B.n278 B.n277 10.6151
R978 B.n279 B.n278 10.6151
R979 B.n279 B.n174 10.6151
R980 B.n283 B.n174 10.6151
R981 B.n284 B.n283 10.6151
R982 B.n285 B.n284 10.6151
R983 B.n285 B.n172 10.6151
R984 B.n289 B.n172 10.6151
R985 B.n290 B.n289 10.6151
R986 B.n291 B.n290 10.6151
R987 B.n291 B.n170 10.6151
R988 B.n295 B.n170 10.6151
R989 B.n296 B.n295 10.6151
R990 B.n297 B.n296 10.6151
R991 B.n297 B.n168 10.6151
R992 B.n301 B.n168 10.6151
R993 B.n302 B.n301 10.6151
R994 B.n303 B.n302 10.6151
R995 B.n303 B.n166 10.6151
R996 B.n307 B.n166 10.6151
R997 B.n308 B.n307 10.6151
R998 B.n309 B.n308 10.6151
R999 B.n309 B.n164 10.6151
R1000 B.n313 B.n164 10.6151
R1001 B.n314 B.n313 10.6151
R1002 B.n315 B.n314 10.6151
R1003 B.n315 B.n162 10.6151
R1004 B.n319 B.n162 10.6151
R1005 B.n320 B.n319 10.6151
R1006 B.n321 B.n320 10.6151
R1007 B.n321 B.n160 10.6151
R1008 B.n325 B.n160 10.6151
R1009 B.n326 B.n325 10.6151
R1010 B.n327 B.n326 10.6151
R1011 B.n327 B.n158 10.6151
R1012 B.n331 B.n158 10.6151
R1013 B.n332 B.n331 10.6151
R1014 B.n333 B.n332 10.6151
R1015 B.n337 B.n336 10.6151
R1016 B.n338 B.n337 10.6151
R1017 B.n338 B.n152 10.6151
R1018 B.n342 B.n152 10.6151
R1019 B.n343 B.n342 10.6151
R1020 B.n344 B.n343 10.6151
R1021 B.n344 B.n150 10.6151
R1022 B.n348 B.n150 10.6151
R1023 B.n349 B.n348 10.6151
R1024 B.n351 B.n146 10.6151
R1025 B.n355 B.n146 10.6151
R1026 B.n356 B.n355 10.6151
R1027 B.n357 B.n356 10.6151
R1028 B.n357 B.n144 10.6151
R1029 B.n361 B.n144 10.6151
R1030 B.n362 B.n361 10.6151
R1031 B.n363 B.n362 10.6151
R1032 B.n363 B.n142 10.6151
R1033 B.n367 B.n142 10.6151
R1034 B.n368 B.n367 10.6151
R1035 B.n369 B.n368 10.6151
R1036 B.n369 B.n140 10.6151
R1037 B.n373 B.n140 10.6151
R1038 B.n374 B.n373 10.6151
R1039 B.n375 B.n374 10.6151
R1040 B.n375 B.n138 10.6151
R1041 B.n379 B.n138 10.6151
R1042 B.n380 B.n379 10.6151
R1043 B.n381 B.n380 10.6151
R1044 B.n381 B.n136 10.6151
R1045 B.n385 B.n136 10.6151
R1046 B.n386 B.n385 10.6151
R1047 B.n387 B.n386 10.6151
R1048 B.n387 B.n134 10.6151
R1049 B.n391 B.n134 10.6151
R1050 B.n392 B.n391 10.6151
R1051 B.n393 B.n392 10.6151
R1052 B.n393 B.n132 10.6151
R1053 B.n397 B.n132 10.6151
R1054 B.n398 B.n397 10.6151
R1055 B.n399 B.n398 10.6151
R1056 B.n399 B.n130 10.6151
R1057 B.n403 B.n130 10.6151
R1058 B.n404 B.n403 10.6151
R1059 B.n405 B.n404 10.6151
R1060 B.n405 B.n128 10.6151
R1061 B.n409 B.n128 10.6151
R1062 B.n410 B.n409 10.6151
R1063 B.n273 B.n272 10.6151
R1064 B.n272 B.n271 10.6151
R1065 B.n271 B.n178 10.6151
R1066 B.n267 B.n178 10.6151
R1067 B.n267 B.n266 10.6151
R1068 B.n266 B.n265 10.6151
R1069 B.n265 B.n180 10.6151
R1070 B.n261 B.n180 10.6151
R1071 B.n261 B.n260 10.6151
R1072 B.n260 B.n259 10.6151
R1073 B.n259 B.n182 10.6151
R1074 B.n255 B.n182 10.6151
R1075 B.n255 B.n254 10.6151
R1076 B.n254 B.n253 10.6151
R1077 B.n253 B.n184 10.6151
R1078 B.n249 B.n184 10.6151
R1079 B.n249 B.n248 10.6151
R1080 B.n248 B.n247 10.6151
R1081 B.n247 B.n186 10.6151
R1082 B.n243 B.n186 10.6151
R1083 B.n243 B.n242 10.6151
R1084 B.n242 B.n241 10.6151
R1085 B.n241 B.n188 10.6151
R1086 B.n237 B.n188 10.6151
R1087 B.n237 B.n236 10.6151
R1088 B.n236 B.n235 10.6151
R1089 B.n235 B.n190 10.6151
R1090 B.n231 B.n190 10.6151
R1091 B.n231 B.n230 10.6151
R1092 B.n230 B.n229 10.6151
R1093 B.n229 B.n192 10.6151
R1094 B.n225 B.n192 10.6151
R1095 B.n225 B.n224 10.6151
R1096 B.n224 B.n223 10.6151
R1097 B.n223 B.n194 10.6151
R1098 B.n219 B.n194 10.6151
R1099 B.n219 B.n218 10.6151
R1100 B.n218 B.n217 10.6151
R1101 B.n217 B.n196 10.6151
R1102 B.n213 B.n196 10.6151
R1103 B.n213 B.n212 10.6151
R1104 B.n212 B.n211 10.6151
R1105 B.n211 B.n198 10.6151
R1106 B.n207 B.n198 10.6151
R1107 B.n207 B.n206 10.6151
R1108 B.n206 B.n205 10.6151
R1109 B.n205 B.n200 10.6151
R1110 B.n201 B.n200 10.6151
R1111 B.n201 B.n0 10.6151
R1112 B.n771 B.n1 10.6151
R1113 B.n771 B.n770 10.6151
R1114 B.n770 B.n769 10.6151
R1115 B.n769 B.n4 10.6151
R1116 B.n765 B.n4 10.6151
R1117 B.n765 B.n764 10.6151
R1118 B.n764 B.n763 10.6151
R1119 B.n763 B.n6 10.6151
R1120 B.n759 B.n6 10.6151
R1121 B.n759 B.n758 10.6151
R1122 B.n758 B.n757 10.6151
R1123 B.n757 B.n8 10.6151
R1124 B.n753 B.n8 10.6151
R1125 B.n753 B.n752 10.6151
R1126 B.n752 B.n751 10.6151
R1127 B.n751 B.n10 10.6151
R1128 B.n747 B.n10 10.6151
R1129 B.n747 B.n746 10.6151
R1130 B.n746 B.n745 10.6151
R1131 B.n745 B.n12 10.6151
R1132 B.n741 B.n12 10.6151
R1133 B.n741 B.n740 10.6151
R1134 B.n740 B.n739 10.6151
R1135 B.n739 B.n14 10.6151
R1136 B.n735 B.n14 10.6151
R1137 B.n735 B.n734 10.6151
R1138 B.n734 B.n733 10.6151
R1139 B.n733 B.n16 10.6151
R1140 B.n729 B.n16 10.6151
R1141 B.n729 B.n728 10.6151
R1142 B.n728 B.n727 10.6151
R1143 B.n727 B.n18 10.6151
R1144 B.n723 B.n18 10.6151
R1145 B.n723 B.n722 10.6151
R1146 B.n722 B.n721 10.6151
R1147 B.n721 B.n20 10.6151
R1148 B.n717 B.n20 10.6151
R1149 B.n717 B.n716 10.6151
R1150 B.n716 B.n715 10.6151
R1151 B.n715 B.n22 10.6151
R1152 B.n711 B.n22 10.6151
R1153 B.n711 B.n710 10.6151
R1154 B.n710 B.n709 10.6151
R1155 B.n709 B.n24 10.6151
R1156 B.n705 B.n24 10.6151
R1157 B.n705 B.n704 10.6151
R1158 B.n704 B.n703 10.6151
R1159 B.n703 B.n26 10.6151
R1160 B.n699 B.n26 10.6151
R1161 B.n639 B.n638 9.36635
R1162 B.n621 B.n56 9.36635
R1163 B.n333 B.n156 9.36635
R1164 B.n351 B.n350 9.36635
R1165 B.n775 B.n0 2.81026
R1166 B.n775 B.n1 2.81026
R1167 B.n638 B.n637 1.24928
R1168 B.n624 B.n56 1.24928
R1169 B.n336 B.n156 1.24928
R1170 B.n350 B.n349 1.24928
R1171 VN.n34 VN.n33 161.3
R1172 VN.n32 VN.n19 161.3
R1173 VN.n31 VN.n30 161.3
R1174 VN.n29 VN.n20 161.3
R1175 VN.n28 VN.n27 161.3
R1176 VN.n26 VN.n21 161.3
R1177 VN.n25 VN.n24 161.3
R1178 VN.n16 VN.n15 161.3
R1179 VN.n14 VN.n1 161.3
R1180 VN.n13 VN.n12 161.3
R1181 VN.n11 VN.n2 161.3
R1182 VN.n10 VN.n9 161.3
R1183 VN.n8 VN.n3 161.3
R1184 VN.n7 VN.n6 161.3
R1185 VN.n23 VN.t0 118.43
R1186 VN.n5 VN.t5 118.43
R1187 VN.n4 VN.t2 85.507
R1188 VN.n0 VN.t4 85.507
R1189 VN.n22 VN.t1 85.507
R1190 VN.n18 VN.t3 85.507
R1191 VN.n17 VN.n0 74.7981
R1192 VN.n35 VN.n18 74.7981
R1193 VN.n5 VN.n4 61.8808
R1194 VN.n23 VN.n22 61.8808
R1195 VN VN.n35 51.0055
R1196 VN.n13 VN.n2 43.3318
R1197 VN.n31 VN.n20 43.3318
R1198 VN.n9 VN.n2 37.4894
R1199 VN.n27 VN.n20 37.4894
R1200 VN.n8 VN.n7 24.3439
R1201 VN.n9 VN.n8 24.3439
R1202 VN.n14 VN.n13 24.3439
R1203 VN.n15 VN.n14 24.3439
R1204 VN.n27 VN.n26 24.3439
R1205 VN.n26 VN.n25 24.3439
R1206 VN.n33 VN.n32 24.3439
R1207 VN.n32 VN.n31 24.3439
R1208 VN.n15 VN.n0 15.0934
R1209 VN.n33 VN.n18 15.0934
R1210 VN.n7 VN.n4 12.1722
R1211 VN.n25 VN.n22 12.1722
R1212 VN.n24 VN.n23 4.14964
R1213 VN.n6 VN.n5 4.14964
R1214 VN.n35 VN.n34 0.355081
R1215 VN.n17 VN.n16 0.355081
R1216 VN VN.n17 0.26685
R1217 VN.n34 VN.n19 0.189894
R1218 VN.n30 VN.n19 0.189894
R1219 VN.n30 VN.n29 0.189894
R1220 VN.n29 VN.n28 0.189894
R1221 VN.n28 VN.n21 0.189894
R1222 VN.n24 VN.n21 0.189894
R1223 VN.n6 VN.n3 0.189894
R1224 VN.n10 VN.n3 0.189894
R1225 VN.n11 VN.n10 0.189894
R1226 VN.n12 VN.n11 0.189894
R1227 VN.n12 VN.n1 0.189894
R1228 VN.n16 VN.n1 0.189894
R1229 VTAIL.n250 VTAIL.n194 756.745
R1230 VTAIL.n58 VTAIL.n2 756.745
R1231 VTAIL.n188 VTAIL.n132 756.745
R1232 VTAIL.n124 VTAIL.n68 756.745
R1233 VTAIL.n215 VTAIL.n214 585
R1234 VTAIL.n217 VTAIL.n216 585
R1235 VTAIL.n210 VTAIL.n209 585
R1236 VTAIL.n223 VTAIL.n222 585
R1237 VTAIL.n225 VTAIL.n224 585
R1238 VTAIL.n206 VTAIL.n205 585
R1239 VTAIL.n232 VTAIL.n231 585
R1240 VTAIL.n233 VTAIL.n204 585
R1241 VTAIL.n235 VTAIL.n234 585
R1242 VTAIL.n202 VTAIL.n201 585
R1243 VTAIL.n241 VTAIL.n240 585
R1244 VTAIL.n243 VTAIL.n242 585
R1245 VTAIL.n198 VTAIL.n197 585
R1246 VTAIL.n249 VTAIL.n248 585
R1247 VTAIL.n251 VTAIL.n250 585
R1248 VTAIL.n23 VTAIL.n22 585
R1249 VTAIL.n25 VTAIL.n24 585
R1250 VTAIL.n18 VTAIL.n17 585
R1251 VTAIL.n31 VTAIL.n30 585
R1252 VTAIL.n33 VTAIL.n32 585
R1253 VTAIL.n14 VTAIL.n13 585
R1254 VTAIL.n40 VTAIL.n39 585
R1255 VTAIL.n41 VTAIL.n12 585
R1256 VTAIL.n43 VTAIL.n42 585
R1257 VTAIL.n10 VTAIL.n9 585
R1258 VTAIL.n49 VTAIL.n48 585
R1259 VTAIL.n51 VTAIL.n50 585
R1260 VTAIL.n6 VTAIL.n5 585
R1261 VTAIL.n57 VTAIL.n56 585
R1262 VTAIL.n59 VTAIL.n58 585
R1263 VTAIL.n189 VTAIL.n188 585
R1264 VTAIL.n187 VTAIL.n186 585
R1265 VTAIL.n136 VTAIL.n135 585
R1266 VTAIL.n181 VTAIL.n180 585
R1267 VTAIL.n179 VTAIL.n178 585
R1268 VTAIL.n140 VTAIL.n139 585
R1269 VTAIL.n144 VTAIL.n142 585
R1270 VTAIL.n173 VTAIL.n172 585
R1271 VTAIL.n171 VTAIL.n170 585
R1272 VTAIL.n146 VTAIL.n145 585
R1273 VTAIL.n165 VTAIL.n164 585
R1274 VTAIL.n163 VTAIL.n162 585
R1275 VTAIL.n150 VTAIL.n149 585
R1276 VTAIL.n157 VTAIL.n156 585
R1277 VTAIL.n155 VTAIL.n154 585
R1278 VTAIL.n125 VTAIL.n124 585
R1279 VTAIL.n123 VTAIL.n122 585
R1280 VTAIL.n72 VTAIL.n71 585
R1281 VTAIL.n117 VTAIL.n116 585
R1282 VTAIL.n115 VTAIL.n114 585
R1283 VTAIL.n76 VTAIL.n75 585
R1284 VTAIL.n80 VTAIL.n78 585
R1285 VTAIL.n109 VTAIL.n108 585
R1286 VTAIL.n107 VTAIL.n106 585
R1287 VTAIL.n82 VTAIL.n81 585
R1288 VTAIL.n101 VTAIL.n100 585
R1289 VTAIL.n99 VTAIL.n98 585
R1290 VTAIL.n86 VTAIL.n85 585
R1291 VTAIL.n93 VTAIL.n92 585
R1292 VTAIL.n91 VTAIL.n90 585
R1293 VTAIL.n213 VTAIL.t9 329.036
R1294 VTAIL.n21 VTAIL.t0 329.036
R1295 VTAIL.n153 VTAIL.t3 329.036
R1296 VTAIL.n89 VTAIL.t11 329.036
R1297 VTAIL.n216 VTAIL.n215 171.744
R1298 VTAIL.n216 VTAIL.n209 171.744
R1299 VTAIL.n223 VTAIL.n209 171.744
R1300 VTAIL.n224 VTAIL.n223 171.744
R1301 VTAIL.n224 VTAIL.n205 171.744
R1302 VTAIL.n232 VTAIL.n205 171.744
R1303 VTAIL.n233 VTAIL.n232 171.744
R1304 VTAIL.n234 VTAIL.n233 171.744
R1305 VTAIL.n234 VTAIL.n201 171.744
R1306 VTAIL.n241 VTAIL.n201 171.744
R1307 VTAIL.n242 VTAIL.n241 171.744
R1308 VTAIL.n242 VTAIL.n197 171.744
R1309 VTAIL.n249 VTAIL.n197 171.744
R1310 VTAIL.n250 VTAIL.n249 171.744
R1311 VTAIL.n24 VTAIL.n23 171.744
R1312 VTAIL.n24 VTAIL.n17 171.744
R1313 VTAIL.n31 VTAIL.n17 171.744
R1314 VTAIL.n32 VTAIL.n31 171.744
R1315 VTAIL.n32 VTAIL.n13 171.744
R1316 VTAIL.n40 VTAIL.n13 171.744
R1317 VTAIL.n41 VTAIL.n40 171.744
R1318 VTAIL.n42 VTAIL.n41 171.744
R1319 VTAIL.n42 VTAIL.n9 171.744
R1320 VTAIL.n49 VTAIL.n9 171.744
R1321 VTAIL.n50 VTAIL.n49 171.744
R1322 VTAIL.n50 VTAIL.n5 171.744
R1323 VTAIL.n57 VTAIL.n5 171.744
R1324 VTAIL.n58 VTAIL.n57 171.744
R1325 VTAIL.n188 VTAIL.n187 171.744
R1326 VTAIL.n187 VTAIL.n135 171.744
R1327 VTAIL.n180 VTAIL.n135 171.744
R1328 VTAIL.n180 VTAIL.n179 171.744
R1329 VTAIL.n179 VTAIL.n139 171.744
R1330 VTAIL.n144 VTAIL.n139 171.744
R1331 VTAIL.n172 VTAIL.n144 171.744
R1332 VTAIL.n172 VTAIL.n171 171.744
R1333 VTAIL.n171 VTAIL.n145 171.744
R1334 VTAIL.n164 VTAIL.n145 171.744
R1335 VTAIL.n164 VTAIL.n163 171.744
R1336 VTAIL.n163 VTAIL.n149 171.744
R1337 VTAIL.n156 VTAIL.n149 171.744
R1338 VTAIL.n156 VTAIL.n155 171.744
R1339 VTAIL.n124 VTAIL.n123 171.744
R1340 VTAIL.n123 VTAIL.n71 171.744
R1341 VTAIL.n116 VTAIL.n71 171.744
R1342 VTAIL.n116 VTAIL.n115 171.744
R1343 VTAIL.n115 VTAIL.n75 171.744
R1344 VTAIL.n80 VTAIL.n75 171.744
R1345 VTAIL.n108 VTAIL.n80 171.744
R1346 VTAIL.n108 VTAIL.n107 171.744
R1347 VTAIL.n107 VTAIL.n81 171.744
R1348 VTAIL.n100 VTAIL.n81 171.744
R1349 VTAIL.n100 VTAIL.n99 171.744
R1350 VTAIL.n99 VTAIL.n85 171.744
R1351 VTAIL.n92 VTAIL.n85 171.744
R1352 VTAIL.n92 VTAIL.n91 171.744
R1353 VTAIL.n215 VTAIL.t9 85.8723
R1354 VTAIL.n23 VTAIL.t0 85.8723
R1355 VTAIL.n155 VTAIL.t3 85.8723
R1356 VTAIL.n91 VTAIL.t11 85.8723
R1357 VTAIL.n131 VTAIL.n130 59.2678
R1358 VTAIL.n67 VTAIL.n66 59.2678
R1359 VTAIL.n1 VTAIL.n0 59.2676
R1360 VTAIL.n65 VTAIL.n64 59.2676
R1361 VTAIL.n255 VTAIL.n254 33.349
R1362 VTAIL.n63 VTAIL.n62 33.349
R1363 VTAIL.n193 VTAIL.n192 33.349
R1364 VTAIL.n129 VTAIL.n128 33.349
R1365 VTAIL.n67 VTAIL.n65 28.3841
R1366 VTAIL.n255 VTAIL.n193 25.3152
R1367 VTAIL.n235 VTAIL.n202 13.1884
R1368 VTAIL.n43 VTAIL.n10 13.1884
R1369 VTAIL.n142 VTAIL.n140 13.1884
R1370 VTAIL.n78 VTAIL.n76 13.1884
R1371 VTAIL.n236 VTAIL.n204 12.8005
R1372 VTAIL.n240 VTAIL.n239 12.8005
R1373 VTAIL.n44 VTAIL.n12 12.8005
R1374 VTAIL.n48 VTAIL.n47 12.8005
R1375 VTAIL.n178 VTAIL.n177 12.8005
R1376 VTAIL.n174 VTAIL.n173 12.8005
R1377 VTAIL.n114 VTAIL.n113 12.8005
R1378 VTAIL.n110 VTAIL.n109 12.8005
R1379 VTAIL.n231 VTAIL.n230 12.0247
R1380 VTAIL.n243 VTAIL.n200 12.0247
R1381 VTAIL.n39 VTAIL.n38 12.0247
R1382 VTAIL.n51 VTAIL.n8 12.0247
R1383 VTAIL.n181 VTAIL.n138 12.0247
R1384 VTAIL.n170 VTAIL.n143 12.0247
R1385 VTAIL.n117 VTAIL.n74 12.0247
R1386 VTAIL.n106 VTAIL.n79 12.0247
R1387 VTAIL.n229 VTAIL.n206 11.249
R1388 VTAIL.n244 VTAIL.n198 11.249
R1389 VTAIL.n37 VTAIL.n14 11.249
R1390 VTAIL.n52 VTAIL.n6 11.249
R1391 VTAIL.n182 VTAIL.n136 11.249
R1392 VTAIL.n169 VTAIL.n146 11.249
R1393 VTAIL.n118 VTAIL.n72 11.249
R1394 VTAIL.n105 VTAIL.n82 11.249
R1395 VTAIL.n214 VTAIL.n213 10.7239
R1396 VTAIL.n22 VTAIL.n21 10.7239
R1397 VTAIL.n154 VTAIL.n153 10.7239
R1398 VTAIL.n90 VTAIL.n89 10.7239
R1399 VTAIL.n226 VTAIL.n225 10.4732
R1400 VTAIL.n248 VTAIL.n247 10.4732
R1401 VTAIL.n34 VTAIL.n33 10.4732
R1402 VTAIL.n56 VTAIL.n55 10.4732
R1403 VTAIL.n186 VTAIL.n185 10.4732
R1404 VTAIL.n166 VTAIL.n165 10.4732
R1405 VTAIL.n122 VTAIL.n121 10.4732
R1406 VTAIL.n102 VTAIL.n101 10.4732
R1407 VTAIL.n222 VTAIL.n208 9.69747
R1408 VTAIL.n251 VTAIL.n196 9.69747
R1409 VTAIL.n30 VTAIL.n16 9.69747
R1410 VTAIL.n59 VTAIL.n4 9.69747
R1411 VTAIL.n189 VTAIL.n134 9.69747
R1412 VTAIL.n162 VTAIL.n148 9.69747
R1413 VTAIL.n125 VTAIL.n70 9.69747
R1414 VTAIL.n98 VTAIL.n84 9.69747
R1415 VTAIL.n254 VTAIL.n253 9.45567
R1416 VTAIL.n62 VTAIL.n61 9.45567
R1417 VTAIL.n192 VTAIL.n191 9.45567
R1418 VTAIL.n128 VTAIL.n127 9.45567
R1419 VTAIL.n253 VTAIL.n252 9.3005
R1420 VTAIL.n196 VTAIL.n195 9.3005
R1421 VTAIL.n247 VTAIL.n246 9.3005
R1422 VTAIL.n245 VTAIL.n244 9.3005
R1423 VTAIL.n200 VTAIL.n199 9.3005
R1424 VTAIL.n239 VTAIL.n238 9.3005
R1425 VTAIL.n212 VTAIL.n211 9.3005
R1426 VTAIL.n219 VTAIL.n218 9.3005
R1427 VTAIL.n221 VTAIL.n220 9.3005
R1428 VTAIL.n208 VTAIL.n207 9.3005
R1429 VTAIL.n227 VTAIL.n226 9.3005
R1430 VTAIL.n229 VTAIL.n228 9.3005
R1431 VTAIL.n230 VTAIL.n203 9.3005
R1432 VTAIL.n237 VTAIL.n236 9.3005
R1433 VTAIL.n61 VTAIL.n60 9.3005
R1434 VTAIL.n4 VTAIL.n3 9.3005
R1435 VTAIL.n55 VTAIL.n54 9.3005
R1436 VTAIL.n53 VTAIL.n52 9.3005
R1437 VTAIL.n8 VTAIL.n7 9.3005
R1438 VTAIL.n47 VTAIL.n46 9.3005
R1439 VTAIL.n20 VTAIL.n19 9.3005
R1440 VTAIL.n27 VTAIL.n26 9.3005
R1441 VTAIL.n29 VTAIL.n28 9.3005
R1442 VTAIL.n16 VTAIL.n15 9.3005
R1443 VTAIL.n35 VTAIL.n34 9.3005
R1444 VTAIL.n37 VTAIL.n36 9.3005
R1445 VTAIL.n38 VTAIL.n11 9.3005
R1446 VTAIL.n45 VTAIL.n44 9.3005
R1447 VTAIL.n152 VTAIL.n151 9.3005
R1448 VTAIL.n159 VTAIL.n158 9.3005
R1449 VTAIL.n161 VTAIL.n160 9.3005
R1450 VTAIL.n148 VTAIL.n147 9.3005
R1451 VTAIL.n167 VTAIL.n166 9.3005
R1452 VTAIL.n169 VTAIL.n168 9.3005
R1453 VTAIL.n143 VTAIL.n141 9.3005
R1454 VTAIL.n175 VTAIL.n174 9.3005
R1455 VTAIL.n191 VTAIL.n190 9.3005
R1456 VTAIL.n134 VTAIL.n133 9.3005
R1457 VTAIL.n185 VTAIL.n184 9.3005
R1458 VTAIL.n183 VTAIL.n182 9.3005
R1459 VTAIL.n138 VTAIL.n137 9.3005
R1460 VTAIL.n177 VTAIL.n176 9.3005
R1461 VTAIL.n88 VTAIL.n87 9.3005
R1462 VTAIL.n95 VTAIL.n94 9.3005
R1463 VTAIL.n97 VTAIL.n96 9.3005
R1464 VTAIL.n84 VTAIL.n83 9.3005
R1465 VTAIL.n103 VTAIL.n102 9.3005
R1466 VTAIL.n105 VTAIL.n104 9.3005
R1467 VTAIL.n79 VTAIL.n77 9.3005
R1468 VTAIL.n111 VTAIL.n110 9.3005
R1469 VTAIL.n127 VTAIL.n126 9.3005
R1470 VTAIL.n70 VTAIL.n69 9.3005
R1471 VTAIL.n121 VTAIL.n120 9.3005
R1472 VTAIL.n119 VTAIL.n118 9.3005
R1473 VTAIL.n74 VTAIL.n73 9.3005
R1474 VTAIL.n113 VTAIL.n112 9.3005
R1475 VTAIL.n221 VTAIL.n210 8.92171
R1476 VTAIL.n252 VTAIL.n194 8.92171
R1477 VTAIL.n29 VTAIL.n18 8.92171
R1478 VTAIL.n60 VTAIL.n2 8.92171
R1479 VTAIL.n190 VTAIL.n132 8.92171
R1480 VTAIL.n161 VTAIL.n150 8.92171
R1481 VTAIL.n126 VTAIL.n68 8.92171
R1482 VTAIL.n97 VTAIL.n86 8.92171
R1483 VTAIL.n218 VTAIL.n217 8.14595
R1484 VTAIL.n26 VTAIL.n25 8.14595
R1485 VTAIL.n158 VTAIL.n157 8.14595
R1486 VTAIL.n94 VTAIL.n93 8.14595
R1487 VTAIL.n214 VTAIL.n212 7.3702
R1488 VTAIL.n22 VTAIL.n20 7.3702
R1489 VTAIL.n154 VTAIL.n152 7.3702
R1490 VTAIL.n90 VTAIL.n88 7.3702
R1491 VTAIL.n217 VTAIL.n212 5.81868
R1492 VTAIL.n25 VTAIL.n20 5.81868
R1493 VTAIL.n157 VTAIL.n152 5.81868
R1494 VTAIL.n93 VTAIL.n88 5.81868
R1495 VTAIL.n218 VTAIL.n210 5.04292
R1496 VTAIL.n254 VTAIL.n194 5.04292
R1497 VTAIL.n26 VTAIL.n18 5.04292
R1498 VTAIL.n62 VTAIL.n2 5.04292
R1499 VTAIL.n192 VTAIL.n132 5.04292
R1500 VTAIL.n158 VTAIL.n150 5.04292
R1501 VTAIL.n128 VTAIL.n68 5.04292
R1502 VTAIL.n94 VTAIL.n86 5.04292
R1503 VTAIL.n222 VTAIL.n221 4.26717
R1504 VTAIL.n252 VTAIL.n251 4.26717
R1505 VTAIL.n30 VTAIL.n29 4.26717
R1506 VTAIL.n60 VTAIL.n59 4.26717
R1507 VTAIL.n190 VTAIL.n189 4.26717
R1508 VTAIL.n162 VTAIL.n161 4.26717
R1509 VTAIL.n126 VTAIL.n125 4.26717
R1510 VTAIL.n98 VTAIL.n97 4.26717
R1511 VTAIL.n225 VTAIL.n208 3.49141
R1512 VTAIL.n248 VTAIL.n196 3.49141
R1513 VTAIL.n33 VTAIL.n16 3.49141
R1514 VTAIL.n56 VTAIL.n4 3.49141
R1515 VTAIL.n186 VTAIL.n134 3.49141
R1516 VTAIL.n165 VTAIL.n148 3.49141
R1517 VTAIL.n122 VTAIL.n70 3.49141
R1518 VTAIL.n101 VTAIL.n84 3.49141
R1519 VTAIL.n129 VTAIL.n67 3.06947
R1520 VTAIL.n193 VTAIL.n131 3.06947
R1521 VTAIL.n65 VTAIL.n63 3.06947
R1522 VTAIL.n0 VTAIL.t10 2.83689
R1523 VTAIL.n0 VTAIL.t8 2.83689
R1524 VTAIL.n64 VTAIL.t5 2.83689
R1525 VTAIL.n64 VTAIL.t2 2.83689
R1526 VTAIL.n130 VTAIL.t1 2.83689
R1527 VTAIL.n130 VTAIL.t4 2.83689
R1528 VTAIL.n66 VTAIL.t6 2.83689
R1529 VTAIL.n66 VTAIL.t7 2.83689
R1530 VTAIL.n226 VTAIL.n206 2.71565
R1531 VTAIL.n247 VTAIL.n198 2.71565
R1532 VTAIL.n34 VTAIL.n14 2.71565
R1533 VTAIL.n55 VTAIL.n6 2.71565
R1534 VTAIL.n185 VTAIL.n136 2.71565
R1535 VTAIL.n166 VTAIL.n146 2.71565
R1536 VTAIL.n121 VTAIL.n72 2.71565
R1537 VTAIL.n102 VTAIL.n82 2.71565
R1538 VTAIL.n213 VTAIL.n211 2.41282
R1539 VTAIL.n21 VTAIL.n19 2.41282
R1540 VTAIL.n153 VTAIL.n151 2.41282
R1541 VTAIL.n89 VTAIL.n87 2.41282
R1542 VTAIL VTAIL.n255 2.24403
R1543 VTAIL.n131 VTAIL.n129 2.00481
R1544 VTAIL.n63 VTAIL.n1 2.00481
R1545 VTAIL.n231 VTAIL.n229 1.93989
R1546 VTAIL.n244 VTAIL.n243 1.93989
R1547 VTAIL.n39 VTAIL.n37 1.93989
R1548 VTAIL.n52 VTAIL.n51 1.93989
R1549 VTAIL.n182 VTAIL.n181 1.93989
R1550 VTAIL.n170 VTAIL.n169 1.93989
R1551 VTAIL.n118 VTAIL.n117 1.93989
R1552 VTAIL.n106 VTAIL.n105 1.93989
R1553 VTAIL.n230 VTAIL.n204 1.16414
R1554 VTAIL.n240 VTAIL.n200 1.16414
R1555 VTAIL.n38 VTAIL.n12 1.16414
R1556 VTAIL.n48 VTAIL.n8 1.16414
R1557 VTAIL.n178 VTAIL.n138 1.16414
R1558 VTAIL.n173 VTAIL.n143 1.16414
R1559 VTAIL.n114 VTAIL.n74 1.16414
R1560 VTAIL.n109 VTAIL.n79 1.16414
R1561 VTAIL VTAIL.n1 0.825931
R1562 VTAIL.n236 VTAIL.n235 0.388379
R1563 VTAIL.n239 VTAIL.n202 0.388379
R1564 VTAIL.n44 VTAIL.n43 0.388379
R1565 VTAIL.n47 VTAIL.n10 0.388379
R1566 VTAIL.n177 VTAIL.n140 0.388379
R1567 VTAIL.n174 VTAIL.n142 0.388379
R1568 VTAIL.n113 VTAIL.n76 0.388379
R1569 VTAIL.n110 VTAIL.n78 0.388379
R1570 VTAIL.n219 VTAIL.n211 0.155672
R1571 VTAIL.n220 VTAIL.n219 0.155672
R1572 VTAIL.n220 VTAIL.n207 0.155672
R1573 VTAIL.n227 VTAIL.n207 0.155672
R1574 VTAIL.n228 VTAIL.n227 0.155672
R1575 VTAIL.n228 VTAIL.n203 0.155672
R1576 VTAIL.n237 VTAIL.n203 0.155672
R1577 VTAIL.n238 VTAIL.n237 0.155672
R1578 VTAIL.n238 VTAIL.n199 0.155672
R1579 VTAIL.n245 VTAIL.n199 0.155672
R1580 VTAIL.n246 VTAIL.n245 0.155672
R1581 VTAIL.n246 VTAIL.n195 0.155672
R1582 VTAIL.n253 VTAIL.n195 0.155672
R1583 VTAIL.n27 VTAIL.n19 0.155672
R1584 VTAIL.n28 VTAIL.n27 0.155672
R1585 VTAIL.n28 VTAIL.n15 0.155672
R1586 VTAIL.n35 VTAIL.n15 0.155672
R1587 VTAIL.n36 VTAIL.n35 0.155672
R1588 VTAIL.n36 VTAIL.n11 0.155672
R1589 VTAIL.n45 VTAIL.n11 0.155672
R1590 VTAIL.n46 VTAIL.n45 0.155672
R1591 VTAIL.n46 VTAIL.n7 0.155672
R1592 VTAIL.n53 VTAIL.n7 0.155672
R1593 VTAIL.n54 VTAIL.n53 0.155672
R1594 VTAIL.n54 VTAIL.n3 0.155672
R1595 VTAIL.n61 VTAIL.n3 0.155672
R1596 VTAIL.n191 VTAIL.n133 0.155672
R1597 VTAIL.n184 VTAIL.n133 0.155672
R1598 VTAIL.n184 VTAIL.n183 0.155672
R1599 VTAIL.n183 VTAIL.n137 0.155672
R1600 VTAIL.n176 VTAIL.n137 0.155672
R1601 VTAIL.n176 VTAIL.n175 0.155672
R1602 VTAIL.n175 VTAIL.n141 0.155672
R1603 VTAIL.n168 VTAIL.n141 0.155672
R1604 VTAIL.n168 VTAIL.n167 0.155672
R1605 VTAIL.n167 VTAIL.n147 0.155672
R1606 VTAIL.n160 VTAIL.n147 0.155672
R1607 VTAIL.n160 VTAIL.n159 0.155672
R1608 VTAIL.n159 VTAIL.n151 0.155672
R1609 VTAIL.n127 VTAIL.n69 0.155672
R1610 VTAIL.n120 VTAIL.n69 0.155672
R1611 VTAIL.n120 VTAIL.n119 0.155672
R1612 VTAIL.n119 VTAIL.n73 0.155672
R1613 VTAIL.n112 VTAIL.n73 0.155672
R1614 VTAIL.n112 VTAIL.n111 0.155672
R1615 VTAIL.n111 VTAIL.n77 0.155672
R1616 VTAIL.n104 VTAIL.n77 0.155672
R1617 VTAIL.n104 VTAIL.n103 0.155672
R1618 VTAIL.n103 VTAIL.n83 0.155672
R1619 VTAIL.n96 VTAIL.n83 0.155672
R1620 VTAIL.n96 VTAIL.n95 0.155672
R1621 VTAIL.n95 VTAIL.n87 0.155672
R1622 VDD2.n119 VDD2.n63 756.745
R1623 VDD2.n56 VDD2.n0 756.745
R1624 VDD2.n120 VDD2.n119 585
R1625 VDD2.n118 VDD2.n117 585
R1626 VDD2.n67 VDD2.n66 585
R1627 VDD2.n112 VDD2.n111 585
R1628 VDD2.n110 VDD2.n109 585
R1629 VDD2.n71 VDD2.n70 585
R1630 VDD2.n75 VDD2.n73 585
R1631 VDD2.n104 VDD2.n103 585
R1632 VDD2.n102 VDD2.n101 585
R1633 VDD2.n77 VDD2.n76 585
R1634 VDD2.n96 VDD2.n95 585
R1635 VDD2.n94 VDD2.n93 585
R1636 VDD2.n81 VDD2.n80 585
R1637 VDD2.n88 VDD2.n87 585
R1638 VDD2.n86 VDD2.n85 585
R1639 VDD2.n21 VDD2.n20 585
R1640 VDD2.n23 VDD2.n22 585
R1641 VDD2.n16 VDD2.n15 585
R1642 VDD2.n29 VDD2.n28 585
R1643 VDD2.n31 VDD2.n30 585
R1644 VDD2.n12 VDD2.n11 585
R1645 VDD2.n38 VDD2.n37 585
R1646 VDD2.n39 VDD2.n10 585
R1647 VDD2.n41 VDD2.n40 585
R1648 VDD2.n8 VDD2.n7 585
R1649 VDD2.n47 VDD2.n46 585
R1650 VDD2.n49 VDD2.n48 585
R1651 VDD2.n4 VDD2.n3 585
R1652 VDD2.n55 VDD2.n54 585
R1653 VDD2.n57 VDD2.n56 585
R1654 VDD2.n84 VDD2.t2 329.036
R1655 VDD2.n19 VDD2.t0 329.036
R1656 VDD2.n119 VDD2.n118 171.744
R1657 VDD2.n118 VDD2.n66 171.744
R1658 VDD2.n111 VDD2.n66 171.744
R1659 VDD2.n111 VDD2.n110 171.744
R1660 VDD2.n110 VDD2.n70 171.744
R1661 VDD2.n75 VDD2.n70 171.744
R1662 VDD2.n103 VDD2.n75 171.744
R1663 VDD2.n103 VDD2.n102 171.744
R1664 VDD2.n102 VDD2.n76 171.744
R1665 VDD2.n95 VDD2.n76 171.744
R1666 VDD2.n95 VDD2.n94 171.744
R1667 VDD2.n94 VDD2.n80 171.744
R1668 VDD2.n87 VDD2.n80 171.744
R1669 VDD2.n87 VDD2.n86 171.744
R1670 VDD2.n22 VDD2.n21 171.744
R1671 VDD2.n22 VDD2.n15 171.744
R1672 VDD2.n29 VDD2.n15 171.744
R1673 VDD2.n30 VDD2.n29 171.744
R1674 VDD2.n30 VDD2.n11 171.744
R1675 VDD2.n38 VDD2.n11 171.744
R1676 VDD2.n39 VDD2.n38 171.744
R1677 VDD2.n40 VDD2.n39 171.744
R1678 VDD2.n40 VDD2.n7 171.744
R1679 VDD2.n47 VDD2.n7 171.744
R1680 VDD2.n48 VDD2.n47 171.744
R1681 VDD2.n48 VDD2.n3 171.744
R1682 VDD2.n55 VDD2.n3 171.744
R1683 VDD2.n56 VDD2.n55 171.744
R1684 VDD2.n86 VDD2.t2 85.8723
R1685 VDD2.n21 VDD2.t0 85.8723
R1686 VDD2.n62 VDD2.n61 76.6583
R1687 VDD2 VDD2.n125 76.6555
R1688 VDD2.n62 VDD2.n60 52.2742
R1689 VDD2.n124 VDD2.n123 50.0278
R1690 VDD2.n124 VDD2.n62 43.5687
R1691 VDD2.n73 VDD2.n71 13.1884
R1692 VDD2.n41 VDD2.n8 13.1884
R1693 VDD2.n109 VDD2.n108 12.8005
R1694 VDD2.n105 VDD2.n104 12.8005
R1695 VDD2.n42 VDD2.n10 12.8005
R1696 VDD2.n46 VDD2.n45 12.8005
R1697 VDD2.n112 VDD2.n69 12.0247
R1698 VDD2.n101 VDD2.n74 12.0247
R1699 VDD2.n37 VDD2.n36 12.0247
R1700 VDD2.n49 VDD2.n6 12.0247
R1701 VDD2.n113 VDD2.n67 11.249
R1702 VDD2.n100 VDD2.n77 11.249
R1703 VDD2.n35 VDD2.n12 11.249
R1704 VDD2.n50 VDD2.n4 11.249
R1705 VDD2.n85 VDD2.n84 10.7239
R1706 VDD2.n20 VDD2.n19 10.7239
R1707 VDD2.n117 VDD2.n116 10.4732
R1708 VDD2.n97 VDD2.n96 10.4732
R1709 VDD2.n32 VDD2.n31 10.4732
R1710 VDD2.n54 VDD2.n53 10.4732
R1711 VDD2.n120 VDD2.n65 9.69747
R1712 VDD2.n93 VDD2.n79 9.69747
R1713 VDD2.n28 VDD2.n14 9.69747
R1714 VDD2.n57 VDD2.n2 9.69747
R1715 VDD2.n123 VDD2.n122 9.45567
R1716 VDD2.n60 VDD2.n59 9.45567
R1717 VDD2.n83 VDD2.n82 9.3005
R1718 VDD2.n90 VDD2.n89 9.3005
R1719 VDD2.n92 VDD2.n91 9.3005
R1720 VDD2.n79 VDD2.n78 9.3005
R1721 VDD2.n98 VDD2.n97 9.3005
R1722 VDD2.n100 VDD2.n99 9.3005
R1723 VDD2.n74 VDD2.n72 9.3005
R1724 VDD2.n106 VDD2.n105 9.3005
R1725 VDD2.n122 VDD2.n121 9.3005
R1726 VDD2.n65 VDD2.n64 9.3005
R1727 VDD2.n116 VDD2.n115 9.3005
R1728 VDD2.n114 VDD2.n113 9.3005
R1729 VDD2.n69 VDD2.n68 9.3005
R1730 VDD2.n108 VDD2.n107 9.3005
R1731 VDD2.n59 VDD2.n58 9.3005
R1732 VDD2.n2 VDD2.n1 9.3005
R1733 VDD2.n53 VDD2.n52 9.3005
R1734 VDD2.n51 VDD2.n50 9.3005
R1735 VDD2.n6 VDD2.n5 9.3005
R1736 VDD2.n45 VDD2.n44 9.3005
R1737 VDD2.n18 VDD2.n17 9.3005
R1738 VDD2.n25 VDD2.n24 9.3005
R1739 VDD2.n27 VDD2.n26 9.3005
R1740 VDD2.n14 VDD2.n13 9.3005
R1741 VDD2.n33 VDD2.n32 9.3005
R1742 VDD2.n35 VDD2.n34 9.3005
R1743 VDD2.n36 VDD2.n9 9.3005
R1744 VDD2.n43 VDD2.n42 9.3005
R1745 VDD2.n121 VDD2.n63 8.92171
R1746 VDD2.n92 VDD2.n81 8.92171
R1747 VDD2.n27 VDD2.n16 8.92171
R1748 VDD2.n58 VDD2.n0 8.92171
R1749 VDD2.n89 VDD2.n88 8.14595
R1750 VDD2.n24 VDD2.n23 8.14595
R1751 VDD2.n85 VDD2.n83 7.3702
R1752 VDD2.n20 VDD2.n18 7.3702
R1753 VDD2.n88 VDD2.n83 5.81868
R1754 VDD2.n23 VDD2.n18 5.81868
R1755 VDD2.n123 VDD2.n63 5.04292
R1756 VDD2.n89 VDD2.n81 5.04292
R1757 VDD2.n24 VDD2.n16 5.04292
R1758 VDD2.n60 VDD2.n0 5.04292
R1759 VDD2.n121 VDD2.n120 4.26717
R1760 VDD2.n93 VDD2.n92 4.26717
R1761 VDD2.n28 VDD2.n27 4.26717
R1762 VDD2.n58 VDD2.n57 4.26717
R1763 VDD2.n117 VDD2.n65 3.49141
R1764 VDD2.n96 VDD2.n79 3.49141
R1765 VDD2.n31 VDD2.n14 3.49141
R1766 VDD2.n54 VDD2.n2 3.49141
R1767 VDD2.n125 VDD2.t4 2.83689
R1768 VDD2.n125 VDD2.t5 2.83689
R1769 VDD2.n61 VDD2.t3 2.83689
R1770 VDD2.n61 VDD2.t1 2.83689
R1771 VDD2.n116 VDD2.n67 2.71565
R1772 VDD2.n97 VDD2.n77 2.71565
R1773 VDD2.n32 VDD2.n12 2.71565
R1774 VDD2.n53 VDD2.n4 2.71565
R1775 VDD2.n84 VDD2.n82 2.41282
R1776 VDD2.n19 VDD2.n17 2.41282
R1777 VDD2 VDD2.n124 2.36041
R1778 VDD2.n113 VDD2.n112 1.93989
R1779 VDD2.n101 VDD2.n100 1.93989
R1780 VDD2.n37 VDD2.n35 1.93989
R1781 VDD2.n50 VDD2.n49 1.93989
R1782 VDD2.n109 VDD2.n69 1.16414
R1783 VDD2.n104 VDD2.n74 1.16414
R1784 VDD2.n36 VDD2.n10 1.16414
R1785 VDD2.n46 VDD2.n6 1.16414
R1786 VDD2.n108 VDD2.n71 0.388379
R1787 VDD2.n105 VDD2.n73 0.388379
R1788 VDD2.n42 VDD2.n41 0.388379
R1789 VDD2.n45 VDD2.n8 0.388379
R1790 VDD2.n122 VDD2.n64 0.155672
R1791 VDD2.n115 VDD2.n64 0.155672
R1792 VDD2.n115 VDD2.n114 0.155672
R1793 VDD2.n114 VDD2.n68 0.155672
R1794 VDD2.n107 VDD2.n68 0.155672
R1795 VDD2.n107 VDD2.n106 0.155672
R1796 VDD2.n106 VDD2.n72 0.155672
R1797 VDD2.n99 VDD2.n72 0.155672
R1798 VDD2.n99 VDD2.n98 0.155672
R1799 VDD2.n98 VDD2.n78 0.155672
R1800 VDD2.n91 VDD2.n78 0.155672
R1801 VDD2.n91 VDD2.n90 0.155672
R1802 VDD2.n90 VDD2.n82 0.155672
R1803 VDD2.n25 VDD2.n17 0.155672
R1804 VDD2.n26 VDD2.n25 0.155672
R1805 VDD2.n26 VDD2.n13 0.155672
R1806 VDD2.n33 VDD2.n13 0.155672
R1807 VDD2.n34 VDD2.n33 0.155672
R1808 VDD2.n34 VDD2.n9 0.155672
R1809 VDD2.n43 VDD2.n9 0.155672
R1810 VDD2.n44 VDD2.n43 0.155672
R1811 VDD2.n44 VDD2.n5 0.155672
R1812 VDD2.n51 VDD2.n5 0.155672
R1813 VDD2.n52 VDD2.n51 0.155672
R1814 VDD2.n52 VDD2.n1 0.155672
R1815 VDD2.n59 VDD2.n1 0.155672
R1816 VP.n16 VP.n15 161.3
R1817 VP.n17 VP.n12 161.3
R1818 VP.n19 VP.n18 161.3
R1819 VP.n20 VP.n11 161.3
R1820 VP.n22 VP.n21 161.3
R1821 VP.n23 VP.n10 161.3
R1822 VP.n25 VP.n24 161.3
R1823 VP.n49 VP.n48 161.3
R1824 VP.n47 VP.n1 161.3
R1825 VP.n46 VP.n45 161.3
R1826 VP.n44 VP.n2 161.3
R1827 VP.n43 VP.n42 161.3
R1828 VP.n41 VP.n3 161.3
R1829 VP.n40 VP.n39 161.3
R1830 VP.n38 VP.n37 161.3
R1831 VP.n36 VP.n5 161.3
R1832 VP.n35 VP.n34 161.3
R1833 VP.n33 VP.n6 161.3
R1834 VP.n32 VP.n31 161.3
R1835 VP.n30 VP.n7 161.3
R1836 VP.n29 VP.n28 161.3
R1837 VP.n14 VP.t3 118.43
R1838 VP.n8 VP.t4 85.507
R1839 VP.n4 VP.t1 85.507
R1840 VP.n0 VP.t5 85.507
R1841 VP.n9 VP.t0 85.507
R1842 VP.n13 VP.t2 85.507
R1843 VP.n27 VP.n8 74.7981
R1844 VP.n50 VP.n0 74.7981
R1845 VP.n26 VP.n9 74.7981
R1846 VP.n14 VP.n13 61.8808
R1847 VP.n27 VP.n26 50.84
R1848 VP.n31 VP.n6 43.3318
R1849 VP.n46 VP.n2 43.3318
R1850 VP.n22 VP.n11 43.3318
R1851 VP.n35 VP.n6 37.4894
R1852 VP.n42 VP.n2 37.4894
R1853 VP.n18 VP.n11 37.4894
R1854 VP.n30 VP.n29 24.3439
R1855 VP.n31 VP.n30 24.3439
R1856 VP.n36 VP.n35 24.3439
R1857 VP.n37 VP.n36 24.3439
R1858 VP.n41 VP.n40 24.3439
R1859 VP.n42 VP.n41 24.3439
R1860 VP.n47 VP.n46 24.3439
R1861 VP.n48 VP.n47 24.3439
R1862 VP.n23 VP.n22 24.3439
R1863 VP.n24 VP.n23 24.3439
R1864 VP.n17 VP.n16 24.3439
R1865 VP.n18 VP.n17 24.3439
R1866 VP.n29 VP.n8 15.0934
R1867 VP.n48 VP.n0 15.0934
R1868 VP.n24 VP.n9 15.0934
R1869 VP.n37 VP.n4 12.1722
R1870 VP.n40 VP.n4 12.1722
R1871 VP.n16 VP.n13 12.1722
R1872 VP.n15 VP.n14 4.14962
R1873 VP.n26 VP.n25 0.355081
R1874 VP.n28 VP.n27 0.355081
R1875 VP.n50 VP.n49 0.355081
R1876 VP VP.n50 0.26685
R1877 VP.n15 VP.n12 0.189894
R1878 VP.n19 VP.n12 0.189894
R1879 VP.n20 VP.n19 0.189894
R1880 VP.n21 VP.n20 0.189894
R1881 VP.n21 VP.n10 0.189894
R1882 VP.n25 VP.n10 0.189894
R1883 VP.n28 VP.n7 0.189894
R1884 VP.n32 VP.n7 0.189894
R1885 VP.n33 VP.n32 0.189894
R1886 VP.n34 VP.n33 0.189894
R1887 VP.n34 VP.n5 0.189894
R1888 VP.n38 VP.n5 0.189894
R1889 VP.n39 VP.n38 0.189894
R1890 VP.n39 VP.n3 0.189894
R1891 VP.n43 VP.n3 0.189894
R1892 VP.n44 VP.n43 0.189894
R1893 VP.n45 VP.n44 0.189894
R1894 VP.n45 VP.n1 0.189894
R1895 VP.n49 VP.n1 0.189894
R1896 VDD1.n56 VDD1.n0 756.745
R1897 VDD1.n117 VDD1.n61 756.745
R1898 VDD1.n57 VDD1.n56 585
R1899 VDD1.n55 VDD1.n54 585
R1900 VDD1.n4 VDD1.n3 585
R1901 VDD1.n49 VDD1.n48 585
R1902 VDD1.n47 VDD1.n46 585
R1903 VDD1.n8 VDD1.n7 585
R1904 VDD1.n12 VDD1.n10 585
R1905 VDD1.n41 VDD1.n40 585
R1906 VDD1.n39 VDD1.n38 585
R1907 VDD1.n14 VDD1.n13 585
R1908 VDD1.n33 VDD1.n32 585
R1909 VDD1.n31 VDD1.n30 585
R1910 VDD1.n18 VDD1.n17 585
R1911 VDD1.n25 VDD1.n24 585
R1912 VDD1.n23 VDD1.n22 585
R1913 VDD1.n82 VDD1.n81 585
R1914 VDD1.n84 VDD1.n83 585
R1915 VDD1.n77 VDD1.n76 585
R1916 VDD1.n90 VDD1.n89 585
R1917 VDD1.n92 VDD1.n91 585
R1918 VDD1.n73 VDD1.n72 585
R1919 VDD1.n99 VDD1.n98 585
R1920 VDD1.n100 VDD1.n71 585
R1921 VDD1.n102 VDD1.n101 585
R1922 VDD1.n69 VDD1.n68 585
R1923 VDD1.n108 VDD1.n107 585
R1924 VDD1.n110 VDD1.n109 585
R1925 VDD1.n65 VDD1.n64 585
R1926 VDD1.n116 VDD1.n115 585
R1927 VDD1.n118 VDD1.n117 585
R1928 VDD1.n21 VDD1.t2 329.036
R1929 VDD1.n80 VDD1.t1 329.036
R1930 VDD1.n56 VDD1.n55 171.744
R1931 VDD1.n55 VDD1.n3 171.744
R1932 VDD1.n48 VDD1.n3 171.744
R1933 VDD1.n48 VDD1.n47 171.744
R1934 VDD1.n47 VDD1.n7 171.744
R1935 VDD1.n12 VDD1.n7 171.744
R1936 VDD1.n40 VDD1.n12 171.744
R1937 VDD1.n40 VDD1.n39 171.744
R1938 VDD1.n39 VDD1.n13 171.744
R1939 VDD1.n32 VDD1.n13 171.744
R1940 VDD1.n32 VDD1.n31 171.744
R1941 VDD1.n31 VDD1.n17 171.744
R1942 VDD1.n24 VDD1.n17 171.744
R1943 VDD1.n24 VDD1.n23 171.744
R1944 VDD1.n83 VDD1.n82 171.744
R1945 VDD1.n83 VDD1.n76 171.744
R1946 VDD1.n90 VDD1.n76 171.744
R1947 VDD1.n91 VDD1.n90 171.744
R1948 VDD1.n91 VDD1.n72 171.744
R1949 VDD1.n99 VDD1.n72 171.744
R1950 VDD1.n100 VDD1.n99 171.744
R1951 VDD1.n101 VDD1.n100 171.744
R1952 VDD1.n101 VDD1.n68 171.744
R1953 VDD1.n108 VDD1.n68 171.744
R1954 VDD1.n109 VDD1.n108 171.744
R1955 VDD1.n109 VDD1.n64 171.744
R1956 VDD1.n116 VDD1.n64 171.744
R1957 VDD1.n117 VDD1.n116 171.744
R1958 VDD1.n23 VDD1.t2 85.8723
R1959 VDD1.n82 VDD1.t1 85.8723
R1960 VDD1.n123 VDD1.n122 76.6583
R1961 VDD1.n125 VDD1.n124 75.9464
R1962 VDD1 VDD1.n60 52.3877
R1963 VDD1.n123 VDD1.n121 52.2742
R1964 VDD1.n125 VDD1.n123 45.6862
R1965 VDD1.n10 VDD1.n8 13.1884
R1966 VDD1.n102 VDD1.n69 13.1884
R1967 VDD1.n46 VDD1.n45 12.8005
R1968 VDD1.n42 VDD1.n41 12.8005
R1969 VDD1.n103 VDD1.n71 12.8005
R1970 VDD1.n107 VDD1.n106 12.8005
R1971 VDD1.n49 VDD1.n6 12.0247
R1972 VDD1.n38 VDD1.n11 12.0247
R1973 VDD1.n98 VDD1.n97 12.0247
R1974 VDD1.n110 VDD1.n67 12.0247
R1975 VDD1.n50 VDD1.n4 11.249
R1976 VDD1.n37 VDD1.n14 11.249
R1977 VDD1.n96 VDD1.n73 11.249
R1978 VDD1.n111 VDD1.n65 11.249
R1979 VDD1.n22 VDD1.n21 10.7239
R1980 VDD1.n81 VDD1.n80 10.7239
R1981 VDD1.n54 VDD1.n53 10.4732
R1982 VDD1.n34 VDD1.n33 10.4732
R1983 VDD1.n93 VDD1.n92 10.4732
R1984 VDD1.n115 VDD1.n114 10.4732
R1985 VDD1.n57 VDD1.n2 9.69747
R1986 VDD1.n30 VDD1.n16 9.69747
R1987 VDD1.n89 VDD1.n75 9.69747
R1988 VDD1.n118 VDD1.n63 9.69747
R1989 VDD1.n60 VDD1.n59 9.45567
R1990 VDD1.n121 VDD1.n120 9.45567
R1991 VDD1.n20 VDD1.n19 9.3005
R1992 VDD1.n27 VDD1.n26 9.3005
R1993 VDD1.n29 VDD1.n28 9.3005
R1994 VDD1.n16 VDD1.n15 9.3005
R1995 VDD1.n35 VDD1.n34 9.3005
R1996 VDD1.n37 VDD1.n36 9.3005
R1997 VDD1.n11 VDD1.n9 9.3005
R1998 VDD1.n43 VDD1.n42 9.3005
R1999 VDD1.n59 VDD1.n58 9.3005
R2000 VDD1.n2 VDD1.n1 9.3005
R2001 VDD1.n53 VDD1.n52 9.3005
R2002 VDD1.n51 VDD1.n50 9.3005
R2003 VDD1.n6 VDD1.n5 9.3005
R2004 VDD1.n45 VDD1.n44 9.3005
R2005 VDD1.n120 VDD1.n119 9.3005
R2006 VDD1.n63 VDD1.n62 9.3005
R2007 VDD1.n114 VDD1.n113 9.3005
R2008 VDD1.n112 VDD1.n111 9.3005
R2009 VDD1.n67 VDD1.n66 9.3005
R2010 VDD1.n106 VDD1.n105 9.3005
R2011 VDD1.n79 VDD1.n78 9.3005
R2012 VDD1.n86 VDD1.n85 9.3005
R2013 VDD1.n88 VDD1.n87 9.3005
R2014 VDD1.n75 VDD1.n74 9.3005
R2015 VDD1.n94 VDD1.n93 9.3005
R2016 VDD1.n96 VDD1.n95 9.3005
R2017 VDD1.n97 VDD1.n70 9.3005
R2018 VDD1.n104 VDD1.n103 9.3005
R2019 VDD1.n58 VDD1.n0 8.92171
R2020 VDD1.n29 VDD1.n18 8.92171
R2021 VDD1.n88 VDD1.n77 8.92171
R2022 VDD1.n119 VDD1.n61 8.92171
R2023 VDD1.n26 VDD1.n25 8.14595
R2024 VDD1.n85 VDD1.n84 8.14595
R2025 VDD1.n22 VDD1.n20 7.3702
R2026 VDD1.n81 VDD1.n79 7.3702
R2027 VDD1.n25 VDD1.n20 5.81868
R2028 VDD1.n84 VDD1.n79 5.81868
R2029 VDD1.n60 VDD1.n0 5.04292
R2030 VDD1.n26 VDD1.n18 5.04292
R2031 VDD1.n85 VDD1.n77 5.04292
R2032 VDD1.n121 VDD1.n61 5.04292
R2033 VDD1.n58 VDD1.n57 4.26717
R2034 VDD1.n30 VDD1.n29 4.26717
R2035 VDD1.n89 VDD1.n88 4.26717
R2036 VDD1.n119 VDD1.n118 4.26717
R2037 VDD1.n54 VDD1.n2 3.49141
R2038 VDD1.n33 VDD1.n16 3.49141
R2039 VDD1.n92 VDD1.n75 3.49141
R2040 VDD1.n115 VDD1.n63 3.49141
R2041 VDD1.n124 VDD1.t3 2.83689
R2042 VDD1.n124 VDD1.t5 2.83689
R2043 VDD1.n122 VDD1.t4 2.83689
R2044 VDD1.n122 VDD1.t0 2.83689
R2045 VDD1.n53 VDD1.n4 2.71565
R2046 VDD1.n34 VDD1.n14 2.71565
R2047 VDD1.n93 VDD1.n73 2.71565
R2048 VDD1.n114 VDD1.n65 2.71565
R2049 VDD1.n21 VDD1.n19 2.41282
R2050 VDD1.n80 VDD1.n78 2.41282
R2051 VDD1.n50 VDD1.n49 1.93989
R2052 VDD1.n38 VDD1.n37 1.93989
R2053 VDD1.n98 VDD1.n96 1.93989
R2054 VDD1.n111 VDD1.n110 1.93989
R2055 VDD1.n46 VDD1.n6 1.16414
R2056 VDD1.n41 VDD1.n11 1.16414
R2057 VDD1.n97 VDD1.n71 1.16414
R2058 VDD1.n107 VDD1.n67 1.16414
R2059 VDD1 VDD1.n125 0.709552
R2060 VDD1.n45 VDD1.n8 0.388379
R2061 VDD1.n42 VDD1.n10 0.388379
R2062 VDD1.n103 VDD1.n102 0.388379
R2063 VDD1.n106 VDD1.n69 0.388379
R2064 VDD1.n59 VDD1.n1 0.155672
R2065 VDD1.n52 VDD1.n1 0.155672
R2066 VDD1.n52 VDD1.n51 0.155672
R2067 VDD1.n51 VDD1.n5 0.155672
R2068 VDD1.n44 VDD1.n5 0.155672
R2069 VDD1.n44 VDD1.n43 0.155672
R2070 VDD1.n43 VDD1.n9 0.155672
R2071 VDD1.n36 VDD1.n9 0.155672
R2072 VDD1.n36 VDD1.n35 0.155672
R2073 VDD1.n35 VDD1.n15 0.155672
R2074 VDD1.n28 VDD1.n15 0.155672
R2075 VDD1.n28 VDD1.n27 0.155672
R2076 VDD1.n27 VDD1.n19 0.155672
R2077 VDD1.n86 VDD1.n78 0.155672
R2078 VDD1.n87 VDD1.n86 0.155672
R2079 VDD1.n87 VDD1.n74 0.155672
R2080 VDD1.n94 VDD1.n74 0.155672
R2081 VDD1.n95 VDD1.n94 0.155672
R2082 VDD1.n95 VDD1.n70 0.155672
R2083 VDD1.n104 VDD1.n70 0.155672
R2084 VDD1.n105 VDD1.n104 0.155672
R2085 VDD1.n105 VDD1.n66 0.155672
R2086 VDD1.n112 VDD1.n66 0.155672
R2087 VDD1.n113 VDD1.n112 0.155672
R2088 VDD1.n113 VDD1.n62 0.155672
R2089 VDD1.n120 VDD1.n62 0.155672
C0 B VDD2 2.30367f
C1 VTAIL VP 7.03729f
C2 w_n3818_n3260# B 10.3949f
C3 VN B 1.28945f
C4 VTAIL B 3.81148f
C5 VP B 2.11969f
C6 VDD1 VDD2 1.65156f
C7 w_n3818_n3260# VDD1 2.40459f
C8 VN VDD1 0.151109f
C9 VTAIL VDD1 7.72852f
C10 VP VDD1 7.04459f
C11 w_n3818_n3260# VDD2 2.50979f
C12 VN VDD2 6.68749f
C13 VDD1 B 2.21447f
C14 VN w_n3818_n3260# 7.39169f
C15 VTAIL VDD2 7.78426f
C16 VP VDD2 0.51121f
C17 VTAIL w_n3818_n3260# 2.94967f
C18 VP w_n3818_n3260# 7.88705f
C19 VN VTAIL 7.02305f
C20 VN VP 7.44651f
C21 VDD2 VSUBS 2.062479f
C22 VDD1 VSUBS 2.034674f
C23 VTAIL VSUBS 1.294051f
C24 VN VSUBS 6.43241f
C25 VP VSUBS 3.411706f
C26 B VSUBS 5.215275f
C27 w_n3818_n3260# VSUBS 0.153346p
C28 VDD1.n0 VSUBS 0.031293f
C29 VDD1.n1 VSUBS 0.028369f
C30 VDD1.n2 VSUBS 0.015244f
C31 VDD1.n3 VSUBS 0.036031f
C32 VDD1.n4 VSUBS 0.016141f
C33 VDD1.n5 VSUBS 0.028369f
C34 VDD1.n6 VSUBS 0.015244f
C35 VDD1.n7 VSUBS 0.036031f
C36 VDD1.n8 VSUBS 0.015692f
C37 VDD1.n9 VSUBS 0.028369f
C38 VDD1.n10 VSUBS 0.015692f
C39 VDD1.n11 VSUBS 0.015244f
C40 VDD1.n12 VSUBS 0.036031f
C41 VDD1.n13 VSUBS 0.036031f
C42 VDD1.n14 VSUBS 0.016141f
C43 VDD1.n15 VSUBS 0.028369f
C44 VDD1.n16 VSUBS 0.015244f
C45 VDD1.n17 VSUBS 0.036031f
C46 VDD1.n18 VSUBS 0.016141f
C47 VDD1.n19 VSUBS 1.32671f
C48 VDD1.n20 VSUBS 0.015244f
C49 VDD1.t2 VSUBS 0.077597f
C50 VDD1.n21 VSUBS 0.216498f
C51 VDD1.n22 VSUBS 0.027105f
C52 VDD1.n23 VSUBS 0.027024f
C53 VDD1.n24 VSUBS 0.036031f
C54 VDD1.n25 VSUBS 0.016141f
C55 VDD1.n26 VSUBS 0.015244f
C56 VDD1.n27 VSUBS 0.028369f
C57 VDD1.n28 VSUBS 0.028369f
C58 VDD1.n29 VSUBS 0.015244f
C59 VDD1.n30 VSUBS 0.016141f
C60 VDD1.n31 VSUBS 0.036031f
C61 VDD1.n32 VSUBS 0.036031f
C62 VDD1.n33 VSUBS 0.016141f
C63 VDD1.n34 VSUBS 0.015244f
C64 VDD1.n35 VSUBS 0.028369f
C65 VDD1.n36 VSUBS 0.028369f
C66 VDD1.n37 VSUBS 0.015244f
C67 VDD1.n38 VSUBS 0.016141f
C68 VDD1.n39 VSUBS 0.036031f
C69 VDD1.n40 VSUBS 0.036031f
C70 VDD1.n41 VSUBS 0.016141f
C71 VDD1.n42 VSUBS 0.015244f
C72 VDD1.n43 VSUBS 0.028369f
C73 VDD1.n44 VSUBS 0.028369f
C74 VDD1.n45 VSUBS 0.015244f
C75 VDD1.n46 VSUBS 0.016141f
C76 VDD1.n47 VSUBS 0.036031f
C77 VDD1.n48 VSUBS 0.036031f
C78 VDD1.n49 VSUBS 0.016141f
C79 VDD1.n50 VSUBS 0.015244f
C80 VDD1.n51 VSUBS 0.028369f
C81 VDD1.n52 VSUBS 0.028369f
C82 VDD1.n53 VSUBS 0.015244f
C83 VDD1.n54 VSUBS 0.016141f
C84 VDD1.n55 VSUBS 0.036031f
C85 VDD1.n56 VSUBS 0.087643f
C86 VDD1.n57 VSUBS 0.016141f
C87 VDD1.n58 VSUBS 0.015244f
C88 VDD1.n59 VSUBS 0.067898f
C89 VDD1.n60 VSUBS 0.075973f
C90 VDD1.n61 VSUBS 0.031293f
C91 VDD1.n62 VSUBS 0.028369f
C92 VDD1.n63 VSUBS 0.015244f
C93 VDD1.n64 VSUBS 0.036031f
C94 VDD1.n65 VSUBS 0.016141f
C95 VDD1.n66 VSUBS 0.028369f
C96 VDD1.n67 VSUBS 0.015244f
C97 VDD1.n68 VSUBS 0.036031f
C98 VDD1.n69 VSUBS 0.015692f
C99 VDD1.n70 VSUBS 0.028369f
C100 VDD1.n71 VSUBS 0.016141f
C101 VDD1.n72 VSUBS 0.036031f
C102 VDD1.n73 VSUBS 0.016141f
C103 VDD1.n74 VSUBS 0.028369f
C104 VDD1.n75 VSUBS 0.015244f
C105 VDD1.n76 VSUBS 0.036031f
C106 VDD1.n77 VSUBS 0.016141f
C107 VDD1.n78 VSUBS 1.32671f
C108 VDD1.n79 VSUBS 0.015244f
C109 VDD1.t1 VSUBS 0.077597f
C110 VDD1.n80 VSUBS 0.216498f
C111 VDD1.n81 VSUBS 0.027105f
C112 VDD1.n82 VSUBS 0.027024f
C113 VDD1.n83 VSUBS 0.036031f
C114 VDD1.n84 VSUBS 0.016141f
C115 VDD1.n85 VSUBS 0.015244f
C116 VDD1.n86 VSUBS 0.028369f
C117 VDD1.n87 VSUBS 0.028369f
C118 VDD1.n88 VSUBS 0.015244f
C119 VDD1.n89 VSUBS 0.016141f
C120 VDD1.n90 VSUBS 0.036031f
C121 VDD1.n91 VSUBS 0.036031f
C122 VDD1.n92 VSUBS 0.016141f
C123 VDD1.n93 VSUBS 0.015244f
C124 VDD1.n94 VSUBS 0.028369f
C125 VDD1.n95 VSUBS 0.028369f
C126 VDD1.n96 VSUBS 0.015244f
C127 VDD1.n97 VSUBS 0.015244f
C128 VDD1.n98 VSUBS 0.016141f
C129 VDD1.n99 VSUBS 0.036031f
C130 VDD1.n100 VSUBS 0.036031f
C131 VDD1.n101 VSUBS 0.036031f
C132 VDD1.n102 VSUBS 0.015692f
C133 VDD1.n103 VSUBS 0.015244f
C134 VDD1.n104 VSUBS 0.028369f
C135 VDD1.n105 VSUBS 0.028369f
C136 VDD1.n106 VSUBS 0.015244f
C137 VDD1.n107 VSUBS 0.016141f
C138 VDD1.n108 VSUBS 0.036031f
C139 VDD1.n109 VSUBS 0.036031f
C140 VDD1.n110 VSUBS 0.016141f
C141 VDD1.n111 VSUBS 0.015244f
C142 VDD1.n112 VSUBS 0.028369f
C143 VDD1.n113 VSUBS 0.028369f
C144 VDD1.n114 VSUBS 0.015244f
C145 VDD1.n115 VSUBS 0.016141f
C146 VDD1.n116 VSUBS 0.036031f
C147 VDD1.n117 VSUBS 0.087643f
C148 VDD1.n118 VSUBS 0.016141f
C149 VDD1.n119 VSUBS 0.015244f
C150 VDD1.n120 VSUBS 0.067898f
C151 VDD1.n121 VSUBS 0.074976f
C152 VDD1.t4 VSUBS 0.256908f
C153 VDD1.t0 VSUBS 0.256908f
C154 VDD1.n122 VSUBS 2.00105f
C155 VDD1.n123 VSUBS 3.75888f
C156 VDD1.t3 VSUBS 0.256908f
C157 VDD1.t5 VSUBS 0.256908f
C158 VDD1.n124 VSUBS 1.99286f
C159 VDD1.n125 VSUBS 3.61047f
C160 VP.t5 VSUBS 3.05485f
C161 VP.n0 VSUBS 1.19561f
C162 VP.n1 VSUBS 0.030331f
C163 VP.n2 VSUBS 0.024899f
C164 VP.n3 VSUBS 0.030331f
C165 VP.t1 VSUBS 3.05485f
C166 VP.n4 VSUBS 1.07684f
C167 VP.n5 VSUBS 0.030331f
C168 VP.n6 VSUBS 0.024899f
C169 VP.n7 VSUBS 0.030331f
C170 VP.t4 VSUBS 3.05485f
C171 VP.n8 VSUBS 1.19561f
C172 VP.t0 VSUBS 3.05485f
C173 VP.n9 VSUBS 1.19561f
C174 VP.n10 VSUBS 0.030331f
C175 VP.n11 VSUBS 0.024899f
C176 VP.n12 VSUBS 0.030331f
C177 VP.t2 VSUBS 3.05485f
C178 VP.n13 VSUBS 1.17771f
C179 VP.t3 VSUBS 3.4143f
C180 VP.n14 VSUBS 1.12393f
C181 VP.n15 VSUBS 0.353766f
C182 VP.n16 VSUBS 0.042787f
C183 VP.n17 VSUBS 0.056812f
C184 VP.n18 VSUBS 0.061337f
C185 VP.n19 VSUBS 0.030331f
C186 VP.n20 VSUBS 0.030331f
C187 VP.n21 VSUBS 0.030331f
C188 VP.n22 VSUBS 0.059516f
C189 VP.n23 VSUBS 0.056812f
C190 VP.n24 VSUBS 0.046153f
C191 VP.n25 VSUBS 0.048961f
C192 VP.n26 VSUBS 1.76535f
C193 VP.n27 VSUBS 1.78674f
C194 VP.n28 VSUBS 0.048961f
C195 VP.n29 VSUBS 0.046153f
C196 VP.n30 VSUBS 0.056812f
C197 VP.n31 VSUBS 0.059516f
C198 VP.n32 VSUBS 0.030331f
C199 VP.n33 VSUBS 0.030331f
C200 VP.n34 VSUBS 0.030331f
C201 VP.n35 VSUBS 0.061337f
C202 VP.n36 VSUBS 0.056812f
C203 VP.n37 VSUBS 0.042787f
C204 VP.n38 VSUBS 0.030331f
C205 VP.n39 VSUBS 0.030331f
C206 VP.n40 VSUBS 0.042787f
C207 VP.n41 VSUBS 0.056812f
C208 VP.n42 VSUBS 0.061337f
C209 VP.n43 VSUBS 0.030331f
C210 VP.n44 VSUBS 0.030331f
C211 VP.n45 VSUBS 0.030331f
C212 VP.n46 VSUBS 0.059516f
C213 VP.n47 VSUBS 0.056812f
C214 VP.n48 VSUBS 0.046153f
C215 VP.n49 VSUBS 0.048961f
C216 VP.n50 VSUBS 0.072f
C217 VDD2.n0 VSUBS 0.031464f
C218 VDD2.n1 VSUBS 0.028524f
C219 VDD2.n2 VSUBS 0.015327f
C220 VDD2.n3 VSUBS 0.036228f
C221 VDD2.n4 VSUBS 0.016229f
C222 VDD2.n5 VSUBS 0.028524f
C223 VDD2.n6 VSUBS 0.015327f
C224 VDD2.n7 VSUBS 0.036228f
C225 VDD2.n8 VSUBS 0.015778f
C226 VDD2.n9 VSUBS 0.028524f
C227 VDD2.n10 VSUBS 0.016229f
C228 VDD2.n11 VSUBS 0.036228f
C229 VDD2.n12 VSUBS 0.016229f
C230 VDD2.n13 VSUBS 0.028524f
C231 VDD2.n14 VSUBS 0.015327f
C232 VDD2.n15 VSUBS 0.036228f
C233 VDD2.n16 VSUBS 0.016229f
C234 VDD2.n17 VSUBS 1.33395f
C235 VDD2.n18 VSUBS 0.015327f
C236 VDD2.t0 VSUBS 0.078021f
C237 VDD2.n19 VSUBS 0.21768f
C238 VDD2.n20 VSUBS 0.027253f
C239 VDD2.n21 VSUBS 0.027171f
C240 VDD2.n22 VSUBS 0.036228f
C241 VDD2.n23 VSUBS 0.016229f
C242 VDD2.n24 VSUBS 0.015327f
C243 VDD2.n25 VSUBS 0.028524f
C244 VDD2.n26 VSUBS 0.028524f
C245 VDD2.n27 VSUBS 0.015327f
C246 VDD2.n28 VSUBS 0.016229f
C247 VDD2.n29 VSUBS 0.036228f
C248 VDD2.n30 VSUBS 0.036228f
C249 VDD2.n31 VSUBS 0.016229f
C250 VDD2.n32 VSUBS 0.015327f
C251 VDD2.n33 VSUBS 0.028524f
C252 VDD2.n34 VSUBS 0.028524f
C253 VDD2.n35 VSUBS 0.015327f
C254 VDD2.n36 VSUBS 0.015327f
C255 VDD2.n37 VSUBS 0.016229f
C256 VDD2.n38 VSUBS 0.036228f
C257 VDD2.n39 VSUBS 0.036228f
C258 VDD2.n40 VSUBS 0.036228f
C259 VDD2.n41 VSUBS 0.015778f
C260 VDD2.n42 VSUBS 0.015327f
C261 VDD2.n43 VSUBS 0.028524f
C262 VDD2.n44 VSUBS 0.028524f
C263 VDD2.n45 VSUBS 0.015327f
C264 VDD2.n46 VSUBS 0.016229f
C265 VDD2.n47 VSUBS 0.036228f
C266 VDD2.n48 VSUBS 0.036228f
C267 VDD2.n49 VSUBS 0.016229f
C268 VDD2.n50 VSUBS 0.015327f
C269 VDD2.n51 VSUBS 0.028524f
C270 VDD2.n52 VSUBS 0.028524f
C271 VDD2.n53 VSUBS 0.015327f
C272 VDD2.n54 VSUBS 0.016229f
C273 VDD2.n55 VSUBS 0.036228f
C274 VDD2.n56 VSUBS 0.088122f
C275 VDD2.n57 VSUBS 0.016229f
C276 VDD2.n58 VSUBS 0.015327f
C277 VDD2.n59 VSUBS 0.068269f
C278 VDD2.n60 VSUBS 0.075385f
C279 VDD2.t3 VSUBS 0.25831f
C280 VDD2.t1 VSUBS 0.25831f
C281 VDD2.n61 VSUBS 2.01197f
C282 VDD2.n62 VSUBS 3.61934f
C283 VDD2.n63 VSUBS 0.031464f
C284 VDD2.n64 VSUBS 0.028524f
C285 VDD2.n65 VSUBS 0.015327f
C286 VDD2.n66 VSUBS 0.036228f
C287 VDD2.n67 VSUBS 0.016229f
C288 VDD2.n68 VSUBS 0.028524f
C289 VDD2.n69 VSUBS 0.015327f
C290 VDD2.n70 VSUBS 0.036228f
C291 VDD2.n71 VSUBS 0.015778f
C292 VDD2.n72 VSUBS 0.028524f
C293 VDD2.n73 VSUBS 0.015778f
C294 VDD2.n74 VSUBS 0.015327f
C295 VDD2.n75 VSUBS 0.036228f
C296 VDD2.n76 VSUBS 0.036228f
C297 VDD2.n77 VSUBS 0.016229f
C298 VDD2.n78 VSUBS 0.028524f
C299 VDD2.n79 VSUBS 0.015327f
C300 VDD2.n80 VSUBS 0.036228f
C301 VDD2.n81 VSUBS 0.016229f
C302 VDD2.n82 VSUBS 1.33395f
C303 VDD2.n83 VSUBS 0.015327f
C304 VDD2.t2 VSUBS 0.078021f
C305 VDD2.n84 VSUBS 0.217679f
C306 VDD2.n85 VSUBS 0.027253f
C307 VDD2.n86 VSUBS 0.027171f
C308 VDD2.n87 VSUBS 0.036228f
C309 VDD2.n88 VSUBS 0.016229f
C310 VDD2.n89 VSUBS 0.015327f
C311 VDD2.n90 VSUBS 0.028524f
C312 VDD2.n91 VSUBS 0.028524f
C313 VDD2.n92 VSUBS 0.015327f
C314 VDD2.n93 VSUBS 0.016229f
C315 VDD2.n94 VSUBS 0.036228f
C316 VDD2.n95 VSUBS 0.036228f
C317 VDD2.n96 VSUBS 0.016229f
C318 VDD2.n97 VSUBS 0.015327f
C319 VDD2.n98 VSUBS 0.028524f
C320 VDD2.n99 VSUBS 0.028524f
C321 VDD2.n100 VSUBS 0.015327f
C322 VDD2.n101 VSUBS 0.016229f
C323 VDD2.n102 VSUBS 0.036228f
C324 VDD2.n103 VSUBS 0.036228f
C325 VDD2.n104 VSUBS 0.016229f
C326 VDD2.n105 VSUBS 0.015327f
C327 VDD2.n106 VSUBS 0.028524f
C328 VDD2.n107 VSUBS 0.028524f
C329 VDD2.n108 VSUBS 0.015327f
C330 VDD2.n109 VSUBS 0.016229f
C331 VDD2.n110 VSUBS 0.036228f
C332 VDD2.n111 VSUBS 0.036228f
C333 VDD2.n112 VSUBS 0.016229f
C334 VDD2.n113 VSUBS 0.015327f
C335 VDD2.n114 VSUBS 0.028524f
C336 VDD2.n115 VSUBS 0.028524f
C337 VDD2.n116 VSUBS 0.015327f
C338 VDD2.n117 VSUBS 0.016229f
C339 VDD2.n118 VSUBS 0.036228f
C340 VDD2.n119 VSUBS 0.088122f
C341 VDD2.n120 VSUBS 0.016229f
C342 VDD2.n121 VSUBS 0.015327f
C343 VDD2.n122 VSUBS 0.068269f
C344 VDD2.n123 VSUBS 0.064082f
C345 VDD2.n124 VSUBS 3.07262f
C346 VDD2.t4 VSUBS 0.25831f
C347 VDD2.t5 VSUBS 0.25831f
C348 VDD2.n125 VSUBS 2.01193f
C349 VTAIL.t10 VSUBS 0.26959f
C350 VTAIL.t8 VSUBS 0.26959f
C351 VTAIL.n0 VSUBS 1.93813f
C352 VTAIL.n1 VSUBS 0.933777f
C353 VTAIL.n2 VSUBS 0.032838f
C354 VTAIL.n3 VSUBS 0.029769f
C355 VTAIL.n4 VSUBS 0.015997f
C356 VTAIL.n5 VSUBS 0.03781f
C357 VTAIL.n6 VSUBS 0.016938f
C358 VTAIL.n7 VSUBS 0.029769f
C359 VTAIL.n8 VSUBS 0.015997f
C360 VTAIL.n9 VSUBS 0.03781f
C361 VTAIL.n10 VSUBS 0.016467f
C362 VTAIL.n11 VSUBS 0.029769f
C363 VTAIL.n12 VSUBS 0.016938f
C364 VTAIL.n13 VSUBS 0.03781f
C365 VTAIL.n14 VSUBS 0.016938f
C366 VTAIL.n15 VSUBS 0.029769f
C367 VTAIL.n16 VSUBS 0.015997f
C368 VTAIL.n17 VSUBS 0.03781f
C369 VTAIL.n18 VSUBS 0.016938f
C370 VTAIL.n19 VSUBS 1.3922f
C371 VTAIL.n20 VSUBS 0.015997f
C372 VTAIL.t0 VSUBS 0.081428f
C373 VTAIL.n21 VSUBS 0.227185f
C374 VTAIL.n22 VSUBS 0.028443f
C375 VTAIL.n23 VSUBS 0.028358f
C376 VTAIL.n24 VSUBS 0.03781f
C377 VTAIL.n25 VSUBS 0.016938f
C378 VTAIL.n26 VSUBS 0.015997f
C379 VTAIL.n27 VSUBS 0.029769f
C380 VTAIL.n28 VSUBS 0.029769f
C381 VTAIL.n29 VSUBS 0.015997f
C382 VTAIL.n30 VSUBS 0.016938f
C383 VTAIL.n31 VSUBS 0.03781f
C384 VTAIL.n32 VSUBS 0.03781f
C385 VTAIL.n33 VSUBS 0.016938f
C386 VTAIL.n34 VSUBS 0.015997f
C387 VTAIL.n35 VSUBS 0.029769f
C388 VTAIL.n36 VSUBS 0.029769f
C389 VTAIL.n37 VSUBS 0.015997f
C390 VTAIL.n38 VSUBS 0.015997f
C391 VTAIL.n39 VSUBS 0.016938f
C392 VTAIL.n40 VSUBS 0.03781f
C393 VTAIL.n41 VSUBS 0.03781f
C394 VTAIL.n42 VSUBS 0.03781f
C395 VTAIL.n43 VSUBS 0.016467f
C396 VTAIL.n44 VSUBS 0.015997f
C397 VTAIL.n45 VSUBS 0.029769f
C398 VTAIL.n46 VSUBS 0.029769f
C399 VTAIL.n47 VSUBS 0.015997f
C400 VTAIL.n48 VSUBS 0.016938f
C401 VTAIL.n49 VSUBS 0.03781f
C402 VTAIL.n50 VSUBS 0.03781f
C403 VTAIL.n51 VSUBS 0.016938f
C404 VTAIL.n52 VSUBS 0.015997f
C405 VTAIL.n53 VSUBS 0.029769f
C406 VTAIL.n54 VSUBS 0.029769f
C407 VTAIL.n55 VSUBS 0.015997f
C408 VTAIL.n56 VSUBS 0.016938f
C409 VTAIL.n57 VSUBS 0.03781f
C410 VTAIL.n58 VSUBS 0.09197f
C411 VTAIL.n59 VSUBS 0.016938f
C412 VTAIL.n60 VSUBS 0.015997f
C413 VTAIL.n61 VSUBS 0.07125f
C414 VTAIL.n62 VSUBS 0.046344f
C415 VTAIL.n63 VSUBS 0.513445f
C416 VTAIL.t5 VSUBS 0.26959f
C417 VTAIL.t2 VSUBS 0.26959f
C418 VTAIL.n64 VSUBS 1.93813f
C419 VTAIL.n65 VSUBS 2.89752f
C420 VTAIL.t6 VSUBS 0.26959f
C421 VTAIL.t7 VSUBS 0.26959f
C422 VTAIL.n66 VSUBS 1.93815f
C423 VTAIL.n67 VSUBS 2.8975f
C424 VTAIL.n68 VSUBS 0.032838f
C425 VTAIL.n69 VSUBS 0.029769f
C426 VTAIL.n70 VSUBS 0.015997f
C427 VTAIL.n71 VSUBS 0.03781f
C428 VTAIL.n72 VSUBS 0.016938f
C429 VTAIL.n73 VSUBS 0.029769f
C430 VTAIL.n74 VSUBS 0.015997f
C431 VTAIL.n75 VSUBS 0.03781f
C432 VTAIL.n76 VSUBS 0.016467f
C433 VTAIL.n77 VSUBS 0.029769f
C434 VTAIL.n78 VSUBS 0.016467f
C435 VTAIL.n79 VSUBS 0.015997f
C436 VTAIL.n80 VSUBS 0.03781f
C437 VTAIL.n81 VSUBS 0.03781f
C438 VTAIL.n82 VSUBS 0.016938f
C439 VTAIL.n83 VSUBS 0.029769f
C440 VTAIL.n84 VSUBS 0.015997f
C441 VTAIL.n85 VSUBS 0.03781f
C442 VTAIL.n86 VSUBS 0.016938f
C443 VTAIL.n87 VSUBS 1.3922f
C444 VTAIL.n88 VSUBS 0.015997f
C445 VTAIL.t11 VSUBS 0.081428f
C446 VTAIL.n89 VSUBS 0.227185f
C447 VTAIL.n90 VSUBS 0.028443f
C448 VTAIL.n91 VSUBS 0.028358f
C449 VTAIL.n92 VSUBS 0.03781f
C450 VTAIL.n93 VSUBS 0.016938f
C451 VTAIL.n94 VSUBS 0.015997f
C452 VTAIL.n95 VSUBS 0.029769f
C453 VTAIL.n96 VSUBS 0.029769f
C454 VTAIL.n97 VSUBS 0.015997f
C455 VTAIL.n98 VSUBS 0.016938f
C456 VTAIL.n99 VSUBS 0.03781f
C457 VTAIL.n100 VSUBS 0.03781f
C458 VTAIL.n101 VSUBS 0.016938f
C459 VTAIL.n102 VSUBS 0.015997f
C460 VTAIL.n103 VSUBS 0.029769f
C461 VTAIL.n104 VSUBS 0.029769f
C462 VTAIL.n105 VSUBS 0.015997f
C463 VTAIL.n106 VSUBS 0.016938f
C464 VTAIL.n107 VSUBS 0.03781f
C465 VTAIL.n108 VSUBS 0.03781f
C466 VTAIL.n109 VSUBS 0.016938f
C467 VTAIL.n110 VSUBS 0.015997f
C468 VTAIL.n111 VSUBS 0.029769f
C469 VTAIL.n112 VSUBS 0.029769f
C470 VTAIL.n113 VSUBS 0.015997f
C471 VTAIL.n114 VSUBS 0.016938f
C472 VTAIL.n115 VSUBS 0.03781f
C473 VTAIL.n116 VSUBS 0.03781f
C474 VTAIL.n117 VSUBS 0.016938f
C475 VTAIL.n118 VSUBS 0.015997f
C476 VTAIL.n119 VSUBS 0.029769f
C477 VTAIL.n120 VSUBS 0.029769f
C478 VTAIL.n121 VSUBS 0.015997f
C479 VTAIL.n122 VSUBS 0.016938f
C480 VTAIL.n123 VSUBS 0.03781f
C481 VTAIL.n124 VSUBS 0.09197f
C482 VTAIL.n125 VSUBS 0.016938f
C483 VTAIL.n126 VSUBS 0.015997f
C484 VTAIL.n127 VSUBS 0.07125f
C485 VTAIL.n128 VSUBS 0.046344f
C486 VTAIL.n129 VSUBS 0.513445f
C487 VTAIL.t1 VSUBS 0.26959f
C488 VTAIL.t4 VSUBS 0.26959f
C489 VTAIL.n130 VSUBS 1.93815f
C490 VTAIL.n131 VSUBS 1.14897f
C491 VTAIL.n132 VSUBS 0.032838f
C492 VTAIL.n133 VSUBS 0.029769f
C493 VTAIL.n134 VSUBS 0.015997f
C494 VTAIL.n135 VSUBS 0.03781f
C495 VTAIL.n136 VSUBS 0.016938f
C496 VTAIL.n137 VSUBS 0.029769f
C497 VTAIL.n138 VSUBS 0.015997f
C498 VTAIL.n139 VSUBS 0.03781f
C499 VTAIL.n140 VSUBS 0.016467f
C500 VTAIL.n141 VSUBS 0.029769f
C501 VTAIL.n142 VSUBS 0.016467f
C502 VTAIL.n143 VSUBS 0.015997f
C503 VTAIL.n144 VSUBS 0.03781f
C504 VTAIL.n145 VSUBS 0.03781f
C505 VTAIL.n146 VSUBS 0.016938f
C506 VTAIL.n147 VSUBS 0.029769f
C507 VTAIL.n148 VSUBS 0.015997f
C508 VTAIL.n149 VSUBS 0.03781f
C509 VTAIL.n150 VSUBS 0.016938f
C510 VTAIL.n151 VSUBS 1.3922f
C511 VTAIL.n152 VSUBS 0.015997f
C512 VTAIL.t3 VSUBS 0.081428f
C513 VTAIL.n153 VSUBS 0.227185f
C514 VTAIL.n154 VSUBS 0.028443f
C515 VTAIL.n155 VSUBS 0.028358f
C516 VTAIL.n156 VSUBS 0.03781f
C517 VTAIL.n157 VSUBS 0.016938f
C518 VTAIL.n158 VSUBS 0.015997f
C519 VTAIL.n159 VSUBS 0.029769f
C520 VTAIL.n160 VSUBS 0.029769f
C521 VTAIL.n161 VSUBS 0.015997f
C522 VTAIL.n162 VSUBS 0.016938f
C523 VTAIL.n163 VSUBS 0.03781f
C524 VTAIL.n164 VSUBS 0.03781f
C525 VTAIL.n165 VSUBS 0.016938f
C526 VTAIL.n166 VSUBS 0.015997f
C527 VTAIL.n167 VSUBS 0.029769f
C528 VTAIL.n168 VSUBS 0.029769f
C529 VTAIL.n169 VSUBS 0.015997f
C530 VTAIL.n170 VSUBS 0.016938f
C531 VTAIL.n171 VSUBS 0.03781f
C532 VTAIL.n172 VSUBS 0.03781f
C533 VTAIL.n173 VSUBS 0.016938f
C534 VTAIL.n174 VSUBS 0.015997f
C535 VTAIL.n175 VSUBS 0.029769f
C536 VTAIL.n176 VSUBS 0.029769f
C537 VTAIL.n177 VSUBS 0.015997f
C538 VTAIL.n178 VSUBS 0.016938f
C539 VTAIL.n179 VSUBS 0.03781f
C540 VTAIL.n180 VSUBS 0.03781f
C541 VTAIL.n181 VSUBS 0.016938f
C542 VTAIL.n182 VSUBS 0.015997f
C543 VTAIL.n183 VSUBS 0.029769f
C544 VTAIL.n184 VSUBS 0.029769f
C545 VTAIL.n185 VSUBS 0.015997f
C546 VTAIL.n186 VSUBS 0.016938f
C547 VTAIL.n187 VSUBS 0.03781f
C548 VTAIL.n188 VSUBS 0.09197f
C549 VTAIL.n189 VSUBS 0.016938f
C550 VTAIL.n190 VSUBS 0.015997f
C551 VTAIL.n191 VSUBS 0.07125f
C552 VTAIL.n192 VSUBS 0.046344f
C553 VTAIL.n193 VSUBS 1.9676f
C554 VTAIL.n194 VSUBS 0.032838f
C555 VTAIL.n195 VSUBS 0.029769f
C556 VTAIL.n196 VSUBS 0.015997f
C557 VTAIL.n197 VSUBS 0.03781f
C558 VTAIL.n198 VSUBS 0.016938f
C559 VTAIL.n199 VSUBS 0.029769f
C560 VTAIL.n200 VSUBS 0.015997f
C561 VTAIL.n201 VSUBS 0.03781f
C562 VTAIL.n202 VSUBS 0.016467f
C563 VTAIL.n203 VSUBS 0.029769f
C564 VTAIL.n204 VSUBS 0.016938f
C565 VTAIL.n205 VSUBS 0.03781f
C566 VTAIL.n206 VSUBS 0.016938f
C567 VTAIL.n207 VSUBS 0.029769f
C568 VTAIL.n208 VSUBS 0.015997f
C569 VTAIL.n209 VSUBS 0.03781f
C570 VTAIL.n210 VSUBS 0.016938f
C571 VTAIL.n211 VSUBS 1.3922f
C572 VTAIL.n212 VSUBS 0.015997f
C573 VTAIL.t9 VSUBS 0.081428f
C574 VTAIL.n213 VSUBS 0.227185f
C575 VTAIL.n214 VSUBS 0.028443f
C576 VTAIL.n215 VSUBS 0.028358f
C577 VTAIL.n216 VSUBS 0.03781f
C578 VTAIL.n217 VSUBS 0.016938f
C579 VTAIL.n218 VSUBS 0.015997f
C580 VTAIL.n219 VSUBS 0.029769f
C581 VTAIL.n220 VSUBS 0.029769f
C582 VTAIL.n221 VSUBS 0.015997f
C583 VTAIL.n222 VSUBS 0.016938f
C584 VTAIL.n223 VSUBS 0.03781f
C585 VTAIL.n224 VSUBS 0.03781f
C586 VTAIL.n225 VSUBS 0.016938f
C587 VTAIL.n226 VSUBS 0.015997f
C588 VTAIL.n227 VSUBS 0.029769f
C589 VTAIL.n228 VSUBS 0.029769f
C590 VTAIL.n229 VSUBS 0.015997f
C591 VTAIL.n230 VSUBS 0.015997f
C592 VTAIL.n231 VSUBS 0.016938f
C593 VTAIL.n232 VSUBS 0.03781f
C594 VTAIL.n233 VSUBS 0.03781f
C595 VTAIL.n234 VSUBS 0.03781f
C596 VTAIL.n235 VSUBS 0.016467f
C597 VTAIL.n236 VSUBS 0.015997f
C598 VTAIL.n237 VSUBS 0.029769f
C599 VTAIL.n238 VSUBS 0.029769f
C600 VTAIL.n239 VSUBS 0.015997f
C601 VTAIL.n240 VSUBS 0.016938f
C602 VTAIL.n241 VSUBS 0.03781f
C603 VTAIL.n242 VSUBS 0.03781f
C604 VTAIL.n243 VSUBS 0.016938f
C605 VTAIL.n244 VSUBS 0.015997f
C606 VTAIL.n245 VSUBS 0.029769f
C607 VTAIL.n246 VSUBS 0.029769f
C608 VTAIL.n247 VSUBS 0.015997f
C609 VTAIL.n248 VSUBS 0.016938f
C610 VTAIL.n249 VSUBS 0.03781f
C611 VTAIL.n250 VSUBS 0.09197f
C612 VTAIL.n251 VSUBS 0.016938f
C613 VTAIL.n252 VSUBS 0.015997f
C614 VTAIL.n253 VSUBS 0.07125f
C615 VTAIL.n254 VSUBS 0.046344f
C616 VTAIL.n255 VSUBS 1.88842f
C617 VN.t4 VSUBS 2.76896f
C618 VN.n0 VSUBS 1.08372f
C619 VN.n1 VSUBS 0.027492f
C620 VN.n2 VSUBS 0.022569f
C621 VN.n3 VSUBS 0.027492f
C622 VN.t2 VSUBS 2.76896f
C623 VN.n4 VSUBS 1.06749f
C624 VN.t5 VSUBS 3.09477f
C625 VN.n5 VSUBS 1.01874f
C626 VN.n6 VSUBS 0.320657f
C627 VN.n7 VSUBS 0.038783f
C628 VN.n8 VSUBS 0.051495f
C629 VN.n9 VSUBS 0.055596f
C630 VN.n10 VSUBS 0.027492f
C631 VN.n11 VSUBS 0.027492f
C632 VN.n12 VSUBS 0.027492f
C633 VN.n13 VSUBS 0.053946f
C634 VN.n14 VSUBS 0.051495f
C635 VN.n15 VSUBS 0.041834f
C636 VN.n16 VSUBS 0.044379f
C637 VN.n17 VSUBS 0.065262f
C638 VN.t3 VSUBS 2.76896f
C639 VN.n18 VSUBS 1.08372f
C640 VN.n19 VSUBS 0.027492f
C641 VN.n20 VSUBS 0.022569f
C642 VN.n21 VSUBS 0.027492f
C643 VN.t1 VSUBS 2.76896f
C644 VN.n22 VSUBS 1.06749f
C645 VN.t0 VSUBS 3.09477f
C646 VN.n23 VSUBS 1.01874f
C647 VN.n24 VSUBS 0.320657f
C648 VN.n25 VSUBS 0.038783f
C649 VN.n26 VSUBS 0.051495f
C650 VN.n27 VSUBS 0.055596f
C651 VN.n28 VSUBS 0.027492f
C652 VN.n29 VSUBS 0.027492f
C653 VN.n30 VSUBS 0.027492f
C654 VN.n31 VSUBS 0.053946f
C655 VN.n32 VSUBS 0.051495f
C656 VN.n33 VSUBS 0.041834f
C657 VN.n34 VSUBS 0.044379f
C658 VN.n35 VSUBS 1.61133f
C659 B.n0 VSUBS 0.005529f
C660 B.n1 VSUBS 0.005529f
C661 B.n2 VSUBS 0.008744f
C662 B.n3 VSUBS 0.008744f
C663 B.n4 VSUBS 0.008744f
C664 B.n5 VSUBS 0.008744f
C665 B.n6 VSUBS 0.008744f
C666 B.n7 VSUBS 0.008744f
C667 B.n8 VSUBS 0.008744f
C668 B.n9 VSUBS 0.008744f
C669 B.n10 VSUBS 0.008744f
C670 B.n11 VSUBS 0.008744f
C671 B.n12 VSUBS 0.008744f
C672 B.n13 VSUBS 0.008744f
C673 B.n14 VSUBS 0.008744f
C674 B.n15 VSUBS 0.008744f
C675 B.n16 VSUBS 0.008744f
C676 B.n17 VSUBS 0.008744f
C677 B.n18 VSUBS 0.008744f
C678 B.n19 VSUBS 0.008744f
C679 B.n20 VSUBS 0.008744f
C680 B.n21 VSUBS 0.008744f
C681 B.n22 VSUBS 0.008744f
C682 B.n23 VSUBS 0.008744f
C683 B.n24 VSUBS 0.008744f
C684 B.n25 VSUBS 0.008744f
C685 B.n26 VSUBS 0.008744f
C686 B.n27 VSUBS 0.020234f
C687 B.n28 VSUBS 0.008744f
C688 B.n29 VSUBS 0.008744f
C689 B.n30 VSUBS 0.008744f
C690 B.n31 VSUBS 0.008744f
C691 B.n32 VSUBS 0.008744f
C692 B.n33 VSUBS 0.008744f
C693 B.n34 VSUBS 0.008744f
C694 B.n35 VSUBS 0.008744f
C695 B.n36 VSUBS 0.008744f
C696 B.n37 VSUBS 0.008744f
C697 B.n38 VSUBS 0.008744f
C698 B.n39 VSUBS 0.008744f
C699 B.n40 VSUBS 0.008744f
C700 B.n41 VSUBS 0.008744f
C701 B.n42 VSUBS 0.008744f
C702 B.n43 VSUBS 0.008744f
C703 B.n44 VSUBS 0.008744f
C704 B.n45 VSUBS 0.008744f
C705 B.n46 VSUBS 0.008744f
C706 B.n47 VSUBS 0.008744f
C707 B.t5 VSUBS 0.248793f
C708 B.t4 VSUBS 0.29573f
C709 B.t3 VSUBS 2.14124f
C710 B.n48 VSUBS 0.472986f
C711 B.n49 VSUBS 0.308227f
C712 B.n50 VSUBS 0.008744f
C713 B.n51 VSUBS 0.008744f
C714 B.n52 VSUBS 0.008744f
C715 B.n53 VSUBS 0.008744f
C716 B.t8 VSUBS 0.248796f
C717 B.t7 VSUBS 0.295733f
C718 B.t6 VSUBS 2.14124f
C719 B.n54 VSUBS 0.472983f
C720 B.n55 VSUBS 0.308224f
C721 B.n56 VSUBS 0.020258f
C722 B.n57 VSUBS 0.008744f
C723 B.n58 VSUBS 0.008744f
C724 B.n59 VSUBS 0.008744f
C725 B.n60 VSUBS 0.008744f
C726 B.n61 VSUBS 0.008744f
C727 B.n62 VSUBS 0.008744f
C728 B.n63 VSUBS 0.008744f
C729 B.n64 VSUBS 0.008744f
C730 B.n65 VSUBS 0.008744f
C731 B.n66 VSUBS 0.008744f
C732 B.n67 VSUBS 0.008744f
C733 B.n68 VSUBS 0.008744f
C734 B.n69 VSUBS 0.008744f
C735 B.n70 VSUBS 0.008744f
C736 B.n71 VSUBS 0.008744f
C737 B.n72 VSUBS 0.008744f
C738 B.n73 VSUBS 0.008744f
C739 B.n74 VSUBS 0.008744f
C740 B.n75 VSUBS 0.008744f
C741 B.n76 VSUBS 0.019125f
C742 B.n77 VSUBS 0.008744f
C743 B.n78 VSUBS 0.008744f
C744 B.n79 VSUBS 0.008744f
C745 B.n80 VSUBS 0.008744f
C746 B.n81 VSUBS 0.008744f
C747 B.n82 VSUBS 0.008744f
C748 B.n83 VSUBS 0.008744f
C749 B.n84 VSUBS 0.008744f
C750 B.n85 VSUBS 0.008744f
C751 B.n86 VSUBS 0.008744f
C752 B.n87 VSUBS 0.008744f
C753 B.n88 VSUBS 0.008744f
C754 B.n89 VSUBS 0.008744f
C755 B.n90 VSUBS 0.008744f
C756 B.n91 VSUBS 0.008744f
C757 B.n92 VSUBS 0.008744f
C758 B.n93 VSUBS 0.008744f
C759 B.n94 VSUBS 0.008744f
C760 B.n95 VSUBS 0.008744f
C761 B.n96 VSUBS 0.008744f
C762 B.n97 VSUBS 0.008744f
C763 B.n98 VSUBS 0.008744f
C764 B.n99 VSUBS 0.008744f
C765 B.n100 VSUBS 0.008744f
C766 B.n101 VSUBS 0.008744f
C767 B.n102 VSUBS 0.008744f
C768 B.n103 VSUBS 0.008744f
C769 B.n104 VSUBS 0.008744f
C770 B.n105 VSUBS 0.008744f
C771 B.n106 VSUBS 0.008744f
C772 B.n107 VSUBS 0.008744f
C773 B.n108 VSUBS 0.008744f
C774 B.n109 VSUBS 0.008744f
C775 B.n110 VSUBS 0.008744f
C776 B.n111 VSUBS 0.008744f
C777 B.n112 VSUBS 0.008744f
C778 B.n113 VSUBS 0.008744f
C779 B.n114 VSUBS 0.008744f
C780 B.n115 VSUBS 0.008744f
C781 B.n116 VSUBS 0.008744f
C782 B.n117 VSUBS 0.008744f
C783 B.n118 VSUBS 0.008744f
C784 B.n119 VSUBS 0.008744f
C785 B.n120 VSUBS 0.008744f
C786 B.n121 VSUBS 0.008744f
C787 B.n122 VSUBS 0.008744f
C788 B.n123 VSUBS 0.008744f
C789 B.n124 VSUBS 0.008744f
C790 B.n125 VSUBS 0.008744f
C791 B.n126 VSUBS 0.008744f
C792 B.n127 VSUBS 0.020234f
C793 B.n128 VSUBS 0.008744f
C794 B.n129 VSUBS 0.008744f
C795 B.n130 VSUBS 0.008744f
C796 B.n131 VSUBS 0.008744f
C797 B.n132 VSUBS 0.008744f
C798 B.n133 VSUBS 0.008744f
C799 B.n134 VSUBS 0.008744f
C800 B.n135 VSUBS 0.008744f
C801 B.n136 VSUBS 0.008744f
C802 B.n137 VSUBS 0.008744f
C803 B.n138 VSUBS 0.008744f
C804 B.n139 VSUBS 0.008744f
C805 B.n140 VSUBS 0.008744f
C806 B.n141 VSUBS 0.008744f
C807 B.n142 VSUBS 0.008744f
C808 B.n143 VSUBS 0.008744f
C809 B.n144 VSUBS 0.008744f
C810 B.n145 VSUBS 0.008744f
C811 B.n146 VSUBS 0.008744f
C812 B.n147 VSUBS 0.008744f
C813 B.t10 VSUBS 0.248796f
C814 B.t11 VSUBS 0.295733f
C815 B.t9 VSUBS 2.14124f
C816 B.n148 VSUBS 0.472983f
C817 B.n149 VSUBS 0.308224f
C818 B.n150 VSUBS 0.008744f
C819 B.n151 VSUBS 0.008744f
C820 B.n152 VSUBS 0.008744f
C821 B.n153 VSUBS 0.008744f
C822 B.t1 VSUBS 0.248793f
C823 B.t2 VSUBS 0.29573f
C824 B.t0 VSUBS 2.14124f
C825 B.n154 VSUBS 0.472986f
C826 B.n155 VSUBS 0.308227f
C827 B.n156 VSUBS 0.020258f
C828 B.n157 VSUBS 0.008744f
C829 B.n158 VSUBS 0.008744f
C830 B.n159 VSUBS 0.008744f
C831 B.n160 VSUBS 0.008744f
C832 B.n161 VSUBS 0.008744f
C833 B.n162 VSUBS 0.008744f
C834 B.n163 VSUBS 0.008744f
C835 B.n164 VSUBS 0.008744f
C836 B.n165 VSUBS 0.008744f
C837 B.n166 VSUBS 0.008744f
C838 B.n167 VSUBS 0.008744f
C839 B.n168 VSUBS 0.008744f
C840 B.n169 VSUBS 0.008744f
C841 B.n170 VSUBS 0.008744f
C842 B.n171 VSUBS 0.008744f
C843 B.n172 VSUBS 0.008744f
C844 B.n173 VSUBS 0.008744f
C845 B.n174 VSUBS 0.008744f
C846 B.n175 VSUBS 0.008744f
C847 B.n176 VSUBS 0.020234f
C848 B.n177 VSUBS 0.008744f
C849 B.n178 VSUBS 0.008744f
C850 B.n179 VSUBS 0.008744f
C851 B.n180 VSUBS 0.008744f
C852 B.n181 VSUBS 0.008744f
C853 B.n182 VSUBS 0.008744f
C854 B.n183 VSUBS 0.008744f
C855 B.n184 VSUBS 0.008744f
C856 B.n185 VSUBS 0.008744f
C857 B.n186 VSUBS 0.008744f
C858 B.n187 VSUBS 0.008744f
C859 B.n188 VSUBS 0.008744f
C860 B.n189 VSUBS 0.008744f
C861 B.n190 VSUBS 0.008744f
C862 B.n191 VSUBS 0.008744f
C863 B.n192 VSUBS 0.008744f
C864 B.n193 VSUBS 0.008744f
C865 B.n194 VSUBS 0.008744f
C866 B.n195 VSUBS 0.008744f
C867 B.n196 VSUBS 0.008744f
C868 B.n197 VSUBS 0.008744f
C869 B.n198 VSUBS 0.008744f
C870 B.n199 VSUBS 0.008744f
C871 B.n200 VSUBS 0.008744f
C872 B.n201 VSUBS 0.008744f
C873 B.n202 VSUBS 0.008744f
C874 B.n203 VSUBS 0.008744f
C875 B.n204 VSUBS 0.008744f
C876 B.n205 VSUBS 0.008744f
C877 B.n206 VSUBS 0.008744f
C878 B.n207 VSUBS 0.008744f
C879 B.n208 VSUBS 0.008744f
C880 B.n209 VSUBS 0.008744f
C881 B.n210 VSUBS 0.008744f
C882 B.n211 VSUBS 0.008744f
C883 B.n212 VSUBS 0.008744f
C884 B.n213 VSUBS 0.008744f
C885 B.n214 VSUBS 0.008744f
C886 B.n215 VSUBS 0.008744f
C887 B.n216 VSUBS 0.008744f
C888 B.n217 VSUBS 0.008744f
C889 B.n218 VSUBS 0.008744f
C890 B.n219 VSUBS 0.008744f
C891 B.n220 VSUBS 0.008744f
C892 B.n221 VSUBS 0.008744f
C893 B.n222 VSUBS 0.008744f
C894 B.n223 VSUBS 0.008744f
C895 B.n224 VSUBS 0.008744f
C896 B.n225 VSUBS 0.008744f
C897 B.n226 VSUBS 0.008744f
C898 B.n227 VSUBS 0.008744f
C899 B.n228 VSUBS 0.008744f
C900 B.n229 VSUBS 0.008744f
C901 B.n230 VSUBS 0.008744f
C902 B.n231 VSUBS 0.008744f
C903 B.n232 VSUBS 0.008744f
C904 B.n233 VSUBS 0.008744f
C905 B.n234 VSUBS 0.008744f
C906 B.n235 VSUBS 0.008744f
C907 B.n236 VSUBS 0.008744f
C908 B.n237 VSUBS 0.008744f
C909 B.n238 VSUBS 0.008744f
C910 B.n239 VSUBS 0.008744f
C911 B.n240 VSUBS 0.008744f
C912 B.n241 VSUBS 0.008744f
C913 B.n242 VSUBS 0.008744f
C914 B.n243 VSUBS 0.008744f
C915 B.n244 VSUBS 0.008744f
C916 B.n245 VSUBS 0.008744f
C917 B.n246 VSUBS 0.008744f
C918 B.n247 VSUBS 0.008744f
C919 B.n248 VSUBS 0.008744f
C920 B.n249 VSUBS 0.008744f
C921 B.n250 VSUBS 0.008744f
C922 B.n251 VSUBS 0.008744f
C923 B.n252 VSUBS 0.008744f
C924 B.n253 VSUBS 0.008744f
C925 B.n254 VSUBS 0.008744f
C926 B.n255 VSUBS 0.008744f
C927 B.n256 VSUBS 0.008744f
C928 B.n257 VSUBS 0.008744f
C929 B.n258 VSUBS 0.008744f
C930 B.n259 VSUBS 0.008744f
C931 B.n260 VSUBS 0.008744f
C932 B.n261 VSUBS 0.008744f
C933 B.n262 VSUBS 0.008744f
C934 B.n263 VSUBS 0.008744f
C935 B.n264 VSUBS 0.008744f
C936 B.n265 VSUBS 0.008744f
C937 B.n266 VSUBS 0.008744f
C938 B.n267 VSUBS 0.008744f
C939 B.n268 VSUBS 0.008744f
C940 B.n269 VSUBS 0.008744f
C941 B.n270 VSUBS 0.008744f
C942 B.n271 VSUBS 0.008744f
C943 B.n272 VSUBS 0.008744f
C944 B.n273 VSUBS 0.018855f
C945 B.n274 VSUBS 0.018855f
C946 B.n275 VSUBS 0.020234f
C947 B.n276 VSUBS 0.008744f
C948 B.n277 VSUBS 0.008744f
C949 B.n278 VSUBS 0.008744f
C950 B.n279 VSUBS 0.008744f
C951 B.n280 VSUBS 0.008744f
C952 B.n281 VSUBS 0.008744f
C953 B.n282 VSUBS 0.008744f
C954 B.n283 VSUBS 0.008744f
C955 B.n284 VSUBS 0.008744f
C956 B.n285 VSUBS 0.008744f
C957 B.n286 VSUBS 0.008744f
C958 B.n287 VSUBS 0.008744f
C959 B.n288 VSUBS 0.008744f
C960 B.n289 VSUBS 0.008744f
C961 B.n290 VSUBS 0.008744f
C962 B.n291 VSUBS 0.008744f
C963 B.n292 VSUBS 0.008744f
C964 B.n293 VSUBS 0.008744f
C965 B.n294 VSUBS 0.008744f
C966 B.n295 VSUBS 0.008744f
C967 B.n296 VSUBS 0.008744f
C968 B.n297 VSUBS 0.008744f
C969 B.n298 VSUBS 0.008744f
C970 B.n299 VSUBS 0.008744f
C971 B.n300 VSUBS 0.008744f
C972 B.n301 VSUBS 0.008744f
C973 B.n302 VSUBS 0.008744f
C974 B.n303 VSUBS 0.008744f
C975 B.n304 VSUBS 0.008744f
C976 B.n305 VSUBS 0.008744f
C977 B.n306 VSUBS 0.008744f
C978 B.n307 VSUBS 0.008744f
C979 B.n308 VSUBS 0.008744f
C980 B.n309 VSUBS 0.008744f
C981 B.n310 VSUBS 0.008744f
C982 B.n311 VSUBS 0.008744f
C983 B.n312 VSUBS 0.008744f
C984 B.n313 VSUBS 0.008744f
C985 B.n314 VSUBS 0.008744f
C986 B.n315 VSUBS 0.008744f
C987 B.n316 VSUBS 0.008744f
C988 B.n317 VSUBS 0.008744f
C989 B.n318 VSUBS 0.008744f
C990 B.n319 VSUBS 0.008744f
C991 B.n320 VSUBS 0.008744f
C992 B.n321 VSUBS 0.008744f
C993 B.n322 VSUBS 0.008744f
C994 B.n323 VSUBS 0.008744f
C995 B.n324 VSUBS 0.008744f
C996 B.n325 VSUBS 0.008744f
C997 B.n326 VSUBS 0.008744f
C998 B.n327 VSUBS 0.008744f
C999 B.n328 VSUBS 0.008744f
C1000 B.n329 VSUBS 0.008744f
C1001 B.n330 VSUBS 0.008744f
C1002 B.n331 VSUBS 0.008744f
C1003 B.n332 VSUBS 0.008744f
C1004 B.n333 VSUBS 0.008229f
C1005 B.n334 VSUBS 0.008744f
C1006 B.n335 VSUBS 0.008744f
C1007 B.n336 VSUBS 0.004886f
C1008 B.n337 VSUBS 0.008744f
C1009 B.n338 VSUBS 0.008744f
C1010 B.n339 VSUBS 0.008744f
C1011 B.n340 VSUBS 0.008744f
C1012 B.n341 VSUBS 0.008744f
C1013 B.n342 VSUBS 0.008744f
C1014 B.n343 VSUBS 0.008744f
C1015 B.n344 VSUBS 0.008744f
C1016 B.n345 VSUBS 0.008744f
C1017 B.n346 VSUBS 0.008744f
C1018 B.n347 VSUBS 0.008744f
C1019 B.n348 VSUBS 0.008744f
C1020 B.n349 VSUBS 0.004886f
C1021 B.n350 VSUBS 0.020258f
C1022 B.n351 VSUBS 0.008229f
C1023 B.n352 VSUBS 0.008744f
C1024 B.n353 VSUBS 0.008744f
C1025 B.n354 VSUBS 0.008744f
C1026 B.n355 VSUBS 0.008744f
C1027 B.n356 VSUBS 0.008744f
C1028 B.n357 VSUBS 0.008744f
C1029 B.n358 VSUBS 0.008744f
C1030 B.n359 VSUBS 0.008744f
C1031 B.n360 VSUBS 0.008744f
C1032 B.n361 VSUBS 0.008744f
C1033 B.n362 VSUBS 0.008744f
C1034 B.n363 VSUBS 0.008744f
C1035 B.n364 VSUBS 0.008744f
C1036 B.n365 VSUBS 0.008744f
C1037 B.n366 VSUBS 0.008744f
C1038 B.n367 VSUBS 0.008744f
C1039 B.n368 VSUBS 0.008744f
C1040 B.n369 VSUBS 0.008744f
C1041 B.n370 VSUBS 0.008744f
C1042 B.n371 VSUBS 0.008744f
C1043 B.n372 VSUBS 0.008744f
C1044 B.n373 VSUBS 0.008744f
C1045 B.n374 VSUBS 0.008744f
C1046 B.n375 VSUBS 0.008744f
C1047 B.n376 VSUBS 0.008744f
C1048 B.n377 VSUBS 0.008744f
C1049 B.n378 VSUBS 0.008744f
C1050 B.n379 VSUBS 0.008744f
C1051 B.n380 VSUBS 0.008744f
C1052 B.n381 VSUBS 0.008744f
C1053 B.n382 VSUBS 0.008744f
C1054 B.n383 VSUBS 0.008744f
C1055 B.n384 VSUBS 0.008744f
C1056 B.n385 VSUBS 0.008744f
C1057 B.n386 VSUBS 0.008744f
C1058 B.n387 VSUBS 0.008744f
C1059 B.n388 VSUBS 0.008744f
C1060 B.n389 VSUBS 0.008744f
C1061 B.n390 VSUBS 0.008744f
C1062 B.n391 VSUBS 0.008744f
C1063 B.n392 VSUBS 0.008744f
C1064 B.n393 VSUBS 0.008744f
C1065 B.n394 VSUBS 0.008744f
C1066 B.n395 VSUBS 0.008744f
C1067 B.n396 VSUBS 0.008744f
C1068 B.n397 VSUBS 0.008744f
C1069 B.n398 VSUBS 0.008744f
C1070 B.n399 VSUBS 0.008744f
C1071 B.n400 VSUBS 0.008744f
C1072 B.n401 VSUBS 0.008744f
C1073 B.n402 VSUBS 0.008744f
C1074 B.n403 VSUBS 0.008744f
C1075 B.n404 VSUBS 0.008744f
C1076 B.n405 VSUBS 0.008744f
C1077 B.n406 VSUBS 0.008744f
C1078 B.n407 VSUBS 0.008744f
C1079 B.n408 VSUBS 0.008744f
C1080 B.n409 VSUBS 0.008744f
C1081 B.n410 VSUBS 0.020234f
C1082 B.n411 VSUBS 0.018855f
C1083 B.n412 VSUBS 0.018855f
C1084 B.n413 VSUBS 0.008744f
C1085 B.n414 VSUBS 0.008744f
C1086 B.n415 VSUBS 0.008744f
C1087 B.n416 VSUBS 0.008744f
C1088 B.n417 VSUBS 0.008744f
C1089 B.n418 VSUBS 0.008744f
C1090 B.n419 VSUBS 0.008744f
C1091 B.n420 VSUBS 0.008744f
C1092 B.n421 VSUBS 0.008744f
C1093 B.n422 VSUBS 0.008744f
C1094 B.n423 VSUBS 0.008744f
C1095 B.n424 VSUBS 0.008744f
C1096 B.n425 VSUBS 0.008744f
C1097 B.n426 VSUBS 0.008744f
C1098 B.n427 VSUBS 0.008744f
C1099 B.n428 VSUBS 0.008744f
C1100 B.n429 VSUBS 0.008744f
C1101 B.n430 VSUBS 0.008744f
C1102 B.n431 VSUBS 0.008744f
C1103 B.n432 VSUBS 0.008744f
C1104 B.n433 VSUBS 0.008744f
C1105 B.n434 VSUBS 0.008744f
C1106 B.n435 VSUBS 0.008744f
C1107 B.n436 VSUBS 0.008744f
C1108 B.n437 VSUBS 0.008744f
C1109 B.n438 VSUBS 0.008744f
C1110 B.n439 VSUBS 0.008744f
C1111 B.n440 VSUBS 0.008744f
C1112 B.n441 VSUBS 0.008744f
C1113 B.n442 VSUBS 0.008744f
C1114 B.n443 VSUBS 0.008744f
C1115 B.n444 VSUBS 0.008744f
C1116 B.n445 VSUBS 0.008744f
C1117 B.n446 VSUBS 0.008744f
C1118 B.n447 VSUBS 0.008744f
C1119 B.n448 VSUBS 0.008744f
C1120 B.n449 VSUBS 0.008744f
C1121 B.n450 VSUBS 0.008744f
C1122 B.n451 VSUBS 0.008744f
C1123 B.n452 VSUBS 0.008744f
C1124 B.n453 VSUBS 0.008744f
C1125 B.n454 VSUBS 0.008744f
C1126 B.n455 VSUBS 0.008744f
C1127 B.n456 VSUBS 0.008744f
C1128 B.n457 VSUBS 0.008744f
C1129 B.n458 VSUBS 0.008744f
C1130 B.n459 VSUBS 0.008744f
C1131 B.n460 VSUBS 0.008744f
C1132 B.n461 VSUBS 0.008744f
C1133 B.n462 VSUBS 0.008744f
C1134 B.n463 VSUBS 0.008744f
C1135 B.n464 VSUBS 0.008744f
C1136 B.n465 VSUBS 0.008744f
C1137 B.n466 VSUBS 0.008744f
C1138 B.n467 VSUBS 0.008744f
C1139 B.n468 VSUBS 0.008744f
C1140 B.n469 VSUBS 0.008744f
C1141 B.n470 VSUBS 0.008744f
C1142 B.n471 VSUBS 0.008744f
C1143 B.n472 VSUBS 0.008744f
C1144 B.n473 VSUBS 0.008744f
C1145 B.n474 VSUBS 0.008744f
C1146 B.n475 VSUBS 0.008744f
C1147 B.n476 VSUBS 0.008744f
C1148 B.n477 VSUBS 0.008744f
C1149 B.n478 VSUBS 0.008744f
C1150 B.n479 VSUBS 0.008744f
C1151 B.n480 VSUBS 0.008744f
C1152 B.n481 VSUBS 0.008744f
C1153 B.n482 VSUBS 0.008744f
C1154 B.n483 VSUBS 0.008744f
C1155 B.n484 VSUBS 0.008744f
C1156 B.n485 VSUBS 0.008744f
C1157 B.n486 VSUBS 0.008744f
C1158 B.n487 VSUBS 0.008744f
C1159 B.n488 VSUBS 0.008744f
C1160 B.n489 VSUBS 0.008744f
C1161 B.n490 VSUBS 0.008744f
C1162 B.n491 VSUBS 0.008744f
C1163 B.n492 VSUBS 0.008744f
C1164 B.n493 VSUBS 0.008744f
C1165 B.n494 VSUBS 0.008744f
C1166 B.n495 VSUBS 0.008744f
C1167 B.n496 VSUBS 0.008744f
C1168 B.n497 VSUBS 0.008744f
C1169 B.n498 VSUBS 0.008744f
C1170 B.n499 VSUBS 0.008744f
C1171 B.n500 VSUBS 0.008744f
C1172 B.n501 VSUBS 0.008744f
C1173 B.n502 VSUBS 0.008744f
C1174 B.n503 VSUBS 0.008744f
C1175 B.n504 VSUBS 0.008744f
C1176 B.n505 VSUBS 0.008744f
C1177 B.n506 VSUBS 0.008744f
C1178 B.n507 VSUBS 0.008744f
C1179 B.n508 VSUBS 0.008744f
C1180 B.n509 VSUBS 0.008744f
C1181 B.n510 VSUBS 0.008744f
C1182 B.n511 VSUBS 0.008744f
C1183 B.n512 VSUBS 0.008744f
C1184 B.n513 VSUBS 0.008744f
C1185 B.n514 VSUBS 0.008744f
C1186 B.n515 VSUBS 0.008744f
C1187 B.n516 VSUBS 0.008744f
C1188 B.n517 VSUBS 0.008744f
C1189 B.n518 VSUBS 0.008744f
C1190 B.n519 VSUBS 0.008744f
C1191 B.n520 VSUBS 0.008744f
C1192 B.n521 VSUBS 0.008744f
C1193 B.n522 VSUBS 0.008744f
C1194 B.n523 VSUBS 0.008744f
C1195 B.n524 VSUBS 0.008744f
C1196 B.n525 VSUBS 0.008744f
C1197 B.n526 VSUBS 0.008744f
C1198 B.n527 VSUBS 0.008744f
C1199 B.n528 VSUBS 0.008744f
C1200 B.n529 VSUBS 0.008744f
C1201 B.n530 VSUBS 0.008744f
C1202 B.n531 VSUBS 0.008744f
C1203 B.n532 VSUBS 0.008744f
C1204 B.n533 VSUBS 0.008744f
C1205 B.n534 VSUBS 0.008744f
C1206 B.n535 VSUBS 0.008744f
C1207 B.n536 VSUBS 0.008744f
C1208 B.n537 VSUBS 0.008744f
C1209 B.n538 VSUBS 0.008744f
C1210 B.n539 VSUBS 0.008744f
C1211 B.n540 VSUBS 0.008744f
C1212 B.n541 VSUBS 0.008744f
C1213 B.n542 VSUBS 0.008744f
C1214 B.n543 VSUBS 0.008744f
C1215 B.n544 VSUBS 0.008744f
C1216 B.n545 VSUBS 0.008744f
C1217 B.n546 VSUBS 0.008744f
C1218 B.n547 VSUBS 0.008744f
C1219 B.n548 VSUBS 0.008744f
C1220 B.n549 VSUBS 0.008744f
C1221 B.n550 VSUBS 0.008744f
C1222 B.n551 VSUBS 0.008744f
C1223 B.n552 VSUBS 0.008744f
C1224 B.n553 VSUBS 0.008744f
C1225 B.n554 VSUBS 0.008744f
C1226 B.n555 VSUBS 0.008744f
C1227 B.n556 VSUBS 0.008744f
C1228 B.n557 VSUBS 0.008744f
C1229 B.n558 VSUBS 0.008744f
C1230 B.n559 VSUBS 0.008744f
C1231 B.n560 VSUBS 0.008744f
C1232 B.n561 VSUBS 0.019963f
C1233 B.n562 VSUBS 0.018855f
C1234 B.n563 VSUBS 0.020234f
C1235 B.n564 VSUBS 0.008744f
C1236 B.n565 VSUBS 0.008744f
C1237 B.n566 VSUBS 0.008744f
C1238 B.n567 VSUBS 0.008744f
C1239 B.n568 VSUBS 0.008744f
C1240 B.n569 VSUBS 0.008744f
C1241 B.n570 VSUBS 0.008744f
C1242 B.n571 VSUBS 0.008744f
C1243 B.n572 VSUBS 0.008744f
C1244 B.n573 VSUBS 0.008744f
C1245 B.n574 VSUBS 0.008744f
C1246 B.n575 VSUBS 0.008744f
C1247 B.n576 VSUBS 0.008744f
C1248 B.n577 VSUBS 0.008744f
C1249 B.n578 VSUBS 0.008744f
C1250 B.n579 VSUBS 0.008744f
C1251 B.n580 VSUBS 0.008744f
C1252 B.n581 VSUBS 0.008744f
C1253 B.n582 VSUBS 0.008744f
C1254 B.n583 VSUBS 0.008744f
C1255 B.n584 VSUBS 0.008744f
C1256 B.n585 VSUBS 0.008744f
C1257 B.n586 VSUBS 0.008744f
C1258 B.n587 VSUBS 0.008744f
C1259 B.n588 VSUBS 0.008744f
C1260 B.n589 VSUBS 0.008744f
C1261 B.n590 VSUBS 0.008744f
C1262 B.n591 VSUBS 0.008744f
C1263 B.n592 VSUBS 0.008744f
C1264 B.n593 VSUBS 0.008744f
C1265 B.n594 VSUBS 0.008744f
C1266 B.n595 VSUBS 0.008744f
C1267 B.n596 VSUBS 0.008744f
C1268 B.n597 VSUBS 0.008744f
C1269 B.n598 VSUBS 0.008744f
C1270 B.n599 VSUBS 0.008744f
C1271 B.n600 VSUBS 0.008744f
C1272 B.n601 VSUBS 0.008744f
C1273 B.n602 VSUBS 0.008744f
C1274 B.n603 VSUBS 0.008744f
C1275 B.n604 VSUBS 0.008744f
C1276 B.n605 VSUBS 0.008744f
C1277 B.n606 VSUBS 0.008744f
C1278 B.n607 VSUBS 0.008744f
C1279 B.n608 VSUBS 0.008744f
C1280 B.n609 VSUBS 0.008744f
C1281 B.n610 VSUBS 0.008744f
C1282 B.n611 VSUBS 0.008744f
C1283 B.n612 VSUBS 0.008744f
C1284 B.n613 VSUBS 0.008744f
C1285 B.n614 VSUBS 0.008744f
C1286 B.n615 VSUBS 0.008744f
C1287 B.n616 VSUBS 0.008744f
C1288 B.n617 VSUBS 0.008744f
C1289 B.n618 VSUBS 0.008744f
C1290 B.n619 VSUBS 0.008744f
C1291 B.n620 VSUBS 0.008744f
C1292 B.n621 VSUBS 0.008229f
C1293 B.n622 VSUBS 0.008744f
C1294 B.n623 VSUBS 0.008744f
C1295 B.n624 VSUBS 0.004886f
C1296 B.n625 VSUBS 0.008744f
C1297 B.n626 VSUBS 0.008744f
C1298 B.n627 VSUBS 0.008744f
C1299 B.n628 VSUBS 0.008744f
C1300 B.n629 VSUBS 0.008744f
C1301 B.n630 VSUBS 0.008744f
C1302 B.n631 VSUBS 0.008744f
C1303 B.n632 VSUBS 0.008744f
C1304 B.n633 VSUBS 0.008744f
C1305 B.n634 VSUBS 0.008744f
C1306 B.n635 VSUBS 0.008744f
C1307 B.n636 VSUBS 0.008744f
C1308 B.n637 VSUBS 0.004886f
C1309 B.n638 VSUBS 0.020258f
C1310 B.n639 VSUBS 0.008229f
C1311 B.n640 VSUBS 0.008744f
C1312 B.n641 VSUBS 0.008744f
C1313 B.n642 VSUBS 0.008744f
C1314 B.n643 VSUBS 0.008744f
C1315 B.n644 VSUBS 0.008744f
C1316 B.n645 VSUBS 0.008744f
C1317 B.n646 VSUBS 0.008744f
C1318 B.n647 VSUBS 0.008744f
C1319 B.n648 VSUBS 0.008744f
C1320 B.n649 VSUBS 0.008744f
C1321 B.n650 VSUBS 0.008744f
C1322 B.n651 VSUBS 0.008744f
C1323 B.n652 VSUBS 0.008744f
C1324 B.n653 VSUBS 0.008744f
C1325 B.n654 VSUBS 0.008744f
C1326 B.n655 VSUBS 0.008744f
C1327 B.n656 VSUBS 0.008744f
C1328 B.n657 VSUBS 0.008744f
C1329 B.n658 VSUBS 0.008744f
C1330 B.n659 VSUBS 0.008744f
C1331 B.n660 VSUBS 0.008744f
C1332 B.n661 VSUBS 0.008744f
C1333 B.n662 VSUBS 0.008744f
C1334 B.n663 VSUBS 0.008744f
C1335 B.n664 VSUBS 0.008744f
C1336 B.n665 VSUBS 0.008744f
C1337 B.n666 VSUBS 0.008744f
C1338 B.n667 VSUBS 0.008744f
C1339 B.n668 VSUBS 0.008744f
C1340 B.n669 VSUBS 0.008744f
C1341 B.n670 VSUBS 0.008744f
C1342 B.n671 VSUBS 0.008744f
C1343 B.n672 VSUBS 0.008744f
C1344 B.n673 VSUBS 0.008744f
C1345 B.n674 VSUBS 0.008744f
C1346 B.n675 VSUBS 0.008744f
C1347 B.n676 VSUBS 0.008744f
C1348 B.n677 VSUBS 0.008744f
C1349 B.n678 VSUBS 0.008744f
C1350 B.n679 VSUBS 0.008744f
C1351 B.n680 VSUBS 0.008744f
C1352 B.n681 VSUBS 0.008744f
C1353 B.n682 VSUBS 0.008744f
C1354 B.n683 VSUBS 0.008744f
C1355 B.n684 VSUBS 0.008744f
C1356 B.n685 VSUBS 0.008744f
C1357 B.n686 VSUBS 0.008744f
C1358 B.n687 VSUBS 0.008744f
C1359 B.n688 VSUBS 0.008744f
C1360 B.n689 VSUBS 0.008744f
C1361 B.n690 VSUBS 0.008744f
C1362 B.n691 VSUBS 0.008744f
C1363 B.n692 VSUBS 0.008744f
C1364 B.n693 VSUBS 0.008744f
C1365 B.n694 VSUBS 0.008744f
C1366 B.n695 VSUBS 0.008744f
C1367 B.n696 VSUBS 0.008744f
C1368 B.n697 VSUBS 0.008744f
C1369 B.n698 VSUBS 0.020234f
C1370 B.n699 VSUBS 0.018855f
C1371 B.n700 VSUBS 0.018855f
C1372 B.n701 VSUBS 0.008744f
C1373 B.n702 VSUBS 0.008744f
C1374 B.n703 VSUBS 0.008744f
C1375 B.n704 VSUBS 0.008744f
C1376 B.n705 VSUBS 0.008744f
C1377 B.n706 VSUBS 0.008744f
C1378 B.n707 VSUBS 0.008744f
C1379 B.n708 VSUBS 0.008744f
C1380 B.n709 VSUBS 0.008744f
C1381 B.n710 VSUBS 0.008744f
C1382 B.n711 VSUBS 0.008744f
C1383 B.n712 VSUBS 0.008744f
C1384 B.n713 VSUBS 0.008744f
C1385 B.n714 VSUBS 0.008744f
C1386 B.n715 VSUBS 0.008744f
C1387 B.n716 VSUBS 0.008744f
C1388 B.n717 VSUBS 0.008744f
C1389 B.n718 VSUBS 0.008744f
C1390 B.n719 VSUBS 0.008744f
C1391 B.n720 VSUBS 0.008744f
C1392 B.n721 VSUBS 0.008744f
C1393 B.n722 VSUBS 0.008744f
C1394 B.n723 VSUBS 0.008744f
C1395 B.n724 VSUBS 0.008744f
C1396 B.n725 VSUBS 0.008744f
C1397 B.n726 VSUBS 0.008744f
C1398 B.n727 VSUBS 0.008744f
C1399 B.n728 VSUBS 0.008744f
C1400 B.n729 VSUBS 0.008744f
C1401 B.n730 VSUBS 0.008744f
C1402 B.n731 VSUBS 0.008744f
C1403 B.n732 VSUBS 0.008744f
C1404 B.n733 VSUBS 0.008744f
C1405 B.n734 VSUBS 0.008744f
C1406 B.n735 VSUBS 0.008744f
C1407 B.n736 VSUBS 0.008744f
C1408 B.n737 VSUBS 0.008744f
C1409 B.n738 VSUBS 0.008744f
C1410 B.n739 VSUBS 0.008744f
C1411 B.n740 VSUBS 0.008744f
C1412 B.n741 VSUBS 0.008744f
C1413 B.n742 VSUBS 0.008744f
C1414 B.n743 VSUBS 0.008744f
C1415 B.n744 VSUBS 0.008744f
C1416 B.n745 VSUBS 0.008744f
C1417 B.n746 VSUBS 0.008744f
C1418 B.n747 VSUBS 0.008744f
C1419 B.n748 VSUBS 0.008744f
C1420 B.n749 VSUBS 0.008744f
C1421 B.n750 VSUBS 0.008744f
C1422 B.n751 VSUBS 0.008744f
C1423 B.n752 VSUBS 0.008744f
C1424 B.n753 VSUBS 0.008744f
C1425 B.n754 VSUBS 0.008744f
C1426 B.n755 VSUBS 0.008744f
C1427 B.n756 VSUBS 0.008744f
C1428 B.n757 VSUBS 0.008744f
C1429 B.n758 VSUBS 0.008744f
C1430 B.n759 VSUBS 0.008744f
C1431 B.n760 VSUBS 0.008744f
C1432 B.n761 VSUBS 0.008744f
C1433 B.n762 VSUBS 0.008744f
C1434 B.n763 VSUBS 0.008744f
C1435 B.n764 VSUBS 0.008744f
C1436 B.n765 VSUBS 0.008744f
C1437 B.n766 VSUBS 0.008744f
C1438 B.n767 VSUBS 0.008744f
C1439 B.n768 VSUBS 0.008744f
C1440 B.n769 VSUBS 0.008744f
C1441 B.n770 VSUBS 0.008744f
C1442 B.n771 VSUBS 0.008744f
C1443 B.n772 VSUBS 0.008744f
C1444 B.n773 VSUBS 0.008744f
C1445 B.n774 VSUBS 0.008744f
C1446 B.n775 VSUBS 0.019798f
.ends

