* NGSPICE file created from diff_pair_sample_1361.ext - technology: sky130A

.subckt diff_pair_sample_1361 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t13 VN.t0 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=1.6302 ps=10.21 w=9.88 l=0.48
X1 VDD1.t7 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=0 ps=0 w=9.88 l=0.48
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=0 ps=0 w=9.88 l=0.48
X4 VDD1.t6 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=3.8532 ps=20.54 w=9.88 l=0.48
X5 VDD1.t5 VP.t2 VTAIL.t14 B.t21 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X6 VTAIL.t12 VN.t1 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=0 ps=0 w=9.88 l=0.48
X8 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=1.6302 ps=10.21 w=9.88 l=0.48
X9 VTAIL.t0 VP.t4 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X10 VDD1.t2 VP.t5 VTAIL.t15 B.t20 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=3.8532 ps=20.54 w=9.88 l=0.48
X11 VTAIL.t2 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=1.6302 ps=10.21 w=9.88 l=0.48
X12 VDD2.t5 VN.t2 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=3.8532 ps=20.54 w=9.88 l=0.48
X13 VTAIL.t10 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=1.6302 ps=10.21 w=9.88 l=0.48
X14 VTAIL.t3 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X15 VTAIL.t9 VN.t4 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X16 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8532 pd=20.54 as=0 ps=0 w=9.88 l=0.48
X17 VDD2.t3 VN.t5 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X18 VDD2.t6 VN.t6 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=1.6302 ps=10.21 w=9.88 l=0.48
X19 VDD2.t2 VN.t7 VTAIL.t6 B.t20 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=10.21 as=3.8532 ps=20.54 w=9.88 l=0.48
R0 VN.n2 VN.t0 599.885
R1 VN.n10 VN.t2 599.885
R2 VN.n1 VN.t5 578.903
R3 VN.n5 VN.t4 578.903
R4 VN.n6 VN.t7 578.903
R5 VN.n9 VN.t1 578.903
R6 VN.n13 VN.t6 578.903
R7 VN.n14 VN.t3 578.903
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.4033
R15 VN.n3 VN.n2 70.4033
R16 VN.n6 VN.n5 48.2005
R17 VN.n14 VN.n13 48.2005
R18 VN VN.n15 39.813
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.9576
R24 VN.n2 VN.n1 20.9576
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VDD2.n2 VDD2.n1 61.3824
R31 VDD2.n2 VDD2.n0 61.3824
R32 VDD2 VDD2.n5 61.3796
R33 VDD2.n4 VDD2.n3 61.0888
R34 VDD2.n4 VDD2.n2 35.3748
R35 VDD2.n5 VDD2.t0 2.00455
R36 VDD2.n5 VDD2.t5 2.00455
R37 VDD2.n3 VDD2.t4 2.00455
R38 VDD2.n3 VDD2.t6 2.00455
R39 VDD2.n1 VDD2.t7 2.00455
R40 VDD2.n1 VDD2.t2 2.00455
R41 VDD2.n0 VDD2.t1 2.00455
R42 VDD2.n0 VDD2.t3 2.00455
R43 VDD2 VDD2.n4 0.407828
R44 VTAIL.n434 VTAIL.n386 289.615
R45 VTAIL.n50 VTAIL.n2 289.615
R46 VTAIL.n104 VTAIL.n56 289.615
R47 VTAIL.n160 VTAIL.n112 289.615
R48 VTAIL.n380 VTAIL.n332 289.615
R49 VTAIL.n324 VTAIL.n276 289.615
R50 VTAIL.n270 VTAIL.n222 289.615
R51 VTAIL.n214 VTAIL.n166 289.615
R52 VTAIL.n402 VTAIL.n401 185
R53 VTAIL.n407 VTAIL.n406 185
R54 VTAIL.n409 VTAIL.n408 185
R55 VTAIL.n398 VTAIL.n397 185
R56 VTAIL.n415 VTAIL.n414 185
R57 VTAIL.n417 VTAIL.n416 185
R58 VTAIL.n394 VTAIL.n393 185
R59 VTAIL.n424 VTAIL.n423 185
R60 VTAIL.n425 VTAIL.n392 185
R61 VTAIL.n427 VTAIL.n426 185
R62 VTAIL.n390 VTAIL.n389 185
R63 VTAIL.n433 VTAIL.n432 185
R64 VTAIL.n435 VTAIL.n434 185
R65 VTAIL.n18 VTAIL.n17 185
R66 VTAIL.n23 VTAIL.n22 185
R67 VTAIL.n25 VTAIL.n24 185
R68 VTAIL.n14 VTAIL.n13 185
R69 VTAIL.n31 VTAIL.n30 185
R70 VTAIL.n33 VTAIL.n32 185
R71 VTAIL.n10 VTAIL.n9 185
R72 VTAIL.n40 VTAIL.n39 185
R73 VTAIL.n41 VTAIL.n8 185
R74 VTAIL.n43 VTAIL.n42 185
R75 VTAIL.n6 VTAIL.n5 185
R76 VTAIL.n49 VTAIL.n48 185
R77 VTAIL.n51 VTAIL.n50 185
R78 VTAIL.n72 VTAIL.n71 185
R79 VTAIL.n77 VTAIL.n76 185
R80 VTAIL.n79 VTAIL.n78 185
R81 VTAIL.n68 VTAIL.n67 185
R82 VTAIL.n85 VTAIL.n84 185
R83 VTAIL.n87 VTAIL.n86 185
R84 VTAIL.n64 VTAIL.n63 185
R85 VTAIL.n94 VTAIL.n93 185
R86 VTAIL.n95 VTAIL.n62 185
R87 VTAIL.n97 VTAIL.n96 185
R88 VTAIL.n60 VTAIL.n59 185
R89 VTAIL.n103 VTAIL.n102 185
R90 VTAIL.n105 VTAIL.n104 185
R91 VTAIL.n128 VTAIL.n127 185
R92 VTAIL.n133 VTAIL.n132 185
R93 VTAIL.n135 VTAIL.n134 185
R94 VTAIL.n124 VTAIL.n123 185
R95 VTAIL.n141 VTAIL.n140 185
R96 VTAIL.n143 VTAIL.n142 185
R97 VTAIL.n120 VTAIL.n119 185
R98 VTAIL.n150 VTAIL.n149 185
R99 VTAIL.n151 VTAIL.n118 185
R100 VTAIL.n153 VTAIL.n152 185
R101 VTAIL.n116 VTAIL.n115 185
R102 VTAIL.n159 VTAIL.n158 185
R103 VTAIL.n161 VTAIL.n160 185
R104 VTAIL.n381 VTAIL.n380 185
R105 VTAIL.n379 VTAIL.n378 185
R106 VTAIL.n336 VTAIL.n335 185
R107 VTAIL.n373 VTAIL.n372 185
R108 VTAIL.n371 VTAIL.n338 185
R109 VTAIL.n370 VTAIL.n369 185
R110 VTAIL.n341 VTAIL.n339 185
R111 VTAIL.n364 VTAIL.n363 185
R112 VTAIL.n362 VTAIL.n361 185
R113 VTAIL.n345 VTAIL.n344 185
R114 VTAIL.n356 VTAIL.n355 185
R115 VTAIL.n354 VTAIL.n353 185
R116 VTAIL.n349 VTAIL.n348 185
R117 VTAIL.n325 VTAIL.n324 185
R118 VTAIL.n323 VTAIL.n322 185
R119 VTAIL.n280 VTAIL.n279 185
R120 VTAIL.n317 VTAIL.n316 185
R121 VTAIL.n315 VTAIL.n282 185
R122 VTAIL.n314 VTAIL.n313 185
R123 VTAIL.n285 VTAIL.n283 185
R124 VTAIL.n308 VTAIL.n307 185
R125 VTAIL.n306 VTAIL.n305 185
R126 VTAIL.n289 VTAIL.n288 185
R127 VTAIL.n300 VTAIL.n299 185
R128 VTAIL.n298 VTAIL.n297 185
R129 VTAIL.n293 VTAIL.n292 185
R130 VTAIL.n271 VTAIL.n270 185
R131 VTAIL.n269 VTAIL.n268 185
R132 VTAIL.n226 VTAIL.n225 185
R133 VTAIL.n263 VTAIL.n262 185
R134 VTAIL.n261 VTAIL.n228 185
R135 VTAIL.n260 VTAIL.n259 185
R136 VTAIL.n231 VTAIL.n229 185
R137 VTAIL.n254 VTAIL.n253 185
R138 VTAIL.n252 VTAIL.n251 185
R139 VTAIL.n235 VTAIL.n234 185
R140 VTAIL.n246 VTAIL.n245 185
R141 VTAIL.n244 VTAIL.n243 185
R142 VTAIL.n239 VTAIL.n238 185
R143 VTAIL.n215 VTAIL.n214 185
R144 VTAIL.n213 VTAIL.n212 185
R145 VTAIL.n170 VTAIL.n169 185
R146 VTAIL.n207 VTAIL.n206 185
R147 VTAIL.n205 VTAIL.n172 185
R148 VTAIL.n204 VTAIL.n203 185
R149 VTAIL.n175 VTAIL.n173 185
R150 VTAIL.n198 VTAIL.n197 185
R151 VTAIL.n196 VTAIL.n195 185
R152 VTAIL.n179 VTAIL.n178 185
R153 VTAIL.n190 VTAIL.n189 185
R154 VTAIL.n188 VTAIL.n187 185
R155 VTAIL.n183 VTAIL.n182 185
R156 VTAIL.n403 VTAIL.t6 149.524
R157 VTAIL.n19 VTAIL.t13 149.524
R158 VTAIL.n73 VTAIL.t1 149.524
R159 VTAIL.n129 VTAIL.t2 149.524
R160 VTAIL.n350 VTAIL.t15 149.524
R161 VTAIL.n294 VTAIL.t4 149.524
R162 VTAIL.n240 VTAIL.t11 149.524
R163 VTAIL.n184 VTAIL.t10 149.524
R164 VTAIL.n407 VTAIL.n401 104.615
R165 VTAIL.n408 VTAIL.n407 104.615
R166 VTAIL.n408 VTAIL.n397 104.615
R167 VTAIL.n415 VTAIL.n397 104.615
R168 VTAIL.n416 VTAIL.n415 104.615
R169 VTAIL.n416 VTAIL.n393 104.615
R170 VTAIL.n424 VTAIL.n393 104.615
R171 VTAIL.n425 VTAIL.n424 104.615
R172 VTAIL.n426 VTAIL.n425 104.615
R173 VTAIL.n426 VTAIL.n389 104.615
R174 VTAIL.n433 VTAIL.n389 104.615
R175 VTAIL.n434 VTAIL.n433 104.615
R176 VTAIL.n23 VTAIL.n17 104.615
R177 VTAIL.n24 VTAIL.n23 104.615
R178 VTAIL.n24 VTAIL.n13 104.615
R179 VTAIL.n31 VTAIL.n13 104.615
R180 VTAIL.n32 VTAIL.n31 104.615
R181 VTAIL.n32 VTAIL.n9 104.615
R182 VTAIL.n40 VTAIL.n9 104.615
R183 VTAIL.n41 VTAIL.n40 104.615
R184 VTAIL.n42 VTAIL.n41 104.615
R185 VTAIL.n42 VTAIL.n5 104.615
R186 VTAIL.n49 VTAIL.n5 104.615
R187 VTAIL.n50 VTAIL.n49 104.615
R188 VTAIL.n77 VTAIL.n71 104.615
R189 VTAIL.n78 VTAIL.n77 104.615
R190 VTAIL.n78 VTAIL.n67 104.615
R191 VTAIL.n85 VTAIL.n67 104.615
R192 VTAIL.n86 VTAIL.n85 104.615
R193 VTAIL.n86 VTAIL.n63 104.615
R194 VTAIL.n94 VTAIL.n63 104.615
R195 VTAIL.n95 VTAIL.n94 104.615
R196 VTAIL.n96 VTAIL.n95 104.615
R197 VTAIL.n96 VTAIL.n59 104.615
R198 VTAIL.n103 VTAIL.n59 104.615
R199 VTAIL.n104 VTAIL.n103 104.615
R200 VTAIL.n133 VTAIL.n127 104.615
R201 VTAIL.n134 VTAIL.n133 104.615
R202 VTAIL.n134 VTAIL.n123 104.615
R203 VTAIL.n141 VTAIL.n123 104.615
R204 VTAIL.n142 VTAIL.n141 104.615
R205 VTAIL.n142 VTAIL.n119 104.615
R206 VTAIL.n150 VTAIL.n119 104.615
R207 VTAIL.n151 VTAIL.n150 104.615
R208 VTAIL.n152 VTAIL.n151 104.615
R209 VTAIL.n152 VTAIL.n115 104.615
R210 VTAIL.n159 VTAIL.n115 104.615
R211 VTAIL.n160 VTAIL.n159 104.615
R212 VTAIL.n380 VTAIL.n379 104.615
R213 VTAIL.n379 VTAIL.n335 104.615
R214 VTAIL.n372 VTAIL.n335 104.615
R215 VTAIL.n372 VTAIL.n371 104.615
R216 VTAIL.n371 VTAIL.n370 104.615
R217 VTAIL.n370 VTAIL.n339 104.615
R218 VTAIL.n363 VTAIL.n339 104.615
R219 VTAIL.n363 VTAIL.n362 104.615
R220 VTAIL.n362 VTAIL.n344 104.615
R221 VTAIL.n355 VTAIL.n344 104.615
R222 VTAIL.n355 VTAIL.n354 104.615
R223 VTAIL.n354 VTAIL.n348 104.615
R224 VTAIL.n324 VTAIL.n323 104.615
R225 VTAIL.n323 VTAIL.n279 104.615
R226 VTAIL.n316 VTAIL.n279 104.615
R227 VTAIL.n316 VTAIL.n315 104.615
R228 VTAIL.n315 VTAIL.n314 104.615
R229 VTAIL.n314 VTAIL.n283 104.615
R230 VTAIL.n307 VTAIL.n283 104.615
R231 VTAIL.n307 VTAIL.n306 104.615
R232 VTAIL.n306 VTAIL.n288 104.615
R233 VTAIL.n299 VTAIL.n288 104.615
R234 VTAIL.n299 VTAIL.n298 104.615
R235 VTAIL.n298 VTAIL.n292 104.615
R236 VTAIL.n270 VTAIL.n269 104.615
R237 VTAIL.n269 VTAIL.n225 104.615
R238 VTAIL.n262 VTAIL.n225 104.615
R239 VTAIL.n262 VTAIL.n261 104.615
R240 VTAIL.n261 VTAIL.n260 104.615
R241 VTAIL.n260 VTAIL.n229 104.615
R242 VTAIL.n253 VTAIL.n229 104.615
R243 VTAIL.n253 VTAIL.n252 104.615
R244 VTAIL.n252 VTAIL.n234 104.615
R245 VTAIL.n245 VTAIL.n234 104.615
R246 VTAIL.n245 VTAIL.n244 104.615
R247 VTAIL.n244 VTAIL.n238 104.615
R248 VTAIL.n214 VTAIL.n213 104.615
R249 VTAIL.n213 VTAIL.n169 104.615
R250 VTAIL.n206 VTAIL.n169 104.615
R251 VTAIL.n206 VTAIL.n205 104.615
R252 VTAIL.n205 VTAIL.n204 104.615
R253 VTAIL.n204 VTAIL.n173 104.615
R254 VTAIL.n197 VTAIL.n173 104.615
R255 VTAIL.n197 VTAIL.n196 104.615
R256 VTAIL.n196 VTAIL.n178 104.615
R257 VTAIL.n189 VTAIL.n178 104.615
R258 VTAIL.n189 VTAIL.n188 104.615
R259 VTAIL.n188 VTAIL.n182 104.615
R260 VTAIL.t6 VTAIL.n401 52.3082
R261 VTAIL.t13 VTAIL.n17 52.3082
R262 VTAIL.t1 VTAIL.n71 52.3082
R263 VTAIL.t2 VTAIL.n127 52.3082
R264 VTAIL.t15 VTAIL.n348 52.3082
R265 VTAIL.t4 VTAIL.n292 52.3082
R266 VTAIL.t11 VTAIL.n238 52.3082
R267 VTAIL.t10 VTAIL.n182 52.3082
R268 VTAIL.n331 VTAIL.n330 44.41
R269 VTAIL.n221 VTAIL.n220 44.41
R270 VTAIL.n1 VTAIL.n0 44.4099
R271 VTAIL.n111 VTAIL.n110 44.4099
R272 VTAIL.n439 VTAIL.n438 30.6338
R273 VTAIL.n55 VTAIL.n54 30.6338
R274 VTAIL.n109 VTAIL.n108 30.6338
R275 VTAIL.n165 VTAIL.n164 30.6338
R276 VTAIL.n385 VTAIL.n384 30.6338
R277 VTAIL.n329 VTAIL.n328 30.6338
R278 VTAIL.n275 VTAIL.n274 30.6338
R279 VTAIL.n219 VTAIL.n218 30.6338
R280 VTAIL.n439 VTAIL.n385 21.5824
R281 VTAIL.n219 VTAIL.n165 21.5824
R282 VTAIL.n427 VTAIL.n392 13.1884
R283 VTAIL.n43 VTAIL.n8 13.1884
R284 VTAIL.n97 VTAIL.n62 13.1884
R285 VTAIL.n153 VTAIL.n118 13.1884
R286 VTAIL.n373 VTAIL.n338 13.1884
R287 VTAIL.n317 VTAIL.n282 13.1884
R288 VTAIL.n263 VTAIL.n228 13.1884
R289 VTAIL.n207 VTAIL.n172 13.1884
R290 VTAIL.n423 VTAIL.n422 12.8005
R291 VTAIL.n428 VTAIL.n390 12.8005
R292 VTAIL.n39 VTAIL.n38 12.8005
R293 VTAIL.n44 VTAIL.n6 12.8005
R294 VTAIL.n93 VTAIL.n92 12.8005
R295 VTAIL.n98 VTAIL.n60 12.8005
R296 VTAIL.n149 VTAIL.n148 12.8005
R297 VTAIL.n154 VTAIL.n116 12.8005
R298 VTAIL.n374 VTAIL.n336 12.8005
R299 VTAIL.n369 VTAIL.n340 12.8005
R300 VTAIL.n318 VTAIL.n280 12.8005
R301 VTAIL.n313 VTAIL.n284 12.8005
R302 VTAIL.n264 VTAIL.n226 12.8005
R303 VTAIL.n259 VTAIL.n230 12.8005
R304 VTAIL.n208 VTAIL.n170 12.8005
R305 VTAIL.n203 VTAIL.n174 12.8005
R306 VTAIL.n421 VTAIL.n394 12.0247
R307 VTAIL.n432 VTAIL.n431 12.0247
R308 VTAIL.n37 VTAIL.n10 12.0247
R309 VTAIL.n48 VTAIL.n47 12.0247
R310 VTAIL.n91 VTAIL.n64 12.0247
R311 VTAIL.n102 VTAIL.n101 12.0247
R312 VTAIL.n147 VTAIL.n120 12.0247
R313 VTAIL.n158 VTAIL.n157 12.0247
R314 VTAIL.n378 VTAIL.n377 12.0247
R315 VTAIL.n368 VTAIL.n341 12.0247
R316 VTAIL.n322 VTAIL.n321 12.0247
R317 VTAIL.n312 VTAIL.n285 12.0247
R318 VTAIL.n268 VTAIL.n267 12.0247
R319 VTAIL.n258 VTAIL.n231 12.0247
R320 VTAIL.n212 VTAIL.n211 12.0247
R321 VTAIL.n202 VTAIL.n175 12.0247
R322 VTAIL.n418 VTAIL.n417 11.249
R323 VTAIL.n435 VTAIL.n388 11.249
R324 VTAIL.n34 VTAIL.n33 11.249
R325 VTAIL.n51 VTAIL.n4 11.249
R326 VTAIL.n88 VTAIL.n87 11.249
R327 VTAIL.n105 VTAIL.n58 11.249
R328 VTAIL.n144 VTAIL.n143 11.249
R329 VTAIL.n161 VTAIL.n114 11.249
R330 VTAIL.n381 VTAIL.n334 11.249
R331 VTAIL.n365 VTAIL.n364 11.249
R332 VTAIL.n325 VTAIL.n278 11.249
R333 VTAIL.n309 VTAIL.n308 11.249
R334 VTAIL.n271 VTAIL.n224 11.249
R335 VTAIL.n255 VTAIL.n254 11.249
R336 VTAIL.n215 VTAIL.n168 11.249
R337 VTAIL.n199 VTAIL.n198 11.249
R338 VTAIL.n414 VTAIL.n396 10.4732
R339 VTAIL.n436 VTAIL.n386 10.4732
R340 VTAIL.n30 VTAIL.n12 10.4732
R341 VTAIL.n52 VTAIL.n2 10.4732
R342 VTAIL.n84 VTAIL.n66 10.4732
R343 VTAIL.n106 VTAIL.n56 10.4732
R344 VTAIL.n140 VTAIL.n122 10.4732
R345 VTAIL.n162 VTAIL.n112 10.4732
R346 VTAIL.n382 VTAIL.n332 10.4732
R347 VTAIL.n361 VTAIL.n343 10.4732
R348 VTAIL.n326 VTAIL.n276 10.4732
R349 VTAIL.n305 VTAIL.n287 10.4732
R350 VTAIL.n272 VTAIL.n222 10.4732
R351 VTAIL.n251 VTAIL.n233 10.4732
R352 VTAIL.n216 VTAIL.n166 10.4732
R353 VTAIL.n195 VTAIL.n177 10.4732
R354 VTAIL.n403 VTAIL.n402 10.2747
R355 VTAIL.n19 VTAIL.n18 10.2747
R356 VTAIL.n73 VTAIL.n72 10.2747
R357 VTAIL.n129 VTAIL.n128 10.2747
R358 VTAIL.n350 VTAIL.n349 10.2747
R359 VTAIL.n294 VTAIL.n293 10.2747
R360 VTAIL.n240 VTAIL.n239 10.2747
R361 VTAIL.n184 VTAIL.n183 10.2747
R362 VTAIL.n413 VTAIL.n398 9.69747
R363 VTAIL.n29 VTAIL.n14 9.69747
R364 VTAIL.n83 VTAIL.n68 9.69747
R365 VTAIL.n139 VTAIL.n124 9.69747
R366 VTAIL.n360 VTAIL.n345 9.69747
R367 VTAIL.n304 VTAIL.n289 9.69747
R368 VTAIL.n250 VTAIL.n235 9.69747
R369 VTAIL.n194 VTAIL.n179 9.69747
R370 VTAIL.n438 VTAIL.n437 9.45567
R371 VTAIL.n54 VTAIL.n53 9.45567
R372 VTAIL.n108 VTAIL.n107 9.45567
R373 VTAIL.n164 VTAIL.n163 9.45567
R374 VTAIL.n384 VTAIL.n383 9.45567
R375 VTAIL.n328 VTAIL.n327 9.45567
R376 VTAIL.n274 VTAIL.n273 9.45567
R377 VTAIL.n218 VTAIL.n217 9.45567
R378 VTAIL.n437 VTAIL.n436 9.3005
R379 VTAIL.n388 VTAIL.n387 9.3005
R380 VTAIL.n431 VTAIL.n430 9.3005
R381 VTAIL.n429 VTAIL.n428 9.3005
R382 VTAIL.n405 VTAIL.n404 9.3005
R383 VTAIL.n400 VTAIL.n399 9.3005
R384 VTAIL.n411 VTAIL.n410 9.3005
R385 VTAIL.n413 VTAIL.n412 9.3005
R386 VTAIL.n396 VTAIL.n395 9.3005
R387 VTAIL.n419 VTAIL.n418 9.3005
R388 VTAIL.n421 VTAIL.n420 9.3005
R389 VTAIL.n422 VTAIL.n391 9.3005
R390 VTAIL.n53 VTAIL.n52 9.3005
R391 VTAIL.n4 VTAIL.n3 9.3005
R392 VTAIL.n47 VTAIL.n46 9.3005
R393 VTAIL.n45 VTAIL.n44 9.3005
R394 VTAIL.n21 VTAIL.n20 9.3005
R395 VTAIL.n16 VTAIL.n15 9.3005
R396 VTAIL.n27 VTAIL.n26 9.3005
R397 VTAIL.n29 VTAIL.n28 9.3005
R398 VTAIL.n12 VTAIL.n11 9.3005
R399 VTAIL.n35 VTAIL.n34 9.3005
R400 VTAIL.n37 VTAIL.n36 9.3005
R401 VTAIL.n38 VTAIL.n7 9.3005
R402 VTAIL.n107 VTAIL.n106 9.3005
R403 VTAIL.n58 VTAIL.n57 9.3005
R404 VTAIL.n101 VTAIL.n100 9.3005
R405 VTAIL.n99 VTAIL.n98 9.3005
R406 VTAIL.n75 VTAIL.n74 9.3005
R407 VTAIL.n70 VTAIL.n69 9.3005
R408 VTAIL.n81 VTAIL.n80 9.3005
R409 VTAIL.n83 VTAIL.n82 9.3005
R410 VTAIL.n66 VTAIL.n65 9.3005
R411 VTAIL.n89 VTAIL.n88 9.3005
R412 VTAIL.n91 VTAIL.n90 9.3005
R413 VTAIL.n92 VTAIL.n61 9.3005
R414 VTAIL.n163 VTAIL.n162 9.3005
R415 VTAIL.n114 VTAIL.n113 9.3005
R416 VTAIL.n157 VTAIL.n156 9.3005
R417 VTAIL.n155 VTAIL.n154 9.3005
R418 VTAIL.n131 VTAIL.n130 9.3005
R419 VTAIL.n126 VTAIL.n125 9.3005
R420 VTAIL.n137 VTAIL.n136 9.3005
R421 VTAIL.n139 VTAIL.n138 9.3005
R422 VTAIL.n122 VTAIL.n121 9.3005
R423 VTAIL.n145 VTAIL.n144 9.3005
R424 VTAIL.n147 VTAIL.n146 9.3005
R425 VTAIL.n148 VTAIL.n117 9.3005
R426 VTAIL.n352 VTAIL.n351 9.3005
R427 VTAIL.n347 VTAIL.n346 9.3005
R428 VTAIL.n358 VTAIL.n357 9.3005
R429 VTAIL.n360 VTAIL.n359 9.3005
R430 VTAIL.n343 VTAIL.n342 9.3005
R431 VTAIL.n366 VTAIL.n365 9.3005
R432 VTAIL.n368 VTAIL.n367 9.3005
R433 VTAIL.n340 VTAIL.n337 9.3005
R434 VTAIL.n383 VTAIL.n382 9.3005
R435 VTAIL.n334 VTAIL.n333 9.3005
R436 VTAIL.n377 VTAIL.n376 9.3005
R437 VTAIL.n375 VTAIL.n374 9.3005
R438 VTAIL.n296 VTAIL.n295 9.3005
R439 VTAIL.n291 VTAIL.n290 9.3005
R440 VTAIL.n302 VTAIL.n301 9.3005
R441 VTAIL.n304 VTAIL.n303 9.3005
R442 VTAIL.n287 VTAIL.n286 9.3005
R443 VTAIL.n310 VTAIL.n309 9.3005
R444 VTAIL.n312 VTAIL.n311 9.3005
R445 VTAIL.n284 VTAIL.n281 9.3005
R446 VTAIL.n327 VTAIL.n326 9.3005
R447 VTAIL.n278 VTAIL.n277 9.3005
R448 VTAIL.n321 VTAIL.n320 9.3005
R449 VTAIL.n319 VTAIL.n318 9.3005
R450 VTAIL.n242 VTAIL.n241 9.3005
R451 VTAIL.n237 VTAIL.n236 9.3005
R452 VTAIL.n248 VTAIL.n247 9.3005
R453 VTAIL.n250 VTAIL.n249 9.3005
R454 VTAIL.n233 VTAIL.n232 9.3005
R455 VTAIL.n256 VTAIL.n255 9.3005
R456 VTAIL.n258 VTAIL.n257 9.3005
R457 VTAIL.n230 VTAIL.n227 9.3005
R458 VTAIL.n273 VTAIL.n272 9.3005
R459 VTAIL.n224 VTAIL.n223 9.3005
R460 VTAIL.n267 VTAIL.n266 9.3005
R461 VTAIL.n265 VTAIL.n264 9.3005
R462 VTAIL.n186 VTAIL.n185 9.3005
R463 VTAIL.n181 VTAIL.n180 9.3005
R464 VTAIL.n192 VTAIL.n191 9.3005
R465 VTAIL.n194 VTAIL.n193 9.3005
R466 VTAIL.n177 VTAIL.n176 9.3005
R467 VTAIL.n200 VTAIL.n199 9.3005
R468 VTAIL.n202 VTAIL.n201 9.3005
R469 VTAIL.n174 VTAIL.n171 9.3005
R470 VTAIL.n217 VTAIL.n216 9.3005
R471 VTAIL.n168 VTAIL.n167 9.3005
R472 VTAIL.n211 VTAIL.n210 9.3005
R473 VTAIL.n209 VTAIL.n208 9.3005
R474 VTAIL.n410 VTAIL.n409 8.92171
R475 VTAIL.n26 VTAIL.n25 8.92171
R476 VTAIL.n80 VTAIL.n79 8.92171
R477 VTAIL.n136 VTAIL.n135 8.92171
R478 VTAIL.n357 VTAIL.n356 8.92171
R479 VTAIL.n301 VTAIL.n300 8.92171
R480 VTAIL.n247 VTAIL.n246 8.92171
R481 VTAIL.n191 VTAIL.n190 8.92171
R482 VTAIL.n406 VTAIL.n400 8.14595
R483 VTAIL.n22 VTAIL.n16 8.14595
R484 VTAIL.n76 VTAIL.n70 8.14595
R485 VTAIL.n132 VTAIL.n126 8.14595
R486 VTAIL.n353 VTAIL.n347 8.14595
R487 VTAIL.n297 VTAIL.n291 8.14595
R488 VTAIL.n243 VTAIL.n237 8.14595
R489 VTAIL.n187 VTAIL.n181 8.14595
R490 VTAIL.n405 VTAIL.n402 7.3702
R491 VTAIL.n21 VTAIL.n18 7.3702
R492 VTAIL.n75 VTAIL.n72 7.3702
R493 VTAIL.n131 VTAIL.n128 7.3702
R494 VTAIL.n352 VTAIL.n349 7.3702
R495 VTAIL.n296 VTAIL.n293 7.3702
R496 VTAIL.n242 VTAIL.n239 7.3702
R497 VTAIL.n186 VTAIL.n183 7.3702
R498 VTAIL.n406 VTAIL.n405 5.81868
R499 VTAIL.n22 VTAIL.n21 5.81868
R500 VTAIL.n76 VTAIL.n75 5.81868
R501 VTAIL.n132 VTAIL.n131 5.81868
R502 VTAIL.n353 VTAIL.n352 5.81868
R503 VTAIL.n297 VTAIL.n296 5.81868
R504 VTAIL.n243 VTAIL.n242 5.81868
R505 VTAIL.n187 VTAIL.n186 5.81868
R506 VTAIL.n409 VTAIL.n400 5.04292
R507 VTAIL.n25 VTAIL.n16 5.04292
R508 VTAIL.n79 VTAIL.n70 5.04292
R509 VTAIL.n135 VTAIL.n126 5.04292
R510 VTAIL.n356 VTAIL.n347 5.04292
R511 VTAIL.n300 VTAIL.n291 5.04292
R512 VTAIL.n246 VTAIL.n237 5.04292
R513 VTAIL.n190 VTAIL.n181 5.04292
R514 VTAIL.n410 VTAIL.n398 4.26717
R515 VTAIL.n26 VTAIL.n14 4.26717
R516 VTAIL.n80 VTAIL.n68 4.26717
R517 VTAIL.n136 VTAIL.n124 4.26717
R518 VTAIL.n357 VTAIL.n345 4.26717
R519 VTAIL.n301 VTAIL.n289 4.26717
R520 VTAIL.n247 VTAIL.n235 4.26717
R521 VTAIL.n191 VTAIL.n179 4.26717
R522 VTAIL.n414 VTAIL.n413 3.49141
R523 VTAIL.n438 VTAIL.n386 3.49141
R524 VTAIL.n30 VTAIL.n29 3.49141
R525 VTAIL.n54 VTAIL.n2 3.49141
R526 VTAIL.n84 VTAIL.n83 3.49141
R527 VTAIL.n108 VTAIL.n56 3.49141
R528 VTAIL.n140 VTAIL.n139 3.49141
R529 VTAIL.n164 VTAIL.n112 3.49141
R530 VTAIL.n384 VTAIL.n332 3.49141
R531 VTAIL.n361 VTAIL.n360 3.49141
R532 VTAIL.n328 VTAIL.n276 3.49141
R533 VTAIL.n305 VTAIL.n304 3.49141
R534 VTAIL.n274 VTAIL.n222 3.49141
R535 VTAIL.n251 VTAIL.n250 3.49141
R536 VTAIL.n218 VTAIL.n166 3.49141
R537 VTAIL.n195 VTAIL.n194 3.49141
R538 VTAIL.n404 VTAIL.n403 2.84303
R539 VTAIL.n20 VTAIL.n19 2.84303
R540 VTAIL.n74 VTAIL.n73 2.84303
R541 VTAIL.n130 VTAIL.n129 2.84303
R542 VTAIL.n351 VTAIL.n350 2.84303
R543 VTAIL.n295 VTAIL.n294 2.84303
R544 VTAIL.n241 VTAIL.n240 2.84303
R545 VTAIL.n185 VTAIL.n184 2.84303
R546 VTAIL.n417 VTAIL.n396 2.71565
R547 VTAIL.n436 VTAIL.n435 2.71565
R548 VTAIL.n33 VTAIL.n12 2.71565
R549 VTAIL.n52 VTAIL.n51 2.71565
R550 VTAIL.n87 VTAIL.n66 2.71565
R551 VTAIL.n106 VTAIL.n105 2.71565
R552 VTAIL.n143 VTAIL.n122 2.71565
R553 VTAIL.n162 VTAIL.n161 2.71565
R554 VTAIL.n382 VTAIL.n381 2.71565
R555 VTAIL.n364 VTAIL.n343 2.71565
R556 VTAIL.n326 VTAIL.n325 2.71565
R557 VTAIL.n308 VTAIL.n287 2.71565
R558 VTAIL.n272 VTAIL.n271 2.71565
R559 VTAIL.n254 VTAIL.n233 2.71565
R560 VTAIL.n216 VTAIL.n215 2.71565
R561 VTAIL.n198 VTAIL.n177 2.71565
R562 VTAIL.n0 VTAIL.t8 2.00455
R563 VTAIL.n0 VTAIL.t9 2.00455
R564 VTAIL.n110 VTAIL.t14 2.00455
R565 VTAIL.n110 VTAIL.t0 2.00455
R566 VTAIL.n330 VTAIL.t5 2.00455
R567 VTAIL.n330 VTAIL.t3 2.00455
R568 VTAIL.n220 VTAIL.t7 2.00455
R569 VTAIL.n220 VTAIL.t12 2.00455
R570 VTAIL.n418 VTAIL.n394 1.93989
R571 VTAIL.n432 VTAIL.n388 1.93989
R572 VTAIL.n34 VTAIL.n10 1.93989
R573 VTAIL.n48 VTAIL.n4 1.93989
R574 VTAIL.n88 VTAIL.n64 1.93989
R575 VTAIL.n102 VTAIL.n58 1.93989
R576 VTAIL.n144 VTAIL.n120 1.93989
R577 VTAIL.n158 VTAIL.n114 1.93989
R578 VTAIL.n378 VTAIL.n334 1.93989
R579 VTAIL.n365 VTAIL.n341 1.93989
R580 VTAIL.n322 VTAIL.n278 1.93989
R581 VTAIL.n309 VTAIL.n285 1.93989
R582 VTAIL.n268 VTAIL.n224 1.93989
R583 VTAIL.n255 VTAIL.n231 1.93989
R584 VTAIL.n212 VTAIL.n168 1.93989
R585 VTAIL.n199 VTAIL.n175 1.93989
R586 VTAIL.n423 VTAIL.n421 1.16414
R587 VTAIL.n431 VTAIL.n390 1.16414
R588 VTAIL.n39 VTAIL.n37 1.16414
R589 VTAIL.n47 VTAIL.n6 1.16414
R590 VTAIL.n93 VTAIL.n91 1.16414
R591 VTAIL.n101 VTAIL.n60 1.16414
R592 VTAIL.n149 VTAIL.n147 1.16414
R593 VTAIL.n157 VTAIL.n116 1.16414
R594 VTAIL.n377 VTAIL.n336 1.16414
R595 VTAIL.n369 VTAIL.n368 1.16414
R596 VTAIL.n321 VTAIL.n280 1.16414
R597 VTAIL.n313 VTAIL.n312 1.16414
R598 VTAIL.n267 VTAIL.n226 1.16414
R599 VTAIL.n259 VTAIL.n258 1.16414
R600 VTAIL.n211 VTAIL.n170 1.16414
R601 VTAIL.n203 VTAIL.n202 1.16414
R602 VTAIL.n221 VTAIL.n219 0.698776
R603 VTAIL.n275 VTAIL.n221 0.698776
R604 VTAIL.n331 VTAIL.n329 0.698776
R605 VTAIL.n385 VTAIL.n331 0.698776
R606 VTAIL.n165 VTAIL.n111 0.698776
R607 VTAIL.n111 VTAIL.n109 0.698776
R608 VTAIL.n55 VTAIL.n1 0.698776
R609 VTAIL VTAIL.n439 0.640586
R610 VTAIL.n329 VTAIL.n275 0.470328
R611 VTAIL.n109 VTAIL.n55 0.470328
R612 VTAIL.n422 VTAIL.n392 0.388379
R613 VTAIL.n428 VTAIL.n427 0.388379
R614 VTAIL.n38 VTAIL.n8 0.388379
R615 VTAIL.n44 VTAIL.n43 0.388379
R616 VTAIL.n92 VTAIL.n62 0.388379
R617 VTAIL.n98 VTAIL.n97 0.388379
R618 VTAIL.n148 VTAIL.n118 0.388379
R619 VTAIL.n154 VTAIL.n153 0.388379
R620 VTAIL.n374 VTAIL.n373 0.388379
R621 VTAIL.n340 VTAIL.n338 0.388379
R622 VTAIL.n318 VTAIL.n317 0.388379
R623 VTAIL.n284 VTAIL.n282 0.388379
R624 VTAIL.n264 VTAIL.n263 0.388379
R625 VTAIL.n230 VTAIL.n228 0.388379
R626 VTAIL.n208 VTAIL.n207 0.388379
R627 VTAIL.n174 VTAIL.n172 0.388379
R628 VTAIL.n404 VTAIL.n399 0.155672
R629 VTAIL.n411 VTAIL.n399 0.155672
R630 VTAIL.n412 VTAIL.n411 0.155672
R631 VTAIL.n412 VTAIL.n395 0.155672
R632 VTAIL.n419 VTAIL.n395 0.155672
R633 VTAIL.n420 VTAIL.n419 0.155672
R634 VTAIL.n420 VTAIL.n391 0.155672
R635 VTAIL.n429 VTAIL.n391 0.155672
R636 VTAIL.n430 VTAIL.n429 0.155672
R637 VTAIL.n430 VTAIL.n387 0.155672
R638 VTAIL.n437 VTAIL.n387 0.155672
R639 VTAIL.n20 VTAIL.n15 0.155672
R640 VTAIL.n27 VTAIL.n15 0.155672
R641 VTAIL.n28 VTAIL.n27 0.155672
R642 VTAIL.n28 VTAIL.n11 0.155672
R643 VTAIL.n35 VTAIL.n11 0.155672
R644 VTAIL.n36 VTAIL.n35 0.155672
R645 VTAIL.n36 VTAIL.n7 0.155672
R646 VTAIL.n45 VTAIL.n7 0.155672
R647 VTAIL.n46 VTAIL.n45 0.155672
R648 VTAIL.n46 VTAIL.n3 0.155672
R649 VTAIL.n53 VTAIL.n3 0.155672
R650 VTAIL.n74 VTAIL.n69 0.155672
R651 VTAIL.n81 VTAIL.n69 0.155672
R652 VTAIL.n82 VTAIL.n81 0.155672
R653 VTAIL.n82 VTAIL.n65 0.155672
R654 VTAIL.n89 VTAIL.n65 0.155672
R655 VTAIL.n90 VTAIL.n89 0.155672
R656 VTAIL.n90 VTAIL.n61 0.155672
R657 VTAIL.n99 VTAIL.n61 0.155672
R658 VTAIL.n100 VTAIL.n99 0.155672
R659 VTAIL.n100 VTAIL.n57 0.155672
R660 VTAIL.n107 VTAIL.n57 0.155672
R661 VTAIL.n130 VTAIL.n125 0.155672
R662 VTAIL.n137 VTAIL.n125 0.155672
R663 VTAIL.n138 VTAIL.n137 0.155672
R664 VTAIL.n138 VTAIL.n121 0.155672
R665 VTAIL.n145 VTAIL.n121 0.155672
R666 VTAIL.n146 VTAIL.n145 0.155672
R667 VTAIL.n146 VTAIL.n117 0.155672
R668 VTAIL.n155 VTAIL.n117 0.155672
R669 VTAIL.n156 VTAIL.n155 0.155672
R670 VTAIL.n156 VTAIL.n113 0.155672
R671 VTAIL.n163 VTAIL.n113 0.155672
R672 VTAIL.n383 VTAIL.n333 0.155672
R673 VTAIL.n376 VTAIL.n333 0.155672
R674 VTAIL.n376 VTAIL.n375 0.155672
R675 VTAIL.n375 VTAIL.n337 0.155672
R676 VTAIL.n367 VTAIL.n337 0.155672
R677 VTAIL.n367 VTAIL.n366 0.155672
R678 VTAIL.n366 VTAIL.n342 0.155672
R679 VTAIL.n359 VTAIL.n342 0.155672
R680 VTAIL.n359 VTAIL.n358 0.155672
R681 VTAIL.n358 VTAIL.n346 0.155672
R682 VTAIL.n351 VTAIL.n346 0.155672
R683 VTAIL.n327 VTAIL.n277 0.155672
R684 VTAIL.n320 VTAIL.n277 0.155672
R685 VTAIL.n320 VTAIL.n319 0.155672
R686 VTAIL.n319 VTAIL.n281 0.155672
R687 VTAIL.n311 VTAIL.n281 0.155672
R688 VTAIL.n311 VTAIL.n310 0.155672
R689 VTAIL.n310 VTAIL.n286 0.155672
R690 VTAIL.n303 VTAIL.n286 0.155672
R691 VTAIL.n303 VTAIL.n302 0.155672
R692 VTAIL.n302 VTAIL.n290 0.155672
R693 VTAIL.n295 VTAIL.n290 0.155672
R694 VTAIL.n273 VTAIL.n223 0.155672
R695 VTAIL.n266 VTAIL.n223 0.155672
R696 VTAIL.n266 VTAIL.n265 0.155672
R697 VTAIL.n265 VTAIL.n227 0.155672
R698 VTAIL.n257 VTAIL.n227 0.155672
R699 VTAIL.n257 VTAIL.n256 0.155672
R700 VTAIL.n256 VTAIL.n232 0.155672
R701 VTAIL.n249 VTAIL.n232 0.155672
R702 VTAIL.n249 VTAIL.n248 0.155672
R703 VTAIL.n248 VTAIL.n236 0.155672
R704 VTAIL.n241 VTAIL.n236 0.155672
R705 VTAIL.n217 VTAIL.n167 0.155672
R706 VTAIL.n210 VTAIL.n167 0.155672
R707 VTAIL.n210 VTAIL.n209 0.155672
R708 VTAIL.n209 VTAIL.n171 0.155672
R709 VTAIL.n201 VTAIL.n171 0.155672
R710 VTAIL.n201 VTAIL.n200 0.155672
R711 VTAIL.n200 VTAIL.n176 0.155672
R712 VTAIL.n193 VTAIL.n176 0.155672
R713 VTAIL.n193 VTAIL.n192 0.155672
R714 VTAIL.n192 VTAIL.n180 0.155672
R715 VTAIL.n185 VTAIL.n180 0.155672
R716 VTAIL VTAIL.n1 0.0586897
R717 B.n298 B.t10 702.968
R718 B.n307 B.t14 702.968
R719 B.n83 B.t6 702.968
R720 B.n81 B.t17 702.968
R721 B.n572 B.n571 585
R722 B.n241 B.n80 585
R723 B.n240 B.n239 585
R724 B.n238 B.n237 585
R725 B.n236 B.n235 585
R726 B.n234 B.n233 585
R727 B.n232 B.n231 585
R728 B.n230 B.n229 585
R729 B.n228 B.n227 585
R730 B.n226 B.n225 585
R731 B.n224 B.n223 585
R732 B.n222 B.n221 585
R733 B.n220 B.n219 585
R734 B.n218 B.n217 585
R735 B.n216 B.n215 585
R736 B.n214 B.n213 585
R737 B.n212 B.n211 585
R738 B.n210 B.n209 585
R739 B.n208 B.n207 585
R740 B.n206 B.n205 585
R741 B.n204 B.n203 585
R742 B.n202 B.n201 585
R743 B.n200 B.n199 585
R744 B.n198 B.n197 585
R745 B.n196 B.n195 585
R746 B.n194 B.n193 585
R747 B.n192 B.n191 585
R748 B.n190 B.n189 585
R749 B.n188 B.n187 585
R750 B.n186 B.n185 585
R751 B.n184 B.n183 585
R752 B.n182 B.n181 585
R753 B.n180 B.n179 585
R754 B.n178 B.n177 585
R755 B.n176 B.n175 585
R756 B.n173 B.n172 585
R757 B.n171 B.n170 585
R758 B.n169 B.n168 585
R759 B.n167 B.n166 585
R760 B.n165 B.n164 585
R761 B.n163 B.n162 585
R762 B.n161 B.n160 585
R763 B.n159 B.n158 585
R764 B.n157 B.n156 585
R765 B.n155 B.n154 585
R766 B.n152 B.n151 585
R767 B.n150 B.n149 585
R768 B.n148 B.n147 585
R769 B.n146 B.n145 585
R770 B.n144 B.n143 585
R771 B.n142 B.n141 585
R772 B.n140 B.n139 585
R773 B.n138 B.n137 585
R774 B.n136 B.n135 585
R775 B.n134 B.n133 585
R776 B.n132 B.n131 585
R777 B.n130 B.n129 585
R778 B.n128 B.n127 585
R779 B.n126 B.n125 585
R780 B.n124 B.n123 585
R781 B.n122 B.n121 585
R782 B.n120 B.n119 585
R783 B.n118 B.n117 585
R784 B.n116 B.n115 585
R785 B.n114 B.n113 585
R786 B.n112 B.n111 585
R787 B.n110 B.n109 585
R788 B.n108 B.n107 585
R789 B.n106 B.n105 585
R790 B.n104 B.n103 585
R791 B.n102 B.n101 585
R792 B.n100 B.n99 585
R793 B.n98 B.n97 585
R794 B.n96 B.n95 585
R795 B.n94 B.n93 585
R796 B.n92 B.n91 585
R797 B.n90 B.n89 585
R798 B.n88 B.n87 585
R799 B.n86 B.n85 585
R800 B.n39 B.n38 585
R801 B.n570 B.n40 585
R802 B.n575 B.n40 585
R803 B.n569 B.n568 585
R804 B.n568 B.n36 585
R805 B.n567 B.n35 585
R806 B.n581 B.n35 585
R807 B.n566 B.n34 585
R808 B.n582 B.n34 585
R809 B.n565 B.n33 585
R810 B.n583 B.n33 585
R811 B.n564 B.n563 585
R812 B.n563 B.n29 585
R813 B.n562 B.n28 585
R814 B.n589 B.n28 585
R815 B.n561 B.n27 585
R816 B.n590 B.n27 585
R817 B.n560 B.n26 585
R818 B.n591 B.n26 585
R819 B.n559 B.n558 585
R820 B.n558 B.n22 585
R821 B.n557 B.n21 585
R822 B.n597 B.n21 585
R823 B.n556 B.n20 585
R824 B.n598 B.n20 585
R825 B.n555 B.n19 585
R826 B.n599 B.n19 585
R827 B.n554 B.n553 585
R828 B.n553 B.n15 585
R829 B.n552 B.n14 585
R830 B.n605 B.n14 585
R831 B.n551 B.n13 585
R832 B.n606 B.n13 585
R833 B.n550 B.n12 585
R834 B.n607 B.n12 585
R835 B.n549 B.n548 585
R836 B.n548 B.n11 585
R837 B.n547 B.n7 585
R838 B.n613 B.n7 585
R839 B.n546 B.n6 585
R840 B.n614 B.n6 585
R841 B.n545 B.n5 585
R842 B.n615 B.n5 585
R843 B.n544 B.n543 585
R844 B.n543 B.n4 585
R845 B.n542 B.n242 585
R846 B.n542 B.n541 585
R847 B.n531 B.n243 585
R848 B.n534 B.n243 585
R849 B.n533 B.n532 585
R850 B.n535 B.n533 585
R851 B.n530 B.n248 585
R852 B.n248 B.n247 585
R853 B.n529 B.n528 585
R854 B.n528 B.n527 585
R855 B.n250 B.n249 585
R856 B.n251 B.n250 585
R857 B.n520 B.n519 585
R858 B.n521 B.n520 585
R859 B.n518 B.n256 585
R860 B.n256 B.n255 585
R861 B.n517 B.n516 585
R862 B.n516 B.n515 585
R863 B.n258 B.n257 585
R864 B.n259 B.n258 585
R865 B.n508 B.n507 585
R866 B.n509 B.n508 585
R867 B.n506 B.n264 585
R868 B.n264 B.n263 585
R869 B.n505 B.n504 585
R870 B.n504 B.n503 585
R871 B.n266 B.n265 585
R872 B.n267 B.n266 585
R873 B.n496 B.n495 585
R874 B.n497 B.n496 585
R875 B.n494 B.n272 585
R876 B.n272 B.n271 585
R877 B.n493 B.n492 585
R878 B.n492 B.n491 585
R879 B.n274 B.n273 585
R880 B.n275 B.n274 585
R881 B.n484 B.n483 585
R882 B.n485 B.n484 585
R883 B.n278 B.n277 585
R884 B.n327 B.n326 585
R885 B.n328 B.n324 585
R886 B.n324 B.n279 585
R887 B.n330 B.n329 585
R888 B.n332 B.n323 585
R889 B.n335 B.n334 585
R890 B.n336 B.n322 585
R891 B.n338 B.n337 585
R892 B.n340 B.n321 585
R893 B.n343 B.n342 585
R894 B.n344 B.n320 585
R895 B.n346 B.n345 585
R896 B.n348 B.n319 585
R897 B.n351 B.n350 585
R898 B.n352 B.n318 585
R899 B.n354 B.n353 585
R900 B.n356 B.n317 585
R901 B.n359 B.n358 585
R902 B.n360 B.n316 585
R903 B.n362 B.n361 585
R904 B.n364 B.n315 585
R905 B.n367 B.n366 585
R906 B.n368 B.n314 585
R907 B.n370 B.n369 585
R908 B.n372 B.n313 585
R909 B.n375 B.n374 585
R910 B.n376 B.n312 585
R911 B.n378 B.n377 585
R912 B.n380 B.n311 585
R913 B.n383 B.n382 585
R914 B.n384 B.n310 585
R915 B.n386 B.n385 585
R916 B.n388 B.n309 585
R917 B.n391 B.n390 585
R918 B.n392 B.n306 585
R919 B.n395 B.n394 585
R920 B.n397 B.n305 585
R921 B.n400 B.n399 585
R922 B.n401 B.n304 585
R923 B.n403 B.n402 585
R924 B.n405 B.n303 585
R925 B.n408 B.n407 585
R926 B.n409 B.n302 585
R927 B.n411 B.n410 585
R928 B.n413 B.n301 585
R929 B.n416 B.n415 585
R930 B.n417 B.n297 585
R931 B.n419 B.n418 585
R932 B.n421 B.n296 585
R933 B.n424 B.n423 585
R934 B.n425 B.n295 585
R935 B.n427 B.n426 585
R936 B.n429 B.n294 585
R937 B.n432 B.n431 585
R938 B.n433 B.n293 585
R939 B.n435 B.n434 585
R940 B.n437 B.n292 585
R941 B.n440 B.n439 585
R942 B.n441 B.n291 585
R943 B.n443 B.n442 585
R944 B.n445 B.n290 585
R945 B.n448 B.n447 585
R946 B.n449 B.n289 585
R947 B.n451 B.n450 585
R948 B.n453 B.n288 585
R949 B.n456 B.n455 585
R950 B.n457 B.n287 585
R951 B.n459 B.n458 585
R952 B.n461 B.n286 585
R953 B.n464 B.n463 585
R954 B.n465 B.n285 585
R955 B.n467 B.n466 585
R956 B.n469 B.n284 585
R957 B.n472 B.n471 585
R958 B.n473 B.n283 585
R959 B.n475 B.n474 585
R960 B.n477 B.n282 585
R961 B.n478 B.n281 585
R962 B.n481 B.n480 585
R963 B.n482 B.n280 585
R964 B.n280 B.n279 585
R965 B.n487 B.n486 585
R966 B.n486 B.n485 585
R967 B.n488 B.n276 585
R968 B.n276 B.n275 585
R969 B.n490 B.n489 585
R970 B.n491 B.n490 585
R971 B.n270 B.n269 585
R972 B.n271 B.n270 585
R973 B.n499 B.n498 585
R974 B.n498 B.n497 585
R975 B.n500 B.n268 585
R976 B.n268 B.n267 585
R977 B.n502 B.n501 585
R978 B.n503 B.n502 585
R979 B.n262 B.n261 585
R980 B.n263 B.n262 585
R981 B.n511 B.n510 585
R982 B.n510 B.n509 585
R983 B.n512 B.n260 585
R984 B.n260 B.n259 585
R985 B.n514 B.n513 585
R986 B.n515 B.n514 585
R987 B.n254 B.n253 585
R988 B.n255 B.n254 585
R989 B.n523 B.n522 585
R990 B.n522 B.n521 585
R991 B.n524 B.n252 585
R992 B.n252 B.n251 585
R993 B.n526 B.n525 585
R994 B.n527 B.n526 585
R995 B.n246 B.n245 585
R996 B.n247 B.n246 585
R997 B.n537 B.n536 585
R998 B.n536 B.n535 585
R999 B.n538 B.n244 585
R1000 B.n534 B.n244 585
R1001 B.n540 B.n539 585
R1002 B.n541 B.n540 585
R1003 B.n2 B.n0 585
R1004 B.n4 B.n2 585
R1005 B.n3 B.n1 585
R1006 B.n614 B.n3 585
R1007 B.n612 B.n611 585
R1008 B.n613 B.n612 585
R1009 B.n610 B.n8 585
R1010 B.n11 B.n8 585
R1011 B.n609 B.n608 585
R1012 B.n608 B.n607 585
R1013 B.n10 B.n9 585
R1014 B.n606 B.n10 585
R1015 B.n604 B.n603 585
R1016 B.n605 B.n604 585
R1017 B.n602 B.n16 585
R1018 B.n16 B.n15 585
R1019 B.n601 B.n600 585
R1020 B.n600 B.n599 585
R1021 B.n18 B.n17 585
R1022 B.n598 B.n18 585
R1023 B.n596 B.n595 585
R1024 B.n597 B.n596 585
R1025 B.n594 B.n23 585
R1026 B.n23 B.n22 585
R1027 B.n593 B.n592 585
R1028 B.n592 B.n591 585
R1029 B.n25 B.n24 585
R1030 B.n590 B.n25 585
R1031 B.n588 B.n587 585
R1032 B.n589 B.n588 585
R1033 B.n586 B.n30 585
R1034 B.n30 B.n29 585
R1035 B.n585 B.n584 585
R1036 B.n584 B.n583 585
R1037 B.n32 B.n31 585
R1038 B.n582 B.n32 585
R1039 B.n580 B.n579 585
R1040 B.n581 B.n580 585
R1041 B.n578 B.n37 585
R1042 B.n37 B.n36 585
R1043 B.n577 B.n576 585
R1044 B.n576 B.n575 585
R1045 B.n617 B.n616 585
R1046 B.n616 B.n615 585
R1047 B.n486 B.n278 530.939
R1048 B.n576 B.n39 530.939
R1049 B.n484 B.n280 530.939
R1050 B.n572 B.n40 530.939
R1051 B.n298 B.t13 261.029
R1052 B.n81 B.t18 261.029
R1053 B.n307 B.t16 261.029
R1054 B.n83 B.t8 261.029
R1055 B.n574 B.n573 256.663
R1056 B.n574 B.n79 256.663
R1057 B.n574 B.n78 256.663
R1058 B.n574 B.n77 256.663
R1059 B.n574 B.n76 256.663
R1060 B.n574 B.n75 256.663
R1061 B.n574 B.n74 256.663
R1062 B.n574 B.n73 256.663
R1063 B.n574 B.n72 256.663
R1064 B.n574 B.n71 256.663
R1065 B.n574 B.n70 256.663
R1066 B.n574 B.n69 256.663
R1067 B.n574 B.n68 256.663
R1068 B.n574 B.n67 256.663
R1069 B.n574 B.n66 256.663
R1070 B.n574 B.n65 256.663
R1071 B.n574 B.n64 256.663
R1072 B.n574 B.n63 256.663
R1073 B.n574 B.n62 256.663
R1074 B.n574 B.n61 256.663
R1075 B.n574 B.n60 256.663
R1076 B.n574 B.n59 256.663
R1077 B.n574 B.n58 256.663
R1078 B.n574 B.n57 256.663
R1079 B.n574 B.n56 256.663
R1080 B.n574 B.n55 256.663
R1081 B.n574 B.n54 256.663
R1082 B.n574 B.n53 256.663
R1083 B.n574 B.n52 256.663
R1084 B.n574 B.n51 256.663
R1085 B.n574 B.n50 256.663
R1086 B.n574 B.n49 256.663
R1087 B.n574 B.n48 256.663
R1088 B.n574 B.n47 256.663
R1089 B.n574 B.n46 256.663
R1090 B.n574 B.n45 256.663
R1091 B.n574 B.n44 256.663
R1092 B.n574 B.n43 256.663
R1093 B.n574 B.n42 256.663
R1094 B.n574 B.n41 256.663
R1095 B.n325 B.n279 256.663
R1096 B.n331 B.n279 256.663
R1097 B.n333 B.n279 256.663
R1098 B.n339 B.n279 256.663
R1099 B.n341 B.n279 256.663
R1100 B.n347 B.n279 256.663
R1101 B.n349 B.n279 256.663
R1102 B.n355 B.n279 256.663
R1103 B.n357 B.n279 256.663
R1104 B.n363 B.n279 256.663
R1105 B.n365 B.n279 256.663
R1106 B.n371 B.n279 256.663
R1107 B.n373 B.n279 256.663
R1108 B.n379 B.n279 256.663
R1109 B.n381 B.n279 256.663
R1110 B.n387 B.n279 256.663
R1111 B.n389 B.n279 256.663
R1112 B.n396 B.n279 256.663
R1113 B.n398 B.n279 256.663
R1114 B.n404 B.n279 256.663
R1115 B.n406 B.n279 256.663
R1116 B.n412 B.n279 256.663
R1117 B.n414 B.n279 256.663
R1118 B.n420 B.n279 256.663
R1119 B.n422 B.n279 256.663
R1120 B.n428 B.n279 256.663
R1121 B.n430 B.n279 256.663
R1122 B.n436 B.n279 256.663
R1123 B.n438 B.n279 256.663
R1124 B.n444 B.n279 256.663
R1125 B.n446 B.n279 256.663
R1126 B.n452 B.n279 256.663
R1127 B.n454 B.n279 256.663
R1128 B.n460 B.n279 256.663
R1129 B.n462 B.n279 256.663
R1130 B.n468 B.n279 256.663
R1131 B.n470 B.n279 256.663
R1132 B.n476 B.n279 256.663
R1133 B.n479 B.n279 256.663
R1134 B.n299 B.t12 245.32
R1135 B.n82 B.t19 245.32
R1136 B.n308 B.t15 245.32
R1137 B.n84 B.t9 245.32
R1138 B.n486 B.n276 163.367
R1139 B.n490 B.n276 163.367
R1140 B.n490 B.n270 163.367
R1141 B.n498 B.n270 163.367
R1142 B.n498 B.n268 163.367
R1143 B.n502 B.n268 163.367
R1144 B.n502 B.n262 163.367
R1145 B.n510 B.n262 163.367
R1146 B.n510 B.n260 163.367
R1147 B.n514 B.n260 163.367
R1148 B.n514 B.n254 163.367
R1149 B.n522 B.n254 163.367
R1150 B.n522 B.n252 163.367
R1151 B.n526 B.n252 163.367
R1152 B.n526 B.n246 163.367
R1153 B.n536 B.n246 163.367
R1154 B.n536 B.n244 163.367
R1155 B.n540 B.n244 163.367
R1156 B.n540 B.n2 163.367
R1157 B.n616 B.n2 163.367
R1158 B.n616 B.n3 163.367
R1159 B.n612 B.n3 163.367
R1160 B.n612 B.n8 163.367
R1161 B.n608 B.n8 163.367
R1162 B.n608 B.n10 163.367
R1163 B.n604 B.n10 163.367
R1164 B.n604 B.n16 163.367
R1165 B.n600 B.n16 163.367
R1166 B.n600 B.n18 163.367
R1167 B.n596 B.n18 163.367
R1168 B.n596 B.n23 163.367
R1169 B.n592 B.n23 163.367
R1170 B.n592 B.n25 163.367
R1171 B.n588 B.n25 163.367
R1172 B.n588 B.n30 163.367
R1173 B.n584 B.n30 163.367
R1174 B.n584 B.n32 163.367
R1175 B.n580 B.n32 163.367
R1176 B.n580 B.n37 163.367
R1177 B.n576 B.n37 163.367
R1178 B.n326 B.n324 163.367
R1179 B.n330 B.n324 163.367
R1180 B.n334 B.n332 163.367
R1181 B.n338 B.n322 163.367
R1182 B.n342 B.n340 163.367
R1183 B.n346 B.n320 163.367
R1184 B.n350 B.n348 163.367
R1185 B.n354 B.n318 163.367
R1186 B.n358 B.n356 163.367
R1187 B.n362 B.n316 163.367
R1188 B.n366 B.n364 163.367
R1189 B.n370 B.n314 163.367
R1190 B.n374 B.n372 163.367
R1191 B.n378 B.n312 163.367
R1192 B.n382 B.n380 163.367
R1193 B.n386 B.n310 163.367
R1194 B.n390 B.n388 163.367
R1195 B.n395 B.n306 163.367
R1196 B.n399 B.n397 163.367
R1197 B.n403 B.n304 163.367
R1198 B.n407 B.n405 163.367
R1199 B.n411 B.n302 163.367
R1200 B.n415 B.n413 163.367
R1201 B.n419 B.n297 163.367
R1202 B.n423 B.n421 163.367
R1203 B.n427 B.n295 163.367
R1204 B.n431 B.n429 163.367
R1205 B.n435 B.n293 163.367
R1206 B.n439 B.n437 163.367
R1207 B.n443 B.n291 163.367
R1208 B.n447 B.n445 163.367
R1209 B.n451 B.n289 163.367
R1210 B.n455 B.n453 163.367
R1211 B.n459 B.n287 163.367
R1212 B.n463 B.n461 163.367
R1213 B.n467 B.n285 163.367
R1214 B.n471 B.n469 163.367
R1215 B.n475 B.n283 163.367
R1216 B.n478 B.n477 163.367
R1217 B.n480 B.n280 163.367
R1218 B.n484 B.n274 163.367
R1219 B.n492 B.n274 163.367
R1220 B.n492 B.n272 163.367
R1221 B.n496 B.n272 163.367
R1222 B.n496 B.n266 163.367
R1223 B.n504 B.n266 163.367
R1224 B.n504 B.n264 163.367
R1225 B.n508 B.n264 163.367
R1226 B.n508 B.n258 163.367
R1227 B.n516 B.n258 163.367
R1228 B.n516 B.n256 163.367
R1229 B.n520 B.n256 163.367
R1230 B.n520 B.n250 163.367
R1231 B.n528 B.n250 163.367
R1232 B.n528 B.n248 163.367
R1233 B.n533 B.n248 163.367
R1234 B.n533 B.n243 163.367
R1235 B.n542 B.n243 163.367
R1236 B.n543 B.n542 163.367
R1237 B.n543 B.n5 163.367
R1238 B.n6 B.n5 163.367
R1239 B.n7 B.n6 163.367
R1240 B.n548 B.n7 163.367
R1241 B.n548 B.n12 163.367
R1242 B.n13 B.n12 163.367
R1243 B.n14 B.n13 163.367
R1244 B.n553 B.n14 163.367
R1245 B.n553 B.n19 163.367
R1246 B.n20 B.n19 163.367
R1247 B.n21 B.n20 163.367
R1248 B.n558 B.n21 163.367
R1249 B.n558 B.n26 163.367
R1250 B.n27 B.n26 163.367
R1251 B.n28 B.n27 163.367
R1252 B.n563 B.n28 163.367
R1253 B.n563 B.n33 163.367
R1254 B.n34 B.n33 163.367
R1255 B.n35 B.n34 163.367
R1256 B.n568 B.n35 163.367
R1257 B.n568 B.n40 163.367
R1258 B.n87 B.n86 163.367
R1259 B.n91 B.n90 163.367
R1260 B.n95 B.n94 163.367
R1261 B.n99 B.n98 163.367
R1262 B.n103 B.n102 163.367
R1263 B.n107 B.n106 163.367
R1264 B.n111 B.n110 163.367
R1265 B.n115 B.n114 163.367
R1266 B.n119 B.n118 163.367
R1267 B.n123 B.n122 163.367
R1268 B.n127 B.n126 163.367
R1269 B.n131 B.n130 163.367
R1270 B.n135 B.n134 163.367
R1271 B.n139 B.n138 163.367
R1272 B.n143 B.n142 163.367
R1273 B.n147 B.n146 163.367
R1274 B.n151 B.n150 163.367
R1275 B.n156 B.n155 163.367
R1276 B.n160 B.n159 163.367
R1277 B.n164 B.n163 163.367
R1278 B.n168 B.n167 163.367
R1279 B.n172 B.n171 163.367
R1280 B.n177 B.n176 163.367
R1281 B.n181 B.n180 163.367
R1282 B.n185 B.n184 163.367
R1283 B.n189 B.n188 163.367
R1284 B.n193 B.n192 163.367
R1285 B.n197 B.n196 163.367
R1286 B.n201 B.n200 163.367
R1287 B.n205 B.n204 163.367
R1288 B.n209 B.n208 163.367
R1289 B.n213 B.n212 163.367
R1290 B.n217 B.n216 163.367
R1291 B.n221 B.n220 163.367
R1292 B.n225 B.n224 163.367
R1293 B.n229 B.n228 163.367
R1294 B.n233 B.n232 163.367
R1295 B.n237 B.n236 163.367
R1296 B.n239 B.n80 163.367
R1297 B.n485 B.n279 90.7296
R1298 B.n575 B.n574 90.7296
R1299 B.n325 B.n278 71.676
R1300 B.n331 B.n330 71.676
R1301 B.n334 B.n333 71.676
R1302 B.n339 B.n338 71.676
R1303 B.n342 B.n341 71.676
R1304 B.n347 B.n346 71.676
R1305 B.n350 B.n349 71.676
R1306 B.n355 B.n354 71.676
R1307 B.n358 B.n357 71.676
R1308 B.n363 B.n362 71.676
R1309 B.n366 B.n365 71.676
R1310 B.n371 B.n370 71.676
R1311 B.n374 B.n373 71.676
R1312 B.n379 B.n378 71.676
R1313 B.n382 B.n381 71.676
R1314 B.n387 B.n386 71.676
R1315 B.n390 B.n389 71.676
R1316 B.n396 B.n395 71.676
R1317 B.n399 B.n398 71.676
R1318 B.n404 B.n403 71.676
R1319 B.n407 B.n406 71.676
R1320 B.n412 B.n411 71.676
R1321 B.n415 B.n414 71.676
R1322 B.n420 B.n419 71.676
R1323 B.n423 B.n422 71.676
R1324 B.n428 B.n427 71.676
R1325 B.n431 B.n430 71.676
R1326 B.n436 B.n435 71.676
R1327 B.n439 B.n438 71.676
R1328 B.n444 B.n443 71.676
R1329 B.n447 B.n446 71.676
R1330 B.n452 B.n451 71.676
R1331 B.n455 B.n454 71.676
R1332 B.n460 B.n459 71.676
R1333 B.n463 B.n462 71.676
R1334 B.n468 B.n467 71.676
R1335 B.n471 B.n470 71.676
R1336 B.n476 B.n475 71.676
R1337 B.n479 B.n478 71.676
R1338 B.n41 B.n39 71.676
R1339 B.n87 B.n42 71.676
R1340 B.n91 B.n43 71.676
R1341 B.n95 B.n44 71.676
R1342 B.n99 B.n45 71.676
R1343 B.n103 B.n46 71.676
R1344 B.n107 B.n47 71.676
R1345 B.n111 B.n48 71.676
R1346 B.n115 B.n49 71.676
R1347 B.n119 B.n50 71.676
R1348 B.n123 B.n51 71.676
R1349 B.n127 B.n52 71.676
R1350 B.n131 B.n53 71.676
R1351 B.n135 B.n54 71.676
R1352 B.n139 B.n55 71.676
R1353 B.n143 B.n56 71.676
R1354 B.n147 B.n57 71.676
R1355 B.n151 B.n58 71.676
R1356 B.n156 B.n59 71.676
R1357 B.n160 B.n60 71.676
R1358 B.n164 B.n61 71.676
R1359 B.n168 B.n62 71.676
R1360 B.n172 B.n63 71.676
R1361 B.n177 B.n64 71.676
R1362 B.n181 B.n65 71.676
R1363 B.n185 B.n66 71.676
R1364 B.n189 B.n67 71.676
R1365 B.n193 B.n68 71.676
R1366 B.n197 B.n69 71.676
R1367 B.n201 B.n70 71.676
R1368 B.n205 B.n71 71.676
R1369 B.n209 B.n72 71.676
R1370 B.n213 B.n73 71.676
R1371 B.n217 B.n74 71.676
R1372 B.n221 B.n75 71.676
R1373 B.n225 B.n76 71.676
R1374 B.n229 B.n77 71.676
R1375 B.n233 B.n78 71.676
R1376 B.n237 B.n79 71.676
R1377 B.n573 B.n80 71.676
R1378 B.n573 B.n572 71.676
R1379 B.n239 B.n79 71.676
R1380 B.n236 B.n78 71.676
R1381 B.n232 B.n77 71.676
R1382 B.n228 B.n76 71.676
R1383 B.n224 B.n75 71.676
R1384 B.n220 B.n74 71.676
R1385 B.n216 B.n73 71.676
R1386 B.n212 B.n72 71.676
R1387 B.n208 B.n71 71.676
R1388 B.n204 B.n70 71.676
R1389 B.n200 B.n69 71.676
R1390 B.n196 B.n68 71.676
R1391 B.n192 B.n67 71.676
R1392 B.n188 B.n66 71.676
R1393 B.n184 B.n65 71.676
R1394 B.n180 B.n64 71.676
R1395 B.n176 B.n63 71.676
R1396 B.n171 B.n62 71.676
R1397 B.n167 B.n61 71.676
R1398 B.n163 B.n60 71.676
R1399 B.n159 B.n59 71.676
R1400 B.n155 B.n58 71.676
R1401 B.n150 B.n57 71.676
R1402 B.n146 B.n56 71.676
R1403 B.n142 B.n55 71.676
R1404 B.n138 B.n54 71.676
R1405 B.n134 B.n53 71.676
R1406 B.n130 B.n52 71.676
R1407 B.n126 B.n51 71.676
R1408 B.n122 B.n50 71.676
R1409 B.n118 B.n49 71.676
R1410 B.n114 B.n48 71.676
R1411 B.n110 B.n47 71.676
R1412 B.n106 B.n46 71.676
R1413 B.n102 B.n45 71.676
R1414 B.n98 B.n44 71.676
R1415 B.n94 B.n43 71.676
R1416 B.n90 B.n42 71.676
R1417 B.n86 B.n41 71.676
R1418 B.n326 B.n325 71.676
R1419 B.n332 B.n331 71.676
R1420 B.n333 B.n322 71.676
R1421 B.n340 B.n339 71.676
R1422 B.n341 B.n320 71.676
R1423 B.n348 B.n347 71.676
R1424 B.n349 B.n318 71.676
R1425 B.n356 B.n355 71.676
R1426 B.n357 B.n316 71.676
R1427 B.n364 B.n363 71.676
R1428 B.n365 B.n314 71.676
R1429 B.n372 B.n371 71.676
R1430 B.n373 B.n312 71.676
R1431 B.n380 B.n379 71.676
R1432 B.n381 B.n310 71.676
R1433 B.n388 B.n387 71.676
R1434 B.n389 B.n306 71.676
R1435 B.n397 B.n396 71.676
R1436 B.n398 B.n304 71.676
R1437 B.n405 B.n404 71.676
R1438 B.n406 B.n302 71.676
R1439 B.n413 B.n412 71.676
R1440 B.n414 B.n297 71.676
R1441 B.n421 B.n420 71.676
R1442 B.n422 B.n295 71.676
R1443 B.n429 B.n428 71.676
R1444 B.n430 B.n293 71.676
R1445 B.n437 B.n436 71.676
R1446 B.n438 B.n291 71.676
R1447 B.n445 B.n444 71.676
R1448 B.n446 B.n289 71.676
R1449 B.n453 B.n452 71.676
R1450 B.n454 B.n287 71.676
R1451 B.n461 B.n460 71.676
R1452 B.n462 B.n285 71.676
R1453 B.n469 B.n468 71.676
R1454 B.n470 B.n283 71.676
R1455 B.n477 B.n476 71.676
R1456 B.n480 B.n479 71.676
R1457 B.n300 B.n299 59.5399
R1458 B.n393 B.n308 59.5399
R1459 B.n153 B.n84 59.5399
R1460 B.n174 B.n82 59.5399
R1461 B.n485 B.n275 49.3571
R1462 B.n491 B.n275 49.3571
R1463 B.n491 B.n271 49.3571
R1464 B.n497 B.n271 49.3571
R1465 B.n503 B.n267 49.3571
R1466 B.n503 B.n263 49.3571
R1467 B.n509 B.n263 49.3571
R1468 B.n509 B.n259 49.3571
R1469 B.n515 B.n259 49.3571
R1470 B.n521 B.n255 49.3571
R1471 B.n527 B.n251 49.3571
R1472 B.n535 B.n247 49.3571
R1473 B.n535 B.n534 49.3571
R1474 B.n541 B.n4 49.3571
R1475 B.n615 B.n4 49.3571
R1476 B.n615 B.n614 49.3571
R1477 B.n614 B.n613 49.3571
R1478 B.n607 B.n11 49.3571
R1479 B.n607 B.n606 49.3571
R1480 B.n605 B.n15 49.3571
R1481 B.n599 B.n598 49.3571
R1482 B.n597 B.n22 49.3571
R1483 B.n591 B.n22 49.3571
R1484 B.n591 B.n590 49.3571
R1485 B.n590 B.n589 49.3571
R1486 B.n589 B.n29 49.3571
R1487 B.n583 B.n582 49.3571
R1488 B.n582 B.n581 49.3571
R1489 B.n581 B.n36 49.3571
R1490 B.n575 B.n36 49.3571
R1491 B.t2 B.n255 46.4538
R1492 B.n598 B.t20 46.4538
R1493 B.n527 B.t0 40.6472
R1494 B.t5 B.n605 40.6472
R1495 B.n541 B.t1 39.1955
R1496 B.n613 B.t4 39.1955
R1497 B.n577 B.n38 34.4981
R1498 B.n571 B.n570 34.4981
R1499 B.n483 B.n482 34.4981
R1500 B.n487 B.n277 34.4981
R1501 B.t21 B.n251 27.5822
R1502 B.t3 B.n15 27.5822
R1503 B.t11 B.n267 26.1305
R1504 B.t7 B.n29 26.1305
R1505 B.n497 B.t11 23.2272
R1506 B.n583 B.t7 23.2272
R1507 B.n521 B.t21 21.7755
R1508 B.n599 B.t3 21.7755
R1509 B B.n617 18.0485
R1510 B.n299 B.n298 15.7096
R1511 B.n308 B.n307 15.7096
R1512 B.n84 B.n83 15.7096
R1513 B.n82 B.n81 15.7096
R1514 B.n85 B.n38 10.6151
R1515 B.n88 B.n85 10.6151
R1516 B.n89 B.n88 10.6151
R1517 B.n92 B.n89 10.6151
R1518 B.n93 B.n92 10.6151
R1519 B.n96 B.n93 10.6151
R1520 B.n97 B.n96 10.6151
R1521 B.n100 B.n97 10.6151
R1522 B.n101 B.n100 10.6151
R1523 B.n104 B.n101 10.6151
R1524 B.n105 B.n104 10.6151
R1525 B.n108 B.n105 10.6151
R1526 B.n109 B.n108 10.6151
R1527 B.n112 B.n109 10.6151
R1528 B.n113 B.n112 10.6151
R1529 B.n116 B.n113 10.6151
R1530 B.n117 B.n116 10.6151
R1531 B.n120 B.n117 10.6151
R1532 B.n121 B.n120 10.6151
R1533 B.n124 B.n121 10.6151
R1534 B.n125 B.n124 10.6151
R1535 B.n128 B.n125 10.6151
R1536 B.n129 B.n128 10.6151
R1537 B.n132 B.n129 10.6151
R1538 B.n133 B.n132 10.6151
R1539 B.n136 B.n133 10.6151
R1540 B.n137 B.n136 10.6151
R1541 B.n140 B.n137 10.6151
R1542 B.n141 B.n140 10.6151
R1543 B.n144 B.n141 10.6151
R1544 B.n145 B.n144 10.6151
R1545 B.n148 B.n145 10.6151
R1546 B.n149 B.n148 10.6151
R1547 B.n152 B.n149 10.6151
R1548 B.n157 B.n154 10.6151
R1549 B.n158 B.n157 10.6151
R1550 B.n161 B.n158 10.6151
R1551 B.n162 B.n161 10.6151
R1552 B.n165 B.n162 10.6151
R1553 B.n166 B.n165 10.6151
R1554 B.n169 B.n166 10.6151
R1555 B.n170 B.n169 10.6151
R1556 B.n173 B.n170 10.6151
R1557 B.n178 B.n175 10.6151
R1558 B.n179 B.n178 10.6151
R1559 B.n182 B.n179 10.6151
R1560 B.n183 B.n182 10.6151
R1561 B.n186 B.n183 10.6151
R1562 B.n187 B.n186 10.6151
R1563 B.n190 B.n187 10.6151
R1564 B.n191 B.n190 10.6151
R1565 B.n194 B.n191 10.6151
R1566 B.n195 B.n194 10.6151
R1567 B.n198 B.n195 10.6151
R1568 B.n199 B.n198 10.6151
R1569 B.n202 B.n199 10.6151
R1570 B.n203 B.n202 10.6151
R1571 B.n206 B.n203 10.6151
R1572 B.n207 B.n206 10.6151
R1573 B.n210 B.n207 10.6151
R1574 B.n211 B.n210 10.6151
R1575 B.n214 B.n211 10.6151
R1576 B.n215 B.n214 10.6151
R1577 B.n218 B.n215 10.6151
R1578 B.n219 B.n218 10.6151
R1579 B.n222 B.n219 10.6151
R1580 B.n223 B.n222 10.6151
R1581 B.n226 B.n223 10.6151
R1582 B.n227 B.n226 10.6151
R1583 B.n230 B.n227 10.6151
R1584 B.n231 B.n230 10.6151
R1585 B.n234 B.n231 10.6151
R1586 B.n235 B.n234 10.6151
R1587 B.n238 B.n235 10.6151
R1588 B.n240 B.n238 10.6151
R1589 B.n241 B.n240 10.6151
R1590 B.n571 B.n241 10.6151
R1591 B.n483 B.n273 10.6151
R1592 B.n493 B.n273 10.6151
R1593 B.n494 B.n493 10.6151
R1594 B.n495 B.n494 10.6151
R1595 B.n495 B.n265 10.6151
R1596 B.n505 B.n265 10.6151
R1597 B.n506 B.n505 10.6151
R1598 B.n507 B.n506 10.6151
R1599 B.n507 B.n257 10.6151
R1600 B.n517 B.n257 10.6151
R1601 B.n518 B.n517 10.6151
R1602 B.n519 B.n518 10.6151
R1603 B.n519 B.n249 10.6151
R1604 B.n529 B.n249 10.6151
R1605 B.n530 B.n529 10.6151
R1606 B.n532 B.n530 10.6151
R1607 B.n532 B.n531 10.6151
R1608 B.n531 B.n242 10.6151
R1609 B.n544 B.n242 10.6151
R1610 B.n545 B.n544 10.6151
R1611 B.n546 B.n545 10.6151
R1612 B.n547 B.n546 10.6151
R1613 B.n549 B.n547 10.6151
R1614 B.n550 B.n549 10.6151
R1615 B.n551 B.n550 10.6151
R1616 B.n552 B.n551 10.6151
R1617 B.n554 B.n552 10.6151
R1618 B.n555 B.n554 10.6151
R1619 B.n556 B.n555 10.6151
R1620 B.n557 B.n556 10.6151
R1621 B.n559 B.n557 10.6151
R1622 B.n560 B.n559 10.6151
R1623 B.n561 B.n560 10.6151
R1624 B.n562 B.n561 10.6151
R1625 B.n564 B.n562 10.6151
R1626 B.n565 B.n564 10.6151
R1627 B.n566 B.n565 10.6151
R1628 B.n567 B.n566 10.6151
R1629 B.n569 B.n567 10.6151
R1630 B.n570 B.n569 10.6151
R1631 B.n327 B.n277 10.6151
R1632 B.n328 B.n327 10.6151
R1633 B.n329 B.n328 10.6151
R1634 B.n329 B.n323 10.6151
R1635 B.n335 B.n323 10.6151
R1636 B.n336 B.n335 10.6151
R1637 B.n337 B.n336 10.6151
R1638 B.n337 B.n321 10.6151
R1639 B.n343 B.n321 10.6151
R1640 B.n344 B.n343 10.6151
R1641 B.n345 B.n344 10.6151
R1642 B.n345 B.n319 10.6151
R1643 B.n351 B.n319 10.6151
R1644 B.n352 B.n351 10.6151
R1645 B.n353 B.n352 10.6151
R1646 B.n353 B.n317 10.6151
R1647 B.n359 B.n317 10.6151
R1648 B.n360 B.n359 10.6151
R1649 B.n361 B.n360 10.6151
R1650 B.n361 B.n315 10.6151
R1651 B.n367 B.n315 10.6151
R1652 B.n368 B.n367 10.6151
R1653 B.n369 B.n368 10.6151
R1654 B.n369 B.n313 10.6151
R1655 B.n375 B.n313 10.6151
R1656 B.n376 B.n375 10.6151
R1657 B.n377 B.n376 10.6151
R1658 B.n377 B.n311 10.6151
R1659 B.n383 B.n311 10.6151
R1660 B.n384 B.n383 10.6151
R1661 B.n385 B.n384 10.6151
R1662 B.n385 B.n309 10.6151
R1663 B.n391 B.n309 10.6151
R1664 B.n392 B.n391 10.6151
R1665 B.n394 B.n305 10.6151
R1666 B.n400 B.n305 10.6151
R1667 B.n401 B.n400 10.6151
R1668 B.n402 B.n401 10.6151
R1669 B.n402 B.n303 10.6151
R1670 B.n408 B.n303 10.6151
R1671 B.n409 B.n408 10.6151
R1672 B.n410 B.n409 10.6151
R1673 B.n410 B.n301 10.6151
R1674 B.n417 B.n416 10.6151
R1675 B.n418 B.n417 10.6151
R1676 B.n418 B.n296 10.6151
R1677 B.n424 B.n296 10.6151
R1678 B.n425 B.n424 10.6151
R1679 B.n426 B.n425 10.6151
R1680 B.n426 B.n294 10.6151
R1681 B.n432 B.n294 10.6151
R1682 B.n433 B.n432 10.6151
R1683 B.n434 B.n433 10.6151
R1684 B.n434 B.n292 10.6151
R1685 B.n440 B.n292 10.6151
R1686 B.n441 B.n440 10.6151
R1687 B.n442 B.n441 10.6151
R1688 B.n442 B.n290 10.6151
R1689 B.n448 B.n290 10.6151
R1690 B.n449 B.n448 10.6151
R1691 B.n450 B.n449 10.6151
R1692 B.n450 B.n288 10.6151
R1693 B.n456 B.n288 10.6151
R1694 B.n457 B.n456 10.6151
R1695 B.n458 B.n457 10.6151
R1696 B.n458 B.n286 10.6151
R1697 B.n464 B.n286 10.6151
R1698 B.n465 B.n464 10.6151
R1699 B.n466 B.n465 10.6151
R1700 B.n466 B.n284 10.6151
R1701 B.n472 B.n284 10.6151
R1702 B.n473 B.n472 10.6151
R1703 B.n474 B.n473 10.6151
R1704 B.n474 B.n282 10.6151
R1705 B.n282 B.n281 10.6151
R1706 B.n481 B.n281 10.6151
R1707 B.n482 B.n481 10.6151
R1708 B.n488 B.n487 10.6151
R1709 B.n489 B.n488 10.6151
R1710 B.n489 B.n269 10.6151
R1711 B.n499 B.n269 10.6151
R1712 B.n500 B.n499 10.6151
R1713 B.n501 B.n500 10.6151
R1714 B.n501 B.n261 10.6151
R1715 B.n511 B.n261 10.6151
R1716 B.n512 B.n511 10.6151
R1717 B.n513 B.n512 10.6151
R1718 B.n513 B.n253 10.6151
R1719 B.n523 B.n253 10.6151
R1720 B.n524 B.n523 10.6151
R1721 B.n525 B.n524 10.6151
R1722 B.n525 B.n245 10.6151
R1723 B.n537 B.n245 10.6151
R1724 B.n538 B.n537 10.6151
R1725 B.n539 B.n538 10.6151
R1726 B.n539 B.n0 10.6151
R1727 B.n611 B.n1 10.6151
R1728 B.n611 B.n610 10.6151
R1729 B.n610 B.n609 10.6151
R1730 B.n609 B.n9 10.6151
R1731 B.n603 B.n9 10.6151
R1732 B.n603 B.n602 10.6151
R1733 B.n602 B.n601 10.6151
R1734 B.n601 B.n17 10.6151
R1735 B.n595 B.n17 10.6151
R1736 B.n595 B.n594 10.6151
R1737 B.n594 B.n593 10.6151
R1738 B.n593 B.n24 10.6151
R1739 B.n587 B.n24 10.6151
R1740 B.n587 B.n586 10.6151
R1741 B.n586 B.n585 10.6151
R1742 B.n585 B.n31 10.6151
R1743 B.n579 B.n31 10.6151
R1744 B.n579 B.n578 10.6151
R1745 B.n578 B.n577 10.6151
R1746 B.n534 B.t1 10.1622
R1747 B.n11 B.t4 10.1622
R1748 B.n153 B.n152 9.36635
R1749 B.n175 B.n174 9.36635
R1750 B.n393 B.n392 9.36635
R1751 B.n416 B.n300 9.36635
R1752 B.t0 B.n247 8.7105
R1753 B.n606 B.t5 8.7105
R1754 B.n515 B.t2 2.90383
R1755 B.t20 B.n597 2.90383
R1756 B.n617 B.n0 2.81026
R1757 B.n617 B.n1 2.81026
R1758 B.n154 B.n153 1.24928
R1759 B.n174 B.n173 1.24928
R1760 B.n394 B.n393 1.24928
R1761 B.n301 B.n300 1.24928
R1762 VP.n4 VP.t3 599.885
R1763 VP.n10 VP.t6 578.903
R1764 VP.n1 VP.t2 578.903
R1765 VP.n15 VP.t4 578.903
R1766 VP.n16 VP.t1 578.903
R1767 VP.n8 VP.t5 578.903
R1768 VP.n7 VP.t7 578.903
R1769 VP.n3 VP.t0 578.903
R1770 VP.n17 VP.n16 161.3
R1771 VP.n6 VP.n5 161.3
R1772 VP.n7 VP.n2 161.3
R1773 VP.n9 VP.n8 161.3
R1774 VP.n15 VP.n0 161.3
R1775 VP.n14 VP.n13 161.3
R1776 VP.n12 VP.n1 161.3
R1777 VP.n11 VP.n10 161.3
R1778 VP.n5 VP.n4 70.4033
R1779 VP.n10 VP.n1 48.2005
R1780 VP.n16 VP.n15 48.2005
R1781 VP.n8 VP.n7 48.2005
R1782 VP.n11 VP.n9 39.4323
R1783 VP.n14 VP.n1 24.1005
R1784 VP.n15 VP.n14 24.1005
R1785 VP.n6 VP.n3 24.1005
R1786 VP.n7 VP.n6 24.1005
R1787 VP.n4 VP.n3 20.9576
R1788 VP.n5 VP.n2 0.189894
R1789 VP.n9 VP.n2 0.189894
R1790 VP.n12 VP.n11 0.189894
R1791 VP.n13 VP.n12 0.189894
R1792 VP.n13 VP.n0 0.189894
R1793 VP.n17 VP.n0 0.189894
R1794 VP VP.n17 0.0516364
R1795 VDD1 VDD1.n0 61.4961
R1796 VDD1.n3 VDD1.n2 61.3824
R1797 VDD1.n3 VDD1.n1 61.3824
R1798 VDD1.n5 VDD1.n4 61.0886
R1799 VDD1.n5 VDD1.n3 35.9578
R1800 VDD1.n4 VDD1.t0 2.00455
R1801 VDD1.n4 VDD1.t2 2.00455
R1802 VDD1.n0 VDD1.t4 2.00455
R1803 VDD1.n0 VDD1.t7 2.00455
R1804 VDD1.n2 VDD1.t3 2.00455
R1805 VDD1.n2 VDD1.t6 2.00455
R1806 VDD1.n1 VDD1.t1 2.00455
R1807 VDD1.n1 VDD1.t5 2.00455
R1808 VDD1 VDD1.n5 0.291448
C0 VN VTAIL 3.49325f
C1 VN VDD1 0.147599f
C2 VP VN 4.67907f
C3 VN VDD2 3.73614f
C4 VDD1 VTAIL 11.198701f
C5 VP VTAIL 3.50736f
C6 VDD2 VTAIL 11.238901f
C7 VP VDD1 3.882f
C8 VDD2 VDD1 0.71873f
C9 VP VDD2 0.293785f
C10 VDD2 B 3.126164f
C11 VDD1 B 3.340829f
C12 VTAIL B 7.521987f
C13 VN B 7.59354f
C14 VP B 5.62648f
C15 VDD1.t4 B 0.229696f
C16 VDD1.t7 B 0.229696f
C17 VDD1.n0 B 2.02136f
C18 VDD1.t1 B 0.229696f
C19 VDD1.t5 B 0.229696f
C20 VDD1.n1 B 2.02066f
C21 VDD1.t3 B 0.229696f
C22 VDD1.t6 B 0.229696f
C23 VDD1.n2 B 2.02066f
C24 VDD1.n3 B 2.31517f
C25 VDD1.t0 B 0.229696f
C26 VDD1.t2 B 0.229696f
C27 VDD1.n4 B 2.01898f
C28 VDD1.n5 B 2.44367f
C29 VP.n0 B 0.050709f
C30 VP.t2 B 0.688727f
C31 VP.n1 B 0.293839f
C32 VP.n2 B 0.050709f
C33 VP.t5 B 0.688727f
C34 VP.t7 B 0.688727f
C35 VP.t0 B 0.688727f
C36 VP.n3 B 0.293839f
C37 VP.t3 B 0.698827f
C38 VP.n4 B 0.278963f
C39 VP.n5 B 0.164565f
C40 VP.n6 B 0.011507f
C41 VP.n7 B 0.293839f
C42 VP.n8 B 0.28868f
C43 VP.n9 B 1.87984f
C44 VP.t6 B 0.688727f
C45 VP.n10 B 0.28868f
C46 VP.n11 B 1.92594f
C47 VP.n12 B 0.050709f
C48 VP.n13 B 0.050709f
C49 VP.n14 B 0.011507f
C50 VP.t4 B 0.688727f
C51 VP.n15 B 0.293839f
C52 VP.t1 B 0.688727f
C53 VP.n16 B 0.28868f
C54 VP.n17 B 0.039298f
C55 VTAIL.t8 B 0.169569f
C56 VTAIL.t9 B 0.169569f
C57 VTAIL.n0 B 1.42508f
C58 VTAIL.n1 B 0.267073f
C59 VTAIL.n2 B 0.027597f
C60 VTAIL.n3 B 0.021719f
C61 VTAIL.n4 B 0.011671f
C62 VTAIL.n5 B 0.027585f
C63 VTAIL.n6 B 0.012357f
C64 VTAIL.n7 B 0.021719f
C65 VTAIL.n8 B 0.012014f
C66 VTAIL.n9 B 0.027585f
C67 VTAIL.n10 B 0.012357f
C68 VTAIL.n11 B 0.021719f
C69 VTAIL.n12 B 0.011671f
C70 VTAIL.n13 B 0.027585f
C71 VTAIL.n14 B 0.012357f
C72 VTAIL.n15 B 0.021719f
C73 VTAIL.n16 B 0.011671f
C74 VTAIL.n17 B 0.020689f
C75 VTAIL.n18 B 0.019501f
C76 VTAIL.t13 B 0.046343f
C77 VTAIL.n19 B 0.138915f
C78 VTAIL.n20 B 0.890874f
C79 VTAIL.n21 B 0.011671f
C80 VTAIL.n22 B 0.012357f
C81 VTAIL.n23 B 0.027585f
C82 VTAIL.n24 B 0.027585f
C83 VTAIL.n25 B 0.012357f
C84 VTAIL.n26 B 0.011671f
C85 VTAIL.n27 B 0.021719f
C86 VTAIL.n28 B 0.021719f
C87 VTAIL.n29 B 0.011671f
C88 VTAIL.n30 B 0.012357f
C89 VTAIL.n31 B 0.027585f
C90 VTAIL.n32 B 0.027585f
C91 VTAIL.n33 B 0.012357f
C92 VTAIL.n34 B 0.011671f
C93 VTAIL.n35 B 0.021719f
C94 VTAIL.n36 B 0.021719f
C95 VTAIL.n37 B 0.011671f
C96 VTAIL.n38 B 0.011671f
C97 VTAIL.n39 B 0.012357f
C98 VTAIL.n40 B 0.027585f
C99 VTAIL.n41 B 0.027585f
C100 VTAIL.n42 B 0.027585f
C101 VTAIL.n43 B 0.012014f
C102 VTAIL.n44 B 0.011671f
C103 VTAIL.n45 B 0.021719f
C104 VTAIL.n46 B 0.021719f
C105 VTAIL.n47 B 0.011671f
C106 VTAIL.n48 B 0.012357f
C107 VTAIL.n49 B 0.027585f
C108 VTAIL.n50 B 0.054535f
C109 VTAIL.n51 B 0.012357f
C110 VTAIL.n52 B 0.011671f
C111 VTAIL.n53 B 0.047828f
C112 VTAIL.n54 B 0.029907f
C113 VTAIL.n55 B 0.098958f
C114 VTAIL.n56 B 0.027597f
C115 VTAIL.n57 B 0.021719f
C116 VTAIL.n58 B 0.011671f
C117 VTAIL.n59 B 0.027585f
C118 VTAIL.n60 B 0.012357f
C119 VTAIL.n61 B 0.021719f
C120 VTAIL.n62 B 0.012014f
C121 VTAIL.n63 B 0.027585f
C122 VTAIL.n64 B 0.012357f
C123 VTAIL.n65 B 0.021719f
C124 VTAIL.n66 B 0.011671f
C125 VTAIL.n67 B 0.027585f
C126 VTAIL.n68 B 0.012357f
C127 VTAIL.n69 B 0.021719f
C128 VTAIL.n70 B 0.011671f
C129 VTAIL.n71 B 0.020689f
C130 VTAIL.n72 B 0.019501f
C131 VTAIL.t1 B 0.046343f
C132 VTAIL.n73 B 0.138915f
C133 VTAIL.n74 B 0.890874f
C134 VTAIL.n75 B 0.011671f
C135 VTAIL.n76 B 0.012357f
C136 VTAIL.n77 B 0.027585f
C137 VTAIL.n78 B 0.027585f
C138 VTAIL.n79 B 0.012357f
C139 VTAIL.n80 B 0.011671f
C140 VTAIL.n81 B 0.021719f
C141 VTAIL.n82 B 0.021719f
C142 VTAIL.n83 B 0.011671f
C143 VTAIL.n84 B 0.012357f
C144 VTAIL.n85 B 0.027585f
C145 VTAIL.n86 B 0.027585f
C146 VTAIL.n87 B 0.012357f
C147 VTAIL.n88 B 0.011671f
C148 VTAIL.n89 B 0.021719f
C149 VTAIL.n90 B 0.021719f
C150 VTAIL.n91 B 0.011671f
C151 VTAIL.n92 B 0.011671f
C152 VTAIL.n93 B 0.012357f
C153 VTAIL.n94 B 0.027585f
C154 VTAIL.n95 B 0.027585f
C155 VTAIL.n96 B 0.027585f
C156 VTAIL.n97 B 0.012014f
C157 VTAIL.n98 B 0.011671f
C158 VTAIL.n99 B 0.021719f
C159 VTAIL.n100 B 0.021719f
C160 VTAIL.n101 B 0.011671f
C161 VTAIL.n102 B 0.012357f
C162 VTAIL.n103 B 0.027585f
C163 VTAIL.n104 B 0.054535f
C164 VTAIL.n105 B 0.012357f
C165 VTAIL.n106 B 0.011671f
C166 VTAIL.n107 B 0.047828f
C167 VTAIL.n108 B 0.029907f
C168 VTAIL.n109 B 0.098958f
C169 VTAIL.t14 B 0.169569f
C170 VTAIL.t0 B 0.169569f
C171 VTAIL.n110 B 1.42508f
C172 VTAIL.n111 B 0.311868f
C173 VTAIL.n112 B 0.027597f
C174 VTAIL.n113 B 0.021719f
C175 VTAIL.n114 B 0.011671f
C176 VTAIL.n115 B 0.027585f
C177 VTAIL.n116 B 0.012357f
C178 VTAIL.n117 B 0.021719f
C179 VTAIL.n118 B 0.012014f
C180 VTAIL.n119 B 0.027585f
C181 VTAIL.n120 B 0.012357f
C182 VTAIL.n121 B 0.021719f
C183 VTAIL.n122 B 0.011671f
C184 VTAIL.n123 B 0.027585f
C185 VTAIL.n124 B 0.012357f
C186 VTAIL.n125 B 0.021719f
C187 VTAIL.n126 B 0.011671f
C188 VTAIL.n127 B 0.020689f
C189 VTAIL.n128 B 0.019501f
C190 VTAIL.t2 B 0.046343f
C191 VTAIL.n129 B 0.138915f
C192 VTAIL.n130 B 0.890874f
C193 VTAIL.n131 B 0.011671f
C194 VTAIL.n132 B 0.012357f
C195 VTAIL.n133 B 0.027585f
C196 VTAIL.n134 B 0.027585f
C197 VTAIL.n135 B 0.012357f
C198 VTAIL.n136 B 0.011671f
C199 VTAIL.n137 B 0.021719f
C200 VTAIL.n138 B 0.021719f
C201 VTAIL.n139 B 0.011671f
C202 VTAIL.n140 B 0.012357f
C203 VTAIL.n141 B 0.027585f
C204 VTAIL.n142 B 0.027585f
C205 VTAIL.n143 B 0.012357f
C206 VTAIL.n144 B 0.011671f
C207 VTAIL.n145 B 0.021719f
C208 VTAIL.n146 B 0.021719f
C209 VTAIL.n147 B 0.011671f
C210 VTAIL.n148 B 0.011671f
C211 VTAIL.n149 B 0.012357f
C212 VTAIL.n150 B 0.027585f
C213 VTAIL.n151 B 0.027585f
C214 VTAIL.n152 B 0.027585f
C215 VTAIL.n153 B 0.012014f
C216 VTAIL.n154 B 0.011671f
C217 VTAIL.n155 B 0.021719f
C218 VTAIL.n156 B 0.021719f
C219 VTAIL.n157 B 0.011671f
C220 VTAIL.n158 B 0.012357f
C221 VTAIL.n159 B 0.027585f
C222 VTAIL.n160 B 0.054535f
C223 VTAIL.n161 B 0.012357f
C224 VTAIL.n162 B 0.011671f
C225 VTAIL.n163 B 0.047828f
C226 VTAIL.n164 B 0.029907f
C227 VTAIL.n165 B 1.00603f
C228 VTAIL.n166 B 0.027597f
C229 VTAIL.n167 B 0.021719f
C230 VTAIL.n168 B 0.011671f
C231 VTAIL.n169 B 0.027585f
C232 VTAIL.n170 B 0.012357f
C233 VTAIL.n171 B 0.021719f
C234 VTAIL.n172 B 0.012014f
C235 VTAIL.n173 B 0.027585f
C236 VTAIL.n174 B 0.011671f
C237 VTAIL.n175 B 0.012357f
C238 VTAIL.n176 B 0.021719f
C239 VTAIL.n177 B 0.011671f
C240 VTAIL.n178 B 0.027585f
C241 VTAIL.n179 B 0.012357f
C242 VTAIL.n180 B 0.021719f
C243 VTAIL.n181 B 0.011671f
C244 VTAIL.n182 B 0.020689f
C245 VTAIL.n183 B 0.019501f
C246 VTAIL.t10 B 0.046343f
C247 VTAIL.n184 B 0.138915f
C248 VTAIL.n185 B 0.890874f
C249 VTAIL.n186 B 0.011671f
C250 VTAIL.n187 B 0.012357f
C251 VTAIL.n188 B 0.027585f
C252 VTAIL.n189 B 0.027585f
C253 VTAIL.n190 B 0.012357f
C254 VTAIL.n191 B 0.011671f
C255 VTAIL.n192 B 0.021719f
C256 VTAIL.n193 B 0.021719f
C257 VTAIL.n194 B 0.011671f
C258 VTAIL.n195 B 0.012357f
C259 VTAIL.n196 B 0.027585f
C260 VTAIL.n197 B 0.027585f
C261 VTAIL.n198 B 0.012357f
C262 VTAIL.n199 B 0.011671f
C263 VTAIL.n200 B 0.021719f
C264 VTAIL.n201 B 0.021719f
C265 VTAIL.n202 B 0.011671f
C266 VTAIL.n203 B 0.012357f
C267 VTAIL.n204 B 0.027585f
C268 VTAIL.n205 B 0.027585f
C269 VTAIL.n206 B 0.027585f
C270 VTAIL.n207 B 0.012014f
C271 VTAIL.n208 B 0.011671f
C272 VTAIL.n209 B 0.021719f
C273 VTAIL.n210 B 0.021719f
C274 VTAIL.n211 B 0.011671f
C275 VTAIL.n212 B 0.012357f
C276 VTAIL.n213 B 0.027585f
C277 VTAIL.n214 B 0.054535f
C278 VTAIL.n215 B 0.012357f
C279 VTAIL.n216 B 0.011671f
C280 VTAIL.n217 B 0.047828f
C281 VTAIL.n218 B 0.029907f
C282 VTAIL.n219 B 1.00603f
C283 VTAIL.t7 B 0.169569f
C284 VTAIL.t12 B 0.169569f
C285 VTAIL.n220 B 1.42509f
C286 VTAIL.n221 B 0.311858f
C287 VTAIL.n222 B 0.027597f
C288 VTAIL.n223 B 0.021719f
C289 VTAIL.n224 B 0.011671f
C290 VTAIL.n225 B 0.027585f
C291 VTAIL.n226 B 0.012357f
C292 VTAIL.n227 B 0.021719f
C293 VTAIL.n228 B 0.012014f
C294 VTAIL.n229 B 0.027585f
C295 VTAIL.n230 B 0.011671f
C296 VTAIL.n231 B 0.012357f
C297 VTAIL.n232 B 0.021719f
C298 VTAIL.n233 B 0.011671f
C299 VTAIL.n234 B 0.027585f
C300 VTAIL.n235 B 0.012357f
C301 VTAIL.n236 B 0.021719f
C302 VTAIL.n237 B 0.011671f
C303 VTAIL.n238 B 0.020689f
C304 VTAIL.n239 B 0.019501f
C305 VTAIL.t11 B 0.046343f
C306 VTAIL.n240 B 0.138915f
C307 VTAIL.n241 B 0.890874f
C308 VTAIL.n242 B 0.011671f
C309 VTAIL.n243 B 0.012357f
C310 VTAIL.n244 B 0.027585f
C311 VTAIL.n245 B 0.027585f
C312 VTAIL.n246 B 0.012357f
C313 VTAIL.n247 B 0.011671f
C314 VTAIL.n248 B 0.021719f
C315 VTAIL.n249 B 0.021719f
C316 VTAIL.n250 B 0.011671f
C317 VTAIL.n251 B 0.012357f
C318 VTAIL.n252 B 0.027585f
C319 VTAIL.n253 B 0.027585f
C320 VTAIL.n254 B 0.012357f
C321 VTAIL.n255 B 0.011671f
C322 VTAIL.n256 B 0.021719f
C323 VTAIL.n257 B 0.021719f
C324 VTAIL.n258 B 0.011671f
C325 VTAIL.n259 B 0.012357f
C326 VTAIL.n260 B 0.027585f
C327 VTAIL.n261 B 0.027585f
C328 VTAIL.n262 B 0.027585f
C329 VTAIL.n263 B 0.012014f
C330 VTAIL.n264 B 0.011671f
C331 VTAIL.n265 B 0.021719f
C332 VTAIL.n266 B 0.021719f
C333 VTAIL.n267 B 0.011671f
C334 VTAIL.n268 B 0.012357f
C335 VTAIL.n269 B 0.027585f
C336 VTAIL.n270 B 0.054535f
C337 VTAIL.n271 B 0.012357f
C338 VTAIL.n272 B 0.011671f
C339 VTAIL.n273 B 0.047828f
C340 VTAIL.n274 B 0.029907f
C341 VTAIL.n275 B 0.098958f
C342 VTAIL.n276 B 0.027597f
C343 VTAIL.n277 B 0.021719f
C344 VTAIL.n278 B 0.011671f
C345 VTAIL.n279 B 0.027585f
C346 VTAIL.n280 B 0.012357f
C347 VTAIL.n281 B 0.021719f
C348 VTAIL.n282 B 0.012014f
C349 VTAIL.n283 B 0.027585f
C350 VTAIL.n284 B 0.011671f
C351 VTAIL.n285 B 0.012357f
C352 VTAIL.n286 B 0.021719f
C353 VTAIL.n287 B 0.011671f
C354 VTAIL.n288 B 0.027585f
C355 VTAIL.n289 B 0.012357f
C356 VTAIL.n290 B 0.021719f
C357 VTAIL.n291 B 0.011671f
C358 VTAIL.n292 B 0.020689f
C359 VTAIL.n293 B 0.019501f
C360 VTAIL.t4 B 0.046343f
C361 VTAIL.n294 B 0.138915f
C362 VTAIL.n295 B 0.890874f
C363 VTAIL.n296 B 0.011671f
C364 VTAIL.n297 B 0.012357f
C365 VTAIL.n298 B 0.027585f
C366 VTAIL.n299 B 0.027585f
C367 VTAIL.n300 B 0.012357f
C368 VTAIL.n301 B 0.011671f
C369 VTAIL.n302 B 0.021719f
C370 VTAIL.n303 B 0.021719f
C371 VTAIL.n304 B 0.011671f
C372 VTAIL.n305 B 0.012357f
C373 VTAIL.n306 B 0.027585f
C374 VTAIL.n307 B 0.027585f
C375 VTAIL.n308 B 0.012357f
C376 VTAIL.n309 B 0.011671f
C377 VTAIL.n310 B 0.021719f
C378 VTAIL.n311 B 0.021719f
C379 VTAIL.n312 B 0.011671f
C380 VTAIL.n313 B 0.012357f
C381 VTAIL.n314 B 0.027585f
C382 VTAIL.n315 B 0.027585f
C383 VTAIL.n316 B 0.027585f
C384 VTAIL.n317 B 0.012014f
C385 VTAIL.n318 B 0.011671f
C386 VTAIL.n319 B 0.021719f
C387 VTAIL.n320 B 0.021719f
C388 VTAIL.n321 B 0.011671f
C389 VTAIL.n322 B 0.012357f
C390 VTAIL.n323 B 0.027585f
C391 VTAIL.n324 B 0.054535f
C392 VTAIL.n325 B 0.012357f
C393 VTAIL.n326 B 0.011671f
C394 VTAIL.n327 B 0.047828f
C395 VTAIL.n328 B 0.029907f
C396 VTAIL.n329 B 0.098958f
C397 VTAIL.t5 B 0.169569f
C398 VTAIL.t3 B 0.169569f
C399 VTAIL.n330 B 1.42509f
C400 VTAIL.n331 B 0.311858f
C401 VTAIL.n332 B 0.027597f
C402 VTAIL.n333 B 0.021719f
C403 VTAIL.n334 B 0.011671f
C404 VTAIL.n335 B 0.027585f
C405 VTAIL.n336 B 0.012357f
C406 VTAIL.n337 B 0.021719f
C407 VTAIL.n338 B 0.012014f
C408 VTAIL.n339 B 0.027585f
C409 VTAIL.n340 B 0.011671f
C410 VTAIL.n341 B 0.012357f
C411 VTAIL.n342 B 0.021719f
C412 VTAIL.n343 B 0.011671f
C413 VTAIL.n344 B 0.027585f
C414 VTAIL.n345 B 0.012357f
C415 VTAIL.n346 B 0.021719f
C416 VTAIL.n347 B 0.011671f
C417 VTAIL.n348 B 0.020689f
C418 VTAIL.n349 B 0.019501f
C419 VTAIL.t15 B 0.046343f
C420 VTAIL.n350 B 0.138915f
C421 VTAIL.n351 B 0.890874f
C422 VTAIL.n352 B 0.011671f
C423 VTAIL.n353 B 0.012357f
C424 VTAIL.n354 B 0.027585f
C425 VTAIL.n355 B 0.027585f
C426 VTAIL.n356 B 0.012357f
C427 VTAIL.n357 B 0.011671f
C428 VTAIL.n358 B 0.021719f
C429 VTAIL.n359 B 0.021719f
C430 VTAIL.n360 B 0.011671f
C431 VTAIL.n361 B 0.012357f
C432 VTAIL.n362 B 0.027585f
C433 VTAIL.n363 B 0.027585f
C434 VTAIL.n364 B 0.012357f
C435 VTAIL.n365 B 0.011671f
C436 VTAIL.n366 B 0.021719f
C437 VTAIL.n367 B 0.021719f
C438 VTAIL.n368 B 0.011671f
C439 VTAIL.n369 B 0.012357f
C440 VTAIL.n370 B 0.027585f
C441 VTAIL.n371 B 0.027585f
C442 VTAIL.n372 B 0.027585f
C443 VTAIL.n373 B 0.012014f
C444 VTAIL.n374 B 0.011671f
C445 VTAIL.n375 B 0.021719f
C446 VTAIL.n376 B 0.021719f
C447 VTAIL.n377 B 0.011671f
C448 VTAIL.n378 B 0.012357f
C449 VTAIL.n379 B 0.027585f
C450 VTAIL.n380 B 0.054535f
C451 VTAIL.n381 B 0.012357f
C452 VTAIL.n382 B 0.011671f
C453 VTAIL.n383 B 0.047828f
C454 VTAIL.n384 B 0.029907f
C455 VTAIL.n385 B 1.00603f
C456 VTAIL.n386 B 0.027597f
C457 VTAIL.n387 B 0.021719f
C458 VTAIL.n388 B 0.011671f
C459 VTAIL.n389 B 0.027585f
C460 VTAIL.n390 B 0.012357f
C461 VTAIL.n391 B 0.021719f
C462 VTAIL.n392 B 0.012014f
C463 VTAIL.n393 B 0.027585f
C464 VTAIL.n394 B 0.012357f
C465 VTAIL.n395 B 0.021719f
C466 VTAIL.n396 B 0.011671f
C467 VTAIL.n397 B 0.027585f
C468 VTAIL.n398 B 0.012357f
C469 VTAIL.n399 B 0.021719f
C470 VTAIL.n400 B 0.011671f
C471 VTAIL.n401 B 0.020689f
C472 VTAIL.n402 B 0.019501f
C473 VTAIL.t6 B 0.046343f
C474 VTAIL.n403 B 0.138915f
C475 VTAIL.n404 B 0.890874f
C476 VTAIL.n405 B 0.011671f
C477 VTAIL.n406 B 0.012357f
C478 VTAIL.n407 B 0.027585f
C479 VTAIL.n408 B 0.027585f
C480 VTAIL.n409 B 0.012357f
C481 VTAIL.n410 B 0.011671f
C482 VTAIL.n411 B 0.021719f
C483 VTAIL.n412 B 0.021719f
C484 VTAIL.n413 B 0.011671f
C485 VTAIL.n414 B 0.012357f
C486 VTAIL.n415 B 0.027585f
C487 VTAIL.n416 B 0.027585f
C488 VTAIL.n417 B 0.012357f
C489 VTAIL.n418 B 0.011671f
C490 VTAIL.n419 B 0.021719f
C491 VTAIL.n420 B 0.021719f
C492 VTAIL.n421 B 0.011671f
C493 VTAIL.n422 B 0.011671f
C494 VTAIL.n423 B 0.012357f
C495 VTAIL.n424 B 0.027585f
C496 VTAIL.n425 B 0.027585f
C497 VTAIL.n426 B 0.027585f
C498 VTAIL.n427 B 0.012014f
C499 VTAIL.n428 B 0.011671f
C500 VTAIL.n429 B 0.021719f
C501 VTAIL.n430 B 0.021719f
C502 VTAIL.n431 B 0.011671f
C503 VTAIL.n432 B 0.012357f
C504 VTAIL.n433 B 0.027585f
C505 VTAIL.n434 B 0.054535f
C506 VTAIL.n435 B 0.012357f
C507 VTAIL.n436 B 0.011671f
C508 VTAIL.n437 B 0.047828f
C509 VTAIL.n438 B 0.029907f
C510 VTAIL.n439 B 1.00196f
C511 VDD2.t1 B 0.228296f
C512 VDD2.t3 B 0.228296f
C513 VDD2.n0 B 2.00835f
C514 VDD2.t7 B 0.228296f
C515 VDD2.t2 B 0.228296f
C516 VDD2.n1 B 2.00835f
C517 VDD2.n2 B 2.23832f
C518 VDD2.t4 B 0.228296f
C519 VDD2.t6 B 0.228296f
C520 VDD2.n3 B 2.00669f
C521 VDD2.n4 B 2.39448f
C522 VDD2.t0 B 0.228296f
C523 VDD2.t5 B 0.228296f
C524 VDD2.n5 B 2.00832f
C525 VN.n0 B 0.049579f
C526 VN.t5 B 0.673376f
C527 VN.n1 B 0.28729f
C528 VN.t0 B 0.683251f
C529 VN.n2 B 0.272745f
C530 VN.n3 B 0.160897f
C531 VN.n4 B 0.01125f
C532 VN.t4 B 0.673376f
C533 VN.n5 B 0.28729f
C534 VN.t7 B 0.673376f
C535 VN.n6 B 0.282246f
C536 VN.n7 B 0.038422f
C537 VN.n8 B 0.049579f
C538 VN.t1 B 0.673376f
C539 VN.n9 B 0.28729f
C540 VN.t2 B 0.683251f
C541 VN.n10 B 0.272745f
C542 VN.n11 B 0.160897f
C543 VN.n12 B 0.01125f
C544 VN.t6 B 0.673376f
C545 VN.n13 B 0.28729f
C546 VN.t3 B 0.673376f
C547 VN.n14 B 0.282246f
C548 VN.n15 B 1.87062f
.ends

