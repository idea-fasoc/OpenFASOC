* NGSPICE file created from diff_pair_sample_1739.ext - technology: sky130A

.subckt diff_pair_sample_1739 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=0 ps=0 w=4.78 l=3.74
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=1.8642 ps=10.34 w=4.78 l=3.74
X2 B.t8 B.t6 B.t7 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=0 ps=0 w=4.78 l=3.74
X3 B.t5 B.t3 B.t4 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=0 ps=0 w=4.78 l=3.74
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=1.8642 ps=10.34 w=4.78 l=3.74
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=1.8642 ps=10.34 w=4.78 l=3.74
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=1.8642 ps=10.34 w=4.78 l=3.74
X7 B.t2 B.t0 B.t1 w_n2598_n1924# sky130_fd_pr__pfet_01v8 ad=1.8642 pd=10.34 as=0 ps=0 w=4.78 l=3.74
R0 B.n346 B.n47 585
R1 B.n348 B.n347 585
R2 B.n349 B.n46 585
R3 B.n351 B.n350 585
R4 B.n352 B.n45 585
R5 B.n354 B.n353 585
R6 B.n355 B.n44 585
R7 B.n357 B.n356 585
R8 B.n358 B.n43 585
R9 B.n360 B.n359 585
R10 B.n361 B.n42 585
R11 B.n363 B.n362 585
R12 B.n364 B.n41 585
R13 B.n366 B.n365 585
R14 B.n367 B.n40 585
R15 B.n369 B.n368 585
R16 B.n370 B.n39 585
R17 B.n372 B.n371 585
R18 B.n373 B.n38 585
R19 B.n375 B.n374 585
R20 B.n377 B.n35 585
R21 B.n379 B.n378 585
R22 B.n380 B.n34 585
R23 B.n382 B.n381 585
R24 B.n383 B.n33 585
R25 B.n385 B.n384 585
R26 B.n386 B.n32 585
R27 B.n388 B.n387 585
R28 B.n389 B.n31 585
R29 B.n391 B.n390 585
R30 B.n393 B.n392 585
R31 B.n394 B.n27 585
R32 B.n396 B.n395 585
R33 B.n397 B.n26 585
R34 B.n399 B.n398 585
R35 B.n400 B.n25 585
R36 B.n402 B.n401 585
R37 B.n403 B.n24 585
R38 B.n405 B.n404 585
R39 B.n406 B.n23 585
R40 B.n408 B.n407 585
R41 B.n409 B.n22 585
R42 B.n411 B.n410 585
R43 B.n412 B.n21 585
R44 B.n414 B.n413 585
R45 B.n415 B.n20 585
R46 B.n417 B.n416 585
R47 B.n418 B.n19 585
R48 B.n420 B.n419 585
R49 B.n421 B.n18 585
R50 B.n345 B.n344 585
R51 B.n343 B.n48 585
R52 B.n342 B.n341 585
R53 B.n340 B.n49 585
R54 B.n339 B.n338 585
R55 B.n337 B.n50 585
R56 B.n336 B.n335 585
R57 B.n334 B.n51 585
R58 B.n333 B.n332 585
R59 B.n331 B.n52 585
R60 B.n330 B.n329 585
R61 B.n328 B.n53 585
R62 B.n327 B.n326 585
R63 B.n325 B.n54 585
R64 B.n324 B.n323 585
R65 B.n322 B.n55 585
R66 B.n321 B.n320 585
R67 B.n319 B.n56 585
R68 B.n318 B.n317 585
R69 B.n316 B.n57 585
R70 B.n315 B.n314 585
R71 B.n313 B.n58 585
R72 B.n312 B.n311 585
R73 B.n310 B.n59 585
R74 B.n309 B.n308 585
R75 B.n307 B.n60 585
R76 B.n306 B.n305 585
R77 B.n304 B.n61 585
R78 B.n303 B.n302 585
R79 B.n301 B.n62 585
R80 B.n300 B.n299 585
R81 B.n298 B.n63 585
R82 B.n297 B.n296 585
R83 B.n295 B.n64 585
R84 B.n294 B.n293 585
R85 B.n292 B.n65 585
R86 B.n291 B.n290 585
R87 B.n289 B.n66 585
R88 B.n288 B.n287 585
R89 B.n286 B.n67 585
R90 B.n285 B.n284 585
R91 B.n283 B.n68 585
R92 B.n282 B.n281 585
R93 B.n280 B.n69 585
R94 B.n279 B.n278 585
R95 B.n277 B.n70 585
R96 B.n276 B.n275 585
R97 B.n274 B.n71 585
R98 B.n273 B.n272 585
R99 B.n271 B.n72 585
R100 B.n270 B.n269 585
R101 B.n268 B.n73 585
R102 B.n267 B.n266 585
R103 B.n265 B.n74 585
R104 B.n264 B.n263 585
R105 B.n262 B.n75 585
R106 B.n261 B.n260 585
R107 B.n259 B.n76 585
R108 B.n258 B.n257 585
R109 B.n256 B.n77 585
R110 B.n255 B.n254 585
R111 B.n253 B.n78 585
R112 B.n252 B.n251 585
R113 B.n250 B.n79 585
R114 B.n249 B.n248 585
R115 B.n172 B.n109 585
R116 B.n174 B.n173 585
R117 B.n175 B.n108 585
R118 B.n177 B.n176 585
R119 B.n178 B.n107 585
R120 B.n180 B.n179 585
R121 B.n181 B.n106 585
R122 B.n183 B.n182 585
R123 B.n184 B.n105 585
R124 B.n186 B.n185 585
R125 B.n187 B.n104 585
R126 B.n189 B.n188 585
R127 B.n190 B.n103 585
R128 B.n192 B.n191 585
R129 B.n193 B.n102 585
R130 B.n195 B.n194 585
R131 B.n196 B.n101 585
R132 B.n198 B.n197 585
R133 B.n199 B.n100 585
R134 B.n201 B.n200 585
R135 B.n203 B.n97 585
R136 B.n205 B.n204 585
R137 B.n206 B.n96 585
R138 B.n208 B.n207 585
R139 B.n209 B.n95 585
R140 B.n211 B.n210 585
R141 B.n212 B.n94 585
R142 B.n214 B.n213 585
R143 B.n215 B.n93 585
R144 B.n217 B.n216 585
R145 B.n219 B.n218 585
R146 B.n220 B.n89 585
R147 B.n222 B.n221 585
R148 B.n223 B.n88 585
R149 B.n225 B.n224 585
R150 B.n226 B.n87 585
R151 B.n228 B.n227 585
R152 B.n229 B.n86 585
R153 B.n231 B.n230 585
R154 B.n232 B.n85 585
R155 B.n234 B.n233 585
R156 B.n235 B.n84 585
R157 B.n237 B.n236 585
R158 B.n238 B.n83 585
R159 B.n240 B.n239 585
R160 B.n241 B.n82 585
R161 B.n243 B.n242 585
R162 B.n244 B.n81 585
R163 B.n246 B.n245 585
R164 B.n247 B.n80 585
R165 B.n171 B.n170 585
R166 B.n169 B.n110 585
R167 B.n168 B.n167 585
R168 B.n166 B.n111 585
R169 B.n165 B.n164 585
R170 B.n163 B.n112 585
R171 B.n162 B.n161 585
R172 B.n160 B.n113 585
R173 B.n159 B.n158 585
R174 B.n157 B.n114 585
R175 B.n156 B.n155 585
R176 B.n154 B.n115 585
R177 B.n153 B.n152 585
R178 B.n151 B.n116 585
R179 B.n150 B.n149 585
R180 B.n148 B.n117 585
R181 B.n147 B.n146 585
R182 B.n145 B.n118 585
R183 B.n144 B.n143 585
R184 B.n142 B.n119 585
R185 B.n141 B.n140 585
R186 B.n139 B.n120 585
R187 B.n138 B.n137 585
R188 B.n136 B.n121 585
R189 B.n135 B.n134 585
R190 B.n133 B.n122 585
R191 B.n132 B.n131 585
R192 B.n130 B.n123 585
R193 B.n129 B.n128 585
R194 B.n127 B.n124 585
R195 B.n126 B.n125 585
R196 B.n2 B.n0 585
R197 B.n469 B.n1 585
R198 B.n468 B.n467 585
R199 B.n466 B.n3 585
R200 B.n465 B.n464 585
R201 B.n463 B.n4 585
R202 B.n462 B.n461 585
R203 B.n460 B.n5 585
R204 B.n459 B.n458 585
R205 B.n457 B.n6 585
R206 B.n456 B.n455 585
R207 B.n454 B.n7 585
R208 B.n453 B.n452 585
R209 B.n451 B.n8 585
R210 B.n450 B.n449 585
R211 B.n448 B.n9 585
R212 B.n447 B.n446 585
R213 B.n445 B.n10 585
R214 B.n444 B.n443 585
R215 B.n442 B.n11 585
R216 B.n441 B.n440 585
R217 B.n439 B.n12 585
R218 B.n438 B.n437 585
R219 B.n436 B.n13 585
R220 B.n435 B.n434 585
R221 B.n433 B.n14 585
R222 B.n432 B.n431 585
R223 B.n430 B.n15 585
R224 B.n429 B.n428 585
R225 B.n427 B.n16 585
R226 B.n426 B.n425 585
R227 B.n424 B.n17 585
R228 B.n423 B.n422 585
R229 B.n471 B.n470 585
R230 B.n170 B.n109 535.745
R231 B.n422 B.n421 535.745
R232 B.n248 B.n247 535.745
R233 B.n344 B.n47 535.745
R234 B.n90 B.t3 240.099
R235 B.n98 B.t9 240.099
R236 B.n28 B.t6 240.099
R237 B.n36 B.t0 240.099
R238 B.n90 B.t5 194.139
R239 B.n36 B.t1 194.139
R240 B.n98 B.t11 194.136
R241 B.n28 B.t7 194.136
R242 B.n170 B.n169 163.367
R243 B.n169 B.n168 163.367
R244 B.n168 B.n111 163.367
R245 B.n164 B.n111 163.367
R246 B.n164 B.n163 163.367
R247 B.n163 B.n162 163.367
R248 B.n162 B.n113 163.367
R249 B.n158 B.n113 163.367
R250 B.n158 B.n157 163.367
R251 B.n157 B.n156 163.367
R252 B.n156 B.n115 163.367
R253 B.n152 B.n115 163.367
R254 B.n152 B.n151 163.367
R255 B.n151 B.n150 163.367
R256 B.n150 B.n117 163.367
R257 B.n146 B.n117 163.367
R258 B.n146 B.n145 163.367
R259 B.n145 B.n144 163.367
R260 B.n144 B.n119 163.367
R261 B.n140 B.n119 163.367
R262 B.n140 B.n139 163.367
R263 B.n139 B.n138 163.367
R264 B.n138 B.n121 163.367
R265 B.n134 B.n121 163.367
R266 B.n134 B.n133 163.367
R267 B.n133 B.n132 163.367
R268 B.n132 B.n123 163.367
R269 B.n128 B.n123 163.367
R270 B.n128 B.n127 163.367
R271 B.n127 B.n126 163.367
R272 B.n126 B.n2 163.367
R273 B.n470 B.n2 163.367
R274 B.n470 B.n469 163.367
R275 B.n469 B.n468 163.367
R276 B.n468 B.n3 163.367
R277 B.n464 B.n3 163.367
R278 B.n464 B.n463 163.367
R279 B.n463 B.n462 163.367
R280 B.n462 B.n5 163.367
R281 B.n458 B.n5 163.367
R282 B.n458 B.n457 163.367
R283 B.n457 B.n456 163.367
R284 B.n456 B.n7 163.367
R285 B.n452 B.n7 163.367
R286 B.n452 B.n451 163.367
R287 B.n451 B.n450 163.367
R288 B.n450 B.n9 163.367
R289 B.n446 B.n9 163.367
R290 B.n446 B.n445 163.367
R291 B.n445 B.n444 163.367
R292 B.n444 B.n11 163.367
R293 B.n440 B.n11 163.367
R294 B.n440 B.n439 163.367
R295 B.n439 B.n438 163.367
R296 B.n438 B.n13 163.367
R297 B.n434 B.n13 163.367
R298 B.n434 B.n433 163.367
R299 B.n433 B.n432 163.367
R300 B.n432 B.n15 163.367
R301 B.n428 B.n15 163.367
R302 B.n428 B.n427 163.367
R303 B.n427 B.n426 163.367
R304 B.n426 B.n17 163.367
R305 B.n422 B.n17 163.367
R306 B.n174 B.n109 163.367
R307 B.n175 B.n174 163.367
R308 B.n176 B.n175 163.367
R309 B.n176 B.n107 163.367
R310 B.n180 B.n107 163.367
R311 B.n181 B.n180 163.367
R312 B.n182 B.n181 163.367
R313 B.n182 B.n105 163.367
R314 B.n186 B.n105 163.367
R315 B.n187 B.n186 163.367
R316 B.n188 B.n187 163.367
R317 B.n188 B.n103 163.367
R318 B.n192 B.n103 163.367
R319 B.n193 B.n192 163.367
R320 B.n194 B.n193 163.367
R321 B.n194 B.n101 163.367
R322 B.n198 B.n101 163.367
R323 B.n199 B.n198 163.367
R324 B.n200 B.n199 163.367
R325 B.n200 B.n97 163.367
R326 B.n205 B.n97 163.367
R327 B.n206 B.n205 163.367
R328 B.n207 B.n206 163.367
R329 B.n207 B.n95 163.367
R330 B.n211 B.n95 163.367
R331 B.n212 B.n211 163.367
R332 B.n213 B.n212 163.367
R333 B.n213 B.n93 163.367
R334 B.n217 B.n93 163.367
R335 B.n218 B.n217 163.367
R336 B.n218 B.n89 163.367
R337 B.n222 B.n89 163.367
R338 B.n223 B.n222 163.367
R339 B.n224 B.n223 163.367
R340 B.n224 B.n87 163.367
R341 B.n228 B.n87 163.367
R342 B.n229 B.n228 163.367
R343 B.n230 B.n229 163.367
R344 B.n230 B.n85 163.367
R345 B.n234 B.n85 163.367
R346 B.n235 B.n234 163.367
R347 B.n236 B.n235 163.367
R348 B.n236 B.n83 163.367
R349 B.n240 B.n83 163.367
R350 B.n241 B.n240 163.367
R351 B.n242 B.n241 163.367
R352 B.n242 B.n81 163.367
R353 B.n246 B.n81 163.367
R354 B.n247 B.n246 163.367
R355 B.n248 B.n79 163.367
R356 B.n252 B.n79 163.367
R357 B.n253 B.n252 163.367
R358 B.n254 B.n253 163.367
R359 B.n254 B.n77 163.367
R360 B.n258 B.n77 163.367
R361 B.n259 B.n258 163.367
R362 B.n260 B.n259 163.367
R363 B.n260 B.n75 163.367
R364 B.n264 B.n75 163.367
R365 B.n265 B.n264 163.367
R366 B.n266 B.n265 163.367
R367 B.n266 B.n73 163.367
R368 B.n270 B.n73 163.367
R369 B.n271 B.n270 163.367
R370 B.n272 B.n271 163.367
R371 B.n272 B.n71 163.367
R372 B.n276 B.n71 163.367
R373 B.n277 B.n276 163.367
R374 B.n278 B.n277 163.367
R375 B.n278 B.n69 163.367
R376 B.n282 B.n69 163.367
R377 B.n283 B.n282 163.367
R378 B.n284 B.n283 163.367
R379 B.n284 B.n67 163.367
R380 B.n288 B.n67 163.367
R381 B.n289 B.n288 163.367
R382 B.n290 B.n289 163.367
R383 B.n290 B.n65 163.367
R384 B.n294 B.n65 163.367
R385 B.n295 B.n294 163.367
R386 B.n296 B.n295 163.367
R387 B.n296 B.n63 163.367
R388 B.n300 B.n63 163.367
R389 B.n301 B.n300 163.367
R390 B.n302 B.n301 163.367
R391 B.n302 B.n61 163.367
R392 B.n306 B.n61 163.367
R393 B.n307 B.n306 163.367
R394 B.n308 B.n307 163.367
R395 B.n308 B.n59 163.367
R396 B.n312 B.n59 163.367
R397 B.n313 B.n312 163.367
R398 B.n314 B.n313 163.367
R399 B.n314 B.n57 163.367
R400 B.n318 B.n57 163.367
R401 B.n319 B.n318 163.367
R402 B.n320 B.n319 163.367
R403 B.n320 B.n55 163.367
R404 B.n324 B.n55 163.367
R405 B.n325 B.n324 163.367
R406 B.n326 B.n325 163.367
R407 B.n326 B.n53 163.367
R408 B.n330 B.n53 163.367
R409 B.n331 B.n330 163.367
R410 B.n332 B.n331 163.367
R411 B.n332 B.n51 163.367
R412 B.n336 B.n51 163.367
R413 B.n337 B.n336 163.367
R414 B.n338 B.n337 163.367
R415 B.n338 B.n49 163.367
R416 B.n342 B.n49 163.367
R417 B.n343 B.n342 163.367
R418 B.n344 B.n343 163.367
R419 B.n421 B.n420 163.367
R420 B.n420 B.n19 163.367
R421 B.n416 B.n19 163.367
R422 B.n416 B.n415 163.367
R423 B.n415 B.n414 163.367
R424 B.n414 B.n21 163.367
R425 B.n410 B.n21 163.367
R426 B.n410 B.n409 163.367
R427 B.n409 B.n408 163.367
R428 B.n408 B.n23 163.367
R429 B.n404 B.n23 163.367
R430 B.n404 B.n403 163.367
R431 B.n403 B.n402 163.367
R432 B.n402 B.n25 163.367
R433 B.n398 B.n25 163.367
R434 B.n398 B.n397 163.367
R435 B.n397 B.n396 163.367
R436 B.n396 B.n27 163.367
R437 B.n392 B.n27 163.367
R438 B.n392 B.n391 163.367
R439 B.n391 B.n31 163.367
R440 B.n387 B.n31 163.367
R441 B.n387 B.n386 163.367
R442 B.n386 B.n385 163.367
R443 B.n385 B.n33 163.367
R444 B.n381 B.n33 163.367
R445 B.n381 B.n380 163.367
R446 B.n380 B.n379 163.367
R447 B.n379 B.n35 163.367
R448 B.n374 B.n35 163.367
R449 B.n374 B.n373 163.367
R450 B.n373 B.n372 163.367
R451 B.n372 B.n39 163.367
R452 B.n368 B.n39 163.367
R453 B.n368 B.n367 163.367
R454 B.n367 B.n366 163.367
R455 B.n366 B.n41 163.367
R456 B.n362 B.n41 163.367
R457 B.n362 B.n361 163.367
R458 B.n361 B.n360 163.367
R459 B.n360 B.n43 163.367
R460 B.n356 B.n43 163.367
R461 B.n356 B.n355 163.367
R462 B.n355 B.n354 163.367
R463 B.n354 B.n45 163.367
R464 B.n350 B.n45 163.367
R465 B.n350 B.n349 163.367
R466 B.n349 B.n348 163.367
R467 B.n348 B.n47 163.367
R468 B.n91 B.t4 115.207
R469 B.n37 B.t2 115.207
R470 B.n99 B.t10 115.203
R471 B.n29 B.t8 115.203
R472 B.n91 B.n90 78.9338
R473 B.n99 B.n98 78.9338
R474 B.n29 B.n28 78.9338
R475 B.n37 B.n36 78.9338
R476 B.n92 B.n91 59.5399
R477 B.n202 B.n99 59.5399
R478 B.n30 B.n29 59.5399
R479 B.n376 B.n37 59.5399
R480 B.n423 B.n18 34.8103
R481 B.n346 B.n345 34.8103
R482 B.n249 B.n80 34.8103
R483 B.n172 B.n171 34.8103
R484 B B.n471 18.0485
R485 B.n419 B.n18 10.6151
R486 B.n419 B.n418 10.6151
R487 B.n418 B.n417 10.6151
R488 B.n417 B.n20 10.6151
R489 B.n413 B.n20 10.6151
R490 B.n413 B.n412 10.6151
R491 B.n412 B.n411 10.6151
R492 B.n411 B.n22 10.6151
R493 B.n407 B.n22 10.6151
R494 B.n407 B.n406 10.6151
R495 B.n406 B.n405 10.6151
R496 B.n405 B.n24 10.6151
R497 B.n401 B.n24 10.6151
R498 B.n401 B.n400 10.6151
R499 B.n400 B.n399 10.6151
R500 B.n399 B.n26 10.6151
R501 B.n395 B.n26 10.6151
R502 B.n395 B.n394 10.6151
R503 B.n394 B.n393 10.6151
R504 B.n390 B.n389 10.6151
R505 B.n389 B.n388 10.6151
R506 B.n388 B.n32 10.6151
R507 B.n384 B.n32 10.6151
R508 B.n384 B.n383 10.6151
R509 B.n383 B.n382 10.6151
R510 B.n382 B.n34 10.6151
R511 B.n378 B.n34 10.6151
R512 B.n378 B.n377 10.6151
R513 B.n375 B.n38 10.6151
R514 B.n371 B.n38 10.6151
R515 B.n371 B.n370 10.6151
R516 B.n370 B.n369 10.6151
R517 B.n369 B.n40 10.6151
R518 B.n365 B.n40 10.6151
R519 B.n365 B.n364 10.6151
R520 B.n364 B.n363 10.6151
R521 B.n363 B.n42 10.6151
R522 B.n359 B.n42 10.6151
R523 B.n359 B.n358 10.6151
R524 B.n358 B.n357 10.6151
R525 B.n357 B.n44 10.6151
R526 B.n353 B.n44 10.6151
R527 B.n353 B.n352 10.6151
R528 B.n352 B.n351 10.6151
R529 B.n351 B.n46 10.6151
R530 B.n347 B.n46 10.6151
R531 B.n347 B.n346 10.6151
R532 B.n250 B.n249 10.6151
R533 B.n251 B.n250 10.6151
R534 B.n251 B.n78 10.6151
R535 B.n255 B.n78 10.6151
R536 B.n256 B.n255 10.6151
R537 B.n257 B.n256 10.6151
R538 B.n257 B.n76 10.6151
R539 B.n261 B.n76 10.6151
R540 B.n262 B.n261 10.6151
R541 B.n263 B.n262 10.6151
R542 B.n263 B.n74 10.6151
R543 B.n267 B.n74 10.6151
R544 B.n268 B.n267 10.6151
R545 B.n269 B.n268 10.6151
R546 B.n269 B.n72 10.6151
R547 B.n273 B.n72 10.6151
R548 B.n274 B.n273 10.6151
R549 B.n275 B.n274 10.6151
R550 B.n275 B.n70 10.6151
R551 B.n279 B.n70 10.6151
R552 B.n280 B.n279 10.6151
R553 B.n281 B.n280 10.6151
R554 B.n281 B.n68 10.6151
R555 B.n285 B.n68 10.6151
R556 B.n286 B.n285 10.6151
R557 B.n287 B.n286 10.6151
R558 B.n287 B.n66 10.6151
R559 B.n291 B.n66 10.6151
R560 B.n292 B.n291 10.6151
R561 B.n293 B.n292 10.6151
R562 B.n293 B.n64 10.6151
R563 B.n297 B.n64 10.6151
R564 B.n298 B.n297 10.6151
R565 B.n299 B.n298 10.6151
R566 B.n299 B.n62 10.6151
R567 B.n303 B.n62 10.6151
R568 B.n304 B.n303 10.6151
R569 B.n305 B.n304 10.6151
R570 B.n305 B.n60 10.6151
R571 B.n309 B.n60 10.6151
R572 B.n310 B.n309 10.6151
R573 B.n311 B.n310 10.6151
R574 B.n311 B.n58 10.6151
R575 B.n315 B.n58 10.6151
R576 B.n316 B.n315 10.6151
R577 B.n317 B.n316 10.6151
R578 B.n317 B.n56 10.6151
R579 B.n321 B.n56 10.6151
R580 B.n322 B.n321 10.6151
R581 B.n323 B.n322 10.6151
R582 B.n323 B.n54 10.6151
R583 B.n327 B.n54 10.6151
R584 B.n328 B.n327 10.6151
R585 B.n329 B.n328 10.6151
R586 B.n329 B.n52 10.6151
R587 B.n333 B.n52 10.6151
R588 B.n334 B.n333 10.6151
R589 B.n335 B.n334 10.6151
R590 B.n335 B.n50 10.6151
R591 B.n339 B.n50 10.6151
R592 B.n340 B.n339 10.6151
R593 B.n341 B.n340 10.6151
R594 B.n341 B.n48 10.6151
R595 B.n345 B.n48 10.6151
R596 B.n173 B.n172 10.6151
R597 B.n173 B.n108 10.6151
R598 B.n177 B.n108 10.6151
R599 B.n178 B.n177 10.6151
R600 B.n179 B.n178 10.6151
R601 B.n179 B.n106 10.6151
R602 B.n183 B.n106 10.6151
R603 B.n184 B.n183 10.6151
R604 B.n185 B.n184 10.6151
R605 B.n185 B.n104 10.6151
R606 B.n189 B.n104 10.6151
R607 B.n190 B.n189 10.6151
R608 B.n191 B.n190 10.6151
R609 B.n191 B.n102 10.6151
R610 B.n195 B.n102 10.6151
R611 B.n196 B.n195 10.6151
R612 B.n197 B.n196 10.6151
R613 B.n197 B.n100 10.6151
R614 B.n201 B.n100 10.6151
R615 B.n204 B.n203 10.6151
R616 B.n204 B.n96 10.6151
R617 B.n208 B.n96 10.6151
R618 B.n209 B.n208 10.6151
R619 B.n210 B.n209 10.6151
R620 B.n210 B.n94 10.6151
R621 B.n214 B.n94 10.6151
R622 B.n215 B.n214 10.6151
R623 B.n216 B.n215 10.6151
R624 B.n220 B.n219 10.6151
R625 B.n221 B.n220 10.6151
R626 B.n221 B.n88 10.6151
R627 B.n225 B.n88 10.6151
R628 B.n226 B.n225 10.6151
R629 B.n227 B.n226 10.6151
R630 B.n227 B.n86 10.6151
R631 B.n231 B.n86 10.6151
R632 B.n232 B.n231 10.6151
R633 B.n233 B.n232 10.6151
R634 B.n233 B.n84 10.6151
R635 B.n237 B.n84 10.6151
R636 B.n238 B.n237 10.6151
R637 B.n239 B.n238 10.6151
R638 B.n239 B.n82 10.6151
R639 B.n243 B.n82 10.6151
R640 B.n244 B.n243 10.6151
R641 B.n245 B.n244 10.6151
R642 B.n245 B.n80 10.6151
R643 B.n171 B.n110 10.6151
R644 B.n167 B.n110 10.6151
R645 B.n167 B.n166 10.6151
R646 B.n166 B.n165 10.6151
R647 B.n165 B.n112 10.6151
R648 B.n161 B.n112 10.6151
R649 B.n161 B.n160 10.6151
R650 B.n160 B.n159 10.6151
R651 B.n159 B.n114 10.6151
R652 B.n155 B.n114 10.6151
R653 B.n155 B.n154 10.6151
R654 B.n154 B.n153 10.6151
R655 B.n153 B.n116 10.6151
R656 B.n149 B.n116 10.6151
R657 B.n149 B.n148 10.6151
R658 B.n148 B.n147 10.6151
R659 B.n147 B.n118 10.6151
R660 B.n143 B.n118 10.6151
R661 B.n143 B.n142 10.6151
R662 B.n142 B.n141 10.6151
R663 B.n141 B.n120 10.6151
R664 B.n137 B.n120 10.6151
R665 B.n137 B.n136 10.6151
R666 B.n136 B.n135 10.6151
R667 B.n135 B.n122 10.6151
R668 B.n131 B.n122 10.6151
R669 B.n131 B.n130 10.6151
R670 B.n130 B.n129 10.6151
R671 B.n129 B.n124 10.6151
R672 B.n125 B.n124 10.6151
R673 B.n125 B.n0 10.6151
R674 B.n467 B.n1 10.6151
R675 B.n467 B.n466 10.6151
R676 B.n466 B.n465 10.6151
R677 B.n465 B.n4 10.6151
R678 B.n461 B.n4 10.6151
R679 B.n461 B.n460 10.6151
R680 B.n460 B.n459 10.6151
R681 B.n459 B.n6 10.6151
R682 B.n455 B.n6 10.6151
R683 B.n455 B.n454 10.6151
R684 B.n454 B.n453 10.6151
R685 B.n453 B.n8 10.6151
R686 B.n449 B.n8 10.6151
R687 B.n449 B.n448 10.6151
R688 B.n448 B.n447 10.6151
R689 B.n447 B.n10 10.6151
R690 B.n443 B.n10 10.6151
R691 B.n443 B.n442 10.6151
R692 B.n442 B.n441 10.6151
R693 B.n441 B.n12 10.6151
R694 B.n437 B.n12 10.6151
R695 B.n437 B.n436 10.6151
R696 B.n436 B.n435 10.6151
R697 B.n435 B.n14 10.6151
R698 B.n431 B.n14 10.6151
R699 B.n431 B.n430 10.6151
R700 B.n430 B.n429 10.6151
R701 B.n429 B.n16 10.6151
R702 B.n425 B.n16 10.6151
R703 B.n425 B.n424 10.6151
R704 B.n424 B.n423 10.6151
R705 B.n393 B.n30 9.36635
R706 B.n376 B.n375 9.36635
R707 B.n202 B.n201 9.36635
R708 B.n219 B.n92 9.36635
R709 B.n471 B.n0 2.81026
R710 B.n471 B.n1 2.81026
R711 B.n390 B.n30 1.24928
R712 B.n377 B.n376 1.24928
R713 B.n203 B.n202 1.24928
R714 B.n216 B.n92 1.24928
R715 VN VN.t1 107.915
R716 VN VN.t0 66.5144
R717 VTAIL.n1 VTAIL.t2 93.9032
R718 VTAIL.n2 VTAIL.t0 93.9023
R719 VTAIL.n3 VTAIL.t3 93.9023
R720 VTAIL.n0 VTAIL.t1 93.9023
R721 VTAIL.n1 VTAIL.n0 23.5048
R722 VTAIL.n3 VTAIL.n2 19.9962
R723 VTAIL.n2 VTAIL.n1 2.22464
R724 VTAIL VTAIL.n0 1.40567
R725 VTAIL VTAIL.n3 0.819465
R726 VDD2.n0 VDD2.t1 145.379
R727 VDD2.n0 VDD2.t0 110.582
R728 VDD2 VDD2.n0 0.935845
R729 VP.n0 VP.t0 108.103
R730 VP.n0 VP.t1 65.8937
R731 VP VP.n0 0.62124
R732 VDD1 VDD1.t0 146.78
R733 VDD1 VDD1.t1 111.516
C0 VN VP 4.65317f
C1 VDD2 VP 0.384934f
C2 VN VDD1 0.152832f
C3 VDD2 VDD1 0.799782f
C4 VN B 1.16126f
C5 VDD2 B 1.31322f
C6 VN w_n2598_n1924# 3.56383f
C7 VDD2 w_n2598_n1924# 1.45454f
C8 VTAIL VP 1.54521f
C9 VTAIL VDD1 3.4959f
C10 VTAIL B 2.31795f
C11 VP VDD1 1.54977f
C12 VP B 1.71387f
C13 VTAIL w_n2598_n1924# 1.79013f
C14 VP w_n2598_n1924# 3.89713f
C15 VN VDD2 1.31908f
C16 B VDD1 1.27276f
C17 w_n2598_n1924# VDD1 1.41492f
C18 w_n2598_n1924# B 8.03609f
C19 VTAIL VN 1.53091f
C20 VTAIL VDD2 3.55622f
C21 VDD2 VSUBS 0.735385f
C22 VDD1 VSUBS 3.156335f
C23 VTAIL VSUBS 0.537752f
C24 VN VSUBS 5.94073f
C25 VP VSUBS 1.614811f
C26 B VSUBS 3.919073f
C27 w_n2598_n1924# VSUBS 62.6949f
C28 VDD1.t1 VSUBS 0.501134f
C29 VDD1.t0 VSUBS 0.753862f
C30 VP.t0 VSUBS 2.95161f
C31 VP.t1 VSUBS 2.09738f
C32 VP.n0 VSUBS 3.40584f
C33 VDD2.t1 VSUBS 0.765977f
C34 VDD2.t0 VSUBS 0.521284f
C35 VDD2.n0 VSUBS 2.17318f
C36 VTAIL.t1 VSUBS 0.70708f
C37 VTAIL.n0 VSUBS 1.71489f
C38 VTAIL.t2 VSUBS 0.707083f
C39 VTAIL.n1 VSUBS 1.7779f
C40 VTAIL.t0 VSUBS 0.707078f
C41 VTAIL.n2 VSUBS 1.50794f
C42 VTAIL.t3 VSUBS 0.70708f
C43 VTAIL.n3 VSUBS 1.39982f
C44 VN.t0 VSUBS 2.01901f
C45 VN.t1 VSUBS 2.83098f
C46 B.n0 VSUBS 0.005178f
C47 B.n1 VSUBS 0.005178f
C48 B.n2 VSUBS 0.008189f
C49 B.n3 VSUBS 0.008189f
C50 B.n4 VSUBS 0.008189f
C51 B.n5 VSUBS 0.008189f
C52 B.n6 VSUBS 0.008189f
C53 B.n7 VSUBS 0.008189f
C54 B.n8 VSUBS 0.008189f
C55 B.n9 VSUBS 0.008189f
C56 B.n10 VSUBS 0.008189f
C57 B.n11 VSUBS 0.008189f
C58 B.n12 VSUBS 0.008189f
C59 B.n13 VSUBS 0.008189f
C60 B.n14 VSUBS 0.008189f
C61 B.n15 VSUBS 0.008189f
C62 B.n16 VSUBS 0.008189f
C63 B.n17 VSUBS 0.008189f
C64 B.n18 VSUBS 0.020333f
C65 B.n19 VSUBS 0.008189f
C66 B.n20 VSUBS 0.008189f
C67 B.n21 VSUBS 0.008189f
C68 B.n22 VSUBS 0.008189f
C69 B.n23 VSUBS 0.008189f
C70 B.n24 VSUBS 0.008189f
C71 B.n25 VSUBS 0.008189f
C72 B.n26 VSUBS 0.008189f
C73 B.n27 VSUBS 0.008189f
C74 B.t8 VSUBS 0.154583f
C75 B.t7 VSUBS 0.185221f
C76 B.t6 VSUBS 1.01254f
C77 B.n28 VSUBS 0.128174f
C78 B.n29 VSUBS 0.087033f
C79 B.n30 VSUBS 0.018972f
C80 B.n31 VSUBS 0.008189f
C81 B.n32 VSUBS 0.008189f
C82 B.n33 VSUBS 0.008189f
C83 B.n34 VSUBS 0.008189f
C84 B.n35 VSUBS 0.008189f
C85 B.t2 VSUBS 0.154583f
C86 B.t1 VSUBS 0.18522f
C87 B.t0 VSUBS 1.01254f
C88 B.n36 VSUBS 0.128175f
C89 B.n37 VSUBS 0.087033f
C90 B.n38 VSUBS 0.008189f
C91 B.n39 VSUBS 0.008189f
C92 B.n40 VSUBS 0.008189f
C93 B.n41 VSUBS 0.008189f
C94 B.n42 VSUBS 0.008189f
C95 B.n43 VSUBS 0.008189f
C96 B.n44 VSUBS 0.008189f
C97 B.n45 VSUBS 0.008189f
C98 B.n46 VSUBS 0.008189f
C99 B.n47 VSUBS 0.020333f
C100 B.n48 VSUBS 0.008189f
C101 B.n49 VSUBS 0.008189f
C102 B.n50 VSUBS 0.008189f
C103 B.n51 VSUBS 0.008189f
C104 B.n52 VSUBS 0.008189f
C105 B.n53 VSUBS 0.008189f
C106 B.n54 VSUBS 0.008189f
C107 B.n55 VSUBS 0.008189f
C108 B.n56 VSUBS 0.008189f
C109 B.n57 VSUBS 0.008189f
C110 B.n58 VSUBS 0.008189f
C111 B.n59 VSUBS 0.008189f
C112 B.n60 VSUBS 0.008189f
C113 B.n61 VSUBS 0.008189f
C114 B.n62 VSUBS 0.008189f
C115 B.n63 VSUBS 0.008189f
C116 B.n64 VSUBS 0.008189f
C117 B.n65 VSUBS 0.008189f
C118 B.n66 VSUBS 0.008189f
C119 B.n67 VSUBS 0.008189f
C120 B.n68 VSUBS 0.008189f
C121 B.n69 VSUBS 0.008189f
C122 B.n70 VSUBS 0.008189f
C123 B.n71 VSUBS 0.008189f
C124 B.n72 VSUBS 0.008189f
C125 B.n73 VSUBS 0.008189f
C126 B.n74 VSUBS 0.008189f
C127 B.n75 VSUBS 0.008189f
C128 B.n76 VSUBS 0.008189f
C129 B.n77 VSUBS 0.008189f
C130 B.n78 VSUBS 0.008189f
C131 B.n79 VSUBS 0.008189f
C132 B.n80 VSUBS 0.020333f
C133 B.n81 VSUBS 0.008189f
C134 B.n82 VSUBS 0.008189f
C135 B.n83 VSUBS 0.008189f
C136 B.n84 VSUBS 0.008189f
C137 B.n85 VSUBS 0.008189f
C138 B.n86 VSUBS 0.008189f
C139 B.n87 VSUBS 0.008189f
C140 B.n88 VSUBS 0.008189f
C141 B.n89 VSUBS 0.008189f
C142 B.t4 VSUBS 0.154583f
C143 B.t5 VSUBS 0.18522f
C144 B.t3 VSUBS 1.01254f
C145 B.n90 VSUBS 0.128175f
C146 B.n91 VSUBS 0.087033f
C147 B.n92 VSUBS 0.018972f
C148 B.n93 VSUBS 0.008189f
C149 B.n94 VSUBS 0.008189f
C150 B.n95 VSUBS 0.008189f
C151 B.n96 VSUBS 0.008189f
C152 B.n97 VSUBS 0.008189f
C153 B.t10 VSUBS 0.154583f
C154 B.t11 VSUBS 0.185221f
C155 B.t9 VSUBS 1.01254f
C156 B.n98 VSUBS 0.128174f
C157 B.n99 VSUBS 0.087033f
C158 B.n100 VSUBS 0.008189f
C159 B.n101 VSUBS 0.008189f
C160 B.n102 VSUBS 0.008189f
C161 B.n103 VSUBS 0.008189f
C162 B.n104 VSUBS 0.008189f
C163 B.n105 VSUBS 0.008189f
C164 B.n106 VSUBS 0.008189f
C165 B.n107 VSUBS 0.008189f
C166 B.n108 VSUBS 0.008189f
C167 B.n109 VSUBS 0.020333f
C168 B.n110 VSUBS 0.008189f
C169 B.n111 VSUBS 0.008189f
C170 B.n112 VSUBS 0.008189f
C171 B.n113 VSUBS 0.008189f
C172 B.n114 VSUBS 0.008189f
C173 B.n115 VSUBS 0.008189f
C174 B.n116 VSUBS 0.008189f
C175 B.n117 VSUBS 0.008189f
C176 B.n118 VSUBS 0.008189f
C177 B.n119 VSUBS 0.008189f
C178 B.n120 VSUBS 0.008189f
C179 B.n121 VSUBS 0.008189f
C180 B.n122 VSUBS 0.008189f
C181 B.n123 VSUBS 0.008189f
C182 B.n124 VSUBS 0.008189f
C183 B.n125 VSUBS 0.008189f
C184 B.n126 VSUBS 0.008189f
C185 B.n127 VSUBS 0.008189f
C186 B.n128 VSUBS 0.008189f
C187 B.n129 VSUBS 0.008189f
C188 B.n130 VSUBS 0.008189f
C189 B.n131 VSUBS 0.008189f
C190 B.n132 VSUBS 0.008189f
C191 B.n133 VSUBS 0.008189f
C192 B.n134 VSUBS 0.008189f
C193 B.n135 VSUBS 0.008189f
C194 B.n136 VSUBS 0.008189f
C195 B.n137 VSUBS 0.008189f
C196 B.n138 VSUBS 0.008189f
C197 B.n139 VSUBS 0.008189f
C198 B.n140 VSUBS 0.008189f
C199 B.n141 VSUBS 0.008189f
C200 B.n142 VSUBS 0.008189f
C201 B.n143 VSUBS 0.008189f
C202 B.n144 VSUBS 0.008189f
C203 B.n145 VSUBS 0.008189f
C204 B.n146 VSUBS 0.008189f
C205 B.n147 VSUBS 0.008189f
C206 B.n148 VSUBS 0.008189f
C207 B.n149 VSUBS 0.008189f
C208 B.n150 VSUBS 0.008189f
C209 B.n151 VSUBS 0.008189f
C210 B.n152 VSUBS 0.008189f
C211 B.n153 VSUBS 0.008189f
C212 B.n154 VSUBS 0.008189f
C213 B.n155 VSUBS 0.008189f
C214 B.n156 VSUBS 0.008189f
C215 B.n157 VSUBS 0.008189f
C216 B.n158 VSUBS 0.008189f
C217 B.n159 VSUBS 0.008189f
C218 B.n160 VSUBS 0.008189f
C219 B.n161 VSUBS 0.008189f
C220 B.n162 VSUBS 0.008189f
C221 B.n163 VSUBS 0.008189f
C222 B.n164 VSUBS 0.008189f
C223 B.n165 VSUBS 0.008189f
C224 B.n166 VSUBS 0.008189f
C225 B.n167 VSUBS 0.008189f
C226 B.n168 VSUBS 0.008189f
C227 B.n169 VSUBS 0.008189f
C228 B.n170 VSUBS 0.019647f
C229 B.n171 VSUBS 0.019647f
C230 B.n172 VSUBS 0.020333f
C231 B.n173 VSUBS 0.008189f
C232 B.n174 VSUBS 0.008189f
C233 B.n175 VSUBS 0.008189f
C234 B.n176 VSUBS 0.008189f
C235 B.n177 VSUBS 0.008189f
C236 B.n178 VSUBS 0.008189f
C237 B.n179 VSUBS 0.008189f
C238 B.n180 VSUBS 0.008189f
C239 B.n181 VSUBS 0.008189f
C240 B.n182 VSUBS 0.008189f
C241 B.n183 VSUBS 0.008189f
C242 B.n184 VSUBS 0.008189f
C243 B.n185 VSUBS 0.008189f
C244 B.n186 VSUBS 0.008189f
C245 B.n187 VSUBS 0.008189f
C246 B.n188 VSUBS 0.008189f
C247 B.n189 VSUBS 0.008189f
C248 B.n190 VSUBS 0.008189f
C249 B.n191 VSUBS 0.008189f
C250 B.n192 VSUBS 0.008189f
C251 B.n193 VSUBS 0.008189f
C252 B.n194 VSUBS 0.008189f
C253 B.n195 VSUBS 0.008189f
C254 B.n196 VSUBS 0.008189f
C255 B.n197 VSUBS 0.008189f
C256 B.n198 VSUBS 0.008189f
C257 B.n199 VSUBS 0.008189f
C258 B.n200 VSUBS 0.008189f
C259 B.n201 VSUBS 0.007707f
C260 B.n202 VSUBS 0.018972f
C261 B.n203 VSUBS 0.004576f
C262 B.n204 VSUBS 0.008189f
C263 B.n205 VSUBS 0.008189f
C264 B.n206 VSUBS 0.008189f
C265 B.n207 VSUBS 0.008189f
C266 B.n208 VSUBS 0.008189f
C267 B.n209 VSUBS 0.008189f
C268 B.n210 VSUBS 0.008189f
C269 B.n211 VSUBS 0.008189f
C270 B.n212 VSUBS 0.008189f
C271 B.n213 VSUBS 0.008189f
C272 B.n214 VSUBS 0.008189f
C273 B.n215 VSUBS 0.008189f
C274 B.n216 VSUBS 0.004576f
C275 B.n217 VSUBS 0.008189f
C276 B.n218 VSUBS 0.008189f
C277 B.n219 VSUBS 0.007707f
C278 B.n220 VSUBS 0.008189f
C279 B.n221 VSUBS 0.008189f
C280 B.n222 VSUBS 0.008189f
C281 B.n223 VSUBS 0.008189f
C282 B.n224 VSUBS 0.008189f
C283 B.n225 VSUBS 0.008189f
C284 B.n226 VSUBS 0.008189f
C285 B.n227 VSUBS 0.008189f
C286 B.n228 VSUBS 0.008189f
C287 B.n229 VSUBS 0.008189f
C288 B.n230 VSUBS 0.008189f
C289 B.n231 VSUBS 0.008189f
C290 B.n232 VSUBS 0.008189f
C291 B.n233 VSUBS 0.008189f
C292 B.n234 VSUBS 0.008189f
C293 B.n235 VSUBS 0.008189f
C294 B.n236 VSUBS 0.008189f
C295 B.n237 VSUBS 0.008189f
C296 B.n238 VSUBS 0.008189f
C297 B.n239 VSUBS 0.008189f
C298 B.n240 VSUBS 0.008189f
C299 B.n241 VSUBS 0.008189f
C300 B.n242 VSUBS 0.008189f
C301 B.n243 VSUBS 0.008189f
C302 B.n244 VSUBS 0.008189f
C303 B.n245 VSUBS 0.008189f
C304 B.n246 VSUBS 0.008189f
C305 B.n247 VSUBS 0.020333f
C306 B.n248 VSUBS 0.019647f
C307 B.n249 VSUBS 0.019647f
C308 B.n250 VSUBS 0.008189f
C309 B.n251 VSUBS 0.008189f
C310 B.n252 VSUBS 0.008189f
C311 B.n253 VSUBS 0.008189f
C312 B.n254 VSUBS 0.008189f
C313 B.n255 VSUBS 0.008189f
C314 B.n256 VSUBS 0.008189f
C315 B.n257 VSUBS 0.008189f
C316 B.n258 VSUBS 0.008189f
C317 B.n259 VSUBS 0.008189f
C318 B.n260 VSUBS 0.008189f
C319 B.n261 VSUBS 0.008189f
C320 B.n262 VSUBS 0.008189f
C321 B.n263 VSUBS 0.008189f
C322 B.n264 VSUBS 0.008189f
C323 B.n265 VSUBS 0.008189f
C324 B.n266 VSUBS 0.008189f
C325 B.n267 VSUBS 0.008189f
C326 B.n268 VSUBS 0.008189f
C327 B.n269 VSUBS 0.008189f
C328 B.n270 VSUBS 0.008189f
C329 B.n271 VSUBS 0.008189f
C330 B.n272 VSUBS 0.008189f
C331 B.n273 VSUBS 0.008189f
C332 B.n274 VSUBS 0.008189f
C333 B.n275 VSUBS 0.008189f
C334 B.n276 VSUBS 0.008189f
C335 B.n277 VSUBS 0.008189f
C336 B.n278 VSUBS 0.008189f
C337 B.n279 VSUBS 0.008189f
C338 B.n280 VSUBS 0.008189f
C339 B.n281 VSUBS 0.008189f
C340 B.n282 VSUBS 0.008189f
C341 B.n283 VSUBS 0.008189f
C342 B.n284 VSUBS 0.008189f
C343 B.n285 VSUBS 0.008189f
C344 B.n286 VSUBS 0.008189f
C345 B.n287 VSUBS 0.008189f
C346 B.n288 VSUBS 0.008189f
C347 B.n289 VSUBS 0.008189f
C348 B.n290 VSUBS 0.008189f
C349 B.n291 VSUBS 0.008189f
C350 B.n292 VSUBS 0.008189f
C351 B.n293 VSUBS 0.008189f
C352 B.n294 VSUBS 0.008189f
C353 B.n295 VSUBS 0.008189f
C354 B.n296 VSUBS 0.008189f
C355 B.n297 VSUBS 0.008189f
C356 B.n298 VSUBS 0.008189f
C357 B.n299 VSUBS 0.008189f
C358 B.n300 VSUBS 0.008189f
C359 B.n301 VSUBS 0.008189f
C360 B.n302 VSUBS 0.008189f
C361 B.n303 VSUBS 0.008189f
C362 B.n304 VSUBS 0.008189f
C363 B.n305 VSUBS 0.008189f
C364 B.n306 VSUBS 0.008189f
C365 B.n307 VSUBS 0.008189f
C366 B.n308 VSUBS 0.008189f
C367 B.n309 VSUBS 0.008189f
C368 B.n310 VSUBS 0.008189f
C369 B.n311 VSUBS 0.008189f
C370 B.n312 VSUBS 0.008189f
C371 B.n313 VSUBS 0.008189f
C372 B.n314 VSUBS 0.008189f
C373 B.n315 VSUBS 0.008189f
C374 B.n316 VSUBS 0.008189f
C375 B.n317 VSUBS 0.008189f
C376 B.n318 VSUBS 0.008189f
C377 B.n319 VSUBS 0.008189f
C378 B.n320 VSUBS 0.008189f
C379 B.n321 VSUBS 0.008189f
C380 B.n322 VSUBS 0.008189f
C381 B.n323 VSUBS 0.008189f
C382 B.n324 VSUBS 0.008189f
C383 B.n325 VSUBS 0.008189f
C384 B.n326 VSUBS 0.008189f
C385 B.n327 VSUBS 0.008189f
C386 B.n328 VSUBS 0.008189f
C387 B.n329 VSUBS 0.008189f
C388 B.n330 VSUBS 0.008189f
C389 B.n331 VSUBS 0.008189f
C390 B.n332 VSUBS 0.008189f
C391 B.n333 VSUBS 0.008189f
C392 B.n334 VSUBS 0.008189f
C393 B.n335 VSUBS 0.008189f
C394 B.n336 VSUBS 0.008189f
C395 B.n337 VSUBS 0.008189f
C396 B.n338 VSUBS 0.008189f
C397 B.n339 VSUBS 0.008189f
C398 B.n340 VSUBS 0.008189f
C399 B.n341 VSUBS 0.008189f
C400 B.n342 VSUBS 0.008189f
C401 B.n343 VSUBS 0.008189f
C402 B.n344 VSUBS 0.019647f
C403 B.n345 VSUBS 0.020555f
C404 B.n346 VSUBS 0.019425f
C405 B.n347 VSUBS 0.008189f
C406 B.n348 VSUBS 0.008189f
C407 B.n349 VSUBS 0.008189f
C408 B.n350 VSUBS 0.008189f
C409 B.n351 VSUBS 0.008189f
C410 B.n352 VSUBS 0.008189f
C411 B.n353 VSUBS 0.008189f
C412 B.n354 VSUBS 0.008189f
C413 B.n355 VSUBS 0.008189f
C414 B.n356 VSUBS 0.008189f
C415 B.n357 VSUBS 0.008189f
C416 B.n358 VSUBS 0.008189f
C417 B.n359 VSUBS 0.008189f
C418 B.n360 VSUBS 0.008189f
C419 B.n361 VSUBS 0.008189f
C420 B.n362 VSUBS 0.008189f
C421 B.n363 VSUBS 0.008189f
C422 B.n364 VSUBS 0.008189f
C423 B.n365 VSUBS 0.008189f
C424 B.n366 VSUBS 0.008189f
C425 B.n367 VSUBS 0.008189f
C426 B.n368 VSUBS 0.008189f
C427 B.n369 VSUBS 0.008189f
C428 B.n370 VSUBS 0.008189f
C429 B.n371 VSUBS 0.008189f
C430 B.n372 VSUBS 0.008189f
C431 B.n373 VSUBS 0.008189f
C432 B.n374 VSUBS 0.008189f
C433 B.n375 VSUBS 0.007707f
C434 B.n376 VSUBS 0.018972f
C435 B.n377 VSUBS 0.004576f
C436 B.n378 VSUBS 0.008189f
C437 B.n379 VSUBS 0.008189f
C438 B.n380 VSUBS 0.008189f
C439 B.n381 VSUBS 0.008189f
C440 B.n382 VSUBS 0.008189f
C441 B.n383 VSUBS 0.008189f
C442 B.n384 VSUBS 0.008189f
C443 B.n385 VSUBS 0.008189f
C444 B.n386 VSUBS 0.008189f
C445 B.n387 VSUBS 0.008189f
C446 B.n388 VSUBS 0.008189f
C447 B.n389 VSUBS 0.008189f
C448 B.n390 VSUBS 0.004576f
C449 B.n391 VSUBS 0.008189f
C450 B.n392 VSUBS 0.008189f
C451 B.n393 VSUBS 0.007707f
C452 B.n394 VSUBS 0.008189f
C453 B.n395 VSUBS 0.008189f
C454 B.n396 VSUBS 0.008189f
C455 B.n397 VSUBS 0.008189f
C456 B.n398 VSUBS 0.008189f
C457 B.n399 VSUBS 0.008189f
C458 B.n400 VSUBS 0.008189f
C459 B.n401 VSUBS 0.008189f
C460 B.n402 VSUBS 0.008189f
C461 B.n403 VSUBS 0.008189f
C462 B.n404 VSUBS 0.008189f
C463 B.n405 VSUBS 0.008189f
C464 B.n406 VSUBS 0.008189f
C465 B.n407 VSUBS 0.008189f
C466 B.n408 VSUBS 0.008189f
C467 B.n409 VSUBS 0.008189f
C468 B.n410 VSUBS 0.008189f
C469 B.n411 VSUBS 0.008189f
C470 B.n412 VSUBS 0.008189f
C471 B.n413 VSUBS 0.008189f
C472 B.n414 VSUBS 0.008189f
C473 B.n415 VSUBS 0.008189f
C474 B.n416 VSUBS 0.008189f
C475 B.n417 VSUBS 0.008189f
C476 B.n418 VSUBS 0.008189f
C477 B.n419 VSUBS 0.008189f
C478 B.n420 VSUBS 0.008189f
C479 B.n421 VSUBS 0.020333f
C480 B.n422 VSUBS 0.019647f
C481 B.n423 VSUBS 0.019647f
C482 B.n424 VSUBS 0.008189f
C483 B.n425 VSUBS 0.008189f
C484 B.n426 VSUBS 0.008189f
C485 B.n427 VSUBS 0.008189f
C486 B.n428 VSUBS 0.008189f
C487 B.n429 VSUBS 0.008189f
C488 B.n430 VSUBS 0.008189f
C489 B.n431 VSUBS 0.008189f
C490 B.n432 VSUBS 0.008189f
C491 B.n433 VSUBS 0.008189f
C492 B.n434 VSUBS 0.008189f
C493 B.n435 VSUBS 0.008189f
C494 B.n436 VSUBS 0.008189f
C495 B.n437 VSUBS 0.008189f
C496 B.n438 VSUBS 0.008189f
C497 B.n439 VSUBS 0.008189f
C498 B.n440 VSUBS 0.008189f
C499 B.n441 VSUBS 0.008189f
C500 B.n442 VSUBS 0.008189f
C501 B.n443 VSUBS 0.008189f
C502 B.n444 VSUBS 0.008189f
C503 B.n445 VSUBS 0.008189f
C504 B.n446 VSUBS 0.008189f
C505 B.n447 VSUBS 0.008189f
C506 B.n448 VSUBS 0.008189f
C507 B.n449 VSUBS 0.008189f
C508 B.n450 VSUBS 0.008189f
C509 B.n451 VSUBS 0.008189f
C510 B.n452 VSUBS 0.008189f
C511 B.n453 VSUBS 0.008189f
C512 B.n454 VSUBS 0.008189f
C513 B.n455 VSUBS 0.008189f
C514 B.n456 VSUBS 0.008189f
C515 B.n457 VSUBS 0.008189f
C516 B.n458 VSUBS 0.008189f
C517 B.n459 VSUBS 0.008189f
C518 B.n460 VSUBS 0.008189f
C519 B.n461 VSUBS 0.008189f
C520 B.n462 VSUBS 0.008189f
C521 B.n463 VSUBS 0.008189f
C522 B.n464 VSUBS 0.008189f
C523 B.n465 VSUBS 0.008189f
C524 B.n466 VSUBS 0.008189f
C525 B.n467 VSUBS 0.008189f
C526 B.n468 VSUBS 0.008189f
C527 B.n469 VSUBS 0.008189f
C528 B.n470 VSUBS 0.008189f
C529 B.n471 VSUBS 0.018542f
.ends

