* NGSPICE file created from diff_pair_sample_0452.ext - technology: sky130A

.subckt diff_pair_sample_0452 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=2.29185 ps=14.22 w=13.89 l=3.11
X1 VTAIL.t4 VP.t0 VDD1.t5 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=2.29185 ps=14.22 w=13.89 l=3.11
X2 VDD2.t4 VN.t1 VTAIL.t11 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=2.29185 ps=14.22 w=13.89 l=3.11
X3 VTAIL.t10 VN.t2 VDD2.t3 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=2.29185 ps=14.22 w=13.89 l=3.11
X4 B.t11 B.t9 B.t10 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=0 ps=0 w=13.89 l=3.11
X5 VTAIL.t8 VN.t3 VDD2.t2 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=2.29185 ps=14.22 w=13.89 l=3.11
X6 VDD1.t4 VP.t1 VTAIL.t5 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=2.29185 ps=14.22 w=13.89 l=3.11
X7 VDD2.t1 VN.t4 VTAIL.t7 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=5.4171 ps=28.56 w=13.89 l=3.11
X8 VDD1.t3 VP.t2 VTAIL.t0 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=5.4171 ps=28.56 w=13.89 l=3.11
X9 VDD2.t0 VN.t5 VTAIL.t6 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=5.4171 ps=28.56 w=13.89 l=3.11
X10 B.t8 B.t6 B.t7 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=0 ps=0 w=13.89 l=3.11
X11 VTAIL.t3 VP.t3 VDD1.t2 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=2.29185 ps=14.22 w=13.89 l=3.11
X12 VDD1.t1 VP.t4 VTAIL.t1 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=2.29185 pd=14.22 as=5.4171 ps=28.56 w=13.89 l=3.11
X13 B.t5 B.t3 B.t4 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=0 ps=0 w=13.89 l=3.11
X14 VDD1.t0 VP.t5 VTAIL.t2 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=2.29185 ps=14.22 w=13.89 l=3.11
X15 B.t2 B.t0 B.t1 w_n3722_n3746# sky130_fd_pr__pfet_01v8 ad=5.4171 pd=28.56 as=0 ps=0 w=13.89 l=3.11
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t4 141.054
R13 VN.n4 VN.t0 141.054
R14 VN.n5 VN.t3 107.636
R15 VN.n0 VN.t5 107.636
R16 VN.n21 VN.t2 107.636
R17 VN.n16 VN.t1 107.636
R18 VN.n15 VN.n0 68.5364
R19 VN.n31 VN.n16 68.5364
R20 VN.n11 VN.n2 56.5193
R21 VN.n27 VN.n18 56.5193
R22 VN VN.n31 52.445
R23 VN.n5 VN.n4 49.4728
R24 VN.n21 VN.n20 49.4728
R25 VN.n6 VN.n5 24.4675
R26 VN.n7 VN.n6 24.4675
R27 VN.n7 VN.n2 24.4675
R28 VN.n12 VN.n11 24.4675
R29 VN.n13 VN.n12 24.4675
R30 VN.n23 VN.n18 24.4675
R31 VN.n23 VN.n22 24.4675
R32 VN.n22 VN.n21 24.4675
R33 VN.n29 VN.n28 24.4675
R34 VN.n28 VN.n27 24.4675
R35 VN.n13 VN.n0 21.5315
R36 VN.n29 VN.n16 21.5315
R37 VN.n20 VN.n19 3.84099
R38 VN.n4 VN.n3 3.84099
R39 VN.n31 VN.n30 0.354971
R40 VN.n15 VN.n14 0.354971
R41 VN VN.n15 0.26696
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n10 VTAIL.t1 57.0267
R53 VTAIL.n7 VTAIL.t7 57.0267
R54 VTAIL.n11 VTAIL.t6 57.0265
R55 VTAIL.n2 VTAIL.t0 57.0265
R56 VTAIL.n9 VTAIL.n8 54.6866
R57 VTAIL.n6 VTAIL.n5 54.6866
R58 VTAIL.n1 VTAIL.n0 54.6865
R59 VTAIL.n4 VTAIL.n3 54.6865
R60 VTAIL.n6 VTAIL.n4 30.2721
R61 VTAIL.n11 VTAIL.n10 27.3065
R62 VTAIL.n7 VTAIL.n6 2.96602
R63 VTAIL.n10 VTAIL.n9 2.96602
R64 VTAIL.n4 VTAIL.n2 2.96602
R65 VTAIL.n0 VTAIL.t9 2.34067
R66 VTAIL.n0 VTAIL.t8 2.34067
R67 VTAIL.n3 VTAIL.t2 2.34067
R68 VTAIL.n3 VTAIL.t3 2.34067
R69 VTAIL.n8 VTAIL.t5 2.34067
R70 VTAIL.n8 VTAIL.t4 2.34067
R71 VTAIL.n5 VTAIL.t11 2.34067
R72 VTAIL.n5 VTAIL.t10 2.34067
R73 VTAIL VTAIL.n11 2.16645
R74 VTAIL.n9 VTAIL.n7 1.95309
R75 VTAIL.n2 VTAIL.n1 1.95309
R76 VTAIL VTAIL.n1 0.800069
R77 VDD2.n1 VDD2.t5 75.8741
R78 VDD2.n2 VDD2.t4 73.7055
R79 VDD2.n1 VDD2.n0 72.0513
R80 VDD2 VDD2.n3 72.0485
R81 VDD2.n2 VDD2.n1 45.3274
R82 VDD2.n3 VDD2.t3 2.34067
R83 VDD2.n3 VDD2.t1 2.34067
R84 VDD2.n0 VDD2.t2 2.34067
R85 VDD2.n0 VDD2.t0 2.34067
R86 VDD2 VDD2.n2 2.28283
R87 VP.n13 VP.n10 161.3
R88 VP.n15 VP.n14 161.3
R89 VP.n16 VP.n9 161.3
R90 VP.n18 VP.n17 161.3
R91 VP.n19 VP.n8 161.3
R92 VP.n21 VP.n20 161.3
R93 VP.n44 VP.n43 161.3
R94 VP.n42 VP.n1 161.3
R95 VP.n41 VP.n40 161.3
R96 VP.n39 VP.n2 161.3
R97 VP.n38 VP.n37 161.3
R98 VP.n36 VP.n3 161.3
R99 VP.n35 VP.n34 161.3
R100 VP.n33 VP.n4 161.3
R101 VP.n32 VP.n31 161.3
R102 VP.n30 VP.n5 161.3
R103 VP.n29 VP.n28 161.3
R104 VP.n27 VP.n6 161.3
R105 VP.n26 VP.n25 161.3
R106 VP.n11 VP.t1 141.054
R107 VP.n35 VP.t3 107.636
R108 VP.n24 VP.t5 107.636
R109 VP.n0 VP.t2 107.636
R110 VP.n12 VP.t0 107.636
R111 VP.n7 VP.t4 107.636
R112 VP.n24 VP.n23 68.5364
R113 VP.n45 VP.n0 68.5364
R114 VP.n22 VP.n7 68.5364
R115 VP.n30 VP.n29 56.5193
R116 VP.n41 VP.n2 56.5193
R117 VP.n18 VP.n9 56.5193
R118 VP.n23 VP.n22 52.2796
R119 VP.n12 VP.n11 49.4728
R120 VP.n25 VP.n6 24.4675
R121 VP.n29 VP.n6 24.4675
R122 VP.n31 VP.n30 24.4675
R123 VP.n31 VP.n4 24.4675
R124 VP.n35 VP.n4 24.4675
R125 VP.n36 VP.n35 24.4675
R126 VP.n37 VP.n36 24.4675
R127 VP.n37 VP.n2 24.4675
R128 VP.n42 VP.n41 24.4675
R129 VP.n43 VP.n42 24.4675
R130 VP.n19 VP.n18 24.4675
R131 VP.n20 VP.n19 24.4675
R132 VP.n13 VP.n12 24.4675
R133 VP.n14 VP.n13 24.4675
R134 VP.n14 VP.n9 24.4675
R135 VP.n25 VP.n24 21.5315
R136 VP.n43 VP.n0 21.5315
R137 VP.n20 VP.n7 21.5315
R138 VP.n11 VP.n10 3.84097
R139 VP.n22 VP.n21 0.354971
R140 VP.n26 VP.n23 0.354971
R141 VP.n45 VP.n44 0.354971
R142 VP VP.n45 0.26696
R143 VP.n15 VP.n10 0.189894
R144 VP.n16 VP.n15 0.189894
R145 VP.n17 VP.n16 0.189894
R146 VP.n17 VP.n8 0.189894
R147 VP.n21 VP.n8 0.189894
R148 VP.n27 VP.n26 0.189894
R149 VP.n28 VP.n27 0.189894
R150 VP.n28 VP.n5 0.189894
R151 VP.n32 VP.n5 0.189894
R152 VP.n33 VP.n32 0.189894
R153 VP.n34 VP.n33 0.189894
R154 VP.n34 VP.n3 0.189894
R155 VP.n38 VP.n3 0.189894
R156 VP.n39 VP.n38 0.189894
R157 VP.n40 VP.n39 0.189894
R158 VP.n40 VP.n1 0.189894
R159 VP.n44 VP.n1 0.189894
R160 VDD1 VDD1.t4 75.9878
R161 VDD1.n1 VDD1.t0 75.8741
R162 VDD1.n1 VDD1.n0 72.0513
R163 VDD1.n3 VDD1.n2 71.3653
R164 VDD1.n3 VDD1.n1 47.3931
R165 VDD1.n2 VDD1.t5 2.34067
R166 VDD1.n2 VDD1.t1 2.34067
R167 VDD1.n0 VDD1.t2 2.34067
R168 VDD1.n0 VDD1.t3 2.34067
R169 VDD1 VDD1.n3 0.68369
R170 B.n439 B.n132 585
R171 B.n438 B.n437 585
R172 B.n436 B.n133 585
R173 B.n435 B.n434 585
R174 B.n433 B.n134 585
R175 B.n432 B.n431 585
R176 B.n430 B.n135 585
R177 B.n429 B.n428 585
R178 B.n427 B.n136 585
R179 B.n426 B.n425 585
R180 B.n424 B.n137 585
R181 B.n423 B.n422 585
R182 B.n421 B.n138 585
R183 B.n420 B.n419 585
R184 B.n418 B.n139 585
R185 B.n417 B.n416 585
R186 B.n415 B.n140 585
R187 B.n414 B.n413 585
R188 B.n412 B.n141 585
R189 B.n411 B.n410 585
R190 B.n409 B.n142 585
R191 B.n408 B.n407 585
R192 B.n406 B.n143 585
R193 B.n405 B.n404 585
R194 B.n403 B.n144 585
R195 B.n402 B.n401 585
R196 B.n400 B.n145 585
R197 B.n399 B.n398 585
R198 B.n397 B.n146 585
R199 B.n396 B.n395 585
R200 B.n394 B.n147 585
R201 B.n393 B.n392 585
R202 B.n391 B.n148 585
R203 B.n390 B.n389 585
R204 B.n388 B.n149 585
R205 B.n387 B.n386 585
R206 B.n385 B.n150 585
R207 B.n384 B.n383 585
R208 B.n382 B.n151 585
R209 B.n381 B.n380 585
R210 B.n379 B.n152 585
R211 B.n378 B.n377 585
R212 B.n376 B.n153 585
R213 B.n375 B.n374 585
R214 B.n373 B.n154 585
R215 B.n372 B.n371 585
R216 B.n370 B.n155 585
R217 B.n369 B.n368 585
R218 B.n364 B.n156 585
R219 B.n363 B.n362 585
R220 B.n361 B.n157 585
R221 B.n360 B.n359 585
R222 B.n358 B.n158 585
R223 B.n357 B.n356 585
R224 B.n355 B.n159 585
R225 B.n354 B.n353 585
R226 B.n352 B.n160 585
R227 B.n350 B.n349 585
R228 B.n348 B.n163 585
R229 B.n347 B.n346 585
R230 B.n345 B.n164 585
R231 B.n344 B.n343 585
R232 B.n342 B.n165 585
R233 B.n341 B.n340 585
R234 B.n339 B.n166 585
R235 B.n338 B.n337 585
R236 B.n336 B.n167 585
R237 B.n335 B.n334 585
R238 B.n333 B.n168 585
R239 B.n332 B.n331 585
R240 B.n330 B.n169 585
R241 B.n329 B.n328 585
R242 B.n327 B.n170 585
R243 B.n326 B.n325 585
R244 B.n324 B.n171 585
R245 B.n323 B.n322 585
R246 B.n321 B.n172 585
R247 B.n320 B.n319 585
R248 B.n318 B.n173 585
R249 B.n317 B.n316 585
R250 B.n315 B.n174 585
R251 B.n314 B.n313 585
R252 B.n312 B.n175 585
R253 B.n311 B.n310 585
R254 B.n309 B.n176 585
R255 B.n308 B.n307 585
R256 B.n306 B.n177 585
R257 B.n305 B.n304 585
R258 B.n303 B.n178 585
R259 B.n302 B.n301 585
R260 B.n300 B.n179 585
R261 B.n299 B.n298 585
R262 B.n297 B.n180 585
R263 B.n296 B.n295 585
R264 B.n294 B.n181 585
R265 B.n293 B.n292 585
R266 B.n291 B.n182 585
R267 B.n290 B.n289 585
R268 B.n288 B.n183 585
R269 B.n287 B.n286 585
R270 B.n285 B.n184 585
R271 B.n284 B.n283 585
R272 B.n282 B.n185 585
R273 B.n281 B.n280 585
R274 B.n441 B.n440 585
R275 B.n442 B.n131 585
R276 B.n444 B.n443 585
R277 B.n445 B.n130 585
R278 B.n447 B.n446 585
R279 B.n448 B.n129 585
R280 B.n450 B.n449 585
R281 B.n451 B.n128 585
R282 B.n453 B.n452 585
R283 B.n454 B.n127 585
R284 B.n456 B.n455 585
R285 B.n457 B.n126 585
R286 B.n459 B.n458 585
R287 B.n460 B.n125 585
R288 B.n462 B.n461 585
R289 B.n463 B.n124 585
R290 B.n465 B.n464 585
R291 B.n466 B.n123 585
R292 B.n468 B.n467 585
R293 B.n469 B.n122 585
R294 B.n471 B.n470 585
R295 B.n472 B.n121 585
R296 B.n474 B.n473 585
R297 B.n475 B.n120 585
R298 B.n477 B.n476 585
R299 B.n478 B.n119 585
R300 B.n480 B.n479 585
R301 B.n481 B.n118 585
R302 B.n483 B.n482 585
R303 B.n484 B.n117 585
R304 B.n486 B.n485 585
R305 B.n487 B.n116 585
R306 B.n489 B.n488 585
R307 B.n490 B.n115 585
R308 B.n492 B.n491 585
R309 B.n493 B.n114 585
R310 B.n495 B.n494 585
R311 B.n496 B.n113 585
R312 B.n498 B.n497 585
R313 B.n499 B.n112 585
R314 B.n501 B.n500 585
R315 B.n502 B.n111 585
R316 B.n504 B.n503 585
R317 B.n505 B.n110 585
R318 B.n507 B.n506 585
R319 B.n508 B.n109 585
R320 B.n510 B.n509 585
R321 B.n511 B.n108 585
R322 B.n513 B.n512 585
R323 B.n514 B.n107 585
R324 B.n516 B.n515 585
R325 B.n517 B.n106 585
R326 B.n519 B.n518 585
R327 B.n520 B.n105 585
R328 B.n522 B.n521 585
R329 B.n523 B.n104 585
R330 B.n525 B.n524 585
R331 B.n526 B.n103 585
R332 B.n528 B.n527 585
R333 B.n529 B.n102 585
R334 B.n531 B.n530 585
R335 B.n532 B.n101 585
R336 B.n534 B.n533 585
R337 B.n535 B.n100 585
R338 B.n537 B.n536 585
R339 B.n538 B.n99 585
R340 B.n540 B.n539 585
R341 B.n541 B.n98 585
R342 B.n543 B.n542 585
R343 B.n544 B.n97 585
R344 B.n546 B.n545 585
R345 B.n547 B.n96 585
R346 B.n549 B.n548 585
R347 B.n550 B.n95 585
R348 B.n552 B.n551 585
R349 B.n553 B.n94 585
R350 B.n555 B.n554 585
R351 B.n556 B.n93 585
R352 B.n558 B.n557 585
R353 B.n559 B.n92 585
R354 B.n561 B.n560 585
R355 B.n562 B.n91 585
R356 B.n564 B.n563 585
R357 B.n565 B.n90 585
R358 B.n567 B.n566 585
R359 B.n568 B.n89 585
R360 B.n570 B.n569 585
R361 B.n571 B.n88 585
R362 B.n573 B.n572 585
R363 B.n574 B.n87 585
R364 B.n576 B.n575 585
R365 B.n577 B.n86 585
R366 B.n579 B.n578 585
R367 B.n580 B.n85 585
R368 B.n582 B.n581 585
R369 B.n583 B.n84 585
R370 B.n585 B.n584 585
R371 B.n586 B.n83 585
R372 B.n743 B.n26 585
R373 B.n742 B.n741 585
R374 B.n740 B.n27 585
R375 B.n739 B.n738 585
R376 B.n737 B.n28 585
R377 B.n736 B.n735 585
R378 B.n734 B.n29 585
R379 B.n733 B.n732 585
R380 B.n731 B.n30 585
R381 B.n730 B.n729 585
R382 B.n728 B.n31 585
R383 B.n727 B.n726 585
R384 B.n725 B.n32 585
R385 B.n724 B.n723 585
R386 B.n722 B.n33 585
R387 B.n721 B.n720 585
R388 B.n719 B.n34 585
R389 B.n718 B.n717 585
R390 B.n716 B.n35 585
R391 B.n715 B.n714 585
R392 B.n713 B.n36 585
R393 B.n712 B.n711 585
R394 B.n710 B.n37 585
R395 B.n709 B.n708 585
R396 B.n707 B.n38 585
R397 B.n706 B.n705 585
R398 B.n704 B.n39 585
R399 B.n703 B.n702 585
R400 B.n701 B.n40 585
R401 B.n700 B.n699 585
R402 B.n698 B.n41 585
R403 B.n697 B.n696 585
R404 B.n695 B.n42 585
R405 B.n694 B.n693 585
R406 B.n692 B.n43 585
R407 B.n691 B.n690 585
R408 B.n689 B.n44 585
R409 B.n688 B.n687 585
R410 B.n686 B.n45 585
R411 B.n685 B.n684 585
R412 B.n683 B.n46 585
R413 B.n682 B.n681 585
R414 B.n680 B.n47 585
R415 B.n679 B.n678 585
R416 B.n677 B.n48 585
R417 B.n676 B.n675 585
R418 B.n674 B.n49 585
R419 B.n672 B.n671 585
R420 B.n670 B.n52 585
R421 B.n669 B.n668 585
R422 B.n667 B.n53 585
R423 B.n666 B.n665 585
R424 B.n664 B.n54 585
R425 B.n663 B.n662 585
R426 B.n661 B.n55 585
R427 B.n660 B.n659 585
R428 B.n658 B.n56 585
R429 B.n657 B.n656 585
R430 B.n655 B.n57 585
R431 B.n654 B.n653 585
R432 B.n652 B.n61 585
R433 B.n651 B.n650 585
R434 B.n649 B.n62 585
R435 B.n648 B.n647 585
R436 B.n646 B.n63 585
R437 B.n645 B.n644 585
R438 B.n643 B.n64 585
R439 B.n642 B.n641 585
R440 B.n640 B.n65 585
R441 B.n639 B.n638 585
R442 B.n637 B.n66 585
R443 B.n636 B.n635 585
R444 B.n634 B.n67 585
R445 B.n633 B.n632 585
R446 B.n631 B.n68 585
R447 B.n630 B.n629 585
R448 B.n628 B.n69 585
R449 B.n627 B.n626 585
R450 B.n625 B.n70 585
R451 B.n624 B.n623 585
R452 B.n622 B.n71 585
R453 B.n621 B.n620 585
R454 B.n619 B.n72 585
R455 B.n618 B.n617 585
R456 B.n616 B.n73 585
R457 B.n615 B.n614 585
R458 B.n613 B.n74 585
R459 B.n612 B.n611 585
R460 B.n610 B.n75 585
R461 B.n609 B.n608 585
R462 B.n607 B.n76 585
R463 B.n606 B.n605 585
R464 B.n604 B.n77 585
R465 B.n603 B.n602 585
R466 B.n601 B.n78 585
R467 B.n600 B.n599 585
R468 B.n598 B.n79 585
R469 B.n597 B.n596 585
R470 B.n595 B.n80 585
R471 B.n594 B.n593 585
R472 B.n592 B.n81 585
R473 B.n591 B.n590 585
R474 B.n589 B.n82 585
R475 B.n588 B.n587 585
R476 B.n745 B.n744 585
R477 B.n746 B.n25 585
R478 B.n748 B.n747 585
R479 B.n749 B.n24 585
R480 B.n751 B.n750 585
R481 B.n752 B.n23 585
R482 B.n754 B.n753 585
R483 B.n755 B.n22 585
R484 B.n757 B.n756 585
R485 B.n758 B.n21 585
R486 B.n760 B.n759 585
R487 B.n761 B.n20 585
R488 B.n763 B.n762 585
R489 B.n764 B.n19 585
R490 B.n766 B.n765 585
R491 B.n767 B.n18 585
R492 B.n769 B.n768 585
R493 B.n770 B.n17 585
R494 B.n772 B.n771 585
R495 B.n773 B.n16 585
R496 B.n775 B.n774 585
R497 B.n776 B.n15 585
R498 B.n778 B.n777 585
R499 B.n779 B.n14 585
R500 B.n781 B.n780 585
R501 B.n782 B.n13 585
R502 B.n784 B.n783 585
R503 B.n785 B.n12 585
R504 B.n787 B.n786 585
R505 B.n788 B.n11 585
R506 B.n790 B.n789 585
R507 B.n791 B.n10 585
R508 B.n793 B.n792 585
R509 B.n794 B.n9 585
R510 B.n796 B.n795 585
R511 B.n797 B.n8 585
R512 B.n799 B.n798 585
R513 B.n800 B.n7 585
R514 B.n802 B.n801 585
R515 B.n803 B.n6 585
R516 B.n805 B.n804 585
R517 B.n806 B.n5 585
R518 B.n808 B.n807 585
R519 B.n809 B.n4 585
R520 B.n811 B.n810 585
R521 B.n812 B.n3 585
R522 B.n814 B.n813 585
R523 B.n815 B.n0 585
R524 B.n2 B.n1 585
R525 B.n210 B.n209 585
R526 B.n212 B.n211 585
R527 B.n213 B.n208 585
R528 B.n215 B.n214 585
R529 B.n216 B.n207 585
R530 B.n218 B.n217 585
R531 B.n219 B.n206 585
R532 B.n221 B.n220 585
R533 B.n222 B.n205 585
R534 B.n224 B.n223 585
R535 B.n225 B.n204 585
R536 B.n227 B.n226 585
R537 B.n228 B.n203 585
R538 B.n230 B.n229 585
R539 B.n231 B.n202 585
R540 B.n233 B.n232 585
R541 B.n234 B.n201 585
R542 B.n236 B.n235 585
R543 B.n237 B.n200 585
R544 B.n239 B.n238 585
R545 B.n240 B.n199 585
R546 B.n242 B.n241 585
R547 B.n243 B.n198 585
R548 B.n245 B.n244 585
R549 B.n246 B.n197 585
R550 B.n248 B.n247 585
R551 B.n249 B.n196 585
R552 B.n251 B.n250 585
R553 B.n252 B.n195 585
R554 B.n254 B.n253 585
R555 B.n255 B.n194 585
R556 B.n257 B.n256 585
R557 B.n258 B.n193 585
R558 B.n260 B.n259 585
R559 B.n261 B.n192 585
R560 B.n263 B.n262 585
R561 B.n264 B.n191 585
R562 B.n266 B.n265 585
R563 B.n267 B.n190 585
R564 B.n269 B.n268 585
R565 B.n270 B.n189 585
R566 B.n272 B.n271 585
R567 B.n273 B.n188 585
R568 B.n275 B.n274 585
R569 B.n276 B.n187 585
R570 B.n278 B.n277 585
R571 B.n279 B.n186 585
R572 B.n281 B.n186 506.916
R573 B.n441 B.n132 506.916
R574 B.n587 B.n586 506.916
R575 B.n744 B.n743 506.916
R576 B.n161 B.t3 316.342
R577 B.n365 B.t6 316.342
R578 B.n58 B.t0 316.342
R579 B.n50 B.t9 316.342
R580 B.n817 B.n816 256.663
R581 B.n816 B.n815 235.042
R582 B.n816 B.n2 235.042
R583 B.n365 B.t7 179.072
R584 B.n58 B.t2 179.072
R585 B.n161 B.t4 179.055
R586 B.n50 B.t11 179.055
R587 B.n282 B.n281 163.367
R588 B.n283 B.n282 163.367
R589 B.n283 B.n184 163.367
R590 B.n287 B.n184 163.367
R591 B.n288 B.n287 163.367
R592 B.n289 B.n288 163.367
R593 B.n289 B.n182 163.367
R594 B.n293 B.n182 163.367
R595 B.n294 B.n293 163.367
R596 B.n295 B.n294 163.367
R597 B.n295 B.n180 163.367
R598 B.n299 B.n180 163.367
R599 B.n300 B.n299 163.367
R600 B.n301 B.n300 163.367
R601 B.n301 B.n178 163.367
R602 B.n305 B.n178 163.367
R603 B.n306 B.n305 163.367
R604 B.n307 B.n306 163.367
R605 B.n307 B.n176 163.367
R606 B.n311 B.n176 163.367
R607 B.n312 B.n311 163.367
R608 B.n313 B.n312 163.367
R609 B.n313 B.n174 163.367
R610 B.n317 B.n174 163.367
R611 B.n318 B.n317 163.367
R612 B.n319 B.n318 163.367
R613 B.n319 B.n172 163.367
R614 B.n323 B.n172 163.367
R615 B.n324 B.n323 163.367
R616 B.n325 B.n324 163.367
R617 B.n325 B.n170 163.367
R618 B.n329 B.n170 163.367
R619 B.n330 B.n329 163.367
R620 B.n331 B.n330 163.367
R621 B.n331 B.n168 163.367
R622 B.n335 B.n168 163.367
R623 B.n336 B.n335 163.367
R624 B.n337 B.n336 163.367
R625 B.n337 B.n166 163.367
R626 B.n341 B.n166 163.367
R627 B.n342 B.n341 163.367
R628 B.n343 B.n342 163.367
R629 B.n343 B.n164 163.367
R630 B.n347 B.n164 163.367
R631 B.n348 B.n347 163.367
R632 B.n349 B.n348 163.367
R633 B.n349 B.n160 163.367
R634 B.n354 B.n160 163.367
R635 B.n355 B.n354 163.367
R636 B.n356 B.n355 163.367
R637 B.n356 B.n158 163.367
R638 B.n360 B.n158 163.367
R639 B.n361 B.n360 163.367
R640 B.n362 B.n361 163.367
R641 B.n362 B.n156 163.367
R642 B.n369 B.n156 163.367
R643 B.n370 B.n369 163.367
R644 B.n371 B.n370 163.367
R645 B.n371 B.n154 163.367
R646 B.n375 B.n154 163.367
R647 B.n376 B.n375 163.367
R648 B.n377 B.n376 163.367
R649 B.n377 B.n152 163.367
R650 B.n381 B.n152 163.367
R651 B.n382 B.n381 163.367
R652 B.n383 B.n382 163.367
R653 B.n383 B.n150 163.367
R654 B.n387 B.n150 163.367
R655 B.n388 B.n387 163.367
R656 B.n389 B.n388 163.367
R657 B.n389 B.n148 163.367
R658 B.n393 B.n148 163.367
R659 B.n394 B.n393 163.367
R660 B.n395 B.n394 163.367
R661 B.n395 B.n146 163.367
R662 B.n399 B.n146 163.367
R663 B.n400 B.n399 163.367
R664 B.n401 B.n400 163.367
R665 B.n401 B.n144 163.367
R666 B.n405 B.n144 163.367
R667 B.n406 B.n405 163.367
R668 B.n407 B.n406 163.367
R669 B.n407 B.n142 163.367
R670 B.n411 B.n142 163.367
R671 B.n412 B.n411 163.367
R672 B.n413 B.n412 163.367
R673 B.n413 B.n140 163.367
R674 B.n417 B.n140 163.367
R675 B.n418 B.n417 163.367
R676 B.n419 B.n418 163.367
R677 B.n419 B.n138 163.367
R678 B.n423 B.n138 163.367
R679 B.n424 B.n423 163.367
R680 B.n425 B.n424 163.367
R681 B.n425 B.n136 163.367
R682 B.n429 B.n136 163.367
R683 B.n430 B.n429 163.367
R684 B.n431 B.n430 163.367
R685 B.n431 B.n134 163.367
R686 B.n435 B.n134 163.367
R687 B.n436 B.n435 163.367
R688 B.n437 B.n436 163.367
R689 B.n437 B.n132 163.367
R690 B.n586 B.n585 163.367
R691 B.n585 B.n84 163.367
R692 B.n581 B.n84 163.367
R693 B.n581 B.n580 163.367
R694 B.n580 B.n579 163.367
R695 B.n579 B.n86 163.367
R696 B.n575 B.n86 163.367
R697 B.n575 B.n574 163.367
R698 B.n574 B.n573 163.367
R699 B.n573 B.n88 163.367
R700 B.n569 B.n88 163.367
R701 B.n569 B.n568 163.367
R702 B.n568 B.n567 163.367
R703 B.n567 B.n90 163.367
R704 B.n563 B.n90 163.367
R705 B.n563 B.n562 163.367
R706 B.n562 B.n561 163.367
R707 B.n561 B.n92 163.367
R708 B.n557 B.n92 163.367
R709 B.n557 B.n556 163.367
R710 B.n556 B.n555 163.367
R711 B.n555 B.n94 163.367
R712 B.n551 B.n94 163.367
R713 B.n551 B.n550 163.367
R714 B.n550 B.n549 163.367
R715 B.n549 B.n96 163.367
R716 B.n545 B.n96 163.367
R717 B.n545 B.n544 163.367
R718 B.n544 B.n543 163.367
R719 B.n543 B.n98 163.367
R720 B.n539 B.n98 163.367
R721 B.n539 B.n538 163.367
R722 B.n538 B.n537 163.367
R723 B.n537 B.n100 163.367
R724 B.n533 B.n100 163.367
R725 B.n533 B.n532 163.367
R726 B.n532 B.n531 163.367
R727 B.n531 B.n102 163.367
R728 B.n527 B.n102 163.367
R729 B.n527 B.n526 163.367
R730 B.n526 B.n525 163.367
R731 B.n525 B.n104 163.367
R732 B.n521 B.n104 163.367
R733 B.n521 B.n520 163.367
R734 B.n520 B.n519 163.367
R735 B.n519 B.n106 163.367
R736 B.n515 B.n106 163.367
R737 B.n515 B.n514 163.367
R738 B.n514 B.n513 163.367
R739 B.n513 B.n108 163.367
R740 B.n509 B.n108 163.367
R741 B.n509 B.n508 163.367
R742 B.n508 B.n507 163.367
R743 B.n507 B.n110 163.367
R744 B.n503 B.n110 163.367
R745 B.n503 B.n502 163.367
R746 B.n502 B.n501 163.367
R747 B.n501 B.n112 163.367
R748 B.n497 B.n112 163.367
R749 B.n497 B.n496 163.367
R750 B.n496 B.n495 163.367
R751 B.n495 B.n114 163.367
R752 B.n491 B.n114 163.367
R753 B.n491 B.n490 163.367
R754 B.n490 B.n489 163.367
R755 B.n489 B.n116 163.367
R756 B.n485 B.n116 163.367
R757 B.n485 B.n484 163.367
R758 B.n484 B.n483 163.367
R759 B.n483 B.n118 163.367
R760 B.n479 B.n118 163.367
R761 B.n479 B.n478 163.367
R762 B.n478 B.n477 163.367
R763 B.n477 B.n120 163.367
R764 B.n473 B.n120 163.367
R765 B.n473 B.n472 163.367
R766 B.n472 B.n471 163.367
R767 B.n471 B.n122 163.367
R768 B.n467 B.n122 163.367
R769 B.n467 B.n466 163.367
R770 B.n466 B.n465 163.367
R771 B.n465 B.n124 163.367
R772 B.n461 B.n124 163.367
R773 B.n461 B.n460 163.367
R774 B.n460 B.n459 163.367
R775 B.n459 B.n126 163.367
R776 B.n455 B.n126 163.367
R777 B.n455 B.n454 163.367
R778 B.n454 B.n453 163.367
R779 B.n453 B.n128 163.367
R780 B.n449 B.n128 163.367
R781 B.n449 B.n448 163.367
R782 B.n448 B.n447 163.367
R783 B.n447 B.n130 163.367
R784 B.n443 B.n130 163.367
R785 B.n443 B.n442 163.367
R786 B.n442 B.n441 163.367
R787 B.n743 B.n742 163.367
R788 B.n742 B.n27 163.367
R789 B.n738 B.n27 163.367
R790 B.n738 B.n737 163.367
R791 B.n737 B.n736 163.367
R792 B.n736 B.n29 163.367
R793 B.n732 B.n29 163.367
R794 B.n732 B.n731 163.367
R795 B.n731 B.n730 163.367
R796 B.n730 B.n31 163.367
R797 B.n726 B.n31 163.367
R798 B.n726 B.n725 163.367
R799 B.n725 B.n724 163.367
R800 B.n724 B.n33 163.367
R801 B.n720 B.n33 163.367
R802 B.n720 B.n719 163.367
R803 B.n719 B.n718 163.367
R804 B.n718 B.n35 163.367
R805 B.n714 B.n35 163.367
R806 B.n714 B.n713 163.367
R807 B.n713 B.n712 163.367
R808 B.n712 B.n37 163.367
R809 B.n708 B.n37 163.367
R810 B.n708 B.n707 163.367
R811 B.n707 B.n706 163.367
R812 B.n706 B.n39 163.367
R813 B.n702 B.n39 163.367
R814 B.n702 B.n701 163.367
R815 B.n701 B.n700 163.367
R816 B.n700 B.n41 163.367
R817 B.n696 B.n41 163.367
R818 B.n696 B.n695 163.367
R819 B.n695 B.n694 163.367
R820 B.n694 B.n43 163.367
R821 B.n690 B.n43 163.367
R822 B.n690 B.n689 163.367
R823 B.n689 B.n688 163.367
R824 B.n688 B.n45 163.367
R825 B.n684 B.n45 163.367
R826 B.n684 B.n683 163.367
R827 B.n683 B.n682 163.367
R828 B.n682 B.n47 163.367
R829 B.n678 B.n47 163.367
R830 B.n678 B.n677 163.367
R831 B.n677 B.n676 163.367
R832 B.n676 B.n49 163.367
R833 B.n671 B.n49 163.367
R834 B.n671 B.n670 163.367
R835 B.n670 B.n669 163.367
R836 B.n669 B.n53 163.367
R837 B.n665 B.n53 163.367
R838 B.n665 B.n664 163.367
R839 B.n664 B.n663 163.367
R840 B.n663 B.n55 163.367
R841 B.n659 B.n55 163.367
R842 B.n659 B.n658 163.367
R843 B.n658 B.n657 163.367
R844 B.n657 B.n57 163.367
R845 B.n653 B.n57 163.367
R846 B.n653 B.n652 163.367
R847 B.n652 B.n651 163.367
R848 B.n651 B.n62 163.367
R849 B.n647 B.n62 163.367
R850 B.n647 B.n646 163.367
R851 B.n646 B.n645 163.367
R852 B.n645 B.n64 163.367
R853 B.n641 B.n64 163.367
R854 B.n641 B.n640 163.367
R855 B.n640 B.n639 163.367
R856 B.n639 B.n66 163.367
R857 B.n635 B.n66 163.367
R858 B.n635 B.n634 163.367
R859 B.n634 B.n633 163.367
R860 B.n633 B.n68 163.367
R861 B.n629 B.n68 163.367
R862 B.n629 B.n628 163.367
R863 B.n628 B.n627 163.367
R864 B.n627 B.n70 163.367
R865 B.n623 B.n70 163.367
R866 B.n623 B.n622 163.367
R867 B.n622 B.n621 163.367
R868 B.n621 B.n72 163.367
R869 B.n617 B.n72 163.367
R870 B.n617 B.n616 163.367
R871 B.n616 B.n615 163.367
R872 B.n615 B.n74 163.367
R873 B.n611 B.n74 163.367
R874 B.n611 B.n610 163.367
R875 B.n610 B.n609 163.367
R876 B.n609 B.n76 163.367
R877 B.n605 B.n76 163.367
R878 B.n605 B.n604 163.367
R879 B.n604 B.n603 163.367
R880 B.n603 B.n78 163.367
R881 B.n599 B.n78 163.367
R882 B.n599 B.n598 163.367
R883 B.n598 B.n597 163.367
R884 B.n597 B.n80 163.367
R885 B.n593 B.n80 163.367
R886 B.n593 B.n592 163.367
R887 B.n592 B.n591 163.367
R888 B.n591 B.n82 163.367
R889 B.n587 B.n82 163.367
R890 B.n744 B.n25 163.367
R891 B.n748 B.n25 163.367
R892 B.n749 B.n748 163.367
R893 B.n750 B.n749 163.367
R894 B.n750 B.n23 163.367
R895 B.n754 B.n23 163.367
R896 B.n755 B.n754 163.367
R897 B.n756 B.n755 163.367
R898 B.n756 B.n21 163.367
R899 B.n760 B.n21 163.367
R900 B.n761 B.n760 163.367
R901 B.n762 B.n761 163.367
R902 B.n762 B.n19 163.367
R903 B.n766 B.n19 163.367
R904 B.n767 B.n766 163.367
R905 B.n768 B.n767 163.367
R906 B.n768 B.n17 163.367
R907 B.n772 B.n17 163.367
R908 B.n773 B.n772 163.367
R909 B.n774 B.n773 163.367
R910 B.n774 B.n15 163.367
R911 B.n778 B.n15 163.367
R912 B.n779 B.n778 163.367
R913 B.n780 B.n779 163.367
R914 B.n780 B.n13 163.367
R915 B.n784 B.n13 163.367
R916 B.n785 B.n784 163.367
R917 B.n786 B.n785 163.367
R918 B.n786 B.n11 163.367
R919 B.n790 B.n11 163.367
R920 B.n791 B.n790 163.367
R921 B.n792 B.n791 163.367
R922 B.n792 B.n9 163.367
R923 B.n796 B.n9 163.367
R924 B.n797 B.n796 163.367
R925 B.n798 B.n797 163.367
R926 B.n798 B.n7 163.367
R927 B.n802 B.n7 163.367
R928 B.n803 B.n802 163.367
R929 B.n804 B.n803 163.367
R930 B.n804 B.n5 163.367
R931 B.n808 B.n5 163.367
R932 B.n809 B.n808 163.367
R933 B.n810 B.n809 163.367
R934 B.n810 B.n3 163.367
R935 B.n814 B.n3 163.367
R936 B.n815 B.n814 163.367
R937 B.n210 B.n2 163.367
R938 B.n211 B.n210 163.367
R939 B.n211 B.n208 163.367
R940 B.n215 B.n208 163.367
R941 B.n216 B.n215 163.367
R942 B.n217 B.n216 163.367
R943 B.n217 B.n206 163.367
R944 B.n221 B.n206 163.367
R945 B.n222 B.n221 163.367
R946 B.n223 B.n222 163.367
R947 B.n223 B.n204 163.367
R948 B.n227 B.n204 163.367
R949 B.n228 B.n227 163.367
R950 B.n229 B.n228 163.367
R951 B.n229 B.n202 163.367
R952 B.n233 B.n202 163.367
R953 B.n234 B.n233 163.367
R954 B.n235 B.n234 163.367
R955 B.n235 B.n200 163.367
R956 B.n239 B.n200 163.367
R957 B.n240 B.n239 163.367
R958 B.n241 B.n240 163.367
R959 B.n241 B.n198 163.367
R960 B.n245 B.n198 163.367
R961 B.n246 B.n245 163.367
R962 B.n247 B.n246 163.367
R963 B.n247 B.n196 163.367
R964 B.n251 B.n196 163.367
R965 B.n252 B.n251 163.367
R966 B.n253 B.n252 163.367
R967 B.n253 B.n194 163.367
R968 B.n257 B.n194 163.367
R969 B.n258 B.n257 163.367
R970 B.n259 B.n258 163.367
R971 B.n259 B.n192 163.367
R972 B.n263 B.n192 163.367
R973 B.n264 B.n263 163.367
R974 B.n265 B.n264 163.367
R975 B.n265 B.n190 163.367
R976 B.n269 B.n190 163.367
R977 B.n270 B.n269 163.367
R978 B.n271 B.n270 163.367
R979 B.n271 B.n188 163.367
R980 B.n275 B.n188 163.367
R981 B.n276 B.n275 163.367
R982 B.n277 B.n276 163.367
R983 B.n277 B.n186 163.367
R984 B.n366 B.t8 112.358
R985 B.n59 B.t1 112.358
R986 B.n162 B.t5 112.341
R987 B.n51 B.t10 112.341
R988 B.n162 B.n161 66.7156
R989 B.n366 B.n365 66.7156
R990 B.n59 B.n58 66.7156
R991 B.n51 B.n50 66.7156
R992 B.n351 B.n162 59.5399
R993 B.n367 B.n366 59.5399
R994 B.n60 B.n59 59.5399
R995 B.n673 B.n51 59.5399
R996 B.n745 B.n26 32.9371
R997 B.n588 B.n83 32.9371
R998 B.n440 B.n439 32.9371
R999 B.n280 B.n279 32.9371
R1000 B B.n817 18.0485
R1001 B.n746 B.n745 10.6151
R1002 B.n747 B.n746 10.6151
R1003 B.n747 B.n24 10.6151
R1004 B.n751 B.n24 10.6151
R1005 B.n752 B.n751 10.6151
R1006 B.n753 B.n752 10.6151
R1007 B.n753 B.n22 10.6151
R1008 B.n757 B.n22 10.6151
R1009 B.n758 B.n757 10.6151
R1010 B.n759 B.n758 10.6151
R1011 B.n759 B.n20 10.6151
R1012 B.n763 B.n20 10.6151
R1013 B.n764 B.n763 10.6151
R1014 B.n765 B.n764 10.6151
R1015 B.n765 B.n18 10.6151
R1016 B.n769 B.n18 10.6151
R1017 B.n770 B.n769 10.6151
R1018 B.n771 B.n770 10.6151
R1019 B.n771 B.n16 10.6151
R1020 B.n775 B.n16 10.6151
R1021 B.n776 B.n775 10.6151
R1022 B.n777 B.n776 10.6151
R1023 B.n777 B.n14 10.6151
R1024 B.n781 B.n14 10.6151
R1025 B.n782 B.n781 10.6151
R1026 B.n783 B.n782 10.6151
R1027 B.n783 B.n12 10.6151
R1028 B.n787 B.n12 10.6151
R1029 B.n788 B.n787 10.6151
R1030 B.n789 B.n788 10.6151
R1031 B.n789 B.n10 10.6151
R1032 B.n793 B.n10 10.6151
R1033 B.n794 B.n793 10.6151
R1034 B.n795 B.n794 10.6151
R1035 B.n795 B.n8 10.6151
R1036 B.n799 B.n8 10.6151
R1037 B.n800 B.n799 10.6151
R1038 B.n801 B.n800 10.6151
R1039 B.n801 B.n6 10.6151
R1040 B.n805 B.n6 10.6151
R1041 B.n806 B.n805 10.6151
R1042 B.n807 B.n806 10.6151
R1043 B.n807 B.n4 10.6151
R1044 B.n811 B.n4 10.6151
R1045 B.n812 B.n811 10.6151
R1046 B.n813 B.n812 10.6151
R1047 B.n813 B.n0 10.6151
R1048 B.n741 B.n26 10.6151
R1049 B.n741 B.n740 10.6151
R1050 B.n740 B.n739 10.6151
R1051 B.n739 B.n28 10.6151
R1052 B.n735 B.n28 10.6151
R1053 B.n735 B.n734 10.6151
R1054 B.n734 B.n733 10.6151
R1055 B.n733 B.n30 10.6151
R1056 B.n729 B.n30 10.6151
R1057 B.n729 B.n728 10.6151
R1058 B.n728 B.n727 10.6151
R1059 B.n727 B.n32 10.6151
R1060 B.n723 B.n32 10.6151
R1061 B.n723 B.n722 10.6151
R1062 B.n722 B.n721 10.6151
R1063 B.n721 B.n34 10.6151
R1064 B.n717 B.n34 10.6151
R1065 B.n717 B.n716 10.6151
R1066 B.n716 B.n715 10.6151
R1067 B.n715 B.n36 10.6151
R1068 B.n711 B.n36 10.6151
R1069 B.n711 B.n710 10.6151
R1070 B.n710 B.n709 10.6151
R1071 B.n709 B.n38 10.6151
R1072 B.n705 B.n38 10.6151
R1073 B.n705 B.n704 10.6151
R1074 B.n704 B.n703 10.6151
R1075 B.n703 B.n40 10.6151
R1076 B.n699 B.n40 10.6151
R1077 B.n699 B.n698 10.6151
R1078 B.n698 B.n697 10.6151
R1079 B.n697 B.n42 10.6151
R1080 B.n693 B.n42 10.6151
R1081 B.n693 B.n692 10.6151
R1082 B.n692 B.n691 10.6151
R1083 B.n691 B.n44 10.6151
R1084 B.n687 B.n44 10.6151
R1085 B.n687 B.n686 10.6151
R1086 B.n686 B.n685 10.6151
R1087 B.n685 B.n46 10.6151
R1088 B.n681 B.n46 10.6151
R1089 B.n681 B.n680 10.6151
R1090 B.n680 B.n679 10.6151
R1091 B.n679 B.n48 10.6151
R1092 B.n675 B.n48 10.6151
R1093 B.n675 B.n674 10.6151
R1094 B.n672 B.n52 10.6151
R1095 B.n668 B.n52 10.6151
R1096 B.n668 B.n667 10.6151
R1097 B.n667 B.n666 10.6151
R1098 B.n666 B.n54 10.6151
R1099 B.n662 B.n54 10.6151
R1100 B.n662 B.n661 10.6151
R1101 B.n661 B.n660 10.6151
R1102 B.n660 B.n56 10.6151
R1103 B.n656 B.n655 10.6151
R1104 B.n655 B.n654 10.6151
R1105 B.n654 B.n61 10.6151
R1106 B.n650 B.n61 10.6151
R1107 B.n650 B.n649 10.6151
R1108 B.n649 B.n648 10.6151
R1109 B.n648 B.n63 10.6151
R1110 B.n644 B.n63 10.6151
R1111 B.n644 B.n643 10.6151
R1112 B.n643 B.n642 10.6151
R1113 B.n642 B.n65 10.6151
R1114 B.n638 B.n65 10.6151
R1115 B.n638 B.n637 10.6151
R1116 B.n637 B.n636 10.6151
R1117 B.n636 B.n67 10.6151
R1118 B.n632 B.n67 10.6151
R1119 B.n632 B.n631 10.6151
R1120 B.n631 B.n630 10.6151
R1121 B.n630 B.n69 10.6151
R1122 B.n626 B.n69 10.6151
R1123 B.n626 B.n625 10.6151
R1124 B.n625 B.n624 10.6151
R1125 B.n624 B.n71 10.6151
R1126 B.n620 B.n71 10.6151
R1127 B.n620 B.n619 10.6151
R1128 B.n619 B.n618 10.6151
R1129 B.n618 B.n73 10.6151
R1130 B.n614 B.n73 10.6151
R1131 B.n614 B.n613 10.6151
R1132 B.n613 B.n612 10.6151
R1133 B.n612 B.n75 10.6151
R1134 B.n608 B.n75 10.6151
R1135 B.n608 B.n607 10.6151
R1136 B.n607 B.n606 10.6151
R1137 B.n606 B.n77 10.6151
R1138 B.n602 B.n77 10.6151
R1139 B.n602 B.n601 10.6151
R1140 B.n601 B.n600 10.6151
R1141 B.n600 B.n79 10.6151
R1142 B.n596 B.n79 10.6151
R1143 B.n596 B.n595 10.6151
R1144 B.n595 B.n594 10.6151
R1145 B.n594 B.n81 10.6151
R1146 B.n590 B.n81 10.6151
R1147 B.n590 B.n589 10.6151
R1148 B.n589 B.n588 10.6151
R1149 B.n584 B.n83 10.6151
R1150 B.n584 B.n583 10.6151
R1151 B.n583 B.n582 10.6151
R1152 B.n582 B.n85 10.6151
R1153 B.n578 B.n85 10.6151
R1154 B.n578 B.n577 10.6151
R1155 B.n577 B.n576 10.6151
R1156 B.n576 B.n87 10.6151
R1157 B.n572 B.n87 10.6151
R1158 B.n572 B.n571 10.6151
R1159 B.n571 B.n570 10.6151
R1160 B.n570 B.n89 10.6151
R1161 B.n566 B.n89 10.6151
R1162 B.n566 B.n565 10.6151
R1163 B.n565 B.n564 10.6151
R1164 B.n564 B.n91 10.6151
R1165 B.n560 B.n91 10.6151
R1166 B.n560 B.n559 10.6151
R1167 B.n559 B.n558 10.6151
R1168 B.n558 B.n93 10.6151
R1169 B.n554 B.n93 10.6151
R1170 B.n554 B.n553 10.6151
R1171 B.n553 B.n552 10.6151
R1172 B.n552 B.n95 10.6151
R1173 B.n548 B.n95 10.6151
R1174 B.n548 B.n547 10.6151
R1175 B.n547 B.n546 10.6151
R1176 B.n546 B.n97 10.6151
R1177 B.n542 B.n97 10.6151
R1178 B.n542 B.n541 10.6151
R1179 B.n541 B.n540 10.6151
R1180 B.n540 B.n99 10.6151
R1181 B.n536 B.n99 10.6151
R1182 B.n536 B.n535 10.6151
R1183 B.n535 B.n534 10.6151
R1184 B.n534 B.n101 10.6151
R1185 B.n530 B.n101 10.6151
R1186 B.n530 B.n529 10.6151
R1187 B.n529 B.n528 10.6151
R1188 B.n528 B.n103 10.6151
R1189 B.n524 B.n103 10.6151
R1190 B.n524 B.n523 10.6151
R1191 B.n523 B.n522 10.6151
R1192 B.n522 B.n105 10.6151
R1193 B.n518 B.n105 10.6151
R1194 B.n518 B.n517 10.6151
R1195 B.n517 B.n516 10.6151
R1196 B.n516 B.n107 10.6151
R1197 B.n512 B.n107 10.6151
R1198 B.n512 B.n511 10.6151
R1199 B.n511 B.n510 10.6151
R1200 B.n510 B.n109 10.6151
R1201 B.n506 B.n109 10.6151
R1202 B.n506 B.n505 10.6151
R1203 B.n505 B.n504 10.6151
R1204 B.n504 B.n111 10.6151
R1205 B.n500 B.n111 10.6151
R1206 B.n500 B.n499 10.6151
R1207 B.n499 B.n498 10.6151
R1208 B.n498 B.n113 10.6151
R1209 B.n494 B.n113 10.6151
R1210 B.n494 B.n493 10.6151
R1211 B.n493 B.n492 10.6151
R1212 B.n492 B.n115 10.6151
R1213 B.n488 B.n115 10.6151
R1214 B.n488 B.n487 10.6151
R1215 B.n487 B.n486 10.6151
R1216 B.n486 B.n117 10.6151
R1217 B.n482 B.n117 10.6151
R1218 B.n482 B.n481 10.6151
R1219 B.n481 B.n480 10.6151
R1220 B.n480 B.n119 10.6151
R1221 B.n476 B.n119 10.6151
R1222 B.n476 B.n475 10.6151
R1223 B.n475 B.n474 10.6151
R1224 B.n474 B.n121 10.6151
R1225 B.n470 B.n121 10.6151
R1226 B.n470 B.n469 10.6151
R1227 B.n469 B.n468 10.6151
R1228 B.n468 B.n123 10.6151
R1229 B.n464 B.n123 10.6151
R1230 B.n464 B.n463 10.6151
R1231 B.n463 B.n462 10.6151
R1232 B.n462 B.n125 10.6151
R1233 B.n458 B.n125 10.6151
R1234 B.n458 B.n457 10.6151
R1235 B.n457 B.n456 10.6151
R1236 B.n456 B.n127 10.6151
R1237 B.n452 B.n127 10.6151
R1238 B.n452 B.n451 10.6151
R1239 B.n451 B.n450 10.6151
R1240 B.n450 B.n129 10.6151
R1241 B.n446 B.n129 10.6151
R1242 B.n446 B.n445 10.6151
R1243 B.n445 B.n444 10.6151
R1244 B.n444 B.n131 10.6151
R1245 B.n440 B.n131 10.6151
R1246 B.n209 B.n1 10.6151
R1247 B.n212 B.n209 10.6151
R1248 B.n213 B.n212 10.6151
R1249 B.n214 B.n213 10.6151
R1250 B.n214 B.n207 10.6151
R1251 B.n218 B.n207 10.6151
R1252 B.n219 B.n218 10.6151
R1253 B.n220 B.n219 10.6151
R1254 B.n220 B.n205 10.6151
R1255 B.n224 B.n205 10.6151
R1256 B.n225 B.n224 10.6151
R1257 B.n226 B.n225 10.6151
R1258 B.n226 B.n203 10.6151
R1259 B.n230 B.n203 10.6151
R1260 B.n231 B.n230 10.6151
R1261 B.n232 B.n231 10.6151
R1262 B.n232 B.n201 10.6151
R1263 B.n236 B.n201 10.6151
R1264 B.n237 B.n236 10.6151
R1265 B.n238 B.n237 10.6151
R1266 B.n238 B.n199 10.6151
R1267 B.n242 B.n199 10.6151
R1268 B.n243 B.n242 10.6151
R1269 B.n244 B.n243 10.6151
R1270 B.n244 B.n197 10.6151
R1271 B.n248 B.n197 10.6151
R1272 B.n249 B.n248 10.6151
R1273 B.n250 B.n249 10.6151
R1274 B.n250 B.n195 10.6151
R1275 B.n254 B.n195 10.6151
R1276 B.n255 B.n254 10.6151
R1277 B.n256 B.n255 10.6151
R1278 B.n256 B.n193 10.6151
R1279 B.n260 B.n193 10.6151
R1280 B.n261 B.n260 10.6151
R1281 B.n262 B.n261 10.6151
R1282 B.n262 B.n191 10.6151
R1283 B.n266 B.n191 10.6151
R1284 B.n267 B.n266 10.6151
R1285 B.n268 B.n267 10.6151
R1286 B.n268 B.n189 10.6151
R1287 B.n272 B.n189 10.6151
R1288 B.n273 B.n272 10.6151
R1289 B.n274 B.n273 10.6151
R1290 B.n274 B.n187 10.6151
R1291 B.n278 B.n187 10.6151
R1292 B.n279 B.n278 10.6151
R1293 B.n280 B.n185 10.6151
R1294 B.n284 B.n185 10.6151
R1295 B.n285 B.n284 10.6151
R1296 B.n286 B.n285 10.6151
R1297 B.n286 B.n183 10.6151
R1298 B.n290 B.n183 10.6151
R1299 B.n291 B.n290 10.6151
R1300 B.n292 B.n291 10.6151
R1301 B.n292 B.n181 10.6151
R1302 B.n296 B.n181 10.6151
R1303 B.n297 B.n296 10.6151
R1304 B.n298 B.n297 10.6151
R1305 B.n298 B.n179 10.6151
R1306 B.n302 B.n179 10.6151
R1307 B.n303 B.n302 10.6151
R1308 B.n304 B.n303 10.6151
R1309 B.n304 B.n177 10.6151
R1310 B.n308 B.n177 10.6151
R1311 B.n309 B.n308 10.6151
R1312 B.n310 B.n309 10.6151
R1313 B.n310 B.n175 10.6151
R1314 B.n314 B.n175 10.6151
R1315 B.n315 B.n314 10.6151
R1316 B.n316 B.n315 10.6151
R1317 B.n316 B.n173 10.6151
R1318 B.n320 B.n173 10.6151
R1319 B.n321 B.n320 10.6151
R1320 B.n322 B.n321 10.6151
R1321 B.n322 B.n171 10.6151
R1322 B.n326 B.n171 10.6151
R1323 B.n327 B.n326 10.6151
R1324 B.n328 B.n327 10.6151
R1325 B.n328 B.n169 10.6151
R1326 B.n332 B.n169 10.6151
R1327 B.n333 B.n332 10.6151
R1328 B.n334 B.n333 10.6151
R1329 B.n334 B.n167 10.6151
R1330 B.n338 B.n167 10.6151
R1331 B.n339 B.n338 10.6151
R1332 B.n340 B.n339 10.6151
R1333 B.n340 B.n165 10.6151
R1334 B.n344 B.n165 10.6151
R1335 B.n345 B.n344 10.6151
R1336 B.n346 B.n345 10.6151
R1337 B.n346 B.n163 10.6151
R1338 B.n350 B.n163 10.6151
R1339 B.n353 B.n352 10.6151
R1340 B.n353 B.n159 10.6151
R1341 B.n357 B.n159 10.6151
R1342 B.n358 B.n357 10.6151
R1343 B.n359 B.n358 10.6151
R1344 B.n359 B.n157 10.6151
R1345 B.n363 B.n157 10.6151
R1346 B.n364 B.n363 10.6151
R1347 B.n368 B.n364 10.6151
R1348 B.n372 B.n155 10.6151
R1349 B.n373 B.n372 10.6151
R1350 B.n374 B.n373 10.6151
R1351 B.n374 B.n153 10.6151
R1352 B.n378 B.n153 10.6151
R1353 B.n379 B.n378 10.6151
R1354 B.n380 B.n379 10.6151
R1355 B.n380 B.n151 10.6151
R1356 B.n384 B.n151 10.6151
R1357 B.n385 B.n384 10.6151
R1358 B.n386 B.n385 10.6151
R1359 B.n386 B.n149 10.6151
R1360 B.n390 B.n149 10.6151
R1361 B.n391 B.n390 10.6151
R1362 B.n392 B.n391 10.6151
R1363 B.n392 B.n147 10.6151
R1364 B.n396 B.n147 10.6151
R1365 B.n397 B.n396 10.6151
R1366 B.n398 B.n397 10.6151
R1367 B.n398 B.n145 10.6151
R1368 B.n402 B.n145 10.6151
R1369 B.n403 B.n402 10.6151
R1370 B.n404 B.n403 10.6151
R1371 B.n404 B.n143 10.6151
R1372 B.n408 B.n143 10.6151
R1373 B.n409 B.n408 10.6151
R1374 B.n410 B.n409 10.6151
R1375 B.n410 B.n141 10.6151
R1376 B.n414 B.n141 10.6151
R1377 B.n415 B.n414 10.6151
R1378 B.n416 B.n415 10.6151
R1379 B.n416 B.n139 10.6151
R1380 B.n420 B.n139 10.6151
R1381 B.n421 B.n420 10.6151
R1382 B.n422 B.n421 10.6151
R1383 B.n422 B.n137 10.6151
R1384 B.n426 B.n137 10.6151
R1385 B.n427 B.n426 10.6151
R1386 B.n428 B.n427 10.6151
R1387 B.n428 B.n135 10.6151
R1388 B.n432 B.n135 10.6151
R1389 B.n433 B.n432 10.6151
R1390 B.n434 B.n433 10.6151
R1391 B.n434 B.n133 10.6151
R1392 B.n438 B.n133 10.6151
R1393 B.n439 B.n438 10.6151
R1394 B.n674 B.n673 9.36635
R1395 B.n656 B.n60 9.36635
R1396 B.n351 B.n350 9.36635
R1397 B.n367 B.n155 9.36635
R1398 B.n817 B.n0 8.11757
R1399 B.n817 B.n1 8.11757
R1400 B.n673 B.n672 1.24928
R1401 B.n60 B.n56 1.24928
R1402 B.n352 B.n351 1.24928
R1403 B.n368 B.n367 1.24928
C0 VDD2 VP 0.50178f
C1 w_n3722_n3746# VTAIL 3.27979f
C2 VDD1 B 2.3775f
C3 VN B 1.29692f
C4 w_n3722_n3746# VDD2 2.64807f
C5 VN VDD1 0.151525f
C6 w_n3722_n3746# VP 7.68717f
C7 B VTAIL 4.32986f
C8 VDD1 VTAIL 8.50765f
C9 VN VTAIL 8.163401f
C10 VDD2 B 2.46383f
C11 VDD1 VDD2 1.60669f
C12 VP B 2.10528f
C13 VDD1 VP 8.31451f
C14 VN VDD2 7.96764f
C15 VN VP 7.77176f
C16 w_n3722_n3746# B 10.910599f
C17 w_n3722_n3746# VDD1 2.54671f
C18 VDD2 VTAIL 8.56202f
C19 VN w_n3722_n3746# 7.20454f
C20 VP VTAIL 8.17768f
C21 VDD2 VSUBS 2.106896f
C22 VDD1 VSUBS 2.63141f
C23 VTAIL VSUBS 1.360798f
C24 VN VSUBS 6.40411f
C25 VP VSUBS 3.414034f
C26 B VSUBS 5.30198f
C27 w_n3722_n3746# VSUBS 0.171197p
C28 B.n0 VSUBS 0.007251f
C29 B.n1 VSUBS 0.007251f
C30 B.n2 VSUBS 0.010724f
C31 B.n3 VSUBS 0.008218f
C32 B.n4 VSUBS 0.008218f
C33 B.n5 VSUBS 0.008218f
C34 B.n6 VSUBS 0.008218f
C35 B.n7 VSUBS 0.008218f
C36 B.n8 VSUBS 0.008218f
C37 B.n9 VSUBS 0.008218f
C38 B.n10 VSUBS 0.008218f
C39 B.n11 VSUBS 0.008218f
C40 B.n12 VSUBS 0.008218f
C41 B.n13 VSUBS 0.008218f
C42 B.n14 VSUBS 0.008218f
C43 B.n15 VSUBS 0.008218f
C44 B.n16 VSUBS 0.008218f
C45 B.n17 VSUBS 0.008218f
C46 B.n18 VSUBS 0.008218f
C47 B.n19 VSUBS 0.008218f
C48 B.n20 VSUBS 0.008218f
C49 B.n21 VSUBS 0.008218f
C50 B.n22 VSUBS 0.008218f
C51 B.n23 VSUBS 0.008218f
C52 B.n24 VSUBS 0.008218f
C53 B.n25 VSUBS 0.008218f
C54 B.n26 VSUBS 0.019888f
C55 B.n27 VSUBS 0.008218f
C56 B.n28 VSUBS 0.008218f
C57 B.n29 VSUBS 0.008218f
C58 B.n30 VSUBS 0.008218f
C59 B.n31 VSUBS 0.008218f
C60 B.n32 VSUBS 0.008218f
C61 B.n33 VSUBS 0.008218f
C62 B.n34 VSUBS 0.008218f
C63 B.n35 VSUBS 0.008218f
C64 B.n36 VSUBS 0.008218f
C65 B.n37 VSUBS 0.008218f
C66 B.n38 VSUBS 0.008218f
C67 B.n39 VSUBS 0.008218f
C68 B.n40 VSUBS 0.008218f
C69 B.n41 VSUBS 0.008218f
C70 B.n42 VSUBS 0.008218f
C71 B.n43 VSUBS 0.008218f
C72 B.n44 VSUBS 0.008218f
C73 B.n45 VSUBS 0.008218f
C74 B.n46 VSUBS 0.008218f
C75 B.n47 VSUBS 0.008218f
C76 B.n48 VSUBS 0.008218f
C77 B.n49 VSUBS 0.008218f
C78 B.t10 VSUBS 0.539191f
C79 B.t11 VSUBS 0.567201f
C80 B.t9 VSUBS 2.31687f
C81 B.n50 VSUBS 0.316755f
C82 B.n51 VSUBS 0.086895f
C83 B.n52 VSUBS 0.008218f
C84 B.n53 VSUBS 0.008218f
C85 B.n54 VSUBS 0.008218f
C86 B.n55 VSUBS 0.008218f
C87 B.n56 VSUBS 0.004592f
C88 B.n57 VSUBS 0.008218f
C89 B.t1 VSUBS 0.539178f
C90 B.t2 VSUBS 0.56719f
C91 B.t0 VSUBS 2.31687f
C92 B.n58 VSUBS 0.316765f
C93 B.n59 VSUBS 0.086908f
C94 B.n60 VSUBS 0.01904f
C95 B.n61 VSUBS 0.008218f
C96 B.n62 VSUBS 0.008218f
C97 B.n63 VSUBS 0.008218f
C98 B.n64 VSUBS 0.008218f
C99 B.n65 VSUBS 0.008218f
C100 B.n66 VSUBS 0.008218f
C101 B.n67 VSUBS 0.008218f
C102 B.n68 VSUBS 0.008218f
C103 B.n69 VSUBS 0.008218f
C104 B.n70 VSUBS 0.008218f
C105 B.n71 VSUBS 0.008218f
C106 B.n72 VSUBS 0.008218f
C107 B.n73 VSUBS 0.008218f
C108 B.n74 VSUBS 0.008218f
C109 B.n75 VSUBS 0.008218f
C110 B.n76 VSUBS 0.008218f
C111 B.n77 VSUBS 0.008218f
C112 B.n78 VSUBS 0.008218f
C113 B.n79 VSUBS 0.008218f
C114 B.n80 VSUBS 0.008218f
C115 B.n81 VSUBS 0.008218f
C116 B.n82 VSUBS 0.008218f
C117 B.n83 VSUBS 0.018784f
C118 B.n84 VSUBS 0.008218f
C119 B.n85 VSUBS 0.008218f
C120 B.n86 VSUBS 0.008218f
C121 B.n87 VSUBS 0.008218f
C122 B.n88 VSUBS 0.008218f
C123 B.n89 VSUBS 0.008218f
C124 B.n90 VSUBS 0.008218f
C125 B.n91 VSUBS 0.008218f
C126 B.n92 VSUBS 0.008218f
C127 B.n93 VSUBS 0.008218f
C128 B.n94 VSUBS 0.008218f
C129 B.n95 VSUBS 0.008218f
C130 B.n96 VSUBS 0.008218f
C131 B.n97 VSUBS 0.008218f
C132 B.n98 VSUBS 0.008218f
C133 B.n99 VSUBS 0.008218f
C134 B.n100 VSUBS 0.008218f
C135 B.n101 VSUBS 0.008218f
C136 B.n102 VSUBS 0.008218f
C137 B.n103 VSUBS 0.008218f
C138 B.n104 VSUBS 0.008218f
C139 B.n105 VSUBS 0.008218f
C140 B.n106 VSUBS 0.008218f
C141 B.n107 VSUBS 0.008218f
C142 B.n108 VSUBS 0.008218f
C143 B.n109 VSUBS 0.008218f
C144 B.n110 VSUBS 0.008218f
C145 B.n111 VSUBS 0.008218f
C146 B.n112 VSUBS 0.008218f
C147 B.n113 VSUBS 0.008218f
C148 B.n114 VSUBS 0.008218f
C149 B.n115 VSUBS 0.008218f
C150 B.n116 VSUBS 0.008218f
C151 B.n117 VSUBS 0.008218f
C152 B.n118 VSUBS 0.008218f
C153 B.n119 VSUBS 0.008218f
C154 B.n120 VSUBS 0.008218f
C155 B.n121 VSUBS 0.008218f
C156 B.n122 VSUBS 0.008218f
C157 B.n123 VSUBS 0.008218f
C158 B.n124 VSUBS 0.008218f
C159 B.n125 VSUBS 0.008218f
C160 B.n126 VSUBS 0.008218f
C161 B.n127 VSUBS 0.008218f
C162 B.n128 VSUBS 0.008218f
C163 B.n129 VSUBS 0.008218f
C164 B.n130 VSUBS 0.008218f
C165 B.n131 VSUBS 0.008218f
C166 B.n132 VSUBS 0.019888f
C167 B.n133 VSUBS 0.008218f
C168 B.n134 VSUBS 0.008218f
C169 B.n135 VSUBS 0.008218f
C170 B.n136 VSUBS 0.008218f
C171 B.n137 VSUBS 0.008218f
C172 B.n138 VSUBS 0.008218f
C173 B.n139 VSUBS 0.008218f
C174 B.n140 VSUBS 0.008218f
C175 B.n141 VSUBS 0.008218f
C176 B.n142 VSUBS 0.008218f
C177 B.n143 VSUBS 0.008218f
C178 B.n144 VSUBS 0.008218f
C179 B.n145 VSUBS 0.008218f
C180 B.n146 VSUBS 0.008218f
C181 B.n147 VSUBS 0.008218f
C182 B.n148 VSUBS 0.008218f
C183 B.n149 VSUBS 0.008218f
C184 B.n150 VSUBS 0.008218f
C185 B.n151 VSUBS 0.008218f
C186 B.n152 VSUBS 0.008218f
C187 B.n153 VSUBS 0.008218f
C188 B.n154 VSUBS 0.008218f
C189 B.n155 VSUBS 0.007734f
C190 B.n156 VSUBS 0.008218f
C191 B.n157 VSUBS 0.008218f
C192 B.n158 VSUBS 0.008218f
C193 B.n159 VSUBS 0.008218f
C194 B.n160 VSUBS 0.008218f
C195 B.t5 VSUBS 0.539191f
C196 B.t4 VSUBS 0.567201f
C197 B.t3 VSUBS 2.31687f
C198 B.n161 VSUBS 0.316755f
C199 B.n162 VSUBS 0.086895f
C200 B.n163 VSUBS 0.008218f
C201 B.n164 VSUBS 0.008218f
C202 B.n165 VSUBS 0.008218f
C203 B.n166 VSUBS 0.008218f
C204 B.n167 VSUBS 0.008218f
C205 B.n168 VSUBS 0.008218f
C206 B.n169 VSUBS 0.008218f
C207 B.n170 VSUBS 0.008218f
C208 B.n171 VSUBS 0.008218f
C209 B.n172 VSUBS 0.008218f
C210 B.n173 VSUBS 0.008218f
C211 B.n174 VSUBS 0.008218f
C212 B.n175 VSUBS 0.008218f
C213 B.n176 VSUBS 0.008218f
C214 B.n177 VSUBS 0.008218f
C215 B.n178 VSUBS 0.008218f
C216 B.n179 VSUBS 0.008218f
C217 B.n180 VSUBS 0.008218f
C218 B.n181 VSUBS 0.008218f
C219 B.n182 VSUBS 0.008218f
C220 B.n183 VSUBS 0.008218f
C221 B.n184 VSUBS 0.008218f
C222 B.n185 VSUBS 0.008218f
C223 B.n186 VSUBS 0.018784f
C224 B.n187 VSUBS 0.008218f
C225 B.n188 VSUBS 0.008218f
C226 B.n189 VSUBS 0.008218f
C227 B.n190 VSUBS 0.008218f
C228 B.n191 VSUBS 0.008218f
C229 B.n192 VSUBS 0.008218f
C230 B.n193 VSUBS 0.008218f
C231 B.n194 VSUBS 0.008218f
C232 B.n195 VSUBS 0.008218f
C233 B.n196 VSUBS 0.008218f
C234 B.n197 VSUBS 0.008218f
C235 B.n198 VSUBS 0.008218f
C236 B.n199 VSUBS 0.008218f
C237 B.n200 VSUBS 0.008218f
C238 B.n201 VSUBS 0.008218f
C239 B.n202 VSUBS 0.008218f
C240 B.n203 VSUBS 0.008218f
C241 B.n204 VSUBS 0.008218f
C242 B.n205 VSUBS 0.008218f
C243 B.n206 VSUBS 0.008218f
C244 B.n207 VSUBS 0.008218f
C245 B.n208 VSUBS 0.008218f
C246 B.n209 VSUBS 0.008218f
C247 B.n210 VSUBS 0.008218f
C248 B.n211 VSUBS 0.008218f
C249 B.n212 VSUBS 0.008218f
C250 B.n213 VSUBS 0.008218f
C251 B.n214 VSUBS 0.008218f
C252 B.n215 VSUBS 0.008218f
C253 B.n216 VSUBS 0.008218f
C254 B.n217 VSUBS 0.008218f
C255 B.n218 VSUBS 0.008218f
C256 B.n219 VSUBS 0.008218f
C257 B.n220 VSUBS 0.008218f
C258 B.n221 VSUBS 0.008218f
C259 B.n222 VSUBS 0.008218f
C260 B.n223 VSUBS 0.008218f
C261 B.n224 VSUBS 0.008218f
C262 B.n225 VSUBS 0.008218f
C263 B.n226 VSUBS 0.008218f
C264 B.n227 VSUBS 0.008218f
C265 B.n228 VSUBS 0.008218f
C266 B.n229 VSUBS 0.008218f
C267 B.n230 VSUBS 0.008218f
C268 B.n231 VSUBS 0.008218f
C269 B.n232 VSUBS 0.008218f
C270 B.n233 VSUBS 0.008218f
C271 B.n234 VSUBS 0.008218f
C272 B.n235 VSUBS 0.008218f
C273 B.n236 VSUBS 0.008218f
C274 B.n237 VSUBS 0.008218f
C275 B.n238 VSUBS 0.008218f
C276 B.n239 VSUBS 0.008218f
C277 B.n240 VSUBS 0.008218f
C278 B.n241 VSUBS 0.008218f
C279 B.n242 VSUBS 0.008218f
C280 B.n243 VSUBS 0.008218f
C281 B.n244 VSUBS 0.008218f
C282 B.n245 VSUBS 0.008218f
C283 B.n246 VSUBS 0.008218f
C284 B.n247 VSUBS 0.008218f
C285 B.n248 VSUBS 0.008218f
C286 B.n249 VSUBS 0.008218f
C287 B.n250 VSUBS 0.008218f
C288 B.n251 VSUBS 0.008218f
C289 B.n252 VSUBS 0.008218f
C290 B.n253 VSUBS 0.008218f
C291 B.n254 VSUBS 0.008218f
C292 B.n255 VSUBS 0.008218f
C293 B.n256 VSUBS 0.008218f
C294 B.n257 VSUBS 0.008218f
C295 B.n258 VSUBS 0.008218f
C296 B.n259 VSUBS 0.008218f
C297 B.n260 VSUBS 0.008218f
C298 B.n261 VSUBS 0.008218f
C299 B.n262 VSUBS 0.008218f
C300 B.n263 VSUBS 0.008218f
C301 B.n264 VSUBS 0.008218f
C302 B.n265 VSUBS 0.008218f
C303 B.n266 VSUBS 0.008218f
C304 B.n267 VSUBS 0.008218f
C305 B.n268 VSUBS 0.008218f
C306 B.n269 VSUBS 0.008218f
C307 B.n270 VSUBS 0.008218f
C308 B.n271 VSUBS 0.008218f
C309 B.n272 VSUBS 0.008218f
C310 B.n273 VSUBS 0.008218f
C311 B.n274 VSUBS 0.008218f
C312 B.n275 VSUBS 0.008218f
C313 B.n276 VSUBS 0.008218f
C314 B.n277 VSUBS 0.008218f
C315 B.n278 VSUBS 0.008218f
C316 B.n279 VSUBS 0.018784f
C317 B.n280 VSUBS 0.019888f
C318 B.n281 VSUBS 0.019888f
C319 B.n282 VSUBS 0.008218f
C320 B.n283 VSUBS 0.008218f
C321 B.n284 VSUBS 0.008218f
C322 B.n285 VSUBS 0.008218f
C323 B.n286 VSUBS 0.008218f
C324 B.n287 VSUBS 0.008218f
C325 B.n288 VSUBS 0.008218f
C326 B.n289 VSUBS 0.008218f
C327 B.n290 VSUBS 0.008218f
C328 B.n291 VSUBS 0.008218f
C329 B.n292 VSUBS 0.008218f
C330 B.n293 VSUBS 0.008218f
C331 B.n294 VSUBS 0.008218f
C332 B.n295 VSUBS 0.008218f
C333 B.n296 VSUBS 0.008218f
C334 B.n297 VSUBS 0.008218f
C335 B.n298 VSUBS 0.008218f
C336 B.n299 VSUBS 0.008218f
C337 B.n300 VSUBS 0.008218f
C338 B.n301 VSUBS 0.008218f
C339 B.n302 VSUBS 0.008218f
C340 B.n303 VSUBS 0.008218f
C341 B.n304 VSUBS 0.008218f
C342 B.n305 VSUBS 0.008218f
C343 B.n306 VSUBS 0.008218f
C344 B.n307 VSUBS 0.008218f
C345 B.n308 VSUBS 0.008218f
C346 B.n309 VSUBS 0.008218f
C347 B.n310 VSUBS 0.008218f
C348 B.n311 VSUBS 0.008218f
C349 B.n312 VSUBS 0.008218f
C350 B.n313 VSUBS 0.008218f
C351 B.n314 VSUBS 0.008218f
C352 B.n315 VSUBS 0.008218f
C353 B.n316 VSUBS 0.008218f
C354 B.n317 VSUBS 0.008218f
C355 B.n318 VSUBS 0.008218f
C356 B.n319 VSUBS 0.008218f
C357 B.n320 VSUBS 0.008218f
C358 B.n321 VSUBS 0.008218f
C359 B.n322 VSUBS 0.008218f
C360 B.n323 VSUBS 0.008218f
C361 B.n324 VSUBS 0.008218f
C362 B.n325 VSUBS 0.008218f
C363 B.n326 VSUBS 0.008218f
C364 B.n327 VSUBS 0.008218f
C365 B.n328 VSUBS 0.008218f
C366 B.n329 VSUBS 0.008218f
C367 B.n330 VSUBS 0.008218f
C368 B.n331 VSUBS 0.008218f
C369 B.n332 VSUBS 0.008218f
C370 B.n333 VSUBS 0.008218f
C371 B.n334 VSUBS 0.008218f
C372 B.n335 VSUBS 0.008218f
C373 B.n336 VSUBS 0.008218f
C374 B.n337 VSUBS 0.008218f
C375 B.n338 VSUBS 0.008218f
C376 B.n339 VSUBS 0.008218f
C377 B.n340 VSUBS 0.008218f
C378 B.n341 VSUBS 0.008218f
C379 B.n342 VSUBS 0.008218f
C380 B.n343 VSUBS 0.008218f
C381 B.n344 VSUBS 0.008218f
C382 B.n345 VSUBS 0.008218f
C383 B.n346 VSUBS 0.008218f
C384 B.n347 VSUBS 0.008218f
C385 B.n348 VSUBS 0.008218f
C386 B.n349 VSUBS 0.008218f
C387 B.n350 VSUBS 0.007734f
C388 B.n351 VSUBS 0.01904f
C389 B.n352 VSUBS 0.004592f
C390 B.n353 VSUBS 0.008218f
C391 B.n354 VSUBS 0.008218f
C392 B.n355 VSUBS 0.008218f
C393 B.n356 VSUBS 0.008218f
C394 B.n357 VSUBS 0.008218f
C395 B.n358 VSUBS 0.008218f
C396 B.n359 VSUBS 0.008218f
C397 B.n360 VSUBS 0.008218f
C398 B.n361 VSUBS 0.008218f
C399 B.n362 VSUBS 0.008218f
C400 B.n363 VSUBS 0.008218f
C401 B.n364 VSUBS 0.008218f
C402 B.t8 VSUBS 0.539178f
C403 B.t7 VSUBS 0.56719f
C404 B.t6 VSUBS 2.31687f
C405 B.n365 VSUBS 0.316765f
C406 B.n366 VSUBS 0.086908f
C407 B.n367 VSUBS 0.01904f
C408 B.n368 VSUBS 0.004592f
C409 B.n369 VSUBS 0.008218f
C410 B.n370 VSUBS 0.008218f
C411 B.n371 VSUBS 0.008218f
C412 B.n372 VSUBS 0.008218f
C413 B.n373 VSUBS 0.008218f
C414 B.n374 VSUBS 0.008218f
C415 B.n375 VSUBS 0.008218f
C416 B.n376 VSUBS 0.008218f
C417 B.n377 VSUBS 0.008218f
C418 B.n378 VSUBS 0.008218f
C419 B.n379 VSUBS 0.008218f
C420 B.n380 VSUBS 0.008218f
C421 B.n381 VSUBS 0.008218f
C422 B.n382 VSUBS 0.008218f
C423 B.n383 VSUBS 0.008218f
C424 B.n384 VSUBS 0.008218f
C425 B.n385 VSUBS 0.008218f
C426 B.n386 VSUBS 0.008218f
C427 B.n387 VSUBS 0.008218f
C428 B.n388 VSUBS 0.008218f
C429 B.n389 VSUBS 0.008218f
C430 B.n390 VSUBS 0.008218f
C431 B.n391 VSUBS 0.008218f
C432 B.n392 VSUBS 0.008218f
C433 B.n393 VSUBS 0.008218f
C434 B.n394 VSUBS 0.008218f
C435 B.n395 VSUBS 0.008218f
C436 B.n396 VSUBS 0.008218f
C437 B.n397 VSUBS 0.008218f
C438 B.n398 VSUBS 0.008218f
C439 B.n399 VSUBS 0.008218f
C440 B.n400 VSUBS 0.008218f
C441 B.n401 VSUBS 0.008218f
C442 B.n402 VSUBS 0.008218f
C443 B.n403 VSUBS 0.008218f
C444 B.n404 VSUBS 0.008218f
C445 B.n405 VSUBS 0.008218f
C446 B.n406 VSUBS 0.008218f
C447 B.n407 VSUBS 0.008218f
C448 B.n408 VSUBS 0.008218f
C449 B.n409 VSUBS 0.008218f
C450 B.n410 VSUBS 0.008218f
C451 B.n411 VSUBS 0.008218f
C452 B.n412 VSUBS 0.008218f
C453 B.n413 VSUBS 0.008218f
C454 B.n414 VSUBS 0.008218f
C455 B.n415 VSUBS 0.008218f
C456 B.n416 VSUBS 0.008218f
C457 B.n417 VSUBS 0.008218f
C458 B.n418 VSUBS 0.008218f
C459 B.n419 VSUBS 0.008218f
C460 B.n420 VSUBS 0.008218f
C461 B.n421 VSUBS 0.008218f
C462 B.n422 VSUBS 0.008218f
C463 B.n423 VSUBS 0.008218f
C464 B.n424 VSUBS 0.008218f
C465 B.n425 VSUBS 0.008218f
C466 B.n426 VSUBS 0.008218f
C467 B.n427 VSUBS 0.008218f
C468 B.n428 VSUBS 0.008218f
C469 B.n429 VSUBS 0.008218f
C470 B.n430 VSUBS 0.008218f
C471 B.n431 VSUBS 0.008218f
C472 B.n432 VSUBS 0.008218f
C473 B.n433 VSUBS 0.008218f
C474 B.n434 VSUBS 0.008218f
C475 B.n435 VSUBS 0.008218f
C476 B.n436 VSUBS 0.008218f
C477 B.n437 VSUBS 0.008218f
C478 B.n438 VSUBS 0.008218f
C479 B.n439 VSUBS 0.018925f
C480 B.n440 VSUBS 0.019747f
C481 B.n441 VSUBS 0.018784f
C482 B.n442 VSUBS 0.008218f
C483 B.n443 VSUBS 0.008218f
C484 B.n444 VSUBS 0.008218f
C485 B.n445 VSUBS 0.008218f
C486 B.n446 VSUBS 0.008218f
C487 B.n447 VSUBS 0.008218f
C488 B.n448 VSUBS 0.008218f
C489 B.n449 VSUBS 0.008218f
C490 B.n450 VSUBS 0.008218f
C491 B.n451 VSUBS 0.008218f
C492 B.n452 VSUBS 0.008218f
C493 B.n453 VSUBS 0.008218f
C494 B.n454 VSUBS 0.008218f
C495 B.n455 VSUBS 0.008218f
C496 B.n456 VSUBS 0.008218f
C497 B.n457 VSUBS 0.008218f
C498 B.n458 VSUBS 0.008218f
C499 B.n459 VSUBS 0.008218f
C500 B.n460 VSUBS 0.008218f
C501 B.n461 VSUBS 0.008218f
C502 B.n462 VSUBS 0.008218f
C503 B.n463 VSUBS 0.008218f
C504 B.n464 VSUBS 0.008218f
C505 B.n465 VSUBS 0.008218f
C506 B.n466 VSUBS 0.008218f
C507 B.n467 VSUBS 0.008218f
C508 B.n468 VSUBS 0.008218f
C509 B.n469 VSUBS 0.008218f
C510 B.n470 VSUBS 0.008218f
C511 B.n471 VSUBS 0.008218f
C512 B.n472 VSUBS 0.008218f
C513 B.n473 VSUBS 0.008218f
C514 B.n474 VSUBS 0.008218f
C515 B.n475 VSUBS 0.008218f
C516 B.n476 VSUBS 0.008218f
C517 B.n477 VSUBS 0.008218f
C518 B.n478 VSUBS 0.008218f
C519 B.n479 VSUBS 0.008218f
C520 B.n480 VSUBS 0.008218f
C521 B.n481 VSUBS 0.008218f
C522 B.n482 VSUBS 0.008218f
C523 B.n483 VSUBS 0.008218f
C524 B.n484 VSUBS 0.008218f
C525 B.n485 VSUBS 0.008218f
C526 B.n486 VSUBS 0.008218f
C527 B.n487 VSUBS 0.008218f
C528 B.n488 VSUBS 0.008218f
C529 B.n489 VSUBS 0.008218f
C530 B.n490 VSUBS 0.008218f
C531 B.n491 VSUBS 0.008218f
C532 B.n492 VSUBS 0.008218f
C533 B.n493 VSUBS 0.008218f
C534 B.n494 VSUBS 0.008218f
C535 B.n495 VSUBS 0.008218f
C536 B.n496 VSUBS 0.008218f
C537 B.n497 VSUBS 0.008218f
C538 B.n498 VSUBS 0.008218f
C539 B.n499 VSUBS 0.008218f
C540 B.n500 VSUBS 0.008218f
C541 B.n501 VSUBS 0.008218f
C542 B.n502 VSUBS 0.008218f
C543 B.n503 VSUBS 0.008218f
C544 B.n504 VSUBS 0.008218f
C545 B.n505 VSUBS 0.008218f
C546 B.n506 VSUBS 0.008218f
C547 B.n507 VSUBS 0.008218f
C548 B.n508 VSUBS 0.008218f
C549 B.n509 VSUBS 0.008218f
C550 B.n510 VSUBS 0.008218f
C551 B.n511 VSUBS 0.008218f
C552 B.n512 VSUBS 0.008218f
C553 B.n513 VSUBS 0.008218f
C554 B.n514 VSUBS 0.008218f
C555 B.n515 VSUBS 0.008218f
C556 B.n516 VSUBS 0.008218f
C557 B.n517 VSUBS 0.008218f
C558 B.n518 VSUBS 0.008218f
C559 B.n519 VSUBS 0.008218f
C560 B.n520 VSUBS 0.008218f
C561 B.n521 VSUBS 0.008218f
C562 B.n522 VSUBS 0.008218f
C563 B.n523 VSUBS 0.008218f
C564 B.n524 VSUBS 0.008218f
C565 B.n525 VSUBS 0.008218f
C566 B.n526 VSUBS 0.008218f
C567 B.n527 VSUBS 0.008218f
C568 B.n528 VSUBS 0.008218f
C569 B.n529 VSUBS 0.008218f
C570 B.n530 VSUBS 0.008218f
C571 B.n531 VSUBS 0.008218f
C572 B.n532 VSUBS 0.008218f
C573 B.n533 VSUBS 0.008218f
C574 B.n534 VSUBS 0.008218f
C575 B.n535 VSUBS 0.008218f
C576 B.n536 VSUBS 0.008218f
C577 B.n537 VSUBS 0.008218f
C578 B.n538 VSUBS 0.008218f
C579 B.n539 VSUBS 0.008218f
C580 B.n540 VSUBS 0.008218f
C581 B.n541 VSUBS 0.008218f
C582 B.n542 VSUBS 0.008218f
C583 B.n543 VSUBS 0.008218f
C584 B.n544 VSUBS 0.008218f
C585 B.n545 VSUBS 0.008218f
C586 B.n546 VSUBS 0.008218f
C587 B.n547 VSUBS 0.008218f
C588 B.n548 VSUBS 0.008218f
C589 B.n549 VSUBS 0.008218f
C590 B.n550 VSUBS 0.008218f
C591 B.n551 VSUBS 0.008218f
C592 B.n552 VSUBS 0.008218f
C593 B.n553 VSUBS 0.008218f
C594 B.n554 VSUBS 0.008218f
C595 B.n555 VSUBS 0.008218f
C596 B.n556 VSUBS 0.008218f
C597 B.n557 VSUBS 0.008218f
C598 B.n558 VSUBS 0.008218f
C599 B.n559 VSUBS 0.008218f
C600 B.n560 VSUBS 0.008218f
C601 B.n561 VSUBS 0.008218f
C602 B.n562 VSUBS 0.008218f
C603 B.n563 VSUBS 0.008218f
C604 B.n564 VSUBS 0.008218f
C605 B.n565 VSUBS 0.008218f
C606 B.n566 VSUBS 0.008218f
C607 B.n567 VSUBS 0.008218f
C608 B.n568 VSUBS 0.008218f
C609 B.n569 VSUBS 0.008218f
C610 B.n570 VSUBS 0.008218f
C611 B.n571 VSUBS 0.008218f
C612 B.n572 VSUBS 0.008218f
C613 B.n573 VSUBS 0.008218f
C614 B.n574 VSUBS 0.008218f
C615 B.n575 VSUBS 0.008218f
C616 B.n576 VSUBS 0.008218f
C617 B.n577 VSUBS 0.008218f
C618 B.n578 VSUBS 0.008218f
C619 B.n579 VSUBS 0.008218f
C620 B.n580 VSUBS 0.008218f
C621 B.n581 VSUBS 0.008218f
C622 B.n582 VSUBS 0.008218f
C623 B.n583 VSUBS 0.008218f
C624 B.n584 VSUBS 0.008218f
C625 B.n585 VSUBS 0.008218f
C626 B.n586 VSUBS 0.018784f
C627 B.n587 VSUBS 0.019888f
C628 B.n588 VSUBS 0.019888f
C629 B.n589 VSUBS 0.008218f
C630 B.n590 VSUBS 0.008218f
C631 B.n591 VSUBS 0.008218f
C632 B.n592 VSUBS 0.008218f
C633 B.n593 VSUBS 0.008218f
C634 B.n594 VSUBS 0.008218f
C635 B.n595 VSUBS 0.008218f
C636 B.n596 VSUBS 0.008218f
C637 B.n597 VSUBS 0.008218f
C638 B.n598 VSUBS 0.008218f
C639 B.n599 VSUBS 0.008218f
C640 B.n600 VSUBS 0.008218f
C641 B.n601 VSUBS 0.008218f
C642 B.n602 VSUBS 0.008218f
C643 B.n603 VSUBS 0.008218f
C644 B.n604 VSUBS 0.008218f
C645 B.n605 VSUBS 0.008218f
C646 B.n606 VSUBS 0.008218f
C647 B.n607 VSUBS 0.008218f
C648 B.n608 VSUBS 0.008218f
C649 B.n609 VSUBS 0.008218f
C650 B.n610 VSUBS 0.008218f
C651 B.n611 VSUBS 0.008218f
C652 B.n612 VSUBS 0.008218f
C653 B.n613 VSUBS 0.008218f
C654 B.n614 VSUBS 0.008218f
C655 B.n615 VSUBS 0.008218f
C656 B.n616 VSUBS 0.008218f
C657 B.n617 VSUBS 0.008218f
C658 B.n618 VSUBS 0.008218f
C659 B.n619 VSUBS 0.008218f
C660 B.n620 VSUBS 0.008218f
C661 B.n621 VSUBS 0.008218f
C662 B.n622 VSUBS 0.008218f
C663 B.n623 VSUBS 0.008218f
C664 B.n624 VSUBS 0.008218f
C665 B.n625 VSUBS 0.008218f
C666 B.n626 VSUBS 0.008218f
C667 B.n627 VSUBS 0.008218f
C668 B.n628 VSUBS 0.008218f
C669 B.n629 VSUBS 0.008218f
C670 B.n630 VSUBS 0.008218f
C671 B.n631 VSUBS 0.008218f
C672 B.n632 VSUBS 0.008218f
C673 B.n633 VSUBS 0.008218f
C674 B.n634 VSUBS 0.008218f
C675 B.n635 VSUBS 0.008218f
C676 B.n636 VSUBS 0.008218f
C677 B.n637 VSUBS 0.008218f
C678 B.n638 VSUBS 0.008218f
C679 B.n639 VSUBS 0.008218f
C680 B.n640 VSUBS 0.008218f
C681 B.n641 VSUBS 0.008218f
C682 B.n642 VSUBS 0.008218f
C683 B.n643 VSUBS 0.008218f
C684 B.n644 VSUBS 0.008218f
C685 B.n645 VSUBS 0.008218f
C686 B.n646 VSUBS 0.008218f
C687 B.n647 VSUBS 0.008218f
C688 B.n648 VSUBS 0.008218f
C689 B.n649 VSUBS 0.008218f
C690 B.n650 VSUBS 0.008218f
C691 B.n651 VSUBS 0.008218f
C692 B.n652 VSUBS 0.008218f
C693 B.n653 VSUBS 0.008218f
C694 B.n654 VSUBS 0.008218f
C695 B.n655 VSUBS 0.008218f
C696 B.n656 VSUBS 0.007734f
C697 B.n657 VSUBS 0.008218f
C698 B.n658 VSUBS 0.008218f
C699 B.n659 VSUBS 0.008218f
C700 B.n660 VSUBS 0.008218f
C701 B.n661 VSUBS 0.008218f
C702 B.n662 VSUBS 0.008218f
C703 B.n663 VSUBS 0.008218f
C704 B.n664 VSUBS 0.008218f
C705 B.n665 VSUBS 0.008218f
C706 B.n666 VSUBS 0.008218f
C707 B.n667 VSUBS 0.008218f
C708 B.n668 VSUBS 0.008218f
C709 B.n669 VSUBS 0.008218f
C710 B.n670 VSUBS 0.008218f
C711 B.n671 VSUBS 0.008218f
C712 B.n672 VSUBS 0.004592f
C713 B.n673 VSUBS 0.01904f
C714 B.n674 VSUBS 0.007734f
C715 B.n675 VSUBS 0.008218f
C716 B.n676 VSUBS 0.008218f
C717 B.n677 VSUBS 0.008218f
C718 B.n678 VSUBS 0.008218f
C719 B.n679 VSUBS 0.008218f
C720 B.n680 VSUBS 0.008218f
C721 B.n681 VSUBS 0.008218f
C722 B.n682 VSUBS 0.008218f
C723 B.n683 VSUBS 0.008218f
C724 B.n684 VSUBS 0.008218f
C725 B.n685 VSUBS 0.008218f
C726 B.n686 VSUBS 0.008218f
C727 B.n687 VSUBS 0.008218f
C728 B.n688 VSUBS 0.008218f
C729 B.n689 VSUBS 0.008218f
C730 B.n690 VSUBS 0.008218f
C731 B.n691 VSUBS 0.008218f
C732 B.n692 VSUBS 0.008218f
C733 B.n693 VSUBS 0.008218f
C734 B.n694 VSUBS 0.008218f
C735 B.n695 VSUBS 0.008218f
C736 B.n696 VSUBS 0.008218f
C737 B.n697 VSUBS 0.008218f
C738 B.n698 VSUBS 0.008218f
C739 B.n699 VSUBS 0.008218f
C740 B.n700 VSUBS 0.008218f
C741 B.n701 VSUBS 0.008218f
C742 B.n702 VSUBS 0.008218f
C743 B.n703 VSUBS 0.008218f
C744 B.n704 VSUBS 0.008218f
C745 B.n705 VSUBS 0.008218f
C746 B.n706 VSUBS 0.008218f
C747 B.n707 VSUBS 0.008218f
C748 B.n708 VSUBS 0.008218f
C749 B.n709 VSUBS 0.008218f
C750 B.n710 VSUBS 0.008218f
C751 B.n711 VSUBS 0.008218f
C752 B.n712 VSUBS 0.008218f
C753 B.n713 VSUBS 0.008218f
C754 B.n714 VSUBS 0.008218f
C755 B.n715 VSUBS 0.008218f
C756 B.n716 VSUBS 0.008218f
C757 B.n717 VSUBS 0.008218f
C758 B.n718 VSUBS 0.008218f
C759 B.n719 VSUBS 0.008218f
C760 B.n720 VSUBS 0.008218f
C761 B.n721 VSUBS 0.008218f
C762 B.n722 VSUBS 0.008218f
C763 B.n723 VSUBS 0.008218f
C764 B.n724 VSUBS 0.008218f
C765 B.n725 VSUBS 0.008218f
C766 B.n726 VSUBS 0.008218f
C767 B.n727 VSUBS 0.008218f
C768 B.n728 VSUBS 0.008218f
C769 B.n729 VSUBS 0.008218f
C770 B.n730 VSUBS 0.008218f
C771 B.n731 VSUBS 0.008218f
C772 B.n732 VSUBS 0.008218f
C773 B.n733 VSUBS 0.008218f
C774 B.n734 VSUBS 0.008218f
C775 B.n735 VSUBS 0.008218f
C776 B.n736 VSUBS 0.008218f
C777 B.n737 VSUBS 0.008218f
C778 B.n738 VSUBS 0.008218f
C779 B.n739 VSUBS 0.008218f
C780 B.n740 VSUBS 0.008218f
C781 B.n741 VSUBS 0.008218f
C782 B.n742 VSUBS 0.008218f
C783 B.n743 VSUBS 0.019888f
C784 B.n744 VSUBS 0.018784f
C785 B.n745 VSUBS 0.018784f
C786 B.n746 VSUBS 0.008218f
C787 B.n747 VSUBS 0.008218f
C788 B.n748 VSUBS 0.008218f
C789 B.n749 VSUBS 0.008218f
C790 B.n750 VSUBS 0.008218f
C791 B.n751 VSUBS 0.008218f
C792 B.n752 VSUBS 0.008218f
C793 B.n753 VSUBS 0.008218f
C794 B.n754 VSUBS 0.008218f
C795 B.n755 VSUBS 0.008218f
C796 B.n756 VSUBS 0.008218f
C797 B.n757 VSUBS 0.008218f
C798 B.n758 VSUBS 0.008218f
C799 B.n759 VSUBS 0.008218f
C800 B.n760 VSUBS 0.008218f
C801 B.n761 VSUBS 0.008218f
C802 B.n762 VSUBS 0.008218f
C803 B.n763 VSUBS 0.008218f
C804 B.n764 VSUBS 0.008218f
C805 B.n765 VSUBS 0.008218f
C806 B.n766 VSUBS 0.008218f
C807 B.n767 VSUBS 0.008218f
C808 B.n768 VSUBS 0.008218f
C809 B.n769 VSUBS 0.008218f
C810 B.n770 VSUBS 0.008218f
C811 B.n771 VSUBS 0.008218f
C812 B.n772 VSUBS 0.008218f
C813 B.n773 VSUBS 0.008218f
C814 B.n774 VSUBS 0.008218f
C815 B.n775 VSUBS 0.008218f
C816 B.n776 VSUBS 0.008218f
C817 B.n777 VSUBS 0.008218f
C818 B.n778 VSUBS 0.008218f
C819 B.n779 VSUBS 0.008218f
C820 B.n780 VSUBS 0.008218f
C821 B.n781 VSUBS 0.008218f
C822 B.n782 VSUBS 0.008218f
C823 B.n783 VSUBS 0.008218f
C824 B.n784 VSUBS 0.008218f
C825 B.n785 VSUBS 0.008218f
C826 B.n786 VSUBS 0.008218f
C827 B.n787 VSUBS 0.008218f
C828 B.n788 VSUBS 0.008218f
C829 B.n789 VSUBS 0.008218f
C830 B.n790 VSUBS 0.008218f
C831 B.n791 VSUBS 0.008218f
C832 B.n792 VSUBS 0.008218f
C833 B.n793 VSUBS 0.008218f
C834 B.n794 VSUBS 0.008218f
C835 B.n795 VSUBS 0.008218f
C836 B.n796 VSUBS 0.008218f
C837 B.n797 VSUBS 0.008218f
C838 B.n798 VSUBS 0.008218f
C839 B.n799 VSUBS 0.008218f
C840 B.n800 VSUBS 0.008218f
C841 B.n801 VSUBS 0.008218f
C842 B.n802 VSUBS 0.008218f
C843 B.n803 VSUBS 0.008218f
C844 B.n804 VSUBS 0.008218f
C845 B.n805 VSUBS 0.008218f
C846 B.n806 VSUBS 0.008218f
C847 B.n807 VSUBS 0.008218f
C848 B.n808 VSUBS 0.008218f
C849 B.n809 VSUBS 0.008218f
C850 B.n810 VSUBS 0.008218f
C851 B.n811 VSUBS 0.008218f
C852 B.n812 VSUBS 0.008218f
C853 B.n813 VSUBS 0.008218f
C854 B.n814 VSUBS 0.008218f
C855 B.n815 VSUBS 0.010724f
C856 B.n816 VSUBS 0.011424f
C857 B.n817 VSUBS 0.022717f
C858 VDD1.t4 VSUBS 3.19694f
C859 VDD1.t0 VSUBS 3.19541f
C860 VDD1.t2 VSUBS 0.305013f
C861 VDD1.t3 VSUBS 0.305013f
C862 VDD1.n0 VSUBS 2.44194f
C863 VDD1.n1 VSUBS 4.392509f
C864 VDD1.t5 VSUBS 0.305013f
C865 VDD1.t1 VSUBS 0.305013f
C866 VDD1.n2 VSUBS 2.43358f
C867 VDD1.n3 VSUBS 3.73061f
C868 VP.t2 VSUBS 3.43099f
C869 VP.n0 VSUBS 1.32015f
C870 VP.n1 VSUBS 0.029038f
C871 VP.n2 VSUBS 0.039963f
C872 VP.n3 VSUBS 0.029038f
C873 VP.t3 VSUBS 3.43099f
C874 VP.n4 VSUBS 0.054119f
C875 VP.n5 VSUBS 0.029038f
C876 VP.n6 VSUBS 0.054119f
C877 VP.t4 VSUBS 3.43099f
C878 VP.n7 VSUBS 1.32015f
C879 VP.n8 VSUBS 0.029038f
C880 VP.n9 VSUBS 0.039963f
C881 VP.n10 VSUBS 0.330329f
C882 VP.t0 VSUBS 3.43099f
C883 VP.t1 VSUBS 3.76446f
C884 VP.n11 VSUBS 1.24387f
C885 VP.n12 VSUBS 1.308f
C886 VP.n13 VSUBS 0.054119f
C887 VP.n14 VSUBS 0.054119f
C888 VP.n15 VSUBS 0.029038f
C889 VP.n16 VSUBS 0.029038f
C890 VP.n17 VSUBS 0.029038f
C891 VP.n18 VSUBS 0.044818f
C892 VP.n19 VSUBS 0.054119f
C893 VP.n20 VSUBS 0.050913f
C894 VP.n21 VSUBS 0.046867f
C895 VP.n22 VSUBS 1.75017f
C896 VP.n23 VSUBS 1.77014f
C897 VP.t5 VSUBS 3.43099f
C898 VP.n24 VSUBS 1.32015f
C899 VP.n25 VSUBS 0.050913f
C900 VP.n26 VSUBS 0.046867f
C901 VP.n27 VSUBS 0.029038f
C902 VP.n28 VSUBS 0.029038f
C903 VP.n29 VSUBS 0.044818f
C904 VP.n30 VSUBS 0.039963f
C905 VP.n31 VSUBS 0.054119f
C906 VP.n32 VSUBS 0.029038f
C907 VP.n33 VSUBS 0.029038f
C908 VP.n34 VSUBS 0.029038f
C909 VP.n35 VSUBS 1.2259f
C910 VP.n36 VSUBS 0.054119f
C911 VP.n37 VSUBS 0.054119f
C912 VP.n38 VSUBS 0.029038f
C913 VP.n39 VSUBS 0.029038f
C914 VP.n40 VSUBS 0.029038f
C915 VP.n41 VSUBS 0.044818f
C916 VP.n42 VSUBS 0.054119f
C917 VP.n43 VSUBS 0.050913f
C918 VP.n44 VSUBS 0.046867f
C919 VP.n45 VSUBS 0.059314f
C920 VDD2.t5 VSUBS 3.2106f
C921 VDD2.t2 VSUBS 0.306463f
C922 VDD2.t0 VSUBS 0.306463f
C923 VDD2.n0 VSUBS 2.45354f
C924 VDD2.n1 VSUBS 4.25804f
C925 VDD2.t4 VSUBS 3.18651f
C926 VDD2.n2 VSUBS 3.77208f
C927 VDD2.t3 VSUBS 0.306463f
C928 VDD2.t1 VSUBS 0.306463f
C929 VDD2.n3 VSUBS 2.4535f
C930 VTAIL.t9 VSUBS 0.317655f
C931 VTAIL.t8 VSUBS 0.317655f
C932 VTAIL.n0 VSUBS 2.36479f
C933 VTAIL.n1 VSUBS 0.948689f
C934 VTAIL.t0 VSUBS 3.11155f
C935 VTAIL.n2 VSUBS 1.27024f
C936 VTAIL.t2 VSUBS 0.317655f
C937 VTAIL.t3 VSUBS 0.317655f
C938 VTAIL.n3 VSUBS 2.36479f
C939 VTAIL.n4 VSUBS 3.03138f
C940 VTAIL.t11 VSUBS 0.317655f
C941 VTAIL.t10 VSUBS 0.317655f
C942 VTAIL.n5 VSUBS 2.36479f
C943 VTAIL.n6 VSUBS 3.03138f
C944 VTAIL.t7 VSUBS 3.11157f
C945 VTAIL.n7 VSUBS 1.27022f
C946 VTAIL.t5 VSUBS 0.317655f
C947 VTAIL.t4 VSUBS 0.317655f
C948 VTAIL.n8 VSUBS 2.36479f
C949 VTAIL.n9 VSUBS 1.15066f
C950 VTAIL.t1 VSUBS 3.11157f
C951 VTAIL.n10 VSUBS 2.8744f
C952 VTAIL.t6 VSUBS 3.11155f
C953 VTAIL.n11 VSUBS 2.79985f
C954 VN.t5 VSUBS 3.13545f
C955 VN.n0 VSUBS 1.20644f
C956 VN.n1 VSUBS 0.026537f
C957 VN.n2 VSUBS 0.03652f
C958 VN.n3 VSUBS 0.301874f
C959 VN.t3 VSUBS 3.13545f
C960 VN.t0 VSUBS 3.4402f
C961 VN.n4 VSUBS 1.13672f
C962 VN.n5 VSUBS 1.19533f
C963 VN.n6 VSUBS 0.049458f
C964 VN.n7 VSUBS 0.049458f
C965 VN.n8 VSUBS 0.026537f
C966 VN.n9 VSUBS 0.026537f
C967 VN.n10 VSUBS 0.026537f
C968 VN.n11 VSUBS 0.040957f
C969 VN.n12 VSUBS 0.049458f
C970 VN.n13 VSUBS 0.046528f
C971 VN.n14 VSUBS 0.042829f
C972 VN.n15 VSUBS 0.054204f
C973 VN.t1 VSUBS 3.13545f
C974 VN.n16 VSUBS 1.20644f
C975 VN.n17 VSUBS 0.026537f
C976 VN.n18 VSUBS 0.03652f
C977 VN.n19 VSUBS 0.301874f
C978 VN.t2 VSUBS 3.13545f
C979 VN.t4 VSUBS 3.4402f
C980 VN.n20 VSUBS 1.13672f
C981 VN.n21 VSUBS 1.19533f
C982 VN.n22 VSUBS 0.049458f
C983 VN.n23 VSUBS 0.049458f
C984 VN.n24 VSUBS 0.026537f
C985 VN.n25 VSUBS 0.026537f
C986 VN.n26 VSUBS 0.026537f
C987 VN.n27 VSUBS 0.040957f
C988 VN.n28 VSUBS 0.049458f
C989 VN.n29 VSUBS 0.046528f
C990 VN.n30 VSUBS 0.042829f
C991 VN.n31 VSUBS 1.6101f
.ends

