* NGSPICE file created from diff_pair_sample_0396.ext - technology: sky130A

.subckt diff_pair_sample_0396 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=1.59
X1 VTAIL.t15 VN.t0 VDD2.t0 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=1.59
X2 VTAIL.t14 VN.t1 VDD2.t5 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=1.59
X3 VDD2.t1 VN.t2 VTAIL.t13 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=1.59
X4 VTAIL.t12 VN.t3 VDD2.t2 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X5 VDD2.t7 VN.t4 VTAIL.t11 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X6 VDD1.t7 VP.t0 VTAIL.t3 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X7 VDD1.t6 VP.t1 VTAIL.t7 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=1.59
X8 VDD2.t6 VN.t5 VTAIL.t10 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=1.59
X9 VTAIL.t5 VP.t2 VDD1.t5 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X10 VDD1.t4 VP.t3 VTAIL.t4 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X11 VTAIL.t6 VP.t4 VDD1.t3 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=1.59
X12 B.t8 B.t6 B.t7 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=1.59
X13 B.t5 B.t3 B.t4 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=1.59
X14 VTAIL.t2 VP.t5 VDD1.t2 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X15 B.t2 B.t0 B.t1 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=1.59
X16 VTAIL.t9 VN.t6 VDD2.t3 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
X17 VDD1.t1 VP.t6 VTAIL.t1 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=1.59
X18 VTAIL.t0 VP.t7 VDD1.t0 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=1.59
X19 VDD2.t4 VN.t7 VTAIL.t8 w_n2890_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=1.59
R0 B.n259 B.n86 585
R1 B.n258 B.n257 585
R2 B.n256 B.n87 585
R3 B.n255 B.n254 585
R4 B.n253 B.n88 585
R5 B.n252 B.n251 585
R6 B.n250 B.n89 585
R7 B.n249 B.n248 585
R8 B.n247 B.n90 585
R9 B.n246 B.n245 585
R10 B.n244 B.n91 585
R11 B.n243 B.n242 585
R12 B.n241 B.n92 585
R13 B.n240 B.n239 585
R14 B.n238 B.n93 585
R15 B.n237 B.n236 585
R16 B.n235 B.n94 585
R17 B.n234 B.n233 585
R18 B.n232 B.n95 585
R19 B.n231 B.n230 585
R20 B.n229 B.n228 585
R21 B.n227 B.n99 585
R22 B.n226 B.n225 585
R23 B.n224 B.n100 585
R24 B.n223 B.n222 585
R25 B.n221 B.n101 585
R26 B.n220 B.n219 585
R27 B.n218 B.n102 585
R28 B.n217 B.n216 585
R29 B.n214 B.n103 585
R30 B.n213 B.n212 585
R31 B.n211 B.n106 585
R32 B.n210 B.n209 585
R33 B.n208 B.n107 585
R34 B.n207 B.n206 585
R35 B.n205 B.n108 585
R36 B.n204 B.n203 585
R37 B.n202 B.n109 585
R38 B.n201 B.n200 585
R39 B.n199 B.n110 585
R40 B.n198 B.n197 585
R41 B.n196 B.n111 585
R42 B.n195 B.n194 585
R43 B.n193 B.n112 585
R44 B.n192 B.n191 585
R45 B.n190 B.n113 585
R46 B.n189 B.n188 585
R47 B.n187 B.n114 585
R48 B.n186 B.n185 585
R49 B.n261 B.n260 585
R50 B.n262 B.n85 585
R51 B.n264 B.n263 585
R52 B.n265 B.n84 585
R53 B.n267 B.n266 585
R54 B.n268 B.n83 585
R55 B.n270 B.n269 585
R56 B.n271 B.n82 585
R57 B.n273 B.n272 585
R58 B.n274 B.n81 585
R59 B.n276 B.n275 585
R60 B.n277 B.n80 585
R61 B.n279 B.n278 585
R62 B.n280 B.n79 585
R63 B.n282 B.n281 585
R64 B.n283 B.n78 585
R65 B.n285 B.n284 585
R66 B.n286 B.n77 585
R67 B.n288 B.n287 585
R68 B.n289 B.n76 585
R69 B.n291 B.n290 585
R70 B.n292 B.n75 585
R71 B.n294 B.n293 585
R72 B.n295 B.n74 585
R73 B.n297 B.n296 585
R74 B.n298 B.n73 585
R75 B.n300 B.n299 585
R76 B.n301 B.n72 585
R77 B.n303 B.n302 585
R78 B.n304 B.n71 585
R79 B.n306 B.n305 585
R80 B.n307 B.n70 585
R81 B.n309 B.n308 585
R82 B.n310 B.n69 585
R83 B.n312 B.n311 585
R84 B.n313 B.n68 585
R85 B.n315 B.n314 585
R86 B.n316 B.n67 585
R87 B.n318 B.n317 585
R88 B.n319 B.n66 585
R89 B.n321 B.n320 585
R90 B.n322 B.n65 585
R91 B.n324 B.n323 585
R92 B.n325 B.n64 585
R93 B.n327 B.n326 585
R94 B.n328 B.n63 585
R95 B.n330 B.n329 585
R96 B.n331 B.n62 585
R97 B.n333 B.n332 585
R98 B.n334 B.n61 585
R99 B.n336 B.n335 585
R100 B.n337 B.n60 585
R101 B.n339 B.n338 585
R102 B.n340 B.n59 585
R103 B.n342 B.n341 585
R104 B.n343 B.n58 585
R105 B.n345 B.n344 585
R106 B.n346 B.n57 585
R107 B.n348 B.n347 585
R108 B.n349 B.n56 585
R109 B.n351 B.n350 585
R110 B.n352 B.n55 585
R111 B.n354 B.n353 585
R112 B.n355 B.n54 585
R113 B.n357 B.n356 585
R114 B.n358 B.n53 585
R115 B.n360 B.n359 585
R116 B.n361 B.n52 585
R117 B.n363 B.n362 585
R118 B.n364 B.n51 585
R119 B.n366 B.n365 585
R120 B.n367 B.n50 585
R121 B.n369 B.n368 585
R122 B.n370 B.n49 585
R123 B.n445 B.n20 585
R124 B.n444 B.n443 585
R125 B.n442 B.n21 585
R126 B.n441 B.n440 585
R127 B.n439 B.n22 585
R128 B.n438 B.n437 585
R129 B.n436 B.n23 585
R130 B.n435 B.n434 585
R131 B.n433 B.n24 585
R132 B.n432 B.n431 585
R133 B.n430 B.n25 585
R134 B.n429 B.n428 585
R135 B.n427 B.n26 585
R136 B.n426 B.n425 585
R137 B.n424 B.n27 585
R138 B.n423 B.n422 585
R139 B.n421 B.n28 585
R140 B.n420 B.n419 585
R141 B.n418 B.n29 585
R142 B.n417 B.n416 585
R143 B.n415 B.n414 585
R144 B.n413 B.n33 585
R145 B.n412 B.n411 585
R146 B.n410 B.n34 585
R147 B.n409 B.n408 585
R148 B.n407 B.n35 585
R149 B.n406 B.n405 585
R150 B.n404 B.n36 585
R151 B.n403 B.n402 585
R152 B.n400 B.n37 585
R153 B.n399 B.n398 585
R154 B.n397 B.n40 585
R155 B.n396 B.n395 585
R156 B.n394 B.n41 585
R157 B.n393 B.n392 585
R158 B.n391 B.n42 585
R159 B.n390 B.n389 585
R160 B.n388 B.n43 585
R161 B.n387 B.n386 585
R162 B.n385 B.n44 585
R163 B.n384 B.n383 585
R164 B.n382 B.n45 585
R165 B.n381 B.n380 585
R166 B.n379 B.n46 585
R167 B.n378 B.n377 585
R168 B.n376 B.n47 585
R169 B.n375 B.n374 585
R170 B.n373 B.n48 585
R171 B.n372 B.n371 585
R172 B.n447 B.n446 585
R173 B.n448 B.n19 585
R174 B.n450 B.n449 585
R175 B.n451 B.n18 585
R176 B.n453 B.n452 585
R177 B.n454 B.n17 585
R178 B.n456 B.n455 585
R179 B.n457 B.n16 585
R180 B.n459 B.n458 585
R181 B.n460 B.n15 585
R182 B.n462 B.n461 585
R183 B.n463 B.n14 585
R184 B.n465 B.n464 585
R185 B.n466 B.n13 585
R186 B.n468 B.n467 585
R187 B.n469 B.n12 585
R188 B.n471 B.n470 585
R189 B.n472 B.n11 585
R190 B.n474 B.n473 585
R191 B.n475 B.n10 585
R192 B.n477 B.n476 585
R193 B.n478 B.n9 585
R194 B.n480 B.n479 585
R195 B.n481 B.n8 585
R196 B.n483 B.n482 585
R197 B.n484 B.n7 585
R198 B.n486 B.n485 585
R199 B.n487 B.n6 585
R200 B.n489 B.n488 585
R201 B.n490 B.n5 585
R202 B.n492 B.n491 585
R203 B.n493 B.n4 585
R204 B.n495 B.n494 585
R205 B.n496 B.n3 585
R206 B.n498 B.n497 585
R207 B.n499 B.n0 585
R208 B.n2 B.n1 585
R209 B.n133 B.n132 585
R210 B.n135 B.n134 585
R211 B.n136 B.n131 585
R212 B.n138 B.n137 585
R213 B.n139 B.n130 585
R214 B.n141 B.n140 585
R215 B.n142 B.n129 585
R216 B.n144 B.n143 585
R217 B.n145 B.n128 585
R218 B.n147 B.n146 585
R219 B.n148 B.n127 585
R220 B.n150 B.n149 585
R221 B.n151 B.n126 585
R222 B.n153 B.n152 585
R223 B.n154 B.n125 585
R224 B.n156 B.n155 585
R225 B.n157 B.n124 585
R226 B.n159 B.n158 585
R227 B.n160 B.n123 585
R228 B.n162 B.n161 585
R229 B.n163 B.n122 585
R230 B.n165 B.n164 585
R231 B.n166 B.n121 585
R232 B.n168 B.n167 585
R233 B.n169 B.n120 585
R234 B.n171 B.n170 585
R235 B.n172 B.n119 585
R236 B.n174 B.n173 585
R237 B.n175 B.n118 585
R238 B.n177 B.n176 585
R239 B.n178 B.n117 585
R240 B.n180 B.n179 585
R241 B.n181 B.n116 585
R242 B.n183 B.n182 585
R243 B.n184 B.n115 585
R244 B.n186 B.n115 439.647
R245 B.n260 B.n259 439.647
R246 B.n372 B.n49 439.647
R247 B.n446 B.n445 439.647
R248 B.n96 B.t10 279.253
R249 B.n38 B.t8 279.253
R250 B.n104 B.t4 279.253
R251 B.n30 B.t2 279.253
R252 B.n104 B.t3 273.664
R253 B.n96 B.t9 273.664
R254 B.n38 B.t6 273.664
R255 B.n30 B.t0 273.664
R256 B.n501 B.n500 256.663
R257 B.n97 B.t11 242.018
R258 B.n39 B.t7 242.018
R259 B.n105 B.t5 242.018
R260 B.n31 B.t1 242.018
R261 B.n500 B.n499 235.042
R262 B.n500 B.n2 235.042
R263 B.n187 B.n186 163.367
R264 B.n188 B.n187 163.367
R265 B.n188 B.n113 163.367
R266 B.n192 B.n113 163.367
R267 B.n193 B.n192 163.367
R268 B.n194 B.n193 163.367
R269 B.n194 B.n111 163.367
R270 B.n198 B.n111 163.367
R271 B.n199 B.n198 163.367
R272 B.n200 B.n199 163.367
R273 B.n200 B.n109 163.367
R274 B.n204 B.n109 163.367
R275 B.n205 B.n204 163.367
R276 B.n206 B.n205 163.367
R277 B.n206 B.n107 163.367
R278 B.n210 B.n107 163.367
R279 B.n211 B.n210 163.367
R280 B.n212 B.n211 163.367
R281 B.n212 B.n103 163.367
R282 B.n217 B.n103 163.367
R283 B.n218 B.n217 163.367
R284 B.n219 B.n218 163.367
R285 B.n219 B.n101 163.367
R286 B.n223 B.n101 163.367
R287 B.n224 B.n223 163.367
R288 B.n225 B.n224 163.367
R289 B.n225 B.n99 163.367
R290 B.n229 B.n99 163.367
R291 B.n230 B.n229 163.367
R292 B.n230 B.n95 163.367
R293 B.n234 B.n95 163.367
R294 B.n235 B.n234 163.367
R295 B.n236 B.n235 163.367
R296 B.n236 B.n93 163.367
R297 B.n240 B.n93 163.367
R298 B.n241 B.n240 163.367
R299 B.n242 B.n241 163.367
R300 B.n242 B.n91 163.367
R301 B.n246 B.n91 163.367
R302 B.n247 B.n246 163.367
R303 B.n248 B.n247 163.367
R304 B.n248 B.n89 163.367
R305 B.n252 B.n89 163.367
R306 B.n253 B.n252 163.367
R307 B.n254 B.n253 163.367
R308 B.n254 B.n87 163.367
R309 B.n258 B.n87 163.367
R310 B.n259 B.n258 163.367
R311 B.n368 B.n49 163.367
R312 B.n368 B.n367 163.367
R313 B.n367 B.n366 163.367
R314 B.n366 B.n51 163.367
R315 B.n362 B.n51 163.367
R316 B.n362 B.n361 163.367
R317 B.n361 B.n360 163.367
R318 B.n360 B.n53 163.367
R319 B.n356 B.n53 163.367
R320 B.n356 B.n355 163.367
R321 B.n355 B.n354 163.367
R322 B.n354 B.n55 163.367
R323 B.n350 B.n55 163.367
R324 B.n350 B.n349 163.367
R325 B.n349 B.n348 163.367
R326 B.n348 B.n57 163.367
R327 B.n344 B.n57 163.367
R328 B.n344 B.n343 163.367
R329 B.n343 B.n342 163.367
R330 B.n342 B.n59 163.367
R331 B.n338 B.n59 163.367
R332 B.n338 B.n337 163.367
R333 B.n337 B.n336 163.367
R334 B.n336 B.n61 163.367
R335 B.n332 B.n61 163.367
R336 B.n332 B.n331 163.367
R337 B.n331 B.n330 163.367
R338 B.n330 B.n63 163.367
R339 B.n326 B.n63 163.367
R340 B.n326 B.n325 163.367
R341 B.n325 B.n324 163.367
R342 B.n324 B.n65 163.367
R343 B.n320 B.n65 163.367
R344 B.n320 B.n319 163.367
R345 B.n319 B.n318 163.367
R346 B.n318 B.n67 163.367
R347 B.n314 B.n67 163.367
R348 B.n314 B.n313 163.367
R349 B.n313 B.n312 163.367
R350 B.n312 B.n69 163.367
R351 B.n308 B.n69 163.367
R352 B.n308 B.n307 163.367
R353 B.n307 B.n306 163.367
R354 B.n306 B.n71 163.367
R355 B.n302 B.n71 163.367
R356 B.n302 B.n301 163.367
R357 B.n301 B.n300 163.367
R358 B.n300 B.n73 163.367
R359 B.n296 B.n73 163.367
R360 B.n296 B.n295 163.367
R361 B.n295 B.n294 163.367
R362 B.n294 B.n75 163.367
R363 B.n290 B.n75 163.367
R364 B.n290 B.n289 163.367
R365 B.n289 B.n288 163.367
R366 B.n288 B.n77 163.367
R367 B.n284 B.n77 163.367
R368 B.n284 B.n283 163.367
R369 B.n283 B.n282 163.367
R370 B.n282 B.n79 163.367
R371 B.n278 B.n79 163.367
R372 B.n278 B.n277 163.367
R373 B.n277 B.n276 163.367
R374 B.n276 B.n81 163.367
R375 B.n272 B.n81 163.367
R376 B.n272 B.n271 163.367
R377 B.n271 B.n270 163.367
R378 B.n270 B.n83 163.367
R379 B.n266 B.n83 163.367
R380 B.n266 B.n265 163.367
R381 B.n265 B.n264 163.367
R382 B.n264 B.n85 163.367
R383 B.n260 B.n85 163.367
R384 B.n445 B.n444 163.367
R385 B.n444 B.n21 163.367
R386 B.n440 B.n21 163.367
R387 B.n440 B.n439 163.367
R388 B.n439 B.n438 163.367
R389 B.n438 B.n23 163.367
R390 B.n434 B.n23 163.367
R391 B.n434 B.n433 163.367
R392 B.n433 B.n432 163.367
R393 B.n432 B.n25 163.367
R394 B.n428 B.n25 163.367
R395 B.n428 B.n427 163.367
R396 B.n427 B.n426 163.367
R397 B.n426 B.n27 163.367
R398 B.n422 B.n27 163.367
R399 B.n422 B.n421 163.367
R400 B.n421 B.n420 163.367
R401 B.n420 B.n29 163.367
R402 B.n416 B.n29 163.367
R403 B.n416 B.n415 163.367
R404 B.n415 B.n33 163.367
R405 B.n411 B.n33 163.367
R406 B.n411 B.n410 163.367
R407 B.n410 B.n409 163.367
R408 B.n409 B.n35 163.367
R409 B.n405 B.n35 163.367
R410 B.n405 B.n404 163.367
R411 B.n404 B.n403 163.367
R412 B.n403 B.n37 163.367
R413 B.n398 B.n37 163.367
R414 B.n398 B.n397 163.367
R415 B.n397 B.n396 163.367
R416 B.n396 B.n41 163.367
R417 B.n392 B.n41 163.367
R418 B.n392 B.n391 163.367
R419 B.n391 B.n390 163.367
R420 B.n390 B.n43 163.367
R421 B.n386 B.n43 163.367
R422 B.n386 B.n385 163.367
R423 B.n385 B.n384 163.367
R424 B.n384 B.n45 163.367
R425 B.n380 B.n45 163.367
R426 B.n380 B.n379 163.367
R427 B.n379 B.n378 163.367
R428 B.n378 B.n47 163.367
R429 B.n374 B.n47 163.367
R430 B.n374 B.n373 163.367
R431 B.n373 B.n372 163.367
R432 B.n446 B.n19 163.367
R433 B.n450 B.n19 163.367
R434 B.n451 B.n450 163.367
R435 B.n452 B.n451 163.367
R436 B.n452 B.n17 163.367
R437 B.n456 B.n17 163.367
R438 B.n457 B.n456 163.367
R439 B.n458 B.n457 163.367
R440 B.n458 B.n15 163.367
R441 B.n462 B.n15 163.367
R442 B.n463 B.n462 163.367
R443 B.n464 B.n463 163.367
R444 B.n464 B.n13 163.367
R445 B.n468 B.n13 163.367
R446 B.n469 B.n468 163.367
R447 B.n470 B.n469 163.367
R448 B.n470 B.n11 163.367
R449 B.n474 B.n11 163.367
R450 B.n475 B.n474 163.367
R451 B.n476 B.n475 163.367
R452 B.n476 B.n9 163.367
R453 B.n480 B.n9 163.367
R454 B.n481 B.n480 163.367
R455 B.n482 B.n481 163.367
R456 B.n482 B.n7 163.367
R457 B.n486 B.n7 163.367
R458 B.n487 B.n486 163.367
R459 B.n488 B.n487 163.367
R460 B.n488 B.n5 163.367
R461 B.n492 B.n5 163.367
R462 B.n493 B.n492 163.367
R463 B.n494 B.n493 163.367
R464 B.n494 B.n3 163.367
R465 B.n498 B.n3 163.367
R466 B.n499 B.n498 163.367
R467 B.n133 B.n2 163.367
R468 B.n134 B.n133 163.367
R469 B.n134 B.n131 163.367
R470 B.n138 B.n131 163.367
R471 B.n139 B.n138 163.367
R472 B.n140 B.n139 163.367
R473 B.n140 B.n129 163.367
R474 B.n144 B.n129 163.367
R475 B.n145 B.n144 163.367
R476 B.n146 B.n145 163.367
R477 B.n146 B.n127 163.367
R478 B.n150 B.n127 163.367
R479 B.n151 B.n150 163.367
R480 B.n152 B.n151 163.367
R481 B.n152 B.n125 163.367
R482 B.n156 B.n125 163.367
R483 B.n157 B.n156 163.367
R484 B.n158 B.n157 163.367
R485 B.n158 B.n123 163.367
R486 B.n162 B.n123 163.367
R487 B.n163 B.n162 163.367
R488 B.n164 B.n163 163.367
R489 B.n164 B.n121 163.367
R490 B.n168 B.n121 163.367
R491 B.n169 B.n168 163.367
R492 B.n170 B.n169 163.367
R493 B.n170 B.n119 163.367
R494 B.n174 B.n119 163.367
R495 B.n175 B.n174 163.367
R496 B.n176 B.n175 163.367
R497 B.n176 B.n117 163.367
R498 B.n180 B.n117 163.367
R499 B.n181 B.n180 163.367
R500 B.n182 B.n181 163.367
R501 B.n182 B.n115 163.367
R502 B.n215 B.n105 59.5399
R503 B.n98 B.n97 59.5399
R504 B.n401 B.n39 59.5399
R505 B.n32 B.n31 59.5399
R506 B.n105 B.n104 37.2369
R507 B.n97 B.n96 37.2369
R508 B.n39 B.n38 37.2369
R509 B.n31 B.n30 37.2369
R510 B.n261 B.n86 28.5664
R511 B.n447 B.n20 28.5664
R512 B.n371 B.n370 28.5664
R513 B.n185 B.n184 28.5664
R514 B B.n501 18.0485
R515 B.n448 B.n447 10.6151
R516 B.n449 B.n448 10.6151
R517 B.n449 B.n18 10.6151
R518 B.n453 B.n18 10.6151
R519 B.n454 B.n453 10.6151
R520 B.n455 B.n454 10.6151
R521 B.n455 B.n16 10.6151
R522 B.n459 B.n16 10.6151
R523 B.n460 B.n459 10.6151
R524 B.n461 B.n460 10.6151
R525 B.n461 B.n14 10.6151
R526 B.n465 B.n14 10.6151
R527 B.n466 B.n465 10.6151
R528 B.n467 B.n466 10.6151
R529 B.n467 B.n12 10.6151
R530 B.n471 B.n12 10.6151
R531 B.n472 B.n471 10.6151
R532 B.n473 B.n472 10.6151
R533 B.n473 B.n10 10.6151
R534 B.n477 B.n10 10.6151
R535 B.n478 B.n477 10.6151
R536 B.n479 B.n478 10.6151
R537 B.n479 B.n8 10.6151
R538 B.n483 B.n8 10.6151
R539 B.n484 B.n483 10.6151
R540 B.n485 B.n484 10.6151
R541 B.n485 B.n6 10.6151
R542 B.n489 B.n6 10.6151
R543 B.n490 B.n489 10.6151
R544 B.n491 B.n490 10.6151
R545 B.n491 B.n4 10.6151
R546 B.n495 B.n4 10.6151
R547 B.n496 B.n495 10.6151
R548 B.n497 B.n496 10.6151
R549 B.n497 B.n0 10.6151
R550 B.n443 B.n20 10.6151
R551 B.n443 B.n442 10.6151
R552 B.n442 B.n441 10.6151
R553 B.n441 B.n22 10.6151
R554 B.n437 B.n22 10.6151
R555 B.n437 B.n436 10.6151
R556 B.n436 B.n435 10.6151
R557 B.n435 B.n24 10.6151
R558 B.n431 B.n24 10.6151
R559 B.n431 B.n430 10.6151
R560 B.n430 B.n429 10.6151
R561 B.n429 B.n26 10.6151
R562 B.n425 B.n26 10.6151
R563 B.n425 B.n424 10.6151
R564 B.n424 B.n423 10.6151
R565 B.n423 B.n28 10.6151
R566 B.n419 B.n28 10.6151
R567 B.n419 B.n418 10.6151
R568 B.n418 B.n417 10.6151
R569 B.n414 B.n413 10.6151
R570 B.n413 B.n412 10.6151
R571 B.n412 B.n34 10.6151
R572 B.n408 B.n34 10.6151
R573 B.n408 B.n407 10.6151
R574 B.n407 B.n406 10.6151
R575 B.n406 B.n36 10.6151
R576 B.n402 B.n36 10.6151
R577 B.n400 B.n399 10.6151
R578 B.n399 B.n40 10.6151
R579 B.n395 B.n40 10.6151
R580 B.n395 B.n394 10.6151
R581 B.n394 B.n393 10.6151
R582 B.n393 B.n42 10.6151
R583 B.n389 B.n42 10.6151
R584 B.n389 B.n388 10.6151
R585 B.n388 B.n387 10.6151
R586 B.n387 B.n44 10.6151
R587 B.n383 B.n44 10.6151
R588 B.n383 B.n382 10.6151
R589 B.n382 B.n381 10.6151
R590 B.n381 B.n46 10.6151
R591 B.n377 B.n46 10.6151
R592 B.n377 B.n376 10.6151
R593 B.n376 B.n375 10.6151
R594 B.n375 B.n48 10.6151
R595 B.n371 B.n48 10.6151
R596 B.n370 B.n369 10.6151
R597 B.n369 B.n50 10.6151
R598 B.n365 B.n50 10.6151
R599 B.n365 B.n364 10.6151
R600 B.n364 B.n363 10.6151
R601 B.n363 B.n52 10.6151
R602 B.n359 B.n52 10.6151
R603 B.n359 B.n358 10.6151
R604 B.n358 B.n357 10.6151
R605 B.n357 B.n54 10.6151
R606 B.n353 B.n54 10.6151
R607 B.n353 B.n352 10.6151
R608 B.n352 B.n351 10.6151
R609 B.n351 B.n56 10.6151
R610 B.n347 B.n56 10.6151
R611 B.n347 B.n346 10.6151
R612 B.n346 B.n345 10.6151
R613 B.n345 B.n58 10.6151
R614 B.n341 B.n58 10.6151
R615 B.n341 B.n340 10.6151
R616 B.n340 B.n339 10.6151
R617 B.n339 B.n60 10.6151
R618 B.n335 B.n60 10.6151
R619 B.n335 B.n334 10.6151
R620 B.n334 B.n333 10.6151
R621 B.n333 B.n62 10.6151
R622 B.n329 B.n62 10.6151
R623 B.n329 B.n328 10.6151
R624 B.n328 B.n327 10.6151
R625 B.n327 B.n64 10.6151
R626 B.n323 B.n64 10.6151
R627 B.n323 B.n322 10.6151
R628 B.n322 B.n321 10.6151
R629 B.n321 B.n66 10.6151
R630 B.n317 B.n66 10.6151
R631 B.n317 B.n316 10.6151
R632 B.n316 B.n315 10.6151
R633 B.n315 B.n68 10.6151
R634 B.n311 B.n68 10.6151
R635 B.n311 B.n310 10.6151
R636 B.n310 B.n309 10.6151
R637 B.n309 B.n70 10.6151
R638 B.n305 B.n70 10.6151
R639 B.n305 B.n304 10.6151
R640 B.n304 B.n303 10.6151
R641 B.n303 B.n72 10.6151
R642 B.n299 B.n72 10.6151
R643 B.n299 B.n298 10.6151
R644 B.n298 B.n297 10.6151
R645 B.n297 B.n74 10.6151
R646 B.n293 B.n74 10.6151
R647 B.n293 B.n292 10.6151
R648 B.n292 B.n291 10.6151
R649 B.n291 B.n76 10.6151
R650 B.n287 B.n76 10.6151
R651 B.n287 B.n286 10.6151
R652 B.n286 B.n285 10.6151
R653 B.n285 B.n78 10.6151
R654 B.n281 B.n78 10.6151
R655 B.n281 B.n280 10.6151
R656 B.n280 B.n279 10.6151
R657 B.n279 B.n80 10.6151
R658 B.n275 B.n80 10.6151
R659 B.n275 B.n274 10.6151
R660 B.n274 B.n273 10.6151
R661 B.n273 B.n82 10.6151
R662 B.n269 B.n82 10.6151
R663 B.n269 B.n268 10.6151
R664 B.n268 B.n267 10.6151
R665 B.n267 B.n84 10.6151
R666 B.n263 B.n84 10.6151
R667 B.n263 B.n262 10.6151
R668 B.n262 B.n261 10.6151
R669 B.n132 B.n1 10.6151
R670 B.n135 B.n132 10.6151
R671 B.n136 B.n135 10.6151
R672 B.n137 B.n136 10.6151
R673 B.n137 B.n130 10.6151
R674 B.n141 B.n130 10.6151
R675 B.n142 B.n141 10.6151
R676 B.n143 B.n142 10.6151
R677 B.n143 B.n128 10.6151
R678 B.n147 B.n128 10.6151
R679 B.n148 B.n147 10.6151
R680 B.n149 B.n148 10.6151
R681 B.n149 B.n126 10.6151
R682 B.n153 B.n126 10.6151
R683 B.n154 B.n153 10.6151
R684 B.n155 B.n154 10.6151
R685 B.n155 B.n124 10.6151
R686 B.n159 B.n124 10.6151
R687 B.n160 B.n159 10.6151
R688 B.n161 B.n160 10.6151
R689 B.n161 B.n122 10.6151
R690 B.n165 B.n122 10.6151
R691 B.n166 B.n165 10.6151
R692 B.n167 B.n166 10.6151
R693 B.n167 B.n120 10.6151
R694 B.n171 B.n120 10.6151
R695 B.n172 B.n171 10.6151
R696 B.n173 B.n172 10.6151
R697 B.n173 B.n118 10.6151
R698 B.n177 B.n118 10.6151
R699 B.n178 B.n177 10.6151
R700 B.n179 B.n178 10.6151
R701 B.n179 B.n116 10.6151
R702 B.n183 B.n116 10.6151
R703 B.n184 B.n183 10.6151
R704 B.n185 B.n114 10.6151
R705 B.n189 B.n114 10.6151
R706 B.n190 B.n189 10.6151
R707 B.n191 B.n190 10.6151
R708 B.n191 B.n112 10.6151
R709 B.n195 B.n112 10.6151
R710 B.n196 B.n195 10.6151
R711 B.n197 B.n196 10.6151
R712 B.n197 B.n110 10.6151
R713 B.n201 B.n110 10.6151
R714 B.n202 B.n201 10.6151
R715 B.n203 B.n202 10.6151
R716 B.n203 B.n108 10.6151
R717 B.n207 B.n108 10.6151
R718 B.n208 B.n207 10.6151
R719 B.n209 B.n208 10.6151
R720 B.n209 B.n106 10.6151
R721 B.n213 B.n106 10.6151
R722 B.n214 B.n213 10.6151
R723 B.n216 B.n102 10.6151
R724 B.n220 B.n102 10.6151
R725 B.n221 B.n220 10.6151
R726 B.n222 B.n221 10.6151
R727 B.n222 B.n100 10.6151
R728 B.n226 B.n100 10.6151
R729 B.n227 B.n226 10.6151
R730 B.n228 B.n227 10.6151
R731 B.n232 B.n231 10.6151
R732 B.n233 B.n232 10.6151
R733 B.n233 B.n94 10.6151
R734 B.n237 B.n94 10.6151
R735 B.n238 B.n237 10.6151
R736 B.n239 B.n238 10.6151
R737 B.n239 B.n92 10.6151
R738 B.n243 B.n92 10.6151
R739 B.n244 B.n243 10.6151
R740 B.n245 B.n244 10.6151
R741 B.n245 B.n90 10.6151
R742 B.n249 B.n90 10.6151
R743 B.n250 B.n249 10.6151
R744 B.n251 B.n250 10.6151
R745 B.n251 B.n88 10.6151
R746 B.n255 B.n88 10.6151
R747 B.n256 B.n255 10.6151
R748 B.n257 B.n256 10.6151
R749 B.n257 B.n86 10.6151
R750 B.n501 B.n0 8.11757
R751 B.n501 B.n1 8.11757
R752 B.n414 B.n32 6.5566
R753 B.n402 B.n401 6.5566
R754 B.n216 B.n215 6.5566
R755 B.n228 B.n98 6.5566
R756 B.n417 B.n32 4.05904
R757 B.n401 B.n400 4.05904
R758 B.n215 B.n214 4.05904
R759 B.n231 B.n98 4.05904
R760 VN.n20 VN.n19 179.499
R761 VN.n41 VN.n40 179.499
R762 VN.n39 VN.n21 161.3
R763 VN.n38 VN.n37 161.3
R764 VN.n36 VN.n22 161.3
R765 VN.n35 VN.n34 161.3
R766 VN.n32 VN.n23 161.3
R767 VN.n31 VN.n30 161.3
R768 VN.n29 VN.n24 161.3
R769 VN.n28 VN.n27 161.3
R770 VN.n18 VN.n0 161.3
R771 VN.n17 VN.n16 161.3
R772 VN.n15 VN.n1 161.3
R773 VN.n14 VN.n13 161.3
R774 VN.n11 VN.n2 161.3
R775 VN.n10 VN.n9 161.3
R776 VN.n8 VN.n3 161.3
R777 VN.n7 VN.n6 161.3
R778 VN.n4 VN.t0 99.7665
R779 VN.n25 VN.t2 99.7665
R780 VN.n5 VN.t7 67.9049
R781 VN.n12 VN.t6 67.9049
R782 VN.n19 VN.t5 67.9049
R783 VN.n26 VN.t3 67.9049
R784 VN.n33 VN.t4 67.9049
R785 VN.n40 VN.t1 67.9049
R786 VN.n10 VN.n3 56.5617
R787 VN.n31 VN.n24 56.5617
R788 VN.n17 VN.n1 56.5617
R789 VN.n38 VN.n22 56.5617
R790 VN.n5 VN.n4 55.8951
R791 VN.n26 VN.n25 55.8951
R792 VN VN.n41 40.7448
R793 VN.n6 VN.n3 24.5923
R794 VN.n11 VN.n10 24.5923
R795 VN.n13 VN.n1 24.5923
R796 VN.n18 VN.n17 24.5923
R797 VN.n27 VN.n24 24.5923
R798 VN.n34 VN.n22 24.5923
R799 VN.n32 VN.n31 24.5923
R800 VN.n39 VN.n38 24.5923
R801 VN.n28 VN.n25 18.12
R802 VN.n7 VN.n4 18.12
R803 VN.n13 VN.n12 14.2638
R804 VN.n34 VN.n33 14.2638
R805 VN.n6 VN.n5 10.3291
R806 VN.n12 VN.n11 10.3291
R807 VN.n27 VN.n26 10.3291
R808 VN.n33 VN.n32 10.3291
R809 VN.n19 VN.n18 6.39438
R810 VN.n40 VN.n39 6.39438
R811 VN.n41 VN.n21 0.189894
R812 VN.n37 VN.n21 0.189894
R813 VN.n37 VN.n36 0.189894
R814 VN.n36 VN.n35 0.189894
R815 VN.n35 VN.n23 0.189894
R816 VN.n30 VN.n23 0.189894
R817 VN.n30 VN.n29 0.189894
R818 VN.n29 VN.n28 0.189894
R819 VN.n8 VN.n7 0.189894
R820 VN.n9 VN.n8 0.189894
R821 VN.n9 VN.n2 0.189894
R822 VN.n14 VN.n2 0.189894
R823 VN.n15 VN.n14 0.189894
R824 VN.n16 VN.n15 0.189894
R825 VN.n16 VN.n0 0.189894
R826 VN.n20 VN.n0 0.189894
R827 VN VN.n20 0.0516364
R828 VDD2.n2 VDD2.n1 103.3
R829 VDD2.n2 VDD2.n0 103.3
R830 VDD2 VDD2.n5 103.297
R831 VDD2.n4 VDD2.n3 102.528
R832 VDD2.n4 VDD2.n2 35.0256
R833 VDD2.n5 VDD2.t2 7.25608
R834 VDD2.n5 VDD2.t1 7.25608
R835 VDD2.n3 VDD2.t5 7.25608
R836 VDD2.n3 VDD2.t7 7.25608
R837 VDD2.n1 VDD2.t3 7.25608
R838 VDD2.n1 VDD2.t6 7.25608
R839 VDD2.n0 VDD2.t0 7.25608
R840 VDD2.n0 VDD2.t4 7.25608
R841 VDD2 VDD2.n4 0.886276
R842 VTAIL.n194 VTAIL.n176 756.745
R843 VTAIL.n20 VTAIL.n2 756.745
R844 VTAIL.n44 VTAIL.n26 756.745
R845 VTAIL.n70 VTAIL.n52 756.745
R846 VTAIL.n170 VTAIL.n152 756.745
R847 VTAIL.n144 VTAIL.n126 756.745
R848 VTAIL.n120 VTAIL.n102 756.745
R849 VTAIL.n94 VTAIL.n76 756.745
R850 VTAIL.n185 VTAIL.n184 585
R851 VTAIL.n187 VTAIL.n186 585
R852 VTAIL.n180 VTAIL.n179 585
R853 VTAIL.n193 VTAIL.n192 585
R854 VTAIL.n195 VTAIL.n194 585
R855 VTAIL.n11 VTAIL.n10 585
R856 VTAIL.n13 VTAIL.n12 585
R857 VTAIL.n6 VTAIL.n5 585
R858 VTAIL.n19 VTAIL.n18 585
R859 VTAIL.n21 VTAIL.n20 585
R860 VTAIL.n35 VTAIL.n34 585
R861 VTAIL.n37 VTAIL.n36 585
R862 VTAIL.n30 VTAIL.n29 585
R863 VTAIL.n43 VTAIL.n42 585
R864 VTAIL.n45 VTAIL.n44 585
R865 VTAIL.n61 VTAIL.n60 585
R866 VTAIL.n63 VTAIL.n62 585
R867 VTAIL.n56 VTAIL.n55 585
R868 VTAIL.n69 VTAIL.n68 585
R869 VTAIL.n71 VTAIL.n70 585
R870 VTAIL.n171 VTAIL.n170 585
R871 VTAIL.n169 VTAIL.n168 585
R872 VTAIL.n156 VTAIL.n155 585
R873 VTAIL.n163 VTAIL.n162 585
R874 VTAIL.n161 VTAIL.n160 585
R875 VTAIL.n145 VTAIL.n144 585
R876 VTAIL.n143 VTAIL.n142 585
R877 VTAIL.n130 VTAIL.n129 585
R878 VTAIL.n137 VTAIL.n136 585
R879 VTAIL.n135 VTAIL.n134 585
R880 VTAIL.n121 VTAIL.n120 585
R881 VTAIL.n119 VTAIL.n118 585
R882 VTAIL.n106 VTAIL.n105 585
R883 VTAIL.n113 VTAIL.n112 585
R884 VTAIL.n111 VTAIL.n110 585
R885 VTAIL.n95 VTAIL.n94 585
R886 VTAIL.n93 VTAIL.n92 585
R887 VTAIL.n80 VTAIL.n79 585
R888 VTAIL.n87 VTAIL.n86 585
R889 VTAIL.n85 VTAIL.n84 585
R890 VTAIL.n183 VTAIL.t10 328.587
R891 VTAIL.n9 VTAIL.t15 328.587
R892 VTAIL.n33 VTAIL.t1 328.587
R893 VTAIL.n59 VTAIL.t0 328.587
R894 VTAIL.n159 VTAIL.t7 328.587
R895 VTAIL.n133 VTAIL.t6 328.587
R896 VTAIL.n109 VTAIL.t13 328.587
R897 VTAIL.n83 VTAIL.t14 328.587
R898 VTAIL.n186 VTAIL.n185 171.744
R899 VTAIL.n186 VTAIL.n179 171.744
R900 VTAIL.n193 VTAIL.n179 171.744
R901 VTAIL.n194 VTAIL.n193 171.744
R902 VTAIL.n12 VTAIL.n11 171.744
R903 VTAIL.n12 VTAIL.n5 171.744
R904 VTAIL.n19 VTAIL.n5 171.744
R905 VTAIL.n20 VTAIL.n19 171.744
R906 VTAIL.n36 VTAIL.n35 171.744
R907 VTAIL.n36 VTAIL.n29 171.744
R908 VTAIL.n43 VTAIL.n29 171.744
R909 VTAIL.n44 VTAIL.n43 171.744
R910 VTAIL.n62 VTAIL.n61 171.744
R911 VTAIL.n62 VTAIL.n55 171.744
R912 VTAIL.n69 VTAIL.n55 171.744
R913 VTAIL.n70 VTAIL.n69 171.744
R914 VTAIL.n170 VTAIL.n169 171.744
R915 VTAIL.n169 VTAIL.n155 171.744
R916 VTAIL.n162 VTAIL.n155 171.744
R917 VTAIL.n162 VTAIL.n161 171.744
R918 VTAIL.n144 VTAIL.n143 171.744
R919 VTAIL.n143 VTAIL.n129 171.744
R920 VTAIL.n136 VTAIL.n129 171.744
R921 VTAIL.n136 VTAIL.n135 171.744
R922 VTAIL.n120 VTAIL.n119 171.744
R923 VTAIL.n119 VTAIL.n105 171.744
R924 VTAIL.n112 VTAIL.n105 171.744
R925 VTAIL.n112 VTAIL.n111 171.744
R926 VTAIL.n94 VTAIL.n93 171.744
R927 VTAIL.n93 VTAIL.n79 171.744
R928 VTAIL.n86 VTAIL.n79 171.744
R929 VTAIL.n86 VTAIL.n85 171.744
R930 VTAIL.n185 VTAIL.t10 85.8723
R931 VTAIL.n11 VTAIL.t15 85.8723
R932 VTAIL.n35 VTAIL.t1 85.8723
R933 VTAIL.n61 VTAIL.t0 85.8723
R934 VTAIL.n161 VTAIL.t7 85.8723
R935 VTAIL.n135 VTAIL.t6 85.8723
R936 VTAIL.n111 VTAIL.t13 85.8723
R937 VTAIL.n85 VTAIL.t14 85.8723
R938 VTAIL.n151 VTAIL.n150 85.8495
R939 VTAIL.n101 VTAIL.n100 85.8495
R940 VTAIL.n1 VTAIL.n0 85.8494
R941 VTAIL.n51 VTAIL.n50 85.8494
R942 VTAIL.n199 VTAIL.n198 30.6338
R943 VTAIL.n25 VTAIL.n24 30.6338
R944 VTAIL.n49 VTAIL.n48 30.6338
R945 VTAIL.n75 VTAIL.n74 30.6338
R946 VTAIL.n175 VTAIL.n174 30.6338
R947 VTAIL.n149 VTAIL.n148 30.6338
R948 VTAIL.n125 VTAIL.n124 30.6338
R949 VTAIL.n99 VTAIL.n98 30.6338
R950 VTAIL.n199 VTAIL.n175 17.8841
R951 VTAIL.n99 VTAIL.n75 17.8841
R952 VTAIL.n184 VTAIL.n183 16.3651
R953 VTAIL.n10 VTAIL.n9 16.3651
R954 VTAIL.n34 VTAIL.n33 16.3651
R955 VTAIL.n60 VTAIL.n59 16.3651
R956 VTAIL.n160 VTAIL.n159 16.3651
R957 VTAIL.n134 VTAIL.n133 16.3651
R958 VTAIL.n110 VTAIL.n109 16.3651
R959 VTAIL.n84 VTAIL.n83 16.3651
R960 VTAIL.n187 VTAIL.n182 12.8005
R961 VTAIL.n13 VTAIL.n8 12.8005
R962 VTAIL.n37 VTAIL.n32 12.8005
R963 VTAIL.n63 VTAIL.n58 12.8005
R964 VTAIL.n163 VTAIL.n158 12.8005
R965 VTAIL.n137 VTAIL.n132 12.8005
R966 VTAIL.n113 VTAIL.n108 12.8005
R967 VTAIL.n87 VTAIL.n82 12.8005
R968 VTAIL.n188 VTAIL.n180 12.0247
R969 VTAIL.n14 VTAIL.n6 12.0247
R970 VTAIL.n38 VTAIL.n30 12.0247
R971 VTAIL.n64 VTAIL.n56 12.0247
R972 VTAIL.n164 VTAIL.n156 12.0247
R973 VTAIL.n138 VTAIL.n130 12.0247
R974 VTAIL.n114 VTAIL.n106 12.0247
R975 VTAIL.n88 VTAIL.n80 12.0247
R976 VTAIL.n192 VTAIL.n191 11.249
R977 VTAIL.n18 VTAIL.n17 11.249
R978 VTAIL.n42 VTAIL.n41 11.249
R979 VTAIL.n68 VTAIL.n67 11.249
R980 VTAIL.n168 VTAIL.n167 11.249
R981 VTAIL.n142 VTAIL.n141 11.249
R982 VTAIL.n118 VTAIL.n117 11.249
R983 VTAIL.n92 VTAIL.n91 11.249
R984 VTAIL.n195 VTAIL.n178 10.4732
R985 VTAIL.n21 VTAIL.n4 10.4732
R986 VTAIL.n45 VTAIL.n28 10.4732
R987 VTAIL.n71 VTAIL.n54 10.4732
R988 VTAIL.n171 VTAIL.n154 10.4732
R989 VTAIL.n145 VTAIL.n128 10.4732
R990 VTAIL.n121 VTAIL.n104 10.4732
R991 VTAIL.n95 VTAIL.n78 10.4732
R992 VTAIL.n196 VTAIL.n176 9.69747
R993 VTAIL.n22 VTAIL.n2 9.69747
R994 VTAIL.n46 VTAIL.n26 9.69747
R995 VTAIL.n72 VTAIL.n52 9.69747
R996 VTAIL.n172 VTAIL.n152 9.69747
R997 VTAIL.n146 VTAIL.n126 9.69747
R998 VTAIL.n122 VTAIL.n102 9.69747
R999 VTAIL.n96 VTAIL.n76 9.69747
R1000 VTAIL.n198 VTAIL.n197 9.45567
R1001 VTAIL.n24 VTAIL.n23 9.45567
R1002 VTAIL.n48 VTAIL.n47 9.45567
R1003 VTAIL.n74 VTAIL.n73 9.45567
R1004 VTAIL.n174 VTAIL.n173 9.45567
R1005 VTAIL.n148 VTAIL.n147 9.45567
R1006 VTAIL.n124 VTAIL.n123 9.45567
R1007 VTAIL.n98 VTAIL.n97 9.45567
R1008 VTAIL.n197 VTAIL.n196 9.3005
R1009 VTAIL.n178 VTAIL.n177 9.3005
R1010 VTAIL.n191 VTAIL.n190 9.3005
R1011 VTAIL.n189 VTAIL.n188 9.3005
R1012 VTAIL.n182 VTAIL.n181 9.3005
R1013 VTAIL.n23 VTAIL.n22 9.3005
R1014 VTAIL.n4 VTAIL.n3 9.3005
R1015 VTAIL.n17 VTAIL.n16 9.3005
R1016 VTAIL.n15 VTAIL.n14 9.3005
R1017 VTAIL.n8 VTAIL.n7 9.3005
R1018 VTAIL.n47 VTAIL.n46 9.3005
R1019 VTAIL.n28 VTAIL.n27 9.3005
R1020 VTAIL.n41 VTAIL.n40 9.3005
R1021 VTAIL.n39 VTAIL.n38 9.3005
R1022 VTAIL.n32 VTAIL.n31 9.3005
R1023 VTAIL.n73 VTAIL.n72 9.3005
R1024 VTAIL.n54 VTAIL.n53 9.3005
R1025 VTAIL.n67 VTAIL.n66 9.3005
R1026 VTAIL.n65 VTAIL.n64 9.3005
R1027 VTAIL.n58 VTAIL.n57 9.3005
R1028 VTAIL.n173 VTAIL.n172 9.3005
R1029 VTAIL.n154 VTAIL.n153 9.3005
R1030 VTAIL.n167 VTAIL.n166 9.3005
R1031 VTAIL.n165 VTAIL.n164 9.3005
R1032 VTAIL.n158 VTAIL.n157 9.3005
R1033 VTAIL.n147 VTAIL.n146 9.3005
R1034 VTAIL.n128 VTAIL.n127 9.3005
R1035 VTAIL.n141 VTAIL.n140 9.3005
R1036 VTAIL.n139 VTAIL.n138 9.3005
R1037 VTAIL.n132 VTAIL.n131 9.3005
R1038 VTAIL.n123 VTAIL.n122 9.3005
R1039 VTAIL.n104 VTAIL.n103 9.3005
R1040 VTAIL.n117 VTAIL.n116 9.3005
R1041 VTAIL.n115 VTAIL.n114 9.3005
R1042 VTAIL.n108 VTAIL.n107 9.3005
R1043 VTAIL.n97 VTAIL.n96 9.3005
R1044 VTAIL.n78 VTAIL.n77 9.3005
R1045 VTAIL.n91 VTAIL.n90 9.3005
R1046 VTAIL.n89 VTAIL.n88 9.3005
R1047 VTAIL.n82 VTAIL.n81 9.3005
R1048 VTAIL.n0 VTAIL.t8 7.25608
R1049 VTAIL.n0 VTAIL.t9 7.25608
R1050 VTAIL.n50 VTAIL.t3 7.25608
R1051 VTAIL.n50 VTAIL.t2 7.25608
R1052 VTAIL.n150 VTAIL.t4 7.25608
R1053 VTAIL.n150 VTAIL.t5 7.25608
R1054 VTAIL.n100 VTAIL.t11 7.25608
R1055 VTAIL.n100 VTAIL.t12 7.25608
R1056 VTAIL.n198 VTAIL.n176 4.26717
R1057 VTAIL.n24 VTAIL.n2 4.26717
R1058 VTAIL.n48 VTAIL.n26 4.26717
R1059 VTAIL.n74 VTAIL.n52 4.26717
R1060 VTAIL.n174 VTAIL.n152 4.26717
R1061 VTAIL.n148 VTAIL.n126 4.26717
R1062 VTAIL.n124 VTAIL.n102 4.26717
R1063 VTAIL.n98 VTAIL.n76 4.26717
R1064 VTAIL.n183 VTAIL.n181 3.73474
R1065 VTAIL.n9 VTAIL.n7 3.73474
R1066 VTAIL.n33 VTAIL.n31 3.73474
R1067 VTAIL.n59 VTAIL.n57 3.73474
R1068 VTAIL.n159 VTAIL.n157 3.73474
R1069 VTAIL.n133 VTAIL.n131 3.73474
R1070 VTAIL.n109 VTAIL.n107 3.73474
R1071 VTAIL.n83 VTAIL.n81 3.73474
R1072 VTAIL.n196 VTAIL.n195 3.49141
R1073 VTAIL.n22 VTAIL.n21 3.49141
R1074 VTAIL.n46 VTAIL.n45 3.49141
R1075 VTAIL.n72 VTAIL.n71 3.49141
R1076 VTAIL.n172 VTAIL.n171 3.49141
R1077 VTAIL.n146 VTAIL.n145 3.49141
R1078 VTAIL.n122 VTAIL.n121 3.49141
R1079 VTAIL.n96 VTAIL.n95 3.49141
R1080 VTAIL.n192 VTAIL.n178 2.71565
R1081 VTAIL.n18 VTAIL.n4 2.71565
R1082 VTAIL.n42 VTAIL.n28 2.71565
R1083 VTAIL.n68 VTAIL.n54 2.71565
R1084 VTAIL.n168 VTAIL.n154 2.71565
R1085 VTAIL.n142 VTAIL.n128 2.71565
R1086 VTAIL.n118 VTAIL.n104 2.71565
R1087 VTAIL.n92 VTAIL.n78 2.71565
R1088 VTAIL.n191 VTAIL.n180 1.93989
R1089 VTAIL.n17 VTAIL.n6 1.93989
R1090 VTAIL.n41 VTAIL.n30 1.93989
R1091 VTAIL.n67 VTAIL.n56 1.93989
R1092 VTAIL.n167 VTAIL.n156 1.93989
R1093 VTAIL.n141 VTAIL.n130 1.93989
R1094 VTAIL.n117 VTAIL.n106 1.93989
R1095 VTAIL.n91 VTAIL.n80 1.93989
R1096 VTAIL.n101 VTAIL.n99 1.65567
R1097 VTAIL.n125 VTAIL.n101 1.65567
R1098 VTAIL.n151 VTAIL.n149 1.65567
R1099 VTAIL.n175 VTAIL.n151 1.65567
R1100 VTAIL.n75 VTAIL.n51 1.65567
R1101 VTAIL.n51 VTAIL.n49 1.65567
R1102 VTAIL.n25 VTAIL.n1 1.65567
R1103 VTAIL VTAIL.n199 1.59748
R1104 VTAIL.n188 VTAIL.n187 1.16414
R1105 VTAIL.n14 VTAIL.n13 1.16414
R1106 VTAIL.n38 VTAIL.n37 1.16414
R1107 VTAIL.n64 VTAIL.n63 1.16414
R1108 VTAIL.n164 VTAIL.n163 1.16414
R1109 VTAIL.n138 VTAIL.n137 1.16414
R1110 VTAIL.n114 VTAIL.n113 1.16414
R1111 VTAIL.n88 VTAIL.n87 1.16414
R1112 VTAIL.n149 VTAIL.n125 0.470328
R1113 VTAIL.n49 VTAIL.n25 0.470328
R1114 VTAIL.n184 VTAIL.n182 0.388379
R1115 VTAIL.n10 VTAIL.n8 0.388379
R1116 VTAIL.n34 VTAIL.n32 0.388379
R1117 VTAIL.n60 VTAIL.n58 0.388379
R1118 VTAIL.n160 VTAIL.n158 0.388379
R1119 VTAIL.n134 VTAIL.n132 0.388379
R1120 VTAIL.n110 VTAIL.n108 0.388379
R1121 VTAIL.n84 VTAIL.n82 0.388379
R1122 VTAIL.n189 VTAIL.n181 0.155672
R1123 VTAIL.n190 VTAIL.n189 0.155672
R1124 VTAIL.n190 VTAIL.n177 0.155672
R1125 VTAIL.n197 VTAIL.n177 0.155672
R1126 VTAIL.n15 VTAIL.n7 0.155672
R1127 VTAIL.n16 VTAIL.n15 0.155672
R1128 VTAIL.n16 VTAIL.n3 0.155672
R1129 VTAIL.n23 VTAIL.n3 0.155672
R1130 VTAIL.n39 VTAIL.n31 0.155672
R1131 VTAIL.n40 VTAIL.n39 0.155672
R1132 VTAIL.n40 VTAIL.n27 0.155672
R1133 VTAIL.n47 VTAIL.n27 0.155672
R1134 VTAIL.n65 VTAIL.n57 0.155672
R1135 VTAIL.n66 VTAIL.n65 0.155672
R1136 VTAIL.n66 VTAIL.n53 0.155672
R1137 VTAIL.n73 VTAIL.n53 0.155672
R1138 VTAIL.n173 VTAIL.n153 0.155672
R1139 VTAIL.n166 VTAIL.n153 0.155672
R1140 VTAIL.n166 VTAIL.n165 0.155672
R1141 VTAIL.n165 VTAIL.n157 0.155672
R1142 VTAIL.n147 VTAIL.n127 0.155672
R1143 VTAIL.n140 VTAIL.n127 0.155672
R1144 VTAIL.n140 VTAIL.n139 0.155672
R1145 VTAIL.n139 VTAIL.n131 0.155672
R1146 VTAIL.n123 VTAIL.n103 0.155672
R1147 VTAIL.n116 VTAIL.n103 0.155672
R1148 VTAIL.n116 VTAIL.n115 0.155672
R1149 VTAIL.n115 VTAIL.n107 0.155672
R1150 VTAIL.n97 VTAIL.n77 0.155672
R1151 VTAIL.n90 VTAIL.n77 0.155672
R1152 VTAIL.n90 VTAIL.n89 0.155672
R1153 VTAIL.n89 VTAIL.n81 0.155672
R1154 VTAIL VTAIL.n1 0.0586897
R1155 VP.n28 VP.n27 179.499
R1156 VP.n50 VP.n49 179.499
R1157 VP.n26 VP.n25 179.499
R1158 VP.n13 VP.n12 161.3
R1159 VP.n14 VP.n9 161.3
R1160 VP.n16 VP.n15 161.3
R1161 VP.n17 VP.n8 161.3
R1162 VP.n20 VP.n19 161.3
R1163 VP.n21 VP.n7 161.3
R1164 VP.n23 VP.n22 161.3
R1165 VP.n24 VP.n6 161.3
R1166 VP.n48 VP.n0 161.3
R1167 VP.n47 VP.n46 161.3
R1168 VP.n45 VP.n1 161.3
R1169 VP.n44 VP.n43 161.3
R1170 VP.n41 VP.n2 161.3
R1171 VP.n40 VP.n39 161.3
R1172 VP.n38 VP.n3 161.3
R1173 VP.n37 VP.n36 161.3
R1174 VP.n34 VP.n4 161.3
R1175 VP.n33 VP.n32 161.3
R1176 VP.n31 VP.n5 161.3
R1177 VP.n30 VP.n29 161.3
R1178 VP.n10 VP.t4 99.7665
R1179 VP.n28 VP.t7 67.9049
R1180 VP.n35 VP.t0 67.9049
R1181 VP.n42 VP.t5 67.9049
R1182 VP.n49 VP.t6 67.9049
R1183 VP.n25 VP.t1 67.9049
R1184 VP.n18 VP.t2 67.9049
R1185 VP.n11 VP.t3 67.9049
R1186 VP.n40 VP.n3 56.5617
R1187 VP.n16 VP.n9 56.5617
R1188 VP.n33 VP.n5 56.5617
R1189 VP.n47 VP.n1 56.5617
R1190 VP.n23 VP.n7 56.5617
R1191 VP.n11 VP.n10 55.8951
R1192 VP.n27 VP.n26 40.3641
R1193 VP.n29 VP.n5 24.5923
R1194 VP.n34 VP.n33 24.5923
R1195 VP.n36 VP.n3 24.5923
R1196 VP.n41 VP.n40 24.5923
R1197 VP.n43 VP.n1 24.5923
R1198 VP.n48 VP.n47 24.5923
R1199 VP.n24 VP.n23 24.5923
R1200 VP.n17 VP.n16 24.5923
R1201 VP.n19 VP.n7 24.5923
R1202 VP.n12 VP.n9 24.5923
R1203 VP.n13 VP.n10 18.12
R1204 VP.n35 VP.n34 14.2638
R1205 VP.n43 VP.n42 14.2638
R1206 VP.n19 VP.n18 14.2638
R1207 VP.n36 VP.n35 10.3291
R1208 VP.n42 VP.n41 10.3291
R1209 VP.n18 VP.n17 10.3291
R1210 VP.n12 VP.n11 10.3291
R1211 VP.n29 VP.n28 6.39438
R1212 VP.n49 VP.n48 6.39438
R1213 VP.n25 VP.n24 6.39438
R1214 VP.n14 VP.n13 0.189894
R1215 VP.n15 VP.n14 0.189894
R1216 VP.n15 VP.n8 0.189894
R1217 VP.n20 VP.n8 0.189894
R1218 VP.n21 VP.n20 0.189894
R1219 VP.n22 VP.n21 0.189894
R1220 VP.n22 VP.n6 0.189894
R1221 VP.n26 VP.n6 0.189894
R1222 VP.n30 VP.n27 0.189894
R1223 VP.n31 VP.n30 0.189894
R1224 VP.n32 VP.n31 0.189894
R1225 VP.n32 VP.n4 0.189894
R1226 VP.n37 VP.n4 0.189894
R1227 VP.n38 VP.n37 0.189894
R1228 VP.n39 VP.n38 0.189894
R1229 VP.n39 VP.n2 0.189894
R1230 VP.n44 VP.n2 0.189894
R1231 VP.n45 VP.n44 0.189894
R1232 VP.n46 VP.n45 0.189894
R1233 VP.n46 VP.n0 0.189894
R1234 VP.n50 VP.n0 0.189894
R1235 VP VP.n50 0.0516364
R1236 VDD1 VDD1.n0 103.415
R1237 VDD1.n3 VDD1.n2 103.3
R1238 VDD1.n3 VDD1.n1 103.3
R1239 VDD1.n5 VDD1.n4 102.528
R1240 VDD1.n5 VDD1.n3 35.6086
R1241 VDD1.n4 VDD1.t5 7.25608
R1242 VDD1.n4 VDD1.t6 7.25608
R1243 VDD1.n0 VDD1.t3 7.25608
R1244 VDD1.n0 VDD1.t4 7.25608
R1245 VDD1.n2 VDD1.t2 7.25608
R1246 VDD1.n2 VDD1.t1 7.25608
R1247 VDD1.n1 VDD1.t0 7.25608
R1248 VDD1.n1 VDD1.t7 7.25608
R1249 VDD1 VDD1.n5 0.769897
C0 VDD2 w_n2890_n1864# 1.49385f
C1 VN B 0.922466f
C2 VDD1 w_n2890_n1864# 1.4218f
C3 VDD2 VP 0.417067f
C4 VTAIL w_n2890_n1864# 2.38376f
C5 VDD1 VP 3.39878f
C6 VDD1 VDD2 1.2552f
C7 VN w_n2890_n1864# 5.45317f
C8 VTAIL VP 3.65967f
C9 VTAIL VDD2 5.056839f
C10 w_n2890_n1864# B 6.46714f
C11 VN VP 5.03638f
C12 VDD1 VTAIL 5.009201f
C13 VN VDD2 3.13743f
C14 VDD1 VN 0.154347f
C15 VP B 1.54091f
C16 VDD2 B 1.20356f
C17 VTAIL VN 3.64557f
C18 VDD1 B 1.13921f
C19 VTAIL B 2.15447f
C20 VP w_n2890_n1864# 5.8251f
C21 VDD2 VSUBS 1.249632f
C22 VDD1 VSUBS 1.720068f
C23 VTAIL VSUBS 0.553731f
C24 VN VSUBS 5.10399f
C25 VP VSUBS 2.073892f
C26 B VSUBS 3.066845f
C27 w_n2890_n1864# VSUBS 67.6607f
C28 VDD1.t3 VSUBS 0.088496f
C29 VDD1.t4 VSUBS 0.088496f
C30 VDD1.n0 VSUBS 0.541179f
C31 VDD1.t0 VSUBS 0.088496f
C32 VDD1.t7 VSUBS 0.088496f
C33 VDD1.n1 VSUBS 0.540477f
C34 VDD1.t2 VSUBS 0.088496f
C35 VDD1.t1 VSUBS 0.088496f
C36 VDD1.n2 VSUBS 0.540477f
C37 VDD1.n3 VSUBS 2.61811f
C38 VDD1.t5 VSUBS 0.088496f
C39 VDD1.t6 VSUBS 0.088496f
C40 VDD1.n4 VSUBS 0.536172f
C41 VDD1.n5 VSUBS 2.20309f
C42 VP.n0 VSUBS 0.050388f
C43 VP.t6 VSUBS 0.931027f
C44 VP.n1 VSUBS 0.062094f
C45 VP.n2 VSUBS 0.050388f
C46 VP.t5 VSUBS 0.931027f
C47 VP.n3 VSUBS 0.073246f
C48 VP.n4 VSUBS 0.050388f
C49 VP.t0 VSUBS 0.931027f
C50 VP.n5 VSUBS 0.084399f
C51 VP.n6 VSUBS 0.050388f
C52 VP.t1 VSUBS 0.931027f
C53 VP.n7 VSUBS 0.062094f
C54 VP.n8 VSUBS 0.050388f
C55 VP.t2 VSUBS 0.931027f
C56 VP.n9 VSUBS 0.073246f
C57 VP.t4 VSUBS 1.11742f
C58 VP.n10 VSUBS 0.488754f
C59 VP.t3 VSUBS 0.931027f
C60 VP.n11 VSUBS 0.475098f
C61 VP.n12 VSUBS 0.066685f
C62 VP.n13 VSUBS 0.319388f
C63 VP.n14 VSUBS 0.050388f
C64 VP.n15 VSUBS 0.050388f
C65 VP.n16 VSUBS 0.073246f
C66 VP.n17 VSUBS 0.066685f
C67 VP.n18 VSUBS 0.381418f
C68 VP.n19 VSUBS 0.074065f
C69 VP.n20 VSUBS 0.050388f
C70 VP.n21 VSUBS 0.050388f
C71 VP.n22 VSUBS 0.050388f
C72 VP.n23 VSUBS 0.084399f
C73 VP.n24 VSUBS 0.059304f
C74 VP.n25 VSUBS 0.483623f
C75 VP.n26 VSUBS 1.95628f
C76 VP.n27 VSUBS 2.00128f
C77 VP.t7 VSUBS 0.931027f
C78 VP.n28 VSUBS 0.483623f
C79 VP.n29 VSUBS 0.059304f
C80 VP.n30 VSUBS 0.050388f
C81 VP.n31 VSUBS 0.050388f
C82 VP.n32 VSUBS 0.050388f
C83 VP.n33 VSUBS 0.062094f
C84 VP.n34 VSUBS 0.074065f
C85 VP.n35 VSUBS 0.381418f
C86 VP.n36 VSUBS 0.066685f
C87 VP.n37 VSUBS 0.050388f
C88 VP.n38 VSUBS 0.050388f
C89 VP.n39 VSUBS 0.050388f
C90 VP.n40 VSUBS 0.073246f
C91 VP.n41 VSUBS 0.066685f
C92 VP.n42 VSUBS 0.381418f
C93 VP.n43 VSUBS 0.074065f
C94 VP.n44 VSUBS 0.050388f
C95 VP.n45 VSUBS 0.050388f
C96 VP.n46 VSUBS 0.050388f
C97 VP.n47 VSUBS 0.084399f
C98 VP.n48 VSUBS 0.059304f
C99 VP.n49 VSUBS 0.483623f
C100 VP.n50 VSUBS 0.050579f
C101 VTAIL.t8 VSUBS 0.105129f
C102 VTAIL.t9 VSUBS 0.105129f
C103 VTAIL.n0 VSUBS 0.552772f
C104 VTAIL.n1 VSUBS 0.64669f
C105 VTAIL.n2 VSUBS 0.030491f
C106 VTAIL.n3 VSUBS 0.029695f
C107 VTAIL.n4 VSUBS 0.015957f
C108 VTAIL.n5 VSUBS 0.037717f
C109 VTAIL.n6 VSUBS 0.016896f
C110 VTAIL.n7 VSUBS 0.475254f
C111 VTAIL.n8 VSUBS 0.015957f
C112 VTAIL.t15 VSUBS 0.081527f
C113 VTAIL.n9 VSUBS 0.118393f
C114 VTAIL.n10 VSUBS 0.023894f
C115 VTAIL.n11 VSUBS 0.028287f
C116 VTAIL.n12 VSUBS 0.037717f
C117 VTAIL.n13 VSUBS 0.016896f
C118 VTAIL.n14 VSUBS 0.015957f
C119 VTAIL.n15 VSUBS 0.029695f
C120 VTAIL.n16 VSUBS 0.029695f
C121 VTAIL.n17 VSUBS 0.015957f
C122 VTAIL.n18 VSUBS 0.016896f
C123 VTAIL.n19 VSUBS 0.037717f
C124 VTAIL.n20 VSUBS 0.084025f
C125 VTAIL.n21 VSUBS 0.016896f
C126 VTAIL.n22 VSUBS 0.015957f
C127 VTAIL.n23 VSUBS 0.065394f
C128 VTAIL.n24 VSUBS 0.04183f
C129 VTAIL.n25 VSUBS 0.226864f
C130 VTAIL.n26 VSUBS 0.030491f
C131 VTAIL.n27 VSUBS 0.029695f
C132 VTAIL.n28 VSUBS 0.015957f
C133 VTAIL.n29 VSUBS 0.037717f
C134 VTAIL.n30 VSUBS 0.016896f
C135 VTAIL.n31 VSUBS 0.475254f
C136 VTAIL.n32 VSUBS 0.015957f
C137 VTAIL.t1 VSUBS 0.081527f
C138 VTAIL.n33 VSUBS 0.118393f
C139 VTAIL.n34 VSUBS 0.023894f
C140 VTAIL.n35 VSUBS 0.028287f
C141 VTAIL.n36 VSUBS 0.037717f
C142 VTAIL.n37 VSUBS 0.016896f
C143 VTAIL.n38 VSUBS 0.015957f
C144 VTAIL.n39 VSUBS 0.029695f
C145 VTAIL.n40 VSUBS 0.029695f
C146 VTAIL.n41 VSUBS 0.015957f
C147 VTAIL.n42 VSUBS 0.016896f
C148 VTAIL.n43 VSUBS 0.037717f
C149 VTAIL.n44 VSUBS 0.084025f
C150 VTAIL.n45 VSUBS 0.016896f
C151 VTAIL.n46 VSUBS 0.015957f
C152 VTAIL.n47 VSUBS 0.065394f
C153 VTAIL.n48 VSUBS 0.04183f
C154 VTAIL.n49 VSUBS 0.226864f
C155 VTAIL.t3 VSUBS 0.105129f
C156 VTAIL.t2 VSUBS 0.105129f
C157 VTAIL.n50 VSUBS 0.552772f
C158 VTAIL.n51 VSUBS 0.799498f
C159 VTAIL.n52 VSUBS 0.030491f
C160 VTAIL.n53 VSUBS 0.029695f
C161 VTAIL.n54 VSUBS 0.015957f
C162 VTAIL.n55 VSUBS 0.037717f
C163 VTAIL.n56 VSUBS 0.016896f
C164 VTAIL.n57 VSUBS 0.475254f
C165 VTAIL.n58 VSUBS 0.015957f
C166 VTAIL.t0 VSUBS 0.081527f
C167 VTAIL.n59 VSUBS 0.118393f
C168 VTAIL.n60 VSUBS 0.023894f
C169 VTAIL.n61 VSUBS 0.028287f
C170 VTAIL.n62 VSUBS 0.037717f
C171 VTAIL.n63 VSUBS 0.016896f
C172 VTAIL.n64 VSUBS 0.015957f
C173 VTAIL.n65 VSUBS 0.029695f
C174 VTAIL.n66 VSUBS 0.029695f
C175 VTAIL.n67 VSUBS 0.015957f
C176 VTAIL.n68 VSUBS 0.016896f
C177 VTAIL.n69 VSUBS 0.037717f
C178 VTAIL.n70 VSUBS 0.084025f
C179 VTAIL.n71 VSUBS 0.016896f
C180 VTAIL.n72 VSUBS 0.015957f
C181 VTAIL.n73 VSUBS 0.065394f
C182 VTAIL.n74 VSUBS 0.04183f
C183 VTAIL.n75 VSUBS 1.11321f
C184 VTAIL.n76 VSUBS 0.030491f
C185 VTAIL.n77 VSUBS 0.029695f
C186 VTAIL.n78 VSUBS 0.015957f
C187 VTAIL.n79 VSUBS 0.037717f
C188 VTAIL.n80 VSUBS 0.016896f
C189 VTAIL.n81 VSUBS 0.475254f
C190 VTAIL.n82 VSUBS 0.015957f
C191 VTAIL.t14 VSUBS 0.081527f
C192 VTAIL.n83 VSUBS 0.118393f
C193 VTAIL.n84 VSUBS 0.023894f
C194 VTAIL.n85 VSUBS 0.028287f
C195 VTAIL.n86 VSUBS 0.037717f
C196 VTAIL.n87 VSUBS 0.016896f
C197 VTAIL.n88 VSUBS 0.015957f
C198 VTAIL.n89 VSUBS 0.029695f
C199 VTAIL.n90 VSUBS 0.029695f
C200 VTAIL.n91 VSUBS 0.015957f
C201 VTAIL.n92 VSUBS 0.016896f
C202 VTAIL.n93 VSUBS 0.037717f
C203 VTAIL.n94 VSUBS 0.084025f
C204 VTAIL.n95 VSUBS 0.016896f
C205 VTAIL.n96 VSUBS 0.015957f
C206 VTAIL.n97 VSUBS 0.065394f
C207 VTAIL.n98 VSUBS 0.04183f
C208 VTAIL.n99 VSUBS 1.11321f
C209 VTAIL.t11 VSUBS 0.105129f
C210 VTAIL.t12 VSUBS 0.105129f
C211 VTAIL.n100 VSUBS 0.552776f
C212 VTAIL.n101 VSUBS 0.799494f
C213 VTAIL.n102 VSUBS 0.030491f
C214 VTAIL.n103 VSUBS 0.029695f
C215 VTAIL.n104 VSUBS 0.015957f
C216 VTAIL.n105 VSUBS 0.037717f
C217 VTAIL.n106 VSUBS 0.016896f
C218 VTAIL.n107 VSUBS 0.475254f
C219 VTAIL.n108 VSUBS 0.015957f
C220 VTAIL.t13 VSUBS 0.081527f
C221 VTAIL.n109 VSUBS 0.118393f
C222 VTAIL.n110 VSUBS 0.023894f
C223 VTAIL.n111 VSUBS 0.028287f
C224 VTAIL.n112 VSUBS 0.037717f
C225 VTAIL.n113 VSUBS 0.016896f
C226 VTAIL.n114 VSUBS 0.015957f
C227 VTAIL.n115 VSUBS 0.029695f
C228 VTAIL.n116 VSUBS 0.029695f
C229 VTAIL.n117 VSUBS 0.015957f
C230 VTAIL.n118 VSUBS 0.016896f
C231 VTAIL.n119 VSUBS 0.037717f
C232 VTAIL.n120 VSUBS 0.084025f
C233 VTAIL.n121 VSUBS 0.016896f
C234 VTAIL.n122 VSUBS 0.015957f
C235 VTAIL.n123 VSUBS 0.065394f
C236 VTAIL.n124 VSUBS 0.04183f
C237 VTAIL.n125 VSUBS 0.226864f
C238 VTAIL.n126 VSUBS 0.030491f
C239 VTAIL.n127 VSUBS 0.029695f
C240 VTAIL.n128 VSUBS 0.015957f
C241 VTAIL.n129 VSUBS 0.037717f
C242 VTAIL.n130 VSUBS 0.016896f
C243 VTAIL.n131 VSUBS 0.475254f
C244 VTAIL.n132 VSUBS 0.015957f
C245 VTAIL.t6 VSUBS 0.081527f
C246 VTAIL.n133 VSUBS 0.118393f
C247 VTAIL.n134 VSUBS 0.023894f
C248 VTAIL.n135 VSUBS 0.028287f
C249 VTAIL.n136 VSUBS 0.037717f
C250 VTAIL.n137 VSUBS 0.016896f
C251 VTAIL.n138 VSUBS 0.015957f
C252 VTAIL.n139 VSUBS 0.029695f
C253 VTAIL.n140 VSUBS 0.029695f
C254 VTAIL.n141 VSUBS 0.015957f
C255 VTAIL.n142 VSUBS 0.016896f
C256 VTAIL.n143 VSUBS 0.037717f
C257 VTAIL.n144 VSUBS 0.084025f
C258 VTAIL.n145 VSUBS 0.016896f
C259 VTAIL.n146 VSUBS 0.015957f
C260 VTAIL.n147 VSUBS 0.065394f
C261 VTAIL.n148 VSUBS 0.04183f
C262 VTAIL.n149 VSUBS 0.226864f
C263 VTAIL.t4 VSUBS 0.105129f
C264 VTAIL.t5 VSUBS 0.105129f
C265 VTAIL.n150 VSUBS 0.552776f
C266 VTAIL.n151 VSUBS 0.799494f
C267 VTAIL.n152 VSUBS 0.030491f
C268 VTAIL.n153 VSUBS 0.029695f
C269 VTAIL.n154 VSUBS 0.015957f
C270 VTAIL.n155 VSUBS 0.037717f
C271 VTAIL.n156 VSUBS 0.016896f
C272 VTAIL.n157 VSUBS 0.475254f
C273 VTAIL.n158 VSUBS 0.015957f
C274 VTAIL.t7 VSUBS 0.081527f
C275 VTAIL.n159 VSUBS 0.118393f
C276 VTAIL.n160 VSUBS 0.023894f
C277 VTAIL.n161 VSUBS 0.028287f
C278 VTAIL.n162 VSUBS 0.037717f
C279 VTAIL.n163 VSUBS 0.016896f
C280 VTAIL.n164 VSUBS 0.015957f
C281 VTAIL.n165 VSUBS 0.029695f
C282 VTAIL.n166 VSUBS 0.029695f
C283 VTAIL.n167 VSUBS 0.015957f
C284 VTAIL.n168 VSUBS 0.016896f
C285 VTAIL.n169 VSUBS 0.037717f
C286 VTAIL.n170 VSUBS 0.084025f
C287 VTAIL.n171 VSUBS 0.016896f
C288 VTAIL.n172 VSUBS 0.015957f
C289 VTAIL.n173 VSUBS 0.065394f
C290 VTAIL.n174 VSUBS 0.04183f
C291 VTAIL.n175 VSUBS 1.11321f
C292 VTAIL.n176 VSUBS 0.030491f
C293 VTAIL.n177 VSUBS 0.029695f
C294 VTAIL.n178 VSUBS 0.015957f
C295 VTAIL.n179 VSUBS 0.037717f
C296 VTAIL.n180 VSUBS 0.016896f
C297 VTAIL.n181 VSUBS 0.475254f
C298 VTAIL.n182 VSUBS 0.015957f
C299 VTAIL.t10 VSUBS 0.081527f
C300 VTAIL.n183 VSUBS 0.118393f
C301 VTAIL.n184 VSUBS 0.023894f
C302 VTAIL.n185 VSUBS 0.028287f
C303 VTAIL.n186 VSUBS 0.037717f
C304 VTAIL.n187 VSUBS 0.016896f
C305 VTAIL.n188 VSUBS 0.015957f
C306 VTAIL.n189 VSUBS 0.029695f
C307 VTAIL.n190 VSUBS 0.029695f
C308 VTAIL.n191 VSUBS 0.015957f
C309 VTAIL.n192 VSUBS 0.016896f
C310 VTAIL.n193 VSUBS 0.037717f
C311 VTAIL.n194 VSUBS 0.084025f
C312 VTAIL.n195 VSUBS 0.016896f
C313 VTAIL.n196 VSUBS 0.015957f
C314 VTAIL.n197 VSUBS 0.065394f
C315 VTAIL.n198 VSUBS 0.04183f
C316 VTAIL.n199 VSUBS 1.10764f
C317 VDD2.t0 VSUBS 0.087349f
C318 VDD2.t4 VSUBS 0.087349f
C319 VDD2.n0 VSUBS 0.533472f
C320 VDD2.t3 VSUBS 0.087349f
C321 VDD2.t6 VSUBS 0.087349f
C322 VDD2.n1 VSUBS 0.533472f
C323 VDD2.n2 VSUBS 2.53195f
C324 VDD2.t5 VSUBS 0.087349f
C325 VDD2.t7 VSUBS 0.087349f
C326 VDD2.n3 VSUBS 0.529226f
C327 VDD2.n4 VSUBS 2.14489f
C328 VDD2.t2 VSUBS 0.087349f
C329 VDD2.t1 VSUBS 0.087349f
C330 VDD2.n5 VSUBS 0.533449f
C331 VN.n0 VSUBS 0.048227f
C332 VN.t5 VSUBS 0.891092f
C333 VN.n1 VSUBS 0.05943f
C334 VN.n2 VSUBS 0.048227f
C335 VN.t6 VSUBS 0.891092f
C336 VN.n3 VSUBS 0.070105f
C337 VN.t0 VSUBS 1.06949f
C338 VN.n4 VSUBS 0.46779f
C339 VN.t7 VSUBS 0.891092f
C340 VN.n5 VSUBS 0.45472f
C341 VN.n6 VSUBS 0.063825f
C342 VN.n7 VSUBS 0.305688f
C343 VN.n8 VSUBS 0.048227f
C344 VN.n9 VSUBS 0.048227f
C345 VN.n10 VSUBS 0.070105f
C346 VN.n11 VSUBS 0.063825f
C347 VN.n12 VSUBS 0.365058f
C348 VN.n13 VSUBS 0.070888f
C349 VN.n14 VSUBS 0.048227f
C350 VN.n15 VSUBS 0.048227f
C351 VN.n16 VSUBS 0.048227f
C352 VN.n17 VSUBS 0.080779f
C353 VN.n18 VSUBS 0.056761f
C354 VN.n19 VSUBS 0.462879f
C355 VN.n20 VSUBS 0.04841f
C356 VN.n21 VSUBS 0.048227f
C357 VN.t1 VSUBS 0.891092f
C358 VN.n22 VSUBS 0.05943f
C359 VN.n23 VSUBS 0.048227f
C360 VN.t4 VSUBS 0.891092f
C361 VN.n24 VSUBS 0.070105f
C362 VN.t2 VSUBS 1.06949f
C363 VN.n25 VSUBS 0.46779f
C364 VN.t3 VSUBS 0.891092f
C365 VN.n26 VSUBS 0.45472f
C366 VN.n27 VSUBS 0.063825f
C367 VN.n28 VSUBS 0.305688f
C368 VN.n29 VSUBS 0.048227f
C369 VN.n30 VSUBS 0.048227f
C370 VN.n31 VSUBS 0.070105f
C371 VN.n32 VSUBS 0.063825f
C372 VN.n33 VSUBS 0.365058f
C373 VN.n34 VSUBS 0.070888f
C374 VN.n35 VSUBS 0.048227f
C375 VN.n36 VSUBS 0.048227f
C376 VN.n37 VSUBS 0.048227f
C377 VN.n38 VSUBS 0.080779f
C378 VN.n39 VSUBS 0.056761f
C379 VN.n40 VSUBS 0.462879f
C380 VN.n41 VSUBS 1.90411f
C381 B.n0 VSUBS 0.008134f
C382 B.n1 VSUBS 0.008134f
C383 B.n2 VSUBS 0.012029f
C384 B.n3 VSUBS 0.009218f
C385 B.n4 VSUBS 0.009218f
C386 B.n5 VSUBS 0.009218f
C387 B.n6 VSUBS 0.009218f
C388 B.n7 VSUBS 0.009218f
C389 B.n8 VSUBS 0.009218f
C390 B.n9 VSUBS 0.009218f
C391 B.n10 VSUBS 0.009218f
C392 B.n11 VSUBS 0.009218f
C393 B.n12 VSUBS 0.009218f
C394 B.n13 VSUBS 0.009218f
C395 B.n14 VSUBS 0.009218f
C396 B.n15 VSUBS 0.009218f
C397 B.n16 VSUBS 0.009218f
C398 B.n17 VSUBS 0.009218f
C399 B.n18 VSUBS 0.009218f
C400 B.n19 VSUBS 0.009218f
C401 B.n20 VSUBS 0.020445f
C402 B.n21 VSUBS 0.009218f
C403 B.n22 VSUBS 0.009218f
C404 B.n23 VSUBS 0.009218f
C405 B.n24 VSUBS 0.009218f
C406 B.n25 VSUBS 0.009218f
C407 B.n26 VSUBS 0.009218f
C408 B.n27 VSUBS 0.009218f
C409 B.n28 VSUBS 0.009218f
C410 B.n29 VSUBS 0.009218f
C411 B.t1 VSUBS 0.084803f
C412 B.t2 VSUBS 0.104541f
C413 B.t0 VSUBS 0.438975f
C414 B.n30 VSUBS 0.188501f
C415 B.n31 VSUBS 0.161175f
C416 B.n32 VSUBS 0.021357f
C417 B.n33 VSUBS 0.009218f
C418 B.n34 VSUBS 0.009218f
C419 B.n35 VSUBS 0.009218f
C420 B.n36 VSUBS 0.009218f
C421 B.n37 VSUBS 0.009218f
C422 B.t7 VSUBS 0.084804f
C423 B.t8 VSUBS 0.104543f
C424 B.t6 VSUBS 0.438975f
C425 B.n38 VSUBS 0.1885f
C426 B.n39 VSUBS 0.161173f
C427 B.n40 VSUBS 0.009218f
C428 B.n41 VSUBS 0.009218f
C429 B.n42 VSUBS 0.009218f
C430 B.n43 VSUBS 0.009218f
C431 B.n44 VSUBS 0.009218f
C432 B.n45 VSUBS 0.009218f
C433 B.n46 VSUBS 0.009218f
C434 B.n47 VSUBS 0.009218f
C435 B.n48 VSUBS 0.009218f
C436 B.n49 VSUBS 0.019139f
C437 B.n50 VSUBS 0.009218f
C438 B.n51 VSUBS 0.009218f
C439 B.n52 VSUBS 0.009218f
C440 B.n53 VSUBS 0.009218f
C441 B.n54 VSUBS 0.009218f
C442 B.n55 VSUBS 0.009218f
C443 B.n56 VSUBS 0.009218f
C444 B.n57 VSUBS 0.009218f
C445 B.n58 VSUBS 0.009218f
C446 B.n59 VSUBS 0.009218f
C447 B.n60 VSUBS 0.009218f
C448 B.n61 VSUBS 0.009218f
C449 B.n62 VSUBS 0.009218f
C450 B.n63 VSUBS 0.009218f
C451 B.n64 VSUBS 0.009218f
C452 B.n65 VSUBS 0.009218f
C453 B.n66 VSUBS 0.009218f
C454 B.n67 VSUBS 0.009218f
C455 B.n68 VSUBS 0.009218f
C456 B.n69 VSUBS 0.009218f
C457 B.n70 VSUBS 0.009218f
C458 B.n71 VSUBS 0.009218f
C459 B.n72 VSUBS 0.009218f
C460 B.n73 VSUBS 0.009218f
C461 B.n74 VSUBS 0.009218f
C462 B.n75 VSUBS 0.009218f
C463 B.n76 VSUBS 0.009218f
C464 B.n77 VSUBS 0.009218f
C465 B.n78 VSUBS 0.009218f
C466 B.n79 VSUBS 0.009218f
C467 B.n80 VSUBS 0.009218f
C468 B.n81 VSUBS 0.009218f
C469 B.n82 VSUBS 0.009218f
C470 B.n83 VSUBS 0.009218f
C471 B.n84 VSUBS 0.009218f
C472 B.n85 VSUBS 0.009218f
C473 B.n86 VSUBS 0.0192f
C474 B.n87 VSUBS 0.009218f
C475 B.n88 VSUBS 0.009218f
C476 B.n89 VSUBS 0.009218f
C477 B.n90 VSUBS 0.009218f
C478 B.n91 VSUBS 0.009218f
C479 B.n92 VSUBS 0.009218f
C480 B.n93 VSUBS 0.009218f
C481 B.n94 VSUBS 0.009218f
C482 B.n95 VSUBS 0.009218f
C483 B.t11 VSUBS 0.084804f
C484 B.t10 VSUBS 0.104543f
C485 B.t9 VSUBS 0.438975f
C486 B.n96 VSUBS 0.1885f
C487 B.n97 VSUBS 0.161173f
C488 B.n98 VSUBS 0.021357f
C489 B.n99 VSUBS 0.009218f
C490 B.n100 VSUBS 0.009218f
C491 B.n101 VSUBS 0.009218f
C492 B.n102 VSUBS 0.009218f
C493 B.n103 VSUBS 0.009218f
C494 B.t5 VSUBS 0.084803f
C495 B.t4 VSUBS 0.104541f
C496 B.t3 VSUBS 0.438975f
C497 B.n104 VSUBS 0.188501f
C498 B.n105 VSUBS 0.161175f
C499 B.n106 VSUBS 0.009218f
C500 B.n107 VSUBS 0.009218f
C501 B.n108 VSUBS 0.009218f
C502 B.n109 VSUBS 0.009218f
C503 B.n110 VSUBS 0.009218f
C504 B.n111 VSUBS 0.009218f
C505 B.n112 VSUBS 0.009218f
C506 B.n113 VSUBS 0.009218f
C507 B.n114 VSUBS 0.009218f
C508 B.n115 VSUBS 0.019139f
C509 B.n116 VSUBS 0.009218f
C510 B.n117 VSUBS 0.009218f
C511 B.n118 VSUBS 0.009218f
C512 B.n119 VSUBS 0.009218f
C513 B.n120 VSUBS 0.009218f
C514 B.n121 VSUBS 0.009218f
C515 B.n122 VSUBS 0.009218f
C516 B.n123 VSUBS 0.009218f
C517 B.n124 VSUBS 0.009218f
C518 B.n125 VSUBS 0.009218f
C519 B.n126 VSUBS 0.009218f
C520 B.n127 VSUBS 0.009218f
C521 B.n128 VSUBS 0.009218f
C522 B.n129 VSUBS 0.009218f
C523 B.n130 VSUBS 0.009218f
C524 B.n131 VSUBS 0.009218f
C525 B.n132 VSUBS 0.009218f
C526 B.n133 VSUBS 0.009218f
C527 B.n134 VSUBS 0.009218f
C528 B.n135 VSUBS 0.009218f
C529 B.n136 VSUBS 0.009218f
C530 B.n137 VSUBS 0.009218f
C531 B.n138 VSUBS 0.009218f
C532 B.n139 VSUBS 0.009218f
C533 B.n140 VSUBS 0.009218f
C534 B.n141 VSUBS 0.009218f
C535 B.n142 VSUBS 0.009218f
C536 B.n143 VSUBS 0.009218f
C537 B.n144 VSUBS 0.009218f
C538 B.n145 VSUBS 0.009218f
C539 B.n146 VSUBS 0.009218f
C540 B.n147 VSUBS 0.009218f
C541 B.n148 VSUBS 0.009218f
C542 B.n149 VSUBS 0.009218f
C543 B.n150 VSUBS 0.009218f
C544 B.n151 VSUBS 0.009218f
C545 B.n152 VSUBS 0.009218f
C546 B.n153 VSUBS 0.009218f
C547 B.n154 VSUBS 0.009218f
C548 B.n155 VSUBS 0.009218f
C549 B.n156 VSUBS 0.009218f
C550 B.n157 VSUBS 0.009218f
C551 B.n158 VSUBS 0.009218f
C552 B.n159 VSUBS 0.009218f
C553 B.n160 VSUBS 0.009218f
C554 B.n161 VSUBS 0.009218f
C555 B.n162 VSUBS 0.009218f
C556 B.n163 VSUBS 0.009218f
C557 B.n164 VSUBS 0.009218f
C558 B.n165 VSUBS 0.009218f
C559 B.n166 VSUBS 0.009218f
C560 B.n167 VSUBS 0.009218f
C561 B.n168 VSUBS 0.009218f
C562 B.n169 VSUBS 0.009218f
C563 B.n170 VSUBS 0.009218f
C564 B.n171 VSUBS 0.009218f
C565 B.n172 VSUBS 0.009218f
C566 B.n173 VSUBS 0.009218f
C567 B.n174 VSUBS 0.009218f
C568 B.n175 VSUBS 0.009218f
C569 B.n176 VSUBS 0.009218f
C570 B.n177 VSUBS 0.009218f
C571 B.n178 VSUBS 0.009218f
C572 B.n179 VSUBS 0.009218f
C573 B.n180 VSUBS 0.009218f
C574 B.n181 VSUBS 0.009218f
C575 B.n182 VSUBS 0.009218f
C576 B.n183 VSUBS 0.009218f
C577 B.n184 VSUBS 0.019139f
C578 B.n185 VSUBS 0.020445f
C579 B.n186 VSUBS 0.020445f
C580 B.n187 VSUBS 0.009218f
C581 B.n188 VSUBS 0.009218f
C582 B.n189 VSUBS 0.009218f
C583 B.n190 VSUBS 0.009218f
C584 B.n191 VSUBS 0.009218f
C585 B.n192 VSUBS 0.009218f
C586 B.n193 VSUBS 0.009218f
C587 B.n194 VSUBS 0.009218f
C588 B.n195 VSUBS 0.009218f
C589 B.n196 VSUBS 0.009218f
C590 B.n197 VSUBS 0.009218f
C591 B.n198 VSUBS 0.009218f
C592 B.n199 VSUBS 0.009218f
C593 B.n200 VSUBS 0.009218f
C594 B.n201 VSUBS 0.009218f
C595 B.n202 VSUBS 0.009218f
C596 B.n203 VSUBS 0.009218f
C597 B.n204 VSUBS 0.009218f
C598 B.n205 VSUBS 0.009218f
C599 B.n206 VSUBS 0.009218f
C600 B.n207 VSUBS 0.009218f
C601 B.n208 VSUBS 0.009218f
C602 B.n209 VSUBS 0.009218f
C603 B.n210 VSUBS 0.009218f
C604 B.n211 VSUBS 0.009218f
C605 B.n212 VSUBS 0.009218f
C606 B.n213 VSUBS 0.009218f
C607 B.n214 VSUBS 0.006371f
C608 B.n215 VSUBS 0.021357f
C609 B.n216 VSUBS 0.007456f
C610 B.n217 VSUBS 0.009218f
C611 B.n218 VSUBS 0.009218f
C612 B.n219 VSUBS 0.009218f
C613 B.n220 VSUBS 0.009218f
C614 B.n221 VSUBS 0.009218f
C615 B.n222 VSUBS 0.009218f
C616 B.n223 VSUBS 0.009218f
C617 B.n224 VSUBS 0.009218f
C618 B.n225 VSUBS 0.009218f
C619 B.n226 VSUBS 0.009218f
C620 B.n227 VSUBS 0.009218f
C621 B.n228 VSUBS 0.007456f
C622 B.n229 VSUBS 0.009218f
C623 B.n230 VSUBS 0.009218f
C624 B.n231 VSUBS 0.006371f
C625 B.n232 VSUBS 0.009218f
C626 B.n233 VSUBS 0.009218f
C627 B.n234 VSUBS 0.009218f
C628 B.n235 VSUBS 0.009218f
C629 B.n236 VSUBS 0.009218f
C630 B.n237 VSUBS 0.009218f
C631 B.n238 VSUBS 0.009218f
C632 B.n239 VSUBS 0.009218f
C633 B.n240 VSUBS 0.009218f
C634 B.n241 VSUBS 0.009218f
C635 B.n242 VSUBS 0.009218f
C636 B.n243 VSUBS 0.009218f
C637 B.n244 VSUBS 0.009218f
C638 B.n245 VSUBS 0.009218f
C639 B.n246 VSUBS 0.009218f
C640 B.n247 VSUBS 0.009218f
C641 B.n248 VSUBS 0.009218f
C642 B.n249 VSUBS 0.009218f
C643 B.n250 VSUBS 0.009218f
C644 B.n251 VSUBS 0.009218f
C645 B.n252 VSUBS 0.009218f
C646 B.n253 VSUBS 0.009218f
C647 B.n254 VSUBS 0.009218f
C648 B.n255 VSUBS 0.009218f
C649 B.n256 VSUBS 0.009218f
C650 B.n257 VSUBS 0.009218f
C651 B.n258 VSUBS 0.009218f
C652 B.n259 VSUBS 0.020445f
C653 B.n260 VSUBS 0.019139f
C654 B.n261 VSUBS 0.020384f
C655 B.n262 VSUBS 0.009218f
C656 B.n263 VSUBS 0.009218f
C657 B.n264 VSUBS 0.009218f
C658 B.n265 VSUBS 0.009218f
C659 B.n266 VSUBS 0.009218f
C660 B.n267 VSUBS 0.009218f
C661 B.n268 VSUBS 0.009218f
C662 B.n269 VSUBS 0.009218f
C663 B.n270 VSUBS 0.009218f
C664 B.n271 VSUBS 0.009218f
C665 B.n272 VSUBS 0.009218f
C666 B.n273 VSUBS 0.009218f
C667 B.n274 VSUBS 0.009218f
C668 B.n275 VSUBS 0.009218f
C669 B.n276 VSUBS 0.009218f
C670 B.n277 VSUBS 0.009218f
C671 B.n278 VSUBS 0.009218f
C672 B.n279 VSUBS 0.009218f
C673 B.n280 VSUBS 0.009218f
C674 B.n281 VSUBS 0.009218f
C675 B.n282 VSUBS 0.009218f
C676 B.n283 VSUBS 0.009218f
C677 B.n284 VSUBS 0.009218f
C678 B.n285 VSUBS 0.009218f
C679 B.n286 VSUBS 0.009218f
C680 B.n287 VSUBS 0.009218f
C681 B.n288 VSUBS 0.009218f
C682 B.n289 VSUBS 0.009218f
C683 B.n290 VSUBS 0.009218f
C684 B.n291 VSUBS 0.009218f
C685 B.n292 VSUBS 0.009218f
C686 B.n293 VSUBS 0.009218f
C687 B.n294 VSUBS 0.009218f
C688 B.n295 VSUBS 0.009218f
C689 B.n296 VSUBS 0.009218f
C690 B.n297 VSUBS 0.009218f
C691 B.n298 VSUBS 0.009218f
C692 B.n299 VSUBS 0.009218f
C693 B.n300 VSUBS 0.009218f
C694 B.n301 VSUBS 0.009218f
C695 B.n302 VSUBS 0.009218f
C696 B.n303 VSUBS 0.009218f
C697 B.n304 VSUBS 0.009218f
C698 B.n305 VSUBS 0.009218f
C699 B.n306 VSUBS 0.009218f
C700 B.n307 VSUBS 0.009218f
C701 B.n308 VSUBS 0.009218f
C702 B.n309 VSUBS 0.009218f
C703 B.n310 VSUBS 0.009218f
C704 B.n311 VSUBS 0.009218f
C705 B.n312 VSUBS 0.009218f
C706 B.n313 VSUBS 0.009218f
C707 B.n314 VSUBS 0.009218f
C708 B.n315 VSUBS 0.009218f
C709 B.n316 VSUBS 0.009218f
C710 B.n317 VSUBS 0.009218f
C711 B.n318 VSUBS 0.009218f
C712 B.n319 VSUBS 0.009218f
C713 B.n320 VSUBS 0.009218f
C714 B.n321 VSUBS 0.009218f
C715 B.n322 VSUBS 0.009218f
C716 B.n323 VSUBS 0.009218f
C717 B.n324 VSUBS 0.009218f
C718 B.n325 VSUBS 0.009218f
C719 B.n326 VSUBS 0.009218f
C720 B.n327 VSUBS 0.009218f
C721 B.n328 VSUBS 0.009218f
C722 B.n329 VSUBS 0.009218f
C723 B.n330 VSUBS 0.009218f
C724 B.n331 VSUBS 0.009218f
C725 B.n332 VSUBS 0.009218f
C726 B.n333 VSUBS 0.009218f
C727 B.n334 VSUBS 0.009218f
C728 B.n335 VSUBS 0.009218f
C729 B.n336 VSUBS 0.009218f
C730 B.n337 VSUBS 0.009218f
C731 B.n338 VSUBS 0.009218f
C732 B.n339 VSUBS 0.009218f
C733 B.n340 VSUBS 0.009218f
C734 B.n341 VSUBS 0.009218f
C735 B.n342 VSUBS 0.009218f
C736 B.n343 VSUBS 0.009218f
C737 B.n344 VSUBS 0.009218f
C738 B.n345 VSUBS 0.009218f
C739 B.n346 VSUBS 0.009218f
C740 B.n347 VSUBS 0.009218f
C741 B.n348 VSUBS 0.009218f
C742 B.n349 VSUBS 0.009218f
C743 B.n350 VSUBS 0.009218f
C744 B.n351 VSUBS 0.009218f
C745 B.n352 VSUBS 0.009218f
C746 B.n353 VSUBS 0.009218f
C747 B.n354 VSUBS 0.009218f
C748 B.n355 VSUBS 0.009218f
C749 B.n356 VSUBS 0.009218f
C750 B.n357 VSUBS 0.009218f
C751 B.n358 VSUBS 0.009218f
C752 B.n359 VSUBS 0.009218f
C753 B.n360 VSUBS 0.009218f
C754 B.n361 VSUBS 0.009218f
C755 B.n362 VSUBS 0.009218f
C756 B.n363 VSUBS 0.009218f
C757 B.n364 VSUBS 0.009218f
C758 B.n365 VSUBS 0.009218f
C759 B.n366 VSUBS 0.009218f
C760 B.n367 VSUBS 0.009218f
C761 B.n368 VSUBS 0.009218f
C762 B.n369 VSUBS 0.009218f
C763 B.n370 VSUBS 0.019139f
C764 B.n371 VSUBS 0.020445f
C765 B.n372 VSUBS 0.020445f
C766 B.n373 VSUBS 0.009218f
C767 B.n374 VSUBS 0.009218f
C768 B.n375 VSUBS 0.009218f
C769 B.n376 VSUBS 0.009218f
C770 B.n377 VSUBS 0.009218f
C771 B.n378 VSUBS 0.009218f
C772 B.n379 VSUBS 0.009218f
C773 B.n380 VSUBS 0.009218f
C774 B.n381 VSUBS 0.009218f
C775 B.n382 VSUBS 0.009218f
C776 B.n383 VSUBS 0.009218f
C777 B.n384 VSUBS 0.009218f
C778 B.n385 VSUBS 0.009218f
C779 B.n386 VSUBS 0.009218f
C780 B.n387 VSUBS 0.009218f
C781 B.n388 VSUBS 0.009218f
C782 B.n389 VSUBS 0.009218f
C783 B.n390 VSUBS 0.009218f
C784 B.n391 VSUBS 0.009218f
C785 B.n392 VSUBS 0.009218f
C786 B.n393 VSUBS 0.009218f
C787 B.n394 VSUBS 0.009218f
C788 B.n395 VSUBS 0.009218f
C789 B.n396 VSUBS 0.009218f
C790 B.n397 VSUBS 0.009218f
C791 B.n398 VSUBS 0.009218f
C792 B.n399 VSUBS 0.009218f
C793 B.n400 VSUBS 0.006371f
C794 B.n401 VSUBS 0.021357f
C795 B.n402 VSUBS 0.007456f
C796 B.n403 VSUBS 0.009218f
C797 B.n404 VSUBS 0.009218f
C798 B.n405 VSUBS 0.009218f
C799 B.n406 VSUBS 0.009218f
C800 B.n407 VSUBS 0.009218f
C801 B.n408 VSUBS 0.009218f
C802 B.n409 VSUBS 0.009218f
C803 B.n410 VSUBS 0.009218f
C804 B.n411 VSUBS 0.009218f
C805 B.n412 VSUBS 0.009218f
C806 B.n413 VSUBS 0.009218f
C807 B.n414 VSUBS 0.007456f
C808 B.n415 VSUBS 0.009218f
C809 B.n416 VSUBS 0.009218f
C810 B.n417 VSUBS 0.006371f
C811 B.n418 VSUBS 0.009218f
C812 B.n419 VSUBS 0.009218f
C813 B.n420 VSUBS 0.009218f
C814 B.n421 VSUBS 0.009218f
C815 B.n422 VSUBS 0.009218f
C816 B.n423 VSUBS 0.009218f
C817 B.n424 VSUBS 0.009218f
C818 B.n425 VSUBS 0.009218f
C819 B.n426 VSUBS 0.009218f
C820 B.n427 VSUBS 0.009218f
C821 B.n428 VSUBS 0.009218f
C822 B.n429 VSUBS 0.009218f
C823 B.n430 VSUBS 0.009218f
C824 B.n431 VSUBS 0.009218f
C825 B.n432 VSUBS 0.009218f
C826 B.n433 VSUBS 0.009218f
C827 B.n434 VSUBS 0.009218f
C828 B.n435 VSUBS 0.009218f
C829 B.n436 VSUBS 0.009218f
C830 B.n437 VSUBS 0.009218f
C831 B.n438 VSUBS 0.009218f
C832 B.n439 VSUBS 0.009218f
C833 B.n440 VSUBS 0.009218f
C834 B.n441 VSUBS 0.009218f
C835 B.n442 VSUBS 0.009218f
C836 B.n443 VSUBS 0.009218f
C837 B.n444 VSUBS 0.009218f
C838 B.n445 VSUBS 0.020445f
C839 B.n446 VSUBS 0.019139f
C840 B.n447 VSUBS 0.019139f
C841 B.n448 VSUBS 0.009218f
C842 B.n449 VSUBS 0.009218f
C843 B.n450 VSUBS 0.009218f
C844 B.n451 VSUBS 0.009218f
C845 B.n452 VSUBS 0.009218f
C846 B.n453 VSUBS 0.009218f
C847 B.n454 VSUBS 0.009218f
C848 B.n455 VSUBS 0.009218f
C849 B.n456 VSUBS 0.009218f
C850 B.n457 VSUBS 0.009218f
C851 B.n458 VSUBS 0.009218f
C852 B.n459 VSUBS 0.009218f
C853 B.n460 VSUBS 0.009218f
C854 B.n461 VSUBS 0.009218f
C855 B.n462 VSUBS 0.009218f
C856 B.n463 VSUBS 0.009218f
C857 B.n464 VSUBS 0.009218f
C858 B.n465 VSUBS 0.009218f
C859 B.n466 VSUBS 0.009218f
C860 B.n467 VSUBS 0.009218f
C861 B.n468 VSUBS 0.009218f
C862 B.n469 VSUBS 0.009218f
C863 B.n470 VSUBS 0.009218f
C864 B.n471 VSUBS 0.009218f
C865 B.n472 VSUBS 0.009218f
C866 B.n473 VSUBS 0.009218f
C867 B.n474 VSUBS 0.009218f
C868 B.n475 VSUBS 0.009218f
C869 B.n476 VSUBS 0.009218f
C870 B.n477 VSUBS 0.009218f
C871 B.n478 VSUBS 0.009218f
C872 B.n479 VSUBS 0.009218f
C873 B.n480 VSUBS 0.009218f
C874 B.n481 VSUBS 0.009218f
C875 B.n482 VSUBS 0.009218f
C876 B.n483 VSUBS 0.009218f
C877 B.n484 VSUBS 0.009218f
C878 B.n485 VSUBS 0.009218f
C879 B.n486 VSUBS 0.009218f
C880 B.n487 VSUBS 0.009218f
C881 B.n488 VSUBS 0.009218f
C882 B.n489 VSUBS 0.009218f
C883 B.n490 VSUBS 0.009218f
C884 B.n491 VSUBS 0.009218f
C885 B.n492 VSUBS 0.009218f
C886 B.n493 VSUBS 0.009218f
C887 B.n494 VSUBS 0.009218f
C888 B.n495 VSUBS 0.009218f
C889 B.n496 VSUBS 0.009218f
C890 B.n497 VSUBS 0.009218f
C891 B.n498 VSUBS 0.009218f
C892 B.n499 VSUBS 0.012029f
C893 B.n500 VSUBS 0.012814f
C894 B.n501 VSUBS 0.025482f
.ends

