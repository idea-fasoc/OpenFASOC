* NGSPICE file created from diff_pair_sample_0694.ext - technology: sky130A

.subckt diff_pair_sample_0694 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X1 VDD2.t9 VN.t0 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=1.2792 ps=7.34 w=3.28 l=0.84
X2 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X3 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X4 VTAIL.t8 VN.t3 VDD2.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X5 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0 ps=0 w=3.28 l=0.84
X6 VDD2.t5 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0.5412 ps=3.61 w=3.28 l=0.84
X7 VDD1.t8 VP.t1 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0.5412 ps=3.61 w=3.28 l=0.84
X8 VDD1.t7 VP.t2 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0.5412 ps=3.61 w=3.28 l=0.84
X9 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0 ps=0 w=3.28 l=0.84
X10 VTAIL.t15 VP.t3 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X11 VDD2.t4 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X12 VDD2.t3 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0.5412 ps=3.61 w=3.28 l=0.84
X13 VDD2.t2 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=1.2792 ps=7.34 w=3.28 l=0.84
X14 VTAIL.t13 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X15 VTAIL.t17 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X16 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0 ps=0 w=3.28 l=0.84
X17 VDD1.t3 VP.t6 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X18 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.2792 pd=7.34 as=0 ps=0 w=3.28 l=0.84
X19 VTAIL.t16 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X20 VDD1.t1 VP.t8 VTAIL.t10 B.t23 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=1.2792 ps=7.34 w=3.28 l=0.84
X21 VTAIL.t1 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
X22 VDD1.t0 VP.t9 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=1.2792 ps=7.34 w=3.28 l=0.84
X23 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5412 pd=3.61 as=0.5412 ps=3.61 w=3.28 l=0.84
R0 VP.n10 VP.t1 165.869
R1 VP.n40 VP.n39 161.3
R2 VP.n11 VP.n8 161.3
R3 VP.n13 VP.n12 161.3
R4 VP.n15 VP.n7 161.3
R5 VP.n17 VP.n16 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n20 VP.n5 161.3
R8 VP.n22 VP.n21 161.3
R9 VP.n38 VP.n0 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n35 VP.n34 161.3
R12 VP.n33 VP.n2 161.3
R13 VP.n31 VP.n30 161.3
R14 VP.n29 VP.n3 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n25 VP.n4 161.3
R17 VP.n24 VP.n23 161.3
R18 VP.n24 VP.t2 140.87
R19 VP.n39 VP.t9 140.87
R20 VP.n21 VP.t8 140.87
R21 VP.n26 VP.t5 94.1053
R22 VP.n32 VP.t6 94.1053
R23 VP.n1 VP.t7 94.1053
R24 VP.n6 VP.t3 94.1053
R25 VP.n14 VP.t0 94.1053
R26 VP.n9 VP.t4 94.1053
R27 VP.n31 VP.n3 56.5617
R28 VP.n34 VP.n33 56.5617
R29 VP.n16 VP.n15 56.5617
R30 VP.n13 VP.n8 56.5617
R31 VP.n11 VP.n10 42.2591
R32 VP.n27 VP.n25 40.0926
R33 VP.n38 VP.n37 40.0926
R34 VP.n20 VP.n19 40.0926
R35 VP.n23 VP.n22 36.9967
R36 VP.n10 VP.n9 32.8395
R37 VP.n25 VP.n24 24.8308
R38 VP.n39 VP.n38 24.8308
R39 VP.n21 VP.n20 24.8308
R40 VP.n26 VP.n3 20.6576
R41 VP.n34 VP.n1 20.6576
R42 VP.n16 VP.n6 20.6576
R43 VP.n9 VP.n8 20.6576
R44 VP.n32 VP.n31 12.2964
R45 VP.n33 VP.n32 12.2964
R46 VP.n14 VP.n13 12.2964
R47 VP.n15 VP.n14 12.2964
R48 VP.n27 VP.n26 3.93519
R49 VP.n37 VP.n1 3.93519
R50 VP.n19 VP.n6 3.93519
R51 VP.n12 VP.n11 0.189894
R52 VP.n12 VP.n7 0.189894
R53 VP.n17 VP.n7 0.189894
R54 VP.n18 VP.n17 0.189894
R55 VP.n18 VP.n5 0.189894
R56 VP.n22 VP.n5 0.189894
R57 VP.n23 VP.n4 0.189894
R58 VP.n28 VP.n4 0.189894
R59 VP.n29 VP.n28 0.189894
R60 VP.n30 VP.n29 0.189894
R61 VP.n30 VP.n2 0.189894
R62 VP.n35 VP.n2 0.189894
R63 VP.n36 VP.n35 0.189894
R64 VP.n36 VP.n0 0.189894
R65 VP.n40 VP.n0 0.189894
R66 VP VP.n40 0.0516364
R67 VTAIL.n72 VTAIL.n62 289.615
R68 VTAIL.n12 VTAIL.n2 289.615
R69 VTAIL.n56 VTAIL.n46 289.615
R70 VTAIL.n36 VTAIL.n26 289.615
R71 VTAIL.n66 VTAIL.n65 185
R72 VTAIL.n71 VTAIL.n70 185
R73 VTAIL.n73 VTAIL.n72 185
R74 VTAIL.n6 VTAIL.n5 185
R75 VTAIL.n11 VTAIL.n10 185
R76 VTAIL.n13 VTAIL.n12 185
R77 VTAIL.n57 VTAIL.n56 185
R78 VTAIL.n55 VTAIL.n54 185
R79 VTAIL.n50 VTAIL.n49 185
R80 VTAIL.n37 VTAIL.n36 185
R81 VTAIL.n35 VTAIL.n34 185
R82 VTAIL.n30 VTAIL.n29 185
R83 VTAIL.n67 VTAIL.t19 148.606
R84 VTAIL.n7 VTAIL.t18 148.606
R85 VTAIL.n51 VTAIL.t10 148.606
R86 VTAIL.n31 VTAIL.t3 148.606
R87 VTAIL.n71 VTAIL.n65 104.615
R88 VTAIL.n72 VTAIL.n71 104.615
R89 VTAIL.n11 VTAIL.n5 104.615
R90 VTAIL.n12 VTAIL.n11 104.615
R91 VTAIL.n56 VTAIL.n55 104.615
R92 VTAIL.n55 VTAIL.n49 104.615
R93 VTAIL.n36 VTAIL.n35 104.615
R94 VTAIL.n35 VTAIL.n29 104.615
R95 VTAIL.n45 VTAIL.n44 64.1734
R96 VTAIL.n43 VTAIL.n42 64.1734
R97 VTAIL.n25 VTAIL.n24 64.1734
R98 VTAIL.n23 VTAIL.n22 64.1734
R99 VTAIL.n79 VTAIL.n78 64.1733
R100 VTAIL.n1 VTAIL.n0 64.1733
R101 VTAIL.n19 VTAIL.n18 64.1733
R102 VTAIL.n21 VTAIL.n20 64.1733
R103 VTAIL.t19 VTAIL.n65 52.3082
R104 VTAIL.t18 VTAIL.n5 52.3082
R105 VTAIL.t10 VTAIL.n49 52.3082
R106 VTAIL.t3 VTAIL.n29 52.3082
R107 VTAIL.n77 VTAIL.n76 35.2884
R108 VTAIL.n17 VTAIL.n16 35.2884
R109 VTAIL.n61 VTAIL.n60 35.2884
R110 VTAIL.n41 VTAIL.n40 35.2884
R111 VTAIL.n23 VTAIL.n21 17.2117
R112 VTAIL.n77 VTAIL.n61 16.2031
R113 VTAIL.n67 VTAIL.n66 15.5966
R114 VTAIL.n7 VTAIL.n6 15.5966
R115 VTAIL.n51 VTAIL.n50 15.5966
R116 VTAIL.n31 VTAIL.n30 15.5966
R117 VTAIL.n70 VTAIL.n69 12.8005
R118 VTAIL.n10 VTAIL.n9 12.8005
R119 VTAIL.n54 VTAIL.n53 12.8005
R120 VTAIL.n34 VTAIL.n33 12.8005
R121 VTAIL.n73 VTAIL.n64 12.0247
R122 VTAIL.n13 VTAIL.n4 12.0247
R123 VTAIL.n57 VTAIL.n48 12.0247
R124 VTAIL.n37 VTAIL.n28 12.0247
R125 VTAIL.n74 VTAIL.n62 11.249
R126 VTAIL.n14 VTAIL.n2 11.249
R127 VTAIL.n58 VTAIL.n46 11.249
R128 VTAIL.n38 VTAIL.n26 11.249
R129 VTAIL.n76 VTAIL.n75 9.45567
R130 VTAIL.n16 VTAIL.n15 9.45567
R131 VTAIL.n60 VTAIL.n59 9.45567
R132 VTAIL.n40 VTAIL.n39 9.45567
R133 VTAIL.n75 VTAIL.n74 9.3005
R134 VTAIL.n64 VTAIL.n63 9.3005
R135 VTAIL.n69 VTAIL.n68 9.3005
R136 VTAIL.n15 VTAIL.n14 9.3005
R137 VTAIL.n4 VTAIL.n3 9.3005
R138 VTAIL.n9 VTAIL.n8 9.3005
R139 VTAIL.n59 VTAIL.n58 9.3005
R140 VTAIL.n48 VTAIL.n47 9.3005
R141 VTAIL.n53 VTAIL.n52 9.3005
R142 VTAIL.n39 VTAIL.n38 9.3005
R143 VTAIL.n28 VTAIL.n27 9.3005
R144 VTAIL.n33 VTAIL.n32 9.3005
R145 VTAIL.n78 VTAIL.t6 6.03709
R146 VTAIL.n78 VTAIL.t2 6.03709
R147 VTAIL.n0 VTAIL.t4 6.03709
R148 VTAIL.n0 VTAIL.t8 6.03709
R149 VTAIL.n18 VTAIL.t11 6.03709
R150 VTAIL.n18 VTAIL.t16 6.03709
R151 VTAIL.n20 VTAIL.t9 6.03709
R152 VTAIL.n20 VTAIL.t17 6.03709
R153 VTAIL.n44 VTAIL.t14 6.03709
R154 VTAIL.n44 VTAIL.t15 6.03709
R155 VTAIL.n42 VTAIL.t12 6.03709
R156 VTAIL.n42 VTAIL.t13 6.03709
R157 VTAIL.n24 VTAIL.t5 6.03709
R158 VTAIL.n24 VTAIL.t0 6.03709
R159 VTAIL.n22 VTAIL.t7 6.03709
R160 VTAIL.n22 VTAIL.t1 6.03709
R161 VTAIL.n68 VTAIL.n67 4.46457
R162 VTAIL.n8 VTAIL.n7 4.46457
R163 VTAIL.n52 VTAIL.n51 4.46457
R164 VTAIL.n32 VTAIL.n31 4.46457
R165 VTAIL.n76 VTAIL.n62 2.71565
R166 VTAIL.n16 VTAIL.n2 2.71565
R167 VTAIL.n60 VTAIL.n46 2.71565
R168 VTAIL.n40 VTAIL.n26 2.71565
R169 VTAIL.n74 VTAIL.n73 1.93989
R170 VTAIL.n14 VTAIL.n13 1.93989
R171 VTAIL.n58 VTAIL.n57 1.93989
R172 VTAIL.n38 VTAIL.n37 1.93989
R173 VTAIL.n70 VTAIL.n64 1.16414
R174 VTAIL.n10 VTAIL.n4 1.16414
R175 VTAIL.n54 VTAIL.n48 1.16414
R176 VTAIL.n34 VTAIL.n28 1.16414
R177 VTAIL.n25 VTAIL.n23 1.00912
R178 VTAIL.n41 VTAIL.n25 1.00912
R179 VTAIL.n45 VTAIL.n43 1.00912
R180 VTAIL.n61 VTAIL.n45 1.00912
R181 VTAIL.n21 VTAIL.n19 1.00912
R182 VTAIL.n19 VTAIL.n17 1.00912
R183 VTAIL.n79 VTAIL.n77 1.00912
R184 VTAIL.n43 VTAIL.n41 0.974638
R185 VTAIL.n17 VTAIL.n1 0.974638
R186 VTAIL VTAIL.n1 0.815155
R187 VTAIL.n69 VTAIL.n66 0.388379
R188 VTAIL.n9 VTAIL.n6 0.388379
R189 VTAIL.n53 VTAIL.n50 0.388379
R190 VTAIL.n33 VTAIL.n30 0.388379
R191 VTAIL VTAIL.n79 0.194466
R192 VTAIL.n68 VTAIL.n63 0.155672
R193 VTAIL.n75 VTAIL.n63 0.155672
R194 VTAIL.n8 VTAIL.n3 0.155672
R195 VTAIL.n15 VTAIL.n3 0.155672
R196 VTAIL.n59 VTAIL.n47 0.155672
R197 VTAIL.n52 VTAIL.n47 0.155672
R198 VTAIL.n39 VTAIL.n27 0.155672
R199 VTAIL.n32 VTAIL.n27 0.155672
R200 VDD1.n10 VDD1.n0 289.615
R201 VDD1.n27 VDD1.n17 289.615
R202 VDD1.n11 VDD1.n10 185
R203 VDD1.n9 VDD1.n8 185
R204 VDD1.n4 VDD1.n3 185
R205 VDD1.n21 VDD1.n20 185
R206 VDD1.n26 VDD1.n25 185
R207 VDD1.n28 VDD1.n27 185
R208 VDD1.n5 VDD1.t8 148.606
R209 VDD1.n22 VDD1.t7 148.606
R210 VDD1.n10 VDD1.n9 104.615
R211 VDD1.n9 VDD1.n3 104.615
R212 VDD1.n26 VDD1.n20 104.615
R213 VDD1.n27 VDD1.n26 104.615
R214 VDD1.n35 VDD1.n34 81.5532
R215 VDD1.n16 VDD1.n15 80.8522
R216 VDD1.n37 VDD1.n36 80.8521
R217 VDD1.n33 VDD1.n32 80.8521
R218 VDD1.n16 VDD1.n14 52.9758
R219 VDD1.n33 VDD1.n31 52.9758
R220 VDD1.t8 VDD1.n3 52.3082
R221 VDD1.t7 VDD1.n20 52.3082
R222 VDD1.n37 VDD1.n35 32.4212
R223 VDD1.n5 VDD1.n4 15.5966
R224 VDD1.n22 VDD1.n21 15.5966
R225 VDD1.n8 VDD1.n7 12.8005
R226 VDD1.n25 VDD1.n24 12.8005
R227 VDD1.n11 VDD1.n2 12.0247
R228 VDD1.n28 VDD1.n19 12.0247
R229 VDD1.n12 VDD1.n0 11.249
R230 VDD1.n29 VDD1.n17 11.249
R231 VDD1.n14 VDD1.n13 9.45567
R232 VDD1.n31 VDD1.n30 9.45567
R233 VDD1.n13 VDD1.n12 9.3005
R234 VDD1.n2 VDD1.n1 9.3005
R235 VDD1.n7 VDD1.n6 9.3005
R236 VDD1.n30 VDD1.n29 9.3005
R237 VDD1.n19 VDD1.n18 9.3005
R238 VDD1.n24 VDD1.n23 9.3005
R239 VDD1.n36 VDD1.t6 6.03709
R240 VDD1.n36 VDD1.t1 6.03709
R241 VDD1.n15 VDD1.t5 6.03709
R242 VDD1.n15 VDD1.t9 6.03709
R243 VDD1.n34 VDD1.t2 6.03709
R244 VDD1.n34 VDD1.t0 6.03709
R245 VDD1.n32 VDD1.t4 6.03709
R246 VDD1.n32 VDD1.t3 6.03709
R247 VDD1.n6 VDD1.n5 4.46457
R248 VDD1.n23 VDD1.n22 4.46457
R249 VDD1.n14 VDD1.n0 2.71565
R250 VDD1.n31 VDD1.n17 2.71565
R251 VDD1.n12 VDD1.n11 1.93989
R252 VDD1.n29 VDD1.n28 1.93989
R253 VDD1.n8 VDD1.n2 1.16414
R254 VDD1.n25 VDD1.n19 1.16414
R255 VDD1 VDD1.n37 0.698776
R256 VDD1.n7 VDD1.n4 0.388379
R257 VDD1.n24 VDD1.n21 0.388379
R258 VDD1 VDD1.n16 0.310845
R259 VDD1.n35 VDD1.n33 0.197309
R260 VDD1.n13 VDD1.n1 0.155672
R261 VDD1.n6 VDD1.n1 0.155672
R262 VDD1.n23 VDD1.n18 0.155672
R263 VDD1.n30 VDD1.n18 0.155672
R264 B.n445 B.n444 585
R265 B.n446 B.n445 585
R266 B.n159 B.n76 585
R267 B.n158 B.n157 585
R268 B.n156 B.n155 585
R269 B.n154 B.n153 585
R270 B.n152 B.n151 585
R271 B.n150 B.n149 585
R272 B.n148 B.n147 585
R273 B.n146 B.n145 585
R274 B.n144 B.n143 585
R275 B.n142 B.n141 585
R276 B.n140 B.n139 585
R277 B.n138 B.n137 585
R278 B.n136 B.n135 585
R279 B.n134 B.n133 585
R280 B.n132 B.n131 585
R281 B.n129 B.n128 585
R282 B.n127 B.n126 585
R283 B.n125 B.n124 585
R284 B.n123 B.n122 585
R285 B.n121 B.n120 585
R286 B.n119 B.n118 585
R287 B.n117 B.n116 585
R288 B.n115 B.n114 585
R289 B.n113 B.n112 585
R290 B.n111 B.n110 585
R291 B.n109 B.n108 585
R292 B.n107 B.n106 585
R293 B.n105 B.n104 585
R294 B.n103 B.n102 585
R295 B.n101 B.n100 585
R296 B.n99 B.n98 585
R297 B.n97 B.n96 585
R298 B.n95 B.n94 585
R299 B.n93 B.n92 585
R300 B.n91 B.n90 585
R301 B.n89 B.n88 585
R302 B.n87 B.n86 585
R303 B.n85 B.n84 585
R304 B.n83 B.n82 585
R305 B.n54 B.n53 585
R306 B.n443 B.n55 585
R307 B.n447 B.n55 585
R308 B.n442 B.n441 585
R309 B.n441 B.n51 585
R310 B.n440 B.n50 585
R311 B.n453 B.n50 585
R312 B.n439 B.n49 585
R313 B.n454 B.n49 585
R314 B.n438 B.n48 585
R315 B.n455 B.n48 585
R316 B.n437 B.n436 585
R317 B.n436 B.n44 585
R318 B.n435 B.n43 585
R319 B.n461 B.n43 585
R320 B.n434 B.n42 585
R321 B.n462 B.n42 585
R322 B.n433 B.n41 585
R323 B.n463 B.n41 585
R324 B.n432 B.n431 585
R325 B.n431 B.n37 585
R326 B.n430 B.n36 585
R327 B.n469 B.n36 585
R328 B.n429 B.n35 585
R329 B.n470 B.n35 585
R330 B.n428 B.n34 585
R331 B.n471 B.n34 585
R332 B.n427 B.n426 585
R333 B.n426 B.n30 585
R334 B.n425 B.n29 585
R335 B.n477 B.n29 585
R336 B.n424 B.n28 585
R337 B.n478 B.n28 585
R338 B.n423 B.n27 585
R339 B.n479 B.n27 585
R340 B.n422 B.n421 585
R341 B.n421 B.n23 585
R342 B.n420 B.n22 585
R343 B.n485 B.n22 585
R344 B.n419 B.n21 585
R345 B.n486 B.n21 585
R346 B.n418 B.n20 585
R347 B.n487 B.n20 585
R348 B.n417 B.n416 585
R349 B.n416 B.n19 585
R350 B.n415 B.n15 585
R351 B.n493 B.n15 585
R352 B.n414 B.n14 585
R353 B.n494 B.n14 585
R354 B.n413 B.n13 585
R355 B.n495 B.n13 585
R356 B.n412 B.n411 585
R357 B.n411 B.n12 585
R358 B.n410 B.n409 585
R359 B.n410 B.n8 585
R360 B.n408 B.n7 585
R361 B.n502 B.n7 585
R362 B.n407 B.n6 585
R363 B.n503 B.n6 585
R364 B.n406 B.n5 585
R365 B.n504 B.n5 585
R366 B.n405 B.n404 585
R367 B.n404 B.n4 585
R368 B.n403 B.n160 585
R369 B.n403 B.n402 585
R370 B.n392 B.n161 585
R371 B.n395 B.n161 585
R372 B.n394 B.n393 585
R373 B.n396 B.n394 585
R374 B.n391 B.n166 585
R375 B.n166 B.n165 585
R376 B.n390 B.n389 585
R377 B.n389 B.n388 585
R378 B.n168 B.n167 585
R379 B.n381 B.n168 585
R380 B.n380 B.n379 585
R381 B.n382 B.n380 585
R382 B.n378 B.n173 585
R383 B.n173 B.n172 585
R384 B.n377 B.n376 585
R385 B.n376 B.n375 585
R386 B.n175 B.n174 585
R387 B.n176 B.n175 585
R388 B.n368 B.n367 585
R389 B.n369 B.n368 585
R390 B.n366 B.n181 585
R391 B.n181 B.n180 585
R392 B.n365 B.n364 585
R393 B.n364 B.n363 585
R394 B.n183 B.n182 585
R395 B.n184 B.n183 585
R396 B.n356 B.n355 585
R397 B.n357 B.n356 585
R398 B.n354 B.n188 585
R399 B.n192 B.n188 585
R400 B.n353 B.n352 585
R401 B.n352 B.n351 585
R402 B.n190 B.n189 585
R403 B.n191 B.n190 585
R404 B.n344 B.n343 585
R405 B.n345 B.n344 585
R406 B.n342 B.n197 585
R407 B.n197 B.n196 585
R408 B.n341 B.n340 585
R409 B.n340 B.n339 585
R410 B.n199 B.n198 585
R411 B.n200 B.n199 585
R412 B.n332 B.n331 585
R413 B.n333 B.n332 585
R414 B.n330 B.n205 585
R415 B.n205 B.n204 585
R416 B.n329 B.n328 585
R417 B.n328 B.n327 585
R418 B.n207 B.n206 585
R419 B.n208 B.n207 585
R420 B.n320 B.n319 585
R421 B.n321 B.n320 585
R422 B.n211 B.n210 585
R423 B.n239 B.n237 585
R424 B.n240 B.n236 585
R425 B.n240 B.n212 585
R426 B.n243 B.n242 585
R427 B.n244 B.n235 585
R428 B.n246 B.n245 585
R429 B.n248 B.n234 585
R430 B.n251 B.n250 585
R431 B.n252 B.n233 585
R432 B.n254 B.n253 585
R433 B.n256 B.n232 585
R434 B.n259 B.n258 585
R435 B.n260 B.n231 585
R436 B.n262 B.n261 585
R437 B.n264 B.n230 585
R438 B.n267 B.n266 585
R439 B.n269 B.n227 585
R440 B.n271 B.n270 585
R441 B.n273 B.n226 585
R442 B.n276 B.n275 585
R443 B.n277 B.n225 585
R444 B.n279 B.n278 585
R445 B.n281 B.n224 585
R446 B.n284 B.n283 585
R447 B.n285 B.n221 585
R448 B.n288 B.n287 585
R449 B.n290 B.n220 585
R450 B.n293 B.n292 585
R451 B.n294 B.n219 585
R452 B.n296 B.n295 585
R453 B.n298 B.n218 585
R454 B.n301 B.n300 585
R455 B.n302 B.n217 585
R456 B.n304 B.n303 585
R457 B.n306 B.n216 585
R458 B.n309 B.n308 585
R459 B.n310 B.n215 585
R460 B.n312 B.n311 585
R461 B.n314 B.n214 585
R462 B.n317 B.n316 585
R463 B.n318 B.n213 585
R464 B.n323 B.n322 585
R465 B.n322 B.n321 585
R466 B.n324 B.n209 585
R467 B.n209 B.n208 585
R468 B.n326 B.n325 585
R469 B.n327 B.n326 585
R470 B.n203 B.n202 585
R471 B.n204 B.n203 585
R472 B.n335 B.n334 585
R473 B.n334 B.n333 585
R474 B.n336 B.n201 585
R475 B.n201 B.n200 585
R476 B.n338 B.n337 585
R477 B.n339 B.n338 585
R478 B.n195 B.n194 585
R479 B.n196 B.n195 585
R480 B.n347 B.n346 585
R481 B.n346 B.n345 585
R482 B.n348 B.n193 585
R483 B.n193 B.n191 585
R484 B.n350 B.n349 585
R485 B.n351 B.n350 585
R486 B.n187 B.n186 585
R487 B.n192 B.n187 585
R488 B.n359 B.n358 585
R489 B.n358 B.n357 585
R490 B.n360 B.n185 585
R491 B.n185 B.n184 585
R492 B.n362 B.n361 585
R493 B.n363 B.n362 585
R494 B.n179 B.n178 585
R495 B.n180 B.n179 585
R496 B.n371 B.n370 585
R497 B.n370 B.n369 585
R498 B.n372 B.n177 585
R499 B.n177 B.n176 585
R500 B.n374 B.n373 585
R501 B.n375 B.n374 585
R502 B.n171 B.n170 585
R503 B.n172 B.n171 585
R504 B.n384 B.n383 585
R505 B.n383 B.n382 585
R506 B.n385 B.n169 585
R507 B.n381 B.n169 585
R508 B.n387 B.n386 585
R509 B.n388 B.n387 585
R510 B.n164 B.n163 585
R511 B.n165 B.n164 585
R512 B.n398 B.n397 585
R513 B.n397 B.n396 585
R514 B.n399 B.n162 585
R515 B.n395 B.n162 585
R516 B.n401 B.n400 585
R517 B.n402 B.n401 585
R518 B.n3 B.n0 585
R519 B.n4 B.n3 585
R520 B.n501 B.n1 585
R521 B.n502 B.n501 585
R522 B.n500 B.n499 585
R523 B.n500 B.n8 585
R524 B.n498 B.n9 585
R525 B.n12 B.n9 585
R526 B.n497 B.n496 585
R527 B.n496 B.n495 585
R528 B.n11 B.n10 585
R529 B.n494 B.n11 585
R530 B.n492 B.n491 585
R531 B.n493 B.n492 585
R532 B.n490 B.n16 585
R533 B.n19 B.n16 585
R534 B.n489 B.n488 585
R535 B.n488 B.n487 585
R536 B.n18 B.n17 585
R537 B.n486 B.n18 585
R538 B.n484 B.n483 585
R539 B.n485 B.n484 585
R540 B.n482 B.n24 585
R541 B.n24 B.n23 585
R542 B.n481 B.n480 585
R543 B.n480 B.n479 585
R544 B.n26 B.n25 585
R545 B.n478 B.n26 585
R546 B.n476 B.n475 585
R547 B.n477 B.n476 585
R548 B.n474 B.n31 585
R549 B.n31 B.n30 585
R550 B.n473 B.n472 585
R551 B.n472 B.n471 585
R552 B.n33 B.n32 585
R553 B.n470 B.n33 585
R554 B.n468 B.n467 585
R555 B.n469 B.n468 585
R556 B.n466 B.n38 585
R557 B.n38 B.n37 585
R558 B.n465 B.n464 585
R559 B.n464 B.n463 585
R560 B.n40 B.n39 585
R561 B.n462 B.n40 585
R562 B.n460 B.n459 585
R563 B.n461 B.n460 585
R564 B.n458 B.n45 585
R565 B.n45 B.n44 585
R566 B.n457 B.n456 585
R567 B.n456 B.n455 585
R568 B.n47 B.n46 585
R569 B.n454 B.n47 585
R570 B.n452 B.n451 585
R571 B.n453 B.n452 585
R572 B.n450 B.n52 585
R573 B.n52 B.n51 585
R574 B.n449 B.n448 585
R575 B.n448 B.n447 585
R576 B.n505 B.n504 585
R577 B.n503 B.n2 585
R578 B.n448 B.n54 583.793
R579 B.n445 B.n55 583.793
R580 B.n320 B.n213 583.793
R581 B.n322 B.n211 583.793
R582 B.n79 B.t13 295.807
R583 B.n77 B.t9 295.807
R584 B.n222 B.t20 295.807
R585 B.n228 B.t16 295.807
R586 B.n446 B.n75 256.663
R587 B.n446 B.n74 256.663
R588 B.n446 B.n73 256.663
R589 B.n446 B.n72 256.663
R590 B.n446 B.n71 256.663
R591 B.n446 B.n70 256.663
R592 B.n446 B.n69 256.663
R593 B.n446 B.n68 256.663
R594 B.n446 B.n67 256.663
R595 B.n446 B.n66 256.663
R596 B.n446 B.n65 256.663
R597 B.n446 B.n64 256.663
R598 B.n446 B.n63 256.663
R599 B.n446 B.n62 256.663
R600 B.n446 B.n61 256.663
R601 B.n446 B.n60 256.663
R602 B.n446 B.n59 256.663
R603 B.n446 B.n58 256.663
R604 B.n446 B.n57 256.663
R605 B.n446 B.n56 256.663
R606 B.n238 B.n212 256.663
R607 B.n241 B.n212 256.663
R608 B.n247 B.n212 256.663
R609 B.n249 B.n212 256.663
R610 B.n255 B.n212 256.663
R611 B.n257 B.n212 256.663
R612 B.n263 B.n212 256.663
R613 B.n265 B.n212 256.663
R614 B.n272 B.n212 256.663
R615 B.n274 B.n212 256.663
R616 B.n280 B.n212 256.663
R617 B.n282 B.n212 256.663
R618 B.n289 B.n212 256.663
R619 B.n291 B.n212 256.663
R620 B.n297 B.n212 256.663
R621 B.n299 B.n212 256.663
R622 B.n305 B.n212 256.663
R623 B.n307 B.n212 256.663
R624 B.n313 B.n212 256.663
R625 B.n315 B.n212 256.663
R626 B.n507 B.n506 256.663
R627 B.n321 B.n212 181.298
R628 B.n447 B.n446 181.298
R629 B.n84 B.n83 163.367
R630 B.n88 B.n87 163.367
R631 B.n92 B.n91 163.367
R632 B.n96 B.n95 163.367
R633 B.n100 B.n99 163.367
R634 B.n104 B.n103 163.367
R635 B.n108 B.n107 163.367
R636 B.n112 B.n111 163.367
R637 B.n116 B.n115 163.367
R638 B.n120 B.n119 163.367
R639 B.n124 B.n123 163.367
R640 B.n128 B.n127 163.367
R641 B.n133 B.n132 163.367
R642 B.n137 B.n136 163.367
R643 B.n141 B.n140 163.367
R644 B.n145 B.n144 163.367
R645 B.n149 B.n148 163.367
R646 B.n153 B.n152 163.367
R647 B.n157 B.n156 163.367
R648 B.n445 B.n76 163.367
R649 B.n320 B.n207 163.367
R650 B.n328 B.n207 163.367
R651 B.n328 B.n205 163.367
R652 B.n332 B.n205 163.367
R653 B.n332 B.n199 163.367
R654 B.n340 B.n199 163.367
R655 B.n340 B.n197 163.367
R656 B.n344 B.n197 163.367
R657 B.n344 B.n190 163.367
R658 B.n352 B.n190 163.367
R659 B.n352 B.n188 163.367
R660 B.n356 B.n188 163.367
R661 B.n356 B.n183 163.367
R662 B.n364 B.n183 163.367
R663 B.n364 B.n181 163.367
R664 B.n368 B.n181 163.367
R665 B.n368 B.n175 163.367
R666 B.n376 B.n175 163.367
R667 B.n376 B.n173 163.367
R668 B.n380 B.n173 163.367
R669 B.n380 B.n168 163.367
R670 B.n389 B.n168 163.367
R671 B.n389 B.n166 163.367
R672 B.n394 B.n166 163.367
R673 B.n394 B.n161 163.367
R674 B.n403 B.n161 163.367
R675 B.n404 B.n403 163.367
R676 B.n404 B.n5 163.367
R677 B.n6 B.n5 163.367
R678 B.n7 B.n6 163.367
R679 B.n410 B.n7 163.367
R680 B.n411 B.n410 163.367
R681 B.n411 B.n13 163.367
R682 B.n14 B.n13 163.367
R683 B.n15 B.n14 163.367
R684 B.n416 B.n15 163.367
R685 B.n416 B.n20 163.367
R686 B.n21 B.n20 163.367
R687 B.n22 B.n21 163.367
R688 B.n421 B.n22 163.367
R689 B.n421 B.n27 163.367
R690 B.n28 B.n27 163.367
R691 B.n29 B.n28 163.367
R692 B.n426 B.n29 163.367
R693 B.n426 B.n34 163.367
R694 B.n35 B.n34 163.367
R695 B.n36 B.n35 163.367
R696 B.n431 B.n36 163.367
R697 B.n431 B.n41 163.367
R698 B.n42 B.n41 163.367
R699 B.n43 B.n42 163.367
R700 B.n436 B.n43 163.367
R701 B.n436 B.n48 163.367
R702 B.n49 B.n48 163.367
R703 B.n50 B.n49 163.367
R704 B.n441 B.n50 163.367
R705 B.n441 B.n55 163.367
R706 B.n240 B.n239 163.367
R707 B.n242 B.n240 163.367
R708 B.n246 B.n235 163.367
R709 B.n250 B.n248 163.367
R710 B.n254 B.n233 163.367
R711 B.n258 B.n256 163.367
R712 B.n262 B.n231 163.367
R713 B.n266 B.n264 163.367
R714 B.n271 B.n227 163.367
R715 B.n275 B.n273 163.367
R716 B.n279 B.n225 163.367
R717 B.n283 B.n281 163.367
R718 B.n288 B.n221 163.367
R719 B.n292 B.n290 163.367
R720 B.n296 B.n219 163.367
R721 B.n300 B.n298 163.367
R722 B.n304 B.n217 163.367
R723 B.n308 B.n306 163.367
R724 B.n312 B.n215 163.367
R725 B.n316 B.n314 163.367
R726 B.n322 B.n209 163.367
R727 B.n326 B.n209 163.367
R728 B.n326 B.n203 163.367
R729 B.n334 B.n203 163.367
R730 B.n334 B.n201 163.367
R731 B.n338 B.n201 163.367
R732 B.n338 B.n195 163.367
R733 B.n346 B.n195 163.367
R734 B.n346 B.n193 163.367
R735 B.n350 B.n193 163.367
R736 B.n350 B.n187 163.367
R737 B.n358 B.n187 163.367
R738 B.n358 B.n185 163.367
R739 B.n362 B.n185 163.367
R740 B.n362 B.n179 163.367
R741 B.n370 B.n179 163.367
R742 B.n370 B.n177 163.367
R743 B.n374 B.n177 163.367
R744 B.n374 B.n171 163.367
R745 B.n383 B.n171 163.367
R746 B.n383 B.n169 163.367
R747 B.n387 B.n169 163.367
R748 B.n387 B.n164 163.367
R749 B.n397 B.n164 163.367
R750 B.n397 B.n162 163.367
R751 B.n401 B.n162 163.367
R752 B.n401 B.n3 163.367
R753 B.n505 B.n3 163.367
R754 B.n501 B.n2 163.367
R755 B.n501 B.n500 163.367
R756 B.n500 B.n9 163.367
R757 B.n496 B.n9 163.367
R758 B.n496 B.n11 163.367
R759 B.n492 B.n11 163.367
R760 B.n492 B.n16 163.367
R761 B.n488 B.n16 163.367
R762 B.n488 B.n18 163.367
R763 B.n484 B.n18 163.367
R764 B.n484 B.n24 163.367
R765 B.n480 B.n24 163.367
R766 B.n480 B.n26 163.367
R767 B.n476 B.n26 163.367
R768 B.n476 B.n31 163.367
R769 B.n472 B.n31 163.367
R770 B.n472 B.n33 163.367
R771 B.n468 B.n33 163.367
R772 B.n468 B.n38 163.367
R773 B.n464 B.n38 163.367
R774 B.n464 B.n40 163.367
R775 B.n460 B.n40 163.367
R776 B.n460 B.n45 163.367
R777 B.n456 B.n45 163.367
R778 B.n456 B.n47 163.367
R779 B.n452 B.n47 163.367
R780 B.n452 B.n52 163.367
R781 B.n448 B.n52 163.367
R782 B.n77 B.t11 156.422
R783 B.n222 B.t22 156.422
R784 B.n79 B.t14 156.422
R785 B.n228 B.t19 156.422
R786 B.n78 B.t12 133.731
R787 B.n223 B.t21 133.731
R788 B.n80 B.t15 133.731
R789 B.n229 B.t18 133.731
R790 B.n321 B.n208 87.4347
R791 B.n327 B.n208 87.4347
R792 B.n327 B.n204 87.4347
R793 B.n333 B.n204 87.4347
R794 B.n339 B.n200 87.4347
R795 B.n339 B.n196 87.4347
R796 B.n345 B.n196 87.4347
R797 B.n345 B.n191 87.4347
R798 B.n351 B.n191 87.4347
R799 B.n351 B.n192 87.4347
R800 B.n357 B.n184 87.4347
R801 B.n363 B.n184 87.4347
R802 B.n369 B.n180 87.4347
R803 B.n369 B.n176 87.4347
R804 B.n375 B.n176 87.4347
R805 B.n382 B.n172 87.4347
R806 B.n382 B.n381 87.4347
R807 B.n388 B.n165 87.4347
R808 B.n396 B.n165 87.4347
R809 B.n396 B.n395 87.4347
R810 B.n402 B.n4 87.4347
R811 B.n504 B.n4 87.4347
R812 B.n504 B.n503 87.4347
R813 B.n503 B.n502 87.4347
R814 B.n502 B.n8 87.4347
R815 B.n495 B.n12 87.4347
R816 B.n495 B.n494 87.4347
R817 B.n494 B.n493 87.4347
R818 B.n487 B.n19 87.4347
R819 B.n487 B.n486 87.4347
R820 B.n485 B.n23 87.4347
R821 B.n479 B.n23 87.4347
R822 B.n479 B.n478 87.4347
R823 B.n477 B.n30 87.4347
R824 B.n471 B.n30 87.4347
R825 B.n470 B.n469 87.4347
R826 B.n469 B.n37 87.4347
R827 B.n463 B.n37 87.4347
R828 B.n463 B.n462 87.4347
R829 B.n462 B.n461 87.4347
R830 B.n461 B.n44 87.4347
R831 B.n455 B.n454 87.4347
R832 B.n454 B.n453 87.4347
R833 B.n453 B.n51 87.4347
R834 B.n447 B.n51 87.4347
R835 B.n363 B.t1 74.5768
R836 B.t2 B.n477 74.5768
R837 B.n402 B.t3 72.0052
R838 B.t4 B.n8 72.0052
R839 B.n56 B.n54 71.676
R840 B.n84 B.n57 71.676
R841 B.n88 B.n58 71.676
R842 B.n92 B.n59 71.676
R843 B.n96 B.n60 71.676
R844 B.n100 B.n61 71.676
R845 B.n104 B.n62 71.676
R846 B.n108 B.n63 71.676
R847 B.n112 B.n64 71.676
R848 B.n116 B.n65 71.676
R849 B.n120 B.n66 71.676
R850 B.n124 B.n67 71.676
R851 B.n128 B.n68 71.676
R852 B.n133 B.n69 71.676
R853 B.n137 B.n70 71.676
R854 B.n141 B.n71 71.676
R855 B.n145 B.n72 71.676
R856 B.n149 B.n73 71.676
R857 B.n153 B.n74 71.676
R858 B.n157 B.n75 71.676
R859 B.n76 B.n75 71.676
R860 B.n156 B.n74 71.676
R861 B.n152 B.n73 71.676
R862 B.n148 B.n72 71.676
R863 B.n144 B.n71 71.676
R864 B.n140 B.n70 71.676
R865 B.n136 B.n69 71.676
R866 B.n132 B.n68 71.676
R867 B.n127 B.n67 71.676
R868 B.n123 B.n66 71.676
R869 B.n119 B.n65 71.676
R870 B.n115 B.n64 71.676
R871 B.n111 B.n63 71.676
R872 B.n107 B.n62 71.676
R873 B.n103 B.n61 71.676
R874 B.n99 B.n60 71.676
R875 B.n95 B.n59 71.676
R876 B.n91 B.n58 71.676
R877 B.n87 B.n57 71.676
R878 B.n83 B.n56 71.676
R879 B.n238 B.n211 71.676
R880 B.n242 B.n241 71.676
R881 B.n247 B.n246 71.676
R882 B.n250 B.n249 71.676
R883 B.n255 B.n254 71.676
R884 B.n258 B.n257 71.676
R885 B.n263 B.n262 71.676
R886 B.n266 B.n265 71.676
R887 B.n272 B.n271 71.676
R888 B.n275 B.n274 71.676
R889 B.n280 B.n279 71.676
R890 B.n283 B.n282 71.676
R891 B.n289 B.n288 71.676
R892 B.n292 B.n291 71.676
R893 B.n297 B.n296 71.676
R894 B.n300 B.n299 71.676
R895 B.n305 B.n304 71.676
R896 B.n308 B.n307 71.676
R897 B.n313 B.n312 71.676
R898 B.n316 B.n315 71.676
R899 B.n239 B.n238 71.676
R900 B.n241 B.n235 71.676
R901 B.n248 B.n247 71.676
R902 B.n249 B.n233 71.676
R903 B.n256 B.n255 71.676
R904 B.n257 B.n231 71.676
R905 B.n264 B.n263 71.676
R906 B.n265 B.n227 71.676
R907 B.n273 B.n272 71.676
R908 B.n274 B.n225 71.676
R909 B.n281 B.n280 71.676
R910 B.n282 B.n221 71.676
R911 B.n290 B.n289 71.676
R912 B.n291 B.n219 71.676
R913 B.n298 B.n297 71.676
R914 B.n299 B.n217 71.676
R915 B.n306 B.n305 71.676
R916 B.n307 B.n215 71.676
R917 B.n314 B.n313 71.676
R918 B.n315 B.n213 71.676
R919 B.n506 B.n505 71.676
R920 B.n506 B.n2 71.676
R921 B.n333 B.t17 66.862
R922 B.n455 B.t10 66.862
R923 B.n381 B.t0 64.2904
R924 B.n19 B.t8 64.2904
R925 B.t5 B.n172 61.7188
R926 B.n486 B.t6 61.7188
R927 B.n81 B.n80 59.5399
R928 B.n130 B.n78 59.5399
R929 B.n286 B.n223 59.5399
R930 B.n268 B.n229 59.5399
R931 B.n357 B.t7 51.4324
R932 B.n471 B.t23 51.4324
R933 B.n323 B.n210 37.9322
R934 B.n319 B.n318 37.9322
R935 B.n444 B.n443 37.9322
R936 B.n449 B.n53 37.9322
R937 B.n192 B.t7 36.0028
R938 B.t23 B.n470 36.0028
R939 B.n375 B.t5 25.7165
R940 B.t6 B.n485 25.7165
R941 B.n388 B.t0 23.1449
R942 B.n493 B.t8 23.1449
R943 B.n80 B.n79 22.6914
R944 B.n78 B.n77 22.6914
R945 B.n223 B.n222 22.6914
R946 B.n229 B.n228 22.6914
R947 B.t17 B.n200 20.5733
R948 B.t10 B.n44 20.5733
R949 B B.n507 18.0485
R950 B.n395 B.t3 15.4301
R951 B.n12 B.t4 15.4301
R952 B.t1 B.n180 12.8585
R953 B.n478 B.t2 12.8585
R954 B.n324 B.n323 10.6151
R955 B.n325 B.n324 10.6151
R956 B.n325 B.n202 10.6151
R957 B.n335 B.n202 10.6151
R958 B.n336 B.n335 10.6151
R959 B.n337 B.n336 10.6151
R960 B.n337 B.n194 10.6151
R961 B.n347 B.n194 10.6151
R962 B.n348 B.n347 10.6151
R963 B.n349 B.n348 10.6151
R964 B.n349 B.n186 10.6151
R965 B.n359 B.n186 10.6151
R966 B.n360 B.n359 10.6151
R967 B.n361 B.n360 10.6151
R968 B.n361 B.n178 10.6151
R969 B.n371 B.n178 10.6151
R970 B.n372 B.n371 10.6151
R971 B.n373 B.n372 10.6151
R972 B.n373 B.n170 10.6151
R973 B.n384 B.n170 10.6151
R974 B.n385 B.n384 10.6151
R975 B.n386 B.n385 10.6151
R976 B.n386 B.n163 10.6151
R977 B.n398 B.n163 10.6151
R978 B.n399 B.n398 10.6151
R979 B.n400 B.n399 10.6151
R980 B.n400 B.n0 10.6151
R981 B.n237 B.n210 10.6151
R982 B.n237 B.n236 10.6151
R983 B.n243 B.n236 10.6151
R984 B.n244 B.n243 10.6151
R985 B.n245 B.n244 10.6151
R986 B.n245 B.n234 10.6151
R987 B.n251 B.n234 10.6151
R988 B.n252 B.n251 10.6151
R989 B.n253 B.n252 10.6151
R990 B.n253 B.n232 10.6151
R991 B.n259 B.n232 10.6151
R992 B.n260 B.n259 10.6151
R993 B.n261 B.n260 10.6151
R994 B.n261 B.n230 10.6151
R995 B.n267 B.n230 10.6151
R996 B.n270 B.n269 10.6151
R997 B.n270 B.n226 10.6151
R998 B.n276 B.n226 10.6151
R999 B.n277 B.n276 10.6151
R1000 B.n278 B.n277 10.6151
R1001 B.n278 B.n224 10.6151
R1002 B.n284 B.n224 10.6151
R1003 B.n285 B.n284 10.6151
R1004 B.n287 B.n220 10.6151
R1005 B.n293 B.n220 10.6151
R1006 B.n294 B.n293 10.6151
R1007 B.n295 B.n294 10.6151
R1008 B.n295 B.n218 10.6151
R1009 B.n301 B.n218 10.6151
R1010 B.n302 B.n301 10.6151
R1011 B.n303 B.n302 10.6151
R1012 B.n303 B.n216 10.6151
R1013 B.n309 B.n216 10.6151
R1014 B.n310 B.n309 10.6151
R1015 B.n311 B.n310 10.6151
R1016 B.n311 B.n214 10.6151
R1017 B.n317 B.n214 10.6151
R1018 B.n318 B.n317 10.6151
R1019 B.n319 B.n206 10.6151
R1020 B.n329 B.n206 10.6151
R1021 B.n330 B.n329 10.6151
R1022 B.n331 B.n330 10.6151
R1023 B.n331 B.n198 10.6151
R1024 B.n341 B.n198 10.6151
R1025 B.n342 B.n341 10.6151
R1026 B.n343 B.n342 10.6151
R1027 B.n343 B.n189 10.6151
R1028 B.n353 B.n189 10.6151
R1029 B.n354 B.n353 10.6151
R1030 B.n355 B.n354 10.6151
R1031 B.n355 B.n182 10.6151
R1032 B.n365 B.n182 10.6151
R1033 B.n366 B.n365 10.6151
R1034 B.n367 B.n366 10.6151
R1035 B.n367 B.n174 10.6151
R1036 B.n377 B.n174 10.6151
R1037 B.n378 B.n377 10.6151
R1038 B.n379 B.n378 10.6151
R1039 B.n379 B.n167 10.6151
R1040 B.n390 B.n167 10.6151
R1041 B.n391 B.n390 10.6151
R1042 B.n393 B.n391 10.6151
R1043 B.n393 B.n392 10.6151
R1044 B.n392 B.n160 10.6151
R1045 B.n405 B.n160 10.6151
R1046 B.n406 B.n405 10.6151
R1047 B.n407 B.n406 10.6151
R1048 B.n408 B.n407 10.6151
R1049 B.n409 B.n408 10.6151
R1050 B.n412 B.n409 10.6151
R1051 B.n413 B.n412 10.6151
R1052 B.n414 B.n413 10.6151
R1053 B.n415 B.n414 10.6151
R1054 B.n417 B.n415 10.6151
R1055 B.n418 B.n417 10.6151
R1056 B.n419 B.n418 10.6151
R1057 B.n420 B.n419 10.6151
R1058 B.n422 B.n420 10.6151
R1059 B.n423 B.n422 10.6151
R1060 B.n424 B.n423 10.6151
R1061 B.n425 B.n424 10.6151
R1062 B.n427 B.n425 10.6151
R1063 B.n428 B.n427 10.6151
R1064 B.n429 B.n428 10.6151
R1065 B.n430 B.n429 10.6151
R1066 B.n432 B.n430 10.6151
R1067 B.n433 B.n432 10.6151
R1068 B.n434 B.n433 10.6151
R1069 B.n435 B.n434 10.6151
R1070 B.n437 B.n435 10.6151
R1071 B.n438 B.n437 10.6151
R1072 B.n439 B.n438 10.6151
R1073 B.n440 B.n439 10.6151
R1074 B.n442 B.n440 10.6151
R1075 B.n443 B.n442 10.6151
R1076 B.n499 B.n1 10.6151
R1077 B.n499 B.n498 10.6151
R1078 B.n498 B.n497 10.6151
R1079 B.n497 B.n10 10.6151
R1080 B.n491 B.n10 10.6151
R1081 B.n491 B.n490 10.6151
R1082 B.n490 B.n489 10.6151
R1083 B.n489 B.n17 10.6151
R1084 B.n483 B.n17 10.6151
R1085 B.n483 B.n482 10.6151
R1086 B.n482 B.n481 10.6151
R1087 B.n481 B.n25 10.6151
R1088 B.n475 B.n25 10.6151
R1089 B.n475 B.n474 10.6151
R1090 B.n474 B.n473 10.6151
R1091 B.n473 B.n32 10.6151
R1092 B.n467 B.n32 10.6151
R1093 B.n467 B.n466 10.6151
R1094 B.n466 B.n465 10.6151
R1095 B.n465 B.n39 10.6151
R1096 B.n459 B.n39 10.6151
R1097 B.n459 B.n458 10.6151
R1098 B.n458 B.n457 10.6151
R1099 B.n457 B.n46 10.6151
R1100 B.n451 B.n46 10.6151
R1101 B.n451 B.n450 10.6151
R1102 B.n450 B.n449 10.6151
R1103 B.n82 B.n53 10.6151
R1104 B.n85 B.n82 10.6151
R1105 B.n86 B.n85 10.6151
R1106 B.n89 B.n86 10.6151
R1107 B.n90 B.n89 10.6151
R1108 B.n93 B.n90 10.6151
R1109 B.n94 B.n93 10.6151
R1110 B.n97 B.n94 10.6151
R1111 B.n98 B.n97 10.6151
R1112 B.n101 B.n98 10.6151
R1113 B.n102 B.n101 10.6151
R1114 B.n105 B.n102 10.6151
R1115 B.n106 B.n105 10.6151
R1116 B.n109 B.n106 10.6151
R1117 B.n110 B.n109 10.6151
R1118 B.n114 B.n113 10.6151
R1119 B.n117 B.n114 10.6151
R1120 B.n118 B.n117 10.6151
R1121 B.n121 B.n118 10.6151
R1122 B.n122 B.n121 10.6151
R1123 B.n125 B.n122 10.6151
R1124 B.n126 B.n125 10.6151
R1125 B.n129 B.n126 10.6151
R1126 B.n134 B.n131 10.6151
R1127 B.n135 B.n134 10.6151
R1128 B.n138 B.n135 10.6151
R1129 B.n139 B.n138 10.6151
R1130 B.n142 B.n139 10.6151
R1131 B.n143 B.n142 10.6151
R1132 B.n146 B.n143 10.6151
R1133 B.n147 B.n146 10.6151
R1134 B.n150 B.n147 10.6151
R1135 B.n151 B.n150 10.6151
R1136 B.n154 B.n151 10.6151
R1137 B.n155 B.n154 10.6151
R1138 B.n158 B.n155 10.6151
R1139 B.n159 B.n158 10.6151
R1140 B.n444 B.n159 10.6151
R1141 B.n507 B.n0 8.11757
R1142 B.n507 B.n1 8.11757
R1143 B.n269 B.n268 6.5566
R1144 B.n286 B.n285 6.5566
R1145 B.n113 B.n81 6.5566
R1146 B.n130 B.n129 6.5566
R1147 B.n268 B.n267 4.05904
R1148 B.n287 B.n286 4.05904
R1149 B.n110 B.n81 4.05904
R1150 B.n131 B.n130 4.05904
R1151 VN.n5 VN.t6 165.869
R1152 VN.n23 VN.t7 165.869
R1153 VN.n17 VN.n16 161.3
R1154 VN.n35 VN.n34 161.3
R1155 VN.n33 VN.n18 161.3
R1156 VN.n32 VN.n31 161.3
R1157 VN.n30 VN.n29 161.3
R1158 VN.n28 VN.n20 161.3
R1159 VN.n26 VN.n25 161.3
R1160 VN.n24 VN.n21 161.3
R1161 VN.n15 VN.n0 161.3
R1162 VN.n14 VN.n13 161.3
R1163 VN.n12 VN.n11 161.3
R1164 VN.n10 VN.n2 161.3
R1165 VN.n8 VN.n7 161.3
R1166 VN.n6 VN.n3 161.3
R1167 VN.n16 VN.t0 140.87
R1168 VN.n34 VN.t4 140.87
R1169 VN.n4 VN.t3 94.1053
R1170 VN.n9 VN.t2 94.1053
R1171 VN.n1 VN.t1 94.1053
R1172 VN.n22 VN.t9 94.1053
R1173 VN.n27 VN.t5 94.1053
R1174 VN.n19 VN.t8 94.1053
R1175 VN.n8 VN.n3 56.5617
R1176 VN.n11 VN.n10 56.5617
R1177 VN.n26 VN.n21 56.5617
R1178 VN.n29 VN.n28 56.5617
R1179 VN.n24 VN.n23 42.2591
R1180 VN.n6 VN.n5 42.2591
R1181 VN.n15 VN.n14 40.0926
R1182 VN.n33 VN.n32 40.0926
R1183 VN VN.n35 37.3774
R1184 VN.n5 VN.n4 32.8395
R1185 VN.n23 VN.n22 32.8395
R1186 VN.n16 VN.n15 24.8308
R1187 VN.n34 VN.n33 24.8308
R1188 VN.n4 VN.n3 20.6576
R1189 VN.n11 VN.n1 20.6576
R1190 VN.n22 VN.n21 20.6576
R1191 VN.n29 VN.n19 20.6576
R1192 VN.n9 VN.n8 12.2964
R1193 VN.n10 VN.n9 12.2964
R1194 VN.n28 VN.n27 12.2964
R1195 VN.n27 VN.n26 12.2964
R1196 VN.n14 VN.n1 3.93519
R1197 VN.n32 VN.n19 3.93519
R1198 VN.n35 VN.n18 0.189894
R1199 VN.n31 VN.n18 0.189894
R1200 VN.n31 VN.n30 0.189894
R1201 VN.n30 VN.n20 0.189894
R1202 VN.n25 VN.n20 0.189894
R1203 VN.n25 VN.n24 0.189894
R1204 VN.n7 VN.n6 0.189894
R1205 VN.n7 VN.n2 0.189894
R1206 VN.n12 VN.n2 0.189894
R1207 VN.n13 VN.n12 0.189894
R1208 VN.n13 VN.n0 0.189894
R1209 VN.n17 VN.n0 0.189894
R1210 VN VN.n17 0.0516364
R1211 VDD2.n29 VDD2.n19 289.615
R1212 VDD2.n10 VDD2.n0 289.615
R1213 VDD2.n30 VDD2.n29 185
R1214 VDD2.n28 VDD2.n27 185
R1215 VDD2.n23 VDD2.n22 185
R1216 VDD2.n4 VDD2.n3 185
R1217 VDD2.n9 VDD2.n8 185
R1218 VDD2.n11 VDD2.n10 185
R1219 VDD2.n24 VDD2.t5 148.606
R1220 VDD2.n5 VDD2.t3 148.606
R1221 VDD2.n29 VDD2.n28 104.615
R1222 VDD2.n28 VDD2.n22 104.615
R1223 VDD2.n9 VDD2.n3 104.615
R1224 VDD2.n10 VDD2.n9 104.615
R1225 VDD2.n18 VDD2.n17 81.5532
R1226 VDD2 VDD2.n37 81.5504
R1227 VDD2.n36 VDD2.n35 80.8522
R1228 VDD2.n16 VDD2.n15 80.8521
R1229 VDD2.n16 VDD2.n14 52.9758
R1230 VDD2.t5 VDD2.n22 52.3082
R1231 VDD2.t3 VDD2.n3 52.3082
R1232 VDD2.n34 VDD2.n33 51.9672
R1233 VDD2.n34 VDD2.n18 31.3338
R1234 VDD2.n24 VDD2.n23 15.5966
R1235 VDD2.n5 VDD2.n4 15.5966
R1236 VDD2.n27 VDD2.n26 12.8005
R1237 VDD2.n8 VDD2.n7 12.8005
R1238 VDD2.n30 VDD2.n21 12.0247
R1239 VDD2.n11 VDD2.n2 12.0247
R1240 VDD2.n31 VDD2.n19 11.249
R1241 VDD2.n12 VDD2.n0 11.249
R1242 VDD2.n33 VDD2.n32 9.45567
R1243 VDD2.n14 VDD2.n13 9.45567
R1244 VDD2.n32 VDD2.n31 9.3005
R1245 VDD2.n21 VDD2.n20 9.3005
R1246 VDD2.n26 VDD2.n25 9.3005
R1247 VDD2.n13 VDD2.n12 9.3005
R1248 VDD2.n2 VDD2.n1 9.3005
R1249 VDD2.n7 VDD2.n6 9.3005
R1250 VDD2.n37 VDD2.t0 6.03709
R1251 VDD2.n37 VDD2.t2 6.03709
R1252 VDD2.n35 VDD2.t1 6.03709
R1253 VDD2.n35 VDD2.t4 6.03709
R1254 VDD2.n17 VDD2.t8 6.03709
R1255 VDD2.n17 VDD2.t9 6.03709
R1256 VDD2.n15 VDD2.t6 6.03709
R1257 VDD2.n15 VDD2.t7 6.03709
R1258 VDD2.n25 VDD2.n24 4.46457
R1259 VDD2.n6 VDD2.n5 4.46457
R1260 VDD2.n33 VDD2.n19 2.71565
R1261 VDD2.n14 VDD2.n0 2.71565
R1262 VDD2.n31 VDD2.n30 1.93989
R1263 VDD2.n12 VDD2.n11 1.93989
R1264 VDD2.n27 VDD2.n21 1.16414
R1265 VDD2.n8 VDD2.n2 1.16414
R1266 VDD2.n36 VDD2.n34 1.00912
R1267 VDD2.n26 VDD2.n23 0.388379
R1268 VDD2.n7 VDD2.n4 0.388379
R1269 VDD2 VDD2.n36 0.310845
R1270 VDD2.n18 VDD2.n16 0.197309
R1271 VDD2.n32 VDD2.n20 0.155672
R1272 VDD2.n25 VDD2.n20 0.155672
R1273 VDD2.n6 VDD2.n1 0.155672
R1274 VDD2.n13 VDD2.n1 0.155672
C0 VDD2 VP 0.363707f
C1 VDD2 VTAIL 5.58912f
C2 VDD2 VN 2.3314f
C3 VDD1 VP 2.53841f
C4 VDD1 VTAIL 5.54899f
C5 VDD1 VN 0.154412f
C6 VDD1 VDD2 1.05686f
C7 VP VTAIL 2.69632f
C8 VP VN 4.18902f
C9 VN VTAIL 2.68209f
C10 VDD2 B 3.559369f
C11 VDD1 B 3.505346f
C12 VTAIL B 3.240263f
C13 VN B 8.995939f
C14 VP B 7.433147f
C15 VDD2.n0 B 0.033793f
C16 VDD2.n1 B 0.024042f
C17 VDD2.n2 B 0.012919f
C18 VDD2.n3 B 0.022902f
C19 VDD2.n4 B 0.017806f
C20 VDD2.t3 B 0.051873f
C21 VDD2.n5 B 0.090143f
C22 VDD2.n6 B 0.266598f
C23 VDD2.n7 B 0.012919f
C24 VDD2.n8 B 0.013679f
C25 VDD2.n9 B 0.030536f
C26 VDD2.n10 B 0.066105f
C27 VDD2.n11 B 0.013679f
C28 VDD2.n12 B 0.012919f
C29 VDD2.n13 B 0.060826f
C30 VDD2.n14 B 0.056133f
C31 VDD2.t6 B 0.062315f
C32 VDD2.t7 B 0.062315f
C33 VDD2.n15 B 0.470427f
C34 VDD2.n16 B 0.404915f
C35 VDD2.t8 B 0.062315f
C36 VDD2.t9 B 0.062315f
C37 VDD2.n17 B 0.473235f
C38 VDD2.n18 B 1.39519f
C39 VDD2.n19 B 0.033793f
C40 VDD2.n20 B 0.024042f
C41 VDD2.n21 B 0.012919f
C42 VDD2.n22 B 0.022902f
C43 VDD2.n23 B 0.017806f
C44 VDD2.t5 B 0.051873f
C45 VDD2.n24 B 0.090143f
C46 VDD2.n25 B 0.266598f
C47 VDD2.n26 B 0.012919f
C48 VDD2.n27 B 0.013679f
C49 VDD2.n28 B 0.030536f
C50 VDD2.n29 B 0.066105f
C51 VDD2.n30 B 0.013679f
C52 VDD2.n31 B 0.012919f
C53 VDD2.n32 B 0.060826f
C54 VDD2.n33 B 0.053706f
C55 VDD2.n34 B 1.45594f
C56 VDD2.t1 B 0.062315f
C57 VDD2.t4 B 0.062315f
C58 VDD2.n35 B 0.470429f
C59 VDD2.n36 B 0.285863f
C60 VDD2.t0 B 0.062315f
C61 VDD2.t2 B 0.062315f
C62 VDD2.n37 B 0.473215f
C63 VN.n0 B 0.042444f
C64 VN.t1 B 0.294417f
C65 VN.n1 B 0.148097f
C66 VN.n2 B 0.042444f
C67 VN.t2 B 0.294417f
C68 VN.n3 B 0.0455f
C69 VN.t6 B 0.378925f
C70 VN.t3 B 0.294417f
C71 VN.n4 B 0.197807f
C72 VN.n5 B 0.185843f
C73 VN.n6 B 0.182438f
C74 VN.n7 B 0.042444f
C75 VN.n8 B 0.052252f
C76 VN.n9 B 0.148097f
C77 VN.n10 B 0.052252f
C78 VN.n11 B 0.0455f
C79 VN.n12 B 0.042444f
C80 VN.n13 B 0.042444f
C81 VN.n14 B 0.051477f
C82 VN.n15 B 0.022398f
C83 VN.t0 B 0.348705f
C84 VN.n16 B 0.190954f
C85 VN.n17 B 0.032892f
C86 VN.n18 B 0.042444f
C87 VN.t8 B 0.294417f
C88 VN.n19 B 0.148097f
C89 VN.n20 B 0.042444f
C90 VN.t5 B 0.294417f
C91 VN.n21 B 0.0455f
C92 VN.t7 B 0.378925f
C93 VN.t9 B 0.294417f
C94 VN.n22 B 0.197807f
C95 VN.n23 B 0.185843f
C96 VN.n24 B 0.182438f
C97 VN.n25 B 0.042444f
C98 VN.n26 B 0.052252f
C99 VN.n27 B 0.148097f
C100 VN.n28 B 0.052252f
C101 VN.n29 B 0.0455f
C102 VN.n30 B 0.042444f
C103 VN.n31 B 0.042444f
C104 VN.n32 B 0.051477f
C105 VN.n33 B 0.022398f
C106 VN.t4 B 0.348705f
C107 VN.n34 B 0.190954f
C108 VN.n35 B 1.43187f
C109 VDD1.n0 B 0.03384f
C110 VDD1.n1 B 0.024076f
C111 VDD1.n2 B 0.012937f
C112 VDD1.n3 B 0.022934f
C113 VDD1.n4 B 0.017831f
C114 VDD1.t8 B 0.051946f
C115 VDD1.n5 B 0.090269f
C116 VDD1.n6 B 0.266972f
C117 VDD1.n7 B 0.012937f
C118 VDD1.n8 B 0.013698f
C119 VDD1.n9 B 0.030579f
C120 VDD1.n10 B 0.066198f
C121 VDD1.n11 B 0.013698f
C122 VDD1.n12 B 0.012937f
C123 VDD1.n13 B 0.060912f
C124 VDD1.n14 B 0.056211f
C125 VDD1.t5 B 0.062403f
C126 VDD1.t9 B 0.062403f
C127 VDD1.n15 B 0.471089f
C128 VDD1.n16 B 0.411453f
C129 VDD1.n17 B 0.03384f
C130 VDD1.n18 B 0.024076f
C131 VDD1.n19 B 0.012937f
C132 VDD1.n20 B 0.022934f
C133 VDD1.n21 B 0.017831f
C134 VDD1.t7 B 0.051946f
C135 VDD1.n22 B 0.090269f
C136 VDD1.n23 B 0.266972f
C137 VDD1.n24 B 0.012937f
C138 VDD1.n25 B 0.013698f
C139 VDD1.n26 B 0.030579f
C140 VDD1.n27 B 0.066198f
C141 VDD1.n28 B 0.013698f
C142 VDD1.n29 B 0.012937f
C143 VDD1.n30 B 0.060912f
C144 VDD1.n31 B 0.056211f
C145 VDD1.t4 B 0.062403f
C146 VDD1.t3 B 0.062403f
C147 VDD1.n32 B 0.471086f
C148 VDD1.n33 B 0.405483f
C149 VDD1.t2 B 0.062403f
C150 VDD1.t0 B 0.062403f
C151 VDD1.n34 B 0.473898f
C152 VDD1.n35 B 1.47023f
C153 VDD1.t6 B 0.062403f
C154 VDD1.t1 B 0.062403f
C155 VDD1.n36 B 0.471086f
C156 VDD1.n37 B 1.67226f
C157 VTAIL.t4 B 0.077091f
C158 VTAIL.t8 B 0.077091f
C159 VTAIL.n0 B 0.524384f
C160 VTAIL.n1 B 0.41584f
C161 VTAIL.n2 B 0.041806f
C162 VTAIL.n3 B 0.029743f
C163 VTAIL.n4 B 0.015982f
C164 VTAIL.n5 B 0.028332f
C165 VTAIL.n6 B 0.022028f
C166 VTAIL.t18 B 0.064173f
C167 VTAIL.n7 B 0.111517f
C168 VTAIL.n8 B 0.329814f
C169 VTAIL.n9 B 0.015982f
C170 VTAIL.n10 B 0.016922f
C171 VTAIL.n11 B 0.037776f
C172 VTAIL.n12 B 0.08178f
C173 VTAIL.n13 B 0.016922f
C174 VTAIL.n14 B 0.015982f
C175 VTAIL.n15 B 0.075249f
C176 VTAIL.n16 B 0.045951f
C177 VTAIL.n17 B 0.219101f
C178 VTAIL.t11 B 0.077091f
C179 VTAIL.t16 B 0.077091f
C180 VTAIL.n18 B 0.524384f
C181 VTAIL.n19 B 0.437734f
C182 VTAIL.t9 B 0.077091f
C183 VTAIL.t17 B 0.077091f
C184 VTAIL.n20 B 0.524384f
C185 VTAIL.n21 B 1.2094f
C186 VTAIL.t7 B 0.077091f
C187 VTAIL.t1 B 0.077091f
C188 VTAIL.n22 B 0.524387f
C189 VTAIL.n23 B 1.2094f
C190 VTAIL.t5 B 0.077091f
C191 VTAIL.t0 B 0.077091f
C192 VTAIL.n24 B 0.524387f
C193 VTAIL.n25 B 0.43773f
C194 VTAIL.n26 B 0.041806f
C195 VTAIL.n27 B 0.029743f
C196 VTAIL.n28 B 0.015982f
C197 VTAIL.n29 B 0.028332f
C198 VTAIL.n30 B 0.022028f
C199 VTAIL.t3 B 0.064173f
C200 VTAIL.n31 B 0.111517f
C201 VTAIL.n32 B 0.329814f
C202 VTAIL.n33 B 0.015982f
C203 VTAIL.n34 B 0.016922f
C204 VTAIL.n35 B 0.037776f
C205 VTAIL.n36 B 0.08178f
C206 VTAIL.n37 B 0.016922f
C207 VTAIL.n38 B 0.015982f
C208 VTAIL.n39 B 0.075249f
C209 VTAIL.n40 B 0.045951f
C210 VTAIL.n41 B 0.219101f
C211 VTAIL.t12 B 0.077091f
C212 VTAIL.t13 B 0.077091f
C213 VTAIL.n42 B 0.524387f
C214 VTAIL.n43 B 0.434426f
C215 VTAIL.t14 B 0.077091f
C216 VTAIL.t15 B 0.077091f
C217 VTAIL.n44 B 0.524387f
C218 VTAIL.n45 B 0.43773f
C219 VTAIL.n46 B 0.041806f
C220 VTAIL.n47 B 0.029743f
C221 VTAIL.n48 B 0.015982f
C222 VTAIL.n49 B 0.028332f
C223 VTAIL.n50 B 0.022028f
C224 VTAIL.t10 B 0.064173f
C225 VTAIL.n51 B 0.111517f
C226 VTAIL.n52 B 0.329814f
C227 VTAIL.n53 B 0.015982f
C228 VTAIL.n54 B 0.016922f
C229 VTAIL.n55 B 0.037776f
C230 VTAIL.n56 B 0.08178f
C231 VTAIL.n57 B 0.016922f
C232 VTAIL.n58 B 0.015982f
C233 VTAIL.n59 B 0.075249f
C234 VTAIL.n60 B 0.045951f
C235 VTAIL.n61 B 0.897411f
C236 VTAIL.n62 B 0.041806f
C237 VTAIL.n63 B 0.029743f
C238 VTAIL.n64 B 0.015982f
C239 VTAIL.n65 B 0.028332f
C240 VTAIL.n66 B 0.022028f
C241 VTAIL.t19 B 0.064173f
C242 VTAIL.n67 B 0.111517f
C243 VTAIL.n68 B 0.329814f
C244 VTAIL.n69 B 0.015982f
C245 VTAIL.n70 B 0.016922f
C246 VTAIL.n71 B 0.037776f
C247 VTAIL.n72 B 0.08178f
C248 VTAIL.n73 B 0.016922f
C249 VTAIL.n74 B 0.015982f
C250 VTAIL.n75 B 0.075249f
C251 VTAIL.n76 B 0.045951f
C252 VTAIL.n77 B 0.897411f
C253 VTAIL.t6 B 0.077091f
C254 VTAIL.t2 B 0.077091f
C255 VTAIL.n78 B 0.524384f
C256 VTAIL.n79 B 0.35966f
C257 VP.n0 B 0.043649f
C258 VP.t7 B 0.302781f
C259 VP.n1 B 0.152304f
C260 VP.n2 B 0.043649f
C261 VP.t6 B 0.302781f
C262 VP.n3 B 0.046792f
C263 VP.n4 B 0.043649f
C264 VP.n5 B 0.043649f
C265 VP.t8 B 0.358611f
C266 VP.t3 B 0.302781f
C267 VP.n6 B 0.152304f
C268 VP.n7 B 0.043649f
C269 VP.t0 B 0.302781f
C270 VP.n8 B 0.046792f
C271 VP.t4 B 0.302781f
C272 VP.n9 B 0.203426f
C273 VP.t1 B 0.38969f
C274 VP.n10 B 0.191122f
C275 VP.n11 B 0.187621f
C276 VP.n12 B 0.043649f
C277 VP.n13 B 0.053736f
C278 VP.n14 B 0.152304f
C279 VP.n15 B 0.053736f
C280 VP.n16 B 0.046792f
C281 VP.n17 B 0.043649f
C282 VP.n18 B 0.043649f
C283 VP.n19 B 0.052939f
C284 VP.n20 B 0.023035f
C285 VP.n21 B 0.196379f
C286 VP.n22 B 1.44366f
C287 VP.n23 B 1.48619f
C288 VP.t2 B 0.358611f
C289 VP.n24 B 0.196379f
C290 VP.n25 B 0.023035f
C291 VP.t5 B 0.302781f
C292 VP.n26 B 0.152304f
C293 VP.n27 B 0.052939f
C294 VP.n28 B 0.043649f
C295 VP.n29 B 0.043649f
C296 VP.n30 B 0.043649f
C297 VP.n31 B 0.053736f
C298 VP.n32 B 0.152304f
C299 VP.n33 B 0.053736f
C300 VP.n34 B 0.046792f
C301 VP.n35 B 0.043649f
C302 VP.n36 B 0.043649f
C303 VP.n37 B 0.052939f
C304 VP.n38 B 0.023035f
C305 VP.t9 B 0.358611f
C306 VP.n39 B 0.196379f
C307 VP.n40 B 0.033827f
.ends

