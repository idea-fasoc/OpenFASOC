* NGSPICE file created from diff_pair_sample_1585.ext - technology: sky130A

.subckt diff_pair_sample_1585 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=1.59
X1 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=1.59
X2 VDD1.t7 VP.t0 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X3 VDD2.t7 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=1.59
X4 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=1.59
X5 VTAIL.t8 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X6 VTAIL.t5 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=1.59
X7 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X8 VDD1.t5 VP.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=1.59
X9 VTAIL.t11 VP.t3 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=1.59
X10 VDD2.t4 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X11 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=1.59
X12 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X13 VTAIL.t3 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X14 VDD1.t3 VP.t4 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=1.59
X15 VTAIL.t14 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X16 VDD1.t1 VP.t6 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=1.59
X17 VTAIL.t12 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=1.59
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=1.59
X19 VTAIL.t6 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=1.59
R0 B.n633 B.n632 585
R1 B.n234 B.n101 585
R2 B.n233 B.n232 585
R3 B.n231 B.n230 585
R4 B.n229 B.n228 585
R5 B.n227 B.n226 585
R6 B.n225 B.n224 585
R7 B.n223 B.n222 585
R8 B.n221 B.n220 585
R9 B.n219 B.n218 585
R10 B.n217 B.n216 585
R11 B.n215 B.n214 585
R12 B.n213 B.n212 585
R13 B.n211 B.n210 585
R14 B.n209 B.n208 585
R15 B.n207 B.n206 585
R16 B.n205 B.n204 585
R17 B.n203 B.n202 585
R18 B.n201 B.n200 585
R19 B.n199 B.n198 585
R20 B.n197 B.n196 585
R21 B.n195 B.n194 585
R22 B.n193 B.n192 585
R23 B.n191 B.n190 585
R24 B.n189 B.n188 585
R25 B.n187 B.n186 585
R26 B.n185 B.n184 585
R27 B.n183 B.n182 585
R28 B.n181 B.n180 585
R29 B.n179 B.n178 585
R30 B.n177 B.n176 585
R31 B.n175 B.n174 585
R32 B.n173 B.n172 585
R33 B.n171 B.n170 585
R34 B.n169 B.n168 585
R35 B.n167 B.n166 585
R36 B.n165 B.n164 585
R37 B.n163 B.n162 585
R38 B.n161 B.n160 585
R39 B.n159 B.n158 585
R40 B.n157 B.n156 585
R41 B.n155 B.n154 585
R42 B.n153 B.n152 585
R43 B.n151 B.n150 585
R44 B.n149 B.n148 585
R45 B.n147 B.n146 585
R46 B.n145 B.n144 585
R47 B.n143 B.n142 585
R48 B.n141 B.n140 585
R49 B.n139 B.n138 585
R50 B.n137 B.n136 585
R51 B.n135 B.n134 585
R52 B.n133 B.n132 585
R53 B.n131 B.n130 585
R54 B.n129 B.n128 585
R55 B.n127 B.n126 585
R56 B.n125 B.n124 585
R57 B.n123 B.n122 585
R58 B.n121 B.n120 585
R59 B.n119 B.n118 585
R60 B.n117 B.n116 585
R61 B.n115 B.n114 585
R62 B.n113 B.n112 585
R63 B.n111 B.n110 585
R64 B.n109 B.n108 585
R65 B.n67 B.n66 585
R66 B.n631 B.n68 585
R67 B.n636 B.n68 585
R68 B.n630 B.n629 585
R69 B.n629 B.n64 585
R70 B.n628 B.n63 585
R71 B.n642 B.n63 585
R72 B.n627 B.n62 585
R73 B.n643 B.n62 585
R74 B.n626 B.n61 585
R75 B.n644 B.n61 585
R76 B.n625 B.n624 585
R77 B.n624 B.n57 585
R78 B.n623 B.n56 585
R79 B.n650 B.n56 585
R80 B.n622 B.n55 585
R81 B.n651 B.n55 585
R82 B.n621 B.n54 585
R83 B.n652 B.n54 585
R84 B.n620 B.n619 585
R85 B.n619 B.n50 585
R86 B.n618 B.n49 585
R87 B.n658 B.n49 585
R88 B.n617 B.n48 585
R89 B.n659 B.n48 585
R90 B.n616 B.n47 585
R91 B.n660 B.n47 585
R92 B.n615 B.n614 585
R93 B.n614 B.n43 585
R94 B.n613 B.n42 585
R95 B.n666 B.n42 585
R96 B.n612 B.n41 585
R97 B.n667 B.n41 585
R98 B.n611 B.n40 585
R99 B.n668 B.n40 585
R100 B.n610 B.n609 585
R101 B.n609 B.n36 585
R102 B.n608 B.n35 585
R103 B.n674 B.n35 585
R104 B.n607 B.n34 585
R105 B.n675 B.n34 585
R106 B.n606 B.n33 585
R107 B.n676 B.n33 585
R108 B.n605 B.n604 585
R109 B.n604 B.n29 585
R110 B.n603 B.n28 585
R111 B.n682 B.n28 585
R112 B.n602 B.n27 585
R113 B.n683 B.n27 585
R114 B.n601 B.n26 585
R115 B.n684 B.n26 585
R116 B.n600 B.n599 585
R117 B.n599 B.n22 585
R118 B.n598 B.n21 585
R119 B.n690 B.n21 585
R120 B.n597 B.n20 585
R121 B.n691 B.n20 585
R122 B.n596 B.n19 585
R123 B.n692 B.n19 585
R124 B.n595 B.n594 585
R125 B.n594 B.n15 585
R126 B.n593 B.n14 585
R127 B.n698 B.n14 585
R128 B.n592 B.n13 585
R129 B.n699 B.n13 585
R130 B.n591 B.n12 585
R131 B.n700 B.n12 585
R132 B.n590 B.n589 585
R133 B.n589 B.n588 585
R134 B.n587 B.n586 585
R135 B.n587 B.n8 585
R136 B.n585 B.n7 585
R137 B.n707 B.n7 585
R138 B.n584 B.n6 585
R139 B.n708 B.n6 585
R140 B.n583 B.n5 585
R141 B.n709 B.n5 585
R142 B.n582 B.n581 585
R143 B.n581 B.n4 585
R144 B.n580 B.n235 585
R145 B.n580 B.n579 585
R146 B.n570 B.n236 585
R147 B.n237 B.n236 585
R148 B.n572 B.n571 585
R149 B.n573 B.n572 585
R150 B.n569 B.n242 585
R151 B.n242 B.n241 585
R152 B.n568 B.n567 585
R153 B.n567 B.n566 585
R154 B.n244 B.n243 585
R155 B.n245 B.n244 585
R156 B.n559 B.n558 585
R157 B.n560 B.n559 585
R158 B.n557 B.n250 585
R159 B.n250 B.n249 585
R160 B.n556 B.n555 585
R161 B.n555 B.n554 585
R162 B.n252 B.n251 585
R163 B.n253 B.n252 585
R164 B.n547 B.n546 585
R165 B.n548 B.n547 585
R166 B.n545 B.n258 585
R167 B.n258 B.n257 585
R168 B.n544 B.n543 585
R169 B.n543 B.n542 585
R170 B.n260 B.n259 585
R171 B.n261 B.n260 585
R172 B.n535 B.n534 585
R173 B.n536 B.n535 585
R174 B.n533 B.n266 585
R175 B.n266 B.n265 585
R176 B.n532 B.n531 585
R177 B.n531 B.n530 585
R178 B.n268 B.n267 585
R179 B.n269 B.n268 585
R180 B.n523 B.n522 585
R181 B.n524 B.n523 585
R182 B.n521 B.n273 585
R183 B.n277 B.n273 585
R184 B.n520 B.n519 585
R185 B.n519 B.n518 585
R186 B.n275 B.n274 585
R187 B.n276 B.n275 585
R188 B.n511 B.n510 585
R189 B.n512 B.n511 585
R190 B.n509 B.n282 585
R191 B.n282 B.n281 585
R192 B.n508 B.n507 585
R193 B.n507 B.n506 585
R194 B.n284 B.n283 585
R195 B.n285 B.n284 585
R196 B.n499 B.n498 585
R197 B.n500 B.n499 585
R198 B.n497 B.n290 585
R199 B.n290 B.n289 585
R200 B.n496 B.n495 585
R201 B.n495 B.n494 585
R202 B.n292 B.n291 585
R203 B.n293 B.n292 585
R204 B.n487 B.n486 585
R205 B.n488 B.n487 585
R206 B.n485 B.n298 585
R207 B.n298 B.n297 585
R208 B.n484 B.n483 585
R209 B.n483 B.n482 585
R210 B.n300 B.n299 585
R211 B.n301 B.n300 585
R212 B.n475 B.n474 585
R213 B.n476 B.n475 585
R214 B.n304 B.n303 585
R215 B.n343 B.n341 585
R216 B.n344 B.n340 585
R217 B.n344 B.n305 585
R218 B.n347 B.n346 585
R219 B.n348 B.n339 585
R220 B.n350 B.n349 585
R221 B.n352 B.n338 585
R222 B.n355 B.n354 585
R223 B.n356 B.n337 585
R224 B.n358 B.n357 585
R225 B.n360 B.n336 585
R226 B.n363 B.n362 585
R227 B.n364 B.n335 585
R228 B.n366 B.n365 585
R229 B.n368 B.n334 585
R230 B.n371 B.n370 585
R231 B.n372 B.n333 585
R232 B.n374 B.n373 585
R233 B.n376 B.n332 585
R234 B.n379 B.n378 585
R235 B.n380 B.n331 585
R236 B.n382 B.n381 585
R237 B.n384 B.n330 585
R238 B.n387 B.n386 585
R239 B.n388 B.n329 585
R240 B.n390 B.n389 585
R241 B.n392 B.n328 585
R242 B.n395 B.n394 585
R243 B.n397 B.n325 585
R244 B.n399 B.n398 585
R245 B.n401 B.n324 585
R246 B.n404 B.n403 585
R247 B.n405 B.n323 585
R248 B.n407 B.n406 585
R249 B.n409 B.n322 585
R250 B.n412 B.n411 585
R251 B.n413 B.n321 585
R252 B.n418 B.n417 585
R253 B.n420 B.n320 585
R254 B.n423 B.n422 585
R255 B.n424 B.n319 585
R256 B.n426 B.n425 585
R257 B.n428 B.n318 585
R258 B.n431 B.n430 585
R259 B.n432 B.n317 585
R260 B.n434 B.n433 585
R261 B.n436 B.n316 585
R262 B.n439 B.n438 585
R263 B.n440 B.n315 585
R264 B.n442 B.n441 585
R265 B.n444 B.n314 585
R266 B.n447 B.n446 585
R267 B.n448 B.n313 585
R268 B.n450 B.n449 585
R269 B.n452 B.n312 585
R270 B.n455 B.n454 585
R271 B.n456 B.n311 585
R272 B.n458 B.n457 585
R273 B.n460 B.n310 585
R274 B.n463 B.n462 585
R275 B.n464 B.n309 585
R276 B.n466 B.n465 585
R277 B.n468 B.n308 585
R278 B.n469 B.n307 585
R279 B.n472 B.n471 585
R280 B.n473 B.n306 585
R281 B.n306 B.n305 585
R282 B.n478 B.n477 585
R283 B.n477 B.n476 585
R284 B.n479 B.n302 585
R285 B.n302 B.n301 585
R286 B.n481 B.n480 585
R287 B.n482 B.n481 585
R288 B.n296 B.n295 585
R289 B.n297 B.n296 585
R290 B.n490 B.n489 585
R291 B.n489 B.n488 585
R292 B.n491 B.n294 585
R293 B.n294 B.n293 585
R294 B.n493 B.n492 585
R295 B.n494 B.n493 585
R296 B.n288 B.n287 585
R297 B.n289 B.n288 585
R298 B.n502 B.n501 585
R299 B.n501 B.n500 585
R300 B.n503 B.n286 585
R301 B.n286 B.n285 585
R302 B.n505 B.n504 585
R303 B.n506 B.n505 585
R304 B.n280 B.n279 585
R305 B.n281 B.n280 585
R306 B.n514 B.n513 585
R307 B.n513 B.n512 585
R308 B.n515 B.n278 585
R309 B.n278 B.n276 585
R310 B.n517 B.n516 585
R311 B.n518 B.n517 585
R312 B.n272 B.n271 585
R313 B.n277 B.n272 585
R314 B.n526 B.n525 585
R315 B.n525 B.n524 585
R316 B.n527 B.n270 585
R317 B.n270 B.n269 585
R318 B.n529 B.n528 585
R319 B.n530 B.n529 585
R320 B.n264 B.n263 585
R321 B.n265 B.n264 585
R322 B.n538 B.n537 585
R323 B.n537 B.n536 585
R324 B.n539 B.n262 585
R325 B.n262 B.n261 585
R326 B.n541 B.n540 585
R327 B.n542 B.n541 585
R328 B.n256 B.n255 585
R329 B.n257 B.n256 585
R330 B.n550 B.n549 585
R331 B.n549 B.n548 585
R332 B.n551 B.n254 585
R333 B.n254 B.n253 585
R334 B.n553 B.n552 585
R335 B.n554 B.n553 585
R336 B.n248 B.n247 585
R337 B.n249 B.n248 585
R338 B.n562 B.n561 585
R339 B.n561 B.n560 585
R340 B.n563 B.n246 585
R341 B.n246 B.n245 585
R342 B.n565 B.n564 585
R343 B.n566 B.n565 585
R344 B.n240 B.n239 585
R345 B.n241 B.n240 585
R346 B.n575 B.n574 585
R347 B.n574 B.n573 585
R348 B.n576 B.n238 585
R349 B.n238 B.n237 585
R350 B.n578 B.n577 585
R351 B.n579 B.n578 585
R352 B.n3 B.n0 585
R353 B.n4 B.n3 585
R354 B.n706 B.n1 585
R355 B.n707 B.n706 585
R356 B.n705 B.n704 585
R357 B.n705 B.n8 585
R358 B.n703 B.n9 585
R359 B.n588 B.n9 585
R360 B.n702 B.n701 585
R361 B.n701 B.n700 585
R362 B.n11 B.n10 585
R363 B.n699 B.n11 585
R364 B.n697 B.n696 585
R365 B.n698 B.n697 585
R366 B.n695 B.n16 585
R367 B.n16 B.n15 585
R368 B.n694 B.n693 585
R369 B.n693 B.n692 585
R370 B.n18 B.n17 585
R371 B.n691 B.n18 585
R372 B.n689 B.n688 585
R373 B.n690 B.n689 585
R374 B.n687 B.n23 585
R375 B.n23 B.n22 585
R376 B.n686 B.n685 585
R377 B.n685 B.n684 585
R378 B.n25 B.n24 585
R379 B.n683 B.n25 585
R380 B.n681 B.n680 585
R381 B.n682 B.n681 585
R382 B.n679 B.n30 585
R383 B.n30 B.n29 585
R384 B.n678 B.n677 585
R385 B.n677 B.n676 585
R386 B.n32 B.n31 585
R387 B.n675 B.n32 585
R388 B.n673 B.n672 585
R389 B.n674 B.n673 585
R390 B.n671 B.n37 585
R391 B.n37 B.n36 585
R392 B.n670 B.n669 585
R393 B.n669 B.n668 585
R394 B.n39 B.n38 585
R395 B.n667 B.n39 585
R396 B.n665 B.n664 585
R397 B.n666 B.n665 585
R398 B.n663 B.n44 585
R399 B.n44 B.n43 585
R400 B.n662 B.n661 585
R401 B.n661 B.n660 585
R402 B.n46 B.n45 585
R403 B.n659 B.n46 585
R404 B.n657 B.n656 585
R405 B.n658 B.n657 585
R406 B.n655 B.n51 585
R407 B.n51 B.n50 585
R408 B.n654 B.n653 585
R409 B.n653 B.n652 585
R410 B.n53 B.n52 585
R411 B.n651 B.n53 585
R412 B.n649 B.n648 585
R413 B.n650 B.n649 585
R414 B.n647 B.n58 585
R415 B.n58 B.n57 585
R416 B.n646 B.n645 585
R417 B.n645 B.n644 585
R418 B.n60 B.n59 585
R419 B.n643 B.n60 585
R420 B.n641 B.n640 585
R421 B.n642 B.n641 585
R422 B.n639 B.n65 585
R423 B.n65 B.n64 585
R424 B.n638 B.n637 585
R425 B.n637 B.n636 585
R426 B.n710 B.n709 585
R427 B.n708 B.n2 585
R428 B.n637 B.n67 487.695
R429 B.n633 B.n68 487.695
R430 B.n475 B.n306 487.695
R431 B.n477 B.n304 487.695
R432 B.n105 B.t19 318.985
R433 B.n102 B.t8 318.985
R434 B.n414 B.t12 318.985
R435 B.n326 B.t16 318.985
R436 B.n635 B.n634 256.663
R437 B.n635 B.n100 256.663
R438 B.n635 B.n99 256.663
R439 B.n635 B.n98 256.663
R440 B.n635 B.n97 256.663
R441 B.n635 B.n96 256.663
R442 B.n635 B.n95 256.663
R443 B.n635 B.n94 256.663
R444 B.n635 B.n93 256.663
R445 B.n635 B.n92 256.663
R446 B.n635 B.n91 256.663
R447 B.n635 B.n90 256.663
R448 B.n635 B.n89 256.663
R449 B.n635 B.n88 256.663
R450 B.n635 B.n87 256.663
R451 B.n635 B.n86 256.663
R452 B.n635 B.n85 256.663
R453 B.n635 B.n84 256.663
R454 B.n635 B.n83 256.663
R455 B.n635 B.n82 256.663
R456 B.n635 B.n81 256.663
R457 B.n635 B.n80 256.663
R458 B.n635 B.n79 256.663
R459 B.n635 B.n78 256.663
R460 B.n635 B.n77 256.663
R461 B.n635 B.n76 256.663
R462 B.n635 B.n75 256.663
R463 B.n635 B.n74 256.663
R464 B.n635 B.n73 256.663
R465 B.n635 B.n72 256.663
R466 B.n635 B.n71 256.663
R467 B.n635 B.n70 256.663
R468 B.n635 B.n69 256.663
R469 B.n342 B.n305 256.663
R470 B.n345 B.n305 256.663
R471 B.n351 B.n305 256.663
R472 B.n353 B.n305 256.663
R473 B.n359 B.n305 256.663
R474 B.n361 B.n305 256.663
R475 B.n367 B.n305 256.663
R476 B.n369 B.n305 256.663
R477 B.n375 B.n305 256.663
R478 B.n377 B.n305 256.663
R479 B.n383 B.n305 256.663
R480 B.n385 B.n305 256.663
R481 B.n391 B.n305 256.663
R482 B.n393 B.n305 256.663
R483 B.n400 B.n305 256.663
R484 B.n402 B.n305 256.663
R485 B.n408 B.n305 256.663
R486 B.n410 B.n305 256.663
R487 B.n419 B.n305 256.663
R488 B.n421 B.n305 256.663
R489 B.n427 B.n305 256.663
R490 B.n429 B.n305 256.663
R491 B.n435 B.n305 256.663
R492 B.n437 B.n305 256.663
R493 B.n443 B.n305 256.663
R494 B.n445 B.n305 256.663
R495 B.n451 B.n305 256.663
R496 B.n453 B.n305 256.663
R497 B.n459 B.n305 256.663
R498 B.n461 B.n305 256.663
R499 B.n467 B.n305 256.663
R500 B.n470 B.n305 256.663
R501 B.n712 B.n711 256.663
R502 B.n102 B.t10 241.732
R503 B.n414 B.t15 241.732
R504 B.n105 B.t20 241.732
R505 B.n326 B.t18 241.732
R506 B.n103 B.t11 204.494
R507 B.n415 B.t14 204.494
R508 B.n106 B.t21 204.494
R509 B.n327 B.t17 204.494
R510 B.n110 B.n109 163.367
R511 B.n114 B.n113 163.367
R512 B.n118 B.n117 163.367
R513 B.n122 B.n121 163.367
R514 B.n126 B.n125 163.367
R515 B.n130 B.n129 163.367
R516 B.n134 B.n133 163.367
R517 B.n138 B.n137 163.367
R518 B.n142 B.n141 163.367
R519 B.n146 B.n145 163.367
R520 B.n150 B.n149 163.367
R521 B.n154 B.n153 163.367
R522 B.n158 B.n157 163.367
R523 B.n162 B.n161 163.367
R524 B.n166 B.n165 163.367
R525 B.n170 B.n169 163.367
R526 B.n174 B.n173 163.367
R527 B.n178 B.n177 163.367
R528 B.n182 B.n181 163.367
R529 B.n186 B.n185 163.367
R530 B.n190 B.n189 163.367
R531 B.n194 B.n193 163.367
R532 B.n198 B.n197 163.367
R533 B.n202 B.n201 163.367
R534 B.n206 B.n205 163.367
R535 B.n210 B.n209 163.367
R536 B.n214 B.n213 163.367
R537 B.n218 B.n217 163.367
R538 B.n222 B.n221 163.367
R539 B.n226 B.n225 163.367
R540 B.n230 B.n229 163.367
R541 B.n232 B.n101 163.367
R542 B.n475 B.n300 163.367
R543 B.n483 B.n300 163.367
R544 B.n483 B.n298 163.367
R545 B.n487 B.n298 163.367
R546 B.n487 B.n292 163.367
R547 B.n495 B.n292 163.367
R548 B.n495 B.n290 163.367
R549 B.n499 B.n290 163.367
R550 B.n499 B.n284 163.367
R551 B.n507 B.n284 163.367
R552 B.n507 B.n282 163.367
R553 B.n511 B.n282 163.367
R554 B.n511 B.n275 163.367
R555 B.n519 B.n275 163.367
R556 B.n519 B.n273 163.367
R557 B.n523 B.n273 163.367
R558 B.n523 B.n268 163.367
R559 B.n531 B.n268 163.367
R560 B.n531 B.n266 163.367
R561 B.n535 B.n266 163.367
R562 B.n535 B.n260 163.367
R563 B.n543 B.n260 163.367
R564 B.n543 B.n258 163.367
R565 B.n547 B.n258 163.367
R566 B.n547 B.n252 163.367
R567 B.n555 B.n252 163.367
R568 B.n555 B.n250 163.367
R569 B.n559 B.n250 163.367
R570 B.n559 B.n244 163.367
R571 B.n567 B.n244 163.367
R572 B.n567 B.n242 163.367
R573 B.n572 B.n242 163.367
R574 B.n572 B.n236 163.367
R575 B.n580 B.n236 163.367
R576 B.n581 B.n580 163.367
R577 B.n581 B.n5 163.367
R578 B.n6 B.n5 163.367
R579 B.n7 B.n6 163.367
R580 B.n587 B.n7 163.367
R581 B.n589 B.n587 163.367
R582 B.n589 B.n12 163.367
R583 B.n13 B.n12 163.367
R584 B.n14 B.n13 163.367
R585 B.n594 B.n14 163.367
R586 B.n594 B.n19 163.367
R587 B.n20 B.n19 163.367
R588 B.n21 B.n20 163.367
R589 B.n599 B.n21 163.367
R590 B.n599 B.n26 163.367
R591 B.n27 B.n26 163.367
R592 B.n28 B.n27 163.367
R593 B.n604 B.n28 163.367
R594 B.n604 B.n33 163.367
R595 B.n34 B.n33 163.367
R596 B.n35 B.n34 163.367
R597 B.n609 B.n35 163.367
R598 B.n609 B.n40 163.367
R599 B.n41 B.n40 163.367
R600 B.n42 B.n41 163.367
R601 B.n614 B.n42 163.367
R602 B.n614 B.n47 163.367
R603 B.n48 B.n47 163.367
R604 B.n49 B.n48 163.367
R605 B.n619 B.n49 163.367
R606 B.n619 B.n54 163.367
R607 B.n55 B.n54 163.367
R608 B.n56 B.n55 163.367
R609 B.n624 B.n56 163.367
R610 B.n624 B.n61 163.367
R611 B.n62 B.n61 163.367
R612 B.n63 B.n62 163.367
R613 B.n629 B.n63 163.367
R614 B.n629 B.n68 163.367
R615 B.n344 B.n343 163.367
R616 B.n346 B.n344 163.367
R617 B.n350 B.n339 163.367
R618 B.n354 B.n352 163.367
R619 B.n358 B.n337 163.367
R620 B.n362 B.n360 163.367
R621 B.n366 B.n335 163.367
R622 B.n370 B.n368 163.367
R623 B.n374 B.n333 163.367
R624 B.n378 B.n376 163.367
R625 B.n382 B.n331 163.367
R626 B.n386 B.n384 163.367
R627 B.n390 B.n329 163.367
R628 B.n394 B.n392 163.367
R629 B.n399 B.n325 163.367
R630 B.n403 B.n401 163.367
R631 B.n407 B.n323 163.367
R632 B.n411 B.n409 163.367
R633 B.n418 B.n321 163.367
R634 B.n422 B.n420 163.367
R635 B.n426 B.n319 163.367
R636 B.n430 B.n428 163.367
R637 B.n434 B.n317 163.367
R638 B.n438 B.n436 163.367
R639 B.n442 B.n315 163.367
R640 B.n446 B.n444 163.367
R641 B.n450 B.n313 163.367
R642 B.n454 B.n452 163.367
R643 B.n458 B.n311 163.367
R644 B.n462 B.n460 163.367
R645 B.n466 B.n309 163.367
R646 B.n469 B.n468 163.367
R647 B.n471 B.n306 163.367
R648 B.n477 B.n302 163.367
R649 B.n481 B.n302 163.367
R650 B.n481 B.n296 163.367
R651 B.n489 B.n296 163.367
R652 B.n489 B.n294 163.367
R653 B.n493 B.n294 163.367
R654 B.n493 B.n288 163.367
R655 B.n501 B.n288 163.367
R656 B.n501 B.n286 163.367
R657 B.n505 B.n286 163.367
R658 B.n505 B.n280 163.367
R659 B.n513 B.n280 163.367
R660 B.n513 B.n278 163.367
R661 B.n517 B.n278 163.367
R662 B.n517 B.n272 163.367
R663 B.n525 B.n272 163.367
R664 B.n525 B.n270 163.367
R665 B.n529 B.n270 163.367
R666 B.n529 B.n264 163.367
R667 B.n537 B.n264 163.367
R668 B.n537 B.n262 163.367
R669 B.n541 B.n262 163.367
R670 B.n541 B.n256 163.367
R671 B.n549 B.n256 163.367
R672 B.n549 B.n254 163.367
R673 B.n553 B.n254 163.367
R674 B.n553 B.n248 163.367
R675 B.n561 B.n248 163.367
R676 B.n561 B.n246 163.367
R677 B.n565 B.n246 163.367
R678 B.n565 B.n240 163.367
R679 B.n574 B.n240 163.367
R680 B.n574 B.n238 163.367
R681 B.n578 B.n238 163.367
R682 B.n578 B.n3 163.367
R683 B.n710 B.n3 163.367
R684 B.n706 B.n2 163.367
R685 B.n706 B.n705 163.367
R686 B.n705 B.n9 163.367
R687 B.n701 B.n9 163.367
R688 B.n701 B.n11 163.367
R689 B.n697 B.n11 163.367
R690 B.n697 B.n16 163.367
R691 B.n693 B.n16 163.367
R692 B.n693 B.n18 163.367
R693 B.n689 B.n18 163.367
R694 B.n689 B.n23 163.367
R695 B.n685 B.n23 163.367
R696 B.n685 B.n25 163.367
R697 B.n681 B.n25 163.367
R698 B.n681 B.n30 163.367
R699 B.n677 B.n30 163.367
R700 B.n677 B.n32 163.367
R701 B.n673 B.n32 163.367
R702 B.n673 B.n37 163.367
R703 B.n669 B.n37 163.367
R704 B.n669 B.n39 163.367
R705 B.n665 B.n39 163.367
R706 B.n665 B.n44 163.367
R707 B.n661 B.n44 163.367
R708 B.n661 B.n46 163.367
R709 B.n657 B.n46 163.367
R710 B.n657 B.n51 163.367
R711 B.n653 B.n51 163.367
R712 B.n653 B.n53 163.367
R713 B.n649 B.n53 163.367
R714 B.n649 B.n58 163.367
R715 B.n645 B.n58 163.367
R716 B.n645 B.n60 163.367
R717 B.n641 B.n60 163.367
R718 B.n641 B.n65 163.367
R719 B.n637 B.n65 163.367
R720 B.n476 B.n305 97.5289
R721 B.n636 B.n635 97.5289
R722 B.n69 B.n67 71.676
R723 B.n110 B.n70 71.676
R724 B.n114 B.n71 71.676
R725 B.n118 B.n72 71.676
R726 B.n122 B.n73 71.676
R727 B.n126 B.n74 71.676
R728 B.n130 B.n75 71.676
R729 B.n134 B.n76 71.676
R730 B.n138 B.n77 71.676
R731 B.n142 B.n78 71.676
R732 B.n146 B.n79 71.676
R733 B.n150 B.n80 71.676
R734 B.n154 B.n81 71.676
R735 B.n158 B.n82 71.676
R736 B.n162 B.n83 71.676
R737 B.n166 B.n84 71.676
R738 B.n170 B.n85 71.676
R739 B.n174 B.n86 71.676
R740 B.n178 B.n87 71.676
R741 B.n182 B.n88 71.676
R742 B.n186 B.n89 71.676
R743 B.n190 B.n90 71.676
R744 B.n194 B.n91 71.676
R745 B.n198 B.n92 71.676
R746 B.n202 B.n93 71.676
R747 B.n206 B.n94 71.676
R748 B.n210 B.n95 71.676
R749 B.n214 B.n96 71.676
R750 B.n218 B.n97 71.676
R751 B.n222 B.n98 71.676
R752 B.n226 B.n99 71.676
R753 B.n230 B.n100 71.676
R754 B.n634 B.n101 71.676
R755 B.n634 B.n633 71.676
R756 B.n232 B.n100 71.676
R757 B.n229 B.n99 71.676
R758 B.n225 B.n98 71.676
R759 B.n221 B.n97 71.676
R760 B.n217 B.n96 71.676
R761 B.n213 B.n95 71.676
R762 B.n209 B.n94 71.676
R763 B.n205 B.n93 71.676
R764 B.n201 B.n92 71.676
R765 B.n197 B.n91 71.676
R766 B.n193 B.n90 71.676
R767 B.n189 B.n89 71.676
R768 B.n185 B.n88 71.676
R769 B.n181 B.n87 71.676
R770 B.n177 B.n86 71.676
R771 B.n173 B.n85 71.676
R772 B.n169 B.n84 71.676
R773 B.n165 B.n83 71.676
R774 B.n161 B.n82 71.676
R775 B.n157 B.n81 71.676
R776 B.n153 B.n80 71.676
R777 B.n149 B.n79 71.676
R778 B.n145 B.n78 71.676
R779 B.n141 B.n77 71.676
R780 B.n137 B.n76 71.676
R781 B.n133 B.n75 71.676
R782 B.n129 B.n74 71.676
R783 B.n125 B.n73 71.676
R784 B.n121 B.n72 71.676
R785 B.n117 B.n71 71.676
R786 B.n113 B.n70 71.676
R787 B.n109 B.n69 71.676
R788 B.n342 B.n304 71.676
R789 B.n346 B.n345 71.676
R790 B.n351 B.n350 71.676
R791 B.n354 B.n353 71.676
R792 B.n359 B.n358 71.676
R793 B.n362 B.n361 71.676
R794 B.n367 B.n366 71.676
R795 B.n370 B.n369 71.676
R796 B.n375 B.n374 71.676
R797 B.n378 B.n377 71.676
R798 B.n383 B.n382 71.676
R799 B.n386 B.n385 71.676
R800 B.n391 B.n390 71.676
R801 B.n394 B.n393 71.676
R802 B.n400 B.n399 71.676
R803 B.n403 B.n402 71.676
R804 B.n408 B.n407 71.676
R805 B.n411 B.n410 71.676
R806 B.n419 B.n418 71.676
R807 B.n422 B.n421 71.676
R808 B.n427 B.n426 71.676
R809 B.n430 B.n429 71.676
R810 B.n435 B.n434 71.676
R811 B.n438 B.n437 71.676
R812 B.n443 B.n442 71.676
R813 B.n446 B.n445 71.676
R814 B.n451 B.n450 71.676
R815 B.n454 B.n453 71.676
R816 B.n459 B.n458 71.676
R817 B.n462 B.n461 71.676
R818 B.n467 B.n466 71.676
R819 B.n470 B.n469 71.676
R820 B.n343 B.n342 71.676
R821 B.n345 B.n339 71.676
R822 B.n352 B.n351 71.676
R823 B.n353 B.n337 71.676
R824 B.n360 B.n359 71.676
R825 B.n361 B.n335 71.676
R826 B.n368 B.n367 71.676
R827 B.n369 B.n333 71.676
R828 B.n376 B.n375 71.676
R829 B.n377 B.n331 71.676
R830 B.n384 B.n383 71.676
R831 B.n385 B.n329 71.676
R832 B.n392 B.n391 71.676
R833 B.n393 B.n325 71.676
R834 B.n401 B.n400 71.676
R835 B.n402 B.n323 71.676
R836 B.n409 B.n408 71.676
R837 B.n410 B.n321 71.676
R838 B.n420 B.n419 71.676
R839 B.n421 B.n319 71.676
R840 B.n428 B.n427 71.676
R841 B.n429 B.n317 71.676
R842 B.n436 B.n435 71.676
R843 B.n437 B.n315 71.676
R844 B.n444 B.n443 71.676
R845 B.n445 B.n313 71.676
R846 B.n452 B.n451 71.676
R847 B.n453 B.n311 71.676
R848 B.n460 B.n459 71.676
R849 B.n461 B.n309 71.676
R850 B.n468 B.n467 71.676
R851 B.n471 B.n470 71.676
R852 B.n711 B.n710 71.676
R853 B.n711 B.n2 71.676
R854 B.n107 B.n106 59.5399
R855 B.n104 B.n103 59.5399
R856 B.n416 B.n415 59.5399
R857 B.n396 B.n327 59.5399
R858 B.n476 B.n301 58.6902
R859 B.n482 B.n301 58.6902
R860 B.n482 B.n297 58.6902
R861 B.n488 B.n297 58.6902
R862 B.n488 B.n293 58.6902
R863 B.n494 B.n293 58.6902
R864 B.n500 B.n289 58.6902
R865 B.n500 B.n285 58.6902
R866 B.n506 B.n285 58.6902
R867 B.n506 B.n281 58.6902
R868 B.n512 B.n281 58.6902
R869 B.n512 B.n276 58.6902
R870 B.n518 B.n276 58.6902
R871 B.n518 B.n277 58.6902
R872 B.n524 B.n269 58.6902
R873 B.n530 B.n269 58.6902
R874 B.n530 B.n265 58.6902
R875 B.n536 B.n265 58.6902
R876 B.n542 B.n261 58.6902
R877 B.n542 B.n257 58.6902
R878 B.n548 B.n257 58.6902
R879 B.n548 B.n253 58.6902
R880 B.n554 B.n253 58.6902
R881 B.n560 B.n249 58.6902
R882 B.n560 B.n245 58.6902
R883 B.n566 B.n245 58.6902
R884 B.n566 B.n241 58.6902
R885 B.n573 B.n241 58.6902
R886 B.n579 B.n237 58.6902
R887 B.n579 B.n4 58.6902
R888 B.n709 B.n4 58.6902
R889 B.n709 B.n708 58.6902
R890 B.n708 B.n707 58.6902
R891 B.n707 B.n8 58.6902
R892 B.n588 B.n8 58.6902
R893 B.n700 B.n699 58.6902
R894 B.n699 B.n698 58.6902
R895 B.n698 B.n15 58.6902
R896 B.n692 B.n15 58.6902
R897 B.n692 B.n691 58.6902
R898 B.n690 B.n22 58.6902
R899 B.n684 B.n22 58.6902
R900 B.n684 B.n683 58.6902
R901 B.n683 B.n682 58.6902
R902 B.n682 B.n29 58.6902
R903 B.n676 B.n675 58.6902
R904 B.n675 B.n674 58.6902
R905 B.n674 B.n36 58.6902
R906 B.n668 B.n36 58.6902
R907 B.n667 B.n666 58.6902
R908 B.n666 B.n43 58.6902
R909 B.n660 B.n43 58.6902
R910 B.n660 B.n659 58.6902
R911 B.n659 B.n658 58.6902
R912 B.n658 B.n50 58.6902
R913 B.n652 B.n50 58.6902
R914 B.n652 B.n651 58.6902
R915 B.n650 B.n57 58.6902
R916 B.n644 B.n57 58.6902
R917 B.n644 B.n643 58.6902
R918 B.n643 B.n642 58.6902
R919 B.n642 B.n64 58.6902
R920 B.n636 B.n64 58.6902
R921 B.t4 B.n237 54.3748
R922 B.n588 B.t5 54.3748
R923 B.n524 B.t6 50.9224
R924 B.n668 B.t2 50.9224
R925 B.n536 B.t1 45.7439
R926 B.n676 B.t0 45.7439
R927 B.t13 B.n289 42.2916
R928 B.n651 B.t9 42.2916
R929 B.n106 B.n105 37.2369
R930 B.n103 B.n102 37.2369
R931 B.n415 B.n414 37.2369
R932 B.n327 B.n326 37.2369
R933 B.t3 B.n249 33.6608
R934 B.n691 B.t7 33.6608
R935 B.n478 B.n303 31.6883
R936 B.n474 B.n473 31.6883
R937 B.n632 B.n631 31.6883
R938 B.n638 B.n66 31.6883
R939 B.n554 B.t3 25.0299
R940 B.t7 B.n690 25.0299
R941 B B.n712 18.0485
R942 B.n494 B.t13 16.3991
R943 B.t9 B.n650 16.3991
R944 B.t1 B.n261 12.9468
R945 B.t0 B.n29 12.9468
R946 B.n479 B.n478 10.6151
R947 B.n480 B.n479 10.6151
R948 B.n480 B.n295 10.6151
R949 B.n490 B.n295 10.6151
R950 B.n491 B.n490 10.6151
R951 B.n492 B.n491 10.6151
R952 B.n492 B.n287 10.6151
R953 B.n502 B.n287 10.6151
R954 B.n503 B.n502 10.6151
R955 B.n504 B.n503 10.6151
R956 B.n504 B.n279 10.6151
R957 B.n514 B.n279 10.6151
R958 B.n515 B.n514 10.6151
R959 B.n516 B.n515 10.6151
R960 B.n516 B.n271 10.6151
R961 B.n526 B.n271 10.6151
R962 B.n527 B.n526 10.6151
R963 B.n528 B.n527 10.6151
R964 B.n528 B.n263 10.6151
R965 B.n538 B.n263 10.6151
R966 B.n539 B.n538 10.6151
R967 B.n540 B.n539 10.6151
R968 B.n540 B.n255 10.6151
R969 B.n550 B.n255 10.6151
R970 B.n551 B.n550 10.6151
R971 B.n552 B.n551 10.6151
R972 B.n552 B.n247 10.6151
R973 B.n562 B.n247 10.6151
R974 B.n563 B.n562 10.6151
R975 B.n564 B.n563 10.6151
R976 B.n564 B.n239 10.6151
R977 B.n575 B.n239 10.6151
R978 B.n576 B.n575 10.6151
R979 B.n577 B.n576 10.6151
R980 B.n577 B.n0 10.6151
R981 B.n341 B.n303 10.6151
R982 B.n341 B.n340 10.6151
R983 B.n347 B.n340 10.6151
R984 B.n348 B.n347 10.6151
R985 B.n349 B.n348 10.6151
R986 B.n349 B.n338 10.6151
R987 B.n355 B.n338 10.6151
R988 B.n356 B.n355 10.6151
R989 B.n357 B.n356 10.6151
R990 B.n357 B.n336 10.6151
R991 B.n363 B.n336 10.6151
R992 B.n364 B.n363 10.6151
R993 B.n365 B.n364 10.6151
R994 B.n365 B.n334 10.6151
R995 B.n371 B.n334 10.6151
R996 B.n372 B.n371 10.6151
R997 B.n373 B.n372 10.6151
R998 B.n373 B.n332 10.6151
R999 B.n379 B.n332 10.6151
R1000 B.n380 B.n379 10.6151
R1001 B.n381 B.n380 10.6151
R1002 B.n381 B.n330 10.6151
R1003 B.n387 B.n330 10.6151
R1004 B.n388 B.n387 10.6151
R1005 B.n389 B.n388 10.6151
R1006 B.n389 B.n328 10.6151
R1007 B.n395 B.n328 10.6151
R1008 B.n398 B.n397 10.6151
R1009 B.n398 B.n324 10.6151
R1010 B.n404 B.n324 10.6151
R1011 B.n405 B.n404 10.6151
R1012 B.n406 B.n405 10.6151
R1013 B.n406 B.n322 10.6151
R1014 B.n412 B.n322 10.6151
R1015 B.n413 B.n412 10.6151
R1016 B.n417 B.n413 10.6151
R1017 B.n423 B.n320 10.6151
R1018 B.n424 B.n423 10.6151
R1019 B.n425 B.n424 10.6151
R1020 B.n425 B.n318 10.6151
R1021 B.n431 B.n318 10.6151
R1022 B.n432 B.n431 10.6151
R1023 B.n433 B.n432 10.6151
R1024 B.n433 B.n316 10.6151
R1025 B.n439 B.n316 10.6151
R1026 B.n440 B.n439 10.6151
R1027 B.n441 B.n440 10.6151
R1028 B.n441 B.n314 10.6151
R1029 B.n447 B.n314 10.6151
R1030 B.n448 B.n447 10.6151
R1031 B.n449 B.n448 10.6151
R1032 B.n449 B.n312 10.6151
R1033 B.n455 B.n312 10.6151
R1034 B.n456 B.n455 10.6151
R1035 B.n457 B.n456 10.6151
R1036 B.n457 B.n310 10.6151
R1037 B.n463 B.n310 10.6151
R1038 B.n464 B.n463 10.6151
R1039 B.n465 B.n464 10.6151
R1040 B.n465 B.n308 10.6151
R1041 B.n308 B.n307 10.6151
R1042 B.n472 B.n307 10.6151
R1043 B.n473 B.n472 10.6151
R1044 B.n474 B.n299 10.6151
R1045 B.n484 B.n299 10.6151
R1046 B.n485 B.n484 10.6151
R1047 B.n486 B.n485 10.6151
R1048 B.n486 B.n291 10.6151
R1049 B.n496 B.n291 10.6151
R1050 B.n497 B.n496 10.6151
R1051 B.n498 B.n497 10.6151
R1052 B.n498 B.n283 10.6151
R1053 B.n508 B.n283 10.6151
R1054 B.n509 B.n508 10.6151
R1055 B.n510 B.n509 10.6151
R1056 B.n510 B.n274 10.6151
R1057 B.n520 B.n274 10.6151
R1058 B.n521 B.n520 10.6151
R1059 B.n522 B.n521 10.6151
R1060 B.n522 B.n267 10.6151
R1061 B.n532 B.n267 10.6151
R1062 B.n533 B.n532 10.6151
R1063 B.n534 B.n533 10.6151
R1064 B.n534 B.n259 10.6151
R1065 B.n544 B.n259 10.6151
R1066 B.n545 B.n544 10.6151
R1067 B.n546 B.n545 10.6151
R1068 B.n546 B.n251 10.6151
R1069 B.n556 B.n251 10.6151
R1070 B.n557 B.n556 10.6151
R1071 B.n558 B.n557 10.6151
R1072 B.n558 B.n243 10.6151
R1073 B.n568 B.n243 10.6151
R1074 B.n569 B.n568 10.6151
R1075 B.n571 B.n569 10.6151
R1076 B.n571 B.n570 10.6151
R1077 B.n570 B.n235 10.6151
R1078 B.n582 B.n235 10.6151
R1079 B.n583 B.n582 10.6151
R1080 B.n584 B.n583 10.6151
R1081 B.n585 B.n584 10.6151
R1082 B.n586 B.n585 10.6151
R1083 B.n590 B.n586 10.6151
R1084 B.n591 B.n590 10.6151
R1085 B.n592 B.n591 10.6151
R1086 B.n593 B.n592 10.6151
R1087 B.n595 B.n593 10.6151
R1088 B.n596 B.n595 10.6151
R1089 B.n597 B.n596 10.6151
R1090 B.n598 B.n597 10.6151
R1091 B.n600 B.n598 10.6151
R1092 B.n601 B.n600 10.6151
R1093 B.n602 B.n601 10.6151
R1094 B.n603 B.n602 10.6151
R1095 B.n605 B.n603 10.6151
R1096 B.n606 B.n605 10.6151
R1097 B.n607 B.n606 10.6151
R1098 B.n608 B.n607 10.6151
R1099 B.n610 B.n608 10.6151
R1100 B.n611 B.n610 10.6151
R1101 B.n612 B.n611 10.6151
R1102 B.n613 B.n612 10.6151
R1103 B.n615 B.n613 10.6151
R1104 B.n616 B.n615 10.6151
R1105 B.n617 B.n616 10.6151
R1106 B.n618 B.n617 10.6151
R1107 B.n620 B.n618 10.6151
R1108 B.n621 B.n620 10.6151
R1109 B.n622 B.n621 10.6151
R1110 B.n623 B.n622 10.6151
R1111 B.n625 B.n623 10.6151
R1112 B.n626 B.n625 10.6151
R1113 B.n627 B.n626 10.6151
R1114 B.n628 B.n627 10.6151
R1115 B.n630 B.n628 10.6151
R1116 B.n631 B.n630 10.6151
R1117 B.n704 B.n1 10.6151
R1118 B.n704 B.n703 10.6151
R1119 B.n703 B.n702 10.6151
R1120 B.n702 B.n10 10.6151
R1121 B.n696 B.n10 10.6151
R1122 B.n696 B.n695 10.6151
R1123 B.n695 B.n694 10.6151
R1124 B.n694 B.n17 10.6151
R1125 B.n688 B.n17 10.6151
R1126 B.n688 B.n687 10.6151
R1127 B.n687 B.n686 10.6151
R1128 B.n686 B.n24 10.6151
R1129 B.n680 B.n24 10.6151
R1130 B.n680 B.n679 10.6151
R1131 B.n679 B.n678 10.6151
R1132 B.n678 B.n31 10.6151
R1133 B.n672 B.n31 10.6151
R1134 B.n672 B.n671 10.6151
R1135 B.n671 B.n670 10.6151
R1136 B.n670 B.n38 10.6151
R1137 B.n664 B.n38 10.6151
R1138 B.n664 B.n663 10.6151
R1139 B.n663 B.n662 10.6151
R1140 B.n662 B.n45 10.6151
R1141 B.n656 B.n45 10.6151
R1142 B.n656 B.n655 10.6151
R1143 B.n655 B.n654 10.6151
R1144 B.n654 B.n52 10.6151
R1145 B.n648 B.n52 10.6151
R1146 B.n648 B.n647 10.6151
R1147 B.n647 B.n646 10.6151
R1148 B.n646 B.n59 10.6151
R1149 B.n640 B.n59 10.6151
R1150 B.n640 B.n639 10.6151
R1151 B.n639 B.n638 10.6151
R1152 B.n108 B.n66 10.6151
R1153 B.n111 B.n108 10.6151
R1154 B.n112 B.n111 10.6151
R1155 B.n115 B.n112 10.6151
R1156 B.n116 B.n115 10.6151
R1157 B.n119 B.n116 10.6151
R1158 B.n120 B.n119 10.6151
R1159 B.n123 B.n120 10.6151
R1160 B.n124 B.n123 10.6151
R1161 B.n127 B.n124 10.6151
R1162 B.n128 B.n127 10.6151
R1163 B.n131 B.n128 10.6151
R1164 B.n132 B.n131 10.6151
R1165 B.n135 B.n132 10.6151
R1166 B.n136 B.n135 10.6151
R1167 B.n139 B.n136 10.6151
R1168 B.n140 B.n139 10.6151
R1169 B.n143 B.n140 10.6151
R1170 B.n144 B.n143 10.6151
R1171 B.n147 B.n144 10.6151
R1172 B.n148 B.n147 10.6151
R1173 B.n151 B.n148 10.6151
R1174 B.n152 B.n151 10.6151
R1175 B.n155 B.n152 10.6151
R1176 B.n156 B.n155 10.6151
R1177 B.n159 B.n156 10.6151
R1178 B.n160 B.n159 10.6151
R1179 B.n164 B.n163 10.6151
R1180 B.n167 B.n164 10.6151
R1181 B.n168 B.n167 10.6151
R1182 B.n171 B.n168 10.6151
R1183 B.n172 B.n171 10.6151
R1184 B.n175 B.n172 10.6151
R1185 B.n176 B.n175 10.6151
R1186 B.n179 B.n176 10.6151
R1187 B.n180 B.n179 10.6151
R1188 B.n184 B.n183 10.6151
R1189 B.n187 B.n184 10.6151
R1190 B.n188 B.n187 10.6151
R1191 B.n191 B.n188 10.6151
R1192 B.n192 B.n191 10.6151
R1193 B.n195 B.n192 10.6151
R1194 B.n196 B.n195 10.6151
R1195 B.n199 B.n196 10.6151
R1196 B.n200 B.n199 10.6151
R1197 B.n203 B.n200 10.6151
R1198 B.n204 B.n203 10.6151
R1199 B.n207 B.n204 10.6151
R1200 B.n208 B.n207 10.6151
R1201 B.n211 B.n208 10.6151
R1202 B.n212 B.n211 10.6151
R1203 B.n215 B.n212 10.6151
R1204 B.n216 B.n215 10.6151
R1205 B.n219 B.n216 10.6151
R1206 B.n220 B.n219 10.6151
R1207 B.n223 B.n220 10.6151
R1208 B.n224 B.n223 10.6151
R1209 B.n227 B.n224 10.6151
R1210 B.n228 B.n227 10.6151
R1211 B.n231 B.n228 10.6151
R1212 B.n233 B.n231 10.6151
R1213 B.n234 B.n233 10.6151
R1214 B.n632 B.n234 10.6151
R1215 B.n396 B.n395 9.36635
R1216 B.n416 B.n320 9.36635
R1217 B.n160 B.n107 9.36635
R1218 B.n183 B.n104 9.36635
R1219 B.n712 B.n0 8.11757
R1220 B.n712 B.n1 8.11757
R1221 B.n277 B.t6 7.76825
R1222 B.t2 B.n667 7.76825
R1223 B.n573 B.t4 4.31592
R1224 B.n700 B.t5 4.31592
R1225 B.n397 B.n396 1.24928
R1226 B.n417 B.n416 1.24928
R1227 B.n163 B.n107 1.24928
R1228 B.n180 B.n104 1.24928
R1229 VP.n28 VP.n27 179.406
R1230 VP.n50 VP.n49 179.406
R1231 VP.n26 VP.n25 179.406
R1232 VP.n13 VP.n12 161.3
R1233 VP.n14 VP.n9 161.3
R1234 VP.n16 VP.n15 161.3
R1235 VP.n17 VP.n8 161.3
R1236 VP.n20 VP.n19 161.3
R1237 VP.n21 VP.n7 161.3
R1238 VP.n23 VP.n22 161.3
R1239 VP.n24 VP.n6 161.3
R1240 VP.n48 VP.n0 161.3
R1241 VP.n47 VP.n46 161.3
R1242 VP.n45 VP.n1 161.3
R1243 VP.n44 VP.n43 161.3
R1244 VP.n41 VP.n2 161.3
R1245 VP.n40 VP.n39 161.3
R1246 VP.n38 VP.n3 161.3
R1247 VP.n37 VP.n36 161.3
R1248 VP.n34 VP.n4 161.3
R1249 VP.n33 VP.n32 161.3
R1250 VP.n31 VP.n5 161.3
R1251 VP.n30 VP.n29 161.3
R1252 VP.n10 VP.t7 145.01
R1253 VP.n28 VP.t3 113.225
R1254 VP.n35 VP.t0 113.225
R1255 VP.n42 VP.t1 113.225
R1256 VP.n49 VP.t2 113.225
R1257 VP.n25 VP.t4 113.225
R1258 VP.n18 VP.t5 113.225
R1259 VP.n11 VP.t6 113.225
R1260 VP.n33 VP.n5 56.5193
R1261 VP.n47 VP.n1 56.5193
R1262 VP.n23 VP.n7 56.5193
R1263 VP.n40 VP.n3 56.5193
R1264 VP.n16 VP.n9 56.5193
R1265 VP.n11 VP.n10 55.7366
R1266 VP.n27 VP.n26 42.6293
R1267 VP.n29 VP.n5 24.4675
R1268 VP.n34 VP.n33 24.4675
R1269 VP.n36 VP.n3 24.4675
R1270 VP.n41 VP.n40 24.4675
R1271 VP.n43 VP.n1 24.4675
R1272 VP.n48 VP.n47 24.4675
R1273 VP.n24 VP.n23 24.4675
R1274 VP.n17 VP.n16 24.4675
R1275 VP.n19 VP.n7 24.4675
R1276 VP.n12 VP.n9 24.4675
R1277 VP.n13 VP.n10 18.144
R1278 VP.n35 VP.n34 14.1914
R1279 VP.n43 VP.n42 14.1914
R1280 VP.n19 VP.n18 14.1914
R1281 VP.n36 VP.n35 10.2766
R1282 VP.n42 VP.n41 10.2766
R1283 VP.n18 VP.n17 10.2766
R1284 VP.n12 VP.n11 10.2766
R1285 VP.n29 VP.n28 6.36192
R1286 VP.n49 VP.n48 6.36192
R1287 VP.n25 VP.n24 6.36192
R1288 VP.n14 VP.n13 0.189894
R1289 VP.n15 VP.n14 0.189894
R1290 VP.n15 VP.n8 0.189894
R1291 VP.n20 VP.n8 0.189894
R1292 VP.n21 VP.n20 0.189894
R1293 VP.n22 VP.n21 0.189894
R1294 VP.n22 VP.n6 0.189894
R1295 VP.n26 VP.n6 0.189894
R1296 VP.n30 VP.n27 0.189894
R1297 VP.n31 VP.n30 0.189894
R1298 VP.n32 VP.n31 0.189894
R1299 VP.n32 VP.n4 0.189894
R1300 VP.n37 VP.n4 0.189894
R1301 VP.n38 VP.n37 0.189894
R1302 VP.n39 VP.n38 0.189894
R1303 VP.n39 VP.n2 0.189894
R1304 VP.n44 VP.n2 0.189894
R1305 VP.n45 VP.n44 0.189894
R1306 VP.n46 VP.n45 0.189894
R1307 VP.n46 VP.n0 0.189894
R1308 VP.n50 VP.n0 0.189894
R1309 VP VP.n50 0.0516364
R1310 VTAIL.n322 VTAIL.n288 289.615
R1311 VTAIL.n36 VTAIL.n2 289.615
R1312 VTAIL.n76 VTAIL.n42 289.615
R1313 VTAIL.n118 VTAIL.n84 289.615
R1314 VTAIL.n282 VTAIL.n248 289.615
R1315 VTAIL.n240 VTAIL.n206 289.615
R1316 VTAIL.n200 VTAIL.n166 289.615
R1317 VTAIL.n158 VTAIL.n124 289.615
R1318 VTAIL.n300 VTAIL.n299 185
R1319 VTAIL.n305 VTAIL.n304 185
R1320 VTAIL.n307 VTAIL.n306 185
R1321 VTAIL.n296 VTAIL.n295 185
R1322 VTAIL.n313 VTAIL.n312 185
R1323 VTAIL.n315 VTAIL.n314 185
R1324 VTAIL.n292 VTAIL.n291 185
R1325 VTAIL.n321 VTAIL.n320 185
R1326 VTAIL.n323 VTAIL.n322 185
R1327 VTAIL.n14 VTAIL.n13 185
R1328 VTAIL.n19 VTAIL.n18 185
R1329 VTAIL.n21 VTAIL.n20 185
R1330 VTAIL.n10 VTAIL.n9 185
R1331 VTAIL.n27 VTAIL.n26 185
R1332 VTAIL.n29 VTAIL.n28 185
R1333 VTAIL.n6 VTAIL.n5 185
R1334 VTAIL.n35 VTAIL.n34 185
R1335 VTAIL.n37 VTAIL.n36 185
R1336 VTAIL.n54 VTAIL.n53 185
R1337 VTAIL.n59 VTAIL.n58 185
R1338 VTAIL.n61 VTAIL.n60 185
R1339 VTAIL.n50 VTAIL.n49 185
R1340 VTAIL.n67 VTAIL.n66 185
R1341 VTAIL.n69 VTAIL.n68 185
R1342 VTAIL.n46 VTAIL.n45 185
R1343 VTAIL.n75 VTAIL.n74 185
R1344 VTAIL.n77 VTAIL.n76 185
R1345 VTAIL.n96 VTAIL.n95 185
R1346 VTAIL.n101 VTAIL.n100 185
R1347 VTAIL.n103 VTAIL.n102 185
R1348 VTAIL.n92 VTAIL.n91 185
R1349 VTAIL.n109 VTAIL.n108 185
R1350 VTAIL.n111 VTAIL.n110 185
R1351 VTAIL.n88 VTAIL.n87 185
R1352 VTAIL.n117 VTAIL.n116 185
R1353 VTAIL.n119 VTAIL.n118 185
R1354 VTAIL.n283 VTAIL.n282 185
R1355 VTAIL.n281 VTAIL.n280 185
R1356 VTAIL.n252 VTAIL.n251 185
R1357 VTAIL.n275 VTAIL.n274 185
R1358 VTAIL.n273 VTAIL.n272 185
R1359 VTAIL.n256 VTAIL.n255 185
R1360 VTAIL.n267 VTAIL.n266 185
R1361 VTAIL.n265 VTAIL.n264 185
R1362 VTAIL.n260 VTAIL.n259 185
R1363 VTAIL.n241 VTAIL.n240 185
R1364 VTAIL.n239 VTAIL.n238 185
R1365 VTAIL.n210 VTAIL.n209 185
R1366 VTAIL.n233 VTAIL.n232 185
R1367 VTAIL.n231 VTAIL.n230 185
R1368 VTAIL.n214 VTAIL.n213 185
R1369 VTAIL.n225 VTAIL.n224 185
R1370 VTAIL.n223 VTAIL.n222 185
R1371 VTAIL.n218 VTAIL.n217 185
R1372 VTAIL.n201 VTAIL.n200 185
R1373 VTAIL.n199 VTAIL.n198 185
R1374 VTAIL.n170 VTAIL.n169 185
R1375 VTAIL.n193 VTAIL.n192 185
R1376 VTAIL.n191 VTAIL.n190 185
R1377 VTAIL.n174 VTAIL.n173 185
R1378 VTAIL.n185 VTAIL.n184 185
R1379 VTAIL.n183 VTAIL.n182 185
R1380 VTAIL.n178 VTAIL.n177 185
R1381 VTAIL.n159 VTAIL.n158 185
R1382 VTAIL.n157 VTAIL.n156 185
R1383 VTAIL.n128 VTAIL.n127 185
R1384 VTAIL.n151 VTAIL.n150 185
R1385 VTAIL.n149 VTAIL.n148 185
R1386 VTAIL.n132 VTAIL.n131 185
R1387 VTAIL.n143 VTAIL.n142 185
R1388 VTAIL.n141 VTAIL.n140 185
R1389 VTAIL.n136 VTAIL.n135 185
R1390 VTAIL.n301 VTAIL.t2 147.659
R1391 VTAIL.n15 VTAIL.t6 147.659
R1392 VTAIL.n55 VTAIL.t10 147.659
R1393 VTAIL.n97 VTAIL.t11 147.659
R1394 VTAIL.n261 VTAIL.t13 147.659
R1395 VTAIL.n219 VTAIL.t12 147.659
R1396 VTAIL.n179 VTAIL.t4 147.659
R1397 VTAIL.n137 VTAIL.t5 147.659
R1398 VTAIL.n305 VTAIL.n299 104.615
R1399 VTAIL.n306 VTAIL.n305 104.615
R1400 VTAIL.n306 VTAIL.n295 104.615
R1401 VTAIL.n313 VTAIL.n295 104.615
R1402 VTAIL.n314 VTAIL.n313 104.615
R1403 VTAIL.n314 VTAIL.n291 104.615
R1404 VTAIL.n321 VTAIL.n291 104.615
R1405 VTAIL.n322 VTAIL.n321 104.615
R1406 VTAIL.n19 VTAIL.n13 104.615
R1407 VTAIL.n20 VTAIL.n19 104.615
R1408 VTAIL.n20 VTAIL.n9 104.615
R1409 VTAIL.n27 VTAIL.n9 104.615
R1410 VTAIL.n28 VTAIL.n27 104.615
R1411 VTAIL.n28 VTAIL.n5 104.615
R1412 VTAIL.n35 VTAIL.n5 104.615
R1413 VTAIL.n36 VTAIL.n35 104.615
R1414 VTAIL.n59 VTAIL.n53 104.615
R1415 VTAIL.n60 VTAIL.n59 104.615
R1416 VTAIL.n60 VTAIL.n49 104.615
R1417 VTAIL.n67 VTAIL.n49 104.615
R1418 VTAIL.n68 VTAIL.n67 104.615
R1419 VTAIL.n68 VTAIL.n45 104.615
R1420 VTAIL.n75 VTAIL.n45 104.615
R1421 VTAIL.n76 VTAIL.n75 104.615
R1422 VTAIL.n101 VTAIL.n95 104.615
R1423 VTAIL.n102 VTAIL.n101 104.615
R1424 VTAIL.n102 VTAIL.n91 104.615
R1425 VTAIL.n109 VTAIL.n91 104.615
R1426 VTAIL.n110 VTAIL.n109 104.615
R1427 VTAIL.n110 VTAIL.n87 104.615
R1428 VTAIL.n117 VTAIL.n87 104.615
R1429 VTAIL.n118 VTAIL.n117 104.615
R1430 VTAIL.n282 VTAIL.n281 104.615
R1431 VTAIL.n281 VTAIL.n251 104.615
R1432 VTAIL.n274 VTAIL.n251 104.615
R1433 VTAIL.n274 VTAIL.n273 104.615
R1434 VTAIL.n273 VTAIL.n255 104.615
R1435 VTAIL.n266 VTAIL.n255 104.615
R1436 VTAIL.n266 VTAIL.n265 104.615
R1437 VTAIL.n265 VTAIL.n259 104.615
R1438 VTAIL.n240 VTAIL.n239 104.615
R1439 VTAIL.n239 VTAIL.n209 104.615
R1440 VTAIL.n232 VTAIL.n209 104.615
R1441 VTAIL.n232 VTAIL.n231 104.615
R1442 VTAIL.n231 VTAIL.n213 104.615
R1443 VTAIL.n224 VTAIL.n213 104.615
R1444 VTAIL.n224 VTAIL.n223 104.615
R1445 VTAIL.n223 VTAIL.n217 104.615
R1446 VTAIL.n200 VTAIL.n199 104.615
R1447 VTAIL.n199 VTAIL.n169 104.615
R1448 VTAIL.n192 VTAIL.n169 104.615
R1449 VTAIL.n192 VTAIL.n191 104.615
R1450 VTAIL.n191 VTAIL.n173 104.615
R1451 VTAIL.n184 VTAIL.n173 104.615
R1452 VTAIL.n184 VTAIL.n183 104.615
R1453 VTAIL.n183 VTAIL.n177 104.615
R1454 VTAIL.n158 VTAIL.n157 104.615
R1455 VTAIL.n157 VTAIL.n127 104.615
R1456 VTAIL.n150 VTAIL.n127 104.615
R1457 VTAIL.n150 VTAIL.n149 104.615
R1458 VTAIL.n149 VTAIL.n131 104.615
R1459 VTAIL.n142 VTAIL.n131 104.615
R1460 VTAIL.n142 VTAIL.n141 104.615
R1461 VTAIL.n141 VTAIL.n135 104.615
R1462 VTAIL.t2 VTAIL.n299 52.3082
R1463 VTAIL.t6 VTAIL.n13 52.3082
R1464 VTAIL.t10 VTAIL.n53 52.3082
R1465 VTAIL.t11 VTAIL.n95 52.3082
R1466 VTAIL.t13 VTAIL.n259 52.3082
R1467 VTAIL.t12 VTAIL.n217 52.3082
R1468 VTAIL.t4 VTAIL.n177 52.3082
R1469 VTAIL.t5 VTAIL.n135 52.3082
R1470 VTAIL.n247 VTAIL.n246 49.1035
R1471 VTAIL.n165 VTAIL.n164 49.1035
R1472 VTAIL.n1 VTAIL.n0 49.1034
R1473 VTAIL.n83 VTAIL.n82 49.1034
R1474 VTAIL.n327 VTAIL.n326 32.7672
R1475 VTAIL.n41 VTAIL.n40 32.7672
R1476 VTAIL.n81 VTAIL.n80 32.7672
R1477 VTAIL.n123 VTAIL.n122 32.7672
R1478 VTAIL.n287 VTAIL.n286 32.7672
R1479 VTAIL.n245 VTAIL.n244 32.7672
R1480 VTAIL.n205 VTAIL.n204 32.7672
R1481 VTAIL.n163 VTAIL.n162 32.7672
R1482 VTAIL.n327 VTAIL.n287 20.4617
R1483 VTAIL.n163 VTAIL.n123 20.4617
R1484 VTAIL.n301 VTAIL.n300 15.6677
R1485 VTAIL.n15 VTAIL.n14 15.6677
R1486 VTAIL.n55 VTAIL.n54 15.6677
R1487 VTAIL.n97 VTAIL.n96 15.6677
R1488 VTAIL.n261 VTAIL.n260 15.6677
R1489 VTAIL.n219 VTAIL.n218 15.6677
R1490 VTAIL.n179 VTAIL.n178 15.6677
R1491 VTAIL.n137 VTAIL.n136 15.6677
R1492 VTAIL.n304 VTAIL.n303 12.8005
R1493 VTAIL.n18 VTAIL.n17 12.8005
R1494 VTAIL.n58 VTAIL.n57 12.8005
R1495 VTAIL.n100 VTAIL.n99 12.8005
R1496 VTAIL.n264 VTAIL.n263 12.8005
R1497 VTAIL.n222 VTAIL.n221 12.8005
R1498 VTAIL.n182 VTAIL.n181 12.8005
R1499 VTAIL.n140 VTAIL.n139 12.8005
R1500 VTAIL.n307 VTAIL.n298 12.0247
R1501 VTAIL.n21 VTAIL.n12 12.0247
R1502 VTAIL.n61 VTAIL.n52 12.0247
R1503 VTAIL.n103 VTAIL.n94 12.0247
R1504 VTAIL.n267 VTAIL.n258 12.0247
R1505 VTAIL.n225 VTAIL.n216 12.0247
R1506 VTAIL.n185 VTAIL.n176 12.0247
R1507 VTAIL.n143 VTAIL.n134 12.0247
R1508 VTAIL.n308 VTAIL.n296 11.249
R1509 VTAIL.n22 VTAIL.n10 11.249
R1510 VTAIL.n62 VTAIL.n50 11.249
R1511 VTAIL.n104 VTAIL.n92 11.249
R1512 VTAIL.n268 VTAIL.n256 11.249
R1513 VTAIL.n226 VTAIL.n214 11.249
R1514 VTAIL.n186 VTAIL.n174 11.249
R1515 VTAIL.n144 VTAIL.n132 11.249
R1516 VTAIL.n312 VTAIL.n311 10.4732
R1517 VTAIL.n26 VTAIL.n25 10.4732
R1518 VTAIL.n66 VTAIL.n65 10.4732
R1519 VTAIL.n108 VTAIL.n107 10.4732
R1520 VTAIL.n272 VTAIL.n271 10.4732
R1521 VTAIL.n230 VTAIL.n229 10.4732
R1522 VTAIL.n190 VTAIL.n189 10.4732
R1523 VTAIL.n148 VTAIL.n147 10.4732
R1524 VTAIL.n315 VTAIL.n294 9.69747
R1525 VTAIL.n29 VTAIL.n8 9.69747
R1526 VTAIL.n69 VTAIL.n48 9.69747
R1527 VTAIL.n111 VTAIL.n90 9.69747
R1528 VTAIL.n275 VTAIL.n254 9.69747
R1529 VTAIL.n233 VTAIL.n212 9.69747
R1530 VTAIL.n193 VTAIL.n172 9.69747
R1531 VTAIL.n151 VTAIL.n130 9.69747
R1532 VTAIL.n326 VTAIL.n325 9.45567
R1533 VTAIL.n40 VTAIL.n39 9.45567
R1534 VTAIL.n80 VTAIL.n79 9.45567
R1535 VTAIL.n122 VTAIL.n121 9.45567
R1536 VTAIL.n286 VTAIL.n285 9.45567
R1537 VTAIL.n244 VTAIL.n243 9.45567
R1538 VTAIL.n204 VTAIL.n203 9.45567
R1539 VTAIL.n162 VTAIL.n161 9.45567
R1540 VTAIL.n325 VTAIL.n324 9.3005
R1541 VTAIL.n319 VTAIL.n318 9.3005
R1542 VTAIL.n317 VTAIL.n316 9.3005
R1543 VTAIL.n294 VTAIL.n293 9.3005
R1544 VTAIL.n311 VTAIL.n310 9.3005
R1545 VTAIL.n309 VTAIL.n308 9.3005
R1546 VTAIL.n298 VTAIL.n297 9.3005
R1547 VTAIL.n303 VTAIL.n302 9.3005
R1548 VTAIL.n290 VTAIL.n289 9.3005
R1549 VTAIL.n39 VTAIL.n38 9.3005
R1550 VTAIL.n33 VTAIL.n32 9.3005
R1551 VTAIL.n31 VTAIL.n30 9.3005
R1552 VTAIL.n8 VTAIL.n7 9.3005
R1553 VTAIL.n25 VTAIL.n24 9.3005
R1554 VTAIL.n23 VTAIL.n22 9.3005
R1555 VTAIL.n12 VTAIL.n11 9.3005
R1556 VTAIL.n17 VTAIL.n16 9.3005
R1557 VTAIL.n4 VTAIL.n3 9.3005
R1558 VTAIL.n79 VTAIL.n78 9.3005
R1559 VTAIL.n73 VTAIL.n72 9.3005
R1560 VTAIL.n71 VTAIL.n70 9.3005
R1561 VTAIL.n48 VTAIL.n47 9.3005
R1562 VTAIL.n65 VTAIL.n64 9.3005
R1563 VTAIL.n63 VTAIL.n62 9.3005
R1564 VTAIL.n52 VTAIL.n51 9.3005
R1565 VTAIL.n57 VTAIL.n56 9.3005
R1566 VTAIL.n44 VTAIL.n43 9.3005
R1567 VTAIL.n121 VTAIL.n120 9.3005
R1568 VTAIL.n115 VTAIL.n114 9.3005
R1569 VTAIL.n113 VTAIL.n112 9.3005
R1570 VTAIL.n90 VTAIL.n89 9.3005
R1571 VTAIL.n107 VTAIL.n106 9.3005
R1572 VTAIL.n105 VTAIL.n104 9.3005
R1573 VTAIL.n94 VTAIL.n93 9.3005
R1574 VTAIL.n99 VTAIL.n98 9.3005
R1575 VTAIL.n86 VTAIL.n85 9.3005
R1576 VTAIL.n285 VTAIL.n284 9.3005
R1577 VTAIL.n250 VTAIL.n249 9.3005
R1578 VTAIL.n279 VTAIL.n278 9.3005
R1579 VTAIL.n277 VTAIL.n276 9.3005
R1580 VTAIL.n254 VTAIL.n253 9.3005
R1581 VTAIL.n271 VTAIL.n270 9.3005
R1582 VTAIL.n269 VTAIL.n268 9.3005
R1583 VTAIL.n258 VTAIL.n257 9.3005
R1584 VTAIL.n263 VTAIL.n262 9.3005
R1585 VTAIL.n243 VTAIL.n242 9.3005
R1586 VTAIL.n208 VTAIL.n207 9.3005
R1587 VTAIL.n237 VTAIL.n236 9.3005
R1588 VTAIL.n235 VTAIL.n234 9.3005
R1589 VTAIL.n212 VTAIL.n211 9.3005
R1590 VTAIL.n229 VTAIL.n228 9.3005
R1591 VTAIL.n227 VTAIL.n226 9.3005
R1592 VTAIL.n216 VTAIL.n215 9.3005
R1593 VTAIL.n221 VTAIL.n220 9.3005
R1594 VTAIL.n203 VTAIL.n202 9.3005
R1595 VTAIL.n168 VTAIL.n167 9.3005
R1596 VTAIL.n197 VTAIL.n196 9.3005
R1597 VTAIL.n195 VTAIL.n194 9.3005
R1598 VTAIL.n172 VTAIL.n171 9.3005
R1599 VTAIL.n189 VTAIL.n188 9.3005
R1600 VTAIL.n187 VTAIL.n186 9.3005
R1601 VTAIL.n176 VTAIL.n175 9.3005
R1602 VTAIL.n181 VTAIL.n180 9.3005
R1603 VTAIL.n161 VTAIL.n160 9.3005
R1604 VTAIL.n126 VTAIL.n125 9.3005
R1605 VTAIL.n155 VTAIL.n154 9.3005
R1606 VTAIL.n153 VTAIL.n152 9.3005
R1607 VTAIL.n130 VTAIL.n129 9.3005
R1608 VTAIL.n147 VTAIL.n146 9.3005
R1609 VTAIL.n145 VTAIL.n144 9.3005
R1610 VTAIL.n134 VTAIL.n133 9.3005
R1611 VTAIL.n139 VTAIL.n138 9.3005
R1612 VTAIL.n316 VTAIL.n292 8.92171
R1613 VTAIL.n30 VTAIL.n6 8.92171
R1614 VTAIL.n70 VTAIL.n46 8.92171
R1615 VTAIL.n112 VTAIL.n88 8.92171
R1616 VTAIL.n276 VTAIL.n252 8.92171
R1617 VTAIL.n234 VTAIL.n210 8.92171
R1618 VTAIL.n194 VTAIL.n170 8.92171
R1619 VTAIL.n152 VTAIL.n128 8.92171
R1620 VTAIL.n320 VTAIL.n319 8.14595
R1621 VTAIL.n34 VTAIL.n33 8.14595
R1622 VTAIL.n74 VTAIL.n73 8.14595
R1623 VTAIL.n116 VTAIL.n115 8.14595
R1624 VTAIL.n280 VTAIL.n279 8.14595
R1625 VTAIL.n238 VTAIL.n237 8.14595
R1626 VTAIL.n198 VTAIL.n197 8.14595
R1627 VTAIL.n156 VTAIL.n155 8.14595
R1628 VTAIL.n323 VTAIL.n290 7.3702
R1629 VTAIL.n326 VTAIL.n288 7.3702
R1630 VTAIL.n37 VTAIL.n4 7.3702
R1631 VTAIL.n40 VTAIL.n2 7.3702
R1632 VTAIL.n77 VTAIL.n44 7.3702
R1633 VTAIL.n80 VTAIL.n42 7.3702
R1634 VTAIL.n119 VTAIL.n86 7.3702
R1635 VTAIL.n122 VTAIL.n84 7.3702
R1636 VTAIL.n286 VTAIL.n248 7.3702
R1637 VTAIL.n283 VTAIL.n250 7.3702
R1638 VTAIL.n244 VTAIL.n206 7.3702
R1639 VTAIL.n241 VTAIL.n208 7.3702
R1640 VTAIL.n204 VTAIL.n166 7.3702
R1641 VTAIL.n201 VTAIL.n168 7.3702
R1642 VTAIL.n162 VTAIL.n124 7.3702
R1643 VTAIL.n159 VTAIL.n126 7.3702
R1644 VTAIL.n324 VTAIL.n323 6.59444
R1645 VTAIL.n324 VTAIL.n288 6.59444
R1646 VTAIL.n38 VTAIL.n37 6.59444
R1647 VTAIL.n38 VTAIL.n2 6.59444
R1648 VTAIL.n78 VTAIL.n77 6.59444
R1649 VTAIL.n78 VTAIL.n42 6.59444
R1650 VTAIL.n120 VTAIL.n119 6.59444
R1651 VTAIL.n120 VTAIL.n84 6.59444
R1652 VTAIL.n284 VTAIL.n248 6.59444
R1653 VTAIL.n284 VTAIL.n283 6.59444
R1654 VTAIL.n242 VTAIL.n206 6.59444
R1655 VTAIL.n242 VTAIL.n241 6.59444
R1656 VTAIL.n202 VTAIL.n166 6.59444
R1657 VTAIL.n202 VTAIL.n201 6.59444
R1658 VTAIL.n160 VTAIL.n124 6.59444
R1659 VTAIL.n160 VTAIL.n159 6.59444
R1660 VTAIL.n320 VTAIL.n290 5.81868
R1661 VTAIL.n34 VTAIL.n4 5.81868
R1662 VTAIL.n74 VTAIL.n44 5.81868
R1663 VTAIL.n116 VTAIL.n86 5.81868
R1664 VTAIL.n280 VTAIL.n250 5.81868
R1665 VTAIL.n238 VTAIL.n208 5.81868
R1666 VTAIL.n198 VTAIL.n168 5.81868
R1667 VTAIL.n156 VTAIL.n126 5.81868
R1668 VTAIL.n319 VTAIL.n292 5.04292
R1669 VTAIL.n33 VTAIL.n6 5.04292
R1670 VTAIL.n73 VTAIL.n46 5.04292
R1671 VTAIL.n115 VTAIL.n88 5.04292
R1672 VTAIL.n279 VTAIL.n252 5.04292
R1673 VTAIL.n237 VTAIL.n210 5.04292
R1674 VTAIL.n197 VTAIL.n170 5.04292
R1675 VTAIL.n155 VTAIL.n128 5.04292
R1676 VTAIL.n262 VTAIL.n261 4.38565
R1677 VTAIL.n220 VTAIL.n219 4.38565
R1678 VTAIL.n180 VTAIL.n179 4.38565
R1679 VTAIL.n138 VTAIL.n137 4.38565
R1680 VTAIL.n302 VTAIL.n301 4.38565
R1681 VTAIL.n16 VTAIL.n15 4.38565
R1682 VTAIL.n56 VTAIL.n55 4.38565
R1683 VTAIL.n98 VTAIL.n97 4.38565
R1684 VTAIL.n316 VTAIL.n315 4.26717
R1685 VTAIL.n30 VTAIL.n29 4.26717
R1686 VTAIL.n70 VTAIL.n69 4.26717
R1687 VTAIL.n112 VTAIL.n111 4.26717
R1688 VTAIL.n276 VTAIL.n275 4.26717
R1689 VTAIL.n234 VTAIL.n233 4.26717
R1690 VTAIL.n194 VTAIL.n193 4.26717
R1691 VTAIL.n152 VTAIL.n151 4.26717
R1692 VTAIL.n312 VTAIL.n294 3.49141
R1693 VTAIL.n26 VTAIL.n8 3.49141
R1694 VTAIL.n66 VTAIL.n48 3.49141
R1695 VTAIL.n108 VTAIL.n90 3.49141
R1696 VTAIL.n272 VTAIL.n254 3.49141
R1697 VTAIL.n230 VTAIL.n212 3.49141
R1698 VTAIL.n190 VTAIL.n172 3.49141
R1699 VTAIL.n148 VTAIL.n130 3.49141
R1700 VTAIL.n311 VTAIL.n296 2.71565
R1701 VTAIL.n25 VTAIL.n10 2.71565
R1702 VTAIL.n65 VTAIL.n50 2.71565
R1703 VTAIL.n107 VTAIL.n92 2.71565
R1704 VTAIL.n271 VTAIL.n256 2.71565
R1705 VTAIL.n229 VTAIL.n214 2.71565
R1706 VTAIL.n189 VTAIL.n174 2.71565
R1707 VTAIL.n147 VTAIL.n132 2.71565
R1708 VTAIL.n0 VTAIL.t7 2.6511
R1709 VTAIL.n0 VTAIL.t0 2.6511
R1710 VTAIL.n82 VTAIL.t15 2.6511
R1711 VTAIL.n82 VTAIL.t8 2.6511
R1712 VTAIL.n246 VTAIL.t9 2.6511
R1713 VTAIL.n246 VTAIL.t14 2.6511
R1714 VTAIL.n164 VTAIL.t1 2.6511
R1715 VTAIL.n164 VTAIL.t3 2.6511
R1716 VTAIL.n308 VTAIL.n307 1.93989
R1717 VTAIL.n22 VTAIL.n21 1.93989
R1718 VTAIL.n62 VTAIL.n61 1.93989
R1719 VTAIL.n104 VTAIL.n103 1.93989
R1720 VTAIL.n268 VTAIL.n267 1.93989
R1721 VTAIL.n226 VTAIL.n225 1.93989
R1722 VTAIL.n186 VTAIL.n185 1.93989
R1723 VTAIL.n144 VTAIL.n143 1.93989
R1724 VTAIL.n165 VTAIL.n163 1.65567
R1725 VTAIL.n205 VTAIL.n165 1.65567
R1726 VTAIL.n247 VTAIL.n245 1.65567
R1727 VTAIL.n287 VTAIL.n247 1.65567
R1728 VTAIL.n123 VTAIL.n83 1.65567
R1729 VTAIL.n83 VTAIL.n81 1.65567
R1730 VTAIL.n41 VTAIL.n1 1.65567
R1731 VTAIL VTAIL.n327 1.59748
R1732 VTAIL.n304 VTAIL.n298 1.16414
R1733 VTAIL.n18 VTAIL.n12 1.16414
R1734 VTAIL.n58 VTAIL.n52 1.16414
R1735 VTAIL.n100 VTAIL.n94 1.16414
R1736 VTAIL.n264 VTAIL.n258 1.16414
R1737 VTAIL.n222 VTAIL.n216 1.16414
R1738 VTAIL.n182 VTAIL.n176 1.16414
R1739 VTAIL.n140 VTAIL.n134 1.16414
R1740 VTAIL.n245 VTAIL.n205 0.470328
R1741 VTAIL.n81 VTAIL.n41 0.470328
R1742 VTAIL.n303 VTAIL.n300 0.388379
R1743 VTAIL.n17 VTAIL.n14 0.388379
R1744 VTAIL.n57 VTAIL.n54 0.388379
R1745 VTAIL.n99 VTAIL.n96 0.388379
R1746 VTAIL.n263 VTAIL.n260 0.388379
R1747 VTAIL.n221 VTAIL.n218 0.388379
R1748 VTAIL.n181 VTAIL.n178 0.388379
R1749 VTAIL.n139 VTAIL.n136 0.388379
R1750 VTAIL.n302 VTAIL.n297 0.155672
R1751 VTAIL.n309 VTAIL.n297 0.155672
R1752 VTAIL.n310 VTAIL.n309 0.155672
R1753 VTAIL.n310 VTAIL.n293 0.155672
R1754 VTAIL.n317 VTAIL.n293 0.155672
R1755 VTAIL.n318 VTAIL.n317 0.155672
R1756 VTAIL.n318 VTAIL.n289 0.155672
R1757 VTAIL.n325 VTAIL.n289 0.155672
R1758 VTAIL.n16 VTAIL.n11 0.155672
R1759 VTAIL.n23 VTAIL.n11 0.155672
R1760 VTAIL.n24 VTAIL.n23 0.155672
R1761 VTAIL.n24 VTAIL.n7 0.155672
R1762 VTAIL.n31 VTAIL.n7 0.155672
R1763 VTAIL.n32 VTAIL.n31 0.155672
R1764 VTAIL.n32 VTAIL.n3 0.155672
R1765 VTAIL.n39 VTAIL.n3 0.155672
R1766 VTAIL.n56 VTAIL.n51 0.155672
R1767 VTAIL.n63 VTAIL.n51 0.155672
R1768 VTAIL.n64 VTAIL.n63 0.155672
R1769 VTAIL.n64 VTAIL.n47 0.155672
R1770 VTAIL.n71 VTAIL.n47 0.155672
R1771 VTAIL.n72 VTAIL.n71 0.155672
R1772 VTAIL.n72 VTAIL.n43 0.155672
R1773 VTAIL.n79 VTAIL.n43 0.155672
R1774 VTAIL.n98 VTAIL.n93 0.155672
R1775 VTAIL.n105 VTAIL.n93 0.155672
R1776 VTAIL.n106 VTAIL.n105 0.155672
R1777 VTAIL.n106 VTAIL.n89 0.155672
R1778 VTAIL.n113 VTAIL.n89 0.155672
R1779 VTAIL.n114 VTAIL.n113 0.155672
R1780 VTAIL.n114 VTAIL.n85 0.155672
R1781 VTAIL.n121 VTAIL.n85 0.155672
R1782 VTAIL.n285 VTAIL.n249 0.155672
R1783 VTAIL.n278 VTAIL.n249 0.155672
R1784 VTAIL.n278 VTAIL.n277 0.155672
R1785 VTAIL.n277 VTAIL.n253 0.155672
R1786 VTAIL.n270 VTAIL.n253 0.155672
R1787 VTAIL.n270 VTAIL.n269 0.155672
R1788 VTAIL.n269 VTAIL.n257 0.155672
R1789 VTAIL.n262 VTAIL.n257 0.155672
R1790 VTAIL.n243 VTAIL.n207 0.155672
R1791 VTAIL.n236 VTAIL.n207 0.155672
R1792 VTAIL.n236 VTAIL.n235 0.155672
R1793 VTAIL.n235 VTAIL.n211 0.155672
R1794 VTAIL.n228 VTAIL.n211 0.155672
R1795 VTAIL.n228 VTAIL.n227 0.155672
R1796 VTAIL.n227 VTAIL.n215 0.155672
R1797 VTAIL.n220 VTAIL.n215 0.155672
R1798 VTAIL.n203 VTAIL.n167 0.155672
R1799 VTAIL.n196 VTAIL.n167 0.155672
R1800 VTAIL.n196 VTAIL.n195 0.155672
R1801 VTAIL.n195 VTAIL.n171 0.155672
R1802 VTAIL.n188 VTAIL.n171 0.155672
R1803 VTAIL.n188 VTAIL.n187 0.155672
R1804 VTAIL.n187 VTAIL.n175 0.155672
R1805 VTAIL.n180 VTAIL.n175 0.155672
R1806 VTAIL.n161 VTAIL.n125 0.155672
R1807 VTAIL.n154 VTAIL.n125 0.155672
R1808 VTAIL.n154 VTAIL.n153 0.155672
R1809 VTAIL.n153 VTAIL.n129 0.155672
R1810 VTAIL.n146 VTAIL.n129 0.155672
R1811 VTAIL.n146 VTAIL.n145 0.155672
R1812 VTAIL.n145 VTAIL.n133 0.155672
R1813 VTAIL.n138 VTAIL.n133 0.155672
R1814 VTAIL VTAIL.n1 0.0586897
R1815 VDD1 VDD1.n0 66.6681
R1816 VDD1.n3 VDD1.n2 66.5544
R1817 VDD1.n3 VDD1.n1 66.5544
R1818 VDD1.n5 VDD1.n4 65.7822
R1819 VDD1.n5 VDD1.n3 38.1862
R1820 VDD1.n4 VDD1.t2 2.6511
R1821 VDD1.n4 VDD1.t3 2.6511
R1822 VDD1.n0 VDD1.t0 2.6511
R1823 VDD1.n0 VDD1.t1 2.6511
R1824 VDD1.n2 VDD1.t6 2.6511
R1825 VDD1.n2 VDD1.t5 2.6511
R1826 VDD1.n1 VDD1.t4 2.6511
R1827 VDD1.n1 VDD1.t7 2.6511
R1828 VDD1 VDD1.n5 0.769897
R1829 VN.n20 VN.n19 179.406
R1830 VN.n41 VN.n40 179.406
R1831 VN.n39 VN.n21 161.3
R1832 VN.n38 VN.n37 161.3
R1833 VN.n36 VN.n22 161.3
R1834 VN.n35 VN.n34 161.3
R1835 VN.n32 VN.n23 161.3
R1836 VN.n31 VN.n30 161.3
R1837 VN.n29 VN.n24 161.3
R1838 VN.n28 VN.n27 161.3
R1839 VN.n18 VN.n0 161.3
R1840 VN.n17 VN.n16 161.3
R1841 VN.n15 VN.n1 161.3
R1842 VN.n14 VN.n13 161.3
R1843 VN.n11 VN.n2 161.3
R1844 VN.n10 VN.n9 161.3
R1845 VN.n8 VN.n3 161.3
R1846 VN.n7 VN.n6 161.3
R1847 VN.n4 VN.t7 145.01
R1848 VN.n25 VN.t4 145.01
R1849 VN.n5 VN.t3 113.225
R1850 VN.n12 VN.t2 113.225
R1851 VN.n19 VN.t0 113.225
R1852 VN.n26 VN.t6 113.225
R1853 VN.n33 VN.t5 113.225
R1854 VN.n40 VN.t1 113.225
R1855 VN.n17 VN.n1 56.5193
R1856 VN.n38 VN.n22 56.5193
R1857 VN.n10 VN.n3 56.5193
R1858 VN.n31 VN.n24 56.5193
R1859 VN.n5 VN.n4 55.7366
R1860 VN.n26 VN.n25 55.7366
R1861 VN VN.n41 43.01
R1862 VN.n6 VN.n3 24.4675
R1863 VN.n11 VN.n10 24.4675
R1864 VN.n13 VN.n1 24.4675
R1865 VN.n18 VN.n17 24.4675
R1866 VN.n27 VN.n24 24.4675
R1867 VN.n34 VN.n22 24.4675
R1868 VN.n32 VN.n31 24.4675
R1869 VN.n39 VN.n38 24.4675
R1870 VN.n28 VN.n25 18.144
R1871 VN.n7 VN.n4 18.144
R1872 VN.n13 VN.n12 14.1914
R1873 VN.n34 VN.n33 14.1914
R1874 VN.n6 VN.n5 10.2766
R1875 VN.n12 VN.n11 10.2766
R1876 VN.n27 VN.n26 10.2766
R1877 VN.n33 VN.n32 10.2766
R1878 VN.n19 VN.n18 6.36192
R1879 VN.n40 VN.n39 6.36192
R1880 VN.n41 VN.n21 0.189894
R1881 VN.n37 VN.n21 0.189894
R1882 VN.n37 VN.n36 0.189894
R1883 VN.n36 VN.n35 0.189894
R1884 VN.n35 VN.n23 0.189894
R1885 VN.n30 VN.n23 0.189894
R1886 VN.n30 VN.n29 0.189894
R1887 VN.n29 VN.n28 0.189894
R1888 VN.n8 VN.n7 0.189894
R1889 VN.n9 VN.n8 0.189894
R1890 VN.n9 VN.n2 0.189894
R1891 VN.n14 VN.n2 0.189894
R1892 VN.n15 VN.n14 0.189894
R1893 VN.n16 VN.n15 0.189894
R1894 VN.n16 VN.n0 0.189894
R1895 VN.n20 VN.n0 0.189894
R1896 VN VN.n20 0.0516364
R1897 VDD2.n2 VDD2.n1 66.5544
R1898 VDD2.n2 VDD2.n0 66.5544
R1899 VDD2 VDD2.n5 66.5516
R1900 VDD2.n4 VDD2.n3 65.7823
R1901 VDD2.n4 VDD2.n2 37.6032
R1902 VDD2.n5 VDD2.t1 2.6511
R1903 VDD2.n5 VDD2.t3 2.6511
R1904 VDD2.n3 VDD2.t6 2.6511
R1905 VDD2.n3 VDD2.t2 2.6511
R1906 VDD2.n1 VDD2.t5 2.6511
R1907 VDD2.n1 VDD2.t7 2.6511
R1908 VDD2.n0 VDD2.t0 2.6511
R1909 VDD2.n0 VDD2.t4 2.6511
R1910 VDD2 VDD2.n4 0.886276
C0 VN VP 5.58923f
C1 VDD1 VN 0.149974f
C2 VDD2 VP 0.412268f
C3 VTAIL VN 5.20096f
C4 VDD1 VDD2 1.2552f
C5 VTAIL VDD2 6.393f
C6 VDD1 VP 5.20807f
C7 VTAIL VP 5.21506f
C8 VTAIL VDD1 6.34535f
C9 VN VDD2 4.94666f
C10 VDD2 B 4.02685f
C11 VDD1 B 4.356495f
C12 VTAIL B 7.080961f
C13 VN B 11.276569f
C14 VP B 9.808548f
C15 VDD2.t0 B 0.14571f
C16 VDD2.t4 B 0.14571f
C17 VDD2.n0 B 1.25004f
C18 VDD2.t5 B 0.14571f
C19 VDD2.t7 B 0.14571f
C20 VDD2.n1 B 1.25004f
C21 VDD2.n2 B 2.38603f
C22 VDD2.t6 B 0.14571f
C23 VDD2.t2 B 0.14571f
C24 VDD2.n3 B 1.24532f
C25 VDD2.n4 B 2.2192f
C26 VDD2.t1 B 0.14571f
C27 VDD2.t3 B 0.14571f
C28 VDD2.n5 B 1.25001f
C29 VN.n0 B 0.031005f
C30 VN.t0 B 0.985962f
C31 VN.n1 B 0.038349f
C32 VN.n2 B 0.031005f
C33 VN.t2 B 0.985962f
C34 VN.n3 B 0.045261f
C35 VN.t7 B 1.09505f
C36 VN.n4 B 0.445003f
C37 VN.t3 B 0.985962f
C38 VN.n5 B 0.430502f
C39 VN.n6 B 0.041238f
C40 VN.n7 B 0.196533f
C41 VN.n8 B 0.031005f
C42 VN.n9 B 0.031005f
C43 VN.n10 B 0.045261f
C44 VN.n11 B 0.041238f
C45 VN.n12 B 0.372533f
C46 VN.n13 B 0.045803f
C47 VN.n14 B 0.031005f
C48 VN.n15 B 0.031005f
C49 VN.n16 B 0.031005f
C50 VN.n17 B 0.052173f
C51 VN.n18 B 0.036674f
C52 VN.n19 B 0.435772f
C53 VN.n20 B 0.031126f
C54 VN.n21 B 0.031005f
C55 VN.t1 B 0.985962f
C56 VN.n22 B 0.038349f
C57 VN.n23 B 0.031005f
C58 VN.t5 B 0.985962f
C59 VN.n24 B 0.045261f
C60 VN.t4 B 1.09505f
C61 VN.n25 B 0.445003f
C62 VN.t6 B 0.985962f
C63 VN.n26 B 0.430502f
C64 VN.n27 B 0.041238f
C65 VN.n28 B 0.196533f
C66 VN.n29 B 0.031005f
C67 VN.n30 B 0.031005f
C68 VN.n31 B 0.045261f
C69 VN.n32 B 0.041238f
C70 VN.n33 B 0.372533f
C71 VN.n34 B 0.045803f
C72 VN.n35 B 0.031005f
C73 VN.n36 B 0.031005f
C74 VN.n37 B 0.031005f
C75 VN.n38 B 0.052173f
C76 VN.n39 B 0.036674f
C77 VN.n40 B 0.435772f
C78 VN.n41 B 1.33916f
C79 VDD1.t0 B 0.147102f
C80 VDD1.t1 B 0.147102f
C81 VDD1.n0 B 1.26279f
C82 VDD1.t4 B 0.147102f
C83 VDD1.t7 B 0.147102f
C84 VDD1.n1 B 1.26198f
C85 VDD1.t6 B 0.147102f
C86 VDD1.t5 B 0.147102f
C87 VDD1.n2 B 1.26198f
C88 VDD1.n3 B 2.46152f
C89 VDD1.t2 B 0.147102f
C90 VDD1.t3 B 0.147102f
C91 VDD1.n4 B 1.25721f
C92 VDD1.n5 B 2.27041f
C93 VTAIL.t7 B 0.122371f
C94 VTAIL.t0 B 0.122371f
C95 VTAIL.n0 B 0.989005f
C96 VTAIL.n1 B 0.314392f
C97 VTAIL.n2 B 0.030677f
C98 VTAIL.n3 B 0.02073f
C99 VTAIL.n4 B 0.011139f
C100 VTAIL.n5 B 0.02633f
C101 VTAIL.n6 B 0.011795f
C102 VTAIL.n7 B 0.02073f
C103 VTAIL.n8 B 0.011139f
C104 VTAIL.n9 B 0.02633f
C105 VTAIL.n10 B 0.011795f
C106 VTAIL.n11 B 0.02073f
C107 VTAIL.n12 B 0.011139f
C108 VTAIL.n13 B 0.019747f
C109 VTAIL.n14 B 0.015554f
C110 VTAIL.t6 B 0.04292f
C111 VTAIL.n15 B 0.096155f
C112 VTAIL.n16 B 0.633208f
C113 VTAIL.n17 B 0.011139f
C114 VTAIL.n18 B 0.011795f
C115 VTAIL.n19 B 0.02633f
C116 VTAIL.n20 B 0.02633f
C117 VTAIL.n21 B 0.011795f
C118 VTAIL.n22 B 0.011139f
C119 VTAIL.n23 B 0.02073f
C120 VTAIL.n24 B 0.02073f
C121 VTAIL.n25 B 0.011139f
C122 VTAIL.n26 B 0.011795f
C123 VTAIL.n27 B 0.02633f
C124 VTAIL.n28 B 0.02633f
C125 VTAIL.n29 B 0.011795f
C126 VTAIL.n30 B 0.011139f
C127 VTAIL.n31 B 0.02073f
C128 VTAIL.n32 B 0.02073f
C129 VTAIL.n33 B 0.011139f
C130 VTAIL.n34 B 0.011795f
C131 VTAIL.n35 B 0.02633f
C132 VTAIL.n36 B 0.05972f
C133 VTAIL.n37 B 0.011795f
C134 VTAIL.n38 B 0.011139f
C135 VTAIL.n39 B 0.048766f
C136 VTAIL.n40 B 0.033721f
C137 VTAIL.n41 B 0.160129f
C138 VTAIL.n42 B 0.030677f
C139 VTAIL.n43 B 0.02073f
C140 VTAIL.n44 B 0.011139f
C141 VTAIL.n45 B 0.02633f
C142 VTAIL.n46 B 0.011795f
C143 VTAIL.n47 B 0.02073f
C144 VTAIL.n48 B 0.011139f
C145 VTAIL.n49 B 0.02633f
C146 VTAIL.n50 B 0.011795f
C147 VTAIL.n51 B 0.02073f
C148 VTAIL.n52 B 0.011139f
C149 VTAIL.n53 B 0.019747f
C150 VTAIL.n54 B 0.015554f
C151 VTAIL.t10 B 0.04292f
C152 VTAIL.n55 B 0.096155f
C153 VTAIL.n56 B 0.633208f
C154 VTAIL.n57 B 0.011139f
C155 VTAIL.n58 B 0.011795f
C156 VTAIL.n59 B 0.02633f
C157 VTAIL.n60 B 0.02633f
C158 VTAIL.n61 B 0.011795f
C159 VTAIL.n62 B 0.011139f
C160 VTAIL.n63 B 0.02073f
C161 VTAIL.n64 B 0.02073f
C162 VTAIL.n65 B 0.011139f
C163 VTAIL.n66 B 0.011795f
C164 VTAIL.n67 B 0.02633f
C165 VTAIL.n68 B 0.02633f
C166 VTAIL.n69 B 0.011795f
C167 VTAIL.n70 B 0.011139f
C168 VTAIL.n71 B 0.02073f
C169 VTAIL.n72 B 0.02073f
C170 VTAIL.n73 B 0.011139f
C171 VTAIL.n74 B 0.011795f
C172 VTAIL.n75 B 0.02633f
C173 VTAIL.n76 B 0.05972f
C174 VTAIL.n77 B 0.011795f
C175 VTAIL.n78 B 0.011139f
C176 VTAIL.n79 B 0.048766f
C177 VTAIL.n80 B 0.033721f
C178 VTAIL.n81 B 0.160129f
C179 VTAIL.t15 B 0.122371f
C180 VTAIL.t8 B 0.122371f
C181 VTAIL.n82 B 0.989005f
C182 VTAIL.n83 B 0.421066f
C183 VTAIL.n84 B 0.030677f
C184 VTAIL.n85 B 0.02073f
C185 VTAIL.n86 B 0.011139f
C186 VTAIL.n87 B 0.02633f
C187 VTAIL.n88 B 0.011795f
C188 VTAIL.n89 B 0.02073f
C189 VTAIL.n90 B 0.011139f
C190 VTAIL.n91 B 0.02633f
C191 VTAIL.n92 B 0.011795f
C192 VTAIL.n93 B 0.02073f
C193 VTAIL.n94 B 0.011139f
C194 VTAIL.n95 B 0.019747f
C195 VTAIL.n96 B 0.015554f
C196 VTAIL.t11 B 0.04292f
C197 VTAIL.n97 B 0.096155f
C198 VTAIL.n98 B 0.633208f
C199 VTAIL.n99 B 0.011139f
C200 VTAIL.n100 B 0.011795f
C201 VTAIL.n101 B 0.02633f
C202 VTAIL.n102 B 0.02633f
C203 VTAIL.n103 B 0.011795f
C204 VTAIL.n104 B 0.011139f
C205 VTAIL.n105 B 0.02073f
C206 VTAIL.n106 B 0.02073f
C207 VTAIL.n107 B 0.011139f
C208 VTAIL.n108 B 0.011795f
C209 VTAIL.n109 B 0.02633f
C210 VTAIL.n110 B 0.02633f
C211 VTAIL.n111 B 0.011795f
C212 VTAIL.n112 B 0.011139f
C213 VTAIL.n113 B 0.02073f
C214 VTAIL.n114 B 0.02073f
C215 VTAIL.n115 B 0.011139f
C216 VTAIL.n116 B 0.011795f
C217 VTAIL.n117 B 0.02633f
C218 VTAIL.n118 B 0.05972f
C219 VTAIL.n119 B 0.011795f
C220 VTAIL.n120 B 0.011139f
C221 VTAIL.n121 B 0.048766f
C222 VTAIL.n122 B 0.033721f
C223 VTAIL.n123 B 0.951054f
C224 VTAIL.n124 B 0.030677f
C225 VTAIL.n125 B 0.02073f
C226 VTAIL.n126 B 0.011139f
C227 VTAIL.n127 B 0.02633f
C228 VTAIL.n128 B 0.011795f
C229 VTAIL.n129 B 0.02073f
C230 VTAIL.n130 B 0.011139f
C231 VTAIL.n131 B 0.02633f
C232 VTAIL.n132 B 0.011795f
C233 VTAIL.n133 B 0.02073f
C234 VTAIL.n134 B 0.011139f
C235 VTAIL.n135 B 0.019747f
C236 VTAIL.n136 B 0.015554f
C237 VTAIL.t5 B 0.04292f
C238 VTAIL.n137 B 0.096155f
C239 VTAIL.n138 B 0.633208f
C240 VTAIL.n139 B 0.011139f
C241 VTAIL.n140 B 0.011795f
C242 VTAIL.n141 B 0.02633f
C243 VTAIL.n142 B 0.02633f
C244 VTAIL.n143 B 0.011795f
C245 VTAIL.n144 B 0.011139f
C246 VTAIL.n145 B 0.02073f
C247 VTAIL.n146 B 0.02073f
C248 VTAIL.n147 B 0.011139f
C249 VTAIL.n148 B 0.011795f
C250 VTAIL.n149 B 0.02633f
C251 VTAIL.n150 B 0.02633f
C252 VTAIL.n151 B 0.011795f
C253 VTAIL.n152 B 0.011139f
C254 VTAIL.n153 B 0.02073f
C255 VTAIL.n154 B 0.02073f
C256 VTAIL.n155 B 0.011139f
C257 VTAIL.n156 B 0.011795f
C258 VTAIL.n157 B 0.02633f
C259 VTAIL.n158 B 0.05972f
C260 VTAIL.n159 B 0.011795f
C261 VTAIL.n160 B 0.011139f
C262 VTAIL.n161 B 0.048766f
C263 VTAIL.n162 B 0.033721f
C264 VTAIL.n163 B 0.951054f
C265 VTAIL.t1 B 0.122371f
C266 VTAIL.t3 B 0.122371f
C267 VTAIL.n164 B 0.989011f
C268 VTAIL.n165 B 0.42106f
C269 VTAIL.n166 B 0.030677f
C270 VTAIL.n167 B 0.02073f
C271 VTAIL.n168 B 0.011139f
C272 VTAIL.n169 B 0.02633f
C273 VTAIL.n170 B 0.011795f
C274 VTAIL.n171 B 0.02073f
C275 VTAIL.n172 B 0.011139f
C276 VTAIL.n173 B 0.02633f
C277 VTAIL.n174 B 0.011795f
C278 VTAIL.n175 B 0.02073f
C279 VTAIL.n176 B 0.011139f
C280 VTAIL.n177 B 0.019747f
C281 VTAIL.n178 B 0.015554f
C282 VTAIL.t4 B 0.04292f
C283 VTAIL.n179 B 0.096155f
C284 VTAIL.n180 B 0.633208f
C285 VTAIL.n181 B 0.011139f
C286 VTAIL.n182 B 0.011795f
C287 VTAIL.n183 B 0.02633f
C288 VTAIL.n184 B 0.02633f
C289 VTAIL.n185 B 0.011795f
C290 VTAIL.n186 B 0.011139f
C291 VTAIL.n187 B 0.02073f
C292 VTAIL.n188 B 0.02073f
C293 VTAIL.n189 B 0.011139f
C294 VTAIL.n190 B 0.011795f
C295 VTAIL.n191 B 0.02633f
C296 VTAIL.n192 B 0.02633f
C297 VTAIL.n193 B 0.011795f
C298 VTAIL.n194 B 0.011139f
C299 VTAIL.n195 B 0.02073f
C300 VTAIL.n196 B 0.02073f
C301 VTAIL.n197 B 0.011139f
C302 VTAIL.n198 B 0.011795f
C303 VTAIL.n199 B 0.02633f
C304 VTAIL.n200 B 0.05972f
C305 VTAIL.n201 B 0.011795f
C306 VTAIL.n202 B 0.011139f
C307 VTAIL.n203 B 0.048766f
C308 VTAIL.n204 B 0.033721f
C309 VTAIL.n205 B 0.160129f
C310 VTAIL.n206 B 0.030677f
C311 VTAIL.n207 B 0.02073f
C312 VTAIL.n208 B 0.011139f
C313 VTAIL.n209 B 0.02633f
C314 VTAIL.n210 B 0.011795f
C315 VTAIL.n211 B 0.02073f
C316 VTAIL.n212 B 0.011139f
C317 VTAIL.n213 B 0.02633f
C318 VTAIL.n214 B 0.011795f
C319 VTAIL.n215 B 0.02073f
C320 VTAIL.n216 B 0.011139f
C321 VTAIL.n217 B 0.019747f
C322 VTAIL.n218 B 0.015554f
C323 VTAIL.t12 B 0.04292f
C324 VTAIL.n219 B 0.096155f
C325 VTAIL.n220 B 0.633208f
C326 VTAIL.n221 B 0.011139f
C327 VTAIL.n222 B 0.011795f
C328 VTAIL.n223 B 0.02633f
C329 VTAIL.n224 B 0.02633f
C330 VTAIL.n225 B 0.011795f
C331 VTAIL.n226 B 0.011139f
C332 VTAIL.n227 B 0.02073f
C333 VTAIL.n228 B 0.02073f
C334 VTAIL.n229 B 0.011139f
C335 VTAIL.n230 B 0.011795f
C336 VTAIL.n231 B 0.02633f
C337 VTAIL.n232 B 0.02633f
C338 VTAIL.n233 B 0.011795f
C339 VTAIL.n234 B 0.011139f
C340 VTAIL.n235 B 0.02073f
C341 VTAIL.n236 B 0.02073f
C342 VTAIL.n237 B 0.011139f
C343 VTAIL.n238 B 0.011795f
C344 VTAIL.n239 B 0.02633f
C345 VTAIL.n240 B 0.05972f
C346 VTAIL.n241 B 0.011795f
C347 VTAIL.n242 B 0.011139f
C348 VTAIL.n243 B 0.048766f
C349 VTAIL.n244 B 0.033721f
C350 VTAIL.n245 B 0.160129f
C351 VTAIL.t9 B 0.122371f
C352 VTAIL.t14 B 0.122371f
C353 VTAIL.n246 B 0.989011f
C354 VTAIL.n247 B 0.42106f
C355 VTAIL.n248 B 0.030677f
C356 VTAIL.n249 B 0.02073f
C357 VTAIL.n250 B 0.011139f
C358 VTAIL.n251 B 0.02633f
C359 VTAIL.n252 B 0.011795f
C360 VTAIL.n253 B 0.02073f
C361 VTAIL.n254 B 0.011139f
C362 VTAIL.n255 B 0.02633f
C363 VTAIL.n256 B 0.011795f
C364 VTAIL.n257 B 0.02073f
C365 VTAIL.n258 B 0.011139f
C366 VTAIL.n259 B 0.019747f
C367 VTAIL.n260 B 0.015554f
C368 VTAIL.t13 B 0.04292f
C369 VTAIL.n261 B 0.096155f
C370 VTAIL.n262 B 0.633208f
C371 VTAIL.n263 B 0.011139f
C372 VTAIL.n264 B 0.011795f
C373 VTAIL.n265 B 0.02633f
C374 VTAIL.n266 B 0.02633f
C375 VTAIL.n267 B 0.011795f
C376 VTAIL.n268 B 0.011139f
C377 VTAIL.n269 B 0.02073f
C378 VTAIL.n270 B 0.02073f
C379 VTAIL.n271 B 0.011139f
C380 VTAIL.n272 B 0.011795f
C381 VTAIL.n273 B 0.02633f
C382 VTAIL.n274 B 0.02633f
C383 VTAIL.n275 B 0.011795f
C384 VTAIL.n276 B 0.011139f
C385 VTAIL.n277 B 0.02073f
C386 VTAIL.n278 B 0.02073f
C387 VTAIL.n279 B 0.011139f
C388 VTAIL.n280 B 0.011795f
C389 VTAIL.n281 B 0.02633f
C390 VTAIL.n282 B 0.05972f
C391 VTAIL.n283 B 0.011795f
C392 VTAIL.n284 B 0.011139f
C393 VTAIL.n285 B 0.048766f
C394 VTAIL.n286 B 0.033721f
C395 VTAIL.n287 B 0.951054f
C396 VTAIL.n288 B 0.030677f
C397 VTAIL.n289 B 0.02073f
C398 VTAIL.n290 B 0.011139f
C399 VTAIL.n291 B 0.02633f
C400 VTAIL.n292 B 0.011795f
C401 VTAIL.n293 B 0.02073f
C402 VTAIL.n294 B 0.011139f
C403 VTAIL.n295 B 0.02633f
C404 VTAIL.n296 B 0.011795f
C405 VTAIL.n297 B 0.02073f
C406 VTAIL.n298 B 0.011139f
C407 VTAIL.n299 B 0.019747f
C408 VTAIL.n300 B 0.015554f
C409 VTAIL.t2 B 0.04292f
C410 VTAIL.n301 B 0.096155f
C411 VTAIL.n302 B 0.633208f
C412 VTAIL.n303 B 0.011139f
C413 VTAIL.n304 B 0.011795f
C414 VTAIL.n305 B 0.02633f
C415 VTAIL.n306 B 0.02633f
C416 VTAIL.n307 B 0.011795f
C417 VTAIL.n308 B 0.011139f
C418 VTAIL.n309 B 0.02073f
C419 VTAIL.n310 B 0.02073f
C420 VTAIL.n311 B 0.011139f
C421 VTAIL.n312 B 0.011795f
C422 VTAIL.n313 B 0.02633f
C423 VTAIL.n314 B 0.02633f
C424 VTAIL.n315 B 0.011795f
C425 VTAIL.n316 B 0.011139f
C426 VTAIL.n317 B 0.02073f
C427 VTAIL.n318 B 0.02073f
C428 VTAIL.n319 B 0.011139f
C429 VTAIL.n320 B 0.011795f
C430 VTAIL.n321 B 0.02633f
C431 VTAIL.n322 B 0.05972f
C432 VTAIL.n323 B 0.011795f
C433 VTAIL.n324 B 0.011139f
C434 VTAIL.n325 B 0.048766f
C435 VTAIL.n326 B 0.033721f
C436 VTAIL.n327 B 0.947167f
C437 VP.n0 B 0.031685f
C438 VP.t2 B 1.0076f
C439 VP.n1 B 0.039191f
C440 VP.n2 B 0.031685f
C441 VP.t1 B 1.0076f
C442 VP.n3 B 0.046255f
C443 VP.n4 B 0.031685f
C444 VP.t0 B 1.0076f
C445 VP.n5 B 0.053318f
C446 VP.n6 B 0.031685f
C447 VP.t4 B 1.0076f
C448 VP.n7 B 0.039191f
C449 VP.n8 B 0.031685f
C450 VP.t5 B 1.0076f
C451 VP.n9 B 0.046255f
C452 VP.t7 B 1.11908f
C453 VP.n10 B 0.454769f
C454 VP.t6 B 1.0076f
C455 VP.n11 B 0.43995f
C456 VP.n12 B 0.042143f
C457 VP.n13 B 0.200846f
C458 VP.n14 B 0.031685f
C459 VP.n15 B 0.031685f
C460 VP.n16 B 0.046255f
C461 VP.n17 B 0.042143f
C462 VP.n18 B 0.380709f
C463 VP.n19 B 0.046808f
C464 VP.n20 B 0.031685f
C465 VP.n21 B 0.031685f
C466 VP.n22 B 0.031685f
C467 VP.n23 B 0.053318f
C468 VP.n24 B 0.037479f
C469 VP.n25 B 0.445336f
C470 VP.n26 B 1.34777f
C471 VP.n27 B 1.37449f
C472 VP.t3 B 1.0076f
C473 VP.n28 B 0.445336f
C474 VP.n29 B 0.037479f
C475 VP.n30 B 0.031685f
C476 VP.n31 B 0.031685f
C477 VP.n32 B 0.031685f
C478 VP.n33 B 0.039191f
C479 VP.n34 B 0.046808f
C480 VP.n35 B 0.380709f
C481 VP.n36 B 0.042143f
C482 VP.n37 B 0.031685f
C483 VP.n38 B 0.031685f
C484 VP.n39 B 0.031685f
C485 VP.n40 B 0.046255f
C486 VP.n41 B 0.042143f
C487 VP.n42 B 0.380709f
C488 VP.n43 B 0.046808f
C489 VP.n44 B 0.031685f
C490 VP.n45 B 0.031685f
C491 VP.n46 B 0.031685f
C492 VP.n47 B 0.053318f
C493 VP.n48 B 0.037479f
C494 VP.n49 B 0.445336f
C495 VP.n50 B 0.031809f
.ends

