* NGSPICE file created from diff_pair_sample_0559.ext - technology: sky130A

.subckt diff_pair_sample_0559 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X1 VDD1.t8 VP.t1 VTAIL.t11 B.t22 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=0.36
X2 VDD2.t9 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=0.36
X3 VDD2.t8 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=0.36
X4 VTAIL.t8 VP.t2 VDD1.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X5 VDD1.t6 VP.t3 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=0.36
X6 VDD2.t7 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=0.36
X7 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=0.36
X8 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=0.36
X9 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X10 VTAIL.t12 VP.t4 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X11 VDD2.t5 VN.t4 VTAIL.t16 B.t20 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X12 VTAIL.t15 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X13 VDD2.t4 VN.t5 VTAIL.t17 B.t22 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=0.36
X14 VTAIL.t13 VP.t6 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X15 VDD2.t3 VN.t6 VTAIL.t18 B.t23 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X16 VDD1.t2 VP.t7 VTAIL.t14 B.t20 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X17 VDD1.t1 VP.t8 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=0.36
X18 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=0.36
X19 VTAIL.t19 VN.t7 VDD2.t2 B.t21 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X20 VTAIL.t1 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
X21 VDD1.t0 VP.t9 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=0.36
X22 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=0.36
X23 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=0.36
R0 VP.n5 VP.t3 820.968
R1 VP.n15 VP.t8 799.986
R2 VP.n16 VP.t2 799.986
R3 VP.n1 VP.t7 799.986
R4 VP.n21 VP.t4 799.986
R5 VP.n22 VP.t1 799.986
R6 VP.n12 VP.t9 799.986
R7 VP.n11 VP.t5 799.986
R8 VP.n4 VP.t0 799.986
R9 VP.n6 VP.t6 799.986
R10 VP.n23 VP.n22 161.3
R11 VP.n8 VP.n7 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n11 VP.n3 161.3
R14 VP.n13 VP.n12 161.3
R15 VP.n21 VP.n0 161.3
R16 VP.n20 VP.n19 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n2 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n8 VP.n5 70.4033
R21 VP.n16 VP.n15 48.2005
R22 VP.n22 VP.n21 48.2005
R23 VP.n12 VP.n11 48.2005
R24 VP.n14 VP.n13 39.6179
R25 VP.n17 VP.n16 37.9763
R26 VP.n21 VP.n20 37.9763
R27 VP.n11 VP.n10 37.9763
R28 VP.n7 VP.n6 37.9763
R29 VP.n6 VP.n5 20.9576
R30 VP.n17 VP.n1 10.2247
R31 VP.n20 VP.n1 10.2247
R32 VP.n10 VP.n4 10.2247
R33 VP.n7 VP.n4 10.2247
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n3 0.189894
R36 VP.n13 VP.n3 0.189894
R37 VP.n14 VP.n2 0.189894
R38 VP.n18 VP.n2 0.189894
R39 VP.n19 VP.n18 0.189894
R40 VP.n19 VP.n0 0.189894
R41 VP.n23 VP.n0 0.189894
R42 VP VP.n23 0.0516364
R43 VTAIL.n11 VTAIL.t17 47.3387
R44 VTAIL.n17 VTAIL.t3 47.3384
R45 VTAIL.n2 VTAIL.t11 47.3384
R46 VTAIL.n16 VTAIL.t7 47.3384
R47 VTAIL.n15 VTAIL.n14 45.4163
R48 VTAIL.n13 VTAIL.n12 45.4163
R49 VTAIL.n10 VTAIL.n9 45.4163
R50 VTAIL.n8 VTAIL.n7 45.4163
R51 VTAIL.n19 VTAIL.n18 45.4161
R52 VTAIL.n1 VTAIL.n0 45.4161
R53 VTAIL.n4 VTAIL.n3 45.4161
R54 VTAIL.n6 VTAIL.n5 45.4161
R55 VTAIL.n8 VTAIL.n6 22.4358
R56 VTAIL.n17 VTAIL.n16 21.841
R57 VTAIL.n18 VTAIL.t18 1.92283
R58 VTAIL.n18 VTAIL.t2 1.92283
R59 VTAIL.n0 VTAIL.t5 1.92283
R60 VTAIL.n0 VTAIL.t1 1.92283
R61 VTAIL.n3 VTAIL.t14 1.92283
R62 VTAIL.n3 VTAIL.t12 1.92283
R63 VTAIL.n5 VTAIL.t10 1.92283
R64 VTAIL.n5 VTAIL.t8 1.92283
R65 VTAIL.n14 VTAIL.t9 1.92283
R66 VTAIL.n14 VTAIL.t15 1.92283
R67 VTAIL.n12 VTAIL.t6 1.92283
R68 VTAIL.n12 VTAIL.t13 1.92283
R69 VTAIL.n9 VTAIL.t16 1.92283
R70 VTAIL.n9 VTAIL.t0 1.92283
R71 VTAIL.n7 VTAIL.t4 1.92283
R72 VTAIL.n7 VTAIL.t19 1.92283
R73 VTAIL.n13 VTAIL.n11 0.767741
R74 VTAIL.n2 VTAIL.n1 0.767741
R75 VTAIL.n10 VTAIL.n8 0.595328
R76 VTAIL.n11 VTAIL.n10 0.595328
R77 VTAIL.n15 VTAIL.n13 0.595328
R78 VTAIL.n16 VTAIL.n15 0.595328
R79 VTAIL.n6 VTAIL.n4 0.595328
R80 VTAIL.n4 VTAIL.n2 0.595328
R81 VTAIL.n19 VTAIL.n17 0.595328
R82 VTAIL VTAIL.n1 0.50481
R83 VTAIL VTAIL.n19 0.0910172
R84 VDD1.n1 VDD1.t6 64.6123
R85 VDD1.n3 VDD1.t1 64.612
R86 VDD1.n5 VDD1.n4 62.4857
R87 VDD1.n1 VDD1.n0 62.0951
R88 VDD1.n7 VDD1.n6 62.0949
R89 VDD1.n3 VDD1.n2 62.0949
R90 VDD1.n7 VDD1.n5 36.3005
R91 VDD1.n6 VDD1.t4 1.92283
R92 VDD1.n6 VDD1.t0 1.92283
R93 VDD1.n0 VDD1.t3 1.92283
R94 VDD1.n0 VDD1.t9 1.92283
R95 VDD1.n4 VDD1.t5 1.92283
R96 VDD1.n4 VDD1.t8 1.92283
R97 VDD1.n2 VDD1.t7 1.92283
R98 VDD1.n2 VDD1.t2 1.92283
R99 VDD1 VDD1.n7 0.388431
R100 VDD1 VDD1.n1 0.207397
R101 VDD1.n5 VDD1.n3 0.0938609
R102 B.n305 B.t17 900.621
R103 B.n311 B.t13 900.621
R104 B.n86 B.t6 900.621
R105 B.n83 B.t10 900.621
R106 B.n588 B.n587 585
R107 B.n589 B.n588 585
R108 B.n249 B.n82 585
R109 B.n248 B.n247 585
R110 B.n246 B.n245 585
R111 B.n244 B.n243 585
R112 B.n242 B.n241 585
R113 B.n240 B.n239 585
R114 B.n238 B.n237 585
R115 B.n236 B.n235 585
R116 B.n234 B.n233 585
R117 B.n232 B.n231 585
R118 B.n230 B.n229 585
R119 B.n228 B.n227 585
R120 B.n226 B.n225 585
R121 B.n224 B.n223 585
R122 B.n222 B.n221 585
R123 B.n220 B.n219 585
R124 B.n218 B.n217 585
R125 B.n216 B.n215 585
R126 B.n214 B.n213 585
R127 B.n212 B.n211 585
R128 B.n210 B.n209 585
R129 B.n208 B.n207 585
R130 B.n206 B.n205 585
R131 B.n204 B.n203 585
R132 B.n202 B.n201 585
R133 B.n200 B.n199 585
R134 B.n198 B.n197 585
R135 B.n196 B.n195 585
R136 B.n194 B.n193 585
R137 B.n192 B.n191 585
R138 B.n190 B.n189 585
R139 B.n188 B.n187 585
R140 B.n186 B.n185 585
R141 B.n184 B.n183 585
R142 B.n182 B.n181 585
R143 B.n180 B.n179 585
R144 B.n178 B.n177 585
R145 B.n176 B.n175 585
R146 B.n174 B.n173 585
R147 B.n172 B.n171 585
R148 B.n170 B.n169 585
R149 B.n168 B.n167 585
R150 B.n166 B.n165 585
R151 B.n164 B.n163 585
R152 B.n162 B.n161 585
R153 B.n159 B.n158 585
R154 B.n157 B.n156 585
R155 B.n155 B.n154 585
R156 B.n153 B.n152 585
R157 B.n151 B.n150 585
R158 B.n149 B.n148 585
R159 B.n147 B.n146 585
R160 B.n145 B.n144 585
R161 B.n143 B.n142 585
R162 B.n141 B.n140 585
R163 B.n139 B.n138 585
R164 B.n137 B.n136 585
R165 B.n135 B.n134 585
R166 B.n133 B.n132 585
R167 B.n131 B.n130 585
R168 B.n129 B.n128 585
R169 B.n127 B.n126 585
R170 B.n125 B.n124 585
R171 B.n123 B.n122 585
R172 B.n121 B.n120 585
R173 B.n119 B.n118 585
R174 B.n117 B.n116 585
R175 B.n115 B.n114 585
R176 B.n113 B.n112 585
R177 B.n111 B.n110 585
R178 B.n109 B.n108 585
R179 B.n107 B.n106 585
R180 B.n105 B.n104 585
R181 B.n103 B.n102 585
R182 B.n101 B.n100 585
R183 B.n99 B.n98 585
R184 B.n97 B.n96 585
R185 B.n95 B.n94 585
R186 B.n93 B.n92 585
R187 B.n91 B.n90 585
R188 B.n89 B.n88 585
R189 B.n39 B.n38 585
R190 B.n586 B.n40 585
R191 B.n590 B.n40 585
R192 B.n585 B.n584 585
R193 B.n584 B.n36 585
R194 B.n583 B.n35 585
R195 B.n596 B.n35 585
R196 B.n582 B.n34 585
R197 B.n597 B.n34 585
R198 B.n581 B.n33 585
R199 B.n598 B.n33 585
R200 B.n580 B.n579 585
R201 B.n579 B.n29 585
R202 B.n578 B.n28 585
R203 B.n604 B.n28 585
R204 B.n577 B.n27 585
R205 B.n605 B.n27 585
R206 B.n576 B.n26 585
R207 B.n606 B.n26 585
R208 B.n575 B.n574 585
R209 B.n574 B.n25 585
R210 B.n573 B.n21 585
R211 B.n612 B.n21 585
R212 B.n572 B.n20 585
R213 B.n613 B.n20 585
R214 B.n571 B.n19 585
R215 B.n614 B.n19 585
R216 B.n570 B.n569 585
R217 B.n569 B.n18 585
R218 B.n568 B.n14 585
R219 B.n620 B.n14 585
R220 B.n567 B.n13 585
R221 B.n621 B.n13 585
R222 B.n566 B.n12 585
R223 B.n622 B.n12 585
R224 B.n565 B.n564 585
R225 B.n564 B.n11 585
R226 B.n563 B.n7 585
R227 B.n628 B.n7 585
R228 B.n562 B.n6 585
R229 B.n629 B.n6 585
R230 B.n561 B.n5 585
R231 B.n630 B.n5 585
R232 B.n560 B.n559 585
R233 B.n559 B.n4 585
R234 B.n558 B.n250 585
R235 B.n558 B.n557 585
R236 B.n547 B.n251 585
R237 B.n550 B.n251 585
R238 B.n549 B.n548 585
R239 B.n551 B.n549 585
R240 B.n546 B.n255 585
R241 B.n258 B.n255 585
R242 B.n545 B.n544 585
R243 B.n544 B.n543 585
R244 B.n257 B.n256 585
R245 B.n536 B.n257 585
R246 B.n535 B.n534 585
R247 B.n537 B.n535 585
R248 B.n533 B.n262 585
R249 B.n265 B.n262 585
R250 B.n532 B.n531 585
R251 B.n531 B.n530 585
R252 B.n264 B.n263 585
R253 B.n523 B.n264 585
R254 B.n522 B.n521 585
R255 B.n524 B.n522 585
R256 B.n520 B.n270 585
R257 B.n270 B.n269 585
R258 B.n519 B.n518 585
R259 B.n518 B.n517 585
R260 B.n272 B.n271 585
R261 B.n273 B.n272 585
R262 B.n510 B.n509 585
R263 B.n511 B.n510 585
R264 B.n508 B.n278 585
R265 B.n278 B.n277 585
R266 B.n507 B.n506 585
R267 B.n506 B.n505 585
R268 B.n280 B.n279 585
R269 B.n281 B.n280 585
R270 B.n498 B.n497 585
R271 B.n499 B.n498 585
R272 B.n284 B.n283 585
R273 B.n334 B.n333 585
R274 B.n335 B.n331 585
R275 B.n331 B.n285 585
R276 B.n337 B.n336 585
R277 B.n339 B.n330 585
R278 B.n342 B.n341 585
R279 B.n343 B.n329 585
R280 B.n345 B.n344 585
R281 B.n347 B.n328 585
R282 B.n350 B.n349 585
R283 B.n351 B.n327 585
R284 B.n353 B.n352 585
R285 B.n355 B.n326 585
R286 B.n358 B.n357 585
R287 B.n359 B.n325 585
R288 B.n361 B.n360 585
R289 B.n363 B.n324 585
R290 B.n366 B.n365 585
R291 B.n367 B.n323 585
R292 B.n369 B.n368 585
R293 B.n371 B.n322 585
R294 B.n374 B.n373 585
R295 B.n375 B.n321 585
R296 B.n377 B.n376 585
R297 B.n379 B.n320 585
R298 B.n382 B.n381 585
R299 B.n383 B.n319 585
R300 B.n385 B.n384 585
R301 B.n387 B.n318 585
R302 B.n390 B.n389 585
R303 B.n391 B.n317 585
R304 B.n393 B.n392 585
R305 B.n395 B.n316 585
R306 B.n398 B.n397 585
R307 B.n399 B.n315 585
R308 B.n401 B.n400 585
R309 B.n403 B.n314 585
R310 B.n406 B.n405 585
R311 B.n407 B.n310 585
R312 B.n409 B.n408 585
R313 B.n411 B.n309 585
R314 B.n414 B.n413 585
R315 B.n415 B.n308 585
R316 B.n417 B.n416 585
R317 B.n419 B.n307 585
R318 B.n422 B.n421 585
R319 B.n424 B.n304 585
R320 B.n426 B.n425 585
R321 B.n428 B.n303 585
R322 B.n431 B.n430 585
R323 B.n432 B.n302 585
R324 B.n434 B.n433 585
R325 B.n436 B.n301 585
R326 B.n439 B.n438 585
R327 B.n440 B.n300 585
R328 B.n442 B.n441 585
R329 B.n444 B.n299 585
R330 B.n447 B.n446 585
R331 B.n448 B.n298 585
R332 B.n450 B.n449 585
R333 B.n452 B.n297 585
R334 B.n455 B.n454 585
R335 B.n456 B.n296 585
R336 B.n458 B.n457 585
R337 B.n460 B.n295 585
R338 B.n463 B.n462 585
R339 B.n464 B.n294 585
R340 B.n466 B.n465 585
R341 B.n468 B.n293 585
R342 B.n471 B.n470 585
R343 B.n472 B.n292 585
R344 B.n474 B.n473 585
R345 B.n476 B.n291 585
R346 B.n479 B.n478 585
R347 B.n480 B.n290 585
R348 B.n482 B.n481 585
R349 B.n484 B.n289 585
R350 B.n487 B.n486 585
R351 B.n488 B.n288 585
R352 B.n490 B.n489 585
R353 B.n492 B.n287 585
R354 B.n495 B.n494 585
R355 B.n496 B.n286 585
R356 B.n501 B.n500 585
R357 B.n500 B.n499 585
R358 B.n502 B.n282 585
R359 B.n282 B.n281 585
R360 B.n504 B.n503 585
R361 B.n505 B.n504 585
R362 B.n276 B.n275 585
R363 B.n277 B.n276 585
R364 B.n513 B.n512 585
R365 B.n512 B.n511 585
R366 B.n514 B.n274 585
R367 B.n274 B.n273 585
R368 B.n516 B.n515 585
R369 B.n517 B.n516 585
R370 B.n268 B.n267 585
R371 B.n269 B.n268 585
R372 B.n526 B.n525 585
R373 B.n525 B.n524 585
R374 B.n527 B.n266 585
R375 B.n523 B.n266 585
R376 B.n529 B.n528 585
R377 B.n530 B.n529 585
R378 B.n261 B.n260 585
R379 B.n265 B.n261 585
R380 B.n539 B.n538 585
R381 B.n538 B.n537 585
R382 B.n540 B.n259 585
R383 B.n536 B.n259 585
R384 B.n542 B.n541 585
R385 B.n543 B.n542 585
R386 B.n254 B.n253 585
R387 B.n258 B.n254 585
R388 B.n553 B.n552 585
R389 B.n552 B.n551 585
R390 B.n554 B.n252 585
R391 B.n550 B.n252 585
R392 B.n556 B.n555 585
R393 B.n557 B.n556 585
R394 B.n2 B.n0 585
R395 B.n4 B.n2 585
R396 B.n3 B.n1 585
R397 B.n629 B.n3 585
R398 B.n627 B.n626 585
R399 B.n628 B.n627 585
R400 B.n625 B.n8 585
R401 B.n11 B.n8 585
R402 B.n624 B.n623 585
R403 B.n623 B.n622 585
R404 B.n10 B.n9 585
R405 B.n621 B.n10 585
R406 B.n619 B.n618 585
R407 B.n620 B.n619 585
R408 B.n617 B.n15 585
R409 B.n18 B.n15 585
R410 B.n616 B.n615 585
R411 B.n615 B.n614 585
R412 B.n17 B.n16 585
R413 B.n613 B.n17 585
R414 B.n611 B.n610 585
R415 B.n612 B.n611 585
R416 B.n609 B.n22 585
R417 B.n25 B.n22 585
R418 B.n608 B.n607 585
R419 B.n607 B.n606 585
R420 B.n24 B.n23 585
R421 B.n605 B.n24 585
R422 B.n603 B.n602 585
R423 B.n604 B.n603 585
R424 B.n601 B.n30 585
R425 B.n30 B.n29 585
R426 B.n600 B.n599 585
R427 B.n599 B.n598 585
R428 B.n32 B.n31 585
R429 B.n597 B.n32 585
R430 B.n595 B.n594 585
R431 B.n596 B.n595 585
R432 B.n593 B.n37 585
R433 B.n37 B.n36 585
R434 B.n592 B.n591 585
R435 B.n591 B.n590 585
R436 B.n632 B.n631 585
R437 B.n631 B.n630 585
R438 B.n500 B.n284 530.939
R439 B.n591 B.n39 530.939
R440 B.n498 B.n286 530.939
R441 B.n588 B.n40 530.939
R442 B.n589 B.n81 256.663
R443 B.n589 B.n80 256.663
R444 B.n589 B.n79 256.663
R445 B.n589 B.n78 256.663
R446 B.n589 B.n77 256.663
R447 B.n589 B.n76 256.663
R448 B.n589 B.n75 256.663
R449 B.n589 B.n74 256.663
R450 B.n589 B.n73 256.663
R451 B.n589 B.n72 256.663
R452 B.n589 B.n71 256.663
R453 B.n589 B.n70 256.663
R454 B.n589 B.n69 256.663
R455 B.n589 B.n68 256.663
R456 B.n589 B.n67 256.663
R457 B.n589 B.n66 256.663
R458 B.n589 B.n65 256.663
R459 B.n589 B.n64 256.663
R460 B.n589 B.n63 256.663
R461 B.n589 B.n62 256.663
R462 B.n589 B.n61 256.663
R463 B.n589 B.n60 256.663
R464 B.n589 B.n59 256.663
R465 B.n589 B.n58 256.663
R466 B.n589 B.n57 256.663
R467 B.n589 B.n56 256.663
R468 B.n589 B.n55 256.663
R469 B.n589 B.n54 256.663
R470 B.n589 B.n53 256.663
R471 B.n589 B.n52 256.663
R472 B.n589 B.n51 256.663
R473 B.n589 B.n50 256.663
R474 B.n589 B.n49 256.663
R475 B.n589 B.n48 256.663
R476 B.n589 B.n47 256.663
R477 B.n589 B.n46 256.663
R478 B.n589 B.n45 256.663
R479 B.n589 B.n44 256.663
R480 B.n589 B.n43 256.663
R481 B.n589 B.n42 256.663
R482 B.n589 B.n41 256.663
R483 B.n332 B.n285 256.663
R484 B.n338 B.n285 256.663
R485 B.n340 B.n285 256.663
R486 B.n346 B.n285 256.663
R487 B.n348 B.n285 256.663
R488 B.n354 B.n285 256.663
R489 B.n356 B.n285 256.663
R490 B.n362 B.n285 256.663
R491 B.n364 B.n285 256.663
R492 B.n370 B.n285 256.663
R493 B.n372 B.n285 256.663
R494 B.n378 B.n285 256.663
R495 B.n380 B.n285 256.663
R496 B.n386 B.n285 256.663
R497 B.n388 B.n285 256.663
R498 B.n394 B.n285 256.663
R499 B.n396 B.n285 256.663
R500 B.n402 B.n285 256.663
R501 B.n404 B.n285 256.663
R502 B.n410 B.n285 256.663
R503 B.n412 B.n285 256.663
R504 B.n418 B.n285 256.663
R505 B.n420 B.n285 256.663
R506 B.n427 B.n285 256.663
R507 B.n429 B.n285 256.663
R508 B.n435 B.n285 256.663
R509 B.n437 B.n285 256.663
R510 B.n443 B.n285 256.663
R511 B.n445 B.n285 256.663
R512 B.n451 B.n285 256.663
R513 B.n453 B.n285 256.663
R514 B.n459 B.n285 256.663
R515 B.n461 B.n285 256.663
R516 B.n467 B.n285 256.663
R517 B.n469 B.n285 256.663
R518 B.n475 B.n285 256.663
R519 B.n477 B.n285 256.663
R520 B.n483 B.n285 256.663
R521 B.n485 B.n285 256.663
R522 B.n491 B.n285 256.663
R523 B.n493 B.n285 256.663
R524 B.n500 B.n282 163.367
R525 B.n504 B.n282 163.367
R526 B.n504 B.n276 163.367
R527 B.n512 B.n276 163.367
R528 B.n512 B.n274 163.367
R529 B.n516 B.n274 163.367
R530 B.n516 B.n268 163.367
R531 B.n525 B.n268 163.367
R532 B.n525 B.n266 163.367
R533 B.n529 B.n266 163.367
R534 B.n529 B.n261 163.367
R535 B.n538 B.n261 163.367
R536 B.n538 B.n259 163.367
R537 B.n542 B.n259 163.367
R538 B.n542 B.n254 163.367
R539 B.n552 B.n254 163.367
R540 B.n552 B.n252 163.367
R541 B.n556 B.n252 163.367
R542 B.n556 B.n2 163.367
R543 B.n631 B.n2 163.367
R544 B.n631 B.n3 163.367
R545 B.n627 B.n3 163.367
R546 B.n627 B.n8 163.367
R547 B.n623 B.n8 163.367
R548 B.n623 B.n10 163.367
R549 B.n619 B.n10 163.367
R550 B.n619 B.n15 163.367
R551 B.n615 B.n15 163.367
R552 B.n615 B.n17 163.367
R553 B.n611 B.n17 163.367
R554 B.n611 B.n22 163.367
R555 B.n607 B.n22 163.367
R556 B.n607 B.n24 163.367
R557 B.n603 B.n24 163.367
R558 B.n603 B.n30 163.367
R559 B.n599 B.n30 163.367
R560 B.n599 B.n32 163.367
R561 B.n595 B.n32 163.367
R562 B.n595 B.n37 163.367
R563 B.n591 B.n37 163.367
R564 B.n333 B.n331 163.367
R565 B.n337 B.n331 163.367
R566 B.n341 B.n339 163.367
R567 B.n345 B.n329 163.367
R568 B.n349 B.n347 163.367
R569 B.n353 B.n327 163.367
R570 B.n357 B.n355 163.367
R571 B.n361 B.n325 163.367
R572 B.n365 B.n363 163.367
R573 B.n369 B.n323 163.367
R574 B.n373 B.n371 163.367
R575 B.n377 B.n321 163.367
R576 B.n381 B.n379 163.367
R577 B.n385 B.n319 163.367
R578 B.n389 B.n387 163.367
R579 B.n393 B.n317 163.367
R580 B.n397 B.n395 163.367
R581 B.n401 B.n315 163.367
R582 B.n405 B.n403 163.367
R583 B.n409 B.n310 163.367
R584 B.n413 B.n411 163.367
R585 B.n417 B.n308 163.367
R586 B.n421 B.n419 163.367
R587 B.n426 B.n304 163.367
R588 B.n430 B.n428 163.367
R589 B.n434 B.n302 163.367
R590 B.n438 B.n436 163.367
R591 B.n442 B.n300 163.367
R592 B.n446 B.n444 163.367
R593 B.n450 B.n298 163.367
R594 B.n454 B.n452 163.367
R595 B.n458 B.n296 163.367
R596 B.n462 B.n460 163.367
R597 B.n466 B.n294 163.367
R598 B.n470 B.n468 163.367
R599 B.n474 B.n292 163.367
R600 B.n478 B.n476 163.367
R601 B.n482 B.n290 163.367
R602 B.n486 B.n484 163.367
R603 B.n490 B.n288 163.367
R604 B.n494 B.n492 163.367
R605 B.n498 B.n280 163.367
R606 B.n506 B.n280 163.367
R607 B.n506 B.n278 163.367
R608 B.n510 B.n278 163.367
R609 B.n510 B.n272 163.367
R610 B.n518 B.n272 163.367
R611 B.n518 B.n270 163.367
R612 B.n522 B.n270 163.367
R613 B.n522 B.n264 163.367
R614 B.n531 B.n264 163.367
R615 B.n531 B.n262 163.367
R616 B.n535 B.n262 163.367
R617 B.n535 B.n257 163.367
R618 B.n544 B.n257 163.367
R619 B.n544 B.n255 163.367
R620 B.n549 B.n255 163.367
R621 B.n549 B.n251 163.367
R622 B.n558 B.n251 163.367
R623 B.n559 B.n558 163.367
R624 B.n559 B.n5 163.367
R625 B.n6 B.n5 163.367
R626 B.n7 B.n6 163.367
R627 B.n564 B.n7 163.367
R628 B.n564 B.n12 163.367
R629 B.n13 B.n12 163.367
R630 B.n14 B.n13 163.367
R631 B.n569 B.n14 163.367
R632 B.n569 B.n19 163.367
R633 B.n20 B.n19 163.367
R634 B.n21 B.n20 163.367
R635 B.n574 B.n21 163.367
R636 B.n574 B.n26 163.367
R637 B.n27 B.n26 163.367
R638 B.n28 B.n27 163.367
R639 B.n579 B.n28 163.367
R640 B.n579 B.n33 163.367
R641 B.n34 B.n33 163.367
R642 B.n35 B.n34 163.367
R643 B.n584 B.n35 163.367
R644 B.n584 B.n40 163.367
R645 B.n90 B.n89 163.367
R646 B.n94 B.n93 163.367
R647 B.n98 B.n97 163.367
R648 B.n102 B.n101 163.367
R649 B.n106 B.n105 163.367
R650 B.n110 B.n109 163.367
R651 B.n114 B.n113 163.367
R652 B.n118 B.n117 163.367
R653 B.n122 B.n121 163.367
R654 B.n126 B.n125 163.367
R655 B.n130 B.n129 163.367
R656 B.n134 B.n133 163.367
R657 B.n138 B.n137 163.367
R658 B.n142 B.n141 163.367
R659 B.n146 B.n145 163.367
R660 B.n150 B.n149 163.367
R661 B.n154 B.n153 163.367
R662 B.n158 B.n157 163.367
R663 B.n163 B.n162 163.367
R664 B.n167 B.n166 163.367
R665 B.n171 B.n170 163.367
R666 B.n175 B.n174 163.367
R667 B.n179 B.n178 163.367
R668 B.n183 B.n182 163.367
R669 B.n187 B.n186 163.367
R670 B.n191 B.n190 163.367
R671 B.n195 B.n194 163.367
R672 B.n199 B.n198 163.367
R673 B.n203 B.n202 163.367
R674 B.n207 B.n206 163.367
R675 B.n211 B.n210 163.367
R676 B.n215 B.n214 163.367
R677 B.n219 B.n218 163.367
R678 B.n223 B.n222 163.367
R679 B.n227 B.n226 163.367
R680 B.n231 B.n230 163.367
R681 B.n235 B.n234 163.367
R682 B.n239 B.n238 163.367
R683 B.n243 B.n242 163.367
R684 B.n247 B.n246 163.367
R685 B.n588 B.n82 163.367
R686 B.n499 B.n285 100.996
R687 B.n590 B.n589 100.996
R688 B.n305 B.t19 83.381
R689 B.n83 B.t11 83.381
R690 B.n311 B.t16 83.3682
R691 B.n86 B.t8 83.3682
R692 B.n332 B.n284 71.676
R693 B.n338 B.n337 71.676
R694 B.n341 B.n340 71.676
R695 B.n346 B.n345 71.676
R696 B.n349 B.n348 71.676
R697 B.n354 B.n353 71.676
R698 B.n357 B.n356 71.676
R699 B.n362 B.n361 71.676
R700 B.n365 B.n364 71.676
R701 B.n370 B.n369 71.676
R702 B.n373 B.n372 71.676
R703 B.n378 B.n377 71.676
R704 B.n381 B.n380 71.676
R705 B.n386 B.n385 71.676
R706 B.n389 B.n388 71.676
R707 B.n394 B.n393 71.676
R708 B.n397 B.n396 71.676
R709 B.n402 B.n401 71.676
R710 B.n405 B.n404 71.676
R711 B.n410 B.n409 71.676
R712 B.n413 B.n412 71.676
R713 B.n418 B.n417 71.676
R714 B.n421 B.n420 71.676
R715 B.n427 B.n426 71.676
R716 B.n430 B.n429 71.676
R717 B.n435 B.n434 71.676
R718 B.n438 B.n437 71.676
R719 B.n443 B.n442 71.676
R720 B.n446 B.n445 71.676
R721 B.n451 B.n450 71.676
R722 B.n454 B.n453 71.676
R723 B.n459 B.n458 71.676
R724 B.n462 B.n461 71.676
R725 B.n467 B.n466 71.676
R726 B.n470 B.n469 71.676
R727 B.n475 B.n474 71.676
R728 B.n478 B.n477 71.676
R729 B.n483 B.n482 71.676
R730 B.n486 B.n485 71.676
R731 B.n491 B.n490 71.676
R732 B.n494 B.n493 71.676
R733 B.n41 B.n39 71.676
R734 B.n90 B.n42 71.676
R735 B.n94 B.n43 71.676
R736 B.n98 B.n44 71.676
R737 B.n102 B.n45 71.676
R738 B.n106 B.n46 71.676
R739 B.n110 B.n47 71.676
R740 B.n114 B.n48 71.676
R741 B.n118 B.n49 71.676
R742 B.n122 B.n50 71.676
R743 B.n126 B.n51 71.676
R744 B.n130 B.n52 71.676
R745 B.n134 B.n53 71.676
R746 B.n138 B.n54 71.676
R747 B.n142 B.n55 71.676
R748 B.n146 B.n56 71.676
R749 B.n150 B.n57 71.676
R750 B.n154 B.n58 71.676
R751 B.n158 B.n59 71.676
R752 B.n163 B.n60 71.676
R753 B.n167 B.n61 71.676
R754 B.n171 B.n62 71.676
R755 B.n175 B.n63 71.676
R756 B.n179 B.n64 71.676
R757 B.n183 B.n65 71.676
R758 B.n187 B.n66 71.676
R759 B.n191 B.n67 71.676
R760 B.n195 B.n68 71.676
R761 B.n199 B.n69 71.676
R762 B.n203 B.n70 71.676
R763 B.n207 B.n71 71.676
R764 B.n211 B.n72 71.676
R765 B.n215 B.n73 71.676
R766 B.n219 B.n74 71.676
R767 B.n223 B.n75 71.676
R768 B.n227 B.n76 71.676
R769 B.n231 B.n77 71.676
R770 B.n235 B.n78 71.676
R771 B.n239 B.n79 71.676
R772 B.n243 B.n80 71.676
R773 B.n247 B.n81 71.676
R774 B.n82 B.n81 71.676
R775 B.n246 B.n80 71.676
R776 B.n242 B.n79 71.676
R777 B.n238 B.n78 71.676
R778 B.n234 B.n77 71.676
R779 B.n230 B.n76 71.676
R780 B.n226 B.n75 71.676
R781 B.n222 B.n74 71.676
R782 B.n218 B.n73 71.676
R783 B.n214 B.n72 71.676
R784 B.n210 B.n71 71.676
R785 B.n206 B.n70 71.676
R786 B.n202 B.n69 71.676
R787 B.n198 B.n68 71.676
R788 B.n194 B.n67 71.676
R789 B.n190 B.n66 71.676
R790 B.n186 B.n65 71.676
R791 B.n182 B.n64 71.676
R792 B.n178 B.n63 71.676
R793 B.n174 B.n62 71.676
R794 B.n170 B.n61 71.676
R795 B.n166 B.n60 71.676
R796 B.n162 B.n59 71.676
R797 B.n157 B.n58 71.676
R798 B.n153 B.n57 71.676
R799 B.n149 B.n56 71.676
R800 B.n145 B.n55 71.676
R801 B.n141 B.n54 71.676
R802 B.n137 B.n53 71.676
R803 B.n133 B.n52 71.676
R804 B.n129 B.n51 71.676
R805 B.n125 B.n50 71.676
R806 B.n121 B.n49 71.676
R807 B.n117 B.n48 71.676
R808 B.n113 B.n47 71.676
R809 B.n109 B.n46 71.676
R810 B.n105 B.n45 71.676
R811 B.n101 B.n44 71.676
R812 B.n97 B.n43 71.676
R813 B.n93 B.n42 71.676
R814 B.n89 B.n41 71.676
R815 B.n333 B.n332 71.676
R816 B.n339 B.n338 71.676
R817 B.n340 B.n329 71.676
R818 B.n347 B.n346 71.676
R819 B.n348 B.n327 71.676
R820 B.n355 B.n354 71.676
R821 B.n356 B.n325 71.676
R822 B.n363 B.n362 71.676
R823 B.n364 B.n323 71.676
R824 B.n371 B.n370 71.676
R825 B.n372 B.n321 71.676
R826 B.n379 B.n378 71.676
R827 B.n380 B.n319 71.676
R828 B.n387 B.n386 71.676
R829 B.n388 B.n317 71.676
R830 B.n395 B.n394 71.676
R831 B.n396 B.n315 71.676
R832 B.n403 B.n402 71.676
R833 B.n404 B.n310 71.676
R834 B.n411 B.n410 71.676
R835 B.n412 B.n308 71.676
R836 B.n419 B.n418 71.676
R837 B.n420 B.n304 71.676
R838 B.n428 B.n427 71.676
R839 B.n429 B.n302 71.676
R840 B.n436 B.n435 71.676
R841 B.n437 B.n300 71.676
R842 B.n444 B.n443 71.676
R843 B.n445 B.n298 71.676
R844 B.n452 B.n451 71.676
R845 B.n453 B.n296 71.676
R846 B.n460 B.n459 71.676
R847 B.n461 B.n294 71.676
R848 B.n468 B.n467 71.676
R849 B.n469 B.n292 71.676
R850 B.n476 B.n475 71.676
R851 B.n477 B.n290 71.676
R852 B.n484 B.n483 71.676
R853 B.n485 B.n288 71.676
R854 B.n492 B.n491 71.676
R855 B.n493 B.n286 71.676
R856 B.n306 B.t18 69.9991
R857 B.n84 B.t12 69.9991
R858 B.n312 B.t15 69.9864
R859 B.n87 B.t9 69.9864
R860 B.n423 B.n306 59.5399
R861 B.n313 B.n312 59.5399
R862 B.n160 B.n87 59.5399
R863 B.n85 B.n84 59.5399
R864 B.n499 B.n281 48.0262
R865 B.n505 B.n281 48.0262
R866 B.n505 B.n277 48.0262
R867 B.n511 B.n277 48.0262
R868 B.n517 B.n273 48.0262
R869 B.n517 B.n269 48.0262
R870 B.n524 B.n269 48.0262
R871 B.n524 B.n523 48.0262
R872 B.n530 B.n265 48.0262
R873 B.n537 B.n536 48.0262
R874 B.n543 B.n258 48.0262
R875 B.n551 B.n550 48.0262
R876 B.n557 B.n4 48.0262
R877 B.n630 B.n4 48.0262
R878 B.n630 B.n629 48.0262
R879 B.n629 B.n628 48.0262
R880 B.n622 B.n11 48.0262
R881 B.n621 B.n620 48.0262
R882 B.n614 B.n18 48.0262
R883 B.n613 B.n612 48.0262
R884 B.n606 B.n25 48.0262
R885 B.n606 B.n605 48.0262
R886 B.n605 B.n604 48.0262
R887 B.n604 B.n29 48.0262
R888 B.n598 B.n597 48.0262
R889 B.n597 B.n596 48.0262
R890 B.n596 B.n36 48.0262
R891 B.n590 B.n36 48.0262
R892 B.t14 B.n273 46.6137
R893 B.t7 B.n29 46.6137
R894 B.n530 B.t4 35.3135
R895 B.n612 B.t3 35.3135
R896 B.n592 B.n38 34.4981
R897 B.n587 B.n586 34.4981
R898 B.n497 B.n496 34.4981
R899 B.n501 B.n283 34.4981
R900 B.n537 B.t21 33.901
R901 B.n614 B.t2 33.901
R902 B.n543 B.t20 32.4885
R903 B.n620 B.t23 32.4885
R904 B.n551 B.t0 31.0759
R905 B.n622 B.t1 31.0759
R906 B.n557 B.t22 29.6634
R907 B.n628 B.t5 29.6634
R908 B.n550 B.t22 18.3633
R909 B.n11 B.t5 18.3633
R910 B B.n632 18.0485
R911 B.n258 B.t0 16.9507
R912 B.t1 B.n621 16.9507
R913 B.n536 B.t20 15.5382
R914 B.n18 B.t23 15.5382
R915 B.n265 B.t21 14.1257
R916 B.t2 B.n613 14.1257
R917 B.n306 B.n305 13.3823
R918 B.n312 B.n311 13.3823
R919 B.n87 B.n86 13.3823
R920 B.n84 B.n83 13.3823
R921 B.n523 B.t4 12.7132
R922 B.n25 B.t3 12.7132
R923 B.n88 B.n38 10.6151
R924 B.n91 B.n88 10.6151
R925 B.n92 B.n91 10.6151
R926 B.n95 B.n92 10.6151
R927 B.n96 B.n95 10.6151
R928 B.n99 B.n96 10.6151
R929 B.n100 B.n99 10.6151
R930 B.n103 B.n100 10.6151
R931 B.n104 B.n103 10.6151
R932 B.n107 B.n104 10.6151
R933 B.n108 B.n107 10.6151
R934 B.n111 B.n108 10.6151
R935 B.n112 B.n111 10.6151
R936 B.n115 B.n112 10.6151
R937 B.n116 B.n115 10.6151
R938 B.n119 B.n116 10.6151
R939 B.n120 B.n119 10.6151
R940 B.n123 B.n120 10.6151
R941 B.n124 B.n123 10.6151
R942 B.n127 B.n124 10.6151
R943 B.n128 B.n127 10.6151
R944 B.n131 B.n128 10.6151
R945 B.n132 B.n131 10.6151
R946 B.n135 B.n132 10.6151
R947 B.n136 B.n135 10.6151
R948 B.n139 B.n136 10.6151
R949 B.n140 B.n139 10.6151
R950 B.n143 B.n140 10.6151
R951 B.n144 B.n143 10.6151
R952 B.n147 B.n144 10.6151
R953 B.n148 B.n147 10.6151
R954 B.n151 B.n148 10.6151
R955 B.n152 B.n151 10.6151
R956 B.n155 B.n152 10.6151
R957 B.n156 B.n155 10.6151
R958 B.n159 B.n156 10.6151
R959 B.n164 B.n161 10.6151
R960 B.n165 B.n164 10.6151
R961 B.n168 B.n165 10.6151
R962 B.n169 B.n168 10.6151
R963 B.n172 B.n169 10.6151
R964 B.n173 B.n172 10.6151
R965 B.n176 B.n173 10.6151
R966 B.n177 B.n176 10.6151
R967 B.n181 B.n180 10.6151
R968 B.n184 B.n181 10.6151
R969 B.n185 B.n184 10.6151
R970 B.n188 B.n185 10.6151
R971 B.n189 B.n188 10.6151
R972 B.n192 B.n189 10.6151
R973 B.n193 B.n192 10.6151
R974 B.n196 B.n193 10.6151
R975 B.n197 B.n196 10.6151
R976 B.n200 B.n197 10.6151
R977 B.n201 B.n200 10.6151
R978 B.n204 B.n201 10.6151
R979 B.n205 B.n204 10.6151
R980 B.n208 B.n205 10.6151
R981 B.n209 B.n208 10.6151
R982 B.n212 B.n209 10.6151
R983 B.n213 B.n212 10.6151
R984 B.n216 B.n213 10.6151
R985 B.n217 B.n216 10.6151
R986 B.n220 B.n217 10.6151
R987 B.n221 B.n220 10.6151
R988 B.n224 B.n221 10.6151
R989 B.n225 B.n224 10.6151
R990 B.n228 B.n225 10.6151
R991 B.n229 B.n228 10.6151
R992 B.n232 B.n229 10.6151
R993 B.n233 B.n232 10.6151
R994 B.n236 B.n233 10.6151
R995 B.n237 B.n236 10.6151
R996 B.n240 B.n237 10.6151
R997 B.n241 B.n240 10.6151
R998 B.n244 B.n241 10.6151
R999 B.n245 B.n244 10.6151
R1000 B.n248 B.n245 10.6151
R1001 B.n249 B.n248 10.6151
R1002 B.n587 B.n249 10.6151
R1003 B.n497 B.n279 10.6151
R1004 B.n507 B.n279 10.6151
R1005 B.n508 B.n507 10.6151
R1006 B.n509 B.n508 10.6151
R1007 B.n509 B.n271 10.6151
R1008 B.n519 B.n271 10.6151
R1009 B.n520 B.n519 10.6151
R1010 B.n521 B.n520 10.6151
R1011 B.n521 B.n263 10.6151
R1012 B.n532 B.n263 10.6151
R1013 B.n533 B.n532 10.6151
R1014 B.n534 B.n533 10.6151
R1015 B.n534 B.n256 10.6151
R1016 B.n545 B.n256 10.6151
R1017 B.n546 B.n545 10.6151
R1018 B.n548 B.n546 10.6151
R1019 B.n548 B.n547 10.6151
R1020 B.n547 B.n250 10.6151
R1021 B.n560 B.n250 10.6151
R1022 B.n561 B.n560 10.6151
R1023 B.n562 B.n561 10.6151
R1024 B.n563 B.n562 10.6151
R1025 B.n565 B.n563 10.6151
R1026 B.n566 B.n565 10.6151
R1027 B.n567 B.n566 10.6151
R1028 B.n568 B.n567 10.6151
R1029 B.n570 B.n568 10.6151
R1030 B.n571 B.n570 10.6151
R1031 B.n572 B.n571 10.6151
R1032 B.n573 B.n572 10.6151
R1033 B.n575 B.n573 10.6151
R1034 B.n576 B.n575 10.6151
R1035 B.n577 B.n576 10.6151
R1036 B.n578 B.n577 10.6151
R1037 B.n580 B.n578 10.6151
R1038 B.n581 B.n580 10.6151
R1039 B.n582 B.n581 10.6151
R1040 B.n583 B.n582 10.6151
R1041 B.n585 B.n583 10.6151
R1042 B.n586 B.n585 10.6151
R1043 B.n334 B.n283 10.6151
R1044 B.n335 B.n334 10.6151
R1045 B.n336 B.n335 10.6151
R1046 B.n336 B.n330 10.6151
R1047 B.n342 B.n330 10.6151
R1048 B.n343 B.n342 10.6151
R1049 B.n344 B.n343 10.6151
R1050 B.n344 B.n328 10.6151
R1051 B.n350 B.n328 10.6151
R1052 B.n351 B.n350 10.6151
R1053 B.n352 B.n351 10.6151
R1054 B.n352 B.n326 10.6151
R1055 B.n358 B.n326 10.6151
R1056 B.n359 B.n358 10.6151
R1057 B.n360 B.n359 10.6151
R1058 B.n360 B.n324 10.6151
R1059 B.n366 B.n324 10.6151
R1060 B.n367 B.n366 10.6151
R1061 B.n368 B.n367 10.6151
R1062 B.n368 B.n322 10.6151
R1063 B.n374 B.n322 10.6151
R1064 B.n375 B.n374 10.6151
R1065 B.n376 B.n375 10.6151
R1066 B.n376 B.n320 10.6151
R1067 B.n382 B.n320 10.6151
R1068 B.n383 B.n382 10.6151
R1069 B.n384 B.n383 10.6151
R1070 B.n384 B.n318 10.6151
R1071 B.n390 B.n318 10.6151
R1072 B.n391 B.n390 10.6151
R1073 B.n392 B.n391 10.6151
R1074 B.n392 B.n316 10.6151
R1075 B.n398 B.n316 10.6151
R1076 B.n399 B.n398 10.6151
R1077 B.n400 B.n399 10.6151
R1078 B.n400 B.n314 10.6151
R1079 B.n407 B.n406 10.6151
R1080 B.n408 B.n407 10.6151
R1081 B.n408 B.n309 10.6151
R1082 B.n414 B.n309 10.6151
R1083 B.n415 B.n414 10.6151
R1084 B.n416 B.n415 10.6151
R1085 B.n416 B.n307 10.6151
R1086 B.n422 B.n307 10.6151
R1087 B.n425 B.n424 10.6151
R1088 B.n425 B.n303 10.6151
R1089 B.n431 B.n303 10.6151
R1090 B.n432 B.n431 10.6151
R1091 B.n433 B.n432 10.6151
R1092 B.n433 B.n301 10.6151
R1093 B.n439 B.n301 10.6151
R1094 B.n440 B.n439 10.6151
R1095 B.n441 B.n440 10.6151
R1096 B.n441 B.n299 10.6151
R1097 B.n447 B.n299 10.6151
R1098 B.n448 B.n447 10.6151
R1099 B.n449 B.n448 10.6151
R1100 B.n449 B.n297 10.6151
R1101 B.n455 B.n297 10.6151
R1102 B.n456 B.n455 10.6151
R1103 B.n457 B.n456 10.6151
R1104 B.n457 B.n295 10.6151
R1105 B.n463 B.n295 10.6151
R1106 B.n464 B.n463 10.6151
R1107 B.n465 B.n464 10.6151
R1108 B.n465 B.n293 10.6151
R1109 B.n471 B.n293 10.6151
R1110 B.n472 B.n471 10.6151
R1111 B.n473 B.n472 10.6151
R1112 B.n473 B.n291 10.6151
R1113 B.n479 B.n291 10.6151
R1114 B.n480 B.n479 10.6151
R1115 B.n481 B.n480 10.6151
R1116 B.n481 B.n289 10.6151
R1117 B.n487 B.n289 10.6151
R1118 B.n488 B.n487 10.6151
R1119 B.n489 B.n488 10.6151
R1120 B.n489 B.n287 10.6151
R1121 B.n495 B.n287 10.6151
R1122 B.n496 B.n495 10.6151
R1123 B.n502 B.n501 10.6151
R1124 B.n503 B.n502 10.6151
R1125 B.n503 B.n275 10.6151
R1126 B.n513 B.n275 10.6151
R1127 B.n514 B.n513 10.6151
R1128 B.n515 B.n514 10.6151
R1129 B.n515 B.n267 10.6151
R1130 B.n526 B.n267 10.6151
R1131 B.n527 B.n526 10.6151
R1132 B.n528 B.n527 10.6151
R1133 B.n528 B.n260 10.6151
R1134 B.n539 B.n260 10.6151
R1135 B.n540 B.n539 10.6151
R1136 B.n541 B.n540 10.6151
R1137 B.n541 B.n253 10.6151
R1138 B.n553 B.n253 10.6151
R1139 B.n554 B.n553 10.6151
R1140 B.n555 B.n554 10.6151
R1141 B.n555 B.n0 10.6151
R1142 B.n626 B.n1 10.6151
R1143 B.n626 B.n625 10.6151
R1144 B.n625 B.n624 10.6151
R1145 B.n624 B.n9 10.6151
R1146 B.n618 B.n9 10.6151
R1147 B.n618 B.n617 10.6151
R1148 B.n617 B.n616 10.6151
R1149 B.n616 B.n16 10.6151
R1150 B.n610 B.n16 10.6151
R1151 B.n610 B.n609 10.6151
R1152 B.n609 B.n608 10.6151
R1153 B.n608 B.n23 10.6151
R1154 B.n602 B.n23 10.6151
R1155 B.n602 B.n601 10.6151
R1156 B.n601 B.n600 10.6151
R1157 B.n600 B.n31 10.6151
R1158 B.n594 B.n31 10.6151
R1159 B.n594 B.n593 10.6151
R1160 B.n593 B.n592 10.6151
R1161 B.n161 B.n160 6.5566
R1162 B.n177 B.n85 6.5566
R1163 B.n406 B.n313 6.5566
R1164 B.n423 B.n422 6.5566
R1165 B.n160 B.n159 4.05904
R1166 B.n180 B.n85 4.05904
R1167 B.n314 B.n313 4.05904
R1168 B.n424 B.n423 4.05904
R1169 B.n632 B.n0 2.81026
R1170 B.n632 B.n1 2.81026
R1171 B.n511 B.t14 1.41302
R1172 B.n598 B.t7 1.41302
R1173 VN.n2 VN.t2 820.968
R1174 VN.n13 VN.t5 820.968
R1175 VN.n3 VN.t8 799.986
R1176 VN.n1 VN.t6 799.986
R1177 VN.n8 VN.t3 799.986
R1178 VN.n9 VN.t0 799.986
R1179 VN.n14 VN.t9 799.986
R1180 VN.n12 VN.t4 799.986
R1181 VN.n19 VN.t7 799.986
R1182 VN.n20 VN.t1 799.986
R1183 VN.n10 VN.n9 161.3
R1184 VN.n21 VN.n20 161.3
R1185 VN.n19 VN.n11 161.3
R1186 VN.n18 VN.n17 161.3
R1187 VN.n16 VN.n15 161.3
R1188 VN.n8 VN.n0 161.3
R1189 VN.n7 VN.n6 161.3
R1190 VN.n5 VN.n4 161.3
R1191 VN.n16 VN.n13 70.4033
R1192 VN.n5 VN.n2 70.4033
R1193 VN.n9 VN.n8 48.2005
R1194 VN.n20 VN.n19 48.2005
R1195 VN VN.n21 39.9986
R1196 VN.n4 VN.n3 37.9763
R1197 VN.n8 VN.n7 37.9763
R1198 VN.n15 VN.n14 37.9763
R1199 VN.n19 VN.n18 37.9763
R1200 VN.n14 VN.n13 20.9576
R1201 VN.n3 VN.n2 20.9576
R1202 VN.n4 VN.n1 10.2247
R1203 VN.n7 VN.n1 10.2247
R1204 VN.n15 VN.n12 10.2247
R1205 VN.n18 VN.n12 10.2247
R1206 VN.n21 VN.n11 0.189894
R1207 VN.n17 VN.n11 0.189894
R1208 VN.n17 VN.n16 0.189894
R1209 VN.n6 VN.n5 0.189894
R1210 VN.n6 VN.n0 0.189894
R1211 VN.n10 VN.n0 0.189894
R1212 VN VN.n10 0.0516364
R1213 VDD2.n1 VDD2.t7 64.612
R1214 VDD2.n4 VDD2.t8 64.0174
R1215 VDD2.n3 VDD2.n2 62.4857
R1216 VDD2 VDD2.n7 62.4829
R1217 VDD2.n6 VDD2.n5 62.0951
R1218 VDD2.n1 VDD2.n0 62.0949
R1219 VDD2.n4 VDD2.n3 35.42
R1220 VDD2.n7 VDD2.t0 1.92283
R1221 VDD2.n7 VDD2.t4 1.92283
R1222 VDD2.n5 VDD2.t2 1.92283
R1223 VDD2.n5 VDD2.t5 1.92283
R1224 VDD2.n2 VDD2.t6 1.92283
R1225 VDD2.n2 VDD2.t9 1.92283
R1226 VDD2.n0 VDD2.t1 1.92283
R1227 VDD2.n0 VDD2.t3 1.92283
R1228 VDD2.n6 VDD2.n4 0.595328
R1229 VDD2 VDD2.n6 0.207397
R1230 VDD2.n3 VDD2.n1 0.0938609
C0 VDD2 VP 0.297754f
C1 VDD2 VTAIL 16.8611f
C2 VN VP 4.78791f
C3 VN VTAIL 3.6205f
C4 VDD2 VDD1 0.761821f
C5 VTAIL VP 3.63514f
C6 VN VDD1 0.147899f
C7 VDD1 VP 4.05123f
C8 VTAIL VDD1 16.8296f
C9 VN VDD2 3.9058f
C10 VDD2 B 4.298054f
C11 VDD1 B 4.173601f
C12 VTAIL B 5.544244f
C13 VN B 7.81184f
C14 VP B 5.750705f
C15 VDD2.t7 B 2.5978f
C16 VDD2.t1 B 0.230986f
C17 VDD2.t3 B 0.230986f
C18 VDD2.n0 B 2.03759f
C19 VDD2.n1 B 0.670532f
C20 VDD2.t6 B 0.230986f
C21 VDD2.t9 B 0.230986f
C22 VDD2.n2 B 2.03969f
C23 VDD2.n3 B 1.83467f
C24 VDD2.t8 B 2.59439f
C25 VDD2.n4 B 2.40828f
C26 VDD2.t2 B 0.230986f
C27 VDD2.t5 B 0.230986f
C28 VDD2.n5 B 2.03759f
C29 VDD2.n6 B 0.3058f
C30 VDD2.t0 B 0.230986f
C31 VDD2.t4 B 0.230986f
C32 VDD2.n7 B 2.03966f
C33 VN.n0 B 0.05141f
C34 VN.t6 B 0.545465f
C35 VN.n1 B 0.222451f
C36 VN.t2 B 0.551337f
C37 VN.n2 B 0.224159f
C38 VN.t8 B 0.545465f
C39 VN.n3 B 0.23792f
C40 VN.n4 B 0.011666f
C41 VN.n5 B 0.157681f
C42 VN.n6 B 0.05141f
C43 VN.n7 B 0.011666f
C44 VN.t3 B 0.545465f
C45 VN.n8 B 0.23792f
C46 VN.t0 B 0.545465f
C47 VN.n9 B 0.229679f
C48 VN.n10 B 0.039841f
C49 VN.n11 B 0.05141f
C50 VN.t4 B 0.545465f
C51 VN.n12 B 0.222451f
C52 VN.t5 B 0.551337f
C53 VN.n13 B 0.224159f
C54 VN.t9 B 0.545465f
C55 VN.n14 B 0.23792f
C56 VN.n15 B 0.011666f
C57 VN.n16 B 0.157681f
C58 VN.n17 B 0.05141f
C59 VN.n18 B 0.011666f
C60 VN.t7 B 0.545465f
C61 VN.n19 B 0.23792f
C62 VN.t1 B 0.545465f
C63 VN.n20 B 0.229679f
C64 VN.n21 B 1.95533f
C65 VDD1.t6 B 2.59721f
C66 VDD1.t3 B 0.230933f
C67 VDD1.t9 B 0.230933f
C68 VDD1.n0 B 2.03712f
C69 VDD1.n1 B 0.673703f
C70 VDD1.t1 B 2.59721f
C71 VDD1.t7 B 0.230933f
C72 VDD1.t2 B 0.230933f
C73 VDD1.n2 B 2.03712f
C74 VDD1.n3 B 0.670377f
C75 VDD1.t5 B 0.230933f
C76 VDD1.t8 B 0.230933f
C77 VDD1.n4 B 2.03922f
C78 VDD1.n5 B 1.91231f
C79 VDD1.t4 B 0.230933f
C80 VDD1.t0 B 0.230933f
C81 VDD1.n6 B 2.03711f
C82 VDD1.n7 B 2.39678f
C83 VTAIL.t5 B 0.24063f
C84 VTAIL.t1 B 0.24063f
C85 VTAIL.n0 B 2.03578f
C86 VTAIL.n1 B 0.410026f
C87 VTAIL.t11 B 2.5925f
C88 VTAIL.n2 B 0.518197f
C89 VTAIL.t14 B 0.24063f
C90 VTAIL.t12 B 0.24063f
C91 VTAIL.n3 B 2.03578f
C92 VTAIL.n4 B 0.402224f
C93 VTAIL.t10 B 0.24063f
C94 VTAIL.t8 B 0.24063f
C95 VTAIL.n5 B 2.03578f
C96 VTAIL.n6 B 1.70633f
C97 VTAIL.t4 B 0.24063f
C98 VTAIL.t19 B 0.24063f
C99 VTAIL.n7 B 2.03579f
C100 VTAIL.n8 B 1.70632f
C101 VTAIL.t16 B 0.24063f
C102 VTAIL.t0 B 0.24063f
C103 VTAIL.n9 B 2.03579f
C104 VTAIL.n10 B 0.402218f
C105 VTAIL.t17 B 2.5925f
C106 VTAIL.n11 B 0.518191f
C107 VTAIL.t6 B 0.24063f
C108 VTAIL.t13 B 0.24063f
C109 VTAIL.n12 B 2.03579f
C110 VTAIL.n13 B 0.418642f
C111 VTAIL.t9 B 0.24063f
C112 VTAIL.t15 B 0.24063f
C113 VTAIL.n14 B 2.03579f
C114 VTAIL.n15 B 0.402218f
C115 VTAIL.t7 B 2.5925f
C116 VTAIL.n16 B 1.74921f
C117 VTAIL.t3 B 2.5925f
C118 VTAIL.n17 B 1.74921f
C119 VTAIL.t18 B 0.24063f
C120 VTAIL.t2 B 0.24063f
C121 VTAIL.n18 B 2.03578f
C122 VTAIL.n19 B 0.354183f
C123 VP.n0 B 0.052554f
C124 VP.t7 B 0.557611f
C125 VP.n1 B 0.227404f
C126 VP.n2 B 0.052554f
C127 VP.n3 B 0.052554f
C128 VP.t9 B 0.557611f
C129 VP.t5 B 0.557611f
C130 VP.t0 B 0.557611f
C131 VP.n4 B 0.227404f
C132 VP.t3 B 0.563613f
C133 VP.n5 B 0.22915f
C134 VP.t6 B 0.557611f
C135 VP.n6 B 0.243218f
C136 VP.n7 B 0.011926f
C137 VP.n8 B 0.161192f
C138 VP.n9 B 0.052554f
C139 VP.n10 B 0.011926f
C140 VP.n11 B 0.243218f
C141 VP.n12 B 0.234793f
C142 VP.n13 B 1.96424f
C143 VP.n14 B 2.01178f
C144 VP.t8 B 0.557611f
C145 VP.n15 B 0.234793f
C146 VP.t2 B 0.557611f
C147 VP.n16 B 0.243218f
C148 VP.n17 B 0.011926f
C149 VP.n18 B 0.052554f
C150 VP.n19 B 0.052554f
C151 VP.n20 B 0.011926f
C152 VP.t4 B 0.557611f
C153 VP.n21 B 0.243218f
C154 VP.t1 B 0.557611f
C155 VP.n22 B 0.234793f
C156 VP.n23 B 0.040728f
.ends

