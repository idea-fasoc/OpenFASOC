* NGSPICE file created from diff_pair_sample_1033.ext - technology: sky130A

.subckt diff_pair_sample_1033 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=0 ps=0 w=17.26 l=2.98
X1 VTAIL.t19 VP.t0 VDD1.t8 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X2 VTAIL.t0 VN.t0 VDD2.t9 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X3 VTAIL.t18 VP.t1 VDD1.t7 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X4 VTAIL.t1 VN.t1 VDD2.t8 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X5 VTAIL.t17 VP.t2 VDD1.t6 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X6 VDD1.t1 VP.t3 VTAIL.t16 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=2.8479 ps=17.59 w=17.26 l=2.98
X7 B.t8 B.t6 B.t7 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=0 ps=0 w=17.26 l=2.98
X8 VDD2.t7 VN.t2 VTAIL.t8 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=6.7314 ps=35.3 w=17.26 l=2.98
X9 B.t5 B.t3 B.t4 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=0 ps=0 w=17.26 l=2.98
X10 VDD2.t6 VN.t3 VTAIL.t7 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X11 VDD1.t9 VP.t4 VTAIL.t15 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X12 VDD2.t5 VN.t4 VTAIL.t6 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=6.7314 ps=35.3 w=17.26 l=2.98
X13 VDD1.t3 VP.t5 VTAIL.t14 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=6.7314 ps=35.3 w=17.26 l=2.98
X14 VTAIL.t5 VN.t5 VDD2.t4 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X15 VDD2.t3 VN.t6 VTAIL.t9 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=2.8479 ps=17.59 w=17.26 l=2.98
X16 VDD1.t4 VP.t6 VTAIL.t13 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X17 VTAIL.t12 VP.t7 VDD1.t0 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X18 B.t2 B.t0 B.t1 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=0 ps=0 w=17.26 l=2.98
X19 VDD2.t2 VN.t7 VTAIL.t4 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X20 VDD1.t5 VP.t8 VTAIL.t11 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=6.7314 ps=35.3 w=17.26 l=2.98
X21 VDD1.t2 VP.t9 VTAIL.t10 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=2.8479 ps=17.59 w=17.26 l=2.98
X22 VTAIL.t3 VN.t8 VDD2.t1 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=2.8479 pd=17.59 as=2.8479 ps=17.59 w=17.26 l=2.98
X23 VDD2.t0 VN.t9 VTAIL.t2 w_n4942_n4420# sky130_fd_pr__pfet_01v8 ad=6.7314 pd=35.3 as=2.8479 ps=17.59 w=17.26 l=2.98
R0 B.n552 B.n169 585
R1 B.n551 B.n550 585
R2 B.n549 B.n170 585
R3 B.n548 B.n547 585
R4 B.n546 B.n171 585
R5 B.n545 B.n544 585
R6 B.n543 B.n172 585
R7 B.n542 B.n541 585
R8 B.n540 B.n173 585
R9 B.n539 B.n538 585
R10 B.n537 B.n174 585
R11 B.n536 B.n535 585
R12 B.n534 B.n175 585
R13 B.n533 B.n532 585
R14 B.n531 B.n176 585
R15 B.n530 B.n529 585
R16 B.n528 B.n177 585
R17 B.n527 B.n526 585
R18 B.n525 B.n178 585
R19 B.n524 B.n523 585
R20 B.n522 B.n179 585
R21 B.n521 B.n520 585
R22 B.n519 B.n180 585
R23 B.n518 B.n517 585
R24 B.n516 B.n181 585
R25 B.n515 B.n514 585
R26 B.n513 B.n182 585
R27 B.n512 B.n511 585
R28 B.n510 B.n183 585
R29 B.n509 B.n508 585
R30 B.n507 B.n184 585
R31 B.n506 B.n505 585
R32 B.n504 B.n185 585
R33 B.n503 B.n502 585
R34 B.n501 B.n186 585
R35 B.n500 B.n499 585
R36 B.n498 B.n187 585
R37 B.n497 B.n496 585
R38 B.n495 B.n188 585
R39 B.n494 B.n493 585
R40 B.n492 B.n189 585
R41 B.n491 B.n490 585
R42 B.n489 B.n190 585
R43 B.n488 B.n487 585
R44 B.n486 B.n191 585
R45 B.n485 B.n484 585
R46 B.n483 B.n192 585
R47 B.n482 B.n481 585
R48 B.n480 B.n193 585
R49 B.n479 B.n478 585
R50 B.n477 B.n194 585
R51 B.n476 B.n475 585
R52 B.n474 B.n195 585
R53 B.n473 B.n472 585
R54 B.n471 B.n196 585
R55 B.n470 B.n469 585
R56 B.n468 B.n197 585
R57 B.n467 B.n466 585
R58 B.n462 B.n198 585
R59 B.n461 B.n460 585
R60 B.n459 B.n199 585
R61 B.n458 B.n457 585
R62 B.n456 B.n200 585
R63 B.n455 B.n454 585
R64 B.n453 B.n201 585
R65 B.n452 B.n451 585
R66 B.n450 B.n202 585
R67 B.n448 B.n447 585
R68 B.n446 B.n205 585
R69 B.n445 B.n444 585
R70 B.n443 B.n206 585
R71 B.n442 B.n441 585
R72 B.n440 B.n207 585
R73 B.n439 B.n438 585
R74 B.n437 B.n208 585
R75 B.n436 B.n435 585
R76 B.n434 B.n209 585
R77 B.n433 B.n432 585
R78 B.n431 B.n210 585
R79 B.n430 B.n429 585
R80 B.n428 B.n211 585
R81 B.n427 B.n426 585
R82 B.n425 B.n212 585
R83 B.n424 B.n423 585
R84 B.n422 B.n213 585
R85 B.n421 B.n420 585
R86 B.n419 B.n214 585
R87 B.n418 B.n417 585
R88 B.n416 B.n215 585
R89 B.n415 B.n414 585
R90 B.n413 B.n216 585
R91 B.n412 B.n411 585
R92 B.n410 B.n217 585
R93 B.n409 B.n408 585
R94 B.n407 B.n218 585
R95 B.n406 B.n405 585
R96 B.n404 B.n219 585
R97 B.n403 B.n402 585
R98 B.n401 B.n220 585
R99 B.n400 B.n399 585
R100 B.n398 B.n221 585
R101 B.n397 B.n396 585
R102 B.n395 B.n222 585
R103 B.n394 B.n393 585
R104 B.n392 B.n223 585
R105 B.n391 B.n390 585
R106 B.n389 B.n224 585
R107 B.n388 B.n387 585
R108 B.n386 B.n225 585
R109 B.n385 B.n384 585
R110 B.n383 B.n226 585
R111 B.n382 B.n381 585
R112 B.n380 B.n227 585
R113 B.n379 B.n378 585
R114 B.n377 B.n228 585
R115 B.n376 B.n375 585
R116 B.n374 B.n229 585
R117 B.n373 B.n372 585
R118 B.n371 B.n230 585
R119 B.n370 B.n369 585
R120 B.n368 B.n231 585
R121 B.n367 B.n366 585
R122 B.n365 B.n232 585
R123 B.n364 B.n363 585
R124 B.n554 B.n553 585
R125 B.n555 B.n168 585
R126 B.n557 B.n556 585
R127 B.n558 B.n167 585
R128 B.n560 B.n559 585
R129 B.n561 B.n166 585
R130 B.n563 B.n562 585
R131 B.n564 B.n165 585
R132 B.n566 B.n565 585
R133 B.n567 B.n164 585
R134 B.n569 B.n568 585
R135 B.n570 B.n163 585
R136 B.n572 B.n571 585
R137 B.n573 B.n162 585
R138 B.n575 B.n574 585
R139 B.n576 B.n161 585
R140 B.n578 B.n577 585
R141 B.n579 B.n160 585
R142 B.n581 B.n580 585
R143 B.n582 B.n159 585
R144 B.n584 B.n583 585
R145 B.n585 B.n158 585
R146 B.n587 B.n586 585
R147 B.n588 B.n157 585
R148 B.n590 B.n589 585
R149 B.n591 B.n156 585
R150 B.n593 B.n592 585
R151 B.n594 B.n155 585
R152 B.n596 B.n595 585
R153 B.n597 B.n154 585
R154 B.n599 B.n598 585
R155 B.n600 B.n153 585
R156 B.n602 B.n601 585
R157 B.n603 B.n152 585
R158 B.n605 B.n604 585
R159 B.n606 B.n151 585
R160 B.n608 B.n607 585
R161 B.n609 B.n150 585
R162 B.n611 B.n610 585
R163 B.n612 B.n149 585
R164 B.n614 B.n613 585
R165 B.n615 B.n148 585
R166 B.n617 B.n616 585
R167 B.n618 B.n147 585
R168 B.n620 B.n619 585
R169 B.n621 B.n146 585
R170 B.n623 B.n622 585
R171 B.n624 B.n145 585
R172 B.n626 B.n625 585
R173 B.n627 B.n144 585
R174 B.n629 B.n628 585
R175 B.n630 B.n143 585
R176 B.n632 B.n631 585
R177 B.n633 B.n142 585
R178 B.n635 B.n634 585
R179 B.n636 B.n141 585
R180 B.n638 B.n637 585
R181 B.n639 B.n140 585
R182 B.n641 B.n640 585
R183 B.n642 B.n139 585
R184 B.n644 B.n643 585
R185 B.n645 B.n138 585
R186 B.n647 B.n646 585
R187 B.n648 B.n137 585
R188 B.n650 B.n649 585
R189 B.n651 B.n136 585
R190 B.n653 B.n652 585
R191 B.n654 B.n135 585
R192 B.n656 B.n655 585
R193 B.n657 B.n134 585
R194 B.n659 B.n658 585
R195 B.n660 B.n133 585
R196 B.n662 B.n661 585
R197 B.n663 B.n132 585
R198 B.n665 B.n664 585
R199 B.n666 B.n131 585
R200 B.n668 B.n667 585
R201 B.n669 B.n130 585
R202 B.n671 B.n670 585
R203 B.n672 B.n129 585
R204 B.n674 B.n673 585
R205 B.n675 B.n128 585
R206 B.n677 B.n676 585
R207 B.n678 B.n127 585
R208 B.n680 B.n679 585
R209 B.n681 B.n126 585
R210 B.n683 B.n682 585
R211 B.n684 B.n125 585
R212 B.n686 B.n685 585
R213 B.n687 B.n124 585
R214 B.n689 B.n688 585
R215 B.n690 B.n123 585
R216 B.n692 B.n691 585
R217 B.n693 B.n122 585
R218 B.n695 B.n694 585
R219 B.n696 B.n121 585
R220 B.n698 B.n697 585
R221 B.n699 B.n120 585
R222 B.n701 B.n700 585
R223 B.n702 B.n119 585
R224 B.n704 B.n703 585
R225 B.n705 B.n118 585
R226 B.n707 B.n706 585
R227 B.n708 B.n117 585
R228 B.n710 B.n709 585
R229 B.n711 B.n116 585
R230 B.n713 B.n712 585
R231 B.n714 B.n115 585
R232 B.n716 B.n715 585
R233 B.n717 B.n114 585
R234 B.n719 B.n718 585
R235 B.n720 B.n113 585
R236 B.n722 B.n721 585
R237 B.n723 B.n112 585
R238 B.n725 B.n724 585
R239 B.n726 B.n111 585
R240 B.n728 B.n727 585
R241 B.n729 B.n110 585
R242 B.n731 B.n730 585
R243 B.n732 B.n109 585
R244 B.n734 B.n733 585
R245 B.n735 B.n108 585
R246 B.n737 B.n736 585
R247 B.n738 B.n107 585
R248 B.n740 B.n739 585
R249 B.n741 B.n106 585
R250 B.n743 B.n742 585
R251 B.n744 B.n105 585
R252 B.n746 B.n745 585
R253 B.n747 B.n104 585
R254 B.n749 B.n748 585
R255 B.n750 B.n103 585
R256 B.n752 B.n751 585
R257 B.n753 B.n102 585
R258 B.n940 B.n35 585
R259 B.n939 B.n938 585
R260 B.n937 B.n36 585
R261 B.n936 B.n935 585
R262 B.n934 B.n37 585
R263 B.n933 B.n932 585
R264 B.n931 B.n38 585
R265 B.n930 B.n929 585
R266 B.n928 B.n39 585
R267 B.n927 B.n926 585
R268 B.n925 B.n40 585
R269 B.n924 B.n923 585
R270 B.n922 B.n41 585
R271 B.n921 B.n920 585
R272 B.n919 B.n42 585
R273 B.n918 B.n917 585
R274 B.n916 B.n43 585
R275 B.n915 B.n914 585
R276 B.n913 B.n44 585
R277 B.n912 B.n911 585
R278 B.n910 B.n45 585
R279 B.n909 B.n908 585
R280 B.n907 B.n46 585
R281 B.n906 B.n905 585
R282 B.n904 B.n47 585
R283 B.n903 B.n902 585
R284 B.n901 B.n48 585
R285 B.n900 B.n899 585
R286 B.n898 B.n49 585
R287 B.n897 B.n896 585
R288 B.n895 B.n50 585
R289 B.n894 B.n893 585
R290 B.n892 B.n51 585
R291 B.n891 B.n890 585
R292 B.n889 B.n52 585
R293 B.n888 B.n887 585
R294 B.n886 B.n53 585
R295 B.n885 B.n884 585
R296 B.n883 B.n54 585
R297 B.n882 B.n881 585
R298 B.n880 B.n55 585
R299 B.n879 B.n878 585
R300 B.n877 B.n56 585
R301 B.n876 B.n875 585
R302 B.n874 B.n57 585
R303 B.n873 B.n872 585
R304 B.n871 B.n58 585
R305 B.n870 B.n869 585
R306 B.n868 B.n59 585
R307 B.n867 B.n866 585
R308 B.n865 B.n60 585
R309 B.n864 B.n863 585
R310 B.n862 B.n61 585
R311 B.n861 B.n860 585
R312 B.n859 B.n62 585
R313 B.n858 B.n857 585
R314 B.n856 B.n63 585
R315 B.n854 B.n853 585
R316 B.n852 B.n66 585
R317 B.n851 B.n850 585
R318 B.n849 B.n67 585
R319 B.n848 B.n847 585
R320 B.n846 B.n68 585
R321 B.n845 B.n844 585
R322 B.n843 B.n69 585
R323 B.n842 B.n841 585
R324 B.n840 B.n70 585
R325 B.n839 B.n838 585
R326 B.n837 B.n71 585
R327 B.n836 B.n835 585
R328 B.n834 B.n75 585
R329 B.n833 B.n832 585
R330 B.n831 B.n76 585
R331 B.n830 B.n829 585
R332 B.n828 B.n77 585
R333 B.n827 B.n826 585
R334 B.n825 B.n78 585
R335 B.n824 B.n823 585
R336 B.n822 B.n79 585
R337 B.n821 B.n820 585
R338 B.n819 B.n80 585
R339 B.n818 B.n817 585
R340 B.n816 B.n81 585
R341 B.n815 B.n814 585
R342 B.n813 B.n82 585
R343 B.n812 B.n811 585
R344 B.n810 B.n83 585
R345 B.n809 B.n808 585
R346 B.n807 B.n84 585
R347 B.n806 B.n805 585
R348 B.n804 B.n85 585
R349 B.n803 B.n802 585
R350 B.n801 B.n86 585
R351 B.n800 B.n799 585
R352 B.n798 B.n87 585
R353 B.n797 B.n796 585
R354 B.n795 B.n88 585
R355 B.n794 B.n793 585
R356 B.n792 B.n89 585
R357 B.n791 B.n790 585
R358 B.n789 B.n90 585
R359 B.n788 B.n787 585
R360 B.n786 B.n91 585
R361 B.n785 B.n784 585
R362 B.n783 B.n92 585
R363 B.n782 B.n781 585
R364 B.n780 B.n93 585
R365 B.n779 B.n778 585
R366 B.n777 B.n94 585
R367 B.n776 B.n775 585
R368 B.n774 B.n95 585
R369 B.n773 B.n772 585
R370 B.n771 B.n96 585
R371 B.n770 B.n769 585
R372 B.n768 B.n97 585
R373 B.n767 B.n766 585
R374 B.n765 B.n98 585
R375 B.n764 B.n763 585
R376 B.n762 B.n99 585
R377 B.n761 B.n760 585
R378 B.n759 B.n100 585
R379 B.n758 B.n757 585
R380 B.n756 B.n101 585
R381 B.n755 B.n754 585
R382 B.n942 B.n941 585
R383 B.n943 B.n34 585
R384 B.n945 B.n944 585
R385 B.n946 B.n33 585
R386 B.n948 B.n947 585
R387 B.n949 B.n32 585
R388 B.n951 B.n950 585
R389 B.n952 B.n31 585
R390 B.n954 B.n953 585
R391 B.n955 B.n30 585
R392 B.n957 B.n956 585
R393 B.n958 B.n29 585
R394 B.n960 B.n959 585
R395 B.n961 B.n28 585
R396 B.n963 B.n962 585
R397 B.n964 B.n27 585
R398 B.n966 B.n965 585
R399 B.n967 B.n26 585
R400 B.n969 B.n968 585
R401 B.n970 B.n25 585
R402 B.n972 B.n971 585
R403 B.n973 B.n24 585
R404 B.n975 B.n974 585
R405 B.n976 B.n23 585
R406 B.n978 B.n977 585
R407 B.n979 B.n22 585
R408 B.n981 B.n980 585
R409 B.n982 B.n21 585
R410 B.n984 B.n983 585
R411 B.n985 B.n20 585
R412 B.n987 B.n986 585
R413 B.n988 B.n19 585
R414 B.n990 B.n989 585
R415 B.n991 B.n18 585
R416 B.n993 B.n992 585
R417 B.n994 B.n17 585
R418 B.n996 B.n995 585
R419 B.n997 B.n16 585
R420 B.n999 B.n998 585
R421 B.n1000 B.n15 585
R422 B.n1002 B.n1001 585
R423 B.n1003 B.n14 585
R424 B.n1005 B.n1004 585
R425 B.n1006 B.n13 585
R426 B.n1008 B.n1007 585
R427 B.n1009 B.n12 585
R428 B.n1011 B.n1010 585
R429 B.n1012 B.n11 585
R430 B.n1014 B.n1013 585
R431 B.n1015 B.n10 585
R432 B.n1017 B.n1016 585
R433 B.n1018 B.n9 585
R434 B.n1020 B.n1019 585
R435 B.n1021 B.n8 585
R436 B.n1023 B.n1022 585
R437 B.n1024 B.n7 585
R438 B.n1026 B.n1025 585
R439 B.n1027 B.n6 585
R440 B.n1029 B.n1028 585
R441 B.n1030 B.n5 585
R442 B.n1032 B.n1031 585
R443 B.n1033 B.n4 585
R444 B.n1035 B.n1034 585
R445 B.n1036 B.n3 585
R446 B.n1038 B.n1037 585
R447 B.n1039 B.n0 585
R448 B.n2 B.n1 585
R449 B.n266 B.n265 585
R450 B.n268 B.n267 585
R451 B.n269 B.n264 585
R452 B.n271 B.n270 585
R453 B.n272 B.n263 585
R454 B.n274 B.n273 585
R455 B.n275 B.n262 585
R456 B.n277 B.n276 585
R457 B.n278 B.n261 585
R458 B.n280 B.n279 585
R459 B.n281 B.n260 585
R460 B.n283 B.n282 585
R461 B.n284 B.n259 585
R462 B.n286 B.n285 585
R463 B.n287 B.n258 585
R464 B.n289 B.n288 585
R465 B.n290 B.n257 585
R466 B.n292 B.n291 585
R467 B.n293 B.n256 585
R468 B.n295 B.n294 585
R469 B.n296 B.n255 585
R470 B.n298 B.n297 585
R471 B.n299 B.n254 585
R472 B.n301 B.n300 585
R473 B.n302 B.n253 585
R474 B.n304 B.n303 585
R475 B.n305 B.n252 585
R476 B.n307 B.n306 585
R477 B.n308 B.n251 585
R478 B.n310 B.n309 585
R479 B.n311 B.n250 585
R480 B.n313 B.n312 585
R481 B.n314 B.n249 585
R482 B.n316 B.n315 585
R483 B.n317 B.n248 585
R484 B.n319 B.n318 585
R485 B.n320 B.n247 585
R486 B.n322 B.n321 585
R487 B.n323 B.n246 585
R488 B.n325 B.n324 585
R489 B.n326 B.n245 585
R490 B.n328 B.n327 585
R491 B.n329 B.n244 585
R492 B.n331 B.n330 585
R493 B.n332 B.n243 585
R494 B.n334 B.n333 585
R495 B.n335 B.n242 585
R496 B.n337 B.n336 585
R497 B.n338 B.n241 585
R498 B.n340 B.n339 585
R499 B.n341 B.n240 585
R500 B.n343 B.n342 585
R501 B.n344 B.n239 585
R502 B.n346 B.n345 585
R503 B.n347 B.n238 585
R504 B.n349 B.n348 585
R505 B.n350 B.n237 585
R506 B.n352 B.n351 585
R507 B.n353 B.n236 585
R508 B.n355 B.n354 585
R509 B.n356 B.n235 585
R510 B.n358 B.n357 585
R511 B.n359 B.n234 585
R512 B.n361 B.n360 585
R513 B.n362 B.n233 585
R514 B.n363 B.n362 482.89
R515 B.n553 B.n552 482.89
R516 B.n755 B.n102 482.89
R517 B.n942 B.n35 482.89
R518 B.n203 B.t6 348.142
R519 B.n463 B.t9 348.142
R520 B.n72 B.t0 348.142
R521 B.n64 B.t3 348.142
R522 B.n1041 B.n1040 256.663
R523 B.n1040 B.n1039 235.042
R524 B.n1040 B.n2 235.042
R525 B.n463 B.t10 175.517
R526 B.n72 B.t2 175.517
R527 B.n203 B.t7 175.494
R528 B.n64 B.t5 175.494
R529 B.n363 B.n232 163.367
R530 B.n367 B.n232 163.367
R531 B.n368 B.n367 163.367
R532 B.n369 B.n368 163.367
R533 B.n369 B.n230 163.367
R534 B.n373 B.n230 163.367
R535 B.n374 B.n373 163.367
R536 B.n375 B.n374 163.367
R537 B.n375 B.n228 163.367
R538 B.n379 B.n228 163.367
R539 B.n380 B.n379 163.367
R540 B.n381 B.n380 163.367
R541 B.n381 B.n226 163.367
R542 B.n385 B.n226 163.367
R543 B.n386 B.n385 163.367
R544 B.n387 B.n386 163.367
R545 B.n387 B.n224 163.367
R546 B.n391 B.n224 163.367
R547 B.n392 B.n391 163.367
R548 B.n393 B.n392 163.367
R549 B.n393 B.n222 163.367
R550 B.n397 B.n222 163.367
R551 B.n398 B.n397 163.367
R552 B.n399 B.n398 163.367
R553 B.n399 B.n220 163.367
R554 B.n403 B.n220 163.367
R555 B.n404 B.n403 163.367
R556 B.n405 B.n404 163.367
R557 B.n405 B.n218 163.367
R558 B.n409 B.n218 163.367
R559 B.n410 B.n409 163.367
R560 B.n411 B.n410 163.367
R561 B.n411 B.n216 163.367
R562 B.n415 B.n216 163.367
R563 B.n416 B.n415 163.367
R564 B.n417 B.n416 163.367
R565 B.n417 B.n214 163.367
R566 B.n421 B.n214 163.367
R567 B.n422 B.n421 163.367
R568 B.n423 B.n422 163.367
R569 B.n423 B.n212 163.367
R570 B.n427 B.n212 163.367
R571 B.n428 B.n427 163.367
R572 B.n429 B.n428 163.367
R573 B.n429 B.n210 163.367
R574 B.n433 B.n210 163.367
R575 B.n434 B.n433 163.367
R576 B.n435 B.n434 163.367
R577 B.n435 B.n208 163.367
R578 B.n439 B.n208 163.367
R579 B.n440 B.n439 163.367
R580 B.n441 B.n440 163.367
R581 B.n441 B.n206 163.367
R582 B.n445 B.n206 163.367
R583 B.n446 B.n445 163.367
R584 B.n447 B.n446 163.367
R585 B.n447 B.n202 163.367
R586 B.n452 B.n202 163.367
R587 B.n453 B.n452 163.367
R588 B.n454 B.n453 163.367
R589 B.n454 B.n200 163.367
R590 B.n458 B.n200 163.367
R591 B.n459 B.n458 163.367
R592 B.n460 B.n459 163.367
R593 B.n460 B.n198 163.367
R594 B.n467 B.n198 163.367
R595 B.n468 B.n467 163.367
R596 B.n469 B.n468 163.367
R597 B.n469 B.n196 163.367
R598 B.n473 B.n196 163.367
R599 B.n474 B.n473 163.367
R600 B.n475 B.n474 163.367
R601 B.n475 B.n194 163.367
R602 B.n479 B.n194 163.367
R603 B.n480 B.n479 163.367
R604 B.n481 B.n480 163.367
R605 B.n481 B.n192 163.367
R606 B.n485 B.n192 163.367
R607 B.n486 B.n485 163.367
R608 B.n487 B.n486 163.367
R609 B.n487 B.n190 163.367
R610 B.n491 B.n190 163.367
R611 B.n492 B.n491 163.367
R612 B.n493 B.n492 163.367
R613 B.n493 B.n188 163.367
R614 B.n497 B.n188 163.367
R615 B.n498 B.n497 163.367
R616 B.n499 B.n498 163.367
R617 B.n499 B.n186 163.367
R618 B.n503 B.n186 163.367
R619 B.n504 B.n503 163.367
R620 B.n505 B.n504 163.367
R621 B.n505 B.n184 163.367
R622 B.n509 B.n184 163.367
R623 B.n510 B.n509 163.367
R624 B.n511 B.n510 163.367
R625 B.n511 B.n182 163.367
R626 B.n515 B.n182 163.367
R627 B.n516 B.n515 163.367
R628 B.n517 B.n516 163.367
R629 B.n517 B.n180 163.367
R630 B.n521 B.n180 163.367
R631 B.n522 B.n521 163.367
R632 B.n523 B.n522 163.367
R633 B.n523 B.n178 163.367
R634 B.n527 B.n178 163.367
R635 B.n528 B.n527 163.367
R636 B.n529 B.n528 163.367
R637 B.n529 B.n176 163.367
R638 B.n533 B.n176 163.367
R639 B.n534 B.n533 163.367
R640 B.n535 B.n534 163.367
R641 B.n535 B.n174 163.367
R642 B.n539 B.n174 163.367
R643 B.n540 B.n539 163.367
R644 B.n541 B.n540 163.367
R645 B.n541 B.n172 163.367
R646 B.n545 B.n172 163.367
R647 B.n546 B.n545 163.367
R648 B.n547 B.n546 163.367
R649 B.n547 B.n170 163.367
R650 B.n551 B.n170 163.367
R651 B.n552 B.n551 163.367
R652 B.n751 B.n102 163.367
R653 B.n751 B.n750 163.367
R654 B.n750 B.n749 163.367
R655 B.n749 B.n104 163.367
R656 B.n745 B.n104 163.367
R657 B.n745 B.n744 163.367
R658 B.n744 B.n743 163.367
R659 B.n743 B.n106 163.367
R660 B.n739 B.n106 163.367
R661 B.n739 B.n738 163.367
R662 B.n738 B.n737 163.367
R663 B.n737 B.n108 163.367
R664 B.n733 B.n108 163.367
R665 B.n733 B.n732 163.367
R666 B.n732 B.n731 163.367
R667 B.n731 B.n110 163.367
R668 B.n727 B.n110 163.367
R669 B.n727 B.n726 163.367
R670 B.n726 B.n725 163.367
R671 B.n725 B.n112 163.367
R672 B.n721 B.n112 163.367
R673 B.n721 B.n720 163.367
R674 B.n720 B.n719 163.367
R675 B.n719 B.n114 163.367
R676 B.n715 B.n114 163.367
R677 B.n715 B.n714 163.367
R678 B.n714 B.n713 163.367
R679 B.n713 B.n116 163.367
R680 B.n709 B.n116 163.367
R681 B.n709 B.n708 163.367
R682 B.n708 B.n707 163.367
R683 B.n707 B.n118 163.367
R684 B.n703 B.n118 163.367
R685 B.n703 B.n702 163.367
R686 B.n702 B.n701 163.367
R687 B.n701 B.n120 163.367
R688 B.n697 B.n120 163.367
R689 B.n697 B.n696 163.367
R690 B.n696 B.n695 163.367
R691 B.n695 B.n122 163.367
R692 B.n691 B.n122 163.367
R693 B.n691 B.n690 163.367
R694 B.n690 B.n689 163.367
R695 B.n689 B.n124 163.367
R696 B.n685 B.n124 163.367
R697 B.n685 B.n684 163.367
R698 B.n684 B.n683 163.367
R699 B.n683 B.n126 163.367
R700 B.n679 B.n126 163.367
R701 B.n679 B.n678 163.367
R702 B.n678 B.n677 163.367
R703 B.n677 B.n128 163.367
R704 B.n673 B.n128 163.367
R705 B.n673 B.n672 163.367
R706 B.n672 B.n671 163.367
R707 B.n671 B.n130 163.367
R708 B.n667 B.n130 163.367
R709 B.n667 B.n666 163.367
R710 B.n666 B.n665 163.367
R711 B.n665 B.n132 163.367
R712 B.n661 B.n132 163.367
R713 B.n661 B.n660 163.367
R714 B.n660 B.n659 163.367
R715 B.n659 B.n134 163.367
R716 B.n655 B.n134 163.367
R717 B.n655 B.n654 163.367
R718 B.n654 B.n653 163.367
R719 B.n653 B.n136 163.367
R720 B.n649 B.n136 163.367
R721 B.n649 B.n648 163.367
R722 B.n648 B.n647 163.367
R723 B.n647 B.n138 163.367
R724 B.n643 B.n138 163.367
R725 B.n643 B.n642 163.367
R726 B.n642 B.n641 163.367
R727 B.n641 B.n140 163.367
R728 B.n637 B.n140 163.367
R729 B.n637 B.n636 163.367
R730 B.n636 B.n635 163.367
R731 B.n635 B.n142 163.367
R732 B.n631 B.n142 163.367
R733 B.n631 B.n630 163.367
R734 B.n630 B.n629 163.367
R735 B.n629 B.n144 163.367
R736 B.n625 B.n144 163.367
R737 B.n625 B.n624 163.367
R738 B.n624 B.n623 163.367
R739 B.n623 B.n146 163.367
R740 B.n619 B.n146 163.367
R741 B.n619 B.n618 163.367
R742 B.n618 B.n617 163.367
R743 B.n617 B.n148 163.367
R744 B.n613 B.n148 163.367
R745 B.n613 B.n612 163.367
R746 B.n612 B.n611 163.367
R747 B.n611 B.n150 163.367
R748 B.n607 B.n150 163.367
R749 B.n607 B.n606 163.367
R750 B.n606 B.n605 163.367
R751 B.n605 B.n152 163.367
R752 B.n601 B.n152 163.367
R753 B.n601 B.n600 163.367
R754 B.n600 B.n599 163.367
R755 B.n599 B.n154 163.367
R756 B.n595 B.n154 163.367
R757 B.n595 B.n594 163.367
R758 B.n594 B.n593 163.367
R759 B.n593 B.n156 163.367
R760 B.n589 B.n156 163.367
R761 B.n589 B.n588 163.367
R762 B.n588 B.n587 163.367
R763 B.n587 B.n158 163.367
R764 B.n583 B.n158 163.367
R765 B.n583 B.n582 163.367
R766 B.n582 B.n581 163.367
R767 B.n581 B.n160 163.367
R768 B.n577 B.n160 163.367
R769 B.n577 B.n576 163.367
R770 B.n576 B.n575 163.367
R771 B.n575 B.n162 163.367
R772 B.n571 B.n162 163.367
R773 B.n571 B.n570 163.367
R774 B.n570 B.n569 163.367
R775 B.n569 B.n164 163.367
R776 B.n565 B.n164 163.367
R777 B.n565 B.n564 163.367
R778 B.n564 B.n563 163.367
R779 B.n563 B.n166 163.367
R780 B.n559 B.n166 163.367
R781 B.n559 B.n558 163.367
R782 B.n558 B.n557 163.367
R783 B.n557 B.n168 163.367
R784 B.n553 B.n168 163.367
R785 B.n938 B.n35 163.367
R786 B.n938 B.n937 163.367
R787 B.n937 B.n936 163.367
R788 B.n936 B.n37 163.367
R789 B.n932 B.n37 163.367
R790 B.n932 B.n931 163.367
R791 B.n931 B.n930 163.367
R792 B.n930 B.n39 163.367
R793 B.n926 B.n39 163.367
R794 B.n926 B.n925 163.367
R795 B.n925 B.n924 163.367
R796 B.n924 B.n41 163.367
R797 B.n920 B.n41 163.367
R798 B.n920 B.n919 163.367
R799 B.n919 B.n918 163.367
R800 B.n918 B.n43 163.367
R801 B.n914 B.n43 163.367
R802 B.n914 B.n913 163.367
R803 B.n913 B.n912 163.367
R804 B.n912 B.n45 163.367
R805 B.n908 B.n45 163.367
R806 B.n908 B.n907 163.367
R807 B.n907 B.n906 163.367
R808 B.n906 B.n47 163.367
R809 B.n902 B.n47 163.367
R810 B.n902 B.n901 163.367
R811 B.n901 B.n900 163.367
R812 B.n900 B.n49 163.367
R813 B.n896 B.n49 163.367
R814 B.n896 B.n895 163.367
R815 B.n895 B.n894 163.367
R816 B.n894 B.n51 163.367
R817 B.n890 B.n51 163.367
R818 B.n890 B.n889 163.367
R819 B.n889 B.n888 163.367
R820 B.n888 B.n53 163.367
R821 B.n884 B.n53 163.367
R822 B.n884 B.n883 163.367
R823 B.n883 B.n882 163.367
R824 B.n882 B.n55 163.367
R825 B.n878 B.n55 163.367
R826 B.n878 B.n877 163.367
R827 B.n877 B.n876 163.367
R828 B.n876 B.n57 163.367
R829 B.n872 B.n57 163.367
R830 B.n872 B.n871 163.367
R831 B.n871 B.n870 163.367
R832 B.n870 B.n59 163.367
R833 B.n866 B.n59 163.367
R834 B.n866 B.n865 163.367
R835 B.n865 B.n864 163.367
R836 B.n864 B.n61 163.367
R837 B.n860 B.n61 163.367
R838 B.n860 B.n859 163.367
R839 B.n859 B.n858 163.367
R840 B.n858 B.n63 163.367
R841 B.n853 B.n63 163.367
R842 B.n853 B.n852 163.367
R843 B.n852 B.n851 163.367
R844 B.n851 B.n67 163.367
R845 B.n847 B.n67 163.367
R846 B.n847 B.n846 163.367
R847 B.n846 B.n845 163.367
R848 B.n845 B.n69 163.367
R849 B.n841 B.n69 163.367
R850 B.n841 B.n840 163.367
R851 B.n840 B.n839 163.367
R852 B.n839 B.n71 163.367
R853 B.n835 B.n71 163.367
R854 B.n835 B.n834 163.367
R855 B.n834 B.n833 163.367
R856 B.n833 B.n76 163.367
R857 B.n829 B.n76 163.367
R858 B.n829 B.n828 163.367
R859 B.n828 B.n827 163.367
R860 B.n827 B.n78 163.367
R861 B.n823 B.n78 163.367
R862 B.n823 B.n822 163.367
R863 B.n822 B.n821 163.367
R864 B.n821 B.n80 163.367
R865 B.n817 B.n80 163.367
R866 B.n817 B.n816 163.367
R867 B.n816 B.n815 163.367
R868 B.n815 B.n82 163.367
R869 B.n811 B.n82 163.367
R870 B.n811 B.n810 163.367
R871 B.n810 B.n809 163.367
R872 B.n809 B.n84 163.367
R873 B.n805 B.n84 163.367
R874 B.n805 B.n804 163.367
R875 B.n804 B.n803 163.367
R876 B.n803 B.n86 163.367
R877 B.n799 B.n86 163.367
R878 B.n799 B.n798 163.367
R879 B.n798 B.n797 163.367
R880 B.n797 B.n88 163.367
R881 B.n793 B.n88 163.367
R882 B.n793 B.n792 163.367
R883 B.n792 B.n791 163.367
R884 B.n791 B.n90 163.367
R885 B.n787 B.n90 163.367
R886 B.n787 B.n786 163.367
R887 B.n786 B.n785 163.367
R888 B.n785 B.n92 163.367
R889 B.n781 B.n92 163.367
R890 B.n781 B.n780 163.367
R891 B.n780 B.n779 163.367
R892 B.n779 B.n94 163.367
R893 B.n775 B.n94 163.367
R894 B.n775 B.n774 163.367
R895 B.n774 B.n773 163.367
R896 B.n773 B.n96 163.367
R897 B.n769 B.n96 163.367
R898 B.n769 B.n768 163.367
R899 B.n768 B.n767 163.367
R900 B.n767 B.n98 163.367
R901 B.n763 B.n98 163.367
R902 B.n763 B.n762 163.367
R903 B.n762 B.n761 163.367
R904 B.n761 B.n100 163.367
R905 B.n757 B.n100 163.367
R906 B.n757 B.n756 163.367
R907 B.n756 B.n755 163.367
R908 B.n943 B.n942 163.367
R909 B.n944 B.n943 163.367
R910 B.n944 B.n33 163.367
R911 B.n948 B.n33 163.367
R912 B.n949 B.n948 163.367
R913 B.n950 B.n949 163.367
R914 B.n950 B.n31 163.367
R915 B.n954 B.n31 163.367
R916 B.n955 B.n954 163.367
R917 B.n956 B.n955 163.367
R918 B.n956 B.n29 163.367
R919 B.n960 B.n29 163.367
R920 B.n961 B.n960 163.367
R921 B.n962 B.n961 163.367
R922 B.n962 B.n27 163.367
R923 B.n966 B.n27 163.367
R924 B.n967 B.n966 163.367
R925 B.n968 B.n967 163.367
R926 B.n968 B.n25 163.367
R927 B.n972 B.n25 163.367
R928 B.n973 B.n972 163.367
R929 B.n974 B.n973 163.367
R930 B.n974 B.n23 163.367
R931 B.n978 B.n23 163.367
R932 B.n979 B.n978 163.367
R933 B.n980 B.n979 163.367
R934 B.n980 B.n21 163.367
R935 B.n984 B.n21 163.367
R936 B.n985 B.n984 163.367
R937 B.n986 B.n985 163.367
R938 B.n986 B.n19 163.367
R939 B.n990 B.n19 163.367
R940 B.n991 B.n990 163.367
R941 B.n992 B.n991 163.367
R942 B.n992 B.n17 163.367
R943 B.n996 B.n17 163.367
R944 B.n997 B.n996 163.367
R945 B.n998 B.n997 163.367
R946 B.n998 B.n15 163.367
R947 B.n1002 B.n15 163.367
R948 B.n1003 B.n1002 163.367
R949 B.n1004 B.n1003 163.367
R950 B.n1004 B.n13 163.367
R951 B.n1008 B.n13 163.367
R952 B.n1009 B.n1008 163.367
R953 B.n1010 B.n1009 163.367
R954 B.n1010 B.n11 163.367
R955 B.n1014 B.n11 163.367
R956 B.n1015 B.n1014 163.367
R957 B.n1016 B.n1015 163.367
R958 B.n1016 B.n9 163.367
R959 B.n1020 B.n9 163.367
R960 B.n1021 B.n1020 163.367
R961 B.n1022 B.n1021 163.367
R962 B.n1022 B.n7 163.367
R963 B.n1026 B.n7 163.367
R964 B.n1027 B.n1026 163.367
R965 B.n1028 B.n1027 163.367
R966 B.n1028 B.n5 163.367
R967 B.n1032 B.n5 163.367
R968 B.n1033 B.n1032 163.367
R969 B.n1034 B.n1033 163.367
R970 B.n1034 B.n3 163.367
R971 B.n1038 B.n3 163.367
R972 B.n1039 B.n1038 163.367
R973 B.n266 B.n2 163.367
R974 B.n267 B.n266 163.367
R975 B.n267 B.n264 163.367
R976 B.n271 B.n264 163.367
R977 B.n272 B.n271 163.367
R978 B.n273 B.n272 163.367
R979 B.n273 B.n262 163.367
R980 B.n277 B.n262 163.367
R981 B.n278 B.n277 163.367
R982 B.n279 B.n278 163.367
R983 B.n279 B.n260 163.367
R984 B.n283 B.n260 163.367
R985 B.n284 B.n283 163.367
R986 B.n285 B.n284 163.367
R987 B.n285 B.n258 163.367
R988 B.n289 B.n258 163.367
R989 B.n290 B.n289 163.367
R990 B.n291 B.n290 163.367
R991 B.n291 B.n256 163.367
R992 B.n295 B.n256 163.367
R993 B.n296 B.n295 163.367
R994 B.n297 B.n296 163.367
R995 B.n297 B.n254 163.367
R996 B.n301 B.n254 163.367
R997 B.n302 B.n301 163.367
R998 B.n303 B.n302 163.367
R999 B.n303 B.n252 163.367
R1000 B.n307 B.n252 163.367
R1001 B.n308 B.n307 163.367
R1002 B.n309 B.n308 163.367
R1003 B.n309 B.n250 163.367
R1004 B.n313 B.n250 163.367
R1005 B.n314 B.n313 163.367
R1006 B.n315 B.n314 163.367
R1007 B.n315 B.n248 163.367
R1008 B.n319 B.n248 163.367
R1009 B.n320 B.n319 163.367
R1010 B.n321 B.n320 163.367
R1011 B.n321 B.n246 163.367
R1012 B.n325 B.n246 163.367
R1013 B.n326 B.n325 163.367
R1014 B.n327 B.n326 163.367
R1015 B.n327 B.n244 163.367
R1016 B.n331 B.n244 163.367
R1017 B.n332 B.n331 163.367
R1018 B.n333 B.n332 163.367
R1019 B.n333 B.n242 163.367
R1020 B.n337 B.n242 163.367
R1021 B.n338 B.n337 163.367
R1022 B.n339 B.n338 163.367
R1023 B.n339 B.n240 163.367
R1024 B.n343 B.n240 163.367
R1025 B.n344 B.n343 163.367
R1026 B.n345 B.n344 163.367
R1027 B.n345 B.n238 163.367
R1028 B.n349 B.n238 163.367
R1029 B.n350 B.n349 163.367
R1030 B.n351 B.n350 163.367
R1031 B.n351 B.n236 163.367
R1032 B.n355 B.n236 163.367
R1033 B.n356 B.n355 163.367
R1034 B.n357 B.n356 163.367
R1035 B.n357 B.n234 163.367
R1036 B.n361 B.n234 163.367
R1037 B.n362 B.n361 163.367
R1038 B.n464 B.t11 111.323
R1039 B.n73 B.t1 111.323
R1040 B.n204 B.t8 111.3
R1041 B.n65 B.t4 111.3
R1042 B.n204 B.n203 64.1944
R1043 B.n464 B.n463 64.1944
R1044 B.n73 B.n72 64.1944
R1045 B.n65 B.n64 64.1944
R1046 B.n449 B.n204 59.5399
R1047 B.n465 B.n464 59.5399
R1048 B.n74 B.n73 59.5399
R1049 B.n855 B.n65 59.5399
R1050 B.n941 B.n940 31.3761
R1051 B.n754 B.n753 31.3761
R1052 B.n554 B.n169 31.3761
R1053 B.n364 B.n233 31.3761
R1054 B B.n1041 18.0485
R1055 B.n941 B.n34 10.6151
R1056 B.n945 B.n34 10.6151
R1057 B.n946 B.n945 10.6151
R1058 B.n947 B.n946 10.6151
R1059 B.n947 B.n32 10.6151
R1060 B.n951 B.n32 10.6151
R1061 B.n952 B.n951 10.6151
R1062 B.n953 B.n952 10.6151
R1063 B.n953 B.n30 10.6151
R1064 B.n957 B.n30 10.6151
R1065 B.n958 B.n957 10.6151
R1066 B.n959 B.n958 10.6151
R1067 B.n959 B.n28 10.6151
R1068 B.n963 B.n28 10.6151
R1069 B.n964 B.n963 10.6151
R1070 B.n965 B.n964 10.6151
R1071 B.n965 B.n26 10.6151
R1072 B.n969 B.n26 10.6151
R1073 B.n970 B.n969 10.6151
R1074 B.n971 B.n970 10.6151
R1075 B.n971 B.n24 10.6151
R1076 B.n975 B.n24 10.6151
R1077 B.n976 B.n975 10.6151
R1078 B.n977 B.n976 10.6151
R1079 B.n977 B.n22 10.6151
R1080 B.n981 B.n22 10.6151
R1081 B.n982 B.n981 10.6151
R1082 B.n983 B.n982 10.6151
R1083 B.n983 B.n20 10.6151
R1084 B.n987 B.n20 10.6151
R1085 B.n988 B.n987 10.6151
R1086 B.n989 B.n988 10.6151
R1087 B.n989 B.n18 10.6151
R1088 B.n993 B.n18 10.6151
R1089 B.n994 B.n993 10.6151
R1090 B.n995 B.n994 10.6151
R1091 B.n995 B.n16 10.6151
R1092 B.n999 B.n16 10.6151
R1093 B.n1000 B.n999 10.6151
R1094 B.n1001 B.n1000 10.6151
R1095 B.n1001 B.n14 10.6151
R1096 B.n1005 B.n14 10.6151
R1097 B.n1006 B.n1005 10.6151
R1098 B.n1007 B.n1006 10.6151
R1099 B.n1007 B.n12 10.6151
R1100 B.n1011 B.n12 10.6151
R1101 B.n1012 B.n1011 10.6151
R1102 B.n1013 B.n1012 10.6151
R1103 B.n1013 B.n10 10.6151
R1104 B.n1017 B.n10 10.6151
R1105 B.n1018 B.n1017 10.6151
R1106 B.n1019 B.n1018 10.6151
R1107 B.n1019 B.n8 10.6151
R1108 B.n1023 B.n8 10.6151
R1109 B.n1024 B.n1023 10.6151
R1110 B.n1025 B.n1024 10.6151
R1111 B.n1025 B.n6 10.6151
R1112 B.n1029 B.n6 10.6151
R1113 B.n1030 B.n1029 10.6151
R1114 B.n1031 B.n1030 10.6151
R1115 B.n1031 B.n4 10.6151
R1116 B.n1035 B.n4 10.6151
R1117 B.n1036 B.n1035 10.6151
R1118 B.n1037 B.n1036 10.6151
R1119 B.n1037 B.n0 10.6151
R1120 B.n940 B.n939 10.6151
R1121 B.n939 B.n36 10.6151
R1122 B.n935 B.n36 10.6151
R1123 B.n935 B.n934 10.6151
R1124 B.n934 B.n933 10.6151
R1125 B.n933 B.n38 10.6151
R1126 B.n929 B.n38 10.6151
R1127 B.n929 B.n928 10.6151
R1128 B.n928 B.n927 10.6151
R1129 B.n927 B.n40 10.6151
R1130 B.n923 B.n40 10.6151
R1131 B.n923 B.n922 10.6151
R1132 B.n922 B.n921 10.6151
R1133 B.n921 B.n42 10.6151
R1134 B.n917 B.n42 10.6151
R1135 B.n917 B.n916 10.6151
R1136 B.n916 B.n915 10.6151
R1137 B.n915 B.n44 10.6151
R1138 B.n911 B.n44 10.6151
R1139 B.n911 B.n910 10.6151
R1140 B.n910 B.n909 10.6151
R1141 B.n909 B.n46 10.6151
R1142 B.n905 B.n46 10.6151
R1143 B.n905 B.n904 10.6151
R1144 B.n904 B.n903 10.6151
R1145 B.n903 B.n48 10.6151
R1146 B.n899 B.n48 10.6151
R1147 B.n899 B.n898 10.6151
R1148 B.n898 B.n897 10.6151
R1149 B.n897 B.n50 10.6151
R1150 B.n893 B.n50 10.6151
R1151 B.n893 B.n892 10.6151
R1152 B.n892 B.n891 10.6151
R1153 B.n891 B.n52 10.6151
R1154 B.n887 B.n52 10.6151
R1155 B.n887 B.n886 10.6151
R1156 B.n886 B.n885 10.6151
R1157 B.n885 B.n54 10.6151
R1158 B.n881 B.n54 10.6151
R1159 B.n881 B.n880 10.6151
R1160 B.n880 B.n879 10.6151
R1161 B.n879 B.n56 10.6151
R1162 B.n875 B.n56 10.6151
R1163 B.n875 B.n874 10.6151
R1164 B.n874 B.n873 10.6151
R1165 B.n873 B.n58 10.6151
R1166 B.n869 B.n58 10.6151
R1167 B.n869 B.n868 10.6151
R1168 B.n868 B.n867 10.6151
R1169 B.n867 B.n60 10.6151
R1170 B.n863 B.n60 10.6151
R1171 B.n863 B.n862 10.6151
R1172 B.n862 B.n861 10.6151
R1173 B.n861 B.n62 10.6151
R1174 B.n857 B.n62 10.6151
R1175 B.n857 B.n856 10.6151
R1176 B.n854 B.n66 10.6151
R1177 B.n850 B.n66 10.6151
R1178 B.n850 B.n849 10.6151
R1179 B.n849 B.n848 10.6151
R1180 B.n848 B.n68 10.6151
R1181 B.n844 B.n68 10.6151
R1182 B.n844 B.n843 10.6151
R1183 B.n843 B.n842 10.6151
R1184 B.n842 B.n70 10.6151
R1185 B.n838 B.n837 10.6151
R1186 B.n837 B.n836 10.6151
R1187 B.n836 B.n75 10.6151
R1188 B.n832 B.n75 10.6151
R1189 B.n832 B.n831 10.6151
R1190 B.n831 B.n830 10.6151
R1191 B.n830 B.n77 10.6151
R1192 B.n826 B.n77 10.6151
R1193 B.n826 B.n825 10.6151
R1194 B.n825 B.n824 10.6151
R1195 B.n824 B.n79 10.6151
R1196 B.n820 B.n79 10.6151
R1197 B.n820 B.n819 10.6151
R1198 B.n819 B.n818 10.6151
R1199 B.n818 B.n81 10.6151
R1200 B.n814 B.n81 10.6151
R1201 B.n814 B.n813 10.6151
R1202 B.n813 B.n812 10.6151
R1203 B.n812 B.n83 10.6151
R1204 B.n808 B.n83 10.6151
R1205 B.n808 B.n807 10.6151
R1206 B.n807 B.n806 10.6151
R1207 B.n806 B.n85 10.6151
R1208 B.n802 B.n85 10.6151
R1209 B.n802 B.n801 10.6151
R1210 B.n801 B.n800 10.6151
R1211 B.n800 B.n87 10.6151
R1212 B.n796 B.n87 10.6151
R1213 B.n796 B.n795 10.6151
R1214 B.n795 B.n794 10.6151
R1215 B.n794 B.n89 10.6151
R1216 B.n790 B.n89 10.6151
R1217 B.n790 B.n789 10.6151
R1218 B.n789 B.n788 10.6151
R1219 B.n788 B.n91 10.6151
R1220 B.n784 B.n91 10.6151
R1221 B.n784 B.n783 10.6151
R1222 B.n783 B.n782 10.6151
R1223 B.n782 B.n93 10.6151
R1224 B.n778 B.n93 10.6151
R1225 B.n778 B.n777 10.6151
R1226 B.n777 B.n776 10.6151
R1227 B.n776 B.n95 10.6151
R1228 B.n772 B.n95 10.6151
R1229 B.n772 B.n771 10.6151
R1230 B.n771 B.n770 10.6151
R1231 B.n770 B.n97 10.6151
R1232 B.n766 B.n97 10.6151
R1233 B.n766 B.n765 10.6151
R1234 B.n765 B.n764 10.6151
R1235 B.n764 B.n99 10.6151
R1236 B.n760 B.n99 10.6151
R1237 B.n760 B.n759 10.6151
R1238 B.n759 B.n758 10.6151
R1239 B.n758 B.n101 10.6151
R1240 B.n754 B.n101 10.6151
R1241 B.n753 B.n752 10.6151
R1242 B.n752 B.n103 10.6151
R1243 B.n748 B.n103 10.6151
R1244 B.n748 B.n747 10.6151
R1245 B.n747 B.n746 10.6151
R1246 B.n746 B.n105 10.6151
R1247 B.n742 B.n105 10.6151
R1248 B.n742 B.n741 10.6151
R1249 B.n741 B.n740 10.6151
R1250 B.n740 B.n107 10.6151
R1251 B.n736 B.n107 10.6151
R1252 B.n736 B.n735 10.6151
R1253 B.n735 B.n734 10.6151
R1254 B.n734 B.n109 10.6151
R1255 B.n730 B.n109 10.6151
R1256 B.n730 B.n729 10.6151
R1257 B.n729 B.n728 10.6151
R1258 B.n728 B.n111 10.6151
R1259 B.n724 B.n111 10.6151
R1260 B.n724 B.n723 10.6151
R1261 B.n723 B.n722 10.6151
R1262 B.n722 B.n113 10.6151
R1263 B.n718 B.n113 10.6151
R1264 B.n718 B.n717 10.6151
R1265 B.n717 B.n716 10.6151
R1266 B.n716 B.n115 10.6151
R1267 B.n712 B.n115 10.6151
R1268 B.n712 B.n711 10.6151
R1269 B.n711 B.n710 10.6151
R1270 B.n710 B.n117 10.6151
R1271 B.n706 B.n117 10.6151
R1272 B.n706 B.n705 10.6151
R1273 B.n705 B.n704 10.6151
R1274 B.n704 B.n119 10.6151
R1275 B.n700 B.n119 10.6151
R1276 B.n700 B.n699 10.6151
R1277 B.n699 B.n698 10.6151
R1278 B.n698 B.n121 10.6151
R1279 B.n694 B.n121 10.6151
R1280 B.n694 B.n693 10.6151
R1281 B.n693 B.n692 10.6151
R1282 B.n692 B.n123 10.6151
R1283 B.n688 B.n123 10.6151
R1284 B.n688 B.n687 10.6151
R1285 B.n687 B.n686 10.6151
R1286 B.n686 B.n125 10.6151
R1287 B.n682 B.n125 10.6151
R1288 B.n682 B.n681 10.6151
R1289 B.n681 B.n680 10.6151
R1290 B.n680 B.n127 10.6151
R1291 B.n676 B.n127 10.6151
R1292 B.n676 B.n675 10.6151
R1293 B.n675 B.n674 10.6151
R1294 B.n674 B.n129 10.6151
R1295 B.n670 B.n129 10.6151
R1296 B.n670 B.n669 10.6151
R1297 B.n669 B.n668 10.6151
R1298 B.n668 B.n131 10.6151
R1299 B.n664 B.n131 10.6151
R1300 B.n664 B.n663 10.6151
R1301 B.n663 B.n662 10.6151
R1302 B.n662 B.n133 10.6151
R1303 B.n658 B.n133 10.6151
R1304 B.n658 B.n657 10.6151
R1305 B.n657 B.n656 10.6151
R1306 B.n656 B.n135 10.6151
R1307 B.n652 B.n135 10.6151
R1308 B.n652 B.n651 10.6151
R1309 B.n651 B.n650 10.6151
R1310 B.n650 B.n137 10.6151
R1311 B.n646 B.n137 10.6151
R1312 B.n646 B.n645 10.6151
R1313 B.n645 B.n644 10.6151
R1314 B.n644 B.n139 10.6151
R1315 B.n640 B.n139 10.6151
R1316 B.n640 B.n639 10.6151
R1317 B.n639 B.n638 10.6151
R1318 B.n638 B.n141 10.6151
R1319 B.n634 B.n141 10.6151
R1320 B.n634 B.n633 10.6151
R1321 B.n633 B.n632 10.6151
R1322 B.n632 B.n143 10.6151
R1323 B.n628 B.n143 10.6151
R1324 B.n628 B.n627 10.6151
R1325 B.n627 B.n626 10.6151
R1326 B.n626 B.n145 10.6151
R1327 B.n622 B.n145 10.6151
R1328 B.n622 B.n621 10.6151
R1329 B.n621 B.n620 10.6151
R1330 B.n620 B.n147 10.6151
R1331 B.n616 B.n147 10.6151
R1332 B.n616 B.n615 10.6151
R1333 B.n615 B.n614 10.6151
R1334 B.n614 B.n149 10.6151
R1335 B.n610 B.n149 10.6151
R1336 B.n610 B.n609 10.6151
R1337 B.n609 B.n608 10.6151
R1338 B.n608 B.n151 10.6151
R1339 B.n604 B.n151 10.6151
R1340 B.n604 B.n603 10.6151
R1341 B.n603 B.n602 10.6151
R1342 B.n602 B.n153 10.6151
R1343 B.n598 B.n153 10.6151
R1344 B.n598 B.n597 10.6151
R1345 B.n597 B.n596 10.6151
R1346 B.n596 B.n155 10.6151
R1347 B.n592 B.n155 10.6151
R1348 B.n592 B.n591 10.6151
R1349 B.n591 B.n590 10.6151
R1350 B.n590 B.n157 10.6151
R1351 B.n586 B.n157 10.6151
R1352 B.n586 B.n585 10.6151
R1353 B.n585 B.n584 10.6151
R1354 B.n584 B.n159 10.6151
R1355 B.n580 B.n159 10.6151
R1356 B.n580 B.n579 10.6151
R1357 B.n579 B.n578 10.6151
R1358 B.n578 B.n161 10.6151
R1359 B.n574 B.n161 10.6151
R1360 B.n574 B.n573 10.6151
R1361 B.n573 B.n572 10.6151
R1362 B.n572 B.n163 10.6151
R1363 B.n568 B.n163 10.6151
R1364 B.n568 B.n567 10.6151
R1365 B.n567 B.n566 10.6151
R1366 B.n566 B.n165 10.6151
R1367 B.n562 B.n165 10.6151
R1368 B.n562 B.n561 10.6151
R1369 B.n561 B.n560 10.6151
R1370 B.n560 B.n167 10.6151
R1371 B.n556 B.n167 10.6151
R1372 B.n556 B.n555 10.6151
R1373 B.n555 B.n554 10.6151
R1374 B.n265 B.n1 10.6151
R1375 B.n268 B.n265 10.6151
R1376 B.n269 B.n268 10.6151
R1377 B.n270 B.n269 10.6151
R1378 B.n270 B.n263 10.6151
R1379 B.n274 B.n263 10.6151
R1380 B.n275 B.n274 10.6151
R1381 B.n276 B.n275 10.6151
R1382 B.n276 B.n261 10.6151
R1383 B.n280 B.n261 10.6151
R1384 B.n281 B.n280 10.6151
R1385 B.n282 B.n281 10.6151
R1386 B.n282 B.n259 10.6151
R1387 B.n286 B.n259 10.6151
R1388 B.n287 B.n286 10.6151
R1389 B.n288 B.n287 10.6151
R1390 B.n288 B.n257 10.6151
R1391 B.n292 B.n257 10.6151
R1392 B.n293 B.n292 10.6151
R1393 B.n294 B.n293 10.6151
R1394 B.n294 B.n255 10.6151
R1395 B.n298 B.n255 10.6151
R1396 B.n299 B.n298 10.6151
R1397 B.n300 B.n299 10.6151
R1398 B.n300 B.n253 10.6151
R1399 B.n304 B.n253 10.6151
R1400 B.n305 B.n304 10.6151
R1401 B.n306 B.n305 10.6151
R1402 B.n306 B.n251 10.6151
R1403 B.n310 B.n251 10.6151
R1404 B.n311 B.n310 10.6151
R1405 B.n312 B.n311 10.6151
R1406 B.n312 B.n249 10.6151
R1407 B.n316 B.n249 10.6151
R1408 B.n317 B.n316 10.6151
R1409 B.n318 B.n317 10.6151
R1410 B.n318 B.n247 10.6151
R1411 B.n322 B.n247 10.6151
R1412 B.n323 B.n322 10.6151
R1413 B.n324 B.n323 10.6151
R1414 B.n324 B.n245 10.6151
R1415 B.n328 B.n245 10.6151
R1416 B.n329 B.n328 10.6151
R1417 B.n330 B.n329 10.6151
R1418 B.n330 B.n243 10.6151
R1419 B.n334 B.n243 10.6151
R1420 B.n335 B.n334 10.6151
R1421 B.n336 B.n335 10.6151
R1422 B.n336 B.n241 10.6151
R1423 B.n340 B.n241 10.6151
R1424 B.n341 B.n340 10.6151
R1425 B.n342 B.n341 10.6151
R1426 B.n342 B.n239 10.6151
R1427 B.n346 B.n239 10.6151
R1428 B.n347 B.n346 10.6151
R1429 B.n348 B.n347 10.6151
R1430 B.n348 B.n237 10.6151
R1431 B.n352 B.n237 10.6151
R1432 B.n353 B.n352 10.6151
R1433 B.n354 B.n353 10.6151
R1434 B.n354 B.n235 10.6151
R1435 B.n358 B.n235 10.6151
R1436 B.n359 B.n358 10.6151
R1437 B.n360 B.n359 10.6151
R1438 B.n360 B.n233 10.6151
R1439 B.n365 B.n364 10.6151
R1440 B.n366 B.n365 10.6151
R1441 B.n366 B.n231 10.6151
R1442 B.n370 B.n231 10.6151
R1443 B.n371 B.n370 10.6151
R1444 B.n372 B.n371 10.6151
R1445 B.n372 B.n229 10.6151
R1446 B.n376 B.n229 10.6151
R1447 B.n377 B.n376 10.6151
R1448 B.n378 B.n377 10.6151
R1449 B.n378 B.n227 10.6151
R1450 B.n382 B.n227 10.6151
R1451 B.n383 B.n382 10.6151
R1452 B.n384 B.n383 10.6151
R1453 B.n384 B.n225 10.6151
R1454 B.n388 B.n225 10.6151
R1455 B.n389 B.n388 10.6151
R1456 B.n390 B.n389 10.6151
R1457 B.n390 B.n223 10.6151
R1458 B.n394 B.n223 10.6151
R1459 B.n395 B.n394 10.6151
R1460 B.n396 B.n395 10.6151
R1461 B.n396 B.n221 10.6151
R1462 B.n400 B.n221 10.6151
R1463 B.n401 B.n400 10.6151
R1464 B.n402 B.n401 10.6151
R1465 B.n402 B.n219 10.6151
R1466 B.n406 B.n219 10.6151
R1467 B.n407 B.n406 10.6151
R1468 B.n408 B.n407 10.6151
R1469 B.n408 B.n217 10.6151
R1470 B.n412 B.n217 10.6151
R1471 B.n413 B.n412 10.6151
R1472 B.n414 B.n413 10.6151
R1473 B.n414 B.n215 10.6151
R1474 B.n418 B.n215 10.6151
R1475 B.n419 B.n418 10.6151
R1476 B.n420 B.n419 10.6151
R1477 B.n420 B.n213 10.6151
R1478 B.n424 B.n213 10.6151
R1479 B.n425 B.n424 10.6151
R1480 B.n426 B.n425 10.6151
R1481 B.n426 B.n211 10.6151
R1482 B.n430 B.n211 10.6151
R1483 B.n431 B.n430 10.6151
R1484 B.n432 B.n431 10.6151
R1485 B.n432 B.n209 10.6151
R1486 B.n436 B.n209 10.6151
R1487 B.n437 B.n436 10.6151
R1488 B.n438 B.n437 10.6151
R1489 B.n438 B.n207 10.6151
R1490 B.n442 B.n207 10.6151
R1491 B.n443 B.n442 10.6151
R1492 B.n444 B.n443 10.6151
R1493 B.n444 B.n205 10.6151
R1494 B.n448 B.n205 10.6151
R1495 B.n451 B.n450 10.6151
R1496 B.n451 B.n201 10.6151
R1497 B.n455 B.n201 10.6151
R1498 B.n456 B.n455 10.6151
R1499 B.n457 B.n456 10.6151
R1500 B.n457 B.n199 10.6151
R1501 B.n461 B.n199 10.6151
R1502 B.n462 B.n461 10.6151
R1503 B.n466 B.n462 10.6151
R1504 B.n470 B.n197 10.6151
R1505 B.n471 B.n470 10.6151
R1506 B.n472 B.n471 10.6151
R1507 B.n472 B.n195 10.6151
R1508 B.n476 B.n195 10.6151
R1509 B.n477 B.n476 10.6151
R1510 B.n478 B.n477 10.6151
R1511 B.n478 B.n193 10.6151
R1512 B.n482 B.n193 10.6151
R1513 B.n483 B.n482 10.6151
R1514 B.n484 B.n483 10.6151
R1515 B.n484 B.n191 10.6151
R1516 B.n488 B.n191 10.6151
R1517 B.n489 B.n488 10.6151
R1518 B.n490 B.n489 10.6151
R1519 B.n490 B.n189 10.6151
R1520 B.n494 B.n189 10.6151
R1521 B.n495 B.n494 10.6151
R1522 B.n496 B.n495 10.6151
R1523 B.n496 B.n187 10.6151
R1524 B.n500 B.n187 10.6151
R1525 B.n501 B.n500 10.6151
R1526 B.n502 B.n501 10.6151
R1527 B.n502 B.n185 10.6151
R1528 B.n506 B.n185 10.6151
R1529 B.n507 B.n506 10.6151
R1530 B.n508 B.n507 10.6151
R1531 B.n508 B.n183 10.6151
R1532 B.n512 B.n183 10.6151
R1533 B.n513 B.n512 10.6151
R1534 B.n514 B.n513 10.6151
R1535 B.n514 B.n181 10.6151
R1536 B.n518 B.n181 10.6151
R1537 B.n519 B.n518 10.6151
R1538 B.n520 B.n519 10.6151
R1539 B.n520 B.n179 10.6151
R1540 B.n524 B.n179 10.6151
R1541 B.n525 B.n524 10.6151
R1542 B.n526 B.n525 10.6151
R1543 B.n526 B.n177 10.6151
R1544 B.n530 B.n177 10.6151
R1545 B.n531 B.n530 10.6151
R1546 B.n532 B.n531 10.6151
R1547 B.n532 B.n175 10.6151
R1548 B.n536 B.n175 10.6151
R1549 B.n537 B.n536 10.6151
R1550 B.n538 B.n537 10.6151
R1551 B.n538 B.n173 10.6151
R1552 B.n542 B.n173 10.6151
R1553 B.n543 B.n542 10.6151
R1554 B.n544 B.n543 10.6151
R1555 B.n544 B.n171 10.6151
R1556 B.n548 B.n171 10.6151
R1557 B.n549 B.n548 10.6151
R1558 B.n550 B.n549 10.6151
R1559 B.n550 B.n169 10.6151
R1560 B.n856 B.n855 9.36635
R1561 B.n838 B.n74 9.36635
R1562 B.n449 B.n448 9.36635
R1563 B.n465 B.n197 9.36635
R1564 B.n1041 B.n0 8.11757
R1565 B.n1041 B.n1 8.11757
R1566 B.n855 B.n854 1.24928
R1567 B.n74 B.n70 1.24928
R1568 B.n450 B.n449 1.24928
R1569 B.n466 B.n465 1.24928
R1570 VP.n26 VP.t9 171.1
R1571 VP.n27 VP.n24 161.3
R1572 VP.n29 VP.n28 161.3
R1573 VP.n30 VP.n23 161.3
R1574 VP.n32 VP.n31 161.3
R1575 VP.n33 VP.n22 161.3
R1576 VP.n35 VP.n34 161.3
R1577 VP.n36 VP.n21 161.3
R1578 VP.n39 VP.n38 161.3
R1579 VP.n40 VP.n20 161.3
R1580 VP.n42 VP.n41 161.3
R1581 VP.n43 VP.n19 161.3
R1582 VP.n45 VP.n44 161.3
R1583 VP.n46 VP.n18 161.3
R1584 VP.n48 VP.n47 161.3
R1585 VP.n50 VP.n17 161.3
R1586 VP.n52 VP.n51 161.3
R1587 VP.n53 VP.n16 161.3
R1588 VP.n55 VP.n54 161.3
R1589 VP.n56 VP.n15 161.3
R1590 VP.n58 VP.n57 161.3
R1591 VP.n103 VP.n102 161.3
R1592 VP.n101 VP.n1 161.3
R1593 VP.n100 VP.n99 161.3
R1594 VP.n98 VP.n2 161.3
R1595 VP.n97 VP.n96 161.3
R1596 VP.n95 VP.n3 161.3
R1597 VP.n93 VP.n92 161.3
R1598 VP.n91 VP.n4 161.3
R1599 VP.n90 VP.n89 161.3
R1600 VP.n88 VP.n5 161.3
R1601 VP.n87 VP.n86 161.3
R1602 VP.n85 VP.n6 161.3
R1603 VP.n84 VP.n83 161.3
R1604 VP.n81 VP.n7 161.3
R1605 VP.n80 VP.n79 161.3
R1606 VP.n78 VP.n8 161.3
R1607 VP.n77 VP.n76 161.3
R1608 VP.n75 VP.n9 161.3
R1609 VP.n74 VP.n73 161.3
R1610 VP.n72 VP.n10 161.3
R1611 VP.n71 VP.n70 161.3
R1612 VP.n68 VP.n11 161.3
R1613 VP.n67 VP.n66 161.3
R1614 VP.n65 VP.n12 161.3
R1615 VP.n64 VP.n63 161.3
R1616 VP.n62 VP.n13 161.3
R1617 VP.n61 VP.t3 139.587
R1618 VP.n69 VP.t1 139.587
R1619 VP.n82 VP.t4 139.587
R1620 VP.n94 VP.t2 139.587
R1621 VP.n0 VP.t5 139.587
R1622 VP.n14 VP.t8 139.587
R1623 VP.n49 VP.t0 139.587
R1624 VP.n37 VP.t6 139.587
R1625 VP.n25 VP.t7 139.587
R1626 VP.n61 VP.n60 71.8769
R1627 VP.n104 VP.n0 71.8769
R1628 VP.n59 VP.n14 71.8769
R1629 VP.n26 VP.n25 70.3732
R1630 VP.n60 VP.n59 59.2529
R1631 VP.n67 VP.n12 56.4773
R1632 VP.n100 VP.n2 56.4773
R1633 VP.n55 VP.n16 56.4773
R1634 VP.n76 VP.n8 49.6611
R1635 VP.n88 VP.n87 49.6611
R1636 VP.n43 VP.n42 49.6611
R1637 VP.n31 VP.n22 49.6611
R1638 VP.n76 VP.n75 31.1601
R1639 VP.n89 VP.n88 31.1601
R1640 VP.n44 VP.n43 31.1601
R1641 VP.n31 VP.n30 31.1601
R1642 VP.n63 VP.n62 24.3439
R1643 VP.n63 VP.n12 24.3439
R1644 VP.n68 VP.n67 24.3439
R1645 VP.n70 VP.n68 24.3439
R1646 VP.n74 VP.n10 24.3439
R1647 VP.n75 VP.n74 24.3439
R1648 VP.n80 VP.n8 24.3439
R1649 VP.n81 VP.n80 24.3439
R1650 VP.n83 VP.n6 24.3439
R1651 VP.n87 VP.n6 24.3439
R1652 VP.n89 VP.n4 24.3439
R1653 VP.n93 VP.n4 24.3439
R1654 VP.n96 VP.n95 24.3439
R1655 VP.n96 VP.n2 24.3439
R1656 VP.n101 VP.n100 24.3439
R1657 VP.n102 VP.n101 24.3439
R1658 VP.n56 VP.n55 24.3439
R1659 VP.n57 VP.n56 24.3439
R1660 VP.n44 VP.n18 24.3439
R1661 VP.n48 VP.n18 24.3439
R1662 VP.n51 VP.n50 24.3439
R1663 VP.n51 VP.n16 24.3439
R1664 VP.n35 VP.n22 24.3439
R1665 VP.n36 VP.n35 24.3439
R1666 VP.n38 VP.n20 24.3439
R1667 VP.n42 VP.n20 24.3439
R1668 VP.n29 VP.n24 24.3439
R1669 VP.n30 VP.n29 24.3439
R1670 VP.n70 VP.n69 21.4227
R1671 VP.n95 VP.n94 21.4227
R1672 VP.n50 VP.n49 21.4227
R1673 VP.n62 VP.n61 18.0146
R1674 VP.n102 VP.n0 18.0146
R1675 VP.n57 VP.n14 18.0146
R1676 VP.n82 VP.n81 12.1722
R1677 VP.n83 VP.n82 12.1722
R1678 VP.n37 VP.n36 12.1722
R1679 VP.n38 VP.n37 12.1722
R1680 VP.n27 VP.n26 5.7067
R1681 VP.n69 VP.n10 2.92171
R1682 VP.n94 VP.n93 2.92171
R1683 VP.n49 VP.n48 2.92171
R1684 VP.n25 VP.n24 2.92171
R1685 VP.n59 VP.n58 0.355081
R1686 VP.n60 VP.n13 0.355081
R1687 VP.n104 VP.n103 0.355081
R1688 VP VP.n104 0.26685
R1689 VP.n28 VP.n27 0.189894
R1690 VP.n28 VP.n23 0.189894
R1691 VP.n32 VP.n23 0.189894
R1692 VP.n33 VP.n32 0.189894
R1693 VP.n34 VP.n33 0.189894
R1694 VP.n34 VP.n21 0.189894
R1695 VP.n39 VP.n21 0.189894
R1696 VP.n40 VP.n39 0.189894
R1697 VP.n41 VP.n40 0.189894
R1698 VP.n41 VP.n19 0.189894
R1699 VP.n45 VP.n19 0.189894
R1700 VP.n46 VP.n45 0.189894
R1701 VP.n47 VP.n46 0.189894
R1702 VP.n47 VP.n17 0.189894
R1703 VP.n52 VP.n17 0.189894
R1704 VP.n53 VP.n52 0.189894
R1705 VP.n54 VP.n53 0.189894
R1706 VP.n54 VP.n15 0.189894
R1707 VP.n58 VP.n15 0.189894
R1708 VP.n64 VP.n13 0.189894
R1709 VP.n65 VP.n64 0.189894
R1710 VP.n66 VP.n65 0.189894
R1711 VP.n66 VP.n11 0.189894
R1712 VP.n71 VP.n11 0.189894
R1713 VP.n72 VP.n71 0.189894
R1714 VP.n73 VP.n72 0.189894
R1715 VP.n73 VP.n9 0.189894
R1716 VP.n77 VP.n9 0.189894
R1717 VP.n78 VP.n77 0.189894
R1718 VP.n79 VP.n78 0.189894
R1719 VP.n79 VP.n7 0.189894
R1720 VP.n84 VP.n7 0.189894
R1721 VP.n85 VP.n84 0.189894
R1722 VP.n86 VP.n85 0.189894
R1723 VP.n86 VP.n5 0.189894
R1724 VP.n90 VP.n5 0.189894
R1725 VP.n91 VP.n90 0.189894
R1726 VP.n92 VP.n91 0.189894
R1727 VP.n92 VP.n3 0.189894
R1728 VP.n97 VP.n3 0.189894
R1729 VP.n98 VP.n97 0.189894
R1730 VP.n99 VP.n98 0.189894
R1731 VP.n99 VP.n1 0.189894
R1732 VP.n103 VP.n1 0.189894
R1733 VDD1.n1 VDD1.t2 75.8782
R1734 VDD1.n3 VDD1.t1 75.8781
R1735 VDD1.n5 VDD1.n4 73.2261
R1736 VDD1.n1 VDD1.n0 71.1416
R1737 VDD1.n7 VDD1.n6 71.1414
R1738 VDD1.n3 VDD1.n2 71.1413
R1739 VDD1.n7 VDD1.n5 54.1582
R1740 VDD1 VDD1.n7 2.0824
R1741 VDD1.n6 VDD1.t8 1.88376
R1742 VDD1.n6 VDD1.t5 1.88376
R1743 VDD1.n0 VDD1.t0 1.88376
R1744 VDD1.n0 VDD1.t4 1.88376
R1745 VDD1.n4 VDD1.t6 1.88376
R1746 VDD1.n4 VDD1.t3 1.88376
R1747 VDD1.n2 VDD1.t7 1.88376
R1748 VDD1.n2 VDD1.t9 1.88376
R1749 VDD1 VDD1.n1 0.772052
R1750 VDD1.n5 VDD1.n3 0.658516
R1751 VTAIL.n11 VTAIL.t8 56.346
R1752 VTAIL.n17 VTAIL.t6 56.3459
R1753 VTAIL.n2 VTAIL.t14 56.3459
R1754 VTAIL.n16 VTAIL.t11 56.3459
R1755 VTAIL.n15 VTAIL.n14 54.4628
R1756 VTAIL.n13 VTAIL.n12 54.4628
R1757 VTAIL.n10 VTAIL.n9 54.4628
R1758 VTAIL.n8 VTAIL.n7 54.4628
R1759 VTAIL.n19 VTAIL.n18 54.4625
R1760 VTAIL.n1 VTAIL.n0 54.4625
R1761 VTAIL.n4 VTAIL.n3 54.4625
R1762 VTAIL.n6 VTAIL.n5 54.4625
R1763 VTAIL.n8 VTAIL.n6 32.9531
R1764 VTAIL.n17 VTAIL.n16 30.0996
R1765 VTAIL.n10 VTAIL.n8 2.85395
R1766 VTAIL.n11 VTAIL.n10 2.85395
R1767 VTAIL.n15 VTAIL.n13 2.85395
R1768 VTAIL.n16 VTAIL.n15 2.85395
R1769 VTAIL.n6 VTAIL.n4 2.85395
R1770 VTAIL.n4 VTAIL.n2 2.85395
R1771 VTAIL.n19 VTAIL.n17 2.85395
R1772 VTAIL VTAIL.n1 2.19878
R1773 VTAIL.n13 VTAIL.n11 1.89705
R1774 VTAIL.n2 VTAIL.n1 1.89705
R1775 VTAIL.n18 VTAIL.t7 1.88376
R1776 VTAIL.n18 VTAIL.t1 1.88376
R1777 VTAIL.n0 VTAIL.t9 1.88376
R1778 VTAIL.n0 VTAIL.t0 1.88376
R1779 VTAIL.n3 VTAIL.t15 1.88376
R1780 VTAIL.n3 VTAIL.t17 1.88376
R1781 VTAIL.n5 VTAIL.t16 1.88376
R1782 VTAIL.n5 VTAIL.t18 1.88376
R1783 VTAIL.n14 VTAIL.t13 1.88376
R1784 VTAIL.n14 VTAIL.t19 1.88376
R1785 VTAIL.n12 VTAIL.t10 1.88376
R1786 VTAIL.n12 VTAIL.t12 1.88376
R1787 VTAIL.n9 VTAIL.t4 1.88376
R1788 VTAIL.n9 VTAIL.t5 1.88376
R1789 VTAIL.n7 VTAIL.t2 1.88376
R1790 VTAIL.n7 VTAIL.t3 1.88376
R1791 VTAIL VTAIL.n19 0.655672
R1792 VN.n58 VN.t2 171.1
R1793 VN.n12 VN.t6 171.1
R1794 VN.n90 VN.n89 161.3
R1795 VN.n88 VN.n47 161.3
R1796 VN.n87 VN.n86 161.3
R1797 VN.n85 VN.n48 161.3
R1798 VN.n84 VN.n83 161.3
R1799 VN.n82 VN.n49 161.3
R1800 VN.n80 VN.n79 161.3
R1801 VN.n78 VN.n50 161.3
R1802 VN.n77 VN.n76 161.3
R1803 VN.n75 VN.n51 161.3
R1804 VN.n74 VN.n73 161.3
R1805 VN.n72 VN.n52 161.3
R1806 VN.n71 VN.n70 161.3
R1807 VN.n68 VN.n53 161.3
R1808 VN.n67 VN.n66 161.3
R1809 VN.n65 VN.n54 161.3
R1810 VN.n64 VN.n63 161.3
R1811 VN.n62 VN.n55 161.3
R1812 VN.n61 VN.n60 161.3
R1813 VN.n59 VN.n56 161.3
R1814 VN.n44 VN.n43 161.3
R1815 VN.n42 VN.n1 161.3
R1816 VN.n41 VN.n40 161.3
R1817 VN.n39 VN.n2 161.3
R1818 VN.n38 VN.n37 161.3
R1819 VN.n36 VN.n3 161.3
R1820 VN.n34 VN.n33 161.3
R1821 VN.n32 VN.n4 161.3
R1822 VN.n31 VN.n30 161.3
R1823 VN.n29 VN.n5 161.3
R1824 VN.n28 VN.n27 161.3
R1825 VN.n26 VN.n6 161.3
R1826 VN.n25 VN.n24 161.3
R1827 VN.n22 VN.n7 161.3
R1828 VN.n21 VN.n20 161.3
R1829 VN.n19 VN.n8 161.3
R1830 VN.n18 VN.n17 161.3
R1831 VN.n16 VN.n9 161.3
R1832 VN.n15 VN.n14 161.3
R1833 VN.n13 VN.n10 161.3
R1834 VN.n11 VN.t0 139.587
R1835 VN.n23 VN.t3 139.587
R1836 VN.n35 VN.t1 139.587
R1837 VN.n0 VN.t4 139.587
R1838 VN.n57 VN.t5 139.587
R1839 VN.n69 VN.t7 139.587
R1840 VN.n81 VN.t8 139.587
R1841 VN.n46 VN.t9 139.587
R1842 VN.n45 VN.n0 71.8769
R1843 VN.n91 VN.n46 71.8769
R1844 VN.n12 VN.n11 70.3732
R1845 VN.n58 VN.n57 70.3732
R1846 VN VN.n91 59.4184
R1847 VN.n41 VN.n2 56.4773
R1848 VN.n87 VN.n48 56.4773
R1849 VN.n17 VN.n8 49.6611
R1850 VN.n29 VN.n28 49.6611
R1851 VN.n63 VN.n54 49.6611
R1852 VN.n75 VN.n74 49.6611
R1853 VN.n17 VN.n16 31.1601
R1854 VN.n30 VN.n29 31.1601
R1855 VN.n63 VN.n62 31.1601
R1856 VN.n76 VN.n75 31.1601
R1857 VN.n15 VN.n10 24.3439
R1858 VN.n16 VN.n15 24.3439
R1859 VN.n21 VN.n8 24.3439
R1860 VN.n22 VN.n21 24.3439
R1861 VN.n24 VN.n6 24.3439
R1862 VN.n28 VN.n6 24.3439
R1863 VN.n30 VN.n4 24.3439
R1864 VN.n34 VN.n4 24.3439
R1865 VN.n37 VN.n36 24.3439
R1866 VN.n37 VN.n2 24.3439
R1867 VN.n42 VN.n41 24.3439
R1868 VN.n43 VN.n42 24.3439
R1869 VN.n62 VN.n61 24.3439
R1870 VN.n61 VN.n56 24.3439
R1871 VN.n74 VN.n52 24.3439
R1872 VN.n70 VN.n52 24.3439
R1873 VN.n68 VN.n67 24.3439
R1874 VN.n67 VN.n54 24.3439
R1875 VN.n83 VN.n48 24.3439
R1876 VN.n83 VN.n82 24.3439
R1877 VN.n80 VN.n50 24.3439
R1878 VN.n76 VN.n50 24.3439
R1879 VN.n89 VN.n88 24.3439
R1880 VN.n88 VN.n87 24.3439
R1881 VN.n36 VN.n35 21.4227
R1882 VN.n82 VN.n81 21.4227
R1883 VN.n43 VN.n0 18.0146
R1884 VN.n89 VN.n46 18.0146
R1885 VN.n23 VN.n22 12.1722
R1886 VN.n24 VN.n23 12.1722
R1887 VN.n70 VN.n69 12.1722
R1888 VN.n69 VN.n68 12.1722
R1889 VN.n59 VN.n58 5.70674
R1890 VN.n13 VN.n12 5.70674
R1891 VN.n11 VN.n10 2.92171
R1892 VN.n35 VN.n34 2.92171
R1893 VN.n57 VN.n56 2.92171
R1894 VN.n81 VN.n80 2.92171
R1895 VN.n91 VN.n90 0.355081
R1896 VN.n45 VN.n44 0.355081
R1897 VN VN.n45 0.26685
R1898 VN.n90 VN.n47 0.189894
R1899 VN.n86 VN.n47 0.189894
R1900 VN.n86 VN.n85 0.189894
R1901 VN.n85 VN.n84 0.189894
R1902 VN.n84 VN.n49 0.189894
R1903 VN.n79 VN.n49 0.189894
R1904 VN.n79 VN.n78 0.189894
R1905 VN.n78 VN.n77 0.189894
R1906 VN.n77 VN.n51 0.189894
R1907 VN.n73 VN.n51 0.189894
R1908 VN.n73 VN.n72 0.189894
R1909 VN.n72 VN.n71 0.189894
R1910 VN.n71 VN.n53 0.189894
R1911 VN.n66 VN.n53 0.189894
R1912 VN.n66 VN.n65 0.189894
R1913 VN.n65 VN.n64 0.189894
R1914 VN.n64 VN.n55 0.189894
R1915 VN.n60 VN.n55 0.189894
R1916 VN.n60 VN.n59 0.189894
R1917 VN.n14 VN.n13 0.189894
R1918 VN.n14 VN.n9 0.189894
R1919 VN.n18 VN.n9 0.189894
R1920 VN.n19 VN.n18 0.189894
R1921 VN.n20 VN.n19 0.189894
R1922 VN.n20 VN.n7 0.189894
R1923 VN.n25 VN.n7 0.189894
R1924 VN.n26 VN.n25 0.189894
R1925 VN.n27 VN.n26 0.189894
R1926 VN.n27 VN.n5 0.189894
R1927 VN.n31 VN.n5 0.189894
R1928 VN.n32 VN.n31 0.189894
R1929 VN.n33 VN.n32 0.189894
R1930 VN.n33 VN.n3 0.189894
R1931 VN.n38 VN.n3 0.189894
R1932 VN.n39 VN.n38 0.189894
R1933 VN.n40 VN.n39 0.189894
R1934 VN.n40 VN.n1 0.189894
R1935 VN.n44 VN.n1 0.189894
R1936 VDD2.n1 VDD2.t3 75.8781
R1937 VDD2.n3 VDD2.n2 73.2261
R1938 VDD2 VDD2.n7 73.2233
R1939 VDD2.n4 VDD2.t0 73.0248
R1940 VDD2.n6 VDD2.n5 71.1416
R1941 VDD2.n1 VDD2.n0 71.1413
R1942 VDD2.n4 VDD2.n3 52.1485
R1943 VDD2.n6 VDD2.n4 2.85395
R1944 VDD2.n7 VDD2.t4 1.88376
R1945 VDD2.n7 VDD2.t7 1.88376
R1946 VDD2.n5 VDD2.t1 1.88376
R1947 VDD2.n5 VDD2.t2 1.88376
R1948 VDD2.n2 VDD2.t8 1.88376
R1949 VDD2.n2 VDD2.t5 1.88376
R1950 VDD2.n0 VDD2.t9 1.88376
R1951 VDD2.n0 VDD2.t6 1.88376
R1952 VDD2 VDD2.n6 0.772052
R1953 VDD2.n3 VDD2.n1 0.658516
C0 VTAIL w_n4942_n4420# 3.98944f
C1 VN VDD2 15.5104f
C2 VN VDD1 0.153929f
C3 VP w_n4942_n4420# 11.4498f
C4 VTAIL VP 16.092499f
C5 VDD2 B 3.18075f
C6 VN w_n4942_n4420# 10.805201f
C7 B VDD1 3.04804f
C8 VTAIL VN 16.0782f
C9 VDD2 VDD1 2.42263f
C10 VN VP 9.94423f
C11 B w_n4942_n4420# 12.660701f
C12 VTAIL B 5.09062f
C13 VDD2 w_n4942_n4420# 3.46028f
C14 VTAIL VDD2 12.838901f
C15 VDD1 w_n4942_n4420# 3.29698f
C16 VTAIL VDD1 12.786099f
C17 VP B 2.52365f
C18 VP VDD2 0.632134f
C19 VP VDD1 15.9839f
C20 VN B 1.43762f
C21 VDD2 VSUBS 2.40806f
C22 VDD1 VSUBS 2.252234f
C23 VTAIL VSUBS 1.579608f
C24 VN VSUBS 8.49818f
C25 VP VSUBS 4.921781f
C26 B VSUBS 6.282527f
C27 w_n4942_n4420# VSUBS 0.267283p
C28 VDD2.t3 VSUBS 4.25075f
C29 VDD2.t9 VSUBS 0.391935f
C30 VDD2.t6 VSUBS 0.391935f
C31 VDD2.n0 VSUBS 3.24804f
C32 VDD2.n1 VSUBS 1.77694f
C33 VDD2.t8 VSUBS 0.391935f
C34 VDD2.t5 VSUBS 0.391935f
C35 VDD2.n2 VSUBS 3.27718f
C36 VDD2.n3 VSUBS 4.25779f
C37 VDD2.t0 VSUBS 4.21574f
C38 VDD2.n4 VSUBS 4.56479f
C39 VDD2.t1 VSUBS 0.391935f
C40 VDD2.t2 VSUBS 0.391935f
C41 VDD2.n5 VSUBS 3.24804f
C42 VDD2.n6 VSUBS 0.890044f
C43 VDD2.t4 VSUBS 0.391935f
C44 VDD2.t7 VSUBS 0.391935f
C45 VDD2.n7 VSUBS 3.27712f
C46 VN.t4 VSUBS 3.34391f
C47 VN.n0 VSUBS 1.24895f
C48 VN.n1 VSUBS 0.023655f
C49 VN.n2 VSUBS 0.032359f
C50 VN.n3 VSUBS 0.023655f
C51 VN.t1 VSUBS 3.34391f
C52 VN.n4 VSUBS 0.044308f
C53 VN.n5 VSUBS 0.023655f
C54 VN.n6 VSUBS 0.044308f
C55 VN.n7 VSUBS 0.023655f
C56 VN.t3 VSUBS 3.34391f
C57 VN.n8 VSUBS 0.043862f
C58 VN.n9 VSUBS 0.023655f
C59 VN.n10 VSUBS 0.025057f
C60 VN.t0 VSUBS 3.34391f
C61 VN.n11 VSUBS 1.22601f
C62 VN.t6 VSUBS 3.58612f
C63 VN.n12 VSUBS 1.19709f
C64 VN.n13 VSUBS 0.256027f
C65 VN.n14 VSUBS 0.023655f
C66 VN.n15 VSUBS 0.044308f
C67 VN.n16 VSUBS 0.047754f
C68 VN.n17 VSUBS 0.022057f
C69 VN.n18 VSUBS 0.023655f
C70 VN.n19 VSUBS 0.023655f
C71 VN.n20 VSUBS 0.023655f
C72 VN.n21 VSUBS 0.044308f
C73 VN.n22 VSUBS 0.03337f
C74 VN.n23 VSUBS 1.15846f
C75 VN.n24 VSUBS 0.03337f
C76 VN.n25 VSUBS 0.023655f
C77 VN.n26 VSUBS 0.023655f
C78 VN.n27 VSUBS 0.023655f
C79 VN.n28 VSUBS 0.043862f
C80 VN.n29 VSUBS 0.022057f
C81 VN.n30 VSUBS 0.047754f
C82 VN.n31 VSUBS 0.023655f
C83 VN.n32 VSUBS 0.023655f
C84 VN.n33 VSUBS 0.023655f
C85 VN.n34 VSUBS 0.025057f
C86 VN.n35 VSUBS 1.15846f
C87 VN.n36 VSUBS 0.041683f
C88 VN.n37 VSUBS 0.044308f
C89 VN.n38 VSUBS 0.023655f
C90 VN.n39 VSUBS 0.023655f
C91 VN.n40 VSUBS 0.023655f
C92 VN.n41 VSUBS 0.037006f
C93 VN.n42 VSUBS 0.044308f
C94 VN.n43 VSUBS 0.03862f
C95 VN.n44 VSUBS 0.038185f
C96 VN.n45 VSUBS 0.05105f
C97 VN.t9 VSUBS 3.34391f
C98 VN.n46 VSUBS 1.24895f
C99 VN.n47 VSUBS 0.023655f
C100 VN.n48 VSUBS 0.032359f
C101 VN.n49 VSUBS 0.023655f
C102 VN.t8 VSUBS 3.34391f
C103 VN.n50 VSUBS 0.044308f
C104 VN.n51 VSUBS 0.023655f
C105 VN.n52 VSUBS 0.044308f
C106 VN.n53 VSUBS 0.023655f
C107 VN.t7 VSUBS 3.34391f
C108 VN.n54 VSUBS 0.043862f
C109 VN.n55 VSUBS 0.023655f
C110 VN.n56 VSUBS 0.025057f
C111 VN.t2 VSUBS 3.58612f
C112 VN.t5 VSUBS 3.34391f
C113 VN.n57 VSUBS 1.22601f
C114 VN.n58 VSUBS 1.19709f
C115 VN.n59 VSUBS 0.256027f
C116 VN.n60 VSUBS 0.023655f
C117 VN.n61 VSUBS 0.044308f
C118 VN.n62 VSUBS 0.047754f
C119 VN.n63 VSUBS 0.022057f
C120 VN.n64 VSUBS 0.023655f
C121 VN.n65 VSUBS 0.023655f
C122 VN.n66 VSUBS 0.023655f
C123 VN.n67 VSUBS 0.044308f
C124 VN.n68 VSUBS 0.03337f
C125 VN.n69 VSUBS 1.15846f
C126 VN.n70 VSUBS 0.03337f
C127 VN.n71 VSUBS 0.023655f
C128 VN.n72 VSUBS 0.023655f
C129 VN.n73 VSUBS 0.023655f
C130 VN.n74 VSUBS 0.043862f
C131 VN.n75 VSUBS 0.022057f
C132 VN.n76 VSUBS 0.047754f
C133 VN.n77 VSUBS 0.023655f
C134 VN.n78 VSUBS 0.023655f
C135 VN.n79 VSUBS 0.023655f
C136 VN.n80 VSUBS 0.025057f
C137 VN.n81 VSUBS 1.15846f
C138 VN.n82 VSUBS 0.041683f
C139 VN.n83 VSUBS 0.044308f
C140 VN.n84 VSUBS 0.023655f
C141 VN.n85 VSUBS 0.023655f
C142 VN.n86 VSUBS 0.023655f
C143 VN.n87 VSUBS 0.037006f
C144 VN.n88 VSUBS 0.044308f
C145 VN.n89 VSUBS 0.03862f
C146 VN.n90 VSUBS 0.038185f
C147 VN.n91 VSUBS 1.70492f
C148 VTAIL.t9 VSUBS 0.378392f
C149 VTAIL.t0 VSUBS 0.378392f
C150 VTAIL.n0 VSUBS 2.97351f
C151 VTAIL.n1 VSUBS 1.02588f
C152 VTAIL.t14 VSUBS 3.88424f
C153 VTAIL.n2 VSUBS 1.20569f
C154 VTAIL.t15 VSUBS 0.378392f
C155 VTAIL.t17 VSUBS 0.378392f
C156 VTAIL.n3 VSUBS 2.97351f
C157 VTAIL.n4 VSUBS 1.16999f
C158 VTAIL.t16 VSUBS 0.378392f
C159 VTAIL.t18 VSUBS 0.378392f
C160 VTAIL.n5 VSUBS 2.97351f
C161 VTAIL.n6 VSUBS 3.13203f
C162 VTAIL.t2 VSUBS 0.378392f
C163 VTAIL.t3 VSUBS 0.378392f
C164 VTAIL.n7 VSUBS 2.97351f
C165 VTAIL.n8 VSUBS 3.13202f
C166 VTAIL.t4 VSUBS 0.378392f
C167 VTAIL.t5 VSUBS 0.378392f
C168 VTAIL.n9 VSUBS 2.97351f
C169 VTAIL.n10 VSUBS 1.16999f
C170 VTAIL.t8 VSUBS 3.88427f
C171 VTAIL.n11 VSUBS 1.20566f
C172 VTAIL.t10 VSUBS 0.378392f
C173 VTAIL.t12 VSUBS 0.378392f
C174 VTAIL.n12 VSUBS 2.97351f
C175 VTAIL.n13 VSUBS 1.08445f
C176 VTAIL.t13 VSUBS 0.378392f
C177 VTAIL.t19 VSUBS 0.378392f
C178 VTAIL.n14 VSUBS 2.97351f
C179 VTAIL.n15 VSUBS 1.16999f
C180 VTAIL.t11 VSUBS 3.88425f
C181 VTAIL.n16 VSUBS 2.99819f
C182 VTAIL.t6 VSUBS 3.88424f
C183 VTAIL.n17 VSUBS 2.99819f
C184 VTAIL.t7 VSUBS 0.378392f
C185 VTAIL.t1 VSUBS 0.378392f
C186 VTAIL.n18 VSUBS 2.97351f
C187 VTAIL.n19 VSUBS 0.973481f
C188 VDD1.t2 VSUBS 4.25007f
C189 VDD1.t0 VSUBS 0.391871f
C190 VDD1.t4 VSUBS 0.391871f
C191 VDD1.n0 VSUBS 3.24751f
C192 VDD1.n1 VSUBS 1.78612f
C193 VDD1.t1 VSUBS 4.25005f
C194 VDD1.t7 VSUBS 0.391871f
C195 VDD1.t9 VSUBS 0.391871f
C196 VDD1.n2 VSUBS 3.24751f
C197 VDD1.n3 VSUBS 1.77665f
C198 VDD1.t6 VSUBS 0.391871f
C199 VDD1.t3 VSUBS 0.391871f
C200 VDD1.n4 VSUBS 3.27664f
C201 VDD1.n5 VSUBS 4.41659f
C202 VDD1.t8 VSUBS 0.391871f
C203 VDD1.t5 VSUBS 0.391871f
C204 VDD1.n6 VSUBS 3.2475f
C205 VDD1.n7 VSUBS 4.60222f
C206 VP.t5 VSUBS 3.57636f
C207 VP.n0 VSUBS 1.33577f
C208 VP.n1 VSUBS 0.025299f
C209 VP.n2 VSUBS 0.034609f
C210 VP.n3 VSUBS 0.025299f
C211 VP.t2 VSUBS 3.57636f
C212 VP.n4 VSUBS 0.047388f
C213 VP.n5 VSUBS 0.025299f
C214 VP.n6 VSUBS 0.047388f
C215 VP.n7 VSUBS 0.025299f
C216 VP.t4 VSUBS 3.57636f
C217 VP.n8 VSUBS 0.046911f
C218 VP.n9 VSUBS 0.025299f
C219 VP.n10 VSUBS 0.026799f
C220 VP.n11 VSUBS 0.025299f
C221 VP.n12 VSUBS 0.039578f
C222 VP.n13 VSUBS 0.040839f
C223 VP.t3 VSUBS 3.57636f
C224 VP.t8 VSUBS 3.57636f
C225 VP.n14 VSUBS 1.33577f
C226 VP.n15 VSUBS 0.025299f
C227 VP.n16 VSUBS 0.034609f
C228 VP.n17 VSUBS 0.025299f
C229 VP.t0 VSUBS 3.57636f
C230 VP.n18 VSUBS 0.047388f
C231 VP.n19 VSUBS 0.025299f
C232 VP.n20 VSUBS 0.047388f
C233 VP.n21 VSUBS 0.025299f
C234 VP.t6 VSUBS 3.57636f
C235 VP.n22 VSUBS 0.046911f
C236 VP.n23 VSUBS 0.025299f
C237 VP.n24 VSUBS 0.026799f
C238 VP.t9 VSUBS 3.8354f
C239 VP.t7 VSUBS 3.57636f
C240 VP.n25 VSUBS 1.31124f
C241 VP.n26 VSUBS 1.28031f
C242 VP.n27 VSUBS 0.273824f
C243 VP.n28 VSUBS 0.025299f
C244 VP.n29 VSUBS 0.047388f
C245 VP.n30 VSUBS 0.051073f
C246 VP.n31 VSUBS 0.023591f
C247 VP.n32 VSUBS 0.025299f
C248 VP.n33 VSUBS 0.025299f
C249 VP.n34 VSUBS 0.025299f
C250 VP.n35 VSUBS 0.047388f
C251 VP.n36 VSUBS 0.03569f
C252 VP.n37 VSUBS 1.23899f
C253 VP.n38 VSUBS 0.03569f
C254 VP.n39 VSUBS 0.025299f
C255 VP.n40 VSUBS 0.025299f
C256 VP.n41 VSUBS 0.025299f
C257 VP.n42 VSUBS 0.046911f
C258 VP.n43 VSUBS 0.023591f
C259 VP.n44 VSUBS 0.051073f
C260 VP.n45 VSUBS 0.025299f
C261 VP.n46 VSUBS 0.025299f
C262 VP.n47 VSUBS 0.025299f
C263 VP.n48 VSUBS 0.026799f
C264 VP.n49 VSUBS 1.23899f
C265 VP.n50 VSUBS 0.044581f
C266 VP.n51 VSUBS 0.047388f
C267 VP.n52 VSUBS 0.025299f
C268 VP.n53 VSUBS 0.025299f
C269 VP.n54 VSUBS 0.025299f
C270 VP.n55 VSUBS 0.039578f
C271 VP.n56 VSUBS 0.047388f
C272 VP.n57 VSUBS 0.041305f
C273 VP.n58 VSUBS 0.040839f
C274 VP.n59 VSUBS 1.81363f
C275 VP.n60 VSUBS 1.82893f
C276 VP.n61 VSUBS 1.33577f
C277 VP.n62 VSUBS 0.041305f
C278 VP.n63 VSUBS 0.047388f
C279 VP.n64 VSUBS 0.025299f
C280 VP.n65 VSUBS 0.025299f
C281 VP.n66 VSUBS 0.025299f
C282 VP.n67 VSUBS 0.034609f
C283 VP.n68 VSUBS 0.047388f
C284 VP.t1 VSUBS 3.57636f
C285 VP.n69 VSUBS 1.23899f
C286 VP.n70 VSUBS 0.044581f
C287 VP.n71 VSUBS 0.025299f
C288 VP.n72 VSUBS 0.025299f
C289 VP.n73 VSUBS 0.025299f
C290 VP.n74 VSUBS 0.047388f
C291 VP.n75 VSUBS 0.051073f
C292 VP.n76 VSUBS 0.023591f
C293 VP.n77 VSUBS 0.025299f
C294 VP.n78 VSUBS 0.025299f
C295 VP.n79 VSUBS 0.025299f
C296 VP.n80 VSUBS 0.047388f
C297 VP.n81 VSUBS 0.03569f
C298 VP.n82 VSUBS 1.23899f
C299 VP.n83 VSUBS 0.03569f
C300 VP.n84 VSUBS 0.025299f
C301 VP.n85 VSUBS 0.025299f
C302 VP.n86 VSUBS 0.025299f
C303 VP.n87 VSUBS 0.046911f
C304 VP.n88 VSUBS 0.023591f
C305 VP.n89 VSUBS 0.051073f
C306 VP.n90 VSUBS 0.025299f
C307 VP.n91 VSUBS 0.025299f
C308 VP.n92 VSUBS 0.025299f
C309 VP.n93 VSUBS 0.026799f
C310 VP.n94 VSUBS 1.23899f
C311 VP.n95 VSUBS 0.044581f
C312 VP.n96 VSUBS 0.047388f
C313 VP.n97 VSUBS 0.025299f
C314 VP.n98 VSUBS 0.025299f
C315 VP.n99 VSUBS 0.025299f
C316 VP.n100 VSUBS 0.039578f
C317 VP.n101 VSUBS 0.047388f
C318 VP.n102 VSUBS 0.041305f
C319 VP.n103 VSUBS 0.040839f
C320 VP.n104 VSUBS 0.054599f
C321 B.n0 VSUBS 0.007088f
C322 B.n1 VSUBS 0.007088f
C323 B.n2 VSUBS 0.010483f
C324 B.n3 VSUBS 0.008034f
C325 B.n4 VSUBS 0.008034f
C326 B.n5 VSUBS 0.008034f
C327 B.n6 VSUBS 0.008034f
C328 B.n7 VSUBS 0.008034f
C329 B.n8 VSUBS 0.008034f
C330 B.n9 VSUBS 0.008034f
C331 B.n10 VSUBS 0.008034f
C332 B.n11 VSUBS 0.008034f
C333 B.n12 VSUBS 0.008034f
C334 B.n13 VSUBS 0.008034f
C335 B.n14 VSUBS 0.008034f
C336 B.n15 VSUBS 0.008034f
C337 B.n16 VSUBS 0.008034f
C338 B.n17 VSUBS 0.008034f
C339 B.n18 VSUBS 0.008034f
C340 B.n19 VSUBS 0.008034f
C341 B.n20 VSUBS 0.008034f
C342 B.n21 VSUBS 0.008034f
C343 B.n22 VSUBS 0.008034f
C344 B.n23 VSUBS 0.008034f
C345 B.n24 VSUBS 0.008034f
C346 B.n25 VSUBS 0.008034f
C347 B.n26 VSUBS 0.008034f
C348 B.n27 VSUBS 0.008034f
C349 B.n28 VSUBS 0.008034f
C350 B.n29 VSUBS 0.008034f
C351 B.n30 VSUBS 0.008034f
C352 B.n31 VSUBS 0.008034f
C353 B.n32 VSUBS 0.008034f
C354 B.n33 VSUBS 0.008034f
C355 B.n34 VSUBS 0.008034f
C356 B.n35 VSUBS 0.018902f
C357 B.n36 VSUBS 0.008034f
C358 B.n37 VSUBS 0.008034f
C359 B.n38 VSUBS 0.008034f
C360 B.n39 VSUBS 0.008034f
C361 B.n40 VSUBS 0.008034f
C362 B.n41 VSUBS 0.008034f
C363 B.n42 VSUBS 0.008034f
C364 B.n43 VSUBS 0.008034f
C365 B.n44 VSUBS 0.008034f
C366 B.n45 VSUBS 0.008034f
C367 B.n46 VSUBS 0.008034f
C368 B.n47 VSUBS 0.008034f
C369 B.n48 VSUBS 0.008034f
C370 B.n49 VSUBS 0.008034f
C371 B.n50 VSUBS 0.008034f
C372 B.n51 VSUBS 0.008034f
C373 B.n52 VSUBS 0.008034f
C374 B.n53 VSUBS 0.008034f
C375 B.n54 VSUBS 0.008034f
C376 B.n55 VSUBS 0.008034f
C377 B.n56 VSUBS 0.008034f
C378 B.n57 VSUBS 0.008034f
C379 B.n58 VSUBS 0.008034f
C380 B.n59 VSUBS 0.008034f
C381 B.n60 VSUBS 0.008034f
C382 B.n61 VSUBS 0.008034f
C383 B.n62 VSUBS 0.008034f
C384 B.n63 VSUBS 0.008034f
C385 B.t4 VSUBS 0.666755f
C386 B.t5 VSUBS 0.693478f
C387 B.t3 VSUBS 2.6521f
C388 B.n64 VSUBS 0.396164f
C389 B.n65 VSUBS 0.084512f
C390 B.n66 VSUBS 0.008034f
C391 B.n67 VSUBS 0.008034f
C392 B.n68 VSUBS 0.008034f
C393 B.n69 VSUBS 0.008034f
C394 B.n70 VSUBS 0.004489f
C395 B.n71 VSUBS 0.008034f
C396 B.t1 VSUBS 0.666733f
C397 B.t2 VSUBS 0.69346f
C398 B.t0 VSUBS 2.6521f
C399 B.n72 VSUBS 0.396182f
C400 B.n73 VSUBS 0.084534f
C401 B.n74 VSUBS 0.018613f
C402 B.n75 VSUBS 0.008034f
C403 B.n76 VSUBS 0.008034f
C404 B.n77 VSUBS 0.008034f
C405 B.n78 VSUBS 0.008034f
C406 B.n79 VSUBS 0.008034f
C407 B.n80 VSUBS 0.008034f
C408 B.n81 VSUBS 0.008034f
C409 B.n82 VSUBS 0.008034f
C410 B.n83 VSUBS 0.008034f
C411 B.n84 VSUBS 0.008034f
C412 B.n85 VSUBS 0.008034f
C413 B.n86 VSUBS 0.008034f
C414 B.n87 VSUBS 0.008034f
C415 B.n88 VSUBS 0.008034f
C416 B.n89 VSUBS 0.008034f
C417 B.n90 VSUBS 0.008034f
C418 B.n91 VSUBS 0.008034f
C419 B.n92 VSUBS 0.008034f
C420 B.n93 VSUBS 0.008034f
C421 B.n94 VSUBS 0.008034f
C422 B.n95 VSUBS 0.008034f
C423 B.n96 VSUBS 0.008034f
C424 B.n97 VSUBS 0.008034f
C425 B.n98 VSUBS 0.008034f
C426 B.n99 VSUBS 0.008034f
C427 B.n100 VSUBS 0.008034f
C428 B.n101 VSUBS 0.008034f
C429 B.n102 VSUBS 0.017722f
C430 B.n103 VSUBS 0.008034f
C431 B.n104 VSUBS 0.008034f
C432 B.n105 VSUBS 0.008034f
C433 B.n106 VSUBS 0.008034f
C434 B.n107 VSUBS 0.008034f
C435 B.n108 VSUBS 0.008034f
C436 B.n109 VSUBS 0.008034f
C437 B.n110 VSUBS 0.008034f
C438 B.n111 VSUBS 0.008034f
C439 B.n112 VSUBS 0.008034f
C440 B.n113 VSUBS 0.008034f
C441 B.n114 VSUBS 0.008034f
C442 B.n115 VSUBS 0.008034f
C443 B.n116 VSUBS 0.008034f
C444 B.n117 VSUBS 0.008034f
C445 B.n118 VSUBS 0.008034f
C446 B.n119 VSUBS 0.008034f
C447 B.n120 VSUBS 0.008034f
C448 B.n121 VSUBS 0.008034f
C449 B.n122 VSUBS 0.008034f
C450 B.n123 VSUBS 0.008034f
C451 B.n124 VSUBS 0.008034f
C452 B.n125 VSUBS 0.008034f
C453 B.n126 VSUBS 0.008034f
C454 B.n127 VSUBS 0.008034f
C455 B.n128 VSUBS 0.008034f
C456 B.n129 VSUBS 0.008034f
C457 B.n130 VSUBS 0.008034f
C458 B.n131 VSUBS 0.008034f
C459 B.n132 VSUBS 0.008034f
C460 B.n133 VSUBS 0.008034f
C461 B.n134 VSUBS 0.008034f
C462 B.n135 VSUBS 0.008034f
C463 B.n136 VSUBS 0.008034f
C464 B.n137 VSUBS 0.008034f
C465 B.n138 VSUBS 0.008034f
C466 B.n139 VSUBS 0.008034f
C467 B.n140 VSUBS 0.008034f
C468 B.n141 VSUBS 0.008034f
C469 B.n142 VSUBS 0.008034f
C470 B.n143 VSUBS 0.008034f
C471 B.n144 VSUBS 0.008034f
C472 B.n145 VSUBS 0.008034f
C473 B.n146 VSUBS 0.008034f
C474 B.n147 VSUBS 0.008034f
C475 B.n148 VSUBS 0.008034f
C476 B.n149 VSUBS 0.008034f
C477 B.n150 VSUBS 0.008034f
C478 B.n151 VSUBS 0.008034f
C479 B.n152 VSUBS 0.008034f
C480 B.n153 VSUBS 0.008034f
C481 B.n154 VSUBS 0.008034f
C482 B.n155 VSUBS 0.008034f
C483 B.n156 VSUBS 0.008034f
C484 B.n157 VSUBS 0.008034f
C485 B.n158 VSUBS 0.008034f
C486 B.n159 VSUBS 0.008034f
C487 B.n160 VSUBS 0.008034f
C488 B.n161 VSUBS 0.008034f
C489 B.n162 VSUBS 0.008034f
C490 B.n163 VSUBS 0.008034f
C491 B.n164 VSUBS 0.008034f
C492 B.n165 VSUBS 0.008034f
C493 B.n166 VSUBS 0.008034f
C494 B.n167 VSUBS 0.008034f
C495 B.n168 VSUBS 0.008034f
C496 B.n169 VSUBS 0.017914f
C497 B.n170 VSUBS 0.008034f
C498 B.n171 VSUBS 0.008034f
C499 B.n172 VSUBS 0.008034f
C500 B.n173 VSUBS 0.008034f
C501 B.n174 VSUBS 0.008034f
C502 B.n175 VSUBS 0.008034f
C503 B.n176 VSUBS 0.008034f
C504 B.n177 VSUBS 0.008034f
C505 B.n178 VSUBS 0.008034f
C506 B.n179 VSUBS 0.008034f
C507 B.n180 VSUBS 0.008034f
C508 B.n181 VSUBS 0.008034f
C509 B.n182 VSUBS 0.008034f
C510 B.n183 VSUBS 0.008034f
C511 B.n184 VSUBS 0.008034f
C512 B.n185 VSUBS 0.008034f
C513 B.n186 VSUBS 0.008034f
C514 B.n187 VSUBS 0.008034f
C515 B.n188 VSUBS 0.008034f
C516 B.n189 VSUBS 0.008034f
C517 B.n190 VSUBS 0.008034f
C518 B.n191 VSUBS 0.008034f
C519 B.n192 VSUBS 0.008034f
C520 B.n193 VSUBS 0.008034f
C521 B.n194 VSUBS 0.008034f
C522 B.n195 VSUBS 0.008034f
C523 B.n196 VSUBS 0.008034f
C524 B.n197 VSUBS 0.007561f
C525 B.n198 VSUBS 0.008034f
C526 B.n199 VSUBS 0.008034f
C527 B.n200 VSUBS 0.008034f
C528 B.n201 VSUBS 0.008034f
C529 B.n202 VSUBS 0.008034f
C530 B.t8 VSUBS 0.666755f
C531 B.t7 VSUBS 0.693478f
C532 B.t6 VSUBS 2.6521f
C533 B.n203 VSUBS 0.396164f
C534 B.n204 VSUBS 0.084512f
C535 B.n205 VSUBS 0.008034f
C536 B.n206 VSUBS 0.008034f
C537 B.n207 VSUBS 0.008034f
C538 B.n208 VSUBS 0.008034f
C539 B.n209 VSUBS 0.008034f
C540 B.n210 VSUBS 0.008034f
C541 B.n211 VSUBS 0.008034f
C542 B.n212 VSUBS 0.008034f
C543 B.n213 VSUBS 0.008034f
C544 B.n214 VSUBS 0.008034f
C545 B.n215 VSUBS 0.008034f
C546 B.n216 VSUBS 0.008034f
C547 B.n217 VSUBS 0.008034f
C548 B.n218 VSUBS 0.008034f
C549 B.n219 VSUBS 0.008034f
C550 B.n220 VSUBS 0.008034f
C551 B.n221 VSUBS 0.008034f
C552 B.n222 VSUBS 0.008034f
C553 B.n223 VSUBS 0.008034f
C554 B.n224 VSUBS 0.008034f
C555 B.n225 VSUBS 0.008034f
C556 B.n226 VSUBS 0.008034f
C557 B.n227 VSUBS 0.008034f
C558 B.n228 VSUBS 0.008034f
C559 B.n229 VSUBS 0.008034f
C560 B.n230 VSUBS 0.008034f
C561 B.n231 VSUBS 0.008034f
C562 B.n232 VSUBS 0.008034f
C563 B.n233 VSUBS 0.017722f
C564 B.n234 VSUBS 0.008034f
C565 B.n235 VSUBS 0.008034f
C566 B.n236 VSUBS 0.008034f
C567 B.n237 VSUBS 0.008034f
C568 B.n238 VSUBS 0.008034f
C569 B.n239 VSUBS 0.008034f
C570 B.n240 VSUBS 0.008034f
C571 B.n241 VSUBS 0.008034f
C572 B.n242 VSUBS 0.008034f
C573 B.n243 VSUBS 0.008034f
C574 B.n244 VSUBS 0.008034f
C575 B.n245 VSUBS 0.008034f
C576 B.n246 VSUBS 0.008034f
C577 B.n247 VSUBS 0.008034f
C578 B.n248 VSUBS 0.008034f
C579 B.n249 VSUBS 0.008034f
C580 B.n250 VSUBS 0.008034f
C581 B.n251 VSUBS 0.008034f
C582 B.n252 VSUBS 0.008034f
C583 B.n253 VSUBS 0.008034f
C584 B.n254 VSUBS 0.008034f
C585 B.n255 VSUBS 0.008034f
C586 B.n256 VSUBS 0.008034f
C587 B.n257 VSUBS 0.008034f
C588 B.n258 VSUBS 0.008034f
C589 B.n259 VSUBS 0.008034f
C590 B.n260 VSUBS 0.008034f
C591 B.n261 VSUBS 0.008034f
C592 B.n262 VSUBS 0.008034f
C593 B.n263 VSUBS 0.008034f
C594 B.n264 VSUBS 0.008034f
C595 B.n265 VSUBS 0.008034f
C596 B.n266 VSUBS 0.008034f
C597 B.n267 VSUBS 0.008034f
C598 B.n268 VSUBS 0.008034f
C599 B.n269 VSUBS 0.008034f
C600 B.n270 VSUBS 0.008034f
C601 B.n271 VSUBS 0.008034f
C602 B.n272 VSUBS 0.008034f
C603 B.n273 VSUBS 0.008034f
C604 B.n274 VSUBS 0.008034f
C605 B.n275 VSUBS 0.008034f
C606 B.n276 VSUBS 0.008034f
C607 B.n277 VSUBS 0.008034f
C608 B.n278 VSUBS 0.008034f
C609 B.n279 VSUBS 0.008034f
C610 B.n280 VSUBS 0.008034f
C611 B.n281 VSUBS 0.008034f
C612 B.n282 VSUBS 0.008034f
C613 B.n283 VSUBS 0.008034f
C614 B.n284 VSUBS 0.008034f
C615 B.n285 VSUBS 0.008034f
C616 B.n286 VSUBS 0.008034f
C617 B.n287 VSUBS 0.008034f
C618 B.n288 VSUBS 0.008034f
C619 B.n289 VSUBS 0.008034f
C620 B.n290 VSUBS 0.008034f
C621 B.n291 VSUBS 0.008034f
C622 B.n292 VSUBS 0.008034f
C623 B.n293 VSUBS 0.008034f
C624 B.n294 VSUBS 0.008034f
C625 B.n295 VSUBS 0.008034f
C626 B.n296 VSUBS 0.008034f
C627 B.n297 VSUBS 0.008034f
C628 B.n298 VSUBS 0.008034f
C629 B.n299 VSUBS 0.008034f
C630 B.n300 VSUBS 0.008034f
C631 B.n301 VSUBS 0.008034f
C632 B.n302 VSUBS 0.008034f
C633 B.n303 VSUBS 0.008034f
C634 B.n304 VSUBS 0.008034f
C635 B.n305 VSUBS 0.008034f
C636 B.n306 VSUBS 0.008034f
C637 B.n307 VSUBS 0.008034f
C638 B.n308 VSUBS 0.008034f
C639 B.n309 VSUBS 0.008034f
C640 B.n310 VSUBS 0.008034f
C641 B.n311 VSUBS 0.008034f
C642 B.n312 VSUBS 0.008034f
C643 B.n313 VSUBS 0.008034f
C644 B.n314 VSUBS 0.008034f
C645 B.n315 VSUBS 0.008034f
C646 B.n316 VSUBS 0.008034f
C647 B.n317 VSUBS 0.008034f
C648 B.n318 VSUBS 0.008034f
C649 B.n319 VSUBS 0.008034f
C650 B.n320 VSUBS 0.008034f
C651 B.n321 VSUBS 0.008034f
C652 B.n322 VSUBS 0.008034f
C653 B.n323 VSUBS 0.008034f
C654 B.n324 VSUBS 0.008034f
C655 B.n325 VSUBS 0.008034f
C656 B.n326 VSUBS 0.008034f
C657 B.n327 VSUBS 0.008034f
C658 B.n328 VSUBS 0.008034f
C659 B.n329 VSUBS 0.008034f
C660 B.n330 VSUBS 0.008034f
C661 B.n331 VSUBS 0.008034f
C662 B.n332 VSUBS 0.008034f
C663 B.n333 VSUBS 0.008034f
C664 B.n334 VSUBS 0.008034f
C665 B.n335 VSUBS 0.008034f
C666 B.n336 VSUBS 0.008034f
C667 B.n337 VSUBS 0.008034f
C668 B.n338 VSUBS 0.008034f
C669 B.n339 VSUBS 0.008034f
C670 B.n340 VSUBS 0.008034f
C671 B.n341 VSUBS 0.008034f
C672 B.n342 VSUBS 0.008034f
C673 B.n343 VSUBS 0.008034f
C674 B.n344 VSUBS 0.008034f
C675 B.n345 VSUBS 0.008034f
C676 B.n346 VSUBS 0.008034f
C677 B.n347 VSUBS 0.008034f
C678 B.n348 VSUBS 0.008034f
C679 B.n349 VSUBS 0.008034f
C680 B.n350 VSUBS 0.008034f
C681 B.n351 VSUBS 0.008034f
C682 B.n352 VSUBS 0.008034f
C683 B.n353 VSUBS 0.008034f
C684 B.n354 VSUBS 0.008034f
C685 B.n355 VSUBS 0.008034f
C686 B.n356 VSUBS 0.008034f
C687 B.n357 VSUBS 0.008034f
C688 B.n358 VSUBS 0.008034f
C689 B.n359 VSUBS 0.008034f
C690 B.n360 VSUBS 0.008034f
C691 B.n361 VSUBS 0.008034f
C692 B.n362 VSUBS 0.017722f
C693 B.n363 VSUBS 0.018902f
C694 B.n364 VSUBS 0.018902f
C695 B.n365 VSUBS 0.008034f
C696 B.n366 VSUBS 0.008034f
C697 B.n367 VSUBS 0.008034f
C698 B.n368 VSUBS 0.008034f
C699 B.n369 VSUBS 0.008034f
C700 B.n370 VSUBS 0.008034f
C701 B.n371 VSUBS 0.008034f
C702 B.n372 VSUBS 0.008034f
C703 B.n373 VSUBS 0.008034f
C704 B.n374 VSUBS 0.008034f
C705 B.n375 VSUBS 0.008034f
C706 B.n376 VSUBS 0.008034f
C707 B.n377 VSUBS 0.008034f
C708 B.n378 VSUBS 0.008034f
C709 B.n379 VSUBS 0.008034f
C710 B.n380 VSUBS 0.008034f
C711 B.n381 VSUBS 0.008034f
C712 B.n382 VSUBS 0.008034f
C713 B.n383 VSUBS 0.008034f
C714 B.n384 VSUBS 0.008034f
C715 B.n385 VSUBS 0.008034f
C716 B.n386 VSUBS 0.008034f
C717 B.n387 VSUBS 0.008034f
C718 B.n388 VSUBS 0.008034f
C719 B.n389 VSUBS 0.008034f
C720 B.n390 VSUBS 0.008034f
C721 B.n391 VSUBS 0.008034f
C722 B.n392 VSUBS 0.008034f
C723 B.n393 VSUBS 0.008034f
C724 B.n394 VSUBS 0.008034f
C725 B.n395 VSUBS 0.008034f
C726 B.n396 VSUBS 0.008034f
C727 B.n397 VSUBS 0.008034f
C728 B.n398 VSUBS 0.008034f
C729 B.n399 VSUBS 0.008034f
C730 B.n400 VSUBS 0.008034f
C731 B.n401 VSUBS 0.008034f
C732 B.n402 VSUBS 0.008034f
C733 B.n403 VSUBS 0.008034f
C734 B.n404 VSUBS 0.008034f
C735 B.n405 VSUBS 0.008034f
C736 B.n406 VSUBS 0.008034f
C737 B.n407 VSUBS 0.008034f
C738 B.n408 VSUBS 0.008034f
C739 B.n409 VSUBS 0.008034f
C740 B.n410 VSUBS 0.008034f
C741 B.n411 VSUBS 0.008034f
C742 B.n412 VSUBS 0.008034f
C743 B.n413 VSUBS 0.008034f
C744 B.n414 VSUBS 0.008034f
C745 B.n415 VSUBS 0.008034f
C746 B.n416 VSUBS 0.008034f
C747 B.n417 VSUBS 0.008034f
C748 B.n418 VSUBS 0.008034f
C749 B.n419 VSUBS 0.008034f
C750 B.n420 VSUBS 0.008034f
C751 B.n421 VSUBS 0.008034f
C752 B.n422 VSUBS 0.008034f
C753 B.n423 VSUBS 0.008034f
C754 B.n424 VSUBS 0.008034f
C755 B.n425 VSUBS 0.008034f
C756 B.n426 VSUBS 0.008034f
C757 B.n427 VSUBS 0.008034f
C758 B.n428 VSUBS 0.008034f
C759 B.n429 VSUBS 0.008034f
C760 B.n430 VSUBS 0.008034f
C761 B.n431 VSUBS 0.008034f
C762 B.n432 VSUBS 0.008034f
C763 B.n433 VSUBS 0.008034f
C764 B.n434 VSUBS 0.008034f
C765 B.n435 VSUBS 0.008034f
C766 B.n436 VSUBS 0.008034f
C767 B.n437 VSUBS 0.008034f
C768 B.n438 VSUBS 0.008034f
C769 B.n439 VSUBS 0.008034f
C770 B.n440 VSUBS 0.008034f
C771 B.n441 VSUBS 0.008034f
C772 B.n442 VSUBS 0.008034f
C773 B.n443 VSUBS 0.008034f
C774 B.n444 VSUBS 0.008034f
C775 B.n445 VSUBS 0.008034f
C776 B.n446 VSUBS 0.008034f
C777 B.n447 VSUBS 0.008034f
C778 B.n448 VSUBS 0.007561f
C779 B.n449 VSUBS 0.018613f
C780 B.n450 VSUBS 0.004489f
C781 B.n451 VSUBS 0.008034f
C782 B.n452 VSUBS 0.008034f
C783 B.n453 VSUBS 0.008034f
C784 B.n454 VSUBS 0.008034f
C785 B.n455 VSUBS 0.008034f
C786 B.n456 VSUBS 0.008034f
C787 B.n457 VSUBS 0.008034f
C788 B.n458 VSUBS 0.008034f
C789 B.n459 VSUBS 0.008034f
C790 B.n460 VSUBS 0.008034f
C791 B.n461 VSUBS 0.008034f
C792 B.n462 VSUBS 0.008034f
C793 B.t11 VSUBS 0.666733f
C794 B.t10 VSUBS 0.69346f
C795 B.t9 VSUBS 2.6521f
C796 B.n463 VSUBS 0.396182f
C797 B.n464 VSUBS 0.084534f
C798 B.n465 VSUBS 0.018613f
C799 B.n466 VSUBS 0.004489f
C800 B.n467 VSUBS 0.008034f
C801 B.n468 VSUBS 0.008034f
C802 B.n469 VSUBS 0.008034f
C803 B.n470 VSUBS 0.008034f
C804 B.n471 VSUBS 0.008034f
C805 B.n472 VSUBS 0.008034f
C806 B.n473 VSUBS 0.008034f
C807 B.n474 VSUBS 0.008034f
C808 B.n475 VSUBS 0.008034f
C809 B.n476 VSUBS 0.008034f
C810 B.n477 VSUBS 0.008034f
C811 B.n478 VSUBS 0.008034f
C812 B.n479 VSUBS 0.008034f
C813 B.n480 VSUBS 0.008034f
C814 B.n481 VSUBS 0.008034f
C815 B.n482 VSUBS 0.008034f
C816 B.n483 VSUBS 0.008034f
C817 B.n484 VSUBS 0.008034f
C818 B.n485 VSUBS 0.008034f
C819 B.n486 VSUBS 0.008034f
C820 B.n487 VSUBS 0.008034f
C821 B.n488 VSUBS 0.008034f
C822 B.n489 VSUBS 0.008034f
C823 B.n490 VSUBS 0.008034f
C824 B.n491 VSUBS 0.008034f
C825 B.n492 VSUBS 0.008034f
C826 B.n493 VSUBS 0.008034f
C827 B.n494 VSUBS 0.008034f
C828 B.n495 VSUBS 0.008034f
C829 B.n496 VSUBS 0.008034f
C830 B.n497 VSUBS 0.008034f
C831 B.n498 VSUBS 0.008034f
C832 B.n499 VSUBS 0.008034f
C833 B.n500 VSUBS 0.008034f
C834 B.n501 VSUBS 0.008034f
C835 B.n502 VSUBS 0.008034f
C836 B.n503 VSUBS 0.008034f
C837 B.n504 VSUBS 0.008034f
C838 B.n505 VSUBS 0.008034f
C839 B.n506 VSUBS 0.008034f
C840 B.n507 VSUBS 0.008034f
C841 B.n508 VSUBS 0.008034f
C842 B.n509 VSUBS 0.008034f
C843 B.n510 VSUBS 0.008034f
C844 B.n511 VSUBS 0.008034f
C845 B.n512 VSUBS 0.008034f
C846 B.n513 VSUBS 0.008034f
C847 B.n514 VSUBS 0.008034f
C848 B.n515 VSUBS 0.008034f
C849 B.n516 VSUBS 0.008034f
C850 B.n517 VSUBS 0.008034f
C851 B.n518 VSUBS 0.008034f
C852 B.n519 VSUBS 0.008034f
C853 B.n520 VSUBS 0.008034f
C854 B.n521 VSUBS 0.008034f
C855 B.n522 VSUBS 0.008034f
C856 B.n523 VSUBS 0.008034f
C857 B.n524 VSUBS 0.008034f
C858 B.n525 VSUBS 0.008034f
C859 B.n526 VSUBS 0.008034f
C860 B.n527 VSUBS 0.008034f
C861 B.n528 VSUBS 0.008034f
C862 B.n529 VSUBS 0.008034f
C863 B.n530 VSUBS 0.008034f
C864 B.n531 VSUBS 0.008034f
C865 B.n532 VSUBS 0.008034f
C866 B.n533 VSUBS 0.008034f
C867 B.n534 VSUBS 0.008034f
C868 B.n535 VSUBS 0.008034f
C869 B.n536 VSUBS 0.008034f
C870 B.n537 VSUBS 0.008034f
C871 B.n538 VSUBS 0.008034f
C872 B.n539 VSUBS 0.008034f
C873 B.n540 VSUBS 0.008034f
C874 B.n541 VSUBS 0.008034f
C875 B.n542 VSUBS 0.008034f
C876 B.n543 VSUBS 0.008034f
C877 B.n544 VSUBS 0.008034f
C878 B.n545 VSUBS 0.008034f
C879 B.n546 VSUBS 0.008034f
C880 B.n547 VSUBS 0.008034f
C881 B.n548 VSUBS 0.008034f
C882 B.n549 VSUBS 0.008034f
C883 B.n550 VSUBS 0.008034f
C884 B.n551 VSUBS 0.008034f
C885 B.n552 VSUBS 0.018902f
C886 B.n553 VSUBS 0.017722f
C887 B.n554 VSUBS 0.01871f
C888 B.n555 VSUBS 0.008034f
C889 B.n556 VSUBS 0.008034f
C890 B.n557 VSUBS 0.008034f
C891 B.n558 VSUBS 0.008034f
C892 B.n559 VSUBS 0.008034f
C893 B.n560 VSUBS 0.008034f
C894 B.n561 VSUBS 0.008034f
C895 B.n562 VSUBS 0.008034f
C896 B.n563 VSUBS 0.008034f
C897 B.n564 VSUBS 0.008034f
C898 B.n565 VSUBS 0.008034f
C899 B.n566 VSUBS 0.008034f
C900 B.n567 VSUBS 0.008034f
C901 B.n568 VSUBS 0.008034f
C902 B.n569 VSUBS 0.008034f
C903 B.n570 VSUBS 0.008034f
C904 B.n571 VSUBS 0.008034f
C905 B.n572 VSUBS 0.008034f
C906 B.n573 VSUBS 0.008034f
C907 B.n574 VSUBS 0.008034f
C908 B.n575 VSUBS 0.008034f
C909 B.n576 VSUBS 0.008034f
C910 B.n577 VSUBS 0.008034f
C911 B.n578 VSUBS 0.008034f
C912 B.n579 VSUBS 0.008034f
C913 B.n580 VSUBS 0.008034f
C914 B.n581 VSUBS 0.008034f
C915 B.n582 VSUBS 0.008034f
C916 B.n583 VSUBS 0.008034f
C917 B.n584 VSUBS 0.008034f
C918 B.n585 VSUBS 0.008034f
C919 B.n586 VSUBS 0.008034f
C920 B.n587 VSUBS 0.008034f
C921 B.n588 VSUBS 0.008034f
C922 B.n589 VSUBS 0.008034f
C923 B.n590 VSUBS 0.008034f
C924 B.n591 VSUBS 0.008034f
C925 B.n592 VSUBS 0.008034f
C926 B.n593 VSUBS 0.008034f
C927 B.n594 VSUBS 0.008034f
C928 B.n595 VSUBS 0.008034f
C929 B.n596 VSUBS 0.008034f
C930 B.n597 VSUBS 0.008034f
C931 B.n598 VSUBS 0.008034f
C932 B.n599 VSUBS 0.008034f
C933 B.n600 VSUBS 0.008034f
C934 B.n601 VSUBS 0.008034f
C935 B.n602 VSUBS 0.008034f
C936 B.n603 VSUBS 0.008034f
C937 B.n604 VSUBS 0.008034f
C938 B.n605 VSUBS 0.008034f
C939 B.n606 VSUBS 0.008034f
C940 B.n607 VSUBS 0.008034f
C941 B.n608 VSUBS 0.008034f
C942 B.n609 VSUBS 0.008034f
C943 B.n610 VSUBS 0.008034f
C944 B.n611 VSUBS 0.008034f
C945 B.n612 VSUBS 0.008034f
C946 B.n613 VSUBS 0.008034f
C947 B.n614 VSUBS 0.008034f
C948 B.n615 VSUBS 0.008034f
C949 B.n616 VSUBS 0.008034f
C950 B.n617 VSUBS 0.008034f
C951 B.n618 VSUBS 0.008034f
C952 B.n619 VSUBS 0.008034f
C953 B.n620 VSUBS 0.008034f
C954 B.n621 VSUBS 0.008034f
C955 B.n622 VSUBS 0.008034f
C956 B.n623 VSUBS 0.008034f
C957 B.n624 VSUBS 0.008034f
C958 B.n625 VSUBS 0.008034f
C959 B.n626 VSUBS 0.008034f
C960 B.n627 VSUBS 0.008034f
C961 B.n628 VSUBS 0.008034f
C962 B.n629 VSUBS 0.008034f
C963 B.n630 VSUBS 0.008034f
C964 B.n631 VSUBS 0.008034f
C965 B.n632 VSUBS 0.008034f
C966 B.n633 VSUBS 0.008034f
C967 B.n634 VSUBS 0.008034f
C968 B.n635 VSUBS 0.008034f
C969 B.n636 VSUBS 0.008034f
C970 B.n637 VSUBS 0.008034f
C971 B.n638 VSUBS 0.008034f
C972 B.n639 VSUBS 0.008034f
C973 B.n640 VSUBS 0.008034f
C974 B.n641 VSUBS 0.008034f
C975 B.n642 VSUBS 0.008034f
C976 B.n643 VSUBS 0.008034f
C977 B.n644 VSUBS 0.008034f
C978 B.n645 VSUBS 0.008034f
C979 B.n646 VSUBS 0.008034f
C980 B.n647 VSUBS 0.008034f
C981 B.n648 VSUBS 0.008034f
C982 B.n649 VSUBS 0.008034f
C983 B.n650 VSUBS 0.008034f
C984 B.n651 VSUBS 0.008034f
C985 B.n652 VSUBS 0.008034f
C986 B.n653 VSUBS 0.008034f
C987 B.n654 VSUBS 0.008034f
C988 B.n655 VSUBS 0.008034f
C989 B.n656 VSUBS 0.008034f
C990 B.n657 VSUBS 0.008034f
C991 B.n658 VSUBS 0.008034f
C992 B.n659 VSUBS 0.008034f
C993 B.n660 VSUBS 0.008034f
C994 B.n661 VSUBS 0.008034f
C995 B.n662 VSUBS 0.008034f
C996 B.n663 VSUBS 0.008034f
C997 B.n664 VSUBS 0.008034f
C998 B.n665 VSUBS 0.008034f
C999 B.n666 VSUBS 0.008034f
C1000 B.n667 VSUBS 0.008034f
C1001 B.n668 VSUBS 0.008034f
C1002 B.n669 VSUBS 0.008034f
C1003 B.n670 VSUBS 0.008034f
C1004 B.n671 VSUBS 0.008034f
C1005 B.n672 VSUBS 0.008034f
C1006 B.n673 VSUBS 0.008034f
C1007 B.n674 VSUBS 0.008034f
C1008 B.n675 VSUBS 0.008034f
C1009 B.n676 VSUBS 0.008034f
C1010 B.n677 VSUBS 0.008034f
C1011 B.n678 VSUBS 0.008034f
C1012 B.n679 VSUBS 0.008034f
C1013 B.n680 VSUBS 0.008034f
C1014 B.n681 VSUBS 0.008034f
C1015 B.n682 VSUBS 0.008034f
C1016 B.n683 VSUBS 0.008034f
C1017 B.n684 VSUBS 0.008034f
C1018 B.n685 VSUBS 0.008034f
C1019 B.n686 VSUBS 0.008034f
C1020 B.n687 VSUBS 0.008034f
C1021 B.n688 VSUBS 0.008034f
C1022 B.n689 VSUBS 0.008034f
C1023 B.n690 VSUBS 0.008034f
C1024 B.n691 VSUBS 0.008034f
C1025 B.n692 VSUBS 0.008034f
C1026 B.n693 VSUBS 0.008034f
C1027 B.n694 VSUBS 0.008034f
C1028 B.n695 VSUBS 0.008034f
C1029 B.n696 VSUBS 0.008034f
C1030 B.n697 VSUBS 0.008034f
C1031 B.n698 VSUBS 0.008034f
C1032 B.n699 VSUBS 0.008034f
C1033 B.n700 VSUBS 0.008034f
C1034 B.n701 VSUBS 0.008034f
C1035 B.n702 VSUBS 0.008034f
C1036 B.n703 VSUBS 0.008034f
C1037 B.n704 VSUBS 0.008034f
C1038 B.n705 VSUBS 0.008034f
C1039 B.n706 VSUBS 0.008034f
C1040 B.n707 VSUBS 0.008034f
C1041 B.n708 VSUBS 0.008034f
C1042 B.n709 VSUBS 0.008034f
C1043 B.n710 VSUBS 0.008034f
C1044 B.n711 VSUBS 0.008034f
C1045 B.n712 VSUBS 0.008034f
C1046 B.n713 VSUBS 0.008034f
C1047 B.n714 VSUBS 0.008034f
C1048 B.n715 VSUBS 0.008034f
C1049 B.n716 VSUBS 0.008034f
C1050 B.n717 VSUBS 0.008034f
C1051 B.n718 VSUBS 0.008034f
C1052 B.n719 VSUBS 0.008034f
C1053 B.n720 VSUBS 0.008034f
C1054 B.n721 VSUBS 0.008034f
C1055 B.n722 VSUBS 0.008034f
C1056 B.n723 VSUBS 0.008034f
C1057 B.n724 VSUBS 0.008034f
C1058 B.n725 VSUBS 0.008034f
C1059 B.n726 VSUBS 0.008034f
C1060 B.n727 VSUBS 0.008034f
C1061 B.n728 VSUBS 0.008034f
C1062 B.n729 VSUBS 0.008034f
C1063 B.n730 VSUBS 0.008034f
C1064 B.n731 VSUBS 0.008034f
C1065 B.n732 VSUBS 0.008034f
C1066 B.n733 VSUBS 0.008034f
C1067 B.n734 VSUBS 0.008034f
C1068 B.n735 VSUBS 0.008034f
C1069 B.n736 VSUBS 0.008034f
C1070 B.n737 VSUBS 0.008034f
C1071 B.n738 VSUBS 0.008034f
C1072 B.n739 VSUBS 0.008034f
C1073 B.n740 VSUBS 0.008034f
C1074 B.n741 VSUBS 0.008034f
C1075 B.n742 VSUBS 0.008034f
C1076 B.n743 VSUBS 0.008034f
C1077 B.n744 VSUBS 0.008034f
C1078 B.n745 VSUBS 0.008034f
C1079 B.n746 VSUBS 0.008034f
C1080 B.n747 VSUBS 0.008034f
C1081 B.n748 VSUBS 0.008034f
C1082 B.n749 VSUBS 0.008034f
C1083 B.n750 VSUBS 0.008034f
C1084 B.n751 VSUBS 0.008034f
C1085 B.n752 VSUBS 0.008034f
C1086 B.n753 VSUBS 0.017722f
C1087 B.n754 VSUBS 0.018902f
C1088 B.n755 VSUBS 0.018902f
C1089 B.n756 VSUBS 0.008034f
C1090 B.n757 VSUBS 0.008034f
C1091 B.n758 VSUBS 0.008034f
C1092 B.n759 VSUBS 0.008034f
C1093 B.n760 VSUBS 0.008034f
C1094 B.n761 VSUBS 0.008034f
C1095 B.n762 VSUBS 0.008034f
C1096 B.n763 VSUBS 0.008034f
C1097 B.n764 VSUBS 0.008034f
C1098 B.n765 VSUBS 0.008034f
C1099 B.n766 VSUBS 0.008034f
C1100 B.n767 VSUBS 0.008034f
C1101 B.n768 VSUBS 0.008034f
C1102 B.n769 VSUBS 0.008034f
C1103 B.n770 VSUBS 0.008034f
C1104 B.n771 VSUBS 0.008034f
C1105 B.n772 VSUBS 0.008034f
C1106 B.n773 VSUBS 0.008034f
C1107 B.n774 VSUBS 0.008034f
C1108 B.n775 VSUBS 0.008034f
C1109 B.n776 VSUBS 0.008034f
C1110 B.n777 VSUBS 0.008034f
C1111 B.n778 VSUBS 0.008034f
C1112 B.n779 VSUBS 0.008034f
C1113 B.n780 VSUBS 0.008034f
C1114 B.n781 VSUBS 0.008034f
C1115 B.n782 VSUBS 0.008034f
C1116 B.n783 VSUBS 0.008034f
C1117 B.n784 VSUBS 0.008034f
C1118 B.n785 VSUBS 0.008034f
C1119 B.n786 VSUBS 0.008034f
C1120 B.n787 VSUBS 0.008034f
C1121 B.n788 VSUBS 0.008034f
C1122 B.n789 VSUBS 0.008034f
C1123 B.n790 VSUBS 0.008034f
C1124 B.n791 VSUBS 0.008034f
C1125 B.n792 VSUBS 0.008034f
C1126 B.n793 VSUBS 0.008034f
C1127 B.n794 VSUBS 0.008034f
C1128 B.n795 VSUBS 0.008034f
C1129 B.n796 VSUBS 0.008034f
C1130 B.n797 VSUBS 0.008034f
C1131 B.n798 VSUBS 0.008034f
C1132 B.n799 VSUBS 0.008034f
C1133 B.n800 VSUBS 0.008034f
C1134 B.n801 VSUBS 0.008034f
C1135 B.n802 VSUBS 0.008034f
C1136 B.n803 VSUBS 0.008034f
C1137 B.n804 VSUBS 0.008034f
C1138 B.n805 VSUBS 0.008034f
C1139 B.n806 VSUBS 0.008034f
C1140 B.n807 VSUBS 0.008034f
C1141 B.n808 VSUBS 0.008034f
C1142 B.n809 VSUBS 0.008034f
C1143 B.n810 VSUBS 0.008034f
C1144 B.n811 VSUBS 0.008034f
C1145 B.n812 VSUBS 0.008034f
C1146 B.n813 VSUBS 0.008034f
C1147 B.n814 VSUBS 0.008034f
C1148 B.n815 VSUBS 0.008034f
C1149 B.n816 VSUBS 0.008034f
C1150 B.n817 VSUBS 0.008034f
C1151 B.n818 VSUBS 0.008034f
C1152 B.n819 VSUBS 0.008034f
C1153 B.n820 VSUBS 0.008034f
C1154 B.n821 VSUBS 0.008034f
C1155 B.n822 VSUBS 0.008034f
C1156 B.n823 VSUBS 0.008034f
C1157 B.n824 VSUBS 0.008034f
C1158 B.n825 VSUBS 0.008034f
C1159 B.n826 VSUBS 0.008034f
C1160 B.n827 VSUBS 0.008034f
C1161 B.n828 VSUBS 0.008034f
C1162 B.n829 VSUBS 0.008034f
C1163 B.n830 VSUBS 0.008034f
C1164 B.n831 VSUBS 0.008034f
C1165 B.n832 VSUBS 0.008034f
C1166 B.n833 VSUBS 0.008034f
C1167 B.n834 VSUBS 0.008034f
C1168 B.n835 VSUBS 0.008034f
C1169 B.n836 VSUBS 0.008034f
C1170 B.n837 VSUBS 0.008034f
C1171 B.n838 VSUBS 0.007561f
C1172 B.n839 VSUBS 0.008034f
C1173 B.n840 VSUBS 0.008034f
C1174 B.n841 VSUBS 0.008034f
C1175 B.n842 VSUBS 0.008034f
C1176 B.n843 VSUBS 0.008034f
C1177 B.n844 VSUBS 0.008034f
C1178 B.n845 VSUBS 0.008034f
C1179 B.n846 VSUBS 0.008034f
C1180 B.n847 VSUBS 0.008034f
C1181 B.n848 VSUBS 0.008034f
C1182 B.n849 VSUBS 0.008034f
C1183 B.n850 VSUBS 0.008034f
C1184 B.n851 VSUBS 0.008034f
C1185 B.n852 VSUBS 0.008034f
C1186 B.n853 VSUBS 0.008034f
C1187 B.n854 VSUBS 0.004489f
C1188 B.n855 VSUBS 0.018613f
C1189 B.n856 VSUBS 0.007561f
C1190 B.n857 VSUBS 0.008034f
C1191 B.n858 VSUBS 0.008034f
C1192 B.n859 VSUBS 0.008034f
C1193 B.n860 VSUBS 0.008034f
C1194 B.n861 VSUBS 0.008034f
C1195 B.n862 VSUBS 0.008034f
C1196 B.n863 VSUBS 0.008034f
C1197 B.n864 VSUBS 0.008034f
C1198 B.n865 VSUBS 0.008034f
C1199 B.n866 VSUBS 0.008034f
C1200 B.n867 VSUBS 0.008034f
C1201 B.n868 VSUBS 0.008034f
C1202 B.n869 VSUBS 0.008034f
C1203 B.n870 VSUBS 0.008034f
C1204 B.n871 VSUBS 0.008034f
C1205 B.n872 VSUBS 0.008034f
C1206 B.n873 VSUBS 0.008034f
C1207 B.n874 VSUBS 0.008034f
C1208 B.n875 VSUBS 0.008034f
C1209 B.n876 VSUBS 0.008034f
C1210 B.n877 VSUBS 0.008034f
C1211 B.n878 VSUBS 0.008034f
C1212 B.n879 VSUBS 0.008034f
C1213 B.n880 VSUBS 0.008034f
C1214 B.n881 VSUBS 0.008034f
C1215 B.n882 VSUBS 0.008034f
C1216 B.n883 VSUBS 0.008034f
C1217 B.n884 VSUBS 0.008034f
C1218 B.n885 VSUBS 0.008034f
C1219 B.n886 VSUBS 0.008034f
C1220 B.n887 VSUBS 0.008034f
C1221 B.n888 VSUBS 0.008034f
C1222 B.n889 VSUBS 0.008034f
C1223 B.n890 VSUBS 0.008034f
C1224 B.n891 VSUBS 0.008034f
C1225 B.n892 VSUBS 0.008034f
C1226 B.n893 VSUBS 0.008034f
C1227 B.n894 VSUBS 0.008034f
C1228 B.n895 VSUBS 0.008034f
C1229 B.n896 VSUBS 0.008034f
C1230 B.n897 VSUBS 0.008034f
C1231 B.n898 VSUBS 0.008034f
C1232 B.n899 VSUBS 0.008034f
C1233 B.n900 VSUBS 0.008034f
C1234 B.n901 VSUBS 0.008034f
C1235 B.n902 VSUBS 0.008034f
C1236 B.n903 VSUBS 0.008034f
C1237 B.n904 VSUBS 0.008034f
C1238 B.n905 VSUBS 0.008034f
C1239 B.n906 VSUBS 0.008034f
C1240 B.n907 VSUBS 0.008034f
C1241 B.n908 VSUBS 0.008034f
C1242 B.n909 VSUBS 0.008034f
C1243 B.n910 VSUBS 0.008034f
C1244 B.n911 VSUBS 0.008034f
C1245 B.n912 VSUBS 0.008034f
C1246 B.n913 VSUBS 0.008034f
C1247 B.n914 VSUBS 0.008034f
C1248 B.n915 VSUBS 0.008034f
C1249 B.n916 VSUBS 0.008034f
C1250 B.n917 VSUBS 0.008034f
C1251 B.n918 VSUBS 0.008034f
C1252 B.n919 VSUBS 0.008034f
C1253 B.n920 VSUBS 0.008034f
C1254 B.n921 VSUBS 0.008034f
C1255 B.n922 VSUBS 0.008034f
C1256 B.n923 VSUBS 0.008034f
C1257 B.n924 VSUBS 0.008034f
C1258 B.n925 VSUBS 0.008034f
C1259 B.n926 VSUBS 0.008034f
C1260 B.n927 VSUBS 0.008034f
C1261 B.n928 VSUBS 0.008034f
C1262 B.n929 VSUBS 0.008034f
C1263 B.n930 VSUBS 0.008034f
C1264 B.n931 VSUBS 0.008034f
C1265 B.n932 VSUBS 0.008034f
C1266 B.n933 VSUBS 0.008034f
C1267 B.n934 VSUBS 0.008034f
C1268 B.n935 VSUBS 0.008034f
C1269 B.n936 VSUBS 0.008034f
C1270 B.n937 VSUBS 0.008034f
C1271 B.n938 VSUBS 0.008034f
C1272 B.n939 VSUBS 0.008034f
C1273 B.n940 VSUBS 0.018902f
C1274 B.n941 VSUBS 0.017722f
C1275 B.n942 VSUBS 0.017722f
C1276 B.n943 VSUBS 0.008034f
C1277 B.n944 VSUBS 0.008034f
C1278 B.n945 VSUBS 0.008034f
C1279 B.n946 VSUBS 0.008034f
C1280 B.n947 VSUBS 0.008034f
C1281 B.n948 VSUBS 0.008034f
C1282 B.n949 VSUBS 0.008034f
C1283 B.n950 VSUBS 0.008034f
C1284 B.n951 VSUBS 0.008034f
C1285 B.n952 VSUBS 0.008034f
C1286 B.n953 VSUBS 0.008034f
C1287 B.n954 VSUBS 0.008034f
C1288 B.n955 VSUBS 0.008034f
C1289 B.n956 VSUBS 0.008034f
C1290 B.n957 VSUBS 0.008034f
C1291 B.n958 VSUBS 0.008034f
C1292 B.n959 VSUBS 0.008034f
C1293 B.n960 VSUBS 0.008034f
C1294 B.n961 VSUBS 0.008034f
C1295 B.n962 VSUBS 0.008034f
C1296 B.n963 VSUBS 0.008034f
C1297 B.n964 VSUBS 0.008034f
C1298 B.n965 VSUBS 0.008034f
C1299 B.n966 VSUBS 0.008034f
C1300 B.n967 VSUBS 0.008034f
C1301 B.n968 VSUBS 0.008034f
C1302 B.n969 VSUBS 0.008034f
C1303 B.n970 VSUBS 0.008034f
C1304 B.n971 VSUBS 0.008034f
C1305 B.n972 VSUBS 0.008034f
C1306 B.n973 VSUBS 0.008034f
C1307 B.n974 VSUBS 0.008034f
C1308 B.n975 VSUBS 0.008034f
C1309 B.n976 VSUBS 0.008034f
C1310 B.n977 VSUBS 0.008034f
C1311 B.n978 VSUBS 0.008034f
C1312 B.n979 VSUBS 0.008034f
C1313 B.n980 VSUBS 0.008034f
C1314 B.n981 VSUBS 0.008034f
C1315 B.n982 VSUBS 0.008034f
C1316 B.n983 VSUBS 0.008034f
C1317 B.n984 VSUBS 0.008034f
C1318 B.n985 VSUBS 0.008034f
C1319 B.n986 VSUBS 0.008034f
C1320 B.n987 VSUBS 0.008034f
C1321 B.n988 VSUBS 0.008034f
C1322 B.n989 VSUBS 0.008034f
C1323 B.n990 VSUBS 0.008034f
C1324 B.n991 VSUBS 0.008034f
C1325 B.n992 VSUBS 0.008034f
C1326 B.n993 VSUBS 0.008034f
C1327 B.n994 VSUBS 0.008034f
C1328 B.n995 VSUBS 0.008034f
C1329 B.n996 VSUBS 0.008034f
C1330 B.n997 VSUBS 0.008034f
C1331 B.n998 VSUBS 0.008034f
C1332 B.n999 VSUBS 0.008034f
C1333 B.n1000 VSUBS 0.008034f
C1334 B.n1001 VSUBS 0.008034f
C1335 B.n1002 VSUBS 0.008034f
C1336 B.n1003 VSUBS 0.008034f
C1337 B.n1004 VSUBS 0.008034f
C1338 B.n1005 VSUBS 0.008034f
C1339 B.n1006 VSUBS 0.008034f
C1340 B.n1007 VSUBS 0.008034f
C1341 B.n1008 VSUBS 0.008034f
C1342 B.n1009 VSUBS 0.008034f
C1343 B.n1010 VSUBS 0.008034f
C1344 B.n1011 VSUBS 0.008034f
C1345 B.n1012 VSUBS 0.008034f
C1346 B.n1013 VSUBS 0.008034f
C1347 B.n1014 VSUBS 0.008034f
C1348 B.n1015 VSUBS 0.008034f
C1349 B.n1016 VSUBS 0.008034f
C1350 B.n1017 VSUBS 0.008034f
C1351 B.n1018 VSUBS 0.008034f
C1352 B.n1019 VSUBS 0.008034f
C1353 B.n1020 VSUBS 0.008034f
C1354 B.n1021 VSUBS 0.008034f
C1355 B.n1022 VSUBS 0.008034f
C1356 B.n1023 VSUBS 0.008034f
C1357 B.n1024 VSUBS 0.008034f
C1358 B.n1025 VSUBS 0.008034f
C1359 B.n1026 VSUBS 0.008034f
C1360 B.n1027 VSUBS 0.008034f
C1361 B.n1028 VSUBS 0.008034f
C1362 B.n1029 VSUBS 0.008034f
C1363 B.n1030 VSUBS 0.008034f
C1364 B.n1031 VSUBS 0.008034f
C1365 B.n1032 VSUBS 0.008034f
C1366 B.n1033 VSUBS 0.008034f
C1367 B.n1034 VSUBS 0.008034f
C1368 B.n1035 VSUBS 0.008034f
C1369 B.n1036 VSUBS 0.008034f
C1370 B.n1037 VSUBS 0.008034f
C1371 B.n1038 VSUBS 0.008034f
C1372 B.n1039 VSUBS 0.010483f
C1373 B.n1040 VSUBS 0.011168f
C1374 B.n1041 VSUBS 0.022208f
.ends

