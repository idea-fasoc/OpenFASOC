* NGSPICE file created from diff_pair_sample_0580.ext - technology: sky130A

.subckt diff_pair_sample_0580 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=3.09
X1 VDD1.t5 VP.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=3.09
X2 VDD1.t4 VP.t1 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=3.09
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=3.09
X4 VDD2.t5 VN.t0 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=3.09
X5 VDD2.t4 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=3.09
X6 VDD2.t3 VN.t2 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=3.09
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=3.09
X8 VTAIL.t0 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=2.53605 ps=15.7 w=15.37 l=3.09
X9 VDD1.t3 VP.t2 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=3.09
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=3.09
X11 VTAIL.t11 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=2.53605 ps=15.7 w=15.37 l=3.09
X12 VDD1.t2 VP.t3 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=3.09
X13 VTAIL.t7 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=2.53605 ps=15.7 w=15.37 l=3.09
X14 VDD2.t0 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=3.09
X15 VTAIL.t5 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=2.53605 ps=15.7 w=15.37 l=3.09
R0 B.n965 B.n964 585
R1 B.n966 B.n965 585
R2 B.n374 B.n147 585
R3 B.n373 B.n372 585
R4 B.n371 B.n370 585
R5 B.n369 B.n368 585
R6 B.n367 B.n366 585
R7 B.n365 B.n364 585
R8 B.n363 B.n362 585
R9 B.n361 B.n360 585
R10 B.n359 B.n358 585
R11 B.n357 B.n356 585
R12 B.n355 B.n354 585
R13 B.n353 B.n352 585
R14 B.n351 B.n350 585
R15 B.n349 B.n348 585
R16 B.n347 B.n346 585
R17 B.n345 B.n344 585
R18 B.n343 B.n342 585
R19 B.n341 B.n340 585
R20 B.n339 B.n338 585
R21 B.n337 B.n336 585
R22 B.n335 B.n334 585
R23 B.n333 B.n332 585
R24 B.n331 B.n330 585
R25 B.n329 B.n328 585
R26 B.n327 B.n326 585
R27 B.n325 B.n324 585
R28 B.n323 B.n322 585
R29 B.n321 B.n320 585
R30 B.n319 B.n318 585
R31 B.n317 B.n316 585
R32 B.n315 B.n314 585
R33 B.n313 B.n312 585
R34 B.n311 B.n310 585
R35 B.n309 B.n308 585
R36 B.n307 B.n306 585
R37 B.n305 B.n304 585
R38 B.n303 B.n302 585
R39 B.n301 B.n300 585
R40 B.n299 B.n298 585
R41 B.n297 B.n296 585
R42 B.n295 B.n294 585
R43 B.n293 B.n292 585
R44 B.n291 B.n290 585
R45 B.n289 B.n288 585
R46 B.n287 B.n286 585
R47 B.n285 B.n284 585
R48 B.n283 B.n282 585
R49 B.n281 B.n280 585
R50 B.n279 B.n278 585
R51 B.n277 B.n276 585
R52 B.n275 B.n274 585
R53 B.n272 B.n271 585
R54 B.n270 B.n269 585
R55 B.n268 B.n267 585
R56 B.n266 B.n265 585
R57 B.n264 B.n263 585
R58 B.n262 B.n261 585
R59 B.n260 B.n259 585
R60 B.n258 B.n257 585
R61 B.n256 B.n255 585
R62 B.n254 B.n253 585
R63 B.n252 B.n251 585
R64 B.n250 B.n249 585
R65 B.n248 B.n247 585
R66 B.n246 B.n245 585
R67 B.n244 B.n243 585
R68 B.n242 B.n241 585
R69 B.n240 B.n239 585
R70 B.n238 B.n237 585
R71 B.n236 B.n235 585
R72 B.n234 B.n233 585
R73 B.n232 B.n231 585
R74 B.n230 B.n229 585
R75 B.n228 B.n227 585
R76 B.n226 B.n225 585
R77 B.n224 B.n223 585
R78 B.n222 B.n221 585
R79 B.n220 B.n219 585
R80 B.n218 B.n217 585
R81 B.n216 B.n215 585
R82 B.n214 B.n213 585
R83 B.n212 B.n211 585
R84 B.n210 B.n209 585
R85 B.n208 B.n207 585
R86 B.n206 B.n205 585
R87 B.n204 B.n203 585
R88 B.n202 B.n201 585
R89 B.n200 B.n199 585
R90 B.n198 B.n197 585
R91 B.n196 B.n195 585
R92 B.n194 B.n193 585
R93 B.n192 B.n191 585
R94 B.n190 B.n189 585
R95 B.n188 B.n187 585
R96 B.n186 B.n185 585
R97 B.n184 B.n183 585
R98 B.n182 B.n181 585
R99 B.n180 B.n179 585
R100 B.n178 B.n177 585
R101 B.n176 B.n175 585
R102 B.n174 B.n173 585
R103 B.n172 B.n171 585
R104 B.n170 B.n169 585
R105 B.n168 B.n167 585
R106 B.n166 B.n165 585
R107 B.n164 B.n163 585
R108 B.n162 B.n161 585
R109 B.n160 B.n159 585
R110 B.n158 B.n157 585
R111 B.n156 B.n155 585
R112 B.n154 B.n153 585
R113 B.n89 B.n88 585
R114 B.n963 B.n90 585
R115 B.n967 B.n90 585
R116 B.n962 B.n961 585
R117 B.n961 B.n86 585
R118 B.n960 B.n85 585
R119 B.n973 B.n85 585
R120 B.n959 B.n84 585
R121 B.n974 B.n84 585
R122 B.n958 B.n83 585
R123 B.n975 B.n83 585
R124 B.n957 B.n956 585
R125 B.n956 B.n79 585
R126 B.n955 B.n78 585
R127 B.n981 B.n78 585
R128 B.n954 B.n77 585
R129 B.n982 B.n77 585
R130 B.n953 B.n76 585
R131 B.n983 B.n76 585
R132 B.n952 B.n951 585
R133 B.n951 B.n72 585
R134 B.n950 B.n71 585
R135 B.n989 B.n71 585
R136 B.n949 B.n70 585
R137 B.n990 B.n70 585
R138 B.n948 B.n69 585
R139 B.n991 B.n69 585
R140 B.n947 B.n946 585
R141 B.n946 B.n65 585
R142 B.n945 B.n64 585
R143 B.n997 B.n64 585
R144 B.n944 B.n63 585
R145 B.n998 B.n63 585
R146 B.n943 B.n62 585
R147 B.n999 B.n62 585
R148 B.n942 B.n941 585
R149 B.n941 B.n58 585
R150 B.n940 B.n57 585
R151 B.n1005 B.n57 585
R152 B.n939 B.n56 585
R153 B.n1006 B.n56 585
R154 B.n938 B.n55 585
R155 B.n1007 B.n55 585
R156 B.n937 B.n936 585
R157 B.n936 B.n54 585
R158 B.n935 B.n50 585
R159 B.n1013 B.n50 585
R160 B.n934 B.n49 585
R161 B.n1014 B.n49 585
R162 B.n933 B.n48 585
R163 B.n1015 B.n48 585
R164 B.n932 B.n931 585
R165 B.n931 B.n44 585
R166 B.n930 B.n43 585
R167 B.n1021 B.n43 585
R168 B.n929 B.n42 585
R169 B.n1022 B.n42 585
R170 B.n928 B.n41 585
R171 B.n1023 B.n41 585
R172 B.n927 B.n926 585
R173 B.n926 B.n37 585
R174 B.n925 B.n36 585
R175 B.n1029 B.n36 585
R176 B.n924 B.n35 585
R177 B.n1030 B.n35 585
R178 B.n923 B.n34 585
R179 B.n1031 B.n34 585
R180 B.n922 B.n921 585
R181 B.n921 B.n30 585
R182 B.n920 B.n29 585
R183 B.n1037 B.n29 585
R184 B.n919 B.n28 585
R185 B.n1038 B.n28 585
R186 B.n918 B.n27 585
R187 B.n1039 B.n27 585
R188 B.n917 B.n916 585
R189 B.n916 B.n23 585
R190 B.n915 B.n22 585
R191 B.n1045 B.n22 585
R192 B.n914 B.n21 585
R193 B.n1046 B.n21 585
R194 B.n913 B.n20 585
R195 B.n1047 B.n20 585
R196 B.n912 B.n911 585
R197 B.n911 B.n19 585
R198 B.n910 B.n15 585
R199 B.n1053 B.n15 585
R200 B.n909 B.n14 585
R201 B.n1054 B.n14 585
R202 B.n908 B.n13 585
R203 B.n1055 B.n13 585
R204 B.n907 B.n906 585
R205 B.n906 B.n12 585
R206 B.n905 B.n904 585
R207 B.n905 B.n8 585
R208 B.n903 B.n7 585
R209 B.n1062 B.n7 585
R210 B.n902 B.n6 585
R211 B.n1063 B.n6 585
R212 B.n901 B.n5 585
R213 B.n1064 B.n5 585
R214 B.n900 B.n899 585
R215 B.n899 B.n4 585
R216 B.n898 B.n375 585
R217 B.n898 B.n897 585
R218 B.n888 B.n376 585
R219 B.n377 B.n376 585
R220 B.n890 B.n889 585
R221 B.n891 B.n890 585
R222 B.n887 B.n382 585
R223 B.n382 B.n381 585
R224 B.n886 B.n885 585
R225 B.n885 B.n884 585
R226 B.n384 B.n383 585
R227 B.n877 B.n384 585
R228 B.n876 B.n875 585
R229 B.n878 B.n876 585
R230 B.n874 B.n389 585
R231 B.n389 B.n388 585
R232 B.n873 B.n872 585
R233 B.n872 B.n871 585
R234 B.n391 B.n390 585
R235 B.n392 B.n391 585
R236 B.n864 B.n863 585
R237 B.n865 B.n864 585
R238 B.n862 B.n397 585
R239 B.n397 B.n396 585
R240 B.n861 B.n860 585
R241 B.n860 B.n859 585
R242 B.n399 B.n398 585
R243 B.n400 B.n399 585
R244 B.n852 B.n851 585
R245 B.n853 B.n852 585
R246 B.n850 B.n404 585
R247 B.n408 B.n404 585
R248 B.n849 B.n848 585
R249 B.n848 B.n847 585
R250 B.n406 B.n405 585
R251 B.n407 B.n406 585
R252 B.n840 B.n839 585
R253 B.n841 B.n840 585
R254 B.n838 B.n413 585
R255 B.n413 B.n412 585
R256 B.n837 B.n836 585
R257 B.n836 B.n835 585
R258 B.n415 B.n414 585
R259 B.n416 B.n415 585
R260 B.n828 B.n827 585
R261 B.n829 B.n828 585
R262 B.n826 B.n421 585
R263 B.n421 B.n420 585
R264 B.n825 B.n824 585
R265 B.n824 B.n823 585
R266 B.n423 B.n422 585
R267 B.n816 B.n423 585
R268 B.n815 B.n814 585
R269 B.n817 B.n815 585
R270 B.n813 B.n428 585
R271 B.n428 B.n427 585
R272 B.n812 B.n811 585
R273 B.n811 B.n810 585
R274 B.n430 B.n429 585
R275 B.n431 B.n430 585
R276 B.n803 B.n802 585
R277 B.n804 B.n803 585
R278 B.n801 B.n436 585
R279 B.n436 B.n435 585
R280 B.n800 B.n799 585
R281 B.n799 B.n798 585
R282 B.n438 B.n437 585
R283 B.n439 B.n438 585
R284 B.n791 B.n790 585
R285 B.n792 B.n791 585
R286 B.n789 B.n444 585
R287 B.n444 B.n443 585
R288 B.n788 B.n787 585
R289 B.n787 B.n786 585
R290 B.n446 B.n445 585
R291 B.n447 B.n446 585
R292 B.n779 B.n778 585
R293 B.n780 B.n779 585
R294 B.n777 B.n452 585
R295 B.n452 B.n451 585
R296 B.n776 B.n775 585
R297 B.n775 B.n774 585
R298 B.n454 B.n453 585
R299 B.n455 B.n454 585
R300 B.n767 B.n766 585
R301 B.n768 B.n767 585
R302 B.n765 B.n460 585
R303 B.n460 B.n459 585
R304 B.n764 B.n763 585
R305 B.n763 B.n762 585
R306 B.n462 B.n461 585
R307 B.n463 B.n462 585
R308 B.n755 B.n754 585
R309 B.n756 B.n755 585
R310 B.n466 B.n465 585
R311 B.n530 B.n528 585
R312 B.n531 B.n527 585
R313 B.n531 B.n467 585
R314 B.n534 B.n533 585
R315 B.n535 B.n526 585
R316 B.n537 B.n536 585
R317 B.n539 B.n525 585
R318 B.n542 B.n541 585
R319 B.n543 B.n524 585
R320 B.n545 B.n544 585
R321 B.n547 B.n523 585
R322 B.n550 B.n549 585
R323 B.n551 B.n522 585
R324 B.n553 B.n552 585
R325 B.n555 B.n521 585
R326 B.n558 B.n557 585
R327 B.n559 B.n520 585
R328 B.n561 B.n560 585
R329 B.n563 B.n519 585
R330 B.n566 B.n565 585
R331 B.n567 B.n518 585
R332 B.n569 B.n568 585
R333 B.n571 B.n517 585
R334 B.n574 B.n573 585
R335 B.n575 B.n516 585
R336 B.n577 B.n576 585
R337 B.n579 B.n515 585
R338 B.n582 B.n581 585
R339 B.n583 B.n514 585
R340 B.n585 B.n584 585
R341 B.n587 B.n513 585
R342 B.n590 B.n589 585
R343 B.n591 B.n512 585
R344 B.n593 B.n592 585
R345 B.n595 B.n511 585
R346 B.n598 B.n597 585
R347 B.n599 B.n510 585
R348 B.n601 B.n600 585
R349 B.n603 B.n509 585
R350 B.n606 B.n605 585
R351 B.n607 B.n508 585
R352 B.n609 B.n608 585
R353 B.n611 B.n507 585
R354 B.n614 B.n613 585
R355 B.n615 B.n506 585
R356 B.n617 B.n616 585
R357 B.n619 B.n505 585
R358 B.n622 B.n621 585
R359 B.n623 B.n504 585
R360 B.n625 B.n624 585
R361 B.n627 B.n503 585
R362 B.n630 B.n629 585
R363 B.n632 B.n500 585
R364 B.n634 B.n633 585
R365 B.n636 B.n499 585
R366 B.n639 B.n638 585
R367 B.n640 B.n498 585
R368 B.n642 B.n641 585
R369 B.n644 B.n497 585
R370 B.n647 B.n646 585
R371 B.n648 B.n494 585
R372 B.n651 B.n650 585
R373 B.n653 B.n493 585
R374 B.n656 B.n655 585
R375 B.n657 B.n492 585
R376 B.n659 B.n658 585
R377 B.n661 B.n491 585
R378 B.n664 B.n663 585
R379 B.n665 B.n490 585
R380 B.n667 B.n666 585
R381 B.n669 B.n489 585
R382 B.n672 B.n671 585
R383 B.n673 B.n488 585
R384 B.n675 B.n674 585
R385 B.n677 B.n487 585
R386 B.n680 B.n679 585
R387 B.n681 B.n486 585
R388 B.n683 B.n682 585
R389 B.n685 B.n485 585
R390 B.n688 B.n687 585
R391 B.n689 B.n484 585
R392 B.n691 B.n690 585
R393 B.n693 B.n483 585
R394 B.n696 B.n695 585
R395 B.n697 B.n482 585
R396 B.n699 B.n698 585
R397 B.n701 B.n481 585
R398 B.n704 B.n703 585
R399 B.n705 B.n480 585
R400 B.n707 B.n706 585
R401 B.n709 B.n479 585
R402 B.n712 B.n711 585
R403 B.n713 B.n478 585
R404 B.n715 B.n714 585
R405 B.n717 B.n477 585
R406 B.n720 B.n719 585
R407 B.n721 B.n476 585
R408 B.n723 B.n722 585
R409 B.n725 B.n475 585
R410 B.n728 B.n727 585
R411 B.n729 B.n474 585
R412 B.n731 B.n730 585
R413 B.n733 B.n473 585
R414 B.n736 B.n735 585
R415 B.n737 B.n472 585
R416 B.n739 B.n738 585
R417 B.n741 B.n471 585
R418 B.n744 B.n743 585
R419 B.n745 B.n470 585
R420 B.n747 B.n746 585
R421 B.n749 B.n469 585
R422 B.n752 B.n751 585
R423 B.n753 B.n468 585
R424 B.n758 B.n757 585
R425 B.n757 B.n756 585
R426 B.n759 B.n464 585
R427 B.n464 B.n463 585
R428 B.n761 B.n760 585
R429 B.n762 B.n761 585
R430 B.n458 B.n457 585
R431 B.n459 B.n458 585
R432 B.n770 B.n769 585
R433 B.n769 B.n768 585
R434 B.n771 B.n456 585
R435 B.n456 B.n455 585
R436 B.n773 B.n772 585
R437 B.n774 B.n773 585
R438 B.n450 B.n449 585
R439 B.n451 B.n450 585
R440 B.n782 B.n781 585
R441 B.n781 B.n780 585
R442 B.n783 B.n448 585
R443 B.n448 B.n447 585
R444 B.n785 B.n784 585
R445 B.n786 B.n785 585
R446 B.n442 B.n441 585
R447 B.n443 B.n442 585
R448 B.n794 B.n793 585
R449 B.n793 B.n792 585
R450 B.n795 B.n440 585
R451 B.n440 B.n439 585
R452 B.n797 B.n796 585
R453 B.n798 B.n797 585
R454 B.n434 B.n433 585
R455 B.n435 B.n434 585
R456 B.n806 B.n805 585
R457 B.n805 B.n804 585
R458 B.n807 B.n432 585
R459 B.n432 B.n431 585
R460 B.n809 B.n808 585
R461 B.n810 B.n809 585
R462 B.n426 B.n425 585
R463 B.n427 B.n426 585
R464 B.n819 B.n818 585
R465 B.n818 B.n817 585
R466 B.n820 B.n424 585
R467 B.n816 B.n424 585
R468 B.n822 B.n821 585
R469 B.n823 B.n822 585
R470 B.n419 B.n418 585
R471 B.n420 B.n419 585
R472 B.n831 B.n830 585
R473 B.n830 B.n829 585
R474 B.n832 B.n417 585
R475 B.n417 B.n416 585
R476 B.n834 B.n833 585
R477 B.n835 B.n834 585
R478 B.n411 B.n410 585
R479 B.n412 B.n411 585
R480 B.n843 B.n842 585
R481 B.n842 B.n841 585
R482 B.n844 B.n409 585
R483 B.n409 B.n407 585
R484 B.n846 B.n845 585
R485 B.n847 B.n846 585
R486 B.n403 B.n402 585
R487 B.n408 B.n403 585
R488 B.n855 B.n854 585
R489 B.n854 B.n853 585
R490 B.n856 B.n401 585
R491 B.n401 B.n400 585
R492 B.n858 B.n857 585
R493 B.n859 B.n858 585
R494 B.n395 B.n394 585
R495 B.n396 B.n395 585
R496 B.n867 B.n866 585
R497 B.n866 B.n865 585
R498 B.n868 B.n393 585
R499 B.n393 B.n392 585
R500 B.n870 B.n869 585
R501 B.n871 B.n870 585
R502 B.n387 B.n386 585
R503 B.n388 B.n387 585
R504 B.n880 B.n879 585
R505 B.n879 B.n878 585
R506 B.n881 B.n385 585
R507 B.n877 B.n385 585
R508 B.n883 B.n882 585
R509 B.n884 B.n883 585
R510 B.n380 B.n379 585
R511 B.n381 B.n380 585
R512 B.n893 B.n892 585
R513 B.n892 B.n891 585
R514 B.n894 B.n378 585
R515 B.n378 B.n377 585
R516 B.n896 B.n895 585
R517 B.n897 B.n896 585
R518 B.n3 B.n0 585
R519 B.n4 B.n3 585
R520 B.n1061 B.n1 585
R521 B.n1062 B.n1061 585
R522 B.n1060 B.n1059 585
R523 B.n1060 B.n8 585
R524 B.n1058 B.n9 585
R525 B.n12 B.n9 585
R526 B.n1057 B.n1056 585
R527 B.n1056 B.n1055 585
R528 B.n11 B.n10 585
R529 B.n1054 B.n11 585
R530 B.n1052 B.n1051 585
R531 B.n1053 B.n1052 585
R532 B.n1050 B.n16 585
R533 B.n19 B.n16 585
R534 B.n1049 B.n1048 585
R535 B.n1048 B.n1047 585
R536 B.n18 B.n17 585
R537 B.n1046 B.n18 585
R538 B.n1044 B.n1043 585
R539 B.n1045 B.n1044 585
R540 B.n1042 B.n24 585
R541 B.n24 B.n23 585
R542 B.n1041 B.n1040 585
R543 B.n1040 B.n1039 585
R544 B.n26 B.n25 585
R545 B.n1038 B.n26 585
R546 B.n1036 B.n1035 585
R547 B.n1037 B.n1036 585
R548 B.n1034 B.n31 585
R549 B.n31 B.n30 585
R550 B.n1033 B.n1032 585
R551 B.n1032 B.n1031 585
R552 B.n33 B.n32 585
R553 B.n1030 B.n33 585
R554 B.n1028 B.n1027 585
R555 B.n1029 B.n1028 585
R556 B.n1026 B.n38 585
R557 B.n38 B.n37 585
R558 B.n1025 B.n1024 585
R559 B.n1024 B.n1023 585
R560 B.n40 B.n39 585
R561 B.n1022 B.n40 585
R562 B.n1020 B.n1019 585
R563 B.n1021 B.n1020 585
R564 B.n1018 B.n45 585
R565 B.n45 B.n44 585
R566 B.n1017 B.n1016 585
R567 B.n1016 B.n1015 585
R568 B.n47 B.n46 585
R569 B.n1014 B.n47 585
R570 B.n1012 B.n1011 585
R571 B.n1013 B.n1012 585
R572 B.n1010 B.n51 585
R573 B.n54 B.n51 585
R574 B.n1009 B.n1008 585
R575 B.n1008 B.n1007 585
R576 B.n53 B.n52 585
R577 B.n1006 B.n53 585
R578 B.n1004 B.n1003 585
R579 B.n1005 B.n1004 585
R580 B.n1002 B.n59 585
R581 B.n59 B.n58 585
R582 B.n1001 B.n1000 585
R583 B.n1000 B.n999 585
R584 B.n61 B.n60 585
R585 B.n998 B.n61 585
R586 B.n996 B.n995 585
R587 B.n997 B.n996 585
R588 B.n994 B.n66 585
R589 B.n66 B.n65 585
R590 B.n993 B.n992 585
R591 B.n992 B.n991 585
R592 B.n68 B.n67 585
R593 B.n990 B.n68 585
R594 B.n988 B.n987 585
R595 B.n989 B.n988 585
R596 B.n986 B.n73 585
R597 B.n73 B.n72 585
R598 B.n985 B.n984 585
R599 B.n984 B.n983 585
R600 B.n75 B.n74 585
R601 B.n982 B.n75 585
R602 B.n980 B.n979 585
R603 B.n981 B.n980 585
R604 B.n978 B.n80 585
R605 B.n80 B.n79 585
R606 B.n977 B.n976 585
R607 B.n976 B.n975 585
R608 B.n82 B.n81 585
R609 B.n974 B.n82 585
R610 B.n972 B.n971 585
R611 B.n973 B.n972 585
R612 B.n970 B.n87 585
R613 B.n87 B.n86 585
R614 B.n969 B.n968 585
R615 B.n968 B.n967 585
R616 B.n1065 B.n1064 585
R617 B.n1063 B.n2 585
R618 B.n968 B.n89 444.452
R619 B.n965 B.n90 444.452
R620 B.n755 B.n468 444.452
R621 B.n757 B.n466 444.452
R622 B.n148 B.t8 406.315
R623 B.n495 B.t13 406.315
R624 B.n150 B.t18 406.315
R625 B.n501 B.t16 406.315
R626 B.n149 B.t9 339.988
R627 B.n496 B.t12 339.988
R628 B.n151 B.t19 339.988
R629 B.n502 B.t15 339.988
R630 B.n150 B.t17 328.56
R631 B.n148 B.t6 328.56
R632 B.n495 B.t10 328.56
R633 B.n501 B.t14 328.56
R634 B.n966 B.n146 256.663
R635 B.n966 B.n145 256.663
R636 B.n966 B.n144 256.663
R637 B.n966 B.n143 256.663
R638 B.n966 B.n142 256.663
R639 B.n966 B.n141 256.663
R640 B.n966 B.n140 256.663
R641 B.n966 B.n139 256.663
R642 B.n966 B.n138 256.663
R643 B.n966 B.n137 256.663
R644 B.n966 B.n136 256.663
R645 B.n966 B.n135 256.663
R646 B.n966 B.n134 256.663
R647 B.n966 B.n133 256.663
R648 B.n966 B.n132 256.663
R649 B.n966 B.n131 256.663
R650 B.n966 B.n130 256.663
R651 B.n966 B.n129 256.663
R652 B.n966 B.n128 256.663
R653 B.n966 B.n127 256.663
R654 B.n966 B.n126 256.663
R655 B.n966 B.n125 256.663
R656 B.n966 B.n124 256.663
R657 B.n966 B.n123 256.663
R658 B.n966 B.n122 256.663
R659 B.n966 B.n121 256.663
R660 B.n966 B.n120 256.663
R661 B.n966 B.n119 256.663
R662 B.n966 B.n118 256.663
R663 B.n966 B.n117 256.663
R664 B.n966 B.n116 256.663
R665 B.n966 B.n115 256.663
R666 B.n966 B.n114 256.663
R667 B.n966 B.n113 256.663
R668 B.n966 B.n112 256.663
R669 B.n966 B.n111 256.663
R670 B.n966 B.n110 256.663
R671 B.n966 B.n109 256.663
R672 B.n966 B.n108 256.663
R673 B.n966 B.n107 256.663
R674 B.n966 B.n106 256.663
R675 B.n966 B.n105 256.663
R676 B.n966 B.n104 256.663
R677 B.n966 B.n103 256.663
R678 B.n966 B.n102 256.663
R679 B.n966 B.n101 256.663
R680 B.n966 B.n100 256.663
R681 B.n966 B.n99 256.663
R682 B.n966 B.n98 256.663
R683 B.n966 B.n97 256.663
R684 B.n966 B.n96 256.663
R685 B.n966 B.n95 256.663
R686 B.n966 B.n94 256.663
R687 B.n966 B.n93 256.663
R688 B.n966 B.n92 256.663
R689 B.n966 B.n91 256.663
R690 B.n529 B.n467 256.663
R691 B.n532 B.n467 256.663
R692 B.n538 B.n467 256.663
R693 B.n540 B.n467 256.663
R694 B.n546 B.n467 256.663
R695 B.n548 B.n467 256.663
R696 B.n554 B.n467 256.663
R697 B.n556 B.n467 256.663
R698 B.n562 B.n467 256.663
R699 B.n564 B.n467 256.663
R700 B.n570 B.n467 256.663
R701 B.n572 B.n467 256.663
R702 B.n578 B.n467 256.663
R703 B.n580 B.n467 256.663
R704 B.n586 B.n467 256.663
R705 B.n588 B.n467 256.663
R706 B.n594 B.n467 256.663
R707 B.n596 B.n467 256.663
R708 B.n602 B.n467 256.663
R709 B.n604 B.n467 256.663
R710 B.n610 B.n467 256.663
R711 B.n612 B.n467 256.663
R712 B.n618 B.n467 256.663
R713 B.n620 B.n467 256.663
R714 B.n626 B.n467 256.663
R715 B.n628 B.n467 256.663
R716 B.n635 B.n467 256.663
R717 B.n637 B.n467 256.663
R718 B.n643 B.n467 256.663
R719 B.n645 B.n467 256.663
R720 B.n652 B.n467 256.663
R721 B.n654 B.n467 256.663
R722 B.n660 B.n467 256.663
R723 B.n662 B.n467 256.663
R724 B.n668 B.n467 256.663
R725 B.n670 B.n467 256.663
R726 B.n676 B.n467 256.663
R727 B.n678 B.n467 256.663
R728 B.n684 B.n467 256.663
R729 B.n686 B.n467 256.663
R730 B.n692 B.n467 256.663
R731 B.n694 B.n467 256.663
R732 B.n700 B.n467 256.663
R733 B.n702 B.n467 256.663
R734 B.n708 B.n467 256.663
R735 B.n710 B.n467 256.663
R736 B.n716 B.n467 256.663
R737 B.n718 B.n467 256.663
R738 B.n724 B.n467 256.663
R739 B.n726 B.n467 256.663
R740 B.n732 B.n467 256.663
R741 B.n734 B.n467 256.663
R742 B.n740 B.n467 256.663
R743 B.n742 B.n467 256.663
R744 B.n748 B.n467 256.663
R745 B.n750 B.n467 256.663
R746 B.n1067 B.n1066 256.663
R747 B.n155 B.n154 163.367
R748 B.n159 B.n158 163.367
R749 B.n163 B.n162 163.367
R750 B.n167 B.n166 163.367
R751 B.n171 B.n170 163.367
R752 B.n175 B.n174 163.367
R753 B.n179 B.n178 163.367
R754 B.n183 B.n182 163.367
R755 B.n187 B.n186 163.367
R756 B.n191 B.n190 163.367
R757 B.n195 B.n194 163.367
R758 B.n199 B.n198 163.367
R759 B.n203 B.n202 163.367
R760 B.n207 B.n206 163.367
R761 B.n211 B.n210 163.367
R762 B.n215 B.n214 163.367
R763 B.n219 B.n218 163.367
R764 B.n223 B.n222 163.367
R765 B.n227 B.n226 163.367
R766 B.n231 B.n230 163.367
R767 B.n235 B.n234 163.367
R768 B.n239 B.n238 163.367
R769 B.n243 B.n242 163.367
R770 B.n247 B.n246 163.367
R771 B.n251 B.n250 163.367
R772 B.n255 B.n254 163.367
R773 B.n259 B.n258 163.367
R774 B.n263 B.n262 163.367
R775 B.n267 B.n266 163.367
R776 B.n271 B.n270 163.367
R777 B.n276 B.n275 163.367
R778 B.n280 B.n279 163.367
R779 B.n284 B.n283 163.367
R780 B.n288 B.n287 163.367
R781 B.n292 B.n291 163.367
R782 B.n296 B.n295 163.367
R783 B.n300 B.n299 163.367
R784 B.n304 B.n303 163.367
R785 B.n308 B.n307 163.367
R786 B.n312 B.n311 163.367
R787 B.n316 B.n315 163.367
R788 B.n320 B.n319 163.367
R789 B.n324 B.n323 163.367
R790 B.n328 B.n327 163.367
R791 B.n332 B.n331 163.367
R792 B.n336 B.n335 163.367
R793 B.n340 B.n339 163.367
R794 B.n344 B.n343 163.367
R795 B.n348 B.n347 163.367
R796 B.n352 B.n351 163.367
R797 B.n356 B.n355 163.367
R798 B.n360 B.n359 163.367
R799 B.n364 B.n363 163.367
R800 B.n368 B.n367 163.367
R801 B.n372 B.n371 163.367
R802 B.n965 B.n147 163.367
R803 B.n755 B.n462 163.367
R804 B.n763 B.n462 163.367
R805 B.n763 B.n460 163.367
R806 B.n767 B.n460 163.367
R807 B.n767 B.n454 163.367
R808 B.n775 B.n454 163.367
R809 B.n775 B.n452 163.367
R810 B.n779 B.n452 163.367
R811 B.n779 B.n446 163.367
R812 B.n787 B.n446 163.367
R813 B.n787 B.n444 163.367
R814 B.n791 B.n444 163.367
R815 B.n791 B.n438 163.367
R816 B.n799 B.n438 163.367
R817 B.n799 B.n436 163.367
R818 B.n803 B.n436 163.367
R819 B.n803 B.n430 163.367
R820 B.n811 B.n430 163.367
R821 B.n811 B.n428 163.367
R822 B.n815 B.n428 163.367
R823 B.n815 B.n423 163.367
R824 B.n824 B.n423 163.367
R825 B.n824 B.n421 163.367
R826 B.n828 B.n421 163.367
R827 B.n828 B.n415 163.367
R828 B.n836 B.n415 163.367
R829 B.n836 B.n413 163.367
R830 B.n840 B.n413 163.367
R831 B.n840 B.n406 163.367
R832 B.n848 B.n406 163.367
R833 B.n848 B.n404 163.367
R834 B.n852 B.n404 163.367
R835 B.n852 B.n399 163.367
R836 B.n860 B.n399 163.367
R837 B.n860 B.n397 163.367
R838 B.n864 B.n397 163.367
R839 B.n864 B.n391 163.367
R840 B.n872 B.n391 163.367
R841 B.n872 B.n389 163.367
R842 B.n876 B.n389 163.367
R843 B.n876 B.n384 163.367
R844 B.n885 B.n384 163.367
R845 B.n885 B.n382 163.367
R846 B.n890 B.n382 163.367
R847 B.n890 B.n376 163.367
R848 B.n898 B.n376 163.367
R849 B.n899 B.n898 163.367
R850 B.n899 B.n5 163.367
R851 B.n6 B.n5 163.367
R852 B.n7 B.n6 163.367
R853 B.n905 B.n7 163.367
R854 B.n906 B.n905 163.367
R855 B.n906 B.n13 163.367
R856 B.n14 B.n13 163.367
R857 B.n15 B.n14 163.367
R858 B.n911 B.n15 163.367
R859 B.n911 B.n20 163.367
R860 B.n21 B.n20 163.367
R861 B.n22 B.n21 163.367
R862 B.n916 B.n22 163.367
R863 B.n916 B.n27 163.367
R864 B.n28 B.n27 163.367
R865 B.n29 B.n28 163.367
R866 B.n921 B.n29 163.367
R867 B.n921 B.n34 163.367
R868 B.n35 B.n34 163.367
R869 B.n36 B.n35 163.367
R870 B.n926 B.n36 163.367
R871 B.n926 B.n41 163.367
R872 B.n42 B.n41 163.367
R873 B.n43 B.n42 163.367
R874 B.n931 B.n43 163.367
R875 B.n931 B.n48 163.367
R876 B.n49 B.n48 163.367
R877 B.n50 B.n49 163.367
R878 B.n936 B.n50 163.367
R879 B.n936 B.n55 163.367
R880 B.n56 B.n55 163.367
R881 B.n57 B.n56 163.367
R882 B.n941 B.n57 163.367
R883 B.n941 B.n62 163.367
R884 B.n63 B.n62 163.367
R885 B.n64 B.n63 163.367
R886 B.n946 B.n64 163.367
R887 B.n946 B.n69 163.367
R888 B.n70 B.n69 163.367
R889 B.n71 B.n70 163.367
R890 B.n951 B.n71 163.367
R891 B.n951 B.n76 163.367
R892 B.n77 B.n76 163.367
R893 B.n78 B.n77 163.367
R894 B.n956 B.n78 163.367
R895 B.n956 B.n83 163.367
R896 B.n84 B.n83 163.367
R897 B.n85 B.n84 163.367
R898 B.n961 B.n85 163.367
R899 B.n961 B.n90 163.367
R900 B.n531 B.n530 163.367
R901 B.n533 B.n531 163.367
R902 B.n537 B.n526 163.367
R903 B.n541 B.n539 163.367
R904 B.n545 B.n524 163.367
R905 B.n549 B.n547 163.367
R906 B.n553 B.n522 163.367
R907 B.n557 B.n555 163.367
R908 B.n561 B.n520 163.367
R909 B.n565 B.n563 163.367
R910 B.n569 B.n518 163.367
R911 B.n573 B.n571 163.367
R912 B.n577 B.n516 163.367
R913 B.n581 B.n579 163.367
R914 B.n585 B.n514 163.367
R915 B.n589 B.n587 163.367
R916 B.n593 B.n512 163.367
R917 B.n597 B.n595 163.367
R918 B.n601 B.n510 163.367
R919 B.n605 B.n603 163.367
R920 B.n609 B.n508 163.367
R921 B.n613 B.n611 163.367
R922 B.n617 B.n506 163.367
R923 B.n621 B.n619 163.367
R924 B.n625 B.n504 163.367
R925 B.n629 B.n627 163.367
R926 B.n634 B.n500 163.367
R927 B.n638 B.n636 163.367
R928 B.n642 B.n498 163.367
R929 B.n646 B.n644 163.367
R930 B.n651 B.n494 163.367
R931 B.n655 B.n653 163.367
R932 B.n659 B.n492 163.367
R933 B.n663 B.n661 163.367
R934 B.n667 B.n490 163.367
R935 B.n671 B.n669 163.367
R936 B.n675 B.n488 163.367
R937 B.n679 B.n677 163.367
R938 B.n683 B.n486 163.367
R939 B.n687 B.n685 163.367
R940 B.n691 B.n484 163.367
R941 B.n695 B.n693 163.367
R942 B.n699 B.n482 163.367
R943 B.n703 B.n701 163.367
R944 B.n707 B.n480 163.367
R945 B.n711 B.n709 163.367
R946 B.n715 B.n478 163.367
R947 B.n719 B.n717 163.367
R948 B.n723 B.n476 163.367
R949 B.n727 B.n725 163.367
R950 B.n731 B.n474 163.367
R951 B.n735 B.n733 163.367
R952 B.n739 B.n472 163.367
R953 B.n743 B.n741 163.367
R954 B.n747 B.n470 163.367
R955 B.n751 B.n749 163.367
R956 B.n757 B.n464 163.367
R957 B.n761 B.n464 163.367
R958 B.n761 B.n458 163.367
R959 B.n769 B.n458 163.367
R960 B.n769 B.n456 163.367
R961 B.n773 B.n456 163.367
R962 B.n773 B.n450 163.367
R963 B.n781 B.n450 163.367
R964 B.n781 B.n448 163.367
R965 B.n785 B.n448 163.367
R966 B.n785 B.n442 163.367
R967 B.n793 B.n442 163.367
R968 B.n793 B.n440 163.367
R969 B.n797 B.n440 163.367
R970 B.n797 B.n434 163.367
R971 B.n805 B.n434 163.367
R972 B.n805 B.n432 163.367
R973 B.n809 B.n432 163.367
R974 B.n809 B.n426 163.367
R975 B.n818 B.n426 163.367
R976 B.n818 B.n424 163.367
R977 B.n822 B.n424 163.367
R978 B.n822 B.n419 163.367
R979 B.n830 B.n419 163.367
R980 B.n830 B.n417 163.367
R981 B.n834 B.n417 163.367
R982 B.n834 B.n411 163.367
R983 B.n842 B.n411 163.367
R984 B.n842 B.n409 163.367
R985 B.n846 B.n409 163.367
R986 B.n846 B.n403 163.367
R987 B.n854 B.n403 163.367
R988 B.n854 B.n401 163.367
R989 B.n858 B.n401 163.367
R990 B.n858 B.n395 163.367
R991 B.n866 B.n395 163.367
R992 B.n866 B.n393 163.367
R993 B.n870 B.n393 163.367
R994 B.n870 B.n387 163.367
R995 B.n879 B.n387 163.367
R996 B.n879 B.n385 163.367
R997 B.n883 B.n385 163.367
R998 B.n883 B.n380 163.367
R999 B.n892 B.n380 163.367
R1000 B.n892 B.n378 163.367
R1001 B.n896 B.n378 163.367
R1002 B.n896 B.n3 163.367
R1003 B.n1065 B.n3 163.367
R1004 B.n1061 B.n2 163.367
R1005 B.n1061 B.n1060 163.367
R1006 B.n1060 B.n9 163.367
R1007 B.n1056 B.n9 163.367
R1008 B.n1056 B.n11 163.367
R1009 B.n1052 B.n11 163.367
R1010 B.n1052 B.n16 163.367
R1011 B.n1048 B.n16 163.367
R1012 B.n1048 B.n18 163.367
R1013 B.n1044 B.n18 163.367
R1014 B.n1044 B.n24 163.367
R1015 B.n1040 B.n24 163.367
R1016 B.n1040 B.n26 163.367
R1017 B.n1036 B.n26 163.367
R1018 B.n1036 B.n31 163.367
R1019 B.n1032 B.n31 163.367
R1020 B.n1032 B.n33 163.367
R1021 B.n1028 B.n33 163.367
R1022 B.n1028 B.n38 163.367
R1023 B.n1024 B.n38 163.367
R1024 B.n1024 B.n40 163.367
R1025 B.n1020 B.n40 163.367
R1026 B.n1020 B.n45 163.367
R1027 B.n1016 B.n45 163.367
R1028 B.n1016 B.n47 163.367
R1029 B.n1012 B.n47 163.367
R1030 B.n1012 B.n51 163.367
R1031 B.n1008 B.n51 163.367
R1032 B.n1008 B.n53 163.367
R1033 B.n1004 B.n53 163.367
R1034 B.n1004 B.n59 163.367
R1035 B.n1000 B.n59 163.367
R1036 B.n1000 B.n61 163.367
R1037 B.n996 B.n61 163.367
R1038 B.n996 B.n66 163.367
R1039 B.n992 B.n66 163.367
R1040 B.n992 B.n68 163.367
R1041 B.n988 B.n68 163.367
R1042 B.n988 B.n73 163.367
R1043 B.n984 B.n73 163.367
R1044 B.n984 B.n75 163.367
R1045 B.n980 B.n75 163.367
R1046 B.n980 B.n80 163.367
R1047 B.n976 B.n80 163.367
R1048 B.n976 B.n82 163.367
R1049 B.n972 B.n82 163.367
R1050 B.n972 B.n87 163.367
R1051 B.n968 B.n87 163.367
R1052 B.n91 B.n89 71.676
R1053 B.n155 B.n92 71.676
R1054 B.n159 B.n93 71.676
R1055 B.n163 B.n94 71.676
R1056 B.n167 B.n95 71.676
R1057 B.n171 B.n96 71.676
R1058 B.n175 B.n97 71.676
R1059 B.n179 B.n98 71.676
R1060 B.n183 B.n99 71.676
R1061 B.n187 B.n100 71.676
R1062 B.n191 B.n101 71.676
R1063 B.n195 B.n102 71.676
R1064 B.n199 B.n103 71.676
R1065 B.n203 B.n104 71.676
R1066 B.n207 B.n105 71.676
R1067 B.n211 B.n106 71.676
R1068 B.n215 B.n107 71.676
R1069 B.n219 B.n108 71.676
R1070 B.n223 B.n109 71.676
R1071 B.n227 B.n110 71.676
R1072 B.n231 B.n111 71.676
R1073 B.n235 B.n112 71.676
R1074 B.n239 B.n113 71.676
R1075 B.n243 B.n114 71.676
R1076 B.n247 B.n115 71.676
R1077 B.n251 B.n116 71.676
R1078 B.n255 B.n117 71.676
R1079 B.n259 B.n118 71.676
R1080 B.n263 B.n119 71.676
R1081 B.n267 B.n120 71.676
R1082 B.n271 B.n121 71.676
R1083 B.n276 B.n122 71.676
R1084 B.n280 B.n123 71.676
R1085 B.n284 B.n124 71.676
R1086 B.n288 B.n125 71.676
R1087 B.n292 B.n126 71.676
R1088 B.n296 B.n127 71.676
R1089 B.n300 B.n128 71.676
R1090 B.n304 B.n129 71.676
R1091 B.n308 B.n130 71.676
R1092 B.n312 B.n131 71.676
R1093 B.n316 B.n132 71.676
R1094 B.n320 B.n133 71.676
R1095 B.n324 B.n134 71.676
R1096 B.n328 B.n135 71.676
R1097 B.n332 B.n136 71.676
R1098 B.n336 B.n137 71.676
R1099 B.n340 B.n138 71.676
R1100 B.n344 B.n139 71.676
R1101 B.n348 B.n140 71.676
R1102 B.n352 B.n141 71.676
R1103 B.n356 B.n142 71.676
R1104 B.n360 B.n143 71.676
R1105 B.n364 B.n144 71.676
R1106 B.n368 B.n145 71.676
R1107 B.n372 B.n146 71.676
R1108 B.n147 B.n146 71.676
R1109 B.n371 B.n145 71.676
R1110 B.n367 B.n144 71.676
R1111 B.n363 B.n143 71.676
R1112 B.n359 B.n142 71.676
R1113 B.n355 B.n141 71.676
R1114 B.n351 B.n140 71.676
R1115 B.n347 B.n139 71.676
R1116 B.n343 B.n138 71.676
R1117 B.n339 B.n137 71.676
R1118 B.n335 B.n136 71.676
R1119 B.n331 B.n135 71.676
R1120 B.n327 B.n134 71.676
R1121 B.n323 B.n133 71.676
R1122 B.n319 B.n132 71.676
R1123 B.n315 B.n131 71.676
R1124 B.n311 B.n130 71.676
R1125 B.n307 B.n129 71.676
R1126 B.n303 B.n128 71.676
R1127 B.n299 B.n127 71.676
R1128 B.n295 B.n126 71.676
R1129 B.n291 B.n125 71.676
R1130 B.n287 B.n124 71.676
R1131 B.n283 B.n123 71.676
R1132 B.n279 B.n122 71.676
R1133 B.n275 B.n121 71.676
R1134 B.n270 B.n120 71.676
R1135 B.n266 B.n119 71.676
R1136 B.n262 B.n118 71.676
R1137 B.n258 B.n117 71.676
R1138 B.n254 B.n116 71.676
R1139 B.n250 B.n115 71.676
R1140 B.n246 B.n114 71.676
R1141 B.n242 B.n113 71.676
R1142 B.n238 B.n112 71.676
R1143 B.n234 B.n111 71.676
R1144 B.n230 B.n110 71.676
R1145 B.n226 B.n109 71.676
R1146 B.n222 B.n108 71.676
R1147 B.n218 B.n107 71.676
R1148 B.n214 B.n106 71.676
R1149 B.n210 B.n105 71.676
R1150 B.n206 B.n104 71.676
R1151 B.n202 B.n103 71.676
R1152 B.n198 B.n102 71.676
R1153 B.n194 B.n101 71.676
R1154 B.n190 B.n100 71.676
R1155 B.n186 B.n99 71.676
R1156 B.n182 B.n98 71.676
R1157 B.n178 B.n97 71.676
R1158 B.n174 B.n96 71.676
R1159 B.n170 B.n95 71.676
R1160 B.n166 B.n94 71.676
R1161 B.n162 B.n93 71.676
R1162 B.n158 B.n92 71.676
R1163 B.n154 B.n91 71.676
R1164 B.n529 B.n466 71.676
R1165 B.n533 B.n532 71.676
R1166 B.n538 B.n537 71.676
R1167 B.n541 B.n540 71.676
R1168 B.n546 B.n545 71.676
R1169 B.n549 B.n548 71.676
R1170 B.n554 B.n553 71.676
R1171 B.n557 B.n556 71.676
R1172 B.n562 B.n561 71.676
R1173 B.n565 B.n564 71.676
R1174 B.n570 B.n569 71.676
R1175 B.n573 B.n572 71.676
R1176 B.n578 B.n577 71.676
R1177 B.n581 B.n580 71.676
R1178 B.n586 B.n585 71.676
R1179 B.n589 B.n588 71.676
R1180 B.n594 B.n593 71.676
R1181 B.n597 B.n596 71.676
R1182 B.n602 B.n601 71.676
R1183 B.n605 B.n604 71.676
R1184 B.n610 B.n609 71.676
R1185 B.n613 B.n612 71.676
R1186 B.n618 B.n617 71.676
R1187 B.n621 B.n620 71.676
R1188 B.n626 B.n625 71.676
R1189 B.n629 B.n628 71.676
R1190 B.n635 B.n634 71.676
R1191 B.n638 B.n637 71.676
R1192 B.n643 B.n642 71.676
R1193 B.n646 B.n645 71.676
R1194 B.n652 B.n651 71.676
R1195 B.n655 B.n654 71.676
R1196 B.n660 B.n659 71.676
R1197 B.n663 B.n662 71.676
R1198 B.n668 B.n667 71.676
R1199 B.n671 B.n670 71.676
R1200 B.n676 B.n675 71.676
R1201 B.n679 B.n678 71.676
R1202 B.n684 B.n683 71.676
R1203 B.n687 B.n686 71.676
R1204 B.n692 B.n691 71.676
R1205 B.n695 B.n694 71.676
R1206 B.n700 B.n699 71.676
R1207 B.n703 B.n702 71.676
R1208 B.n708 B.n707 71.676
R1209 B.n711 B.n710 71.676
R1210 B.n716 B.n715 71.676
R1211 B.n719 B.n718 71.676
R1212 B.n724 B.n723 71.676
R1213 B.n727 B.n726 71.676
R1214 B.n732 B.n731 71.676
R1215 B.n735 B.n734 71.676
R1216 B.n740 B.n739 71.676
R1217 B.n743 B.n742 71.676
R1218 B.n748 B.n747 71.676
R1219 B.n751 B.n750 71.676
R1220 B.n530 B.n529 71.676
R1221 B.n532 B.n526 71.676
R1222 B.n539 B.n538 71.676
R1223 B.n540 B.n524 71.676
R1224 B.n547 B.n546 71.676
R1225 B.n548 B.n522 71.676
R1226 B.n555 B.n554 71.676
R1227 B.n556 B.n520 71.676
R1228 B.n563 B.n562 71.676
R1229 B.n564 B.n518 71.676
R1230 B.n571 B.n570 71.676
R1231 B.n572 B.n516 71.676
R1232 B.n579 B.n578 71.676
R1233 B.n580 B.n514 71.676
R1234 B.n587 B.n586 71.676
R1235 B.n588 B.n512 71.676
R1236 B.n595 B.n594 71.676
R1237 B.n596 B.n510 71.676
R1238 B.n603 B.n602 71.676
R1239 B.n604 B.n508 71.676
R1240 B.n611 B.n610 71.676
R1241 B.n612 B.n506 71.676
R1242 B.n619 B.n618 71.676
R1243 B.n620 B.n504 71.676
R1244 B.n627 B.n626 71.676
R1245 B.n628 B.n500 71.676
R1246 B.n636 B.n635 71.676
R1247 B.n637 B.n498 71.676
R1248 B.n644 B.n643 71.676
R1249 B.n645 B.n494 71.676
R1250 B.n653 B.n652 71.676
R1251 B.n654 B.n492 71.676
R1252 B.n661 B.n660 71.676
R1253 B.n662 B.n490 71.676
R1254 B.n669 B.n668 71.676
R1255 B.n670 B.n488 71.676
R1256 B.n677 B.n676 71.676
R1257 B.n678 B.n486 71.676
R1258 B.n685 B.n684 71.676
R1259 B.n686 B.n484 71.676
R1260 B.n693 B.n692 71.676
R1261 B.n694 B.n482 71.676
R1262 B.n701 B.n700 71.676
R1263 B.n702 B.n480 71.676
R1264 B.n709 B.n708 71.676
R1265 B.n710 B.n478 71.676
R1266 B.n717 B.n716 71.676
R1267 B.n718 B.n476 71.676
R1268 B.n725 B.n724 71.676
R1269 B.n726 B.n474 71.676
R1270 B.n733 B.n732 71.676
R1271 B.n734 B.n472 71.676
R1272 B.n741 B.n740 71.676
R1273 B.n742 B.n470 71.676
R1274 B.n749 B.n748 71.676
R1275 B.n750 B.n468 71.676
R1276 B.n1066 B.n1065 71.676
R1277 B.n1066 B.n2 71.676
R1278 B.n151 B.n150 66.3278
R1279 B.n149 B.n148 66.3278
R1280 B.n496 B.n495 66.3278
R1281 B.n502 B.n501 66.3278
R1282 B.n756 B.n467 60.2088
R1283 B.n967 B.n966 60.2088
R1284 B.n152 B.n151 59.5399
R1285 B.n273 B.n149 59.5399
R1286 B.n649 B.n496 59.5399
R1287 B.n631 B.n502 59.5399
R1288 B.n756 B.n463 36.232
R1289 B.n762 B.n463 36.232
R1290 B.n762 B.n459 36.232
R1291 B.n768 B.n459 36.232
R1292 B.n768 B.n455 36.232
R1293 B.n774 B.n455 36.232
R1294 B.n774 B.n451 36.232
R1295 B.n780 B.n451 36.232
R1296 B.n786 B.n447 36.232
R1297 B.n786 B.n443 36.232
R1298 B.n792 B.n443 36.232
R1299 B.n792 B.n439 36.232
R1300 B.n798 B.n439 36.232
R1301 B.n798 B.n435 36.232
R1302 B.n804 B.n435 36.232
R1303 B.n804 B.n431 36.232
R1304 B.n810 B.n431 36.232
R1305 B.n810 B.n427 36.232
R1306 B.n817 B.n427 36.232
R1307 B.n817 B.n816 36.232
R1308 B.n823 B.n420 36.232
R1309 B.n829 B.n420 36.232
R1310 B.n829 B.n416 36.232
R1311 B.n835 B.n416 36.232
R1312 B.n835 B.n412 36.232
R1313 B.n841 B.n412 36.232
R1314 B.n841 B.n407 36.232
R1315 B.n847 B.n407 36.232
R1316 B.n847 B.n408 36.232
R1317 B.n853 B.n400 36.232
R1318 B.n859 B.n400 36.232
R1319 B.n859 B.n396 36.232
R1320 B.n865 B.n396 36.232
R1321 B.n865 B.n392 36.232
R1322 B.n871 B.n392 36.232
R1323 B.n871 B.n388 36.232
R1324 B.n878 B.n388 36.232
R1325 B.n878 B.n877 36.232
R1326 B.n884 B.n381 36.232
R1327 B.n891 B.n381 36.232
R1328 B.n891 B.n377 36.232
R1329 B.n897 B.n377 36.232
R1330 B.n897 B.n4 36.232
R1331 B.n1064 B.n4 36.232
R1332 B.n1064 B.n1063 36.232
R1333 B.n1063 B.n1062 36.232
R1334 B.n1062 B.n8 36.232
R1335 B.n12 B.n8 36.232
R1336 B.n1055 B.n12 36.232
R1337 B.n1055 B.n1054 36.232
R1338 B.n1054 B.n1053 36.232
R1339 B.n1047 B.n19 36.232
R1340 B.n1047 B.n1046 36.232
R1341 B.n1046 B.n1045 36.232
R1342 B.n1045 B.n23 36.232
R1343 B.n1039 B.n23 36.232
R1344 B.n1039 B.n1038 36.232
R1345 B.n1038 B.n1037 36.232
R1346 B.n1037 B.n30 36.232
R1347 B.n1031 B.n30 36.232
R1348 B.n1030 B.n1029 36.232
R1349 B.n1029 B.n37 36.232
R1350 B.n1023 B.n37 36.232
R1351 B.n1023 B.n1022 36.232
R1352 B.n1022 B.n1021 36.232
R1353 B.n1021 B.n44 36.232
R1354 B.n1015 B.n44 36.232
R1355 B.n1015 B.n1014 36.232
R1356 B.n1014 B.n1013 36.232
R1357 B.n1007 B.n54 36.232
R1358 B.n1007 B.n1006 36.232
R1359 B.n1006 B.n1005 36.232
R1360 B.n1005 B.n58 36.232
R1361 B.n999 B.n58 36.232
R1362 B.n999 B.n998 36.232
R1363 B.n998 B.n997 36.232
R1364 B.n997 B.n65 36.232
R1365 B.n991 B.n65 36.232
R1366 B.n991 B.n990 36.232
R1367 B.n990 B.n989 36.232
R1368 B.n989 B.n72 36.232
R1369 B.n983 B.n982 36.232
R1370 B.n982 B.n981 36.232
R1371 B.n981 B.n79 36.232
R1372 B.n975 B.n79 36.232
R1373 B.n975 B.n974 36.232
R1374 B.n974 B.n973 36.232
R1375 B.n973 B.n86 36.232
R1376 B.n967 B.n86 36.232
R1377 B.n877 B.t3 31.4367
R1378 B.n19 B.t1 31.4367
R1379 B.n408 B.t2 29.3054
R1380 B.t4 B.n1030 29.3054
R1381 B.n758 B.n465 28.8785
R1382 B.n754 B.n753 28.8785
R1383 B.n964 B.n963 28.8785
R1384 B.n969 B.n88 28.8785
R1385 B.n816 B.t0 27.1742
R1386 B.n54 B.t5 27.1742
R1387 B.t11 B.n447 18.6491
R1388 B.t7 B.n72 18.6491
R1389 B B.n1067 18.0485
R1390 B.n780 B.t11 17.5834
R1391 B.n983 B.t7 17.5834
R1392 B.n759 B.n758 10.6151
R1393 B.n760 B.n759 10.6151
R1394 B.n760 B.n457 10.6151
R1395 B.n770 B.n457 10.6151
R1396 B.n771 B.n770 10.6151
R1397 B.n772 B.n771 10.6151
R1398 B.n772 B.n449 10.6151
R1399 B.n782 B.n449 10.6151
R1400 B.n783 B.n782 10.6151
R1401 B.n784 B.n783 10.6151
R1402 B.n784 B.n441 10.6151
R1403 B.n794 B.n441 10.6151
R1404 B.n795 B.n794 10.6151
R1405 B.n796 B.n795 10.6151
R1406 B.n796 B.n433 10.6151
R1407 B.n806 B.n433 10.6151
R1408 B.n807 B.n806 10.6151
R1409 B.n808 B.n807 10.6151
R1410 B.n808 B.n425 10.6151
R1411 B.n819 B.n425 10.6151
R1412 B.n820 B.n819 10.6151
R1413 B.n821 B.n820 10.6151
R1414 B.n821 B.n418 10.6151
R1415 B.n831 B.n418 10.6151
R1416 B.n832 B.n831 10.6151
R1417 B.n833 B.n832 10.6151
R1418 B.n833 B.n410 10.6151
R1419 B.n843 B.n410 10.6151
R1420 B.n844 B.n843 10.6151
R1421 B.n845 B.n844 10.6151
R1422 B.n845 B.n402 10.6151
R1423 B.n855 B.n402 10.6151
R1424 B.n856 B.n855 10.6151
R1425 B.n857 B.n856 10.6151
R1426 B.n857 B.n394 10.6151
R1427 B.n867 B.n394 10.6151
R1428 B.n868 B.n867 10.6151
R1429 B.n869 B.n868 10.6151
R1430 B.n869 B.n386 10.6151
R1431 B.n880 B.n386 10.6151
R1432 B.n881 B.n880 10.6151
R1433 B.n882 B.n881 10.6151
R1434 B.n882 B.n379 10.6151
R1435 B.n893 B.n379 10.6151
R1436 B.n894 B.n893 10.6151
R1437 B.n895 B.n894 10.6151
R1438 B.n895 B.n0 10.6151
R1439 B.n528 B.n465 10.6151
R1440 B.n528 B.n527 10.6151
R1441 B.n534 B.n527 10.6151
R1442 B.n535 B.n534 10.6151
R1443 B.n536 B.n535 10.6151
R1444 B.n536 B.n525 10.6151
R1445 B.n542 B.n525 10.6151
R1446 B.n543 B.n542 10.6151
R1447 B.n544 B.n543 10.6151
R1448 B.n544 B.n523 10.6151
R1449 B.n550 B.n523 10.6151
R1450 B.n551 B.n550 10.6151
R1451 B.n552 B.n551 10.6151
R1452 B.n552 B.n521 10.6151
R1453 B.n558 B.n521 10.6151
R1454 B.n559 B.n558 10.6151
R1455 B.n560 B.n559 10.6151
R1456 B.n560 B.n519 10.6151
R1457 B.n566 B.n519 10.6151
R1458 B.n567 B.n566 10.6151
R1459 B.n568 B.n567 10.6151
R1460 B.n568 B.n517 10.6151
R1461 B.n574 B.n517 10.6151
R1462 B.n575 B.n574 10.6151
R1463 B.n576 B.n575 10.6151
R1464 B.n576 B.n515 10.6151
R1465 B.n582 B.n515 10.6151
R1466 B.n583 B.n582 10.6151
R1467 B.n584 B.n583 10.6151
R1468 B.n584 B.n513 10.6151
R1469 B.n590 B.n513 10.6151
R1470 B.n591 B.n590 10.6151
R1471 B.n592 B.n591 10.6151
R1472 B.n592 B.n511 10.6151
R1473 B.n598 B.n511 10.6151
R1474 B.n599 B.n598 10.6151
R1475 B.n600 B.n599 10.6151
R1476 B.n600 B.n509 10.6151
R1477 B.n606 B.n509 10.6151
R1478 B.n607 B.n606 10.6151
R1479 B.n608 B.n607 10.6151
R1480 B.n608 B.n507 10.6151
R1481 B.n614 B.n507 10.6151
R1482 B.n615 B.n614 10.6151
R1483 B.n616 B.n615 10.6151
R1484 B.n616 B.n505 10.6151
R1485 B.n622 B.n505 10.6151
R1486 B.n623 B.n622 10.6151
R1487 B.n624 B.n623 10.6151
R1488 B.n624 B.n503 10.6151
R1489 B.n630 B.n503 10.6151
R1490 B.n633 B.n632 10.6151
R1491 B.n633 B.n499 10.6151
R1492 B.n639 B.n499 10.6151
R1493 B.n640 B.n639 10.6151
R1494 B.n641 B.n640 10.6151
R1495 B.n641 B.n497 10.6151
R1496 B.n647 B.n497 10.6151
R1497 B.n648 B.n647 10.6151
R1498 B.n650 B.n493 10.6151
R1499 B.n656 B.n493 10.6151
R1500 B.n657 B.n656 10.6151
R1501 B.n658 B.n657 10.6151
R1502 B.n658 B.n491 10.6151
R1503 B.n664 B.n491 10.6151
R1504 B.n665 B.n664 10.6151
R1505 B.n666 B.n665 10.6151
R1506 B.n666 B.n489 10.6151
R1507 B.n672 B.n489 10.6151
R1508 B.n673 B.n672 10.6151
R1509 B.n674 B.n673 10.6151
R1510 B.n674 B.n487 10.6151
R1511 B.n680 B.n487 10.6151
R1512 B.n681 B.n680 10.6151
R1513 B.n682 B.n681 10.6151
R1514 B.n682 B.n485 10.6151
R1515 B.n688 B.n485 10.6151
R1516 B.n689 B.n688 10.6151
R1517 B.n690 B.n689 10.6151
R1518 B.n690 B.n483 10.6151
R1519 B.n696 B.n483 10.6151
R1520 B.n697 B.n696 10.6151
R1521 B.n698 B.n697 10.6151
R1522 B.n698 B.n481 10.6151
R1523 B.n704 B.n481 10.6151
R1524 B.n705 B.n704 10.6151
R1525 B.n706 B.n705 10.6151
R1526 B.n706 B.n479 10.6151
R1527 B.n712 B.n479 10.6151
R1528 B.n713 B.n712 10.6151
R1529 B.n714 B.n713 10.6151
R1530 B.n714 B.n477 10.6151
R1531 B.n720 B.n477 10.6151
R1532 B.n721 B.n720 10.6151
R1533 B.n722 B.n721 10.6151
R1534 B.n722 B.n475 10.6151
R1535 B.n728 B.n475 10.6151
R1536 B.n729 B.n728 10.6151
R1537 B.n730 B.n729 10.6151
R1538 B.n730 B.n473 10.6151
R1539 B.n736 B.n473 10.6151
R1540 B.n737 B.n736 10.6151
R1541 B.n738 B.n737 10.6151
R1542 B.n738 B.n471 10.6151
R1543 B.n744 B.n471 10.6151
R1544 B.n745 B.n744 10.6151
R1545 B.n746 B.n745 10.6151
R1546 B.n746 B.n469 10.6151
R1547 B.n752 B.n469 10.6151
R1548 B.n753 B.n752 10.6151
R1549 B.n754 B.n461 10.6151
R1550 B.n764 B.n461 10.6151
R1551 B.n765 B.n764 10.6151
R1552 B.n766 B.n765 10.6151
R1553 B.n766 B.n453 10.6151
R1554 B.n776 B.n453 10.6151
R1555 B.n777 B.n776 10.6151
R1556 B.n778 B.n777 10.6151
R1557 B.n778 B.n445 10.6151
R1558 B.n788 B.n445 10.6151
R1559 B.n789 B.n788 10.6151
R1560 B.n790 B.n789 10.6151
R1561 B.n790 B.n437 10.6151
R1562 B.n800 B.n437 10.6151
R1563 B.n801 B.n800 10.6151
R1564 B.n802 B.n801 10.6151
R1565 B.n802 B.n429 10.6151
R1566 B.n812 B.n429 10.6151
R1567 B.n813 B.n812 10.6151
R1568 B.n814 B.n813 10.6151
R1569 B.n814 B.n422 10.6151
R1570 B.n825 B.n422 10.6151
R1571 B.n826 B.n825 10.6151
R1572 B.n827 B.n826 10.6151
R1573 B.n827 B.n414 10.6151
R1574 B.n837 B.n414 10.6151
R1575 B.n838 B.n837 10.6151
R1576 B.n839 B.n838 10.6151
R1577 B.n839 B.n405 10.6151
R1578 B.n849 B.n405 10.6151
R1579 B.n850 B.n849 10.6151
R1580 B.n851 B.n850 10.6151
R1581 B.n851 B.n398 10.6151
R1582 B.n861 B.n398 10.6151
R1583 B.n862 B.n861 10.6151
R1584 B.n863 B.n862 10.6151
R1585 B.n863 B.n390 10.6151
R1586 B.n873 B.n390 10.6151
R1587 B.n874 B.n873 10.6151
R1588 B.n875 B.n874 10.6151
R1589 B.n875 B.n383 10.6151
R1590 B.n886 B.n383 10.6151
R1591 B.n887 B.n886 10.6151
R1592 B.n889 B.n887 10.6151
R1593 B.n889 B.n888 10.6151
R1594 B.n888 B.n375 10.6151
R1595 B.n900 B.n375 10.6151
R1596 B.n901 B.n900 10.6151
R1597 B.n902 B.n901 10.6151
R1598 B.n903 B.n902 10.6151
R1599 B.n904 B.n903 10.6151
R1600 B.n907 B.n904 10.6151
R1601 B.n908 B.n907 10.6151
R1602 B.n909 B.n908 10.6151
R1603 B.n910 B.n909 10.6151
R1604 B.n912 B.n910 10.6151
R1605 B.n913 B.n912 10.6151
R1606 B.n914 B.n913 10.6151
R1607 B.n915 B.n914 10.6151
R1608 B.n917 B.n915 10.6151
R1609 B.n918 B.n917 10.6151
R1610 B.n919 B.n918 10.6151
R1611 B.n920 B.n919 10.6151
R1612 B.n922 B.n920 10.6151
R1613 B.n923 B.n922 10.6151
R1614 B.n924 B.n923 10.6151
R1615 B.n925 B.n924 10.6151
R1616 B.n927 B.n925 10.6151
R1617 B.n928 B.n927 10.6151
R1618 B.n929 B.n928 10.6151
R1619 B.n930 B.n929 10.6151
R1620 B.n932 B.n930 10.6151
R1621 B.n933 B.n932 10.6151
R1622 B.n934 B.n933 10.6151
R1623 B.n935 B.n934 10.6151
R1624 B.n937 B.n935 10.6151
R1625 B.n938 B.n937 10.6151
R1626 B.n939 B.n938 10.6151
R1627 B.n940 B.n939 10.6151
R1628 B.n942 B.n940 10.6151
R1629 B.n943 B.n942 10.6151
R1630 B.n944 B.n943 10.6151
R1631 B.n945 B.n944 10.6151
R1632 B.n947 B.n945 10.6151
R1633 B.n948 B.n947 10.6151
R1634 B.n949 B.n948 10.6151
R1635 B.n950 B.n949 10.6151
R1636 B.n952 B.n950 10.6151
R1637 B.n953 B.n952 10.6151
R1638 B.n954 B.n953 10.6151
R1639 B.n955 B.n954 10.6151
R1640 B.n957 B.n955 10.6151
R1641 B.n958 B.n957 10.6151
R1642 B.n959 B.n958 10.6151
R1643 B.n960 B.n959 10.6151
R1644 B.n962 B.n960 10.6151
R1645 B.n963 B.n962 10.6151
R1646 B.n1059 B.n1 10.6151
R1647 B.n1059 B.n1058 10.6151
R1648 B.n1058 B.n1057 10.6151
R1649 B.n1057 B.n10 10.6151
R1650 B.n1051 B.n10 10.6151
R1651 B.n1051 B.n1050 10.6151
R1652 B.n1050 B.n1049 10.6151
R1653 B.n1049 B.n17 10.6151
R1654 B.n1043 B.n17 10.6151
R1655 B.n1043 B.n1042 10.6151
R1656 B.n1042 B.n1041 10.6151
R1657 B.n1041 B.n25 10.6151
R1658 B.n1035 B.n25 10.6151
R1659 B.n1035 B.n1034 10.6151
R1660 B.n1034 B.n1033 10.6151
R1661 B.n1033 B.n32 10.6151
R1662 B.n1027 B.n32 10.6151
R1663 B.n1027 B.n1026 10.6151
R1664 B.n1026 B.n1025 10.6151
R1665 B.n1025 B.n39 10.6151
R1666 B.n1019 B.n39 10.6151
R1667 B.n1019 B.n1018 10.6151
R1668 B.n1018 B.n1017 10.6151
R1669 B.n1017 B.n46 10.6151
R1670 B.n1011 B.n46 10.6151
R1671 B.n1011 B.n1010 10.6151
R1672 B.n1010 B.n1009 10.6151
R1673 B.n1009 B.n52 10.6151
R1674 B.n1003 B.n52 10.6151
R1675 B.n1003 B.n1002 10.6151
R1676 B.n1002 B.n1001 10.6151
R1677 B.n1001 B.n60 10.6151
R1678 B.n995 B.n60 10.6151
R1679 B.n995 B.n994 10.6151
R1680 B.n994 B.n993 10.6151
R1681 B.n993 B.n67 10.6151
R1682 B.n987 B.n67 10.6151
R1683 B.n987 B.n986 10.6151
R1684 B.n986 B.n985 10.6151
R1685 B.n985 B.n74 10.6151
R1686 B.n979 B.n74 10.6151
R1687 B.n979 B.n978 10.6151
R1688 B.n978 B.n977 10.6151
R1689 B.n977 B.n81 10.6151
R1690 B.n971 B.n81 10.6151
R1691 B.n971 B.n970 10.6151
R1692 B.n970 B.n969 10.6151
R1693 B.n153 B.n88 10.6151
R1694 B.n156 B.n153 10.6151
R1695 B.n157 B.n156 10.6151
R1696 B.n160 B.n157 10.6151
R1697 B.n161 B.n160 10.6151
R1698 B.n164 B.n161 10.6151
R1699 B.n165 B.n164 10.6151
R1700 B.n168 B.n165 10.6151
R1701 B.n169 B.n168 10.6151
R1702 B.n172 B.n169 10.6151
R1703 B.n173 B.n172 10.6151
R1704 B.n176 B.n173 10.6151
R1705 B.n177 B.n176 10.6151
R1706 B.n180 B.n177 10.6151
R1707 B.n181 B.n180 10.6151
R1708 B.n184 B.n181 10.6151
R1709 B.n185 B.n184 10.6151
R1710 B.n188 B.n185 10.6151
R1711 B.n189 B.n188 10.6151
R1712 B.n192 B.n189 10.6151
R1713 B.n193 B.n192 10.6151
R1714 B.n196 B.n193 10.6151
R1715 B.n197 B.n196 10.6151
R1716 B.n200 B.n197 10.6151
R1717 B.n201 B.n200 10.6151
R1718 B.n204 B.n201 10.6151
R1719 B.n205 B.n204 10.6151
R1720 B.n208 B.n205 10.6151
R1721 B.n209 B.n208 10.6151
R1722 B.n212 B.n209 10.6151
R1723 B.n213 B.n212 10.6151
R1724 B.n216 B.n213 10.6151
R1725 B.n217 B.n216 10.6151
R1726 B.n220 B.n217 10.6151
R1727 B.n221 B.n220 10.6151
R1728 B.n224 B.n221 10.6151
R1729 B.n225 B.n224 10.6151
R1730 B.n228 B.n225 10.6151
R1731 B.n229 B.n228 10.6151
R1732 B.n232 B.n229 10.6151
R1733 B.n233 B.n232 10.6151
R1734 B.n236 B.n233 10.6151
R1735 B.n237 B.n236 10.6151
R1736 B.n240 B.n237 10.6151
R1737 B.n241 B.n240 10.6151
R1738 B.n244 B.n241 10.6151
R1739 B.n245 B.n244 10.6151
R1740 B.n248 B.n245 10.6151
R1741 B.n249 B.n248 10.6151
R1742 B.n252 B.n249 10.6151
R1743 B.n253 B.n252 10.6151
R1744 B.n257 B.n256 10.6151
R1745 B.n260 B.n257 10.6151
R1746 B.n261 B.n260 10.6151
R1747 B.n264 B.n261 10.6151
R1748 B.n265 B.n264 10.6151
R1749 B.n268 B.n265 10.6151
R1750 B.n269 B.n268 10.6151
R1751 B.n272 B.n269 10.6151
R1752 B.n277 B.n274 10.6151
R1753 B.n278 B.n277 10.6151
R1754 B.n281 B.n278 10.6151
R1755 B.n282 B.n281 10.6151
R1756 B.n285 B.n282 10.6151
R1757 B.n286 B.n285 10.6151
R1758 B.n289 B.n286 10.6151
R1759 B.n290 B.n289 10.6151
R1760 B.n293 B.n290 10.6151
R1761 B.n294 B.n293 10.6151
R1762 B.n297 B.n294 10.6151
R1763 B.n298 B.n297 10.6151
R1764 B.n301 B.n298 10.6151
R1765 B.n302 B.n301 10.6151
R1766 B.n305 B.n302 10.6151
R1767 B.n306 B.n305 10.6151
R1768 B.n309 B.n306 10.6151
R1769 B.n310 B.n309 10.6151
R1770 B.n313 B.n310 10.6151
R1771 B.n314 B.n313 10.6151
R1772 B.n317 B.n314 10.6151
R1773 B.n318 B.n317 10.6151
R1774 B.n321 B.n318 10.6151
R1775 B.n322 B.n321 10.6151
R1776 B.n325 B.n322 10.6151
R1777 B.n326 B.n325 10.6151
R1778 B.n329 B.n326 10.6151
R1779 B.n330 B.n329 10.6151
R1780 B.n333 B.n330 10.6151
R1781 B.n334 B.n333 10.6151
R1782 B.n337 B.n334 10.6151
R1783 B.n338 B.n337 10.6151
R1784 B.n341 B.n338 10.6151
R1785 B.n342 B.n341 10.6151
R1786 B.n345 B.n342 10.6151
R1787 B.n346 B.n345 10.6151
R1788 B.n349 B.n346 10.6151
R1789 B.n350 B.n349 10.6151
R1790 B.n353 B.n350 10.6151
R1791 B.n354 B.n353 10.6151
R1792 B.n357 B.n354 10.6151
R1793 B.n358 B.n357 10.6151
R1794 B.n361 B.n358 10.6151
R1795 B.n362 B.n361 10.6151
R1796 B.n365 B.n362 10.6151
R1797 B.n366 B.n365 10.6151
R1798 B.n369 B.n366 10.6151
R1799 B.n370 B.n369 10.6151
R1800 B.n373 B.n370 10.6151
R1801 B.n374 B.n373 10.6151
R1802 B.n964 B.n374 10.6151
R1803 B.n823 B.t0 9.05838
R1804 B.n1013 B.t5 9.05838
R1805 B.n1067 B.n0 8.11757
R1806 B.n1067 B.n1 8.11757
R1807 B.n853 B.t2 6.92712
R1808 B.n1031 B.t4 6.92712
R1809 B.n632 B.n631 6.5566
R1810 B.n649 B.n648 6.5566
R1811 B.n256 B.n152 6.5566
R1812 B.n273 B.n272 6.5566
R1813 B.n884 B.t3 4.79585
R1814 B.n1053 B.t1 4.79585
R1815 B.n631 B.n630 4.05904
R1816 B.n650 B.n649 4.05904
R1817 B.n253 B.n152 4.05904
R1818 B.n274 B.n273 4.05904
R1819 VP.n13 VP.n10 161.3
R1820 VP.n15 VP.n14 161.3
R1821 VP.n16 VP.n9 161.3
R1822 VP.n18 VP.n17 161.3
R1823 VP.n19 VP.n8 161.3
R1824 VP.n21 VP.n20 161.3
R1825 VP.n44 VP.n43 161.3
R1826 VP.n42 VP.n1 161.3
R1827 VP.n41 VP.n40 161.3
R1828 VP.n39 VP.n2 161.3
R1829 VP.n38 VP.n37 161.3
R1830 VP.n36 VP.n3 161.3
R1831 VP.n35 VP.n34 161.3
R1832 VP.n33 VP.n4 161.3
R1833 VP.n32 VP.n31 161.3
R1834 VP.n30 VP.n5 161.3
R1835 VP.n29 VP.n28 161.3
R1836 VP.n27 VP.n6 161.3
R1837 VP.n26 VP.n25 161.3
R1838 VP.n11 VP.t3 153.286
R1839 VP.n35 VP.t5 119.876
R1840 VP.n24 VP.t0 119.876
R1841 VP.n0 VP.t1 119.876
R1842 VP.n12 VP.t4 119.876
R1843 VP.n7 VP.t2 119.876
R1844 VP.n24 VP.n23 69.5151
R1845 VP.n45 VP.n0 69.5151
R1846 VP.n22 VP.n7 69.5151
R1847 VP.n30 VP.n29 56.5193
R1848 VP.n41 VP.n2 56.5193
R1849 VP.n18 VP.n9 56.5193
R1850 VP.n23 VP.n22 53.3024
R1851 VP.n12 VP.n11 49.4257
R1852 VP.n25 VP.n6 24.4675
R1853 VP.n29 VP.n6 24.4675
R1854 VP.n31 VP.n30 24.4675
R1855 VP.n31 VP.n4 24.4675
R1856 VP.n35 VP.n4 24.4675
R1857 VP.n36 VP.n35 24.4675
R1858 VP.n37 VP.n36 24.4675
R1859 VP.n37 VP.n2 24.4675
R1860 VP.n42 VP.n41 24.4675
R1861 VP.n43 VP.n42 24.4675
R1862 VP.n19 VP.n18 24.4675
R1863 VP.n20 VP.n19 24.4675
R1864 VP.n13 VP.n12 24.4675
R1865 VP.n14 VP.n13 24.4675
R1866 VP.n14 VP.n9 24.4675
R1867 VP.n25 VP.n24 20.5528
R1868 VP.n43 VP.n0 20.5528
R1869 VP.n20 VP.n7 20.5528
R1870 VP.n11 VP.n10 3.88809
R1871 VP.n22 VP.n21 0.354971
R1872 VP.n26 VP.n23 0.354971
R1873 VP.n45 VP.n44 0.354971
R1874 VP VP.n45 0.26696
R1875 VP.n15 VP.n10 0.189894
R1876 VP.n16 VP.n15 0.189894
R1877 VP.n17 VP.n16 0.189894
R1878 VP.n17 VP.n8 0.189894
R1879 VP.n21 VP.n8 0.189894
R1880 VP.n27 VP.n26 0.189894
R1881 VP.n28 VP.n27 0.189894
R1882 VP.n28 VP.n5 0.189894
R1883 VP.n32 VP.n5 0.189894
R1884 VP.n33 VP.n32 0.189894
R1885 VP.n34 VP.n33 0.189894
R1886 VP.n34 VP.n3 0.189894
R1887 VP.n38 VP.n3 0.189894
R1888 VP.n39 VP.n38 0.189894
R1889 VP.n40 VP.n39 0.189894
R1890 VP.n40 VP.n1 0.189894
R1891 VP.n44 VP.n1 0.189894
R1892 VTAIL.n346 VTAIL.n266 289.615
R1893 VTAIL.n82 VTAIL.n2 289.615
R1894 VTAIL.n260 VTAIL.n180 289.615
R1895 VTAIL.n172 VTAIL.n92 289.615
R1896 VTAIL.n295 VTAIL.n294 185
R1897 VTAIL.n297 VTAIL.n296 185
R1898 VTAIL.n290 VTAIL.n289 185
R1899 VTAIL.n303 VTAIL.n302 185
R1900 VTAIL.n305 VTAIL.n304 185
R1901 VTAIL.n286 VTAIL.n285 185
R1902 VTAIL.n311 VTAIL.n310 185
R1903 VTAIL.n313 VTAIL.n312 185
R1904 VTAIL.n282 VTAIL.n281 185
R1905 VTAIL.n319 VTAIL.n318 185
R1906 VTAIL.n321 VTAIL.n320 185
R1907 VTAIL.n278 VTAIL.n277 185
R1908 VTAIL.n327 VTAIL.n326 185
R1909 VTAIL.n329 VTAIL.n328 185
R1910 VTAIL.n274 VTAIL.n273 185
R1911 VTAIL.n336 VTAIL.n335 185
R1912 VTAIL.n337 VTAIL.n272 185
R1913 VTAIL.n339 VTAIL.n338 185
R1914 VTAIL.n270 VTAIL.n269 185
R1915 VTAIL.n345 VTAIL.n344 185
R1916 VTAIL.n347 VTAIL.n346 185
R1917 VTAIL.n31 VTAIL.n30 185
R1918 VTAIL.n33 VTAIL.n32 185
R1919 VTAIL.n26 VTAIL.n25 185
R1920 VTAIL.n39 VTAIL.n38 185
R1921 VTAIL.n41 VTAIL.n40 185
R1922 VTAIL.n22 VTAIL.n21 185
R1923 VTAIL.n47 VTAIL.n46 185
R1924 VTAIL.n49 VTAIL.n48 185
R1925 VTAIL.n18 VTAIL.n17 185
R1926 VTAIL.n55 VTAIL.n54 185
R1927 VTAIL.n57 VTAIL.n56 185
R1928 VTAIL.n14 VTAIL.n13 185
R1929 VTAIL.n63 VTAIL.n62 185
R1930 VTAIL.n65 VTAIL.n64 185
R1931 VTAIL.n10 VTAIL.n9 185
R1932 VTAIL.n72 VTAIL.n71 185
R1933 VTAIL.n73 VTAIL.n8 185
R1934 VTAIL.n75 VTAIL.n74 185
R1935 VTAIL.n6 VTAIL.n5 185
R1936 VTAIL.n81 VTAIL.n80 185
R1937 VTAIL.n83 VTAIL.n82 185
R1938 VTAIL.n261 VTAIL.n260 185
R1939 VTAIL.n259 VTAIL.n258 185
R1940 VTAIL.n184 VTAIL.n183 185
R1941 VTAIL.n188 VTAIL.n186 185
R1942 VTAIL.n253 VTAIL.n252 185
R1943 VTAIL.n251 VTAIL.n250 185
R1944 VTAIL.n190 VTAIL.n189 185
R1945 VTAIL.n245 VTAIL.n244 185
R1946 VTAIL.n243 VTAIL.n242 185
R1947 VTAIL.n194 VTAIL.n193 185
R1948 VTAIL.n237 VTAIL.n236 185
R1949 VTAIL.n235 VTAIL.n234 185
R1950 VTAIL.n198 VTAIL.n197 185
R1951 VTAIL.n229 VTAIL.n228 185
R1952 VTAIL.n227 VTAIL.n226 185
R1953 VTAIL.n202 VTAIL.n201 185
R1954 VTAIL.n221 VTAIL.n220 185
R1955 VTAIL.n219 VTAIL.n218 185
R1956 VTAIL.n206 VTAIL.n205 185
R1957 VTAIL.n213 VTAIL.n212 185
R1958 VTAIL.n211 VTAIL.n210 185
R1959 VTAIL.n173 VTAIL.n172 185
R1960 VTAIL.n171 VTAIL.n170 185
R1961 VTAIL.n96 VTAIL.n95 185
R1962 VTAIL.n100 VTAIL.n98 185
R1963 VTAIL.n165 VTAIL.n164 185
R1964 VTAIL.n163 VTAIL.n162 185
R1965 VTAIL.n102 VTAIL.n101 185
R1966 VTAIL.n157 VTAIL.n156 185
R1967 VTAIL.n155 VTAIL.n154 185
R1968 VTAIL.n106 VTAIL.n105 185
R1969 VTAIL.n149 VTAIL.n148 185
R1970 VTAIL.n147 VTAIL.n146 185
R1971 VTAIL.n110 VTAIL.n109 185
R1972 VTAIL.n141 VTAIL.n140 185
R1973 VTAIL.n139 VTAIL.n138 185
R1974 VTAIL.n114 VTAIL.n113 185
R1975 VTAIL.n133 VTAIL.n132 185
R1976 VTAIL.n131 VTAIL.n130 185
R1977 VTAIL.n118 VTAIL.n117 185
R1978 VTAIL.n125 VTAIL.n124 185
R1979 VTAIL.n123 VTAIL.n122 185
R1980 VTAIL.n293 VTAIL.t3 147.659
R1981 VTAIL.n29 VTAIL.t4 147.659
R1982 VTAIL.n209 VTAIL.t8 147.659
R1983 VTAIL.n121 VTAIL.t2 147.659
R1984 VTAIL.n296 VTAIL.n295 104.615
R1985 VTAIL.n296 VTAIL.n289 104.615
R1986 VTAIL.n303 VTAIL.n289 104.615
R1987 VTAIL.n304 VTAIL.n303 104.615
R1988 VTAIL.n304 VTAIL.n285 104.615
R1989 VTAIL.n311 VTAIL.n285 104.615
R1990 VTAIL.n312 VTAIL.n311 104.615
R1991 VTAIL.n312 VTAIL.n281 104.615
R1992 VTAIL.n319 VTAIL.n281 104.615
R1993 VTAIL.n320 VTAIL.n319 104.615
R1994 VTAIL.n320 VTAIL.n277 104.615
R1995 VTAIL.n327 VTAIL.n277 104.615
R1996 VTAIL.n328 VTAIL.n327 104.615
R1997 VTAIL.n328 VTAIL.n273 104.615
R1998 VTAIL.n336 VTAIL.n273 104.615
R1999 VTAIL.n337 VTAIL.n336 104.615
R2000 VTAIL.n338 VTAIL.n337 104.615
R2001 VTAIL.n338 VTAIL.n269 104.615
R2002 VTAIL.n345 VTAIL.n269 104.615
R2003 VTAIL.n346 VTAIL.n345 104.615
R2004 VTAIL.n32 VTAIL.n31 104.615
R2005 VTAIL.n32 VTAIL.n25 104.615
R2006 VTAIL.n39 VTAIL.n25 104.615
R2007 VTAIL.n40 VTAIL.n39 104.615
R2008 VTAIL.n40 VTAIL.n21 104.615
R2009 VTAIL.n47 VTAIL.n21 104.615
R2010 VTAIL.n48 VTAIL.n47 104.615
R2011 VTAIL.n48 VTAIL.n17 104.615
R2012 VTAIL.n55 VTAIL.n17 104.615
R2013 VTAIL.n56 VTAIL.n55 104.615
R2014 VTAIL.n56 VTAIL.n13 104.615
R2015 VTAIL.n63 VTAIL.n13 104.615
R2016 VTAIL.n64 VTAIL.n63 104.615
R2017 VTAIL.n64 VTAIL.n9 104.615
R2018 VTAIL.n72 VTAIL.n9 104.615
R2019 VTAIL.n73 VTAIL.n72 104.615
R2020 VTAIL.n74 VTAIL.n73 104.615
R2021 VTAIL.n74 VTAIL.n5 104.615
R2022 VTAIL.n81 VTAIL.n5 104.615
R2023 VTAIL.n82 VTAIL.n81 104.615
R2024 VTAIL.n260 VTAIL.n259 104.615
R2025 VTAIL.n259 VTAIL.n183 104.615
R2026 VTAIL.n188 VTAIL.n183 104.615
R2027 VTAIL.n252 VTAIL.n188 104.615
R2028 VTAIL.n252 VTAIL.n251 104.615
R2029 VTAIL.n251 VTAIL.n189 104.615
R2030 VTAIL.n244 VTAIL.n189 104.615
R2031 VTAIL.n244 VTAIL.n243 104.615
R2032 VTAIL.n243 VTAIL.n193 104.615
R2033 VTAIL.n236 VTAIL.n193 104.615
R2034 VTAIL.n236 VTAIL.n235 104.615
R2035 VTAIL.n235 VTAIL.n197 104.615
R2036 VTAIL.n228 VTAIL.n197 104.615
R2037 VTAIL.n228 VTAIL.n227 104.615
R2038 VTAIL.n227 VTAIL.n201 104.615
R2039 VTAIL.n220 VTAIL.n201 104.615
R2040 VTAIL.n220 VTAIL.n219 104.615
R2041 VTAIL.n219 VTAIL.n205 104.615
R2042 VTAIL.n212 VTAIL.n205 104.615
R2043 VTAIL.n212 VTAIL.n211 104.615
R2044 VTAIL.n172 VTAIL.n171 104.615
R2045 VTAIL.n171 VTAIL.n95 104.615
R2046 VTAIL.n100 VTAIL.n95 104.615
R2047 VTAIL.n164 VTAIL.n100 104.615
R2048 VTAIL.n164 VTAIL.n163 104.615
R2049 VTAIL.n163 VTAIL.n101 104.615
R2050 VTAIL.n156 VTAIL.n101 104.615
R2051 VTAIL.n156 VTAIL.n155 104.615
R2052 VTAIL.n155 VTAIL.n105 104.615
R2053 VTAIL.n148 VTAIL.n105 104.615
R2054 VTAIL.n148 VTAIL.n147 104.615
R2055 VTAIL.n147 VTAIL.n109 104.615
R2056 VTAIL.n140 VTAIL.n109 104.615
R2057 VTAIL.n140 VTAIL.n139 104.615
R2058 VTAIL.n139 VTAIL.n113 104.615
R2059 VTAIL.n132 VTAIL.n113 104.615
R2060 VTAIL.n132 VTAIL.n131 104.615
R2061 VTAIL.n131 VTAIL.n117 104.615
R2062 VTAIL.n124 VTAIL.n117 104.615
R2063 VTAIL.n124 VTAIL.n123 104.615
R2064 VTAIL.n295 VTAIL.t3 52.3082
R2065 VTAIL.n31 VTAIL.t4 52.3082
R2066 VTAIL.n211 VTAIL.t8 52.3082
R2067 VTAIL.n123 VTAIL.t2 52.3082
R2068 VTAIL.n179 VTAIL.n178 44.3577
R2069 VTAIL.n91 VTAIL.n90 44.3577
R2070 VTAIL.n1 VTAIL.n0 44.3575
R2071 VTAIL.n89 VTAIL.n88 44.3575
R2072 VTAIL.n351 VTAIL.n350 32.3793
R2073 VTAIL.n87 VTAIL.n86 32.3793
R2074 VTAIL.n265 VTAIL.n264 32.3793
R2075 VTAIL.n177 VTAIL.n176 32.3793
R2076 VTAIL.n91 VTAIL.n89 31.5134
R2077 VTAIL.n351 VTAIL.n265 28.5652
R2078 VTAIL.n294 VTAIL.n293 15.6677
R2079 VTAIL.n30 VTAIL.n29 15.6677
R2080 VTAIL.n210 VTAIL.n209 15.6677
R2081 VTAIL.n122 VTAIL.n121 15.6677
R2082 VTAIL.n339 VTAIL.n270 13.1884
R2083 VTAIL.n75 VTAIL.n6 13.1884
R2084 VTAIL.n186 VTAIL.n184 13.1884
R2085 VTAIL.n98 VTAIL.n96 13.1884
R2086 VTAIL.n297 VTAIL.n292 12.8005
R2087 VTAIL.n340 VTAIL.n272 12.8005
R2088 VTAIL.n344 VTAIL.n343 12.8005
R2089 VTAIL.n33 VTAIL.n28 12.8005
R2090 VTAIL.n76 VTAIL.n8 12.8005
R2091 VTAIL.n80 VTAIL.n79 12.8005
R2092 VTAIL.n258 VTAIL.n257 12.8005
R2093 VTAIL.n254 VTAIL.n253 12.8005
R2094 VTAIL.n213 VTAIL.n208 12.8005
R2095 VTAIL.n170 VTAIL.n169 12.8005
R2096 VTAIL.n166 VTAIL.n165 12.8005
R2097 VTAIL.n125 VTAIL.n120 12.8005
R2098 VTAIL.n298 VTAIL.n290 12.0247
R2099 VTAIL.n335 VTAIL.n334 12.0247
R2100 VTAIL.n347 VTAIL.n268 12.0247
R2101 VTAIL.n34 VTAIL.n26 12.0247
R2102 VTAIL.n71 VTAIL.n70 12.0247
R2103 VTAIL.n83 VTAIL.n4 12.0247
R2104 VTAIL.n261 VTAIL.n182 12.0247
R2105 VTAIL.n250 VTAIL.n187 12.0247
R2106 VTAIL.n214 VTAIL.n206 12.0247
R2107 VTAIL.n173 VTAIL.n94 12.0247
R2108 VTAIL.n162 VTAIL.n99 12.0247
R2109 VTAIL.n126 VTAIL.n118 12.0247
R2110 VTAIL.n302 VTAIL.n301 11.249
R2111 VTAIL.n333 VTAIL.n274 11.249
R2112 VTAIL.n348 VTAIL.n266 11.249
R2113 VTAIL.n38 VTAIL.n37 11.249
R2114 VTAIL.n69 VTAIL.n10 11.249
R2115 VTAIL.n84 VTAIL.n2 11.249
R2116 VTAIL.n262 VTAIL.n180 11.249
R2117 VTAIL.n249 VTAIL.n190 11.249
R2118 VTAIL.n218 VTAIL.n217 11.249
R2119 VTAIL.n174 VTAIL.n92 11.249
R2120 VTAIL.n161 VTAIL.n102 11.249
R2121 VTAIL.n130 VTAIL.n129 11.249
R2122 VTAIL.n305 VTAIL.n288 10.4732
R2123 VTAIL.n330 VTAIL.n329 10.4732
R2124 VTAIL.n41 VTAIL.n24 10.4732
R2125 VTAIL.n66 VTAIL.n65 10.4732
R2126 VTAIL.n246 VTAIL.n245 10.4732
R2127 VTAIL.n221 VTAIL.n204 10.4732
R2128 VTAIL.n158 VTAIL.n157 10.4732
R2129 VTAIL.n133 VTAIL.n116 10.4732
R2130 VTAIL.n306 VTAIL.n286 9.69747
R2131 VTAIL.n326 VTAIL.n276 9.69747
R2132 VTAIL.n42 VTAIL.n22 9.69747
R2133 VTAIL.n62 VTAIL.n12 9.69747
R2134 VTAIL.n242 VTAIL.n192 9.69747
R2135 VTAIL.n222 VTAIL.n202 9.69747
R2136 VTAIL.n154 VTAIL.n104 9.69747
R2137 VTAIL.n134 VTAIL.n114 9.69747
R2138 VTAIL.n350 VTAIL.n349 9.45567
R2139 VTAIL.n86 VTAIL.n85 9.45567
R2140 VTAIL.n264 VTAIL.n263 9.45567
R2141 VTAIL.n176 VTAIL.n175 9.45567
R2142 VTAIL.n349 VTAIL.n348 9.3005
R2143 VTAIL.n268 VTAIL.n267 9.3005
R2144 VTAIL.n343 VTAIL.n342 9.3005
R2145 VTAIL.n315 VTAIL.n314 9.3005
R2146 VTAIL.n284 VTAIL.n283 9.3005
R2147 VTAIL.n309 VTAIL.n308 9.3005
R2148 VTAIL.n307 VTAIL.n306 9.3005
R2149 VTAIL.n288 VTAIL.n287 9.3005
R2150 VTAIL.n301 VTAIL.n300 9.3005
R2151 VTAIL.n299 VTAIL.n298 9.3005
R2152 VTAIL.n292 VTAIL.n291 9.3005
R2153 VTAIL.n317 VTAIL.n316 9.3005
R2154 VTAIL.n280 VTAIL.n279 9.3005
R2155 VTAIL.n323 VTAIL.n322 9.3005
R2156 VTAIL.n325 VTAIL.n324 9.3005
R2157 VTAIL.n276 VTAIL.n275 9.3005
R2158 VTAIL.n331 VTAIL.n330 9.3005
R2159 VTAIL.n333 VTAIL.n332 9.3005
R2160 VTAIL.n334 VTAIL.n271 9.3005
R2161 VTAIL.n341 VTAIL.n340 9.3005
R2162 VTAIL.n85 VTAIL.n84 9.3005
R2163 VTAIL.n4 VTAIL.n3 9.3005
R2164 VTAIL.n79 VTAIL.n78 9.3005
R2165 VTAIL.n51 VTAIL.n50 9.3005
R2166 VTAIL.n20 VTAIL.n19 9.3005
R2167 VTAIL.n45 VTAIL.n44 9.3005
R2168 VTAIL.n43 VTAIL.n42 9.3005
R2169 VTAIL.n24 VTAIL.n23 9.3005
R2170 VTAIL.n37 VTAIL.n36 9.3005
R2171 VTAIL.n35 VTAIL.n34 9.3005
R2172 VTAIL.n28 VTAIL.n27 9.3005
R2173 VTAIL.n53 VTAIL.n52 9.3005
R2174 VTAIL.n16 VTAIL.n15 9.3005
R2175 VTAIL.n59 VTAIL.n58 9.3005
R2176 VTAIL.n61 VTAIL.n60 9.3005
R2177 VTAIL.n12 VTAIL.n11 9.3005
R2178 VTAIL.n67 VTAIL.n66 9.3005
R2179 VTAIL.n69 VTAIL.n68 9.3005
R2180 VTAIL.n70 VTAIL.n7 9.3005
R2181 VTAIL.n77 VTAIL.n76 9.3005
R2182 VTAIL.n196 VTAIL.n195 9.3005
R2183 VTAIL.n239 VTAIL.n238 9.3005
R2184 VTAIL.n241 VTAIL.n240 9.3005
R2185 VTAIL.n192 VTAIL.n191 9.3005
R2186 VTAIL.n247 VTAIL.n246 9.3005
R2187 VTAIL.n249 VTAIL.n248 9.3005
R2188 VTAIL.n187 VTAIL.n185 9.3005
R2189 VTAIL.n255 VTAIL.n254 9.3005
R2190 VTAIL.n263 VTAIL.n262 9.3005
R2191 VTAIL.n182 VTAIL.n181 9.3005
R2192 VTAIL.n257 VTAIL.n256 9.3005
R2193 VTAIL.n233 VTAIL.n232 9.3005
R2194 VTAIL.n231 VTAIL.n230 9.3005
R2195 VTAIL.n200 VTAIL.n199 9.3005
R2196 VTAIL.n225 VTAIL.n224 9.3005
R2197 VTAIL.n223 VTAIL.n222 9.3005
R2198 VTAIL.n204 VTAIL.n203 9.3005
R2199 VTAIL.n217 VTAIL.n216 9.3005
R2200 VTAIL.n215 VTAIL.n214 9.3005
R2201 VTAIL.n208 VTAIL.n207 9.3005
R2202 VTAIL.n108 VTAIL.n107 9.3005
R2203 VTAIL.n151 VTAIL.n150 9.3005
R2204 VTAIL.n153 VTAIL.n152 9.3005
R2205 VTAIL.n104 VTAIL.n103 9.3005
R2206 VTAIL.n159 VTAIL.n158 9.3005
R2207 VTAIL.n161 VTAIL.n160 9.3005
R2208 VTAIL.n99 VTAIL.n97 9.3005
R2209 VTAIL.n167 VTAIL.n166 9.3005
R2210 VTAIL.n175 VTAIL.n174 9.3005
R2211 VTAIL.n94 VTAIL.n93 9.3005
R2212 VTAIL.n169 VTAIL.n168 9.3005
R2213 VTAIL.n145 VTAIL.n144 9.3005
R2214 VTAIL.n143 VTAIL.n142 9.3005
R2215 VTAIL.n112 VTAIL.n111 9.3005
R2216 VTAIL.n137 VTAIL.n136 9.3005
R2217 VTAIL.n135 VTAIL.n134 9.3005
R2218 VTAIL.n116 VTAIL.n115 9.3005
R2219 VTAIL.n129 VTAIL.n128 9.3005
R2220 VTAIL.n127 VTAIL.n126 9.3005
R2221 VTAIL.n120 VTAIL.n119 9.3005
R2222 VTAIL.n310 VTAIL.n309 8.92171
R2223 VTAIL.n325 VTAIL.n278 8.92171
R2224 VTAIL.n46 VTAIL.n45 8.92171
R2225 VTAIL.n61 VTAIL.n14 8.92171
R2226 VTAIL.n241 VTAIL.n194 8.92171
R2227 VTAIL.n226 VTAIL.n225 8.92171
R2228 VTAIL.n153 VTAIL.n106 8.92171
R2229 VTAIL.n138 VTAIL.n137 8.92171
R2230 VTAIL.n313 VTAIL.n284 8.14595
R2231 VTAIL.n322 VTAIL.n321 8.14595
R2232 VTAIL.n49 VTAIL.n20 8.14595
R2233 VTAIL.n58 VTAIL.n57 8.14595
R2234 VTAIL.n238 VTAIL.n237 8.14595
R2235 VTAIL.n229 VTAIL.n200 8.14595
R2236 VTAIL.n150 VTAIL.n149 8.14595
R2237 VTAIL.n141 VTAIL.n112 8.14595
R2238 VTAIL.n314 VTAIL.n282 7.3702
R2239 VTAIL.n318 VTAIL.n280 7.3702
R2240 VTAIL.n50 VTAIL.n18 7.3702
R2241 VTAIL.n54 VTAIL.n16 7.3702
R2242 VTAIL.n234 VTAIL.n196 7.3702
R2243 VTAIL.n230 VTAIL.n198 7.3702
R2244 VTAIL.n146 VTAIL.n108 7.3702
R2245 VTAIL.n142 VTAIL.n110 7.3702
R2246 VTAIL.n317 VTAIL.n282 6.59444
R2247 VTAIL.n318 VTAIL.n317 6.59444
R2248 VTAIL.n53 VTAIL.n18 6.59444
R2249 VTAIL.n54 VTAIL.n53 6.59444
R2250 VTAIL.n234 VTAIL.n233 6.59444
R2251 VTAIL.n233 VTAIL.n198 6.59444
R2252 VTAIL.n146 VTAIL.n145 6.59444
R2253 VTAIL.n145 VTAIL.n110 6.59444
R2254 VTAIL.n314 VTAIL.n313 5.81868
R2255 VTAIL.n321 VTAIL.n280 5.81868
R2256 VTAIL.n50 VTAIL.n49 5.81868
R2257 VTAIL.n57 VTAIL.n16 5.81868
R2258 VTAIL.n237 VTAIL.n196 5.81868
R2259 VTAIL.n230 VTAIL.n229 5.81868
R2260 VTAIL.n149 VTAIL.n108 5.81868
R2261 VTAIL.n142 VTAIL.n141 5.81868
R2262 VTAIL.n310 VTAIL.n284 5.04292
R2263 VTAIL.n322 VTAIL.n278 5.04292
R2264 VTAIL.n46 VTAIL.n20 5.04292
R2265 VTAIL.n58 VTAIL.n14 5.04292
R2266 VTAIL.n238 VTAIL.n194 5.04292
R2267 VTAIL.n226 VTAIL.n200 5.04292
R2268 VTAIL.n150 VTAIL.n106 5.04292
R2269 VTAIL.n138 VTAIL.n112 5.04292
R2270 VTAIL.n293 VTAIL.n291 4.38563
R2271 VTAIL.n29 VTAIL.n27 4.38563
R2272 VTAIL.n209 VTAIL.n207 4.38563
R2273 VTAIL.n121 VTAIL.n119 4.38563
R2274 VTAIL.n309 VTAIL.n286 4.26717
R2275 VTAIL.n326 VTAIL.n325 4.26717
R2276 VTAIL.n45 VTAIL.n22 4.26717
R2277 VTAIL.n62 VTAIL.n61 4.26717
R2278 VTAIL.n242 VTAIL.n241 4.26717
R2279 VTAIL.n225 VTAIL.n202 4.26717
R2280 VTAIL.n154 VTAIL.n153 4.26717
R2281 VTAIL.n137 VTAIL.n114 4.26717
R2282 VTAIL.n306 VTAIL.n305 3.49141
R2283 VTAIL.n329 VTAIL.n276 3.49141
R2284 VTAIL.n42 VTAIL.n41 3.49141
R2285 VTAIL.n65 VTAIL.n12 3.49141
R2286 VTAIL.n245 VTAIL.n192 3.49141
R2287 VTAIL.n222 VTAIL.n221 3.49141
R2288 VTAIL.n157 VTAIL.n104 3.49141
R2289 VTAIL.n134 VTAIL.n133 3.49141
R2290 VTAIL.n177 VTAIL.n91 2.94878
R2291 VTAIL.n265 VTAIL.n179 2.94878
R2292 VTAIL.n89 VTAIL.n87 2.94878
R2293 VTAIL.n302 VTAIL.n288 2.71565
R2294 VTAIL.n330 VTAIL.n274 2.71565
R2295 VTAIL.n350 VTAIL.n266 2.71565
R2296 VTAIL.n38 VTAIL.n24 2.71565
R2297 VTAIL.n66 VTAIL.n10 2.71565
R2298 VTAIL.n86 VTAIL.n2 2.71565
R2299 VTAIL.n264 VTAIL.n180 2.71565
R2300 VTAIL.n246 VTAIL.n190 2.71565
R2301 VTAIL.n218 VTAIL.n204 2.71565
R2302 VTAIL.n176 VTAIL.n92 2.71565
R2303 VTAIL.n158 VTAIL.n102 2.71565
R2304 VTAIL.n130 VTAIL.n116 2.71565
R2305 VTAIL VTAIL.n351 2.15352
R2306 VTAIL.n179 VTAIL.n177 1.94447
R2307 VTAIL.n87 VTAIL.n1 1.94447
R2308 VTAIL.n301 VTAIL.n290 1.93989
R2309 VTAIL.n335 VTAIL.n333 1.93989
R2310 VTAIL.n348 VTAIL.n347 1.93989
R2311 VTAIL.n37 VTAIL.n26 1.93989
R2312 VTAIL.n71 VTAIL.n69 1.93989
R2313 VTAIL.n84 VTAIL.n83 1.93989
R2314 VTAIL.n262 VTAIL.n261 1.93989
R2315 VTAIL.n250 VTAIL.n249 1.93989
R2316 VTAIL.n217 VTAIL.n206 1.93989
R2317 VTAIL.n174 VTAIL.n173 1.93989
R2318 VTAIL.n162 VTAIL.n161 1.93989
R2319 VTAIL.n129 VTAIL.n118 1.93989
R2320 VTAIL.n0 VTAIL.t1 1.28872
R2321 VTAIL.n0 VTAIL.t11 1.28872
R2322 VTAIL.n88 VTAIL.t6 1.28872
R2323 VTAIL.n88 VTAIL.t5 1.28872
R2324 VTAIL.n178 VTAIL.t9 1.28872
R2325 VTAIL.n178 VTAIL.t7 1.28872
R2326 VTAIL.n90 VTAIL.t10 1.28872
R2327 VTAIL.n90 VTAIL.t0 1.28872
R2328 VTAIL.n298 VTAIL.n297 1.16414
R2329 VTAIL.n334 VTAIL.n272 1.16414
R2330 VTAIL.n344 VTAIL.n268 1.16414
R2331 VTAIL.n34 VTAIL.n33 1.16414
R2332 VTAIL.n70 VTAIL.n8 1.16414
R2333 VTAIL.n80 VTAIL.n4 1.16414
R2334 VTAIL.n258 VTAIL.n182 1.16414
R2335 VTAIL.n253 VTAIL.n187 1.16414
R2336 VTAIL.n214 VTAIL.n213 1.16414
R2337 VTAIL.n170 VTAIL.n94 1.16414
R2338 VTAIL.n165 VTAIL.n99 1.16414
R2339 VTAIL.n126 VTAIL.n125 1.16414
R2340 VTAIL VTAIL.n1 0.795759
R2341 VTAIL.n294 VTAIL.n292 0.388379
R2342 VTAIL.n340 VTAIL.n339 0.388379
R2343 VTAIL.n343 VTAIL.n270 0.388379
R2344 VTAIL.n30 VTAIL.n28 0.388379
R2345 VTAIL.n76 VTAIL.n75 0.388379
R2346 VTAIL.n79 VTAIL.n6 0.388379
R2347 VTAIL.n257 VTAIL.n184 0.388379
R2348 VTAIL.n254 VTAIL.n186 0.388379
R2349 VTAIL.n210 VTAIL.n208 0.388379
R2350 VTAIL.n169 VTAIL.n96 0.388379
R2351 VTAIL.n166 VTAIL.n98 0.388379
R2352 VTAIL.n122 VTAIL.n120 0.388379
R2353 VTAIL.n299 VTAIL.n291 0.155672
R2354 VTAIL.n300 VTAIL.n299 0.155672
R2355 VTAIL.n300 VTAIL.n287 0.155672
R2356 VTAIL.n307 VTAIL.n287 0.155672
R2357 VTAIL.n308 VTAIL.n307 0.155672
R2358 VTAIL.n308 VTAIL.n283 0.155672
R2359 VTAIL.n315 VTAIL.n283 0.155672
R2360 VTAIL.n316 VTAIL.n315 0.155672
R2361 VTAIL.n316 VTAIL.n279 0.155672
R2362 VTAIL.n323 VTAIL.n279 0.155672
R2363 VTAIL.n324 VTAIL.n323 0.155672
R2364 VTAIL.n324 VTAIL.n275 0.155672
R2365 VTAIL.n331 VTAIL.n275 0.155672
R2366 VTAIL.n332 VTAIL.n331 0.155672
R2367 VTAIL.n332 VTAIL.n271 0.155672
R2368 VTAIL.n341 VTAIL.n271 0.155672
R2369 VTAIL.n342 VTAIL.n341 0.155672
R2370 VTAIL.n342 VTAIL.n267 0.155672
R2371 VTAIL.n349 VTAIL.n267 0.155672
R2372 VTAIL.n35 VTAIL.n27 0.155672
R2373 VTAIL.n36 VTAIL.n35 0.155672
R2374 VTAIL.n36 VTAIL.n23 0.155672
R2375 VTAIL.n43 VTAIL.n23 0.155672
R2376 VTAIL.n44 VTAIL.n43 0.155672
R2377 VTAIL.n44 VTAIL.n19 0.155672
R2378 VTAIL.n51 VTAIL.n19 0.155672
R2379 VTAIL.n52 VTAIL.n51 0.155672
R2380 VTAIL.n52 VTAIL.n15 0.155672
R2381 VTAIL.n59 VTAIL.n15 0.155672
R2382 VTAIL.n60 VTAIL.n59 0.155672
R2383 VTAIL.n60 VTAIL.n11 0.155672
R2384 VTAIL.n67 VTAIL.n11 0.155672
R2385 VTAIL.n68 VTAIL.n67 0.155672
R2386 VTAIL.n68 VTAIL.n7 0.155672
R2387 VTAIL.n77 VTAIL.n7 0.155672
R2388 VTAIL.n78 VTAIL.n77 0.155672
R2389 VTAIL.n78 VTAIL.n3 0.155672
R2390 VTAIL.n85 VTAIL.n3 0.155672
R2391 VTAIL.n263 VTAIL.n181 0.155672
R2392 VTAIL.n256 VTAIL.n181 0.155672
R2393 VTAIL.n256 VTAIL.n255 0.155672
R2394 VTAIL.n255 VTAIL.n185 0.155672
R2395 VTAIL.n248 VTAIL.n185 0.155672
R2396 VTAIL.n248 VTAIL.n247 0.155672
R2397 VTAIL.n247 VTAIL.n191 0.155672
R2398 VTAIL.n240 VTAIL.n191 0.155672
R2399 VTAIL.n240 VTAIL.n239 0.155672
R2400 VTAIL.n239 VTAIL.n195 0.155672
R2401 VTAIL.n232 VTAIL.n195 0.155672
R2402 VTAIL.n232 VTAIL.n231 0.155672
R2403 VTAIL.n231 VTAIL.n199 0.155672
R2404 VTAIL.n224 VTAIL.n199 0.155672
R2405 VTAIL.n224 VTAIL.n223 0.155672
R2406 VTAIL.n223 VTAIL.n203 0.155672
R2407 VTAIL.n216 VTAIL.n203 0.155672
R2408 VTAIL.n216 VTAIL.n215 0.155672
R2409 VTAIL.n215 VTAIL.n207 0.155672
R2410 VTAIL.n175 VTAIL.n93 0.155672
R2411 VTAIL.n168 VTAIL.n93 0.155672
R2412 VTAIL.n168 VTAIL.n167 0.155672
R2413 VTAIL.n167 VTAIL.n97 0.155672
R2414 VTAIL.n160 VTAIL.n97 0.155672
R2415 VTAIL.n160 VTAIL.n159 0.155672
R2416 VTAIL.n159 VTAIL.n103 0.155672
R2417 VTAIL.n152 VTAIL.n103 0.155672
R2418 VTAIL.n152 VTAIL.n151 0.155672
R2419 VTAIL.n151 VTAIL.n107 0.155672
R2420 VTAIL.n144 VTAIL.n107 0.155672
R2421 VTAIL.n144 VTAIL.n143 0.155672
R2422 VTAIL.n143 VTAIL.n111 0.155672
R2423 VTAIL.n136 VTAIL.n111 0.155672
R2424 VTAIL.n136 VTAIL.n135 0.155672
R2425 VTAIL.n135 VTAIL.n115 0.155672
R2426 VTAIL.n128 VTAIL.n115 0.155672
R2427 VTAIL.n128 VTAIL.n127 0.155672
R2428 VTAIL.n127 VTAIL.n119 0.155672
R2429 VDD1.n80 VDD1.n0 289.615
R2430 VDD1.n165 VDD1.n85 289.615
R2431 VDD1.n81 VDD1.n80 185
R2432 VDD1.n79 VDD1.n78 185
R2433 VDD1.n4 VDD1.n3 185
R2434 VDD1.n8 VDD1.n6 185
R2435 VDD1.n73 VDD1.n72 185
R2436 VDD1.n71 VDD1.n70 185
R2437 VDD1.n10 VDD1.n9 185
R2438 VDD1.n65 VDD1.n64 185
R2439 VDD1.n63 VDD1.n62 185
R2440 VDD1.n14 VDD1.n13 185
R2441 VDD1.n57 VDD1.n56 185
R2442 VDD1.n55 VDD1.n54 185
R2443 VDD1.n18 VDD1.n17 185
R2444 VDD1.n49 VDD1.n48 185
R2445 VDD1.n47 VDD1.n46 185
R2446 VDD1.n22 VDD1.n21 185
R2447 VDD1.n41 VDD1.n40 185
R2448 VDD1.n39 VDD1.n38 185
R2449 VDD1.n26 VDD1.n25 185
R2450 VDD1.n33 VDD1.n32 185
R2451 VDD1.n31 VDD1.n30 185
R2452 VDD1.n114 VDD1.n113 185
R2453 VDD1.n116 VDD1.n115 185
R2454 VDD1.n109 VDD1.n108 185
R2455 VDD1.n122 VDD1.n121 185
R2456 VDD1.n124 VDD1.n123 185
R2457 VDD1.n105 VDD1.n104 185
R2458 VDD1.n130 VDD1.n129 185
R2459 VDD1.n132 VDD1.n131 185
R2460 VDD1.n101 VDD1.n100 185
R2461 VDD1.n138 VDD1.n137 185
R2462 VDD1.n140 VDD1.n139 185
R2463 VDD1.n97 VDD1.n96 185
R2464 VDD1.n146 VDD1.n145 185
R2465 VDD1.n148 VDD1.n147 185
R2466 VDD1.n93 VDD1.n92 185
R2467 VDD1.n155 VDD1.n154 185
R2468 VDD1.n156 VDD1.n91 185
R2469 VDD1.n158 VDD1.n157 185
R2470 VDD1.n89 VDD1.n88 185
R2471 VDD1.n164 VDD1.n163 185
R2472 VDD1.n166 VDD1.n165 185
R2473 VDD1.n29 VDD1.t2 147.659
R2474 VDD1.n112 VDD1.t5 147.659
R2475 VDD1.n80 VDD1.n79 104.615
R2476 VDD1.n79 VDD1.n3 104.615
R2477 VDD1.n8 VDD1.n3 104.615
R2478 VDD1.n72 VDD1.n8 104.615
R2479 VDD1.n72 VDD1.n71 104.615
R2480 VDD1.n71 VDD1.n9 104.615
R2481 VDD1.n64 VDD1.n9 104.615
R2482 VDD1.n64 VDD1.n63 104.615
R2483 VDD1.n63 VDD1.n13 104.615
R2484 VDD1.n56 VDD1.n13 104.615
R2485 VDD1.n56 VDD1.n55 104.615
R2486 VDD1.n55 VDD1.n17 104.615
R2487 VDD1.n48 VDD1.n17 104.615
R2488 VDD1.n48 VDD1.n47 104.615
R2489 VDD1.n47 VDD1.n21 104.615
R2490 VDD1.n40 VDD1.n21 104.615
R2491 VDD1.n40 VDD1.n39 104.615
R2492 VDD1.n39 VDD1.n25 104.615
R2493 VDD1.n32 VDD1.n25 104.615
R2494 VDD1.n32 VDD1.n31 104.615
R2495 VDD1.n115 VDD1.n114 104.615
R2496 VDD1.n115 VDD1.n108 104.615
R2497 VDD1.n122 VDD1.n108 104.615
R2498 VDD1.n123 VDD1.n122 104.615
R2499 VDD1.n123 VDD1.n104 104.615
R2500 VDD1.n130 VDD1.n104 104.615
R2501 VDD1.n131 VDD1.n130 104.615
R2502 VDD1.n131 VDD1.n100 104.615
R2503 VDD1.n138 VDD1.n100 104.615
R2504 VDD1.n139 VDD1.n138 104.615
R2505 VDD1.n139 VDD1.n96 104.615
R2506 VDD1.n146 VDD1.n96 104.615
R2507 VDD1.n147 VDD1.n146 104.615
R2508 VDD1.n147 VDD1.n92 104.615
R2509 VDD1.n155 VDD1.n92 104.615
R2510 VDD1.n156 VDD1.n155 104.615
R2511 VDD1.n157 VDD1.n156 104.615
R2512 VDD1.n157 VDD1.n88 104.615
R2513 VDD1.n164 VDD1.n88 104.615
R2514 VDD1.n165 VDD1.n164 104.615
R2515 VDD1.n171 VDD1.n170 61.7181
R2516 VDD1.n173 VDD1.n172 61.0363
R2517 VDD1.n31 VDD1.t2 52.3082
R2518 VDD1.n114 VDD1.t5 52.3082
R2519 VDD1 VDD1.n84 51.3275
R2520 VDD1.n171 VDD1.n169 51.2139
R2521 VDD1.n173 VDD1.n171 48.6043
R2522 VDD1.n30 VDD1.n29 15.6677
R2523 VDD1.n113 VDD1.n112 15.6677
R2524 VDD1.n6 VDD1.n4 13.1884
R2525 VDD1.n158 VDD1.n89 13.1884
R2526 VDD1.n78 VDD1.n77 12.8005
R2527 VDD1.n74 VDD1.n73 12.8005
R2528 VDD1.n33 VDD1.n28 12.8005
R2529 VDD1.n116 VDD1.n111 12.8005
R2530 VDD1.n159 VDD1.n91 12.8005
R2531 VDD1.n163 VDD1.n162 12.8005
R2532 VDD1.n81 VDD1.n2 12.0247
R2533 VDD1.n70 VDD1.n7 12.0247
R2534 VDD1.n34 VDD1.n26 12.0247
R2535 VDD1.n117 VDD1.n109 12.0247
R2536 VDD1.n154 VDD1.n153 12.0247
R2537 VDD1.n166 VDD1.n87 12.0247
R2538 VDD1.n82 VDD1.n0 11.249
R2539 VDD1.n69 VDD1.n10 11.249
R2540 VDD1.n38 VDD1.n37 11.249
R2541 VDD1.n121 VDD1.n120 11.249
R2542 VDD1.n152 VDD1.n93 11.249
R2543 VDD1.n167 VDD1.n85 11.249
R2544 VDD1.n66 VDD1.n65 10.4732
R2545 VDD1.n41 VDD1.n24 10.4732
R2546 VDD1.n124 VDD1.n107 10.4732
R2547 VDD1.n149 VDD1.n148 10.4732
R2548 VDD1.n62 VDD1.n12 9.69747
R2549 VDD1.n42 VDD1.n22 9.69747
R2550 VDD1.n125 VDD1.n105 9.69747
R2551 VDD1.n145 VDD1.n95 9.69747
R2552 VDD1.n84 VDD1.n83 9.45567
R2553 VDD1.n169 VDD1.n168 9.45567
R2554 VDD1.n16 VDD1.n15 9.3005
R2555 VDD1.n59 VDD1.n58 9.3005
R2556 VDD1.n61 VDD1.n60 9.3005
R2557 VDD1.n12 VDD1.n11 9.3005
R2558 VDD1.n67 VDD1.n66 9.3005
R2559 VDD1.n69 VDD1.n68 9.3005
R2560 VDD1.n7 VDD1.n5 9.3005
R2561 VDD1.n75 VDD1.n74 9.3005
R2562 VDD1.n83 VDD1.n82 9.3005
R2563 VDD1.n2 VDD1.n1 9.3005
R2564 VDD1.n77 VDD1.n76 9.3005
R2565 VDD1.n53 VDD1.n52 9.3005
R2566 VDD1.n51 VDD1.n50 9.3005
R2567 VDD1.n20 VDD1.n19 9.3005
R2568 VDD1.n45 VDD1.n44 9.3005
R2569 VDD1.n43 VDD1.n42 9.3005
R2570 VDD1.n24 VDD1.n23 9.3005
R2571 VDD1.n37 VDD1.n36 9.3005
R2572 VDD1.n35 VDD1.n34 9.3005
R2573 VDD1.n28 VDD1.n27 9.3005
R2574 VDD1.n168 VDD1.n167 9.3005
R2575 VDD1.n87 VDD1.n86 9.3005
R2576 VDD1.n162 VDD1.n161 9.3005
R2577 VDD1.n134 VDD1.n133 9.3005
R2578 VDD1.n103 VDD1.n102 9.3005
R2579 VDD1.n128 VDD1.n127 9.3005
R2580 VDD1.n126 VDD1.n125 9.3005
R2581 VDD1.n107 VDD1.n106 9.3005
R2582 VDD1.n120 VDD1.n119 9.3005
R2583 VDD1.n118 VDD1.n117 9.3005
R2584 VDD1.n111 VDD1.n110 9.3005
R2585 VDD1.n136 VDD1.n135 9.3005
R2586 VDD1.n99 VDD1.n98 9.3005
R2587 VDD1.n142 VDD1.n141 9.3005
R2588 VDD1.n144 VDD1.n143 9.3005
R2589 VDD1.n95 VDD1.n94 9.3005
R2590 VDD1.n150 VDD1.n149 9.3005
R2591 VDD1.n152 VDD1.n151 9.3005
R2592 VDD1.n153 VDD1.n90 9.3005
R2593 VDD1.n160 VDD1.n159 9.3005
R2594 VDD1.n61 VDD1.n14 8.92171
R2595 VDD1.n46 VDD1.n45 8.92171
R2596 VDD1.n129 VDD1.n128 8.92171
R2597 VDD1.n144 VDD1.n97 8.92171
R2598 VDD1.n58 VDD1.n57 8.14595
R2599 VDD1.n49 VDD1.n20 8.14595
R2600 VDD1.n132 VDD1.n103 8.14595
R2601 VDD1.n141 VDD1.n140 8.14595
R2602 VDD1.n54 VDD1.n16 7.3702
R2603 VDD1.n50 VDD1.n18 7.3702
R2604 VDD1.n133 VDD1.n101 7.3702
R2605 VDD1.n137 VDD1.n99 7.3702
R2606 VDD1.n54 VDD1.n53 6.59444
R2607 VDD1.n53 VDD1.n18 6.59444
R2608 VDD1.n136 VDD1.n101 6.59444
R2609 VDD1.n137 VDD1.n136 6.59444
R2610 VDD1.n57 VDD1.n16 5.81868
R2611 VDD1.n50 VDD1.n49 5.81868
R2612 VDD1.n133 VDD1.n132 5.81868
R2613 VDD1.n140 VDD1.n99 5.81868
R2614 VDD1.n58 VDD1.n14 5.04292
R2615 VDD1.n46 VDD1.n20 5.04292
R2616 VDD1.n129 VDD1.n103 5.04292
R2617 VDD1.n141 VDD1.n97 5.04292
R2618 VDD1.n29 VDD1.n27 4.38563
R2619 VDD1.n112 VDD1.n110 4.38563
R2620 VDD1.n62 VDD1.n61 4.26717
R2621 VDD1.n45 VDD1.n22 4.26717
R2622 VDD1.n128 VDD1.n105 4.26717
R2623 VDD1.n145 VDD1.n144 4.26717
R2624 VDD1.n65 VDD1.n12 3.49141
R2625 VDD1.n42 VDD1.n41 3.49141
R2626 VDD1.n125 VDD1.n124 3.49141
R2627 VDD1.n148 VDD1.n95 3.49141
R2628 VDD1.n84 VDD1.n0 2.71565
R2629 VDD1.n66 VDD1.n10 2.71565
R2630 VDD1.n38 VDD1.n24 2.71565
R2631 VDD1.n121 VDD1.n107 2.71565
R2632 VDD1.n149 VDD1.n93 2.71565
R2633 VDD1.n169 VDD1.n85 2.71565
R2634 VDD1.n82 VDD1.n81 1.93989
R2635 VDD1.n70 VDD1.n69 1.93989
R2636 VDD1.n37 VDD1.n26 1.93989
R2637 VDD1.n120 VDD1.n109 1.93989
R2638 VDD1.n154 VDD1.n152 1.93989
R2639 VDD1.n167 VDD1.n166 1.93989
R2640 VDD1.n172 VDD1.t1 1.28872
R2641 VDD1.n172 VDD1.t3 1.28872
R2642 VDD1.n170 VDD1.t0 1.28872
R2643 VDD1.n170 VDD1.t4 1.28872
R2644 VDD1.n78 VDD1.n2 1.16414
R2645 VDD1.n73 VDD1.n7 1.16414
R2646 VDD1.n34 VDD1.n33 1.16414
R2647 VDD1.n117 VDD1.n116 1.16414
R2648 VDD1.n153 VDD1.n91 1.16414
R2649 VDD1.n163 VDD1.n87 1.16414
R2650 VDD1 VDD1.n173 0.679379
R2651 VDD1.n77 VDD1.n4 0.388379
R2652 VDD1.n74 VDD1.n6 0.388379
R2653 VDD1.n30 VDD1.n28 0.388379
R2654 VDD1.n113 VDD1.n111 0.388379
R2655 VDD1.n159 VDD1.n158 0.388379
R2656 VDD1.n162 VDD1.n89 0.388379
R2657 VDD1.n83 VDD1.n1 0.155672
R2658 VDD1.n76 VDD1.n1 0.155672
R2659 VDD1.n76 VDD1.n75 0.155672
R2660 VDD1.n75 VDD1.n5 0.155672
R2661 VDD1.n68 VDD1.n5 0.155672
R2662 VDD1.n68 VDD1.n67 0.155672
R2663 VDD1.n67 VDD1.n11 0.155672
R2664 VDD1.n60 VDD1.n11 0.155672
R2665 VDD1.n60 VDD1.n59 0.155672
R2666 VDD1.n59 VDD1.n15 0.155672
R2667 VDD1.n52 VDD1.n15 0.155672
R2668 VDD1.n52 VDD1.n51 0.155672
R2669 VDD1.n51 VDD1.n19 0.155672
R2670 VDD1.n44 VDD1.n19 0.155672
R2671 VDD1.n44 VDD1.n43 0.155672
R2672 VDD1.n43 VDD1.n23 0.155672
R2673 VDD1.n36 VDD1.n23 0.155672
R2674 VDD1.n36 VDD1.n35 0.155672
R2675 VDD1.n35 VDD1.n27 0.155672
R2676 VDD1.n118 VDD1.n110 0.155672
R2677 VDD1.n119 VDD1.n118 0.155672
R2678 VDD1.n119 VDD1.n106 0.155672
R2679 VDD1.n126 VDD1.n106 0.155672
R2680 VDD1.n127 VDD1.n126 0.155672
R2681 VDD1.n127 VDD1.n102 0.155672
R2682 VDD1.n134 VDD1.n102 0.155672
R2683 VDD1.n135 VDD1.n134 0.155672
R2684 VDD1.n135 VDD1.n98 0.155672
R2685 VDD1.n142 VDD1.n98 0.155672
R2686 VDD1.n143 VDD1.n142 0.155672
R2687 VDD1.n143 VDD1.n94 0.155672
R2688 VDD1.n150 VDD1.n94 0.155672
R2689 VDD1.n151 VDD1.n150 0.155672
R2690 VDD1.n151 VDD1.n90 0.155672
R2691 VDD1.n160 VDD1.n90 0.155672
R2692 VDD1.n161 VDD1.n160 0.155672
R2693 VDD1.n161 VDD1.n86 0.155672
R2694 VDD1.n168 VDD1.n86 0.155672
R2695 VN.n30 VN.n29 161.3
R2696 VN.n28 VN.n17 161.3
R2697 VN.n27 VN.n26 161.3
R2698 VN.n25 VN.n18 161.3
R2699 VN.n24 VN.n23 161.3
R2700 VN.n22 VN.n19 161.3
R2701 VN.n14 VN.n13 161.3
R2702 VN.n12 VN.n1 161.3
R2703 VN.n11 VN.n10 161.3
R2704 VN.n9 VN.n2 161.3
R2705 VN.n8 VN.n7 161.3
R2706 VN.n6 VN.n3 161.3
R2707 VN.n20 VN.t2 153.286
R2708 VN.n4 VN.t1 153.286
R2709 VN.n5 VN.t4 119.876
R2710 VN.n0 VN.t0 119.876
R2711 VN.n21 VN.t3 119.876
R2712 VN.n16 VN.t5 119.876
R2713 VN.n15 VN.n0 69.5151
R2714 VN.n31 VN.n16 69.5151
R2715 VN.n11 VN.n2 56.5193
R2716 VN.n27 VN.n18 56.5193
R2717 VN VN.n31 53.4677
R2718 VN.n5 VN.n4 49.4256
R2719 VN.n21 VN.n20 49.4256
R2720 VN.n6 VN.n5 24.4675
R2721 VN.n7 VN.n6 24.4675
R2722 VN.n7 VN.n2 24.4675
R2723 VN.n12 VN.n11 24.4675
R2724 VN.n13 VN.n12 24.4675
R2725 VN.n23 VN.n18 24.4675
R2726 VN.n23 VN.n22 24.4675
R2727 VN.n22 VN.n21 24.4675
R2728 VN.n29 VN.n28 24.4675
R2729 VN.n28 VN.n27 24.4675
R2730 VN.n13 VN.n0 20.5528
R2731 VN.n29 VN.n16 20.5528
R2732 VN.n20 VN.n19 3.88811
R2733 VN.n4 VN.n3 3.88811
R2734 VN.n31 VN.n30 0.354971
R2735 VN.n15 VN.n14 0.354971
R2736 VN VN.n15 0.26696
R2737 VN.n30 VN.n17 0.189894
R2738 VN.n26 VN.n17 0.189894
R2739 VN.n26 VN.n25 0.189894
R2740 VN.n25 VN.n24 0.189894
R2741 VN.n24 VN.n19 0.189894
R2742 VN.n8 VN.n3 0.189894
R2743 VN.n9 VN.n8 0.189894
R2744 VN.n10 VN.n9 0.189894
R2745 VN.n10 VN.n1 0.189894
R2746 VN.n14 VN.n1 0.189894
R2747 VDD2.n167 VDD2.n87 289.615
R2748 VDD2.n80 VDD2.n0 289.615
R2749 VDD2.n168 VDD2.n167 185
R2750 VDD2.n166 VDD2.n165 185
R2751 VDD2.n91 VDD2.n90 185
R2752 VDD2.n95 VDD2.n93 185
R2753 VDD2.n160 VDD2.n159 185
R2754 VDD2.n158 VDD2.n157 185
R2755 VDD2.n97 VDD2.n96 185
R2756 VDD2.n152 VDD2.n151 185
R2757 VDD2.n150 VDD2.n149 185
R2758 VDD2.n101 VDD2.n100 185
R2759 VDD2.n144 VDD2.n143 185
R2760 VDD2.n142 VDD2.n141 185
R2761 VDD2.n105 VDD2.n104 185
R2762 VDD2.n136 VDD2.n135 185
R2763 VDD2.n134 VDD2.n133 185
R2764 VDD2.n109 VDD2.n108 185
R2765 VDD2.n128 VDD2.n127 185
R2766 VDD2.n126 VDD2.n125 185
R2767 VDD2.n113 VDD2.n112 185
R2768 VDD2.n120 VDD2.n119 185
R2769 VDD2.n118 VDD2.n117 185
R2770 VDD2.n29 VDD2.n28 185
R2771 VDD2.n31 VDD2.n30 185
R2772 VDD2.n24 VDD2.n23 185
R2773 VDD2.n37 VDD2.n36 185
R2774 VDD2.n39 VDD2.n38 185
R2775 VDD2.n20 VDD2.n19 185
R2776 VDD2.n45 VDD2.n44 185
R2777 VDD2.n47 VDD2.n46 185
R2778 VDD2.n16 VDD2.n15 185
R2779 VDD2.n53 VDD2.n52 185
R2780 VDD2.n55 VDD2.n54 185
R2781 VDD2.n12 VDD2.n11 185
R2782 VDD2.n61 VDD2.n60 185
R2783 VDD2.n63 VDD2.n62 185
R2784 VDD2.n8 VDD2.n7 185
R2785 VDD2.n70 VDD2.n69 185
R2786 VDD2.n71 VDD2.n6 185
R2787 VDD2.n73 VDD2.n72 185
R2788 VDD2.n4 VDD2.n3 185
R2789 VDD2.n79 VDD2.n78 185
R2790 VDD2.n81 VDD2.n80 185
R2791 VDD2.n116 VDD2.t0 147.659
R2792 VDD2.n27 VDD2.t4 147.659
R2793 VDD2.n167 VDD2.n166 104.615
R2794 VDD2.n166 VDD2.n90 104.615
R2795 VDD2.n95 VDD2.n90 104.615
R2796 VDD2.n159 VDD2.n95 104.615
R2797 VDD2.n159 VDD2.n158 104.615
R2798 VDD2.n158 VDD2.n96 104.615
R2799 VDD2.n151 VDD2.n96 104.615
R2800 VDD2.n151 VDD2.n150 104.615
R2801 VDD2.n150 VDD2.n100 104.615
R2802 VDD2.n143 VDD2.n100 104.615
R2803 VDD2.n143 VDD2.n142 104.615
R2804 VDD2.n142 VDD2.n104 104.615
R2805 VDD2.n135 VDD2.n104 104.615
R2806 VDD2.n135 VDD2.n134 104.615
R2807 VDD2.n134 VDD2.n108 104.615
R2808 VDD2.n127 VDD2.n108 104.615
R2809 VDD2.n127 VDD2.n126 104.615
R2810 VDD2.n126 VDD2.n112 104.615
R2811 VDD2.n119 VDD2.n112 104.615
R2812 VDD2.n119 VDD2.n118 104.615
R2813 VDD2.n30 VDD2.n29 104.615
R2814 VDD2.n30 VDD2.n23 104.615
R2815 VDD2.n37 VDD2.n23 104.615
R2816 VDD2.n38 VDD2.n37 104.615
R2817 VDD2.n38 VDD2.n19 104.615
R2818 VDD2.n45 VDD2.n19 104.615
R2819 VDD2.n46 VDD2.n45 104.615
R2820 VDD2.n46 VDD2.n15 104.615
R2821 VDD2.n53 VDD2.n15 104.615
R2822 VDD2.n54 VDD2.n53 104.615
R2823 VDD2.n54 VDD2.n11 104.615
R2824 VDD2.n61 VDD2.n11 104.615
R2825 VDD2.n62 VDD2.n61 104.615
R2826 VDD2.n62 VDD2.n7 104.615
R2827 VDD2.n70 VDD2.n7 104.615
R2828 VDD2.n71 VDD2.n70 104.615
R2829 VDD2.n72 VDD2.n71 104.615
R2830 VDD2.n72 VDD2.n3 104.615
R2831 VDD2.n79 VDD2.n3 104.615
R2832 VDD2.n80 VDD2.n79 104.615
R2833 VDD2.n86 VDD2.n85 61.7181
R2834 VDD2 VDD2.n173 61.7152
R2835 VDD2.n118 VDD2.t0 52.3082
R2836 VDD2.n29 VDD2.t4 52.3082
R2837 VDD2.n86 VDD2.n84 51.2139
R2838 VDD2.n172 VDD2.n171 49.0581
R2839 VDD2.n172 VDD2.n86 46.5472
R2840 VDD2.n117 VDD2.n116 15.6677
R2841 VDD2.n28 VDD2.n27 15.6677
R2842 VDD2.n93 VDD2.n91 13.1884
R2843 VDD2.n73 VDD2.n4 13.1884
R2844 VDD2.n165 VDD2.n164 12.8005
R2845 VDD2.n161 VDD2.n160 12.8005
R2846 VDD2.n120 VDD2.n115 12.8005
R2847 VDD2.n31 VDD2.n26 12.8005
R2848 VDD2.n74 VDD2.n6 12.8005
R2849 VDD2.n78 VDD2.n77 12.8005
R2850 VDD2.n168 VDD2.n89 12.0247
R2851 VDD2.n157 VDD2.n94 12.0247
R2852 VDD2.n121 VDD2.n113 12.0247
R2853 VDD2.n32 VDD2.n24 12.0247
R2854 VDD2.n69 VDD2.n68 12.0247
R2855 VDD2.n81 VDD2.n2 12.0247
R2856 VDD2.n169 VDD2.n87 11.249
R2857 VDD2.n156 VDD2.n97 11.249
R2858 VDD2.n125 VDD2.n124 11.249
R2859 VDD2.n36 VDD2.n35 11.249
R2860 VDD2.n67 VDD2.n8 11.249
R2861 VDD2.n82 VDD2.n0 11.249
R2862 VDD2.n153 VDD2.n152 10.4732
R2863 VDD2.n128 VDD2.n111 10.4732
R2864 VDD2.n39 VDD2.n22 10.4732
R2865 VDD2.n64 VDD2.n63 10.4732
R2866 VDD2.n149 VDD2.n99 9.69747
R2867 VDD2.n129 VDD2.n109 9.69747
R2868 VDD2.n40 VDD2.n20 9.69747
R2869 VDD2.n60 VDD2.n10 9.69747
R2870 VDD2.n171 VDD2.n170 9.45567
R2871 VDD2.n84 VDD2.n83 9.45567
R2872 VDD2.n103 VDD2.n102 9.3005
R2873 VDD2.n146 VDD2.n145 9.3005
R2874 VDD2.n148 VDD2.n147 9.3005
R2875 VDD2.n99 VDD2.n98 9.3005
R2876 VDD2.n154 VDD2.n153 9.3005
R2877 VDD2.n156 VDD2.n155 9.3005
R2878 VDD2.n94 VDD2.n92 9.3005
R2879 VDD2.n162 VDD2.n161 9.3005
R2880 VDD2.n170 VDD2.n169 9.3005
R2881 VDD2.n89 VDD2.n88 9.3005
R2882 VDD2.n164 VDD2.n163 9.3005
R2883 VDD2.n140 VDD2.n139 9.3005
R2884 VDD2.n138 VDD2.n137 9.3005
R2885 VDD2.n107 VDD2.n106 9.3005
R2886 VDD2.n132 VDD2.n131 9.3005
R2887 VDD2.n130 VDD2.n129 9.3005
R2888 VDD2.n111 VDD2.n110 9.3005
R2889 VDD2.n124 VDD2.n123 9.3005
R2890 VDD2.n122 VDD2.n121 9.3005
R2891 VDD2.n115 VDD2.n114 9.3005
R2892 VDD2.n83 VDD2.n82 9.3005
R2893 VDD2.n2 VDD2.n1 9.3005
R2894 VDD2.n77 VDD2.n76 9.3005
R2895 VDD2.n49 VDD2.n48 9.3005
R2896 VDD2.n18 VDD2.n17 9.3005
R2897 VDD2.n43 VDD2.n42 9.3005
R2898 VDD2.n41 VDD2.n40 9.3005
R2899 VDD2.n22 VDD2.n21 9.3005
R2900 VDD2.n35 VDD2.n34 9.3005
R2901 VDD2.n33 VDD2.n32 9.3005
R2902 VDD2.n26 VDD2.n25 9.3005
R2903 VDD2.n51 VDD2.n50 9.3005
R2904 VDD2.n14 VDD2.n13 9.3005
R2905 VDD2.n57 VDD2.n56 9.3005
R2906 VDD2.n59 VDD2.n58 9.3005
R2907 VDD2.n10 VDD2.n9 9.3005
R2908 VDD2.n65 VDD2.n64 9.3005
R2909 VDD2.n67 VDD2.n66 9.3005
R2910 VDD2.n68 VDD2.n5 9.3005
R2911 VDD2.n75 VDD2.n74 9.3005
R2912 VDD2.n148 VDD2.n101 8.92171
R2913 VDD2.n133 VDD2.n132 8.92171
R2914 VDD2.n44 VDD2.n43 8.92171
R2915 VDD2.n59 VDD2.n12 8.92171
R2916 VDD2.n145 VDD2.n144 8.14595
R2917 VDD2.n136 VDD2.n107 8.14595
R2918 VDD2.n47 VDD2.n18 8.14595
R2919 VDD2.n56 VDD2.n55 8.14595
R2920 VDD2.n141 VDD2.n103 7.3702
R2921 VDD2.n137 VDD2.n105 7.3702
R2922 VDD2.n48 VDD2.n16 7.3702
R2923 VDD2.n52 VDD2.n14 7.3702
R2924 VDD2.n141 VDD2.n140 6.59444
R2925 VDD2.n140 VDD2.n105 6.59444
R2926 VDD2.n51 VDD2.n16 6.59444
R2927 VDD2.n52 VDD2.n51 6.59444
R2928 VDD2.n144 VDD2.n103 5.81868
R2929 VDD2.n137 VDD2.n136 5.81868
R2930 VDD2.n48 VDD2.n47 5.81868
R2931 VDD2.n55 VDD2.n14 5.81868
R2932 VDD2.n145 VDD2.n101 5.04292
R2933 VDD2.n133 VDD2.n107 5.04292
R2934 VDD2.n44 VDD2.n18 5.04292
R2935 VDD2.n56 VDD2.n12 5.04292
R2936 VDD2.n116 VDD2.n114 4.38563
R2937 VDD2.n27 VDD2.n25 4.38563
R2938 VDD2.n149 VDD2.n148 4.26717
R2939 VDD2.n132 VDD2.n109 4.26717
R2940 VDD2.n43 VDD2.n20 4.26717
R2941 VDD2.n60 VDD2.n59 4.26717
R2942 VDD2.n152 VDD2.n99 3.49141
R2943 VDD2.n129 VDD2.n128 3.49141
R2944 VDD2.n40 VDD2.n39 3.49141
R2945 VDD2.n63 VDD2.n10 3.49141
R2946 VDD2.n171 VDD2.n87 2.71565
R2947 VDD2.n153 VDD2.n97 2.71565
R2948 VDD2.n125 VDD2.n111 2.71565
R2949 VDD2.n36 VDD2.n22 2.71565
R2950 VDD2.n64 VDD2.n8 2.71565
R2951 VDD2.n84 VDD2.n0 2.71565
R2952 VDD2 VDD2.n172 2.2699
R2953 VDD2.n169 VDD2.n168 1.93989
R2954 VDD2.n157 VDD2.n156 1.93989
R2955 VDD2.n124 VDD2.n113 1.93989
R2956 VDD2.n35 VDD2.n24 1.93989
R2957 VDD2.n69 VDD2.n67 1.93989
R2958 VDD2.n82 VDD2.n81 1.93989
R2959 VDD2.n173 VDD2.t2 1.28872
R2960 VDD2.n173 VDD2.t3 1.28872
R2961 VDD2.n85 VDD2.t1 1.28872
R2962 VDD2.n85 VDD2.t5 1.28872
R2963 VDD2.n165 VDD2.n89 1.16414
R2964 VDD2.n160 VDD2.n94 1.16414
R2965 VDD2.n121 VDD2.n120 1.16414
R2966 VDD2.n32 VDD2.n31 1.16414
R2967 VDD2.n68 VDD2.n6 1.16414
R2968 VDD2.n78 VDD2.n2 1.16414
R2969 VDD2.n164 VDD2.n91 0.388379
R2970 VDD2.n161 VDD2.n93 0.388379
R2971 VDD2.n117 VDD2.n115 0.388379
R2972 VDD2.n28 VDD2.n26 0.388379
R2973 VDD2.n74 VDD2.n73 0.388379
R2974 VDD2.n77 VDD2.n4 0.388379
R2975 VDD2.n170 VDD2.n88 0.155672
R2976 VDD2.n163 VDD2.n88 0.155672
R2977 VDD2.n163 VDD2.n162 0.155672
R2978 VDD2.n162 VDD2.n92 0.155672
R2979 VDD2.n155 VDD2.n92 0.155672
R2980 VDD2.n155 VDD2.n154 0.155672
R2981 VDD2.n154 VDD2.n98 0.155672
R2982 VDD2.n147 VDD2.n98 0.155672
R2983 VDD2.n147 VDD2.n146 0.155672
R2984 VDD2.n146 VDD2.n102 0.155672
R2985 VDD2.n139 VDD2.n102 0.155672
R2986 VDD2.n139 VDD2.n138 0.155672
R2987 VDD2.n138 VDD2.n106 0.155672
R2988 VDD2.n131 VDD2.n106 0.155672
R2989 VDD2.n131 VDD2.n130 0.155672
R2990 VDD2.n130 VDD2.n110 0.155672
R2991 VDD2.n123 VDD2.n110 0.155672
R2992 VDD2.n123 VDD2.n122 0.155672
R2993 VDD2.n122 VDD2.n114 0.155672
R2994 VDD2.n33 VDD2.n25 0.155672
R2995 VDD2.n34 VDD2.n33 0.155672
R2996 VDD2.n34 VDD2.n21 0.155672
R2997 VDD2.n41 VDD2.n21 0.155672
R2998 VDD2.n42 VDD2.n41 0.155672
R2999 VDD2.n42 VDD2.n17 0.155672
R3000 VDD2.n49 VDD2.n17 0.155672
R3001 VDD2.n50 VDD2.n49 0.155672
R3002 VDD2.n50 VDD2.n13 0.155672
R3003 VDD2.n57 VDD2.n13 0.155672
R3004 VDD2.n58 VDD2.n57 0.155672
R3005 VDD2.n58 VDD2.n9 0.155672
R3006 VDD2.n65 VDD2.n9 0.155672
R3007 VDD2.n66 VDD2.n65 0.155672
R3008 VDD2.n66 VDD2.n5 0.155672
R3009 VDD2.n75 VDD2.n5 0.155672
R3010 VDD2.n76 VDD2.n75 0.155672
R3011 VDD2.n76 VDD2.n1 0.155672
R3012 VDD2.n83 VDD2.n1 0.155672
C0 VDD1 VP 9.111269f
C1 VTAIL VN 8.88949f
C2 VDD2 VTAIL 9.06001f
C3 VDD1 VN 0.151498f
C4 VDD2 VDD1 1.59902f
C5 VP VN 8.02738f
C6 VDD2 VP 0.500187f
C7 VDD2 VN 8.766179f
C8 VTAIL VDD1 9.006081f
C9 VTAIL VP 8.90379f
C10 VDD2 B 6.960328f
C11 VDD1 B 7.109957f
C12 VTAIL B 9.505937f
C13 VN B 14.598689f
C14 VP B 13.229697f
C15 VDD2.n0 B 0.027786f
C16 VDD2.n1 B 0.021302f
C17 VDD2.n2 B 0.011447f
C18 VDD2.n3 B 0.027056f
C19 VDD2.n4 B 0.011783f
C20 VDD2.n5 B 0.021302f
C21 VDD2.n6 B 0.01212f
C22 VDD2.n7 B 0.027056f
C23 VDD2.n8 B 0.01212f
C24 VDD2.n9 B 0.021302f
C25 VDD2.n10 B 0.011447f
C26 VDD2.n11 B 0.027056f
C27 VDD2.n12 B 0.01212f
C28 VDD2.n13 B 0.021302f
C29 VDD2.n14 B 0.011447f
C30 VDD2.n15 B 0.027056f
C31 VDD2.n16 B 0.01212f
C32 VDD2.n17 B 0.021302f
C33 VDD2.n18 B 0.011447f
C34 VDD2.n19 B 0.027056f
C35 VDD2.n20 B 0.01212f
C36 VDD2.n21 B 0.021302f
C37 VDD2.n22 B 0.011447f
C38 VDD2.n23 B 0.027056f
C39 VDD2.n24 B 0.01212f
C40 VDD2.n25 B 1.42204f
C41 VDD2.n26 B 0.011447f
C42 VDD2.t4 B 0.044638f
C43 VDD2.n27 B 0.14091f
C44 VDD2.n28 B 0.015983f
C45 VDD2.n29 B 0.020292f
C46 VDD2.n30 B 0.027056f
C47 VDD2.n31 B 0.01212f
C48 VDD2.n32 B 0.011447f
C49 VDD2.n33 B 0.021302f
C50 VDD2.n34 B 0.021302f
C51 VDD2.n35 B 0.011447f
C52 VDD2.n36 B 0.01212f
C53 VDD2.n37 B 0.027056f
C54 VDD2.n38 B 0.027056f
C55 VDD2.n39 B 0.01212f
C56 VDD2.n40 B 0.011447f
C57 VDD2.n41 B 0.021302f
C58 VDD2.n42 B 0.021302f
C59 VDD2.n43 B 0.011447f
C60 VDD2.n44 B 0.01212f
C61 VDD2.n45 B 0.027056f
C62 VDD2.n46 B 0.027056f
C63 VDD2.n47 B 0.01212f
C64 VDD2.n48 B 0.011447f
C65 VDD2.n49 B 0.021302f
C66 VDD2.n50 B 0.021302f
C67 VDD2.n51 B 0.011447f
C68 VDD2.n52 B 0.01212f
C69 VDD2.n53 B 0.027056f
C70 VDD2.n54 B 0.027056f
C71 VDD2.n55 B 0.01212f
C72 VDD2.n56 B 0.011447f
C73 VDD2.n57 B 0.021302f
C74 VDD2.n58 B 0.021302f
C75 VDD2.n59 B 0.011447f
C76 VDD2.n60 B 0.01212f
C77 VDD2.n61 B 0.027056f
C78 VDD2.n62 B 0.027056f
C79 VDD2.n63 B 0.01212f
C80 VDD2.n64 B 0.011447f
C81 VDD2.n65 B 0.021302f
C82 VDD2.n66 B 0.021302f
C83 VDD2.n67 B 0.011447f
C84 VDD2.n68 B 0.011447f
C85 VDD2.n69 B 0.01212f
C86 VDD2.n70 B 0.027056f
C87 VDD2.n71 B 0.027056f
C88 VDD2.n72 B 0.027056f
C89 VDD2.n73 B 0.011783f
C90 VDD2.n74 B 0.011447f
C91 VDD2.n75 B 0.021302f
C92 VDD2.n76 B 0.021302f
C93 VDD2.n77 B 0.011447f
C94 VDD2.n78 B 0.01212f
C95 VDD2.n79 B 0.027056f
C96 VDD2.n80 B 0.054759f
C97 VDD2.n81 B 0.01212f
C98 VDD2.n82 B 0.011447f
C99 VDD2.n83 B 0.049529f
C100 VDD2.n84 B 0.052935f
C101 VDD2.t1 B 0.258727f
C102 VDD2.t5 B 0.258727f
C103 VDD2.n85 B 2.34616f
C104 VDD2.n86 B 2.64036f
C105 VDD2.n87 B 0.027786f
C106 VDD2.n88 B 0.021302f
C107 VDD2.n89 B 0.011447f
C108 VDD2.n90 B 0.027056f
C109 VDD2.n91 B 0.011783f
C110 VDD2.n92 B 0.021302f
C111 VDD2.n93 B 0.011783f
C112 VDD2.n94 B 0.011447f
C113 VDD2.n95 B 0.027056f
C114 VDD2.n96 B 0.027056f
C115 VDD2.n97 B 0.01212f
C116 VDD2.n98 B 0.021302f
C117 VDD2.n99 B 0.011447f
C118 VDD2.n100 B 0.027056f
C119 VDD2.n101 B 0.01212f
C120 VDD2.n102 B 0.021302f
C121 VDD2.n103 B 0.011447f
C122 VDD2.n104 B 0.027056f
C123 VDD2.n105 B 0.01212f
C124 VDD2.n106 B 0.021302f
C125 VDD2.n107 B 0.011447f
C126 VDD2.n108 B 0.027056f
C127 VDD2.n109 B 0.01212f
C128 VDD2.n110 B 0.021302f
C129 VDD2.n111 B 0.011447f
C130 VDD2.n112 B 0.027056f
C131 VDD2.n113 B 0.01212f
C132 VDD2.n114 B 1.42204f
C133 VDD2.n115 B 0.011447f
C134 VDD2.t0 B 0.044638f
C135 VDD2.n116 B 0.14091f
C136 VDD2.n117 B 0.015983f
C137 VDD2.n118 B 0.020292f
C138 VDD2.n119 B 0.027056f
C139 VDD2.n120 B 0.01212f
C140 VDD2.n121 B 0.011447f
C141 VDD2.n122 B 0.021302f
C142 VDD2.n123 B 0.021302f
C143 VDD2.n124 B 0.011447f
C144 VDD2.n125 B 0.01212f
C145 VDD2.n126 B 0.027056f
C146 VDD2.n127 B 0.027056f
C147 VDD2.n128 B 0.01212f
C148 VDD2.n129 B 0.011447f
C149 VDD2.n130 B 0.021302f
C150 VDD2.n131 B 0.021302f
C151 VDD2.n132 B 0.011447f
C152 VDD2.n133 B 0.01212f
C153 VDD2.n134 B 0.027056f
C154 VDD2.n135 B 0.027056f
C155 VDD2.n136 B 0.01212f
C156 VDD2.n137 B 0.011447f
C157 VDD2.n138 B 0.021302f
C158 VDD2.n139 B 0.021302f
C159 VDD2.n140 B 0.011447f
C160 VDD2.n141 B 0.01212f
C161 VDD2.n142 B 0.027056f
C162 VDD2.n143 B 0.027056f
C163 VDD2.n144 B 0.01212f
C164 VDD2.n145 B 0.011447f
C165 VDD2.n146 B 0.021302f
C166 VDD2.n147 B 0.021302f
C167 VDD2.n148 B 0.011447f
C168 VDD2.n149 B 0.01212f
C169 VDD2.n150 B 0.027056f
C170 VDD2.n151 B 0.027056f
C171 VDD2.n152 B 0.01212f
C172 VDD2.n153 B 0.011447f
C173 VDD2.n154 B 0.021302f
C174 VDD2.n155 B 0.021302f
C175 VDD2.n156 B 0.011447f
C176 VDD2.n157 B 0.01212f
C177 VDD2.n158 B 0.027056f
C178 VDD2.n159 B 0.027056f
C179 VDD2.n160 B 0.01212f
C180 VDD2.n161 B 0.011447f
C181 VDD2.n162 B 0.021302f
C182 VDD2.n163 B 0.021302f
C183 VDD2.n164 B 0.011447f
C184 VDD2.n165 B 0.01212f
C185 VDD2.n166 B 0.027056f
C186 VDD2.n167 B 0.054759f
C187 VDD2.n168 B 0.01212f
C188 VDD2.n169 B 0.011447f
C189 VDD2.n170 B 0.049529f
C190 VDD2.n171 B 0.044963f
C191 VDD2.n172 B 2.51656f
C192 VDD2.t2 B 0.258727f
C193 VDD2.t3 B 0.258727f
C194 VDD2.n173 B 2.34613f
C195 VN.t0 B 2.62474f
C196 VN.n0 B 0.995394f
C197 VN.n1 B 0.020157f
C198 VN.n2 B 0.027179f
C199 VN.n3 B 0.229378f
C200 VN.t4 B 2.62474f
C201 VN.t1 B 2.85501f
C202 VN.n4 B 0.942798f
C203 VN.n5 B 0.988602f
C204 VN.n6 B 0.037569f
C205 VN.n7 B 0.037569f
C206 VN.n8 B 0.020157f
C207 VN.n9 B 0.020157f
C208 VN.n10 B 0.020157f
C209 VN.n11 B 0.031673f
C210 VN.n12 B 0.037569f
C211 VN.n13 B 0.034601f
C212 VN.n14 B 0.032534f
C213 VN.n15 B 0.042019f
C214 VN.t5 B 2.62474f
C215 VN.n16 B 0.995394f
C216 VN.n17 B 0.020157f
C217 VN.n18 B 0.027179f
C218 VN.n19 B 0.229378f
C219 VN.t3 B 2.62474f
C220 VN.t2 B 2.85501f
C221 VN.n20 B 0.942798f
C222 VN.n21 B 0.988602f
C223 VN.n22 B 0.037569f
C224 VN.n23 B 0.037569f
C225 VN.n24 B 0.020157f
C226 VN.n25 B 0.020157f
C227 VN.n26 B 0.020157f
C228 VN.n27 B 0.031673f
C229 VN.n28 B 0.037569f
C230 VN.n29 B 0.034601f
C231 VN.n30 B 0.032534f
C232 VN.n31 B 1.25711f
C233 VDD1.n0 B 0.027973f
C234 VDD1.n1 B 0.021445f
C235 VDD1.n2 B 0.011524f
C236 VDD1.n3 B 0.027238f
C237 VDD1.n4 B 0.011863f
C238 VDD1.n5 B 0.021445f
C239 VDD1.n6 B 0.011863f
C240 VDD1.n7 B 0.011524f
C241 VDD1.n8 B 0.027238f
C242 VDD1.n9 B 0.027238f
C243 VDD1.n10 B 0.012202f
C244 VDD1.n11 B 0.021445f
C245 VDD1.n12 B 0.011524f
C246 VDD1.n13 B 0.027238f
C247 VDD1.n14 B 0.012202f
C248 VDD1.n15 B 0.021445f
C249 VDD1.n16 B 0.011524f
C250 VDD1.n17 B 0.027238f
C251 VDD1.n18 B 0.012202f
C252 VDD1.n19 B 0.021445f
C253 VDD1.n20 B 0.011524f
C254 VDD1.n21 B 0.027238f
C255 VDD1.n22 B 0.012202f
C256 VDD1.n23 B 0.021445f
C257 VDD1.n24 B 0.011524f
C258 VDD1.n25 B 0.027238f
C259 VDD1.n26 B 0.012202f
C260 VDD1.n27 B 1.43164f
C261 VDD1.n28 B 0.011524f
C262 VDD1.t2 B 0.04494f
C263 VDD1.n29 B 0.141861f
C264 VDD1.n30 B 0.01609f
C265 VDD1.n31 B 0.020429f
C266 VDD1.n32 B 0.027238f
C267 VDD1.n33 B 0.012202f
C268 VDD1.n34 B 0.011524f
C269 VDD1.n35 B 0.021445f
C270 VDD1.n36 B 0.021445f
C271 VDD1.n37 B 0.011524f
C272 VDD1.n38 B 0.012202f
C273 VDD1.n39 B 0.027238f
C274 VDD1.n40 B 0.027238f
C275 VDD1.n41 B 0.012202f
C276 VDD1.n42 B 0.011524f
C277 VDD1.n43 B 0.021445f
C278 VDD1.n44 B 0.021445f
C279 VDD1.n45 B 0.011524f
C280 VDD1.n46 B 0.012202f
C281 VDD1.n47 B 0.027238f
C282 VDD1.n48 B 0.027238f
C283 VDD1.n49 B 0.012202f
C284 VDD1.n50 B 0.011524f
C285 VDD1.n51 B 0.021445f
C286 VDD1.n52 B 0.021445f
C287 VDD1.n53 B 0.011524f
C288 VDD1.n54 B 0.012202f
C289 VDD1.n55 B 0.027238f
C290 VDD1.n56 B 0.027238f
C291 VDD1.n57 B 0.012202f
C292 VDD1.n58 B 0.011524f
C293 VDD1.n59 B 0.021445f
C294 VDD1.n60 B 0.021445f
C295 VDD1.n61 B 0.011524f
C296 VDD1.n62 B 0.012202f
C297 VDD1.n63 B 0.027238f
C298 VDD1.n64 B 0.027238f
C299 VDD1.n65 B 0.012202f
C300 VDD1.n66 B 0.011524f
C301 VDD1.n67 B 0.021445f
C302 VDD1.n68 B 0.021445f
C303 VDD1.n69 B 0.011524f
C304 VDD1.n70 B 0.012202f
C305 VDD1.n71 B 0.027238f
C306 VDD1.n72 B 0.027238f
C307 VDD1.n73 B 0.012202f
C308 VDD1.n74 B 0.011524f
C309 VDD1.n75 B 0.021445f
C310 VDD1.n76 B 0.021445f
C311 VDD1.n77 B 0.011524f
C312 VDD1.n78 B 0.012202f
C313 VDD1.n79 B 0.027238f
C314 VDD1.n80 B 0.055128f
C315 VDD1.n81 B 0.012202f
C316 VDD1.n82 B 0.011524f
C317 VDD1.n83 B 0.049863f
C318 VDD1.n84 B 0.054033f
C319 VDD1.n85 B 0.027973f
C320 VDD1.n86 B 0.021445f
C321 VDD1.n87 B 0.011524f
C322 VDD1.n88 B 0.027238f
C323 VDD1.n89 B 0.011863f
C324 VDD1.n90 B 0.021445f
C325 VDD1.n91 B 0.012202f
C326 VDD1.n92 B 0.027238f
C327 VDD1.n93 B 0.012202f
C328 VDD1.n94 B 0.021445f
C329 VDD1.n95 B 0.011524f
C330 VDD1.n96 B 0.027238f
C331 VDD1.n97 B 0.012202f
C332 VDD1.n98 B 0.021445f
C333 VDD1.n99 B 0.011524f
C334 VDD1.n100 B 0.027238f
C335 VDD1.n101 B 0.012202f
C336 VDD1.n102 B 0.021445f
C337 VDD1.n103 B 0.011524f
C338 VDD1.n104 B 0.027238f
C339 VDD1.n105 B 0.012202f
C340 VDD1.n106 B 0.021445f
C341 VDD1.n107 B 0.011524f
C342 VDD1.n108 B 0.027238f
C343 VDD1.n109 B 0.012202f
C344 VDD1.n110 B 1.43164f
C345 VDD1.n111 B 0.011524f
C346 VDD1.t5 B 0.04494f
C347 VDD1.n112 B 0.141861f
C348 VDD1.n113 B 0.01609f
C349 VDD1.n114 B 0.020429f
C350 VDD1.n115 B 0.027238f
C351 VDD1.n116 B 0.012202f
C352 VDD1.n117 B 0.011524f
C353 VDD1.n118 B 0.021445f
C354 VDD1.n119 B 0.021445f
C355 VDD1.n120 B 0.011524f
C356 VDD1.n121 B 0.012202f
C357 VDD1.n122 B 0.027238f
C358 VDD1.n123 B 0.027238f
C359 VDD1.n124 B 0.012202f
C360 VDD1.n125 B 0.011524f
C361 VDD1.n126 B 0.021445f
C362 VDD1.n127 B 0.021445f
C363 VDD1.n128 B 0.011524f
C364 VDD1.n129 B 0.012202f
C365 VDD1.n130 B 0.027238f
C366 VDD1.n131 B 0.027238f
C367 VDD1.n132 B 0.012202f
C368 VDD1.n133 B 0.011524f
C369 VDD1.n134 B 0.021445f
C370 VDD1.n135 B 0.021445f
C371 VDD1.n136 B 0.011524f
C372 VDD1.n137 B 0.012202f
C373 VDD1.n138 B 0.027238f
C374 VDD1.n139 B 0.027238f
C375 VDD1.n140 B 0.012202f
C376 VDD1.n141 B 0.011524f
C377 VDD1.n142 B 0.021445f
C378 VDD1.n143 B 0.021445f
C379 VDD1.n144 B 0.011524f
C380 VDD1.n145 B 0.012202f
C381 VDD1.n146 B 0.027238f
C382 VDD1.n147 B 0.027238f
C383 VDD1.n148 B 0.012202f
C384 VDD1.n149 B 0.011524f
C385 VDD1.n150 B 0.021445f
C386 VDD1.n151 B 0.021445f
C387 VDD1.n152 B 0.011524f
C388 VDD1.n153 B 0.011524f
C389 VDD1.n154 B 0.012202f
C390 VDD1.n155 B 0.027238f
C391 VDD1.n156 B 0.027238f
C392 VDD1.n157 B 0.027238f
C393 VDD1.n158 B 0.011863f
C394 VDD1.n159 B 0.011524f
C395 VDD1.n160 B 0.021445f
C396 VDD1.n161 B 0.021445f
C397 VDD1.n162 B 0.011524f
C398 VDD1.n163 B 0.012202f
C399 VDD1.n164 B 0.027238f
C400 VDD1.n165 B 0.055128f
C401 VDD1.n166 B 0.012202f
C402 VDD1.n167 B 0.011524f
C403 VDD1.n168 B 0.049863f
C404 VDD1.n169 B 0.053292f
C405 VDD1.t0 B 0.260473f
C406 VDD1.t4 B 0.260473f
C407 VDD1.n170 B 2.362f
C408 VDD1.n171 B 2.77799f
C409 VDD1.t1 B 0.260473f
C410 VDD1.t3 B 0.260473f
C411 VDD1.n172 B 2.35718f
C412 VDD1.n173 B 2.72977f
C413 VTAIL.t1 B 0.281882f
C414 VTAIL.t11 B 0.281882f
C415 VTAIL.n0 B 2.48103f
C416 VTAIL.n1 B 0.433469f
C417 VTAIL.n2 B 0.030272f
C418 VTAIL.n3 B 0.023208f
C419 VTAIL.n4 B 0.012471f
C420 VTAIL.n5 B 0.029477f
C421 VTAIL.n6 B 0.012838f
C422 VTAIL.n7 B 0.023208f
C423 VTAIL.n8 B 0.013205f
C424 VTAIL.n9 B 0.029477f
C425 VTAIL.n10 B 0.013205f
C426 VTAIL.n11 B 0.023208f
C427 VTAIL.n12 B 0.012471f
C428 VTAIL.n13 B 0.029477f
C429 VTAIL.n14 B 0.013205f
C430 VTAIL.n15 B 0.023208f
C431 VTAIL.n16 B 0.012471f
C432 VTAIL.n17 B 0.029477f
C433 VTAIL.n18 B 0.013205f
C434 VTAIL.n19 B 0.023208f
C435 VTAIL.n20 B 0.012471f
C436 VTAIL.n21 B 0.029477f
C437 VTAIL.n22 B 0.013205f
C438 VTAIL.n23 B 0.023208f
C439 VTAIL.n24 B 0.012471f
C440 VTAIL.n25 B 0.029477f
C441 VTAIL.n26 B 0.013205f
C442 VTAIL.n27 B 1.54931f
C443 VTAIL.n28 B 0.012471f
C444 VTAIL.t4 B 0.048633f
C445 VTAIL.n29 B 0.153521f
C446 VTAIL.n30 B 0.017413f
C447 VTAIL.n31 B 0.022108f
C448 VTAIL.n32 B 0.029477f
C449 VTAIL.n33 B 0.013205f
C450 VTAIL.n34 B 0.012471f
C451 VTAIL.n35 B 0.023208f
C452 VTAIL.n36 B 0.023208f
C453 VTAIL.n37 B 0.012471f
C454 VTAIL.n38 B 0.013205f
C455 VTAIL.n39 B 0.029477f
C456 VTAIL.n40 B 0.029477f
C457 VTAIL.n41 B 0.013205f
C458 VTAIL.n42 B 0.012471f
C459 VTAIL.n43 B 0.023208f
C460 VTAIL.n44 B 0.023208f
C461 VTAIL.n45 B 0.012471f
C462 VTAIL.n46 B 0.013205f
C463 VTAIL.n47 B 0.029477f
C464 VTAIL.n48 B 0.029477f
C465 VTAIL.n49 B 0.013205f
C466 VTAIL.n50 B 0.012471f
C467 VTAIL.n51 B 0.023208f
C468 VTAIL.n52 B 0.023208f
C469 VTAIL.n53 B 0.012471f
C470 VTAIL.n54 B 0.013205f
C471 VTAIL.n55 B 0.029477f
C472 VTAIL.n56 B 0.029477f
C473 VTAIL.n57 B 0.013205f
C474 VTAIL.n58 B 0.012471f
C475 VTAIL.n59 B 0.023208f
C476 VTAIL.n60 B 0.023208f
C477 VTAIL.n61 B 0.012471f
C478 VTAIL.n62 B 0.013205f
C479 VTAIL.n63 B 0.029477f
C480 VTAIL.n64 B 0.029477f
C481 VTAIL.n65 B 0.013205f
C482 VTAIL.n66 B 0.012471f
C483 VTAIL.n67 B 0.023208f
C484 VTAIL.n68 B 0.023208f
C485 VTAIL.n69 B 0.012471f
C486 VTAIL.n70 B 0.012471f
C487 VTAIL.n71 B 0.013205f
C488 VTAIL.n72 B 0.029477f
C489 VTAIL.n73 B 0.029477f
C490 VTAIL.n74 B 0.029477f
C491 VTAIL.n75 B 0.012838f
C492 VTAIL.n76 B 0.012471f
C493 VTAIL.n77 B 0.023208f
C494 VTAIL.n78 B 0.023208f
C495 VTAIL.n79 B 0.012471f
C496 VTAIL.n80 B 0.013205f
C497 VTAIL.n81 B 0.029477f
C498 VTAIL.n82 B 0.059659f
C499 VTAIL.n83 B 0.013205f
C500 VTAIL.n84 B 0.012471f
C501 VTAIL.n85 B 0.053961f
C502 VTAIL.n86 B 0.032965f
C503 VTAIL.n87 B 0.38585f
C504 VTAIL.t6 B 0.281882f
C505 VTAIL.t5 B 0.281882f
C506 VTAIL.n88 B 2.48103f
C507 VTAIL.n89 B 2.19617f
C508 VTAIL.t10 B 0.281882f
C509 VTAIL.t0 B 0.281882f
C510 VTAIL.n90 B 2.48104f
C511 VTAIL.n91 B 2.19616f
C512 VTAIL.n92 B 0.030272f
C513 VTAIL.n93 B 0.023208f
C514 VTAIL.n94 B 0.012471f
C515 VTAIL.n95 B 0.029477f
C516 VTAIL.n96 B 0.012838f
C517 VTAIL.n97 B 0.023208f
C518 VTAIL.n98 B 0.012838f
C519 VTAIL.n99 B 0.012471f
C520 VTAIL.n100 B 0.029477f
C521 VTAIL.n101 B 0.029477f
C522 VTAIL.n102 B 0.013205f
C523 VTAIL.n103 B 0.023208f
C524 VTAIL.n104 B 0.012471f
C525 VTAIL.n105 B 0.029477f
C526 VTAIL.n106 B 0.013205f
C527 VTAIL.n107 B 0.023208f
C528 VTAIL.n108 B 0.012471f
C529 VTAIL.n109 B 0.029477f
C530 VTAIL.n110 B 0.013205f
C531 VTAIL.n111 B 0.023208f
C532 VTAIL.n112 B 0.012471f
C533 VTAIL.n113 B 0.029477f
C534 VTAIL.n114 B 0.013205f
C535 VTAIL.n115 B 0.023208f
C536 VTAIL.n116 B 0.012471f
C537 VTAIL.n117 B 0.029477f
C538 VTAIL.n118 B 0.013205f
C539 VTAIL.n119 B 1.54931f
C540 VTAIL.n120 B 0.012471f
C541 VTAIL.t2 B 0.048633f
C542 VTAIL.n121 B 0.153521f
C543 VTAIL.n122 B 0.017413f
C544 VTAIL.n123 B 0.022108f
C545 VTAIL.n124 B 0.029477f
C546 VTAIL.n125 B 0.013205f
C547 VTAIL.n126 B 0.012471f
C548 VTAIL.n127 B 0.023208f
C549 VTAIL.n128 B 0.023208f
C550 VTAIL.n129 B 0.012471f
C551 VTAIL.n130 B 0.013205f
C552 VTAIL.n131 B 0.029477f
C553 VTAIL.n132 B 0.029477f
C554 VTAIL.n133 B 0.013205f
C555 VTAIL.n134 B 0.012471f
C556 VTAIL.n135 B 0.023208f
C557 VTAIL.n136 B 0.023208f
C558 VTAIL.n137 B 0.012471f
C559 VTAIL.n138 B 0.013205f
C560 VTAIL.n139 B 0.029477f
C561 VTAIL.n140 B 0.029477f
C562 VTAIL.n141 B 0.013205f
C563 VTAIL.n142 B 0.012471f
C564 VTAIL.n143 B 0.023208f
C565 VTAIL.n144 B 0.023208f
C566 VTAIL.n145 B 0.012471f
C567 VTAIL.n146 B 0.013205f
C568 VTAIL.n147 B 0.029477f
C569 VTAIL.n148 B 0.029477f
C570 VTAIL.n149 B 0.013205f
C571 VTAIL.n150 B 0.012471f
C572 VTAIL.n151 B 0.023208f
C573 VTAIL.n152 B 0.023208f
C574 VTAIL.n153 B 0.012471f
C575 VTAIL.n154 B 0.013205f
C576 VTAIL.n155 B 0.029477f
C577 VTAIL.n156 B 0.029477f
C578 VTAIL.n157 B 0.013205f
C579 VTAIL.n158 B 0.012471f
C580 VTAIL.n159 B 0.023208f
C581 VTAIL.n160 B 0.023208f
C582 VTAIL.n161 B 0.012471f
C583 VTAIL.n162 B 0.013205f
C584 VTAIL.n163 B 0.029477f
C585 VTAIL.n164 B 0.029477f
C586 VTAIL.n165 B 0.013205f
C587 VTAIL.n166 B 0.012471f
C588 VTAIL.n167 B 0.023208f
C589 VTAIL.n168 B 0.023208f
C590 VTAIL.n169 B 0.012471f
C591 VTAIL.n170 B 0.013205f
C592 VTAIL.n171 B 0.029477f
C593 VTAIL.n172 B 0.059659f
C594 VTAIL.n173 B 0.013205f
C595 VTAIL.n174 B 0.012471f
C596 VTAIL.n175 B 0.053961f
C597 VTAIL.n176 B 0.032965f
C598 VTAIL.n177 B 0.38585f
C599 VTAIL.t9 B 0.281882f
C600 VTAIL.t7 B 0.281882f
C601 VTAIL.n178 B 2.48104f
C602 VTAIL.n179 B 0.594463f
C603 VTAIL.n180 B 0.030272f
C604 VTAIL.n181 B 0.023208f
C605 VTAIL.n182 B 0.012471f
C606 VTAIL.n183 B 0.029477f
C607 VTAIL.n184 B 0.012838f
C608 VTAIL.n185 B 0.023208f
C609 VTAIL.n186 B 0.012838f
C610 VTAIL.n187 B 0.012471f
C611 VTAIL.n188 B 0.029477f
C612 VTAIL.n189 B 0.029477f
C613 VTAIL.n190 B 0.013205f
C614 VTAIL.n191 B 0.023208f
C615 VTAIL.n192 B 0.012471f
C616 VTAIL.n193 B 0.029477f
C617 VTAIL.n194 B 0.013205f
C618 VTAIL.n195 B 0.023208f
C619 VTAIL.n196 B 0.012471f
C620 VTAIL.n197 B 0.029477f
C621 VTAIL.n198 B 0.013205f
C622 VTAIL.n199 B 0.023208f
C623 VTAIL.n200 B 0.012471f
C624 VTAIL.n201 B 0.029477f
C625 VTAIL.n202 B 0.013205f
C626 VTAIL.n203 B 0.023208f
C627 VTAIL.n204 B 0.012471f
C628 VTAIL.n205 B 0.029477f
C629 VTAIL.n206 B 0.013205f
C630 VTAIL.n207 B 1.54931f
C631 VTAIL.n208 B 0.012471f
C632 VTAIL.t8 B 0.048633f
C633 VTAIL.n209 B 0.153521f
C634 VTAIL.n210 B 0.017413f
C635 VTAIL.n211 B 0.022108f
C636 VTAIL.n212 B 0.029477f
C637 VTAIL.n213 B 0.013205f
C638 VTAIL.n214 B 0.012471f
C639 VTAIL.n215 B 0.023208f
C640 VTAIL.n216 B 0.023208f
C641 VTAIL.n217 B 0.012471f
C642 VTAIL.n218 B 0.013205f
C643 VTAIL.n219 B 0.029477f
C644 VTAIL.n220 B 0.029477f
C645 VTAIL.n221 B 0.013205f
C646 VTAIL.n222 B 0.012471f
C647 VTAIL.n223 B 0.023208f
C648 VTAIL.n224 B 0.023208f
C649 VTAIL.n225 B 0.012471f
C650 VTAIL.n226 B 0.013205f
C651 VTAIL.n227 B 0.029477f
C652 VTAIL.n228 B 0.029477f
C653 VTAIL.n229 B 0.013205f
C654 VTAIL.n230 B 0.012471f
C655 VTAIL.n231 B 0.023208f
C656 VTAIL.n232 B 0.023208f
C657 VTAIL.n233 B 0.012471f
C658 VTAIL.n234 B 0.013205f
C659 VTAIL.n235 B 0.029477f
C660 VTAIL.n236 B 0.029477f
C661 VTAIL.n237 B 0.013205f
C662 VTAIL.n238 B 0.012471f
C663 VTAIL.n239 B 0.023208f
C664 VTAIL.n240 B 0.023208f
C665 VTAIL.n241 B 0.012471f
C666 VTAIL.n242 B 0.013205f
C667 VTAIL.n243 B 0.029477f
C668 VTAIL.n244 B 0.029477f
C669 VTAIL.n245 B 0.013205f
C670 VTAIL.n246 B 0.012471f
C671 VTAIL.n247 B 0.023208f
C672 VTAIL.n248 B 0.023208f
C673 VTAIL.n249 B 0.012471f
C674 VTAIL.n250 B 0.013205f
C675 VTAIL.n251 B 0.029477f
C676 VTAIL.n252 B 0.029477f
C677 VTAIL.n253 B 0.013205f
C678 VTAIL.n254 B 0.012471f
C679 VTAIL.n255 B 0.023208f
C680 VTAIL.n256 B 0.023208f
C681 VTAIL.n257 B 0.012471f
C682 VTAIL.n258 B 0.013205f
C683 VTAIL.n259 B 0.029477f
C684 VTAIL.n260 B 0.059659f
C685 VTAIL.n261 B 0.013205f
C686 VTAIL.n262 B 0.012471f
C687 VTAIL.n263 B 0.053961f
C688 VTAIL.n264 B 0.032965f
C689 VTAIL.n265 B 1.76707f
C690 VTAIL.n266 B 0.030272f
C691 VTAIL.n267 B 0.023208f
C692 VTAIL.n268 B 0.012471f
C693 VTAIL.n269 B 0.029477f
C694 VTAIL.n270 B 0.012838f
C695 VTAIL.n271 B 0.023208f
C696 VTAIL.n272 B 0.013205f
C697 VTAIL.n273 B 0.029477f
C698 VTAIL.n274 B 0.013205f
C699 VTAIL.n275 B 0.023208f
C700 VTAIL.n276 B 0.012471f
C701 VTAIL.n277 B 0.029477f
C702 VTAIL.n278 B 0.013205f
C703 VTAIL.n279 B 0.023208f
C704 VTAIL.n280 B 0.012471f
C705 VTAIL.n281 B 0.029477f
C706 VTAIL.n282 B 0.013205f
C707 VTAIL.n283 B 0.023208f
C708 VTAIL.n284 B 0.012471f
C709 VTAIL.n285 B 0.029477f
C710 VTAIL.n286 B 0.013205f
C711 VTAIL.n287 B 0.023208f
C712 VTAIL.n288 B 0.012471f
C713 VTAIL.n289 B 0.029477f
C714 VTAIL.n290 B 0.013205f
C715 VTAIL.n291 B 1.54931f
C716 VTAIL.n292 B 0.012471f
C717 VTAIL.t3 B 0.048633f
C718 VTAIL.n293 B 0.153521f
C719 VTAIL.n294 B 0.017413f
C720 VTAIL.n295 B 0.022108f
C721 VTAIL.n296 B 0.029477f
C722 VTAIL.n297 B 0.013205f
C723 VTAIL.n298 B 0.012471f
C724 VTAIL.n299 B 0.023208f
C725 VTAIL.n300 B 0.023208f
C726 VTAIL.n301 B 0.012471f
C727 VTAIL.n302 B 0.013205f
C728 VTAIL.n303 B 0.029477f
C729 VTAIL.n304 B 0.029477f
C730 VTAIL.n305 B 0.013205f
C731 VTAIL.n306 B 0.012471f
C732 VTAIL.n307 B 0.023208f
C733 VTAIL.n308 B 0.023208f
C734 VTAIL.n309 B 0.012471f
C735 VTAIL.n310 B 0.013205f
C736 VTAIL.n311 B 0.029477f
C737 VTAIL.n312 B 0.029477f
C738 VTAIL.n313 B 0.013205f
C739 VTAIL.n314 B 0.012471f
C740 VTAIL.n315 B 0.023208f
C741 VTAIL.n316 B 0.023208f
C742 VTAIL.n317 B 0.012471f
C743 VTAIL.n318 B 0.013205f
C744 VTAIL.n319 B 0.029477f
C745 VTAIL.n320 B 0.029477f
C746 VTAIL.n321 B 0.013205f
C747 VTAIL.n322 B 0.012471f
C748 VTAIL.n323 B 0.023208f
C749 VTAIL.n324 B 0.023208f
C750 VTAIL.n325 B 0.012471f
C751 VTAIL.n326 B 0.013205f
C752 VTAIL.n327 B 0.029477f
C753 VTAIL.n328 B 0.029477f
C754 VTAIL.n329 B 0.013205f
C755 VTAIL.n330 B 0.012471f
C756 VTAIL.n331 B 0.023208f
C757 VTAIL.n332 B 0.023208f
C758 VTAIL.n333 B 0.012471f
C759 VTAIL.n334 B 0.012471f
C760 VTAIL.n335 B 0.013205f
C761 VTAIL.n336 B 0.029477f
C762 VTAIL.n337 B 0.029477f
C763 VTAIL.n338 B 0.029477f
C764 VTAIL.n339 B 0.012838f
C765 VTAIL.n340 B 0.012471f
C766 VTAIL.n341 B 0.023208f
C767 VTAIL.n342 B 0.023208f
C768 VTAIL.n343 B 0.012471f
C769 VTAIL.n344 B 0.013205f
C770 VTAIL.n345 B 0.029477f
C771 VTAIL.n346 B 0.059659f
C772 VTAIL.n347 B 0.013205f
C773 VTAIL.n348 B 0.012471f
C774 VTAIL.n349 B 0.053961f
C775 VTAIL.n350 B 0.032965f
C776 VTAIL.n351 B 1.7076f
C777 VP.t1 B 2.65831f
C778 VP.n0 B 1.00813f
C779 VP.n1 B 0.020415f
C780 VP.n2 B 0.027527f
C781 VP.n3 B 0.020415f
C782 VP.t5 B 2.65831f
C783 VP.n4 B 0.038049f
C784 VP.n5 B 0.020415f
C785 VP.n6 B 0.038049f
C786 VP.t2 B 2.65831f
C787 VP.n7 B 1.00813f
C788 VP.n8 B 0.020415f
C789 VP.n9 B 0.027527f
C790 VP.n10 B 0.232312f
C791 VP.t4 B 2.65831f
C792 VP.t3 B 2.89152f
C793 VP.n11 B 0.954857f
C794 VP.n12 B 1.00125f
C795 VP.n13 B 0.038049f
C796 VP.n14 B 0.038049f
C797 VP.n15 B 0.020415f
C798 VP.n16 B 0.020415f
C799 VP.n17 B 0.020415f
C800 VP.n18 B 0.032078f
C801 VP.n19 B 0.038049f
C802 VP.n20 B 0.035043f
C803 VP.n21 B 0.03295f
C804 VP.n22 B 1.26502f
C805 VP.n23 B 1.27879f
C806 VP.t0 B 2.65831f
C807 VP.n24 B 1.00813f
C808 VP.n25 B 0.035043f
C809 VP.n26 B 0.03295f
C810 VP.n27 B 0.020415f
C811 VP.n28 B 0.020415f
C812 VP.n29 B 0.032078f
C813 VP.n30 B 0.027527f
C814 VP.n31 B 0.038049f
C815 VP.n32 B 0.020415f
C816 VP.n33 B 0.020415f
C817 VP.n34 B 0.020415f
C818 VP.n35 B 0.943796f
C819 VP.n36 B 0.038049f
C820 VP.n37 B 0.038049f
C821 VP.n38 B 0.020415f
C822 VP.n39 B 0.020415f
C823 VP.n40 B 0.020415f
C824 VP.n41 B 0.032078f
C825 VP.n42 B 0.038049f
C826 VP.n43 B 0.035043f
C827 VP.n44 B 0.03295f
C828 VP.n45 B 0.042556f
.ends

