* NGSPICE file created from diff_pair_sample_0777.ext - technology: sky130A

.subckt diff_pair_sample_0777 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=3.042 ps=16.38 w=7.8 l=3.32
X1 VDD1.t5 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=3.042 ps=16.38 w=7.8 l=3.32
X2 VTAIL.t2 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=1.287 ps=8.13 w=7.8 l=3.32
X3 VDD1.t3 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=1.287 ps=8.13 w=7.8 l=3.32
X4 VTAIL.t4 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=1.287 ps=8.13 w=7.8 l=3.32
X5 VDD2.t4 VN.t1 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=1.287 ps=8.13 w=7.8 l=3.32
X6 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=0 ps=0 w=7.8 l=3.32
X7 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=3.042 ps=16.38 w=7.8 l=3.32
X8 VTAIL.t7 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=1.287 ps=8.13 w=7.8 l=3.32
X9 VDD2.t2 VN.t3 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=3.042 ps=16.38 w=7.8 l=3.32
X10 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=0 ps=0 w=7.8 l=3.32
X11 VTAIL.t11 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.287 pd=8.13 as=1.287 ps=8.13 w=7.8 l=3.32
X12 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=0 ps=0 w=7.8 l=3.32
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=0 ps=0 w=7.8 l=3.32
X14 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=1.287 ps=8.13 w=7.8 l=3.32
X15 VDD2.t0 VN.t5 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=3.042 pd=16.38 as=1.287 ps=8.13 w=7.8 l=3.32
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n23 VN.t3 89.4682
R15 VN.n5 VN.t5 89.4682
R16 VN.n17 VN.n0 82.588
R17 VN.n35 VN.n18 82.588
R18 VN.n4 VN.t2 56.621
R19 VN.n0 VN.t0 56.621
R20 VN.n22 VN.t4 56.621
R21 VN.n18 VN.t1 56.621
R22 VN.n9 VN.n2 56.4773
R23 VN.n27 VN.n20 56.4773
R24 VN.n5 VN.n4 49.9437
R25 VN.n23 VN.n22 49.9437
R26 VN VN.n35 48.4865
R27 VN.n7 VN.n4 24.3439
R28 VN.n8 VN.n7 24.3439
R29 VN.n9 VN.n8 24.3439
R30 VN.n13 VN.n2 24.3439
R31 VN.n14 VN.n13 24.3439
R32 VN.n15 VN.n14 24.3439
R33 VN.n27 VN.n26 24.3439
R34 VN.n26 VN.n25 24.3439
R35 VN.n25 VN.n22 24.3439
R36 VN.n33 VN.n32 24.3439
R37 VN.n32 VN.n31 24.3439
R38 VN.n31 VN.n20 24.3439
R39 VN.n15 VN.n0 7.30353
R40 VN.n33 VN.n18 7.30353
R41 VN.n24 VN.n23 3.25664
R42 VN.n6 VN.n5 3.25664
R43 VN.n35 VN.n34 0.355081
R44 VN.n17 VN.n16 0.355081
R45 VN VN.n17 0.26685
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VTAIL.n10 VTAIL.t5 50.6923
R59 VTAIL.n7 VTAIL.t10 50.6922
R60 VTAIL.n11 VTAIL.t6 50.6921
R61 VTAIL.n2 VTAIL.t1 50.6921
R62 VTAIL.n9 VTAIL.n8 48.1538
R63 VTAIL.n6 VTAIL.n5 48.1538
R64 VTAIL.n1 VTAIL.n0 48.1538
R65 VTAIL.n4 VTAIL.n3 48.1538
R66 VTAIL.n6 VTAIL.n4 25.3841
R67 VTAIL.n11 VTAIL.n10 22.2376
R68 VTAIL.n7 VTAIL.n6 3.14705
R69 VTAIL.n10 VTAIL.n9 3.14705
R70 VTAIL.n4 VTAIL.n2 3.14705
R71 VTAIL.n0 VTAIL.t8 2.53896
R72 VTAIL.n0 VTAIL.t7 2.53896
R73 VTAIL.n3 VTAIL.t0 2.53896
R74 VTAIL.n3 VTAIL.t2 2.53896
R75 VTAIL.n8 VTAIL.t3 2.53896
R76 VTAIL.n8 VTAIL.t4 2.53896
R77 VTAIL.n5 VTAIL.t9 2.53896
R78 VTAIL.n5 VTAIL.t11 2.53896
R79 VTAIL VTAIL.n11 2.30222
R80 VTAIL.n9 VTAIL.n7 2.0436
R81 VTAIL.n2 VTAIL.n1 2.0436
R82 VTAIL VTAIL.n1 0.845328
R83 VDD2.n1 VDD2.t0 69.6755
R84 VDD2.n2 VDD2.t4 67.371
R85 VDD2.n1 VDD2.n0 65.5639
R86 VDD2 VDD2.n3 65.5611
R87 VDD2.n2 VDD2.n1 40.6657
R88 VDD2.n3 VDD2.t1 2.53896
R89 VDD2.n3 VDD2.t2 2.53896
R90 VDD2.n0 VDD2.t3 2.53896
R91 VDD2.n0 VDD2.t5 2.53896
R92 VDD2 VDD2.n2 2.4186
R93 B.n758 B.n757 585
R94 B.n264 B.n128 585
R95 B.n263 B.n262 585
R96 B.n261 B.n260 585
R97 B.n259 B.n258 585
R98 B.n257 B.n256 585
R99 B.n255 B.n254 585
R100 B.n253 B.n252 585
R101 B.n251 B.n250 585
R102 B.n249 B.n248 585
R103 B.n247 B.n246 585
R104 B.n245 B.n244 585
R105 B.n243 B.n242 585
R106 B.n241 B.n240 585
R107 B.n239 B.n238 585
R108 B.n237 B.n236 585
R109 B.n235 B.n234 585
R110 B.n233 B.n232 585
R111 B.n231 B.n230 585
R112 B.n229 B.n228 585
R113 B.n227 B.n226 585
R114 B.n225 B.n224 585
R115 B.n223 B.n222 585
R116 B.n221 B.n220 585
R117 B.n219 B.n218 585
R118 B.n217 B.n216 585
R119 B.n215 B.n214 585
R120 B.n213 B.n212 585
R121 B.n211 B.n210 585
R122 B.n208 B.n207 585
R123 B.n206 B.n205 585
R124 B.n204 B.n203 585
R125 B.n202 B.n201 585
R126 B.n200 B.n199 585
R127 B.n198 B.n197 585
R128 B.n196 B.n195 585
R129 B.n194 B.n193 585
R130 B.n192 B.n191 585
R131 B.n190 B.n189 585
R132 B.n187 B.n186 585
R133 B.n185 B.n184 585
R134 B.n183 B.n182 585
R135 B.n181 B.n180 585
R136 B.n179 B.n178 585
R137 B.n177 B.n176 585
R138 B.n175 B.n174 585
R139 B.n173 B.n172 585
R140 B.n171 B.n170 585
R141 B.n169 B.n168 585
R142 B.n167 B.n166 585
R143 B.n165 B.n164 585
R144 B.n163 B.n162 585
R145 B.n161 B.n160 585
R146 B.n159 B.n158 585
R147 B.n157 B.n156 585
R148 B.n155 B.n154 585
R149 B.n153 B.n152 585
R150 B.n151 B.n150 585
R151 B.n149 B.n148 585
R152 B.n147 B.n146 585
R153 B.n145 B.n144 585
R154 B.n143 B.n142 585
R155 B.n141 B.n140 585
R156 B.n139 B.n138 585
R157 B.n137 B.n136 585
R158 B.n135 B.n134 585
R159 B.n95 B.n94 585
R160 B.n763 B.n762 585
R161 B.n756 B.n129 585
R162 B.n129 B.n92 585
R163 B.n755 B.n91 585
R164 B.n767 B.n91 585
R165 B.n754 B.n90 585
R166 B.n768 B.n90 585
R167 B.n753 B.n89 585
R168 B.n769 B.n89 585
R169 B.n752 B.n751 585
R170 B.n751 B.n85 585
R171 B.n750 B.n84 585
R172 B.n775 B.n84 585
R173 B.n749 B.n83 585
R174 B.n776 B.n83 585
R175 B.n748 B.n82 585
R176 B.n777 B.n82 585
R177 B.n747 B.n746 585
R178 B.n746 B.n81 585
R179 B.n745 B.n77 585
R180 B.n783 B.n77 585
R181 B.n744 B.n76 585
R182 B.n784 B.n76 585
R183 B.n743 B.n75 585
R184 B.n785 B.n75 585
R185 B.n742 B.n741 585
R186 B.n741 B.n71 585
R187 B.n740 B.n70 585
R188 B.n791 B.n70 585
R189 B.n739 B.n69 585
R190 B.n792 B.n69 585
R191 B.n738 B.n68 585
R192 B.n793 B.n68 585
R193 B.n737 B.n736 585
R194 B.n736 B.n64 585
R195 B.n735 B.n63 585
R196 B.n799 B.n63 585
R197 B.n734 B.n62 585
R198 B.n800 B.n62 585
R199 B.n733 B.n61 585
R200 B.n801 B.n61 585
R201 B.n732 B.n731 585
R202 B.n731 B.n57 585
R203 B.n730 B.n56 585
R204 B.n807 B.n56 585
R205 B.n729 B.n55 585
R206 B.n808 B.n55 585
R207 B.n728 B.n54 585
R208 B.n809 B.n54 585
R209 B.n727 B.n726 585
R210 B.n726 B.n50 585
R211 B.n725 B.n49 585
R212 B.n815 B.n49 585
R213 B.n724 B.n48 585
R214 B.n816 B.n48 585
R215 B.n723 B.n47 585
R216 B.n817 B.n47 585
R217 B.n722 B.n721 585
R218 B.n721 B.n43 585
R219 B.n720 B.n42 585
R220 B.n823 B.n42 585
R221 B.n719 B.n41 585
R222 B.n824 B.n41 585
R223 B.n718 B.n40 585
R224 B.n825 B.n40 585
R225 B.n717 B.n716 585
R226 B.n716 B.n36 585
R227 B.n715 B.n35 585
R228 B.n831 B.n35 585
R229 B.n714 B.n34 585
R230 B.n832 B.n34 585
R231 B.n713 B.n33 585
R232 B.n833 B.n33 585
R233 B.n712 B.n711 585
R234 B.n711 B.n29 585
R235 B.n710 B.n28 585
R236 B.n839 B.n28 585
R237 B.n709 B.n27 585
R238 B.n840 B.n27 585
R239 B.n708 B.n26 585
R240 B.n841 B.n26 585
R241 B.n707 B.n706 585
R242 B.n706 B.n22 585
R243 B.n705 B.n21 585
R244 B.n847 B.n21 585
R245 B.n704 B.n20 585
R246 B.n848 B.n20 585
R247 B.n703 B.n19 585
R248 B.n849 B.n19 585
R249 B.n702 B.n701 585
R250 B.n701 B.n18 585
R251 B.n700 B.n14 585
R252 B.n855 B.n14 585
R253 B.n699 B.n13 585
R254 B.n856 B.n13 585
R255 B.n698 B.n12 585
R256 B.n857 B.n12 585
R257 B.n697 B.n696 585
R258 B.n696 B.n8 585
R259 B.n695 B.n7 585
R260 B.n863 B.n7 585
R261 B.n694 B.n6 585
R262 B.n864 B.n6 585
R263 B.n693 B.n5 585
R264 B.n865 B.n5 585
R265 B.n692 B.n691 585
R266 B.n691 B.n4 585
R267 B.n690 B.n265 585
R268 B.n690 B.n689 585
R269 B.n680 B.n266 585
R270 B.n267 B.n266 585
R271 B.n682 B.n681 585
R272 B.n683 B.n682 585
R273 B.n679 B.n272 585
R274 B.n272 B.n271 585
R275 B.n678 B.n677 585
R276 B.n677 B.n676 585
R277 B.n274 B.n273 585
R278 B.n669 B.n274 585
R279 B.n668 B.n667 585
R280 B.n670 B.n668 585
R281 B.n666 B.n279 585
R282 B.n279 B.n278 585
R283 B.n665 B.n664 585
R284 B.n664 B.n663 585
R285 B.n281 B.n280 585
R286 B.n282 B.n281 585
R287 B.n656 B.n655 585
R288 B.n657 B.n656 585
R289 B.n654 B.n287 585
R290 B.n287 B.n286 585
R291 B.n653 B.n652 585
R292 B.n652 B.n651 585
R293 B.n289 B.n288 585
R294 B.n290 B.n289 585
R295 B.n644 B.n643 585
R296 B.n645 B.n644 585
R297 B.n642 B.n295 585
R298 B.n295 B.n294 585
R299 B.n641 B.n640 585
R300 B.n640 B.n639 585
R301 B.n297 B.n296 585
R302 B.n298 B.n297 585
R303 B.n632 B.n631 585
R304 B.n633 B.n632 585
R305 B.n630 B.n303 585
R306 B.n303 B.n302 585
R307 B.n629 B.n628 585
R308 B.n628 B.n627 585
R309 B.n305 B.n304 585
R310 B.n306 B.n305 585
R311 B.n620 B.n619 585
R312 B.n621 B.n620 585
R313 B.n618 B.n311 585
R314 B.n311 B.n310 585
R315 B.n617 B.n616 585
R316 B.n616 B.n615 585
R317 B.n313 B.n312 585
R318 B.n314 B.n313 585
R319 B.n608 B.n607 585
R320 B.n609 B.n608 585
R321 B.n606 B.n318 585
R322 B.n322 B.n318 585
R323 B.n605 B.n604 585
R324 B.n604 B.n603 585
R325 B.n320 B.n319 585
R326 B.n321 B.n320 585
R327 B.n596 B.n595 585
R328 B.n597 B.n596 585
R329 B.n594 B.n327 585
R330 B.n327 B.n326 585
R331 B.n593 B.n592 585
R332 B.n592 B.n591 585
R333 B.n329 B.n328 585
R334 B.n330 B.n329 585
R335 B.n584 B.n583 585
R336 B.n585 B.n584 585
R337 B.n582 B.n335 585
R338 B.n335 B.n334 585
R339 B.n581 B.n580 585
R340 B.n580 B.n579 585
R341 B.n337 B.n336 585
R342 B.n338 B.n337 585
R343 B.n572 B.n571 585
R344 B.n573 B.n572 585
R345 B.n570 B.n343 585
R346 B.n343 B.n342 585
R347 B.n569 B.n568 585
R348 B.n568 B.n567 585
R349 B.n345 B.n344 585
R350 B.n560 B.n345 585
R351 B.n559 B.n558 585
R352 B.n561 B.n559 585
R353 B.n557 B.n350 585
R354 B.n350 B.n349 585
R355 B.n556 B.n555 585
R356 B.n555 B.n554 585
R357 B.n352 B.n351 585
R358 B.n353 B.n352 585
R359 B.n547 B.n546 585
R360 B.n548 B.n547 585
R361 B.n545 B.n358 585
R362 B.n358 B.n357 585
R363 B.n544 B.n543 585
R364 B.n543 B.n542 585
R365 B.n360 B.n359 585
R366 B.n361 B.n360 585
R367 B.n538 B.n537 585
R368 B.n364 B.n363 585
R369 B.n534 B.n533 585
R370 B.n535 B.n534 585
R371 B.n532 B.n398 585
R372 B.n531 B.n530 585
R373 B.n529 B.n528 585
R374 B.n527 B.n526 585
R375 B.n525 B.n524 585
R376 B.n523 B.n522 585
R377 B.n521 B.n520 585
R378 B.n519 B.n518 585
R379 B.n517 B.n516 585
R380 B.n515 B.n514 585
R381 B.n513 B.n512 585
R382 B.n511 B.n510 585
R383 B.n509 B.n508 585
R384 B.n507 B.n506 585
R385 B.n505 B.n504 585
R386 B.n503 B.n502 585
R387 B.n501 B.n500 585
R388 B.n499 B.n498 585
R389 B.n497 B.n496 585
R390 B.n495 B.n494 585
R391 B.n493 B.n492 585
R392 B.n491 B.n490 585
R393 B.n489 B.n488 585
R394 B.n487 B.n486 585
R395 B.n485 B.n484 585
R396 B.n483 B.n482 585
R397 B.n481 B.n480 585
R398 B.n479 B.n478 585
R399 B.n477 B.n476 585
R400 B.n475 B.n474 585
R401 B.n473 B.n472 585
R402 B.n471 B.n470 585
R403 B.n469 B.n468 585
R404 B.n467 B.n466 585
R405 B.n465 B.n464 585
R406 B.n463 B.n462 585
R407 B.n461 B.n460 585
R408 B.n459 B.n458 585
R409 B.n457 B.n456 585
R410 B.n455 B.n454 585
R411 B.n453 B.n452 585
R412 B.n451 B.n450 585
R413 B.n449 B.n448 585
R414 B.n447 B.n446 585
R415 B.n445 B.n444 585
R416 B.n443 B.n442 585
R417 B.n441 B.n440 585
R418 B.n439 B.n438 585
R419 B.n437 B.n436 585
R420 B.n435 B.n434 585
R421 B.n433 B.n432 585
R422 B.n431 B.n430 585
R423 B.n429 B.n428 585
R424 B.n427 B.n426 585
R425 B.n425 B.n424 585
R426 B.n423 B.n422 585
R427 B.n421 B.n420 585
R428 B.n419 B.n418 585
R429 B.n417 B.n416 585
R430 B.n415 B.n414 585
R431 B.n413 B.n412 585
R432 B.n411 B.n410 585
R433 B.n409 B.n408 585
R434 B.n407 B.n406 585
R435 B.n405 B.n397 585
R436 B.n535 B.n397 585
R437 B.n539 B.n362 585
R438 B.n362 B.n361 585
R439 B.n541 B.n540 585
R440 B.n542 B.n541 585
R441 B.n356 B.n355 585
R442 B.n357 B.n356 585
R443 B.n550 B.n549 585
R444 B.n549 B.n548 585
R445 B.n551 B.n354 585
R446 B.n354 B.n353 585
R447 B.n553 B.n552 585
R448 B.n554 B.n553 585
R449 B.n348 B.n347 585
R450 B.n349 B.n348 585
R451 B.n563 B.n562 585
R452 B.n562 B.n561 585
R453 B.n564 B.n346 585
R454 B.n560 B.n346 585
R455 B.n566 B.n565 585
R456 B.n567 B.n566 585
R457 B.n341 B.n340 585
R458 B.n342 B.n341 585
R459 B.n575 B.n574 585
R460 B.n574 B.n573 585
R461 B.n576 B.n339 585
R462 B.n339 B.n338 585
R463 B.n578 B.n577 585
R464 B.n579 B.n578 585
R465 B.n333 B.n332 585
R466 B.n334 B.n333 585
R467 B.n587 B.n586 585
R468 B.n586 B.n585 585
R469 B.n588 B.n331 585
R470 B.n331 B.n330 585
R471 B.n590 B.n589 585
R472 B.n591 B.n590 585
R473 B.n325 B.n324 585
R474 B.n326 B.n325 585
R475 B.n599 B.n598 585
R476 B.n598 B.n597 585
R477 B.n600 B.n323 585
R478 B.n323 B.n321 585
R479 B.n602 B.n601 585
R480 B.n603 B.n602 585
R481 B.n317 B.n316 585
R482 B.n322 B.n317 585
R483 B.n611 B.n610 585
R484 B.n610 B.n609 585
R485 B.n612 B.n315 585
R486 B.n315 B.n314 585
R487 B.n614 B.n613 585
R488 B.n615 B.n614 585
R489 B.n309 B.n308 585
R490 B.n310 B.n309 585
R491 B.n623 B.n622 585
R492 B.n622 B.n621 585
R493 B.n624 B.n307 585
R494 B.n307 B.n306 585
R495 B.n626 B.n625 585
R496 B.n627 B.n626 585
R497 B.n301 B.n300 585
R498 B.n302 B.n301 585
R499 B.n635 B.n634 585
R500 B.n634 B.n633 585
R501 B.n636 B.n299 585
R502 B.n299 B.n298 585
R503 B.n638 B.n637 585
R504 B.n639 B.n638 585
R505 B.n293 B.n292 585
R506 B.n294 B.n293 585
R507 B.n647 B.n646 585
R508 B.n646 B.n645 585
R509 B.n648 B.n291 585
R510 B.n291 B.n290 585
R511 B.n650 B.n649 585
R512 B.n651 B.n650 585
R513 B.n285 B.n284 585
R514 B.n286 B.n285 585
R515 B.n659 B.n658 585
R516 B.n658 B.n657 585
R517 B.n660 B.n283 585
R518 B.n283 B.n282 585
R519 B.n662 B.n661 585
R520 B.n663 B.n662 585
R521 B.n277 B.n276 585
R522 B.n278 B.n277 585
R523 B.n672 B.n671 585
R524 B.n671 B.n670 585
R525 B.n673 B.n275 585
R526 B.n669 B.n275 585
R527 B.n675 B.n674 585
R528 B.n676 B.n675 585
R529 B.n270 B.n269 585
R530 B.n271 B.n270 585
R531 B.n685 B.n684 585
R532 B.n684 B.n683 585
R533 B.n686 B.n268 585
R534 B.n268 B.n267 585
R535 B.n688 B.n687 585
R536 B.n689 B.n688 585
R537 B.n2 B.n0 585
R538 B.n4 B.n2 585
R539 B.n3 B.n1 585
R540 B.n864 B.n3 585
R541 B.n862 B.n861 585
R542 B.n863 B.n862 585
R543 B.n860 B.n9 585
R544 B.n9 B.n8 585
R545 B.n859 B.n858 585
R546 B.n858 B.n857 585
R547 B.n11 B.n10 585
R548 B.n856 B.n11 585
R549 B.n854 B.n853 585
R550 B.n855 B.n854 585
R551 B.n852 B.n15 585
R552 B.n18 B.n15 585
R553 B.n851 B.n850 585
R554 B.n850 B.n849 585
R555 B.n17 B.n16 585
R556 B.n848 B.n17 585
R557 B.n846 B.n845 585
R558 B.n847 B.n846 585
R559 B.n844 B.n23 585
R560 B.n23 B.n22 585
R561 B.n843 B.n842 585
R562 B.n842 B.n841 585
R563 B.n25 B.n24 585
R564 B.n840 B.n25 585
R565 B.n838 B.n837 585
R566 B.n839 B.n838 585
R567 B.n836 B.n30 585
R568 B.n30 B.n29 585
R569 B.n835 B.n834 585
R570 B.n834 B.n833 585
R571 B.n32 B.n31 585
R572 B.n832 B.n32 585
R573 B.n830 B.n829 585
R574 B.n831 B.n830 585
R575 B.n828 B.n37 585
R576 B.n37 B.n36 585
R577 B.n827 B.n826 585
R578 B.n826 B.n825 585
R579 B.n39 B.n38 585
R580 B.n824 B.n39 585
R581 B.n822 B.n821 585
R582 B.n823 B.n822 585
R583 B.n820 B.n44 585
R584 B.n44 B.n43 585
R585 B.n819 B.n818 585
R586 B.n818 B.n817 585
R587 B.n46 B.n45 585
R588 B.n816 B.n46 585
R589 B.n814 B.n813 585
R590 B.n815 B.n814 585
R591 B.n812 B.n51 585
R592 B.n51 B.n50 585
R593 B.n811 B.n810 585
R594 B.n810 B.n809 585
R595 B.n53 B.n52 585
R596 B.n808 B.n53 585
R597 B.n806 B.n805 585
R598 B.n807 B.n806 585
R599 B.n804 B.n58 585
R600 B.n58 B.n57 585
R601 B.n803 B.n802 585
R602 B.n802 B.n801 585
R603 B.n60 B.n59 585
R604 B.n800 B.n60 585
R605 B.n798 B.n797 585
R606 B.n799 B.n798 585
R607 B.n796 B.n65 585
R608 B.n65 B.n64 585
R609 B.n795 B.n794 585
R610 B.n794 B.n793 585
R611 B.n67 B.n66 585
R612 B.n792 B.n67 585
R613 B.n790 B.n789 585
R614 B.n791 B.n790 585
R615 B.n788 B.n72 585
R616 B.n72 B.n71 585
R617 B.n787 B.n786 585
R618 B.n786 B.n785 585
R619 B.n74 B.n73 585
R620 B.n784 B.n74 585
R621 B.n782 B.n781 585
R622 B.n783 B.n782 585
R623 B.n780 B.n78 585
R624 B.n81 B.n78 585
R625 B.n779 B.n778 585
R626 B.n778 B.n777 585
R627 B.n80 B.n79 585
R628 B.n776 B.n80 585
R629 B.n774 B.n773 585
R630 B.n775 B.n774 585
R631 B.n772 B.n86 585
R632 B.n86 B.n85 585
R633 B.n771 B.n770 585
R634 B.n770 B.n769 585
R635 B.n88 B.n87 585
R636 B.n768 B.n88 585
R637 B.n766 B.n765 585
R638 B.n767 B.n766 585
R639 B.n764 B.n93 585
R640 B.n93 B.n92 585
R641 B.n867 B.n866 585
R642 B.n866 B.n865 585
R643 B.n537 B.n362 516.524
R644 B.n762 B.n93 516.524
R645 B.n397 B.n360 516.524
R646 B.n758 B.n129 516.524
R647 B.n402 B.t17 265.546
R648 B.n399 B.t13 265.546
R649 B.n132 B.t10 265.546
R650 B.n130 B.t6 265.546
R651 B.n760 B.n759 256.663
R652 B.n760 B.n127 256.663
R653 B.n760 B.n126 256.663
R654 B.n760 B.n125 256.663
R655 B.n760 B.n124 256.663
R656 B.n760 B.n123 256.663
R657 B.n760 B.n122 256.663
R658 B.n760 B.n121 256.663
R659 B.n760 B.n120 256.663
R660 B.n760 B.n119 256.663
R661 B.n760 B.n118 256.663
R662 B.n760 B.n117 256.663
R663 B.n760 B.n116 256.663
R664 B.n760 B.n115 256.663
R665 B.n760 B.n114 256.663
R666 B.n760 B.n113 256.663
R667 B.n760 B.n112 256.663
R668 B.n760 B.n111 256.663
R669 B.n760 B.n110 256.663
R670 B.n760 B.n109 256.663
R671 B.n760 B.n108 256.663
R672 B.n760 B.n107 256.663
R673 B.n760 B.n106 256.663
R674 B.n760 B.n105 256.663
R675 B.n760 B.n104 256.663
R676 B.n760 B.n103 256.663
R677 B.n760 B.n102 256.663
R678 B.n760 B.n101 256.663
R679 B.n760 B.n100 256.663
R680 B.n760 B.n99 256.663
R681 B.n760 B.n98 256.663
R682 B.n760 B.n97 256.663
R683 B.n760 B.n96 256.663
R684 B.n761 B.n760 256.663
R685 B.n536 B.n535 256.663
R686 B.n535 B.n365 256.663
R687 B.n535 B.n366 256.663
R688 B.n535 B.n367 256.663
R689 B.n535 B.n368 256.663
R690 B.n535 B.n369 256.663
R691 B.n535 B.n370 256.663
R692 B.n535 B.n371 256.663
R693 B.n535 B.n372 256.663
R694 B.n535 B.n373 256.663
R695 B.n535 B.n374 256.663
R696 B.n535 B.n375 256.663
R697 B.n535 B.n376 256.663
R698 B.n535 B.n377 256.663
R699 B.n535 B.n378 256.663
R700 B.n535 B.n379 256.663
R701 B.n535 B.n380 256.663
R702 B.n535 B.n381 256.663
R703 B.n535 B.n382 256.663
R704 B.n535 B.n383 256.663
R705 B.n535 B.n384 256.663
R706 B.n535 B.n385 256.663
R707 B.n535 B.n386 256.663
R708 B.n535 B.n387 256.663
R709 B.n535 B.n388 256.663
R710 B.n535 B.n389 256.663
R711 B.n535 B.n390 256.663
R712 B.n535 B.n391 256.663
R713 B.n535 B.n392 256.663
R714 B.n535 B.n393 256.663
R715 B.n535 B.n394 256.663
R716 B.n535 B.n395 256.663
R717 B.n535 B.n396 256.663
R718 B.n541 B.n362 163.367
R719 B.n541 B.n356 163.367
R720 B.n549 B.n356 163.367
R721 B.n549 B.n354 163.367
R722 B.n553 B.n354 163.367
R723 B.n553 B.n348 163.367
R724 B.n562 B.n348 163.367
R725 B.n562 B.n346 163.367
R726 B.n566 B.n346 163.367
R727 B.n566 B.n341 163.367
R728 B.n574 B.n341 163.367
R729 B.n574 B.n339 163.367
R730 B.n578 B.n339 163.367
R731 B.n578 B.n333 163.367
R732 B.n586 B.n333 163.367
R733 B.n586 B.n331 163.367
R734 B.n590 B.n331 163.367
R735 B.n590 B.n325 163.367
R736 B.n598 B.n325 163.367
R737 B.n598 B.n323 163.367
R738 B.n602 B.n323 163.367
R739 B.n602 B.n317 163.367
R740 B.n610 B.n317 163.367
R741 B.n610 B.n315 163.367
R742 B.n614 B.n315 163.367
R743 B.n614 B.n309 163.367
R744 B.n622 B.n309 163.367
R745 B.n622 B.n307 163.367
R746 B.n626 B.n307 163.367
R747 B.n626 B.n301 163.367
R748 B.n634 B.n301 163.367
R749 B.n634 B.n299 163.367
R750 B.n638 B.n299 163.367
R751 B.n638 B.n293 163.367
R752 B.n646 B.n293 163.367
R753 B.n646 B.n291 163.367
R754 B.n650 B.n291 163.367
R755 B.n650 B.n285 163.367
R756 B.n658 B.n285 163.367
R757 B.n658 B.n283 163.367
R758 B.n662 B.n283 163.367
R759 B.n662 B.n277 163.367
R760 B.n671 B.n277 163.367
R761 B.n671 B.n275 163.367
R762 B.n675 B.n275 163.367
R763 B.n675 B.n270 163.367
R764 B.n684 B.n270 163.367
R765 B.n684 B.n268 163.367
R766 B.n688 B.n268 163.367
R767 B.n688 B.n2 163.367
R768 B.n866 B.n2 163.367
R769 B.n866 B.n3 163.367
R770 B.n862 B.n3 163.367
R771 B.n862 B.n9 163.367
R772 B.n858 B.n9 163.367
R773 B.n858 B.n11 163.367
R774 B.n854 B.n11 163.367
R775 B.n854 B.n15 163.367
R776 B.n850 B.n15 163.367
R777 B.n850 B.n17 163.367
R778 B.n846 B.n17 163.367
R779 B.n846 B.n23 163.367
R780 B.n842 B.n23 163.367
R781 B.n842 B.n25 163.367
R782 B.n838 B.n25 163.367
R783 B.n838 B.n30 163.367
R784 B.n834 B.n30 163.367
R785 B.n834 B.n32 163.367
R786 B.n830 B.n32 163.367
R787 B.n830 B.n37 163.367
R788 B.n826 B.n37 163.367
R789 B.n826 B.n39 163.367
R790 B.n822 B.n39 163.367
R791 B.n822 B.n44 163.367
R792 B.n818 B.n44 163.367
R793 B.n818 B.n46 163.367
R794 B.n814 B.n46 163.367
R795 B.n814 B.n51 163.367
R796 B.n810 B.n51 163.367
R797 B.n810 B.n53 163.367
R798 B.n806 B.n53 163.367
R799 B.n806 B.n58 163.367
R800 B.n802 B.n58 163.367
R801 B.n802 B.n60 163.367
R802 B.n798 B.n60 163.367
R803 B.n798 B.n65 163.367
R804 B.n794 B.n65 163.367
R805 B.n794 B.n67 163.367
R806 B.n790 B.n67 163.367
R807 B.n790 B.n72 163.367
R808 B.n786 B.n72 163.367
R809 B.n786 B.n74 163.367
R810 B.n782 B.n74 163.367
R811 B.n782 B.n78 163.367
R812 B.n778 B.n78 163.367
R813 B.n778 B.n80 163.367
R814 B.n774 B.n80 163.367
R815 B.n774 B.n86 163.367
R816 B.n770 B.n86 163.367
R817 B.n770 B.n88 163.367
R818 B.n766 B.n88 163.367
R819 B.n766 B.n93 163.367
R820 B.n534 B.n364 163.367
R821 B.n534 B.n398 163.367
R822 B.n530 B.n529 163.367
R823 B.n526 B.n525 163.367
R824 B.n522 B.n521 163.367
R825 B.n518 B.n517 163.367
R826 B.n514 B.n513 163.367
R827 B.n510 B.n509 163.367
R828 B.n506 B.n505 163.367
R829 B.n502 B.n501 163.367
R830 B.n498 B.n497 163.367
R831 B.n494 B.n493 163.367
R832 B.n490 B.n489 163.367
R833 B.n486 B.n485 163.367
R834 B.n482 B.n481 163.367
R835 B.n478 B.n477 163.367
R836 B.n474 B.n473 163.367
R837 B.n470 B.n469 163.367
R838 B.n466 B.n465 163.367
R839 B.n462 B.n461 163.367
R840 B.n458 B.n457 163.367
R841 B.n454 B.n453 163.367
R842 B.n450 B.n449 163.367
R843 B.n446 B.n445 163.367
R844 B.n442 B.n441 163.367
R845 B.n438 B.n437 163.367
R846 B.n434 B.n433 163.367
R847 B.n430 B.n429 163.367
R848 B.n426 B.n425 163.367
R849 B.n422 B.n421 163.367
R850 B.n418 B.n417 163.367
R851 B.n414 B.n413 163.367
R852 B.n410 B.n409 163.367
R853 B.n406 B.n397 163.367
R854 B.n543 B.n360 163.367
R855 B.n543 B.n358 163.367
R856 B.n547 B.n358 163.367
R857 B.n547 B.n352 163.367
R858 B.n555 B.n352 163.367
R859 B.n555 B.n350 163.367
R860 B.n559 B.n350 163.367
R861 B.n559 B.n345 163.367
R862 B.n568 B.n345 163.367
R863 B.n568 B.n343 163.367
R864 B.n572 B.n343 163.367
R865 B.n572 B.n337 163.367
R866 B.n580 B.n337 163.367
R867 B.n580 B.n335 163.367
R868 B.n584 B.n335 163.367
R869 B.n584 B.n329 163.367
R870 B.n592 B.n329 163.367
R871 B.n592 B.n327 163.367
R872 B.n596 B.n327 163.367
R873 B.n596 B.n320 163.367
R874 B.n604 B.n320 163.367
R875 B.n604 B.n318 163.367
R876 B.n608 B.n318 163.367
R877 B.n608 B.n313 163.367
R878 B.n616 B.n313 163.367
R879 B.n616 B.n311 163.367
R880 B.n620 B.n311 163.367
R881 B.n620 B.n305 163.367
R882 B.n628 B.n305 163.367
R883 B.n628 B.n303 163.367
R884 B.n632 B.n303 163.367
R885 B.n632 B.n297 163.367
R886 B.n640 B.n297 163.367
R887 B.n640 B.n295 163.367
R888 B.n644 B.n295 163.367
R889 B.n644 B.n289 163.367
R890 B.n652 B.n289 163.367
R891 B.n652 B.n287 163.367
R892 B.n656 B.n287 163.367
R893 B.n656 B.n281 163.367
R894 B.n664 B.n281 163.367
R895 B.n664 B.n279 163.367
R896 B.n668 B.n279 163.367
R897 B.n668 B.n274 163.367
R898 B.n677 B.n274 163.367
R899 B.n677 B.n272 163.367
R900 B.n682 B.n272 163.367
R901 B.n682 B.n266 163.367
R902 B.n690 B.n266 163.367
R903 B.n691 B.n690 163.367
R904 B.n691 B.n5 163.367
R905 B.n6 B.n5 163.367
R906 B.n7 B.n6 163.367
R907 B.n696 B.n7 163.367
R908 B.n696 B.n12 163.367
R909 B.n13 B.n12 163.367
R910 B.n14 B.n13 163.367
R911 B.n701 B.n14 163.367
R912 B.n701 B.n19 163.367
R913 B.n20 B.n19 163.367
R914 B.n21 B.n20 163.367
R915 B.n706 B.n21 163.367
R916 B.n706 B.n26 163.367
R917 B.n27 B.n26 163.367
R918 B.n28 B.n27 163.367
R919 B.n711 B.n28 163.367
R920 B.n711 B.n33 163.367
R921 B.n34 B.n33 163.367
R922 B.n35 B.n34 163.367
R923 B.n716 B.n35 163.367
R924 B.n716 B.n40 163.367
R925 B.n41 B.n40 163.367
R926 B.n42 B.n41 163.367
R927 B.n721 B.n42 163.367
R928 B.n721 B.n47 163.367
R929 B.n48 B.n47 163.367
R930 B.n49 B.n48 163.367
R931 B.n726 B.n49 163.367
R932 B.n726 B.n54 163.367
R933 B.n55 B.n54 163.367
R934 B.n56 B.n55 163.367
R935 B.n731 B.n56 163.367
R936 B.n731 B.n61 163.367
R937 B.n62 B.n61 163.367
R938 B.n63 B.n62 163.367
R939 B.n736 B.n63 163.367
R940 B.n736 B.n68 163.367
R941 B.n69 B.n68 163.367
R942 B.n70 B.n69 163.367
R943 B.n741 B.n70 163.367
R944 B.n741 B.n75 163.367
R945 B.n76 B.n75 163.367
R946 B.n77 B.n76 163.367
R947 B.n746 B.n77 163.367
R948 B.n746 B.n82 163.367
R949 B.n83 B.n82 163.367
R950 B.n84 B.n83 163.367
R951 B.n751 B.n84 163.367
R952 B.n751 B.n89 163.367
R953 B.n90 B.n89 163.367
R954 B.n91 B.n90 163.367
R955 B.n129 B.n91 163.367
R956 B.n134 B.n95 163.367
R957 B.n138 B.n137 163.367
R958 B.n142 B.n141 163.367
R959 B.n146 B.n145 163.367
R960 B.n150 B.n149 163.367
R961 B.n154 B.n153 163.367
R962 B.n158 B.n157 163.367
R963 B.n162 B.n161 163.367
R964 B.n166 B.n165 163.367
R965 B.n170 B.n169 163.367
R966 B.n174 B.n173 163.367
R967 B.n178 B.n177 163.367
R968 B.n182 B.n181 163.367
R969 B.n186 B.n185 163.367
R970 B.n191 B.n190 163.367
R971 B.n195 B.n194 163.367
R972 B.n199 B.n198 163.367
R973 B.n203 B.n202 163.367
R974 B.n207 B.n206 163.367
R975 B.n212 B.n211 163.367
R976 B.n216 B.n215 163.367
R977 B.n220 B.n219 163.367
R978 B.n224 B.n223 163.367
R979 B.n228 B.n227 163.367
R980 B.n232 B.n231 163.367
R981 B.n236 B.n235 163.367
R982 B.n240 B.n239 163.367
R983 B.n244 B.n243 163.367
R984 B.n248 B.n247 163.367
R985 B.n252 B.n251 163.367
R986 B.n256 B.n255 163.367
R987 B.n260 B.n259 163.367
R988 B.n262 B.n128 163.367
R989 B.n402 B.t19 145.667
R990 B.n130 B.t8 145.667
R991 B.n399 B.t16 145.659
R992 B.n132 B.t11 145.659
R993 B.n535 B.n361 106.846
R994 B.n760 B.n92 106.846
R995 B.n403 B.t18 74.8793
R996 B.n131 B.t9 74.8793
R997 B.n400 B.t15 74.8706
R998 B.n133 B.t12 74.8706
R999 B.n537 B.n536 71.676
R1000 B.n398 B.n365 71.676
R1001 B.n529 B.n366 71.676
R1002 B.n525 B.n367 71.676
R1003 B.n521 B.n368 71.676
R1004 B.n517 B.n369 71.676
R1005 B.n513 B.n370 71.676
R1006 B.n509 B.n371 71.676
R1007 B.n505 B.n372 71.676
R1008 B.n501 B.n373 71.676
R1009 B.n497 B.n374 71.676
R1010 B.n493 B.n375 71.676
R1011 B.n489 B.n376 71.676
R1012 B.n485 B.n377 71.676
R1013 B.n481 B.n378 71.676
R1014 B.n477 B.n379 71.676
R1015 B.n473 B.n380 71.676
R1016 B.n469 B.n381 71.676
R1017 B.n465 B.n382 71.676
R1018 B.n461 B.n383 71.676
R1019 B.n457 B.n384 71.676
R1020 B.n453 B.n385 71.676
R1021 B.n449 B.n386 71.676
R1022 B.n445 B.n387 71.676
R1023 B.n441 B.n388 71.676
R1024 B.n437 B.n389 71.676
R1025 B.n433 B.n390 71.676
R1026 B.n429 B.n391 71.676
R1027 B.n425 B.n392 71.676
R1028 B.n421 B.n393 71.676
R1029 B.n417 B.n394 71.676
R1030 B.n413 B.n395 71.676
R1031 B.n409 B.n396 71.676
R1032 B.n762 B.n761 71.676
R1033 B.n134 B.n96 71.676
R1034 B.n138 B.n97 71.676
R1035 B.n142 B.n98 71.676
R1036 B.n146 B.n99 71.676
R1037 B.n150 B.n100 71.676
R1038 B.n154 B.n101 71.676
R1039 B.n158 B.n102 71.676
R1040 B.n162 B.n103 71.676
R1041 B.n166 B.n104 71.676
R1042 B.n170 B.n105 71.676
R1043 B.n174 B.n106 71.676
R1044 B.n178 B.n107 71.676
R1045 B.n182 B.n108 71.676
R1046 B.n186 B.n109 71.676
R1047 B.n191 B.n110 71.676
R1048 B.n195 B.n111 71.676
R1049 B.n199 B.n112 71.676
R1050 B.n203 B.n113 71.676
R1051 B.n207 B.n114 71.676
R1052 B.n212 B.n115 71.676
R1053 B.n216 B.n116 71.676
R1054 B.n220 B.n117 71.676
R1055 B.n224 B.n118 71.676
R1056 B.n228 B.n119 71.676
R1057 B.n232 B.n120 71.676
R1058 B.n236 B.n121 71.676
R1059 B.n240 B.n122 71.676
R1060 B.n244 B.n123 71.676
R1061 B.n248 B.n124 71.676
R1062 B.n252 B.n125 71.676
R1063 B.n256 B.n126 71.676
R1064 B.n260 B.n127 71.676
R1065 B.n759 B.n128 71.676
R1066 B.n759 B.n758 71.676
R1067 B.n262 B.n127 71.676
R1068 B.n259 B.n126 71.676
R1069 B.n255 B.n125 71.676
R1070 B.n251 B.n124 71.676
R1071 B.n247 B.n123 71.676
R1072 B.n243 B.n122 71.676
R1073 B.n239 B.n121 71.676
R1074 B.n235 B.n120 71.676
R1075 B.n231 B.n119 71.676
R1076 B.n227 B.n118 71.676
R1077 B.n223 B.n117 71.676
R1078 B.n219 B.n116 71.676
R1079 B.n215 B.n115 71.676
R1080 B.n211 B.n114 71.676
R1081 B.n206 B.n113 71.676
R1082 B.n202 B.n112 71.676
R1083 B.n198 B.n111 71.676
R1084 B.n194 B.n110 71.676
R1085 B.n190 B.n109 71.676
R1086 B.n185 B.n108 71.676
R1087 B.n181 B.n107 71.676
R1088 B.n177 B.n106 71.676
R1089 B.n173 B.n105 71.676
R1090 B.n169 B.n104 71.676
R1091 B.n165 B.n103 71.676
R1092 B.n161 B.n102 71.676
R1093 B.n157 B.n101 71.676
R1094 B.n153 B.n100 71.676
R1095 B.n149 B.n99 71.676
R1096 B.n145 B.n98 71.676
R1097 B.n141 B.n97 71.676
R1098 B.n137 B.n96 71.676
R1099 B.n761 B.n95 71.676
R1100 B.n536 B.n364 71.676
R1101 B.n530 B.n365 71.676
R1102 B.n526 B.n366 71.676
R1103 B.n522 B.n367 71.676
R1104 B.n518 B.n368 71.676
R1105 B.n514 B.n369 71.676
R1106 B.n510 B.n370 71.676
R1107 B.n506 B.n371 71.676
R1108 B.n502 B.n372 71.676
R1109 B.n498 B.n373 71.676
R1110 B.n494 B.n374 71.676
R1111 B.n490 B.n375 71.676
R1112 B.n486 B.n376 71.676
R1113 B.n482 B.n377 71.676
R1114 B.n478 B.n378 71.676
R1115 B.n474 B.n379 71.676
R1116 B.n470 B.n380 71.676
R1117 B.n466 B.n381 71.676
R1118 B.n462 B.n382 71.676
R1119 B.n458 B.n383 71.676
R1120 B.n454 B.n384 71.676
R1121 B.n450 B.n385 71.676
R1122 B.n446 B.n386 71.676
R1123 B.n442 B.n387 71.676
R1124 B.n438 B.n388 71.676
R1125 B.n434 B.n389 71.676
R1126 B.n430 B.n390 71.676
R1127 B.n426 B.n391 71.676
R1128 B.n422 B.n392 71.676
R1129 B.n418 B.n393 71.676
R1130 B.n414 B.n394 71.676
R1131 B.n410 B.n395 71.676
R1132 B.n406 B.n396 71.676
R1133 B.n403 B.n402 70.7884
R1134 B.n400 B.n399 70.7884
R1135 B.n133 B.n132 70.7884
R1136 B.n131 B.n130 70.7884
R1137 B.n404 B.n403 59.5399
R1138 B.n401 B.n400 59.5399
R1139 B.n188 B.n133 59.5399
R1140 B.n209 B.n131 59.5399
R1141 B.n542 B.n361 57.2089
R1142 B.n542 B.n357 57.2089
R1143 B.n548 B.n357 57.2089
R1144 B.n548 B.n353 57.2089
R1145 B.n554 B.n353 57.2089
R1146 B.n554 B.n349 57.2089
R1147 B.n561 B.n349 57.2089
R1148 B.n561 B.n560 57.2089
R1149 B.n567 B.n342 57.2089
R1150 B.n573 B.n342 57.2089
R1151 B.n573 B.n338 57.2089
R1152 B.n579 B.n338 57.2089
R1153 B.n579 B.n334 57.2089
R1154 B.n585 B.n334 57.2089
R1155 B.n585 B.n330 57.2089
R1156 B.n591 B.n330 57.2089
R1157 B.n591 B.n326 57.2089
R1158 B.n597 B.n326 57.2089
R1159 B.n597 B.n321 57.2089
R1160 B.n603 B.n321 57.2089
R1161 B.n603 B.n322 57.2089
R1162 B.n609 B.n314 57.2089
R1163 B.n615 B.n314 57.2089
R1164 B.n615 B.n310 57.2089
R1165 B.n621 B.n310 57.2089
R1166 B.n621 B.n306 57.2089
R1167 B.n627 B.n306 57.2089
R1168 B.n627 B.n302 57.2089
R1169 B.n633 B.n302 57.2089
R1170 B.n633 B.n298 57.2089
R1171 B.n639 B.n298 57.2089
R1172 B.n645 B.n294 57.2089
R1173 B.n645 B.n290 57.2089
R1174 B.n651 B.n290 57.2089
R1175 B.n651 B.n286 57.2089
R1176 B.n657 B.n286 57.2089
R1177 B.n657 B.n282 57.2089
R1178 B.n663 B.n282 57.2089
R1179 B.n663 B.n278 57.2089
R1180 B.n670 B.n278 57.2089
R1181 B.n670 B.n669 57.2089
R1182 B.n676 B.n271 57.2089
R1183 B.n683 B.n271 57.2089
R1184 B.n683 B.n267 57.2089
R1185 B.n689 B.n267 57.2089
R1186 B.n689 B.n4 57.2089
R1187 B.n865 B.n4 57.2089
R1188 B.n865 B.n864 57.2089
R1189 B.n864 B.n863 57.2089
R1190 B.n863 B.n8 57.2089
R1191 B.n857 B.n8 57.2089
R1192 B.n857 B.n856 57.2089
R1193 B.n856 B.n855 57.2089
R1194 B.n849 B.n18 57.2089
R1195 B.n849 B.n848 57.2089
R1196 B.n848 B.n847 57.2089
R1197 B.n847 B.n22 57.2089
R1198 B.n841 B.n22 57.2089
R1199 B.n841 B.n840 57.2089
R1200 B.n840 B.n839 57.2089
R1201 B.n839 B.n29 57.2089
R1202 B.n833 B.n29 57.2089
R1203 B.n833 B.n832 57.2089
R1204 B.n831 B.n36 57.2089
R1205 B.n825 B.n36 57.2089
R1206 B.n825 B.n824 57.2089
R1207 B.n824 B.n823 57.2089
R1208 B.n823 B.n43 57.2089
R1209 B.n817 B.n43 57.2089
R1210 B.n817 B.n816 57.2089
R1211 B.n816 B.n815 57.2089
R1212 B.n815 B.n50 57.2089
R1213 B.n809 B.n50 57.2089
R1214 B.n808 B.n807 57.2089
R1215 B.n807 B.n57 57.2089
R1216 B.n801 B.n57 57.2089
R1217 B.n801 B.n800 57.2089
R1218 B.n800 B.n799 57.2089
R1219 B.n799 B.n64 57.2089
R1220 B.n793 B.n64 57.2089
R1221 B.n793 B.n792 57.2089
R1222 B.n792 B.n791 57.2089
R1223 B.n791 B.n71 57.2089
R1224 B.n785 B.n71 57.2089
R1225 B.n785 B.n784 57.2089
R1226 B.n784 B.n783 57.2089
R1227 B.n777 B.n81 57.2089
R1228 B.n777 B.n776 57.2089
R1229 B.n776 B.n775 57.2089
R1230 B.n775 B.n85 57.2089
R1231 B.n769 B.n85 57.2089
R1232 B.n769 B.n768 57.2089
R1233 B.n768 B.n767 57.2089
R1234 B.n767 B.n92 57.2089
R1235 B.n676 B.t1 55.5263
R1236 B.n855 B.t3 55.5263
R1237 B.t2 B.n294 40.3829
R1238 B.n832 B.t4 40.3829
R1239 B.n560 B.t14 35.3351
R1240 B.n81 B.t7 35.3351
R1241 B.n764 B.n763 33.5615
R1242 B.n757 B.n756 33.5615
R1243 B.n405 B.n359 33.5615
R1244 B.n539 B.n538 33.5615
R1245 B.n322 B.t0 31.9699
R1246 B.t5 B.n808 31.9699
R1247 B.n609 B.t0 25.2395
R1248 B.n809 B.t5 25.2395
R1249 B.n567 B.t14 21.8743
R1250 B.n783 B.t7 21.8743
R1251 B B.n867 18.0485
R1252 B.n639 B.t2 16.8265
R1253 B.t4 B.n831 16.8265
R1254 B.n763 B.n94 10.6151
R1255 B.n135 B.n94 10.6151
R1256 B.n136 B.n135 10.6151
R1257 B.n139 B.n136 10.6151
R1258 B.n140 B.n139 10.6151
R1259 B.n143 B.n140 10.6151
R1260 B.n144 B.n143 10.6151
R1261 B.n147 B.n144 10.6151
R1262 B.n148 B.n147 10.6151
R1263 B.n151 B.n148 10.6151
R1264 B.n152 B.n151 10.6151
R1265 B.n155 B.n152 10.6151
R1266 B.n156 B.n155 10.6151
R1267 B.n159 B.n156 10.6151
R1268 B.n160 B.n159 10.6151
R1269 B.n163 B.n160 10.6151
R1270 B.n164 B.n163 10.6151
R1271 B.n167 B.n164 10.6151
R1272 B.n168 B.n167 10.6151
R1273 B.n171 B.n168 10.6151
R1274 B.n172 B.n171 10.6151
R1275 B.n175 B.n172 10.6151
R1276 B.n176 B.n175 10.6151
R1277 B.n179 B.n176 10.6151
R1278 B.n180 B.n179 10.6151
R1279 B.n183 B.n180 10.6151
R1280 B.n184 B.n183 10.6151
R1281 B.n187 B.n184 10.6151
R1282 B.n192 B.n189 10.6151
R1283 B.n193 B.n192 10.6151
R1284 B.n196 B.n193 10.6151
R1285 B.n197 B.n196 10.6151
R1286 B.n200 B.n197 10.6151
R1287 B.n201 B.n200 10.6151
R1288 B.n204 B.n201 10.6151
R1289 B.n205 B.n204 10.6151
R1290 B.n208 B.n205 10.6151
R1291 B.n213 B.n210 10.6151
R1292 B.n214 B.n213 10.6151
R1293 B.n217 B.n214 10.6151
R1294 B.n218 B.n217 10.6151
R1295 B.n221 B.n218 10.6151
R1296 B.n222 B.n221 10.6151
R1297 B.n225 B.n222 10.6151
R1298 B.n226 B.n225 10.6151
R1299 B.n229 B.n226 10.6151
R1300 B.n230 B.n229 10.6151
R1301 B.n233 B.n230 10.6151
R1302 B.n234 B.n233 10.6151
R1303 B.n237 B.n234 10.6151
R1304 B.n238 B.n237 10.6151
R1305 B.n241 B.n238 10.6151
R1306 B.n242 B.n241 10.6151
R1307 B.n245 B.n242 10.6151
R1308 B.n246 B.n245 10.6151
R1309 B.n249 B.n246 10.6151
R1310 B.n250 B.n249 10.6151
R1311 B.n253 B.n250 10.6151
R1312 B.n254 B.n253 10.6151
R1313 B.n257 B.n254 10.6151
R1314 B.n258 B.n257 10.6151
R1315 B.n261 B.n258 10.6151
R1316 B.n263 B.n261 10.6151
R1317 B.n264 B.n263 10.6151
R1318 B.n757 B.n264 10.6151
R1319 B.n544 B.n359 10.6151
R1320 B.n545 B.n544 10.6151
R1321 B.n546 B.n545 10.6151
R1322 B.n546 B.n351 10.6151
R1323 B.n556 B.n351 10.6151
R1324 B.n557 B.n556 10.6151
R1325 B.n558 B.n557 10.6151
R1326 B.n558 B.n344 10.6151
R1327 B.n569 B.n344 10.6151
R1328 B.n570 B.n569 10.6151
R1329 B.n571 B.n570 10.6151
R1330 B.n571 B.n336 10.6151
R1331 B.n581 B.n336 10.6151
R1332 B.n582 B.n581 10.6151
R1333 B.n583 B.n582 10.6151
R1334 B.n583 B.n328 10.6151
R1335 B.n593 B.n328 10.6151
R1336 B.n594 B.n593 10.6151
R1337 B.n595 B.n594 10.6151
R1338 B.n595 B.n319 10.6151
R1339 B.n605 B.n319 10.6151
R1340 B.n606 B.n605 10.6151
R1341 B.n607 B.n606 10.6151
R1342 B.n607 B.n312 10.6151
R1343 B.n617 B.n312 10.6151
R1344 B.n618 B.n617 10.6151
R1345 B.n619 B.n618 10.6151
R1346 B.n619 B.n304 10.6151
R1347 B.n629 B.n304 10.6151
R1348 B.n630 B.n629 10.6151
R1349 B.n631 B.n630 10.6151
R1350 B.n631 B.n296 10.6151
R1351 B.n641 B.n296 10.6151
R1352 B.n642 B.n641 10.6151
R1353 B.n643 B.n642 10.6151
R1354 B.n643 B.n288 10.6151
R1355 B.n653 B.n288 10.6151
R1356 B.n654 B.n653 10.6151
R1357 B.n655 B.n654 10.6151
R1358 B.n655 B.n280 10.6151
R1359 B.n665 B.n280 10.6151
R1360 B.n666 B.n665 10.6151
R1361 B.n667 B.n666 10.6151
R1362 B.n667 B.n273 10.6151
R1363 B.n678 B.n273 10.6151
R1364 B.n679 B.n678 10.6151
R1365 B.n681 B.n679 10.6151
R1366 B.n681 B.n680 10.6151
R1367 B.n680 B.n265 10.6151
R1368 B.n692 B.n265 10.6151
R1369 B.n693 B.n692 10.6151
R1370 B.n694 B.n693 10.6151
R1371 B.n695 B.n694 10.6151
R1372 B.n697 B.n695 10.6151
R1373 B.n698 B.n697 10.6151
R1374 B.n699 B.n698 10.6151
R1375 B.n700 B.n699 10.6151
R1376 B.n702 B.n700 10.6151
R1377 B.n703 B.n702 10.6151
R1378 B.n704 B.n703 10.6151
R1379 B.n705 B.n704 10.6151
R1380 B.n707 B.n705 10.6151
R1381 B.n708 B.n707 10.6151
R1382 B.n709 B.n708 10.6151
R1383 B.n710 B.n709 10.6151
R1384 B.n712 B.n710 10.6151
R1385 B.n713 B.n712 10.6151
R1386 B.n714 B.n713 10.6151
R1387 B.n715 B.n714 10.6151
R1388 B.n717 B.n715 10.6151
R1389 B.n718 B.n717 10.6151
R1390 B.n719 B.n718 10.6151
R1391 B.n720 B.n719 10.6151
R1392 B.n722 B.n720 10.6151
R1393 B.n723 B.n722 10.6151
R1394 B.n724 B.n723 10.6151
R1395 B.n725 B.n724 10.6151
R1396 B.n727 B.n725 10.6151
R1397 B.n728 B.n727 10.6151
R1398 B.n729 B.n728 10.6151
R1399 B.n730 B.n729 10.6151
R1400 B.n732 B.n730 10.6151
R1401 B.n733 B.n732 10.6151
R1402 B.n734 B.n733 10.6151
R1403 B.n735 B.n734 10.6151
R1404 B.n737 B.n735 10.6151
R1405 B.n738 B.n737 10.6151
R1406 B.n739 B.n738 10.6151
R1407 B.n740 B.n739 10.6151
R1408 B.n742 B.n740 10.6151
R1409 B.n743 B.n742 10.6151
R1410 B.n744 B.n743 10.6151
R1411 B.n745 B.n744 10.6151
R1412 B.n747 B.n745 10.6151
R1413 B.n748 B.n747 10.6151
R1414 B.n749 B.n748 10.6151
R1415 B.n750 B.n749 10.6151
R1416 B.n752 B.n750 10.6151
R1417 B.n753 B.n752 10.6151
R1418 B.n754 B.n753 10.6151
R1419 B.n755 B.n754 10.6151
R1420 B.n756 B.n755 10.6151
R1421 B.n538 B.n363 10.6151
R1422 B.n533 B.n363 10.6151
R1423 B.n533 B.n532 10.6151
R1424 B.n532 B.n531 10.6151
R1425 B.n531 B.n528 10.6151
R1426 B.n528 B.n527 10.6151
R1427 B.n527 B.n524 10.6151
R1428 B.n524 B.n523 10.6151
R1429 B.n523 B.n520 10.6151
R1430 B.n520 B.n519 10.6151
R1431 B.n519 B.n516 10.6151
R1432 B.n516 B.n515 10.6151
R1433 B.n515 B.n512 10.6151
R1434 B.n512 B.n511 10.6151
R1435 B.n511 B.n508 10.6151
R1436 B.n508 B.n507 10.6151
R1437 B.n507 B.n504 10.6151
R1438 B.n504 B.n503 10.6151
R1439 B.n503 B.n500 10.6151
R1440 B.n500 B.n499 10.6151
R1441 B.n499 B.n496 10.6151
R1442 B.n496 B.n495 10.6151
R1443 B.n495 B.n492 10.6151
R1444 B.n492 B.n491 10.6151
R1445 B.n491 B.n488 10.6151
R1446 B.n488 B.n487 10.6151
R1447 B.n487 B.n484 10.6151
R1448 B.n484 B.n483 10.6151
R1449 B.n480 B.n479 10.6151
R1450 B.n479 B.n476 10.6151
R1451 B.n476 B.n475 10.6151
R1452 B.n475 B.n472 10.6151
R1453 B.n472 B.n471 10.6151
R1454 B.n471 B.n468 10.6151
R1455 B.n468 B.n467 10.6151
R1456 B.n467 B.n464 10.6151
R1457 B.n464 B.n463 10.6151
R1458 B.n460 B.n459 10.6151
R1459 B.n459 B.n456 10.6151
R1460 B.n456 B.n455 10.6151
R1461 B.n455 B.n452 10.6151
R1462 B.n452 B.n451 10.6151
R1463 B.n451 B.n448 10.6151
R1464 B.n448 B.n447 10.6151
R1465 B.n447 B.n444 10.6151
R1466 B.n444 B.n443 10.6151
R1467 B.n443 B.n440 10.6151
R1468 B.n440 B.n439 10.6151
R1469 B.n439 B.n436 10.6151
R1470 B.n436 B.n435 10.6151
R1471 B.n435 B.n432 10.6151
R1472 B.n432 B.n431 10.6151
R1473 B.n431 B.n428 10.6151
R1474 B.n428 B.n427 10.6151
R1475 B.n427 B.n424 10.6151
R1476 B.n424 B.n423 10.6151
R1477 B.n423 B.n420 10.6151
R1478 B.n420 B.n419 10.6151
R1479 B.n419 B.n416 10.6151
R1480 B.n416 B.n415 10.6151
R1481 B.n415 B.n412 10.6151
R1482 B.n412 B.n411 10.6151
R1483 B.n411 B.n408 10.6151
R1484 B.n408 B.n407 10.6151
R1485 B.n407 B.n405 10.6151
R1486 B.n540 B.n539 10.6151
R1487 B.n540 B.n355 10.6151
R1488 B.n550 B.n355 10.6151
R1489 B.n551 B.n550 10.6151
R1490 B.n552 B.n551 10.6151
R1491 B.n552 B.n347 10.6151
R1492 B.n563 B.n347 10.6151
R1493 B.n564 B.n563 10.6151
R1494 B.n565 B.n564 10.6151
R1495 B.n565 B.n340 10.6151
R1496 B.n575 B.n340 10.6151
R1497 B.n576 B.n575 10.6151
R1498 B.n577 B.n576 10.6151
R1499 B.n577 B.n332 10.6151
R1500 B.n587 B.n332 10.6151
R1501 B.n588 B.n587 10.6151
R1502 B.n589 B.n588 10.6151
R1503 B.n589 B.n324 10.6151
R1504 B.n599 B.n324 10.6151
R1505 B.n600 B.n599 10.6151
R1506 B.n601 B.n600 10.6151
R1507 B.n601 B.n316 10.6151
R1508 B.n611 B.n316 10.6151
R1509 B.n612 B.n611 10.6151
R1510 B.n613 B.n612 10.6151
R1511 B.n613 B.n308 10.6151
R1512 B.n623 B.n308 10.6151
R1513 B.n624 B.n623 10.6151
R1514 B.n625 B.n624 10.6151
R1515 B.n625 B.n300 10.6151
R1516 B.n635 B.n300 10.6151
R1517 B.n636 B.n635 10.6151
R1518 B.n637 B.n636 10.6151
R1519 B.n637 B.n292 10.6151
R1520 B.n647 B.n292 10.6151
R1521 B.n648 B.n647 10.6151
R1522 B.n649 B.n648 10.6151
R1523 B.n649 B.n284 10.6151
R1524 B.n659 B.n284 10.6151
R1525 B.n660 B.n659 10.6151
R1526 B.n661 B.n660 10.6151
R1527 B.n661 B.n276 10.6151
R1528 B.n672 B.n276 10.6151
R1529 B.n673 B.n672 10.6151
R1530 B.n674 B.n673 10.6151
R1531 B.n674 B.n269 10.6151
R1532 B.n685 B.n269 10.6151
R1533 B.n686 B.n685 10.6151
R1534 B.n687 B.n686 10.6151
R1535 B.n687 B.n0 10.6151
R1536 B.n861 B.n1 10.6151
R1537 B.n861 B.n860 10.6151
R1538 B.n860 B.n859 10.6151
R1539 B.n859 B.n10 10.6151
R1540 B.n853 B.n10 10.6151
R1541 B.n853 B.n852 10.6151
R1542 B.n852 B.n851 10.6151
R1543 B.n851 B.n16 10.6151
R1544 B.n845 B.n16 10.6151
R1545 B.n845 B.n844 10.6151
R1546 B.n844 B.n843 10.6151
R1547 B.n843 B.n24 10.6151
R1548 B.n837 B.n24 10.6151
R1549 B.n837 B.n836 10.6151
R1550 B.n836 B.n835 10.6151
R1551 B.n835 B.n31 10.6151
R1552 B.n829 B.n31 10.6151
R1553 B.n829 B.n828 10.6151
R1554 B.n828 B.n827 10.6151
R1555 B.n827 B.n38 10.6151
R1556 B.n821 B.n38 10.6151
R1557 B.n821 B.n820 10.6151
R1558 B.n820 B.n819 10.6151
R1559 B.n819 B.n45 10.6151
R1560 B.n813 B.n45 10.6151
R1561 B.n813 B.n812 10.6151
R1562 B.n812 B.n811 10.6151
R1563 B.n811 B.n52 10.6151
R1564 B.n805 B.n52 10.6151
R1565 B.n805 B.n804 10.6151
R1566 B.n804 B.n803 10.6151
R1567 B.n803 B.n59 10.6151
R1568 B.n797 B.n59 10.6151
R1569 B.n797 B.n796 10.6151
R1570 B.n796 B.n795 10.6151
R1571 B.n795 B.n66 10.6151
R1572 B.n789 B.n66 10.6151
R1573 B.n789 B.n788 10.6151
R1574 B.n788 B.n787 10.6151
R1575 B.n787 B.n73 10.6151
R1576 B.n781 B.n73 10.6151
R1577 B.n781 B.n780 10.6151
R1578 B.n780 B.n779 10.6151
R1579 B.n779 B.n79 10.6151
R1580 B.n773 B.n79 10.6151
R1581 B.n773 B.n772 10.6151
R1582 B.n772 B.n771 10.6151
R1583 B.n771 B.n87 10.6151
R1584 B.n765 B.n87 10.6151
R1585 B.n765 B.n764 10.6151
R1586 B.n188 B.n187 9.36635
R1587 B.n210 B.n209 9.36635
R1588 B.n483 B.n401 9.36635
R1589 B.n460 B.n404 9.36635
R1590 B.n867 B.n0 2.81026
R1591 B.n867 B.n1 2.81026
R1592 B.n669 B.t1 1.6831
R1593 B.n18 B.t3 1.6831
R1594 B.n189 B.n188 1.24928
R1595 B.n209 B.n208 1.24928
R1596 B.n480 B.n401 1.24928
R1597 B.n463 B.n404 1.24928
R1598 VP.n16 VP.n15 161.3
R1599 VP.n17 VP.n12 161.3
R1600 VP.n19 VP.n18 161.3
R1601 VP.n20 VP.n11 161.3
R1602 VP.n22 VP.n21 161.3
R1603 VP.n23 VP.n10 161.3
R1604 VP.n25 VP.n24 161.3
R1605 VP.n50 VP.n49 161.3
R1606 VP.n48 VP.n1 161.3
R1607 VP.n47 VP.n46 161.3
R1608 VP.n45 VP.n2 161.3
R1609 VP.n44 VP.n43 161.3
R1610 VP.n42 VP.n3 161.3
R1611 VP.n41 VP.n40 161.3
R1612 VP.n39 VP.n4 161.3
R1613 VP.n38 VP.n37 161.3
R1614 VP.n36 VP.n5 161.3
R1615 VP.n35 VP.n34 161.3
R1616 VP.n33 VP.n6 161.3
R1617 VP.n32 VP.n31 161.3
R1618 VP.n30 VP.n7 161.3
R1619 VP.n29 VP.n28 161.3
R1620 VP.n14 VP.t2 89.468
R1621 VP.n27 VP.n8 82.588
R1622 VP.n51 VP.n0 82.588
R1623 VP.n26 VP.n9 82.588
R1624 VP.n4 VP.t1 56.621
R1625 VP.n8 VP.t5 56.621
R1626 VP.n0 VP.t4 56.621
R1627 VP.n13 VP.t3 56.621
R1628 VP.n9 VP.t0 56.621
R1629 VP.n35 VP.n6 56.4773
R1630 VP.n43 VP.n2 56.4773
R1631 VP.n18 VP.n11 56.4773
R1632 VP.n14 VP.n13 49.9437
R1633 VP.n27 VP.n26 48.3211
R1634 VP.n30 VP.n29 24.3439
R1635 VP.n31 VP.n30 24.3439
R1636 VP.n31 VP.n6 24.3439
R1637 VP.n36 VP.n35 24.3439
R1638 VP.n37 VP.n36 24.3439
R1639 VP.n37 VP.n4 24.3439
R1640 VP.n41 VP.n4 24.3439
R1641 VP.n42 VP.n41 24.3439
R1642 VP.n43 VP.n42 24.3439
R1643 VP.n47 VP.n2 24.3439
R1644 VP.n48 VP.n47 24.3439
R1645 VP.n49 VP.n48 24.3439
R1646 VP.n22 VP.n11 24.3439
R1647 VP.n23 VP.n22 24.3439
R1648 VP.n24 VP.n23 24.3439
R1649 VP.n16 VP.n13 24.3439
R1650 VP.n17 VP.n16 24.3439
R1651 VP.n18 VP.n17 24.3439
R1652 VP.n29 VP.n8 7.30353
R1653 VP.n49 VP.n0 7.30353
R1654 VP.n24 VP.n9 7.30353
R1655 VP.n15 VP.n14 3.25662
R1656 VP.n26 VP.n25 0.355081
R1657 VP.n28 VP.n27 0.355081
R1658 VP.n51 VP.n50 0.355081
R1659 VP VP.n51 0.26685
R1660 VP.n15 VP.n12 0.189894
R1661 VP.n19 VP.n12 0.189894
R1662 VP.n20 VP.n19 0.189894
R1663 VP.n21 VP.n20 0.189894
R1664 VP.n21 VP.n10 0.189894
R1665 VP.n25 VP.n10 0.189894
R1666 VP.n28 VP.n7 0.189894
R1667 VP.n32 VP.n7 0.189894
R1668 VP.n33 VP.n32 0.189894
R1669 VP.n34 VP.n33 0.189894
R1670 VP.n34 VP.n5 0.189894
R1671 VP.n38 VP.n5 0.189894
R1672 VP.n39 VP.n38 0.189894
R1673 VP.n40 VP.n39 0.189894
R1674 VP.n40 VP.n3 0.189894
R1675 VP.n44 VP.n3 0.189894
R1676 VP.n45 VP.n44 0.189894
R1677 VP.n46 VP.n45 0.189894
R1678 VP.n46 VP.n1 0.189894
R1679 VP.n50 VP.n1 0.189894
R1680 VDD1 VDD1.t3 69.7891
R1681 VDD1.n1 VDD1.t0 69.6755
R1682 VDD1.n1 VDD1.n0 65.5639
R1683 VDD1.n3 VDD1.n2 64.8326
R1684 VDD1.n3 VDD1.n1 42.822
R1685 VDD1.n2 VDD1.t2 2.53896
R1686 VDD1.n2 VDD1.t5 2.53896
R1687 VDD1.n0 VDD1.t4 2.53896
R1688 VDD1.n0 VDD1.t1 2.53896
R1689 VDD1 VDD1.n3 0.728948
C0 VP VDD2 0.518856f
C1 VP VDD1 5.05639f
C2 VDD1 VDD2 1.6881f
C3 VP VTAIL 5.23365f
C4 VTAIL VDD2 6.60652f
C5 VTAIL VDD1 6.54946f
C6 VN VP 6.86011f
C7 VN VDD2 4.6915f
C8 VN VDD1 0.151482f
C9 VN VTAIL 5.21946f
C10 VDD2 B 5.797511f
C11 VDD1 B 6.154675f
C12 VTAIL B 6.584038f
C13 VN B 14.710939f
C14 VP B 13.427878f
C15 VDD1.t3 B 1.4996f
C16 VDD1.t0 B 1.49868f
C17 VDD1.t4 B 0.136011f
C18 VDD1.t1 B 0.136011f
C19 VDD1.n0 B 1.17226f
C20 VDD1.n1 B 2.73344f
C21 VDD1.t2 B 0.136011f
C22 VDD1.t5 B 0.136011f
C23 VDD1.n2 B 1.16704f
C24 VDD1.n3 B 2.35875f
C25 VP.t4 B 1.52995f
C26 VP.n0 B 0.631356f
C27 VP.n1 B 0.022023f
C28 VP.n2 B 0.027654f
C29 VP.n3 B 0.022023f
C30 VP.t1 B 1.52995f
C31 VP.n4 B 0.574002f
C32 VP.n5 B 0.022023f
C33 VP.n6 B 0.027654f
C34 VP.n7 B 0.022023f
C35 VP.t5 B 1.52995f
C36 VP.n8 B 0.631356f
C37 VP.t0 B 1.52995f
C38 VP.n9 B 0.631356f
C39 VP.n10 B 0.022023f
C40 VP.n11 B 0.027654f
C41 VP.n12 B 0.022023f
C42 VP.t3 B 1.52995f
C43 VP.n13 B 0.639804f
C44 VP.t2 B 1.79169f
C45 VP.n14 B 0.60219f
C46 VP.n15 B 0.268391f
C47 VP.n16 B 0.041251f
C48 VP.n17 B 0.041251f
C49 VP.n18 B 0.036924f
C50 VP.n19 B 0.022023f
C51 VP.n20 B 0.022023f
C52 VP.n21 B 0.022023f
C53 VP.n22 B 0.041251f
C54 VP.n23 B 0.041251f
C55 VP.n24 B 0.026994f
C56 VP.n25 B 0.03555f
C57 VP.n26 B 1.19625f
C58 VP.n27 B 1.21259f
C59 VP.n28 B 0.03555f
C60 VP.n29 B 0.026994f
C61 VP.n30 B 0.041251f
C62 VP.n31 B 0.041251f
C63 VP.n32 B 0.022023f
C64 VP.n33 B 0.022023f
C65 VP.n34 B 0.022023f
C66 VP.n35 B 0.036924f
C67 VP.n36 B 0.041251f
C68 VP.n37 B 0.041251f
C69 VP.n38 B 0.022023f
C70 VP.n39 B 0.022023f
C71 VP.n40 B 0.022023f
C72 VP.n41 B 0.041251f
C73 VP.n42 B 0.041251f
C74 VP.n43 B 0.036924f
C75 VP.n44 B 0.022023f
C76 VP.n45 B 0.022023f
C77 VP.n46 B 0.022023f
C78 VP.n47 B 0.041251f
C79 VP.n48 B 0.041251f
C80 VP.n49 B 0.026994f
C81 VP.n50 B 0.03555f
C82 VP.n51 B 0.059183f
C83 VDD2.t0 B 1.47025f
C84 VDD2.t3 B 0.133431f
C85 VDD2.t5 B 0.133431f
C86 VDD2.n0 B 1.15003f
C87 VDD2.n1 B 2.56122f
C88 VDD2.t4 B 1.45698f
C89 VDD2.n2 B 2.30461f
C90 VDD2.t1 B 0.133431f
C91 VDD2.t2 B 0.133431f
C92 VDD2.n3 B 1.15f
C93 VTAIL.t8 B 0.160141f
C94 VTAIL.t7 B 0.160141f
C95 VTAIL.n0 B 1.30106f
C96 VTAIL.n1 B 0.495272f
C97 VTAIL.t1 B 1.6588f
C98 VTAIL.n2 B 0.766974f
C99 VTAIL.t0 B 0.160141f
C100 VTAIL.t2 B 0.160141f
C101 VTAIL.n3 B 1.30106f
C102 VTAIL.n4 B 1.9596f
C103 VTAIL.t9 B 0.160141f
C104 VTAIL.t11 B 0.160141f
C105 VTAIL.n5 B 1.30106f
C106 VTAIL.n6 B 1.9596f
C107 VTAIL.t10 B 1.65881f
C108 VTAIL.n7 B 0.766964f
C109 VTAIL.t3 B 0.160141f
C110 VTAIL.t4 B 0.160141f
C111 VTAIL.n8 B 1.30106f
C112 VTAIL.n9 B 0.687962f
C113 VTAIL.t5 B 1.6588f
C114 VTAIL.n10 B 1.77518f
C115 VTAIL.t6 B 1.6588f
C116 VTAIL.n11 B 1.70446f
C117 VN.t0 B 1.49169f
C118 VN.n0 B 0.615565f
C119 VN.n1 B 0.021472f
C120 VN.n2 B 0.026962f
C121 VN.n3 B 0.021472f
C122 VN.t2 B 1.49169f
C123 VN.n4 B 0.623802f
C124 VN.t5 B 1.74688f
C125 VN.n5 B 0.587129f
C126 VN.n6 B 0.261678f
C127 VN.n7 B 0.040219f
C128 VN.n8 B 0.040219f
C129 VN.n9 B 0.036001f
C130 VN.n10 B 0.021472f
C131 VN.n11 B 0.021472f
C132 VN.n12 B 0.021472f
C133 VN.n13 B 0.040219f
C134 VN.n14 B 0.040219f
C135 VN.n15 B 0.026319f
C136 VN.n16 B 0.034661f
C137 VN.n17 B 0.057703f
C138 VN.t1 B 1.49169f
C139 VN.n18 B 0.615565f
C140 VN.n19 B 0.021472f
C141 VN.n20 B 0.026962f
C142 VN.n21 B 0.021472f
C143 VN.t4 B 1.49169f
C144 VN.n22 B 0.623802f
C145 VN.t3 B 1.74688f
C146 VN.n23 B 0.587129f
C147 VN.n24 B 0.261678f
C148 VN.n25 B 0.040219f
C149 VN.n26 B 0.040219f
C150 VN.n27 B 0.036001f
C151 VN.n28 B 0.021472f
C152 VN.n29 B 0.021472f
C153 VN.n30 B 0.021472f
C154 VN.n31 B 0.040219f
C155 VN.n32 B 0.040219f
C156 VN.n33 B 0.026319f
C157 VN.n34 B 0.034661f
C158 VN.n35 B 1.17524f
.ends

