* NGSPICE file created from diff_pair_sample_1471.ext - technology: sky130A

.subckt diff_pair_sample_1471 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=0.53
X1 B.t11 B.t9 B.t10 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=0.53
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=0.53
X3 VDD1.t0 VP.t1 VTAIL.t2 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=0.53
X4 B.t8 B.t6 B.t7 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=0.53
X5 B.t5 B.t3 B.t4 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=0.53
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=0.53
X7 B.t2 B.t0 B.t1 w_n1314_n1562# sky130_fd_pr__pfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=0.53
R0 VP.n0 VP.t1 402.341
R1 VP.n0 VP.t0 370.015
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t0 136.095
R4 VTAIL.n3 VTAIL.t3 136.095
R5 VTAIL.n0 VTAIL.t1 136.095
R6 VTAIL.n2 VTAIL.t2 136.095
R7 VTAIL.n1 VTAIL.n0 16.41
R8 VTAIL.n3 VTAIL.n2 15.6686
R9 VTAIL.n2 VTAIL.n1 0.841017
R10 VTAIL VTAIL.n0 0.713862
R11 VTAIL VTAIL.n3 0.127655
R12 VDD1 VDD1.t1 181.186
R13 VDD1 VDD1.t0 153.017
R14 B.n198 B.n197 585
R15 B.n199 B.n32 585
R16 B.n201 B.n200 585
R17 B.n202 B.n31 585
R18 B.n204 B.n203 585
R19 B.n205 B.n30 585
R20 B.n207 B.n206 585
R21 B.n208 B.n29 585
R22 B.n210 B.n209 585
R23 B.n211 B.n28 585
R24 B.n213 B.n212 585
R25 B.n214 B.n27 585
R26 B.n216 B.n215 585
R27 B.n217 B.n26 585
R28 B.n219 B.n218 585
R29 B.n221 B.n23 585
R30 B.n223 B.n222 585
R31 B.n224 B.n22 585
R32 B.n226 B.n225 585
R33 B.n227 B.n21 585
R34 B.n229 B.n228 585
R35 B.n230 B.n20 585
R36 B.n232 B.n231 585
R37 B.n233 B.n19 585
R38 B.n235 B.n234 585
R39 B.n237 B.n236 585
R40 B.n238 B.n15 585
R41 B.n240 B.n239 585
R42 B.n241 B.n14 585
R43 B.n243 B.n242 585
R44 B.n244 B.n13 585
R45 B.n246 B.n245 585
R46 B.n247 B.n12 585
R47 B.n249 B.n248 585
R48 B.n250 B.n11 585
R49 B.n252 B.n251 585
R50 B.n253 B.n10 585
R51 B.n255 B.n254 585
R52 B.n256 B.n9 585
R53 B.n258 B.n257 585
R54 B.n196 B.n33 585
R55 B.n195 B.n194 585
R56 B.n193 B.n34 585
R57 B.n192 B.n191 585
R58 B.n190 B.n35 585
R59 B.n189 B.n188 585
R60 B.n187 B.n36 585
R61 B.n186 B.n185 585
R62 B.n184 B.n37 585
R63 B.n183 B.n182 585
R64 B.n181 B.n38 585
R65 B.n180 B.n179 585
R66 B.n178 B.n39 585
R67 B.n177 B.n176 585
R68 B.n175 B.n40 585
R69 B.n174 B.n173 585
R70 B.n172 B.n41 585
R71 B.n171 B.n170 585
R72 B.n169 B.n42 585
R73 B.n168 B.n167 585
R74 B.n166 B.n43 585
R75 B.n165 B.n164 585
R76 B.n163 B.n44 585
R77 B.n162 B.n161 585
R78 B.n160 B.n45 585
R79 B.n159 B.n158 585
R80 B.n157 B.n46 585
R81 B.n96 B.n95 585
R82 B.n97 B.n70 585
R83 B.n99 B.n98 585
R84 B.n100 B.n69 585
R85 B.n102 B.n101 585
R86 B.n103 B.n68 585
R87 B.n105 B.n104 585
R88 B.n106 B.n67 585
R89 B.n108 B.n107 585
R90 B.n109 B.n66 585
R91 B.n111 B.n110 585
R92 B.n112 B.n65 585
R93 B.n114 B.n113 585
R94 B.n115 B.n64 585
R95 B.n117 B.n116 585
R96 B.n119 B.n61 585
R97 B.n121 B.n120 585
R98 B.n122 B.n60 585
R99 B.n124 B.n123 585
R100 B.n125 B.n59 585
R101 B.n127 B.n126 585
R102 B.n128 B.n58 585
R103 B.n130 B.n129 585
R104 B.n131 B.n57 585
R105 B.n133 B.n132 585
R106 B.n135 B.n134 585
R107 B.n136 B.n53 585
R108 B.n138 B.n137 585
R109 B.n139 B.n52 585
R110 B.n141 B.n140 585
R111 B.n142 B.n51 585
R112 B.n144 B.n143 585
R113 B.n145 B.n50 585
R114 B.n147 B.n146 585
R115 B.n148 B.n49 585
R116 B.n150 B.n149 585
R117 B.n151 B.n48 585
R118 B.n153 B.n152 585
R119 B.n154 B.n47 585
R120 B.n156 B.n155 585
R121 B.n94 B.n71 585
R122 B.n93 B.n92 585
R123 B.n91 B.n72 585
R124 B.n90 B.n89 585
R125 B.n88 B.n73 585
R126 B.n87 B.n86 585
R127 B.n85 B.n74 585
R128 B.n84 B.n83 585
R129 B.n82 B.n75 585
R130 B.n81 B.n80 585
R131 B.n79 B.n76 585
R132 B.n78 B.n77 585
R133 B.n2 B.n0 585
R134 B.n277 B.n1 585
R135 B.n276 B.n275 585
R136 B.n274 B.n3 585
R137 B.n273 B.n272 585
R138 B.n271 B.n4 585
R139 B.n270 B.n269 585
R140 B.n268 B.n5 585
R141 B.n267 B.n266 585
R142 B.n265 B.n6 585
R143 B.n264 B.n263 585
R144 B.n262 B.n7 585
R145 B.n261 B.n260 585
R146 B.n259 B.n8 585
R147 B.n279 B.n278 585
R148 B.n96 B.n71 502.111
R149 B.n259 B.n258 502.111
R150 B.n157 B.n156 502.111
R151 B.n198 B.n33 502.111
R152 B.n54 B.t9 339.868
R153 B.n62 B.t0 339.868
R154 B.n16 B.t6 339.868
R155 B.n24 B.t3 339.868
R156 B.n92 B.n71 163.367
R157 B.n92 B.n91 163.367
R158 B.n91 B.n90 163.367
R159 B.n90 B.n73 163.367
R160 B.n86 B.n73 163.367
R161 B.n86 B.n85 163.367
R162 B.n85 B.n84 163.367
R163 B.n84 B.n75 163.367
R164 B.n80 B.n75 163.367
R165 B.n80 B.n79 163.367
R166 B.n79 B.n78 163.367
R167 B.n78 B.n2 163.367
R168 B.n278 B.n2 163.367
R169 B.n278 B.n277 163.367
R170 B.n277 B.n276 163.367
R171 B.n276 B.n3 163.367
R172 B.n272 B.n3 163.367
R173 B.n272 B.n271 163.367
R174 B.n271 B.n270 163.367
R175 B.n270 B.n5 163.367
R176 B.n266 B.n5 163.367
R177 B.n266 B.n265 163.367
R178 B.n265 B.n264 163.367
R179 B.n264 B.n7 163.367
R180 B.n260 B.n7 163.367
R181 B.n260 B.n259 163.367
R182 B.n97 B.n96 163.367
R183 B.n98 B.n97 163.367
R184 B.n98 B.n69 163.367
R185 B.n102 B.n69 163.367
R186 B.n103 B.n102 163.367
R187 B.n104 B.n103 163.367
R188 B.n104 B.n67 163.367
R189 B.n108 B.n67 163.367
R190 B.n109 B.n108 163.367
R191 B.n110 B.n109 163.367
R192 B.n110 B.n65 163.367
R193 B.n114 B.n65 163.367
R194 B.n115 B.n114 163.367
R195 B.n116 B.n115 163.367
R196 B.n116 B.n61 163.367
R197 B.n121 B.n61 163.367
R198 B.n122 B.n121 163.367
R199 B.n123 B.n122 163.367
R200 B.n123 B.n59 163.367
R201 B.n127 B.n59 163.367
R202 B.n128 B.n127 163.367
R203 B.n129 B.n128 163.367
R204 B.n129 B.n57 163.367
R205 B.n133 B.n57 163.367
R206 B.n134 B.n133 163.367
R207 B.n134 B.n53 163.367
R208 B.n138 B.n53 163.367
R209 B.n139 B.n138 163.367
R210 B.n140 B.n139 163.367
R211 B.n140 B.n51 163.367
R212 B.n144 B.n51 163.367
R213 B.n145 B.n144 163.367
R214 B.n146 B.n145 163.367
R215 B.n146 B.n49 163.367
R216 B.n150 B.n49 163.367
R217 B.n151 B.n150 163.367
R218 B.n152 B.n151 163.367
R219 B.n152 B.n47 163.367
R220 B.n156 B.n47 163.367
R221 B.n158 B.n157 163.367
R222 B.n158 B.n45 163.367
R223 B.n162 B.n45 163.367
R224 B.n163 B.n162 163.367
R225 B.n164 B.n163 163.367
R226 B.n164 B.n43 163.367
R227 B.n168 B.n43 163.367
R228 B.n169 B.n168 163.367
R229 B.n170 B.n169 163.367
R230 B.n170 B.n41 163.367
R231 B.n174 B.n41 163.367
R232 B.n175 B.n174 163.367
R233 B.n176 B.n175 163.367
R234 B.n176 B.n39 163.367
R235 B.n180 B.n39 163.367
R236 B.n181 B.n180 163.367
R237 B.n182 B.n181 163.367
R238 B.n182 B.n37 163.367
R239 B.n186 B.n37 163.367
R240 B.n187 B.n186 163.367
R241 B.n188 B.n187 163.367
R242 B.n188 B.n35 163.367
R243 B.n192 B.n35 163.367
R244 B.n193 B.n192 163.367
R245 B.n194 B.n193 163.367
R246 B.n194 B.n33 163.367
R247 B.n258 B.n9 163.367
R248 B.n254 B.n9 163.367
R249 B.n254 B.n253 163.367
R250 B.n253 B.n252 163.367
R251 B.n252 B.n11 163.367
R252 B.n248 B.n11 163.367
R253 B.n248 B.n247 163.367
R254 B.n247 B.n246 163.367
R255 B.n246 B.n13 163.367
R256 B.n242 B.n13 163.367
R257 B.n242 B.n241 163.367
R258 B.n241 B.n240 163.367
R259 B.n240 B.n15 163.367
R260 B.n236 B.n15 163.367
R261 B.n236 B.n235 163.367
R262 B.n235 B.n19 163.367
R263 B.n231 B.n19 163.367
R264 B.n231 B.n230 163.367
R265 B.n230 B.n229 163.367
R266 B.n229 B.n21 163.367
R267 B.n225 B.n21 163.367
R268 B.n225 B.n224 163.367
R269 B.n224 B.n223 163.367
R270 B.n223 B.n23 163.367
R271 B.n218 B.n23 163.367
R272 B.n218 B.n217 163.367
R273 B.n217 B.n216 163.367
R274 B.n216 B.n27 163.367
R275 B.n212 B.n27 163.367
R276 B.n212 B.n211 163.367
R277 B.n211 B.n210 163.367
R278 B.n210 B.n29 163.367
R279 B.n206 B.n29 163.367
R280 B.n206 B.n205 163.367
R281 B.n205 B.n204 163.367
R282 B.n204 B.n31 163.367
R283 B.n200 B.n31 163.367
R284 B.n200 B.n199 163.367
R285 B.n199 B.n198 163.367
R286 B.n54 B.t11 161.115
R287 B.n24 B.t4 161.115
R288 B.n62 B.t2 161.113
R289 B.n16 B.t7 161.113
R290 B.n55 B.t10 144.436
R291 B.n25 B.t5 144.436
R292 B.n63 B.t1 144.435
R293 B.n17 B.t8 144.435
R294 B.n56 B.n55 59.5399
R295 B.n118 B.n63 59.5399
R296 B.n18 B.n17 59.5399
R297 B.n220 B.n25 59.5399
R298 B.n257 B.n8 32.6249
R299 B.n197 B.n196 32.6249
R300 B.n155 B.n46 32.6249
R301 B.n95 B.n94 32.6249
R302 B B.n279 18.0485
R303 B.n55 B.n54 16.6793
R304 B.n63 B.n62 16.6793
R305 B.n17 B.n16 16.6793
R306 B.n25 B.n24 16.6793
R307 B.n257 B.n256 10.6151
R308 B.n256 B.n255 10.6151
R309 B.n255 B.n10 10.6151
R310 B.n251 B.n10 10.6151
R311 B.n251 B.n250 10.6151
R312 B.n250 B.n249 10.6151
R313 B.n249 B.n12 10.6151
R314 B.n245 B.n12 10.6151
R315 B.n245 B.n244 10.6151
R316 B.n244 B.n243 10.6151
R317 B.n243 B.n14 10.6151
R318 B.n239 B.n14 10.6151
R319 B.n239 B.n238 10.6151
R320 B.n238 B.n237 10.6151
R321 B.n234 B.n233 10.6151
R322 B.n233 B.n232 10.6151
R323 B.n232 B.n20 10.6151
R324 B.n228 B.n20 10.6151
R325 B.n228 B.n227 10.6151
R326 B.n227 B.n226 10.6151
R327 B.n226 B.n22 10.6151
R328 B.n222 B.n22 10.6151
R329 B.n222 B.n221 10.6151
R330 B.n219 B.n26 10.6151
R331 B.n215 B.n26 10.6151
R332 B.n215 B.n214 10.6151
R333 B.n214 B.n213 10.6151
R334 B.n213 B.n28 10.6151
R335 B.n209 B.n28 10.6151
R336 B.n209 B.n208 10.6151
R337 B.n208 B.n207 10.6151
R338 B.n207 B.n30 10.6151
R339 B.n203 B.n30 10.6151
R340 B.n203 B.n202 10.6151
R341 B.n202 B.n201 10.6151
R342 B.n201 B.n32 10.6151
R343 B.n197 B.n32 10.6151
R344 B.n159 B.n46 10.6151
R345 B.n160 B.n159 10.6151
R346 B.n161 B.n160 10.6151
R347 B.n161 B.n44 10.6151
R348 B.n165 B.n44 10.6151
R349 B.n166 B.n165 10.6151
R350 B.n167 B.n166 10.6151
R351 B.n167 B.n42 10.6151
R352 B.n171 B.n42 10.6151
R353 B.n172 B.n171 10.6151
R354 B.n173 B.n172 10.6151
R355 B.n173 B.n40 10.6151
R356 B.n177 B.n40 10.6151
R357 B.n178 B.n177 10.6151
R358 B.n179 B.n178 10.6151
R359 B.n179 B.n38 10.6151
R360 B.n183 B.n38 10.6151
R361 B.n184 B.n183 10.6151
R362 B.n185 B.n184 10.6151
R363 B.n185 B.n36 10.6151
R364 B.n189 B.n36 10.6151
R365 B.n190 B.n189 10.6151
R366 B.n191 B.n190 10.6151
R367 B.n191 B.n34 10.6151
R368 B.n195 B.n34 10.6151
R369 B.n196 B.n195 10.6151
R370 B.n95 B.n70 10.6151
R371 B.n99 B.n70 10.6151
R372 B.n100 B.n99 10.6151
R373 B.n101 B.n100 10.6151
R374 B.n101 B.n68 10.6151
R375 B.n105 B.n68 10.6151
R376 B.n106 B.n105 10.6151
R377 B.n107 B.n106 10.6151
R378 B.n107 B.n66 10.6151
R379 B.n111 B.n66 10.6151
R380 B.n112 B.n111 10.6151
R381 B.n113 B.n112 10.6151
R382 B.n113 B.n64 10.6151
R383 B.n117 B.n64 10.6151
R384 B.n120 B.n119 10.6151
R385 B.n120 B.n60 10.6151
R386 B.n124 B.n60 10.6151
R387 B.n125 B.n124 10.6151
R388 B.n126 B.n125 10.6151
R389 B.n126 B.n58 10.6151
R390 B.n130 B.n58 10.6151
R391 B.n131 B.n130 10.6151
R392 B.n132 B.n131 10.6151
R393 B.n136 B.n135 10.6151
R394 B.n137 B.n136 10.6151
R395 B.n137 B.n52 10.6151
R396 B.n141 B.n52 10.6151
R397 B.n142 B.n141 10.6151
R398 B.n143 B.n142 10.6151
R399 B.n143 B.n50 10.6151
R400 B.n147 B.n50 10.6151
R401 B.n148 B.n147 10.6151
R402 B.n149 B.n148 10.6151
R403 B.n149 B.n48 10.6151
R404 B.n153 B.n48 10.6151
R405 B.n154 B.n153 10.6151
R406 B.n155 B.n154 10.6151
R407 B.n94 B.n93 10.6151
R408 B.n93 B.n72 10.6151
R409 B.n89 B.n72 10.6151
R410 B.n89 B.n88 10.6151
R411 B.n88 B.n87 10.6151
R412 B.n87 B.n74 10.6151
R413 B.n83 B.n74 10.6151
R414 B.n83 B.n82 10.6151
R415 B.n82 B.n81 10.6151
R416 B.n81 B.n76 10.6151
R417 B.n77 B.n76 10.6151
R418 B.n77 B.n0 10.6151
R419 B.n275 B.n1 10.6151
R420 B.n275 B.n274 10.6151
R421 B.n274 B.n273 10.6151
R422 B.n273 B.n4 10.6151
R423 B.n269 B.n4 10.6151
R424 B.n269 B.n268 10.6151
R425 B.n268 B.n267 10.6151
R426 B.n267 B.n6 10.6151
R427 B.n263 B.n6 10.6151
R428 B.n263 B.n262 10.6151
R429 B.n262 B.n261 10.6151
R430 B.n261 B.n8 10.6151
R431 B.n237 B.n18 8.74196
R432 B.n220 B.n219 8.74196
R433 B.n118 B.n117 8.74196
R434 B.n135 B.n56 8.74196
R435 B.n279 B.n0 2.81026
R436 B.n279 B.n1 2.81026
R437 B.n234 B.n18 1.87367
R438 B.n221 B.n220 1.87367
R439 B.n119 B.n118 1.87367
R440 B.n132 B.n56 1.87367
R441 VN VN.t1 402.723
R442 VN VN.t0 370.067
R443 VDD2.n0 VDD2.t1 180.476
R444 VDD2.n0 VDD2.t0 152.774
R445 VDD2 VDD2.n0 0.244034
C0 VDD1 VTAIL 2.36445f
C1 VDD1 B 0.733363f
C2 VTAIL VDD2 2.40201f
C3 VDD2 B 0.746802f
C4 VTAIL B 1.00852f
C5 VP VN 2.81532f
C6 VN w_n1314_n1562# 1.45236f
C7 VN VDD1 0.153643f
C8 VN VDD2 0.617457f
C9 VN VTAIL 0.557609f
C10 VN B 0.583852f
C11 VP w_n1314_n1562# 1.61286f
C12 VP VDD1 0.714144f
C13 VP VDD2 0.252067f
C14 VP VTAIL 0.571853f
C15 VP B 0.842948f
C16 w_n1314_n1562# VDD1 0.876764f
C17 w_n1314_n1562# VDD2 0.879187f
C18 w_n1314_n1562# VTAIL 1.39067f
C19 w_n1314_n1562# B 4.02608f
C20 VDD1 VDD2 0.443558f
C21 VDD2 VSUBS 0.414991f
C22 VDD1 VSUBS 2.21731f
C23 VTAIL VSUBS 0.146649f
C24 VN VSUBS 3.39776f
C25 VP VSUBS 0.652088f
C26 B VSUBS 1.5356f
C27 w_n1314_n1562# VSUBS 26.0014f
C28 VDD2.t1 VSUBS 0.414797f
C29 VDD2.t0 VSUBS 0.299673f
C30 VDD2.n0 VSUBS 1.6508f
C31 VN.t0 VSUBS 0.240547f
C32 VN.t1 VSUBS 0.332705f
C33 B.n0 VSUBS 0.005161f
C34 B.n1 VSUBS 0.005161f
C35 B.n2 VSUBS 0.008162f
C36 B.n3 VSUBS 0.008162f
C37 B.n4 VSUBS 0.008162f
C38 B.n5 VSUBS 0.008162f
C39 B.n6 VSUBS 0.008162f
C40 B.n7 VSUBS 0.008162f
C41 B.n8 VSUBS 0.018367f
C42 B.n9 VSUBS 0.008162f
C43 B.n10 VSUBS 0.008162f
C44 B.n11 VSUBS 0.008162f
C45 B.n12 VSUBS 0.008162f
C46 B.n13 VSUBS 0.008162f
C47 B.n14 VSUBS 0.008162f
C48 B.n15 VSUBS 0.008162f
C49 B.t8 VSUBS 0.082259f
C50 B.t7 VSUBS 0.087878f
C51 B.t6 VSUBS 0.082157f
C52 B.n16 VSUBS 0.072735f
C53 B.n17 VSUBS 0.065921f
C54 B.n18 VSUBS 0.018911f
C55 B.n19 VSUBS 0.008162f
C56 B.n20 VSUBS 0.008162f
C57 B.n21 VSUBS 0.008162f
C58 B.n22 VSUBS 0.008162f
C59 B.n23 VSUBS 0.008162f
C60 B.t5 VSUBS 0.082259f
C61 B.t4 VSUBS 0.087878f
C62 B.t3 VSUBS 0.082157f
C63 B.n24 VSUBS 0.072735f
C64 B.n25 VSUBS 0.065921f
C65 B.n26 VSUBS 0.008162f
C66 B.n27 VSUBS 0.008162f
C67 B.n28 VSUBS 0.008162f
C68 B.n29 VSUBS 0.008162f
C69 B.n30 VSUBS 0.008162f
C70 B.n31 VSUBS 0.008162f
C71 B.n32 VSUBS 0.008162f
C72 B.n33 VSUBS 0.018367f
C73 B.n34 VSUBS 0.008162f
C74 B.n35 VSUBS 0.008162f
C75 B.n36 VSUBS 0.008162f
C76 B.n37 VSUBS 0.008162f
C77 B.n38 VSUBS 0.008162f
C78 B.n39 VSUBS 0.008162f
C79 B.n40 VSUBS 0.008162f
C80 B.n41 VSUBS 0.008162f
C81 B.n42 VSUBS 0.008162f
C82 B.n43 VSUBS 0.008162f
C83 B.n44 VSUBS 0.008162f
C84 B.n45 VSUBS 0.008162f
C85 B.n46 VSUBS 0.018367f
C86 B.n47 VSUBS 0.008162f
C87 B.n48 VSUBS 0.008162f
C88 B.n49 VSUBS 0.008162f
C89 B.n50 VSUBS 0.008162f
C90 B.n51 VSUBS 0.008162f
C91 B.n52 VSUBS 0.008162f
C92 B.n53 VSUBS 0.008162f
C93 B.t10 VSUBS 0.082259f
C94 B.t11 VSUBS 0.087878f
C95 B.t9 VSUBS 0.082157f
C96 B.n54 VSUBS 0.072735f
C97 B.n55 VSUBS 0.065921f
C98 B.n56 VSUBS 0.018911f
C99 B.n57 VSUBS 0.008162f
C100 B.n58 VSUBS 0.008162f
C101 B.n59 VSUBS 0.008162f
C102 B.n60 VSUBS 0.008162f
C103 B.n61 VSUBS 0.008162f
C104 B.t1 VSUBS 0.082259f
C105 B.t2 VSUBS 0.087878f
C106 B.t0 VSUBS 0.082157f
C107 B.n62 VSUBS 0.072735f
C108 B.n63 VSUBS 0.065921f
C109 B.n64 VSUBS 0.008162f
C110 B.n65 VSUBS 0.008162f
C111 B.n66 VSUBS 0.008162f
C112 B.n67 VSUBS 0.008162f
C113 B.n68 VSUBS 0.008162f
C114 B.n69 VSUBS 0.008162f
C115 B.n70 VSUBS 0.008162f
C116 B.n71 VSUBS 0.018367f
C117 B.n72 VSUBS 0.008162f
C118 B.n73 VSUBS 0.008162f
C119 B.n74 VSUBS 0.008162f
C120 B.n75 VSUBS 0.008162f
C121 B.n76 VSUBS 0.008162f
C122 B.n77 VSUBS 0.008162f
C123 B.n78 VSUBS 0.008162f
C124 B.n79 VSUBS 0.008162f
C125 B.n80 VSUBS 0.008162f
C126 B.n81 VSUBS 0.008162f
C127 B.n82 VSUBS 0.008162f
C128 B.n83 VSUBS 0.008162f
C129 B.n84 VSUBS 0.008162f
C130 B.n85 VSUBS 0.008162f
C131 B.n86 VSUBS 0.008162f
C132 B.n87 VSUBS 0.008162f
C133 B.n88 VSUBS 0.008162f
C134 B.n89 VSUBS 0.008162f
C135 B.n90 VSUBS 0.008162f
C136 B.n91 VSUBS 0.008162f
C137 B.n92 VSUBS 0.008162f
C138 B.n93 VSUBS 0.008162f
C139 B.n94 VSUBS 0.018367f
C140 B.n95 VSUBS 0.019803f
C141 B.n96 VSUBS 0.019803f
C142 B.n97 VSUBS 0.008162f
C143 B.n98 VSUBS 0.008162f
C144 B.n99 VSUBS 0.008162f
C145 B.n100 VSUBS 0.008162f
C146 B.n101 VSUBS 0.008162f
C147 B.n102 VSUBS 0.008162f
C148 B.n103 VSUBS 0.008162f
C149 B.n104 VSUBS 0.008162f
C150 B.n105 VSUBS 0.008162f
C151 B.n106 VSUBS 0.008162f
C152 B.n107 VSUBS 0.008162f
C153 B.n108 VSUBS 0.008162f
C154 B.n109 VSUBS 0.008162f
C155 B.n110 VSUBS 0.008162f
C156 B.n111 VSUBS 0.008162f
C157 B.n112 VSUBS 0.008162f
C158 B.n113 VSUBS 0.008162f
C159 B.n114 VSUBS 0.008162f
C160 B.n115 VSUBS 0.008162f
C161 B.n116 VSUBS 0.008162f
C162 B.n117 VSUBS 0.007442f
C163 B.n118 VSUBS 0.018911f
C164 B.n119 VSUBS 0.004801f
C165 B.n120 VSUBS 0.008162f
C166 B.n121 VSUBS 0.008162f
C167 B.n122 VSUBS 0.008162f
C168 B.n123 VSUBS 0.008162f
C169 B.n124 VSUBS 0.008162f
C170 B.n125 VSUBS 0.008162f
C171 B.n126 VSUBS 0.008162f
C172 B.n127 VSUBS 0.008162f
C173 B.n128 VSUBS 0.008162f
C174 B.n129 VSUBS 0.008162f
C175 B.n130 VSUBS 0.008162f
C176 B.n131 VSUBS 0.008162f
C177 B.n132 VSUBS 0.004801f
C178 B.n133 VSUBS 0.008162f
C179 B.n134 VSUBS 0.008162f
C180 B.n135 VSUBS 0.007442f
C181 B.n136 VSUBS 0.008162f
C182 B.n137 VSUBS 0.008162f
C183 B.n138 VSUBS 0.008162f
C184 B.n139 VSUBS 0.008162f
C185 B.n140 VSUBS 0.008162f
C186 B.n141 VSUBS 0.008162f
C187 B.n142 VSUBS 0.008162f
C188 B.n143 VSUBS 0.008162f
C189 B.n144 VSUBS 0.008162f
C190 B.n145 VSUBS 0.008162f
C191 B.n146 VSUBS 0.008162f
C192 B.n147 VSUBS 0.008162f
C193 B.n148 VSUBS 0.008162f
C194 B.n149 VSUBS 0.008162f
C195 B.n150 VSUBS 0.008162f
C196 B.n151 VSUBS 0.008162f
C197 B.n152 VSUBS 0.008162f
C198 B.n153 VSUBS 0.008162f
C199 B.n154 VSUBS 0.008162f
C200 B.n155 VSUBS 0.019803f
C201 B.n156 VSUBS 0.019803f
C202 B.n157 VSUBS 0.018367f
C203 B.n158 VSUBS 0.008162f
C204 B.n159 VSUBS 0.008162f
C205 B.n160 VSUBS 0.008162f
C206 B.n161 VSUBS 0.008162f
C207 B.n162 VSUBS 0.008162f
C208 B.n163 VSUBS 0.008162f
C209 B.n164 VSUBS 0.008162f
C210 B.n165 VSUBS 0.008162f
C211 B.n166 VSUBS 0.008162f
C212 B.n167 VSUBS 0.008162f
C213 B.n168 VSUBS 0.008162f
C214 B.n169 VSUBS 0.008162f
C215 B.n170 VSUBS 0.008162f
C216 B.n171 VSUBS 0.008162f
C217 B.n172 VSUBS 0.008162f
C218 B.n173 VSUBS 0.008162f
C219 B.n174 VSUBS 0.008162f
C220 B.n175 VSUBS 0.008162f
C221 B.n176 VSUBS 0.008162f
C222 B.n177 VSUBS 0.008162f
C223 B.n178 VSUBS 0.008162f
C224 B.n179 VSUBS 0.008162f
C225 B.n180 VSUBS 0.008162f
C226 B.n181 VSUBS 0.008162f
C227 B.n182 VSUBS 0.008162f
C228 B.n183 VSUBS 0.008162f
C229 B.n184 VSUBS 0.008162f
C230 B.n185 VSUBS 0.008162f
C231 B.n186 VSUBS 0.008162f
C232 B.n187 VSUBS 0.008162f
C233 B.n188 VSUBS 0.008162f
C234 B.n189 VSUBS 0.008162f
C235 B.n190 VSUBS 0.008162f
C236 B.n191 VSUBS 0.008162f
C237 B.n192 VSUBS 0.008162f
C238 B.n193 VSUBS 0.008162f
C239 B.n194 VSUBS 0.008162f
C240 B.n195 VSUBS 0.008162f
C241 B.n196 VSUBS 0.019332f
C242 B.n197 VSUBS 0.018838f
C243 B.n198 VSUBS 0.019803f
C244 B.n199 VSUBS 0.008162f
C245 B.n200 VSUBS 0.008162f
C246 B.n201 VSUBS 0.008162f
C247 B.n202 VSUBS 0.008162f
C248 B.n203 VSUBS 0.008162f
C249 B.n204 VSUBS 0.008162f
C250 B.n205 VSUBS 0.008162f
C251 B.n206 VSUBS 0.008162f
C252 B.n207 VSUBS 0.008162f
C253 B.n208 VSUBS 0.008162f
C254 B.n209 VSUBS 0.008162f
C255 B.n210 VSUBS 0.008162f
C256 B.n211 VSUBS 0.008162f
C257 B.n212 VSUBS 0.008162f
C258 B.n213 VSUBS 0.008162f
C259 B.n214 VSUBS 0.008162f
C260 B.n215 VSUBS 0.008162f
C261 B.n216 VSUBS 0.008162f
C262 B.n217 VSUBS 0.008162f
C263 B.n218 VSUBS 0.008162f
C264 B.n219 VSUBS 0.007442f
C265 B.n220 VSUBS 0.018911f
C266 B.n221 VSUBS 0.004801f
C267 B.n222 VSUBS 0.008162f
C268 B.n223 VSUBS 0.008162f
C269 B.n224 VSUBS 0.008162f
C270 B.n225 VSUBS 0.008162f
C271 B.n226 VSUBS 0.008162f
C272 B.n227 VSUBS 0.008162f
C273 B.n228 VSUBS 0.008162f
C274 B.n229 VSUBS 0.008162f
C275 B.n230 VSUBS 0.008162f
C276 B.n231 VSUBS 0.008162f
C277 B.n232 VSUBS 0.008162f
C278 B.n233 VSUBS 0.008162f
C279 B.n234 VSUBS 0.004801f
C280 B.n235 VSUBS 0.008162f
C281 B.n236 VSUBS 0.008162f
C282 B.n237 VSUBS 0.007442f
C283 B.n238 VSUBS 0.008162f
C284 B.n239 VSUBS 0.008162f
C285 B.n240 VSUBS 0.008162f
C286 B.n241 VSUBS 0.008162f
C287 B.n242 VSUBS 0.008162f
C288 B.n243 VSUBS 0.008162f
C289 B.n244 VSUBS 0.008162f
C290 B.n245 VSUBS 0.008162f
C291 B.n246 VSUBS 0.008162f
C292 B.n247 VSUBS 0.008162f
C293 B.n248 VSUBS 0.008162f
C294 B.n249 VSUBS 0.008162f
C295 B.n250 VSUBS 0.008162f
C296 B.n251 VSUBS 0.008162f
C297 B.n252 VSUBS 0.008162f
C298 B.n253 VSUBS 0.008162f
C299 B.n254 VSUBS 0.008162f
C300 B.n255 VSUBS 0.008162f
C301 B.n256 VSUBS 0.008162f
C302 B.n257 VSUBS 0.019803f
C303 B.n258 VSUBS 0.019803f
C304 B.n259 VSUBS 0.018367f
C305 B.n260 VSUBS 0.008162f
C306 B.n261 VSUBS 0.008162f
C307 B.n262 VSUBS 0.008162f
C308 B.n263 VSUBS 0.008162f
C309 B.n264 VSUBS 0.008162f
C310 B.n265 VSUBS 0.008162f
C311 B.n266 VSUBS 0.008162f
C312 B.n267 VSUBS 0.008162f
C313 B.n268 VSUBS 0.008162f
C314 B.n269 VSUBS 0.008162f
C315 B.n270 VSUBS 0.008162f
C316 B.n271 VSUBS 0.008162f
C317 B.n272 VSUBS 0.008162f
C318 B.n273 VSUBS 0.008162f
C319 B.n274 VSUBS 0.008162f
C320 B.n275 VSUBS 0.008162f
C321 B.n276 VSUBS 0.008162f
C322 B.n277 VSUBS 0.008162f
C323 B.n278 VSUBS 0.008162f
C324 B.n279 VSUBS 0.018482f
C325 VDD1.t0 VSUBS 0.2923f
C326 VDD1.t1 VSUBS 0.412725f
C327 VTAIL.t1 VSUBS 0.324694f
C328 VTAIL.n0 VSUBS 0.891584f
C329 VTAIL.t0 VSUBS 0.324695f
C330 VTAIL.n1 VSUBS 0.900082f
C331 VTAIL.t2 VSUBS 0.324694f
C332 VTAIL.n2 VSUBS 0.850529f
C333 VTAIL.t3 VSUBS 0.324694f
C334 VTAIL.n3 VSUBS 0.802849f
C335 VP.t1 VSUBS 0.33646f
C336 VP.t0 VSUBS 0.245611f
C337 VP.n0 VSUBS 2.20769f
.ends

