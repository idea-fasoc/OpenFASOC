* NGSPICE file created from opamp_sample_0008.ext - technology: sky130A

.subckt opamp_sample_0008 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VDD.t128 VDD.t126 VDD.t127 VDD.t120 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X1 VOUT.t41 CS_BIAS.t24 GND.t79 GND.t65 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X2 GND.t78 CS_BIAS.t25 VOUT.t40 GND.t53 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0.6204 ps=4.09 w=3.76 l=5.93
X3 a_n6364_n172.t22 VN.t5 a_n18960_7900.t17 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X4 a_n7729_8946.t17 a_n7651_8750.t30 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X5 VP.t4 GND.t169 GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X6 a_n7729_8946.t16 a_n7651_8750.t31 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X7 a_n7651_8750.t13 a_n7651_8750.t12 a_n7729_8946.t9 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X8 DIFFPAIR_BIAS.t11 DIFFPAIR_BIAS.t10 GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X9 DIFFPAIR_BIAS.t9 DIFFPAIR_BIAS.t8 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X10 a_n6364_n172.t21 VN.t6 a_n18960_7900.t15 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X11 a_n6364_n172.t1 VP.t5 a_n7651_8750.t0 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X12 VP.t3 GND.t166 GND.t168 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 a_n8793_8946# a_n8793_8946# a_n8793_8946# VDD.t140 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=3.198 ps=17.96 w=4.1 l=3.9
X14 GND.t165 GND.t162 GND.t164 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0 ps=0 w=2.48 l=3.75
X15 a_n7651_8750.t11 a_n7651_8750.t10 a_n7729_8946.t8 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X16 VDD.t44 a_n7651_8750.t32 a_n5900_7192.t18 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X17 GND.t77 CS_BIAS.t26 VOUT.t39 GND.t55 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X18 GND.t161 GND.t159 GND.t160 GND.t91 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X19 a_n7651_8750.t23 a_n7651_8750.t22 a_n7729_8946.t7 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X20 VOUT.t44 a_n18960_7900.t20 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=1.9188 ps=10.62 w=4.92 l=5.29
X21 GND.t76 CS_BIAS.t27 VOUT.t38 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0.6204 ps=4.09 w=3.76 l=5.93
X22 VDD.t125 VDD.t123 VDD.t124 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X23 VDD.t122 VDD.t119 VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X24 CS_BIAS.t21 CS_BIAS.t20 GND.t75 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X25 a_n6364_n172.t12 VP.t6 a_n7651_8750.t7 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X26 GND.t74 CS_BIAS.t14 CS_BIAS.t15 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0.6204 ps=4.09 w=3.76 l=5.93
X27 VOUT.t37 CS_BIAS.t28 GND.t73 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=1.4664 ps=8.3 w=3.76 l=5.93
X28 GND.t72 CS_BIAS.t4 CS_BIAS.t5 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X29 a_n18960_7900.t18 a_n7651_8750.t33 a_n5900_7192.t10 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X30 VOUT.t51 a_n18960_7900.t21 VDD.t141 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X31 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X32 a_n6364_n172.t20 VN.t7 a_n18960_7900.t16 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X33 a_n7651_8750.t2 VP.t7 a_n6364_n172.t4 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=5.88
X34 VOUT.t8 a_n18960_7900.t22 VDD.t39 VDD.t37 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0.8118 ps=5.25 w=4.92 l=5.29
X35 VOUT.t42 a_n18960_7900.t23 VDD.t66 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X36 VDD.t10 a_n7651_8750.t34 a_n7729_8946.t15 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X37 VN.t4 GND.t156 GND.t158 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X38 GND.t71 CS_BIAS.t0 CS_BIAS.t1 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X39 GND.t70 CS_BIAS.t29 VOUT.t36 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X40 GND.t155 GND.t153 VP.t2 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X41 a_n6364_n172.t9 DIFFPAIR_BIAS.t12 GND.t20 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X42 VDD.t56 a_n18960_7900.t24 VOUT.t15 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X43 VDD.t118 VDD.t116 VDD.t117 VDD.t74 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X44 CS_BIAS.t9 CS_BIAS.t8 GND.t59 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=1.4664 ps=8.3 w=3.76 l=5.93
X45 VOUT.t52 a_n5900_7192.t0 sky130_fd_pr__cap_mim_m3_1 l=5.72 w=6.01
X46 VDD.t115 VDD.t113 VDD.t114 VDD.t78 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X47 VOUT.t53 a_n5900_7192.t0 sky130_fd_pr__cap_mim_m3_1 l=5.72 w=6.01
X48 GND.t152 GND.t150 GND.t151 GND.t101 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X49 a_n18960_7900.t10 VN.t8 a_n6364_n172.t19 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=5.88
X50 VDD.t24 a_n18960_7900.t25 VOUT.t4 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X51 a_n7729_8946.t6 a_n7651_8750.t18 a_n7651_8750.t19 VDD.t36 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X52 GND.t68 CS_BIAS.t30 VOUT.t35 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X53 VDD.t112 VDD.t110 VDD.t111 VDD.t90 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X54 a_n18960_7900.t11 VN.t9 a_n6364_n172.t18 GND.t31 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=5.88
X55 GND.t69 CS_BIAS.t31 VOUT.t34 GND.t55 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X56 VOUT.t33 CS_BIAS.t32 GND.t67 GND.t65 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X57 GND.t149 GND.t147 GND.t148 GND.t114 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X58 a_n7729_8946.t14 a_n7651_8750.t35 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X59 a_n7729_8946.t13 a_n7651_8750.t36 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X60 CS_BIAS.t7 CS_BIAS.t6 GND.t66 GND.t65 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X61 a_n5900_7192.t9 a_n7651_8750.t37 a_n18960_7900.t5 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X62 VDD.t109 VDD.t107 VDD.t108 VDD.t94 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X63 GND.t64 CS_BIAS.t33 VOUT.t32 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0.6204 ps=4.09 w=3.76 l=5.93
X64 VOUT.t11 a_n18960_7900.t26 VDD.t49 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X65 CS_BIAS.t13 CS_BIAS.t12 GND.t62 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X66 GND.t61 CS_BIAS.t34 VOUT.t31 GND.t53 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0.6204 ps=4.09 w=3.76 l=5.93
X67 a_n18960_7900.t4 a_n7651_8750.t38 a_n5900_7192.t8 VDD.t36 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X68 a_n7729_8946.t5 a_n7651_8750.t16 a_n7651_8750.t17 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X69 GND.t60 CS_BIAS.t22 CS_BIAS.t23 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X70 a_n7651_8750.t9 VP.t8 a_n6364_n172.t24 GND.t31 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=5.88
X71 GND.t146 GND.t144 GND.t145 GND.t135 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=5.88
X72 VOUT.t30 CS_BIAS.t35 GND.t58 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X73 VDD.t6 a_n18960_7900.t27 VOUT.t0 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X74 GND.t143 GND.t141 VP.t1 GND.t142 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X75 CS_BIAS.t11 CS_BIAS.t10 GND.t57 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=1.4664 ps=8.3 w=3.76 l=5.93
X76 GND.t140 GND.t138 GND.t139 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=5.88
X77 VDD.t71 a_n18960_7900.t28 VOUT.t45 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X78 a_n6364_n172.t8 DIFFPAIR_BIAS.t13 GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X79 GND.t56 CS_BIAS.t16 CS_BIAS.t17 GND.t55 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X80 VDD.t3 a_n7651_8750.t39 a_n5900_7192.t17 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X81 a_n6364_n172.t25 DIFFPAIR_BIAS.t14 GND.t173 GND.t172 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X82 GND.t137 GND.t134 GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=5.88
X83 VOUT.t9 a_n18960_7900.t29 VDD.t46 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=1.9188 ps=10.62 w=4.92 l=5.29
X84 GND.t133 GND.t131 GND.t132 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X85 VOUT.t47 a_n18960_7900.t30 VDD.t129 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=1.9188 ps=10.62 w=4.92 l=5.29
X86 a_n6364_n172.t2 DIFFPAIR_BIAS.t15 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X87 GND.t130 GND.t128 GND.t129 GND.t114 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X88 a_n7651_8750.t5 VP.t9 a_n6364_n172.t7 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X89 GND.t127 GND.t124 GND.t126 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=5.88
X90 VDD.t106 VDD.t103 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X91 a_n5900_7192.t16 a_n7651_8750.t40 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X92 VDD.t102 VDD.t100 VDD.t101 VDD.t86 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X93 a_n18960_7900.t6 a_n7651_8750.t41 a_n5900_7192.t7 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X94 GND.t123 GND.t120 GND.t122 GND.t121 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0 ps=0 w=2.48 l=3.75
X95 VDD.t99 VDD.t97 VDD.t98 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X96 GND.t54 CS_BIAS.t2 CS_BIAS.t3 GND.t53 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0.6204 ps=4.09 w=3.76 l=5.93
X97 VDD.t27 a_n18960_7900.t31 VOUT.t5 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X98 CS_BIAS.t19 CS_BIAS.t18 GND.t52 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X99 a_n18960_7900.t12 VN.t10 a_n6364_n172.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X100 a_n18960_7900.t14 VN.t11 a_n6364_n172.t16 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=5.88
X101 VOUT.t29 CS_BIAS.t36 GND.t51 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=1.4664 ps=8.3 w=3.76 l=5.93
X102 a_n5900_7192.t6 a_n7651_8750.t42 a_n18960_7900.t7 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X103 a_n5900_7192.t5 a_n7651_8750.t43 a_n18960_7900.t1 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X104 VOUT.t13 a_n18960_7900.t32 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X105 GND.t116 GND.t113 GND.t115 GND.t114 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X106 VOUT.t28 CS_BIAS.t37 GND.t50 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=1.4664 ps=8.3 w=3.76 l=5.93
X107 VOUT.t43 a_n18960_7900.t33 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X108 a_n7729_8946.t4 a_n7651_8750.t14 a_n7651_8750.t15 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X109 a_n7651_8750.t8 VP.t10 a_n6364_n172.t23 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=5.88
X110 VOUT.t10 a_n18960_7900.t34 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X111 GND.t48 CS_BIAS.t38 VOUT.t27 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X112 a_n18960_7900.t0 a_n7651_8750.t44 a_n5900_7192.t4 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X113 VDD.t72 a_n18960_7900.t35 VOUT.t46 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X114 GND.t47 CS_BIAS.t39 VOUT.t26 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X115 VOUT.t25 CS_BIAS.t40 GND.t45 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=1.4664 ps=8.3 w=3.76 l=5.93
X116 VDD.t65 a_n18960_7900.t36 VOUT.t17 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X117 a_n7651_8750.t29 a_n7651_8750.t28 a_n7729_8946.t3 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X118 GND.t112 GND.t110 GND.t111 GND.t101 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X119 a_n7651_8750.t6 VP.t11 a_n6364_n172.t10 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=5.88
X120 VN.t3 GND.t117 GND.t119 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X121 VDD.t60 a_n7651_8750.t45 a_n7729_8946.t12 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X122 VOUT.t50 a_n18960_7900.t37 VDD.t139 VDD.t54 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0.8118 ps=5.25 w=4.92 l=5.29
X123 VDD.t96 VDD.t93 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X124 VOUT.t24 CS_BIAS.t41 GND.t43 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X125 VOUT.t2 a_n18960_7900.t38 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X126 GND.t109 GND.t107 VN.t2 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X127 VDD.t31 a_n7651_8750.t46 a_n7729_8946.t11 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X128 a_n18960_7900.t9 VN.t12 a_n6364_n172.t15 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=5.88
X129 VDD.t34 a_n7651_8750.t47 a_n7729_8946.t10 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X130 VDD.t35 a_n18960_7900.t39 VOUT.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X131 GND.t89 GND.t87 VP.t0 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X132 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X133 a_n18960_7900.t13 VN.t13 a_n6364_n172.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X134 VDD.t64 a_n18960_7900.t40 VOUT.t16 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X135 a_n6364_n172.t11 DIFFPAIR_BIAS.t16 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X136 GND.t106 GND.t104 GND.t105 GND.t91 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X137 a_n5900_7192.t15 a_n7651_8750.t48 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X138 VOUT.t23 CS_BIAS.t42 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X139 VOUT.t1 a_n18960_7900.t41 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=1.9188 ps=10.62 w=4.92 l=5.29
X140 VDD.t92 VDD.t89 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X141 GND.t40 CS_BIAS.t43 VOUT.t22 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X142 VOUT.t21 CS_BIAS.t44 GND.t38 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X143 VDD.t88 VDD.t85 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X144 a_n6364_n172.t13 VN.t14 a_n18960_7900.t8 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X145 a_n5900_7192.t14 a_n7651_8750.t49 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X146 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X147 GND.t103 GND.t100 GND.t102 GND.t101 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X148 a_n7651_8750.t4 VP.t12 a_n6364_n172.t6 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X149 VDD.t84 VDD.t81 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=5.29
X150 GND.t99 GND.t97 VN.t1 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X151 a_n7729_8946.t2 a_n7651_8750.t26 a_n7651_8750.t27 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X152 VDD.t138 a_n18960_7900.t42 VOUT.t49 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X153 a_7857_8946# a_7857_8946# a_7857_8946# VDD.t42 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=3.198 ps=17.96 w=4.1 l=3.9
X154 GND.t37 CS_BIAS.t45 VOUT.t20 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X155 VOUT.t19 CS_BIAS.t46 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X156 a_n18960_7900.t3 a_n7651_8750.t50 a_n5900_7192.t3 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X157 a_n6364_n172.t5 VP.t13 a_n7651_8750.t3 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X158 GND.t96 GND.t94 GND.t95 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X159 a_n5900_7192.t2 a_n7651_8750.t51 a_n18960_7900.t19 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X160 VDD.t1 a_n7651_8750.t52 a_n5900_7192.t13 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X161 VOUT.t48 a_n18960_7900.t43 VDD.t133 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X162 VDD.t80 VDD.t77 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X163 VDD.t76 VDD.t73 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=3.9
X164 VOUT.t7 a_n18960_7900.t44 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0.8118 ps=5.25 w=4.92 l=5.29
X165 VDD.t58 a_n7651_8750.t53 a_n5900_7192.t12 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=3.9
X166 a_n6364_n172.t0 DIFFPAIR_BIAS.t17 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X167 VDD.t22 a_n18960_7900.t45 VOUT.t3 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X168 GND.t93 GND.t90 GND.t92 GND.t91 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X169 GND.t86 GND.t83 GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=5.93
X170 VOUT.t18 CS_BIAS.t47 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6204 pd=4.09 as=0.6204 ps=4.09 w=3.76 l=5.93
X171 a_n18960_7900.t2 a_n7651_8750.t54 a_n5900_7192.t1 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X172 VDD.t51 a_n18960_7900.t46 VOUT.t12 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.8118 pd=5.25 as=0.8118 ps=5.25 w=4.92 l=5.29
X173 GND.t82 GND.t80 VN.t0 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X174 a_n7729_8946.t1 a_n7651_8750.t24 a_n7651_8750.t25 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=3.9
X175 a_n7729_8946.t0 a_n7651_8750.t20 a_n7651_8750.t21 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
X176 VOUT.t14 a_n18960_7900.t47 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=1.9188 pd=10.62 as=0.8118 ps=5.25 w=4.92 l=5.29
X177 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t30 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.9672 pd=5.74 as=0.9672 ps=5.74 w=2.48 l=3.75
X178 a_n6364_n172.t3 VP.t14 a_n7651_8750.t1 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=5.88
X179 a_n5900_7192.t11 a_n7651_8750.t55 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=3.9
R0 VDD.n215 VDD.n177 466.829
R1 VDD.n4048 VDD.n179 466.829
R2 VDD.n513 VDD.n467 466.829
R3 VDD.n603 VDD.n465 466.829
R4 VDD.n2521 VDD.n1243 466.829
R5 VDD.n2524 VDD.n2523 466.829
R6 VDD.n1640 VDD.n1620 466.829
R7 VDD.n1731 VDD.n1622 466.829
R8 VDD.n3296 VDD.n903 304.39
R9 VDD.n3717 VDD.n489 304.39
R10 VDD.n3681 VDD.n486 304.39
R11 VDD.n3170 VDD.n2977 304.39
R12 VDD.n3660 VDD.n487 304.39
R13 VDD.n3720 VDD.n3719 304.39
R14 VDD.n3253 VDD.n2978 304.39
R15 VDD.n3294 VDD.n2979 304.39
R16 VDD.n2902 VDD.n2901 304.39
R17 VDD.n2973 VDD.n925 304.39
R18 VDD.n2483 VDD.n2482 304.39
R19 VDD.n2160 VDD.n1213 304.39
R20 VDD.n2963 VDD.n933 304.39
R21 VDD.n2924 VDD.n2923 304.39
R22 VDD.n2329 VDD.n1228 304.39
R23 VDD.n2590 VDD.n1217 304.39
R24 VDD.n2308 VDD.t126 234.756
R25 VDD.n935 VDD.t116 234.756
R26 VDD.n2988 VDD.t89 234.756
R27 VDD.n614 VDD.t77 234.756
R28 VDD.n3124 VDD.t110 234.756
R29 VDD.n479 VDD.t113 234.756
R30 VDD.n2179 VDD.t119 234.756
R31 VDD.n2863 VDD.t73 234.756
R32 VDD.n1259 VDD.t81 232.611
R33 VDD.n1281 VDD.t97 232.611
R34 VDD.n1681 VDD.t100 232.611
R35 VDD.n1708 VDD.t85 232.611
R36 VDD.n527 VDD.t93 232.611
R37 VDD.n545 VDD.t107 232.611
R38 VDD.n195 VDD.t123 232.611
R39 VDD.n205 VDD.t103 232.611
R40 VDD.n1259 VDD.t83 226.718
R41 VDD.n1281 VDD.t98 226.718
R42 VDD.n1681 VDD.t102 226.718
R43 VDD.n1708 VDD.t88 226.718
R44 VDD.n527 VDD.t96 226.718
R45 VDD.n545 VDD.t109 226.718
R46 VDD.n195 VDD.t124 226.718
R47 VDD.n205 VDD.t105 226.718
R48 VDD.n1308 VDD.t42 221.085
R49 VDD.n601 VDD.t140 221.085
R50 VDD.n2308 VDD.t128 201.472
R51 VDD.n935 VDD.t117 201.472
R52 VDD.n2988 VDD.t92 201.472
R53 VDD.n614 VDD.t79 201.472
R54 VDD.n3124 VDD.t112 201.472
R55 VDD.n479 VDD.t114 201.472
R56 VDD.n2179 VDD.t122 201.472
R57 VDD.n2863 VDD.t75 201.472
R58 VDD.t42 VDD.t28 185.81
R59 VDD.t140 VDD.t9 185.81
R60 VDD.n2903 VDD.n2902 185
R61 VDD.n2902 VDD.n904 185
R62 VDD.n2904 VDD.n931 185
R63 VDD.n2968 VDD.n931 185
R64 VDD.n2906 VDD.n2905 185
R65 VDD.n2905 VDD.n929 185
R66 VDD.n2907 VDD.n941 185
R67 VDD.n2917 VDD.n941 185
R68 VDD.n2908 VDD.n949 185
R69 VDD.n949 VDD.n939 185
R70 VDD.n2910 VDD.n2909 185
R71 VDD.n2911 VDD.n2910 185
R72 VDD.n2862 VDD.n948 185
R73 VDD.n948 VDD.n945 185
R74 VDD.n2861 VDD.n2860 185
R75 VDD.n2860 VDD.n2859 185
R76 VDD.n951 VDD.n950 185
R77 VDD.n960 VDD.n951 185
R78 VDD.n2852 VDD.n2851 185
R79 VDD.n2853 VDD.n2852 185
R80 VDD.n2850 VDD.n961 185
R81 VDD.n961 VDD.n957 185
R82 VDD.n2849 VDD.n2848 185
R83 VDD.n2848 VDD.n2847 185
R84 VDD.n963 VDD.n962 185
R85 VDD.n964 VDD.n963 185
R86 VDD.n2840 VDD.n2839 185
R87 VDD.n2841 VDD.n2840 185
R88 VDD.n2838 VDD.n973 185
R89 VDD.n973 VDD.n970 185
R90 VDD.n2837 VDD.n2836 185
R91 VDD.n2836 VDD.n2835 185
R92 VDD.n975 VDD.n974 185
R93 VDD.n976 VDD.n975 185
R94 VDD.n2828 VDD.n2827 185
R95 VDD.n2829 VDD.n2828 185
R96 VDD.n2826 VDD.n985 185
R97 VDD.n985 VDD.n982 185
R98 VDD.n2825 VDD.n2824 185
R99 VDD.n2824 VDD.n2823 185
R100 VDD.n987 VDD.n986 185
R101 VDD.n988 VDD.n987 185
R102 VDD.n2816 VDD.n2815 185
R103 VDD.n2817 VDD.n2816 185
R104 VDD.n2814 VDD.n997 185
R105 VDD.n997 VDD.n994 185
R106 VDD.n2813 VDD.n2812 185
R107 VDD.n2812 VDD.n2811 185
R108 VDD.n999 VDD.n998 185
R109 VDD.n1008 VDD.n999 185
R110 VDD.n2804 VDD.n2803 185
R111 VDD.n2805 VDD.n2804 185
R112 VDD.n2802 VDD.n1009 185
R113 VDD.n1009 VDD.n1005 185
R114 VDD.n2801 VDD.n2800 185
R115 VDD.n2800 VDD.n2799 185
R116 VDD.n1011 VDD.n1010 185
R117 VDD.n1012 VDD.n1011 185
R118 VDD.n2792 VDD.n2791 185
R119 VDD.n2793 VDD.n2792 185
R120 VDD.n2790 VDD.n1021 185
R121 VDD.n1021 VDD.n1018 185
R122 VDD.n2789 VDD.n2788 185
R123 VDD.n2788 VDD.n2787 185
R124 VDD.n1023 VDD.n1022 185
R125 VDD.n1032 VDD.n1023 185
R126 VDD.n2780 VDD.n2779 185
R127 VDD.n2781 VDD.n2780 185
R128 VDD.n2778 VDD.n1033 185
R129 VDD.n1033 VDD.n1029 185
R130 VDD.n2777 VDD.n2776 185
R131 VDD.n2776 VDD.n2775 185
R132 VDD.n1035 VDD.n1034 185
R133 VDD.n1044 VDD.n1035 185
R134 VDD.n2768 VDD.n2767 185
R135 VDD.n2769 VDD.n2768 185
R136 VDD.n2766 VDD.n1045 185
R137 VDD.n1045 VDD.n1041 185
R138 VDD.n2765 VDD.n2764 185
R139 VDD.n2764 VDD.n2763 185
R140 VDD.n1047 VDD.n1046 185
R141 VDD.n1048 VDD.n1047 185
R142 VDD.n2756 VDD.n2755 185
R143 VDD.n2757 VDD.n2756 185
R144 VDD.n2754 VDD.n1057 185
R145 VDD.n1057 VDD.n1054 185
R146 VDD.n2753 VDD.n2752 185
R147 VDD.n2752 VDD.n2751 185
R148 VDD.n1059 VDD.n1058 185
R149 VDD.n1068 VDD.n1059 185
R150 VDD.n2744 VDD.n2743 185
R151 VDD.n2745 VDD.n2744 185
R152 VDD.n2742 VDD.n1069 185
R153 VDD.n1069 VDD.n1065 185
R154 VDD.n2741 VDD.n2740 185
R155 VDD.n2740 VDD.n2739 185
R156 VDD.n1071 VDD.n1070 185
R157 VDD.t25 VDD.n1071 185
R158 VDD.n2732 VDD.n2731 185
R159 VDD.n2733 VDD.n2732 185
R160 VDD.n2730 VDD.n1080 185
R161 VDD.n1080 VDD.n1077 185
R162 VDD.n2729 VDD.n2728 185
R163 VDD.n2728 VDD.n2727 185
R164 VDD.n1082 VDD.n1081 185
R165 VDD.n1083 VDD.n1082 185
R166 VDD.n2720 VDD.n2719 185
R167 VDD.n2721 VDD.n2720 185
R168 VDD.n2718 VDD.n1092 185
R169 VDD.n1092 VDD.n1089 185
R170 VDD.n2717 VDD.n2716 185
R171 VDD.n2716 VDD.n2715 185
R172 VDD.n1094 VDD.n1093 185
R173 VDD.n1095 VDD.n1094 185
R174 VDD.n2708 VDD.n2707 185
R175 VDD.n2709 VDD.n2708 185
R176 VDD.n2706 VDD.n1104 185
R177 VDD.n1104 VDD.n1101 185
R178 VDD.n2705 VDD.n2704 185
R179 VDD.n2704 VDD.n2703 185
R180 VDD.n1106 VDD.n1105 185
R181 VDD.n1107 VDD.n1106 185
R182 VDD.n2696 VDD.n2695 185
R183 VDD.n2697 VDD.n2696 185
R184 VDD.n2694 VDD.n1116 185
R185 VDD.n1116 VDD.n1113 185
R186 VDD.n2693 VDD.n2692 185
R187 VDD.n2692 VDD.n2691 185
R188 VDD.n1118 VDD.n1117 185
R189 VDD.n1119 VDD.n1118 185
R190 VDD.n2684 VDD.n2683 185
R191 VDD.n2685 VDD.n2684 185
R192 VDD.n2682 VDD.n1128 185
R193 VDD.n1128 VDD.n1125 185
R194 VDD.n2681 VDD.n2680 185
R195 VDD.n2680 VDD.n2679 185
R196 VDD.n1130 VDD.n1129 185
R197 VDD.n1131 VDD.n1130 185
R198 VDD.n2672 VDD.n2671 185
R199 VDD.n2673 VDD.n2672 185
R200 VDD.n2670 VDD.n1140 185
R201 VDD.n1140 VDD.n1137 185
R202 VDD.n2669 VDD.n2668 185
R203 VDD.n2668 VDD.n2667 185
R204 VDD.n1142 VDD.n1141 185
R205 VDD.n1143 VDD.n1142 185
R206 VDD.n2660 VDD.n2659 185
R207 VDD.n2661 VDD.n2660 185
R208 VDD.n2658 VDD.n1152 185
R209 VDD.n1152 VDD.n1149 185
R210 VDD.n2657 VDD.n2656 185
R211 VDD.n2656 VDD.n2655 185
R212 VDD.n1154 VDD.n1153 185
R213 VDD.n1155 VDD.n1154 185
R214 VDD.n2648 VDD.n2647 185
R215 VDD.n2649 VDD.n2648 185
R216 VDD.n2646 VDD.n1164 185
R217 VDD.n1164 VDD.n1161 185
R218 VDD.n2645 VDD.n2644 185
R219 VDD.n2644 VDD.n2643 185
R220 VDD.n1166 VDD.n1165 185
R221 VDD.n1167 VDD.n1166 185
R222 VDD.n2636 VDD.n2635 185
R223 VDD.n2637 VDD.n2636 185
R224 VDD.n2634 VDD.n1176 185
R225 VDD.n1176 VDD.n1173 185
R226 VDD.n2633 VDD.n2632 185
R227 VDD.n2632 VDD.n2631 185
R228 VDD.n1178 VDD.n1177 185
R229 VDD.n1179 VDD.n1178 185
R230 VDD.n2624 VDD.n2623 185
R231 VDD.n2625 VDD.n2624 185
R232 VDD.n2622 VDD.n1188 185
R233 VDD.n1188 VDD.n1185 185
R234 VDD.n2621 VDD.n2620 185
R235 VDD.n2620 VDD.n2619 185
R236 VDD.n1190 VDD.n1189 185
R237 VDD.n2468 VDD.n1190 185
R238 VDD.n2612 VDD.n2611 185
R239 VDD.n2613 VDD.n2612 185
R240 VDD.n2610 VDD.n1199 185
R241 VDD.n1199 VDD.n1196 185
R242 VDD.n2609 VDD.n2608 185
R243 VDD.n2608 VDD.n2607 185
R244 VDD.n1201 VDD.n1200 185
R245 VDD.n1202 VDD.n1201 185
R246 VDD.n2600 VDD.n2599 185
R247 VDD.n2601 VDD.n2600 185
R248 VDD.n2598 VDD.n1211 185
R249 VDD.n1211 VDD.n1208 185
R250 VDD.n2597 VDD.n2596 185
R251 VDD.n2596 VDD.n2595 185
R252 VDD.n1213 VDD.n1212 185
R253 VDD.n1214 VDD.n1213 185
R254 VDD.n2161 VDD.n2160 185
R255 VDD.n2163 VDD.n2162 185
R256 VDD.n2165 VDD.n2164 185
R257 VDD.n2167 VDD.n2166 185
R258 VDD.n2169 VDD.n2168 185
R259 VDD.n2171 VDD.n2170 185
R260 VDD.n2173 VDD.n2172 185
R261 VDD.n2175 VDD.n2174 185
R262 VDD.n2177 VDD.n2176 185
R263 VDD.n2502 VDD.n2178 185
R264 VDD.n2504 VDD.n2503 185
R265 VDD.n2501 VDD.n2500 185
R266 VDD.n2499 VDD.n2498 185
R267 VDD.n2497 VDD.n2496 185
R268 VDD.n2495 VDD.n2494 185
R269 VDD.n2493 VDD.n2492 185
R270 VDD.n2491 VDD.n2490 185
R271 VDD.n2488 VDD.n2487 185
R272 VDD.n2486 VDD.n2485 185
R273 VDD.n2484 VDD.n2483 185
R274 VDD.n2973 VDD.n2972 185
R275 VDD.n926 VDD.n924 185
R276 VDD.n2866 VDD.n2865 185
R277 VDD.n2869 VDD.n2868 185
R278 VDD.n2871 VDD.n2870 185
R279 VDD.n2873 VDD.n2872 185
R280 VDD.n2875 VDD.n2874 185
R281 VDD.n2877 VDD.n2876 185
R282 VDD.n2879 VDD.n2878 185
R283 VDD.n2881 VDD.n2880 185
R284 VDD.n2883 VDD.n2882 185
R285 VDD.n2885 VDD.n2884 185
R286 VDD.n2887 VDD.n2886 185
R287 VDD.n2889 VDD.n2888 185
R288 VDD.n2891 VDD.n2890 185
R289 VDD.n2893 VDD.n2892 185
R290 VDD.n2895 VDD.n2894 185
R291 VDD.n2897 VDD.n2896 185
R292 VDD.n2899 VDD.n2898 185
R293 VDD.n2901 VDD.n2900 185
R294 VDD.n2971 VDD.n925 185
R295 VDD.n925 VDD.n904 185
R296 VDD.n2970 VDD.n2969 185
R297 VDD.n2969 VDD.n2968 185
R298 VDD.n928 VDD.n927 185
R299 VDD.n929 VDD.n928 185
R300 VDD.n2181 VDD.n940 185
R301 VDD.n2917 VDD.n940 185
R302 VDD.n2183 VDD.n2182 185
R303 VDD.n2182 VDD.n939 185
R304 VDD.n2184 VDD.n947 185
R305 VDD.n2911 VDD.n947 185
R306 VDD.n2186 VDD.n2185 185
R307 VDD.n2185 VDD.n945 185
R308 VDD.n2187 VDD.n953 185
R309 VDD.n2859 VDD.n953 185
R310 VDD.n2189 VDD.n2188 185
R311 VDD.n2188 VDD.n960 185
R312 VDD.n2190 VDD.n959 185
R313 VDD.n2853 VDD.n959 185
R314 VDD.n2192 VDD.n2191 185
R315 VDD.n2191 VDD.n957 185
R316 VDD.n2193 VDD.n966 185
R317 VDD.n2847 VDD.n966 185
R318 VDD.n2195 VDD.n2194 185
R319 VDD.n2194 VDD.n964 185
R320 VDD.n2196 VDD.n972 185
R321 VDD.n2841 VDD.n972 185
R322 VDD.n2198 VDD.n2197 185
R323 VDD.n2197 VDD.n970 185
R324 VDD.n2199 VDD.n978 185
R325 VDD.n2835 VDD.n978 185
R326 VDD.n2201 VDD.n2200 185
R327 VDD.n2200 VDD.n976 185
R328 VDD.n2202 VDD.n984 185
R329 VDD.n2829 VDD.n984 185
R330 VDD.n2204 VDD.n2203 185
R331 VDD.n2203 VDD.n982 185
R332 VDD.n2205 VDD.n990 185
R333 VDD.n2823 VDD.n990 185
R334 VDD.n2207 VDD.n2206 185
R335 VDD.n2206 VDD.n988 185
R336 VDD.n2208 VDD.n996 185
R337 VDD.n2817 VDD.n996 185
R338 VDD.n2210 VDD.n2209 185
R339 VDD.n2209 VDD.n994 185
R340 VDD.n2211 VDD.n1001 185
R341 VDD.n2811 VDD.n1001 185
R342 VDD.n2213 VDD.n2212 185
R343 VDD.n2212 VDD.n1008 185
R344 VDD.n2214 VDD.n1007 185
R345 VDD.n2805 VDD.n1007 185
R346 VDD.n2216 VDD.n2215 185
R347 VDD.n2215 VDD.n1005 185
R348 VDD.n2217 VDD.n1014 185
R349 VDD.n2799 VDD.n1014 185
R350 VDD.n2219 VDD.n2218 185
R351 VDD.n2218 VDD.n1012 185
R352 VDD.n2220 VDD.n1020 185
R353 VDD.n2793 VDD.n1020 185
R354 VDD.n2222 VDD.n2221 185
R355 VDD.n2221 VDD.n1018 185
R356 VDD.n2223 VDD.n1025 185
R357 VDD.n2787 VDD.n1025 185
R358 VDD.n2225 VDD.n2224 185
R359 VDD.n2224 VDD.n1032 185
R360 VDD.n2226 VDD.n1031 185
R361 VDD.n2781 VDD.n1031 185
R362 VDD.n2228 VDD.n2227 185
R363 VDD.n2227 VDD.n1029 185
R364 VDD.n2229 VDD.n1037 185
R365 VDD.n2775 VDD.n1037 185
R366 VDD.n2231 VDD.n2230 185
R367 VDD.n2230 VDD.n1044 185
R368 VDD.n2232 VDD.n1043 185
R369 VDD.n2769 VDD.n1043 185
R370 VDD.n2234 VDD.n2233 185
R371 VDD.n2233 VDD.n1041 185
R372 VDD.n2235 VDD.n1050 185
R373 VDD.n2763 VDD.n1050 185
R374 VDD.n2237 VDD.n2236 185
R375 VDD.n2236 VDD.n1048 185
R376 VDD.n2238 VDD.n1056 185
R377 VDD.n2757 VDD.n1056 185
R378 VDD.n2240 VDD.n2239 185
R379 VDD.n2239 VDD.n1054 185
R380 VDD.n2241 VDD.n1061 185
R381 VDD.n2751 VDD.n1061 185
R382 VDD.n2243 VDD.n2242 185
R383 VDD.n2242 VDD.n1068 185
R384 VDD.n2244 VDD.n1067 185
R385 VDD.n2745 VDD.n1067 185
R386 VDD.n2246 VDD.n2245 185
R387 VDD.n2245 VDD.n1065 185
R388 VDD.n2247 VDD.n1073 185
R389 VDD.n2739 VDD.n1073 185
R390 VDD.n2249 VDD.n2248 185
R391 VDD.n2248 VDD.t25 185
R392 VDD.n2250 VDD.n1079 185
R393 VDD.n2733 VDD.n1079 185
R394 VDD.n2252 VDD.n2251 185
R395 VDD.n2251 VDD.n1077 185
R396 VDD.n2253 VDD.n1085 185
R397 VDD.n2727 VDD.n1085 185
R398 VDD.n2255 VDD.n2254 185
R399 VDD.n2254 VDD.n1083 185
R400 VDD.n2256 VDD.n1091 185
R401 VDD.n2721 VDD.n1091 185
R402 VDD.n2258 VDD.n2257 185
R403 VDD.n2257 VDD.n1089 185
R404 VDD.n2259 VDD.n1097 185
R405 VDD.n2715 VDD.n1097 185
R406 VDD.n2261 VDD.n2260 185
R407 VDD.n2260 VDD.n1095 185
R408 VDD.n2262 VDD.n1103 185
R409 VDD.n2709 VDD.n1103 185
R410 VDD.n2264 VDD.n2263 185
R411 VDD.n2263 VDD.n1101 185
R412 VDD.n2265 VDD.n1109 185
R413 VDD.n2703 VDD.n1109 185
R414 VDD.n2267 VDD.n2266 185
R415 VDD.n2266 VDD.n1107 185
R416 VDD.n2268 VDD.n1115 185
R417 VDD.n2697 VDD.n1115 185
R418 VDD.n2270 VDD.n2269 185
R419 VDD.n2269 VDD.n1113 185
R420 VDD.n2271 VDD.n1121 185
R421 VDD.n2691 VDD.n1121 185
R422 VDD.n2273 VDD.n2272 185
R423 VDD.n2272 VDD.n1119 185
R424 VDD.n2274 VDD.n1127 185
R425 VDD.n2685 VDD.n1127 185
R426 VDD.n2276 VDD.n2275 185
R427 VDD.n2275 VDD.n1125 185
R428 VDD.n2277 VDD.n1133 185
R429 VDD.n2679 VDD.n1133 185
R430 VDD.n2279 VDD.n2278 185
R431 VDD.n2278 VDD.n1131 185
R432 VDD.n2280 VDD.n1139 185
R433 VDD.n2673 VDD.n1139 185
R434 VDD.n2282 VDD.n2281 185
R435 VDD.n2281 VDD.n1137 185
R436 VDD.n2283 VDD.n1145 185
R437 VDD.n2667 VDD.n1145 185
R438 VDD.n2285 VDD.n2284 185
R439 VDD.n2284 VDD.n1143 185
R440 VDD.n2286 VDD.n1151 185
R441 VDD.n2661 VDD.n1151 185
R442 VDD.n2288 VDD.n2287 185
R443 VDD.n2287 VDD.n1149 185
R444 VDD.n2289 VDD.n1157 185
R445 VDD.n2655 VDD.n1157 185
R446 VDD.n2291 VDD.n2290 185
R447 VDD.n2290 VDD.n1155 185
R448 VDD.n2292 VDD.n1163 185
R449 VDD.n2649 VDD.n1163 185
R450 VDD.n2294 VDD.n2293 185
R451 VDD.n2293 VDD.n1161 185
R452 VDD.n2295 VDD.n1169 185
R453 VDD.n2643 VDD.n1169 185
R454 VDD.n2297 VDD.n2296 185
R455 VDD.n2296 VDD.n1167 185
R456 VDD.n2298 VDD.n1175 185
R457 VDD.n2637 VDD.n1175 185
R458 VDD.n2300 VDD.n2299 185
R459 VDD.n2299 VDD.n1173 185
R460 VDD.n2301 VDD.n1181 185
R461 VDD.n2631 VDD.n1181 185
R462 VDD.n2303 VDD.n2302 185
R463 VDD.n2302 VDD.n1179 185
R464 VDD.n2304 VDD.n1187 185
R465 VDD.n2625 VDD.n1187 185
R466 VDD.n2306 VDD.n2305 185
R467 VDD.n2305 VDD.n1185 185
R468 VDD.n2307 VDD.n1192 185
R469 VDD.n2619 VDD.n1192 185
R470 VDD.n2470 VDD.n2469 185
R471 VDD.n2469 VDD.n2468 185
R472 VDD.n2471 VDD.n1198 185
R473 VDD.n2613 VDD.n1198 185
R474 VDD.n2473 VDD.n2472 185
R475 VDD.n2472 VDD.n1196 185
R476 VDD.n2474 VDD.n1204 185
R477 VDD.n2607 VDD.n1204 185
R478 VDD.n2476 VDD.n2475 185
R479 VDD.n2475 VDD.n1202 185
R480 VDD.n2477 VDD.n1210 185
R481 VDD.n2601 VDD.n1210 185
R482 VDD.n2479 VDD.n2478 185
R483 VDD.n2478 VDD.n1208 185
R484 VDD.n2480 VDD.n1216 185
R485 VDD.n2595 VDD.n1216 185
R486 VDD.n2482 VDD.n2481 185
R487 VDD.n2482 VDD.n1214 185
R488 VDD.n3662 VDD.n487 185
R489 VDD.n3718 VDD.n487 185
R490 VDD.n3664 VDD.n3663 185
R491 VDD.n3663 VDD.n485 185
R492 VDD.n3665 VDD.n622 185
R493 VDD.n3675 VDD.n622 185
R494 VDD.n3666 VDD.n630 185
R495 VDD.n630 VDD.n620 185
R496 VDD.n3668 VDD.n3667 185
R497 VDD.n3669 VDD.n3668 185
R498 VDD.n3638 VDD.n629 185
R499 VDD.n629 VDD.n626 185
R500 VDD.n3637 VDD.n3636 185
R501 VDD.n3636 VDD.n3635 185
R502 VDD.n632 VDD.n631 185
R503 VDD.n633 VDD.n632 185
R504 VDD.n3628 VDD.n3627 185
R505 VDD.n3629 VDD.n3628 185
R506 VDD.n3626 VDD.n641 185
R507 VDD.n647 VDD.n641 185
R508 VDD.n3625 VDD.n3624 185
R509 VDD.n3624 VDD.n3623 185
R510 VDD.n643 VDD.n642 185
R511 VDD.n644 VDD.n643 185
R512 VDD.n3616 VDD.n3615 185
R513 VDD.n3617 VDD.n3616 185
R514 VDD.n3614 VDD.n654 185
R515 VDD.n654 VDD.n651 185
R516 VDD.n3613 VDD.n3612 185
R517 VDD.n3612 VDD.n3611 185
R518 VDD.n656 VDD.n655 185
R519 VDD.n657 VDD.n656 185
R520 VDD.n3604 VDD.n3603 185
R521 VDD.n3605 VDD.n3604 185
R522 VDD.n3602 VDD.n666 185
R523 VDD.n666 VDD.n663 185
R524 VDD.n3601 VDD.n3600 185
R525 VDD.n3600 VDD.n3599 185
R526 VDD.n668 VDD.n667 185
R527 VDD.n669 VDD.n668 185
R528 VDD.n3592 VDD.n3591 185
R529 VDD.n3593 VDD.n3592 185
R530 VDD.n3590 VDD.n678 185
R531 VDD.n678 VDD.n675 185
R532 VDD.n3589 VDD.n3588 185
R533 VDD.n3588 VDD.n3587 185
R534 VDD.n680 VDD.n679 185
R535 VDD.n681 VDD.n680 185
R536 VDD.n3580 VDD.n3579 185
R537 VDD.n3581 VDD.n3580 185
R538 VDD.n3578 VDD.n690 185
R539 VDD.n690 VDD.n687 185
R540 VDD.n3577 VDD.n3576 185
R541 VDD.n3576 VDD.n3575 185
R542 VDD.n692 VDD.n691 185
R543 VDD.n693 VDD.n692 185
R544 VDD.n3568 VDD.n3567 185
R545 VDD.n3569 VDD.n3568 185
R546 VDD.n3566 VDD.n702 185
R547 VDD.n702 VDD.n699 185
R548 VDD.n3565 VDD.n3564 185
R549 VDD.n3564 VDD.n3563 185
R550 VDD.n704 VDD.n703 185
R551 VDD.n705 VDD.n704 185
R552 VDD.n3556 VDD.n3555 185
R553 VDD.n3557 VDD.n3556 185
R554 VDD.n3554 VDD.n714 185
R555 VDD.n714 VDD.n711 185
R556 VDD.n3553 VDD.n3552 185
R557 VDD.n3552 VDD.n3551 185
R558 VDD.n716 VDD.n715 185
R559 VDD.n717 VDD.n716 185
R560 VDD.n3544 VDD.n3543 185
R561 VDD.n3545 VDD.n3544 185
R562 VDD.n3542 VDD.n726 185
R563 VDD.n726 VDD.n723 185
R564 VDD.n3541 VDD.n3540 185
R565 VDD.n3540 VDD.n3539 185
R566 VDD.n728 VDD.n727 185
R567 VDD.n729 VDD.n728 185
R568 VDD.n3532 VDD.n3531 185
R569 VDD.n3533 VDD.n3532 185
R570 VDD.n3530 VDD.n738 185
R571 VDD.n738 VDD.n735 185
R572 VDD.n3529 VDD.n3528 185
R573 VDD.n3528 VDD.n3527 185
R574 VDD.n740 VDD.n739 185
R575 VDD.n741 VDD.n740 185
R576 VDD.n3520 VDD.n3519 185
R577 VDD.n3521 VDD.n3520 185
R578 VDD.n3518 VDD.n750 185
R579 VDD.n750 VDD.n747 185
R580 VDD.n3517 VDD.n3516 185
R581 VDD.n3516 VDD.n3515 185
R582 VDD.n752 VDD.n751 185
R583 VDD.n753 VDD.n752 185
R584 VDD.n3425 VDD.n760 185
R585 VDD.t16 VDD.n760 185
R586 VDD.n3427 VDD.n3426 185
R587 VDD.n3426 VDD.n759 185
R588 VDD.n3428 VDD.n768 185
R589 VDD.n3438 VDD.n768 185
R590 VDD.n3429 VDD.n775 185
R591 VDD.n775 VDD.n766 185
R592 VDD.n3431 VDD.n3430 185
R593 VDD.n3432 VDD.n3431 185
R594 VDD.n3424 VDD.n774 185
R595 VDD.n781 VDD.n774 185
R596 VDD.n3423 VDD.n3422 185
R597 VDD.n3422 VDD.n3421 185
R598 VDD.n777 VDD.n776 185
R599 VDD.n778 VDD.n777 185
R600 VDD.n3414 VDD.n3413 185
R601 VDD.n3415 VDD.n3414 185
R602 VDD.n3412 VDD.n788 185
R603 VDD.n788 VDD.n785 185
R604 VDD.n3411 VDD.n3410 185
R605 VDD.n3410 VDD.n3409 185
R606 VDD.n790 VDD.n789 185
R607 VDD.n791 VDD.n790 185
R608 VDD.n3402 VDD.n3401 185
R609 VDD.n3403 VDD.n3402 185
R610 VDD.n3400 VDD.n799 185
R611 VDD.n805 VDD.n799 185
R612 VDD.n3399 VDD.n3398 185
R613 VDD.n3398 VDD.n3397 185
R614 VDD.n801 VDD.n800 185
R615 VDD.n802 VDD.n801 185
R616 VDD.n3390 VDD.n3389 185
R617 VDD.n3391 VDD.n3390 185
R618 VDD.n3388 VDD.n811 185
R619 VDD.n817 VDD.n811 185
R620 VDD.n3387 VDD.n3386 185
R621 VDD.n3386 VDD.n3385 185
R622 VDD.n813 VDD.n812 185
R623 VDD.n814 VDD.n813 185
R624 VDD.n3378 VDD.n3377 185
R625 VDD.n3379 VDD.n3378 185
R626 VDD.n3376 VDD.n824 185
R627 VDD.n824 VDD.n821 185
R628 VDD.n3375 VDD.n3374 185
R629 VDD.n3374 VDD.n3373 185
R630 VDD.n826 VDD.n825 185
R631 VDD.n827 VDD.n826 185
R632 VDD.n3366 VDD.n3365 185
R633 VDD.n3367 VDD.n3366 185
R634 VDD.n3364 VDD.n835 185
R635 VDD.n841 VDD.n835 185
R636 VDD.n3363 VDD.n3362 185
R637 VDD.n3362 VDD.n3361 185
R638 VDD.n837 VDD.n836 185
R639 VDD.n838 VDD.n837 185
R640 VDD.n3354 VDD.n3353 185
R641 VDD.n3355 VDD.n3354 185
R642 VDD.n3352 VDD.n848 185
R643 VDD.n848 VDD.n845 185
R644 VDD.n3351 VDD.n3350 185
R645 VDD.n3350 VDD.n3349 185
R646 VDD.n850 VDD.n849 185
R647 VDD.n851 VDD.n850 185
R648 VDD.n3342 VDD.n3341 185
R649 VDD.n3343 VDD.n3342 185
R650 VDD.n3340 VDD.n860 185
R651 VDD.n860 VDD.n857 185
R652 VDD.n3339 VDD.n3338 185
R653 VDD.n3338 VDD.n3337 185
R654 VDD.n862 VDD.n861 185
R655 VDD.n863 VDD.n862 185
R656 VDD.n3330 VDD.n3329 185
R657 VDD.n3331 VDD.n3330 185
R658 VDD.n3328 VDD.n872 185
R659 VDD.n872 VDD.n869 185
R660 VDD.n3327 VDD.n3326 185
R661 VDD.n3326 VDD.n3325 185
R662 VDD.n874 VDD.n873 185
R663 VDD.n875 VDD.n874 185
R664 VDD.n3318 VDD.n3317 185
R665 VDD.n3319 VDD.n3318 185
R666 VDD.n3316 VDD.n883 185
R667 VDD.n3239 VDD.n883 185
R668 VDD.n3315 VDD.n3314 185
R669 VDD.n3314 VDD.n3313 185
R670 VDD.n885 VDD.n884 185
R671 VDD.n886 VDD.n885 185
R672 VDD.n3306 VDD.n3305 185
R673 VDD.n3307 VDD.n3306 185
R674 VDD.n3304 VDD.n895 185
R675 VDD.n895 VDD.n892 185
R676 VDD.n3303 VDD.n3302 185
R677 VDD.n3302 VDD.n3301 185
R678 VDD.n897 VDD.n896 185
R679 VDD.n898 VDD.n897 185
R680 VDD.n3294 VDD.n3293 185
R681 VDD.n3295 VDD.n3294 185
R682 VDD.n3292 VDD.n2979 185
R683 VDD.n3291 VDD.n3290 185
R684 VDD.n3288 VDD.n2980 185
R685 VDD.n3286 VDD.n3285 185
R686 VDD.n3284 VDD.n2981 185
R687 VDD.n3283 VDD.n3282 185
R688 VDD.n3280 VDD.n2982 185
R689 VDD.n3278 VDD.n3277 185
R690 VDD.n3276 VDD.n2983 185
R691 VDD.n3275 VDD.n3274 185
R692 VDD.n3272 VDD.n2984 185
R693 VDD.n3270 VDD.n3269 185
R694 VDD.n3268 VDD.n2985 185
R695 VDD.n3267 VDD.n3266 185
R696 VDD.n3264 VDD.n2986 185
R697 VDD.n3262 VDD.n3261 185
R698 VDD.n3260 VDD.n2987 185
R699 VDD.n3258 VDD.n3257 185
R700 VDD.n3255 VDD.n2990 185
R701 VDD.n3253 VDD.n3252 185
R702 VDD.n3721 VDD.n3720 185
R703 VDD.n3722 VDD.n478 185
R704 VDD.n3724 VDD.n3723 185
R705 VDD.n3726 VDD.n476 185
R706 VDD.n3728 VDD.n3727 185
R707 VDD.n3729 VDD.n475 185
R708 VDD.n3731 VDD.n3730 185
R709 VDD.n3733 VDD.n474 185
R710 VDD.n3734 VDD.n471 185
R711 VDD.n3737 VDD.n3736 185
R712 VDD.n472 VDD.n470 185
R713 VDD.n3646 VDD.n3645 185
R714 VDD.n3648 VDD.n3647 185
R715 VDD.n3650 VDD.n3642 185
R716 VDD.n3652 VDD.n3651 185
R717 VDD.n3653 VDD.n3641 185
R718 VDD.n3655 VDD.n3654 185
R719 VDD.n3657 VDD.n3640 185
R720 VDD.n3658 VDD.n3639 185
R721 VDD.n3661 VDD.n3660 185
R722 VDD.n3719 VDD.n482 185
R723 VDD.n3719 VDD.n3718 185
R724 VDD.n2991 VDD.n484 185
R725 VDD.n485 VDD.n484 185
R726 VDD.n2992 VDD.n621 185
R727 VDD.n3675 VDD.n621 185
R728 VDD.n2994 VDD.n2993 185
R729 VDD.n2993 VDD.n620 185
R730 VDD.n2995 VDD.n628 185
R731 VDD.n3669 VDD.n628 185
R732 VDD.n2997 VDD.n2996 185
R733 VDD.n2996 VDD.n626 185
R734 VDD.n2998 VDD.n635 185
R735 VDD.n3635 VDD.n635 185
R736 VDD.n3000 VDD.n2999 185
R737 VDD.n2999 VDD.n633 185
R738 VDD.n3001 VDD.n640 185
R739 VDD.n3629 VDD.n640 185
R740 VDD.n3003 VDD.n3002 185
R741 VDD.n3002 VDD.n647 185
R742 VDD.n3004 VDD.n646 185
R743 VDD.n3623 VDD.n646 185
R744 VDD.n3006 VDD.n3005 185
R745 VDD.n3005 VDD.n644 185
R746 VDD.n3007 VDD.n653 185
R747 VDD.n3617 VDD.n653 185
R748 VDD.n3009 VDD.n3008 185
R749 VDD.n3008 VDD.n651 185
R750 VDD.n3010 VDD.n659 185
R751 VDD.n3611 VDD.n659 185
R752 VDD.n3012 VDD.n3011 185
R753 VDD.n3011 VDD.n657 185
R754 VDD.n3013 VDD.n665 185
R755 VDD.n3605 VDD.n665 185
R756 VDD.n3015 VDD.n3014 185
R757 VDD.n3014 VDD.n663 185
R758 VDD.n3016 VDD.n671 185
R759 VDD.n3599 VDD.n671 185
R760 VDD.n3018 VDD.n3017 185
R761 VDD.n3017 VDD.n669 185
R762 VDD.n3019 VDD.n677 185
R763 VDD.n3593 VDD.n677 185
R764 VDD.n3021 VDD.n3020 185
R765 VDD.n3020 VDD.n675 185
R766 VDD.n3022 VDD.n683 185
R767 VDD.n3587 VDD.n683 185
R768 VDD.n3024 VDD.n3023 185
R769 VDD.n3023 VDD.n681 185
R770 VDD.n3025 VDD.n689 185
R771 VDD.n3581 VDD.n689 185
R772 VDD.n3027 VDD.n3026 185
R773 VDD.n3026 VDD.n687 185
R774 VDD.n3028 VDD.n695 185
R775 VDD.n3575 VDD.n695 185
R776 VDD.n3030 VDD.n3029 185
R777 VDD.n3029 VDD.n693 185
R778 VDD.n3031 VDD.n701 185
R779 VDD.n3569 VDD.n701 185
R780 VDD.n3033 VDD.n3032 185
R781 VDD.n3032 VDD.n699 185
R782 VDD.n3034 VDD.n707 185
R783 VDD.n3563 VDD.n707 185
R784 VDD.n3036 VDD.n3035 185
R785 VDD.n3035 VDD.n705 185
R786 VDD.n3037 VDD.n713 185
R787 VDD.n3557 VDD.n713 185
R788 VDD.n3039 VDD.n3038 185
R789 VDD.n3038 VDD.n711 185
R790 VDD.n3040 VDD.n719 185
R791 VDD.n3551 VDD.n719 185
R792 VDD.n3042 VDD.n3041 185
R793 VDD.n3041 VDD.n717 185
R794 VDD.n3043 VDD.n725 185
R795 VDD.n3545 VDD.n725 185
R796 VDD.n3045 VDD.n3044 185
R797 VDD.n3044 VDD.n723 185
R798 VDD.n3046 VDD.n731 185
R799 VDD.n3539 VDD.n731 185
R800 VDD.n3048 VDD.n3047 185
R801 VDD.n3047 VDD.n729 185
R802 VDD.n3049 VDD.n737 185
R803 VDD.n3533 VDD.n737 185
R804 VDD.n3051 VDD.n3050 185
R805 VDD.n3050 VDD.n735 185
R806 VDD.n3052 VDD.n743 185
R807 VDD.n3527 VDD.n743 185
R808 VDD.n3054 VDD.n3053 185
R809 VDD.n3053 VDD.n741 185
R810 VDD.n3055 VDD.n749 185
R811 VDD.n3521 VDD.n749 185
R812 VDD.n3057 VDD.n3056 185
R813 VDD.n3056 VDD.n747 185
R814 VDD.n3058 VDD.n755 185
R815 VDD.n3515 VDD.n755 185
R816 VDD.n3060 VDD.n3059 185
R817 VDD.n3059 VDD.n753 185
R818 VDD.n3061 VDD.n761 185
R819 VDD.t16 VDD.n761 185
R820 VDD.n3063 VDD.n3062 185
R821 VDD.n3062 VDD.n759 185
R822 VDD.n3064 VDD.n767 185
R823 VDD.n3438 VDD.n767 185
R824 VDD.n3066 VDD.n3065 185
R825 VDD.n3065 VDD.n766 185
R826 VDD.n3067 VDD.n773 185
R827 VDD.n3432 VDD.n773 185
R828 VDD.n3069 VDD.n3068 185
R829 VDD.n3068 VDD.n781 185
R830 VDD.n3070 VDD.n780 185
R831 VDD.n3421 VDD.n780 185
R832 VDD.n3072 VDD.n3071 185
R833 VDD.n3071 VDD.n778 185
R834 VDD.n3073 VDD.n787 185
R835 VDD.n3415 VDD.n787 185
R836 VDD.n3075 VDD.n3074 185
R837 VDD.n3074 VDD.n785 185
R838 VDD.n3076 VDD.n793 185
R839 VDD.n3409 VDD.n793 185
R840 VDD.n3078 VDD.n3077 185
R841 VDD.n3077 VDD.n791 185
R842 VDD.n3079 VDD.n798 185
R843 VDD.n3403 VDD.n798 185
R844 VDD.n3081 VDD.n3080 185
R845 VDD.n3080 VDD.n805 185
R846 VDD.n3082 VDD.n804 185
R847 VDD.n3397 VDD.n804 185
R848 VDD.n3084 VDD.n3083 185
R849 VDD.n3083 VDD.n802 185
R850 VDD.n3085 VDD.n810 185
R851 VDD.n3391 VDD.n810 185
R852 VDD.n3087 VDD.n3086 185
R853 VDD.n3086 VDD.n817 185
R854 VDD.n3088 VDD.n816 185
R855 VDD.n3385 VDD.n816 185
R856 VDD.n3090 VDD.n3089 185
R857 VDD.n3089 VDD.n814 185
R858 VDD.n3091 VDD.n823 185
R859 VDD.n3379 VDD.n823 185
R860 VDD.n3093 VDD.n3092 185
R861 VDD.n3092 VDD.n821 185
R862 VDD.n3094 VDD.n829 185
R863 VDD.n3373 VDD.n829 185
R864 VDD.n3096 VDD.n3095 185
R865 VDD.n3095 VDD.n827 185
R866 VDD.n3097 VDD.n834 185
R867 VDD.n3367 VDD.n834 185
R868 VDD.n3099 VDD.n3098 185
R869 VDD.n3098 VDD.n841 185
R870 VDD.n3100 VDD.n840 185
R871 VDD.n3361 VDD.n840 185
R872 VDD.n3102 VDD.n3101 185
R873 VDD.n3101 VDD.n838 185
R874 VDD.n3103 VDD.n847 185
R875 VDD.n3355 VDD.n847 185
R876 VDD.n3105 VDD.n3104 185
R877 VDD.n3104 VDD.n845 185
R878 VDD.n3106 VDD.n853 185
R879 VDD.n3349 VDD.n853 185
R880 VDD.n3108 VDD.n3107 185
R881 VDD.n3107 VDD.n851 185
R882 VDD.n3109 VDD.n859 185
R883 VDD.n3343 VDD.n859 185
R884 VDD.n3111 VDD.n3110 185
R885 VDD.n3110 VDD.n857 185
R886 VDD.n3112 VDD.n865 185
R887 VDD.n3337 VDD.n865 185
R888 VDD.n3114 VDD.n3113 185
R889 VDD.n3113 VDD.n863 185
R890 VDD.n3115 VDD.n871 185
R891 VDD.n3331 VDD.n871 185
R892 VDD.n3117 VDD.n3116 185
R893 VDD.n3116 VDD.n869 185
R894 VDD.n3118 VDD.n877 185
R895 VDD.n3325 VDD.n877 185
R896 VDD.n3120 VDD.n3119 185
R897 VDD.n3119 VDD.n875 185
R898 VDD.n3121 VDD.n882 185
R899 VDD.n3319 VDD.n882 185
R900 VDD.n3241 VDD.n3240 185
R901 VDD.n3240 VDD.n3239 185
R902 VDD.n3242 VDD.n888 185
R903 VDD.n3313 VDD.n888 185
R904 VDD.n3244 VDD.n3243 185
R905 VDD.n3243 VDD.n886 185
R906 VDD.n3245 VDD.n894 185
R907 VDD.n3307 VDD.n894 185
R908 VDD.n3247 VDD.n3246 185
R909 VDD.n3246 VDD.n892 185
R910 VDD.n3248 VDD.n900 185
R911 VDD.n3301 VDD.n900 185
R912 VDD.n3250 VDD.n3249 185
R913 VDD.n3249 VDD.n898 185
R914 VDD.n3251 VDD.n2978 185
R915 VDD.n3295 VDD.n2978 185
R916 VDD.n2521 VDD.n2520 185
R917 VDD.n2522 VDD.n2521 185
R918 VDD.n2519 VDD.n1309 185
R919 VDD.n1309 VDD.n1286 185
R920 VDD.n1314 VDD.n1310 185
R921 VDD.n2512 VDD.n1314 185
R922 VDD.n2515 VDD.n2514 185
R923 VDD.n2514 VDD.n2513 185
R924 VDD.n1313 VDD.n1312 185
R925 VDD.n1315 VDD.n1313 185
R926 VDD.n2153 VDD.n2152 185
R927 VDD.n2154 VDD.n2153 185
R928 VDD.n1323 VDD.n1322 185
R929 VDD.n2145 VDD.n1322 185
R930 VDD.n2148 VDD.n2147 185
R931 VDD.n2147 VDD.n2146 185
R932 VDD.n1326 VDD.n1325 185
R933 VDD.n1327 VDD.n1326 185
R934 VDD.n2135 VDD.n2134 185
R935 VDD.n2136 VDD.n2135 185
R936 VDD.n1336 VDD.n1335 185
R937 VDD.n1335 VDD.n1334 185
R938 VDD.n2130 VDD.n2129 185
R939 VDD.n2129 VDD.n2128 185
R940 VDD.n1339 VDD.n1338 185
R941 VDD.n1340 VDD.n1339 185
R942 VDD.n2119 VDD.n2118 185
R943 VDD.n2120 VDD.n2119 185
R944 VDD.n1348 VDD.n1347 185
R945 VDD.n1347 VDD.n1346 185
R946 VDD.n2114 VDD.n2113 185
R947 VDD.n2113 VDD.n2112 185
R948 VDD.n1351 VDD.n1350 185
R949 VDD.n1352 VDD.n1351 185
R950 VDD.n2103 VDD.n2102 185
R951 VDD.n2104 VDD.n2103 185
R952 VDD.n1360 VDD.n1359 185
R953 VDD.n1359 VDD.n1358 185
R954 VDD.n2098 VDD.n2097 185
R955 VDD.n2097 VDD.n2096 185
R956 VDD.n1363 VDD.n1362 185
R957 VDD.n1370 VDD.n1363 185
R958 VDD.n2087 VDD.n2086 185
R959 VDD.n2088 VDD.n2087 185
R960 VDD.n1372 VDD.n1371 185
R961 VDD.n1371 VDD.n1369 185
R962 VDD.n2082 VDD.n2081 185
R963 VDD.n2081 VDD.n2080 185
R964 VDD.n1375 VDD.n1374 185
R965 VDD.n1376 VDD.n1375 185
R966 VDD.n2071 VDD.n2070 185
R967 VDD.n2072 VDD.n2071 185
R968 VDD.n1384 VDD.n1383 185
R969 VDD.n1383 VDD.n1382 185
R970 VDD.n2066 VDD.n2065 185
R971 VDD.n2065 VDD.n2064 185
R972 VDD.n1387 VDD.n1386 185
R973 VDD.n1388 VDD.n1387 185
R974 VDD.n2055 VDD.n2054 185
R975 VDD.n2056 VDD.n2055 185
R976 VDD.n1396 VDD.n1395 185
R977 VDD.n1395 VDD.n1394 185
R978 VDD.n2050 VDD.n2049 185
R979 VDD.n2049 VDD.n2048 185
R980 VDD.n1399 VDD.n1398 185
R981 VDD.n1400 VDD.n1399 185
R982 VDD.n2039 VDD.n2038 185
R983 VDD.n2040 VDD.n2039 185
R984 VDD.n1408 VDD.n1407 185
R985 VDD.n1407 VDD.n1406 185
R986 VDD.n2034 VDD.n2033 185
R987 VDD.n2033 VDD.n2032 185
R988 VDD.n1411 VDD.n1410 185
R989 VDD.n1412 VDD.n1411 185
R990 VDD.n2023 VDD.n2022 185
R991 VDD.n2024 VDD.n2023 185
R992 VDD.n1420 VDD.n1419 185
R993 VDD.n1419 VDD.n1418 185
R994 VDD.n2018 VDD.n2017 185
R995 VDD.n2017 VDD.n2016 185
R996 VDD.n1423 VDD.n1422 185
R997 VDD.n1424 VDD.n1423 185
R998 VDD.n2007 VDD.n2006 185
R999 VDD.n2008 VDD.n2007 185
R1000 VDD.n1431 VDD.n1430 185
R1001 VDD.n1999 VDD.n1430 185
R1002 VDD.n2002 VDD.n2001 185
R1003 VDD.n2001 VDD.n2000 185
R1004 VDD.n1434 VDD.n1433 185
R1005 VDD.n1435 VDD.n1434 185
R1006 VDD.n1990 VDD.n1989 185
R1007 VDD.n1991 VDD.n1990 185
R1008 VDD.n1443 VDD.n1442 185
R1009 VDD.n1442 VDD.n1441 185
R1010 VDD.n1985 VDD.n1984 185
R1011 VDD.n1984 VDD.n1983 185
R1012 VDD.n1446 VDD.n1445 185
R1013 VDD.n1447 VDD.n1446 185
R1014 VDD.n1974 VDD.n1973 185
R1015 VDD.n1975 VDD.n1974 185
R1016 VDD.n1455 VDD.n1454 185
R1017 VDD.n1454 VDD.n1453 185
R1018 VDD.n1969 VDD.n1968 185
R1019 VDD.n1968 VDD.n1967 185
R1020 VDD.n1458 VDD.n1457 185
R1021 VDD.n1459 VDD.n1458 185
R1022 VDD.n1959 VDD.n1958 185
R1023 VDD.t26 VDD.n1959 185
R1024 VDD.n1467 VDD.n1466 185
R1025 VDD.n1466 VDD.n1465 185
R1026 VDD.n1940 VDD.n1939 185
R1027 VDD.n1939 VDD.n1938 185
R1028 VDD.n1470 VDD.n1469 185
R1029 VDD.n1471 VDD.n1470 185
R1030 VDD.n1929 VDD.n1928 185
R1031 VDD.n1930 VDD.n1929 185
R1032 VDD.n1479 VDD.n1478 185
R1033 VDD.n1478 VDD.n1477 185
R1034 VDD.n1924 VDD.n1923 185
R1035 VDD.n1923 VDD.n1922 185
R1036 VDD.n1482 VDD.n1481 185
R1037 VDD.n1483 VDD.n1482 185
R1038 VDD.n1913 VDD.n1912 185
R1039 VDD.n1914 VDD.n1913 185
R1040 VDD.n1491 VDD.n1490 185
R1041 VDD.n1490 VDD.n1489 185
R1042 VDD.n1908 VDD.n1907 185
R1043 VDD.n1907 VDD.n1906 185
R1044 VDD.n1494 VDD.n1493 185
R1045 VDD.n1495 VDD.n1494 185
R1046 VDD.n1897 VDD.n1896 185
R1047 VDD.n1898 VDD.n1897 185
R1048 VDD.n1503 VDD.n1502 185
R1049 VDD.n1502 VDD.n1501 185
R1050 VDD.n1892 VDD.n1891 185
R1051 VDD.n1891 VDD.n1890 185
R1052 VDD.n1506 VDD.n1505 185
R1053 VDD.n1507 VDD.n1506 185
R1054 VDD.n1881 VDD.n1880 185
R1055 VDD.n1882 VDD.n1881 185
R1056 VDD.n1515 VDD.n1514 185
R1057 VDD.n1514 VDD.n1513 185
R1058 VDD.n1876 VDD.n1875 185
R1059 VDD.n1875 VDD.n1874 185
R1060 VDD.n1518 VDD.n1517 185
R1061 VDD.n1519 VDD.n1518 185
R1062 VDD.n1865 VDD.n1864 185
R1063 VDD.n1866 VDD.n1865 185
R1064 VDD.n1527 VDD.n1526 185
R1065 VDD.n1526 VDD.n1525 185
R1066 VDD.n1860 VDD.n1859 185
R1067 VDD.n1859 VDD.n1858 185
R1068 VDD.n1530 VDD.n1529 185
R1069 VDD.n1537 VDD.n1530 185
R1070 VDD.n1849 VDD.n1848 185
R1071 VDD.n1850 VDD.n1849 185
R1072 VDD.n1539 VDD.n1538 185
R1073 VDD.n1538 VDD.n1536 185
R1074 VDD.n1844 VDD.n1843 185
R1075 VDD.n1843 VDD.n1842 185
R1076 VDD.n1542 VDD.n1541 185
R1077 VDD.n1543 VDD.n1542 185
R1078 VDD.n1833 VDD.n1832 185
R1079 VDD.n1834 VDD.n1833 185
R1080 VDD.n1551 VDD.n1550 185
R1081 VDD.n1550 VDD.n1549 185
R1082 VDD.n1828 VDD.n1827 185
R1083 VDD.n1827 VDD.n1826 185
R1084 VDD.n1554 VDD.n1553 185
R1085 VDD.n1555 VDD.n1554 185
R1086 VDD.n1817 VDD.n1816 185
R1087 VDD.n1818 VDD.n1817 185
R1088 VDD.n1563 VDD.n1562 185
R1089 VDD.n1562 VDD.n1561 185
R1090 VDD.n1812 VDD.n1811 185
R1091 VDD.n1811 VDD.n1810 185
R1092 VDD.n1566 VDD.n1565 185
R1093 VDD.n1567 VDD.n1566 185
R1094 VDD.n1801 VDD.n1800 185
R1095 VDD.n1802 VDD.n1801 185
R1096 VDD.n1575 VDD.n1574 185
R1097 VDD.n1574 VDD.n1573 185
R1098 VDD.n1796 VDD.n1795 185
R1099 VDD.n1795 VDD.n1794 185
R1100 VDD.n1578 VDD.n1577 185
R1101 VDD.n1579 VDD.n1578 185
R1102 VDD.n1785 VDD.n1784 185
R1103 VDD.n1786 VDD.n1785 185
R1104 VDD.n1587 VDD.n1586 185
R1105 VDD.n1586 VDD.n1585 185
R1106 VDD.n1780 VDD.n1779 185
R1107 VDD.n1779 VDD.n1778 185
R1108 VDD.n1590 VDD.n1589 185
R1109 VDD.n1591 VDD.n1590 185
R1110 VDD.n1769 VDD.n1768 185
R1111 VDD.n1770 VDD.n1769 185
R1112 VDD.n1599 VDD.n1598 185
R1113 VDD.n1598 VDD.n1597 185
R1114 VDD.n1764 VDD.n1763 185
R1115 VDD.n1763 VDD.n1762 185
R1116 VDD.n1602 VDD.n1601 185
R1117 VDD.n1603 VDD.n1602 185
R1118 VDD.n1753 VDD.n1752 185
R1119 VDD.n1754 VDD.n1753 185
R1120 VDD.n1611 VDD.n1610 185
R1121 VDD.n1610 VDD.n1609 185
R1122 VDD.n1748 VDD.n1747 185
R1123 VDD.n1747 VDD.n1746 185
R1124 VDD.n1614 VDD.n1613 185
R1125 VDD.n1615 VDD.n1614 185
R1126 VDD.n1737 VDD.n1736 185
R1127 VDD.n1738 VDD.n1737 185
R1128 VDD.n1623 VDD.n1622 185
R1129 VDD.n1622 VDD.n1621 185
R1130 VDD.n1732 VDD.n1731 185
R1131 VDD.n1626 VDD.n1625 185
R1132 VDD.n1728 VDD.n1727 185
R1133 VDD.n1729 VDD.n1728 185
R1134 VDD.n1642 VDD.n1641 185
R1135 VDD.n1723 VDD.n1644 185
R1136 VDD.n1722 VDD.n1645 185
R1137 VDD.n1721 VDD.n1646 185
R1138 VDD.n1648 VDD.n1647 185
R1139 VDD.n1717 VDD.n1650 185
R1140 VDD.n1716 VDD.n1651 185
R1141 VDD.n1715 VDD.n1652 185
R1142 VDD.n1654 VDD.n1653 185
R1143 VDD.n1711 VDD.n1656 185
R1144 VDD.n1710 VDD.n1707 185
R1145 VDD.n1706 VDD.n1657 185
R1146 VDD.n1659 VDD.n1658 185
R1147 VDD.n1702 VDD.n1661 185
R1148 VDD.n1701 VDD.n1662 185
R1149 VDD.n1700 VDD.n1663 185
R1150 VDD.n1665 VDD.n1664 185
R1151 VDD.n1696 VDD.n1667 185
R1152 VDD.n1695 VDD.n1668 185
R1153 VDD.n1694 VDD.n1669 185
R1154 VDD.n1671 VDD.n1670 185
R1155 VDD.n1690 VDD.n1673 185
R1156 VDD.n1689 VDD.n1674 185
R1157 VDD.n1688 VDD.n1675 185
R1158 VDD.n1677 VDD.n1676 185
R1159 VDD.n1684 VDD.n1679 185
R1160 VDD.n1680 VDD.n1640 185
R1161 VDD.n1729 VDD.n1640 185
R1162 VDD.n2525 VDD.n2524 185
R1163 VDD.n2527 VDD.n1280 185
R1164 VDD.n1306 VDD.n1278 185
R1165 VDD.n2531 VDD.n1277 185
R1166 VDD.n2532 VDD.n1276 185
R1167 VDD.n2533 VDD.n1275 185
R1168 VDD.n1303 VDD.n1273 185
R1169 VDD.n2537 VDD.n1272 185
R1170 VDD.n2538 VDD.n1271 185
R1171 VDD.n2539 VDD.n1270 185
R1172 VDD.n1300 VDD.n1268 185
R1173 VDD.n2543 VDD.n1267 185
R1174 VDD.n2544 VDD.n1266 185
R1175 VDD.n2545 VDD.n1265 185
R1176 VDD.n1297 VDD.n1263 185
R1177 VDD.n2549 VDD.n1262 185
R1178 VDD.n2550 VDD.n1261 185
R1179 VDD.n2551 VDD.n1258 185
R1180 VDD.n1294 VDD.n1256 185
R1181 VDD.n2555 VDD.n1255 185
R1182 VDD.n2556 VDD.n1254 185
R1183 VDD.n2557 VDD.n1253 185
R1184 VDD.n1291 VDD.n1251 185
R1185 VDD.n2561 VDD.n1250 185
R1186 VDD.n2562 VDD.n1249 185
R1187 VDD.n2563 VDD.n1248 185
R1188 VDD.n1288 VDD.n1246 185
R1189 VDD.n2567 VDD.n1245 185
R1190 VDD.n2568 VDD.n1244 185
R1191 VDD.n2569 VDD.n1243 185
R1192 VDD.n2523 VDD.n1285 185
R1193 VDD.n2523 VDD.n2522 185
R1194 VDD.n1318 VDD.n1284 185
R1195 VDD.n1286 VDD.n1284 185
R1196 VDD.n2511 VDD.n2510 185
R1197 VDD.n2512 VDD.n2511 185
R1198 VDD.n1317 VDD.n1316 185
R1199 VDD.n2513 VDD.n1316 185
R1200 VDD.n2157 VDD.n2156 185
R1201 VDD.n2156 VDD.n1315 185
R1202 VDD.n2155 VDD.n1320 185
R1203 VDD.n2155 VDD.n2154 185
R1204 VDD.n1330 VDD.n1321 185
R1205 VDD.n2145 VDD.n1321 185
R1206 VDD.n2144 VDD.n2143 185
R1207 VDD.n2146 VDD.n2144 185
R1208 VDD.n1329 VDD.n1328 185
R1209 VDD.n1328 VDD.n1327 185
R1210 VDD.n2138 VDD.n2137 185
R1211 VDD.n2137 VDD.n2136 185
R1212 VDD.n1333 VDD.n1332 185
R1213 VDD.n1334 VDD.n1333 185
R1214 VDD.n2127 VDD.n2126 185
R1215 VDD.n2128 VDD.n2127 185
R1216 VDD.n1342 VDD.n1341 185
R1217 VDD.n1341 VDD.n1340 185
R1218 VDD.n2122 VDD.n2121 185
R1219 VDD.n2121 VDD.n2120 185
R1220 VDD.n1345 VDD.n1344 185
R1221 VDD.n1346 VDD.n1345 185
R1222 VDD.n2111 VDD.n2110 185
R1223 VDD.n2112 VDD.n2111 185
R1224 VDD.n1354 VDD.n1353 185
R1225 VDD.n1353 VDD.n1352 185
R1226 VDD.n2106 VDD.n2105 185
R1227 VDD.n2105 VDD.n2104 185
R1228 VDD.n1357 VDD.n1356 185
R1229 VDD.n1358 VDD.n1357 185
R1230 VDD.n2095 VDD.n2094 185
R1231 VDD.n2096 VDD.n2095 185
R1232 VDD.n1365 VDD.n1364 185
R1233 VDD.n1370 VDD.n1364 185
R1234 VDD.n2090 VDD.n2089 185
R1235 VDD.n2089 VDD.n2088 185
R1236 VDD.n1368 VDD.n1367 185
R1237 VDD.n1369 VDD.n1368 185
R1238 VDD.n2079 VDD.n2078 185
R1239 VDD.n2080 VDD.n2079 185
R1240 VDD.n1378 VDD.n1377 185
R1241 VDD.n1377 VDD.n1376 185
R1242 VDD.n2074 VDD.n2073 185
R1243 VDD.n2073 VDD.n2072 185
R1244 VDD.n1381 VDD.n1380 185
R1245 VDD.n1382 VDD.n1381 185
R1246 VDD.n2063 VDD.n2062 185
R1247 VDD.n2064 VDD.n2063 185
R1248 VDD.n1390 VDD.n1389 185
R1249 VDD.n1389 VDD.n1388 185
R1250 VDD.n2058 VDD.n2057 185
R1251 VDD.n2057 VDD.n2056 185
R1252 VDD.n1393 VDD.n1392 185
R1253 VDD.n1394 VDD.n1393 185
R1254 VDD.n2047 VDD.n2046 185
R1255 VDD.n2048 VDD.n2047 185
R1256 VDD.n1402 VDD.n1401 185
R1257 VDD.n1401 VDD.n1400 185
R1258 VDD.n2042 VDD.n2041 185
R1259 VDD.n2041 VDD.n2040 185
R1260 VDD.n1405 VDD.n1404 185
R1261 VDD.n1406 VDD.n1405 185
R1262 VDD.n2031 VDD.n2030 185
R1263 VDD.n2032 VDD.n2031 185
R1264 VDD.n1414 VDD.n1413 185
R1265 VDD.n1413 VDD.n1412 185
R1266 VDD.n2026 VDD.n2025 185
R1267 VDD.n2025 VDD.n2024 185
R1268 VDD.n1417 VDD.n1416 185
R1269 VDD.n1418 VDD.n1417 185
R1270 VDD.n2015 VDD.n2014 185
R1271 VDD.n2016 VDD.n2015 185
R1272 VDD.n1426 VDD.n1425 185
R1273 VDD.n1425 VDD.n1424 185
R1274 VDD.n2010 VDD.n2009 185
R1275 VDD.n2009 VDD.n2008 185
R1276 VDD.n1429 VDD.n1428 185
R1277 VDD.n1999 VDD.n1429 185
R1278 VDD.n1998 VDD.n1997 185
R1279 VDD.n2000 VDD.n1998 185
R1280 VDD.n1437 VDD.n1436 185
R1281 VDD.n1436 VDD.n1435 185
R1282 VDD.n1993 VDD.n1992 185
R1283 VDD.n1992 VDD.n1991 185
R1284 VDD.n1440 VDD.n1439 185
R1285 VDD.n1441 VDD.n1440 185
R1286 VDD.n1982 VDD.n1981 185
R1287 VDD.n1983 VDD.n1982 185
R1288 VDD.n1449 VDD.n1448 185
R1289 VDD.n1448 VDD.n1447 185
R1290 VDD.n1977 VDD.n1976 185
R1291 VDD.n1976 VDD.n1975 185
R1292 VDD.n1452 VDD.n1451 185
R1293 VDD.n1453 VDD.n1452 185
R1294 VDD.n1966 VDD.n1965 185
R1295 VDD.n1967 VDD.n1966 185
R1296 VDD.n1461 VDD.n1460 185
R1297 VDD.n1460 VDD.n1459 185
R1298 VDD.n1961 VDD.n1960 185
R1299 VDD.n1960 VDD.t26 185
R1300 VDD.n1464 VDD.n1463 185
R1301 VDD.n1465 VDD.n1464 185
R1302 VDD.n1937 VDD.n1936 185
R1303 VDD.n1938 VDD.n1937 185
R1304 VDD.n1473 VDD.n1472 185
R1305 VDD.n1472 VDD.n1471 185
R1306 VDD.n1932 VDD.n1931 185
R1307 VDD.n1931 VDD.n1930 185
R1308 VDD.n1476 VDD.n1475 185
R1309 VDD.n1477 VDD.n1476 185
R1310 VDD.n1921 VDD.n1920 185
R1311 VDD.n1922 VDD.n1921 185
R1312 VDD.n1485 VDD.n1484 185
R1313 VDD.n1484 VDD.n1483 185
R1314 VDD.n1916 VDD.n1915 185
R1315 VDD.n1915 VDD.n1914 185
R1316 VDD.n1488 VDD.n1487 185
R1317 VDD.n1489 VDD.n1488 185
R1318 VDD.n1905 VDD.n1904 185
R1319 VDD.n1906 VDD.n1905 185
R1320 VDD.n1497 VDD.n1496 185
R1321 VDD.n1496 VDD.n1495 185
R1322 VDD.n1900 VDD.n1899 185
R1323 VDD.n1899 VDD.n1898 185
R1324 VDD.n1500 VDD.n1499 185
R1325 VDD.n1501 VDD.n1500 185
R1326 VDD.n1889 VDD.n1888 185
R1327 VDD.n1890 VDD.n1889 185
R1328 VDD.n1509 VDD.n1508 185
R1329 VDD.n1508 VDD.n1507 185
R1330 VDD.n1884 VDD.n1883 185
R1331 VDD.n1883 VDD.n1882 185
R1332 VDD.n1512 VDD.n1511 185
R1333 VDD.n1513 VDD.n1512 185
R1334 VDD.n1873 VDD.n1872 185
R1335 VDD.n1874 VDD.n1873 185
R1336 VDD.n1521 VDD.n1520 185
R1337 VDD.n1520 VDD.n1519 185
R1338 VDD.n1868 VDD.n1867 185
R1339 VDD.n1867 VDD.n1866 185
R1340 VDD.n1524 VDD.n1523 185
R1341 VDD.n1525 VDD.n1524 185
R1342 VDD.n1857 VDD.n1856 185
R1343 VDD.n1858 VDD.n1857 185
R1344 VDD.n1532 VDD.n1531 185
R1345 VDD.n1537 VDD.n1531 185
R1346 VDD.n1852 VDD.n1851 185
R1347 VDD.n1851 VDD.n1850 185
R1348 VDD.n1535 VDD.n1534 185
R1349 VDD.n1536 VDD.n1535 185
R1350 VDD.n1841 VDD.n1840 185
R1351 VDD.n1842 VDD.n1841 185
R1352 VDD.n1545 VDD.n1544 185
R1353 VDD.n1544 VDD.n1543 185
R1354 VDD.n1836 VDD.n1835 185
R1355 VDD.n1835 VDD.n1834 185
R1356 VDD.n1548 VDD.n1547 185
R1357 VDD.n1549 VDD.n1548 185
R1358 VDD.n1825 VDD.n1824 185
R1359 VDD.n1826 VDD.n1825 185
R1360 VDD.n1557 VDD.n1556 185
R1361 VDD.n1556 VDD.n1555 185
R1362 VDD.n1820 VDD.n1819 185
R1363 VDD.n1819 VDD.n1818 185
R1364 VDD.n1560 VDD.n1559 185
R1365 VDD.n1561 VDD.n1560 185
R1366 VDD.n1809 VDD.n1808 185
R1367 VDD.n1810 VDD.n1809 185
R1368 VDD.n1569 VDD.n1568 185
R1369 VDD.n1568 VDD.n1567 185
R1370 VDD.n1804 VDD.n1803 185
R1371 VDD.n1803 VDD.n1802 185
R1372 VDD.n1572 VDD.n1571 185
R1373 VDD.n1573 VDD.n1572 185
R1374 VDD.n1793 VDD.n1792 185
R1375 VDD.n1794 VDD.n1793 185
R1376 VDD.n1581 VDD.n1580 185
R1377 VDD.n1580 VDD.n1579 185
R1378 VDD.n1788 VDD.n1787 185
R1379 VDD.n1787 VDD.n1786 185
R1380 VDD.n1584 VDD.n1583 185
R1381 VDD.n1585 VDD.n1584 185
R1382 VDD.n1777 VDD.n1776 185
R1383 VDD.n1778 VDD.n1777 185
R1384 VDD.n1593 VDD.n1592 185
R1385 VDD.n1592 VDD.n1591 185
R1386 VDD.n1772 VDD.n1771 185
R1387 VDD.n1771 VDD.n1770 185
R1388 VDD.n1596 VDD.n1595 185
R1389 VDD.n1597 VDD.n1596 185
R1390 VDD.n1761 VDD.n1760 185
R1391 VDD.n1762 VDD.n1761 185
R1392 VDD.n1605 VDD.n1604 185
R1393 VDD.n1604 VDD.n1603 185
R1394 VDD.n1756 VDD.n1755 185
R1395 VDD.n1755 VDD.n1754 185
R1396 VDD.n1608 VDD.n1607 185
R1397 VDD.n1609 VDD.n1608 185
R1398 VDD.n1745 VDD.n1744 185
R1399 VDD.n1746 VDD.n1745 185
R1400 VDD.n1617 VDD.n1616 185
R1401 VDD.n1616 VDD.n1615 185
R1402 VDD.n1740 VDD.n1739 185
R1403 VDD.n1739 VDD.n1738 185
R1404 VDD.n1620 VDD.n1619 185
R1405 VDD.n1621 VDD.n1620 185
R1406 VDD.n177 VDD.n176 185
R1407 VDD.n4051 VDD.n177 185
R1408 VDD.n4054 VDD.n4053 185
R1409 VDD.n4053 VDD.n4052 185
R1410 VDD.n4055 VDD.n171 185
R1411 VDD.n171 VDD.n170 185
R1412 VDD.n4057 VDD.n4056 185
R1413 VDD.n4058 VDD.n4057 185
R1414 VDD.n166 VDD.n165 185
R1415 VDD.n4059 VDD.n166 185
R1416 VDD.n4062 VDD.n4061 185
R1417 VDD.n4061 VDD.n4060 185
R1418 VDD.n4063 VDD.n160 185
R1419 VDD.n160 VDD.n159 185
R1420 VDD.n4065 VDD.n4064 185
R1421 VDD.n4066 VDD.n4065 185
R1422 VDD.n155 VDD.n154 185
R1423 VDD.n4067 VDD.n155 185
R1424 VDD.n4070 VDD.n4069 185
R1425 VDD.n4069 VDD.n4068 185
R1426 VDD.n4071 VDD.n149 185
R1427 VDD.n149 VDD.n148 185
R1428 VDD.n4073 VDD.n4072 185
R1429 VDD.n4074 VDD.n4073 185
R1430 VDD.n144 VDD.n143 185
R1431 VDD.n4075 VDD.n144 185
R1432 VDD.n4078 VDD.n4077 185
R1433 VDD.n4077 VDD.n4076 185
R1434 VDD.n4079 VDD.n138 185
R1435 VDD.n138 VDD.n137 185
R1436 VDD.n4081 VDD.n4080 185
R1437 VDD.n4082 VDD.n4081 185
R1438 VDD.n133 VDD.n132 185
R1439 VDD.n4083 VDD.n133 185
R1440 VDD.n4086 VDD.n4085 185
R1441 VDD.n4085 VDD.n4084 185
R1442 VDD.n4087 VDD.n127 185
R1443 VDD.n127 VDD.n126 185
R1444 VDD.n4089 VDD.n4088 185
R1445 VDD.n4090 VDD.n4089 185
R1446 VDD.n122 VDD.n121 185
R1447 VDD.n4091 VDD.n122 185
R1448 VDD.n4094 VDD.n4093 185
R1449 VDD.n4093 VDD.n4092 185
R1450 VDD.n4095 VDD.n116 185
R1451 VDD.n116 VDD.n115 185
R1452 VDD.n4097 VDD.n4096 185
R1453 VDD.n4098 VDD.n4097 185
R1454 VDD.n111 VDD.n110 185
R1455 VDD.n4099 VDD.n111 185
R1456 VDD.n4102 VDD.n4101 185
R1457 VDD.n4101 VDD.n4100 185
R1458 VDD.n4103 VDD.n105 185
R1459 VDD.n105 VDD.n104 185
R1460 VDD.n4105 VDD.n4104 185
R1461 VDD.n4106 VDD.n4105 185
R1462 VDD.n99 VDD.n98 185
R1463 VDD.n4107 VDD.n99 185
R1464 VDD.n4110 VDD.n4109 185
R1465 VDD.n4109 VDD.n4108 185
R1466 VDD.n4111 VDD.n93 185
R1467 VDD.n100 VDD.n93 185
R1468 VDD.n4113 VDD.n4112 185
R1469 VDD.n4114 VDD.n4113 185
R1470 VDD.n89 VDD.n88 185
R1471 VDD.n4115 VDD.n89 185
R1472 VDD.n4118 VDD.n4117 185
R1473 VDD.n4117 VDD.n4116 185
R1474 VDD.n4119 VDD.n83 185
R1475 VDD.n83 VDD.n82 185
R1476 VDD.n4121 VDD.n4120 185
R1477 VDD.n4122 VDD.n4121 185
R1478 VDD.n78 VDD.n77 185
R1479 VDD.n4123 VDD.n78 185
R1480 VDD.n4126 VDD.n4125 185
R1481 VDD.n4125 VDD.n4124 185
R1482 VDD.n4127 VDD.n72 185
R1483 VDD.n72 VDD.n71 185
R1484 VDD.n4129 VDD.n4128 185
R1485 VDD.n4130 VDD.n4129 185
R1486 VDD.n67 VDD.n66 185
R1487 VDD.n4131 VDD.n67 185
R1488 VDD.n4134 VDD.n4133 185
R1489 VDD.n4133 VDD.n4132 185
R1490 VDD.n4135 VDD.n61 185
R1491 VDD.n61 VDD.n60 185
R1492 VDD.n4137 VDD.n4136 185
R1493 VDD.n4138 VDD.n4137 185
R1494 VDD.n56 VDD.n55 185
R1495 VDD.n4139 VDD.n56 185
R1496 VDD.n4142 VDD.n4141 185
R1497 VDD.n4141 VDD.n4140 185
R1498 VDD.n4143 VDD.n50 185
R1499 VDD.n50 VDD.n49 185
R1500 VDD.n4145 VDD.n4144 185
R1501 VDD.n4146 VDD.n4145 185
R1502 VDD.n45 VDD.n44 185
R1503 VDD.n4147 VDD.n45 185
R1504 VDD.n4150 VDD.n4149 185
R1505 VDD.n4149 VDD.n4148 185
R1506 VDD.n4151 VDD.n40 185
R1507 VDD.n40 VDD.n39 185
R1508 VDD.n4153 VDD.n4152 185
R1509 VDD.n4154 VDD.n4153 185
R1510 VDD.n34 VDD.n32 185
R1511 VDD.n4155 VDD.n34 185
R1512 VDD.n4157 VDD.n4156 185
R1513 VDD.n4156 VDD.t23 185
R1514 VDD.n33 VDD.n31 185
R1515 VDD.n35 VDD.n33 185
R1516 VDD.n3947 VDD.n3946 185
R1517 VDD.n3948 VDD.n3947 185
R1518 VDD.n319 VDD.n318 185
R1519 VDD.n318 VDD.n317 185
R1520 VDD.n3942 VDD.n3941 185
R1521 VDD.n3941 VDD.n3940 185
R1522 VDD.n322 VDD.n321 185
R1523 VDD.n323 VDD.n322 185
R1524 VDD.n3928 VDD.n3927 185
R1525 VDD.n3929 VDD.n3928 185
R1526 VDD.n331 VDD.n330 185
R1527 VDD.n330 VDD.n329 185
R1528 VDD.n3923 VDD.n3922 185
R1529 VDD.n3922 VDD.n3921 185
R1530 VDD.n334 VDD.n333 185
R1531 VDD.n335 VDD.n334 185
R1532 VDD.n3912 VDD.n3911 185
R1533 VDD.n3913 VDD.n3912 185
R1534 VDD.n343 VDD.n342 185
R1535 VDD.n342 VDD.n341 185
R1536 VDD.n3907 VDD.n3906 185
R1537 VDD.n3906 VDD.n3905 185
R1538 VDD.n346 VDD.n345 185
R1539 VDD.n347 VDD.n346 185
R1540 VDD.n3896 VDD.n3895 185
R1541 VDD.n3897 VDD.n3896 185
R1542 VDD.n355 VDD.n354 185
R1543 VDD.n354 VDD.n353 185
R1544 VDD.n3891 VDD.n3890 185
R1545 VDD.n3890 VDD.n3889 185
R1546 VDD.n358 VDD.n357 185
R1547 VDD.n359 VDD.n358 185
R1548 VDD.n3880 VDD.n3879 185
R1549 VDD.n3881 VDD.n3880 185
R1550 VDD.n367 VDD.n366 185
R1551 VDD.n366 VDD.n365 185
R1552 VDD.n3875 VDD.n3874 185
R1553 VDD.n3874 VDD.n3873 185
R1554 VDD.n370 VDD.n369 185
R1555 VDD.n371 VDD.n370 185
R1556 VDD.n3864 VDD.n3863 185
R1557 VDD.n3865 VDD.n3864 185
R1558 VDD.n378 VDD.n377 185
R1559 VDD.n3856 VDD.n377 185
R1560 VDD.n3859 VDD.n3858 185
R1561 VDD.n3858 VDD.n3857 185
R1562 VDD.n381 VDD.n380 185
R1563 VDD.n382 VDD.n381 185
R1564 VDD.n3847 VDD.n3846 185
R1565 VDD.n3848 VDD.n3847 185
R1566 VDD.n390 VDD.n389 185
R1567 VDD.n389 VDD.n388 185
R1568 VDD.n3842 VDD.n3841 185
R1569 VDD.n3841 VDD.n3840 185
R1570 VDD.n393 VDD.n392 185
R1571 VDD.n394 VDD.n393 185
R1572 VDD.n3831 VDD.n3830 185
R1573 VDD.n3832 VDD.n3831 185
R1574 VDD.n402 VDD.n401 185
R1575 VDD.n401 VDD.n400 185
R1576 VDD.n3826 VDD.n3825 185
R1577 VDD.n3825 VDD.n3824 185
R1578 VDD.n405 VDD.n404 185
R1579 VDD.n406 VDD.n405 185
R1580 VDD.n3815 VDD.n3814 185
R1581 VDD.n3816 VDD.n3815 185
R1582 VDD.n414 VDD.n413 185
R1583 VDD.n413 VDD.n412 185
R1584 VDD.n3810 VDD.n3809 185
R1585 VDD.n3809 VDD.n3808 185
R1586 VDD.n417 VDD.n416 185
R1587 VDD.n418 VDD.n417 185
R1588 VDD.n3799 VDD.n3798 185
R1589 VDD.n3800 VDD.n3799 185
R1590 VDD.n426 VDD.n425 185
R1591 VDD.n425 VDD.n424 185
R1592 VDD.n3794 VDD.n3793 185
R1593 VDD.n3793 VDD.n3792 185
R1594 VDD.n429 VDD.n428 185
R1595 VDD.n430 VDD.n429 185
R1596 VDD.n3783 VDD.n3782 185
R1597 VDD.n3784 VDD.n3783 185
R1598 VDD.n438 VDD.n437 185
R1599 VDD.n437 VDD.n436 185
R1600 VDD.n3778 VDD.n3777 185
R1601 VDD.n3777 VDD.n3776 185
R1602 VDD.n441 VDD.n440 185
R1603 VDD.n442 VDD.n441 185
R1604 VDD.n3767 VDD.n3766 185
R1605 VDD.n3768 VDD.n3767 185
R1606 VDD.n450 VDD.n449 185
R1607 VDD.n449 VDD.n448 185
R1608 VDD.n3762 VDD.n3761 185
R1609 VDD.n3761 VDD.n3760 185
R1610 VDD.n453 VDD.n452 185
R1611 VDD.n454 VDD.n453 185
R1612 VDD.n3751 VDD.n3750 185
R1613 VDD.n3752 VDD.n3751 185
R1614 VDD.n462 VDD.n461 185
R1615 VDD.n461 VDD.n460 185
R1616 VDD.n3746 VDD.n3745 185
R1617 VDD.n3745 VDD.n3744 185
R1618 VDD.n465 VDD.n464 185
R1619 VDD.n466 VDD.n465 185
R1620 VDD.n604 VDD.n603 185
R1621 VDD.n499 VDD.n498 185
R1622 VDD.n600 VDD.n599 185
R1623 VDD.n601 VDD.n600 185
R1624 VDD.n598 VDD.n514 185
R1625 VDD.n597 VDD.n596 185
R1626 VDD.n595 VDD.n594 185
R1627 VDD.n593 VDD.n592 185
R1628 VDD.n591 VDD.n590 185
R1629 VDD.n589 VDD.n588 185
R1630 VDD.n587 VDD.n586 185
R1631 VDD.n585 VDD.n584 185
R1632 VDD.n583 VDD.n582 185
R1633 VDD.n581 VDD.n580 185
R1634 VDD.n579 VDD.n578 185
R1635 VDD.n577 VDD.n576 185
R1636 VDD.n575 VDD.n574 185
R1637 VDD.n573 VDD.n572 185
R1638 VDD.n571 VDD.n570 185
R1639 VDD.n569 VDD.n568 185
R1640 VDD.n567 VDD.n566 185
R1641 VDD.n565 VDD.n564 185
R1642 VDD.n563 VDD.n562 185
R1643 VDD.n561 VDD.n560 185
R1644 VDD.n559 VDD.n558 185
R1645 VDD.n557 VDD.n556 185
R1646 VDD.n555 VDD.n554 185
R1647 VDD.n553 VDD.n552 185
R1648 VDD.n551 VDD.n550 185
R1649 VDD.n549 VDD.n543 185
R1650 VDD.n544 VDD.n513 185
R1651 VDD.n601 VDD.n513 185
R1652 VDD.n4048 VDD.n4047 185
R1653 VDD.n285 VDD.n194 185
R1654 VDD.n284 VDD.n283 185
R1655 VDD.n282 VDD.n281 185
R1656 VDD.n280 VDD.n199 185
R1657 VDD.n276 VDD.n275 185
R1658 VDD.n274 VDD.n273 185
R1659 VDD.n272 VDD.n271 185
R1660 VDD.n270 VDD.n201 185
R1661 VDD.n266 VDD.n265 185
R1662 VDD.n264 VDD.n263 185
R1663 VDD.n262 VDD.n261 185
R1664 VDD.n260 VDD.n203 185
R1665 VDD.n256 VDD.n255 185
R1666 VDD.n254 VDD.n253 185
R1667 VDD.n252 VDD.n251 185
R1668 VDD.n250 VDD.n207 185
R1669 VDD.n246 VDD.n245 185
R1670 VDD.n244 VDD.n243 185
R1671 VDD.n242 VDD.n241 185
R1672 VDD.n240 VDD.n209 185
R1673 VDD.n236 VDD.n235 185
R1674 VDD.n234 VDD.n233 185
R1675 VDD.n232 VDD.n231 185
R1676 VDD.n230 VDD.n211 185
R1677 VDD.n226 VDD.n225 185
R1678 VDD.n224 VDD.n223 185
R1679 VDD.n222 VDD.n221 185
R1680 VDD.n220 VDD.n213 185
R1681 VDD.n216 VDD.n215 185
R1682 VDD.n4044 VDD.n179 185
R1683 VDD.n4051 VDD.n179 185
R1684 VDD.n4043 VDD.n178 185
R1685 VDD.n4052 VDD.n178 185
R1686 VDD.n4042 VDD.n4041 185
R1687 VDD.n4041 VDD.n170 185
R1688 VDD.n288 VDD.n169 185
R1689 VDD.n4058 VDD.n169 185
R1690 VDD.n4037 VDD.n168 185
R1691 VDD.n4059 VDD.n168 185
R1692 VDD.n4036 VDD.n167 185
R1693 VDD.n4060 VDD.n167 185
R1694 VDD.n4035 VDD.n4034 185
R1695 VDD.n4034 VDD.n159 185
R1696 VDD.n290 VDD.n158 185
R1697 VDD.n4066 VDD.n158 185
R1698 VDD.n4030 VDD.n157 185
R1699 VDD.n4067 VDD.n157 185
R1700 VDD.n4029 VDD.n156 185
R1701 VDD.n4068 VDD.n156 185
R1702 VDD.n4028 VDD.n4027 185
R1703 VDD.n4027 VDD.n148 185
R1704 VDD.n292 VDD.n147 185
R1705 VDD.n4074 VDD.n147 185
R1706 VDD.n4023 VDD.n146 185
R1707 VDD.n4075 VDD.n146 185
R1708 VDD.n4022 VDD.n145 185
R1709 VDD.n4076 VDD.n145 185
R1710 VDD.n4021 VDD.n4020 185
R1711 VDD.n4020 VDD.n137 185
R1712 VDD.n294 VDD.n136 185
R1713 VDD.n4082 VDD.n136 185
R1714 VDD.n4016 VDD.n135 185
R1715 VDD.n4083 VDD.n135 185
R1716 VDD.n4015 VDD.n134 185
R1717 VDD.n4084 VDD.n134 185
R1718 VDD.n4014 VDD.n4013 185
R1719 VDD.n4013 VDD.n126 185
R1720 VDD.n296 VDD.n125 185
R1721 VDD.n4090 VDD.n125 185
R1722 VDD.n4009 VDD.n124 185
R1723 VDD.n4091 VDD.n124 185
R1724 VDD.n4008 VDD.n123 185
R1725 VDD.n4092 VDD.n123 185
R1726 VDD.n4007 VDD.n4006 185
R1727 VDD.n4006 VDD.n115 185
R1728 VDD.n298 VDD.n114 185
R1729 VDD.n4098 VDD.n114 185
R1730 VDD.n4002 VDD.n113 185
R1731 VDD.n4099 VDD.n113 185
R1732 VDD.n4001 VDD.n112 185
R1733 VDD.n4100 VDD.n112 185
R1734 VDD.n4000 VDD.n3999 185
R1735 VDD.n3999 VDD.n104 185
R1736 VDD.n300 VDD.n103 185
R1737 VDD.n4106 VDD.n103 185
R1738 VDD.n3995 VDD.n102 185
R1739 VDD.n4107 VDD.n102 185
R1740 VDD.n3994 VDD.n101 185
R1741 VDD.n4108 VDD.n101 185
R1742 VDD.n3993 VDD.n3992 185
R1743 VDD.n3992 VDD.n100 185
R1744 VDD.n302 VDD.n92 185
R1745 VDD.n4114 VDD.n92 185
R1746 VDD.n3988 VDD.n91 185
R1747 VDD.n4115 VDD.n91 185
R1748 VDD.n3987 VDD.n90 185
R1749 VDD.n4116 VDD.n90 185
R1750 VDD.n3986 VDD.n3985 185
R1751 VDD.n3985 VDD.n82 185
R1752 VDD.n304 VDD.n81 185
R1753 VDD.n4122 VDD.n81 185
R1754 VDD.n3981 VDD.n80 185
R1755 VDD.n4123 VDD.n80 185
R1756 VDD.n3980 VDD.n79 185
R1757 VDD.n4124 VDD.n79 185
R1758 VDD.n3979 VDD.n3978 185
R1759 VDD.n3978 VDD.n71 185
R1760 VDD.n306 VDD.n70 185
R1761 VDD.n4130 VDD.n70 185
R1762 VDD.n3974 VDD.n69 185
R1763 VDD.n4131 VDD.n69 185
R1764 VDD.n3973 VDD.n68 185
R1765 VDD.n4132 VDD.n68 185
R1766 VDD.n3972 VDD.n3971 185
R1767 VDD.n3971 VDD.n60 185
R1768 VDD.n308 VDD.n59 185
R1769 VDD.n4138 VDD.n59 185
R1770 VDD.n3967 VDD.n58 185
R1771 VDD.n4139 VDD.n58 185
R1772 VDD.n3966 VDD.n57 185
R1773 VDD.n4140 VDD.n57 185
R1774 VDD.n3965 VDD.n3964 185
R1775 VDD.n3964 VDD.n49 185
R1776 VDD.n310 VDD.n48 185
R1777 VDD.n4146 VDD.n48 185
R1778 VDD.n3960 VDD.n47 185
R1779 VDD.n4147 VDD.n47 185
R1780 VDD.n3959 VDD.n46 185
R1781 VDD.n4148 VDD.n46 185
R1782 VDD.n3958 VDD.n3957 185
R1783 VDD.n3957 VDD.n39 185
R1784 VDD.n312 VDD.n38 185
R1785 VDD.n4154 VDD.n38 185
R1786 VDD.n3953 VDD.n37 185
R1787 VDD.n4155 VDD.n37 185
R1788 VDD.n3952 VDD.n36 185
R1789 VDD.t23 VDD.n36 185
R1790 VDD.n3951 VDD.n3950 185
R1791 VDD.n3950 VDD.n35 185
R1792 VDD.n3949 VDD.n314 185
R1793 VDD.n3949 VDD.n3948 185
R1794 VDD.n3937 VDD.n316 185
R1795 VDD.n317 VDD.n316 185
R1796 VDD.n3939 VDD.n3938 185
R1797 VDD.n3940 VDD.n3939 185
R1798 VDD.n325 VDD.n324 185
R1799 VDD.n324 VDD.n323 185
R1800 VDD.n3931 VDD.n3930 185
R1801 VDD.n3930 VDD.n3929 185
R1802 VDD.n328 VDD.n327 185
R1803 VDD.n329 VDD.n328 185
R1804 VDD.n3920 VDD.n3919 185
R1805 VDD.n3921 VDD.n3920 185
R1806 VDD.n337 VDD.n336 185
R1807 VDD.n336 VDD.n335 185
R1808 VDD.n3915 VDD.n3914 185
R1809 VDD.n3914 VDD.n3913 185
R1810 VDD.n340 VDD.n339 185
R1811 VDD.n341 VDD.n340 185
R1812 VDD.n3904 VDD.n3903 185
R1813 VDD.n3905 VDD.n3904 185
R1814 VDD.n349 VDD.n348 185
R1815 VDD.n348 VDD.n347 185
R1816 VDD.n3899 VDD.n3898 185
R1817 VDD.n3898 VDD.n3897 185
R1818 VDD.n352 VDD.n351 185
R1819 VDD.n353 VDD.n352 185
R1820 VDD.n3888 VDD.n3887 185
R1821 VDD.n3889 VDD.n3888 185
R1822 VDD.n361 VDD.n360 185
R1823 VDD.n360 VDD.n359 185
R1824 VDD.n3883 VDD.n3882 185
R1825 VDD.n3882 VDD.n3881 185
R1826 VDD.n364 VDD.n363 185
R1827 VDD.n365 VDD.n364 185
R1828 VDD.n3872 VDD.n3871 185
R1829 VDD.n3873 VDD.n3872 185
R1830 VDD.n373 VDD.n372 185
R1831 VDD.n372 VDD.n371 185
R1832 VDD.n3867 VDD.n3866 185
R1833 VDD.n3866 VDD.n3865 185
R1834 VDD.n376 VDD.n375 185
R1835 VDD.n3856 VDD.n376 185
R1836 VDD.n3855 VDD.n3854 185
R1837 VDD.n3857 VDD.n3855 185
R1838 VDD.n384 VDD.n383 185
R1839 VDD.n383 VDD.n382 185
R1840 VDD.n3850 VDD.n3849 185
R1841 VDD.n3849 VDD.n3848 185
R1842 VDD.n387 VDD.n386 185
R1843 VDD.n388 VDD.n387 185
R1844 VDD.n3839 VDD.n3838 185
R1845 VDD.n3840 VDD.n3839 185
R1846 VDD.n396 VDD.n395 185
R1847 VDD.n395 VDD.n394 185
R1848 VDD.n3834 VDD.n3833 185
R1849 VDD.n3833 VDD.n3832 185
R1850 VDD.n399 VDD.n398 185
R1851 VDD.n400 VDD.n399 185
R1852 VDD.n3823 VDD.n3822 185
R1853 VDD.n3824 VDD.n3823 185
R1854 VDD.n408 VDD.n407 185
R1855 VDD.n407 VDD.n406 185
R1856 VDD.n3818 VDD.n3817 185
R1857 VDD.n3817 VDD.n3816 185
R1858 VDD.n411 VDD.n410 185
R1859 VDD.n412 VDD.n411 185
R1860 VDD.n3807 VDD.n3806 185
R1861 VDD.n3808 VDD.n3807 185
R1862 VDD.n420 VDD.n419 185
R1863 VDD.n419 VDD.n418 185
R1864 VDD.n3802 VDD.n3801 185
R1865 VDD.n3801 VDD.n3800 185
R1866 VDD.n423 VDD.n422 185
R1867 VDD.n424 VDD.n423 185
R1868 VDD.n3791 VDD.n3790 185
R1869 VDD.n3792 VDD.n3791 185
R1870 VDD.n432 VDD.n431 185
R1871 VDD.n431 VDD.n430 185
R1872 VDD.n3786 VDD.n3785 185
R1873 VDD.n3785 VDD.n3784 185
R1874 VDD.n435 VDD.n434 185
R1875 VDD.n436 VDD.n435 185
R1876 VDD.n3775 VDD.n3774 185
R1877 VDD.n3776 VDD.n3775 185
R1878 VDD.n444 VDD.n443 185
R1879 VDD.n443 VDD.n442 185
R1880 VDD.n3770 VDD.n3769 185
R1881 VDD.n3769 VDD.n3768 185
R1882 VDD.n447 VDD.n446 185
R1883 VDD.n448 VDD.n447 185
R1884 VDD.n3759 VDD.n3758 185
R1885 VDD.n3760 VDD.n3759 185
R1886 VDD.n456 VDD.n455 185
R1887 VDD.n455 VDD.n454 185
R1888 VDD.n3754 VDD.n3753 185
R1889 VDD.n3753 VDD.n3752 185
R1890 VDD.n459 VDD.n458 185
R1891 VDD.n460 VDD.n459 185
R1892 VDD.n3743 VDD.n3742 185
R1893 VDD.n3744 VDD.n3743 185
R1894 VDD.n468 VDD.n467 185
R1895 VDD.n467 VDD.n466 185
R1896 VDD.n903 VDD.n902 185
R1897 VDD.n3135 VDD.n3133 185
R1898 VDD.n3136 VDD.n3132 185
R1899 VDD.n3136 VDD.n2976 185
R1900 VDD.n3139 VDD.n3138 185
R1901 VDD.n3140 VDD.n3131 185
R1902 VDD.n3142 VDD.n3141 185
R1903 VDD.n3144 VDD.n3130 185
R1904 VDD.n3147 VDD.n3146 185
R1905 VDD.n3148 VDD.n3129 185
R1906 VDD.n3150 VDD.n3149 185
R1907 VDD.n3152 VDD.n3128 185
R1908 VDD.n3155 VDD.n3154 185
R1909 VDD.n3156 VDD.n3127 185
R1910 VDD.n3158 VDD.n3157 185
R1911 VDD.n3160 VDD.n3126 185
R1912 VDD.n3163 VDD.n3162 185
R1913 VDD.n3164 VDD.n3123 185
R1914 VDD.n3167 VDD.n3166 185
R1915 VDD.n3169 VDD.n3122 185
R1916 VDD.n3171 VDD.n3170 185
R1917 VDD.n3170 VDD.n2976 185
R1918 VDD.n3681 VDD.n3680 185
R1919 VDD.n3683 VDD.n616 185
R1920 VDD.n3685 VDD.n3684 185
R1921 VDD.n3687 VDD.n613 185
R1922 VDD.n3689 VDD.n3688 185
R1923 VDD.n3691 VDD.n611 185
R1924 VDD.n3693 VDD.n3692 185
R1925 VDD.n3694 VDD.n610 185
R1926 VDD.n3696 VDD.n3695 185
R1927 VDD.n3698 VDD.n609 185
R1928 VDD.n3700 VDD.n3699 185
R1929 VDD.n3701 VDD.n496 185
R1930 VDD.n3703 VDD.n3702 185
R1931 VDD.n3705 VDD.n494 185
R1932 VDD.n3707 VDD.n3706 185
R1933 VDD.n3708 VDD.n493 185
R1934 VDD.n3710 VDD.n3709 185
R1935 VDD.n3712 VDD.n491 185
R1936 VDD.n3714 VDD.n3713 185
R1937 VDD.n3715 VDD.n489 185
R1938 VDD.n3679 VDD.n486 185
R1939 VDD.n3718 VDD.n486 185
R1940 VDD.n3678 VDD.n3677 185
R1941 VDD.n3677 VDD.n485 185
R1942 VDD.n3676 VDD.n618 185
R1943 VDD.n3676 VDD.n3675 185
R1944 VDD.n3442 VDD.n619 185
R1945 VDD.n620 VDD.n619 185
R1946 VDD.n3443 VDD.n627 185
R1947 VDD.n3669 VDD.n627 185
R1948 VDD.n3445 VDD.n3444 185
R1949 VDD.n3444 VDD.n626 185
R1950 VDD.n3446 VDD.n634 185
R1951 VDD.n3635 VDD.n634 185
R1952 VDD.n3448 VDD.n3447 185
R1953 VDD.n3447 VDD.n633 185
R1954 VDD.n3449 VDD.n639 185
R1955 VDD.n3629 VDD.n639 185
R1956 VDD.n3451 VDD.n3450 185
R1957 VDD.n3450 VDD.n647 185
R1958 VDD.n3452 VDD.n645 185
R1959 VDD.n3623 VDD.n645 185
R1960 VDD.n3454 VDD.n3453 185
R1961 VDD.n3453 VDD.n644 185
R1962 VDD.n3455 VDD.n652 185
R1963 VDD.n3617 VDD.n652 185
R1964 VDD.n3457 VDD.n3456 185
R1965 VDD.n3456 VDD.n651 185
R1966 VDD.n3458 VDD.n658 185
R1967 VDD.n3611 VDD.n658 185
R1968 VDD.n3460 VDD.n3459 185
R1969 VDD.n3459 VDD.n657 185
R1970 VDD.n3461 VDD.n664 185
R1971 VDD.n3605 VDD.n664 185
R1972 VDD.n3463 VDD.n3462 185
R1973 VDD.n3462 VDD.n663 185
R1974 VDD.n3464 VDD.n670 185
R1975 VDD.n3599 VDD.n670 185
R1976 VDD.n3466 VDD.n3465 185
R1977 VDD.n3465 VDD.n669 185
R1978 VDD.n3467 VDD.n676 185
R1979 VDD.n3593 VDD.n676 185
R1980 VDD.n3469 VDD.n3468 185
R1981 VDD.n3468 VDD.n675 185
R1982 VDD.n3470 VDD.n682 185
R1983 VDD.n3587 VDD.n682 185
R1984 VDD.n3472 VDD.n3471 185
R1985 VDD.n3471 VDD.n681 185
R1986 VDD.n3473 VDD.n688 185
R1987 VDD.n3581 VDD.n688 185
R1988 VDD.n3475 VDD.n3474 185
R1989 VDD.n3474 VDD.n687 185
R1990 VDD.n3476 VDD.n694 185
R1991 VDD.n3575 VDD.n694 185
R1992 VDD.n3478 VDD.n3477 185
R1993 VDD.n3477 VDD.n693 185
R1994 VDD.n3479 VDD.n700 185
R1995 VDD.n3569 VDD.n700 185
R1996 VDD.n3481 VDD.n3480 185
R1997 VDD.n3480 VDD.n699 185
R1998 VDD.n3482 VDD.n706 185
R1999 VDD.n3563 VDD.n706 185
R2000 VDD.n3484 VDD.n3483 185
R2001 VDD.n3483 VDD.n705 185
R2002 VDD.n3485 VDD.n712 185
R2003 VDD.n3557 VDD.n712 185
R2004 VDD.n3487 VDD.n3486 185
R2005 VDD.n3486 VDD.n711 185
R2006 VDD.n3488 VDD.n718 185
R2007 VDD.n3551 VDD.n718 185
R2008 VDD.n3490 VDD.n3489 185
R2009 VDD.n3489 VDD.n717 185
R2010 VDD.n3491 VDD.n724 185
R2011 VDD.n3545 VDD.n724 185
R2012 VDD.n3493 VDD.n3492 185
R2013 VDD.n3492 VDD.n723 185
R2014 VDD.n3494 VDD.n730 185
R2015 VDD.n3539 VDD.n730 185
R2016 VDD.n3496 VDD.n3495 185
R2017 VDD.n3495 VDD.n729 185
R2018 VDD.n3497 VDD.n736 185
R2019 VDD.n3533 VDD.n736 185
R2020 VDD.n3499 VDD.n3498 185
R2021 VDD.n3498 VDD.n735 185
R2022 VDD.n3500 VDD.n742 185
R2023 VDD.n3527 VDD.n742 185
R2024 VDD.n3502 VDD.n3501 185
R2025 VDD.n3501 VDD.n741 185
R2026 VDD.n3503 VDD.n748 185
R2027 VDD.n3521 VDD.n748 185
R2028 VDD.n3505 VDD.n3504 185
R2029 VDD.n3504 VDD.n747 185
R2030 VDD.n3506 VDD.n754 185
R2031 VDD.n3515 VDD.n754 185
R2032 VDD.n3507 VDD.n763 185
R2033 VDD.n763 VDD.n753 185
R2034 VDD.n3509 VDD.n3508 185
R2035 VDD.t16 VDD.n3509 185
R2036 VDD.n3441 VDD.n762 185
R2037 VDD.n762 VDD.n759 185
R2038 VDD.n3440 VDD.n3439 185
R2039 VDD.n3439 VDD.n3438 185
R2040 VDD.n765 VDD.n764 185
R2041 VDD.n766 VDD.n765 185
R2042 VDD.n3182 VDD.n772 185
R2043 VDD.n3432 VDD.n772 185
R2044 VDD.n3184 VDD.n3183 185
R2045 VDD.n3183 VDD.n781 185
R2046 VDD.n3185 VDD.n779 185
R2047 VDD.n3421 VDD.n779 185
R2048 VDD.n3187 VDD.n3186 185
R2049 VDD.n3186 VDD.n778 185
R2050 VDD.n3188 VDD.n786 185
R2051 VDD.n3415 VDD.n786 185
R2052 VDD.n3190 VDD.n3189 185
R2053 VDD.n3189 VDD.n785 185
R2054 VDD.n3191 VDD.n792 185
R2055 VDD.n3409 VDD.n792 185
R2056 VDD.n3193 VDD.n3192 185
R2057 VDD.n3192 VDD.n791 185
R2058 VDD.n3194 VDD.n797 185
R2059 VDD.n3403 VDD.n797 185
R2060 VDD.n3196 VDD.n3195 185
R2061 VDD.n3195 VDD.n805 185
R2062 VDD.n3197 VDD.n803 185
R2063 VDD.n3397 VDD.n803 185
R2064 VDD.n3199 VDD.n3198 185
R2065 VDD.n3198 VDD.n802 185
R2066 VDD.n3200 VDD.n809 185
R2067 VDD.n3391 VDD.n809 185
R2068 VDD.n3202 VDD.n3201 185
R2069 VDD.n3201 VDD.n817 185
R2070 VDD.n3203 VDD.n815 185
R2071 VDD.n3385 VDD.n815 185
R2072 VDD.n3205 VDD.n3204 185
R2073 VDD.n3204 VDD.n814 185
R2074 VDD.n3206 VDD.n822 185
R2075 VDD.n3379 VDD.n822 185
R2076 VDD.n3208 VDD.n3207 185
R2077 VDD.n3207 VDD.n821 185
R2078 VDD.n3209 VDD.n828 185
R2079 VDD.n3373 VDD.n828 185
R2080 VDD.n3211 VDD.n3210 185
R2081 VDD.n3210 VDD.n827 185
R2082 VDD.n3212 VDD.n833 185
R2083 VDD.n3367 VDD.n833 185
R2084 VDD.n3214 VDD.n3213 185
R2085 VDD.n3213 VDD.n841 185
R2086 VDD.n3215 VDD.n839 185
R2087 VDD.n3361 VDD.n839 185
R2088 VDD.n3217 VDD.n3216 185
R2089 VDD.n3216 VDD.n838 185
R2090 VDD.n3218 VDD.n846 185
R2091 VDD.n3355 VDD.n846 185
R2092 VDD.n3220 VDD.n3219 185
R2093 VDD.n3219 VDD.n845 185
R2094 VDD.n3221 VDD.n852 185
R2095 VDD.n3349 VDD.n852 185
R2096 VDD.n3223 VDD.n3222 185
R2097 VDD.n3222 VDD.n851 185
R2098 VDD.n3224 VDD.n858 185
R2099 VDD.n3343 VDD.n858 185
R2100 VDD.n3226 VDD.n3225 185
R2101 VDD.n3225 VDD.n857 185
R2102 VDD.n3227 VDD.n864 185
R2103 VDD.n3337 VDD.n864 185
R2104 VDD.n3229 VDD.n3228 185
R2105 VDD.n3228 VDD.n863 185
R2106 VDD.n3230 VDD.n870 185
R2107 VDD.n3331 VDD.n870 185
R2108 VDD.n3232 VDD.n3231 185
R2109 VDD.n3231 VDD.n869 185
R2110 VDD.n3233 VDD.n876 185
R2111 VDD.n3325 VDD.n876 185
R2112 VDD.n3235 VDD.n3234 185
R2113 VDD.n3234 VDD.n875 185
R2114 VDD.n3236 VDD.n881 185
R2115 VDD.n3319 VDD.n881 185
R2116 VDD.n3238 VDD.n3237 185
R2117 VDD.n3239 VDD.n3238 185
R2118 VDD.n3181 VDD.n887 185
R2119 VDD.n3313 VDD.n887 185
R2120 VDD.n3180 VDD.n3179 185
R2121 VDD.n3179 VDD.n886 185
R2122 VDD.n3178 VDD.n893 185
R2123 VDD.n3307 VDD.n893 185
R2124 VDD.n3177 VDD.n3176 185
R2125 VDD.n3176 VDD.n892 185
R2126 VDD.n3175 VDD.n899 185
R2127 VDD.n3301 VDD.n899 185
R2128 VDD.n3174 VDD.n3173 185
R2129 VDD.n3173 VDD.n898 185
R2130 VDD.n3172 VDD.n2977 185
R2131 VDD.n3295 VDD.n2977 185
R2132 VDD.n3297 VDD.n3296 185
R2133 VDD.n3296 VDD.n3295 185
R2134 VDD.n3298 VDD.n901 185
R2135 VDD.n901 VDD.n898 185
R2136 VDD.n3300 VDD.n3299 185
R2137 VDD.n3301 VDD.n3300 185
R2138 VDD.n891 VDD.n890 185
R2139 VDD.n892 VDD.n891 185
R2140 VDD.n3309 VDD.n3308 185
R2141 VDD.n3308 VDD.n3307 185
R2142 VDD.n3310 VDD.n889 185
R2143 VDD.n889 VDD.n886 185
R2144 VDD.n3312 VDD.n3311 185
R2145 VDD.n3313 VDD.n3312 185
R2146 VDD.n880 VDD.n879 185
R2147 VDD.n3239 VDD.n880 185
R2148 VDD.n3321 VDD.n3320 185
R2149 VDD.n3320 VDD.n3319 185
R2150 VDD.n3322 VDD.n878 185
R2151 VDD.n878 VDD.n875 185
R2152 VDD.n3324 VDD.n3323 185
R2153 VDD.n3325 VDD.n3324 185
R2154 VDD.n868 VDD.n867 185
R2155 VDD.n869 VDD.n868 185
R2156 VDD.n3333 VDD.n3332 185
R2157 VDD.n3332 VDD.n3331 185
R2158 VDD.n3334 VDD.n866 185
R2159 VDD.n866 VDD.n863 185
R2160 VDD.n3336 VDD.n3335 185
R2161 VDD.n3337 VDD.n3336 185
R2162 VDD.n856 VDD.n855 185
R2163 VDD.n857 VDD.n856 185
R2164 VDD.n3345 VDD.n3344 185
R2165 VDD.n3344 VDD.n3343 185
R2166 VDD.n3346 VDD.n854 185
R2167 VDD.n854 VDD.n851 185
R2168 VDD.n3348 VDD.n3347 185
R2169 VDD.n3349 VDD.n3348 185
R2170 VDD.n844 VDD.n843 185
R2171 VDD.n845 VDD.n844 185
R2172 VDD.n3357 VDD.n3356 185
R2173 VDD.n3356 VDD.n3355 185
R2174 VDD.n3358 VDD.n842 185
R2175 VDD.n842 VDD.n838 185
R2176 VDD.n3360 VDD.n3359 185
R2177 VDD.n3361 VDD.n3360 185
R2178 VDD.n832 VDD.n831 185
R2179 VDD.n841 VDD.n832 185
R2180 VDD.n3369 VDD.n3368 185
R2181 VDD.n3368 VDD.n3367 185
R2182 VDD.n3370 VDD.n830 185
R2183 VDD.n830 VDD.n827 185
R2184 VDD.n3372 VDD.n3371 185
R2185 VDD.n3373 VDD.n3372 185
R2186 VDD.n820 VDD.n819 185
R2187 VDD.n821 VDD.n820 185
R2188 VDD.n3381 VDD.n3380 185
R2189 VDD.n3380 VDD.n3379 185
R2190 VDD.n3382 VDD.n818 185
R2191 VDD.n818 VDD.n814 185
R2192 VDD.n3384 VDD.n3383 185
R2193 VDD.n3385 VDD.n3384 185
R2194 VDD.n808 VDD.n807 185
R2195 VDD.n817 VDD.n808 185
R2196 VDD.n3393 VDD.n3392 185
R2197 VDD.n3392 VDD.n3391 185
R2198 VDD.n3394 VDD.n806 185
R2199 VDD.n806 VDD.n802 185
R2200 VDD.n3396 VDD.n3395 185
R2201 VDD.n3397 VDD.n3396 185
R2202 VDD.n796 VDD.n795 185
R2203 VDD.n805 VDD.n796 185
R2204 VDD.n3405 VDD.n3404 185
R2205 VDD.n3404 VDD.n3403 185
R2206 VDD.n3406 VDD.n794 185
R2207 VDD.n794 VDD.n791 185
R2208 VDD.n3408 VDD.n3407 185
R2209 VDD.n3409 VDD.n3408 185
R2210 VDD.n784 VDD.n783 185
R2211 VDD.n785 VDD.n784 185
R2212 VDD.n3417 VDD.n3416 185
R2213 VDD.n3416 VDD.n3415 185
R2214 VDD.n3418 VDD.n782 185
R2215 VDD.n782 VDD.n778 185
R2216 VDD.n3420 VDD.n3419 185
R2217 VDD.n3421 VDD.n3420 185
R2218 VDD.n771 VDD.n770 185
R2219 VDD.n781 VDD.n771 185
R2220 VDD.n3434 VDD.n3433 185
R2221 VDD.n3433 VDD.n3432 185
R2222 VDD.n3435 VDD.n769 185
R2223 VDD.n769 VDD.n766 185
R2224 VDD.n3437 VDD.n3436 185
R2225 VDD.n3438 VDD.n3437 185
R2226 VDD.n758 VDD.n757 185
R2227 VDD.n759 VDD.n758 185
R2228 VDD.n3511 VDD.n3510 185
R2229 VDD.n3510 VDD.t16 185
R2230 VDD.n3512 VDD.n756 185
R2231 VDD.n756 VDD.n753 185
R2232 VDD.n3514 VDD.n3513 185
R2233 VDD.n3515 VDD.n3514 185
R2234 VDD.n746 VDD.n745 185
R2235 VDD.n747 VDD.n746 185
R2236 VDD.n3523 VDD.n3522 185
R2237 VDD.n3522 VDD.n3521 185
R2238 VDD.n3524 VDD.n744 185
R2239 VDD.n744 VDD.n741 185
R2240 VDD.n3526 VDD.n3525 185
R2241 VDD.n3527 VDD.n3526 185
R2242 VDD.n734 VDD.n733 185
R2243 VDD.n735 VDD.n734 185
R2244 VDD.n3535 VDD.n3534 185
R2245 VDD.n3534 VDD.n3533 185
R2246 VDD.n3536 VDD.n732 185
R2247 VDD.n732 VDD.n729 185
R2248 VDD.n3538 VDD.n3537 185
R2249 VDD.n3539 VDD.n3538 185
R2250 VDD.n722 VDD.n721 185
R2251 VDD.n723 VDD.n722 185
R2252 VDD.n3547 VDD.n3546 185
R2253 VDD.n3546 VDD.n3545 185
R2254 VDD.n3548 VDD.n720 185
R2255 VDD.n720 VDD.n717 185
R2256 VDD.n3550 VDD.n3549 185
R2257 VDD.n3551 VDD.n3550 185
R2258 VDD.n710 VDD.n709 185
R2259 VDD.n711 VDD.n710 185
R2260 VDD.n3559 VDD.n3558 185
R2261 VDD.n3558 VDD.n3557 185
R2262 VDD.n3560 VDD.n708 185
R2263 VDD.n708 VDD.n705 185
R2264 VDD.n3562 VDD.n3561 185
R2265 VDD.n3563 VDD.n3562 185
R2266 VDD.n698 VDD.n697 185
R2267 VDD.n699 VDD.n698 185
R2268 VDD.n3571 VDD.n3570 185
R2269 VDD.n3570 VDD.n3569 185
R2270 VDD.n3572 VDD.n696 185
R2271 VDD.n696 VDD.n693 185
R2272 VDD.n3574 VDD.n3573 185
R2273 VDD.n3575 VDD.n3574 185
R2274 VDD.n686 VDD.n685 185
R2275 VDD.n687 VDD.n686 185
R2276 VDD.n3583 VDD.n3582 185
R2277 VDD.n3582 VDD.n3581 185
R2278 VDD.n3584 VDD.n684 185
R2279 VDD.n684 VDD.n681 185
R2280 VDD.n3586 VDD.n3585 185
R2281 VDD.n3587 VDD.n3586 185
R2282 VDD.n674 VDD.n673 185
R2283 VDD.n675 VDD.n674 185
R2284 VDD.n3595 VDD.n3594 185
R2285 VDD.n3594 VDD.n3593 185
R2286 VDD.n3596 VDD.n672 185
R2287 VDD.n672 VDD.n669 185
R2288 VDD.n3598 VDD.n3597 185
R2289 VDD.n3599 VDD.n3598 185
R2290 VDD.n662 VDD.n661 185
R2291 VDD.n663 VDD.n662 185
R2292 VDD.n3607 VDD.n3606 185
R2293 VDD.n3606 VDD.n3605 185
R2294 VDD.n3608 VDD.n660 185
R2295 VDD.n660 VDD.n657 185
R2296 VDD.n3610 VDD.n3609 185
R2297 VDD.n3611 VDD.n3610 185
R2298 VDD.n650 VDD.n649 185
R2299 VDD.n651 VDD.n650 185
R2300 VDD.n3619 VDD.n3618 185
R2301 VDD.n3618 VDD.n3617 185
R2302 VDD.n3620 VDD.n648 185
R2303 VDD.n648 VDD.n644 185
R2304 VDD.n3622 VDD.n3621 185
R2305 VDD.n3623 VDD.n3622 185
R2306 VDD.n638 VDD.n637 185
R2307 VDD.n647 VDD.n638 185
R2308 VDD.n3631 VDD.n3630 185
R2309 VDD.n3630 VDD.n3629 185
R2310 VDD.n3632 VDD.n636 185
R2311 VDD.n636 VDD.n633 185
R2312 VDD.n3634 VDD.n3633 185
R2313 VDD.n3635 VDD.n3634 185
R2314 VDD.n625 VDD.n624 185
R2315 VDD.n626 VDD.n625 185
R2316 VDD.n3671 VDD.n3670 185
R2317 VDD.n3670 VDD.n3669 185
R2318 VDD.n3672 VDD.n623 185
R2319 VDD.n623 VDD.n620 185
R2320 VDD.n3674 VDD.n3673 185
R2321 VDD.n3675 VDD.n3674 185
R2322 VDD.n490 VDD.n488 185
R2323 VDD.n488 VDD.n485 185
R2324 VDD.n3717 VDD.n3716 185
R2325 VDD.n3718 VDD.n3717 185
R2326 VDD.n2965 VDD.n933 185
R2327 VDD.n933 VDD.n904 185
R2328 VDD.n2967 VDD.n2966 185
R2329 VDD.n2968 VDD.n2967 185
R2330 VDD.n934 VDD.n932 185
R2331 VDD.n932 VDD.n929 185
R2332 VDD.n2916 VDD.n2915 185
R2333 VDD.n2917 VDD.n2916 185
R2334 VDD.n2914 VDD.n942 185
R2335 VDD.n942 VDD.n939 185
R2336 VDD.n2913 VDD.n2912 185
R2337 VDD.n2912 VDD.n2911 185
R2338 VDD.n944 VDD.n943 185
R2339 VDD.n945 VDD.n944 185
R2340 VDD.n2858 VDD.n2857 185
R2341 VDD.n2859 VDD.n2858 185
R2342 VDD.n2856 VDD.n954 185
R2343 VDD.n960 VDD.n954 185
R2344 VDD.n2855 VDD.n2854 185
R2345 VDD.n2854 VDD.n2853 185
R2346 VDD.n956 VDD.n955 185
R2347 VDD.n957 VDD.n956 185
R2348 VDD.n2846 VDD.n2845 185
R2349 VDD.n2847 VDD.n2846 185
R2350 VDD.n2844 VDD.n967 185
R2351 VDD.n967 VDD.n964 185
R2352 VDD.n2843 VDD.n2842 185
R2353 VDD.n2842 VDD.n2841 185
R2354 VDD.n969 VDD.n968 185
R2355 VDD.n970 VDD.n969 185
R2356 VDD.n2834 VDD.n2833 185
R2357 VDD.n2835 VDD.n2834 185
R2358 VDD.n2832 VDD.n979 185
R2359 VDD.n979 VDD.n976 185
R2360 VDD.n2831 VDD.n2830 185
R2361 VDD.n2830 VDD.n2829 185
R2362 VDD.n981 VDD.n980 185
R2363 VDD.n982 VDD.n981 185
R2364 VDD.n2822 VDD.n2821 185
R2365 VDD.n2823 VDD.n2822 185
R2366 VDD.n2820 VDD.n991 185
R2367 VDD.n991 VDD.n988 185
R2368 VDD.n2819 VDD.n2818 185
R2369 VDD.n2818 VDD.n2817 185
R2370 VDD.n993 VDD.n992 185
R2371 VDD.n994 VDD.n993 185
R2372 VDD.n2810 VDD.n2809 185
R2373 VDD.n2811 VDD.n2810 185
R2374 VDD.n2808 VDD.n1002 185
R2375 VDD.n1008 VDD.n1002 185
R2376 VDD.n2807 VDD.n2806 185
R2377 VDD.n2806 VDD.n2805 185
R2378 VDD.n1004 VDD.n1003 185
R2379 VDD.n1005 VDD.n1004 185
R2380 VDD.n2798 VDD.n2797 185
R2381 VDD.n2799 VDD.n2798 185
R2382 VDD.n2796 VDD.n1015 185
R2383 VDD.n1015 VDD.n1012 185
R2384 VDD.n2795 VDD.n2794 185
R2385 VDD.n2794 VDD.n2793 185
R2386 VDD.n1017 VDD.n1016 185
R2387 VDD.n1018 VDD.n1017 185
R2388 VDD.n2786 VDD.n2785 185
R2389 VDD.n2787 VDD.n2786 185
R2390 VDD.n2784 VDD.n1026 185
R2391 VDD.n1032 VDD.n1026 185
R2392 VDD.n2783 VDD.n2782 185
R2393 VDD.n2782 VDD.n2781 185
R2394 VDD.n1028 VDD.n1027 185
R2395 VDD.n1029 VDD.n1028 185
R2396 VDD.n2774 VDD.n2773 185
R2397 VDD.n2775 VDD.n2774 185
R2398 VDD.n2772 VDD.n1038 185
R2399 VDD.n1044 VDD.n1038 185
R2400 VDD.n2771 VDD.n2770 185
R2401 VDD.n2770 VDD.n2769 185
R2402 VDD.n1040 VDD.n1039 185
R2403 VDD.n1041 VDD.n1040 185
R2404 VDD.n2762 VDD.n2761 185
R2405 VDD.n2763 VDD.n2762 185
R2406 VDD.n2760 VDD.n1051 185
R2407 VDD.n1051 VDD.n1048 185
R2408 VDD.n2759 VDD.n2758 185
R2409 VDD.n2758 VDD.n2757 185
R2410 VDD.n1053 VDD.n1052 185
R2411 VDD.n1054 VDD.n1053 185
R2412 VDD.n2750 VDD.n2749 185
R2413 VDD.n2751 VDD.n2750 185
R2414 VDD.n2748 VDD.n1062 185
R2415 VDD.n1068 VDD.n1062 185
R2416 VDD.n2747 VDD.n2746 185
R2417 VDD.n2746 VDD.n2745 185
R2418 VDD.n1064 VDD.n1063 185
R2419 VDD.n1065 VDD.n1064 185
R2420 VDD.n2738 VDD.n2737 185
R2421 VDD.n2739 VDD.n2738 185
R2422 VDD.n2736 VDD.n1074 185
R2423 VDD.n1074 VDD.t25 185
R2424 VDD.n2735 VDD.n2734 185
R2425 VDD.n2734 VDD.n2733 185
R2426 VDD.n1076 VDD.n1075 185
R2427 VDD.n1077 VDD.n1076 185
R2428 VDD.n2726 VDD.n2725 185
R2429 VDD.n2727 VDD.n2726 185
R2430 VDD.n2724 VDD.n1086 185
R2431 VDD.n1086 VDD.n1083 185
R2432 VDD.n2723 VDD.n2722 185
R2433 VDD.n2722 VDD.n2721 185
R2434 VDD.n1088 VDD.n1087 185
R2435 VDD.n1089 VDD.n1088 185
R2436 VDD.n2714 VDD.n2713 185
R2437 VDD.n2715 VDD.n2714 185
R2438 VDD.n2712 VDD.n1098 185
R2439 VDD.n1098 VDD.n1095 185
R2440 VDD.n2711 VDD.n2710 185
R2441 VDD.n2710 VDD.n2709 185
R2442 VDD.n1100 VDD.n1099 185
R2443 VDD.n1101 VDD.n1100 185
R2444 VDD.n2702 VDD.n2701 185
R2445 VDD.n2703 VDD.n2702 185
R2446 VDD.n2700 VDD.n1110 185
R2447 VDD.n1110 VDD.n1107 185
R2448 VDD.n2699 VDD.n2698 185
R2449 VDD.n2698 VDD.n2697 185
R2450 VDD.n1112 VDD.n1111 185
R2451 VDD.n1113 VDD.n1112 185
R2452 VDD.n2690 VDD.n2689 185
R2453 VDD.n2691 VDD.n2690 185
R2454 VDD.n2688 VDD.n1122 185
R2455 VDD.n1122 VDD.n1119 185
R2456 VDD.n2687 VDD.n2686 185
R2457 VDD.n2686 VDD.n2685 185
R2458 VDD.n1124 VDD.n1123 185
R2459 VDD.n1125 VDD.n1124 185
R2460 VDD.n2678 VDD.n2677 185
R2461 VDD.n2679 VDD.n2678 185
R2462 VDD.n2676 VDD.n1134 185
R2463 VDD.n1134 VDD.n1131 185
R2464 VDD.n2675 VDD.n2674 185
R2465 VDD.n2674 VDD.n2673 185
R2466 VDD.n1136 VDD.n1135 185
R2467 VDD.n1137 VDD.n1136 185
R2468 VDD.n2666 VDD.n2665 185
R2469 VDD.n2667 VDD.n2666 185
R2470 VDD.n2664 VDD.n1146 185
R2471 VDD.n1146 VDD.n1143 185
R2472 VDD.n2663 VDD.n2662 185
R2473 VDD.n2662 VDD.n2661 185
R2474 VDD.n1148 VDD.n1147 185
R2475 VDD.n1149 VDD.n1148 185
R2476 VDD.n2654 VDD.n2653 185
R2477 VDD.n2655 VDD.n2654 185
R2478 VDD.n2652 VDD.n1158 185
R2479 VDD.n1158 VDD.n1155 185
R2480 VDD.n2651 VDD.n2650 185
R2481 VDD.n2650 VDD.n2649 185
R2482 VDD.n1160 VDD.n1159 185
R2483 VDD.n1161 VDD.n1160 185
R2484 VDD.n2642 VDD.n2641 185
R2485 VDD.n2643 VDD.n2642 185
R2486 VDD.n2640 VDD.n1170 185
R2487 VDD.n1170 VDD.n1167 185
R2488 VDD.n2639 VDD.n2638 185
R2489 VDD.n2638 VDD.n2637 185
R2490 VDD.n1172 VDD.n1171 185
R2491 VDD.n1173 VDD.n1172 185
R2492 VDD.n2630 VDD.n2629 185
R2493 VDD.n2631 VDD.n2630 185
R2494 VDD.n2628 VDD.n1182 185
R2495 VDD.n1182 VDD.n1179 185
R2496 VDD.n2627 VDD.n2626 185
R2497 VDD.n2626 VDD.n2625 185
R2498 VDD.n1184 VDD.n1183 185
R2499 VDD.n1185 VDD.n1184 185
R2500 VDD.n2618 VDD.n2617 185
R2501 VDD.n2619 VDD.n2618 185
R2502 VDD.n2616 VDD.n1193 185
R2503 VDD.n2468 VDD.n1193 185
R2504 VDD.n2615 VDD.n2614 185
R2505 VDD.n2614 VDD.n2613 185
R2506 VDD.n1195 VDD.n1194 185
R2507 VDD.n1196 VDD.n1195 185
R2508 VDD.n2606 VDD.n2605 185
R2509 VDD.n2607 VDD.n2606 185
R2510 VDD.n2604 VDD.n1205 185
R2511 VDD.n1205 VDD.n1202 185
R2512 VDD.n2603 VDD.n2602 185
R2513 VDD.n2602 VDD.n2601 185
R2514 VDD.n1207 VDD.n1206 185
R2515 VDD.n1208 VDD.n1207 185
R2516 VDD.n2594 VDD.n2593 185
R2517 VDD.n2595 VDD.n2594 185
R2518 VDD.n2592 VDD.n1217 185
R2519 VDD.n1217 VDD.n1214 185
R2520 VDD.n2925 VDD.n2924 185
R2521 VDD.n2927 VDD.n2926 185
R2522 VDD.n2929 VDD.n2928 185
R2523 VDD.n2932 VDD.n2931 185
R2524 VDD.n2934 VDD.n2933 185
R2525 VDD.n2936 VDD.n2935 185
R2526 VDD.n2938 VDD.n2937 185
R2527 VDD.n2940 VDD.n2939 185
R2528 VDD.n2942 VDD.n2941 185
R2529 VDD.n2944 VDD.n2943 185
R2530 VDD.n2946 VDD.n2945 185
R2531 VDD.n2948 VDD.n2947 185
R2532 VDD.n2950 VDD.n2949 185
R2533 VDD.n2952 VDD.n2951 185
R2534 VDD.n2954 VDD.n2953 185
R2535 VDD.n2956 VDD.n2955 185
R2536 VDD.n2958 VDD.n2957 185
R2537 VDD.n2960 VDD.n2959 185
R2538 VDD.n2962 VDD.n2961 185
R2539 VDD.n2964 VDD.n2963 185
R2540 VDD.n2923 VDD.n2922 185
R2541 VDD.n2923 VDD.n904 185
R2542 VDD.n2921 VDD.n930 185
R2543 VDD.n2968 VDD.n930 185
R2544 VDD.n2920 VDD.n2919 185
R2545 VDD.n2919 VDD.n929 185
R2546 VDD.n2918 VDD.n937 185
R2547 VDD.n2918 VDD.n2917 185
R2548 VDD.n2341 VDD.n938 185
R2549 VDD.n939 VDD.n938 185
R2550 VDD.n2342 VDD.n946 185
R2551 VDD.n2911 VDD.n946 185
R2552 VDD.n2344 VDD.n2343 185
R2553 VDD.n2343 VDD.n945 185
R2554 VDD.n2345 VDD.n952 185
R2555 VDD.n2859 VDD.n952 185
R2556 VDD.n2347 VDD.n2346 185
R2557 VDD.n2346 VDD.n960 185
R2558 VDD.n2348 VDD.n958 185
R2559 VDD.n2853 VDD.n958 185
R2560 VDD.n2350 VDD.n2349 185
R2561 VDD.n2349 VDD.n957 185
R2562 VDD.n2351 VDD.n965 185
R2563 VDD.n2847 VDD.n965 185
R2564 VDD.n2353 VDD.n2352 185
R2565 VDD.n2352 VDD.n964 185
R2566 VDD.n2354 VDD.n971 185
R2567 VDD.n2841 VDD.n971 185
R2568 VDD.n2356 VDD.n2355 185
R2569 VDD.n2355 VDD.n970 185
R2570 VDD.n2357 VDD.n977 185
R2571 VDD.n2835 VDD.n977 185
R2572 VDD.n2359 VDD.n2358 185
R2573 VDD.n2358 VDD.n976 185
R2574 VDD.n2360 VDD.n983 185
R2575 VDD.n2829 VDD.n983 185
R2576 VDD.n2362 VDD.n2361 185
R2577 VDD.n2361 VDD.n982 185
R2578 VDD.n2363 VDD.n989 185
R2579 VDD.n2823 VDD.n989 185
R2580 VDD.n2365 VDD.n2364 185
R2581 VDD.n2364 VDD.n988 185
R2582 VDD.n2366 VDD.n995 185
R2583 VDD.n2817 VDD.n995 185
R2584 VDD.n2368 VDD.n2367 185
R2585 VDD.n2367 VDD.n994 185
R2586 VDD.n2369 VDD.n1000 185
R2587 VDD.n2811 VDD.n1000 185
R2588 VDD.n2371 VDD.n2370 185
R2589 VDD.n2370 VDD.n1008 185
R2590 VDD.n2372 VDD.n1006 185
R2591 VDD.n2805 VDD.n1006 185
R2592 VDD.n2374 VDD.n2373 185
R2593 VDD.n2373 VDD.n1005 185
R2594 VDD.n2375 VDD.n1013 185
R2595 VDD.n2799 VDD.n1013 185
R2596 VDD.n2377 VDD.n2376 185
R2597 VDD.n2376 VDD.n1012 185
R2598 VDD.n2378 VDD.n1019 185
R2599 VDD.n2793 VDD.n1019 185
R2600 VDD.n2380 VDD.n2379 185
R2601 VDD.n2379 VDD.n1018 185
R2602 VDD.n2381 VDD.n1024 185
R2603 VDD.n2787 VDD.n1024 185
R2604 VDD.n2383 VDD.n2382 185
R2605 VDD.n2382 VDD.n1032 185
R2606 VDD.n2384 VDD.n1030 185
R2607 VDD.n2781 VDD.n1030 185
R2608 VDD.n2386 VDD.n2385 185
R2609 VDD.n2385 VDD.n1029 185
R2610 VDD.n2387 VDD.n1036 185
R2611 VDD.n2775 VDD.n1036 185
R2612 VDD.n2389 VDD.n2388 185
R2613 VDD.n2388 VDD.n1044 185
R2614 VDD.n2390 VDD.n1042 185
R2615 VDD.n2769 VDD.n1042 185
R2616 VDD.n2392 VDD.n2391 185
R2617 VDD.n2391 VDD.n1041 185
R2618 VDD.n2393 VDD.n1049 185
R2619 VDD.n2763 VDD.n1049 185
R2620 VDD.n2395 VDD.n2394 185
R2621 VDD.n2394 VDD.n1048 185
R2622 VDD.n2396 VDD.n1055 185
R2623 VDD.n2757 VDD.n1055 185
R2624 VDD.n2398 VDD.n2397 185
R2625 VDD.n2397 VDD.n1054 185
R2626 VDD.n2399 VDD.n1060 185
R2627 VDD.n2751 VDD.n1060 185
R2628 VDD.n2401 VDD.n2400 185
R2629 VDD.n2400 VDD.n1068 185
R2630 VDD.n2402 VDD.n1066 185
R2631 VDD.n2745 VDD.n1066 185
R2632 VDD.n2404 VDD.n2403 185
R2633 VDD.n2403 VDD.n1065 185
R2634 VDD.n2405 VDD.n1072 185
R2635 VDD.n2739 VDD.n1072 185
R2636 VDD.n2407 VDD.n2406 185
R2637 VDD.n2406 VDD.t25 185
R2638 VDD.n2408 VDD.n1078 185
R2639 VDD.n2733 VDD.n1078 185
R2640 VDD.n2410 VDD.n2409 185
R2641 VDD.n2409 VDD.n1077 185
R2642 VDD.n2411 VDD.n1084 185
R2643 VDD.n2727 VDD.n1084 185
R2644 VDD.n2413 VDD.n2412 185
R2645 VDD.n2412 VDD.n1083 185
R2646 VDD.n2414 VDD.n1090 185
R2647 VDD.n2721 VDD.n1090 185
R2648 VDD.n2416 VDD.n2415 185
R2649 VDD.n2415 VDD.n1089 185
R2650 VDD.n2417 VDD.n1096 185
R2651 VDD.n2715 VDD.n1096 185
R2652 VDD.n2419 VDD.n2418 185
R2653 VDD.n2418 VDD.n1095 185
R2654 VDD.n2420 VDD.n1102 185
R2655 VDD.n2709 VDD.n1102 185
R2656 VDD.n2422 VDD.n2421 185
R2657 VDD.n2421 VDD.n1101 185
R2658 VDD.n2423 VDD.n1108 185
R2659 VDD.n2703 VDD.n1108 185
R2660 VDD.n2425 VDD.n2424 185
R2661 VDD.n2424 VDD.n1107 185
R2662 VDD.n2426 VDD.n1114 185
R2663 VDD.n2697 VDD.n1114 185
R2664 VDD.n2428 VDD.n2427 185
R2665 VDD.n2427 VDD.n1113 185
R2666 VDD.n2429 VDD.n1120 185
R2667 VDD.n2691 VDD.n1120 185
R2668 VDD.n2431 VDD.n2430 185
R2669 VDD.n2430 VDD.n1119 185
R2670 VDD.n2432 VDD.n1126 185
R2671 VDD.n2685 VDD.n1126 185
R2672 VDD.n2434 VDD.n2433 185
R2673 VDD.n2433 VDD.n1125 185
R2674 VDD.n2435 VDD.n1132 185
R2675 VDD.n2679 VDD.n1132 185
R2676 VDD.n2437 VDD.n2436 185
R2677 VDD.n2436 VDD.n1131 185
R2678 VDD.n2438 VDD.n1138 185
R2679 VDD.n2673 VDD.n1138 185
R2680 VDD.n2440 VDD.n2439 185
R2681 VDD.n2439 VDD.n1137 185
R2682 VDD.n2441 VDD.n1144 185
R2683 VDD.n2667 VDD.n1144 185
R2684 VDD.n2443 VDD.n2442 185
R2685 VDD.n2442 VDD.n1143 185
R2686 VDD.n2444 VDD.n1150 185
R2687 VDD.n2661 VDD.n1150 185
R2688 VDD.n2446 VDD.n2445 185
R2689 VDD.n2445 VDD.n1149 185
R2690 VDD.n2447 VDD.n1156 185
R2691 VDD.n2655 VDD.n1156 185
R2692 VDD.n2449 VDD.n2448 185
R2693 VDD.n2448 VDD.n1155 185
R2694 VDD.n2450 VDD.n1162 185
R2695 VDD.n2649 VDD.n1162 185
R2696 VDD.n2452 VDD.n2451 185
R2697 VDD.n2451 VDD.n1161 185
R2698 VDD.n2453 VDD.n1168 185
R2699 VDD.n2643 VDD.n1168 185
R2700 VDD.n2455 VDD.n2454 185
R2701 VDD.n2454 VDD.n1167 185
R2702 VDD.n2456 VDD.n1174 185
R2703 VDD.n2637 VDD.n1174 185
R2704 VDD.n2458 VDD.n2457 185
R2705 VDD.n2457 VDD.n1173 185
R2706 VDD.n2459 VDD.n1180 185
R2707 VDD.n2631 VDD.n1180 185
R2708 VDD.n2461 VDD.n2460 185
R2709 VDD.n2460 VDD.n1179 185
R2710 VDD.n2462 VDD.n1186 185
R2711 VDD.n2625 VDD.n1186 185
R2712 VDD.n2464 VDD.n2463 185
R2713 VDD.n2463 VDD.n1185 185
R2714 VDD.n2465 VDD.n1191 185
R2715 VDD.n2619 VDD.n1191 185
R2716 VDD.n2467 VDD.n2466 185
R2717 VDD.n2468 VDD.n2467 185
R2718 VDD.n2340 VDD.n1197 185
R2719 VDD.n2613 VDD.n1197 185
R2720 VDD.n2339 VDD.n2338 185
R2721 VDD.n2338 VDD.n1196 185
R2722 VDD.n2337 VDD.n1203 185
R2723 VDD.n2607 VDD.n1203 185
R2724 VDD.n2336 VDD.n2335 185
R2725 VDD.n2335 VDD.n1202 185
R2726 VDD.n2334 VDD.n1209 185
R2727 VDD.n2601 VDD.n1209 185
R2728 VDD.n2333 VDD.n2332 185
R2729 VDD.n2332 VDD.n1208 185
R2730 VDD.n2331 VDD.n1215 185
R2731 VDD.n2595 VDD.n1215 185
R2732 VDD.n2330 VDD.n2329 185
R2733 VDD.n2329 VDD.n1214 185
R2734 VDD.n2591 VDD.n2590 185
R2735 VDD.n1219 VDD.n1218 185
R2736 VDD.n2587 VDD.n2586 185
R2737 VDD.n2588 VDD.n2587 185
R2738 VDD.n2585 VDD.n1239 185
R2739 VDD.n2584 VDD.n2583 185
R2740 VDD.n2582 VDD.n2581 185
R2741 VDD.n2580 VDD.n2579 185
R2742 VDD.n2578 VDD.n2577 185
R2743 VDD.n2576 VDD.n2575 185
R2744 VDD.n2574 VDD.n2573 185
R2745 VDD.n2311 VDD.n1240 185
R2746 VDD.n2313 VDD.n2312 185
R2747 VDD.n2315 VDD.n2314 185
R2748 VDD.n2317 VDD.n2316 185
R2749 VDD.n2319 VDD.n2318 185
R2750 VDD.n2321 VDD.n2320 185
R2751 VDD.n2323 VDD.n2322 185
R2752 VDD.n2325 VDD.n2324 185
R2753 VDD.n2327 VDD.n2326 185
R2754 VDD.n2328 VDD.n1228 185
R2755 VDD.n2588 VDD.n1228 185
R2756 VDD.n221 VDD.n220 146.341
R2757 VDD.n225 VDD.n224 146.341
R2758 VDD.n231 VDD.n230 146.341
R2759 VDD.n235 VDD.n234 146.341
R2760 VDD.n241 VDD.n240 146.341
R2761 VDD.n245 VDD.n244 146.341
R2762 VDD.n251 VDD.n250 146.341
R2763 VDD.n255 VDD.n254 146.341
R2764 VDD.n261 VDD.n260 146.341
R2765 VDD.n265 VDD.n264 146.341
R2766 VDD.n271 VDD.n270 146.341
R2767 VDD.n275 VDD.n274 146.341
R2768 VDD.n281 VDD.n280 146.341
R2769 VDD.n283 VDD.n194 146.341
R2770 VDD.n3743 VDD.n467 146.341
R2771 VDD.n3743 VDD.n459 146.341
R2772 VDD.n3753 VDD.n459 146.341
R2773 VDD.n3753 VDD.n455 146.341
R2774 VDD.n3759 VDD.n455 146.341
R2775 VDD.n3759 VDD.n447 146.341
R2776 VDD.n3769 VDD.n447 146.341
R2777 VDD.n3769 VDD.n443 146.341
R2778 VDD.n3775 VDD.n443 146.341
R2779 VDD.n3775 VDD.n435 146.341
R2780 VDD.n3785 VDD.n435 146.341
R2781 VDD.n3785 VDD.n431 146.341
R2782 VDD.n3791 VDD.n431 146.341
R2783 VDD.n3791 VDD.n423 146.341
R2784 VDD.n3801 VDD.n423 146.341
R2785 VDD.n3801 VDD.n419 146.341
R2786 VDD.n3807 VDD.n419 146.341
R2787 VDD.n3807 VDD.n411 146.341
R2788 VDD.n3817 VDD.n411 146.341
R2789 VDD.n3817 VDD.n407 146.341
R2790 VDD.n3823 VDD.n407 146.341
R2791 VDD.n3823 VDD.n399 146.341
R2792 VDD.n3833 VDD.n399 146.341
R2793 VDD.n3833 VDD.n395 146.341
R2794 VDD.n3839 VDD.n395 146.341
R2795 VDD.n3839 VDD.n387 146.341
R2796 VDD.n3849 VDD.n387 146.341
R2797 VDD.n3849 VDD.n383 146.341
R2798 VDD.n3855 VDD.n383 146.341
R2799 VDD.n3855 VDD.n376 146.341
R2800 VDD.n3866 VDD.n376 146.341
R2801 VDD.n3866 VDD.n372 146.341
R2802 VDD.n3872 VDD.n372 146.341
R2803 VDD.n3872 VDD.n364 146.341
R2804 VDD.n3882 VDD.n364 146.341
R2805 VDD.n3882 VDD.n360 146.341
R2806 VDD.n3888 VDD.n360 146.341
R2807 VDD.n3888 VDD.n352 146.341
R2808 VDD.n3898 VDD.n352 146.341
R2809 VDD.n3898 VDD.n348 146.341
R2810 VDD.n3904 VDD.n348 146.341
R2811 VDD.n3904 VDD.n340 146.341
R2812 VDD.n3914 VDD.n340 146.341
R2813 VDD.n3914 VDD.n336 146.341
R2814 VDD.n3920 VDD.n336 146.341
R2815 VDD.n3920 VDD.n328 146.341
R2816 VDD.n3930 VDD.n328 146.341
R2817 VDD.n3930 VDD.n324 146.341
R2818 VDD.n3939 VDD.n324 146.341
R2819 VDD.n3939 VDD.n316 146.341
R2820 VDD.n3949 VDD.n316 146.341
R2821 VDD.n3950 VDD.n3949 146.341
R2822 VDD.n3950 VDD.n36 146.341
R2823 VDD.n37 VDD.n36 146.341
R2824 VDD.n38 VDD.n37 146.341
R2825 VDD.n3957 VDD.n38 146.341
R2826 VDD.n3957 VDD.n46 146.341
R2827 VDD.n47 VDD.n46 146.341
R2828 VDD.n48 VDD.n47 146.341
R2829 VDD.n3964 VDD.n48 146.341
R2830 VDD.n3964 VDD.n57 146.341
R2831 VDD.n58 VDD.n57 146.341
R2832 VDD.n59 VDD.n58 146.341
R2833 VDD.n3971 VDD.n59 146.341
R2834 VDD.n3971 VDD.n68 146.341
R2835 VDD.n69 VDD.n68 146.341
R2836 VDD.n70 VDD.n69 146.341
R2837 VDD.n3978 VDD.n70 146.341
R2838 VDD.n3978 VDD.n79 146.341
R2839 VDD.n80 VDD.n79 146.341
R2840 VDD.n81 VDD.n80 146.341
R2841 VDD.n3985 VDD.n81 146.341
R2842 VDD.n3985 VDD.n90 146.341
R2843 VDD.n91 VDD.n90 146.341
R2844 VDD.n92 VDD.n91 146.341
R2845 VDD.n3992 VDD.n92 146.341
R2846 VDD.n3992 VDD.n101 146.341
R2847 VDD.n102 VDD.n101 146.341
R2848 VDD.n103 VDD.n102 146.341
R2849 VDD.n3999 VDD.n103 146.341
R2850 VDD.n3999 VDD.n112 146.341
R2851 VDD.n113 VDD.n112 146.341
R2852 VDD.n114 VDD.n113 146.341
R2853 VDD.n4006 VDD.n114 146.341
R2854 VDD.n4006 VDD.n123 146.341
R2855 VDD.n124 VDD.n123 146.341
R2856 VDD.n125 VDD.n124 146.341
R2857 VDD.n4013 VDD.n125 146.341
R2858 VDD.n4013 VDD.n134 146.341
R2859 VDD.n135 VDD.n134 146.341
R2860 VDD.n136 VDD.n135 146.341
R2861 VDD.n4020 VDD.n136 146.341
R2862 VDD.n4020 VDD.n145 146.341
R2863 VDD.n146 VDD.n145 146.341
R2864 VDD.n147 VDD.n146 146.341
R2865 VDD.n4027 VDD.n147 146.341
R2866 VDD.n4027 VDD.n156 146.341
R2867 VDD.n157 VDD.n156 146.341
R2868 VDD.n158 VDD.n157 146.341
R2869 VDD.n4034 VDD.n158 146.341
R2870 VDD.n4034 VDD.n167 146.341
R2871 VDD.n168 VDD.n167 146.341
R2872 VDD.n169 VDD.n168 146.341
R2873 VDD.n4041 VDD.n169 146.341
R2874 VDD.n4041 VDD.n178 146.341
R2875 VDD.n179 VDD.n178 146.341
R2876 VDD.n600 VDD.n499 146.341
R2877 VDD.n600 VDD.n514 146.341
R2878 VDD.n596 VDD.n595 146.341
R2879 VDD.n592 VDD.n591 146.341
R2880 VDD.n588 VDD.n587 146.341
R2881 VDD.n584 VDD.n583 146.341
R2882 VDD.n580 VDD.n579 146.341
R2883 VDD.n576 VDD.n575 146.341
R2884 VDD.n572 VDD.n571 146.341
R2885 VDD.n568 VDD.n567 146.341
R2886 VDD.n564 VDD.n563 146.341
R2887 VDD.n560 VDD.n559 146.341
R2888 VDD.n556 VDD.n555 146.341
R2889 VDD.n552 VDD.n551 146.341
R2890 VDD.n543 VDD.n513 146.341
R2891 VDD.n3745 VDD.n465 146.341
R2892 VDD.n3745 VDD.n461 146.341
R2893 VDD.n3751 VDD.n461 146.341
R2894 VDD.n3751 VDD.n453 146.341
R2895 VDD.n3761 VDD.n453 146.341
R2896 VDD.n3761 VDD.n449 146.341
R2897 VDD.n3767 VDD.n449 146.341
R2898 VDD.n3767 VDD.n441 146.341
R2899 VDD.n3777 VDD.n441 146.341
R2900 VDD.n3777 VDD.n437 146.341
R2901 VDD.n3783 VDD.n437 146.341
R2902 VDD.n3783 VDD.n429 146.341
R2903 VDD.n3793 VDD.n429 146.341
R2904 VDD.n3793 VDD.n425 146.341
R2905 VDD.n3799 VDD.n425 146.341
R2906 VDD.n3799 VDD.n417 146.341
R2907 VDD.n3809 VDD.n417 146.341
R2908 VDD.n3809 VDD.n413 146.341
R2909 VDD.n3815 VDD.n413 146.341
R2910 VDD.n3815 VDD.n405 146.341
R2911 VDD.n3825 VDD.n405 146.341
R2912 VDD.n3825 VDD.n401 146.341
R2913 VDD.n3831 VDD.n401 146.341
R2914 VDD.n3831 VDD.n393 146.341
R2915 VDD.n3841 VDD.n393 146.341
R2916 VDD.n3841 VDD.n389 146.341
R2917 VDD.n3847 VDD.n389 146.341
R2918 VDD.n3847 VDD.n381 146.341
R2919 VDD.n3858 VDD.n381 146.341
R2920 VDD.n3858 VDD.n377 146.341
R2921 VDD.n3864 VDD.n377 146.341
R2922 VDD.n3864 VDD.n370 146.341
R2923 VDD.n3874 VDD.n370 146.341
R2924 VDD.n3874 VDD.n366 146.341
R2925 VDD.n3880 VDD.n366 146.341
R2926 VDD.n3880 VDD.n358 146.341
R2927 VDD.n3890 VDD.n358 146.341
R2928 VDD.n3890 VDD.n354 146.341
R2929 VDD.n3896 VDD.n354 146.341
R2930 VDD.n3896 VDD.n346 146.341
R2931 VDD.n3906 VDD.n346 146.341
R2932 VDD.n3906 VDD.n342 146.341
R2933 VDD.n3912 VDD.n342 146.341
R2934 VDD.n3912 VDD.n334 146.341
R2935 VDD.n3922 VDD.n334 146.341
R2936 VDD.n3922 VDD.n330 146.341
R2937 VDD.n3928 VDD.n330 146.341
R2938 VDD.n3928 VDD.n322 146.341
R2939 VDD.n3941 VDD.n322 146.341
R2940 VDD.n3941 VDD.n318 146.341
R2941 VDD.n3947 VDD.n318 146.341
R2942 VDD.n3947 VDD.n33 146.341
R2943 VDD.n4156 VDD.n33 146.341
R2944 VDD.n4156 VDD.n34 146.341
R2945 VDD.n4153 VDD.n34 146.341
R2946 VDD.n4153 VDD.n40 146.341
R2947 VDD.n4149 VDD.n40 146.341
R2948 VDD.n4149 VDD.n45 146.341
R2949 VDD.n4145 VDD.n45 146.341
R2950 VDD.n4145 VDD.n50 146.341
R2951 VDD.n4141 VDD.n50 146.341
R2952 VDD.n4141 VDD.n56 146.341
R2953 VDD.n4137 VDD.n56 146.341
R2954 VDD.n4137 VDD.n61 146.341
R2955 VDD.n4133 VDD.n61 146.341
R2956 VDD.n4133 VDD.n67 146.341
R2957 VDD.n4129 VDD.n67 146.341
R2958 VDD.n4129 VDD.n72 146.341
R2959 VDD.n4125 VDD.n72 146.341
R2960 VDD.n4125 VDD.n78 146.341
R2961 VDD.n4121 VDD.n78 146.341
R2962 VDD.n4121 VDD.n83 146.341
R2963 VDD.n4117 VDD.n83 146.341
R2964 VDD.n4117 VDD.n89 146.341
R2965 VDD.n4113 VDD.n89 146.341
R2966 VDD.n4113 VDD.n93 146.341
R2967 VDD.n4109 VDD.n93 146.341
R2968 VDD.n4109 VDD.n99 146.341
R2969 VDD.n4105 VDD.n99 146.341
R2970 VDD.n4105 VDD.n105 146.341
R2971 VDD.n4101 VDD.n105 146.341
R2972 VDD.n4101 VDD.n111 146.341
R2973 VDD.n4097 VDD.n111 146.341
R2974 VDD.n4097 VDD.n116 146.341
R2975 VDD.n4093 VDD.n116 146.341
R2976 VDD.n4093 VDD.n122 146.341
R2977 VDD.n4089 VDD.n122 146.341
R2978 VDD.n4089 VDD.n127 146.341
R2979 VDD.n4085 VDD.n127 146.341
R2980 VDD.n4085 VDD.n133 146.341
R2981 VDD.n4081 VDD.n133 146.341
R2982 VDD.n4081 VDD.n138 146.341
R2983 VDD.n4077 VDD.n138 146.341
R2984 VDD.n4077 VDD.n144 146.341
R2985 VDD.n4073 VDD.n144 146.341
R2986 VDD.n4073 VDD.n149 146.341
R2987 VDD.n4069 VDD.n149 146.341
R2988 VDD.n4069 VDD.n155 146.341
R2989 VDD.n4065 VDD.n155 146.341
R2990 VDD.n4065 VDD.n160 146.341
R2991 VDD.n4061 VDD.n160 146.341
R2992 VDD.n4061 VDD.n166 146.341
R2993 VDD.n4057 VDD.n166 146.341
R2994 VDD.n4057 VDD.n171 146.341
R2995 VDD.n4053 VDD.n171 146.341
R2996 VDD.n4053 VDD.n177 146.341
R2997 VDD.n1245 VDD.n1244 146.341
R2998 VDD.n1288 VDD.n1248 146.341
R2999 VDD.n1250 VDD.n1249 146.341
R3000 VDD.n1291 VDD.n1253 146.341
R3001 VDD.n1255 VDD.n1254 146.341
R3002 VDD.n1294 VDD.n1258 146.341
R3003 VDD.n1262 VDD.n1261 146.341
R3004 VDD.n1297 VDD.n1265 146.341
R3005 VDD.n1267 VDD.n1266 146.341
R3006 VDD.n1300 VDD.n1270 146.341
R3007 VDD.n1272 VDD.n1271 146.341
R3008 VDD.n1303 VDD.n1275 146.341
R3009 VDD.n1277 VDD.n1276 146.341
R3010 VDD.n1306 VDD.n1280 146.341
R3011 VDD.n1739 VDD.n1620 146.341
R3012 VDD.n1739 VDD.n1616 146.341
R3013 VDD.n1745 VDD.n1616 146.341
R3014 VDD.n1745 VDD.n1608 146.341
R3015 VDD.n1755 VDD.n1608 146.341
R3016 VDD.n1755 VDD.n1604 146.341
R3017 VDD.n1761 VDD.n1604 146.341
R3018 VDD.n1761 VDD.n1596 146.341
R3019 VDD.n1771 VDD.n1596 146.341
R3020 VDD.n1771 VDD.n1592 146.341
R3021 VDD.n1777 VDD.n1592 146.341
R3022 VDD.n1777 VDD.n1584 146.341
R3023 VDD.n1787 VDD.n1584 146.341
R3024 VDD.n1787 VDD.n1580 146.341
R3025 VDD.n1793 VDD.n1580 146.341
R3026 VDD.n1793 VDD.n1572 146.341
R3027 VDD.n1803 VDD.n1572 146.341
R3028 VDD.n1803 VDD.n1568 146.341
R3029 VDD.n1809 VDD.n1568 146.341
R3030 VDD.n1809 VDD.n1560 146.341
R3031 VDD.n1819 VDD.n1560 146.341
R3032 VDD.n1819 VDD.n1556 146.341
R3033 VDD.n1825 VDD.n1556 146.341
R3034 VDD.n1825 VDD.n1548 146.341
R3035 VDD.n1835 VDD.n1548 146.341
R3036 VDD.n1835 VDD.n1544 146.341
R3037 VDD.n1841 VDD.n1544 146.341
R3038 VDD.n1841 VDD.n1535 146.341
R3039 VDD.n1851 VDD.n1535 146.341
R3040 VDD.n1851 VDD.n1531 146.341
R3041 VDD.n1857 VDD.n1531 146.341
R3042 VDD.n1857 VDD.n1524 146.341
R3043 VDD.n1867 VDD.n1524 146.341
R3044 VDD.n1867 VDD.n1520 146.341
R3045 VDD.n1873 VDD.n1520 146.341
R3046 VDD.n1873 VDD.n1512 146.341
R3047 VDD.n1883 VDD.n1512 146.341
R3048 VDD.n1883 VDD.n1508 146.341
R3049 VDD.n1889 VDD.n1508 146.341
R3050 VDD.n1889 VDD.n1500 146.341
R3051 VDD.n1899 VDD.n1500 146.341
R3052 VDD.n1899 VDD.n1496 146.341
R3053 VDD.n1905 VDD.n1496 146.341
R3054 VDD.n1905 VDD.n1488 146.341
R3055 VDD.n1915 VDD.n1488 146.341
R3056 VDD.n1915 VDD.n1484 146.341
R3057 VDD.n1921 VDD.n1484 146.341
R3058 VDD.n1921 VDD.n1476 146.341
R3059 VDD.n1931 VDD.n1476 146.341
R3060 VDD.n1931 VDD.n1472 146.341
R3061 VDD.n1937 VDD.n1472 146.341
R3062 VDD.n1937 VDD.n1464 146.341
R3063 VDD.n1960 VDD.n1464 146.341
R3064 VDD.n1960 VDD.n1460 146.341
R3065 VDD.n1966 VDD.n1460 146.341
R3066 VDD.n1966 VDD.n1452 146.341
R3067 VDD.n1976 VDD.n1452 146.341
R3068 VDD.n1976 VDD.n1448 146.341
R3069 VDD.n1982 VDD.n1448 146.341
R3070 VDD.n1982 VDD.n1440 146.341
R3071 VDD.n1992 VDD.n1440 146.341
R3072 VDD.n1992 VDD.n1436 146.341
R3073 VDD.n1998 VDD.n1436 146.341
R3074 VDD.n1998 VDD.n1429 146.341
R3075 VDD.n2009 VDD.n1429 146.341
R3076 VDD.n2009 VDD.n1425 146.341
R3077 VDD.n2015 VDD.n1425 146.341
R3078 VDD.n2015 VDD.n1417 146.341
R3079 VDD.n2025 VDD.n1417 146.341
R3080 VDD.n2025 VDD.n1413 146.341
R3081 VDD.n2031 VDD.n1413 146.341
R3082 VDD.n2031 VDD.n1405 146.341
R3083 VDD.n2041 VDD.n1405 146.341
R3084 VDD.n2041 VDD.n1401 146.341
R3085 VDD.n2047 VDD.n1401 146.341
R3086 VDD.n2047 VDD.n1393 146.341
R3087 VDD.n2057 VDD.n1393 146.341
R3088 VDD.n2057 VDD.n1389 146.341
R3089 VDD.n2063 VDD.n1389 146.341
R3090 VDD.n2063 VDD.n1381 146.341
R3091 VDD.n2073 VDD.n1381 146.341
R3092 VDD.n2073 VDD.n1377 146.341
R3093 VDD.n2079 VDD.n1377 146.341
R3094 VDD.n2079 VDD.n1368 146.341
R3095 VDD.n2089 VDD.n1368 146.341
R3096 VDD.n2089 VDD.n1364 146.341
R3097 VDD.n2095 VDD.n1364 146.341
R3098 VDD.n2095 VDD.n1357 146.341
R3099 VDD.n2105 VDD.n1357 146.341
R3100 VDD.n2105 VDD.n1353 146.341
R3101 VDD.n2111 VDD.n1353 146.341
R3102 VDD.n2111 VDD.n1345 146.341
R3103 VDD.n2121 VDD.n1345 146.341
R3104 VDD.n2121 VDD.n1341 146.341
R3105 VDD.n2127 VDD.n1341 146.341
R3106 VDD.n2127 VDD.n1333 146.341
R3107 VDD.n2137 VDD.n1333 146.341
R3108 VDD.n2137 VDD.n1328 146.341
R3109 VDD.n2144 VDD.n1328 146.341
R3110 VDD.n2144 VDD.n1321 146.341
R3111 VDD.n2155 VDD.n1321 146.341
R3112 VDD.n2156 VDD.n2155 146.341
R3113 VDD.n2156 VDD.n1316 146.341
R3114 VDD.n2511 VDD.n1316 146.341
R3115 VDD.n2511 VDD.n1284 146.341
R3116 VDD.n2523 VDD.n1284 146.341
R3117 VDD.n1728 VDD.n1626 146.341
R3118 VDD.n1728 VDD.n1641 146.341
R3119 VDD.n1645 VDD.n1644 146.341
R3120 VDD.n1647 VDD.n1646 146.341
R3121 VDD.n1651 VDD.n1650 146.341
R3122 VDD.n1653 VDD.n1652 146.341
R3123 VDD.n1707 VDD.n1656 146.341
R3124 VDD.n1658 VDD.n1657 146.341
R3125 VDD.n1662 VDD.n1661 146.341
R3126 VDD.n1664 VDD.n1663 146.341
R3127 VDD.n1668 VDD.n1667 146.341
R3128 VDD.n1670 VDD.n1669 146.341
R3129 VDD.n1674 VDD.n1673 146.341
R3130 VDD.n1676 VDD.n1675 146.341
R3131 VDD.n1679 VDD.n1640 146.341
R3132 VDD.n1737 VDD.n1622 146.341
R3133 VDD.n1737 VDD.n1614 146.341
R3134 VDD.n1747 VDD.n1614 146.341
R3135 VDD.n1747 VDD.n1610 146.341
R3136 VDD.n1753 VDD.n1610 146.341
R3137 VDD.n1753 VDD.n1602 146.341
R3138 VDD.n1763 VDD.n1602 146.341
R3139 VDD.n1763 VDD.n1598 146.341
R3140 VDD.n1769 VDD.n1598 146.341
R3141 VDD.n1769 VDD.n1590 146.341
R3142 VDD.n1779 VDD.n1590 146.341
R3143 VDD.n1779 VDD.n1586 146.341
R3144 VDD.n1785 VDD.n1586 146.341
R3145 VDD.n1785 VDD.n1578 146.341
R3146 VDD.n1795 VDD.n1578 146.341
R3147 VDD.n1795 VDD.n1574 146.341
R3148 VDD.n1801 VDD.n1574 146.341
R3149 VDD.n1801 VDD.n1566 146.341
R3150 VDD.n1811 VDD.n1566 146.341
R3151 VDD.n1811 VDD.n1562 146.341
R3152 VDD.n1817 VDD.n1562 146.341
R3153 VDD.n1817 VDD.n1554 146.341
R3154 VDD.n1827 VDD.n1554 146.341
R3155 VDD.n1827 VDD.n1550 146.341
R3156 VDD.n1833 VDD.n1550 146.341
R3157 VDD.n1833 VDD.n1542 146.341
R3158 VDD.n1843 VDD.n1542 146.341
R3159 VDD.n1843 VDD.n1538 146.341
R3160 VDD.n1849 VDD.n1538 146.341
R3161 VDD.n1849 VDD.n1530 146.341
R3162 VDD.n1859 VDD.n1530 146.341
R3163 VDD.n1859 VDD.n1526 146.341
R3164 VDD.n1865 VDD.n1526 146.341
R3165 VDD.n1865 VDD.n1518 146.341
R3166 VDD.n1875 VDD.n1518 146.341
R3167 VDD.n1875 VDD.n1514 146.341
R3168 VDD.n1881 VDD.n1514 146.341
R3169 VDD.n1881 VDD.n1506 146.341
R3170 VDD.n1891 VDD.n1506 146.341
R3171 VDD.n1891 VDD.n1502 146.341
R3172 VDD.n1897 VDD.n1502 146.341
R3173 VDD.n1897 VDD.n1494 146.341
R3174 VDD.n1907 VDD.n1494 146.341
R3175 VDD.n1907 VDD.n1490 146.341
R3176 VDD.n1913 VDD.n1490 146.341
R3177 VDD.n1913 VDD.n1482 146.341
R3178 VDD.n1923 VDD.n1482 146.341
R3179 VDD.n1923 VDD.n1478 146.341
R3180 VDD.n1929 VDD.n1478 146.341
R3181 VDD.n1929 VDD.n1470 146.341
R3182 VDD.n1939 VDD.n1470 146.341
R3183 VDD.n1939 VDD.n1466 146.341
R3184 VDD.n1959 VDD.n1466 146.341
R3185 VDD.n1959 VDD.n1458 146.341
R3186 VDD.n1968 VDD.n1458 146.341
R3187 VDD.n1968 VDD.n1454 146.341
R3188 VDD.n1974 VDD.n1454 146.341
R3189 VDD.n1974 VDD.n1446 146.341
R3190 VDD.n1984 VDD.n1446 146.341
R3191 VDD.n1984 VDD.n1442 146.341
R3192 VDD.n1990 VDD.n1442 146.341
R3193 VDD.n1990 VDD.n1434 146.341
R3194 VDD.n2001 VDD.n1434 146.341
R3195 VDD.n2001 VDD.n1430 146.341
R3196 VDD.n2007 VDD.n1430 146.341
R3197 VDD.n2007 VDD.n1423 146.341
R3198 VDD.n2017 VDD.n1423 146.341
R3199 VDD.n2017 VDD.n1419 146.341
R3200 VDD.n2023 VDD.n1419 146.341
R3201 VDD.n2023 VDD.n1411 146.341
R3202 VDD.n2033 VDD.n1411 146.341
R3203 VDD.n2033 VDD.n1407 146.341
R3204 VDD.n2039 VDD.n1407 146.341
R3205 VDD.n2039 VDD.n1399 146.341
R3206 VDD.n2049 VDD.n1399 146.341
R3207 VDD.n2049 VDD.n1395 146.341
R3208 VDD.n2055 VDD.n1395 146.341
R3209 VDD.n2055 VDD.n1387 146.341
R3210 VDD.n2065 VDD.n1387 146.341
R3211 VDD.n2065 VDD.n1383 146.341
R3212 VDD.n2071 VDD.n1383 146.341
R3213 VDD.n2071 VDD.n1375 146.341
R3214 VDD.n2081 VDD.n1375 146.341
R3215 VDD.n2081 VDD.n1371 146.341
R3216 VDD.n2087 VDD.n1371 146.341
R3217 VDD.n2087 VDD.n1363 146.341
R3218 VDD.n2097 VDD.n1363 146.341
R3219 VDD.n2097 VDD.n1359 146.341
R3220 VDD.n2103 VDD.n1359 146.341
R3221 VDD.n2103 VDD.n1351 146.341
R3222 VDD.n2113 VDD.n1351 146.341
R3223 VDD.n2113 VDD.n1347 146.341
R3224 VDD.n2119 VDD.n1347 146.341
R3225 VDD.n2119 VDD.n1339 146.341
R3226 VDD.n2129 VDD.n1339 146.341
R3227 VDD.n2129 VDD.n1335 146.341
R3228 VDD.n2135 VDD.n1335 146.341
R3229 VDD.n2135 VDD.n1326 146.341
R3230 VDD.n2147 VDD.n1326 146.341
R3231 VDD.n2147 VDD.n1322 146.341
R3232 VDD.n2153 VDD.n1322 146.341
R3233 VDD.n2153 VDD.n1313 146.341
R3234 VDD.n2514 VDD.n1313 146.341
R3235 VDD.n2514 VDD.n1314 146.341
R3236 VDD.n1314 VDD.n1309 146.341
R3237 VDD.n2521 VDD.n1309 146.341
R3238 VDD.n2976 VDD.n2975 126.784
R3239 VDD.n9 VDD.n7 125.144
R3240 VDD.n2 VDD.n0 125.144
R3241 VDD.n9 VDD.n8 123.32
R3242 VDD.n11 VDD.n10 123.32
R3243 VDD.n13 VDD.n12 123.32
R3244 VDD.n6 VDD.n5 123.32
R3245 VDD.n4 VDD.n3 123.32
R3246 VDD.n2 VDD.n1 123.32
R3247 VDD.n2309 VDD.t127 119.436
R3248 VDD.n936 VDD.t118 119.436
R3249 VDD.n2989 VDD.t91 119.436
R3250 VDD.n615 VDD.t80 119.436
R3251 VDD.n3125 VDD.t111 119.436
R3252 VDD.n480 VDD.t115 119.436
R3253 VDD.n2180 VDD.t121 119.436
R3254 VDD.n2864 VDD.t76 119.436
R3255 VDD.n1260 VDD.t84 117.724
R3256 VDD.n1282 VDD.t99 117.724
R3257 VDD.n1682 VDD.t101 117.724
R3258 VDD.n1709 VDD.t87 117.724
R3259 VDD.n528 VDD.t95 117.724
R3260 VDD.n546 VDD.t108 117.724
R3261 VDD.n196 VDD.t125 117.724
R3262 VDD.n206 VDD.t106 117.724
R3263 VDD.n1260 VDD.n1259 108.995
R3264 VDD.n1282 VDD.n1281 108.995
R3265 VDD.n1682 VDD.n1681 108.995
R3266 VDD.n1709 VDD.n1708 108.995
R3267 VDD.n528 VDD.n527 108.995
R3268 VDD.n546 VDD.n545 108.995
R3269 VDD.n196 VDD.n195 108.995
R3270 VDD.n206 VDD.n205 108.995
R3271 VDD.n3296 VDD.n901 99.5127
R3272 VDD.n3300 VDD.n901 99.5127
R3273 VDD.n3300 VDD.n891 99.5127
R3274 VDD.n3308 VDD.n891 99.5127
R3275 VDD.n3308 VDD.n889 99.5127
R3276 VDD.n3312 VDD.n889 99.5127
R3277 VDD.n3312 VDD.n880 99.5127
R3278 VDD.n3320 VDD.n880 99.5127
R3279 VDD.n3320 VDD.n878 99.5127
R3280 VDD.n3324 VDD.n878 99.5127
R3281 VDD.n3324 VDD.n868 99.5127
R3282 VDD.n3332 VDD.n868 99.5127
R3283 VDD.n3332 VDD.n866 99.5127
R3284 VDD.n3336 VDD.n866 99.5127
R3285 VDD.n3336 VDD.n856 99.5127
R3286 VDD.n3344 VDD.n856 99.5127
R3287 VDD.n3344 VDD.n854 99.5127
R3288 VDD.n3348 VDD.n854 99.5127
R3289 VDD.n3348 VDD.n844 99.5127
R3290 VDD.n3356 VDD.n844 99.5127
R3291 VDD.n3356 VDD.n842 99.5127
R3292 VDD.n3360 VDD.n842 99.5127
R3293 VDD.n3360 VDD.n832 99.5127
R3294 VDD.n3368 VDD.n832 99.5127
R3295 VDD.n3368 VDD.n830 99.5127
R3296 VDD.n3372 VDD.n830 99.5127
R3297 VDD.n3372 VDD.n820 99.5127
R3298 VDD.n3380 VDD.n820 99.5127
R3299 VDD.n3380 VDD.n818 99.5127
R3300 VDD.n3384 VDD.n818 99.5127
R3301 VDD.n3384 VDD.n808 99.5127
R3302 VDD.n3392 VDD.n808 99.5127
R3303 VDD.n3392 VDD.n806 99.5127
R3304 VDD.n3396 VDD.n806 99.5127
R3305 VDD.n3396 VDD.n796 99.5127
R3306 VDD.n3404 VDD.n796 99.5127
R3307 VDD.n3404 VDD.n794 99.5127
R3308 VDD.n3408 VDD.n794 99.5127
R3309 VDD.n3408 VDD.n784 99.5127
R3310 VDD.n3416 VDD.n784 99.5127
R3311 VDD.n3416 VDD.n782 99.5127
R3312 VDD.n3420 VDD.n782 99.5127
R3313 VDD.n3420 VDD.n771 99.5127
R3314 VDD.n3433 VDD.n771 99.5127
R3315 VDD.n3433 VDD.n769 99.5127
R3316 VDD.n3437 VDD.n769 99.5127
R3317 VDD.n3437 VDD.n758 99.5127
R3318 VDD.n3510 VDD.n758 99.5127
R3319 VDD.n3510 VDD.n756 99.5127
R3320 VDD.n3514 VDD.n756 99.5127
R3321 VDD.n3514 VDD.n746 99.5127
R3322 VDD.n3522 VDD.n746 99.5127
R3323 VDD.n3522 VDD.n744 99.5127
R3324 VDD.n3526 VDD.n744 99.5127
R3325 VDD.n3526 VDD.n734 99.5127
R3326 VDD.n3534 VDD.n734 99.5127
R3327 VDD.n3534 VDD.n732 99.5127
R3328 VDD.n3538 VDD.n732 99.5127
R3329 VDD.n3538 VDD.n722 99.5127
R3330 VDD.n3546 VDD.n722 99.5127
R3331 VDD.n3546 VDD.n720 99.5127
R3332 VDD.n3550 VDD.n720 99.5127
R3333 VDD.n3550 VDD.n710 99.5127
R3334 VDD.n3558 VDD.n710 99.5127
R3335 VDD.n3558 VDD.n708 99.5127
R3336 VDD.n3562 VDD.n708 99.5127
R3337 VDD.n3562 VDD.n698 99.5127
R3338 VDD.n3570 VDD.n698 99.5127
R3339 VDD.n3570 VDD.n696 99.5127
R3340 VDD.n3574 VDD.n696 99.5127
R3341 VDD.n3574 VDD.n686 99.5127
R3342 VDD.n3582 VDD.n686 99.5127
R3343 VDD.n3582 VDD.n684 99.5127
R3344 VDD.n3586 VDD.n684 99.5127
R3345 VDD.n3586 VDD.n674 99.5127
R3346 VDD.n3594 VDD.n674 99.5127
R3347 VDD.n3594 VDD.n672 99.5127
R3348 VDD.n3598 VDD.n672 99.5127
R3349 VDD.n3598 VDD.n662 99.5127
R3350 VDD.n3606 VDD.n662 99.5127
R3351 VDD.n3606 VDD.n660 99.5127
R3352 VDD.n3610 VDD.n660 99.5127
R3353 VDD.n3610 VDD.n650 99.5127
R3354 VDD.n3618 VDD.n650 99.5127
R3355 VDD.n3618 VDD.n648 99.5127
R3356 VDD.n3622 VDD.n648 99.5127
R3357 VDD.n3622 VDD.n638 99.5127
R3358 VDD.n3630 VDD.n638 99.5127
R3359 VDD.n3630 VDD.n636 99.5127
R3360 VDD.n3634 VDD.n636 99.5127
R3361 VDD.n3634 VDD.n625 99.5127
R3362 VDD.n3670 VDD.n625 99.5127
R3363 VDD.n3670 VDD.n623 99.5127
R3364 VDD.n3674 VDD.n623 99.5127
R3365 VDD.n3674 VDD.n488 99.5127
R3366 VDD.n3717 VDD.n488 99.5127
R3367 VDD.n3713 VDD.n3712 99.5127
R3368 VDD.n3710 VDD.n493 99.5127
R3369 VDD.n3706 VDD.n3705 99.5127
R3370 VDD.n3703 VDD.n496 99.5127
R3371 VDD.n3699 VDD.n3698 99.5127
R3372 VDD.n3696 VDD.n610 99.5127
R3373 VDD.n3692 VDD.n3691 99.5127
R3374 VDD.n3689 VDD.n613 99.5127
R3375 VDD.n3684 VDD.n3683 99.5127
R3376 VDD.n3173 VDD.n2977 99.5127
R3377 VDD.n3173 VDD.n899 99.5127
R3378 VDD.n3176 VDD.n899 99.5127
R3379 VDD.n3176 VDD.n893 99.5127
R3380 VDD.n3179 VDD.n893 99.5127
R3381 VDD.n3179 VDD.n887 99.5127
R3382 VDD.n3238 VDD.n887 99.5127
R3383 VDD.n3238 VDD.n881 99.5127
R3384 VDD.n3234 VDD.n881 99.5127
R3385 VDD.n3234 VDD.n876 99.5127
R3386 VDD.n3231 VDD.n876 99.5127
R3387 VDD.n3231 VDD.n870 99.5127
R3388 VDD.n3228 VDD.n870 99.5127
R3389 VDD.n3228 VDD.n864 99.5127
R3390 VDD.n3225 VDD.n864 99.5127
R3391 VDD.n3225 VDD.n858 99.5127
R3392 VDD.n3222 VDD.n858 99.5127
R3393 VDD.n3222 VDD.n852 99.5127
R3394 VDD.n3219 VDD.n852 99.5127
R3395 VDD.n3219 VDD.n846 99.5127
R3396 VDD.n3216 VDD.n846 99.5127
R3397 VDD.n3216 VDD.n839 99.5127
R3398 VDD.n3213 VDD.n839 99.5127
R3399 VDD.n3213 VDD.n833 99.5127
R3400 VDD.n3210 VDD.n833 99.5127
R3401 VDD.n3210 VDD.n828 99.5127
R3402 VDD.n3207 VDD.n828 99.5127
R3403 VDD.n3207 VDD.n822 99.5127
R3404 VDD.n3204 VDD.n822 99.5127
R3405 VDD.n3204 VDD.n815 99.5127
R3406 VDD.n3201 VDD.n815 99.5127
R3407 VDD.n3201 VDD.n809 99.5127
R3408 VDD.n3198 VDD.n809 99.5127
R3409 VDD.n3198 VDD.n803 99.5127
R3410 VDD.n3195 VDD.n803 99.5127
R3411 VDD.n3195 VDD.n797 99.5127
R3412 VDD.n3192 VDD.n797 99.5127
R3413 VDD.n3192 VDD.n792 99.5127
R3414 VDD.n3189 VDD.n792 99.5127
R3415 VDD.n3189 VDD.n786 99.5127
R3416 VDD.n3186 VDD.n786 99.5127
R3417 VDD.n3186 VDD.n779 99.5127
R3418 VDD.n3183 VDD.n779 99.5127
R3419 VDD.n3183 VDD.n772 99.5127
R3420 VDD.n772 VDD.n765 99.5127
R3421 VDD.n3439 VDD.n765 99.5127
R3422 VDD.n3439 VDD.n762 99.5127
R3423 VDD.n3509 VDD.n762 99.5127
R3424 VDD.n3509 VDD.n763 99.5127
R3425 VDD.n763 VDD.n754 99.5127
R3426 VDD.n3504 VDD.n754 99.5127
R3427 VDD.n3504 VDD.n748 99.5127
R3428 VDD.n3501 VDD.n748 99.5127
R3429 VDD.n3501 VDD.n742 99.5127
R3430 VDD.n3498 VDD.n742 99.5127
R3431 VDD.n3498 VDD.n736 99.5127
R3432 VDD.n3495 VDD.n736 99.5127
R3433 VDD.n3495 VDD.n730 99.5127
R3434 VDD.n3492 VDD.n730 99.5127
R3435 VDD.n3492 VDD.n724 99.5127
R3436 VDD.n3489 VDD.n724 99.5127
R3437 VDD.n3489 VDD.n718 99.5127
R3438 VDD.n3486 VDD.n718 99.5127
R3439 VDD.n3486 VDD.n712 99.5127
R3440 VDD.n3483 VDD.n712 99.5127
R3441 VDD.n3483 VDD.n706 99.5127
R3442 VDD.n3480 VDD.n706 99.5127
R3443 VDD.n3480 VDD.n700 99.5127
R3444 VDD.n3477 VDD.n700 99.5127
R3445 VDD.n3477 VDD.n694 99.5127
R3446 VDD.n3474 VDD.n694 99.5127
R3447 VDD.n3474 VDD.n688 99.5127
R3448 VDD.n3471 VDD.n688 99.5127
R3449 VDD.n3471 VDD.n682 99.5127
R3450 VDD.n3468 VDD.n682 99.5127
R3451 VDD.n3468 VDD.n676 99.5127
R3452 VDD.n3465 VDD.n676 99.5127
R3453 VDD.n3465 VDD.n670 99.5127
R3454 VDD.n3462 VDD.n670 99.5127
R3455 VDD.n3462 VDD.n664 99.5127
R3456 VDD.n3459 VDD.n664 99.5127
R3457 VDD.n3459 VDD.n658 99.5127
R3458 VDD.n3456 VDD.n658 99.5127
R3459 VDD.n3456 VDD.n652 99.5127
R3460 VDD.n3453 VDD.n652 99.5127
R3461 VDD.n3453 VDD.n645 99.5127
R3462 VDD.n3450 VDD.n645 99.5127
R3463 VDD.n3450 VDD.n639 99.5127
R3464 VDD.n3447 VDD.n639 99.5127
R3465 VDD.n3447 VDD.n634 99.5127
R3466 VDD.n3444 VDD.n634 99.5127
R3467 VDD.n3444 VDD.n627 99.5127
R3468 VDD.n627 VDD.n619 99.5127
R3469 VDD.n3676 VDD.n619 99.5127
R3470 VDD.n3677 VDD.n3676 99.5127
R3471 VDD.n3677 VDD.n486 99.5127
R3472 VDD.n3136 VDD.n3135 99.5127
R3473 VDD.n3138 VDD.n3136 99.5127
R3474 VDD.n3142 VDD.n3131 99.5127
R3475 VDD.n3146 VDD.n3144 99.5127
R3476 VDD.n3150 VDD.n3129 99.5127
R3477 VDD.n3154 VDD.n3152 99.5127
R3478 VDD.n3158 VDD.n3127 99.5127
R3479 VDD.n3162 VDD.n3160 99.5127
R3480 VDD.n3167 VDD.n3123 99.5127
R3481 VDD.n3170 VDD.n3169 99.5127
R3482 VDD.n3658 VDD.n3657 99.5127
R3483 VDD.n3655 VDD.n3641 99.5127
R3484 VDD.n3651 VDD.n3650 99.5127
R3485 VDD.n3648 VDD.n3645 99.5127
R3486 VDD.n3736 VDD.n472 99.5127
R3487 VDD.n3734 VDD.n3733 99.5127
R3488 VDD.n3731 VDD.n475 99.5127
R3489 VDD.n3727 VDD.n3726 99.5127
R3490 VDD.n3724 VDD.n478 99.5127
R3491 VDD.n3249 VDD.n2978 99.5127
R3492 VDD.n3249 VDD.n900 99.5127
R3493 VDD.n3246 VDD.n900 99.5127
R3494 VDD.n3246 VDD.n894 99.5127
R3495 VDD.n3243 VDD.n894 99.5127
R3496 VDD.n3243 VDD.n888 99.5127
R3497 VDD.n3240 VDD.n888 99.5127
R3498 VDD.n3240 VDD.n882 99.5127
R3499 VDD.n3119 VDD.n882 99.5127
R3500 VDD.n3119 VDD.n877 99.5127
R3501 VDD.n3116 VDD.n877 99.5127
R3502 VDD.n3116 VDD.n871 99.5127
R3503 VDD.n3113 VDD.n871 99.5127
R3504 VDD.n3113 VDD.n865 99.5127
R3505 VDD.n3110 VDD.n865 99.5127
R3506 VDD.n3110 VDD.n859 99.5127
R3507 VDD.n3107 VDD.n859 99.5127
R3508 VDD.n3107 VDD.n853 99.5127
R3509 VDD.n3104 VDD.n853 99.5127
R3510 VDD.n3104 VDD.n847 99.5127
R3511 VDD.n3101 VDD.n847 99.5127
R3512 VDD.n3101 VDD.n840 99.5127
R3513 VDD.n3098 VDD.n840 99.5127
R3514 VDD.n3098 VDD.n834 99.5127
R3515 VDD.n3095 VDD.n834 99.5127
R3516 VDD.n3095 VDD.n829 99.5127
R3517 VDD.n3092 VDD.n829 99.5127
R3518 VDD.n3092 VDD.n823 99.5127
R3519 VDD.n3089 VDD.n823 99.5127
R3520 VDD.n3089 VDD.n816 99.5127
R3521 VDD.n3086 VDD.n816 99.5127
R3522 VDD.n3086 VDD.n810 99.5127
R3523 VDD.n3083 VDD.n810 99.5127
R3524 VDD.n3083 VDD.n804 99.5127
R3525 VDD.n3080 VDD.n804 99.5127
R3526 VDD.n3080 VDD.n798 99.5127
R3527 VDD.n3077 VDD.n798 99.5127
R3528 VDD.n3077 VDD.n793 99.5127
R3529 VDD.n3074 VDD.n793 99.5127
R3530 VDD.n3074 VDD.n787 99.5127
R3531 VDD.n3071 VDD.n787 99.5127
R3532 VDD.n3071 VDD.n780 99.5127
R3533 VDD.n3068 VDD.n780 99.5127
R3534 VDD.n3068 VDD.n773 99.5127
R3535 VDD.n3065 VDD.n773 99.5127
R3536 VDD.n3065 VDD.n767 99.5127
R3537 VDD.n3062 VDD.n767 99.5127
R3538 VDD.n3062 VDD.n761 99.5127
R3539 VDD.n3059 VDD.n761 99.5127
R3540 VDD.n3059 VDD.n755 99.5127
R3541 VDD.n3056 VDD.n755 99.5127
R3542 VDD.n3056 VDD.n749 99.5127
R3543 VDD.n3053 VDD.n749 99.5127
R3544 VDD.n3053 VDD.n743 99.5127
R3545 VDD.n3050 VDD.n743 99.5127
R3546 VDD.n3050 VDD.n737 99.5127
R3547 VDD.n3047 VDD.n737 99.5127
R3548 VDD.n3047 VDD.n731 99.5127
R3549 VDD.n3044 VDD.n731 99.5127
R3550 VDD.n3044 VDD.n725 99.5127
R3551 VDD.n3041 VDD.n725 99.5127
R3552 VDD.n3041 VDD.n719 99.5127
R3553 VDD.n3038 VDD.n719 99.5127
R3554 VDD.n3038 VDD.n713 99.5127
R3555 VDD.n3035 VDD.n713 99.5127
R3556 VDD.n3035 VDD.n707 99.5127
R3557 VDD.n3032 VDD.n707 99.5127
R3558 VDD.n3032 VDD.n701 99.5127
R3559 VDD.n3029 VDD.n701 99.5127
R3560 VDD.n3029 VDD.n695 99.5127
R3561 VDD.n3026 VDD.n695 99.5127
R3562 VDD.n3026 VDD.n689 99.5127
R3563 VDD.n3023 VDD.n689 99.5127
R3564 VDD.n3023 VDD.n683 99.5127
R3565 VDD.n3020 VDD.n683 99.5127
R3566 VDD.n3020 VDD.n677 99.5127
R3567 VDD.n3017 VDD.n677 99.5127
R3568 VDD.n3017 VDD.n671 99.5127
R3569 VDD.n3014 VDD.n671 99.5127
R3570 VDD.n3014 VDD.n665 99.5127
R3571 VDD.n3011 VDD.n665 99.5127
R3572 VDD.n3011 VDD.n659 99.5127
R3573 VDD.n3008 VDD.n659 99.5127
R3574 VDD.n3008 VDD.n653 99.5127
R3575 VDD.n3005 VDD.n653 99.5127
R3576 VDD.n3005 VDD.n646 99.5127
R3577 VDD.n3002 VDD.n646 99.5127
R3578 VDD.n3002 VDD.n640 99.5127
R3579 VDD.n2999 VDD.n640 99.5127
R3580 VDD.n2999 VDD.n635 99.5127
R3581 VDD.n2996 VDD.n635 99.5127
R3582 VDD.n2996 VDD.n628 99.5127
R3583 VDD.n2993 VDD.n628 99.5127
R3584 VDD.n2993 VDD.n621 99.5127
R3585 VDD.n621 VDD.n484 99.5127
R3586 VDD.n3719 VDD.n484 99.5127
R3587 VDD.n3290 VDD.n3288 99.5127
R3588 VDD.n3286 VDD.n2981 99.5127
R3589 VDD.n3282 VDD.n3280 99.5127
R3590 VDD.n3278 VDD.n2983 99.5127
R3591 VDD.n3274 VDD.n3272 99.5127
R3592 VDD.n3270 VDD.n2985 99.5127
R3593 VDD.n3266 VDD.n3264 99.5127
R3594 VDD.n3262 VDD.n2987 99.5127
R3595 VDD.n3257 VDD.n3255 99.5127
R3596 VDD.n3294 VDD.n897 99.5127
R3597 VDD.n3302 VDD.n897 99.5127
R3598 VDD.n3302 VDD.n895 99.5127
R3599 VDD.n3306 VDD.n895 99.5127
R3600 VDD.n3306 VDD.n885 99.5127
R3601 VDD.n3314 VDD.n885 99.5127
R3602 VDD.n3314 VDD.n883 99.5127
R3603 VDD.n3318 VDD.n883 99.5127
R3604 VDD.n3318 VDD.n874 99.5127
R3605 VDD.n3326 VDD.n874 99.5127
R3606 VDD.n3326 VDD.n872 99.5127
R3607 VDD.n3330 VDD.n872 99.5127
R3608 VDD.n3330 VDD.n862 99.5127
R3609 VDD.n3338 VDD.n862 99.5127
R3610 VDD.n3338 VDD.n860 99.5127
R3611 VDD.n3342 VDD.n860 99.5127
R3612 VDD.n3342 VDD.n850 99.5127
R3613 VDD.n3350 VDD.n850 99.5127
R3614 VDD.n3350 VDD.n848 99.5127
R3615 VDD.n3354 VDD.n848 99.5127
R3616 VDD.n3354 VDD.n837 99.5127
R3617 VDD.n3362 VDD.n837 99.5127
R3618 VDD.n3362 VDD.n835 99.5127
R3619 VDD.n3366 VDD.n835 99.5127
R3620 VDD.n3366 VDD.n826 99.5127
R3621 VDD.n3374 VDD.n826 99.5127
R3622 VDD.n3374 VDD.n824 99.5127
R3623 VDD.n3378 VDD.n824 99.5127
R3624 VDD.n3378 VDD.n813 99.5127
R3625 VDD.n3386 VDD.n813 99.5127
R3626 VDD.n3386 VDD.n811 99.5127
R3627 VDD.n3390 VDD.n811 99.5127
R3628 VDD.n3390 VDD.n801 99.5127
R3629 VDD.n3398 VDD.n801 99.5127
R3630 VDD.n3398 VDD.n799 99.5127
R3631 VDD.n3402 VDD.n799 99.5127
R3632 VDD.n3402 VDD.n790 99.5127
R3633 VDD.n3410 VDD.n790 99.5127
R3634 VDD.n3410 VDD.n788 99.5127
R3635 VDD.n3414 VDD.n788 99.5127
R3636 VDD.n3414 VDD.n777 99.5127
R3637 VDD.n3422 VDD.n777 99.5127
R3638 VDD.n3422 VDD.n774 99.5127
R3639 VDD.n3431 VDD.n774 99.5127
R3640 VDD.n3431 VDD.n775 99.5127
R3641 VDD.n775 VDD.n768 99.5127
R3642 VDD.n3426 VDD.n768 99.5127
R3643 VDD.n3426 VDD.n760 99.5127
R3644 VDD.n760 VDD.n752 99.5127
R3645 VDD.n3516 VDD.n752 99.5127
R3646 VDD.n3516 VDD.n750 99.5127
R3647 VDD.n3520 VDD.n750 99.5127
R3648 VDD.n3520 VDD.n740 99.5127
R3649 VDD.n3528 VDD.n740 99.5127
R3650 VDD.n3528 VDD.n738 99.5127
R3651 VDD.n3532 VDD.n738 99.5127
R3652 VDD.n3532 VDD.n728 99.5127
R3653 VDD.n3540 VDD.n728 99.5127
R3654 VDD.n3540 VDD.n726 99.5127
R3655 VDD.n3544 VDD.n726 99.5127
R3656 VDD.n3544 VDD.n716 99.5127
R3657 VDD.n3552 VDD.n716 99.5127
R3658 VDD.n3552 VDD.n714 99.5127
R3659 VDD.n3556 VDD.n714 99.5127
R3660 VDD.n3556 VDD.n704 99.5127
R3661 VDD.n3564 VDD.n704 99.5127
R3662 VDD.n3564 VDD.n702 99.5127
R3663 VDD.n3568 VDD.n702 99.5127
R3664 VDD.n3568 VDD.n692 99.5127
R3665 VDD.n3576 VDD.n692 99.5127
R3666 VDD.n3576 VDD.n690 99.5127
R3667 VDD.n3580 VDD.n690 99.5127
R3668 VDD.n3580 VDD.n680 99.5127
R3669 VDD.n3588 VDD.n680 99.5127
R3670 VDD.n3588 VDD.n678 99.5127
R3671 VDD.n3592 VDD.n678 99.5127
R3672 VDD.n3592 VDD.n668 99.5127
R3673 VDD.n3600 VDD.n668 99.5127
R3674 VDD.n3600 VDD.n666 99.5127
R3675 VDD.n3604 VDD.n666 99.5127
R3676 VDD.n3604 VDD.n656 99.5127
R3677 VDD.n3612 VDD.n656 99.5127
R3678 VDD.n3612 VDD.n654 99.5127
R3679 VDD.n3616 VDD.n654 99.5127
R3680 VDD.n3616 VDD.n643 99.5127
R3681 VDD.n3624 VDD.n643 99.5127
R3682 VDD.n3624 VDD.n641 99.5127
R3683 VDD.n3628 VDD.n641 99.5127
R3684 VDD.n3628 VDD.n632 99.5127
R3685 VDD.n3636 VDD.n632 99.5127
R3686 VDD.n3636 VDD.n629 99.5127
R3687 VDD.n3668 VDD.n629 99.5127
R3688 VDD.n3668 VDD.n630 99.5127
R3689 VDD.n630 VDD.n622 99.5127
R3690 VDD.n3663 VDD.n622 99.5127
R3691 VDD.n3663 VDD.n487 99.5127
R3692 VDD.n2898 VDD.n2897 99.5127
R3693 VDD.n2894 VDD.n2893 99.5127
R3694 VDD.n2890 VDD.n2889 99.5127
R3695 VDD.n2886 VDD.n2885 99.5127
R3696 VDD.n2882 VDD.n2881 99.5127
R3697 VDD.n2878 VDD.n2877 99.5127
R3698 VDD.n2874 VDD.n2873 99.5127
R3699 VDD.n2870 VDD.n2869 99.5127
R3700 VDD.n2865 VDD.n924 99.5127
R3701 VDD.n2482 VDD.n1216 99.5127
R3702 VDD.n2478 VDD.n1216 99.5127
R3703 VDD.n2478 VDD.n1210 99.5127
R3704 VDD.n2475 VDD.n1210 99.5127
R3705 VDD.n2475 VDD.n1204 99.5127
R3706 VDD.n2472 VDD.n1204 99.5127
R3707 VDD.n2472 VDD.n1198 99.5127
R3708 VDD.n2469 VDD.n1198 99.5127
R3709 VDD.n2469 VDD.n1192 99.5127
R3710 VDD.n2305 VDD.n1192 99.5127
R3711 VDD.n2305 VDD.n1187 99.5127
R3712 VDD.n2302 VDD.n1187 99.5127
R3713 VDD.n2302 VDD.n1181 99.5127
R3714 VDD.n2299 VDD.n1181 99.5127
R3715 VDD.n2299 VDD.n1175 99.5127
R3716 VDD.n2296 VDD.n1175 99.5127
R3717 VDD.n2296 VDD.n1169 99.5127
R3718 VDD.n2293 VDD.n1169 99.5127
R3719 VDD.n2293 VDD.n1163 99.5127
R3720 VDD.n2290 VDD.n1163 99.5127
R3721 VDD.n2290 VDD.n1157 99.5127
R3722 VDD.n2287 VDD.n1157 99.5127
R3723 VDD.n2287 VDD.n1151 99.5127
R3724 VDD.n2284 VDD.n1151 99.5127
R3725 VDD.n2284 VDD.n1145 99.5127
R3726 VDD.n2281 VDD.n1145 99.5127
R3727 VDD.n2281 VDD.n1139 99.5127
R3728 VDD.n2278 VDD.n1139 99.5127
R3729 VDD.n2278 VDD.n1133 99.5127
R3730 VDD.n2275 VDD.n1133 99.5127
R3731 VDD.n2275 VDD.n1127 99.5127
R3732 VDD.n2272 VDD.n1127 99.5127
R3733 VDD.n2272 VDD.n1121 99.5127
R3734 VDD.n2269 VDD.n1121 99.5127
R3735 VDD.n2269 VDD.n1115 99.5127
R3736 VDD.n2266 VDD.n1115 99.5127
R3737 VDD.n2266 VDD.n1109 99.5127
R3738 VDD.n2263 VDD.n1109 99.5127
R3739 VDD.n2263 VDD.n1103 99.5127
R3740 VDD.n2260 VDD.n1103 99.5127
R3741 VDD.n2260 VDD.n1097 99.5127
R3742 VDD.n2257 VDD.n1097 99.5127
R3743 VDD.n2257 VDD.n1091 99.5127
R3744 VDD.n2254 VDD.n1091 99.5127
R3745 VDD.n2254 VDD.n1085 99.5127
R3746 VDD.n2251 VDD.n1085 99.5127
R3747 VDD.n2251 VDD.n1079 99.5127
R3748 VDD.n2248 VDD.n1079 99.5127
R3749 VDD.n2248 VDD.n1073 99.5127
R3750 VDD.n2245 VDD.n1073 99.5127
R3751 VDD.n2245 VDD.n1067 99.5127
R3752 VDD.n2242 VDD.n1067 99.5127
R3753 VDD.n2242 VDD.n1061 99.5127
R3754 VDD.n2239 VDD.n1061 99.5127
R3755 VDD.n2239 VDD.n1056 99.5127
R3756 VDD.n2236 VDD.n1056 99.5127
R3757 VDD.n2236 VDD.n1050 99.5127
R3758 VDD.n2233 VDD.n1050 99.5127
R3759 VDD.n2233 VDD.n1043 99.5127
R3760 VDD.n2230 VDD.n1043 99.5127
R3761 VDD.n2230 VDD.n1037 99.5127
R3762 VDD.n2227 VDD.n1037 99.5127
R3763 VDD.n2227 VDD.n1031 99.5127
R3764 VDD.n2224 VDD.n1031 99.5127
R3765 VDD.n2224 VDD.n1025 99.5127
R3766 VDD.n2221 VDD.n1025 99.5127
R3767 VDD.n2221 VDD.n1020 99.5127
R3768 VDD.n2218 VDD.n1020 99.5127
R3769 VDD.n2218 VDD.n1014 99.5127
R3770 VDD.n2215 VDD.n1014 99.5127
R3771 VDD.n2215 VDD.n1007 99.5127
R3772 VDD.n2212 VDD.n1007 99.5127
R3773 VDD.n2212 VDD.n1001 99.5127
R3774 VDD.n2209 VDD.n1001 99.5127
R3775 VDD.n2209 VDD.n996 99.5127
R3776 VDD.n2206 VDD.n996 99.5127
R3777 VDD.n2206 VDD.n990 99.5127
R3778 VDD.n2203 VDD.n990 99.5127
R3779 VDD.n2203 VDD.n984 99.5127
R3780 VDD.n2200 VDD.n984 99.5127
R3781 VDD.n2200 VDD.n978 99.5127
R3782 VDD.n2197 VDD.n978 99.5127
R3783 VDD.n2197 VDD.n972 99.5127
R3784 VDD.n2194 VDD.n972 99.5127
R3785 VDD.n2194 VDD.n966 99.5127
R3786 VDD.n2191 VDD.n966 99.5127
R3787 VDD.n2191 VDD.n959 99.5127
R3788 VDD.n2188 VDD.n959 99.5127
R3789 VDD.n2188 VDD.n953 99.5127
R3790 VDD.n2185 VDD.n953 99.5127
R3791 VDD.n2185 VDD.n947 99.5127
R3792 VDD.n2182 VDD.n947 99.5127
R3793 VDD.n2182 VDD.n940 99.5127
R3794 VDD.n940 VDD.n928 99.5127
R3795 VDD.n2969 VDD.n928 99.5127
R3796 VDD.n2969 VDD.n925 99.5127
R3797 VDD.n2164 VDD.n2163 99.5127
R3798 VDD.n2168 VDD.n2167 99.5127
R3799 VDD.n2172 VDD.n2171 99.5127
R3800 VDD.n2176 VDD.n2175 99.5127
R3801 VDD.n2503 VDD.n2502 99.5127
R3802 VDD.n2500 VDD.n2499 99.5127
R3803 VDD.n2496 VDD.n2495 99.5127
R3804 VDD.n2492 VDD.n2491 99.5127
R3805 VDD.n2487 VDD.n2486 99.5127
R3806 VDD.n2596 VDD.n1213 99.5127
R3807 VDD.n2596 VDD.n1211 99.5127
R3808 VDD.n2600 VDD.n1211 99.5127
R3809 VDD.n2600 VDD.n1201 99.5127
R3810 VDD.n2608 VDD.n1201 99.5127
R3811 VDD.n2608 VDD.n1199 99.5127
R3812 VDD.n2612 VDD.n1199 99.5127
R3813 VDD.n2612 VDD.n1190 99.5127
R3814 VDD.n2620 VDD.n1190 99.5127
R3815 VDD.n2620 VDD.n1188 99.5127
R3816 VDD.n2624 VDD.n1188 99.5127
R3817 VDD.n2624 VDD.n1178 99.5127
R3818 VDD.n2632 VDD.n1178 99.5127
R3819 VDD.n2632 VDD.n1176 99.5127
R3820 VDD.n2636 VDD.n1176 99.5127
R3821 VDD.n2636 VDD.n1166 99.5127
R3822 VDD.n2644 VDD.n1166 99.5127
R3823 VDD.n2644 VDD.n1164 99.5127
R3824 VDD.n2648 VDD.n1164 99.5127
R3825 VDD.n2648 VDD.n1154 99.5127
R3826 VDD.n2656 VDD.n1154 99.5127
R3827 VDD.n2656 VDD.n1152 99.5127
R3828 VDD.n2660 VDD.n1152 99.5127
R3829 VDD.n2660 VDD.n1142 99.5127
R3830 VDD.n2668 VDD.n1142 99.5127
R3831 VDD.n2668 VDD.n1140 99.5127
R3832 VDD.n2672 VDD.n1140 99.5127
R3833 VDD.n2672 VDD.n1130 99.5127
R3834 VDD.n2680 VDD.n1130 99.5127
R3835 VDD.n2680 VDD.n1128 99.5127
R3836 VDD.n2684 VDD.n1128 99.5127
R3837 VDD.n2684 VDD.n1118 99.5127
R3838 VDD.n2692 VDD.n1118 99.5127
R3839 VDD.n2692 VDD.n1116 99.5127
R3840 VDD.n2696 VDD.n1116 99.5127
R3841 VDD.n2696 VDD.n1106 99.5127
R3842 VDD.n2704 VDD.n1106 99.5127
R3843 VDD.n2704 VDD.n1104 99.5127
R3844 VDD.n2708 VDD.n1104 99.5127
R3845 VDD.n2708 VDD.n1094 99.5127
R3846 VDD.n2716 VDD.n1094 99.5127
R3847 VDD.n2716 VDD.n1092 99.5127
R3848 VDD.n2720 VDD.n1092 99.5127
R3849 VDD.n2720 VDD.n1082 99.5127
R3850 VDD.n2728 VDD.n1082 99.5127
R3851 VDD.n2728 VDD.n1080 99.5127
R3852 VDD.n2732 VDD.n1080 99.5127
R3853 VDD.n2732 VDD.n1071 99.5127
R3854 VDD.n2740 VDD.n1071 99.5127
R3855 VDD.n2740 VDD.n1069 99.5127
R3856 VDD.n2744 VDD.n1069 99.5127
R3857 VDD.n2744 VDD.n1059 99.5127
R3858 VDD.n2752 VDD.n1059 99.5127
R3859 VDD.n2752 VDD.n1057 99.5127
R3860 VDD.n2756 VDD.n1057 99.5127
R3861 VDD.n2756 VDD.n1047 99.5127
R3862 VDD.n2764 VDD.n1047 99.5127
R3863 VDD.n2764 VDD.n1045 99.5127
R3864 VDD.n2768 VDD.n1045 99.5127
R3865 VDD.n2768 VDD.n1035 99.5127
R3866 VDD.n2776 VDD.n1035 99.5127
R3867 VDD.n2776 VDD.n1033 99.5127
R3868 VDD.n2780 VDD.n1033 99.5127
R3869 VDD.n2780 VDD.n1023 99.5127
R3870 VDD.n2788 VDD.n1023 99.5127
R3871 VDD.n2788 VDD.n1021 99.5127
R3872 VDD.n2792 VDD.n1021 99.5127
R3873 VDD.n2792 VDD.n1011 99.5127
R3874 VDD.n2800 VDD.n1011 99.5127
R3875 VDD.n2800 VDD.n1009 99.5127
R3876 VDD.n2804 VDD.n1009 99.5127
R3877 VDD.n2804 VDD.n999 99.5127
R3878 VDD.n2812 VDD.n999 99.5127
R3879 VDD.n2812 VDD.n997 99.5127
R3880 VDD.n2816 VDD.n997 99.5127
R3881 VDD.n2816 VDD.n987 99.5127
R3882 VDD.n2824 VDD.n987 99.5127
R3883 VDD.n2824 VDD.n985 99.5127
R3884 VDD.n2828 VDD.n985 99.5127
R3885 VDD.n2828 VDD.n975 99.5127
R3886 VDD.n2836 VDD.n975 99.5127
R3887 VDD.n2836 VDD.n973 99.5127
R3888 VDD.n2840 VDD.n973 99.5127
R3889 VDD.n2840 VDD.n963 99.5127
R3890 VDD.n2848 VDD.n963 99.5127
R3891 VDD.n2848 VDD.n961 99.5127
R3892 VDD.n2852 VDD.n961 99.5127
R3893 VDD.n2852 VDD.n951 99.5127
R3894 VDD.n2860 VDD.n951 99.5127
R3895 VDD.n2860 VDD.n948 99.5127
R3896 VDD.n2910 VDD.n948 99.5127
R3897 VDD.n2910 VDD.n949 99.5127
R3898 VDD.n949 VDD.n941 99.5127
R3899 VDD.n2905 VDD.n941 99.5127
R3900 VDD.n2905 VDD.n931 99.5127
R3901 VDD.n2902 VDD.n931 99.5127
R3902 VDD.n2961 VDD.n2960 99.5127
R3903 VDD.n2957 VDD.n2956 99.5127
R3904 VDD.n2953 VDD.n2952 99.5127
R3905 VDD.n2949 VDD.n2948 99.5127
R3906 VDD.n2945 VDD.n2944 99.5127
R3907 VDD.n2941 VDD.n2940 99.5127
R3908 VDD.n2937 VDD.n2936 99.5127
R3909 VDD.n2933 VDD.n2932 99.5127
R3910 VDD.n2928 VDD.n2927 99.5127
R3911 VDD.n2329 VDD.n1215 99.5127
R3912 VDD.n2332 VDD.n1215 99.5127
R3913 VDD.n2332 VDD.n1209 99.5127
R3914 VDD.n2335 VDD.n1209 99.5127
R3915 VDD.n2335 VDD.n1203 99.5127
R3916 VDD.n2338 VDD.n1203 99.5127
R3917 VDD.n2338 VDD.n1197 99.5127
R3918 VDD.n2467 VDD.n1197 99.5127
R3919 VDD.n2467 VDD.n1191 99.5127
R3920 VDD.n2463 VDD.n1191 99.5127
R3921 VDD.n2463 VDD.n1186 99.5127
R3922 VDD.n2460 VDD.n1186 99.5127
R3923 VDD.n2460 VDD.n1180 99.5127
R3924 VDD.n2457 VDD.n1180 99.5127
R3925 VDD.n2457 VDD.n1174 99.5127
R3926 VDD.n2454 VDD.n1174 99.5127
R3927 VDD.n2454 VDD.n1168 99.5127
R3928 VDD.n2451 VDD.n1168 99.5127
R3929 VDD.n2451 VDD.n1162 99.5127
R3930 VDD.n2448 VDD.n1162 99.5127
R3931 VDD.n2448 VDD.n1156 99.5127
R3932 VDD.n2445 VDD.n1156 99.5127
R3933 VDD.n2445 VDD.n1150 99.5127
R3934 VDD.n2442 VDD.n1150 99.5127
R3935 VDD.n2442 VDD.n1144 99.5127
R3936 VDD.n2439 VDD.n1144 99.5127
R3937 VDD.n2439 VDD.n1138 99.5127
R3938 VDD.n2436 VDD.n1138 99.5127
R3939 VDD.n2436 VDD.n1132 99.5127
R3940 VDD.n2433 VDD.n1132 99.5127
R3941 VDD.n2433 VDD.n1126 99.5127
R3942 VDD.n2430 VDD.n1126 99.5127
R3943 VDD.n2430 VDD.n1120 99.5127
R3944 VDD.n2427 VDD.n1120 99.5127
R3945 VDD.n2427 VDD.n1114 99.5127
R3946 VDD.n2424 VDD.n1114 99.5127
R3947 VDD.n2424 VDD.n1108 99.5127
R3948 VDD.n2421 VDD.n1108 99.5127
R3949 VDD.n2421 VDD.n1102 99.5127
R3950 VDD.n2418 VDD.n1102 99.5127
R3951 VDD.n2418 VDD.n1096 99.5127
R3952 VDD.n2415 VDD.n1096 99.5127
R3953 VDD.n2415 VDD.n1090 99.5127
R3954 VDD.n2412 VDD.n1090 99.5127
R3955 VDD.n2412 VDD.n1084 99.5127
R3956 VDD.n2409 VDD.n1084 99.5127
R3957 VDD.n2409 VDD.n1078 99.5127
R3958 VDD.n2406 VDD.n1078 99.5127
R3959 VDD.n2406 VDD.n1072 99.5127
R3960 VDD.n2403 VDD.n1072 99.5127
R3961 VDD.n2403 VDD.n1066 99.5127
R3962 VDD.n2400 VDD.n1066 99.5127
R3963 VDD.n2400 VDD.n1060 99.5127
R3964 VDD.n2397 VDD.n1060 99.5127
R3965 VDD.n2397 VDD.n1055 99.5127
R3966 VDD.n2394 VDD.n1055 99.5127
R3967 VDD.n2394 VDD.n1049 99.5127
R3968 VDD.n2391 VDD.n1049 99.5127
R3969 VDD.n2391 VDD.n1042 99.5127
R3970 VDD.n2388 VDD.n1042 99.5127
R3971 VDD.n2388 VDD.n1036 99.5127
R3972 VDD.n2385 VDD.n1036 99.5127
R3973 VDD.n2385 VDD.n1030 99.5127
R3974 VDD.n2382 VDD.n1030 99.5127
R3975 VDD.n2382 VDD.n1024 99.5127
R3976 VDD.n2379 VDD.n1024 99.5127
R3977 VDD.n2379 VDD.n1019 99.5127
R3978 VDD.n2376 VDD.n1019 99.5127
R3979 VDD.n2376 VDD.n1013 99.5127
R3980 VDD.n2373 VDD.n1013 99.5127
R3981 VDD.n2373 VDD.n1006 99.5127
R3982 VDD.n2370 VDD.n1006 99.5127
R3983 VDD.n2370 VDD.n1000 99.5127
R3984 VDD.n2367 VDD.n1000 99.5127
R3985 VDD.n2367 VDD.n995 99.5127
R3986 VDD.n2364 VDD.n995 99.5127
R3987 VDD.n2364 VDD.n989 99.5127
R3988 VDD.n2361 VDD.n989 99.5127
R3989 VDD.n2361 VDD.n983 99.5127
R3990 VDD.n2358 VDD.n983 99.5127
R3991 VDD.n2358 VDD.n977 99.5127
R3992 VDD.n2355 VDD.n977 99.5127
R3993 VDD.n2355 VDD.n971 99.5127
R3994 VDD.n2352 VDD.n971 99.5127
R3995 VDD.n2352 VDD.n965 99.5127
R3996 VDD.n2349 VDD.n965 99.5127
R3997 VDD.n2349 VDD.n958 99.5127
R3998 VDD.n2346 VDD.n958 99.5127
R3999 VDD.n2346 VDD.n952 99.5127
R4000 VDD.n2343 VDD.n952 99.5127
R4001 VDD.n2343 VDD.n946 99.5127
R4002 VDD.n946 VDD.n938 99.5127
R4003 VDD.n2918 VDD.n938 99.5127
R4004 VDD.n2919 VDD.n2918 99.5127
R4005 VDD.n2919 VDD.n930 99.5127
R4006 VDD.n2923 VDD.n930 99.5127
R4007 VDD.n2587 VDD.n1219 99.5127
R4008 VDD.n2587 VDD.n1239 99.5127
R4009 VDD.n2583 VDD.n2582 99.5127
R4010 VDD.n2579 VDD.n2578 99.5127
R4011 VDD.n2575 VDD.n2574 99.5127
R4012 VDD.n2312 VDD.n2311 99.5127
R4013 VDD.n2316 VDD.n2315 99.5127
R4014 VDD.n2320 VDD.n2319 99.5127
R4015 VDD.n2324 VDD.n2323 99.5127
R4016 VDD.n2326 VDD.n1228 99.5127
R4017 VDD.n2594 VDD.n1217 99.5127
R4018 VDD.n2594 VDD.n1207 99.5127
R4019 VDD.n2602 VDD.n1207 99.5127
R4020 VDD.n2602 VDD.n1205 99.5127
R4021 VDD.n2606 VDD.n1205 99.5127
R4022 VDD.n2606 VDD.n1195 99.5127
R4023 VDD.n2614 VDD.n1195 99.5127
R4024 VDD.n2614 VDD.n1193 99.5127
R4025 VDD.n2618 VDD.n1193 99.5127
R4026 VDD.n2618 VDD.n1184 99.5127
R4027 VDD.n2626 VDD.n1184 99.5127
R4028 VDD.n2626 VDD.n1182 99.5127
R4029 VDD.n2630 VDD.n1182 99.5127
R4030 VDD.n2630 VDD.n1172 99.5127
R4031 VDD.n2638 VDD.n1172 99.5127
R4032 VDD.n2638 VDD.n1170 99.5127
R4033 VDD.n2642 VDD.n1170 99.5127
R4034 VDD.n2642 VDD.n1160 99.5127
R4035 VDD.n2650 VDD.n1160 99.5127
R4036 VDD.n2650 VDD.n1158 99.5127
R4037 VDD.n2654 VDD.n1158 99.5127
R4038 VDD.n2654 VDD.n1148 99.5127
R4039 VDD.n2662 VDD.n1148 99.5127
R4040 VDD.n2662 VDD.n1146 99.5127
R4041 VDD.n2666 VDD.n1146 99.5127
R4042 VDD.n2666 VDD.n1136 99.5127
R4043 VDD.n2674 VDD.n1136 99.5127
R4044 VDD.n2674 VDD.n1134 99.5127
R4045 VDD.n2678 VDD.n1134 99.5127
R4046 VDD.n2678 VDD.n1124 99.5127
R4047 VDD.n2686 VDD.n1124 99.5127
R4048 VDD.n2686 VDD.n1122 99.5127
R4049 VDD.n2690 VDD.n1122 99.5127
R4050 VDD.n2690 VDD.n1112 99.5127
R4051 VDD.n2698 VDD.n1112 99.5127
R4052 VDD.n2698 VDD.n1110 99.5127
R4053 VDD.n2702 VDD.n1110 99.5127
R4054 VDD.n2702 VDD.n1100 99.5127
R4055 VDD.n2710 VDD.n1100 99.5127
R4056 VDD.n2710 VDD.n1098 99.5127
R4057 VDD.n2714 VDD.n1098 99.5127
R4058 VDD.n2714 VDD.n1088 99.5127
R4059 VDD.n2722 VDD.n1088 99.5127
R4060 VDD.n2722 VDD.n1086 99.5127
R4061 VDD.n2726 VDD.n1086 99.5127
R4062 VDD.n2726 VDD.n1076 99.5127
R4063 VDD.n2734 VDD.n1076 99.5127
R4064 VDD.n2734 VDD.n1074 99.5127
R4065 VDD.n2738 VDD.n1074 99.5127
R4066 VDD.n2738 VDD.n1064 99.5127
R4067 VDD.n2746 VDD.n1064 99.5127
R4068 VDD.n2746 VDD.n1062 99.5127
R4069 VDD.n2750 VDD.n1062 99.5127
R4070 VDD.n2750 VDD.n1053 99.5127
R4071 VDD.n2758 VDD.n1053 99.5127
R4072 VDD.n2758 VDD.n1051 99.5127
R4073 VDD.n2762 VDD.n1051 99.5127
R4074 VDD.n2762 VDD.n1040 99.5127
R4075 VDD.n2770 VDD.n1040 99.5127
R4076 VDD.n2770 VDD.n1038 99.5127
R4077 VDD.n2774 VDD.n1038 99.5127
R4078 VDD.n2774 VDD.n1028 99.5127
R4079 VDD.n2782 VDD.n1028 99.5127
R4080 VDD.n2782 VDD.n1026 99.5127
R4081 VDD.n2786 VDD.n1026 99.5127
R4082 VDD.n2786 VDD.n1017 99.5127
R4083 VDD.n2794 VDD.n1017 99.5127
R4084 VDD.n2794 VDD.n1015 99.5127
R4085 VDD.n2798 VDD.n1015 99.5127
R4086 VDD.n2798 VDD.n1004 99.5127
R4087 VDD.n2806 VDD.n1004 99.5127
R4088 VDD.n2806 VDD.n1002 99.5127
R4089 VDD.n2810 VDD.n1002 99.5127
R4090 VDD.n2810 VDD.n993 99.5127
R4091 VDD.n2818 VDD.n993 99.5127
R4092 VDD.n2818 VDD.n991 99.5127
R4093 VDD.n2822 VDD.n991 99.5127
R4094 VDD.n2822 VDD.n981 99.5127
R4095 VDD.n2830 VDD.n981 99.5127
R4096 VDD.n2830 VDD.n979 99.5127
R4097 VDD.n2834 VDD.n979 99.5127
R4098 VDD.n2834 VDD.n969 99.5127
R4099 VDD.n2842 VDD.n969 99.5127
R4100 VDD.n2842 VDD.n967 99.5127
R4101 VDD.n2846 VDD.n967 99.5127
R4102 VDD.n2846 VDD.n956 99.5127
R4103 VDD.n2854 VDD.n956 99.5127
R4104 VDD.n2854 VDD.n954 99.5127
R4105 VDD.n2858 VDD.n954 99.5127
R4106 VDD.n2858 VDD.n944 99.5127
R4107 VDD.n2912 VDD.n944 99.5127
R4108 VDD.n2912 VDD.n942 99.5127
R4109 VDD.n2916 VDD.n942 99.5127
R4110 VDD.n2916 VDD.n932 99.5127
R4111 VDD.n2967 VDD.n932 99.5127
R4112 VDD.n2967 VDD.n933 99.5127
R4113 VDD.n1950 VDD.t129 98.4153
R4114 VDD.n1944 VDD.t70 98.4153
R4115 VDD.n27 VDD.t8 95.9929
R4116 VDD.n21 VDD.t46 95.9929
R4117 VDD.n24 VDD.n22 91.8087
R4118 VDD.n18 VDD.n16 91.8087
R4119 VDD.n26 VDD.n25 89.3863
R4120 VDD.n24 VDD.n23 89.3863
R4121 VDD.n20 VDD.n19 89.3863
R4122 VDD.n18 VDD.n17 89.3863
R4123 VDD.n1950 VDD.n1949 89.3863
R4124 VDD.n1952 VDD.n1951 89.3863
R4125 VDD.n1954 VDD.n1953 89.3863
R4126 VDD.n1944 VDD.n1943 89.3863
R4127 VDD.n1946 VDD.n1945 89.3863
R4128 VDD.n1948 VDD.n1947 89.3863
R4129 VDD.n2309 VDD.n2308 82.0369
R4130 VDD.n936 VDD.n935 82.0369
R4131 VDD.n2989 VDD.n2988 82.0369
R4132 VDD.n615 VDD.n614 82.0369
R4133 VDD.n3125 VDD.n3124 82.0369
R4134 VDD.n480 VDD.n479 82.0369
R4135 VDD.n2180 VDD.n2179 82.0369
R4136 VDD.n2864 VDD.n2863 82.0369
R4137 VDD.n2588 VDD.n1238 72.8958
R4138 VDD.n2588 VDD.n1237 72.8958
R4139 VDD.n2588 VDD.n1236 72.8958
R4140 VDD.n2588 VDD.n1235 72.8958
R4141 VDD.n2588 VDD.n1234 72.8958
R4142 VDD.n2588 VDD.n1233 72.8958
R4143 VDD.n2588 VDD.n1232 72.8958
R4144 VDD.n2588 VDD.n1231 72.8958
R4145 VDD.n2588 VDD.n1230 72.8958
R4146 VDD.n2588 VDD.n1229 72.8958
R4147 VDD.n2975 VDD.n2974 72.8958
R4148 VDD.n2975 VDD.n923 72.8958
R4149 VDD.n2975 VDD.n922 72.8958
R4150 VDD.n2975 VDD.n921 72.8958
R4151 VDD.n2975 VDD.n920 72.8958
R4152 VDD.n2975 VDD.n919 72.8958
R4153 VDD.n2975 VDD.n918 72.8958
R4154 VDD.n2975 VDD.n917 72.8958
R4155 VDD.n2975 VDD.n916 72.8958
R4156 VDD.n2975 VDD.n915 72.8958
R4157 VDD.n3289 VDD.n2976 72.8958
R4158 VDD.n3287 VDD.n2976 72.8958
R4159 VDD.n3281 VDD.n2976 72.8958
R4160 VDD.n3279 VDD.n2976 72.8958
R4161 VDD.n3273 VDD.n2976 72.8958
R4162 VDD.n3271 VDD.n2976 72.8958
R4163 VDD.n3265 VDD.n2976 72.8958
R4164 VDD.n3263 VDD.n2976 72.8958
R4165 VDD.n3256 VDD.n2976 72.8958
R4166 VDD.n3254 VDD.n2976 72.8958
R4167 VDD.n483 VDD.n473 72.8958
R4168 VDD.n3725 VDD.n473 72.8958
R4169 VDD.n477 VDD.n473 72.8958
R4170 VDD.n3732 VDD.n473 72.8958
R4171 VDD.n3735 VDD.n473 72.8958
R4172 VDD.n3644 VDD.n473 72.8958
R4173 VDD.n3649 VDD.n473 72.8958
R4174 VDD.n3643 VDD.n473 72.8958
R4175 VDD.n3656 VDD.n473 72.8958
R4176 VDD.n3659 VDD.n473 72.8958
R4177 VDD.n3134 VDD.n2976 72.8958
R4178 VDD.n3137 VDD.n2976 72.8958
R4179 VDD.n3143 VDD.n2976 72.8958
R4180 VDD.n3145 VDD.n2976 72.8958
R4181 VDD.n3151 VDD.n2976 72.8958
R4182 VDD.n3153 VDD.n2976 72.8958
R4183 VDD.n3159 VDD.n2976 72.8958
R4184 VDD.n3161 VDD.n2976 72.8958
R4185 VDD.n3168 VDD.n2976 72.8958
R4186 VDD.n3682 VDD.n473 72.8958
R4187 VDD.n617 VDD.n473 72.8958
R4188 VDD.n3690 VDD.n473 72.8958
R4189 VDD.n612 VDD.n473 72.8958
R4190 VDD.n3697 VDD.n473 72.8958
R4191 VDD.n608 VDD.n473 72.8958
R4192 VDD.n3704 VDD.n473 72.8958
R4193 VDD.n495 VDD.n473 72.8958
R4194 VDD.n3711 VDD.n473 72.8958
R4195 VDD.n492 VDD.n473 72.8958
R4196 VDD.n2975 VDD.n914 72.8958
R4197 VDD.n2975 VDD.n913 72.8958
R4198 VDD.n2975 VDD.n912 72.8958
R4199 VDD.n2975 VDD.n911 72.8958
R4200 VDD.n2975 VDD.n910 72.8958
R4201 VDD.n2975 VDD.n909 72.8958
R4202 VDD.n2975 VDD.n908 72.8958
R4203 VDD.n2975 VDD.n907 72.8958
R4204 VDD.n2975 VDD.n906 72.8958
R4205 VDD.n2975 VDD.n905 72.8958
R4206 VDD.n2589 VDD.n2588 72.8958
R4207 VDD.n2588 VDD.n1220 72.8958
R4208 VDD.n2588 VDD.n1221 72.8958
R4209 VDD.n2588 VDD.n1222 72.8958
R4210 VDD.n2588 VDD.n1223 72.8958
R4211 VDD.n2588 VDD.n1224 72.8958
R4212 VDD.n2588 VDD.n1225 72.8958
R4213 VDD.n2588 VDD.n1226 72.8958
R4214 VDD.n2588 VDD.n1227 72.8958
R4215 VDD.n1730 VDD.n1729 66.2847
R4216 VDD.n1729 VDD.n1627 66.2847
R4217 VDD.n1729 VDD.n1628 66.2847
R4218 VDD.n1729 VDD.n1629 66.2847
R4219 VDD.n1729 VDD.n1630 66.2847
R4220 VDD.n1729 VDD.n1631 66.2847
R4221 VDD.n1729 VDD.n1632 66.2847
R4222 VDD.n1729 VDD.n1633 66.2847
R4223 VDD.n1729 VDD.n1634 66.2847
R4224 VDD.n1729 VDD.n1635 66.2847
R4225 VDD.n1729 VDD.n1636 66.2847
R4226 VDD.n1729 VDD.n1637 66.2847
R4227 VDD.n1729 VDD.n1638 66.2847
R4228 VDD.n1729 VDD.n1639 66.2847
R4229 VDD.n1308 VDD.n1283 66.2847
R4230 VDD.n1308 VDD.n1307 66.2847
R4231 VDD.n1308 VDD.n1305 66.2847
R4232 VDD.n1308 VDD.n1304 66.2847
R4233 VDD.n1308 VDD.n1302 66.2847
R4234 VDD.n1308 VDD.n1301 66.2847
R4235 VDD.n1308 VDD.n1299 66.2847
R4236 VDD.n1308 VDD.n1298 66.2847
R4237 VDD.n1308 VDD.n1296 66.2847
R4238 VDD.n1308 VDD.n1295 66.2847
R4239 VDD.n1308 VDD.n1293 66.2847
R4240 VDD.n1308 VDD.n1292 66.2847
R4241 VDD.n1308 VDD.n1290 66.2847
R4242 VDD.n1308 VDD.n1289 66.2847
R4243 VDD.n1308 VDD.n1287 66.2847
R4244 VDD.n602 VDD.n601 66.2847
R4245 VDD.n601 VDD.n500 66.2847
R4246 VDD.n601 VDD.n501 66.2847
R4247 VDD.n601 VDD.n502 66.2847
R4248 VDD.n601 VDD.n503 66.2847
R4249 VDD.n601 VDD.n504 66.2847
R4250 VDD.n601 VDD.n505 66.2847
R4251 VDD.n601 VDD.n506 66.2847
R4252 VDD.n601 VDD.n507 66.2847
R4253 VDD.n601 VDD.n508 66.2847
R4254 VDD.n601 VDD.n509 66.2847
R4255 VDD.n601 VDD.n510 66.2847
R4256 VDD.n601 VDD.n511 66.2847
R4257 VDD.n601 VDD.n512 66.2847
R4258 VDD.n4050 VDD.n4049 66.2847
R4259 VDD.n4050 VDD.n193 66.2847
R4260 VDD.n4050 VDD.n192 66.2847
R4261 VDD.n4050 VDD.n191 66.2847
R4262 VDD.n4050 VDD.n190 66.2847
R4263 VDD.n4050 VDD.n189 66.2847
R4264 VDD.n4050 VDD.n188 66.2847
R4265 VDD.n4050 VDD.n187 66.2847
R4266 VDD.n4050 VDD.n186 66.2847
R4267 VDD.n4050 VDD.n185 66.2847
R4268 VDD.n4050 VDD.n184 66.2847
R4269 VDD.n4050 VDD.n183 66.2847
R4270 VDD.n4050 VDD.n182 66.2847
R4271 VDD.n4050 VDD.n181 66.2847
R4272 VDD.n4050 VDD.n180 66.2847
R4273 VDD.n220 VDD.n180 52.4337
R4274 VDD.n224 VDD.n181 52.4337
R4275 VDD.n230 VDD.n182 52.4337
R4276 VDD.n234 VDD.n183 52.4337
R4277 VDD.n240 VDD.n184 52.4337
R4278 VDD.n244 VDD.n185 52.4337
R4279 VDD.n250 VDD.n186 52.4337
R4280 VDD.n254 VDD.n187 52.4337
R4281 VDD.n260 VDD.n188 52.4337
R4282 VDD.n264 VDD.n189 52.4337
R4283 VDD.n270 VDD.n190 52.4337
R4284 VDD.n274 VDD.n191 52.4337
R4285 VDD.n280 VDD.n192 52.4337
R4286 VDD.n283 VDD.n193 52.4337
R4287 VDD.n4049 VDD.n4048 52.4337
R4288 VDD.n603 VDD.n602 52.4337
R4289 VDD.n514 VDD.n500 52.4337
R4290 VDD.n595 VDD.n501 52.4337
R4291 VDD.n591 VDD.n502 52.4337
R4292 VDD.n587 VDD.n503 52.4337
R4293 VDD.n583 VDD.n504 52.4337
R4294 VDD.n579 VDD.n505 52.4337
R4295 VDD.n575 VDD.n506 52.4337
R4296 VDD.n571 VDD.n507 52.4337
R4297 VDD.n567 VDD.n508 52.4337
R4298 VDD.n563 VDD.n509 52.4337
R4299 VDD.n559 VDD.n510 52.4337
R4300 VDD.n555 VDD.n511 52.4337
R4301 VDD.n551 VDD.n512 52.4337
R4302 VDD.n1287 VDD.n1244 52.4337
R4303 VDD.n1289 VDD.n1288 52.4337
R4304 VDD.n1290 VDD.n1249 52.4337
R4305 VDD.n1292 VDD.n1291 52.4337
R4306 VDD.n1293 VDD.n1254 52.4337
R4307 VDD.n1295 VDD.n1294 52.4337
R4308 VDD.n1296 VDD.n1261 52.4337
R4309 VDD.n1298 VDD.n1297 52.4337
R4310 VDD.n1299 VDD.n1266 52.4337
R4311 VDD.n1301 VDD.n1300 52.4337
R4312 VDD.n1302 VDD.n1271 52.4337
R4313 VDD.n1304 VDD.n1303 52.4337
R4314 VDD.n1305 VDD.n1276 52.4337
R4315 VDD.n1307 VDD.n1306 52.4337
R4316 VDD.n2524 VDD.n1283 52.4337
R4317 VDD.n1731 VDD.n1730 52.4337
R4318 VDD.n1641 VDD.n1627 52.4337
R4319 VDD.n1645 VDD.n1628 52.4337
R4320 VDD.n1647 VDD.n1629 52.4337
R4321 VDD.n1651 VDD.n1630 52.4337
R4322 VDD.n1653 VDD.n1631 52.4337
R4323 VDD.n1707 VDD.n1632 52.4337
R4324 VDD.n1658 VDD.n1633 52.4337
R4325 VDD.n1662 VDD.n1634 52.4337
R4326 VDD.n1664 VDD.n1635 52.4337
R4327 VDD.n1668 VDD.n1636 52.4337
R4328 VDD.n1670 VDD.n1637 52.4337
R4329 VDD.n1674 VDD.n1638 52.4337
R4330 VDD.n1676 VDD.n1639 52.4337
R4331 VDD.n1730 VDD.n1626 52.4337
R4332 VDD.n1644 VDD.n1627 52.4337
R4333 VDD.n1646 VDD.n1628 52.4337
R4334 VDD.n1650 VDD.n1629 52.4337
R4335 VDD.n1652 VDD.n1630 52.4337
R4336 VDD.n1656 VDD.n1631 52.4337
R4337 VDD.n1657 VDD.n1632 52.4337
R4338 VDD.n1661 VDD.n1633 52.4337
R4339 VDD.n1663 VDD.n1634 52.4337
R4340 VDD.n1667 VDD.n1635 52.4337
R4341 VDD.n1669 VDD.n1636 52.4337
R4342 VDD.n1673 VDD.n1637 52.4337
R4343 VDD.n1675 VDD.n1638 52.4337
R4344 VDD.n1679 VDD.n1639 52.4337
R4345 VDD.n1283 VDD.n1280 52.4337
R4346 VDD.n1307 VDD.n1277 52.4337
R4347 VDD.n1305 VDD.n1275 52.4337
R4348 VDD.n1304 VDD.n1272 52.4337
R4349 VDD.n1302 VDD.n1270 52.4337
R4350 VDD.n1301 VDD.n1267 52.4337
R4351 VDD.n1299 VDD.n1265 52.4337
R4352 VDD.n1298 VDD.n1262 52.4337
R4353 VDD.n1296 VDD.n1258 52.4337
R4354 VDD.n1295 VDD.n1255 52.4337
R4355 VDD.n1293 VDD.n1253 52.4337
R4356 VDD.n1292 VDD.n1250 52.4337
R4357 VDD.n1290 VDD.n1248 52.4337
R4358 VDD.n1289 VDD.n1245 52.4337
R4359 VDD.n1287 VDD.n1243 52.4337
R4360 VDD.n602 VDD.n499 52.4337
R4361 VDD.n596 VDD.n500 52.4337
R4362 VDD.n592 VDD.n501 52.4337
R4363 VDD.n588 VDD.n502 52.4337
R4364 VDD.n584 VDD.n503 52.4337
R4365 VDD.n580 VDD.n504 52.4337
R4366 VDD.n576 VDD.n505 52.4337
R4367 VDD.n572 VDD.n506 52.4337
R4368 VDD.n568 VDD.n507 52.4337
R4369 VDD.n564 VDD.n508 52.4337
R4370 VDD.n560 VDD.n509 52.4337
R4371 VDD.n556 VDD.n510 52.4337
R4372 VDD.n552 VDD.n511 52.4337
R4373 VDD.n543 VDD.n512 52.4337
R4374 VDD.n4049 VDD.n194 52.4337
R4375 VDD.n281 VDD.n193 52.4337
R4376 VDD.n275 VDD.n192 52.4337
R4377 VDD.n271 VDD.n191 52.4337
R4378 VDD.n265 VDD.n190 52.4337
R4379 VDD.n261 VDD.n189 52.4337
R4380 VDD.n255 VDD.n188 52.4337
R4381 VDD.n251 VDD.n187 52.4337
R4382 VDD.n245 VDD.n186 52.4337
R4383 VDD.n241 VDD.n185 52.4337
R4384 VDD.n235 VDD.n184 52.4337
R4385 VDD.n231 VDD.n183 52.4337
R4386 VDD.n225 VDD.n182 52.4337
R4387 VDD.n221 VDD.n181 52.4337
R4388 VDD.n215 VDD.n180 52.4337
R4389 VDD.n3713 VDD.n492 39.2114
R4390 VDD.n3711 VDD.n3710 39.2114
R4391 VDD.n3706 VDD.n495 39.2114
R4392 VDD.n3704 VDD.n3703 39.2114
R4393 VDD.n3699 VDD.n608 39.2114
R4394 VDD.n3697 VDD.n3696 39.2114
R4395 VDD.n3692 VDD.n612 39.2114
R4396 VDD.n3690 VDD.n3689 39.2114
R4397 VDD.n3684 VDD.n617 39.2114
R4398 VDD.n3682 VDD.n3681 39.2114
R4399 VDD.n3134 VDD.n903 39.2114
R4400 VDD.n3138 VDD.n3137 39.2114
R4401 VDD.n3143 VDD.n3142 39.2114
R4402 VDD.n3146 VDD.n3145 39.2114
R4403 VDD.n3151 VDD.n3150 39.2114
R4404 VDD.n3154 VDD.n3153 39.2114
R4405 VDD.n3159 VDD.n3158 39.2114
R4406 VDD.n3162 VDD.n3161 39.2114
R4407 VDD.n3168 VDD.n3167 39.2114
R4408 VDD.n3659 VDD.n3658 39.2114
R4409 VDD.n3656 VDD.n3655 39.2114
R4410 VDD.n3651 VDD.n3643 39.2114
R4411 VDD.n3649 VDD.n3648 39.2114
R4412 VDD.n3644 VDD.n472 39.2114
R4413 VDD.n3735 VDD.n3734 39.2114
R4414 VDD.n3732 VDD.n3731 39.2114
R4415 VDD.n3727 VDD.n477 39.2114
R4416 VDD.n3725 VDD.n3724 39.2114
R4417 VDD.n3720 VDD.n483 39.2114
R4418 VDD.n3289 VDD.n2979 39.2114
R4419 VDD.n3288 VDD.n3287 39.2114
R4420 VDD.n3281 VDD.n2981 39.2114
R4421 VDD.n3280 VDD.n3279 39.2114
R4422 VDD.n3273 VDD.n2983 39.2114
R4423 VDD.n3272 VDD.n3271 39.2114
R4424 VDD.n3265 VDD.n2985 39.2114
R4425 VDD.n3264 VDD.n3263 39.2114
R4426 VDD.n3256 VDD.n2987 39.2114
R4427 VDD.n3255 VDD.n3254 39.2114
R4428 VDD.n2898 VDD.n915 39.2114
R4429 VDD.n2894 VDD.n916 39.2114
R4430 VDD.n2890 VDD.n917 39.2114
R4431 VDD.n2886 VDD.n918 39.2114
R4432 VDD.n2882 VDD.n919 39.2114
R4433 VDD.n2878 VDD.n920 39.2114
R4434 VDD.n2874 VDD.n921 39.2114
R4435 VDD.n2870 VDD.n922 39.2114
R4436 VDD.n2865 VDD.n923 39.2114
R4437 VDD.n2974 VDD.n2973 39.2114
R4438 VDD.n2160 VDD.n1238 39.2114
R4439 VDD.n2164 VDD.n1237 39.2114
R4440 VDD.n2168 VDD.n1236 39.2114
R4441 VDD.n2172 VDD.n1235 39.2114
R4442 VDD.n2176 VDD.n1234 39.2114
R4443 VDD.n2503 VDD.n1233 39.2114
R4444 VDD.n2499 VDD.n1232 39.2114
R4445 VDD.n2495 VDD.n1231 39.2114
R4446 VDD.n2491 VDD.n1230 39.2114
R4447 VDD.n2486 VDD.n1229 39.2114
R4448 VDD.n2163 VDD.n1238 39.2114
R4449 VDD.n2167 VDD.n1237 39.2114
R4450 VDD.n2171 VDD.n1236 39.2114
R4451 VDD.n2175 VDD.n1235 39.2114
R4452 VDD.n2502 VDD.n1234 39.2114
R4453 VDD.n2500 VDD.n1233 39.2114
R4454 VDD.n2496 VDD.n1232 39.2114
R4455 VDD.n2492 VDD.n1231 39.2114
R4456 VDD.n2487 VDD.n1230 39.2114
R4457 VDD.n2483 VDD.n1229 39.2114
R4458 VDD.n2974 VDD.n924 39.2114
R4459 VDD.n2869 VDD.n923 39.2114
R4460 VDD.n2873 VDD.n922 39.2114
R4461 VDD.n2877 VDD.n921 39.2114
R4462 VDD.n2881 VDD.n920 39.2114
R4463 VDD.n2885 VDD.n919 39.2114
R4464 VDD.n2889 VDD.n918 39.2114
R4465 VDD.n2893 VDD.n917 39.2114
R4466 VDD.n2897 VDD.n916 39.2114
R4467 VDD.n2901 VDD.n915 39.2114
R4468 VDD.n3290 VDD.n3289 39.2114
R4469 VDD.n3287 VDD.n3286 39.2114
R4470 VDD.n3282 VDD.n3281 39.2114
R4471 VDD.n3279 VDD.n3278 39.2114
R4472 VDD.n3274 VDD.n3273 39.2114
R4473 VDD.n3271 VDD.n3270 39.2114
R4474 VDD.n3266 VDD.n3265 39.2114
R4475 VDD.n3263 VDD.n3262 39.2114
R4476 VDD.n3257 VDD.n3256 39.2114
R4477 VDD.n3254 VDD.n3253 39.2114
R4478 VDD.n483 VDD.n478 39.2114
R4479 VDD.n3726 VDD.n3725 39.2114
R4480 VDD.n477 VDD.n475 39.2114
R4481 VDD.n3733 VDD.n3732 39.2114
R4482 VDD.n3736 VDD.n3735 39.2114
R4483 VDD.n3645 VDD.n3644 39.2114
R4484 VDD.n3650 VDD.n3649 39.2114
R4485 VDD.n3643 VDD.n3641 39.2114
R4486 VDD.n3657 VDD.n3656 39.2114
R4487 VDD.n3660 VDD.n3659 39.2114
R4488 VDD.n3135 VDD.n3134 39.2114
R4489 VDD.n3137 VDD.n3131 39.2114
R4490 VDD.n3144 VDD.n3143 39.2114
R4491 VDD.n3145 VDD.n3129 39.2114
R4492 VDD.n3152 VDD.n3151 39.2114
R4493 VDD.n3153 VDD.n3127 39.2114
R4494 VDD.n3160 VDD.n3159 39.2114
R4495 VDD.n3161 VDD.n3123 39.2114
R4496 VDD.n3169 VDD.n3168 39.2114
R4497 VDD.n3683 VDD.n3682 39.2114
R4498 VDD.n617 VDD.n613 39.2114
R4499 VDD.n3691 VDD.n3690 39.2114
R4500 VDD.n612 VDD.n610 39.2114
R4501 VDD.n3698 VDD.n3697 39.2114
R4502 VDD.n608 VDD.n496 39.2114
R4503 VDD.n3705 VDD.n3704 39.2114
R4504 VDD.n495 VDD.n493 39.2114
R4505 VDD.n3712 VDD.n3711 39.2114
R4506 VDD.n492 VDD.n489 39.2114
R4507 VDD.n2961 VDD.n905 39.2114
R4508 VDD.n2957 VDD.n906 39.2114
R4509 VDD.n2953 VDD.n907 39.2114
R4510 VDD.n2949 VDD.n908 39.2114
R4511 VDD.n2945 VDD.n909 39.2114
R4512 VDD.n2941 VDD.n910 39.2114
R4513 VDD.n2937 VDD.n911 39.2114
R4514 VDD.n2933 VDD.n912 39.2114
R4515 VDD.n2928 VDD.n913 39.2114
R4516 VDD.n2924 VDD.n914 39.2114
R4517 VDD.n2590 VDD.n2589 39.2114
R4518 VDD.n1239 VDD.n1220 39.2114
R4519 VDD.n2582 VDD.n1221 39.2114
R4520 VDD.n2578 VDD.n1222 39.2114
R4521 VDD.n2574 VDD.n1223 39.2114
R4522 VDD.n2312 VDD.n1224 39.2114
R4523 VDD.n2316 VDD.n1225 39.2114
R4524 VDD.n2320 VDD.n1226 39.2114
R4525 VDD.n2324 VDD.n1227 39.2114
R4526 VDD.n2927 VDD.n914 39.2114
R4527 VDD.n2932 VDD.n913 39.2114
R4528 VDD.n2936 VDD.n912 39.2114
R4529 VDD.n2940 VDD.n911 39.2114
R4530 VDD.n2944 VDD.n910 39.2114
R4531 VDD.n2948 VDD.n909 39.2114
R4532 VDD.n2952 VDD.n908 39.2114
R4533 VDD.n2956 VDD.n907 39.2114
R4534 VDD.n2960 VDD.n906 39.2114
R4535 VDD.n2963 VDD.n905 39.2114
R4536 VDD.n2589 VDD.n1219 39.2114
R4537 VDD.n2583 VDD.n1220 39.2114
R4538 VDD.n2579 VDD.n1221 39.2114
R4539 VDD.n2575 VDD.n1222 39.2114
R4540 VDD.n2311 VDD.n1223 39.2114
R4541 VDD.n2315 VDD.n1224 39.2114
R4542 VDD.n2319 VDD.n1225 39.2114
R4543 VDD.n2323 VDD.n1226 39.2114
R4544 VDD.n2326 VDD.n1227 39.2114
R4545 VDD.n2550 VDD.n1260 37.2369
R4546 VDD.n2526 VDD.n1282 37.2369
R4547 VDD.n1683 VDD.n1682 37.2369
R4548 VDD.n1710 VDD.n1709 37.2369
R4549 VDD.n578 VDD.n528 37.2369
R4550 VDD.n547 VDD.n546 37.2369
R4551 VDD.n197 VDD.n196 37.2369
R4552 VDD.n207 VDD.n206 37.2369
R4553 VDD.n3172 VDD.n3171 32.4688
R4554 VDD.n3680 VDD.n3679 32.4688
R4555 VDD.n3297 VDD.n902 32.4688
R4556 VDD.n3716 VDD.n3715 32.4688
R4557 VDD.n3662 VDD.n3661 32.4688
R4558 VDD.n3721 VDD.n482 32.4688
R4559 VDD.n3252 VDD.n3251 32.4688
R4560 VDD.n3293 VDD.n3292 32.4688
R4561 VDD.n2903 VDD.n2900 32.4688
R4562 VDD.n2972 VDD.n2971 32.4688
R4563 VDD.n2484 VDD.n2481 32.4688
R4564 VDD.n2161 VDD.n1212 32.4688
R4565 VDD.n2592 VDD.n2591 32.4688
R4566 VDD.n2965 VDD.n2964 32.4688
R4567 VDD.n2925 VDD.n2922 32.4688
R4568 VDD.n2330 VDD.n2328 32.4688
R4569 VDD.n2310 VDD.n2309 30.449
R4570 VDD.n2930 VDD.n936 30.449
R4571 VDD.n3259 VDD.n2989 30.449
R4572 VDD.n3686 VDD.n615 30.449
R4573 VDD.n3165 VDD.n3125 30.449
R4574 VDD.n481 VDD.n480 30.449
R4575 VDD.n2489 VDD.n2180 30.449
R4576 VDD.n2867 VDD.n2864 30.449
R4577 VDD.n1729 VDD.n1621 29.3387
R4578 VDD.n2522 VDD.n1308 29.3387
R4579 VDD.n601 VDD.n466 29.3387
R4580 VDD.n4051 VDD.n4050 29.3387
R4581 VDD.n2588 VDD.t28 25.1476
R4582 VDD.t9 VDD.n473 25.1476
R4583 VDD.n2588 VDD.n1214 19.734
R4584 VDD.n2975 VDD.n904 19.734
R4585 VDD.n3295 VDD.n2976 19.734
R4586 VDD.n3718 VDD.n473 19.734
R4587 VDD.n1740 VDD.n1619 19.3944
R4588 VDD.n1740 VDD.n1617 19.3944
R4589 VDD.n1744 VDD.n1617 19.3944
R4590 VDD.n1744 VDD.n1607 19.3944
R4591 VDD.n1756 VDD.n1607 19.3944
R4592 VDD.n1756 VDD.n1605 19.3944
R4593 VDD.n1760 VDD.n1605 19.3944
R4594 VDD.n1760 VDD.n1595 19.3944
R4595 VDD.n1772 VDD.n1595 19.3944
R4596 VDD.n1772 VDD.n1593 19.3944
R4597 VDD.n1776 VDD.n1593 19.3944
R4598 VDD.n1776 VDD.n1583 19.3944
R4599 VDD.n1788 VDD.n1583 19.3944
R4600 VDD.n1788 VDD.n1581 19.3944
R4601 VDD.n1792 VDD.n1581 19.3944
R4602 VDD.n1792 VDD.n1571 19.3944
R4603 VDD.n1804 VDD.n1571 19.3944
R4604 VDD.n1804 VDD.n1569 19.3944
R4605 VDD.n1808 VDD.n1569 19.3944
R4606 VDD.n1808 VDD.n1559 19.3944
R4607 VDD.n1820 VDD.n1559 19.3944
R4608 VDD.n1820 VDD.n1557 19.3944
R4609 VDD.n1824 VDD.n1557 19.3944
R4610 VDD.n1824 VDD.n1547 19.3944
R4611 VDD.n1836 VDD.n1547 19.3944
R4612 VDD.n1836 VDD.n1545 19.3944
R4613 VDD.n1840 VDD.n1545 19.3944
R4614 VDD.n1840 VDD.n1534 19.3944
R4615 VDD.n1852 VDD.n1534 19.3944
R4616 VDD.n1852 VDD.n1532 19.3944
R4617 VDD.n1856 VDD.n1532 19.3944
R4618 VDD.n1856 VDD.n1523 19.3944
R4619 VDD.n1868 VDD.n1523 19.3944
R4620 VDD.n1868 VDD.n1521 19.3944
R4621 VDD.n1872 VDD.n1521 19.3944
R4622 VDD.n1872 VDD.n1511 19.3944
R4623 VDD.n1884 VDD.n1511 19.3944
R4624 VDD.n1884 VDD.n1509 19.3944
R4625 VDD.n1888 VDD.n1509 19.3944
R4626 VDD.n1888 VDD.n1499 19.3944
R4627 VDD.n1900 VDD.n1499 19.3944
R4628 VDD.n1900 VDD.n1497 19.3944
R4629 VDD.n1904 VDD.n1497 19.3944
R4630 VDD.n1904 VDD.n1487 19.3944
R4631 VDD.n1916 VDD.n1487 19.3944
R4632 VDD.n1916 VDD.n1485 19.3944
R4633 VDD.n1920 VDD.n1485 19.3944
R4634 VDD.n1920 VDD.n1475 19.3944
R4635 VDD.n1932 VDD.n1475 19.3944
R4636 VDD.n1932 VDD.n1473 19.3944
R4637 VDD.n1936 VDD.n1473 19.3944
R4638 VDD.n1936 VDD.n1463 19.3944
R4639 VDD.n1961 VDD.n1463 19.3944
R4640 VDD.n1961 VDD.n1461 19.3944
R4641 VDD.n1965 VDD.n1461 19.3944
R4642 VDD.n1965 VDD.n1451 19.3944
R4643 VDD.n1977 VDD.n1451 19.3944
R4644 VDD.n1977 VDD.n1449 19.3944
R4645 VDD.n1981 VDD.n1449 19.3944
R4646 VDD.n1981 VDD.n1439 19.3944
R4647 VDD.n1993 VDD.n1439 19.3944
R4648 VDD.n1993 VDD.n1437 19.3944
R4649 VDD.n1997 VDD.n1437 19.3944
R4650 VDD.n1997 VDD.n1428 19.3944
R4651 VDD.n2010 VDD.n1428 19.3944
R4652 VDD.n2010 VDD.n1426 19.3944
R4653 VDD.n2014 VDD.n1426 19.3944
R4654 VDD.n2014 VDD.n1416 19.3944
R4655 VDD.n2026 VDD.n1416 19.3944
R4656 VDD.n2026 VDD.n1414 19.3944
R4657 VDD.n2030 VDD.n1414 19.3944
R4658 VDD.n2030 VDD.n1404 19.3944
R4659 VDD.n2042 VDD.n1404 19.3944
R4660 VDD.n2042 VDD.n1402 19.3944
R4661 VDD.n2046 VDD.n1402 19.3944
R4662 VDD.n2046 VDD.n1392 19.3944
R4663 VDD.n2058 VDD.n1392 19.3944
R4664 VDD.n2058 VDD.n1390 19.3944
R4665 VDD.n2062 VDD.n1390 19.3944
R4666 VDD.n2062 VDD.n1380 19.3944
R4667 VDD.n2074 VDD.n1380 19.3944
R4668 VDD.n2074 VDD.n1378 19.3944
R4669 VDD.n2078 VDD.n1378 19.3944
R4670 VDD.n2078 VDD.n1367 19.3944
R4671 VDD.n2090 VDD.n1367 19.3944
R4672 VDD.n2090 VDD.n1365 19.3944
R4673 VDD.n2094 VDD.n1365 19.3944
R4674 VDD.n2094 VDD.n1356 19.3944
R4675 VDD.n2106 VDD.n1356 19.3944
R4676 VDD.n2106 VDD.n1354 19.3944
R4677 VDD.n2110 VDD.n1354 19.3944
R4678 VDD.n2110 VDD.n1344 19.3944
R4679 VDD.n2122 VDD.n1344 19.3944
R4680 VDD.n2122 VDD.n1342 19.3944
R4681 VDD.n2126 VDD.n1342 19.3944
R4682 VDD.n2126 VDD.n1332 19.3944
R4683 VDD.n2138 VDD.n1332 19.3944
R4684 VDD.n2138 VDD.n1329 19.3944
R4685 VDD.n2143 VDD.n1329 19.3944
R4686 VDD.n2143 VDD.n1330 19.3944
R4687 VDD.n1330 VDD.n1320 19.3944
R4688 VDD.n2157 VDD.n1320 19.3944
R4689 VDD.n2157 VDD.n1317 19.3944
R4690 VDD.n2510 VDD.n1317 19.3944
R4691 VDD.n2510 VDD.n1318 19.3944
R4692 VDD.n1318 VDD.n1285 19.3944
R4693 VDD.n2569 VDD.n2568 19.3944
R4694 VDD.n2568 VDD.n2567 19.3944
R4695 VDD.n2567 VDD.n1246 19.3944
R4696 VDD.n2563 VDD.n1246 19.3944
R4697 VDD.n2563 VDD.n2562 19.3944
R4698 VDD.n2562 VDD.n2561 19.3944
R4699 VDD.n2561 VDD.n1251 19.3944
R4700 VDD.n2557 VDD.n1251 19.3944
R4701 VDD.n2557 VDD.n2556 19.3944
R4702 VDD.n2556 VDD.n2555 19.3944
R4703 VDD.n2555 VDD.n1256 19.3944
R4704 VDD.n2551 VDD.n1256 19.3944
R4705 VDD.n2549 VDD.n1263 19.3944
R4706 VDD.n2545 VDD.n1263 19.3944
R4707 VDD.n2545 VDD.n2544 19.3944
R4708 VDD.n2544 VDD.n2543 19.3944
R4709 VDD.n2543 VDD.n1268 19.3944
R4710 VDD.n2539 VDD.n1268 19.3944
R4711 VDD.n2539 VDD.n2538 19.3944
R4712 VDD.n2538 VDD.n2537 19.3944
R4713 VDD.n2537 VDD.n1273 19.3944
R4714 VDD.n2533 VDD.n1273 19.3944
R4715 VDD.n2533 VDD.n2532 19.3944
R4716 VDD.n2532 VDD.n2531 19.3944
R4717 VDD.n2531 VDD.n1278 19.3944
R4718 VDD.n2527 VDD.n1278 19.3944
R4719 VDD.n1706 VDD.n1659 19.3944
R4720 VDD.n1702 VDD.n1659 19.3944
R4721 VDD.n1702 VDD.n1701 19.3944
R4722 VDD.n1701 VDD.n1700 19.3944
R4723 VDD.n1700 VDD.n1665 19.3944
R4724 VDD.n1696 VDD.n1665 19.3944
R4725 VDD.n1696 VDD.n1695 19.3944
R4726 VDD.n1695 VDD.n1694 19.3944
R4727 VDD.n1694 VDD.n1671 19.3944
R4728 VDD.n1690 VDD.n1671 19.3944
R4729 VDD.n1690 VDD.n1689 19.3944
R4730 VDD.n1689 VDD.n1688 19.3944
R4731 VDD.n1688 VDD.n1677 19.3944
R4732 VDD.n1684 VDD.n1677 19.3944
R4733 VDD.n1732 VDD.n1625 19.3944
R4734 VDD.n1727 VDD.n1625 19.3944
R4735 VDD.n1727 VDD.n1642 19.3944
R4736 VDD.n1723 VDD.n1642 19.3944
R4737 VDD.n1723 VDD.n1722 19.3944
R4738 VDD.n1722 VDD.n1721 19.3944
R4739 VDD.n1721 VDD.n1648 19.3944
R4740 VDD.n1717 VDD.n1648 19.3944
R4741 VDD.n1717 VDD.n1716 19.3944
R4742 VDD.n1716 VDD.n1715 19.3944
R4743 VDD.n1715 VDD.n1654 19.3944
R4744 VDD.n1711 VDD.n1654 19.3944
R4745 VDD.n1736 VDD.n1623 19.3944
R4746 VDD.n1736 VDD.n1613 19.3944
R4747 VDD.n1748 VDD.n1613 19.3944
R4748 VDD.n1748 VDD.n1611 19.3944
R4749 VDD.n1752 VDD.n1611 19.3944
R4750 VDD.n1752 VDD.n1601 19.3944
R4751 VDD.n1764 VDD.n1601 19.3944
R4752 VDD.n1764 VDD.n1599 19.3944
R4753 VDD.n1768 VDD.n1599 19.3944
R4754 VDD.n1768 VDD.n1589 19.3944
R4755 VDD.n1780 VDD.n1589 19.3944
R4756 VDD.n1780 VDD.n1587 19.3944
R4757 VDD.n1784 VDD.n1587 19.3944
R4758 VDD.n1784 VDD.n1577 19.3944
R4759 VDD.n1796 VDD.n1577 19.3944
R4760 VDD.n1796 VDD.n1575 19.3944
R4761 VDD.n1800 VDD.n1575 19.3944
R4762 VDD.n1800 VDD.n1565 19.3944
R4763 VDD.n1812 VDD.n1565 19.3944
R4764 VDD.n1812 VDD.n1563 19.3944
R4765 VDD.n1816 VDD.n1563 19.3944
R4766 VDD.n1816 VDD.n1553 19.3944
R4767 VDD.n1828 VDD.n1553 19.3944
R4768 VDD.n1828 VDD.n1551 19.3944
R4769 VDD.n1832 VDD.n1551 19.3944
R4770 VDD.n1832 VDD.n1541 19.3944
R4771 VDD.n1844 VDD.n1541 19.3944
R4772 VDD.n1844 VDD.n1539 19.3944
R4773 VDD.n1848 VDD.n1539 19.3944
R4774 VDD.n1848 VDD.n1529 19.3944
R4775 VDD.n1860 VDD.n1529 19.3944
R4776 VDD.n1860 VDD.n1527 19.3944
R4777 VDD.n1864 VDD.n1527 19.3944
R4778 VDD.n1864 VDD.n1517 19.3944
R4779 VDD.n1876 VDD.n1517 19.3944
R4780 VDD.n1876 VDD.n1515 19.3944
R4781 VDD.n1880 VDD.n1515 19.3944
R4782 VDD.n1880 VDD.n1505 19.3944
R4783 VDD.n1892 VDD.n1505 19.3944
R4784 VDD.n1892 VDD.n1503 19.3944
R4785 VDD.n1896 VDD.n1503 19.3944
R4786 VDD.n1896 VDD.n1493 19.3944
R4787 VDD.n1908 VDD.n1493 19.3944
R4788 VDD.n1908 VDD.n1491 19.3944
R4789 VDD.n1912 VDD.n1491 19.3944
R4790 VDD.n1912 VDD.n1481 19.3944
R4791 VDD.n1924 VDD.n1481 19.3944
R4792 VDD.n1924 VDD.n1479 19.3944
R4793 VDD.n1928 VDD.n1479 19.3944
R4794 VDD.n1928 VDD.n1469 19.3944
R4795 VDD.n1940 VDD.n1469 19.3944
R4796 VDD.n1940 VDD.n1467 19.3944
R4797 VDD.n1958 VDD.n1467 19.3944
R4798 VDD.n1958 VDD.n1457 19.3944
R4799 VDD.n1969 VDD.n1457 19.3944
R4800 VDD.n1969 VDD.n1455 19.3944
R4801 VDD.n1973 VDD.n1455 19.3944
R4802 VDD.n1973 VDD.n1445 19.3944
R4803 VDD.n1985 VDD.n1445 19.3944
R4804 VDD.n1985 VDD.n1443 19.3944
R4805 VDD.n1989 VDD.n1443 19.3944
R4806 VDD.n1989 VDD.n1433 19.3944
R4807 VDD.n2002 VDD.n1433 19.3944
R4808 VDD.n2002 VDD.n1431 19.3944
R4809 VDD.n2006 VDD.n1431 19.3944
R4810 VDD.n2006 VDD.n1422 19.3944
R4811 VDD.n2018 VDD.n1422 19.3944
R4812 VDD.n2018 VDD.n1420 19.3944
R4813 VDD.n2022 VDD.n1420 19.3944
R4814 VDD.n2022 VDD.n1410 19.3944
R4815 VDD.n2034 VDD.n1410 19.3944
R4816 VDD.n2034 VDD.n1408 19.3944
R4817 VDD.n2038 VDD.n1408 19.3944
R4818 VDD.n2038 VDD.n1398 19.3944
R4819 VDD.n2050 VDD.n1398 19.3944
R4820 VDD.n2050 VDD.n1396 19.3944
R4821 VDD.n2054 VDD.n1396 19.3944
R4822 VDD.n2054 VDD.n1386 19.3944
R4823 VDD.n2066 VDD.n1386 19.3944
R4824 VDD.n2066 VDD.n1384 19.3944
R4825 VDD.n2070 VDD.n1384 19.3944
R4826 VDD.n2070 VDD.n1374 19.3944
R4827 VDD.n2082 VDD.n1374 19.3944
R4828 VDD.n2082 VDD.n1372 19.3944
R4829 VDD.n2086 VDD.n1372 19.3944
R4830 VDD.n2086 VDD.n1362 19.3944
R4831 VDD.n2098 VDD.n1362 19.3944
R4832 VDD.n2098 VDD.n1360 19.3944
R4833 VDD.n2102 VDD.n1360 19.3944
R4834 VDD.n2102 VDD.n1350 19.3944
R4835 VDD.n2114 VDD.n1350 19.3944
R4836 VDD.n2114 VDD.n1348 19.3944
R4837 VDD.n2118 VDD.n1348 19.3944
R4838 VDD.n2118 VDD.n1338 19.3944
R4839 VDD.n2130 VDD.n1338 19.3944
R4840 VDD.n2130 VDD.n1336 19.3944
R4841 VDD.n2134 VDD.n1336 19.3944
R4842 VDD.n2134 VDD.n1325 19.3944
R4843 VDD.n2148 VDD.n1325 19.3944
R4844 VDD.n2148 VDD.n1323 19.3944
R4845 VDD.n2152 VDD.n1323 19.3944
R4846 VDD.n2152 VDD.n1312 19.3944
R4847 VDD.n2515 VDD.n1312 19.3944
R4848 VDD.n2515 VDD.n1310 19.3944
R4849 VDD.n2519 VDD.n1310 19.3944
R4850 VDD.n2520 VDD.n2519 19.3944
R4851 VDD.n604 VDD.n498 19.3944
R4852 VDD.n599 VDD.n498 19.3944
R4853 VDD.n599 VDD.n598 19.3944
R4854 VDD.n598 VDD.n597 19.3944
R4855 VDD.n597 VDD.n594 19.3944
R4856 VDD.n594 VDD.n593 19.3944
R4857 VDD.n593 VDD.n590 19.3944
R4858 VDD.n590 VDD.n589 19.3944
R4859 VDD.n589 VDD.n586 19.3944
R4860 VDD.n586 VDD.n585 19.3944
R4861 VDD.n585 VDD.n582 19.3944
R4862 VDD.n582 VDD.n581 19.3944
R4863 VDD.n577 VDD.n574 19.3944
R4864 VDD.n574 VDD.n573 19.3944
R4865 VDD.n573 VDD.n570 19.3944
R4866 VDD.n570 VDD.n569 19.3944
R4867 VDD.n569 VDD.n566 19.3944
R4868 VDD.n566 VDD.n565 19.3944
R4869 VDD.n565 VDD.n562 19.3944
R4870 VDD.n562 VDD.n561 19.3944
R4871 VDD.n561 VDD.n558 19.3944
R4872 VDD.n558 VDD.n557 19.3944
R4873 VDD.n557 VDD.n554 19.3944
R4874 VDD.n554 VDD.n553 19.3944
R4875 VDD.n553 VDD.n550 19.3944
R4876 VDD.n550 VDD.n549 19.3944
R4877 VDD.n3746 VDD.n464 19.3944
R4878 VDD.n3746 VDD.n462 19.3944
R4879 VDD.n3750 VDD.n462 19.3944
R4880 VDD.n3750 VDD.n452 19.3944
R4881 VDD.n3762 VDD.n452 19.3944
R4882 VDD.n3762 VDD.n450 19.3944
R4883 VDD.n3766 VDD.n450 19.3944
R4884 VDD.n3766 VDD.n440 19.3944
R4885 VDD.n3778 VDD.n440 19.3944
R4886 VDD.n3778 VDD.n438 19.3944
R4887 VDD.n3782 VDD.n438 19.3944
R4888 VDD.n3782 VDD.n428 19.3944
R4889 VDD.n3794 VDD.n428 19.3944
R4890 VDD.n3794 VDD.n426 19.3944
R4891 VDD.n3798 VDD.n426 19.3944
R4892 VDD.n3798 VDD.n416 19.3944
R4893 VDD.n3810 VDD.n416 19.3944
R4894 VDD.n3810 VDD.n414 19.3944
R4895 VDD.n3814 VDD.n414 19.3944
R4896 VDD.n3814 VDD.n404 19.3944
R4897 VDD.n3826 VDD.n404 19.3944
R4898 VDD.n3826 VDD.n402 19.3944
R4899 VDD.n3830 VDD.n402 19.3944
R4900 VDD.n3830 VDD.n392 19.3944
R4901 VDD.n3842 VDD.n392 19.3944
R4902 VDD.n3842 VDD.n390 19.3944
R4903 VDD.n3846 VDD.n390 19.3944
R4904 VDD.n3846 VDD.n380 19.3944
R4905 VDD.n3859 VDD.n380 19.3944
R4906 VDD.n3859 VDD.n378 19.3944
R4907 VDD.n3863 VDD.n378 19.3944
R4908 VDD.n3863 VDD.n369 19.3944
R4909 VDD.n3875 VDD.n369 19.3944
R4910 VDD.n3875 VDD.n367 19.3944
R4911 VDD.n3879 VDD.n367 19.3944
R4912 VDD.n3879 VDD.n357 19.3944
R4913 VDD.n3891 VDD.n357 19.3944
R4914 VDD.n3891 VDD.n355 19.3944
R4915 VDD.n3895 VDD.n355 19.3944
R4916 VDD.n3895 VDD.n345 19.3944
R4917 VDD.n3907 VDD.n345 19.3944
R4918 VDD.n3907 VDD.n343 19.3944
R4919 VDD.n3911 VDD.n343 19.3944
R4920 VDD.n3911 VDD.n333 19.3944
R4921 VDD.n3923 VDD.n333 19.3944
R4922 VDD.n3923 VDD.n331 19.3944
R4923 VDD.n3927 VDD.n331 19.3944
R4924 VDD.n3927 VDD.n321 19.3944
R4925 VDD.n3942 VDD.n321 19.3944
R4926 VDD.n3942 VDD.n319 19.3944
R4927 VDD.n3946 VDD.n319 19.3944
R4928 VDD.n3946 VDD.n31 19.3944
R4929 VDD.n4157 VDD.n31 19.3944
R4930 VDD.n4157 VDD.n32 19.3944
R4931 VDD.n4152 VDD.n32 19.3944
R4932 VDD.n4152 VDD.n4151 19.3944
R4933 VDD.n4151 VDD.n4150 19.3944
R4934 VDD.n4150 VDD.n44 19.3944
R4935 VDD.n4144 VDD.n44 19.3944
R4936 VDD.n4144 VDD.n4143 19.3944
R4937 VDD.n4143 VDD.n4142 19.3944
R4938 VDD.n4142 VDD.n55 19.3944
R4939 VDD.n4136 VDD.n55 19.3944
R4940 VDD.n4136 VDD.n4135 19.3944
R4941 VDD.n4135 VDD.n4134 19.3944
R4942 VDD.n4134 VDD.n66 19.3944
R4943 VDD.n4128 VDD.n66 19.3944
R4944 VDD.n4128 VDD.n4127 19.3944
R4945 VDD.n4127 VDD.n4126 19.3944
R4946 VDD.n4126 VDD.n77 19.3944
R4947 VDD.n4120 VDD.n77 19.3944
R4948 VDD.n4120 VDD.n4119 19.3944
R4949 VDD.n4119 VDD.n4118 19.3944
R4950 VDD.n4118 VDD.n88 19.3944
R4951 VDD.n4112 VDD.n88 19.3944
R4952 VDD.n4112 VDD.n4111 19.3944
R4953 VDD.n4111 VDD.n4110 19.3944
R4954 VDD.n4110 VDD.n98 19.3944
R4955 VDD.n4104 VDD.n98 19.3944
R4956 VDD.n4104 VDD.n4103 19.3944
R4957 VDD.n4103 VDD.n4102 19.3944
R4958 VDD.n4102 VDD.n110 19.3944
R4959 VDD.n4096 VDD.n110 19.3944
R4960 VDD.n4096 VDD.n4095 19.3944
R4961 VDD.n4095 VDD.n4094 19.3944
R4962 VDD.n4094 VDD.n121 19.3944
R4963 VDD.n4088 VDD.n121 19.3944
R4964 VDD.n4088 VDD.n4087 19.3944
R4965 VDD.n4087 VDD.n4086 19.3944
R4966 VDD.n4086 VDD.n132 19.3944
R4967 VDD.n4080 VDD.n132 19.3944
R4968 VDD.n4080 VDD.n4079 19.3944
R4969 VDD.n4079 VDD.n4078 19.3944
R4970 VDD.n4078 VDD.n143 19.3944
R4971 VDD.n4072 VDD.n143 19.3944
R4972 VDD.n4072 VDD.n4071 19.3944
R4973 VDD.n4071 VDD.n4070 19.3944
R4974 VDD.n4070 VDD.n154 19.3944
R4975 VDD.n4064 VDD.n154 19.3944
R4976 VDD.n4064 VDD.n4063 19.3944
R4977 VDD.n4063 VDD.n4062 19.3944
R4978 VDD.n4062 VDD.n165 19.3944
R4979 VDD.n4056 VDD.n165 19.3944
R4980 VDD.n4056 VDD.n4055 19.3944
R4981 VDD.n4055 VDD.n4054 19.3944
R4982 VDD.n4054 VDD.n176 19.3944
R4983 VDD.n253 VDD.n252 19.3944
R4984 VDD.n256 VDD.n253 19.3944
R4985 VDD.n256 VDD.n203 19.3944
R4986 VDD.n262 VDD.n203 19.3944
R4987 VDD.n263 VDD.n262 19.3944
R4988 VDD.n266 VDD.n263 19.3944
R4989 VDD.n266 VDD.n201 19.3944
R4990 VDD.n272 VDD.n201 19.3944
R4991 VDD.n273 VDD.n272 19.3944
R4992 VDD.n276 VDD.n273 19.3944
R4993 VDD.n276 VDD.n199 19.3944
R4994 VDD.n282 VDD.n199 19.3944
R4995 VDD.n284 VDD.n282 19.3944
R4996 VDD.n285 VDD.n284 19.3944
R4997 VDD.n216 VDD.n213 19.3944
R4998 VDD.n222 VDD.n213 19.3944
R4999 VDD.n223 VDD.n222 19.3944
R5000 VDD.n226 VDD.n223 19.3944
R5001 VDD.n226 VDD.n211 19.3944
R5002 VDD.n232 VDD.n211 19.3944
R5003 VDD.n233 VDD.n232 19.3944
R5004 VDD.n236 VDD.n233 19.3944
R5005 VDD.n236 VDD.n209 19.3944
R5006 VDD.n242 VDD.n209 19.3944
R5007 VDD.n243 VDD.n242 19.3944
R5008 VDD.n246 VDD.n243 19.3944
R5009 VDD.n3742 VDD.n468 19.3944
R5010 VDD.n3742 VDD.n458 19.3944
R5011 VDD.n3754 VDD.n458 19.3944
R5012 VDD.n3754 VDD.n456 19.3944
R5013 VDD.n3758 VDD.n456 19.3944
R5014 VDD.n3758 VDD.n446 19.3944
R5015 VDD.n3770 VDD.n446 19.3944
R5016 VDD.n3770 VDD.n444 19.3944
R5017 VDD.n3774 VDD.n444 19.3944
R5018 VDD.n3774 VDD.n434 19.3944
R5019 VDD.n3786 VDD.n434 19.3944
R5020 VDD.n3786 VDD.n432 19.3944
R5021 VDD.n3790 VDD.n432 19.3944
R5022 VDD.n3790 VDD.n422 19.3944
R5023 VDD.n3802 VDD.n422 19.3944
R5024 VDD.n3802 VDD.n420 19.3944
R5025 VDD.n3806 VDD.n420 19.3944
R5026 VDD.n3806 VDD.n410 19.3944
R5027 VDD.n3818 VDD.n410 19.3944
R5028 VDD.n3818 VDD.n408 19.3944
R5029 VDD.n3822 VDD.n408 19.3944
R5030 VDD.n3822 VDD.n398 19.3944
R5031 VDD.n3834 VDD.n398 19.3944
R5032 VDD.n3834 VDD.n396 19.3944
R5033 VDD.n3838 VDD.n396 19.3944
R5034 VDD.n3838 VDD.n386 19.3944
R5035 VDD.n3850 VDD.n386 19.3944
R5036 VDD.n3850 VDD.n384 19.3944
R5037 VDD.n3854 VDD.n384 19.3944
R5038 VDD.n3854 VDD.n375 19.3944
R5039 VDD.n3867 VDD.n375 19.3944
R5040 VDD.n3867 VDD.n373 19.3944
R5041 VDD.n3871 VDD.n373 19.3944
R5042 VDD.n3871 VDD.n363 19.3944
R5043 VDD.n3883 VDD.n363 19.3944
R5044 VDD.n3883 VDD.n361 19.3944
R5045 VDD.n3887 VDD.n361 19.3944
R5046 VDD.n3887 VDD.n351 19.3944
R5047 VDD.n3899 VDD.n351 19.3944
R5048 VDD.n3899 VDD.n349 19.3944
R5049 VDD.n3903 VDD.n349 19.3944
R5050 VDD.n3903 VDD.n339 19.3944
R5051 VDD.n3915 VDD.n339 19.3944
R5052 VDD.n3915 VDD.n337 19.3944
R5053 VDD.n3919 VDD.n337 19.3944
R5054 VDD.n3919 VDD.n327 19.3944
R5055 VDD.n3931 VDD.n327 19.3944
R5056 VDD.n3931 VDD.n325 19.3944
R5057 VDD.n3938 VDD.n325 19.3944
R5058 VDD.n3938 VDD.n3937 19.3944
R5059 VDD.n3937 VDD.n314 19.3944
R5060 VDD.n3951 VDD.n314 19.3944
R5061 VDD.n3952 VDD.n3951 19.3944
R5062 VDD.n3953 VDD.n3952 19.3944
R5063 VDD.n3953 VDD.n312 19.3944
R5064 VDD.n3958 VDD.n312 19.3944
R5065 VDD.n3959 VDD.n3958 19.3944
R5066 VDD.n3960 VDD.n3959 19.3944
R5067 VDD.n3960 VDD.n310 19.3944
R5068 VDD.n3965 VDD.n310 19.3944
R5069 VDD.n3966 VDD.n3965 19.3944
R5070 VDD.n3967 VDD.n3966 19.3944
R5071 VDD.n3967 VDD.n308 19.3944
R5072 VDD.n3972 VDD.n308 19.3944
R5073 VDD.n3973 VDD.n3972 19.3944
R5074 VDD.n3974 VDD.n3973 19.3944
R5075 VDD.n3974 VDD.n306 19.3944
R5076 VDD.n3979 VDD.n306 19.3944
R5077 VDD.n3980 VDD.n3979 19.3944
R5078 VDD.n3981 VDD.n3980 19.3944
R5079 VDD.n3981 VDD.n304 19.3944
R5080 VDD.n3986 VDD.n304 19.3944
R5081 VDD.n3987 VDD.n3986 19.3944
R5082 VDD.n3988 VDD.n3987 19.3944
R5083 VDD.n3988 VDD.n302 19.3944
R5084 VDD.n3993 VDD.n302 19.3944
R5085 VDD.n3994 VDD.n3993 19.3944
R5086 VDD.n3995 VDD.n3994 19.3944
R5087 VDD.n3995 VDD.n300 19.3944
R5088 VDD.n4000 VDD.n300 19.3944
R5089 VDD.n4001 VDD.n4000 19.3944
R5090 VDD.n4002 VDD.n4001 19.3944
R5091 VDD.n4002 VDD.n298 19.3944
R5092 VDD.n4007 VDD.n298 19.3944
R5093 VDD.n4008 VDD.n4007 19.3944
R5094 VDD.n4009 VDD.n4008 19.3944
R5095 VDD.n4009 VDD.n296 19.3944
R5096 VDD.n4014 VDD.n296 19.3944
R5097 VDD.n4015 VDD.n4014 19.3944
R5098 VDD.n4016 VDD.n4015 19.3944
R5099 VDD.n4016 VDD.n294 19.3944
R5100 VDD.n4021 VDD.n294 19.3944
R5101 VDD.n4022 VDD.n4021 19.3944
R5102 VDD.n4023 VDD.n4022 19.3944
R5103 VDD.n4023 VDD.n292 19.3944
R5104 VDD.n4028 VDD.n292 19.3944
R5105 VDD.n4029 VDD.n4028 19.3944
R5106 VDD.n4030 VDD.n4029 19.3944
R5107 VDD.n4030 VDD.n290 19.3944
R5108 VDD.n4035 VDD.n290 19.3944
R5109 VDD.n4036 VDD.n4035 19.3944
R5110 VDD.n4037 VDD.n4036 19.3944
R5111 VDD.n4037 VDD.n288 19.3944
R5112 VDD.n4042 VDD.n288 19.3944
R5113 VDD.n4043 VDD.n4042 19.3944
R5114 VDD.n4044 VDD.n4043 19.3944
R5115 VDD.n1738 VDD.n1621 17.4637
R5116 VDD.n1738 VDD.n1615 17.4637
R5117 VDD.n1746 VDD.n1615 17.4637
R5118 VDD.n1746 VDD.n1609 17.4637
R5119 VDD.n1754 VDD.n1609 17.4637
R5120 VDD.n1762 VDD.n1603 17.4637
R5121 VDD.n1762 VDD.n1597 17.4637
R5122 VDD.n1770 VDD.n1597 17.4637
R5123 VDD.n1770 VDD.n1591 17.4637
R5124 VDD.n1778 VDD.n1591 17.4637
R5125 VDD.n1778 VDD.n1585 17.4637
R5126 VDD.n1786 VDD.n1585 17.4637
R5127 VDD.n1786 VDD.n1579 17.4637
R5128 VDD.n1794 VDD.n1579 17.4637
R5129 VDD.n1794 VDD.n1573 17.4637
R5130 VDD.n1802 VDD.n1573 17.4637
R5131 VDD.n1802 VDD.n1567 17.4637
R5132 VDD.n1810 VDD.n1567 17.4637
R5133 VDD.n1818 VDD.n1561 17.4637
R5134 VDD.n1818 VDD.n1555 17.4637
R5135 VDD.n1826 VDD.n1555 17.4637
R5136 VDD.n1826 VDD.n1549 17.4637
R5137 VDD.n1834 VDD.n1549 17.4637
R5138 VDD.n1834 VDD.n1543 17.4637
R5139 VDD.n1842 VDD.n1543 17.4637
R5140 VDD.n1842 VDD.n1536 17.4637
R5141 VDD.n1850 VDD.n1536 17.4637
R5142 VDD.n1850 VDD.n1537 17.4637
R5143 VDD.n1858 VDD.n1525 17.4637
R5144 VDD.n1866 VDD.n1525 17.4637
R5145 VDD.n1866 VDD.n1519 17.4637
R5146 VDD.n1874 VDD.n1519 17.4637
R5147 VDD.n1874 VDD.n1513 17.4637
R5148 VDD.n1882 VDD.n1513 17.4637
R5149 VDD.n1882 VDD.n1507 17.4637
R5150 VDD.n1890 VDD.n1507 17.4637
R5151 VDD.n1890 VDD.n1501 17.4637
R5152 VDD.n1898 VDD.n1501 17.4637
R5153 VDD.n1906 VDD.n1495 17.4637
R5154 VDD.n1906 VDD.n1489 17.4637
R5155 VDD.n1914 VDD.n1489 17.4637
R5156 VDD.n1914 VDD.n1483 17.4637
R5157 VDD.n1922 VDD.n1483 17.4637
R5158 VDD.n1922 VDD.n1477 17.4637
R5159 VDD.n1930 VDD.n1477 17.4637
R5160 VDD.n1930 VDD.n1471 17.4637
R5161 VDD.n1938 VDD.n1471 17.4637
R5162 VDD.n1938 VDD.n1465 17.4637
R5163 VDD.t26 VDD.n1465 17.4637
R5164 VDD.t26 VDD.n1459 17.4637
R5165 VDD.n1967 VDD.n1459 17.4637
R5166 VDD.n1967 VDD.n1453 17.4637
R5167 VDD.n1975 VDD.n1453 17.4637
R5168 VDD.n1975 VDD.n1447 17.4637
R5169 VDD.n1983 VDD.n1447 17.4637
R5170 VDD.n1983 VDD.n1441 17.4637
R5171 VDD.n1991 VDD.n1441 17.4637
R5172 VDD.n1991 VDD.n1435 17.4637
R5173 VDD.n2000 VDD.n1435 17.4637
R5174 VDD.n2000 VDD.n1999 17.4637
R5175 VDD.n2008 VDD.n1424 17.4637
R5176 VDD.n2016 VDD.n1424 17.4637
R5177 VDD.n2016 VDD.n1418 17.4637
R5178 VDD.n2024 VDD.n1418 17.4637
R5179 VDD.n2024 VDD.n1412 17.4637
R5180 VDD.n2032 VDD.n1412 17.4637
R5181 VDD.n2032 VDD.n1406 17.4637
R5182 VDD.n2040 VDD.n1406 17.4637
R5183 VDD.n2040 VDD.n1400 17.4637
R5184 VDD.n2048 VDD.n1400 17.4637
R5185 VDD.n2056 VDD.n1394 17.4637
R5186 VDD.n2056 VDD.n1388 17.4637
R5187 VDD.n2064 VDD.n1388 17.4637
R5188 VDD.n2064 VDD.n1382 17.4637
R5189 VDD.n2072 VDD.n1382 17.4637
R5190 VDD.n2072 VDD.n1376 17.4637
R5191 VDD.n2080 VDD.n1376 17.4637
R5192 VDD.n2080 VDD.n1369 17.4637
R5193 VDD.n2088 VDD.n1369 17.4637
R5194 VDD.n2088 VDD.n1370 17.4637
R5195 VDD.n2096 VDD.n1358 17.4637
R5196 VDD.n2104 VDD.n1358 17.4637
R5197 VDD.n2104 VDD.n1352 17.4637
R5198 VDD.n2112 VDD.n1352 17.4637
R5199 VDD.n2112 VDD.n1346 17.4637
R5200 VDD.n2120 VDD.n1346 17.4637
R5201 VDD.n2120 VDD.n1340 17.4637
R5202 VDD.n2128 VDD.n1340 17.4637
R5203 VDD.n2128 VDD.n1334 17.4637
R5204 VDD.n2136 VDD.n1334 17.4637
R5205 VDD.n2136 VDD.n1327 17.4637
R5206 VDD.n2146 VDD.n1327 17.4637
R5207 VDD.n2146 VDD.n2145 17.4637
R5208 VDD.n2154 VDD.n1315 17.4637
R5209 VDD.n2513 VDD.n1315 17.4637
R5210 VDD.n2513 VDD.n2512 17.4637
R5211 VDD.n2512 VDD.n1286 17.4637
R5212 VDD.n2522 VDD.n1286 17.4637
R5213 VDD.n3744 VDD.n466 17.4637
R5214 VDD.n3744 VDD.n460 17.4637
R5215 VDD.n3752 VDD.n460 17.4637
R5216 VDD.n3752 VDD.n454 17.4637
R5217 VDD.n3760 VDD.n454 17.4637
R5218 VDD.n3768 VDD.n448 17.4637
R5219 VDD.n3768 VDD.n442 17.4637
R5220 VDD.n3776 VDD.n442 17.4637
R5221 VDD.n3776 VDD.n436 17.4637
R5222 VDD.n3784 VDD.n436 17.4637
R5223 VDD.n3784 VDD.n430 17.4637
R5224 VDD.n3792 VDD.n430 17.4637
R5225 VDD.n3792 VDD.n424 17.4637
R5226 VDD.n3800 VDD.n424 17.4637
R5227 VDD.n3800 VDD.n418 17.4637
R5228 VDD.n3808 VDD.n418 17.4637
R5229 VDD.n3808 VDD.n412 17.4637
R5230 VDD.n3816 VDD.n412 17.4637
R5231 VDD.n3824 VDD.n406 17.4637
R5232 VDD.n3824 VDD.n400 17.4637
R5233 VDD.n3832 VDD.n400 17.4637
R5234 VDD.n3832 VDD.n394 17.4637
R5235 VDD.n3840 VDD.n394 17.4637
R5236 VDD.n3840 VDD.n388 17.4637
R5237 VDD.n3848 VDD.n388 17.4637
R5238 VDD.n3848 VDD.n382 17.4637
R5239 VDD.n3857 VDD.n382 17.4637
R5240 VDD.n3857 VDD.n3856 17.4637
R5241 VDD.n3865 VDD.n371 17.4637
R5242 VDD.n3873 VDD.n371 17.4637
R5243 VDD.n3873 VDD.n365 17.4637
R5244 VDD.n3881 VDD.n365 17.4637
R5245 VDD.n3881 VDD.n359 17.4637
R5246 VDD.n3889 VDD.n359 17.4637
R5247 VDD.n3889 VDD.n353 17.4637
R5248 VDD.n3897 VDD.n353 17.4637
R5249 VDD.n3897 VDD.n347 17.4637
R5250 VDD.n3905 VDD.n347 17.4637
R5251 VDD.n3913 VDD.n341 17.4637
R5252 VDD.n3913 VDD.n335 17.4637
R5253 VDD.n3921 VDD.n335 17.4637
R5254 VDD.n3921 VDD.n329 17.4637
R5255 VDD.n3929 VDD.n329 17.4637
R5256 VDD.n3929 VDD.n323 17.4637
R5257 VDD.n3940 VDD.n323 17.4637
R5258 VDD.n3940 VDD.n317 17.4637
R5259 VDD.n3948 VDD.n317 17.4637
R5260 VDD.n3948 VDD.n35 17.4637
R5261 VDD.t23 VDD.n35 17.4637
R5262 VDD.t23 VDD.n4155 17.4637
R5263 VDD.n4155 VDD.n4154 17.4637
R5264 VDD.n4154 VDD.n39 17.4637
R5265 VDD.n4148 VDD.n39 17.4637
R5266 VDD.n4148 VDD.n4147 17.4637
R5267 VDD.n4147 VDD.n4146 17.4637
R5268 VDD.n4146 VDD.n49 17.4637
R5269 VDD.n4140 VDD.n49 17.4637
R5270 VDD.n4140 VDD.n4139 17.4637
R5271 VDD.n4139 VDD.n4138 17.4637
R5272 VDD.n4138 VDD.n60 17.4637
R5273 VDD.n4132 VDD.n4131 17.4637
R5274 VDD.n4131 VDD.n4130 17.4637
R5275 VDD.n4130 VDD.n71 17.4637
R5276 VDD.n4124 VDD.n71 17.4637
R5277 VDD.n4124 VDD.n4123 17.4637
R5278 VDD.n4123 VDD.n4122 17.4637
R5279 VDD.n4122 VDD.n82 17.4637
R5280 VDD.n4116 VDD.n82 17.4637
R5281 VDD.n4116 VDD.n4115 17.4637
R5282 VDD.n4115 VDD.n4114 17.4637
R5283 VDD.n4108 VDD.n100 17.4637
R5284 VDD.n4108 VDD.n4107 17.4637
R5285 VDD.n4107 VDD.n4106 17.4637
R5286 VDD.n4106 VDD.n104 17.4637
R5287 VDD.n4100 VDD.n104 17.4637
R5288 VDD.n4100 VDD.n4099 17.4637
R5289 VDD.n4099 VDD.n4098 17.4637
R5290 VDD.n4098 VDD.n115 17.4637
R5291 VDD.n4092 VDD.n115 17.4637
R5292 VDD.n4092 VDD.n4091 17.4637
R5293 VDD.n4090 VDD.n126 17.4637
R5294 VDD.n4084 VDD.n126 17.4637
R5295 VDD.n4084 VDD.n4083 17.4637
R5296 VDD.n4083 VDD.n4082 17.4637
R5297 VDD.n4082 VDD.n137 17.4637
R5298 VDD.n4076 VDD.n137 17.4637
R5299 VDD.n4076 VDD.n4075 17.4637
R5300 VDD.n4075 VDD.n4074 17.4637
R5301 VDD.n4074 VDD.n148 17.4637
R5302 VDD.n4068 VDD.n148 17.4637
R5303 VDD.n4068 VDD.n4067 17.4637
R5304 VDD.n4067 VDD.n4066 17.4637
R5305 VDD.n4066 VDD.n159 17.4637
R5306 VDD.n4060 VDD.n4059 17.4637
R5307 VDD.n4059 VDD.n4058 17.4637
R5308 VDD.n4058 VDD.n170 17.4637
R5309 VDD.n4052 VDD.n170 17.4637
R5310 VDD.n4052 VDD.n4051 17.4637
R5311 VDD.n2550 VDD.n2549 15.9035
R5312 VDD.n1710 VDD.n1706 15.9035
R5313 VDD.n578 VDD.n577 15.9035
R5314 VDD.n252 VDD.n207 15.9035
R5315 VDD.n1754 VDD.t86 15.0189
R5316 VDD.n2154 VDD.t82 15.0189
R5317 VDD.n3760 VDD.t94 15.0189
R5318 VDD.n4060 VDD.t104 15.0189
R5319 VDD.n1898 VDD.t67 13.2726
R5320 VDD.n2008 VDD.t52 13.2726
R5321 VDD.n3905 VDD.t47 13.2726
R5322 VDD.n4132 VDD.t17 13.2726
R5323 VDD.t54 VDD.n1561 12.574
R5324 VDD.n1370 VDD.t69 12.574
R5325 VDD.t37 VDD.n406 12.574
R5326 VDD.n4091 VDD.t7 12.574
R5327 VDD.n2595 VDD.n1214 11.8755
R5328 VDD.n2595 VDD.n1208 11.8755
R5329 VDD.n2601 VDD.n1208 11.8755
R5330 VDD.n2601 VDD.n1202 11.8755
R5331 VDD.n2607 VDD.n1202 11.8755
R5332 VDD.n2607 VDD.n1196 11.8755
R5333 VDD.n2613 VDD.n1196 11.8755
R5334 VDD.n2619 VDD.n1185 11.8755
R5335 VDD.n2625 VDD.n1185 11.8755
R5336 VDD.n2625 VDD.n1179 11.8755
R5337 VDD.n2631 VDD.n1179 11.8755
R5338 VDD.n2631 VDD.n1173 11.8755
R5339 VDD.n2637 VDD.n1173 11.8755
R5340 VDD.n2637 VDD.n1167 11.8755
R5341 VDD.n2643 VDD.n1167 11.8755
R5342 VDD.n2643 VDD.n1161 11.8755
R5343 VDD.n2649 VDD.n1161 11.8755
R5344 VDD.n2649 VDD.n1155 11.8755
R5345 VDD.n2655 VDD.n1155 11.8755
R5346 VDD.n2661 VDD.n1149 11.8755
R5347 VDD.n2667 VDD.n1143 11.8755
R5348 VDD.n2667 VDD.n1137 11.8755
R5349 VDD.n2673 VDD.n1137 11.8755
R5350 VDD.n2673 VDD.n1131 11.8755
R5351 VDD.n2679 VDD.n1131 11.8755
R5352 VDD.n2679 VDD.n1125 11.8755
R5353 VDD.n2685 VDD.n1125 11.8755
R5354 VDD.n2685 VDD.n1119 11.8755
R5355 VDD.n2691 VDD.n1119 11.8755
R5356 VDD.n2697 VDD.n1113 11.8755
R5357 VDD.n2703 VDD.n1107 11.8755
R5358 VDD.n2703 VDD.n1101 11.8755
R5359 VDD.n2709 VDD.n1101 11.8755
R5360 VDD.n2709 VDD.n1095 11.8755
R5361 VDD.n2715 VDD.n1095 11.8755
R5362 VDD.n2715 VDD.n1089 11.8755
R5363 VDD.n2721 VDD.n1089 11.8755
R5364 VDD.n2721 VDD.n1083 11.8755
R5365 VDD.n2727 VDD.n1083 11.8755
R5366 VDD.n2727 VDD.n1077 11.8755
R5367 VDD.n2733 VDD.n1077 11.8755
R5368 VDD.n2733 VDD.t25 11.8755
R5369 VDD.n2739 VDD.t25 11.8755
R5370 VDD.n2739 VDD.n1065 11.8755
R5371 VDD.n2745 VDD.n1065 11.8755
R5372 VDD.n2745 VDD.n1068 11.8755
R5373 VDD.n2751 VDD.n1054 11.8755
R5374 VDD.n2757 VDD.n1054 11.8755
R5375 VDD.n2757 VDD.n1048 11.8755
R5376 VDD.n2763 VDD.n1048 11.8755
R5377 VDD.n2763 VDD.n1041 11.8755
R5378 VDD.n2769 VDD.n1041 11.8755
R5379 VDD.n2769 VDD.n1044 11.8755
R5380 VDD.n2775 VDD.n1029 11.8755
R5381 VDD.n2781 VDD.n1029 11.8755
R5382 VDD.n2781 VDD.n1032 11.8755
R5383 VDD.n2787 VDD.n1018 11.8755
R5384 VDD.n2793 VDD.n1018 11.8755
R5385 VDD.n2793 VDD.n1012 11.8755
R5386 VDD.n2799 VDD.n1012 11.8755
R5387 VDD.n2799 VDD.n1005 11.8755
R5388 VDD.n2805 VDD.n1005 11.8755
R5389 VDD.n2805 VDD.n1008 11.8755
R5390 VDD.n2811 VDD.n994 11.8755
R5391 VDD.n2817 VDD.n994 11.8755
R5392 VDD.n2817 VDD.n988 11.8755
R5393 VDD.n2823 VDD.n988 11.8755
R5394 VDD.n2829 VDD.n982 11.8755
R5395 VDD.n2829 VDD.n976 11.8755
R5396 VDD.n2835 VDD.n976 11.8755
R5397 VDD.n2835 VDD.n970 11.8755
R5398 VDD.n2841 VDD.n970 11.8755
R5399 VDD.n2841 VDD.n964 11.8755
R5400 VDD.n2847 VDD.n964 11.8755
R5401 VDD.n2847 VDD.n957 11.8755
R5402 VDD.n2853 VDD.n957 11.8755
R5403 VDD.n2853 VDD.n960 11.8755
R5404 VDD.n2911 VDD.n945 11.8755
R5405 VDD.n2911 VDD.n939 11.8755
R5406 VDD.n2917 VDD.n939 11.8755
R5407 VDD.n2917 VDD.n929 11.8755
R5408 VDD.n2968 VDD.n929 11.8755
R5409 VDD.n2968 VDD.n904 11.8755
R5410 VDD.n3295 VDD.n898 11.8755
R5411 VDD.n3301 VDD.n898 11.8755
R5412 VDD.n3301 VDD.n892 11.8755
R5413 VDD.n3307 VDD.n892 11.8755
R5414 VDD.n3307 VDD.n886 11.8755
R5415 VDD.n3313 VDD.n886 11.8755
R5416 VDD.n3319 VDD.n875 11.8755
R5417 VDD.n3325 VDD.n875 11.8755
R5418 VDD.n3325 VDD.n869 11.8755
R5419 VDD.n3331 VDD.n869 11.8755
R5420 VDD.n3331 VDD.n863 11.8755
R5421 VDD.n3337 VDD.n863 11.8755
R5422 VDD.n3337 VDD.n857 11.8755
R5423 VDD.n3343 VDD.n857 11.8755
R5424 VDD.n3343 VDD.n851 11.8755
R5425 VDD.n3349 VDD.n851 11.8755
R5426 VDD.n3355 VDD.n845 11.8755
R5427 VDD.n3355 VDD.n838 11.8755
R5428 VDD.n3361 VDD.n838 11.8755
R5429 VDD.n3361 VDD.n841 11.8755
R5430 VDD.n3367 VDD.n827 11.8755
R5431 VDD.n3373 VDD.n827 11.8755
R5432 VDD.n3373 VDD.n821 11.8755
R5433 VDD.n3379 VDD.n821 11.8755
R5434 VDD.n3379 VDD.n814 11.8755
R5435 VDD.n3385 VDD.n814 11.8755
R5436 VDD.n3385 VDD.n817 11.8755
R5437 VDD.n3391 VDD.n802 11.8755
R5438 VDD.n3397 VDD.n802 11.8755
R5439 VDD.n3397 VDD.n805 11.8755
R5440 VDD.n3403 VDD.n791 11.8755
R5441 VDD.n3409 VDD.n791 11.8755
R5442 VDD.n3409 VDD.n785 11.8755
R5443 VDD.n3415 VDD.n785 11.8755
R5444 VDD.n3415 VDD.n778 11.8755
R5445 VDD.n3421 VDD.n778 11.8755
R5446 VDD.n3421 VDD.n781 11.8755
R5447 VDD.n3432 VDD.n766 11.8755
R5448 VDD.n3438 VDD.n766 11.8755
R5449 VDD.n3438 VDD.n759 11.8755
R5450 VDD.t16 VDD.n759 11.8755
R5451 VDD.t16 VDD.n753 11.8755
R5452 VDD.n3515 VDD.n753 11.8755
R5453 VDD.n3515 VDD.n747 11.8755
R5454 VDD.n3521 VDD.n747 11.8755
R5455 VDD.n3521 VDD.n741 11.8755
R5456 VDD.n3527 VDD.n741 11.8755
R5457 VDD.n3527 VDD.n735 11.8755
R5458 VDD.n3533 VDD.n735 11.8755
R5459 VDD.n3533 VDD.n729 11.8755
R5460 VDD.n3539 VDD.n729 11.8755
R5461 VDD.n3539 VDD.n723 11.8755
R5462 VDD.n3545 VDD.n723 11.8755
R5463 VDD.n3551 VDD.n717 11.8755
R5464 VDD.n3557 VDD.n711 11.8755
R5465 VDD.n3557 VDD.n705 11.8755
R5466 VDD.n3563 VDD.n705 11.8755
R5467 VDD.n3563 VDD.n699 11.8755
R5468 VDD.n3569 VDD.n699 11.8755
R5469 VDD.n3569 VDD.n693 11.8755
R5470 VDD.n3575 VDD.n693 11.8755
R5471 VDD.n3575 VDD.n687 11.8755
R5472 VDD.n3581 VDD.n687 11.8755
R5473 VDD.n3587 VDD.n681 11.8755
R5474 VDD.n3593 VDD.n675 11.8755
R5475 VDD.n3593 VDD.n669 11.8755
R5476 VDD.n3599 VDD.n669 11.8755
R5477 VDD.n3599 VDD.n663 11.8755
R5478 VDD.n3605 VDD.n663 11.8755
R5479 VDD.n3605 VDD.n657 11.8755
R5480 VDD.n3611 VDD.n657 11.8755
R5481 VDD.n3611 VDD.n651 11.8755
R5482 VDD.n3617 VDD.n651 11.8755
R5483 VDD.n3617 VDD.n644 11.8755
R5484 VDD.n3623 VDD.n644 11.8755
R5485 VDD.n3623 VDD.n647 11.8755
R5486 VDD.n3635 VDD.n633 11.8755
R5487 VDD.n3635 VDD.n626 11.8755
R5488 VDD.n3669 VDD.n626 11.8755
R5489 VDD.n3669 VDD.n620 11.8755
R5490 VDD.n3675 VDD.n620 11.8755
R5491 VDD.n3675 VDD.n485 11.8755
R5492 VDD.n3718 VDD.n485 11.8755
R5493 VDD.n2572 VDD.n2571 11.5727
R5494 VDD.n607 VDD.n606 11.5717
R5495 VDD.t130 VDD.n1149 10.6531
R5496 VDD.n3587 VDD.t59 10.6531
R5497 VDD.n3174 VDD.n3172 10.6151
R5498 VDD.n3175 VDD.n3174 10.6151
R5499 VDD.n3177 VDD.n3175 10.6151
R5500 VDD.n3178 VDD.n3177 10.6151
R5501 VDD.n3180 VDD.n3178 10.6151
R5502 VDD.n3181 VDD.n3180 10.6151
R5503 VDD.n3237 VDD.n3181 10.6151
R5504 VDD.n3237 VDD.n3236 10.6151
R5505 VDD.n3236 VDD.n3235 10.6151
R5506 VDD.n3235 VDD.n3233 10.6151
R5507 VDD.n3233 VDD.n3232 10.6151
R5508 VDD.n3232 VDD.n3230 10.6151
R5509 VDD.n3230 VDD.n3229 10.6151
R5510 VDD.n3229 VDD.n3227 10.6151
R5511 VDD.n3227 VDD.n3226 10.6151
R5512 VDD.n3226 VDD.n3224 10.6151
R5513 VDD.n3224 VDD.n3223 10.6151
R5514 VDD.n3223 VDD.n3221 10.6151
R5515 VDD.n3221 VDD.n3220 10.6151
R5516 VDD.n3220 VDD.n3218 10.6151
R5517 VDD.n3218 VDD.n3217 10.6151
R5518 VDD.n3217 VDD.n3215 10.6151
R5519 VDD.n3215 VDD.n3214 10.6151
R5520 VDD.n3214 VDD.n3212 10.6151
R5521 VDD.n3212 VDD.n3211 10.6151
R5522 VDD.n3211 VDD.n3209 10.6151
R5523 VDD.n3209 VDD.n3208 10.6151
R5524 VDD.n3208 VDD.n3206 10.6151
R5525 VDD.n3206 VDD.n3205 10.6151
R5526 VDD.n3205 VDD.n3203 10.6151
R5527 VDD.n3203 VDD.n3202 10.6151
R5528 VDD.n3202 VDD.n3200 10.6151
R5529 VDD.n3200 VDD.n3199 10.6151
R5530 VDD.n3199 VDD.n3197 10.6151
R5531 VDD.n3197 VDD.n3196 10.6151
R5532 VDD.n3196 VDD.n3194 10.6151
R5533 VDD.n3194 VDD.n3193 10.6151
R5534 VDD.n3193 VDD.n3191 10.6151
R5535 VDD.n3191 VDD.n3190 10.6151
R5536 VDD.n3190 VDD.n3188 10.6151
R5537 VDD.n3188 VDD.n3187 10.6151
R5538 VDD.n3187 VDD.n3185 10.6151
R5539 VDD.n3185 VDD.n3184 10.6151
R5540 VDD.n3184 VDD.n3182 10.6151
R5541 VDD.n3182 VDD.n764 10.6151
R5542 VDD.n3440 VDD.n764 10.6151
R5543 VDD.n3441 VDD.n3440 10.6151
R5544 VDD.n3508 VDD.n3441 10.6151
R5545 VDD.n3508 VDD.n3507 10.6151
R5546 VDD.n3507 VDD.n3506 10.6151
R5547 VDD.n3506 VDD.n3505 10.6151
R5548 VDD.n3505 VDD.n3503 10.6151
R5549 VDD.n3503 VDD.n3502 10.6151
R5550 VDD.n3502 VDD.n3500 10.6151
R5551 VDD.n3500 VDD.n3499 10.6151
R5552 VDD.n3499 VDD.n3497 10.6151
R5553 VDD.n3497 VDD.n3496 10.6151
R5554 VDD.n3496 VDD.n3494 10.6151
R5555 VDD.n3494 VDD.n3493 10.6151
R5556 VDD.n3493 VDD.n3491 10.6151
R5557 VDD.n3491 VDD.n3490 10.6151
R5558 VDD.n3490 VDD.n3488 10.6151
R5559 VDD.n3488 VDD.n3487 10.6151
R5560 VDD.n3487 VDD.n3485 10.6151
R5561 VDD.n3485 VDD.n3484 10.6151
R5562 VDD.n3484 VDD.n3482 10.6151
R5563 VDD.n3482 VDD.n3481 10.6151
R5564 VDD.n3481 VDD.n3479 10.6151
R5565 VDD.n3479 VDD.n3478 10.6151
R5566 VDD.n3478 VDD.n3476 10.6151
R5567 VDD.n3476 VDD.n3475 10.6151
R5568 VDD.n3475 VDD.n3473 10.6151
R5569 VDD.n3473 VDD.n3472 10.6151
R5570 VDD.n3472 VDD.n3470 10.6151
R5571 VDD.n3470 VDD.n3469 10.6151
R5572 VDD.n3469 VDD.n3467 10.6151
R5573 VDD.n3467 VDD.n3466 10.6151
R5574 VDD.n3466 VDD.n3464 10.6151
R5575 VDD.n3464 VDD.n3463 10.6151
R5576 VDD.n3463 VDD.n3461 10.6151
R5577 VDD.n3461 VDD.n3460 10.6151
R5578 VDD.n3460 VDD.n3458 10.6151
R5579 VDD.n3458 VDD.n3457 10.6151
R5580 VDD.n3457 VDD.n3455 10.6151
R5581 VDD.n3455 VDD.n3454 10.6151
R5582 VDD.n3454 VDD.n3452 10.6151
R5583 VDD.n3452 VDD.n3451 10.6151
R5584 VDD.n3451 VDD.n3449 10.6151
R5585 VDD.n3449 VDD.n3448 10.6151
R5586 VDD.n3448 VDD.n3446 10.6151
R5587 VDD.n3446 VDD.n3445 10.6151
R5588 VDD.n3445 VDD.n3443 10.6151
R5589 VDD.n3443 VDD.n3442 10.6151
R5590 VDD.n3442 VDD.n618 10.6151
R5591 VDD.n3678 VDD.n618 10.6151
R5592 VDD.n3679 VDD.n3678 10.6151
R5593 VDD.n3133 VDD.n902 10.6151
R5594 VDD.n3133 VDD.n3132 10.6151
R5595 VDD.n3139 VDD.n3132 10.6151
R5596 VDD.n3140 VDD.n3139 10.6151
R5597 VDD.n3141 VDD.n3140 10.6151
R5598 VDD.n3141 VDD.n3130 10.6151
R5599 VDD.n3147 VDD.n3130 10.6151
R5600 VDD.n3148 VDD.n3147 10.6151
R5601 VDD.n3149 VDD.n3148 10.6151
R5602 VDD.n3149 VDD.n3128 10.6151
R5603 VDD.n3155 VDD.n3128 10.6151
R5604 VDD.n3156 VDD.n3155 10.6151
R5605 VDD.n3157 VDD.n3156 10.6151
R5606 VDD.n3157 VDD.n3126 10.6151
R5607 VDD.n3163 VDD.n3126 10.6151
R5608 VDD.n3164 VDD.n3163 10.6151
R5609 VDD.n3166 VDD.n3122 10.6151
R5610 VDD.n3171 VDD.n3122 10.6151
R5611 VDD.n3298 VDD.n3297 10.6151
R5612 VDD.n3299 VDD.n3298 10.6151
R5613 VDD.n3299 VDD.n890 10.6151
R5614 VDD.n3309 VDD.n890 10.6151
R5615 VDD.n3310 VDD.n3309 10.6151
R5616 VDD.n3311 VDD.n3310 10.6151
R5617 VDD.n3311 VDD.n879 10.6151
R5618 VDD.n3321 VDD.n879 10.6151
R5619 VDD.n3322 VDD.n3321 10.6151
R5620 VDD.n3323 VDD.n3322 10.6151
R5621 VDD.n3323 VDD.n867 10.6151
R5622 VDD.n3333 VDD.n867 10.6151
R5623 VDD.n3334 VDD.n3333 10.6151
R5624 VDD.n3335 VDD.n3334 10.6151
R5625 VDD.n3335 VDD.n855 10.6151
R5626 VDD.n3345 VDD.n855 10.6151
R5627 VDD.n3346 VDD.n3345 10.6151
R5628 VDD.n3347 VDD.n3346 10.6151
R5629 VDD.n3347 VDD.n843 10.6151
R5630 VDD.n3357 VDD.n843 10.6151
R5631 VDD.n3358 VDD.n3357 10.6151
R5632 VDD.n3359 VDD.n3358 10.6151
R5633 VDD.n3359 VDD.n831 10.6151
R5634 VDD.n3369 VDD.n831 10.6151
R5635 VDD.n3370 VDD.n3369 10.6151
R5636 VDD.n3371 VDD.n3370 10.6151
R5637 VDD.n3371 VDD.n819 10.6151
R5638 VDD.n3381 VDD.n819 10.6151
R5639 VDD.n3382 VDD.n3381 10.6151
R5640 VDD.n3383 VDD.n3382 10.6151
R5641 VDD.n3383 VDD.n807 10.6151
R5642 VDD.n3393 VDD.n807 10.6151
R5643 VDD.n3394 VDD.n3393 10.6151
R5644 VDD.n3395 VDD.n3394 10.6151
R5645 VDD.n3395 VDD.n795 10.6151
R5646 VDD.n3405 VDD.n795 10.6151
R5647 VDD.n3406 VDD.n3405 10.6151
R5648 VDD.n3407 VDD.n3406 10.6151
R5649 VDD.n3407 VDD.n783 10.6151
R5650 VDD.n3417 VDD.n783 10.6151
R5651 VDD.n3418 VDD.n3417 10.6151
R5652 VDD.n3419 VDD.n3418 10.6151
R5653 VDD.n3419 VDD.n770 10.6151
R5654 VDD.n3434 VDD.n770 10.6151
R5655 VDD.n3435 VDD.n3434 10.6151
R5656 VDD.n3436 VDD.n3435 10.6151
R5657 VDD.n3436 VDD.n757 10.6151
R5658 VDD.n3511 VDD.n757 10.6151
R5659 VDD.n3512 VDD.n3511 10.6151
R5660 VDD.n3513 VDD.n3512 10.6151
R5661 VDD.n3513 VDD.n745 10.6151
R5662 VDD.n3523 VDD.n745 10.6151
R5663 VDD.n3524 VDD.n3523 10.6151
R5664 VDD.n3525 VDD.n3524 10.6151
R5665 VDD.n3525 VDD.n733 10.6151
R5666 VDD.n3535 VDD.n733 10.6151
R5667 VDD.n3536 VDD.n3535 10.6151
R5668 VDD.n3537 VDD.n3536 10.6151
R5669 VDD.n3537 VDD.n721 10.6151
R5670 VDD.n3547 VDD.n721 10.6151
R5671 VDD.n3548 VDD.n3547 10.6151
R5672 VDD.n3549 VDD.n3548 10.6151
R5673 VDD.n3549 VDD.n709 10.6151
R5674 VDD.n3559 VDD.n709 10.6151
R5675 VDD.n3560 VDD.n3559 10.6151
R5676 VDD.n3561 VDD.n3560 10.6151
R5677 VDD.n3561 VDD.n697 10.6151
R5678 VDD.n3571 VDD.n697 10.6151
R5679 VDD.n3572 VDD.n3571 10.6151
R5680 VDD.n3573 VDD.n3572 10.6151
R5681 VDD.n3573 VDD.n685 10.6151
R5682 VDD.n3583 VDD.n685 10.6151
R5683 VDD.n3584 VDD.n3583 10.6151
R5684 VDD.n3585 VDD.n3584 10.6151
R5685 VDD.n3585 VDD.n673 10.6151
R5686 VDD.n3595 VDD.n673 10.6151
R5687 VDD.n3596 VDD.n3595 10.6151
R5688 VDD.n3597 VDD.n3596 10.6151
R5689 VDD.n3597 VDD.n661 10.6151
R5690 VDD.n3607 VDD.n661 10.6151
R5691 VDD.n3608 VDD.n3607 10.6151
R5692 VDD.n3609 VDD.n3608 10.6151
R5693 VDD.n3609 VDD.n649 10.6151
R5694 VDD.n3619 VDD.n649 10.6151
R5695 VDD.n3620 VDD.n3619 10.6151
R5696 VDD.n3621 VDD.n3620 10.6151
R5697 VDD.n3621 VDD.n637 10.6151
R5698 VDD.n3631 VDD.n637 10.6151
R5699 VDD.n3632 VDD.n3631 10.6151
R5700 VDD.n3633 VDD.n3632 10.6151
R5701 VDD.n3633 VDD.n624 10.6151
R5702 VDD.n3671 VDD.n624 10.6151
R5703 VDD.n3672 VDD.n3671 10.6151
R5704 VDD.n3673 VDD.n3672 10.6151
R5705 VDD.n3673 VDD.n490 10.6151
R5706 VDD.n3716 VDD.n490 10.6151
R5707 VDD.n3715 VDD.n3714 10.6151
R5708 VDD.n3714 VDD.n491 10.6151
R5709 VDD.n3709 VDD.n491 10.6151
R5710 VDD.n3709 VDD.n3708 10.6151
R5711 VDD.n3708 VDD.n3707 10.6151
R5712 VDD.n3707 VDD.n494 10.6151
R5713 VDD.n3702 VDD.n494 10.6151
R5714 VDD.n3702 VDD.n3701 10.6151
R5715 VDD.n3701 VDD.n3700 10.6151
R5716 VDD.n3695 VDD.n609 10.6151
R5717 VDD.n3695 VDD.n3694 10.6151
R5718 VDD.n3694 VDD.n3693 10.6151
R5719 VDD.n3693 VDD.n611 10.6151
R5720 VDD.n3688 VDD.n611 10.6151
R5721 VDD.n3688 VDD.n3687 10.6151
R5722 VDD.n3685 VDD.n616 10.6151
R5723 VDD.n3680 VDD.n616 10.6151
R5724 VDD.n3661 VDD.n3639 10.6151
R5725 VDD.n3640 VDD.n3639 10.6151
R5726 VDD.n3654 VDD.n3640 10.6151
R5727 VDD.n3654 VDD.n3653 10.6151
R5728 VDD.n3653 VDD.n3652 10.6151
R5729 VDD.n3652 VDD.n3642 10.6151
R5730 VDD.n3647 VDD.n3642 10.6151
R5731 VDD.n3647 VDD.n3646 10.6151
R5732 VDD.n3646 VDD.n470 10.6151
R5733 VDD.n3737 VDD.n471 10.6151
R5734 VDD.n474 VDD.n471 10.6151
R5735 VDD.n3730 VDD.n474 10.6151
R5736 VDD.n3730 VDD.n3729 10.6151
R5737 VDD.n3729 VDD.n3728 10.6151
R5738 VDD.n3728 VDD.n476 10.6151
R5739 VDD.n3723 VDD.n3722 10.6151
R5740 VDD.n3722 VDD.n3721 10.6151
R5741 VDD.n3251 VDD.n3250 10.6151
R5742 VDD.n3250 VDD.n3248 10.6151
R5743 VDD.n3248 VDD.n3247 10.6151
R5744 VDD.n3247 VDD.n3245 10.6151
R5745 VDD.n3245 VDD.n3244 10.6151
R5746 VDD.n3244 VDD.n3242 10.6151
R5747 VDD.n3242 VDD.n3241 10.6151
R5748 VDD.n3241 VDD.n3121 10.6151
R5749 VDD.n3121 VDD.n3120 10.6151
R5750 VDD.n3120 VDD.n3118 10.6151
R5751 VDD.n3118 VDD.n3117 10.6151
R5752 VDD.n3117 VDD.n3115 10.6151
R5753 VDD.n3115 VDD.n3114 10.6151
R5754 VDD.n3114 VDD.n3112 10.6151
R5755 VDD.n3112 VDD.n3111 10.6151
R5756 VDD.n3111 VDD.n3109 10.6151
R5757 VDD.n3109 VDD.n3108 10.6151
R5758 VDD.n3108 VDD.n3106 10.6151
R5759 VDD.n3106 VDD.n3105 10.6151
R5760 VDD.n3105 VDD.n3103 10.6151
R5761 VDD.n3103 VDD.n3102 10.6151
R5762 VDD.n3102 VDD.n3100 10.6151
R5763 VDD.n3100 VDD.n3099 10.6151
R5764 VDD.n3099 VDD.n3097 10.6151
R5765 VDD.n3097 VDD.n3096 10.6151
R5766 VDD.n3096 VDD.n3094 10.6151
R5767 VDD.n3094 VDD.n3093 10.6151
R5768 VDD.n3093 VDD.n3091 10.6151
R5769 VDD.n3091 VDD.n3090 10.6151
R5770 VDD.n3090 VDD.n3088 10.6151
R5771 VDD.n3088 VDD.n3087 10.6151
R5772 VDD.n3087 VDD.n3085 10.6151
R5773 VDD.n3085 VDD.n3084 10.6151
R5774 VDD.n3084 VDD.n3082 10.6151
R5775 VDD.n3082 VDD.n3081 10.6151
R5776 VDD.n3081 VDD.n3079 10.6151
R5777 VDD.n3079 VDD.n3078 10.6151
R5778 VDD.n3078 VDD.n3076 10.6151
R5779 VDD.n3076 VDD.n3075 10.6151
R5780 VDD.n3075 VDD.n3073 10.6151
R5781 VDD.n3073 VDD.n3072 10.6151
R5782 VDD.n3072 VDD.n3070 10.6151
R5783 VDD.n3070 VDD.n3069 10.6151
R5784 VDD.n3069 VDD.n3067 10.6151
R5785 VDD.n3067 VDD.n3066 10.6151
R5786 VDD.n3066 VDD.n3064 10.6151
R5787 VDD.n3064 VDD.n3063 10.6151
R5788 VDD.n3063 VDD.n3061 10.6151
R5789 VDD.n3061 VDD.n3060 10.6151
R5790 VDD.n3060 VDD.n3058 10.6151
R5791 VDD.n3058 VDD.n3057 10.6151
R5792 VDD.n3057 VDD.n3055 10.6151
R5793 VDD.n3055 VDD.n3054 10.6151
R5794 VDD.n3054 VDD.n3052 10.6151
R5795 VDD.n3052 VDD.n3051 10.6151
R5796 VDD.n3051 VDD.n3049 10.6151
R5797 VDD.n3049 VDD.n3048 10.6151
R5798 VDD.n3048 VDD.n3046 10.6151
R5799 VDD.n3046 VDD.n3045 10.6151
R5800 VDD.n3045 VDD.n3043 10.6151
R5801 VDD.n3043 VDD.n3042 10.6151
R5802 VDD.n3042 VDD.n3040 10.6151
R5803 VDD.n3040 VDD.n3039 10.6151
R5804 VDD.n3039 VDD.n3037 10.6151
R5805 VDD.n3037 VDD.n3036 10.6151
R5806 VDD.n3036 VDD.n3034 10.6151
R5807 VDD.n3034 VDD.n3033 10.6151
R5808 VDD.n3033 VDD.n3031 10.6151
R5809 VDD.n3031 VDD.n3030 10.6151
R5810 VDD.n3030 VDD.n3028 10.6151
R5811 VDD.n3028 VDD.n3027 10.6151
R5812 VDD.n3027 VDD.n3025 10.6151
R5813 VDD.n3025 VDD.n3024 10.6151
R5814 VDD.n3024 VDD.n3022 10.6151
R5815 VDD.n3022 VDD.n3021 10.6151
R5816 VDD.n3021 VDD.n3019 10.6151
R5817 VDD.n3019 VDD.n3018 10.6151
R5818 VDD.n3018 VDD.n3016 10.6151
R5819 VDD.n3016 VDD.n3015 10.6151
R5820 VDD.n3015 VDD.n3013 10.6151
R5821 VDD.n3013 VDD.n3012 10.6151
R5822 VDD.n3012 VDD.n3010 10.6151
R5823 VDD.n3010 VDD.n3009 10.6151
R5824 VDD.n3009 VDD.n3007 10.6151
R5825 VDD.n3007 VDD.n3006 10.6151
R5826 VDD.n3006 VDD.n3004 10.6151
R5827 VDD.n3004 VDD.n3003 10.6151
R5828 VDD.n3003 VDD.n3001 10.6151
R5829 VDD.n3001 VDD.n3000 10.6151
R5830 VDD.n3000 VDD.n2998 10.6151
R5831 VDD.n2998 VDD.n2997 10.6151
R5832 VDD.n2997 VDD.n2995 10.6151
R5833 VDD.n2995 VDD.n2994 10.6151
R5834 VDD.n2994 VDD.n2992 10.6151
R5835 VDD.n2992 VDD.n2991 10.6151
R5836 VDD.n2991 VDD.n482 10.6151
R5837 VDD.n3292 VDD.n3291 10.6151
R5838 VDD.n3291 VDD.n2980 10.6151
R5839 VDD.n3285 VDD.n2980 10.6151
R5840 VDD.n3285 VDD.n3284 10.6151
R5841 VDD.n3284 VDD.n3283 10.6151
R5842 VDD.n3283 VDD.n2982 10.6151
R5843 VDD.n3277 VDD.n2982 10.6151
R5844 VDD.n3277 VDD.n3276 10.6151
R5845 VDD.n3276 VDD.n3275 10.6151
R5846 VDD.n3275 VDD.n2984 10.6151
R5847 VDD.n3269 VDD.n2984 10.6151
R5848 VDD.n3269 VDD.n3268 10.6151
R5849 VDD.n3268 VDD.n3267 10.6151
R5850 VDD.n3267 VDD.n2986 10.6151
R5851 VDD.n3261 VDD.n2986 10.6151
R5852 VDD.n3261 VDD.n3260 10.6151
R5853 VDD.n3258 VDD.n2990 10.6151
R5854 VDD.n3252 VDD.n2990 10.6151
R5855 VDD.n3293 VDD.n896 10.6151
R5856 VDD.n3303 VDD.n896 10.6151
R5857 VDD.n3304 VDD.n3303 10.6151
R5858 VDD.n3305 VDD.n3304 10.6151
R5859 VDD.n3305 VDD.n884 10.6151
R5860 VDD.n3315 VDD.n884 10.6151
R5861 VDD.n3316 VDD.n3315 10.6151
R5862 VDD.n3317 VDD.n3316 10.6151
R5863 VDD.n3317 VDD.n873 10.6151
R5864 VDD.n3327 VDD.n873 10.6151
R5865 VDD.n3328 VDD.n3327 10.6151
R5866 VDD.n3329 VDD.n3328 10.6151
R5867 VDD.n3329 VDD.n861 10.6151
R5868 VDD.n3339 VDD.n861 10.6151
R5869 VDD.n3340 VDD.n3339 10.6151
R5870 VDD.n3341 VDD.n3340 10.6151
R5871 VDD.n3341 VDD.n849 10.6151
R5872 VDD.n3351 VDD.n849 10.6151
R5873 VDD.n3352 VDD.n3351 10.6151
R5874 VDD.n3353 VDD.n3352 10.6151
R5875 VDD.n3353 VDD.n836 10.6151
R5876 VDD.n3363 VDD.n836 10.6151
R5877 VDD.n3364 VDD.n3363 10.6151
R5878 VDD.n3365 VDD.n3364 10.6151
R5879 VDD.n3365 VDD.n825 10.6151
R5880 VDD.n3375 VDD.n825 10.6151
R5881 VDD.n3376 VDD.n3375 10.6151
R5882 VDD.n3377 VDD.n3376 10.6151
R5883 VDD.n3377 VDD.n812 10.6151
R5884 VDD.n3387 VDD.n812 10.6151
R5885 VDD.n3388 VDD.n3387 10.6151
R5886 VDD.n3389 VDD.n3388 10.6151
R5887 VDD.n3389 VDD.n800 10.6151
R5888 VDD.n3399 VDD.n800 10.6151
R5889 VDD.n3400 VDD.n3399 10.6151
R5890 VDD.n3401 VDD.n3400 10.6151
R5891 VDD.n3401 VDD.n789 10.6151
R5892 VDD.n3411 VDD.n789 10.6151
R5893 VDD.n3412 VDD.n3411 10.6151
R5894 VDD.n3413 VDD.n3412 10.6151
R5895 VDD.n3413 VDD.n776 10.6151
R5896 VDD.n3423 VDD.n776 10.6151
R5897 VDD.n3424 VDD.n3423 10.6151
R5898 VDD.n3430 VDD.n3424 10.6151
R5899 VDD.n3430 VDD.n3429 10.6151
R5900 VDD.n3429 VDD.n3428 10.6151
R5901 VDD.n3428 VDD.n3427 10.6151
R5902 VDD.n3427 VDD.n3425 10.6151
R5903 VDD.n3425 VDD.n751 10.6151
R5904 VDD.n3517 VDD.n751 10.6151
R5905 VDD.n3518 VDD.n3517 10.6151
R5906 VDD.n3519 VDD.n3518 10.6151
R5907 VDD.n3519 VDD.n739 10.6151
R5908 VDD.n3529 VDD.n739 10.6151
R5909 VDD.n3530 VDD.n3529 10.6151
R5910 VDD.n3531 VDD.n3530 10.6151
R5911 VDD.n3531 VDD.n727 10.6151
R5912 VDD.n3541 VDD.n727 10.6151
R5913 VDD.n3542 VDD.n3541 10.6151
R5914 VDD.n3543 VDD.n3542 10.6151
R5915 VDD.n3543 VDD.n715 10.6151
R5916 VDD.n3553 VDD.n715 10.6151
R5917 VDD.n3554 VDD.n3553 10.6151
R5918 VDD.n3555 VDD.n3554 10.6151
R5919 VDD.n3555 VDD.n703 10.6151
R5920 VDD.n3565 VDD.n703 10.6151
R5921 VDD.n3566 VDD.n3565 10.6151
R5922 VDD.n3567 VDD.n3566 10.6151
R5923 VDD.n3567 VDD.n691 10.6151
R5924 VDD.n3577 VDD.n691 10.6151
R5925 VDD.n3578 VDD.n3577 10.6151
R5926 VDD.n3579 VDD.n3578 10.6151
R5927 VDD.n3579 VDD.n679 10.6151
R5928 VDD.n3589 VDD.n679 10.6151
R5929 VDD.n3590 VDD.n3589 10.6151
R5930 VDD.n3591 VDD.n3590 10.6151
R5931 VDD.n3591 VDD.n667 10.6151
R5932 VDD.n3601 VDD.n667 10.6151
R5933 VDD.n3602 VDD.n3601 10.6151
R5934 VDD.n3603 VDD.n3602 10.6151
R5935 VDD.n3603 VDD.n655 10.6151
R5936 VDD.n3613 VDD.n655 10.6151
R5937 VDD.n3614 VDD.n3613 10.6151
R5938 VDD.n3615 VDD.n3614 10.6151
R5939 VDD.n3615 VDD.n642 10.6151
R5940 VDD.n3625 VDD.n642 10.6151
R5941 VDD.n3626 VDD.n3625 10.6151
R5942 VDD.n3627 VDD.n3626 10.6151
R5943 VDD.n3627 VDD.n631 10.6151
R5944 VDD.n3637 VDD.n631 10.6151
R5945 VDD.n3638 VDD.n3637 10.6151
R5946 VDD.n3667 VDD.n3638 10.6151
R5947 VDD.n3667 VDD.n3666 10.6151
R5948 VDD.n3666 VDD.n3665 10.6151
R5949 VDD.n3665 VDD.n3664 10.6151
R5950 VDD.n3664 VDD.n3662 10.6151
R5951 VDD.n2900 VDD.n2899 10.6151
R5952 VDD.n2899 VDD.n2896 10.6151
R5953 VDD.n2896 VDD.n2895 10.6151
R5954 VDD.n2895 VDD.n2892 10.6151
R5955 VDD.n2892 VDD.n2891 10.6151
R5956 VDD.n2891 VDD.n2888 10.6151
R5957 VDD.n2888 VDD.n2887 10.6151
R5958 VDD.n2887 VDD.n2884 10.6151
R5959 VDD.n2884 VDD.n2883 10.6151
R5960 VDD.n2883 VDD.n2880 10.6151
R5961 VDD.n2880 VDD.n2879 10.6151
R5962 VDD.n2879 VDD.n2876 10.6151
R5963 VDD.n2876 VDD.n2875 10.6151
R5964 VDD.n2875 VDD.n2872 10.6151
R5965 VDD.n2872 VDD.n2871 10.6151
R5966 VDD.n2871 VDD.n2868 10.6151
R5967 VDD.n2866 VDD.n926 10.6151
R5968 VDD.n2972 VDD.n926 10.6151
R5969 VDD.n2481 VDD.n2480 10.6151
R5970 VDD.n2480 VDD.n2479 10.6151
R5971 VDD.n2479 VDD.n2477 10.6151
R5972 VDD.n2477 VDD.n2476 10.6151
R5973 VDD.n2476 VDD.n2474 10.6151
R5974 VDD.n2474 VDD.n2473 10.6151
R5975 VDD.n2473 VDD.n2471 10.6151
R5976 VDD.n2471 VDD.n2470 10.6151
R5977 VDD.n2470 VDD.n2307 10.6151
R5978 VDD.n2307 VDD.n2306 10.6151
R5979 VDD.n2306 VDD.n2304 10.6151
R5980 VDD.n2304 VDD.n2303 10.6151
R5981 VDD.n2303 VDD.n2301 10.6151
R5982 VDD.n2301 VDD.n2300 10.6151
R5983 VDD.n2300 VDD.n2298 10.6151
R5984 VDD.n2298 VDD.n2297 10.6151
R5985 VDD.n2297 VDD.n2295 10.6151
R5986 VDD.n2295 VDD.n2294 10.6151
R5987 VDD.n2294 VDD.n2292 10.6151
R5988 VDD.n2292 VDD.n2291 10.6151
R5989 VDD.n2291 VDD.n2289 10.6151
R5990 VDD.n2289 VDD.n2288 10.6151
R5991 VDD.n2288 VDD.n2286 10.6151
R5992 VDD.n2286 VDD.n2285 10.6151
R5993 VDD.n2285 VDD.n2283 10.6151
R5994 VDD.n2283 VDD.n2282 10.6151
R5995 VDD.n2282 VDD.n2280 10.6151
R5996 VDD.n2280 VDD.n2279 10.6151
R5997 VDD.n2279 VDD.n2277 10.6151
R5998 VDD.n2277 VDD.n2276 10.6151
R5999 VDD.n2276 VDD.n2274 10.6151
R6000 VDD.n2274 VDD.n2273 10.6151
R6001 VDD.n2273 VDD.n2271 10.6151
R6002 VDD.n2271 VDD.n2270 10.6151
R6003 VDD.n2270 VDD.n2268 10.6151
R6004 VDD.n2268 VDD.n2267 10.6151
R6005 VDD.n2267 VDD.n2265 10.6151
R6006 VDD.n2265 VDD.n2264 10.6151
R6007 VDD.n2264 VDD.n2262 10.6151
R6008 VDD.n2262 VDD.n2261 10.6151
R6009 VDD.n2261 VDD.n2259 10.6151
R6010 VDD.n2259 VDD.n2258 10.6151
R6011 VDD.n2258 VDD.n2256 10.6151
R6012 VDD.n2256 VDD.n2255 10.6151
R6013 VDD.n2255 VDD.n2253 10.6151
R6014 VDD.n2253 VDD.n2252 10.6151
R6015 VDD.n2252 VDD.n2250 10.6151
R6016 VDD.n2250 VDD.n2249 10.6151
R6017 VDD.n2249 VDD.n2247 10.6151
R6018 VDD.n2247 VDD.n2246 10.6151
R6019 VDD.n2246 VDD.n2244 10.6151
R6020 VDD.n2244 VDD.n2243 10.6151
R6021 VDD.n2243 VDD.n2241 10.6151
R6022 VDD.n2241 VDD.n2240 10.6151
R6023 VDD.n2240 VDD.n2238 10.6151
R6024 VDD.n2238 VDD.n2237 10.6151
R6025 VDD.n2237 VDD.n2235 10.6151
R6026 VDD.n2235 VDD.n2234 10.6151
R6027 VDD.n2234 VDD.n2232 10.6151
R6028 VDD.n2232 VDD.n2231 10.6151
R6029 VDD.n2231 VDD.n2229 10.6151
R6030 VDD.n2229 VDD.n2228 10.6151
R6031 VDD.n2228 VDD.n2226 10.6151
R6032 VDD.n2226 VDD.n2225 10.6151
R6033 VDD.n2225 VDD.n2223 10.6151
R6034 VDD.n2223 VDD.n2222 10.6151
R6035 VDD.n2222 VDD.n2220 10.6151
R6036 VDD.n2220 VDD.n2219 10.6151
R6037 VDD.n2219 VDD.n2217 10.6151
R6038 VDD.n2217 VDD.n2216 10.6151
R6039 VDD.n2216 VDD.n2214 10.6151
R6040 VDD.n2214 VDD.n2213 10.6151
R6041 VDD.n2213 VDD.n2211 10.6151
R6042 VDD.n2211 VDD.n2210 10.6151
R6043 VDD.n2210 VDD.n2208 10.6151
R6044 VDD.n2208 VDD.n2207 10.6151
R6045 VDD.n2207 VDD.n2205 10.6151
R6046 VDD.n2205 VDD.n2204 10.6151
R6047 VDD.n2204 VDD.n2202 10.6151
R6048 VDD.n2202 VDD.n2201 10.6151
R6049 VDD.n2201 VDD.n2199 10.6151
R6050 VDD.n2199 VDD.n2198 10.6151
R6051 VDD.n2198 VDD.n2196 10.6151
R6052 VDD.n2196 VDD.n2195 10.6151
R6053 VDD.n2195 VDD.n2193 10.6151
R6054 VDD.n2193 VDD.n2192 10.6151
R6055 VDD.n2192 VDD.n2190 10.6151
R6056 VDD.n2190 VDD.n2189 10.6151
R6057 VDD.n2189 VDD.n2187 10.6151
R6058 VDD.n2187 VDD.n2186 10.6151
R6059 VDD.n2186 VDD.n2184 10.6151
R6060 VDD.n2184 VDD.n2183 10.6151
R6061 VDD.n2183 VDD.n2181 10.6151
R6062 VDD.n2181 VDD.n927 10.6151
R6063 VDD.n2970 VDD.n927 10.6151
R6064 VDD.n2971 VDD.n2970 10.6151
R6065 VDD.n2162 VDD.n2161 10.6151
R6066 VDD.n2165 VDD.n2162 10.6151
R6067 VDD.n2166 VDD.n2165 10.6151
R6068 VDD.n2169 VDD.n2166 10.6151
R6069 VDD.n2170 VDD.n2169 10.6151
R6070 VDD.n2173 VDD.n2170 10.6151
R6071 VDD.n2174 VDD.n2173 10.6151
R6072 VDD.n2177 VDD.n2174 10.6151
R6073 VDD.n2178 VDD.n2177 10.6151
R6074 VDD.n2504 VDD.n2501 10.6151
R6075 VDD.n2501 VDD.n2498 10.6151
R6076 VDD.n2498 VDD.n2497 10.6151
R6077 VDD.n2497 VDD.n2494 10.6151
R6078 VDD.n2494 VDD.n2493 10.6151
R6079 VDD.n2493 VDD.n2490 10.6151
R6080 VDD.n2488 VDD.n2485 10.6151
R6081 VDD.n2485 VDD.n2484 10.6151
R6082 VDD.n2597 VDD.n1212 10.6151
R6083 VDD.n2598 VDD.n2597 10.6151
R6084 VDD.n2599 VDD.n2598 10.6151
R6085 VDD.n2599 VDD.n1200 10.6151
R6086 VDD.n2609 VDD.n1200 10.6151
R6087 VDD.n2610 VDD.n2609 10.6151
R6088 VDD.n2611 VDD.n2610 10.6151
R6089 VDD.n2611 VDD.n1189 10.6151
R6090 VDD.n2621 VDD.n1189 10.6151
R6091 VDD.n2622 VDD.n2621 10.6151
R6092 VDD.n2623 VDD.n2622 10.6151
R6093 VDD.n2623 VDD.n1177 10.6151
R6094 VDD.n2633 VDD.n1177 10.6151
R6095 VDD.n2634 VDD.n2633 10.6151
R6096 VDD.n2635 VDD.n2634 10.6151
R6097 VDD.n2635 VDD.n1165 10.6151
R6098 VDD.n2645 VDD.n1165 10.6151
R6099 VDD.n2646 VDD.n2645 10.6151
R6100 VDD.n2647 VDD.n2646 10.6151
R6101 VDD.n2647 VDD.n1153 10.6151
R6102 VDD.n2657 VDD.n1153 10.6151
R6103 VDD.n2658 VDD.n2657 10.6151
R6104 VDD.n2659 VDD.n2658 10.6151
R6105 VDD.n2659 VDD.n1141 10.6151
R6106 VDD.n2669 VDD.n1141 10.6151
R6107 VDD.n2670 VDD.n2669 10.6151
R6108 VDD.n2671 VDD.n2670 10.6151
R6109 VDD.n2671 VDD.n1129 10.6151
R6110 VDD.n2681 VDD.n1129 10.6151
R6111 VDD.n2682 VDD.n2681 10.6151
R6112 VDD.n2683 VDD.n2682 10.6151
R6113 VDD.n2683 VDD.n1117 10.6151
R6114 VDD.n2693 VDD.n1117 10.6151
R6115 VDD.n2694 VDD.n2693 10.6151
R6116 VDD.n2695 VDD.n2694 10.6151
R6117 VDD.n2695 VDD.n1105 10.6151
R6118 VDD.n2705 VDD.n1105 10.6151
R6119 VDD.n2706 VDD.n2705 10.6151
R6120 VDD.n2707 VDD.n2706 10.6151
R6121 VDD.n2707 VDD.n1093 10.6151
R6122 VDD.n2717 VDD.n1093 10.6151
R6123 VDD.n2718 VDD.n2717 10.6151
R6124 VDD.n2719 VDD.n2718 10.6151
R6125 VDD.n2719 VDD.n1081 10.6151
R6126 VDD.n2729 VDD.n1081 10.6151
R6127 VDD.n2730 VDD.n2729 10.6151
R6128 VDD.n2731 VDD.n2730 10.6151
R6129 VDD.n2731 VDD.n1070 10.6151
R6130 VDD.n2741 VDD.n1070 10.6151
R6131 VDD.n2742 VDD.n2741 10.6151
R6132 VDD.n2743 VDD.n2742 10.6151
R6133 VDD.n2743 VDD.n1058 10.6151
R6134 VDD.n2753 VDD.n1058 10.6151
R6135 VDD.n2754 VDD.n2753 10.6151
R6136 VDD.n2755 VDD.n2754 10.6151
R6137 VDD.n2755 VDD.n1046 10.6151
R6138 VDD.n2765 VDD.n1046 10.6151
R6139 VDD.n2766 VDD.n2765 10.6151
R6140 VDD.n2767 VDD.n2766 10.6151
R6141 VDD.n2767 VDD.n1034 10.6151
R6142 VDD.n2777 VDD.n1034 10.6151
R6143 VDD.n2778 VDD.n2777 10.6151
R6144 VDD.n2779 VDD.n2778 10.6151
R6145 VDD.n2779 VDD.n1022 10.6151
R6146 VDD.n2789 VDD.n1022 10.6151
R6147 VDD.n2790 VDD.n2789 10.6151
R6148 VDD.n2791 VDD.n2790 10.6151
R6149 VDD.n2791 VDD.n1010 10.6151
R6150 VDD.n2801 VDD.n1010 10.6151
R6151 VDD.n2802 VDD.n2801 10.6151
R6152 VDD.n2803 VDD.n2802 10.6151
R6153 VDD.n2803 VDD.n998 10.6151
R6154 VDD.n2813 VDD.n998 10.6151
R6155 VDD.n2814 VDD.n2813 10.6151
R6156 VDD.n2815 VDD.n2814 10.6151
R6157 VDD.n2815 VDD.n986 10.6151
R6158 VDD.n2825 VDD.n986 10.6151
R6159 VDD.n2826 VDD.n2825 10.6151
R6160 VDD.n2827 VDD.n2826 10.6151
R6161 VDD.n2827 VDD.n974 10.6151
R6162 VDD.n2837 VDD.n974 10.6151
R6163 VDD.n2838 VDD.n2837 10.6151
R6164 VDD.n2839 VDD.n2838 10.6151
R6165 VDD.n2839 VDD.n962 10.6151
R6166 VDD.n2849 VDD.n962 10.6151
R6167 VDD.n2850 VDD.n2849 10.6151
R6168 VDD.n2851 VDD.n2850 10.6151
R6169 VDD.n2851 VDD.n950 10.6151
R6170 VDD.n2861 VDD.n950 10.6151
R6171 VDD.n2862 VDD.n2861 10.6151
R6172 VDD.n2909 VDD.n2862 10.6151
R6173 VDD.n2909 VDD.n2908 10.6151
R6174 VDD.n2908 VDD.n2907 10.6151
R6175 VDD.n2907 VDD.n2906 10.6151
R6176 VDD.n2906 VDD.n2904 10.6151
R6177 VDD.n2904 VDD.n2903 10.6151
R6178 VDD.n2593 VDD.n2592 10.6151
R6179 VDD.n2593 VDD.n1206 10.6151
R6180 VDD.n2603 VDD.n1206 10.6151
R6181 VDD.n2604 VDD.n2603 10.6151
R6182 VDD.n2605 VDD.n2604 10.6151
R6183 VDD.n2605 VDD.n1194 10.6151
R6184 VDD.n2615 VDD.n1194 10.6151
R6185 VDD.n2616 VDD.n2615 10.6151
R6186 VDD.n2617 VDD.n2616 10.6151
R6187 VDD.n2617 VDD.n1183 10.6151
R6188 VDD.n2627 VDD.n1183 10.6151
R6189 VDD.n2628 VDD.n2627 10.6151
R6190 VDD.n2629 VDD.n2628 10.6151
R6191 VDD.n2629 VDD.n1171 10.6151
R6192 VDD.n2639 VDD.n1171 10.6151
R6193 VDD.n2640 VDD.n2639 10.6151
R6194 VDD.n2641 VDD.n2640 10.6151
R6195 VDD.n2641 VDD.n1159 10.6151
R6196 VDD.n2651 VDD.n1159 10.6151
R6197 VDD.n2652 VDD.n2651 10.6151
R6198 VDD.n2653 VDD.n2652 10.6151
R6199 VDD.n2653 VDD.n1147 10.6151
R6200 VDD.n2663 VDD.n1147 10.6151
R6201 VDD.n2664 VDD.n2663 10.6151
R6202 VDD.n2665 VDD.n2664 10.6151
R6203 VDD.n2665 VDD.n1135 10.6151
R6204 VDD.n2675 VDD.n1135 10.6151
R6205 VDD.n2676 VDD.n2675 10.6151
R6206 VDD.n2677 VDD.n2676 10.6151
R6207 VDD.n2677 VDD.n1123 10.6151
R6208 VDD.n2687 VDD.n1123 10.6151
R6209 VDD.n2688 VDD.n2687 10.6151
R6210 VDD.n2689 VDD.n2688 10.6151
R6211 VDD.n2689 VDD.n1111 10.6151
R6212 VDD.n2699 VDD.n1111 10.6151
R6213 VDD.n2700 VDD.n2699 10.6151
R6214 VDD.n2701 VDD.n2700 10.6151
R6215 VDD.n2701 VDD.n1099 10.6151
R6216 VDD.n2711 VDD.n1099 10.6151
R6217 VDD.n2712 VDD.n2711 10.6151
R6218 VDD.n2713 VDD.n2712 10.6151
R6219 VDD.n2713 VDD.n1087 10.6151
R6220 VDD.n2723 VDD.n1087 10.6151
R6221 VDD.n2724 VDD.n2723 10.6151
R6222 VDD.n2725 VDD.n2724 10.6151
R6223 VDD.n2725 VDD.n1075 10.6151
R6224 VDD.n2735 VDD.n1075 10.6151
R6225 VDD.n2736 VDD.n2735 10.6151
R6226 VDD.n2737 VDD.n2736 10.6151
R6227 VDD.n2737 VDD.n1063 10.6151
R6228 VDD.n2747 VDD.n1063 10.6151
R6229 VDD.n2748 VDD.n2747 10.6151
R6230 VDD.n2749 VDD.n2748 10.6151
R6231 VDD.n2749 VDD.n1052 10.6151
R6232 VDD.n2759 VDD.n1052 10.6151
R6233 VDD.n2760 VDD.n2759 10.6151
R6234 VDD.n2761 VDD.n2760 10.6151
R6235 VDD.n2761 VDD.n1039 10.6151
R6236 VDD.n2771 VDD.n1039 10.6151
R6237 VDD.n2772 VDD.n2771 10.6151
R6238 VDD.n2773 VDD.n2772 10.6151
R6239 VDD.n2773 VDD.n1027 10.6151
R6240 VDD.n2783 VDD.n1027 10.6151
R6241 VDD.n2784 VDD.n2783 10.6151
R6242 VDD.n2785 VDD.n2784 10.6151
R6243 VDD.n2785 VDD.n1016 10.6151
R6244 VDD.n2795 VDD.n1016 10.6151
R6245 VDD.n2796 VDD.n2795 10.6151
R6246 VDD.n2797 VDD.n2796 10.6151
R6247 VDD.n2797 VDD.n1003 10.6151
R6248 VDD.n2807 VDD.n1003 10.6151
R6249 VDD.n2808 VDD.n2807 10.6151
R6250 VDD.n2809 VDD.n2808 10.6151
R6251 VDD.n2809 VDD.n992 10.6151
R6252 VDD.n2819 VDD.n992 10.6151
R6253 VDD.n2820 VDD.n2819 10.6151
R6254 VDD.n2821 VDD.n2820 10.6151
R6255 VDD.n2821 VDD.n980 10.6151
R6256 VDD.n2831 VDD.n980 10.6151
R6257 VDD.n2832 VDD.n2831 10.6151
R6258 VDD.n2833 VDD.n2832 10.6151
R6259 VDD.n2833 VDD.n968 10.6151
R6260 VDD.n2843 VDD.n968 10.6151
R6261 VDD.n2844 VDD.n2843 10.6151
R6262 VDD.n2845 VDD.n2844 10.6151
R6263 VDD.n2845 VDD.n955 10.6151
R6264 VDD.n2855 VDD.n955 10.6151
R6265 VDD.n2856 VDD.n2855 10.6151
R6266 VDD.n2857 VDD.n2856 10.6151
R6267 VDD.n2857 VDD.n943 10.6151
R6268 VDD.n2913 VDD.n943 10.6151
R6269 VDD.n2914 VDD.n2913 10.6151
R6270 VDD.n2915 VDD.n2914 10.6151
R6271 VDD.n2915 VDD.n934 10.6151
R6272 VDD.n2966 VDD.n934 10.6151
R6273 VDD.n2966 VDD.n2965 10.6151
R6274 VDD.n2964 VDD.n2962 10.6151
R6275 VDD.n2962 VDD.n2959 10.6151
R6276 VDD.n2959 VDD.n2958 10.6151
R6277 VDD.n2958 VDD.n2955 10.6151
R6278 VDD.n2955 VDD.n2954 10.6151
R6279 VDD.n2954 VDD.n2951 10.6151
R6280 VDD.n2951 VDD.n2950 10.6151
R6281 VDD.n2950 VDD.n2947 10.6151
R6282 VDD.n2947 VDD.n2946 10.6151
R6283 VDD.n2946 VDD.n2943 10.6151
R6284 VDD.n2943 VDD.n2942 10.6151
R6285 VDD.n2942 VDD.n2939 10.6151
R6286 VDD.n2939 VDD.n2938 10.6151
R6287 VDD.n2938 VDD.n2935 10.6151
R6288 VDD.n2935 VDD.n2934 10.6151
R6289 VDD.n2934 VDD.n2931 10.6151
R6290 VDD.n2929 VDD.n2926 10.6151
R6291 VDD.n2926 VDD.n2925 10.6151
R6292 VDD.n2331 VDD.n2330 10.6151
R6293 VDD.n2333 VDD.n2331 10.6151
R6294 VDD.n2334 VDD.n2333 10.6151
R6295 VDD.n2336 VDD.n2334 10.6151
R6296 VDD.n2337 VDD.n2336 10.6151
R6297 VDD.n2339 VDD.n2337 10.6151
R6298 VDD.n2340 VDD.n2339 10.6151
R6299 VDD.n2466 VDD.n2340 10.6151
R6300 VDD.n2466 VDD.n2465 10.6151
R6301 VDD.n2465 VDD.n2464 10.6151
R6302 VDD.n2464 VDD.n2462 10.6151
R6303 VDD.n2462 VDD.n2461 10.6151
R6304 VDD.n2461 VDD.n2459 10.6151
R6305 VDD.n2459 VDD.n2458 10.6151
R6306 VDD.n2458 VDD.n2456 10.6151
R6307 VDD.n2456 VDD.n2455 10.6151
R6308 VDD.n2455 VDD.n2453 10.6151
R6309 VDD.n2453 VDD.n2452 10.6151
R6310 VDD.n2452 VDD.n2450 10.6151
R6311 VDD.n2450 VDD.n2449 10.6151
R6312 VDD.n2449 VDD.n2447 10.6151
R6313 VDD.n2447 VDD.n2446 10.6151
R6314 VDD.n2446 VDD.n2444 10.6151
R6315 VDD.n2444 VDD.n2443 10.6151
R6316 VDD.n2443 VDD.n2441 10.6151
R6317 VDD.n2441 VDD.n2440 10.6151
R6318 VDD.n2440 VDD.n2438 10.6151
R6319 VDD.n2438 VDD.n2437 10.6151
R6320 VDD.n2437 VDD.n2435 10.6151
R6321 VDD.n2435 VDD.n2434 10.6151
R6322 VDD.n2434 VDD.n2432 10.6151
R6323 VDD.n2432 VDD.n2431 10.6151
R6324 VDD.n2431 VDD.n2429 10.6151
R6325 VDD.n2429 VDD.n2428 10.6151
R6326 VDD.n2428 VDD.n2426 10.6151
R6327 VDD.n2426 VDD.n2425 10.6151
R6328 VDD.n2425 VDD.n2423 10.6151
R6329 VDD.n2423 VDD.n2422 10.6151
R6330 VDD.n2422 VDD.n2420 10.6151
R6331 VDD.n2420 VDD.n2419 10.6151
R6332 VDD.n2419 VDD.n2417 10.6151
R6333 VDD.n2417 VDD.n2416 10.6151
R6334 VDD.n2416 VDD.n2414 10.6151
R6335 VDD.n2414 VDD.n2413 10.6151
R6336 VDD.n2413 VDD.n2411 10.6151
R6337 VDD.n2411 VDD.n2410 10.6151
R6338 VDD.n2410 VDD.n2408 10.6151
R6339 VDD.n2408 VDD.n2407 10.6151
R6340 VDD.n2407 VDD.n2405 10.6151
R6341 VDD.n2405 VDD.n2404 10.6151
R6342 VDD.n2404 VDD.n2402 10.6151
R6343 VDD.n2402 VDD.n2401 10.6151
R6344 VDD.n2401 VDD.n2399 10.6151
R6345 VDD.n2399 VDD.n2398 10.6151
R6346 VDD.n2398 VDD.n2396 10.6151
R6347 VDD.n2396 VDD.n2395 10.6151
R6348 VDD.n2395 VDD.n2393 10.6151
R6349 VDD.n2393 VDD.n2392 10.6151
R6350 VDD.n2392 VDD.n2390 10.6151
R6351 VDD.n2390 VDD.n2389 10.6151
R6352 VDD.n2389 VDD.n2387 10.6151
R6353 VDD.n2387 VDD.n2386 10.6151
R6354 VDD.n2386 VDD.n2384 10.6151
R6355 VDD.n2384 VDD.n2383 10.6151
R6356 VDD.n2383 VDD.n2381 10.6151
R6357 VDD.n2381 VDD.n2380 10.6151
R6358 VDD.n2380 VDD.n2378 10.6151
R6359 VDD.n2378 VDD.n2377 10.6151
R6360 VDD.n2377 VDD.n2375 10.6151
R6361 VDD.n2375 VDD.n2374 10.6151
R6362 VDD.n2374 VDD.n2372 10.6151
R6363 VDD.n2372 VDD.n2371 10.6151
R6364 VDD.n2371 VDD.n2369 10.6151
R6365 VDD.n2369 VDD.n2368 10.6151
R6366 VDD.n2368 VDD.n2366 10.6151
R6367 VDD.n2366 VDD.n2365 10.6151
R6368 VDD.n2365 VDD.n2363 10.6151
R6369 VDD.n2363 VDD.n2362 10.6151
R6370 VDD.n2362 VDD.n2360 10.6151
R6371 VDD.n2360 VDD.n2359 10.6151
R6372 VDD.n2359 VDD.n2357 10.6151
R6373 VDD.n2357 VDD.n2356 10.6151
R6374 VDD.n2356 VDD.n2354 10.6151
R6375 VDD.n2354 VDD.n2353 10.6151
R6376 VDD.n2353 VDD.n2351 10.6151
R6377 VDD.n2351 VDD.n2350 10.6151
R6378 VDD.n2350 VDD.n2348 10.6151
R6379 VDD.n2348 VDD.n2347 10.6151
R6380 VDD.n2347 VDD.n2345 10.6151
R6381 VDD.n2345 VDD.n2344 10.6151
R6382 VDD.n2344 VDD.n2342 10.6151
R6383 VDD.n2342 VDD.n2341 10.6151
R6384 VDD.n2341 VDD.n937 10.6151
R6385 VDD.n2920 VDD.n937 10.6151
R6386 VDD.n2921 VDD.n2920 10.6151
R6387 VDD.n2922 VDD.n2921 10.6151
R6388 VDD.n2591 VDD.n1218 10.6151
R6389 VDD.n2586 VDD.n1218 10.6151
R6390 VDD.n2586 VDD.n2585 10.6151
R6391 VDD.n2585 VDD.n2584 10.6151
R6392 VDD.n2584 VDD.n2581 10.6151
R6393 VDD.n2581 VDD.n2580 10.6151
R6394 VDD.n2580 VDD.n2577 10.6151
R6395 VDD.n2577 VDD.n2576 10.6151
R6396 VDD.n2576 VDD.n2573 10.6151
R6397 VDD.n2313 VDD.n1240 10.6151
R6398 VDD.n2314 VDD.n2313 10.6151
R6399 VDD.n2317 VDD.n2314 10.6151
R6400 VDD.n2318 VDD.n2317 10.6151
R6401 VDD.n2321 VDD.n2318 10.6151
R6402 VDD.n2322 VDD.n2321 10.6151
R6403 VDD.n2327 VDD.n2325 10.6151
R6404 VDD.n2328 VDD.n2327 10.6151
R6405 VDD.t36 VDD.n1143 10.4784
R6406 VDD.n1008 VDD.t14 10.4784
R6407 VDD.n3367 VDD.t11 10.4784
R6408 VDD.n3581 VDD.t45 10.4784
R6409 VDD.n2551 VDD.n2550 10.0853
R6410 VDD.n1711 VDD.n1710 10.0853
R6411 VDD.n581 VDD.n578 10.0853
R6412 VDD.n246 VDD.n207 10.0853
R6413 VDD.n3739 VDD.n3738 10.0608
R6414 VDD.n2506 VDD.n2505 10.0608
R6415 VDD.n1457 VDD.n1456 9.3005
R6416 VDD.n1970 VDD.n1969 9.3005
R6417 VDD.n1971 VDD.n1455 9.3005
R6418 VDD.n1973 VDD.n1972 9.3005
R6419 VDD.n1445 VDD.n1444 9.3005
R6420 VDD.n1986 VDD.n1985 9.3005
R6421 VDD.n1987 VDD.n1443 9.3005
R6422 VDD.n1989 VDD.n1988 9.3005
R6423 VDD.n1433 VDD.n1432 9.3005
R6424 VDD.n2003 VDD.n2002 9.3005
R6425 VDD.n2004 VDD.n1431 9.3005
R6426 VDD.n2006 VDD.n2005 9.3005
R6427 VDD.n1422 VDD.n1421 9.3005
R6428 VDD.n2019 VDD.n2018 9.3005
R6429 VDD.n2020 VDD.n1420 9.3005
R6430 VDD.n2022 VDD.n2021 9.3005
R6431 VDD.n1410 VDD.n1409 9.3005
R6432 VDD.n2035 VDD.n2034 9.3005
R6433 VDD.n2036 VDD.n1408 9.3005
R6434 VDD.n2038 VDD.n2037 9.3005
R6435 VDD.n1398 VDD.n1397 9.3005
R6436 VDD.n2051 VDD.n2050 9.3005
R6437 VDD.n2052 VDD.n1396 9.3005
R6438 VDD.n2054 VDD.n2053 9.3005
R6439 VDD.n1386 VDD.n1385 9.3005
R6440 VDD.n2067 VDD.n2066 9.3005
R6441 VDD.n2068 VDD.n1384 9.3005
R6442 VDD.n2070 VDD.n2069 9.3005
R6443 VDD.n1374 VDD.n1373 9.3005
R6444 VDD.n2083 VDD.n2082 9.3005
R6445 VDD.n2084 VDD.n1372 9.3005
R6446 VDD.n2086 VDD.n2085 9.3005
R6447 VDD.n1362 VDD.n1361 9.3005
R6448 VDD.n2099 VDD.n2098 9.3005
R6449 VDD.n2100 VDD.n1360 9.3005
R6450 VDD.n2102 VDD.n2101 9.3005
R6451 VDD.n1350 VDD.n1349 9.3005
R6452 VDD.n2115 VDD.n2114 9.3005
R6453 VDD.n2116 VDD.n1348 9.3005
R6454 VDD.n2118 VDD.n2117 9.3005
R6455 VDD.n1338 VDD.n1337 9.3005
R6456 VDD.n2131 VDD.n2130 9.3005
R6457 VDD.n2132 VDD.n1336 9.3005
R6458 VDD.n2134 VDD.n2133 9.3005
R6459 VDD.n1325 VDD.n1324 9.3005
R6460 VDD.n2149 VDD.n2148 9.3005
R6461 VDD.n2150 VDD.n1323 9.3005
R6462 VDD.n2152 VDD.n2151 9.3005
R6463 VDD.n1312 VDD.n1311 9.3005
R6464 VDD.n2516 VDD.n2515 9.3005
R6465 VDD.n2517 VDD.n1310 9.3005
R6466 VDD.n2519 VDD.n2518 9.3005
R6467 VDD.n2520 VDD.n1241 9.3005
R6468 VDD.n3742 VDD.n3741 9.3005
R6469 VDD.n458 VDD.n457 9.3005
R6470 VDD.n3755 VDD.n3754 9.3005
R6471 VDD.n3756 VDD.n456 9.3005
R6472 VDD.n3758 VDD.n3757 9.3005
R6473 VDD.n446 VDD.n445 9.3005
R6474 VDD.n3771 VDD.n3770 9.3005
R6475 VDD.n3772 VDD.n444 9.3005
R6476 VDD.n3774 VDD.n3773 9.3005
R6477 VDD.n434 VDD.n433 9.3005
R6478 VDD.n3787 VDD.n3786 9.3005
R6479 VDD.n3788 VDD.n432 9.3005
R6480 VDD.n3790 VDD.n3789 9.3005
R6481 VDD.n422 VDD.n421 9.3005
R6482 VDD.n3803 VDD.n3802 9.3005
R6483 VDD.n3804 VDD.n420 9.3005
R6484 VDD.n3806 VDD.n3805 9.3005
R6485 VDD.n410 VDD.n409 9.3005
R6486 VDD.n3819 VDD.n3818 9.3005
R6487 VDD.n3820 VDD.n408 9.3005
R6488 VDD.n3822 VDD.n3821 9.3005
R6489 VDD.n398 VDD.n397 9.3005
R6490 VDD.n3835 VDD.n3834 9.3005
R6491 VDD.n3836 VDD.n396 9.3005
R6492 VDD.n3838 VDD.n3837 9.3005
R6493 VDD.n386 VDD.n385 9.3005
R6494 VDD.n3851 VDD.n3850 9.3005
R6495 VDD.n3852 VDD.n384 9.3005
R6496 VDD.n3854 VDD.n3853 9.3005
R6497 VDD.n375 VDD.n374 9.3005
R6498 VDD.n3868 VDD.n3867 9.3005
R6499 VDD.n3869 VDD.n373 9.3005
R6500 VDD.n3871 VDD.n3870 9.3005
R6501 VDD.n363 VDD.n362 9.3005
R6502 VDD.n3884 VDD.n3883 9.3005
R6503 VDD.n3885 VDD.n361 9.3005
R6504 VDD.n3887 VDD.n3886 9.3005
R6505 VDD.n351 VDD.n350 9.3005
R6506 VDD.n3900 VDD.n3899 9.3005
R6507 VDD.n3901 VDD.n349 9.3005
R6508 VDD.n3903 VDD.n3902 9.3005
R6509 VDD.n339 VDD.n338 9.3005
R6510 VDD.n3916 VDD.n3915 9.3005
R6511 VDD.n3917 VDD.n337 9.3005
R6512 VDD.n3919 VDD.n3918 9.3005
R6513 VDD.n327 VDD.n326 9.3005
R6514 VDD.n3932 VDD.n3931 9.3005
R6515 VDD.n3933 VDD.n325 9.3005
R6516 VDD.n3938 VDD.n3934 9.3005
R6517 VDD.n3937 VDD.n3936 9.3005
R6518 VDD.n3935 VDD.n314 9.3005
R6519 VDD.n3951 VDD.n315 9.3005
R6520 VDD.n3952 VDD.n313 9.3005
R6521 VDD.n3954 VDD.n3953 9.3005
R6522 VDD.n3955 VDD.n312 9.3005
R6523 VDD.n3958 VDD.n3956 9.3005
R6524 VDD.n3959 VDD.n311 9.3005
R6525 VDD.n3961 VDD.n3960 9.3005
R6526 VDD.n3962 VDD.n310 9.3005
R6527 VDD.n3965 VDD.n3963 9.3005
R6528 VDD.n3966 VDD.n309 9.3005
R6529 VDD.n3968 VDD.n3967 9.3005
R6530 VDD.n3969 VDD.n308 9.3005
R6531 VDD.n3972 VDD.n3970 9.3005
R6532 VDD.n3973 VDD.n307 9.3005
R6533 VDD.n3975 VDD.n3974 9.3005
R6534 VDD.n3976 VDD.n306 9.3005
R6535 VDD.n3979 VDD.n3977 9.3005
R6536 VDD.n3980 VDD.n305 9.3005
R6537 VDD.n3982 VDD.n3981 9.3005
R6538 VDD.n3983 VDD.n304 9.3005
R6539 VDD.n3986 VDD.n3984 9.3005
R6540 VDD.n3987 VDD.n303 9.3005
R6541 VDD.n3989 VDD.n3988 9.3005
R6542 VDD.n3990 VDD.n302 9.3005
R6543 VDD.n3993 VDD.n3991 9.3005
R6544 VDD.n3994 VDD.n301 9.3005
R6545 VDD.n3996 VDD.n3995 9.3005
R6546 VDD.n3997 VDD.n300 9.3005
R6547 VDD.n4000 VDD.n3998 9.3005
R6548 VDD.n4001 VDD.n299 9.3005
R6549 VDD.n4003 VDD.n4002 9.3005
R6550 VDD.n4004 VDD.n298 9.3005
R6551 VDD.n4007 VDD.n4005 9.3005
R6552 VDD.n4008 VDD.n297 9.3005
R6553 VDD.n4010 VDD.n4009 9.3005
R6554 VDD.n4011 VDD.n296 9.3005
R6555 VDD.n4014 VDD.n4012 9.3005
R6556 VDD.n4015 VDD.n295 9.3005
R6557 VDD.n4017 VDD.n4016 9.3005
R6558 VDD.n4018 VDD.n294 9.3005
R6559 VDD.n4021 VDD.n4019 9.3005
R6560 VDD.n4022 VDD.n293 9.3005
R6561 VDD.n4024 VDD.n4023 9.3005
R6562 VDD.n4025 VDD.n292 9.3005
R6563 VDD.n4028 VDD.n4026 9.3005
R6564 VDD.n4029 VDD.n291 9.3005
R6565 VDD.n4031 VDD.n4030 9.3005
R6566 VDD.n4032 VDD.n290 9.3005
R6567 VDD.n4035 VDD.n4033 9.3005
R6568 VDD.n4036 VDD.n289 9.3005
R6569 VDD.n4038 VDD.n4037 9.3005
R6570 VDD.n4039 VDD.n288 9.3005
R6571 VDD.n4042 VDD.n4040 9.3005
R6572 VDD.n4043 VDD.n287 9.3005
R6573 VDD.n4045 VDD.n4044 9.3005
R6574 VDD.n3740 VDD.n468 9.3005
R6575 VDD.n218 VDD.n213 9.3005
R6576 VDD.n222 VDD.n219 9.3005
R6577 VDD.n223 VDD.n212 9.3005
R6578 VDD.n227 VDD.n226 9.3005
R6579 VDD.n228 VDD.n211 9.3005
R6580 VDD.n232 VDD.n229 9.3005
R6581 VDD.n233 VDD.n210 9.3005
R6582 VDD.n237 VDD.n236 9.3005
R6583 VDD.n238 VDD.n209 9.3005
R6584 VDD.n242 VDD.n239 9.3005
R6585 VDD.n243 VDD.n208 9.3005
R6586 VDD.n247 VDD.n246 9.3005
R6587 VDD.n248 VDD.n207 9.3005
R6588 VDD.n252 VDD.n249 9.3005
R6589 VDD.n253 VDD.n204 9.3005
R6590 VDD.n257 VDD.n256 9.3005
R6591 VDD.n258 VDD.n203 9.3005
R6592 VDD.n262 VDD.n259 9.3005
R6593 VDD.n263 VDD.n202 9.3005
R6594 VDD.n267 VDD.n266 9.3005
R6595 VDD.n268 VDD.n201 9.3005
R6596 VDD.n272 VDD.n269 9.3005
R6597 VDD.n273 VDD.n200 9.3005
R6598 VDD.n277 VDD.n276 9.3005
R6599 VDD.n278 VDD.n199 9.3005
R6600 VDD.n282 VDD.n279 9.3005
R6601 VDD.n284 VDD.n198 9.3005
R6602 VDD.n286 VDD.n285 9.3005
R6603 VDD.n4047 VDD.n4046 9.3005
R6604 VDD.n217 VDD.n216 9.3005
R6605 VDD.n32 VDD.n30 9.3005
R6606 VDD.n4152 VDD.n41 9.3005
R6607 VDD.n4151 VDD.n42 9.3005
R6608 VDD.n4150 VDD.n43 9.3005
R6609 VDD.n51 VDD.n44 9.3005
R6610 VDD.n4144 VDD.n52 9.3005
R6611 VDD.n4143 VDD.n53 9.3005
R6612 VDD.n4142 VDD.n54 9.3005
R6613 VDD.n62 VDD.n55 9.3005
R6614 VDD.n4136 VDD.n63 9.3005
R6615 VDD.n4135 VDD.n64 9.3005
R6616 VDD.n4134 VDD.n65 9.3005
R6617 VDD.n73 VDD.n66 9.3005
R6618 VDD.n4128 VDD.n74 9.3005
R6619 VDD.n4127 VDD.n75 9.3005
R6620 VDD.n4126 VDD.n76 9.3005
R6621 VDD.n84 VDD.n77 9.3005
R6622 VDD.n4120 VDD.n85 9.3005
R6623 VDD.n4119 VDD.n86 9.3005
R6624 VDD.n4118 VDD.n87 9.3005
R6625 VDD.n94 VDD.n88 9.3005
R6626 VDD.n4112 VDD.n95 9.3005
R6627 VDD.n4111 VDD.n96 9.3005
R6628 VDD.n4110 VDD.n97 9.3005
R6629 VDD.n106 VDD.n98 9.3005
R6630 VDD.n4104 VDD.n107 9.3005
R6631 VDD.n4103 VDD.n108 9.3005
R6632 VDD.n4102 VDD.n109 9.3005
R6633 VDD.n117 VDD.n110 9.3005
R6634 VDD.n4096 VDD.n118 9.3005
R6635 VDD.n4095 VDD.n119 9.3005
R6636 VDD.n4094 VDD.n120 9.3005
R6637 VDD.n128 VDD.n121 9.3005
R6638 VDD.n4088 VDD.n129 9.3005
R6639 VDD.n4087 VDD.n130 9.3005
R6640 VDD.n4086 VDD.n131 9.3005
R6641 VDD.n139 VDD.n132 9.3005
R6642 VDD.n4080 VDD.n140 9.3005
R6643 VDD.n4079 VDD.n141 9.3005
R6644 VDD.n4078 VDD.n142 9.3005
R6645 VDD.n150 VDD.n143 9.3005
R6646 VDD.n4072 VDD.n151 9.3005
R6647 VDD.n4071 VDD.n152 9.3005
R6648 VDD.n4070 VDD.n153 9.3005
R6649 VDD.n161 VDD.n154 9.3005
R6650 VDD.n4064 VDD.n162 9.3005
R6651 VDD.n4063 VDD.n163 9.3005
R6652 VDD.n4062 VDD.n164 9.3005
R6653 VDD.n172 VDD.n165 9.3005
R6654 VDD.n4056 VDD.n173 9.3005
R6655 VDD.n4055 VDD.n174 9.3005
R6656 VDD.n4054 VDD.n175 9.3005
R6657 VDD.n214 VDD.n176 9.3005
R6658 VDD.n4158 VDD.n4157 9.3005
R6659 VDD.n3747 VDD.n3746 9.3005
R6660 VDD.n3748 VDD.n462 9.3005
R6661 VDD.n3750 VDD.n3749 9.3005
R6662 VDD.n452 VDD.n451 9.3005
R6663 VDD.n3763 VDD.n3762 9.3005
R6664 VDD.n3764 VDD.n450 9.3005
R6665 VDD.n3766 VDD.n3765 9.3005
R6666 VDD.n440 VDD.n439 9.3005
R6667 VDD.n3779 VDD.n3778 9.3005
R6668 VDD.n3780 VDD.n438 9.3005
R6669 VDD.n3782 VDD.n3781 9.3005
R6670 VDD.n428 VDD.n427 9.3005
R6671 VDD.n3795 VDD.n3794 9.3005
R6672 VDD.n3796 VDD.n426 9.3005
R6673 VDD.n3798 VDD.n3797 9.3005
R6674 VDD.n416 VDD.n415 9.3005
R6675 VDD.n3811 VDD.n3810 9.3005
R6676 VDD.n3812 VDD.n414 9.3005
R6677 VDD.n3814 VDD.n3813 9.3005
R6678 VDD.n404 VDD.n403 9.3005
R6679 VDD.n3827 VDD.n3826 9.3005
R6680 VDD.n3828 VDD.n402 9.3005
R6681 VDD.n3830 VDD.n3829 9.3005
R6682 VDD.n392 VDD.n391 9.3005
R6683 VDD.n3843 VDD.n3842 9.3005
R6684 VDD.n3844 VDD.n390 9.3005
R6685 VDD.n3846 VDD.n3845 9.3005
R6686 VDD.n380 VDD.n379 9.3005
R6687 VDD.n3860 VDD.n3859 9.3005
R6688 VDD.n3861 VDD.n378 9.3005
R6689 VDD.n3863 VDD.n3862 9.3005
R6690 VDD.n369 VDD.n368 9.3005
R6691 VDD.n3876 VDD.n3875 9.3005
R6692 VDD.n3877 VDD.n367 9.3005
R6693 VDD.n3879 VDD.n3878 9.3005
R6694 VDD.n357 VDD.n356 9.3005
R6695 VDD.n3892 VDD.n3891 9.3005
R6696 VDD.n3893 VDD.n355 9.3005
R6697 VDD.n3895 VDD.n3894 9.3005
R6698 VDD.n345 VDD.n344 9.3005
R6699 VDD.n3908 VDD.n3907 9.3005
R6700 VDD.n3909 VDD.n343 9.3005
R6701 VDD.n3911 VDD.n3910 9.3005
R6702 VDD.n333 VDD.n332 9.3005
R6703 VDD.n3924 VDD.n3923 9.3005
R6704 VDD.n3925 VDD.n331 9.3005
R6705 VDD.n3927 VDD.n3926 9.3005
R6706 VDD.n321 VDD.n320 9.3005
R6707 VDD.n3943 VDD.n3942 9.3005
R6708 VDD.n3944 VDD.n319 9.3005
R6709 VDD.n3946 VDD.n3945 9.3005
R6710 VDD.n31 VDD.n29 9.3005
R6711 VDD.n464 VDD.n463 9.3005
R6712 VDD.n549 VDD.n548 9.3005
R6713 VDD.n550 VDD.n542 9.3005
R6714 VDD.n553 VDD.n541 9.3005
R6715 VDD.n554 VDD.n540 9.3005
R6716 VDD.n557 VDD.n539 9.3005
R6717 VDD.n558 VDD.n538 9.3005
R6718 VDD.n561 VDD.n537 9.3005
R6719 VDD.n562 VDD.n536 9.3005
R6720 VDD.n565 VDD.n535 9.3005
R6721 VDD.n566 VDD.n534 9.3005
R6722 VDD.n569 VDD.n533 9.3005
R6723 VDD.n570 VDD.n532 9.3005
R6724 VDD.n573 VDD.n531 9.3005
R6725 VDD.n574 VDD.n530 9.3005
R6726 VDD.n577 VDD.n529 9.3005
R6727 VDD.n578 VDD.n526 9.3005
R6728 VDD.n581 VDD.n525 9.3005
R6729 VDD.n582 VDD.n524 9.3005
R6730 VDD.n585 VDD.n523 9.3005
R6731 VDD.n586 VDD.n522 9.3005
R6732 VDD.n589 VDD.n521 9.3005
R6733 VDD.n590 VDD.n520 9.3005
R6734 VDD.n593 VDD.n519 9.3005
R6735 VDD.n594 VDD.n518 9.3005
R6736 VDD.n597 VDD.n517 9.3005
R6737 VDD.n598 VDD.n516 9.3005
R6738 VDD.n599 VDD.n515 9.3005
R6739 VDD.n498 VDD.n497 9.3005
R6740 VDD.n605 VDD.n604 9.3005
R6741 VDD.n544 VDD.n469 9.3005
R6742 VDD.n2568 VDD.n1242 9.3005
R6743 VDD.n2567 VDD.n2566 9.3005
R6744 VDD.n2565 VDD.n1246 9.3005
R6745 VDD.n2564 VDD.n2563 9.3005
R6746 VDD.n2562 VDD.n1247 9.3005
R6747 VDD.n2561 VDD.n2560 9.3005
R6748 VDD.n2559 VDD.n1251 9.3005
R6749 VDD.n2558 VDD.n2557 9.3005
R6750 VDD.n2556 VDD.n1252 9.3005
R6751 VDD.n2555 VDD.n2554 9.3005
R6752 VDD.n2553 VDD.n1256 9.3005
R6753 VDD.n2552 VDD.n2551 9.3005
R6754 VDD.n2550 VDD.n1257 9.3005
R6755 VDD.n2549 VDD.n2548 9.3005
R6756 VDD.n2547 VDD.n1263 9.3005
R6757 VDD.n2546 VDD.n2545 9.3005
R6758 VDD.n2544 VDD.n1264 9.3005
R6759 VDD.n2543 VDD.n2542 9.3005
R6760 VDD.n2541 VDD.n1268 9.3005
R6761 VDD.n2540 VDD.n2539 9.3005
R6762 VDD.n2538 VDD.n1269 9.3005
R6763 VDD.n2537 VDD.n2536 9.3005
R6764 VDD.n2535 VDD.n1273 9.3005
R6765 VDD.n2534 VDD.n2533 9.3005
R6766 VDD.n2532 VDD.n1274 9.3005
R6767 VDD.n2531 VDD.n2530 9.3005
R6768 VDD.n2529 VDD.n1278 9.3005
R6769 VDD.n2528 VDD.n2527 9.3005
R6770 VDD.n2525 VDD.n1279 9.3005
R6771 VDD.n2570 VDD.n2569 9.3005
R6772 VDD.n1741 VDD.n1740 9.3005
R6773 VDD.n1742 VDD.n1617 9.3005
R6774 VDD.n1744 VDD.n1743 9.3005
R6775 VDD.n1607 VDD.n1606 9.3005
R6776 VDD.n1757 VDD.n1756 9.3005
R6777 VDD.n1758 VDD.n1605 9.3005
R6778 VDD.n1760 VDD.n1759 9.3005
R6779 VDD.n1595 VDD.n1594 9.3005
R6780 VDD.n1773 VDD.n1772 9.3005
R6781 VDD.n1774 VDD.n1593 9.3005
R6782 VDD.n1776 VDD.n1775 9.3005
R6783 VDD.n1583 VDD.n1582 9.3005
R6784 VDD.n1789 VDD.n1788 9.3005
R6785 VDD.n1790 VDD.n1581 9.3005
R6786 VDD.n1792 VDD.n1791 9.3005
R6787 VDD.n1571 VDD.n1570 9.3005
R6788 VDD.n1805 VDD.n1804 9.3005
R6789 VDD.n1806 VDD.n1569 9.3005
R6790 VDD.n1808 VDD.n1807 9.3005
R6791 VDD.n1559 VDD.n1558 9.3005
R6792 VDD.n1821 VDD.n1820 9.3005
R6793 VDD.n1822 VDD.n1557 9.3005
R6794 VDD.n1824 VDD.n1823 9.3005
R6795 VDD.n1547 VDD.n1546 9.3005
R6796 VDD.n1837 VDD.n1836 9.3005
R6797 VDD.n1838 VDD.n1545 9.3005
R6798 VDD.n1840 VDD.n1839 9.3005
R6799 VDD.n1534 VDD.n1533 9.3005
R6800 VDD.n1853 VDD.n1852 9.3005
R6801 VDD.n1854 VDD.n1532 9.3005
R6802 VDD.n1856 VDD.n1855 9.3005
R6803 VDD.n1523 VDD.n1522 9.3005
R6804 VDD.n1869 VDD.n1868 9.3005
R6805 VDD.n1870 VDD.n1521 9.3005
R6806 VDD.n1872 VDD.n1871 9.3005
R6807 VDD.n1511 VDD.n1510 9.3005
R6808 VDD.n1885 VDD.n1884 9.3005
R6809 VDD.n1886 VDD.n1509 9.3005
R6810 VDD.n1888 VDD.n1887 9.3005
R6811 VDD.n1499 VDD.n1498 9.3005
R6812 VDD.n1901 VDD.n1900 9.3005
R6813 VDD.n1902 VDD.n1497 9.3005
R6814 VDD.n1904 VDD.n1903 9.3005
R6815 VDD.n1487 VDD.n1486 9.3005
R6816 VDD.n1917 VDD.n1916 9.3005
R6817 VDD.n1918 VDD.n1485 9.3005
R6818 VDD.n1920 VDD.n1919 9.3005
R6819 VDD.n1475 VDD.n1474 9.3005
R6820 VDD.n1933 VDD.n1932 9.3005
R6821 VDD.n1934 VDD.n1473 9.3005
R6822 VDD.n1936 VDD.n1935 9.3005
R6823 VDD.n1463 VDD.n1462 9.3005
R6824 VDD.n1962 VDD.n1961 9.3005
R6825 VDD.n1963 VDD.n1461 9.3005
R6826 VDD.n1965 VDD.n1964 9.3005
R6827 VDD.n1451 VDD.n1450 9.3005
R6828 VDD.n1978 VDD.n1977 9.3005
R6829 VDD.n1979 VDD.n1449 9.3005
R6830 VDD.n1981 VDD.n1980 9.3005
R6831 VDD.n1439 VDD.n1438 9.3005
R6832 VDD.n1994 VDD.n1993 9.3005
R6833 VDD.n1995 VDD.n1437 9.3005
R6834 VDD.n1997 VDD.n1996 9.3005
R6835 VDD.n1428 VDD.n1427 9.3005
R6836 VDD.n2011 VDD.n2010 9.3005
R6837 VDD.n2012 VDD.n1426 9.3005
R6838 VDD.n2014 VDD.n2013 9.3005
R6839 VDD.n1416 VDD.n1415 9.3005
R6840 VDD.n2027 VDD.n2026 9.3005
R6841 VDD.n2028 VDD.n1414 9.3005
R6842 VDD.n2030 VDD.n2029 9.3005
R6843 VDD.n1404 VDD.n1403 9.3005
R6844 VDD.n2043 VDD.n2042 9.3005
R6845 VDD.n2044 VDD.n1402 9.3005
R6846 VDD.n2046 VDD.n2045 9.3005
R6847 VDD.n1392 VDD.n1391 9.3005
R6848 VDD.n2059 VDD.n2058 9.3005
R6849 VDD.n2060 VDD.n1390 9.3005
R6850 VDD.n2062 VDD.n2061 9.3005
R6851 VDD.n1380 VDD.n1379 9.3005
R6852 VDD.n2075 VDD.n2074 9.3005
R6853 VDD.n2076 VDD.n1378 9.3005
R6854 VDD.n2078 VDD.n2077 9.3005
R6855 VDD.n1367 VDD.n1366 9.3005
R6856 VDD.n2091 VDD.n2090 9.3005
R6857 VDD.n2092 VDD.n1365 9.3005
R6858 VDD.n2094 VDD.n2093 9.3005
R6859 VDD.n1356 VDD.n1355 9.3005
R6860 VDD.n2107 VDD.n2106 9.3005
R6861 VDD.n2108 VDD.n1354 9.3005
R6862 VDD.n2110 VDD.n2109 9.3005
R6863 VDD.n1344 VDD.n1343 9.3005
R6864 VDD.n2123 VDD.n2122 9.3005
R6865 VDD.n2124 VDD.n1342 9.3005
R6866 VDD.n2126 VDD.n2125 9.3005
R6867 VDD.n1332 VDD.n1331 9.3005
R6868 VDD.n2139 VDD.n2138 9.3005
R6869 VDD.n2140 VDD.n1329 9.3005
R6870 VDD.n2143 VDD.n2142 9.3005
R6871 VDD.n2141 VDD.n1330 9.3005
R6872 VDD.n1320 VDD.n1319 9.3005
R6873 VDD.n2158 VDD.n2157 9.3005
R6874 VDD.n2159 VDD.n1317 9.3005
R6875 VDD.n2510 VDD.n2509 9.3005
R6876 VDD.n2508 VDD.n1318 9.3005
R6877 VDD.n2507 VDD.n1285 9.3005
R6878 VDD.n1619 VDD.n1618 9.3005
R6879 VDD.n1685 VDD.n1684 9.3005
R6880 VDD.n1686 VDD.n1677 9.3005
R6881 VDD.n1688 VDD.n1687 9.3005
R6882 VDD.n1689 VDD.n1672 9.3005
R6883 VDD.n1691 VDD.n1690 9.3005
R6884 VDD.n1692 VDD.n1671 9.3005
R6885 VDD.n1694 VDD.n1693 9.3005
R6886 VDD.n1695 VDD.n1666 9.3005
R6887 VDD.n1697 VDD.n1696 9.3005
R6888 VDD.n1698 VDD.n1665 9.3005
R6889 VDD.n1700 VDD.n1699 9.3005
R6890 VDD.n1701 VDD.n1660 9.3005
R6891 VDD.n1703 VDD.n1702 9.3005
R6892 VDD.n1704 VDD.n1659 9.3005
R6893 VDD.n1706 VDD.n1705 9.3005
R6894 VDD.n1710 VDD.n1655 9.3005
R6895 VDD.n1712 VDD.n1711 9.3005
R6896 VDD.n1713 VDD.n1654 9.3005
R6897 VDD.n1715 VDD.n1714 9.3005
R6898 VDD.n1716 VDD.n1649 9.3005
R6899 VDD.n1718 VDD.n1717 9.3005
R6900 VDD.n1719 VDD.n1648 9.3005
R6901 VDD.n1721 VDD.n1720 9.3005
R6902 VDD.n1722 VDD.n1643 9.3005
R6903 VDD.n1724 VDD.n1723 9.3005
R6904 VDD.n1725 VDD.n1642 9.3005
R6905 VDD.n1727 VDD.n1726 9.3005
R6906 VDD.n1625 VDD.n1624 9.3005
R6907 VDD.n1733 VDD.n1732 9.3005
R6908 VDD.n1680 VDD.n1678 9.3005
R6909 VDD.n1736 VDD.n1735 9.3005
R6910 VDD.n1613 VDD.n1612 9.3005
R6911 VDD.n1749 VDD.n1748 9.3005
R6912 VDD.n1750 VDD.n1611 9.3005
R6913 VDD.n1752 VDD.n1751 9.3005
R6914 VDD.n1601 VDD.n1600 9.3005
R6915 VDD.n1765 VDD.n1764 9.3005
R6916 VDD.n1766 VDD.n1599 9.3005
R6917 VDD.n1768 VDD.n1767 9.3005
R6918 VDD.n1589 VDD.n1588 9.3005
R6919 VDD.n1781 VDD.n1780 9.3005
R6920 VDD.n1782 VDD.n1587 9.3005
R6921 VDD.n1784 VDD.n1783 9.3005
R6922 VDD.n1577 VDD.n1576 9.3005
R6923 VDD.n1797 VDD.n1796 9.3005
R6924 VDD.n1798 VDD.n1575 9.3005
R6925 VDD.n1800 VDD.n1799 9.3005
R6926 VDD.n1565 VDD.n1564 9.3005
R6927 VDD.n1813 VDD.n1812 9.3005
R6928 VDD.n1814 VDD.n1563 9.3005
R6929 VDD.n1816 VDD.n1815 9.3005
R6930 VDD.n1553 VDD.n1552 9.3005
R6931 VDD.n1829 VDD.n1828 9.3005
R6932 VDD.n1830 VDD.n1551 9.3005
R6933 VDD.n1832 VDD.n1831 9.3005
R6934 VDD.n1541 VDD.n1540 9.3005
R6935 VDD.n1845 VDD.n1844 9.3005
R6936 VDD.n1846 VDD.n1539 9.3005
R6937 VDD.n1848 VDD.n1847 9.3005
R6938 VDD.n1529 VDD.n1528 9.3005
R6939 VDD.n1861 VDD.n1860 9.3005
R6940 VDD.n1862 VDD.n1527 9.3005
R6941 VDD.n1864 VDD.n1863 9.3005
R6942 VDD.n1517 VDD.n1516 9.3005
R6943 VDD.n1877 VDD.n1876 9.3005
R6944 VDD.n1878 VDD.n1515 9.3005
R6945 VDD.n1880 VDD.n1879 9.3005
R6946 VDD.n1505 VDD.n1504 9.3005
R6947 VDD.n1893 VDD.n1892 9.3005
R6948 VDD.n1894 VDD.n1503 9.3005
R6949 VDD.n1896 VDD.n1895 9.3005
R6950 VDD.n1493 VDD.n1492 9.3005
R6951 VDD.n1909 VDD.n1908 9.3005
R6952 VDD.n1910 VDD.n1491 9.3005
R6953 VDD.n1912 VDD.n1911 9.3005
R6954 VDD.n1481 VDD.n1480 9.3005
R6955 VDD.n1925 VDD.n1924 9.3005
R6956 VDD.n1926 VDD.n1479 9.3005
R6957 VDD.n1928 VDD.n1927 9.3005
R6958 VDD.n1469 VDD.n1468 9.3005
R6959 VDD.n1941 VDD.n1940 9.3005
R6960 VDD.n1942 VDD.n1467 9.3005
R6961 VDD.n1734 VDD.n1623 9.3005
R6962 VDD.n1958 VDD.n1957 9.3005
R6963 VDD.n1032 VDD.t0 9.25602
R6964 VDD.t61 VDD.n982 9.25602
R6965 VDD.n3349 VDD.t33 9.25602
R6966 VDD.n3391 VDD.t136 9.25602
R6967 VDD.n1537 VDD.t21 9.08138
R6968 VDD.t63 VDD.n1394 9.08138
R6969 VDD.n3856 VDD.t50 9.08138
R6970 VDD.n100 VDD.t5 9.08138
R6971 VDD.n1858 VDD.t21 8.38285
R6972 VDD.n2048 VDD.t63 8.38285
R6973 VDD.n3865 VDD.t50 8.38285
R6974 VDD.n4114 VDD.t5 8.38285
R6975 VDD.n15 VDD.n14 8.26895
R6976 VDD.n4159 VDD.n4158 8.19113
R6977 VDD.n1957 VDD.n1956 8.19113
R6978 VDD.n3165 VDD.n3164 7.96148
R6979 VDD.n3687 VDD.n3686 7.96148
R6980 VDD.n481 VDD.n476 7.96148
R6981 VDD.n3260 VDD.n3259 7.96148
R6982 VDD.n2868 VDD.n2867 7.96148
R6983 VDD.n2490 VDD.n2489 7.96148
R6984 VDD.n2931 VDD.n2930 7.96148
R6985 VDD.n2322 VDD.n2310 7.96148
R6986 VDD.n7 VDD.t13 7.92855
R6987 VDD.n7 VDD.t10 7.92855
R6988 VDD.n8 VDD.t20 7.92855
R6989 VDD.n8 VDD.t60 7.92855
R6990 VDD.n10 VDD.t137 7.92855
R6991 VDD.n10 VDD.t31 7.92855
R6992 VDD.n12 VDD.t41 7.92855
R6993 VDD.n12 VDD.t34 7.92855
R6994 VDD.n5 VDD.t62 7.92855
R6995 VDD.n5 VDD.t58 7.92855
R6996 VDD.n3 VDD.t135 7.92855
R6997 VDD.n3 VDD.t1 7.92855
R6998 VDD.n1 VDD.t131 7.92855
R6999 VDD.n1 VDD.t44 7.92855
R7000 VDD.n0 VDD.t29 7.92855
R7001 VDD.n0 VDD.t3 7.92855
R7002 VDD.n2468 VDD.t2 7.85896
R7003 VDD.n2751 VDD.t134 7.85896
R7004 VDD.n2859 VDD.t57 7.85896
R7005 VDD.n3239 VDD.t40 7.85896
R7006 VDD.n781 VDD.t30 7.85896
R7007 VDD.n3629 VDD.t12 7.85896
R7008 VDD.n1955 VDD.n1948 7.59102
R7009 VDD.n2697 VDD.t132 6.63653
R7010 VDD.n2775 VDD.t32 6.63653
R7011 VDD.n805 VDD.t15 6.63653
R7012 VDD.t4 VDD.n717 6.63653
R7013 VDD.n25 VDD.t18 6.60721
R7014 VDD.n25 VDD.t35 6.60721
R7015 VDD.n23 VDD.t48 6.60721
R7016 VDD.n23 VDD.t65 6.60721
R7017 VDD.n22 VDD.t39 6.60721
R7018 VDD.n22 VDD.t56 6.60721
R7019 VDD.n19 VDD.t49 6.60721
R7020 VDD.n19 VDD.t6 6.60721
R7021 VDD.n17 VDD.t66 6.60721
R7022 VDD.n17 VDD.t24 6.60721
R7023 VDD.n16 VDD.t38 6.60721
R7024 VDD.n16 VDD.t51 6.60721
R7025 VDD.n1949 VDD.t53 6.60721
R7026 VDD.n1949 VDD.t64 6.60721
R7027 VDD.n1951 VDD.t133 6.60721
R7028 VDD.n1951 VDD.t138 6.60721
R7029 VDD.n1953 VDD.t55 6.60721
R7030 VDD.n1953 VDD.t22 6.60721
R7031 VDD.n1943 VDD.t141 6.60721
R7032 VDD.n1943 VDD.t71 6.60721
R7033 VDD.n1945 VDD.t68 6.60721
R7034 VDD.n1945 VDD.t27 6.60721
R7035 VDD.n1947 VDD.t139 6.60721
R7036 VDD.n1947 VDD.t72 6.60721
R7037 VDD.n2691 VDD.t43 6.4619
R7038 VDD.t19 VDD.n711 6.4619
R7039 VDD.n28 VDD.n21 6.37981
R7040 VDD.n2468 VDD.t120 6.28726
R7041 VDD.n960 VDD.t74 6.28726
R7042 VDD.n3319 VDD.t90 6.28726
R7043 VDD.n3629 VDD.t78 6.28726
R7044 VDD.n1955 VDD.n1954 5.9186
R7045 VDD.n4159 VDD.n28 5.85499
R7046 VDD.n1956 VDD.n1955 5.85499
R7047 VDD.n2526 VDD.n2525 5.81868
R7048 VDD.n1683 VDD.n1680 5.81868
R7049 VDD.n547 VDD.n544 5.81868
R7050 VDD.n4047 VDD.n197 5.81868
R7051 VDD.n2613 VDD.t120 5.58874
R7052 VDD.n2859 VDD.t74 5.58874
R7053 VDD.n3239 VDD.t90 5.58874
R7054 VDD.t78 VDD.n633 5.58874
R7055 VDD.t43 VDD.n1113 5.4141
R7056 VDD.n3551 VDD.t19 5.4141
R7057 VDD.n3700 VDD.n607 5.30782
R7058 VDD.n609 VDD.n607 5.30782
R7059 VDD.n3738 VDD.n470 5.30782
R7060 VDD.n3738 VDD.n3737 5.30782
R7061 VDD.n2505 VDD.n2178 5.30782
R7062 VDD.n2505 VDD.n2504 5.30782
R7063 VDD.n2573 VDD.n2572 5.30782
R7064 VDD.n2572 VDD.n1240 5.30782
R7065 VDD.t132 VDD.n1107 5.23947
R7066 VDD.n1044 VDD.t32 5.23947
R7067 VDD.n3403 VDD.t15 5.23947
R7068 VDD.n3545 VDD.t4 5.23947
R7069 VDD.n1810 VDD.t54 4.89021
R7070 VDD.n2096 VDD.t69 4.89021
R7071 VDD.n3816 VDD.t37 4.89021
R7072 VDD.t7 VDD.n4090 4.89021
R7073 VDD.n28 VDD.n27 4.7074
R7074 VDD.t67 VDD.n1495 4.19168
R7075 VDD.n1999 VDD.t52 4.19168
R7076 VDD.t47 VDD.n341 4.19168
R7077 VDD.t17 VDD.n60 4.19168
R7078 VDD.n2619 VDD.t2 4.01704
R7079 VDD.n1068 VDD.t134 4.01704
R7080 VDD.t57 VDD.n945 4.01704
R7081 VDD.n3313 VDD.t40 4.01704
R7082 VDD.n3432 VDD.t30 4.01704
R7083 VDD.n647 VDD.t12 4.01704
R7084 VDD.n3166 VDD.n3165 2.65416
R7085 VDD.n3686 VDD.n3685 2.65416
R7086 VDD.n3723 VDD.n481 2.65416
R7087 VDD.n3259 VDD.n3258 2.65416
R7088 VDD.n2867 VDD.n2866 2.65416
R7089 VDD.n2489 VDD.n2488 2.65416
R7090 VDD.n2930 VDD.n2929 2.65416
R7091 VDD.n2325 VDD.n2310 2.65416
R7092 VDD.n2787 VDD.t0 2.61999
R7093 VDD.n2823 VDD.t61 2.61999
R7094 VDD.t33 VDD.n845 2.61999
R7095 VDD.n817 VDD.t136 2.61999
R7096 VDD.t86 VDD.n1603 2.44535
R7097 VDD.n2145 VDD.t82 2.44535
R7098 VDD.t94 VDD.n448 2.44535
R7099 VDD.t104 VDD.n159 2.44535
R7100 VDD.n26 VDD.n24 2.42291
R7101 VDD.n27 VDD.n26 2.42291
R7102 VDD.n20 VDD.n18 2.42291
R7103 VDD.n21 VDD.n20 2.42291
R7104 VDD.n1954 VDD.n1952 2.42291
R7105 VDD.n1952 VDD.n1950 2.42291
R7106 VDD.n1948 VDD.n1946 2.42291
R7107 VDD.n1946 VDD.n1944 2.42291
R7108 VDD.n1956 VDD.n15 2.32058
R7109 VDD VDD.n4159 2.31274
R7110 VDD.n4 VDD.n2 2.28929
R7111 VDD.n11 VDD.n9 2.28929
R7112 VDD.n6 VDD.n4 1.82378
R7113 VDD.n13 VDD.n11 1.82378
R7114 VDD.n14 VDD.n6 1.43369
R7115 VDD.n14 VDD.n13 1.43369
R7116 VDD.n2661 VDD.t36 1.39756
R7117 VDD.n2811 VDD.t14 1.39756
R7118 VDD.n841 VDD.t11 1.39756
R7119 VDD.t45 VDD.n681 1.39756
R7120 VDD.n2655 VDD.t130 1.22293
R7121 VDD.t59 VDD.n675 1.22293
R7122 VDD.n2527 VDD.n2526 0.776258
R7123 VDD.n1684 VDD.n1683 0.776258
R7124 VDD.n549 VDD.n547 0.776258
R7125 VDD.n285 VDD.n197 0.776258
R7126 VDD.n4046 VDD.n4045 0.486781
R7127 VDD.n217 VDD.n214 0.486781
R7128 VDD.n1678 VDD.n1618 0.486781
R7129 VDD.n1734 VDD.n1733 0.486781
R7130 VDD.n2571 VDD.n1241 0.254392
R7131 VDD.n606 VDD.n463 0.254392
R7132 VDD.n606 VDD.n605 0.22611
R7133 VDD.n3739 VDD.n469 0.22611
R7134 VDD.n2571 VDD.n2570 0.22611
R7135 VDD.n2506 VDD.n1279 0.22611
R7136 VDD.n3740 VDD.n3739 0.20691
R7137 VDD.n2507 VDD.n2506 0.20691
R7138 VDD.n1970 VDD.n1456 0.152939
R7139 VDD.n1971 VDD.n1970 0.152939
R7140 VDD.n1972 VDD.n1971 0.152939
R7141 VDD.n1972 VDD.n1444 0.152939
R7142 VDD.n1986 VDD.n1444 0.152939
R7143 VDD.n1987 VDD.n1986 0.152939
R7144 VDD.n1988 VDD.n1987 0.152939
R7145 VDD.n1988 VDD.n1432 0.152939
R7146 VDD.n2003 VDD.n1432 0.152939
R7147 VDD.n2004 VDD.n2003 0.152939
R7148 VDD.n2005 VDD.n2004 0.152939
R7149 VDD.n2005 VDD.n1421 0.152939
R7150 VDD.n2019 VDD.n1421 0.152939
R7151 VDD.n2020 VDD.n2019 0.152939
R7152 VDD.n2021 VDD.n2020 0.152939
R7153 VDD.n2021 VDD.n1409 0.152939
R7154 VDD.n2035 VDD.n1409 0.152939
R7155 VDD.n2036 VDD.n2035 0.152939
R7156 VDD.n2037 VDD.n2036 0.152939
R7157 VDD.n2037 VDD.n1397 0.152939
R7158 VDD.n2051 VDD.n1397 0.152939
R7159 VDD.n2052 VDD.n2051 0.152939
R7160 VDD.n2053 VDD.n2052 0.152939
R7161 VDD.n2053 VDD.n1385 0.152939
R7162 VDD.n2067 VDD.n1385 0.152939
R7163 VDD.n2068 VDD.n2067 0.152939
R7164 VDD.n2069 VDD.n2068 0.152939
R7165 VDD.n2069 VDD.n1373 0.152939
R7166 VDD.n2083 VDD.n1373 0.152939
R7167 VDD.n2084 VDD.n2083 0.152939
R7168 VDD.n2085 VDD.n2084 0.152939
R7169 VDD.n2085 VDD.n1361 0.152939
R7170 VDD.n2099 VDD.n1361 0.152939
R7171 VDD.n2100 VDD.n2099 0.152939
R7172 VDD.n2101 VDD.n2100 0.152939
R7173 VDD.n2101 VDD.n1349 0.152939
R7174 VDD.n2115 VDD.n1349 0.152939
R7175 VDD.n2116 VDD.n2115 0.152939
R7176 VDD.n2117 VDD.n2116 0.152939
R7177 VDD.n2117 VDD.n1337 0.152939
R7178 VDD.n2131 VDD.n1337 0.152939
R7179 VDD.n2132 VDD.n2131 0.152939
R7180 VDD.n2133 VDD.n2132 0.152939
R7181 VDD.n2133 VDD.n1324 0.152939
R7182 VDD.n2149 VDD.n1324 0.152939
R7183 VDD.n2150 VDD.n2149 0.152939
R7184 VDD.n2151 VDD.n2150 0.152939
R7185 VDD.n2151 VDD.n1311 0.152939
R7186 VDD.n2516 VDD.n1311 0.152939
R7187 VDD.n2517 VDD.n2516 0.152939
R7188 VDD.n2518 VDD.n2517 0.152939
R7189 VDD.n2518 VDD.n1241 0.152939
R7190 VDD.n3741 VDD.n3740 0.152939
R7191 VDD.n3741 VDD.n457 0.152939
R7192 VDD.n3755 VDD.n457 0.152939
R7193 VDD.n3756 VDD.n3755 0.152939
R7194 VDD.n3757 VDD.n3756 0.152939
R7195 VDD.n3757 VDD.n445 0.152939
R7196 VDD.n3771 VDD.n445 0.152939
R7197 VDD.n3772 VDD.n3771 0.152939
R7198 VDD.n3773 VDD.n3772 0.152939
R7199 VDD.n3773 VDD.n433 0.152939
R7200 VDD.n3787 VDD.n433 0.152939
R7201 VDD.n3788 VDD.n3787 0.152939
R7202 VDD.n3789 VDD.n3788 0.152939
R7203 VDD.n3789 VDD.n421 0.152939
R7204 VDD.n3803 VDD.n421 0.152939
R7205 VDD.n3804 VDD.n3803 0.152939
R7206 VDD.n3805 VDD.n3804 0.152939
R7207 VDD.n3805 VDD.n409 0.152939
R7208 VDD.n3819 VDD.n409 0.152939
R7209 VDD.n3820 VDD.n3819 0.152939
R7210 VDD.n3821 VDD.n3820 0.152939
R7211 VDD.n3821 VDD.n397 0.152939
R7212 VDD.n3835 VDD.n397 0.152939
R7213 VDD.n3836 VDD.n3835 0.152939
R7214 VDD.n3837 VDD.n3836 0.152939
R7215 VDD.n3837 VDD.n385 0.152939
R7216 VDD.n3851 VDD.n385 0.152939
R7217 VDD.n3852 VDD.n3851 0.152939
R7218 VDD.n3853 VDD.n3852 0.152939
R7219 VDD.n3853 VDD.n374 0.152939
R7220 VDD.n3868 VDD.n374 0.152939
R7221 VDD.n3869 VDD.n3868 0.152939
R7222 VDD.n3870 VDD.n3869 0.152939
R7223 VDD.n3870 VDD.n362 0.152939
R7224 VDD.n3884 VDD.n362 0.152939
R7225 VDD.n3885 VDD.n3884 0.152939
R7226 VDD.n3886 VDD.n3885 0.152939
R7227 VDD.n3886 VDD.n350 0.152939
R7228 VDD.n3900 VDD.n350 0.152939
R7229 VDD.n3901 VDD.n3900 0.152939
R7230 VDD.n3902 VDD.n3901 0.152939
R7231 VDD.n3902 VDD.n338 0.152939
R7232 VDD.n3916 VDD.n338 0.152939
R7233 VDD.n3917 VDD.n3916 0.152939
R7234 VDD.n3918 VDD.n3917 0.152939
R7235 VDD.n3918 VDD.n326 0.152939
R7236 VDD.n3932 VDD.n326 0.152939
R7237 VDD.n3933 VDD.n3932 0.152939
R7238 VDD.n3934 VDD.n3933 0.152939
R7239 VDD.n3936 VDD.n3934 0.152939
R7240 VDD.n3936 VDD.n3935 0.152939
R7241 VDD.n3935 VDD.n315 0.152939
R7242 VDD.n315 VDD.n313 0.152939
R7243 VDD.n3954 VDD.n313 0.152939
R7244 VDD.n3955 VDD.n3954 0.152939
R7245 VDD.n3956 VDD.n3955 0.152939
R7246 VDD.n3956 VDD.n311 0.152939
R7247 VDD.n3961 VDD.n311 0.152939
R7248 VDD.n3962 VDD.n3961 0.152939
R7249 VDD.n3963 VDD.n3962 0.152939
R7250 VDD.n3963 VDD.n309 0.152939
R7251 VDD.n3968 VDD.n309 0.152939
R7252 VDD.n3969 VDD.n3968 0.152939
R7253 VDD.n3970 VDD.n3969 0.152939
R7254 VDD.n3970 VDD.n307 0.152939
R7255 VDD.n3975 VDD.n307 0.152939
R7256 VDD.n3976 VDD.n3975 0.152939
R7257 VDD.n3977 VDD.n3976 0.152939
R7258 VDD.n3977 VDD.n305 0.152939
R7259 VDD.n3982 VDD.n305 0.152939
R7260 VDD.n3983 VDD.n3982 0.152939
R7261 VDD.n3984 VDD.n3983 0.152939
R7262 VDD.n3984 VDD.n303 0.152939
R7263 VDD.n3989 VDD.n303 0.152939
R7264 VDD.n3990 VDD.n3989 0.152939
R7265 VDD.n3991 VDD.n3990 0.152939
R7266 VDD.n3991 VDD.n301 0.152939
R7267 VDD.n3996 VDD.n301 0.152939
R7268 VDD.n3997 VDD.n3996 0.152939
R7269 VDD.n3998 VDD.n3997 0.152939
R7270 VDD.n3998 VDD.n299 0.152939
R7271 VDD.n4003 VDD.n299 0.152939
R7272 VDD.n4004 VDD.n4003 0.152939
R7273 VDD.n4005 VDD.n4004 0.152939
R7274 VDD.n4005 VDD.n297 0.152939
R7275 VDD.n4010 VDD.n297 0.152939
R7276 VDD.n4011 VDD.n4010 0.152939
R7277 VDD.n4012 VDD.n4011 0.152939
R7278 VDD.n4012 VDD.n295 0.152939
R7279 VDD.n4017 VDD.n295 0.152939
R7280 VDD.n4018 VDD.n4017 0.152939
R7281 VDD.n4019 VDD.n4018 0.152939
R7282 VDD.n4019 VDD.n293 0.152939
R7283 VDD.n4024 VDD.n293 0.152939
R7284 VDD.n4025 VDD.n4024 0.152939
R7285 VDD.n4026 VDD.n4025 0.152939
R7286 VDD.n4026 VDD.n291 0.152939
R7287 VDD.n4031 VDD.n291 0.152939
R7288 VDD.n4032 VDD.n4031 0.152939
R7289 VDD.n4033 VDD.n4032 0.152939
R7290 VDD.n4033 VDD.n289 0.152939
R7291 VDD.n4038 VDD.n289 0.152939
R7292 VDD.n4039 VDD.n4038 0.152939
R7293 VDD.n4040 VDD.n4039 0.152939
R7294 VDD.n4040 VDD.n287 0.152939
R7295 VDD.n4045 VDD.n287 0.152939
R7296 VDD.n218 VDD.n217 0.152939
R7297 VDD.n219 VDD.n218 0.152939
R7298 VDD.n219 VDD.n212 0.152939
R7299 VDD.n227 VDD.n212 0.152939
R7300 VDD.n228 VDD.n227 0.152939
R7301 VDD.n229 VDD.n228 0.152939
R7302 VDD.n229 VDD.n210 0.152939
R7303 VDD.n237 VDD.n210 0.152939
R7304 VDD.n238 VDD.n237 0.152939
R7305 VDD.n239 VDD.n238 0.152939
R7306 VDD.n239 VDD.n208 0.152939
R7307 VDD.n247 VDD.n208 0.152939
R7308 VDD.n248 VDD.n247 0.152939
R7309 VDD.n249 VDD.n248 0.152939
R7310 VDD.n249 VDD.n204 0.152939
R7311 VDD.n257 VDD.n204 0.152939
R7312 VDD.n258 VDD.n257 0.152939
R7313 VDD.n259 VDD.n258 0.152939
R7314 VDD.n259 VDD.n202 0.152939
R7315 VDD.n267 VDD.n202 0.152939
R7316 VDD.n268 VDD.n267 0.152939
R7317 VDD.n269 VDD.n268 0.152939
R7318 VDD.n269 VDD.n200 0.152939
R7319 VDD.n277 VDD.n200 0.152939
R7320 VDD.n278 VDD.n277 0.152939
R7321 VDD.n279 VDD.n278 0.152939
R7322 VDD.n279 VDD.n198 0.152939
R7323 VDD.n286 VDD.n198 0.152939
R7324 VDD.n4046 VDD.n286 0.152939
R7325 VDD.n41 VDD.n30 0.152939
R7326 VDD.n42 VDD.n41 0.152939
R7327 VDD.n43 VDD.n42 0.152939
R7328 VDD.n51 VDD.n43 0.152939
R7329 VDD.n52 VDD.n51 0.152939
R7330 VDD.n53 VDD.n52 0.152939
R7331 VDD.n54 VDD.n53 0.152939
R7332 VDD.n62 VDD.n54 0.152939
R7333 VDD.n63 VDD.n62 0.152939
R7334 VDD.n64 VDD.n63 0.152939
R7335 VDD.n65 VDD.n64 0.152939
R7336 VDD.n73 VDD.n65 0.152939
R7337 VDD.n74 VDD.n73 0.152939
R7338 VDD.n75 VDD.n74 0.152939
R7339 VDD.n76 VDD.n75 0.152939
R7340 VDD.n84 VDD.n76 0.152939
R7341 VDD.n85 VDD.n84 0.152939
R7342 VDD.n86 VDD.n85 0.152939
R7343 VDD.n87 VDD.n86 0.152939
R7344 VDD.n94 VDD.n87 0.152939
R7345 VDD.n95 VDD.n94 0.152939
R7346 VDD.n96 VDD.n95 0.152939
R7347 VDD.n97 VDD.n96 0.152939
R7348 VDD.n106 VDD.n97 0.152939
R7349 VDD.n107 VDD.n106 0.152939
R7350 VDD.n108 VDD.n107 0.152939
R7351 VDD.n109 VDD.n108 0.152939
R7352 VDD.n117 VDD.n109 0.152939
R7353 VDD.n118 VDD.n117 0.152939
R7354 VDD.n119 VDD.n118 0.152939
R7355 VDD.n120 VDD.n119 0.152939
R7356 VDD.n128 VDD.n120 0.152939
R7357 VDD.n129 VDD.n128 0.152939
R7358 VDD.n130 VDD.n129 0.152939
R7359 VDD.n131 VDD.n130 0.152939
R7360 VDD.n139 VDD.n131 0.152939
R7361 VDD.n140 VDD.n139 0.152939
R7362 VDD.n141 VDD.n140 0.152939
R7363 VDD.n142 VDD.n141 0.152939
R7364 VDD.n150 VDD.n142 0.152939
R7365 VDD.n151 VDD.n150 0.152939
R7366 VDD.n152 VDD.n151 0.152939
R7367 VDD.n153 VDD.n152 0.152939
R7368 VDD.n161 VDD.n153 0.152939
R7369 VDD.n162 VDD.n161 0.152939
R7370 VDD.n163 VDD.n162 0.152939
R7371 VDD.n164 VDD.n163 0.152939
R7372 VDD.n172 VDD.n164 0.152939
R7373 VDD.n173 VDD.n172 0.152939
R7374 VDD.n174 VDD.n173 0.152939
R7375 VDD.n175 VDD.n174 0.152939
R7376 VDD.n214 VDD.n175 0.152939
R7377 VDD.n3747 VDD.n463 0.152939
R7378 VDD.n3748 VDD.n3747 0.152939
R7379 VDD.n3749 VDD.n3748 0.152939
R7380 VDD.n3749 VDD.n451 0.152939
R7381 VDD.n3763 VDD.n451 0.152939
R7382 VDD.n3764 VDD.n3763 0.152939
R7383 VDD.n3765 VDD.n3764 0.152939
R7384 VDD.n3765 VDD.n439 0.152939
R7385 VDD.n3779 VDD.n439 0.152939
R7386 VDD.n3780 VDD.n3779 0.152939
R7387 VDD.n3781 VDD.n3780 0.152939
R7388 VDD.n3781 VDD.n427 0.152939
R7389 VDD.n3795 VDD.n427 0.152939
R7390 VDD.n3796 VDD.n3795 0.152939
R7391 VDD.n3797 VDD.n3796 0.152939
R7392 VDD.n3797 VDD.n415 0.152939
R7393 VDD.n3811 VDD.n415 0.152939
R7394 VDD.n3812 VDD.n3811 0.152939
R7395 VDD.n3813 VDD.n3812 0.152939
R7396 VDD.n3813 VDD.n403 0.152939
R7397 VDD.n3827 VDD.n403 0.152939
R7398 VDD.n3828 VDD.n3827 0.152939
R7399 VDD.n3829 VDD.n3828 0.152939
R7400 VDD.n3829 VDD.n391 0.152939
R7401 VDD.n3843 VDD.n391 0.152939
R7402 VDD.n3844 VDD.n3843 0.152939
R7403 VDD.n3845 VDD.n3844 0.152939
R7404 VDD.n3845 VDD.n379 0.152939
R7405 VDD.n3860 VDD.n379 0.152939
R7406 VDD.n3861 VDD.n3860 0.152939
R7407 VDD.n3862 VDD.n3861 0.152939
R7408 VDD.n3862 VDD.n368 0.152939
R7409 VDD.n3876 VDD.n368 0.152939
R7410 VDD.n3877 VDD.n3876 0.152939
R7411 VDD.n3878 VDD.n3877 0.152939
R7412 VDD.n3878 VDD.n356 0.152939
R7413 VDD.n3892 VDD.n356 0.152939
R7414 VDD.n3893 VDD.n3892 0.152939
R7415 VDD.n3894 VDD.n3893 0.152939
R7416 VDD.n3894 VDD.n344 0.152939
R7417 VDD.n3908 VDD.n344 0.152939
R7418 VDD.n3909 VDD.n3908 0.152939
R7419 VDD.n3910 VDD.n3909 0.152939
R7420 VDD.n3910 VDD.n332 0.152939
R7421 VDD.n3924 VDD.n332 0.152939
R7422 VDD.n3925 VDD.n3924 0.152939
R7423 VDD.n3926 VDD.n3925 0.152939
R7424 VDD.n3926 VDD.n320 0.152939
R7425 VDD.n3943 VDD.n320 0.152939
R7426 VDD.n3944 VDD.n3943 0.152939
R7427 VDD.n3945 VDD.n3944 0.152939
R7428 VDD.n3945 VDD.n29 0.152939
R7429 VDD.n605 VDD.n497 0.152939
R7430 VDD.n515 VDD.n497 0.152939
R7431 VDD.n516 VDD.n515 0.152939
R7432 VDD.n517 VDD.n516 0.152939
R7433 VDD.n518 VDD.n517 0.152939
R7434 VDD.n519 VDD.n518 0.152939
R7435 VDD.n520 VDD.n519 0.152939
R7436 VDD.n521 VDD.n520 0.152939
R7437 VDD.n522 VDD.n521 0.152939
R7438 VDD.n523 VDD.n522 0.152939
R7439 VDD.n524 VDD.n523 0.152939
R7440 VDD.n525 VDD.n524 0.152939
R7441 VDD.n526 VDD.n525 0.152939
R7442 VDD.n529 VDD.n526 0.152939
R7443 VDD.n530 VDD.n529 0.152939
R7444 VDD.n531 VDD.n530 0.152939
R7445 VDD.n532 VDD.n531 0.152939
R7446 VDD.n533 VDD.n532 0.152939
R7447 VDD.n534 VDD.n533 0.152939
R7448 VDD.n535 VDD.n534 0.152939
R7449 VDD.n536 VDD.n535 0.152939
R7450 VDD.n537 VDD.n536 0.152939
R7451 VDD.n538 VDD.n537 0.152939
R7452 VDD.n539 VDD.n538 0.152939
R7453 VDD.n540 VDD.n539 0.152939
R7454 VDD.n541 VDD.n540 0.152939
R7455 VDD.n542 VDD.n541 0.152939
R7456 VDD.n548 VDD.n542 0.152939
R7457 VDD.n548 VDD.n469 0.152939
R7458 VDD.n2570 VDD.n1242 0.152939
R7459 VDD.n2566 VDD.n1242 0.152939
R7460 VDD.n2566 VDD.n2565 0.152939
R7461 VDD.n2565 VDD.n2564 0.152939
R7462 VDD.n2564 VDD.n1247 0.152939
R7463 VDD.n2560 VDD.n1247 0.152939
R7464 VDD.n2560 VDD.n2559 0.152939
R7465 VDD.n2559 VDD.n2558 0.152939
R7466 VDD.n2558 VDD.n1252 0.152939
R7467 VDD.n2554 VDD.n1252 0.152939
R7468 VDD.n2554 VDD.n2553 0.152939
R7469 VDD.n2553 VDD.n2552 0.152939
R7470 VDD.n2552 VDD.n1257 0.152939
R7471 VDD.n2548 VDD.n1257 0.152939
R7472 VDD.n2548 VDD.n2547 0.152939
R7473 VDD.n2547 VDD.n2546 0.152939
R7474 VDD.n2546 VDD.n1264 0.152939
R7475 VDD.n2542 VDD.n1264 0.152939
R7476 VDD.n2542 VDD.n2541 0.152939
R7477 VDD.n2541 VDD.n2540 0.152939
R7478 VDD.n2540 VDD.n1269 0.152939
R7479 VDD.n2536 VDD.n1269 0.152939
R7480 VDD.n2536 VDD.n2535 0.152939
R7481 VDD.n2535 VDD.n2534 0.152939
R7482 VDD.n2534 VDD.n1274 0.152939
R7483 VDD.n2530 VDD.n1274 0.152939
R7484 VDD.n2530 VDD.n2529 0.152939
R7485 VDD.n2529 VDD.n2528 0.152939
R7486 VDD.n2528 VDD.n1279 0.152939
R7487 VDD.n1741 VDD.n1618 0.152939
R7488 VDD.n1742 VDD.n1741 0.152939
R7489 VDD.n1743 VDD.n1742 0.152939
R7490 VDD.n1743 VDD.n1606 0.152939
R7491 VDD.n1757 VDD.n1606 0.152939
R7492 VDD.n1758 VDD.n1757 0.152939
R7493 VDD.n1759 VDD.n1758 0.152939
R7494 VDD.n1759 VDD.n1594 0.152939
R7495 VDD.n1773 VDD.n1594 0.152939
R7496 VDD.n1774 VDD.n1773 0.152939
R7497 VDD.n1775 VDD.n1774 0.152939
R7498 VDD.n1775 VDD.n1582 0.152939
R7499 VDD.n1789 VDD.n1582 0.152939
R7500 VDD.n1790 VDD.n1789 0.152939
R7501 VDD.n1791 VDD.n1790 0.152939
R7502 VDD.n1791 VDD.n1570 0.152939
R7503 VDD.n1805 VDD.n1570 0.152939
R7504 VDD.n1806 VDD.n1805 0.152939
R7505 VDD.n1807 VDD.n1806 0.152939
R7506 VDD.n1807 VDD.n1558 0.152939
R7507 VDD.n1821 VDD.n1558 0.152939
R7508 VDD.n1822 VDD.n1821 0.152939
R7509 VDD.n1823 VDD.n1822 0.152939
R7510 VDD.n1823 VDD.n1546 0.152939
R7511 VDD.n1837 VDD.n1546 0.152939
R7512 VDD.n1838 VDD.n1837 0.152939
R7513 VDD.n1839 VDD.n1838 0.152939
R7514 VDD.n1839 VDD.n1533 0.152939
R7515 VDD.n1853 VDD.n1533 0.152939
R7516 VDD.n1854 VDD.n1853 0.152939
R7517 VDD.n1855 VDD.n1854 0.152939
R7518 VDD.n1855 VDD.n1522 0.152939
R7519 VDD.n1869 VDD.n1522 0.152939
R7520 VDD.n1870 VDD.n1869 0.152939
R7521 VDD.n1871 VDD.n1870 0.152939
R7522 VDD.n1871 VDD.n1510 0.152939
R7523 VDD.n1885 VDD.n1510 0.152939
R7524 VDD.n1886 VDD.n1885 0.152939
R7525 VDD.n1887 VDD.n1886 0.152939
R7526 VDD.n1887 VDD.n1498 0.152939
R7527 VDD.n1901 VDD.n1498 0.152939
R7528 VDD.n1902 VDD.n1901 0.152939
R7529 VDD.n1903 VDD.n1902 0.152939
R7530 VDD.n1903 VDD.n1486 0.152939
R7531 VDD.n1917 VDD.n1486 0.152939
R7532 VDD.n1918 VDD.n1917 0.152939
R7533 VDD.n1919 VDD.n1918 0.152939
R7534 VDD.n1919 VDD.n1474 0.152939
R7535 VDD.n1933 VDD.n1474 0.152939
R7536 VDD.n1934 VDD.n1933 0.152939
R7537 VDD.n1935 VDD.n1934 0.152939
R7538 VDD.n1935 VDD.n1462 0.152939
R7539 VDD.n1962 VDD.n1462 0.152939
R7540 VDD.n1963 VDD.n1962 0.152939
R7541 VDD.n1964 VDD.n1963 0.152939
R7542 VDD.n1964 VDD.n1450 0.152939
R7543 VDD.n1978 VDD.n1450 0.152939
R7544 VDD.n1979 VDD.n1978 0.152939
R7545 VDD.n1980 VDD.n1979 0.152939
R7546 VDD.n1980 VDD.n1438 0.152939
R7547 VDD.n1994 VDD.n1438 0.152939
R7548 VDD.n1995 VDD.n1994 0.152939
R7549 VDD.n1996 VDD.n1995 0.152939
R7550 VDD.n1996 VDD.n1427 0.152939
R7551 VDD.n2011 VDD.n1427 0.152939
R7552 VDD.n2012 VDD.n2011 0.152939
R7553 VDD.n2013 VDD.n2012 0.152939
R7554 VDD.n2013 VDD.n1415 0.152939
R7555 VDD.n2027 VDD.n1415 0.152939
R7556 VDD.n2028 VDD.n2027 0.152939
R7557 VDD.n2029 VDD.n2028 0.152939
R7558 VDD.n2029 VDD.n1403 0.152939
R7559 VDD.n2043 VDD.n1403 0.152939
R7560 VDD.n2044 VDD.n2043 0.152939
R7561 VDD.n2045 VDD.n2044 0.152939
R7562 VDD.n2045 VDD.n1391 0.152939
R7563 VDD.n2059 VDD.n1391 0.152939
R7564 VDD.n2060 VDD.n2059 0.152939
R7565 VDD.n2061 VDD.n2060 0.152939
R7566 VDD.n2061 VDD.n1379 0.152939
R7567 VDD.n2075 VDD.n1379 0.152939
R7568 VDD.n2076 VDD.n2075 0.152939
R7569 VDD.n2077 VDD.n2076 0.152939
R7570 VDD.n2077 VDD.n1366 0.152939
R7571 VDD.n2091 VDD.n1366 0.152939
R7572 VDD.n2092 VDD.n2091 0.152939
R7573 VDD.n2093 VDD.n2092 0.152939
R7574 VDD.n2093 VDD.n1355 0.152939
R7575 VDD.n2107 VDD.n1355 0.152939
R7576 VDD.n2108 VDD.n2107 0.152939
R7577 VDD.n2109 VDD.n2108 0.152939
R7578 VDD.n2109 VDD.n1343 0.152939
R7579 VDD.n2123 VDD.n1343 0.152939
R7580 VDD.n2124 VDD.n2123 0.152939
R7581 VDD.n2125 VDD.n2124 0.152939
R7582 VDD.n2125 VDD.n1331 0.152939
R7583 VDD.n2139 VDD.n1331 0.152939
R7584 VDD.n2140 VDD.n2139 0.152939
R7585 VDD.n2142 VDD.n2140 0.152939
R7586 VDD.n2142 VDD.n2141 0.152939
R7587 VDD.n2141 VDD.n1319 0.152939
R7588 VDD.n2158 VDD.n1319 0.152939
R7589 VDD.n2159 VDD.n2158 0.152939
R7590 VDD.n2509 VDD.n2159 0.152939
R7591 VDD.n2509 VDD.n2508 0.152939
R7592 VDD.n2508 VDD.n2507 0.152939
R7593 VDD.n1733 VDD.n1624 0.152939
R7594 VDD.n1726 VDD.n1624 0.152939
R7595 VDD.n1726 VDD.n1725 0.152939
R7596 VDD.n1725 VDD.n1724 0.152939
R7597 VDD.n1724 VDD.n1643 0.152939
R7598 VDD.n1720 VDD.n1643 0.152939
R7599 VDD.n1720 VDD.n1719 0.152939
R7600 VDD.n1719 VDD.n1718 0.152939
R7601 VDD.n1718 VDD.n1649 0.152939
R7602 VDD.n1714 VDD.n1649 0.152939
R7603 VDD.n1714 VDD.n1713 0.152939
R7604 VDD.n1713 VDD.n1712 0.152939
R7605 VDD.n1712 VDD.n1655 0.152939
R7606 VDD.n1705 VDD.n1655 0.152939
R7607 VDD.n1705 VDD.n1704 0.152939
R7608 VDD.n1704 VDD.n1703 0.152939
R7609 VDD.n1703 VDD.n1660 0.152939
R7610 VDD.n1699 VDD.n1660 0.152939
R7611 VDD.n1699 VDD.n1698 0.152939
R7612 VDD.n1698 VDD.n1697 0.152939
R7613 VDD.n1697 VDD.n1666 0.152939
R7614 VDD.n1693 VDD.n1666 0.152939
R7615 VDD.n1693 VDD.n1692 0.152939
R7616 VDD.n1692 VDD.n1691 0.152939
R7617 VDD.n1691 VDD.n1672 0.152939
R7618 VDD.n1687 VDD.n1672 0.152939
R7619 VDD.n1687 VDD.n1686 0.152939
R7620 VDD.n1686 VDD.n1685 0.152939
R7621 VDD.n1685 VDD.n1678 0.152939
R7622 VDD.n1735 VDD.n1734 0.152939
R7623 VDD.n1735 VDD.n1612 0.152939
R7624 VDD.n1749 VDD.n1612 0.152939
R7625 VDD.n1750 VDD.n1749 0.152939
R7626 VDD.n1751 VDD.n1750 0.152939
R7627 VDD.n1751 VDD.n1600 0.152939
R7628 VDD.n1765 VDD.n1600 0.152939
R7629 VDD.n1766 VDD.n1765 0.152939
R7630 VDD.n1767 VDD.n1766 0.152939
R7631 VDD.n1767 VDD.n1588 0.152939
R7632 VDD.n1781 VDD.n1588 0.152939
R7633 VDD.n1782 VDD.n1781 0.152939
R7634 VDD.n1783 VDD.n1782 0.152939
R7635 VDD.n1783 VDD.n1576 0.152939
R7636 VDD.n1797 VDD.n1576 0.152939
R7637 VDD.n1798 VDD.n1797 0.152939
R7638 VDD.n1799 VDD.n1798 0.152939
R7639 VDD.n1799 VDD.n1564 0.152939
R7640 VDD.n1813 VDD.n1564 0.152939
R7641 VDD.n1814 VDD.n1813 0.152939
R7642 VDD.n1815 VDD.n1814 0.152939
R7643 VDD.n1815 VDD.n1552 0.152939
R7644 VDD.n1829 VDD.n1552 0.152939
R7645 VDD.n1830 VDD.n1829 0.152939
R7646 VDD.n1831 VDD.n1830 0.152939
R7647 VDD.n1831 VDD.n1540 0.152939
R7648 VDD.n1845 VDD.n1540 0.152939
R7649 VDD.n1846 VDD.n1845 0.152939
R7650 VDD.n1847 VDD.n1846 0.152939
R7651 VDD.n1847 VDD.n1528 0.152939
R7652 VDD.n1861 VDD.n1528 0.152939
R7653 VDD.n1862 VDD.n1861 0.152939
R7654 VDD.n1863 VDD.n1862 0.152939
R7655 VDD.n1863 VDD.n1516 0.152939
R7656 VDD.n1877 VDD.n1516 0.152939
R7657 VDD.n1878 VDD.n1877 0.152939
R7658 VDD.n1879 VDD.n1878 0.152939
R7659 VDD.n1879 VDD.n1504 0.152939
R7660 VDD.n1893 VDD.n1504 0.152939
R7661 VDD.n1894 VDD.n1893 0.152939
R7662 VDD.n1895 VDD.n1894 0.152939
R7663 VDD.n1895 VDD.n1492 0.152939
R7664 VDD.n1909 VDD.n1492 0.152939
R7665 VDD.n1910 VDD.n1909 0.152939
R7666 VDD.n1911 VDD.n1910 0.152939
R7667 VDD.n1911 VDD.n1480 0.152939
R7668 VDD.n1925 VDD.n1480 0.152939
R7669 VDD.n1926 VDD.n1925 0.152939
R7670 VDD.n1927 VDD.n1926 0.152939
R7671 VDD.n1927 VDD.n1468 0.152939
R7672 VDD.n1941 VDD.n1468 0.152939
R7673 VDD.n1942 VDD.n1941 0.152939
R7674 VDD.n1957 VDD.n1456 0.145814
R7675 VDD.n4158 VDD.n30 0.145814
R7676 VDD.n4158 VDD.n29 0.145814
R7677 VDD.n1957 VDD.n1942 0.145814
R7678 VDD VDD.n15 0.00833333
R7679 CS_BIAS.n324 CS_BIAS.n220 161.3
R7680 CS_BIAS.n323 CS_BIAS.n322 161.3
R7681 CS_BIAS.n321 CS_BIAS.n221 161.3
R7682 CS_BIAS.n320 CS_BIAS.n319 161.3
R7683 CS_BIAS.n318 CS_BIAS.n222 161.3
R7684 CS_BIAS.n317 CS_BIAS.n316 161.3
R7685 CS_BIAS.n315 CS_BIAS.n223 161.3
R7686 CS_BIAS.n314 CS_BIAS.n313 161.3
R7687 CS_BIAS.n312 CS_BIAS.n224 161.3
R7688 CS_BIAS.n311 CS_BIAS.n310 161.3
R7689 CS_BIAS.n309 CS_BIAS.n225 161.3
R7690 CS_BIAS.n308 CS_BIAS.n307 161.3
R7691 CS_BIAS.n305 CS_BIAS.n226 161.3
R7692 CS_BIAS.n304 CS_BIAS.n303 161.3
R7693 CS_BIAS.n302 CS_BIAS.n227 161.3
R7694 CS_BIAS.n301 CS_BIAS.n300 161.3
R7695 CS_BIAS.n299 CS_BIAS.n228 161.3
R7696 CS_BIAS.n298 CS_BIAS.n297 161.3
R7697 CS_BIAS.n296 CS_BIAS.n229 161.3
R7698 CS_BIAS.n295 CS_BIAS.n294 161.3
R7699 CS_BIAS.n293 CS_BIAS.n230 161.3
R7700 CS_BIAS.n292 CS_BIAS.n291 161.3
R7701 CS_BIAS.n290 CS_BIAS.n231 161.3
R7702 CS_BIAS.n289 CS_BIAS.n288 161.3
R7703 CS_BIAS.n287 CS_BIAS.n232 161.3
R7704 CS_BIAS.n285 CS_BIAS.n284 161.3
R7705 CS_BIAS.n283 CS_BIAS.n233 161.3
R7706 CS_BIAS.n282 CS_BIAS.n281 161.3
R7707 CS_BIAS.n280 CS_BIAS.n234 161.3
R7708 CS_BIAS.n279 CS_BIAS.n278 161.3
R7709 CS_BIAS.n277 CS_BIAS.n235 161.3
R7710 CS_BIAS.n276 CS_BIAS.n275 161.3
R7711 CS_BIAS.n274 CS_BIAS.n236 161.3
R7712 CS_BIAS.n273 CS_BIAS.n272 161.3
R7713 CS_BIAS.n271 CS_BIAS.n237 161.3
R7714 CS_BIAS.n270 CS_BIAS.n269 161.3
R7715 CS_BIAS.n268 CS_BIAS.n238 161.3
R7716 CS_BIAS.n266 CS_BIAS.n265 161.3
R7717 CS_BIAS.n264 CS_BIAS.n239 161.3
R7718 CS_BIAS.n263 CS_BIAS.n262 161.3
R7719 CS_BIAS.n261 CS_BIAS.n240 161.3
R7720 CS_BIAS.n260 CS_BIAS.n259 161.3
R7721 CS_BIAS.n258 CS_BIAS.n241 161.3
R7722 CS_BIAS.n257 CS_BIAS.n256 161.3
R7723 CS_BIAS.n255 CS_BIAS.n242 161.3
R7724 CS_BIAS.n254 CS_BIAS.n253 161.3
R7725 CS_BIAS.n252 CS_BIAS.n243 161.3
R7726 CS_BIAS.n251 CS_BIAS.n250 161.3
R7727 CS_BIAS.n249 CS_BIAS.n244 161.3
R7728 CS_BIAS.n248 CS_BIAS.n247 161.3
R7729 CS_BIAS.n85 CS_BIAS.n84 161.3
R7730 CS_BIAS.n86 CS_BIAS.n81 161.3
R7731 CS_BIAS.n88 CS_BIAS.n87 161.3
R7732 CS_BIAS.n89 CS_BIAS.n80 161.3
R7733 CS_BIAS.n91 CS_BIAS.n90 161.3
R7734 CS_BIAS.n92 CS_BIAS.n79 161.3
R7735 CS_BIAS.n94 CS_BIAS.n93 161.3
R7736 CS_BIAS.n95 CS_BIAS.n78 161.3
R7737 CS_BIAS.n97 CS_BIAS.n96 161.3
R7738 CS_BIAS.n98 CS_BIAS.n77 161.3
R7739 CS_BIAS.n100 CS_BIAS.n99 161.3
R7740 CS_BIAS.n101 CS_BIAS.n76 161.3
R7741 CS_BIAS.n103 CS_BIAS.n102 161.3
R7742 CS_BIAS.n105 CS_BIAS.n75 161.3
R7743 CS_BIAS.n107 CS_BIAS.n106 161.3
R7744 CS_BIAS.n108 CS_BIAS.n74 161.3
R7745 CS_BIAS.n110 CS_BIAS.n109 161.3
R7746 CS_BIAS.n111 CS_BIAS.n73 161.3
R7747 CS_BIAS.n113 CS_BIAS.n112 161.3
R7748 CS_BIAS.n114 CS_BIAS.n72 161.3
R7749 CS_BIAS.n116 CS_BIAS.n115 161.3
R7750 CS_BIAS.n117 CS_BIAS.n71 161.3
R7751 CS_BIAS.n119 CS_BIAS.n118 161.3
R7752 CS_BIAS.n120 CS_BIAS.n70 161.3
R7753 CS_BIAS.n122 CS_BIAS.n121 161.3
R7754 CS_BIAS.n124 CS_BIAS.n69 161.3
R7755 CS_BIAS.n126 CS_BIAS.n125 161.3
R7756 CS_BIAS.n127 CS_BIAS.n68 161.3
R7757 CS_BIAS.n129 CS_BIAS.n128 161.3
R7758 CS_BIAS.n130 CS_BIAS.n67 161.3
R7759 CS_BIAS.n132 CS_BIAS.n131 161.3
R7760 CS_BIAS.n133 CS_BIAS.n66 161.3
R7761 CS_BIAS.n135 CS_BIAS.n134 161.3
R7762 CS_BIAS.n136 CS_BIAS.n65 161.3
R7763 CS_BIAS.n138 CS_BIAS.n137 161.3
R7764 CS_BIAS.n139 CS_BIAS.n64 161.3
R7765 CS_BIAS.n141 CS_BIAS.n140 161.3
R7766 CS_BIAS.n142 CS_BIAS.n63 161.3
R7767 CS_BIAS.n145 CS_BIAS.n144 161.3
R7768 CS_BIAS.n146 CS_BIAS.n62 161.3
R7769 CS_BIAS.n148 CS_BIAS.n147 161.3
R7770 CS_BIAS.n149 CS_BIAS.n61 161.3
R7771 CS_BIAS.n151 CS_BIAS.n150 161.3
R7772 CS_BIAS.n152 CS_BIAS.n60 161.3
R7773 CS_BIAS.n154 CS_BIAS.n153 161.3
R7774 CS_BIAS.n155 CS_BIAS.n59 161.3
R7775 CS_BIAS.n157 CS_BIAS.n156 161.3
R7776 CS_BIAS.n158 CS_BIAS.n58 161.3
R7777 CS_BIAS.n160 CS_BIAS.n159 161.3
R7778 CS_BIAS.n161 CS_BIAS.n57 161.3
R7779 CS_BIAS.n28 CS_BIAS.n27 161.3
R7780 CS_BIAS.n29 CS_BIAS.n24 161.3
R7781 CS_BIAS.n31 CS_BIAS.n30 161.3
R7782 CS_BIAS.n32 CS_BIAS.n23 161.3
R7783 CS_BIAS.n34 CS_BIAS.n33 161.3
R7784 CS_BIAS.n35 CS_BIAS.n22 161.3
R7785 CS_BIAS.n37 CS_BIAS.n36 161.3
R7786 CS_BIAS.n38 CS_BIAS.n21 161.3
R7787 CS_BIAS.n40 CS_BIAS.n39 161.3
R7788 CS_BIAS.n41 CS_BIAS.n20 161.3
R7789 CS_BIAS.n43 CS_BIAS.n42 161.3
R7790 CS_BIAS.n44 CS_BIAS.n19 161.3
R7791 CS_BIAS.n46 CS_BIAS.n45 161.3
R7792 CS_BIAS.n48 CS_BIAS.n18 161.3
R7793 CS_BIAS.n50 CS_BIAS.n49 161.3
R7794 CS_BIAS.n51 CS_BIAS.n17 161.3
R7795 CS_BIAS.n53 CS_BIAS.n52 161.3
R7796 CS_BIAS.n54 CS_BIAS.n16 161.3
R7797 CS_BIAS.n56 CS_BIAS.n55 161.3
R7798 CS_BIAS.n170 CS_BIAS.n15 161.3
R7799 CS_BIAS.n172 CS_BIAS.n171 161.3
R7800 CS_BIAS.n173 CS_BIAS.n14 161.3
R7801 CS_BIAS.n175 CS_BIAS.n174 161.3
R7802 CS_BIAS.n176 CS_BIAS.n13 161.3
R7803 CS_BIAS.n178 CS_BIAS.n177 161.3
R7804 CS_BIAS.n180 CS_BIAS.n12 161.3
R7805 CS_BIAS.n182 CS_BIAS.n181 161.3
R7806 CS_BIAS.n183 CS_BIAS.n11 161.3
R7807 CS_BIAS.n185 CS_BIAS.n184 161.3
R7808 CS_BIAS.n186 CS_BIAS.n10 161.3
R7809 CS_BIAS.n188 CS_BIAS.n187 161.3
R7810 CS_BIAS.n189 CS_BIAS.n9 161.3
R7811 CS_BIAS.n191 CS_BIAS.n190 161.3
R7812 CS_BIAS.n192 CS_BIAS.n8 161.3
R7813 CS_BIAS.n194 CS_BIAS.n193 161.3
R7814 CS_BIAS.n195 CS_BIAS.n7 161.3
R7815 CS_BIAS.n197 CS_BIAS.n196 161.3
R7816 CS_BIAS.n198 CS_BIAS.n6 161.3
R7817 CS_BIAS.n201 CS_BIAS.n200 161.3
R7818 CS_BIAS.n202 CS_BIAS.n5 161.3
R7819 CS_BIAS.n204 CS_BIAS.n203 161.3
R7820 CS_BIAS.n205 CS_BIAS.n4 161.3
R7821 CS_BIAS.n207 CS_BIAS.n206 161.3
R7822 CS_BIAS.n208 CS_BIAS.n3 161.3
R7823 CS_BIAS.n210 CS_BIAS.n209 161.3
R7824 CS_BIAS.n211 CS_BIAS.n2 161.3
R7825 CS_BIAS.n213 CS_BIAS.n212 161.3
R7826 CS_BIAS.n214 CS_BIAS.n1 161.3
R7827 CS_BIAS.n216 CS_BIAS.n215 161.3
R7828 CS_BIAS.n217 CS_BIAS.n0 161.3
R7829 CS_BIAS.n652 CS_BIAS.n548 161.3
R7830 CS_BIAS.n651 CS_BIAS.n650 161.3
R7831 CS_BIAS.n649 CS_BIAS.n549 161.3
R7832 CS_BIAS.n648 CS_BIAS.n647 161.3
R7833 CS_BIAS.n646 CS_BIAS.n550 161.3
R7834 CS_BIAS.n645 CS_BIAS.n644 161.3
R7835 CS_BIAS.n643 CS_BIAS.n551 161.3
R7836 CS_BIAS.n642 CS_BIAS.n641 161.3
R7837 CS_BIAS.n640 CS_BIAS.n552 161.3
R7838 CS_BIAS.n639 CS_BIAS.n638 161.3
R7839 CS_BIAS.n637 CS_BIAS.n553 161.3
R7840 CS_BIAS.n636 CS_BIAS.n635 161.3
R7841 CS_BIAS.n633 CS_BIAS.n554 161.3
R7842 CS_BIAS.n632 CS_BIAS.n631 161.3
R7843 CS_BIAS.n630 CS_BIAS.n555 161.3
R7844 CS_BIAS.n629 CS_BIAS.n628 161.3
R7845 CS_BIAS.n627 CS_BIAS.n556 161.3
R7846 CS_BIAS.n626 CS_BIAS.n625 161.3
R7847 CS_BIAS.n624 CS_BIAS.n557 161.3
R7848 CS_BIAS.n623 CS_BIAS.n622 161.3
R7849 CS_BIAS.n621 CS_BIAS.n558 161.3
R7850 CS_BIAS.n620 CS_BIAS.n619 161.3
R7851 CS_BIAS.n618 CS_BIAS.n559 161.3
R7852 CS_BIAS.n617 CS_BIAS.n616 161.3
R7853 CS_BIAS.n615 CS_BIAS.n560 161.3
R7854 CS_BIAS.n613 CS_BIAS.n612 161.3
R7855 CS_BIAS.n611 CS_BIAS.n561 161.3
R7856 CS_BIAS.n610 CS_BIAS.n609 161.3
R7857 CS_BIAS.n608 CS_BIAS.n562 161.3
R7858 CS_BIAS.n607 CS_BIAS.n606 161.3
R7859 CS_BIAS.n605 CS_BIAS.n563 161.3
R7860 CS_BIAS.n604 CS_BIAS.n603 161.3
R7861 CS_BIAS.n602 CS_BIAS.n564 161.3
R7862 CS_BIAS.n601 CS_BIAS.n600 161.3
R7863 CS_BIAS.n599 CS_BIAS.n565 161.3
R7864 CS_BIAS.n598 CS_BIAS.n597 161.3
R7865 CS_BIAS.n596 CS_BIAS.n566 161.3
R7866 CS_BIAS.n594 CS_BIAS.n593 161.3
R7867 CS_BIAS.n592 CS_BIAS.n567 161.3
R7868 CS_BIAS.n591 CS_BIAS.n590 161.3
R7869 CS_BIAS.n589 CS_BIAS.n568 161.3
R7870 CS_BIAS.n588 CS_BIAS.n587 161.3
R7871 CS_BIAS.n586 CS_BIAS.n569 161.3
R7872 CS_BIAS.n585 CS_BIAS.n584 161.3
R7873 CS_BIAS.n583 CS_BIAS.n570 161.3
R7874 CS_BIAS.n582 CS_BIAS.n581 161.3
R7875 CS_BIAS.n580 CS_BIAS.n571 161.3
R7876 CS_BIAS.n579 CS_BIAS.n578 161.3
R7877 CS_BIAS.n577 CS_BIAS.n572 161.3
R7878 CS_BIAS.n576 CS_BIAS.n575 161.3
R7879 CS_BIAS.n491 CS_BIAS.n387 161.3
R7880 CS_BIAS.n490 CS_BIAS.n489 161.3
R7881 CS_BIAS.n488 CS_BIAS.n388 161.3
R7882 CS_BIAS.n487 CS_BIAS.n486 161.3
R7883 CS_BIAS.n485 CS_BIAS.n389 161.3
R7884 CS_BIAS.n484 CS_BIAS.n483 161.3
R7885 CS_BIAS.n482 CS_BIAS.n390 161.3
R7886 CS_BIAS.n481 CS_BIAS.n480 161.3
R7887 CS_BIAS.n479 CS_BIAS.n391 161.3
R7888 CS_BIAS.n478 CS_BIAS.n477 161.3
R7889 CS_BIAS.n476 CS_BIAS.n392 161.3
R7890 CS_BIAS.n475 CS_BIAS.n474 161.3
R7891 CS_BIAS.n472 CS_BIAS.n393 161.3
R7892 CS_BIAS.n471 CS_BIAS.n470 161.3
R7893 CS_BIAS.n469 CS_BIAS.n394 161.3
R7894 CS_BIAS.n468 CS_BIAS.n467 161.3
R7895 CS_BIAS.n466 CS_BIAS.n395 161.3
R7896 CS_BIAS.n465 CS_BIAS.n464 161.3
R7897 CS_BIAS.n463 CS_BIAS.n396 161.3
R7898 CS_BIAS.n462 CS_BIAS.n461 161.3
R7899 CS_BIAS.n460 CS_BIAS.n397 161.3
R7900 CS_BIAS.n459 CS_BIAS.n458 161.3
R7901 CS_BIAS.n457 CS_BIAS.n398 161.3
R7902 CS_BIAS.n456 CS_BIAS.n455 161.3
R7903 CS_BIAS.n454 CS_BIAS.n399 161.3
R7904 CS_BIAS.n452 CS_BIAS.n451 161.3
R7905 CS_BIAS.n450 CS_BIAS.n400 161.3
R7906 CS_BIAS.n449 CS_BIAS.n448 161.3
R7907 CS_BIAS.n447 CS_BIAS.n401 161.3
R7908 CS_BIAS.n446 CS_BIAS.n445 161.3
R7909 CS_BIAS.n444 CS_BIAS.n402 161.3
R7910 CS_BIAS.n443 CS_BIAS.n442 161.3
R7911 CS_BIAS.n441 CS_BIAS.n403 161.3
R7912 CS_BIAS.n440 CS_BIAS.n439 161.3
R7913 CS_BIAS.n438 CS_BIAS.n404 161.3
R7914 CS_BIAS.n437 CS_BIAS.n436 161.3
R7915 CS_BIAS.n435 CS_BIAS.n405 161.3
R7916 CS_BIAS.n433 CS_BIAS.n432 161.3
R7917 CS_BIAS.n431 CS_BIAS.n406 161.3
R7918 CS_BIAS.n430 CS_BIAS.n429 161.3
R7919 CS_BIAS.n428 CS_BIAS.n407 161.3
R7920 CS_BIAS.n427 CS_BIAS.n426 161.3
R7921 CS_BIAS.n425 CS_BIAS.n408 161.3
R7922 CS_BIAS.n424 CS_BIAS.n423 161.3
R7923 CS_BIAS.n422 CS_BIAS.n409 161.3
R7924 CS_BIAS.n421 CS_BIAS.n420 161.3
R7925 CS_BIAS.n419 CS_BIAS.n410 161.3
R7926 CS_BIAS.n418 CS_BIAS.n417 161.3
R7927 CS_BIAS.n416 CS_BIAS.n411 161.3
R7928 CS_BIAS.n415 CS_BIAS.n414 161.3
R7929 CS_BIAS.n384 CS_BIAS.n383 161.3
R7930 CS_BIAS.n382 CS_BIAS.n344 161.3
R7931 CS_BIAS.n381 CS_BIAS.n380 161.3
R7932 CS_BIAS.n379 CS_BIAS.n345 161.3
R7933 CS_BIAS.n378 CS_BIAS.n377 161.3
R7934 CS_BIAS.n376 CS_BIAS.n346 161.3
R7935 CS_BIAS.n374 CS_BIAS.n373 161.3
R7936 CS_BIAS.n372 CS_BIAS.n347 161.3
R7937 CS_BIAS.n371 CS_BIAS.n370 161.3
R7938 CS_BIAS.n369 CS_BIAS.n348 161.3
R7939 CS_BIAS.n368 CS_BIAS.n367 161.3
R7940 CS_BIAS.n366 CS_BIAS.n349 161.3
R7941 CS_BIAS.n365 CS_BIAS.n364 161.3
R7942 CS_BIAS.n363 CS_BIAS.n350 161.3
R7943 CS_BIAS.n362 CS_BIAS.n361 161.3
R7944 CS_BIAS.n360 CS_BIAS.n351 161.3
R7945 CS_BIAS.n359 CS_BIAS.n358 161.3
R7946 CS_BIAS.n357 CS_BIAS.n352 161.3
R7947 CS_BIAS.n356 CS_BIAS.n355 161.3
R7948 CS_BIAS.n545 CS_BIAS.n328 161.3
R7949 CS_BIAS.n544 CS_BIAS.n543 161.3
R7950 CS_BIAS.n542 CS_BIAS.n329 161.3
R7951 CS_BIAS.n541 CS_BIAS.n540 161.3
R7952 CS_BIAS.n539 CS_BIAS.n330 161.3
R7953 CS_BIAS.n538 CS_BIAS.n537 161.3
R7954 CS_BIAS.n536 CS_BIAS.n331 161.3
R7955 CS_BIAS.n535 CS_BIAS.n534 161.3
R7956 CS_BIAS.n533 CS_BIAS.n332 161.3
R7957 CS_BIAS.n532 CS_BIAS.n531 161.3
R7958 CS_BIAS.n530 CS_BIAS.n333 161.3
R7959 CS_BIAS.n529 CS_BIAS.n528 161.3
R7960 CS_BIAS.n526 CS_BIAS.n334 161.3
R7961 CS_BIAS.n525 CS_BIAS.n524 161.3
R7962 CS_BIAS.n523 CS_BIAS.n335 161.3
R7963 CS_BIAS.n522 CS_BIAS.n521 161.3
R7964 CS_BIAS.n520 CS_BIAS.n336 161.3
R7965 CS_BIAS.n519 CS_BIAS.n518 161.3
R7966 CS_BIAS.n517 CS_BIAS.n337 161.3
R7967 CS_BIAS.n516 CS_BIAS.n515 161.3
R7968 CS_BIAS.n514 CS_BIAS.n338 161.3
R7969 CS_BIAS.n513 CS_BIAS.n512 161.3
R7970 CS_BIAS.n511 CS_BIAS.n339 161.3
R7971 CS_BIAS.n510 CS_BIAS.n509 161.3
R7972 CS_BIAS.n508 CS_BIAS.n340 161.3
R7973 CS_BIAS.n506 CS_BIAS.n505 161.3
R7974 CS_BIAS.n504 CS_BIAS.n341 161.3
R7975 CS_BIAS.n503 CS_BIAS.n502 161.3
R7976 CS_BIAS.n501 CS_BIAS.n342 161.3
R7977 CS_BIAS.n500 CS_BIAS.n499 161.3
R7978 CS_BIAS.n498 CS_BIAS.n343 161.3
R7979 CS_BIAS.n168 CS_BIAS.n167 91.4836
R7980 CS_BIAS.n496 CS_BIAS.n385 91.4836
R7981 CS_BIAS.n168 CS_BIAS.n166 88.7853
R7982 CS_BIAS.n165 CS_BIAS.n164 88.7853
R7983 CS_BIAS.n495 CS_BIAS.n494 88.7853
R7984 CS_BIAS.n496 CS_BIAS.n386 88.7853
R7985 CS_BIAS.n83 CS_BIAS.n82 69.1729
R7986 CS_BIAS.n26 CS_BIAS.n25 69.1729
R7987 CS_BIAS.n246 CS_BIAS.n245 69.1729
R7988 CS_BIAS.n574 CS_BIAS.n573 69.1729
R7989 CS_BIAS.n413 CS_BIAS.n412 69.1729
R7990 CS_BIAS.n354 CS_BIAS.n353 69.1729
R7991 CS_BIAS.n326 CS_BIAS.n325 57.8583
R7992 CS_BIAS.n163 CS_BIAS.n162 57.8583
R7993 CS_BIAS.n219 CS_BIAS.n218 57.8583
R7994 CS_BIAS.n654 CS_BIAS.n653 57.8583
R7995 CS_BIAS.n493 CS_BIAS.n492 57.8583
R7996 CS_BIAS.n547 CS_BIAS.n546 57.8583
R7997 CS_BIAS.n275 CS_BIAS.n235 56.5617
R7998 CS_BIAS.n112 CS_BIAS.n72 56.5617
R7999 CS_BIAS.n55 CS_BIAS.n15 56.5617
R8000 CS_BIAS.n603 CS_BIAS.n563 56.5617
R8001 CS_BIAS.n442 CS_BIAS.n402 56.5617
R8002 CS_BIAS.n383 CS_BIAS.n343 56.5617
R8003 CS_BIAS.n317 CS_BIAS.n223 56.5617
R8004 CS_BIAS.n154 CS_BIAS.n60 56.5617
R8005 CS_BIAS.n210 CS_BIAS.n3 56.5617
R8006 CS_BIAS.n645 CS_BIAS.n551 56.5617
R8007 CS_BIAS.n484 CS_BIAS.n390 56.5617
R8008 CS_BIAS.n538 CS_BIAS.n331 56.5617
R8009 CS_BIAS.n246 CS_BIAS.t37 48.4449
R8010 CS_BIAS.n574 CS_BIAS.t25 48.4449
R8011 CS_BIAS.n413 CS_BIAS.t2 48.4449
R8012 CS_BIAS.n354 CS_BIAS.t34 48.4449
R8013 CS_BIAS.n83 CS_BIAS.t10 48.4445
R8014 CS_BIAS.n26 CS_BIAS.t36 48.4445
R8015 CS_BIAS.n256 CS_BIAS.n255 41.5458
R8016 CS_BIAS.n298 CS_BIAS.n229 41.5458
R8017 CS_BIAS.n135 CS_BIAS.n66 41.5458
R8018 CS_BIAS.n93 CS_BIAS.n92 41.5458
R8019 CS_BIAS.n191 CS_BIAS.n9 41.5458
R8020 CS_BIAS.n36 CS_BIAS.n35 41.5458
R8021 CS_BIAS.n584 CS_BIAS.n583 41.5458
R8022 CS_BIAS.n626 CS_BIAS.n557 41.5458
R8023 CS_BIAS.n423 CS_BIAS.n422 41.5458
R8024 CS_BIAS.n465 CS_BIAS.n396 41.5458
R8025 CS_BIAS.n519 CS_BIAS.n337 41.5458
R8026 CS_BIAS.n364 CS_BIAS.n363 41.5458
R8027 CS_BIAS.n256 CS_BIAS.n241 39.6083
R8028 CS_BIAS.n294 CS_BIAS.n229 39.6083
R8029 CS_BIAS.n131 CS_BIAS.n66 39.6083
R8030 CS_BIAS.n93 CS_BIAS.n78 39.6083
R8031 CS_BIAS.n187 CS_BIAS.n9 39.6083
R8032 CS_BIAS.n36 CS_BIAS.n21 39.6083
R8033 CS_BIAS.n584 CS_BIAS.n569 39.6083
R8034 CS_BIAS.n622 CS_BIAS.n557 39.6083
R8035 CS_BIAS.n423 CS_BIAS.n408 39.6083
R8036 CS_BIAS.n461 CS_BIAS.n396 39.6083
R8037 CS_BIAS.n515 CS_BIAS.n337 39.6083
R8038 CS_BIAS.n364 CS_BIAS.n349 39.6083
R8039 CS_BIAS.n255 CS_BIAS.n254 24.5923
R8040 CS_BIAS.n254 CS_BIAS.n243 24.5923
R8041 CS_BIAS.n250 CS_BIAS.n243 24.5923
R8042 CS_BIAS.n250 CS_BIAS.n249 24.5923
R8043 CS_BIAS.n249 CS_BIAS.n248 24.5923
R8044 CS_BIAS.n275 CS_BIAS.n274 24.5923
R8045 CS_BIAS.n274 CS_BIAS.n273 24.5923
R8046 CS_BIAS.n273 CS_BIAS.n237 24.5923
R8047 CS_BIAS.n269 CS_BIAS.n237 24.5923
R8048 CS_BIAS.n269 CS_BIAS.n268 24.5923
R8049 CS_BIAS.n266 CS_BIAS.n239 24.5923
R8050 CS_BIAS.n262 CS_BIAS.n239 24.5923
R8051 CS_BIAS.n262 CS_BIAS.n261 24.5923
R8052 CS_BIAS.n261 CS_BIAS.n260 24.5923
R8053 CS_BIAS.n260 CS_BIAS.n241 24.5923
R8054 CS_BIAS.n294 CS_BIAS.n293 24.5923
R8055 CS_BIAS.n293 CS_BIAS.n292 24.5923
R8056 CS_BIAS.n292 CS_BIAS.n231 24.5923
R8057 CS_BIAS.n288 CS_BIAS.n231 24.5923
R8058 CS_BIAS.n288 CS_BIAS.n287 24.5923
R8059 CS_BIAS.n285 CS_BIAS.n233 24.5923
R8060 CS_BIAS.n281 CS_BIAS.n233 24.5923
R8061 CS_BIAS.n281 CS_BIAS.n280 24.5923
R8062 CS_BIAS.n280 CS_BIAS.n279 24.5923
R8063 CS_BIAS.n279 CS_BIAS.n235 24.5923
R8064 CS_BIAS.n313 CS_BIAS.n223 24.5923
R8065 CS_BIAS.n313 CS_BIAS.n312 24.5923
R8066 CS_BIAS.n312 CS_BIAS.n311 24.5923
R8067 CS_BIAS.n311 CS_BIAS.n225 24.5923
R8068 CS_BIAS.n307 CS_BIAS.n225 24.5923
R8069 CS_BIAS.n305 CS_BIAS.n304 24.5923
R8070 CS_BIAS.n304 CS_BIAS.n227 24.5923
R8071 CS_BIAS.n300 CS_BIAS.n227 24.5923
R8072 CS_BIAS.n300 CS_BIAS.n299 24.5923
R8073 CS_BIAS.n299 CS_BIAS.n298 24.5923
R8074 CS_BIAS.n324 CS_BIAS.n323 24.5923
R8075 CS_BIAS.n323 CS_BIAS.n221 24.5923
R8076 CS_BIAS.n319 CS_BIAS.n221 24.5923
R8077 CS_BIAS.n319 CS_BIAS.n318 24.5923
R8078 CS_BIAS.n318 CS_BIAS.n317 24.5923
R8079 CS_BIAS.n161 CS_BIAS.n160 24.5923
R8080 CS_BIAS.n160 CS_BIAS.n58 24.5923
R8081 CS_BIAS.n156 CS_BIAS.n58 24.5923
R8082 CS_BIAS.n156 CS_BIAS.n155 24.5923
R8083 CS_BIAS.n155 CS_BIAS.n154 24.5923
R8084 CS_BIAS.n150 CS_BIAS.n60 24.5923
R8085 CS_BIAS.n150 CS_BIAS.n149 24.5923
R8086 CS_BIAS.n149 CS_BIAS.n148 24.5923
R8087 CS_BIAS.n148 CS_BIAS.n62 24.5923
R8088 CS_BIAS.n144 CS_BIAS.n62 24.5923
R8089 CS_BIAS.n142 CS_BIAS.n141 24.5923
R8090 CS_BIAS.n141 CS_BIAS.n64 24.5923
R8091 CS_BIAS.n137 CS_BIAS.n64 24.5923
R8092 CS_BIAS.n137 CS_BIAS.n136 24.5923
R8093 CS_BIAS.n136 CS_BIAS.n135 24.5923
R8094 CS_BIAS.n131 CS_BIAS.n130 24.5923
R8095 CS_BIAS.n130 CS_BIAS.n129 24.5923
R8096 CS_BIAS.n129 CS_BIAS.n68 24.5923
R8097 CS_BIAS.n125 CS_BIAS.n68 24.5923
R8098 CS_BIAS.n125 CS_BIAS.n124 24.5923
R8099 CS_BIAS.n122 CS_BIAS.n70 24.5923
R8100 CS_BIAS.n118 CS_BIAS.n70 24.5923
R8101 CS_BIAS.n118 CS_BIAS.n117 24.5923
R8102 CS_BIAS.n117 CS_BIAS.n116 24.5923
R8103 CS_BIAS.n116 CS_BIAS.n72 24.5923
R8104 CS_BIAS.n112 CS_BIAS.n111 24.5923
R8105 CS_BIAS.n111 CS_BIAS.n110 24.5923
R8106 CS_BIAS.n110 CS_BIAS.n74 24.5923
R8107 CS_BIAS.n106 CS_BIAS.n74 24.5923
R8108 CS_BIAS.n106 CS_BIAS.n105 24.5923
R8109 CS_BIAS.n103 CS_BIAS.n76 24.5923
R8110 CS_BIAS.n99 CS_BIAS.n76 24.5923
R8111 CS_BIAS.n99 CS_BIAS.n98 24.5923
R8112 CS_BIAS.n98 CS_BIAS.n97 24.5923
R8113 CS_BIAS.n97 CS_BIAS.n78 24.5923
R8114 CS_BIAS.n92 CS_BIAS.n91 24.5923
R8115 CS_BIAS.n91 CS_BIAS.n80 24.5923
R8116 CS_BIAS.n87 CS_BIAS.n80 24.5923
R8117 CS_BIAS.n87 CS_BIAS.n86 24.5923
R8118 CS_BIAS.n86 CS_BIAS.n85 24.5923
R8119 CS_BIAS.n217 CS_BIAS.n216 24.5923
R8120 CS_BIAS.n216 CS_BIAS.n1 24.5923
R8121 CS_BIAS.n212 CS_BIAS.n1 24.5923
R8122 CS_BIAS.n212 CS_BIAS.n211 24.5923
R8123 CS_BIAS.n211 CS_BIAS.n210 24.5923
R8124 CS_BIAS.n206 CS_BIAS.n3 24.5923
R8125 CS_BIAS.n206 CS_BIAS.n205 24.5923
R8126 CS_BIAS.n205 CS_BIAS.n204 24.5923
R8127 CS_BIAS.n204 CS_BIAS.n5 24.5923
R8128 CS_BIAS.n200 CS_BIAS.n5 24.5923
R8129 CS_BIAS.n198 CS_BIAS.n197 24.5923
R8130 CS_BIAS.n197 CS_BIAS.n7 24.5923
R8131 CS_BIAS.n193 CS_BIAS.n7 24.5923
R8132 CS_BIAS.n193 CS_BIAS.n192 24.5923
R8133 CS_BIAS.n192 CS_BIAS.n191 24.5923
R8134 CS_BIAS.n187 CS_BIAS.n186 24.5923
R8135 CS_BIAS.n186 CS_BIAS.n185 24.5923
R8136 CS_BIAS.n185 CS_BIAS.n11 24.5923
R8137 CS_BIAS.n181 CS_BIAS.n11 24.5923
R8138 CS_BIAS.n181 CS_BIAS.n180 24.5923
R8139 CS_BIAS.n178 CS_BIAS.n13 24.5923
R8140 CS_BIAS.n174 CS_BIAS.n13 24.5923
R8141 CS_BIAS.n174 CS_BIAS.n173 24.5923
R8142 CS_BIAS.n173 CS_BIAS.n172 24.5923
R8143 CS_BIAS.n172 CS_BIAS.n15 24.5923
R8144 CS_BIAS.n55 CS_BIAS.n54 24.5923
R8145 CS_BIAS.n54 CS_BIAS.n53 24.5923
R8146 CS_BIAS.n53 CS_BIAS.n17 24.5923
R8147 CS_BIAS.n49 CS_BIAS.n17 24.5923
R8148 CS_BIAS.n49 CS_BIAS.n48 24.5923
R8149 CS_BIAS.n46 CS_BIAS.n19 24.5923
R8150 CS_BIAS.n42 CS_BIAS.n19 24.5923
R8151 CS_BIAS.n42 CS_BIAS.n41 24.5923
R8152 CS_BIAS.n41 CS_BIAS.n40 24.5923
R8153 CS_BIAS.n40 CS_BIAS.n21 24.5923
R8154 CS_BIAS.n35 CS_BIAS.n34 24.5923
R8155 CS_BIAS.n34 CS_BIAS.n23 24.5923
R8156 CS_BIAS.n30 CS_BIAS.n23 24.5923
R8157 CS_BIAS.n30 CS_BIAS.n29 24.5923
R8158 CS_BIAS.n29 CS_BIAS.n28 24.5923
R8159 CS_BIAS.n577 CS_BIAS.n576 24.5923
R8160 CS_BIAS.n578 CS_BIAS.n577 24.5923
R8161 CS_BIAS.n578 CS_BIAS.n571 24.5923
R8162 CS_BIAS.n582 CS_BIAS.n571 24.5923
R8163 CS_BIAS.n583 CS_BIAS.n582 24.5923
R8164 CS_BIAS.n588 CS_BIAS.n569 24.5923
R8165 CS_BIAS.n589 CS_BIAS.n588 24.5923
R8166 CS_BIAS.n590 CS_BIAS.n589 24.5923
R8167 CS_BIAS.n590 CS_BIAS.n567 24.5923
R8168 CS_BIAS.n594 CS_BIAS.n567 24.5923
R8169 CS_BIAS.n597 CS_BIAS.n596 24.5923
R8170 CS_BIAS.n597 CS_BIAS.n565 24.5923
R8171 CS_BIAS.n601 CS_BIAS.n565 24.5923
R8172 CS_BIAS.n602 CS_BIAS.n601 24.5923
R8173 CS_BIAS.n603 CS_BIAS.n602 24.5923
R8174 CS_BIAS.n607 CS_BIAS.n563 24.5923
R8175 CS_BIAS.n608 CS_BIAS.n607 24.5923
R8176 CS_BIAS.n609 CS_BIAS.n608 24.5923
R8177 CS_BIAS.n609 CS_BIAS.n561 24.5923
R8178 CS_BIAS.n613 CS_BIAS.n561 24.5923
R8179 CS_BIAS.n616 CS_BIAS.n615 24.5923
R8180 CS_BIAS.n616 CS_BIAS.n559 24.5923
R8181 CS_BIAS.n620 CS_BIAS.n559 24.5923
R8182 CS_BIAS.n621 CS_BIAS.n620 24.5923
R8183 CS_BIAS.n622 CS_BIAS.n621 24.5923
R8184 CS_BIAS.n627 CS_BIAS.n626 24.5923
R8185 CS_BIAS.n628 CS_BIAS.n627 24.5923
R8186 CS_BIAS.n628 CS_BIAS.n555 24.5923
R8187 CS_BIAS.n632 CS_BIAS.n555 24.5923
R8188 CS_BIAS.n633 CS_BIAS.n632 24.5923
R8189 CS_BIAS.n635 CS_BIAS.n553 24.5923
R8190 CS_BIAS.n639 CS_BIAS.n553 24.5923
R8191 CS_BIAS.n640 CS_BIAS.n639 24.5923
R8192 CS_BIAS.n641 CS_BIAS.n640 24.5923
R8193 CS_BIAS.n641 CS_BIAS.n551 24.5923
R8194 CS_BIAS.n646 CS_BIAS.n645 24.5923
R8195 CS_BIAS.n647 CS_BIAS.n646 24.5923
R8196 CS_BIAS.n647 CS_BIAS.n549 24.5923
R8197 CS_BIAS.n651 CS_BIAS.n549 24.5923
R8198 CS_BIAS.n652 CS_BIAS.n651 24.5923
R8199 CS_BIAS.n416 CS_BIAS.n415 24.5923
R8200 CS_BIAS.n417 CS_BIAS.n416 24.5923
R8201 CS_BIAS.n417 CS_BIAS.n410 24.5923
R8202 CS_BIAS.n421 CS_BIAS.n410 24.5923
R8203 CS_BIAS.n422 CS_BIAS.n421 24.5923
R8204 CS_BIAS.n427 CS_BIAS.n408 24.5923
R8205 CS_BIAS.n428 CS_BIAS.n427 24.5923
R8206 CS_BIAS.n429 CS_BIAS.n428 24.5923
R8207 CS_BIAS.n429 CS_BIAS.n406 24.5923
R8208 CS_BIAS.n433 CS_BIAS.n406 24.5923
R8209 CS_BIAS.n436 CS_BIAS.n435 24.5923
R8210 CS_BIAS.n436 CS_BIAS.n404 24.5923
R8211 CS_BIAS.n440 CS_BIAS.n404 24.5923
R8212 CS_BIAS.n441 CS_BIAS.n440 24.5923
R8213 CS_BIAS.n442 CS_BIAS.n441 24.5923
R8214 CS_BIAS.n446 CS_BIAS.n402 24.5923
R8215 CS_BIAS.n447 CS_BIAS.n446 24.5923
R8216 CS_BIAS.n448 CS_BIAS.n447 24.5923
R8217 CS_BIAS.n448 CS_BIAS.n400 24.5923
R8218 CS_BIAS.n452 CS_BIAS.n400 24.5923
R8219 CS_BIAS.n455 CS_BIAS.n454 24.5923
R8220 CS_BIAS.n455 CS_BIAS.n398 24.5923
R8221 CS_BIAS.n459 CS_BIAS.n398 24.5923
R8222 CS_BIAS.n460 CS_BIAS.n459 24.5923
R8223 CS_BIAS.n461 CS_BIAS.n460 24.5923
R8224 CS_BIAS.n466 CS_BIAS.n465 24.5923
R8225 CS_BIAS.n467 CS_BIAS.n466 24.5923
R8226 CS_BIAS.n467 CS_BIAS.n394 24.5923
R8227 CS_BIAS.n471 CS_BIAS.n394 24.5923
R8228 CS_BIAS.n472 CS_BIAS.n471 24.5923
R8229 CS_BIAS.n474 CS_BIAS.n392 24.5923
R8230 CS_BIAS.n478 CS_BIAS.n392 24.5923
R8231 CS_BIAS.n479 CS_BIAS.n478 24.5923
R8232 CS_BIAS.n480 CS_BIAS.n479 24.5923
R8233 CS_BIAS.n480 CS_BIAS.n390 24.5923
R8234 CS_BIAS.n485 CS_BIAS.n484 24.5923
R8235 CS_BIAS.n486 CS_BIAS.n485 24.5923
R8236 CS_BIAS.n486 CS_BIAS.n388 24.5923
R8237 CS_BIAS.n490 CS_BIAS.n388 24.5923
R8238 CS_BIAS.n491 CS_BIAS.n490 24.5923
R8239 CS_BIAS.n539 CS_BIAS.n538 24.5923
R8240 CS_BIAS.n540 CS_BIAS.n539 24.5923
R8241 CS_BIAS.n540 CS_BIAS.n329 24.5923
R8242 CS_BIAS.n544 CS_BIAS.n329 24.5923
R8243 CS_BIAS.n545 CS_BIAS.n544 24.5923
R8244 CS_BIAS.n520 CS_BIAS.n519 24.5923
R8245 CS_BIAS.n521 CS_BIAS.n520 24.5923
R8246 CS_BIAS.n521 CS_BIAS.n335 24.5923
R8247 CS_BIAS.n525 CS_BIAS.n335 24.5923
R8248 CS_BIAS.n526 CS_BIAS.n525 24.5923
R8249 CS_BIAS.n528 CS_BIAS.n333 24.5923
R8250 CS_BIAS.n532 CS_BIAS.n333 24.5923
R8251 CS_BIAS.n533 CS_BIAS.n532 24.5923
R8252 CS_BIAS.n534 CS_BIAS.n533 24.5923
R8253 CS_BIAS.n534 CS_BIAS.n331 24.5923
R8254 CS_BIAS.n500 CS_BIAS.n343 24.5923
R8255 CS_BIAS.n501 CS_BIAS.n500 24.5923
R8256 CS_BIAS.n502 CS_BIAS.n501 24.5923
R8257 CS_BIAS.n502 CS_BIAS.n341 24.5923
R8258 CS_BIAS.n506 CS_BIAS.n341 24.5923
R8259 CS_BIAS.n509 CS_BIAS.n508 24.5923
R8260 CS_BIAS.n509 CS_BIAS.n339 24.5923
R8261 CS_BIAS.n513 CS_BIAS.n339 24.5923
R8262 CS_BIAS.n514 CS_BIAS.n513 24.5923
R8263 CS_BIAS.n515 CS_BIAS.n514 24.5923
R8264 CS_BIAS.n357 CS_BIAS.n356 24.5923
R8265 CS_BIAS.n358 CS_BIAS.n357 24.5923
R8266 CS_BIAS.n358 CS_BIAS.n351 24.5923
R8267 CS_BIAS.n362 CS_BIAS.n351 24.5923
R8268 CS_BIAS.n363 CS_BIAS.n362 24.5923
R8269 CS_BIAS.n368 CS_BIAS.n349 24.5923
R8270 CS_BIAS.n369 CS_BIAS.n368 24.5923
R8271 CS_BIAS.n370 CS_BIAS.n369 24.5923
R8272 CS_BIAS.n370 CS_BIAS.n347 24.5923
R8273 CS_BIAS.n374 CS_BIAS.n347 24.5923
R8274 CS_BIAS.n377 CS_BIAS.n376 24.5923
R8275 CS_BIAS.n377 CS_BIAS.n345 24.5923
R8276 CS_BIAS.n381 CS_BIAS.n345 24.5923
R8277 CS_BIAS.n382 CS_BIAS.n381 24.5923
R8278 CS_BIAS.n383 CS_BIAS.n382 24.5923
R8279 CS_BIAS.n325 CS_BIAS.n324 19.674
R8280 CS_BIAS.n162 CS_BIAS.n161 19.674
R8281 CS_BIAS.n218 CS_BIAS.n217 19.674
R8282 CS_BIAS.n653 CS_BIAS.n652 19.674
R8283 CS_BIAS.n492 CS_BIAS.n491 19.674
R8284 CS_BIAS.n546 CS_BIAS.n545 19.674
R8285 CS_BIAS.n268 CS_BIAS.n267 18.6903
R8286 CS_BIAS.n286 CS_BIAS.n285 18.6903
R8287 CS_BIAS.n123 CS_BIAS.n122 18.6903
R8288 CS_BIAS.n105 CS_BIAS.n104 18.6903
R8289 CS_BIAS.n179 CS_BIAS.n178 18.6903
R8290 CS_BIAS.n48 CS_BIAS.n47 18.6903
R8291 CS_BIAS.n596 CS_BIAS.n595 18.6903
R8292 CS_BIAS.n614 CS_BIAS.n613 18.6903
R8293 CS_BIAS.n435 CS_BIAS.n434 18.6903
R8294 CS_BIAS.n453 CS_BIAS.n452 18.6903
R8295 CS_BIAS.n507 CS_BIAS.n506 18.6903
R8296 CS_BIAS.n376 CS_BIAS.n375 18.6903
R8297 CS_BIAS.n307 CS_BIAS.n306 17.7066
R8298 CS_BIAS.n144 CS_BIAS.n143 17.7066
R8299 CS_BIAS.n200 CS_BIAS.n199 17.7066
R8300 CS_BIAS.n635 CS_BIAS.n634 17.7066
R8301 CS_BIAS.n474 CS_BIAS.n473 17.7066
R8302 CS_BIAS.n528 CS_BIAS.n527 17.7066
R8303 CS_BIAS.n245 CS_BIAS.t31 15.2814
R8304 CS_BIAS.n267 CS_BIAS.t46 15.2814
R8305 CS_BIAS.n286 CS_BIAS.t39 15.2814
R8306 CS_BIAS.n306 CS_BIAS.t35 15.2814
R8307 CS_BIAS.n325 CS_BIAS.t27 15.2814
R8308 CS_BIAS.n162 CS_BIAS.t14 15.2814
R8309 CS_BIAS.n143 CS_BIAS.t20 15.2814
R8310 CS_BIAS.n123 CS_BIAS.t22 15.2814
R8311 CS_BIAS.n104 CS_BIAS.t12 15.2814
R8312 CS_BIAS.n82 CS_BIAS.t16 15.2814
R8313 CS_BIAS.n218 CS_BIAS.t33 15.2814
R8314 CS_BIAS.n199 CS_BIAS.t42 15.2814
R8315 CS_BIAS.n179 CS_BIAS.t29 15.2814
R8316 CS_BIAS.n47 CS_BIAS.t41 15.2814
R8317 CS_BIAS.n25 CS_BIAS.t26 15.2814
R8318 CS_BIAS.n573 CS_BIAS.t44 15.2814
R8319 CS_BIAS.n595 CS_BIAS.t30 15.2814
R8320 CS_BIAS.n614 CS_BIAS.t32 15.2814
R8321 CS_BIAS.n634 CS_BIAS.t45 15.2814
R8322 CS_BIAS.n653 CS_BIAS.t40 15.2814
R8323 CS_BIAS.n412 CS_BIAS.t18 15.2814
R8324 CS_BIAS.n434 CS_BIAS.t4 15.2814
R8325 CS_BIAS.n453 CS_BIAS.t6 15.2814
R8326 CS_BIAS.n473 CS_BIAS.t0 15.2814
R8327 CS_BIAS.n492 CS_BIAS.t8 15.2814
R8328 CS_BIAS.n546 CS_BIAS.t28 15.2814
R8329 CS_BIAS.n527 CS_BIAS.t38 15.2814
R8330 CS_BIAS.n507 CS_BIAS.t24 15.2814
R8331 CS_BIAS.n353 CS_BIAS.t47 15.2814
R8332 CS_BIAS.n375 CS_BIAS.t43 15.2814
R8333 CS_BIAS.n495 CS_BIAS.n493 13.602
R8334 CS_BIAS.n165 CS_BIAS.n163 13.6019
R8335 CS_BIAS.n656 CS_BIAS.n327 12.1432
R8336 CS_BIAS.n169 CS_BIAS.n168 9.50425
R8337 CS_BIAS.n497 CS_BIAS.n496 9.50425
R8338 CS_BIAS.n656 CS_BIAS.n655 8.92186
R8339 CS_BIAS.n655 CS_BIAS.n547 8.02792
R8340 CS_BIAS.n327 CS_BIAS.n219 8.02792
R8341 CS_BIAS.n248 CS_BIAS.n245 6.88621
R8342 CS_BIAS.n306 CS_BIAS.n305 6.88621
R8343 CS_BIAS.n143 CS_BIAS.n142 6.88621
R8344 CS_BIAS.n85 CS_BIAS.n82 6.88621
R8345 CS_BIAS.n199 CS_BIAS.n198 6.88621
R8346 CS_BIAS.n28 CS_BIAS.n25 6.88621
R8347 CS_BIAS.n576 CS_BIAS.n573 6.88621
R8348 CS_BIAS.n634 CS_BIAS.n633 6.88621
R8349 CS_BIAS.n415 CS_BIAS.n412 6.88621
R8350 CS_BIAS.n473 CS_BIAS.n472 6.88621
R8351 CS_BIAS.n527 CS_BIAS.n526 6.88621
R8352 CS_BIAS.n356 CS_BIAS.n353 6.88621
R8353 CS_BIAS.n267 CS_BIAS.n266 5.90254
R8354 CS_BIAS.n287 CS_BIAS.n286 5.90254
R8355 CS_BIAS.n124 CS_BIAS.n123 5.90254
R8356 CS_BIAS.n104 CS_BIAS.n103 5.90254
R8357 CS_BIAS.n180 CS_BIAS.n179 5.90254
R8358 CS_BIAS.n47 CS_BIAS.n46 5.90254
R8359 CS_BIAS.n595 CS_BIAS.n594 5.90254
R8360 CS_BIAS.n615 CS_BIAS.n614 5.90254
R8361 CS_BIAS.n434 CS_BIAS.n433 5.90254
R8362 CS_BIAS.n454 CS_BIAS.n453 5.90254
R8363 CS_BIAS.n508 CS_BIAS.n507 5.90254
R8364 CS_BIAS.n375 CS_BIAS.n374 5.90254
R8365 CS_BIAS.n327 CS_BIAS.n326 5.5658
R8366 CS_BIAS.n655 CS_BIAS.n654 5.5658
R8367 CS_BIAS.n167 CS_BIAS.t17 5.26646
R8368 CS_BIAS.n167 CS_BIAS.t11 5.26646
R8369 CS_BIAS.n166 CS_BIAS.t23 5.26646
R8370 CS_BIAS.n166 CS_BIAS.t13 5.26646
R8371 CS_BIAS.n164 CS_BIAS.t15 5.26646
R8372 CS_BIAS.n164 CS_BIAS.t21 5.26646
R8373 CS_BIAS.n494 CS_BIAS.t1 5.26646
R8374 CS_BIAS.n494 CS_BIAS.t9 5.26646
R8375 CS_BIAS.n386 CS_BIAS.t5 5.26646
R8376 CS_BIAS.n386 CS_BIAS.t7 5.26646
R8377 CS_BIAS.n385 CS_BIAS.t3 5.26646
R8378 CS_BIAS.n385 CS_BIAS.t19 5.26646
R8379 CS_BIAS CS_BIAS.n656 4.62792
R8380 CS_BIAS.n168 CS_BIAS.n165 2.69878
R8381 CS_BIAS.n496 CS_BIAS.n495 2.69878
R8382 CS_BIAS.n247 CS_BIAS.n246 1.00073
R8383 CS_BIAS.n575 CS_BIAS.n574 1.00073
R8384 CS_BIAS.n414 CS_BIAS.n413 1.00073
R8385 CS_BIAS.n355 CS_BIAS.n354 1.00073
R8386 CS_BIAS.n84 CS_BIAS.n83 1.00072
R8387 CS_BIAS.n27 CS_BIAS.n26 1.00072
R8388 CS_BIAS.n326 CS_BIAS.n220 0.502096
R8389 CS_BIAS.n163 CS_BIAS.n57 0.502096
R8390 CS_BIAS.n219 CS_BIAS.n0 0.502096
R8391 CS_BIAS.n654 CS_BIAS.n548 0.502096
R8392 CS_BIAS.n493 CS_BIAS.n387 0.502096
R8393 CS_BIAS.n547 CS_BIAS.n328 0.502096
R8394 CS_BIAS.n322 CS_BIAS.n220 0.189894
R8395 CS_BIAS.n322 CS_BIAS.n321 0.189894
R8396 CS_BIAS.n321 CS_BIAS.n320 0.189894
R8397 CS_BIAS.n320 CS_BIAS.n222 0.189894
R8398 CS_BIAS.n316 CS_BIAS.n222 0.189894
R8399 CS_BIAS.n316 CS_BIAS.n315 0.189894
R8400 CS_BIAS.n315 CS_BIAS.n314 0.189894
R8401 CS_BIAS.n314 CS_BIAS.n224 0.189894
R8402 CS_BIAS.n310 CS_BIAS.n224 0.189894
R8403 CS_BIAS.n310 CS_BIAS.n309 0.189894
R8404 CS_BIAS.n309 CS_BIAS.n308 0.189894
R8405 CS_BIAS.n308 CS_BIAS.n226 0.189894
R8406 CS_BIAS.n303 CS_BIAS.n226 0.189894
R8407 CS_BIAS.n303 CS_BIAS.n302 0.189894
R8408 CS_BIAS.n302 CS_BIAS.n301 0.189894
R8409 CS_BIAS.n301 CS_BIAS.n228 0.189894
R8410 CS_BIAS.n297 CS_BIAS.n228 0.189894
R8411 CS_BIAS.n297 CS_BIAS.n296 0.189894
R8412 CS_BIAS.n296 CS_BIAS.n295 0.189894
R8413 CS_BIAS.n295 CS_BIAS.n230 0.189894
R8414 CS_BIAS.n291 CS_BIAS.n230 0.189894
R8415 CS_BIAS.n291 CS_BIAS.n290 0.189894
R8416 CS_BIAS.n290 CS_BIAS.n289 0.189894
R8417 CS_BIAS.n289 CS_BIAS.n232 0.189894
R8418 CS_BIAS.n284 CS_BIAS.n232 0.189894
R8419 CS_BIAS.n284 CS_BIAS.n283 0.189894
R8420 CS_BIAS.n283 CS_BIAS.n282 0.189894
R8421 CS_BIAS.n282 CS_BIAS.n234 0.189894
R8422 CS_BIAS.n278 CS_BIAS.n234 0.189894
R8423 CS_BIAS.n278 CS_BIAS.n277 0.189894
R8424 CS_BIAS.n277 CS_BIAS.n276 0.189894
R8425 CS_BIAS.n276 CS_BIAS.n236 0.189894
R8426 CS_BIAS.n272 CS_BIAS.n236 0.189894
R8427 CS_BIAS.n272 CS_BIAS.n271 0.189894
R8428 CS_BIAS.n271 CS_BIAS.n270 0.189894
R8429 CS_BIAS.n270 CS_BIAS.n238 0.189894
R8430 CS_BIAS.n265 CS_BIAS.n238 0.189894
R8431 CS_BIAS.n265 CS_BIAS.n264 0.189894
R8432 CS_BIAS.n264 CS_BIAS.n263 0.189894
R8433 CS_BIAS.n263 CS_BIAS.n240 0.189894
R8434 CS_BIAS.n259 CS_BIAS.n240 0.189894
R8435 CS_BIAS.n259 CS_BIAS.n258 0.189894
R8436 CS_BIAS.n258 CS_BIAS.n257 0.189894
R8437 CS_BIAS.n257 CS_BIAS.n242 0.189894
R8438 CS_BIAS.n253 CS_BIAS.n242 0.189894
R8439 CS_BIAS.n253 CS_BIAS.n252 0.189894
R8440 CS_BIAS.n252 CS_BIAS.n251 0.189894
R8441 CS_BIAS.n251 CS_BIAS.n244 0.189894
R8442 CS_BIAS.n247 CS_BIAS.n244 0.189894
R8443 CS_BIAS.n159 CS_BIAS.n57 0.189894
R8444 CS_BIAS.n159 CS_BIAS.n158 0.189894
R8445 CS_BIAS.n158 CS_BIAS.n157 0.189894
R8446 CS_BIAS.n157 CS_BIAS.n59 0.189894
R8447 CS_BIAS.n153 CS_BIAS.n59 0.189894
R8448 CS_BIAS.n153 CS_BIAS.n152 0.189894
R8449 CS_BIAS.n152 CS_BIAS.n151 0.189894
R8450 CS_BIAS.n151 CS_BIAS.n61 0.189894
R8451 CS_BIAS.n147 CS_BIAS.n61 0.189894
R8452 CS_BIAS.n147 CS_BIAS.n146 0.189894
R8453 CS_BIAS.n146 CS_BIAS.n145 0.189894
R8454 CS_BIAS.n145 CS_BIAS.n63 0.189894
R8455 CS_BIAS.n140 CS_BIAS.n63 0.189894
R8456 CS_BIAS.n140 CS_BIAS.n139 0.189894
R8457 CS_BIAS.n139 CS_BIAS.n138 0.189894
R8458 CS_BIAS.n138 CS_BIAS.n65 0.189894
R8459 CS_BIAS.n134 CS_BIAS.n65 0.189894
R8460 CS_BIAS.n134 CS_BIAS.n133 0.189894
R8461 CS_BIAS.n133 CS_BIAS.n132 0.189894
R8462 CS_BIAS.n132 CS_BIAS.n67 0.189894
R8463 CS_BIAS.n128 CS_BIAS.n67 0.189894
R8464 CS_BIAS.n128 CS_BIAS.n127 0.189894
R8465 CS_BIAS.n127 CS_BIAS.n126 0.189894
R8466 CS_BIAS.n126 CS_BIAS.n69 0.189894
R8467 CS_BIAS.n121 CS_BIAS.n69 0.189894
R8468 CS_BIAS.n121 CS_BIAS.n120 0.189894
R8469 CS_BIAS.n120 CS_BIAS.n119 0.189894
R8470 CS_BIAS.n119 CS_BIAS.n71 0.189894
R8471 CS_BIAS.n115 CS_BIAS.n71 0.189894
R8472 CS_BIAS.n115 CS_BIAS.n114 0.189894
R8473 CS_BIAS.n114 CS_BIAS.n113 0.189894
R8474 CS_BIAS.n113 CS_BIAS.n73 0.189894
R8475 CS_BIAS.n109 CS_BIAS.n73 0.189894
R8476 CS_BIAS.n109 CS_BIAS.n108 0.189894
R8477 CS_BIAS.n108 CS_BIAS.n107 0.189894
R8478 CS_BIAS.n107 CS_BIAS.n75 0.189894
R8479 CS_BIAS.n102 CS_BIAS.n75 0.189894
R8480 CS_BIAS.n102 CS_BIAS.n101 0.189894
R8481 CS_BIAS.n101 CS_BIAS.n100 0.189894
R8482 CS_BIAS.n100 CS_BIAS.n77 0.189894
R8483 CS_BIAS.n96 CS_BIAS.n77 0.189894
R8484 CS_BIAS.n96 CS_BIAS.n95 0.189894
R8485 CS_BIAS.n95 CS_BIAS.n94 0.189894
R8486 CS_BIAS.n94 CS_BIAS.n79 0.189894
R8487 CS_BIAS.n90 CS_BIAS.n79 0.189894
R8488 CS_BIAS.n90 CS_BIAS.n89 0.189894
R8489 CS_BIAS.n89 CS_BIAS.n88 0.189894
R8490 CS_BIAS.n88 CS_BIAS.n81 0.189894
R8491 CS_BIAS.n84 CS_BIAS.n81 0.189894
R8492 CS_BIAS.n56 CS_BIAS.n16 0.189894
R8493 CS_BIAS.n52 CS_BIAS.n16 0.189894
R8494 CS_BIAS.n52 CS_BIAS.n51 0.189894
R8495 CS_BIAS.n51 CS_BIAS.n50 0.189894
R8496 CS_BIAS.n50 CS_BIAS.n18 0.189894
R8497 CS_BIAS.n45 CS_BIAS.n18 0.189894
R8498 CS_BIAS.n45 CS_BIAS.n44 0.189894
R8499 CS_BIAS.n44 CS_BIAS.n43 0.189894
R8500 CS_BIAS.n43 CS_BIAS.n20 0.189894
R8501 CS_BIAS.n39 CS_BIAS.n20 0.189894
R8502 CS_BIAS.n39 CS_BIAS.n38 0.189894
R8503 CS_BIAS.n38 CS_BIAS.n37 0.189894
R8504 CS_BIAS.n37 CS_BIAS.n22 0.189894
R8505 CS_BIAS.n33 CS_BIAS.n22 0.189894
R8506 CS_BIAS.n33 CS_BIAS.n32 0.189894
R8507 CS_BIAS.n32 CS_BIAS.n31 0.189894
R8508 CS_BIAS.n31 CS_BIAS.n24 0.189894
R8509 CS_BIAS.n27 CS_BIAS.n24 0.189894
R8510 CS_BIAS.n215 CS_BIAS.n0 0.189894
R8511 CS_BIAS.n215 CS_BIAS.n214 0.189894
R8512 CS_BIAS.n214 CS_BIAS.n213 0.189894
R8513 CS_BIAS.n213 CS_BIAS.n2 0.189894
R8514 CS_BIAS.n209 CS_BIAS.n2 0.189894
R8515 CS_BIAS.n209 CS_BIAS.n208 0.189894
R8516 CS_BIAS.n208 CS_BIAS.n207 0.189894
R8517 CS_BIAS.n207 CS_BIAS.n4 0.189894
R8518 CS_BIAS.n203 CS_BIAS.n4 0.189894
R8519 CS_BIAS.n203 CS_BIAS.n202 0.189894
R8520 CS_BIAS.n202 CS_BIAS.n201 0.189894
R8521 CS_BIAS.n201 CS_BIAS.n6 0.189894
R8522 CS_BIAS.n196 CS_BIAS.n6 0.189894
R8523 CS_BIAS.n196 CS_BIAS.n195 0.189894
R8524 CS_BIAS.n195 CS_BIAS.n194 0.189894
R8525 CS_BIAS.n194 CS_BIAS.n8 0.189894
R8526 CS_BIAS.n190 CS_BIAS.n8 0.189894
R8527 CS_BIAS.n190 CS_BIAS.n189 0.189894
R8528 CS_BIAS.n189 CS_BIAS.n188 0.189894
R8529 CS_BIAS.n188 CS_BIAS.n10 0.189894
R8530 CS_BIAS.n184 CS_BIAS.n10 0.189894
R8531 CS_BIAS.n184 CS_BIAS.n183 0.189894
R8532 CS_BIAS.n183 CS_BIAS.n182 0.189894
R8533 CS_BIAS.n182 CS_BIAS.n12 0.189894
R8534 CS_BIAS.n177 CS_BIAS.n12 0.189894
R8535 CS_BIAS.n177 CS_BIAS.n176 0.189894
R8536 CS_BIAS.n176 CS_BIAS.n175 0.189894
R8537 CS_BIAS.n175 CS_BIAS.n14 0.189894
R8538 CS_BIAS.n171 CS_BIAS.n14 0.189894
R8539 CS_BIAS.n171 CS_BIAS.n170 0.189894
R8540 CS_BIAS.n575 CS_BIAS.n572 0.189894
R8541 CS_BIAS.n579 CS_BIAS.n572 0.189894
R8542 CS_BIAS.n580 CS_BIAS.n579 0.189894
R8543 CS_BIAS.n581 CS_BIAS.n580 0.189894
R8544 CS_BIAS.n581 CS_BIAS.n570 0.189894
R8545 CS_BIAS.n585 CS_BIAS.n570 0.189894
R8546 CS_BIAS.n586 CS_BIAS.n585 0.189894
R8547 CS_BIAS.n587 CS_BIAS.n586 0.189894
R8548 CS_BIAS.n587 CS_BIAS.n568 0.189894
R8549 CS_BIAS.n591 CS_BIAS.n568 0.189894
R8550 CS_BIAS.n592 CS_BIAS.n591 0.189894
R8551 CS_BIAS.n593 CS_BIAS.n592 0.189894
R8552 CS_BIAS.n593 CS_BIAS.n566 0.189894
R8553 CS_BIAS.n598 CS_BIAS.n566 0.189894
R8554 CS_BIAS.n599 CS_BIAS.n598 0.189894
R8555 CS_BIAS.n600 CS_BIAS.n599 0.189894
R8556 CS_BIAS.n600 CS_BIAS.n564 0.189894
R8557 CS_BIAS.n604 CS_BIAS.n564 0.189894
R8558 CS_BIAS.n605 CS_BIAS.n604 0.189894
R8559 CS_BIAS.n606 CS_BIAS.n605 0.189894
R8560 CS_BIAS.n606 CS_BIAS.n562 0.189894
R8561 CS_BIAS.n610 CS_BIAS.n562 0.189894
R8562 CS_BIAS.n611 CS_BIAS.n610 0.189894
R8563 CS_BIAS.n612 CS_BIAS.n611 0.189894
R8564 CS_BIAS.n612 CS_BIAS.n560 0.189894
R8565 CS_BIAS.n617 CS_BIAS.n560 0.189894
R8566 CS_BIAS.n618 CS_BIAS.n617 0.189894
R8567 CS_BIAS.n619 CS_BIAS.n618 0.189894
R8568 CS_BIAS.n619 CS_BIAS.n558 0.189894
R8569 CS_BIAS.n623 CS_BIAS.n558 0.189894
R8570 CS_BIAS.n624 CS_BIAS.n623 0.189894
R8571 CS_BIAS.n625 CS_BIAS.n624 0.189894
R8572 CS_BIAS.n625 CS_BIAS.n556 0.189894
R8573 CS_BIAS.n629 CS_BIAS.n556 0.189894
R8574 CS_BIAS.n630 CS_BIAS.n629 0.189894
R8575 CS_BIAS.n631 CS_BIAS.n630 0.189894
R8576 CS_BIAS.n631 CS_BIAS.n554 0.189894
R8577 CS_BIAS.n636 CS_BIAS.n554 0.189894
R8578 CS_BIAS.n637 CS_BIAS.n636 0.189894
R8579 CS_BIAS.n638 CS_BIAS.n637 0.189894
R8580 CS_BIAS.n638 CS_BIAS.n552 0.189894
R8581 CS_BIAS.n642 CS_BIAS.n552 0.189894
R8582 CS_BIAS.n643 CS_BIAS.n642 0.189894
R8583 CS_BIAS.n644 CS_BIAS.n643 0.189894
R8584 CS_BIAS.n644 CS_BIAS.n550 0.189894
R8585 CS_BIAS.n648 CS_BIAS.n550 0.189894
R8586 CS_BIAS.n649 CS_BIAS.n648 0.189894
R8587 CS_BIAS.n650 CS_BIAS.n649 0.189894
R8588 CS_BIAS.n650 CS_BIAS.n548 0.189894
R8589 CS_BIAS.n414 CS_BIAS.n411 0.189894
R8590 CS_BIAS.n418 CS_BIAS.n411 0.189894
R8591 CS_BIAS.n419 CS_BIAS.n418 0.189894
R8592 CS_BIAS.n420 CS_BIAS.n419 0.189894
R8593 CS_BIAS.n420 CS_BIAS.n409 0.189894
R8594 CS_BIAS.n424 CS_BIAS.n409 0.189894
R8595 CS_BIAS.n425 CS_BIAS.n424 0.189894
R8596 CS_BIAS.n426 CS_BIAS.n425 0.189894
R8597 CS_BIAS.n426 CS_BIAS.n407 0.189894
R8598 CS_BIAS.n430 CS_BIAS.n407 0.189894
R8599 CS_BIAS.n431 CS_BIAS.n430 0.189894
R8600 CS_BIAS.n432 CS_BIAS.n431 0.189894
R8601 CS_BIAS.n432 CS_BIAS.n405 0.189894
R8602 CS_BIAS.n437 CS_BIAS.n405 0.189894
R8603 CS_BIAS.n438 CS_BIAS.n437 0.189894
R8604 CS_BIAS.n439 CS_BIAS.n438 0.189894
R8605 CS_BIAS.n439 CS_BIAS.n403 0.189894
R8606 CS_BIAS.n443 CS_BIAS.n403 0.189894
R8607 CS_BIAS.n444 CS_BIAS.n443 0.189894
R8608 CS_BIAS.n445 CS_BIAS.n444 0.189894
R8609 CS_BIAS.n445 CS_BIAS.n401 0.189894
R8610 CS_BIAS.n449 CS_BIAS.n401 0.189894
R8611 CS_BIAS.n450 CS_BIAS.n449 0.189894
R8612 CS_BIAS.n451 CS_BIAS.n450 0.189894
R8613 CS_BIAS.n451 CS_BIAS.n399 0.189894
R8614 CS_BIAS.n456 CS_BIAS.n399 0.189894
R8615 CS_BIAS.n457 CS_BIAS.n456 0.189894
R8616 CS_BIAS.n458 CS_BIAS.n457 0.189894
R8617 CS_BIAS.n458 CS_BIAS.n397 0.189894
R8618 CS_BIAS.n462 CS_BIAS.n397 0.189894
R8619 CS_BIAS.n463 CS_BIAS.n462 0.189894
R8620 CS_BIAS.n464 CS_BIAS.n463 0.189894
R8621 CS_BIAS.n464 CS_BIAS.n395 0.189894
R8622 CS_BIAS.n468 CS_BIAS.n395 0.189894
R8623 CS_BIAS.n469 CS_BIAS.n468 0.189894
R8624 CS_BIAS.n470 CS_BIAS.n469 0.189894
R8625 CS_BIAS.n470 CS_BIAS.n393 0.189894
R8626 CS_BIAS.n475 CS_BIAS.n393 0.189894
R8627 CS_BIAS.n476 CS_BIAS.n475 0.189894
R8628 CS_BIAS.n477 CS_BIAS.n476 0.189894
R8629 CS_BIAS.n477 CS_BIAS.n391 0.189894
R8630 CS_BIAS.n481 CS_BIAS.n391 0.189894
R8631 CS_BIAS.n482 CS_BIAS.n481 0.189894
R8632 CS_BIAS.n483 CS_BIAS.n482 0.189894
R8633 CS_BIAS.n483 CS_BIAS.n389 0.189894
R8634 CS_BIAS.n487 CS_BIAS.n389 0.189894
R8635 CS_BIAS.n488 CS_BIAS.n487 0.189894
R8636 CS_BIAS.n489 CS_BIAS.n488 0.189894
R8637 CS_BIAS.n489 CS_BIAS.n387 0.189894
R8638 CS_BIAS.n355 CS_BIAS.n352 0.189894
R8639 CS_BIAS.n359 CS_BIAS.n352 0.189894
R8640 CS_BIAS.n360 CS_BIAS.n359 0.189894
R8641 CS_BIAS.n361 CS_BIAS.n360 0.189894
R8642 CS_BIAS.n361 CS_BIAS.n350 0.189894
R8643 CS_BIAS.n365 CS_BIAS.n350 0.189894
R8644 CS_BIAS.n366 CS_BIAS.n365 0.189894
R8645 CS_BIAS.n367 CS_BIAS.n366 0.189894
R8646 CS_BIAS.n367 CS_BIAS.n348 0.189894
R8647 CS_BIAS.n371 CS_BIAS.n348 0.189894
R8648 CS_BIAS.n372 CS_BIAS.n371 0.189894
R8649 CS_BIAS.n373 CS_BIAS.n372 0.189894
R8650 CS_BIAS.n373 CS_BIAS.n346 0.189894
R8651 CS_BIAS.n378 CS_BIAS.n346 0.189894
R8652 CS_BIAS.n379 CS_BIAS.n378 0.189894
R8653 CS_BIAS.n380 CS_BIAS.n379 0.189894
R8654 CS_BIAS.n380 CS_BIAS.n344 0.189894
R8655 CS_BIAS.n384 CS_BIAS.n344 0.189894
R8656 CS_BIAS.n499 CS_BIAS.n498 0.189894
R8657 CS_BIAS.n499 CS_BIAS.n342 0.189894
R8658 CS_BIAS.n503 CS_BIAS.n342 0.189894
R8659 CS_BIAS.n504 CS_BIAS.n503 0.189894
R8660 CS_BIAS.n505 CS_BIAS.n504 0.189894
R8661 CS_BIAS.n505 CS_BIAS.n340 0.189894
R8662 CS_BIAS.n510 CS_BIAS.n340 0.189894
R8663 CS_BIAS.n511 CS_BIAS.n510 0.189894
R8664 CS_BIAS.n512 CS_BIAS.n511 0.189894
R8665 CS_BIAS.n512 CS_BIAS.n338 0.189894
R8666 CS_BIAS.n516 CS_BIAS.n338 0.189894
R8667 CS_BIAS.n517 CS_BIAS.n516 0.189894
R8668 CS_BIAS.n518 CS_BIAS.n517 0.189894
R8669 CS_BIAS.n518 CS_BIAS.n336 0.189894
R8670 CS_BIAS.n522 CS_BIAS.n336 0.189894
R8671 CS_BIAS.n523 CS_BIAS.n522 0.189894
R8672 CS_BIAS.n524 CS_BIAS.n523 0.189894
R8673 CS_BIAS.n524 CS_BIAS.n334 0.189894
R8674 CS_BIAS.n529 CS_BIAS.n334 0.189894
R8675 CS_BIAS.n530 CS_BIAS.n529 0.189894
R8676 CS_BIAS.n531 CS_BIAS.n530 0.189894
R8677 CS_BIAS.n531 CS_BIAS.n332 0.189894
R8678 CS_BIAS.n535 CS_BIAS.n332 0.189894
R8679 CS_BIAS.n536 CS_BIAS.n535 0.189894
R8680 CS_BIAS.n537 CS_BIAS.n536 0.189894
R8681 CS_BIAS.n537 CS_BIAS.n330 0.189894
R8682 CS_BIAS.n541 CS_BIAS.n330 0.189894
R8683 CS_BIAS.n542 CS_BIAS.n541 0.189894
R8684 CS_BIAS.n543 CS_BIAS.n542 0.189894
R8685 CS_BIAS.n543 CS_BIAS.n328 0.189894
R8686 CS_BIAS.n169 CS_BIAS.n56 0.0762576
R8687 CS_BIAS.n170 CS_BIAS.n169 0.0762576
R8688 CS_BIAS.n497 CS_BIAS.n384 0.0762576
R8689 CS_BIAS.n498 CS_BIAS.n497 0.0762576
R8690 GND.n9323 GND.n9322 2247.06
R8691 GND.n8179 GND.n8178 1108.29
R8692 GND.n9611 GND.n481 816.83
R8693 GND.n9569 GND.n477 816.83
R8694 GND.n3357 GND.n3305 816.83
R8695 GND.n7255 GND.n3359 816.83
R8696 GND.n7923 GND.n1776 816.83
R8697 GND.n7925 GND.n1770 816.83
R8698 GND.n1510 GND.n1463 816.83
R8699 GND.n8149 GND.n1474 816.83
R8700 GND.n7873 GND.n1774 771.183
R8701 GND.n7836 GND.n1772 771.183
R8702 GND.n1511 GND.n1465 771.183
R8703 GND.n8096 GND.n8095 771.183
R8704 GND.n7292 GND.n3313 771.183
R8705 GND.n7258 GND.n7257 771.183
R8706 GND.n9566 GND.n479 771.183
R8707 GND.n9613 GND.n475 771.183
R8708 GND.n8285 GND.n1319 742.355
R8709 GND.n9321 GND.n699 742.355
R8710 GND.n9462 GND.n617 742.355
R8711 GND.n8177 GND.n1428 742.355
R8712 GND.n6401 GND.n3231 727.939
R8713 GND.n7342 GND.n3229 727.939
R8714 GND.n3052 GND.n1848 727.939
R8715 GND.n7868 GND.n1837 727.939
R8716 GND.n8284 GND.n1318 693.51
R8717 GND.n8286 GND.n8285 585
R8718 GND.n8285 GND.n8284 585
R8719 GND.n1323 GND.n1322 585
R8720 GND.n8283 GND.n1323 585
R8721 GND.n8281 GND.n8280 585
R8722 GND.n8282 GND.n8281 585
R8723 GND.n8279 GND.n1325 585
R8724 GND.n1325 GND.n1324 585
R8725 GND.n8278 GND.n8277 585
R8726 GND.n8277 GND.n8276 585
R8727 GND.n1330 GND.n1329 585
R8728 GND.n8275 GND.n1330 585
R8729 GND.n8273 GND.n8272 585
R8730 GND.n8274 GND.n8273 585
R8731 GND.n8271 GND.n1332 585
R8732 GND.n1332 GND.n1331 585
R8733 GND.n8270 GND.n8269 585
R8734 GND.n8269 GND.n8268 585
R8735 GND.n1338 GND.n1337 585
R8736 GND.n8267 GND.n1338 585
R8737 GND.n8265 GND.n8264 585
R8738 GND.n8266 GND.n8265 585
R8739 GND.n8263 GND.n1340 585
R8740 GND.n1340 GND.n1339 585
R8741 GND.n8262 GND.n8261 585
R8742 GND.n8261 GND.n8260 585
R8743 GND.n1346 GND.n1345 585
R8744 GND.n8259 GND.n1346 585
R8745 GND.n8257 GND.n8256 585
R8746 GND.n8258 GND.n8257 585
R8747 GND.n8255 GND.n1348 585
R8748 GND.n1348 GND.n1347 585
R8749 GND.n8254 GND.n8253 585
R8750 GND.n8253 GND.n8252 585
R8751 GND.n1354 GND.n1353 585
R8752 GND.n8251 GND.n1354 585
R8753 GND.n8249 GND.n8248 585
R8754 GND.n8250 GND.n8249 585
R8755 GND.n8247 GND.n1356 585
R8756 GND.n1356 GND.n1355 585
R8757 GND.n8246 GND.n8245 585
R8758 GND.n8245 GND.n8244 585
R8759 GND.n1362 GND.n1361 585
R8760 GND.n8243 GND.n1362 585
R8761 GND.n8241 GND.n8240 585
R8762 GND.n8242 GND.n8241 585
R8763 GND.n8239 GND.n1364 585
R8764 GND.n1364 GND.n1363 585
R8765 GND.n8238 GND.n8237 585
R8766 GND.n8237 GND.n8236 585
R8767 GND.n1370 GND.n1369 585
R8768 GND.n8235 GND.n1370 585
R8769 GND.n8233 GND.n8232 585
R8770 GND.n8234 GND.n8233 585
R8771 GND.n8231 GND.n1372 585
R8772 GND.n1372 GND.n1371 585
R8773 GND.n8230 GND.n8229 585
R8774 GND.n8229 GND.n8228 585
R8775 GND.n1378 GND.n1377 585
R8776 GND.n8227 GND.n1378 585
R8777 GND.n8225 GND.n8224 585
R8778 GND.n8226 GND.n8225 585
R8779 GND.n8223 GND.n1380 585
R8780 GND.n1380 GND.n1379 585
R8781 GND.n8222 GND.n8221 585
R8782 GND.n8221 GND.n8220 585
R8783 GND.n1386 GND.n1385 585
R8784 GND.n8219 GND.n1386 585
R8785 GND.n8217 GND.n8216 585
R8786 GND.n8218 GND.n8217 585
R8787 GND.n8215 GND.n1388 585
R8788 GND.n1388 GND.n1387 585
R8789 GND.n8214 GND.n8213 585
R8790 GND.n8213 GND.n8212 585
R8791 GND.n1394 GND.n1393 585
R8792 GND.n8211 GND.n1394 585
R8793 GND.n8209 GND.n8208 585
R8794 GND.n8210 GND.n8209 585
R8795 GND.n8207 GND.n1396 585
R8796 GND.n1396 GND.n1395 585
R8797 GND.n8206 GND.n8205 585
R8798 GND.n8205 GND.n8204 585
R8799 GND.n1402 GND.n1401 585
R8800 GND.n8203 GND.n1402 585
R8801 GND.n8201 GND.n8200 585
R8802 GND.n8202 GND.n8201 585
R8803 GND.n8199 GND.n1404 585
R8804 GND.n1404 GND.n1403 585
R8805 GND.n8198 GND.n8197 585
R8806 GND.n8197 GND.n8196 585
R8807 GND.n1410 GND.n1409 585
R8808 GND.n8195 GND.n1410 585
R8809 GND.n8193 GND.n8192 585
R8810 GND.n8194 GND.n8193 585
R8811 GND.n8191 GND.n1412 585
R8812 GND.n1412 GND.n1411 585
R8813 GND.n8190 GND.n8189 585
R8814 GND.n8189 GND.n8188 585
R8815 GND.n1418 GND.n1417 585
R8816 GND.n8187 GND.n1418 585
R8817 GND.n8185 GND.n8184 585
R8818 GND.n8186 GND.n8185 585
R8819 GND.n8183 GND.n1420 585
R8820 GND.n1420 GND.n1419 585
R8821 GND.n8182 GND.n8181 585
R8822 GND.n8181 GND.n8180 585
R8823 GND.n1426 GND.n1425 585
R8824 GND.n8179 GND.n1426 585
R8825 GND.n1320 GND.n1319 585
R8826 GND.n1319 GND.n1318 585
R8827 GND.n8291 GND.n8290 585
R8828 GND.n8292 GND.n8291 585
R8829 GND.n1317 GND.n1316 585
R8830 GND.n8293 GND.n1317 585
R8831 GND.n8296 GND.n8295 585
R8832 GND.n8295 GND.n8294 585
R8833 GND.n1314 GND.n1313 585
R8834 GND.n1313 GND.n1312 585
R8835 GND.n8301 GND.n8300 585
R8836 GND.n8302 GND.n8301 585
R8837 GND.n1311 GND.n1310 585
R8838 GND.n8303 GND.n1311 585
R8839 GND.n8306 GND.n8305 585
R8840 GND.n8305 GND.n8304 585
R8841 GND.n1308 GND.n1307 585
R8842 GND.n1307 GND.n1306 585
R8843 GND.n8311 GND.n8310 585
R8844 GND.n8312 GND.n8311 585
R8845 GND.n1305 GND.n1304 585
R8846 GND.n8313 GND.n1305 585
R8847 GND.n8316 GND.n8315 585
R8848 GND.n8315 GND.n8314 585
R8849 GND.n1302 GND.n1301 585
R8850 GND.n1301 GND.n1300 585
R8851 GND.n8321 GND.n8320 585
R8852 GND.n8322 GND.n8321 585
R8853 GND.n1299 GND.n1298 585
R8854 GND.n8323 GND.n1299 585
R8855 GND.n8326 GND.n8325 585
R8856 GND.n8325 GND.n8324 585
R8857 GND.n1296 GND.n1295 585
R8858 GND.n1295 GND.n1294 585
R8859 GND.n8331 GND.n8330 585
R8860 GND.n8332 GND.n8331 585
R8861 GND.n1293 GND.n1292 585
R8862 GND.n8333 GND.n1293 585
R8863 GND.n8336 GND.n8335 585
R8864 GND.n8335 GND.n8334 585
R8865 GND.n1290 GND.n1289 585
R8866 GND.n1289 GND.n1288 585
R8867 GND.n8341 GND.n8340 585
R8868 GND.n8342 GND.n8341 585
R8869 GND.n1287 GND.n1286 585
R8870 GND.n8343 GND.n1287 585
R8871 GND.n8346 GND.n8345 585
R8872 GND.n8345 GND.n8344 585
R8873 GND.n1284 GND.n1283 585
R8874 GND.n1283 GND.n1282 585
R8875 GND.n8351 GND.n8350 585
R8876 GND.n8352 GND.n8351 585
R8877 GND.n1281 GND.n1280 585
R8878 GND.n8353 GND.n1281 585
R8879 GND.n8356 GND.n8355 585
R8880 GND.n8355 GND.n8354 585
R8881 GND.n1278 GND.n1277 585
R8882 GND.n1277 GND.n1276 585
R8883 GND.n8361 GND.n8360 585
R8884 GND.n8362 GND.n8361 585
R8885 GND.n1275 GND.n1274 585
R8886 GND.n8363 GND.n1275 585
R8887 GND.n8366 GND.n8365 585
R8888 GND.n8365 GND.n8364 585
R8889 GND.n1272 GND.n1271 585
R8890 GND.n1271 GND.n1270 585
R8891 GND.n8371 GND.n8370 585
R8892 GND.n8372 GND.n8371 585
R8893 GND.n1269 GND.n1268 585
R8894 GND.n8373 GND.n1269 585
R8895 GND.n8376 GND.n8375 585
R8896 GND.n8375 GND.n8374 585
R8897 GND.n1266 GND.n1265 585
R8898 GND.n1265 GND.n1264 585
R8899 GND.n8381 GND.n8380 585
R8900 GND.n8382 GND.n8381 585
R8901 GND.n1263 GND.n1262 585
R8902 GND.n8383 GND.n1263 585
R8903 GND.n8386 GND.n8385 585
R8904 GND.n8385 GND.n8384 585
R8905 GND.n1260 GND.n1259 585
R8906 GND.n1259 GND.n1258 585
R8907 GND.n8391 GND.n8390 585
R8908 GND.n8392 GND.n8391 585
R8909 GND.n1257 GND.n1256 585
R8910 GND.n8393 GND.n1257 585
R8911 GND.n8396 GND.n8395 585
R8912 GND.n8395 GND.n8394 585
R8913 GND.n1254 GND.n1253 585
R8914 GND.n1253 GND.n1252 585
R8915 GND.n8401 GND.n8400 585
R8916 GND.n8402 GND.n8401 585
R8917 GND.n1251 GND.n1250 585
R8918 GND.n8403 GND.n1251 585
R8919 GND.n8406 GND.n8405 585
R8920 GND.n8405 GND.n8404 585
R8921 GND.n1248 GND.n1247 585
R8922 GND.n1247 GND.n1246 585
R8923 GND.n8411 GND.n8410 585
R8924 GND.n8412 GND.n8411 585
R8925 GND.n1245 GND.n1244 585
R8926 GND.n8413 GND.n1245 585
R8927 GND.n8416 GND.n8415 585
R8928 GND.n8415 GND.n8414 585
R8929 GND.n1242 GND.n1241 585
R8930 GND.n1241 GND.n1240 585
R8931 GND.n8421 GND.n8420 585
R8932 GND.n8422 GND.n8421 585
R8933 GND.n1239 GND.n1238 585
R8934 GND.n8423 GND.n1239 585
R8935 GND.n8426 GND.n8425 585
R8936 GND.n8425 GND.n8424 585
R8937 GND.n1236 GND.n1235 585
R8938 GND.n1235 GND.n1234 585
R8939 GND.n8431 GND.n8430 585
R8940 GND.n8432 GND.n8431 585
R8941 GND.n1233 GND.n1232 585
R8942 GND.n8433 GND.n1233 585
R8943 GND.n8436 GND.n8435 585
R8944 GND.n8435 GND.n8434 585
R8945 GND.n1230 GND.n1229 585
R8946 GND.n1229 GND.n1228 585
R8947 GND.n8441 GND.n8440 585
R8948 GND.n8442 GND.n8441 585
R8949 GND.n1227 GND.n1226 585
R8950 GND.n8443 GND.n1227 585
R8951 GND.n8446 GND.n8445 585
R8952 GND.n8445 GND.n8444 585
R8953 GND.n1224 GND.n1223 585
R8954 GND.n1223 GND.n1222 585
R8955 GND.n8451 GND.n8450 585
R8956 GND.n8452 GND.n8451 585
R8957 GND.n1221 GND.n1220 585
R8958 GND.n8453 GND.n1221 585
R8959 GND.n8456 GND.n8455 585
R8960 GND.n8455 GND.n8454 585
R8961 GND.n1218 GND.n1217 585
R8962 GND.n1217 GND.n1216 585
R8963 GND.n8461 GND.n8460 585
R8964 GND.n8462 GND.n8461 585
R8965 GND.n1215 GND.n1214 585
R8966 GND.n8463 GND.n1215 585
R8967 GND.n8466 GND.n8465 585
R8968 GND.n8465 GND.n8464 585
R8969 GND.n1212 GND.n1211 585
R8970 GND.n1211 GND.n1210 585
R8971 GND.n8471 GND.n8470 585
R8972 GND.n8472 GND.n8471 585
R8973 GND.n1209 GND.n1208 585
R8974 GND.n8473 GND.n1209 585
R8975 GND.n8476 GND.n8475 585
R8976 GND.n8475 GND.n8474 585
R8977 GND.n1206 GND.n1205 585
R8978 GND.n1205 GND.n1204 585
R8979 GND.n8481 GND.n8480 585
R8980 GND.n8482 GND.n8481 585
R8981 GND.n1203 GND.n1202 585
R8982 GND.n8483 GND.n1203 585
R8983 GND.n8486 GND.n8485 585
R8984 GND.n8485 GND.n8484 585
R8985 GND.n1200 GND.n1199 585
R8986 GND.n1199 GND.n1198 585
R8987 GND.n8491 GND.n8490 585
R8988 GND.n8492 GND.n8491 585
R8989 GND.n1197 GND.n1196 585
R8990 GND.n8493 GND.n1197 585
R8991 GND.n8496 GND.n8495 585
R8992 GND.n8495 GND.n8494 585
R8993 GND.n1194 GND.n1193 585
R8994 GND.n1193 GND.n1192 585
R8995 GND.n8501 GND.n8500 585
R8996 GND.n8502 GND.n8501 585
R8997 GND.n1191 GND.n1190 585
R8998 GND.n8503 GND.n1191 585
R8999 GND.n8506 GND.n8505 585
R9000 GND.n8505 GND.n8504 585
R9001 GND.n1188 GND.n1187 585
R9002 GND.n1187 GND.n1186 585
R9003 GND.n8511 GND.n8510 585
R9004 GND.n8512 GND.n8511 585
R9005 GND.n1185 GND.n1184 585
R9006 GND.n8513 GND.n1185 585
R9007 GND.n8516 GND.n8515 585
R9008 GND.n8515 GND.n8514 585
R9009 GND.n1182 GND.n1181 585
R9010 GND.n1181 GND.n1180 585
R9011 GND.n8521 GND.n8520 585
R9012 GND.n8522 GND.n8521 585
R9013 GND.n1179 GND.n1178 585
R9014 GND.n8523 GND.n1179 585
R9015 GND.n8526 GND.n8525 585
R9016 GND.n8525 GND.n8524 585
R9017 GND.n1176 GND.n1175 585
R9018 GND.n1175 GND.n1174 585
R9019 GND.n8531 GND.n8530 585
R9020 GND.n8532 GND.n8531 585
R9021 GND.n1173 GND.n1172 585
R9022 GND.n8533 GND.n1173 585
R9023 GND.n8536 GND.n8535 585
R9024 GND.n8535 GND.n8534 585
R9025 GND.n1170 GND.n1169 585
R9026 GND.n1169 GND.n1168 585
R9027 GND.n8541 GND.n8540 585
R9028 GND.n8542 GND.n8541 585
R9029 GND.n1167 GND.n1166 585
R9030 GND.n8543 GND.n1167 585
R9031 GND.n8546 GND.n8545 585
R9032 GND.n8545 GND.n8544 585
R9033 GND.n1164 GND.n1163 585
R9034 GND.n1163 GND.n1162 585
R9035 GND.n8551 GND.n8550 585
R9036 GND.n8552 GND.n8551 585
R9037 GND.n1161 GND.n1160 585
R9038 GND.n8553 GND.n1161 585
R9039 GND.n8556 GND.n8555 585
R9040 GND.n8555 GND.n8554 585
R9041 GND.n1158 GND.n1157 585
R9042 GND.n1157 GND.n1156 585
R9043 GND.n8561 GND.n8560 585
R9044 GND.n8562 GND.n8561 585
R9045 GND.n1155 GND.n1154 585
R9046 GND.n8563 GND.n1155 585
R9047 GND.n8566 GND.n8565 585
R9048 GND.n8565 GND.n8564 585
R9049 GND.n1152 GND.n1151 585
R9050 GND.n1151 GND.n1150 585
R9051 GND.n8571 GND.n8570 585
R9052 GND.n8572 GND.n8571 585
R9053 GND.n1149 GND.n1148 585
R9054 GND.n8573 GND.n1149 585
R9055 GND.n8576 GND.n8575 585
R9056 GND.n8575 GND.n8574 585
R9057 GND.n1146 GND.n1145 585
R9058 GND.n1145 GND.n1144 585
R9059 GND.n8581 GND.n8580 585
R9060 GND.n8582 GND.n8581 585
R9061 GND.n1143 GND.n1142 585
R9062 GND.n8583 GND.n1143 585
R9063 GND.n8586 GND.n8585 585
R9064 GND.n8585 GND.n8584 585
R9065 GND.n1140 GND.n1139 585
R9066 GND.n1139 GND.n1138 585
R9067 GND.n8591 GND.n8590 585
R9068 GND.n8592 GND.n8591 585
R9069 GND.n1137 GND.n1136 585
R9070 GND.n8593 GND.n1137 585
R9071 GND.n8596 GND.n8595 585
R9072 GND.n8595 GND.n8594 585
R9073 GND.n1134 GND.n1133 585
R9074 GND.n1133 GND.n1132 585
R9075 GND.n8601 GND.n8600 585
R9076 GND.n8602 GND.n8601 585
R9077 GND.n1131 GND.n1130 585
R9078 GND.n8603 GND.n1131 585
R9079 GND.n8606 GND.n8605 585
R9080 GND.n8605 GND.n8604 585
R9081 GND.n1128 GND.n1127 585
R9082 GND.n1127 GND.n1126 585
R9083 GND.n8611 GND.n8610 585
R9084 GND.n8612 GND.n8611 585
R9085 GND.n1125 GND.n1124 585
R9086 GND.n8613 GND.n1125 585
R9087 GND.n8616 GND.n8615 585
R9088 GND.n8615 GND.n8614 585
R9089 GND.n1122 GND.n1121 585
R9090 GND.n1121 GND.n1120 585
R9091 GND.n8621 GND.n8620 585
R9092 GND.n8622 GND.n8621 585
R9093 GND.n1119 GND.n1118 585
R9094 GND.n8623 GND.n1119 585
R9095 GND.n8626 GND.n8625 585
R9096 GND.n8625 GND.n8624 585
R9097 GND.n1116 GND.n1115 585
R9098 GND.n1115 GND.n1114 585
R9099 GND.n8631 GND.n8630 585
R9100 GND.n8632 GND.n8631 585
R9101 GND.n1113 GND.n1112 585
R9102 GND.n8633 GND.n1113 585
R9103 GND.n8636 GND.n8635 585
R9104 GND.n8635 GND.n8634 585
R9105 GND.n1110 GND.n1109 585
R9106 GND.n1109 GND.n1108 585
R9107 GND.n8641 GND.n8640 585
R9108 GND.n8642 GND.n8641 585
R9109 GND.n1107 GND.n1106 585
R9110 GND.n8643 GND.n1107 585
R9111 GND.n8646 GND.n8645 585
R9112 GND.n8645 GND.n8644 585
R9113 GND.n1104 GND.n1103 585
R9114 GND.n1103 GND.n1102 585
R9115 GND.n8651 GND.n8650 585
R9116 GND.n8652 GND.n8651 585
R9117 GND.n1101 GND.n1100 585
R9118 GND.n8653 GND.n1101 585
R9119 GND.n8656 GND.n8655 585
R9120 GND.n8655 GND.n8654 585
R9121 GND.n1098 GND.n1097 585
R9122 GND.n1097 GND.n1096 585
R9123 GND.n8661 GND.n8660 585
R9124 GND.n8662 GND.n8661 585
R9125 GND.n1095 GND.n1094 585
R9126 GND.n8663 GND.n1095 585
R9127 GND.n8666 GND.n8665 585
R9128 GND.n8665 GND.n8664 585
R9129 GND.n1092 GND.n1091 585
R9130 GND.n1091 GND.n1090 585
R9131 GND.n8671 GND.n8670 585
R9132 GND.n8672 GND.n8671 585
R9133 GND.n1089 GND.n1088 585
R9134 GND.n8673 GND.n1089 585
R9135 GND.n8676 GND.n8675 585
R9136 GND.n8675 GND.n8674 585
R9137 GND.n1086 GND.n1085 585
R9138 GND.n1085 GND.n1084 585
R9139 GND.n8681 GND.n8680 585
R9140 GND.n8682 GND.n8681 585
R9141 GND.n1083 GND.n1082 585
R9142 GND.n8683 GND.n1083 585
R9143 GND.n8686 GND.n8685 585
R9144 GND.n8685 GND.n8684 585
R9145 GND.n1080 GND.n1079 585
R9146 GND.n1079 GND.n1078 585
R9147 GND.n8691 GND.n8690 585
R9148 GND.n8692 GND.n8691 585
R9149 GND.n1077 GND.n1076 585
R9150 GND.n8693 GND.n1077 585
R9151 GND.n8696 GND.n8695 585
R9152 GND.n8695 GND.n8694 585
R9153 GND.n1074 GND.n1073 585
R9154 GND.n1073 GND.n1072 585
R9155 GND.n8701 GND.n8700 585
R9156 GND.n8702 GND.n8701 585
R9157 GND.n1071 GND.n1070 585
R9158 GND.n8703 GND.n1071 585
R9159 GND.n8706 GND.n8705 585
R9160 GND.n8705 GND.n8704 585
R9161 GND.n1068 GND.n1067 585
R9162 GND.n1067 GND.n1066 585
R9163 GND.n8711 GND.n8710 585
R9164 GND.n8712 GND.n8711 585
R9165 GND.n1065 GND.n1064 585
R9166 GND.n8713 GND.n1065 585
R9167 GND.n8716 GND.n8715 585
R9168 GND.n8715 GND.n8714 585
R9169 GND.n1062 GND.n1061 585
R9170 GND.n1061 GND.n1060 585
R9171 GND.n8721 GND.n8720 585
R9172 GND.n8722 GND.n8721 585
R9173 GND.n1059 GND.n1058 585
R9174 GND.n8723 GND.n1059 585
R9175 GND.n8726 GND.n8725 585
R9176 GND.n8725 GND.n8724 585
R9177 GND.n1056 GND.n1055 585
R9178 GND.n1055 GND.n1054 585
R9179 GND.n8731 GND.n8730 585
R9180 GND.n8732 GND.n8731 585
R9181 GND.n1053 GND.n1052 585
R9182 GND.n8733 GND.n1053 585
R9183 GND.n8736 GND.n8735 585
R9184 GND.n8735 GND.n8734 585
R9185 GND.n1050 GND.n1049 585
R9186 GND.n1049 GND.n1048 585
R9187 GND.n8741 GND.n8740 585
R9188 GND.n8742 GND.n8741 585
R9189 GND.n1047 GND.n1046 585
R9190 GND.n8743 GND.n1047 585
R9191 GND.n8746 GND.n8745 585
R9192 GND.n8745 GND.n8744 585
R9193 GND.n1044 GND.n1043 585
R9194 GND.n1043 GND.n1042 585
R9195 GND.n8751 GND.n8750 585
R9196 GND.n8752 GND.n8751 585
R9197 GND.n1041 GND.n1040 585
R9198 GND.n8753 GND.n1041 585
R9199 GND.n8756 GND.n8755 585
R9200 GND.n8755 GND.n8754 585
R9201 GND.n1038 GND.n1037 585
R9202 GND.n1037 GND.n1036 585
R9203 GND.n8761 GND.n8760 585
R9204 GND.n8762 GND.n8761 585
R9205 GND.n1035 GND.n1034 585
R9206 GND.n8763 GND.n1035 585
R9207 GND.n8766 GND.n8765 585
R9208 GND.n8765 GND.n8764 585
R9209 GND.n1032 GND.n1031 585
R9210 GND.n1031 GND.n1030 585
R9211 GND.n8771 GND.n8770 585
R9212 GND.n8772 GND.n8771 585
R9213 GND.n1029 GND.n1028 585
R9214 GND.n8773 GND.n1029 585
R9215 GND.n8776 GND.n8775 585
R9216 GND.n8775 GND.n8774 585
R9217 GND.n1026 GND.n1025 585
R9218 GND.n1025 GND.n1024 585
R9219 GND.n8781 GND.n8780 585
R9220 GND.n8782 GND.n8781 585
R9221 GND.n1023 GND.n1022 585
R9222 GND.n8783 GND.n1023 585
R9223 GND.n8786 GND.n8785 585
R9224 GND.n8785 GND.n8784 585
R9225 GND.n1020 GND.n1019 585
R9226 GND.n1019 GND.n1018 585
R9227 GND.n8791 GND.n8790 585
R9228 GND.n8792 GND.n8791 585
R9229 GND.n1017 GND.n1016 585
R9230 GND.n8793 GND.n1017 585
R9231 GND.n8796 GND.n8795 585
R9232 GND.n8795 GND.n8794 585
R9233 GND.n1014 GND.n1013 585
R9234 GND.n1013 GND.n1012 585
R9235 GND.n8801 GND.n8800 585
R9236 GND.n8802 GND.n8801 585
R9237 GND.n1011 GND.n1010 585
R9238 GND.n8803 GND.n1011 585
R9239 GND.n8806 GND.n8805 585
R9240 GND.n8805 GND.n8804 585
R9241 GND.n1008 GND.n1007 585
R9242 GND.n1007 GND.n1006 585
R9243 GND.n8811 GND.n8810 585
R9244 GND.n8812 GND.n8811 585
R9245 GND.n1005 GND.n1004 585
R9246 GND.n8813 GND.n1005 585
R9247 GND.n8816 GND.n8815 585
R9248 GND.n8815 GND.n8814 585
R9249 GND.n1002 GND.n1001 585
R9250 GND.n1001 GND.n1000 585
R9251 GND.n8821 GND.n8820 585
R9252 GND.n8822 GND.n8821 585
R9253 GND.n999 GND.n998 585
R9254 GND.n8823 GND.n999 585
R9255 GND.n8826 GND.n8825 585
R9256 GND.n8825 GND.n8824 585
R9257 GND.n996 GND.n995 585
R9258 GND.n995 GND.n994 585
R9259 GND.n8831 GND.n8830 585
R9260 GND.n8832 GND.n8831 585
R9261 GND.n993 GND.n992 585
R9262 GND.n8833 GND.n993 585
R9263 GND.n8836 GND.n8835 585
R9264 GND.n8835 GND.n8834 585
R9265 GND.n990 GND.n989 585
R9266 GND.n989 GND.n988 585
R9267 GND.n8841 GND.n8840 585
R9268 GND.n8842 GND.n8841 585
R9269 GND.n987 GND.n986 585
R9270 GND.n8843 GND.n987 585
R9271 GND.n8846 GND.n8845 585
R9272 GND.n8845 GND.n8844 585
R9273 GND.n984 GND.n983 585
R9274 GND.n983 GND.n982 585
R9275 GND.n8851 GND.n8850 585
R9276 GND.n8852 GND.n8851 585
R9277 GND.n981 GND.n980 585
R9278 GND.n8853 GND.n981 585
R9279 GND.n8856 GND.n8855 585
R9280 GND.n8855 GND.n8854 585
R9281 GND.n978 GND.n977 585
R9282 GND.n977 GND.n976 585
R9283 GND.n8861 GND.n8860 585
R9284 GND.n8862 GND.n8861 585
R9285 GND.n975 GND.n974 585
R9286 GND.n8863 GND.n975 585
R9287 GND.n8866 GND.n8865 585
R9288 GND.n8865 GND.n8864 585
R9289 GND.n972 GND.n971 585
R9290 GND.n971 GND.n970 585
R9291 GND.n8871 GND.n8870 585
R9292 GND.n8872 GND.n8871 585
R9293 GND.n969 GND.n968 585
R9294 GND.n8873 GND.n969 585
R9295 GND.n8876 GND.n8875 585
R9296 GND.n8875 GND.n8874 585
R9297 GND.n966 GND.n965 585
R9298 GND.n965 GND.n964 585
R9299 GND.n8881 GND.n8880 585
R9300 GND.n8882 GND.n8881 585
R9301 GND.n963 GND.n962 585
R9302 GND.n8883 GND.n963 585
R9303 GND.n8886 GND.n8885 585
R9304 GND.n8885 GND.n8884 585
R9305 GND.n960 GND.n959 585
R9306 GND.n959 GND.n958 585
R9307 GND.n8891 GND.n8890 585
R9308 GND.n8892 GND.n8891 585
R9309 GND.n957 GND.n956 585
R9310 GND.n8893 GND.n957 585
R9311 GND.n8896 GND.n8895 585
R9312 GND.n8895 GND.n8894 585
R9313 GND.n954 GND.n953 585
R9314 GND.n953 GND.n952 585
R9315 GND.n8901 GND.n8900 585
R9316 GND.n8902 GND.n8901 585
R9317 GND.n951 GND.n950 585
R9318 GND.n8903 GND.n951 585
R9319 GND.n8906 GND.n8905 585
R9320 GND.n8905 GND.n8904 585
R9321 GND.n948 GND.n947 585
R9322 GND.n947 GND.n946 585
R9323 GND.n8911 GND.n8910 585
R9324 GND.n8912 GND.n8911 585
R9325 GND.n945 GND.n944 585
R9326 GND.n8913 GND.n945 585
R9327 GND.n8916 GND.n8915 585
R9328 GND.n8915 GND.n8914 585
R9329 GND.n942 GND.n941 585
R9330 GND.n941 GND.n940 585
R9331 GND.n8921 GND.n8920 585
R9332 GND.n8922 GND.n8921 585
R9333 GND.n939 GND.n938 585
R9334 GND.n8923 GND.n939 585
R9335 GND.n8926 GND.n8925 585
R9336 GND.n8925 GND.n8924 585
R9337 GND.n936 GND.n935 585
R9338 GND.n935 GND.n934 585
R9339 GND.n8931 GND.n8930 585
R9340 GND.n8932 GND.n8931 585
R9341 GND.n933 GND.n932 585
R9342 GND.n8933 GND.n933 585
R9343 GND.n8936 GND.n8935 585
R9344 GND.n8935 GND.n8934 585
R9345 GND.n930 GND.n929 585
R9346 GND.n929 GND.n928 585
R9347 GND.n8941 GND.n8940 585
R9348 GND.n8942 GND.n8941 585
R9349 GND.n927 GND.n926 585
R9350 GND.n8943 GND.n927 585
R9351 GND.n8946 GND.n8945 585
R9352 GND.n8945 GND.n8944 585
R9353 GND.n924 GND.n923 585
R9354 GND.n923 GND.n922 585
R9355 GND.n8951 GND.n8950 585
R9356 GND.n8952 GND.n8951 585
R9357 GND.n921 GND.n920 585
R9358 GND.n8953 GND.n921 585
R9359 GND.n8956 GND.n8955 585
R9360 GND.n8955 GND.n8954 585
R9361 GND.n918 GND.n917 585
R9362 GND.n917 GND.n916 585
R9363 GND.n8961 GND.n8960 585
R9364 GND.n8962 GND.n8961 585
R9365 GND.n915 GND.n914 585
R9366 GND.n8963 GND.n915 585
R9367 GND.n8966 GND.n8965 585
R9368 GND.n8965 GND.n8964 585
R9369 GND.n912 GND.n911 585
R9370 GND.n911 GND.n910 585
R9371 GND.n8971 GND.n8970 585
R9372 GND.n8972 GND.n8971 585
R9373 GND.n909 GND.n908 585
R9374 GND.n8973 GND.n909 585
R9375 GND.n8976 GND.n8975 585
R9376 GND.n8975 GND.n8974 585
R9377 GND.n906 GND.n905 585
R9378 GND.n905 GND.n904 585
R9379 GND.n8981 GND.n8980 585
R9380 GND.n8982 GND.n8981 585
R9381 GND.n903 GND.n902 585
R9382 GND.n8983 GND.n903 585
R9383 GND.n8986 GND.n8985 585
R9384 GND.n8985 GND.n8984 585
R9385 GND.n900 GND.n899 585
R9386 GND.n899 GND.n898 585
R9387 GND.n8991 GND.n8990 585
R9388 GND.n8992 GND.n8991 585
R9389 GND.n897 GND.n896 585
R9390 GND.n8993 GND.n897 585
R9391 GND.n8996 GND.n8995 585
R9392 GND.n8995 GND.n8994 585
R9393 GND.n894 GND.n893 585
R9394 GND.n893 GND.n892 585
R9395 GND.n9001 GND.n9000 585
R9396 GND.n9002 GND.n9001 585
R9397 GND.n891 GND.n890 585
R9398 GND.n9003 GND.n891 585
R9399 GND.n9006 GND.n9005 585
R9400 GND.n9005 GND.n9004 585
R9401 GND.n888 GND.n887 585
R9402 GND.n887 GND.n886 585
R9403 GND.n9011 GND.n9010 585
R9404 GND.n9012 GND.n9011 585
R9405 GND.n885 GND.n884 585
R9406 GND.n9013 GND.n885 585
R9407 GND.n9016 GND.n9015 585
R9408 GND.n9015 GND.n9014 585
R9409 GND.n882 GND.n881 585
R9410 GND.n881 GND.n880 585
R9411 GND.n9021 GND.n9020 585
R9412 GND.n9022 GND.n9021 585
R9413 GND.n879 GND.n878 585
R9414 GND.n9023 GND.n879 585
R9415 GND.n9026 GND.n9025 585
R9416 GND.n9025 GND.n9024 585
R9417 GND.n876 GND.n875 585
R9418 GND.n875 GND.n874 585
R9419 GND.n9031 GND.n9030 585
R9420 GND.n9032 GND.n9031 585
R9421 GND.n873 GND.n872 585
R9422 GND.n9033 GND.n873 585
R9423 GND.n9036 GND.n9035 585
R9424 GND.n9035 GND.n9034 585
R9425 GND.n870 GND.n869 585
R9426 GND.n869 GND.n868 585
R9427 GND.n9041 GND.n9040 585
R9428 GND.n9042 GND.n9041 585
R9429 GND.n867 GND.n866 585
R9430 GND.n9043 GND.n867 585
R9431 GND.n9046 GND.n9045 585
R9432 GND.n9045 GND.n9044 585
R9433 GND.n864 GND.n863 585
R9434 GND.n863 GND.n862 585
R9435 GND.n9051 GND.n9050 585
R9436 GND.n9052 GND.n9051 585
R9437 GND.n861 GND.n860 585
R9438 GND.n9053 GND.n861 585
R9439 GND.n9056 GND.n9055 585
R9440 GND.n9055 GND.n9054 585
R9441 GND.n858 GND.n857 585
R9442 GND.n857 GND.n856 585
R9443 GND.n9061 GND.n9060 585
R9444 GND.n9062 GND.n9061 585
R9445 GND.n855 GND.n854 585
R9446 GND.n9063 GND.n855 585
R9447 GND.n9066 GND.n9065 585
R9448 GND.n9065 GND.n9064 585
R9449 GND.n852 GND.n851 585
R9450 GND.n851 GND.n850 585
R9451 GND.n9071 GND.n9070 585
R9452 GND.n9072 GND.n9071 585
R9453 GND.n849 GND.n848 585
R9454 GND.n9073 GND.n849 585
R9455 GND.n9076 GND.n9075 585
R9456 GND.n9075 GND.n9074 585
R9457 GND.n846 GND.n845 585
R9458 GND.n845 GND.n844 585
R9459 GND.n9081 GND.n9080 585
R9460 GND.n9082 GND.n9081 585
R9461 GND.n843 GND.n842 585
R9462 GND.n9083 GND.n843 585
R9463 GND.n9086 GND.n9085 585
R9464 GND.n9085 GND.n9084 585
R9465 GND.n840 GND.n839 585
R9466 GND.n839 GND.n838 585
R9467 GND.n9091 GND.n9090 585
R9468 GND.n9092 GND.n9091 585
R9469 GND.n837 GND.n836 585
R9470 GND.n9093 GND.n837 585
R9471 GND.n9096 GND.n9095 585
R9472 GND.n9095 GND.n9094 585
R9473 GND.n834 GND.n833 585
R9474 GND.n833 GND.n832 585
R9475 GND.n9101 GND.n9100 585
R9476 GND.n9102 GND.n9101 585
R9477 GND.n831 GND.n830 585
R9478 GND.n9103 GND.n831 585
R9479 GND.n9106 GND.n9105 585
R9480 GND.n9105 GND.n9104 585
R9481 GND.n828 GND.n827 585
R9482 GND.n827 GND.n826 585
R9483 GND.n9111 GND.n9110 585
R9484 GND.n9112 GND.n9111 585
R9485 GND.n825 GND.n824 585
R9486 GND.n9113 GND.n825 585
R9487 GND.n9116 GND.n9115 585
R9488 GND.n9115 GND.n9114 585
R9489 GND.n822 GND.n821 585
R9490 GND.n821 GND.n820 585
R9491 GND.n9121 GND.n9120 585
R9492 GND.n9122 GND.n9121 585
R9493 GND.n819 GND.n818 585
R9494 GND.n9123 GND.n819 585
R9495 GND.n9126 GND.n9125 585
R9496 GND.n9125 GND.n9124 585
R9497 GND.n816 GND.n815 585
R9498 GND.n815 GND.n814 585
R9499 GND.n9131 GND.n9130 585
R9500 GND.n9132 GND.n9131 585
R9501 GND.n813 GND.n812 585
R9502 GND.n9133 GND.n813 585
R9503 GND.n9136 GND.n9135 585
R9504 GND.n9135 GND.n9134 585
R9505 GND.n810 GND.n809 585
R9506 GND.n809 GND.n808 585
R9507 GND.n9141 GND.n9140 585
R9508 GND.n9142 GND.n9141 585
R9509 GND.n807 GND.n806 585
R9510 GND.n9143 GND.n807 585
R9511 GND.n9146 GND.n9145 585
R9512 GND.n9145 GND.n9144 585
R9513 GND.n804 GND.n803 585
R9514 GND.n803 GND.n802 585
R9515 GND.n9151 GND.n9150 585
R9516 GND.n9152 GND.n9151 585
R9517 GND.n801 GND.n800 585
R9518 GND.n9153 GND.n801 585
R9519 GND.n9156 GND.n9155 585
R9520 GND.n9155 GND.n9154 585
R9521 GND.n798 GND.n797 585
R9522 GND.n797 GND.n796 585
R9523 GND.n9161 GND.n9160 585
R9524 GND.n9162 GND.n9161 585
R9525 GND.n795 GND.n794 585
R9526 GND.n9163 GND.n795 585
R9527 GND.n9166 GND.n9165 585
R9528 GND.n9165 GND.n9164 585
R9529 GND.n792 GND.n791 585
R9530 GND.n791 GND.n790 585
R9531 GND.n9171 GND.n9170 585
R9532 GND.n9172 GND.n9171 585
R9533 GND.n789 GND.n788 585
R9534 GND.n9173 GND.n789 585
R9535 GND.n9176 GND.n9175 585
R9536 GND.n9175 GND.n9174 585
R9537 GND.n786 GND.n785 585
R9538 GND.n785 GND.n784 585
R9539 GND.n9181 GND.n9180 585
R9540 GND.n9182 GND.n9181 585
R9541 GND.n783 GND.n782 585
R9542 GND.n9183 GND.n783 585
R9543 GND.n9186 GND.n9185 585
R9544 GND.n9185 GND.n9184 585
R9545 GND.n780 GND.n779 585
R9546 GND.n779 GND.n778 585
R9547 GND.n9191 GND.n9190 585
R9548 GND.n9192 GND.n9191 585
R9549 GND.n777 GND.n776 585
R9550 GND.n9193 GND.n777 585
R9551 GND.n9196 GND.n9195 585
R9552 GND.n9195 GND.n9194 585
R9553 GND.n774 GND.n773 585
R9554 GND.n773 GND.n772 585
R9555 GND.n9201 GND.n9200 585
R9556 GND.n9202 GND.n9201 585
R9557 GND.n771 GND.n770 585
R9558 GND.n9203 GND.n771 585
R9559 GND.n9206 GND.n9205 585
R9560 GND.n9205 GND.n9204 585
R9561 GND.n768 GND.n767 585
R9562 GND.n767 GND.n766 585
R9563 GND.n9211 GND.n9210 585
R9564 GND.n9212 GND.n9211 585
R9565 GND.n765 GND.n764 585
R9566 GND.n9213 GND.n765 585
R9567 GND.n9216 GND.n9215 585
R9568 GND.n9215 GND.n9214 585
R9569 GND.n762 GND.n761 585
R9570 GND.n761 GND.n760 585
R9571 GND.n9221 GND.n9220 585
R9572 GND.n9222 GND.n9221 585
R9573 GND.n759 GND.n758 585
R9574 GND.n9223 GND.n759 585
R9575 GND.n9226 GND.n9225 585
R9576 GND.n9225 GND.n9224 585
R9577 GND.n756 GND.n755 585
R9578 GND.n755 GND.n754 585
R9579 GND.n9231 GND.n9230 585
R9580 GND.n9232 GND.n9231 585
R9581 GND.n753 GND.n752 585
R9582 GND.n9233 GND.n753 585
R9583 GND.n9236 GND.n9235 585
R9584 GND.n9235 GND.n9234 585
R9585 GND.n750 GND.n749 585
R9586 GND.n749 GND.n748 585
R9587 GND.n9241 GND.n9240 585
R9588 GND.n9242 GND.n9241 585
R9589 GND.n747 GND.n746 585
R9590 GND.n9243 GND.n747 585
R9591 GND.n9246 GND.n9245 585
R9592 GND.n9245 GND.n9244 585
R9593 GND.n744 GND.n743 585
R9594 GND.n743 GND.n742 585
R9595 GND.n9251 GND.n9250 585
R9596 GND.n9252 GND.n9251 585
R9597 GND.n741 GND.n740 585
R9598 GND.n9253 GND.n741 585
R9599 GND.n9256 GND.n9255 585
R9600 GND.n9255 GND.n9254 585
R9601 GND.n738 GND.n737 585
R9602 GND.n737 GND.n736 585
R9603 GND.n9261 GND.n9260 585
R9604 GND.n9262 GND.n9261 585
R9605 GND.n735 GND.n734 585
R9606 GND.n9263 GND.n735 585
R9607 GND.n9266 GND.n9265 585
R9608 GND.n9265 GND.n9264 585
R9609 GND.n732 GND.n731 585
R9610 GND.n731 GND.n730 585
R9611 GND.n9271 GND.n9270 585
R9612 GND.n9272 GND.n9271 585
R9613 GND.n729 GND.n728 585
R9614 GND.n9273 GND.n729 585
R9615 GND.n9276 GND.n9275 585
R9616 GND.n9275 GND.n9274 585
R9617 GND.n726 GND.n725 585
R9618 GND.n725 GND.n724 585
R9619 GND.n9281 GND.n9280 585
R9620 GND.n9282 GND.n9281 585
R9621 GND.n723 GND.n722 585
R9622 GND.n9283 GND.n723 585
R9623 GND.n9286 GND.n9285 585
R9624 GND.n9285 GND.n9284 585
R9625 GND.n720 GND.n719 585
R9626 GND.n719 GND.n718 585
R9627 GND.n9291 GND.n9290 585
R9628 GND.n9292 GND.n9291 585
R9629 GND.n717 GND.n716 585
R9630 GND.n9293 GND.n717 585
R9631 GND.n9296 GND.n9295 585
R9632 GND.n9295 GND.n9294 585
R9633 GND.n714 GND.n713 585
R9634 GND.n713 GND.n712 585
R9635 GND.n9301 GND.n9300 585
R9636 GND.n9302 GND.n9301 585
R9637 GND.n711 GND.n710 585
R9638 GND.n9303 GND.n711 585
R9639 GND.n9306 GND.n9305 585
R9640 GND.n9305 GND.n9304 585
R9641 GND.n708 GND.n707 585
R9642 GND.n707 GND.n706 585
R9643 GND.n9311 GND.n9310 585
R9644 GND.n9312 GND.n9311 585
R9645 GND.n705 GND.n704 585
R9646 GND.n9313 GND.n705 585
R9647 GND.n9316 GND.n9315 585
R9648 GND.n9315 GND.n9314 585
R9649 GND.n702 GND.n701 585
R9650 GND.n701 GND.n700 585
R9651 GND.n9321 GND.n9320 585
R9652 GND.n9322 GND.n9321 585
R9653 GND.n9457 GND.n9456 585
R9654 GND.n9456 GND.n9455 585
R9655 GND.n621 GND.n620 585
R9656 GND.n9454 GND.n621 585
R9657 GND.n9452 GND.n9451 585
R9658 GND.n9453 GND.n9452 585
R9659 GND.n624 GND.n623 585
R9660 GND.n623 GND.n622 585
R9661 GND.n9446 GND.n9445 585
R9662 GND.n9445 GND.n9444 585
R9663 GND.n627 GND.n626 585
R9664 GND.n9443 GND.n627 585
R9665 GND.n9441 GND.n9440 585
R9666 GND.n9442 GND.n9441 585
R9667 GND.n630 GND.n629 585
R9668 GND.n629 GND.n628 585
R9669 GND.n9436 GND.n9435 585
R9670 GND.n9435 GND.n9434 585
R9671 GND.n633 GND.n632 585
R9672 GND.n9433 GND.n633 585
R9673 GND.n9431 GND.n9430 585
R9674 GND.n9432 GND.n9431 585
R9675 GND.n636 GND.n635 585
R9676 GND.n635 GND.n634 585
R9677 GND.n9426 GND.n9425 585
R9678 GND.n9425 GND.n9424 585
R9679 GND.n639 GND.n638 585
R9680 GND.n9423 GND.n639 585
R9681 GND.n9421 GND.n9420 585
R9682 GND.n9422 GND.n9421 585
R9683 GND.n642 GND.n641 585
R9684 GND.n641 GND.n640 585
R9685 GND.n9416 GND.n9415 585
R9686 GND.n9415 GND.n9414 585
R9687 GND.n645 GND.n644 585
R9688 GND.n9413 GND.n645 585
R9689 GND.n9411 GND.n9410 585
R9690 GND.n9412 GND.n9411 585
R9691 GND.n648 GND.n647 585
R9692 GND.n647 GND.n646 585
R9693 GND.n9406 GND.n9405 585
R9694 GND.n9405 GND.n9404 585
R9695 GND.n651 GND.n650 585
R9696 GND.n9403 GND.n651 585
R9697 GND.n9401 GND.n9400 585
R9698 GND.n9402 GND.n9401 585
R9699 GND.n654 GND.n653 585
R9700 GND.n653 GND.n652 585
R9701 GND.n9396 GND.n9395 585
R9702 GND.n9395 GND.n9394 585
R9703 GND.n657 GND.n656 585
R9704 GND.n9393 GND.n657 585
R9705 GND.n9391 GND.n9390 585
R9706 GND.n9392 GND.n9391 585
R9707 GND.n660 GND.n659 585
R9708 GND.n659 GND.n658 585
R9709 GND.n9386 GND.n9385 585
R9710 GND.n9385 GND.n9384 585
R9711 GND.n663 GND.n662 585
R9712 GND.n9383 GND.n663 585
R9713 GND.n9381 GND.n9380 585
R9714 GND.n9382 GND.n9381 585
R9715 GND.n666 GND.n665 585
R9716 GND.n665 GND.n664 585
R9717 GND.n9376 GND.n9375 585
R9718 GND.n9375 GND.n9374 585
R9719 GND.n669 GND.n668 585
R9720 GND.n9373 GND.n669 585
R9721 GND.n9371 GND.n9370 585
R9722 GND.n9372 GND.n9371 585
R9723 GND.n672 GND.n671 585
R9724 GND.n671 GND.n670 585
R9725 GND.n9366 GND.n9365 585
R9726 GND.n9365 GND.n9364 585
R9727 GND.n675 GND.n674 585
R9728 GND.n9363 GND.n675 585
R9729 GND.n9361 GND.n9360 585
R9730 GND.n9362 GND.n9361 585
R9731 GND.n678 GND.n677 585
R9732 GND.n677 GND.n676 585
R9733 GND.n9356 GND.n9355 585
R9734 GND.n9355 GND.n9354 585
R9735 GND.n681 GND.n680 585
R9736 GND.n9353 GND.n681 585
R9737 GND.n9351 GND.n9350 585
R9738 GND.n9352 GND.n9351 585
R9739 GND.n684 GND.n683 585
R9740 GND.n683 GND.n682 585
R9741 GND.n9346 GND.n9345 585
R9742 GND.n9345 GND.n9344 585
R9743 GND.n687 GND.n686 585
R9744 GND.n9343 GND.n687 585
R9745 GND.n9341 GND.n9340 585
R9746 GND.n9342 GND.n9341 585
R9747 GND.n690 GND.n689 585
R9748 GND.n689 GND.n688 585
R9749 GND.n9336 GND.n9335 585
R9750 GND.n9335 GND.n9334 585
R9751 GND.n693 GND.n692 585
R9752 GND.n9333 GND.n693 585
R9753 GND.n9331 GND.n9330 585
R9754 GND.n9332 GND.n9331 585
R9755 GND.n696 GND.n695 585
R9756 GND.n695 GND.n694 585
R9757 GND.n9326 GND.n9325 585
R9758 GND.n9325 GND.n9324 585
R9759 GND.n699 GND.n698 585
R9760 GND.n9323 GND.n699 585
R9761 GND.n6330 GND.n3231 585
R9762 GND.n7341 GND.n3231 585
R9763 GND.n6332 GND.n6331 585
R9764 GND.n6332 GND.n3978 585
R9765 GND.n6334 GND.n6333 585
R9766 GND.n6333 GND.n3985 585
R9767 GND.n6335 GND.n3991 585
R9768 GND.n6361 GND.n3991 585
R9769 GND.n6337 GND.n6336 585
R9770 GND.n6336 GND.n3989 585
R9771 GND.n6338 GND.n3999 585
R9772 GND.n6350 GND.n3999 585
R9773 GND.n6340 GND.n6339 585
R9774 GND.n6341 GND.n6340 585
R9775 GND.n4007 GND.n4006 585
R9776 GND.n4014 GND.n4006 585
R9777 GND.n6097 GND.n6096 585
R9778 GND.n6096 GND.n6095 585
R9779 GND.n4010 GND.n4009 585
R9780 GND.n4024 GND.n4010 585
R9781 GND.n5987 GND.n4021 585
R9782 GND.n6085 GND.n4021 585
R9783 GND.n5988 GND.n4030 585
R9784 GND.n6073 GND.n4030 585
R9785 GND.n5989 GND.n5981 585
R9786 GND.n5981 GND.n4037 585
R9787 GND.n5991 GND.n5990 585
R9788 GND.n5991 GND.n4036 585
R9789 GND.n5992 GND.n5980 585
R9790 GND.n5992 GND.n4041 585
R9791 GND.n5994 GND.n5993 585
R9792 GND.n5993 GND.n4047 585
R9793 GND.n5995 GND.n4054 585
R9794 GND.n6028 GND.n4054 585
R9795 GND.n5997 GND.n5996 585
R9796 GND.n5996 GND.n4052 585
R9797 GND.n5998 GND.n4062 585
R9798 GND.n6009 GND.n4062 585
R9799 GND.n6000 GND.n5999 585
R9800 GND.n6001 GND.n6000 585
R9801 GND.n4071 GND.n4070 585
R9802 GND.n4079 GND.n4070 585
R9803 GND.n5972 GND.n5971 585
R9804 GND.n5971 GND.n5970 585
R9805 GND.n4074 GND.n4073 585
R9806 GND.n4088 GND.n4074 585
R9807 GND.n5761 GND.n4086 585
R9808 GND.n5960 GND.n4086 585
R9809 GND.n5763 GND.n5762 585
R9810 GND.n5763 GND.n4093 585
R9811 GND.n5765 GND.n5764 585
R9812 GND.n5764 GND.n4100 585
R9813 GND.n5766 GND.n4106 585
R9814 GND.n5917 GND.n4106 585
R9815 GND.n5768 GND.n5767 585
R9816 GND.n5767 GND.n4104 585
R9817 GND.n5769 GND.n4116 585
R9818 GND.n5907 GND.n4116 585
R9819 GND.n5770 GND.n5751 585
R9820 GND.n5751 GND.n4124 585
R9821 GND.n5772 GND.n5771 585
R9822 GND.n5772 GND.n4122 585
R9823 GND.n5773 GND.n5750 585
R9824 GND.n5773 GND.n4129 585
R9825 GND.n5775 GND.n5774 585
R9826 GND.n5774 GND.n4135 585
R9827 GND.n5776 GND.n4141 585
R9828 GND.n5877 GND.n4141 585
R9829 GND.n5778 GND.n5777 585
R9830 GND.n5777 GND.n4139 585
R9831 GND.n5779 GND.n4149 585
R9832 GND.n5861 GND.n4149 585
R9833 GND.n5780 GND.n4157 585
R9834 GND.n5853 GND.n4157 585
R9835 GND.n5781 GND.n5741 585
R9836 GND.n5741 GND.n4162 585
R9837 GND.n5783 GND.n5782 585
R9838 GND.n5783 GND.n4160 585
R9839 GND.n5784 GND.n5740 585
R9840 GND.n5784 GND.n4166 585
R9841 GND.n5786 GND.n5785 585
R9842 GND.n5785 GND.n4172 585
R9843 GND.n5787 GND.n4178 585
R9844 GND.n5820 GND.n4178 585
R9845 GND.n5789 GND.n5788 585
R9846 GND.n5788 GND.n4176 585
R9847 GND.n5790 GND.n4187 585
R9848 GND.n5801 GND.n4187 585
R9849 GND.n5792 GND.n5791 585
R9850 GND.n5793 GND.n5792 585
R9851 GND.n4197 GND.n4196 585
R9852 GND.n4196 GND.n4194 585
R9853 GND.n5732 GND.n5731 585
R9854 GND.n5731 GND.n5730 585
R9855 GND.n4200 GND.n4199 585
R9856 GND.n4212 GND.n4200 585
R9857 GND.n5703 GND.n4210 585
R9858 GND.n5720 GND.n4210 585
R9859 GND.n5705 GND.n5704 585
R9860 GND.n5707 GND.n5705 585
R9861 GND.n4221 GND.n4220 585
R9862 GND.n5676 GND.n4220 585
R9863 GND.n5698 GND.n5697 585
R9864 GND.n5697 GND.n5696 585
R9865 GND.n4224 GND.n4223 585
R9866 GND.n4235 GND.n4224 585
R9867 GND.n5510 GND.n4233 585
R9868 GND.n5686 GND.n4233 585
R9869 GND.n5512 GND.n5511 585
R9870 GND.n5511 GND.n4244 585
R9871 GND.n5513 GND.n4249 585
R9872 GND.n5638 GND.n4249 585
R9873 GND.n5515 GND.n5514 585
R9874 GND.n5514 GND.n4259 585
R9875 GND.n5516 GND.n4257 585
R9876 GND.n5630 GND.n4257 585
R9877 GND.n5518 GND.n5517 585
R9878 GND.n5518 GND.n4263 585
R9879 GND.n5520 GND.n5519 585
R9880 GND.n5519 GND.n4270 585
R9881 GND.n5521 GND.n4277 585
R9882 GND.n5602 GND.n4277 585
R9883 GND.n5523 GND.n5522 585
R9884 GND.n5522 GND.n4275 585
R9885 GND.n5524 GND.n4286 585
R9886 GND.n5592 GND.n4286 585
R9887 GND.n5525 GND.n5496 585
R9888 GND.n5496 GND.n5495 585
R9889 GND.n5527 GND.n5526 585
R9890 GND.n5527 GND.n4292 585
R9891 GND.n5528 GND.n5494 585
R9892 GND.n5528 GND.n4298 585
R9893 GND.n5530 GND.n5529 585
R9894 GND.n5529 GND.n4304 585
R9895 GND.n5531 GND.n4310 585
R9896 GND.n5562 GND.n4310 585
R9897 GND.n5533 GND.n5532 585
R9898 GND.n5532 GND.n4308 585
R9899 GND.n5534 GND.n4318 585
R9900 GND.n5546 GND.n4318 585
R9901 GND.n5536 GND.n5535 585
R9902 GND.n5537 GND.n5536 585
R9903 GND.n4327 GND.n4326 585
R9904 GND.n4334 GND.n4326 585
R9905 GND.n5486 GND.n5485 585
R9906 GND.n5485 GND.n5484 585
R9907 GND.n4330 GND.n4329 585
R9908 GND.n4344 GND.n4330 585
R9909 GND.n5345 GND.n4341 585
R9910 GND.n5474 GND.n4341 585
R9911 GND.n5347 GND.n5346 585
R9912 GND.n5347 GND.n4349 585
R9913 GND.n5349 GND.n5348 585
R9914 GND.n5348 GND.n4356 585
R9915 GND.n5350 GND.n4361 585
R9916 GND.n5431 GND.n4361 585
R9917 GND.n5353 GND.n5352 585
R9918 GND.n5352 GND.n5351 585
R9919 GND.n5354 GND.n4371 585
R9920 GND.n5421 GND.n4371 585
R9921 GND.n5355 GND.n5335 585
R9922 GND.n5335 GND.n4379 585
R9923 GND.n5357 GND.n5356 585
R9924 GND.n5357 GND.n4378 585
R9925 GND.n5358 GND.n5334 585
R9926 GND.n5358 GND.n4384 585
R9927 GND.n5360 GND.n5359 585
R9928 GND.n5359 GND.n4390 585
R9929 GND.n5361 GND.n4397 585
R9930 GND.n5391 GND.n4397 585
R9931 GND.n5363 GND.n5362 585
R9932 GND.n5362 GND.n4395 585
R9933 GND.n5364 GND.n4405 585
R9934 GND.n5375 GND.n4405 585
R9935 GND.n5366 GND.n5365 585
R9936 GND.n5367 GND.n5366 585
R9937 GND.n4413 GND.n4412 585
R9938 GND.n4421 GND.n4412 585
R9939 GND.n5326 GND.n5325 585
R9940 GND.n5325 GND.n5324 585
R9941 GND.n4416 GND.n4415 585
R9942 GND.n5294 GND.n4416 585
R9943 GND.n5184 GND.n4428 585
R9944 GND.n5314 GND.n4428 585
R9945 GND.n5186 GND.n5185 585
R9946 GND.n5186 GND.n4434 585
R9947 GND.n5188 GND.n5187 585
R9948 GND.n5187 GND.n4442 585
R9949 GND.n5189 GND.n4448 585
R9950 GND.n5269 GND.n4448 585
R9951 GND.n5191 GND.n5190 585
R9952 GND.n5190 GND.n4446 585
R9953 GND.n5192 GND.n4457 585
R9954 GND.n5259 GND.n4457 585
R9955 GND.n5193 GND.n5174 585
R9956 GND.n5174 GND.n4465 585
R9957 GND.n5195 GND.n5194 585
R9958 GND.n5195 GND.n4463 585
R9959 GND.n5196 GND.n5173 585
R9960 GND.n5196 GND.n4470 585
R9961 GND.n5198 GND.n5197 585
R9962 GND.n5197 GND.n4476 585
R9963 GND.n5199 GND.n4482 585
R9964 GND.n5229 GND.n4482 585
R9965 GND.n5201 GND.n5200 585
R9966 GND.n5200 GND.n4480 585
R9967 GND.n5202 GND.n4491 585
R9968 GND.n5213 GND.n4491 585
R9969 GND.n5204 GND.n5203 585
R9970 GND.n5205 GND.n5204 585
R9971 GND.n4499 GND.n4498 585
R9972 GND.n5144 GND.n4498 585
R9973 GND.n5165 GND.n5164 585
R9974 GND.n5164 GND.n5163 585
R9975 GND.n4502 GND.n4501 585
R9976 GND.n4513 GND.n4502 585
R9977 GND.n5021 GND.n4511 585
R9978 GND.n5153 GND.n4511 585
R9979 GND.n5023 GND.n5022 585
R9980 GND.n5022 GND.n4523 585
R9981 GND.n5024 GND.n4529 585
R9982 GND.n5116 GND.n4529 585
R9983 GND.n5026 GND.n5025 585
R9984 GND.n5025 GND.n4539 585
R9985 GND.n5027 GND.n4537 585
R9986 GND.n5108 GND.n4537 585
R9987 GND.n5028 GND.n4544 585
R9988 GND.n5101 GND.n4544 585
R9989 GND.n5029 GND.n5011 585
R9990 GND.n5011 GND.n4551 585
R9991 GND.n5031 GND.n5030 585
R9992 GND.n5031 GND.n4550 585
R9993 GND.n5032 GND.n5010 585
R9994 GND.n5032 GND.n4555 585
R9995 GND.n5034 GND.n5033 585
R9996 GND.n5033 GND.n4562 585
R9997 GND.n5035 GND.n4568 585
R9998 GND.n5069 GND.n4568 585
R9999 GND.n5037 GND.n5036 585
R10000 GND.n5036 GND.n4566 585
R10001 GND.n5038 GND.n4576 585
R10002 GND.n5050 GND.n4576 585
R10003 GND.n5040 GND.n5039 585
R10004 GND.n5042 GND.n5040 585
R10005 GND.n4585 GND.n4584 585
R10006 GND.n4592 GND.n4584 585
R10007 GND.n5002 GND.n5001 585
R10008 GND.n5001 GND.n5000 585
R10009 GND.n4588 GND.n4587 585
R10010 GND.n4601 GND.n4588 585
R10011 GND.n4873 GND.n4599 585
R10012 GND.n4990 GND.n4599 585
R10013 GND.n4875 GND.n4874 585
R10014 GND.n4875 GND.n4606 585
R10015 GND.n4877 GND.n4876 585
R10016 GND.n4876 GND.n4612 585
R10017 GND.n4878 GND.n4619 585
R10018 GND.n4946 GND.n4619 585
R10019 GND.n4880 GND.n4879 585
R10020 GND.n4879 GND.n4617 585
R10021 GND.n4881 GND.n4629 585
R10022 GND.n4936 GND.n4629 585
R10023 GND.n4883 GND.n4882 585
R10024 GND.n4883 GND.n4636 585
R10025 GND.n4884 GND.n4864 585
R10026 GND.n4884 GND.n4635 585
R10027 GND.n4886 GND.n4885 585
R10028 GND.n4885 GND.n4642 585
R10029 GND.n4887 GND.n4655 585
R10030 GND.n4655 GND.n4648 585
R10031 GND.n4889 GND.n4888 585
R10032 GND.n4906 GND.n4889 585
R10033 GND.n4656 GND.n4654 585
R10034 GND.n4654 GND.n4652 585
R10035 GND.n4858 GND.n4857 585
R10036 GND.n4857 GND.n4856 585
R10037 GND.n4658 GND.n3022 585
R10038 GND.n7553 GND.n3022 585
R10039 GND.n4668 GND.n4667 585
R10040 GND.n4669 GND.n4668 585
R10041 GND.n4662 GND.n3011 585
R10042 GND.n7559 GND.n3011 585
R10043 GND.n4663 GND.n1837 585
R10044 GND.n3001 GND.n1837 585
R10045 GND.n7869 GND.n7868 585
R10046 GND.n1838 GND.n1836 585
R10047 GND.n7865 GND.n7864 585
R10048 GND.n7866 GND.n7865 585
R10049 GND.n1851 GND.n1850 585
R10050 GND.n7857 GND.n1862 585
R10051 GND.n7856 GND.n1863 585
R10052 GND.n1870 GND.n1864 585
R10053 GND.n7849 GND.n1871 585
R10054 GND.n7848 GND.n1872 585
R10055 GND.n1874 GND.n1873 585
R10056 GND.n7841 GND.n1884 585
R10057 GND.n7840 GND.n1885 585
R10058 GND.n3033 GND.n1886 585
R10059 GND.n3035 GND.n3034 585
R10060 GND.n3037 GND.n3036 585
R10061 GND.n3042 GND.n3038 585
R10062 GND.n3030 GND.n3029 585
R10063 GND.n3046 GND.n3031 585
R10064 GND.n3048 GND.n3047 585
R10065 GND.n3049 GND.n1848 585
R10066 GND.n7866 GND.n1848 585
R10067 GND.n6418 GND.n3229 585
R10068 GND.n6420 GND.n6417 585
R10069 GND.n6421 GND.n3972 585
R10070 GND.n6422 GND.n3971 585
R10071 GND.n6425 GND.n3966 585
R10072 GND.n6426 GND.n3965 585
R10073 GND.n6427 GND.n3964 585
R10074 GND.n6411 GND.n3352 585
R10075 GND.n7262 GND.n3351 585
R10076 GND.n7263 GND.n3350 585
R10077 GND.n6408 GND.n3340 585
R10078 GND.n7270 GND.n3339 585
R10079 GND.n7271 GND.n3338 585
R10080 GND.n6406 GND.n3332 585
R10081 GND.n7278 GND.n3331 585
R10082 GND.n7279 GND.n3330 585
R10083 GND.n6403 GND.n3322 585
R10084 GND.n7286 GND.n3321 585
R10085 GND.n7287 GND.n3320 585
R10086 GND.n6401 GND.n3319 585
R10087 GND.n7343 GND.n7342 585
R10088 GND.n7342 GND.n7341 585
R10089 GND.n3228 GND.n3226 585
R10090 GND.n3978 GND.n3228 585
R10091 GND.n7347 GND.n3225 585
R10092 GND.n3985 GND.n3225 585
R10093 GND.n7348 GND.n3224 585
R10094 GND.n6361 GND.n3224 585
R10095 GND.n7349 GND.n3223 585
R10096 GND.n3989 GND.n3223 585
R10097 GND.n6349 GND.n3221 585
R10098 GND.n6350 GND.n6349 585
R10099 GND.n7353 GND.n3220 585
R10100 GND.n6341 GND.n3220 585
R10101 GND.n7354 GND.n3219 585
R10102 GND.n4014 GND.n3219 585
R10103 GND.n7355 GND.n3218 585
R10104 GND.n6095 GND.n3218 585
R10105 GND.n4023 GND.n3216 585
R10106 GND.n4024 GND.n4023 585
R10107 GND.n7359 GND.n3215 585
R10108 GND.n6085 GND.n3215 585
R10109 GND.n7360 GND.n3214 585
R10110 GND.n6073 GND.n3214 585
R10111 GND.n7361 GND.n3213 585
R10112 GND.n4037 GND.n3213 585
R10113 GND.n4035 GND.n3211 585
R10114 GND.n4036 GND.n4035 585
R10115 GND.n7365 GND.n3210 585
R10116 GND.n4041 GND.n3210 585
R10117 GND.n7366 GND.n3209 585
R10118 GND.n4047 GND.n3209 585
R10119 GND.n7367 GND.n3208 585
R10120 GND.n6028 GND.n3208 585
R10121 GND.n4051 GND.n3206 585
R10122 GND.n4052 GND.n4051 585
R10123 GND.n7371 GND.n3205 585
R10124 GND.n6009 GND.n3205 585
R10125 GND.n7372 GND.n3204 585
R10126 GND.n6001 GND.n3204 585
R10127 GND.n7373 GND.n3203 585
R10128 GND.n4079 GND.n3203 585
R10129 GND.n4077 GND.n3201 585
R10130 GND.n5970 GND.n4077 585
R10131 GND.n7377 GND.n3200 585
R10132 GND.n4088 GND.n3200 585
R10133 GND.n7378 GND.n3199 585
R10134 GND.n5960 GND.n3199 585
R10135 GND.n7379 GND.n3198 585
R10136 GND.n4093 GND.n3198 585
R10137 GND.n4099 GND.n3196 585
R10138 GND.n4100 GND.n4099 585
R10139 GND.n7383 GND.n3195 585
R10140 GND.n5917 GND.n3195 585
R10141 GND.n7384 GND.n3194 585
R10142 GND.n4104 GND.n3194 585
R10143 GND.n7385 GND.n3193 585
R10144 GND.n5907 GND.n3193 585
R10145 GND.n4123 GND.n3191 585
R10146 GND.n4124 GND.n4123 585
R10147 GND.n7389 GND.n3190 585
R10148 GND.n4122 GND.n3190 585
R10149 GND.n7390 GND.n3189 585
R10150 GND.n4129 GND.n3189 585
R10151 GND.n7391 GND.n3188 585
R10152 GND.n4135 GND.n3188 585
R10153 GND.n4142 GND.n3186 585
R10154 GND.n5877 GND.n4142 585
R10155 GND.n7395 GND.n3185 585
R10156 GND.n4139 GND.n3185 585
R10157 GND.n7396 GND.n3184 585
R10158 GND.n5861 GND.n3184 585
R10159 GND.n7397 GND.n3183 585
R10160 GND.n5853 GND.n3183 585
R10161 GND.n4161 GND.n3181 585
R10162 GND.n4162 GND.n4161 585
R10163 GND.n7401 GND.n3180 585
R10164 GND.n4160 GND.n3180 585
R10165 GND.n7402 GND.n3179 585
R10166 GND.n4166 GND.n3179 585
R10167 GND.n7403 GND.n3178 585
R10168 GND.n4172 GND.n3178 585
R10169 GND.n4179 GND.n3176 585
R10170 GND.n5820 GND.n4179 585
R10171 GND.n7407 GND.n3175 585
R10172 GND.n4176 GND.n3175 585
R10173 GND.n7408 GND.n3174 585
R10174 GND.n5801 GND.n3174 585
R10175 GND.n7409 GND.n3173 585
R10176 GND.n5793 GND.n3173 585
R10177 GND.n4193 GND.n3171 585
R10178 GND.n4194 GND.n4193 585
R10179 GND.n7413 GND.n3170 585
R10180 GND.n5730 GND.n3170 585
R10181 GND.n7414 GND.n3169 585
R10182 GND.n4212 GND.n3169 585
R10183 GND.n7415 GND.n3168 585
R10184 GND.n5720 GND.n3168 585
R10185 GND.n5706 GND.n3166 585
R10186 GND.n5707 GND.n5706 585
R10187 GND.n7419 GND.n3165 585
R10188 GND.n5676 GND.n3165 585
R10189 GND.n7420 GND.n3164 585
R10190 GND.n5696 GND.n3164 585
R10191 GND.n7421 GND.n3163 585
R10192 GND.n4235 GND.n3163 585
R10193 GND.n5685 GND.n3161 585
R10194 GND.n5686 GND.n5685 585
R10195 GND.n7425 GND.n3160 585
R10196 GND.n4244 GND.n3160 585
R10197 GND.n7426 GND.n3159 585
R10198 GND.n5638 GND.n3159 585
R10199 GND.n7427 GND.n3158 585
R10200 GND.n4259 GND.n3158 585
R10201 GND.n5629 GND.n3156 585
R10202 GND.n5630 GND.n5629 585
R10203 GND.n7431 GND.n3155 585
R10204 GND.n4263 GND.n3155 585
R10205 GND.n7432 GND.n3154 585
R10206 GND.n4270 GND.n3154 585
R10207 GND.n7433 GND.n3153 585
R10208 GND.n5602 GND.n3153 585
R10209 GND.n4274 GND.n3151 585
R10210 GND.n4275 GND.n4274 585
R10211 GND.n7437 GND.n3150 585
R10212 GND.n5592 GND.n3150 585
R10213 GND.n7438 GND.n3149 585
R10214 GND.n5495 GND.n3149 585
R10215 GND.n7439 GND.n3148 585
R10216 GND.n4292 GND.n3148 585
R10217 GND.n4297 GND.n3146 585
R10218 GND.n4298 GND.n4297 585
R10219 GND.n7443 GND.n3145 585
R10220 GND.n4304 GND.n3145 585
R10221 GND.n7444 GND.n3144 585
R10222 GND.n5562 GND.n3144 585
R10223 GND.n7445 GND.n3143 585
R10224 GND.n4308 GND.n3143 585
R10225 GND.n5545 GND.n3141 585
R10226 GND.n5546 GND.n5545 585
R10227 GND.n7449 GND.n3140 585
R10228 GND.n5537 GND.n3140 585
R10229 GND.n7450 GND.n3139 585
R10230 GND.n4334 GND.n3139 585
R10231 GND.n7451 GND.n3138 585
R10232 GND.n5484 GND.n3138 585
R10233 GND.n4343 GND.n3136 585
R10234 GND.n4344 GND.n4343 585
R10235 GND.n7455 GND.n3135 585
R10236 GND.n5474 GND.n3135 585
R10237 GND.n7456 GND.n3134 585
R10238 GND.n4349 GND.n3134 585
R10239 GND.n7457 GND.n3133 585
R10240 GND.n4356 GND.n3133 585
R10241 GND.n4362 GND.n3131 585
R10242 GND.n5431 GND.n4362 585
R10243 GND.n7461 GND.n3130 585
R10244 GND.n5351 GND.n3130 585
R10245 GND.n7462 GND.n3129 585
R10246 GND.n5421 GND.n3129 585
R10247 GND.n7463 GND.n3128 585
R10248 GND.n4379 GND.n3128 585
R10249 GND.n4377 GND.n3126 585
R10250 GND.n4378 GND.n4377 585
R10251 GND.n7467 GND.n3125 585
R10252 GND.n4384 GND.n3125 585
R10253 GND.n7468 GND.n3124 585
R10254 GND.n4390 GND.n3124 585
R10255 GND.n7469 GND.n3123 585
R10256 GND.n5391 GND.n3123 585
R10257 GND.n4394 GND.n3121 585
R10258 GND.n4395 GND.n4394 585
R10259 GND.n7473 GND.n3120 585
R10260 GND.n5375 GND.n3120 585
R10261 GND.n7474 GND.n3119 585
R10262 GND.n5367 GND.n3119 585
R10263 GND.n7475 GND.n3118 585
R10264 GND.n4421 GND.n3118 585
R10265 GND.n4419 GND.n3116 585
R10266 GND.n5324 GND.n4419 585
R10267 GND.n7479 GND.n3115 585
R10268 GND.n5294 GND.n3115 585
R10269 GND.n7480 GND.n3114 585
R10270 GND.n5314 GND.n3114 585
R10271 GND.n7481 GND.n3113 585
R10272 GND.n4434 GND.n3113 585
R10273 GND.n4441 GND.n3111 585
R10274 GND.n4442 GND.n4441 585
R10275 GND.n7485 GND.n3110 585
R10276 GND.n5269 GND.n3110 585
R10277 GND.n7486 GND.n3109 585
R10278 GND.n4446 GND.n3109 585
R10279 GND.n7487 GND.n3108 585
R10280 GND.n5259 GND.n3108 585
R10281 GND.n4464 GND.n3106 585
R10282 GND.n4465 GND.n4464 585
R10283 GND.n7491 GND.n3105 585
R10284 GND.n4463 GND.n3105 585
R10285 GND.n7492 GND.n3104 585
R10286 GND.n4470 GND.n3104 585
R10287 GND.n7493 GND.n3103 585
R10288 GND.n4476 GND.n3103 585
R10289 GND.n4483 GND.n3101 585
R10290 GND.n5229 GND.n4483 585
R10291 GND.n7497 GND.n3100 585
R10292 GND.n4480 GND.n3100 585
R10293 GND.n7498 GND.n3099 585
R10294 GND.n5213 GND.n3099 585
R10295 GND.n7499 GND.n3098 585
R10296 GND.n5205 GND.n3098 585
R10297 GND.n5143 GND.n3096 585
R10298 GND.n5144 GND.n5143 585
R10299 GND.n7503 GND.n3095 585
R10300 GND.n5163 GND.n3095 585
R10301 GND.n7504 GND.n3094 585
R10302 GND.n4513 GND.n3094 585
R10303 GND.n7505 GND.n3093 585
R10304 GND.n5153 GND.n3093 585
R10305 GND.n4522 GND.n3091 585
R10306 GND.n4523 GND.n4522 585
R10307 GND.n7509 GND.n3090 585
R10308 GND.n5116 GND.n3090 585
R10309 GND.n7510 GND.n3089 585
R10310 GND.n4539 GND.n3089 585
R10311 GND.n7511 GND.n3088 585
R10312 GND.n5108 GND.n3088 585
R10313 GND.n4545 GND.n3086 585
R10314 GND.n5101 GND.n4545 585
R10315 GND.n7515 GND.n3085 585
R10316 GND.n4551 GND.n3085 585
R10317 GND.n7516 GND.n3084 585
R10318 GND.n4550 GND.n3084 585
R10319 GND.n7517 GND.n3083 585
R10320 GND.n4555 GND.n3083 585
R10321 GND.n4561 GND.n3081 585
R10322 GND.n4562 GND.n4561 585
R10323 GND.n7521 GND.n3080 585
R10324 GND.n5069 GND.n3080 585
R10325 GND.n7522 GND.n3079 585
R10326 GND.n4566 GND.n3079 585
R10327 GND.n7523 GND.n3078 585
R10328 GND.n5050 GND.n3078 585
R10329 GND.n5041 GND.n3076 585
R10330 GND.n5042 GND.n5041 585
R10331 GND.n7527 GND.n3075 585
R10332 GND.n4592 GND.n3075 585
R10333 GND.n7528 GND.n3074 585
R10334 GND.n5000 GND.n3074 585
R10335 GND.n7529 GND.n3073 585
R10336 GND.n4601 GND.n3073 585
R10337 GND.n4989 GND.n3071 585
R10338 GND.n4990 GND.n4989 585
R10339 GND.n7533 GND.n3070 585
R10340 GND.n4606 GND.n3070 585
R10341 GND.n7534 GND.n3069 585
R10342 GND.n4612 GND.n3069 585
R10343 GND.n7535 GND.n3068 585
R10344 GND.n4946 GND.n3068 585
R10345 GND.n4616 GND.n3066 585
R10346 GND.n4617 GND.n4616 585
R10347 GND.n7539 GND.n3065 585
R10348 GND.n4936 GND.n3065 585
R10349 GND.n7540 GND.n3064 585
R10350 GND.n4636 GND.n3064 585
R10351 GND.n7541 GND.n3063 585
R10352 GND.n4635 GND.n3063 585
R10353 GND.n4641 GND.n3061 585
R10354 GND.n4642 GND.n4641 585
R10355 GND.n7545 GND.n3060 585
R10356 GND.n4648 GND.n3060 585
R10357 GND.n7546 GND.n3059 585
R10358 GND.n4906 GND.n3059 585
R10359 GND.n7547 GND.n3058 585
R10360 GND.n4652 GND.n3058 585
R10361 GND.n3027 GND.n3025 585
R10362 GND.n4856 GND.n3025 585
R10363 GND.n7552 GND.n7551 585
R10364 GND.n7553 GND.n7552 585
R10365 GND.n3026 GND.n3024 585
R10366 GND.n4669 GND.n3024 585
R10367 GND.n3054 GND.n3013 585
R10368 GND.n7559 GND.n3013 585
R10369 GND.n3053 GND.n3052 585
R10370 GND.n3052 GND.n3001 585
R10371 GND.n1774 GND.n1767 585
R10372 GND.n7924 GND.n1774 585
R10373 GND.n7828 GND.n1766 585
R10374 GND.n7829 GND.n7828 585
R10375 GND.n7827 GND.n1765 585
R10376 GND.n7827 GND.n7826 585
R10377 GND.n1893 GND.n1892 585
R10378 GND.n7807 GND.n1893 585
R10379 GND.n7817 GND.n1759 585
R10380 GND.n7818 GND.n7817 585
R10381 GND.n7816 GND.n1758 585
R10382 GND.n7816 GND.n7815 585
R10383 GND.n1903 GND.n1757 585
R10384 GND.n1916 GND.n1903 585
R10385 GND.n1914 GND.n1913 585
R10386 GND.n7801 GND.n1914 585
R10387 GND.n7789 GND.n1751 585
R10388 GND.n7789 GND.n7788 585
R10389 GND.n7790 GND.n1750 585
R10390 GND.n7791 GND.n7790 585
R10391 GND.n7787 GND.n1749 585
R10392 GND.n7787 GND.n7786 585
R10393 GND.n1927 GND.n1926 585
R10394 GND.n1939 GND.n1927 585
R10395 GND.n1937 GND.n1743 585
R10396 GND.n7777 GND.n1937 585
R10397 GND.n7765 GND.n1742 585
R10398 GND.n7765 GND.n7764 585
R10399 GND.n7766 GND.n1741 585
R10400 GND.n7767 GND.n7766 585
R10401 GND.n7762 GND.n1949 585
R10402 GND.n7762 GND.n7761 585
R10403 GND.n1948 GND.n1735 585
R10404 GND.n1962 GND.n1948 585
R10405 GND.n1960 GND.n1734 585
R10406 GND.n7752 GND.n1960 585
R10407 GND.n7739 GND.n1733 585
R10408 GND.n7739 GND.n7738 585
R10409 GND.n7741 GND.n7740 585
R10410 GND.n7742 GND.n7741 585
R10411 GND.n7737 GND.n1727 585
R10412 GND.n7737 GND.n7736 585
R10413 GND.n1971 GND.n1726 585
R10414 GND.n1984 GND.n1971 585
R10415 GND.n1981 GND.n1725 585
R10416 GND.n7727 GND.n1981 585
R10417 GND.n7715 GND.n7713 585
R10418 GND.n7715 GND.n7714 585
R10419 GND.n7716 GND.n1719 585
R10420 GND.n7717 GND.n7716 585
R10421 GND.n7712 GND.n1718 585
R10422 GND.n7712 GND.n7711 585
R10423 GND.n1993 GND.n1717 585
R10424 GND.n2007 GND.n1993 585
R10425 GND.n2005 GND.n2004 585
R10426 GND.n7702 GND.n2005 585
R10427 GND.n7690 GND.n1711 585
R10428 GND.n7690 GND.n7689 585
R10429 GND.n7691 GND.n1710 585
R10430 GND.n7692 GND.n7691 585
R10431 GND.n7688 GND.n1709 585
R10432 GND.n7688 GND.n7687 585
R10433 GND.n2018 GND.n2017 585
R10434 GND.n2030 GND.n2018 585
R10435 GND.n2028 GND.n1703 585
R10436 GND.n7678 GND.n2028 585
R10437 GND.n7666 GND.n1702 585
R10438 GND.n7666 GND.n7665 585
R10439 GND.n7667 GND.n1701 585
R10440 GND.n7668 GND.n7667 585
R10441 GND.n2039 GND.n2038 585
R10442 GND.n2889 GND.n2039 585
R10443 GND.n2056 GND.n1695 585
R10444 GND.n2056 GND.n2046 585
R10445 GND.n2057 GND.n1694 585
R10446 GND.n2880 GND.n2057 585
R10447 GND.n2867 GND.n1693 585
R10448 GND.n2867 GND.n2866 585
R10449 GND.n2869 GND.n2868 585
R10450 GND.n2870 GND.n2869 585
R10451 GND.n2865 GND.n1687 585
R10452 GND.n2865 GND.n2864 585
R10453 GND.n2067 GND.n1686 585
R10454 GND.n2080 GND.n2067 585
R10455 GND.n2077 GND.n1685 585
R10456 GND.n2855 GND.n2077 585
R10457 GND.n2843 GND.n2841 585
R10458 GND.n2843 GND.n2842 585
R10459 GND.n2844 GND.n1679 585
R10460 GND.n2845 GND.n2844 585
R10461 GND.n2840 GND.n1678 585
R10462 GND.n2840 GND.n2839 585
R10463 GND.n2089 GND.n1677 585
R10464 GND.n2103 GND.n2089 585
R10465 GND.n2101 GND.n2100 585
R10466 GND.n2830 GND.n2101 585
R10467 GND.n2790 GND.n1671 585
R10468 GND.n2791 GND.n2790 585
R10469 GND.n2789 GND.n1670 585
R10470 GND.n2789 GND.n2788 585
R10471 GND.n2143 GND.n1669 585
R10472 GND.n2146 GND.n2143 585
R10473 GND.n2801 GND.n2144 585
R10474 GND.n2801 GND.n2800 585
R10475 GND.n2802 GND.n1663 585
R10476 GND.n2803 GND.n2802 585
R10477 GND.n2136 GND.n1662 585
R10478 GND.n2808 GND.n2136 585
R10479 GND.n2135 GND.n1661 585
R10480 GND.n2135 GND.n2131 585
R10481 GND.n2122 GND.n2121 585
R10482 GND.n2124 GND.n2122 585
R10483 GND.n2818 GND.n1655 585
R10484 GND.n2818 GND.n2817 585
R10485 GND.n2819 GND.n1654 585
R10486 GND.n2820 GND.n2819 585
R10487 GND.n2120 GND.n1653 585
R10488 GND.n2666 GND.n2120 585
R10489 GND.n2198 GND.n2197 585
R10490 GND.n2760 GND.n2198 585
R10491 GND.n2750 GND.n1647 585
R10492 GND.n2750 GND.n2749 585
R10493 GND.n2751 GND.n1646 585
R10494 GND.n2752 GND.n2751 585
R10495 GND.n2748 GND.n1645 585
R10496 GND.n2748 GND.n2747 585
R10497 GND.n2209 GND.n2208 585
R10498 GND.n2221 GND.n2209 585
R10499 GND.n2219 GND.n1639 585
R10500 GND.n2738 GND.n2219 585
R10501 GND.n2726 GND.n1638 585
R10502 GND.n2726 GND.n2725 585
R10503 GND.n2727 GND.n1637 585
R10504 GND.n2728 GND.n2727 585
R10505 GND.n2723 GND.n2231 585
R10506 GND.n2723 GND.n2722 585
R10507 GND.n2230 GND.n1631 585
R10508 GND.n2244 GND.n2230 585
R10509 GND.n2242 GND.n1630 585
R10510 GND.n2713 GND.n2242 585
R10511 GND.n2700 GND.n1629 585
R10512 GND.n2700 GND.n2699 585
R10513 GND.n2702 GND.n2701 585
R10514 GND.n2703 GND.n2702 585
R10515 GND.n2698 GND.n1623 585
R10516 GND.n2698 GND.n2697 585
R10517 GND.n2252 GND.n1622 585
R10518 GND.n2644 GND.n2252 585
R10519 GND.n2633 GND.n1621 585
R10520 GND.n2633 GND.n2261 585
R10521 GND.n2635 GND.n2634 585
R10522 GND.n2636 GND.n2635 585
R10523 GND.n2632 GND.n1615 585
R10524 GND.n2632 GND.n2631 585
R10525 GND.n2272 GND.n1614 585
R10526 GND.n2285 GND.n2272 585
R10527 GND.n2282 GND.n1613 585
R10528 GND.n2613 GND.n2282 585
R10529 GND.n2601 GND.n2599 585
R10530 GND.n2601 GND.n2600 585
R10531 GND.n2602 GND.n1607 585
R10532 GND.n2603 GND.n2602 585
R10533 GND.n2598 GND.n1606 585
R10534 GND.n2598 GND.n2597 585
R10535 GND.n2294 GND.n1605 585
R10536 GND.n2308 GND.n2294 585
R10537 GND.n2306 GND.n2305 585
R10538 GND.n2588 GND.n2306 585
R10539 GND.n2576 GND.n1599 585
R10540 GND.n2576 GND.n2575 585
R10541 GND.n2577 GND.n1598 585
R10542 GND.n2578 GND.n2577 585
R10543 GND.n2574 GND.n1597 585
R10544 GND.n2574 GND.n2573 585
R10545 GND.n2319 GND.n2318 585
R10546 GND.n2331 GND.n2319 585
R10547 GND.n2329 GND.n1591 585
R10548 GND.n2564 GND.n2329 585
R10549 GND.n2552 GND.n1590 585
R10550 GND.n2552 GND.n2551 585
R10551 GND.n2553 GND.n1589 585
R10552 GND.n2554 GND.n2553 585
R10553 GND.n2549 GND.n2341 585
R10554 GND.n2549 GND.n2548 585
R10555 GND.n2340 GND.n1583 585
R10556 GND.n2354 GND.n2340 585
R10557 GND.n2352 GND.n1582 585
R10558 GND.n2539 GND.n2352 585
R10559 GND.n2526 GND.n1581 585
R10560 GND.n2526 GND.n2525 585
R10561 GND.n2528 GND.n2527 585
R10562 GND.n2529 GND.n2528 585
R10563 GND.n2524 GND.n1575 585
R10564 GND.n2524 GND.n2523 585
R10565 GND.n2363 GND.n1574 585
R10566 GND.n2506 GND.n2363 585
R10567 GND.n2504 GND.n1573 585
R10568 GND.n2514 GND.n2504 585
R10569 GND.n1553 GND.n1551 585
R10570 GND.n2423 GND.n1551 585
R10571 GND.n8079 GND.n8078 585
R10572 GND.n8080 GND.n8079 585
R10573 GND.n1552 GND.n1550 585
R10574 GND.n2370 GND.n1550 585
R10575 GND.n1566 GND.n1531 585
R10576 GND.n8086 GND.n1531 585
R10577 GND.n1565 GND.n1564 585
R10578 GND.n1564 GND.n1527 585
R10579 GND.n1563 GND.n1507 585
R10580 GND.n1512 GND.n1507 585
R10581 GND.n8095 GND.n1508 585
R10582 GND.n8095 GND.n8094 585
R10583 GND.n8097 GND.n8096 585
R10584 GND.n2387 GND.n1506 585
R10585 GND.n2390 GND.n2388 585
R10586 GND.n2392 GND.n2391 585
R10587 GND.n2394 GND.n2393 585
R10588 GND.n2384 GND.n2383 585
R10589 GND.n2398 GND.n2385 585
R10590 GND.n2400 GND.n2399 585
R10591 GND.n2402 GND.n2401 585
R10592 GND.n2380 GND.n2379 585
R10593 GND.n2406 GND.n2381 585
R10594 GND.n2407 GND.n2376 585
R10595 GND.n2408 GND.n1465 585
R10596 GND.n8151 GND.n1465 585
R10597 GND.n7837 GND.n7836 585
R10598 GND.n1882 GND.n1881 585
R10599 GND.n7844 GND.n1878 585
R10600 GND.n7845 GND.n1877 585
R10601 GND.n1876 GND.n1868 585
R10602 GND.n7852 GND.n1867 585
R10603 GND.n7853 GND.n1866 585
R10604 GND.n1860 GND.n1859 585
R10605 GND.n7860 GND.n1858 585
R10606 GND.n7861 GND.n1857 585
R10607 GND.n1856 GND.n1855 585
R10608 GND.n1833 GND.n1832 585
R10609 GND.n7873 GND.n7872 585
R10610 GND.n7881 GND.n7873 585
R10611 GND.n7832 GND.n1772 585
R10612 GND.n7924 GND.n1772 585
R10613 GND.n7831 GND.n7830 585
R10614 GND.n7830 GND.n7829 585
R10615 GND.n1890 GND.n1889 585
R10616 GND.n7826 GND.n1890 585
R10617 GND.n7809 GND.n7808 585
R10618 GND.n7808 GND.n7807 585
R10619 GND.n1908 GND.n1901 585
R10620 GND.n7818 GND.n1901 585
R10621 GND.n7814 GND.n7813 585
R10622 GND.n7815 GND.n7814 585
R10623 GND.n1907 GND.n1906 585
R10624 GND.n1916 GND.n1906 585
R10625 GND.n7803 GND.n7802 585
R10626 GND.n7802 GND.n7801 585
R10627 GND.n1911 GND.n1910 585
R10628 GND.n7788 GND.n1911 585
R10629 GND.n1931 GND.n1924 585
R10630 GND.n7791 GND.n1924 585
R10631 GND.n7785 GND.n7784 585
R10632 GND.n7786 GND.n7785 585
R10633 GND.n1930 GND.n1929 585
R10634 GND.n1939 GND.n1929 585
R10635 GND.n7779 GND.n7778 585
R10636 GND.n7778 GND.n7777 585
R10637 GND.n1934 GND.n1933 585
R10638 GND.n7764 GND.n1934 585
R10639 GND.n1953 GND.n1946 585
R10640 GND.n7767 GND.n1946 585
R10641 GND.n7760 GND.n7759 585
R10642 GND.n7761 GND.n7760 585
R10643 GND.n1952 GND.n1951 585
R10644 GND.n1962 GND.n1951 585
R10645 GND.n7754 GND.n7753 585
R10646 GND.n7753 GND.n7752 585
R10647 GND.n1956 GND.n1955 585
R10648 GND.n7738 GND.n1956 585
R10649 GND.n1975 GND.n1969 585
R10650 GND.n7742 GND.n1969 585
R10651 GND.n7735 GND.n7734 585
R10652 GND.n7736 GND.n7735 585
R10653 GND.n1974 GND.n1973 585
R10654 GND.n1984 GND.n1973 585
R10655 GND.n7729 GND.n7728 585
R10656 GND.n7728 GND.n7727 585
R10657 GND.n1978 GND.n1977 585
R10658 GND.n7714 GND.n1978 585
R10659 GND.n1998 GND.n1991 585
R10660 GND.n7717 GND.n1991 585
R10661 GND.n7710 GND.n7709 585
R10662 GND.n7711 GND.n7710 585
R10663 GND.n1997 GND.n1996 585
R10664 GND.n2007 GND.n1996 585
R10665 GND.n7704 GND.n7703 585
R10666 GND.n7703 GND.n7702 585
R10667 GND.n2001 GND.n2000 585
R10668 GND.n7689 GND.n2001 585
R10669 GND.n2022 GND.n2015 585
R10670 GND.n7692 GND.n2015 585
R10671 GND.n7686 GND.n7685 585
R10672 GND.n7687 GND.n7686 585
R10673 GND.n2021 GND.n2020 585
R10674 GND.n2030 GND.n2020 585
R10675 GND.n7680 GND.n7679 585
R10676 GND.n7679 GND.n7678 585
R10677 GND.n2025 GND.n2024 585
R10678 GND.n7665 GND.n2025 585
R10679 GND.n2049 GND.n2037 585
R10680 GND.n7668 GND.n2037 585
R10681 GND.n2888 GND.n2887 585
R10682 GND.n2889 GND.n2888 585
R10683 GND.n2048 GND.n2047 585
R10684 GND.n2047 GND.n2046 585
R10685 GND.n2882 GND.n2881 585
R10686 GND.n2881 GND.n2880 585
R10687 GND.n2052 GND.n2051 585
R10688 GND.n2866 GND.n2052 585
R10689 GND.n2071 GND.n2065 585
R10690 GND.n2870 GND.n2065 585
R10691 GND.n2863 GND.n2862 585
R10692 GND.n2864 GND.n2863 585
R10693 GND.n2070 GND.n2069 585
R10694 GND.n2080 GND.n2069 585
R10695 GND.n2857 GND.n2856 585
R10696 GND.n2856 GND.n2855 585
R10697 GND.n2074 GND.n2073 585
R10698 GND.n2842 GND.n2074 585
R10699 GND.n2094 GND.n2087 585
R10700 GND.n2845 GND.n2087 585
R10701 GND.n2838 GND.n2837 585
R10702 GND.n2839 GND.n2838 585
R10703 GND.n2093 GND.n2092 585
R10704 GND.n2103 GND.n2092 585
R10705 GND.n2832 GND.n2831 585
R10706 GND.n2831 GND.n2830 585
R10707 GND.n2097 GND.n2096 585
R10708 GND.n2791 GND.n2097 585
R10709 GND.n2782 GND.n2781 585
R10710 GND.n2788 GND.n2782 585
R10711 GND.n2187 GND.n2186 585
R10712 GND.n2186 GND.n2146 585
R10713 GND.n2777 GND.n2145 585
R10714 GND.n2800 GND.n2145 585
R10715 GND.n2776 GND.n2141 585
R10716 GND.n2803 GND.n2141 585
R10717 GND.n2775 GND.n2133 585
R10718 GND.n2808 GND.n2133 585
R10719 GND.n2768 GND.n2189 585
R10720 GND.n2768 GND.n2131 585
R10721 GND.n2770 GND.n2769 585
R10722 GND.n2769 GND.n2124 585
R10723 GND.n2767 GND.n2123 585
R10724 GND.n2817 GND.n2123 585
R10725 GND.n2766 GND.n2118 585
R10726 GND.n2820 GND.n2118 585
R10727 GND.n2195 GND.n2191 585
R10728 GND.n2666 GND.n2195 585
R10729 GND.n2762 GND.n2761 585
R10730 GND.n2761 GND.n2760 585
R10731 GND.n2194 GND.n2193 585
R10732 GND.n2749 GND.n2194 585
R10733 GND.n2213 GND.n2206 585
R10734 GND.n2752 GND.n2206 585
R10735 GND.n2746 GND.n2745 585
R10736 GND.n2747 GND.n2746 585
R10737 GND.n2212 GND.n2211 585
R10738 GND.n2221 GND.n2211 585
R10739 GND.n2740 GND.n2739 585
R10740 GND.n2739 GND.n2738 585
R10741 GND.n2216 GND.n2215 585
R10742 GND.n2725 GND.n2216 585
R10743 GND.n2235 GND.n2228 585
R10744 GND.n2728 GND.n2228 585
R10745 GND.n2721 GND.n2720 585
R10746 GND.n2722 GND.n2721 585
R10747 GND.n2234 GND.n2233 585
R10748 GND.n2244 GND.n2233 585
R10749 GND.n2715 GND.n2714 585
R10750 GND.n2714 GND.n2713 585
R10751 GND.n2238 GND.n2237 585
R10752 GND.n2699 GND.n2238 585
R10753 GND.n2620 GND.n2250 585
R10754 GND.n2703 GND.n2250 585
R10755 GND.n2623 GND.n2254 585
R10756 GND.n2697 GND.n2254 585
R10757 GND.n2624 GND.n2263 585
R10758 GND.n2644 GND.n2263 585
R10759 GND.n2625 GND.n2619 585
R10760 GND.n2619 GND.n2261 585
R10761 GND.n2276 GND.n2270 585
R10762 GND.n2636 GND.n2270 585
R10763 GND.n2630 GND.n2629 585
R10764 GND.n2631 GND.n2630 585
R10765 GND.n2275 GND.n2274 585
R10766 GND.n2285 GND.n2274 585
R10767 GND.n2615 GND.n2614 585
R10768 GND.n2614 GND.n2613 585
R10769 GND.n2279 GND.n2278 585
R10770 GND.n2600 GND.n2279 585
R10771 GND.n2299 GND.n2292 585
R10772 GND.n2603 GND.n2292 585
R10773 GND.n2596 GND.n2595 585
R10774 GND.n2597 GND.n2596 585
R10775 GND.n2298 GND.n2297 585
R10776 GND.n2308 GND.n2297 585
R10777 GND.n2590 GND.n2589 585
R10778 GND.n2589 GND.n2588 585
R10779 GND.n2302 GND.n2301 585
R10780 GND.n2575 GND.n2302 585
R10781 GND.n2323 GND.n2316 585
R10782 GND.n2578 GND.n2316 585
R10783 GND.n2572 GND.n2571 585
R10784 GND.n2573 GND.n2572 585
R10785 GND.n2322 GND.n2321 585
R10786 GND.n2331 GND.n2321 585
R10787 GND.n2566 GND.n2565 585
R10788 GND.n2565 GND.n2564 585
R10789 GND.n2326 GND.n2325 585
R10790 GND.n2551 GND.n2326 585
R10791 GND.n2345 GND.n2338 585
R10792 GND.n2554 GND.n2338 585
R10793 GND.n2547 GND.n2546 585
R10794 GND.n2548 GND.n2547 585
R10795 GND.n2344 GND.n2343 585
R10796 GND.n2354 GND.n2343 585
R10797 GND.n2541 GND.n2540 585
R10798 GND.n2540 GND.n2539 585
R10799 GND.n2348 GND.n2347 585
R10800 GND.n2525 GND.n2348 585
R10801 GND.n2367 GND.n2361 585
R10802 GND.n2529 GND.n2361 585
R10803 GND.n2522 GND.n2521 585
R10804 GND.n2523 GND.n2522 585
R10805 GND.n2366 GND.n2365 585
R10806 GND.n2506 GND.n2365 585
R10807 GND.n2516 GND.n2515 585
R10808 GND.n2515 GND.n2514 585
R10809 GND.n2422 GND.n2421 585
R10810 GND.n2423 GND.n2422 585
R10811 GND.n2420 GND.n1548 585
R10812 GND.n8080 GND.n1548 585
R10813 GND.n2372 GND.n2371 585
R10814 GND.n2371 GND.n2370 585
R10815 GND.n2416 GND.n1529 585
R10816 GND.n8086 GND.n1529 585
R10817 GND.n2415 GND.n2414 585
R10818 GND.n2414 GND.n1527 585
R10819 GND.n2413 GND.n2412 585
R10820 GND.n2413 GND.n1512 585
R10821 GND.n2374 GND.n1511 585
R10822 GND.n8094 GND.n1511 585
R10823 GND.n7923 GND.n7922 585
R10824 GND.n7924 GND.n7923 585
R10825 GND.n1777 GND.n1775 585
R10826 GND.n7829 GND.n1775 585
R10827 GND.n7825 GND.n7824 585
R10828 GND.n7826 GND.n7825 585
R10829 GND.n1896 GND.n1895 585
R10830 GND.n7807 GND.n1895 585
R10831 GND.n7820 GND.n7819 585
R10832 GND.n7819 GND.n7818 585
R10833 GND.n1899 GND.n1898 585
R10834 GND.n7815 GND.n1899 585
R10835 GND.n7798 GND.n1917 585
R10836 GND.n1917 GND.n1916 585
R10837 GND.n7800 GND.n7799 585
R10838 GND.n7801 GND.n7800 585
R10839 GND.n1918 GND.n1915 585
R10840 GND.n7788 GND.n1915 585
R10841 GND.n7793 GND.n7792 585
R10842 GND.n7792 GND.n7791 585
R10843 GND.n1921 GND.n1920 585
R10844 GND.n7786 GND.n1921 585
R10845 GND.n7774 GND.n1940 585
R10846 GND.n1940 GND.n1939 585
R10847 GND.n7776 GND.n7775 585
R10848 GND.n7777 GND.n7776 585
R10849 GND.n1941 GND.n1938 585
R10850 GND.n7764 GND.n1938 585
R10851 GND.n7769 GND.n7768 585
R10852 GND.n7768 GND.n7767 585
R10853 GND.n1944 GND.n1943 585
R10854 GND.n7761 GND.n1944 585
R10855 GND.n7749 GND.n1963 585
R10856 GND.n1963 GND.n1962 585
R10857 GND.n7751 GND.n7750 585
R10858 GND.n7752 GND.n7751 585
R10859 GND.n1964 GND.n1961 585
R10860 GND.n7738 GND.n1961 585
R10861 GND.n7744 GND.n7743 585
R10862 GND.n7743 GND.n7742 585
R10863 GND.n1967 GND.n1966 585
R10864 GND.n7736 GND.n1967 585
R10865 GND.n7724 GND.n1985 585
R10866 GND.n1985 GND.n1984 585
R10867 GND.n7726 GND.n7725 585
R10868 GND.n7727 GND.n7726 585
R10869 GND.n1986 GND.n1982 585
R10870 GND.n7714 GND.n1982 585
R10871 GND.n7719 GND.n7718 585
R10872 GND.n7718 GND.n7717 585
R10873 GND.n1989 GND.n1988 585
R10874 GND.n7711 GND.n1989 585
R10875 GND.n7699 GND.n2008 585
R10876 GND.n2008 GND.n2007 585
R10877 GND.n7701 GND.n7700 585
R10878 GND.n7702 GND.n7701 585
R10879 GND.n2009 GND.n2006 585
R10880 GND.n7689 GND.n2006 585
R10881 GND.n7694 GND.n7693 585
R10882 GND.n7693 GND.n7692 585
R10883 GND.n2012 GND.n2011 585
R10884 GND.n7687 GND.n2012 585
R10885 GND.n7675 GND.n2031 585
R10886 GND.n2031 GND.n2030 585
R10887 GND.n7677 GND.n7676 585
R10888 GND.n7678 GND.n7677 585
R10889 GND.n2032 GND.n2029 585
R10890 GND.n7665 GND.n2029 585
R10891 GND.n7670 GND.n7669 585
R10892 GND.n7669 GND.n7668 585
R10893 GND.n2035 GND.n2034 585
R10894 GND.n2889 GND.n2035 585
R10895 GND.n2877 GND.n2059 585
R10896 GND.n2059 GND.n2046 585
R10897 GND.n2879 GND.n2878 585
R10898 GND.n2880 GND.n2879 585
R10899 GND.n2060 GND.n2058 585
R10900 GND.n2866 GND.n2058 585
R10901 GND.n2872 GND.n2871 585
R10902 GND.n2871 GND.n2870 585
R10903 GND.n2063 GND.n2062 585
R10904 GND.n2864 GND.n2063 585
R10905 GND.n2852 GND.n2081 585
R10906 GND.n2081 GND.n2080 585
R10907 GND.n2854 GND.n2853 585
R10908 GND.n2855 GND.n2854 585
R10909 GND.n2082 GND.n2078 585
R10910 GND.n2842 GND.n2078 585
R10911 GND.n2847 GND.n2846 585
R10912 GND.n2846 GND.n2845 585
R10913 GND.n2085 GND.n2084 585
R10914 GND.n2839 GND.n2085 585
R10915 GND.n2827 GND.n2104 585
R10916 GND.n2104 GND.n2103 585
R10917 GND.n2829 GND.n2828 585
R10918 GND.n2830 GND.n2829 585
R10919 GND.n2105 GND.n2102 585
R10920 GND.n2791 GND.n2102 585
R10921 GND.n2787 GND.n2786 585
R10922 GND.n2788 GND.n2787 585
R10923 GND.n2785 GND.n2784 585
R10924 GND.n2785 GND.n2146 585
R10925 GND.n2783 GND.n2140 585
R10926 GND.n2800 GND.n2140 585
R10927 GND.n2805 GND.n2804 585
R10928 GND.n2804 GND.n2803 585
R10929 GND.n2807 GND.n2806 585
R10930 GND.n2808 GND.n2807 585
R10931 GND.n2139 GND.n2138 585
R10932 GND.n2139 GND.n2131 585
R10933 GND.n2137 GND.n2111 585
R10934 GND.n2137 GND.n2124 585
R10935 GND.n2115 GND.n2112 585
R10936 GND.n2817 GND.n2115 585
R10937 GND.n2822 GND.n2821 585
R10938 GND.n2821 GND.n2820 585
R10939 GND.n2114 GND.n2113 585
R10940 GND.n2666 GND.n2114 585
R10941 GND.n2759 GND.n2758 585
R10942 GND.n2760 GND.n2759 585
R10943 GND.n2200 GND.n2199 585
R10944 GND.n2749 GND.n2199 585
R10945 GND.n2754 GND.n2753 585
R10946 GND.n2753 GND.n2752 585
R10947 GND.n2203 GND.n2202 585
R10948 GND.n2747 GND.n2203 585
R10949 GND.n2735 GND.n2222 585
R10950 GND.n2222 GND.n2221 585
R10951 GND.n2737 GND.n2736 585
R10952 GND.n2738 GND.n2737 585
R10953 GND.n2223 GND.n2220 585
R10954 GND.n2725 GND.n2220 585
R10955 GND.n2730 GND.n2729 585
R10956 GND.n2729 GND.n2728 585
R10957 GND.n2226 GND.n2225 585
R10958 GND.n2722 GND.n2226 585
R10959 GND.n2710 GND.n2245 585
R10960 GND.n2245 GND.n2244 585
R10961 GND.n2712 GND.n2711 585
R10962 GND.n2713 GND.n2712 585
R10963 GND.n2246 GND.n2243 585
R10964 GND.n2699 GND.n2243 585
R10965 GND.n2705 GND.n2704 585
R10966 GND.n2704 GND.n2703 585
R10967 GND.n2249 GND.n2248 585
R10968 GND.n2697 GND.n2249 585
R10969 GND.n2643 GND.n2642 585
R10970 GND.n2644 GND.n2643 585
R10971 GND.n2265 GND.n2264 585
R10972 GND.n2264 GND.n2261 585
R10973 GND.n2638 GND.n2637 585
R10974 GND.n2637 GND.n2636 585
R10975 GND.n2268 GND.n2267 585
R10976 GND.n2631 GND.n2268 585
R10977 GND.n2610 GND.n2286 585
R10978 GND.n2286 GND.n2285 585
R10979 GND.n2612 GND.n2611 585
R10980 GND.n2613 GND.n2612 585
R10981 GND.n2287 GND.n2283 585
R10982 GND.n2600 GND.n2283 585
R10983 GND.n2605 GND.n2604 585
R10984 GND.n2604 GND.n2603 585
R10985 GND.n2290 GND.n2289 585
R10986 GND.n2597 GND.n2290 585
R10987 GND.n2585 GND.n2309 585
R10988 GND.n2309 GND.n2308 585
R10989 GND.n2587 GND.n2586 585
R10990 GND.n2588 GND.n2587 585
R10991 GND.n2310 GND.n2307 585
R10992 GND.n2575 GND.n2307 585
R10993 GND.n2580 GND.n2579 585
R10994 GND.n2579 GND.n2578 585
R10995 GND.n2313 GND.n2312 585
R10996 GND.n2573 GND.n2313 585
R10997 GND.n2561 GND.n2332 585
R10998 GND.n2332 GND.n2331 585
R10999 GND.n2563 GND.n2562 585
R11000 GND.n2564 GND.n2563 585
R11001 GND.n2333 GND.n2330 585
R11002 GND.n2551 GND.n2330 585
R11003 GND.n2556 GND.n2555 585
R11004 GND.n2555 GND.n2554 585
R11005 GND.n2336 GND.n2335 585
R11006 GND.n2548 GND.n2336 585
R11007 GND.n2536 GND.n2355 585
R11008 GND.n2355 GND.n2354 585
R11009 GND.n2538 GND.n2537 585
R11010 GND.n2539 GND.n2538 585
R11011 GND.n2356 GND.n2353 585
R11012 GND.n2525 GND.n2353 585
R11013 GND.n2531 GND.n2530 585
R11014 GND.n2530 GND.n2529 585
R11015 GND.n2359 GND.n2358 585
R11016 GND.n2523 GND.n2359 585
R11017 GND.n2511 GND.n2507 585
R11018 GND.n2507 GND.n2506 585
R11019 GND.n2513 GND.n2512 585
R11020 GND.n2514 GND.n2513 585
R11021 GND.n1545 GND.n1544 585
R11022 GND.n2423 GND.n1545 585
R11023 GND.n8082 GND.n8081 585
R11024 GND.n8081 GND.n8080 585
R11025 GND.n8083 GND.n1533 585
R11026 GND.n2370 GND.n1533 585
R11027 GND.n8085 GND.n8084 585
R11028 GND.n8086 GND.n8085 585
R11029 GND.n1534 GND.n1532 585
R11030 GND.n1532 GND.n1527 585
R11031 GND.n1538 GND.n1537 585
R11032 GND.n1537 GND.n1512 585
R11033 GND.n1536 GND.n1474 585
R11034 GND.n8094 GND.n1474 585
R11035 GND.n8149 GND.n8148 585
R11036 GND.n8147 GND.n1473 585
R11037 GND.n8146 GND.n1472 585
R11038 GND.n8151 GND.n1472 585
R11039 GND.n8145 GND.n8144 585
R11040 GND.n8143 GND.n8142 585
R11041 GND.n8141 GND.n8140 585
R11042 GND.n8139 GND.n8138 585
R11043 GND.n8137 GND.n8136 585
R11044 GND.n8135 GND.n8134 585
R11045 GND.n8133 GND.n8132 585
R11046 GND.n8131 GND.n8130 585
R11047 GND.n8129 GND.n8128 585
R11048 GND.n8127 GND.n8126 585
R11049 GND.n8125 GND.n8124 585
R11050 GND.n8123 GND.n8122 585
R11051 GND.n8121 GND.n8120 585
R11052 GND.n8119 GND.n8118 585
R11053 GND.n8117 GND.n8116 585
R11054 GND.n8115 GND.n8114 585
R11055 GND.n8113 GND.n8112 585
R11056 GND.n8111 GND.n8110 585
R11057 GND.n8109 GND.n8108 585
R11058 GND.n8107 GND.n8106 585
R11059 GND.n8105 GND.n8104 585
R11060 GND.n1503 GND.n1500 585
R11061 GND.n8100 GND.n1463 585
R11062 GND.n8151 GND.n1463 585
R11063 GND.n7885 GND.n1770 585
R11064 GND.n7886 GND.n7883 585
R11065 GND.n7887 GND.n1810 585
R11066 GND.n7888 GND.n1809 585
R11067 GND.n1822 GND.n1807 585
R11068 GND.n7892 GND.n1806 585
R11069 GND.n7893 GND.n1805 585
R11070 GND.n7894 GND.n1804 585
R11071 GND.n1819 GND.n1802 585
R11072 GND.n7898 GND.n1801 585
R11073 GND.n7899 GND.n1800 585
R11074 GND.n7900 GND.n1799 585
R11075 GND.n1816 GND.n1797 585
R11076 GND.n7904 GND.n1796 585
R11077 GND.n7881 GND.n1815 585
R11078 GND.n7906 GND.n1790 585
R11079 GND.n7907 GND.n1789 585
R11080 GND.n7875 GND.n1787 585
R11081 GND.n7911 GND.n1786 585
R11082 GND.n7912 GND.n1785 585
R11083 GND.n7913 GND.n1784 585
R11084 GND.n7878 GND.n1782 585
R11085 GND.n7917 GND.n1781 585
R11086 GND.n7918 GND.n1780 585
R11087 GND.n7919 GND.n1776 585
R11088 GND.n7881 GND.n1776 585
R11089 GND.n7926 GND.n7925 585
R11090 GND.n7925 GND.n7924 585
R11091 GND.n1769 GND.n1764 585
R11092 GND.n7829 GND.n1769 585
R11093 GND.n7930 GND.n1763 585
R11094 GND.n7826 GND.n1763 585
R11095 GND.n7931 GND.n1762 585
R11096 GND.n7807 GND.n1762 585
R11097 GND.n7932 GND.n1761 585
R11098 GND.n7818 GND.n1761 585
R11099 GND.n1905 GND.n1756 585
R11100 GND.n7815 GND.n1905 585
R11101 GND.n7936 GND.n1755 585
R11102 GND.n1916 GND.n1755 585
R11103 GND.n7937 GND.n1754 585
R11104 GND.n7801 GND.n1754 585
R11105 GND.n7938 GND.n1753 585
R11106 GND.n7788 GND.n1753 585
R11107 GND.n1923 GND.n1748 585
R11108 GND.n7791 GND.n1923 585
R11109 GND.n7942 GND.n1747 585
R11110 GND.n7786 GND.n1747 585
R11111 GND.n7943 GND.n1746 585
R11112 GND.n1939 GND.n1746 585
R11113 GND.n7944 GND.n1745 585
R11114 GND.n7777 GND.n1745 585
R11115 GND.n7763 GND.n1740 585
R11116 GND.n7764 GND.n7763 585
R11117 GND.n7948 GND.n1739 585
R11118 GND.n7767 GND.n1739 585
R11119 GND.n7949 GND.n1738 585
R11120 GND.n7761 GND.n1738 585
R11121 GND.n7950 GND.n1737 585
R11122 GND.n1962 GND.n1737 585
R11123 GND.n1958 GND.n1732 585
R11124 GND.n7752 GND.n1958 585
R11125 GND.n7954 GND.n1731 585
R11126 GND.n7738 GND.n1731 585
R11127 GND.n7955 GND.n1730 585
R11128 GND.n7742 GND.n1730 585
R11129 GND.n7956 GND.n1729 585
R11130 GND.n7736 GND.n1729 585
R11131 GND.n1983 GND.n1724 585
R11132 GND.n1984 GND.n1983 585
R11133 GND.n7960 GND.n1723 585
R11134 GND.n7727 GND.n1723 585
R11135 GND.n7961 GND.n1722 585
R11136 GND.n7714 GND.n1722 585
R11137 GND.n7962 GND.n1721 585
R11138 GND.n7717 GND.n1721 585
R11139 GND.n1995 GND.n1716 585
R11140 GND.n7711 GND.n1995 585
R11141 GND.n7966 GND.n1715 585
R11142 GND.n2007 GND.n1715 585
R11143 GND.n7967 GND.n1714 585
R11144 GND.n7702 GND.n1714 585
R11145 GND.n7968 GND.n1713 585
R11146 GND.n7689 GND.n1713 585
R11147 GND.n2014 GND.n1708 585
R11148 GND.n7692 GND.n2014 585
R11149 GND.n7972 GND.n1707 585
R11150 GND.n7687 GND.n1707 585
R11151 GND.n7973 GND.n1706 585
R11152 GND.n2030 GND.n1706 585
R11153 GND.n7974 GND.n1705 585
R11154 GND.n7678 GND.n1705 585
R11155 GND.n7664 GND.n1700 585
R11156 GND.n7665 GND.n7664 585
R11157 GND.n7978 GND.n1699 585
R11158 GND.n7668 GND.n1699 585
R11159 GND.n7979 GND.n1698 585
R11160 GND.n2889 GND.n1698 585
R11161 GND.n7980 GND.n1697 585
R11162 GND.n2046 GND.n1697 585
R11163 GND.n2054 GND.n1692 585
R11164 GND.n2880 GND.n2054 585
R11165 GND.n7984 GND.n1691 585
R11166 GND.n2866 GND.n1691 585
R11167 GND.n7985 GND.n1690 585
R11168 GND.n2870 GND.n1690 585
R11169 GND.n7986 GND.n1689 585
R11170 GND.n2864 GND.n1689 585
R11171 GND.n2079 GND.n1684 585
R11172 GND.n2080 GND.n2079 585
R11173 GND.n7990 GND.n1683 585
R11174 GND.n2855 GND.n1683 585
R11175 GND.n7991 GND.n1682 585
R11176 GND.n2842 GND.n1682 585
R11177 GND.n7992 GND.n1681 585
R11178 GND.n2845 GND.n1681 585
R11179 GND.n2091 GND.n1676 585
R11180 GND.n2839 GND.n2091 585
R11181 GND.n7996 GND.n1675 585
R11182 GND.n2103 GND.n1675 585
R11183 GND.n7997 GND.n1674 585
R11184 GND.n2830 GND.n1674 585
R11185 GND.n7998 GND.n1673 585
R11186 GND.n2791 GND.n1673 585
R11187 GND.n2185 GND.n1668 585
R11188 GND.n2788 GND.n2185 585
R11189 GND.n8002 GND.n1667 585
R11190 GND.n2146 GND.n1667 585
R11191 GND.n8003 GND.n1666 585
R11192 GND.n2800 GND.n1666 585
R11193 GND.n8004 GND.n1665 585
R11194 GND.n2803 GND.n1665 585
R11195 GND.n2132 GND.n1660 585
R11196 GND.n2808 GND.n2132 585
R11197 GND.n8008 GND.n1659 585
R11198 GND.n2131 GND.n1659 585
R11199 GND.n8009 GND.n1658 585
R11200 GND.n2124 GND.n1658 585
R11201 GND.n8010 GND.n1657 585
R11202 GND.n2817 GND.n1657 585
R11203 GND.n2117 GND.n1652 585
R11204 GND.n2820 GND.n2117 585
R11205 GND.n8014 GND.n1651 585
R11206 GND.n2666 GND.n1651 585
R11207 GND.n8015 GND.n1650 585
R11208 GND.n2760 GND.n1650 585
R11209 GND.n8016 GND.n1649 585
R11210 GND.n2749 GND.n1649 585
R11211 GND.n2205 GND.n1644 585
R11212 GND.n2752 GND.n2205 585
R11213 GND.n8020 GND.n1643 585
R11214 GND.n2747 GND.n1643 585
R11215 GND.n8021 GND.n1642 585
R11216 GND.n2221 GND.n1642 585
R11217 GND.n8022 GND.n1641 585
R11218 GND.n2738 GND.n1641 585
R11219 GND.n2724 GND.n1636 585
R11220 GND.n2725 GND.n2724 585
R11221 GND.n8026 GND.n1635 585
R11222 GND.n2728 GND.n1635 585
R11223 GND.n8027 GND.n1634 585
R11224 GND.n2722 GND.n1634 585
R11225 GND.n8028 GND.n1633 585
R11226 GND.n2244 GND.n1633 585
R11227 GND.n2240 GND.n1628 585
R11228 GND.n2713 GND.n2240 585
R11229 GND.n8032 GND.n1627 585
R11230 GND.n2699 GND.n1627 585
R11231 GND.n8033 GND.n1626 585
R11232 GND.n2703 GND.n1626 585
R11233 GND.n8034 GND.n1625 585
R11234 GND.n2697 GND.n1625 585
R11235 GND.n2262 GND.n1620 585
R11236 GND.n2644 GND.n2262 585
R11237 GND.n8038 GND.n1619 585
R11238 GND.n2261 GND.n1619 585
R11239 GND.n8039 GND.n1618 585
R11240 GND.n2636 GND.n1618 585
R11241 GND.n8040 GND.n1617 585
R11242 GND.n2631 GND.n1617 585
R11243 GND.n2284 GND.n1612 585
R11244 GND.n2285 GND.n2284 585
R11245 GND.n8044 GND.n1611 585
R11246 GND.n2613 GND.n1611 585
R11247 GND.n8045 GND.n1610 585
R11248 GND.n2600 GND.n1610 585
R11249 GND.n8046 GND.n1609 585
R11250 GND.n2603 GND.n1609 585
R11251 GND.n2296 GND.n1604 585
R11252 GND.n2597 GND.n2296 585
R11253 GND.n8050 GND.n1603 585
R11254 GND.n2308 GND.n1603 585
R11255 GND.n8051 GND.n1602 585
R11256 GND.n2588 GND.n1602 585
R11257 GND.n8052 GND.n1601 585
R11258 GND.n2575 GND.n1601 585
R11259 GND.n2315 GND.n1596 585
R11260 GND.n2578 GND.n2315 585
R11261 GND.n8056 GND.n1595 585
R11262 GND.n2573 GND.n1595 585
R11263 GND.n8057 GND.n1594 585
R11264 GND.n2331 GND.n1594 585
R11265 GND.n8058 GND.n1593 585
R11266 GND.n2564 GND.n1593 585
R11267 GND.n2550 GND.n1588 585
R11268 GND.n2551 GND.n2550 585
R11269 GND.n8062 GND.n1587 585
R11270 GND.n2554 GND.n1587 585
R11271 GND.n8063 GND.n1586 585
R11272 GND.n2548 GND.n1586 585
R11273 GND.n8064 GND.n1585 585
R11274 GND.n2354 GND.n1585 585
R11275 GND.n2350 GND.n1580 585
R11276 GND.n2539 GND.n2350 585
R11277 GND.n8068 GND.n1579 585
R11278 GND.n2525 GND.n1579 585
R11279 GND.n8069 GND.n1578 585
R11280 GND.n2529 GND.n1578 585
R11281 GND.n8070 GND.n1577 585
R11282 GND.n2523 GND.n1577 585
R11283 GND.n2505 GND.n1572 585
R11284 GND.n2506 GND.n2505 585
R11285 GND.n8074 GND.n1571 585
R11286 GND.n2514 GND.n1571 585
R11287 GND.n8075 GND.n1570 585
R11288 GND.n2423 GND.n1570 585
R11289 GND.n8076 GND.n1547 585
R11290 GND.n8080 GND.n1547 585
R11291 GND.n2369 GND.n1569 585
R11292 GND.n2370 GND.n2369 585
R11293 GND.n1568 GND.n1528 585
R11294 GND.n8086 GND.n1528 585
R11295 GND.n1559 GND.n1556 585
R11296 GND.n1559 GND.n1527 585
R11297 GND.n1561 GND.n1560 585
R11298 GND.n1560 GND.n1512 585
R11299 GND.n1558 GND.n1510 585
R11300 GND.n8094 GND.n1510 585
R11301 GND.n9611 GND.n9610 585
R11302 GND.n9612 GND.n9611 585
R11303 GND.n482 GND.n480 585
R11304 GND.n9524 GND.n480 585
R11305 GND.n9513 GND.n562 585
R11306 GND.n562 GND.n561 585
R11307 GND.n9515 GND.n9514 585
R11308 GND.n9516 GND.n9515 585
R11309 GND.n563 GND.n560 585
R11310 GND.n572 GND.n560 585
R11311 GND.n9508 GND.n9507 585
R11312 GND.n9507 GND.n9506 585
R11313 GND.n566 GND.n565 585
R11314 GND.n9499 GND.n566 585
R11315 GND.n7096 GND.n3573 585
R11316 GND.n3573 GND.n579 585
R11317 GND.n7098 GND.n7097 585
R11318 GND.n7099 GND.n7098 585
R11319 GND.n3574 GND.n3572 585
R11320 GND.n3580 GND.n3572 585
R11321 GND.n7091 GND.n7090 585
R11322 GND.n7090 GND.n7089 585
R11323 GND.n3577 GND.n3576 585
R11324 GND.n7085 GND.n3577 585
R11325 GND.n7063 GND.n3596 585
R11326 GND.n3596 GND.n3584 585
R11327 GND.n7065 GND.n7064 585
R11328 GND.n7066 GND.n7065 585
R11329 GND.n3597 GND.n3595 585
R11330 GND.n3595 GND.n3591 585
R11331 GND.n7058 GND.n7057 585
R11332 GND.n7057 GND.n7056 585
R11333 GND.n3600 GND.n3599 585
R11334 GND.n7051 GND.n3600 585
R11335 GND.n7035 GND.n3617 585
R11336 GND.n3617 GND.n3605 585
R11337 GND.n7037 GND.n7036 585
R11338 GND.n7038 GND.n7037 585
R11339 GND.n3618 GND.n3616 585
R11340 GND.n3616 GND.n3612 585
R11341 GND.n7030 GND.n7029 585
R11342 GND.n7029 GND.n7028 585
R11343 GND.n3621 GND.n3620 585
R11344 GND.n7024 GND.n3621 585
R11345 GND.n7008 GND.n3639 585
R11346 GND.n3639 GND.n3627 585
R11347 GND.n7010 GND.n7009 585
R11348 GND.n7011 GND.n7010 585
R11349 GND.n3640 GND.n3638 585
R11350 GND.n3638 GND.n3635 585
R11351 GND.n7003 GND.n7002 585
R11352 GND.n7002 GND.n7001 585
R11353 GND.n3643 GND.n3642 585
R11354 GND.n6997 GND.n3643 585
R11355 GND.n6982 GND.n3662 585
R11356 GND.n3662 GND.n3649 585
R11357 GND.n6984 GND.n6983 585
R11358 GND.n6985 GND.n6984 585
R11359 GND.n3663 GND.n3661 585
R11360 GND.n3661 GND.n3657 585
R11361 GND.n6977 GND.n6976 585
R11362 GND.n6976 GND.n6975 585
R11363 GND.n3666 GND.n3665 585
R11364 GND.n6970 GND.n3666 585
R11365 GND.n6955 GND.n3682 585
R11366 GND.n3682 GND.n3671 585
R11367 GND.n6957 GND.n6956 585
R11368 GND.n6958 GND.n6957 585
R11369 GND.n3683 GND.n3681 585
R11370 GND.n6945 GND.n3681 585
R11371 GND.n6950 GND.n6949 585
R11372 GND.n6949 GND.n6948 585
R11373 GND.n3686 GND.n3685 585
R11374 GND.n6942 GND.n3686 585
R11375 GND.n6926 GND.n3703 585
R11376 GND.n3703 GND.n3691 585
R11377 GND.n6928 GND.n6927 585
R11378 GND.n6929 GND.n6928 585
R11379 GND.n3704 GND.n3702 585
R11380 GND.n3702 GND.n3698 585
R11381 GND.n6921 GND.n6920 585
R11382 GND.n6920 GND.n6919 585
R11383 GND.n3707 GND.n3706 585
R11384 GND.n6915 GND.n3707 585
R11385 GND.n6899 GND.n3725 585
R11386 GND.n3725 GND.n3713 585
R11387 GND.n6901 GND.n6900 585
R11388 GND.n6902 GND.n6901 585
R11389 GND.n3726 GND.n3724 585
R11390 GND.n3724 GND.n3721 585
R11391 GND.n6894 GND.n6893 585
R11392 GND.n6893 GND.n6892 585
R11393 GND.n3729 GND.n3728 585
R11394 GND.n6888 GND.n3729 585
R11395 GND.n6837 GND.n6834 585
R11396 GND.n6834 GND.n3735 585
R11397 GND.n6839 GND.n6838 585
R11398 GND.n6840 GND.n6839 585
R11399 GND.n6835 GND.n6825 585
R11400 GND.n6849 GND.n6825 585
R11401 GND.n6855 GND.n6854 585
R11402 GND.n6854 GND.n6853 585
R11403 GND.n6856 GND.n6821 585
R11404 GND.n6828 GND.n6821 585
R11405 GND.n6859 GND.n6858 585
R11406 GND.n6860 GND.n6859 585
R11407 GND.n6823 GND.n6820 585
R11408 GND.n6820 GND.n6811 585
R11409 GND.n3758 GND.n3757 585
R11410 GND.n6867 GND.n3758 585
R11411 GND.n6872 GND.n6871 585
R11412 GND.n6871 GND.n6870 585
R11413 GND.n6873 GND.n3755 585
R11414 GND.n6802 GND.n3755 585
R11415 GND.n6876 GND.n6875 585
R11416 GND.n6877 GND.n6876 585
R11417 GND.n3756 GND.n3754 585
R11418 GND.n3754 GND.n3750 585
R11419 GND.n6790 GND.n3783 585
R11420 GND.n3783 GND.n3782 585
R11421 GND.n6792 GND.n6791 585
R11422 GND.n6793 GND.n6792 585
R11423 GND.n3784 GND.n3777 585
R11424 GND.n6778 GND.n3777 585
R11425 GND.n6784 GND.n6783 585
R11426 GND.n6783 GND.n6782 585
R11427 GND.n3787 GND.n3786 585
R11428 GND.n6776 GND.n3787 585
R11429 GND.n6764 GND.n3805 585
R11430 GND.n3805 GND.n3804 585
R11431 GND.n6766 GND.n6765 585
R11432 GND.n6767 GND.n6766 585
R11433 GND.n3806 GND.n3802 585
R11434 GND.n6754 GND.n3802 585
R11435 GND.n6759 GND.n6758 585
R11436 GND.n6758 GND.n6757 585
R11437 GND.n3809 GND.n3808 585
R11438 GND.n6751 GND.n3809 585
R11439 GND.n6739 GND.n3828 585
R11440 GND.n3828 GND.n3827 585
R11441 GND.n6741 GND.n6740 585
R11442 GND.n6742 GND.n6741 585
R11443 GND.n3829 GND.n3826 585
R11444 GND.n6729 GND.n3826 585
R11445 GND.n6734 GND.n6733 585
R11446 GND.n6733 GND.n6732 585
R11447 GND.n3832 GND.n3831 585
R11448 GND.n6727 GND.n3832 585
R11449 GND.n6715 GND.n3851 585
R11450 GND.n3851 GND.n3850 585
R11451 GND.n6717 GND.n6716 585
R11452 GND.n6718 GND.n6717 585
R11453 GND.n3852 GND.n3849 585
R11454 GND.n6705 GND.n3849 585
R11455 GND.n6710 GND.n6709 585
R11456 GND.n6709 GND.n6708 585
R11457 GND.n3855 GND.n3854 585
R11458 GND.n6702 GND.n3855 585
R11459 GND.n6690 GND.n3874 585
R11460 GND.n3874 GND.n3873 585
R11461 GND.n6692 GND.n6691 585
R11462 GND.n6693 GND.n6692 585
R11463 GND.n3875 GND.n3872 585
R11464 GND.n6679 GND.n3872 585
R11465 GND.n6685 GND.n6684 585
R11466 GND.n6684 GND.n6683 585
R11467 GND.n3878 GND.n3877 585
R11468 GND.n6677 GND.n3878 585
R11469 GND.n6665 GND.n3896 585
R11470 GND.n3896 GND.n3895 585
R11471 GND.n6667 GND.n6666 585
R11472 GND.n6668 GND.n6667 585
R11473 GND.n3897 GND.n3893 585
R11474 GND.n6655 GND.n3893 585
R11475 GND.n6660 GND.n6659 585
R11476 GND.n6659 GND.n6658 585
R11477 GND.n3900 GND.n3899 585
R11478 GND.n6652 GND.n3900 585
R11479 GND.n6640 GND.n3919 585
R11480 GND.n3919 GND.n3918 585
R11481 GND.n6642 GND.n6641 585
R11482 GND.n6643 GND.n6642 585
R11483 GND.n3920 GND.n3917 585
R11484 GND.n6630 GND.n3917 585
R11485 GND.n6635 GND.n6634 585
R11486 GND.n6634 GND.n6633 585
R11487 GND.n3923 GND.n3922 585
R11488 GND.n6628 GND.n3923 585
R11489 GND.n6616 GND.n3942 585
R11490 GND.n3942 GND.n3941 585
R11491 GND.n6618 GND.n6617 585
R11492 GND.n6619 GND.n6618 585
R11493 GND.n3943 GND.n3940 585
R11494 GND.n6606 GND.n3940 585
R11495 GND.n6611 GND.n6610 585
R11496 GND.n6610 GND.n6609 585
R11497 GND.n3946 GND.n3945 585
R11498 GND.n6603 GND.n3946 585
R11499 GND.n6591 GND.n6585 585
R11500 GND.n6585 GND.n6584 585
R11501 GND.n6593 GND.n6592 585
R11502 GND.n6594 GND.n6593 585
R11503 GND.n6586 GND.n6583 585
R11504 GND.n6583 GND.n6582 585
R11505 GND.n3365 GND.n3364 585
R11506 GND.n6437 GND.n3365 585
R11507 GND.n7252 GND.n7251 585
R11508 GND.n7251 GND.n7250 585
R11509 GND.n7253 GND.n3360 585
R11510 GND.n3376 GND.n3360 585
R11511 GND.n7255 GND.n7254 585
R11512 GND.n7256 GND.n7255 585
R11513 GND.n6266 GND.n3359 585
R11514 GND.n6270 GND.n6265 585
R11515 GND.n6272 GND.n6271 585
R11516 GND.n6274 GND.n6273 585
R11517 GND.n6276 GND.n6275 585
R11518 GND.n6280 GND.n6263 585
R11519 GND.n6282 GND.n6281 585
R11520 GND.n6284 GND.n6283 585
R11521 GND.n6286 GND.n6285 585
R11522 GND.n6119 GND.n6118 585
R11523 GND.n7293 GND.n3297 585
R11524 GND.n6294 GND.n6293 585
R11525 GND.n6296 GND.n6295 585
R11526 GND.n6300 GND.n6116 585
R11527 GND.n6302 GND.n6301 585
R11528 GND.n6304 GND.n6303 585
R11529 GND.n6306 GND.n6305 585
R11530 GND.n6310 GND.n6114 585
R11531 GND.n6312 GND.n6311 585
R11532 GND.n6314 GND.n6313 585
R11533 GND.n6316 GND.n6315 585
R11534 GND.n6111 GND.n6110 585
R11535 GND.n6320 GND.n6112 585
R11536 GND.n6321 GND.n6107 585
R11537 GND.n6322 GND.n3305 585
R11538 GND.n7293 GND.n3305 585
R11539 GND.n9570 GND.n9569 585
R11540 GND.n9571 GND.n518 585
R11541 GND.n536 GND.n514 585
R11542 GND.n9575 GND.n513 585
R11543 GND.n9576 GND.n512 585
R11544 GND.n9577 GND.n511 585
R11545 GND.n533 GND.n509 585
R11546 GND.n9581 GND.n508 585
R11547 GND.n9582 GND.n507 585
R11548 GND.n9583 GND.n506 585
R11549 GND.n530 GND.n504 585
R11550 GND.n9587 GND.n503 585
R11551 GND.n9588 GND.n502 585
R11552 GND.n9589 GND.n501 585
R11553 GND.n527 GND.n499 585
R11554 GND.n9593 GND.n496 585
R11555 GND.n9594 GND.n495 585
R11556 GND.n9595 GND.n494 585
R11557 GND.n524 GND.n492 585
R11558 GND.n9599 GND.n491 585
R11559 GND.n9600 GND.n490 585
R11560 GND.n9601 GND.n489 585
R11561 GND.n521 GND.n487 585
R11562 GND.n9605 GND.n486 585
R11563 GND.n9606 GND.n485 585
R11564 GND.n9607 GND.n481 585
R11565 GND.n9527 GND.n477 585
R11566 GND.n9612 GND.n477 585
R11567 GND.n9526 GND.n9525 585
R11568 GND.n9525 GND.n9524 585
R11569 GND.n550 GND.n549 585
R11570 GND.n561 GND.n550 585
R11571 GND.n9518 GND.n9517 585
R11572 GND.n9517 GND.n9516 585
R11573 GND.n556 GND.n555 585
R11574 GND.n572 GND.n556 585
R11575 GND.n9502 GND.n568 585
R11576 GND.n9506 GND.n568 585
R11577 GND.n9501 GND.n9500 585
R11578 GND.n9500 GND.n9499 585
R11579 GND.n578 GND.n577 585
R11580 GND.n579 GND.n578 585
R11581 GND.n3570 GND.n3565 585
R11582 GND.n7099 GND.n3570 585
R11583 GND.n7106 GND.n3564 585
R11584 GND.n3580 GND.n3564 585
R11585 GND.n7107 GND.n3563 585
R11586 GND.n7089 GND.n3563 585
R11587 GND.n7108 GND.n3562 585
R11588 GND.n7085 GND.n3562 585
R11589 GND.n3583 GND.n3557 585
R11590 GND.n3584 GND.n3583 585
R11591 GND.n7112 GND.n3556 585
R11592 GND.n7066 GND.n3556 585
R11593 GND.n7113 GND.n3555 585
R11594 GND.n3591 GND.n3555 585
R11595 GND.n7114 GND.n3554 585
R11596 GND.n7056 GND.n3554 585
R11597 GND.n7050 GND.n3549 585
R11598 GND.n7051 GND.n7050 585
R11599 GND.n7118 GND.n3548 585
R11600 GND.n3605 GND.n3548 585
R11601 GND.n7119 GND.n3547 585
R11602 GND.n7038 GND.n3547 585
R11603 GND.n7120 GND.n3546 585
R11604 GND.n3612 GND.n3546 585
R11605 GND.n3623 GND.n3541 585
R11606 GND.n7028 GND.n3623 585
R11607 GND.n7124 GND.n3540 585
R11608 GND.n7024 GND.n3540 585
R11609 GND.n7125 GND.n3539 585
R11610 GND.n3627 GND.n3539 585
R11611 GND.n7126 GND.n3538 585
R11612 GND.n7011 GND.n3538 585
R11613 GND.n3634 GND.n3533 585
R11614 GND.n3635 GND.n3634 585
R11615 GND.n7130 GND.n3532 585
R11616 GND.n7001 GND.n3532 585
R11617 GND.n7131 GND.n3531 585
R11618 GND.n6997 GND.n3531 585
R11619 GND.n7132 GND.n3530 585
R11620 GND.n3649 GND.n3530 585
R11621 GND.n3658 GND.n3525 585
R11622 GND.n6985 GND.n3658 585
R11623 GND.n7136 GND.n3524 585
R11624 GND.n3657 GND.n3524 585
R11625 GND.n7137 GND.n3523 585
R11626 GND.n6975 GND.n3523 585
R11627 GND.n7138 GND.n3522 585
R11628 GND.n6970 GND.n3522 585
R11629 GND.n3670 GND.n3517 585
R11630 GND.n3671 GND.n3670 585
R11631 GND.n7142 GND.n3516 585
R11632 GND.n6958 GND.n3516 585
R11633 GND.n7143 GND.n3515 585
R11634 GND.n6945 GND.n3515 585
R11635 GND.n7144 GND.n3514 585
R11636 GND.n6948 GND.n3514 585
R11637 GND.n6941 GND.n3509 585
R11638 GND.n6942 GND.n6941 585
R11639 GND.n7148 GND.n3508 585
R11640 GND.n3691 GND.n3508 585
R11641 GND.n7149 GND.n3507 585
R11642 GND.n6929 GND.n3507 585
R11643 GND.n7150 GND.n3506 585
R11644 GND.n3698 GND.n3506 585
R11645 GND.n3709 GND.n3501 585
R11646 GND.n6919 GND.n3709 585
R11647 GND.n7154 GND.n3500 585
R11648 GND.n6915 GND.n3500 585
R11649 GND.n7155 GND.n3499 585
R11650 GND.n3713 GND.n3499 585
R11651 GND.n7156 GND.n3498 585
R11652 GND.n6902 GND.n3498 585
R11653 GND.n3720 GND.n3493 585
R11654 GND.n3721 GND.n3720 585
R11655 GND.n7160 GND.n3492 585
R11656 GND.n6892 GND.n3492 585
R11657 GND.n7161 GND.n3491 585
R11658 GND.n6888 GND.n3491 585
R11659 GND.n7162 GND.n3490 585
R11660 GND.n3735 GND.n3490 585
R11661 GND.n6832 GND.n3485 585
R11662 GND.n6840 GND.n6832 585
R11663 GND.n7166 GND.n3484 585
R11664 GND.n6849 GND.n3484 585
R11665 GND.n7167 GND.n3483 585
R11666 GND.n6853 GND.n3483 585
R11667 GND.n7168 GND.n3482 585
R11668 GND.n6828 GND.n3482 585
R11669 GND.n6817 GND.n3477 585
R11670 GND.n6860 GND.n6817 585
R11671 GND.n7172 GND.n3476 585
R11672 GND.n6811 GND.n3476 585
R11673 GND.n7173 GND.n3475 585
R11674 GND.n6867 GND.n3475 585
R11675 GND.n7174 GND.n3474 585
R11676 GND.n6870 GND.n3474 585
R11677 GND.n6801 GND.n3469 585
R11678 GND.n6802 GND.n6801 585
R11679 GND.n7178 GND.n3468 585
R11680 GND.n6877 GND.n3468 585
R11681 GND.n7179 GND.n3467 585
R11682 GND.n3750 GND.n3467 585
R11683 GND.n7180 GND.n3466 585
R11684 GND.n3782 GND.n3466 585
R11685 GND.n3774 GND.n3461 585
R11686 GND.n6793 GND.n3774 585
R11687 GND.n7184 GND.n3460 585
R11688 GND.n6778 GND.n3460 585
R11689 GND.n7185 GND.n3459 585
R11690 GND.n6782 GND.n3459 585
R11691 GND.n7186 GND.n3458 585
R11692 GND.n6776 GND.n3458 585
R11693 GND.n3803 GND.n3453 585
R11694 GND.n3804 GND.n3803 585
R11695 GND.n7190 GND.n3452 585
R11696 GND.n6767 GND.n3452 585
R11697 GND.n7191 GND.n3451 585
R11698 GND.n6754 GND.n3451 585
R11699 GND.n7192 GND.n3450 585
R11700 GND.n6757 GND.n3450 585
R11701 GND.n3815 GND.n3445 585
R11702 GND.n6751 GND.n3815 585
R11703 GND.n7196 GND.n3444 585
R11704 GND.n3827 GND.n3444 585
R11705 GND.n7197 GND.n3443 585
R11706 GND.n6742 GND.n3443 585
R11707 GND.n7198 GND.n3442 585
R11708 GND.n6729 GND.n3442 585
R11709 GND.n3834 GND.n3437 585
R11710 GND.n6732 GND.n3834 585
R11711 GND.n7202 GND.n3436 585
R11712 GND.n6727 GND.n3436 585
R11713 GND.n7203 GND.n3435 585
R11714 GND.n3850 GND.n3435 585
R11715 GND.n7204 GND.n3434 585
R11716 GND.n6718 GND.n3434 585
R11717 GND.n6704 GND.n3429 585
R11718 GND.n6705 GND.n6704 585
R11719 GND.n7208 GND.n3428 585
R11720 GND.n6708 GND.n3428 585
R11721 GND.n7209 GND.n3427 585
R11722 GND.n6702 GND.n3427 585
R11723 GND.n7210 GND.n3426 585
R11724 GND.n3873 GND.n3426 585
R11725 GND.n3869 GND.n3421 585
R11726 GND.n6693 GND.n3869 585
R11727 GND.n7214 GND.n3420 585
R11728 GND.n6679 GND.n3420 585
R11729 GND.n7215 GND.n3419 585
R11730 GND.n6683 GND.n3419 585
R11731 GND.n7216 GND.n3418 585
R11732 GND.n6677 GND.n3418 585
R11733 GND.n3894 GND.n3413 585
R11734 GND.n3895 GND.n3894 585
R11735 GND.n7220 GND.n3412 585
R11736 GND.n6668 GND.n3412 585
R11737 GND.n7221 GND.n3411 585
R11738 GND.n6655 GND.n3411 585
R11739 GND.n7222 GND.n3410 585
R11740 GND.n6658 GND.n3410 585
R11741 GND.n3906 GND.n3405 585
R11742 GND.n6652 GND.n3906 585
R11743 GND.n7226 GND.n3404 585
R11744 GND.n3918 GND.n3404 585
R11745 GND.n7227 GND.n3403 585
R11746 GND.n6643 GND.n3403 585
R11747 GND.n7228 GND.n3402 585
R11748 GND.n6630 GND.n3402 585
R11749 GND.n3925 GND.n3397 585
R11750 GND.n6633 GND.n3925 585
R11751 GND.n7232 GND.n3396 585
R11752 GND.n6628 GND.n3396 585
R11753 GND.n7233 GND.n3395 585
R11754 GND.n3941 GND.n3395 585
R11755 GND.n7234 GND.n3394 585
R11756 GND.n6619 GND.n3394 585
R11757 GND.n6605 GND.n3389 585
R11758 GND.n6606 GND.n6605 585
R11759 GND.n7238 GND.n3388 585
R11760 GND.n6609 GND.n3388 585
R11761 GND.n7239 GND.n3387 585
R11762 GND.n6603 GND.n3387 585
R11763 GND.n7240 GND.n3386 585
R11764 GND.n6584 GND.n3386 585
R11765 GND.n3959 GND.n3381 585
R11766 GND.n6594 GND.n3959 585
R11767 GND.n7244 GND.n3380 585
R11768 GND.n6582 GND.n3380 585
R11769 GND.n7245 GND.n3379 585
R11770 GND.n6437 GND.n3379 585
R11771 GND.n7246 GND.n3367 585
R11772 GND.n7250 GND.n3367 585
R11773 GND.n3378 GND.n3377 585
R11774 GND.n3377 GND.n3376 585
R11775 GND.n6325 GND.n3357 585
R11776 GND.n7256 GND.n3357 585
R11777 GND.n3270 GND.n3269 585
R11778 GND.n6140 GND.n3270 585
R11779 GND.n7311 GND.n7310 585
R11780 GND.n7310 GND.n7309 585
R11781 GND.n7312 GND.n3267 585
R11782 GND.n3271 GND.n3267 585
R11783 GND.n7314 GND.n7313 585
R11784 GND.n7315 GND.n7314 585
R11785 GND.n3268 GND.n3266 585
R11786 GND.n3266 GND.n3259 585
R11787 GND.n6373 GND.n3258 585
R11788 GND.n7321 GND.n3258 585
R11789 GND.n6375 GND.n6374 585
R11790 GND.n6376 GND.n6375 585
R11791 GND.n3248 GND.n3247 585
R11792 GND.n6378 GND.n3248 585
R11793 GND.n7330 GND.n7329 585
R11794 GND.n7329 GND.n7328 585
R11795 GND.n7331 GND.n3245 585
R11796 GND.n3249 GND.n3245 585
R11797 GND.n7333 GND.n7332 585
R11798 GND.n7334 GND.n7333 585
R11799 GND.n3246 GND.n3244 585
R11800 GND.n3244 GND.n3241 585
R11801 GND.n6399 GND.n6398 585
R11802 GND.n6400 GND.n6399 585
R11803 GND.n6397 GND.n3975 585
R11804 GND.n3975 GND.n3232 585
R11805 GND.n6396 GND.n6395 585
R11806 GND.n6395 GND.n3230 585
R11807 GND.n6394 GND.n3976 585
R11808 GND.n6394 GND.n6393 585
R11809 GND.n6366 GND.n3977 585
R11810 GND.n3984 GND.n3977 585
R11811 GND.n6368 GND.n6367 585
R11812 GND.n6369 GND.n6368 585
R11813 GND.n6365 GND.n3986 585
R11814 GND.n3986 GND.n3983 585
R11815 GND.n6364 GND.n6363 585
R11816 GND.n6363 GND.n6362 585
R11817 GND.n3988 GND.n3987 585
R11818 GND.n6055 GND.n3988 585
R11819 GND.n6347 GND.n6346 585
R11820 GND.n6348 GND.n6347 585
R11821 GND.n6345 GND.n4001 585
R11822 GND.n4001 GND.n3998 585
R11823 GND.n6344 GND.n6343 585
R11824 GND.n6343 GND.n6342 585
R11825 GND.n4003 GND.n4002 585
R11826 GND.n4004 GND.n4003 585
R11827 GND.n6078 GND.n6077 585
R11828 GND.n6078 GND.n4012 585
R11829 GND.n6080 GND.n6079 585
R11830 GND.n6079 GND.n4011 585
R11831 GND.n6081 GND.n4026 585
R11832 GND.n6066 GND.n4026 585
R11833 GND.n6083 GND.n6082 585
R11834 GND.n6084 GND.n6083 585
R11835 GND.n6076 GND.n4025 585
R11836 GND.n4025 GND.n4020 585
R11837 GND.n6075 GND.n6074 585
R11838 GND.n6074 GND.n6073 585
R11839 GND.n4028 GND.n4027 585
R11840 GND.n4029 GND.n4028 585
R11841 GND.n6047 GND.n6046 585
R11842 GND.n6048 GND.n6047 585
R11843 GND.n6045 GND.n4038 585
R11844 GND.n6041 GND.n4038 585
R11845 GND.n6044 GND.n6043 585
R11846 GND.n6043 GND.n6042 585
R11847 GND.n4040 GND.n4039 585
R11848 GND.n4046 GND.n4040 585
R11849 GND.n6034 GND.n6033 585
R11850 GND.n6035 GND.n6034 585
R11851 GND.n6032 GND.n4048 585
R11852 GND.n4048 GND.n4045 585
R11853 GND.n6031 GND.n6030 585
R11854 GND.n6030 GND.n6029 585
R11855 GND.n4050 GND.n4049 585
R11856 GND.n4064 GND.n4050 585
R11857 GND.n6007 GND.n6006 585
R11858 GND.n6008 GND.n6007 585
R11859 GND.n6005 GND.n4065 585
R11860 GND.n4065 GND.n4061 585
R11861 GND.n6004 GND.n6003 585
R11862 GND.n6003 GND.n6002 585
R11863 GND.n4067 GND.n4066 585
R11864 GND.n4068 GND.n4067 585
R11865 GND.n5953 GND.n5952 585
R11866 GND.n5953 GND.n4076 585
R11867 GND.n5955 GND.n5954 585
R11868 GND.n5954 GND.n4075 585
R11869 GND.n5956 GND.n4090 585
R11870 GND.n5941 GND.n4090 585
R11871 GND.n5958 GND.n5957 585
R11872 GND.n5959 GND.n5958 585
R11873 GND.n5951 GND.n4089 585
R11874 GND.n4089 GND.n4085 585
R11875 GND.n5950 GND.n5949 585
R11876 GND.n5949 GND.n5948 585
R11877 GND.n4092 GND.n4091 585
R11878 GND.n4098 GND.n4092 585
R11879 GND.n5923 GND.n5922 585
R11880 GND.n5924 GND.n5923 585
R11881 GND.n5921 GND.n4101 585
R11882 GND.n4107 GND.n4101 585
R11883 GND.n5920 GND.n5919 585
R11884 GND.n5919 GND.n5918 585
R11885 GND.n4103 GND.n4102 585
R11886 GND.n4117 GND.n4103 585
R11887 GND.n5895 GND.n4115 585
R11888 GND.n5907 GND.n4115 585
R11889 GND.n5896 GND.n4126 585
R11890 GND.n4126 GND.n4114 585
R11891 GND.n5898 GND.n5897 585
R11892 GND.n5899 GND.n5898 585
R11893 GND.n5894 GND.n4125 585
R11894 GND.n5890 GND.n4125 585
R11895 GND.n5893 GND.n5892 585
R11896 GND.n5892 GND.n5891 585
R11897 GND.n4128 GND.n4127 585
R11898 GND.n4134 GND.n4128 585
R11899 GND.n5883 GND.n5882 585
R11900 GND.n5884 GND.n5883 585
R11901 GND.n5881 GND.n4136 585
R11902 GND.n4136 GND.n4133 585
R11903 GND.n5880 GND.n5879 585
R11904 GND.n5879 GND.n5878 585
R11905 GND.n4138 GND.n4137 585
R11906 GND.n4151 GND.n4138 585
R11907 GND.n5859 GND.n5858 585
R11908 GND.n5860 GND.n5859 585
R11909 GND.n5857 GND.n4152 585
R11910 GND.n5852 GND.n4152 585
R11911 GND.n5856 GND.n5855 585
R11912 GND.n5855 GND.n5854 585
R11913 GND.n4154 GND.n4153 585
R11914 GND.n4155 GND.n4154 585
R11915 GND.n5840 GND.n5839 585
R11916 GND.n5841 GND.n5840 585
R11917 GND.n5838 GND.n4163 585
R11918 GND.n5834 GND.n4163 585
R11919 GND.n5837 GND.n5836 585
R11920 GND.n5836 GND.n5835 585
R11921 GND.n4165 GND.n4164 585
R11922 GND.n4171 GND.n4165 585
R11923 GND.n5826 GND.n5825 585
R11924 GND.n5827 GND.n5826 585
R11925 GND.n5824 GND.n4173 585
R11926 GND.n4173 GND.n4170 585
R11927 GND.n5823 GND.n5822 585
R11928 GND.n5822 GND.n5821 585
R11929 GND.n4175 GND.n4174 585
R11930 GND.n4189 GND.n4175 585
R11931 GND.n5799 GND.n5798 585
R11932 GND.n5800 GND.n5799 585
R11933 GND.n5797 GND.n4190 585
R11934 GND.n4190 GND.n4186 585
R11935 GND.n5796 GND.n5795 585
R11936 GND.n5795 GND.n5794 585
R11937 GND.n4192 GND.n4191 585
R11938 GND.n4194 GND.n4192 585
R11939 GND.n5713 GND.n5712 585
R11940 GND.n5713 GND.n4202 585
R11941 GND.n5715 GND.n5714 585
R11942 GND.n5714 GND.n4201 585
R11943 GND.n5716 GND.n4215 585
R11944 GND.n4215 GND.n4213 585
R11945 GND.n5718 GND.n5717 585
R11946 GND.n5719 GND.n5718 585
R11947 GND.n5711 GND.n4214 585
R11948 GND.n4214 GND.n4209 585
R11949 GND.n5710 GND.n5709 585
R11950 GND.n5709 GND.n5708 585
R11951 GND.n4217 GND.n4216 585
R11952 GND.n4218 GND.n4217 585
R11953 GND.n5678 GND.n4239 585
R11954 GND.n5678 GND.n5677 585
R11955 GND.n5680 GND.n5679 585
R11956 GND.n5679 GND.n4225 585
R11957 GND.n5681 GND.n4237 585
R11958 GND.n5650 GND.n4237 585
R11959 GND.n5683 GND.n5682 585
R11960 GND.n5684 GND.n5683 585
R11961 GND.n4238 GND.n4236 585
R11962 GND.n4236 GND.n4232 585
R11963 GND.n5644 GND.n5643 585
R11964 GND.n5645 GND.n5644 585
R11965 GND.n5642 GND.n4245 585
R11966 GND.n4250 GND.n4245 585
R11967 GND.n5641 GND.n5640 585
R11968 GND.n5640 GND.n5639 585
R11969 GND.n4247 GND.n4246 585
R11970 GND.n5615 GND.n4247 585
R11971 GND.n5627 GND.n5626 585
R11972 GND.n5628 GND.n5627 585
R11973 GND.n5625 GND.n4260 585
R11974 GND.n4260 GND.n4256 585
R11975 GND.n5624 GND.n5623 585
R11976 GND.n5623 GND.n5622 585
R11977 GND.n4262 GND.n4261 585
R11978 GND.n4269 GND.n4262 585
R11979 GND.n5608 GND.n5607 585
R11980 GND.n5609 GND.n5608 585
R11981 GND.n5606 GND.n4271 585
R11982 GND.n4271 GND.n4268 585
R11983 GND.n5605 GND.n5604 585
R11984 GND.n5604 GND.n5603 585
R11985 GND.n4273 GND.n4272 585
R11986 GND.n4287 GND.n4273 585
R11987 GND.n5580 GND.n4285 585
R11988 GND.n5592 GND.n4285 585
R11989 GND.n5581 GND.n4294 585
R11990 GND.n4294 GND.n4284 585
R11991 GND.n5583 GND.n5582 585
R11992 GND.n5584 GND.n5583 585
R11993 GND.n5579 GND.n4293 585
R11994 GND.n5575 GND.n4293 585
R11995 GND.n5578 GND.n5577 585
R11996 GND.n5577 GND.n5576 585
R11997 GND.n4296 GND.n4295 585
R11998 GND.n4303 GND.n4296 585
R11999 GND.n5568 GND.n5567 585
R12000 GND.n5569 GND.n5568 585
R12001 GND.n5566 GND.n4305 585
R12002 GND.n4305 GND.n4302 585
R12003 GND.n5565 GND.n5564 585
R12004 GND.n5564 GND.n5563 585
R12005 GND.n4307 GND.n4306 585
R12006 GND.n4320 GND.n4307 585
R12007 GND.n5543 GND.n5542 585
R12008 GND.n5544 GND.n5543 585
R12009 GND.n5541 GND.n4321 585
R12010 GND.n4321 GND.n4317 585
R12011 GND.n5540 GND.n5539 585
R12012 GND.n5539 GND.n5538 585
R12013 GND.n4323 GND.n4322 585
R12014 GND.n4324 GND.n4323 585
R12015 GND.n5467 GND.n5466 585
R12016 GND.n5467 GND.n4332 585
R12017 GND.n5469 GND.n5468 585
R12018 GND.n5468 GND.n4331 585
R12019 GND.n5470 GND.n4346 585
R12020 GND.n5455 GND.n4346 585
R12021 GND.n5472 GND.n5471 585
R12022 GND.n5473 GND.n5472 585
R12023 GND.n5465 GND.n4345 585
R12024 GND.n4345 GND.n4340 585
R12025 GND.n5464 GND.n5463 585
R12026 GND.n5463 GND.n5462 585
R12027 GND.n4348 GND.n4347 585
R12028 GND.n4355 GND.n4348 585
R12029 GND.n5437 GND.n5436 585
R12030 GND.n5438 GND.n5437 585
R12031 GND.n5435 GND.n4357 585
R12032 GND.n4357 GND.n4354 585
R12033 GND.n5434 GND.n5433 585
R12034 GND.n5433 GND.n5432 585
R12035 GND.n4359 GND.n4358 585
R12036 GND.n4372 GND.n4359 585
R12037 GND.n5409 GND.n4370 585
R12038 GND.n5421 GND.n4370 585
R12039 GND.n5410 GND.n4381 585
R12040 GND.n4381 GND.n4369 585
R12041 GND.n5412 GND.n5411 585
R12042 GND.n5413 GND.n5412 585
R12043 GND.n5408 GND.n4380 585
R12044 GND.n5404 GND.n4380 585
R12045 GND.n5407 GND.n5406 585
R12046 GND.n5406 GND.n5405 585
R12047 GND.n4383 GND.n4382 585
R12048 GND.n4389 GND.n4383 585
R12049 GND.n5397 GND.n5396 585
R12050 GND.n5398 GND.n5397 585
R12051 GND.n5395 GND.n4391 585
R12052 GND.n4391 GND.n4388 585
R12053 GND.n5394 GND.n5393 585
R12054 GND.n5393 GND.n5392 585
R12055 GND.n4393 GND.n4392 585
R12056 GND.n5283 GND.n4393 585
R12057 GND.n5373 GND.n5372 585
R12058 GND.n5374 GND.n5373 585
R12059 GND.n5371 GND.n4407 585
R12060 GND.n4407 GND.n4404 585
R12061 GND.n5370 GND.n5369 585
R12062 GND.n5369 GND.n5368 585
R12063 GND.n4409 GND.n4408 585
R12064 GND.n4410 GND.n4409 585
R12065 GND.n5307 GND.n5306 585
R12066 GND.n5307 GND.n4418 585
R12067 GND.n5309 GND.n5308 585
R12068 GND.n5308 GND.n4417 585
R12069 GND.n5310 GND.n4431 585
R12070 GND.n5295 GND.n4431 585
R12071 GND.n5312 GND.n5311 585
R12072 GND.n5313 GND.n5312 585
R12073 GND.n5305 GND.n4430 585
R12074 GND.n4430 GND.n4427 585
R12075 GND.n5304 GND.n5303 585
R12076 GND.n5303 GND.n5302 585
R12077 GND.n4433 GND.n4432 585
R12078 GND.n4440 GND.n4433 585
R12079 GND.n5275 GND.n5274 585
R12080 GND.n5276 GND.n5275 585
R12081 GND.n5273 GND.n4443 585
R12082 GND.n4443 GND.n4439 585
R12083 GND.n5272 GND.n5271 585
R12084 GND.n5271 GND.n5270 585
R12085 GND.n4445 GND.n4444 585
R12086 GND.n4459 GND.n4445 585
R12087 GND.n5247 GND.n4456 585
R12088 GND.n5259 GND.n4456 585
R12089 GND.n5248 GND.n4467 585
R12090 GND.n4467 GND.n4455 585
R12091 GND.n5250 GND.n5249 585
R12092 GND.n5251 GND.n5250 585
R12093 GND.n5246 GND.n4466 585
R12094 GND.n5242 GND.n4466 585
R12095 GND.n5245 GND.n5244 585
R12096 GND.n5244 GND.n5243 585
R12097 GND.n4469 GND.n4468 585
R12098 GND.n4475 GND.n4469 585
R12099 GND.n5235 GND.n5234 585
R12100 GND.n5236 GND.n5235 585
R12101 GND.n5233 GND.n4477 585
R12102 GND.n4477 GND.n4474 585
R12103 GND.n5232 GND.n5231 585
R12104 GND.n5231 GND.n5230 585
R12105 GND.n4479 GND.n4478 585
R12106 GND.n5133 GND.n4479 585
R12107 GND.n5211 GND.n5210 585
R12108 GND.n5212 GND.n5211 585
R12109 GND.n5209 GND.n4493 585
R12110 GND.n4493 GND.n4490 585
R12111 GND.n5208 GND.n5207 585
R12112 GND.n5207 GND.n5206 585
R12113 GND.n4495 GND.n4494 585
R12114 GND.n4496 GND.n4495 585
R12115 GND.n5146 GND.n4517 585
R12116 GND.n5146 GND.n5145 585
R12117 GND.n5148 GND.n5147 585
R12118 GND.n5147 GND.n4503 585
R12119 GND.n5149 GND.n4515 585
R12120 GND.n5128 GND.n4515 585
R12121 GND.n5151 GND.n5150 585
R12122 GND.n5152 GND.n5151 585
R12123 GND.n4516 GND.n4514 585
R12124 GND.n4514 GND.n4510 585
R12125 GND.n5122 GND.n5121 585
R12126 GND.n5123 GND.n5122 585
R12127 GND.n5120 GND.n4524 585
R12128 GND.n4530 GND.n4524 585
R12129 GND.n5119 GND.n5118 585
R12130 GND.n5118 GND.n5117 585
R12131 GND.n4526 GND.n4525 585
R12132 GND.n4527 GND.n4526 585
R12133 GND.n5106 GND.n5105 585
R12134 GND.n5107 GND.n5106 585
R12135 GND.n5104 GND.n4540 585
R12136 GND.n4540 GND.n4536 585
R12137 GND.n5103 GND.n5102 585
R12138 GND.n5102 GND.n5101 585
R12139 GND.n4542 GND.n4541 585
R12140 GND.n4543 GND.n4542 585
R12141 GND.n5088 GND.n5087 585
R12142 GND.n5089 GND.n5088 585
R12143 GND.n5086 GND.n4552 585
R12144 GND.n5082 GND.n4552 585
R12145 GND.n5085 GND.n5084 585
R12146 GND.n5084 GND.n5083 585
R12147 GND.n4554 GND.n4553 585
R12148 GND.n4560 GND.n4554 585
R12149 GND.n5075 GND.n5074 585
R12150 GND.n5076 GND.n5075 585
R12151 GND.n5073 GND.n4563 585
R12152 GND.n4563 GND.n4559 585
R12153 GND.n5072 GND.n5071 585
R12154 GND.n5071 GND.n5070 585
R12155 GND.n4565 GND.n4564 585
R12156 GND.n4578 GND.n4565 585
R12157 GND.n5048 GND.n5047 585
R12158 GND.n5049 GND.n5048 585
R12159 GND.n5046 GND.n4579 585
R12160 GND.n4579 GND.n4575 585
R12161 GND.n5045 GND.n5044 585
R12162 GND.n5044 GND.n5043 585
R12163 GND.n4581 GND.n4580 585
R12164 GND.n4582 GND.n4581 585
R12165 GND.n4982 GND.n4981 585
R12166 GND.n4982 GND.n4590 585
R12167 GND.n4984 GND.n4983 585
R12168 GND.n4983 GND.n4589 585
R12169 GND.n4985 GND.n4603 585
R12170 GND.n4970 GND.n4603 585
R12171 GND.n4987 GND.n4986 585
R12172 GND.n4988 GND.n4987 585
R12173 GND.n4980 GND.n4602 585
R12174 GND.n4602 GND.n4598 585
R12175 GND.n4979 GND.n4978 585
R12176 GND.n4978 GND.n4977 585
R12177 GND.n4605 GND.n4604 585
R12178 GND.n4611 GND.n4605 585
R12179 GND.n4952 GND.n4951 585
R12180 GND.n4953 GND.n4952 585
R12181 GND.n4950 GND.n4613 585
R12182 GND.n4620 GND.n4613 585
R12183 GND.n4949 GND.n4948 585
R12184 GND.n4948 GND.n4947 585
R12185 GND.n4615 GND.n4614 585
R12186 GND.n4630 GND.n4615 585
R12187 GND.n4924 GND.n4628 585
R12188 GND.n4936 GND.n4628 585
R12189 GND.n4925 GND.n4638 585
R12190 GND.n4638 GND.n4627 585
R12191 GND.n4927 GND.n4926 585
R12192 GND.n4928 GND.n4927 585
R12193 GND.n4923 GND.n4637 585
R12194 GND.n4919 GND.n4637 585
R12195 GND.n4922 GND.n4921 585
R12196 GND.n4921 GND.n4920 585
R12197 GND.n4640 GND.n4639 585
R12198 GND.n4647 GND.n4640 585
R12199 GND.n4912 GND.n4911 585
R12200 GND.n4913 GND.n4912 585
R12201 GND.n4910 GND.n4649 585
R12202 GND.n4649 GND.n4646 585
R12203 GND.n4909 GND.n4908 585
R12204 GND.n4908 GND.n4907 585
R12205 GND.n4651 GND.n4650 585
R12206 GND.n4839 GND.n4651 585
R12207 GND.n4854 GND.n4853 585
R12208 GND.n4855 GND.n4854 585
R12209 GND.n4852 GND.n4660 585
R12210 GND.n4660 GND.n3023 585
R12211 GND.n4851 GND.n4850 585
R12212 GND.n4850 GND.n3021 585
R12213 GND.n4849 GND.n4661 585
R12214 GND.n4849 GND.n4848 585
R12215 GND.n3008 GND.n3007 585
R12216 GND.n3012 GND.n3008 585
R12217 GND.n7562 GND.n7561 585
R12218 GND.n7561 GND.n7560 585
R12219 GND.n7563 GND.n3003 585
R12220 GND.n3009 GND.n3003 585
R12221 GND.n7565 GND.n7564 585
R12222 GND.n7566 GND.n7565 585
R12223 GND.n3006 GND.n3002 585
R12224 GND.n3002 GND.n1849 585
R12225 GND.n3005 GND.n3004 585
R12226 GND.n3004 GND.n1839 585
R12227 GND.n2988 GND.n2987 585
R12228 GND.n2991 GND.n2988 585
R12229 GND.n7576 GND.n7575 585
R12230 GND.n7575 GND.n7574 585
R12231 GND.n7577 GND.n2985 585
R12232 GND.n2989 GND.n2985 585
R12233 GND.n7579 GND.n7578 585
R12234 GND.n7580 GND.n7579 585
R12235 GND.n2986 GND.n2984 585
R12236 GND.n2984 GND.n2981 585
R12237 GND.n4819 GND.n4818 585
R12238 GND.n4820 GND.n4819 585
R12239 GND.n2970 GND.n2969 585
R12240 GND.n2973 GND.n2970 585
R12241 GND.n7590 GND.n7589 585
R12242 GND.n7589 GND.n7588 585
R12243 GND.n7591 GND.n2967 585
R12244 GND.n4812 GND.n2967 585
R12245 GND.n7593 GND.n7592 585
R12246 GND.n7594 GND.n7593 585
R12247 GND.n2968 GND.n2966 585
R12248 GND.n2966 GND.n2964 585
R12249 GND.n4721 GND.n4720 585
R12250 GND.n4724 GND.n4723 585
R12251 GND.n4725 GND.n4698 585
R12252 GND.n4698 GND.n2955 585
R12253 GND.n4727 GND.n4726 585
R12254 GND.n4729 GND.n4697 585
R12255 GND.n4732 GND.n4731 585
R12256 GND.n4733 GND.n4696 585
R12257 GND.n4735 GND.n4734 585
R12258 GND.n4737 GND.n4695 585
R12259 GND.n4740 GND.n4739 585
R12260 GND.n4741 GND.n4694 585
R12261 GND.n4743 GND.n4742 585
R12262 GND.n4745 GND.n4693 585
R12263 GND.n4748 GND.n4747 585
R12264 GND.n4749 GND.n4692 585
R12265 GND.n4751 GND.n4750 585
R12266 GND.n4753 GND.n4691 585
R12267 GND.n4756 GND.n4755 585
R12268 GND.n4758 GND.n4688 585
R12269 GND.n4760 GND.n4759 585
R12270 GND.n4762 GND.n4687 585
R12271 GND.n4763 GND.n1795 585
R12272 GND.n4767 GND.n4686 585
R12273 GND.n4770 GND.n4769 585
R12274 GND.n4771 GND.n4683 585
R12275 GND.n4774 GND.n4773 585
R12276 GND.n4776 GND.n4682 585
R12277 GND.n4779 GND.n4778 585
R12278 GND.n4780 GND.n4681 585
R12279 GND.n4782 GND.n4781 585
R12280 GND.n4784 GND.n4680 585
R12281 GND.n4787 GND.n4786 585
R12282 GND.n4788 GND.n4679 585
R12283 GND.n4790 GND.n4789 585
R12284 GND.n4792 GND.n4678 585
R12285 GND.n4795 GND.n4794 585
R12286 GND.n4796 GND.n4677 585
R12287 GND.n4798 GND.n4797 585
R12288 GND.n4800 GND.n4676 585
R12289 GND.n4803 GND.n4802 585
R12290 GND.n4804 GND.n4675 585
R12291 GND.n4806 GND.n4805 585
R12292 GND.n4808 GND.n4674 585
R12293 GND.n6143 GND.n6142 585
R12294 GND.n6145 GND.n6144 585
R12295 GND.n6147 GND.n6146 585
R12296 GND.n6149 GND.n6148 585
R12297 GND.n6151 GND.n6150 585
R12298 GND.n6153 GND.n6152 585
R12299 GND.n6155 GND.n6154 585
R12300 GND.n6157 GND.n6156 585
R12301 GND.n6159 GND.n6158 585
R12302 GND.n6161 GND.n6160 585
R12303 GND.n6163 GND.n6162 585
R12304 GND.n6165 GND.n6164 585
R12305 GND.n6167 GND.n6166 585
R12306 GND.n6169 GND.n6168 585
R12307 GND.n6171 GND.n6170 585
R12308 GND.n6173 GND.n6172 585
R12309 GND.n6175 GND.n6174 585
R12310 GND.n6177 GND.n6176 585
R12311 GND.n6179 GND.n6178 585
R12312 GND.n6181 GND.n6180 585
R12313 GND.n6182 GND.n6120 585
R12314 GND.n6260 GND.n6259 585
R12315 GND.n6123 GND.n6121 585
R12316 GND.n6218 GND.n6217 585
R12317 GND.n6220 GND.n6219 585
R12318 GND.n6223 GND.n6222 585
R12319 GND.n6225 GND.n6224 585
R12320 GND.n6227 GND.n6226 585
R12321 GND.n6229 GND.n6228 585
R12322 GND.n6231 GND.n6230 585
R12323 GND.n6233 GND.n6232 585
R12324 GND.n6235 GND.n6234 585
R12325 GND.n6237 GND.n6236 585
R12326 GND.n6239 GND.n6238 585
R12327 GND.n6241 GND.n6240 585
R12328 GND.n6243 GND.n6242 585
R12329 GND.n6245 GND.n6244 585
R12330 GND.n6247 GND.n6246 585
R12331 GND.n6249 GND.n6248 585
R12332 GND.n6251 GND.n6250 585
R12333 GND.n6253 GND.n6252 585
R12334 GND.n6254 GND.n6194 585
R12335 GND.n6256 GND.n6255 585
R12336 GND.n6257 GND.n6256 585
R12337 GND.n6141 GND.n6139 585
R12338 GND.n6141 GND.n6140 585
R12339 GND.n6138 GND.n3272 585
R12340 GND.n7309 GND.n3272 585
R12341 GND.n3264 GND.n3263 585
R12342 GND.n3271 GND.n3264 585
R12343 GND.n7317 GND.n7316 585
R12344 GND.n7316 GND.n7315 585
R12345 GND.n7318 GND.n3261 585
R12346 GND.n3261 GND.n3259 585
R12347 GND.n7320 GND.n7319 585
R12348 GND.n7321 GND.n7320 585
R12349 GND.n3262 GND.n3260 585
R12350 GND.n6376 GND.n3260 585
R12351 GND.n6380 GND.n6379 585
R12352 GND.n6379 GND.n6378 585
R12353 GND.n6381 GND.n3250 585
R12354 GND.n7328 GND.n3250 585
R12355 GND.n6383 GND.n6382 585
R12356 GND.n6382 GND.n3249 585
R12357 GND.n6384 GND.n3242 585
R12358 GND.n7334 GND.n3242 585
R12359 GND.n6386 GND.n6385 585
R12360 GND.n6385 GND.n3241 585
R12361 GND.n6387 GND.n3974 585
R12362 GND.n6400 GND.n3974 585
R12363 GND.n6389 GND.n6388 585
R12364 GND.n6388 GND.n3232 585
R12365 GND.n6390 GND.n3980 585
R12366 GND.n3980 GND.n3230 585
R12367 GND.n6392 GND.n6391 585
R12368 GND.n6393 GND.n6392 585
R12369 GND.n6372 GND.n3979 585
R12370 GND.n3984 GND.n3979 585
R12371 GND.n6371 GND.n6370 585
R12372 GND.n6370 GND.n6369 585
R12373 GND.n3982 GND.n3981 585
R12374 GND.n3983 GND.n3982 585
R12375 GND.n6054 GND.n3990 585
R12376 GND.n6362 GND.n3990 585
R12377 GND.n6057 GND.n6056 585
R12378 GND.n6056 GND.n6055 585
R12379 GND.n6058 GND.n4000 585
R12380 GND.n6348 GND.n4000 585
R12381 GND.n6060 GND.n6059 585
R12382 GND.n6059 GND.n3998 585
R12383 GND.n6061 GND.n4005 585
R12384 GND.n6342 GND.n4005 585
R12385 GND.n6062 GND.n6053 585
R12386 GND.n6053 GND.n4004 585
R12387 GND.n6064 GND.n6063 585
R12388 GND.n6064 GND.n4012 585
R12389 GND.n6065 GND.n6052 585
R12390 GND.n6065 GND.n4011 585
R12391 GND.n6068 GND.n6067 585
R12392 GND.n6067 GND.n6066 585
R12393 GND.n6069 GND.n4022 585
R12394 GND.n6084 GND.n4022 585
R12395 GND.n6070 GND.n4032 585
R12396 GND.n4032 GND.n4020 585
R12397 GND.n6072 GND.n6071 585
R12398 GND.n6073 GND.n6072 585
R12399 GND.n6051 GND.n4031 585
R12400 GND.n4031 GND.n4029 585
R12401 GND.n6050 GND.n6049 585
R12402 GND.n6049 GND.n6048 585
R12403 GND.n4034 GND.n4033 585
R12404 GND.n6041 GND.n4034 585
R12405 GND.n6040 GND.n6039 585
R12406 GND.n6042 GND.n6040 585
R12407 GND.n6038 GND.n4042 585
R12408 GND.n4046 GND.n4042 585
R12409 GND.n6037 GND.n6036 585
R12410 GND.n6036 GND.n6035 585
R12411 GND.n4044 GND.n4043 585
R12412 GND.n4045 GND.n4044 585
R12413 GND.n5930 GND.n4053 585
R12414 GND.n6029 GND.n4053 585
R12415 GND.n5932 GND.n5931 585
R12416 GND.n5931 GND.n4064 585
R12417 GND.n5933 GND.n4063 585
R12418 GND.n6008 GND.n4063 585
R12419 GND.n5935 GND.n5934 585
R12420 GND.n5934 GND.n4061 585
R12421 GND.n5936 GND.n4069 585
R12422 GND.n6002 GND.n4069 585
R12423 GND.n5937 GND.n5929 585
R12424 GND.n5929 GND.n4068 585
R12425 GND.n5939 GND.n5938 585
R12426 GND.n5939 GND.n4076 585
R12427 GND.n5940 GND.n5928 585
R12428 GND.n5940 GND.n4075 585
R12429 GND.n5943 GND.n5942 585
R12430 GND.n5942 GND.n5941 585
R12431 GND.n5944 GND.n4087 585
R12432 GND.n5959 GND.n4087 585
R12433 GND.n5945 GND.n4095 585
R12434 GND.n4095 GND.n4085 585
R12435 GND.n5947 GND.n5946 585
R12436 GND.n5948 GND.n5947 585
R12437 GND.n5927 GND.n4094 585
R12438 GND.n4098 GND.n4094 585
R12439 GND.n5926 GND.n5925 585
R12440 GND.n5925 GND.n5924 585
R12441 GND.n4097 GND.n4096 585
R12442 GND.n4107 GND.n4097 585
R12443 GND.n5903 GND.n4105 585
R12444 GND.n5918 GND.n4105 585
R12445 GND.n5904 GND.n4119 585
R12446 GND.n4119 GND.n4117 585
R12447 GND.n5906 GND.n5905 585
R12448 GND.n5907 GND.n5906 585
R12449 GND.n5902 GND.n4118 585
R12450 GND.n4118 GND.n4114 585
R12451 GND.n5901 GND.n5900 585
R12452 GND.n5900 GND.n5899 585
R12453 GND.n4121 GND.n4120 585
R12454 GND.n5890 GND.n4121 585
R12455 GND.n5889 GND.n5888 585
R12456 GND.n5891 GND.n5889 585
R12457 GND.n5887 GND.n4130 585
R12458 GND.n4134 GND.n4130 585
R12459 GND.n5886 GND.n5885 585
R12460 GND.n5885 GND.n5884 585
R12461 GND.n4132 GND.n4131 585
R12462 GND.n4133 GND.n4132 585
R12463 GND.n5846 GND.n4140 585
R12464 GND.n5878 GND.n4140 585
R12465 GND.n5848 GND.n5847 585
R12466 GND.n5847 GND.n4151 585
R12467 GND.n5849 GND.n4150 585
R12468 GND.n5860 GND.n4150 585
R12469 GND.n5851 GND.n5850 585
R12470 GND.n5852 GND.n5851 585
R12471 GND.n5845 GND.n4156 585
R12472 GND.n5854 GND.n4156 585
R12473 GND.n5844 GND.n5843 585
R12474 GND.n5843 GND.n4155 585
R12475 GND.n5842 GND.n4158 585
R12476 GND.n5842 GND.n5841 585
R12477 GND.n5831 GND.n4159 585
R12478 GND.n5834 GND.n4159 585
R12479 GND.n5833 GND.n5832 585
R12480 GND.n5835 GND.n5833 585
R12481 GND.n5830 GND.n4167 585
R12482 GND.n4171 GND.n4167 585
R12483 GND.n5829 GND.n5828 585
R12484 GND.n5828 GND.n5827 585
R12485 GND.n4169 GND.n4168 585
R12486 GND.n4170 GND.n4169 585
R12487 GND.n5656 GND.n4177 585
R12488 GND.n5821 GND.n4177 585
R12489 GND.n5658 GND.n5657 585
R12490 GND.n5657 GND.n4189 585
R12491 GND.n5659 GND.n4188 585
R12492 GND.n5800 GND.n4188 585
R12493 GND.n5661 GND.n5660 585
R12494 GND.n5660 GND.n4186 585
R12495 GND.n5662 GND.n4195 585
R12496 GND.n5794 GND.n4195 585
R12497 GND.n5663 GND.n5655 585
R12498 GND.n5655 GND.n4194 585
R12499 GND.n5665 GND.n5664 585
R12500 GND.n5665 GND.n4202 585
R12501 GND.n5666 GND.n5654 585
R12502 GND.n5666 GND.n4201 585
R12503 GND.n5668 GND.n5667 585
R12504 GND.n5667 GND.n4213 585
R12505 GND.n5669 GND.n4211 585
R12506 GND.n5719 GND.n4211 585
R12507 GND.n5671 GND.n5670 585
R12508 GND.n5670 GND.n4209 585
R12509 GND.n5672 GND.n4219 585
R12510 GND.n5708 GND.n4219 585
R12511 GND.n5673 GND.n4241 585
R12512 GND.n4241 GND.n4218 585
R12513 GND.n5675 GND.n5674 585
R12514 GND.n5677 GND.n5675 585
R12515 GND.n5653 GND.n4240 585
R12516 GND.n4240 GND.n4225 585
R12517 GND.n5652 GND.n5651 585
R12518 GND.n5651 GND.n5650 585
R12519 GND.n5649 GND.n4234 585
R12520 GND.n5684 GND.n4234 585
R12521 GND.n5648 GND.n5647 585
R12522 GND.n5647 GND.n4232 585
R12523 GND.n5646 GND.n4242 585
R12524 GND.n5646 GND.n5645 585
R12525 GND.n5613 GND.n4243 585
R12526 GND.n4250 GND.n4243 585
R12527 GND.n5614 GND.n4248 585
R12528 GND.n5639 GND.n4248 585
R12529 GND.n5617 GND.n5616 585
R12530 GND.n5616 GND.n5615 585
R12531 GND.n5618 GND.n4258 585
R12532 GND.n5628 GND.n4258 585
R12533 GND.n5619 GND.n4265 585
R12534 GND.n4265 GND.n4256 585
R12535 GND.n5621 GND.n5620 585
R12536 GND.n5622 GND.n5621 585
R12537 GND.n5612 GND.n4264 585
R12538 GND.n4269 GND.n4264 585
R12539 GND.n5611 GND.n5610 585
R12540 GND.n5610 GND.n5609 585
R12541 GND.n4267 GND.n4266 585
R12542 GND.n4268 GND.n4267 585
R12543 GND.n5588 GND.n4276 585
R12544 GND.n5603 GND.n4276 585
R12545 GND.n5589 GND.n4289 585
R12546 GND.n4289 GND.n4287 585
R12547 GND.n5591 GND.n5590 585
R12548 GND.n5592 GND.n5591 585
R12549 GND.n5587 GND.n4288 585
R12550 GND.n4288 GND.n4284 585
R12551 GND.n5586 GND.n5585 585
R12552 GND.n5585 GND.n5584 585
R12553 GND.n4291 GND.n4290 585
R12554 GND.n5575 GND.n4291 585
R12555 GND.n5574 GND.n5573 585
R12556 GND.n5576 GND.n5574 585
R12557 GND.n5572 GND.n4299 585
R12558 GND.n4303 GND.n4299 585
R12559 GND.n5571 GND.n5570 585
R12560 GND.n5570 GND.n5569 585
R12561 GND.n4301 GND.n4300 585
R12562 GND.n4302 GND.n4301 585
R12563 GND.n5444 GND.n4309 585
R12564 GND.n5563 GND.n4309 585
R12565 GND.n5446 GND.n5445 585
R12566 GND.n5445 GND.n4320 585
R12567 GND.n5447 GND.n4319 585
R12568 GND.n5544 GND.n4319 585
R12569 GND.n5449 GND.n5448 585
R12570 GND.n5448 GND.n4317 585
R12571 GND.n5450 GND.n4325 585
R12572 GND.n5538 GND.n4325 585
R12573 GND.n5451 GND.n5443 585
R12574 GND.n5443 GND.n4324 585
R12575 GND.n5453 GND.n5452 585
R12576 GND.n5453 GND.n4332 585
R12577 GND.n5454 GND.n5442 585
R12578 GND.n5454 GND.n4331 585
R12579 GND.n5457 GND.n5456 585
R12580 GND.n5456 GND.n5455 585
R12581 GND.n5458 GND.n4342 585
R12582 GND.n5473 GND.n4342 585
R12583 GND.n5459 GND.n4351 585
R12584 GND.n4351 GND.n4340 585
R12585 GND.n5461 GND.n5460 585
R12586 GND.n5462 GND.n5461 585
R12587 GND.n5441 GND.n4350 585
R12588 GND.n4355 GND.n4350 585
R12589 GND.n5440 GND.n5439 585
R12590 GND.n5439 GND.n5438 585
R12591 GND.n4353 GND.n4352 585
R12592 GND.n4354 GND.n4353 585
R12593 GND.n5417 GND.n4360 585
R12594 GND.n5432 GND.n4360 585
R12595 GND.n5418 GND.n4374 585
R12596 GND.n4374 GND.n4372 585
R12597 GND.n5420 GND.n5419 585
R12598 GND.n5421 GND.n5420 585
R12599 GND.n5416 GND.n4373 585
R12600 GND.n4373 GND.n4369 585
R12601 GND.n5415 GND.n5414 585
R12602 GND.n5414 GND.n5413 585
R12603 GND.n4376 GND.n4375 585
R12604 GND.n5404 GND.n4376 585
R12605 GND.n5403 GND.n5402 585
R12606 GND.n5405 GND.n5403 585
R12607 GND.n5401 GND.n4385 585
R12608 GND.n4389 GND.n4385 585
R12609 GND.n5400 GND.n5399 585
R12610 GND.n5399 GND.n5398 585
R12611 GND.n4387 GND.n4386 585
R12612 GND.n4388 GND.n4387 585
R12613 GND.n5282 GND.n4396 585
R12614 GND.n5392 GND.n4396 585
R12615 GND.n5285 GND.n5284 585
R12616 GND.n5284 GND.n5283 585
R12617 GND.n5286 GND.n4406 585
R12618 GND.n5374 GND.n4406 585
R12619 GND.n5288 GND.n5287 585
R12620 GND.n5287 GND.n4404 585
R12621 GND.n5289 GND.n4411 585
R12622 GND.n5368 GND.n4411 585
R12623 GND.n5290 GND.n5281 585
R12624 GND.n5281 GND.n4410 585
R12625 GND.n5292 GND.n5291 585
R12626 GND.n5292 GND.n4418 585
R12627 GND.n5293 GND.n5280 585
R12628 GND.n5293 GND.n4417 585
R12629 GND.n5297 GND.n5296 585
R12630 GND.n5296 GND.n5295 585
R12631 GND.n5298 GND.n4429 585
R12632 GND.n5313 GND.n4429 585
R12633 GND.n5299 GND.n4436 585
R12634 GND.n4436 GND.n4427 585
R12635 GND.n5301 GND.n5300 585
R12636 GND.n5302 GND.n5301 585
R12637 GND.n5279 GND.n4435 585
R12638 GND.n4440 GND.n4435 585
R12639 GND.n5278 GND.n5277 585
R12640 GND.n5277 GND.n5276 585
R12641 GND.n4438 GND.n4437 585
R12642 GND.n4439 GND.n4438 585
R12643 GND.n5255 GND.n4447 585
R12644 GND.n5270 GND.n4447 585
R12645 GND.n5256 GND.n4460 585
R12646 GND.n4460 GND.n4459 585
R12647 GND.n5258 GND.n5257 585
R12648 GND.n5259 GND.n5258 585
R12649 GND.n5254 GND.n4458 585
R12650 GND.n4458 GND.n4455 585
R12651 GND.n5253 GND.n5252 585
R12652 GND.n5252 GND.n5251 585
R12653 GND.n4462 GND.n4461 585
R12654 GND.n5242 GND.n4462 585
R12655 GND.n5241 GND.n5240 585
R12656 GND.n5243 GND.n5241 585
R12657 GND.n5239 GND.n4471 585
R12658 GND.n4475 GND.n4471 585
R12659 GND.n5238 GND.n5237 585
R12660 GND.n5237 GND.n5236 585
R12661 GND.n4473 GND.n4472 585
R12662 GND.n4474 GND.n4473 585
R12663 GND.n5132 GND.n4481 585
R12664 GND.n5230 GND.n4481 585
R12665 GND.n5135 GND.n5134 585
R12666 GND.n5134 GND.n5133 585
R12667 GND.n5136 GND.n4492 585
R12668 GND.n5212 GND.n4492 585
R12669 GND.n5138 GND.n5137 585
R12670 GND.n5137 GND.n4490 585
R12671 GND.n5139 GND.n4497 585
R12672 GND.n5206 GND.n4497 585
R12673 GND.n5140 GND.n4519 585
R12674 GND.n4519 GND.n4496 585
R12675 GND.n5142 GND.n5141 585
R12676 GND.n5145 GND.n5142 585
R12677 GND.n5131 GND.n4518 585
R12678 GND.n4518 GND.n4503 585
R12679 GND.n5130 GND.n5129 585
R12680 GND.n5129 GND.n5128 585
R12681 GND.n5127 GND.n4512 585
R12682 GND.n5152 GND.n4512 585
R12683 GND.n5126 GND.n5125 585
R12684 GND.n5125 GND.n4510 585
R12685 GND.n5124 GND.n4520 585
R12686 GND.n5124 GND.n5123 585
R12687 GND.n5093 GND.n4521 585
R12688 GND.n4530 GND.n4521 585
R12689 GND.n5094 GND.n4528 585
R12690 GND.n5117 GND.n4528 585
R12691 GND.n5096 GND.n5095 585
R12692 GND.n5095 GND.n4527 585
R12693 GND.n5097 GND.n4538 585
R12694 GND.n5107 GND.n4538 585
R12695 GND.n5098 GND.n4547 585
R12696 GND.n4547 GND.n4536 585
R12697 GND.n5100 GND.n5099 585
R12698 GND.n5101 GND.n5100 585
R12699 GND.n5092 GND.n4546 585
R12700 GND.n4546 GND.n4543 585
R12701 GND.n5091 GND.n5090 585
R12702 GND.n5090 GND.n5089 585
R12703 GND.n4549 GND.n4548 585
R12704 GND.n5082 GND.n4549 585
R12705 GND.n5081 GND.n5080 585
R12706 GND.n5083 GND.n5081 585
R12707 GND.n5079 GND.n4556 585
R12708 GND.n4560 GND.n4556 585
R12709 GND.n5078 GND.n5077 585
R12710 GND.n5077 GND.n5076 585
R12711 GND.n4558 GND.n4557 585
R12712 GND.n4559 GND.n4558 585
R12713 GND.n4959 GND.n4567 585
R12714 GND.n5070 GND.n4567 585
R12715 GND.n4961 GND.n4960 585
R12716 GND.n4960 GND.n4578 585
R12717 GND.n4962 GND.n4577 585
R12718 GND.n5049 GND.n4577 585
R12719 GND.n4964 GND.n4963 585
R12720 GND.n4963 GND.n4575 585
R12721 GND.n4965 GND.n4583 585
R12722 GND.n5043 GND.n4583 585
R12723 GND.n4966 GND.n4958 585
R12724 GND.n4958 GND.n4582 585
R12725 GND.n4968 GND.n4967 585
R12726 GND.n4968 GND.n4590 585
R12727 GND.n4969 GND.n4957 585
R12728 GND.n4969 GND.n4589 585
R12729 GND.n4972 GND.n4971 585
R12730 GND.n4971 GND.n4970 585
R12731 GND.n4973 GND.n4600 585
R12732 GND.n4988 GND.n4600 585
R12733 GND.n4974 GND.n4608 585
R12734 GND.n4608 GND.n4598 585
R12735 GND.n4976 GND.n4975 585
R12736 GND.n4977 GND.n4976 585
R12737 GND.n4956 GND.n4607 585
R12738 GND.n4611 GND.n4607 585
R12739 GND.n4955 GND.n4954 585
R12740 GND.n4954 GND.n4953 585
R12741 GND.n4610 GND.n4609 585
R12742 GND.n4620 GND.n4610 585
R12743 GND.n4932 GND.n4618 585
R12744 GND.n4947 GND.n4618 585
R12745 GND.n4933 GND.n4632 585
R12746 GND.n4632 GND.n4630 585
R12747 GND.n4935 GND.n4934 585
R12748 GND.n4936 GND.n4935 585
R12749 GND.n4931 GND.n4631 585
R12750 GND.n4631 GND.n4627 585
R12751 GND.n4930 GND.n4929 585
R12752 GND.n4929 GND.n4928 585
R12753 GND.n4634 GND.n4633 585
R12754 GND.n4919 GND.n4634 585
R12755 GND.n4918 GND.n4917 585
R12756 GND.n4920 GND.n4918 585
R12757 GND.n4916 GND.n4643 585
R12758 GND.n4647 GND.n4643 585
R12759 GND.n4915 GND.n4914 585
R12760 GND.n4914 GND.n4913 585
R12761 GND.n4645 GND.n4644 585
R12762 GND.n4646 GND.n4645 585
R12763 GND.n4838 GND.n4653 585
R12764 GND.n4907 GND.n4653 585
R12765 GND.n4841 GND.n4840 585
R12766 GND.n4840 GND.n4839 585
R12767 GND.n4842 GND.n4659 585
R12768 GND.n4855 GND.n4659 585
R12769 GND.n4844 GND.n4843 585
R12770 GND.n4843 GND.n3023 585
R12771 GND.n4845 GND.n4671 585
R12772 GND.n4671 GND.n3021 585
R12773 GND.n4847 GND.n4846 585
R12774 GND.n4848 GND.n4847 585
R12775 GND.n4837 GND.n4670 585
R12776 GND.n4670 GND.n3012 585
R12777 GND.n4836 GND.n3010 585
R12778 GND.n7560 GND.n3010 585
R12779 GND.n4835 GND.n4834 585
R12780 GND.n4834 GND.n3009 585
R12781 GND.n4833 GND.n3000 585
R12782 GND.n7566 GND.n3000 585
R12783 GND.n4832 GND.n4831 585
R12784 GND.n4831 GND.n1849 585
R12785 GND.n4830 GND.n4672 585
R12786 GND.n4830 GND.n1839 585
R12787 GND.n4829 GND.n4828 585
R12788 GND.n4829 GND.n2991 585
R12789 GND.n4827 GND.n2990 585
R12790 GND.n7574 GND.n2990 585
R12791 GND.n4826 GND.n4825 585
R12792 GND.n4825 GND.n2989 585
R12793 GND.n4824 GND.n2982 585
R12794 GND.n7580 GND.n2982 585
R12795 GND.n4823 GND.n4822 585
R12796 GND.n4822 GND.n2981 585
R12797 GND.n4821 GND.n4673 585
R12798 GND.n4821 GND.n4820 585
R12799 GND.n4817 GND.n4816 585
R12800 GND.n4817 GND.n2973 585
R12801 GND.n4815 GND.n2972 585
R12802 GND.n7588 GND.n2972 585
R12803 GND.n4814 GND.n4813 585
R12804 GND.n4813 GND.n4812 585
R12805 GND.n4811 GND.n2965 585
R12806 GND.n7594 GND.n2965 585
R12807 GND.n4810 GND.n4809 585
R12808 GND.n4809 GND.n2964 585
R12809 GND.n8177 GND.n8176 585
R12810 GND.n8178 GND.n8177 585
R12811 GND.n9458 GND.n617 585
R12812 GND.n617 GND.n616 585
R12813 GND.n9462 GND.n9461 585
R12814 GND.n9463 GND.n9462 585
R12815 GND.n615 GND.n614 585
R12816 GND.n9464 GND.n615 585
R12817 GND.n9467 GND.n9466 585
R12818 GND.n9466 GND.n9465 585
R12819 GND.n9468 GND.n609 585
R12820 GND.n609 GND.n608 585
R12821 GND.n9470 GND.n9469 585
R12822 GND.n9471 GND.n9470 585
R12823 GND.n607 GND.n606 585
R12824 GND.n9472 GND.n607 585
R12825 GND.n9475 GND.n9474 585
R12826 GND.n9474 GND.n9473 585
R12827 GND.n9476 GND.n601 585
R12828 GND.n601 GND.n600 585
R12829 GND.n9478 GND.n9477 585
R12830 GND.n9479 GND.n9478 585
R12831 GND.n599 GND.n598 585
R12832 GND.n9480 GND.n599 585
R12833 GND.n9483 GND.n9482 585
R12834 GND.n9482 GND.n9481 585
R12835 GND.n9484 GND.n593 585
R12836 GND.n593 GND.n544 585
R12837 GND.n9486 GND.n9485 585
R12838 GND.n9486 GND.n519 585
R12839 GND.n9487 GND.n592 585
R12840 GND.n9487 GND.n478 585
R12841 GND.n9489 GND.n9488 585
R12842 GND.n9488 GND.n476 585
R12843 GND.n9490 GND.n587 585
R12844 GND.n587 GND.n551 585
R12845 GND.n9492 GND.n9491 585
R12846 GND.n9492 GND.n558 585
R12847 GND.n9493 GND.n586 585
R12848 GND.n9493 GND.n557 585
R12849 GND.n9495 GND.n9494 585
R12850 GND.n9494 GND.n570 585
R12851 GND.n9496 GND.n581 585
R12852 GND.n581 GND.n567 585
R12853 GND.n9498 GND.n9497 585
R12854 GND.t114 GND.n9498 585
R12855 GND.n582 GND.n580 585
R12856 GND.n3571 GND.n580 585
R12857 GND.n7078 GND.n7077 585
R12858 GND.n7078 GND.n3569 585
R12859 GND.n7080 GND.n7079 585
R12860 GND.n7079 GND.n3581 585
R12861 GND.n7081 GND.n3586 585
R12862 GND.n3586 GND.n3578 585
R12863 GND.n7083 GND.n7082 585
R12864 GND.n7084 GND.n7083 585
R12865 GND.n3587 GND.n3585 585
R12866 GND.n3593 GND.n3585 585
R12867 GND.n7069 GND.n7068 585
R12868 GND.n7068 GND.n7067 585
R12869 GND.n3590 GND.n3589 585
R12870 GND.n3602 GND.n3590 585
R12871 GND.n7046 GND.n3607 585
R12872 GND.n3607 GND.n3601 585
R12873 GND.n7048 GND.n7047 585
R12874 GND.n7049 GND.n7048 585
R12875 GND.n3608 GND.n3606 585
R12876 GND.n3613 GND.n3606 585
R12877 GND.n7041 GND.n7040 585
R12878 GND.n7040 GND.n7039 585
R12879 GND.n3611 GND.n3610 585
R12880 GND.n3624 GND.n3611 585
R12881 GND.n7019 GND.n3629 585
R12882 GND.n3629 GND.n3622 585
R12883 GND.n7021 GND.n7020 585
R12884 GND.n7022 GND.n7021 585
R12885 GND.n3630 GND.n3628 585
R12886 GND.n3636 GND.n3628 585
R12887 GND.n7014 GND.n7013 585
R12888 GND.n7013 GND.n7012 585
R12889 GND.n3633 GND.n3632 585
R12890 GND.n3646 GND.n3633 585
R12891 GND.n6993 GND.n3651 585
R12892 GND.n3651 GND.n3644 585
R12893 GND.n6995 GND.n6994 585
R12894 GND.n6996 GND.n6995 585
R12895 GND.n3652 GND.n3650 585
R12896 GND.n3659 GND.n3650 585
R12897 GND.n6988 GND.n6987 585
R12898 GND.n6987 GND.n6986 585
R12899 GND.n3655 GND.n3654 585
R12900 GND.n3668 GND.n3655 585
R12901 GND.n6966 GND.n3673 585
R12902 GND.n3673 GND.n3667 585
R12903 GND.n6968 GND.n6967 585
R12904 GND.n6969 GND.n6968 585
R12905 GND.n3674 GND.n3672 585
R12906 GND.n3679 GND.n3672 585
R12907 GND.n6961 GND.n6960 585
R12908 GND.n6960 GND.n6959 585
R12909 GND.n3677 GND.n3676 585
R12910 GND.n3688 GND.n3677 585
R12911 GND.n6937 GND.n3693 585
R12912 GND.n3693 GND.n3687 585
R12913 GND.n6939 GND.n6938 585
R12914 GND.n6940 GND.n6939 585
R12915 GND.n3694 GND.n3692 585
R12916 GND.n3699 GND.n3692 585
R12917 GND.n6932 GND.n6931 585
R12918 GND.n6931 GND.n6930 585
R12919 GND.n3697 GND.n3696 585
R12920 GND.n3710 GND.n3697 585
R12921 GND.n6910 GND.n3715 585
R12922 GND.n3715 GND.n3708 585
R12923 GND.n6912 GND.n6911 585
R12924 GND.n6913 GND.n6912 585
R12925 GND.n3716 GND.n3714 585
R12926 GND.n3722 GND.n3714 585
R12927 GND.n6905 GND.n6904 585
R12928 GND.n6904 GND.n6903 585
R12929 GND.n3719 GND.n3718 585
R12930 GND.n3732 GND.n3719 585
R12931 GND.n6884 GND.n3737 585
R12932 GND.n3737 GND.n3730 585
R12933 GND.n6886 GND.n6885 585
R12934 GND.n6887 GND.n6886 585
R12935 GND.n3738 GND.n3736 585
R12936 GND.n6833 GND.n3736 585
R12937 GND.n6847 GND.n6846 585
R12938 GND.n6848 GND.n6847 585
R12939 GND.n6845 GND.n6844 585
R12940 GND.n6844 GND.n6827 585
R12941 GND.n6843 GND.n6842 585
R12942 GND.n6843 GND.n6826 585
R12943 GND.n6841 GND.n6816 585
R12944 GND.n6818 GND.n6816 585
R12945 GND.n6863 GND.n6862 585
R12946 GND.n6862 GND.n6861 585
R12947 GND.n6865 GND.n6864 585
R12948 GND.n6866 GND.n6865 585
R12949 GND.n6815 GND.n6814 585
R12950 GND.n6815 GND.n3761 585
R12951 GND.n6813 GND.n6812 585
R12952 GND.n6812 GND.n3759 585
R12953 GND.n3749 GND.n3747 585
R12954 GND.n3752 GND.n3749 585
R12955 GND.n6880 GND.n6879 585
R12956 GND.n6879 GND.n6878 585
R12957 GND.n3748 GND.n3746 585
R12958 GND.n3778 GND.n3748 585
R12959 GND.n6516 GND.n6515 585
R12960 GND.n6515 GND.n3775 585
R12961 GND.n6517 GND.n6510 585
R12962 GND.n6510 GND.n3773 585
R12963 GND.n6519 GND.n6518 585
R12964 GND.n6519 GND.n3790 585
R12965 GND.n6520 GND.n6509 585
R12966 GND.n6520 GND.n3788 585
R12967 GND.n6522 GND.n6521 585
R12968 GND.n6521 GND.n3792 585
R12969 GND.n6523 GND.n6504 585
R12970 GND.n6504 GND.n3800 585
R12971 GND.n6525 GND.n6524 585
R12972 GND.n6525 GND.n3799 585
R12973 GND.n6526 GND.n6503 585
R12974 GND.n6526 GND.n3812 585
R12975 GND.n6528 GND.n6527 585
R12976 GND.n6527 GND.n3810 585
R12977 GND.n6529 GND.n6498 585
R12978 GND.n6498 GND.n3814 585
R12979 GND.n6531 GND.n6530 585
R12980 GND.n6531 GND.n3823 585
R12981 GND.n6532 GND.n6497 585
R12982 GND.n6532 GND.n3822 585
R12983 GND.n6534 GND.n6533 585
R12984 GND.n6533 GND.n3836 585
R12985 GND.n6535 GND.n6492 585
R12986 GND.n6492 GND.n3833 585
R12987 GND.n6537 GND.n6536 585
R12988 GND.n6537 GND.n3839 585
R12989 GND.n6538 GND.n6491 585
R12990 GND.n6538 GND.n3847 585
R12991 GND.n6540 GND.n6539 585
R12992 GND.n6539 GND.n3846 585
R12993 GND.n6541 GND.n6486 585
R12994 GND.n6486 GND.n3858 585
R12995 GND.n6543 GND.n6542 585
R12996 GND.n6543 GND.n3856 585
R12997 GND.n6544 GND.n6485 585
R12998 GND.n6544 GND.n3861 585
R12999 GND.n6546 GND.n6545 585
R13000 GND.n6545 GND.n3870 585
R13001 GND.n6547 GND.n6480 585
R13002 GND.n6480 GND.n3868 585
R13003 GND.n6549 GND.n6548 585
R13004 GND.n6549 GND.n3881 585
R13005 GND.n6550 GND.n6479 585
R13006 GND.n6550 GND.n3879 585
R13007 GND.n6552 GND.n6551 585
R13008 GND.n6551 GND.n3883 585
R13009 GND.n6553 GND.n6474 585
R13010 GND.n6474 GND.n3891 585
R13011 GND.n6555 GND.n6554 585
R13012 GND.n6555 GND.n3890 585
R13013 GND.n6556 GND.n6473 585
R13014 GND.n6556 GND.n3903 585
R13015 GND.n6558 GND.n6557 585
R13016 GND.n6557 GND.n3901 585
R13017 GND.n6559 GND.n6468 585
R13018 GND.n6468 GND.n3905 585
R13019 GND.n6561 GND.n6560 585
R13020 GND.n6561 GND.n3914 585
R13021 GND.n6562 GND.n6467 585
R13022 GND.n6562 GND.n3913 585
R13023 GND.n6564 GND.n6563 585
R13024 GND.n6563 GND.n3927 585
R13025 GND.n6565 GND.n6462 585
R13026 GND.n6462 GND.n3924 585
R13027 GND.n6567 GND.n6566 585
R13028 GND.n6567 GND.n3930 585
R13029 GND.n6568 GND.n6461 585
R13030 GND.n6568 GND.n3938 585
R13031 GND.n6570 GND.n6569 585
R13032 GND.n6569 GND.n3937 585
R13033 GND.n6571 GND.n6456 585
R13034 GND.n6456 GND.n3949 585
R13035 GND.n6573 GND.n6572 585
R13036 GND.n6573 GND.n3947 585
R13037 GND.n6574 GND.n6455 585
R13038 GND.n6574 GND.t91 585
R13039 GND.n6576 GND.n6575 585
R13040 GND.n6575 GND.n3960 585
R13041 GND.n6577 GND.n6439 585
R13042 GND.n6439 GND.n3958 585
R13043 GND.n6579 GND.n6578 585
R13044 GND.n6580 GND.n6579 585
R13045 GND.n6440 GND.n6438 585
R13046 GND.n6438 GND.n3369 585
R13047 GND.n6449 GND.n6448 585
R13048 GND.n6448 GND.n3366 585
R13049 GND.n6447 GND.n6442 585
R13050 GND.n6447 GND.n3358 585
R13051 GND.n6446 GND.n6445 585
R13052 GND.n6446 GND.n3356 585
R13053 GND.n3291 GND.n3290 585
R13054 GND.n3312 GND.n3291 585
R13055 GND.n7296 GND.n7295 585
R13056 GND.n7295 GND.n7294 585
R13057 GND.n7297 GND.n3285 585
R13058 GND.n3285 GND.n3284 585
R13059 GND.n7299 GND.n7298 585
R13060 GND.n7300 GND.n7299 585
R13061 GND.n3283 GND.n3282 585
R13062 GND.n7301 GND.n3283 585
R13063 GND.n7304 GND.n7303 585
R13064 GND.n7303 GND.n7302 585
R13065 GND.n7305 GND.n3275 585
R13066 GND.n6124 GND.n3275 585
R13067 GND.n7307 GND.n7306 585
R13068 GND.n7308 GND.n7307 585
R13069 GND.n3276 GND.n3274 585
R13070 GND.n3274 GND.n3273 585
R13071 GND.n3257 GND.n3256 585
R13072 GND.n3265 GND.n3257 585
R13073 GND.n7323 GND.n7322 585
R13074 GND.n7322 GND.n7321 585
R13075 GND.n7324 GND.n3251 585
R13076 GND.n6377 GND.n3251 585
R13077 GND.n7326 GND.n7325 585
R13078 GND.n7327 GND.n7326 585
R13079 GND.n3240 GND.n3239 585
R13080 GND.n3243 GND.n3240 585
R13081 GND.n7337 GND.n7336 585
R13082 GND.n7336 GND.n7335 585
R13083 GND.n7338 GND.n3234 585
R13084 GND.n3973 GND.n3234 585
R13085 GND.n7340 GND.n7339 585
R13086 GND.n7341 GND.n7340 585
R13087 GND.n3235 GND.n3233 585
R13088 GND.n3978 GND.n3233 585
R13089 GND.n6358 GND.n3993 585
R13090 GND.n3993 GND.n3985 585
R13091 GND.n6360 GND.n6359 585
R13092 GND.n6361 GND.n6360 585
R13093 GND.n3994 GND.n3992 585
R13094 GND.n3992 GND.n3989 585
R13095 GND.n6352 GND.n6351 585
R13096 GND.n6351 GND.n6350 585
R13097 GND.n3997 GND.n3996 585
R13098 GND.n6341 GND.n3997 585
R13099 GND.n6092 GND.n4015 585
R13100 GND.n4015 GND.n4014 585
R13101 GND.n6094 GND.n6093 585
R13102 GND.n6095 GND.n6094 585
R13103 GND.n4016 GND.n4013 585
R13104 GND.n4024 GND.n4013 585
R13105 GND.n6087 GND.n6086 585
R13106 GND.n6086 GND.n6085 585
R13107 GND.n4019 GND.n4018 585
R13108 GND.n6073 GND.n4019 585
R13109 GND.n6021 GND.n6020 585
R13110 GND.n6021 GND.n4037 585
R13111 GND.n6022 GND.n6017 585
R13112 GND.n6022 GND.n4036 585
R13113 GND.n6024 GND.n6023 585
R13114 GND.n6023 GND.n4041 585
R13115 GND.n6025 GND.n4056 585
R13116 GND.n4056 GND.n4047 585
R13117 GND.n6027 GND.n6026 585
R13118 GND.n6028 GND.n6027 585
R13119 GND.n4057 GND.n4055 585
R13120 GND.n4055 GND.n4052 585
R13121 GND.n6011 GND.n6010 585
R13122 GND.n6010 GND.n6009 585
R13123 GND.n4060 GND.n4059 585
R13124 GND.n6001 GND.n4060 585
R13125 GND.n5967 GND.n4080 585
R13126 GND.n4080 GND.n4079 585
R13127 GND.n5969 GND.n5968 585
R13128 GND.n5970 GND.n5969 585
R13129 GND.n4081 GND.n4078 585
R13130 GND.n4088 GND.n4078 585
R13131 GND.n5962 GND.n5961 585
R13132 GND.n5961 GND.n5960 585
R13133 GND.n4084 GND.n4083 585
R13134 GND.n4093 GND.n4084 585
R13135 GND.n5914 GND.n4109 585
R13136 GND.n4109 GND.n4100 585
R13137 GND.n5916 GND.n5915 585
R13138 GND.n5917 GND.n5916 585
R13139 GND.n4110 GND.n4108 585
R13140 GND.n4108 GND.n4104 585
R13141 GND.n5909 GND.n5908 585
R13142 GND.n5908 GND.n5907 585
R13143 GND.n4113 GND.n4112 585
R13144 GND.n4124 GND.n4113 585
R13145 GND.n5871 GND.n5870 585
R13146 GND.n5871 GND.n4122 585
R13147 GND.n5873 GND.n5872 585
R13148 GND.n5872 GND.n4129 585
R13149 GND.n5874 GND.n4144 585
R13150 GND.n4144 GND.n4135 585
R13151 GND.n5876 GND.n5875 585
R13152 GND.n5877 GND.n5876 585
R13153 GND.n4145 GND.n4143 585
R13154 GND.n4143 GND.n4139 585
R13155 GND.n5863 GND.n5862 585
R13156 GND.n5862 GND.n5861 585
R13157 GND.n4148 GND.n4147 585
R13158 GND.n5853 GND.n4148 585
R13159 GND.n5813 GND.n5812 585
R13160 GND.n5813 GND.n4162 585
R13161 GND.n5814 GND.n5809 585
R13162 GND.n5814 GND.n4160 585
R13163 GND.n5816 GND.n5815 585
R13164 GND.n5815 GND.n4166 585
R13165 GND.n5817 GND.n4181 585
R13166 GND.n4181 GND.n4172 585
R13167 GND.n5819 GND.n5818 585
R13168 GND.n5820 GND.n5819 585
R13169 GND.n4182 GND.n4180 585
R13170 GND.n4180 GND.n4176 585
R13171 GND.n5803 GND.n5802 585
R13172 GND.n5802 GND.n5801 585
R13173 GND.n4185 GND.n4184 585
R13174 GND.n5793 GND.n4185 585
R13175 GND.n5727 GND.n4204 585
R13176 GND.n4204 GND.n4194 585
R13177 GND.n5729 GND.n5728 585
R13178 GND.n5730 GND.n5729 585
R13179 GND.n4205 GND.n4203 585
R13180 GND.n4212 GND.n4203 585
R13181 GND.n5722 GND.n5721 585
R13182 GND.n5721 GND.n5720 585
R13183 GND.n4208 GND.n4207 585
R13184 GND.n5707 GND.n4208 585
R13185 GND.n5693 GND.n4227 585
R13186 GND.n5676 GND.n4227 585
R13187 GND.n5695 GND.n5694 585
R13188 GND.n5696 GND.n5695 585
R13189 GND.n4228 GND.n4226 585
R13190 GND.n4235 GND.n4226 585
R13191 GND.n5688 GND.n5687 585
R13192 GND.n5687 GND.n5686 585
R13193 GND.n4231 GND.n4230 585
R13194 GND.n4244 GND.n4231 585
R13195 GND.n5637 GND.n5636 585
R13196 GND.n5638 GND.n5637 585
R13197 GND.n4252 GND.n4251 585
R13198 GND.n4259 GND.n4251 585
R13199 GND.n5632 GND.n5631 585
R13200 GND.n5631 GND.n5630 585
R13201 GND.n4255 GND.n4254 585
R13202 GND.n4263 GND.n4255 585
R13203 GND.n5599 GND.n4279 585
R13204 GND.n4279 GND.n4270 585
R13205 GND.n5601 GND.n5600 585
R13206 GND.n5602 GND.n5601 585
R13207 GND.n4280 GND.n4278 585
R13208 GND.n4278 GND.n4275 585
R13209 GND.n5594 GND.n5593 585
R13210 GND.n5593 GND.n5592 585
R13211 GND.n4283 GND.n4282 585
R13212 GND.n5495 GND.n4283 585
R13213 GND.n5556 GND.n5555 585
R13214 GND.n5556 GND.n4292 585
R13215 GND.n5558 GND.n5557 585
R13216 GND.n5557 GND.n4298 585
R13217 GND.n5559 GND.n4312 585
R13218 GND.n4312 GND.n4304 585
R13219 GND.n5561 GND.n5560 585
R13220 GND.n5562 GND.n5561 585
R13221 GND.n4313 GND.n4311 585
R13222 GND.n4311 GND.n4308 585
R13223 GND.n5548 GND.n5547 585
R13224 GND.n5547 GND.n5546 585
R13225 GND.n4316 GND.n4315 585
R13226 GND.n5537 GND.n4316 585
R13227 GND.n5481 GND.n4335 585
R13228 GND.n4335 GND.n4334 585
R13229 GND.n5483 GND.n5482 585
R13230 GND.n5484 GND.n5483 585
R13231 GND.n4336 GND.n4333 585
R13232 GND.n4344 GND.n4333 585
R13233 GND.n5476 GND.n5475 585
R13234 GND.n5475 GND.n5474 585
R13235 GND.n4339 GND.n4338 585
R13236 GND.n4349 GND.n4339 585
R13237 GND.n5428 GND.n4364 585
R13238 GND.n4364 GND.n4356 585
R13239 GND.n5430 GND.n5429 585
R13240 GND.n5431 GND.n5430 585
R13241 GND.n4365 GND.n4363 585
R13242 GND.n5351 GND.n4363 585
R13243 GND.n5423 GND.n5422 585
R13244 GND.n5422 GND.n5421 585
R13245 GND.n4368 GND.n4367 585
R13246 GND.n4379 GND.n4368 585
R13247 GND.n5385 GND.n5384 585
R13248 GND.n5385 GND.n4378 585
R13249 GND.n5387 GND.n5386 585
R13250 GND.n5386 GND.n4384 585
R13251 GND.n5388 GND.n4399 585
R13252 GND.n4399 GND.n4390 585
R13253 GND.n5390 GND.n5389 585
R13254 GND.n5391 GND.n5390 585
R13255 GND.n4400 GND.n4398 585
R13256 GND.n4398 GND.n4395 585
R13257 GND.n5377 GND.n5376 585
R13258 GND.n5376 GND.n5375 585
R13259 GND.n4403 GND.n4402 585
R13260 GND.n5367 GND.n4403 585
R13261 GND.n5321 GND.n4422 585
R13262 GND.n4422 GND.n4421 585
R13263 GND.n5323 GND.n5322 585
R13264 GND.n5324 GND.n5323 585
R13265 GND.n4423 GND.n4420 585
R13266 GND.n5294 GND.n4420 585
R13267 GND.n5316 GND.n5315 585
R13268 GND.n5315 GND.n5314 585
R13269 GND.n4426 GND.n4425 585
R13270 GND.n4434 GND.n4426 585
R13271 GND.n5266 GND.n4450 585
R13272 GND.n4450 GND.n4442 585
R13273 GND.n5268 GND.n5267 585
R13274 GND.n5269 GND.n5268 585
R13275 GND.n4451 GND.n4449 585
R13276 GND.n4449 GND.n4446 585
R13277 GND.n5261 GND.n5260 585
R13278 GND.n5260 GND.n5259 585
R13279 GND.n4454 GND.n4453 585
R13280 GND.n4465 GND.n4454 585
R13281 GND.n5223 GND.n5222 585
R13282 GND.n5223 GND.n4463 585
R13283 GND.n5225 GND.n5224 585
R13284 GND.n5224 GND.n4470 585
R13285 GND.n5226 GND.n4485 585
R13286 GND.n4485 GND.n4476 585
R13287 GND.n5228 GND.n5227 585
R13288 GND.n5229 GND.n5228 585
R13289 GND.n4486 GND.n4484 585
R13290 GND.n4484 GND.n4480 585
R13291 GND.n5215 GND.n5214 585
R13292 GND.n5214 GND.n5213 585
R13293 GND.n4489 GND.n4488 585
R13294 GND.n5205 GND.n4489 585
R13295 GND.n5160 GND.n4505 585
R13296 GND.n5144 GND.n4505 585
R13297 GND.n5162 GND.n5161 585
R13298 GND.n5163 GND.n5162 585
R13299 GND.n4506 GND.n4504 585
R13300 GND.n4513 GND.n4504 585
R13301 GND.n5155 GND.n5154 585
R13302 GND.n5154 GND.n5153 585
R13303 GND.n4509 GND.n4508 585
R13304 GND.n4523 GND.n4509 585
R13305 GND.n5115 GND.n5114 585
R13306 GND.n5116 GND.n5115 585
R13307 GND.n4532 GND.n4531 585
R13308 GND.n4539 GND.n4531 585
R13309 GND.n5110 GND.n5109 585
R13310 GND.n5109 GND.n5108 585
R13311 GND.n4535 GND.n4534 585
R13312 GND.n5101 GND.n4535 585
R13313 GND.n5062 GND.n5061 585
R13314 GND.n5062 GND.n4551 585
R13315 GND.n5063 GND.n5058 585
R13316 GND.n5063 GND.n4550 585
R13317 GND.n5065 GND.n5064 585
R13318 GND.n5064 GND.n4555 585
R13319 GND.n5066 GND.n4570 585
R13320 GND.n4570 GND.n4562 585
R13321 GND.n5068 GND.n5067 585
R13322 GND.n5069 GND.n5068 585
R13323 GND.n4571 GND.n4569 585
R13324 GND.n4569 GND.n4566 585
R13325 GND.n5052 GND.n5051 585
R13326 GND.n5051 GND.n5050 585
R13327 GND.n4574 GND.n4573 585
R13328 GND.n5042 GND.n4574 585
R13329 GND.n4997 GND.n4593 585
R13330 GND.n4593 GND.n4592 585
R13331 GND.n4999 GND.n4998 585
R13332 GND.n5000 GND.n4999 585
R13333 GND.n4594 GND.n4591 585
R13334 GND.n4601 GND.n4591 585
R13335 GND.n4992 GND.n4991 585
R13336 GND.n4991 GND.n4990 585
R13337 GND.n4597 GND.n4596 585
R13338 GND.n4606 GND.n4597 585
R13339 GND.n4943 GND.n4622 585
R13340 GND.n4622 GND.n4612 585
R13341 GND.n4945 GND.n4944 585
R13342 GND.n4946 GND.n4945 585
R13343 GND.n4623 GND.n4621 585
R13344 GND.n4621 GND.n4617 585
R13345 GND.n4938 GND.n4937 585
R13346 GND.n4937 GND.n4936 585
R13347 GND.n4626 GND.n4625 585
R13348 GND.n4636 GND.n4626 585
R13349 GND.n4900 GND.n4899 585
R13350 GND.n4900 GND.n4635 585
R13351 GND.n4902 GND.n4901 585
R13352 GND.n4901 GND.n4642 585
R13353 GND.n4903 GND.n4891 585
R13354 GND.n4891 GND.n4648 585
R13355 GND.n4905 GND.n4904 585
R13356 GND.n4906 GND.n4905 585
R13357 GND.n4892 GND.n4890 585
R13358 GND.n4890 GND.n4652 585
R13359 GND.n3020 GND.n3019 585
R13360 GND.n4856 GND.n3020 585
R13361 GND.n7555 GND.n7554 585
R13362 GND.n7554 GND.n7553 585
R13363 GND.n7556 GND.n3014 585
R13364 GND.n4669 GND.n3014 585
R13365 GND.n7558 GND.n7557 585
R13366 GND.n7559 GND.n7558 585
R13367 GND.n2999 GND.n2998 585
R13368 GND.n3001 GND.n2999 585
R13369 GND.n7569 GND.n7568 585
R13370 GND.n7568 GND.n7567 585
R13371 GND.n7570 GND.n2993 585
R13372 GND.n2993 GND.n2992 585
R13373 GND.n7572 GND.n7571 585
R13374 GND.n7573 GND.n7572 585
R13375 GND.n2980 GND.n2979 585
R13376 GND.n2983 GND.n2980 585
R13377 GND.n7583 GND.n7582 585
R13378 GND.n7582 GND.n7581 585
R13379 GND.n7584 GND.n2974 585
R13380 GND.n4820 GND.n2974 585
R13381 GND.n7586 GND.n7585 585
R13382 GND.n7587 GND.n7586 585
R13383 GND.n2962 GND.n2961 585
R13384 GND.n2971 GND.n2962 585
R13385 GND.n7597 GND.n7596 585
R13386 GND.n7596 GND.n7595 585
R13387 GND.n7598 GND.n2956 585
R13388 GND.n2963 GND.n2956 585
R13389 GND.n7600 GND.n7599 585
R13390 GND.n7601 GND.n7600 585
R13391 GND.n2953 GND.n2952 585
R13392 GND.n7602 GND.n2953 585
R13393 GND.n7605 GND.n7604 585
R13394 GND.n7604 GND.n7603 585
R13395 GND.n7606 GND.n2947 585
R13396 GND.n2954 GND.n2947 585
R13397 GND.n7608 GND.n7607 585
R13398 GND.n7608 GND.n1825 585
R13399 GND.n7609 GND.n2946 585
R13400 GND.n7609 GND.n1814 585
R13401 GND.n7611 GND.n7610 585
R13402 GND.n7610 GND.n1773 585
R13403 GND.n7612 GND.n2941 585
R13404 GND.n2941 GND.n1771 585
R13405 GND.n7614 GND.n7613 585
R13406 GND.n7614 GND.n1891 585
R13407 GND.n7615 GND.n2940 585
R13408 GND.n7615 GND.n1894 585
R13409 GND.n7617 GND.n7616 585
R13410 GND.n7616 GND.n1902 585
R13411 GND.n7618 GND.n2935 585
R13412 GND.n2935 GND.n1900 585
R13413 GND.n7620 GND.n7619 585
R13414 GND.n7620 GND.n1904 585
R13415 GND.n7621 GND.n2934 585
R13416 GND.n7621 GND.t84 585
R13417 GND.n7623 GND.n7622 585
R13418 GND.n7622 GND.n1912 585
R13419 GND.n7624 GND.n2929 585
R13420 GND.n2929 GND.n1925 585
R13421 GND.n7626 GND.n7625 585
R13422 GND.n7626 GND.n1922 585
R13423 GND.n7627 GND.n2928 585
R13424 GND.n7627 GND.n1928 585
R13425 GND.n7629 GND.n7628 585
R13426 GND.n7628 GND.n1936 585
R13427 GND.n7630 GND.n2923 585
R13428 GND.n2923 GND.n1935 585
R13429 GND.n7632 GND.n7631 585
R13430 GND.n7632 GND.n1947 585
R13431 GND.n7633 GND.n2922 585
R13432 GND.n7633 GND.n1945 585
R13433 GND.n7635 GND.n7634 585
R13434 GND.n7634 GND.n1950 585
R13435 GND.n7636 GND.n2917 585
R13436 GND.n2917 GND.n1959 585
R13437 GND.n7638 GND.n7637 585
R13438 GND.n7638 GND.n1957 585
R13439 GND.n7639 GND.n2916 585
R13440 GND.n7639 GND.n1970 585
R13441 GND.n7641 GND.n7640 585
R13442 GND.n7640 GND.n1968 585
R13443 GND.n7642 GND.n2911 585
R13444 GND.n2911 GND.n1972 585
R13445 GND.n7644 GND.n7643 585
R13446 GND.n7644 GND.n1980 585
R13447 GND.n7645 GND.n2910 585
R13448 GND.n7645 GND.n1979 585
R13449 GND.n7647 GND.n7646 585
R13450 GND.n7646 GND.n1992 585
R13451 GND.n7648 GND.n2905 585
R13452 GND.n2905 GND.n1990 585
R13453 GND.n7650 GND.n7649 585
R13454 GND.n7650 GND.n1994 585
R13455 GND.n7651 GND.n2904 585
R13456 GND.n7651 GND.n2003 585
R13457 GND.n7653 GND.n7652 585
R13458 GND.n7652 GND.n2002 585
R13459 GND.n7654 GND.n2899 585
R13460 GND.n2899 GND.n2016 585
R13461 GND.n7656 GND.n7655 585
R13462 GND.n7656 GND.n2013 585
R13463 GND.n7657 GND.n2898 585
R13464 GND.n7657 GND.n2019 585
R13465 GND.n7659 GND.n7658 585
R13466 GND.n7658 GND.n2027 585
R13467 GND.n7660 GND.n2041 585
R13468 GND.n2041 GND.n2026 585
R13469 GND.n7662 GND.n7661 585
R13470 GND.n7663 GND.n7662 585
R13471 GND.n2042 GND.n2040 585
R13472 GND.n2040 GND.n2036 585
R13473 GND.n2892 GND.n2891 585
R13474 GND.n2891 GND.n2890 585
R13475 GND.n2045 GND.n2044 585
R13476 GND.n2055 GND.n2045 585
R13477 GND.n2168 GND.n2167 585
R13478 GND.n2167 GND.n2053 585
R13479 GND.n2169 GND.n2162 585
R13480 GND.n2162 GND.n2066 585
R13481 GND.n2171 GND.n2170 585
R13482 GND.n2171 GND.n2064 585
R13483 GND.n2172 GND.n2161 585
R13484 GND.n2172 GND.n2068 585
R13485 GND.n2174 GND.n2173 585
R13486 GND.n2173 GND.n2076 585
R13487 GND.n2175 GND.n2156 585
R13488 GND.n2156 GND.n2075 585
R13489 GND.n2177 GND.n2176 585
R13490 GND.n2177 GND.n2088 585
R13491 GND.n2178 GND.n2155 585
R13492 GND.n2178 GND.n2086 585
R13493 GND.n2180 GND.n2179 585
R13494 GND.n2179 GND.n2090 585
R13495 GND.n2181 GND.n2152 585
R13496 GND.n2152 GND.n2099 585
R13497 GND.n2183 GND.n2182 585
R13498 GND.n2183 GND.n2098 585
R13499 GND.n2794 GND.n2793 585
R13500 GND.n2793 GND.n2792 585
R13501 GND.n2795 GND.n2148 585
R13502 GND.n2184 GND.n2148 585
R13503 GND.n2798 GND.n2797 585
R13504 GND.n2799 GND.n2798 585
R13505 GND.n2150 GND.n2147 585
R13506 GND.n2147 GND.n2142 585
R13507 GND.n2129 GND.n2128 585
R13508 GND.n2134 GND.n2129 585
R13509 GND.n2811 GND.n2810 585
R13510 GND.n2810 GND.n2809 585
R13511 GND.n2813 GND.n2126 585
R13512 GND.n2130 GND.n2126 585
R13513 GND.n2815 GND.n2814 585
R13514 GND.n2816 GND.n2815 585
R13515 GND.n2127 GND.n2125 585
R13516 GND.n2125 GND.n2119 585
R13517 GND.n2674 GND.n2673 585
R13518 GND.n2673 GND.n2116 585
R13519 GND.n2675 GND.n2668 585
R13520 GND.n2668 GND.n2667 585
R13521 GND.n2677 GND.n2676 585
R13522 GND.n2677 GND.n2196 585
R13523 GND.n2678 GND.n2665 585
R13524 GND.n2678 GND.n2207 585
R13525 GND.n2680 GND.n2679 585
R13526 GND.n2679 GND.n2204 585
R13527 GND.n2681 GND.n2660 585
R13528 GND.n2660 GND.n2210 585
R13529 GND.n2683 GND.n2682 585
R13530 GND.n2683 GND.n2218 585
R13531 GND.n2684 GND.n2659 585
R13532 GND.n2684 GND.n2217 585
R13533 GND.n2686 GND.n2685 585
R13534 GND.n2685 GND.n2229 585
R13535 GND.n2687 GND.n2654 585
R13536 GND.n2654 GND.n2227 585
R13537 GND.n2689 GND.n2688 585
R13538 GND.n2689 GND.n2232 585
R13539 GND.n2690 GND.n2653 585
R13540 GND.n2690 GND.n2241 585
R13541 GND.n2692 GND.n2691 585
R13542 GND.n2691 GND.n2239 585
R13543 GND.n2693 GND.n2256 585
R13544 GND.n2256 GND.n2251 585
R13545 GND.n2695 GND.n2694 585
R13546 GND.n2696 GND.n2695 585
R13547 GND.n2257 GND.n2255 585
R13548 GND.n2255 GND.n2253 585
R13549 GND.n2647 GND.n2646 585
R13550 GND.n2646 GND.n2645 585
R13551 GND.n2260 GND.n2259 585
R13552 GND.n2271 GND.n2260 585
R13553 GND.n2469 GND.n2468 585
R13554 GND.n2468 GND.n2269 585
R13555 GND.n2470 GND.n2463 585
R13556 GND.n2463 GND.n2273 585
R13557 GND.n2472 GND.n2471 585
R13558 GND.n2472 GND.n2281 585
R13559 GND.n2473 GND.n2462 585
R13560 GND.n2473 GND.n2280 585
R13561 GND.n2475 GND.n2474 585
R13562 GND.n2474 GND.n2293 585
R13563 GND.n2476 GND.n2457 585
R13564 GND.n2457 GND.n2291 585
R13565 GND.n2478 GND.n2477 585
R13566 GND.n2478 GND.n2295 585
R13567 GND.n2479 GND.n2456 585
R13568 GND.n2479 GND.n2304 585
R13569 GND.n2481 GND.n2480 585
R13570 GND.n2480 GND.n2303 585
R13571 GND.n2482 GND.n2451 585
R13572 GND.n2451 GND.n2317 585
R13573 GND.n2484 GND.n2483 585
R13574 GND.n2484 GND.n2314 585
R13575 GND.n2485 GND.n2450 585
R13576 GND.n2485 GND.n2320 585
R13577 GND.n2487 GND.n2486 585
R13578 GND.n2486 GND.n2328 585
R13579 GND.n2488 GND.n2445 585
R13580 GND.n2445 GND.n2327 585
R13581 GND.n2490 GND.n2489 585
R13582 GND.n2490 GND.n2339 585
R13583 GND.n2491 GND.n2444 585
R13584 GND.n2491 GND.n2337 585
R13585 GND.n2493 GND.n2492 585
R13586 GND.n2492 GND.n2342 585
R13587 GND.n2494 GND.n2439 585
R13588 GND.n2439 GND.n2351 585
R13589 GND.n2496 GND.n2495 585
R13590 GND.n2496 GND.n2349 585
R13591 GND.n2497 GND.n2438 585
R13592 GND.n2497 GND.n2362 585
R13593 GND.n2499 GND.n2498 585
R13594 GND.n2498 GND.n2360 585
R13595 GND.n2500 GND.n2425 585
R13596 GND.n2425 GND.n2364 585
R13597 GND.n2502 GND.n2501 585
R13598 GND.n2503 GND.n2502 585
R13599 GND.n2426 GND.n2424 585
R13600 GND.n2424 GND.t101 585
R13601 GND.n2432 GND.n2431 585
R13602 GND.n2431 GND.n1549 585
R13603 GND.n2430 GND.n2429 585
R13604 GND.n2430 GND.n1546 585
R13605 GND.n1525 GND.n1524 585
R13606 GND.n1530 GND.n1525 585
R13607 GND.n8089 GND.n8088 585
R13608 GND.n8088 GND.n8087 585
R13609 GND.n8090 GND.n1514 585
R13610 GND.n1526 GND.n1514 585
R13611 GND.n8092 GND.n8091 585
R13612 GND.n8093 GND.n8092 585
R13613 GND.n1515 GND.n1513 585
R13614 GND.n1513 GND.n1509 585
R13615 GND.n1518 GND.n1517 585
R13616 GND.n1517 GND.n1464 585
R13617 GND.n1451 GND.n1450 585
R13618 GND.n8152 GND.n1451 585
R13619 GND.n8155 GND.n8154 585
R13620 GND.n8154 GND.n8153 585
R13621 GND.n8156 GND.n1445 585
R13622 GND.n1445 GND.n1444 585
R13623 GND.n8158 GND.n8157 585
R13624 GND.n8159 GND.n8158 585
R13625 GND.n1443 GND.n1442 585
R13626 GND.n8160 GND.n1443 585
R13627 GND.n8163 GND.n8162 585
R13628 GND.n8162 GND.n8161 585
R13629 GND.n8164 GND.n1437 585
R13630 GND.n1437 GND.n1436 585
R13631 GND.n8166 GND.n8165 585
R13632 GND.n8167 GND.n8166 585
R13633 GND.n1434 GND.n1433 585
R13634 GND.n8168 GND.n1434 585
R13635 GND.n8171 GND.n8170 585
R13636 GND.n8170 GND.n8169 585
R13637 GND.n8172 GND.n1431 585
R13638 GND.n1435 GND.n1431 585
R13639 GND.n8173 GND.n1428 585
R13640 GND.n1428 GND.n1427 585
R13641 GND.n7292 GND.n7291 585
R13642 GND.n7293 GND.n7292 585
R13643 GND.n7290 GND.n3314 585
R13644 GND.n3324 GND.n3316 585
R13645 GND.n7283 GND.n3325 585
R13646 GND.n7282 GND.n3326 585
R13647 GND.n3328 GND.n3327 585
R13648 GND.n7275 GND.n3334 585
R13649 GND.n7274 GND.n3335 585
R13650 GND.n3342 GND.n3336 585
R13651 GND.n7267 GND.n3343 585
R13652 GND.n7266 GND.n3344 585
R13653 GND.n3348 GND.n3345 585
R13654 GND.n7259 GND.n7258 585
R13655 GND.n548 GND.n479 585
R13656 GND.n9612 GND.n479 585
R13657 GND.n9523 GND.n9522 585
R13658 GND.n9524 GND.n9523 585
R13659 GND.n9521 GND.n552 585
R13660 GND.n561 GND.n552 585
R13661 GND.n559 GND.n553 585
R13662 GND.n9516 GND.n559 585
R13663 GND.n575 GND.n573 585
R13664 GND.n573 GND.n572 585
R13665 GND.n9505 GND.n9504 585
R13666 GND.n9506 GND.n9505 585
R13667 GND.n574 GND.n571 585
R13668 GND.n9499 GND.n571 585
R13669 GND.n7102 GND.n7101 585
R13670 GND.n7101 GND.n579 585
R13671 GND.n7100 GND.n3567 585
R13672 GND.n7100 GND.n7099 585
R13673 GND.n3568 GND.n3566 585
R13674 GND.n3580 GND.n3568 585
R13675 GND.n7088 GND.n7087 585
R13676 GND.n7089 GND.n7088 585
R13677 GND.n7086 GND.n3560 585
R13678 GND.n7086 GND.n7085 585
R13679 GND.n3582 GND.n3559 585
R13680 GND.n3584 GND.n3582 585
R13681 GND.n3594 GND.n3558 585
R13682 GND.n7066 GND.n3594 585
R13683 GND.n7054 GND.n7053 585
R13684 GND.n7054 GND.n3591 585
R13685 GND.n7055 GND.n3552 585
R13686 GND.n7056 GND.n7055 585
R13687 GND.n7052 GND.n3551 585
R13688 GND.n7052 GND.n7051 585
R13689 GND.n3603 GND.n3550 585
R13690 GND.n3605 GND.n3603 585
R13691 GND.n3615 GND.n3614 585
R13692 GND.n7038 GND.n3615 585
R13693 GND.n7026 GND.n3544 585
R13694 GND.n7026 GND.n3612 585
R13695 GND.n7027 GND.n3543 585
R13696 GND.n7028 GND.n7027 585
R13697 GND.n7025 GND.n3542 585
R13698 GND.n7025 GND.n7024 585
R13699 GND.n3626 GND.n3625 585
R13700 GND.n3627 GND.n3626 585
R13701 GND.n3637 GND.n3536 585
R13702 GND.n7011 GND.n3637 585
R13703 GND.n6999 GND.n3535 585
R13704 GND.n6999 GND.n3635 585
R13705 GND.n7000 GND.n3534 585
R13706 GND.n7001 GND.n7000 585
R13707 GND.n6998 GND.n3648 585
R13708 GND.n6998 GND.n6997 585
R13709 GND.n3647 GND.n3528 585
R13710 GND.n3649 GND.n3647 585
R13711 GND.n3660 GND.n3527 585
R13712 GND.n6985 GND.n3660 585
R13713 GND.n6972 GND.n3526 585
R13714 GND.n6972 GND.n3657 585
R13715 GND.n6974 GND.n6973 585
R13716 GND.n6975 GND.n6974 585
R13717 GND.n6971 GND.n3520 585
R13718 GND.n6971 GND.n6970 585
R13719 GND.n3669 GND.n3519 585
R13720 GND.n3671 GND.n3669 585
R13721 GND.n3680 GND.n3518 585
R13722 GND.n6958 GND.n3680 585
R13723 GND.n6946 GND.n6944 585
R13724 GND.n6946 GND.n6945 585
R13725 GND.n6947 GND.n3512 585
R13726 GND.n6948 GND.n6947 585
R13727 GND.n6943 GND.n3511 585
R13728 GND.n6943 GND.n6942 585
R13729 GND.n3689 GND.n3510 585
R13730 GND.n3691 GND.n3689 585
R13731 GND.n3701 GND.n3700 585
R13732 GND.n6929 GND.n3701 585
R13733 GND.n6917 GND.n3504 585
R13734 GND.n6917 GND.n3698 585
R13735 GND.n6918 GND.n3503 585
R13736 GND.n6919 GND.n6918 585
R13737 GND.n6916 GND.n3502 585
R13738 GND.n6916 GND.n6915 585
R13739 GND.n3712 GND.n3711 585
R13740 GND.n3713 GND.n3712 585
R13741 GND.n3723 GND.n3496 585
R13742 GND.n6902 GND.n3723 585
R13743 GND.n6890 GND.n3495 585
R13744 GND.n6890 GND.n3721 585
R13745 GND.n6891 GND.n3494 585
R13746 GND.n6892 GND.n6891 585
R13747 GND.n6889 GND.n3734 585
R13748 GND.n6889 GND.n6888 585
R13749 GND.n3733 GND.n3488 585
R13750 GND.n3735 GND.n3733 585
R13751 GND.n6830 GND.n3487 585
R13752 GND.n6840 GND.n6830 585
R13753 GND.n6850 GND.n3486 585
R13754 GND.n6850 GND.n6849 585
R13755 GND.n6852 GND.n6851 585
R13756 GND.n6853 GND.n6852 585
R13757 GND.n6829 GND.n3480 585
R13758 GND.n6829 GND.n6828 585
R13759 GND.n6819 GND.n3479 585
R13760 GND.n6860 GND.n6819 585
R13761 GND.n3763 GND.n3478 585
R13762 GND.n6811 GND.n3763 585
R13763 GND.n6868 GND.n3764 585
R13764 GND.n6868 GND.n6867 585
R13765 GND.n6869 GND.n3472 585
R13766 GND.n6870 GND.n6869 585
R13767 GND.n3762 GND.n3471 585
R13768 GND.n6802 GND.n3762 585
R13769 GND.n3753 GND.n3470 585
R13770 GND.n6877 GND.n3753 585
R13771 GND.n3780 GND.n3779 585
R13772 GND.n3780 GND.n3750 585
R13773 GND.n3781 GND.n3464 585
R13774 GND.n3782 GND.n3781 585
R13775 GND.n3776 GND.n3463 585
R13776 GND.n6793 GND.n3776 585
R13777 GND.n6779 GND.n3462 585
R13778 GND.n6779 GND.n6778 585
R13779 GND.n6781 GND.n6780 585
R13780 GND.n6782 GND.n6781 585
R13781 GND.n6777 GND.n3456 585
R13782 GND.n6777 GND.n6776 585
R13783 GND.n3791 GND.n3455 585
R13784 GND.n3804 GND.n3791 585
R13785 GND.n3801 GND.n3454 585
R13786 GND.n6767 GND.n3801 585
R13787 GND.n6755 GND.n6753 585
R13788 GND.n6755 GND.n6754 585
R13789 GND.n6756 GND.n3448 585
R13790 GND.n6757 GND.n6756 585
R13791 GND.n6752 GND.n3447 585
R13792 GND.n6752 GND.n6751 585
R13793 GND.n3813 GND.n3446 585
R13794 GND.n3827 GND.n3813 585
R13795 GND.n3825 GND.n3824 585
R13796 GND.n6742 GND.n3825 585
R13797 GND.n6730 GND.n3440 585
R13798 GND.n6730 GND.n6729 585
R13799 GND.n6731 GND.n3439 585
R13800 GND.n6732 GND.n6731 585
R13801 GND.n6728 GND.n3438 585
R13802 GND.n6728 GND.n6727 585
R13803 GND.n3838 GND.n3837 585
R13804 GND.n3850 GND.n3838 585
R13805 GND.n3848 GND.n3432 585
R13806 GND.n6718 GND.n3848 585
R13807 GND.n6706 GND.n3431 585
R13808 GND.n6706 GND.n6705 585
R13809 GND.n6707 GND.n3430 585
R13810 GND.n6708 GND.n6707 585
R13811 GND.n6703 GND.n3860 585
R13812 GND.n6703 GND.n6702 585
R13813 GND.n3859 GND.n3424 585
R13814 GND.n3873 GND.n3859 585
R13815 GND.n3871 GND.n3423 585
R13816 GND.n6693 GND.n3871 585
R13817 GND.n6680 GND.n3422 585
R13818 GND.n6680 GND.n6679 585
R13819 GND.n6682 GND.n6681 585
R13820 GND.n6683 GND.n6682 585
R13821 GND.n6678 GND.n3416 585
R13822 GND.n6678 GND.n6677 585
R13823 GND.n3882 GND.n3415 585
R13824 GND.n3895 GND.n3882 585
R13825 GND.n3892 GND.n3414 585
R13826 GND.n6668 GND.n3892 585
R13827 GND.n6656 GND.n6654 585
R13828 GND.n6656 GND.n6655 585
R13829 GND.n6657 GND.n3408 585
R13830 GND.n6658 GND.n6657 585
R13831 GND.n6653 GND.n3407 585
R13832 GND.n6653 GND.n6652 585
R13833 GND.n3904 GND.n3406 585
R13834 GND.n3918 GND.n3904 585
R13835 GND.n3916 GND.n3915 585
R13836 GND.n6643 GND.n3916 585
R13837 GND.n6631 GND.n3400 585
R13838 GND.n6631 GND.n6630 585
R13839 GND.n6632 GND.n3399 585
R13840 GND.n6633 GND.n6632 585
R13841 GND.n6629 GND.n3398 585
R13842 GND.n6629 GND.n6628 585
R13843 GND.n3929 GND.n3928 585
R13844 GND.n3941 GND.n3929 585
R13845 GND.n3939 GND.n3392 585
R13846 GND.n6619 GND.n3939 585
R13847 GND.n6607 GND.n3391 585
R13848 GND.n6607 GND.n6606 585
R13849 GND.n6608 GND.n3390 585
R13850 GND.n6609 GND.n6608 585
R13851 GND.n6604 GND.n3951 585
R13852 GND.n6604 GND.n6603 585
R13853 GND.n3950 GND.n3384 585
R13854 GND.n6584 GND.n3950 585
R13855 GND.n3961 GND.n3383 585
R13856 GND.n6594 GND.n3961 585
R13857 GND.n6581 GND.n3382 585
R13858 GND.n6582 GND.n6581 585
R13859 GND.n3373 GND.n3371 585
R13860 GND.n6437 GND.n3371 585
R13861 GND.n7249 GND.n7248 585
R13862 GND.n7250 GND.n7249 585
R13863 GND.n3372 GND.n3370 585
R13864 GND.n3376 GND.n3370 585
R13865 GND.n6324 GND.n3313 585
R13866 GND.n7256 GND.n3313 585
R13867 GND.n9547 GND.n475 585
R13868 GND.n9548 GND.n9546 585
R13869 GND.n9549 GND.n9543 585
R13870 GND.n9541 GND.n9540 585
R13871 GND.n9553 GND.n9539 585
R13872 GND.n9554 GND.n9538 585
R13873 GND.n9555 GND.n9537 585
R13874 GND.n9535 GND.n9534 585
R13875 GND.n9559 GND.n9533 585
R13876 GND.n9560 GND.n9532 585
R13877 GND.n9561 GND.n9531 585
R13878 GND.n546 GND.n545 585
R13879 GND.n9566 GND.n9565 585
R13880 GND.n9567 GND.n9566 585
R13881 GND.n9614 GND.n9613 585
R13882 GND.n9613 GND.n9612 585
R13883 GND.n474 GND.n472 585
R13884 GND.n9524 GND.n474 585
R13885 GND.n9618 GND.n471 585
R13886 GND.n561 GND.n471 585
R13887 GND.n9619 GND.n470 585
R13888 GND.n9516 GND.n470 585
R13889 GND.n9620 GND.n469 585
R13890 GND.n572 GND.n469 585
R13891 GND.n569 GND.n467 585
R13892 GND.n9506 GND.n569 585
R13893 GND.n9624 GND.n466 585
R13894 GND.n9499 GND.n466 585
R13895 GND.n9625 GND.n465 585
R13896 GND.n579 GND.n465 585
R13897 GND.n9626 GND.n464 585
R13898 GND.n7099 GND.n464 585
R13899 GND.n3579 GND.n462 585
R13900 GND.n3580 GND.n3579 585
R13901 GND.n9630 GND.n461 585
R13902 GND.n7089 GND.n461 585
R13903 GND.n9631 GND.n460 585
R13904 GND.n7085 GND.n460 585
R13905 GND.n9632 GND.n459 585
R13906 GND.n3584 GND.n459 585
R13907 GND.n3592 GND.n457 585
R13908 GND.n7066 GND.n3592 585
R13909 GND.n9636 GND.n456 585
R13910 GND.n3591 GND.n456 585
R13911 GND.n9637 GND.n455 585
R13912 GND.n7056 GND.n455 585
R13913 GND.n9638 GND.n454 585
R13914 GND.n7051 GND.n454 585
R13915 GND.n3604 GND.n452 585
R13916 GND.n3605 GND.n3604 585
R13917 GND.n9642 GND.n451 585
R13918 GND.n7038 GND.n451 585
R13919 GND.n9643 GND.n450 585
R13920 GND.n3612 GND.n450 585
R13921 GND.n9644 GND.n449 585
R13922 GND.n7028 GND.n449 585
R13923 GND.n7023 GND.n447 585
R13924 GND.n7024 GND.n7023 585
R13925 GND.n9648 GND.n446 585
R13926 GND.n3627 GND.n446 585
R13927 GND.n9649 GND.n445 585
R13928 GND.n7011 GND.n445 585
R13929 GND.n9650 GND.n444 585
R13930 GND.n3635 GND.n444 585
R13931 GND.n3645 GND.n442 585
R13932 GND.n7001 GND.n3645 585
R13933 GND.n9654 GND.n441 585
R13934 GND.n6997 GND.n441 585
R13935 GND.n9655 GND.n440 585
R13936 GND.n3649 GND.n440 585
R13937 GND.n9656 GND.n439 585
R13938 GND.n6985 GND.n439 585
R13939 GND.n3656 GND.n437 585
R13940 GND.n3657 GND.n3656 585
R13941 GND.n9660 GND.n436 585
R13942 GND.n6975 GND.n436 585
R13943 GND.n9661 GND.n435 585
R13944 GND.n6970 GND.n435 585
R13945 GND.n9662 GND.n434 585
R13946 GND.n3671 GND.n434 585
R13947 GND.n3678 GND.n432 585
R13948 GND.n6958 GND.n3678 585
R13949 GND.n9666 GND.n431 585
R13950 GND.n6945 GND.n431 585
R13951 GND.n9667 GND.n430 585
R13952 GND.n6948 GND.n430 585
R13953 GND.n9668 GND.n429 585
R13954 GND.n6942 GND.n429 585
R13955 GND.n3690 GND.n427 585
R13956 GND.n3691 GND.n3690 585
R13957 GND.n9672 GND.n426 585
R13958 GND.n6929 GND.n426 585
R13959 GND.n9673 GND.n425 585
R13960 GND.n3698 GND.n425 585
R13961 GND.n9674 GND.n424 585
R13962 GND.n6919 GND.n424 585
R13963 GND.n6914 GND.n422 585
R13964 GND.n6915 GND.n6914 585
R13965 GND.n9678 GND.n421 585
R13966 GND.n3713 GND.n421 585
R13967 GND.n9679 GND.n420 585
R13968 GND.n6902 GND.n420 585
R13969 GND.n9680 GND.n419 585
R13970 GND.n3721 GND.n419 585
R13971 GND.n3731 GND.n417 585
R13972 GND.n6892 GND.n3731 585
R13973 GND.n9684 GND.n416 585
R13974 GND.n6888 GND.n416 585
R13975 GND.n9685 GND.n415 585
R13976 GND.n3735 GND.n415 585
R13977 GND.n9686 GND.n414 585
R13978 GND.n6840 GND.n414 585
R13979 GND.n6831 GND.n412 585
R13980 GND.n6849 GND.n6831 585
R13981 GND.n9690 GND.n411 585
R13982 GND.n6853 GND.n411 585
R13983 GND.n9691 GND.n410 585
R13984 GND.n6828 GND.n410 585
R13985 GND.n9692 GND.n409 585
R13986 GND.n6860 GND.n409 585
R13987 GND.n6810 GND.n408 585
R13988 GND.n6811 GND.n6810 585
R13989 GND.n6809 GND.n6808 585
R13990 GND.n6867 GND.n6809 585
R13991 GND.n3765 GND.n3760 585
R13992 GND.n6870 GND.n3760 585
R13993 GND.n6804 GND.n6803 585
R13994 GND.n6803 GND.n6802 585
R13995 GND.n6800 GND.n3751 585
R13996 GND.n6877 GND.n3751 585
R13997 GND.n6799 GND.n3768 585
R13998 GND.n3768 GND.n3750 585
R13999 GND.n3772 GND.n3767 585
R14000 GND.n3782 GND.n3772 585
R14001 GND.n6795 GND.n6794 585
R14002 GND.n6794 GND.n6793 585
R14003 GND.n3771 GND.n3770 585
R14004 GND.n6778 GND.n3771 585
R14005 GND.n3795 GND.n3789 585
R14006 GND.n6782 GND.n3789 585
R14007 GND.n6775 GND.n6774 585
R14008 GND.n6776 GND.n6775 585
R14009 GND.n3794 GND.n3793 585
R14010 GND.n3804 GND.n3793 585
R14011 GND.n6769 GND.n6768 585
R14012 GND.n6768 GND.n6767 585
R14013 GND.n3798 GND.n3797 585
R14014 GND.n6754 GND.n3798 585
R14015 GND.n3818 GND.n3811 585
R14016 GND.n6757 GND.n3811 585
R14017 GND.n6750 GND.n6749 585
R14018 GND.n6751 GND.n6750 585
R14019 GND.n3817 GND.n3816 585
R14020 GND.n3827 GND.n3816 585
R14021 GND.n6744 GND.n6743 585
R14022 GND.n6743 GND.n6742 585
R14023 GND.n3821 GND.n3820 585
R14024 GND.n6729 GND.n3821 585
R14025 GND.n3842 GND.n3835 585
R14026 GND.n6732 GND.n3835 585
R14027 GND.n6726 GND.n6725 585
R14028 GND.n6727 GND.n6726 585
R14029 GND.n3841 GND.n3840 585
R14030 GND.n3850 GND.n3840 585
R14031 GND.n6720 GND.n6719 585
R14032 GND.n6719 GND.n6718 585
R14033 GND.n3845 GND.n3844 585
R14034 GND.n6705 GND.n3845 585
R14035 GND.n3864 GND.n3857 585
R14036 GND.n6708 GND.n3857 585
R14037 GND.n6701 GND.n6700 585
R14038 GND.n6702 GND.n6701 585
R14039 GND.n3863 GND.n3862 585
R14040 GND.n3873 GND.n3862 585
R14041 GND.n6695 GND.n6694 585
R14042 GND.n6694 GND.n6693 585
R14043 GND.n3867 GND.n3866 585
R14044 GND.n6679 GND.n3867 585
R14045 GND.n3886 GND.n3880 585
R14046 GND.n6683 GND.n3880 585
R14047 GND.n6676 GND.n6675 585
R14048 GND.n6677 GND.n6676 585
R14049 GND.n3885 GND.n3884 585
R14050 GND.n3895 GND.n3884 585
R14051 GND.n6670 GND.n6669 585
R14052 GND.n6669 GND.n6668 585
R14053 GND.n3889 GND.n3888 585
R14054 GND.n6655 GND.n3889 585
R14055 GND.n3909 GND.n3902 585
R14056 GND.n6658 GND.n3902 585
R14057 GND.n6651 GND.n6650 585
R14058 GND.n6652 GND.n6651 585
R14059 GND.n3908 GND.n3907 585
R14060 GND.n3918 GND.n3907 585
R14061 GND.n6645 GND.n6644 585
R14062 GND.n6644 GND.n6643 585
R14063 GND.n3912 GND.n3911 585
R14064 GND.n6630 GND.n3912 585
R14065 GND.n3933 GND.n3926 585
R14066 GND.n6633 GND.n3926 585
R14067 GND.n6627 GND.n6626 585
R14068 GND.n6628 GND.n6627 585
R14069 GND.n3932 GND.n3931 585
R14070 GND.n3941 GND.n3931 585
R14071 GND.n6621 GND.n6620 585
R14072 GND.n6620 GND.n6619 585
R14073 GND.n3936 GND.n3935 585
R14074 GND.n6606 GND.n3936 585
R14075 GND.n3954 GND.n3948 585
R14076 GND.n6609 GND.n3948 585
R14077 GND.n6602 GND.n6601 585
R14078 GND.n6603 GND.n6602 585
R14079 GND.n3953 GND.n3952 585
R14080 GND.n6584 GND.n3952 585
R14081 GND.n6596 GND.n6595 585
R14082 GND.n6595 GND.n6594 585
R14083 GND.n3957 GND.n3956 585
R14084 GND.n6582 GND.n3957 585
R14085 GND.n6436 GND.n6435 585
R14086 GND.n6437 GND.n6436 585
R14087 GND.n3962 GND.n3368 585
R14088 GND.n7250 GND.n3368 585
R14089 GND.n6431 GND.n3354 585
R14090 GND.n3376 GND.n3354 585
R14091 GND.n7257 GND.n3355 585
R14092 GND.n7257 GND.n7256 585
R14093 GND.n6256 GND.n3270 545.355
R14094 GND.n6142 GND.n6141 545.355
R14095 GND.n4809 GND.n4808 545.355
R14096 GND.n4721 GND.n2966 545.355
R14097 GND.n9455 GND.n616 496.853
R14098 GND.n9324 GND.n9323 301.784
R14099 GND.n9324 GND.n694 301.784
R14100 GND.n9332 GND.n694 301.784
R14101 GND.n9333 GND.n9332 301.784
R14102 GND.n9334 GND.n9333 301.784
R14103 GND.n9334 GND.n688 301.784
R14104 GND.n9342 GND.n688 301.784
R14105 GND.n9343 GND.n9342 301.784
R14106 GND.n9344 GND.n9343 301.784
R14107 GND.n9344 GND.n682 301.784
R14108 GND.n9352 GND.n682 301.784
R14109 GND.n9353 GND.n9352 301.784
R14110 GND.n9354 GND.n9353 301.784
R14111 GND.n9354 GND.n676 301.784
R14112 GND.n9362 GND.n676 301.784
R14113 GND.n9363 GND.n9362 301.784
R14114 GND.n9364 GND.n9363 301.784
R14115 GND.n9364 GND.n670 301.784
R14116 GND.n9372 GND.n670 301.784
R14117 GND.n9373 GND.n9372 301.784
R14118 GND.n9374 GND.n9373 301.784
R14119 GND.n9374 GND.n664 301.784
R14120 GND.n9382 GND.n664 301.784
R14121 GND.n9383 GND.n9382 301.784
R14122 GND.n9384 GND.n9383 301.784
R14123 GND.n9384 GND.n658 301.784
R14124 GND.n9392 GND.n658 301.784
R14125 GND.n9393 GND.n9392 301.784
R14126 GND.n9394 GND.n9393 301.784
R14127 GND.n9394 GND.n652 301.784
R14128 GND.n9402 GND.n652 301.784
R14129 GND.n9403 GND.n9402 301.784
R14130 GND.n9404 GND.n9403 301.784
R14131 GND.n9404 GND.n646 301.784
R14132 GND.n9412 GND.n646 301.784
R14133 GND.n9413 GND.n9412 301.784
R14134 GND.n9414 GND.n9413 301.784
R14135 GND.n9414 GND.n640 301.784
R14136 GND.n9422 GND.n640 301.784
R14137 GND.n9423 GND.n9422 301.784
R14138 GND.n9424 GND.n9423 301.784
R14139 GND.n9424 GND.n634 301.784
R14140 GND.n9432 GND.n634 301.784
R14141 GND.n9433 GND.n9432 301.784
R14142 GND.n9434 GND.n9433 301.784
R14143 GND.n9434 GND.n628 301.784
R14144 GND.n9442 GND.n628 301.784
R14145 GND.n9443 GND.n9442 301.784
R14146 GND.n9444 GND.n9443 301.784
R14147 GND.n9444 GND.n622 301.784
R14148 GND.n9453 GND.n622 301.784
R14149 GND.n9454 GND.n9453 301.784
R14150 GND.n9455 GND.n9454 301.784
R14151 GND.n57 GND.n43 289.615
R14152 GND.n80 GND.n66 289.615
R14153 GND.n100 GND.n86 289.615
R14154 GND.n123 GND.n109 289.615
R14155 GND.n14 GND.n0 289.615
R14156 GND.n37 GND.n23 289.615
R14157 GND.n312 GND.n298 289.615
R14158 GND.n289 GND.n275 289.615
R14159 GND.n355 GND.n341 289.615
R14160 GND.n332 GND.n318 289.615
R14161 GND.n399 GND.n385 289.615
R14162 GND.n376 GND.n362 289.615
R14163 GND.n197 GND.n191 289.615
R14164 GND.n185 GND.n179 289.615
R14165 GND.n173 GND.n167 289.615
R14166 GND.n161 GND.n155 289.615
R14167 GND.n149 GND.n143 289.615
R14168 GND.n138 GND.n132 289.615
R14169 GND.n268 GND.n262 289.615
R14170 GND.n256 GND.n250 289.615
R14171 GND.n244 GND.n238 289.615
R14172 GND.n232 GND.n226 289.615
R14173 GND.n220 GND.n214 289.615
R14174 GND.n209 GND.n203 289.615
R14175 GND.n8292 GND.n1318 280.613
R14176 GND.n8293 GND.n8292 280.613
R14177 GND.n8294 GND.n8293 280.613
R14178 GND.n8294 GND.n1312 280.613
R14179 GND.n8302 GND.n1312 280.613
R14180 GND.n8303 GND.n8302 280.613
R14181 GND.n8304 GND.n8303 280.613
R14182 GND.n8304 GND.n1306 280.613
R14183 GND.n8312 GND.n1306 280.613
R14184 GND.n8313 GND.n8312 280.613
R14185 GND.n8314 GND.n8313 280.613
R14186 GND.n8314 GND.n1300 280.613
R14187 GND.n8322 GND.n1300 280.613
R14188 GND.n8323 GND.n8322 280.613
R14189 GND.n8324 GND.n8323 280.613
R14190 GND.n8324 GND.n1294 280.613
R14191 GND.n8332 GND.n1294 280.613
R14192 GND.n8333 GND.n8332 280.613
R14193 GND.n8334 GND.n8333 280.613
R14194 GND.n8334 GND.n1288 280.613
R14195 GND.n8342 GND.n1288 280.613
R14196 GND.n8343 GND.n8342 280.613
R14197 GND.n8344 GND.n8343 280.613
R14198 GND.n8344 GND.n1282 280.613
R14199 GND.n8352 GND.n1282 280.613
R14200 GND.n8353 GND.n8352 280.613
R14201 GND.n8354 GND.n8353 280.613
R14202 GND.n8354 GND.n1276 280.613
R14203 GND.n8362 GND.n1276 280.613
R14204 GND.n8363 GND.n8362 280.613
R14205 GND.n8364 GND.n8363 280.613
R14206 GND.n8364 GND.n1270 280.613
R14207 GND.n8372 GND.n1270 280.613
R14208 GND.n8373 GND.n8372 280.613
R14209 GND.n8374 GND.n8373 280.613
R14210 GND.n8374 GND.n1264 280.613
R14211 GND.n8382 GND.n1264 280.613
R14212 GND.n8383 GND.n8382 280.613
R14213 GND.n8384 GND.n8383 280.613
R14214 GND.n8384 GND.n1258 280.613
R14215 GND.n8392 GND.n1258 280.613
R14216 GND.n8393 GND.n8392 280.613
R14217 GND.n8394 GND.n8393 280.613
R14218 GND.n8394 GND.n1252 280.613
R14219 GND.n8402 GND.n1252 280.613
R14220 GND.n8403 GND.n8402 280.613
R14221 GND.n8404 GND.n8403 280.613
R14222 GND.n8404 GND.n1246 280.613
R14223 GND.n8412 GND.n1246 280.613
R14224 GND.n8413 GND.n8412 280.613
R14225 GND.n8414 GND.n8413 280.613
R14226 GND.n8414 GND.n1240 280.613
R14227 GND.n8422 GND.n1240 280.613
R14228 GND.n8423 GND.n8422 280.613
R14229 GND.n8424 GND.n8423 280.613
R14230 GND.n8424 GND.n1234 280.613
R14231 GND.n8432 GND.n1234 280.613
R14232 GND.n8433 GND.n8432 280.613
R14233 GND.n8434 GND.n8433 280.613
R14234 GND.n8434 GND.n1228 280.613
R14235 GND.n8442 GND.n1228 280.613
R14236 GND.n8443 GND.n8442 280.613
R14237 GND.n8444 GND.n8443 280.613
R14238 GND.n8444 GND.n1222 280.613
R14239 GND.n8452 GND.n1222 280.613
R14240 GND.n8453 GND.n8452 280.613
R14241 GND.n8454 GND.n8453 280.613
R14242 GND.n8454 GND.n1216 280.613
R14243 GND.n8462 GND.n1216 280.613
R14244 GND.n8463 GND.n8462 280.613
R14245 GND.n8464 GND.n8463 280.613
R14246 GND.n8464 GND.n1210 280.613
R14247 GND.n8472 GND.n1210 280.613
R14248 GND.n8473 GND.n8472 280.613
R14249 GND.n8474 GND.n8473 280.613
R14250 GND.n8474 GND.n1204 280.613
R14251 GND.n8482 GND.n1204 280.613
R14252 GND.n8483 GND.n8482 280.613
R14253 GND.n8484 GND.n8483 280.613
R14254 GND.n8484 GND.n1198 280.613
R14255 GND.n8492 GND.n1198 280.613
R14256 GND.n8493 GND.n8492 280.613
R14257 GND.n8494 GND.n8493 280.613
R14258 GND.n8494 GND.n1192 280.613
R14259 GND.n8502 GND.n1192 280.613
R14260 GND.n8503 GND.n8502 280.613
R14261 GND.n8504 GND.n8503 280.613
R14262 GND.n8504 GND.n1186 280.613
R14263 GND.n8512 GND.n1186 280.613
R14264 GND.n8513 GND.n8512 280.613
R14265 GND.n8514 GND.n8513 280.613
R14266 GND.n8514 GND.n1180 280.613
R14267 GND.n8522 GND.n1180 280.613
R14268 GND.n8523 GND.n8522 280.613
R14269 GND.n8524 GND.n8523 280.613
R14270 GND.n8524 GND.n1174 280.613
R14271 GND.n8532 GND.n1174 280.613
R14272 GND.n8533 GND.n8532 280.613
R14273 GND.n8534 GND.n8533 280.613
R14274 GND.n8534 GND.n1168 280.613
R14275 GND.n8542 GND.n1168 280.613
R14276 GND.n8543 GND.n8542 280.613
R14277 GND.n8544 GND.n8543 280.613
R14278 GND.n8544 GND.n1162 280.613
R14279 GND.n8552 GND.n1162 280.613
R14280 GND.n8553 GND.n8552 280.613
R14281 GND.n8554 GND.n8553 280.613
R14282 GND.n8554 GND.n1156 280.613
R14283 GND.n8562 GND.n1156 280.613
R14284 GND.n8563 GND.n8562 280.613
R14285 GND.n8564 GND.n8563 280.613
R14286 GND.n8564 GND.n1150 280.613
R14287 GND.n8572 GND.n1150 280.613
R14288 GND.n8573 GND.n8572 280.613
R14289 GND.n8574 GND.n8573 280.613
R14290 GND.n8574 GND.n1144 280.613
R14291 GND.n8582 GND.n1144 280.613
R14292 GND.n8583 GND.n8582 280.613
R14293 GND.n8584 GND.n8583 280.613
R14294 GND.n8584 GND.n1138 280.613
R14295 GND.n8592 GND.n1138 280.613
R14296 GND.n8593 GND.n8592 280.613
R14297 GND.n8594 GND.n8593 280.613
R14298 GND.n8594 GND.n1132 280.613
R14299 GND.n8602 GND.n1132 280.613
R14300 GND.n8603 GND.n8602 280.613
R14301 GND.n8604 GND.n8603 280.613
R14302 GND.n8604 GND.n1126 280.613
R14303 GND.n8612 GND.n1126 280.613
R14304 GND.n8613 GND.n8612 280.613
R14305 GND.n8614 GND.n8613 280.613
R14306 GND.n8614 GND.n1120 280.613
R14307 GND.n8622 GND.n1120 280.613
R14308 GND.n8623 GND.n8622 280.613
R14309 GND.n8624 GND.n8623 280.613
R14310 GND.n8624 GND.n1114 280.613
R14311 GND.n8632 GND.n1114 280.613
R14312 GND.n8633 GND.n8632 280.613
R14313 GND.n8634 GND.n8633 280.613
R14314 GND.n8634 GND.n1108 280.613
R14315 GND.n8642 GND.n1108 280.613
R14316 GND.n8643 GND.n8642 280.613
R14317 GND.n8644 GND.n8643 280.613
R14318 GND.n8644 GND.n1102 280.613
R14319 GND.n8652 GND.n1102 280.613
R14320 GND.n8653 GND.n8652 280.613
R14321 GND.n8654 GND.n8653 280.613
R14322 GND.n8654 GND.n1096 280.613
R14323 GND.n8662 GND.n1096 280.613
R14324 GND.n8663 GND.n8662 280.613
R14325 GND.n8664 GND.n8663 280.613
R14326 GND.n8664 GND.n1090 280.613
R14327 GND.n8672 GND.n1090 280.613
R14328 GND.n8673 GND.n8672 280.613
R14329 GND.n8674 GND.n8673 280.613
R14330 GND.n8674 GND.n1084 280.613
R14331 GND.n8682 GND.n1084 280.613
R14332 GND.n8683 GND.n8682 280.613
R14333 GND.n8684 GND.n8683 280.613
R14334 GND.n8684 GND.n1078 280.613
R14335 GND.n8692 GND.n1078 280.613
R14336 GND.n8693 GND.n8692 280.613
R14337 GND.n8694 GND.n8693 280.613
R14338 GND.n8694 GND.n1072 280.613
R14339 GND.n8702 GND.n1072 280.613
R14340 GND.n8703 GND.n8702 280.613
R14341 GND.n8704 GND.n8703 280.613
R14342 GND.n8704 GND.n1066 280.613
R14343 GND.n8712 GND.n1066 280.613
R14344 GND.n8713 GND.n8712 280.613
R14345 GND.n8714 GND.n8713 280.613
R14346 GND.n8714 GND.n1060 280.613
R14347 GND.n8722 GND.n1060 280.613
R14348 GND.n8723 GND.n8722 280.613
R14349 GND.n8724 GND.n8723 280.613
R14350 GND.n8724 GND.n1054 280.613
R14351 GND.n8732 GND.n1054 280.613
R14352 GND.n8733 GND.n8732 280.613
R14353 GND.n8734 GND.n8733 280.613
R14354 GND.n8734 GND.n1048 280.613
R14355 GND.n8742 GND.n1048 280.613
R14356 GND.n8743 GND.n8742 280.613
R14357 GND.n8744 GND.n8743 280.613
R14358 GND.n8744 GND.n1042 280.613
R14359 GND.n8752 GND.n1042 280.613
R14360 GND.n8753 GND.n8752 280.613
R14361 GND.n8754 GND.n8753 280.613
R14362 GND.n8754 GND.n1036 280.613
R14363 GND.n8762 GND.n1036 280.613
R14364 GND.n8763 GND.n8762 280.613
R14365 GND.n8764 GND.n8763 280.613
R14366 GND.n8764 GND.n1030 280.613
R14367 GND.n8772 GND.n1030 280.613
R14368 GND.n8773 GND.n8772 280.613
R14369 GND.n8774 GND.n8773 280.613
R14370 GND.n8774 GND.n1024 280.613
R14371 GND.n8782 GND.n1024 280.613
R14372 GND.n8783 GND.n8782 280.613
R14373 GND.n8784 GND.n8783 280.613
R14374 GND.n8784 GND.n1018 280.613
R14375 GND.n8792 GND.n1018 280.613
R14376 GND.n8793 GND.n8792 280.613
R14377 GND.n8794 GND.n8793 280.613
R14378 GND.n8794 GND.n1012 280.613
R14379 GND.n8802 GND.n1012 280.613
R14380 GND.n8803 GND.n8802 280.613
R14381 GND.n8804 GND.n8803 280.613
R14382 GND.n8804 GND.n1006 280.613
R14383 GND.n8812 GND.n1006 280.613
R14384 GND.n8813 GND.n8812 280.613
R14385 GND.n8814 GND.n8813 280.613
R14386 GND.n8814 GND.n1000 280.613
R14387 GND.n8822 GND.n1000 280.613
R14388 GND.n8823 GND.n8822 280.613
R14389 GND.n8824 GND.n8823 280.613
R14390 GND.n8824 GND.n994 280.613
R14391 GND.n8832 GND.n994 280.613
R14392 GND.n8833 GND.n8832 280.613
R14393 GND.n8834 GND.n8833 280.613
R14394 GND.n8834 GND.n988 280.613
R14395 GND.n8842 GND.n988 280.613
R14396 GND.n8843 GND.n8842 280.613
R14397 GND.n8844 GND.n8843 280.613
R14398 GND.n8844 GND.n982 280.613
R14399 GND.n8852 GND.n982 280.613
R14400 GND.n8853 GND.n8852 280.613
R14401 GND.n8854 GND.n8853 280.613
R14402 GND.n8854 GND.n976 280.613
R14403 GND.n8862 GND.n976 280.613
R14404 GND.n8863 GND.n8862 280.613
R14405 GND.n8864 GND.n8863 280.613
R14406 GND.n8864 GND.n970 280.613
R14407 GND.n8872 GND.n970 280.613
R14408 GND.n8873 GND.n8872 280.613
R14409 GND.n8874 GND.n8873 280.613
R14410 GND.n8874 GND.n964 280.613
R14411 GND.n8882 GND.n964 280.613
R14412 GND.n8883 GND.n8882 280.613
R14413 GND.n8884 GND.n8883 280.613
R14414 GND.n8884 GND.n958 280.613
R14415 GND.n8892 GND.n958 280.613
R14416 GND.n8893 GND.n8892 280.613
R14417 GND.n8894 GND.n8893 280.613
R14418 GND.n8894 GND.n952 280.613
R14419 GND.n8902 GND.n952 280.613
R14420 GND.n8903 GND.n8902 280.613
R14421 GND.n8904 GND.n8903 280.613
R14422 GND.n8904 GND.n946 280.613
R14423 GND.n8912 GND.n946 280.613
R14424 GND.n8913 GND.n8912 280.613
R14425 GND.n8914 GND.n8913 280.613
R14426 GND.n8914 GND.n940 280.613
R14427 GND.n8922 GND.n940 280.613
R14428 GND.n8923 GND.n8922 280.613
R14429 GND.n8924 GND.n8923 280.613
R14430 GND.n8924 GND.n934 280.613
R14431 GND.n8932 GND.n934 280.613
R14432 GND.n8933 GND.n8932 280.613
R14433 GND.n8934 GND.n8933 280.613
R14434 GND.n8934 GND.n928 280.613
R14435 GND.n8942 GND.n928 280.613
R14436 GND.n8943 GND.n8942 280.613
R14437 GND.n8944 GND.n8943 280.613
R14438 GND.n8944 GND.n922 280.613
R14439 GND.n8952 GND.n922 280.613
R14440 GND.n8953 GND.n8952 280.613
R14441 GND.n8954 GND.n8953 280.613
R14442 GND.n8954 GND.n916 280.613
R14443 GND.n8962 GND.n916 280.613
R14444 GND.n8963 GND.n8962 280.613
R14445 GND.n8964 GND.n8963 280.613
R14446 GND.n8964 GND.n910 280.613
R14447 GND.n8972 GND.n910 280.613
R14448 GND.n8973 GND.n8972 280.613
R14449 GND.n8974 GND.n8973 280.613
R14450 GND.n8974 GND.n904 280.613
R14451 GND.n8982 GND.n904 280.613
R14452 GND.n8983 GND.n8982 280.613
R14453 GND.n8984 GND.n8983 280.613
R14454 GND.n8984 GND.n898 280.613
R14455 GND.n8992 GND.n898 280.613
R14456 GND.n8993 GND.n8992 280.613
R14457 GND.n8994 GND.n8993 280.613
R14458 GND.n8994 GND.n892 280.613
R14459 GND.n9002 GND.n892 280.613
R14460 GND.n9003 GND.n9002 280.613
R14461 GND.n9004 GND.n9003 280.613
R14462 GND.n9004 GND.n886 280.613
R14463 GND.n9012 GND.n886 280.613
R14464 GND.n9013 GND.n9012 280.613
R14465 GND.n9014 GND.n9013 280.613
R14466 GND.n9014 GND.n880 280.613
R14467 GND.n9022 GND.n880 280.613
R14468 GND.n9023 GND.n9022 280.613
R14469 GND.n9024 GND.n9023 280.613
R14470 GND.n9024 GND.n874 280.613
R14471 GND.n9032 GND.n874 280.613
R14472 GND.n9033 GND.n9032 280.613
R14473 GND.n9034 GND.n9033 280.613
R14474 GND.n9034 GND.n868 280.613
R14475 GND.n9042 GND.n868 280.613
R14476 GND.n9043 GND.n9042 280.613
R14477 GND.n9044 GND.n9043 280.613
R14478 GND.n9044 GND.n862 280.613
R14479 GND.n9052 GND.n862 280.613
R14480 GND.n9053 GND.n9052 280.613
R14481 GND.n9054 GND.n9053 280.613
R14482 GND.n9054 GND.n856 280.613
R14483 GND.n9062 GND.n856 280.613
R14484 GND.n9063 GND.n9062 280.613
R14485 GND.n9064 GND.n9063 280.613
R14486 GND.n9064 GND.n850 280.613
R14487 GND.n9072 GND.n850 280.613
R14488 GND.n9073 GND.n9072 280.613
R14489 GND.n9074 GND.n9073 280.613
R14490 GND.n9074 GND.n844 280.613
R14491 GND.n9082 GND.n844 280.613
R14492 GND.n9083 GND.n9082 280.613
R14493 GND.n9084 GND.n9083 280.613
R14494 GND.n9084 GND.n838 280.613
R14495 GND.n9092 GND.n838 280.613
R14496 GND.n9093 GND.n9092 280.613
R14497 GND.n9094 GND.n9093 280.613
R14498 GND.n9094 GND.n832 280.613
R14499 GND.n9102 GND.n832 280.613
R14500 GND.n9103 GND.n9102 280.613
R14501 GND.n9104 GND.n9103 280.613
R14502 GND.n9104 GND.n826 280.613
R14503 GND.n9112 GND.n826 280.613
R14504 GND.n9113 GND.n9112 280.613
R14505 GND.n9114 GND.n9113 280.613
R14506 GND.n9114 GND.n820 280.613
R14507 GND.n9122 GND.n820 280.613
R14508 GND.n9123 GND.n9122 280.613
R14509 GND.n9124 GND.n9123 280.613
R14510 GND.n9124 GND.n814 280.613
R14511 GND.n9132 GND.n814 280.613
R14512 GND.n9133 GND.n9132 280.613
R14513 GND.n9134 GND.n9133 280.613
R14514 GND.n9134 GND.n808 280.613
R14515 GND.n9142 GND.n808 280.613
R14516 GND.n9143 GND.n9142 280.613
R14517 GND.n9144 GND.n9143 280.613
R14518 GND.n9144 GND.n802 280.613
R14519 GND.n9152 GND.n802 280.613
R14520 GND.n9153 GND.n9152 280.613
R14521 GND.n9154 GND.n9153 280.613
R14522 GND.n9154 GND.n796 280.613
R14523 GND.n9162 GND.n796 280.613
R14524 GND.n9163 GND.n9162 280.613
R14525 GND.n9164 GND.n9163 280.613
R14526 GND.n9164 GND.n790 280.613
R14527 GND.n9172 GND.n790 280.613
R14528 GND.n9173 GND.n9172 280.613
R14529 GND.n9174 GND.n9173 280.613
R14530 GND.n9174 GND.n784 280.613
R14531 GND.n9182 GND.n784 280.613
R14532 GND.n9183 GND.n9182 280.613
R14533 GND.n9184 GND.n9183 280.613
R14534 GND.n9184 GND.n778 280.613
R14535 GND.n9192 GND.n778 280.613
R14536 GND.n9193 GND.n9192 280.613
R14537 GND.n9194 GND.n9193 280.613
R14538 GND.n9194 GND.n772 280.613
R14539 GND.n9202 GND.n772 280.613
R14540 GND.n9203 GND.n9202 280.613
R14541 GND.n9204 GND.n9203 280.613
R14542 GND.n9204 GND.n766 280.613
R14543 GND.n9212 GND.n766 280.613
R14544 GND.n9213 GND.n9212 280.613
R14545 GND.n9214 GND.n9213 280.613
R14546 GND.n9214 GND.n760 280.613
R14547 GND.n9222 GND.n760 280.613
R14548 GND.n9223 GND.n9222 280.613
R14549 GND.n9224 GND.n9223 280.613
R14550 GND.n9224 GND.n754 280.613
R14551 GND.n9232 GND.n754 280.613
R14552 GND.n9233 GND.n9232 280.613
R14553 GND.n9234 GND.n9233 280.613
R14554 GND.n9234 GND.n748 280.613
R14555 GND.n9242 GND.n748 280.613
R14556 GND.n9243 GND.n9242 280.613
R14557 GND.n9244 GND.n9243 280.613
R14558 GND.n9244 GND.n742 280.613
R14559 GND.n9252 GND.n742 280.613
R14560 GND.n9253 GND.n9252 280.613
R14561 GND.n9254 GND.n9253 280.613
R14562 GND.n9254 GND.n736 280.613
R14563 GND.n9262 GND.n736 280.613
R14564 GND.n9263 GND.n9262 280.613
R14565 GND.n9264 GND.n9263 280.613
R14566 GND.n9264 GND.n730 280.613
R14567 GND.n9272 GND.n730 280.613
R14568 GND.n9273 GND.n9272 280.613
R14569 GND.n9274 GND.n9273 280.613
R14570 GND.n9274 GND.n724 280.613
R14571 GND.n9282 GND.n724 280.613
R14572 GND.n9283 GND.n9282 280.613
R14573 GND.n9284 GND.n9283 280.613
R14574 GND.n9284 GND.n718 280.613
R14575 GND.n9292 GND.n718 280.613
R14576 GND.n9293 GND.n9292 280.613
R14577 GND.n9294 GND.n9293 280.613
R14578 GND.n9294 GND.n712 280.613
R14579 GND.n9302 GND.n712 280.613
R14580 GND.n9303 GND.n9302 280.613
R14581 GND.n9304 GND.n9303 280.613
R14582 GND.n9304 GND.n706 280.613
R14583 GND.n9312 GND.n706 280.613
R14584 GND.n9313 GND.n9312 280.613
R14585 GND.n9314 GND.n9313 280.613
R14586 GND.n9314 GND.n700 280.613
R14587 GND.n9322 GND.n700 280.613
R14588 GND.n9544 GND.t115 262.012
R14589 GND.n497 GND.t148 262.012
R14590 GND.n516 GND.t129 262.012
R14591 GND.n1791 GND.t95 262.012
R14592 GND.n1811 GND.t132 262.012
R14593 GND.n1879 GND.t85 262.012
R14594 GND.n2377 GND.t112 262.012
R14595 GND.n6290 GND.t161 262.012
R14596 GND.n6108 GND.t106 262.012
R14597 GND.n1487 GND.t103 262.012
R14598 GND.n1501 GND.t152 262.012
R14599 GND.n3346 GND.t93 262.012
R14600 GND.n4705 GND.t109 260.649
R14601 GND.n6206 GND.t143 260.649
R14602 GND.n4722 GND.n2955 256.663
R14603 GND.n4728 GND.n2955 256.663
R14604 GND.n4730 GND.n2955 256.663
R14605 GND.n4736 GND.n2955 256.663
R14606 GND.n4738 GND.n2955 256.663
R14607 GND.n4744 GND.n2955 256.663
R14608 GND.n4746 GND.n2955 256.663
R14609 GND.n4752 GND.n2955 256.663
R14610 GND.n4754 GND.n2955 256.663
R14611 GND.n4761 GND.n2955 256.663
R14612 GND.n4764 GND.n2955 256.663
R14613 GND.n4765 GND.n1795 256.663
R14614 GND.n4766 GND.n2955 256.663
R14615 GND.n4768 GND.n2955 256.663
R14616 GND.n4775 GND.n2955 256.663
R14617 GND.n4777 GND.n2955 256.663
R14618 GND.n4783 GND.n2955 256.663
R14619 GND.n4785 GND.n2955 256.663
R14620 GND.n4791 GND.n2955 256.663
R14621 GND.n4793 GND.n2955 256.663
R14622 GND.n4799 GND.n2955 256.663
R14623 GND.n4801 GND.n2955 256.663
R14624 GND.n4807 GND.n2955 256.663
R14625 GND.n6257 GND.n6125 256.663
R14626 GND.n6257 GND.n6126 256.663
R14627 GND.n6257 GND.n6127 256.663
R14628 GND.n6257 GND.n6128 256.663
R14629 GND.n6257 GND.n6129 256.663
R14630 GND.n6257 GND.n6130 256.663
R14631 GND.n6257 GND.n6131 256.663
R14632 GND.n6257 GND.n6132 256.663
R14633 GND.n6257 GND.n6133 256.663
R14634 GND.n6257 GND.n6134 256.663
R14635 GND.n6257 GND.n6183 256.663
R14636 GND.n6260 GND.n6122 256.663
R14637 GND.n6258 GND.n6257 256.663
R14638 GND.n6257 GND.n6184 256.663
R14639 GND.n6257 GND.n6185 256.663
R14640 GND.n6257 GND.n6186 256.663
R14641 GND.n6257 GND.n6187 256.663
R14642 GND.n6257 GND.n6188 256.663
R14643 GND.n6257 GND.n6189 256.663
R14644 GND.n6257 GND.n6190 256.663
R14645 GND.n6257 GND.n6191 256.663
R14646 GND.n6257 GND.n6192 256.663
R14647 GND.n6257 GND.n6193 256.663
R14648 GND.n4684 GND.t137 254.942
R14649 GND.n6135 GND.t126 254.942
R14650 GND.n4689 GND.t146 254.942
R14651 GND.n6215 GND.t139 254.942
R14652 GND.n7867 GND.n7866 242.672
R14653 GND.n7866 GND.n1840 242.672
R14654 GND.n7866 GND.n1841 242.672
R14655 GND.n7866 GND.n1842 242.672
R14656 GND.n7866 GND.n1843 242.672
R14657 GND.n7866 GND.n1844 242.672
R14658 GND.n7866 GND.n1845 242.672
R14659 GND.n7866 GND.n1846 242.672
R14660 GND.n7866 GND.n1847 242.672
R14661 GND.n6416 GND.n6415 242.672
R14662 GND.n6415 GND.n6414 242.672
R14663 GND.n6415 GND.n6413 242.672
R14664 GND.n6415 GND.n6412 242.672
R14665 GND.n6415 GND.n6410 242.672
R14666 GND.n6415 GND.n6409 242.672
R14667 GND.n6415 GND.n6407 242.672
R14668 GND.n6415 GND.n6405 242.672
R14669 GND.n6415 GND.n6404 242.672
R14670 GND.n6415 GND.n6402 242.672
R14671 GND.n8151 GND.n1471 242.672
R14672 GND.n8151 GND.n1470 242.672
R14673 GND.n8151 GND.n1469 242.672
R14674 GND.n8151 GND.n1468 242.672
R14675 GND.n8151 GND.n1467 242.672
R14676 GND.n8151 GND.n1466 242.672
R14677 GND.n7881 GND.n1826 242.672
R14678 GND.n7881 GND.n1827 242.672
R14679 GND.n7881 GND.n1828 242.672
R14680 GND.n7881 GND.n1829 242.672
R14681 GND.n7881 GND.n1830 242.672
R14682 GND.n7881 GND.n1831 242.672
R14683 GND.n8151 GND.n8150 242.672
R14684 GND.n8151 GND.n1452 242.672
R14685 GND.n8151 GND.n1453 242.672
R14686 GND.n8151 GND.n1454 242.672
R14687 GND.n8151 GND.n1455 242.672
R14688 GND.n8151 GND.n1456 242.672
R14689 GND.n8151 GND.n1457 242.672
R14690 GND.n8151 GND.n1458 242.672
R14691 GND.n8151 GND.n1459 242.672
R14692 GND.n8151 GND.n1460 242.672
R14693 GND.n8151 GND.n1461 242.672
R14694 GND.n8151 GND.n1462 242.672
R14695 GND.n7882 GND.n7881 242.672
R14696 GND.n7881 GND.n1824 242.672
R14697 GND.n7881 GND.n1823 242.672
R14698 GND.n7881 GND.n1821 242.672
R14699 GND.n7881 GND.n1820 242.672
R14700 GND.n7881 GND.n1818 242.672
R14701 GND.n7881 GND.n1817 242.672
R14702 GND.n7905 GND.n1794 242.672
R14703 GND.n7881 GND.n7874 242.672
R14704 GND.n7881 GND.n7876 242.672
R14705 GND.n7881 GND.n7877 242.672
R14706 GND.n7881 GND.n7879 242.672
R14707 GND.n7881 GND.n7880 242.672
R14708 GND.n7293 GND.n3292 242.672
R14709 GND.n7293 GND.n3293 242.672
R14710 GND.n7293 GND.n3294 242.672
R14711 GND.n7293 GND.n3295 242.672
R14712 GND.n7293 GND.n3296 242.672
R14713 GND.n6292 GND.n6261 242.672
R14714 GND.n7293 GND.n3298 242.672
R14715 GND.n7293 GND.n3299 242.672
R14716 GND.n7293 GND.n3300 242.672
R14717 GND.n7293 GND.n3301 242.672
R14718 GND.n7293 GND.n3302 242.672
R14719 GND.n7293 GND.n3303 242.672
R14720 GND.n7293 GND.n3304 242.672
R14721 GND.n9568 GND.n9567 242.672
R14722 GND.n9567 GND.n537 242.672
R14723 GND.n9567 GND.n535 242.672
R14724 GND.n9567 GND.n534 242.672
R14725 GND.n9567 GND.n532 242.672
R14726 GND.n9567 GND.n531 242.672
R14727 GND.n9567 GND.n529 242.672
R14728 GND.n9567 GND.n528 242.672
R14729 GND.n9567 GND.n526 242.672
R14730 GND.n9567 GND.n525 242.672
R14731 GND.n9567 GND.n523 242.672
R14732 GND.n9567 GND.n522 242.672
R14733 GND.n9567 GND.n520 242.672
R14734 GND.n7293 GND.n3306 242.672
R14735 GND.n7293 GND.n3307 242.672
R14736 GND.n7293 GND.n3308 242.672
R14737 GND.n7293 GND.n3309 242.672
R14738 GND.n7293 GND.n3310 242.672
R14739 GND.n7293 GND.n3311 242.672
R14740 GND.n9567 GND.n543 242.672
R14741 GND.n9567 GND.n542 242.672
R14742 GND.n9567 GND.n541 242.672
R14743 GND.n9567 GND.n540 242.672
R14744 GND.n9567 GND.n539 242.672
R14745 GND.n9567 GND.n538 242.672
R14746 GND.n486 GND.n485 240.244
R14747 GND.n521 GND.n489 240.244
R14748 GND.n491 GND.n490 240.244
R14749 GND.n524 GND.n494 240.244
R14750 GND.n496 GND.n495 240.244
R14751 GND.n527 GND.n501 240.244
R14752 GND.n503 GND.n502 240.244
R14753 GND.n530 GND.n506 240.244
R14754 GND.n508 GND.n507 240.244
R14755 GND.n533 GND.n511 240.244
R14756 GND.n513 GND.n512 240.244
R14757 GND.n536 GND.n518 240.244
R14758 GND.n3377 GND.n3357 240.244
R14759 GND.n3377 GND.n3367 240.244
R14760 GND.n3379 GND.n3367 240.244
R14761 GND.n3380 GND.n3379 240.244
R14762 GND.n3959 GND.n3380 240.244
R14763 GND.n3959 GND.n3386 240.244
R14764 GND.n3387 GND.n3386 240.244
R14765 GND.n3388 GND.n3387 240.244
R14766 GND.n6605 GND.n3388 240.244
R14767 GND.n6605 GND.n3394 240.244
R14768 GND.n3395 GND.n3394 240.244
R14769 GND.n3396 GND.n3395 240.244
R14770 GND.n3925 GND.n3396 240.244
R14771 GND.n3925 GND.n3402 240.244
R14772 GND.n3403 GND.n3402 240.244
R14773 GND.n3404 GND.n3403 240.244
R14774 GND.n3906 GND.n3404 240.244
R14775 GND.n3906 GND.n3410 240.244
R14776 GND.n3411 GND.n3410 240.244
R14777 GND.n3412 GND.n3411 240.244
R14778 GND.n3894 GND.n3412 240.244
R14779 GND.n3894 GND.n3418 240.244
R14780 GND.n3419 GND.n3418 240.244
R14781 GND.n3420 GND.n3419 240.244
R14782 GND.n3869 GND.n3420 240.244
R14783 GND.n3869 GND.n3426 240.244
R14784 GND.n3427 GND.n3426 240.244
R14785 GND.n3428 GND.n3427 240.244
R14786 GND.n6704 GND.n3428 240.244
R14787 GND.n6704 GND.n3434 240.244
R14788 GND.n3435 GND.n3434 240.244
R14789 GND.n3436 GND.n3435 240.244
R14790 GND.n3834 GND.n3436 240.244
R14791 GND.n3834 GND.n3442 240.244
R14792 GND.n3443 GND.n3442 240.244
R14793 GND.n3444 GND.n3443 240.244
R14794 GND.n3815 GND.n3444 240.244
R14795 GND.n3815 GND.n3450 240.244
R14796 GND.n3451 GND.n3450 240.244
R14797 GND.n3452 GND.n3451 240.244
R14798 GND.n3803 GND.n3452 240.244
R14799 GND.n3803 GND.n3458 240.244
R14800 GND.n3459 GND.n3458 240.244
R14801 GND.n3460 GND.n3459 240.244
R14802 GND.n3774 GND.n3460 240.244
R14803 GND.n3774 GND.n3466 240.244
R14804 GND.n3467 GND.n3466 240.244
R14805 GND.n3468 GND.n3467 240.244
R14806 GND.n6801 GND.n3468 240.244
R14807 GND.n6801 GND.n3474 240.244
R14808 GND.n3475 GND.n3474 240.244
R14809 GND.n3476 GND.n3475 240.244
R14810 GND.n6817 GND.n3476 240.244
R14811 GND.n6817 GND.n3482 240.244
R14812 GND.n3483 GND.n3482 240.244
R14813 GND.n3484 GND.n3483 240.244
R14814 GND.n6832 GND.n3484 240.244
R14815 GND.n6832 GND.n3490 240.244
R14816 GND.n3491 GND.n3490 240.244
R14817 GND.n3492 GND.n3491 240.244
R14818 GND.n3720 GND.n3492 240.244
R14819 GND.n3720 GND.n3498 240.244
R14820 GND.n3499 GND.n3498 240.244
R14821 GND.n3500 GND.n3499 240.244
R14822 GND.n3709 GND.n3500 240.244
R14823 GND.n3709 GND.n3506 240.244
R14824 GND.n3507 GND.n3506 240.244
R14825 GND.n3508 GND.n3507 240.244
R14826 GND.n6941 GND.n3508 240.244
R14827 GND.n6941 GND.n3514 240.244
R14828 GND.n3515 GND.n3514 240.244
R14829 GND.n3516 GND.n3515 240.244
R14830 GND.n3670 GND.n3516 240.244
R14831 GND.n3670 GND.n3522 240.244
R14832 GND.n3523 GND.n3522 240.244
R14833 GND.n3524 GND.n3523 240.244
R14834 GND.n3658 GND.n3524 240.244
R14835 GND.n3658 GND.n3530 240.244
R14836 GND.n3531 GND.n3530 240.244
R14837 GND.n3532 GND.n3531 240.244
R14838 GND.n3634 GND.n3532 240.244
R14839 GND.n3634 GND.n3538 240.244
R14840 GND.n3539 GND.n3538 240.244
R14841 GND.n3540 GND.n3539 240.244
R14842 GND.n3623 GND.n3540 240.244
R14843 GND.n3623 GND.n3546 240.244
R14844 GND.n3547 GND.n3546 240.244
R14845 GND.n3548 GND.n3547 240.244
R14846 GND.n7050 GND.n3548 240.244
R14847 GND.n7050 GND.n3554 240.244
R14848 GND.n3555 GND.n3554 240.244
R14849 GND.n3556 GND.n3555 240.244
R14850 GND.n3583 GND.n3556 240.244
R14851 GND.n3583 GND.n3562 240.244
R14852 GND.n3563 GND.n3562 240.244
R14853 GND.n3564 GND.n3563 240.244
R14854 GND.n3570 GND.n3564 240.244
R14855 GND.n3570 GND.n578 240.244
R14856 GND.n9500 GND.n578 240.244
R14857 GND.n9500 GND.n568 240.244
R14858 GND.n568 GND.n556 240.244
R14859 GND.n9517 GND.n556 240.244
R14860 GND.n9517 GND.n550 240.244
R14861 GND.n9525 GND.n550 240.244
R14862 GND.n9525 GND.n477 240.244
R14863 GND.n6271 GND.n6270 240.244
R14864 GND.n6275 GND.n6274 240.244
R14865 GND.n6281 GND.n6280 240.244
R14866 GND.n6285 GND.n6284 240.244
R14867 GND.n6118 GND.n3297 240.244
R14868 GND.n6295 GND.n6294 240.244
R14869 GND.n6301 GND.n6300 240.244
R14870 GND.n6305 GND.n6304 240.244
R14871 GND.n6311 GND.n6310 240.244
R14872 GND.n6315 GND.n6314 240.244
R14873 GND.n6112 GND.n6111 240.244
R14874 GND.n6107 GND.n3305 240.244
R14875 GND.n7255 GND.n3360 240.244
R14876 GND.n7251 GND.n3360 240.244
R14877 GND.n7251 GND.n3365 240.244
R14878 GND.n6583 GND.n3365 240.244
R14879 GND.n6593 GND.n6583 240.244
R14880 GND.n6593 GND.n6585 240.244
R14881 GND.n6585 GND.n3946 240.244
R14882 GND.n6610 GND.n3946 240.244
R14883 GND.n6610 GND.n3940 240.244
R14884 GND.n6618 GND.n3940 240.244
R14885 GND.n6618 GND.n3942 240.244
R14886 GND.n3942 GND.n3923 240.244
R14887 GND.n6634 GND.n3923 240.244
R14888 GND.n6634 GND.n3917 240.244
R14889 GND.n6642 GND.n3917 240.244
R14890 GND.n6642 GND.n3919 240.244
R14891 GND.n3919 GND.n3900 240.244
R14892 GND.n6659 GND.n3900 240.244
R14893 GND.n6659 GND.n3893 240.244
R14894 GND.n6667 GND.n3893 240.244
R14895 GND.n6667 GND.n3896 240.244
R14896 GND.n3896 GND.n3878 240.244
R14897 GND.n6684 GND.n3878 240.244
R14898 GND.n6684 GND.n3872 240.244
R14899 GND.n6692 GND.n3872 240.244
R14900 GND.n6692 GND.n3874 240.244
R14901 GND.n3874 GND.n3855 240.244
R14902 GND.n6709 GND.n3855 240.244
R14903 GND.n6709 GND.n3849 240.244
R14904 GND.n6717 GND.n3849 240.244
R14905 GND.n6717 GND.n3851 240.244
R14906 GND.n3851 GND.n3832 240.244
R14907 GND.n6733 GND.n3832 240.244
R14908 GND.n6733 GND.n3826 240.244
R14909 GND.n6741 GND.n3826 240.244
R14910 GND.n6741 GND.n3828 240.244
R14911 GND.n3828 GND.n3809 240.244
R14912 GND.n6758 GND.n3809 240.244
R14913 GND.n6758 GND.n3802 240.244
R14914 GND.n6766 GND.n3802 240.244
R14915 GND.n6766 GND.n3805 240.244
R14916 GND.n3805 GND.n3787 240.244
R14917 GND.n6783 GND.n3787 240.244
R14918 GND.n6783 GND.n3777 240.244
R14919 GND.n6792 GND.n3777 240.244
R14920 GND.n6792 GND.n3783 240.244
R14921 GND.n3783 GND.n3754 240.244
R14922 GND.n6876 GND.n3754 240.244
R14923 GND.n6876 GND.n3755 240.244
R14924 GND.n6871 GND.n3755 240.244
R14925 GND.n6871 GND.n3758 240.244
R14926 GND.n6820 GND.n3758 240.244
R14927 GND.n6859 GND.n6820 240.244
R14928 GND.n6859 GND.n6821 240.244
R14929 GND.n6854 GND.n6821 240.244
R14930 GND.n6854 GND.n6825 240.244
R14931 GND.n6839 GND.n6825 240.244
R14932 GND.n6839 GND.n6834 240.244
R14933 GND.n6834 GND.n3729 240.244
R14934 GND.n6893 GND.n3729 240.244
R14935 GND.n6893 GND.n3724 240.244
R14936 GND.n6901 GND.n3724 240.244
R14937 GND.n6901 GND.n3725 240.244
R14938 GND.n3725 GND.n3707 240.244
R14939 GND.n6920 GND.n3707 240.244
R14940 GND.n6920 GND.n3702 240.244
R14941 GND.n6928 GND.n3702 240.244
R14942 GND.n6928 GND.n3703 240.244
R14943 GND.n3703 GND.n3686 240.244
R14944 GND.n6949 GND.n3686 240.244
R14945 GND.n6949 GND.n3681 240.244
R14946 GND.n6957 GND.n3681 240.244
R14947 GND.n6957 GND.n3682 240.244
R14948 GND.n3682 GND.n3666 240.244
R14949 GND.n6976 GND.n3666 240.244
R14950 GND.n6976 GND.n3661 240.244
R14951 GND.n6984 GND.n3661 240.244
R14952 GND.n6984 GND.n3662 240.244
R14953 GND.n3662 GND.n3643 240.244
R14954 GND.n7002 GND.n3643 240.244
R14955 GND.n7002 GND.n3638 240.244
R14956 GND.n7010 GND.n3638 240.244
R14957 GND.n7010 GND.n3639 240.244
R14958 GND.n3639 GND.n3621 240.244
R14959 GND.n7029 GND.n3621 240.244
R14960 GND.n7029 GND.n3616 240.244
R14961 GND.n7037 GND.n3616 240.244
R14962 GND.n7037 GND.n3617 240.244
R14963 GND.n3617 GND.n3600 240.244
R14964 GND.n7057 GND.n3600 240.244
R14965 GND.n7057 GND.n3595 240.244
R14966 GND.n7065 GND.n3595 240.244
R14967 GND.n7065 GND.n3596 240.244
R14968 GND.n3596 GND.n3577 240.244
R14969 GND.n7090 GND.n3577 240.244
R14970 GND.n7090 GND.n3572 240.244
R14971 GND.n7098 GND.n3572 240.244
R14972 GND.n7098 GND.n3573 240.244
R14973 GND.n3573 GND.n566 240.244
R14974 GND.n9507 GND.n566 240.244
R14975 GND.n9507 GND.n560 240.244
R14976 GND.n9515 GND.n560 240.244
R14977 GND.n9515 GND.n562 240.244
R14978 GND.n562 GND.n480 240.244
R14979 GND.n9611 GND.n480 240.244
R14980 GND.n1780 GND.n1776 240.244
R14981 GND.n7878 GND.n1781 240.244
R14982 GND.n1785 GND.n1784 240.244
R14983 GND.n7875 GND.n1786 240.244
R14984 GND.n1790 GND.n1789 240.244
R14985 GND.n1815 GND.n1796 240.244
R14986 GND.n1816 GND.n1799 240.244
R14987 GND.n1801 GND.n1800 240.244
R14988 GND.n1819 GND.n1804 240.244
R14989 GND.n1806 GND.n1805 240.244
R14990 GND.n1822 GND.n1809 240.244
R14991 GND.n7883 GND.n1810 240.244
R14992 GND.n1560 GND.n1510 240.244
R14993 GND.n1560 GND.n1559 240.244
R14994 GND.n1559 GND.n1528 240.244
R14995 GND.n2369 GND.n1528 240.244
R14996 GND.n2369 GND.n1547 240.244
R14997 GND.n1570 GND.n1547 240.244
R14998 GND.n1571 GND.n1570 240.244
R14999 GND.n2505 GND.n1571 240.244
R15000 GND.n2505 GND.n1577 240.244
R15001 GND.n1578 GND.n1577 240.244
R15002 GND.n1579 GND.n1578 240.244
R15003 GND.n2350 GND.n1579 240.244
R15004 GND.n2350 GND.n1585 240.244
R15005 GND.n1586 GND.n1585 240.244
R15006 GND.n1587 GND.n1586 240.244
R15007 GND.n2550 GND.n1587 240.244
R15008 GND.n2550 GND.n1593 240.244
R15009 GND.n1594 GND.n1593 240.244
R15010 GND.n1595 GND.n1594 240.244
R15011 GND.n2315 GND.n1595 240.244
R15012 GND.n2315 GND.n1601 240.244
R15013 GND.n1602 GND.n1601 240.244
R15014 GND.n1603 GND.n1602 240.244
R15015 GND.n2296 GND.n1603 240.244
R15016 GND.n2296 GND.n1609 240.244
R15017 GND.n1610 GND.n1609 240.244
R15018 GND.n1611 GND.n1610 240.244
R15019 GND.n2284 GND.n1611 240.244
R15020 GND.n2284 GND.n1617 240.244
R15021 GND.n1618 GND.n1617 240.244
R15022 GND.n1619 GND.n1618 240.244
R15023 GND.n2262 GND.n1619 240.244
R15024 GND.n2262 GND.n1625 240.244
R15025 GND.n1626 GND.n1625 240.244
R15026 GND.n1627 GND.n1626 240.244
R15027 GND.n2240 GND.n1627 240.244
R15028 GND.n2240 GND.n1633 240.244
R15029 GND.n1634 GND.n1633 240.244
R15030 GND.n1635 GND.n1634 240.244
R15031 GND.n2724 GND.n1635 240.244
R15032 GND.n2724 GND.n1641 240.244
R15033 GND.n1642 GND.n1641 240.244
R15034 GND.n1643 GND.n1642 240.244
R15035 GND.n2205 GND.n1643 240.244
R15036 GND.n2205 GND.n1649 240.244
R15037 GND.n1650 GND.n1649 240.244
R15038 GND.n1651 GND.n1650 240.244
R15039 GND.n2117 GND.n1651 240.244
R15040 GND.n2117 GND.n1657 240.244
R15041 GND.n1658 GND.n1657 240.244
R15042 GND.n1659 GND.n1658 240.244
R15043 GND.n2132 GND.n1659 240.244
R15044 GND.n2132 GND.n1665 240.244
R15045 GND.n1666 GND.n1665 240.244
R15046 GND.n1667 GND.n1666 240.244
R15047 GND.n2185 GND.n1667 240.244
R15048 GND.n2185 GND.n1673 240.244
R15049 GND.n1674 GND.n1673 240.244
R15050 GND.n1675 GND.n1674 240.244
R15051 GND.n2091 GND.n1675 240.244
R15052 GND.n2091 GND.n1681 240.244
R15053 GND.n1682 GND.n1681 240.244
R15054 GND.n1683 GND.n1682 240.244
R15055 GND.n2079 GND.n1683 240.244
R15056 GND.n2079 GND.n1689 240.244
R15057 GND.n1690 GND.n1689 240.244
R15058 GND.n1691 GND.n1690 240.244
R15059 GND.n2054 GND.n1691 240.244
R15060 GND.n2054 GND.n1697 240.244
R15061 GND.n1698 GND.n1697 240.244
R15062 GND.n1699 GND.n1698 240.244
R15063 GND.n7664 GND.n1699 240.244
R15064 GND.n7664 GND.n1705 240.244
R15065 GND.n1706 GND.n1705 240.244
R15066 GND.n1707 GND.n1706 240.244
R15067 GND.n2014 GND.n1707 240.244
R15068 GND.n2014 GND.n1713 240.244
R15069 GND.n1714 GND.n1713 240.244
R15070 GND.n1715 GND.n1714 240.244
R15071 GND.n1995 GND.n1715 240.244
R15072 GND.n1995 GND.n1721 240.244
R15073 GND.n1722 GND.n1721 240.244
R15074 GND.n1723 GND.n1722 240.244
R15075 GND.n1983 GND.n1723 240.244
R15076 GND.n1983 GND.n1729 240.244
R15077 GND.n1730 GND.n1729 240.244
R15078 GND.n1731 GND.n1730 240.244
R15079 GND.n1958 GND.n1731 240.244
R15080 GND.n1958 GND.n1737 240.244
R15081 GND.n1738 GND.n1737 240.244
R15082 GND.n1739 GND.n1738 240.244
R15083 GND.n7763 GND.n1739 240.244
R15084 GND.n7763 GND.n1745 240.244
R15085 GND.n1746 GND.n1745 240.244
R15086 GND.n1747 GND.n1746 240.244
R15087 GND.n1923 GND.n1747 240.244
R15088 GND.n1923 GND.n1753 240.244
R15089 GND.n1754 GND.n1753 240.244
R15090 GND.n1755 GND.n1754 240.244
R15091 GND.n1905 GND.n1755 240.244
R15092 GND.n1905 GND.n1761 240.244
R15093 GND.n1762 GND.n1761 240.244
R15094 GND.n1763 GND.n1762 240.244
R15095 GND.n1769 GND.n1763 240.244
R15096 GND.n7925 GND.n1769 240.244
R15097 GND.n1473 GND.n1472 240.244
R15098 GND.n8144 GND.n1472 240.244
R15099 GND.n8142 GND.n8141 240.244
R15100 GND.n8138 GND.n8137 240.244
R15101 GND.n8134 GND.n8133 240.244
R15102 GND.n8130 GND.n8129 240.244
R15103 GND.n8126 GND.n8125 240.244
R15104 GND.n8122 GND.n8121 240.244
R15105 GND.n8118 GND.n8117 240.244
R15106 GND.n8114 GND.n8113 240.244
R15107 GND.n8110 GND.n8109 240.244
R15108 GND.n8106 GND.n8105 240.244
R15109 GND.n1500 GND.n1463 240.244
R15110 GND.n1537 GND.n1474 240.244
R15111 GND.n1537 GND.n1532 240.244
R15112 GND.n8085 GND.n1532 240.244
R15113 GND.n8085 GND.n1533 240.244
R15114 GND.n8081 GND.n1533 240.244
R15115 GND.n8081 GND.n1545 240.244
R15116 GND.n2513 GND.n1545 240.244
R15117 GND.n2513 GND.n2507 240.244
R15118 GND.n2507 GND.n2359 240.244
R15119 GND.n2530 GND.n2359 240.244
R15120 GND.n2530 GND.n2353 240.244
R15121 GND.n2538 GND.n2353 240.244
R15122 GND.n2538 GND.n2355 240.244
R15123 GND.n2355 GND.n2336 240.244
R15124 GND.n2555 GND.n2336 240.244
R15125 GND.n2555 GND.n2330 240.244
R15126 GND.n2563 GND.n2330 240.244
R15127 GND.n2563 GND.n2332 240.244
R15128 GND.n2332 GND.n2313 240.244
R15129 GND.n2579 GND.n2313 240.244
R15130 GND.n2579 GND.n2307 240.244
R15131 GND.n2587 GND.n2307 240.244
R15132 GND.n2587 GND.n2309 240.244
R15133 GND.n2309 GND.n2290 240.244
R15134 GND.n2604 GND.n2290 240.244
R15135 GND.n2604 GND.n2283 240.244
R15136 GND.n2612 GND.n2283 240.244
R15137 GND.n2612 GND.n2286 240.244
R15138 GND.n2286 GND.n2268 240.244
R15139 GND.n2637 GND.n2268 240.244
R15140 GND.n2637 GND.n2264 240.244
R15141 GND.n2643 GND.n2264 240.244
R15142 GND.n2643 GND.n2249 240.244
R15143 GND.n2704 GND.n2249 240.244
R15144 GND.n2704 GND.n2243 240.244
R15145 GND.n2712 GND.n2243 240.244
R15146 GND.n2712 GND.n2245 240.244
R15147 GND.n2245 GND.n2226 240.244
R15148 GND.n2729 GND.n2226 240.244
R15149 GND.n2729 GND.n2220 240.244
R15150 GND.n2737 GND.n2220 240.244
R15151 GND.n2737 GND.n2222 240.244
R15152 GND.n2222 GND.n2203 240.244
R15153 GND.n2753 GND.n2203 240.244
R15154 GND.n2753 GND.n2199 240.244
R15155 GND.n2759 GND.n2199 240.244
R15156 GND.n2759 GND.n2114 240.244
R15157 GND.n2821 GND.n2114 240.244
R15158 GND.n2821 GND.n2115 240.244
R15159 GND.n2137 GND.n2115 240.244
R15160 GND.n2139 GND.n2137 240.244
R15161 GND.n2807 GND.n2139 240.244
R15162 GND.n2807 GND.n2804 240.244
R15163 GND.n2804 GND.n2140 240.244
R15164 GND.n2785 GND.n2140 240.244
R15165 GND.n2787 GND.n2785 240.244
R15166 GND.n2787 GND.n2102 240.244
R15167 GND.n2829 GND.n2102 240.244
R15168 GND.n2829 GND.n2104 240.244
R15169 GND.n2104 GND.n2085 240.244
R15170 GND.n2846 GND.n2085 240.244
R15171 GND.n2846 GND.n2078 240.244
R15172 GND.n2854 GND.n2078 240.244
R15173 GND.n2854 GND.n2081 240.244
R15174 GND.n2081 GND.n2063 240.244
R15175 GND.n2871 GND.n2063 240.244
R15176 GND.n2871 GND.n2058 240.244
R15177 GND.n2879 GND.n2058 240.244
R15178 GND.n2879 GND.n2059 240.244
R15179 GND.n2059 GND.n2035 240.244
R15180 GND.n7669 GND.n2035 240.244
R15181 GND.n7669 GND.n2029 240.244
R15182 GND.n7677 GND.n2029 240.244
R15183 GND.n7677 GND.n2031 240.244
R15184 GND.n2031 GND.n2012 240.244
R15185 GND.n7693 GND.n2012 240.244
R15186 GND.n7693 GND.n2006 240.244
R15187 GND.n7701 GND.n2006 240.244
R15188 GND.n7701 GND.n2008 240.244
R15189 GND.n2008 GND.n1989 240.244
R15190 GND.n7718 GND.n1989 240.244
R15191 GND.n7718 GND.n1982 240.244
R15192 GND.n7726 GND.n1982 240.244
R15193 GND.n7726 GND.n1985 240.244
R15194 GND.n1985 GND.n1967 240.244
R15195 GND.n7743 GND.n1967 240.244
R15196 GND.n7743 GND.n1961 240.244
R15197 GND.n7751 GND.n1961 240.244
R15198 GND.n7751 GND.n1963 240.244
R15199 GND.n1963 GND.n1944 240.244
R15200 GND.n7768 GND.n1944 240.244
R15201 GND.n7768 GND.n1938 240.244
R15202 GND.n7776 GND.n1938 240.244
R15203 GND.n7776 GND.n1940 240.244
R15204 GND.n1940 GND.n1921 240.244
R15205 GND.n7792 GND.n1921 240.244
R15206 GND.n7792 GND.n1915 240.244
R15207 GND.n7800 GND.n1915 240.244
R15208 GND.n7800 GND.n1917 240.244
R15209 GND.n1917 GND.n1899 240.244
R15210 GND.n7819 GND.n1899 240.244
R15211 GND.n7819 GND.n1895 240.244
R15212 GND.n7825 GND.n1895 240.244
R15213 GND.n7825 GND.n1775 240.244
R15214 GND.n7923 GND.n1775 240.244
R15215 GND.n7873 GND.n1832 240.244
R15216 GND.n1857 GND.n1856 240.244
R15217 GND.n1859 GND.n1858 240.244
R15218 GND.n1867 GND.n1866 240.244
R15219 GND.n1877 GND.n1876 240.244
R15220 GND.n1881 GND.n1878 240.244
R15221 GND.n2413 GND.n1511 240.244
R15222 GND.n2414 GND.n2413 240.244
R15223 GND.n2414 GND.n1529 240.244
R15224 GND.n2371 GND.n1529 240.244
R15225 GND.n2371 GND.n1548 240.244
R15226 GND.n2422 GND.n1548 240.244
R15227 GND.n2515 GND.n2422 240.244
R15228 GND.n2515 GND.n2365 240.244
R15229 GND.n2522 GND.n2365 240.244
R15230 GND.n2522 GND.n2361 240.244
R15231 GND.n2361 GND.n2348 240.244
R15232 GND.n2540 GND.n2348 240.244
R15233 GND.n2540 GND.n2343 240.244
R15234 GND.n2547 GND.n2343 240.244
R15235 GND.n2547 GND.n2338 240.244
R15236 GND.n2338 GND.n2326 240.244
R15237 GND.n2565 GND.n2326 240.244
R15238 GND.n2565 GND.n2321 240.244
R15239 GND.n2572 GND.n2321 240.244
R15240 GND.n2572 GND.n2316 240.244
R15241 GND.n2316 GND.n2302 240.244
R15242 GND.n2589 GND.n2302 240.244
R15243 GND.n2589 GND.n2297 240.244
R15244 GND.n2596 GND.n2297 240.244
R15245 GND.n2596 GND.n2292 240.244
R15246 GND.n2292 GND.n2279 240.244
R15247 GND.n2614 GND.n2279 240.244
R15248 GND.n2614 GND.n2274 240.244
R15249 GND.n2630 GND.n2274 240.244
R15250 GND.n2630 GND.n2270 240.244
R15251 GND.n2619 GND.n2270 240.244
R15252 GND.n2619 GND.n2263 240.244
R15253 GND.n2263 GND.n2254 240.244
R15254 GND.n2254 GND.n2250 240.244
R15255 GND.n2250 GND.n2238 240.244
R15256 GND.n2714 GND.n2238 240.244
R15257 GND.n2714 GND.n2233 240.244
R15258 GND.n2721 GND.n2233 240.244
R15259 GND.n2721 GND.n2228 240.244
R15260 GND.n2228 GND.n2216 240.244
R15261 GND.n2739 GND.n2216 240.244
R15262 GND.n2739 GND.n2211 240.244
R15263 GND.n2746 GND.n2211 240.244
R15264 GND.n2746 GND.n2206 240.244
R15265 GND.n2206 GND.n2194 240.244
R15266 GND.n2761 GND.n2194 240.244
R15267 GND.n2761 GND.n2195 240.244
R15268 GND.n2195 GND.n2118 240.244
R15269 GND.n2123 GND.n2118 240.244
R15270 GND.n2769 GND.n2123 240.244
R15271 GND.n2769 GND.n2768 240.244
R15272 GND.n2768 GND.n2133 240.244
R15273 GND.n2141 GND.n2133 240.244
R15274 GND.n2145 GND.n2141 240.244
R15275 GND.n2186 GND.n2145 240.244
R15276 GND.n2782 GND.n2186 240.244
R15277 GND.n2782 GND.n2097 240.244
R15278 GND.n2831 GND.n2097 240.244
R15279 GND.n2831 GND.n2092 240.244
R15280 GND.n2838 GND.n2092 240.244
R15281 GND.n2838 GND.n2087 240.244
R15282 GND.n2087 GND.n2074 240.244
R15283 GND.n2856 GND.n2074 240.244
R15284 GND.n2856 GND.n2069 240.244
R15285 GND.n2863 GND.n2069 240.244
R15286 GND.n2863 GND.n2065 240.244
R15287 GND.n2065 GND.n2052 240.244
R15288 GND.n2881 GND.n2052 240.244
R15289 GND.n2881 GND.n2047 240.244
R15290 GND.n2888 GND.n2047 240.244
R15291 GND.n2888 GND.n2037 240.244
R15292 GND.n2037 GND.n2025 240.244
R15293 GND.n7679 GND.n2025 240.244
R15294 GND.n7679 GND.n2020 240.244
R15295 GND.n7686 GND.n2020 240.244
R15296 GND.n7686 GND.n2015 240.244
R15297 GND.n2015 GND.n2001 240.244
R15298 GND.n7703 GND.n2001 240.244
R15299 GND.n7703 GND.n1996 240.244
R15300 GND.n7710 GND.n1996 240.244
R15301 GND.n7710 GND.n1991 240.244
R15302 GND.n1991 GND.n1978 240.244
R15303 GND.n7728 GND.n1978 240.244
R15304 GND.n7728 GND.n1973 240.244
R15305 GND.n7735 GND.n1973 240.244
R15306 GND.n7735 GND.n1969 240.244
R15307 GND.n1969 GND.n1956 240.244
R15308 GND.n7753 GND.n1956 240.244
R15309 GND.n7753 GND.n1951 240.244
R15310 GND.n7760 GND.n1951 240.244
R15311 GND.n7760 GND.n1946 240.244
R15312 GND.n1946 GND.n1934 240.244
R15313 GND.n7778 GND.n1934 240.244
R15314 GND.n7778 GND.n1929 240.244
R15315 GND.n7785 GND.n1929 240.244
R15316 GND.n7785 GND.n1924 240.244
R15317 GND.n1924 GND.n1911 240.244
R15318 GND.n7802 GND.n1911 240.244
R15319 GND.n7802 GND.n1906 240.244
R15320 GND.n7814 GND.n1906 240.244
R15321 GND.n7814 GND.n1901 240.244
R15322 GND.n7808 GND.n1901 240.244
R15323 GND.n7808 GND.n1890 240.244
R15324 GND.n7830 GND.n1890 240.244
R15325 GND.n7830 GND.n1772 240.244
R15326 GND.n2388 GND.n2387 240.244
R15327 GND.n2393 GND.n2392 240.244
R15328 GND.n2385 GND.n2384 240.244
R15329 GND.n2401 GND.n2400 240.244
R15330 GND.n2381 GND.n2380 240.244
R15331 GND.n2376 GND.n1465 240.244
R15332 GND.n8095 GND.n1507 240.244
R15333 GND.n1564 GND.n1507 240.244
R15334 GND.n1564 GND.n1531 240.244
R15335 GND.n1550 GND.n1531 240.244
R15336 GND.n8079 GND.n1550 240.244
R15337 GND.n8079 GND.n1551 240.244
R15338 GND.n2504 GND.n1551 240.244
R15339 GND.n2504 GND.n2363 240.244
R15340 GND.n2524 GND.n2363 240.244
R15341 GND.n2528 GND.n2524 240.244
R15342 GND.n2528 GND.n2526 240.244
R15343 GND.n2526 GND.n2352 240.244
R15344 GND.n2352 GND.n2340 240.244
R15345 GND.n2549 GND.n2340 240.244
R15346 GND.n2553 GND.n2549 240.244
R15347 GND.n2553 GND.n2552 240.244
R15348 GND.n2552 GND.n2329 240.244
R15349 GND.n2329 GND.n2319 240.244
R15350 GND.n2574 GND.n2319 240.244
R15351 GND.n2577 GND.n2574 240.244
R15352 GND.n2577 GND.n2576 240.244
R15353 GND.n2576 GND.n2306 240.244
R15354 GND.n2306 GND.n2294 240.244
R15355 GND.n2598 GND.n2294 240.244
R15356 GND.n2602 GND.n2598 240.244
R15357 GND.n2602 GND.n2601 240.244
R15358 GND.n2601 GND.n2282 240.244
R15359 GND.n2282 GND.n2272 240.244
R15360 GND.n2632 GND.n2272 240.244
R15361 GND.n2635 GND.n2632 240.244
R15362 GND.n2635 GND.n2633 240.244
R15363 GND.n2633 GND.n2252 240.244
R15364 GND.n2698 GND.n2252 240.244
R15365 GND.n2702 GND.n2698 240.244
R15366 GND.n2702 GND.n2700 240.244
R15367 GND.n2700 GND.n2242 240.244
R15368 GND.n2242 GND.n2230 240.244
R15369 GND.n2723 GND.n2230 240.244
R15370 GND.n2727 GND.n2723 240.244
R15371 GND.n2727 GND.n2726 240.244
R15372 GND.n2726 GND.n2219 240.244
R15373 GND.n2219 GND.n2209 240.244
R15374 GND.n2748 GND.n2209 240.244
R15375 GND.n2751 GND.n2748 240.244
R15376 GND.n2751 GND.n2750 240.244
R15377 GND.n2750 GND.n2198 240.244
R15378 GND.n2198 GND.n2120 240.244
R15379 GND.n2819 GND.n2120 240.244
R15380 GND.n2819 GND.n2818 240.244
R15381 GND.n2818 GND.n2122 240.244
R15382 GND.n2135 GND.n2122 240.244
R15383 GND.n2136 GND.n2135 240.244
R15384 GND.n2802 GND.n2136 240.244
R15385 GND.n2802 GND.n2801 240.244
R15386 GND.n2801 GND.n2143 240.244
R15387 GND.n2789 GND.n2143 240.244
R15388 GND.n2790 GND.n2789 240.244
R15389 GND.n2790 GND.n2101 240.244
R15390 GND.n2101 GND.n2089 240.244
R15391 GND.n2840 GND.n2089 240.244
R15392 GND.n2844 GND.n2840 240.244
R15393 GND.n2844 GND.n2843 240.244
R15394 GND.n2843 GND.n2077 240.244
R15395 GND.n2077 GND.n2067 240.244
R15396 GND.n2865 GND.n2067 240.244
R15397 GND.n2869 GND.n2865 240.244
R15398 GND.n2869 GND.n2867 240.244
R15399 GND.n2867 GND.n2057 240.244
R15400 GND.n2057 GND.n2056 240.244
R15401 GND.n2056 GND.n2039 240.244
R15402 GND.n7667 GND.n2039 240.244
R15403 GND.n7667 GND.n7666 240.244
R15404 GND.n7666 GND.n2028 240.244
R15405 GND.n2028 GND.n2018 240.244
R15406 GND.n7688 GND.n2018 240.244
R15407 GND.n7691 GND.n7688 240.244
R15408 GND.n7691 GND.n7690 240.244
R15409 GND.n7690 GND.n2005 240.244
R15410 GND.n2005 GND.n1993 240.244
R15411 GND.n7712 GND.n1993 240.244
R15412 GND.n7716 GND.n7712 240.244
R15413 GND.n7716 GND.n7715 240.244
R15414 GND.n7715 GND.n1981 240.244
R15415 GND.n1981 GND.n1971 240.244
R15416 GND.n7737 GND.n1971 240.244
R15417 GND.n7741 GND.n7737 240.244
R15418 GND.n7741 GND.n7739 240.244
R15419 GND.n7739 GND.n1960 240.244
R15420 GND.n1960 GND.n1948 240.244
R15421 GND.n7762 GND.n1948 240.244
R15422 GND.n7766 GND.n7762 240.244
R15423 GND.n7766 GND.n7765 240.244
R15424 GND.n7765 GND.n1937 240.244
R15425 GND.n1937 GND.n1927 240.244
R15426 GND.n7787 GND.n1927 240.244
R15427 GND.n7790 GND.n7787 240.244
R15428 GND.n7790 GND.n7789 240.244
R15429 GND.n7789 GND.n1914 240.244
R15430 GND.n1914 GND.n1903 240.244
R15431 GND.n7816 GND.n1903 240.244
R15432 GND.n7817 GND.n7816 240.244
R15433 GND.n7817 GND.n1893 240.244
R15434 GND.n7827 GND.n1893 240.244
R15435 GND.n7828 GND.n7827 240.244
R15436 GND.n7828 GND.n1774 240.244
R15437 GND.n3321 GND.n3320 240.244
R15438 GND.n6403 GND.n3330 240.244
R15439 GND.n6406 GND.n3331 240.244
R15440 GND.n3339 GND.n3338 240.244
R15441 GND.n6408 GND.n3350 240.244
R15442 GND.n6411 GND.n3351 240.244
R15443 GND.n3965 GND.n3964 240.244
R15444 GND.n3971 GND.n3966 240.244
R15445 GND.n6417 GND.n3972 240.244
R15446 GND.n3052 GND.n3013 240.244
R15447 GND.n3024 GND.n3013 240.244
R15448 GND.n7552 GND.n3024 240.244
R15449 GND.n7552 GND.n3025 240.244
R15450 GND.n3058 GND.n3025 240.244
R15451 GND.n3059 GND.n3058 240.244
R15452 GND.n3060 GND.n3059 240.244
R15453 GND.n4641 GND.n3060 240.244
R15454 GND.n4641 GND.n3063 240.244
R15455 GND.n3064 GND.n3063 240.244
R15456 GND.n3065 GND.n3064 240.244
R15457 GND.n4616 GND.n3065 240.244
R15458 GND.n4616 GND.n3068 240.244
R15459 GND.n3069 GND.n3068 240.244
R15460 GND.n3070 GND.n3069 240.244
R15461 GND.n4989 GND.n3070 240.244
R15462 GND.n4989 GND.n3073 240.244
R15463 GND.n3074 GND.n3073 240.244
R15464 GND.n3075 GND.n3074 240.244
R15465 GND.n5041 GND.n3075 240.244
R15466 GND.n5041 GND.n3078 240.244
R15467 GND.n3079 GND.n3078 240.244
R15468 GND.n3080 GND.n3079 240.244
R15469 GND.n4561 GND.n3080 240.244
R15470 GND.n4561 GND.n3083 240.244
R15471 GND.n3084 GND.n3083 240.244
R15472 GND.n3085 GND.n3084 240.244
R15473 GND.n4545 GND.n3085 240.244
R15474 GND.n4545 GND.n3088 240.244
R15475 GND.n3089 GND.n3088 240.244
R15476 GND.n3090 GND.n3089 240.244
R15477 GND.n4522 GND.n3090 240.244
R15478 GND.n4522 GND.n3093 240.244
R15479 GND.n3094 GND.n3093 240.244
R15480 GND.n3095 GND.n3094 240.244
R15481 GND.n5143 GND.n3095 240.244
R15482 GND.n5143 GND.n3098 240.244
R15483 GND.n3099 GND.n3098 240.244
R15484 GND.n3100 GND.n3099 240.244
R15485 GND.n4483 GND.n3100 240.244
R15486 GND.n4483 GND.n3103 240.244
R15487 GND.n3104 GND.n3103 240.244
R15488 GND.n3105 GND.n3104 240.244
R15489 GND.n4464 GND.n3105 240.244
R15490 GND.n4464 GND.n3108 240.244
R15491 GND.n3109 GND.n3108 240.244
R15492 GND.n3110 GND.n3109 240.244
R15493 GND.n4441 GND.n3110 240.244
R15494 GND.n4441 GND.n3113 240.244
R15495 GND.n3114 GND.n3113 240.244
R15496 GND.n3115 GND.n3114 240.244
R15497 GND.n4419 GND.n3115 240.244
R15498 GND.n4419 GND.n3118 240.244
R15499 GND.n3119 GND.n3118 240.244
R15500 GND.n3120 GND.n3119 240.244
R15501 GND.n4394 GND.n3120 240.244
R15502 GND.n4394 GND.n3123 240.244
R15503 GND.n3124 GND.n3123 240.244
R15504 GND.n3125 GND.n3124 240.244
R15505 GND.n4377 GND.n3125 240.244
R15506 GND.n4377 GND.n3128 240.244
R15507 GND.n3129 GND.n3128 240.244
R15508 GND.n3130 GND.n3129 240.244
R15509 GND.n4362 GND.n3130 240.244
R15510 GND.n4362 GND.n3133 240.244
R15511 GND.n3134 GND.n3133 240.244
R15512 GND.n3135 GND.n3134 240.244
R15513 GND.n4343 GND.n3135 240.244
R15514 GND.n4343 GND.n3138 240.244
R15515 GND.n3139 GND.n3138 240.244
R15516 GND.n3140 GND.n3139 240.244
R15517 GND.n5545 GND.n3140 240.244
R15518 GND.n5545 GND.n3143 240.244
R15519 GND.n3144 GND.n3143 240.244
R15520 GND.n3145 GND.n3144 240.244
R15521 GND.n4297 GND.n3145 240.244
R15522 GND.n4297 GND.n3148 240.244
R15523 GND.n3149 GND.n3148 240.244
R15524 GND.n3150 GND.n3149 240.244
R15525 GND.n4274 GND.n3150 240.244
R15526 GND.n4274 GND.n3153 240.244
R15527 GND.n3154 GND.n3153 240.244
R15528 GND.n3155 GND.n3154 240.244
R15529 GND.n5629 GND.n3155 240.244
R15530 GND.n5629 GND.n3158 240.244
R15531 GND.n3159 GND.n3158 240.244
R15532 GND.n3160 GND.n3159 240.244
R15533 GND.n5685 GND.n3160 240.244
R15534 GND.n5685 GND.n3163 240.244
R15535 GND.n3164 GND.n3163 240.244
R15536 GND.n3165 GND.n3164 240.244
R15537 GND.n5706 GND.n3165 240.244
R15538 GND.n5706 GND.n3168 240.244
R15539 GND.n3169 GND.n3168 240.244
R15540 GND.n3170 GND.n3169 240.244
R15541 GND.n4193 GND.n3170 240.244
R15542 GND.n4193 GND.n3173 240.244
R15543 GND.n3174 GND.n3173 240.244
R15544 GND.n3175 GND.n3174 240.244
R15545 GND.n4179 GND.n3175 240.244
R15546 GND.n4179 GND.n3178 240.244
R15547 GND.n3179 GND.n3178 240.244
R15548 GND.n3180 GND.n3179 240.244
R15549 GND.n4161 GND.n3180 240.244
R15550 GND.n4161 GND.n3183 240.244
R15551 GND.n3184 GND.n3183 240.244
R15552 GND.n3185 GND.n3184 240.244
R15553 GND.n4142 GND.n3185 240.244
R15554 GND.n4142 GND.n3188 240.244
R15555 GND.n3189 GND.n3188 240.244
R15556 GND.n3190 GND.n3189 240.244
R15557 GND.n4123 GND.n3190 240.244
R15558 GND.n4123 GND.n3193 240.244
R15559 GND.n3194 GND.n3193 240.244
R15560 GND.n3195 GND.n3194 240.244
R15561 GND.n4099 GND.n3195 240.244
R15562 GND.n4099 GND.n3198 240.244
R15563 GND.n3199 GND.n3198 240.244
R15564 GND.n3200 GND.n3199 240.244
R15565 GND.n4077 GND.n3200 240.244
R15566 GND.n4077 GND.n3203 240.244
R15567 GND.n3204 GND.n3203 240.244
R15568 GND.n3205 GND.n3204 240.244
R15569 GND.n4051 GND.n3205 240.244
R15570 GND.n4051 GND.n3208 240.244
R15571 GND.n3209 GND.n3208 240.244
R15572 GND.n3210 GND.n3209 240.244
R15573 GND.n4035 GND.n3210 240.244
R15574 GND.n4035 GND.n3213 240.244
R15575 GND.n3214 GND.n3213 240.244
R15576 GND.n3215 GND.n3214 240.244
R15577 GND.n4023 GND.n3215 240.244
R15578 GND.n4023 GND.n3218 240.244
R15579 GND.n3219 GND.n3218 240.244
R15580 GND.n3220 GND.n3219 240.244
R15581 GND.n6349 GND.n3220 240.244
R15582 GND.n6349 GND.n3223 240.244
R15583 GND.n3224 GND.n3223 240.244
R15584 GND.n3225 GND.n3224 240.244
R15585 GND.n3228 GND.n3225 240.244
R15586 GND.n7342 GND.n3228 240.244
R15587 GND.n7865 GND.n1838 240.244
R15588 GND.n7865 GND.n1850 240.244
R15589 GND.n1863 GND.n1862 240.244
R15590 GND.n1871 GND.n1870 240.244
R15591 GND.n1873 GND.n1872 240.244
R15592 GND.n1885 GND.n1884 240.244
R15593 GND.n3034 GND.n3033 240.244
R15594 GND.n3038 GND.n3037 240.244
R15595 GND.n3031 GND.n3030 240.244
R15596 GND.n3047 GND.n1848 240.244
R15597 GND.n3011 GND.n1837 240.244
R15598 GND.n4668 GND.n3011 240.244
R15599 GND.n4668 GND.n3022 240.244
R15600 GND.n4857 GND.n3022 240.244
R15601 GND.n4857 GND.n4654 240.244
R15602 GND.n4889 GND.n4654 240.244
R15603 GND.n4889 GND.n4655 240.244
R15604 GND.n4885 GND.n4655 240.244
R15605 GND.n4885 GND.n4884 240.244
R15606 GND.n4884 GND.n4883 240.244
R15607 GND.n4883 GND.n4629 240.244
R15608 GND.n4879 GND.n4629 240.244
R15609 GND.n4879 GND.n4619 240.244
R15610 GND.n4876 GND.n4619 240.244
R15611 GND.n4876 GND.n4875 240.244
R15612 GND.n4875 GND.n4599 240.244
R15613 GND.n4599 GND.n4588 240.244
R15614 GND.n5001 GND.n4588 240.244
R15615 GND.n5001 GND.n4584 240.244
R15616 GND.n5040 GND.n4584 240.244
R15617 GND.n5040 GND.n4576 240.244
R15618 GND.n5036 GND.n4576 240.244
R15619 GND.n5036 GND.n4568 240.244
R15620 GND.n5033 GND.n4568 240.244
R15621 GND.n5033 GND.n5032 240.244
R15622 GND.n5032 GND.n5031 240.244
R15623 GND.n5031 GND.n5011 240.244
R15624 GND.n5011 GND.n4544 240.244
R15625 GND.n4544 GND.n4537 240.244
R15626 GND.n5025 GND.n4537 240.244
R15627 GND.n5025 GND.n4529 240.244
R15628 GND.n5022 GND.n4529 240.244
R15629 GND.n5022 GND.n4511 240.244
R15630 GND.n4511 GND.n4502 240.244
R15631 GND.n5164 GND.n4502 240.244
R15632 GND.n5164 GND.n4498 240.244
R15633 GND.n5204 GND.n4498 240.244
R15634 GND.n5204 GND.n4491 240.244
R15635 GND.n5200 GND.n4491 240.244
R15636 GND.n5200 GND.n4482 240.244
R15637 GND.n5197 GND.n4482 240.244
R15638 GND.n5197 GND.n5196 240.244
R15639 GND.n5196 GND.n5195 240.244
R15640 GND.n5195 GND.n5174 240.244
R15641 GND.n5174 GND.n4457 240.244
R15642 GND.n5190 GND.n4457 240.244
R15643 GND.n5190 GND.n4448 240.244
R15644 GND.n5187 GND.n4448 240.244
R15645 GND.n5187 GND.n5186 240.244
R15646 GND.n5186 GND.n4428 240.244
R15647 GND.n4428 GND.n4416 240.244
R15648 GND.n5325 GND.n4416 240.244
R15649 GND.n5325 GND.n4412 240.244
R15650 GND.n5366 GND.n4412 240.244
R15651 GND.n5366 GND.n4405 240.244
R15652 GND.n5362 GND.n4405 240.244
R15653 GND.n5362 GND.n4397 240.244
R15654 GND.n5359 GND.n4397 240.244
R15655 GND.n5359 GND.n5358 240.244
R15656 GND.n5358 GND.n5357 240.244
R15657 GND.n5357 GND.n5335 240.244
R15658 GND.n5335 GND.n4371 240.244
R15659 GND.n5352 GND.n4371 240.244
R15660 GND.n5352 GND.n4361 240.244
R15661 GND.n5348 GND.n4361 240.244
R15662 GND.n5348 GND.n5347 240.244
R15663 GND.n5347 GND.n4341 240.244
R15664 GND.n4341 GND.n4330 240.244
R15665 GND.n5485 GND.n4330 240.244
R15666 GND.n5485 GND.n4326 240.244
R15667 GND.n5536 GND.n4326 240.244
R15668 GND.n5536 GND.n4318 240.244
R15669 GND.n5532 GND.n4318 240.244
R15670 GND.n5532 GND.n4310 240.244
R15671 GND.n5529 GND.n4310 240.244
R15672 GND.n5529 GND.n5528 240.244
R15673 GND.n5528 GND.n5527 240.244
R15674 GND.n5527 GND.n5496 240.244
R15675 GND.n5496 GND.n4286 240.244
R15676 GND.n5522 GND.n4286 240.244
R15677 GND.n5522 GND.n4277 240.244
R15678 GND.n5519 GND.n4277 240.244
R15679 GND.n5519 GND.n5518 240.244
R15680 GND.n5518 GND.n4257 240.244
R15681 GND.n5514 GND.n4257 240.244
R15682 GND.n5514 GND.n4249 240.244
R15683 GND.n5511 GND.n4249 240.244
R15684 GND.n5511 GND.n4233 240.244
R15685 GND.n4233 GND.n4224 240.244
R15686 GND.n5697 GND.n4224 240.244
R15687 GND.n5697 GND.n4220 240.244
R15688 GND.n5705 GND.n4220 240.244
R15689 GND.n5705 GND.n4210 240.244
R15690 GND.n4210 GND.n4200 240.244
R15691 GND.n5731 GND.n4200 240.244
R15692 GND.n5731 GND.n4196 240.244
R15693 GND.n5792 GND.n4196 240.244
R15694 GND.n5792 GND.n4187 240.244
R15695 GND.n5788 GND.n4187 240.244
R15696 GND.n5788 GND.n4178 240.244
R15697 GND.n5785 GND.n4178 240.244
R15698 GND.n5785 GND.n5784 240.244
R15699 GND.n5784 GND.n5783 240.244
R15700 GND.n5783 GND.n5741 240.244
R15701 GND.n5741 GND.n4157 240.244
R15702 GND.n4157 GND.n4149 240.244
R15703 GND.n5777 GND.n4149 240.244
R15704 GND.n5777 GND.n4141 240.244
R15705 GND.n5774 GND.n4141 240.244
R15706 GND.n5774 GND.n5773 240.244
R15707 GND.n5773 GND.n5772 240.244
R15708 GND.n5772 GND.n5751 240.244
R15709 GND.n5751 GND.n4116 240.244
R15710 GND.n5767 GND.n4116 240.244
R15711 GND.n5767 GND.n4106 240.244
R15712 GND.n5764 GND.n4106 240.244
R15713 GND.n5764 GND.n5763 240.244
R15714 GND.n5763 GND.n4086 240.244
R15715 GND.n4086 GND.n4074 240.244
R15716 GND.n5971 GND.n4074 240.244
R15717 GND.n5971 GND.n4070 240.244
R15718 GND.n6000 GND.n4070 240.244
R15719 GND.n6000 GND.n4062 240.244
R15720 GND.n5996 GND.n4062 240.244
R15721 GND.n5996 GND.n4054 240.244
R15722 GND.n5993 GND.n4054 240.244
R15723 GND.n5993 GND.n5992 240.244
R15724 GND.n5992 GND.n5991 240.244
R15725 GND.n5991 GND.n5981 240.244
R15726 GND.n5981 GND.n4030 240.244
R15727 GND.n4030 GND.n4021 240.244
R15728 GND.n4021 GND.n4010 240.244
R15729 GND.n6096 GND.n4010 240.244
R15730 GND.n6096 GND.n4006 240.244
R15731 GND.n6340 GND.n4006 240.244
R15732 GND.n6340 GND.n3999 240.244
R15733 GND.n6336 GND.n3999 240.244
R15734 GND.n6336 GND.n3991 240.244
R15735 GND.n6333 GND.n3991 240.244
R15736 GND.n6333 GND.n6332 240.244
R15737 GND.n6332 GND.n3231 240.244
R15738 GND.n8291 GND.n1319 240.244
R15739 GND.n8291 GND.n1317 240.244
R15740 GND.n8295 GND.n1317 240.244
R15741 GND.n8295 GND.n1313 240.244
R15742 GND.n8301 GND.n1313 240.244
R15743 GND.n8301 GND.n1311 240.244
R15744 GND.n8305 GND.n1311 240.244
R15745 GND.n8305 GND.n1307 240.244
R15746 GND.n8311 GND.n1307 240.244
R15747 GND.n8311 GND.n1305 240.244
R15748 GND.n8315 GND.n1305 240.244
R15749 GND.n8315 GND.n1301 240.244
R15750 GND.n8321 GND.n1301 240.244
R15751 GND.n8321 GND.n1299 240.244
R15752 GND.n8325 GND.n1299 240.244
R15753 GND.n8325 GND.n1295 240.244
R15754 GND.n8331 GND.n1295 240.244
R15755 GND.n8331 GND.n1293 240.244
R15756 GND.n8335 GND.n1293 240.244
R15757 GND.n8335 GND.n1289 240.244
R15758 GND.n8341 GND.n1289 240.244
R15759 GND.n8341 GND.n1287 240.244
R15760 GND.n8345 GND.n1287 240.244
R15761 GND.n8345 GND.n1283 240.244
R15762 GND.n8351 GND.n1283 240.244
R15763 GND.n8351 GND.n1281 240.244
R15764 GND.n8355 GND.n1281 240.244
R15765 GND.n8355 GND.n1277 240.244
R15766 GND.n8361 GND.n1277 240.244
R15767 GND.n8361 GND.n1275 240.244
R15768 GND.n8365 GND.n1275 240.244
R15769 GND.n8365 GND.n1271 240.244
R15770 GND.n8371 GND.n1271 240.244
R15771 GND.n8371 GND.n1269 240.244
R15772 GND.n8375 GND.n1269 240.244
R15773 GND.n8375 GND.n1265 240.244
R15774 GND.n8381 GND.n1265 240.244
R15775 GND.n8381 GND.n1263 240.244
R15776 GND.n8385 GND.n1263 240.244
R15777 GND.n8385 GND.n1259 240.244
R15778 GND.n8391 GND.n1259 240.244
R15779 GND.n8391 GND.n1257 240.244
R15780 GND.n8395 GND.n1257 240.244
R15781 GND.n8395 GND.n1253 240.244
R15782 GND.n8401 GND.n1253 240.244
R15783 GND.n8401 GND.n1251 240.244
R15784 GND.n8405 GND.n1251 240.244
R15785 GND.n8405 GND.n1247 240.244
R15786 GND.n8411 GND.n1247 240.244
R15787 GND.n8411 GND.n1245 240.244
R15788 GND.n8415 GND.n1245 240.244
R15789 GND.n8415 GND.n1241 240.244
R15790 GND.n8421 GND.n1241 240.244
R15791 GND.n8421 GND.n1239 240.244
R15792 GND.n8425 GND.n1239 240.244
R15793 GND.n8425 GND.n1235 240.244
R15794 GND.n8431 GND.n1235 240.244
R15795 GND.n8431 GND.n1233 240.244
R15796 GND.n8435 GND.n1233 240.244
R15797 GND.n8435 GND.n1229 240.244
R15798 GND.n8441 GND.n1229 240.244
R15799 GND.n8441 GND.n1227 240.244
R15800 GND.n8445 GND.n1227 240.244
R15801 GND.n8445 GND.n1223 240.244
R15802 GND.n8451 GND.n1223 240.244
R15803 GND.n8451 GND.n1221 240.244
R15804 GND.n8455 GND.n1221 240.244
R15805 GND.n8455 GND.n1217 240.244
R15806 GND.n8461 GND.n1217 240.244
R15807 GND.n8461 GND.n1215 240.244
R15808 GND.n8465 GND.n1215 240.244
R15809 GND.n8465 GND.n1211 240.244
R15810 GND.n8471 GND.n1211 240.244
R15811 GND.n8471 GND.n1209 240.244
R15812 GND.n8475 GND.n1209 240.244
R15813 GND.n8475 GND.n1205 240.244
R15814 GND.n8481 GND.n1205 240.244
R15815 GND.n8481 GND.n1203 240.244
R15816 GND.n8485 GND.n1203 240.244
R15817 GND.n8485 GND.n1199 240.244
R15818 GND.n8491 GND.n1199 240.244
R15819 GND.n8491 GND.n1197 240.244
R15820 GND.n8495 GND.n1197 240.244
R15821 GND.n8495 GND.n1193 240.244
R15822 GND.n8501 GND.n1193 240.244
R15823 GND.n8501 GND.n1191 240.244
R15824 GND.n8505 GND.n1191 240.244
R15825 GND.n8505 GND.n1187 240.244
R15826 GND.n8511 GND.n1187 240.244
R15827 GND.n8511 GND.n1185 240.244
R15828 GND.n8515 GND.n1185 240.244
R15829 GND.n8515 GND.n1181 240.244
R15830 GND.n8521 GND.n1181 240.244
R15831 GND.n8521 GND.n1179 240.244
R15832 GND.n8525 GND.n1179 240.244
R15833 GND.n8525 GND.n1175 240.244
R15834 GND.n8531 GND.n1175 240.244
R15835 GND.n8531 GND.n1173 240.244
R15836 GND.n8535 GND.n1173 240.244
R15837 GND.n8535 GND.n1169 240.244
R15838 GND.n8541 GND.n1169 240.244
R15839 GND.n8541 GND.n1167 240.244
R15840 GND.n8545 GND.n1167 240.244
R15841 GND.n8545 GND.n1163 240.244
R15842 GND.n8551 GND.n1163 240.244
R15843 GND.n8551 GND.n1161 240.244
R15844 GND.n8555 GND.n1161 240.244
R15845 GND.n8555 GND.n1157 240.244
R15846 GND.n8561 GND.n1157 240.244
R15847 GND.n8561 GND.n1155 240.244
R15848 GND.n8565 GND.n1155 240.244
R15849 GND.n8565 GND.n1151 240.244
R15850 GND.n8571 GND.n1151 240.244
R15851 GND.n8571 GND.n1149 240.244
R15852 GND.n8575 GND.n1149 240.244
R15853 GND.n8575 GND.n1145 240.244
R15854 GND.n8581 GND.n1145 240.244
R15855 GND.n8581 GND.n1143 240.244
R15856 GND.n8585 GND.n1143 240.244
R15857 GND.n8585 GND.n1139 240.244
R15858 GND.n8591 GND.n1139 240.244
R15859 GND.n8591 GND.n1137 240.244
R15860 GND.n8595 GND.n1137 240.244
R15861 GND.n8595 GND.n1133 240.244
R15862 GND.n8601 GND.n1133 240.244
R15863 GND.n8601 GND.n1131 240.244
R15864 GND.n8605 GND.n1131 240.244
R15865 GND.n8605 GND.n1127 240.244
R15866 GND.n8611 GND.n1127 240.244
R15867 GND.n8611 GND.n1125 240.244
R15868 GND.n8615 GND.n1125 240.244
R15869 GND.n8615 GND.n1121 240.244
R15870 GND.n8621 GND.n1121 240.244
R15871 GND.n8621 GND.n1119 240.244
R15872 GND.n8625 GND.n1119 240.244
R15873 GND.n8625 GND.n1115 240.244
R15874 GND.n8631 GND.n1115 240.244
R15875 GND.n8631 GND.n1113 240.244
R15876 GND.n8635 GND.n1113 240.244
R15877 GND.n8635 GND.n1109 240.244
R15878 GND.n8641 GND.n1109 240.244
R15879 GND.n8641 GND.n1107 240.244
R15880 GND.n8645 GND.n1107 240.244
R15881 GND.n8645 GND.n1103 240.244
R15882 GND.n8651 GND.n1103 240.244
R15883 GND.n8651 GND.n1101 240.244
R15884 GND.n8655 GND.n1101 240.244
R15885 GND.n8655 GND.n1097 240.244
R15886 GND.n8661 GND.n1097 240.244
R15887 GND.n8661 GND.n1095 240.244
R15888 GND.n8665 GND.n1095 240.244
R15889 GND.n8665 GND.n1091 240.244
R15890 GND.n8671 GND.n1091 240.244
R15891 GND.n8671 GND.n1089 240.244
R15892 GND.n8675 GND.n1089 240.244
R15893 GND.n8675 GND.n1085 240.244
R15894 GND.n8681 GND.n1085 240.244
R15895 GND.n8681 GND.n1083 240.244
R15896 GND.n8685 GND.n1083 240.244
R15897 GND.n8685 GND.n1079 240.244
R15898 GND.n8691 GND.n1079 240.244
R15899 GND.n8691 GND.n1077 240.244
R15900 GND.n8695 GND.n1077 240.244
R15901 GND.n8695 GND.n1073 240.244
R15902 GND.n8701 GND.n1073 240.244
R15903 GND.n8701 GND.n1071 240.244
R15904 GND.n8705 GND.n1071 240.244
R15905 GND.n8705 GND.n1067 240.244
R15906 GND.n8711 GND.n1067 240.244
R15907 GND.n8711 GND.n1065 240.244
R15908 GND.n8715 GND.n1065 240.244
R15909 GND.n8715 GND.n1061 240.244
R15910 GND.n8721 GND.n1061 240.244
R15911 GND.n8721 GND.n1059 240.244
R15912 GND.n8725 GND.n1059 240.244
R15913 GND.n8725 GND.n1055 240.244
R15914 GND.n8731 GND.n1055 240.244
R15915 GND.n8731 GND.n1053 240.244
R15916 GND.n8735 GND.n1053 240.244
R15917 GND.n8735 GND.n1049 240.244
R15918 GND.n8741 GND.n1049 240.244
R15919 GND.n8741 GND.n1047 240.244
R15920 GND.n8745 GND.n1047 240.244
R15921 GND.n8745 GND.n1043 240.244
R15922 GND.n8751 GND.n1043 240.244
R15923 GND.n8751 GND.n1041 240.244
R15924 GND.n8755 GND.n1041 240.244
R15925 GND.n8755 GND.n1037 240.244
R15926 GND.n8761 GND.n1037 240.244
R15927 GND.n8761 GND.n1035 240.244
R15928 GND.n8765 GND.n1035 240.244
R15929 GND.n8765 GND.n1031 240.244
R15930 GND.n8771 GND.n1031 240.244
R15931 GND.n8771 GND.n1029 240.244
R15932 GND.n8775 GND.n1029 240.244
R15933 GND.n8775 GND.n1025 240.244
R15934 GND.n8781 GND.n1025 240.244
R15935 GND.n8781 GND.n1023 240.244
R15936 GND.n8785 GND.n1023 240.244
R15937 GND.n8785 GND.n1019 240.244
R15938 GND.n8791 GND.n1019 240.244
R15939 GND.n8791 GND.n1017 240.244
R15940 GND.n8795 GND.n1017 240.244
R15941 GND.n8795 GND.n1013 240.244
R15942 GND.n8801 GND.n1013 240.244
R15943 GND.n8801 GND.n1011 240.244
R15944 GND.n8805 GND.n1011 240.244
R15945 GND.n8805 GND.n1007 240.244
R15946 GND.n8811 GND.n1007 240.244
R15947 GND.n8811 GND.n1005 240.244
R15948 GND.n8815 GND.n1005 240.244
R15949 GND.n8815 GND.n1001 240.244
R15950 GND.n8821 GND.n1001 240.244
R15951 GND.n8821 GND.n999 240.244
R15952 GND.n8825 GND.n999 240.244
R15953 GND.n8825 GND.n995 240.244
R15954 GND.n8831 GND.n995 240.244
R15955 GND.n8831 GND.n993 240.244
R15956 GND.n8835 GND.n993 240.244
R15957 GND.n8835 GND.n989 240.244
R15958 GND.n8841 GND.n989 240.244
R15959 GND.n8841 GND.n987 240.244
R15960 GND.n8845 GND.n987 240.244
R15961 GND.n8845 GND.n983 240.244
R15962 GND.n8851 GND.n983 240.244
R15963 GND.n8851 GND.n981 240.244
R15964 GND.n8855 GND.n981 240.244
R15965 GND.n8855 GND.n977 240.244
R15966 GND.n8861 GND.n977 240.244
R15967 GND.n8861 GND.n975 240.244
R15968 GND.n8865 GND.n975 240.244
R15969 GND.n8865 GND.n971 240.244
R15970 GND.n8871 GND.n971 240.244
R15971 GND.n8871 GND.n969 240.244
R15972 GND.n8875 GND.n969 240.244
R15973 GND.n8875 GND.n965 240.244
R15974 GND.n8881 GND.n965 240.244
R15975 GND.n8881 GND.n963 240.244
R15976 GND.n8885 GND.n963 240.244
R15977 GND.n8885 GND.n959 240.244
R15978 GND.n8891 GND.n959 240.244
R15979 GND.n8891 GND.n957 240.244
R15980 GND.n8895 GND.n957 240.244
R15981 GND.n8895 GND.n953 240.244
R15982 GND.n8901 GND.n953 240.244
R15983 GND.n8901 GND.n951 240.244
R15984 GND.n8905 GND.n951 240.244
R15985 GND.n8905 GND.n947 240.244
R15986 GND.n8911 GND.n947 240.244
R15987 GND.n8911 GND.n945 240.244
R15988 GND.n8915 GND.n945 240.244
R15989 GND.n8915 GND.n941 240.244
R15990 GND.n8921 GND.n941 240.244
R15991 GND.n8921 GND.n939 240.244
R15992 GND.n8925 GND.n939 240.244
R15993 GND.n8925 GND.n935 240.244
R15994 GND.n8931 GND.n935 240.244
R15995 GND.n8931 GND.n933 240.244
R15996 GND.n8935 GND.n933 240.244
R15997 GND.n8935 GND.n929 240.244
R15998 GND.n8941 GND.n929 240.244
R15999 GND.n8941 GND.n927 240.244
R16000 GND.n8945 GND.n927 240.244
R16001 GND.n8945 GND.n923 240.244
R16002 GND.n8951 GND.n923 240.244
R16003 GND.n8951 GND.n921 240.244
R16004 GND.n8955 GND.n921 240.244
R16005 GND.n8955 GND.n917 240.244
R16006 GND.n8961 GND.n917 240.244
R16007 GND.n8961 GND.n915 240.244
R16008 GND.n8965 GND.n915 240.244
R16009 GND.n8965 GND.n911 240.244
R16010 GND.n8971 GND.n911 240.244
R16011 GND.n8971 GND.n909 240.244
R16012 GND.n8975 GND.n909 240.244
R16013 GND.n8975 GND.n905 240.244
R16014 GND.n8981 GND.n905 240.244
R16015 GND.n8981 GND.n903 240.244
R16016 GND.n8985 GND.n903 240.244
R16017 GND.n8985 GND.n899 240.244
R16018 GND.n8991 GND.n899 240.244
R16019 GND.n8991 GND.n897 240.244
R16020 GND.n8995 GND.n897 240.244
R16021 GND.n8995 GND.n893 240.244
R16022 GND.n9001 GND.n893 240.244
R16023 GND.n9001 GND.n891 240.244
R16024 GND.n9005 GND.n891 240.244
R16025 GND.n9005 GND.n887 240.244
R16026 GND.n9011 GND.n887 240.244
R16027 GND.n9011 GND.n885 240.244
R16028 GND.n9015 GND.n885 240.244
R16029 GND.n9015 GND.n881 240.244
R16030 GND.n9021 GND.n881 240.244
R16031 GND.n9021 GND.n879 240.244
R16032 GND.n9025 GND.n879 240.244
R16033 GND.n9025 GND.n875 240.244
R16034 GND.n9031 GND.n875 240.244
R16035 GND.n9031 GND.n873 240.244
R16036 GND.n9035 GND.n873 240.244
R16037 GND.n9035 GND.n869 240.244
R16038 GND.n9041 GND.n869 240.244
R16039 GND.n9041 GND.n867 240.244
R16040 GND.n9045 GND.n867 240.244
R16041 GND.n9045 GND.n863 240.244
R16042 GND.n9051 GND.n863 240.244
R16043 GND.n9051 GND.n861 240.244
R16044 GND.n9055 GND.n861 240.244
R16045 GND.n9055 GND.n857 240.244
R16046 GND.n9061 GND.n857 240.244
R16047 GND.n9061 GND.n855 240.244
R16048 GND.n9065 GND.n855 240.244
R16049 GND.n9065 GND.n851 240.244
R16050 GND.n9071 GND.n851 240.244
R16051 GND.n9071 GND.n849 240.244
R16052 GND.n9075 GND.n849 240.244
R16053 GND.n9075 GND.n845 240.244
R16054 GND.n9081 GND.n845 240.244
R16055 GND.n9081 GND.n843 240.244
R16056 GND.n9085 GND.n843 240.244
R16057 GND.n9085 GND.n839 240.244
R16058 GND.n9091 GND.n839 240.244
R16059 GND.n9091 GND.n837 240.244
R16060 GND.n9095 GND.n837 240.244
R16061 GND.n9095 GND.n833 240.244
R16062 GND.n9101 GND.n833 240.244
R16063 GND.n9101 GND.n831 240.244
R16064 GND.n9105 GND.n831 240.244
R16065 GND.n9105 GND.n827 240.244
R16066 GND.n9111 GND.n827 240.244
R16067 GND.n9111 GND.n825 240.244
R16068 GND.n9115 GND.n825 240.244
R16069 GND.n9115 GND.n821 240.244
R16070 GND.n9121 GND.n821 240.244
R16071 GND.n9121 GND.n819 240.244
R16072 GND.n9125 GND.n819 240.244
R16073 GND.n9125 GND.n815 240.244
R16074 GND.n9131 GND.n815 240.244
R16075 GND.n9131 GND.n813 240.244
R16076 GND.n9135 GND.n813 240.244
R16077 GND.n9135 GND.n809 240.244
R16078 GND.n9141 GND.n809 240.244
R16079 GND.n9141 GND.n807 240.244
R16080 GND.n9145 GND.n807 240.244
R16081 GND.n9145 GND.n803 240.244
R16082 GND.n9151 GND.n803 240.244
R16083 GND.n9151 GND.n801 240.244
R16084 GND.n9155 GND.n801 240.244
R16085 GND.n9155 GND.n797 240.244
R16086 GND.n9161 GND.n797 240.244
R16087 GND.n9161 GND.n795 240.244
R16088 GND.n9165 GND.n795 240.244
R16089 GND.n9165 GND.n791 240.244
R16090 GND.n9171 GND.n791 240.244
R16091 GND.n9171 GND.n789 240.244
R16092 GND.n9175 GND.n789 240.244
R16093 GND.n9175 GND.n785 240.244
R16094 GND.n9181 GND.n785 240.244
R16095 GND.n9181 GND.n783 240.244
R16096 GND.n9185 GND.n783 240.244
R16097 GND.n9185 GND.n779 240.244
R16098 GND.n9191 GND.n779 240.244
R16099 GND.n9191 GND.n777 240.244
R16100 GND.n9195 GND.n777 240.244
R16101 GND.n9195 GND.n773 240.244
R16102 GND.n9201 GND.n773 240.244
R16103 GND.n9201 GND.n771 240.244
R16104 GND.n9205 GND.n771 240.244
R16105 GND.n9205 GND.n767 240.244
R16106 GND.n9211 GND.n767 240.244
R16107 GND.n9211 GND.n765 240.244
R16108 GND.n9215 GND.n765 240.244
R16109 GND.n9215 GND.n761 240.244
R16110 GND.n9221 GND.n761 240.244
R16111 GND.n9221 GND.n759 240.244
R16112 GND.n9225 GND.n759 240.244
R16113 GND.n9225 GND.n755 240.244
R16114 GND.n9231 GND.n755 240.244
R16115 GND.n9231 GND.n753 240.244
R16116 GND.n9235 GND.n753 240.244
R16117 GND.n9235 GND.n749 240.244
R16118 GND.n9241 GND.n749 240.244
R16119 GND.n9241 GND.n747 240.244
R16120 GND.n9245 GND.n747 240.244
R16121 GND.n9245 GND.n743 240.244
R16122 GND.n9251 GND.n743 240.244
R16123 GND.n9251 GND.n741 240.244
R16124 GND.n9255 GND.n741 240.244
R16125 GND.n9255 GND.n737 240.244
R16126 GND.n9261 GND.n737 240.244
R16127 GND.n9261 GND.n735 240.244
R16128 GND.n9265 GND.n735 240.244
R16129 GND.n9265 GND.n731 240.244
R16130 GND.n9271 GND.n731 240.244
R16131 GND.n9271 GND.n729 240.244
R16132 GND.n9275 GND.n729 240.244
R16133 GND.n9275 GND.n725 240.244
R16134 GND.n9281 GND.n725 240.244
R16135 GND.n9281 GND.n723 240.244
R16136 GND.n9285 GND.n723 240.244
R16137 GND.n9285 GND.n719 240.244
R16138 GND.n9291 GND.n719 240.244
R16139 GND.n9291 GND.n717 240.244
R16140 GND.n9295 GND.n717 240.244
R16141 GND.n9295 GND.n713 240.244
R16142 GND.n9301 GND.n713 240.244
R16143 GND.n9301 GND.n711 240.244
R16144 GND.n9305 GND.n711 240.244
R16145 GND.n9305 GND.n707 240.244
R16146 GND.n9311 GND.n707 240.244
R16147 GND.n9311 GND.n705 240.244
R16148 GND.n9315 GND.n705 240.244
R16149 GND.n9315 GND.n701 240.244
R16150 GND.n9321 GND.n701 240.244
R16151 GND.n9325 GND.n699 240.244
R16152 GND.n9325 GND.n695 240.244
R16153 GND.n9331 GND.n695 240.244
R16154 GND.n9331 GND.n693 240.244
R16155 GND.n9335 GND.n693 240.244
R16156 GND.n9335 GND.n689 240.244
R16157 GND.n9341 GND.n689 240.244
R16158 GND.n9341 GND.n687 240.244
R16159 GND.n9345 GND.n687 240.244
R16160 GND.n9345 GND.n683 240.244
R16161 GND.n9351 GND.n683 240.244
R16162 GND.n9351 GND.n681 240.244
R16163 GND.n9355 GND.n681 240.244
R16164 GND.n9355 GND.n677 240.244
R16165 GND.n9361 GND.n677 240.244
R16166 GND.n9361 GND.n675 240.244
R16167 GND.n9365 GND.n675 240.244
R16168 GND.n9365 GND.n671 240.244
R16169 GND.n9371 GND.n671 240.244
R16170 GND.n9371 GND.n669 240.244
R16171 GND.n9375 GND.n669 240.244
R16172 GND.n9375 GND.n665 240.244
R16173 GND.n9381 GND.n665 240.244
R16174 GND.n9381 GND.n663 240.244
R16175 GND.n9385 GND.n663 240.244
R16176 GND.n9385 GND.n659 240.244
R16177 GND.n9391 GND.n659 240.244
R16178 GND.n9391 GND.n657 240.244
R16179 GND.n9395 GND.n657 240.244
R16180 GND.n9395 GND.n653 240.244
R16181 GND.n9401 GND.n653 240.244
R16182 GND.n9401 GND.n651 240.244
R16183 GND.n9405 GND.n651 240.244
R16184 GND.n9405 GND.n647 240.244
R16185 GND.n9411 GND.n647 240.244
R16186 GND.n9411 GND.n645 240.244
R16187 GND.n9415 GND.n645 240.244
R16188 GND.n9415 GND.n641 240.244
R16189 GND.n9421 GND.n641 240.244
R16190 GND.n9421 GND.n639 240.244
R16191 GND.n9425 GND.n639 240.244
R16192 GND.n9425 GND.n635 240.244
R16193 GND.n9431 GND.n635 240.244
R16194 GND.n9431 GND.n633 240.244
R16195 GND.n9435 GND.n633 240.244
R16196 GND.n9435 GND.n629 240.244
R16197 GND.n9441 GND.n629 240.244
R16198 GND.n9441 GND.n627 240.244
R16199 GND.n9445 GND.n627 240.244
R16200 GND.n9445 GND.n623 240.244
R16201 GND.n9452 GND.n623 240.244
R16202 GND.n9452 GND.n621 240.244
R16203 GND.n9456 GND.n621 240.244
R16204 GND.n9456 GND.n617 240.244
R16205 GND.n1431 GND.n1428 240.244
R16206 GND.n8170 GND.n1431 240.244
R16207 GND.n8170 GND.n1434 240.244
R16208 GND.n8166 GND.n1434 240.244
R16209 GND.n8166 GND.n1437 240.244
R16210 GND.n8162 GND.n1437 240.244
R16211 GND.n8162 GND.n1443 240.244
R16212 GND.n8158 GND.n1443 240.244
R16213 GND.n8158 GND.n1445 240.244
R16214 GND.n8154 GND.n1445 240.244
R16215 GND.n8154 GND.n1451 240.244
R16216 GND.n1517 GND.n1451 240.244
R16217 GND.n1517 GND.n1513 240.244
R16218 GND.n8092 GND.n1513 240.244
R16219 GND.n8092 GND.n1514 240.244
R16220 GND.n8088 GND.n1514 240.244
R16221 GND.n8088 GND.n1525 240.244
R16222 GND.n2430 GND.n1525 240.244
R16223 GND.n2431 GND.n2430 240.244
R16224 GND.n2431 GND.n2424 240.244
R16225 GND.n2502 GND.n2424 240.244
R16226 GND.n2502 GND.n2425 240.244
R16227 GND.n2498 GND.n2425 240.244
R16228 GND.n2498 GND.n2497 240.244
R16229 GND.n2497 GND.n2496 240.244
R16230 GND.n2496 GND.n2439 240.244
R16231 GND.n2492 GND.n2439 240.244
R16232 GND.n2492 GND.n2491 240.244
R16233 GND.n2491 GND.n2490 240.244
R16234 GND.n2490 GND.n2445 240.244
R16235 GND.n2486 GND.n2445 240.244
R16236 GND.n2486 GND.n2485 240.244
R16237 GND.n2485 GND.n2484 240.244
R16238 GND.n2484 GND.n2451 240.244
R16239 GND.n2480 GND.n2451 240.244
R16240 GND.n2480 GND.n2479 240.244
R16241 GND.n2479 GND.n2478 240.244
R16242 GND.n2478 GND.n2457 240.244
R16243 GND.n2474 GND.n2457 240.244
R16244 GND.n2474 GND.n2473 240.244
R16245 GND.n2473 GND.n2472 240.244
R16246 GND.n2472 GND.n2463 240.244
R16247 GND.n2468 GND.n2463 240.244
R16248 GND.n2468 GND.n2260 240.244
R16249 GND.n2646 GND.n2260 240.244
R16250 GND.n2646 GND.n2255 240.244
R16251 GND.n2695 GND.n2255 240.244
R16252 GND.n2695 GND.n2256 240.244
R16253 GND.n2691 GND.n2256 240.244
R16254 GND.n2691 GND.n2690 240.244
R16255 GND.n2690 GND.n2689 240.244
R16256 GND.n2689 GND.n2654 240.244
R16257 GND.n2685 GND.n2654 240.244
R16258 GND.n2685 GND.n2684 240.244
R16259 GND.n2684 GND.n2683 240.244
R16260 GND.n2683 GND.n2660 240.244
R16261 GND.n2679 GND.n2660 240.244
R16262 GND.n2679 GND.n2678 240.244
R16263 GND.n2678 GND.n2677 240.244
R16264 GND.n2677 GND.n2668 240.244
R16265 GND.n2673 GND.n2668 240.244
R16266 GND.n2673 GND.n2125 240.244
R16267 GND.n2815 GND.n2125 240.244
R16268 GND.n2815 GND.n2126 240.244
R16269 GND.n2810 GND.n2126 240.244
R16270 GND.n2810 GND.n2129 240.244
R16271 GND.n2147 GND.n2129 240.244
R16272 GND.n2798 GND.n2147 240.244
R16273 GND.n2798 GND.n2148 240.244
R16274 GND.n2793 GND.n2148 240.244
R16275 GND.n2793 GND.n2183 240.244
R16276 GND.n2183 GND.n2152 240.244
R16277 GND.n2179 GND.n2152 240.244
R16278 GND.n2179 GND.n2178 240.244
R16279 GND.n2178 GND.n2177 240.244
R16280 GND.n2177 GND.n2156 240.244
R16281 GND.n2173 GND.n2156 240.244
R16282 GND.n2173 GND.n2172 240.244
R16283 GND.n2172 GND.n2171 240.244
R16284 GND.n2171 GND.n2162 240.244
R16285 GND.n2167 GND.n2162 240.244
R16286 GND.n2167 GND.n2045 240.244
R16287 GND.n2891 GND.n2045 240.244
R16288 GND.n2891 GND.n2040 240.244
R16289 GND.n7662 GND.n2040 240.244
R16290 GND.n7662 GND.n2041 240.244
R16291 GND.n7658 GND.n2041 240.244
R16292 GND.n7658 GND.n7657 240.244
R16293 GND.n7657 GND.n7656 240.244
R16294 GND.n7656 GND.n2899 240.244
R16295 GND.n7652 GND.n2899 240.244
R16296 GND.n7652 GND.n7651 240.244
R16297 GND.n7651 GND.n7650 240.244
R16298 GND.n7650 GND.n2905 240.244
R16299 GND.n7646 GND.n2905 240.244
R16300 GND.n7646 GND.n7645 240.244
R16301 GND.n7645 GND.n7644 240.244
R16302 GND.n7644 GND.n2911 240.244
R16303 GND.n7640 GND.n2911 240.244
R16304 GND.n7640 GND.n7639 240.244
R16305 GND.n7639 GND.n7638 240.244
R16306 GND.n7638 GND.n2917 240.244
R16307 GND.n7634 GND.n2917 240.244
R16308 GND.n7634 GND.n7633 240.244
R16309 GND.n7633 GND.n7632 240.244
R16310 GND.n7632 GND.n2923 240.244
R16311 GND.n7628 GND.n2923 240.244
R16312 GND.n7628 GND.n7627 240.244
R16313 GND.n7627 GND.n7626 240.244
R16314 GND.n7626 GND.n2929 240.244
R16315 GND.n7622 GND.n2929 240.244
R16316 GND.n7622 GND.n7621 240.244
R16317 GND.n7621 GND.n7620 240.244
R16318 GND.n7620 GND.n2935 240.244
R16319 GND.n7616 GND.n2935 240.244
R16320 GND.n7616 GND.n7615 240.244
R16321 GND.n7615 GND.n7614 240.244
R16322 GND.n7614 GND.n2941 240.244
R16323 GND.n7610 GND.n2941 240.244
R16324 GND.n7610 GND.n7609 240.244
R16325 GND.n7609 GND.n7608 240.244
R16326 GND.n7608 GND.n2947 240.244
R16327 GND.n7604 GND.n2947 240.244
R16328 GND.n7604 GND.n2953 240.244
R16329 GND.n7600 GND.n2953 240.244
R16330 GND.n7600 GND.n2956 240.244
R16331 GND.n7596 GND.n2956 240.244
R16332 GND.n7596 GND.n2962 240.244
R16333 GND.n7586 GND.n2962 240.244
R16334 GND.n7586 GND.n2974 240.244
R16335 GND.n7582 GND.n2974 240.244
R16336 GND.n7582 GND.n2980 240.244
R16337 GND.n7572 GND.n2980 240.244
R16338 GND.n7572 GND.n2993 240.244
R16339 GND.n7568 GND.n2993 240.244
R16340 GND.n7568 GND.n2999 240.244
R16341 GND.n7558 GND.n2999 240.244
R16342 GND.n7558 GND.n3014 240.244
R16343 GND.n7554 GND.n3014 240.244
R16344 GND.n7554 GND.n3020 240.244
R16345 GND.n4890 GND.n3020 240.244
R16346 GND.n4905 GND.n4890 240.244
R16347 GND.n4905 GND.n4891 240.244
R16348 GND.n4901 GND.n4891 240.244
R16349 GND.n4901 GND.n4900 240.244
R16350 GND.n4900 GND.n4626 240.244
R16351 GND.n4937 GND.n4626 240.244
R16352 GND.n4937 GND.n4621 240.244
R16353 GND.n4945 GND.n4621 240.244
R16354 GND.n4945 GND.n4622 240.244
R16355 GND.n4622 GND.n4597 240.244
R16356 GND.n4991 GND.n4597 240.244
R16357 GND.n4991 GND.n4591 240.244
R16358 GND.n4999 GND.n4591 240.244
R16359 GND.n4999 GND.n4593 240.244
R16360 GND.n4593 GND.n4574 240.244
R16361 GND.n5051 GND.n4574 240.244
R16362 GND.n5051 GND.n4569 240.244
R16363 GND.n5068 GND.n4569 240.244
R16364 GND.n5068 GND.n4570 240.244
R16365 GND.n5064 GND.n4570 240.244
R16366 GND.n5064 GND.n5063 240.244
R16367 GND.n5063 GND.n5062 240.244
R16368 GND.n5062 GND.n4535 240.244
R16369 GND.n5109 GND.n4535 240.244
R16370 GND.n5109 GND.n4531 240.244
R16371 GND.n5115 GND.n4531 240.244
R16372 GND.n5115 GND.n4509 240.244
R16373 GND.n5154 GND.n4509 240.244
R16374 GND.n5154 GND.n4504 240.244
R16375 GND.n5162 GND.n4504 240.244
R16376 GND.n5162 GND.n4505 240.244
R16377 GND.n4505 GND.n4489 240.244
R16378 GND.n5214 GND.n4489 240.244
R16379 GND.n5214 GND.n4484 240.244
R16380 GND.n5228 GND.n4484 240.244
R16381 GND.n5228 GND.n4485 240.244
R16382 GND.n5224 GND.n4485 240.244
R16383 GND.n5224 GND.n5223 240.244
R16384 GND.n5223 GND.n4454 240.244
R16385 GND.n5260 GND.n4454 240.244
R16386 GND.n5260 GND.n4449 240.244
R16387 GND.n5268 GND.n4449 240.244
R16388 GND.n5268 GND.n4450 240.244
R16389 GND.n4450 GND.n4426 240.244
R16390 GND.n5315 GND.n4426 240.244
R16391 GND.n5315 GND.n4420 240.244
R16392 GND.n5323 GND.n4420 240.244
R16393 GND.n5323 GND.n4422 240.244
R16394 GND.n4422 GND.n4403 240.244
R16395 GND.n5376 GND.n4403 240.244
R16396 GND.n5376 GND.n4398 240.244
R16397 GND.n5390 GND.n4398 240.244
R16398 GND.n5390 GND.n4399 240.244
R16399 GND.n5386 GND.n4399 240.244
R16400 GND.n5386 GND.n5385 240.244
R16401 GND.n5385 GND.n4368 240.244
R16402 GND.n5422 GND.n4368 240.244
R16403 GND.n5422 GND.n4363 240.244
R16404 GND.n5430 GND.n4363 240.244
R16405 GND.n5430 GND.n4364 240.244
R16406 GND.n4364 GND.n4339 240.244
R16407 GND.n5475 GND.n4339 240.244
R16408 GND.n5475 GND.n4333 240.244
R16409 GND.n5483 GND.n4333 240.244
R16410 GND.n5483 GND.n4335 240.244
R16411 GND.n4335 GND.n4316 240.244
R16412 GND.n5547 GND.n4316 240.244
R16413 GND.n5547 GND.n4311 240.244
R16414 GND.n5561 GND.n4311 240.244
R16415 GND.n5561 GND.n4312 240.244
R16416 GND.n5557 GND.n4312 240.244
R16417 GND.n5557 GND.n5556 240.244
R16418 GND.n5556 GND.n4283 240.244
R16419 GND.n5593 GND.n4283 240.244
R16420 GND.n5593 GND.n4278 240.244
R16421 GND.n5601 GND.n4278 240.244
R16422 GND.n5601 GND.n4279 240.244
R16423 GND.n4279 GND.n4255 240.244
R16424 GND.n5631 GND.n4255 240.244
R16425 GND.n5631 GND.n4251 240.244
R16426 GND.n5637 GND.n4251 240.244
R16427 GND.n5637 GND.n4231 240.244
R16428 GND.n5687 GND.n4231 240.244
R16429 GND.n5687 GND.n4226 240.244
R16430 GND.n5695 GND.n4226 240.244
R16431 GND.n5695 GND.n4227 240.244
R16432 GND.n4227 GND.n4208 240.244
R16433 GND.n5721 GND.n4208 240.244
R16434 GND.n5721 GND.n4203 240.244
R16435 GND.n5729 GND.n4203 240.244
R16436 GND.n5729 GND.n4204 240.244
R16437 GND.n4204 GND.n4185 240.244
R16438 GND.n5802 GND.n4185 240.244
R16439 GND.n5802 GND.n4180 240.244
R16440 GND.n5819 GND.n4180 240.244
R16441 GND.n5819 GND.n4181 240.244
R16442 GND.n5815 GND.n4181 240.244
R16443 GND.n5815 GND.n5814 240.244
R16444 GND.n5814 GND.n5813 240.244
R16445 GND.n5813 GND.n4148 240.244
R16446 GND.n5862 GND.n4148 240.244
R16447 GND.n5862 GND.n4143 240.244
R16448 GND.n5876 GND.n4143 240.244
R16449 GND.n5876 GND.n4144 240.244
R16450 GND.n5872 GND.n4144 240.244
R16451 GND.n5872 GND.n5871 240.244
R16452 GND.n5871 GND.n4113 240.244
R16453 GND.n5908 GND.n4113 240.244
R16454 GND.n5908 GND.n4108 240.244
R16455 GND.n5916 GND.n4108 240.244
R16456 GND.n5916 GND.n4109 240.244
R16457 GND.n4109 GND.n4084 240.244
R16458 GND.n5961 GND.n4084 240.244
R16459 GND.n5961 GND.n4078 240.244
R16460 GND.n5969 GND.n4078 240.244
R16461 GND.n5969 GND.n4080 240.244
R16462 GND.n4080 GND.n4060 240.244
R16463 GND.n6010 GND.n4060 240.244
R16464 GND.n6010 GND.n4055 240.244
R16465 GND.n6027 GND.n4055 240.244
R16466 GND.n6027 GND.n4056 240.244
R16467 GND.n6023 GND.n4056 240.244
R16468 GND.n6023 GND.n6022 240.244
R16469 GND.n6022 GND.n6021 240.244
R16470 GND.n6021 GND.n4019 240.244
R16471 GND.n6086 GND.n4019 240.244
R16472 GND.n6086 GND.n4013 240.244
R16473 GND.n6094 GND.n4013 240.244
R16474 GND.n6094 GND.n4015 240.244
R16475 GND.n4015 GND.n3997 240.244
R16476 GND.n6351 GND.n3997 240.244
R16477 GND.n6351 GND.n3992 240.244
R16478 GND.n6360 GND.n3992 240.244
R16479 GND.n6360 GND.n3993 240.244
R16480 GND.n3993 GND.n3233 240.244
R16481 GND.n7340 GND.n3233 240.244
R16482 GND.n7340 GND.n3234 240.244
R16483 GND.n7336 GND.n3234 240.244
R16484 GND.n7336 GND.n3240 240.244
R16485 GND.n7326 GND.n3240 240.244
R16486 GND.n7326 GND.n3251 240.244
R16487 GND.n7322 GND.n3251 240.244
R16488 GND.n7322 GND.n3257 240.244
R16489 GND.n3274 GND.n3257 240.244
R16490 GND.n7307 GND.n3274 240.244
R16491 GND.n7307 GND.n3275 240.244
R16492 GND.n7303 GND.n3275 240.244
R16493 GND.n7303 GND.n3283 240.244
R16494 GND.n7299 GND.n3283 240.244
R16495 GND.n7299 GND.n3285 240.244
R16496 GND.n7295 GND.n3285 240.244
R16497 GND.n7295 GND.n3291 240.244
R16498 GND.n6446 GND.n3291 240.244
R16499 GND.n6447 GND.n6446 240.244
R16500 GND.n6448 GND.n6447 240.244
R16501 GND.n6448 GND.n6438 240.244
R16502 GND.n6579 GND.n6438 240.244
R16503 GND.n6579 GND.n6439 240.244
R16504 GND.n6575 GND.n6439 240.244
R16505 GND.n6575 GND.n6574 240.244
R16506 GND.n6574 GND.n6573 240.244
R16507 GND.n6573 GND.n6456 240.244
R16508 GND.n6569 GND.n6456 240.244
R16509 GND.n6569 GND.n6568 240.244
R16510 GND.n6568 GND.n6567 240.244
R16511 GND.n6567 GND.n6462 240.244
R16512 GND.n6563 GND.n6462 240.244
R16513 GND.n6563 GND.n6562 240.244
R16514 GND.n6562 GND.n6561 240.244
R16515 GND.n6561 GND.n6468 240.244
R16516 GND.n6557 GND.n6468 240.244
R16517 GND.n6557 GND.n6556 240.244
R16518 GND.n6556 GND.n6555 240.244
R16519 GND.n6555 GND.n6474 240.244
R16520 GND.n6551 GND.n6474 240.244
R16521 GND.n6551 GND.n6550 240.244
R16522 GND.n6550 GND.n6549 240.244
R16523 GND.n6549 GND.n6480 240.244
R16524 GND.n6545 GND.n6480 240.244
R16525 GND.n6545 GND.n6544 240.244
R16526 GND.n6544 GND.n6543 240.244
R16527 GND.n6543 GND.n6486 240.244
R16528 GND.n6539 GND.n6486 240.244
R16529 GND.n6539 GND.n6538 240.244
R16530 GND.n6538 GND.n6537 240.244
R16531 GND.n6537 GND.n6492 240.244
R16532 GND.n6533 GND.n6492 240.244
R16533 GND.n6533 GND.n6532 240.244
R16534 GND.n6532 GND.n6531 240.244
R16535 GND.n6531 GND.n6498 240.244
R16536 GND.n6527 GND.n6498 240.244
R16537 GND.n6527 GND.n6526 240.244
R16538 GND.n6526 GND.n6525 240.244
R16539 GND.n6525 GND.n6504 240.244
R16540 GND.n6521 GND.n6504 240.244
R16541 GND.n6521 GND.n6520 240.244
R16542 GND.n6520 GND.n6519 240.244
R16543 GND.n6519 GND.n6510 240.244
R16544 GND.n6515 GND.n6510 240.244
R16545 GND.n6515 GND.n3748 240.244
R16546 GND.n6879 GND.n3748 240.244
R16547 GND.n6879 GND.n3749 240.244
R16548 GND.n6812 GND.n3749 240.244
R16549 GND.n6815 GND.n6812 240.244
R16550 GND.n6865 GND.n6815 240.244
R16551 GND.n6865 GND.n6862 240.244
R16552 GND.n6862 GND.n6816 240.244
R16553 GND.n6843 GND.n6816 240.244
R16554 GND.n6844 GND.n6843 240.244
R16555 GND.n6847 GND.n6844 240.244
R16556 GND.n6847 GND.n3736 240.244
R16557 GND.n6886 GND.n3736 240.244
R16558 GND.n6886 GND.n3737 240.244
R16559 GND.n3737 GND.n3719 240.244
R16560 GND.n6904 GND.n3719 240.244
R16561 GND.n6904 GND.n3714 240.244
R16562 GND.n6912 GND.n3714 240.244
R16563 GND.n6912 GND.n3715 240.244
R16564 GND.n3715 GND.n3697 240.244
R16565 GND.n6931 GND.n3697 240.244
R16566 GND.n6931 GND.n3692 240.244
R16567 GND.n6939 GND.n3692 240.244
R16568 GND.n6939 GND.n3693 240.244
R16569 GND.n3693 GND.n3677 240.244
R16570 GND.n6960 GND.n3677 240.244
R16571 GND.n6960 GND.n3672 240.244
R16572 GND.n6968 GND.n3672 240.244
R16573 GND.n6968 GND.n3673 240.244
R16574 GND.n3673 GND.n3655 240.244
R16575 GND.n6987 GND.n3655 240.244
R16576 GND.n6987 GND.n3650 240.244
R16577 GND.n6995 GND.n3650 240.244
R16578 GND.n6995 GND.n3651 240.244
R16579 GND.n3651 GND.n3633 240.244
R16580 GND.n7013 GND.n3633 240.244
R16581 GND.n7013 GND.n3628 240.244
R16582 GND.n7021 GND.n3628 240.244
R16583 GND.n7021 GND.n3629 240.244
R16584 GND.n3629 GND.n3611 240.244
R16585 GND.n7040 GND.n3611 240.244
R16586 GND.n7040 GND.n3606 240.244
R16587 GND.n7048 GND.n3606 240.244
R16588 GND.n7048 GND.n3607 240.244
R16589 GND.n3607 GND.n3590 240.244
R16590 GND.n7068 GND.n3590 240.244
R16591 GND.n7068 GND.n3585 240.244
R16592 GND.n7083 GND.n3585 240.244
R16593 GND.n7083 GND.n3586 240.244
R16594 GND.n7079 GND.n3586 240.244
R16595 GND.n7079 GND.n7078 240.244
R16596 GND.n7078 GND.n580 240.244
R16597 GND.n9498 GND.n580 240.244
R16598 GND.n9498 GND.n581 240.244
R16599 GND.n9494 GND.n581 240.244
R16600 GND.n9494 GND.n9493 240.244
R16601 GND.n9493 GND.n9492 240.244
R16602 GND.n9492 GND.n587 240.244
R16603 GND.n9488 GND.n587 240.244
R16604 GND.n9488 GND.n9487 240.244
R16605 GND.n9487 GND.n9486 240.244
R16606 GND.n9486 GND.n593 240.244
R16607 GND.n9482 GND.n593 240.244
R16608 GND.n9482 GND.n599 240.244
R16609 GND.n9478 GND.n599 240.244
R16610 GND.n9478 GND.n601 240.244
R16611 GND.n9474 GND.n601 240.244
R16612 GND.n9474 GND.n607 240.244
R16613 GND.n9470 GND.n607 240.244
R16614 GND.n9470 GND.n609 240.244
R16615 GND.n9466 GND.n609 240.244
R16616 GND.n9466 GND.n615 240.244
R16617 GND.n9462 GND.n615 240.244
R16618 GND.n8285 GND.n1323 240.244
R16619 GND.n8281 GND.n1323 240.244
R16620 GND.n8281 GND.n1325 240.244
R16621 GND.n8277 GND.n1325 240.244
R16622 GND.n8277 GND.n1330 240.244
R16623 GND.n8273 GND.n1330 240.244
R16624 GND.n8273 GND.n1332 240.244
R16625 GND.n8269 GND.n1332 240.244
R16626 GND.n8269 GND.n1338 240.244
R16627 GND.n8265 GND.n1338 240.244
R16628 GND.n8265 GND.n1340 240.244
R16629 GND.n8261 GND.n1340 240.244
R16630 GND.n8261 GND.n1346 240.244
R16631 GND.n8257 GND.n1346 240.244
R16632 GND.n8257 GND.n1348 240.244
R16633 GND.n8253 GND.n1348 240.244
R16634 GND.n8253 GND.n1354 240.244
R16635 GND.n8249 GND.n1354 240.244
R16636 GND.n8249 GND.n1356 240.244
R16637 GND.n8245 GND.n1356 240.244
R16638 GND.n8245 GND.n1362 240.244
R16639 GND.n8241 GND.n1362 240.244
R16640 GND.n8241 GND.n1364 240.244
R16641 GND.n8237 GND.n1364 240.244
R16642 GND.n8237 GND.n1370 240.244
R16643 GND.n8233 GND.n1370 240.244
R16644 GND.n8233 GND.n1372 240.244
R16645 GND.n8229 GND.n1372 240.244
R16646 GND.n8229 GND.n1378 240.244
R16647 GND.n8225 GND.n1378 240.244
R16648 GND.n8225 GND.n1380 240.244
R16649 GND.n8221 GND.n1380 240.244
R16650 GND.n8221 GND.n1386 240.244
R16651 GND.n8217 GND.n1386 240.244
R16652 GND.n8217 GND.n1388 240.244
R16653 GND.n8213 GND.n1388 240.244
R16654 GND.n8213 GND.n1394 240.244
R16655 GND.n8209 GND.n1394 240.244
R16656 GND.n8209 GND.n1396 240.244
R16657 GND.n8205 GND.n1396 240.244
R16658 GND.n8205 GND.n1402 240.244
R16659 GND.n8201 GND.n1402 240.244
R16660 GND.n8201 GND.n1404 240.244
R16661 GND.n8197 GND.n1404 240.244
R16662 GND.n8197 GND.n1410 240.244
R16663 GND.n8193 GND.n1410 240.244
R16664 GND.n8193 GND.n1412 240.244
R16665 GND.n8189 GND.n1412 240.244
R16666 GND.n8189 GND.n1418 240.244
R16667 GND.n8185 GND.n1418 240.244
R16668 GND.n8185 GND.n1420 240.244
R16669 GND.n8181 GND.n1420 240.244
R16670 GND.n8181 GND.n1426 240.244
R16671 GND.n8177 GND.n1426 240.244
R16672 GND.n7292 GND.n3314 240.244
R16673 GND.n3325 GND.n3324 240.244
R16674 GND.n3327 GND.n3326 240.244
R16675 GND.n3335 GND.n3334 240.244
R16676 GND.n3343 GND.n3342 240.244
R16677 GND.n3345 GND.n3344 240.244
R16678 GND.n3370 GND.n3313 240.244
R16679 GND.n7249 GND.n3370 240.244
R16680 GND.n7249 GND.n3371 240.244
R16681 GND.n6581 GND.n3371 240.244
R16682 GND.n6581 GND.n3961 240.244
R16683 GND.n3961 GND.n3950 240.244
R16684 GND.n6604 GND.n3950 240.244
R16685 GND.n6608 GND.n6604 240.244
R16686 GND.n6608 GND.n6607 240.244
R16687 GND.n6607 GND.n3939 240.244
R16688 GND.n3939 GND.n3929 240.244
R16689 GND.n6629 GND.n3929 240.244
R16690 GND.n6632 GND.n6629 240.244
R16691 GND.n6632 GND.n6631 240.244
R16692 GND.n6631 GND.n3916 240.244
R16693 GND.n3916 GND.n3904 240.244
R16694 GND.n6653 GND.n3904 240.244
R16695 GND.n6657 GND.n6653 240.244
R16696 GND.n6657 GND.n6656 240.244
R16697 GND.n6656 GND.n3892 240.244
R16698 GND.n3892 GND.n3882 240.244
R16699 GND.n6678 GND.n3882 240.244
R16700 GND.n6682 GND.n6678 240.244
R16701 GND.n6682 GND.n6680 240.244
R16702 GND.n6680 GND.n3871 240.244
R16703 GND.n3871 GND.n3859 240.244
R16704 GND.n6703 GND.n3859 240.244
R16705 GND.n6707 GND.n6703 240.244
R16706 GND.n6707 GND.n6706 240.244
R16707 GND.n6706 GND.n3848 240.244
R16708 GND.n3848 GND.n3838 240.244
R16709 GND.n6728 GND.n3838 240.244
R16710 GND.n6731 GND.n6728 240.244
R16711 GND.n6731 GND.n6730 240.244
R16712 GND.n6730 GND.n3825 240.244
R16713 GND.n3825 GND.n3813 240.244
R16714 GND.n6752 GND.n3813 240.244
R16715 GND.n6756 GND.n6752 240.244
R16716 GND.n6756 GND.n6755 240.244
R16717 GND.n6755 GND.n3801 240.244
R16718 GND.n3801 GND.n3791 240.244
R16719 GND.n6777 GND.n3791 240.244
R16720 GND.n6781 GND.n6777 240.244
R16721 GND.n6781 GND.n6779 240.244
R16722 GND.n6779 GND.n3776 240.244
R16723 GND.n3781 GND.n3776 240.244
R16724 GND.n3781 GND.n3780 240.244
R16725 GND.n3780 GND.n3753 240.244
R16726 GND.n3762 GND.n3753 240.244
R16727 GND.n6869 GND.n3762 240.244
R16728 GND.n6869 GND.n6868 240.244
R16729 GND.n6868 GND.n3763 240.244
R16730 GND.n6819 GND.n3763 240.244
R16731 GND.n6829 GND.n6819 240.244
R16732 GND.n6852 GND.n6829 240.244
R16733 GND.n6852 GND.n6850 240.244
R16734 GND.n6850 GND.n6830 240.244
R16735 GND.n6830 GND.n3733 240.244
R16736 GND.n6889 GND.n3733 240.244
R16737 GND.n6891 GND.n6889 240.244
R16738 GND.n6891 GND.n6890 240.244
R16739 GND.n6890 GND.n3723 240.244
R16740 GND.n3723 GND.n3712 240.244
R16741 GND.n6916 GND.n3712 240.244
R16742 GND.n6918 GND.n6916 240.244
R16743 GND.n6918 GND.n6917 240.244
R16744 GND.n6917 GND.n3701 240.244
R16745 GND.n3701 GND.n3689 240.244
R16746 GND.n6943 GND.n3689 240.244
R16747 GND.n6947 GND.n6943 240.244
R16748 GND.n6947 GND.n6946 240.244
R16749 GND.n6946 GND.n3680 240.244
R16750 GND.n3680 GND.n3669 240.244
R16751 GND.n6971 GND.n3669 240.244
R16752 GND.n6974 GND.n6971 240.244
R16753 GND.n6974 GND.n6972 240.244
R16754 GND.n6972 GND.n3660 240.244
R16755 GND.n3660 GND.n3647 240.244
R16756 GND.n6998 GND.n3647 240.244
R16757 GND.n7000 GND.n6998 240.244
R16758 GND.n7000 GND.n6999 240.244
R16759 GND.n6999 GND.n3637 240.244
R16760 GND.n3637 GND.n3626 240.244
R16761 GND.n7025 GND.n3626 240.244
R16762 GND.n7027 GND.n7025 240.244
R16763 GND.n7027 GND.n7026 240.244
R16764 GND.n7026 GND.n3615 240.244
R16765 GND.n3615 GND.n3603 240.244
R16766 GND.n7052 GND.n3603 240.244
R16767 GND.n7055 GND.n7052 240.244
R16768 GND.n7055 GND.n7054 240.244
R16769 GND.n7054 GND.n3594 240.244
R16770 GND.n3594 GND.n3582 240.244
R16771 GND.n7086 GND.n3582 240.244
R16772 GND.n7088 GND.n7086 240.244
R16773 GND.n7088 GND.n3568 240.244
R16774 GND.n7100 GND.n3568 240.244
R16775 GND.n7101 GND.n7100 240.244
R16776 GND.n7101 GND.n571 240.244
R16777 GND.n9505 GND.n571 240.244
R16778 GND.n9505 GND.n573 240.244
R16779 GND.n573 GND.n559 240.244
R16780 GND.n559 GND.n552 240.244
R16781 GND.n9523 GND.n552 240.244
R16782 GND.n9523 GND.n479 240.244
R16783 GND.n9566 GND.n545 240.244
R16784 GND.n9532 GND.n9531 240.244
R16785 GND.n9534 GND.n9533 240.244
R16786 GND.n9538 GND.n9537 240.244
R16787 GND.n9540 GND.n9539 240.244
R16788 GND.n9546 GND.n9543 240.244
R16789 GND.n7257 GND.n3354 240.244
R16790 GND.n3368 GND.n3354 240.244
R16791 GND.n6436 GND.n3368 240.244
R16792 GND.n6436 GND.n3957 240.244
R16793 GND.n6595 GND.n3957 240.244
R16794 GND.n6595 GND.n3952 240.244
R16795 GND.n6602 GND.n3952 240.244
R16796 GND.n6602 GND.n3948 240.244
R16797 GND.n3948 GND.n3936 240.244
R16798 GND.n6620 GND.n3936 240.244
R16799 GND.n6620 GND.n3931 240.244
R16800 GND.n6627 GND.n3931 240.244
R16801 GND.n6627 GND.n3926 240.244
R16802 GND.n3926 GND.n3912 240.244
R16803 GND.n6644 GND.n3912 240.244
R16804 GND.n6644 GND.n3907 240.244
R16805 GND.n6651 GND.n3907 240.244
R16806 GND.n6651 GND.n3902 240.244
R16807 GND.n3902 GND.n3889 240.244
R16808 GND.n6669 GND.n3889 240.244
R16809 GND.n6669 GND.n3884 240.244
R16810 GND.n6676 GND.n3884 240.244
R16811 GND.n6676 GND.n3880 240.244
R16812 GND.n3880 GND.n3867 240.244
R16813 GND.n6694 GND.n3867 240.244
R16814 GND.n6694 GND.n3862 240.244
R16815 GND.n6701 GND.n3862 240.244
R16816 GND.n6701 GND.n3857 240.244
R16817 GND.n3857 GND.n3845 240.244
R16818 GND.n6719 GND.n3845 240.244
R16819 GND.n6719 GND.n3840 240.244
R16820 GND.n6726 GND.n3840 240.244
R16821 GND.n6726 GND.n3835 240.244
R16822 GND.n3835 GND.n3821 240.244
R16823 GND.n6743 GND.n3821 240.244
R16824 GND.n6743 GND.n3816 240.244
R16825 GND.n6750 GND.n3816 240.244
R16826 GND.n6750 GND.n3811 240.244
R16827 GND.n3811 GND.n3798 240.244
R16828 GND.n6768 GND.n3798 240.244
R16829 GND.n6768 GND.n3793 240.244
R16830 GND.n6775 GND.n3793 240.244
R16831 GND.n6775 GND.n3789 240.244
R16832 GND.n3789 GND.n3771 240.244
R16833 GND.n6794 GND.n3771 240.244
R16834 GND.n6794 GND.n3772 240.244
R16835 GND.n3772 GND.n3768 240.244
R16836 GND.n3768 GND.n3751 240.244
R16837 GND.n6803 GND.n3751 240.244
R16838 GND.n6803 GND.n3760 240.244
R16839 GND.n6809 GND.n3760 240.244
R16840 GND.n6810 GND.n6809 240.244
R16841 GND.n6810 GND.n409 240.244
R16842 GND.n410 GND.n409 240.244
R16843 GND.n411 GND.n410 240.244
R16844 GND.n6831 GND.n411 240.244
R16845 GND.n6831 GND.n414 240.244
R16846 GND.n415 GND.n414 240.244
R16847 GND.n416 GND.n415 240.244
R16848 GND.n3731 GND.n416 240.244
R16849 GND.n3731 GND.n419 240.244
R16850 GND.n420 GND.n419 240.244
R16851 GND.n421 GND.n420 240.244
R16852 GND.n6914 GND.n421 240.244
R16853 GND.n6914 GND.n424 240.244
R16854 GND.n425 GND.n424 240.244
R16855 GND.n426 GND.n425 240.244
R16856 GND.n3690 GND.n426 240.244
R16857 GND.n3690 GND.n429 240.244
R16858 GND.n430 GND.n429 240.244
R16859 GND.n431 GND.n430 240.244
R16860 GND.n3678 GND.n431 240.244
R16861 GND.n3678 GND.n434 240.244
R16862 GND.n435 GND.n434 240.244
R16863 GND.n436 GND.n435 240.244
R16864 GND.n3656 GND.n436 240.244
R16865 GND.n3656 GND.n439 240.244
R16866 GND.n440 GND.n439 240.244
R16867 GND.n441 GND.n440 240.244
R16868 GND.n3645 GND.n441 240.244
R16869 GND.n3645 GND.n444 240.244
R16870 GND.n445 GND.n444 240.244
R16871 GND.n446 GND.n445 240.244
R16872 GND.n7023 GND.n446 240.244
R16873 GND.n7023 GND.n449 240.244
R16874 GND.n450 GND.n449 240.244
R16875 GND.n451 GND.n450 240.244
R16876 GND.n3604 GND.n451 240.244
R16877 GND.n3604 GND.n454 240.244
R16878 GND.n455 GND.n454 240.244
R16879 GND.n456 GND.n455 240.244
R16880 GND.n3592 GND.n456 240.244
R16881 GND.n3592 GND.n459 240.244
R16882 GND.n460 GND.n459 240.244
R16883 GND.n461 GND.n460 240.244
R16884 GND.n3579 GND.n461 240.244
R16885 GND.n3579 GND.n464 240.244
R16886 GND.n465 GND.n464 240.244
R16887 GND.n466 GND.n465 240.244
R16888 GND.n569 GND.n466 240.244
R16889 GND.n569 GND.n469 240.244
R16890 GND.n470 GND.n469 240.244
R16891 GND.n471 GND.n470 240.244
R16892 GND.n474 GND.n471 240.244
R16893 GND.n9613 GND.n474 240.244
R16894 GND.n4705 GND.n4704 240.132
R16895 GND.n6206 GND.n6205 240.132
R16896 GND.n9544 GND.t113 225.721
R16897 GND.n497 GND.t147 225.721
R16898 GND.n516 GND.t128 225.721
R16899 GND.n1791 GND.t94 225.721
R16900 GND.n1811 GND.t131 225.721
R16901 GND.n1879 GND.t83 225.721
R16902 GND.n2377 GND.t110 225.721
R16903 GND.n6290 GND.t159 225.721
R16904 GND.n6108 GND.t104 225.721
R16905 GND.n1487 GND.t100 225.721
R16906 GND.n1501 GND.t150 225.721
R16907 GND.n3346 GND.t90 225.721
R16908 GND.n3967 GND.t162 225.243
R16909 GND.n3039 GND.t120 225.243
R16910 GND.n4684 GND.t134 224.03
R16911 GND.n6135 GND.t124 224.03
R16912 GND.n4689 GND.t144 224.03
R16913 GND.n6215 GND.t138 224.03
R16914 GND.n3967 GND.t164 201.439
R16915 GND.n3039 GND.t123 201.439
R16916 GND.n6261 GND.n3298 199.319
R16917 GND.n7874 GND.n1794 199.319
R16918 GND.n4706 GND.n4703 186.49
R16919 GND.n6207 GND.n6204 186.49
R16920 GND.n58 GND.n57 185
R16921 GND.n56 GND.n55 185
R16922 GND.n47 GND.n46 185
R16923 GND.n50 GND.n49 185
R16924 GND.n81 GND.n80 185
R16925 GND.n79 GND.n78 185
R16926 GND.n70 GND.n69 185
R16927 GND.n73 GND.n72 185
R16928 GND.n101 GND.n100 185
R16929 GND.n99 GND.n98 185
R16930 GND.n90 GND.n89 185
R16931 GND.n93 GND.n92 185
R16932 GND.n124 GND.n123 185
R16933 GND.n122 GND.n121 185
R16934 GND.n113 GND.n112 185
R16935 GND.n116 GND.n115 185
R16936 GND.n15 GND.n14 185
R16937 GND.n13 GND.n12 185
R16938 GND.n4 GND.n3 185
R16939 GND.n7 GND.n6 185
R16940 GND.n38 GND.n37 185
R16941 GND.n36 GND.n35 185
R16942 GND.n27 GND.n26 185
R16943 GND.n30 GND.n29 185
R16944 GND.n313 GND.n312 185
R16945 GND.n311 GND.n310 185
R16946 GND.n302 GND.n301 185
R16947 GND.n305 GND.n304 185
R16948 GND.n290 GND.n289 185
R16949 GND.n288 GND.n287 185
R16950 GND.n279 GND.n278 185
R16951 GND.n282 GND.n281 185
R16952 GND.n356 GND.n355 185
R16953 GND.n354 GND.n353 185
R16954 GND.n345 GND.n344 185
R16955 GND.n348 GND.n347 185
R16956 GND.n333 GND.n332 185
R16957 GND.n331 GND.n330 185
R16958 GND.n322 GND.n321 185
R16959 GND.n325 GND.n324 185
R16960 GND.n400 GND.n399 185
R16961 GND.n398 GND.n397 185
R16962 GND.n389 GND.n388 185
R16963 GND.n392 GND.n391 185
R16964 GND.n377 GND.n376 185
R16965 GND.n375 GND.n374 185
R16966 GND.n366 GND.n365 185
R16967 GND.n369 GND.n368 185
R16968 GND.n198 GND.n197 185
R16969 GND.n196 GND.n195 185
R16970 GND.n186 GND.n185 185
R16971 GND.n184 GND.n183 185
R16972 GND.n174 GND.n173 185
R16973 GND.n172 GND.n171 185
R16974 GND.n162 GND.n161 185
R16975 GND.n160 GND.n159 185
R16976 GND.n150 GND.n149 185
R16977 GND.n148 GND.n147 185
R16978 GND.n139 GND.n138 185
R16979 GND.n137 GND.n136 185
R16980 GND.n269 GND.n268 185
R16981 GND.n267 GND.n266 185
R16982 GND.n257 GND.n256 185
R16983 GND.n255 GND.n254 185
R16984 GND.n245 GND.n244 185
R16985 GND.n243 GND.n242 185
R16986 GND.n233 GND.n232 185
R16987 GND.n231 GND.n230 185
R16988 GND.n221 GND.n220 185
R16989 GND.n219 GND.n218 185
R16990 GND.n210 GND.n209 185
R16991 GND.n208 GND.n207 185
R16992 GND.n6256 GND.n6194 163.367
R16993 GND.n6252 GND.n6251 163.367
R16994 GND.n6248 GND.n6247 163.367
R16995 GND.n6244 GND.n6243 163.367
R16996 GND.n6240 GND.n6239 163.367
R16997 GND.n6236 GND.n6235 163.367
R16998 GND.n6232 GND.n6231 163.367
R16999 GND.n6228 GND.n6227 163.367
R17000 GND.n6224 GND.n6223 163.367
R17001 GND.n6219 GND.n6218 163.367
R17002 GND.n6259 GND.n6123 163.367
R17003 GND.n6182 GND.n6181 163.367
R17004 GND.n6178 GND.n6177 163.367
R17005 GND.n6174 GND.n6173 163.367
R17006 GND.n6170 GND.n6169 163.367
R17007 GND.n6166 GND.n6165 163.367
R17008 GND.n6162 GND.n6161 163.367
R17009 GND.n6158 GND.n6157 163.367
R17010 GND.n6154 GND.n6153 163.367
R17011 GND.n6150 GND.n6149 163.367
R17012 GND.n6146 GND.n6145 163.367
R17013 GND.n4809 GND.n2965 163.367
R17014 GND.n4813 GND.n2965 163.367
R17015 GND.n4813 GND.n2972 163.367
R17016 GND.n4817 GND.n2972 163.367
R17017 GND.n4821 GND.n4817 163.367
R17018 GND.n4822 GND.n4821 163.367
R17019 GND.n4822 GND.n2982 163.367
R17020 GND.n4825 GND.n2982 163.367
R17021 GND.n4825 GND.n2990 163.367
R17022 GND.n4829 GND.n2990 163.367
R17023 GND.n4830 GND.n4829 163.367
R17024 GND.n4831 GND.n4830 163.367
R17025 GND.n4831 GND.n3000 163.367
R17026 GND.n4834 GND.n3000 163.367
R17027 GND.n4834 GND.n3010 163.367
R17028 GND.n4670 GND.n3010 163.367
R17029 GND.n4847 GND.n4670 163.367
R17030 GND.n4847 GND.n4671 163.367
R17031 GND.n4843 GND.n4671 163.367
R17032 GND.n4843 GND.n4659 163.367
R17033 GND.n4840 GND.n4659 163.367
R17034 GND.n4840 GND.n4653 163.367
R17035 GND.n4653 GND.n4645 163.367
R17036 GND.n4914 GND.n4645 163.367
R17037 GND.n4914 GND.n4643 163.367
R17038 GND.n4918 GND.n4643 163.367
R17039 GND.n4918 GND.n4634 163.367
R17040 GND.n4929 GND.n4634 163.367
R17041 GND.n4929 GND.n4631 163.367
R17042 GND.n4935 GND.n4631 163.367
R17043 GND.n4935 GND.n4632 163.367
R17044 GND.n4632 GND.n4618 163.367
R17045 GND.n4618 GND.n4610 163.367
R17046 GND.n4954 GND.n4610 163.367
R17047 GND.n4954 GND.n4607 163.367
R17048 GND.n4976 GND.n4607 163.367
R17049 GND.n4976 GND.n4608 163.367
R17050 GND.n4608 GND.n4600 163.367
R17051 GND.n4971 GND.n4600 163.367
R17052 GND.n4971 GND.n4969 163.367
R17053 GND.n4969 GND.n4968 163.367
R17054 GND.n4968 GND.n4958 163.367
R17055 GND.n4958 GND.n4583 163.367
R17056 GND.n4963 GND.n4583 163.367
R17057 GND.n4963 GND.n4577 163.367
R17058 GND.n4960 GND.n4577 163.367
R17059 GND.n4960 GND.n4567 163.367
R17060 GND.n4567 GND.n4558 163.367
R17061 GND.n5077 GND.n4558 163.367
R17062 GND.n5077 GND.n4556 163.367
R17063 GND.n5081 GND.n4556 163.367
R17064 GND.n5081 GND.n4549 163.367
R17065 GND.n5090 GND.n4549 163.367
R17066 GND.n5090 GND.n4546 163.367
R17067 GND.n5100 GND.n4546 163.367
R17068 GND.n5100 GND.n4547 163.367
R17069 GND.n4547 GND.n4538 163.367
R17070 GND.n5095 GND.n4538 163.367
R17071 GND.n5095 GND.n4528 163.367
R17072 GND.n4528 GND.n4521 163.367
R17073 GND.n5124 GND.n4521 163.367
R17074 GND.n5125 GND.n5124 163.367
R17075 GND.n5125 GND.n4512 163.367
R17076 GND.n5129 GND.n4512 163.367
R17077 GND.n5129 GND.n4518 163.367
R17078 GND.n5142 GND.n4518 163.367
R17079 GND.n5142 GND.n4519 163.367
R17080 GND.n4519 GND.n4497 163.367
R17081 GND.n5137 GND.n4497 163.367
R17082 GND.n5137 GND.n4492 163.367
R17083 GND.n5134 GND.n4492 163.367
R17084 GND.n5134 GND.n4481 163.367
R17085 GND.n4481 GND.n4473 163.367
R17086 GND.n5237 GND.n4473 163.367
R17087 GND.n5237 GND.n4471 163.367
R17088 GND.n5241 GND.n4471 163.367
R17089 GND.n5241 GND.n4462 163.367
R17090 GND.n5252 GND.n4462 163.367
R17091 GND.n5252 GND.n4458 163.367
R17092 GND.n5258 GND.n4458 163.367
R17093 GND.n5258 GND.n4460 163.367
R17094 GND.n4460 GND.n4447 163.367
R17095 GND.n4447 GND.n4438 163.367
R17096 GND.n5277 GND.n4438 163.367
R17097 GND.n5277 GND.n4435 163.367
R17098 GND.n5301 GND.n4435 163.367
R17099 GND.n5301 GND.n4436 163.367
R17100 GND.n4436 GND.n4429 163.367
R17101 GND.n5296 GND.n4429 163.367
R17102 GND.n5296 GND.n5293 163.367
R17103 GND.n5293 GND.n5292 163.367
R17104 GND.n5292 GND.n5281 163.367
R17105 GND.n5281 GND.n4411 163.367
R17106 GND.n5287 GND.n4411 163.367
R17107 GND.n5287 GND.n4406 163.367
R17108 GND.n5284 GND.n4406 163.367
R17109 GND.n5284 GND.n4396 163.367
R17110 GND.n4396 GND.n4387 163.367
R17111 GND.n5399 GND.n4387 163.367
R17112 GND.n5399 GND.n4385 163.367
R17113 GND.n5403 GND.n4385 163.367
R17114 GND.n5403 GND.n4376 163.367
R17115 GND.n5414 GND.n4376 163.367
R17116 GND.n5414 GND.n4373 163.367
R17117 GND.n5420 GND.n4373 163.367
R17118 GND.n5420 GND.n4374 163.367
R17119 GND.n4374 GND.n4360 163.367
R17120 GND.n4360 GND.n4353 163.367
R17121 GND.n5439 GND.n4353 163.367
R17122 GND.n5439 GND.n4350 163.367
R17123 GND.n5461 GND.n4350 163.367
R17124 GND.n5461 GND.n4351 163.367
R17125 GND.n4351 GND.n4342 163.367
R17126 GND.n5456 GND.n4342 163.367
R17127 GND.n5456 GND.n5454 163.367
R17128 GND.n5454 GND.n5453 163.367
R17129 GND.n5453 GND.n5443 163.367
R17130 GND.n5443 GND.n4325 163.367
R17131 GND.n5448 GND.n4325 163.367
R17132 GND.n5448 GND.n4319 163.367
R17133 GND.n5445 GND.n4319 163.367
R17134 GND.n5445 GND.n4309 163.367
R17135 GND.n4309 GND.n4301 163.367
R17136 GND.n5570 GND.n4301 163.367
R17137 GND.n5570 GND.n4299 163.367
R17138 GND.n5574 GND.n4299 163.367
R17139 GND.n5574 GND.n4291 163.367
R17140 GND.n5585 GND.n4291 163.367
R17141 GND.n5585 GND.n4288 163.367
R17142 GND.n5591 GND.n4288 163.367
R17143 GND.n5591 GND.n4289 163.367
R17144 GND.n4289 GND.n4276 163.367
R17145 GND.n4276 GND.n4267 163.367
R17146 GND.n5610 GND.n4267 163.367
R17147 GND.n5610 GND.n4264 163.367
R17148 GND.n5621 GND.n4264 163.367
R17149 GND.n5621 GND.n4265 163.367
R17150 GND.n4265 GND.n4258 163.367
R17151 GND.n5616 GND.n4258 163.367
R17152 GND.n5616 GND.n4248 163.367
R17153 GND.n4248 GND.n4243 163.367
R17154 GND.n5646 GND.n4243 163.367
R17155 GND.n5647 GND.n5646 163.367
R17156 GND.n5647 GND.n4234 163.367
R17157 GND.n5651 GND.n4234 163.367
R17158 GND.n5651 GND.n4240 163.367
R17159 GND.n5675 GND.n4240 163.367
R17160 GND.n5675 GND.n4241 163.367
R17161 GND.n4241 GND.n4219 163.367
R17162 GND.n5670 GND.n4219 163.367
R17163 GND.n5670 GND.n4211 163.367
R17164 GND.n5667 GND.n4211 163.367
R17165 GND.n5667 GND.n5666 163.367
R17166 GND.n5666 GND.n5665 163.367
R17167 GND.n5665 GND.n5655 163.367
R17168 GND.n5655 GND.n4195 163.367
R17169 GND.n5660 GND.n4195 163.367
R17170 GND.n5660 GND.n4188 163.367
R17171 GND.n5657 GND.n4188 163.367
R17172 GND.n5657 GND.n4177 163.367
R17173 GND.n4177 GND.n4169 163.367
R17174 GND.n5828 GND.n4169 163.367
R17175 GND.n5828 GND.n4167 163.367
R17176 GND.n5833 GND.n4167 163.367
R17177 GND.n5833 GND.n4159 163.367
R17178 GND.n5842 GND.n4159 163.367
R17179 GND.n5843 GND.n5842 163.367
R17180 GND.n5843 GND.n4156 163.367
R17181 GND.n5851 GND.n4156 163.367
R17182 GND.n5851 GND.n4150 163.367
R17183 GND.n5847 GND.n4150 163.367
R17184 GND.n5847 GND.n4140 163.367
R17185 GND.n4140 GND.n4132 163.367
R17186 GND.n5885 GND.n4132 163.367
R17187 GND.n5885 GND.n4130 163.367
R17188 GND.n5889 GND.n4130 163.367
R17189 GND.n5889 GND.n4121 163.367
R17190 GND.n5900 GND.n4121 163.367
R17191 GND.n5900 GND.n4118 163.367
R17192 GND.n5906 GND.n4118 163.367
R17193 GND.n5906 GND.n4119 163.367
R17194 GND.n4119 GND.n4105 163.367
R17195 GND.n4105 GND.n4097 163.367
R17196 GND.n5925 GND.n4097 163.367
R17197 GND.n5925 GND.n4094 163.367
R17198 GND.n5947 GND.n4094 163.367
R17199 GND.n5947 GND.n4095 163.367
R17200 GND.n4095 GND.n4087 163.367
R17201 GND.n5942 GND.n4087 163.367
R17202 GND.n5942 GND.n5940 163.367
R17203 GND.n5940 GND.n5939 163.367
R17204 GND.n5939 GND.n5929 163.367
R17205 GND.n5929 GND.n4069 163.367
R17206 GND.n5934 GND.n4069 163.367
R17207 GND.n5934 GND.n4063 163.367
R17208 GND.n5931 GND.n4063 163.367
R17209 GND.n5931 GND.n4053 163.367
R17210 GND.n4053 GND.n4044 163.367
R17211 GND.n6036 GND.n4044 163.367
R17212 GND.n6036 GND.n4042 163.367
R17213 GND.n6040 GND.n4042 163.367
R17214 GND.n6040 GND.n4034 163.367
R17215 GND.n6049 GND.n4034 163.367
R17216 GND.n6049 GND.n4031 163.367
R17217 GND.n6072 GND.n4031 163.367
R17218 GND.n6072 GND.n4032 163.367
R17219 GND.n4032 GND.n4022 163.367
R17220 GND.n6067 GND.n4022 163.367
R17221 GND.n6067 GND.n6065 163.367
R17222 GND.n6065 GND.n6064 163.367
R17223 GND.n6064 GND.n6053 163.367
R17224 GND.n6053 GND.n4005 163.367
R17225 GND.n6059 GND.n4005 163.367
R17226 GND.n6059 GND.n4000 163.367
R17227 GND.n6056 GND.n4000 163.367
R17228 GND.n6056 GND.n3990 163.367
R17229 GND.n3990 GND.n3982 163.367
R17230 GND.n6370 GND.n3982 163.367
R17231 GND.n6370 GND.n3979 163.367
R17232 GND.n6392 GND.n3979 163.367
R17233 GND.n6392 GND.n3980 163.367
R17234 GND.n6388 GND.n3980 163.367
R17235 GND.n6388 GND.n3974 163.367
R17236 GND.n6385 GND.n3974 163.367
R17237 GND.n6385 GND.n3242 163.367
R17238 GND.n6382 GND.n3242 163.367
R17239 GND.n6382 GND.n3250 163.367
R17240 GND.n6379 GND.n3250 163.367
R17241 GND.n6379 GND.n3260 163.367
R17242 GND.n7320 GND.n3260 163.367
R17243 GND.n7320 GND.n3261 163.367
R17244 GND.n7316 GND.n3261 163.367
R17245 GND.n7316 GND.n3264 163.367
R17246 GND.n3272 GND.n3264 163.367
R17247 GND.n6141 GND.n3272 163.367
R17248 GND.n4723 GND.n4698 163.367
R17249 GND.n4727 GND.n4698 163.367
R17250 GND.n4731 GND.n4729 163.367
R17251 GND.n4735 GND.n4696 163.367
R17252 GND.n4739 GND.n4737 163.367
R17253 GND.n4743 GND.n4694 163.367
R17254 GND.n4747 GND.n4745 163.367
R17255 GND.n4751 GND.n4692 163.367
R17256 GND.n4755 GND.n4753 163.367
R17257 GND.n4760 GND.n4688 163.367
R17258 GND.n4763 GND.n4762 163.367
R17259 GND.n4769 GND.n4767 163.367
R17260 GND.n4774 GND.n4683 163.367
R17261 GND.n4778 GND.n4776 163.367
R17262 GND.n4782 GND.n4681 163.367
R17263 GND.n4786 GND.n4784 163.367
R17264 GND.n4790 GND.n4679 163.367
R17265 GND.n4794 GND.n4792 163.367
R17266 GND.n4798 GND.n4677 163.367
R17267 GND.n4802 GND.n4800 163.367
R17268 GND.n4806 GND.n4675 163.367
R17269 GND.n7593 GND.n2966 163.367
R17270 GND.n7593 GND.n2967 163.367
R17271 GND.n7589 GND.n2967 163.367
R17272 GND.n7589 GND.n2970 163.367
R17273 GND.n4819 GND.n2970 163.367
R17274 GND.n4819 GND.n2984 163.367
R17275 GND.n7579 GND.n2984 163.367
R17276 GND.n7579 GND.n2985 163.367
R17277 GND.n7575 GND.n2985 163.367
R17278 GND.n7575 GND.n2988 163.367
R17279 GND.n3004 GND.n2988 163.367
R17280 GND.n3004 GND.n3002 163.367
R17281 GND.n7565 GND.n3002 163.367
R17282 GND.n7565 GND.n3003 163.367
R17283 GND.n7561 GND.n3003 163.367
R17284 GND.n7561 GND.n3008 163.367
R17285 GND.n4849 GND.n3008 163.367
R17286 GND.n4850 GND.n4849 163.367
R17287 GND.n4850 GND.n4660 163.367
R17288 GND.n4854 GND.n4660 163.367
R17289 GND.n4854 GND.n4651 163.367
R17290 GND.n4908 GND.n4651 163.367
R17291 GND.n4908 GND.n4649 163.367
R17292 GND.n4912 GND.n4649 163.367
R17293 GND.n4912 GND.n4640 163.367
R17294 GND.n4921 GND.n4640 163.367
R17295 GND.n4921 GND.n4637 163.367
R17296 GND.n4927 GND.n4637 163.367
R17297 GND.n4927 GND.n4638 163.367
R17298 GND.n4638 GND.n4628 163.367
R17299 GND.n4628 GND.n4615 163.367
R17300 GND.n4948 GND.n4615 163.367
R17301 GND.n4948 GND.n4613 163.367
R17302 GND.n4952 GND.n4613 163.367
R17303 GND.n4952 GND.n4605 163.367
R17304 GND.n4978 GND.n4605 163.367
R17305 GND.n4978 GND.n4602 163.367
R17306 GND.n4987 GND.n4602 163.367
R17307 GND.n4987 GND.n4603 163.367
R17308 GND.n4983 GND.n4603 163.367
R17309 GND.n4983 GND.n4982 163.367
R17310 GND.n4982 GND.n4581 163.367
R17311 GND.n5044 GND.n4581 163.367
R17312 GND.n5044 GND.n4579 163.367
R17313 GND.n5048 GND.n4579 163.367
R17314 GND.n5048 GND.n4565 163.367
R17315 GND.n5071 GND.n4565 163.367
R17316 GND.n5071 GND.n4563 163.367
R17317 GND.n5075 GND.n4563 163.367
R17318 GND.n5075 GND.n4554 163.367
R17319 GND.n5084 GND.n4554 163.367
R17320 GND.n5084 GND.n4552 163.367
R17321 GND.n5088 GND.n4552 163.367
R17322 GND.n5088 GND.n4542 163.367
R17323 GND.n5102 GND.n4542 163.367
R17324 GND.n5102 GND.n4540 163.367
R17325 GND.n5106 GND.n4540 163.367
R17326 GND.n5106 GND.n4526 163.367
R17327 GND.n5118 GND.n4526 163.367
R17328 GND.n5118 GND.n4524 163.367
R17329 GND.n5122 GND.n4524 163.367
R17330 GND.n5122 GND.n4514 163.367
R17331 GND.n5151 GND.n4514 163.367
R17332 GND.n5151 GND.n4515 163.367
R17333 GND.n5147 GND.n4515 163.367
R17334 GND.n5147 GND.n5146 163.367
R17335 GND.n5146 GND.n4495 163.367
R17336 GND.n5207 GND.n4495 163.367
R17337 GND.n5207 GND.n4493 163.367
R17338 GND.n5211 GND.n4493 163.367
R17339 GND.n5211 GND.n4479 163.367
R17340 GND.n5231 GND.n4479 163.367
R17341 GND.n5231 GND.n4477 163.367
R17342 GND.n5235 GND.n4477 163.367
R17343 GND.n5235 GND.n4469 163.367
R17344 GND.n5244 GND.n4469 163.367
R17345 GND.n5244 GND.n4466 163.367
R17346 GND.n5250 GND.n4466 163.367
R17347 GND.n5250 GND.n4467 163.367
R17348 GND.n4467 GND.n4456 163.367
R17349 GND.n4456 GND.n4445 163.367
R17350 GND.n5271 GND.n4445 163.367
R17351 GND.n5271 GND.n4443 163.367
R17352 GND.n5275 GND.n4443 163.367
R17353 GND.n5275 GND.n4433 163.367
R17354 GND.n5303 GND.n4433 163.367
R17355 GND.n5303 GND.n4430 163.367
R17356 GND.n5312 GND.n4430 163.367
R17357 GND.n5312 GND.n4431 163.367
R17358 GND.n5308 GND.n4431 163.367
R17359 GND.n5308 GND.n5307 163.367
R17360 GND.n5307 GND.n4409 163.367
R17361 GND.n5369 GND.n4409 163.367
R17362 GND.n5369 GND.n4407 163.367
R17363 GND.n5373 GND.n4407 163.367
R17364 GND.n5373 GND.n4393 163.367
R17365 GND.n5393 GND.n4393 163.367
R17366 GND.n5393 GND.n4391 163.367
R17367 GND.n5397 GND.n4391 163.367
R17368 GND.n5397 GND.n4383 163.367
R17369 GND.n5406 GND.n4383 163.367
R17370 GND.n5406 GND.n4380 163.367
R17371 GND.n5412 GND.n4380 163.367
R17372 GND.n5412 GND.n4381 163.367
R17373 GND.n4381 GND.n4370 163.367
R17374 GND.n4370 GND.n4359 163.367
R17375 GND.n5433 GND.n4359 163.367
R17376 GND.n5433 GND.n4357 163.367
R17377 GND.n5437 GND.n4357 163.367
R17378 GND.n5437 GND.n4348 163.367
R17379 GND.n5463 GND.n4348 163.367
R17380 GND.n5463 GND.n4345 163.367
R17381 GND.n5472 GND.n4345 163.367
R17382 GND.n5472 GND.n4346 163.367
R17383 GND.n5468 GND.n4346 163.367
R17384 GND.n5468 GND.n5467 163.367
R17385 GND.n5467 GND.n4323 163.367
R17386 GND.n5539 GND.n4323 163.367
R17387 GND.n5539 GND.n4321 163.367
R17388 GND.n5543 GND.n4321 163.367
R17389 GND.n5543 GND.n4307 163.367
R17390 GND.n5564 GND.n4307 163.367
R17391 GND.n5564 GND.n4305 163.367
R17392 GND.n5568 GND.n4305 163.367
R17393 GND.n5568 GND.n4296 163.367
R17394 GND.n5577 GND.n4296 163.367
R17395 GND.n5577 GND.n4293 163.367
R17396 GND.n5583 GND.n4293 163.367
R17397 GND.n5583 GND.n4294 163.367
R17398 GND.n4294 GND.n4285 163.367
R17399 GND.n4285 GND.n4273 163.367
R17400 GND.n5604 GND.n4273 163.367
R17401 GND.n5604 GND.n4271 163.367
R17402 GND.n5608 GND.n4271 163.367
R17403 GND.n5608 GND.n4262 163.367
R17404 GND.n5623 GND.n4262 163.367
R17405 GND.n5623 GND.n4260 163.367
R17406 GND.n5627 GND.n4260 163.367
R17407 GND.n5627 GND.n4247 163.367
R17408 GND.n5640 GND.n4247 163.367
R17409 GND.n5640 GND.n4245 163.367
R17410 GND.n5644 GND.n4245 163.367
R17411 GND.n5644 GND.n4236 163.367
R17412 GND.n5683 GND.n4236 163.367
R17413 GND.n5683 GND.n4237 163.367
R17414 GND.n5679 GND.n4237 163.367
R17415 GND.n5679 GND.n5678 163.367
R17416 GND.n5678 GND.n4217 163.367
R17417 GND.n5709 GND.n4217 163.367
R17418 GND.n5709 GND.n4214 163.367
R17419 GND.n5718 GND.n4214 163.367
R17420 GND.n5718 GND.n4215 163.367
R17421 GND.n5714 GND.n4215 163.367
R17422 GND.n5714 GND.n5713 163.367
R17423 GND.n5713 GND.n4192 163.367
R17424 GND.n5795 GND.n4192 163.367
R17425 GND.n5795 GND.n4190 163.367
R17426 GND.n5799 GND.n4190 163.367
R17427 GND.n5799 GND.n4175 163.367
R17428 GND.n5822 GND.n4175 163.367
R17429 GND.n5822 GND.n4173 163.367
R17430 GND.n5826 GND.n4173 163.367
R17431 GND.n5826 GND.n4165 163.367
R17432 GND.n5836 GND.n4165 163.367
R17433 GND.n5836 GND.n4163 163.367
R17434 GND.n5840 GND.n4163 163.367
R17435 GND.n5840 GND.n4154 163.367
R17436 GND.n5855 GND.n4154 163.367
R17437 GND.n5855 GND.n4152 163.367
R17438 GND.n5859 GND.n4152 163.367
R17439 GND.n5859 GND.n4138 163.367
R17440 GND.n5879 GND.n4138 163.367
R17441 GND.n5879 GND.n4136 163.367
R17442 GND.n5883 GND.n4136 163.367
R17443 GND.n5883 GND.n4128 163.367
R17444 GND.n5892 GND.n4128 163.367
R17445 GND.n5892 GND.n4125 163.367
R17446 GND.n5898 GND.n4125 163.367
R17447 GND.n5898 GND.n4126 163.367
R17448 GND.n4126 GND.n4115 163.367
R17449 GND.n4115 GND.n4103 163.367
R17450 GND.n5919 GND.n4103 163.367
R17451 GND.n5919 GND.n4101 163.367
R17452 GND.n5923 GND.n4101 163.367
R17453 GND.n5923 GND.n4092 163.367
R17454 GND.n5949 GND.n4092 163.367
R17455 GND.n5949 GND.n4089 163.367
R17456 GND.n5958 GND.n4089 163.367
R17457 GND.n5958 GND.n4090 163.367
R17458 GND.n5954 GND.n4090 163.367
R17459 GND.n5954 GND.n5953 163.367
R17460 GND.n5953 GND.n4067 163.367
R17461 GND.n6003 GND.n4067 163.367
R17462 GND.n6003 GND.n4065 163.367
R17463 GND.n6007 GND.n4065 163.367
R17464 GND.n6007 GND.n4050 163.367
R17465 GND.n6030 GND.n4050 163.367
R17466 GND.n6030 GND.n4048 163.367
R17467 GND.n6034 GND.n4048 163.367
R17468 GND.n6034 GND.n4040 163.367
R17469 GND.n6043 GND.n4040 163.367
R17470 GND.n6043 GND.n4038 163.367
R17471 GND.n6047 GND.n4038 163.367
R17472 GND.n6047 GND.n4028 163.367
R17473 GND.n6074 GND.n4028 163.367
R17474 GND.n6074 GND.n4025 163.367
R17475 GND.n6083 GND.n4025 163.367
R17476 GND.n6083 GND.n4026 163.367
R17477 GND.n6079 GND.n4026 163.367
R17478 GND.n6079 GND.n6078 163.367
R17479 GND.n6078 GND.n4003 163.367
R17480 GND.n6343 GND.n4003 163.367
R17481 GND.n6343 GND.n4001 163.367
R17482 GND.n6347 GND.n4001 163.367
R17483 GND.n6347 GND.n3988 163.367
R17484 GND.n6363 GND.n3988 163.367
R17485 GND.n6363 GND.n3986 163.367
R17486 GND.n6368 GND.n3986 163.367
R17487 GND.n6368 GND.n3977 163.367
R17488 GND.n6394 GND.n3977 163.367
R17489 GND.n6395 GND.n6394 163.367
R17490 GND.n6395 GND.n3975 163.367
R17491 GND.n6399 GND.n3975 163.367
R17492 GND.n6399 GND.n3244 163.367
R17493 GND.n7333 GND.n3244 163.367
R17494 GND.n7333 GND.n3245 163.367
R17495 GND.n7329 GND.n3245 163.367
R17496 GND.n7329 GND.n3248 163.367
R17497 GND.n6375 GND.n3248 163.367
R17498 GND.n6375 GND.n3258 163.367
R17499 GND.n3266 GND.n3258 163.367
R17500 GND.n7314 GND.n3266 163.367
R17501 GND.n7314 GND.n3267 163.367
R17502 GND.n7310 GND.n3267 163.367
R17503 GND.n7310 GND.n3270 163.367
R17504 GND.n6213 GND.n6212 156.462
R17505 GND.n154 GND.n142 155.105
R17506 GND.n202 GND.n201 153.631
R17507 GND.n190 GND.n189 153.631
R17508 GND.n178 GND.n177 153.631
R17509 GND.n166 GND.n165 153.631
R17510 GND.n154 GND.n153 153.631
R17511 GND.n4711 GND.n4710 152
R17512 GND.n4712 GND.n4701 152
R17513 GND.n4714 GND.n4713 152
R17514 GND.n4716 GND.n4699 152
R17515 GND.n4718 GND.n4717 152
R17516 GND.n6211 GND.n6195 152
R17517 GND.n6203 GND.n6196 152
R17518 GND.n6202 GND.n6201 152
R17519 GND.n6200 GND.n6197 152
R17520 GND.n194 GND.t25 151.613
R17521 GND.n182 GND.t1 151.613
R17522 GND.n170 GND.t18 151.613
R17523 GND.n158 GND.t5 151.613
R17524 GND.n146 GND.t20 151.613
R17525 GND.n135 GND.t173 151.613
R17526 GND.n265 GND.t22 151.613
R17527 GND.n253 GND.t15 151.613
R17528 GND.n241 GND.t7 151.613
R17529 GND.n229 GND.t30 151.613
R17530 GND.n217 GND.t12 151.613
R17531 GND.n206 GND.t28 151.613
R17532 GND.n6198 GND.t141 150.546
R17533 GND.t45 GND.n48 147.888
R17534 GND.t78 GND.n71 147.888
R17535 GND.t73 GND.n91 147.888
R17536 GND.t61 GND.n114 147.888
R17537 GND.t59 GND.n5 147.888
R17538 GND.t54 GND.n28 147.888
R17539 GND.t50 GND.n303 147.888
R17540 GND.t76 GND.n280 147.888
R17541 GND.t51 GND.n346 147.888
R17542 GND.t64 GND.n323 147.888
R17543 GND.t57 GND.n390 147.888
R17544 GND.t74 GND.n367 147.888
R17545 GND.n6258 GND.n6122 143.351
R17546 GND.n6183 GND.n6122 143.351
R17547 GND.n4765 GND.n4764 143.351
R17548 GND.n4766 GND.n4765 143.351
R17549 GND.n9545 GND.t116 140.606
R17550 GND.n498 GND.t149 140.606
R17551 GND.n517 GND.t130 140.606
R17552 GND.n1792 GND.t96 140.606
R17553 GND.n1812 GND.t133 140.606
R17554 GND.n1880 GND.t86 140.606
R17555 GND.n2378 GND.t111 140.606
R17556 GND.n6291 GND.t160 140.606
R17557 GND.n6109 GND.t105 140.606
R17558 GND.n1488 GND.t102 140.606
R17559 GND.n1502 GND.t151 140.606
R17560 GND.n3347 GND.t92 140.606
R17561 GND.n4685 GND.t136 134.506
R17562 GND.n6136 GND.t127 134.506
R17563 GND.n4690 GND.t145 134.506
R17564 GND.n6216 GND.t140 134.506
R17565 GND.n4708 GND.t80 130.484
R17566 GND.n4717 GND.t107 126.766
R17567 GND.n4715 GND.t156 126.766
R17568 GND.n4701 GND.t97 126.766
R17569 GND.n4709 GND.t117 126.766
R17570 GND.n6199 GND.t166 126.766
R17571 GND.n6201 GND.t153 126.766
R17572 GND.n6210 GND.t169 126.766
R17573 GND.n6212 GND.t87 126.766
R17574 GND.n3968 GND.t165 122.311
R17575 GND.n3040 GND.t122 122.311
R17576 GND.n9545 GND.n9544 121.406
R17577 GND.n498 GND.n497 121.406
R17578 GND.n517 GND.n516 121.406
R17579 GND.n1792 GND.n1791 121.406
R17580 GND.n1812 GND.n1811 121.406
R17581 GND.n1880 GND.n1879 121.406
R17582 GND.n2378 GND.n2377 121.406
R17583 GND.n6291 GND.n6290 121.406
R17584 GND.n6109 GND.n6108 121.406
R17585 GND.n1488 GND.n1487 121.406
R17586 GND.n1502 GND.n1501 121.406
R17587 GND.n3347 GND.n3346 121.406
R17588 GND.n4685 GND.n4684 120.436
R17589 GND.n6136 GND.n6135 120.436
R17590 GND.n4690 GND.n4689 120.436
R17591 GND.n6216 GND.n6215 120.436
R17592 GND.n57 GND.n56 104.615
R17593 GND.n56 GND.n46 104.615
R17594 GND.n49 GND.n46 104.615
R17595 GND.n80 GND.n79 104.615
R17596 GND.n79 GND.n69 104.615
R17597 GND.n72 GND.n69 104.615
R17598 GND.n100 GND.n99 104.615
R17599 GND.n99 GND.n89 104.615
R17600 GND.n92 GND.n89 104.615
R17601 GND.n123 GND.n122 104.615
R17602 GND.n122 GND.n112 104.615
R17603 GND.n115 GND.n112 104.615
R17604 GND.n14 GND.n13 104.615
R17605 GND.n13 GND.n3 104.615
R17606 GND.n6 GND.n3 104.615
R17607 GND.n37 GND.n36 104.615
R17608 GND.n36 GND.n26 104.615
R17609 GND.n29 GND.n26 104.615
R17610 GND.n312 GND.n311 104.615
R17611 GND.n311 GND.n301 104.615
R17612 GND.n304 GND.n301 104.615
R17613 GND.n289 GND.n288 104.615
R17614 GND.n288 GND.n278 104.615
R17615 GND.n281 GND.n278 104.615
R17616 GND.n355 GND.n354 104.615
R17617 GND.n354 GND.n344 104.615
R17618 GND.n347 GND.n344 104.615
R17619 GND.n332 GND.n331 104.615
R17620 GND.n331 GND.n321 104.615
R17621 GND.n324 GND.n321 104.615
R17622 GND.n399 GND.n398 104.615
R17623 GND.n398 GND.n388 104.615
R17624 GND.n391 GND.n388 104.615
R17625 GND.n376 GND.n375 104.615
R17626 GND.n375 GND.n365 104.615
R17627 GND.n368 GND.n365 104.615
R17628 GND.n197 GND.n196 104.615
R17629 GND.n185 GND.n184 104.615
R17630 GND.n173 GND.n172 104.615
R17631 GND.n161 GND.n160 104.615
R17632 GND.n149 GND.n148 104.615
R17633 GND.n138 GND.n137 104.615
R17634 GND.n268 GND.n267 104.615
R17635 GND.n256 GND.n255 104.615
R17636 GND.n244 GND.n243 104.615
R17637 GND.n232 GND.n231 104.615
R17638 GND.n220 GND.n219 104.615
R17639 GND.n209 GND.n208 104.615
R17640 GND.n520 GND.n485 99.6594
R17641 GND.n522 GND.n521 99.6594
R17642 GND.n523 GND.n490 99.6594
R17643 GND.n525 GND.n524 99.6594
R17644 GND.n526 GND.n495 99.6594
R17645 GND.n528 GND.n527 99.6594
R17646 GND.n529 GND.n502 99.6594
R17647 GND.n531 GND.n530 99.6594
R17648 GND.n532 GND.n507 99.6594
R17649 GND.n534 GND.n533 99.6594
R17650 GND.n535 GND.n512 99.6594
R17651 GND.n537 GND.n536 99.6594
R17652 GND.n9569 GND.n9568 99.6594
R17653 GND.n3359 GND.n3292 99.6594
R17654 GND.n6271 GND.n3293 99.6594
R17655 GND.n6275 GND.n3294 99.6594
R17656 GND.n6281 GND.n3295 99.6594
R17657 GND.n6285 GND.n3296 99.6594
R17658 GND.n6261 GND.n3297 99.6594
R17659 GND.n6295 GND.n3299 99.6594
R17660 GND.n6301 GND.n3300 99.6594
R17661 GND.n6305 GND.n3301 99.6594
R17662 GND.n6311 GND.n3302 99.6594
R17663 GND.n6315 GND.n3303 99.6594
R17664 GND.n6112 GND.n3304 99.6594
R17665 GND.n7880 GND.n1781 99.6594
R17666 GND.n7879 GND.n1784 99.6594
R17667 GND.n7877 GND.n1786 99.6594
R17668 GND.n7876 GND.n1789 99.6594
R17669 GND.n1817 GND.n1816 99.6594
R17670 GND.n1818 GND.n1800 99.6594
R17671 GND.n1820 GND.n1819 99.6594
R17672 GND.n1821 GND.n1805 99.6594
R17673 GND.n1823 GND.n1822 99.6594
R17674 GND.n1824 GND.n1810 99.6594
R17675 GND.n7882 GND.n1770 99.6594
R17676 GND.n8150 GND.n8149 99.6594
R17677 GND.n8144 GND.n1452 99.6594
R17678 GND.n8141 GND.n1453 99.6594
R17679 GND.n8137 GND.n1454 99.6594
R17680 GND.n8133 GND.n1455 99.6594
R17681 GND.n8129 GND.n1456 99.6594
R17682 GND.n8125 GND.n1457 99.6594
R17683 GND.n8121 GND.n1458 99.6594
R17684 GND.n8117 GND.n1459 99.6594
R17685 GND.n8113 GND.n1460 99.6594
R17686 GND.n8109 GND.n1461 99.6594
R17687 GND.n8105 GND.n1462 99.6594
R17688 GND.n1856 GND.n1831 99.6594
R17689 GND.n1858 GND.n1830 99.6594
R17690 GND.n1866 GND.n1829 99.6594
R17691 GND.n1876 GND.n1828 99.6594
R17692 GND.n1878 GND.n1827 99.6594
R17693 GND.n7836 GND.n1826 99.6594
R17694 GND.n8096 GND.n1471 99.6594
R17695 GND.n2388 GND.n1470 99.6594
R17696 GND.n2393 GND.n1469 99.6594
R17697 GND.n2385 GND.n1468 99.6594
R17698 GND.n2401 GND.n1467 99.6594
R17699 GND.n2381 GND.n1466 99.6594
R17700 GND.n6402 GND.n3320 99.6594
R17701 GND.n6404 GND.n6403 99.6594
R17702 GND.n6405 GND.n3331 99.6594
R17703 GND.n6407 GND.n3338 99.6594
R17704 GND.n6409 GND.n6408 99.6594
R17705 GND.n6410 GND.n3351 99.6594
R17706 GND.n6412 GND.n3964 99.6594
R17707 GND.n6413 GND.n3966 99.6594
R17708 GND.n6414 GND.n3972 99.6594
R17709 GND.n6416 GND.n3229 99.6594
R17710 GND.n7868 GND.n7867 99.6594
R17711 GND.n1850 GND.n1840 99.6594
R17712 GND.n1863 GND.n1841 99.6594
R17713 GND.n1871 GND.n1842 99.6594
R17714 GND.n1873 GND.n1843 99.6594
R17715 GND.n1885 GND.n1844 99.6594
R17716 GND.n3034 GND.n1845 99.6594
R17717 GND.n3038 GND.n1846 99.6594
R17718 GND.n3031 GND.n1847 99.6594
R17719 GND.n7867 GND.n1838 99.6594
R17720 GND.n1862 GND.n1840 99.6594
R17721 GND.n1870 GND.n1841 99.6594
R17722 GND.n1872 GND.n1842 99.6594
R17723 GND.n1884 GND.n1843 99.6594
R17724 GND.n3033 GND.n1844 99.6594
R17725 GND.n3037 GND.n1845 99.6594
R17726 GND.n3030 GND.n1846 99.6594
R17727 GND.n3047 GND.n1847 99.6594
R17728 GND.n6417 GND.n6416 99.6594
R17729 GND.n6414 GND.n3971 99.6594
R17730 GND.n6413 GND.n3965 99.6594
R17731 GND.n6412 GND.n6411 99.6594
R17732 GND.n6410 GND.n3350 99.6594
R17733 GND.n6409 GND.n3339 99.6594
R17734 GND.n6407 GND.n6406 99.6594
R17735 GND.n6405 GND.n3330 99.6594
R17736 GND.n6404 GND.n3321 99.6594
R17737 GND.n6402 GND.n6401 99.6594
R17738 GND.n2387 GND.n1471 99.6594
R17739 GND.n2392 GND.n1470 99.6594
R17740 GND.n2384 GND.n1469 99.6594
R17741 GND.n2400 GND.n1468 99.6594
R17742 GND.n2380 GND.n1467 99.6594
R17743 GND.n2376 GND.n1466 99.6594
R17744 GND.n1881 GND.n1826 99.6594
R17745 GND.n1877 GND.n1827 99.6594
R17746 GND.n1867 GND.n1828 99.6594
R17747 GND.n1859 GND.n1829 99.6594
R17748 GND.n1857 GND.n1830 99.6594
R17749 GND.n1832 GND.n1831 99.6594
R17750 GND.n8150 GND.n1473 99.6594
R17751 GND.n8142 GND.n1452 99.6594
R17752 GND.n8138 GND.n1453 99.6594
R17753 GND.n8134 GND.n1454 99.6594
R17754 GND.n8130 GND.n1455 99.6594
R17755 GND.n8126 GND.n1456 99.6594
R17756 GND.n8122 GND.n1457 99.6594
R17757 GND.n8118 GND.n1458 99.6594
R17758 GND.n8114 GND.n1459 99.6594
R17759 GND.n8110 GND.n1460 99.6594
R17760 GND.n8106 GND.n1461 99.6594
R17761 GND.n1500 GND.n1462 99.6594
R17762 GND.n7883 GND.n7882 99.6594
R17763 GND.n1824 GND.n1809 99.6594
R17764 GND.n1823 GND.n1806 99.6594
R17765 GND.n1821 GND.n1804 99.6594
R17766 GND.n1820 GND.n1801 99.6594
R17767 GND.n1818 GND.n1799 99.6594
R17768 GND.n1817 GND.n1796 99.6594
R17769 GND.n1815 GND.n1794 99.6594
R17770 GND.n7874 GND.n1790 99.6594
R17771 GND.n7876 GND.n7875 99.6594
R17772 GND.n7877 GND.n1785 99.6594
R17773 GND.n7879 GND.n7878 99.6594
R17774 GND.n7880 GND.n1780 99.6594
R17775 GND.n6270 GND.n3292 99.6594
R17776 GND.n6274 GND.n3293 99.6594
R17777 GND.n6280 GND.n3294 99.6594
R17778 GND.n6284 GND.n3295 99.6594
R17779 GND.n6118 GND.n3296 99.6594
R17780 GND.n6294 GND.n3298 99.6594
R17781 GND.n6300 GND.n3299 99.6594
R17782 GND.n6304 GND.n3300 99.6594
R17783 GND.n6310 GND.n3301 99.6594
R17784 GND.n6314 GND.n3302 99.6594
R17785 GND.n6111 GND.n3303 99.6594
R17786 GND.n6107 GND.n3304 99.6594
R17787 GND.n9568 GND.n518 99.6594
R17788 GND.n537 GND.n513 99.6594
R17789 GND.n535 GND.n511 99.6594
R17790 GND.n534 GND.n508 99.6594
R17791 GND.n532 GND.n506 99.6594
R17792 GND.n531 GND.n503 99.6594
R17793 GND.n529 GND.n501 99.6594
R17794 GND.n528 GND.n496 99.6594
R17795 GND.n526 GND.n494 99.6594
R17796 GND.n525 GND.n491 99.6594
R17797 GND.n523 GND.n489 99.6594
R17798 GND.n522 GND.n486 99.6594
R17799 GND.n520 GND.n481 99.6594
R17800 GND.n3314 GND.n3306 99.6594
R17801 GND.n3325 GND.n3307 99.6594
R17802 GND.n3327 GND.n3308 99.6594
R17803 GND.n3335 GND.n3309 99.6594
R17804 GND.n3343 GND.n3310 99.6594
R17805 GND.n3345 GND.n3311 99.6594
R17806 GND.n3324 GND.n3306 99.6594
R17807 GND.n3326 GND.n3307 99.6594
R17808 GND.n3334 GND.n3308 99.6594
R17809 GND.n3342 GND.n3309 99.6594
R17810 GND.n3344 GND.n3310 99.6594
R17811 GND.n7258 GND.n3311 99.6594
R17812 GND.n545 GND.n538 99.6594
R17813 GND.n9532 GND.n539 99.6594
R17814 GND.n9534 GND.n540 99.6594
R17815 GND.n9538 GND.n541 99.6594
R17816 GND.n9540 GND.n542 99.6594
R17817 GND.n9546 GND.n543 99.6594
R17818 GND.n543 GND.n475 99.6594
R17819 GND.n9543 GND.n542 99.6594
R17820 GND.n9539 GND.n541 99.6594
R17821 GND.n9537 GND.n540 99.6594
R17822 GND.n9533 GND.n539 99.6594
R17823 GND.n9531 GND.n538 99.6594
R17824 GND.n4708 GND.n4707 81.8399
R17825 GND.n3968 GND.n3967 79.1278
R17826 GND.n3040 GND.n3039 79.1278
R17827 GND.n8284 GND.n8283 77.0988
R17828 GND.n8283 GND.n8282 77.0988
R17829 GND.n8282 GND.n1324 77.0988
R17830 GND.n8276 GND.n1324 77.0988
R17831 GND.n8276 GND.n8275 77.0988
R17832 GND.n8275 GND.n8274 77.0988
R17833 GND.n8274 GND.n1331 77.0988
R17834 GND.n8268 GND.n1331 77.0988
R17835 GND.n8268 GND.n8267 77.0988
R17836 GND.n8267 GND.n8266 77.0988
R17837 GND.n8266 GND.n1339 77.0988
R17838 GND.n8260 GND.n1339 77.0988
R17839 GND.n8260 GND.n8259 77.0988
R17840 GND.n8259 GND.n8258 77.0988
R17841 GND.n8258 GND.n1347 77.0988
R17842 GND.n8252 GND.n1347 77.0988
R17843 GND.n8252 GND.n8251 77.0988
R17844 GND.n8251 GND.n8250 77.0988
R17845 GND.n8250 GND.n1355 77.0988
R17846 GND.n8244 GND.n1355 77.0988
R17847 GND.n8244 GND.n8243 77.0988
R17848 GND.n8243 GND.n8242 77.0988
R17849 GND.n8242 GND.n1363 77.0988
R17850 GND.n8236 GND.n1363 77.0988
R17851 GND.n8236 GND.n8235 77.0988
R17852 GND.n8235 GND.n8234 77.0988
R17853 GND.n8234 GND.n1371 77.0988
R17854 GND.n8228 GND.n1371 77.0988
R17855 GND.n8228 GND.n8227 77.0988
R17856 GND.n8227 GND.n8226 77.0988
R17857 GND.n8226 GND.n1379 77.0988
R17858 GND.n8220 GND.n1379 77.0988
R17859 GND.n8220 GND.n8219 77.0988
R17860 GND.n8219 GND.n8218 77.0988
R17861 GND.n8218 GND.n1387 77.0988
R17862 GND.n8212 GND.n1387 77.0988
R17863 GND.n8212 GND.n8211 77.0988
R17864 GND.n8211 GND.n8210 77.0988
R17865 GND.n8210 GND.n1395 77.0988
R17866 GND.n8204 GND.n1395 77.0988
R17867 GND.n8204 GND.n8203 77.0988
R17868 GND.n8203 GND.n8202 77.0988
R17869 GND.n8202 GND.n1403 77.0988
R17870 GND.n8196 GND.n1403 77.0988
R17871 GND.n8196 GND.n8195 77.0988
R17872 GND.n8195 GND.n8194 77.0988
R17873 GND.n8194 GND.n1411 77.0988
R17874 GND.n8188 GND.n1411 77.0988
R17875 GND.n8188 GND.n8187 77.0988
R17876 GND.n8187 GND.n8186 77.0988
R17877 GND.n8186 GND.n1419 77.0988
R17878 GND.n8180 GND.n1419 77.0988
R17879 GND.n8180 GND.n8179 77.0988
R17880 GND.n4709 GND.n4702 72.8411
R17881 GND.n4715 GND.n4700 72.8411
R17882 GND.n6210 GND.n6209 72.8411
R17883 GND.n6252 GND.n6193 71.676
R17884 GND.n6248 GND.n6192 71.676
R17885 GND.n6244 GND.n6191 71.676
R17886 GND.n6240 GND.n6190 71.676
R17887 GND.n6236 GND.n6189 71.676
R17888 GND.n6232 GND.n6188 71.676
R17889 GND.n6228 GND.n6187 71.676
R17890 GND.n6224 GND.n6186 71.676
R17891 GND.n6219 GND.n6185 71.676
R17892 GND.n6184 GND.n6123 71.676
R17893 GND.n6183 GND.n6182 71.676
R17894 GND.n6178 GND.n6134 71.676
R17895 GND.n6174 GND.n6133 71.676
R17896 GND.n6170 GND.n6132 71.676
R17897 GND.n6166 GND.n6131 71.676
R17898 GND.n6162 GND.n6130 71.676
R17899 GND.n6158 GND.n6129 71.676
R17900 GND.n6154 GND.n6128 71.676
R17901 GND.n6150 GND.n6127 71.676
R17902 GND.n6146 GND.n6126 71.676
R17903 GND.n6142 GND.n6125 71.676
R17904 GND.n4722 GND.n4721 71.676
R17905 GND.n4728 GND.n4727 71.676
R17906 GND.n4731 GND.n4730 71.676
R17907 GND.n4736 GND.n4735 71.676
R17908 GND.n4739 GND.n4738 71.676
R17909 GND.n4744 GND.n4743 71.676
R17910 GND.n4747 GND.n4746 71.676
R17911 GND.n4752 GND.n4751 71.676
R17912 GND.n4755 GND.n4754 71.676
R17913 GND.n4761 GND.n4760 71.676
R17914 GND.n4764 GND.n4763 71.676
R17915 GND.n4769 GND.n4768 71.676
R17916 GND.n4775 GND.n4774 71.676
R17917 GND.n4778 GND.n4777 71.676
R17918 GND.n4783 GND.n4782 71.676
R17919 GND.n4786 GND.n4785 71.676
R17920 GND.n4791 GND.n4790 71.676
R17921 GND.n4794 GND.n4793 71.676
R17922 GND.n4799 GND.n4798 71.676
R17923 GND.n4802 GND.n4801 71.676
R17924 GND.n4807 GND.n4806 71.676
R17925 GND.n4723 GND.n4722 71.676
R17926 GND.n4729 GND.n4728 71.676
R17927 GND.n4730 GND.n4696 71.676
R17928 GND.n4737 GND.n4736 71.676
R17929 GND.n4738 GND.n4694 71.676
R17930 GND.n4745 GND.n4744 71.676
R17931 GND.n4746 GND.n4692 71.676
R17932 GND.n4753 GND.n4752 71.676
R17933 GND.n4754 GND.n4688 71.676
R17934 GND.n4762 GND.n4761 71.676
R17935 GND.n4767 GND.n4766 71.676
R17936 GND.n4768 GND.n4683 71.676
R17937 GND.n4776 GND.n4775 71.676
R17938 GND.n4777 GND.n4681 71.676
R17939 GND.n4784 GND.n4783 71.676
R17940 GND.n4785 GND.n4679 71.676
R17941 GND.n4792 GND.n4791 71.676
R17942 GND.n4793 GND.n4677 71.676
R17943 GND.n4800 GND.n4799 71.676
R17944 GND.n4801 GND.n4675 71.676
R17945 GND.n4808 GND.n4807 71.676
R17946 GND.n6145 GND.n6125 71.676
R17947 GND.n6149 GND.n6126 71.676
R17948 GND.n6153 GND.n6127 71.676
R17949 GND.n6157 GND.n6128 71.676
R17950 GND.n6161 GND.n6129 71.676
R17951 GND.n6165 GND.n6130 71.676
R17952 GND.n6169 GND.n6131 71.676
R17953 GND.n6173 GND.n6132 71.676
R17954 GND.n6177 GND.n6133 71.676
R17955 GND.n6181 GND.n6134 71.676
R17956 GND.n6259 GND.n6258 71.676
R17957 GND.n6218 GND.n6184 71.676
R17958 GND.n6223 GND.n6185 71.676
R17959 GND.n6227 GND.n6186 71.676
R17960 GND.n6231 GND.n6187 71.676
R17961 GND.n6235 GND.n6188 71.676
R17962 GND.n6239 GND.n6189 71.676
R17963 GND.n6243 GND.n6190 71.676
R17964 GND.n6247 GND.n6191 71.676
R17965 GND.n6251 GND.n6192 71.676
R17966 GND.n6194 GND.n6193 71.676
R17967 GND.n8178 GND.n1427 60.9094
R17968 GND.n9463 GND.n616 60.9094
R17969 GND.n63 GND.n62 60.858
R17970 GND.n65 GND.n64 60.858
R17971 GND.n106 GND.n105 60.858
R17972 GND.n108 GND.n107 60.858
R17973 GND.n20 GND.n19 60.858
R17974 GND.n22 GND.n21 60.858
R17975 GND.n297 GND.n296 60.858
R17976 GND.n295 GND.n294 60.858
R17977 GND.n340 GND.n339 60.858
R17978 GND.n338 GND.n337 60.858
R17979 GND.n384 GND.n383 60.858
R17980 GND.n382 GND.n381 60.858
R17981 GND.n4772 GND.n4685 59.5399
R17982 GND.n6137 GND.n6136 59.5399
R17983 GND.n4757 GND.n4690 59.5399
R17984 GND.n6221 GND.n6216 59.5399
R17985 GND.n4719 GND.n4718 59.1804
R17986 GND.n4706 GND.n4705 54.358
R17987 GND.n6207 GND.n6206 54.358
R17988 GND.n225 GND.n213 53.4804
R17989 GND.n6198 GND.n6197 52.4801
R17990 GND.n49 GND.t45 52.3082
R17991 GND.n72 GND.t78 52.3082
R17992 GND.n92 GND.t73 52.3082
R17993 GND.n115 GND.t61 52.3082
R17994 GND.n6 GND.t59 52.3082
R17995 GND.n29 GND.t54 52.3082
R17996 GND.n304 GND.t50 52.3082
R17997 GND.n281 GND.t76 52.3082
R17998 GND.n347 GND.t51 52.3082
R17999 GND.n324 GND.t64 52.3082
R18000 GND.n391 GND.t57 52.3082
R18001 GND.n368 GND.t74 52.3082
R18002 GND.n196 GND.t25 52.3082
R18003 GND.n184 GND.t1 52.3082
R18004 GND.n172 GND.t18 52.3082
R18005 GND.n160 GND.t5 52.3082
R18006 GND.n148 GND.t20 52.3082
R18007 GND.n137 GND.t173 52.3082
R18008 GND.n267 GND.t22 52.3082
R18009 GND.n255 GND.t15 52.3082
R18010 GND.n243 GND.t7 52.3082
R18011 GND.n231 GND.t30 52.3082
R18012 GND.n219 GND.t12 52.3082
R18013 GND.n208 GND.t28 52.3082
R18014 GND.n273 GND.n272 52.0066
R18015 GND.n261 GND.n260 52.0066
R18016 GND.n249 GND.n248 52.0066
R18017 GND.n237 GND.n236 52.0066
R18018 GND.n225 GND.n224 52.0066
R18019 GND.n6214 GND.n6213 44.3322
R18020 GND.n4709 GND.n4708 44.3189
R18021 GND.n3969 GND.n3968 42.4732
R18022 GND.n3041 GND.n3040 42.4732
R18023 GND.n9548 GND.n9545 42.2793
R18024 GND.n499 GND.n498 42.2793
R18025 GND.n9571 GND.n517 42.2793
R18026 GND.n7886 GND.n1812 42.2793
R18027 GND.n1882 GND.n1880 42.2793
R18028 GND.n2407 GND.n2378 42.2793
R18029 GND.n6321 GND.n6109 42.2793
R18030 GND.n8128 GND.n1488 42.2793
R18031 GND.n1503 GND.n1502 42.2793
R18032 GND.n3348 GND.n3347 42.2793
R18033 GND.n4707 GND.n4706 41.6274
R18034 GND.n6208 GND.n6207 41.6274
R18035 GND.n4716 GND.n4715 40.8975
R18036 GND.n6211 GND.n6210 40.8975
R18037 GND.n63 GND.n61 38.9564
R18038 GND.n106 GND.n104 38.9564
R18039 GND.n20 GND.n18 38.9564
R18040 GND.n295 GND.n293 38.9564
R18041 GND.n338 GND.n336 38.9564
R18042 GND.n382 GND.n380 38.9564
R18043 GND.n1435 GND.n1427 38.308
R18044 GND.n8169 GND.n1435 38.308
R18045 GND.n8169 GND.n8168 38.308
R18046 GND.n8168 GND.n8167 38.308
R18047 GND.n8167 GND.n1436 38.308
R18048 GND.n8161 GND.n1436 38.308
R18049 GND.n8161 GND.n8160 38.308
R18050 GND.n8160 GND.n8159 38.308
R18051 GND.n8159 GND.n1444 38.308
R18052 GND.n8153 GND.n1444 38.308
R18053 GND.n8153 GND.n8152 38.308
R18054 GND.n1509 GND.n1464 38.308
R18055 GND.n1814 GND.n1773 38.308
R18056 GND.n2954 GND.n1825 38.308
R18057 GND.n7603 GND.n2954 38.308
R18058 GND.n7603 GND.n7602 38.308
R18059 GND.n7602 GND.n7601 38.308
R18060 GND.n7302 GND.n7301 38.308
R18061 GND.n7301 GND.n7300 38.308
R18062 GND.n7300 GND.n3284 38.308
R18063 GND.n7294 GND.n3284 38.308
R18064 GND.n3356 GND.n3312 38.308
R18065 GND.n519 GND.n478 38.308
R18066 GND.n9481 GND.n544 38.308
R18067 GND.n9481 GND.n9480 38.308
R18068 GND.n9480 GND.n9479 38.308
R18069 GND.n9479 GND.n600 38.308
R18070 GND.n9473 GND.n600 38.308
R18071 GND.n9473 GND.n9472 38.308
R18072 GND.n9472 GND.n9471 38.308
R18073 GND.n9471 GND.n608 38.308
R18074 GND.n9465 GND.n608 38.308
R18075 GND.n9465 GND.n9464 38.308
R18076 GND.n9464 GND.n9463 38.308
R18077 GND.n7905 GND.n1792 36.9518
R18078 GND.n6292 GND.n6291 36.9518
R18079 GND.n85 GND.n84 36.2581
R18080 GND.n128 GND.n127 36.2581
R18081 GND.n42 GND.n41 36.2581
R18082 GND.n317 GND.n316 36.2581
R18083 GND.n360 GND.n359 36.2581
R18084 GND.n404 GND.n403 36.2581
R18085 GND.n6143 GND.n6139 35.4346
R18086 GND.n4810 GND.n4674 35.4346
R18087 GND.n4715 GND.n4714 35.055
R18088 GND.n4710 GND.n4709 35.055
R18089 GND.n6200 GND.n6199 35.055
R18090 GND.n6210 GND.n6196 35.055
R18091 GND.n7905 GND.n1795 30.6565
R18092 GND.n6292 GND.n6260 30.6565
R18093 GND.n2963 GND.n2955 29.4973
R18094 GND.n6257 GND.n6124 29.4973
R18095 GND.n4820 GND.n2981 26.0496
R18096 GND.n7574 GND.n2989 26.0496
R18097 GND.n7560 GND.n3009 26.0496
R18098 GND.n4848 GND.n3021 26.0496
R18099 GND.n4913 GND.n4646 26.0496
R18100 GND.n4920 GND.n4919 26.0496
R18101 GND.n4936 GND.n4627 26.0496
R18102 GND.n4936 GND.n4630 26.0496
R18103 GND.n4977 GND.n4598 26.0496
R18104 GND.n4970 GND.n4589 26.0496
R18105 GND.n5043 GND.n4582 26.0496
R18106 GND.n5049 GND.n4578 26.0496
R18107 GND.n5076 GND.n4559 26.0496
R18108 GND.n5101 GND.n4543 26.0496
R18109 GND.n5101 GND.n4536 26.0496
R18110 GND.n5117 GND.n4527 26.0496
R18111 GND.n5123 GND.n4510 26.0496
R18112 GND.n5128 GND.n4503 26.0496
R18113 GND.n5206 GND.n4496 26.0496
R18114 GND.n5236 GND.n4474 26.0496
R18115 GND.n5243 GND.n5242 26.0496
R18116 GND.n5259 GND.n4455 26.0496
R18117 GND.n5276 GND.n4439 26.0496
R18118 GND.n5302 GND.n4427 26.0496
R18119 GND.n5295 GND.n4417 26.0496
R18120 GND.n5368 GND.n4410 26.0496
R18121 GND.n5398 GND.n4388 26.0496
R18122 GND.n5405 GND.n5404 26.0496
R18123 GND.n5421 GND.n4369 26.0496
R18124 GND.n5421 GND.n4372 26.0496
R18125 GND.n5438 GND.n4354 26.0496
R18126 GND.n5462 GND.n4340 26.0496
R18127 GND.n5455 GND.n4331 26.0496
R18128 GND.n5538 GND.n4324 26.0496
R18129 GND.n5544 GND.n4320 26.0496
R18130 GND.n5569 GND.n4302 26.0496
R18131 GND.n5576 GND.n5575 26.0496
R18132 GND.n5592 GND.n4284 26.0496
R18133 GND.n5592 GND.n4287 26.0496
R18134 GND.n5609 GND.n4268 26.0496
R18135 GND.n5622 GND.n4256 26.0496
R18136 GND.n5645 GND.n4232 26.0496
R18137 GND.n5650 GND.n4225 26.0496
R18138 GND.n5708 GND.n4218 26.0496
R18139 GND.n5719 GND.n4213 26.0496
R18140 GND.n5794 GND.n4194 26.0496
R18141 GND.n5800 GND.n4189 26.0496
R18142 GND.n5827 GND.n4170 26.0496
R18143 GND.n5854 GND.n4155 26.0496
R18144 GND.n5860 GND.n4151 26.0496
R18145 GND.n5884 GND.n4133 26.0496
R18146 GND.n5891 GND.n5890 26.0496
R18147 GND.n5907 GND.n4114 26.0496
R18148 GND.n5907 GND.n4117 26.0496
R18149 GND.n5948 GND.n4085 26.0496
R18150 GND.n5941 GND.n4075 26.0496
R18151 GND.n6002 GND.n4068 26.0496
R18152 GND.n6008 GND.n4064 26.0496
R18153 GND.n6035 GND.n4045 26.0496
R18154 GND.n6073 GND.n4029 26.0496
R18155 GND.n6073 GND.n4020 26.0496
R18156 GND.n6066 GND.n4011 26.0496
R18157 GND.n6342 GND.n4004 26.0496
R18158 GND.n6369 GND.n3983 26.0496
R18159 GND.n6393 GND.n3230 26.0496
R18160 GND.n7328 GND.n3249 26.0496
R18161 GND.n7321 GND.n3259 26.0496
R18162 GND.n7309 GND.n3271 26.0496
R18163 GND.n5083 GND.t2 25.2835
R18164 GND.n5924 GND.t10 25.2835
R18165 GND.n7588 GND.n2971 24.5173
R18166 GND.n7580 GND.n2983 24.5173
R18167 GND.n7866 GND.n1849 24.5173
R18168 GND.n4928 GND.n4635 24.5173
R18169 GND.n4947 GND.n4946 24.5173
R18170 GND.n5089 GND.n4550 24.5173
R18171 GND.n5107 GND.n4539 24.5173
R18172 GND.n5251 GND.n4463 24.5173
R18173 GND.n5270 GND.n5269 24.5173
R18174 GND.n5413 GND.n4378 24.5173
R18175 GND.n5432 GND.n5431 24.5173
R18176 GND.n5584 GND.n4292 24.5173
R18177 GND.n5603 GND.n5602 24.5173
R18178 GND.n4212 GND.n4201 24.5173
R18179 GND.n5801 GND.n4186 24.5173
R18180 GND.n5899 GND.n4122 24.5173
R18181 GND.n5918 GND.n5917 24.5173
R18182 GND.n6048 GND.n4036 24.5173
R18183 GND.n6084 GND.n4024 24.5173
R18184 GND.n6415 GND.n6400 24.5173
R18185 GND.n6376 GND.t167 23.7512
R18186 GND.n7594 GND.t157 22.985
R18187 GND.n2992 GND.n2991 22.985
R18188 GND.n4648 GND.n4647 22.985
R18189 GND.n4562 GND.n4560 22.985
R18190 GND.n4530 GND.n4523 22.985
R18191 GND.n4476 GND.n4475 22.985
R18192 GND.n4440 GND.n4434 22.985
R18193 GND.n4390 GND.n4389 22.985
R18194 GND.n4269 GND.n4263 22.985
R18195 GND.n5707 GND.n4209 22.985
R18196 GND.n5821 GND.n5820 22.985
R18197 GND.n4135 GND.n4134 22.985
R18198 GND.n4098 GND.n4093 22.985
R18199 GND.n4014 GND.n4012 22.985
R18200 GND.n7335 GND.n7334 22.985
R18201 GND.n6140 GND.n6124 22.985
R18202 GND.n5283 GND.t4 22.6019
R18203 GND.n5615 GND.t6 22.6019
R18204 GND.t29 GND.n4349 21.8358
R18205 GND.n4304 GND.t17 21.8358
R18206 GND.n8152 GND.n8151 21.4527
R18207 GND.n7881 GND.n1825 21.4527
R18208 GND.n7566 GND.n3001 21.4527
R18209 GND.n4907 GND.n4652 21.4527
R18210 GND.n4988 GND.n4601 21.4527
R18211 GND.n5070 GND.n4566 21.4527
R18212 GND.n5152 GND.n4513 21.4527
R18213 GND.n5230 GND.n4480 21.4527
R18214 GND.n5392 GND.n4395 21.4527
R18215 GND.n5473 GND.n4344 21.4527
R18216 GND.n5563 GND.n4308 21.4527
R18217 GND.n5628 GND.n4259 21.4527
R18218 GND.n4171 GND.n4166 21.4527
R18219 GND.n5878 GND.n4139 21.4527
R18220 GND.n5959 GND.n4088 21.4527
R18221 GND.n6029 GND.n4052 21.4527
R18222 GND.n6350 GND.n3998 21.4527
R18223 GND.n7341 GND.n3232 21.4527
R18224 GND.n7294 GND.n7293 21.4527
R18225 GND.n9567 GND.n544 21.4527
R18226 GND.n4719 GND.n2968 21.3859
R18227 GND.n6214 GND.n3269 21.3859
R18228 GND.n4459 GND.t11 20.3035
R18229 GND.n4202 GND.t0 20.3035
R18230 GND.n4669 GND.n3012 19.9204
R18231 GND.n7553 GND.n3023 19.9204
R18232 GND.n4592 GND.n4590 19.9204
R18233 GND.n5042 GND.n4575 19.9204
R18234 GND.n5145 GND.n5144 19.9204
R18235 GND.n5205 GND.n4490 19.9204
R18236 GND.n5133 GND.t16 19.9204
R18237 GND.n4421 GND.n4418 19.9204
R18238 GND.n5367 GND.n4404 19.9204
R18239 GND.n4334 GND.n4332 19.9204
R18240 GND.n5537 GND.n4317 19.9204
R18241 GND.n4250 GND.n4244 19.9204
R18242 GND.n5686 GND.n5684 19.9204
R18243 GND.n5835 GND.t13 19.9204
R18244 GND.n5841 GND.n4162 19.9204
R18245 GND.n5853 GND.n5852 19.9204
R18246 GND.n4079 GND.n4076 19.9204
R18247 GND.n6001 GND.n4061 19.9204
R18248 GND.n6362 GND.n6361 19.9204
R18249 GND.n3985 GND.n3984 19.9204
R18250 GND.n4703 GND.t119 19.8005
R18251 GND.n4703 GND.t82 19.8005
R18252 GND.n4704 GND.t158 19.8005
R18253 GND.n4704 GND.t99 19.8005
R18254 GND.n6204 GND.t171 19.8005
R18255 GND.n6204 GND.t89 19.8005
R18256 GND.n6205 GND.t168 19.8005
R18257 GND.n6205 GND.t155 19.8005
R18258 GND.n4700 GND.n4699 19.5087
R18259 GND.n4713 GND.n4700 19.5087
R18260 GND.n4711 GND.n4702 19.5087
R18261 GND.n6209 GND.n6203 19.5087
R18262 GND.n9565 GND.n546 19.3944
R18263 GND.n9561 GND.n546 19.3944
R18264 GND.n9561 GND.n9560 19.3944
R18265 GND.n9560 GND.n9559 19.3944
R18266 GND.n9559 GND.n9535 19.3944
R18267 GND.n9555 GND.n9535 19.3944
R18268 GND.n9555 GND.n9554 19.3944
R18269 GND.n9554 GND.n9553 19.3944
R18270 GND.n9553 GND.n9541 19.3944
R18271 GND.n9549 GND.n9541 19.3944
R18272 GND.n6324 GND.n3372 19.3944
R18273 GND.n7248 GND.n3372 19.3944
R18274 GND.n7248 GND.n3373 19.3944
R18275 GND.n3382 GND.n3373 19.3944
R18276 GND.n3383 GND.n3382 19.3944
R18277 GND.n3384 GND.n3383 19.3944
R18278 GND.n3951 GND.n3384 19.3944
R18279 GND.n3951 GND.n3390 19.3944
R18280 GND.n3391 GND.n3390 19.3944
R18281 GND.n3392 GND.n3391 19.3944
R18282 GND.n3928 GND.n3392 19.3944
R18283 GND.n3928 GND.n3398 19.3944
R18284 GND.n3399 GND.n3398 19.3944
R18285 GND.n3400 GND.n3399 19.3944
R18286 GND.n3915 GND.n3400 19.3944
R18287 GND.n3915 GND.n3406 19.3944
R18288 GND.n3407 GND.n3406 19.3944
R18289 GND.n3408 GND.n3407 19.3944
R18290 GND.n6654 GND.n3408 19.3944
R18291 GND.n6654 GND.n3414 19.3944
R18292 GND.n3415 GND.n3414 19.3944
R18293 GND.n3416 GND.n3415 19.3944
R18294 GND.n6681 GND.n3416 19.3944
R18295 GND.n6681 GND.n3422 19.3944
R18296 GND.n3423 GND.n3422 19.3944
R18297 GND.n3424 GND.n3423 19.3944
R18298 GND.n3860 GND.n3424 19.3944
R18299 GND.n3860 GND.n3430 19.3944
R18300 GND.n3431 GND.n3430 19.3944
R18301 GND.n3432 GND.n3431 19.3944
R18302 GND.n3837 GND.n3432 19.3944
R18303 GND.n3837 GND.n3438 19.3944
R18304 GND.n3439 GND.n3438 19.3944
R18305 GND.n3440 GND.n3439 19.3944
R18306 GND.n3824 GND.n3440 19.3944
R18307 GND.n3824 GND.n3446 19.3944
R18308 GND.n3447 GND.n3446 19.3944
R18309 GND.n3448 GND.n3447 19.3944
R18310 GND.n6753 GND.n3448 19.3944
R18311 GND.n6753 GND.n3454 19.3944
R18312 GND.n3455 GND.n3454 19.3944
R18313 GND.n3456 GND.n3455 19.3944
R18314 GND.n6780 GND.n3456 19.3944
R18315 GND.n6780 GND.n3462 19.3944
R18316 GND.n3463 GND.n3462 19.3944
R18317 GND.n3464 GND.n3463 19.3944
R18318 GND.n3779 GND.n3464 19.3944
R18319 GND.n3779 GND.n3470 19.3944
R18320 GND.n3471 GND.n3470 19.3944
R18321 GND.n3472 GND.n3471 19.3944
R18322 GND.n3764 GND.n3472 19.3944
R18323 GND.n3764 GND.n3478 19.3944
R18324 GND.n3479 GND.n3478 19.3944
R18325 GND.n3480 GND.n3479 19.3944
R18326 GND.n6851 GND.n3480 19.3944
R18327 GND.n6851 GND.n3486 19.3944
R18328 GND.n3487 GND.n3486 19.3944
R18329 GND.n3488 GND.n3487 19.3944
R18330 GND.n3734 GND.n3488 19.3944
R18331 GND.n3734 GND.n3494 19.3944
R18332 GND.n3495 GND.n3494 19.3944
R18333 GND.n3496 GND.n3495 19.3944
R18334 GND.n3711 GND.n3496 19.3944
R18335 GND.n3711 GND.n3502 19.3944
R18336 GND.n3503 GND.n3502 19.3944
R18337 GND.n3504 GND.n3503 19.3944
R18338 GND.n3700 GND.n3504 19.3944
R18339 GND.n3700 GND.n3510 19.3944
R18340 GND.n3511 GND.n3510 19.3944
R18341 GND.n3512 GND.n3511 19.3944
R18342 GND.n6944 GND.n3512 19.3944
R18343 GND.n6944 GND.n3518 19.3944
R18344 GND.n3519 GND.n3518 19.3944
R18345 GND.n3520 GND.n3519 19.3944
R18346 GND.n6973 GND.n3520 19.3944
R18347 GND.n6973 GND.n3526 19.3944
R18348 GND.n3527 GND.n3526 19.3944
R18349 GND.n3528 GND.n3527 19.3944
R18350 GND.n3648 GND.n3528 19.3944
R18351 GND.n3648 GND.n3534 19.3944
R18352 GND.n3535 GND.n3534 19.3944
R18353 GND.n3536 GND.n3535 19.3944
R18354 GND.n3625 GND.n3536 19.3944
R18355 GND.n3625 GND.n3542 19.3944
R18356 GND.n3543 GND.n3542 19.3944
R18357 GND.n3544 GND.n3543 19.3944
R18358 GND.n3614 GND.n3544 19.3944
R18359 GND.n3614 GND.n3550 19.3944
R18360 GND.n3551 GND.n3550 19.3944
R18361 GND.n3552 GND.n3551 19.3944
R18362 GND.n7053 GND.n3552 19.3944
R18363 GND.n7053 GND.n3558 19.3944
R18364 GND.n3559 GND.n3558 19.3944
R18365 GND.n3560 GND.n3559 19.3944
R18366 GND.n7087 GND.n3560 19.3944
R18367 GND.n7087 GND.n3566 19.3944
R18368 GND.n3567 GND.n3566 19.3944
R18369 GND.n7102 GND.n3567 19.3944
R18370 GND.n7102 GND.n574 19.3944
R18371 GND.n9504 GND.n574 19.3944
R18372 GND.n9504 GND.n575 19.3944
R18373 GND.n575 GND.n553 19.3944
R18374 GND.n9521 GND.n553 19.3944
R18375 GND.n9522 GND.n9521 19.3944
R18376 GND.n9522 GND.n548 19.3944
R18377 GND.n6325 GND.n3378 19.3944
R18378 GND.n7246 GND.n3378 19.3944
R18379 GND.n7246 GND.n7245 19.3944
R18380 GND.n7245 GND.n7244 19.3944
R18381 GND.n7244 GND.n3381 19.3944
R18382 GND.n7240 GND.n3381 19.3944
R18383 GND.n7240 GND.n7239 19.3944
R18384 GND.n7239 GND.n7238 19.3944
R18385 GND.n7238 GND.n3389 19.3944
R18386 GND.n7234 GND.n3389 19.3944
R18387 GND.n7234 GND.n7233 19.3944
R18388 GND.n7233 GND.n7232 19.3944
R18389 GND.n7232 GND.n3397 19.3944
R18390 GND.n7228 GND.n3397 19.3944
R18391 GND.n7228 GND.n7227 19.3944
R18392 GND.n7227 GND.n7226 19.3944
R18393 GND.n7226 GND.n3405 19.3944
R18394 GND.n7222 GND.n3405 19.3944
R18395 GND.n7222 GND.n7221 19.3944
R18396 GND.n7221 GND.n7220 19.3944
R18397 GND.n7220 GND.n3413 19.3944
R18398 GND.n7216 GND.n3413 19.3944
R18399 GND.n7216 GND.n7215 19.3944
R18400 GND.n7215 GND.n7214 19.3944
R18401 GND.n7214 GND.n3421 19.3944
R18402 GND.n7210 GND.n3421 19.3944
R18403 GND.n7210 GND.n7209 19.3944
R18404 GND.n7209 GND.n7208 19.3944
R18405 GND.n7208 GND.n3429 19.3944
R18406 GND.n7204 GND.n3429 19.3944
R18407 GND.n7204 GND.n7203 19.3944
R18408 GND.n7203 GND.n7202 19.3944
R18409 GND.n7202 GND.n3437 19.3944
R18410 GND.n7198 GND.n3437 19.3944
R18411 GND.n7198 GND.n7197 19.3944
R18412 GND.n7197 GND.n7196 19.3944
R18413 GND.n7196 GND.n3445 19.3944
R18414 GND.n7192 GND.n3445 19.3944
R18415 GND.n7192 GND.n7191 19.3944
R18416 GND.n7191 GND.n7190 19.3944
R18417 GND.n7190 GND.n3453 19.3944
R18418 GND.n7186 GND.n3453 19.3944
R18419 GND.n7186 GND.n7185 19.3944
R18420 GND.n7185 GND.n7184 19.3944
R18421 GND.n7184 GND.n3461 19.3944
R18422 GND.n7180 GND.n3461 19.3944
R18423 GND.n7180 GND.n7179 19.3944
R18424 GND.n7179 GND.n7178 19.3944
R18425 GND.n7178 GND.n3469 19.3944
R18426 GND.n7174 GND.n3469 19.3944
R18427 GND.n7174 GND.n7173 19.3944
R18428 GND.n7173 GND.n7172 19.3944
R18429 GND.n7172 GND.n3477 19.3944
R18430 GND.n7168 GND.n3477 19.3944
R18431 GND.n7168 GND.n7167 19.3944
R18432 GND.n7167 GND.n7166 19.3944
R18433 GND.n7166 GND.n3485 19.3944
R18434 GND.n7162 GND.n3485 19.3944
R18435 GND.n7162 GND.n7161 19.3944
R18436 GND.n7161 GND.n7160 19.3944
R18437 GND.n7160 GND.n3493 19.3944
R18438 GND.n7156 GND.n3493 19.3944
R18439 GND.n7156 GND.n7155 19.3944
R18440 GND.n7155 GND.n7154 19.3944
R18441 GND.n7154 GND.n3501 19.3944
R18442 GND.n7150 GND.n3501 19.3944
R18443 GND.n7150 GND.n7149 19.3944
R18444 GND.n7149 GND.n7148 19.3944
R18445 GND.n7148 GND.n3509 19.3944
R18446 GND.n7144 GND.n3509 19.3944
R18447 GND.n7144 GND.n7143 19.3944
R18448 GND.n7143 GND.n7142 19.3944
R18449 GND.n7142 GND.n3517 19.3944
R18450 GND.n7138 GND.n3517 19.3944
R18451 GND.n7138 GND.n7137 19.3944
R18452 GND.n7137 GND.n7136 19.3944
R18453 GND.n7136 GND.n3525 19.3944
R18454 GND.n7132 GND.n3525 19.3944
R18455 GND.n7132 GND.n7131 19.3944
R18456 GND.n7131 GND.n7130 19.3944
R18457 GND.n7130 GND.n3533 19.3944
R18458 GND.n7126 GND.n3533 19.3944
R18459 GND.n7126 GND.n7125 19.3944
R18460 GND.n7125 GND.n7124 19.3944
R18461 GND.n7124 GND.n3541 19.3944
R18462 GND.n7120 GND.n3541 19.3944
R18463 GND.n7120 GND.n7119 19.3944
R18464 GND.n7119 GND.n7118 19.3944
R18465 GND.n7118 GND.n3549 19.3944
R18466 GND.n7114 GND.n3549 19.3944
R18467 GND.n7114 GND.n7113 19.3944
R18468 GND.n7113 GND.n7112 19.3944
R18469 GND.n7112 GND.n3557 19.3944
R18470 GND.n7108 GND.n3557 19.3944
R18471 GND.n7108 GND.n7107 19.3944
R18472 GND.n7107 GND.n7106 19.3944
R18473 GND.n7106 GND.n3565 19.3944
R18474 GND.n3565 GND.n577 19.3944
R18475 GND.n9501 GND.n577 19.3944
R18476 GND.n9502 GND.n9501 19.3944
R18477 GND.n9502 GND.n555 19.3944
R18478 GND.n9518 GND.n555 19.3944
R18479 GND.n9518 GND.n549 19.3944
R18480 GND.n9526 GND.n549 19.3944
R18481 GND.n9527 GND.n9526 19.3944
R18482 GND.n9607 GND.n9606 19.3944
R18483 GND.n9606 GND.n9605 19.3944
R18484 GND.n9605 GND.n487 19.3944
R18485 GND.n9601 GND.n487 19.3944
R18486 GND.n9601 GND.n9600 19.3944
R18487 GND.n9600 GND.n9599 19.3944
R18488 GND.n9599 GND.n492 19.3944
R18489 GND.n9595 GND.n492 19.3944
R18490 GND.n9595 GND.n9594 19.3944
R18491 GND.n9594 GND.n9593 19.3944
R18492 GND.n9589 GND.n9588 19.3944
R18493 GND.n9588 GND.n9587 19.3944
R18494 GND.n9587 GND.n504 19.3944
R18495 GND.n9583 GND.n504 19.3944
R18496 GND.n9583 GND.n9582 19.3944
R18497 GND.n9582 GND.n9581 19.3944
R18498 GND.n9581 GND.n509 19.3944
R18499 GND.n9577 GND.n509 19.3944
R18500 GND.n9577 GND.n9576 19.3944
R18501 GND.n9576 GND.n9575 19.3944
R18502 GND.n9575 GND.n514 19.3944
R18503 GND.n1561 GND.n1558 19.3944
R18504 GND.n1561 GND.n1556 19.3944
R18505 GND.n1568 GND.n1556 19.3944
R18506 GND.n1569 GND.n1568 19.3944
R18507 GND.n8076 GND.n1569 19.3944
R18508 GND.n8076 GND.n8075 19.3944
R18509 GND.n8075 GND.n8074 19.3944
R18510 GND.n8074 GND.n1572 19.3944
R18511 GND.n8070 GND.n1572 19.3944
R18512 GND.n8070 GND.n8069 19.3944
R18513 GND.n8069 GND.n8068 19.3944
R18514 GND.n8068 GND.n1580 19.3944
R18515 GND.n8064 GND.n1580 19.3944
R18516 GND.n8064 GND.n8063 19.3944
R18517 GND.n8063 GND.n8062 19.3944
R18518 GND.n8062 GND.n1588 19.3944
R18519 GND.n8058 GND.n1588 19.3944
R18520 GND.n8058 GND.n8057 19.3944
R18521 GND.n8057 GND.n8056 19.3944
R18522 GND.n8056 GND.n1596 19.3944
R18523 GND.n8052 GND.n1596 19.3944
R18524 GND.n8052 GND.n8051 19.3944
R18525 GND.n8051 GND.n8050 19.3944
R18526 GND.n8050 GND.n1604 19.3944
R18527 GND.n8046 GND.n1604 19.3944
R18528 GND.n8046 GND.n8045 19.3944
R18529 GND.n8045 GND.n8044 19.3944
R18530 GND.n8044 GND.n1612 19.3944
R18531 GND.n8040 GND.n1612 19.3944
R18532 GND.n8040 GND.n8039 19.3944
R18533 GND.n8039 GND.n8038 19.3944
R18534 GND.n8038 GND.n1620 19.3944
R18535 GND.n8034 GND.n1620 19.3944
R18536 GND.n8034 GND.n8033 19.3944
R18537 GND.n8033 GND.n8032 19.3944
R18538 GND.n8032 GND.n1628 19.3944
R18539 GND.n8028 GND.n1628 19.3944
R18540 GND.n8028 GND.n8027 19.3944
R18541 GND.n8027 GND.n8026 19.3944
R18542 GND.n8026 GND.n1636 19.3944
R18543 GND.n8022 GND.n1636 19.3944
R18544 GND.n8022 GND.n8021 19.3944
R18545 GND.n8021 GND.n8020 19.3944
R18546 GND.n8020 GND.n1644 19.3944
R18547 GND.n8016 GND.n1644 19.3944
R18548 GND.n8016 GND.n8015 19.3944
R18549 GND.n8015 GND.n8014 19.3944
R18550 GND.n8014 GND.n1652 19.3944
R18551 GND.n8010 GND.n1652 19.3944
R18552 GND.n8010 GND.n8009 19.3944
R18553 GND.n8009 GND.n8008 19.3944
R18554 GND.n8008 GND.n1660 19.3944
R18555 GND.n8004 GND.n1660 19.3944
R18556 GND.n8004 GND.n8003 19.3944
R18557 GND.n8003 GND.n8002 19.3944
R18558 GND.n8002 GND.n1668 19.3944
R18559 GND.n7998 GND.n1668 19.3944
R18560 GND.n7998 GND.n7997 19.3944
R18561 GND.n7997 GND.n7996 19.3944
R18562 GND.n7996 GND.n1676 19.3944
R18563 GND.n7992 GND.n1676 19.3944
R18564 GND.n7992 GND.n7991 19.3944
R18565 GND.n7991 GND.n7990 19.3944
R18566 GND.n7990 GND.n1684 19.3944
R18567 GND.n7986 GND.n1684 19.3944
R18568 GND.n7986 GND.n7985 19.3944
R18569 GND.n7985 GND.n7984 19.3944
R18570 GND.n7984 GND.n1692 19.3944
R18571 GND.n7980 GND.n1692 19.3944
R18572 GND.n7980 GND.n7979 19.3944
R18573 GND.n7979 GND.n7978 19.3944
R18574 GND.n7978 GND.n1700 19.3944
R18575 GND.n7974 GND.n1700 19.3944
R18576 GND.n7974 GND.n7973 19.3944
R18577 GND.n7973 GND.n7972 19.3944
R18578 GND.n7972 GND.n1708 19.3944
R18579 GND.n7968 GND.n1708 19.3944
R18580 GND.n7968 GND.n7967 19.3944
R18581 GND.n7967 GND.n7966 19.3944
R18582 GND.n7966 GND.n1716 19.3944
R18583 GND.n7962 GND.n1716 19.3944
R18584 GND.n7962 GND.n7961 19.3944
R18585 GND.n7961 GND.n7960 19.3944
R18586 GND.n7960 GND.n1724 19.3944
R18587 GND.n7956 GND.n1724 19.3944
R18588 GND.n7956 GND.n7955 19.3944
R18589 GND.n7955 GND.n7954 19.3944
R18590 GND.n7954 GND.n1732 19.3944
R18591 GND.n7950 GND.n1732 19.3944
R18592 GND.n7950 GND.n7949 19.3944
R18593 GND.n7949 GND.n7948 19.3944
R18594 GND.n7948 GND.n1740 19.3944
R18595 GND.n7944 GND.n1740 19.3944
R18596 GND.n7944 GND.n7943 19.3944
R18597 GND.n7943 GND.n7942 19.3944
R18598 GND.n7942 GND.n1748 19.3944
R18599 GND.n7938 GND.n1748 19.3944
R18600 GND.n7938 GND.n7937 19.3944
R18601 GND.n7937 GND.n7936 19.3944
R18602 GND.n7936 GND.n1756 19.3944
R18603 GND.n7932 GND.n1756 19.3944
R18604 GND.n7932 GND.n7931 19.3944
R18605 GND.n7931 GND.n7930 19.3944
R18606 GND.n7930 GND.n1764 19.3944
R18607 GND.n7926 GND.n1764 19.3944
R18608 GND.n7919 GND.n7918 19.3944
R18609 GND.n7918 GND.n7917 19.3944
R18610 GND.n7917 GND.n1782 19.3944
R18611 GND.n7913 GND.n1782 19.3944
R18612 GND.n7913 GND.n7912 19.3944
R18613 GND.n7912 GND.n7911 19.3944
R18614 GND.n7911 GND.n1787 19.3944
R18615 GND.n7907 GND.n1787 19.3944
R18616 GND.n7907 GND.n7906 19.3944
R18617 GND.n7904 GND.n1797 19.3944
R18618 GND.n7900 GND.n1797 19.3944
R18619 GND.n7900 GND.n7899 19.3944
R18620 GND.n7899 GND.n7898 19.3944
R18621 GND.n7898 GND.n1802 19.3944
R18622 GND.n7894 GND.n1802 19.3944
R18623 GND.n7894 GND.n7893 19.3944
R18624 GND.n7893 GND.n7892 19.3944
R18625 GND.n7892 GND.n1807 19.3944
R18626 GND.n7888 GND.n1807 19.3944
R18627 GND.n7888 GND.n7887 19.3944
R18628 GND.n2412 GND.n2374 19.3944
R18629 GND.n2415 GND.n2412 19.3944
R18630 GND.n2416 GND.n2415 19.3944
R18631 GND.n2416 GND.n2372 19.3944
R18632 GND.n2420 GND.n2372 19.3944
R18633 GND.n2421 GND.n2420 19.3944
R18634 GND.n2516 GND.n2421 19.3944
R18635 GND.n2516 GND.n2366 19.3944
R18636 GND.n2521 GND.n2366 19.3944
R18637 GND.n2521 GND.n2367 19.3944
R18638 GND.n2367 GND.n2347 19.3944
R18639 GND.n2541 GND.n2347 19.3944
R18640 GND.n2541 GND.n2344 19.3944
R18641 GND.n2546 GND.n2344 19.3944
R18642 GND.n2546 GND.n2345 19.3944
R18643 GND.n2345 GND.n2325 19.3944
R18644 GND.n2566 GND.n2325 19.3944
R18645 GND.n2566 GND.n2322 19.3944
R18646 GND.n2571 GND.n2322 19.3944
R18647 GND.n2571 GND.n2323 19.3944
R18648 GND.n2323 GND.n2301 19.3944
R18649 GND.n2590 GND.n2301 19.3944
R18650 GND.n2590 GND.n2298 19.3944
R18651 GND.n2595 GND.n2298 19.3944
R18652 GND.n2595 GND.n2299 19.3944
R18653 GND.n2299 GND.n2278 19.3944
R18654 GND.n2615 GND.n2278 19.3944
R18655 GND.n2615 GND.n2275 19.3944
R18656 GND.n2629 GND.n2275 19.3944
R18657 GND.n2629 GND.n2276 19.3944
R18658 GND.n2625 GND.n2276 19.3944
R18659 GND.n2625 GND.n2624 19.3944
R18660 GND.n2624 GND.n2623 19.3944
R18661 GND.n2623 GND.n2620 19.3944
R18662 GND.n2620 GND.n2237 19.3944
R18663 GND.n2715 GND.n2237 19.3944
R18664 GND.n2715 GND.n2234 19.3944
R18665 GND.n2720 GND.n2234 19.3944
R18666 GND.n2720 GND.n2235 19.3944
R18667 GND.n2235 GND.n2215 19.3944
R18668 GND.n2740 GND.n2215 19.3944
R18669 GND.n2740 GND.n2212 19.3944
R18670 GND.n2745 GND.n2212 19.3944
R18671 GND.n2745 GND.n2213 19.3944
R18672 GND.n2213 GND.n2193 19.3944
R18673 GND.n2762 GND.n2193 19.3944
R18674 GND.n2762 GND.n2191 19.3944
R18675 GND.n2766 GND.n2191 19.3944
R18676 GND.n2767 GND.n2766 19.3944
R18677 GND.n2770 GND.n2767 19.3944
R18678 GND.n2770 GND.n2189 19.3944
R18679 GND.n2775 GND.n2189 19.3944
R18680 GND.n2776 GND.n2775 19.3944
R18681 GND.n2777 GND.n2776 19.3944
R18682 GND.n2777 GND.n2187 19.3944
R18683 GND.n2781 GND.n2187 19.3944
R18684 GND.n2781 GND.n2096 19.3944
R18685 GND.n2832 GND.n2096 19.3944
R18686 GND.n2832 GND.n2093 19.3944
R18687 GND.n2837 GND.n2093 19.3944
R18688 GND.n2837 GND.n2094 19.3944
R18689 GND.n2094 GND.n2073 19.3944
R18690 GND.n2857 GND.n2073 19.3944
R18691 GND.n2857 GND.n2070 19.3944
R18692 GND.n2862 GND.n2070 19.3944
R18693 GND.n2862 GND.n2071 19.3944
R18694 GND.n2071 GND.n2051 19.3944
R18695 GND.n2882 GND.n2051 19.3944
R18696 GND.n2882 GND.n2048 19.3944
R18697 GND.n2887 GND.n2048 19.3944
R18698 GND.n2887 GND.n2049 19.3944
R18699 GND.n2049 GND.n2024 19.3944
R18700 GND.n7680 GND.n2024 19.3944
R18701 GND.n7680 GND.n2021 19.3944
R18702 GND.n7685 GND.n2021 19.3944
R18703 GND.n7685 GND.n2022 19.3944
R18704 GND.n2022 GND.n2000 19.3944
R18705 GND.n7704 GND.n2000 19.3944
R18706 GND.n7704 GND.n1997 19.3944
R18707 GND.n7709 GND.n1997 19.3944
R18708 GND.n7709 GND.n1998 19.3944
R18709 GND.n1998 GND.n1977 19.3944
R18710 GND.n7729 GND.n1977 19.3944
R18711 GND.n7729 GND.n1974 19.3944
R18712 GND.n7734 GND.n1974 19.3944
R18713 GND.n7734 GND.n1975 19.3944
R18714 GND.n1975 GND.n1955 19.3944
R18715 GND.n7754 GND.n1955 19.3944
R18716 GND.n7754 GND.n1952 19.3944
R18717 GND.n7759 GND.n1952 19.3944
R18718 GND.n7759 GND.n1953 19.3944
R18719 GND.n1953 GND.n1933 19.3944
R18720 GND.n7779 GND.n1933 19.3944
R18721 GND.n7779 GND.n1930 19.3944
R18722 GND.n7784 GND.n1930 19.3944
R18723 GND.n7784 GND.n1931 19.3944
R18724 GND.n1931 GND.n1910 19.3944
R18725 GND.n7803 GND.n1910 19.3944
R18726 GND.n7803 GND.n1907 19.3944
R18727 GND.n7813 GND.n1907 19.3944
R18728 GND.n7813 GND.n1908 19.3944
R18729 GND.n7809 GND.n1908 19.3944
R18730 GND.n7809 GND.n1889 19.3944
R18731 GND.n7831 GND.n1889 19.3944
R18732 GND.n7832 GND.n7831 19.3944
R18733 GND.n7872 GND.n1833 19.3944
R18734 GND.n1855 GND.n1833 19.3944
R18735 GND.n7861 GND.n1855 19.3944
R18736 GND.n7861 GND.n7860 19.3944
R18737 GND.n7860 GND.n1860 19.3944
R18738 GND.n7853 GND.n1860 19.3944
R18739 GND.n7853 GND.n7852 19.3944
R18740 GND.n7852 GND.n1868 19.3944
R18741 GND.n7845 GND.n1868 19.3944
R18742 GND.n7845 GND.n7844 19.3944
R18743 GND.n8097 GND.n1506 19.3944
R18744 GND.n2390 GND.n1506 19.3944
R18745 GND.n2391 GND.n2390 19.3944
R18746 GND.n2394 GND.n2391 19.3944
R18747 GND.n2394 GND.n2383 19.3944
R18748 GND.n2398 GND.n2383 19.3944
R18749 GND.n2399 GND.n2398 19.3944
R18750 GND.n2402 GND.n2399 19.3944
R18751 GND.n2402 GND.n2379 19.3944
R18752 GND.n2406 GND.n2379 19.3944
R18753 GND.n1563 GND.n1508 19.3944
R18754 GND.n1565 GND.n1563 19.3944
R18755 GND.n1566 GND.n1565 19.3944
R18756 GND.n1566 GND.n1552 19.3944
R18757 GND.n8078 GND.n1552 19.3944
R18758 GND.n8078 GND.n1553 19.3944
R18759 GND.n1573 GND.n1553 19.3944
R18760 GND.n1574 GND.n1573 19.3944
R18761 GND.n1575 GND.n1574 19.3944
R18762 GND.n2527 GND.n1575 19.3944
R18763 GND.n2527 GND.n1581 19.3944
R18764 GND.n1582 GND.n1581 19.3944
R18765 GND.n1583 GND.n1582 19.3944
R18766 GND.n2341 GND.n1583 19.3944
R18767 GND.n2341 GND.n1589 19.3944
R18768 GND.n1590 GND.n1589 19.3944
R18769 GND.n1591 GND.n1590 19.3944
R18770 GND.n2318 GND.n1591 19.3944
R18771 GND.n2318 GND.n1597 19.3944
R18772 GND.n1598 GND.n1597 19.3944
R18773 GND.n1599 GND.n1598 19.3944
R18774 GND.n2305 GND.n1599 19.3944
R18775 GND.n2305 GND.n1605 19.3944
R18776 GND.n1606 GND.n1605 19.3944
R18777 GND.n1607 GND.n1606 19.3944
R18778 GND.n2599 GND.n1607 19.3944
R18779 GND.n2599 GND.n1613 19.3944
R18780 GND.n1614 GND.n1613 19.3944
R18781 GND.n1615 GND.n1614 19.3944
R18782 GND.n2634 GND.n1615 19.3944
R18783 GND.n2634 GND.n1621 19.3944
R18784 GND.n1622 GND.n1621 19.3944
R18785 GND.n1623 GND.n1622 19.3944
R18786 GND.n2701 GND.n1623 19.3944
R18787 GND.n2701 GND.n1629 19.3944
R18788 GND.n1630 GND.n1629 19.3944
R18789 GND.n1631 GND.n1630 19.3944
R18790 GND.n2231 GND.n1631 19.3944
R18791 GND.n2231 GND.n1637 19.3944
R18792 GND.n1638 GND.n1637 19.3944
R18793 GND.n1639 GND.n1638 19.3944
R18794 GND.n2208 GND.n1639 19.3944
R18795 GND.n2208 GND.n1645 19.3944
R18796 GND.n1646 GND.n1645 19.3944
R18797 GND.n1647 GND.n1646 19.3944
R18798 GND.n2197 GND.n1647 19.3944
R18799 GND.n2197 GND.n1653 19.3944
R18800 GND.n1654 GND.n1653 19.3944
R18801 GND.n1655 GND.n1654 19.3944
R18802 GND.n2121 GND.n1655 19.3944
R18803 GND.n2121 GND.n1661 19.3944
R18804 GND.n1662 GND.n1661 19.3944
R18805 GND.n1663 GND.n1662 19.3944
R18806 GND.n2144 GND.n1663 19.3944
R18807 GND.n2144 GND.n1669 19.3944
R18808 GND.n1670 GND.n1669 19.3944
R18809 GND.n1671 GND.n1670 19.3944
R18810 GND.n2100 GND.n1671 19.3944
R18811 GND.n2100 GND.n1677 19.3944
R18812 GND.n1678 GND.n1677 19.3944
R18813 GND.n1679 GND.n1678 19.3944
R18814 GND.n2841 GND.n1679 19.3944
R18815 GND.n2841 GND.n1685 19.3944
R18816 GND.n1686 GND.n1685 19.3944
R18817 GND.n1687 GND.n1686 19.3944
R18818 GND.n2868 GND.n1687 19.3944
R18819 GND.n2868 GND.n1693 19.3944
R18820 GND.n1694 GND.n1693 19.3944
R18821 GND.n1695 GND.n1694 19.3944
R18822 GND.n2038 GND.n1695 19.3944
R18823 GND.n2038 GND.n1701 19.3944
R18824 GND.n1702 GND.n1701 19.3944
R18825 GND.n1703 GND.n1702 19.3944
R18826 GND.n2017 GND.n1703 19.3944
R18827 GND.n2017 GND.n1709 19.3944
R18828 GND.n1710 GND.n1709 19.3944
R18829 GND.n1711 GND.n1710 19.3944
R18830 GND.n2004 GND.n1711 19.3944
R18831 GND.n2004 GND.n1717 19.3944
R18832 GND.n1718 GND.n1717 19.3944
R18833 GND.n1719 GND.n1718 19.3944
R18834 GND.n7713 GND.n1719 19.3944
R18835 GND.n7713 GND.n1725 19.3944
R18836 GND.n1726 GND.n1725 19.3944
R18837 GND.n1727 GND.n1726 19.3944
R18838 GND.n7740 GND.n1727 19.3944
R18839 GND.n7740 GND.n1733 19.3944
R18840 GND.n1734 GND.n1733 19.3944
R18841 GND.n1735 GND.n1734 19.3944
R18842 GND.n1949 GND.n1735 19.3944
R18843 GND.n1949 GND.n1741 19.3944
R18844 GND.n1742 GND.n1741 19.3944
R18845 GND.n1743 GND.n1742 19.3944
R18846 GND.n1926 GND.n1743 19.3944
R18847 GND.n1926 GND.n1749 19.3944
R18848 GND.n1750 GND.n1749 19.3944
R18849 GND.n1751 GND.n1750 19.3944
R18850 GND.n1913 GND.n1751 19.3944
R18851 GND.n1913 GND.n1757 19.3944
R18852 GND.n1758 GND.n1757 19.3944
R18853 GND.n1759 GND.n1758 19.3944
R18854 GND.n1892 GND.n1759 19.3944
R18855 GND.n1892 GND.n1765 19.3944
R18856 GND.n1766 GND.n1765 19.3944
R18857 GND.n1767 GND.n1766 19.3944
R18858 GND.n3054 GND.n3053 19.3944
R18859 GND.n3054 GND.n3026 19.3944
R18860 GND.n7551 GND.n3026 19.3944
R18861 GND.n7551 GND.n3027 19.3944
R18862 GND.n7547 GND.n3027 19.3944
R18863 GND.n7547 GND.n7546 19.3944
R18864 GND.n7546 GND.n7545 19.3944
R18865 GND.n7545 GND.n3061 19.3944
R18866 GND.n7541 GND.n3061 19.3944
R18867 GND.n7541 GND.n7540 19.3944
R18868 GND.n7540 GND.n7539 19.3944
R18869 GND.n7539 GND.n3066 19.3944
R18870 GND.n7535 GND.n3066 19.3944
R18871 GND.n7535 GND.n7534 19.3944
R18872 GND.n7534 GND.n7533 19.3944
R18873 GND.n7533 GND.n3071 19.3944
R18874 GND.n7529 GND.n3071 19.3944
R18875 GND.n7529 GND.n7528 19.3944
R18876 GND.n7528 GND.n7527 19.3944
R18877 GND.n7527 GND.n3076 19.3944
R18878 GND.n7523 GND.n3076 19.3944
R18879 GND.n7523 GND.n7522 19.3944
R18880 GND.n7522 GND.n7521 19.3944
R18881 GND.n7521 GND.n3081 19.3944
R18882 GND.n7517 GND.n3081 19.3944
R18883 GND.n7517 GND.n7516 19.3944
R18884 GND.n7516 GND.n7515 19.3944
R18885 GND.n7515 GND.n3086 19.3944
R18886 GND.n7511 GND.n3086 19.3944
R18887 GND.n7511 GND.n7510 19.3944
R18888 GND.n7510 GND.n7509 19.3944
R18889 GND.n7509 GND.n3091 19.3944
R18890 GND.n7505 GND.n3091 19.3944
R18891 GND.n7505 GND.n7504 19.3944
R18892 GND.n7504 GND.n7503 19.3944
R18893 GND.n7503 GND.n3096 19.3944
R18894 GND.n7499 GND.n3096 19.3944
R18895 GND.n7499 GND.n7498 19.3944
R18896 GND.n7498 GND.n7497 19.3944
R18897 GND.n7497 GND.n3101 19.3944
R18898 GND.n7493 GND.n3101 19.3944
R18899 GND.n7493 GND.n7492 19.3944
R18900 GND.n7492 GND.n7491 19.3944
R18901 GND.n7491 GND.n3106 19.3944
R18902 GND.n7487 GND.n3106 19.3944
R18903 GND.n7487 GND.n7486 19.3944
R18904 GND.n7486 GND.n7485 19.3944
R18905 GND.n7485 GND.n3111 19.3944
R18906 GND.n7481 GND.n3111 19.3944
R18907 GND.n7481 GND.n7480 19.3944
R18908 GND.n7480 GND.n7479 19.3944
R18909 GND.n7479 GND.n3116 19.3944
R18910 GND.n7475 GND.n3116 19.3944
R18911 GND.n7475 GND.n7474 19.3944
R18912 GND.n7474 GND.n7473 19.3944
R18913 GND.n7473 GND.n3121 19.3944
R18914 GND.n7469 GND.n3121 19.3944
R18915 GND.n7469 GND.n7468 19.3944
R18916 GND.n7468 GND.n7467 19.3944
R18917 GND.n7467 GND.n3126 19.3944
R18918 GND.n7463 GND.n3126 19.3944
R18919 GND.n7463 GND.n7462 19.3944
R18920 GND.n7462 GND.n7461 19.3944
R18921 GND.n7461 GND.n3131 19.3944
R18922 GND.n7457 GND.n3131 19.3944
R18923 GND.n7457 GND.n7456 19.3944
R18924 GND.n7456 GND.n7455 19.3944
R18925 GND.n7455 GND.n3136 19.3944
R18926 GND.n7451 GND.n3136 19.3944
R18927 GND.n7451 GND.n7450 19.3944
R18928 GND.n7450 GND.n7449 19.3944
R18929 GND.n7449 GND.n3141 19.3944
R18930 GND.n7445 GND.n3141 19.3944
R18931 GND.n7445 GND.n7444 19.3944
R18932 GND.n7444 GND.n7443 19.3944
R18933 GND.n7443 GND.n3146 19.3944
R18934 GND.n7439 GND.n3146 19.3944
R18935 GND.n7439 GND.n7438 19.3944
R18936 GND.n7438 GND.n7437 19.3944
R18937 GND.n7437 GND.n3151 19.3944
R18938 GND.n7433 GND.n3151 19.3944
R18939 GND.n7433 GND.n7432 19.3944
R18940 GND.n7432 GND.n7431 19.3944
R18941 GND.n7431 GND.n3156 19.3944
R18942 GND.n7427 GND.n3156 19.3944
R18943 GND.n7427 GND.n7426 19.3944
R18944 GND.n7426 GND.n7425 19.3944
R18945 GND.n7425 GND.n3161 19.3944
R18946 GND.n7421 GND.n3161 19.3944
R18947 GND.n7421 GND.n7420 19.3944
R18948 GND.n7420 GND.n7419 19.3944
R18949 GND.n7419 GND.n3166 19.3944
R18950 GND.n7415 GND.n3166 19.3944
R18951 GND.n7415 GND.n7414 19.3944
R18952 GND.n7414 GND.n7413 19.3944
R18953 GND.n7413 GND.n3171 19.3944
R18954 GND.n7409 GND.n3171 19.3944
R18955 GND.n7409 GND.n7408 19.3944
R18956 GND.n7408 GND.n7407 19.3944
R18957 GND.n7407 GND.n3176 19.3944
R18958 GND.n7403 GND.n3176 19.3944
R18959 GND.n7403 GND.n7402 19.3944
R18960 GND.n7402 GND.n7401 19.3944
R18961 GND.n7401 GND.n3181 19.3944
R18962 GND.n7397 GND.n3181 19.3944
R18963 GND.n7397 GND.n7396 19.3944
R18964 GND.n7396 GND.n7395 19.3944
R18965 GND.n7395 GND.n3186 19.3944
R18966 GND.n7391 GND.n3186 19.3944
R18967 GND.n7391 GND.n7390 19.3944
R18968 GND.n7390 GND.n7389 19.3944
R18969 GND.n7389 GND.n3191 19.3944
R18970 GND.n7385 GND.n3191 19.3944
R18971 GND.n7385 GND.n7384 19.3944
R18972 GND.n7384 GND.n7383 19.3944
R18973 GND.n7383 GND.n3196 19.3944
R18974 GND.n7379 GND.n3196 19.3944
R18975 GND.n7379 GND.n7378 19.3944
R18976 GND.n7378 GND.n7377 19.3944
R18977 GND.n7377 GND.n3201 19.3944
R18978 GND.n7373 GND.n3201 19.3944
R18979 GND.n7373 GND.n7372 19.3944
R18980 GND.n7372 GND.n7371 19.3944
R18981 GND.n7371 GND.n3206 19.3944
R18982 GND.n7367 GND.n3206 19.3944
R18983 GND.n7367 GND.n7366 19.3944
R18984 GND.n7366 GND.n7365 19.3944
R18985 GND.n7365 GND.n3211 19.3944
R18986 GND.n7361 GND.n3211 19.3944
R18987 GND.n7361 GND.n7360 19.3944
R18988 GND.n7360 GND.n7359 19.3944
R18989 GND.n7359 GND.n3216 19.3944
R18990 GND.n7355 GND.n3216 19.3944
R18991 GND.n7355 GND.n7354 19.3944
R18992 GND.n7354 GND.n7353 19.3944
R18993 GND.n7353 GND.n3221 19.3944
R18994 GND.n7349 GND.n3221 19.3944
R18995 GND.n7349 GND.n7348 19.3944
R18996 GND.n7348 GND.n7347 19.3944
R18997 GND.n7347 GND.n3226 19.3944
R18998 GND.n7343 GND.n3226 19.3944
R18999 GND.n7287 GND.n3319 19.3944
R19000 GND.n7287 GND.n7286 19.3944
R19001 GND.n7286 GND.n3322 19.3944
R19002 GND.n7279 GND.n3322 19.3944
R19003 GND.n7279 GND.n7278 19.3944
R19004 GND.n7278 GND.n3332 19.3944
R19005 GND.n7271 GND.n3332 19.3944
R19006 GND.n7271 GND.n7270 19.3944
R19007 GND.n7270 GND.n3340 19.3944
R19008 GND.n7263 GND.n3340 19.3944
R19009 GND.n7263 GND.n7262 19.3944
R19010 GND.n7262 GND.n3352 19.3944
R19011 GND.n6427 GND.n3352 19.3944
R19012 GND.n6427 GND.n6426 19.3944
R19013 GND.n6426 GND.n6425 19.3944
R19014 GND.n6422 GND.n6421 19.3944
R19015 GND.n6421 GND.n6420 19.3944
R19016 GND.n6420 GND.n6418 19.3944
R19017 GND.n3046 GND.n3029 19.3944
R19018 GND.n3048 GND.n3046 19.3944
R19019 GND.n3049 GND.n3048 19.3944
R19020 GND.n7869 GND.n1836 19.3944
R19021 GND.n7864 GND.n1836 19.3944
R19022 GND.n7864 GND.n1851 19.3944
R19023 GND.n7857 GND.n1851 19.3944
R19024 GND.n7857 GND.n7856 19.3944
R19025 GND.n7856 GND.n1864 19.3944
R19026 GND.n7849 GND.n1864 19.3944
R19027 GND.n7849 GND.n7848 19.3944
R19028 GND.n7848 GND.n1874 19.3944
R19029 GND.n7841 GND.n1874 19.3944
R19030 GND.n7841 GND.n7840 19.3944
R19031 GND.n7840 GND.n1886 19.3944
R19032 GND.n3035 GND.n1886 19.3944
R19033 GND.n3036 GND.n3035 19.3944
R19034 GND.n3042 GND.n3036 19.3944
R19035 GND.n4663 GND.n4662 19.3944
R19036 GND.n4667 GND.n4662 19.3944
R19037 GND.n4667 GND.n4658 19.3944
R19038 GND.n4858 GND.n4658 19.3944
R19039 GND.n4858 GND.n4656 19.3944
R19040 GND.n4888 GND.n4656 19.3944
R19041 GND.n4888 GND.n4887 19.3944
R19042 GND.n4887 GND.n4886 19.3944
R19043 GND.n4886 GND.n4864 19.3944
R19044 GND.n4882 GND.n4864 19.3944
R19045 GND.n4882 GND.n4881 19.3944
R19046 GND.n4881 GND.n4880 19.3944
R19047 GND.n4880 GND.n4878 19.3944
R19048 GND.n4878 GND.n4877 19.3944
R19049 GND.n4877 GND.n4874 19.3944
R19050 GND.n4874 GND.n4873 19.3944
R19051 GND.n4873 GND.n4587 19.3944
R19052 GND.n5002 GND.n4587 19.3944
R19053 GND.n5002 GND.n4585 19.3944
R19054 GND.n5039 GND.n4585 19.3944
R19055 GND.n5039 GND.n5038 19.3944
R19056 GND.n5038 GND.n5037 19.3944
R19057 GND.n5037 GND.n5035 19.3944
R19058 GND.n5035 GND.n5034 19.3944
R19059 GND.n5034 GND.n5010 19.3944
R19060 GND.n5030 GND.n5010 19.3944
R19061 GND.n5030 GND.n5029 19.3944
R19062 GND.n5029 GND.n5028 19.3944
R19063 GND.n5028 GND.n5027 19.3944
R19064 GND.n5027 GND.n5026 19.3944
R19065 GND.n5026 GND.n5024 19.3944
R19066 GND.n5024 GND.n5023 19.3944
R19067 GND.n5023 GND.n5021 19.3944
R19068 GND.n5021 GND.n4501 19.3944
R19069 GND.n5165 GND.n4501 19.3944
R19070 GND.n5165 GND.n4499 19.3944
R19071 GND.n5203 GND.n4499 19.3944
R19072 GND.n5203 GND.n5202 19.3944
R19073 GND.n5202 GND.n5201 19.3944
R19074 GND.n5201 GND.n5199 19.3944
R19075 GND.n5199 GND.n5198 19.3944
R19076 GND.n5198 GND.n5173 19.3944
R19077 GND.n5194 GND.n5173 19.3944
R19078 GND.n5194 GND.n5193 19.3944
R19079 GND.n5193 GND.n5192 19.3944
R19080 GND.n5192 GND.n5191 19.3944
R19081 GND.n5191 GND.n5189 19.3944
R19082 GND.n5189 GND.n5188 19.3944
R19083 GND.n5188 GND.n5185 19.3944
R19084 GND.n5185 GND.n5184 19.3944
R19085 GND.n5184 GND.n4415 19.3944
R19086 GND.n5326 GND.n4415 19.3944
R19087 GND.n5326 GND.n4413 19.3944
R19088 GND.n5365 GND.n4413 19.3944
R19089 GND.n5365 GND.n5364 19.3944
R19090 GND.n5364 GND.n5363 19.3944
R19091 GND.n5363 GND.n5361 19.3944
R19092 GND.n5361 GND.n5360 19.3944
R19093 GND.n5360 GND.n5334 19.3944
R19094 GND.n5356 GND.n5334 19.3944
R19095 GND.n5356 GND.n5355 19.3944
R19096 GND.n5355 GND.n5354 19.3944
R19097 GND.n5354 GND.n5353 19.3944
R19098 GND.n5353 GND.n5350 19.3944
R19099 GND.n5350 GND.n5349 19.3944
R19100 GND.n5349 GND.n5346 19.3944
R19101 GND.n5346 GND.n5345 19.3944
R19102 GND.n5345 GND.n4329 19.3944
R19103 GND.n5486 GND.n4329 19.3944
R19104 GND.n5486 GND.n4327 19.3944
R19105 GND.n5535 GND.n4327 19.3944
R19106 GND.n5535 GND.n5534 19.3944
R19107 GND.n5534 GND.n5533 19.3944
R19108 GND.n5533 GND.n5531 19.3944
R19109 GND.n5531 GND.n5530 19.3944
R19110 GND.n5530 GND.n5494 19.3944
R19111 GND.n5526 GND.n5494 19.3944
R19112 GND.n5526 GND.n5525 19.3944
R19113 GND.n5525 GND.n5524 19.3944
R19114 GND.n5524 GND.n5523 19.3944
R19115 GND.n5523 GND.n5521 19.3944
R19116 GND.n5521 GND.n5520 19.3944
R19117 GND.n5520 GND.n5517 19.3944
R19118 GND.n5517 GND.n5516 19.3944
R19119 GND.n5516 GND.n5515 19.3944
R19120 GND.n5515 GND.n5513 19.3944
R19121 GND.n5513 GND.n5512 19.3944
R19122 GND.n5512 GND.n5510 19.3944
R19123 GND.n5510 GND.n4223 19.3944
R19124 GND.n5698 GND.n4223 19.3944
R19125 GND.n5698 GND.n4221 19.3944
R19126 GND.n5704 GND.n4221 19.3944
R19127 GND.n5704 GND.n5703 19.3944
R19128 GND.n5703 GND.n4199 19.3944
R19129 GND.n5732 GND.n4199 19.3944
R19130 GND.n5732 GND.n4197 19.3944
R19131 GND.n5791 GND.n4197 19.3944
R19132 GND.n5791 GND.n5790 19.3944
R19133 GND.n5790 GND.n5789 19.3944
R19134 GND.n5789 GND.n5787 19.3944
R19135 GND.n5787 GND.n5786 19.3944
R19136 GND.n5786 GND.n5740 19.3944
R19137 GND.n5782 GND.n5740 19.3944
R19138 GND.n5782 GND.n5781 19.3944
R19139 GND.n5781 GND.n5780 19.3944
R19140 GND.n5780 GND.n5779 19.3944
R19141 GND.n5779 GND.n5778 19.3944
R19142 GND.n5778 GND.n5776 19.3944
R19143 GND.n5776 GND.n5775 19.3944
R19144 GND.n5775 GND.n5750 19.3944
R19145 GND.n5771 GND.n5750 19.3944
R19146 GND.n5771 GND.n5770 19.3944
R19147 GND.n5770 GND.n5769 19.3944
R19148 GND.n5769 GND.n5768 19.3944
R19149 GND.n5768 GND.n5766 19.3944
R19150 GND.n5766 GND.n5765 19.3944
R19151 GND.n5765 GND.n5762 19.3944
R19152 GND.n5762 GND.n5761 19.3944
R19153 GND.n5761 GND.n4073 19.3944
R19154 GND.n5972 GND.n4073 19.3944
R19155 GND.n5972 GND.n4071 19.3944
R19156 GND.n5999 GND.n4071 19.3944
R19157 GND.n5999 GND.n5998 19.3944
R19158 GND.n5998 GND.n5997 19.3944
R19159 GND.n5997 GND.n5995 19.3944
R19160 GND.n5995 GND.n5994 19.3944
R19161 GND.n5994 GND.n5980 19.3944
R19162 GND.n5990 GND.n5980 19.3944
R19163 GND.n5990 GND.n5989 19.3944
R19164 GND.n5989 GND.n5988 19.3944
R19165 GND.n5988 GND.n5987 19.3944
R19166 GND.n5987 GND.n4009 19.3944
R19167 GND.n6097 GND.n4009 19.3944
R19168 GND.n6097 GND.n4007 19.3944
R19169 GND.n6339 GND.n4007 19.3944
R19170 GND.n6339 GND.n6338 19.3944
R19171 GND.n6338 GND.n6337 19.3944
R19172 GND.n6337 GND.n6335 19.3944
R19173 GND.n6335 GND.n6334 19.3944
R19174 GND.n6334 GND.n6331 19.3944
R19175 GND.n6331 GND.n6330 19.3944
R19176 GND.n9326 GND.n698 19.3944
R19177 GND.n9326 GND.n696 19.3944
R19178 GND.n9330 GND.n696 19.3944
R19179 GND.n9330 GND.n692 19.3944
R19180 GND.n9336 GND.n692 19.3944
R19181 GND.n9336 GND.n690 19.3944
R19182 GND.n9340 GND.n690 19.3944
R19183 GND.n9340 GND.n686 19.3944
R19184 GND.n9346 GND.n686 19.3944
R19185 GND.n9346 GND.n684 19.3944
R19186 GND.n9350 GND.n684 19.3944
R19187 GND.n9350 GND.n680 19.3944
R19188 GND.n9356 GND.n680 19.3944
R19189 GND.n9356 GND.n678 19.3944
R19190 GND.n9360 GND.n678 19.3944
R19191 GND.n9360 GND.n674 19.3944
R19192 GND.n9366 GND.n674 19.3944
R19193 GND.n9366 GND.n672 19.3944
R19194 GND.n9370 GND.n672 19.3944
R19195 GND.n9370 GND.n668 19.3944
R19196 GND.n9376 GND.n668 19.3944
R19197 GND.n9376 GND.n666 19.3944
R19198 GND.n9380 GND.n666 19.3944
R19199 GND.n9380 GND.n662 19.3944
R19200 GND.n9386 GND.n662 19.3944
R19201 GND.n9386 GND.n660 19.3944
R19202 GND.n9390 GND.n660 19.3944
R19203 GND.n9390 GND.n656 19.3944
R19204 GND.n9396 GND.n656 19.3944
R19205 GND.n9396 GND.n654 19.3944
R19206 GND.n9400 GND.n654 19.3944
R19207 GND.n9400 GND.n650 19.3944
R19208 GND.n9406 GND.n650 19.3944
R19209 GND.n9406 GND.n648 19.3944
R19210 GND.n9410 GND.n648 19.3944
R19211 GND.n9410 GND.n644 19.3944
R19212 GND.n9416 GND.n644 19.3944
R19213 GND.n9416 GND.n642 19.3944
R19214 GND.n9420 GND.n642 19.3944
R19215 GND.n9420 GND.n638 19.3944
R19216 GND.n9426 GND.n638 19.3944
R19217 GND.n9426 GND.n636 19.3944
R19218 GND.n9430 GND.n636 19.3944
R19219 GND.n9430 GND.n632 19.3944
R19220 GND.n9436 GND.n632 19.3944
R19221 GND.n9436 GND.n630 19.3944
R19222 GND.n9440 GND.n630 19.3944
R19223 GND.n9440 GND.n626 19.3944
R19224 GND.n9446 GND.n626 19.3944
R19225 GND.n9446 GND.n624 19.3944
R19226 GND.n9451 GND.n624 19.3944
R19227 GND.n9451 GND.n620 19.3944
R19228 GND.n9457 GND.n620 19.3944
R19229 GND.n9458 GND.n9457 19.3944
R19230 GND.n8290 GND.n1320 19.3944
R19231 GND.n8290 GND.n1316 19.3944
R19232 GND.n8296 GND.n1316 19.3944
R19233 GND.n8296 GND.n1314 19.3944
R19234 GND.n8300 GND.n1314 19.3944
R19235 GND.n8300 GND.n1310 19.3944
R19236 GND.n8306 GND.n1310 19.3944
R19237 GND.n8306 GND.n1308 19.3944
R19238 GND.n8310 GND.n1308 19.3944
R19239 GND.n8310 GND.n1304 19.3944
R19240 GND.n8316 GND.n1304 19.3944
R19241 GND.n8316 GND.n1302 19.3944
R19242 GND.n8320 GND.n1302 19.3944
R19243 GND.n8320 GND.n1298 19.3944
R19244 GND.n8326 GND.n1298 19.3944
R19245 GND.n8326 GND.n1296 19.3944
R19246 GND.n8330 GND.n1296 19.3944
R19247 GND.n8330 GND.n1292 19.3944
R19248 GND.n8336 GND.n1292 19.3944
R19249 GND.n8336 GND.n1290 19.3944
R19250 GND.n8340 GND.n1290 19.3944
R19251 GND.n8340 GND.n1286 19.3944
R19252 GND.n8346 GND.n1286 19.3944
R19253 GND.n8346 GND.n1284 19.3944
R19254 GND.n8350 GND.n1284 19.3944
R19255 GND.n8350 GND.n1280 19.3944
R19256 GND.n8356 GND.n1280 19.3944
R19257 GND.n8356 GND.n1278 19.3944
R19258 GND.n8360 GND.n1278 19.3944
R19259 GND.n8360 GND.n1274 19.3944
R19260 GND.n8366 GND.n1274 19.3944
R19261 GND.n8366 GND.n1272 19.3944
R19262 GND.n8370 GND.n1272 19.3944
R19263 GND.n8370 GND.n1268 19.3944
R19264 GND.n8376 GND.n1268 19.3944
R19265 GND.n8376 GND.n1266 19.3944
R19266 GND.n8380 GND.n1266 19.3944
R19267 GND.n8380 GND.n1262 19.3944
R19268 GND.n8386 GND.n1262 19.3944
R19269 GND.n8386 GND.n1260 19.3944
R19270 GND.n8390 GND.n1260 19.3944
R19271 GND.n8390 GND.n1256 19.3944
R19272 GND.n8396 GND.n1256 19.3944
R19273 GND.n8396 GND.n1254 19.3944
R19274 GND.n8400 GND.n1254 19.3944
R19275 GND.n8400 GND.n1250 19.3944
R19276 GND.n8406 GND.n1250 19.3944
R19277 GND.n8406 GND.n1248 19.3944
R19278 GND.n8410 GND.n1248 19.3944
R19279 GND.n8410 GND.n1244 19.3944
R19280 GND.n8416 GND.n1244 19.3944
R19281 GND.n8416 GND.n1242 19.3944
R19282 GND.n8420 GND.n1242 19.3944
R19283 GND.n8420 GND.n1238 19.3944
R19284 GND.n8426 GND.n1238 19.3944
R19285 GND.n8426 GND.n1236 19.3944
R19286 GND.n8430 GND.n1236 19.3944
R19287 GND.n8430 GND.n1232 19.3944
R19288 GND.n8436 GND.n1232 19.3944
R19289 GND.n8436 GND.n1230 19.3944
R19290 GND.n8440 GND.n1230 19.3944
R19291 GND.n8440 GND.n1226 19.3944
R19292 GND.n8446 GND.n1226 19.3944
R19293 GND.n8446 GND.n1224 19.3944
R19294 GND.n8450 GND.n1224 19.3944
R19295 GND.n8450 GND.n1220 19.3944
R19296 GND.n8456 GND.n1220 19.3944
R19297 GND.n8456 GND.n1218 19.3944
R19298 GND.n8460 GND.n1218 19.3944
R19299 GND.n8460 GND.n1214 19.3944
R19300 GND.n8466 GND.n1214 19.3944
R19301 GND.n8466 GND.n1212 19.3944
R19302 GND.n8470 GND.n1212 19.3944
R19303 GND.n8470 GND.n1208 19.3944
R19304 GND.n8476 GND.n1208 19.3944
R19305 GND.n8476 GND.n1206 19.3944
R19306 GND.n8480 GND.n1206 19.3944
R19307 GND.n8480 GND.n1202 19.3944
R19308 GND.n8486 GND.n1202 19.3944
R19309 GND.n8486 GND.n1200 19.3944
R19310 GND.n8490 GND.n1200 19.3944
R19311 GND.n8490 GND.n1196 19.3944
R19312 GND.n8496 GND.n1196 19.3944
R19313 GND.n8496 GND.n1194 19.3944
R19314 GND.n8500 GND.n1194 19.3944
R19315 GND.n8500 GND.n1190 19.3944
R19316 GND.n8506 GND.n1190 19.3944
R19317 GND.n8506 GND.n1188 19.3944
R19318 GND.n8510 GND.n1188 19.3944
R19319 GND.n8510 GND.n1184 19.3944
R19320 GND.n8516 GND.n1184 19.3944
R19321 GND.n8516 GND.n1182 19.3944
R19322 GND.n8520 GND.n1182 19.3944
R19323 GND.n8520 GND.n1178 19.3944
R19324 GND.n8526 GND.n1178 19.3944
R19325 GND.n8526 GND.n1176 19.3944
R19326 GND.n8530 GND.n1176 19.3944
R19327 GND.n8530 GND.n1172 19.3944
R19328 GND.n8536 GND.n1172 19.3944
R19329 GND.n8536 GND.n1170 19.3944
R19330 GND.n8540 GND.n1170 19.3944
R19331 GND.n8540 GND.n1166 19.3944
R19332 GND.n8546 GND.n1166 19.3944
R19333 GND.n8546 GND.n1164 19.3944
R19334 GND.n8550 GND.n1164 19.3944
R19335 GND.n8550 GND.n1160 19.3944
R19336 GND.n8556 GND.n1160 19.3944
R19337 GND.n8556 GND.n1158 19.3944
R19338 GND.n8560 GND.n1158 19.3944
R19339 GND.n8560 GND.n1154 19.3944
R19340 GND.n8566 GND.n1154 19.3944
R19341 GND.n8566 GND.n1152 19.3944
R19342 GND.n8570 GND.n1152 19.3944
R19343 GND.n8570 GND.n1148 19.3944
R19344 GND.n8576 GND.n1148 19.3944
R19345 GND.n8576 GND.n1146 19.3944
R19346 GND.n8580 GND.n1146 19.3944
R19347 GND.n8580 GND.n1142 19.3944
R19348 GND.n8586 GND.n1142 19.3944
R19349 GND.n8586 GND.n1140 19.3944
R19350 GND.n8590 GND.n1140 19.3944
R19351 GND.n8590 GND.n1136 19.3944
R19352 GND.n8596 GND.n1136 19.3944
R19353 GND.n8596 GND.n1134 19.3944
R19354 GND.n8600 GND.n1134 19.3944
R19355 GND.n8600 GND.n1130 19.3944
R19356 GND.n8606 GND.n1130 19.3944
R19357 GND.n8606 GND.n1128 19.3944
R19358 GND.n8610 GND.n1128 19.3944
R19359 GND.n8610 GND.n1124 19.3944
R19360 GND.n8616 GND.n1124 19.3944
R19361 GND.n8616 GND.n1122 19.3944
R19362 GND.n8620 GND.n1122 19.3944
R19363 GND.n8620 GND.n1118 19.3944
R19364 GND.n8626 GND.n1118 19.3944
R19365 GND.n8626 GND.n1116 19.3944
R19366 GND.n8630 GND.n1116 19.3944
R19367 GND.n8630 GND.n1112 19.3944
R19368 GND.n8636 GND.n1112 19.3944
R19369 GND.n8636 GND.n1110 19.3944
R19370 GND.n8640 GND.n1110 19.3944
R19371 GND.n8640 GND.n1106 19.3944
R19372 GND.n8646 GND.n1106 19.3944
R19373 GND.n8646 GND.n1104 19.3944
R19374 GND.n8650 GND.n1104 19.3944
R19375 GND.n8650 GND.n1100 19.3944
R19376 GND.n8656 GND.n1100 19.3944
R19377 GND.n8656 GND.n1098 19.3944
R19378 GND.n8660 GND.n1098 19.3944
R19379 GND.n8660 GND.n1094 19.3944
R19380 GND.n8666 GND.n1094 19.3944
R19381 GND.n8666 GND.n1092 19.3944
R19382 GND.n8670 GND.n1092 19.3944
R19383 GND.n8670 GND.n1088 19.3944
R19384 GND.n8676 GND.n1088 19.3944
R19385 GND.n8676 GND.n1086 19.3944
R19386 GND.n8680 GND.n1086 19.3944
R19387 GND.n8680 GND.n1082 19.3944
R19388 GND.n8686 GND.n1082 19.3944
R19389 GND.n8686 GND.n1080 19.3944
R19390 GND.n8690 GND.n1080 19.3944
R19391 GND.n8690 GND.n1076 19.3944
R19392 GND.n8696 GND.n1076 19.3944
R19393 GND.n8696 GND.n1074 19.3944
R19394 GND.n8700 GND.n1074 19.3944
R19395 GND.n8700 GND.n1070 19.3944
R19396 GND.n8706 GND.n1070 19.3944
R19397 GND.n8706 GND.n1068 19.3944
R19398 GND.n8710 GND.n1068 19.3944
R19399 GND.n8710 GND.n1064 19.3944
R19400 GND.n8716 GND.n1064 19.3944
R19401 GND.n8716 GND.n1062 19.3944
R19402 GND.n8720 GND.n1062 19.3944
R19403 GND.n8720 GND.n1058 19.3944
R19404 GND.n8726 GND.n1058 19.3944
R19405 GND.n8726 GND.n1056 19.3944
R19406 GND.n8730 GND.n1056 19.3944
R19407 GND.n8730 GND.n1052 19.3944
R19408 GND.n8736 GND.n1052 19.3944
R19409 GND.n8736 GND.n1050 19.3944
R19410 GND.n8740 GND.n1050 19.3944
R19411 GND.n8740 GND.n1046 19.3944
R19412 GND.n8746 GND.n1046 19.3944
R19413 GND.n8746 GND.n1044 19.3944
R19414 GND.n8750 GND.n1044 19.3944
R19415 GND.n8750 GND.n1040 19.3944
R19416 GND.n8756 GND.n1040 19.3944
R19417 GND.n8756 GND.n1038 19.3944
R19418 GND.n8760 GND.n1038 19.3944
R19419 GND.n8760 GND.n1034 19.3944
R19420 GND.n8766 GND.n1034 19.3944
R19421 GND.n8766 GND.n1032 19.3944
R19422 GND.n8770 GND.n1032 19.3944
R19423 GND.n8770 GND.n1028 19.3944
R19424 GND.n8776 GND.n1028 19.3944
R19425 GND.n8776 GND.n1026 19.3944
R19426 GND.n8780 GND.n1026 19.3944
R19427 GND.n8780 GND.n1022 19.3944
R19428 GND.n8786 GND.n1022 19.3944
R19429 GND.n8786 GND.n1020 19.3944
R19430 GND.n8790 GND.n1020 19.3944
R19431 GND.n8790 GND.n1016 19.3944
R19432 GND.n8796 GND.n1016 19.3944
R19433 GND.n8796 GND.n1014 19.3944
R19434 GND.n8800 GND.n1014 19.3944
R19435 GND.n8800 GND.n1010 19.3944
R19436 GND.n8806 GND.n1010 19.3944
R19437 GND.n8806 GND.n1008 19.3944
R19438 GND.n8810 GND.n1008 19.3944
R19439 GND.n8810 GND.n1004 19.3944
R19440 GND.n8816 GND.n1004 19.3944
R19441 GND.n8816 GND.n1002 19.3944
R19442 GND.n8820 GND.n1002 19.3944
R19443 GND.n8820 GND.n998 19.3944
R19444 GND.n8826 GND.n998 19.3944
R19445 GND.n8826 GND.n996 19.3944
R19446 GND.n8830 GND.n996 19.3944
R19447 GND.n8830 GND.n992 19.3944
R19448 GND.n8836 GND.n992 19.3944
R19449 GND.n8836 GND.n990 19.3944
R19450 GND.n8840 GND.n990 19.3944
R19451 GND.n8840 GND.n986 19.3944
R19452 GND.n8846 GND.n986 19.3944
R19453 GND.n8846 GND.n984 19.3944
R19454 GND.n8850 GND.n984 19.3944
R19455 GND.n8850 GND.n980 19.3944
R19456 GND.n8856 GND.n980 19.3944
R19457 GND.n8856 GND.n978 19.3944
R19458 GND.n8860 GND.n978 19.3944
R19459 GND.n8860 GND.n974 19.3944
R19460 GND.n8866 GND.n974 19.3944
R19461 GND.n8866 GND.n972 19.3944
R19462 GND.n8870 GND.n972 19.3944
R19463 GND.n8870 GND.n968 19.3944
R19464 GND.n8876 GND.n968 19.3944
R19465 GND.n8876 GND.n966 19.3944
R19466 GND.n8880 GND.n966 19.3944
R19467 GND.n8880 GND.n962 19.3944
R19468 GND.n8886 GND.n962 19.3944
R19469 GND.n8886 GND.n960 19.3944
R19470 GND.n8890 GND.n960 19.3944
R19471 GND.n8890 GND.n956 19.3944
R19472 GND.n8896 GND.n956 19.3944
R19473 GND.n8896 GND.n954 19.3944
R19474 GND.n8900 GND.n954 19.3944
R19475 GND.n8900 GND.n950 19.3944
R19476 GND.n8906 GND.n950 19.3944
R19477 GND.n8906 GND.n948 19.3944
R19478 GND.n8910 GND.n948 19.3944
R19479 GND.n8910 GND.n944 19.3944
R19480 GND.n8916 GND.n944 19.3944
R19481 GND.n8916 GND.n942 19.3944
R19482 GND.n8920 GND.n942 19.3944
R19483 GND.n8920 GND.n938 19.3944
R19484 GND.n8926 GND.n938 19.3944
R19485 GND.n8926 GND.n936 19.3944
R19486 GND.n8930 GND.n936 19.3944
R19487 GND.n8930 GND.n932 19.3944
R19488 GND.n8936 GND.n932 19.3944
R19489 GND.n8936 GND.n930 19.3944
R19490 GND.n8940 GND.n930 19.3944
R19491 GND.n8940 GND.n926 19.3944
R19492 GND.n8946 GND.n926 19.3944
R19493 GND.n8946 GND.n924 19.3944
R19494 GND.n8950 GND.n924 19.3944
R19495 GND.n8950 GND.n920 19.3944
R19496 GND.n8956 GND.n920 19.3944
R19497 GND.n8956 GND.n918 19.3944
R19498 GND.n8960 GND.n918 19.3944
R19499 GND.n8960 GND.n914 19.3944
R19500 GND.n8966 GND.n914 19.3944
R19501 GND.n8966 GND.n912 19.3944
R19502 GND.n8970 GND.n912 19.3944
R19503 GND.n8970 GND.n908 19.3944
R19504 GND.n8976 GND.n908 19.3944
R19505 GND.n8976 GND.n906 19.3944
R19506 GND.n8980 GND.n906 19.3944
R19507 GND.n8980 GND.n902 19.3944
R19508 GND.n8986 GND.n902 19.3944
R19509 GND.n8986 GND.n900 19.3944
R19510 GND.n8990 GND.n900 19.3944
R19511 GND.n8990 GND.n896 19.3944
R19512 GND.n8996 GND.n896 19.3944
R19513 GND.n8996 GND.n894 19.3944
R19514 GND.n9000 GND.n894 19.3944
R19515 GND.n9000 GND.n890 19.3944
R19516 GND.n9006 GND.n890 19.3944
R19517 GND.n9006 GND.n888 19.3944
R19518 GND.n9010 GND.n888 19.3944
R19519 GND.n9010 GND.n884 19.3944
R19520 GND.n9016 GND.n884 19.3944
R19521 GND.n9016 GND.n882 19.3944
R19522 GND.n9020 GND.n882 19.3944
R19523 GND.n9020 GND.n878 19.3944
R19524 GND.n9026 GND.n878 19.3944
R19525 GND.n9026 GND.n876 19.3944
R19526 GND.n9030 GND.n876 19.3944
R19527 GND.n9030 GND.n872 19.3944
R19528 GND.n9036 GND.n872 19.3944
R19529 GND.n9036 GND.n870 19.3944
R19530 GND.n9040 GND.n870 19.3944
R19531 GND.n9040 GND.n866 19.3944
R19532 GND.n9046 GND.n866 19.3944
R19533 GND.n9046 GND.n864 19.3944
R19534 GND.n9050 GND.n864 19.3944
R19535 GND.n9050 GND.n860 19.3944
R19536 GND.n9056 GND.n860 19.3944
R19537 GND.n9056 GND.n858 19.3944
R19538 GND.n9060 GND.n858 19.3944
R19539 GND.n9060 GND.n854 19.3944
R19540 GND.n9066 GND.n854 19.3944
R19541 GND.n9066 GND.n852 19.3944
R19542 GND.n9070 GND.n852 19.3944
R19543 GND.n9070 GND.n848 19.3944
R19544 GND.n9076 GND.n848 19.3944
R19545 GND.n9076 GND.n846 19.3944
R19546 GND.n9080 GND.n846 19.3944
R19547 GND.n9080 GND.n842 19.3944
R19548 GND.n9086 GND.n842 19.3944
R19549 GND.n9086 GND.n840 19.3944
R19550 GND.n9090 GND.n840 19.3944
R19551 GND.n9090 GND.n836 19.3944
R19552 GND.n9096 GND.n836 19.3944
R19553 GND.n9096 GND.n834 19.3944
R19554 GND.n9100 GND.n834 19.3944
R19555 GND.n9100 GND.n830 19.3944
R19556 GND.n9106 GND.n830 19.3944
R19557 GND.n9106 GND.n828 19.3944
R19558 GND.n9110 GND.n828 19.3944
R19559 GND.n9110 GND.n824 19.3944
R19560 GND.n9116 GND.n824 19.3944
R19561 GND.n9116 GND.n822 19.3944
R19562 GND.n9120 GND.n822 19.3944
R19563 GND.n9120 GND.n818 19.3944
R19564 GND.n9126 GND.n818 19.3944
R19565 GND.n9126 GND.n816 19.3944
R19566 GND.n9130 GND.n816 19.3944
R19567 GND.n9130 GND.n812 19.3944
R19568 GND.n9136 GND.n812 19.3944
R19569 GND.n9136 GND.n810 19.3944
R19570 GND.n9140 GND.n810 19.3944
R19571 GND.n9140 GND.n806 19.3944
R19572 GND.n9146 GND.n806 19.3944
R19573 GND.n9146 GND.n804 19.3944
R19574 GND.n9150 GND.n804 19.3944
R19575 GND.n9150 GND.n800 19.3944
R19576 GND.n9156 GND.n800 19.3944
R19577 GND.n9156 GND.n798 19.3944
R19578 GND.n9160 GND.n798 19.3944
R19579 GND.n9160 GND.n794 19.3944
R19580 GND.n9166 GND.n794 19.3944
R19581 GND.n9166 GND.n792 19.3944
R19582 GND.n9170 GND.n792 19.3944
R19583 GND.n9170 GND.n788 19.3944
R19584 GND.n9176 GND.n788 19.3944
R19585 GND.n9176 GND.n786 19.3944
R19586 GND.n9180 GND.n786 19.3944
R19587 GND.n9180 GND.n782 19.3944
R19588 GND.n9186 GND.n782 19.3944
R19589 GND.n9186 GND.n780 19.3944
R19590 GND.n9190 GND.n780 19.3944
R19591 GND.n9190 GND.n776 19.3944
R19592 GND.n9196 GND.n776 19.3944
R19593 GND.n9196 GND.n774 19.3944
R19594 GND.n9200 GND.n774 19.3944
R19595 GND.n9200 GND.n770 19.3944
R19596 GND.n9206 GND.n770 19.3944
R19597 GND.n9206 GND.n768 19.3944
R19598 GND.n9210 GND.n768 19.3944
R19599 GND.n9210 GND.n764 19.3944
R19600 GND.n9216 GND.n764 19.3944
R19601 GND.n9216 GND.n762 19.3944
R19602 GND.n9220 GND.n762 19.3944
R19603 GND.n9220 GND.n758 19.3944
R19604 GND.n9226 GND.n758 19.3944
R19605 GND.n9226 GND.n756 19.3944
R19606 GND.n9230 GND.n756 19.3944
R19607 GND.n9230 GND.n752 19.3944
R19608 GND.n9236 GND.n752 19.3944
R19609 GND.n9236 GND.n750 19.3944
R19610 GND.n9240 GND.n750 19.3944
R19611 GND.n9240 GND.n746 19.3944
R19612 GND.n9246 GND.n746 19.3944
R19613 GND.n9246 GND.n744 19.3944
R19614 GND.n9250 GND.n744 19.3944
R19615 GND.n9250 GND.n740 19.3944
R19616 GND.n9256 GND.n740 19.3944
R19617 GND.n9256 GND.n738 19.3944
R19618 GND.n9260 GND.n738 19.3944
R19619 GND.n9260 GND.n734 19.3944
R19620 GND.n9266 GND.n734 19.3944
R19621 GND.n9266 GND.n732 19.3944
R19622 GND.n9270 GND.n732 19.3944
R19623 GND.n9270 GND.n728 19.3944
R19624 GND.n9276 GND.n728 19.3944
R19625 GND.n9276 GND.n726 19.3944
R19626 GND.n9280 GND.n726 19.3944
R19627 GND.n9280 GND.n722 19.3944
R19628 GND.n9286 GND.n722 19.3944
R19629 GND.n9286 GND.n720 19.3944
R19630 GND.n9290 GND.n720 19.3944
R19631 GND.n9290 GND.n716 19.3944
R19632 GND.n9296 GND.n716 19.3944
R19633 GND.n9296 GND.n714 19.3944
R19634 GND.n9300 GND.n714 19.3944
R19635 GND.n9300 GND.n710 19.3944
R19636 GND.n9306 GND.n710 19.3944
R19637 GND.n9306 GND.n708 19.3944
R19638 GND.n9310 GND.n708 19.3944
R19639 GND.n9310 GND.n704 19.3944
R19640 GND.n9316 GND.n704 19.3944
R19641 GND.n9316 GND.n702 19.3944
R19642 GND.n9320 GND.n702 19.3944
R19643 GND.n6266 GND.n6265 19.3944
R19644 GND.n6272 GND.n6265 19.3944
R19645 GND.n6273 GND.n6272 19.3944
R19646 GND.n6276 GND.n6273 19.3944
R19647 GND.n6276 GND.n6263 19.3944
R19648 GND.n6282 GND.n6263 19.3944
R19649 GND.n6283 GND.n6282 19.3944
R19650 GND.n6286 GND.n6283 19.3944
R19651 GND.n6286 GND.n6119 19.3944
R19652 GND.n6296 GND.n6293 19.3944
R19653 GND.n6296 GND.n6116 19.3944
R19654 GND.n6302 GND.n6116 19.3944
R19655 GND.n6303 GND.n6302 19.3944
R19656 GND.n6306 GND.n6303 19.3944
R19657 GND.n6306 GND.n6114 19.3944
R19658 GND.n6312 GND.n6114 19.3944
R19659 GND.n6313 GND.n6312 19.3944
R19660 GND.n6316 GND.n6313 19.3944
R19661 GND.n6316 GND.n6110 19.3944
R19662 GND.n6320 GND.n6110 19.3944
R19663 GND.n7254 GND.n7253 19.3944
R19664 GND.n7253 GND.n7252 19.3944
R19665 GND.n7252 GND.n3364 19.3944
R19666 GND.n6586 GND.n3364 19.3944
R19667 GND.n6592 GND.n6586 19.3944
R19668 GND.n6592 GND.n6591 19.3944
R19669 GND.n6591 GND.n3945 19.3944
R19670 GND.n6611 GND.n3945 19.3944
R19671 GND.n6611 GND.n3943 19.3944
R19672 GND.n6617 GND.n3943 19.3944
R19673 GND.n6617 GND.n6616 19.3944
R19674 GND.n6616 GND.n3922 19.3944
R19675 GND.n6635 GND.n3922 19.3944
R19676 GND.n6635 GND.n3920 19.3944
R19677 GND.n6641 GND.n3920 19.3944
R19678 GND.n6641 GND.n6640 19.3944
R19679 GND.n6640 GND.n3899 19.3944
R19680 GND.n6660 GND.n3899 19.3944
R19681 GND.n6660 GND.n3897 19.3944
R19682 GND.n6666 GND.n3897 19.3944
R19683 GND.n6666 GND.n6665 19.3944
R19684 GND.n6665 GND.n3877 19.3944
R19685 GND.n6685 GND.n3877 19.3944
R19686 GND.n6685 GND.n3875 19.3944
R19687 GND.n6691 GND.n3875 19.3944
R19688 GND.n6691 GND.n6690 19.3944
R19689 GND.n6690 GND.n3854 19.3944
R19690 GND.n6710 GND.n3854 19.3944
R19691 GND.n6710 GND.n3852 19.3944
R19692 GND.n6716 GND.n3852 19.3944
R19693 GND.n6716 GND.n6715 19.3944
R19694 GND.n6715 GND.n3831 19.3944
R19695 GND.n6734 GND.n3831 19.3944
R19696 GND.n6734 GND.n3829 19.3944
R19697 GND.n6740 GND.n3829 19.3944
R19698 GND.n6740 GND.n6739 19.3944
R19699 GND.n6739 GND.n3808 19.3944
R19700 GND.n6759 GND.n3808 19.3944
R19701 GND.n6759 GND.n3806 19.3944
R19702 GND.n6765 GND.n3806 19.3944
R19703 GND.n6765 GND.n6764 19.3944
R19704 GND.n6764 GND.n3786 19.3944
R19705 GND.n6784 GND.n3786 19.3944
R19706 GND.n6784 GND.n3784 19.3944
R19707 GND.n6791 GND.n3784 19.3944
R19708 GND.n6791 GND.n6790 19.3944
R19709 GND.n6790 GND.n3756 19.3944
R19710 GND.n6875 GND.n3756 19.3944
R19711 GND.n6873 GND.n6872 19.3944
R19712 GND.n6872 GND.n3757 19.3944
R19713 GND.n6858 GND.n6823 19.3944
R19714 GND.n6856 GND.n6855 19.3944
R19715 GND.n6838 GND.n6835 19.3944
R19716 GND.n6838 GND.n6837 19.3944
R19717 GND.n6837 GND.n3728 19.3944
R19718 GND.n6894 GND.n3728 19.3944
R19719 GND.n6894 GND.n3726 19.3944
R19720 GND.n6900 GND.n3726 19.3944
R19721 GND.n6900 GND.n6899 19.3944
R19722 GND.n6899 GND.n3706 19.3944
R19723 GND.n6921 GND.n3706 19.3944
R19724 GND.n6921 GND.n3704 19.3944
R19725 GND.n6927 GND.n3704 19.3944
R19726 GND.n6927 GND.n6926 19.3944
R19727 GND.n6926 GND.n3685 19.3944
R19728 GND.n6950 GND.n3685 19.3944
R19729 GND.n6950 GND.n3683 19.3944
R19730 GND.n6956 GND.n3683 19.3944
R19731 GND.n6956 GND.n6955 19.3944
R19732 GND.n6955 GND.n3665 19.3944
R19733 GND.n6977 GND.n3665 19.3944
R19734 GND.n6977 GND.n3663 19.3944
R19735 GND.n6983 GND.n3663 19.3944
R19736 GND.n6983 GND.n6982 19.3944
R19737 GND.n6982 GND.n3642 19.3944
R19738 GND.n7003 GND.n3642 19.3944
R19739 GND.n7003 GND.n3640 19.3944
R19740 GND.n7009 GND.n3640 19.3944
R19741 GND.n7009 GND.n7008 19.3944
R19742 GND.n7008 GND.n3620 19.3944
R19743 GND.n7030 GND.n3620 19.3944
R19744 GND.n7030 GND.n3618 19.3944
R19745 GND.n7036 GND.n3618 19.3944
R19746 GND.n7036 GND.n7035 19.3944
R19747 GND.n7035 GND.n3599 19.3944
R19748 GND.n7058 GND.n3599 19.3944
R19749 GND.n7058 GND.n3597 19.3944
R19750 GND.n7064 GND.n3597 19.3944
R19751 GND.n7064 GND.n7063 19.3944
R19752 GND.n7063 GND.n3576 19.3944
R19753 GND.n7091 GND.n3576 19.3944
R19754 GND.n7091 GND.n3574 19.3944
R19755 GND.n7097 GND.n3574 19.3944
R19756 GND.n7097 GND.n7096 19.3944
R19757 GND.n7096 GND.n565 19.3944
R19758 GND.n9508 GND.n565 19.3944
R19759 GND.n9508 GND.n563 19.3944
R19760 GND.n9514 GND.n563 19.3944
R19761 GND.n9514 GND.n9513 19.3944
R19762 GND.n9513 GND.n482 19.3944
R19763 GND.n9610 GND.n482 19.3944
R19764 GND.n8148 GND.n8147 19.3944
R19765 GND.n8147 GND.n8146 19.3944
R19766 GND.n8146 GND.n8145 19.3944
R19767 GND.n8145 GND.n8143 19.3944
R19768 GND.n8143 GND.n8140 19.3944
R19769 GND.n8140 GND.n8139 19.3944
R19770 GND.n8139 GND.n8136 19.3944
R19771 GND.n8136 GND.n8135 19.3944
R19772 GND.n8135 GND.n8132 19.3944
R19773 GND.n8132 GND.n8131 19.3944
R19774 GND.n8127 GND.n8124 19.3944
R19775 GND.n8124 GND.n8123 19.3944
R19776 GND.n8123 GND.n8120 19.3944
R19777 GND.n8120 GND.n8119 19.3944
R19778 GND.n8119 GND.n8116 19.3944
R19779 GND.n8116 GND.n8115 19.3944
R19780 GND.n8115 GND.n8112 19.3944
R19781 GND.n8112 GND.n8111 19.3944
R19782 GND.n8111 GND.n8108 19.3944
R19783 GND.n8108 GND.n8107 19.3944
R19784 GND.n8107 GND.n8104 19.3944
R19785 GND.n1538 GND.n1536 19.3944
R19786 GND.n1538 GND.n1534 19.3944
R19787 GND.n8084 GND.n1534 19.3944
R19788 GND.n8084 GND.n8083 19.3944
R19789 GND.n8083 GND.n8082 19.3944
R19790 GND.n8082 GND.n1544 19.3944
R19791 GND.n2512 GND.n1544 19.3944
R19792 GND.n2512 GND.n2511 19.3944
R19793 GND.n2511 GND.n2358 19.3944
R19794 GND.n2531 GND.n2358 19.3944
R19795 GND.n2531 GND.n2356 19.3944
R19796 GND.n2537 GND.n2356 19.3944
R19797 GND.n2537 GND.n2536 19.3944
R19798 GND.n2536 GND.n2335 19.3944
R19799 GND.n2556 GND.n2335 19.3944
R19800 GND.n2556 GND.n2333 19.3944
R19801 GND.n2562 GND.n2333 19.3944
R19802 GND.n2562 GND.n2561 19.3944
R19803 GND.n2561 GND.n2312 19.3944
R19804 GND.n2580 GND.n2312 19.3944
R19805 GND.n2580 GND.n2310 19.3944
R19806 GND.n2586 GND.n2310 19.3944
R19807 GND.n2586 GND.n2585 19.3944
R19808 GND.n2585 GND.n2289 19.3944
R19809 GND.n2605 GND.n2289 19.3944
R19810 GND.n2605 GND.n2287 19.3944
R19811 GND.n2611 GND.n2287 19.3944
R19812 GND.n2611 GND.n2610 19.3944
R19813 GND.n2610 GND.n2267 19.3944
R19814 GND.n2638 GND.n2267 19.3944
R19815 GND.n2638 GND.n2265 19.3944
R19816 GND.n2642 GND.n2265 19.3944
R19817 GND.n2642 GND.n2248 19.3944
R19818 GND.n2705 GND.n2248 19.3944
R19819 GND.n2705 GND.n2246 19.3944
R19820 GND.n2711 GND.n2246 19.3944
R19821 GND.n2711 GND.n2710 19.3944
R19822 GND.n2710 GND.n2225 19.3944
R19823 GND.n2730 GND.n2225 19.3944
R19824 GND.n2730 GND.n2223 19.3944
R19825 GND.n2736 GND.n2223 19.3944
R19826 GND.n2736 GND.n2735 19.3944
R19827 GND.n2735 GND.n2202 19.3944
R19828 GND.n2754 GND.n2202 19.3944
R19829 GND.n2754 GND.n2200 19.3944
R19830 GND.n2758 GND.n2200 19.3944
R19831 GND.n2758 GND.n2113 19.3944
R19832 GND.n2822 GND.n2113 19.3944
R19833 GND.n2112 GND.n2111 19.3944
R19834 GND.n2138 GND.n2111 19.3944
R19835 GND.n2806 GND.n2805 19.3944
R19836 GND.n2784 GND.n2783 19.3944
R19837 GND.n2786 GND.n2105 19.3944
R19838 GND.n2828 GND.n2105 19.3944
R19839 GND.n2828 GND.n2827 19.3944
R19840 GND.n2827 GND.n2084 19.3944
R19841 GND.n2847 GND.n2084 19.3944
R19842 GND.n2847 GND.n2082 19.3944
R19843 GND.n2853 GND.n2082 19.3944
R19844 GND.n2853 GND.n2852 19.3944
R19845 GND.n2852 GND.n2062 19.3944
R19846 GND.n2872 GND.n2062 19.3944
R19847 GND.n2872 GND.n2060 19.3944
R19848 GND.n2878 GND.n2060 19.3944
R19849 GND.n2878 GND.n2877 19.3944
R19850 GND.n2877 GND.n2034 19.3944
R19851 GND.n7670 GND.n2034 19.3944
R19852 GND.n7670 GND.n2032 19.3944
R19853 GND.n7676 GND.n2032 19.3944
R19854 GND.n7676 GND.n7675 19.3944
R19855 GND.n7675 GND.n2011 19.3944
R19856 GND.n7694 GND.n2011 19.3944
R19857 GND.n7694 GND.n2009 19.3944
R19858 GND.n7700 GND.n2009 19.3944
R19859 GND.n7700 GND.n7699 19.3944
R19860 GND.n7699 GND.n1988 19.3944
R19861 GND.n7719 GND.n1988 19.3944
R19862 GND.n7719 GND.n1986 19.3944
R19863 GND.n7725 GND.n1986 19.3944
R19864 GND.n7725 GND.n7724 19.3944
R19865 GND.n7724 GND.n1966 19.3944
R19866 GND.n7744 GND.n1966 19.3944
R19867 GND.n7744 GND.n1964 19.3944
R19868 GND.n7750 GND.n1964 19.3944
R19869 GND.n7750 GND.n7749 19.3944
R19870 GND.n7749 GND.n1943 19.3944
R19871 GND.n7769 GND.n1943 19.3944
R19872 GND.n7769 GND.n1941 19.3944
R19873 GND.n7775 GND.n1941 19.3944
R19874 GND.n7775 GND.n7774 19.3944
R19875 GND.n7774 GND.n1920 19.3944
R19876 GND.n7793 GND.n1920 19.3944
R19877 GND.n7793 GND.n1918 19.3944
R19878 GND.n7799 GND.n1918 19.3944
R19879 GND.n7799 GND.n7798 19.3944
R19880 GND.n7798 GND.n1898 19.3944
R19881 GND.n7820 GND.n1898 19.3944
R19882 GND.n7820 GND.n1896 19.3944
R19883 GND.n7824 GND.n1896 19.3944
R19884 GND.n7824 GND.n1777 19.3944
R19885 GND.n7922 GND.n1777 19.3944
R19886 GND.n8173 GND.n8172 19.3944
R19887 GND.n8172 GND.n8171 19.3944
R19888 GND.n8171 GND.n1433 19.3944
R19889 GND.n8165 GND.n1433 19.3944
R19890 GND.n8165 GND.n8164 19.3944
R19891 GND.n8164 GND.n8163 19.3944
R19892 GND.n8163 GND.n1442 19.3944
R19893 GND.n8157 GND.n1442 19.3944
R19894 GND.n8157 GND.n8156 19.3944
R19895 GND.n8156 GND.n8155 19.3944
R19896 GND.n8155 GND.n1450 19.3944
R19897 GND.n1518 GND.n1450 19.3944
R19898 GND.n1518 GND.n1515 19.3944
R19899 GND.n8091 GND.n1515 19.3944
R19900 GND.n8091 GND.n8090 19.3944
R19901 GND.n8090 GND.n8089 19.3944
R19902 GND.n8089 GND.n1524 19.3944
R19903 GND.n2429 GND.n1524 19.3944
R19904 GND.n2432 GND.n2429 19.3944
R19905 GND.n2432 GND.n2426 19.3944
R19906 GND.n2501 GND.n2426 19.3944
R19907 GND.n2501 GND.n2500 19.3944
R19908 GND.n2500 GND.n2499 19.3944
R19909 GND.n2499 GND.n2438 19.3944
R19910 GND.n2495 GND.n2438 19.3944
R19911 GND.n2495 GND.n2494 19.3944
R19912 GND.n2494 GND.n2493 19.3944
R19913 GND.n2493 GND.n2444 19.3944
R19914 GND.n2489 GND.n2444 19.3944
R19915 GND.n2489 GND.n2488 19.3944
R19916 GND.n2488 GND.n2487 19.3944
R19917 GND.n2487 GND.n2450 19.3944
R19918 GND.n2483 GND.n2450 19.3944
R19919 GND.n2483 GND.n2482 19.3944
R19920 GND.n2482 GND.n2481 19.3944
R19921 GND.n2481 GND.n2456 19.3944
R19922 GND.n2477 GND.n2456 19.3944
R19923 GND.n2477 GND.n2476 19.3944
R19924 GND.n2476 GND.n2475 19.3944
R19925 GND.n2475 GND.n2462 19.3944
R19926 GND.n2471 GND.n2462 19.3944
R19927 GND.n2471 GND.n2470 19.3944
R19928 GND.n2470 GND.n2469 19.3944
R19929 GND.n2469 GND.n2259 19.3944
R19930 GND.n2647 GND.n2259 19.3944
R19931 GND.n2647 GND.n2257 19.3944
R19932 GND.n2694 GND.n2257 19.3944
R19933 GND.n2694 GND.n2693 19.3944
R19934 GND.n2693 GND.n2692 19.3944
R19935 GND.n2692 GND.n2653 19.3944
R19936 GND.n2688 GND.n2653 19.3944
R19937 GND.n2688 GND.n2687 19.3944
R19938 GND.n2687 GND.n2686 19.3944
R19939 GND.n2686 GND.n2659 19.3944
R19940 GND.n2682 GND.n2659 19.3944
R19941 GND.n2682 GND.n2681 19.3944
R19942 GND.n2681 GND.n2680 19.3944
R19943 GND.n2680 GND.n2665 19.3944
R19944 GND.n2676 GND.n2665 19.3944
R19945 GND.n2676 GND.n2675 19.3944
R19946 GND.n2675 GND.n2674 19.3944
R19947 GND.n2814 GND.n2127 19.3944
R19948 GND.n2814 GND.n2813 19.3944
R19949 GND.n2811 GND.n2128 19.3944
R19950 GND.n2797 GND.n2150 19.3944
R19951 GND.n2795 GND.n2794 19.3944
R19952 GND.n2182 GND.n2181 19.3944
R19953 GND.n2181 GND.n2180 19.3944
R19954 GND.n2180 GND.n2155 19.3944
R19955 GND.n2176 GND.n2155 19.3944
R19956 GND.n2176 GND.n2175 19.3944
R19957 GND.n2175 GND.n2174 19.3944
R19958 GND.n2174 GND.n2161 19.3944
R19959 GND.n2170 GND.n2161 19.3944
R19960 GND.n2170 GND.n2169 19.3944
R19961 GND.n2169 GND.n2168 19.3944
R19962 GND.n2168 GND.n2044 19.3944
R19963 GND.n2892 GND.n2044 19.3944
R19964 GND.n2892 GND.n2042 19.3944
R19965 GND.n7661 GND.n2042 19.3944
R19966 GND.n7661 GND.n7660 19.3944
R19967 GND.n7660 GND.n7659 19.3944
R19968 GND.n7659 GND.n2898 19.3944
R19969 GND.n7655 GND.n2898 19.3944
R19970 GND.n7655 GND.n7654 19.3944
R19971 GND.n7654 GND.n7653 19.3944
R19972 GND.n7653 GND.n2904 19.3944
R19973 GND.n7649 GND.n2904 19.3944
R19974 GND.n7649 GND.n7648 19.3944
R19975 GND.n7648 GND.n7647 19.3944
R19976 GND.n7647 GND.n2910 19.3944
R19977 GND.n7643 GND.n2910 19.3944
R19978 GND.n7643 GND.n7642 19.3944
R19979 GND.n7642 GND.n7641 19.3944
R19980 GND.n7641 GND.n2916 19.3944
R19981 GND.n7637 GND.n2916 19.3944
R19982 GND.n7637 GND.n7636 19.3944
R19983 GND.n7636 GND.n7635 19.3944
R19984 GND.n7635 GND.n2922 19.3944
R19985 GND.n7631 GND.n2922 19.3944
R19986 GND.n7631 GND.n7630 19.3944
R19987 GND.n7630 GND.n7629 19.3944
R19988 GND.n7629 GND.n2928 19.3944
R19989 GND.n7625 GND.n2928 19.3944
R19990 GND.n7625 GND.n7624 19.3944
R19991 GND.n7624 GND.n7623 19.3944
R19992 GND.n7623 GND.n2934 19.3944
R19993 GND.n7619 GND.n2934 19.3944
R19994 GND.n7619 GND.n7618 19.3944
R19995 GND.n7618 GND.n7617 19.3944
R19996 GND.n7617 GND.n2940 19.3944
R19997 GND.n7613 GND.n2940 19.3944
R19998 GND.n7613 GND.n7612 19.3944
R19999 GND.n7612 GND.n7611 19.3944
R20000 GND.n7611 GND.n2946 19.3944
R20001 GND.n7607 GND.n2946 19.3944
R20002 GND.n7607 GND.n7606 19.3944
R20003 GND.n7606 GND.n7605 19.3944
R20004 GND.n7605 GND.n2952 19.3944
R20005 GND.n7599 GND.n2952 19.3944
R20006 GND.n7599 GND.n7598 19.3944
R20007 GND.n7598 GND.n7597 19.3944
R20008 GND.n7597 GND.n2961 19.3944
R20009 GND.n7585 GND.n2961 19.3944
R20010 GND.n7585 GND.n7584 19.3944
R20011 GND.n7584 GND.n7583 19.3944
R20012 GND.n7583 GND.n2979 19.3944
R20013 GND.n7571 GND.n2979 19.3944
R20014 GND.n7571 GND.n7570 19.3944
R20015 GND.n7570 GND.n7569 19.3944
R20016 GND.n7569 GND.n2998 19.3944
R20017 GND.n7557 GND.n2998 19.3944
R20018 GND.n7557 GND.n7556 19.3944
R20019 GND.n7556 GND.n7555 19.3944
R20020 GND.n7555 GND.n3019 19.3944
R20021 GND.n4892 GND.n3019 19.3944
R20022 GND.n4904 GND.n4892 19.3944
R20023 GND.n4904 GND.n4903 19.3944
R20024 GND.n4903 GND.n4902 19.3944
R20025 GND.n4902 GND.n4899 19.3944
R20026 GND.n4899 GND.n4625 19.3944
R20027 GND.n4938 GND.n4625 19.3944
R20028 GND.n4938 GND.n4623 19.3944
R20029 GND.n4944 GND.n4623 19.3944
R20030 GND.n4944 GND.n4943 19.3944
R20031 GND.n4943 GND.n4596 19.3944
R20032 GND.n4992 GND.n4596 19.3944
R20033 GND.n4992 GND.n4594 19.3944
R20034 GND.n4998 GND.n4594 19.3944
R20035 GND.n4998 GND.n4997 19.3944
R20036 GND.n4997 GND.n4573 19.3944
R20037 GND.n5052 GND.n4573 19.3944
R20038 GND.n5052 GND.n4571 19.3944
R20039 GND.n5067 GND.n4571 19.3944
R20040 GND.n5067 GND.n5066 19.3944
R20041 GND.n5066 GND.n5065 19.3944
R20042 GND.n5065 GND.n5058 19.3944
R20043 GND.n5061 GND.n5058 19.3944
R20044 GND.n5061 GND.n4534 19.3944
R20045 GND.n5110 GND.n4534 19.3944
R20046 GND.n5110 GND.n4532 19.3944
R20047 GND.n5114 GND.n4532 19.3944
R20048 GND.n5114 GND.n4508 19.3944
R20049 GND.n5155 GND.n4508 19.3944
R20050 GND.n5155 GND.n4506 19.3944
R20051 GND.n5161 GND.n4506 19.3944
R20052 GND.n5161 GND.n5160 19.3944
R20053 GND.n5160 GND.n4488 19.3944
R20054 GND.n5215 GND.n4488 19.3944
R20055 GND.n5215 GND.n4486 19.3944
R20056 GND.n5227 GND.n4486 19.3944
R20057 GND.n5227 GND.n5226 19.3944
R20058 GND.n5226 GND.n5225 19.3944
R20059 GND.n5225 GND.n5222 19.3944
R20060 GND.n5222 GND.n4453 19.3944
R20061 GND.n5261 GND.n4453 19.3944
R20062 GND.n5261 GND.n4451 19.3944
R20063 GND.n5267 GND.n4451 19.3944
R20064 GND.n5267 GND.n5266 19.3944
R20065 GND.n5266 GND.n4425 19.3944
R20066 GND.n5316 GND.n4425 19.3944
R20067 GND.n5316 GND.n4423 19.3944
R20068 GND.n5322 GND.n4423 19.3944
R20069 GND.n5322 GND.n5321 19.3944
R20070 GND.n5321 GND.n4402 19.3944
R20071 GND.n5377 GND.n4402 19.3944
R20072 GND.n5377 GND.n4400 19.3944
R20073 GND.n5389 GND.n4400 19.3944
R20074 GND.n5389 GND.n5388 19.3944
R20075 GND.n5388 GND.n5387 19.3944
R20076 GND.n5387 GND.n5384 19.3944
R20077 GND.n5384 GND.n4367 19.3944
R20078 GND.n5423 GND.n4367 19.3944
R20079 GND.n5423 GND.n4365 19.3944
R20080 GND.n5429 GND.n4365 19.3944
R20081 GND.n5429 GND.n5428 19.3944
R20082 GND.n5428 GND.n4338 19.3944
R20083 GND.n5476 GND.n4338 19.3944
R20084 GND.n5476 GND.n4336 19.3944
R20085 GND.n5482 GND.n4336 19.3944
R20086 GND.n5482 GND.n5481 19.3944
R20087 GND.n5481 GND.n4315 19.3944
R20088 GND.n5548 GND.n4315 19.3944
R20089 GND.n5548 GND.n4313 19.3944
R20090 GND.n5560 GND.n4313 19.3944
R20091 GND.n5560 GND.n5559 19.3944
R20092 GND.n5559 GND.n5558 19.3944
R20093 GND.n5558 GND.n5555 19.3944
R20094 GND.n5555 GND.n4282 19.3944
R20095 GND.n5594 GND.n4282 19.3944
R20096 GND.n5594 GND.n4280 19.3944
R20097 GND.n5600 GND.n4280 19.3944
R20098 GND.n5600 GND.n5599 19.3944
R20099 GND.n5599 GND.n4254 19.3944
R20100 GND.n5632 GND.n4254 19.3944
R20101 GND.n5632 GND.n4252 19.3944
R20102 GND.n5636 GND.n4252 19.3944
R20103 GND.n5636 GND.n4230 19.3944
R20104 GND.n5688 GND.n4230 19.3944
R20105 GND.n5688 GND.n4228 19.3944
R20106 GND.n5694 GND.n4228 19.3944
R20107 GND.n5694 GND.n5693 19.3944
R20108 GND.n5693 GND.n4207 19.3944
R20109 GND.n5722 GND.n4207 19.3944
R20110 GND.n5722 GND.n4205 19.3944
R20111 GND.n5728 GND.n4205 19.3944
R20112 GND.n5728 GND.n5727 19.3944
R20113 GND.n5727 GND.n4184 19.3944
R20114 GND.n5803 GND.n4184 19.3944
R20115 GND.n5803 GND.n4182 19.3944
R20116 GND.n5818 GND.n4182 19.3944
R20117 GND.n5818 GND.n5817 19.3944
R20118 GND.n5817 GND.n5816 19.3944
R20119 GND.n5816 GND.n5809 19.3944
R20120 GND.n5812 GND.n5809 19.3944
R20121 GND.n5812 GND.n4147 19.3944
R20122 GND.n5863 GND.n4147 19.3944
R20123 GND.n5863 GND.n4145 19.3944
R20124 GND.n5875 GND.n4145 19.3944
R20125 GND.n5875 GND.n5874 19.3944
R20126 GND.n5874 GND.n5873 19.3944
R20127 GND.n5873 GND.n5870 19.3944
R20128 GND.n5870 GND.n4112 19.3944
R20129 GND.n5909 GND.n4112 19.3944
R20130 GND.n5909 GND.n4110 19.3944
R20131 GND.n5915 GND.n4110 19.3944
R20132 GND.n5915 GND.n5914 19.3944
R20133 GND.n5914 GND.n4083 19.3944
R20134 GND.n5962 GND.n4083 19.3944
R20135 GND.n5962 GND.n4081 19.3944
R20136 GND.n5968 GND.n4081 19.3944
R20137 GND.n5968 GND.n5967 19.3944
R20138 GND.n5967 GND.n4059 19.3944
R20139 GND.n6011 GND.n4059 19.3944
R20140 GND.n6011 GND.n4057 19.3944
R20141 GND.n6026 GND.n4057 19.3944
R20142 GND.n6026 GND.n6025 19.3944
R20143 GND.n6025 GND.n6024 19.3944
R20144 GND.n6024 GND.n6017 19.3944
R20145 GND.n6020 GND.n6017 19.3944
R20146 GND.n6020 GND.n4018 19.3944
R20147 GND.n6087 GND.n4018 19.3944
R20148 GND.n6087 GND.n4016 19.3944
R20149 GND.n6093 GND.n4016 19.3944
R20150 GND.n6093 GND.n6092 19.3944
R20151 GND.n6092 GND.n3996 19.3944
R20152 GND.n6352 GND.n3996 19.3944
R20153 GND.n6352 GND.n3994 19.3944
R20154 GND.n6359 GND.n3994 19.3944
R20155 GND.n6359 GND.n6358 19.3944
R20156 GND.n6358 GND.n3235 19.3944
R20157 GND.n7339 GND.n3235 19.3944
R20158 GND.n7339 GND.n7338 19.3944
R20159 GND.n7338 GND.n7337 19.3944
R20160 GND.n7337 GND.n3239 19.3944
R20161 GND.n7325 GND.n3239 19.3944
R20162 GND.n7325 GND.n7324 19.3944
R20163 GND.n7324 GND.n7323 19.3944
R20164 GND.n7323 GND.n3256 19.3944
R20165 GND.n3276 GND.n3256 19.3944
R20166 GND.n7306 GND.n3276 19.3944
R20167 GND.n7306 GND.n7305 19.3944
R20168 GND.n7305 GND.n7304 19.3944
R20169 GND.n7304 GND.n3282 19.3944
R20170 GND.n7298 GND.n3282 19.3944
R20171 GND.n7298 GND.n7297 19.3944
R20172 GND.n7297 GND.n7296 19.3944
R20173 GND.n7296 GND.n3290 19.3944
R20174 GND.n6445 GND.n3290 19.3944
R20175 GND.n6445 GND.n6442 19.3944
R20176 GND.n6449 GND.n6442 19.3944
R20177 GND.n6449 GND.n6440 19.3944
R20178 GND.n6578 GND.n6440 19.3944
R20179 GND.n6578 GND.n6577 19.3944
R20180 GND.n6577 GND.n6576 19.3944
R20181 GND.n6576 GND.n6455 19.3944
R20182 GND.n6572 GND.n6455 19.3944
R20183 GND.n6572 GND.n6571 19.3944
R20184 GND.n6571 GND.n6570 19.3944
R20185 GND.n6570 GND.n6461 19.3944
R20186 GND.n6566 GND.n6461 19.3944
R20187 GND.n6566 GND.n6565 19.3944
R20188 GND.n6565 GND.n6564 19.3944
R20189 GND.n6564 GND.n6467 19.3944
R20190 GND.n6560 GND.n6467 19.3944
R20191 GND.n6560 GND.n6559 19.3944
R20192 GND.n6559 GND.n6558 19.3944
R20193 GND.n6558 GND.n6473 19.3944
R20194 GND.n6554 GND.n6473 19.3944
R20195 GND.n6554 GND.n6553 19.3944
R20196 GND.n6553 GND.n6552 19.3944
R20197 GND.n6552 GND.n6479 19.3944
R20198 GND.n6548 GND.n6479 19.3944
R20199 GND.n6548 GND.n6547 19.3944
R20200 GND.n6547 GND.n6546 19.3944
R20201 GND.n6546 GND.n6485 19.3944
R20202 GND.n6542 GND.n6485 19.3944
R20203 GND.n6542 GND.n6541 19.3944
R20204 GND.n6541 GND.n6540 19.3944
R20205 GND.n6540 GND.n6491 19.3944
R20206 GND.n6536 GND.n6491 19.3944
R20207 GND.n6536 GND.n6535 19.3944
R20208 GND.n6535 GND.n6534 19.3944
R20209 GND.n6534 GND.n6497 19.3944
R20210 GND.n6530 GND.n6497 19.3944
R20211 GND.n6530 GND.n6529 19.3944
R20212 GND.n6529 GND.n6528 19.3944
R20213 GND.n6528 GND.n6503 19.3944
R20214 GND.n6524 GND.n6503 19.3944
R20215 GND.n6524 GND.n6523 19.3944
R20216 GND.n6523 GND.n6522 19.3944
R20217 GND.n6522 GND.n6509 19.3944
R20218 GND.n6518 GND.n6509 19.3944
R20219 GND.n6518 GND.n6517 19.3944
R20220 GND.n6517 GND.n6516 19.3944
R20221 GND.n6516 GND.n3746 19.3944
R20222 GND.n6880 GND.n3746 19.3944
R20223 GND.n6880 GND.n3747 19.3944
R20224 GND.n6814 GND.n6813 19.3944
R20225 GND.n6864 GND.n6863 19.3944
R20226 GND.n6842 GND.n6841 19.3944
R20227 GND.n6846 GND.n6845 19.3944
R20228 GND.n6885 GND.n3738 19.3944
R20229 GND.n6885 GND.n6884 19.3944
R20230 GND.n6884 GND.n3718 19.3944
R20231 GND.n6905 GND.n3718 19.3944
R20232 GND.n6905 GND.n3716 19.3944
R20233 GND.n6911 GND.n3716 19.3944
R20234 GND.n6911 GND.n6910 19.3944
R20235 GND.n6910 GND.n3696 19.3944
R20236 GND.n6932 GND.n3696 19.3944
R20237 GND.n6932 GND.n3694 19.3944
R20238 GND.n6938 GND.n3694 19.3944
R20239 GND.n6938 GND.n6937 19.3944
R20240 GND.n6937 GND.n3676 19.3944
R20241 GND.n6961 GND.n3676 19.3944
R20242 GND.n6961 GND.n3674 19.3944
R20243 GND.n6967 GND.n3674 19.3944
R20244 GND.n6967 GND.n6966 19.3944
R20245 GND.n6966 GND.n3654 19.3944
R20246 GND.n6988 GND.n3654 19.3944
R20247 GND.n6988 GND.n3652 19.3944
R20248 GND.n6994 GND.n3652 19.3944
R20249 GND.n6994 GND.n6993 19.3944
R20250 GND.n6993 GND.n3632 19.3944
R20251 GND.n7014 GND.n3632 19.3944
R20252 GND.n7014 GND.n3630 19.3944
R20253 GND.n7020 GND.n3630 19.3944
R20254 GND.n7020 GND.n7019 19.3944
R20255 GND.n7019 GND.n3610 19.3944
R20256 GND.n7041 GND.n3610 19.3944
R20257 GND.n7041 GND.n3608 19.3944
R20258 GND.n7047 GND.n3608 19.3944
R20259 GND.n7047 GND.n7046 19.3944
R20260 GND.n7046 GND.n3589 19.3944
R20261 GND.n7069 GND.n3589 19.3944
R20262 GND.n7069 GND.n3587 19.3944
R20263 GND.n7082 GND.n3587 19.3944
R20264 GND.n7082 GND.n7081 19.3944
R20265 GND.n7081 GND.n7080 19.3944
R20266 GND.n7080 GND.n7077 19.3944
R20267 GND.n7077 GND.n582 19.3944
R20268 GND.n9497 GND.n582 19.3944
R20269 GND.n9497 GND.n9496 19.3944
R20270 GND.n9496 GND.n9495 19.3944
R20271 GND.n9495 GND.n586 19.3944
R20272 GND.n9491 GND.n586 19.3944
R20273 GND.n9491 GND.n9490 19.3944
R20274 GND.n9490 GND.n9489 19.3944
R20275 GND.n9489 GND.n592 19.3944
R20276 GND.n9485 GND.n592 19.3944
R20277 GND.n9485 GND.n9484 19.3944
R20278 GND.n9484 GND.n9483 19.3944
R20279 GND.n9483 GND.n598 19.3944
R20280 GND.n9477 GND.n598 19.3944
R20281 GND.n9477 GND.n9476 19.3944
R20282 GND.n9476 GND.n9475 19.3944
R20283 GND.n9475 GND.n606 19.3944
R20284 GND.n9469 GND.n606 19.3944
R20285 GND.n9469 GND.n9468 19.3944
R20286 GND.n9468 GND.n9467 19.3944
R20287 GND.n9467 GND.n614 19.3944
R20288 GND.n9461 GND.n614 19.3944
R20289 GND.n8286 GND.n1322 19.3944
R20290 GND.n8280 GND.n1322 19.3944
R20291 GND.n8280 GND.n8279 19.3944
R20292 GND.n8279 GND.n8278 19.3944
R20293 GND.n8278 GND.n1329 19.3944
R20294 GND.n8272 GND.n1329 19.3944
R20295 GND.n8272 GND.n8271 19.3944
R20296 GND.n8271 GND.n8270 19.3944
R20297 GND.n8270 GND.n1337 19.3944
R20298 GND.n8264 GND.n1337 19.3944
R20299 GND.n8264 GND.n8263 19.3944
R20300 GND.n8263 GND.n8262 19.3944
R20301 GND.n8262 GND.n1345 19.3944
R20302 GND.n8256 GND.n1345 19.3944
R20303 GND.n8256 GND.n8255 19.3944
R20304 GND.n8255 GND.n8254 19.3944
R20305 GND.n8254 GND.n1353 19.3944
R20306 GND.n8248 GND.n1353 19.3944
R20307 GND.n8248 GND.n8247 19.3944
R20308 GND.n8247 GND.n8246 19.3944
R20309 GND.n8246 GND.n1361 19.3944
R20310 GND.n8240 GND.n1361 19.3944
R20311 GND.n8240 GND.n8239 19.3944
R20312 GND.n8239 GND.n8238 19.3944
R20313 GND.n8238 GND.n1369 19.3944
R20314 GND.n8232 GND.n1369 19.3944
R20315 GND.n8232 GND.n8231 19.3944
R20316 GND.n8231 GND.n8230 19.3944
R20317 GND.n8230 GND.n1377 19.3944
R20318 GND.n8224 GND.n1377 19.3944
R20319 GND.n8224 GND.n8223 19.3944
R20320 GND.n8223 GND.n8222 19.3944
R20321 GND.n8222 GND.n1385 19.3944
R20322 GND.n8216 GND.n1385 19.3944
R20323 GND.n8216 GND.n8215 19.3944
R20324 GND.n8215 GND.n8214 19.3944
R20325 GND.n8214 GND.n1393 19.3944
R20326 GND.n8208 GND.n1393 19.3944
R20327 GND.n8208 GND.n8207 19.3944
R20328 GND.n8207 GND.n8206 19.3944
R20329 GND.n8206 GND.n1401 19.3944
R20330 GND.n8200 GND.n1401 19.3944
R20331 GND.n8200 GND.n8199 19.3944
R20332 GND.n8199 GND.n8198 19.3944
R20333 GND.n8198 GND.n1409 19.3944
R20334 GND.n8192 GND.n1409 19.3944
R20335 GND.n8192 GND.n8191 19.3944
R20336 GND.n8191 GND.n8190 19.3944
R20337 GND.n8190 GND.n1417 19.3944
R20338 GND.n8184 GND.n1417 19.3944
R20339 GND.n8184 GND.n8183 19.3944
R20340 GND.n8183 GND.n8182 19.3944
R20341 GND.n8182 GND.n1425 19.3944
R20342 GND.n8176 GND.n1425 19.3944
R20343 GND.n7291 GND.n7290 19.3944
R20344 GND.n7290 GND.n3316 19.3944
R20345 GND.n7283 GND.n3316 19.3944
R20346 GND.n7283 GND.n7282 19.3944
R20347 GND.n7282 GND.n3328 19.3944
R20348 GND.n7275 GND.n3328 19.3944
R20349 GND.n7275 GND.n7274 19.3944
R20350 GND.n7274 GND.n3336 19.3944
R20351 GND.n7267 GND.n3336 19.3944
R20352 GND.n7267 GND.n7266 19.3944
R20353 GND.n6431 GND.n3355 19.3944
R20354 GND.n6431 GND.n3962 19.3944
R20355 GND.n6435 GND.n3962 19.3944
R20356 GND.n6435 GND.n3956 19.3944
R20357 GND.n6596 GND.n3956 19.3944
R20358 GND.n6596 GND.n3953 19.3944
R20359 GND.n6601 GND.n3953 19.3944
R20360 GND.n6601 GND.n3954 19.3944
R20361 GND.n3954 GND.n3935 19.3944
R20362 GND.n6621 GND.n3935 19.3944
R20363 GND.n6621 GND.n3932 19.3944
R20364 GND.n6626 GND.n3932 19.3944
R20365 GND.n6626 GND.n3933 19.3944
R20366 GND.n3933 GND.n3911 19.3944
R20367 GND.n6645 GND.n3911 19.3944
R20368 GND.n6645 GND.n3908 19.3944
R20369 GND.n6650 GND.n3908 19.3944
R20370 GND.n6650 GND.n3909 19.3944
R20371 GND.n3909 GND.n3888 19.3944
R20372 GND.n6670 GND.n3888 19.3944
R20373 GND.n6670 GND.n3885 19.3944
R20374 GND.n6675 GND.n3885 19.3944
R20375 GND.n6675 GND.n3886 19.3944
R20376 GND.n3886 GND.n3866 19.3944
R20377 GND.n6695 GND.n3866 19.3944
R20378 GND.n6695 GND.n3863 19.3944
R20379 GND.n6700 GND.n3863 19.3944
R20380 GND.n6700 GND.n3864 19.3944
R20381 GND.n3864 GND.n3844 19.3944
R20382 GND.n6720 GND.n3844 19.3944
R20383 GND.n6720 GND.n3841 19.3944
R20384 GND.n6725 GND.n3841 19.3944
R20385 GND.n6725 GND.n3842 19.3944
R20386 GND.n3842 GND.n3820 19.3944
R20387 GND.n6744 GND.n3820 19.3944
R20388 GND.n6744 GND.n3817 19.3944
R20389 GND.n6749 GND.n3817 19.3944
R20390 GND.n6749 GND.n3818 19.3944
R20391 GND.n3818 GND.n3797 19.3944
R20392 GND.n6769 GND.n3797 19.3944
R20393 GND.n6769 GND.n3794 19.3944
R20394 GND.n6774 GND.n3794 19.3944
R20395 GND.n6774 GND.n3795 19.3944
R20396 GND.n3795 GND.n3770 19.3944
R20397 GND.n6795 GND.n3770 19.3944
R20398 GND.n6795 GND.n3767 19.3944
R20399 GND.n6799 GND.n3767 19.3944
R20400 GND.n6800 GND.n6799 19.3944
R20401 GND.n6804 GND.n6800 19.3944
R20402 GND.n6804 GND.n3765 19.3944
R20403 GND.n6808 GND.n3765 19.3944
R20404 GND.n6808 GND.n408 19.3944
R20405 GND.n9692 GND.n408 19.3944
R20406 GND.n9692 GND.n9691 19.3944
R20407 GND.n9691 GND.n9690 19.3944
R20408 GND.n9690 GND.n412 19.3944
R20409 GND.n9686 GND.n412 19.3944
R20410 GND.n9686 GND.n9685 19.3944
R20411 GND.n9685 GND.n9684 19.3944
R20412 GND.n9684 GND.n417 19.3944
R20413 GND.n9680 GND.n417 19.3944
R20414 GND.n9680 GND.n9679 19.3944
R20415 GND.n9679 GND.n9678 19.3944
R20416 GND.n9678 GND.n422 19.3944
R20417 GND.n9674 GND.n422 19.3944
R20418 GND.n9674 GND.n9673 19.3944
R20419 GND.n9673 GND.n9672 19.3944
R20420 GND.n9672 GND.n427 19.3944
R20421 GND.n9668 GND.n427 19.3944
R20422 GND.n9668 GND.n9667 19.3944
R20423 GND.n9667 GND.n9666 19.3944
R20424 GND.n9666 GND.n432 19.3944
R20425 GND.n9662 GND.n432 19.3944
R20426 GND.n9662 GND.n9661 19.3944
R20427 GND.n9661 GND.n9660 19.3944
R20428 GND.n9660 GND.n437 19.3944
R20429 GND.n9656 GND.n437 19.3944
R20430 GND.n9656 GND.n9655 19.3944
R20431 GND.n9655 GND.n9654 19.3944
R20432 GND.n9654 GND.n442 19.3944
R20433 GND.n9650 GND.n442 19.3944
R20434 GND.n9650 GND.n9649 19.3944
R20435 GND.n9649 GND.n9648 19.3944
R20436 GND.n9648 GND.n447 19.3944
R20437 GND.n9644 GND.n447 19.3944
R20438 GND.n9644 GND.n9643 19.3944
R20439 GND.n9643 GND.n9642 19.3944
R20440 GND.n9642 GND.n452 19.3944
R20441 GND.n9638 GND.n452 19.3944
R20442 GND.n9638 GND.n9637 19.3944
R20443 GND.n9637 GND.n9636 19.3944
R20444 GND.n9636 GND.n457 19.3944
R20445 GND.n9632 GND.n457 19.3944
R20446 GND.n9632 GND.n9631 19.3944
R20447 GND.n9631 GND.n9630 19.3944
R20448 GND.n9630 GND.n462 19.3944
R20449 GND.n9626 GND.n462 19.3944
R20450 GND.n9626 GND.n9625 19.3944
R20451 GND.n9625 GND.n9624 19.3944
R20452 GND.n9624 GND.n467 19.3944
R20453 GND.n9620 GND.n467 19.3944
R20454 GND.n9620 GND.n9619 19.3944
R20455 GND.n9619 GND.n9618 19.3944
R20456 GND.n9618 GND.n472 19.3944
R20457 GND.n9614 GND.n472 19.3944
R20458 GND.n8094 GND.n1509 19.1543
R20459 GND.n8094 GND.n8093 19.1543
R20460 GND.n8093 GND.n1512 19.1543
R20461 GND.n1526 GND.n1512 19.1543
R20462 GND.n1527 GND.n1526 19.1543
R20463 GND.n8087 GND.n1527 19.1543
R20464 GND.n8087 GND.n8086 19.1543
R20465 GND.n8086 GND.n1530 19.1543
R20466 GND.n2370 GND.n1530 19.1543
R20467 GND.n2370 GND.n1546 19.1543
R20468 GND.n8080 GND.n1546 19.1543
R20469 GND.n8080 GND.n1549 19.1543
R20470 GND.n2423 GND.n1549 19.1543
R20471 GND.t101 GND.n2423 19.1543
R20472 GND.n2514 GND.t101 19.1543
R20473 GND.n2514 GND.n2503 19.1543
R20474 GND.n2506 GND.n2503 19.1543
R20475 GND.n2506 GND.n2364 19.1543
R20476 GND.n2523 GND.n2364 19.1543
R20477 GND.n2523 GND.n2360 19.1543
R20478 GND.n2529 GND.n2360 19.1543
R20479 GND.n2529 GND.n2362 19.1543
R20480 GND.n2525 GND.n2362 19.1543
R20481 GND.n2525 GND.n2349 19.1543
R20482 GND.n2539 GND.n2349 19.1543
R20483 GND.n2539 GND.n2351 19.1543
R20484 GND.n2354 GND.n2351 19.1543
R20485 GND.n2354 GND.n2342 19.1543
R20486 GND.n2548 GND.n2342 19.1543
R20487 GND.n2548 GND.n2337 19.1543
R20488 GND.n2554 GND.n2337 19.1543
R20489 GND.n2554 GND.n2339 19.1543
R20490 GND.n2551 GND.n2339 19.1543
R20491 GND.n2551 GND.n2327 19.1543
R20492 GND.n2564 GND.n2327 19.1543
R20493 GND.n2564 GND.n2328 19.1543
R20494 GND.n2331 GND.n2328 19.1543
R20495 GND.n2331 GND.n2320 19.1543
R20496 GND.n2573 GND.n2320 19.1543
R20497 GND.n2573 GND.n2314 19.1543
R20498 GND.n2578 GND.n2314 19.1543
R20499 GND.n2578 GND.n2317 19.1543
R20500 GND.n2575 GND.n2317 19.1543
R20501 GND.n2588 GND.n2303 19.1543
R20502 GND.n2588 GND.n2304 19.1543
R20503 GND.n2308 GND.n2304 19.1543
R20504 GND.n2308 GND.n2295 19.1543
R20505 GND.n2597 GND.n2295 19.1543
R20506 GND.n2597 GND.n2291 19.1543
R20507 GND.n2603 GND.n2291 19.1543
R20508 GND.n2603 GND.n2293 19.1543
R20509 GND.n2600 GND.n2293 19.1543
R20510 GND.n2600 GND.n2280 19.1543
R20511 GND.n2613 GND.n2280 19.1543
R20512 GND.n2613 GND.n2281 19.1543
R20513 GND.n2285 GND.n2281 19.1543
R20514 GND.n2285 GND.n2273 19.1543
R20515 GND.n2631 GND.n2273 19.1543
R20516 GND.n2631 GND.n2269 19.1543
R20517 GND.n2636 GND.n2269 19.1543
R20518 GND.n2636 GND.n2271 19.1543
R20519 GND.n2271 GND.n2261 19.1543
R20520 GND.n2645 GND.n2261 19.1543
R20521 GND.n2645 GND.n2644 19.1543
R20522 GND.n2644 GND.n2253 19.1543
R20523 GND.n2697 GND.n2253 19.1543
R20524 GND.n2697 GND.n2696 19.1543
R20525 GND.n2703 GND.n2251 19.1543
R20526 GND.n2699 GND.n2251 19.1543
R20527 GND.n2699 GND.n2239 19.1543
R20528 GND.n2713 GND.n2239 19.1543
R20529 GND.n2713 GND.n2241 19.1543
R20530 GND.n2244 GND.n2241 19.1543
R20531 GND.n2244 GND.n2232 19.1543
R20532 GND.n2722 GND.n2232 19.1543
R20533 GND.n2722 GND.n2227 19.1543
R20534 GND.n2728 GND.n2227 19.1543
R20535 GND.n2728 GND.n2229 19.1543
R20536 GND.n2725 GND.n2229 19.1543
R20537 GND.n2725 GND.n2217 19.1543
R20538 GND.n2738 GND.n2217 19.1543
R20539 GND.n2738 GND.n2218 19.1543
R20540 GND.n2221 GND.n2218 19.1543
R20541 GND.n2221 GND.n2210 19.1543
R20542 GND.n2747 GND.n2210 19.1543
R20543 GND.n2747 GND.n2204 19.1543
R20544 GND.n2752 GND.n2204 19.1543
R20545 GND.n2752 GND.n2207 19.1543
R20546 GND.n2749 GND.n2207 19.1543
R20547 GND.n2749 GND.n2196 19.1543
R20548 GND.n2760 GND.n2196 19.1543
R20549 GND.n2667 GND.n2666 19.1543
R20550 GND.n2666 GND.n2116 19.1543
R20551 GND.n2820 GND.n2116 19.1543
R20552 GND.n2820 GND.n2119 19.1543
R20553 GND.n2817 GND.n2119 19.1543
R20554 GND.n2817 GND.n2816 19.1543
R20555 GND.n2816 GND.n2124 19.1543
R20556 GND.n2130 GND.n2124 19.1543
R20557 GND.n2131 GND.n2130 19.1543
R20558 GND.n2809 GND.n2131 19.1543
R20559 GND.n2809 GND.n2808 19.1543
R20560 GND.n2808 GND.n2134 19.1543
R20561 GND.n2803 GND.n2134 19.1543
R20562 GND.n2803 GND.n2142 19.1543
R20563 GND.n2800 GND.n2142 19.1543
R20564 GND.n2800 GND.n2799 19.1543
R20565 GND.n2799 GND.n2146 19.1543
R20566 GND.n2184 GND.n2146 19.1543
R20567 GND.n2788 GND.n2184 19.1543
R20568 GND.n2792 GND.n2788 19.1543
R20569 GND.n2792 GND.n2791 19.1543
R20570 GND.n2791 GND.n2098 19.1543
R20571 GND.n2830 GND.n2098 19.1543
R20572 GND.n2830 GND.n2099 19.1543
R20573 GND.n2103 GND.n2090 19.1543
R20574 GND.n2839 GND.n2090 19.1543
R20575 GND.n2839 GND.n2086 19.1543
R20576 GND.n2845 GND.n2086 19.1543
R20577 GND.n2845 GND.n2088 19.1543
R20578 GND.n2842 GND.n2088 19.1543
R20579 GND.n2842 GND.n2075 19.1543
R20580 GND.n2855 GND.n2075 19.1543
R20581 GND.n2855 GND.n2076 19.1543
R20582 GND.n2080 GND.n2076 19.1543
R20583 GND.n2080 GND.n2068 19.1543
R20584 GND.n2864 GND.n2068 19.1543
R20585 GND.n2864 GND.n2064 19.1543
R20586 GND.n2870 GND.n2064 19.1543
R20587 GND.n2870 GND.n2066 19.1543
R20588 GND.n2866 GND.n2066 19.1543
R20589 GND.n2866 GND.n2053 19.1543
R20590 GND.n2880 GND.n2053 19.1543
R20591 GND.n2880 GND.n2055 19.1543
R20592 GND.n2055 GND.n2046 19.1543
R20593 GND.n2890 GND.n2046 19.1543
R20594 GND.n2890 GND.n2889 19.1543
R20595 GND.n2889 GND.n2036 19.1543
R20596 GND.n7668 GND.n2036 19.1543
R20597 GND.n7665 GND.n7663 19.1543
R20598 GND.n7665 GND.n2026 19.1543
R20599 GND.n7678 GND.n2026 19.1543
R20600 GND.n7678 GND.n2027 19.1543
R20601 GND.n2030 GND.n2027 19.1543
R20602 GND.n2030 GND.n2019 19.1543
R20603 GND.n7687 GND.n2019 19.1543
R20604 GND.n7687 GND.n2013 19.1543
R20605 GND.n7692 GND.n2013 19.1543
R20606 GND.n7692 GND.n2016 19.1543
R20607 GND.n7689 GND.n2016 19.1543
R20608 GND.n7689 GND.n2002 19.1543
R20609 GND.n7702 GND.n2002 19.1543
R20610 GND.n7702 GND.n2003 19.1543
R20611 GND.n2007 GND.n2003 19.1543
R20612 GND.n2007 GND.n1994 19.1543
R20613 GND.n7711 GND.n1994 19.1543
R20614 GND.n7711 GND.n1990 19.1543
R20615 GND.n7717 GND.n1990 19.1543
R20616 GND.n7717 GND.n1992 19.1543
R20617 GND.n7714 GND.n1992 19.1543
R20618 GND.n7714 GND.n1979 19.1543
R20619 GND.n7727 GND.n1979 19.1543
R20620 GND.n7727 GND.n1980 19.1543
R20621 GND.n1984 GND.n1972 19.1543
R20622 GND.n7736 GND.n1972 19.1543
R20623 GND.n7736 GND.n1968 19.1543
R20624 GND.n7742 GND.n1968 19.1543
R20625 GND.n7742 GND.n1970 19.1543
R20626 GND.n7738 GND.n1970 19.1543
R20627 GND.n7738 GND.n1957 19.1543
R20628 GND.n7752 GND.n1957 19.1543
R20629 GND.n7752 GND.n1959 19.1543
R20630 GND.n1962 GND.n1959 19.1543
R20631 GND.n1962 GND.n1950 19.1543
R20632 GND.n7761 GND.n1950 19.1543
R20633 GND.n7761 GND.n1945 19.1543
R20634 GND.n7767 GND.n1945 19.1543
R20635 GND.n7767 GND.n1947 19.1543
R20636 GND.n7764 GND.n1947 19.1543
R20637 GND.n7764 GND.n1935 19.1543
R20638 GND.n7777 GND.n1935 19.1543
R20639 GND.n7777 GND.n1936 19.1543
R20640 GND.n1939 GND.n1936 19.1543
R20641 GND.n1939 GND.n1928 19.1543
R20642 GND.n7786 GND.n1928 19.1543
R20643 GND.n7786 GND.n1922 19.1543
R20644 GND.n7791 GND.n1922 19.1543
R20645 GND.n7791 GND.n1925 19.1543
R20646 GND.n7788 GND.n1925 19.1543
R20647 GND.n7788 GND.n1912 19.1543
R20648 GND.n7801 GND.n1912 19.1543
R20649 GND.n7801 GND.t84 19.1543
R20650 GND.n1916 GND.t84 19.1543
R20651 GND.n1916 GND.n1904 19.1543
R20652 GND.n7815 GND.n1904 19.1543
R20653 GND.n7815 GND.n1900 19.1543
R20654 GND.n7818 GND.n1900 19.1543
R20655 GND.n7818 GND.n1902 19.1543
R20656 GND.n7807 GND.n1902 19.1543
R20657 GND.n7807 GND.n1894 19.1543
R20658 GND.n7826 GND.n1894 19.1543
R20659 GND.n7826 GND.n1891 19.1543
R20660 GND.n7829 GND.n1891 19.1543
R20661 GND.n7829 GND.n1771 19.1543
R20662 GND.n7924 GND.n1771 19.1543
R20663 GND.n7924 GND.n1773 19.1543
R20664 GND.n7256 GND.n3356 19.1543
R20665 GND.n7256 GND.n3358 19.1543
R20666 GND.n3376 GND.n3358 19.1543
R20667 GND.n3376 GND.n3366 19.1543
R20668 GND.n7250 GND.n3366 19.1543
R20669 GND.n7250 GND.n3369 19.1543
R20670 GND.n6437 GND.n3369 19.1543
R20671 GND.n6580 GND.n6437 19.1543
R20672 GND.n6582 GND.n6580 19.1543
R20673 GND.n6582 GND.n3958 19.1543
R20674 GND.n6594 GND.n3958 19.1543
R20675 GND.n6594 GND.n3960 19.1543
R20676 GND.n6584 GND.n3960 19.1543
R20677 GND.n6584 GND.t91 19.1543
R20678 GND.n6603 GND.t91 19.1543
R20679 GND.n6603 GND.n3947 19.1543
R20680 GND.n6609 GND.n3947 19.1543
R20681 GND.n6609 GND.n3949 19.1543
R20682 GND.n6606 GND.n3949 19.1543
R20683 GND.n6606 GND.n3937 19.1543
R20684 GND.n6619 GND.n3937 19.1543
R20685 GND.n6619 GND.n3938 19.1543
R20686 GND.n3941 GND.n3938 19.1543
R20687 GND.n3941 GND.n3930 19.1543
R20688 GND.n6628 GND.n3930 19.1543
R20689 GND.n6628 GND.n3924 19.1543
R20690 GND.n6633 GND.n3924 19.1543
R20691 GND.n6633 GND.n3927 19.1543
R20692 GND.n6630 GND.n3927 19.1543
R20693 GND.n6630 GND.n3913 19.1543
R20694 GND.n6643 GND.n3913 19.1543
R20695 GND.n6643 GND.n3914 19.1543
R20696 GND.n3918 GND.n3914 19.1543
R20697 GND.n3918 GND.n3905 19.1543
R20698 GND.n6652 GND.n3905 19.1543
R20699 GND.n6652 GND.n3901 19.1543
R20700 GND.n6658 GND.n3901 19.1543
R20701 GND.n6658 GND.n3903 19.1543
R20702 GND.n6655 GND.n3903 19.1543
R20703 GND.n6655 GND.n3890 19.1543
R20704 GND.n6668 GND.n3890 19.1543
R20705 GND.n6668 GND.n3891 19.1543
R20706 GND.n3895 GND.n3891 19.1543
R20707 GND.n6677 GND.n3883 19.1543
R20708 GND.n6677 GND.n3879 19.1543
R20709 GND.n6683 GND.n3879 19.1543
R20710 GND.n6683 GND.n3881 19.1543
R20711 GND.n6679 GND.n3881 19.1543
R20712 GND.n6679 GND.n3868 19.1543
R20713 GND.n6693 GND.n3868 19.1543
R20714 GND.n6693 GND.n3870 19.1543
R20715 GND.n3873 GND.n3870 19.1543
R20716 GND.n3873 GND.n3861 19.1543
R20717 GND.n6702 GND.n3861 19.1543
R20718 GND.n6702 GND.n3856 19.1543
R20719 GND.n6708 GND.n3856 19.1543
R20720 GND.n6708 GND.n3858 19.1543
R20721 GND.n6705 GND.n3858 19.1543
R20722 GND.n6705 GND.n3846 19.1543
R20723 GND.n6718 GND.n3846 19.1543
R20724 GND.n6718 GND.n3847 19.1543
R20725 GND.n3850 GND.n3847 19.1543
R20726 GND.n3850 GND.n3839 19.1543
R20727 GND.n6727 GND.n3839 19.1543
R20728 GND.n6727 GND.n3833 19.1543
R20729 GND.n6732 GND.n3833 19.1543
R20730 GND.n6732 GND.n3836 19.1543
R20731 GND.n6729 GND.n3822 19.1543
R20732 GND.n6742 GND.n3822 19.1543
R20733 GND.n6742 GND.n3823 19.1543
R20734 GND.n3827 GND.n3823 19.1543
R20735 GND.n3827 GND.n3814 19.1543
R20736 GND.n6751 GND.n3814 19.1543
R20737 GND.n6751 GND.n3810 19.1543
R20738 GND.n6757 GND.n3810 19.1543
R20739 GND.n6757 GND.n3812 19.1543
R20740 GND.n6754 GND.n3812 19.1543
R20741 GND.n6754 GND.n3799 19.1543
R20742 GND.n6767 GND.n3799 19.1543
R20743 GND.n6767 GND.n3800 19.1543
R20744 GND.n3804 GND.n3800 19.1543
R20745 GND.n3804 GND.n3792 19.1543
R20746 GND.n6776 GND.n3792 19.1543
R20747 GND.n6776 GND.n3788 19.1543
R20748 GND.n6782 GND.n3788 19.1543
R20749 GND.n6782 GND.n3790 19.1543
R20750 GND.n6778 GND.n3790 19.1543
R20751 GND.n6778 GND.n3773 19.1543
R20752 GND.n6793 GND.n3773 19.1543
R20753 GND.n6793 GND.n3775 19.1543
R20754 GND.n3782 GND.n3775 19.1543
R20755 GND.n3778 GND.n3750 19.1543
R20756 GND.n6878 GND.n3750 19.1543
R20757 GND.n6878 GND.n6877 19.1543
R20758 GND.n6877 GND.n3752 19.1543
R20759 GND.n6802 GND.n3752 19.1543
R20760 GND.n6802 GND.n3759 19.1543
R20761 GND.n6870 GND.n3759 19.1543
R20762 GND.n6870 GND.n3761 19.1543
R20763 GND.n6867 GND.n3761 19.1543
R20764 GND.n6867 GND.n6866 19.1543
R20765 GND.n6866 GND.n6811 19.1543
R20766 GND.n6861 GND.n6811 19.1543
R20767 GND.n6861 GND.n6860 19.1543
R20768 GND.n6860 GND.n6818 19.1543
R20769 GND.n6828 GND.n6818 19.1543
R20770 GND.n6828 GND.n6826 19.1543
R20771 GND.n6853 GND.n6826 19.1543
R20772 GND.n6853 GND.n6827 19.1543
R20773 GND.n6849 GND.n6827 19.1543
R20774 GND.n6849 GND.n6848 19.1543
R20775 GND.n6848 GND.n6840 19.1543
R20776 GND.n6840 GND.n6833 19.1543
R20777 GND.n6833 GND.n3735 19.1543
R20778 GND.n6887 GND.n3735 19.1543
R20779 GND.n6888 GND.n3730 19.1543
R20780 GND.n6892 GND.n3730 19.1543
R20781 GND.n6892 GND.n3732 19.1543
R20782 GND.n3732 GND.n3721 19.1543
R20783 GND.n6903 GND.n3721 19.1543
R20784 GND.n6903 GND.n6902 19.1543
R20785 GND.n6902 GND.n3722 19.1543
R20786 GND.n3722 GND.n3713 19.1543
R20787 GND.n6913 GND.n3713 19.1543
R20788 GND.n6915 GND.n6913 19.1543
R20789 GND.n6915 GND.n3708 19.1543
R20790 GND.n6919 GND.n3708 19.1543
R20791 GND.n6919 GND.n3710 19.1543
R20792 GND.n3710 GND.n3698 19.1543
R20793 GND.n6930 GND.n3698 19.1543
R20794 GND.n6930 GND.n6929 19.1543
R20795 GND.n6929 GND.n3699 19.1543
R20796 GND.n3699 GND.n3691 19.1543
R20797 GND.n6940 GND.n3691 19.1543
R20798 GND.n6942 GND.n6940 19.1543
R20799 GND.n6942 GND.n3687 19.1543
R20800 GND.n6948 GND.n3687 19.1543
R20801 GND.n6948 GND.n3688 19.1543
R20802 GND.n6945 GND.n3688 19.1543
R20803 GND.n6959 GND.n6958 19.1543
R20804 GND.n6958 GND.n3679 19.1543
R20805 GND.n3679 GND.n3671 19.1543
R20806 GND.n6969 GND.n3671 19.1543
R20807 GND.n6970 GND.n6969 19.1543
R20808 GND.n6970 GND.n3667 19.1543
R20809 GND.n6975 GND.n3667 19.1543
R20810 GND.n6975 GND.n3668 19.1543
R20811 GND.n3668 GND.n3657 19.1543
R20812 GND.n6986 GND.n3657 19.1543
R20813 GND.n6986 GND.n6985 19.1543
R20814 GND.n6985 GND.n3659 19.1543
R20815 GND.n3659 GND.n3649 19.1543
R20816 GND.n6996 GND.n3649 19.1543
R20817 GND.n6997 GND.n6996 19.1543
R20818 GND.n6997 GND.n3644 19.1543
R20819 GND.n7001 GND.n3644 19.1543
R20820 GND.n7001 GND.n3646 19.1543
R20821 GND.n3646 GND.n3635 19.1543
R20822 GND.n7012 GND.n3635 19.1543
R20823 GND.n7012 GND.n7011 19.1543
R20824 GND.n7011 GND.n3636 19.1543
R20825 GND.n3636 GND.n3627 19.1543
R20826 GND.n7022 GND.n3627 19.1543
R20827 GND.n7024 GND.n3622 19.1543
R20828 GND.n7028 GND.n3622 19.1543
R20829 GND.n7028 GND.n3624 19.1543
R20830 GND.n3624 GND.n3612 19.1543
R20831 GND.n7039 GND.n3612 19.1543
R20832 GND.n7039 GND.n7038 19.1543
R20833 GND.n7038 GND.n3613 19.1543
R20834 GND.n3613 GND.n3605 19.1543
R20835 GND.n7049 GND.n3605 19.1543
R20836 GND.n7051 GND.n7049 19.1543
R20837 GND.n7051 GND.n3601 19.1543
R20838 GND.n7056 GND.n3601 19.1543
R20839 GND.n7056 GND.n3602 19.1543
R20840 GND.n3602 GND.n3591 19.1543
R20841 GND.n7067 GND.n3591 19.1543
R20842 GND.n7067 GND.n7066 19.1543
R20843 GND.n7066 GND.n3593 19.1543
R20844 GND.n3593 GND.n3584 19.1543
R20845 GND.n7084 GND.n3584 19.1543
R20846 GND.n7085 GND.n7084 19.1543
R20847 GND.n7085 GND.n3578 19.1543
R20848 GND.n7089 GND.n3578 19.1543
R20849 GND.n7089 GND.n3581 19.1543
R20850 GND.n3581 GND.n3580 19.1543
R20851 GND.n3580 GND.n3569 19.1543
R20852 GND.n7099 GND.n3569 19.1543
R20853 GND.n7099 GND.n3571 19.1543
R20854 GND.n3571 GND.n579 19.1543
R20855 GND.t114 GND.n579 19.1543
R20856 GND.n9499 GND.t114 19.1543
R20857 GND.n9499 GND.n567 19.1543
R20858 GND.n9506 GND.n567 19.1543
R20859 GND.n9506 GND.n570 19.1543
R20860 GND.n572 GND.n570 19.1543
R20861 GND.n572 GND.n557 19.1543
R20862 GND.n9516 GND.n557 19.1543
R20863 GND.n9516 GND.n558 19.1543
R20864 GND.n561 GND.n558 19.1543
R20865 GND.n561 GND.n551 19.1543
R20866 GND.n9524 GND.n551 19.1543
R20867 GND.n9524 GND.n476 19.1543
R20868 GND.n9612 GND.n476 19.1543
R20869 GND.n9612 GND.n478 19.1543
R20870 GND.n4839 GND.t121 18.7712
R20871 GND.n6348 GND.t163 18.7712
R20872 GND.n7559 GND.n3012 18.3881
R20873 GND.n4856 GND.n3023 18.3881
R20874 GND.n4620 GND.t9 18.3881
R20875 GND.n5000 GND.n4590 18.3881
R20876 GND.n5050 GND.n4575 18.3881
R20877 GND.n5213 GND.n4490 18.3881
R20878 GND.n5324 GND.n4418 18.3881
R20879 GND.n5375 GND.n4404 18.3881
R20880 GND.n5484 GND.n4332 18.3881
R20881 GND.n5546 GND.n4317 18.3881
R20882 GND.n5638 GND.n4250 18.3881
R20883 GND.n5684 GND.n4235 18.3881
R20884 GND.n5841 GND.n4160 18.3881
R20885 GND.n5970 GND.n4076 18.3881
R20886 GND.n6009 GND.n4061 18.3881
R20887 GND.t26 GND.n6041 18.3881
R20888 GND.n6362 GND.n3989 18.3881
R20889 GND.n3984 GND.n3978 18.3881
R20890 GND.n5145 GND.t19 18.005
R20891 GND.n5852 GND.t14 18.005
R20892 GND.n4820 GND.t98 17.622
R20893 GND.n8151 GND.n1464 16.8558
R20894 GND.n7881 GND.n1814 16.8558
R20895 GND.n7567 GND.n7566 16.8558
R20896 GND.n4907 GND.n4906 16.8558
R20897 GND.n4990 GND.n4988 16.8558
R20898 GND.n5070 GND.n5069 16.8558
R20899 GND.n5153 GND.n5152 16.8558
R20900 GND.n5230 GND.n5229 16.8558
R20901 GND.n5314 GND.n5313 16.8558
R20902 GND.n5392 GND.n5391 16.8558
R20903 GND.n5474 GND.n5473 16.8558
R20904 GND.n5563 GND.n5562 16.8558
R20905 GND.n5630 GND.n5628 16.8558
R20906 GND.n5677 GND.n5676 16.8558
R20907 GND.n4172 GND.n4171 16.8558
R20908 GND.n5878 GND.n5877 16.8558
R20909 GND.n5960 GND.n5959 16.8558
R20910 GND.n6029 GND.n6028 16.8558
R20911 GND.n6341 GND.n3998 16.8558
R20912 GND.n3973 GND.n3232 16.8558
R20913 GND.n7293 GND.n3312 16.8558
R20914 GND.n9567 GND.n519 16.8558
R20915 GND.n9589 GND.n499 15.9035
R20916 GND.n8128 GND.n8127 15.9035
R20917 GND.n50 GND.n48 15.6496
R20918 GND.n73 GND.n71 15.6496
R20919 GND.n93 GND.n91 15.6496
R20920 GND.n116 GND.n114 15.6496
R20921 GND.n7 GND.n5 15.6496
R20922 GND.n30 GND.n28 15.6496
R20923 GND.n305 GND.n303 15.6496
R20924 GND.n282 GND.n280 15.6496
R20925 GND.n348 GND.n346 15.6496
R20926 GND.n325 GND.n323 15.6496
R20927 GND.n392 GND.n390 15.6496
R20928 GND.n369 GND.n367 15.6496
R20929 GND.n195 GND.n194 15.3979
R20930 GND.n183 GND.n182 15.3979
R20931 GND.n171 GND.n170 15.3979
R20932 GND.n159 GND.n158 15.3979
R20933 GND.n147 GND.n146 15.3979
R20934 GND.n136 GND.n135 15.3979
R20935 GND.n266 GND.n265 15.3979
R20936 GND.n254 GND.n253 15.3979
R20937 GND.n242 GND.n241 15.3979
R20938 GND.n230 GND.n229 15.3979
R20939 GND.n218 GND.n217 15.3979
R20940 GND.n207 GND.n206 15.3979
R20941 GND.n7595 GND.n2964 15.3235
R20942 GND.n7573 GND.n2991 15.3235
R20943 GND.n4647 GND.n4642 15.3235
R20944 GND.n4612 GND.n4611 15.3235
R20945 GND.n5116 GND.n4530 15.3235
R20946 GND.n4475 GND.n4470 15.3235
R20947 GND.n4442 GND.n4440 15.3235
R20948 GND.n4389 GND.n4384 15.3235
R20949 GND.n4356 GND.n4355 15.3235
R20950 GND.n4303 GND.n4298 15.3235
R20951 GND.n4270 GND.n4269 15.3235
R20952 GND.n5720 GND.n4209 15.3235
R20953 GND.n5821 GND.n4176 15.3235
R20954 GND.n4134 GND.n4129 15.3235
R20955 GND.n4046 GND.n4041 15.3235
R20956 GND.n6095 GND.n4012 15.3235
R20957 GND.n7334 GND.n3243 15.3235
R20958 GND.n3273 GND.t154 15.3235
R20959 GND.n6199 GND.n6198 15.0827
R20960 GND.n4707 GND.n4702 15.0481
R20961 GND.n6209 GND.n6208 15.0481
R20962 GND.n2964 GND.t108 14.5574
R20963 GND.n4720 GND.n4719 14.0493
R20964 GND.n6255 GND.n6214 14.0493
R20965 GND.n9571 GND.n514 13.9641
R20966 GND.n7887 GND.n7886 13.9641
R20967 GND.n6321 GND.n6320 13.9641
R20968 GND.n8104 GND.n1503 13.9641
R20969 GND.n7588 GND.n7587 13.7912
R20970 GND.n4928 GND.n4636 13.7912
R20971 GND.n4947 GND.n4617 13.7912
R20972 GND.n5089 GND.n4551 13.7912
R20973 GND.n5108 GND.n5107 13.7912
R20974 GND.n5251 GND.n4465 13.7912
R20975 GND.n5270 GND.n4446 13.7912
R20976 GND.n5413 GND.n4379 13.7912
R20977 GND.n5603 GND.n4275 13.7912
R20978 GND.n5730 GND.n4201 13.7912
R20979 GND.n5793 GND.n4186 13.7912
R20980 GND.n5899 GND.n4124 13.7912
R20981 GND.n5918 GND.n4104 13.7912
R20982 GND.n6048 GND.n4037 13.7912
R20983 GND.n6085 GND.n6084 13.7912
R20984 GND.n6378 GND.t142 13.7912
R20985 GND.n6378 GND.n6377 13.7912
R20986 GND.n7315 GND.n3265 13.7912
R20987 GND.n9549 GND.n9548 13.5763
R20988 GND.n7844 GND.n1882 13.5763
R20989 GND.n2407 GND.n2406 13.5763
R20990 GND.n7266 GND.n3348 13.5763
R20991 GND.n4718 GND.n4699 13.1884
R20992 GND.n4713 GND.n4712 13.1884
R20993 GND.n4712 GND.n4711 13.1884
R20994 GND.n6202 GND.n6197 13.1884
R20995 GND.n6203 GND.n6202 13.1884
R20996 GND.n4714 GND.n4701 13.146
R20997 GND.n4710 GND.n4701 13.146
R20998 GND.n6201 GND.n6200 13.146
R20999 GND.n6201 GND.n6196 13.146
R21000 GND.n5313 GND.t8 13.0251
R21001 GND.n5677 GND.t3 13.0251
R21002 GND.n51 GND.n47 12.8005
R21003 GND.n74 GND.n70 12.8005
R21004 GND.n94 GND.n90 12.8005
R21005 GND.n117 GND.n113 12.8005
R21006 GND.n8 GND.n4 12.8005
R21007 GND.n31 GND.n27 12.8005
R21008 GND.n306 GND.n302 12.8005
R21009 GND.n283 GND.n279 12.8005
R21010 GND.n349 GND.n345 12.8005
R21011 GND.n326 GND.n322 12.8005
R21012 GND.n393 GND.n389 12.8005
R21013 GND.n370 GND.n366 12.8005
R21014 GND.n198 GND.n193 12.8005
R21015 GND.n186 GND.n181 12.8005
R21016 GND.n174 GND.n169 12.8005
R21017 GND.n162 GND.n157 12.8005
R21018 GND.n150 GND.n145 12.8005
R21019 GND.n139 GND.n134 12.8005
R21020 GND.n269 GND.n264 12.8005
R21021 GND.n257 GND.n252 12.8005
R21022 GND.n245 GND.n240 12.8005
R21023 GND.n233 GND.n228 12.8005
R21024 GND.n221 GND.n216 12.8005
R21025 GND.n210 GND.n205 12.8005
R21026 GND.n4611 GND.t172 12.642
R21027 GND.t21 GND.n4046 12.642
R21028 GND.n9548 GND.n9547 12.4126
R21029 GND.n7837 GND.n1882 12.4126
R21030 GND.n2408 GND.n2407 12.4126
R21031 GND.n7259 GND.n3348 12.4126
R21032 GND.n7587 GND.n2973 12.2589
R21033 GND.n7581 GND.n2981 12.2589
R21034 GND.n4636 GND.n4627 12.2589
R21035 GND.n4630 GND.n4617 12.2589
R21036 GND.n4551 GND.n4543 12.2589
R21037 GND.n5108 GND.n4536 12.2589
R21038 GND.n4465 GND.n4455 12.2589
R21039 GND.n4459 GND.n4446 12.2589
R21040 GND.n4379 GND.n4369 12.2589
R21041 GND.n5351 GND.n4372 12.2589
R21042 GND.n5495 GND.n4284 12.2589
R21043 GND.n4287 GND.n4275 12.2589
R21044 GND.n5730 GND.n4202 12.2589
R21045 GND.n5794 GND.n5793 12.2589
R21046 GND.n4124 GND.n4114 12.2589
R21047 GND.n4117 GND.n4104 12.2589
R21048 GND.n4037 GND.n4029 12.2589
R21049 GND.n6085 GND.n4020 12.2589
R21050 GND.n6377 GND.n6376 12.2589
R21051 GND.n3265 GND.n3259 12.2589
R21052 GND.n55 GND.n54 12.0247
R21053 GND.n78 GND.n77 12.0247
R21054 GND.n98 GND.n97 12.0247
R21055 GND.n121 GND.n120 12.0247
R21056 GND.n12 GND.n11 12.0247
R21057 GND.n35 GND.n34 12.0247
R21058 GND.n310 GND.n309 12.0247
R21059 GND.n287 GND.n286 12.0247
R21060 GND.n353 GND.n352 12.0247
R21061 GND.n330 GND.n329 12.0247
R21062 GND.n397 GND.n396 12.0247
R21063 GND.n374 GND.n373 12.0247
R21064 GND.n9571 GND.n9570 12.0247
R21065 GND.n7886 GND.n7885 12.0247
R21066 GND.n6322 GND.n6321 12.0247
R21067 GND.n8100 GND.n1503 12.0247
R21068 GND.n199 GND.n191 12.0247
R21069 GND.n187 GND.n179 12.0247
R21070 GND.n175 GND.n167 12.0247
R21071 GND.n163 GND.n155 12.0247
R21072 GND.n151 GND.n143 12.0247
R21073 GND.n140 GND.n132 12.0247
R21074 GND.n270 GND.n262 12.0247
R21075 GND.n258 GND.n250 12.0247
R21076 GND.n246 GND.n238 12.0247
R21077 GND.n234 GND.n226 12.0247
R21078 GND.n222 GND.n214 12.0247
R21079 GND.n211 GND.n203 12.0247
R21080 GND.t53 GND.n2303 11.4928
R21081 GND.t44 GND.n1980 11.4928
R21082 GND.t63 GND.n3883 11.4928
R21083 GND.t49 GND.n7022 11.4928
R21084 GND.n58 GND.n45 11.249
R21085 GND.n81 GND.n68 11.249
R21086 GND.n101 GND.n88 11.249
R21087 GND.n124 GND.n111 11.249
R21088 GND.n15 GND.n2 11.249
R21089 GND.n38 GND.n25 11.249
R21090 GND.n313 GND.n300 11.249
R21091 GND.n290 GND.n277 11.249
R21092 GND.n356 GND.n343 11.249
R21093 GND.n333 GND.n320 11.249
R21094 GND.n400 GND.n387 11.249
R21095 GND.n377 GND.n364 11.249
R21096 GND.n2703 GND.t32 10.7266
R21097 GND.n7668 GND.t36 10.7266
R21098 GND.n7595 GND.n7594 10.7266
R21099 GND.n4920 GND.n4642 10.7266
R21100 GND.n4953 GND.n4612 10.7266
R21101 GND.n5083 GND.n4555 10.7266
R21102 GND.n5117 GND.n5116 10.7266
R21103 GND.n5243 GND.n4470 10.7266
R21104 GND.n5276 GND.n4442 10.7266
R21105 GND.n5405 GND.n4384 10.7266
R21106 GND.n5438 GND.n4356 10.7266
R21107 GND.n5576 GND.n4298 10.7266
R21108 GND.n5609 GND.n4270 10.7266
R21109 GND.n5720 GND.n5719 10.7266
R21110 GND.n4189 GND.n4176 10.7266
R21111 GND.n5891 GND.n4129 10.7266
R21112 GND.n5924 GND.n4100 10.7266
R21113 GND.n6042 GND.n4041 10.7266
R21114 GND.n6095 GND.n4011 10.7266
R21115 GND.n3249 GND.n3243 10.7266
R21116 GND.n7327 GND.t142 10.7266
R21117 GND.n7309 GND.n7308 10.7266
R21118 GND.n6729 GND.t41 10.7266
R21119 GND.n6945 GND.t55 10.7266
R21120 GND.n7905 GND.n7904 10.6672
R21121 GND.n6293 GND.n6292 10.6672
R21122 GND.n6180 GND.n6120 10.6151
R21123 GND.n6180 GND.n6179 10.6151
R21124 GND.n6176 GND.n6175 10.6151
R21125 GND.n6175 GND.n6172 10.6151
R21126 GND.n6172 GND.n6171 10.6151
R21127 GND.n6171 GND.n6168 10.6151
R21128 GND.n6168 GND.n6167 10.6151
R21129 GND.n6167 GND.n6164 10.6151
R21130 GND.n6164 GND.n6163 10.6151
R21131 GND.n6163 GND.n6160 10.6151
R21132 GND.n6160 GND.n6159 10.6151
R21133 GND.n6159 GND.n6156 10.6151
R21134 GND.n6156 GND.n6155 10.6151
R21135 GND.n6155 GND.n6152 10.6151
R21136 GND.n6152 GND.n6151 10.6151
R21137 GND.n6151 GND.n6148 10.6151
R21138 GND.n6148 GND.n6147 10.6151
R21139 GND.n6147 GND.n6144 10.6151
R21140 GND.n6144 GND.n6143 10.6151
R21141 GND.n4811 GND.n4810 10.6151
R21142 GND.n4814 GND.n4811 10.6151
R21143 GND.n4815 GND.n4814 10.6151
R21144 GND.n4816 GND.n4815 10.6151
R21145 GND.n4816 GND.n4673 10.6151
R21146 GND.n4823 GND.n4673 10.6151
R21147 GND.n4824 GND.n4823 10.6151
R21148 GND.n4826 GND.n4824 10.6151
R21149 GND.n4827 GND.n4826 10.6151
R21150 GND.n4828 GND.n4827 10.6151
R21151 GND.n4828 GND.n4672 10.6151
R21152 GND.n4832 GND.n4672 10.6151
R21153 GND.n4833 GND.n4832 10.6151
R21154 GND.n4835 GND.n4833 10.6151
R21155 GND.n4836 GND.n4835 10.6151
R21156 GND.n4837 GND.n4836 10.6151
R21157 GND.n4846 GND.n4837 10.6151
R21158 GND.n4846 GND.n4845 10.6151
R21159 GND.n4845 GND.n4844 10.6151
R21160 GND.n4844 GND.n4842 10.6151
R21161 GND.n4842 GND.n4841 10.6151
R21162 GND.n4841 GND.n4838 10.6151
R21163 GND.n4838 GND.n4644 10.6151
R21164 GND.n4915 GND.n4644 10.6151
R21165 GND.n4916 GND.n4915 10.6151
R21166 GND.n4917 GND.n4916 10.6151
R21167 GND.n4917 GND.n4633 10.6151
R21168 GND.n4930 GND.n4633 10.6151
R21169 GND.n4931 GND.n4930 10.6151
R21170 GND.n4934 GND.n4931 10.6151
R21171 GND.n4934 GND.n4933 10.6151
R21172 GND.n4933 GND.n4932 10.6151
R21173 GND.n4932 GND.n4609 10.6151
R21174 GND.n4955 GND.n4609 10.6151
R21175 GND.n4956 GND.n4955 10.6151
R21176 GND.n4975 GND.n4956 10.6151
R21177 GND.n4975 GND.n4974 10.6151
R21178 GND.n4974 GND.n4973 10.6151
R21179 GND.n4973 GND.n4972 10.6151
R21180 GND.n4972 GND.n4957 10.6151
R21181 GND.n4967 GND.n4957 10.6151
R21182 GND.n4967 GND.n4966 10.6151
R21183 GND.n4966 GND.n4965 10.6151
R21184 GND.n4965 GND.n4964 10.6151
R21185 GND.n4964 GND.n4962 10.6151
R21186 GND.n4962 GND.n4961 10.6151
R21187 GND.n4961 GND.n4959 10.6151
R21188 GND.n4959 GND.n4557 10.6151
R21189 GND.n5078 GND.n4557 10.6151
R21190 GND.n5079 GND.n5078 10.6151
R21191 GND.n5080 GND.n5079 10.6151
R21192 GND.n5080 GND.n4548 10.6151
R21193 GND.n5091 GND.n4548 10.6151
R21194 GND.n5092 GND.n5091 10.6151
R21195 GND.n5099 GND.n5092 10.6151
R21196 GND.n5099 GND.n5098 10.6151
R21197 GND.n5098 GND.n5097 10.6151
R21198 GND.n5097 GND.n5096 10.6151
R21199 GND.n5096 GND.n5094 10.6151
R21200 GND.n5094 GND.n5093 10.6151
R21201 GND.n5093 GND.n4520 10.6151
R21202 GND.n5126 GND.n4520 10.6151
R21203 GND.n5127 GND.n5126 10.6151
R21204 GND.n5130 GND.n5127 10.6151
R21205 GND.n5131 GND.n5130 10.6151
R21206 GND.n5141 GND.n5131 10.6151
R21207 GND.n5141 GND.n5140 10.6151
R21208 GND.n5140 GND.n5139 10.6151
R21209 GND.n5139 GND.n5138 10.6151
R21210 GND.n5138 GND.n5136 10.6151
R21211 GND.n5136 GND.n5135 10.6151
R21212 GND.n5135 GND.n5132 10.6151
R21213 GND.n5132 GND.n4472 10.6151
R21214 GND.n5238 GND.n4472 10.6151
R21215 GND.n5239 GND.n5238 10.6151
R21216 GND.n5240 GND.n5239 10.6151
R21217 GND.n5240 GND.n4461 10.6151
R21218 GND.n5253 GND.n4461 10.6151
R21219 GND.n5254 GND.n5253 10.6151
R21220 GND.n5257 GND.n5254 10.6151
R21221 GND.n5257 GND.n5256 10.6151
R21222 GND.n5256 GND.n5255 10.6151
R21223 GND.n5255 GND.n4437 10.6151
R21224 GND.n5278 GND.n4437 10.6151
R21225 GND.n5279 GND.n5278 10.6151
R21226 GND.n5300 GND.n5279 10.6151
R21227 GND.n5300 GND.n5299 10.6151
R21228 GND.n5299 GND.n5298 10.6151
R21229 GND.n5298 GND.n5297 10.6151
R21230 GND.n5297 GND.n5280 10.6151
R21231 GND.n5291 GND.n5280 10.6151
R21232 GND.n5291 GND.n5290 10.6151
R21233 GND.n5290 GND.n5289 10.6151
R21234 GND.n5289 GND.n5288 10.6151
R21235 GND.n5288 GND.n5286 10.6151
R21236 GND.n5286 GND.n5285 10.6151
R21237 GND.n5285 GND.n5282 10.6151
R21238 GND.n5282 GND.n4386 10.6151
R21239 GND.n5400 GND.n4386 10.6151
R21240 GND.n5401 GND.n5400 10.6151
R21241 GND.n5402 GND.n5401 10.6151
R21242 GND.n5402 GND.n4375 10.6151
R21243 GND.n5415 GND.n4375 10.6151
R21244 GND.n5416 GND.n5415 10.6151
R21245 GND.n5419 GND.n5416 10.6151
R21246 GND.n5419 GND.n5418 10.6151
R21247 GND.n5418 GND.n5417 10.6151
R21248 GND.n5417 GND.n4352 10.6151
R21249 GND.n5440 GND.n4352 10.6151
R21250 GND.n5441 GND.n5440 10.6151
R21251 GND.n5460 GND.n5441 10.6151
R21252 GND.n5460 GND.n5459 10.6151
R21253 GND.n5459 GND.n5458 10.6151
R21254 GND.n5458 GND.n5457 10.6151
R21255 GND.n5457 GND.n5442 10.6151
R21256 GND.n5452 GND.n5442 10.6151
R21257 GND.n5452 GND.n5451 10.6151
R21258 GND.n5451 GND.n5450 10.6151
R21259 GND.n5450 GND.n5449 10.6151
R21260 GND.n5449 GND.n5447 10.6151
R21261 GND.n5447 GND.n5446 10.6151
R21262 GND.n5446 GND.n5444 10.6151
R21263 GND.n5444 GND.n4300 10.6151
R21264 GND.n5571 GND.n4300 10.6151
R21265 GND.n5572 GND.n5571 10.6151
R21266 GND.n5573 GND.n5572 10.6151
R21267 GND.n5573 GND.n4290 10.6151
R21268 GND.n5586 GND.n4290 10.6151
R21269 GND.n5587 GND.n5586 10.6151
R21270 GND.n5590 GND.n5587 10.6151
R21271 GND.n5590 GND.n5589 10.6151
R21272 GND.n5589 GND.n5588 10.6151
R21273 GND.n5588 GND.n4266 10.6151
R21274 GND.n5611 GND.n4266 10.6151
R21275 GND.n5612 GND.n5611 10.6151
R21276 GND.n5620 GND.n5612 10.6151
R21277 GND.n5620 GND.n5619 10.6151
R21278 GND.n5619 GND.n5618 10.6151
R21279 GND.n5618 GND.n5617 10.6151
R21280 GND.n5617 GND.n5614 10.6151
R21281 GND.n5614 GND.n5613 10.6151
R21282 GND.n5613 GND.n4242 10.6151
R21283 GND.n5648 GND.n4242 10.6151
R21284 GND.n5649 GND.n5648 10.6151
R21285 GND.n5652 GND.n5649 10.6151
R21286 GND.n5653 GND.n5652 10.6151
R21287 GND.n5674 GND.n5653 10.6151
R21288 GND.n5674 GND.n5673 10.6151
R21289 GND.n5673 GND.n5672 10.6151
R21290 GND.n5672 GND.n5671 10.6151
R21291 GND.n5671 GND.n5669 10.6151
R21292 GND.n5669 GND.n5668 10.6151
R21293 GND.n5668 GND.n5654 10.6151
R21294 GND.n5664 GND.n5654 10.6151
R21295 GND.n5664 GND.n5663 10.6151
R21296 GND.n5663 GND.n5662 10.6151
R21297 GND.n5662 GND.n5661 10.6151
R21298 GND.n5661 GND.n5659 10.6151
R21299 GND.n5659 GND.n5658 10.6151
R21300 GND.n5658 GND.n5656 10.6151
R21301 GND.n5656 GND.n4168 10.6151
R21302 GND.n5829 GND.n4168 10.6151
R21303 GND.n5830 GND.n5829 10.6151
R21304 GND.n5832 GND.n5830 10.6151
R21305 GND.n5832 GND.n5831 10.6151
R21306 GND.n5831 GND.n4158 10.6151
R21307 GND.n5844 GND.n4158 10.6151
R21308 GND.n5845 GND.n5844 10.6151
R21309 GND.n5850 GND.n5845 10.6151
R21310 GND.n5850 GND.n5849 10.6151
R21311 GND.n5849 GND.n5848 10.6151
R21312 GND.n5848 GND.n5846 10.6151
R21313 GND.n5846 GND.n4131 10.6151
R21314 GND.n5886 GND.n4131 10.6151
R21315 GND.n5887 GND.n5886 10.6151
R21316 GND.n5888 GND.n5887 10.6151
R21317 GND.n5888 GND.n4120 10.6151
R21318 GND.n5901 GND.n4120 10.6151
R21319 GND.n5902 GND.n5901 10.6151
R21320 GND.n5905 GND.n5902 10.6151
R21321 GND.n5905 GND.n5904 10.6151
R21322 GND.n5904 GND.n5903 10.6151
R21323 GND.n5903 GND.n4096 10.6151
R21324 GND.n5926 GND.n4096 10.6151
R21325 GND.n5927 GND.n5926 10.6151
R21326 GND.n5946 GND.n5927 10.6151
R21327 GND.n5946 GND.n5945 10.6151
R21328 GND.n5945 GND.n5944 10.6151
R21329 GND.n5944 GND.n5943 10.6151
R21330 GND.n5943 GND.n5928 10.6151
R21331 GND.n5938 GND.n5928 10.6151
R21332 GND.n5938 GND.n5937 10.6151
R21333 GND.n5937 GND.n5936 10.6151
R21334 GND.n5936 GND.n5935 10.6151
R21335 GND.n5935 GND.n5933 10.6151
R21336 GND.n5933 GND.n5932 10.6151
R21337 GND.n5932 GND.n5930 10.6151
R21338 GND.n5930 GND.n4043 10.6151
R21339 GND.n6037 GND.n4043 10.6151
R21340 GND.n6038 GND.n6037 10.6151
R21341 GND.n6039 GND.n6038 10.6151
R21342 GND.n6039 GND.n4033 10.6151
R21343 GND.n6050 GND.n4033 10.6151
R21344 GND.n6051 GND.n6050 10.6151
R21345 GND.n6071 GND.n6051 10.6151
R21346 GND.n6071 GND.n6070 10.6151
R21347 GND.n6070 GND.n6069 10.6151
R21348 GND.n6069 GND.n6068 10.6151
R21349 GND.n6068 GND.n6052 10.6151
R21350 GND.n6063 GND.n6052 10.6151
R21351 GND.n6063 GND.n6062 10.6151
R21352 GND.n6062 GND.n6061 10.6151
R21353 GND.n6061 GND.n6060 10.6151
R21354 GND.n6060 GND.n6058 10.6151
R21355 GND.n6058 GND.n6057 10.6151
R21356 GND.n6057 GND.n6054 10.6151
R21357 GND.n6054 GND.n3981 10.6151
R21358 GND.n6371 GND.n3981 10.6151
R21359 GND.n6372 GND.n6371 10.6151
R21360 GND.n6391 GND.n6372 10.6151
R21361 GND.n6391 GND.n6390 10.6151
R21362 GND.n6390 GND.n6389 10.6151
R21363 GND.n6389 GND.n6387 10.6151
R21364 GND.n6387 GND.n6386 10.6151
R21365 GND.n6386 GND.n6384 10.6151
R21366 GND.n6384 GND.n6383 10.6151
R21367 GND.n6383 GND.n6381 10.6151
R21368 GND.n6381 GND.n6380 10.6151
R21369 GND.n6380 GND.n3262 10.6151
R21370 GND.n7319 GND.n3262 10.6151
R21371 GND.n7319 GND.n7318 10.6151
R21372 GND.n7318 GND.n7317 10.6151
R21373 GND.n7317 GND.n3263 10.6151
R21374 GND.n6138 GND.n3263 10.6151
R21375 GND.n6139 GND.n6138 10.6151
R21376 GND.n4770 GND.n4686 10.6151
R21377 GND.n4771 GND.n4770 10.6151
R21378 GND.n4773 GND.n4682 10.6151
R21379 GND.n4779 GND.n4682 10.6151
R21380 GND.n4780 GND.n4779 10.6151
R21381 GND.n4781 GND.n4780 10.6151
R21382 GND.n4781 GND.n4680 10.6151
R21383 GND.n4787 GND.n4680 10.6151
R21384 GND.n4788 GND.n4787 10.6151
R21385 GND.n4789 GND.n4788 10.6151
R21386 GND.n4789 GND.n4678 10.6151
R21387 GND.n4795 GND.n4678 10.6151
R21388 GND.n4796 GND.n4795 10.6151
R21389 GND.n4797 GND.n4796 10.6151
R21390 GND.n4797 GND.n4676 10.6151
R21391 GND.n4803 GND.n4676 10.6151
R21392 GND.n4804 GND.n4803 10.6151
R21393 GND.n4805 GND.n4804 10.6151
R21394 GND.n4805 GND.n4674 10.6151
R21395 GND.n4724 GND.n4720 10.6151
R21396 GND.n4725 GND.n4724 10.6151
R21397 GND.n4726 GND.n4725 10.6151
R21398 GND.n4726 GND.n4697 10.6151
R21399 GND.n4732 GND.n4697 10.6151
R21400 GND.n4733 GND.n4732 10.6151
R21401 GND.n4734 GND.n4733 10.6151
R21402 GND.n4734 GND.n4695 10.6151
R21403 GND.n4740 GND.n4695 10.6151
R21404 GND.n4741 GND.n4740 10.6151
R21405 GND.n4742 GND.n4741 10.6151
R21406 GND.n4742 GND.n4693 10.6151
R21407 GND.n4748 GND.n4693 10.6151
R21408 GND.n4749 GND.n4748 10.6151
R21409 GND.n4750 GND.n4749 10.6151
R21410 GND.n4750 GND.n4691 10.6151
R21411 GND.n4756 GND.n4691 10.6151
R21412 GND.n4759 GND.n4758 10.6151
R21413 GND.n4759 GND.n4687 10.6151
R21414 GND.n6255 GND.n6254 10.6151
R21415 GND.n6254 GND.n6253 10.6151
R21416 GND.n6253 GND.n6250 10.6151
R21417 GND.n6250 GND.n6249 10.6151
R21418 GND.n6249 GND.n6246 10.6151
R21419 GND.n6246 GND.n6245 10.6151
R21420 GND.n6245 GND.n6242 10.6151
R21421 GND.n6242 GND.n6241 10.6151
R21422 GND.n6241 GND.n6238 10.6151
R21423 GND.n6238 GND.n6237 10.6151
R21424 GND.n6237 GND.n6234 10.6151
R21425 GND.n6234 GND.n6233 10.6151
R21426 GND.n6233 GND.n6230 10.6151
R21427 GND.n6230 GND.n6229 10.6151
R21428 GND.n6229 GND.n6226 10.6151
R21429 GND.n6226 GND.n6225 10.6151
R21430 GND.n6225 GND.n6222 10.6151
R21431 GND.n6220 GND.n6217 10.6151
R21432 GND.n6217 GND.n6121 10.6151
R21433 GND.n7592 GND.n2968 10.6151
R21434 GND.n7592 GND.n7591 10.6151
R21435 GND.n7591 GND.n7590 10.6151
R21436 GND.n7590 GND.n2969 10.6151
R21437 GND.n4818 GND.n2969 10.6151
R21438 GND.n4818 GND.n2986 10.6151
R21439 GND.n7578 GND.n2986 10.6151
R21440 GND.n7578 GND.n7577 10.6151
R21441 GND.n7577 GND.n7576 10.6151
R21442 GND.n7576 GND.n2987 10.6151
R21443 GND.n3005 GND.n2987 10.6151
R21444 GND.n3006 GND.n3005 10.6151
R21445 GND.n7564 GND.n3006 10.6151
R21446 GND.n7564 GND.n7563 10.6151
R21447 GND.n7563 GND.n7562 10.6151
R21448 GND.n7562 GND.n3007 10.6151
R21449 GND.n4661 GND.n3007 10.6151
R21450 GND.n4851 GND.n4661 10.6151
R21451 GND.n4852 GND.n4851 10.6151
R21452 GND.n4853 GND.n4852 10.6151
R21453 GND.n4853 GND.n4650 10.6151
R21454 GND.n4909 GND.n4650 10.6151
R21455 GND.n4910 GND.n4909 10.6151
R21456 GND.n4911 GND.n4910 10.6151
R21457 GND.n4911 GND.n4639 10.6151
R21458 GND.n4922 GND.n4639 10.6151
R21459 GND.n4923 GND.n4922 10.6151
R21460 GND.n4926 GND.n4923 10.6151
R21461 GND.n4926 GND.n4925 10.6151
R21462 GND.n4925 GND.n4924 10.6151
R21463 GND.n4924 GND.n4614 10.6151
R21464 GND.n4949 GND.n4614 10.6151
R21465 GND.n4950 GND.n4949 10.6151
R21466 GND.n4951 GND.n4950 10.6151
R21467 GND.n4951 GND.n4604 10.6151
R21468 GND.n4979 GND.n4604 10.6151
R21469 GND.n4980 GND.n4979 10.6151
R21470 GND.n4986 GND.n4980 10.6151
R21471 GND.n4986 GND.n4985 10.6151
R21472 GND.n4985 GND.n4984 10.6151
R21473 GND.n4984 GND.n4981 10.6151
R21474 GND.n4981 GND.n4580 10.6151
R21475 GND.n5045 GND.n4580 10.6151
R21476 GND.n5046 GND.n5045 10.6151
R21477 GND.n5047 GND.n5046 10.6151
R21478 GND.n5047 GND.n4564 10.6151
R21479 GND.n5072 GND.n4564 10.6151
R21480 GND.n5073 GND.n5072 10.6151
R21481 GND.n5074 GND.n5073 10.6151
R21482 GND.n5074 GND.n4553 10.6151
R21483 GND.n5085 GND.n4553 10.6151
R21484 GND.n5086 GND.n5085 10.6151
R21485 GND.n5087 GND.n5086 10.6151
R21486 GND.n5087 GND.n4541 10.6151
R21487 GND.n5103 GND.n4541 10.6151
R21488 GND.n5104 GND.n5103 10.6151
R21489 GND.n5105 GND.n5104 10.6151
R21490 GND.n5105 GND.n4525 10.6151
R21491 GND.n5119 GND.n4525 10.6151
R21492 GND.n5120 GND.n5119 10.6151
R21493 GND.n5121 GND.n5120 10.6151
R21494 GND.n5121 GND.n4516 10.6151
R21495 GND.n5150 GND.n4516 10.6151
R21496 GND.n5150 GND.n5149 10.6151
R21497 GND.n5149 GND.n5148 10.6151
R21498 GND.n5148 GND.n4517 10.6151
R21499 GND.n4517 GND.n4494 10.6151
R21500 GND.n5208 GND.n4494 10.6151
R21501 GND.n5209 GND.n5208 10.6151
R21502 GND.n5210 GND.n5209 10.6151
R21503 GND.n5210 GND.n4478 10.6151
R21504 GND.n5232 GND.n4478 10.6151
R21505 GND.n5233 GND.n5232 10.6151
R21506 GND.n5234 GND.n5233 10.6151
R21507 GND.n5234 GND.n4468 10.6151
R21508 GND.n5245 GND.n4468 10.6151
R21509 GND.n5246 GND.n5245 10.6151
R21510 GND.n5249 GND.n5246 10.6151
R21511 GND.n5249 GND.n5248 10.6151
R21512 GND.n5248 GND.n5247 10.6151
R21513 GND.n5247 GND.n4444 10.6151
R21514 GND.n5272 GND.n4444 10.6151
R21515 GND.n5273 GND.n5272 10.6151
R21516 GND.n5274 GND.n5273 10.6151
R21517 GND.n5274 GND.n4432 10.6151
R21518 GND.n5304 GND.n4432 10.6151
R21519 GND.n5305 GND.n5304 10.6151
R21520 GND.n5311 GND.n5305 10.6151
R21521 GND.n5311 GND.n5310 10.6151
R21522 GND.n5310 GND.n5309 10.6151
R21523 GND.n5309 GND.n5306 10.6151
R21524 GND.n5306 GND.n4408 10.6151
R21525 GND.n5370 GND.n4408 10.6151
R21526 GND.n5371 GND.n5370 10.6151
R21527 GND.n5372 GND.n5371 10.6151
R21528 GND.n5372 GND.n4392 10.6151
R21529 GND.n5394 GND.n4392 10.6151
R21530 GND.n5395 GND.n5394 10.6151
R21531 GND.n5396 GND.n5395 10.6151
R21532 GND.n5396 GND.n4382 10.6151
R21533 GND.n5407 GND.n4382 10.6151
R21534 GND.n5408 GND.n5407 10.6151
R21535 GND.n5411 GND.n5408 10.6151
R21536 GND.n5411 GND.n5410 10.6151
R21537 GND.n5410 GND.n5409 10.6151
R21538 GND.n5409 GND.n4358 10.6151
R21539 GND.n5434 GND.n4358 10.6151
R21540 GND.n5435 GND.n5434 10.6151
R21541 GND.n5436 GND.n5435 10.6151
R21542 GND.n5436 GND.n4347 10.6151
R21543 GND.n5464 GND.n4347 10.6151
R21544 GND.n5465 GND.n5464 10.6151
R21545 GND.n5471 GND.n5465 10.6151
R21546 GND.n5471 GND.n5470 10.6151
R21547 GND.n5470 GND.n5469 10.6151
R21548 GND.n5469 GND.n5466 10.6151
R21549 GND.n5466 GND.n4322 10.6151
R21550 GND.n5540 GND.n4322 10.6151
R21551 GND.n5541 GND.n5540 10.6151
R21552 GND.n5542 GND.n5541 10.6151
R21553 GND.n5542 GND.n4306 10.6151
R21554 GND.n5565 GND.n4306 10.6151
R21555 GND.n5566 GND.n5565 10.6151
R21556 GND.n5567 GND.n5566 10.6151
R21557 GND.n5567 GND.n4295 10.6151
R21558 GND.n5578 GND.n4295 10.6151
R21559 GND.n5579 GND.n5578 10.6151
R21560 GND.n5582 GND.n5579 10.6151
R21561 GND.n5582 GND.n5581 10.6151
R21562 GND.n5581 GND.n5580 10.6151
R21563 GND.n5580 GND.n4272 10.6151
R21564 GND.n5605 GND.n4272 10.6151
R21565 GND.n5606 GND.n5605 10.6151
R21566 GND.n5607 GND.n5606 10.6151
R21567 GND.n5607 GND.n4261 10.6151
R21568 GND.n5624 GND.n4261 10.6151
R21569 GND.n5625 GND.n5624 10.6151
R21570 GND.n5626 GND.n5625 10.6151
R21571 GND.n5626 GND.n4246 10.6151
R21572 GND.n5641 GND.n4246 10.6151
R21573 GND.n5642 GND.n5641 10.6151
R21574 GND.n5643 GND.n5642 10.6151
R21575 GND.n5643 GND.n4238 10.6151
R21576 GND.n5682 GND.n4238 10.6151
R21577 GND.n5682 GND.n5681 10.6151
R21578 GND.n5681 GND.n5680 10.6151
R21579 GND.n5680 GND.n4239 10.6151
R21580 GND.n4239 GND.n4216 10.6151
R21581 GND.n5710 GND.n4216 10.6151
R21582 GND.n5711 GND.n5710 10.6151
R21583 GND.n5717 GND.n5711 10.6151
R21584 GND.n5717 GND.n5716 10.6151
R21585 GND.n5716 GND.n5715 10.6151
R21586 GND.n5715 GND.n5712 10.6151
R21587 GND.n5712 GND.n4191 10.6151
R21588 GND.n5796 GND.n4191 10.6151
R21589 GND.n5797 GND.n5796 10.6151
R21590 GND.n5798 GND.n5797 10.6151
R21591 GND.n5798 GND.n4174 10.6151
R21592 GND.n5823 GND.n4174 10.6151
R21593 GND.n5824 GND.n5823 10.6151
R21594 GND.n5825 GND.n5824 10.6151
R21595 GND.n5825 GND.n4164 10.6151
R21596 GND.n5837 GND.n4164 10.6151
R21597 GND.n5838 GND.n5837 10.6151
R21598 GND.n5839 GND.n5838 10.6151
R21599 GND.n5839 GND.n4153 10.6151
R21600 GND.n5856 GND.n4153 10.6151
R21601 GND.n5857 GND.n5856 10.6151
R21602 GND.n5858 GND.n5857 10.6151
R21603 GND.n5858 GND.n4137 10.6151
R21604 GND.n5880 GND.n4137 10.6151
R21605 GND.n5881 GND.n5880 10.6151
R21606 GND.n5882 GND.n5881 10.6151
R21607 GND.n5882 GND.n4127 10.6151
R21608 GND.n5893 GND.n4127 10.6151
R21609 GND.n5894 GND.n5893 10.6151
R21610 GND.n5897 GND.n5894 10.6151
R21611 GND.n5897 GND.n5896 10.6151
R21612 GND.n5896 GND.n5895 10.6151
R21613 GND.n5895 GND.n4102 10.6151
R21614 GND.n5920 GND.n4102 10.6151
R21615 GND.n5921 GND.n5920 10.6151
R21616 GND.n5922 GND.n5921 10.6151
R21617 GND.n5922 GND.n4091 10.6151
R21618 GND.n5950 GND.n4091 10.6151
R21619 GND.n5951 GND.n5950 10.6151
R21620 GND.n5957 GND.n5951 10.6151
R21621 GND.n5957 GND.n5956 10.6151
R21622 GND.n5956 GND.n5955 10.6151
R21623 GND.n5955 GND.n5952 10.6151
R21624 GND.n5952 GND.n4066 10.6151
R21625 GND.n6004 GND.n4066 10.6151
R21626 GND.n6005 GND.n6004 10.6151
R21627 GND.n6006 GND.n6005 10.6151
R21628 GND.n6006 GND.n4049 10.6151
R21629 GND.n6031 GND.n4049 10.6151
R21630 GND.n6032 GND.n6031 10.6151
R21631 GND.n6033 GND.n6032 10.6151
R21632 GND.n6033 GND.n4039 10.6151
R21633 GND.n6044 GND.n4039 10.6151
R21634 GND.n6045 GND.n6044 10.6151
R21635 GND.n6046 GND.n6045 10.6151
R21636 GND.n6046 GND.n4027 10.6151
R21637 GND.n6075 GND.n4027 10.6151
R21638 GND.n6076 GND.n6075 10.6151
R21639 GND.n6082 GND.n6076 10.6151
R21640 GND.n6082 GND.n6081 10.6151
R21641 GND.n6081 GND.n6080 10.6151
R21642 GND.n6080 GND.n6077 10.6151
R21643 GND.n6077 GND.n4002 10.6151
R21644 GND.n6344 GND.n4002 10.6151
R21645 GND.n6345 GND.n6344 10.6151
R21646 GND.n6346 GND.n6345 10.6151
R21647 GND.n6346 GND.n3987 10.6151
R21648 GND.n6364 GND.n3987 10.6151
R21649 GND.n6365 GND.n6364 10.6151
R21650 GND.n6367 GND.n6365 10.6151
R21651 GND.n6367 GND.n6366 10.6151
R21652 GND.n6366 GND.n3976 10.6151
R21653 GND.n6396 GND.n3976 10.6151
R21654 GND.n6397 GND.n6396 10.6151
R21655 GND.n6398 GND.n6397 10.6151
R21656 GND.n6398 GND.n3246 10.6151
R21657 GND.n7332 GND.n3246 10.6151
R21658 GND.n7332 GND.n7331 10.6151
R21659 GND.n7331 GND.n7330 10.6151
R21660 GND.n7330 GND.n3247 10.6151
R21661 GND.n6374 GND.n3247 10.6151
R21662 GND.n6374 GND.n6373 10.6151
R21663 GND.n6373 GND.n3268 10.6151
R21664 GND.n7313 GND.n3268 10.6151
R21665 GND.n7313 GND.n7312 10.6151
R21666 GND.n7312 GND.n7311 10.6151
R21667 GND.n7311 GND.n3269 10.6151
R21668 GND.n59 GND.n43 10.4732
R21669 GND.n82 GND.n66 10.4732
R21670 GND.n102 GND.n86 10.4732
R21671 GND.n125 GND.n109 10.4732
R21672 GND.n16 GND.n0 10.4732
R21673 GND.n39 GND.n23 10.4732
R21674 GND.n314 GND.n298 10.4732
R21675 GND.n291 GND.n275 10.4732
R21676 GND.n357 GND.n341 10.4732
R21677 GND.n334 GND.n318 10.4732
R21678 GND.n401 GND.n385 10.4732
R21679 GND.n378 GND.n362 10.4732
R21680 GND.t172 GND.n4606 10.3435
R21681 GND.n4560 GND.t27 10.3435
R21682 GND.t24 GND.n4098 10.3435
R21683 GND.n4047 GND.t21 10.3435
R21684 GND.n9593 GND.n499 10.0853
R21685 GND.n8131 GND.n8128 10.0853
R21686 GND.n2667 GND.t39 9.96045
R21687 GND.t65 GND.n2099 9.96045
R21688 GND.n7308 GND.t170 9.96045
R21689 GND.t46 GND.n3778 9.96045
R21690 GND.t34 GND.n6887 9.96045
R21691 GND.n61 GND.n60 9.45567
R21692 GND.n84 GND.n83 9.45567
R21693 GND.n104 GND.n103 9.45567
R21694 GND.n127 GND.n126 9.45567
R21695 GND.n18 GND.n17 9.45567
R21696 GND.n41 GND.n40 9.45567
R21697 GND.n316 GND.n315 9.45567
R21698 GND.n293 GND.n292 9.45567
R21699 GND.n359 GND.n358 9.45567
R21700 GND.n336 GND.n335 9.45567
R21701 GND.n403 GND.n402 9.45567
R21702 GND.n380 GND.n379 9.45567
R21703 GND.n201 GND.n200 9.45567
R21704 GND.n189 GND.n188 9.45567
R21705 GND.n177 GND.n176 9.45567
R21706 GND.n165 GND.n164 9.45567
R21707 GND.n153 GND.n152 9.45567
R21708 GND.n142 GND.n141 9.45567
R21709 GND.n272 GND.n271 9.45567
R21710 GND.n260 GND.n259 9.45567
R21711 GND.n248 GND.n247 9.45567
R21712 GND.n236 GND.n235 9.45567
R21713 GND.n224 GND.n223 9.45567
R21714 GND.n213 GND.n212 9.45567
R21715 GND.n60 GND.n59 9.3005
R21716 GND.n45 GND.n44 9.3005
R21717 GND.n54 GND.n53 9.3005
R21718 GND.n52 GND.n51 9.3005
R21719 GND.n83 GND.n82 9.3005
R21720 GND.n68 GND.n67 9.3005
R21721 GND.n77 GND.n76 9.3005
R21722 GND.n75 GND.n74 9.3005
R21723 GND.n103 GND.n102 9.3005
R21724 GND.n88 GND.n87 9.3005
R21725 GND.n97 GND.n96 9.3005
R21726 GND.n95 GND.n94 9.3005
R21727 GND.n126 GND.n125 9.3005
R21728 GND.n111 GND.n110 9.3005
R21729 GND.n120 GND.n119 9.3005
R21730 GND.n118 GND.n117 9.3005
R21731 GND.n17 GND.n16 9.3005
R21732 GND.n2 GND.n1 9.3005
R21733 GND.n11 GND.n10 9.3005
R21734 GND.n9 GND.n8 9.3005
R21735 GND.n40 GND.n39 9.3005
R21736 GND.n25 GND.n24 9.3005
R21737 GND.n34 GND.n33 9.3005
R21738 GND.n32 GND.n31 9.3005
R21739 GND.n315 GND.n314 9.3005
R21740 GND.n300 GND.n299 9.3005
R21741 GND.n309 GND.n308 9.3005
R21742 GND.n307 GND.n306 9.3005
R21743 GND.n292 GND.n291 9.3005
R21744 GND.n277 GND.n276 9.3005
R21745 GND.n286 GND.n285 9.3005
R21746 GND.n284 GND.n283 9.3005
R21747 GND.n358 GND.n357 9.3005
R21748 GND.n343 GND.n342 9.3005
R21749 GND.n352 GND.n351 9.3005
R21750 GND.n350 GND.n349 9.3005
R21751 GND.n335 GND.n334 9.3005
R21752 GND.n320 GND.n319 9.3005
R21753 GND.n329 GND.n328 9.3005
R21754 GND.n327 GND.n326 9.3005
R21755 GND.n402 GND.n401 9.3005
R21756 GND.n387 GND.n386 9.3005
R21757 GND.n396 GND.n395 9.3005
R21758 GND.n394 GND.n393 9.3005
R21759 GND.n379 GND.n378 9.3005
R21760 GND.n364 GND.n363 9.3005
R21761 GND.n373 GND.n372 9.3005
R21762 GND.n371 GND.n370 9.3005
R21763 GND.n4665 GND.n4662 9.3005
R21764 GND.n4667 GND.n4666 9.3005
R21765 GND.n4658 GND.n4657 9.3005
R21766 GND.n4859 GND.n4858 9.3005
R21767 GND.n4860 GND.n4656 9.3005
R21768 GND.n4888 GND.n4861 9.3005
R21769 GND.n4887 GND.n4862 9.3005
R21770 GND.n4886 GND.n4863 9.3005
R21771 GND.n4865 GND.n4864 9.3005
R21772 GND.n4882 GND.n4866 9.3005
R21773 GND.n4881 GND.n4867 9.3005
R21774 GND.n4880 GND.n4868 9.3005
R21775 GND.n4878 GND.n4869 9.3005
R21776 GND.n4877 GND.n4870 9.3005
R21777 GND.n4874 GND.n4871 9.3005
R21778 GND.n4873 GND.n4872 9.3005
R21779 GND.n4587 GND.n4586 9.3005
R21780 GND.n5003 GND.n5002 9.3005
R21781 GND.n5004 GND.n4585 9.3005
R21782 GND.n5039 GND.n5005 9.3005
R21783 GND.n5038 GND.n5006 9.3005
R21784 GND.n5037 GND.n5007 9.3005
R21785 GND.n5035 GND.n5008 9.3005
R21786 GND.n5034 GND.n5009 9.3005
R21787 GND.n5012 GND.n5010 9.3005
R21788 GND.n5030 GND.n5013 9.3005
R21789 GND.n5029 GND.n5014 9.3005
R21790 GND.n5028 GND.n5015 9.3005
R21791 GND.n5027 GND.n5016 9.3005
R21792 GND.n5026 GND.n5017 9.3005
R21793 GND.n5024 GND.n5018 9.3005
R21794 GND.n5023 GND.n5019 9.3005
R21795 GND.n5021 GND.n5020 9.3005
R21796 GND.n4501 GND.n4500 9.3005
R21797 GND.n5166 GND.n5165 9.3005
R21798 GND.n5167 GND.n4499 9.3005
R21799 GND.n5203 GND.n5168 9.3005
R21800 GND.n5202 GND.n5169 9.3005
R21801 GND.n5201 GND.n5170 9.3005
R21802 GND.n5199 GND.n5171 9.3005
R21803 GND.n5198 GND.n5172 9.3005
R21804 GND.n5175 GND.n5173 9.3005
R21805 GND.n5194 GND.n5176 9.3005
R21806 GND.n5193 GND.n5177 9.3005
R21807 GND.n5192 GND.n5178 9.3005
R21808 GND.n5191 GND.n5179 9.3005
R21809 GND.n5189 GND.n5180 9.3005
R21810 GND.n5188 GND.n5181 9.3005
R21811 GND.n5185 GND.n5182 9.3005
R21812 GND.n5184 GND.n5183 9.3005
R21813 GND.n4415 GND.n4414 9.3005
R21814 GND.n5327 GND.n5326 9.3005
R21815 GND.n5328 GND.n4413 9.3005
R21816 GND.n5365 GND.n5329 9.3005
R21817 GND.n5364 GND.n5330 9.3005
R21818 GND.n5363 GND.n5331 9.3005
R21819 GND.n5361 GND.n5332 9.3005
R21820 GND.n5360 GND.n5333 9.3005
R21821 GND.n5336 GND.n5334 9.3005
R21822 GND.n5356 GND.n5337 9.3005
R21823 GND.n5355 GND.n5338 9.3005
R21824 GND.n5354 GND.n5339 9.3005
R21825 GND.n5353 GND.n5340 9.3005
R21826 GND.n5350 GND.n5341 9.3005
R21827 GND.n5349 GND.n5342 9.3005
R21828 GND.n5346 GND.n5343 9.3005
R21829 GND.n5345 GND.n5344 9.3005
R21830 GND.n4329 GND.n4328 9.3005
R21831 GND.n5487 GND.n5486 9.3005
R21832 GND.n5488 GND.n4327 9.3005
R21833 GND.n5535 GND.n5489 9.3005
R21834 GND.n5534 GND.n5490 9.3005
R21835 GND.n5533 GND.n5491 9.3005
R21836 GND.n5531 GND.n5492 9.3005
R21837 GND.n5530 GND.n5493 9.3005
R21838 GND.n5497 GND.n5494 9.3005
R21839 GND.n5526 GND.n5498 9.3005
R21840 GND.n5525 GND.n5499 9.3005
R21841 GND.n5524 GND.n5500 9.3005
R21842 GND.n5523 GND.n5501 9.3005
R21843 GND.n5521 GND.n5502 9.3005
R21844 GND.n5520 GND.n5503 9.3005
R21845 GND.n5517 GND.n5504 9.3005
R21846 GND.n5516 GND.n5505 9.3005
R21847 GND.n5515 GND.n5506 9.3005
R21848 GND.n5513 GND.n5507 9.3005
R21849 GND.n5512 GND.n5508 9.3005
R21850 GND.n5510 GND.n5509 9.3005
R21851 GND.n4223 GND.n4222 9.3005
R21852 GND.n5699 GND.n5698 9.3005
R21853 GND.n5700 GND.n4221 9.3005
R21854 GND.n5704 GND.n5701 9.3005
R21855 GND.n5703 GND.n5702 9.3005
R21856 GND.n4199 GND.n4198 9.3005
R21857 GND.n5733 GND.n5732 9.3005
R21858 GND.n5734 GND.n4197 9.3005
R21859 GND.n5791 GND.n5735 9.3005
R21860 GND.n5790 GND.n5736 9.3005
R21861 GND.n5789 GND.n5737 9.3005
R21862 GND.n5787 GND.n5738 9.3005
R21863 GND.n5786 GND.n5739 9.3005
R21864 GND.n5742 GND.n5740 9.3005
R21865 GND.n5782 GND.n5743 9.3005
R21866 GND.n5781 GND.n5744 9.3005
R21867 GND.n5780 GND.n5745 9.3005
R21868 GND.n5779 GND.n5746 9.3005
R21869 GND.n5778 GND.n5747 9.3005
R21870 GND.n5776 GND.n5748 9.3005
R21871 GND.n5775 GND.n5749 9.3005
R21872 GND.n5752 GND.n5750 9.3005
R21873 GND.n5771 GND.n5753 9.3005
R21874 GND.n5770 GND.n5754 9.3005
R21875 GND.n5769 GND.n5755 9.3005
R21876 GND.n5768 GND.n5756 9.3005
R21877 GND.n5766 GND.n5757 9.3005
R21878 GND.n5765 GND.n5758 9.3005
R21879 GND.n5762 GND.n5759 9.3005
R21880 GND.n5761 GND.n5760 9.3005
R21881 GND.n4073 GND.n4072 9.3005
R21882 GND.n5973 GND.n5972 9.3005
R21883 GND.n5974 GND.n4071 9.3005
R21884 GND.n5999 GND.n5975 9.3005
R21885 GND.n5998 GND.n5976 9.3005
R21886 GND.n5997 GND.n5977 9.3005
R21887 GND.n5995 GND.n5978 9.3005
R21888 GND.n5994 GND.n5979 9.3005
R21889 GND.n5982 GND.n5980 9.3005
R21890 GND.n5990 GND.n5983 9.3005
R21891 GND.n5989 GND.n5984 9.3005
R21892 GND.n5988 GND.n5985 9.3005
R21893 GND.n5987 GND.n5986 9.3005
R21894 GND.n4009 GND.n4008 9.3005
R21895 GND.n6098 GND.n6097 9.3005
R21896 GND.n6099 GND.n4007 9.3005
R21897 GND.n6339 GND.n6100 9.3005
R21898 GND.n6338 GND.n6101 9.3005
R21899 GND.n6337 GND.n6102 9.3005
R21900 GND.n6335 GND.n6103 9.3005
R21901 GND.n6334 GND.n6104 9.3005
R21902 GND.n6331 GND.n6105 9.3005
R21903 GND.n6330 GND.n6329 9.3005
R21904 GND.n4664 GND.n4663 9.3005
R21905 GND.n8288 GND.n1320 9.3005
R21906 GND.n8290 GND.n8289 9.3005
R21907 GND.n1316 GND.n1315 9.3005
R21908 GND.n8297 GND.n8296 9.3005
R21909 GND.n8298 GND.n1314 9.3005
R21910 GND.n8300 GND.n8299 9.3005
R21911 GND.n1310 GND.n1309 9.3005
R21912 GND.n8307 GND.n8306 9.3005
R21913 GND.n8308 GND.n1308 9.3005
R21914 GND.n8310 GND.n8309 9.3005
R21915 GND.n1304 GND.n1303 9.3005
R21916 GND.n8317 GND.n8316 9.3005
R21917 GND.n8318 GND.n1302 9.3005
R21918 GND.n8320 GND.n8319 9.3005
R21919 GND.n1298 GND.n1297 9.3005
R21920 GND.n8327 GND.n8326 9.3005
R21921 GND.n8328 GND.n1296 9.3005
R21922 GND.n8330 GND.n8329 9.3005
R21923 GND.n1292 GND.n1291 9.3005
R21924 GND.n8337 GND.n8336 9.3005
R21925 GND.n8338 GND.n1290 9.3005
R21926 GND.n8340 GND.n8339 9.3005
R21927 GND.n1286 GND.n1285 9.3005
R21928 GND.n8347 GND.n8346 9.3005
R21929 GND.n8348 GND.n1284 9.3005
R21930 GND.n8350 GND.n8349 9.3005
R21931 GND.n1280 GND.n1279 9.3005
R21932 GND.n8357 GND.n8356 9.3005
R21933 GND.n8358 GND.n1278 9.3005
R21934 GND.n8360 GND.n8359 9.3005
R21935 GND.n1274 GND.n1273 9.3005
R21936 GND.n8367 GND.n8366 9.3005
R21937 GND.n8368 GND.n1272 9.3005
R21938 GND.n8370 GND.n8369 9.3005
R21939 GND.n1268 GND.n1267 9.3005
R21940 GND.n8377 GND.n8376 9.3005
R21941 GND.n8378 GND.n1266 9.3005
R21942 GND.n8380 GND.n8379 9.3005
R21943 GND.n1262 GND.n1261 9.3005
R21944 GND.n8387 GND.n8386 9.3005
R21945 GND.n8388 GND.n1260 9.3005
R21946 GND.n8390 GND.n8389 9.3005
R21947 GND.n1256 GND.n1255 9.3005
R21948 GND.n8397 GND.n8396 9.3005
R21949 GND.n8398 GND.n1254 9.3005
R21950 GND.n8400 GND.n8399 9.3005
R21951 GND.n1250 GND.n1249 9.3005
R21952 GND.n8407 GND.n8406 9.3005
R21953 GND.n8408 GND.n1248 9.3005
R21954 GND.n8410 GND.n8409 9.3005
R21955 GND.n1244 GND.n1243 9.3005
R21956 GND.n8417 GND.n8416 9.3005
R21957 GND.n8418 GND.n1242 9.3005
R21958 GND.n8420 GND.n8419 9.3005
R21959 GND.n1238 GND.n1237 9.3005
R21960 GND.n8427 GND.n8426 9.3005
R21961 GND.n8428 GND.n1236 9.3005
R21962 GND.n8430 GND.n8429 9.3005
R21963 GND.n1232 GND.n1231 9.3005
R21964 GND.n8437 GND.n8436 9.3005
R21965 GND.n8438 GND.n1230 9.3005
R21966 GND.n8440 GND.n8439 9.3005
R21967 GND.n1226 GND.n1225 9.3005
R21968 GND.n8447 GND.n8446 9.3005
R21969 GND.n8448 GND.n1224 9.3005
R21970 GND.n8450 GND.n8449 9.3005
R21971 GND.n1220 GND.n1219 9.3005
R21972 GND.n8457 GND.n8456 9.3005
R21973 GND.n8458 GND.n1218 9.3005
R21974 GND.n8460 GND.n8459 9.3005
R21975 GND.n1214 GND.n1213 9.3005
R21976 GND.n8467 GND.n8466 9.3005
R21977 GND.n8468 GND.n1212 9.3005
R21978 GND.n8470 GND.n8469 9.3005
R21979 GND.n1208 GND.n1207 9.3005
R21980 GND.n8477 GND.n8476 9.3005
R21981 GND.n8478 GND.n1206 9.3005
R21982 GND.n8480 GND.n8479 9.3005
R21983 GND.n1202 GND.n1201 9.3005
R21984 GND.n8487 GND.n8486 9.3005
R21985 GND.n8488 GND.n1200 9.3005
R21986 GND.n8490 GND.n8489 9.3005
R21987 GND.n1196 GND.n1195 9.3005
R21988 GND.n8497 GND.n8496 9.3005
R21989 GND.n8498 GND.n1194 9.3005
R21990 GND.n8500 GND.n8499 9.3005
R21991 GND.n1190 GND.n1189 9.3005
R21992 GND.n8507 GND.n8506 9.3005
R21993 GND.n8508 GND.n1188 9.3005
R21994 GND.n8510 GND.n8509 9.3005
R21995 GND.n1184 GND.n1183 9.3005
R21996 GND.n8517 GND.n8516 9.3005
R21997 GND.n8518 GND.n1182 9.3005
R21998 GND.n8520 GND.n8519 9.3005
R21999 GND.n1178 GND.n1177 9.3005
R22000 GND.n8527 GND.n8526 9.3005
R22001 GND.n8528 GND.n1176 9.3005
R22002 GND.n8530 GND.n8529 9.3005
R22003 GND.n1172 GND.n1171 9.3005
R22004 GND.n8537 GND.n8536 9.3005
R22005 GND.n8538 GND.n1170 9.3005
R22006 GND.n8540 GND.n8539 9.3005
R22007 GND.n1166 GND.n1165 9.3005
R22008 GND.n8547 GND.n8546 9.3005
R22009 GND.n8548 GND.n1164 9.3005
R22010 GND.n8550 GND.n8549 9.3005
R22011 GND.n1160 GND.n1159 9.3005
R22012 GND.n8557 GND.n8556 9.3005
R22013 GND.n8558 GND.n1158 9.3005
R22014 GND.n8560 GND.n8559 9.3005
R22015 GND.n1154 GND.n1153 9.3005
R22016 GND.n8567 GND.n8566 9.3005
R22017 GND.n8568 GND.n1152 9.3005
R22018 GND.n8570 GND.n8569 9.3005
R22019 GND.n1148 GND.n1147 9.3005
R22020 GND.n8577 GND.n8576 9.3005
R22021 GND.n8578 GND.n1146 9.3005
R22022 GND.n8580 GND.n8579 9.3005
R22023 GND.n1142 GND.n1141 9.3005
R22024 GND.n8587 GND.n8586 9.3005
R22025 GND.n8588 GND.n1140 9.3005
R22026 GND.n8590 GND.n8589 9.3005
R22027 GND.n1136 GND.n1135 9.3005
R22028 GND.n8597 GND.n8596 9.3005
R22029 GND.n8598 GND.n1134 9.3005
R22030 GND.n8600 GND.n8599 9.3005
R22031 GND.n1130 GND.n1129 9.3005
R22032 GND.n8607 GND.n8606 9.3005
R22033 GND.n8608 GND.n1128 9.3005
R22034 GND.n8610 GND.n8609 9.3005
R22035 GND.n1124 GND.n1123 9.3005
R22036 GND.n8617 GND.n8616 9.3005
R22037 GND.n8618 GND.n1122 9.3005
R22038 GND.n8620 GND.n8619 9.3005
R22039 GND.n1118 GND.n1117 9.3005
R22040 GND.n8627 GND.n8626 9.3005
R22041 GND.n8628 GND.n1116 9.3005
R22042 GND.n8630 GND.n8629 9.3005
R22043 GND.n1112 GND.n1111 9.3005
R22044 GND.n8637 GND.n8636 9.3005
R22045 GND.n8638 GND.n1110 9.3005
R22046 GND.n8640 GND.n8639 9.3005
R22047 GND.n1106 GND.n1105 9.3005
R22048 GND.n8647 GND.n8646 9.3005
R22049 GND.n8648 GND.n1104 9.3005
R22050 GND.n8650 GND.n8649 9.3005
R22051 GND.n1100 GND.n1099 9.3005
R22052 GND.n8657 GND.n8656 9.3005
R22053 GND.n8658 GND.n1098 9.3005
R22054 GND.n8660 GND.n8659 9.3005
R22055 GND.n1094 GND.n1093 9.3005
R22056 GND.n8667 GND.n8666 9.3005
R22057 GND.n8668 GND.n1092 9.3005
R22058 GND.n8670 GND.n8669 9.3005
R22059 GND.n1088 GND.n1087 9.3005
R22060 GND.n8677 GND.n8676 9.3005
R22061 GND.n8678 GND.n1086 9.3005
R22062 GND.n8680 GND.n8679 9.3005
R22063 GND.n1082 GND.n1081 9.3005
R22064 GND.n8687 GND.n8686 9.3005
R22065 GND.n8688 GND.n1080 9.3005
R22066 GND.n8690 GND.n8689 9.3005
R22067 GND.n1076 GND.n1075 9.3005
R22068 GND.n8697 GND.n8696 9.3005
R22069 GND.n8698 GND.n1074 9.3005
R22070 GND.n8700 GND.n8699 9.3005
R22071 GND.n1070 GND.n1069 9.3005
R22072 GND.n8707 GND.n8706 9.3005
R22073 GND.n8708 GND.n1068 9.3005
R22074 GND.n8710 GND.n8709 9.3005
R22075 GND.n1064 GND.n1063 9.3005
R22076 GND.n8717 GND.n8716 9.3005
R22077 GND.n8718 GND.n1062 9.3005
R22078 GND.n8720 GND.n8719 9.3005
R22079 GND.n1058 GND.n1057 9.3005
R22080 GND.n8727 GND.n8726 9.3005
R22081 GND.n8728 GND.n1056 9.3005
R22082 GND.n8730 GND.n8729 9.3005
R22083 GND.n1052 GND.n1051 9.3005
R22084 GND.n8737 GND.n8736 9.3005
R22085 GND.n8738 GND.n1050 9.3005
R22086 GND.n8740 GND.n8739 9.3005
R22087 GND.n1046 GND.n1045 9.3005
R22088 GND.n8747 GND.n8746 9.3005
R22089 GND.n8748 GND.n1044 9.3005
R22090 GND.n8750 GND.n8749 9.3005
R22091 GND.n1040 GND.n1039 9.3005
R22092 GND.n8757 GND.n8756 9.3005
R22093 GND.n8758 GND.n1038 9.3005
R22094 GND.n8760 GND.n8759 9.3005
R22095 GND.n1034 GND.n1033 9.3005
R22096 GND.n8767 GND.n8766 9.3005
R22097 GND.n8768 GND.n1032 9.3005
R22098 GND.n8770 GND.n8769 9.3005
R22099 GND.n1028 GND.n1027 9.3005
R22100 GND.n8777 GND.n8776 9.3005
R22101 GND.n8778 GND.n1026 9.3005
R22102 GND.n8780 GND.n8779 9.3005
R22103 GND.n1022 GND.n1021 9.3005
R22104 GND.n8787 GND.n8786 9.3005
R22105 GND.n8788 GND.n1020 9.3005
R22106 GND.n8790 GND.n8789 9.3005
R22107 GND.n1016 GND.n1015 9.3005
R22108 GND.n8797 GND.n8796 9.3005
R22109 GND.n8798 GND.n1014 9.3005
R22110 GND.n8800 GND.n8799 9.3005
R22111 GND.n1010 GND.n1009 9.3005
R22112 GND.n8807 GND.n8806 9.3005
R22113 GND.n8808 GND.n1008 9.3005
R22114 GND.n8810 GND.n8809 9.3005
R22115 GND.n1004 GND.n1003 9.3005
R22116 GND.n8817 GND.n8816 9.3005
R22117 GND.n8818 GND.n1002 9.3005
R22118 GND.n8820 GND.n8819 9.3005
R22119 GND.n998 GND.n997 9.3005
R22120 GND.n8827 GND.n8826 9.3005
R22121 GND.n8828 GND.n996 9.3005
R22122 GND.n8830 GND.n8829 9.3005
R22123 GND.n992 GND.n991 9.3005
R22124 GND.n8837 GND.n8836 9.3005
R22125 GND.n8838 GND.n990 9.3005
R22126 GND.n8840 GND.n8839 9.3005
R22127 GND.n986 GND.n985 9.3005
R22128 GND.n8847 GND.n8846 9.3005
R22129 GND.n8848 GND.n984 9.3005
R22130 GND.n8850 GND.n8849 9.3005
R22131 GND.n980 GND.n979 9.3005
R22132 GND.n8857 GND.n8856 9.3005
R22133 GND.n8858 GND.n978 9.3005
R22134 GND.n8860 GND.n8859 9.3005
R22135 GND.n974 GND.n973 9.3005
R22136 GND.n8867 GND.n8866 9.3005
R22137 GND.n8868 GND.n972 9.3005
R22138 GND.n8870 GND.n8869 9.3005
R22139 GND.n968 GND.n967 9.3005
R22140 GND.n8877 GND.n8876 9.3005
R22141 GND.n8878 GND.n966 9.3005
R22142 GND.n8880 GND.n8879 9.3005
R22143 GND.n962 GND.n961 9.3005
R22144 GND.n8887 GND.n8886 9.3005
R22145 GND.n8888 GND.n960 9.3005
R22146 GND.n8890 GND.n8889 9.3005
R22147 GND.n956 GND.n955 9.3005
R22148 GND.n8897 GND.n8896 9.3005
R22149 GND.n8898 GND.n954 9.3005
R22150 GND.n8900 GND.n8899 9.3005
R22151 GND.n950 GND.n949 9.3005
R22152 GND.n8907 GND.n8906 9.3005
R22153 GND.n8908 GND.n948 9.3005
R22154 GND.n8910 GND.n8909 9.3005
R22155 GND.n944 GND.n943 9.3005
R22156 GND.n8917 GND.n8916 9.3005
R22157 GND.n8918 GND.n942 9.3005
R22158 GND.n8920 GND.n8919 9.3005
R22159 GND.n938 GND.n937 9.3005
R22160 GND.n8927 GND.n8926 9.3005
R22161 GND.n8928 GND.n936 9.3005
R22162 GND.n8930 GND.n8929 9.3005
R22163 GND.n932 GND.n931 9.3005
R22164 GND.n8937 GND.n8936 9.3005
R22165 GND.n8938 GND.n930 9.3005
R22166 GND.n8940 GND.n8939 9.3005
R22167 GND.n926 GND.n925 9.3005
R22168 GND.n8947 GND.n8946 9.3005
R22169 GND.n8948 GND.n924 9.3005
R22170 GND.n8950 GND.n8949 9.3005
R22171 GND.n920 GND.n919 9.3005
R22172 GND.n8957 GND.n8956 9.3005
R22173 GND.n8958 GND.n918 9.3005
R22174 GND.n8960 GND.n8959 9.3005
R22175 GND.n914 GND.n913 9.3005
R22176 GND.n8967 GND.n8966 9.3005
R22177 GND.n8968 GND.n912 9.3005
R22178 GND.n8970 GND.n8969 9.3005
R22179 GND.n908 GND.n907 9.3005
R22180 GND.n8977 GND.n8976 9.3005
R22181 GND.n8978 GND.n906 9.3005
R22182 GND.n8980 GND.n8979 9.3005
R22183 GND.n902 GND.n901 9.3005
R22184 GND.n8987 GND.n8986 9.3005
R22185 GND.n8988 GND.n900 9.3005
R22186 GND.n8990 GND.n8989 9.3005
R22187 GND.n896 GND.n895 9.3005
R22188 GND.n8997 GND.n8996 9.3005
R22189 GND.n8998 GND.n894 9.3005
R22190 GND.n9000 GND.n8999 9.3005
R22191 GND.n890 GND.n889 9.3005
R22192 GND.n9007 GND.n9006 9.3005
R22193 GND.n9008 GND.n888 9.3005
R22194 GND.n9010 GND.n9009 9.3005
R22195 GND.n884 GND.n883 9.3005
R22196 GND.n9017 GND.n9016 9.3005
R22197 GND.n9018 GND.n882 9.3005
R22198 GND.n9020 GND.n9019 9.3005
R22199 GND.n878 GND.n877 9.3005
R22200 GND.n9027 GND.n9026 9.3005
R22201 GND.n9028 GND.n876 9.3005
R22202 GND.n9030 GND.n9029 9.3005
R22203 GND.n872 GND.n871 9.3005
R22204 GND.n9037 GND.n9036 9.3005
R22205 GND.n9038 GND.n870 9.3005
R22206 GND.n9040 GND.n9039 9.3005
R22207 GND.n866 GND.n865 9.3005
R22208 GND.n9047 GND.n9046 9.3005
R22209 GND.n9048 GND.n864 9.3005
R22210 GND.n9050 GND.n9049 9.3005
R22211 GND.n860 GND.n859 9.3005
R22212 GND.n9057 GND.n9056 9.3005
R22213 GND.n9058 GND.n858 9.3005
R22214 GND.n9060 GND.n9059 9.3005
R22215 GND.n854 GND.n853 9.3005
R22216 GND.n9067 GND.n9066 9.3005
R22217 GND.n9068 GND.n852 9.3005
R22218 GND.n9070 GND.n9069 9.3005
R22219 GND.n848 GND.n847 9.3005
R22220 GND.n9077 GND.n9076 9.3005
R22221 GND.n9078 GND.n846 9.3005
R22222 GND.n9080 GND.n9079 9.3005
R22223 GND.n842 GND.n841 9.3005
R22224 GND.n9087 GND.n9086 9.3005
R22225 GND.n9088 GND.n840 9.3005
R22226 GND.n9090 GND.n9089 9.3005
R22227 GND.n836 GND.n835 9.3005
R22228 GND.n9097 GND.n9096 9.3005
R22229 GND.n9098 GND.n834 9.3005
R22230 GND.n9100 GND.n9099 9.3005
R22231 GND.n830 GND.n829 9.3005
R22232 GND.n9107 GND.n9106 9.3005
R22233 GND.n9108 GND.n828 9.3005
R22234 GND.n9110 GND.n9109 9.3005
R22235 GND.n824 GND.n823 9.3005
R22236 GND.n9117 GND.n9116 9.3005
R22237 GND.n9118 GND.n822 9.3005
R22238 GND.n9120 GND.n9119 9.3005
R22239 GND.n818 GND.n817 9.3005
R22240 GND.n9127 GND.n9126 9.3005
R22241 GND.n9128 GND.n816 9.3005
R22242 GND.n9130 GND.n9129 9.3005
R22243 GND.n812 GND.n811 9.3005
R22244 GND.n9137 GND.n9136 9.3005
R22245 GND.n9138 GND.n810 9.3005
R22246 GND.n9140 GND.n9139 9.3005
R22247 GND.n806 GND.n805 9.3005
R22248 GND.n9147 GND.n9146 9.3005
R22249 GND.n9148 GND.n804 9.3005
R22250 GND.n9150 GND.n9149 9.3005
R22251 GND.n800 GND.n799 9.3005
R22252 GND.n9157 GND.n9156 9.3005
R22253 GND.n9158 GND.n798 9.3005
R22254 GND.n9160 GND.n9159 9.3005
R22255 GND.n794 GND.n793 9.3005
R22256 GND.n9167 GND.n9166 9.3005
R22257 GND.n9168 GND.n792 9.3005
R22258 GND.n9170 GND.n9169 9.3005
R22259 GND.n788 GND.n787 9.3005
R22260 GND.n9177 GND.n9176 9.3005
R22261 GND.n9178 GND.n786 9.3005
R22262 GND.n9180 GND.n9179 9.3005
R22263 GND.n782 GND.n781 9.3005
R22264 GND.n9187 GND.n9186 9.3005
R22265 GND.n9188 GND.n780 9.3005
R22266 GND.n9190 GND.n9189 9.3005
R22267 GND.n776 GND.n775 9.3005
R22268 GND.n9197 GND.n9196 9.3005
R22269 GND.n9198 GND.n774 9.3005
R22270 GND.n9200 GND.n9199 9.3005
R22271 GND.n770 GND.n769 9.3005
R22272 GND.n9207 GND.n9206 9.3005
R22273 GND.n9208 GND.n768 9.3005
R22274 GND.n9210 GND.n9209 9.3005
R22275 GND.n764 GND.n763 9.3005
R22276 GND.n9217 GND.n9216 9.3005
R22277 GND.n9218 GND.n762 9.3005
R22278 GND.n9220 GND.n9219 9.3005
R22279 GND.n758 GND.n757 9.3005
R22280 GND.n9227 GND.n9226 9.3005
R22281 GND.n9228 GND.n756 9.3005
R22282 GND.n9230 GND.n9229 9.3005
R22283 GND.n752 GND.n751 9.3005
R22284 GND.n9237 GND.n9236 9.3005
R22285 GND.n9238 GND.n750 9.3005
R22286 GND.n9240 GND.n9239 9.3005
R22287 GND.n746 GND.n745 9.3005
R22288 GND.n9247 GND.n9246 9.3005
R22289 GND.n9248 GND.n744 9.3005
R22290 GND.n9250 GND.n9249 9.3005
R22291 GND.n740 GND.n739 9.3005
R22292 GND.n9257 GND.n9256 9.3005
R22293 GND.n9258 GND.n738 9.3005
R22294 GND.n9260 GND.n9259 9.3005
R22295 GND.n734 GND.n733 9.3005
R22296 GND.n9267 GND.n9266 9.3005
R22297 GND.n9268 GND.n732 9.3005
R22298 GND.n9270 GND.n9269 9.3005
R22299 GND.n728 GND.n727 9.3005
R22300 GND.n9277 GND.n9276 9.3005
R22301 GND.n9278 GND.n726 9.3005
R22302 GND.n9280 GND.n9279 9.3005
R22303 GND.n722 GND.n721 9.3005
R22304 GND.n9287 GND.n9286 9.3005
R22305 GND.n9288 GND.n720 9.3005
R22306 GND.n9290 GND.n9289 9.3005
R22307 GND.n716 GND.n715 9.3005
R22308 GND.n9297 GND.n9296 9.3005
R22309 GND.n9298 GND.n714 9.3005
R22310 GND.n9300 GND.n9299 9.3005
R22311 GND.n710 GND.n709 9.3005
R22312 GND.n9307 GND.n9306 9.3005
R22313 GND.n9308 GND.n708 9.3005
R22314 GND.n9310 GND.n9309 9.3005
R22315 GND.n704 GND.n703 9.3005
R22316 GND.n9317 GND.n9316 9.3005
R22317 GND.n9318 GND.n702 9.3005
R22318 GND.n9320 GND.n9319 9.3005
R22319 GND.n9327 GND.n9326 9.3005
R22320 GND.n9328 GND.n696 9.3005
R22321 GND.n9330 GND.n9329 9.3005
R22322 GND.n692 GND.n691 9.3005
R22323 GND.n9337 GND.n9336 9.3005
R22324 GND.n9338 GND.n690 9.3005
R22325 GND.n9340 GND.n9339 9.3005
R22326 GND.n686 GND.n685 9.3005
R22327 GND.n9347 GND.n9346 9.3005
R22328 GND.n9348 GND.n684 9.3005
R22329 GND.n9350 GND.n9349 9.3005
R22330 GND.n680 GND.n679 9.3005
R22331 GND.n9357 GND.n9356 9.3005
R22332 GND.n9358 GND.n678 9.3005
R22333 GND.n9360 GND.n9359 9.3005
R22334 GND.n674 GND.n673 9.3005
R22335 GND.n9367 GND.n9366 9.3005
R22336 GND.n9368 GND.n672 9.3005
R22337 GND.n9370 GND.n9369 9.3005
R22338 GND.n668 GND.n667 9.3005
R22339 GND.n9377 GND.n9376 9.3005
R22340 GND.n9378 GND.n666 9.3005
R22341 GND.n9380 GND.n9379 9.3005
R22342 GND.n662 GND.n661 9.3005
R22343 GND.n9387 GND.n9386 9.3005
R22344 GND.n9388 GND.n660 9.3005
R22345 GND.n9390 GND.n9389 9.3005
R22346 GND.n656 GND.n655 9.3005
R22347 GND.n9397 GND.n9396 9.3005
R22348 GND.n9398 GND.n654 9.3005
R22349 GND.n9400 GND.n9399 9.3005
R22350 GND.n650 GND.n649 9.3005
R22351 GND.n9407 GND.n9406 9.3005
R22352 GND.n9408 GND.n648 9.3005
R22353 GND.n9410 GND.n9409 9.3005
R22354 GND.n644 GND.n643 9.3005
R22355 GND.n9417 GND.n9416 9.3005
R22356 GND.n9418 GND.n642 9.3005
R22357 GND.n9420 GND.n9419 9.3005
R22358 GND.n638 GND.n637 9.3005
R22359 GND.n9427 GND.n9426 9.3005
R22360 GND.n9428 GND.n636 9.3005
R22361 GND.n9430 GND.n9429 9.3005
R22362 GND.n632 GND.n631 9.3005
R22363 GND.n9437 GND.n9436 9.3005
R22364 GND.n9438 GND.n630 9.3005
R22365 GND.n9440 GND.n9439 9.3005
R22366 GND.n626 GND.n625 9.3005
R22367 GND.n9447 GND.n9446 9.3005
R22368 GND.n9448 GND.n624 9.3005
R22369 GND.n9451 GND.n9450 9.3005
R22370 GND.n9449 GND.n620 9.3005
R22371 GND.n9457 GND.n619 9.3005
R22372 GND.n9459 GND.n9458 9.3005
R22373 GND.n698 GND.n697 9.3005
R22374 GND.n6320 GND.n6319 9.3005
R22375 GND.n6318 GND.n6110 9.3005
R22376 GND.n6317 GND.n6316 9.3005
R22377 GND.n6313 GND.n6113 9.3005
R22378 GND.n6312 GND.n6309 9.3005
R22379 GND.n6308 GND.n6114 9.3005
R22380 GND.n6307 GND.n6306 9.3005
R22381 GND.n6303 GND.n6115 9.3005
R22382 GND.n6302 GND.n6299 9.3005
R22383 GND.n6298 GND.n6116 9.3005
R22384 GND.n6297 GND.n6296 9.3005
R22385 GND.n6293 GND.n6117 9.3005
R22386 GND.n6288 GND.n6119 9.3005
R22387 GND.n6287 GND.n6286 9.3005
R22388 GND.n6283 GND.n6262 9.3005
R22389 GND.n6282 GND.n6279 9.3005
R22390 GND.n6278 GND.n6263 9.3005
R22391 GND.n6277 GND.n6276 9.3005
R22392 GND.n6273 GND.n6264 9.3005
R22393 GND.n6272 GND.n6269 9.3005
R22394 GND.n6268 GND.n6265 9.3005
R22395 GND.n6267 GND.n6266 9.3005
R22396 GND.n6321 GND.n6106 9.3005
R22397 GND.n6323 GND.n6322 9.3005
R22398 GND.n7253 GND.n3362 9.3005
R22399 GND.n7252 GND.n3363 9.3005
R22400 GND.n6587 GND.n3364 9.3005
R22401 GND.n6588 GND.n6586 9.3005
R22402 GND.n6592 GND.n6589 9.3005
R22403 GND.n6591 GND.n6590 9.3005
R22404 GND.n3945 GND.n3944 9.3005
R22405 GND.n6612 GND.n6611 9.3005
R22406 GND.n6613 GND.n3943 9.3005
R22407 GND.n6617 GND.n6614 9.3005
R22408 GND.n6616 GND.n6615 9.3005
R22409 GND.n3922 GND.n3921 9.3005
R22410 GND.n6636 GND.n6635 9.3005
R22411 GND.n6637 GND.n3920 9.3005
R22412 GND.n6641 GND.n6638 9.3005
R22413 GND.n6640 GND.n6639 9.3005
R22414 GND.n3899 GND.n3898 9.3005
R22415 GND.n6661 GND.n6660 9.3005
R22416 GND.n6662 GND.n3897 9.3005
R22417 GND.n6666 GND.n6663 9.3005
R22418 GND.n6665 GND.n6664 9.3005
R22419 GND.n3877 GND.n3876 9.3005
R22420 GND.n6686 GND.n6685 9.3005
R22421 GND.n6687 GND.n3875 9.3005
R22422 GND.n6691 GND.n6688 9.3005
R22423 GND.n6690 GND.n6689 9.3005
R22424 GND.n3854 GND.n3853 9.3005
R22425 GND.n6711 GND.n6710 9.3005
R22426 GND.n6712 GND.n3852 9.3005
R22427 GND.n6716 GND.n6713 9.3005
R22428 GND.n6715 GND.n6714 9.3005
R22429 GND.n3831 GND.n3830 9.3005
R22430 GND.n6735 GND.n6734 9.3005
R22431 GND.n6736 GND.n3829 9.3005
R22432 GND.n6740 GND.n6737 9.3005
R22433 GND.n6739 GND.n6738 9.3005
R22434 GND.n3808 GND.n3807 9.3005
R22435 GND.n6760 GND.n6759 9.3005
R22436 GND.n6761 GND.n3806 9.3005
R22437 GND.n6765 GND.n6762 9.3005
R22438 GND.n6764 GND.n6763 9.3005
R22439 GND.n3786 GND.n3785 9.3005
R22440 GND.n6785 GND.n6784 9.3005
R22441 GND.n6786 GND.n3784 9.3005
R22442 GND.n6791 GND.n6787 9.3005
R22443 GND.n6790 GND.n6789 9.3005
R22444 GND.n6788 GND.n3756 9.3005
R22445 GND.n6837 GND.n6836 9.3005
R22446 GND.n3728 GND.n3727 9.3005
R22447 GND.n6895 GND.n6894 9.3005
R22448 GND.n6896 GND.n3726 9.3005
R22449 GND.n6900 GND.n6897 9.3005
R22450 GND.n6899 GND.n6898 9.3005
R22451 GND.n3706 GND.n3705 9.3005
R22452 GND.n6922 GND.n6921 9.3005
R22453 GND.n6923 GND.n3704 9.3005
R22454 GND.n6927 GND.n6924 9.3005
R22455 GND.n6926 GND.n6925 9.3005
R22456 GND.n3685 GND.n3684 9.3005
R22457 GND.n6951 GND.n6950 9.3005
R22458 GND.n6952 GND.n3683 9.3005
R22459 GND.n6956 GND.n6953 9.3005
R22460 GND.n6955 GND.n6954 9.3005
R22461 GND.n3665 GND.n3664 9.3005
R22462 GND.n6978 GND.n6977 9.3005
R22463 GND.n6979 GND.n3663 9.3005
R22464 GND.n6983 GND.n6980 9.3005
R22465 GND.n6982 GND.n6981 9.3005
R22466 GND.n3642 GND.n3641 9.3005
R22467 GND.n7004 GND.n7003 9.3005
R22468 GND.n7005 GND.n3640 9.3005
R22469 GND.n7009 GND.n7006 9.3005
R22470 GND.n7008 GND.n7007 9.3005
R22471 GND.n3620 GND.n3619 9.3005
R22472 GND.n7031 GND.n7030 9.3005
R22473 GND.n7032 GND.n3618 9.3005
R22474 GND.n7036 GND.n7033 9.3005
R22475 GND.n7035 GND.n7034 9.3005
R22476 GND.n3599 GND.n3598 9.3005
R22477 GND.n7059 GND.n7058 9.3005
R22478 GND.n7060 GND.n3597 9.3005
R22479 GND.n7064 GND.n7061 9.3005
R22480 GND.n7063 GND.n7062 9.3005
R22481 GND.n3576 GND.n3575 9.3005
R22482 GND.n7092 GND.n7091 9.3005
R22483 GND.n7093 GND.n3574 9.3005
R22484 GND.n7097 GND.n7094 9.3005
R22485 GND.n7096 GND.n7095 9.3005
R22486 GND.n565 GND.n564 9.3005
R22487 GND.n9509 GND.n9508 9.3005
R22488 GND.n9510 GND.n563 9.3005
R22489 GND.n9514 GND.n9511 9.3005
R22490 GND.n9513 GND.n9512 9.3005
R22491 GND.n483 GND.n482 9.3005
R22492 GND.n9610 GND.n9609 9.3005
R22493 GND.n7254 GND.n3361 9.3005
R22494 GND.n6872 GND.n3744 9.3005
R22495 GND.n6838 GND.n3744 9.3005
R22496 GND.n8104 GND.n8103 9.3005
R22497 GND.n8107 GND.n1499 9.3005
R22498 GND.n8108 GND.n1498 9.3005
R22499 GND.n8111 GND.n1497 9.3005
R22500 GND.n8112 GND.n1496 9.3005
R22501 GND.n8115 GND.n1495 9.3005
R22502 GND.n8116 GND.n1494 9.3005
R22503 GND.n8119 GND.n1493 9.3005
R22504 GND.n8120 GND.n1492 9.3005
R22505 GND.n8123 GND.n1491 9.3005
R22506 GND.n8124 GND.n1490 9.3005
R22507 GND.n8127 GND.n1489 9.3005
R22508 GND.n8128 GND.n1486 9.3005
R22509 GND.n8131 GND.n1485 9.3005
R22510 GND.n8132 GND.n1484 9.3005
R22511 GND.n8135 GND.n1483 9.3005
R22512 GND.n8136 GND.n1482 9.3005
R22513 GND.n8139 GND.n1481 9.3005
R22514 GND.n8140 GND.n1480 9.3005
R22515 GND.n8143 GND.n1479 9.3005
R22516 GND.n8145 GND.n1478 9.3005
R22517 GND.n8146 GND.n1477 9.3005
R22518 GND.n8147 GND.n1476 9.3005
R22519 GND.n8148 GND.n1475 9.3005
R22520 GND.n8102 GND.n1503 9.3005
R22521 GND.n8101 GND.n8100 9.3005
R22522 GND.n1539 GND.n1538 9.3005
R22523 GND.n1540 GND.n1534 9.3005
R22524 GND.n8084 GND.n1541 9.3005
R22525 GND.n8083 GND.n1542 9.3005
R22526 GND.n8082 GND.n1543 9.3005
R22527 GND.n2508 GND.n1544 9.3005
R22528 GND.n2512 GND.n2509 9.3005
R22529 GND.n2511 GND.n2510 9.3005
R22530 GND.n2358 GND.n2357 9.3005
R22531 GND.n2532 GND.n2531 9.3005
R22532 GND.n2533 GND.n2356 9.3005
R22533 GND.n2537 GND.n2534 9.3005
R22534 GND.n2536 GND.n2535 9.3005
R22535 GND.n2335 GND.n2334 9.3005
R22536 GND.n2557 GND.n2556 9.3005
R22537 GND.n2558 GND.n2333 9.3005
R22538 GND.n2562 GND.n2559 9.3005
R22539 GND.n2561 GND.n2560 9.3005
R22540 GND.n2312 GND.n2311 9.3005
R22541 GND.n2581 GND.n2580 9.3005
R22542 GND.n2582 GND.n2310 9.3005
R22543 GND.n2586 GND.n2583 9.3005
R22544 GND.n2585 GND.n2584 9.3005
R22545 GND.n2289 GND.n2288 9.3005
R22546 GND.n2606 GND.n2605 9.3005
R22547 GND.n2607 GND.n2287 9.3005
R22548 GND.n2611 GND.n2608 9.3005
R22549 GND.n2610 GND.n2609 9.3005
R22550 GND.n2267 GND.n2266 9.3005
R22551 GND.n2639 GND.n2638 9.3005
R22552 GND.n2640 GND.n2265 9.3005
R22553 GND.n2642 GND.n2641 9.3005
R22554 GND.n2248 GND.n2247 9.3005
R22555 GND.n2706 GND.n2705 9.3005
R22556 GND.n2707 GND.n2246 9.3005
R22557 GND.n2711 GND.n2708 9.3005
R22558 GND.n2710 GND.n2709 9.3005
R22559 GND.n2225 GND.n2224 9.3005
R22560 GND.n2731 GND.n2730 9.3005
R22561 GND.n2732 GND.n2223 9.3005
R22562 GND.n2736 GND.n2733 9.3005
R22563 GND.n2735 GND.n2734 9.3005
R22564 GND.n2202 GND.n2201 9.3005
R22565 GND.n2755 GND.n2754 9.3005
R22566 GND.n2756 GND.n2200 9.3005
R22567 GND.n2758 GND.n2757 9.3005
R22568 GND.n2113 GND.n2106 9.3005
R22569 GND.n2828 GND.n2825 9.3005
R22570 GND.n2827 GND.n2826 9.3005
R22571 GND.n2084 GND.n2083 9.3005
R22572 GND.n2848 GND.n2847 9.3005
R22573 GND.n2849 GND.n2082 9.3005
R22574 GND.n2853 GND.n2850 9.3005
R22575 GND.n2852 GND.n2851 9.3005
R22576 GND.n2062 GND.n2061 9.3005
R22577 GND.n2873 GND.n2872 9.3005
R22578 GND.n2874 GND.n2060 9.3005
R22579 GND.n2878 GND.n2875 9.3005
R22580 GND.n2877 GND.n2876 9.3005
R22581 GND.n2034 GND.n2033 9.3005
R22582 GND.n7671 GND.n7670 9.3005
R22583 GND.n7672 GND.n2032 9.3005
R22584 GND.n7676 GND.n7673 9.3005
R22585 GND.n7675 GND.n7674 9.3005
R22586 GND.n2011 GND.n2010 9.3005
R22587 GND.n7695 GND.n7694 9.3005
R22588 GND.n7696 GND.n2009 9.3005
R22589 GND.n7700 GND.n7697 9.3005
R22590 GND.n7699 GND.n7698 9.3005
R22591 GND.n1988 GND.n1987 9.3005
R22592 GND.n7720 GND.n7719 9.3005
R22593 GND.n7721 GND.n1986 9.3005
R22594 GND.n7725 GND.n7722 9.3005
R22595 GND.n7724 GND.n7723 9.3005
R22596 GND.n1966 GND.n1965 9.3005
R22597 GND.n7745 GND.n7744 9.3005
R22598 GND.n7746 GND.n1964 9.3005
R22599 GND.n7750 GND.n7747 9.3005
R22600 GND.n7749 GND.n7748 9.3005
R22601 GND.n1943 GND.n1942 9.3005
R22602 GND.n7770 GND.n7769 9.3005
R22603 GND.n7771 GND.n1941 9.3005
R22604 GND.n7775 GND.n7772 9.3005
R22605 GND.n7774 GND.n7773 9.3005
R22606 GND.n1920 GND.n1919 9.3005
R22607 GND.n7794 GND.n7793 9.3005
R22608 GND.n7795 GND.n1918 9.3005
R22609 GND.n7799 GND.n7796 9.3005
R22610 GND.n7798 GND.n7797 9.3005
R22611 GND.n1898 GND.n1897 9.3005
R22612 GND.n7821 GND.n7820 9.3005
R22613 GND.n7822 GND.n1896 9.3005
R22614 GND.n7824 GND.n7823 9.3005
R22615 GND.n1778 GND.n1777 9.3005
R22616 GND.n7922 GND.n7921 9.3005
R22617 GND.n1536 GND.n1535 9.3005
R22618 GND.n2824 GND.n2111 9.3005
R22619 GND.n2824 GND.n2105 9.3005
R22620 GND.n2814 GND.n2107 9.3005
R22621 GND.n2181 GND.n2153 9.3005
R22622 GND.n2180 GND.n2154 9.3005
R22623 GND.n2157 GND.n2155 9.3005
R22624 GND.n2176 GND.n2158 9.3005
R22625 GND.n2175 GND.n2159 9.3005
R22626 GND.n2174 GND.n2160 9.3005
R22627 GND.n2163 GND.n2161 9.3005
R22628 GND.n2170 GND.n2164 9.3005
R22629 GND.n2169 GND.n2165 9.3005
R22630 GND.n2168 GND.n2166 9.3005
R22631 GND.n2044 GND.n2043 9.3005
R22632 GND.n2893 GND.n2892 9.3005
R22633 GND.n2894 GND.n2042 9.3005
R22634 GND.n7661 GND.n2895 9.3005
R22635 GND.n7660 GND.n2896 9.3005
R22636 GND.n7659 GND.n2897 9.3005
R22637 GND.n2900 GND.n2898 9.3005
R22638 GND.n7655 GND.n2901 9.3005
R22639 GND.n7654 GND.n2902 9.3005
R22640 GND.n7653 GND.n2903 9.3005
R22641 GND.n2906 GND.n2904 9.3005
R22642 GND.n7649 GND.n2907 9.3005
R22643 GND.n7648 GND.n2908 9.3005
R22644 GND.n7647 GND.n2909 9.3005
R22645 GND.n2912 GND.n2910 9.3005
R22646 GND.n7643 GND.n2913 9.3005
R22647 GND.n7642 GND.n2914 9.3005
R22648 GND.n7641 GND.n2915 9.3005
R22649 GND.n2918 GND.n2916 9.3005
R22650 GND.n7637 GND.n2919 9.3005
R22651 GND.n7636 GND.n2920 9.3005
R22652 GND.n7635 GND.n2921 9.3005
R22653 GND.n2924 GND.n2922 9.3005
R22654 GND.n7631 GND.n2925 9.3005
R22655 GND.n7630 GND.n2926 9.3005
R22656 GND.n7629 GND.n2927 9.3005
R22657 GND.n2930 GND.n2928 9.3005
R22658 GND.n7625 GND.n2931 9.3005
R22659 GND.n7624 GND.n2932 9.3005
R22660 GND.n7623 GND.n2933 9.3005
R22661 GND.n2936 GND.n2934 9.3005
R22662 GND.n7619 GND.n2937 9.3005
R22663 GND.n7618 GND.n2938 9.3005
R22664 GND.n7617 GND.n2939 9.3005
R22665 GND.n2942 GND.n2940 9.3005
R22666 GND.n7613 GND.n2943 9.3005
R22667 GND.n7612 GND.n2944 9.3005
R22668 GND.n7611 GND.n2945 9.3005
R22669 GND.n2948 GND.n2946 9.3005
R22670 GND.n7607 GND.n2949 9.3005
R22671 GND.n7606 GND.n2950 9.3005
R22672 GND.n7605 GND.n2951 9.3005
R22673 GND.n2957 GND.n2952 9.3005
R22674 GND.n7599 GND.n2958 9.3005
R22675 GND.n7598 GND.n2959 9.3005
R22676 GND.n7597 GND.n2960 9.3005
R22677 GND.n2975 GND.n2961 9.3005
R22678 GND.n7585 GND.n2976 9.3005
R22679 GND.n7584 GND.n2977 9.3005
R22680 GND.n7583 GND.n2978 9.3005
R22681 GND.n2994 GND.n2979 9.3005
R22682 GND.n7571 GND.n2995 9.3005
R22683 GND.n7570 GND.n2996 9.3005
R22684 GND.n7569 GND.n2997 9.3005
R22685 GND.n3015 GND.n2998 9.3005
R22686 GND.n7557 GND.n3016 9.3005
R22687 GND.n7556 GND.n3017 9.3005
R22688 GND.n7555 GND.n3018 9.3005
R22689 GND.n4893 GND.n3019 9.3005
R22690 GND.n4894 GND.n4892 9.3005
R22691 GND.n4904 GND.n4895 9.3005
R22692 GND.n4903 GND.n4896 9.3005
R22693 GND.n4902 GND.n4897 9.3005
R22694 GND.n4899 GND.n4898 9.3005
R22695 GND.n4625 GND.n4624 9.3005
R22696 GND.n4939 GND.n4938 9.3005
R22697 GND.n4940 GND.n4623 9.3005
R22698 GND.n4944 GND.n4941 9.3005
R22699 GND.n4943 GND.n4942 9.3005
R22700 GND.n4596 GND.n4595 9.3005
R22701 GND.n4993 GND.n4992 9.3005
R22702 GND.n4994 GND.n4594 9.3005
R22703 GND.n4998 GND.n4995 9.3005
R22704 GND.n4997 GND.n4996 9.3005
R22705 GND.n4573 GND.n4572 9.3005
R22706 GND.n5053 GND.n5052 9.3005
R22707 GND.n5054 GND.n4571 9.3005
R22708 GND.n5067 GND.n5055 9.3005
R22709 GND.n5066 GND.n5056 9.3005
R22710 GND.n5065 GND.n5057 9.3005
R22711 GND.n5059 GND.n5058 9.3005
R22712 GND.n5061 GND.n5060 9.3005
R22713 GND.n4534 GND.n4533 9.3005
R22714 GND.n5111 GND.n5110 9.3005
R22715 GND.n5112 GND.n4532 9.3005
R22716 GND.n5114 GND.n5113 9.3005
R22717 GND.n4508 GND.n4507 9.3005
R22718 GND.n5156 GND.n5155 9.3005
R22719 GND.n5157 GND.n4506 9.3005
R22720 GND.n5161 GND.n5158 9.3005
R22721 GND.n5160 GND.n5159 9.3005
R22722 GND.n4488 GND.n4487 9.3005
R22723 GND.n5216 GND.n5215 9.3005
R22724 GND.n5217 GND.n4486 9.3005
R22725 GND.n5227 GND.n5218 9.3005
R22726 GND.n5226 GND.n5219 9.3005
R22727 GND.n5225 GND.n5220 9.3005
R22728 GND.n5222 GND.n5221 9.3005
R22729 GND.n4453 GND.n4452 9.3005
R22730 GND.n5262 GND.n5261 9.3005
R22731 GND.n5263 GND.n4451 9.3005
R22732 GND.n5267 GND.n5264 9.3005
R22733 GND.n5266 GND.n5265 9.3005
R22734 GND.n4425 GND.n4424 9.3005
R22735 GND.n5317 GND.n5316 9.3005
R22736 GND.n5318 GND.n4423 9.3005
R22737 GND.n5322 GND.n5319 9.3005
R22738 GND.n5321 GND.n5320 9.3005
R22739 GND.n4402 GND.n4401 9.3005
R22740 GND.n5378 GND.n5377 9.3005
R22741 GND.n5379 GND.n4400 9.3005
R22742 GND.n5389 GND.n5380 9.3005
R22743 GND.n5388 GND.n5381 9.3005
R22744 GND.n5387 GND.n5382 9.3005
R22745 GND.n5384 GND.n5383 9.3005
R22746 GND.n4367 GND.n4366 9.3005
R22747 GND.n5424 GND.n5423 9.3005
R22748 GND.n5425 GND.n4365 9.3005
R22749 GND.n5429 GND.n5426 9.3005
R22750 GND.n5428 GND.n5427 9.3005
R22751 GND.n4338 GND.n4337 9.3005
R22752 GND.n5477 GND.n5476 9.3005
R22753 GND.n5478 GND.n4336 9.3005
R22754 GND.n5482 GND.n5479 9.3005
R22755 GND.n5481 GND.n5480 9.3005
R22756 GND.n4315 GND.n4314 9.3005
R22757 GND.n5549 GND.n5548 9.3005
R22758 GND.n5550 GND.n4313 9.3005
R22759 GND.n5560 GND.n5551 9.3005
R22760 GND.n5559 GND.n5552 9.3005
R22761 GND.n5558 GND.n5553 9.3005
R22762 GND.n5555 GND.n5554 9.3005
R22763 GND.n4282 GND.n4281 9.3005
R22764 GND.n5595 GND.n5594 9.3005
R22765 GND.n5596 GND.n4280 9.3005
R22766 GND.n5600 GND.n5597 9.3005
R22767 GND.n5599 GND.n5598 9.3005
R22768 GND.n4254 GND.n4253 9.3005
R22769 GND.n5633 GND.n5632 9.3005
R22770 GND.n5634 GND.n4252 9.3005
R22771 GND.n5636 GND.n5635 9.3005
R22772 GND.n4230 GND.n4229 9.3005
R22773 GND.n5689 GND.n5688 9.3005
R22774 GND.n5690 GND.n4228 9.3005
R22775 GND.n5694 GND.n5691 9.3005
R22776 GND.n5693 GND.n5692 9.3005
R22777 GND.n4207 GND.n4206 9.3005
R22778 GND.n5723 GND.n5722 9.3005
R22779 GND.n5724 GND.n4205 9.3005
R22780 GND.n5728 GND.n5725 9.3005
R22781 GND.n5727 GND.n5726 9.3005
R22782 GND.n4184 GND.n4183 9.3005
R22783 GND.n5804 GND.n5803 9.3005
R22784 GND.n5805 GND.n4182 9.3005
R22785 GND.n5818 GND.n5806 9.3005
R22786 GND.n5817 GND.n5807 9.3005
R22787 GND.n5816 GND.n5808 9.3005
R22788 GND.n5810 GND.n5809 9.3005
R22789 GND.n5812 GND.n5811 9.3005
R22790 GND.n4147 GND.n4146 9.3005
R22791 GND.n5864 GND.n5863 9.3005
R22792 GND.n5865 GND.n4145 9.3005
R22793 GND.n5875 GND.n5866 9.3005
R22794 GND.n5874 GND.n5867 9.3005
R22795 GND.n5873 GND.n5868 9.3005
R22796 GND.n5870 GND.n5869 9.3005
R22797 GND.n4112 GND.n4111 9.3005
R22798 GND.n5910 GND.n5909 9.3005
R22799 GND.n5911 GND.n4110 9.3005
R22800 GND.n5915 GND.n5912 9.3005
R22801 GND.n5914 GND.n5913 9.3005
R22802 GND.n4083 GND.n4082 9.3005
R22803 GND.n5963 GND.n5962 9.3005
R22804 GND.n5964 GND.n4081 9.3005
R22805 GND.n5968 GND.n5965 9.3005
R22806 GND.n5967 GND.n5966 9.3005
R22807 GND.n4059 GND.n4058 9.3005
R22808 GND.n6012 GND.n6011 9.3005
R22809 GND.n6013 GND.n4057 9.3005
R22810 GND.n6026 GND.n6014 9.3005
R22811 GND.n6025 GND.n6015 9.3005
R22812 GND.n6024 GND.n6016 9.3005
R22813 GND.n6018 GND.n6017 9.3005
R22814 GND.n6020 GND.n6019 9.3005
R22815 GND.n4018 GND.n4017 9.3005
R22816 GND.n6088 GND.n6087 9.3005
R22817 GND.n6089 GND.n4016 9.3005
R22818 GND.n6093 GND.n6090 9.3005
R22819 GND.n6092 GND.n6091 9.3005
R22820 GND.n3996 GND.n3995 9.3005
R22821 GND.n6353 GND.n6352 9.3005
R22822 GND.n6354 GND.n3994 9.3005
R22823 GND.n6359 GND.n6355 9.3005
R22824 GND.n6358 GND.n6357 9.3005
R22825 GND.n6356 GND.n3235 9.3005
R22826 GND.n7339 GND.n3236 9.3005
R22827 GND.n7338 GND.n3237 9.3005
R22828 GND.n7337 GND.n3238 9.3005
R22829 GND.n3252 GND.n3239 9.3005
R22830 GND.n7325 GND.n3253 9.3005
R22831 GND.n7324 GND.n3254 9.3005
R22832 GND.n7323 GND.n3255 9.3005
R22833 GND.n3277 GND.n3256 9.3005
R22834 GND.n3278 GND.n3276 9.3005
R22835 GND.n7306 GND.n3279 9.3005
R22836 GND.n7305 GND.n3280 9.3005
R22837 GND.n7304 GND.n3281 9.3005
R22838 GND.n3286 GND.n3282 9.3005
R22839 GND.n7298 GND.n3287 9.3005
R22840 GND.n7297 GND.n3288 9.3005
R22841 GND.n7296 GND.n3289 9.3005
R22842 GND.n6443 GND.n3290 9.3005
R22843 GND.n6445 GND.n6444 9.3005
R22844 GND.n6442 GND.n6441 9.3005
R22845 GND.n6450 GND.n6449 9.3005
R22846 GND.n6451 GND.n6440 9.3005
R22847 GND.n6578 GND.n6452 9.3005
R22848 GND.n6577 GND.n6453 9.3005
R22849 GND.n6576 GND.n6454 9.3005
R22850 GND.n6457 GND.n6455 9.3005
R22851 GND.n6572 GND.n6458 9.3005
R22852 GND.n6571 GND.n6459 9.3005
R22853 GND.n6570 GND.n6460 9.3005
R22854 GND.n6463 GND.n6461 9.3005
R22855 GND.n6566 GND.n6464 9.3005
R22856 GND.n6565 GND.n6465 9.3005
R22857 GND.n6564 GND.n6466 9.3005
R22858 GND.n6469 GND.n6467 9.3005
R22859 GND.n6560 GND.n6470 9.3005
R22860 GND.n6559 GND.n6471 9.3005
R22861 GND.n6558 GND.n6472 9.3005
R22862 GND.n6475 GND.n6473 9.3005
R22863 GND.n6554 GND.n6476 9.3005
R22864 GND.n6553 GND.n6477 9.3005
R22865 GND.n6552 GND.n6478 9.3005
R22866 GND.n6481 GND.n6479 9.3005
R22867 GND.n6548 GND.n6482 9.3005
R22868 GND.n6547 GND.n6483 9.3005
R22869 GND.n6546 GND.n6484 9.3005
R22870 GND.n6487 GND.n6485 9.3005
R22871 GND.n6542 GND.n6488 9.3005
R22872 GND.n6541 GND.n6489 9.3005
R22873 GND.n6540 GND.n6490 9.3005
R22874 GND.n6493 GND.n6491 9.3005
R22875 GND.n6536 GND.n6494 9.3005
R22876 GND.n6535 GND.n6495 9.3005
R22877 GND.n6534 GND.n6496 9.3005
R22878 GND.n6499 GND.n6497 9.3005
R22879 GND.n6530 GND.n6500 9.3005
R22880 GND.n6529 GND.n6501 9.3005
R22881 GND.n6528 GND.n6502 9.3005
R22882 GND.n6505 GND.n6503 9.3005
R22883 GND.n6524 GND.n6506 9.3005
R22884 GND.n6523 GND.n6507 9.3005
R22885 GND.n6522 GND.n6508 9.3005
R22886 GND.n6511 GND.n6509 9.3005
R22887 GND.n6518 GND.n6512 9.3005
R22888 GND.n6517 GND.n6513 9.3005
R22889 GND.n6516 GND.n6514 9.3005
R22890 GND.n3746 GND.n3745 9.3005
R22891 GND.n6881 GND.n6880 9.3005
R22892 GND.n6885 GND.n6882 9.3005
R22893 GND.n6884 GND.n6883 9.3005
R22894 GND.n3718 GND.n3717 9.3005
R22895 GND.n6906 GND.n6905 9.3005
R22896 GND.n6907 GND.n3716 9.3005
R22897 GND.n6911 GND.n6908 9.3005
R22898 GND.n6910 GND.n6909 9.3005
R22899 GND.n3696 GND.n3695 9.3005
R22900 GND.n6933 GND.n6932 9.3005
R22901 GND.n6934 GND.n3694 9.3005
R22902 GND.n6938 GND.n6935 9.3005
R22903 GND.n6937 GND.n6936 9.3005
R22904 GND.n3676 GND.n3675 9.3005
R22905 GND.n6962 GND.n6961 9.3005
R22906 GND.n6963 GND.n3674 9.3005
R22907 GND.n6967 GND.n6964 9.3005
R22908 GND.n6966 GND.n6965 9.3005
R22909 GND.n3654 GND.n3653 9.3005
R22910 GND.n6989 GND.n6988 9.3005
R22911 GND.n6990 GND.n3652 9.3005
R22912 GND.n6994 GND.n6991 9.3005
R22913 GND.n6993 GND.n6992 9.3005
R22914 GND.n3632 GND.n3631 9.3005
R22915 GND.n7015 GND.n7014 9.3005
R22916 GND.n7016 GND.n3630 9.3005
R22917 GND.n7020 GND.n7017 9.3005
R22918 GND.n7019 GND.n7018 9.3005
R22919 GND.n3610 GND.n3609 9.3005
R22920 GND.n7042 GND.n7041 9.3005
R22921 GND.n7043 GND.n3608 9.3005
R22922 GND.n7047 GND.n7044 9.3005
R22923 GND.n7046 GND.n7045 9.3005
R22924 GND.n3589 GND.n3588 9.3005
R22925 GND.n7070 GND.n7069 9.3005
R22926 GND.n7071 GND.n3587 9.3005
R22927 GND.n7082 GND.n7072 9.3005
R22928 GND.n7081 GND.n7073 9.3005
R22929 GND.n7080 GND.n7074 9.3005
R22930 GND.n7077 GND.n7076 9.3005
R22931 GND.n7075 GND.n582 9.3005
R22932 GND.n9497 GND.n583 9.3005
R22933 GND.n9496 GND.n584 9.3005
R22934 GND.n9495 GND.n585 9.3005
R22935 GND.n588 GND.n586 9.3005
R22936 GND.n9491 GND.n589 9.3005
R22937 GND.n9490 GND.n590 9.3005
R22938 GND.n9489 GND.n591 9.3005
R22939 GND.n594 GND.n592 9.3005
R22940 GND.n9485 GND.n595 9.3005
R22941 GND.n9484 GND.n596 9.3005
R22942 GND.n9483 GND.n597 9.3005
R22943 GND.n602 GND.n598 9.3005
R22944 GND.n9477 GND.n603 9.3005
R22945 GND.n9476 GND.n604 9.3005
R22946 GND.n9475 GND.n605 9.3005
R22947 GND.n610 GND.n606 9.3005
R22948 GND.n9469 GND.n611 9.3005
R22949 GND.n9468 GND.n612 9.3005
R22950 GND.n9467 GND.n613 9.3005
R22951 GND.n618 GND.n614 9.3005
R22952 GND.n9461 GND.n9460 9.3005
R22953 GND.n8172 GND.n1430 9.3005
R22954 GND.n8171 GND.n1432 9.3005
R22955 GND.n1438 GND.n1433 9.3005
R22956 GND.n8165 GND.n1439 9.3005
R22957 GND.n8164 GND.n1440 9.3005
R22958 GND.n8163 GND.n1441 9.3005
R22959 GND.n1446 GND.n1442 9.3005
R22960 GND.n8157 GND.n1447 9.3005
R22961 GND.n8156 GND.n1448 9.3005
R22962 GND.n8155 GND.n1449 9.3005
R22963 GND.n1516 GND.n1450 9.3005
R22964 GND.n1519 GND.n1518 9.3005
R22965 GND.n1520 GND.n1515 9.3005
R22966 GND.n8091 GND.n1521 9.3005
R22967 GND.n8090 GND.n1522 9.3005
R22968 GND.n8089 GND.n1523 9.3005
R22969 GND.n2427 GND.n1524 9.3005
R22970 GND.n2429 GND.n2428 9.3005
R22971 GND.n2433 GND.n2432 9.3005
R22972 GND.n2434 GND.n2426 9.3005
R22973 GND.n2501 GND.n2435 9.3005
R22974 GND.n2500 GND.n2436 9.3005
R22975 GND.n2499 GND.n2437 9.3005
R22976 GND.n2440 GND.n2438 9.3005
R22977 GND.n2495 GND.n2441 9.3005
R22978 GND.n2494 GND.n2442 9.3005
R22979 GND.n2493 GND.n2443 9.3005
R22980 GND.n2446 GND.n2444 9.3005
R22981 GND.n2489 GND.n2447 9.3005
R22982 GND.n2488 GND.n2448 9.3005
R22983 GND.n2487 GND.n2449 9.3005
R22984 GND.n2452 GND.n2450 9.3005
R22985 GND.n2483 GND.n2453 9.3005
R22986 GND.n2482 GND.n2454 9.3005
R22987 GND.n2481 GND.n2455 9.3005
R22988 GND.n2458 GND.n2456 9.3005
R22989 GND.n2477 GND.n2459 9.3005
R22990 GND.n2476 GND.n2460 9.3005
R22991 GND.n2475 GND.n2461 9.3005
R22992 GND.n2464 GND.n2462 9.3005
R22993 GND.n2471 GND.n2465 9.3005
R22994 GND.n2470 GND.n2466 9.3005
R22995 GND.n2469 GND.n2467 9.3005
R22996 GND.n2259 GND.n2258 9.3005
R22997 GND.n2648 GND.n2647 9.3005
R22998 GND.n2649 GND.n2257 9.3005
R22999 GND.n2694 GND.n2650 9.3005
R23000 GND.n2693 GND.n2651 9.3005
R23001 GND.n2692 GND.n2652 9.3005
R23002 GND.n2655 GND.n2653 9.3005
R23003 GND.n2688 GND.n2656 9.3005
R23004 GND.n2687 GND.n2657 9.3005
R23005 GND.n2686 GND.n2658 9.3005
R23006 GND.n2661 GND.n2659 9.3005
R23007 GND.n2682 GND.n2662 9.3005
R23008 GND.n2681 GND.n2663 9.3005
R23009 GND.n2680 GND.n2664 9.3005
R23010 GND.n2669 GND.n2665 9.3005
R23011 GND.n2676 GND.n2670 9.3005
R23012 GND.n2675 GND.n2671 9.3005
R23013 GND.n8174 GND.n8173 9.3005
R23014 GND.n1429 GND.n1425 9.3005
R23015 GND.n8182 GND.n1424 9.3005
R23016 GND.n8183 GND.n1423 9.3005
R23017 GND.n8184 GND.n1422 9.3005
R23018 GND.n1421 GND.n1417 9.3005
R23019 GND.n8190 GND.n1416 9.3005
R23020 GND.n8191 GND.n1415 9.3005
R23021 GND.n8192 GND.n1414 9.3005
R23022 GND.n1413 GND.n1409 9.3005
R23023 GND.n8198 GND.n1408 9.3005
R23024 GND.n8199 GND.n1407 9.3005
R23025 GND.n8200 GND.n1406 9.3005
R23026 GND.n1405 GND.n1401 9.3005
R23027 GND.n8206 GND.n1400 9.3005
R23028 GND.n8207 GND.n1399 9.3005
R23029 GND.n8208 GND.n1398 9.3005
R23030 GND.n1397 GND.n1393 9.3005
R23031 GND.n8214 GND.n1392 9.3005
R23032 GND.n8215 GND.n1391 9.3005
R23033 GND.n8216 GND.n1390 9.3005
R23034 GND.n1389 GND.n1385 9.3005
R23035 GND.n8222 GND.n1384 9.3005
R23036 GND.n8223 GND.n1383 9.3005
R23037 GND.n8224 GND.n1382 9.3005
R23038 GND.n1381 GND.n1377 9.3005
R23039 GND.n8230 GND.n1376 9.3005
R23040 GND.n8231 GND.n1375 9.3005
R23041 GND.n8232 GND.n1374 9.3005
R23042 GND.n1373 GND.n1369 9.3005
R23043 GND.n8238 GND.n1368 9.3005
R23044 GND.n8239 GND.n1367 9.3005
R23045 GND.n8240 GND.n1366 9.3005
R23046 GND.n1365 GND.n1361 9.3005
R23047 GND.n8246 GND.n1360 9.3005
R23048 GND.n8247 GND.n1359 9.3005
R23049 GND.n8248 GND.n1358 9.3005
R23050 GND.n1357 GND.n1353 9.3005
R23051 GND.n8254 GND.n1352 9.3005
R23052 GND.n8255 GND.n1351 9.3005
R23053 GND.n8256 GND.n1350 9.3005
R23054 GND.n1349 GND.n1345 9.3005
R23055 GND.n8262 GND.n1344 9.3005
R23056 GND.n8263 GND.n1343 9.3005
R23057 GND.n8264 GND.n1342 9.3005
R23058 GND.n1341 GND.n1337 9.3005
R23059 GND.n8270 GND.n1336 9.3005
R23060 GND.n8271 GND.n1335 9.3005
R23061 GND.n8272 GND.n1334 9.3005
R23062 GND.n1333 GND.n1329 9.3005
R23063 GND.n8278 GND.n1328 9.3005
R23064 GND.n8279 GND.n1327 9.3005
R23065 GND.n8280 GND.n1326 9.3005
R23066 GND.n1322 GND.n1321 9.3005
R23067 GND.n8287 GND.n8286 9.3005
R23068 GND.n8176 GND.n8175 9.3005
R23069 GND.n6432 GND.n6431 9.3005
R23070 GND.n6433 GND.n3962 9.3005
R23071 GND.n6435 GND.n6434 9.3005
R23072 GND.n3956 GND.n3955 9.3005
R23073 GND.n6597 GND.n6596 9.3005
R23074 GND.n6598 GND.n3953 9.3005
R23075 GND.n6601 GND.n6600 9.3005
R23076 GND.n6599 GND.n3954 9.3005
R23077 GND.n3935 GND.n3934 9.3005
R23078 GND.n6622 GND.n6621 9.3005
R23079 GND.n6623 GND.n3932 9.3005
R23080 GND.n6626 GND.n6625 9.3005
R23081 GND.n6624 GND.n3933 9.3005
R23082 GND.n3911 GND.n3910 9.3005
R23083 GND.n6646 GND.n6645 9.3005
R23084 GND.n6647 GND.n3908 9.3005
R23085 GND.n6650 GND.n6649 9.3005
R23086 GND.n6648 GND.n3909 9.3005
R23087 GND.n3888 GND.n3887 9.3005
R23088 GND.n6671 GND.n6670 9.3005
R23089 GND.n6672 GND.n3885 9.3005
R23090 GND.n6675 GND.n6674 9.3005
R23091 GND.n6673 GND.n3886 9.3005
R23092 GND.n3866 GND.n3865 9.3005
R23093 GND.n6696 GND.n6695 9.3005
R23094 GND.n6697 GND.n3863 9.3005
R23095 GND.n6700 GND.n6699 9.3005
R23096 GND.n6698 GND.n3864 9.3005
R23097 GND.n3844 GND.n3843 9.3005
R23098 GND.n6721 GND.n6720 9.3005
R23099 GND.n6722 GND.n3841 9.3005
R23100 GND.n6725 GND.n6724 9.3005
R23101 GND.n6723 GND.n3842 9.3005
R23102 GND.n3820 GND.n3819 9.3005
R23103 GND.n6745 GND.n6744 9.3005
R23104 GND.n6746 GND.n3817 9.3005
R23105 GND.n6749 GND.n6748 9.3005
R23106 GND.n6747 GND.n3818 9.3005
R23107 GND.n3797 GND.n3796 9.3005
R23108 GND.n6770 GND.n6769 9.3005
R23109 GND.n6771 GND.n3794 9.3005
R23110 GND.n6774 GND.n6773 9.3005
R23111 GND.n6772 GND.n3795 9.3005
R23112 GND.n3770 GND.n3769 9.3005
R23113 GND.n6796 GND.n6795 9.3005
R23114 GND.n6797 GND.n3767 9.3005
R23115 GND.n6799 GND.n6798 9.3005
R23116 GND.n6800 GND.n3766 9.3005
R23117 GND.n6805 GND.n6804 9.3005
R23118 GND.n6806 GND.n3765 9.3005
R23119 GND.n6808 GND.n6807 9.3005
R23120 GND.n408 GND.n406 9.3005
R23121 GND.n6430 GND.n3355 9.3005
R23122 GND.n9693 GND.n9692 9.3005
R23123 GND.n9691 GND.n407 9.3005
R23124 GND.n9690 GND.n9689 9.3005
R23125 GND.n9688 GND.n412 9.3005
R23126 GND.n9687 GND.n9686 9.3005
R23127 GND.n9685 GND.n413 9.3005
R23128 GND.n9684 GND.n9683 9.3005
R23129 GND.n9682 GND.n417 9.3005
R23130 GND.n9681 GND.n9680 9.3005
R23131 GND.n9679 GND.n418 9.3005
R23132 GND.n9678 GND.n9677 9.3005
R23133 GND.n9676 GND.n422 9.3005
R23134 GND.n9675 GND.n9674 9.3005
R23135 GND.n9673 GND.n423 9.3005
R23136 GND.n9672 GND.n9671 9.3005
R23137 GND.n9670 GND.n427 9.3005
R23138 GND.n9669 GND.n9668 9.3005
R23139 GND.n9667 GND.n428 9.3005
R23140 GND.n9666 GND.n9665 9.3005
R23141 GND.n9664 GND.n432 9.3005
R23142 GND.n9663 GND.n9662 9.3005
R23143 GND.n9661 GND.n433 9.3005
R23144 GND.n9660 GND.n9659 9.3005
R23145 GND.n9658 GND.n437 9.3005
R23146 GND.n9657 GND.n9656 9.3005
R23147 GND.n9655 GND.n438 9.3005
R23148 GND.n9654 GND.n9653 9.3005
R23149 GND.n9652 GND.n442 9.3005
R23150 GND.n9651 GND.n9650 9.3005
R23151 GND.n9649 GND.n443 9.3005
R23152 GND.n9648 GND.n9647 9.3005
R23153 GND.n9646 GND.n447 9.3005
R23154 GND.n9645 GND.n9644 9.3005
R23155 GND.n9643 GND.n448 9.3005
R23156 GND.n9642 GND.n9641 9.3005
R23157 GND.n9640 GND.n452 9.3005
R23158 GND.n9639 GND.n9638 9.3005
R23159 GND.n9637 GND.n453 9.3005
R23160 GND.n9636 GND.n9635 9.3005
R23161 GND.n9634 GND.n457 9.3005
R23162 GND.n9633 GND.n9632 9.3005
R23163 GND.n9631 GND.n458 9.3005
R23164 GND.n9630 GND.n9629 9.3005
R23165 GND.n9628 GND.n462 9.3005
R23166 GND.n9627 GND.n9626 9.3005
R23167 GND.n9625 GND.n463 9.3005
R23168 GND.n9624 GND.n9623 9.3005
R23169 GND.n9622 GND.n467 9.3005
R23170 GND.n9621 GND.n9620 9.3005
R23171 GND.n9619 GND.n468 9.3005
R23172 GND.n9618 GND.n9617 9.3005
R23173 GND.n9616 GND.n472 9.3005
R23174 GND.n9615 GND.n9614 9.3005
R23175 GND.n9563 GND.n546 9.3005
R23176 GND.n9562 GND.n9561 9.3005
R23177 GND.n9560 GND.n9530 9.3005
R23178 GND.n9559 GND.n9558 9.3005
R23179 GND.n9557 GND.n9535 9.3005
R23180 GND.n9556 GND.n9555 9.3005
R23181 GND.n9554 GND.n9536 9.3005
R23182 GND.n9553 GND.n9552 9.3005
R23183 GND.n9551 GND.n9541 9.3005
R23184 GND.n9550 GND.n9549 9.3005
R23185 GND.n9548 GND.n9542 9.3005
R23186 GND.n9547 GND.n473 9.3005
R23187 GND.n9565 GND.n9564 9.3005
R23188 GND.n9606 GND.n484 9.3005
R23189 GND.n9605 GND.n9604 9.3005
R23190 GND.n9603 GND.n487 9.3005
R23191 GND.n9602 GND.n9601 9.3005
R23192 GND.n9600 GND.n488 9.3005
R23193 GND.n9599 GND.n9598 9.3005
R23194 GND.n9597 GND.n492 9.3005
R23195 GND.n9596 GND.n9595 9.3005
R23196 GND.n9594 GND.n493 9.3005
R23197 GND.n9593 GND.n9592 9.3005
R23198 GND.n9591 GND.n499 9.3005
R23199 GND.n9590 GND.n9589 9.3005
R23200 GND.n9588 GND.n500 9.3005
R23201 GND.n9587 GND.n9586 9.3005
R23202 GND.n9585 GND.n504 9.3005
R23203 GND.n9584 GND.n9583 9.3005
R23204 GND.n9582 GND.n505 9.3005
R23205 GND.n9581 GND.n9580 9.3005
R23206 GND.n9579 GND.n509 9.3005
R23207 GND.n9578 GND.n9577 9.3005
R23208 GND.n9576 GND.n510 9.3005
R23209 GND.n9575 GND.n9574 9.3005
R23210 GND.n9573 GND.n514 9.3005
R23211 GND.n9572 GND.n9571 9.3005
R23212 GND.n9570 GND.n515 9.3005
R23213 GND.n9608 GND.n9607 9.3005
R23214 GND.n3374 GND.n3372 9.3005
R23215 GND.n7248 GND.n7247 9.3005
R23216 GND.n3375 GND.n3373 9.3005
R23217 GND.n7243 GND.n3382 9.3005
R23218 GND.n7242 GND.n3383 9.3005
R23219 GND.n7241 GND.n3384 9.3005
R23220 GND.n3951 GND.n3385 9.3005
R23221 GND.n7237 GND.n3390 9.3005
R23222 GND.n7236 GND.n3391 9.3005
R23223 GND.n7235 GND.n3392 9.3005
R23224 GND.n3928 GND.n3393 9.3005
R23225 GND.n7231 GND.n3398 9.3005
R23226 GND.n7230 GND.n3399 9.3005
R23227 GND.n7229 GND.n3400 9.3005
R23228 GND.n3915 GND.n3401 9.3005
R23229 GND.n7225 GND.n3406 9.3005
R23230 GND.n7224 GND.n3407 9.3005
R23231 GND.n7223 GND.n3408 9.3005
R23232 GND.n6654 GND.n3409 9.3005
R23233 GND.n7219 GND.n3414 9.3005
R23234 GND.n7218 GND.n3415 9.3005
R23235 GND.n7217 GND.n3416 9.3005
R23236 GND.n6681 GND.n3417 9.3005
R23237 GND.n7213 GND.n3422 9.3005
R23238 GND.n7212 GND.n3423 9.3005
R23239 GND.n7211 GND.n3424 9.3005
R23240 GND.n3860 GND.n3425 9.3005
R23241 GND.n7207 GND.n3430 9.3005
R23242 GND.n7206 GND.n3431 9.3005
R23243 GND.n7205 GND.n3432 9.3005
R23244 GND.n3837 GND.n3433 9.3005
R23245 GND.n7201 GND.n3438 9.3005
R23246 GND.n7200 GND.n3439 9.3005
R23247 GND.n7199 GND.n3440 9.3005
R23248 GND.n3824 GND.n3441 9.3005
R23249 GND.n7195 GND.n3446 9.3005
R23250 GND.n7194 GND.n3447 9.3005
R23251 GND.n7193 GND.n3448 9.3005
R23252 GND.n6753 GND.n3449 9.3005
R23253 GND.n7189 GND.n3454 9.3005
R23254 GND.n7188 GND.n3455 9.3005
R23255 GND.n7187 GND.n3456 9.3005
R23256 GND.n6780 GND.n3457 9.3005
R23257 GND.n7183 GND.n3462 9.3005
R23258 GND.n7182 GND.n3463 9.3005
R23259 GND.n7181 GND.n3464 9.3005
R23260 GND.n3779 GND.n3465 9.3005
R23261 GND.n7177 GND.n3470 9.3005
R23262 GND.n7176 GND.n3471 9.3005
R23263 GND.n7175 GND.n3472 9.3005
R23264 GND.n3764 GND.n3473 9.3005
R23265 GND.n7171 GND.n3478 9.3005
R23266 GND.n7170 GND.n3479 9.3005
R23267 GND.n7169 GND.n3480 9.3005
R23268 GND.n6851 GND.n3481 9.3005
R23269 GND.n7165 GND.n3486 9.3005
R23270 GND.n7164 GND.n3487 9.3005
R23271 GND.n7163 GND.n3488 9.3005
R23272 GND.n3734 GND.n3489 9.3005
R23273 GND.n7159 GND.n3494 9.3005
R23274 GND.n7158 GND.n3495 9.3005
R23275 GND.n7157 GND.n3496 9.3005
R23276 GND.n3711 GND.n3497 9.3005
R23277 GND.n7153 GND.n3502 9.3005
R23278 GND.n7152 GND.n3503 9.3005
R23279 GND.n7151 GND.n3504 9.3005
R23280 GND.n3700 GND.n3505 9.3005
R23281 GND.n7147 GND.n3510 9.3005
R23282 GND.n7146 GND.n3511 9.3005
R23283 GND.n7145 GND.n3512 9.3005
R23284 GND.n6944 GND.n3513 9.3005
R23285 GND.n7141 GND.n3518 9.3005
R23286 GND.n7140 GND.n3519 9.3005
R23287 GND.n7139 GND.n3520 9.3005
R23288 GND.n6973 GND.n3521 9.3005
R23289 GND.n7135 GND.n3526 9.3005
R23290 GND.n7134 GND.n3527 9.3005
R23291 GND.n7133 GND.n3528 9.3005
R23292 GND.n3648 GND.n3529 9.3005
R23293 GND.n7129 GND.n3534 9.3005
R23294 GND.n7128 GND.n3535 9.3005
R23295 GND.n7127 GND.n3536 9.3005
R23296 GND.n3625 GND.n3537 9.3005
R23297 GND.n7123 GND.n3542 9.3005
R23298 GND.n7122 GND.n3543 9.3005
R23299 GND.n7121 GND.n3544 9.3005
R23300 GND.n3614 GND.n3545 9.3005
R23301 GND.n7117 GND.n3550 9.3005
R23302 GND.n7116 GND.n3551 9.3005
R23303 GND.n7115 GND.n3552 9.3005
R23304 GND.n7053 GND.n3553 9.3005
R23305 GND.n7111 GND.n3558 9.3005
R23306 GND.n7110 GND.n3559 9.3005
R23307 GND.n7109 GND.n3560 9.3005
R23308 GND.n7087 GND.n3561 9.3005
R23309 GND.n7105 GND.n3566 9.3005
R23310 GND.n7104 GND.n3567 9.3005
R23311 GND.n7103 GND.n7102 9.3005
R23312 GND.n576 GND.n574 9.3005
R23313 GND.n9504 GND.n9503 9.3005
R23314 GND.n575 GND.n554 9.3005
R23315 GND.n9519 GND.n553 9.3005
R23316 GND.n9521 GND.n9520 9.3005
R23317 GND.n9522 GND.n547 9.3005
R23318 GND.n9528 GND.n548 9.3005
R23319 GND.n6326 GND.n6324 9.3005
R23320 GND.n3378 GND.n3374 9.3005
R23321 GND.n7247 GND.n7246 9.3005
R23322 GND.n7245 GND.n3375 9.3005
R23323 GND.n7244 GND.n7243 9.3005
R23324 GND.n7242 GND.n3381 9.3005
R23325 GND.n7241 GND.n7240 9.3005
R23326 GND.n7239 GND.n3385 9.3005
R23327 GND.n7238 GND.n7237 9.3005
R23328 GND.n7236 GND.n3389 9.3005
R23329 GND.n7235 GND.n7234 9.3005
R23330 GND.n7233 GND.n3393 9.3005
R23331 GND.n7232 GND.n7231 9.3005
R23332 GND.n7230 GND.n3397 9.3005
R23333 GND.n7229 GND.n7228 9.3005
R23334 GND.n7227 GND.n3401 9.3005
R23335 GND.n7226 GND.n7225 9.3005
R23336 GND.n7224 GND.n3405 9.3005
R23337 GND.n7223 GND.n7222 9.3005
R23338 GND.n7221 GND.n3409 9.3005
R23339 GND.n7220 GND.n7219 9.3005
R23340 GND.n7218 GND.n3413 9.3005
R23341 GND.n7217 GND.n7216 9.3005
R23342 GND.n7215 GND.n3417 9.3005
R23343 GND.n7214 GND.n7213 9.3005
R23344 GND.n7212 GND.n3421 9.3005
R23345 GND.n7211 GND.n7210 9.3005
R23346 GND.n7209 GND.n3425 9.3005
R23347 GND.n7208 GND.n7207 9.3005
R23348 GND.n7206 GND.n3429 9.3005
R23349 GND.n7205 GND.n7204 9.3005
R23350 GND.n7203 GND.n3433 9.3005
R23351 GND.n7202 GND.n7201 9.3005
R23352 GND.n7200 GND.n3437 9.3005
R23353 GND.n7199 GND.n7198 9.3005
R23354 GND.n7197 GND.n3441 9.3005
R23355 GND.n7196 GND.n7195 9.3005
R23356 GND.n7194 GND.n3445 9.3005
R23357 GND.n7193 GND.n7192 9.3005
R23358 GND.n7191 GND.n3449 9.3005
R23359 GND.n7190 GND.n7189 9.3005
R23360 GND.n7188 GND.n3453 9.3005
R23361 GND.n7187 GND.n7186 9.3005
R23362 GND.n7185 GND.n3457 9.3005
R23363 GND.n7184 GND.n7183 9.3005
R23364 GND.n7182 GND.n3461 9.3005
R23365 GND.n7181 GND.n7180 9.3005
R23366 GND.n7179 GND.n3465 9.3005
R23367 GND.n7178 GND.n7177 9.3005
R23368 GND.n7176 GND.n3469 9.3005
R23369 GND.n7175 GND.n7174 9.3005
R23370 GND.n7173 GND.n3473 9.3005
R23371 GND.n7172 GND.n7171 9.3005
R23372 GND.n7170 GND.n3477 9.3005
R23373 GND.n7169 GND.n7168 9.3005
R23374 GND.n7167 GND.n3481 9.3005
R23375 GND.n7166 GND.n7165 9.3005
R23376 GND.n7164 GND.n3485 9.3005
R23377 GND.n7163 GND.n7162 9.3005
R23378 GND.n7161 GND.n3489 9.3005
R23379 GND.n7160 GND.n7159 9.3005
R23380 GND.n7158 GND.n3493 9.3005
R23381 GND.n7157 GND.n7156 9.3005
R23382 GND.n7155 GND.n3497 9.3005
R23383 GND.n7154 GND.n7153 9.3005
R23384 GND.n7152 GND.n3501 9.3005
R23385 GND.n7151 GND.n7150 9.3005
R23386 GND.n7149 GND.n3505 9.3005
R23387 GND.n7148 GND.n7147 9.3005
R23388 GND.n7146 GND.n3509 9.3005
R23389 GND.n7145 GND.n7144 9.3005
R23390 GND.n7143 GND.n3513 9.3005
R23391 GND.n7142 GND.n7141 9.3005
R23392 GND.n7140 GND.n3517 9.3005
R23393 GND.n7139 GND.n7138 9.3005
R23394 GND.n7137 GND.n3521 9.3005
R23395 GND.n7136 GND.n7135 9.3005
R23396 GND.n7134 GND.n3525 9.3005
R23397 GND.n7133 GND.n7132 9.3005
R23398 GND.n7131 GND.n3529 9.3005
R23399 GND.n7130 GND.n7129 9.3005
R23400 GND.n7128 GND.n3533 9.3005
R23401 GND.n7127 GND.n7126 9.3005
R23402 GND.n7125 GND.n3537 9.3005
R23403 GND.n7124 GND.n7123 9.3005
R23404 GND.n7122 GND.n3541 9.3005
R23405 GND.n7121 GND.n7120 9.3005
R23406 GND.n7119 GND.n3545 9.3005
R23407 GND.n7118 GND.n7117 9.3005
R23408 GND.n7116 GND.n3549 9.3005
R23409 GND.n7115 GND.n7114 9.3005
R23410 GND.n7113 GND.n3553 9.3005
R23411 GND.n7112 GND.n7111 9.3005
R23412 GND.n7110 GND.n3557 9.3005
R23413 GND.n7109 GND.n7108 9.3005
R23414 GND.n7107 GND.n3561 9.3005
R23415 GND.n7106 GND.n7105 9.3005
R23416 GND.n7104 GND.n3565 9.3005
R23417 GND.n7103 GND.n577 9.3005
R23418 GND.n9501 GND.n576 9.3005
R23419 GND.n9503 GND.n9502 9.3005
R23420 GND.n555 GND.n554 9.3005
R23421 GND.n9519 GND.n9518 9.3005
R23422 GND.n9520 GND.n549 9.3005
R23423 GND.n9526 GND.n547 9.3005
R23424 GND.n9528 GND.n9527 9.3005
R23425 GND.n6326 GND.n6325 9.3005
R23426 GND.n7288 GND.n7287 9.3005
R23427 GND.n7286 GND.n7285 9.3005
R23428 GND.n3323 GND.n3322 9.3005
R23429 GND.n7280 GND.n7279 9.3005
R23430 GND.n7278 GND.n7277 9.3005
R23431 GND.n3333 GND.n3332 9.3005
R23432 GND.n7272 GND.n7271 9.3005
R23433 GND.n7270 GND.n7269 9.3005
R23434 GND.n3341 GND.n3340 9.3005
R23435 GND.n7264 GND.n7263 9.3005
R23436 GND.n7262 GND.n7261 9.3005
R23437 GND.n3353 GND.n3352 9.3005
R23438 GND.n3319 GND.n3317 9.3005
R23439 GND.n7266 GND.n7265 9.3005
R23440 GND.n7268 GND.n7267 9.3005
R23441 GND.n3337 GND.n3336 9.3005
R23442 GND.n7274 GND.n7273 9.3005
R23443 GND.n7276 GND.n7275 9.3005
R23444 GND.n3329 GND.n3328 9.3005
R23445 GND.n7282 GND.n7281 9.3005
R23446 GND.n7284 GND.n7283 9.3005
R23447 GND.n3318 GND.n3316 9.3005
R23448 GND.n7290 GND.n7289 9.3005
R23449 GND.n7291 GND.n3315 9.3005
R23450 GND.n3349 GND.n3348 9.3005
R23451 GND.n7260 GND.n7259 9.3005
R23452 GND.n6428 GND.n6427 9.3005
R23453 GND.n6426 GND.n3963 9.3005
R23454 GND.n6425 GND.n6424 9.3005
R23455 GND.n6423 GND.n6422 9.3005
R23456 GND.n6421 GND.n3970 9.3005
R23457 GND.n6420 GND.n6419 9.3005
R23458 GND.n6418 GND.n3227 9.3005
R23459 GND.n3055 GND.n3054 9.3005
R23460 GND.n3056 GND.n3026 9.3005
R23461 GND.n7551 GND.n7550 9.3005
R23462 GND.n7549 GND.n3027 9.3005
R23463 GND.n7548 GND.n7547 9.3005
R23464 GND.n7546 GND.n3057 9.3005
R23465 GND.n7545 GND.n7544 9.3005
R23466 GND.n7543 GND.n3061 9.3005
R23467 GND.n7542 GND.n7541 9.3005
R23468 GND.n7540 GND.n3062 9.3005
R23469 GND.n7539 GND.n7538 9.3005
R23470 GND.n7537 GND.n3066 9.3005
R23471 GND.n7536 GND.n7535 9.3005
R23472 GND.n7534 GND.n3067 9.3005
R23473 GND.n7533 GND.n7532 9.3005
R23474 GND.n7531 GND.n3071 9.3005
R23475 GND.n7530 GND.n7529 9.3005
R23476 GND.n7528 GND.n3072 9.3005
R23477 GND.n7527 GND.n7526 9.3005
R23478 GND.n7525 GND.n3076 9.3005
R23479 GND.n7524 GND.n7523 9.3005
R23480 GND.n7522 GND.n3077 9.3005
R23481 GND.n7521 GND.n7520 9.3005
R23482 GND.n7519 GND.n3081 9.3005
R23483 GND.n7518 GND.n7517 9.3005
R23484 GND.n7516 GND.n3082 9.3005
R23485 GND.n7515 GND.n7514 9.3005
R23486 GND.n7513 GND.n3086 9.3005
R23487 GND.n7512 GND.n7511 9.3005
R23488 GND.n7510 GND.n3087 9.3005
R23489 GND.n7509 GND.n7508 9.3005
R23490 GND.n7507 GND.n3091 9.3005
R23491 GND.n7506 GND.n7505 9.3005
R23492 GND.n7504 GND.n3092 9.3005
R23493 GND.n7503 GND.n7502 9.3005
R23494 GND.n7501 GND.n3096 9.3005
R23495 GND.n7500 GND.n7499 9.3005
R23496 GND.n7498 GND.n3097 9.3005
R23497 GND.n7497 GND.n7496 9.3005
R23498 GND.n7495 GND.n3101 9.3005
R23499 GND.n7494 GND.n7493 9.3005
R23500 GND.n7492 GND.n3102 9.3005
R23501 GND.n7491 GND.n7490 9.3005
R23502 GND.n7489 GND.n3106 9.3005
R23503 GND.n7488 GND.n7487 9.3005
R23504 GND.n7486 GND.n3107 9.3005
R23505 GND.n7485 GND.n7484 9.3005
R23506 GND.n7483 GND.n3111 9.3005
R23507 GND.n7482 GND.n7481 9.3005
R23508 GND.n7480 GND.n3112 9.3005
R23509 GND.n7479 GND.n7478 9.3005
R23510 GND.n7477 GND.n3116 9.3005
R23511 GND.n7476 GND.n7475 9.3005
R23512 GND.n7474 GND.n3117 9.3005
R23513 GND.n7473 GND.n7472 9.3005
R23514 GND.n7471 GND.n3121 9.3005
R23515 GND.n7470 GND.n7469 9.3005
R23516 GND.n7468 GND.n3122 9.3005
R23517 GND.n7467 GND.n7466 9.3005
R23518 GND.n7465 GND.n3126 9.3005
R23519 GND.n7464 GND.n7463 9.3005
R23520 GND.n7462 GND.n3127 9.3005
R23521 GND.n7461 GND.n7460 9.3005
R23522 GND.n7459 GND.n3131 9.3005
R23523 GND.n7458 GND.n7457 9.3005
R23524 GND.n7456 GND.n3132 9.3005
R23525 GND.n7455 GND.n7454 9.3005
R23526 GND.n7453 GND.n3136 9.3005
R23527 GND.n7452 GND.n7451 9.3005
R23528 GND.n7450 GND.n3137 9.3005
R23529 GND.n7449 GND.n7448 9.3005
R23530 GND.n7447 GND.n3141 9.3005
R23531 GND.n7446 GND.n7445 9.3005
R23532 GND.n7444 GND.n3142 9.3005
R23533 GND.n7443 GND.n7442 9.3005
R23534 GND.n7441 GND.n3146 9.3005
R23535 GND.n7440 GND.n7439 9.3005
R23536 GND.n7438 GND.n3147 9.3005
R23537 GND.n7437 GND.n7436 9.3005
R23538 GND.n7435 GND.n3151 9.3005
R23539 GND.n7434 GND.n7433 9.3005
R23540 GND.n7432 GND.n3152 9.3005
R23541 GND.n7431 GND.n7430 9.3005
R23542 GND.n7429 GND.n3156 9.3005
R23543 GND.n7428 GND.n7427 9.3005
R23544 GND.n7426 GND.n3157 9.3005
R23545 GND.n7425 GND.n7424 9.3005
R23546 GND.n7423 GND.n3161 9.3005
R23547 GND.n7422 GND.n7421 9.3005
R23548 GND.n7420 GND.n3162 9.3005
R23549 GND.n7419 GND.n7418 9.3005
R23550 GND.n7417 GND.n3166 9.3005
R23551 GND.n7416 GND.n7415 9.3005
R23552 GND.n7414 GND.n3167 9.3005
R23553 GND.n7413 GND.n7412 9.3005
R23554 GND.n7411 GND.n3171 9.3005
R23555 GND.n7410 GND.n7409 9.3005
R23556 GND.n7408 GND.n3172 9.3005
R23557 GND.n7407 GND.n7406 9.3005
R23558 GND.n7405 GND.n3176 9.3005
R23559 GND.n7404 GND.n7403 9.3005
R23560 GND.n7402 GND.n3177 9.3005
R23561 GND.n7401 GND.n7400 9.3005
R23562 GND.n7399 GND.n3181 9.3005
R23563 GND.n7398 GND.n7397 9.3005
R23564 GND.n7396 GND.n3182 9.3005
R23565 GND.n7395 GND.n7394 9.3005
R23566 GND.n7393 GND.n3186 9.3005
R23567 GND.n7392 GND.n7391 9.3005
R23568 GND.n7390 GND.n3187 9.3005
R23569 GND.n7389 GND.n7388 9.3005
R23570 GND.n7387 GND.n3191 9.3005
R23571 GND.n7386 GND.n7385 9.3005
R23572 GND.n7384 GND.n3192 9.3005
R23573 GND.n7383 GND.n7382 9.3005
R23574 GND.n7381 GND.n3196 9.3005
R23575 GND.n7380 GND.n7379 9.3005
R23576 GND.n7378 GND.n3197 9.3005
R23577 GND.n7377 GND.n7376 9.3005
R23578 GND.n7375 GND.n3201 9.3005
R23579 GND.n7374 GND.n7373 9.3005
R23580 GND.n7372 GND.n3202 9.3005
R23581 GND.n7371 GND.n7370 9.3005
R23582 GND.n7369 GND.n3206 9.3005
R23583 GND.n7368 GND.n7367 9.3005
R23584 GND.n7366 GND.n3207 9.3005
R23585 GND.n7365 GND.n7364 9.3005
R23586 GND.n7363 GND.n3211 9.3005
R23587 GND.n7362 GND.n7361 9.3005
R23588 GND.n7360 GND.n3212 9.3005
R23589 GND.n7359 GND.n7358 9.3005
R23590 GND.n7357 GND.n3216 9.3005
R23591 GND.n7356 GND.n7355 9.3005
R23592 GND.n7354 GND.n3217 9.3005
R23593 GND.n7353 GND.n7352 9.3005
R23594 GND.n7351 GND.n3221 9.3005
R23595 GND.n7350 GND.n7349 9.3005
R23596 GND.n7348 GND.n3222 9.3005
R23597 GND.n7347 GND.n7346 9.3005
R23598 GND.n7345 GND.n3226 9.3005
R23599 GND.n7344 GND.n7343 9.3005
R23600 GND.n3053 GND.n3051 9.3005
R23601 GND.n3048 GND.n3028 9.3005
R23602 GND.n3046 GND.n3045 9.3005
R23603 GND.n3044 GND.n3029 9.3005
R23604 GND.n3043 GND.n3042 9.3005
R23605 GND.n3036 GND.n3032 9.3005
R23606 GND.n3035 GND.n1887 9.3005
R23607 GND.n3050 GND.n3049 9.3005
R23608 GND.n2776 GND.n2188 9.3005
R23609 GND.n2778 GND.n2777 9.3005
R23610 GND.n2779 GND.n2187 9.3005
R23611 GND.n2781 GND.n2780 9.3005
R23612 GND.n2096 GND.n2095 9.3005
R23613 GND.n2833 GND.n2832 9.3005
R23614 GND.n2834 GND.n2093 9.3005
R23615 GND.n2837 GND.n2836 9.3005
R23616 GND.n2835 GND.n2094 9.3005
R23617 GND.n2073 GND.n2072 9.3005
R23618 GND.n2858 GND.n2857 9.3005
R23619 GND.n2859 GND.n2070 9.3005
R23620 GND.n2862 GND.n2861 9.3005
R23621 GND.n2860 GND.n2071 9.3005
R23622 GND.n2051 GND.n2050 9.3005
R23623 GND.n2883 GND.n2882 9.3005
R23624 GND.n2884 GND.n2048 9.3005
R23625 GND.n2887 GND.n2886 9.3005
R23626 GND.n2885 GND.n2049 9.3005
R23627 GND.n2024 GND.n2023 9.3005
R23628 GND.n7681 GND.n7680 9.3005
R23629 GND.n7682 GND.n2021 9.3005
R23630 GND.n7685 GND.n7684 9.3005
R23631 GND.n7683 GND.n2022 9.3005
R23632 GND.n2000 GND.n1999 9.3005
R23633 GND.n7705 GND.n7704 9.3005
R23634 GND.n7706 GND.n1997 9.3005
R23635 GND.n7709 GND.n7708 9.3005
R23636 GND.n7707 GND.n1998 9.3005
R23637 GND.n1977 GND.n1976 9.3005
R23638 GND.n7730 GND.n7729 9.3005
R23639 GND.n7731 GND.n1974 9.3005
R23640 GND.n7734 GND.n7733 9.3005
R23641 GND.n7732 GND.n1975 9.3005
R23642 GND.n1955 GND.n1954 9.3005
R23643 GND.n7755 GND.n7754 9.3005
R23644 GND.n7756 GND.n1952 9.3005
R23645 GND.n7759 GND.n7758 9.3005
R23646 GND.n7757 GND.n1953 9.3005
R23647 GND.n1933 GND.n1932 9.3005
R23648 GND.n7780 GND.n7779 9.3005
R23649 GND.n7781 GND.n1930 9.3005
R23650 GND.n7784 GND.n7783 9.3005
R23651 GND.n7782 GND.n1931 9.3005
R23652 GND.n1910 GND.n1909 9.3005
R23653 GND.n7804 GND.n7803 9.3005
R23654 GND.n7805 GND.n1907 9.3005
R23655 GND.n7813 GND.n7812 9.3005
R23656 GND.n7811 GND.n1908 9.3005
R23657 GND.n7810 GND.n7809 9.3005
R23658 GND.n7806 GND.n1889 9.3005
R23659 GND.n7831 GND.n1888 9.3005
R23660 GND.n7833 GND.n7832 9.3005
R23661 GND.n7835 GND.n1886 9.3005
R23662 GND.n7840 GND.n7839 9.3005
R23663 GND.n7842 GND.n7841 9.3005
R23664 GND.n1875 GND.n1874 9.3005
R23665 GND.n7848 GND.n7847 9.3005
R23666 GND.n7850 GND.n7849 9.3005
R23667 GND.n1865 GND.n1864 9.3005
R23668 GND.n7856 GND.n7855 9.3005
R23669 GND.n7858 GND.n7857 9.3005
R23670 GND.n1854 GND.n1851 9.3005
R23671 GND.n7864 GND.n7863 9.3005
R23672 GND.n1852 GND.n1836 9.3005
R23673 GND.n7870 GND.n7869 9.3005
R23674 GND.n1835 GND.n1833 9.3005
R23675 GND.n1855 GND.n1853 9.3005
R23676 GND.n7862 GND.n7861 9.3005
R23677 GND.n7860 GND.n7859 9.3005
R23678 GND.n1861 GND.n1860 9.3005
R23679 GND.n7854 GND.n7853 9.3005
R23680 GND.n7852 GND.n7851 9.3005
R23681 GND.n1869 GND.n1868 9.3005
R23682 GND.n7846 GND.n7845 9.3005
R23683 GND.n7844 GND.n7843 9.3005
R23684 GND.n1883 GND.n1882 9.3005
R23685 GND.n7838 GND.n7837 9.3005
R23686 GND.n7872 GND.n7871 9.3005
R23687 GND.n7906 GND.n1788 9.3005
R23688 GND.n7908 GND.n7907 9.3005
R23689 GND.n7909 GND.n1787 9.3005
R23690 GND.n7911 GND.n7910 9.3005
R23691 GND.n7912 GND.n1783 9.3005
R23692 GND.n7914 GND.n7913 9.3005
R23693 GND.n7915 GND.n1782 9.3005
R23694 GND.n7917 GND.n7916 9.3005
R23695 GND.n7918 GND.n1779 9.3005
R23696 GND.n7920 GND.n7919 9.3005
R23697 GND.n7904 GND.n7903 9.3005
R23698 GND.n7902 GND.n1797 9.3005
R23699 GND.n7901 GND.n7900 9.3005
R23700 GND.n7899 GND.n1798 9.3005
R23701 GND.n7898 GND.n7897 9.3005
R23702 GND.n7896 GND.n1802 9.3005
R23703 GND.n7895 GND.n7894 9.3005
R23704 GND.n7893 GND.n1803 9.3005
R23705 GND.n7892 GND.n7891 9.3005
R23706 GND.n7890 GND.n1807 9.3005
R23707 GND.n7889 GND.n7888 9.3005
R23708 GND.n7887 GND.n1808 9.3005
R23709 GND.n7886 GND.n1813 9.3005
R23710 GND.n7885 GND.n7884 9.3005
R23711 GND.n1563 GND.n1562 9.3005
R23712 GND.n1565 GND.n1557 9.3005
R23713 GND.n1567 GND.n1566 9.3005
R23714 GND.n1554 GND.n1552 9.3005
R23715 GND.n8078 GND.n8077 9.3005
R23716 GND.n1555 GND.n1553 9.3005
R23717 GND.n8073 GND.n1573 9.3005
R23718 GND.n8072 GND.n1574 9.3005
R23719 GND.n8071 GND.n1575 9.3005
R23720 GND.n2527 GND.n1576 9.3005
R23721 GND.n8067 GND.n1581 9.3005
R23722 GND.n8066 GND.n1582 9.3005
R23723 GND.n8065 GND.n1583 9.3005
R23724 GND.n2341 GND.n1584 9.3005
R23725 GND.n8061 GND.n1589 9.3005
R23726 GND.n8060 GND.n1590 9.3005
R23727 GND.n8059 GND.n1591 9.3005
R23728 GND.n2318 GND.n1592 9.3005
R23729 GND.n8055 GND.n1597 9.3005
R23730 GND.n8054 GND.n1598 9.3005
R23731 GND.n8053 GND.n1599 9.3005
R23732 GND.n2305 GND.n1600 9.3005
R23733 GND.n8049 GND.n1605 9.3005
R23734 GND.n8048 GND.n1606 9.3005
R23735 GND.n8047 GND.n1607 9.3005
R23736 GND.n2599 GND.n1608 9.3005
R23737 GND.n8043 GND.n1613 9.3005
R23738 GND.n8042 GND.n1614 9.3005
R23739 GND.n8041 GND.n1615 9.3005
R23740 GND.n2634 GND.n1616 9.3005
R23741 GND.n8037 GND.n1621 9.3005
R23742 GND.n8036 GND.n1622 9.3005
R23743 GND.n8035 GND.n1623 9.3005
R23744 GND.n2701 GND.n1624 9.3005
R23745 GND.n8031 GND.n1629 9.3005
R23746 GND.n8030 GND.n1630 9.3005
R23747 GND.n8029 GND.n1631 9.3005
R23748 GND.n2231 GND.n1632 9.3005
R23749 GND.n8025 GND.n1637 9.3005
R23750 GND.n8024 GND.n1638 9.3005
R23751 GND.n8023 GND.n1639 9.3005
R23752 GND.n2208 GND.n1640 9.3005
R23753 GND.n8019 GND.n1645 9.3005
R23754 GND.n8018 GND.n1646 9.3005
R23755 GND.n8017 GND.n1647 9.3005
R23756 GND.n2197 GND.n1648 9.3005
R23757 GND.n8013 GND.n1653 9.3005
R23758 GND.n8012 GND.n1654 9.3005
R23759 GND.n8011 GND.n1655 9.3005
R23760 GND.n2121 GND.n1656 9.3005
R23761 GND.n8007 GND.n1661 9.3005
R23762 GND.n8006 GND.n1662 9.3005
R23763 GND.n8005 GND.n1663 9.3005
R23764 GND.n2144 GND.n1664 9.3005
R23765 GND.n8001 GND.n1669 9.3005
R23766 GND.n8000 GND.n1670 9.3005
R23767 GND.n7999 GND.n1671 9.3005
R23768 GND.n2100 GND.n1672 9.3005
R23769 GND.n7995 GND.n1677 9.3005
R23770 GND.n7994 GND.n1678 9.3005
R23771 GND.n7993 GND.n1679 9.3005
R23772 GND.n2841 GND.n1680 9.3005
R23773 GND.n7989 GND.n1685 9.3005
R23774 GND.n7988 GND.n1686 9.3005
R23775 GND.n7987 GND.n1687 9.3005
R23776 GND.n2868 GND.n1688 9.3005
R23777 GND.n7983 GND.n1693 9.3005
R23778 GND.n7982 GND.n1694 9.3005
R23779 GND.n7981 GND.n1695 9.3005
R23780 GND.n2038 GND.n1696 9.3005
R23781 GND.n7977 GND.n1701 9.3005
R23782 GND.n7976 GND.n1702 9.3005
R23783 GND.n7975 GND.n1703 9.3005
R23784 GND.n2017 GND.n1704 9.3005
R23785 GND.n7971 GND.n1709 9.3005
R23786 GND.n7970 GND.n1710 9.3005
R23787 GND.n7969 GND.n1711 9.3005
R23788 GND.n2004 GND.n1712 9.3005
R23789 GND.n7965 GND.n1717 9.3005
R23790 GND.n7964 GND.n1718 9.3005
R23791 GND.n7963 GND.n1719 9.3005
R23792 GND.n7713 GND.n1720 9.3005
R23793 GND.n7959 GND.n1725 9.3005
R23794 GND.n7958 GND.n1726 9.3005
R23795 GND.n7957 GND.n1727 9.3005
R23796 GND.n7740 GND.n1728 9.3005
R23797 GND.n7953 GND.n1733 9.3005
R23798 GND.n7952 GND.n1734 9.3005
R23799 GND.n7951 GND.n1735 9.3005
R23800 GND.n1949 GND.n1736 9.3005
R23801 GND.n7947 GND.n1741 9.3005
R23802 GND.n7946 GND.n1742 9.3005
R23803 GND.n7945 GND.n1743 9.3005
R23804 GND.n1926 GND.n1744 9.3005
R23805 GND.n7941 GND.n1749 9.3005
R23806 GND.n7940 GND.n1750 9.3005
R23807 GND.n7939 GND.n1751 9.3005
R23808 GND.n1913 GND.n1752 9.3005
R23809 GND.n7935 GND.n1757 9.3005
R23810 GND.n7934 GND.n1758 9.3005
R23811 GND.n7933 GND.n1759 9.3005
R23812 GND.n1892 GND.n1760 9.3005
R23813 GND.n7929 GND.n1765 9.3005
R23814 GND.n7928 GND.n1766 9.3005
R23815 GND.n7927 GND.n1767 9.3005
R23816 GND.n1508 GND.n1504 9.3005
R23817 GND.n1562 GND.n1561 9.3005
R23818 GND.n1557 GND.n1556 9.3005
R23819 GND.n1568 GND.n1567 9.3005
R23820 GND.n1569 GND.n1554 9.3005
R23821 GND.n8077 GND.n8076 9.3005
R23822 GND.n8075 GND.n1555 9.3005
R23823 GND.n8074 GND.n8073 9.3005
R23824 GND.n8072 GND.n1572 9.3005
R23825 GND.n8071 GND.n8070 9.3005
R23826 GND.n8069 GND.n1576 9.3005
R23827 GND.n8068 GND.n8067 9.3005
R23828 GND.n8066 GND.n1580 9.3005
R23829 GND.n8065 GND.n8064 9.3005
R23830 GND.n8063 GND.n1584 9.3005
R23831 GND.n8062 GND.n8061 9.3005
R23832 GND.n8060 GND.n1588 9.3005
R23833 GND.n8059 GND.n8058 9.3005
R23834 GND.n8057 GND.n1592 9.3005
R23835 GND.n8056 GND.n8055 9.3005
R23836 GND.n8054 GND.n1596 9.3005
R23837 GND.n8053 GND.n8052 9.3005
R23838 GND.n8051 GND.n1600 9.3005
R23839 GND.n8050 GND.n8049 9.3005
R23840 GND.n8048 GND.n1604 9.3005
R23841 GND.n8047 GND.n8046 9.3005
R23842 GND.n8045 GND.n1608 9.3005
R23843 GND.n8044 GND.n8043 9.3005
R23844 GND.n8042 GND.n1612 9.3005
R23845 GND.n8041 GND.n8040 9.3005
R23846 GND.n8039 GND.n1616 9.3005
R23847 GND.n8038 GND.n8037 9.3005
R23848 GND.n8036 GND.n1620 9.3005
R23849 GND.n8035 GND.n8034 9.3005
R23850 GND.n8033 GND.n1624 9.3005
R23851 GND.n8032 GND.n8031 9.3005
R23852 GND.n8030 GND.n1628 9.3005
R23853 GND.n8029 GND.n8028 9.3005
R23854 GND.n8027 GND.n1632 9.3005
R23855 GND.n8026 GND.n8025 9.3005
R23856 GND.n8024 GND.n1636 9.3005
R23857 GND.n8023 GND.n8022 9.3005
R23858 GND.n8021 GND.n1640 9.3005
R23859 GND.n8020 GND.n8019 9.3005
R23860 GND.n8018 GND.n1644 9.3005
R23861 GND.n8017 GND.n8016 9.3005
R23862 GND.n8015 GND.n1648 9.3005
R23863 GND.n8014 GND.n8013 9.3005
R23864 GND.n8012 GND.n1652 9.3005
R23865 GND.n8011 GND.n8010 9.3005
R23866 GND.n8009 GND.n1656 9.3005
R23867 GND.n8008 GND.n8007 9.3005
R23868 GND.n8006 GND.n1660 9.3005
R23869 GND.n8005 GND.n8004 9.3005
R23870 GND.n8003 GND.n1664 9.3005
R23871 GND.n8002 GND.n8001 9.3005
R23872 GND.n8000 GND.n1668 9.3005
R23873 GND.n7999 GND.n7998 9.3005
R23874 GND.n7997 GND.n1672 9.3005
R23875 GND.n7996 GND.n7995 9.3005
R23876 GND.n7994 GND.n1676 9.3005
R23877 GND.n7993 GND.n7992 9.3005
R23878 GND.n7991 GND.n1680 9.3005
R23879 GND.n7990 GND.n7989 9.3005
R23880 GND.n7988 GND.n1684 9.3005
R23881 GND.n7987 GND.n7986 9.3005
R23882 GND.n7985 GND.n1688 9.3005
R23883 GND.n7984 GND.n7983 9.3005
R23884 GND.n7982 GND.n1692 9.3005
R23885 GND.n7981 GND.n7980 9.3005
R23886 GND.n7979 GND.n1696 9.3005
R23887 GND.n7978 GND.n7977 9.3005
R23888 GND.n7976 GND.n1700 9.3005
R23889 GND.n7975 GND.n7974 9.3005
R23890 GND.n7973 GND.n1704 9.3005
R23891 GND.n7972 GND.n7971 9.3005
R23892 GND.n7970 GND.n1708 9.3005
R23893 GND.n7969 GND.n7968 9.3005
R23894 GND.n7967 GND.n1712 9.3005
R23895 GND.n7966 GND.n7965 9.3005
R23896 GND.n7964 GND.n1716 9.3005
R23897 GND.n7963 GND.n7962 9.3005
R23898 GND.n7961 GND.n1720 9.3005
R23899 GND.n7960 GND.n7959 9.3005
R23900 GND.n7958 GND.n1724 9.3005
R23901 GND.n7957 GND.n7956 9.3005
R23902 GND.n7955 GND.n1728 9.3005
R23903 GND.n7954 GND.n7953 9.3005
R23904 GND.n7952 GND.n1732 9.3005
R23905 GND.n7951 GND.n7950 9.3005
R23906 GND.n7949 GND.n1736 9.3005
R23907 GND.n7948 GND.n7947 9.3005
R23908 GND.n7946 GND.n1740 9.3005
R23909 GND.n7945 GND.n7944 9.3005
R23910 GND.n7943 GND.n1744 9.3005
R23911 GND.n7942 GND.n7941 9.3005
R23912 GND.n7940 GND.n1748 9.3005
R23913 GND.n7939 GND.n7938 9.3005
R23914 GND.n7937 GND.n1752 9.3005
R23915 GND.n7936 GND.n7935 9.3005
R23916 GND.n7934 GND.n1756 9.3005
R23917 GND.n7933 GND.n7932 9.3005
R23918 GND.n7931 GND.n1760 9.3005
R23919 GND.n7930 GND.n7929 9.3005
R23920 GND.n7928 GND.n1764 9.3005
R23921 GND.n7927 GND.n7926 9.3005
R23922 GND.n1558 GND.n1504 9.3005
R23923 GND.n2406 GND.n2405 9.3005
R23924 GND.n2404 GND.n2379 9.3005
R23925 GND.n2403 GND.n2402 9.3005
R23926 GND.n2399 GND.n2382 9.3005
R23927 GND.n2398 GND.n2397 9.3005
R23928 GND.n2396 GND.n2383 9.3005
R23929 GND.n2395 GND.n2394 9.3005
R23930 GND.n2391 GND.n2386 9.3005
R23931 GND.n2390 GND.n2389 9.3005
R23932 GND.n1506 GND.n1505 9.3005
R23933 GND.n8098 GND.n8097 9.3005
R23934 GND.n2407 GND.n2375 9.3005
R23935 GND.n2409 GND.n2408 9.3005
R23936 GND.n2412 GND.n2411 9.3005
R23937 GND.n2415 GND.n2373 9.3005
R23938 GND.n2417 GND.n2416 9.3005
R23939 GND.n2418 GND.n2372 9.3005
R23940 GND.n2420 GND.n2419 9.3005
R23941 GND.n2421 GND.n2368 9.3005
R23942 GND.n2517 GND.n2516 9.3005
R23943 GND.n2518 GND.n2366 9.3005
R23944 GND.n2521 GND.n2520 9.3005
R23945 GND.n2519 GND.n2367 9.3005
R23946 GND.n2347 GND.n2346 9.3005
R23947 GND.n2542 GND.n2541 9.3005
R23948 GND.n2543 GND.n2344 9.3005
R23949 GND.n2546 GND.n2545 9.3005
R23950 GND.n2544 GND.n2345 9.3005
R23951 GND.n2325 GND.n2324 9.3005
R23952 GND.n2567 GND.n2566 9.3005
R23953 GND.n2568 GND.n2322 9.3005
R23954 GND.n2571 GND.n2570 9.3005
R23955 GND.n2569 GND.n2323 9.3005
R23956 GND.n2301 GND.n2300 9.3005
R23957 GND.n2591 GND.n2590 9.3005
R23958 GND.n2592 GND.n2298 9.3005
R23959 GND.n2595 GND.n2594 9.3005
R23960 GND.n2593 GND.n2299 9.3005
R23961 GND.n2278 GND.n2277 9.3005
R23962 GND.n2616 GND.n2615 9.3005
R23963 GND.n2617 GND.n2275 9.3005
R23964 GND.n2629 GND.n2628 9.3005
R23965 GND.n2627 GND.n2276 9.3005
R23966 GND.n2626 GND.n2625 9.3005
R23967 GND.n2624 GND.n2618 9.3005
R23968 GND.n2623 GND.n2622 9.3005
R23969 GND.n2621 GND.n2620 9.3005
R23970 GND.n2237 GND.n2236 9.3005
R23971 GND.n2716 GND.n2715 9.3005
R23972 GND.n2717 GND.n2234 9.3005
R23973 GND.n2720 GND.n2719 9.3005
R23974 GND.n2718 GND.n2235 9.3005
R23975 GND.n2215 GND.n2214 9.3005
R23976 GND.n2741 GND.n2740 9.3005
R23977 GND.n2742 GND.n2212 9.3005
R23978 GND.n2745 GND.n2744 9.3005
R23979 GND.n2743 GND.n2213 9.3005
R23980 GND.n2193 GND.n2192 9.3005
R23981 GND.n2763 GND.n2762 9.3005
R23982 GND.n2764 GND.n2191 9.3005
R23983 GND.n2766 GND.n2765 9.3005
R23984 GND.n2767 GND.n2190 9.3005
R23985 GND.n2771 GND.n2770 9.3005
R23986 GND.n2772 GND.n2189 9.3005
R23987 GND.n2775 GND.n2774 9.3005
R23988 GND.n2410 GND.n2374 9.3005
R23989 GND.n200 GND.n199 9.3005
R23990 GND.n193 GND.n192 9.3005
R23991 GND.n188 GND.n187 9.3005
R23992 GND.n181 GND.n180 9.3005
R23993 GND.n176 GND.n175 9.3005
R23994 GND.n169 GND.n168 9.3005
R23995 GND.n164 GND.n163 9.3005
R23996 GND.n157 GND.n156 9.3005
R23997 GND.n152 GND.n151 9.3005
R23998 GND.n145 GND.n144 9.3005
R23999 GND.n141 GND.n140 9.3005
R24000 GND.n134 GND.n133 9.3005
R24001 GND.n271 GND.n270 9.3005
R24002 GND.n264 GND.n263 9.3005
R24003 GND.n259 GND.n258 9.3005
R24004 GND.n252 GND.n251 9.3005
R24005 GND.n247 GND.n246 9.3005
R24006 GND.n240 GND.n239 9.3005
R24007 GND.n235 GND.n234 9.3005
R24008 GND.n228 GND.n227 9.3005
R24009 GND.n223 GND.n222 9.3005
R24010 GND.n216 GND.n215 9.3005
R24011 GND.n212 GND.n211 9.3005
R24012 GND.n205 GND.n204 9.3005
R24013 GND.n2760 GND.t39 9.1943
R24014 GND.n2103 GND.t65 9.1943
R24015 GND.n4906 GND.n4646 9.1943
R24016 GND.n4990 GND.n4598 9.1943
R24017 GND.n5069 GND.n4559 9.1943
R24018 GND.n5153 GND.n4510 9.1943
R24019 GND.n5229 GND.n4474 9.1943
R24020 GND.n5314 GND.n4427 9.1943
R24021 GND.n5391 GND.n4388 9.1943
R24022 GND.n5474 GND.n4340 9.1943
R24023 GND.n5562 GND.n4302 9.1943
R24024 GND.n5630 GND.n4256 9.1943
R24025 GND.n5676 GND.n4218 9.1943
R24026 GND.n5827 GND.n4172 9.1943
R24027 GND.n5877 GND.n4133 9.1943
R24028 GND.n5960 GND.n4085 9.1943
R24029 GND.n6028 GND.n4045 9.1943
R24030 GND.n6342 GND.n6341 9.1943
R24031 GND.n7315 GND.t154 9.1943
R24032 GND.n3782 GND.t46 9.1943
R24033 GND.n6888 GND.t34 9.1943
R24034 GND.n6328 GND.n6327 8.99709
R24035 GND.n1834 GND.n1768 8.99709
R24036 GND.n7601 GND.n2955 8.81123
R24037 GND.n6213 GND.n6195 8.72777
R24038 GND.n7906 GND.n7905 8.72777
R24039 GND.n6292 GND.n6119 8.72777
R24040 GND.n2696 GND.t32 8.42815
R24041 GND.n7663 GND.t36 8.42815
R24042 GND.t108 GND.n2963 8.42815
R24043 GND.t98 GND.n2973 8.42815
R24044 GND.n5294 GND.t8 8.42815
R24045 GND.n5696 GND.t3 8.42815
R24046 GND.t41 GND.n3836 8.42815
R24047 GND.n6959 GND.t55 8.42815
R24048 GND.n9695 GND.n9694 8.30425
R24049 GND.n2773 GND.n131 8.30425
R24050 GND.n2575 GND.t53 7.662
R24051 GND.n1984 GND.t44 7.662
R24052 GND.n7581 GND.t118 7.662
R24053 GND.n7560 GND.n7559 7.662
R24054 GND.n4856 GND.n4855 7.662
R24055 GND.n4953 GND.t9 7.662
R24056 GND.n5000 GND.n4589 7.662
R24057 GND.n5050 GND.n5049 7.662
R24058 GND.n5163 GND.n4503 7.662
R24059 GND.n5213 GND.n5212 7.662
R24060 GND.n5324 GND.n4417 7.662
R24061 GND.n5375 GND.n5374 7.662
R24062 GND.n5351 GND.t23 7.662
R24063 GND.n5484 GND.n4331 7.662
R24064 GND.n5546 GND.n5544 7.662
R24065 GND.n5495 GND.t31 7.662
R24066 GND.n5639 GND.n5638 7.662
R24067 GND.n5650 GND.n4235 7.662
R24068 GND.n5834 GND.n4160 7.662
R24069 GND.n5861 GND.n5860 7.662
R24070 GND.n5970 GND.n4075 7.662
R24071 GND.n6009 GND.n6008 7.662
R24072 GND.n6042 GND.t26 7.662
R24073 GND.n6055 GND.n3989 7.662
R24074 GND.n6393 GND.n3978 7.662
R24075 GND.n3895 GND.t63 7.662
R24076 GND.n7024 GND.t49 7.662
R24077 GND.n4717 GND.n4716 7.30353
R24078 GND.n6212 GND.n6211 7.30353
R24079 GND.n4855 GND.t121 7.27893
R24080 GND.n6055 GND.t163 7.27893
R24081 GND.n6179 GND.n6137 6.5566
R24082 GND.n4772 GND.n4771 6.5566
R24083 GND.n4758 GND.n4757 6.5566
R24084 GND.n6221 GND.n6220 6.5566
R24085 GND.n131 GND.n130 6.37315
R24086 GND.n9695 GND.n405 6.37315
R24087 GND.n129 GND.n85 6.12981
R24088 GND.n361 GND.n317 6.12981
R24089 GND.t118 GND.n7580 6.1297
R24090 GND.t135 GND.n1849 6.1297
R24091 GND.n4848 GND.n4669 6.1297
R24092 GND.n7553 GND.n3021 6.1297
R24093 GND.n4592 GND.n4582 6.1297
R24094 GND.n5043 GND.n5042 6.1297
R24095 GND.n5144 GND.n4496 6.1297
R24096 GND.n5206 GND.n5205 6.1297
R24097 GND.n5212 GND.t16 6.1297
R24098 GND.n4421 GND.n4410 6.1297
R24099 GND.n5368 GND.n5367 6.1297
R24100 GND.n5432 GND.t23 6.1297
R24101 GND.n4334 GND.n4324 6.1297
R24102 GND.n5538 GND.n5537 6.1297
R24103 GND.n5584 GND.t31 6.1297
R24104 GND.n5645 GND.n4244 6.1297
R24105 GND.n5686 GND.n4232 6.1297
R24106 GND.t13 GND.n5834 6.1297
R24107 GND.n4162 GND.n4155 6.1297
R24108 GND.n5854 GND.n5853 6.1297
R24109 GND.n4079 GND.n4068 6.1297
R24110 GND.n6002 GND.n6001 6.1297
R24111 GND.n6361 GND.n3983 6.1297
R24112 GND.n6369 GND.n3985 6.1297
R24113 GND.n6400 GND.t125 6.1297
R24114 GND.n6422 GND.n3969 5.81868
R24115 GND.n3041 GND.n3029 5.81868
R24116 GND.n5259 GND.t11 5.74663
R24117 GND.t0 GND.n4194 5.74663
R24118 GND.n6257 GND.t88 5.74663
R24119 GND.n6260 GND.n6120 5.62001
R24120 GND.n4686 GND.n1795 5.62001
R24121 GND.n4687 GND.n1795 5.62001
R24122 GND.n6260 GND.n6121 5.62001
R24123 GND.n7574 GND.t81 5.36355
R24124 GND.t81 GND.n7573 5.36355
R24125 GND.n6140 GND.t170 5.36355
R24126 GND.n62 GND.t67 5.26646
R24127 GND.n62 GND.t37 5.26646
R24128 GND.n64 GND.t38 5.26646
R24129 GND.n64 GND.t68 5.26646
R24130 GND.n105 GND.t79 5.26646
R24131 GND.n105 GND.t48 5.26646
R24132 GND.n107 GND.t33 5.26646
R24133 GND.n107 GND.t40 5.26646
R24134 GND.n19 GND.t66 5.26646
R24135 GND.n19 GND.t71 5.26646
R24136 GND.n21 GND.t52 5.26646
R24137 GND.n21 GND.t72 5.26646
R24138 GND.n296 GND.t35 5.26646
R24139 GND.n296 GND.t69 5.26646
R24140 GND.n294 GND.t58 5.26646
R24141 GND.n294 GND.t47 5.26646
R24142 GND.n339 GND.t43 5.26646
R24143 GND.n339 GND.t77 5.26646
R24144 GND.n337 GND.t42 5.26646
R24145 GND.n337 GND.t70 5.26646
R24146 GND.n383 GND.t62 5.26646
R24147 GND.n383 GND.t56 5.26646
R24148 GND.n381 GND.t75 5.26646
R24149 GND.n381 GND.t60 5.26646
R24150 GND.t27 GND.n4555 4.98048
R24151 GND.n4100 GND.t24 4.98048
R24152 GND.n130 GND.n42 4.7699
R24153 GND.n405 GND.n404 4.7699
R24154 GND.n6875 GND.n6874 4.74817
R24155 GND.n6823 GND.n6822 4.74817
R24156 GND.n6857 GND.n6856 4.74817
R24157 GND.n6835 GND.n6824 4.74817
R24158 GND.n6874 GND.n6873 4.74817
R24159 GND.n6822 GND.n3757 4.74817
R24160 GND.n6858 GND.n6857 4.74817
R24161 GND.n6855 GND.n6824 4.74817
R24162 GND.n2823 GND.n2822 4.74817
R24163 GND.n2806 GND.n2110 4.74817
R24164 GND.n2783 GND.n2109 4.74817
R24165 GND.n2786 GND.n2108 4.74817
R24166 GND.n2823 GND.n2112 4.74817
R24167 GND.n2138 GND.n2110 4.74817
R24168 GND.n2805 GND.n2109 4.74817
R24169 GND.n2784 GND.n2108 4.74817
R24170 GND.n2674 GND.n2672 4.74817
R24171 GND.n2812 GND.n2811 4.74817
R24172 GND.n2150 GND.n2149 4.74817
R24173 GND.n2796 GND.n2795 4.74817
R24174 GND.n2182 GND.n2151 4.74817
R24175 GND.n6813 GND.n3743 4.74817
R24176 GND.n6864 GND.n3742 4.74817
R24177 GND.n6841 GND.n3741 4.74817
R24178 GND.n6845 GND.n3740 4.74817
R24179 GND.n3739 GND.n3738 4.74817
R24180 GND.n2672 GND.n2127 4.74817
R24181 GND.n2813 GND.n2812 4.74817
R24182 GND.n2149 GND.n2128 4.74817
R24183 GND.n2797 GND.n2796 4.74817
R24184 GND.n2794 GND.n2151 4.74817
R24185 GND.n3747 GND.n3743 4.74817
R24186 GND.n6814 GND.n3742 4.74817
R24187 GND.n6863 GND.n3741 4.74817
R24188 GND.n6842 GND.n3740 4.74817
R24189 GND.n6846 GND.n3739 4.74817
R24190 GND.n129 GND.n128 4.7074
R24191 GND.n361 GND.n360 4.7074
R24192 GND.n194 GND.n192 4.69785
R24193 GND.n182 GND.n180 4.69785
R24194 GND.n170 GND.n168 4.69785
R24195 GND.n158 GND.n156 4.69785
R24196 GND.n146 GND.n144 4.69785
R24197 GND.n135 GND.n133 4.69785
R24198 GND.n265 GND.n263 4.69785
R24199 GND.n253 GND.n251 4.69785
R24200 GND.n241 GND.n239 4.69785
R24201 GND.n229 GND.n227 4.69785
R24202 GND.n217 GND.n215 4.69785
R24203 GND.n206 GND.n204 4.69785
R24204 GND.n6292 GND.n6289 4.6132
R24205 GND.n7905 GND.n1793 4.6132
R24206 GND.n3009 GND.n3001 4.5974
R24207 GND.n4839 GND.n4652 4.5974
R24208 GND.n4970 GND.n4601 4.5974
R24209 GND.n4578 GND.n4566 4.5974
R24210 GND.n5128 GND.n4513 4.5974
R24211 GND.n5133 GND.n4480 4.5974
R24212 GND.n5295 GND.n5294 4.5974
R24213 GND.n5283 GND.n4395 4.5974
R24214 GND.n5455 GND.n4344 4.5974
R24215 GND.n4320 GND.n4308 4.5974
R24216 GND.n5615 GND.n4259 4.5974
R24217 GND.n5696 GND.n4225 4.5974
R24218 GND.n5835 GND.n4166 4.5974
R24219 GND.n4151 GND.n4139 4.5974
R24220 GND.n5941 GND.n4088 4.5974
R24221 GND.n4064 GND.n4052 4.5974
R24222 GND.n6350 GND.n6348 4.5974
R24223 GND.n7341 GND.n3230 4.5974
R24224 GND.n6208 GND.n6195 4.46111
R24225 GND.n52 GND.n48 4.40546
R24226 GND.n75 GND.n71 4.40546
R24227 GND.n95 GND.n91 4.40546
R24228 GND.n118 GND.n114 4.40546
R24229 GND.n9 GND.n5 4.40546
R24230 GND.n32 GND.n28 4.40546
R24231 GND.n307 GND.n303 4.40546
R24232 GND.n284 GND.n280 4.40546
R24233 GND.n350 GND.n346 4.40546
R24234 GND.n327 GND.n323 4.40546
R24235 GND.n394 GND.n390 4.40546
R24236 GND.n371 GND.n367 4.40546
R24237 GND.n274 GND.n202 4.40059
R24238 GND.n6176 GND.n6137 4.05904
R24239 GND.n4773 GND.n4772 4.05904
R24240 GND.n4757 GND.n4756 4.05904
R24241 GND.n6222 GND.n6221 4.05904
R24242 GND.n274 GND.n273 3.60163
R24243 GND.n61 GND.n43 3.49141
R24244 GND.n84 GND.n66 3.49141
R24245 GND.n104 GND.n86 3.49141
R24246 GND.n127 GND.n109 3.49141
R24247 GND.n18 GND.n0 3.49141
R24248 GND.n41 GND.n23 3.49141
R24249 GND.n316 GND.n298 3.49141
R24250 GND.n293 GND.n275 3.49141
R24251 GND.n359 GND.n341 3.49141
R24252 GND.n336 GND.n318 3.49141
R24253 GND.n403 GND.n385 3.49141
R24254 GND.n380 GND.n362 3.49141
R24255 GND.n5374 GND.t4 3.44818
R24256 GND.n5639 GND.t6 3.44818
R24257 GND.n4812 GND.t157 3.0651
R24258 GND.n2992 GND.n1839 3.0651
R24259 GND.n7567 GND.t135 3.0651
R24260 GND.n4913 GND.n4648 3.0651
R24261 GND.n4977 GND.n4606 3.0651
R24262 GND.n5076 GND.n4562 3.0651
R24263 GND.n5123 GND.n4523 3.0651
R24264 GND.n5236 GND.n4476 3.0651
R24265 GND.n5302 GND.n4434 3.0651
R24266 GND.n5398 GND.n4390 3.0651
R24267 GND.n5462 GND.n4349 3.0651
R24268 GND.n5569 GND.n4304 3.0651
R24269 GND.n5622 GND.n4263 3.0651
R24270 GND.n5708 GND.n5707 3.0651
R24271 GND.n5820 GND.n4170 3.0651
R24272 GND.n5884 GND.n4135 3.0651
R24273 GND.n5948 GND.n4093 3.0651
R24274 GND.n6035 GND.n4047 3.0651
R24275 GND.n4014 GND.n4004 3.0651
R24276 GND.t125 GND.n3973 3.0651
R24277 GND.n7335 GND.n3241 3.0651
R24278 GND.n7302 GND.t88 3.0651
R24279 GND.n59 GND.n58 2.71565
R24280 GND.n82 GND.n81 2.71565
R24281 GND.n102 GND.n101 2.71565
R24282 GND.n125 GND.n124 2.71565
R24283 GND.n16 GND.n15 2.71565
R24284 GND.n39 GND.n38 2.71565
R24285 GND.n314 GND.n313 2.71565
R24286 GND.n291 GND.n290 2.71565
R24287 GND.n357 GND.n356 2.71565
R24288 GND.n334 GND.n333 2.71565
R24289 GND.n401 GND.n400 2.71565
R24290 GND.n378 GND.n377 2.71565
R24291 GND.n85 GND.n65 2.69878
R24292 GND.n65 GND.n63 2.69878
R24293 GND.n128 GND.n108 2.69878
R24294 GND.n108 GND.n106 2.69878
R24295 GND.n42 GND.n22 2.69878
R24296 GND.n22 GND.n20 2.69878
R24297 GND.n297 GND.n295 2.69878
R24298 GND.n317 GND.n297 2.69878
R24299 GND.n340 GND.n338 2.69878
R24300 GND.n360 GND.n340 2.69878
R24301 GND.n384 GND.n382 2.69878
R24302 GND.n404 GND.n384 2.69878
R24303 GND.n7321 GND.t167 2.29895
R24304 GND.n6874 GND.n3744 2.27742
R24305 GND.n6822 GND.n3744 2.27742
R24306 GND.n6857 GND.n3744 2.27742
R24307 GND.n6824 GND.n3744 2.27742
R24308 GND.n2824 GND.n2823 2.27742
R24309 GND.n2824 GND.n2110 2.27742
R24310 GND.n2824 GND.n2109 2.27742
R24311 GND.n2824 GND.n2108 2.27742
R24312 GND.n2812 GND.n2107 2.27742
R24313 GND.n2149 GND.n2107 2.27742
R24314 GND.n2796 GND.n2107 2.27742
R24315 GND.n2151 GND.n2107 2.27742
R24316 GND.n6881 GND.n3743 2.27742
R24317 GND.n6881 GND.n3742 2.27742
R24318 GND.n6881 GND.n3741 2.27742
R24319 GND.n6881 GND.n3740 2.27742
R24320 GND.n6881 GND.n3739 2.27742
R24321 GND.n2672 GND.n2107 2.27742
R24322 GND GND.n131 2.17817
R24323 GND.n130 GND.n129 1.96602
R24324 GND.n405 GND.n361 1.96602
R24325 GND.n55 GND.n45 1.93989
R24326 GND.n78 GND.n68 1.93989
R24327 GND.n98 GND.n88 1.93989
R24328 GND.n121 GND.n111 1.93989
R24329 GND.n12 GND.n2 1.93989
R24330 GND.n35 GND.n25 1.93989
R24331 GND.n310 GND.n300 1.93989
R24332 GND.n287 GND.n277 1.93989
R24333 GND.n353 GND.n343 1.93989
R24334 GND.n330 GND.n320 1.93989
R24335 GND.n397 GND.n387 1.93989
R24336 GND.n374 GND.n364 1.93989
R24337 GND.n201 GND.n191 1.93989
R24338 GND.n189 GND.n179 1.93989
R24339 GND.n177 GND.n167 1.93989
R24340 GND.n165 GND.n155 1.93989
R24341 GND.n153 GND.n143 1.93989
R24342 GND.n142 GND.n132 1.93989
R24343 GND.n272 GND.n262 1.93989
R24344 GND.n260 GND.n250 1.93989
R24345 GND.n248 GND.n238 1.93989
R24346 GND.n236 GND.n226 1.93989
R24347 GND.n224 GND.n214 1.93989
R24348 GND.n213 GND.n203 1.93989
R24349 GND.n4812 GND.n2971 1.5328
R24350 GND.n2989 GND.n2983 1.5328
R24351 GND.n7866 GND.n1839 1.5328
R24352 GND.n4919 GND.n4635 1.5328
R24353 GND.n4946 GND.n4620 1.5328
R24354 GND.n5082 GND.n4550 1.5328
R24355 GND.n4539 GND.n4527 1.5328
R24356 GND.n5242 GND.n4463 1.5328
R24357 GND.n5269 GND.n4439 1.5328
R24358 GND.n5404 GND.n4378 1.5328
R24359 GND.n5431 GND.n4354 1.5328
R24360 GND.n5575 GND.n4292 1.5328
R24361 GND.n5602 GND.n4268 1.5328
R24362 GND.n4213 GND.n4212 1.5328
R24363 GND.n5801 GND.n5800 1.5328
R24364 GND.n5890 GND.n4122 1.5328
R24365 GND.n5917 GND.n4107 1.5328
R24366 GND.n6041 GND.n4036 1.5328
R24367 GND.n6066 GND.n4024 1.5328
R24368 GND.n6415 GND.n3241 1.5328
R24369 GND.n7328 GND.n7327 1.5328
R24370 GND.n3273 GND.n3271 1.5328
R24371 GND.n166 GND.n154 1.47434
R24372 GND.n178 GND.n166 1.47434
R24373 GND.n190 GND.n178 1.47434
R24374 GND.n202 GND.n190 1.47434
R24375 GND.n237 GND.n225 1.47434
R24376 GND.n249 GND.n237 1.47434
R24377 GND.n261 GND.n249 1.47434
R24378 GND.n273 GND.n261 1.47434
R24379 GND.n9696 GND.n9695 1.2189
R24380 GND.n54 GND.n47 1.16414
R24381 GND.n77 GND.n70 1.16414
R24382 GND.n97 GND.n90 1.16414
R24383 GND.n120 GND.n113 1.16414
R24384 GND.n11 GND.n4 1.16414
R24385 GND.n34 GND.n27 1.16414
R24386 GND.n309 GND.n302 1.16414
R24387 GND.n286 GND.n279 1.16414
R24388 GND.n352 GND.n345 1.16414
R24389 GND.n329 GND.n322 1.16414
R24390 GND.n396 GND.n389 1.16414
R24391 GND.n373 GND.n366 1.16414
R24392 GND.n199 GND.n198 1.16414
R24393 GND.n187 GND.n186 1.16414
R24394 GND.n175 GND.n174 1.16414
R24395 GND.n163 GND.n162 1.16414
R24396 GND.n151 GND.n150 1.16414
R24397 GND.n140 GND.n139 1.16414
R24398 GND.n270 GND.n269 1.16414
R24399 GND.n258 GND.n257 1.16414
R24400 GND.n246 GND.n245 1.16414
R24401 GND.n234 GND.n233 1.16414
R24402 GND.n222 GND.n221 1.16414
R24403 GND.n211 GND.n210 1.16414
R24404 GND.n4355 GND.t29 1.14973
R24405 GND.t17 GND.n4303 1.14973
R24406 GND.n6425 GND.n3969 0.776258
R24407 GND.n3042 GND.n3041 0.776258
R24408 GND.t2 GND.n5082 0.76665
R24409 GND.n4107 GND.t10 0.76665
R24410 GND.n6881 GND.n3744 0.54525
R24411 GND.n2824 GND.n2107 0.54525
R24412 GND.n6267 GND.n3361 0.518793
R24413 GND.n1535 GND.n1475 0.518793
R24414 GND.n9609 GND.n9608 0.518793
R24415 GND.n7921 GND.n7920 0.518793
R24416 GND.n9615 GND.n473 0.489829
R24417 GND.n2410 GND.n2409 0.489829
R24418 GND GND.n9696 0.482093
R24419 GND.n8288 GND.n8287 0.471537
R24420 GND.n9319 GND.n697 0.471537
R24421 GND.n9460 GND.n9459 0.471537
R24422 GND.n8175 GND.n8174 0.471537
R24423 GND.n7344 GND.n3227 0.46239
R24424 GND.n3051 GND.n3050 0.46239
R24425 GND.n51 GND.n50 0.388379
R24426 GND.n74 GND.n73 0.388379
R24427 GND.n94 GND.n93 0.388379
R24428 GND.n117 GND.n116 0.388379
R24429 GND.n8 GND.n7 0.388379
R24430 GND.n31 GND.n30 0.388379
R24431 GND.n306 GND.n305 0.388379
R24432 GND.n283 GND.n282 0.388379
R24433 GND.n349 GND.n348 0.388379
R24434 GND.n326 GND.n325 0.388379
R24435 GND.n393 GND.n392 0.388379
R24436 GND.n370 GND.n369 0.388379
R24437 GND.n195 GND.n193 0.388379
R24438 GND.n183 GND.n181 0.388379
R24439 GND.n171 GND.n169 0.388379
R24440 GND.n159 GND.n157 0.388379
R24441 GND.n147 GND.n145 0.388379
R24442 GND.n136 GND.n134 0.388379
R24443 GND.n266 GND.n264 0.388379
R24444 GND.n254 GND.n252 0.388379
R24445 GND.n242 GND.n240 0.388379
R24446 GND.n230 GND.n228 0.388379
R24447 GND.n218 GND.n216 0.388379
R24448 GND.n207 GND.n205 0.388379
R24449 GND.n5163 GND.t19 0.383575
R24450 GND.n5861 GND.t14 0.383575
R24451 GND.n6430 GND.n6429 0.296232
R24452 GND.n7834 GND.n7833 0.296232
R24453 GND.n6327 GND.n6323 0.285561
R24454 GND.n8101 GND.n8099 0.285561
R24455 GND.n9529 GND.n515 0.285561
R24456 GND.n7884 GND.n1768 0.285561
R24457 GND.n9564 GND.n9529 0.256598
R24458 GND.n8099 GND.n8098 0.256598
R24459 GND.n9696 GND.n274 0.231583
R24460 GND.n6289 GND.n6288 0.229039
R24461 GND.n6289 GND.n6117 0.229039
R24462 GND.n1793 GND.n1788 0.229039
R24463 GND.n7903 GND.n1793 0.229039
R24464 GND.n4664 GND.n1834 0.224585
R24465 GND.n6329 GND.n6328 0.224585
R24466 GND.n60 GND.n44 0.155672
R24467 GND.n53 GND.n44 0.155672
R24468 GND.n53 GND.n52 0.155672
R24469 GND.n83 GND.n67 0.155672
R24470 GND.n76 GND.n67 0.155672
R24471 GND.n76 GND.n75 0.155672
R24472 GND.n103 GND.n87 0.155672
R24473 GND.n96 GND.n87 0.155672
R24474 GND.n96 GND.n95 0.155672
R24475 GND.n126 GND.n110 0.155672
R24476 GND.n119 GND.n110 0.155672
R24477 GND.n119 GND.n118 0.155672
R24478 GND.n17 GND.n1 0.155672
R24479 GND.n10 GND.n1 0.155672
R24480 GND.n10 GND.n9 0.155672
R24481 GND.n40 GND.n24 0.155672
R24482 GND.n33 GND.n24 0.155672
R24483 GND.n33 GND.n32 0.155672
R24484 GND.n315 GND.n299 0.155672
R24485 GND.n308 GND.n299 0.155672
R24486 GND.n308 GND.n307 0.155672
R24487 GND.n292 GND.n276 0.155672
R24488 GND.n285 GND.n276 0.155672
R24489 GND.n285 GND.n284 0.155672
R24490 GND.n358 GND.n342 0.155672
R24491 GND.n351 GND.n342 0.155672
R24492 GND.n351 GND.n350 0.155672
R24493 GND.n335 GND.n319 0.155672
R24494 GND.n328 GND.n319 0.155672
R24495 GND.n328 GND.n327 0.155672
R24496 GND.n402 GND.n386 0.155672
R24497 GND.n395 GND.n386 0.155672
R24498 GND.n395 GND.n394 0.155672
R24499 GND.n379 GND.n363 0.155672
R24500 GND.n372 GND.n363 0.155672
R24501 GND.n372 GND.n371 0.155672
R24502 GND.n200 GND.n192 0.155672
R24503 GND.n188 GND.n180 0.155672
R24504 GND.n176 GND.n168 0.155672
R24505 GND.n164 GND.n156 0.155672
R24506 GND.n152 GND.n144 0.155672
R24507 GND.n141 GND.n133 0.155672
R24508 GND.n271 GND.n263 0.155672
R24509 GND.n259 GND.n251 0.155672
R24510 GND.n247 GND.n239 0.155672
R24511 GND.n235 GND.n227 0.155672
R24512 GND.n223 GND.n215 0.155672
R24513 GND.n212 GND.n204 0.155672
R24514 GND.n4665 GND.n4664 0.152939
R24515 GND.n4666 GND.n4665 0.152939
R24516 GND.n4666 GND.n4657 0.152939
R24517 GND.n4859 GND.n4657 0.152939
R24518 GND.n4860 GND.n4859 0.152939
R24519 GND.n4861 GND.n4860 0.152939
R24520 GND.n4862 GND.n4861 0.152939
R24521 GND.n4863 GND.n4862 0.152939
R24522 GND.n4865 GND.n4863 0.152939
R24523 GND.n4866 GND.n4865 0.152939
R24524 GND.n4867 GND.n4866 0.152939
R24525 GND.n4868 GND.n4867 0.152939
R24526 GND.n4869 GND.n4868 0.152939
R24527 GND.n4870 GND.n4869 0.152939
R24528 GND.n4871 GND.n4870 0.152939
R24529 GND.n4872 GND.n4871 0.152939
R24530 GND.n4872 GND.n4586 0.152939
R24531 GND.n5003 GND.n4586 0.152939
R24532 GND.n5004 GND.n5003 0.152939
R24533 GND.n5005 GND.n5004 0.152939
R24534 GND.n5006 GND.n5005 0.152939
R24535 GND.n5007 GND.n5006 0.152939
R24536 GND.n5008 GND.n5007 0.152939
R24537 GND.n5009 GND.n5008 0.152939
R24538 GND.n5012 GND.n5009 0.152939
R24539 GND.n5013 GND.n5012 0.152939
R24540 GND.n5014 GND.n5013 0.152939
R24541 GND.n5015 GND.n5014 0.152939
R24542 GND.n5016 GND.n5015 0.152939
R24543 GND.n5017 GND.n5016 0.152939
R24544 GND.n5018 GND.n5017 0.152939
R24545 GND.n5019 GND.n5018 0.152939
R24546 GND.n5020 GND.n5019 0.152939
R24547 GND.n5020 GND.n4500 0.152939
R24548 GND.n5166 GND.n4500 0.152939
R24549 GND.n5167 GND.n5166 0.152939
R24550 GND.n5168 GND.n5167 0.152939
R24551 GND.n5169 GND.n5168 0.152939
R24552 GND.n5170 GND.n5169 0.152939
R24553 GND.n5171 GND.n5170 0.152939
R24554 GND.n5172 GND.n5171 0.152939
R24555 GND.n5175 GND.n5172 0.152939
R24556 GND.n5176 GND.n5175 0.152939
R24557 GND.n5177 GND.n5176 0.152939
R24558 GND.n5178 GND.n5177 0.152939
R24559 GND.n5179 GND.n5178 0.152939
R24560 GND.n5180 GND.n5179 0.152939
R24561 GND.n5181 GND.n5180 0.152939
R24562 GND.n5182 GND.n5181 0.152939
R24563 GND.n5183 GND.n5182 0.152939
R24564 GND.n5183 GND.n4414 0.152939
R24565 GND.n5327 GND.n4414 0.152939
R24566 GND.n5328 GND.n5327 0.152939
R24567 GND.n5329 GND.n5328 0.152939
R24568 GND.n5330 GND.n5329 0.152939
R24569 GND.n5331 GND.n5330 0.152939
R24570 GND.n5332 GND.n5331 0.152939
R24571 GND.n5333 GND.n5332 0.152939
R24572 GND.n5336 GND.n5333 0.152939
R24573 GND.n5337 GND.n5336 0.152939
R24574 GND.n5338 GND.n5337 0.152939
R24575 GND.n5339 GND.n5338 0.152939
R24576 GND.n5340 GND.n5339 0.152939
R24577 GND.n5341 GND.n5340 0.152939
R24578 GND.n5342 GND.n5341 0.152939
R24579 GND.n5343 GND.n5342 0.152939
R24580 GND.n5344 GND.n5343 0.152939
R24581 GND.n5344 GND.n4328 0.152939
R24582 GND.n5487 GND.n4328 0.152939
R24583 GND.n5488 GND.n5487 0.152939
R24584 GND.n5489 GND.n5488 0.152939
R24585 GND.n5490 GND.n5489 0.152939
R24586 GND.n5491 GND.n5490 0.152939
R24587 GND.n5492 GND.n5491 0.152939
R24588 GND.n5493 GND.n5492 0.152939
R24589 GND.n5497 GND.n5493 0.152939
R24590 GND.n5498 GND.n5497 0.152939
R24591 GND.n5499 GND.n5498 0.152939
R24592 GND.n5500 GND.n5499 0.152939
R24593 GND.n5501 GND.n5500 0.152939
R24594 GND.n5502 GND.n5501 0.152939
R24595 GND.n5503 GND.n5502 0.152939
R24596 GND.n5504 GND.n5503 0.152939
R24597 GND.n5505 GND.n5504 0.152939
R24598 GND.n5506 GND.n5505 0.152939
R24599 GND.n5507 GND.n5506 0.152939
R24600 GND.n5508 GND.n5507 0.152939
R24601 GND.n5509 GND.n5508 0.152939
R24602 GND.n5509 GND.n4222 0.152939
R24603 GND.n5699 GND.n4222 0.152939
R24604 GND.n5700 GND.n5699 0.152939
R24605 GND.n5701 GND.n5700 0.152939
R24606 GND.n5702 GND.n5701 0.152939
R24607 GND.n5702 GND.n4198 0.152939
R24608 GND.n5733 GND.n4198 0.152939
R24609 GND.n5734 GND.n5733 0.152939
R24610 GND.n5735 GND.n5734 0.152939
R24611 GND.n5736 GND.n5735 0.152939
R24612 GND.n5737 GND.n5736 0.152939
R24613 GND.n5738 GND.n5737 0.152939
R24614 GND.n5739 GND.n5738 0.152939
R24615 GND.n5742 GND.n5739 0.152939
R24616 GND.n5743 GND.n5742 0.152939
R24617 GND.n5744 GND.n5743 0.152939
R24618 GND.n5745 GND.n5744 0.152939
R24619 GND.n5746 GND.n5745 0.152939
R24620 GND.n5747 GND.n5746 0.152939
R24621 GND.n5748 GND.n5747 0.152939
R24622 GND.n5749 GND.n5748 0.152939
R24623 GND.n5752 GND.n5749 0.152939
R24624 GND.n5753 GND.n5752 0.152939
R24625 GND.n5754 GND.n5753 0.152939
R24626 GND.n5755 GND.n5754 0.152939
R24627 GND.n5756 GND.n5755 0.152939
R24628 GND.n5757 GND.n5756 0.152939
R24629 GND.n5758 GND.n5757 0.152939
R24630 GND.n5759 GND.n5758 0.152939
R24631 GND.n5760 GND.n5759 0.152939
R24632 GND.n5760 GND.n4072 0.152939
R24633 GND.n5973 GND.n4072 0.152939
R24634 GND.n5974 GND.n5973 0.152939
R24635 GND.n5975 GND.n5974 0.152939
R24636 GND.n5976 GND.n5975 0.152939
R24637 GND.n5977 GND.n5976 0.152939
R24638 GND.n5978 GND.n5977 0.152939
R24639 GND.n5979 GND.n5978 0.152939
R24640 GND.n5982 GND.n5979 0.152939
R24641 GND.n5983 GND.n5982 0.152939
R24642 GND.n5984 GND.n5983 0.152939
R24643 GND.n5985 GND.n5984 0.152939
R24644 GND.n5986 GND.n5985 0.152939
R24645 GND.n5986 GND.n4008 0.152939
R24646 GND.n6098 GND.n4008 0.152939
R24647 GND.n6099 GND.n6098 0.152939
R24648 GND.n6100 GND.n6099 0.152939
R24649 GND.n6101 GND.n6100 0.152939
R24650 GND.n6102 GND.n6101 0.152939
R24651 GND.n6103 GND.n6102 0.152939
R24652 GND.n6104 GND.n6103 0.152939
R24653 GND.n6105 GND.n6104 0.152939
R24654 GND.n6329 GND.n6105 0.152939
R24655 GND.n8289 GND.n8288 0.152939
R24656 GND.n8289 GND.n1315 0.152939
R24657 GND.n8297 GND.n1315 0.152939
R24658 GND.n8298 GND.n8297 0.152939
R24659 GND.n8299 GND.n8298 0.152939
R24660 GND.n8299 GND.n1309 0.152939
R24661 GND.n8307 GND.n1309 0.152939
R24662 GND.n8308 GND.n8307 0.152939
R24663 GND.n8309 GND.n8308 0.152939
R24664 GND.n8309 GND.n1303 0.152939
R24665 GND.n8317 GND.n1303 0.152939
R24666 GND.n8318 GND.n8317 0.152939
R24667 GND.n8319 GND.n8318 0.152939
R24668 GND.n8319 GND.n1297 0.152939
R24669 GND.n8327 GND.n1297 0.152939
R24670 GND.n8328 GND.n8327 0.152939
R24671 GND.n8329 GND.n8328 0.152939
R24672 GND.n8329 GND.n1291 0.152939
R24673 GND.n8337 GND.n1291 0.152939
R24674 GND.n8338 GND.n8337 0.152939
R24675 GND.n8339 GND.n8338 0.152939
R24676 GND.n8339 GND.n1285 0.152939
R24677 GND.n8347 GND.n1285 0.152939
R24678 GND.n8348 GND.n8347 0.152939
R24679 GND.n8349 GND.n8348 0.152939
R24680 GND.n8349 GND.n1279 0.152939
R24681 GND.n8357 GND.n1279 0.152939
R24682 GND.n8358 GND.n8357 0.152939
R24683 GND.n8359 GND.n8358 0.152939
R24684 GND.n8359 GND.n1273 0.152939
R24685 GND.n8367 GND.n1273 0.152939
R24686 GND.n8368 GND.n8367 0.152939
R24687 GND.n8369 GND.n8368 0.152939
R24688 GND.n8369 GND.n1267 0.152939
R24689 GND.n8377 GND.n1267 0.152939
R24690 GND.n8378 GND.n8377 0.152939
R24691 GND.n8379 GND.n8378 0.152939
R24692 GND.n8379 GND.n1261 0.152939
R24693 GND.n8387 GND.n1261 0.152939
R24694 GND.n8388 GND.n8387 0.152939
R24695 GND.n8389 GND.n8388 0.152939
R24696 GND.n8389 GND.n1255 0.152939
R24697 GND.n8397 GND.n1255 0.152939
R24698 GND.n8398 GND.n8397 0.152939
R24699 GND.n8399 GND.n8398 0.152939
R24700 GND.n8399 GND.n1249 0.152939
R24701 GND.n8407 GND.n1249 0.152939
R24702 GND.n8408 GND.n8407 0.152939
R24703 GND.n8409 GND.n8408 0.152939
R24704 GND.n8409 GND.n1243 0.152939
R24705 GND.n8417 GND.n1243 0.152939
R24706 GND.n8418 GND.n8417 0.152939
R24707 GND.n8419 GND.n8418 0.152939
R24708 GND.n8419 GND.n1237 0.152939
R24709 GND.n8427 GND.n1237 0.152939
R24710 GND.n8428 GND.n8427 0.152939
R24711 GND.n8429 GND.n8428 0.152939
R24712 GND.n8429 GND.n1231 0.152939
R24713 GND.n8437 GND.n1231 0.152939
R24714 GND.n8438 GND.n8437 0.152939
R24715 GND.n8439 GND.n8438 0.152939
R24716 GND.n8439 GND.n1225 0.152939
R24717 GND.n8447 GND.n1225 0.152939
R24718 GND.n8448 GND.n8447 0.152939
R24719 GND.n8449 GND.n8448 0.152939
R24720 GND.n8449 GND.n1219 0.152939
R24721 GND.n8457 GND.n1219 0.152939
R24722 GND.n8458 GND.n8457 0.152939
R24723 GND.n8459 GND.n8458 0.152939
R24724 GND.n8459 GND.n1213 0.152939
R24725 GND.n8467 GND.n1213 0.152939
R24726 GND.n8468 GND.n8467 0.152939
R24727 GND.n8469 GND.n8468 0.152939
R24728 GND.n8469 GND.n1207 0.152939
R24729 GND.n8477 GND.n1207 0.152939
R24730 GND.n8478 GND.n8477 0.152939
R24731 GND.n8479 GND.n8478 0.152939
R24732 GND.n8479 GND.n1201 0.152939
R24733 GND.n8487 GND.n1201 0.152939
R24734 GND.n8488 GND.n8487 0.152939
R24735 GND.n8489 GND.n8488 0.152939
R24736 GND.n8489 GND.n1195 0.152939
R24737 GND.n8497 GND.n1195 0.152939
R24738 GND.n8498 GND.n8497 0.152939
R24739 GND.n8499 GND.n8498 0.152939
R24740 GND.n8499 GND.n1189 0.152939
R24741 GND.n8507 GND.n1189 0.152939
R24742 GND.n8508 GND.n8507 0.152939
R24743 GND.n8509 GND.n8508 0.152939
R24744 GND.n8509 GND.n1183 0.152939
R24745 GND.n8517 GND.n1183 0.152939
R24746 GND.n8518 GND.n8517 0.152939
R24747 GND.n8519 GND.n8518 0.152939
R24748 GND.n8519 GND.n1177 0.152939
R24749 GND.n8527 GND.n1177 0.152939
R24750 GND.n8528 GND.n8527 0.152939
R24751 GND.n8529 GND.n8528 0.152939
R24752 GND.n8529 GND.n1171 0.152939
R24753 GND.n8537 GND.n1171 0.152939
R24754 GND.n8538 GND.n8537 0.152939
R24755 GND.n8539 GND.n8538 0.152939
R24756 GND.n8539 GND.n1165 0.152939
R24757 GND.n8547 GND.n1165 0.152939
R24758 GND.n8548 GND.n8547 0.152939
R24759 GND.n8549 GND.n8548 0.152939
R24760 GND.n8549 GND.n1159 0.152939
R24761 GND.n8557 GND.n1159 0.152939
R24762 GND.n8558 GND.n8557 0.152939
R24763 GND.n8559 GND.n8558 0.152939
R24764 GND.n8559 GND.n1153 0.152939
R24765 GND.n8567 GND.n1153 0.152939
R24766 GND.n8568 GND.n8567 0.152939
R24767 GND.n8569 GND.n8568 0.152939
R24768 GND.n8569 GND.n1147 0.152939
R24769 GND.n8577 GND.n1147 0.152939
R24770 GND.n8578 GND.n8577 0.152939
R24771 GND.n8579 GND.n8578 0.152939
R24772 GND.n8579 GND.n1141 0.152939
R24773 GND.n8587 GND.n1141 0.152939
R24774 GND.n8588 GND.n8587 0.152939
R24775 GND.n8589 GND.n8588 0.152939
R24776 GND.n8589 GND.n1135 0.152939
R24777 GND.n8597 GND.n1135 0.152939
R24778 GND.n8598 GND.n8597 0.152939
R24779 GND.n8599 GND.n8598 0.152939
R24780 GND.n8599 GND.n1129 0.152939
R24781 GND.n8607 GND.n1129 0.152939
R24782 GND.n8608 GND.n8607 0.152939
R24783 GND.n8609 GND.n8608 0.152939
R24784 GND.n8609 GND.n1123 0.152939
R24785 GND.n8617 GND.n1123 0.152939
R24786 GND.n8618 GND.n8617 0.152939
R24787 GND.n8619 GND.n8618 0.152939
R24788 GND.n8619 GND.n1117 0.152939
R24789 GND.n8627 GND.n1117 0.152939
R24790 GND.n8628 GND.n8627 0.152939
R24791 GND.n8629 GND.n8628 0.152939
R24792 GND.n8629 GND.n1111 0.152939
R24793 GND.n8637 GND.n1111 0.152939
R24794 GND.n8638 GND.n8637 0.152939
R24795 GND.n8639 GND.n8638 0.152939
R24796 GND.n8639 GND.n1105 0.152939
R24797 GND.n8647 GND.n1105 0.152939
R24798 GND.n8648 GND.n8647 0.152939
R24799 GND.n8649 GND.n8648 0.152939
R24800 GND.n8649 GND.n1099 0.152939
R24801 GND.n8657 GND.n1099 0.152939
R24802 GND.n8658 GND.n8657 0.152939
R24803 GND.n8659 GND.n8658 0.152939
R24804 GND.n8659 GND.n1093 0.152939
R24805 GND.n8667 GND.n1093 0.152939
R24806 GND.n8668 GND.n8667 0.152939
R24807 GND.n8669 GND.n8668 0.152939
R24808 GND.n8669 GND.n1087 0.152939
R24809 GND.n8677 GND.n1087 0.152939
R24810 GND.n8678 GND.n8677 0.152939
R24811 GND.n8679 GND.n8678 0.152939
R24812 GND.n8679 GND.n1081 0.152939
R24813 GND.n8687 GND.n1081 0.152939
R24814 GND.n8688 GND.n8687 0.152939
R24815 GND.n8689 GND.n8688 0.152939
R24816 GND.n8689 GND.n1075 0.152939
R24817 GND.n8697 GND.n1075 0.152939
R24818 GND.n8698 GND.n8697 0.152939
R24819 GND.n8699 GND.n8698 0.152939
R24820 GND.n8699 GND.n1069 0.152939
R24821 GND.n8707 GND.n1069 0.152939
R24822 GND.n8708 GND.n8707 0.152939
R24823 GND.n8709 GND.n8708 0.152939
R24824 GND.n8709 GND.n1063 0.152939
R24825 GND.n8717 GND.n1063 0.152939
R24826 GND.n8718 GND.n8717 0.152939
R24827 GND.n8719 GND.n8718 0.152939
R24828 GND.n8719 GND.n1057 0.152939
R24829 GND.n8727 GND.n1057 0.152939
R24830 GND.n8728 GND.n8727 0.152939
R24831 GND.n8729 GND.n8728 0.152939
R24832 GND.n8729 GND.n1051 0.152939
R24833 GND.n8737 GND.n1051 0.152939
R24834 GND.n8738 GND.n8737 0.152939
R24835 GND.n8739 GND.n8738 0.152939
R24836 GND.n8739 GND.n1045 0.152939
R24837 GND.n8747 GND.n1045 0.152939
R24838 GND.n8748 GND.n8747 0.152939
R24839 GND.n8749 GND.n8748 0.152939
R24840 GND.n8749 GND.n1039 0.152939
R24841 GND.n8757 GND.n1039 0.152939
R24842 GND.n8758 GND.n8757 0.152939
R24843 GND.n8759 GND.n8758 0.152939
R24844 GND.n8759 GND.n1033 0.152939
R24845 GND.n8767 GND.n1033 0.152939
R24846 GND.n8768 GND.n8767 0.152939
R24847 GND.n8769 GND.n8768 0.152939
R24848 GND.n8769 GND.n1027 0.152939
R24849 GND.n8777 GND.n1027 0.152939
R24850 GND.n8778 GND.n8777 0.152939
R24851 GND.n8779 GND.n8778 0.152939
R24852 GND.n8779 GND.n1021 0.152939
R24853 GND.n8787 GND.n1021 0.152939
R24854 GND.n8788 GND.n8787 0.152939
R24855 GND.n8789 GND.n8788 0.152939
R24856 GND.n8789 GND.n1015 0.152939
R24857 GND.n8797 GND.n1015 0.152939
R24858 GND.n8798 GND.n8797 0.152939
R24859 GND.n8799 GND.n8798 0.152939
R24860 GND.n8799 GND.n1009 0.152939
R24861 GND.n8807 GND.n1009 0.152939
R24862 GND.n8808 GND.n8807 0.152939
R24863 GND.n8809 GND.n8808 0.152939
R24864 GND.n8809 GND.n1003 0.152939
R24865 GND.n8817 GND.n1003 0.152939
R24866 GND.n8818 GND.n8817 0.152939
R24867 GND.n8819 GND.n8818 0.152939
R24868 GND.n8819 GND.n997 0.152939
R24869 GND.n8827 GND.n997 0.152939
R24870 GND.n8828 GND.n8827 0.152939
R24871 GND.n8829 GND.n8828 0.152939
R24872 GND.n8829 GND.n991 0.152939
R24873 GND.n8837 GND.n991 0.152939
R24874 GND.n8838 GND.n8837 0.152939
R24875 GND.n8839 GND.n8838 0.152939
R24876 GND.n8839 GND.n985 0.152939
R24877 GND.n8847 GND.n985 0.152939
R24878 GND.n8848 GND.n8847 0.152939
R24879 GND.n8849 GND.n8848 0.152939
R24880 GND.n8849 GND.n979 0.152939
R24881 GND.n8857 GND.n979 0.152939
R24882 GND.n8858 GND.n8857 0.152939
R24883 GND.n8859 GND.n8858 0.152939
R24884 GND.n8859 GND.n973 0.152939
R24885 GND.n8867 GND.n973 0.152939
R24886 GND.n8868 GND.n8867 0.152939
R24887 GND.n8869 GND.n8868 0.152939
R24888 GND.n8869 GND.n967 0.152939
R24889 GND.n8877 GND.n967 0.152939
R24890 GND.n8878 GND.n8877 0.152939
R24891 GND.n8879 GND.n8878 0.152939
R24892 GND.n8879 GND.n961 0.152939
R24893 GND.n8887 GND.n961 0.152939
R24894 GND.n8888 GND.n8887 0.152939
R24895 GND.n8889 GND.n8888 0.152939
R24896 GND.n8889 GND.n955 0.152939
R24897 GND.n8897 GND.n955 0.152939
R24898 GND.n8898 GND.n8897 0.152939
R24899 GND.n8899 GND.n8898 0.152939
R24900 GND.n8899 GND.n949 0.152939
R24901 GND.n8907 GND.n949 0.152939
R24902 GND.n8908 GND.n8907 0.152939
R24903 GND.n8909 GND.n8908 0.152939
R24904 GND.n8909 GND.n943 0.152939
R24905 GND.n8917 GND.n943 0.152939
R24906 GND.n8918 GND.n8917 0.152939
R24907 GND.n8919 GND.n8918 0.152939
R24908 GND.n8919 GND.n937 0.152939
R24909 GND.n8927 GND.n937 0.152939
R24910 GND.n8928 GND.n8927 0.152939
R24911 GND.n8929 GND.n8928 0.152939
R24912 GND.n8929 GND.n931 0.152939
R24913 GND.n8937 GND.n931 0.152939
R24914 GND.n8938 GND.n8937 0.152939
R24915 GND.n8939 GND.n8938 0.152939
R24916 GND.n8939 GND.n925 0.152939
R24917 GND.n8947 GND.n925 0.152939
R24918 GND.n8948 GND.n8947 0.152939
R24919 GND.n8949 GND.n8948 0.152939
R24920 GND.n8949 GND.n919 0.152939
R24921 GND.n8957 GND.n919 0.152939
R24922 GND.n8958 GND.n8957 0.152939
R24923 GND.n8959 GND.n8958 0.152939
R24924 GND.n8959 GND.n913 0.152939
R24925 GND.n8967 GND.n913 0.152939
R24926 GND.n8968 GND.n8967 0.152939
R24927 GND.n8969 GND.n8968 0.152939
R24928 GND.n8969 GND.n907 0.152939
R24929 GND.n8977 GND.n907 0.152939
R24930 GND.n8978 GND.n8977 0.152939
R24931 GND.n8979 GND.n8978 0.152939
R24932 GND.n8979 GND.n901 0.152939
R24933 GND.n8987 GND.n901 0.152939
R24934 GND.n8988 GND.n8987 0.152939
R24935 GND.n8989 GND.n8988 0.152939
R24936 GND.n8989 GND.n895 0.152939
R24937 GND.n8997 GND.n895 0.152939
R24938 GND.n8998 GND.n8997 0.152939
R24939 GND.n8999 GND.n8998 0.152939
R24940 GND.n8999 GND.n889 0.152939
R24941 GND.n9007 GND.n889 0.152939
R24942 GND.n9008 GND.n9007 0.152939
R24943 GND.n9009 GND.n9008 0.152939
R24944 GND.n9009 GND.n883 0.152939
R24945 GND.n9017 GND.n883 0.152939
R24946 GND.n9018 GND.n9017 0.152939
R24947 GND.n9019 GND.n9018 0.152939
R24948 GND.n9019 GND.n877 0.152939
R24949 GND.n9027 GND.n877 0.152939
R24950 GND.n9028 GND.n9027 0.152939
R24951 GND.n9029 GND.n9028 0.152939
R24952 GND.n9029 GND.n871 0.152939
R24953 GND.n9037 GND.n871 0.152939
R24954 GND.n9038 GND.n9037 0.152939
R24955 GND.n9039 GND.n9038 0.152939
R24956 GND.n9039 GND.n865 0.152939
R24957 GND.n9047 GND.n865 0.152939
R24958 GND.n9048 GND.n9047 0.152939
R24959 GND.n9049 GND.n9048 0.152939
R24960 GND.n9049 GND.n859 0.152939
R24961 GND.n9057 GND.n859 0.152939
R24962 GND.n9058 GND.n9057 0.152939
R24963 GND.n9059 GND.n9058 0.152939
R24964 GND.n9059 GND.n853 0.152939
R24965 GND.n9067 GND.n853 0.152939
R24966 GND.n9068 GND.n9067 0.152939
R24967 GND.n9069 GND.n9068 0.152939
R24968 GND.n9069 GND.n847 0.152939
R24969 GND.n9077 GND.n847 0.152939
R24970 GND.n9078 GND.n9077 0.152939
R24971 GND.n9079 GND.n9078 0.152939
R24972 GND.n9079 GND.n841 0.152939
R24973 GND.n9087 GND.n841 0.152939
R24974 GND.n9088 GND.n9087 0.152939
R24975 GND.n9089 GND.n9088 0.152939
R24976 GND.n9089 GND.n835 0.152939
R24977 GND.n9097 GND.n835 0.152939
R24978 GND.n9098 GND.n9097 0.152939
R24979 GND.n9099 GND.n9098 0.152939
R24980 GND.n9099 GND.n829 0.152939
R24981 GND.n9107 GND.n829 0.152939
R24982 GND.n9108 GND.n9107 0.152939
R24983 GND.n9109 GND.n9108 0.152939
R24984 GND.n9109 GND.n823 0.152939
R24985 GND.n9117 GND.n823 0.152939
R24986 GND.n9118 GND.n9117 0.152939
R24987 GND.n9119 GND.n9118 0.152939
R24988 GND.n9119 GND.n817 0.152939
R24989 GND.n9127 GND.n817 0.152939
R24990 GND.n9128 GND.n9127 0.152939
R24991 GND.n9129 GND.n9128 0.152939
R24992 GND.n9129 GND.n811 0.152939
R24993 GND.n9137 GND.n811 0.152939
R24994 GND.n9138 GND.n9137 0.152939
R24995 GND.n9139 GND.n9138 0.152939
R24996 GND.n9139 GND.n805 0.152939
R24997 GND.n9147 GND.n805 0.152939
R24998 GND.n9148 GND.n9147 0.152939
R24999 GND.n9149 GND.n9148 0.152939
R25000 GND.n9149 GND.n799 0.152939
R25001 GND.n9157 GND.n799 0.152939
R25002 GND.n9158 GND.n9157 0.152939
R25003 GND.n9159 GND.n9158 0.152939
R25004 GND.n9159 GND.n793 0.152939
R25005 GND.n9167 GND.n793 0.152939
R25006 GND.n9168 GND.n9167 0.152939
R25007 GND.n9169 GND.n9168 0.152939
R25008 GND.n9169 GND.n787 0.152939
R25009 GND.n9177 GND.n787 0.152939
R25010 GND.n9178 GND.n9177 0.152939
R25011 GND.n9179 GND.n9178 0.152939
R25012 GND.n9179 GND.n781 0.152939
R25013 GND.n9187 GND.n781 0.152939
R25014 GND.n9188 GND.n9187 0.152939
R25015 GND.n9189 GND.n9188 0.152939
R25016 GND.n9189 GND.n775 0.152939
R25017 GND.n9197 GND.n775 0.152939
R25018 GND.n9198 GND.n9197 0.152939
R25019 GND.n9199 GND.n9198 0.152939
R25020 GND.n9199 GND.n769 0.152939
R25021 GND.n9207 GND.n769 0.152939
R25022 GND.n9208 GND.n9207 0.152939
R25023 GND.n9209 GND.n9208 0.152939
R25024 GND.n9209 GND.n763 0.152939
R25025 GND.n9217 GND.n763 0.152939
R25026 GND.n9218 GND.n9217 0.152939
R25027 GND.n9219 GND.n9218 0.152939
R25028 GND.n9219 GND.n757 0.152939
R25029 GND.n9227 GND.n757 0.152939
R25030 GND.n9228 GND.n9227 0.152939
R25031 GND.n9229 GND.n9228 0.152939
R25032 GND.n9229 GND.n751 0.152939
R25033 GND.n9237 GND.n751 0.152939
R25034 GND.n9238 GND.n9237 0.152939
R25035 GND.n9239 GND.n9238 0.152939
R25036 GND.n9239 GND.n745 0.152939
R25037 GND.n9247 GND.n745 0.152939
R25038 GND.n9248 GND.n9247 0.152939
R25039 GND.n9249 GND.n9248 0.152939
R25040 GND.n9249 GND.n739 0.152939
R25041 GND.n9257 GND.n739 0.152939
R25042 GND.n9258 GND.n9257 0.152939
R25043 GND.n9259 GND.n9258 0.152939
R25044 GND.n9259 GND.n733 0.152939
R25045 GND.n9267 GND.n733 0.152939
R25046 GND.n9268 GND.n9267 0.152939
R25047 GND.n9269 GND.n9268 0.152939
R25048 GND.n9269 GND.n727 0.152939
R25049 GND.n9277 GND.n727 0.152939
R25050 GND.n9278 GND.n9277 0.152939
R25051 GND.n9279 GND.n9278 0.152939
R25052 GND.n9279 GND.n721 0.152939
R25053 GND.n9287 GND.n721 0.152939
R25054 GND.n9288 GND.n9287 0.152939
R25055 GND.n9289 GND.n9288 0.152939
R25056 GND.n9289 GND.n715 0.152939
R25057 GND.n9297 GND.n715 0.152939
R25058 GND.n9298 GND.n9297 0.152939
R25059 GND.n9299 GND.n9298 0.152939
R25060 GND.n9299 GND.n709 0.152939
R25061 GND.n9307 GND.n709 0.152939
R25062 GND.n9308 GND.n9307 0.152939
R25063 GND.n9309 GND.n9308 0.152939
R25064 GND.n9309 GND.n703 0.152939
R25065 GND.n9317 GND.n703 0.152939
R25066 GND.n9318 GND.n9317 0.152939
R25067 GND.n9319 GND.n9318 0.152939
R25068 GND.n9327 GND.n697 0.152939
R25069 GND.n9328 GND.n9327 0.152939
R25070 GND.n9329 GND.n9328 0.152939
R25071 GND.n9329 GND.n691 0.152939
R25072 GND.n9337 GND.n691 0.152939
R25073 GND.n9338 GND.n9337 0.152939
R25074 GND.n9339 GND.n9338 0.152939
R25075 GND.n9339 GND.n685 0.152939
R25076 GND.n9347 GND.n685 0.152939
R25077 GND.n9348 GND.n9347 0.152939
R25078 GND.n9349 GND.n9348 0.152939
R25079 GND.n9349 GND.n679 0.152939
R25080 GND.n9357 GND.n679 0.152939
R25081 GND.n9358 GND.n9357 0.152939
R25082 GND.n9359 GND.n9358 0.152939
R25083 GND.n9359 GND.n673 0.152939
R25084 GND.n9367 GND.n673 0.152939
R25085 GND.n9368 GND.n9367 0.152939
R25086 GND.n9369 GND.n9368 0.152939
R25087 GND.n9369 GND.n667 0.152939
R25088 GND.n9377 GND.n667 0.152939
R25089 GND.n9378 GND.n9377 0.152939
R25090 GND.n9379 GND.n9378 0.152939
R25091 GND.n9379 GND.n661 0.152939
R25092 GND.n9387 GND.n661 0.152939
R25093 GND.n9388 GND.n9387 0.152939
R25094 GND.n9389 GND.n9388 0.152939
R25095 GND.n9389 GND.n655 0.152939
R25096 GND.n9397 GND.n655 0.152939
R25097 GND.n9398 GND.n9397 0.152939
R25098 GND.n9399 GND.n9398 0.152939
R25099 GND.n9399 GND.n649 0.152939
R25100 GND.n9407 GND.n649 0.152939
R25101 GND.n9408 GND.n9407 0.152939
R25102 GND.n9409 GND.n9408 0.152939
R25103 GND.n9409 GND.n643 0.152939
R25104 GND.n9417 GND.n643 0.152939
R25105 GND.n9418 GND.n9417 0.152939
R25106 GND.n9419 GND.n9418 0.152939
R25107 GND.n9419 GND.n637 0.152939
R25108 GND.n9427 GND.n637 0.152939
R25109 GND.n9428 GND.n9427 0.152939
R25110 GND.n9429 GND.n9428 0.152939
R25111 GND.n9429 GND.n631 0.152939
R25112 GND.n9437 GND.n631 0.152939
R25113 GND.n9438 GND.n9437 0.152939
R25114 GND.n9439 GND.n9438 0.152939
R25115 GND.n9439 GND.n625 0.152939
R25116 GND.n9447 GND.n625 0.152939
R25117 GND.n9448 GND.n9447 0.152939
R25118 GND.n9450 GND.n9448 0.152939
R25119 GND.n9450 GND.n9449 0.152939
R25120 GND.n9449 GND.n619 0.152939
R25121 GND.n9459 GND.n619 0.152939
R25122 GND.n6882 GND.n6881 0.152939
R25123 GND.n6883 GND.n6882 0.152939
R25124 GND.n6883 GND.n3717 0.152939
R25125 GND.n6906 GND.n3717 0.152939
R25126 GND.n6907 GND.n6906 0.152939
R25127 GND.n6908 GND.n6907 0.152939
R25128 GND.n6909 GND.n6908 0.152939
R25129 GND.n6909 GND.n3695 0.152939
R25130 GND.n6933 GND.n3695 0.152939
R25131 GND.n6934 GND.n6933 0.152939
R25132 GND.n6935 GND.n6934 0.152939
R25133 GND.n6936 GND.n6935 0.152939
R25134 GND.n6936 GND.n3675 0.152939
R25135 GND.n6962 GND.n3675 0.152939
R25136 GND.n6963 GND.n6962 0.152939
R25137 GND.n6964 GND.n6963 0.152939
R25138 GND.n6965 GND.n6964 0.152939
R25139 GND.n6965 GND.n3653 0.152939
R25140 GND.n6989 GND.n3653 0.152939
R25141 GND.n6990 GND.n6989 0.152939
R25142 GND.n6991 GND.n6990 0.152939
R25143 GND.n6992 GND.n6991 0.152939
R25144 GND.n6992 GND.n3631 0.152939
R25145 GND.n7015 GND.n3631 0.152939
R25146 GND.n7016 GND.n7015 0.152939
R25147 GND.n7017 GND.n7016 0.152939
R25148 GND.n7018 GND.n7017 0.152939
R25149 GND.n7018 GND.n3609 0.152939
R25150 GND.n7042 GND.n3609 0.152939
R25151 GND.n7043 GND.n7042 0.152939
R25152 GND.n7044 GND.n7043 0.152939
R25153 GND.n7045 GND.n7044 0.152939
R25154 GND.n7045 GND.n3588 0.152939
R25155 GND.n7070 GND.n3588 0.152939
R25156 GND.n7071 GND.n7070 0.152939
R25157 GND.n7072 GND.n7071 0.152939
R25158 GND.n7073 GND.n7072 0.152939
R25159 GND.n7074 GND.n7073 0.152939
R25160 GND.n7076 GND.n7074 0.152939
R25161 GND.n7076 GND.n7075 0.152939
R25162 GND.n7075 GND.n583 0.152939
R25163 GND.n584 GND.n583 0.152939
R25164 GND.n585 GND.n584 0.152939
R25165 GND.n588 GND.n585 0.152939
R25166 GND.n589 GND.n588 0.152939
R25167 GND.n590 GND.n589 0.152939
R25168 GND.n591 GND.n590 0.152939
R25169 GND.n594 GND.n591 0.152939
R25170 GND.n595 GND.n594 0.152939
R25171 GND.n596 GND.n595 0.152939
R25172 GND.n597 GND.n596 0.152939
R25173 GND.n602 GND.n597 0.152939
R25174 GND.n603 GND.n602 0.152939
R25175 GND.n604 GND.n603 0.152939
R25176 GND.n605 GND.n604 0.152939
R25177 GND.n610 GND.n605 0.152939
R25178 GND.n611 GND.n610 0.152939
R25179 GND.n612 GND.n611 0.152939
R25180 GND.n613 GND.n612 0.152939
R25181 GND.n618 GND.n613 0.152939
R25182 GND.n9460 GND.n618 0.152939
R25183 GND.n6836 GND.n3727 0.152939
R25184 GND.n6895 GND.n3727 0.152939
R25185 GND.n6896 GND.n6895 0.152939
R25186 GND.n6897 GND.n6896 0.152939
R25187 GND.n6898 GND.n6897 0.152939
R25188 GND.n6898 GND.n3705 0.152939
R25189 GND.n6922 GND.n3705 0.152939
R25190 GND.n6923 GND.n6922 0.152939
R25191 GND.n6924 GND.n6923 0.152939
R25192 GND.n6925 GND.n6924 0.152939
R25193 GND.n6925 GND.n3684 0.152939
R25194 GND.n6951 GND.n3684 0.152939
R25195 GND.n6952 GND.n6951 0.152939
R25196 GND.n6953 GND.n6952 0.152939
R25197 GND.n6954 GND.n6953 0.152939
R25198 GND.n6954 GND.n3664 0.152939
R25199 GND.n6978 GND.n3664 0.152939
R25200 GND.n6979 GND.n6978 0.152939
R25201 GND.n6980 GND.n6979 0.152939
R25202 GND.n6981 GND.n6980 0.152939
R25203 GND.n6981 GND.n3641 0.152939
R25204 GND.n7004 GND.n3641 0.152939
R25205 GND.n7005 GND.n7004 0.152939
R25206 GND.n7006 GND.n7005 0.152939
R25207 GND.n7007 GND.n7006 0.152939
R25208 GND.n7007 GND.n3619 0.152939
R25209 GND.n7031 GND.n3619 0.152939
R25210 GND.n7032 GND.n7031 0.152939
R25211 GND.n7033 GND.n7032 0.152939
R25212 GND.n7034 GND.n7033 0.152939
R25213 GND.n7034 GND.n3598 0.152939
R25214 GND.n7059 GND.n3598 0.152939
R25215 GND.n7060 GND.n7059 0.152939
R25216 GND.n7061 GND.n7060 0.152939
R25217 GND.n7062 GND.n7061 0.152939
R25218 GND.n7062 GND.n3575 0.152939
R25219 GND.n7092 GND.n3575 0.152939
R25220 GND.n7093 GND.n7092 0.152939
R25221 GND.n7094 GND.n7093 0.152939
R25222 GND.n7095 GND.n7094 0.152939
R25223 GND.n7095 GND.n564 0.152939
R25224 GND.n9509 GND.n564 0.152939
R25225 GND.n9510 GND.n9509 0.152939
R25226 GND.n9511 GND.n9510 0.152939
R25227 GND.n9512 GND.n9511 0.152939
R25228 GND.n9512 GND.n483 0.152939
R25229 GND.n9609 GND.n483 0.152939
R25230 GND.n6268 GND.n6267 0.152939
R25231 GND.n6269 GND.n6268 0.152939
R25232 GND.n6269 GND.n6264 0.152939
R25233 GND.n6277 GND.n6264 0.152939
R25234 GND.n6278 GND.n6277 0.152939
R25235 GND.n6279 GND.n6278 0.152939
R25236 GND.n6279 GND.n6262 0.152939
R25237 GND.n6287 GND.n6262 0.152939
R25238 GND.n6288 GND.n6287 0.152939
R25239 GND.n6297 GND.n6117 0.152939
R25240 GND.n6298 GND.n6297 0.152939
R25241 GND.n6299 GND.n6298 0.152939
R25242 GND.n6299 GND.n6115 0.152939
R25243 GND.n6307 GND.n6115 0.152939
R25244 GND.n6308 GND.n6307 0.152939
R25245 GND.n6309 GND.n6308 0.152939
R25246 GND.n6309 GND.n6113 0.152939
R25247 GND.n6317 GND.n6113 0.152939
R25248 GND.n6318 GND.n6317 0.152939
R25249 GND.n6319 GND.n6318 0.152939
R25250 GND.n6319 GND.n6106 0.152939
R25251 GND.n6323 GND.n6106 0.152939
R25252 GND.n3362 GND.n3361 0.152939
R25253 GND.n3363 GND.n3362 0.152939
R25254 GND.n6587 GND.n3363 0.152939
R25255 GND.n6588 GND.n6587 0.152939
R25256 GND.n6589 GND.n6588 0.152939
R25257 GND.n6590 GND.n6589 0.152939
R25258 GND.n6590 GND.n3944 0.152939
R25259 GND.n6612 GND.n3944 0.152939
R25260 GND.n6613 GND.n6612 0.152939
R25261 GND.n6614 GND.n6613 0.152939
R25262 GND.n6615 GND.n6614 0.152939
R25263 GND.n6615 GND.n3921 0.152939
R25264 GND.n6636 GND.n3921 0.152939
R25265 GND.n6637 GND.n6636 0.152939
R25266 GND.n6638 GND.n6637 0.152939
R25267 GND.n6639 GND.n6638 0.152939
R25268 GND.n6639 GND.n3898 0.152939
R25269 GND.n6661 GND.n3898 0.152939
R25270 GND.n6662 GND.n6661 0.152939
R25271 GND.n6663 GND.n6662 0.152939
R25272 GND.n6664 GND.n6663 0.152939
R25273 GND.n6664 GND.n3876 0.152939
R25274 GND.n6686 GND.n3876 0.152939
R25275 GND.n6687 GND.n6686 0.152939
R25276 GND.n6688 GND.n6687 0.152939
R25277 GND.n6689 GND.n6688 0.152939
R25278 GND.n6689 GND.n3853 0.152939
R25279 GND.n6711 GND.n3853 0.152939
R25280 GND.n6712 GND.n6711 0.152939
R25281 GND.n6713 GND.n6712 0.152939
R25282 GND.n6714 GND.n6713 0.152939
R25283 GND.n6714 GND.n3830 0.152939
R25284 GND.n6735 GND.n3830 0.152939
R25285 GND.n6736 GND.n6735 0.152939
R25286 GND.n6737 GND.n6736 0.152939
R25287 GND.n6738 GND.n6737 0.152939
R25288 GND.n6738 GND.n3807 0.152939
R25289 GND.n6760 GND.n3807 0.152939
R25290 GND.n6761 GND.n6760 0.152939
R25291 GND.n6762 GND.n6761 0.152939
R25292 GND.n6763 GND.n6762 0.152939
R25293 GND.n6763 GND.n3785 0.152939
R25294 GND.n6785 GND.n3785 0.152939
R25295 GND.n6786 GND.n6785 0.152939
R25296 GND.n6787 GND.n6786 0.152939
R25297 GND.n6789 GND.n6787 0.152939
R25298 GND.n6789 GND.n6788 0.152939
R25299 GND.n2153 GND.n2107 0.152939
R25300 GND.n2154 GND.n2153 0.152939
R25301 GND.n2157 GND.n2154 0.152939
R25302 GND.n2158 GND.n2157 0.152939
R25303 GND.n2159 GND.n2158 0.152939
R25304 GND.n2160 GND.n2159 0.152939
R25305 GND.n2163 GND.n2160 0.152939
R25306 GND.n2164 GND.n2163 0.152939
R25307 GND.n2165 GND.n2164 0.152939
R25308 GND.n2166 GND.n2165 0.152939
R25309 GND.n2166 GND.n2043 0.152939
R25310 GND.n2893 GND.n2043 0.152939
R25311 GND.n2894 GND.n2893 0.152939
R25312 GND.n2895 GND.n2894 0.152939
R25313 GND.n2896 GND.n2895 0.152939
R25314 GND.n2897 GND.n2896 0.152939
R25315 GND.n2900 GND.n2897 0.152939
R25316 GND.n2901 GND.n2900 0.152939
R25317 GND.n2902 GND.n2901 0.152939
R25318 GND.n2903 GND.n2902 0.152939
R25319 GND.n2906 GND.n2903 0.152939
R25320 GND.n2907 GND.n2906 0.152939
R25321 GND.n2908 GND.n2907 0.152939
R25322 GND.n2909 GND.n2908 0.152939
R25323 GND.n2912 GND.n2909 0.152939
R25324 GND.n2913 GND.n2912 0.152939
R25325 GND.n2914 GND.n2913 0.152939
R25326 GND.n2915 GND.n2914 0.152939
R25327 GND.n2918 GND.n2915 0.152939
R25328 GND.n2919 GND.n2918 0.152939
R25329 GND.n2920 GND.n2919 0.152939
R25330 GND.n2921 GND.n2920 0.152939
R25331 GND.n2924 GND.n2921 0.152939
R25332 GND.n2925 GND.n2924 0.152939
R25333 GND.n2926 GND.n2925 0.152939
R25334 GND.n2927 GND.n2926 0.152939
R25335 GND.n2930 GND.n2927 0.152939
R25336 GND.n2931 GND.n2930 0.152939
R25337 GND.n2932 GND.n2931 0.152939
R25338 GND.n2933 GND.n2932 0.152939
R25339 GND.n2936 GND.n2933 0.152939
R25340 GND.n2937 GND.n2936 0.152939
R25341 GND.n2938 GND.n2937 0.152939
R25342 GND.n2939 GND.n2938 0.152939
R25343 GND.n2942 GND.n2939 0.152939
R25344 GND.n2943 GND.n2942 0.152939
R25345 GND.n2944 GND.n2943 0.152939
R25346 GND.n2945 GND.n2944 0.152939
R25347 GND.n2948 GND.n2945 0.152939
R25348 GND.n2949 GND.n2948 0.152939
R25349 GND.n2950 GND.n2949 0.152939
R25350 GND.n2951 GND.n2950 0.152939
R25351 GND.n2957 GND.n2951 0.152939
R25352 GND.n2958 GND.n2957 0.152939
R25353 GND.n2959 GND.n2958 0.152939
R25354 GND.n2960 GND.n2959 0.152939
R25355 GND.n2975 GND.n2960 0.152939
R25356 GND.n2976 GND.n2975 0.152939
R25357 GND.n2977 GND.n2976 0.152939
R25358 GND.n2978 GND.n2977 0.152939
R25359 GND.n2994 GND.n2978 0.152939
R25360 GND.n2995 GND.n2994 0.152939
R25361 GND.n2996 GND.n2995 0.152939
R25362 GND.n2997 GND.n2996 0.152939
R25363 GND.n3015 GND.n2997 0.152939
R25364 GND.n3016 GND.n3015 0.152939
R25365 GND.n3017 GND.n3016 0.152939
R25366 GND.n3018 GND.n3017 0.152939
R25367 GND.n4893 GND.n3018 0.152939
R25368 GND.n4894 GND.n4893 0.152939
R25369 GND.n4895 GND.n4894 0.152939
R25370 GND.n4896 GND.n4895 0.152939
R25371 GND.n4897 GND.n4896 0.152939
R25372 GND.n4898 GND.n4897 0.152939
R25373 GND.n4898 GND.n4624 0.152939
R25374 GND.n4939 GND.n4624 0.152939
R25375 GND.n4940 GND.n4939 0.152939
R25376 GND.n4941 GND.n4940 0.152939
R25377 GND.n4942 GND.n4941 0.152939
R25378 GND.n4942 GND.n4595 0.152939
R25379 GND.n4993 GND.n4595 0.152939
R25380 GND.n4994 GND.n4993 0.152939
R25381 GND.n4995 GND.n4994 0.152939
R25382 GND.n4996 GND.n4995 0.152939
R25383 GND.n4996 GND.n4572 0.152939
R25384 GND.n5053 GND.n4572 0.152939
R25385 GND.n5054 GND.n5053 0.152939
R25386 GND.n5055 GND.n5054 0.152939
R25387 GND.n5056 GND.n5055 0.152939
R25388 GND.n5057 GND.n5056 0.152939
R25389 GND.n5059 GND.n5057 0.152939
R25390 GND.n5060 GND.n5059 0.152939
R25391 GND.n5060 GND.n4533 0.152939
R25392 GND.n5111 GND.n4533 0.152939
R25393 GND.n5112 GND.n5111 0.152939
R25394 GND.n5113 GND.n5112 0.152939
R25395 GND.n5113 GND.n4507 0.152939
R25396 GND.n5156 GND.n4507 0.152939
R25397 GND.n5157 GND.n5156 0.152939
R25398 GND.n5158 GND.n5157 0.152939
R25399 GND.n5159 GND.n5158 0.152939
R25400 GND.n5159 GND.n4487 0.152939
R25401 GND.n5216 GND.n4487 0.152939
R25402 GND.n5217 GND.n5216 0.152939
R25403 GND.n5218 GND.n5217 0.152939
R25404 GND.n5219 GND.n5218 0.152939
R25405 GND.n5220 GND.n5219 0.152939
R25406 GND.n5221 GND.n5220 0.152939
R25407 GND.n5221 GND.n4452 0.152939
R25408 GND.n5262 GND.n4452 0.152939
R25409 GND.n5263 GND.n5262 0.152939
R25410 GND.n5264 GND.n5263 0.152939
R25411 GND.n5265 GND.n5264 0.152939
R25412 GND.n5265 GND.n4424 0.152939
R25413 GND.n5317 GND.n4424 0.152939
R25414 GND.n5318 GND.n5317 0.152939
R25415 GND.n5319 GND.n5318 0.152939
R25416 GND.n5320 GND.n5319 0.152939
R25417 GND.n5320 GND.n4401 0.152939
R25418 GND.n5378 GND.n4401 0.152939
R25419 GND.n5379 GND.n5378 0.152939
R25420 GND.n5380 GND.n5379 0.152939
R25421 GND.n5381 GND.n5380 0.152939
R25422 GND.n5382 GND.n5381 0.152939
R25423 GND.n5383 GND.n5382 0.152939
R25424 GND.n5383 GND.n4366 0.152939
R25425 GND.n5424 GND.n4366 0.152939
R25426 GND.n5425 GND.n5424 0.152939
R25427 GND.n5426 GND.n5425 0.152939
R25428 GND.n5427 GND.n5426 0.152939
R25429 GND.n5427 GND.n4337 0.152939
R25430 GND.n5477 GND.n4337 0.152939
R25431 GND.n5478 GND.n5477 0.152939
R25432 GND.n5479 GND.n5478 0.152939
R25433 GND.n5480 GND.n5479 0.152939
R25434 GND.n5480 GND.n4314 0.152939
R25435 GND.n5549 GND.n4314 0.152939
R25436 GND.n5550 GND.n5549 0.152939
R25437 GND.n5551 GND.n5550 0.152939
R25438 GND.n5552 GND.n5551 0.152939
R25439 GND.n5553 GND.n5552 0.152939
R25440 GND.n5554 GND.n5553 0.152939
R25441 GND.n5554 GND.n4281 0.152939
R25442 GND.n5595 GND.n4281 0.152939
R25443 GND.n5596 GND.n5595 0.152939
R25444 GND.n5597 GND.n5596 0.152939
R25445 GND.n5598 GND.n5597 0.152939
R25446 GND.n5598 GND.n4253 0.152939
R25447 GND.n5633 GND.n4253 0.152939
R25448 GND.n5634 GND.n5633 0.152939
R25449 GND.n5635 GND.n5634 0.152939
R25450 GND.n5635 GND.n4229 0.152939
R25451 GND.n5689 GND.n4229 0.152939
R25452 GND.n5690 GND.n5689 0.152939
R25453 GND.n5691 GND.n5690 0.152939
R25454 GND.n5692 GND.n5691 0.152939
R25455 GND.n5692 GND.n4206 0.152939
R25456 GND.n5723 GND.n4206 0.152939
R25457 GND.n5724 GND.n5723 0.152939
R25458 GND.n5725 GND.n5724 0.152939
R25459 GND.n5726 GND.n5725 0.152939
R25460 GND.n5726 GND.n4183 0.152939
R25461 GND.n5804 GND.n4183 0.152939
R25462 GND.n5805 GND.n5804 0.152939
R25463 GND.n5806 GND.n5805 0.152939
R25464 GND.n5807 GND.n5806 0.152939
R25465 GND.n5808 GND.n5807 0.152939
R25466 GND.n5810 GND.n5808 0.152939
R25467 GND.n5811 GND.n5810 0.152939
R25468 GND.n5811 GND.n4146 0.152939
R25469 GND.n5864 GND.n4146 0.152939
R25470 GND.n5865 GND.n5864 0.152939
R25471 GND.n5866 GND.n5865 0.152939
R25472 GND.n5867 GND.n5866 0.152939
R25473 GND.n5868 GND.n5867 0.152939
R25474 GND.n5869 GND.n5868 0.152939
R25475 GND.n5869 GND.n4111 0.152939
R25476 GND.n5910 GND.n4111 0.152939
R25477 GND.n5911 GND.n5910 0.152939
R25478 GND.n5912 GND.n5911 0.152939
R25479 GND.n5913 GND.n5912 0.152939
R25480 GND.n5913 GND.n4082 0.152939
R25481 GND.n5963 GND.n4082 0.152939
R25482 GND.n5964 GND.n5963 0.152939
R25483 GND.n5965 GND.n5964 0.152939
R25484 GND.n5966 GND.n5965 0.152939
R25485 GND.n5966 GND.n4058 0.152939
R25486 GND.n6012 GND.n4058 0.152939
R25487 GND.n6013 GND.n6012 0.152939
R25488 GND.n6014 GND.n6013 0.152939
R25489 GND.n6015 GND.n6014 0.152939
R25490 GND.n6016 GND.n6015 0.152939
R25491 GND.n6018 GND.n6016 0.152939
R25492 GND.n6019 GND.n6018 0.152939
R25493 GND.n6019 GND.n4017 0.152939
R25494 GND.n6088 GND.n4017 0.152939
R25495 GND.n6089 GND.n6088 0.152939
R25496 GND.n6090 GND.n6089 0.152939
R25497 GND.n6091 GND.n6090 0.152939
R25498 GND.n6091 GND.n3995 0.152939
R25499 GND.n6353 GND.n3995 0.152939
R25500 GND.n6354 GND.n6353 0.152939
R25501 GND.n6355 GND.n6354 0.152939
R25502 GND.n6357 GND.n6355 0.152939
R25503 GND.n6357 GND.n6356 0.152939
R25504 GND.n6356 GND.n3236 0.152939
R25505 GND.n3237 GND.n3236 0.152939
R25506 GND.n3238 GND.n3237 0.152939
R25507 GND.n3252 GND.n3238 0.152939
R25508 GND.n3253 GND.n3252 0.152939
R25509 GND.n3254 GND.n3253 0.152939
R25510 GND.n3255 GND.n3254 0.152939
R25511 GND.n3277 GND.n3255 0.152939
R25512 GND.n3278 GND.n3277 0.152939
R25513 GND.n3279 GND.n3278 0.152939
R25514 GND.n3280 GND.n3279 0.152939
R25515 GND.n3281 GND.n3280 0.152939
R25516 GND.n3286 GND.n3281 0.152939
R25517 GND.n3287 GND.n3286 0.152939
R25518 GND.n3288 GND.n3287 0.152939
R25519 GND.n3289 GND.n3288 0.152939
R25520 GND.n6443 GND.n3289 0.152939
R25521 GND.n6444 GND.n6443 0.152939
R25522 GND.n6444 GND.n6441 0.152939
R25523 GND.n6450 GND.n6441 0.152939
R25524 GND.n6451 GND.n6450 0.152939
R25525 GND.n6452 GND.n6451 0.152939
R25526 GND.n6453 GND.n6452 0.152939
R25527 GND.n6454 GND.n6453 0.152939
R25528 GND.n6457 GND.n6454 0.152939
R25529 GND.n6458 GND.n6457 0.152939
R25530 GND.n6459 GND.n6458 0.152939
R25531 GND.n6460 GND.n6459 0.152939
R25532 GND.n6463 GND.n6460 0.152939
R25533 GND.n6464 GND.n6463 0.152939
R25534 GND.n6465 GND.n6464 0.152939
R25535 GND.n6466 GND.n6465 0.152939
R25536 GND.n6469 GND.n6466 0.152939
R25537 GND.n6470 GND.n6469 0.152939
R25538 GND.n6471 GND.n6470 0.152939
R25539 GND.n6472 GND.n6471 0.152939
R25540 GND.n6475 GND.n6472 0.152939
R25541 GND.n6476 GND.n6475 0.152939
R25542 GND.n6477 GND.n6476 0.152939
R25543 GND.n6478 GND.n6477 0.152939
R25544 GND.n6481 GND.n6478 0.152939
R25545 GND.n6482 GND.n6481 0.152939
R25546 GND.n6483 GND.n6482 0.152939
R25547 GND.n6484 GND.n6483 0.152939
R25548 GND.n6487 GND.n6484 0.152939
R25549 GND.n6488 GND.n6487 0.152939
R25550 GND.n6489 GND.n6488 0.152939
R25551 GND.n6490 GND.n6489 0.152939
R25552 GND.n6493 GND.n6490 0.152939
R25553 GND.n6494 GND.n6493 0.152939
R25554 GND.n6495 GND.n6494 0.152939
R25555 GND.n6496 GND.n6495 0.152939
R25556 GND.n6499 GND.n6496 0.152939
R25557 GND.n6500 GND.n6499 0.152939
R25558 GND.n6501 GND.n6500 0.152939
R25559 GND.n6502 GND.n6501 0.152939
R25560 GND.n6505 GND.n6502 0.152939
R25561 GND.n6506 GND.n6505 0.152939
R25562 GND.n6507 GND.n6506 0.152939
R25563 GND.n6508 GND.n6507 0.152939
R25564 GND.n6511 GND.n6508 0.152939
R25565 GND.n6512 GND.n6511 0.152939
R25566 GND.n6513 GND.n6512 0.152939
R25567 GND.n6514 GND.n6513 0.152939
R25568 GND.n6514 GND.n3745 0.152939
R25569 GND.n6881 GND.n3745 0.152939
R25570 GND.n2826 GND.n2825 0.152939
R25571 GND.n2826 GND.n2083 0.152939
R25572 GND.n2848 GND.n2083 0.152939
R25573 GND.n2849 GND.n2848 0.152939
R25574 GND.n2850 GND.n2849 0.152939
R25575 GND.n2851 GND.n2850 0.152939
R25576 GND.n2851 GND.n2061 0.152939
R25577 GND.n2873 GND.n2061 0.152939
R25578 GND.n2874 GND.n2873 0.152939
R25579 GND.n2875 GND.n2874 0.152939
R25580 GND.n2876 GND.n2875 0.152939
R25581 GND.n2876 GND.n2033 0.152939
R25582 GND.n7671 GND.n2033 0.152939
R25583 GND.n7672 GND.n7671 0.152939
R25584 GND.n7673 GND.n7672 0.152939
R25585 GND.n7674 GND.n7673 0.152939
R25586 GND.n7674 GND.n2010 0.152939
R25587 GND.n7695 GND.n2010 0.152939
R25588 GND.n7696 GND.n7695 0.152939
R25589 GND.n7697 GND.n7696 0.152939
R25590 GND.n7698 GND.n7697 0.152939
R25591 GND.n7698 GND.n1987 0.152939
R25592 GND.n7720 GND.n1987 0.152939
R25593 GND.n7721 GND.n7720 0.152939
R25594 GND.n7722 GND.n7721 0.152939
R25595 GND.n7723 GND.n7722 0.152939
R25596 GND.n7723 GND.n1965 0.152939
R25597 GND.n7745 GND.n1965 0.152939
R25598 GND.n7746 GND.n7745 0.152939
R25599 GND.n7747 GND.n7746 0.152939
R25600 GND.n7748 GND.n7747 0.152939
R25601 GND.n7748 GND.n1942 0.152939
R25602 GND.n7770 GND.n1942 0.152939
R25603 GND.n7771 GND.n7770 0.152939
R25604 GND.n7772 GND.n7771 0.152939
R25605 GND.n7773 GND.n7772 0.152939
R25606 GND.n7773 GND.n1919 0.152939
R25607 GND.n7794 GND.n1919 0.152939
R25608 GND.n7795 GND.n7794 0.152939
R25609 GND.n7796 GND.n7795 0.152939
R25610 GND.n7797 GND.n7796 0.152939
R25611 GND.n7797 GND.n1897 0.152939
R25612 GND.n7821 GND.n1897 0.152939
R25613 GND.n7822 GND.n7821 0.152939
R25614 GND.n7823 GND.n7822 0.152939
R25615 GND.n7823 GND.n1778 0.152939
R25616 GND.n7921 GND.n1778 0.152939
R25617 GND.n1476 GND.n1475 0.152939
R25618 GND.n1477 GND.n1476 0.152939
R25619 GND.n1478 GND.n1477 0.152939
R25620 GND.n1479 GND.n1478 0.152939
R25621 GND.n1480 GND.n1479 0.152939
R25622 GND.n1481 GND.n1480 0.152939
R25623 GND.n1482 GND.n1481 0.152939
R25624 GND.n1483 GND.n1482 0.152939
R25625 GND.n1484 GND.n1483 0.152939
R25626 GND.n1485 GND.n1484 0.152939
R25627 GND.n1486 GND.n1485 0.152939
R25628 GND.n1489 GND.n1486 0.152939
R25629 GND.n1490 GND.n1489 0.152939
R25630 GND.n1491 GND.n1490 0.152939
R25631 GND.n1492 GND.n1491 0.152939
R25632 GND.n1493 GND.n1492 0.152939
R25633 GND.n1494 GND.n1493 0.152939
R25634 GND.n1495 GND.n1494 0.152939
R25635 GND.n1496 GND.n1495 0.152939
R25636 GND.n1497 GND.n1496 0.152939
R25637 GND.n1498 GND.n1497 0.152939
R25638 GND.n1499 GND.n1498 0.152939
R25639 GND.n8103 GND.n1499 0.152939
R25640 GND.n8103 GND.n8102 0.152939
R25641 GND.n8102 GND.n8101 0.152939
R25642 GND.n1539 GND.n1535 0.152939
R25643 GND.n1540 GND.n1539 0.152939
R25644 GND.n1541 GND.n1540 0.152939
R25645 GND.n1542 GND.n1541 0.152939
R25646 GND.n1543 GND.n1542 0.152939
R25647 GND.n2508 GND.n1543 0.152939
R25648 GND.n2509 GND.n2508 0.152939
R25649 GND.n2510 GND.n2509 0.152939
R25650 GND.n2510 GND.n2357 0.152939
R25651 GND.n2532 GND.n2357 0.152939
R25652 GND.n2533 GND.n2532 0.152939
R25653 GND.n2534 GND.n2533 0.152939
R25654 GND.n2535 GND.n2534 0.152939
R25655 GND.n2535 GND.n2334 0.152939
R25656 GND.n2557 GND.n2334 0.152939
R25657 GND.n2558 GND.n2557 0.152939
R25658 GND.n2559 GND.n2558 0.152939
R25659 GND.n2560 GND.n2559 0.152939
R25660 GND.n2560 GND.n2311 0.152939
R25661 GND.n2581 GND.n2311 0.152939
R25662 GND.n2582 GND.n2581 0.152939
R25663 GND.n2583 GND.n2582 0.152939
R25664 GND.n2584 GND.n2583 0.152939
R25665 GND.n2584 GND.n2288 0.152939
R25666 GND.n2606 GND.n2288 0.152939
R25667 GND.n2607 GND.n2606 0.152939
R25668 GND.n2608 GND.n2607 0.152939
R25669 GND.n2609 GND.n2608 0.152939
R25670 GND.n2609 GND.n2266 0.152939
R25671 GND.n2639 GND.n2266 0.152939
R25672 GND.n2640 GND.n2639 0.152939
R25673 GND.n2641 GND.n2640 0.152939
R25674 GND.n2641 GND.n2247 0.152939
R25675 GND.n2706 GND.n2247 0.152939
R25676 GND.n2707 GND.n2706 0.152939
R25677 GND.n2708 GND.n2707 0.152939
R25678 GND.n2709 GND.n2708 0.152939
R25679 GND.n2709 GND.n2224 0.152939
R25680 GND.n2731 GND.n2224 0.152939
R25681 GND.n2732 GND.n2731 0.152939
R25682 GND.n2733 GND.n2732 0.152939
R25683 GND.n2734 GND.n2733 0.152939
R25684 GND.n2734 GND.n2201 0.152939
R25685 GND.n2755 GND.n2201 0.152939
R25686 GND.n2756 GND.n2755 0.152939
R25687 GND.n2757 GND.n2756 0.152939
R25688 GND.n2757 GND.n2106 0.152939
R25689 GND.n8174 GND.n1430 0.152939
R25690 GND.n1432 GND.n1430 0.152939
R25691 GND.n1438 GND.n1432 0.152939
R25692 GND.n1439 GND.n1438 0.152939
R25693 GND.n1440 GND.n1439 0.152939
R25694 GND.n1441 GND.n1440 0.152939
R25695 GND.n1446 GND.n1441 0.152939
R25696 GND.n1447 GND.n1446 0.152939
R25697 GND.n1448 GND.n1447 0.152939
R25698 GND.n1449 GND.n1448 0.152939
R25699 GND.n1516 GND.n1449 0.152939
R25700 GND.n1519 GND.n1516 0.152939
R25701 GND.n1520 GND.n1519 0.152939
R25702 GND.n1521 GND.n1520 0.152939
R25703 GND.n1522 GND.n1521 0.152939
R25704 GND.n1523 GND.n1522 0.152939
R25705 GND.n2427 GND.n1523 0.152939
R25706 GND.n2428 GND.n2427 0.152939
R25707 GND.n2433 GND.n2428 0.152939
R25708 GND.n2434 GND.n2433 0.152939
R25709 GND.n2435 GND.n2434 0.152939
R25710 GND.n2436 GND.n2435 0.152939
R25711 GND.n2437 GND.n2436 0.152939
R25712 GND.n2440 GND.n2437 0.152939
R25713 GND.n2441 GND.n2440 0.152939
R25714 GND.n2442 GND.n2441 0.152939
R25715 GND.n2443 GND.n2442 0.152939
R25716 GND.n2446 GND.n2443 0.152939
R25717 GND.n2447 GND.n2446 0.152939
R25718 GND.n2448 GND.n2447 0.152939
R25719 GND.n2449 GND.n2448 0.152939
R25720 GND.n2452 GND.n2449 0.152939
R25721 GND.n2453 GND.n2452 0.152939
R25722 GND.n2454 GND.n2453 0.152939
R25723 GND.n2455 GND.n2454 0.152939
R25724 GND.n2458 GND.n2455 0.152939
R25725 GND.n2459 GND.n2458 0.152939
R25726 GND.n2460 GND.n2459 0.152939
R25727 GND.n2461 GND.n2460 0.152939
R25728 GND.n2464 GND.n2461 0.152939
R25729 GND.n2465 GND.n2464 0.152939
R25730 GND.n2466 GND.n2465 0.152939
R25731 GND.n2467 GND.n2466 0.152939
R25732 GND.n2467 GND.n2258 0.152939
R25733 GND.n2648 GND.n2258 0.152939
R25734 GND.n2649 GND.n2648 0.152939
R25735 GND.n2650 GND.n2649 0.152939
R25736 GND.n2651 GND.n2650 0.152939
R25737 GND.n2652 GND.n2651 0.152939
R25738 GND.n2655 GND.n2652 0.152939
R25739 GND.n2656 GND.n2655 0.152939
R25740 GND.n2657 GND.n2656 0.152939
R25741 GND.n2658 GND.n2657 0.152939
R25742 GND.n2661 GND.n2658 0.152939
R25743 GND.n2662 GND.n2661 0.152939
R25744 GND.n2663 GND.n2662 0.152939
R25745 GND.n2664 GND.n2663 0.152939
R25746 GND.n2669 GND.n2664 0.152939
R25747 GND.n2670 GND.n2669 0.152939
R25748 GND.n2671 GND.n2670 0.152939
R25749 GND.n2671 GND.n2107 0.152939
R25750 GND.n8287 GND.n1321 0.152939
R25751 GND.n1326 GND.n1321 0.152939
R25752 GND.n1327 GND.n1326 0.152939
R25753 GND.n1328 GND.n1327 0.152939
R25754 GND.n1333 GND.n1328 0.152939
R25755 GND.n1334 GND.n1333 0.152939
R25756 GND.n1335 GND.n1334 0.152939
R25757 GND.n1336 GND.n1335 0.152939
R25758 GND.n1341 GND.n1336 0.152939
R25759 GND.n1342 GND.n1341 0.152939
R25760 GND.n1343 GND.n1342 0.152939
R25761 GND.n1344 GND.n1343 0.152939
R25762 GND.n1349 GND.n1344 0.152939
R25763 GND.n1350 GND.n1349 0.152939
R25764 GND.n1351 GND.n1350 0.152939
R25765 GND.n1352 GND.n1351 0.152939
R25766 GND.n1357 GND.n1352 0.152939
R25767 GND.n1358 GND.n1357 0.152939
R25768 GND.n1359 GND.n1358 0.152939
R25769 GND.n1360 GND.n1359 0.152939
R25770 GND.n1365 GND.n1360 0.152939
R25771 GND.n1366 GND.n1365 0.152939
R25772 GND.n1367 GND.n1366 0.152939
R25773 GND.n1368 GND.n1367 0.152939
R25774 GND.n1373 GND.n1368 0.152939
R25775 GND.n1374 GND.n1373 0.152939
R25776 GND.n1375 GND.n1374 0.152939
R25777 GND.n1376 GND.n1375 0.152939
R25778 GND.n1381 GND.n1376 0.152939
R25779 GND.n1382 GND.n1381 0.152939
R25780 GND.n1383 GND.n1382 0.152939
R25781 GND.n1384 GND.n1383 0.152939
R25782 GND.n1389 GND.n1384 0.152939
R25783 GND.n1390 GND.n1389 0.152939
R25784 GND.n1391 GND.n1390 0.152939
R25785 GND.n1392 GND.n1391 0.152939
R25786 GND.n1397 GND.n1392 0.152939
R25787 GND.n1398 GND.n1397 0.152939
R25788 GND.n1399 GND.n1398 0.152939
R25789 GND.n1400 GND.n1399 0.152939
R25790 GND.n1405 GND.n1400 0.152939
R25791 GND.n1406 GND.n1405 0.152939
R25792 GND.n1407 GND.n1406 0.152939
R25793 GND.n1408 GND.n1407 0.152939
R25794 GND.n1413 GND.n1408 0.152939
R25795 GND.n1414 GND.n1413 0.152939
R25796 GND.n1415 GND.n1414 0.152939
R25797 GND.n1416 GND.n1415 0.152939
R25798 GND.n1421 GND.n1416 0.152939
R25799 GND.n1422 GND.n1421 0.152939
R25800 GND.n1423 GND.n1422 0.152939
R25801 GND.n1424 GND.n1423 0.152939
R25802 GND.n1429 GND.n1424 0.152939
R25803 GND.n8175 GND.n1429 0.152939
R25804 GND.n6432 GND.n6430 0.152939
R25805 GND.n6433 GND.n6432 0.152939
R25806 GND.n6434 GND.n6433 0.152939
R25807 GND.n6434 GND.n3955 0.152939
R25808 GND.n6597 GND.n3955 0.152939
R25809 GND.n6598 GND.n6597 0.152939
R25810 GND.n6600 GND.n6598 0.152939
R25811 GND.n6600 GND.n6599 0.152939
R25812 GND.n6599 GND.n3934 0.152939
R25813 GND.n6622 GND.n3934 0.152939
R25814 GND.n6623 GND.n6622 0.152939
R25815 GND.n6625 GND.n6623 0.152939
R25816 GND.n6625 GND.n6624 0.152939
R25817 GND.n6624 GND.n3910 0.152939
R25818 GND.n6646 GND.n3910 0.152939
R25819 GND.n6647 GND.n6646 0.152939
R25820 GND.n6649 GND.n6647 0.152939
R25821 GND.n6649 GND.n6648 0.152939
R25822 GND.n6648 GND.n3887 0.152939
R25823 GND.n6671 GND.n3887 0.152939
R25824 GND.n6672 GND.n6671 0.152939
R25825 GND.n6674 GND.n6672 0.152939
R25826 GND.n6674 GND.n6673 0.152939
R25827 GND.n6673 GND.n3865 0.152939
R25828 GND.n6696 GND.n3865 0.152939
R25829 GND.n6697 GND.n6696 0.152939
R25830 GND.n6699 GND.n6697 0.152939
R25831 GND.n6699 GND.n6698 0.152939
R25832 GND.n6698 GND.n3843 0.152939
R25833 GND.n6721 GND.n3843 0.152939
R25834 GND.n6722 GND.n6721 0.152939
R25835 GND.n6724 GND.n6722 0.152939
R25836 GND.n6724 GND.n6723 0.152939
R25837 GND.n6723 GND.n3819 0.152939
R25838 GND.n6745 GND.n3819 0.152939
R25839 GND.n6746 GND.n6745 0.152939
R25840 GND.n6748 GND.n6746 0.152939
R25841 GND.n6748 GND.n6747 0.152939
R25842 GND.n6747 GND.n3796 0.152939
R25843 GND.n6770 GND.n3796 0.152939
R25844 GND.n6771 GND.n6770 0.152939
R25845 GND.n6773 GND.n6771 0.152939
R25846 GND.n6773 GND.n6772 0.152939
R25847 GND.n6772 GND.n3769 0.152939
R25848 GND.n6796 GND.n3769 0.152939
R25849 GND.n6797 GND.n6796 0.152939
R25850 GND.n6798 GND.n6797 0.152939
R25851 GND.n6798 GND.n3766 0.152939
R25852 GND.n6805 GND.n3766 0.152939
R25853 GND.n6806 GND.n6805 0.152939
R25854 GND.n6807 GND.n6806 0.152939
R25855 GND.n6807 GND.n406 0.152939
R25856 GND.n9693 GND.n407 0.152939
R25857 GND.n9689 GND.n407 0.152939
R25858 GND.n9689 GND.n9688 0.152939
R25859 GND.n9688 GND.n9687 0.152939
R25860 GND.n9687 GND.n413 0.152939
R25861 GND.n9683 GND.n413 0.152939
R25862 GND.n9683 GND.n9682 0.152939
R25863 GND.n9682 GND.n9681 0.152939
R25864 GND.n9681 GND.n418 0.152939
R25865 GND.n9677 GND.n418 0.152939
R25866 GND.n9677 GND.n9676 0.152939
R25867 GND.n9676 GND.n9675 0.152939
R25868 GND.n9675 GND.n423 0.152939
R25869 GND.n9671 GND.n423 0.152939
R25870 GND.n9671 GND.n9670 0.152939
R25871 GND.n9670 GND.n9669 0.152939
R25872 GND.n9669 GND.n428 0.152939
R25873 GND.n9665 GND.n428 0.152939
R25874 GND.n9665 GND.n9664 0.152939
R25875 GND.n9664 GND.n9663 0.152939
R25876 GND.n9663 GND.n433 0.152939
R25877 GND.n9659 GND.n433 0.152939
R25878 GND.n9659 GND.n9658 0.152939
R25879 GND.n9658 GND.n9657 0.152939
R25880 GND.n9657 GND.n438 0.152939
R25881 GND.n9653 GND.n438 0.152939
R25882 GND.n9653 GND.n9652 0.152939
R25883 GND.n9652 GND.n9651 0.152939
R25884 GND.n9651 GND.n443 0.152939
R25885 GND.n9647 GND.n443 0.152939
R25886 GND.n9647 GND.n9646 0.152939
R25887 GND.n9646 GND.n9645 0.152939
R25888 GND.n9645 GND.n448 0.152939
R25889 GND.n9641 GND.n448 0.152939
R25890 GND.n9641 GND.n9640 0.152939
R25891 GND.n9640 GND.n9639 0.152939
R25892 GND.n9639 GND.n453 0.152939
R25893 GND.n9635 GND.n453 0.152939
R25894 GND.n9635 GND.n9634 0.152939
R25895 GND.n9634 GND.n9633 0.152939
R25896 GND.n9633 GND.n458 0.152939
R25897 GND.n9629 GND.n458 0.152939
R25898 GND.n9629 GND.n9628 0.152939
R25899 GND.n9628 GND.n9627 0.152939
R25900 GND.n9627 GND.n463 0.152939
R25901 GND.n9623 GND.n463 0.152939
R25902 GND.n9623 GND.n9622 0.152939
R25903 GND.n9622 GND.n9621 0.152939
R25904 GND.n9621 GND.n468 0.152939
R25905 GND.n9617 GND.n468 0.152939
R25906 GND.n9617 GND.n9616 0.152939
R25907 GND.n9616 GND.n9615 0.152939
R25908 GND.n9564 GND.n9563 0.152939
R25909 GND.n9563 GND.n9562 0.152939
R25910 GND.n9562 GND.n9530 0.152939
R25911 GND.n9558 GND.n9530 0.152939
R25912 GND.n9558 GND.n9557 0.152939
R25913 GND.n9557 GND.n9556 0.152939
R25914 GND.n9556 GND.n9536 0.152939
R25915 GND.n9552 GND.n9536 0.152939
R25916 GND.n9552 GND.n9551 0.152939
R25917 GND.n9551 GND.n9550 0.152939
R25918 GND.n9550 GND.n9542 0.152939
R25919 GND.n9542 GND.n473 0.152939
R25920 GND.n9608 GND.n484 0.152939
R25921 GND.n9604 GND.n484 0.152939
R25922 GND.n9604 GND.n9603 0.152939
R25923 GND.n9603 GND.n9602 0.152939
R25924 GND.n9602 GND.n488 0.152939
R25925 GND.n9598 GND.n488 0.152939
R25926 GND.n9598 GND.n9597 0.152939
R25927 GND.n9597 GND.n9596 0.152939
R25928 GND.n9596 GND.n493 0.152939
R25929 GND.n9592 GND.n493 0.152939
R25930 GND.n9592 GND.n9591 0.152939
R25931 GND.n9591 GND.n9590 0.152939
R25932 GND.n9590 GND.n500 0.152939
R25933 GND.n9586 GND.n500 0.152939
R25934 GND.n9586 GND.n9585 0.152939
R25935 GND.n9585 GND.n9584 0.152939
R25936 GND.n9584 GND.n505 0.152939
R25937 GND.n9580 GND.n505 0.152939
R25938 GND.n9580 GND.n9579 0.152939
R25939 GND.n9579 GND.n9578 0.152939
R25940 GND.n9578 GND.n510 0.152939
R25941 GND.n9574 GND.n510 0.152939
R25942 GND.n9574 GND.n9573 0.152939
R25943 GND.n9573 GND.n9572 0.152939
R25944 GND.n9572 GND.n515 0.152939
R25945 GND.n6428 GND.n3963 0.152939
R25946 GND.n6424 GND.n3963 0.152939
R25947 GND.n6424 GND.n6423 0.152939
R25948 GND.n6423 GND.n3970 0.152939
R25949 GND.n6419 GND.n3970 0.152939
R25950 GND.n6419 GND.n3227 0.152939
R25951 GND.n3055 GND.n3051 0.152939
R25952 GND.n3056 GND.n3055 0.152939
R25953 GND.n7550 GND.n3056 0.152939
R25954 GND.n7550 GND.n7549 0.152939
R25955 GND.n7549 GND.n7548 0.152939
R25956 GND.n7548 GND.n3057 0.152939
R25957 GND.n7544 GND.n3057 0.152939
R25958 GND.n7544 GND.n7543 0.152939
R25959 GND.n7543 GND.n7542 0.152939
R25960 GND.n7542 GND.n3062 0.152939
R25961 GND.n7538 GND.n3062 0.152939
R25962 GND.n7538 GND.n7537 0.152939
R25963 GND.n7537 GND.n7536 0.152939
R25964 GND.n7536 GND.n3067 0.152939
R25965 GND.n7532 GND.n3067 0.152939
R25966 GND.n7532 GND.n7531 0.152939
R25967 GND.n7531 GND.n7530 0.152939
R25968 GND.n7530 GND.n3072 0.152939
R25969 GND.n7526 GND.n3072 0.152939
R25970 GND.n7526 GND.n7525 0.152939
R25971 GND.n7525 GND.n7524 0.152939
R25972 GND.n7524 GND.n3077 0.152939
R25973 GND.n7520 GND.n3077 0.152939
R25974 GND.n7520 GND.n7519 0.152939
R25975 GND.n7519 GND.n7518 0.152939
R25976 GND.n7518 GND.n3082 0.152939
R25977 GND.n7514 GND.n3082 0.152939
R25978 GND.n7514 GND.n7513 0.152939
R25979 GND.n7513 GND.n7512 0.152939
R25980 GND.n7512 GND.n3087 0.152939
R25981 GND.n7508 GND.n3087 0.152939
R25982 GND.n7508 GND.n7507 0.152939
R25983 GND.n7507 GND.n7506 0.152939
R25984 GND.n7506 GND.n3092 0.152939
R25985 GND.n7502 GND.n3092 0.152939
R25986 GND.n7502 GND.n7501 0.152939
R25987 GND.n7501 GND.n7500 0.152939
R25988 GND.n7500 GND.n3097 0.152939
R25989 GND.n7496 GND.n3097 0.152939
R25990 GND.n7496 GND.n7495 0.152939
R25991 GND.n7495 GND.n7494 0.152939
R25992 GND.n7494 GND.n3102 0.152939
R25993 GND.n7490 GND.n3102 0.152939
R25994 GND.n7490 GND.n7489 0.152939
R25995 GND.n7489 GND.n7488 0.152939
R25996 GND.n7488 GND.n3107 0.152939
R25997 GND.n7484 GND.n3107 0.152939
R25998 GND.n7484 GND.n7483 0.152939
R25999 GND.n7483 GND.n7482 0.152939
R26000 GND.n7482 GND.n3112 0.152939
R26001 GND.n7478 GND.n3112 0.152939
R26002 GND.n7478 GND.n7477 0.152939
R26003 GND.n7477 GND.n7476 0.152939
R26004 GND.n7476 GND.n3117 0.152939
R26005 GND.n7472 GND.n3117 0.152939
R26006 GND.n7472 GND.n7471 0.152939
R26007 GND.n7471 GND.n7470 0.152939
R26008 GND.n7470 GND.n3122 0.152939
R26009 GND.n7466 GND.n3122 0.152939
R26010 GND.n7466 GND.n7465 0.152939
R26011 GND.n7465 GND.n7464 0.152939
R26012 GND.n7464 GND.n3127 0.152939
R26013 GND.n7460 GND.n3127 0.152939
R26014 GND.n7460 GND.n7459 0.152939
R26015 GND.n7459 GND.n7458 0.152939
R26016 GND.n7458 GND.n3132 0.152939
R26017 GND.n7454 GND.n3132 0.152939
R26018 GND.n7454 GND.n7453 0.152939
R26019 GND.n7453 GND.n7452 0.152939
R26020 GND.n7452 GND.n3137 0.152939
R26021 GND.n7448 GND.n3137 0.152939
R26022 GND.n7448 GND.n7447 0.152939
R26023 GND.n7447 GND.n7446 0.152939
R26024 GND.n7446 GND.n3142 0.152939
R26025 GND.n7442 GND.n3142 0.152939
R26026 GND.n7442 GND.n7441 0.152939
R26027 GND.n7441 GND.n7440 0.152939
R26028 GND.n7440 GND.n3147 0.152939
R26029 GND.n7436 GND.n3147 0.152939
R26030 GND.n7436 GND.n7435 0.152939
R26031 GND.n7435 GND.n7434 0.152939
R26032 GND.n7434 GND.n3152 0.152939
R26033 GND.n7430 GND.n3152 0.152939
R26034 GND.n7430 GND.n7429 0.152939
R26035 GND.n7429 GND.n7428 0.152939
R26036 GND.n7428 GND.n3157 0.152939
R26037 GND.n7424 GND.n3157 0.152939
R26038 GND.n7424 GND.n7423 0.152939
R26039 GND.n7423 GND.n7422 0.152939
R26040 GND.n7422 GND.n3162 0.152939
R26041 GND.n7418 GND.n3162 0.152939
R26042 GND.n7418 GND.n7417 0.152939
R26043 GND.n7417 GND.n7416 0.152939
R26044 GND.n7416 GND.n3167 0.152939
R26045 GND.n7412 GND.n3167 0.152939
R26046 GND.n7412 GND.n7411 0.152939
R26047 GND.n7411 GND.n7410 0.152939
R26048 GND.n7410 GND.n3172 0.152939
R26049 GND.n7406 GND.n3172 0.152939
R26050 GND.n7406 GND.n7405 0.152939
R26051 GND.n7405 GND.n7404 0.152939
R26052 GND.n7404 GND.n3177 0.152939
R26053 GND.n7400 GND.n3177 0.152939
R26054 GND.n7400 GND.n7399 0.152939
R26055 GND.n7399 GND.n7398 0.152939
R26056 GND.n7398 GND.n3182 0.152939
R26057 GND.n7394 GND.n3182 0.152939
R26058 GND.n7394 GND.n7393 0.152939
R26059 GND.n7393 GND.n7392 0.152939
R26060 GND.n7392 GND.n3187 0.152939
R26061 GND.n7388 GND.n3187 0.152939
R26062 GND.n7388 GND.n7387 0.152939
R26063 GND.n7387 GND.n7386 0.152939
R26064 GND.n7386 GND.n3192 0.152939
R26065 GND.n7382 GND.n3192 0.152939
R26066 GND.n7382 GND.n7381 0.152939
R26067 GND.n7381 GND.n7380 0.152939
R26068 GND.n7380 GND.n3197 0.152939
R26069 GND.n7376 GND.n3197 0.152939
R26070 GND.n7376 GND.n7375 0.152939
R26071 GND.n7375 GND.n7374 0.152939
R26072 GND.n7374 GND.n3202 0.152939
R26073 GND.n7370 GND.n3202 0.152939
R26074 GND.n7370 GND.n7369 0.152939
R26075 GND.n7369 GND.n7368 0.152939
R26076 GND.n7368 GND.n3207 0.152939
R26077 GND.n7364 GND.n3207 0.152939
R26078 GND.n7364 GND.n7363 0.152939
R26079 GND.n7363 GND.n7362 0.152939
R26080 GND.n7362 GND.n3212 0.152939
R26081 GND.n7358 GND.n3212 0.152939
R26082 GND.n7358 GND.n7357 0.152939
R26083 GND.n7357 GND.n7356 0.152939
R26084 GND.n7356 GND.n3217 0.152939
R26085 GND.n7352 GND.n3217 0.152939
R26086 GND.n7352 GND.n7351 0.152939
R26087 GND.n7351 GND.n7350 0.152939
R26088 GND.n7350 GND.n3222 0.152939
R26089 GND.n7346 GND.n3222 0.152939
R26090 GND.n7346 GND.n7345 0.152939
R26091 GND.n7345 GND.n7344 0.152939
R26092 GND.n3032 GND.n1887 0.152939
R26093 GND.n3043 GND.n3032 0.152939
R26094 GND.n3044 GND.n3043 0.152939
R26095 GND.n3045 GND.n3044 0.152939
R26096 GND.n3045 GND.n3028 0.152939
R26097 GND.n3050 GND.n3028 0.152939
R26098 GND.n2778 GND.n2188 0.152939
R26099 GND.n2779 GND.n2778 0.152939
R26100 GND.n2780 GND.n2779 0.152939
R26101 GND.n2780 GND.n2095 0.152939
R26102 GND.n2833 GND.n2095 0.152939
R26103 GND.n2834 GND.n2833 0.152939
R26104 GND.n2836 GND.n2834 0.152939
R26105 GND.n2836 GND.n2835 0.152939
R26106 GND.n2835 GND.n2072 0.152939
R26107 GND.n2858 GND.n2072 0.152939
R26108 GND.n2859 GND.n2858 0.152939
R26109 GND.n2861 GND.n2859 0.152939
R26110 GND.n2861 GND.n2860 0.152939
R26111 GND.n2860 GND.n2050 0.152939
R26112 GND.n2883 GND.n2050 0.152939
R26113 GND.n2884 GND.n2883 0.152939
R26114 GND.n2886 GND.n2884 0.152939
R26115 GND.n2886 GND.n2885 0.152939
R26116 GND.n2885 GND.n2023 0.152939
R26117 GND.n7681 GND.n2023 0.152939
R26118 GND.n7682 GND.n7681 0.152939
R26119 GND.n7684 GND.n7682 0.152939
R26120 GND.n7684 GND.n7683 0.152939
R26121 GND.n7683 GND.n1999 0.152939
R26122 GND.n7705 GND.n1999 0.152939
R26123 GND.n7706 GND.n7705 0.152939
R26124 GND.n7708 GND.n7706 0.152939
R26125 GND.n7708 GND.n7707 0.152939
R26126 GND.n7707 GND.n1976 0.152939
R26127 GND.n7730 GND.n1976 0.152939
R26128 GND.n7731 GND.n7730 0.152939
R26129 GND.n7733 GND.n7731 0.152939
R26130 GND.n7733 GND.n7732 0.152939
R26131 GND.n7732 GND.n1954 0.152939
R26132 GND.n7755 GND.n1954 0.152939
R26133 GND.n7756 GND.n7755 0.152939
R26134 GND.n7758 GND.n7756 0.152939
R26135 GND.n7758 GND.n7757 0.152939
R26136 GND.n7757 GND.n1932 0.152939
R26137 GND.n7780 GND.n1932 0.152939
R26138 GND.n7781 GND.n7780 0.152939
R26139 GND.n7783 GND.n7781 0.152939
R26140 GND.n7783 GND.n7782 0.152939
R26141 GND.n7782 GND.n1909 0.152939
R26142 GND.n7804 GND.n1909 0.152939
R26143 GND.n7805 GND.n7804 0.152939
R26144 GND.n7812 GND.n7805 0.152939
R26145 GND.n7812 GND.n7811 0.152939
R26146 GND.n7811 GND.n7810 0.152939
R26147 GND.n7810 GND.n7806 0.152939
R26148 GND.n7806 GND.n1888 0.152939
R26149 GND.n7833 GND.n1888 0.152939
R26150 GND.n7920 GND.n1779 0.152939
R26151 GND.n7916 GND.n1779 0.152939
R26152 GND.n7916 GND.n7915 0.152939
R26153 GND.n7915 GND.n7914 0.152939
R26154 GND.n7914 GND.n1783 0.152939
R26155 GND.n7910 GND.n1783 0.152939
R26156 GND.n7910 GND.n7909 0.152939
R26157 GND.n7909 GND.n7908 0.152939
R26158 GND.n7908 GND.n1788 0.152939
R26159 GND.n7903 GND.n7902 0.152939
R26160 GND.n7902 GND.n7901 0.152939
R26161 GND.n7901 GND.n1798 0.152939
R26162 GND.n7897 GND.n1798 0.152939
R26163 GND.n7897 GND.n7896 0.152939
R26164 GND.n7896 GND.n7895 0.152939
R26165 GND.n7895 GND.n1803 0.152939
R26166 GND.n7891 GND.n1803 0.152939
R26167 GND.n7891 GND.n7890 0.152939
R26168 GND.n7890 GND.n7889 0.152939
R26169 GND.n7889 GND.n1808 0.152939
R26170 GND.n1813 GND.n1808 0.152939
R26171 GND.n7884 GND.n1813 0.152939
R26172 GND.n8098 GND.n1505 0.152939
R26173 GND.n2389 GND.n1505 0.152939
R26174 GND.n2389 GND.n2386 0.152939
R26175 GND.n2395 GND.n2386 0.152939
R26176 GND.n2396 GND.n2395 0.152939
R26177 GND.n2397 GND.n2396 0.152939
R26178 GND.n2397 GND.n2382 0.152939
R26179 GND.n2403 GND.n2382 0.152939
R26180 GND.n2404 GND.n2403 0.152939
R26181 GND.n2405 GND.n2404 0.152939
R26182 GND.n2405 GND.n2375 0.152939
R26183 GND.n2409 GND.n2375 0.152939
R26184 GND.n2411 GND.n2410 0.152939
R26185 GND.n2411 GND.n2373 0.152939
R26186 GND.n2417 GND.n2373 0.152939
R26187 GND.n2418 GND.n2417 0.152939
R26188 GND.n2419 GND.n2418 0.152939
R26189 GND.n2419 GND.n2368 0.152939
R26190 GND.n2517 GND.n2368 0.152939
R26191 GND.n2518 GND.n2517 0.152939
R26192 GND.n2520 GND.n2518 0.152939
R26193 GND.n2520 GND.n2519 0.152939
R26194 GND.n2519 GND.n2346 0.152939
R26195 GND.n2542 GND.n2346 0.152939
R26196 GND.n2543 GND.n2542 0.152939
R26197 GND.n2545 GND.n2543 0.152939
R26198 GND.n2545 GND.n2544 0.152939
R26199 GND.n2544 GND.n2324 0.152939
R26200 GND.n2567 GND.n2324 0.152939
R26201 GND.n2568 GND.n2567 0.152939
R26202 GND.n2570 GND.n2568 0.152939
R26203 GND.n2570 GND.n2569 0.152939
R26204 GND.n2569 GND.n2300 0.152939
R26205 GND.n2591 GND.n2300 0.152939
R26206 GND.n2592 GND.n2591 0.152939
R26207 GND.n2594 GND.n2592 0.152939
R26208 GND.n2594 GND.n2593 0.152939
R26209 GND.n2593 GND.n2277 0.152939
R26210 GND.n2616 GND.n2277 0.152939
R26211 GND.n2617 GND.n2616 0.152939
R26212 GND.n2628 GND.n2617 0.152939
R26213 GND.n2628 GND.n2627 0.152939
R26214 GND.n2627 GND.n2626 0.152939
R26215 GND.n2626 GND.n2618 0.152939
R26216 GND.n2622 GND.n2618 0.152939
R26217 GND.n2622 GND.n2621 0.152939
R26218 GND.n2621 GND.n2236 0.152939
R26219 GND.n2716 GND.n2236 0.152939
R26220 GND.n2717 GND.n2716 0.152939
R26221 GND.n2719 GND.n2717 0.152939
R26222 GND.n2719 GND.n2718 0.152939
R26223 GND.n2718 GND.n2214 0.152939
R26224 GND.n2741 GND.n2214 0.152939
R26225 GND.n2742 GND.n2741 0.152939
R26226 GND.n2744 GND.n2742 0.152939
R26227 GND.n2744 GND.n2743 0.152939
R26228 GND.n2743 GND.n2192 0.152939
R26229 GND.n2763 GND.n2192 0.152939
R26230 GND.n2764 GND.n2763 0.152939
R26231 GND.n2765 GND.n2764 0.152939
R26232 GND.n2765 GND.n2190 0.152939
R26233 GND.n2771 GND.n2190 0.152939
R26234 GND.n2772 GND.n2771 0.152939
R26235 GND.n2774 GND.n2772 0.152939
R26236 GND.n6429 GND.n6428 0.0797683
R26237 GND.n7834 GND.n1887 0.0797683
R26238 GND.n6836 GND.n3744 0.0767195
R26239 GND.n6788 GND.n3744 0.0767195
R26240 GND.n2825 GND.n2824 0.0767195
R26241 GND.n2824 GND.n2106 0.0767195
R26242 GND.n9694 GND.n406 0.0695946
R26243 GND.n9694 GND.n9693 0.0695946
R26244 GND.n2773 GND.n2188 0.0695946
R26245 GND.n2774 GND.n2773 0.0695946
R26246 GND.n6327 GND.n6326 0.0524701
R26247 GND.n9529 GND.n9528 0.0524701
R26248 GND.n8099 GND.n1504 0.0524701
R26249 GND.n7927 GND.n1768 0.0524701
R26250 GND.n6326 GND.n3374 0.0344674
R26251 GND.n7247 GND.n3374 0.0344674
R26252 GND.n7247 GND.n3375 0.0344674
R26253 GND.n7243 GND.n3375 0.0344674
R26254 GND.n7243 GND.n7242 0.0344674
R26255 GND.n7242 GND.n7241 0.0344674
R26256 GND.n7241 GND.n3385 0.0344674
R26257 GND.n7237 GND.n3385 0.0344674
R26258 GND.n7237 GND.n7236 0.0344674
R26259 GND.n7236 GND.n7235 0.0344674
R26260 GND.n7235 GND.n3393 0.0344674
R26261 GND.n7231 GND.n3393 0.0344674
R26262 GND.n7231 GND.n7230 0.0344674
R26263 GND.n7230 GND.n7229 0.0344674
R26264 GND.n7229 GND.n3401 0.0344674
R26265 GND.n7225 GND.n3401 0.0344674
R26266 GND.n7225 GND.n7224 0.0344674
R26267 GND.n7224 GND.n7223 0.0344674
R26268 GND.n7223 GND.n3409 0.0344674
R26269 GND.n7219 GND.n3409 0.0344674
R26270 GND.n7219 GND.n7218 0.0344674
R26271 GND.n7218 GND.n7217 0.0344674
R26272 GND.n7217 GND.n3417 0.0344674
R26273 GND.n7213 GND.n3417 0.0344674
R26274 GND.n7213 GND.n7212 0.0344674
R26275 GND.n7212 GND.n7211 0.0344674
R26276 GND.n7211 GND.n3425 0.0344674
R26277 GND.n7207 GND.n3425 0.0344674
R26278 GND.n7207 GND.n7206 0.0344674
R26279 GND.n7206 GND.n7205 0.0344674
R26280 GND.n7205 GND.n3433 0.0344674
R26281 GND.n7201 GND.n3433 0.0344674
R26282 GND.n7201 GND.n7200 0.0344674
R26283 GND.n7200 GND.n7199 0.0344674
R26284 GND.n7199 GND.n3441 0.0344674
R26285 GND.n7195 GND.n3441 0.0344674
R26286 GND.n7195 GND.n7194 0.0344674
R26287 GND.n7194 GND.n7193 0.0344674
R26288 GND.n7193 GND.n3449 0.0344674
R26289 GND.n7189 GND.n3449 0.0344674
R26290 GND.n7189 GND.n7188 0.0344674
R26291 GND.n7188 GND.n7187 0.0344674
R26292 GND.n7187 GND.n3457 0.0344674
R26293 GND.n7183 GND.n3457 0.0344674
R26294 GND.n7183 GND.n7182 0.0344674
R26295 GND.n7182 GND.n7181 0.0344674
R26296 GND.n7181 GND.n3465 0.0344674
R26297 GND.n7177 GND.n3465 0.0344674
R26298 GND.n7177 GND.n7176 0.0344674
R26299 GND.n7176 GND.n7175 0.0344674
R26300 GND.n7175 GND.n3473 0.0344674
R26301 GND.n7171 GND.n3473 0.0344674
R26302 GND.n7171 GND.n7170 0.0344674
R26303 GND.n7170 GND.n7169 0.0344674
R26304 GND.n7169 GND.n3481 0.0344674
R26305 GND.n7165 GND.n3481 0.0344674
R26306 GND.n7165 GND.n7164 0.0344674
R26307 GND.n7164 GND.n7163 0.0344674
R26308 GND.n7163 GND.n3489 0.0344674
R26309 GND.n7159 GND.n3489 0.0344674
R26310 GND.n7159 GND.n7158 0.0344674
R26311 GND.n7158 GND.n7157 0.0344674
R26312 GND.n7157 GND.n3497 0.0344674
R26313 GND.n7153 GND.n3497 0.0344674
R26314 GND.n7153 GND.n7152 0.0344674
R26315 GND.n7152 GND.n7151 0.0344674
R26316 GND.n7151 GND.n3505 0.0344674
R26317 GND.n7147 GND.n3505 0.0344674
R26318 GND.n7147 GND.n7146 0.0344674
R26319 GND.n7146 GND.n7145 0.0344674
R26320 GND.n7145 GND.n3513 0.0344674
R26321 GND.n7141 GND.n3513 0.0344674
R26322 GND.n7141 GND.n7140 0.0344674
R26323 GND.n7140 GND.n7139 0.0344674
R26324 GND.n7139 GND.n3521 0.0344674
R26325 GND.n7135 GND.n3521 0.0344674
R26326 GND.n7135 GND.n7134 0.0344674
R26327 GND.n7134 GND.n7133 0.0344674
R26328 GND.n7133 GND.n3529 0.0344674
R26329 GND.n7129 GND.n3529 0.0344674
R26330 GND.n7129 GND.n7128 0.0344674
R26331 GND.n7128 GND.n7127 0.0344674
R26332 GND.n7127 GND.n3537 0.0344674
R26333 GND.n7123 GND.n3537 0.0344674
R26334 GND.n7123 GND.n7122 0.0344674
R26335 GND.n7122 GND.n7121 0.0344674
R26336 GND.n7121 GND.n3545 0.0344674
R26337 GND.n7117 GND.n3545 0.0344674
R26338 GND.n7117 GND.n7116 0.0344674
R26339 GND.n7116 GND.n7115 0.0344674
R26340 GND.n7115 GND.n3553 0.0344674
R26341 GND.n7111 GND.n3553 0.0344674
R26342 GND.n7111 GND.n7110 0.0344674
R26343 GND.n7110 GND.n7109 0.0344674
R26344 GND.n7109 GND.n3561 0.0344674
R26345 GND.n7105 GND.n3561 0.0344674
R26346 GND.n7105 GND.n7104 0.0344674
R26347 GND.n7104 GND.n7103 0.0344674
R26348 GND.n7103 GND.n576 0.0344674
R26349 GND.n9503 GND.n576 0.0344674
R26350 GND.n9503 GND.n554 0.0344674
R26351 GND.n9519 GND.n554 0.0344674
R26352 GND.n9520 GND.n9519 0.0344674
R26353 GND.n9520 GND.n547 0.0344674
R26354 GND.n9528 GND.n547 0.0344674
R26355 GND.n1562 GND.n1504 0.0344674
R26356 GND.n1562 GND.n1557 0.0344674
R26357 GND.n1567 GND.n1557 0.0344674
R26358 GND.n1567 GND.n1554 0.0344674
R26359 GND.n8077 GND.n1554 0.0344674
R26360 GND.n8077 GND.n1555 0.0344674
R26361 GND.n8073 GND.n1555 0.0344674
R26362 GND.n8073 GND.n8072 0.0344674
R26363 GND.n8072 GND.n8071 0.0344674
R26364 GND.n8071 GND.n1576 0.0344674
R26365 GND.n8067 GND.n1576 0.0344674
R26366 GND.n8067 GND.n8066 0.0344674
R26367 GND.n8066 GND.n8065 0.0344674
R26368 GND.n8065 GND.n1584 0.0344674
R26369 GND.n8061 GND.n1584 0.0344674
R26370 GND.n8061 GND.n8060 0.0344674
R26371 GND.n8060 GND.n8059 0.0344674
R26372 GND.n8059 GND.n1592 0.0344674
R26373 GND.n8055 GND.n1592 0.0344674
R26374 GND.n8055 GND.n8054 0.0344674
R26375 GND.n8054 GND.n8053 0.0344674
R26376 GND.n8053 GND.n1600 0.0344674
R26377 GND.n8049 GND.n1600 0.0344674
R26378 GND.n8049 GND.n8048 0.0344674
R26379 GND.n8048 GND.n8047 0.0344674
R26380 GND.n8047 GND.n1608 0.0344674
R26381 GND.n8043 GND.n1608 0.0344674
R26382 GND.n8043 GND.n8042 0.0344674
R26383 GND.n8042 GND.n8041 0.0344674
R26384 GND.n8041 GND.n1616 0.0344674
R26385 GND.n8037 GND.n1616 0.0344674
R26386 GND.n8037 GND.n8036 0.0344674
R26387 GND.n8036 GND.n8035 0.0344674
R26388 GND.n8035 GND.n1624 0.0344674
R26389 GND.n8031 GND.n1624 0.0344674
R26390 GND.n8031 GND.n8030 0.0344674
R26391 GND.n8030 GND.n8029 0.0344674
R26392 GND.n8029 GND.n1632 0.0344674
R26393 GND.n8025 GND.n1632 0.0344674
R26394 GND.n8025 GND.n8024 0.0344674
R26395 GND.n8024 GND.n8023 0.0344674
R26396 GND.n8023 GND.n1640 0.0344674
R26397 GND.n8019 GND.n1640 0.0344674
R26398 GND.n8019 GND.n8018 0.0344674
R26399 GND.n8018 GND.n8017 0.0344674
R26400 GND.n8017 GND.n1648 0.0344674
R26401 GND.n8013 GND.n1648 0.0344674
R26402 GND.n8013 GND.n8012 0.0344674
R26403 GND.n8012 GND.n8011 0.0344674
R26404 GND.n8011 GND.n1656 0.0344674
R26405 GND.n8007 GND.n1656 0.0344674
R26406 GND.n8007 GND.n8006 0.0344674
R26407 GND.n8006 GND.n8005 0.0344674
R26408 GND.n8005 GND.n1664 0.0344674
R26409 GND.n8001 GND.n1664 0.0344674
R26410 GND.n8001 GND.n8000 0.0344674
R26411 GND.n8000 GND.n7999 0.0344674
R26412 GND.n7999 GND.n1672 0.0344674
R26413 GND.n7995 GND.n1672 0.0344674
R26414 GND.n7995 GND.n7994 0.0344674
R26415 GND.n7994 GND.n7993 0.0344674
R26416 GND.n7993 GND.n1680 0.0344674
R26417 GND.n7989 GND.n1680 0.0344674
R26418 GND.n7989 GND.n7988 0.0344674
R26419 GND.n7988 GND.n7987 0.0344674
R26420 GND.n7987 GND.n1688 0.0344674
R26421 GND.n7983 GND.n1688 0.0344674
R26422 GND.n7983 GND.n7982 0.0344674
R26423 GND.n7982 GND.n7981 0.0344674
R26424 GND.n7981 GND.n1696 0.0344674
R26425 GND.n7977 GND.n1696 0.0344674
R26426 GND.n7977 GND.n7976 0.0344674
R26427 GND.n7976 GND.n7975 0.0344674
R26428 GND.n7975 GND.n1704 0.0344674
R26429 GND.n7971 GND.n1704 0.0344674
R26430 GND.n7971 GND.n7970 0.0344674
R26431 GND.n7970 GND.n7969 0.0344674
R26432 GND.n7969 GND.n1712 0.0344674
R26433 GND.n7965 GND.n1712 0.0344674
R26434 GND.n7965 GND.n7964 0.0344674
R26435 GND.n7964 GND.n7963 0.0344674
R26436 GND.n7963 GND.n1720 0.0344674
R26437 GND.n7959 GND.n1720 0.0344674
R26438 GND.n7959 GND.n7958 0.0344674
R26439 GND.n7958 GND.n7957 0.0344674
R26440 GND.n7957 GND.n1728 0.0344674
R26441 GND.n7953 GND.n1728 0.0344674
R26442 GND.n7953 GND.n7952 0.0344674
R26443 GND.n7952 GND.n7951 0.0344674
R26444 GND.n7951 GND.n1736 0.0344674
R26445 GND.n7947 GND.n1736 0.0344674
R26446 GND.n7947 GND.n7946 0.0344674
R26447 GND.n7946 GND.n7945 0.0344674
R26448 GND.n7945 GND.n1744 0.0344674
R26449 GND.n7941 GND.n1744 0.0344674
R26450 GND.n7941 GND.n7940 0.0344674
R26451 GND.n7940 GND.n7939 0.0344674
R26452 GND.n7939 GND.n1752 0.0344674
R26453 GND.n7935 GND.n1752 0.0344674
R26454 GND.n7935 GND.n7934 0.0344674
R26455 GND.n7934 GND.n7933 0.0344674
R26456 GND.n7933 GND.n1760 0.0344674
R26457 GND.n7929 GND.n1760 0.0344674
R26458 GND.n7929 GND.n7928 0.0344674
R26459 GND.n7928 GND.n7927 0.0344674
R26460 GND.n3317 GND.n3315 0.00731034
R26461 GND.n7289 GND.n7288 0.00731034
R26462 GND.n7285 GND.n3318 0.00731034
R26463 GND.n7284 GND.n3323 0.00731034
R26464 GND.n7281 GND.n7280 0.00731034
R26465 GND.n7277 GND.n3329 0.00731034
R26466 GND.n7276 GND.n3333 0.00731034
R26467 GND.n7273 GND.n7272 0.00731034
R26468 GND.n7269 GND.n3337 0.00731034
R26469 GND.n7268 GND.n3341 0.00731034
R26470 GND.n7265 GND.n7264 0.00731034
R26471 GND.n7261 GND.n3349 0.00731034
R26472 GND.n7260 GND.n3353 0.00731034
R26473 GND.n7871 GND.n7870 0.00731034
R26474 GND.n1852 GND.n1835 0.00731034
R26475 GND.n7863 GND.n1853 0.00731034
R26476 GND.n7862 GND.n1854 0.00731034
R26477 GND.n7859 GND.n7858 0.00731034
R26478 GND.n7855 GND.n1861 0.00731034
R26479 GND.n7854 GND.n1865 0.00731034
R26480 GND.n7851 GND.n7850 0.00731034
R26481 GND.n7847 GND.n1869 0.00731034
R26482 GND.n7846 GND.n1875 0.00731034
R26483 GND.n7843 GND.n7842 0.00731034
R26484 GND.n7839 GND.n1883 0.00731034
R26485 GND.n7838 GND.n7835 0.00731034
R26486 GND.n6328 GND.n3315 0.00713793
R26487 GND.n7871 GND.n1834 0.00713793
R26488 GND.n6429 GND.n3353 0.00463793
R26489 GND.n7835 GND.n7834 0.00463793
R26490 GND.n7289 GND.n3317 0.00231034
R26491 GND.n7288 GND.n3318 0.00231034
R26492 GND.n7285 GND.n7284 0.00231034
R26493 GND.n7281 GND.n3323 0.00231034
R26494 GND.n7280 GND.n3329 0.00231034
R26495 GND.n7277 GND.n7276 0.00231034
R26496 GND.n7273 GND.n3333 0.00231034
R26497 GND.n7272 GND.n3337 0.00231034
R26498 GND.n7269 GND.n7268 0.00231034
R26499 GND.n7265 GND.n3341 0.00231034
R26500 GND.n7264 GND.n3349 0.00231034
R26501 GND.n7261 GND.n7260 0.00231034
R26502 GND.n7870 GND.n1835 0.00231034
R26503 GND.n1853 GND.n1852 0.00231034
R26504 GND.n7863 GND.n7862 0.00231034
R26505 GND.n7859 GND.n1854 0.00231034
R26506 GND.n7858 GND.n1861 0.00231034
R26507 GND.n7855 GND.n7854 0.00231034
R26508 GND.n7851 GND.n1865 0.00231034
R26509 GND.n7850 GND.n1869 0.00231034
R26510 GND.n7847 GND.n7846 0.00231034
R26511 GND.n7843 GND.n1875 0.00231034
R26512 GND.n7842 GND.n1883 0.00231034
R26513 GND.n7839 GND.n7838 0.00231034
R26514 VOUT.n23 VOUT.t8 126.343
R26515 VOUT.n17 VOUT.t7 126.343
R26516 VOUT.n11 VOUT.t14 123.921
R26517 VOUT.n5 VOUT.t50 123.921
R26518 VOUT.n8 VOUT.n6 119.736
R26519 VOUT.n2 VOUT.n0 119.736
R26520 VOUT.n25 VOUT.n24 117.314
R26521 VOUT.n23 VOUT.n22 117.314
R26522 VOUT.n21 VOUT.n20 117.314
R26523 VOUT.n19 VOUT.n18 117.314
R26524 VOUT.n17 VOUT.n16 117.314
R26525 VOUT.n8 VOUT.n7 117.314
R26526 VOUT.n10 VOUT.n9 117.314
R26527 VOUT.n2 VOUT.n1 117.314
R26528 VOUT.n4 VOUT.n3 117.314
R26529 VOUT.n27 VOUT.n26 117.314
R26530 VOUT.n37 VOUT.n35 91.4836
R26531 VOUT.n32 VOUT.n30 91.4836
R26532 VOUT.n49 VOUT.n47 91.4836
R26533 VOUT.n44 VOUT.n42 91.4836
R26534 VOUT.n39 VOUT.n38 88.7853
R26535 VOUT.n37 VOUT.n36 88.7853
R26536 VOUT.n34 VOUT.n33 88.7853
R26537 VOUT.n32 VOUT.n31 88.7853
R26538 VOUT.n49 VOUT.n48 88.7853
R26539 VOUT.n51 VOUT.n50 88.7853
R26540 VOUT.n44 VOUT.n43 88.7853
R26541 VOUT.n46 VOUT.n45 88.7853
R26542 VOUT.n41 VOUT.n29 8.67473
R26543 VOUT.n28 VOUT.n21 7.84964
R26544 VOUT.n40 VOUT.n34 7.73757
R26545 VOUT.n52 VOUT.n46 7.73757
R26546 VOUT.n12 VOUT.n5 6.63843
R26547 VOUT.n26 VOUT.t6 6.60721
R26548 VOUT.n26 VOUT.t1 6.60721
R26549 VOUT.n24 VOUT.t17 6.60721
R26550 VOUT.n24 VOUT.t2 6.60721
R26551 VOUT.n22 VOUT.t15 6.60721
R26552 VOUT.n22 VOUT.t10 6.60721
R26553 VOUT.n20 VOUT.t0 6.60721
R26554 VOUT.n20 VOUT.t9 6.60721
R26555 VOUT.n18 VOUT.t4 6.60721
R26556 VOUT.n18 VOUT.t11 6.60721
R26557 VOUT.n16 VOUT.t12 6.60721
R26558 VOUT.n16 VOUT.t42 6.60721
R26559 VOUT.n6 VOUT.t16 6.60721
R26560 VOUT.n6 VOUT.t47 6.60721
R26561 VOUT.n7 VOUT.t49 6.60721
R26562 VOUT.n7 VOUT.t13 6.60721
R26563 VOUT.n9 VOUT.t3 6.60721
R26564 VOUT.n9 VOUT.t48 6.60721
R26565 VOUT.n0 VOUT.t45 6.60721
R26566 VOUT.n0 VOUT.t44 6.60721
R26567 VOUT.n1 VOUT.t5 6.60721
R26568 VOUT.n1 VOUT.t51 6.60721
R26569 VOUT.n3 VOUT.t46 6.60721
R26570 VOUT.n3 VOUT.t43 6.60721
R26571 VOUT.n40 VOUT.n39 6.31516
R26572 VOUT.n52 VOUT.n51 6.31516
R26573 VOUT.n28 VOUT.n27 6.17722
R26574 VOUT.n29 VOUT.n13 6.11583
R26575 VOUT.n41 VOUT.n40 5.89326
R26576 VOUT.n53 VOUT.n52 5.89326
R26577 VOUT.n29 VOUT.n28 5.80059
R26578 VOUT.n13 VOUT.n12 5.80059
R26579 VOUT.n53 VOUT.n41 5.68625
R26580 VOUT.n38 VOUT.t34 5.26646
R26581 VOUT.n38 VOUT.t28 5.26646
R26582 VOUT.n36 VOUT.t26 5.26646
R26583 VOUT.n36 VOUT.t19 5.26646
R26584 VOUT.n35 VOUT.t38 5.26646
R26585 VOUT.n35 VOUT.t30 5.26646
R26586 VOUT.n33 VOUT.t39 5.26646
R26587 VOUT.n33 VOUT.t29 5.26646
R26588 VOUT.n31 VOUT.t36 5.26646
R26589 VOUT.n31 VOUT.t24 5.26646
R26590 VOUT.n30 VOUT.t32 5.26646
R26591 VOUT.n30 VOUT.t23 5.26646
R26592 VOUT.n47 VOUT.t20 5.26646
R26593 VOUT.n47 VOUT.t25 5.26646
R26594 VOUT.n48 VOUT.t35 5.26646
R26595 VOUT.n48 VOUT.t33 5.26646
R26596 VOUT.n50 VOUT.t40 5.26646
R26597 VOUT.n50 VOUT.t21 5.26646
R26598 VOUT.n42 VOUT.t27 5.26646
R26599 VOUT.n42 VOUT.t37 5.26646
R26600 VOUT.n43 VOUT.t22 5.26646
R26601 VOUT.n43 VOUT.t41 5.26646
R26602 VOUT.n45 VOUT.t31 5.26646
R26603 VOUT.n45 VOUT.t18 5.26646
R26604 VOUT.n12 VOUT.n11 4.96602
R26605 VOUT.n54 VOUT.n13 4.73136
R26606 VOUT.n54 VOUT.n53 3.92437
R26607 VOUT.n15 VOUT 3.01085
R26608 VOUT.n39 VOUT.n37 2.69878
R26609 VOUT.n34 VOUT.n32 2.69878
R26610 VOUT.n51 VOUT.n49 2.69878
R26611 VOUT.n46 VOUT.n44 2.69878
R26612 VOUT.n25 VOUT.n23 2.42291
R26613 VOUT.n27 VOUT.n25 2.42291
R26614 VOUT.n19 VOUT.n17 2.42291
R26615 VOUT.n21 VOUT.n19 2.42291
R26616 VOUT.n11 VOUT.n10 2.42291
R26617 VOUT.n10 VOUT.n8 2.42291
R26618 VOUT.n5 VOUT.n4 2.42291
R26619 VOUT.n4 VOUT.n2 2.42291
R26620 VOUT.n15 VOUT.n14 0.332206
R26621 VOUT.n54 VOUT.n15 0.292135
R26622 VOUT.n14 VOUT.t53 0.210394
R26623 VOUT.n14 VOUT.t52 0.124973
R26624 VOUT VOUT.n54 0.0099
R26625 VN.n160 VN.t0 243.97
R26626 VN.n160 VN.n159 223.454
R26627 VN.n162 VN.n161 223.454
R26628 VN.n155 VN.n79 161.3
R26629 VN.n154 VN.n153 161.3
R26630 VN.n152 VN.n80 161.3
R26631 VN.n151 VN.n150 161.3
R26632 VN.n149 VN.n81 161.3
R26633 VN.n148 VN.n147 161.3
R26634 VN.n146 VN.n82 161.3
R26635 VN.n145 VN.n144 161.3
R26636 VN.n143 VN.n83 161.3
R26637 VN.n142 VN.n141 161.3
R26638 VN.n140 VN.n84 161.3
R26639 VN.n139 VN.n138 161.3
R26640 VN.n136 VN.n85 161.3
R26641 VN.n135 VN.n134 161.3
R26642 VN.n133 VN.n86 161.3
R26643 VN.n132 VN.n131 161.3
R26644 VN.n130 VN.n87 161.3
R26645 VN.n129 VN.n128 161.3
R26646 VN.n127 VN.n88 161.3
R26647 VN.n126 VN.n125 161.3
R26648 VN.n124 VN.n89 161.3
R26649 VN.n123 VN.n122 161.3
R26650 VN.n121 VN.n90 161.3
R26651 VN.n120 VN.n119 161.3
R26652 VN.n118 VN.n91 161.3
R26653 VN.n117 VN.n116 161.3
R26654 VN.n115 VN.n92 161.3
R26655 VN.n114 VN.n113 161.3
R26656 VN.n112 VN.n93 161.3
R26657 VN.n111 VN.n110 161.3
R26658 VN.n109 VN.n94 161.3
R26659 VN.n108 VN.n107 161.3
R26660 VN.n106 VN.n95 161.3
R26661 VN.n105 VN.n104 161.3
R26662 VN.n103 VN.n96 161.3
R26663 VN.n102 VN.n101 161.3
R26664 VN.n100 VN.n97 161.3
R26665 VN.n21 VN.n18 161.3
R26666 VN.n23 VN.n22 161.3
R26667 VN.n24 VN.n17 161.3
R26668 VN.n26 VN.n25 161.3
R26669 VN.n27 VN.n16 161.3
R26670 VN.n29 VN.n28 161.3
R26671 VN.n30 VN.n15 161.3
R26672 VN.n32 VN.n31 161.3
R26673 VN.n33 VN.n14 161.3
R26674 VN.n35 VN.n34 161.3
R26675 VN.n36 VN.n13 161.3
R26676 VN.n38 VN.n37 161.3
R26677 VN.n39 VN.n12 161.3
R26678 VN.n41 VN.n40 161.3
R26679 VN.n42 VN.n11 161.3
R26680 VN.n44 VN.n43 161.3
R26681 VN.n45 VN.n10 161.3
R26682 VN.n47 VN.n46 161.3
R26683 VN.n48 VN.n9 161.3
R26684 VN.n50 VN.n49 161.3
R26685 VN.n51 VN.n8 161.3
R26686 VN.n53 VN.n52 161.3
R26687 VN.n54 VN.n7 161.3
R26688 VN.n56 VN.n55 161.3
R26689 VN.n57 VN.n6 161.3
R26690 VN.n60 VN.n59 161.3
R26691 VN.n61 VN.n5 161.3
R26692 VN.n63 VN.n62 161.3
R26693 VN.n64 VN.n4 161.3
R26694 VN.n66 VN.n65 161.3
R26695 VN.n67 VN.n3 161.3
R26696 VN.n69 VN.n68 161.3
R26697 VN.n70 VN.n2 161.3
R26698 VN.n72 VN.n71 161.3
R26699 VN.n73 VN.n1 161.3
R26700 VN.n75 VN.n74 161.3
R26701 VN.n76 VN.n0 161.3
R26702 VN.n99 VN.n98 65.7373
R26703 VN.n20 VN.n19 65.7373
R26704 VN.n157 VN.n156 56.8746
R26705 VN.n78 VN.n77 56.8746
R26706 VN.n148 VN.n82 56.5617
R26707 VN.n69 VN.n3 56.5617
R26708 VN.n158 VN.n157 52.4067
R26709 VN.n107 VN.n94 50.7491
R26710 VN.n129 VN.n88 50.7491
R26711 VN.n50 VN.n9 50.7491
R26712 VN.n28 VN.n15 50.7491
R26713 VN.n98 VN.t9 46.6743
R26714 VN.n19 VN.t12 46.6739
R26715 VN.n111 VN.n94 30.405
R26716 VN.n125 VN.n88 30.405
R26717 VN.n46 VN.n9 30.405
R26718 VN.n32 VN.n15 30.405
R26719 VN.n101 VN.n100 24.5923
R26720 VN.n101 VN.n96 24.5923
R26721 VN.n105 VN.n96 24.5923
R26722 VN.n106 VN.n105 24.5923
R26723 VN.n107 VN.n106 24.5923
R26724 VN.n112 VN.n111 24.5923
R26725 VN.n113 VN.n112 24.5923
R26726 VN.n113 VN.n92 24.5923
R26727 VN.n117 VN.n92 24.5923
R26728 VN.n118 VN.n117 24.5923
R26729 VN.n119 VN.n118 24.5923
R26730 VN.n119 VN.n90 24.5923
R26731 VN.n123 VN.n90 24.5923
R26732 VN.n124 VN.n123 24.5923
R26733 VN.n125 VN.n124 24.5923
R26734 VN.n130 VN.n129 24.5923
R26735 VN.n131 VN.n130 24.5923
R26736 VN.n131 VN.n86 24.5923
R26737 VN.n135 VN.n86 24.5923
R26738 VN.n136 VN.n135 24.5923
R26739 VN.n138 VN.n84 24.5923
R26740 VN.n142 VN.n84 24.5923
R26741 VN.n143 VN.n142 24.5923
R26742 VN.n144 VN.n143 24.5923
R26743 VN.n144 VN.n82 24.5923
R26744 VN.n149 VN.n148 24.5923
R26745 VN.n150 VN.n149 24.5923
R26746 VN.n150 VN.n80 24.5923
R26747 VN.n154 VN.n80 24.5923
R26748 VN.n155 VN.n154 24.5923
R26749 VN.n76 VN.n75 24.5923
R26750 VN.n75 VN.n1 24.5923
R26751 VN.n71 VN.n1 24.5923
R26752 VN.n71 VN.n70 24.5923
R26753 VN.n70 VN.n69 24.5923
R26754 VN.n65 VN.n3 24.5923
R26755 VN.n65 VN.n64 24.5923
R26756 VN.n64 VN.n63 24.5923
R26757 VN.n63 VN.n5 24.5923
R26758 VN.n59 VN.n5 24.5923
R26759 VN.n57 VN.n56 24.5923
R26760 VN.n56 VN.n7 24.5923
R26761 VN.n52 VN.n7 24.5923
R26762 VN.n52 VN.n51 24.5923
R26763 VN.n51 VN.n50 24.5923
R26764 VN.n46 VN.n45 24.5923
R26765 VN.n45 VN.n44 24.5923
R26766 VN.n44 VN.n11 24.5923
R26767 VN.n40 VN.n11 24.5923
R26768 VN.n40 VN.n39 24.5923
R26769 VN.n39 VN.n38 24.5923
R26770 VN.n38 VN.n13 24.5923
R26771 VN.n34 VN.n13 24.5923
R26772 VN.n34 VN.n33 24.5923
R26773 VN.n33 VN.n32 24.5923
R26774 VN.n28 VN.n27 24.5923
R26775 VN.n27 VN.n26 24.5923
R26776 VN.n26 VN.n17 24.5923
R26777 VN.n22 VN.n17 24.5923
R26778 VN.n22 VN.n21 24.5923
R26779 VN.n156 VN.n155 20.6576
R26780 VN.n77 VN.n76 20.6576
R26781 VN.n159 VN.t1 19.8005
R26782 VN.n159 VN.t3 19.8005
R26783 VN.n161 VN.t2 19.8005
R26784 VN.n161 VN.t4 19.8005
R26785 VN VN.n163 19.355
R26786 VN.n138 VN.n137 14.2638
R26787 VN.n59 VN.n58 14.2638
R26788 VN.n118 VN.t13 13.608
R26789 VN.n99 VN.t5 13.608
R26790 VN.n137 VN.t14 13.608
R26791 VN.n156 VN.t11 13.608
R26792 VN.n39 VN.t10 13.608
R26793 VN.n77 VN.t8 13.608
R26794 VN.n58 VN.t7 13.608
R26795 VN.n20 VN.t6 13.608
R26796 VN.n158 VN.n78 13.0241
R26797 VN.n100 VN.n99 10.3291
R26798 VN.n137 VN.n136 10.3291
R26799 VN.n58 VN.n57 10.3291
R26800 VN.n21 VN.n20 10.3291
R26801 VN.n163 VN.n162 5.40567
R26802 VN.n163 VN.n158 1.188
R26803 VN.n98 VN.n97 0.993426
R26804 VN.n19 VN.n18 0.993421
R26805 VN.n162 VN.n160 0.716017
R26806 VN.n157 VN.n79 0.502096
R26807 VN.n78 VN.n0 0.502096
R26808 VN.n102 VN.n97 0.189894
R26809 VN.n103 VN.n102 0.189894
R26810 VN.n104 VN.n103 0.189894
R26811 VN.n104 VN.n95 0.189894
R26812 VN.n108 VN.n95 0.189894
R26813 VN.n109 VN.n108 0.189894
R26814 VN.n110 VN.n109 0.189894
R26815 VN.n110 VN.n93 0.189894
R26816 VN.n114 VN.n93 0.189894
R26817 VN.n115 VN.n114 0.189894
R26818 VN.n116 VN.n115 0.189894
R26819 VN.n116 VN.n91 0.189894
R26820 VN.n120 VN.n91 0.189894
R26821 VN.n121 VN.n120 0.189894
R26822 VN.n122 VN.n121 0.189894
R26823 VN.n122 VN.n89 0.189894
R26824 VN.n126 VN.n89 0.189894
R26825 VN.n127 VN.n126 0.189894
R26826 VN.n128 VN.n127 0.189894
R26827 VN.n128 VN.n87 0.189894
R26828 VN.n132 VN.n87 0.189894
R26829 VN.n133 VN.n132 0.189894
R26830 VN.n134 VN.n133 0.189894
R26831 VN.n134 VN.n85 0.189894
R26832 VN.n139 VN.n85 0.189894
R26833 VN.n140 VN.n139 0.189894
R26834 VN.n141 VN.n140 0.189894
R26835 VN.n141 VN.n83 0.189894
R26836 VN.n145 VN.n83 0.189894
R26837 VN.n146 VN.n145 0.189894
R26838 VN.n147 VN.n146 0.189894
R26839 VN.n147 VN.n81 0.189894
R26840 VN.n151 VN.n81 0.189894
R26841 VN.n152 VN.n151 0.189894
R26842 VN.n153 VN.n152 0.189894
R26843 VN.n153 VN.n79 0.189894
R26844 VN.n74 VN.n0 0.189894
R26845 VN.n74 VN.n73 0.189894
R26846 VN.n73 VN.n72 0.189894
R26847 VN.n72 VN.n2 0.189894
R26848 VN.n68 VN.n2 0.189894
R26849 VN.n68 VN.n67 0.189894
R26850 VN.n67 VN.n66 0.189894
R26851 VN.n66 VN.n4 0.189894
R26852 VN.n62 VN.n4 0.189894
R26853 VN.n62 VN.n61 0.189894
R26854 VN.n61 VN.n60 0.189894
R26855 VN.n60 VN.n6 0.189894
R26856 VN.n55 VN.n6 0.189894
R26857 VN.n55 VN.n54 0.189894
R26858 VN.n54 VN.n53 0.189894
R26859 VN.n53 VN.n8 0.189894
R26860 VN.n49 VN.n8 0.189894
R26861 VN.n49 VN.n48 0.189894
R26862 VN.n48 VN.n47 0.189894
R26863 VN.n47 VN.n10 0.189894
R26864 VN.n43 VN.n10 0.189894
R26865 VN.n43 VN.n42 0.189894
R26866 VN.n42 VN.n41 0.189894
R26867 VN.n41 VN.n12 0.189894
R26868 VN.n37 VN.n12 0.189894
R26869 VN.n37 VN.n36 0.189894
R26870 VN.n36 VN.n35 0.189894
R26871 VN.n35 VN.n14 0.189894
R26872 VN.n31 VN.n14 0.189894
R26873 VN.n31 VN.n30 0.189894
R26874 VN.n30 VN.n29 0.189894
R26875 VN.n29 VN.n16 0.189894
R26876 VN.n25 VN.n16 0.189894
R26877 VN.n25 VN.n24 0.189894
R26878 VN.n24 VN.n23 0.189894
R26879 VN.n23 VN.n18 0.189894
R26880 a_n18960_7900.t11 a_n18960_7900.n17 154.475
R26881 a_n18960_7900.n15 a_n18960_7900.n6 2.49614
R26882 a_n18960_7900.n16 a_n18960_7900.n8 2.49614
R26883 a_n18960_7900.t0 a_n18960_7900.n19 133.071
R26884 a_n18960_7900.n18 a_n18960_7900.t4 131.248
R26885 a_n18960_7900.n18 a_n18960_7900.t5 125.144
R26886 a_n18960_7900.n19 a_n18960_7900.t7 123.32
R26887 a_n18960_7900.n19 a_n18960_7900.t1 123.32
R26888 a_n18960_7900.n18 a_n18960_7900.t19 123.32
R26889 a_n18960_7900.n20 a_n18960_7900.t15 100.508
R26890 a_n18960_7900.n17 a_n18960_7900.t8 98.5007
R26891 a_n18960_7900.n17 a_n18960_7900.t17 98.5007
R26892 a_n18960_7900.n20 a_n18960_7900.t16 98.5006
R26893 a_n18960_7900.n20 a_n18960_7900.t10 155.919
R26894 a_n18960_7900.n6 a_n18960_7900.t37 55.7919
R26895 a_n18960_7900.n8 a_n18960_7900.t47 55.7919
R26896 a_n18960_7900.n3 a_n18960_7900.t29 55.7918
R26897 a_n18960_7900.n1 a_n18960_7900.t41 55.7918
R26898 a_n18960_7900.n7 a_n18960_7900.n6 3.39951
R26899 a_n18960_7900.n11 a_n18960_7900.n6 1.94637
R26900 a_n18960_7900.n22 a_n18960_7900.n11 64.9704
R26901 a_n18960_7900.n9 a_n18960_7900.n8 3.39951
R26902 a_n18960_7900.n10 a_n18960_7900.n8 1.94637
R26903 a_n18960_7900.n21 a_n18960_7900.n10 64.9704
R26904 a_n18960_7900.n3 a_n18960_7900.t25 51.6583
R26905 a_n18960_7900.n3 a_n18960_7900.t44 54.4407
R26906 a_n18960_7900.n5 a_n18960_7900.t46 52.8822
R26907 a_n18960_7900.n5 a_n18960_7900.t23 56.3213
R26908 a_n18960_7900.n2 a_n18960_7900.t26 53.0337
R26909 a_n18960_7900.n2 a_n18960_7900.t27 57.3766
R26910 a_n18960_7900.n1 a_n18960_7900.t36 51.6583
R26911 a_n18960_7900.n1 a_n18960_7900.t22 54.4407
R26912 a_n18960_7900.n4 a_n18960_7900.t24 52.8822
R26913 a_n18960_7900.n4 a_n18960_7900.t34 56.3213
R26914 a_n18960_7900.n0 a_n18960_7900.t38 53.0337
R26915 a_n18960_7900.n0 a_n18960_7900.t39 57.3766
R26916 a_n18960_7900.n7 a_n18960_7900.t31 54.6822
R26917 a_n18960_7900.n6 a_n18960_7900.t35 53.7391
R26918 a_n18960_7900.n7 a_n18960_7900.t33 53.0357
R26919 a_n18960_7900.n11 a_n18960_7900.t21 52.6984
R26920 a_n18960_7900.n22 a_n18960_7900.t28 22.4149
R26921 a_n18960_7900.n15 a_n18960_7900.t20 55.3031
R26922 a_n18960_7900.n9 a_n18960_7900.t42 54.6822
R26923 a_n18960_7900.n8 a_n18960_7900.t45 53.7391
R26924 a_n18960_7900.n9 a_n18960_7900.t43 53.0357
R26925 a_n18960_7900.n10 a_n18960_7900.t32 52.6984
R26926 a_n18960_7900.n21 a_n18960_7900.t40 22.4149
R26927 a_n18960_7900.n16 a_n18960_7900.t30 55.3031
R26928 a_n18960_7900.n3 a_n18960_7900.n5 2.9507
R26929 a_n18960_7900.n1 a_n18960_7900.n4 2.9507
R26930 a_n18960_7900.n15 a_n18960_7900.n22 63.7654
R26931 a_n18960_7900.n16 a_n18960_7900.n21 63.7654
R26932 a_n18960_7900.n23 a_n18960_7900.n14 11.4887
R26933 a_n18960_7900.n14 a_n18960_7900.n12 8.67506
R26934 a_n18960_7900.n13 a_n18960_7900.n1 8.36713
R26935 a_n18960_7900.n12 a_n18960_7900.n8 8.36713
R26936 a_n18960_7900.t7 a_n18960_7900.t18 7.92855
R26937 a_n18960_7900.t1 a_n18960_7900.t2 7.92855
R26938 a_n18960_7900.t5 a_n18960_7900.t3 7.92855
R26939 a_n18960_7900.t19 a_n18960_7900.t6 7.92855
R26940 a_n18960_7900.t8 a_n18960_7900.t14 5.96436
R26941 a_n18960_7900.t17 a_n18960_7900.t13 5.96436
R26942 a_n18960_7900.t15 a_n18960_7900.t9 5.96436
R26943 a_n18960_7900.t16 a_n18960_7900.t12 5.96436
R26944 a_n18960_7900.n3 a_n18960_7900.n2 3.08997
R26945 a_n18960_7900.n1 a_n18960_7900.n0 3.08997
R26946 a_n18960_7900.n13 a_n18960_7900.n3 5.46561
R26947 a_n18960_7900.n12 a_n18960_7900.n6 5.46561
R26948 a_n18960_7900.n17 a_n18960_7900.n20 40.691
R26949 a_n18960_7900.n23 a_n18960_7900.n18 37.3469
R26950 a_n18960_7900.n19 a_n18960_7900.n23 24.5212
R26951 a_n18960_7900.n14 a_n18960_7900.n17 15.0268
R26952 a_n18960_7900.n14 a_n18960_7900.n13 11.078
R26953 a_n6364_n172.n101 a_n6364_n172.n99 289.615
R26954 a_n6364_n172.n57 a_n6364_n172.n55 289.615
R26955 a_n6364_n172.n61 a_n6364_n172.n10 214.716
R26956 a_n6364_n172.n67 a_n6364_n172.n12 214.716
R26957 a_n6364_n172.n69 a_n6364_n172.n14 214.716
R26958 a_n6364_n172.n71 a_n6364_n172.n16 214.716
R26959 a_n6364_n172.n73 a_n6364_n172.n18 214.716
R26960 a_n6364_n172.n75 a_n6364_n172.n20 214.716
R26961 a_n6364_n172.n93 a_n6364_n172.n91 289.615
R26962 a_n6364_n172.n84 a_n6364_n172.n82 289.615
R26963 a_n6364_n172.n4 a_n6364_n172.n62 197.849
R26964 a_n6364_n172.n4 a_n6364_n172.n68 197.849
R26965 a_n6364_n172.n2 a_n6364_n172.n70 197.849
R26966 a_n6364_n172.n2 a_n6364_n172.n72 197.849
R26967 a_n6364_n172.n3 a_n6364_n172.n74 197.849
R26968 a_n6364_n172.n3 a_n6364_n172.n76 197.849
R26969 a_n6364_n172.n102 a_n6364_n172.n101 185
R26970 a_n6364_n172.n100 a_n6364_n172.n6 185
R26971 a_n6364_n172.n26 a_n6364_n172.n25 185
R26972 a_n6364_n172.n58 a_n6364_n172.n57 185
R26973 a_n6364_n172.n56 a_n6364_n172.n8 185
R26974 a_n6364_n172.n29 a_n6364_n172.n28 185
R26975 a_n6364_n172.n9 a_n6364_n172.n10 4.57211
R26976 a_n6364_n172.n61 a_n6364_n172.n31 185
R26977 a_n6364_n172.n11 a_n6364_n172.n12 4.57211
R26978 a_n6364_n172.n67 a_n6364_n172.n33 185
R26979 a_n6364_n172.n13 a_n6364_n172.n14 4.57211
R26980 a_n6364_n172.n69 a_n6364_n172.n35 185
R26981 a_n6364_n172.n15 a_n6364_n172.n16 4.57211
R26982 a_n6364_n172.n71 a_n6364_n172.n37 185
R26983 a_n6364_n172.n17 a_n6364_n172.n18 4.57211
R26984 a_n6364_n172.n73 a_n6364_n172.n39 185
R26985 a_n6364_n172.n19 a_n6364_n172.n20 4.57211
R26986 a_n6364_n172.n75 a_n6364_n172.n41 185
R26987 a_n6364_n172.n44 a_n6364_n172.n43 185
R26988 a_n6364_n172.n92 a_n6364_n172.n22 185
R26989 a_n6364_n172.n94 a_n6364_n172.n93 185
R26990 a_n6364_n172.n47 a_n6364_n172.n46 185
R26991 a_n6364_n172.n83 a_n6364_n172.n24 185
R26992 a_n6364_n172.n85 a_n6364_n172.n84 185
R26993 a_n6364_n172.n32 a_n6364_n172.t11 154.111
R26994 a_n6364_n172.n34 a_n6364_n172.t0 154.111
R26995 a_n6364_n172.n36 a_n6364_n172.t8 154.111
R26996 a_n6364_n172.n38 a_n6364_n172.t2 154.111
R26997 a_n6364_n172.n40 a_n6364_n172.t9 154.111
R26998 a_n6364_n172.n42 a_n6364_n172.t25 154.111
R26999 a_n6364_n172.n101 a_n6364_n172.n100 104.615
R27000 a_n6364_n172.n100 a_n6364_n172.n25 104.615
R27001 a_n6364_n172.n57 a_n6364_n172.n56 104.615
R27002 a_n6364_n172.n56 a_n6364_n172.n28 104.615
R27003 a_n6364_n172.n92 a_n6364_n172.n43 104.615
R27004 a_n6364_n172.n93 a_n6364_n172.n92 104.615
R27005 a_n6364_n172.n83 a_n6364_n172.n46 104.615
R27006 a_n6364_n172.n84 a_n6364_n172.n83 104.615
R27007 a_n6364_n172.n107 a_n6364_n172.n106 70.5734
R27008 a_n6364_n172.n64 a_n6364_n172.n63 70.5734
R27009 a_n6364_n172.n66 a_n6364_n172.n65 70.5734
R27010 a_n6364_n172.n108 a_n6364_n172.n1 70.5734
R27011 a_n6364_n172.n90 a_n6364_n172.n89 70.5733
R27012 a_n6364_n172.n0 a_n6364_n172.n88 70.5733
R27013 a_n6364_n172.n81 a_n6364_n172.n80 70.5733
R27014 a_n6364_n172.n79 a_n6364_n172.n78 70.5733
R27015 a_n6364_n172.t16 a_n6364_n172.n25 52.3082
R27016 a_n6364_n172.t10 a_n6364_n172.n28 52.3082
R27017 a_n6364_n172.n61 a_n6364_n172.t11 52.3082
R27018 a_n6364_n172.n67 a_n6364_n172.t0 52.3082
R27019 a_n6364_n172.n69 a_n6364_n172.t8 52.3082
R27020 a_n6364_n172.n71 a_n6364_n172.t2 52.3082
R27021 a_n6364_n172.n73 a_n6364_n172.t9 52.3082
R27022 a_n6364_n172.n75 a_n6364_n172.t25 52.3082
R27023 a_n6364_n172.t23 a_n6364_n172.n43 52.3082
R27024 a_n6364_n172.t15 a_n6364_n172.n46 52.3082
R27025 a_n6364_n172.n105 a_n6364_n172.n104 41.6884
R27026 a_n6364_n172.n1 a_n6364_n172.n60 41.6884
R27027 a_n6364_n172.n97 a_n6364_n172.n96 41.6884
R27028 a_n6364_n172.n0 a_n6364_n172.n87 41.6884
R27029 a_n6364_n172.n27 a_n6364_n172.n26 5.02765
R27030 a_n6364_n172.n30 a_n6364_n172.n29 5.02765
R27031 a_n6364_n172.n45 a_n6364_n172.n44 5.02765
R27032 a_n6364_n172.n48 a_n6364_n172.n47 5.02765
R27033 a_n6364_n172.n31 a_n6364_n172.n32 4.9836
R27034 a_n6364_n172.n33 a_n6364_n172.n34 4.9836
R27035 a_n6364_n172.n35 a_n6364_n172.n36 4.9836
R27036 a_n6364_n172.n37 a_n6364_n172.n38 4.9836
R27037 a_n6364_n172.n39 a_n6364_n172.n40 4.9836
R27038 a_n6364_n172.n41 a_n6364_n172.n42 4.9836
R27039 a_n6364_n172.n6 a_n6364_n172.n26 12.8005
R27040 a_n6364_n172.n8 a_n6364_n172.n29 12.8005
R27041 a_n6364_n172.n9 a_n6364_n172.n31 12.8005
R27042 a_n6364_n172.n11 a_n6364_n172.n33 12.8005
R27043 a_n6364_n172.n13 a_n6364_n172.n35 12.8005
R27044 a_n6364_n172.n15 a_n6364_n172.n37 12.8005
R27045 a_n6364_n172.n17 a_n6364_n172.n39 12.8005
R27046 a_n6364_n172.n19 a_n6364_n172.n41 12.8005
R27047 a_n6364_n172.n22 a_n6364_n172.n44 12.8005
R27048 a_n6364_n172.n24 a_n6364_n172.n47 12.8005
R27049 a_n6364_n172.n102 a_n6364_n172.n6 12.0247
R27050 a_n6364_n172.n58 a_n6364_n172.n8 12.0247
R27051 a_n6364_n172.n94 a_n6364_n172.n22 12.0247
R27052 a_n6364_n172.n85 a_n6364_n172.n24 12.0247
R27053 a_n6364_n172.n77 a_n6364_n172.n66 11.8654
R27054 a_n6364_n172.n103 a_n6364_n172.n99 11.249
R27055 a_n6364_n172.n59 a_n6364_n172.n55 11.249
R27056 a_n6364_n172.n95 a_n6364_n172.n91 11.249
R27057 a_n6364_n172.n86 a_n6364_n172.n82 11.249
R27058 a_n6364_n172.n105 a_n6364_n172.n98 10.5271
R27059 a_n6364_n172.n48 a_n6364_n172.n23 1.5398
R27060 a_n6364_n172.n104 a_n6364_n172.n5 9.45567
R27061 a_n6364_n172.n60 a_n6364_n172.n7 9.45567
R27062 a_n6364_n172.n62 a_n6364_n172.n49 9.45567
R27063 a_n6364_n172.n68 a_n6364_n172.n50 9.45567
R27064 a_n6364_n172.n70 a_n6364_n172.n51 9.45567
R27065 a_n6364_n172.n72 a_n6364_n172.n52 9.45567
R27066 a_n6364_n172.n74 a_n6364_n172.n53 9.45567
R27067 a_n6364_n172.n76 a_n6364_n172.n54 9.45567
R27068 a_n6364_n172.n96 a_n6364_n172.n21 9.45567
R27069 a_n6364_n172.n87 a_n6364_n172.n23 9.45567
R27070 a_n6364_n172.n5 a_n6364_n172.n103 9.3005
R27071 a_n6364_n172.n7 a_n6364_n172.n59 9.3005
R27072 a_n6364_n172.n21 a_n6364_n172.n95 9.3005
R27073 a_n6364_n172.n23 a_n6364_n172.n86 9.3005
R27074 a_n6364_n172.n79 a_n6364_n172.n77 7.57378
R27075 a_n6364_n172.n98 a_n6364_n172.n97 6.23541
R27076 a_n6364_n172.n106 a_n6364_n172.t14 5.96436
R27077 a_n6364_n172.n106 a_n6364_n172.t13 5.96436
R27078 a_n6364_n172.n63 a_n6364_n172.t7 5.96436
R27079 a_n6364_n172.n63 a_n6364_n172.t3 5.96436
R27080 a_n6364_n172.n65 a_n6364_n172.t4 5.96436
R27081 a_n6364_n172.n65 a_n6364_n172.t12 5.96436
R27082 a_n6364_n172.n89 a_n6364_n172.t6 5.96436
R27083 a_n6364_n172.n89 a_n6364_n172.t5 5.96436
R27084 a_n6364_n172.n88 a_n6364_n172.t24 5.96436
R27085 a_n6364_n172.n88 a_n6364_n172.t1 5.96436
R27086 a_n6364_n172.n80 a_n6364_n172.t17 5.96436
R27087 a_n6364_n172.n80 a_n6364_n172.t21 5.96436
R27088 a_n6364_n172.n78 a_n6364_n172.t19 5.96436
R27089 a_n6364_n172.n78 a_n6364_n172.t20 5.96436
R27090 a_n6364_n172.n108 a_n6364_n172.t18 5.96436
R27091 a_n6364_n172.t22 a_n6364_n172.n108 5.96436
R27092 a_n6364_n172.n27 a_n6364_n172.t16 151.083
R27093 a_n6364_n172.n30 a_n6364_n172.t10 151.083
R27094 a_n6364_n172.n45 a_n6364_n172.t23 151.083
R27095 a_n6364_n172.n48 a_n6364_n172.t15 151.083
R27096 a_n6364_n172.n24 a_n6364_n172.n23 10.4641
R27097 a_n6364_n172.n22 a_n6364_n172.n21 10.4641
R27098 a_n6364_n172.n54 a_n6364_n172.n19 10.4641
R27099 a_n6364_n172.n53 a_n6364_n172.n17 10.4641
R27100 a_n6364_n172.n52 a_n6364_n172.n15 10.4641
R27101 a_n6364_n172.n51 a_n6364_n172.n13 10.4641
R27102 a_n6364_n172.n50 a_n6364_n172.n11 10.4641
R27103 a_n6364_n172.n49 a_n6364_n172.n9 10.4641
R27104 a_n6364_n172.n8 a_n6364_n172.n7 10.4641
R27105 a_n6364_n172.n6 a_n6364_n172.n5 10.4641
R27106 a_n6364_n172.n27 a_n6364_n172.n5 1.5398
R27107 a_n6364_n172.n30 a_n6364_n172.n7 1.5398
R27108 a_n6364_n172.n32 a_n6364_n172.n49 1.57128
R27109 a_n6364_n172.n34 a_n6364_n172.n50 1.57128
R27110 a_n6364_n172.n36 a_n6364_n172.n51 1.57128
R27111 a_n6364_n172.n38 a_n6364_n172.n52 1.57128
R27112 a_n6364_n172.n40 a_n6364_n172.n53 1.57128
R27113 a_n6364_n172.n42 a_n6364_n172.n54 1.57128
R27114 a_n6364_n172.n45 a_n6364_n172.n21 1.5398
R27115 a_n6364_n172.n98 a_n6364_n172.n4 4.69967
R27116 a_n6364_n172.n77 a_n6364_n172.n3 3.36973
R27117 a_n6364_n172.n104 a_n6364_n172.n99 2.71565
R27118 a_n6364_n172.n60 a_n6364_n172.n55 2.71565
R27119 a_n6364_n172.n96 a_n6364_n172.n91 2.71565
R27120 a_n6364_n172.n87 a_n6364_n172.n82 2.71565
R27121 a_n6364_n172.n81 a_n6364_n172.n79 2.67722
R27122 a_n6364_n172.n0 a_n6364_n172.n81 2.67722
R27123 a_n6364_n172.n97 a_n6364_n172.n90 2.67722
R27124 a_n6364_n172.n66 a_n6364_n172.n64 2.67722
R27125 a_n6364_n172.n64 a_n6364_n172.n1 2.67722
R27126 a_n6364_n172.n107 a_n6364_n172.n105 2.67722
R27127 a_n6364_n172.n103 a_n6364_n172.n102 1.93989
R27128 a_n6364_n172.n59 a_n6364_n172.n58 1.93989
R27129 a_n6364_n172.n62 a_n6364_n172.n10 9.09642
R27130 a_n6364_n172.n68 a_n6364_n172.n12 9.09642
R27131 a_n6364_n172.n70 a_n6364_n172.n14 9.09642
R27132 a_n6364_n172.n72 a_n6364_n172.n16 9.09642
R27133 a_n6364_n172.n74 a_n6364_n172.n18 9.09642
R27134 a_n6364_n172.n76 a_n6364_n172.n20 9.09642
R27135 a_n6364_n172.n3 a_n6364_n172.n2 4.42201
R27136 a_n6364_n172.n1 a_n6364_n172.n107 4.2505
R27137 a_n6364_n172.n90 a_n6364_n172.n0 4.2505
R27138 a_n6364_n172.n2 a_n6364_n172.n4 2.94817
R27139 a_n6364_n172.n95 a_n6364_n172.n94 1.93989
R27140 a_n6364_n172.n86 a_n6364_n172.n85 1.93989
R27141 a_n7651_8750.n38 a_n7651_8750.n17 214.892
R27142 a_n7651_8750.n38 a_n7651_8750.n25 185
R27143 a_n7651_8750.n30 a_n7651_8750.n29 185
R27144 a_n7651_8750.n33 a_n7651_8750.n32 185
R27145 a_n7651_8750.n36 a_n7651_8750.n27 185
R27146 a_n7651_8750.n20 a_n7651_8750.n21 8.29153
R27147 a_n7651_8750.n24 a_n7651_8750.n7 4.69023
R27148 a_n7651_8750.n10 a_n7651_8750.t17 105.144
R27149 a_n7651_8750.n38 a_n7651_8750.n29 104.615
R27150 a_n7651_8750.n36 a_n7651_8750.n32 104.615
R27151 a_n7651_8750.n21 a_n7651_8750.n36 214.892
R27152 a_n7651_8750.n23 a_n7651_8750.t15 103.32
R27153 a_n7651_8750.n15 a_n7651_8750.t1 100.508
R27154 a_n7651_8750.n28 a_n7651_8750.t3 100.508
R27155 a_n7651_8750.n15 a_n7651_8750.t7 98.5007
R27156 a_n7651_8750.n28 a_n7651_8750.t0 98.5006
R27157 a_n7651_8750.n23 a_n7651_8750.t21 97.216
R27158 a_n7651_8750.n10 a_n7651_8750.t25 95.3927
R27159 a_n7651_8750.n10 a_n7651_8750.t19 95.3927
R27160 a_n7651_8750.t27 a_n7651_8750.n23 95.3926
R27161 a_n7651_8750.n28 a_n7651_8750.n37 72.2924
R27162 a_n7651_8750.n15 a_n7651_8750.n17 69.6157
R27163 a_n7651_8750.t2 a_n7651_8750.n29 52.3082
R27164 a_n7651_8750.t9 a_n7651_8750.n32 52.3082
R27165 a_n7651_8750.n3 a_n7651_8750.n4 1.82316
R27166 a_n7651_8750.n0 a_n7651_8750.n1 1.82316
R27167 a_n7651_8750.n9 a_n7651_8750.t36 56.9465
R27168 a_n7651_8750.n9 a_n7651_8750.t45 54.7818
R27169 a_n7651_8750.n9 a_n7651_8750.t35 58.6647
R27170 a_n7651_8750.n9 a_n7651_8750.t34 57.8307
R27171 a_n7651_8750.n11 a_n7651_8750.t31 62.4753
R27172 a_n7651_8750.n11 a_n7651_8750.t47 54.1629
R27173 a_n7651_8750.n9 a_n7651_8750.t30 55.0537
R27174 a_n7651_8750.n9 a_n7651_8750.t46 57.8307
R27175 a_n7651_8750.n9 a_n7651_8750.t49 56.9465
R27176 a_n7651_8750.n18 a_n7651_8750.t52 54.3195
R27177 a_n7651_8750.n18 a_n7651_8750.t40 60.2658
R27178 a_n7651_8750.n9 a_n7651_8750.t53 57.8307
R27179 a_n7651_8750.n13 a_n7651_8750.t55 62.4469
R27180 a_n7651_8750.n13 a_n7651_8750.t39 54.1784
R27181 a_n7651_8750.n9 a_n7651_8750.t48 55.0537
R27182 a_n7651_8750.n9 a_n7651_8750.t32 57.8307
R27183 a_n7651_8750.n19 a_n7651_8750.t54 52.9495
R27184 a_n7651_8750.n14 a_n7651_8750.t44 60.3423
R27185 a_n7651_8750.n14 a_n7651_8750.t43 55.3078
R27186 a_n7651_8750.n19 a_n7651_8750.t42 60.8968
R27187 a_n7651_8750.n6 a_n7651_8750.t33 56.6979
R27188 a_n7651_8750.n39 a_n7651_8750.t24 25.3364
R27189 a_n7651_8750.n7 a_n7651_8750.t18 56.6979
R27190 a_n7651_8750.n8 a_n7651_8750.t28 55.9038
R27191 a_n7651_8750.n35 a_n7651_8750.t12 25.3364
R27192 a_n7651_8750.n22 a_n7651_8750.t16 56.6979
R27193 a_n7651_8750.n5 a_n7651_8750.t26 52.6435
R27194 a_n7651_8750.n4 a_n7651_8750.t20 59.4248
R27195 a_n7651_8750.n4 a_n7651_8750.t22 55.61
R27196 a_n7651_8750.n5 a_n7651_8750.t10 61.6702
R27197 a_n7651_8750.n3 a_n7651_8750.t14 56.6979
R27198 a_n7651_8750.n2 a_n7651_8750.t41 52.6435
R27199 a_n7651_8750.n1 a_n7651_8750.t38 59.4248
R27200 a_n7651_8750.n1 a_n7651_8750.t51 55.61
R27201 a_n7651_8750.n2 a_n7651_8750.t37 61.6702
R27202 a_n7651_8750.n0 a_n7651_8750.t50 56.6979
R27203 a_n7651_8750.n6 a_n7651_8750.n19 3.75241
R27204 a_n7651_8750.n7 a_n7651_8750.n8 1.58003
R27205 a_n7651_8750.n8 a_n7651_8750.n39 50.9422
R27206 a_n7651_8750.n39 a_n7651_8750.n24 73.3549
R27207 a_n7651_8750.n24 a_n7651_8750.n35 59.7493
R27208 a_n7651_8750.n35 a_n7651_8750.n22 64.2385
R27209 a_n7651_8750.n5 a_n7651_8750.n3 4.25859
R27210 a_n7651_8750.n2 a_n7651_8750.n0 4.25859
R27211 a_n7651_8750.n31 a_n7651_8750.n30 5.02765
R27212 a_n7651_8750.n34 a_n7651_8750.n33 5.02765
R27213 a_n7651_8750.n0 a_n7651_8750.n9 14.171
R27214 a_n7651_8750.n6 a_n7651_8750.n12 13.9665
R27215 a_n7651_8750.n25 a_n7651_8750.n30 12.8005
R27216 a_n7651_8750.n27 a_n7651_8750.n33 12.8005
R27217 a_n7651_8750.n9 a_n7651_8750.n7 12.6616
R27218 a_n7651_8750.n14 a_n7651_8750.n6 2.27518
R27219 a_n7651_8750.n21 a_n7651_8750.n37 9.42119
R27220 a_n7651_8750.n12 a_n7651_8750.n3 10.6824
R27221 a_n7651_8750.n17 a_n7651_8750.n16 5.46409
R27222 a_n7651_8750.n37 a_n7651_8750.n26 9.45567
R27223 a_n7651_8750.t21 a_n7651_8750.t23 7.92855
R27224 a_n7651_8750.t25 a_n7651_8750.t13 7.92855
R27225 a_n7651_8750.t19 a_n7651_8750.t29 7.92855
R27226 a_n7651_8750.t11 a_n7651_8750.t27 7.92855
R27227 a_n7651_8750.n7 a_n7651_8750.n6 7.27718
R27228 a_n7651_8750.n3 a_n7651_8750.n0 7.27718
R27229 a_n7651_8750.n34 a_n7651_8750.n26 1.5398
R27230 a_n7651_8750.t1 a_n7651_8750.t6 5.96436
R27231 a_n7651_8750.t7 a_n7651_8750.t5 5.96436
R27232 a_n7651_8750.t3 a_n7651_8750.t8 5.96436
R27233 a_n7651_8750.t0 a_n7651_8750.t4 5.96436
R27234 a_n7651_8750.n31 a_n7651_8750.t2 151.083
R27235 a_n7651_8750.n34 a_n7651_8750.t9 151.083
R27236 a_n7651_8750.n15 a_n7651_8750.n28 38.614
R27237 a_n7651_8750.n7 a_n7651_8750.n15 27.2531
R27238 a_n7651_8750.n11 a_n7651_8750.n9 14.4697
R27239 a_n7651_8750.n13 a_n7651_8750.n9 13.9709
R27240 a_n7651_8750.n9 a_n7651_8750.n18 12.2318
R27241 a_n7651_8750.n23 a_n7651_8750.n12 11.5202
R27242 a_n7651_8750.n22 a_n7651_8750.n7 10.9964
R27243 a_n7651_8750.n9 a_n7651_8750.n12 10.6307
R27244 a_n7651_8750.n31 a_n7651_8750.n16 2.61599
R27245 a_n7651_8750.n26 a_n7651_8750.n20 3.48794
R27246 a_n7651_8750.n27 a_n7651_8750.n20 3.73143
R27247 a_n7651_8750.n25 a_n7651_8750.n16 5.74693
R27248 a_n7651_8750.n9 a_n7651_8750.n10 10.4445
R27249 a_n7729_8946.n4 a_n7729_8946.t0 133.071
R27250 a_n7729_8946.n0 a_n7729_8946.t6 131.993
R27251 a_n7729_8946.n0 a_n7729_8946.n2 123.32
R27252 a_n7729_8946.n4 a_n7729_8946.n3 123.32
R27253 a_n7729_8946.n13 a_n7729_8946.n0 123.32
R27254 a_n7729_8946.n6 a_n7729_8946.n5 123.32
R27255 a_n7729_8946.n8 a_n7729_8946.t16 105.144
R27256 a_n7729_8946.n11 a_n7729_8946.t15 103.32
R27257 a_n7729_8946.n1 a_n7729_8946.t13 103.32
R27258 a_n7729_8946.n1 a_n7729_8946.t11 103.32
R27259 a_n7729_8946.n10 a_n7729_8946.n9 95.3927
R27260 a_n7729_8946.n8 a_n7729_8946.n7 95.3927
R27261 a_n7729_8946.n0 a_n7729_8946.n12 19.7595
R27262 a_n7729_8946.n12 a_n7729_8946.n6 12.5046
R27263 a_n7729_8946.n2 a_n7729_8946.t3 7.92855
R27264 a_n7729_8946.n2 a_n7729_8946.t1 7.92855
R27265 a_n7729_8946.n5 a_n7729_8946.t8 7.92855
R27266 a_n7729_8946.n5 a_n7729_8946.t4 7.92855
R27267 a_n7729_8946.n3 a_n7729_8946.t7 7.92855
R27268 a_n7729_8946.n3 a_n7729_8946.t2 7.92855
R27269 a_n7729_8946.n9 a_n7729_8946.t12 7.92855
R27270 a_n7729_8946.n9 a_n7729_8946.t14 7.92855
R27271 a_n7729_8946.n7 a_n7729_8946.t10 7.92855
R27272 a_n7729_8946.n7 a_n7729_8946.t17 7.92855
R27273 a_n7729_8946.t9 a_n7729_8946.n13 7.92855
R27274 a_n7729_8946.n13 a_n7729_8946.t5 7.92855
R27275 a_n7729_8946.n12 a_n7729_8946.n11 5.91753
R27276 a_n7729_8946.n10 a_n7729_8946.n1 2.28929
R27277 a_n7729_8946.n6 a_n7729_8946.n4 1.82378
R27278 a_n7729_8946.n1 a_n7729_8946.n8 1.82378
R27279 a_n7729_8946.n11 a_n7729_8946.n10 1.82378
R27280 VP.n162 VP.t0 243.255
R27281 VP.n161 VP.n159 224.169
R27282 VP.n161 VP.n160 223.454
R27283 VP.n100 VP.n97 161.3
R27284 VP.n102 VP.n101 161.3
R27285 VP.n103 VP.n96 161.3
R27286 VP.n105 VP.n104 161.3
R27287 VP.n106 VP.n95 161.3
R27288 VP.n108 VP.n107 161.3
R27289 VP.n109 VP.n94 161.3
R27290 VP.n111 VP.n110 161.3
R27291 VP.n112 VP.n93 161.3
R27292 VP.n114 VP.n113 161.3
R27293 VP.n115 VP.n92 161.3
R27294 VP.n117 VP.n116 161.3
R27295 VP.n118 VP.n91 161.3
R27296 VP.n120 VP.n119 161.3
R27297 VP.n121 VP.n90 161.3
R27298 VP.n123 VP.n122 161.3
R27299 VP.n124 VP.n89 161.3
R27300 VP.n126 VP.n125 161.3
R27301 VP.n127 VP.n88 161.3
R27302 VP.n129 VP.n128 161.3
R27303 VP.n130 VP.n87 161.3
R27304 VP.n132 VP.n131 161.3
R27305 VP.n133 VP.n86 161.3
R27306 VP.n135 VP.n134 161.3
R27307 VP.n136 VP.n85 161.3
R27308 VP.n139 VP.n138 161.3
R27309 VP.n140 VP.n84 161.3
R27310 VP.n142 VP.n141 161.3
R27311 VP.n143 VP.n83 161.3
R27312 VP.n145 VP.n144 161.3
R27313 VP.n146 VP.n82 161.3
R27314 VP.n148 VP.n147 161.3
R27315 VP.n149 VP.n81 161.3
R27316 VP.n151 VP.n150 161.3
R27317 VP.n152 VP.n80 161.3
R27318 VP.n154 VP.n153 161.3
R27319 VP.n155 VP.n79 161.3
R27320 VP.n76 VP.n0 161.3
R27321 VP.n75 VP.n74 161.3
R27322 VP.n73 VP.n1 161.3
R27323 VP.n72 VP.n71 161.3
R27324 VP.n70 VP.n2 161.3
R27325 VP.n69 VP.n68 161.3
R27326 VP.n67 VP.n3 161.3
R27327 VP.n66 VP.n65 161.3
R27328 VP.n64 VP.n4 161.3
R27329 VP.n63 VP.n62 161.3
R27330 VP.n61 VP.n5 161.3
R27331 VP.n60 VP.n59 161.3
R27332 VP.n57 VP.n6 161.3
R27333 VP.n56 VP.n55 161.3
R27334 VP.n54 VP.n7 161.3
R27335 VP.n53 VP.n52 161.3
R27336 VP.n51 VP.n8 161.3
R27337 VP.n50 VP.n49 161.3
R27338 VP.n48 VP.n9 161.3
R27339 VP.n47 VP.n46 161.3
R27340 VP.n45 VP.n10 161.3
R27341 VP.n44 VP.n43 161.3
R27342 VP.n42 VP.n11 161.3
R27343 VP.n41 VP.n40 161.3
R27344 VP.n39 VP.n12 161.3
R27345 VP.n38 VP.n37 161.3
R27346 VP.n36 VP.n13 161.3
R27347 VP.n35 VP.n34 161.3
R27348 VP.n33 VP.n14 161.3
R27349 VP.n32 VP.n31 161.3
R27350 VP.n30 VP.n15 161.3
R27351 VP.n29 VP.n28 161.3
R27352 VP.n27 VP.n16 161.3
R27353 VP.n26 VP.n25 161.3
R27354 VP.n24 VP.n17 161.3
R27355 VP.n23 VP.n22 161.3
R27356 VP.n21 VP.n18 161.3
R27357 VP.n99 VP.n98 65.7373
R27358 VP.n20 VP.n19 65.7373
R27359 VP.n157 VP.n156 56.8746
R27360 VP.n78 VP.n77 56.8746
R27361 VP.n148 VP.n82 56.5617
R27362 VP.n69 VP.n3 56.5617
R27363 VP.n158 VP.n157 52.6226
R27364 VP.n129 VP.n88 50.7491
R27365 VP.n107 VP.n94 50.7491
R27366 VP.n28 VP.n15 50.7491
R27367 VP.n50 VP.n9 50.7491
R27368 VP.n19 VP.t8 46.6743
R27369 VP.n98 VP.t11 46.6739
R27370 VP.n125 VP.n88 30.405
R27371 VP.n111 VP.n94 30.405
R27372 VP.n32 VP.n15 30.405
R27373 VP.n46 VP.n9 30.405
R27374 VP.n155 VP.n154 24.5923
R27375 VP.n154 VP.n80 24.5923
R27376 VP.n150 VP.n80 24.5923
R27377 VP.n150 VP.n149 24.5923
R27378 VP.n149 VP.n148 24.5923
R27379 VP.n144 VP.n82 24.5923
R27380 VP.n144 VP.n143 24.5923
R27381 VP.n143 VP.n142 24.5923
R27382 VP.n142 VP.n84 24.5923
R27383 VP.n138 VP.n84 24.5923
R27384 VP.n136 VP.n135 24.5923
R27385 VP.n135 VP.n86 24.5923
R27386 VP.n131 VP.n86 24.5923
R27387 VP.n131 VP.n130 24.5923
R27388 VP.n130 VP.n129 24.5923
R27389 VP.n125 VP.n124 24.5923
R27390 VP.n124 VP.n123 24.5923
R27391 VP.n123 VP.n90 24.5923
R27392 VP.n119 VP.n90 24.5923
R27393 VP.n119 VP.n118 24.5923
R27394 VP.n118 VP.n117 24.5923
R27395 VP.n117 VP.n92 24.5923
R27396 VP.n113 VP.n92 24.5923
R27397 VP.n113 VP.n112 24.5923
R27398 VP.n112 VP.n111 24.5923
R27399 VP.n107 VP.n106 24.5923
R27400 VP.n106 VP.n105 24.5923
R27401 VP.n105 VP.n96 24.5923
R27402 VP.n101 VP.n96 24.5923
R27403 VP.n101 VP.n100 24.5923
R27404 VP.n22 VP.n21 24.5923
R27405 VP.n22 VP.n17 24.5923
R27406 VP.n26 VP.n17 24.5923
R27407 VP.n27 VP.n26 24.5923
R27408 VP.n28 VP.n27 24.5923
R27409 VP.n33 VP.n32 24.5923
R27410 VP.n34 VP.n33 24.5923
R27411 VP.n34 VP.n13 24.5923
R27412 VP.n38 VP.n13 24.5923
R27413 VP.n39 VP.n38 24.5923
R27414 VP.n40 VP.n39 24.5923
R27415 VP.n40 VP.n11 24.5923
R27416 VP.n44 VP.n11 24.5923
R27417 VP.n45 VP.n44 24.5923
R27418 VP.n46 VP.n45 24.5923
R27419 VP.n51 VP.n50 24.5923
R27420 VP.n52 VP.n51 24.5923
R27421 VP.n52 VP.n7 24.5923
R27422 VP.n56 VP.n7 24.5923
R27423 VP.n57 VP.n56 24.5923
R27424 VP.n59 VP.n5 24.5923
R27425 VP.n63 VP.n5 24.5923
R27426 VP.n64 VP.n63 24.5923
R27427 VP.n65 VP.n64 24.5923
R27428 VP.n65 VP.n3 24.5923
R27429 VP.n70 VP.n69 24.5923
R27430 VP.n71 VP.n70 24.5923
R27431 VP.n71 VP.n1 24.5923
R27432 VP.n75 VP.n1 24.5923
R27433 VP.n76 VP.n75 24.5923
R27434 VP.n156 VP.n155 20.6576
R27435 VP.n77 VP.n76 20.6576
R27436 VP.n160 VP.t2 19.8005
R27437 VP.n160 VP.t4 19.8005
R27438 VP.n159 VP.t1 19.8005
R27439 VP.n159 VP.t3 19.8005
R27440 VP.n138 VP.n137 14.2638
R27441 VP.n59 VP.n58 14.2638
R27442 VP.n118 VP.t9 13.608
R27443 VP.n156 VP.t7 13.608
R27444 VP.n137 VP.t6 13.608
R27445 VP.n99 VP.t14 13.608
R27446 VP.n39 VP.t12 13.608
R27447 VP.n20 VP.t5 13.608
R27448 VP.n58 VP.t13 13.608
R27449 VP.n77 VP.t10 13.608
R27450 VP.n158 VP.n78 13.24
R27451 VP VP.n163 13.209
R27452 VP.n137 VP.n136 10.3291
R27453 VP.n100 VP.n99 10.3291
R27454 VP.n21 VP.n20 10.3291
R27455 VP.n58 VP.n57 10.3291
R27456 VP.n163 VP.n162 4.80222
R27457 VP.n19 VP.n18 0.993426
R27458 VP.n98 VP.n97 0.993421
R27459 VP.n163 VP.n158 0.972091
R27460 VP.n162 VP.n161 0.716017
R27461 VP.n157 VP.n79 0.502096
R27462 VP.n78 VP.n0 0.502096
R27463 VP.n153 VP.n79 0.189894
R27464 VP.n153 VP.n152 0.189894
R27465 VP.n152 VP.n151 0.189894
R27466 VP.n151 VP.n81 0.189894
R27467 VP.n147 VP.n81 0.189894
R27468 VP.n147 VP.n146 0.189894
R27469 VP.n146 VP.n145 0.189894
R27470 VP.n145 VP.n83 0.189894
R27471 VP.n141 VP.n83 0.189894
R27472 VP.n141 VP.n140 0.189894
R27473 VP.n140 VP.n139 0.189894
R27474 VP.n139 VP.n85 0.189894
R27475 VP.n134 VP.n85 0.189894
R27476 VP.n134 VP.n133 0.189894
R27477 VP.n133 VP.n132 0.189894
R27478 VP.n132 VP.n87 0.189894
R27479 VP.n128 VP.n87 0.189894
R27480 VP.n128 VP.n127 0.189894
R27481 VP.n127 VP.n126 0.189894
R27482 VP.n126 VP.n89 0.189894
R27483 VP.n122 VP.n89 0.189894
R27484 VP.n122 VP.n121 0.189894
R27485 VP.n121 VP.n120 0.189894
R27486 VP.n120 VP.n91 0.189894
R27487 VP.n116 VP.n91 0.189894
R27488 VP.n116 VP.n115 0.189894
R27489 VP.n115 VP.n114 0.189894
R27490 VP.n114 VP.n93 0.189894
R27491 VP.n110 VP.n93 0.189894
R27492 VP.n110 VP.n109 0.189894
R27493 VP.n109 VP.n108 0.189894
R27494 VP.n108 VP.n95 0.189894
R27495 VP.n104 VP.n95 0.189894
R27496 VP.n104 VP.n103 0.189894
R27497 VP.n103 VP.n102 0.189894
R27498 VP.n102 VP.n97 0.189894
R27499 VP.n23 VP.n18 0.189894
R27500 VP.n24 VP.n23 0.189894
R27501 VP.n25 VP.n24 0.189894
R27502 VP.n25 VP.n16 0.189894
R27503 VP.n29 VP.n16 0.189894
R27504 VP.n30 VP.n29 0.189894
R27505 VP.n31 VP.n30 0.189894
R27506 VP.n31 VP.n14 0.189894
R27507 VP.n35 VP.n14 0.189894
R27508 VP.n36 VP.n35 0.189894
R27509 VP.n37 VP.n36 0.189894
R27510 VP.n37 VP.n12 0.189894
R27511 VP.n41 VP.n12 0.189894
R27512 VP.n42 VP.n41 0.189894
R27513 VP.n43 VP.n42 0.189894
R27514 VP.n43 VP.n10 0.189894
R27515 VP.n47 VP.n10 0.189894
R27516 VP.n48 VP.n47 0.189894
R27517 VP.n49 VP.n48 0.189894
R27518 VP.n49 VP.n8 0.189894
R27519 VP.n53 VP.n8 0.189894
R27520 VP.n54 VP.n53 0.189894
R27521 VP.n55 VP.n54 0.189894
R27522 VP.n55 VP.n6 0.189894
R27523 VP.n60 VP.n6 0.189894
R27524 VP.n61 VP.n60 0.189894
R27525 VP.n62 VP.n61 0.189894
R27526 VP.n62 VP.n4 0.189894
R27527 VP.n66 VP.n4 0.189894
R27528 VP.n67 VP.n66 0.189894
R27529 VP.n68 VP.n67 0.189894
R27530 VP.n68 VP.n2 0.189894
R27531 VP.n72 VP.n2 0.189894
R27532 VP.n73 VP.n72 0.189894
R27533 VP.n74 VP.n73 0.189894
R27534 VP.n74 VP.n0 0.189894
R27535 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n2 289.615
R27536 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n13 289.615
R27537 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n25 289.615
R27538 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n37 289.615
R27539 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n49 289.615
R27540 DIFFPAIR_BIAS.n67 DIFFPAIR_BIAS.n61 289.615
R27541 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 185
R27542 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 185
R27543 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n19 185
R27544 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 185
R27545 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n31 185
R27546 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n29 185
R27547 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n43 185
R27548 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n41 185
R27549 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 185
R27550 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n53 185
R27551 DIFFPAIR_BIAS.n68 DIFFPAIR_BIAS.n67 185
R27552 DIFFPAIR_BIAS.n66 DIFFPAIR_BIAS.n65 185
R27553 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t11 151.613
R27554 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.t7 151.613
R27555 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.t9 151.613
R27556 DIFFPAIR_BIAS.n40 DIFFPAIR_BIAS.t1 151.613
R27557 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.t5 151.613
R27558 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.t3 151.613
R27559 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 104.615
R27560 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n18 104.615
R27561 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n30 104.615
R27562 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 104.615
R27563 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 104.615
R27564 DIFFPAIR_BIAS.n67 DIFFPAIR_BIAS.n66 104.615
R27565 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n12 97.6986
R27566 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n23 96.2247
R27567 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n35 96.2247
R27568 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n47 96.2247
R27569 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 96.2247
R27570 DIFFPAIR_BIAS.n72 DIFFPAIR_BIAS.n71 96.2247
R27571 DIFFPAIR_BIAS.n73 DIFFPAIR_BIAS.t10 53.2764
R27572 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t16 52.6425
R27573 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.t11 52.3082
R27574 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.t7 52.3082
R27575 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.t9 52.3082
R27576 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.t1 52.3082
R27577 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.t5 52.3082
R27578 DIFFPAIR_BIAS.n66 DIFFPAIR_BIAS.t3 52.3082
R27579 DIFFPAIR_BIAS.n73 DIFFPAIR_BIAS.t6 50.3272
R27580 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.t8 50.3272
R27581 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.t0 50.3272
R27582 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.t4 50.3272
R27583 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.t2 50.3272
R27584 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.t15 49.6934
R27585 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.t12 49.6934
R27586 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.t14 49.6934
R27587 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t17 49.6934
R27588 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t13 49.6934
R27589 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 15.3979
R27590 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 15.3979
R27591 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 15.3979
R27592 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n40 15.3979
R27593 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 15.3979
R27594 DIFFPAIR_BIAS.n65 DIFFPAIR_BIAS.n64 15.3979
R27595 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n4 12.8005
R27596 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n15 12.8005
R27597 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n27 12.8005
R27598 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n39 12.8005
R27599 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n51 12.8005
R27600 DIFFPAIR_BIAS.n68 DIFFPAIR_BIAS.n63 12.8005
R27601 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n2 12.0247
R27602 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n13 12.0247
R27603 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n25 12.0247
R27604 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n37 12.0247
R27605 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n49 12.0247
R27606 DIFFPAIR_BIAS.n69 DIFFPAIR_BIAS.n61 12.0247
R27607 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 9.45567
R27608 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n22 9.45567
R27609 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n34 9.45567
R27610 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n46 9.45567
R27611 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n58 9.45567
R27612 DIFFPAIR_BIAS.n71 DIFFPAIR_BIAS.n70 9.45567
R27613 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 9.3005
R27614 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 9.3005
R27615 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n21 9.3005
R27616 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 9.3005
R27617 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n33 9.3005
R27618 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 9.3005
R27619 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 9.3005
R27620 DIFFPAIR_BIAS.n39 DIFFPAIR_BIAS.n38 9.3005
R27621 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 9.3005
R27622 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 9.3005
R27623 DIFFPAIR_BIAS.n70 DIFFPAIR_BIAS.n69 9.3005
R27624 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n62 9.3005
R27625 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n77 5.9758
R27626 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n3 4.69785
R27627 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n14 4.69785
R27628 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n26 4.69785
R27629 DIFFPAIR_BIAS.n40 DIFFPAIR_BIAS.n38 4.69785
R27630 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n50 4.69785
R27631 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.n62 4.69785
R27632 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n72 4.56792
R27633 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n78 4.53891
R27634 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n76 2.95087
R27635 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n75 2.95087
R27636 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n74 2.95087
R27637 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.n73 2.95087
R27638 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.n0 2.95081
R27639 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n79 2.95081
R27640 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n80 2.95081
R27641 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n81 2.06723
R27642 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n2 1.93989
R27643 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n13 1.93989
R27644 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n25 1.93989
R27645 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n37 1.93989
R27646 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n49 1.93989
R27647 DIFFPAIR_BIAS.n71 DIFFPAIR_BIAS.n61 1.93989
R27648 DIFFPAIR_BIAS.n72 DIFFPAIR_BIAS.n60 1.47434
R27649 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n48 1.47434
R27650 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n36 1.47434
R27651 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n24 1.47434
R27652 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 1.16414
R27653 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 1.16414
R27654 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n32 1.16414
R27655 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n44 1.16414
R27656 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 1.16414
R27657 DIFFPAIR_BIAS.n69 DIFFPAIR_BIAS.n68 1.16414
R27658 DIFFPAIR_BIAS DIFFPAIR_BIAS.n82 0.684875
R27659 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n1 0.593389
R27660 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n4 0.388379
R27661 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n15 0.388379
R27662 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n27 0.388379
R27663 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n39 0.388379
R27664 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n51 0.388379
R27665 DIFFPAIR_BIAS.n65 DIFFPAIR_BIAS.n63 0.388379
R27666 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n3 0.155672
R27667 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n14 0.155672
R27668 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n26 0.155672
R27669 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n38 0.155672
R27670 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n50 0.155672
R27671 DIFFPAIR_BIAS.n70 DIFFPAIR_BIAS.n62 0.155672
R27672 a_n5900_7192.n7 a_n5900_7192.t12 105.144
R27673 a_n5900_7192.t10 a_n5900_7192.n15 105.144
R27674 a_n5900_7192.n2 a_n5900_7192.t3 105.144
R27675 a_n5900_7192.n0 a_n5900_7192.t14 103.32
R27676 a_n5900_7192.n0 a_n5900_7192.t18 103.32
R27677 a_n5900_7192.n10 a_n5900_7192.t11 103.32
R27678 a_n5900_7192.n15 a_n5900_7192.n14 95.3927
R27679 a_n5900_7192.n13 a_n5900_7192.n12 95.3927
R27680 a_n5900_7192.n2 a_n5900_7192.n1 95.3927
R27681 a_n5900_7192.n4 a_n5900_7192.n3 95.3927
R27682 a_n5900_7192.n7 a_n5900_7192.n6 95.3927
R27683 a_n5900_7192.n9 a_n5900_7192.n8 95.3927
R27684 a_n5900_7192.n13 a_n5900_7192.n11 28.8134
R27685 a_n5900_7192.n5 a_n5900_7192.t0 13.2483
R27686 a_n5900_7192.n5 a_n5900_7192.n4 8.80007
R27687 a_n5900_7192.n14 a_n5900_7192.t1 7.92855
R27688 a_n5900_7192.n14 a_n5900_7192.t6 7.92855
R27689 a_n5900_7192.n12 a_n5900_7192.t4 7.92855
R27690 a_n5900_7192.n12 a_n5900_7192.t5 7.92855
R27691 a_n5900_7192.n1 a_n5900_7192.t7 7.92855
R27692 a_n5900_7192.n1 a_n5900_7192.t9 7.92855
R27693 a_n5900_7192.n3 a_n5900_7192.t8 7.92855
R27694 a_n5900_7192.n3 a_n5900_7192.t2 7.92855
R27695 a_n5900_7192.n6 a_n5900_7192.t13 7.92855
R27696 a_n5900_7192.n6 a_n5900_7192.t16 7.92855
R27697 a_n5900_7192.n8 a_n5900_7192.t17 7.92855
R27698 a_n5900_7192.n8 a_n5900_7192.t15 7.92855
R27699 a_n5900_7192.n11 a_n5900_7192.n10 5.91753
R27700 a_n5900_7192.n11 a_n5900_7192.n5 3.48914
R27701 a_n5900_7192.n9 a_n5900_7192.n0 2.28929
R27702 a_n5900_7192.n4 a_n5900_7192.n2 1.82378
R27703 a_n5900_7192.n10 a_n5900_7192.n9 1.82378
R27704 a_n5900_7192.n0 a_n5900_7192.n7 1.82378
R27705 a_n5900_7192.n15 a_n5900_7192.n13 1.82378
C0 VDD VOUT 47.264103f
C1 VOUT VP 4.16339f
C2 VDD VN 0.193956f
C3 a_n8793_8946# VDD 1.44682f
C4 VOUT VN 1.25539f
C5 VP VN 16.7955f
C6 VOUT CS_BIAS 24.2888f
C7 VP CS_BIAS 0.433156f
C8 VP DIFFPAIR_BIAS 9.73e-19
C9 VN CS_BIAS 0.345257f
C10 VN DIFFPAIR_BIAS 0.001338f
C11 a_7857_8946# VDD 1.44682f
C12 DIFFPAIR_BIAS GND 58.677895f
C13 CS_BIAS GND 0.164878p
C14 VN GND 61.4798f
C15 VP GND 49.324013f
C16 VOUT GND 75.79409f
C17 VDD GND 0.690436p
C18 a_7857_8946# GND 0.498415f
C19 a_n8793_8946# GND 0.498415f
C20 a_n5900_7192.n0 GND 1.44567f
C21 a_n5900_7192.t0 GND 23.523401f
C22 a_n5900_7192.t3 GND 0.393149f
C23 a_n5900_7192.t7 GND 0.050554f
C24 a_n5900_7192.t9 GND 0.050554f
C25 a_n5900_7192.n1 GND 0.271693f
C26 a_n5900_7192.n2 GND 1.59901f
C27 a_n5900_7192.t8 GND 0.050554f
C28 a_n5900_7192.t2 GND 0.050554f
C29 a_n5900_7192.n3 GND 0.271693f
C30 a_n5900_7192.n4 GND 1.91809f
C31 a_n5900_7192.n5 GND 8.619889f
C32 a_n5900_7192.t12 GND 0.39315f
C33 a_n5900_7192.t13 GND 0.050554f
C34 a_n5900_7192.t16 GND 0.050554f
C35 a_n5900_7192.n6 GND 0.271693f
C36 a_n5900_7192.n7 GND 1.59901f
C37 a_n5900_7192.t14 GND 0.382021f
C38 a_n5900_7192.t18 GND 0.382021f
C39 a_n5900_7192.t17 GND 0.050554f
C40 a_n5900_7192.t15 GND 0.050554f
C41 a_n5900_7192.n8 GND 0.271693f
C42 a_n5900_7192.n9 GND 0.96835f
C43 a_n5900_7192.t11 GND 0.382021f
C44 a_n5900_7192.n10 GND 1.1451f
C45 a_n5900_7192.n11 GND 3.21898f
C46 a_n5900_7192.t4 GND 0.050554f
C47 a_n5900_7192.t5 GND 0.050554f
C48 a_n5900_7192.n12 GND 0.271693f
C49 a_n5900_7192.n13 GND 3.30117f
C50 a_n5900_7192.t1 GND 0.050554f
C51 a_n5900_7192.t6 GND 0.050554f
C52 a_n5900_7192.n14 GND 0.271693f
C53 a_n5900_7192.n15 GND 1.59901f
C54 a_n5900_7192.t10 GND 0.39315f
C55 VP.n0 GND 0.043338f
C56 VP.t10 GND 0.920762f
C57 VP.n1 GND 0.034694f
C58 VP.n2 GND 0.018709f
C59 VP.n3 GND 0.03056f
C60 VP.n4 GND 0.018709f
C61 VP.n5 GND 0.034694f
C62 VP.n6 GND 0.018709f
C63 VP.t13 GND 0.920762f
C64 VP.n7 GND 0.034694f
C65 VP.n8 GND 0.018709f
C66 VP.n9 GND 0.017916f
C67 VP.n10 GND 0.018709f
C68 VP.n11 GND 0.034694f
C69 VP.n12 GND 0.018709f
C70 VP.t12 GND 0.920762f
C71 VP.n13 GND 0.034694f
C72 VP.n14 GND 0.018709f
C73 VP.n15 GND 0.017916f
C74 VP.n16 GND 0.018709f
C75 VP.n17 GND 0.034694f
C76 VP.n18 GND 0.233228f
C77 VP.t5 GND 0.920762f
C78 VP.t8 GND 1.3003f
C79 VP.n19 GND 0.621729f
C80 VP.n20 GND 0.432812f
C81 VP.n21 GND 0.02476f
C82 VP.n22 GND 0.034694f
C83 VP.n23 GND 0.018709f
C84 VP.n24 GND 0.018709f
C85 VP.n25 GND 0.018709f
C86 VP.n26 GND 0.034694f
C87 VP.n27 GND 0.034694f
C88 VP.n28 GND 0.033987f
C89 VP.n29 GND 0.018709f
C90 VP.n30 GND 0.018709f
C91 VP.n31 GND 0.018709f
C92 VP.n32 GND 0.037182f
C93 VP.n33 GND 0.034694f
C94 VP.n34 GND 0.034694f
C95 VP.n35 GND 0.018709f
C96 VP.n36 GND 0.018709f
C97 VP.n37 GND 0.018709f
C98 VP.n38 GND 0.034694f
C99 VP.n39 GND 0.375869f
C100 VP.n40 GND 0.034694f
C101 VP.n41 GND 0.018709f
C102 VP.n42 GND 0.018709f
C103 VP.n43 GND 0.018709f
C104 VP.n44 GND 0.034694f
C105 VP.n45 GND 0.034694f
C106 VP.n46 GND 0.037182f
C107 VP.n47 GND 0.018709f
C108 VP.n48 GND 0.018709f
C109 VP.n49 GND 0.018709f
C110 VP.n50 GND 0.033987f
C111 VP.n51 GND 0.034694f
C112 VP.n52 GND 0.034694f
C113 VP.n53 GND 0.018709f
C114 VP.n54 GND 0.018709f
C115 VP.n55 GND 0.018709f
C116 VP.n56 GND 0.034694f
C117 VP.n57 GND 0.02476f
C118 VP.n58 GND 0.358303f
C119 VP.n59 GND 0.0275f
C120 VP.n60 GND 0.018709f
C121 VP.n61 GND 0.018709f
C122 VP.n62 GND 0.018709f
C123 VP.n63 GND 0.034694f
C124 VP.n64 GND 0.034694f
C125 VP.n65 GND 0.034694f
C126 VP.n66 GND 0.018709f
C127 VP.n67 GND 0.018709f
C128 VP.n68 GND 0.018709f
C129 VP.n69 GND 0.023831f
C130 VP.n70 GND 0.034694f
C131 VP.n71 GND 0.034694f
C132 VP.n72 GND 0.018709f
C133 VP.n73 GND 0.018709f
C134 VP.n74 GND 0.018709f
C135 VP.n75 GND 0.034694f
C136 VP.n76 GND 0.031953f
C137 VP.n77 GND 0.444571f
C138 VP.n78 GND 0.434642f
C139 VP.n79 GND 0.043338f
C140 VP.t7 GND 0.920762f
C141 VP.n80 GND 0.034694f
C142 VP.n81 GND 0.018709f
C143 VP.n82 GND 0.03056f
C144 VP.n83 GND 0.018709f
C145 VP.n84 GND 0.034694f
C146 VP.n85 GND 0.018709f
C147 VP.t6 GND 0.920762f
C148 VP.n86 GND 0.034694f
C149 VP.n87 GND 0.018709f
C150 VP.n88 GND 0.017916f
C151 VP.n89 GND 0.018709f
C152 VP.n90 GND 0.034694f
C153 VP.n91 GND 0.018709f
C154 VP.t9 GND 0.920762f
C155 VP.n92 GND 0.034694f
C156 VP.n93 GND 0.018709f
C157 VP.n94 GND 0.017916f
C158 VP.n95 GND 0.018709f
C159 VP.n96 GND 0.034694f
C160 VP.n97 GND 0.233228f
C161 VP.t14 GND 0.920762f
C162 VP.t11 GND 1.3003f
C163 VP.n98 GND 0.621732f
C164 VP.n99 GND 0.432812f
C165 VP.n100 GND 0.02476f
C166 VP.n101 GND 0.034694f
C167 VP.n102 GND 0.018709f
C168 VP.n103 GND 0.018709f
C169 VP.n104 GND 0.018709f
C170 VP.n105 GND 0.034694f
C171 VP.n106 GND 0.034694f
C172 VP.n107 GND 0.033987f
C173 VP.n108 GND 0.018709f
C174 VP.n109 GND 0.018709f
C175 VP.n110 GND 0.018709f
C176 VP.n111 GND 0.037182f
C177 VP.n112 GND 0.034694f
C178 VP.n113 GND 0.034694f
C179 VP.n114 GND 0.018709f
C180 VP.n115 GND 0.018709f
C181 VP.n116 GND 0.018709f
C182 VP.n117 GND 0.034694f
C183 VP.n118 GND 0.375869f
C184 VP.n119 GND 0.034694f
C185 VP.n120 GND 0.018709f
C186 VP.n121 GND 0.018709f
C187 VP.n122 GND 0.018709f
C188 VP.n123 GND 0.034694f
C189 VP.n124 GND 0.034694f
C190 VP.n125 GND 0.037182f
C191 VP.n126 GND 0.018709f
C192 VP.n127 GND 0.018709f
C193 VP.n128 GND 0.018709f
C194 VP.n129 GND 0.033987f
C195 VP.n130 GND 0.034694f
C196 VP.n131 GND 0.034694f
C197 VP.n132 GND 0.018709f
C198 VP.n133 GND 0.018709f
C199 VP.n134 GND 0.018709f
C200 VP.n135 GND 0.034694f
C201 VP.n136 GND 0.02476f
C202 VP.n137 GND 0.358303f
C203 VP.n138 GND 0.0275f
C204 VP.n139 GND 0.018709f
C205 VP.n140 GND 0.018709f
C206 VP.n141 GND 0.018709f
C207 VP.n142 GND 0.034694f
C208 VP.n143 GND 0.034694f
C209 VP.n144 GND 0.034694f
C210 VP.n145 GND 0.018709f
C211 VP.n146 GND 0.018709f
C212 VP.n147 GND 0.018709f
C213 VP.n148 GND 0.023831f
C214 VP.n149 GND 0.034694f
C215 VP.n150 GND 0.034694f
C216 VP.n151 GND 0.018709f
C217 VP.n152 GND 0.018709f
C218 VP.n153 GND 0.018709f
C219 VP.n154 GND 0.034694f
C220 VP.n155 GND 0.031953f
C221 VP.n156 GND 0.444571f
C222 VP.n157 GND 1.33124f
C223 VP.n158 GND 1.5427f
C224 VP.t1 GND 0.005767f
C225 VP.t3 GND 0.005767f
C226 VP.n159 GND 0.018964f
C227 VP.t2 GND 0.005767f
C228 VP.t4 GND 0.005767f
C229 VP.n160 GND 0.018704f
C230 VP.n161 GND 0.159634f
C231 VP.t0 GND 0.0321f
C232 VP.n162 GND 0.087111f
C233 VP.n163 GND 1.99476f
C234 a_n7729_8946.n0 GND 14.6051f
C235 a_n7729_8946.n1 GND 2.52994f
C236 a_n7729_8946.t5 GND 0.088471f
C237 a_n7729_8946.t6 GND 0.787261f
C238 a_n7729_8946.t3 GND 0.088471f
C239 a_n7729_8946.t1 GND 0.088471f
C240 a_n7729_8946.n2 GND 0.578656f
C241 a_n7729_8946.t0 GND 0.790526f
C242 a_n7729_8946.t7 GND 0.088471f
C243 a_n7729_8946.t2 GND 0.088471f
C244 a_n7729_8946.n3 GND 0.578656f
C245 a_n7729_8946.n4 GND 2.71687f
C246 a_n7729_8946.t8 GND 0.088471f
C247 a_n7729_8946.t4 GND 0.088471f
C248 a_n7729_8946.n5 GND 0.578654f
C249 a_n7729_8946.n6 GND 3.66867f
C250 a_n7729_8946.t16 GND 0.688016f
C251 a_n7729_8946.t10 GND 0.088471f
C252 a_n7729_8946.t17 GND 0.088471f
C253 a_n7729_8946.n7 GND 0.475466f
C254 a_n7729_8946.n8 GND 2.79828f
C255 a_n7729_8946.t11 GND 0.66854f
C256 a_n7729_8946.t13 GND 0.66854f
C257 a_n7729_8946.t12 GND 0.088471f
C258 a_n7729_8946.t14 GND 0.088471f
C259 a_n7729_8946.n9 GND 0.475466f
C260 a_n7729_8946.n10 GND 1.69462f
C261 a_n7729_8946.t15 GND 0.66854f
C262 a_n7729_8946.n11 GND 2.00394f
C263 a_n7729_8946.n12 GND 4.583971f
C264 a_n7729_8946.n13 GND 0.578657f
C265 a_n7729_8946.t9 GND 0.088471f
C266 a_n7651_8750.n0 GND 3.42019f
C267 a_n7651_8750.n1 GND 0.951635f
C268 a_n7651_8750.n2 GND 0.938637f
C269 a_n7651_8750.n3 GND 3.31569f
C270 a_n7651_8750.n4 GND 0.951635f
C271 a_n7651_8750.n5 GND 0.938637f
C272 a_n7651_8750.n6 GND 3.41275f
C273 a_n7651_8750.n7 GND 4.87931f
C274 a_n7651_8750.n8 GND 0.605577f
C275 a_n7651_8750.n9 GND 13.5029f
C276 a_n7651_8750.n10 GND 3.05261f
C277 a_n7651_8750.n11 GND 0.940635f
C278 a_n7651_8750.n12 GND 1.59093f
C279 a_n7651_8750.n13 GND 0.940781f
C280 a_n7651_8750.n14 GND 0.945104f
C281 a_n7651_8750.n15 GND 7.29866f
C282 a_n7651_8750.n16 GND 0.124941f
C283 a_n7651_8750.n17 GND 0.086333f
C284 a_n7651_8750.n18 GND 0.9411f
C285 a_n7651_8750.n19 GND 0.943357f
C286 a_n7651_8750.n20 GND 0.007848f
C287 a_n7651_8750.n21 GND 0.031708f
C288 a_n7651_8750.n22 GND 0.611075f
C289 a_n7651_8750.n23 GND 3.23469f
C290 a_n7651_8750.n24 GND 0.252741f
C291 a_n7651_8750.n25 GND 0.017942f
C292 a_n7651_8750.n26 GND 0.203634f
C293 a_n7651_8750.n27 GND 0.01519f
C294 a_n7651_8750.n28 GND 5.415009f
C295 a_n7651_8750.n29 GND 0.013079f
C296 a_n7651_8750.n30 GND 0.017546f
C297 a_n7651_8750.n31 GND 0.134786f
C298 a_n7651_8750.n32 GND 0.013079f
C299 a_n7651_8750.n33 GND 0.017546f
C300 a_n7651_8750.n34 GND 0.050998f
C301 a_n7651_8750.t27 GND 0.283552f
C302 a_n7651_8750.t21 GND 0.29974f
C303 a_n7651_8750.t23 GND 0.044484f
C304 a_n7651_8750.t14 GND 1.90346f
C305 a_n7651_8750.t10 GND 1.9472f
C306 a_n7651_8750.t26 GND 1.86893f
C307 a_n7651_8750.t22 GND 1.88848f
C308 a_n7651_8750.t20 GND 1.93106f
C309 a_n7651_8750.t50 GND 1.90346f
C310 a_n7651_8750.t37 GND 1.9472f
C311 a_n7651_8750.t41 GND 1.86893f
C312 a_n7651_8750.t51 GND 1.88848f
C313 a_n7651_8750.t38 GND 1.93106f
C314 a_n7651_8750.t18 GND 1.90346f
C315 a_n7651_8750.t28 GND 1.89057f
C316 a_n7651_8750.t24 GND 1.44893f
C317 a_n7651_8750.t12 GND 1.44893f
C318 a_n7651_8750.t16 GND 1.90346f
C319 a_n7651_8750.t44 GND 1.93969f
C320 a_n7651_8750.t43 GND 1.88638f
C321 a_n7651_8750.t54 GND 1.87118f
C322 a_n7651_8750.t42 GND 1.94023f
C323 a_n7651_8750.t33 GND 1.90346f
C324 a_n7651_8750.n35 GND 0.801773f
C325 a_n7651_8750.t9 GND 0.030593f
C326 a_n7651_8750.n36 GND 0.037147f
C327 a_n7651_8750.n37 GND 0.073774f
C328 a_n7651_8750.t0 GND 0.329141f
C329 a_n7651_8750.t4 GND 0.036021f
C330 a_n7651_8750.t3 GND 0.347985f
C331 a_n7651_8750.t8 GND 0.036021f
C332 a_n7651_8750.t2 GND 0.030593f
C333 a_n7651_8750.n38 GND 0.037147f
C334 a_n7651_8750.t7 GND 0.329142f
C335 a_n7651_8750.t5 GND 0.036021f
C336 a_n7651_8750.t1 GND 0.347986f
C337 a_n7651_8750.t6 GND 0.036021f
C338 a_n7651_8750.n39 GND 0.809687f
C339 a_n7651_8750.t17 GND 0.34594f
C340 a_n7651_8750.t25 GND 0.283552f
C341 a_n7651_8750.t13 GND 0.044484f
C342 a_n7651_8750.t19 GND 0.283552f
C343 a_n7651_8750.t29 GND 0.044484f
C344 a_n7651_8750.t55 GND 1.95887f
C345 a_n7651_8750.t39 GND 1.88157f
C346 a_n7651_8750.t48 GND 1.88278f
C347 a_n7651_8750.t32 GND 1.91411f
C348 a_n7651_8750.t49 GND 1.90498f
C349 a_n7651_8750.t52 GND 1.88256f
C350 a_n7651_8750.t40 GND 1.93599f
C351 a_n7651_8750.t53 GND 1.91411f
C352 a_n7651_8750.t31 GND 1.95912f
C353 a_n7651_8750.t47 GND 1.88146f
C354 a_n7651_8750.t30 GND 1.88278f
C355 a_n7651_8750.t46 GND 1.91411f
C356 a_n7651_8750.t36 GND 1.90498f
C357 a_n7651_8750.t45 GND 1.8856f
C358 a_n7651_8750.t35 GND 1.92065f
C359 a_n7651_8750.t34 GND 1.91411f
C360 a_n7651_8750.t15 GND 0.336146f
C361 a_n7651_8750.t11 GND 0.044484f
C362 a_n6364_n172.n0 GND 1.86772f
C363 a_n6364_n172.n1 GND 1.86772f
C364 a_n6364_n172.n2 GND 2.90872f
C365 a_n6364_n172.n3 GND 3.33404f
C366 a_n6364_n172.n4 GND 4.04533f
C367 a_n6364_n172.n5 GND 0.23323f
C368 a_n6364_n172.n6 GND 0.017397f
C369 a_n6364_n172.n7 GND 0.23323f
C370 a_n6364_n172.n8 GND 0.017397f
C371 a_n6364_n172.n9 GND 0.017397f
C372 a_n6364_n172.n10 GND 0.024411f
C373 a_n6364_n172.n11 GND 0.017397f
C374 a_n6364_n172.n12 GND 0.024411f
C375 a_n6364_n172.n13 GND 0.017397f
C376 a_n6364_n172.n14 GND 0.024411f
C377 a_n6364_n172.n15 GND 0.017397f
C378 a_n6364_n172.n16 GND 0.024411f
C379 a_n6364_n172.n17 GND 0.017397f
C380 a_n6364_n172.n18 GND 0.024411f
C381 a_n6364_n172.n19 GND 0.017397f
C382 a_n6364_n172.n20 GND 0.024411f
C383 a_n6364_n172.n21 GND 0.23323f
C384 a_n6364_n172.n22 GND 0.017397f
C385 a_n6364_n172.n23 GND 0.23323f
C386 a_n6364_n172.n24 GND 0.017397f
C387 a_n6364_n172.n25 GND 0.01498f
C388 a_n6364_n172.n26 GND 0.020096f
C389 a_n6364_n172.n27 GND 0.05841f
C390 a_n6364_n172.n28 GND 0.01498f
C391 a_n6364_n172.n29 GND 0.020096f
C392 a_n6364_n172.n30 GND 0.05841f
C393 a_n6364_n172.n31 GND 0.019756f
C394 a_n6364_n172.n32 GND 0.054282f
C395 a_n6364_n172.n33 GND 0.019756f
C396 a_n6364_n172.n34 GND 0.054282f
C397 a_n6364_n172.n35 GND 0.019756f
C398 a_n6364_n172.n36 GND 0.054282f
C399 a_n6364_n172.n37 GND 0.019756f
C400 a_n6364_n172.n38 GND 0.054282f
C401 a_n6364_n172.n39 GND 0.019756f
C402 a_n6364_n172.n40 GND 0.054282f
C403 a_n6364_n172.n41 GND 0.019756f
C404 a_n6364_n172.n42 GND 0.054282f
C405 a_n6364_n172.n43 GND 0.01498f
C406 a_n6364_n172.n44 GND 0.020096f
C407 a_n6364_n172.n45 GND 0.05841f
C408 a_n6364_n172.n46 GND 0.01498f
C409 a_n6364_n172.n47 GND 0.020096f
C410 a_n6364_n172.n48 GND 0.05841f
C411 a_n6364_n172.n49 GND 0.155273f
C412 a_n6364_n172.n50 GND 0.155273f
C413 a_n6364_n172.n51 GND 0.155273f
C414 a_n6364_n172.n52 GND 0.155273f
C415 a_n6364_n172.n53 GND 0.155273f
C416 a_n6364_n172.n54 GND 0.155273f
C417 a_n6364_n172.t18 GND 0.041256f
C418 a_n6364_n172.n55 GND 0.022528f
C419 a_n6364_n172.t10 GND 0.035039f
C420 a_n6364_n172.n56 GND 0.019973f
C421 a_n6364_n172.n57 GND 0.043988f
C422 a_n6364_n172.n58 GND 0.008947f
C423 a_n6364_n172.n59 GND 0.00845f
C424 a_n6364_n172.n60 GND 0.02848f
C425 a_n6364_n172.t11 GND 0.035266f
C426 a_n6364_n172.n61 GND 0.035996f
C427 a_n6364_n172.n62 GND 0.145086f
C428 a_n6364_n172.t7 GND 0.041256f
C429 a_n6364_n172.t3 GND 0.041256f
C430 a_n6364_n172.n63 GND 0.292878f
C431 a_n6364_n172.n64 GND 1.21057f
C432 a_n6364_n172.t4 GND 0.041256f
C433 a_n6364_n172.t12 GND 0.041256f
C434 a_n6364_n172.n65 GND 0.292878f
C435 a_n6364_n172.n66 GND 1.87123f
C436 a_n6364_n172.t0 GND 0.035266f
C437 a_n6364_n172.n67 GND 0.035996f
C438 a_n6364_n172.n68 GND 0.145086f
C439 a_n6364_n172.t8 GND 0.035266f
C440 a_n6364_n172.n69 GND 0.035996f
C441 a_n6364_n172.n70 GND 0.145086f
C442 a_n6364_n172.t2 GND 0.035266f
C443 a_n6364_n172.n71 GND 0.035996f
C444 a_n6364_n172.n72 GND 0.145086f
C445 a_n6364_n172.t9 GND 0.035266f
C446 a_n6364_n172.n73 GND 0.035996f
C447 a_n6364_n172.n74 GND 0.145086f
C448 a_n6364_n172.t25 GND 0.035266f
C449 a_n6364_n172.n75 GND 0.035996f
C450 a_n6364_n172.n76 GND 0.145086f
C451 a_n6364_n172.n77 GND 1.3483f
C452 a_n6364_n172.t19 GND 0.041256f
C453 a_n6364_n172.t20 GND 0.041256f
C454 a_n6364_n172.n78 GND 0.292876f
C455 a_n6364_n172.n79 GND 1.67223f
C456 a_n6364_n172.t17 GND 0.041256f
C457 a_n6364_n172.t21 GND 0.041256f
C458 a_n6364_n172.n80 GND 0.292876f
C459 a_n6364_n172.n81 GND 1.21057f
C460 a_n6364_n172.n82 GND 0.022528f
C461 a_n6364_n172.t15 GND 0.035039f
C462 a_n6364_n172.n83 GND 0.019973f
C463 a_n6364_n172.n84 GND 0.043988f
C464 a_n6364_n172.n85 GND 0.008947f
C465 a_n6364_n172.n86 GND 0.00845f
C466 a_n6364_n172.n87 GND 0.02848f
C467 a_n6364_n172.t24 GND 0.041256f
C468 a_n6364_n172.t1 GND 0.041256f
C469 a_n6364_n172.n88 GND 0.292876f
C470 a_n6364_n172.t6 GND 0.041256f
C471 a_n6364_n172.t5 GND 0.041256f
C472 a_n6364_n172.n89 GND 0.292876f
C473 a_n6364_n172.n90 GND 1.21057f
C474 a_n6364_n172.n91 GND 0.022528f
C475 a_n6364_n172.t23 GND 0.035039f
C476 a_n6364_n172.n92 GND 0.019973f
C477 a_n6364_n172.n93 GND 0.043988f
C478 a_n6364_n172.n94 GND 0.008947f
C479 a_n6364_n172.n95 GND 0.00845f
C480 a_n6364_n172.n96 GND 0.02848f
C481 a_n6364_n172.n97 GND 1.18091f
C482 a_n6364_n172.n98 GND 1.54646f
C483 a_n6364_n172.n99 GND 0.022528f
C484 a_n6364_n172.t16 GND 0.035039f
C485 a_n6364_n172.n100 GND 0.019973f
C486 a_n6364_n172.n101 GND 0.043988f
C487 a_n6364_n172.n102 GND 0.008947f
C488 a_n6364_n172.n103 GND 0.00845f
C489 a_n6364_n172.n104 GND 0.02848f
C490 a_n6364_n172.n105 GND 1.34107f
C491 a_n6364_n172.t14 GND 0.041256f
C492 a_n6364_n172.t13 GND 0.041256f
C493 a_n6364_n172.n106 GND 0.292878f
C494 a_n6364_n172.n107 GND 1.21057f
C495 a_n6364_n172.n108 GND 0.292878f
C496 a_n6364_n172.t22 GND 0.041256f
C497 a_n18960_7900.n0 GND 1.11186f
C498 a_n18960_7900.n1 GND 5.19338f
C499 a_n18960_7900.n2 GND 1.11186f
C500 a_n18960_7900.n3 GND 5.13325f
C501 a_n18960_7900.n4 GND 1.11758f
C502 a_n18960_7900.n5 GND 1.11758f
C503 a_n18960_7900.n6 GND 4.39183f
C504 a_n18960_7900.n7 GND 1.1221f
C505 a_n18960_7900.n8 GND 4.45195f
C506 a_n18960_7900.n9 GND 1.1221f
C507 a_n18960_7900.n10 GND 0.738446f
C508 a_n18960_7900.n11 GND 0.738446f
C509 a_n18960_7900.n12 GND 2.1937f
C510 a_n18960_7900.n13 GND 1.17718f
C511 a_n18960_7900.n14 GND 19.007599f
C512 a_n18960_7900.n15 GND 0.728193f
C513 a_n18960_7900.n16 GND 0.728193f
C514 a_n18960_7900.n17 GND 4.96886f
C515 a_n18960_7900.n18 GND 4.21559f
C516 a_n18960_7900.n19 GND 3.22039f
C517 a_n18960_7900.n20 GND 4.83279f
C518 a_n18960_7900.t5 GND 0.291444f
C519 a_n18960_7900.t3 GND 0.037285f
C520 a_n18960_7900.t19 GND 0.281156f
C521 a_n18960_7900.t6 GND 0.037285f
C522 a_n18960_7900.t4 GND 0.326937f
C523 a_n18960_7900.t11 GND 0.222889f
C524 a_n18960_7900.t17 GND 0.27588f
C525 a_n18960_7900.t13 GND 0.030192f
C526 a_n18960_7900.t10 GND 0.222185f
C527 a_n18960_7900.t16 GND 0.27588f
C528 a_n18960_7900.t12 GND 0.030192f
C529 a_n18960_7900.t15 GND 0.291675f
C530 a_n18960_7900.t9 GND 0.030192f
C531 a_n18960_7900.t8 GND 0.27588f
C532 a_n18960_7900.t14 GND 0.030192f
C533 a_n18960_7900.t30 GND 2.59781f
C534 a_n18960_7900.t40 GND 2.00593f
C535 a_n18960_7900.n21 GND 0.98648f
C536 a_n18960_7900.t32 GND 2.56583f
C537 a_n18960_7900.t42 GND 2.59998f
C538 a_n18960_7900.t43 GND 2.57777f
C539 a_n18960_7900.t45 GND 2.57374f
C540 a_n18960_7900.t47 GND 2.61211f
C541 a_n18960_7900.t20 GND 2.59781f
C542 a_n18960_7900.t28 GND 2.00593f
C543 a_n18960_7900.n22 GND 0.98648f
C544 a_n18960_7900.t21 GND 2.56583f
C545 a_n18960_7900.t31 GND 2.59998f
C546 a_n18960_7900.t33 GND 2.57777f
C547 a_n18960_7900.t35 GND 2.57374f
C548 a_n18960_7900.t37 GND 2.61211f
C549 a_n18960_7900.t22 GND 2.58673f
C550 a_n18960_7900.t24 GND 2.56975f
C551 a_n18960_7900.t34 GND 2.60963f
C552 a_n18960_7900.t36 GND 2.55976f
C553 a_n18960_7900.t38 GND 2.57895f
C554 a_n18960_7900.t39 GND 2.6206f
C555 a_n18960_7900.t41 GND 2.61211f
C556 a_n18960_7900.t44 GND 2.58673f
C557 a_n18960_7900.t46 GND 2.56975f
C558 a_n18960_7900.t23 GND 2.60963f
C559 a_n18960_7900.t25 GND 2.55976f
C560 a_n18960_7900.t26 GND 2.57895f
C561 a_n18960_7900.t27 GND 2.6206f
C562 a_n18960_7900.t29 GND 2.61211f
C563 a_n18960_7900.n23 GND 5.83353f
C564 a_n18960_7900.t7 GND 0.281156f
C565 a_n18960_7900.t18 GND 0.037285f
C566 a_n18960_7900.t1 GND 0.281156f
C567 a_n18960_7900.t2 GND 0.037285f
C568 a_n18960_7900.t0 GND 0.333162f
C569 VN.n0 GND 0.029143f
C570 VN.t8 GND 0.619175f
C571 VN.n1 GND 0.02333f
C572 VN.n2 GND 0.012581f
C573 VN.n3 GND 0.020551f
C574 VN.n4 GND 0.012581f
C575 VN.n5 GND 0.02333f
C576 VN.n6 GND 0.012581f
C577 VN.t7 GND 0.619175f
C578 VN.n7 GND 0.02333f
C579 VN.n8 GND 0.012581f
C580 VN.n9 GND 0.012048f
C581 VN.n10 GND 0.012581f
C582 VN.n11 GND 0.02333f
C583 VN.n12 GND 0.012581f
C584 VN.t10 GND 0.619175f
C585 VN.n13 GND 0.02333f
C586 VN.n14 GND 0.012581f
C587 VN.n15 GND 0.012048f
C588 VN.n16 GND 0.012581f
C589 VN.n17 GND 0.02333f
C590 VN.n18 GND 0.156837f
C591 VN.t6 GND 0.619175f
C592 VN.t12 GND 0.874399f
C593 VN.n19 GND 0.41809f
C594 VN.n20 GND 0.291049f
C595 VN.n21 GND 0.01665f
C596 VN.n22 GND 0.02333f
C597 VN.n23 GND 0.012581f
C598 VN.n24 GND 0.012581f
C599 VN.n25 GND 0.012581f
C600 VN.n26 GND 0.02333f
C601 VN.n27 GND 0.02333f
C602 VN.n28 GND 0.022855f
C603 VN.n29 GND 0.012581f
C604 VN.n30 GND 0.012581f
C605 VN.n31 GND 0.012581f
C606 VN.n32 GND 0.025003f
C607 VN.n33 GND 0.02333f
C608 VN.n34 GND 0.02333f
C609 VN.n35 GND 0.012581f
C610 VN.n36 GND 0.012581f
C611 VN.n37 GND 0.012581f
C612 VN.n38 GND 0.02333f
C613 VN.n39 GND 0.252756f
C614 VN.n40 GND 0.02333f
C615 VN.n41 GND 0.012581f
C616 VN.n42 GND 0.012581f
C617 VN.n43 GND 0.012581f
C618 VN.n44 GND 0.02333f
C619 VN.n45 GND 0.02333f
C620 VN.n46 GND 0.025003f
C621 VN.n47 GND 0.012581f
C622 VN.n48 GND 0.012581f
C623 VN.n49 GND 0.012581f
C624 VN.n50 GND 0.022855f
C625 VN.n51 GND 0.02333f
C626 VN.n52 GND 0.02333f
C627 VN.n53 GND 0.012581f
C628 VN.n54 GND 0.012581f
C629 VN.n55 GND 0.012581f
C630 VN.n56 GND 0.02333f
C631 VN.n57 GND 0.01665f
C632 VN.n58 GND 0.240944f
C633 VN.n59 GND 0.018493f
C634 VN.n60 GND 0.012581f
C635 VN.n61 GND 0.012581f
C636 VN.n62 GND 0.012581f
C637 VN.n63 GND 0.02333f
C638 VN.n64 GND 0.02333f
C639 VN.n65 GND 0.02333f
C640 VN.n66 GND 0.012581f
C641 VN.n67 GND 0.012581f
C642 VN.n68 GND 0.012581f
C643 VN.n69 GND 0.016026f
C644 VN.n70 GND 0.02333f
C645 VN.n71 GND 0.02333f
C646 VN.n72 GND 0.012581f
C647 VN.n73 GND 0.012581f
C648 VN.n74 GND 0.012581f
C649 VN.n75 GND 0.02333f
C650 VN.n76 GND 0.021487f
C651 VN.n77 GND 0.298956f
C652 VN.n78 GND 0.289357f
C653 VN.n79 GND 0.029143f
C654 VN.t11 GND 0.619175f
C655 VN.n80 GND 0.02333f
C656 VN.n81 GND 0.012581f
C657 VN.n82 GND 0.020551f
C658 VN.n83 GND 0.012581f
C659 VN.n84 GND 0.02333f
C660 VN.n85 GND 0.012581f
C661 VN.t14 GND 0.619175f
C662 VN.n86 GND 0.02333f
C663 VN.n87 GND 0.012581f
C664 VN.n88 GND 0.012048f
C665 VN.n89 GND 0.012581f
C666 VN.n90 GND 0.02333f
C667 VN.n91 GND 0.012581f
C668 VN.t13 GND 0.619175f
C669 VN.n92 GND 0.02333f
C670 VN.n93 GND 0.012581f
C671 VN.n94 GND 0.012048f
C672 VN.n95 GND 0.012581f
C673 VN.n96 GND 0.02333f
C674 VN.n97 GND 0.156837f
C675 VN.t5 GND 0.619175f
C676 VN.t9 GND 0.874401f
C677 VN.n98 GND 0.418087f
C678 VN.n99 GND 0.291049f
C679 VN.n100 GND 0.01665f
C680 VN.n101 GND 0.02333f
C681 VN.n102 GND 0.012581f
C682 VN.n103 GND 0.012581f
C683 VN.n104 GND 0.012581f
C684 VN.n105 GND 0.02333f
C685 VN.n106 GND 0.02333f
C686 VN.n107 GND 0.022855f
C687 VN.n108 GND 0.012581f
C688 VN.n109 GND 0.012581f
C689 VN.n110 GND 0.012581f
C690 VN.n111 GND 0.025003f
C691 VN.n112 GND 0.02333f
C692 VN.n113 GND 0.02333f
C693 VN.n114 GND 0.012581f
C694 VN.n115 GND 0.012581f
C695 VN.n116 GND 0.012581f
C696 VN.n117 GND 0.02333f
C697 VN.n118 GND 0.252756f
C698 VN.n119 GND 0.02333f
C699 VN.n120 GND 0.012581f
C700 VN.n121 GND 0.012581f
C701 VN.n122 GND 0.012581f
C702 VN.n123 GND 0.02333f
C703 VN.n124 GND 0.02333f
C704 VN.n125 GND 0.025003f
C705 VN.n126 GND 0.012581f
C706 VN.n127 GND 0.012581f
C707 VN.n128 GND 0.012581f
C708 VN.n129 GND 0.022855f
C709 VN.n130 GND 0.02333f
C710 VN.n131 GND 0.02333f
C711 VN.n132 GND 0.012581f
C712 VN.n133 GND 0.012581f
C713 VN.n134 GND 0.012581f
C714 VN.n135 GND 0.02333f
C715 VN.n136 GND 0.01665f
C716 VN.n137 GND 0.240944f
C717 VN.n138 GND 0.018493f
C718 VN.n139 GND 0.012581f
C719 VN.n140 GND 0.012581f
C720 VN.n141 GND 0.012581f
C721 VN.n142 GND 0.02333f
C722 VN.n143 GND 0.02333f
C723 VN.n144 GND 0.02333f
C724 VN.n145 GND 0.012581f
C725 VN.n146 GND 0.012581f
C726 VN.n147 GND 0.012581f
C727 VN.n148 GND 0.016026f
C728 VN.n149 GND 0.02333f
C729 VN.n150 GND 0.02333f
C730 VN.n151 GND 0.012581f
C731 VN.n152 GND 0.012581f
C732 VN.n153 GND 0.012581f
C733 VN.n154 GND 0.02333f
C734 VN.n155 GND 0.021487f
C735 VN.n156 GND 0.298956f
C736 VN.n157 GND 0.89032f
C737 VN.n158 GND 1.03195f
C738 VN.t0 GND 0.021718f
C739 VN.t1 GND 0.003878f
C740 VN.t3 GND 0.003878f
C741 VN.n159 GND 0.012578f
C742 VN.n160 GND 0.097644f
C743 VN.t2 GND 0.003878f
C744 VN.t4 GND 0.003878f
C745 VN.n161 GND 0.012578f
C746 VN.n162 GND 0.073294f
C747 VN.n163 GND 3.75938f
C748 VOUT.t45 GND 0.03183f
C749 VOUT.t44 GND 0.03183f
C750 VOUT.n0 GND 0.231089f
C751 VOUT.t5 GND 0.03183f
C752 VOUT.t51 GND 0.03183f
C753 VOUT.n1 GND 0.218252f
C754 VOUT.n2 GND 1.24961f
C755 VOUT.t46 GND 0.03183f
C756 VOUT.t43 GND 0.03183f
C757 VOUT.n3 GND 0.218252f
C758 VOUT.n4 GND 0.627924f
C759 VOUT.t50 GND 0.290493f
C760 VOUT.n5 GND 0.537695f
C761 VOUT.t16 GND 0.03183f
C762 VOUT.t47 GND 0.03183f
C763 VOUT.n6 GND 0.231089f
C764 VOUT.t49 GND 0.03183f
C765 VOUT.t13 GND 0.03183f
C766 VOUT.n7 GND 0.218252f
C767 VOUT.n8 GND 1.24961f
C768 VOUT.t3 GND 0.03183f
C769 VOUT.t48 GND 0.03183f
C770 VOUT.n9 GND 0.218252f
C771 VOUT.n10 GND 0.627924f
C772 VOUT.t14 GND 0.290493f
C773 VOUT.n11 GND 0.489379f
C774 VOUT.n12 GND 0.822305f
C775 VOUT.n13 GND 13.5615f
C776 VOUT.t52 GND 2.73334f
C777 VOUT.t53 GND 3.84558f
C778 VOUT.n14 GND 6.61929f
C779 VOUT.n15 GND 2.26893f
C780 VOUT.t7 GND 0.298038f
C781 VOUT.t12 GND 0.03183f
C782 VOUT.t42 GND 0.03183f
C783 VOUT.n16 GND 0.218252f
C784 VOUT.n17 GND 1.01385f
C785 VOUT.t4 GND 0.03183f
C786 VOUT.t11 GND 0.03183f
C787 VOUT.n18 GND 0.218252f
C788 VOUT.n19 GND 0.627924f
C789 VOUT.t0 GND 0.03183f
C790 VOUT.t9 GND 0.03183f
C791 VOUT.n20 GND 0.218252f
C792 VOUT.n21 GND 0.735745f
C793 VOUT.t8 GND 0.298038f
C794 VOUT.t15 GND 0.03183f
C795 VOUT.t10 GND 0.03183f
C796 VOUT.n22 GND 0.218252f
C797 VOUT.n23 GND 1.01385f
C798 VOUT.t17 GND 0.03183f
C799 VOUT.t2 GND 0.03183f
C800 VOUT.n24 GND 0.218252f
C801 VOUT.n25 GND 0.627924f
C802 VOUT.t6 GND 0.03183f
C803 VOUT.t1 GND 0.03183f
C804 VOUT.n26 GND 0.218251f
C805 VOUT.n27 GND 0.685262f
C806 VOUT.n28 GND 0.91046f
C807 VOUT.n29 GND 16.488401f
C808 VOUT.t32 GND 0.024325f
C809 VOUT.t23 GND 0.024325f
C810 VOUT.n30 GND 0.221969f
C811 VOUT.t36 GND 0.024325f
C812 VOUT.t24 GND 0.024325f
C813 VOUT.n31 GND 0.203199f
C814 VOUT.n32 GND 1.2474f
C815 VOUT.t39 GND 0.024325f
C816 VOUT.t29 GND 0.024325f
C817 VOUT.n33 GND 0.203199f
C818 VOUT.n34 GND 0.719995f
C819 VOUT.t38 GND 0.024325f
C820 VOUT.t30 GND 0.024325f
C821 VOUT.n35 GND 0.221969f
C822 VOUT.t26 GND 0.024325f
C823 VOUT.t19 GND 0.024325f
C824 VOUT.n36 GND 0.203199f
C825 VOUT.n37 GND 1.2474f
C826 VOUT.t34 GND 0.024325f
C827 VOUT.t28 GND 0.024325f
C828 VOUT.n38 GND 0.203199f
C829 VOUT.n39 GND 0.679971f
C830 VOUT.n40 GND 0.894057f
C831 VOUT.n41 GND 16.243f
C832 VOUT.t27 GND 0.024325f
C833 VOUT.t37 GND 0.024325f
C834 VOUT.n42 GND 0.221969f
C835 VOUT.t22 GND 0.024325f
C836 VOUT.t41 GND 0.024325f
C837 VOUT.n43 GND 0.203199f
C838 VOUT.n44 GND 1.2474f
C839 VOUT.t31 GND 0.024325f
C840 VOUT.t18 GND 0.024325f
C841 VOUT.n45 GND 0.203199f
C842 VOUT.n46 GND 0.719995f
C843 VOUT.t20 GND 0.024325f
C844 VOUT.t25 GND 0.024325f
C845 VOUT.n47 GND 0.221969f
C846 VOUT.t35 GND 0.024325f
C847 VOUT.t33 GND 0.024325f
C848 VOUT.n48 GND 0.203199f
C849 VOUT.n49 GND 1.2474f
C850 VOUT.t40 GND 0.024325f
C851 VOUT.t21 GND 0.024325f
C852 VOUT.n50 GND 0.203199f
C853 VOUT.n51 GND 0.679971f
C854 VOUT.n52 GND 0.894057f
C855 VOUT.n53 GND 12.7305f
C856 VOUT.n54 GND 6.53377f
C857 CS_BIAS.n0 GND 0.009829f
C858 CS_BIAS.t33 GND 0.24163f
C859 CS_BIAS.n1 GND 0.007868f
C860 CS_BIAS.n2 GND 0.004243f
C861 CS_BIAS.n3 GND 0.006403f
C862 CS_BIAS.n4 GND 0.004243f
C863 CS_BIAS.n5 GND 0.007868f
C864 CS_BIAS.n6 GND 0.004243f
C865 CS_BIAS.t42 GND 0.24163f
C866 CS_BIAS.n7 GND 0.007868f
C867 CS_BIAS.n8 GND 0.004243f
C868 CS_BIAS.n9 GND 0.003432f
C869 CS_BIAS.n10 GND 0.004243f
C870 CS_BIAS.n11 GND 0.007868f
C871 CS_BIAS.n12 GND 0.004243f
C872 CS_BIAS.t29 GND 0.24163f
C873 CS_BIAS.n13 GND 0.007868f
C874 CS_BIAS.n14 GND 0.004243f
C875 CS_BIAS.n15 GND 0.006168f
C876 CS_BIAS.n16 GND 0.004243f
C877 CS_BIAS.n17 GND 0.007868f
C878 CS_BIAS.n18 GND 0.004243f
C879 CS_BIAS.t41 GND 0.24163f
C880 CS_BIAS.n19 GND 0.007868f
C881 CS_BIAS.n20 GND 0.004243f
C882 CS_BIAS.n21 GND 0.008428f
C883 CS_BIAS.n22 GND 0.004243f
C884 CS_BIAS.n23 GND 0.007868f
C885 CS_BIAS.n24 GND 0.004243f
C886 CS_BIAS.t26 GND 0.24163f
C887 CS_BIAS.n25 GND 0.108683f
C888 CS_BIAS.t36 GND 0.332305f
C889 CS_BIAS.n26 GND 0.147953f
C890 CS_BIAS.n27 GND 0.05348f
C891 CS_BIAS.n28 GND 0.005072f
C892 CS_BIAS.n29 GND 0.007868f
C893 CS_BIAS.n30 GND 0.007868f
C894 CS_BIAS.n31 GND 0.004243f
C895 CS_BIAS.n32 GND 0.004243f
C896 CS_BIAS.n33 GND 0.004243f
C897 CS_BIAS.n34 GND 0.007868f
C898 CS_BIAS.n35 GND 0.008344f
C899 CS_BIAS.n36 GND 0.003432f
C900 CS_BIAS.n37 GND 0.004243f
C901 CS_BIAS.n38 GND 0.004243f
C902 CS_BIAS.n39 GND 0.004243f
C903 CS_BIAS.n40 GND 0.007868f
C904 CS_BIAS.n41 GND 0.007868f
C905 CS_BIAS.n42 GND 0.007868f
C906 CS_BIAS.n43 GND 0.004243f
C907 CS_BIAS.n44 GND 0.004243f
C908 CS_BIAS.n45 GND 0.004243f
C909 CS_BIAS.n46 GND 0.004916f
C910 CS_BIAS.n47 GND 0.092263f
C911 CS_BIAS.n48 GND 0.006936f
C912 CS_BIAS.n49 GND 0.007868f
C913 CS_BIAS.n50 GND 0.004243f
C914 CS_BIAS.n51 GND 0.004243f
C915 CS_BIAS.n52 GND 0.004243f
C916 CS_BIAS.n53 GND 0.007868f
C917 CS_BIAS.n54 GND 0.007868f
C918 CS_BIAS.n55 GND 0.006168f
C919 CS_BIAS.n56 GND 0.003707f
C920 CS_BIAS.n57 GND 0.009829f
C921 CS_BIAS.t14 GND 0.24163f
C922 CS_BIAS.n58 GND 0.007868f
C923 CS_BIAS.n59 GND 0.004243f
C924 CS_BIAS.n60 GND 0.006403f
C925 CS_BIAS.n61 GND 0.004243f
C926 CS_BIAS.n62 GND 0.007868f
C927 CS_BIAS.n63 GND 0.004243f
C928 CS_BIAS.t20 GND 0.24163f
C929 CS_BIAS.n64 GND 0.007868f
C930 CS_BIAS.n65 GND 0.004243f
C931 CS_BIAS.n66 GND 0.003432f
C932 CS_BIAS.n67 GND 0.004243f
C933 CS_BIAS.n68 GND 0.007868f
C934 CS_BIAS.n69 GND 0.004243f
C935 CS_BIAS.t22 GND 0.24163f
C936 CS_BIAS.n70 GND 0.007868f
C937 CS_BIAS.n71 GND 0.004243f
C938 CS_BIAS.n72 GND 0.006168f
C939 CS_BIAS.n73 GND 0.004243f
C940 CS_BIAS.n74 GND 0.007868f
C941 CS_BIAS.n75 GND 0.004243f
C942 CS_BIAS.t12 GND 0.24163f
C943 CS_BIAS.n76 GND 0.007868f
C944 CS_BIAS.n77 GND 0.004243f
C945 CS_BIAS.n78 GND 0.008428f
C946 CS_BIAS.n79 GND 0.004243f
C947 CS_BIAS.n80 GND 0.007868f
C948 CS_BIAS.n81 GND 0.004243f
C949 CS_BIAS.t16 GND 0.24163f
C950 CS_BIAS.n82 GND 0.108683f
C951 CS_BIAS.t10 GND 0.332305f
C952 CS_BIAS.n83 GND 0.147953f
C953 CS_BIAS.n84 GND 0.05348f
C954 CS_BIAS.n85 GND 0.005072f
C955 CS_BIAS.n86 GND 0.007868f
C956 CS_BIAS.n87 GND 0.007868f
C957 CS_BIAS.n88 GND 0.004243f
C958 CS_BIAS.n89 GND 0.004243f
C959 CS_BIAS.n90 GND 0.004243f
C960 CS_BIAS.n91 GND 0.007868f
C961 CS_BIAS.n92 GND 0.008344f
C962 CS_BIAS.n93 GND 0.003432f
C963 CS_BIAS.n94 GND 0.004243f
C964 CS_BIAS.n95 GND 0.004243f
C965 CS_BIAS.n96 GND 0.004243f
C966 CS_BIAS.n97 GND 0.007868f
C967 CS_BIAS.n98 GND 0.007868f
C968 CS_BIAS.n99 GND 0.007868f
C969 CS_BIAS.n100 GND 0.004243f
C970 CS_BIAS.n101 GND 0.004243f
C971 CS_BIAS.n102 GND 0.004243f
C972 CS_BIAS.n103 GND 0.004916f
C973 CS_BIAS.n104 GND 0.092263f
C974 CS_BIAS.n105 GND 0.006936f
C975 CS_BIAS.n106 GND 0.007868f
C976 CS_BIAS.n107 GND 0.004243f
C977 CS_BIAS.n108 GND 0.004243f
C978 CS_BIAS.n109 GND 0.004243f
C979 CS_BIAS.n110 GND 0.007868f
C980 CS_BIAS.n111 GND 0.007868f
C981 CS_BIAS.n112 GND 0.006168f
C982 CS_BIAS.n113 GND 0.004243f
C983 CS_BIAS.n114 GND 0.004243f
C984 CS_BIAS.n115 GND 0.004243f
C985 CS_BIAS.n116 GND 0.007868f
C986 CS_BIAS.n117 GND 0.007868f
C987 CS_BIAS.n118 GND 0.007868f
C988 CS_BIAS.n119 GND 0.004243f
C989 CS_BIAS.n120 GND 0.004243f
C990 CS_BIAS.n121 GND 0.004243f
C991 CS_BIAS.n122 GND 0.006936f
C992 CS_BIAS.n123 GND 0.092263f
C993 CS_BIAS.n124 GND 0.004916f
C994 CS_BIAS.n125 GND 0.007868f
C995 CS_BIAS.n126 GND 0.004243f
C996 CS_BIAS.n127 GND 0.004243f
C997 CS_BIAS.n128 GND 0.004243f
C998 CS_BIAS.n129 GND 0.007868f
C999 CS_BIAS.n130 GND 0.007868f
C1000 CS_BIAS.n131 GND 0.008428f
C1001 CS_BIAS.n132 GND 0.004243f
C1002 CS_BIAS.n133 GND 0.004243f
C1003 CS_BIAS.n134 GND 0.004243f
C1004 CS_BIAS.n135 GND 0.008344f
C1005 CS_BIAS.n136 GND 0.007868f
C1006 CS_BIAS.n137 GND 0.007868f
C1007 CS_BIAS.n138 GND 0.004243f
C1008 CS_BIAS.n139 GND 0.004243f
C1009 CS_BIAS.n140 GND 0.004243f
C1010 CS_BIAS.n141 GND 0.007868f
C1011 CS_BIAS.n142 GND 0.005072f
C1012 CS_BIAS.n143 GND 0.092263f
C1013 CS_BIAS.n144 GND 0.006781f
C1014 CS_BIAS.n145 GND 0.004243f
C1015 CS_BIAS.n146 GND 0.004243f
C1016 CS_BIAS.n147 GND 0.004243f
C1017 CS_BIAS.n148 GND 0.007868f
C1018 CS_BIAS.n149 GND 0.007868f
C1019 CS_BIAS.n150 GND 0.007868f
C1020 CS_BIAS.n151 GND 0.004243f
C1021 CS_BIAS.n152 GND 0.004243f
C1022 CS_BIAS.n153 GND 0.004243f
C1023 CS_BIAS.n154 GND 0.005933f
C1024 CS_BIAS.n155 GND 0.007868f
C1025 CS_BIAS.n156 GND 0.007868f
C1026 CS_BIAS.n157 GND 0.004243f
C1027 CS_BIAS.n158 GND 0.004243f
C1028 CS_BIAS.n159 GND 0.004243f
C1029 CS_BIAS.n160 GND 0.007868f
C1030 CS_BIAS.n161 GND 0.007092f
C1031 CS_BIAS.n162 GND 0.111655f
C1032 CS_BIAS.n163 GND 0.075496f
C1033 CS_BIAS.t15 GND 0.004918f
C1034 CS_BIAS.t21 GND 0.004918f
C1035 CS_BIAS.n164 GND 0.041084f
C1036 CS_BIAS.n165 GND 0.14918f
C1037 CS_BIAS.t23 GND 0.004918f
C1038 CS_BIAS.t13 GND 0.004918f
C1039 CS_BIAS.n166 GND 0.041084f
C1040 CS_BIAS.t17 GND 0.004918f
C1041 CS_BIAS.t11 GND 0.004918f
C1042 CS_BIAS.n167 GND 0.044879f
C1043 CS_BIAS.n168 GND 0.27761f
C1044 CS_BIAS.n169 GND 0.027501f
C1045 CS_BIAS.n170 GND 0.003707f
C1046 CS_BIAS.n171 GND 0.004243f
C1047 CS_BIAS.n172 GND 0.007868f
C1048 CS_BIAS.n173 GND 0.007868f
C1049 CS_BIAS.n174 GND 0.007868f
C1050 CS_BIAS.n175 GND 0.004243f
C1051 CS_BIAS.n176 GND 0.004243f
C1052 CS_BIAS.n177 GND 0.004243f
C1053 CS_BIAS.n178 GND 0.006936f
C1054 CS_BIAS.n179 GND 0.092263f
C1055 CS_BIAS.n180 GND 0.004916f
C1056 CS_BIAS.n181 GND 0.007868f
C1057 CS_BIAS.n182 GND 0.004243f
C1058 CS_BIAS.n183 GND 0.004243f
C1059 CS_BIAS.n184 GND 0.004243f
C1060 CS_BIAS.n185 GND 0.007868f
C1061 CS_BIAS.n186 GND 0.007868f
C1062 CS_BIAS.n187 GND 0.008428f
C1063 CS_BIAS.n188 GND 0.004243f
C1064 CS_BIAS.n189 GND 0.004243f
C1065 CS_BIAS.n190 GND 0.004243f
C1066 CS_BIAS.n191 GND 0.008344f
C1067 CS_BIAS.n192 GND 0.007868f
C1068 CS_BIAS.n193 GND 0.007868f
C1069 CS_BIAS.n194 GND 0.004243f
C1070 CS_BIAS.n195 GND 0.004243f
C1071 CS_BIAS.n196 GND 0.004243f
C1072 CS_BIAS.n197 GND 0.007868f
C1073 CS_BIAS.n198 GND 0.005072f
C1074 CS_BIAS.n199 GND 0.092263f
C1075 CS_BIAS.n200 GND 0.006781f
C1076 CS_BIAS.n201 GND 0.004243f
C1077 CS_BIAS.n202 GND 0.004243f
C1078 CS_BIAS.n203 GND 0.004243f
C1079 CS_BIAS.n204 GND 0.007868f
C1080 CS_BIAS.n205 GND 0.007868f
C1081 CS_BIAS.n206 GND 0.007868f
C1082 CS_BIAS.n207 GND 0.004243f
C1083 CS_BIAS.n208 GND 0.004243f
C1084 CS_BIAS.n209 GND 0.004243f
C1085 CS_BIAS.n210 GND 0.005933f
C1086 CS_BIAS.n211 GND 0.007868f
C1087 CS_BIAS.n212 GND 0.007868f
C1088 CS_BIAS.n213 GND 0.004243f
C1089 CS_BIAS.n214 GND 0.004243f
C1090 CS_BIAS.n215 GND 0.004243f
C1091 CS_BIAS.n216 GND 0.007868f
C1092 CS_BIAS.n217 GND 0.007092f
C1093 CS_BIAS.n218 GND 0.111655f
C1094 CS_BIAS.n219 GND 0.056208f
C1095 CS_BIAS.n220 GND 0.009829f
C1096 CS_BIAS.t27 GND 0.24163f
C1097 CS_BIAS.n221 GND 0.007868f
C1098 CS_BIAS.n222 GND 0.004243f
C1099 CS_BIAS.n223 GND 0.006403f
C1100 CS_BIAS.n224 GND 0.004243f
C1101 CS_BIAS.n225 GND 0.007868f
C1102 CS_BIAS.n226 GND 0.004243f
C1103 CS_BIAS.t35 GND 0.24163f
C1104 CS_BIAS.n227 GND 0.007868f
C1105 CS_BIAS.n228 GND 0.004243f
C1106 CS_BIAS.n229 GND 0.003432f
C1107 CS_BIAS.n230 GND 0.004243f
C1108 CS_BIAS.n231 GND 0.007868f
C1109 CS_BIAS.n232 GND 0.004243f
C1110 CS_BIAS.t39 GND 0.24163f
C1111 CS_BIAS.n233 GND 0.007868f
C1112 CS_BIAS.n234 GND 0.004243f
C1113 CS_BIAS.n235 GND 0.006168f
C1114 CS_BIAS.n236 GND 0.004243f
C1115 CS_BIAS.n237 GND 0.007868f
C1116 CS_BIAS.n238 GND 0.004243f
C1117 CS_BIAS.t46 GND 0.24163f
C1118 CS_BIAS.n239 GND 0.007868f
C1119 CS_BIAS.n240 GND 0.004243f
C1120 CS_BIAS.n241 GND 0.008428f
C1121 CS_BIAS.n242 GND 0.004243f
C1122 CS_BIAS.n243 GND 0.007868f
C1123 CS_BIAS.n244 GND 0.004243f
C1124 CS_BIAS.t31 GND 0.24163f
C1125 CS_BIAS.n245 GND 0.108683f
C1126 CS_BIAS.t37 GND 0.332306f
C1127 CS_BIAS.n246 GND 0.147952f
C1128 CS_BIAS.n247 GND 0.05348f
C1129 CS_BIAS.n248 GND 0.005072f
C1130 CS_BIAS.n249 GND 0.007868f
C1131 CS_BIAS.n250 GND 0.007868f
C1132 CS_BIAS.n251 GND 0.004243f
C1133 CS_BIAS.n252 GND 0.004243f
C1134 CS_BIAS.n253 GND 0.004243f
C1135 CS_BIAS.n254 GND 0.007868f
C1136 CS_BIAS.n255 GND 0.008344f
C1137 CS_BIAS.n256 GND 0.003432f
C1138 CS_BIAS.n257 GND 0.004243f
C1139 CS_BIAS.n258 GND 0.004243f
C1140 CS_BIAS.n259 GND 0.004243f
C1141 CS_BIAS.n260 GND 0.007868f
C1142 CS_BIAS.n261 GND 0.007868f
C1143 CS_BIAS.n262 GND 0.007868f
C1144 CS_BIAS.n263 GND 0.004243f
C1145 CS_BIAS.n264 GND 0.004243f
C1146 CS_BIAS.n265 GND 0.004243f
C1147 CS_BIAS.n266 GND 0.004916f
C1148 CS_BIAS.n267 GND 0.092263f
C1149 CS_BIAS.n268 GND 0.006936f
C1150 CS_BIAS.n269 GND 0.007868f
C1151 CS_BIAS.n270 GND 0.004243f
C1152 CS_BIAS.n271 GND 0.004243f
C1153 CS_BIAS.n272 GND 0.004243f
C1154 CS_BIAS.n273 GND 0.007868f
C1155 CS_BIAS.n274 GND 0.007868f
C1156 CS_BIAS.n275 GND 0.006168f
C1157 CS_BIAS.n276 GND 0.004243f
C1158 CS_BIAS.n277 GND 0.004243f
C1159 CS_BIAS.n278 GND 0.004243f
C1160 CS_BIAS.n279 GND 0.007868f
C1161 CS_BIAS.n280 GND 0.007868f
C1162 CS_BIAS.n281 GND 0.007868f
C1163 CS_BIAS.n282 GND 0.004243f
C1164 CS_BIAS.n283 GND 0.004243f
C1165 CS_BIAS.n284 GND 0.004243f
C1166 CS_BIAS.n285 GND 0.006936f
C1167 CS_BIAS.n286 GND 0.092263f
C1168 CS_BIAS.n287 GND 0.004916f
C1169 CS_BIAS.n288 GND 0.007868f
C1170 CS_BIAS.n289 GND 0.004243f
C1171 CS_BIAS.n290 GND 0.004243f
C1172 CS_BIAS.n291 GND 0.004243f
C1173 CS_BIAS.n292 GND 0.007868f
C1174 CS_BIAS.n293 GND 0.007868f
C1175 CS_BIAS.n294 GND 0.008428f
C1176 CS_BIAS.n295 GND 0.004243f
C1177 CS_BIAS.n296 GND 0.004243f
C1178 CS_BIAS.n297 GND 0.004243f
C1179 CS_BIAS.n298 GND 0.008344f
C1180 CS_BIAS.n299 GND 0.007868f
C1181 CS_BIAS.n300 GND 0.007868f
C1182 CS_BIAS.n301 GND 0.004243f
C1183 CS_BIAS.n302 GND 0.004243f
C1184 CS_BIAS.n303 GND 0.004243f
C1185 CS_BIAS.n304 GND 0.007868f
C1186 CS_BIAS.n305 GND 0.005072f
C1187 CS_BIAS.n306 GND 0.092263f
C1188 CS_BIAS.n307 GND 0.006781f
C1189 CS_BIAS.n308 GND 0.004243f
C1190 CS_BIAS.n309 GND 0.004243f
C1191 CS_BIAS.n310 GND 0.004243f
C1192 CS_BIAS.n311 GND 0.007868f
C1193 CS_BIAS.n312 GND 0.007868f
C1194 CS_BIAS.n313 GND 0.007868f
C1195 CS_BIAS.n314 GND 0.004243f
C1196 CS_BIAS.n315 GND 0.004243f
C1197 CS_BIAS.n316 GND 0.004243f
C1198 CS_BIAS.n317 GND 0.005933f
C1199 CS_BIAS.n318 GND 0.007868f
C1200 CS_BIAS.n319 GND 0.007868f
C1201 CS_BIAS.n320 GND 0.004243f
C1202 CS_BIAS.n321 GND 0.004243f
C1203 CS_BIAS.n322 GND 0.004243f
C1204 CS_BIAS.n323 GND 0.007868f
C1205 CS_BIAS.n324 GND 0.007092f
C1206 CS_BIAS.n325 GND 0.111655f
C1207 CS_BIAS.n326 GND 0.049171f
C1208 CS_BIAS.n327 GND 0.444953f
C1209 CS_BIAS.n328 GND 0.009829f
C1210 CS_BIAS.t28 GND 0.24163f
C1211 CS_BIAS.n329 GND 0.007868f
C1212 CS_BIAS.n330 GND 0.004243f
C1213 CS_BIAS.n331 GND 0.006403f
C1214 CS_BIAS.n332 GND 0.004243f
C1215 CS_BIAS.n333 GND 0.007868f
C1216 CS_BIAS.n334 GND 0.004243f
C1217 CS_BIAS.t38 GND 0.24163f
C1218 CS_BIAS.n335 GND 0.007868f
C1219 CS_BIAS.n336 GND 0.004243f
C1220 CS_BIAS.n337 GND 0.003432f
C1221 CS_BIAS.n338 GND 0.004243f
C1222 CS_BIAS.n339 GND 0.007868f
C1223 CS_BIAS.n340 GND 0.004243f
C1224 CS_BIAS.t24 GND 0.24163f
C1225 CS_BIAS.n341 GND 0.007868f
C1226 CS_BIAS.n342 GND 0.004243f
C1227 CS_BIAS.n343 GND 0.006168f
C1228 CS_BIAS.n344 GND 0.004243f
C1229 CS_BIAS.n345 GND 0.007868f
C1230 CS_BIAS.n346 GND 0.004243f
C1231 CS_BIAS.t43 GND 0.24163f
C1232 CS_BIAS.n347 GND 0.007868f
C1233 CS_BIAS.n348 GND 0.004243f
C1234 CS_BIAS.n349 GND 0.008428f
C1235 CS_BIAS.n350 GND 0.004243f
C1236 CS_BIAS.n351 GND 0.007868f
C1237 CS_BIAS.n352 GND 0.004243f
C1238 CS_BIAS.t47 GND 0.24163f
C1239 CS_BIAS.n353 GND 0.108683f
C1240 CS_BIAS.t34 GND 0.332306f
C1241 CS_BIAS.n354 GND 0.147952f
C1242 CS_BIAS.n355 GND 0.05348f
C1243 CS_BIAS.n356 GND 0.005072f
C1244 CS_BIAS.n357 GND 0.007868f
C1245 CS_BIAS.n358 GND 0.007868f
C1246 CS_BIAS.n359 GND 0.004243f
C1247 CS_BIAS.n360 GND 0.004243f
C1248 CS_BIAS.n361 GND 0.004243f
C1249 CS_BIAS.n362 GND 0.007868f
C1250 CS_BIAS.n363 GND 0.008344f
C1251 CS_BIAS.n364 GND 0.003432f
C1252 CS_BIAS.n365 GND 0.004243f
C1253 CS_BIAS.n366 GND 0.004243f
C1254 CS_BIAS.n367 GND 0.004243f
C1255 CS_BIAS.n368 GND 0.007868f
C1256 CS_BIAS.n369 GND 0.007868f
C1257 CS_BIAS.n370 GND 0.007868f
C1258 CS_BIAS.n371 GND 0.004243f
C1259 CS_BIAS.n372 GND 0.004243f
C1260 CS_BIAS.n373 GND 0.004243f
C1261 CS_BIAS.n374 GND 0.004916f
C1262 CS_BIAS.n375 GND 0.092263f
C1263 CS_BIAS.n376 GND 0.006936f
C1264 CS_BIAS.n377 GND 0.007868f
C1265 CS_BIAS.n378 GND 0.004243f
C1266 CS_BIAS.n379 GND 0.004243f
C1267 CS_BIAS.n380 GND 0.004243f
C1268 CS_BIAS.n381 GND 0.007868f
C1269 CS_BIAS.n382 GND 0.007868f
C1270 CS_BIAS.n383 GND 0.006168f
C1271 CS_BIAS.n384 GND 0.003707f
C1272 CS_BIAS.t3 GND 0.004918f
C1273 CS_BIAS.t19 GND 0.004918f
C1274 CS_BIAS.n385 GND 0.044879f
C1275 CS_BIAS.t5 GND 0.004918f
C1276 CS_BIAS.t7 GND 0.004918f
C1277 CS_BIAS.n386 GND 0.041084f
C1278 CS_BIAS.n387 GND 0.009829f
C1279 CS_BIAS.t8 GND 0.24163f
C1280 CS_BIAS.n388 GND 0.007868f
C1281 CS_BIAS.n389 GND 0.004243f
C1282 CS_BIAS.n390 GND 0.006403f
C1283 CS_BIAS.n391 GND 0.004243f
C1284 CS_BIAS.n392 GND 0.007868f
C1285 CS_BIAS.n393 GND 0.004243f
C1286 CS_BIAS.t0 GND 0.24163f
C1287 CS_BIAS.n394 GND 0.007868f
C1288 CS_BIAS.n395 GND 0.004243f
C1289 CS_BIAS.n396 GND 0.003432f
C1290 CS_BIAS.n397 GND 0.004243f
C1291 CS_BIAS.n398 GND 0.007868f
C1292 CS_BIAS.n399 GND 0.004243f
C1293 CS_BIAS.t6 GND 0.24163f
C1294 CS_BIAS.n400 GND 0.007868f
C1295 CS_BIAS.n401 GND 0.004243f
C1296 CS_BIAS.n402 GND 0.006168f
C1297 CS_BIAS.n403 GND 0.004243f
C1298 CS_BIAS.n404 GND 0.007868f
C1299 CS_BIAS.n405 GND 0.004243f
C1300 CS_BIAS.t4 GND 0.24163f
C1301 CS_BIAS.n406 GND 0.007868f
C1302 CS_BIAS.n407 GND 0.004243f
C1303 CS_BIAS.n408 GND 0.008428f
C1304 CS_BIAS.n409 GND 0.004243f
C1305 CS_BIAS.n410 GND 0.007868f
C1306 CS_BIAS.n411 GND 0.004243f
C1307 CS_BIAS.t18 GND 0.24163f
C1308 CS_BIAS.n412 GND 0.108683f
C1309 CS_BIAS.t2 GND 0.332306f
C1310 CS_BIAS.n413 GND 0.147952f
C1311 CS_BIAS.n414 GND 0.05348f
C1312 CS_BIAS.n415 GND 0.005072f
C1313 CS_BIAS.n416 GND 0.007868f
C1314 CS_BIAS.n417 GND 0.007868f
C1315 CS_BIAS.n418 GND 0.004243f
C1316 CS_BIAS.n419 GND 0.004243f
C1317 CS_BIAS.n420 GND 0.004243f
C1318 CS_BIAS.n421 GND 0.007868f
C1319 CS_BIAS.n422 GND 0.008344f
C1320 CS_BIAS.n423 GND 0.003432f
C1321 CS_BIAS.n424 GND 0.004243f
C1322 CS_BIAS.n425 GND 0.004243f
C1323 CS_BIAS.n426 GND 0.004243f
C1324 CS_BIAS.n427 GND 0.007868f
C1325 CS_BIAS.n428 GND 0.007868f
C1326 CS_BIAS.n429 GND 0.007868f
C1327 CS_BIAS.n430 GND 0.004243f
C1328 CS_BIAS.n431 GND 0.004243f
C1329 CS_BIAS.n432 GND 0.004243f
C1330 CS_BIAS.n433 GND 0.004916f
C1331 CS_BIAS.n434 GND 0.092263f
C1332 CS_BIAS.n435 GND 0.006936f
C1333 CS_BIAS.n436 GND 0.007868f
C1334 CS_BIAS.n437 GND 0.004243f
C1335 CS_BIAS.n438 GND 0.004243f
C1336 CS_BIAS.n439 GND 0.004243f
C1337 CS_BIAS.n440 GND 0.007868f
C1338 CS_BIAS.n441 GND 0.007868f
C1339 CS_BIAS.n442 GND 0.006168f
C1340 CS_BIAS.n443 GND 0.004243f
C1341 CS_BIAS.n444 GND 0.004243f
C1342 CS_BIAS.n445 GND 0.004243f
C1343 CS_BIAS.n446 GND 0.007868f
C1344 CS_BIAS.n447 GND 0.007868f
C1345 CS_BIAS.n448 GND 0.007868f
C1346 CS_BIAS.n449 GND 0.004243f
C1347 CS_BIAS.n450 GND 0.004243f
C1348 CS_BIAS.n451 GND 0.004243f
C1349 CS_BIAS.n452 GND 0.006936f
C1350 CS_BIAS.n453 GND 0.092263f
C1351 CS_BIAS.n454 GND 0.004916f
C1352 CS_BIAS.n455 GND 0.007868f
C1353 CS_BIAS.n456 GND 0.004243f
C1354 CS_BIAS.n457 GND 0.004243f
C1355 CS_BIAS.n458 GND 0.004243f
C1356 CS_BIAS.n459 GND 0.007868f
C1357 CS_BIAS.n460 GND 0.007868f
C1358 CS_BIAS.n461 GND 0.008428f
C1359 CS_BIAS.n462 GND 0.004243f
C1360 CS_BIAS.n463 GND 0.004243f
C1361 CS_BIAS.n464 GND 0.004243f
C1362 CS_BIAS.n465 GND 0.008344f
C1363 CS_BIAS.n466 GND 0.007868f
C1364 CS_BIAS.n467 GND 0.007868f
C1365 CS_BIAS.n468 GND 0.004243f
C1366 CS_BIAS.n469 GND 0.004243f
C1367 CS_BIAS.n470 GND 0.004243f
C1368 CS_BIAS.n471 GND 0.007868f
C1369 CS_BIAS.n472 GND 0.005072f
C1370 CS_BIAS.n473 GND 0.092263f
C1371 CS_BIAS.n474 GND 0.006781f
C1372 CS_BIAS.n475 GND 0.004243f
C1373 CS_BIAS.n476 GND 0.004243f
C1374 CS_BIAS.n477 GND 0.004243f
C1375 CS_BIAS.n478 GND 0.007868f
C1376 CS_BIAS.n479 GND 0.007868f
C1377 CS_BIAS.n480 GND 0.007868f
C1378 CS_BIAS.n481 GND 0.004243f
C1379 CS_BIAS.n482 GND 0.004243f
C1380 CS_BIAS.n483 GND 0.004243f
C1381 CS_BIAS.n484 GND 0.005933f
C1382 CS_BIAS.n485 GND 0.007868f
C1383 CS_BIAS.n486 GND 0.007868f
C1384 CS_BIAS.n487 GND 0.004243f
C1385 CS_BIAS.n488 GND 0.004243f
C1386 CS_BIAS.n489 GND 0.004243f
C1387 CS_BIAS.n490 GND 0.007868f
C1388 CS_BIAS.n491 GND 0.007092f
C1389 CS_BIAS.n492 GND 0.111655f
C1390 CS_BIAS.n493 GND 0.075496f
C1391 CS_BIAS.t1 GND 0.004918f
C1392 CS_BIAS.t9 GND 0.004918f
C1393 CS_BIAS.n494 GND 0.041084f
C1394 CS_BIAS.n495 GND 0.14918f
C1395 CS_BIAS.n496 GND 0.27761f
C1396 CS_BIAS.n497 GND 0.027501f
C1397 CS_BIAS.n498 GND 0.003707f
C1398 CS_BIAS.n499 GND 0.004243f
C1399 CS_BIAS.n500 GND 0.007868f
C1400 CS_BIAS.n501 GND 0.007868f
C1401 CS_BIAS.n502 GND 0.007868f
C1402 CS_BIAS.n503 GND 0.004243f
C1403 CS_BIAS.n504 GND 0.004243f
C1404 CS_BIAS.n505 GND 0.004243f
C1405 CS_BIAS.n506 GND 0.006936f
C1406 CS_BIAS.n507 GND 0.092263f
C1407 CS_BIAS.n508 GND 0.004916f
C1408 CS_BIAS.n509 GND 0.007868f
C1409 CS_BIAS.n510 GND 0.004243f
C1410 CS_BIAS.n511 GND 0.004243f
C1411 CS_BIAS.n512 GND 0.004243f
C1412 CS_BIAS.n513 GND 0.007868f
C1413 CS_BIAS.n514 GND 0.007868f
C1414 CS_BIAS.n515 GND 0.008428f
C1415 CS_BIAS.n516 GND 0.004243f
C1416 CS_BIAS.n517 GND 0.004243f
C1417 CS_BIAS.n518 GND 0.004243f
C1418 CS_BIAS.n519 GND 0.008344f
C1419 CS_BIAS.n520 GND 0.007868f
C1420 CS_BIAS.n521 GND 0.007868f
C1421 CS_BIAS.n522 GND 0.004243f
C1422 CS_BIAS.n523 GND 0.004243f
C1423 CS_BIAS.n524 GND 0.004243f
C1424 CS_BIAS.n525 GND 0.007868f
C1425 CS_BIAS.n526 GND 0.005072f
C1426 CS_BIAS.n527 GND 0.092263f
C1427 CS_BIAS.n528 GND 0.006781f
C1428 CS_BIAS.n529 GND 0.004243f
C1429 CS_BIAS.n530 GND 0.004243f
C1430 CS_BIAS.n531 GND 0.004243f
C1431 CS_BIAS.n532 GND 0.007868f
C1432 CS_BIAS.n533 GND 0.007868f
C1433 CS_BIAS.n534 GND 0.007868f
C1434 CS_BIAS.n535 GND 0.004243f
C1435 CS_BIAS.n536 GND 0.004243f
C1436 CS_BIAS.n537 GND 0.004243f
C1437 CS_BIAS.n538 GND 0.005933f
C1438 CS_BIAS.n539 GND 0.007868f
C1439 CS_BIAS.n540 GND 0.007868f
C1440 CS_BIAS.n541 GND 0.004243f
C1441 CS_BIAS.n542 GND 0.004243f
C1442 CS_BIAS.n543 GND 0.004243f
C1443 CS_BIAS.n544 GND 0.007868f
C1444 CS_BIAS.n545 GND 0.007092f
C1445 CS_BIAS.n546 GND 0.111655f
C1446 CS_BIAS.n547 GND 0.056208f
C1447 CS_BIAS.n548 GND 0.009829f
C1448 CS_BIAS.t40 GND 0.24163f
C1449 CS_BIAS.n549 GND 0.007868f
C1450 CS_BIAS.n550 GND 0.004243f
C1451 CS_BIAS.n551 GND 0.006403f
C1452 CS_BIAS.n552 GND 0.004243f
C1453 CS_BIAS.n553 GND 0.007868f
C1454 CS_BIAS.n554 GND 0.004243f
C1455 CS_BIAS.t45 GND 0.24163f
C1456 CS_BIAS.n555 GND 0.007868f
C1457 CS_BIAS.n556 GND 0.004243f
C1458 CS_BIAS.n557 GND 0.003432f
C1459 CS_BIAS.n558 GND 0.004243f
C1460 CS_BIAS.n559 GND 0.007868f
C1461 CS_BIAS.n560 GND 0.004243f
C1462 CS_BIAS.t32 GND 0.24163f
C1463 CS_BIAS.n561 GND 0.007868f
C1464 CS_BIAS.n562 GND 0.004243f
C1465 CS_BIAS.n563 GND 0.006168f
C1466 CS_BIAS.n564 GND 0.004243f
C1467 CS_BIAS.n565 GND 0.007868f
C1468 CS_BIAS.n566 GND 0.004243f
C1469 CS_BIAS.t30 GND 0.24163f
C1470 CS_BIAS.n567 GND 0.007868f
C1471 CS_BIAS.n568 GND 0.004243f
C1472 CS_BIAS.n569 GND 0.008428f
C1473 CS_BIAS.n570 GND 0.004243f
C1474 CS_BIAS.n571 GND 0.007868f
C1475 CS_BIAS.n572 GND 0.004243f
C1476 CS_BIAS.t44 GND 0.24163f
C1477 CS_BIAS.n573 GND 0.108683f
C1478 CS_BIAS.t25 GND 0.332306f
C1479 CS_BIAS.n574 GND 0.147952f
C1480 CS_BIAS.n575 GND 0.05348f
C1481 CS_BIAS.n576 GND 0.005072f
C1482 CS_BIAS.n577 GND 0.007868f
C1483 CS_BIAS.n578 GND 0.007868f
C1484 CS_BIAS.n579 GND 0.004243f
C1485 CS_BIAS.n580 GND 0.004243f
C1486 CS_BIAS.n581 GND 0.004243f
C1487 CS_BIAS.n582 GND 0.007868f
C1488 CS_BIAS.n583 GND 0.008344f
C1489 CS_BIAS.n584 GND 0.003432f
C1490 CS_BIAS.n585 GND 0.004243f
C1491 CS_BIAS.n586 GND 0.004243f
C1492 CS_BIAS.n587 GND 0.004243f
C1493 CS_BIAS.n588 GND 0.007868f
C1494 CS_BIAS.n589 GND 0.007868f
C1495 CS_BIAS.n590 GND 0.007868f
C1496 CS_BIAS.n591 GND 0.004243f
C1497 CS_BIAS.n592 GND 0.004243f
C1498 CS_BIAS.n593 GND 0.004243f
C1499 CS_BIAS.n594 GND 0.004916f
C1500 CS_BIAS.n595 GND 0.092263f
C1501 CS_BIAS.n596 GND 0.006936f
C1502 CS_BIAS.n597 GND 0.007868f
C1503 CS_BIAS.n598 GND 0.004243f
C1504 CS_BIAS.n599 GND 0.004243f
C1505 CS_BIAS.n600 GND 0.004243f
C1506 CS_BIAS.n601 GND 0.007868f
C1507 CS_BIAS.n602 GND 0.007868f
C1508 CS_BIAS.n603 GND 0.006168f
C1509 CS_BIAS.n604 GND 0.004243f
C1510 CS_BIAS.n605 GND 0.004243f
C1511 CS_BIAS.n606 GND 0.004243f
C1512 CS_BIAS.n607 GND 0.007868f
C1513 CS_BIAS.n608 GND 0.007868f
C1514 CS_BIAS.n609 GND 0.007868f
C1515 CS_BIAS.n610 GND 0.004243f
C1516 CS_BIAS.n611 GND 0.004243f
C1517 CS_BIAS.n612 GND 0.004243f
C1518 CS_BIAS.n613 GND 0.006936f
C1519 CS_BIAS.n614 GND 0.092263f
C1520 CS_BIAS.n615 GND 0.004916f
C1521 CS_BIAS.n616 GND 0.007868f
C1522 CS_BIAS.n617 GND 0.004243f
C1523 CS_BIAS.n618 GND 0.004243f
C1524 CS_BIAS.n619 GND 0.004243f
C1525 CS_BIAS.n620 GND 0.007868f
C1526 CS_BIAS.n621 GND 0.007868f
C1527 CS_BIAS.n622 GND 0.008428f
C1528 CS_BIAS.n623 GND 0.004243f
C1529 CS_BIAS.n624 GND 0.004243f
C1530 CS_BIAS.n625 GND 0.004243f
C1531 CS_BIAS.n626 GND 0.008344f
C1532 CS_BIAS.n627 GND 0.007868f
C1533 CS_BIAS.n628 GND 0.007868f
C1534 CS_BIAS.n629 GND 0.004243f
C1535 CS_BIAS.n630 GND 0.004243f
C1536 CS_BIAS.n631 GND 0.004243f
C1537 CS_BIAS.n632 GND 0.007868f
C1538 CS_BIAS.n633 GND 0.005072f
C1539 CS_BIAS.n634 GND 0.092263f
C1540 CS_BIAS.n635 GND 0.006781f
C1541 CS_BIAS.n636 GND 0.004243f
C1542 CS_BIAS.n637 GND 0.004243f
C1543 CS_BIAS.n638 GND 0.004243f
C1544 CS_BIAS.n639 GND 0.007868f
C1545 CS_BIAS.n640 GND 0.007868f
C1546 CS_BIAS.n641 GND 0.007868f
C1547 CS_BIAS.n642 GND 0.004243f
C1548 CS_BIAS.n643 GND 0.004243f
C1549 CS_BIAS.n644 GND 0.004243f
C1550 CS_BIAS.n645 GND 0.005933f
C1551 CS_BIAS.n646 GND 0.007868f
C1552 CS_BIAS.n647 GND 0.007868f
C1553 CS_BIAS.n648 GND 0.004243f
C1554 CS_BIAS.n649 GND 0.004243f
C1555 CS_BIAS.n650 GND 0.004243f
C1556 CS_BIAS.n651 GND 0.007868f
C1557 CS_BIAS.n652 GND 0.007092f
C1558 CS_BIAS.n653 GND 0.111655f
C1559 CS_BIAS.n654 GND 0.049171f
C1560 CS_BIAS.n655 GND 0.103965f
C1561 CS_BIAS.n656 GND 3.5423f
C1562 VDD.t29 GND 0.010687f
C1563 VDD.t3 GND 0.010687f
C1564 VDD.n0 GND 0.072846f
C1565 VDD.t131 GND 0.010687f
C1566 VDD.t44 GND 0.010687f
C1567 VDD.n1 GND 0.069897f
C1568 VDD.n2 GND 0.418977f
C1569 VDD.t135 GND 0.010687f
C1570 VDD.t1 GND 0.010687f
C1571 VDD.n3 GND 0.069897f
C1572 VDD.n4 GND 0.21953f
C1573 VDD.t62 GND 0.010687f
C1574 VDD.t58 GND 0.010687f
C1575 VDD.n5 GND 0.069897f
C1576 VDD.n6 GND 0.183156f
C1577 VDD.t13 GND 0.010687f
C1578 VDD.t10 GND 0.010687f
C1579 VDD.n7 GND 0.072846f
C1580 VDD.t20 GND 0.010687f
C1581 VDD.t60 GND 0.010687f
C1582 VDD.n8 GND 0.069897f
C1583 VDD.n9 GND 0.418977f
C1584 VDD.t137 GND 0.010687f
C1585 VDD.t31 GND 0.010687f
C1586 VDD.n10 GND 0.069897f
C1587 VDD.n11 GND 0.21953f
C1588 VDD.t41 GND 0.010687f
C1589 VDD.t34 GND 0.010687f
C1590 VDD.n12 GND 0.069897f
C1591 VDD.n13 GND 0.183156f
C1592 VDD.n14 GND 0.138091f
C1593 VDD.n15 GND 2.52461f
C1594 VDD.t38 GND 0.012824f
C1595 VDD.t51 GND 0.012824f
C1596 VDD.n16 GND 0.080827f
C1597 VDD.t66 GND 0.012824f
C1598 VDD.t24 GND 0.012824f
C1599 VDD.n17 GND 0.07391f
C1600 VDD.n18 GND 0.514737f
C1601 VDD.t49 GND 0.012824f
C1602 VDD.t6 GND 0.012824f
C1603 VDD.n19 GND 0.07391f
C1604 VDD.n20 GND 0.259498f
C1605 VDD.t46 GND 0.102273f
C1606 VDD.n21 GND 0.203917f
C1607 VDD.t39 GND 0.012824f
C1608 VDD.t56 GND 0.012824f
C1609 VDD.n22 GND 0.080827f
C1610 VDD.t48 GND 0.012824f
C1611 VDD.t65 GND 0.012824f
C1612 VDD.n23 GND 0.07391f
C1613 VDD.n24 GND 0.514737f
C1614 VDD.t18 GND 0.012824f
C1615 VDD.t35 GND 0.012824f
C1616 VDD.n25 GND 0.07391f
C1617 VDD.n26 GND 0.259498f
C1618 VDD.t8 GND 0.102273f
C1619 VDD.n27 GND 0.184098f
C1620 VDD.n28 GND 0.35869f
C1621 VDD.n29 GND 0.006454f
C1622 VDD.n30 GND 0.006454f
C1623 VDD.n31 GND 0.005213f
C1624 VDD.n32 GND 0.005213f
C1625 VDD.n33 GND 0.006477f
C1626 VDD.n34 GND 0.006477f
C1627 VDD.n35 GND 0.429674f
C1628 VDD.n36 GND 0.006477f
C1629 VDD.n37 GND 0.006477f
C1630 VDD.n38 GND 0.006477f
C1631 VDD.n39 GND 0.429674f
C1632 VDD.n40 GND 0.006477f
C1633 VDD.n41 GND 0.006477f
C1634 VDD.n42 GND 0.006477f
C1635 VDD.n43 GND 0.006477f
C1636 VDD.n44 GND 0.005213f
C1637 VDD.n45 GND 0.006477f
C1638 VDD.n46 GND 0.006477f
C1639 VDD.n47 GND 0.006477f
C1640 VDD.n48 GND 0.006477f
C1641 VDD.n49 GND 0.429674f
C1642 VDD.n50 GND 0.006477f
C1643 VDD.n51 GND 0.006477f
C1644 VDD.n52 GND 0.006477f
C1645 VDD.n53 GND 0.006477f
C1646 VDD.n54 GND 0.006477f
C1647 VDD.n55 GND 0.005213f
C1648 VDD.n56 GND 0.006477f
C1649 VDD.n57 GND 0.006477f
C1650 VDD.n58 GND 0.006477f
C1651 VDD.n59 GND 0.006477f
C1652 VDD.n60 GND 0.266398f
C1653 VDD.n61 GND 0.006477f
C1654 VDD.n62 GND 0.006477f
C1655 VDD.n63 GND 0.006477f
C1656 VDD.n64 GND 0.006477f
C1657 VDD.n65 GND 0.006477f
C1658 VDD.n66 GND 0.005213f
C1659 VDD.n67 GND 0.006477f
C1660 VDD.t17 GND 0.214837f
C1661 VDD.n68 GND 0.006477f
C1662 VDD.n69 GND 0.006477f
C1663 VDD.n70 GND 0.006477f
C1664 VDD.n71 GND 0.429674f
C1665 VDD.n72 GND 0.006477f
C1666 VDD.n73 GND 0.006477f
C1667 VDD.n74 GND 0.006477f
C1668 VDD.n75 GND 0.006477f
C1669 VDD.n76 GND 0.006477f
C1670 VDD.n77 GND 0.005213f
C1671 VDD.n78 GND 0.006477f
C1672 VDD.n79 GND 0.006477f
C1673 VDD.n80 GND 0.006477f
C1674 VDD.n81 GND 0.006477f
C1675 VDD.n82 GND 0.429674f
C1676 VDD.n83 GND 0.006477f
C1677 VDD.n84 GND 0.006477f
C1678 VDD.n85 GND 0.006477f
C1679 VDD.n86 GND 0.006477f
C1680 VDD.n87 GND 0.006477f
C1681 VDD.n88 GND 0.005213f
C1682 VDD.n89 GND 0.006477f
C1683 VDD.n90 GND 0.006477f
C1684 VDD.n91 GND 0.006477f
C1685 VDD.n92 GND 0.006477f
C1686 VDD.t5 GND 0.214837f
C1687 VDD.n93 GND 0.006477f
C1688 VDD.n94 GND 0.006477f
C1689 VDD.n95 GND 0.006477f
C1690 VDD.n96 GND 0.006477f
C1691 VDD.n97 GND 0.006477f
C1692 VDD.n98 GND 0.005213f
C1693 VDD.n99 GND 0.006477f
C1694 VDD.n100 GND 0.326552f
C1695 VDD.n101 GND 0.006477f
C1696 VDD.n102 GND 0.006477f
C1697 VDD.n103 GND 0.006477f
C1698 VDD.n104 GND 0.429674f
C1699 VDD.n105 GND 0.006477f
C1700 VDD.n106 GND 0.006477f
C1701 VDD.n107 GND 0.006477f
C1702 VDD.n108 GND 0.006477f
C1703 VDD.n109 GND 0.006477f
C1704 VDD.n110 GND 0.005213f
C1705 VDD.n111 GND 0.006477f
C1706 VDD.n112 GND 0.006477f
C1707 VDD.n113 GND 0.006477f
C1708 VDD.n114 GND 0.006477f
C1709 VDD.n115 GND 0.429674f
C1710 VDD.n116 GND 0.006477f
C1711 VDD.n117 GND 0.006477f
C1712 VDD.n118 GND 0.006477f
C1713 VDD.n119 GND 0.006477f
C1714 VDD.n120 GND 0.006477f
C1715 VDD.n121 GND 0.005213f
C1716 VDD.n122 GND 0.006477f
C1717 VDD.n123 GND 0.006477f
C1718 VDD.n124 GND 0.006477f
C1719 VDD.n125 GND 0.006477f
C1720 VDD.n126 GND 0.429674f
C1721 VDD.n127 GND 0.006477f
C1722 VDD.n128 GND 0.006477f
C1723 VDD.n129 GND 0.006477f
C1724 VDD.n130 GND 0.006477f
C1725 VDD.n131 GND 0.006477f
C1726 VDD.n132 GND 0.005213f
C1727 VDD.n133 GND 0.006477f
C1728 VDD.n134 GND 0.006477f
C1729 VDD.n135 GND 0.006477f
C1730 VDD.n136 GND 0.006477f
C1731 VDD.n137 GND 0.429674f
C1732 VDD.n138 GND 0.006477f
C1733 VDD.n139 GND 0.006477f
C1734 VDD.n140 GND 0.006477f
C1735 VDD.n141 GND 0.006477f
C1736 VDD.n142 GND 0.006477f
C1737 VDD.n143 GND 0.005213f
C1738 VDD.n144 GND 0.006477f
C1739 VDD.n145 GND 0.006477f
C1740 VDD.n146 GND 0.006477f
C1741 VDD.n147 GND 0.006477f
C1742 VDD.n148 GND 0.429674f
C1743 VDD.n149 GND 0.006477f
C1744 VDD.n150 GND 0.006477f
C1745 VDD.n151 GND 0.006477f
C1746 VDD.n152 GND 0.006477f
C1747 VDD.n153 GND 0.006477f
C1748 VDD.n154 GND 0.005213f
C1749 VDD.n155 GND 0.006477f
C1750 VDD.n156 GND 0.006477f
C1751 VDD.n157 GND 0.006477f
C1752 VDD.n158 GND 0.006477f
C1753 VDD.n159 GND 0.244914f
C1754 VDD.n160 GND 0.006477f
C1755 VDD.n161 GND 0.006477f
C1756 VDD.n162 GND 0.006477f
C1757 VDD.n163 GND 0.006477f
C1758 VDD.n164 GND 0.006477f
C1759 VDD.n165 GND 0.005213f
C1760 VDD.n166 GND 0.006477f
C1761 VDD.t104 GND 0.214837f
C1762 VDD.n167 GND 0.006477f
C1763 VDD.n168 GND 0.006477f
C1764 VDD.n169 GND 0.006477f
C1765 VDD.n170 GND 0.429674f
C1766 VDD.n171 GND 0.006477f
C1767 VDD.n172 GND 0.006477f
C1768 VDD.n173 GND 0.006477f
C1769 VDD.n174 GND 0.006477f
C1770 VDD.n175 GND 0.006477f
C1771 VDD.n176 GND 0.004327f
C1772 VDD.n177 GND 0.014826f
C1773 VDD.n178 GND 0.006477f
C1774 VDD.n179 GND 0.014826f
C1775 VDD.n194 GND 0.006477f
C1776 VDD.t125 GND 0.086094f
C1777 VDD.t124 GND 0.107631f
C1778 VDD.t123 GND 0.799934f
C1779 VDD.n195 GND 0.078348f
C1780 VDD.n196 GND 0.048083f
C1781 VDD.n197 GND 0.008028f
C1782 VDD.n198 GND 0.006477f
C1783 VDD.n199 GND 0.005213f
C1784 VDD.n200 GND 0.006477f
C1785 VDD.n201 GND 0.005213f
C1786 VDD.n202 GND 0.006477f
C1787 VDD.n203 GND 0.005213f
C1788 VDD.n204 GND 0.006477f
C1789 VDD.t106 GND 0.086094f
C1790 VDD.t105 GND 0.107631f
C1791 VDD.t103 GND 0.799934f
C1792 VDD.n205 GND 0.078348f
C1793 VDD.n206 GND 0.048083f
C1794 VDD.n207 GND 0.010634f
C1795 VDD.n208 GND 0.006477f
C1796 VDD.n209 GND 0.005213f
C1797 VDD.n210 GND 0.006477f
C1798 VDD.n211 GND 0.005213f
C1799 VDD.n212 GND 0.006477f
C1800 VDD.n213 GND 0.005213f
C1801 VDD.n214 GND 0.014826f
C1802 VDD.n215 GND 0.014967f
C1803 VDD.n216 GND 0.004327f
C1804 VDD.n217 GND 0.014967f
C1805 VDD.n218 GND 0.006477f
C1806 VDD.n219 GND 0.006477f
C1807 VDD.n220 GND 0.006477f
C1808 VDD.n221 GND 0.006477f
C1809 VDD.n222 GND 0.005213f
C1810 VDD.n223 GND 0.005213f
C1811 VDD.n224 GND 0.006477f
C1812 VDD.n225 GND 0.006477f
C1813 VDD.n226 GND 0.005213f
C1814 VDD.n227 GND 0.006477f
C1815 VDD.n228 GND 0.006477f
C1816 VDD.n229 GND 0.006477f
C1817 VDD.n230 GND 0.006477f
C1818 VDD.n231 GND 0.006477f
C1819 VDD.n232 GND 0.005213f
C1820 VDD.n233 GND 0.005213f
C1821 VDD.n234 GND 0.006477f
C1822 VDD.n235 GND 0.006477f
C1823 VDD.n236 GND 0.005213f
C1824 VDD.n237 GND 0.006477f
C1825 VDD.n238 GND 0.006477f
C1826 VDD.n239 GND 0.006477f
C1827 VDD.n240 GND 0.006477f
C1828 VDD.n241 GND 0.006477f
C1829 VDD.n242 GND 0.005213f
C1830 VDD.n243 GND 0.005213f
C1831 VDD.n244 GND 0.006477f
C1832 VDD.n245 GND 0.006477f
C1833 VDD.n246 GND 0.003962f
C1834 VDD.n247 GND 0.006477f
C1835 VDD.n248 GND 0.006477f
C1836 VDD.n249 GND 0.006477f
C1837 VDD.n250 GND 0.006477f
C1838 VDD.n251 GND 0.006477f
C1839 VDD.n252 GND 0.004744f
C1840 VDD.n253 GND 0.005213f
C1841 VDD.n254 GND 0.006477f
C1842 VDD.n255 GND 0.006477f
C1843 VDD.n256 GND 0.005213f
C1844 VDD.n257 GND 0.006477f
C1845 VDD.n258 GND 0.006477f
C1846 VDD.n259 GND 0.006477f
C1847 VDD.n260 GND 0.006477f
C1848 VDD.n261 GND 0.006477f
C1849 VDD.n262 GND 0.005213f
C1850 VDD.n263 GND 0.005213f
C1851 VDD.n264 GND 0.006477f
C1852 VDD.n265 GND 0.006477f
C1853 VDD.n266 GND 0.005213f
C1854 VDD.n267 GND 0.006477f
C1855 VDD.n268 GND 0.006477f
C1856 VDD.n269 GND 0.006477f
C1857 VDD.n270 GND 0.006477f
C1858 VDD.n271 GND 0.006477f
C1859 VDD.n272 GND 0.005213f
C1860 VDD.n273 GND 0.005213f
C1861 VDD.n274 GND 0.006477f
C1862 VDD.n275 GND 0.006477f
C1863 VDD.n276 GND 0.005213f
C1864 VDD.n277 GND 0.006477f
C1865 VDD.n278 GND 0.006477f
C1866 VDD.n279 GND 0.006477f
C1867 VDD.n280 GND 0.006477f
C1868 VDD.n281 GND 0.006477f
C1869 VDD.n282 GND 0.005213f
C1870 VDD.n283 GND 0.006477f
C1871 VDD.n284 GND 0.005213f
C1872 VDD.n285 GND 0.002711f
C1873 VDD.n286 GND 0.006477f
C1874 VDD.n287 GND 0.006477f
C1875 VDD.n288 GND 0.005213f
C1876 VDD.n289 GND 0.006477f
C1877 VDD.n290 GND 0.005213f
C1878 VDD.n291 GND 0.006477f
C1879 VDD.n292 GND 0.005213f
C1880 VDD.n293 GND 0.006477f
C1881 VDD.n294 GND 0.005213f
C1882 VDD.n295 GND 0.006477f
C1883 VDD.n296 GND 0.005213f
C1884 VDD.n297 GND 0.006477f
C1885 VDD.n298 GND 0.005213f
C1886 VDD.n299 GND 0.006477f
C1887 VDD.n300 GND 0.005213f
C1888 VDD.n301 GND 0.006477f
C1889 VDD.n302 GND 0.005213f
C1890 VDD.n303 GND 0.006477f
C1891 VDD.n304 GND 0.005213f
C1892 VDD.n305 GND 0.006477f
C1893 VDD.n306 GND 0.005213f
C1894 VDD.n307 GND 0.006477f
C1895 VDD.n308 GND 0.005213f
C1896 VDD.n309 GND 0.006477f
C1897 VDD.n310 GND 0.005213f
C1898 VDD.n311 GND 0.006477f
C1899 VDD.n312 GND 0.005213f
C1900 VDD.n313 GND 0.006477f
C1901 VDD.n314 GND 0.005213f
C1902 VDD.n315 GND 0.006477f
C1903 VDD.n316 GND 0.006477f
C1904 VDD.n317 GND 0.429674f
C1905 VDD.n318 GND 0.006477f
C1906 VDD.n319 GND 0.005213f
C1907 VDD.n320 GND 0.006477f
C1908 VDD.n321 GND 0.005213f
C1909 VDD.n322 GND 0.006477f
C1910 VDD.n323 GND 0.429674f
C1911 VDD.n324 GND 0.006477f
C1912 VDD.n325 GND 0.005213f
C1913 VDD.n326 GND 0.006477f
C1914 VDD.n327 GND 0.005213f
C1915 VDD.n328 GND 0.006477f
C1916 VDD.n329 GND 0.429674f
C1917 VDD.n330 GND 0.006477f
C1918 VDD.n331 GND 0.005213f
C1919 VDD.n332 GND 0.006477f
C1920 VDD.n333 GND 0.005213f
C1921 VDD.n334 GND 0.006477f
C1922 VDD.n335 GND 0.429674f
C1923 VDD.n336 GND 0.006477f
C1924 VDD.n337 GND 0.005213f
C1925 VDD.n338 GND 0.006477f
C1926 VDD.n339 GND 0.005213f
C1927 VDD.n340 GND 0.006477f
C1928 VDD.n341 GND 0.266398f
C1929 VDD.n342 GND 0.006477f
C1930 VDD.n343 GND 0.005213f
C1931 VDD.n344 GND 0.006477f
C1932 VDD.n345 GND 0.005213f
C1933 VDD.n346 GND 0.006477f
C1934 VDD.n347 GND 0.429674f
C1935 VDD.n348 GND 0.006477f
C1936 VDD.n349 GND 0.005213f
C1937 VDD.n350 GND 0.006477f
C1938 VDD.n351 GND 0.005213f
C1939 VDD.n352 GND 0.006477f
C1940 VDD.n353 GND 0.429674f
C1941 VDD.n354 GND 0.006477f
C1942 VDD.n355 GND 0.005213f
C1943 VDD.n356 GND 0.006477f
C1944 VDD.n357 GND 0.005213f
C1945 VDD.n358 GND 0.006477f
C1946 VDD.n359 GND 0.429674f
C1947 VDD.n360 GND 0.006477f
C1948 VDD.n361 GND 0.005213f
C1949 VDD.n362 GND 0.006477f
C1950 VDD.n363 GND 0.005213f
C1951 VDD.n364 GND 0.006477f
C1952 VDD.n365 GND 0.429674f
C1953 VDD.n366 GND 0.006477f
C1954 VDD.n367 GND 0.005213f
C1955 VDD.n368 GND 0.006477f
C1956 VDD.n369 GND 0.005213f
C1957 VDD.n370 GND 0.006477f
C1958 VDD.n371 GND 0.429674f
C1959 VDD.n372 GND 0.006477f
C1960 VDD.n373 GND 0.005213f
C1961 VDD.n374 GND 0.006477f
C1962 VDD.n375 GND 0.005213f
C1963 VDD.n376 GND 0.006477f
C1964 VDD.t50 GND 0.214837f
C1965 VDD.n377 GND 0.006477f
C1966 VDD.n378 GND 0.005213f
C1967 VDD.n379 GND 0.006477f
C1968 VDD.n380 GND 0.005213f
C1969 VDD.n381 GND 0.006477f
C1970 VDD.n382 GND 0.429674f
C1971 VDD.n383 GND 0.006477f
C1972 VDD.n384 GND 0.005213f
C1973 VDD.n385 GND 0.006477f
C1974 VDD.n386 GND 0.005213f
C1975 VDD.n387 GND 0.006477f
C1976 VDD.n388 GND 0.429674f
C1977 VDD.n389 GND 0.006477f
C1978 VDD.n390 GND 0.005213f
C1979 VDD.n391 GND 0.006477f
C1980 VDD.n392 GND 0.005213f
C1981 VDD.n393 GND 0.006477f
C1982 VDD.n394 GND 0.429674f
C1983 VDD.n395 GND 0.006477f
C1984 VDD.n396 GND 0.005213f
C1985 VDD.n397 GND 0.006477f
C1986 VDD.n398 GND 0.005213f
C1987 VDD.n399 GND 0.006477f
C1988 VDD.n400 GND 0.429674f
C1989 VDD.n401 GND 0.006477f
C1990 VDD.n402 GND 0.005213f
C1991 VDD.n403 GND 0.006477f
C1992 VDD.n404 GND 0.005213f
C1993 VDD.n405 GND 0.006477f
C1994 VDD.n406 GND 0.36952f
C1995 VDD.n407 GND 0.006477f
C1996 VDD.n408 GND 0.005213f
C1997 VDD.n409 GND 0.006477f
C1998 VDD.n410 GND 0.005213f
C1999 VDD.n411 GND 0.006477f
C2000 VDD.n412 GND 0.429674f
C2001 VDD.t37 GND 0.214837f
C2002 VDD.n413 GND 0.006477f
C2003 VDD.n414 GND 0.005213f
C2004 VDD.n415 GND 0.006477f
C2005 VDD.n416 GND 0.005213f
C2006 VDD.n417 GND 0.006477f
C2007 VDD.n418 GND 0.429674f
C2008 VDD.n419 GND 0.006477f
C2009 VDD.n420 GND 0.005213f
C2010 VDD.n421 GND 0.006477f
C2011 VDD.n422 GND 0.005213f
C2012 VDD.n423 GND 0.006477f
C2013 VDD.n424 GND 0.429674f
C2014 VDD.n425 GND 0.006477f
C2015 VDD.n426 GND 0.005213f
C2016 VDD.n427 GND 0.006477f
C2017 VDD.n428 GND 0.005213f
C2018 VDD.n429 GND 0.006477f
C2019 VDD.n430 GND 0.429674f
C2020 VDD.n431 GND 0.006477f
C2021 VDD.n432 GND 0.005213f
C2022 VDD.n433 GND 0.006477f
C2023 VDD.n434 GND 0.005213f
C2024 VDD.n435 GND 0.006477f
C2025 VDD.n436 GND 0.429674f
C2026 VDD.n437 GND 0.006477f
C2027 VDD.n438 GND 0.005213f
C2028 VDD.n439 GND 0.006477f
C2029 VDD.n440 GND 0.005213f
C2030 VDD.n441 GND 0.006477f
C2031 VDD.n442 GND 0.429674f
C2032 VDD.n443 GND 0.006477f
C2033 VDD.n444 GND 0.005213f
C2034 VDD.n445 GND 0.006477f
C2035 VDD.n446 GND 0.005213f
C2036 VDD.n447 GND 0.006477f
C2037 VDD.n448 GND 0.244914f
C2038 VDD.n449 GND 0.006477f
C2039 VDD.n450 GND 0.005213f
C2040 VDD.n451 GND 0.006477f
C2041 VDD.n452 GND 0.005213f
C2042 VDD.n453 GND 0.006477f
C2043 VDD.n454 GND 0.429674f
C2044 VDD.n455 GND 0.006477f
C2045 VDD.n456 GND 0.005213f
C2046 VDD.n457 GND 0.006477f
C2047 VDD.n458 GND 0.005213f
C2048 VDD.n459 GND 0.006477f
C2049 VDD.n460 GND 0.429674f
C2050 VDD.n461 GND 0.006477f
C2051 VDD.n462 GND 0.005213f
C2052 VDD.n463 GND 0.008655f
C2053 VDD.n464 GND 0.004327f
C2054 VDD.n465 GND 0.014826f
C2055 VDD.n466 GND 0.575763f
C2056 VDD.n467 GND 0.014826f
C2057 VDD.n468 GND 0.004327f
C2058 VDD.n469 GND 0.008031f
C2059 VDD.n470 GND 0.003303f
C2060 VDD.n471 GND 0.004404f
C2061 VDD.n472 GND 0.004404f
C2062 VDD.n473 GND 0.552131f
C2063 VDD.n474 GND 0.004404f
C2064 VDD.n475 GND 0.004404f
C2065 VDD.n476 GND 0.003854f
C2066 VDD.n478 GND 0.004404f
C2067 VDD.t115 GND 0.068381f
C2068 VDD.t114 GND 0.084764f
C2069 VDD.t113 GND 0.489916f
C2070 VDD.n479 GND 0.064611f
C2071 VDD.n480 GND 0.042608f
C2072 VDD.n481 GND 0.006294f
C2073 VDD.n482 GND 0.010674f
C2074 VDD.n484 GND 0.004404f
C2075 VDD.n485 GND 0.292178f
C2076 VDD.n486 GND 0.010151f
C2077 VDD.n487 GND 0.010151f
C2078 VDD.n488 GND 0.004404f
C2079 VDD.n489 GND 0.01038f
C2080 VDD.n490 GND 0.004404f
C2081 VDD.n491 GND 0.004404f
C2082 VDD.n493 GND 0.004404f
C2083 VDD.n494 GND 0.004404f
C2084 VDD.n496 GND 0.004404f
C2085 VDD.n497 GND 0.006477f
C2086 VDD.n498 GND 0.005213f
C2087 VDD.n499 GND 0.006477f
C2088 VDD.t9 GND 2.59523f
C2089 VDD.t140 GND 5.0057f
C2090 VDD.n513 GND 0.014967f
C2091 VDD.n514 GND 0.006477f
C2092 VDD.n515 GND 0.006477f
C2093 VDD.n516 GND 0.006477f
C2094 VDD.n517 GND 0.006477f
C2095 VDD.n518 GND 0.006477f
C2096 VDD.n519 GND 0.006477f
C2097 VDD.n520 GND 0.006477f
C2098 VDD.n521 GND 0.006477f
C2099 VDD.n522 GND 0.006477f
C2100 VDD.n523 GND 0.006477f
C2101 VDD.n524 GND 0.006477f
C2102 VDD.n525 GND 0.006477f
C2103 VDD.n526 GND 0.006477f
C2104 VDD.t95 GND 0.086094f
C2105 VDD.t96 GND 0.107631f
C2106 VDD.t93 GND 0.799934f
C2107 VDD.n527 GND 0.078348f
C2108 VDD.n528 GND 0.048083f
C2109 VDD.n529 GND 0.006477f
C2110 VDD.n530 GND 0.006477f
C2111 VDD.n531 GND 0.006477f
C2112 VDD.n532 GND 0.006477f
C2113 VDD.n533 GND 0.006477f
C2114 VDD.n534 GND 0.006477f
C2115 VDD.n535 GND 0.006477f
C2116 VDD.n536 GND 0.006477f
C2117 VDD.n537 GND 0.006477f
C2118 VDD.n538 GND 0.006477f
C2119 VDD.n539 GND 0.006477f
C2120 VDD.n540 GND 0.006477f
C2121 VDD.n541 GND 0.006477f
C2122 VDD.n542 GND 0.006477f
C2123 VDD.n543 GND 0.006477f
C2124 VDD.n544 GND 0.002502f
C2125 VDD.t108 GND 0.086094f
C2126 VDD.t109 GND 0.107631f
C2127 VDD.t107 GND 0.799934f
C2128 VDD.n545 GND 0.078348f
C2129 VDD.n546 GND 0.048083f
C2130 VDD.n547 GND 0.008028f
C2131 VDD.n548 GND 0.006477f
C2132 VDD.n549 GND 0.002711f
C2133 VDD.n550 GND 0.005213f
C2134 VDD.n551 GND 0.006477f
C2135 VDD.n552 GND 0.006477f
C2136 VDD.n553 GND 0.005213f
C2137 VDD.n554 GND 0.005213f
C2138 VDD.n555 GND 0.006477f
C2139 VDD.n556 GND 0.006477f
C2140 VDD.n557 GND 0.005213f
C2141 VDD.n558 GND 0.005213f
C2142 VDD.n559 GND 0.006477f
C2143 VDD.n560 GND 0.006477f
C2144 VDD.n561 GND 0.005213f
C2145 VDD.n562 GND 0.005213f
C2146 VDD.n563 GND 0.006477f
C2147 VDD.n564 GND 0.006477f
C2148 VDD.n565 GND 0.005213f
C2149 VDD.n566 GND 0.005213f
C2150 VDD.n567 GND 0.006477f
C2151 VDD.n568 GND 0.006477f
C2152 VDD.n569 GND 0.005213f
C2153 VDD.n570 GND 0.005213f
C2154 VDD.n571 GND 0.006477f
C2155 VDD.n572 GND 0.006477f
C2156 VDD.n573 GND 0.005213f
C2157 VDD.n574 GND 0.005213f
C2158 VDD.n575 GND 0.006477f
C2159 VDD.n576 GND 0.006477f
C2160 VDD.n577 GND 0.004744f
C2161 VDD.n578 GND 0.010634f
C2162 VDD.n579 GND 0.006477f
C2163 VDD.n580 GND 0.006477f
C2164 VDD.n581 GND 0.003962f
C2165 VDD.n582 GND 0.005213f
C2166 VDD.n583 GND 0.006477f
C2167 VDD.n584 GND 0.006477f
C2168 VDD.n585 GND 0.005213f
C2169 VDD.n586 GND 0.005213f
C2170 VDD.n587 GND 0.006477f
C2171 VDD.n588 GND 0.006477f
C2172 VDD.n589 GND 0.005213f
C2173 VDD.n590 GND 0.005213f
C2174 VDD.n591 GND 0.006477f
C2175 VDD.n592 GND 0.006477f
C2176 VDD.n593 GND 0.005213f
C2177 VDD.n594 GND 0.005213f
C2178 VDD.n595 GND 0.006477f
C2179 VDD.n596 GND 0.006477f
C2180 VDD.n597 GND 0.005213f
C2181 VDD.n598 GND 0.005213f
C2182 VDD.n599 GND 0.005213f
C2183 VDD.n600 GND 0.006477f
C2184 VDD.n601 GND 3.08076f
C2185 VDD.n603 GND 0.014967f
C2186 VDD.n604 GND 0.004327f
C2187 VDD.n605 GND 0.008031f
C2188 VDD.n606 GND 0.661292f
C2189 VDD.n607 GND 0.119937f
C2190 VDD.n609 GND 0.003303f
C2191 VDD.n610 GND 0.004404f
C2192 VDD.n611 GND 0.004404f
C2193 VDD.n613 GND 0.004404f
C2194 VDD.t80 GND 0.068381f
C2195 VDD.t79 GND 0.084764f
C2196 VDD.t77 GND 0.489916f
C2197 VDD.n614 GND 0.064611f
C2198 VDD.n615 GND 0.042608f
C2199 VDD.n616 GND 0.004404f
C2200 VDD.n618 GND 0.004404f
C2201 VDD.n619 GND 0.004404f
C2202 VDD.n620 GND 0.292178f
C2203 VDD.n621 GND 0.004404f
C2204 VDD.n622 GND 0.004404f
C2205 VDD.n623 GND 0.004404f
C2206 VDD.n624 GND 0.004404f
C2207 VDD.n625 GND 0.004404f
C2208 VDD.n626 GND 0.292178f
C2209 VDD.n627 GND 0.004404f
C2210 VDD.n628 GND 0.004404f
C2211 VDD.n629 GND 0.004404f
C2212 VDD.n630 GND 0.004404f
C2213 VDD.n631 GND 0.004404f
C2214 VDD.n632 GND 0.004404f
C2215 VDD.n633 GND 0.214837f
C2216 VDD.n634 GND 0.004404f
C2217 VDD.n635 GND 0.004404f
C2218 VDD.n636 GND 0.004404f
C2219 VDD.n637 GND 0.004404f
C2220 VDD.n638 GND 0.004404f
C2221 VDD.t12 GND 0.146089f
C2222 VDD.n639 GND 0.004404f
C2223 VDD.n640 GND 0.004404f
C2224 VDD.t78 GND 0.146089f
C2225 VDD.n641 GND 0.004404f
C2226 VDD.n642 GND 0.004404f
C2227 VDD.n643 GND 0.004404f
C2228 VDD.n644 GND 0.292178f
C2229 VDD.n645 GND 0.004404f
C2230 VDD.n646 GND 0.004404f
C2231 VDD.n647 GND 0.195502f
C2232 VDD.n648 GND 0.004404f
C2233 VDD.n649 GND 0.004404f
C2234 VDD.n650 GND 0.004404f
C2235 VDD.n651 GND 0.292178f
C2236 VDD.n652 GND 0.004404f
C2237 VDD.n653 GND 0.004404f
C2238 VDD.n654 GND 0.004404f
C2239 VDD.n655 GND 0.004404f
C2240 VDD.n656 GND 0.004404f
C2241 VDD.n657 GND 0.292178f
C2242 VDD.n658 GND 0.004404f
C2243 VDD.n659 GND 0.004404f
C2244 VDD.n660 GND 0.004404f
C2245 VDD.n661 GND 0.004404f
C2246 VDD.n662 GND 0.004404f
C2247 VDD.n663 GND 0.292178f
C2248 VDD.n664 GND 0.004404f
C2249 VDD.n665 GND 0.004404f
C2250 VDD.n666 GND 0.004404f
C2251 VDD.n667 GND 0.004404f
C2252 VDD.n668 GND 0.004404f
C2253 VDD.n669 GND 0.292178f
C2254 VDD.n670 GND 0.004404f
C2255 VDD.n671 GND 0.004404f
C2256 VDD.n672 GND 0.004404f
C2257 VDD.n673 GND 0.004404f
C2258 VDD.n674 GND 0.004404f
C2259 VDD.n675 GND 0.161128f
C2260 VDD.n676 GND 0.004404f
C2261 VDD.n677 GND 0.004404f
C2262 VDD.n678 GND 0.004404f
C2263 VDD.n679 GND 0.004404f
C2264 VDD.n680 GND 0.004404f
C2265 VDD.n681 GND 0.163276f
C2266 VDD.n682 GND 0.004404f
C2267 VDD.n683 GND 0.004404f
C2268 VDD.t59 GND 0.146089f
C2269 VDD.n684 GND 0.004404f
C2270 VDD.n685 GND 0.004404f
C2271 VDD.n686 GND 0.004404f
C2272 VDD.n687 GND 0.292178f
C2273 VDD.n688 GND 0.004404f
C2274 VDD.n689 GND 0.004404f
C2275 VDD.t45 GND 0.146089f
C2276 VDD.n690 GND 0.004404f
C2277 VDD.n691 GND 0.004404f
C2278 VDD.n692 GND 0.004404f
C2279 VDD.n693 GND 0.292178f
C2280 VDD.n694 GND 0.004404f
C2281 VDD.n695 GND 0.004404f
C2282 VDD.n696 GND 0.004404f
C2283 VDD.n697 GND 0.004404f
C2284 VDD.n698 GND 0.004404f
C2285 VDD.n699 GND 0.292178f
C2286 VDD.n700 GND 0.004404f
C2287 VDD.n701 GND 0.004404f
C2288 VDD.n702 GND 0.004404f
C2289 VDD.n703 GND 0.004404f
C2290 VDD.n704 GND 0.004404f
C2291 VDD.n705 GND 0.292178f
C2292 VDD.n706 GND 0.004404f
C2293 VDD.n707 GND 0.004404f
C2294 VDD.n708 GND 0.004404f
C2295 VDD.n709 GND 0.004404f
C2296 VDD.n710 GND 0.004404f
C2297 VDD.n711 GND 0.225579f
C2298 VDD.n712 GND 0.004404f
C2299 VDD.n713 GND 0.004404f
C2300 VDD.n714 GND 0.004404f
C2301 VDD.n715 GND 0.004404f
C2302 VDD.n716 GND 0.004404f
C2303 VDD.n717 GND 0.227727f
C2304 VDD.n718 GND 0.004404f
C2305 VDD.n719 GND 0.004404f
C2306 VDD.t19 GND 0.146089f
C2307 VDD.n720 GND 0.004404f
C2308 VDD.n721 GND 0.004404f
C2309 VDD.n722 GND 0.004404f
C2310 VDD.n723 GND 0.292178f
C2311 VDD.n724 GND 0.004404f
C2312 VDD.n725 GND 0.004404f
C2313 VDD.t4 GND 0.146089f
C2314 VDD.n726 GND 0.004404f
C2315 VDD.n727 GND 0.004404f
C2316 VDD.n728 GND 0.004404f
C2317 VDD.n729 GND 0.292178f
C2318 VDD.n730 GND 0.004404f
C2319 VDD.n731 GND 0.004404f
C2320 VDD.n732 GND 0.004404f
C2321 VDD.n733 GND 0.004404f
C2322 VDD.n734 GND 0.004404f
C2323 VDD.n735 GND 0.292178f
C2324 VDD.n736 GND 0.004404f
C2325 VDD.n737 GND 0.004404f
C2326 VDD.n738 GND 0.004404f
C2327 VDD.n739 GND 0.004404f
C2328 VDD.n740 GND 0.004404f
C2329 VDD.n741 GND 0.292178f
C2330 VDD.n742 GND 0.004404f
C2331 VDD.n743 GND 0.004404f
C2332 VDD.n744 GND 0.004404f
C2333 VDD.n745 GND 0.004404f
C2334 VDD.n746 GND 0.004404f
C2335 VDD.n747 GND 0.292178f
C2336 VDD.n748 GND 0.004404f
C2337 VDD.n749 GND 0.004404f
C2338 VDD.n750 GND 0.004404f
C2339 VDD.n751 GND 0.004404f
C2340 VDD.n752 GND 0.004404f
C2341 VDD.n753 GND 0.292178f
C2342 VDD.n754 GND 0.004404f
C2343 VDD.n755 GND 0.004404f
C2344 VDD.n756 GND 0.004404f
C2345 VDD.n757 GND 0.004404f
C2346 VDD.n758 GND 0.004404f
C2347 VDD.n759 GND 0.292178f
C2348 VDD.n760 GND 0.004404f
C2349 VDD.n761 GND 0.004404f
C2350 VDD.n762 GND 0.004404f
C2351 VDD.n763 GND 0.004404f
C2352 VDD.n764 GND 0.004404f
C2353 VDD.n765 GND 0.004404f
C2354 VDD.n766 GND 0.292178f
C2355 VDD.n767 GND 0.004404f
C2356 VDD.n768 GND 0.004404f
C2357 VDD.n769 GND 0.004404f
C2358 VDD.n770 GND 0.004404f
C2359 VDD.n771 GND 0.004404f
C2360 VDD.t30 GND 0.146089f
C2361 VDD.n772 GND 0.004404f
C2362 VDD.n773 GND 0.004404f
C2363 VDD.n774 GND 0.004404f
C2364 VDD.n775 GND 0.004404f
C2365 VDD.n776 GND 0.004404f
C2366 VDD.n777 GND 0.004404f
C2367 VDD.n778 GND 0.292178f
C2368 VDD.n779 GND 0.004404f
C2369 VDD.n780 GND 0.004404f
C2370 VDD.n781 GND 0.242766f
C2371 VDD.n782 GND 0.004404f
C2372 VDD.n783 GND 0.004404f
C2373 VDD.n784 GND 0.004404f
C2374 VDD.n785 GND 0.292178f
C2375 VDD.n786 GND 0.004404f
C2376 VDD.n787 GND 0.004404f
C2377 VDD.n788 GND 0.004404f
C2378 VDD.n789 GND 0.004404f
C2379 VDD.n790 GND 0.004404f
C2380 VDD.n791 GND 0.292178f
C2381 VDD.n792 GND 0.004404f
C2382 VDD.n793 GND 0.004404f
C2383 VDD.n794 GND 0.004404f
C2384 VDD.n795 GND 0.004404f
C2385 VDD.n796 GND 0.004404f
C2386 VDD.t15 GND 0.146089f
C2387 VDD.n797 GND 0.004404f
C2388 VDD.n798 GND 0.004404f
C2389 VDD.n799 GND 0.004404f
C2390 VDD.n800 GND 0.004404f
C2391 VDD.n801 GND 0.004404f
C2392 VDD.n802 GND 0.292178f
C2393 VDD.n803 GND 0.004404f
C2394 VDD.n804 GND 0.004404f
C2395 VDD.n805 GND 0.227727f
C2396 VDD.n806 GND 0.004404f
C2397 VDD.n807 GND 0.004404f
C2398 VDD.n808 GND 0.004404f
C2399 VDD.t136 GND 0.146089f
C2400 VDD.n809 GND 0.004404f
C2401 VDD.n810 GND 0.004404f
C2402 VDD.n811 GND 0.004404f
C2403 VDD.n812 GND 0.004404f
C2404 VDD.n813 GND 0.004404f
C2405 VDD.n814 GND 0.292178f
C2406 VDD.n815 GND 0.004404f
C2407 VDD.n816 GND 0.004404f
C2408 VDD.n817 GND 0.178315f
C2409 VDD.n818 GND 0.004404f
C2410 VDD.n819 GND 0.004404f
C2411 VDD.n820 GND 0.004404f
C2412 VDD.n821 GND 0.292178f
C2413 VDD.n822 GND 0.004404f
C2414 VDD.n823 GND 0.004404f
C2415 VDD.n824 GND 0.004404f
C2416 VDD.n825 GND 0.004404f
C2417 VDD.n826 GND 0.004404f
C2418 VDD.n827 GND 0.292178f
C2419 VDD.n828 GND 0.004404f
C2420 VDD.n829 GND 0.004404f
C2421 VDD.n830 GND 0.004404f
C2422 VDD.n831 GND 0.004404f
C2423 VDD.n832 GND 0.004404f
C2424 VDD.t11 GND 0.146089f
C2425 VDD.n833 GND 0.004404f
C2426 VDD.n834 GND 0.004404f
C2427 VDD.n835 GND 0.004404f
C2428 VDD.n836 GND 0.004404f
C2429 VDD.n837 GND 0.004404f
C2430 VDD.n838 GND 0.292178f
C2431 VDD.n839 GND 0.004404f
C2432 VDD.n840 GND 0.004404f
C2433 VDD.n841 GND 0.163276f
C2434 VDD.n842 GND 0.004404f
C2435 VDD.n843 GND 0.004404f
C2436 VDD.n844 GND 0.004404f
C2437 VDD.n845 GND 0.178315f
C2438 VDD.n846 GND 0.004404f
C2439 VDD.n847 GND 0.004404f
C2440 VDD.n848 GND 0.004404f
C2441 VDD.n849 GND 0.004404f
C2442 VDD.n850 GND 0.004404f
C2443 VDD.n851 GND 0.292178f
C2444 VDD.n852 GND 0.004404f
C2445 VDD.n853 GND 0.004404f
C2446 VDD.t33 GND 0.146089f
C2447 VDD.n854 GND 0.004404f
C2448 VDD.n855 GND 0.004404f
C2449 VDD.n856 GND 0.004404f
C2450 VDD.n857 GND 0.292178f
C2451 VDD.n858 GND 0.004404f
C2452 VDD.n859 GND 0.004404f
C2453 VDD.n860 GND 0.004404f
C2454 VDD.n861 GND 0.004404f
C2455 VDD.n862 GND 0.004404f
C2456 VDD.n863 GND 0.292178f
C2457 VDD.n864 GND 0.004404f
C2458 VDD.n865 GND 0.004404f
C2459 VDD.n866 GND 0.004404f
C2460 VDD.n867 GND 0.004404f
C2461 VDD.n868 GND 0.004404f
C2462 VDD.n869 GND 0.292178f
C2463 VDD.n870 GND 0.004404f
C2464 VDD.n871 GND 0.004404f
C2465 VDD.n872 GND 0.004404f
C2466 VDD.n873 GND 0.004404f
C2467 VDD.n874 GND 0.004404f
C2468 VDD.n875 GND 0.292178f
C2469 VDD.n876 GND 0.004404f
C2470 VDD.n877 GND 0.004404f
C2471 VDD.n878 GND 0.004404f
C2472 VDD.n879 GND 0.004404f
C2473 VDD.n880 GND 0.004404f
C2474 VDD.t90 GND 0.146089f
C2475 VDD.n881 GND 0.004404f
C2476 VDD.n882 GND 0.004404f
C2477 VDD.n883 GND 0.004404f
C2478 VDD.n884 GND 0.004404f
C2479 VDD.n885 GND 0.004404f
C2480 VDD.n886 GND 0.292178f
C2481 VDD.n887 GND 0.004404f
C2482 VDD.n888 GND 0.004404f
C2483 VDD.t40 GND 0.146089f
C2484 VDD.n889 GND 0.004404f
C2485 VDD.n890 GND 0.004404f
C2486 VDD.n891 GND 0.004404f
C2487 VDD.n892 GND 0.292178f
C2488 VDD.n893 GND 0.004404f
C2489 VDD.n894 GND 0.004404f
C2490 VDD.n895 GND 0.004404f
C2491 VDD.n896 GND 0.004404f
C2492 VDD.n897 GND 0.004404f
C2493 VDD.n898 GND 0.292178f
C2494 VDD.n899 GND 0.004404f
C2495 VDD.n900 GND 0.004404f
C2496 VDD.n901 GND 0.004404f
C2497 VDD.n902 GND 0.01038f
C2498 VDD.n903 GND 0.01038f
C2499 VDD.n904 GND 0.388855f
C2500 VDD.n924 GND 0.004404f
C2501 VDD.n925 GND 0.010151f
C2502 VDD.n926 GND 0.004404f
C2503 VDD.n927 GND 0.004404f
C2504 VDD.n928 GND 0.004404f
C2505 VDD.n929 GND 0.292178f
C2506 VDD.n930 GND 0.004404f
C2507 VDD.n931 GND 0.004404f
C2508 VDD.n932 GND 0.004404f
C2509 VDD.n933 GND 0.010151f
C2510 VDD.n934 GND 0.004404f
C2511 VDD.t118 GND 0.068381f
C2512 VDD.t117 GND 0.084764f
C2513 VDD.t116 GND 0.489916f
C2514 VDD.n935 GND 0.064611f
C2515 VDD.n936 GND 0.042608f
C2516 VDD.n937 GND 0.004404f
C2517 VDD.n938 GND 0.004404f
C2518 VDD.n939 GND 0.292178f
C2519 VDD.n940 GND 0.004404f
C2520 VDD.n941 GND 0.004404f
C2521 VDD.n942 GND 0.004404f
C2522 VDD.n943 GND 0.004404f
C2523 VDD.n944 GND 0.004404f
C2524 VDD.n945 GND 0.195502f
C2525 VDD.n946 GND 0.004404f
C2526 VDD.n947 GND 0.004404f
C2527 VDD.n948 GND 0.004404f
C2528 VDD.n949 GND 0.004404f
C2529 VDD.n950 GND 0.004404f
C2530 VDD.n951 GND 0.004404f
C2531 VDD.t74 GND 0.146089f
C2532 VDD.n952 GND 0.004404f
C2533 VDD.n953 GND 0.004404f
C2534 VDD.t57 GND 0.146089f
C2535 VDD.n954 GND 0.004404f
C2536 VDD.n955 GND 0.004404f
C2537 VDD.n956 GND 0.004404f
C2538 VDD.n957 GND 0.292178f
C2539 VDD.n958 GND 0.004404f
C2540 VDD.n959 GND 0.004404f
C2541 VDD.n960 GND 0.223431f
C2542 VDD.n961 GND 0.004404f
C2543 VDD.n962 GND 0.004404f
C2544 VDD.n963 GND 0.004404f
C2545 VDD.n964 GND 0.292178f
C2546 VDD.n965 GND 0.004404f
C2547 VDD.n966 GND 0.004404f
C2548 VDD.n967 GND 0.004404f
C2549 VDD.n968 GND 0.004404f
C2550 VDD.n969 GND 0.004404f
C2551 VDD.n970 GND 0.292178f
C2552 VDD.n971 GND 0.004404f
C2553 VDD.n972 GND 0.004404f
C2554 VDD.n973 GND 0.004404f
C2555 VDD.n974 GND 0.004404f
C2556 VDD.n975 GND 0.004404f
C2557 VDD.n976 GND 0.292178f
C2558 VDD.n977 GND 0.004404f
C2559 VDD.n978 GND 0.004404f
C2560 VDD.n979 GND 0.004404f
C2561 VDD.n980 GND 0.004404f
C2562 VDD.n981 GND 0.004404f
C2563 VDD.n982 GND 0.259953f
C2564 VDD.n983 GND 0.004404f
C2565 VDD.n984 GND 0.004404f
C2566 VDD.n985 GND 0.004404f
C2567 VDD.n986 GND 0.004404f
C2568 VDD.n987 GND 0.004404f
C2569 VDD.n988 GND 0.292178f
C2570 VDD.n989 GND 0.004404f
C2571 VDD.n990 GND 0.004404f
C2572 VDD.t61 GND 0.146089f
C2573 VDD.n991 GND 0.004404f
C2574 VDD.n992 GND 0.004404f
C2575 VDD.n993 GND 0.004404f
C2576 VDD.n994 GND 0.292178f
C2577 VDD.n995 GND 0.004404f
C2578 VDD.n996 GND 0.004404f
C2579 VDD.n997 GND 0.004404f
C2580 VDD.n998 GND 0.004404f
C2581 VDD.n999 GND 0.004404f
C2582 VDD.t14 GND 0.146089f
C2583 VDD.n1000 GND 0.004404f
C2584 VDD.n1001 GND 0.004404f
C2585 VDD.n1002 GND 0.004404f
C2586 VDD.n1003 GND 0.004404f
C2587 VDD.n1004 GND 0.004404f
C2588 VDD.n1005 GND 0.292178f
C2589 VDD.n1006 GND 0.004404f
C2590 VDD.n1007 GND 0.004404f
C2591 VDD.n1008 GND 0.274991f
C2592 VDD.n1009 GND 0.004404f
C2593 VDD.n1010 GND 0.004404f
C2594 VDD.n1011 GND 0.004404f
C2595 VDD.n1012 GND 0.292178f
C2596 VDD.n1013 GND 0.004404f
C2597 VDD.n1014 GND 0.004404f
C2598 VDD.n1015 GND 0.004404f
C2599 VDD.n1016 GND 0.004404f
C2600 VDD.n1017 GND 0.004404f
C2601 VDD.n1018 GND 0.292178f
C2602 VDD.n1019 GND 0.004404f
C2603 VDD.n1020 GND 0.004404f
C2604 VDD.n1021 GND 0.004404f
C2605 VDD.n1022 GND 0.004404f
C2606 VDD.n1023 GND 0.004404f
C2607 VDD.t0 GND 0.146089f
C2608 VDD.n1024 GND 0.004404f
C2609 VDD.n1025 GND 0.004404f
C2610 VDD.n1026 GND 0.004404f
C2611 VDD.n1027 GND 0.004404f
C2612 VDD.n1028 GND 0.004404f
C2613 VDD.n1029 GND 0.292178f
C2614 VDD.n1030 GND 0.004404f
C2615 VDD.n1031 GND 0.004404f
C2616 VDD.n1032 GND 0.259953f
C2617 VDD.n1033 GND 0.004404f
C2618 VDD.n1034 GND 0.004404f
C2619 VDD.n1035 GND 0.004404f
C2620 VDD.t32 GND 0.146089f
C2621 VDD.n1036 GND 0.004404f
C2622 VDD.n1037 GND 0.004404f
C2623 VDD.n1038 GND 0.004404f
C2624 VDD.n1039 GND 0.004404f
C2625 VDD.n1040 GND 0.004404f
C2626 VDD.n1041 GND 0.292178f
C2627 VDD.n1042 GND 0.004404f
C2628 VDD.n1043 GND 0.004404f
C2629 VDD.n1044 GND 0.21054f
C2630 VDD.n1045 GND 0.004404f
C2631 VDD.n1046 GND 0.004404f
C2632 VDD.n1047 GND 0.004404f
C2633 VDD.n1048 GND 0.292178f
C2634 VDD.n1049 GND 0.004404f
C2635 VDD.n1050 GND 0.004404f
C2636 VDD.n1051 GND 0.004404f
C2637 VDD.n1052 GND 0.004404f
C2638 VDD.n1053 GND 0.004404f
C2639 VDD.n1054 GND 0.292178f
C2640 VDD.n1055 GND 0.004404f
C2641 VDD.n1056 GND 0.004404f
C2642 VDD.n1057 GND 0.004404f
C2643 VDD.n1058 GND 0.004404f
C2644 VDD.n1059 GND 0.004404f
C2645 VDD.t134 GND 0.146089f
C2646 VDD.n1060 GND 0.004404f
C2647 VDD.n1061 GND 0.004404f
C2648 VDD.n1062 GND 0.004404f
C2649 VDD.n1063 GND 0.004404f
C2650 VDD.n1064 GND 0.004404f
C2651 VDD.n1065 GND 0.292178f
C2652 VDD.n1066 GND 0.004404f
C2653 VDD.n1067 GND 0.004404f
C2654 VDD.n1068 GND 0.195502f
C2655 VDD.n1069 GND 0.004404f
C2656 VDD.n1070 GND 0.004404f
C2657 VDD.n1071 GND 0.004404f
C2658 VDD.t25 GND 0.292178f
C2659 VDD.n1072 GND 0.004404f
C2660 VDD.n1073 GND 0.004404f
C2661 VDD.n1074 GND 0.004404f
C2662 VDD.n1075 GND 0.004404f
C2663 VDD.n1076 GND 0.004404f
C2664 VDD.n1077 GND 0.292178f
C2665 VDD.n1078 GND 0.004404f
C2666 VDD.n1079 GND 0.004404f
C2667 VDD.n1080 GND 0.004404f
C2668 VDD.n1081 GND 0.004404f
C2669 VDD.n1082 GND 0.004404f
C2670 VDD.n1083 GND 0.292178f
C2671 VDD.n1084 GND 0.004404f
C2672 VDD.n1085 GND 0.004404f
C2673 VDD.n1086 GND 0.004404f
C2674 VDD.n1087 GND 0.004404f
C2675 VDD.n1088 GND 0.004404f
C2676 VDD.n1089 GND 0.292178f
C2677 VDD.n1090 GND 0.004404f
C2678 VDD.n1091 GND 0.004404f
C2679 VDD.n1092 GND 0.004404f
C2680 VDD.n1093 GND 0.004404f
C2681 VDD.n1094 GND 0.004404f
C2682 VDD.n1095 GND 0.292178f
C2683 VDD.n1096 GND 0.004404f
C2684 VDD.n1097 GND 0.004404f
C2685 VDD.n1098 GND 0.004404f
C2686 VDD.n1099 GND 0.004404f
C2687 VDD.n1100 GND 0.004404f
C2688 VDD.n1101 GND 0.292178f
C2689 VDD.n1102 GND 0.004404f
C2690 VDD.n1103 GND 0.004404f
C2691 VDD.n1104 GND 0.004404f
C2692 VDD.n1105 GND 0.004404f
C2693 VDD.n1106 GND 0.004404f
C2694 VDD.n1107 GND 0.21054f
C2695 VDD.n1108 GND 0.004404f
C2696 VDD.n1109 GND 0.004404f
C2697 VDD.n1110 GND 0.004404f
C2698 VDD.n1111 GND 0.004404f
C2699 VDD.n1112 GND 0.004404f
C2700 VDD.n1113 GND 0.212689f
C2701 VDD.n1114 GND 0.004404f
C2702 VDD.n1115 GND 0.004404f
C2703 VDD.t132 GND 0.146089f
C2704 VDD.n1116 GND 0.004404f
C2705 VDD.n1117 GND 0.004404f
C2706 VDD.n1118 GND 0.004404f
C2707 VDD.n1119 GND 0.292178f
C2708 VDD.n1120 GND 0.004404f
C2709 VDD.n1121 GND 0.004404f
C2710 VDD.t43 GND 0.146089f
C2711 VDD.n1122 GND 0.004404f
C2712 VDD.n1123 GND 0.004404f
C2713 VDD.n1124 GND 0.004404f
C2714 VDD.n1125 GND 0.292178f
C2715 VDD.n1126 GND 0.004404f
C2716 VDD.n1127 GND 0.004404f
C2717 VDD.n1128 GND 0.004404f
C2718 VDD.n1129 GND 0.004404f
C2719 VDD.n1130 GND 0.004404f
C2720 VDD.n1131 GND 0.292178f
C2721 VDD.n1132 GND 0.004404f
C2722 VDD.n1133 GND 0.004404f
C2723 VDD.n1134 GND 0.004404f
C2724 VDD.n1135 GND 0.004404f
C2725 VDD.n1136 GND 0.004404f
C2726 VDD.n1137 GND 0.292178f
C2727 VDD.n1138 GND 0.004404f
C2728 VDD.n1139 GND 0.004404f
C2729 VDD.n1140 GND 0.004404f
C2730 VDD.n1141 GND 0.004404f
C2731 VDD.n1142 GND 0.004404f
C2732 VDD.n1143 GND 0.274991f
C2733 VDD.n1144 GND 0.004404f
C2734 VDD.n1145 GND 0.004404f
C2735 VDD.n1146 GND 0.004404f
C2736 VDD.n1147 GND 0.004404f
C2737 VDD.n1148 GND 0.004404f
C2738 VDD.n1149 GND 0.27714f
C2739 VDD.n1150 GND 0.004404f
C2740 VDD.n1151 GND 0.004404f
C2741 VDD.t36 GND 0.146089f
C2742 VDD.n1152 GND 0.004404f
C2743 VDD.n1153 GND 0.004404f
C2744 VDD.n1154 GND 0.004404f
C2745 VDD.n1155 GND 0.292178f
C2746 VDD.n1156 GND 0.004404f
C2747 VDD.n1157 GND 0.004404f
C2748 VDD.t130 GND 0.146089f
C2749 VDD.n1158 GND 0.004404f
C2750 VDD.n1159 GND 0.004404f
C2751 VDD.n1160 GND 0.004404f
C2752 VDD.n1161 GND 0.292178f
C2753 VDD.n1162 GND 0.004404f
C2754 VDD.n1163 GND 0.004404f
C2755 VDD.n1164 GND 0.004404f
C2756 VDD.n1165 GND 0.004404f
C2757 VDD.n1166 GND 0.004404f
C2758 VDD.n1167 GND 0.292178f
C2759 VDD.n1168 GND 0.004404f
C2760 VDD.n1169 GND 0.004404f
C2761 VDD.n1170 GND 0.004404f
C2762 VDD.n1171 GND 0.004404f
C2763 VDD.n1172 GND 0.004404f
C2764 VDD.n1173 GND 0.292178f
C2765 VDD.n1174 GND 0.004404f
C2766 VDD.n1175 GND 0.004404f
C2767 VDD.n1176 GND 0.004404f
C2768 VDD.n1177 GND 0.004404f
C2769 VDD.n1178 GND 0.004404f
C2770 VDD.n1179 GND 0.292178f
C2771 VDD.n1180 GND 0.004404f
C2772 VDD.n1181 GND 0.004404f
C2773 VDD.n1182 GND 0.004404f
C2774 VDD.n1183 GND 0.004404f
C2775 VDD.n1184 GND 0.004404f
C2776 VDD.n1185 GND 0.292178f
C2777 VDD.n1186 GND 0.004404f
C2778 VDD.n1187 GND 0.004404f
C2779 VDD.n1188 GND 0.004404f
C2780 VDD.n1189 GND 0.004404f
C2781 VDD.n1190 GND 0.004404f
C2782 VDD.t2 GND 0.146089f
C2783 VDD.n1191 GND 0.004404f
C2784 VDD.n1192 GND 0.004404f
C2785 VDD.n1193 GND 0.004404f
C2786 VDD.n1194 GND 0.004404f
C2787 VDD.n1195 GND 0.004404f
C2788 VDD.n1196 GND 0.292178f
C2789 VDD.n1197 GND 0.004404f
C2790 VDD.n1198 GND 0.004404f
C2791 VDD.t120 GND 0.146089f
C2792 VDD.n1199 GND 0.004404f
C2793 VDD.n1200 GND 0.004404f
C2794 VDD.n1201 GND 0.004404f
C2795 VDD.n1202 GND 0.292178f
C2796 VDD.n1203 GND 0.004404f
C2797 VDD.n1204 GND 0.004404f
C2798 VDD.n1205 GND 0.004404f
C2799 VDD.n1206 GND 0.004404f
C2800 VDD.n1207 GND 0.004404f
C2801 VDD.n1208 GND 0.292178f
C2802 VDD.n1209 GND 0.004404f
C2803 VDD.n1210 GND 0.004404f
C2804 VDD.n1211 GND 0.004404f
C2805 VDD.n1212 GND 0.010151f
C2806 VDD.n1213 GND 0.010151f
C2807 VDD.n1214 GND 0.388855f
C2808 VDD.n1215 GND 0.004404f
C2809 VDD.n1216 GND 0.004404f
C2810 VDD.n1217 GND 0.010151f
C2811 VDD.n1218 GND 0.004404f
C2812 VDD.n1219 GND 0.004404f
C2813 VDD.t28 GND 2.59523f
C2814 VDD.n1228 GND 0.01038f
C2815 VDD.n1239 GND 0.004404f
C2816 VDD.n1240 GND 0.003303f
C2817 VDD.n1241 GND 0.008655f
C2818 VDD.n1242 GND 0.006477f
C2819 VDD.n1243 GND 0.014967f
C2820 VDD.n1244 GND 0.006477f
C2821 VDD.n1245 GND 0.006477f
C2822 VDD.n1246 GND 0.005213f
C2823 VDD.n1247 GND 0.006477f
C2824 VDD.n1248 GND 0.006477f
C2825 VDD.n1249 GND 0.006477f
C2826 VDD.n1250 GND 0.006477f
C2827 VDD.n1251 GND 0.005213f
C2828 VDD.n1252 GND 0.006477f
C2829 VDD.n1253 GND 0.006477f
C2830 VDD.n1254 GND 0.006477f
C2831 VDD.n1255 GND 0.006477f
C2832 VDD.n1256 GND 0.005213f
C2833 VDD.n1257 GND 0.006477f
C2834 VDD.n1258 GND 0.006477f
C2835 VDD.t84 GND 0.086094f
C2836 VDD.t83 GND 0.107631f
C2837 VDD.t81 GND 0.799934f
C2838 VDD.n1259 GND 0.078348f
C2839 VDD.n1260 GND 0.048083f
C2840 VDD.n1261 GND 0.006477f
C2841 VDD.n1262 GND 0.006477f
C2842 VDD.n1263 GND 0.005213f
C2843 VDD.n1264 GND 0.006477f
C2844 VDD.n1265 GND 0.006477f
C2845 VDD.n1266 GND 0.006477f
C2846 VDD.n1267 GND 0.006477f
C2847 VDD.n1268 GND 0.005213f
C2848 VDD.n1269 GND 0.006477f
C2849 VDD.n1270 GND 0.006477f
C2850 VDD.n1271 GND 0.006477f
C2851 VDD.n1272 GND 0.006477f
C2852 VDD.n1273 GND 0.005213f
C2853 VDD.n1274 GND 0.006477f
C2854 VDD.n1275 GND 0.006477f
C2855 VDD.n1276 GND 0.006477f
C2856 VDD.n1277 GND 0.006477f
C2857 VDD.n1278 GND 0.005213f
C2858 VDD.n1279 GND 0.008031f
C2859 VDD.n1280 GND 0.006477f
C2860 VDD.t99 GND 0.086094f
C2861 VDD.t98 GND 0.107631f
C2862 VDD.t97 GND 0.799934f
C2863 VDD.n1281 GND 0.078348f
C2864 VDD.n1282 GND 0.048083f
C2865 VDD.n1284 GND 0.006477f
C2866 VDD.n1285 GND 0.004327f
C2867 VDD.n1286 GND 0.429674f
C2868 VDD.n1288 GND 0.006477f
C2869 VDD.n1291 GND 0.006477f
C2870 VDD.n1294 GND 0.006477f
C2871 VDD.n1297 GND 0.006477f
C2872 VDD.n1300 GND 0.006477f
C2873 VDD.n1303 GND 0.006477f
C2874 VDD.n1306 GND 0.006477f
C2875 VDD.t42 GND 5.0057f
C2876 VDD.n1308 GND 3.08076f
C2877 VDD.n1309 GND 0.006477f
C2878 VDD.n1310 GND 0.005213f
C2879 VDD.n1311 GND 0.006477f
C2880 VDD.n1312 GND 0.005213f
C2881 VDD.n1313 GND 0.006477f
C2882 VDD.n1314 GND 0.006477f
C2883 VDD.n1315 GND 0.429674f
C2884 VDD.n1316 GND 0.006477f
C2885 VDD.n1317 GND 0.005213f
C2886 VDD.n1318 GND 0.005213f
C2887 VDD.n1319 GND 0.006477f
C2888 VDD.n1320 GND 0.005213f
C2889 VDD.n1321 GND 0.006477f
C2890 VDD.t82 GND 0.214837f
C2891 VDD.n1322 GND 0.006477f
C2892 VDD.n1323 GND 0.005213f
C2893 VDD.n1324 GND 0.006477f
C2894 VDD.n1325 GND 0.005213f
C2895 VDD.n1326 GND 0.006477f
C2896 VDD.n1327 GND 0.429674f
C2897 VDD.n1328 GND 0.006477f
C2898 VDD.n1329 GND 0.005213f
C2899 VDD.n1330 GND 0.005213f
C2900 VDD.n1331 GND 0.006477f
C2901 VDD.n1332 GND 0.005213f
C2902 VDD.n1333 GND 0.006477f
C2903 VDD.n1334 GND 0.429674f
C2904 VDD.n1335 GND 0.006477f
C2905 VDD.n1336 GND 0.005213f
C2906 VDD.n1337 GND 0.006477f
C2907 VDD.n1338 GND 0.005213f
C2908 VDD.n1339 GND 0.006477f
C2909 VDD.n1340 GND 0.429674f
C2910 VDD.n1341 GND 0.006477f
C2911 VDD.n1342 GND 0.005213f
C2912 VDD.n1343 GND 0.006477f
C2913 VDD.n1344 GND 0.005213f
C2914 VDD.n1345 GND 0.006477f
C2915 VDD.n1346 GND 0.429674f
C2916 VDD.n1347 GND 0.006477f
C2917 VDD.n1348 GND 0.005213f
C2918 VDD.n1349 GND 0.006477f
C2919 VDD.n1350 GND 0.005213f
C2920 VDD.n1351 GND 0.006477f
C2921 VDD.n1352 GND 0.429674f
C2922 VDD.n1353 GND 0.006477f
C2923 VDD.n1354 GND 0.005213f
C2924 VDD.n1355 GND 0.006477f
C2925 VDD.n1356 GND 0.005213f
C2926 VDD.n1357 GND 0.006477f
C2927 VDD.n1358 GND 0.429674f
C2928 VDD.n1359 GND 0.006477f
C2929 VDD.n1360 GND 0.005213f
C2930 VDD.n1361 GND 0.006477f
C2931 VDD.n1362 GND 0.005213f
C2932 VDD.n1363 GND 0.006477f
C2933 VDD.t69 GND 0.214837f
C2934 VDD.n1364 GND 0.006477f
C2935 VDD.n1365 GND 0.005213f
C2936 VDD.n1366 GND 0.006477f
C2937 VDD.n1367 GND 0.005213f
C2938 VDD.n1368 GND 0.006477f
C2939 VDD.n1369 GND 0.429674f
C2940 VDD.n1370 GND 0.36952f
C2941 VDD.n1371 GND 0.006477f
C2942 VDD.n1372 GND 0.005213f
C2943 VDD.n1373 GND 0.006477f
C2944 VDD.n1374 GND 0.005213f
C2945 VDD.n1375 GND 0.006477f
C2946 VDD.n1376 GND 0.429674f
C2947 VDD.n1377 GND 0.006477f
C2948 VDD.n1378 GND 0.005213f
C2949 VDD.n1379 GND 0.006477f
C2950 VDD.n1380 GND 0.005213f
C2951 VDD.n1381 GND 0.006477f
C2952 VDD.n1382 GND 0.429674f
C2953 VDD.n1383 GND 0.006477f
C2954 VDD.n1384 GND 0.005213f
C2955 VDD.n1385 GND 0.006477f
C2956 VDD.n1386 GND 0.005213f
C2957 VDD.n1387 GND 0.006477f
C2958 VDD.n1388 GND 0.429674f
C2959 VDD.n1389 GND 0.006477f
C2960 VDD.n1390 GND 0.005213f
C2961 VDD.n1391 GND 0.006477f
C2962 VDD.n1392 GND 0.005213f
C2963 VDD.n1393 GND 0.006477f
C2964 VDD.n1394 GND 0.326552f
C2965 VDD.n1395 GND 0.006477f
C2966 VDD.n1396 GND 0.005213f
C2967 VDD.n1397 GND 0.006477f
C2968 VDD.n1398 GND 0.005213f
C2969 VDD.n1399 GND 0.006477f
C2970 VDD.n1400 GND 0.429674f
C2971 VDD.n1401 GND 0.006477f
C2972 VDD.n1402 GND 0.005213f
C2973 VDD.n1403 GND 0.006477f
C2974 VDD.n1404 GND 0.005213f
C2975 VDD.n1405 GND 0.006477f
C2976 VDD.n1406 GND 0.429674f
C2977 VDD.n1407 GND 0.006477f
C2978 VDD.n1408 GND 0.005213f
C2979 VDD.n1409 GND 0.006477f
C2980 VDD.n1410 GND 0.005213f
C2981 VDD.n1411 GND 0.006477f
C2982 VDD.n1412 GND 0.429674f
C2983 VDD.n1413 GND 0.006477f
C2984 VDD.n1414 GND 0.005213f
C2985 VDD.n1415 GND 0.006477f
C2986 VDD.n1416 GND 0.005213f
C2987 VDD.n1417 GND 0.006477f
C2988 VDD.n1418 GND 0.429674f
C2989 VDD.n1419 GND 0.006477f
C2990 VDD.n1420 GND 0.005213f
C2991 VDD.n1421 GND 0.006477f
C2992 VDD.n1422 GND 0.005213f
C2993 VDD.n1423 GND 0.006477f
C2994 VDD.n1424 GND 0.429674f
C2995 VDD.n1425 GND 0.006477f
C2996 VDD.n1426 GND 0.005213f
C2997 VDD.n1427 GND 0.006477f
C2998 VDD.n1428 GND 0.005213f
C2999 VDD.n1429 GND 0.006477f
C3000 VDD.t52 GND 0.214837f
C3001 VDD.n1430 GND 0.006477f
C3002 VDD.n1431 GND 0.005213f
C3003 VDD.n1432 GND 0.006477f
C3004 VDD.n1433 GND 0.005213f
C3005 VDD.n1434 GND 0.006477f
C3006 VDD.n1435 GND 0.429674f
C3007 VDD.n1436 GND 0.006477f
C3008 VDD.n1437 GND 0.005213f
C3009 VDD.n1438 GND 0.006477f
C3010 VDD.n1439 GND 0.005213f
C3011 VDD.n1440 GND 0.006477f
C3012 VDD.n1441 GND 0.429674f
C3013 VDD.n1442 GND 0.006477f
C3014 VDD.n1443 GND 0.005213f
C3015 VDD.n1444 GND 0.006477f
C3016 VDD.n1445 GND 0.005213f
C3017 VDD.n1446 GND 0.006477f
C3018 VDD.n1447 GND 0.429674f
C3019 VDD.n1448 GND 0.006477f
C3020 VDD.n1449 GND 0.005213f
C3021 VDD.n1450 GND 0.006477f
C3022 VDD.n1451 GND 0.005213f
C3023 VDD.n1452 GND 0.006477f
C3024 VDD.n1453 GND 0.429674f
C3025 VDD.n1454 GND 0.006477f
C3026 VDD.n1455 GND 0.005213f
C3027 VDD.n1456 GND 0.006454f
C3028 VDD.n1457 GND 0.005213f
C3029 VDD.n1458 GND 0.006477f
C3030 VDD.n1459 GND 0.429674f
C3031 VDD.n1460 GND 0.006477f
C3032 VDD.n1461 GND 0.005213f
C3033 VDD.n1462 GND 0.006477f
C3034 VDD.n1463 GND 0.005213f
C3035 VDD.n1464 GND 0.006477f
C3036 VDD.n1465 GND 0.429674f
C3037 VDD.n1466 GND 0.006477f
C3038 VDD.n1467 GND 0.005213f
C3039 VDD.n1468 GND 0.006477f
C3040 VDD.n1469 GND 0.005213f
C3041 VDD.n1470 GND 0.006477f
C3042 VDD.n1471 GND 0.429674f
C3043 VDD.n1472 GND 0.006477f
C3044 VDD.n1473 GND 0.005213f
C3045 VDD.n1474 GND 0.006477f
C3046 VDD.n1475 GND 0.005213f
C3047 VDD.n1476 GND 0.006477f
C3048 VDD.n1477 GND 0.429674f
C3049 VDD.n1478 GND 0.006477f
C3050 VDD.n1479 GND 0.005213f
C3051 VDD.n1480 GND 0.006477f
C3052 VDD.n1481 GND 0.005213f
C3053 VDD.n1482 GND 0.006477f
C3054 VDD.n1483 GND 0.429674f
C3055 VDD.n1484 GND 0.006477f
C3056 VDD.n1485 GND 0.005213f
C3057 VDD.n1486 GND 0.006477f
C3058 VDD.n1487 GND 0.005213f
C3059 VDD.n1488 GND 0.006477f
C3060 VDD.n1489 GND 0.429674f
C3061 VDD.n1490 GND 0.006477f
C3062 VDD.n1491 GND 0.005213f
C3063 VDD.n1492 GND 0.006477f
C3064 VDD.n1493 GND 0.005213f
C3065 VDD.n1494 GND 0.006477f
C3066 VDD.n1495 GND 0.266398f
C3067 VDD.n1496 GND 0.006477f
C3068 VDD.n1497 GND 0.005213f
C3069 VDD.n1498 GND 0.006477f
C3070 VDD.n1499 GND 0.005213f
C3071 VDD.n1500 GND 0.006477f
C3072 VDD.n1501 GND 0.429674f
C3073 VDD.t67 GND 0.214837f
C3074 VDD.n1502 GND 0.006477f
C3075 VDD.n1503 GND 0.005213f
C3076 VDD.n1504 GND 0.006477f
C3077 VDD.n1505 GND 0.005213f
C3078 VDD.n1506 GND 0.006477f
C3079 VDD.n1507 GND 0.429674f
C3080 VDD.n1508 GND 0.006477f
C3081 VDD.n1509 GND 0.005213f
C3082 VDD.n1510 GND 0.006477f
C3083 VDD.n1511 GND 0.005213f
C3084 VDD.n1512 GND 0.006477f
C3085 VDD.n1513 GND 0.429674f
C3086 VDD.n1514 GND 0.006477f
C3087 VDD.n1515 GND 0.005213f
C3088 VDD.n1516 GND 0.006477f
C3089 VDD.n1517 GND 0.005213f
C3090 VDD.n1518 GND 0.006477f
C3091 VDD.n1519 GND 0.429674f
C3092 VDD.n1520 GND 0.006477f
C3093 VDD.n1521 GND 0.005213f
C3094 VDD.n1522 GND 0.006477f
C3095 VDD.n1523 GND 0.005213f
C3096 VDD.n1524 GND 0.006477f
C3097 VDD.n1525 GND 0.429674f
C3098 VDD.n1526 GND 0.006477f
C3099 VDD.n1527 GND 0.005213f
C3100 VDD.n1528 GND 0.006477f
C3101 VDD.n1529 GND 0.005213f
C3102 VDD.n1530 GND 0.006477f
C3103 VDD.t21 GND 0.214837f
C3104 VDD.n1531 GND 0.006477f
C3105 VDD.n1532 GND 0.005213f
C3106 VDD.n1533 GND 0.006477f
C3107 VDD.n1534 GND 0.005213f
C3108 VDD.n1535 GND 0.006477f
C3109 VDD.n1536 GND 0.429674f
C3110 VDD.n1537 GND 0.326552f
C3111 VDD.n1538 GND 0.006477f
C3112 VDD.n1539 GND 0.005213f
C3113 VDD.n1540 GND 0.006477f
C3114 VDD.n1541 GND 0.005213f
C3115 VDD.n1542 GND 0.006477f
C3116 VDD.n1543 GND 0.429674f
C3117 VDD.n1544 GND 0.006477f
C3118 VDD.n1545 GND 0.005213f
C3119 VDD.n1546 GND 0.006477f
C3120 VDD.n1547 GND 0.005213f
C3121 VDD.n1548 GND 0.006477f
C3122 VDD.n1549 GND 0.429674f
C3123 VDD.n1550 GND 0.006477f
C3124 VDD.n1551 GND 0.005213f
C3125 VDD.n1552 GND 0.006477f
C3126 VDD.n1553 GND 0.005213f
C3127 VDD.n1554 GND 0.006477f
C3128 VDD.n1555 GND 0.429674f
C3129 VDD.n1556 GND 0.006477f
C3130 VDD.n1557 GND 0.005213f
C3131 VDD.n1558 GND 0.006477f
C3132 VDD.n1559 GND 0.005213f
C3133 VDD.n1560 GND 0.006477f
C3134 VDD.n1561 GND 0.36952f
C3135 VDD.n1562 GND 0.006477f
C3136 VDD.n1563 GND 0.005213f
C3137 VDD.n1564 GND 0.006477f
C3138 VDD.n1565 GND 0.005213f
C3139 VDD.n1566 GND 0.006477f
C3140 VDD.n1567 GND 0.429674f
C3141 VDD.n1568 GND 0.006477f
C3142 VDD.n1569 GND 0.005213f
C3143 VDD.n1570 GND 0.006477f
C3144 VDD.n1571 GND 0.005213f
C3145 VDD.n1572 GND 0.006477f
C3146 VDD.n1573 GND 0.429674f
C3147 VDD.n1574 GND 0.006477f
C3148 VDD.n1575 GND 0.005213f
C3149 VDD.n1576 GND 0.006477f
C3150 VDD.n1577 GND 0.005213f
C3151 VDD.n1578 GND 0.006477f
C3152 VDD.n1579 GND 0.429674f
C3153 VDD.n1580 GND 0.006477f
C3154 VDD.n1581 GND 0.005213f
C3155 VDD.n1582 GND 0.006477f
C3156 VDD.n1583 GND 0.005213f
C3157 VDD.n1584 GND 0.006477f
C3158 VDD.n1585 GND 0.429674f
C3159 VDD.n1586 GND 0.006477f
C3160 VDD.n1587 GND 0.005213f
C3161 VDD.n1588 GND 0.006477f
C3162 VDD.n1589 GND 0.005213f
C3163 VDD.n1590 GND 0.006477f
C3164 VDD.n1591 GND 0.429674f
C3165 VDD.n1592 GND 0.006477f
C3166 VDD.n1593 GND 0.005213f
C3167 VDD.n1594 GND 0.006477f
C3168 VDD.n1595 GND 0.005213f
C3169 VDD.n1596 GND 0.006477f
C3170 VDD.n1597 GND 0.429674f
C3171 VDD.n1598 GND 0.006477f
C3172 VDD.n1599 GND 0.005213f
C3173 VDD.n1600 GND 0.006477f
C3174 VDD.n1601 GND 0.005213f
C3175 VDD.n1602 GND 0.006477f
C3176 VDD.n1603 GND 0.244914f
C3177 VDD.n1604 GND 0.006477f
C3178 VDD.n1605 GND 0.005213f
C3179 VDD.n1606 GND 0.006477f
C3180 VDD.n1607 GND 0.005213f
C3181 VDD.n1608 GND 0.006477f
C3182 VDD.n1609 GND 0.429674f
C3183 VDD.t86 GND 0.214837f
C3184 VDD.n1610 GND 0.006477f
C3185 VDD.n1611 GND 0.005213f
C3186 VDD.n1612 GND 0.006477f
C3187 VDD.n1613 GND 0.005213f
C3188 VDD.n1614 GND 0.006477f
C3189 VDD.n1615 GND 0.429674f
C3190 VDD.n1616 GND 0.006477f
C3191 VDD.n1617 GND 0.005213f
C3192 VDD.n1618 GND 0.014826f
C3193 VDD.n1619 GND 0.004327f
C3194 VDD.n1620 GND 0.014826f
C3195 VDD.n1621 GND 0.575763f
C3196 VDD.n1622 GND 0.014826f
C3197 VDD.n1623 GND 0.004327f
C3198 VDD.n1624 GND 0.006477f
C3199 VDD.n1625 GND 0.005213f
C3200 VDD.n1626 GND 0.006477f
C3201 VDD.n1640 GND 0.014967f
C3202 VDD.n1641 GND 0.006477f
C3203 VDD.n1642 GND 0.005213f
C3204 VDD.n1643 GND 0.006477f
C3205 VDD.n1644 GND 0.006477f
C3206 VDD.n1645 GND 0.006477f
C3207 VDD.n1646 GND 0.006477f
C3208 VDD.n1647 GND 0.006477f
C3209 VDD.n1648 GND 0.005213f
C3210 VDD.n1649 GND 0.006477f
C3211 VDD.n1650 GND 0.006477f
C3212 VDD.n1651 GND 0.006477f
C3213 VDD.n1652 GND 0.006477f
C3214 VDD.n1653 GND 0.006477f
C3215 VDD.n1654 GND 0.005213f
C3216 VDD.n1655 GND 0.006477f
C3217 VDD.n1656 GND 0.006477f
C3218 VDD.n1657 GND 0.006477f
C3219 VDD.n1658 GND 0.006477f
C3220 VDD.n1659 GND 0.005213f
C3221 VDD.n1660 GND 0.006477f
C3222 VDD.n1661 GND 0.006477f
C3223 VDD.n1662 GND 0.006477f
C3224 VDD.n1663 GND 0.006477f
C3225 VDD.n1664 GND 0.006477f
C3226 VDD.n1665 GND 0.005213f
C3227 VDD.n1666 GND 0.006477f
C3228 VDD.n1667 GND 0.006477f
C3229 VDD.n1668 GND 0.006477f
C3230 VDD.n1669 GND 0.006477f
C3231 VDD.n1670 GND 0.006477f
C3232 VDD.n1671 GND 0.005213f
C3233 VDD.n1672 GND 0.006477f
C3234 VDD.n1673 GND 0.006477f
C3235 VDD.n1674 GND 0.006477f
C3236 VDD.n1675 GND 0.006477f
C3237 VDD.n1676 GND 0.006477f
C3238 VDD.n1677 GND 0.005213f
C3239 VDD.n1678 GND 0.014967f
C3240 VDD.n1679 GND 0.006477f
C3241 VDD.n1680 GND 0.002502f
C3242 VDD.t101 GND 0.086094f
C3243 VDD.t102 GND 0.107631f
C3244 VDD.t100 GND 0.799934f
C3245 VDD.n1681 GND 0.078348f
C3246 VDD.n1682 GND 0.048083f
C3247 VDD.n1683 GND 0.008028f
C3248 VDD.n1684 GND 0.002711f
C3249 VDD.n1685 GND 0.006477f
C3250 VDD.n1686 GND 0.006477f
C3251 VDD.n1687 GND 0.006477f
C3252 VDD.n1688 GND 0.005213f
C3253 VDD.n1689 GND 0.005213f
C3254 VDD.n1690 GND 0.005213f
C3255 VDD.n1691 GND 0.006477f
C3256 VDD.n1692 GND 0.006477f
C3257 VDD.n1693 GND 0.006477f
C3258 VDD.n1694 GND 0.005213f
C3259 VDD.n1695 GND 0.005213f
C3260 VDD.n1696 GND 0.005213f
C3261 VDD.n1697 GND 0.006477f
C3262 VDD.n1698 GND 0.006477f
C3263 VDD.n1699 GND 0.006477f
C3264 VDD.n1700 GND 0.005213f
C3265 VDD.n1701 GND 0.005213f
C3266 VDD.n1702 GND 0.005213f
C3267 VDD.n1703 GND 0.006477f
C3268 VDD.n1704 GND 0.006477f
C3269 VDD.n1705 GND 0.006477f
C3270 VDD.n1706 GND 0.004744f
C3271 VDD.n1707 GND 0.006477f
C3272 VDD.t87 GND 0.086094f
C3273 VDD.t88 GND 0.107631f
C3274 VDD.t85 GND 0.799934f
C3275 VDD.n1708 GND 0.078348f
C3276 VDD.n1709 GND 0.048083f
C3277 VDD.n1710 GND 0.010634f
C3278 VDD.n1711 GND 0.003962f
C3279 VDD.n1712 GND 0.006477f
C3280 VDD.n1713 GND 0.006477f
C3281 VDD.n1714 GND 0.006477f
C3282 VDD.n1715 GND 0.005213f
C3283 VDD.n1716 GND 0.005213f
C3284 VDD.n1717 GND 0.005213f
C3285 VDD.n1718 GND 0.006477f
C3286 VDD.n1719 GND 0.006477f
C3287 VDD.n1720 GND 0.006477f
C3288 VDD.n1721 GND 0.005213f
C3289 VDD.n1722 GND 0.005213f
C3290 VDD.n1723 GND 0.005213f
C3291 VDD.n1724 GND 0.006477f
C3292 VDD.n1725 GND 0.006477f
C3293 VDD.n1726 GND 0.006477f
C3294 VDD.n1727 GND 0.005213f
C3295 VDD.n1728 GND 0.006477f
C3296 VDD.n1729 GND 0.966767f
C3297 VDD.n1731 GND 0.014967f
C3298 VDD.n1732 GND 0.004327f
C3299 VDD.n1733 GND 0.014967f
C3300 VDD.n1734 GND 0.014826f
C3301 VDD.n1735 GND 0.006477f
C3302 VDD.n1736 GND 0.005213f
C3303 VDD.n1737 GND 0.006477f
C3304 VDD.n1738 GND 0.429674f
C3305 VDD.n1739 GND 0.006477f
C3306 VDD.n1740 GND 0.005213f
C3307 VDD.n1741 GND 0.006477f
C3308 VDD.n1742 GND 0.006477f
C3309 VDD.n1743 GND 0.006477f
C3310 VDD.n1744 GND 0.005213f
C3311 VDD.n1745 GND 0.006477f
C3312 VDD.n1746 GND 0.429674f
C3313 VDD.n1747 GND 0.006477f
C3314 VDD.n1748 GND 0.005213f
C3315 VDD.n1749 GND 0.006477f
C3316 VDD.n1750 GND 0.006477f
C3317 VDD.n1751 GND 0.006477f
C3318 VDD.n1752 GND 0.005213f
C3319 VDD.n1753 GND 0.006477f
C3320 VDD.n1754 GND 0.399597f
C3321 VDD.n1755 GND 0.006477f
C3322 VDD.n1756 GND 0.005213f
C3323 VDD.n1757 GND 0.006477f
C3324 VDD.n1758 GND 0.006477f
C3325 VDD.n1759 GND 0.006477f
C3326 VDD.n1760 GND 0.005213f
C3327 VDD.n1761 GND 0.006477f
C3328 VDD.n1762 GND 0.429674f
C3329 VDD.n1763 GND 0.006477f
C3330 VDD.n1764 GND 0.005213f
C3331 VDD.n1765 GND 0.006477f
C3332 VDD.n1766 GND 0.006477f
C3333 VDD.n1767 GND 0.006477f
C3334 VDD.n1768 GND 0.005213f
C3335 VDD.n1769 GND 0.006477f
C3336 VDD.n1770 GND 0.429674f
C3337 VDD.n1771 GND 0.006477f
C3338 VDD.n1772 GND 0.005213f
C3339 VDD.n1773 GND 0.006477f
C3340 VDD.n1774 GND 0.006477f
C3341 VDD.n1775 GND 0.006477f
C3342 VDD.n1776 GND 0.005213f
C3343 VDD.n1777 GND 0.006477f
C3344 VDD.n1778 GND 0.429674f
C3345 VDD.n1779 GND 0.006477f
C3346 VDD.n1780 GND 0.005213f
C3347 VDD.n1781 GND 0.006477f
C3348 VDD.n1782 GND 0.006477f
C3349 VDD.n1783 GND 0.006477f
C3350 VDD.n1784 GND 0.005213f
C3351 VDD.n1785 GND 0.006477f
C3352 VDD.n1786 GND 0.429674f
C3353 VDD.n1787 GND 0.006477f
C3354 VDD.n1788 GND 0.005213f
C3355 VDD.n1789 GND 0.006477f
C3356 VDD.n1790 GND 0.006477f
C3357 VDD.n1791 GND 0.006477f
C3358 VDD.n1792 GND 0.005213f
C3359 VDD.n1793 GND 0.006477f
C3360 VDD.n1794 GND 0.429674f
C3361 VDD.n1795 GND 0.006477f
C3362 VDD.n1796 GND 0.005213f
C3363 VDD.n1797 GND 0.006477f
C3364 VDD.n1798 GND 0.006477f
C3365 VDD.n1799 GND 0.006477f
C3366 VDD.n1800 GND 0.005213f
C3367 VDD.n1801 GND 0.006477f
C3368 VDD.n1802 GND 0.429674f
C3369 VDD.n1803 GND 0.006477f
C3370 VDD.n1804 GND 0.005213f
C3371 VDD.n1805 GND 0.006477f
C3372 VDD.n1806 GND 0.006477f
C3373 VDD.n1807 GND 0.006477f
C3374 VDD.n1808 GND 0.005213f
C3375 VDD.n1809 GND 0.006477f
C3376 VDD.t54 GND 0.214837f
C3377 VDD.n1810 GND 0.274991f
C3378 VDD.n1811 GND 0.006477f
C3379 VDD.n1812 GND 0.005213f
C3380 VDD.n1813 GND 0.006477f
C3381 VDD.n1814 GND 0.006477f
C3382 VDD.n1815 GND 0.006477f
C3383 VDD.n1816 GND 0.005213f
C3384 VDD.n1817 GND 0.006477f
C3385 VDD.n1818 GND 0.429674f
C3386 VDD.n1819 GND 0.006477f
C3387 VDD.n1820 GND 0.005213f
C3388 VDD.n1821 GND 0.006477f
C3389 VDD.n1822 GND 0.006477f
C3390 VDD.n1823 GND 0.006477f
C3391 VDD.n1824 GND 0.005213f
C3392 VDD.n1825 GND 0.006477f
C3393 VDD.n1826 GND 0.429674f
C3394 VDD.n1827 GND 0.006477f
C3395 VDD.n1828 GND 0.005213f
C3396 VDD.n1829 GND 0.006477f
C3397 VDD.n1830 GND 0.006477f
C3398 VDD.n1831 GND 0.006477f
C3399 VDD.n1832 GND 0.005213f
C3400 VDD.n1833 GND 0.006477f
C3401 VDD.n1834 GND 0.429674f
C3402 VDD.n1835 GND 0.006477f
C3403 VDD.n1836 GND 0.005213f
C3404 VDD.n1837 GND 0.006477f
C3405 VDD.n1838 GND 0.006477f
C3406 VDD.n1839 GND 0.006477f
C3407 VDD.n1840 GND 0.005213f
C3408 VDD.n1841 GND 0.006477f
C3409 VDD.n1842 GND 0.429674f
C3410 VDD.n1843 GND 0.006477f
C3411 VDD.n1844 GND 0.005213f
C3412 VDD.n1845 GND 0.006477f
C3413 VDD.n1846 GND 0.006477f
C3414 VDD.n1847 GND 0.006477f
C3415 VDD.n1848 GND 0.005213f
C3416 VDD.n1849 GND 0.006477f
C3417 VDD.n1850 GND 0.429674f
C3418 VDD.n1851 GND 0.006477f
C3419 VDD.n1852 GND 0.005213f
C3420 VDD.n1853 GND 0.006477f
C3421 VDD.n1854 GND 0.006477f
C3422 VDD.n1855 GND 0.006477f
C3423 VDD.n1856 GND 0.005213f
C3424 VDD.n1857 GND 0.006477f
C3425 VDD.n1858 GND 0.317959f
C3426 VDD.n1859 GND 0.006477f
C3427 VDD.n1860 GND 0.005213f
C3428 VDD.n1861 GND 0.006477f
C3429 VDD.n1862 GND 0.006477f
C3430 VDD.n1863 GND 0.006477f
C3431 VDD.n1864 GND 0.005213f
C3432 VDD.n1865 GND 0.006477f
C3433 VDD.n1866 GND 0.429674f
C3434 VDD.n1867 GND 0.006477f
C3435 VDD.n1868 GND 0.005213f
C3436 VDD.n1869 GND 0.006477f
C3437 VDD.n1870 GND 0.006477f
C3438 VDD.n1871 GND 0.006477f
C3439 VDD.n1872 GND 0.005213f
C3440 VDD.n1873 GND 0.006477f
C3441 VDD.n1874 GND 0.429674f
C3442 VDD.n1875 GND 0.006477f
C3443 VDD.n1876 GND 0.005213f
C3444 VDD.n1877 GND 0.006477f
C3445 VDD.n1878 GND 0.006477f
C3446 VDD.n1879 GND 0.006477f
C3447 VDD.n1880 GND 0.005213f
C3448 VDD.n1881 GND 0.006477f
C3449 VDD.n1882 GND 0.429674f
C3450 VDD.n1883 GND 0.006477f
C3451 VDD.n1884 GND 0.005213f
C3452 VDD.n1885 GND 0.006477f
C3453 VDD.n1886 GND 0.006477f
C3454 VDD.n1887 GND 0.006477f
C3455 VDD.n1888 GND 0.005213f
C3456 VDD.n1889 GND 0.006477f
C3457 VDD.n1890 GND 0.429674f
C3458 VDD.n1891 GND 0.006477f
C3459 VDD.n1892 GND 0.005213f
C3460 VDD.n1893 GND 0.006477f
C3461 VDD.n1894 GND 0.006477f
C3462 VDD.n1895 GND 0.006477f
C3463 VDD.n1896 GND 0.005213f
C3464 VDD.n1897 GND 0.006477f
C3465 VDD.n1898 GND 0.378113f
C3466 VDD.n1899 GND 0.006477f
C3467 VDD.n1900 GND 0.005213f
C3468 VDD.n1901 GND 0.006477f
C3469 VDD.n1902 GND 0.006477f
C3470 VDD.n1903 GND 0.006477f
C3471 VDD.n1904 GND 0.005213f
C3472 VDD.n1905 GND 0.006477f
C3473 VDD.n1906 GND 0.429674f
C3474 VDD.n1907 GND 0.006477f
C3475 VDD.n1908 GND 0.005213f
C3476 VDD.n1909 GND 0.006477f
C3477 VDD.n1910 GND 0.006477f
C3478 VDD.n1911 GND 0.006477f
C3479 VDD.n1912 GND 0.005213f
C3480 VDD.n1913 GND 0.006477f
C3481 VDD.n1914 GND 0.429674f
C3482 VDD.n1915 GND 0.006477f
C3483 VDD.n1916 GND 0.005213f
C3484 VDD.n1917 GND 0.006477f
C3485 VDD.n1918 GND 0.006477f
C3486 VDD.n1919 GND 0.006477f
C3487 VDD.n1920 GND 0.005213f
C3488 VDD.n1921 GND 0.006477f
C3489 VDD.n1922 GND 0.429674f
C3490 VDD.n1923 GND 0.006477f
C3491 VDD.n1924 GND 0.005213f
C3492 VDD.n1925 GND 0.006477f
C3493 VDD.n1926 GND 0.006477f
C3494 VDD.n1927 GND 0.006477f
C3495 VDD.n1928 GND 0.005213f
C3496 VDD.n1929 GND 0.006477f
C3497 VDD.n1930 GND 0.429674f
C3498 VDD.n1931 GND 0.006477f
C3499 VDD.n1932 GND 0.005213f
C3500 VDD.n1933 GND 0.006477f
C3501 VDD.n1934 GND 0.006477f
C3502 VDD.n1935 GND 0.006477f
C3503 VDD.n1936 GND 0.005213f
C3504 VDD.n1937 GND 0.006477f
C3505 VDD.n1938 GND 0.429674f
C3506 VDD.n1939 GND 0.006477f
C3507 VDD.n1940 GND 0.005213f
C3508 VDD.n1941 GND 0.006477f
C3509 VDD.n1942 GND 0.006454f
C3510 VDD.t70 GND 0.106353f
C3511 VDD.t141 GND 0.012824f
C3512 VDD.t71 GND 0.012824f
C3513 VDD.n1943 GND 0.07391f
C3514 VDD.n1944 GND 0.421202f
C3515 VDD.t68 GND 0.012824f
C3516 VDD.t27 GND 0.012824f
C3517 VDD.n1945 GND 0.07391f
C3518 VDD.n1946 GND 0.259498f
C3519 VDD.t139 GND 0.012824f
C3520 VDD.t72 GND 0.012824f
C3521 VDD.n1947 GND 0.07391f
C3522 VDD.n1948 GND 0.285563f
C3523 VDD.t129 GND 0.106353f
C3524 VDD.t53 GND 0.012824f
C3525 VDD.t64 GND 0.012824f
C3526 VDD.n1949 GND 0.07391f
C3527 VDD.n1950 GND 0.421202f
C3528 VDD.t133 GND 0.012824f
C3529 VDD.t138 GND 0.012824f
C3530 VDD.n1951 GND 0.07391f
C3531 VDD.n1952 GND 0.259498f
C3532 VDD.t55 GND 0.012824f
C3533 VDD.t22 GND 0.012824f
C3534 VDD.n1953 GND 0.07391f
C3535 VDD.n1954 GND 0.265639f
C3536 VDD.n1955 GND 0.388246f
C3537 VDD.n1956 GND 3.33641f
C3538 VDD.n1957 GND 0.46472f
C3539 VDD.n1958 GND 0.005213f
C3540 VDD.n1959 GND 0.006477f
C3541 VDD.t26 GND 0.429674f
C3542 VDD.n1960 GND 0.006477f
C3543 VDD.n1961 GND 0.005213f
C3544 VDD.n1962 GND 0.006477f
C3545 VDD.n1963 GND 0.006477f
C3546 VDD.n1964 GND 0.006477f
C3547 VDD.n1965 GND 0.005213f
C3548 VDD.n1966 GND 0.006477f
C3549 VDD.n1967 GND 0.429674f
C3550 VDD.n1968 GND 0.006477f
C3551 VDD.n1969 GND 0.005213f
C3552 VDD.n1970 GND 0.006477f
C3553 VDD.n1971 GND 0.006477f
C3554 VDD.n1972 GND 0.006477f
C3555 VDD.n1973 GND 0.005213f
C3556 VDD.n1974 GND 0.006477f
C3557 VDD.n1975 GND 0.429674f
C3558 VDD.n1976 GND 0.006477f
C3559 VDD.n1977 GND 0.005213f
C3560 VDD.n1978 GND 0.006477f
C3561 VDD.n1979 GND 0.006477f
C3562 VDD.n1980 GND 0.006477f
C3563 VDD.n1981 GND 0.005213f
C3564 VDD.n1982 GND 0.006477f
C3565 VDD.n1983 GND 0.429674f
C3566 VDD.n1984 GND 0.006477f
C3567 VDD.n1985 GND 0.005213f
C3568 VDD.n1986 GND 0.006477f
C3569 VDD.n1987 GND 0.006477f
C3570 VDD.n1988 GND 0.006477f
C3571 VDD.n1989 GND 0.005213f
C3572 VDD.n1990 GND 0.006477f
C3573 VDD.n1991 GND 0.429674f
C3574 VDD.n1992 GND 0.006477f
C3575 VDD.n1993 GND 0.005213f
C3576 VDD.n1994 GND 0.006477f
C3577 VDD.n1995 GND 0.006477f
C3578 VDD.n1996 GND 0.006477f
C3579 VDD.n1997 GND 0.005213f
C3580 VDD.n1998 GND 0.006477f
C3581 VDD.n1999 GND 0.266398f
C3582 VDD.n2000 GND 0.429674f
C3583 VDD.n2001 GND 0.006477f
C3584 VDD.n2002 GND 0.005213f
C3585 VDD.n2003 GND 0.006477f
C3586 VDD.n2004 GND 0.006477f
C3587 VDD.n2005 GND 0.006477f
C3588 VDD.n2006 GND 0.005213f
C3589 VDD.n2007 GND 0.006477f
C3590 VDD.n2008 GND 0.378113f
C3591 VDD.n2009 GND 0.006477f
C3592 VDD.n2010 GND 0.005213f
C3593 VDD.n2011 GND 0.006477f
C3594 VDD.n2012 GND 0.006477f
C3595 VDD.n2013 GND 0.006477f
C3596 VDD.n2014 GND 0.005213f
C3597 VDD.n2015 GND 0.006477f
C3598 VDD.n2016 GND 0.429674f
C3599 VDD.n2017 GND 0.006477f
C3600 VDD.n2018 GND 0.005213f
C3601 VDD.n2019 GND 0.006477f
C3602 VDD.n2020 GND 0.006477f
C3603 VDD.n2021 GND 0.006477f
C3604 VDD.n2022 GND 0.005213f
C3605 VDD.n2023 GND 0.006477f
C3606 VDD.n2024 GND 0.429674f
C3607 VDD.n2025 GND 0.006477f
C3608 VDD.n2026 GND 0.005213f
C3609 VDD.n2027 GND 0.006477f
C3610 VDD.n2028 GND 0.006477f
C3611 VDD.n2029 GND 0.006477f
C3612 VDD.n2030 GND 0.005213f
C3613 VDD.n2031 GND 0.006477f
C3614 VDD.n2032 GND 0.429674f
C3615 VDD.n2033 GND 0.006477f
C3616 VDD.n2034 GND 0.005213f
C3617 VDD.n2035 GND 0.006477f
C3618 VDD.n2036 GND 0.006477f
C3619 VDD.n2037 GND 0.006477f
C3620 VDD.n2038 GND 0.005213f
C3621 VDD.n2039 GND 0.006477f
C3622 VDD.n2040 GND 0.429674f
C3623 VDD.n2041 GND 0.006477f
C3624 VDD.n2042 GND 0.005213f
C3625 VDD.n2043 GND 0.006477f
C3626 VDD.n2044 GND 0.006477f
C3627 VDD.n2045 GND 0.006477f
C3628 VDD.n2046 GND 0.005213f
C3629 VDD.n2047 GND 0.006477f
C3630 VDD.t63 GND 0.214837f
C3631 VDD.n2048 GND 0.317959f
C3632 VDD.n2049 GND 0.006477f
C3633 VDD.n2050 GND 0.005213f
C3634 VDD.n2051 GND 0.006477f
C3635 VDD.n2052 GND 0.006477f
C3636 VDD.n2053 GND 0.006477f
C3637 VDD.n2054 GND 0.005213f
C3638 VDD.n2055 GND 0.006477f
C3639 VDD.n2056 GND 0.429674f
C3640 VDD.n2057 GND 0.006477f
C3641 VDD.n2058 GND 0.005213f
C3642 VDD.n2059 GND 0.006477f
C3643 VDD.n2060 GND 0.006477f
C3644 VDD.n2061 GND 0.006477f
C3645 VDD.n2062 GND 0.005213f
C3646 VDD.n2063 GND 0.006477f
C3647 VDD.n2064 GND 0.429674f
C3648 VDD.n2065 GND 0.006477f
C3649 VDD.n2066 GND 0.005213f
C3650 VDD.n2067 GND 0.006477f
C3651 VDD.n2068 GND 0.006477f
C3652 VDD.n2069 GND 0.006477f
C3653 VDD.n2070 GND 0.005213f
C3654 VDD.n2071 GND 0.006477f
C3655 VDD.n2072 GND 0.429674f
C3656 VDD.n2073 GND 0.006477f
C3657 VDD.n2074 GND 0.005213f
C3658 VDD.n2075 GND 0.006477f
C3659 VDD.n2076 GND 0.006477f
C3660 VDD.n2077 GND 0.006477f
C3661 VDD.n2078 GND 0.005213f
C3662 VDD.n2079 GND 0.006477f
C3663 VDD.n2080 GND 0.429674f
C3664 VDD.n2081 GND 0.006477f
C3665 VDD.n2082 GND 0.005213f
C3666 VDD.n2083 GND 0.006477f
C3667 VDD.n2084 GND 0.006477f
C3668 VDD.n2085 GND 0.006477f
C3669 VDD.n2086 GND 0.005213f
C3670 VDD.n2087 GND 0.006477f
C3671 VDD.n2088 GND 0.429674f
C3672 VDD.n2089 GND 0.006477f
C3673 VDD.n2090 GND 0.005213f
C3674 VDD.n2091 GND 0.006477f
C3675 VDD.n2092 GND 0.006477f
C3676 VDD.n2093 GND 0.006477f
C3677 VDD.n2094 GND 0.005213f
C3678 VDD.n2095 GND 0.006477f
C3679 VDD.n2096 GND 0.274991f
C3680 VDD.n2097 GND 0.006477f
C3681 VDD.n2098 GND 0.005213f
C3682 VDD.n2099 GND 0.006477f
C3683 VDD.n2100 GND 0.006477f
C3684 VDD.n2101 GND 0.006477f
C3685 VDD.n2102 GND 0.005213f
C3686 VDD.n2103 GND 0.006477f
C3687 VDD.n2104 GND 0.429674f
C3688 VDD.n2105 GND 0.006477f
C3689 VDD.n2106 GND 0.005213f
C3690 VDD.n2107 GND 0.006477f
C3691 VDD.n2108 GND 0.006477f
C3692 VDD.n2109 GND 0.006477f
C3693 VDD.n2110 GND 0.005213f
C3694 VDD.n2111 GND 0.006477f
C3695 VDD.n2112 GND 0.429674f
C3696 VDD.n2113 GND 0.006477f
C3697 VDD.n2114 GND 0.005213f
C3698 VDD.n2115 GND 0.006477f
C3699 VDD.n2116 GND 0.006477f
C3700 VDD.n2117 GND 0.006477f
C3701 VDD.n2118 GND 0.005213f
C3702 VDD.n2119 GND 0.006477f
C3703 VDD.n2120 GND 0.429674f
C3704 VDD.n2121 GND 0.006477f
C3705 VDD.n2122 GND 0.005213f
C3706 VDD.n2123 GND 0.006477f
C3707 VDD.n2124 GND 0.006477f
C3708 VDD.n2125 GND 0.006477f
C3709 VDD.n2126 GND 0.005213f
C3710 VDD.n2127 GND 0.006477f
C3711 VDD.n2128 GND 0.429674f
C3712 VDD.n2129 GND 0.006477f
C3713 VDD.n2130 GND 0.005213f
C3714 VDD.n2131 GND 0.006477f
C3715 VDD.n2132 GND 0.006477f
C3716 VDD.n2133 GND 0.006477f
C3717 VDD.n2134 GND 0.005213f
C3718 VDD.n2135 GND 0.006477f
C3719 VDD.n2136 GND 0.429674f
C3720 VDD.n2137 GND 0.006477f
C3721 VDD.n2138 GND 0.005213f
C3722 VDD.n2139 GND 0.006477f
C3723 VDD.n2140 GND 0.006477f
C3724 VDD.n2141 GND 0.006477f
C3725 VDD.n2142 GND 0.006477f
C3726 VDD.n2143 GND 0.005213f
C3727 VDD.n2144 GND 0.006477f
C3728 VDD.n2145 GND 0.244914f
C3729 VDD.n2146 GND 0.429674f
C3730 VDD.n2147 GND 0.006477f
C3731 VDD.n2148 GND 0.005213f
C3732 VDD.n2149 GND 0.006477f
C3733 VDD.n2150 GND 0.006477f
C3734 VDD.n2151 GND 0.006477f
C3735 VDD.n2152 GND 0.005213f
C3736 VDD.n2153 GND 0.006477f
C3737 VDD.n2154 GND 0.399597f
C3738 VDD.n2155 GND 0.006477f
C3739 VDD.n2156 GND 0.006477f
C3740 VDD.n2157 GND 0.005213f
C3741 VDD.n2158 GND 0.006477f
C3742 VDD.n2159 GND 0.006477f
C3743 VDD.n2160 GND 0.01038f
C3744 VDD.n2161 GND 0.01038f
C3745 VDD.n2162 GND 0.004404f
C3746 VDD.n2163 GND 0.004404f
C3747 VDD.n2164 GND 0.004404f
C3748 VDD.n2165 GND 0.004404f
C3749 VDD.n2166 GND 0.004404f
C3750 VDD.n2167 GND 0.004404f
C3751 VDD.n2168 GND 0.004404f
C3752 VDD.n2169 GND 0.004404f
C3753 VDD.n2170 GND 0.004404f
C3754 VDD.n2171 GND 0.004404f
C3755 VDD.n2172 GND 0.004404f
C3756 VDD.n2173 GND 0.004404f
C3757 VDD.n2174 GND 0.004404f
C3758 VDD.n2175 GND 0.004404f
C3759 VDD.n2176 GND 0.004404f
C3760 VDD.n2177 GND 0.004404f
C3761 VDD.n2178 GND 0.003303f
C3762 VDD.t121 GND 0.068381f
C3763 VDD.t122 GND 0.084764f
C3764 VDD.t119 GND 0.489916f
C3765 VDD.n2179 GND 0.064611f
C3766 VDD.n2180 GND 0.042608f
C3767 VDD.n2181 GND 0.004404f
C3768 VDD.n2182 GND 0.004404f
C3769 VDD.n2183 GND 0.004404f
C3770 VDD.n2184 GND 0.004404f
C3771 VDD.n2185 GND 0.004404f
C3772 VDD.n2186 GND 0.004404f
C3773 VDD.n2187 GND 0.004404f
C3774 VDD.n2188 GND 0.004404f
C3775 VDD.n2189 GND 0.004404f
C3776 VDD.n2190 GND 0.004404f
C3777 VDD.n2191 GND 0.004404f
C3778 VDD.n2192 GND 0.004404f
C3779 VDD.n2193 GND 0.004404f
C3780 VDD.n2194 GND 0.004404f
C3781 VDD.n2195 GND 0.004404f
C3782 VDD.n2196 GND 0.004404f
C3783 VDD.n2197 GND 0.004404f
C3784 VDD.n2198 GND 0.004404f
C3785 VDD.n2199 GND 0.004404f
C3786 VDD.n2200 GND 0.004404f
C3787 VDD.n2201 GND 0.004404f
C3788 VDD.n2202 GND 0.004404f
C3789 VDD.n2203 GND 0.004404f
C3790 VDD.n2204 GND 0.004404f
C3791 VDD.n2205 GND 0.004404f
C3792 VDD.n2206 GND 0.004404f
C3793 VDD.n2207 GND 0.004404f
C3794 VDD.n2208 GND 0.004404f
C3795 VDD.n2209 GND 0.004404f
C3796 VDD.n2210 GND 0.004404f
C3797 VDD.n2211 GND 0.004404f
C3798 VDD.n2212 GND 0.004404f
C3799 VDD.n2213 GND 0.004404f
C3800 VDD.n2214 GND 0.004404f
C3801 VDD.n2215 GND 0.004404f
C3802 VDD.n2216 GND 0.004404f
C3803 VDD.n2217 GND 0.004404f
C3804 VDD.n2218 GND 0.004404f
C3805 VDD.n2219 GND 0.004404f
C3806 VDD.n2220 GND 0.004404f
C3807 VDD.n2221 GND 0.004404f
C3808 VDD.n2222 GND 0.004404f
C3809 VDD.n2223 GND 0.004404f
C3810 VDD.n2224 GND 0.004404f
C3811 VDD.n2225 GND 0.004404f
C3812 VDD.n2226 GND 0.004404f
C3813 VDD.n2227 GND 0.004404f
C3814 VDD.n2228 GND 0.004404f
C3815 VDD.n2229 GND 0.004404f
C3816 VDD.n2230 GND 0.004404f
C3817 VDD.n2231 GND 0.004404f
C3818 VDD.n2232 GND 0.004404f
C3819 VDD.n2233 GND 0.004404f
C3820 VDD.n2234 GND 0.004404f
C3821 VDD.n2235 GND 0.004404f
C3822 VDD.n2236 GND 0.004404f
C3823 VDD.n2237 GND 0.004404f
C3824 VDD.n2238 GND 0.004404f
C3825 VDD.n2239 GND 0.004404f
C3826 VDD.n2240 GND 0.004404f
C3827 VDD.n2241 GND 0.004404f
C3828 VDD.n2242 GND 0.004404f
C3829 VDD.n2243 GND 0.004404f
C3830 VDD.n2244 GND 0.004404f
C3831 VDD.n2245 GND 0.004404f
C3832 VDD.n2246 GND 0.004404f
C3833 VDD.n2247 GND 0.004404f
C3834 VDD.n2248 GND 0.004404f
C3835 VDD.n2249 GND 0.004404f
C3836 VDD.n2250 GND 0.004404f
C3837 VDD.n2251 GND 0.004404f
C3838 VDD.n2252 GND 0.004404f
C3839 VDD.n2253 GND 0.004404f
C3840 VDD.n2254 GND 0.004404f
C3841 VDD.n2255 GND 0.004404f
C3842 VDD.n2256 GND 0.004404f
C3843 VDD.n2257 GND 0.004404f
C3844 VDD.n2258 GND 0.004404f
C3845 VDD.n2259 GND 0.004404f
C3846 VDD.n2260 GND 0.004404f
C3847 VDD.n2261 GND 0.004404f
C3848 VDD.n2262 GND 0.004404f
C3849 VDD.n2263 GND 0.004404f
C3850 VDD.n2264 GND 0.004404f
C3851 VDD.n2265 GND 0.004404f
C3852 VDD.n2266 GND 0.004404f
C3853 VDD.n2267 GND 0.004404f
C3854 VDD.n2268 GND 0.004404f
C3855 VDD.n2269 GND 0.004404f
C3856 VDD.n2270 GND 0.004404f
C3857 VDD.n2271 GND 0.004404f
C3858 VDD.n2272 GND 0.004404f
C3859 VDD.n2273 GND 0.004404f
C3860 VDD.n2274 GND 0.004404f
C3861 VDD.n2275 GND 0.004404f
C3862 VDD.n2276 GND 0.004404f
C3863 VDD.n2277 GND 0.004404f
C3864 VDD.n2278 GND 0.004404f
C3865 VDD.n2279 GND 0.004404f
C3866 VDD.n2280 GND 0.004404f
C3867 VDD.n2281 GND 0.004404f
C3868 VDD.n2282 GND 0.004404f
C3869 VDD.n2283 GND 0.004404f
C3870 VDD.n2284 GND 0.004404f
C3871 VDD.n2285 GND 0.004404f
C3872 VDD.n2286 GND 0.004404f
C3873 VDD.n2287 GND 0.004404f
C3874 VDD.n2288 GND 0.004404f
C3875 VDD.n2289 GND 0.004404f
C3876 VDD.n2290 GND 0.004404f
C3877 VDD.n2291 GND 0.004404f
C3878 VDD.n2292 GND 0.004404f
C3879 VDD.n2293 GND 0.004404f
C3880 VDD.n2294 GND 0.004404f
C3881 VDD.n2295 GND 0.004404f
C3882 VDD.n2296 GND 0.004404f
C3883 VDD.n2297 GND 0.004404f
C3884 VDD.n2298 GND 0.004404f
C3885 VDD.n2299 GND 0.004404f
C3886 VDD.n2300 GND 0.004404f
C3887 VDD.n2301 GND 0.004404f
C3888 VDD.n2302 GND 0.004404f
C3889 VDD.n2303 GND 0.004404f
C3890 VDD.n2304 GND 0.004404f
C3891 VDD.n2305 GND 0.004404f
C3892 VDD.n2306 GND 0.004404f
C3893 VDD.n2307 GND 0.004404f
C3894 VDD.t127 GND 0.068381f
C3895 VDD.t128 GND 0.084764f
C3896 VDD.t126 GND 0.489916f
C3897 VDD.n2308 GND 0.064611f
C3898 VDD.n2309 GND 0.042608f
C3899 VDD.n2310 GND 0.006294f
C3900 VDD.n2311 GND 0.004404f
C3901 VDD.n2312 GND 0.004404f
C3902 VDD.n2313 GND 0.004404f
C3903 VDD.n2314 GND 0.004404f
C3904 VDD.n2315 GND 0.004404f
C3905 VDD.n2316 GND 0.004404f
C3906 VDD.n2317 GND 0.004404f
C3907 VDD.n2318 GND 0.004404f
C3908 VDD.n2319 GND 0.004404f
C3909 VDD.n2320 GND 0.004404f
C3910 VDD.n2321 GND 0.004404f
C3911 VDD.n2322 GND 0.003854f
C3912 VDD.n2323 GND 0.004404f
C3913 VDD.n2324 GND 0.004404f
C3914 VDD.n2325 GND 0.002753f
C3915 VDD.n2326 GND 0.004404f
C3916 VDD.n2327 GND 0.004404f
C3917 VDD.n2328 GND 0.01038f
C3918 VDD.n2329 GND 0.010151f
C3919 VDD.n2330 GND 0.010151f
C3920 VDD.n2331 GND 0.004404f
C3921 VDD.n2332 GND 0.004404f
C3922 VDD.n2333 GND 0.004404f
C3923 VDD.n2334 GND 0.004404f
C3924 VDD.n2335 GND 0.004404f
C3925 VDD.n2336 GND 0.004404f
C3926 VDD.n2337 GND 0.004404f
C3927 VDD.n2338 GND 0.004404f
C3928 VDD.n2339 GND 0.004404f
C3929 VDD.n2340 GND 0.004404f
C3930 VDD.n2341 GND 0.004404f
C3931 VDD.n2342 GND 0.004404f
C3932 VDD.n2343 GND 0.004404f
C3933 VDD.n2344 GND 0.004404f
C3934 VDD.n2345 GND 0.004404f
C3935 VDD.n2346 GND 0.004404f
C3936 VDD.n2347 GND 0.004404f
C3937 VDD.n2348 GND 0.004404f
C3938 VDD.n2349 GND 0.004404f
C3939 VDD.n2350 GND 0.004404f
C3940 VDD.n2351 GND 0.004404f
C3941 VDD.n2352 GND 0.004404f
C3942 VDD.n2353 GND 0.004404f
C3943 VDD.n2354 GND 0.004404f
C3944 VDD.n2355 GND 0.004404f
C3945 VDD.n2356 GND 0.004404f
C3946 VDD.n2357 GND 0.004404f
C3947 VDD.n2358 GND 0.004404f
C3948 VDD.n2359 GND 0.004404f
C3949 VDD.n2360 GND 0.004404f
C3950 VDD.n2361 GND 0.004404f
C3951 VDD.n2362 GND 0.004404f
C3952 VDD.n2363 GND 0.004404f
C3953 VDD.n2364 GND 0.004404f
C3954 VDD.n2365 GND 0.004404f
C3955 VDD.n2366 GND 0.004404f
C3956 VDD.n2367 GND 0.004404f
C3957 VDD.n2368 GND 0.004404f
C3958 VDD.n2369 GND 0.004404f
C3959 VDD.n2370 GND 0.004404f
C3960 VDD.n2371 GND 0.004404f
C3961 VDD.n2372 GND 0.004404f
C3962 VDD.n2373 GND 0.004404f
C3963 VDD.n2374 GND 0.004404f
C3964 VDD.n2375 GND 0.004404f
C3965 VDD.n2376 GND 0.004404f
C3966 VDD.n2377 GND 0.004404f
C3967 VDD.n2378 GND 0.004404f
C3968 VDD.n2379 GND 0.004404f
C3969 VDD.n2380 GND 0.004404f
C3970 VDD.n2381 GND 0.004404f
C3971 VDD.n2382 GND 0.004404f
C3972 VDD.n2383 GND 0.004404f
C3973 VDD.n2384 GND 0.004404f
C3974 VDD.n2385 GND 0.004404f
C3975 VDD.n2386 GND 0.004404f
C3976 VDD.n2387 GND 0.004404f
C3977 VDD.n2388 GND 0.004404f
C3978 VDD.n2389 GND 0.004404f
C3979 VDD.n2390 GND 0.004404f
C3980 VDD.n2391 GND 0.004404f
C3981 VDD.n2392 GND 0.004404f
C3982 VDD.n2393 GND 0.004404f
C3983 VDD.n2394 GND 0.004404f
C3984 VDD.n2395 GND 0.004404f
C3985 VDD.n2396 GND 0.004404f
C3986 VDD.n2397 GND 0.004404f
C3987 VDD.n2398 GND 0.004404f
C3988 VDD.n2399 GND 0.004404f
C3989 VDD.n2400 GND 0.004404f
C3990 VDD.n2401 GND 0.004404f
C3991 VDD.n2402 GND 0.004404f
C3992 VDD.n2403 GND 0.004404f
C3993 VDD.n2404 GND 0.004404f
C3994 VDD.n2405 GND 0.004404f
C3995 VDD.n2406 GND 0.004404f
C3996 VDD.n2407 GND 0.004404f
C3997 VDD.n2408 GND 0.004404f
C3998 VDD.n2409 GND 0.004404f
C3999 VDD.n2410 GND 0.004404f
C4000 VDD.n2411 GND 0.004404f
C4001 VDD.n2412 GND 0.004404f
C4002 VDD.n2413 GND 0.004404f
C4003 VDD.n2414 GND 0.004404f
C4004 VDD.n2415 GND 0.004404f
C4005 VDD.n2416 GND 0.004404f
C4006 VDD.n2417 GND 0.004404f
C4007 VDD.n2418 GND 0.004404f
C4008 VDD.n2419 GND 0.004404f
C4009 VDD.n2420 GND 0.004404f
C4010 VDD.n2421 GND 0.004404f
C4011 VDD.n2422 GND 0.004404f
C4012 VDD.n2423 GND 0.004404f
C4013 VDD.n2424 GND 0.004404f
C4014 VDD.n2425 GND 0.004404f
C4015 VDD.n2426 GND 0.004404f
C4016 VDD.n2427 GND 0.004404f
C4017 VDD.n2428 GND 0.004404f
C4018 VDD.n2429 GND 0.004404f
C4019 VDD.n2430 GND 0.004404f
C4020 VDD.n2431 GND 0.004404f
C4021 VDD.n2432 GND 0.004404f
C4022 VDD.n2433 GND 0.004404f
C4023 VDD.n2434 GND 0.004404f
C4024 VDD.n2435 GND 0.004404f
C4025 VDD.n2436 GND 0.004404f
C4026 VDD.n2437 GND 0.004404f
C4027 VDD.n2438 GND 0.004404f
C4028 VDD.n2439 GND 0.004404f
C4029 VDD.n2440 GND 0.004404f
C4030 VDD.n2441 GND 0.004404f
C4031 VDD.n2442 GND 0.004404f
C4032 VDD.n2443 GND 0.004404f
C4033 VDD.n2444 GND 0.004404f
C4034 VDD.n2445 GND 0.004404f
C4035 VDD.n2446 GND 0.004404f
C4036 VDD.n2447 GND 0.004404f
C4037 VDD.n2448 GND 0.004404f
C4038 VDD.n2449 GND 0.004404f
C4039 VDD.n2450 GND 0.004404f
C4040 VDD.n2451 GND 0.004404f
C4041 VDD.n2452 GND 0.004404f
C4042 VDD.n2453 GND 0.004404f
C4043 VDD.n2454 GND 0.004404f
C4044 VDD.n2455 GND 0.004404f
C4045 VDD.n2456 GND 0.004404f
C4046 VDD.n2457 GND 0.004404f
C4047 VDD.n2458 GND 0.004404f
C4048 VDD.n2459 GND 0.004404f
C4049 VDD.n2460 GND 0.004404f
C4050 VDD.n2461 GND 0.004404f
C4051 VDD.n2462 GND 0.004404f
C4052 VDD.n2463 GND 0.004404f
C4053 VDD.n2464 GND 0.004404f
C4054 VDD.n2465 GND 0.004404f
C4055 VDD.n2466 GND 0.004404f
C4056 VDD.n2467 GND 0.004404f
C4057 VDD.n2468 GND 0.174018f
C4058 VDD.n2469 GND 0.004404f
C4059 VDD.n2470 GND 0.004404f
C4060 VDD.n2471 GND 0.004404f
C4061 VDD.n2472 GND 0.004404f
C4062 VDD.n2473 GND 0.004404f
C4063 VDD.n2474 GND 0.004404f
C4064 VDD.n2475 GND 0.004404f
C4065 VDD.n2476 GND 0.004404f
C4066 VDD.n2477 GND 0.004404f
C4067 VDD.n2478 GND 0.004404f
C4068 VDD.n2479 GND 0.004404f
C4069 VDD.n2480 GND 0.004404f
C4070 VDD.n2481 GND 0.010151f
C4071 VDD.n2482 GND 0.010151f
C4072 VDD.n2483 GND 0.01038f
C4073 VDD.n2484 GND 0.01038f
C4074 VDD.n2485 GND 0.004404f
C4075 VDD.n2486 GND 0.004404f
C4076 VDD.n2487 GND 0.004404f
C4077 VDD.n2488 GND 0.002753f
C4078 VDD.n2489 GND 0.006294f
C4079 VDD.n2490 GND 0.003854f
C4080 VDD.n2491 GND 0.004404f
C4081 VDD.n2492 GND 0.004404f
C4082 VDD.n2493 GND 0.004404f
C4083 VDD.n2494 GND 0.004404f
C4084 VDD.n2495 GND 0.004404f
C4085 VDD.n2496 GND 0.004404f
C4086 VDD.n2497 GND 0.004404f
C4087 VDD.n2498 GND 0.004404f
C4088 VDD.n2499 GND 0.004404f
C4089 VDD.n2500 GND 0.004404f
C4090 VDD.n2501 GND 0.004404f
C4091 VDD.n2502 GND 0.004404f
C4092 VDD.n2503 GND 0.004404f
C4093 VDD.n2504 GND 0.003303f
C4094 VDD.n2505 GND 0.032477f
C4095 VDD.n2506 GND 0.759602f
C4096 VDD.n2507 GND 0.008008f
C4097 VDD.n2508 GND 0.006477f
C4098 VDD.n2509 GND 0.006477f
C4099 VDD.n2510 GND 0.005213f
C4100 VDD.n2511 GND 0.006477f
C4101 VDD.n2512 GND 0.429674f
C4102 VDD.n2513 GND 0.429674f
C4103 VDD.n2514 GND 0.006477f
C4104 VDD.n2515 GND 0.005213f
C4105 VDD.n2516 GND 0.006477f
C4106 VDD.n2517 GND 0.006477f
C4107 VDD.n2518 GND 0.006477f
C4108 VDD.n2519 GND 0.005213f
C4109 VDD.n2520 GND 0.004327f
C4110 VDD.n2521 GND 0.014826f
C4111 VDD.n2522 GND 0.575763f
C4112 VDD.n2523 GND 0.014826f
C4113 VDD.n2524 GND 0.014967f
C4114 VDD.n2525 GND 0.002502f
C4115 VDD.n2526 GND 0.008028f
C4116 VDD.n2527 GND 0.002711f
C4117 VDD.n2528 GND 0.006477f
C4118 VDD.n2529 GND 0.006477f
C4119 VDD.n2530 GND 0.006477f
C4120 VDD.n2531 GND 0.005213f
C4121 VDD.n2532 GND 0.005213f
C4122 VDD.n2533 GND 0.005213f
C4123 VDD.n2534 GND 0.006477f
C4124 VDD.n2535 GND 0.006477f
C4125 VDD.n2536 GND 0.006477f
C4126 VDD.n2537 GND 0.005213f
C4127 VDD.n2538 GND 0.005213f
C4128 VDD.n2539 GND 0.005213f
C4129 VDD.n2540 GND 0.006477f
C4130 VDD.n2541 GND 0.006477f
C4131 VDD.n2542 GND 0.006477f
C4132 VDD.n2543 GND 0.005213f
C4133 VDD.n2544 GND 0.005213f
C4134 VDD.n2545 GND 0.005213f
C4135 VDD.n2546 GND 0.006477f
C4136 VDD.n2547 GND 0.006477f
C4137 VDD.n2548 GND 0.006477f
C4138 VDD.n2549 GND 0.004744f
C4139 VDD.n2550 GND 0.010634f
C4140 VDD.n2551 GND 0.003962f
C4141 VDD.n2552 GND 0.006477f
C4142 VDD.n2553 GND 0.006477f
C4143 VDD.n2554 GND 0.006477f
C4144 VDD.n2555 GND 0.005213f
C4145 VDD.n2556 GND 0.005213f
C4146 VDD.n2557 GND 0.005213f
C4147 VDD.n2558 GND 0.006477f
C4148 VDD.n2559 GND 0.006477f
C4149 VDD.n2560 GND 0.006477f
C4150 VDD.n2561 GND 0.005213f
C4151 VDD.n2562 GND 0.005213f
C4152 VDD.n2563 GND 0.005213f
C4153 VDD.n2564 GND 0.006477f
C4154 VDD.n2565 GND 0.006477f
C4155 VDD.n2566 GND 0.006477f
C4156 VDD.n2567 GND 0.005213f
C4157 VDD.n2568 GND 0.005213f
C4158 VDD.n2569 GND 0.004327f
C4159 VDD.n2570 GND 0.008031f
C4160 VDD.n2571 GND 0.659091f
C4161 VDD.n2572 GND 0.122139f
C4162 VDD.n2573 GND 0.003303f
C4163 VDD.n2574 GND 0.004404f
C4164 VDD.n2575 GND 0.004404f
C4165 VDD.n2576 GND 0.004404f
C4166 VDD.n2577 GND 0.004404f
C4167 VDD.n2578 GND 0.004404f
C4168 VDD.n2579 GND 0.004404f
C4169 VDD.n2580 GND 0.004404f
C4170 VDD.n2581 GND 0.004404f
C4171 VDD.n2582 GND 0.004404f
C4172 VDD.n2583 GND 0.004404f
C4173 VDD.n2584 GND 0.004404f
C4174 VDD.n2585 GND 0.004404f
C4175 VDD.n2586 GND 0.004404f
C4176 VDD.n2587 GND 0.004404f
C4177 VDD.n2588 GND 0.552131f
C4178 VDD.n2590 GND 0.01038f
C4179 VDD.n2591 GND 0.01038f
C4180 VDD.n2592 GND 0.010151f
C4181 VDD.n2593 GND 0.004404f
C4182 VDD.n2594 GND 0.004404f
C4183 VDD.n2595 GND 0.292178f
C4184 VDD.n2596 GND 0.004404f
C4185 VDD.n2597 GND 0.004404f
C4186 VDD.n2598 GND 0.004404f
C4187 VDD.n2599 GND 0.004404f
C4188 VDD.n2600 GND 0.004404f
C4189 VDD.n2601 GND 0.292178f
C4190 VDD.n2602 GND 0.004404f
C4191 VDD.n2603 GND 0.004404f
C4192 VDD.n2604 GND 0.004404f
C4193 VDD.n2605 GND 0.004404f
C4194 VDD.n2606 GND 0.004404f
C4195 VDD.n2607 GND 0.292178f
C4196 VDD.n2608 GND 0.004404f
C4197 VDD.n2609 GND 0.004404f
C4198 VDD.n2610 GND 0.004404f
C4199 VDD.n2611 GND 0.004404f
C4200 VDD.n2612 GND 0.004404f
C4201 VDD.n2613 GND 0.214837f
C4202 VDD.n2614 GND 0.004404f
C4203 VDD.n2615 GND 0.004404f
C4204 VDD.n2616 GND 0.004404f
C4205 VDD.n2617 GND 0.004404f
C4206 VDD.n2618 GND 0.004404f
C4207 VDD.n2619 GND 0.195502f
C4208 VDD.n2620 GND 0.004404f
C4209 VDD.n2621 GND 0.004404f
C4210 VDD.n2622 GND 0.004404f
C4211 VDD.n2623 GND 0.004404f
C4212 VDD.n2624 GND 0.004404f
C4213 VDD.n2625 GND 0.292178f
C4214 VDD.n2626 GND 0.004404f
C4215 VDD.n2627 GND 0.004404f
C4216 VDD.n2628 GND 0.004404f
C4217 VDD.n2629 GND 0.004404f
C4218 VDD.n2630 GND 0.004404f
C4219 VDD.n2631 GND 0.292178f
C4220 VDD.n2632 GND 0.004404f
C4221 VDD.n2633 GND 0.004404f
C4222 VDD.n2634 GND 0.004404f
C4223 VDD.n2635 GND 0.004404f
C4224 VDD.n2636 GND 0.004404f
C4225 VDD.n2637 GND 0.292178f
C4226 VDD.n2638 GND 0.004404f
C4227 VDD.n2639 GND 0.004404f
C4228 VDD.n2640 GND 0.004404f
C4229 VDD.n2641 GND 0.004404f
C4230 VDD.n2642 GND 0.004404f
C4231 VDD.n2643 GND 0.292178f
C4232 VDD.n2644 GND 0.004404f
C4233 VDD.n2645 GND 0.004404f
C4234 VDD.n2646 GND 0.004404f
C4235 VDD.n2647 GND 0.004404f
C4236 VDD.n2648 GND 0.004404f
C4237 VDD.n2649 GND 0.292178f
C4238 VDD.n2650 GND 0.004404f
C4239 VDD.n2651 GND 0.004404f
C4240 VDD.n2652 GND 0.004404f
C4241 VDD.n2653 GND 0.004404f
C4242 VDD.n2654 GND 0.004404f
C4243 VDD.n2655 GND 0.161128f
C4244 VDD.n2656 GND 0.004404f
C4245 VDD.n2657 GND 0.004404f
C4246 VDD.n2658 GND 0.004404f
C4247 VDD.n2659 GND 0.004404f
C4248 VDD.n2660 GND 0.004404f
C4249 VDD.n2661 GND 0.163276f
C4250 VDD.n2662 GND 0.004404f
C4251 VDD.n2663 GND 0.004404f
C4252 VDD.n2664 GND 0.004404f
C4253 VDD.n2665 GND 0.004404f
C4254 VDD.n2666 GND 0.004404f
C4255 VDD.n2667 GND 0.292178f
C4256 VDD.n2668 GND 0.004404f
C4257 VDD.n2669 GND 0.004404f
C4258 VDD.n2670 GND 0.004404f
C4259 VDD.n2671 GND 0.004404f
C4260 VDD.n2672 GND 0.004404f
C4261 VDD.n2673 GND 0.292178f
C4262 VDD.n2674 GND 0.004404f
C4263 VDD.n2675 GND 0.004404f
C4264 VDD.n2676 GND 0.004404f
C4265 VDD.n2677 GND 0.004404f
C4266 VDD.n2678 GND 0.004404f
C4267 VDD.n2679 GND 0.292178f
C4268 VDD.n2680 GND 0.004404f
C4269 VDD.n2681 GND 0.004404f
C4270 VDD.n2682 GND 0.004404f
C4271 VDD.n2683 GND 0.004404f
C4272 VDD.n2684 GND 0.004404f
C4273 VDD.n2685 GND 0.292178f
C4274 VDD.n2686 GND 0.004404f
C4275 VDD.n2687 GND 0.004404f
C4276 VDD.n2688 GND 0.004404f
C4277 VDD.n2689 GND 0.004404f
C4278 VDD.n2690 GND 0.004404f
C4279 VDD.n2691 GND 0.225579f
C4280 VDD.n2692 GND 0.004404f
C4281 VDD.n2693 GND 0.004404f
C4282 VDD.n2694 GND 0.004404f
C4283 VDD.n2695 GND 0.004404f
C4284 VDD.n2696 GND 0.004404f
C4285 VDD.n2697 GND 0.227727f
C4286 VDD.n2698 GND 0.004404f
C4287 VDD.n2699 GND 0.004404f
C4288 VDD.n2700 GND 0.004404f
C4289 VDD.n2701 GND 0.004404f
C4290 VDD.n2702 GND 0.004404f
C4291 VDD.n2703 GND 0.292178f
C4292 VDD.n2704 GND 0.004404f
C4293 VDD.n2705 GND 0.004404f
C4294 VDD.n2706 GND 0.004404f
C4295 VDD.n2707 GND 0.004404f
C4296 VDD.n2708 GND 0.004404f
C4297 VDD.n2709 GND 0.292178f
C4298 VDD.n2710 GND 0.004404f
C4299 VDD.n2711 GND 0.004404f
C4300 VDD.n2712 GND 0.004404f
C4301 VDD.n2713 GND 0.004404f
C4302 VDD.n2714 GND 0.004404f
C4303 VDD.n2715 GND 0.292178f
C4304 VDD.n2716 GND 0.004404f
C4305 VDD.n2717 GND 0.004404f
C4306 VDD.n2718 GND 0.004404f
C4307 VDD.n2719 GND 0.004404f
C4308 VDD.n2720 GND 0.004404f
C4309 VDD.n2721 GND 0.292178f
C4310 VDD.n2722 GND 0.004404f
C4311 VDD.n2723 GND 0.004404f
C4312 VDD.n2724 GND 0.004404f
C4313 VDD.n2725 GND 0.004404f
C4314 VDD.n2726 GND 0.004404f
C4315 VDD.n2727 GND 0.292178f
C4316 VDD.n2728 GND 0.004404f
C4317 VDD.n2729 GND 0.004404f
C4318 VDD.n2730 GND 0.004404f
C4319 VDD.n2731 GND 0.004404f
C4320 VDD.n2732 GND 0.004404f
C4321 VDD.n2733 GND 0.292178f
C4322 VDD.n2734 GND 0.004404f
C4323 VDD.n2735 GND 0.004404f
C4324 VDD.n2736 GND 0.004404f
C4325 VDD.n2737 GND 0.004404f
C4326 VDD.n2738 GND 0.004404f
C4327 VDD.n2739 GND 0.292178f
C4328 VDD.n2740 GND 0.004404f
C4329 VDD.n2741 GND 0.004404f
C4330 VDD.n2742 GND 0.004404f
C4331 VDD.n2743 GND 0.004404f
C4332 VDD.n2744 GND 0.004404f
C4333 VDD.n2745 GND 0.292178f
C4334 VDD.n2746 GND 0.004404f
C4335 VDD.n2747 GND 0.004404f
C4336 VDD.n2748 GND 0.004404f
C4337 VDD.n2749 GND 0.004404f
C4338 VDD.n2750 GND 0.004404f
C4339 VDD.n2751 GND 0.242766f
C4340 VDD.n2752 GND 0.004404f
C4341 VDD.n2753 GND 0.004404f
C4342 VDD.n2754 GND 0.004404f
C4343 VDD.n2755 GND 0.004404f
C4344 VDD.n2756 GND 0.004404f
C4345 VDD.n2757 GND 0.292178f
C4346 VDD.n2758 GND 0.004404f
C4347 VDD.n2759 GND 0.004404f
C4348 VDD.n2760 GND 0.004404f
C4349 VDD.n2761 GND 0.004404f
C4350 VDD.n2762 GND 0.004404f
C4351 VDD.n2763 GND 0.292178f
C4352 VDD.n2764 GND 0.004404f
C4353 VDD.n2765 GND 0.004404f
C4354 VDD.n2766 GND 0.004404f
C4355 VDD.n2767 GND 0.004404f
C4356 VDD.n2768 GND 0.004404f
C4357 VDD.n2769 GND 0.292178f
C4358 VDD.n2770 GND 0.004404f
C4359 VDD.n2771 GND 0.004404f
C4360 VDD.n2772 GND 0.004404f
C4361 VDD.n2773 GND 0.004404f
C4362 VDD.n2774 GND 0.004404f
C4363 VDD.n2775 GND 0.227727f
C4364 VDD.n2776 GND 0.004404f
C4365 VDD.n2777 GND 0.004404f
C4366 VDD.n2778 GND 0.004404f
C4367 VDD.n2779 GND 0.004404f
C4368 VDD.n2780 GND 0.004404f
C4369 VDD.n2781 GND 0.292178f
C4370 VDD.n2782 GND 0.004404f
C4371 VDD.n2783 GND 0.004404f
C4372 VDD.n2784 GND 0.004404f
C4373 VDD.n2785 GND 0.004404f
C4374 VDD.n2786 GND 0.004404f
C4375 VDD.n2787 GND 0.178315f
C4376 VDD.n2788 GND 0.004404f
C4377 VDD.n2789 GND 0.004404f
C4378 VDD.n2790 GND 0.004404f
C4379 VDD.n2791 GND 0.004404f
C4380 VDD.n2792 GND 0.004404f
C4381 VDD.n2793 GND 0.292178f
C4382 VDD.n2794 GND 0.004404f
C4383 VDD.n2795 GND 0.004404f
C4384 VDD.n2796 GND 0.004404f
C4385 VDD.n2797 GND 0.004404f
C4386 VDD.n2798 GND 0.004404f
C4387 VDD.n2799 GND 0.292178f
C4388 VDD.n2800 GND 0.004404f
C4389 VDD.n2801 GND 0.004404f
C4390 VDD.n2802 GND 0.004404f
C4391 VDD.n2803 GND 0.004404f
C4392 VDD.n2804 GND 0.004404f
C4393 VDD.n2805 GND 0.292178f
C4394 VDD.n2806 GND 0.004404f
C4395 VDD.n2807 GND 0.004404f
C4396 VDD.n2808 GND 0.004404f
C4397 VDD.n2809 GND 0.004404f
C4398 VDD.n2810 GND 0.004404f
C4399 VDD.n2811 GND 0.163276f
C4400 VDD.n2812 GND 0.004404f
C4401 VDD.n2813 GND 0.004404f
C4402 VDD.n2814 GND 0.004404f
C4403 VDD.n2815 GND 0.004404f
C4404 VDD.n2816 GND 0.004404f
C4405 VDD.n2817 GND 0.292178f
C4406 VDD.n2818 GND 0.004404f
C4407 VDD.n2819 GND 0.004404f
C4408 VDD.n2820 GND 0.004404f
C4409 VDD.n2821 GND 0.004404f
C4410 VDD.n2822 GND 0.004404f
C4411 VDD.n2823 GND 0.178315f
C4412 VDD.n2824 GND 0.004404f
C4413 VDD.n2825 GND 0.004404f
C4414 VDD.n2826 GND 0.004404f
C4415 VDD.n2827 GND 0.004404f
C4416 VDD.n2828 GND 0.004404f
C4417 VDD.n2829 GND 0.292178f
C4418 VDD.n2830 GND 0.004404f
C4419 VDD.n2831 GND 0.004404f
C4420 VDD.n2832 GND 0.004404f
C4421 VDD.n2833 GND 0.004404f
C4422 VDD.n2834 GND 0.004404f
C4423 VDD.n2835 GND 0.292178f
C4424 VDD.n2836 GND 0.004404f
C4425 VDD.n2837 GND 0.004404f
C4426 VDD.n2838 GND 0.004404f
C4427 VDD.n2839 GND 0.004404f
C4428 VDD.n2840 GND 0.004404f
C4429 VDD.n2841 GND 0.292178f
C4430 VDD.n2842 GND 0.004404f
C4431 VDD.n2843 GND 0.004404f
C4432 VDD.n2844 GND 0.004404f
C4433 VDD.n2845 GND 0.004404f
C4434 VDD.n2846 GND 0.004404f
C4435 VDD.n2847 GND 0.292178f
C4436 VDD.n2848 GND 0.004404f
C4437 VDD.n2849 GND 0.004404f
C4438 VDD.n2850 GND 0.004404f
C4439 VDD.n2851 GND 0.004404f
C4440 VDD.n2852 GND 0.004404f
C4441 VDD.n2853 GND 0.292178f
C4442 VDD.n2854 GND 0.004404f
C4443 VDD.n2855 GND 0.004404f
C4444 VDD.n2856 GND 0.004404f
C4445 VDD.n2857 GND 0.004404f
C4446 VDD.n2858 GND 0.004404f
C4447 VDD.n2859 GND 0.165425f
C4448 VDD.n2860 GND 0.004404f
C4449 VDD.n2861 GND 0.004404f
C4450 VDD.n2862 GND 0.004404f
C4451 VDD.t76 GND 0.068381f
C4452 VDD.t75 GND 0.084764f
C4453 VDD.t73 GND 0.489916f
C4454 VDD.n2863 GND 0.064611f
C4455 VDD.n2864 GND 0.042608f
C4456 VDD.n2865 GND 0.004404f
C4457 VDD.n2866 GND 0.002753f
C4458 VDD.n2867 GND 0.006294f
C4459 VDD.n2868 GND 0.003854f
C4460 VDD.n2869 GND 0.004404f
C4461 VDD.n2870 GND 0.004404f
C4462 VDD.n2871 GND 0.004404f
C4463 VDD.n2872 GND 0.004404f
C4464 VDD.n2873 GND 0.004404f
C4465 VDD.n2874 GND 0.004404f
C4466 VDD.n2875 GND 0.004404f
C4467 VDD.n2876 GND 0.004404f
C4468 VDD.n2877 GND 0.004404f
C4469 VDD.n2878 GND 0.004404f
C4470 VDD.n2879 GND 0.004404f
C4471 VDD.n2880 GND 0.004404f
C4472 VDD.n2881 GND 0.004404f
C4473 VDD.n2882 GND 0.004404f
C4474 VDD.n2883 GND 0.004404f
C4475 VDD.n2884 GND 0.004404f
C4476 VDD.n2885 GND 0.004404f
C4477 VDD.n2886 GND 0.004404f
C4478 VDD.n2887 GND 0.004404f
C4479 VDD.n2888 GND 0.004404f
C4480 VDD.n2889 GND 0.004404f
C4481 VDD.n2890 GND 0.004404f
C4482 VDD.n2891 GND 0.004404f
C4483 VDD.n2892 GND 0.004404f
C4484 VDD.n2893 GND 0.004404f
C4485 VDD.n2894 GND 0.004404f
C4486 VDD.n2895 GND 0.004404f
C4487 VDD.n2896 GND 0.004404f
C4488 VDD.n2897 GND 0.004404f
C4489 VDD.n2898 GND 0.004404f
C4490 VDD.n2899 GND 0.004404f
C4491 VDD.n2900 GND 0.01038f
C4492 VDD.n2901 GND 0.01038f
C4493 VDD.n2902 GND 0.010151f
C4494 VDD.n2903 GND 0.010151f
C4495 VDD.n2904 GND 0.004404f
C4496 VDD.n2905 GND 0.004404f
C4497 VDD.n2906 GND 0.004404f
C4498 VDD.n2907 GND 0.004404f
C4499 VDD.n2908 GND 0.004404f
C4500 VDD.n2909 GND 0.004404f
C4501 VDD.n2910 GND 0.004404f
C4502 VDD.n2911 GND 0.292178f
C4503 VDD.n2912 GND 0.004404f
C4504 VDD.n2913 GND 0.004404f
C4505 VDD.n2914 GND 0.004404f
C4506 VDD.n2915 GND 0.004404f
C4507 VDD.n2916 GND 0.004404f
C4508 VDD.n2917 GND 0.292178f
C4509 VDD.n2918 GND 0.004404f
C4510 VDD.n2919 GND 0.004404f
C4511 VDD.n2920 GND 0.004404f
C4512 VDD.n2921 GND 0.004404f
C4513 VDD.n2922 GND 0.010674f
C4514 VDD.n2923 GND 0.010151f
C4515 VDD.n2924 GND 0.01038f
C4516 VDD.n2925 GND 0.009857f
C4517 VDD.n2926 GND 0.004404f
C4518 VDD.n2927 GND 0.004404f
C4519 VDD.n2928 GND 0.004404f
C4520 VDD.n2929 GND 0.002753f
C4521 VDD.n2930 GND 0.006294f
C4522 VDD.n2931 GND 0.003854f
C4523 VDD.n2932 GND 0.004404f
C4524 VDD.n2933 GND 0.004404f
C4525 VDD.n2934 GND 0.004404f
C4526 VDD.n2935 GND 0.004404f
C4527 VDD.n2936 GND 0.004404f
C4528 VDD.n2937 GND 0.004404f
C4529 VDD.n2938 GND 0.004404f
C4530 VDD.n2939 GND 0.004404f
C4531 VDD.n2940 GND 0.004404f
C4532 VDD.n2941 GND 0.004404f
C4533 VDD.n2942 GND 0.004404f
C4534 VDD.n2943 GND 0.004404f
C4535 VDD.n2944 GND 0.004404f
C4536 VDD.n2945 GND 0.004404f
C4537 VDD.n2946 GND 0.004404f
C4538 VDD.n2947 GND 0.004404f
C4539 VDD.n2948 GND 0.004404f
C4540 VDD.n2949 GND 0.004404f
C4541 VDD.n2950 GND 0.004404f
C4542 VDD.n2951 GND 0.004404f
C4543 VDD.n2952 GND 0.004404f
C4544 VDD.n2953 GND 0.004404f
C4545 VDD.n2954 GND 0.004404f
C4546 VDD.n2955 GND 0.004404f
C4547 VDD.n2956 GND 0.004404f
C4548 VDD.n2957 GND 0.004404f
C4549 VDD.n2958 GND 0.004404f
C4550 VDD.n2959 GND 0.004404f
C4551 VDD.n2960 GND 0.004404f
C4552 VDD.n2961 GND 0.004404f
C4553 VDD.n2962 GND 0.004404f
C4554 VDD.n2963 GND 0.01038f
C4555 VDD.n2964 GND 0.01038f
C4556 VDD.n2965 GND 0.010151f
C4557 VDD.n2966 GND 0.004404f
C4558 VDD.n2967 GND 0.004404f
C4559 VDD.n2968 GND 0.292178f
C4560 VDD.n2969 GND 0.004404f
C4561 VDD.n2970 GND 0.004404f
C4562 VDD.n2971 GND 0.010674f
C4563 VDD.n2972 GND 0.009857f
C4564 VDD.n2973 GND 0.01038f
C4565 VDD.n2975 GND 1.80248f
C4566 VDD.n2976 GND 1.80248f
C4567 VDD.n2977 GND 0.010151f
C4568 VDD.n2978 GND 0.010151f
C4569 VDD.n2979 GND 0.01038f
C4570 VDD.n2980 GND 0.004404f
C4571 VDD.n2981 GND 0.004404f
C4572 VDD.n2982 GND 0.004404f
C4573 VDD.n2983 GND 0.004404f
C4574 VDD.n2984 GND 0.004404f
C4575 VDD.n2985 GND 0.004404f
C4576 VDD.n2986 GND 0.004404f
C4577 VDD.n2987 GND 0.004404f
C4578 VDD.t91 GND 0.068381f
C4579 VDD.t92 GND 0.084764f
C4580 VDD.t89 GND 0.489916f
C4581 VDD.n2988 GND 0.064611f
C4582 VDD.n2989 GND 0.042608f
C4583 VDD.n2990 GND 0.004404f
C4584 VDD.n2991 GND 0.004404f
C4585 VDD.n2992 GND 0.004404f
C4586 VDD.n2993 GND 0.004404f
C4587 VDD.n2994 GND 0.004404f
C4588 VDD.n2995 GND 0.004404f
C4589 VDD.n2996 GND 0.004404f
C4590 VDD.n2997 GND 0.004404f
C4591 VDD.n2998 GND 0.004404f
C4592 VDD.n2999 GND 0.004404f
C4593 VDD.n3000 GND 0.004404f
C4594 VDD.n3001 GND 0.004404f
C4595 VDD.n3002 GND 0.004404f
C4596 VDD.n3003 GND 0.004404f
C4597 VDD.n3004 GND 0.004404f
C4598 VDD.n3005 GND 0.004404f
C4599 VDD.n3006 GND 0.004404f
C4600 VDD.n3007 GND 0.004404f
C4601 VDD.n3008 GND 0.004404f
C4602 VDD.n3009 GND 0.004404f
C4603 VDD.n3010 GND 0.004404f
C4604 VDD.n3011 GND 0.004404f
C4605 VDD.n3012 GND 0.004404f
C4606 VDD.n3013 GND 0.004404f
C4607 VDD.n3014 GND 0.004404f
C4608 VDD.n3015 GND 0.004404f
C4609 VDD.n3016 GND 0.004404f
C4610 VDD.n3017 GND 0.004404f
C4611 VDD.n3018 GND 0.004404f
C4612 VDD.n3019 GND 0.004404f
C4613 VDD.n3020 GND 0.004404f
C4614 VDD.n3021 GND 0.004404f
C4615 VDD.n3022 GND 0.004404f
C4616 VDD.n3023 GND 0.004404f
C4617 VDD.n3024 GND 0.004404f
C4618 VDD.n3025 GND 0.004404f
C4619 VDD.n3026 GND 0.004404f
C4620 VDD.n3027 GND 0.004404f
C4621 VDD.n3028 GND 0.004404f
C4622 VDD.n3029 GND 0.004404f
C4623 VDD.n3030 GND 0.004404f
C4624 VDD.n3031 GND 0.004404f
C4625 VDD.n3032 GND 0.004404f
C4626 VDD.n3033 GND 0.004404f
C4627 VDD.n3034 GND 0.004404f
C4628 VDD.n3035 GND 0.004404f
C4629 VDD.n3036 GND 0.004404f
C4630 VDD.n3037 GND 0.004404f
C4631 VDD.n3038 GND 0.004404f
C4632 VDD.n3039 GND 0.004404f
C4633 VDD.n3040 GND 0.004404f
C4634 VDD.n3041 GND 0.004404f
C4635 VDD.n3042 GND 0.004404f
C4636 VDD.n3043 GND 0.004404f
C4637 VDD.n3044 GND 0.004404f
C4638 VDD.n3045 GND 0.004404f
C4639 VDD.n3046 GND 0.004404f
C4640 VDD.n3047 GND 0.004404f
C4641 VDD.n3048 GND 0.004404f
C4642 VDD.n3049 GND 0.004404f
C4643 VDD.n3050 GND 0.004404f
C4644 VDD.n3051 GND 0.004404f
C4645 VDD.n3052 GND 0.004404f
C4646 VDD.n3053 GND 0.004404f
C4647 VDD.n3054 GND 0.004404f
C4648 VDD.n3055 GND 0.004404f
C4649 VDD.n3056 GND 0.004404f
C4650 VDD.n3057 GND 0.004404f
C4651 VDD.n3058 GND 0.004404f
C4652 VDD.n3059 GND 0.004404f
C4653 VDD.n3060 GND 0.004404f
C4654 VDD.n3061 GND 0.004404f
C4655 VDD.n3062 GND 0.004404f
C4656 VDD.n3063 GND 0.004404f
C4657 VDD.n3064 GND 0.004404f
C4658 VDD.n3065 GND 0.004404f
C4659 VDD.n3066 GND 0.004404f
C4660 VDD.n3067 GND 0.004404f
C4661 VDD.n3068 GND 0.004404f
C4662 VDD.n3069 GND 0.004404f
C4663 VDD.n3070 GND 0.004404f
C4664 VDD.n3071 GND 0.004404f
C4665 VDD.n3072 GND 0.004404f
C4666 VDD.n3073 GND 0.004404f
C4667 VDD.n3074 GND 0.004404f
C4668 VDD.n3075 GND 0.004404f
C4669 VDD.n3076 GND 0.004404f
C4670 VDD.n3077 GND 0.004404f
C4671 VDD.n3078 GND 0.004404f
C4672 VDD.n3079 GND 0.004404f
C4673 VDD.n3080 GND 0.004404f
C4674 VDD.n3081 GND 0.004404f
C4675 VDD.n3082 GND 0.004404f
C4676 VDD.n3083 GND 0.004404f
C4677 VDD.n3084 GND 0.004404f
C4678 VDD.n3085 GND 0.004404f
C4679 VDD.n3086 GND 0.004404f
C4680 VDD.n3087 GND 0.004404f
C4681 VDD.n3088 GND 0.004404f
C4682 VDD.n3089 GND 0.004404f
C4683 VDD.n3090 GND 0.004404f
C4684 VDD.n3091 GND 0.004404f
C4685 VDD.n3092 GND 0.004404f
C4686 VDD.n3093 GND 0.004404f
C4687 VDD.n3094 GND 0.004404f
C4688 VDD.n3095 GND 0.004404f
C4689 VDD.n3096 GND 0.004404f
C4690 VDD.n3097 GND 0.004404f
C4691 VDD.n3098 GND 0.004404f
C4692 VDD.n3099 GND 0.004404f
C4693 VDD.n3100 GND 0.004404f
C4694 VDD.n3101 GND 0.004404f
C4695 VDD.n3102 GND 0.004404f
C4696 VDD.n3103 GND 0.004404f
C4697 VDD.n3104 GND 0.004404f
C4698 VDD.n3105 GND 0.004404f
C4699 VDD.n3106 GND 0.004404f
C4700 VDD.n3107 GND 0.004404f
C4701 VDD.n3108 GND 0.004404f
C4702 VDD.n3109 GND 0.004404f
C4703 VDD.n3110 GND 0.004404f
C4704 VDD.n3111 GND 0.004404f
C4705 VDD.n3112 GND 0.004404f
C4706 VDD.n3113 GND 0.004404f
C4707 VDD.n3114 GND 0.004404f
C4708 VDD.n3115 GND 0.004404f
C4709 VDD.n3116 GND 0.004404f
C4710 VDD.n3117 GND 0.004404f
C4711 VDD.n3118 GND 0.004404f
C4712 VDD.n3119 GND 0.004404f
C4713 VDD.n3120 GND 0.004404f
C4714 VDD.n3121 GND 0.004404f
C4715 VDD.n3122 GND 0.004404f
C4716 VDD.n3123 GND 0.004404f
C4717 VDD.t111 GND 0.068381f
C4718 VDD.t112 GND 0.084764f
C4719 VDD.t110 GND 0.489916f
C4720 VDD.n3124 GND 0.064611f
C4721 VDD.n3125 GND 0.042608f
C4722 VDD.n3126 GND 0.004404f
C4723 VDD.n3127 GND 0.004404f
C4724 VDD.n3128 GND 0.004404f
C4725 VDD.n3129 GND 0.004404f
C4726 VDD.n3130 GND 0.004404f
C4727 VDD.n3131 GND 0.004404f
C4728 VDD.n3132 GND 0.004404f
C4729 VDD.n3133 GND 0.004404f
C4730 VDD.n3135 GND 0.004404f
C4731 VDD.n3136 GND 0.004404f
C4732 VDD.n3138 GND 0.004404f
C4733 VDD.n3139 GND 0.004404f
C4734 VDD.n3140 GND 0.004404f
C4735 VDD.n3141 GND 0.004404f
C4736 VDD.n3142 GND 0.004404f
C4737 VDD.n3144 GND 0.004404f
C4738 VDD.n3146 GND 0.004404f
C4739 VDD.n3147 GND 0.004404f
C4740 VDD.n3148 GND 0.004404f
C4741 VDD.n3149 GND 0.004404f
C4742 VDD.n3150 GND 0.004404f
C4743 VDD.n3152 GND 0.004404f
C4744 VDD.n3154 GND 0.004404f
C4745 VDD.n3155 GND 0.004404f
C4746 VDD.n3156 GND 0.004404f
C4747 VDD.n3157 GND 0.004404f
C4748 VDD.n3158 GND 0.004404f
C4749 VDD.n3160 GND 0.004404f
C4750 VDD.n3162 GND 0.004404f
C4751 VDD.n3163 GND 0.004404f
C4752 VDD.n3164 GND 0.003854f
C4753 VDD.n3165 GND 0.006294f
C4754 VDD.n3166 GND 0.002753f
C4755 VDD.n3167 GND 0.004404f
C4756 VDD.n3169 GND 0.004404f
C4757 VDD.n3170 GND 0.01038f
C4758 VDD.n3171 GND 0.01038f
C4759 VDD.n3172 GND 0.010151f
C4760 VDD.n3173 GND 0.004404f
C4761 VDD.n3174 GND 0.004404f
C4762 VDD.n3175 GND 0.004404f
C4763 VDD.n3176 GND 0.004404f
C4764 VDD.n3177 GND 0.004404f
C4765 VDD.n3178 GND 0.004404f
C4766 VDD.n3179 GND 0.004404f
C4767 VDD.n3180 GND 0.004404f
C4768 VDD.n3181 GND 0.004404f
C4769 VDD.n3182 GND 0.004404f
C4770 VDD.n3183 GND 0.004404f
C4771 VDD.n3184 GND 0.004404f
C4772 VDD.n3185 GND 0.004404f
C4773 VDD.n3186 GND 0.004404f
C4774 VDD.n3187 GND 0.004404f
C4775 VDD.n3188 GND 0.004404f
C4776 VDD.n3189 GND 0.004404f
C4777 VDD.n3190 GND 0.004404f
C4778 VDD.n3191 GND 0.004404f
C4779 VDD.n3192 GND 0.004404f
C4780 VDD.n3193 GND 0.004404f
C4781 VDD.n3194 GND 0.004404f
C4782 VDD.n3195 GND 0.004404f
C4783 VDD.n3196 GND 0.004404f
C4784 VDD.n3197 GND 0.004404f
C4785 VDD.n3198 GND 0.004404f
C4786 VDD.n3199 GND 0.004404f
C4787 VDD.n3200 GND 0.004404f
C4788 VDD.n3201 GND 0.004404f
C4789 VDD.n3202 GND 0.004404f
C4790 VDD.n3203 GND 0.004404f
C4791 VDD.n3204 GND 0.004404f
C4792 VDD.n3205 GND 0.004404f
C4793 VDD.n3206 GND 0.004404f
C4794 VDD.n3207 GND 0.004404f
C4795 VDD.n3208 GND 0.004404f
C4796 VDD.n3209 GND 0.004404f
C4797 VDD.n3210 GND 0.004404f
C4798 VDD.n3211 GND 0.004404f
C4799 VDD.n3212 GND 0.004404f
C4800 VDD.n3213 GND 0.004404f
C4801 VDD.n3214 GND 0.004404f
C4802 VDD.n3215 GND 0.004404f
C4803 VDD.n3216 GND 0.004404f
C4804 VDD.n3217 GND 0.004404f
C4805 VDD.n3218 GND 0.004404f
C4806 VDD.n3219 GND 0.004404f
C4807 VDD.n3220 GND 0.004404f
C4808 VDD.n3221 GND 0.004404f
C4809 VDD.n3222 GND 0.004404f
C4810 VDD.n3223 GND 0.004404f
C4811 VDD.n3224 GND 0.004404f
C4812 VDD.n3225 GND 0.004404f
C4813 VDD.n3226 GND 0.004404f
C4814 VDD.n3227 GND 0.004404f
C4815 VDD.n3228 GND 0.004404f
C4816 VDD.n3229 GND 0.004404f
C4817 VDD.n3230 GND 0.004404f
C4818 VDD.n3231 GND 0.004404f
C4819 VDD.n3232 GND 0.004404f
C4820 VDD.n3233 GND 0.004404f
C4821 VDD.n3234 GND 0.004404f
C4822 VDD.n3235 GND 0.004404f
C4823 VDD.n3236 GND 0.004404f
C4824 VDD.n3237 GND 0.004404f
C4825 VDD.n3238 GND 0.004404f
C4826 VDD.n3239 GND 0.165425f
C4827 VDD.n3240 GND 0.004404f
C4828 VDD.n3241 GND 0.004404f
C4829 VDD.n3242 GND 0.004404f
C4830 VDD.n3243 GND 0.004404f
C4831 VDD.n3244 GND 0.004404f
C4832 VDD.n3245 GND 0.004404f
C4833 VDD.n3246 GND 0.004404f
C4834 VDD.n3247 GND 0.004404f
C4835 VDD.n3248 GND 0.004404f
C4836 VDD.n3249 GND 0.004404f
C4837 VDD.n3250 GND 0.004404f
C4838 VDD.n3251 GND 0.010151f
C4839 VDD.n3252 GND 0.01038f
C4840 VDD.n3253 GND 0.01038f
C4841 VDD.n3255 GND 0.004404f
C4842 VDD.n3257 GND 0.004404f
C4843 VDD.n3258 GND 0.002753f
C4844 VDD.n3259 GND 0.006294f
C4845 VDD.n3260 GND 0.003854f
C4846 VDD.n3261 GND 0.004404f
C4847 VDD.n3262 GND 0.004404f
C4848 VDD.n3264 GND 0.004404f
C4849 VDD.n3266 GND 0.004404f
C4850 VDD.n3267 GND 0.004404f
C4851 VDD.n3268 GND 0.004404f
C4852 VDD.n3269 GND 0.004404f
C4853 VDD.n3270 GND 0.004404f
C4854 VDD.n3272 GND 0.004404f
C4855 VDD.n3274 GND 0.004404f
C4856 VDD.n3275 GND 0.004404f
C4857 VDD.n3276 GND 0.004404f
C4858 VDD.n3277 GND 0.004404f
C4859 VDD.n3278 GND 0.004404f
C4860 VDD.n3280 GND 0.004404f
C4861 VDD.n3282 GND 0.004404f
C4862 VDD.n3283 GND 0.004404f
C4863 VDD.n3284 GND 0.004404f
C4864 VDD.n3285 GND 0.004404f
C4865 VDD.n3286 GND 0.004404f
C4866 VDD.n3288 GND 0.004404f
C4867 VDD.n3290 GND 0.004404f
C4868 VDD.n3291 GND 0.004404f
C4869 VDD.n3292 GND 0.01038f
C4870 VDD.n3293 GND 0.010151f
C4871 VDD.n3294 GND 0.010151f
C4872 VDD.n3295 GND 0.388855f
C4873 VDD.n3296 GND 0.010151f
C4874 VDD.n3297 GND 0.010151f
C4875 VDD.n3298 GND 0.004404f
C4876 VDD.n3299 GND 0.004404f
C4877 VDD.n3300 GND 0.004404f
C4878 VDD.n3301 GND 0.292178f
C4879 VDD.n3302 GND 0.004404f
C4880 VDD.n3303 GND 0.004404f
C4881 VDD.n3304 GND 0.004404f
C4882 VDD.n3305 GND 0.004404f
C4883 VDD.n3306 GND 0.004404f
C4884 VDD.n3307 GND 0.292178f
C4885 VDD.n3308 GND 0.004404f
C4886 VDD.n3309 GND 0.004404f
C4887 VDD.n3310 GND 0.004404f
C4888 VDD.n3311 GND 0.004404f
C4889 VDD.n3312 GND 0.004404f
C4890 VDD.n3313 GND 0.195502f
C4891 VDD.n3314 GND 0.004404f
C4892 VDD.n3315 GND 0.004404f
C4893 VDD.n3316 GND 0.004404f
C4894 VDD.n3317 GND 0.004404f
C4895 VDD.n3318 GND 0.004404f
C4896 VDD.n3319 GND 0.223431f
C4897 VDD.n3320 GND 0.004404f
C4898 VDD.n3321 GND 0.004404f
C4899 VDD.n3322 GND 0.004404f
C4900 VDD.n3323 GND 0.004404f
C4901 VDD.n3324 GND 0.004404f
C4902 VDD.n3325 GND 0.292178f
C4903 VDD.n3326 GND 0.004404f
C4904 VDD.n3327 GND 0.004404f
C4905 VDD.n3328 GND 0.004404f
C4906 VDD.n3329 GND 0.004404f
C4907 VDD.n3330 GND 0.004404f
C4908 VDD.n3331 GND 0.292178f
C4909 VDD.n3332 GND 0.004404f
C4910 VDD.n3333 GND 0.004404f
C4911 VDD.n3334 GND 0.004404f
C4912 VDD.n3335 GND 0.004404f
C4913 VDD.n3336 GND 0.004404f
C4914 VDD.n3337 GND 0.292178f
C4915 VDD.n3338 GND 0.004404f
C4916 VDD.n3339 GND 0.004404f
C4917 VDD.n3340 GND 0.004404f
C4918 VDD.n3341 GND 0.004404f
C4919 VDD.n3342 GND 0.004404f
C4920 VDD.n3343 GND 0.292178f
C4921 VDD.n3344 GND 0.004404f
C4922 VDD.n3345 GND 0.004404f
C4923 VDD.n3346 GND 0.004404f
C4924 VDD.n3347 GND 0.004404f
C4925 VDD.n3348 GND 0.004404f
C4926 VDD.n3349 GND 0.259953f
C4927 VDD.n3350 GND 0.004404f
C4928 VDD.n3351 GND 0.004404f
C4929 VDD.n3352 GND 0.004404f
C4930 VDD.n3353 GND 0.004404f
C4931 VDD.n3354 GND 0.004404f
C4932 VDD.n3355 GND 0.292178f
C4933 VDD.n3356 GND 0.004404f
C4934 VDD.n3357 GND 0.004404f
C4935 VDD.n3358 GND 0.004404f
C4936 VDD.n3359 GND 0.004404f
C4937 VDD.n3360 GND 0.004404f
C4938 VDD.n3361 GND 0.292178f
C4939 VDD.n3362 GND 0.004404f
C4940 VDD.n3363 GND 0.004404f
C4941 VDD.n3364 GND 0.004404f
C4942 VDD.n3365 GND 0.004404f
C4943 VDD.n3366 GND 0.004404f
C4944 VDD.n3367 GND 0.274991f
C4945 VDD.n3368 GND 0.004404f
C4946 VDD.n3369 GND 0.004404f
C4947 VDD.n3370 GND 0.004404f
C4948 VDD.n3371 GND 0.004404f
C4949 VDD.n3372 GND 0.004404f
C4950 VDD.n3373 GND 0.292178f
C4951 VDD.n3374 GND 0.004404f
C4952 VDD.n3375 GND 0.004404f
C4953 VDD.n3376 GND 0.004404f
C4954 VDD.n3377 GND 0.004404f
C4955 VDD.n3378 GND 0.004404f
C4956 VDD.n3379 GND 0.292178f
C4957 VDD.n3380 GND 0.004404f
C4958 VDD.n3381 GND 0.004404f
C4959 VDD.n3382 GND 0.004404f
C4960 VDD.n3383 GND 0.004404f
C4961 VDD.n3384 GND 0.004404f
C4962 VDD.n3385 GND 0.292178f
C4963 VDD.n3386 GND 0.004404f
C4964 VDD.n3387 GND 0.004404f
C4965 VDD.n3388 GND 0.004404f
C4966 VDD.n3389 GND 0.004404f
C4967 VDD.n3390 GND 0.004404f
C4968 VDD.n3391 GND 0.259953f
C4969 VDD.n3392 GND 0.004404f
C4970 VDD.n3393 GND 0.004404f
C4971 VDD.n3394 GND 0.004404f
C4972 VDD.n3395 GND 0.004404f
C4973 VDD.n3396 GND 0.004404f
C4974 VDD.n3397 GND 0.292178f
C4975 VDD.n3398 GND 0.004404f
C4976 VDD.n3399 GND 0.004404f
C4977 VDD.n3400 GND 0.004404f
C4978 VDD.n3401 GND 0.004404f
C4979 VDD.n3402 GND 0.004404f
C4980 VDD.n3403 GND 0.21054f
C4981 VDD.n3404 GND 0.004404f
C4982 VDD.n3405 GND 0.004404f
C4983 VDD.n3406 GND 0.004404f
C4984 VDD.n3407 GND 0.004404f
C4985 VDD.n3408 GND 0.004404f
C4986 VDD.n3409 GND 0.292178f
C4987 VDD.n3410 GND 0.004404f
C4988 VDD.n3411 GND 0.004404f
C4989 VDD.n3412 GND 0.004404f
C4990 VDD.n3413 GND 0.004404f
C4991 VDD.n3414 GND 0.004404f
C4992 VDD.n3415 GND 0.292178f
C4993 VDD.n3416 GND 0.004404f
C4994 VDD.n3417 GND 0.004404f
C4995 VDD.n3418 GND 0.004404f
C4996 VDD.n3419 GND 0.004404f
C4997 VDD.n3420 GND 0.004404f
C4998 VDD.n3421 GND 0.292178f
C4999 VDD.n3422 GND 0.004404f
C5000 VDD.n3423 GND 0.004404f
C5001 VDD.n3424 GND 0.004404f
C5002 VDD.n3425 GND 0.004404f
C5003 VDD.n3426 GND 0.004404f
C5004 VDD.n3427 GND 0.004404f
C5005 VDD.n3428 GND 0.004404f
C5006 VDD.n3429 GND 0.004404f
C5007 VDD.n3430 GND 0.004404f
C5008 VDD.n3431 GND 0.004404f
C5009 VDD.n3432 GND 0.195502f
C5010 VDD.n3433 GND 0.004404f
C5011 VDD.n3434 GND 0.004404f
C5012 VDD.n3435 GND 0.004404f
C5013 VDD.n3436 GND 0.004404f
C5014 VDD.n3437 GND 0.004404f
C5015 VDD.n3438 GND 0.292178f
C5016 VDD.n3439 GND 0.004404f
C5017 VDD.n3440 GND 0.004404f
C5018 VDD.n3441 GND 0.004404f
C5019 VDD.n3442 GND 0.004404f
C5020 VDD.n3443 GND 0.004404f
C5021 VDD.n3444 GND 0.004404f
C5022 VDD.n3445 GND 0.004404f
C5023 VDD.n3446 GND 0.004404f
C5024 VDD.n3447 GND 0.004404f
C5025 VDD.n3448 GND 0.004404f
C5026 VDD.n3449 GND 0.004404f
C5027 VDD.n3450 GND 0.004404f
C5028 VDD.n3451 GND 0.004404f
C5029 VDD.n3452 GND 0.004404f
C5030 VDD.n3453 GND 0.004404f
C5031 VDD.n3454 GND 0.004404f
C5032 VDD.n3455 GND 0.004404f
C5033 VDD.n3456 GND 0.004404f
C5034 VDD.n3457 GND 0.004404f
C5035 VDD.n3458 GND 0.004404f
C5036 VDD.n3459 GND 0.004404f
C5037 VDD.n3460 GND 0.004404f
C5038 VDD.n3461 GND 0.004404f
C5039 VDD.n3462 GND 0.004404f
C5040 VDD.n3463 GND 0.004404f
C5041 VDD.n3464 GND 0.004404f
C5042 VDD.n3465 GND 0.004404f
C5043 VDD.n3466 GND 0.004404f
C5044 VDD.n3467 GND 0.004404f
C5045 VDD.n3468 GND 0.004404f
C5046 VDD.n3469 GND 0.004404f
C5047 VDD.n3470 GND 0.004404f
C5048 VDD.n3471 GND 0.004404f
C5049 VDD.n3472 GND 0.004404f
C5050 VDD.n3473 GND 0.004404f
C5051 VDD.n3474 GND 0.004404f
C5052 VDD.n3475 GND 0.004404f
C5053 VDD.n3476 GND 0.004404f
C5054 VDD.n3477 GND 0.004404f
C5055 VDD.n3478 GND 0.004404f
C5056 VDD.n3479 GND 0.004404f
C5057 VDD.n3480 GND 0.004404f
C5058 VDD.n3481 GND 0.004404f
C5059 VDD.n3482 GND 0.004404f
C5060 VDD.n3483 GND 0.004404f
C5061 VDD.n3484 GND 0.004404f
C5062 VDD.n3485 GND 0.004404f
C5063 VDD.n3486 GND 0.004404f
C5064 VDD.n3487 GND 0.004404f
C5065 VDD.n3488 GND 0.004404f
C5066 VDD.n3489 GND 0.004404f
C5067 VDD.n3490 GND 0.004404f
C5068 VDD.n3491 GND 0.004404f
C5069 VDD.n3492 GND 0.004404f
C5070 VDD.n3493 GND 0.004404f
C5071 VDD.n3494 GND 0.004404f
C5072 VDD.n3495 GND 0.004404f
C5073 VDD.n3496 GND 0.004404f
C5074 VDD.n3497 GND 0.004404f
C5075 VDD.n3498 GND 0.004404f
C5076 VDD.n3499 GND 0.004404f
C5077 VDD.n3500 GND 0.004404f
C5078 VDD.n3501 GND 0.004404f
C5079 VDD.n3502 GND 0.004404f
C5080 VDD.n3503 GND 0.004404f
C5081 VDD.n3504 GND 0.004404f
C5082 VDD.n3505 GND 0.004404f
C5083 VDD.n3506 GND 0.004404f
C5084 VDD.n3507 GND 0.004404f
C5085 VDD.n3508 GND 0.004404f
C5086 VDD.n3509 GND 0.004404f
C5087 VDD.t16 GND 0.292178f
C5088 VDD.n3510 GND 0.004404f
C5089 VDD.n3511 GND 0.004404f
C5090 VDD.n3512 GND 0.004404f
C5091 VDD.n3513 GND 0.004404f
C5092 VDD.n3514 GND 0.004404f
C5093 VDD.n3515 GND 0.292178f
C5094 VDD.n3516 GND 0.004404f
C5095 VDD.n3517 GND 0.004404f
C5096 VDD.n3518 GND 0.004404f
C5097 VDD.n3519 GND 0.004404f
C5098 VDD.n3520 GND 0.004404f
C5099 VDD.n3521 GND 0.292178f
C5100 VDD.n3522 GND 0.004404f
C5101 VDD.n3523 GND 0.004404f
C5102 VDD.n3524 GND 0.004404f
C5103 VDD.n3525 GND 0.004404f
C5104 VDD.n3526 GND 0.004404f
C5105 VDD.n3527 GND 0.292178f
C5106 VDD.n3528 GND 0.004404f
C5107 VDD.n3529 GND 0.004404f
C5108 VDD.n3530 GND 0.004404f
C5109 VDD.n3531 GND 0.004404f
C5110 VDD.n3532 GND 0.004404f
C5111 VDD.n3533 GND 0.292178f
C5112 VDD.n3534 GND 0.004404f
C5113 VDD.n3535 GND 0.004404f
C5114 VDD.n3536 GND 0.004404f
C5115 VDD.n3537 GND 0.004404f
C5116 VDD.n3538 GND 0.004404f
C5117 VDD.n3539 GND 0.292178f
C5118 VDD.n3540 GND 0.004404f
C5119 VDD.n3541 GND 0.004404f
C5120 VDD.n3542 GND 0.004404f
C5121 VDD.n3543 GND 0.004404f
C5122 VDD.n3544 GND 0.004404f
C5123 VDD.n3545 GND 0.21054f
C5124 VDD.n3546 GND 0.004404f
C5125 VDD.n3547 GND 0.004404f
C5126 VDD.n3548 GND 0.004404f
C5127 VDD.n3549 GND 0.004404f
C5128 VDD.n3550 GND 0.004404f
C5129 VDD.n3551 GND 0.212689f
C5130 VDD.n3552 GND 0.004404f
C5131 VDD.n3553 GND 0.004404f
C5132 VDD.n3554 GND 0.004404f
C5133 VDD.n3555 GND 0.004404f
C5134 VDD.n3556 GND 0.004404f
C5135 VDD.n3557 GND 0.292178f
C5136 VDD.n3558 GND 0.004404f
C5137 VDD.n3559 GND 0.004404f
C5138 VDD.n3560 GND 0.004404f
C5139 VDD.n3561 GND 0.004404f
C5140 VDD.n3562 GND 0.004404f
C5141 VDD.n3563 GND 0.292178f
C5142 VDD.n3564 GND 0.004404f
C5143 VDD.n3565 GND 0.004404f
C5144 VDD.n3566 GND 0.004404f
C5145 VDD.n3567 GND 0.004404f
C5146 VDD.n3568 GND 0.004404f
C5147 VDD.n3569 GND 0.292178f
C5148 VDD.n3570 GND 0.004404f
C5149 VDD.n3571 GND 0.004404f
C5150 VDD.n3572 GND 0.004404f
C5151 VDD.n3573 GND 0.004404f
C5152 VDD.n3574 GND 0.004404f
C5153 VDD.n3575 GND 0.292178f
C5154 VDD.n3576 GND 0.004404f
C5155 VDD.n3577 GND 0.004404f
C5156 VDD.n3578 GND 0.004404f
C5157 VDD.n3579 GND 0.004404f
C5158 VDD.n3580 GND 0.004404f
C5159 VDD.n3581 GND 0.274991f
C5160 VDD.n3582 GND 0.004404f
C5161 VDD.n3583 GND 0.004404f
C5162 VDD.n3584 GND 0.004404f
C5163 VDD.n3585 GND 0.004404f
C5164 VDD.n3586 GND 0.004404f
C5165 VDD.n3587 GND 0.27714f
C5166 VDD.n3588 GND 0.004404f
C5167 VDD.n3589 GND 0.004404f
C5168 VDD.n3590 GND 0.004404f
C5169 VDD.n3591 GND 0.004404f
C5170 VDD.n3592 GND 0.004404f
C5171 VDD.n3593 GND 0.292178f
C5172 VDD.n3594 GND 0.004404f
C5173 VDD.n3595 GND 0.004404f
C5174 VDD.n3596 GND 0.004404f
C5175 VDD.n3597 GND 0.004404f
C5176 VDD.n3598 GND 0.004404f
C5177 VDD.n3599 GND 0.292178f
C5178 VDD.n3600 GND 0.004404f
C5179 VDD.n3601 GND 0.004404f
C5180 VDD.n3602 GND 0.004404f
C5181 VDD.n3603 GND 0.004404f
C5182 VDD.n3604 GND 0.004404f
C5183 VDD.n3605 GND 0.292178f
C5184 VDD.n3606 GND 0.004404f
C5185 VDD.n3607 GND 0.004404f
C5186 VDD.n3608 GND 0.004404f
C5187 VDD.n3609 GND 0.004404f
C5188 VDD.n3610 GND 0.004404f
C5189 VDD.n3611 GND 0.292178f
C5190 VDD.n3612 GND 0.004404f
C5191 VDD.n3613 GND 0.004404f
C5192 VDD.n3614 GND 0.004404f
C5193 VDD.n3615 GND 0.004404f
C5194 VDD.n3616 GND 0.004404f
C5195 VDD.n3617 GND 0.292178f
C5196 VDD.n3618 GND 0.004404f
C5197 VDD.n3619 GND 0.004404f
C5198 VDD.n3620 GND 0.004404f
C5199 VDD.n3621 GND 0.004404f
C5200 VDD.n3622 GND 0.004404f
C5201 VDD.n3623 GND 0.292178f
C5202 VDD.n3624 GND 0.004404f
C5203 VDD.n3625 GND 0.004404f
C5204 VDD.n3626 GND 0.004404f
C5205 VDD.n3627 GND 0.004404f
C5206 VDD.n3628 GND 0.004404f
C5207 VDD.n3629 GND 0.174018f
C5208 VDD.n3630 GND 0.004404f
C5209 VDD.n3631 GND 0.004404f
C5210 VDD.n3632 GND 0.004404f
C5211 VDD.n3633 GND 0.004404f
C5212 VDD.n3634 GND 0.004404f
C5213 VDD.n3635 GND 0.292178f
C5214 VDD.n3636 GND 0.004404f
C5215 VDD.n3637 GND 0.004404f
C5216 VDD.n3638 GND 0.004404f
C5217 VDD.n3639 GND 0.004404f
C5218 VDD.n3640 GND 0.004404f
C5219 VDD.n3641 GND 0.004404f
C5220 VDD.n3642 GND 0.004404f
C5221 VDD.n3645 GND 0.004404f
C5222 VDD.n3646 GND 0.004404f
C5223 VDD.n3647 GND 0.004404f
C5224 VDD.n3648 GND 0.004404f
C5225 VDD.n3650 GND 0.004404f
C5226 VDD.n3651 GND 0.004404f
C5227 VDD.n3652 GND 0.004404f
C5228 VDD.n3653 GND 0.004404f
C5229 VDD.n3654 GND 0.004404f
C5230 VDD.n3655 GND 0.004404f
C5231 VDD.n3657 GND 0.004404f
C5232 VDD.n3658 GND 0.004404f
C5233 VDD.n3660 GND 0.01038f
C5234 VDD.n3661 GND 0.01038f
C5235 VDD.n3662 GND 0.010151f
C5236 VDD.n3663 GND 0.004404f
C5237 VDD.n3664 GND 0.004404f
C5238 VDD.n3665 GND 0.004404f
C5239 VDD.n3666 GND 0.004404f
C5240 VDD.n3667 GND 0.004404f
C5241 VDD.n3668 GND 0.004404f
C5242 VDD.n3669 GND 0.292178f
C5243 VDD.n3670 GND 0.004404f
C5244 VDD.n3671 GND 0.004404f
C5245 VDD.n3672 GND 0.004404f
C5246 VDD.n3673 GND 0.004404f
C5247 VDD.n3674 GND 0.004404f
C5248 VDD.n3675 GND 0.292178f
C5249 VDD.n3676 GND 0.004404f
C5250 VDD.n3677 GND 0.004404f
C5251 VDD.n3678 GND 0.004404f
C5252 VDD.n3679 GND 0.010674f
C5253 VDD.n3680 GND 0.009857f
C5254 VDD.n3681 GND 0.01038f
C5255 VDD.n3683 GND 0.004404f
C5256 VDD.n3684 GND 0.004404f
C5257 VDD.n3685 GND 0.002753f
C5258 VDD.n3686 GND 0.006294f
C5259 VDD.n3687 GND 0.003854f
C5260 VDD.n3688 GND 0.004404f
C5261 VDD.n3689 GND 0.004404f
C5262 VDD.n3691 GND 0.004404f
C5263 VDD.n3692 GND 0.004404f
C5264 VDD.n3693 GND 0.004404f
C5265 VDD.n3694 GND 0.004404f
C5266 VDD.n3695 GND 0.004404f
C5267 VDD.n3696 GND 0.004404f
C5268 VDD.n3698 GND 0.004404f
C5269 VDD.n3699 GND 0.004404f
C5270 VDD.n3700 GND 0.003303f
C5271 VDD.n3701 GND 0.004404f
C5272 VDD.n3702 GND 0.004404f
C5273 VDD.n3703 GND 0.004404f
C5274 VDD.n3705 GND 0.004404f
C5275 VDD.n3706 GND 0.004404f
C5276 VDD.n3707 GND 0.004404f
C5277 VDD.n3708 GND 0.004404f
C5278 VDD.n3709 GND 0.004404f
C5279 VDD.n3710 GND 0.004404f
C5280 VDD.n3712 GND 0.004404f
C5281 VDD.n3713 GND 0.004404f
C5282 VDD.n3714 GND 0.004404f
C5283 VDD.n3715 GND 0.01038f
C5284 VDD.n3716 GND 0.010151f
C5285 VDD.n3717 GND 0.010151f
C5286 VDD.n3718 GND 0.388855f
C5287 VDD.n3719 GND 0.010151f
C5288 VDD.n3720 GND 0.01038f
C5289 VDD.n3721 GND 0.009857f
C5290 VDD.n3722 GND 0.004404f
C5291 VDD.n3723 GND 0.002753f
C5292 VDD.n3724 GND 0.004404f
C5293 VDD.n3726 GND 0.004404f
C5294 VDD.n3727 GND 0.004404f
C5295 VDD.n3728 GND 0.004404f
C5296 VDD.n3729 GND 0.004404f
C5297 VDD.n3730 GND 0.004404f
C5298 VDD.n3731 GND 0.004404f
C5299 VDD.n3733 GND 0.004404f
C5300 VDD.n3734 GND 0.004404f
C5301 VDD.n3736 GND 0.004404f
C5302 VDD.n3737 GND 0.003303f
C5303 VDD.n3738 GND 0.03002f
C5304 VDD.n3739 GND 0.762058f
C5305 VDD.n3740 GND 0.008008f
C5306 VDD.n3741 GND 0.006477f
C5307 VDD.n3742 GND 0.005213f
C5308 VDD.n3743 GND 0.006477f
C5309 VDD.n3744 GND 0.429674f
C5310 VDD.n3745 GND 0.006477f
C5311 VDD.n3746 GND 0.005213f
C5312 VDD.n3747 GND 0.006477f
C5313 VDD.n3748 GND 0.006477f
C5314 VDD.n3749 GND 0.006477f
C5315 VDD.n3750 GND 0.005213f
C5316 VDD.n3751 GND 0.006477f
C5317 VDD.n3752 GND 0.429674f
C5318 VDD.n3753 GND 0.006477f
C5319 VDD.n3754 GND 0.005213f
C5320 VDD.n3755 GND 0.006477f
C5321 VDD.n3756 GND 0.006477f
C5322 VDD.n3757 GND 0.006477f
C5323 VDD.n3758 GND 0.005213f
C5324 VDD.n3759 GND 0.006477f
C5325 VDD.t94 GND 0.214837f
C5326 VDD.n3760 GND 0.399597f
C5327 VDD.n3761 GND 0.006477f
C5328 VDD.n3762 GND 0.005213f
C5329 VDD.n3763 GND 0.006477f
C5330 VDD.n3764 GND 0.006477f
C5331 VDD.n3765 GND 0.006477f
C5332 VDD.n3766 GND 0.005213f
C5333 VDD.n3767 GND 0.006477f
C5334 VDD.n3768 GND 0.429674f
C5335 VDD.n3769 GND 0.006477f
C5336 VDD.n3770 GND 0.005213f
C5337 VDD.n3771 GND 0.006477f
C5338 VDD.n3772 GND 0.006477f
C5339 VDD.n3773 GND 0.006477f
C5340 VDD.n3774 GND 0.005213f
C5341 VDD.n3775 GND 0.006477f
C5342 VDD.n3776 GND 0.429674f
C5343 VDD.n3777 GND 0.006477f
C5344 VDD.n3778 GND 0.005213f
C5345 VDD.n3779 GND 0.006477f
C5346 VDD.n3780 GND 0.006477f
C5347 VDD.n3781 GND 0.006477f
C5348 VDD.n3782 GND 0.005213f
C5349 VDD.n3783 GND 0.006477f
C5350 VDD.n3784 GND 0.429674f
C5351 VDD.n3785 GND 0.006477f
C5352 VDD.n3786 GND 0.005213f
C5353 VDD.n3787 GND 0.006477f
C5354 VDD.n3788 GND 0.006477f
C5355 VDD.n3789 GND 0.006477f
C5356 VDD.n3790 GND 0.005213f
C5357 VDD.n3791 GND 0.006477f
C5358 VDD.n3792 GND 0.429674f
C5359 VDD.n3793 GND 0.006477f
C5360 VDD.n3794 GND 0.005213f
C5361 VDD.n3795 GND 0.006477f
C5362 VDD.n3796 GND 0.006477f
C5363 VDD.n3797 GND 0.006477f
C5364 VDD.n3798 GND 0.005213f
C5365 VDD.n3799 GND 0.006477f
C5366 VDD.n3800 GND 0.429674f
C5367 VDD.n3801 GND 0.006477f
C5368 VDD.n3802 GND 0.005213f
C5369 VDD.n3803 GND 0.006477f
C5370 VDD.n3804 GND 0.006477f
C5371 VDD.n3805 GND 0.006477f
C5372 VDD.n3806 GND 0.005213f
C5373 VDD.n3807 GND 0.006477f
C5374 VDD.n3808 GND 0.429674f
C5375 VDD.n3809 GND 0.006477f
C5376 VDD.n3810 GND 0.005213f
C5377 VDD.n3811 GND 0.006477f
C5378 VDD.n3812 GND 0.006477f
C5379 VDD.n3813 GND 0.006477f
C5380 VDD.n3814 GND 0.005213f
C5381 VDD.n3815 GND 0.006477f
C5382 VDD.n3816 GND 0.274991f
C5383 VDD.n3817 GND 0.006477f
C5384 VDD.n3818 GND 0.005213f
C5385 VDD.n3819 GND 0.006477f
C5386 VDD.n3820 GND 0.006477f
C5387 VDD.n3821 GND 0.006477f
C5388 VDD.n3822 GND 0.005213f
C5389 VDD.n3823 GND 0.006477f
C5390 VDD.n3824 GND 0.429674f
C5391 VDD.n3825 GND 0.006477f
C5392 VDD.n3826 GND 0.005213f
C5393 VDD.n3827 GND 0.006477f
C5394 VDD.n3828 GND 0.006477f
C5395 VDD.n3829 GND 0.006477f
C5396 VDD.n3830 GND 0.005213f
C5397 VDD.n3831 GND 0.006477f
C5398 VDD.n3832 GND 0.429674f
C5399 VDD.n3833 GND 0.006477f
C5400 VDD.n3834 GND 0.005213f
C5401 VDD.n3835 GND 0.006477f
C5402 VDD.n3836 GND 0.006477f
C5403 VDD.n3837 GND 0.006477f
C5404 VDD.n3838 GND 0.005213f
C5405 VDD.n3839 GND 0.006477f
C5406 VDD.n3840 GND 0.429674f
C5407 VDD.n3841 GND 0.006477f
C5408 VDD.n3842 GND 0.005213f
C5409 VDD.n3843 GND 0.006477f
C5410 VDD.n3844 GND 0.006477f
C5411 VDD.n3845 GND 0.006477f
C5412 VDD.n3846 GND 0.005213f
C5413 VDD.n3847 GND 0.006477f
C5414 VDD.n3848 GND 0.429674f
C5415 VDD.n3849 GND 0.006477f
C5416 VDD.n3850 GND 0.005213f
C5417 VDD.n3851 GND 0.006477f
C5418 VDD.n3852 GND 0.006477f
C5419 VDD.n3853 GND 0.006477f
C5420 VDD.n3854 GND 0.005213f
C5421 VDD.n3855 GND 0.006477f
C5422 VDD.n3856 GND 0.326552f
C5423 VDD.n3857 GND 0.429674f
C5424 VDD.n3858 GND 0.006477f
C5425 VDD.n3859 GND 0.005213f
C5426 VDD.n3860 GND 0.006477f
C5427 VDD.n3861 GND 0.006477f
C5428 VDD.n3862 GND 0.006477f
C5429 VDD.n3863 GND 0.005213f
C5430 VDD.n3864 GND 0.006477f
C5431 VDD.n3865 GND 0.317959f
C5432 VDD.n3866 GND 0.006477f
C5433 VDD.n3867 GND 0.005213f
C5434 VDD.n3868 GND 0.006477f
C5435 VDD.n3869 GND 0.006477f
C5436 VDD.n3870 GND 0.006477f
C5437 VDD.n3871 GND 0.005213f
C5438 VDD.n3872 GND 0.006477f
C5439 VDD.n3873 GND 0.429674f
C5440 VDD.n3874 GND 0.006477f
C5441 VDD.n3875 GND 0.005213f
C5442 VDD.n3876 GND 0.006477f
C5443 VDD.n3877 GND 0.006477f
C5444 VDD.n3878 GND 0.006477f
C5445 VDD.n3879 GND 0.005213f
C5446 VDD.n3880 GND 0.006477f
C5447 VDD.n3881 GND 0.429674f
C5448 VDD.n3882 GND 0.006477f
C5449 VDD.n3883 GND 0.005213f
C5450 VDD.n3884 GND 0.006477f
C5451 VDD.n3885 GND 0.006477f
C5452 VDD.n3886 GND 0.006477f
C5453 VDD.n3887 GND 0.005213f
C5454 VDD.n3888 GND 0.006477f
C5455 VDD.n3889 GND 0.429674f
C5456 VDD.n3890 GND 0.006477f
C5457 VDD.n3891 GND 0.005213f
C5458 VDD.n3892 GND 0.006477f
C5459 VDD.n3893 GND 0.006477f
C5460 VDD.n3894 GND 0.006477f
C5461 VDD.n3895 GND 0.005213f
C5462 VDD.n3896 GND 0.006477f
C5463 VDD.n3897 GND 0.429674f
C5464 VDD.n3898 GND 0.006477f
C5465 VDD.n3899 GND 0.005213f
C5466 VDD.n3900 GND 0.006477f
C5467 VDD.n3901 GND 0.006477f
C5468 VDD.n3902 GND 0.006477f
C5469 VDD.n3903 GND 0.005213f
C5470 VDD.n3904 GND 0.006477f
C5471 VDD.t47 GND 0.214837f
C5472 VDD.n3905 GND 0.378113f
C5473 VDD.n3906 GND 0.006477f
C5474 VDD.n3907 GND 0.005213f
C5475 VDD.n3908 GND 0.006477f
C5476 VDD.n3909 GND 0.006477f
C5477 VDD.n3910 GND 0.006477f
C5478 VDD.n3911 GND 0.005213f
C5479 VDD.n3912 GND 0.006477f
C5480 VDD.n3913 GND 0.429674f
C5481 VDD.n3914 GND 0.006477f
C5482 VDD.n3915 GND 0.005213f
C5483 VDD.n3916 GND 0.006477f
C5484 VDD.n3917 GND 0.006477f
C5485 VDD.n3918 GND 0.006477f
C5486 VDD.n3919 GND 0.005213f
C5487 VDD.n3920 GND 0.006477f
C5488 VDD.n3921 GND 0.429674f
C5489 VDD.n3922 GND 0.006477f
C5490 VDD.n3923 GND 0.005213f
C5491 VDD.n3924 GND 0.006477f
C5492 VDD.n3925 GND 0.006477f
C5493 VDD.n3926 GND 0.006477f
C5494 VDD.n3927 GND 0.005213f
C5495 VDD.n3928 GND 0.006477f
C5496 VDD.n3929 GND 0.429674f
C5497 VDD.n3930 GND 0.006477f
C5498 VDD.n3931 GND 0.005213f
C5499 VDD.n3932 GND 0.006477f
C5500 VDD.n3933 GND 0.006477f
C5501 VDD.n3934 GND 0.006477f
C5502 VDD.n3935 GND 0.006477f
C5503 VDD.n3936 GND 0.006477f
C5504 VDD.n3937 GND 0.005213f
C5505 VDD.n3938 GND 0.005213f
C5506 VDD.n3939 GND 0.006477f
C5507 VDD.n3940 GND 0.429674f
C5508 VDD.n3941 GND 0.006477f
C5509 VDD.n3942 GND 0.005213f
C5510 VDD.n3943 GND 0.006477f
C5511 VDD.n3944 GND 0.006477f
C5512 VDD.n3945 GND 0.006477f
C5513 VDD.n3946 GND 0.005213f
C5514 VDD.n3947 GND 0.006477f
C5515 VDD.n3948 GND 0.429674f
C5516 VDD.n3949 GND 0.006477f
C5517 VDD.n3950 GND 0.006477f
C5518 VDD.n3951 GND 0.005213f
C5519 VDD.n3952 GND 0.005213f
C5520 VDD.n3953 GND 0.005213f
C5521 VDD.n3954 GND 0.006477f
C5522 VDD.n3955 GND 0.006477f
C5523 VDD.n3956 GND 0.006477f
C5524 VDD.n3957 GND 0.006477f
C5525 VDD.n3958 GND 0.005213f
C5526 VDD.n3959 GND 0.005213f
C5527 VDD.n3960 GND 0.005213f
C5528 VDD.n3961 GND 0.006477f
C5529 VDD.n3962 GND 0.006477f
C5530 VDD.n3963 GND 0.006477f
C5531 VDD.n3964 GND 0.006477f
C5532 VDD.n3965 GND 0.005213f
C5533 VDD.n3966 GND 0.005213f
C5534 VDD.n3967 GND 0.005213f
C5535 VDD.n3968 GND 0.006477f
C5536 VDD.n3969 GND 0.006477f
C5537 VDD.n3970 GND 0.006477f
C5538 VDD.n3971 GND 0.006477f
C5539 VDD.n3972 GND 0.005213f
C5540 VDD.n3973 GND 0.005213f
C5541 VDD.n3974 GND 0.005213f
C5542 VDD.n3975 GND 0.006477f
C5543 VDD.n3976 GND 0.006477f
C5544 VDD.n3977 GND 0.006477f
C5545 VDD.n3978 GND 0.006477f
C5546 VDD.n3979 GND 0.005213f
C5547 VDD.n3980 GND 0.005213f
C5548 VDD.n3981 GND 0.005213f
C5549 VDD.n3982 GND 0.006477f
C5550 VDD.n3983 GND 0.006477f
C5551 VDD.n3984 GND 0.006477f
C5552 VDD.n3985 GND 0.006477f
C5553 VDD.n3986 GND 0.005213f
C5554 VDD.n3987 GND 0.005213f
C5555 VDD.n3988 GND 0.005213f
C5556 VDD.n3989 GND 0.006477f
C5557 VDD.n3990 GND 0.006477f
C5558 VDD.n3991 GND 0.006477f
C5559 VDD.n3992 GND 0.006477f
C5560 VDD.n3993 GND 0.005213f
C5561 VDD.n3994 GND 0.005213f
C5562 VDD.n3995 GND 0.005213f
C5563 VDD.n3996 GND 0.006477f
C5564 VDD.n3997 GND 0.006477f
C5565 VDD.n3998 GND 0.006477f
C5566 VDD.n3999 GND 0.006477f
C5567 VDD.n4000 GND 0.005213f
C5568 VDD.n4001 GND 0.005213f
C5569 VDD.n4002 GND 0.005213f
C5570 VDD.n4003 GND 0.006477f
C5571 VDD.n4004 GND 0.006477f
C5572 VDD.n4005 GND 0.006477f
C5573 VDD.n4006 GND 0.006477f
C5574 VDD.n4007 GND 0.005213f
C5575 VDD.n4008 GND 0.005213f
C5576 VDD.n4009 GND 0.005213f
C5577 VDD.n4010 GND 0.006477f
C5578 VDD.n4011 GND 0.006477f
C5579 VDD.n4012 GND 0.006477f
C5580 VDD.n4013 GND 0.006477f
C5581 VDD.n4014 GND 0.005213f
C5582 VDD.n4015 GND 0.005213f
C5583 VDD.n4016 GND 0.005213f
C5584 VDD.n4017 GND 0.006477f
C5585 VDD.n4018 GND 0.006477f
C5586 VDD.n4019 GND 0.006477f
C5587 VDD.n4020 GND 0.006477f
C5588 VDD.n4021 GND 0.005213f
C5589 VDD.n4022 GND 0.005213f
C5590 VDD.n4023 GND 0.005213f
C5591 VDD.n4024 GND 0.006477f
C5592 VDD.n4025 GND 0.006477f
C5593 VDD.n4026 GND 0.006477f
C5594 VDD.n4027 GND 0.006477f
C5595 VDD.n4028 GND 0.005213f
C5596 VDD.n4029 GND 0.005213f
C5597 VDD.n4030 GND 0.005213f
C5598 VDD.n4031 GND 0.006477f
C5599 VDD.n4032 GND 0.006477f
C5600 VDD.n4033 GND 0.006477f
C5601 VDD.n4034 GND 0.006477f
C5602 VDD.n4035 GND 0.005213f
C5603 VDD.n4036 GND 0.005213f
C5604 VDD.n4037 GND 0.005213f
C5605 VDD.n4038 GND 0.006477f
C5606 VDD.n4039 GND 0.006477f
C5607 VDD.n4040 GND 0.006477f
C5608 VDD.n4041 GND 0.006477f
C5609 VDD.n4042 GND 0.005213f
C5610 VDD.n4043 GND 0.005213f
C5611 VDD.n4044 GND 0.004327f
C5612 VDD.n4045 GND 0.014826f
C5613 VDD.n4046 GND 0.014967f
C5614 VDD.n4047 GND 0.002502f
C5615 VDD.n4048 GND 0.014967f
C5616 VDD.n4050 GND 0.966767f
C5617 VDD.n4051 GND 0.575763f
C5618 VDD.n4052 GND 0.429674f
C5619 VDD.n4053 GND 0.006477f
C5620 VDD.n4054 GND 0.005213f
C5621 VDD.n4055 GND 0.005213f
C5622 VDD.n4056 GND 0.005213f
C5623 VDD.n4057 GND 0.006477f
C5624 VDD.n4058 GND 0.429674f
C5625 VDD.n4059 GND 0.429674f
C5626 VDD.n4060 GND 0.399597f
C5627 VDD.n4061 GND 0.006477f
C5628 VDD.n4062 GND 0.005213f
C5629 VDD.n4063 GND 0.005213f
C5630 VDD.n4064 GND 0.005213f
C5631 VDD.n4065 GND 0.006477f
C5632 VDD.n4066 GND 0.429674f
C5633 VDD.n4067 GND 0.429674f
C5634 VDD.n4068 GND 0.429674f
C5635 VDD.n4069 GND 0.006477f
C5636 VDD.n4070 GND 0.005213f
C5637 VDD.n4071 GND 0.005213f
C5638 VDD.n4072 GND 0.005213f
C5639 VDD.n4073 GND 0.006477f
C5640 VDD.n4074 GND 0.429674f
C5641 VDD.n4075 GND 0.429674f
C5642 VDD.n4076 GND 0.429674f
C5643 VDD.n4077 GND 0.006477f
C5644 VDD.n4078 GND 0.005213f
C5645 VDD.n4079 GND 0.005213f
C5646 VDD.n4080 GND 0.005213f
C5647 VDD.n4081 GND 0.006477f
C5648 VDD.n4082 GND 0.429674f
C5649 VDD.n4083 GND 0.429674f
C5650 VDD.n4084 GND 0.429674f
C5651 VDD.n4085 GND 0.006477f
C5652 VDD.n4086 GND 0.005213f
C5653 VDD.n4087 GND 0.005213f
C5654 VDD.n4088 GND 0.005213f
C5655 VDD.n4089 GND 0.006477f
C5656 VDD.n4090 GND 0.274991f
C5657 VDD.t7 GND 0.214837f
C5658 VDD.n4091 GND 0.36952f
C5659 VDD.n4092 GND 0.429674f
C5660 VDD.n4093 GND 0.006477f
C5661 VDD.n4094 GND 0.005213f
C5662 VDD.n4095 GND 0.005213f
C5663 VDD.n4096 GND 0.005213f
C5664 VDD.n4097 GND 0.006477f
C5665 VDD.n4098 GND 0.429674f
C5666 VDD.n4099 GND 0.429674f
C5667 VDD.n4100 GND 0.429674f
C5668 VDD.n4101 GND 0.006477f
C5669 VDD.n4102 GND 0.005213f
C5670 VDD.n4103 GND 0.005213f
C5671 VDD.n4104 GND 0.005213f
C5672 VDD.n4105 GND 0.006477f
C5673 VDD.n4106 GND 0.429674f
C5674 VDD.n4107 GND 0.429674f
C5675 VDD.n4108 GND 0.429674f
C5676 VDD.n4109 GND 0.006477f
C5677 VDD.n4110 GND 0.005213f
C5678 VDD.n4111 GND 0.005213f
C5679 VDD.n4112 GND 0.005213f
C5680 VDD.n4113 GND 0.006477f
C5681 VDD.n4114 GND 0.317959f
C5682 VDD.n4115 GND 0.429674f
C5683 VDD.n4116 GND 0.429674f
C5684 VDD.n4117 GND 0.006477f
C5685 VDD.n4118 GND 0.005213f
C5686 VDD.n4119 GND 0.005213f
C5687 VDD.n4120 GND 0.005213f
C5688 VDD.n4121 GND 0.006477f
C5689 VDD.n4122 GND 0.429674f
C5690 VDD.n4123 GND 0.429674f
C5691 VDD.n4124 GND 0.429674f
C5692 VDD.n4125 GND 0.006477f
C5693 VDD.n4126 GND 0.005213f
C5694 VDD.n4127 GND 0.005213f
C5695 VDD.n4128 GND 0.005213f
C5696 VDD.n4129 GND 0.006477f
C5697 VDD.n4130 GND 0.429674f
C5698 VDD.n4131 GND 0.429674f
C5699 VDD.n4132 GND 0.378113f
C5700 VDD.n4133 GND 0.006477f
C5701 VDD.n4134 GND 0.005213f
C5702 VDD.n4135 GND 0.005213f
C5703 VDD.n4136 GND 0.005213f
C5704 VDD.n4137 GND 0.006477f
C5705 VDD.n4138 GND 0.429674f
C5706 VDD.n4139 GND 0.429674f
C5707 VDD.n4140 GND 0.429674f
C5708 VDD.n4141 GND 0.006477f
C5709 VDD.n4142 GND 0.005213f
C5710 VDD.n4143 GND 0.005213f
C5711 VDD.n4144 GND 0.005213f
C5712 VDD.n4145 GND 0.006477f
C5713 VDD.n4146 GND 0.429674f
C5714 VDD.n4147 GND 0.429674f
C5715 VDD.n4148 GND 0.429674f
C5716 VDD.n4149 GND 0.006477f
C5717 VDD.n4150 GND 0.005213f
C5718 VDD.n4151 GND 0.005213f
C5719 VDD.n4152 GND 0.005213f
C5720 VDD.n4153 GND 0.006477f
C5721 VDD.n4154 GND 0.429674f
C5722 VDD.n4155 GND 0.429674f
C5723 VDD.t23 GND 0.429674f
C5724 VDD.n4156 GND 0.006477f
C5725 VDD.n4157 GND 0.005213f
C5726 VDD.n4158 GND 0.46472f
C5727 VDD.n4159 GND 3.32995f
.ends

