* NGSPICE file created from diff_pair_sample_1306.ext - technology: sky130A

.subckt diff_pair_sample_1306 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=3.8
X1 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=3.8
X2 VDD1.t3 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=3.8
X3 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=3.8
X4 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=3.8
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=3.8
X6 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=3.8
X7 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=3.8
X8 VTAIL.t5 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=3.8
X9 VDD1.t0 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=3.8
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=3.8
X11 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=3.8
R0 VP.n21 VP.n20 161.3
R1 VP.n19 VP.n1 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n16 VP.n2 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n3 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n4 161.3
R8 VP.n9 VP.n8 161.3
R9 VP.n5 VP.t0 110.745
R10 VP.n5 VP.t1 109.395
R11 VP.n7 VP.n6 86.8867
R12 VP.n22 VP.n0 86.8867
R13 VP.n7 VP.t2 76.8034
R14 VP.n0 VP.t3 76.8034
R15 VP.n6 VP.n5 51.9839
R16 VP.n14 VP.n13 40.4934
R17 VP.n14 VP.n2 40.4934
R18 VP.n8 VP.n4 24.4675
R19 VP.n12 VP.n4 24.4675
R20 VP.n13 VP.n12 24.4675
R21 VP.n18 VP.n2 24.4675
R22 VP.n19 VP.n18 24.4675
R23 VP.n20 VP.n19 24.4675
R24 VP.n8 VP.n7 3.18121
R25 VP.n20 VP.n0 3.18121
R26 VP.n9 VP.n6 0.354971
R27 VP.n22 VP.n21 0.354971
R28 VP VP.n22 0.26696
R29 VP.n10 VP.n9 0.189894
R30 VP.n11 VP.n10 0.189894
R31 VP.n11 VP.n3 0.189894
R32 VP.n15 VP.n3 0.189894
R33 VP.n16 VP.n15 0.189894
R34 VP.n17 VP.n16 0.189894
R35 VP.n17 VP.n1 0.189894
R36 VP.n21 VP.n1 0.189894
R37 VDD1 VDD1.n1 107.046
R38 VDD1 VDD1.n0 61.744
R39 VDD1.n0 VDD1.t2 1.63551
R40 VDD1.n0 VDD1.t3 1.63551
R41 VDD1.n1 VDD1.t1 1.63551
R42 VDD1.n1 VDD1.t0 1.63551
R43 VTAIL.n522 VTAIL.n462 289.615
R44 VTAIL.n60 VTAIL.n0 289.615
R45 VTAIL.n126 VTAIL.n66 289.615
R46 VTAIL.n192 VTAIL.n132 289.615
R47 VTAIL.n456 VTAIL.n396 289.615
R48 VTAIL.n390 VTAIL.n330 289.615
R49 VTAIL.n324 VTAIL.n264 289.615
R50 VTAIL.n258 VTAIL.n198 289.615
R51 VTAIL.n482 VTAIL.n481 185
R52 VTAIL.n487 VTAIL.n486 185
R53 VTAIL.n489 VTAIL.n488 185
R54 VTAIL.n478 VTAIL.n477 185
R55 VTAIL.n495 VTAIL.n494 185
R56 VTAIL.n497 VTAIL.n496 185
R57 VTAIL.n474 VTAIL.n473 185
R58 VTAIL.n504 VTAIL.n503 185
R59 VTAIL.n505 VTAIL.n472 185
R60 VTAIL.n507 VTAIL.n506 185
R61 VTAIL.n470 VTAIL.n469 185
R62 VTAIL.n513 VTAIL.n512 185
R63 VTAIL.n515 VTAIL.n514 185
R64 VTAIL.n466 VTAIL.n465 185
R65 VTAIL.n521 VTAIL.n520 185
R66 VTAIL.n523 VTAIL.n522 185
R67 VTAIL.n20 VTAIL.n19 185
R68 VTAIL.n25 VTAIL.n24 185
R69 VTAIL.n27 VTAIL.n26 185
R70 VTAIL.n16 VTAIL.n15 185
R71 VTAIL.n33 VTAIL.n32 185
R72 VTAIL.n35 VTAIL.n34 185
R73 VTAIL.n12 VTAIL.n11 185
R74 VTAIL.n42 VTAIL.n41 185
R75 VTAIL.n43 VTAIL.n10 185
R76 VTAIL.n45 VTAIL.n44 185
R77 VTAIL.n8 VTAIL.n7 185
R78 VTAIL.n51 VTAIL.n50 185
R79 VTAIL.n53 VTAIL.n52 185
R80 VTAIL.n4 VTAIL.n3 185
R81 VTAIL.n59 VTAIL.n58 185
R82 VTAIL.n61 VTAIL.n60 185
R83 VTAIL.n86 VTAIL.n85 185
R84 VTAIL.n91 VTAIL.n90 185
R85 VTAIL.n93 VTAIL.n92 185
R86 VTAIL.n82 VTAIL.n81 185
R87 VTAIL.n99 VTAIL.n98 185
R88 VTAIL.n101 VTAIL.n100 185
R89 VTAIL.n78 VTAIL.n77 185
R90 VTAIL.n108 VTAIL.n107 185
R91 VTAIL.n109 VTAIL.n76 185
R92 VTAIL.n111 VTAIL.n110 185
R93 VTAIL.n74 VTAIL.n73 185
R94 VTAIL.n117 VTAIL.n116 185
R95 VTAIL.n119 VTAIL.n118 185
R96 VTAIL.n70 VTAIL.n69 185
R97 VTAIL.n125 VTAIL.n124 185
R98 VTAIL.n127 VTAIL.n126 185
R99 VTAIL.n152 VTAIL.n151 185
R100 VTAIL.n157 VTAIL.n156 185
R101 VTAIL.n159 VTAIL.n158 185
R102 VTAIL.n148 VTAIL.n147 185
R103 VTAIL.n165 VTAIL.n164 185
R104 VTAIL.n167 VTAIL.n166 185
R105 VTAIL.n144 VTAIL.n143 185
R106 VTAIL.n174 VTAIL.n173 185
R107 VTAIL.n175 VTAIL.n142 185
R108 VTAIL.n177 VTAIL.n176 185
R109 VTAIL.n140 VTAIL.n139 185
R110 VTAIL.n183 VTAIL.n182 185
R111 VTAIL.n185 VTAIL.n184 185
R112 VTAIL.n136 VTAIL.n135 185
R113 VTAIL.n191 VTAIL.n190 185
R114 VTAIL.n193 VTAIL.n192 185
R115 VTAIL.n457 VTAIL.n456 185
R116 VTAIL.n455 VTAIL.n454 185
R117 VTAIL.n400 VTAIL.n399 185
R118 VTAIL.n449 VTAIL.n448 185
R119 VTAIL.n447 VTAIL.n446 185
R120 VTAIL.n404 VTAIL.n403 185
R121 VTAIL.n441 VTAIL.n440 185
R122 VTAIL.n439 VTAIL.n406 185
R123 VTAIL.n438 VTAIL.n437 185
R124 VTAIL.n409 VTAIL.n407 185
R125 VTAIL.n432 VTAIL.n431 185
R126 VTAIL.n430 VTAIL.n429 185
R127 VTAIL.n413 VTAIL.n412 185
R128 VTAIL.n424 VTAIL.n423 185
R129 VTAIL.n422 VTAIL.n421 185
R130 VTAIL.n417 VTAIL.n416 185
R131 VTAIL.n391 VTAIL.n390 185
R132 VTAIL.n389 VTAIL.n388 185
R133 VTAIL.n334 VTAIL.n333 185
R134 VTAIL.n383 VTAIL.n382 185
R135 VTAIL.n381 VTAIL.n380 185
R136 VTAIL.n338 VTAIL.n337 185
R137 VTAIL.n375 VTAIL.n374 185
R138 VTAIL.n373 VTAIL.n340 185
R139 VTAIL.n372 VTAIL.n371 185
R140 VTAIL.n343 VTAIL.n341 185
R141 VTAIL.n366 VTAIL.n365 185
R142 VTAIL.n364 VTAIL.n363 185
R143 VTAIL.n347 VTAIL.n346 185
R144 VTAIL.n358 VTAIL.n357 185
R145 VTAIL.n356 VTAIL.n355 185
R146 VTAIL.n351 VTAIL.n350 185
R147 VTAIL.n325 VTAIL.n324 185
R148 VTAIL.n323 VTAIL.n322 185
R149 VTAIL.n268 VTAIL.n267 185
R150 VTAIL.n317 VTAIL.n316 185
R151 VTAIL.n315 VTAIL.n314 185
R152 VTAIL.n272 VTAIL.n271 185
R153 VTAIL.n309 VTAIL.n308 185
R154 VTAIL.n307 VTAIL.n274 185
R155 VTAIL.n306 VTAIL.n305 185
R156 VTAIL.n277 VTAIL.n275 185
R157 VTAIL.n300 VTAIL.n299 185
R158 VTAIL.n298 VTAIL.n297 185
R159 VTAIL.n281 VTAIL.n280 185
R160 VTAIL.n292 VTAIL.n291 185
R161 VTAIL.n290 VTAIL.n289 185
R162 VTAIL.n285 VTAIL.n284 185
R163 VTAIL.n259 VTAIL.n258 185
R164 VTAIL.n257 VTAIL.n256 185
R165 VTAIL.n202 VTAIL.n201 185
R166 VTAIL.n251 VTAIL.n250 185
R167 VTAIL.n249 VTAIL.n248 185
R168 VTAIL.n206 VTAIL.n205 185
R169 VTAIL.n243 VTAIL.n242 185
R170 VTAIL.n241 VTAIL.n208 185
R171 VTAIL.n240 VTAIL.n239 185
R172 VTAIL.n211 VTAIL.n209 185
R173 VTAIL.n234 VTAIL.n233 185
R174 VTAIL.n232 VTAIL.n231 185
R175 VTAIL.n215 VTAIL.n214 185
R176 VTAIL.n226 VTAIL.n225 185
R177 VTAIL.n224 VTAIL.n223 185
R178 VTAIL.n219 VTAIL.n218 185
R179 VTAIL.n483 VTAIL.t3 149.524
R180 VTAIL.n21 VTAIL.t2 149.524
R181 VTAIL.n87 VTAIL.t4 149.524
R182 VTAIL.n153 VTAIL.t5 149.524
R183 VTAIL.n418 VTAIL.t6 149.524
R184 VTAIL.n352 VTAIL.t7 149.524
R185 VTAIL.n286 VTAIL.t1 149.524
R186 VTAIL.n220 VTAIL.t0 149.524
R187 VTAIL.n487 VTAIL.n481 104.615
R188 VTAIL.n488 VTAIL.n487 104.615
R189 VTAIL.n488 VTAIL.n477 104.615
R190 VTAIL.n495 VTAIL.n477 104.615
R191 VTAIL.n496 VTAIL.n495 104.615
R192 VTAIL.n496 VTAIL.n473 104.615
R193 VTAIL.n504 VTAIL.n473 104.615
R194 VTAIL.n505 VTAIL.n504 104.615
R195 VTAIL.n506 VTAIL.n505 104.615
R196 VTAIL.n506 VTAIL.n469 104.615
R197 VTAIL.n513 VTAIL.n469 104.615
R198 VTAIL.n514 VTAIL.n513 104.615
R199 VTAIL.n514 VTAIL.n465 104.615
R200 VTAIL.n521 VTAIL.n465 104.615
R201 VTAIL.n522 VTAIL.n521 104.615
R202 VTAIL.n25 VTAIL.n19 104.615
R203 VTAIL.n26 VTAIL.n25 104.615
R204 VTAIL.n26 VTAIL.n15 104.615
R205 VTAIL.n33 VTAIL.n15 104.615
R206 VTAIL.n34 VTAIL.n33 104.615
R207 VTAIL.n34 VTAIL.n11 104.615
R208 VTAIL.n42 VTAIL.n11 104.615
R209 VTAIL.n43 VTAIL.n42 104.615
R210 VTAIL.n44 VTAIL.n43 104.615
R211 VTAIL.n44 VTAIL.n7 104.615
R212 VTAIL.n51 VTAIL.n7 104.615
R213 VTAIL.n52 VTAIL.n51 104.615
R214 VTAIL.n52 VTAIL.n3 104.615
R215 VTAIL.n59 VTAIL.n3 104.615
R216 VTAIL.n60 VTAIL.n59 104.615
R217 VTAIL.n91 VTAIL.n85 104.615
R218 VTAIL.n92 VTAIL.n91 104.615
R219 VTAIL.n92 VTAIL.n81 104.615
R220 VTAIL.n99 VTAIL.n81 104.615
R221 VTAIL.n100 VTAIL.n99 104.615
R222 VTAIL.n100 VTAIL.n77 104.615
R223 VTAIL.n108 VTAIL.n77 104.615
R224 VTAIL.n109 VTAIL.n108 104.615
R225 VTAIL.n110 VTAIL.n109 104.615
R226 VTAIL.n110 VTAIL.n73 104.615
R227 VTAIL.n117 VTAIL.n73 104.615
R228 VTAIL.n118 VTAIL.n117 104.615
R229 VTAIL.n118 VTAIL.n69 104.615
R230 VTAIL.n125 VTAIL.n69 104.615
R231 VTAIL.n126 VTAIL.n125 104.615
R232 VTAIL.n157 VTAIL.n151 104.615
R233 VTAIL.n158 VTAIL.n157 104.615
R234 VTAIL.n158 VTAIL.n147 104.615
R235 VTAIL.n165 VTAIL.n147 104.615
R236 VTAIL.n166 VTAIL.n165 104.615
R237 VTAIL.n166 VTAIL.n143 104.615
R238 VTAIL.n174 VTAIL.n143 104.615
R239 VTAIL.n175 VTAIL.n174 104.615
R240 VTAIL.n176 VTAIL.n175 104.615
R241 VTAIL.n176 VTAIL.n139 104.615
R242 VTAIL.n183 VTAIL.n139 104.615
R243 VTAIL.n184 VTAIL.n183 104.615
R244 VTAIL.n184 VTAIL.n135 104.615
R245 VTAIL.n191 VTAIL.n135 104.615
R246 VTAIL.n192 VTAIL.n191 104.615
R247 VTAIL.n456 VTAIL.n455 104.615
R248 VTAIL.n455 VTAIL.n399 104.615
R249 VTAIL.n448 VTAIL.n399 104.615
R250 VTAIL.n448 VTAIL.n447 104.615
R251 VTAIL.n447 VTAIL.n403 104.615
R252 VTAIL.n440 VTAIL.n403 104.615
R253 VTAIL.n440 VTAIL.n439 104.615
R254 VTAIL.n439 VTAIL.n438 104.615
R255 VTAIL.n438 VTAIL.n407 104.615
R256 VTAIL.n431 VTAIL.n407 104.615
R257 VTAIL.n431 VTAIL.n430 104.615
R258 VTAIL.n430 VTAIL.n412 104.615
R259 VTAIL.n423 VTAIL.n412 104.615
R260 VTAIL.n423 VTAIL.n422 104.615
R261 VTAIL.n422 VTAIL.n416 104.615
R262 VTAIL.n390 VTAIL.n389 104.615
R263 VTAIL.n389 VTAIL.n333 104.615
R264 VTAIL.n382 VTAIL.n333 104.615
R265 VTAIL.n382 VTAIL.n381 104.615
R266 VTAIL.n381 VTAIL.n337 104.615
R267 VTAIL.n374 VTAIL.n337 104.615
R268 VTAIL.n374 VTAIL.n373 104.615
R269 VTAIL.n373 VTAIL.n372 104.615
R270 VTAIL.n372 VTAIL.n341 104.615
R271 VTAIL.n365 VTAIL.n341 104.615
R272 VTAIL.n365 VTAIL.n364 104.615
R273 VTAIL.n364 VTAIL.n346 104.615
R274 VTAIL.n357 VTAIL.n346 104.615
R275 VTAIL.n357 VTAIL.n356 104.615
R276 VTAIL.n356 VTAIL.n350 104.615
R277 VTAIL.n324 VTAIL.n323 104.615
R278 VTAIL.n323 VTAIL.n267 104.615
R279 VTAIL.n316 VTAIL.n267 104.615
R280 VTAIL.n316 VTAIL.n315 104.615
R281 VTAIL.n315 VTAIL.n271 104.615
R282 VTAIL.n308 VTAIL.n271 104.615
R283 VTAIL.n308 VTAIL.n307 104.615
R284 VTAIL.n307 VTAIL.n306 104.615
R285 VTAIL.n306 VTAIL.n275 104.615
R286 VTAIL.n299 VTAIL.n275 104.615
R287 VTAIL.n299 VTAIL.n298 104.615
R288 VTAIL.n298 VTAIL.n280 104.615
R289 VTAIL.n291 VTAIL.n280 104.615
R290 VTAIL.n291 VTAIL.n290 104.615
R291 VTAIL.n290 VTAIL.n284 104.615
R292 VTAIL.n258 VTAIL.n257 104.615
R293 VTAIL.n257 VTAIL.n201 104.615
R294 VTAIL.n250 VTAIL.n201 104.615
R295 VTAIL.n250 VTAIL.n249 104.615
R296 VTAIL.n249 VTAIL.n205 104.615
R297 VTAIL.n242 VTAIL.n205 104.615
R298 VTAIL.n242 VTAIL.n241 104.615
R299 VTAIL.n241 VTAIL.n240 104.615
R300 VTAIL.n240 VTAIL.n209 104.615
R301 VTAIL.n233 VTAIL.n209 104.615
R302 VTAIL.n233 VTAIL.n232 104.615
R303 VTAIL.n232 VTAIL.n214 104.615
R304 VTAIL.n225 VTAIL.n214 104.615
R305 VTAIL.n225 VTAIL.n224 104.615
R306 VTAIL.n224 VTAIL.n218 104.615
R307 VTAIL.t3 VTAIL.n481 52.3082
R308 VTAIL.t2 VTAIL.n19 52.3082
R309 VTAIL.t4 VTAIL.n85 52.3082
R310 VTAIL.t5 VTAIL.n151 52.3082
R311 VTAIL.t6 VTAIL.n416 52.3082
R312 VTAIL.t7 VTAIL.n350 52.3082
R313 VTAIL.t1 VTAIL.n284 52.3082
R314 VTAIL.t0 VTAIL.n218 52.3082
R315 VTAIL.n527 VTAIL.n526 31.9914
R316 VTAIL.n65 VTAIL.n64 31.9914
R317 VTAIL.n131 VTAIL.n130 31.9914
R318 VTAIL.n197 VTAIL.n196 31.9914
R319 VTAIL.n461 VTAIL.n460 31.9914
R320 VTAIL.n395 VTAIL.n394 31.9914
R321 VTAIL.n329 VTAIL.n328 31.9914
R322 VTAIL.n263 VTAIL.n262 31.9914
R323 VTAIL.n527 VTAIL.n461 26.3669
R324 VTAIL.n263 VTAIL.n197 26.3669
R325 VTAIL.n507 VTAIL.n472 13.1884
R326 VTAIL.n45 VTAIL.n10 13.1884
R327 VTAIL.n111 VTAIL.n76 13.1884
R328 VTAIL.n177 VTAIL.n142 13.1884
R329 VTAIL.n441 VTAIL.n406 13.1884
R330 VTAIL.n375 VTAIL.n340 13.1884
R331 VTAIL.n309 VTAIL.n274 13.1884
R332 VTAIL.n243 VTAIL.n208 13.1884
R333 VTAIL.n503 VTAIL.n502 12.8005
R334 VTAIL.n508 VTAIL.n470 12.8005
R335 VTAIL.n41 VTAIL.n40 12.8005
R336 VTAIL.n46 VTAIL.n8 12.8005
R337 VTAIL.n107 VTAIL.n106 12.8005
R338 VTAIL.n112 VTAIL.n74 12.8005
R339 VTAIL.n173 VTAIL.n172 12.8005
R340 VTAIL.n178 VTAIL.n140 12.8005
R341 VTAIL.n442 VTAIL.n404 12.8005
R342 VTAIL.n437 VTAIL.n408 12.8005
R343 VTAIL.n376 VTAIL.n338 12.8005
R344 VTAIL.n371 VTAIL.n342 12.8005
R345 VTAIL.n310 VTAIL.n272 12.8005
R346 VTAIL.n305 VTAIL.n276 12.8005
R347 VTAIL.n244 VTAIL.n206 12.8005
R348 VTAIL.n239 VTAIL.n210 12.8005
R349 VTAIL.n501 VTAIL.n474 12.0247
R350 VTAIL.n512 VTAIL.n511 12.0247
R351 VTAIL.n39 VTAIL.n12 12.0247
R352 VTAIL.n50 VTAIL.n49 12.0247
R353 VTAIL.n105 VTAIL.n78 12.0247
R354 VTAIL.n116 VTAIL.n115 12.0247
R355 VTAIL.n171 VTAIL.n144 12.0247
R356 VTAIL.n182 VTAIL.n181 12.0247
R357 VTAIL.n446 VTAIL.n445 12.0247
R358 VTAIL.n436 VTAIL.n409 12.0247
R359 VTAIL.n380 VTAIL.n379 12.0247
R360 VTAIL.n370 VTAIL.n343 12.0247
R361 VTAIL.n314 VTAIL.n313 12.0247
R362 VTAIL.n304 VTAIL.n277 12.0247
R363 VTAIL.n248 VTAIL.n247 12.0247
R364 VTAIL.n238 VTAIL.n211 12.0247
R365 VTAIL.n498 VTAIL.n497 11.249
R366 VTAIL.n515 VTAIL.n468 11.249
R367 VTAIL.n36 VTAIL.n35 11.249
R368 VTAIL.n53 VTAIL.n6 11.249
R369 VTAIL.n102 VTAIL.n101 11.249
R370 VTAIL.n119 VTAIL.n72 11.249
R371 VTAIL.n168 VTAIL.n167 11.249
R372 VTAIL.n185 VTAIL.n138 11.249
R373 VTAIL.n449 VTAIL.n402 11.249
R374 VTAIL.n433 VTAIL.n432 11.249
R375 VTAIL.n383 VTAIL.n336 11.249
R376 VTAIL.n367 VTAIL.n366 11.249
R377 VTAIL.n317 VTAIL.n270 11.249
R378 VTAIL.n301 VTAIL.n300 11.249
R379 VTAIL.n251 VTAIL.n204 11.249
R380 VTAIL.n235 VTAIL.n234 11.249
R381 VTAIL.n494 VTAIL.n476 10.4732
R382 VTAIL.n516 VTAIL.n466 10.4732
R383 VTAIL.n32 VTAIL.n14 10.4732
R384 VTAIL.n54 VTAIL.n4 10.4732
R385 VTAIL.n98 VTAIL.n80 10.4732
R386 VTAIL.n120 VTAIL.n70 10.4732
R387 VTAIL.n164 VTAIL.n146 10.4732
R388 VTAIL.n186 VTAIL.n136 10.4732
R389 VTAIL.n450 VTAIL.n400 10.4732
R390 VTAIL.n429 VTAIL.n411 10.4732
R391 VTAIL.n384 VTAIL.n334 10.4732
R392 VTAIL.n363 VTAIL.n345 10.4732
R393 VTAIL.n318 VTAIL.n268 10.4732
R394 VTAIL.n297 VTAIL.n279 10.4732
R395 VTAIL.n252 VTAIL.n202 10.4732
R396 VTAIL.n231 VTAIL.n213 10.4732
R397 VTAIL.n483 VTAIL.n482 10.2747
R398 VTAIL.n21 VTAIL.n20 10.2747
R399 VTAIL.n87 VTAIL.n86 10.2747
R400 VTAIL.n153 VTAIL.n152 10.2747
R401 VTAIL.n418 VTAIL.n417 10.2747
R402 VTAIL.n352 VTAIL.n351 10.2747
R403 VTAIL.n286 VTAIL.n285 10.2747
R404 VTAIL.n220 VTAIL.n219 10.2747
R405 VTAIL.n493 VTAIL.n478 9.69747
R406 VTAIL.n520 VTAIL.n519 9.69747
R407 VTAIL.n31 VTAIL.n16 9.69747
R408 VTAIL.n58 VTAIL.n57 9.69747
R409 VTAIL.n97 VTAIL.n82 9.69747
R410 VTAIL.n124 VTAIL.n123 9.69747
R411 VTAIL.n163 VTAIL.n148 9.69747
R412 VTAIL.n190 VTAIL.n189 9.69747
R413 VTAIL.n454 VTAIL.n453 9.69747
R414 VTAIL.n428 VTAIL.n413 9.69747
R415 VTAIL.n388 VTAIL.n387 9.69747
R416 VTAIL.n362 VTAIL.n347 9.69747
R417 VTAIL.n322 VTAIL.n321 9.69747
R418 VTAIL.n296 VTAIL.n281 9.69747
R419 VTAIL.n256 VTAIL.n255 9.69747
R420 VTAIL.n230 VTAIL.n215 9.69747
R421 VTAIL.n526 VTAIL.n525 9.45567
R422 VTAIL.n64 VTAIL.n63 9.45567
R423 VTAIL.n130 VTAIL.n129 9.45567
R424 VTAIL.n196 VTAIL.n195 9.45567
R425 VTAIL.n460 VTAIL.n459 9.45567
R426 VTAIL.n394 VTAIL.n393 9.45567
R427 VTAIL.n328 VTAIL.n327 9.45567
R428 VTAIL.n262 VTAIL.n261 9.45567
R429 VTAIL.n525 VTAIL.n524 9.3005
R430 VTAIL.n464 VTAIL.n463 9.3005
R431 VTAIL.n519 VTAIL.n518 9.3005
R432 VTAIL.n517 VTAIL.n516 9.3005
R433 VTAIL.n468 VTAIL.n467 9.3005
R434 VTAIL.n511 VTAIL.n510 9.3005
R435 VTAIL.n509 VTAIL.n508 9.3005
R436 VTAIL.n485 VTAIL.n484 9.3005
R437 VTAIL.n480 VTAIL.n479 9.3005
R438 VTAIL.n491 VTAIL.n490 9.3005
R439 VTAIL.n493 VTAIL.n492 9.3005
R440 VTAIL.n476 VTAIL.n475 9.3005
R441 VTAIL.n499 VTAIL.n498 9.3005
R442 VTAIL.n501 VTAIL.n500 9.3005
R443 VTAIL.n502 VTAIL.n471 9.3005
R444 VTAIL.n63 VTAIL.n62 9.3005
R445 VTAIL.n2 VTAIL.n1 9.3005
R446 VTAIL.n57 VTAIL.n56 9.3005
R447 VTAIL.n55 VTAIL.n54 9.3005
R448 VTAIL.n6 VTAIL.n5 9.3005
R449 VTAIL.n49 VTAIL.n48 9.3005
R450 VTAIL.n47 VTAIL.n46 9.3005
R451 VTAIL.n23 VTAIL.n22 9.3005
R452 VTAIL.n18 VTAIL.n17 9.3005
R453 VTAIL.n29 VTAIL.n28 9.3005
R454 VTAIL.n31 VTAIL.n30 9.3005
R455 VTAIL.n14 VTAIL.n13 9.3005
R456 VTAIL.n37 VTAIL.n36 9.3005
R457 VTAIL.n39 VTAIL.n38 9.3005
R458 VTAIL.n40 VTAIL.n9 9.3005
R459 VTAIL.n129 VTAIL.n128 9.3005
R460 VTAIL.n68 VTAIL.n67 9.3005
R461 VTAIL.n123 VTAIL.n122 9.3005
R462 VTAIL.n121 VTAIL.n120 9.3005
R463 VTAIL.n72 VTAIL.n71 9.3005
R464 VTAIL.n115 VTAIL.n114 9.3005
R465 VTAIL.n113 VTAIL.n112 9.3005
R466 VTAIL.n89 VTAIL.n88 9.3005
R467 VTAIL.n84 VTAIL.n83 9.3005
R468 VTAIL.n95 VTAIL.n94 9.3005
R469 VTAIL.n97 VTAIL.n96 9.3005
R470 VTAIL.n80 VTAIL.n79 9.3005
R471 VTAIL.n103 VTAIL.n102 9.3005
R472 VTAIL.n105 VTAIL.n104 9.3005
R473 VTAIL.n106 VTAIL.n75 9.3005
R474 VTAIL.n195 VTAIL.n194 9.3005
R475 VTAIL.n134 VTAIL.n133 9.3005
R476 VTAIL.n189 VTAIL.n188 9.3005
R477 VTAIL.n187 VTAIL.n186 9.3005
R478 VTAIL.n138 VTAIL.n137 9.3005
R479 VTAIL.n181 VTAIL.n180 9.3005
R480 VTAIL.n179 VTAIL.n178 9.3005
R481 VTAIL.n155 VTAIL.n154 9.3005
R482 VTAIL.n150 VTAIL.n149 9.3005
R483 VTAIL.n161 VTAIL.n160 9.3005
R484 VTAIL.n163 VTAIL.n162 9.3005
R485 VTAIL.n146 VTAIL.n145 9.3005
R486 VTAIL.n169 VTAIL.n168 9.3005
R487 VTAIL.n171 VTAIL.n170 9.3005
R488 VTAIL.n172 VTAIL.n141 9.3005
R489 VTAIL.n420 VTAIL.n419 9.3005
R490 VTAIL.n415 VTAIL.n414 9.3005
R491 VTAIL.n426 VTAIL.n425 9.3005
R492 VTAIL.n428 VTAIL.n427 9.3005
R493 VTAIL.n411 VTAIL.n410 9.3005
R494 VTAIL.n434 VTAIL.n433 9.3005
R495 VTAIL.n436 VTAIL.n435 9.3005
R496 VTAIL.n408 VTAIL.n405 9.3005
R497 VTAIL.n459 VTAIL.n458 9.3005
R498 VTAIL.n398 VTAIL.n397 9.3005
R499 VTAIL.n453 VTAIL.n452 9.3005
R500 VTAIL.n451 VTAIL.n450 9.3005
R501 VTAIL.n402 VTAIL.n401 9.3005
R502 VTAIL.n445 VTAIL.n444 9.3005
R503 VTAIL.n443 VTAIL.n442 9.3005
R504 VTAIL.n354 VTAIL.n353 9.3005
R505 VTAIL.n349 VTAIL.n348 9.3005
R506 VTAIL.n360 VTAIL.n359 9.3005
R507 VTAIL.n362 VTAIL.n361 9.3005
R508 VTAIL.n345 VTAIL.n344 9.3005
R509 VTAIL.n368 VTAIL.n367 9.3005
R510 VTAIL.n370 VTAIL.n369 9.3005
R511 VTAIL.n342 VTAIL.n339 9.3005
R512 VTAIL.n393 VTAIL.n392 9.3005
R513 VTAIL.n332 VTAIL.n331 9.3005
R514 VTAIL.n387 VTAIL.n386 9.3005
R515 VTAIL.n385 VTAIL.n384 9.3005
R516 VTAIL.n336 VTAIL.n335 9.3005
R517 VTAIL.n379 VTAIL.n378 9.3005
R518 VTAIL.n377 VTAIL.n376 9.3005
R519 VTAIL.n288 VTAIL.n287 9.3005
R520 VTAIL.n283 VTAIL.n282 9.3005
R521 VTAIL.n294 VTAIL.n293 9.3005
R522 VTAIL.n296 VTAIL.n295 9.3005
R523 VTAIL.n279 VTAIL.n278 9.3005
R524 VTAIL.n302 VTAIL.n301 9.3005
R525 VTAIL.n304 VTAIL.n303 9.3005
R526 VTAIL.n276 VTAIL.n273 9.3005
R527 VTAIL.n327 VTAIL.n326 9.3005
R528 VTAIL.n266 VTAIL.n265 9.3005
R529 VTAIL.n321 VTAIL.n320 9.3005
R530 VTAIL.n319 VTAIL.n318 9.3005
R531 VTAIL.n270 VTAIL.n269 9.3005
R532 VTAIL.n313 VTAIL.n312 9.3005
R533 VTAIL.n311 VTAIL.n310 9.3005
R534 VTAIL.n222 VTAIL.n221 9.3005
R535 VTAIL.n217 VTAIL.n216 9.3005
R536 VTAIL.n228 VTAIL.n227 9.3005
R537 VTAIL.n230 VTAIL.n229 9.3005
R538 VTAIL.n213 VTAIL.n212 9.3005
R539 VTAIL.n236 VTAIL.n235 9.3005
R540 VTAIL.n238 VTAIL.n237 9.3005
R541 VTAIL.n210 VTAIL.n207 9.3005
R542 VTAIL.n261 VTAIL.n260 9.3005
R543 VTAIL.n200 VTAIL.n199 9.3005
R544 VTAIL.n255 VTAIL.n254 9.3005
R545 VTAIL.n253 VTAIL.n252 9.3005
R546 VTAIL.n204 VTAIL.n203 9.3005
R547 VTAIL.n247 VTAIL.n246 9.3005
R548 VTAIL.n245 VTAIL.n244 9.3005
R549 VTAIL.n490 VTAIL.n489 8.92171
R550 VTAIL.n523 VTAIL.n464 8.92171
R551 VTAIL.n28 VTAIL.n27 8.92171
R552 VTAIL.n61 VTAIL.n2 8.92171
R553 VTAIL.n94 VTAIL.n93 8.92171
R554 VTAIL.n127 VTAIL.n68 8.92171
R555 VTAIL.n160 VTAIL.n159 8.92171
R556 VTAIL.n193 VTAIL.n134 8.92171
R557 VTAIL.n457 VTAIL.n398 8.92171
R558 VTAIL.n425 VTAIL.n424 8.92171
R559 VTAIL.n391 VTAIL.n332 8.92171
R560 VTAIL.n359 VTAIL.n358 8.92171
R561 VTAIL.n325 VTAIL.n266 8.92171
R562 VTAIL.n293 VTAIL.n292 8.92171
R563 VTAIL.n259 VTAIL.n200 8.92171
R564 VTAIL.n227 VTAIL.n226 8.92171
R565 VTAIL.n486 VTAIL.n480 8.14595
R566 VTAIL.n524 VTAIL.n462 8.14595
R567 VTAIL.n24 VTAIL.n18 8.14595
R568 VTAIL.n62 VTAIL.n0 8.14595
R569 VTAIL.n90 VTAIL.n84 8.14595
R570 VTAIL.n128 VTAIL.n66 8.14595
R571 VTAIL.n156 VTAIL.n150 8.14595
R572 VTAIL.n194 VTAIL.n132 8.14595
R573 VTAIL.n458 VTAIL.n396 8.14595
R574 VTAIL.n421 VTAIL.n415 8.14595
R575 VTAIL.n392 VTAIL.n330 8.14595
R576 VTAIL.n355 VTAIL.n349 8.14595
R577 VTAIL.n326 VTAIL.n264 8.14595
R578 VTAIL.n289 VTAIL.n283 8.14595
R579 VTAIL.n260 VTAIL.n198 8.14595
R580 VTAIL.n223 VTAIL.n217 8.14595
R581 VTAIL.n485 VTAIL.n482 7.3702
R582 VTAIL.n23 VTAIL.n20 7.3702
R583 VTAIL.n89 VTAIL.n86 7.3702
R584 VTAIL.n155 VTAIL.n152 7.3702
R585 VTAIL.n420 VTAIL.n417 7.3702
R586 VTAIL.n354 VTAIL.n351 7.3702
R587 VTAIL.n288 VTAIL.n285 7.3702
R588 VTAIL.n222 VTAIL.n219 7.3702
R589 VTAIL.n486 VTAIL.n485 5.81868
R590 VTAIL.n526 VTAIL.n462 5.81868
R591 VTAIL.n24 VTAIL.n23 5.81868
R592 VTAIL.n64 VTAIL.n0 5.81868
R593 VTAIL.n90 VTAIL.n89 5.81868
R594 VTAIL.n130 VTAIL.n66 5.81868
R595 VTAIL.n156 VTAIL.n155 5.81868
R596 VTAIL.n196 VTAIL.n132 5.81868
R597 VTAIL.n460 VTAIL.n396 5.81868
R598 VTAIL.n421 VTAIL.n420 5.81868
R599 VTAIL.n394 VTAIL.n330 5.81868
R600 VTAIL.n355 VTAIL.n354 5.81868
R601 VTAIL.n328 VTAIL.n264 5.81868
R602 VTAIL.n289 VTAIL.n288 5.81868
R603 VTAIL.n262 VTAIL.n198 5.81868
R604 VTAIL.n223 VTAIL.n222 5.81868
R605 VTAIL.n489 VTAIL.n480 5.04292
R606 VTAIL.n524 VTAIL.n523 5.04292
R607 VTAIL.n27 VTAIL.n18 5.04292
R608 VTAIL.n62 VTAIL.n61 5.04292
R609 VTAIL.n93 VTAIL.n84 5.04292
R610 VTAIL.n128 VTAIL.n127 5.04292
R611 VTAIL.n159 VTAIL.n150 5.04292
R612 VTAIL.n194 VTAIL.n193 5.04292
R613 VTAIL.n458 VTAIL.n457 5.04292
R614 VTAIL.n424 VTAIL.n415 5.04292
R615 VTAIL.n392 VTAIL.n391 5.04292
R616 VTAIL.n358 VTAIL.n349 5.04292
R617 VTAIL.n326 VTAIL.n325 5.04292
R618 VTAIL.n292 VTAIL.n283 5.04292
R619 VTAIL.n260 VTAIL.n259 5.04292
R620 VTAIL.n226 VTAIL.n217 5.04292
R621 VTAIL.n490 VTAIL.n478 4.26717
R622 VTAIL.n520 VTAIL.n464 4.26717
R623 VTAIL.n28 VTAIL.n16 4.26717
R624 VTAIL.n58 VTAIL.n2 4.26717
R625 VTAIL.n94 VTAIL.n82 4.26717
R626 VTAIL.n124 VTAIL.n68 4.26717
R627 VTAIL.n160 VTAIL.n148 4.26717
R628 VTAIL.n190 VTAIL.n134 4.26717
R629 VTAIL.n454 VTAIL.n398 4.26717
R630 VTAIL.n425 VTAIL.n413 4.26717
R631 VTAIL.n388 VTAIL.n332 4.26717
R632 VTAIL.n359 VTAIL.n347 4.26717
R633 VTAIL.n322 VTAIL.n266 4.26717
R634 VTAIL.n293 VTAIL.n281 4.26717
R635 VTAIL.n256 VTAIL.n200 4.26717
R636 VTAIL.n227 VTAIL.n215 4.26717
R637 VTAIL.n329 VTAIL.n263 3.56084
R638 VTAIL.n461 VTAIL.n395 3.56084
R639 VTAIL.n197 VTAIL.n131 3.56084
R640 VTAIL.n494 VTAIL.n493 3.49141
R641 VTAIL.n519 VTAIL.n466 3.49141
R642 VTAIL.n32 VTAIL.n31 3.49141
R643 VTAIL.n57 VTAIL.n4 3.49141
R644 VTAIL.n98 VTAIL.n97 3.49141
R645 VTAIL.n123 VTAIL.n70 3.49141
R646 VTAIL.n164 VTAIL.n163 3.49141
R647 VTAIL.n189 VTAIL.n136 3.49141
R648 VTAIL.n453 VTAIL.n400 3.49141
R649 VTAIL.n429 VTAIL.n428 3.49141
R650 VTAIL.n387 VTAIL.n334 3.49141
R651 VTAIL.n363 VTAIL.n362 3.49141
R652 VTAIL.n321 VTAIL.n268 3.49141
R653 VTAIL.n297 VTAIL.n296 3.49141
R654 VTAIL.n255 VTAIL.n202 3.49141
R655 VTAIL.n231 VTAIL.n230 3.49141
R656 VTAIL.n484 VTAIL.n483 2.84303
R657 VTAIL.n22 VTAIL.n21 2.84303
R658 VTAIL.n88 VTAIL.n87 2.84303
R659 VTAIL.n154 VTAIL.n153 2.84303
R660 VTAIL.n419 VTAIL.n418 2.84303
R661 VTAIL.n353 VTAIL.n352 2.84303
R662 VTAIL.n287 VTAIL.n286 2.84303
R663 VTAIL.n221 VTAIL.n220 2.84303
R664 VTAIL.n497 VTAIL.n476 2.71565
R665 VTAIL.n516 VTAIL.n515 2.71565
R666 VTAIL.n35 VTAIL.n14 2.71565
R667 VTAIL.n54 VTAIL.n53 2.71565
R668 VTAIL.n101 VTAIL.n80 2.71565
R669 VTAIL.n120 VTAIL.n119 2.71565
R670 VTAIL.n167 VTAIL.n146 2.71565
R671 VTAIL.n186 VTAIL.n185 2.71565
R672 VTAIL.n450 VTAIL.n449 2.71565
R673 VTAIL.n432 VTAIL.n411 2.71565
R674 VTAIL.n384 VTAIL.n383 2.71565
R675 VTAIL.n366 VTAIL.n345 2.71565
R676 VTAIL.n318 VTAIL.n317 2.71565
R677 VTAIL.n300 VTAIL.n279 2.71565
R678 VTAIL.n252 VTAIL.n251 2.71565
R679 VTAIL.n234 VTAIL.n213 2.71565
R680 VTAIL.n498 VTAIL.n474 1.93989
R681 VTAIL.n512 VTAIL.n468 1.93989
R682 VTAIL.n36 VTAIL.n12 1.93989
R683 VTAIL.n50 VTAIL.n6 1.93989
R684 VTAIL.n102 VTAIL.n78 1.93989
R685 VTAIL.n116 VTAIL.n72 1.93989
R686 VTAIL.n168 VTAIL.n144 1.93989
R687 VTAIL.n182 VTAIL.n138 1.93989
R688 VTAIL.n446 VTAIL.n402 1.93989
R689 VTAIL.n433 VTAIL.n409 1.93989
R690 VTAIL.n380 VTAIL.n336 1.93989
R691 VTAIL.n367 VTAIL.n343 1.93989
R692 VTAIL.n314 VTAIL.n270 1.93989
R693 VTAIL.n301 VTAIL.n277 1.93989
R694 VTAIL.n248 VTAIL.n204 1.93989
R695 VTAIL.n235 VTAIL.n211 1.93989
R696 VTAIL VTAIL.n65 1.83886
R697 VTAIL VTAIL.n527 1.72248
R698 VTAIL.n503 VTAIL.n501 1.16414
R699 VTAIL.n511 VTAIL.n470 1.16414
R700 VTAIL.n41 VTAIL.n39 1.16414
R701 VTAIL.n49 VTAIL.n8 1.16414
R702 VTAIL.n107 VTAIL.n105 1.16414
R703 VTAIL.n115 VTAIL.n74 1.16414
R704 VTAIL.n173 VTAIL.n171 1.16414
R705 VTAIL.n181 VTAIL.n140 1.16414
R706 VTAIL.n445 VTAIL.n404 1.16414
R707 VTAIL.n437 VTAIL.n436 1.16414
R708 VTAIL.n379 VTAIL.n338 1.16414
R709 VTAIL.n371 VTAIL.n370 1.16414
R710 VTAIL.n313 VTAIL.n272 1.16414
R711 VTAIL.n305 VTAIL.n304 1.16414
R712 VTAIL.n247 VTAIL.n206 1.16414
R713 VTAIL.n239 VTAIL.n238 1.16414
R714 VTAIL.n395 VTAIL.n329 0.470328
R715 VTAIL.n131 VTAIL.n65 0.470328
R716 VTAIL.n502 VTAIL.n472 0.388379
R717 VTAIL.n508 VTAIL.n507 0.388379
R718 VTAIL.n40 VTAIL.n10 0.388379
R719 VTAIL.n46 VTAIL.n45 0.388379
R720 VTAIL.n106 VTAIL.n76 0.388379
R721 VTAIL.n112 VTAIL.n111 0.388379
R722 VTAIL.n172 VTAIL.n142 0.388379
R723 VTAIL.n178 VTAIL.n177 0.388379
R724 VTAIL.n442 VTAIL.n441 0.388379
R725 VTAIL.n408 VTAIL.n406 0.388379
R726 VTAIL.n376 VTAIL.n375 0.388379
R727 VTAIL.n342 VTAIL.n340 0.388379
R728 VTAIL.n310 VTAIL.n309 0.388379
R729 VTAIL.n276 VTAIL.n274 0.388379
R730 VTAIL.n244 VTAIL.n243 0.388379
R731 VTAIL.n210 VTAIL.n208 0.388379
R732 VTAIL.n484 VTAIL.n479 0.155672
R733 VTAIL.n491 VTAIL.n479 0.155672
R734 VTAIL.n492 VTAIL.n491 0.155672
R735 VTAIL.n492 VTAIL.n475 0.155672
R736 VTAIL.n499 VTAIL.n475 0.155672
R737 VTAIL.n500 VTAIL.n499 0.155672
R738 VTAIL.n500 VTAIL.n471 0.155672
R739 VTAIL.n509 VTAIL.n471 0.155672
R740 VTAIL.n510 VTAIL.n509 0.155672
R741 VTAIL.n510 VTAIL.n467 0.155672
R742 VTAIL.n517 VTAIL.n467 0.155672
R743 VTAIL.n518 VTAIL.n517 0.155672
R744 VTAIL.n518 VTAIL.n463 0.155672
R745 VTAIL.n525 VTAIL.n463 0.155672
R746 VTAIL.n22 VTAIL.n17 0.155672
R747 VTAIL.n29 VTAIL.n17 0.155672
R748 VTAIL.n30 VTAIL.n29 0.155672
R749 VTAIL.n30 VTAIL.n13 0.155672
R750 VTAIL.n37 VTAIL.n13 0.155672
R751 VTAIL.n38 VTAIL.n37 0.155672
R752 VTAIL.n38 VTAIL.n9 0.155672
R753 VTAIL.n47 VTAIL.n9 0.155672
R754 VTAIL.n48 VTAIL.n47 0.155672
R755 VTAIL.n48 VTAIL.n5 0.155672
R756 VTAIL.n55 VTAIL.n5 0.155672
R757 VTAIL.n56 VTAIL.n55 0.155672
R758 VTAIL.n56 VTAIL.n1 0.155672
R759 VTAIL.n63 VTAIL.n1 0.155672
R760 VTAIL.n88 VTAIL.n83 0.155672
R761 VTAIL.n95 VTAIL.n83 0.155672
R762 VTAIL.n96 VTAIL.n95 0.155672
R763 VTAIL.n96 VTAIL.n79 0.155672
R764 VTAIL.n103 VTAIL.n79 0.155672
R765 VTAIL.n104 VTAIL.n103 0.155672
R766 VTAIL.n104 VTAIL.n75 0.155672
R767 VTAIL.n113 VTAIL.n75 0.155672
R768 VTAIL.n114 VTAIL.n113 0.155672
R769 VTAIL.n114 VTAIL.n71 0.155672
R770 VTAIL.n121 VTAIL.n71 0.155672
R771 VTAIL.n122 VTAIL.n121 0.155672
R772 VTAIL.n122 VTAIL.n67 0.155672
R773 VTAIL.n129 VTAIL.n67 0.155672
R774 VTAIL.n154 VTAIL.n149 0.155672
R775 VTAIL.n161 VTAIL.n149 0.155672
R776 VTAIL.n162 VTAIL.n161 0.155672
R777 VTAIL.n162 VTAIL.n145 0.155672
R778 VTAIL.n169 VTAIL.n145 0.155672
R779 VTAIL.n170 VTAIL.n169 0.155672
R780 VTAIL.n170 VTAIL.n141 0.155672
R781 VTAIL.n179 VTAIL.n141 0.155672
R782 VTAIL.n180 VTAIL.n179 0.155672
R783 VTAIL.n180 VTAIL.n137 0.155672
R784 VTAIL.n187 VTAIL.n137 0.155672
R785 VTAIL.n188 VTAIL.n187 0.155672
R786 VTAIL.n188 VTAIL.n133 0.155672
R787 VTAIL.n195 VTAIL.n133 0.155672
R788 VTAIL.n459 VTAIL.n397 0.155672
R789 VTAIL.n452 VTAIL.n397 0.155672
R790 VTAIL.n452 VTAIL.n451 0.155672
R791 VTAIL.n451 VTAIL.n401 0.155672
R792 VTAIL.n444 VTAIL.n401 0.155672
R793 VTAIL.n444 VTAIL.n443 0.155672
R794 VTAIL.n443 VTAIL.n405 0.155672
R795 VTAIL.n435 VTAIL.n405 0.155672
R796 VTAIL.n435 VTAIL.n434 0.155672
R797 VTAIL.n434 VTAIL.n410 0.155672
R798 VTAIL.n427 VTAIL.n410 0.155672
R799 VTAIL.n427 VTAIL.n426 0.155672
R800 VTAIL.n426 VTAIL.n414 0.155672
R801 VTAIL.n419 VTAIL.n414 0.155672
R802 VTAIL.n393 VTAIL.n331 0.155672
R803 VTAIL.n386 VTAIL.n331 0.155672
R804 VTAIL.n386 VTAIL.n385 0.155672
R805 VTAIL.n385 VTAIL.n335 0.155672
R806 VTAIL.n378 VTAIL.n335 0.155672
R807 VTAIL.n378 VTAIL.n377 0.155672
R808 VTAIL.n377 VTAIL.n339 0.155672
R809 VTAIL.n369 VTAIL.n339 0.155672
R810 VTAIL.n369 VTAIL.n368 0.155672
R811 VTAIL.n368 VTAIL.n344 0.155672
R812 VTAIL.n361 VTAIL.n344 0.155672
R813 VTAIL.n361 VTAIL.n360 0.155672
R814 VTAIL.n360 VTAIL.n348 0.155672
R815 VTAIL.n353 VTAIL.n348 0.155672
R816 VTAIL.n327 VTAIL.n265 0.155672
R817 VTAIL.n320 VTAIL.n265 0.155672
R818 VTAIL.n320 VTAIL.n319 0.155672
R819 VTAIL.n319 VTAIL.n269 0.155672
R820 VTAIL.n312 VTAIL.n269 0.155672
R821 VTAIL.n312 VTAIL.n311 0.155672
R822 VTAIL.n311 VTAIL.n273 0.155672
R823 VTAIL.n303 VTAIL.n273 0.155672
R824 VTAIL.n303 VTAIL.n302 0.155672
R825 VTAIL.n302 VTAIL.n278 0.155672
R826 VTAIL.n295 VTAIL.n278 0.155672
R827 VTAIL.n295 VTAIL.n294 0.155672
R828 VTAIL.n294 VTAIL.n282 0.155672
R829 VTAIL.n287 VTAIL.n282 0.155672
R830 VTAIL.n261 VTAIL.n199 0.155672
R831 VTAIL.n254 VTAIL.n199 0.155672
R832 VTAIL.n254 VTAIL.n253 0.155672
R833 VTAIL.n253 VTAIL.n203 0.155672
R834 VTAIL.n246 VTAIL.n203 0.155672
R835 VTAIL.n246 VTAIL.n245 0.155672
R836 VTAIL.n245 VTAIL.n207 0.155672
R837 VTAIL.n237 VTAIL.n207 0.155672
R838 VTAIL.n237 VTAIL.n236 0.155672
R839 VTAIL.n236 VTAIL.n212 0.155672
R840 VTAIL.n229 VTAIL.n212 0.155672
R841 VTAIL.n229 VTAIL.n228 0.155672
R842 VTAIL.n228 VTAIL.n216 0.155672
R843 VTAIL.n221 VTAIL.n216 0.155672
R844 B.n833 B.n832 585
R845 B.n834 B.n833 585
R846 B.n317 B.n130 585
R847 B.n316 B.n315 585
R848 B.n314 B.n313 585
R849 B.n312 B.n311 585
R850 B.n310 B.n309 585
R851 B.n308 B.n307 585
R852 B.n306 B.n305 585
R853 B.n304 B.n303 585
R854 B.n302 B.n301 585
R855 B.n300 B.n299 585
R856 B.n298 B.n297 585
R857 B.n296 B.n295 585
R858 B.n294 B.n293 585
R859 B.n292 B.n291 585
R860 B.n290 B.n289 585
R861 B.n288 B.n287 585
R862 B.n286 B.n285 585
R863 B.n284 B.n283 585
R864 B.n282 B.n281 585
R865 B.n280 B.n279 585
R866 B.n278 B.n277 585
R867 B.n276 B.n275 585
R868 B.n274 B.n273 585
R869 B.n272 B.n271 585
R870 B.n270 B.n269 585
R871 B.n268 B.n267 585
R872 B.n266 B.n265 585
R873 B.n264 B.n263 585
R874 B.n262 B.n261 585
R875 B.n260 B.n259 585
R876 B.n258 B.n257 585
R877 B.n256 B.n255 585
R878 B.n254 B.n253 585
R879 B.n252 B.n251 585
R880 B.n250 B.n249 585
R881 B.n248 B.n247 585
R882 B.n246 B.n245 585
R883 B.n244 B.n243 585
R884 B.n242 B.n241 585
R885 B.n240 B.n239 585
R886 B.n238 B.n237 585
R887 B.n235 B.n234 585
R888 B.n233 B.n232 585
R889 B.n231 B.n230 585
R890 B.n229 B.n228 585
R891 B.n227 B.n226 585
R892 B.n225 B.n224 585
R893 B.n223 B.n222 585
R894 B.n221 B.n220 585
R895 B.n219 B.n218 585
R896 B.n217 B.n216 585
R897 B.n215 B.n214 585
R898 B.n213 B.n212 585
R899 B.n211 B.n210 585
R900 B.n209 B.n208 585
R901 B.n207 B.n206 585
R902 B.n205 B.n204 585
R903 B.n203 B.n202 585
R904 B.n201 B.n200 585
R905 B.n199 B.n198 585
R906 B.n197 B.n196 585
R907 B.n195 B.n194 585
R908 B.n193 B.n192 585
R909 B.n191 B.n190 585
R910 B.n189 B.n188 585
R911 B.n187 B.n186 585
R912 B.n185 B.n184 585
R913 B.n183 B.n182 585
R914 B.n181 B.n180 585
R915 B.n179 B.n178 585
R916 B.n177 B.n176 585
R917 B.n175 B.n174 585
R918 B.n173 B.n172 585
R919 B.n171 B.n170 585
R920 B.n169 B.n168 585
R921 B.n167 B.n166 585
R922 B.n165 B.n164 585
R923 B.n163 B.n162 585
R924 B.n161 B.n160 585
R925 B.n159 B.n158 585
R926 B.n157 B.n156 585
R927 B.n155 B.n154 585
R928 B.n153 B.n152 585
R929 B.n151 B.n150 585
R930 B.n149 B.n148 585
R931 B.n147 B.n146 585
R932 B.n145 B.n144 585
R933 B.n143 B.n142 585
R934 B.n141 B.n140 585
R935 B.n139 B.n138 585
R936 B.n137 B.n136 585
R937 B.n82 B.n81 585
R938 B.n831 B.n83 585
R939 B.n835 B.n83 585
R940 B.n830 B.n829 585
R941 B.n829 B.n79 585
R942 B.n828 B.n78 585
R943 B.n841 B.n78 585
R944 B.n827 B.n77 585
R945 B.n842 B.n77 585
R946 B.n826 B.n76 585
R947 B.n843 B.n76 585
R948 B.n825 B.n824 585
R949 B.n824 B.n72 585
R950 B.n823 B.n71 585
R951 B.n849 B.n71 585
R952 B.n822 B.n70 585
R953 B.n850 B.n70 585
R954 B.n821 B.n69 585
R955 B.n851 B.n69 585
R956 B.n820 B.n819 585
R957 B.n819 B.n68 585
R958 B.n818 B.n64 585
R959 B.n857 B.n64 585
R960 B.n817 B.n63 585
R961 B.n858 B.n63 585
R962 B.n816 B.n62 585
R963 B.n859 B.n62 585
R964 B.n815 B.n814 585
R965 B.n814 B.n58 585
R966 B.n813 B.n57 585
R967 B.n865 B.n57 585
R968 B.n812 B.n56 585
R969 B.n866 B.n56 585
R970 B.n811 B.n55 585
R971 B.n867 B.n55 585
R972 B.n810 B.n809 585
R973 B.n809 B.n51 585
R974 B.n808 B.n50 585
R975 B.n873 B.n50 585
R976 B.n807 B.n49 585
R977 B.n874 B.n49 585
R978 B.n806 B.n48 585
R979 B.n875 B.n48 585
R980 B.n805 B.n804 585
R981 B.n804 B.n44 585
R982 B.n803 B.n43 585
R983 B.n881 B.n43 585
R984 B.n802 B.n42 585
R985 B.n882 B.n42 585
R986 B.n801 B.n41 585
R987 B.n883 B.n41 585
R988 B.n800 B.n799 585
R989 B.n799 B.n37 585
R990 B.n798 B.n36 585
R991 B.n889 B.n36 585
R992 B.n797 B.n35 585
R993 B.n890 B.n35 585
R994 B.n796 B.n34 585
R995 B.n891 B.n34 585
R996 B.n795 B.n794 585
R997 B.n794 B.n30 585
R998 B.n793 B.n29 585
R999 B.n897 B.n29 585
R1000 B.n792 B.n28 585
R1001 B.n898 B.n28 585
R1002 B.n791 B.n27 585
R1003 B.n899 B.n27 585
R1004 B.n790 B.n789 585
R1005 B.n789 B.n23 585
R1006 B.n788 B.n22 585
R1007 B.n905 B.n22 585
R1008 B.n787 B.n21 585
R1009 B.n906 B.n21 585
R1010 B.n786 B.n20 585
R1011 B.n907 B.n20 585
R1012 B.n785 B.n784 585
R1013 B.n784 B.n16 585
R1014 B.n783 B.n15 585
R1015 B.n913 B.n15 585
R1016 B.n782 B.n14 585
R1017 B.n914 B.n14 585
R1018 B.n781 B.n13 585
R1019 B.n915 B.n13 585
R1020 B.n780 B.n779 585
R1021 B.n779 B.n12 585
R1022 B.n778 B.n777 585
R1023 B.n778 B.n8 585
R1024 B.n776 B.n7 585
R1025 B.n922 B.n7 585
R1026 B.n775 B.n6 585
R1027 B.n923 B.n6 585
R1028 B.n774 B.n5 585
R1029 B.n924 B.n5 585
R1030 B.n773 B.n772 585
R1031 B.n772 B.n4 585
R1032 B.n771 B.n318 585
R1033 B.n771 B.n770 585
R1034 B.n761 B.n319 585
R1035 B.n320 B.n319 585
R1036 B.n763 B.n762 585
R1037 B.n764 B.n763 585
R1038 B.n760 B.n325 585
R1039 B.n325 B.n324 585
R1040 B.n759 B.n758 585
R1041 B.n758 B.n757 585
R1042 B.n327 B.n326 585
R1043 B.n328 B.n327 585
R1044 B.n750 B.n749 585
R1045 B.n751 B.n750 585
R1046 B.n748 B.n333 585
R1047 B.n333 B.n332 585
R1048 B.n747 B.n746 585
R1049 B.n746 B.n745 585
R1050 B.n335 B.n334 585
R1051 B.n336 B.n335 585
R1052 B.n738 B.n737 585
R1053 B.n739 B.n738 585
R1054 B.n736 B.n341 585
R1055 B.n341 B.n340 585
R1056 B.n735 B.n734 585
R1057 B.n734 B.n733 585
R1058 B.n343 B.n342 585
R1059 B.n344 B.n343 585
R1060 B.n726 B.n725 585
R1061 B.n727 B.n726 585
R1062 B.n724 B.n349 585
R1063 B.n349 B.n348 585
R1064 B.n723 B.n722 585
R1065 B.n722 B.n721 585
R1066 B.n351 B.n350 585
R1067 B.n352 B.n351 585
R1068 B.n714 B.n713 585
R1069 B.n715 B.n714 585
R1070 B.n712 B.n357 585
R1071 B.n357 B.n356 585
R1072 B.n711 B.n710 585
R1073 B.n710 B.n709 585
R1074 B.n359 B.n358 585
R1075 B.n360 B.n359 585
R1076 B.n702 B.n701 585
R1077 B.n703 B.n702 585
R1078 B.n700 B.n365 585
R1079 B.n365 B.n364 585
R1080 B.n699 B.n698 585
R1081 B.n698 B.n697 585
R1082 B.n367 B.n366 585
R1083 B.n368 B.n367 585
R1084 B.n690 B.n689 585
R1085 B.n691 B.n690 585
R1086 B.n688 B.n373 585
R1087 B.n373 B.n372 585
R1088 B.n687 B.n686 585
R1089 B.n686 B.n685 585
R1090 B.n375 B.n374 585
R1091 B.n376 B.n375 585
R1092 B.n678 B.n677 585
R1093 B.n679 B.n678 585
R1094 B.n676 B.n381 585
R1095 B.n381 B.n380 585
R1096 B.n675 B.n674 585
R1097 B.n674 B.n673 585
R1098 B.n383 B.n382 585
R1099 B.n666 B.n383 585
R1100 B.n665 B.n664 585
R1101 B.n667 B.n665 585
R1102 B.n663 B.n388 585
R1103 B.n388 B.n387 585
R1104 B.n662 B.n661 585
R1105 B.n661 B.n660 585
R1106 B.n390 B.n389 585
R1107 B.n391 B.n390 585
R1108 B.n653 B.n652 585
R1109 B.n654 B.n653 585
R1110 B.n651 B.n396 585
R1111 B.n396 B.n395 585
R1112 B.n650 B.n649 585
R1113 B.n649 B.n648 585
R1114 B.n398 B.n397 585
R1115 B.n399 B.n398 585
R1116 B.n641 B.n640 585
R1117 B.n642 B.n641 585
R1118 B.n402 B.n401 585
R1119 B.n455 B.n453 585
R1120 B.n456 B.n452 585
R1121 B.n456 B.n403 585
R1122 B.n459 B.n458 585
R1123 B.n460 B.n451 585
R1124 B.n462 B.n461 585
R1125 B.n464 B.n450 585
R1126 B.n467 B.n466 585
R1127 B.n468 B.n449 585
R1128 B.n470 B.n469 585
R1129 B.n472 B.n448 585
R1130 B.n475 B.n474 585
R1131 B.n476 B.n447 585
R1132 B.n478 B.n477 585
R1133 B.n480 B.n446 585
R1134 B.n483 B.n482 585
R1135 B.n484 B.n445 585
R1136 B.n486 B.n485 585
R1137 B.n488 B.n444 585
R1138 B.n491 B.n490 585
R1139 B.n492 B.n443 585
R1140 B.n494 B.n493 585
R1141 B.n496 B.n442 585
R1142 B.n499 B.n498 585
R1143 B.n500 B.n441 585
R1144 B.n502 B.n501 585
R1145 B.n504 B.n440 585
R1146 B.n507 B.n506 585
R1147 B.n508 B.n439 585
R1148 B.n510 B.n509 585
R1149 B.n512 B.n438 585
R1150 B.n515 B.n514 585
R1151 B.n516 B.n437 585
R1152 B.n518 B.n517 585
R1153 B.n520 B.n436 585
R1154 B.n523 B.n522 585
R1155 B.n524 B.n435 585
R1156 B.n526 B.n525 585
R1157 B.n528 B.n434 585
R1158 B.n531 B.n530 585
R1159 B.n532 B.n433 585
R1160 B.n537 B.n536 585
R1161 B.n539 B.n432 585
R1162 B.n542 B.n541 585
R1163 B.n543 B.n431 585
R1164 B.n545 B.n544 585
R1165 B.n547 B.n430 585
R1166 B.n550 B.n549 585
R1167 B.n551 B.n429 585
R1168 B.n553 B.n552 585
R1169 B.n555 B.n428 585
R1170 B.n558 B.n557 585
R1171 B.n559 B.n424 585
R1172 B.n561 B.n560 585
R1173 B.n563 B.n423 585
R1174 B.n566 B.n565 585
R1175 B.n567 B.n422 585
R1176 B.n569 B.n568 585
R1177 B.n571 B.n421 585
R1178 B.n574 B.n573 585
R1179 B.n575 B.n420 585
R1180 B.n577 B.n576 585
R1181 B.n579 B.n419 585
R1182 B.n582 B.n581 585
R1183 B.n583 B.n418 585
R1184 B.n585 B.n584 585
R1185 B.n587 B.n417 585
R1186 B.n590 B.n589 585
R1187 B.n591 B.n416 585
R1188 B.n593 B.n592 585
R1189 B.n595 B.n415 585
R1190 B.n598 B.n597 585
R1191 B.n599 B.n414 585
R1192 B.n601 B.n600 585
R1193 B.n603 B.n413 585
R1194 B.n606 B.n605 585
R1195 B.n607 B.n412 585
R1196 B.n609 B.n608 585
R1197 B.n611 B.n411 585
R1198 B.n614 B.n613 585
R1199 B.n615 B.n410 585
R1200 B.n617 B.n616 585
R1201 B.n619 B.n409 585
R1202 B.n622 B.n621 585
R1203 B.n623 B.n408 585
R1204 B.n625 B.n624 585
R1205 B.n627 B.n407 585
R1206 B.n630 B.n629 585
R1207 B.n631 B.n406 585
R1208 B.n633 B.n632 585
R1209 B.n635 B.n405 585
R1210 B.n638 B.n637 585
R1211 B.n639 B.n404 585
R1212 B.n644 B.n643 585
R1213 B.n643 B.n642 585
R1214 B.n645 B.n400 585
R1215 B.n400 B.n399 585
R1216 B.n647 B.n646 585
R1217 B.n648 B.n647 585
R1218 B.n394 B.n393 585
R1219 B.n395 B.n394 585
R1220 B.n656 B.n655 585
R1221 B.n655 B.n654 585
R1222 B.n657 B.n392 585
R1223 B.n392 B.n391 585
R1224 B.n659 B.n658 585
R1225 B.n660 B.n659 585
R1226 B.n386 B.n385 585
R1227 B.n387 B.n386 585
R1228 B.n669 B.n668 585
R1229 B.n668 B.n667 585
R1230 B.n670 B.n384 585
R1231 B.n666 B.n384 585
R1232 B.n672 B.n671 585
R1233 B.n673 B.n672 585
R1234 B.n379 B.n378 585
R1235 B.n380 B.n379 585
R1236 B.n681 B.n680 585
R1237 B.n680 B.n679 585
R1238 B.n682 B.n377 585
R1239 B.n377 B.n376 585
R1240 B.n684 B.n683 585
R1241 B.n685 B.n684 585
R1242 B.n371 B.n370 585
R1243 B.n372 B.n371 585
R1244 B.n693 B.n692 585
R1245 B.n692 B.n691 585
R1246 B.n694 B.n369 585
R1247 B.n369 B.n368 585
R1248 B.n696 B.n695 585
R1249 B.n697 B.n696 585
R1250 B.n363 B.n362 585
R1251 B.n364 B.n363 585
R1252 B.n705 B.n704 585
R1253 B.n704 B.n703 585
R1254 B.n706 B.n361 585
R1255 B.n361 B.n360 585
R1256 B.n708 B.n707 585
R1257 B.n709 B.n708 585
R1258 B.n355 B.n354 585
R1259 B.n356 B.n355 585
R1260 B.n717 B.n716 585
R1261 B.n716 B.n715 585
R1262 B.n718 B.n353 585
R1263 B.n353 B.n352 585
R1264 B.n720 B.n719 585
R1265 B.n721 B.n720 585
R1266 B.n347 B.n346 585
R1267 B.n348 B.n347 585
R1268 B.n729 B.n728 585
R1269 B.n728 B.n727 585
R1270 B.n730 B.n345 585
R1271 B.n345 B.n344 585
R1272 B.n732 B.n731 585
R1273 B.n733 B.n732 585
R1274 B.n339 B.n338 585
R1275 B.n340 B.n339 585
R1276 B.n741 B.n740 585
R1277 B.n740 B.n739 585
R1278 B.n742 B.n337 585
R1279 B.n337 B.n336 585
R1280 B.n744 B.n743 585
R1281 B.n745 B.n744 585
R1282 B.n331 B.n330 585
R1283 B.n332 B.n331 585
R1284 B.n753 B.n752 585
R1285 B.n752 B.n751 585
R1286 B.n754 B.n329 585
R1287 B.n329 B.n328 585
R1288 B.n756 B.n755 585
R1289 B.n757 B.n756 585
R1290 B.n323 B.n322 585
R1291 B.n324 B.n323 585
R1292 B.n766 B.n765 585
R1293 B.n765 B.n764 585
R1294 B.n767 B.n321 585
R1295 B.n321 B.n320 585
R1296 B.n769 B.n768 585
R1297 B.n770 B.n769 585
R1298 B.n3 B.n0 585
R1299 B.n4 B.n3 585
R1300 B.n921 B.n1 585
R1301 B.n922 B.n921 585
R1302 B.n920 B.n919 585
R1303 B.n920 B.n8 585
R1304 B.n918 B.n9 585
R1305 B.n12 B.n9 585
R1306 B.n917 B.n916 585
R1307 B.n916 B.n915 585
R1308 B.n11 B.n10 585
R1309 B.n914 B.n11 585
R1310 B.n912 B.n911 585
R1311 B.n913 B.n912 585
R1312 B.n910 B.n17 585
R1313 B.n17 B.n16 585
R1314 B.n909 B.n908 585
R1315 B.n908 B.n907 585
R1316 B.n19 B.n18 585
R1317 B.n906 B.n19 585
R1318 B.n904 B.n903 585
R1319 B.n905 B.n904 585
R1320 B.n902 B.n24 585
R1321 B.n24 B.n23 585
R1322 B.n901 B.n900 585
R1323 B.n900 B.n899 585
R1324 B.n26 B.n25 585
R1325 B.n898 B.n26 585
R1326 B.n896 B.n895 585
R1327 B.n897 B.n896 585
R1328 B.n894 B.n31 585
R1329 B.n31 B.n30 585
R1330 B.n893 B.n892 585
R1331 B.n892 B.n891 585
R1332 B.n33 B.n32 585
R1333 B.n890 B.n33 585
R1334 B.n888 B.n887 585
R1335 B.n889 B.n888 585
R1336 B.n886 B.n38 585
R1337 B.n38 B.n37 585
R1338 B.n885 B.n884 585
R1339 B.n884 B.n883 585
R1340 B.n40 B.n39 585
R1341 B.n882 B.n40 585
R1342 B.n880 B.n879 585
R1343 B.n881 B.n880 585
R1344 B.n878 B.n45 585
R1345 B.n45 B.n44 585
R1346 B.n877 B.n876 585
R1347 B.n876 B.n875 585
R1348 B.n47 B.n46 585
R1349 B.n874 B.n47 585
R1350 B.n872 B.n871 585
R1351 B.n873 B.n872 585
R1352 B.n870 B.n52 585
R1353 B.n52 B.n51 585
R1354 B.n869 B.n868 585
R1355 B.n868 B.n867 585
R1356 B.n54 B.n53 585
R1357 B.n866 B.n54 585
R1358 B.n864 B.n863 585
R1359 B.n865 B.n864 585
R1360 B.n862 B.n59 585
R1361 B.n59 B.n58 585
R1362 B.n861 B.n860 585
R1363 B.n860 B.n859 585
R1364 B.n61 B.n60 585
R1365 B.n858 B.n61 585
R1366 B.n856 B.n855 585
R1367 B.n857 B.n856 585
R1368 B.n854 B.n65 585
R1369 B.n68 B.n65 585
R1370 B.n853 B.n852 585
R1371 B.n852 B.n851 585
R1372 B.n67 B.n66 585
R1373 B.n850 B.n67 585
R1374 B.n848 B.n847 585
R1375 B.n849 B.n848 585
R1376 B.n846 B.n73 585
R1377 B.n73 B.n72 585
R1378 B.n845 B.n844 585
R1379 B.n844 B.n843 585
R1380 B.n75 B.n74 585
R1381 B.n842 B.n75 585
R1382 B.n840 B.n839 585
R1383 B.n841 B.n840 585
R1384 B.n838 B.n80 585
R1385 B.n80 B.n79 585
R1386 B.n837 B.n836 585
R1387 B.n836 B.n835 585
R1388 B.n925 B.n924 585
R1389 B.n923 B.n2 585
R1390 B.n836 B.n82 545.355
R1391 B.n833 B.n83 545.355
R1392 B.n641 B.n404 545.355
R1393 B.n643 B.n402 545.355
R1394 B.n133 B.t9 364.238
R1395 B.n131 B.t6 364.238
R1396 B.n425 B.t17 364.238
R1397 B.n533 B.t14 364.238
R1398 B.n133 B.t8 286.147
R1399 B.n131 B.t4 286.147
R1400 B.n425 B.t15 286.147
R1401 B.n533 B.t11 286.147
R1402 B.n132 B.t7 284.142
R1403 B.n426 B.t16 284.142
R1404 B.n134 B.t10 284.142
R1405 B.n534 B.t13 284.142
R1406 B.n834 B.n129 256.663
R1407 B.n834 B.n128 256.663
R1408 B.n834 B.n127 256.663
R1409 B.n834 B.n126 256.663
R1410 B.n834 B.n125 256.663
R1411 B.n834 B.n124 256.663
R1412 B.n834 B.n123 256.663
R1413 B.n834 B.n122 256.663
R1414 B.n834 B.n121 256.663
R1415 B.n834 B.n120 256.663
R1416 B.n834 B.n119 256.663
R1417 B.n834 B.n118 256.663
R1418 B.n834 B.n117 256.663
R1419 B.n834 B.n116 256.663
R1420 B.n834 B.n115 256.663
R1421 B.n834 B.n114 256.663
R1422 B.n834 B.n113 256.663
R1423 B.n834 B.n112 256.663
R1424 B.n834 B.n111 256.663
R1425 B.n834 B.n110 256.663
R1426 B.n834 B.n109 256.663
R1427 B.n834 B.n108 256.663
R1428 B.n834 B.n107 256.663
R1429 B.n834 B.n106 256.663
R1430 B.n834 B.n105 256.663
R1431 B.n834 B.n104 256.663
R1432 B.n834 B.n103 256.663
R1433 B.n834 B.n102 256.663
R1434 B.n834 B.n101 256.663
R1435 B.n834 B.n100 256.663
R1436 B.n834 B.n99 256.663
R1437 B.n834 B.n98 256.663
R1438 B.n834 B.n97 256.663
R1439 B.n834 B.n96 256.663
R1440 B.n834 B.n95 256.663
R1441 B.n834 B.n94 256.663
R1442 B.n834 B.n93 256.663
R1443 B.n834 B.n92 256.663
R1444 B.n834 B.n91 256.663
R1445 B.n834 B.n90 256.663
R1446 B.n834 B.n89 256.663
R1447 B.n834 B.n88 256.663
R1448 B.n834 B.n87 256.663
R1449 B.n834 B.n86 256.663
R1450 B.n834 B.n85 256.663
R1451 B.n834 B.n84 256.663
R1452 B.n454 B.n403 256.663
R1453 B.n457 B.n403 256.663
R1454 B.n463 B.n403 256.663
R1455 B.n465 B.n403 256.663
R1456 B.n471 B.n403 256.663
R1457 B.n473 B.n403 256.663
R1458 B.n479 B.n403 256.663
R1459 B.n481 B.n403 256.663
R1460 B.n487 B.n403 256.663
R1461 B.n489 B.n403 256.663
R1462 B.n495 B.n403 256.663
R1463 B.n497 B.n403 256.663
R1464 B.n503 B.n403 256.663
R1465 B.n505 B.n403 256.663
R1466 B.n511 B.n403 256.663
R1467 B.n513 B.n403 256.663
R1468 B.n519 B.n403 256.663
R1469 B.n521 B.n403 256.663
R1470 B.n527 B.n403 256.663
R1471 B.n529 B.n403 256.663
R1472 B.n538 B.n403 256.663
R1473 B.n540 B.n403 256.663
R1474 B.n546 B.n403 256.663
R1475 B.n548 B.n403 256.663
R1476 B.n554 B.n403 256.663
R1477 B.n556 B.n403 256.663
R1478 B.n562 B.n403 256.663
R1479 B.n564 B.n403 256.663
R1480 B.n570 B.n403 256.663
R1481 B.n572 B.n403 256.663
R1482 B.n578 B.n403 256.663
R1483 B.n580 B.n403 256.663
R1484 B.n586 B.n403 256.663
R1485 B.n588 B.n403 256.663
R1486 B.n594 B.n403 256.663
R1487 B.n596 B.n403 256.663
R1488 B.n602 B.n403 256.663
R1489 B.n604 B.n403 256.663
R1490 B.n610 B.n403 256.663
R1491 B.n612 B.n403 256.663
R1492 B.n618 B.n403 256.663
R1493 B.n620 B.n403 256.663
R1494 B.n626 B.n403 256.663
R1495 B.n628 B.n403 256.663
R1496 B.n634 B.n403 256.663
R1497 B.n636 B.n403 256.663
R1498 B.n927 B.n926 256.663
R1499 B.n138 B.n137 163.367
R1500 B.n142 B.n141 163.367
R1501 B.n146 B.n145 163.367
R1502 B.n150 B.n149 163.367
R1503 B.n154 B.n153 163.367
R1504 B.n158 B.n157 163.367
R1505 B.n162 B.n161 163.367
R1506 B.n166 B.n165 163.367
R1507 B.n170 B.n169 163.367
R1508 B.n174 B.n173 163.367
R1509 B.n178 B.n177 163.367
R1510 B.n182 B.n181 163.367
R1511 B.n186 B.n185 163.367
R1512 B.n190 B.n189 163.367
R1513 B.n194 B.n193 163.367
R1514 B.n198 B.n197 163.367
R1515 B.n202 B.n201 163.367
R1516 B.n206 B.n205 163.367
R1517 B.n210 B.n209 163.367
R1518 B.n214 B.n213 163.367
R1519 B.n218 B.n217 163.367
R1520 B.n222 B.n221 163.367
R1521 B.n226 B.n225 163.367
R1522 B.n230 B.n229 163.367
R1523 B.n234 B.n233 163.367
R1524 B.n239 B.n238 163.367
R1525 B.n243 B.n242 163.367
R1526 B.n247 B.n246 163.367
R1527 B.n251 B.n250 163.367
R1528 B.n255 B.n254 163.367
R1529 B.n259 B.n258 163.367
R1530 B.n263 B.n262 163.367
R1531 B.n267 B.n266 163.367
R1532 B.n271 B.n270 163.367
R1533 B.n275 B.n274 163.367
R1534 B.n279 B.n278 163.367
R1535 B.n283 B.n282 163.367
R1536 B.n287 B.n286 163.367
R1537 B.n291 B.n290 163.367
R1538 B.n295 B.n294 163.367
R1539 B.n299 B.n298 163.367
R1540 B.n303 B.n302 163.367
R1541 B.n307 B.n306 163.367
R1542 B.n311 B.n310 163.367
R1543 B.n315 B.n314 163.367
R1544 B.n833 B.n130 163.367
R1545 B.n641 B.n398 163.367
R1546 B.n649 B.n398 163.367
R1547 B.n649 B.n396 163.367
R1548 B.n653 B.n396 163.367
R1549 B.n653 B.n390 163.367
R1550 B.n661 B.n390 163.367
R1551 B.n661 B.n388 163.367
R1552 B.n665 B.n388 163.367
R1553 B.n665 B.n383 163.367
R1554 B.n674 B.n383 163.367
R1555 B.n674 B.n381 163.367
R1556 B.n678 B.n381 163.367
R1557 B.n678 B.n375 163.367
R1558 B.n686 B.n375 163.367
R1559 B.n686 B.n373 163.367
R1560 B.n690 B.n373 163.367
R1561 B.n690 B.n367 163.367
R1562 B.n698 B.n367 163.367
R1563 B.n698 B.n365 163.367
R1564 B.n702 B.n365 163.367
R1565 B.n702 B.n359 163.367
R1566 B.n710 B.n359 163.367
R1567 B.n710 B.n357 163.367
R1568 B.n714 B.n357 163.367
R1569 B.n714 B.n351 163.367
R1570 B.n722 B.n351 163.367
R1571 B.n722 B.n349 163.367
R1572 B.n726 B.n349 163.367
R1573 B.n726 B.n343 163.367
R1574 B.n734 B.n343 163.367
R1575 B.n734 B.n341 163.367
R1576 B.n738 B.n341 163.367
R1577 B.n738 B.n335 163.367
R1578 B.n746 B.n335 163.367
R1579 B.n746 B.n333 163.367
R1580 B.n750 B.n333 163.367
R1581 B.n750 B.n327 163.367
R1582 B.n758 B.n327 163.367
R1583 B.n758 B.n325 163.367
R1584 B.n763 B.n325 163.367
R1585 B.n763 B.n319 163.367
R1586 B.n771 B.n319 163.367
R1587 B.n772 B.n771 163.367
R1588 B.n772 B.n5 163.367
R1589 B.n6 B.n5 163.367
R1590 B.n7 B.n6 163.367
R1591 B.n778 B.n7 163.367
R1592 B.n779 B.n778 163.367
R1593 B.n779 B.n13 163.367
R1594 B.n14 B.n13 163.367
R1595 B.n15 B.n14 163.367
R1596 B.n784 B.n15 163.367
R1597 B.n784 B.n20 163.367
R1598 B.n21 B.n20 163.367
R1599 B.n22 B.n21 163.367
R1600 B.n789 B.n22 163.367
R1601 B.n789 B.n27 163.367
R1602 B.n28 B.n27 163.367
R1603 B.n29 B.n28 163.367
R1604 B.n794 B.n29 163.367
R1605 B.n794 B.n34 163.367
R1606 B.n35 B.n34 163.367
R1607 B.n36 B.n35 163.367
R1608 B.n799 B.n36 163.367
R1609 B.n799 B.n41 163.367
R1610 B.n42 B.n41 163.367
R1611 B.n43 B.n42 163.367
R1612 B.n804 B.n43 163.367
R1613 B.n804 B.n48 163.367
R1614 B.n49 B.n48 163.367
R1615 B.n50 B.n49 163.367
R1616 B.n809 B.n50 163.367
R1617 B.n809 B.n55 163.367
R1618 B.n56 B.n55 163.367
R1619 B.n57 B.n56 163.367
R1620 B.n814 B.n57 163.367
R1621 B.n814 B.n62 163.367
R1622 B.n63 B.n62 163.367
R1623 B.n64 B.n63 163.367
R1624 B.n819 B.n64 163.367
R1625 B.n819 B.n69 163.367
R1626 B.n70 B.n69 163.367
R1627 B.n71 B.n70 163.367
R1628 B.n824 B.n71 163.367
R1629 B.n824 B.n76 163.367
R1630 B.n77 B.n76 163.367
R1631 B.n78 B.n77 163.367
R1632 B.n829 B.n78 163.367
R1633 B.n829 B.n83 163.367
R1634 B.n456 B.n455 163.367
R1635 B.n458 B.n456 163.367
R1636 B.n462 B.n451 163.367
R1637 B.n466 B.n464 163.367
R1638 B.n470 B.n449 163.367
R1639 B.n474 B.n472 163.367
R1640 B.n478 B.n447 163.367
R1641 B.n482 B.n480 163.367
R1642 B.n486 B.n445 163.367
R1643 B.n490 B.n488 163.367
R1644 B.n494 B.n443 163.367
R1645 B.n498 B.n496 163.367
R1646 B.n502 B.n441 163.367
R1647 B.n506 B.n504 163.367
R1648 B.n510 B.n439 163.367
R1649 B.n514 B.n512 163.367
R1650 B.n518 B.n437 163.367
R1651 B.n522 B.n520 163.367
R1652 B.n526 B.n435 163.367
R1653 B.n530 B.n528 163.367
R1654 B.n537 B.n433 163.367
R1655 B.n541 B.n539 163.367
R1656 B.n545 B.n431 163.367
R1657 B.n549 B.n547 163.367
R1658 B.n553 B.n429 163.367
R1659 B.n557 B.n555 163.367
R1660 B.n561 B.n424 163.367
R1661 B.n565 B.n563 163.367
R1662 B.n569 B.n422 163.367
R1663 B.n573 B.n571 163.367
R1664 B.n577 B.n420 163.367
R1665 B.n581 B.n579 163.367
R1666 B.n585 B.n418 163.367
R1667 B.n589 B.n587 163.367
R1668 B.n593 B.n416 163.367
R1669 B.n597 B.n595 163.367
R1670 B.n601 B.n414 163.367
R1671 B.n605 B.n603 163.367
R1672 B.n609 B.n412 163.367
R1673 B.n613 B.n611 163.367
R1674 B.n617 B.n410 163.367
R1675 B.n621 B.n619 163.367
R1676 B.n625 B.n408 163.367
R1677 B.n629 B.n627 163.367
R1678 B.n633 B.n406 163.367
R1679 B.n637 B.n635 163.367
R1680 B.n643 B.n400 163.367
R1681 B.n647 B.n400 163.367
R1682 B.n647 B.n394 163.367
R1683 B.n655 B.n394 163.367
R1684 B.n655 B.n392 163.367
R1685 B.n659 B.n392 163.367
R1686 B.n659 B.n386 163.367
R1687 B.n668 B.n386 163.367
R1688 B.n668 B.n384 163.367
R1689 B.n672 B.n384 163.367
R1690 B.n672 B.n379 163.367
R1691 B.n680 B.n379 163.367
R1692 B.n680 B.n377 163.367
R1693 B.n684 B.n377 163.367
R1694 B.n684 B.n371 163.367
R1695 B.n692 B.n371 163.367
R1696 B.n692 B.n369 163.367
R1697 B.n696 B.n369 163.367
R1698 B.n696 B.n363 163.367
R1699 B.n704 B.n363 163.367
R1700 B.n704 B.n361 163.367
R1701 B.n708 B.n361 163.367
R1702 B.n708 B.n355 163.367
R1703 B.n716 B.n355 163.367
R1704 B.n716 B.n353 163.367
R1705 B.n720 B.n353 163.367
R1706 B.n720 B.n347 163.367
R1707 B.n728 B.n347 163.367
R1708 B.n728 B.n345 163.367
R1709 B.n732 B.n345 163.367
R1710 B.n732 B.n339 163.367
R1711 B.n740 B.n339 163.367
R1712 B.n740 B.n337 163.367
R1713 B.n744 B.n337 163.367
R1714 B.n744 B.n331 163.367
R1715 B.n752 B.n331 163.367
R1716 B.n752 B.n329 163.367
R1717 B.n756 B.n329 163.367
R1718 B.n756 B.n323 163.367
R1719 B.n765 B.n323 163.367
R1720 B.n765 B.n321 163.367
R1721 B.n769 B.n321 163.367
R1722 B.n769 B.n3 163.367
R1723 B.n925 B.n3 163.367
R1724 B.n921 B.n2 163.367
R1725 B.n921 B.n920 163.367
R1726 B.n920 B.n9 163.367
R1727 B.n916 B.n9 163.367
R1728 B.n916 B.n11 163.367
R1729 B.n912 B.n11 163.367
R1730 B.n912 B.n17 163.367
R1731 B.n908 B.n17 163.367
R1732 B.n908 B.n19 163.367
R1733 B.n904 B.n19 163.367
R1734 B.n904 B.n24 163.367
R1735 B.n900 B.n24 163.367
R1736 B.n900 B.n26 163.367
R1737 B.n896 B.n26 163.367
R1738 B.n896 B.n31 163.367
R1739 B.n892 B.n31 163.367
R1740 B.n892 B.n33 163.367
R1741 B.n888 B.n33 163.367
R1742 B.n888 B.n38 163.367
R1743 B.n884 B.n38 163.367
R1744 B.n884 B.n40 163.367
R1745 B.n880 B.n40 163.367
R1746 B.n880 B.n45 163.367
R1747 B.n876 B.n45 163.367
R1748 B.n876 B.n47 163.367
R1749 B.n872 B.n47 163.367
R1750 B.n872 B.n52 163.367
R1751 B.n868 B.n52 163.367
R1752 B.n868 B.n54 163.367
R1753 B.n864 B.n54 163.367
R1754 B.n864 B.n59 163.367
R1755 B.n860 B.n59 163.367
R1756 B.n860 B.n61 163.367
R1757 B.n856 B.n61 163.367
R1758 B.n856 B.n65 163.367
R1759 B.n852 B.n65 163.367
R1760 B.n852 B.n67 163.367
R1761 B.n848 B.n67 163.367
R1762 B.n848 B.n73 163.367
R1763 B.n844 B.n73 163.367
R1764 B.n844 B.n75 163.367
R1765 B.n840 B.n75 163.367
R1766 B.n840 B.n80 163.367
R1767 B.n836 B.n80 163.367
R1768 B.n642 B.n403 80.3571
R1769 B.n835 B.n834 80.3571
R1770 B.n134 B.n133 80.0975
R1771 B.n132 B.n131 80.0975
R1772 B.n426 B.n425 80.0975
R1773 B.n534 B.n533 80.0975
R1774 B.n84 B.n82 71.676
R1775 B.n138 B.n85 71.676
R1776 B.n142 B.n86 71.676
R1777 B.n146 B.n87 71.676
R1778 B.n150 B.n88 71.676
R1779 B.n154 B.n89 71.676
R1780 B.n158 B.n90 71.676
R1781 B.n162 B.n91 71.676
R1782 B.n166 B.n92 71.676
R1783 B.n170 B.n93 71.676
R1784 B.n174 B.n94 71.676
R1785 B.n178 B.n95 71.676
R1786 B.n182 B.n96 71.676
R1787 B.n186 B.n97 71.676
R1788 B.n190 B.n98 71.676
R1789 B.n194 B.n99 71.676
R1790 B.n198 B.n100 71.676
R1791 B.n202 B.n101 71.676
R1792 B.n206 B.n102 71.676
R1793 B.n210 B.n103 71.676
R1794 B.n214 B.n104 71.676
R1795 B.n218 B.n105 71.676
R1796 B.n222 B.n106 71.676
R1797 B.n226 B.n107 71.676
R1798 B.n230 B.n108 71.676
R1799 B.n234 B.n109 71.676
R1800 B.n239 B.n110 71.676
R1801 B.n243 B.n111 71.676
R1802 B.n247 B.n112 71.676
R1803 B.n251 B.n113 71.676
R1804 B.n255 B.n114 71.676
R1805 B.n259 B.n115 71.676
R1806 B.n263 B.n116 71.676
R1807 B.n267 B.n117 71.676
R1808 B.n271 B.n118 71.676
R1809 B.n275 B.n119 71.676
R1810 B.n279 B.n120 71.676
R1811 B.n283 B.n121 71.676
R1812 B.n287 B.n122 71.676
R1813 B.n291 B.n123 71.676
R1814 B.n295 B.n124 71.676
R1815 B.n299 B.n125 71.676
R1816 B.n303 B.n126 71.676
R1817 B.n307 B.n127 71.676
R1818 B.n311 B.n128 71.676
R1819 B.n315 B.n129 71.676
R1820 B.n130 B.n129 71.676
R1821 B.n314 B.n128 71.676
R1822 B.n310 B.n127 71.676
R1823 B.n306 B.n126 71.676
R1824 B.n302 B.n125 71.676
R1825 B.n298 B.n124 71.676
R1826 B.n294 B.n123 71.676
R1827 B.n290 B.n122 71.676
R1828 B.n286 B.n121 71.676
R1829 B.n282 B.n120 71.676
R1830 B.n278 B.n119 71.676
R1831 B.n274 B.n118 71.676
R1832 B.n270 B.n117 71.676
R1833 B.n266 B.n116 71.676
R1834 B.n262 B.n115 71.676
R1835 B.n258 B.n114 71.676
R1836 B.n254 B.n113 71.676
R1837 B.n250 B.n112 71.676
R1838 B.n246 B.n111 71.676
R1839 B.n242 B.n110 71.676
R1840 B.n238 B.n109 71.676
R1841 B.n233 B.n108 71.676
R1842 B.n229 B.n107 71.676
R1843 B.n225 B.n106 71.676
R1844 B.n221 B.n105 71.676
R1845 B.n217 B.n104 71.676
R1846 B.n213 B.n103 71.676
R1847 B.n209 B.n102 71.676
R1848 B.n205 B.n101 71.676
R1849 B.n201 B.n100 71.676
R1850 B.n197 B.n99 71.676
R1851 B.n193 B.n98 71.676
R1852 B.n189 B.n97 71.676
R1853 B.n185 B.n96 71.676
R1854 B.n181 B.n95 71.676
R1855 B.n177 B.n94 71.676
R1856 B.n173 B.n93 71.676
R1857 B.n169 B.n92 71.676
R1858 B.n165 B.n91 71.676
R1859 B.n161 B.n90 71.676
R1860 B.n157 B.n89 71.676
R1861 B.n153 B.n88 71.676
R1862 B.n149 B.n87 71.676
R1863 B.n145 B.n86 71.676
R1864 B.n141 B.n85 71.676
R1865 B.n137 B.n84 71.676
R1866 B.n454 B.n402 71.676
R1867 B.n458 B.n457 71.676
R1868 B.n463 B.n462 71.676
R1869 B.n466 B.n465 71.676
R1870 B.n471 B.n470 71.676
R1871 B.n474 B.n473 71.676
R1872 B.n479 B.n478 71.676
R1873 B.n482 B.n481 71.676
R1874 B.n487 B.n486 71.676
R1875 B.n490 B.n489 71.676
R1876 B.n495 B.n494 71.676
R1877 B.n498 B.n497 71.676
R1878 B.n503 B.n502 71.676
R1879 B.n506 B.n505 71.676
R1880 B.n511 B.n510 71.676
R1881 B.n514 B.n513 71.676
R1882 B.n519 B.n518 71.676
R1883 B.n522 B.n521 71.676
R1884 B.n527 B.n526 71.676
R1885 B.n530 B.n529 71.676
R1886 B.n538 B.n537 71.676
R1887 B.n541 B.n540 71.676
R1888 B.n546 B.n545 71.676
R1889 B.n549 B.n548 71.676
R1890 B.n554 B.n553 71.676
R1891 B.n557 B.n556 71.676
R1892 B.n562 B.n561 71.676
R1893 B.n565 B.n564 71.676
R1894 B.n570 B.n569 71.676
R1895 B.n573 B.n572 71.676
R1896 B.n578 B.n577 71.676
R1897 B.n581 B.n580 71.676
R1898 B.n586 B.n585 71.676
R1899 B.n589 B.n588 71.676
R1900 B.n594 B.n593 71.676
R1901 B.n597 B.n596 71.676
R1902 B.n602 B.n601 71.676
R1903 B.n605 B.n604 71.676
R1904 B.n610 B.n609 71.676
R1905 B.n613 B.n612 71.676
R1906 B.n618 B.n617 71.676
R1907 B.n621 B.n620 71.676
R1908 B.n626 B.n625 71.676
R1909 B.n629 B.n628 71.676
R1910 B.n634 B.n633 71.676
R1911 B.n637 B.n636 71.676
R1912 B.n455 B.n454 71.676
R1913 B.n457 B.n451 71.676
R1914 B.n464 B.n463 71.676
R1915 B.n465 B.n449 71.676
R1916 B.n472 B.n471 71.676
R1917 B.n473 B.n447 71.676
R1918 B.n480 B.n479 71.676
R1919 B.n481 B.n445 71.676
R1920 B.n488 B.n487 71.676
R1921 B.n489 B.n443 71.676
R1922 B.n496 B.n495 71.676
R1923 B.n497 B.n441 71.676
R1924 B.n504 B.n503 71.676
R1925 B.n505 B.n439 71.676
R1926 B.n512 B.n511 71.676
R1927 B.n513 B.n437 71.676
R1928 B.n520 B.n519 71.676
R1929 B.n521 B.n435 71.676
R1930 B.n528 B.n527 71.676
R1931 B.n529 B.n433 71.676
R1932 B.n539 B.n538 71.676
R1933 B.n540 B.n431 71.676
R1934 B.n547 B.n546 71.676
R1935 B.n548 B.n429 71.676
R1936 B.n555 B.n554 71.676
R1937 B.n556 B.n424 71.676
R1938 B.n563 B.n562 71.676
R1939 B.n564 B.n422 71.676
R1940 B.n571 B.n570 71.676
R1941 B.n572 B.n420 71.676
R1942 B.n579 B.n578 71.676
R1943 B.n580 B.n418 71.676
R1944 B.n587 B.n586 71.676
R1945 B.n588 B.n416 71.676
R1946 B.n595 B.n594 71.676
R1947 B.n596 B.n414 71.676
R1948 B.n603 B.n602 71.676
R1949 B.n604 B.n412 71.676
R1950 B.n611 B.n610 71.676
R1951 B.n612 B.n410 71.676
R1952 B.n619 B.n618 71.676
R1953 B.n620 B.n408 71.676
R1954 B.n627 B.n626 71.676
R1955 B.n628 B.n406 71.676
R1956 B.n635 B.n634 71.676
R1957 B.n636 B.n404 71.676
R1958 B.n926 B.n925 71.676
R1959 B.n926 B.n2 71.676
R1960 B.n135 B.n134 59.5399
R1961 B.n236 B.n132 59.5399
R1962 B.n427 B.n426 59.5399
R1963 B.n535 B.n534 59.5399
R1964 B.n642 B.n399 43.0261
R1965 B.n648 B.n399 43.0261
R1966 B.n648 B.n395 43.0261
R1967 B.n654 B.n395 43.0261
R1968 B.n654 B.n391 43.0261
R1969 B.n660 B.n391 43.0261
R1970 B.n660 B.n387 43.0261
R1971 B.n667 B.n387 43.0261
R1972 B.n667 B.n666 43.0261
R1973 B.n673 B.n380 43.0261
R1974 B.n679 B.n380 43.0261
R1975 B.n679 B.n376 43.0261
R1976 B.n685 B.n376 43.0261
R1977 B.n685 B.n372 43.0261
R1978 B.n691 B.n372 43.0261
R1979 B.n691 B.n368 43.0261
R1980 B.n697 B.n368 43.0261
R1981 B.n697 B.n364 43.0261
R1982 B.n703 B.n364 43.0261
R1983 B.n703 B.n360 43.0261
R1984 B.n709 B.n360 43.0261
R1985 B.n709 B.n356 43.0261
R1986 B.n715 B.n356 43.0261
R1987 B.n721 B.n352 43.0261
R1988 B.n721 B.n348 43.0261
R1989 B.n727 B.n348 43.0261
R1990 B.n727 B.n344 43.0261
R1991 B.n733 B.n344 43.0261
R1992 B.n733 B.n340 43.0261
R1993 B.n739 B.n340 43.0261
R1994 B.n739 B.n336 43.0261
R1995 B.n745 B.n336 43.0261
R1996 B.n745 B.n332 43.0261
R1997 B.n751 B.n332 43.0261
R1998 B.n757 B.n328 43.0261
R1999 B.n757 B.n324 43.0261
R2000 B.n764 B.n324 43.0261
R2001 B.n764 B.n320 43.0261
R2002 B.n770 B.n320 43.0261
R2003 B.n770 B.n4 43.0261
R2004 B.n924 B.n4 43.0261
R2005 B.n924 B.n923 43.0261
R2006 B.n923 B.n922 43.0261
R2007 B.n922 B.n8 43.0261
R2008 B.n12 B.n8 43.0261
R2009 B.n915 B.n12 43.0261
R2010 B.n915 B.n914 43.0261
R2011 B.n914 B.n913 43.0261
R2012 B.n913 B.n16 43.0261
R2013 B.n907 B.n906 43.0261
R2014 B.n906 B.n905 43.0261
R2015 B.n905 B.n23 43.0261
R2016 B.n899 B.n23 43.0261
R2017 B.n899 B.n898 43.0261
R2018 B.n898 B.n897 43.0261
R2019 B.n897 B.n30 43.0261
R2020 B.n891 B.n30 43.0261
R2021 B.n891 B.n890 43.0261
R2022 B.n890 B.n889 43.0261
R2023 B.n889 B.n37 43.0261
R2024 B.n883 B.n882 43.0261
R2025 B.n882 B.n881 43.0261
R2026 B.n881 B.n44 43.0261
R2027 B.n875 B.n44 43.0261
R2028 B.n875 B.n874 43.0261
R2029 B.n874 B.n873 43.0261
R2030 B.n873 B.n51 43.0261
R2031 B.n867 B.n51 43.0261
R2032 B.n867 B.n866 43.0261
R2033 B.n866 B.n865 43.0261
R2034 B.n865 B.n58 43.0261
R2035 B.n859 B.n58 43.0261
R2036 B.n859 B.n858 43.0261
R2037 B.n858 B.n857 43.0261
R2038 B.n851 B.n68 43.0261
R2039 B.n851 B.n850 43.0261
R2040 B.n850 B.n849 43.0261
R2041 B.n849 B.n72 43.0261
R2042 B.n843 B.n72 43.0261
R2043 B.n843 B.n842 43.0261
R2044 B.n842 B.n841 43.0261
R2045 B.n841 B.n79 43.0261
R2046 B.n835 B.n79 43.0261
R2047 B.n644 B.n401 35.4346
R2048 B.n640 B.n639 35.4346
R2049 B.n832 B.n831 35.4346
R2050 B.n837 B.n81 35.4346
R2051 B.n751 B.t1 35.4333
R2052 B.n907 B.t2 35.4333
R2053 B.n673 B.t12 29.1061
R2054 B.n715 B.t0 29.1061
R2055 B.n883 B.t3 29.1061
R2056 B.n857 B.t5 29.1061
R2057 B B.n927 18.0485
R2058 B.n666 B.t12 13.9205
R2059 B.t0 B.n352 13.9205
R2060 B.t3 B.n37 13.9205
R2061 B.n68 B.t5 13.9205
R2062 B.n645 B.n644 10.6151
R2063 B.n646 B.n645 10.6151
R2064 B.n646 B.n393 10.6151
R2065 B.n656 B.n393 10.6151
R2066 B.n657 B.n656 10.6151
R2067 B.n658 B.n657 10.6151
R2068 B.n658 B.n385 10.6151
R2069 B.n669 B.n385 10.6151
R2070 B.n670 B.n669 10.6151
R2071 B.n671 B.n670 10.6151
R2072 B.n671 B.n378 10.6151
R2073 B.n681 B.n378 10.6151
R2074 B.n682 B.n681 10.6151
R2075 B.n683 B.n682 10.6151
R2076 B.n683 B.n370 10.6151
R2077 B.n693 B.n370 10.6151
R2078 B.n694 B.n693 10.6151
R2079 B.n695 B.n694 10.6151
R2080 B.n695 B.n362 10.6151
R2081 B.n705 B.n362 10.6151
R2082 B.n706 B.n705 10.6151
R2083 B.n707 B.n706 10.6151
R2084 B.n707 B.n354 10.6151
R2085 B.n717 B.n354 10.6151
R2086 B.n718 B.n717 10.6151
R2087 B.n719 B.n718 10.6151
R2088 B.n719 B.n346 10.6151
R2089 B.n729 B.n346 10.6151
R2090 B.n730 B.n729 10.6151
R2091 B.n731 B.n730 10.6151
R2092 B.n731 B.n338 10.6151
R2093 B.n741 B.n338 10.6151
R2094 B.n742 B.n741 10.6151
R2095 B.n743 B.n742 10.6151
R2096 B.n743 B.n330 10.6151
R2097 B.n753 B.n330 10.6151
R2098 B.n754 B.n753 10.6151
R2099 B.n755 B.n754 10.6151
R2100 B.n755 B.n322 10.6151
R2101 B.n766 B.n322 10.6151
R2102 B.n767 B.n766 10.6151
R2103 B.n768 B.n767 10.6151
R2104 B.n768 B.n0 10.6151
R2105 B.n453 B.n401 10.6151
R2106 B.n453 B.n452 10.6151
R2107 B.n459 B.n452 10.6151
R2108 B.n460 B.n459 10.6151
R2109 B.n461 B.n460 10.6151
R2110 B.n461 B.n450 10.6151
R2111 B.n467 B.n450 10.6151
R2112 B.n468 B.n467 10.6151
R2113 B.n469 B.n468 10.6151
R2114 B.n469 B.n448 10.6151
R2115 B.n475 B.n448 10.6151
R2116 B.n476 B.n475 10.6151
R2117 B.n477 B.n476 10.6151
R2118 B.n477 B.n446 10.6151
R2119 B.n483 B.n446 10.6151
R2120 B.n484 B.n483 10.6151
R2121 B.n485 B.n484 10.6151
R2122 B.n485 B.n444 10.6151
R2123 B.n491 B.n444 10.6151
R2124 B.n492 B.n491 10.6151
R2125 B.n493 B.n492 10.6151
R2126 B.n493 B.n442 10.6151
R2127 B.n499 B.n442 10.6151
R2128 B.n500 B.n499 10.6151
R2129 B.n501 B.n500 10.6151
R2130 B.n501 B.n440 10.6151
R2131 B.n507 B.n440 10.6151
R2132 B.n508 B.n507 10.6151
R2133 B.n509 B.n508 10.6151
R2134 B.n509 B.n438 10.6151
R2135 B.n515 B.n438 10.6151
R2136 B.n516 B.n515 10.6151
R2137 B.n517 B.n516 10.6151
R2138 B.n517 B.n436 10.6151
R2139 B.n523 B.n436 10.6151
R2140 B.n524 B.n523 10.6151
R2141 B.n525 B.n524 10.6151
R2142 B.n525 B.n434 10.6151
R2143 B.n531 B.n434 10.6151
R2144 B.n532 B.n531 10.6151
R2145 B.n536 B.n532 10.6151
R2146 B.n542 B.n432 10.6151
R2147 B.n543 B.n542 10.6151
R2148 B.n544 B.n543 10.6151
R2149 B.n544 B.n430 10.6151
R2150 B.n550 B.n430 10.6151
R2151 B.n551 B.n550 10.6151
R2152 B.n552 B.n551 10.6151
R2153 B.n552 B.n428 10.6151
R2154 B.n559 B.n558 10.6151
R2155 B.n560 B.n559 10.6151
R2156 B.n560 B.n423 10.6151
R2157 B.n566 B.n423 10.6151
R2158 B.n567 B.n566 10.6151
R2159 B.n568 B.n567 10.6151
R2160 B.n568 B.n421 10.6151
R2161 B.n574 B.n421 10.6151
R2162 B.n575 B.n574 10.6151
R2163 B.n576 B.n575 10.6151
R2164 B.n576 B.n419 10.6151
R2165 B.n582 B.n419 10.6151
R2166 B.n583 B.n582 10.6151
R2167 B.n584 B.n583 10.6151
R2168 B.n584 B.n417 10.6151
R2169 B.n590 B.n417 10.6151
R2170 B.n591 B.n590 10.6151
R2171 B.n592 B.n591 10.6151
R2172 B.n592 B.n415 10.6151
R2173 B.n598 B.n415 10.6151
R2174 B.n599 B.n598 10.6151
R2175 B.n600 B.n599 10.6151
R2176 B.n600 B.n413 10.6151
R2177 B.n606 B.n413 10.6151
R2178 B.n607 B.n606 10.6151
R2179 B.n608 B.n607 10.6151
R2180 B.n608 B.n411 10.6151
R2181 B.n614 B.n411 10.6151
R2182 B.n615 B.n614 10.6151
R2183 B.n616 B.n615 10.6151
R2184 B.n616 B.n409 10.6151
R2185 B.n622 B.n409 10.6151
R2186 B.n623 B.n622 10.6151
R2187 B.n624 B.n623 10.6151
R2188 B.n624 B.n407 10.6151
R2189 B.n630 B.n407 10.6151
R2190 B.n631 B.n630 10.6151
R2191 B.n632 B.n631 10.6151
R2192 B.n632 B.n405 10.6151
R2193 B.n638 B.n405 10.6151
R2194 B.n639 B.n638 10.6151
R2195 B.n640 B.n397 10.6151
R2196 B.n650 B.n397 10.6151
R2197 B.n651 B.n650 10.6151
R2198 B.n652 B.n651 10.6151
R2199 B.n652 B.n389 10.6151
R2200 B.n662 B.n389 10.6151
R2201 B.n663 B.n662 10.6151
R2202 B.n664 B.n663 10.6151
R2203 B.n664 B.n382 10.6151
R2204 B.n675 B.n382 10.6151
R2205 B.n676 B.n675 10.6151
R2206 B.n677 B.n676 10.6151
R2207 B.n677 B.n374 10.6151
R2208 B.n687 B.n374 10.6151
R2209 B.n688 B.n687 10.6151
R2210 B.n689 B.n688 10.6151
R2211 B.n689 B.n366 10.6151
R2212 B.n699 B.n366 10.6151
R2213 B.n700 B.n699 10.6151
R2214 B.n701 B.n700 10.6151
R2215 B.n701 B.n358 10.6151
R2216 B.n711 B.n358 10.6151
R2217 B.n712 B.n711 10.6151
R2218 B.n713 B.n712 10.6151
R2219 B.n713 B.n350 10.6151
R2220 B.n723 B.n350 10.6151
R2221 B.n724 B.n723 10.6151
R2222 B.n725 B.n724 10.6151
R2223 B.n725 B.n342 10.6151
R2224 B.n735 B.n342 10.6151
R2225 B.n736 B.n735 10.6151
R2226 B.n737 B.n736 10.6151
R2227 B.n737 B.n334 10.6151
R2228 B.n747 B.n334 10.6151
R2229 B.n748 B.n747 10.6151
R2230 B.n749 B.n748 10.6151
R2231 B.n749 B.n326 10.6151
R2232 B.n759 B.n326 10.6151
R2233 B.n760 B.n759 10.6151
R2234 B.n762 B.n760 10.6151
R2235 B.n762 B.n761 10.6151
R2236 B.n761 B.n318 10.6151
R2237 B.n773 B.n318 10.6151
R2238 B.n774 B.n773 10.6151
R2239 B.n775 B.n774 10.6151
R2240 B.n776 B.n775 10.6151
R2241 B.n777 B.n776 10.6151
R2242 B.n780 B.n777 10.6151
R2243 B.n781 B.n780 10.6151
R2244 B.n782 B.n781 10.6151
R2245 B.n783 B.n782 10.6151
R2246 B.n785 B.n783 10.6151
R2247 B.n786 B.n785 10.6151
R2248 B.n787 B.n786 10.6151
R2249 B.n788 B.n787 10.6151
R2250 B.n790 B.n788 10.6151
R2251 B.n791 B.n790 10.6151
R2252 B.n792 B.n791 10.6151
R2253 B.n793 B.n792 10.6151
R2254 B.n795 B.n793 10.6151
R2255 B.n796 B.n795 10.6151
R2256 B.n797 B.n796 10.6151
R2257 B.n798 B.n797 10.6151
R2258 B.n800 B.n798 10.6151
R2259 B.n801 B.n800 10.6151
R2260 B.n802 B.n801 10.6151
R2261 B.n803 B.n802 10.6151
R2262 B.n805 B.n803 10.6151
R2263 B.n806 B.n805 10.6151
R2264 B.n807 B.n806 10.6151
R2265 B.n808 B.n807 10.6151
R2266 B.n810 B.n808 10.6151
R2267 B.n811 B.n810 10.6151
R2268 B.n812 B.n811 10.6151
R2269 B.n813 B.n812 10.6151
R2270 B.n815 B.n813 10.6151
R2271 B.n816 B.n815 10.6151
R2272 B.n817 B.n816 10.6151
R2273 B.n818 B.n817 10.6151
R2274 B.n820 B.n818 10.6151
R2275 B.n821 B.n820 10.6151
R2276 B.n822 B.n821 10.6151
R2277 B.n823 B.n822 10.6151
R2278 B.n825 B.n823 10.6151
R2279 B.n826 B.n825 10.6151
R2280 B.n827 B.n826 10.6151
R2281 B.n828 B.n827 10.6151
R2282 B.n830 B.n828 10.6151
R2283 B.n831 B.n830 10.6151
R2284 B.n919 B.n1 10.6151
R2285 B.n919 B.n918 10.6151
R2286 B.n918 B.n917 10.6151
R2287 B.n917 B.n10 10.6151
R2288 B.n911 B.n10 10.6151
R2289 B.n911 B.n910 10.6151
R2290 B.n910 B.n909 10.6151
R2291 B.n909 B.n18 10.6151
R2292 B.n903 B.n18 10.6151
R2293 B.n903 B.n902 10.6151
R2294 B.n902 B.n901 10.6151
R2295 B.n901 B.n25 10.6151
R2296 B.n895 B.n25 10.6151
R2297 B.n895 B.n894 10.6151
R2298 B.n894 B.n893 10.6151
R2299 B.n893 B.n32 10.6151
R2300 B.n887 B.n32 10.6151
R2301 B.n887 B.n886 10.6151
R2302 B.n886 B.n885 10.6151
R2303 B.n885 B.n39 10.6151
R2304 B.n879 B.n39 10.6151
R2305 B.n879 B.n878 10.6151
R2306 B.n878 B.n877 10.6151
R2307 B.n877 B.n46 10.6151
R2308 B.n871 B.n46 10.6151
R2309 B.n871 B.n870 10.6151
R2310 B.n870 B.n869 10.6151
R2311 B.n869 B.n53 10.6151
R2312 B.n863 B.n53 10.6151
R2313 B.n863 B.n862 10.6151
R2314 B.n862 B.n861 10.6151
R2315 B.n861 B.n60 10.6151
R2316 B.n855 B.n60 10.6151
R2317 B.n855 B.n854 10.6151
R2318 B.n854 B.n853 10.6151
R2319 B.n853 B.n66 10.6151
R2320 B.n847 B.n66 10.6151
R2321 B.n847 B.n846 10.6151
R2322 B.n846 B.n845 10.6151
R2323 B.n845 B.n74 10.6151
R2324 B.n839 B.n74 10.6151
R2325 B.n839 B.n838 10.6151
R2326 B.n838 B.n837 10.6151
R2327 B.n136 B.n81 10.6151
R2328 B.n139 B.n136 10.6151
R2329 B.n140 B.n139 10.6151
R2330 B.n143 B.n140 10.6151
R2331 B.n144 B.n143 10.6151
R2332 B.n147 B.n144 10.6151
R2333 B.n148 B.n147 10.6151
R2334 B.n151 B.n148 10.6151
R2335 B.n152 B.n151 10.6151
R2336 B.n155 B.n152 10.6151
R2337 B.n156 B.n155 10.6151
R2338 B.n159 B.n156 10.6151
R2339 B.n160 B.n159 10.6151
R2340 B.n163 B.n160 10.6151
R2341 B.n164 B.n163 10.6151
R2342 B.n167 B.n164 10.6151
R2343 B.n168 B.n167 10.6151
R2344 B.n171 B.n168 10.6151
R2345 B.n172 B.n171 10.6151
R2346 B.n175 B.n172 10.6151
R2347 B.n176 B.n175 10.6151
R2348 B.n179 B.n176 10.6151
R2349 B.n180 B.n179 10.6151
R2350 B.n183 B.n180 10.6151
R2351 B.n184 B.n183 10.6151
R2352 B.n187 B.n184 10.6151
R2353 B.n188 B.n187 10.6151
R2354 B.n191 B.n188 10.6151
R2355 B.n192 B.n191 10.6151
R2356 B.n195 B.n192 10.6151
R2357 B.n196 B.n195 10.6151
R2358 B.n199 B.n196 10.6151
R2359 B.n200 B.n199 10.6151
R2360 B.n203 B.n200 10.6151
R2361 B.n204 B.n203 10.6151
R2362 B.n207 B.n204 10.6151
R2363 B.n208 B.n207 10.6151
R2364 B.n211 B.n208 10.6151
R2365 B.n212 B.n211 10.6151
R2366 B.n215 B.n212 10.6151
R2367 B.n216 B.n215 10.6151
R2368 B.n220 B.n219 10.6151
R2369 B.n223 B.n220 10.6151
R2370 B.n224 B.n223 10.6151
R2371 B.n227 B.n224 10.6151
R2372 B.n228 B.n227 10.6151
R2373 B.n231 B.n228 10.6151
R2374 B.n232 B.n231 10.6151
R2375 B.n235 B.n232 10.6151
R2376 B.n240 B.n237 10.6151
R2377 B.n241 B.n240 10.6151
R2378 B.n244 B.n241 10.6151
R2379 B.n245 B.n244 10.6151
R2380 B.n248 B.n245 10.6151
R2381 B.n249 B.n248 10.6151
R2382 B.n252 B.n249 10.6151
R2383 B.n253 B.n252 10.6151
R2384 B.n256 B.n253 10.6151
R2385 B.n257 B.n256 10.6151
R2386 B.n260 B.n257 10.6151
R2387 B.n261 B.n260 10.6151
R2388 B.n264 B.n261 10.6151
R2389 B.n265 B.n264 10.6151
R2390 B.n268 B.n265 10.6151
R2391 B.n269 B.n268 10.6151
R2392 B.n272 B.n269 10.6151
R2393 B.n273 B.n272 10.6151
R2394 B.n276 B.n273 10.6151
R2395 B.n277 B.n276 10.6151
R2396 B.n280 B.n277 10.6151
R2397 B.n281 B.n280 10.6151
R2398 B.n284 B.n281 10.6151
R2399 B.n285 B.n284 10.6151
R2400 B.n288 B.n285 10.6151
R2401 B.n289 B.n288 10.6151
R2402 B.n292 B.n289 10.6151
R2403 B.n293 B.n292 10.6151
R2404 B.n296 B.n293 10.6151
R2405 B.n297 B.n296 10.6151
R2406 B.n300 B.n297 10.6151
R2407 B.n301 B.n300 10.6151
R2408 B.n304 B.n301 10.6151
R2409 B.n305 B.n304 10.6151
R2410 B.n308 B.n305 10.6151
R2411 B.n309 B.n308 10.6151
R2412 B.n312 B.n309 10.6151
R2413 B.n313 B.n312 10.6151
R2414 B.n316 B.n313 10.6151
R2415 B.n317 B.n316 10.6151
R2416 B.n832 B.n317 10.6151
R2417 B.n927 B.n0 8.11757
R2418 B.n927 B.n1 8.11757
R2419 B.t1 B.n328 7.59325
R2420 B.t2 B.n16 7.59325
R2421 B.n535 B.n432 6.5566
R2422 B.n428 B.n427 6.5566
R2423 B.n219 B.n135 6.5566
R2424 B.n236 B.n235 6.5566
R2425 B.n536 B.n535 4.05904
R2426 B.n558 B.n427 4.05904
R2427 B.n216 B.n135 4.05904
R2428 B.n237 B.n236 4.05904
R2429 VN.n1 VN.t2 110.746
R2430 VN.n0 VN.t1 110.746
R2431 VN.n0 VN.t0 109.395
R2432 VN.n1 VN.t3 109.395
R2433 VN VN.n1 52.1492
R2434 VN VN.n0 1.85758
R2435 VDD2.n2 VDD2.n0 106.522
R2436 VDD2.n2 VDD2.n1 61.6858
R2437 VDD2.n1 VDD2.t0 1.63551
R2438 VDD2.n1 VDD2.t1 1.63551
R2439 VDD2.n0 VDD2.t2 1.63551
R2440 VDD2.n0 VDD2.t3 1.63551
R2441 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 5.77112f
C1 VTAIL VDD2 5.83338f
C2 VN VDD1 0.149939f
C3 VTAIL VP 5.1727f
C4 VN VDD2 5.07978f
C5 VN VP 7.07667f
C6 VDD1 VDD2 1.31767f
C7 VDD1 VP 5.39932f
C8 VDD2 VP 0.470518f
C9 VN VTAIL 5.15859f
C10 VDD2 B 4.451731f
C11 VDD1 B 9.07682f
C12 VTAIL B 10.79778f
C13 VN B 13.046181f
C14 VP B 11.495604f
C15 VDD2.t2 B 0.260919f
C16 VDD2.t3 B 0.260919f
C17 VDD2.n0 B 3.07964f
C18 VDD2.t0 B 0.260919f
C19 VDD2.t1 B 0.260919f
C20 VDD2.n1 B 2.32578f
C21 VDD2.n2 B 4.13224f
C22 VN.t0 B 2.81491f
C23 VN.t1 B 2.82702f
C24 VN.n0 B 1.68315f
C25 VN.t3 B 2.81491f
C26 VN.t2 B 2.82702f
C27 VN.n1 B 3.00222f
C28 VTAIL.n0 B 0.024055f
C29 VTAIL.n1 B 0.017196f
C30 VTAIL.n2 B 0.009241f
C31 VTAIL.n3 B 0.021841f
C32 VTAIL.n4 B 0.009784f
C33 VTAIL.n5 B 0.017196f
C34 VTAIL.n6 B 0.009241f
C35 VTAIL.n7 B 0.021841f
C36 VTAIL.n8 B 0.009784f
C37 VTAIL.n9 B 0.017196f
C38 VTAIL.n10 B 0.009512f
C39 VTAIL.n11 B 0.021841f
C40 VTAIL.n12 B 0.009784f
C41 VTAIL.n13 B 0.017196f
C42 VTAIL.n14 B 0.009241f
C43 VTAIL.n15 B 0.021841f
C44 VTAIL.n16 B 0.009784f
C45 VTAIL.n17 B 0.017196f
C46 VTAIL.n18 B 0.009241f
C47 VTAIL.n19 B 0.016381f
C48 VTAIL.n20 B 0.01544f
C49 VTAIL.t2 B 0.036899f
C50 VTAIL.n21 B 0.12471f
C51 VTAIL.n22 B 0.875937f
C52 VTAIL.n23 B 0.009241f
C53 VTAIL.n24 B 0.009784f
C54 VTAIL.n25 B 0.021841f
C55 VTAIL.n26 B 0.021841f
C56 VTAIL.n27 B 0.009784f
C57 VTAIL.n28 B 0.009241f
C58 VTAIL.n29 B 0.017196f
C59 VTAIL.n30 B 0.017196f
C60 VTAIL.n31 B 0.009241f
C61 VTAIL.n32 B 0.009784f
C62 VTAIL.n33 B 0.021841f
C63 VTAIL.n34 B 0.021841f
C64 VTAIL.n35 B 0.009784f
C65 VTAIL.n36 B 0.009241f
C66 VTAIL.n37 B 0.017196f
C67 VTAIL.n38 B 0.017196f
C68 VTAIL.n39 B 0.009241f
C69 VTAIL.n40 B 0.009241f
C70 VTAIL.n41 B 0.009784f
C71 VTAIL.n42 B 0.021841f
C72 VTAIL.n43 B 0.021841f
C73 VTAIL.n44 B 0.021841f
C74 VTAIL.n45 B 0.009512f
C75 VTAIL.n46 B 0.009241f
C76 VTAIL.n47 B 0.017196f
C77 VTAIL.n48 B 0.017196f
C78 VTAIL.n49 B 0.009241f
C79 VTAIL.n50 B 0.009784f
C80 VTAIL.n51 B 0.021841f
C81 VTAIL.n52 B 0.021841f
C82 VTAIL.n53 B 0.009784f
C83 VTAIL.n54 B 0.009241f
C84 VTAIL.n55 B 0.017196f
C85 VTAIL.n56 B 0.017196f
C86 VTAIL.n57 B 0.009241f
C87 VTAIL.n58 B 0.009784f
C88 VTAIL.n59 B 0.021841f
C89 VTAIL.n60 B 0.047077f
C90 VTAIL.n61 B 0.009784f
C91 VTAIL.n62 B 0.009241f
C92 VTAIL.n63 B 0.039514f
C93 VTAIL.n64 B 0.026313f
C94 VTAIL.n65 B 0.142452f
C95 VTAIL.n66 B 0.024055f
C96 VTAIL.n67 B 0.017196f
C97 VTAIL.n68 B 0.009241f
C98 VTAIL.n69 B 0.021841f
C99 VTAIL.n70 B 0.009784f
C100 VTAIL.n71 B 0.017196f
C101 VTAIL.n72 B 0.009241f
C102 VTAIL.n73 B 0.021841f
C103 VTAIL.n74 B 0.009784f
C104 VTAIL.n75 B 0.017196f
C105 VTAIL.n76 B 0.009512f
C106 VTAIL.n77 B 0.021841f
C107 VTAIL.n78 B 0.009784f
C108 VTAIL.n79 B 0.017196f
C109 VTAIL.n80 B 0.009241f
C110 VTAIL.n81 B 0.021841f
C111 VTAIL.n82 B 0.009784f
C112 VTAIL.n83 B 0.017196f
C113 VTAIL.n84 B 0.009241f
C114 VTAIL.n85 B 0.016381f
C115 VTAIL.n86 B 0.01544f
C116 VTAIL.t4 B 0.036899f
C117 VTAIL.n87 B 0.12471f
C118 VTAIL.n88 B 0.875937f
C119 VTAIL.n89 B 0.009241f
C120 VTAIL.n90 B 0.009784f
C121 VTAIL.n91 B 0.021841f
C122 VTAIL.n92 B 0.021841f
C123 VTAIL.n93 B 0.009784f
C124 VTAIL.n94 B 0.009241f
C125 VTAIL.n95 B 0.017196f
C126 VTAIL.n96 B 0.017196f
C127 VTAIL.n97 B 0.009241f
C128 VTAIL.n98 B 0.009784f
C129 VTAIL.n99 B 0.021841f
C130 VTAIL.n100 B 0.021841f
C131 VTAIL.n101 B 0.009784f
C132 VTAIL.n102 B 0.009241f
C133 VTAIL.n103 B 0.017196f
C134 VTAIL.n104 B 0.017196f
C135 VTAIL.n105 B 0.009241f
C136 VTAIL.n106 B 0.009241f
C137 VTAIL.n107 B 0.009784f
C138 VTAIL.n108 B 0.021841f
C139 VTAIL.n109 B 0.021841f
C140 VTAIL.n110 B 0.021841f
C141 VTAIL.n111 B 0.009512f
C142 VTAIL.n112 B 0.009241f
C143 VTAIL.n113 B 0.017196f
C144 VTAIL.n114 B 0.017196f
C145 VTAIL.n115 B 0.009241f
C146 VTAIL.n116 B 0.009784f
C147 VTAIL.n117 B 0.021841f
C148 VTAIL.n118 B 0.021841f
C149 VTAIL.n119 B 0.009784f
C150 VTAIL.n120 B 0.009241f
C151 VTAIL.n121 B 0.017196f
C152 VTAIL.n122 B 0.017196f
C153 VTAIL.n123 B 0.009241f
C154 VTAIL.n124 B 0.009784f
C155 VTAIL.n125 B 0.021841f
C156 VTAIL.n126 B 0.047077f
C157 VTAIL.n127 B 0.009784f
C158 VTAIL.n128 B 0.009241f
C159 VTAIL.n129 B 0.039514f
C160 VTAIL.n130 B 0.026313f
C161 VTAIL.n131 B 0.237867f
C162 VTAIL.n132 B 0.024055f
C163 VTAIL.n133 B 0.017196f
C164 VTAIL.n134 B 0.009241f
C165 VTAIL.n135 B 0.021841f
C166 VTAIL.n136 B 0.009784f
C167 VTAIL.n137 B 0.017196f
C168 VTAIL.n138 B 0.009241f
C169 VTAIL.n139 B 0.021841f
C170 VTAIL.n140 B 0.009784f
C171 VTAIL.n141 B 0.017196f
C172 VTAIL.n142 B 0.009512f
C173 VTAIL.n143 B 0.021841f
C174 VTAIL.n144 B 0.009784f
C175 VTAIL.n145 B 0.017196f
C176 VTAIL.n146 B 0.009241f
C177 VTAIL.n147 B 0.021841f
C178 VTAIL.n148 B 0.009784f
C179 VTAIL.n149 B 0.017196f
C180 VTAIL.n150 B 0.009241f
C181 VTAIL.n151 B 0.016381f
C182 VTAIL.n152 B 0.01544f
C183 VTAIL.t5 B 0.036899f
C184 VTAIL.n153 B 0.12471f
C185 VTAIL.n154 B 0.875937f
C186 VTAIL.n155 B 0.009241f
C187 VTAIL.n156 B 0.009784f
C188 VTAIL.n157 B 0.021841f
C189 VTAIL.n158 B 0.021841f
C190 VTAIL.n159 B 0.009784f
C191 VTAIL.n160 B 0.009241f
C192 VTAIL.n161 B 0.017196f
C193 VTAIL.n162 B 0.017196f
C194 VTAIL.n163 B 0.009241f
C195 VTAIL.n164 B 0.009784f
C196 VTAIL.n165 B 0.021841f
C197 VTAIL.n166 B 0.021841f
C198 VTAIL.n167 B 0.009784f
C199 VTAIL.n168 B 0.009241f
C200 VTAIL.n169 B 0.017196f
C201 VTAIL.n170 B 0.017196f
C202 VTAIL.n171 B 0.009241f
C203 VTAIL.n172 B 0.009241f
C204 VTAIL.n173 B 0.009784f
C205 VTAIL.n174 B 0.021841f
C206 VTAIL.n175 B 0.021841f
C207 VTAIL.n176 B 0.021841f
C208 VTAIL.n177 B 0.009512f
C209 VTAIL.n178 B 0.009241f
C210 VTAIL.n179 B 0.017196f
C211 VTAIL.n180 B 0.017196f
C212 VTAIL.n181 B 0.009241f
C213 VTAIL.n182 B 0.009784f
C214 VTAIL.n183 B 0.021841f
C215 VTAIL.n184 B 0.021841f
C216 VTAIL.n185 B 0.009784f
C217 VTAIL.n186 B 0.009241f
C218 VTAIL.n187 B 0.017196f
C219 VTAIL.n188 B 0.017196f
C220 VTAIL.n189 B 0.009241f
C221 VTAIL.n190 B 0.009784f
C222 VTAIL.n191 B 0.021841f
C223 VTAIL.n192 B 0.047077f
C224 VTAIL.n193 B 0.009784f
C225 VTAIL.n194 B 0.009241f
C226 VTAIL.n195 B 0.039514f
C227 VTAIL.n196 B 0.026313f
C228 VTAIL.n197 B 1.22117f
C229 VTAIL.n198 B 0.024055f
C230 VTAIL.n199 B 0.017196f
C231 VTAIL.n200 B 0.009241f
C232 VTAIL.n201 B 0.021841f
C233 VTAIL.n202 B 0.009784f
C234 VTAIL.n203 B 0.017196f
C235 VTAIL.n204 B 0.009241f
C236 VTAIL.n205 B 0.021841f
C237 VTAIL.n206 B 0.009784f
C238 VTAIL.n207 B 0.017196f
C239 VTAIL.n208 B 0.009512f
C240 VTAIL.n209 B 0.021841f
C241 VTAIL.n210 B 0.009241f
C242 VTAIL.n211 B 0.009784f
C243 VTAIL.n212 B 0.017196f
C244 VTAIL.n213 B 0.009241f
C245 VTAIL.n214 B 0.021841f
C246 VTAIL.n215 B 0.009784f
C247 VTAIL.n216 B 0.017196f
C248 VTAIL.n217 B 0.009241f
C249 VTAIL.n218 B 0.016381f
C250 VTAIL.n219 B 0.01544f
C251 VTAIL.t0 B 0.036899f
C252 VTAIL.n220 B 0.12471f
C253 VTAIL.n221 B 0.875937f
C254 VTAIL.n222 B 0.009241f
C255 VTAIL.n223 B 0.009784f
C256 VTAIL.n224 B 0.021841f
C257 VTAIL.n225 B 0.021841f
C258 VTAIL.n226 B 0.009784f
C259 VTAIL.n227 B 0.009241f
C260 VTAIL.n228 B 0.017196f
C261 VTAIL.n229 B 0.017196f
C262 VTAIL.n230 B 0.009241f
C263 VTAIL.n231 B 0.009784f
C264 VTAIL.n232 B 0.021841f
C265 VTAIL.n233 B 0.021841f
C266 VTAIL.n234 B 0.009784f
C267 VTAIL.n235 B 0.009241f
C268 VTAIL.n236 B 0.017196f
C269 VTAIL.n237 B 0.017196f
C270 VTAIL.n238 B 0.009241f
C271 VTAIL.n239 B 0.009784f
C272 VTAIL.n240 B 0.021841f
C273 VTAIL.n241 B 0.021841f
C274 VTAIL.n242 B 0.021841f
C275 VTAIL.n243 B 0.009512f
C276 VTAIL.n244 B 0.009241f
C277 VTAIL.n245 B 0.017196f
C278 VTAIL.n246 B 0.017196f
C279 VTAIL.n247 B 0.009241f
C280 VTAIL.n248 B 0.009784f
C281 VTAIL.n249 B 0.021841f
C282 VTAIL.n250 B 0.021841f
C283 VTAIL.n251 B 0.009784f
C284 VTAIL.n252 B 0.009241f
C285 VTAIL.n253 B 0.017196f
C286 VTAIL.n254 B 0.017196f
C287 VTAIL.n255 B 0.009241f
C288 VTAIL.n256 B 0.009784f
C289 VTAIL.n257 B 0.021841f
C290 VTAIL.n258 B 0.047077f
C291 VTAIL.n259 B 0.009784f
C292 VTAIL.n260 B 0.009241f
C293 VTAIL.n261 B 0.039514f
C294 VTAIL.n262 B 0.026313f
C295 VTAIL.n263 B 1.22117f
C296 VTAIL.n264 B 0.024055f
C297 VTAIL.n265 B 0.017196f
C298 VTAIL.n266 B 0.009241f
C299 VTAIL.n267 B 0.021841f
C300 VTAIL.n268 B 0.009784f
C301 VTAIL.n269 B 0.017196f
C302 VTAIL.n270 B 0.009241f
C303 VTAIL.n271 B 0.021841f
C304 VTAIL.n272 B 0.009784f
C305 VTAIL.n273 B 0.017196f
C306 VTAIL.n274 B 0.009512f
C307 VTAIL.n275 B 0.021841f
C308 VTAIL.n276 B 0.009241f
C309 VTAIL.n277 B 0.009784f
C310 VTAIL.n278 B 0.017196f
C311 VTAIL.n279 B 0.009241f
C312 VTAIL.n280 B 0.021841f
C313 VTAIL.n281 B 0.009784f
C314 VTAIL.n282 B 0.017196f
C315 VTAIL.n283 B 0.009241f
C316 VTAIL.n284 B 0.016381f
C317 VTAIL.n285 B 0.01544f
C318 VTAIL.t1 B 0.036899f
C319 VTAIL.n286 B 0.12471f
C320 VTAIL.n287 B 0.875937f
C321 VTAIL.n288 B 0.009241f
C322 VTAIL.n289 B 0.009784f
C323 VTAIL.n290 B 0.021841f
C324 VTAIL.n291 B 0.021841f
C325 VTAIL.n292 B 0.009784f
C326 VTAIL.n293 B 0.009241f
C327 VTAIL.n294 B 0.017196f
C328 VTAIL.n295 B 0.017196f
C329 VTAIL.n296 B 0.009241f
C330 VTAIL.n297 B 0.009784f
C331 VTAIL.n298 B 0.021841f
C332 VTAIL.n299 B 0.021841f
C333 VTAIL.n300 B 0.009784f
C334 VTAIL.n301 B 0.009241f
C335 VTAIL.n302 B 0.017196f
C336 VTAIL.n303 B 0.017196f
C337 VTAIL.n304 B 0.009241f
C338 VTAIL.n305 B 0.009784f
C339 VTAIL.n306 B 0.021841f
C340 VTAIL.n307 B 0.021841f
C341 VTAIL.n308 B 0.021841f
C342 VTAIL.n309 B 0.009512f
C343 VTAIL.n310 B 0.009241f
C344 VTAIL.n311 B 0.017196f
C345 VTAIL.n312 B 0.017196f
C346 VTAIL.n313 B 0.009241f
C347 VTAIL.n314 B 0.009784f
C348 VTAIL.n315 B 0.021841f
C349 VTAIL.n316 B 0.021841f
C350 VTAIL.n317 B 0.009784f
C351 VTAIL.n318 B 0.009241f
C352 VTAIL.n319 B 0.017196f
C353 VTAIL.n320 B 0.017196f
C354 VTAIL.n321 B 0.009241f
C355 VTAIL.n322 B 0.009784f
C356 VTAIL.n323 B 0.021841f
C357 VTAIL.n324 B 0.047077f
C358 VTAIL.n325 B 0.009784f
C359 VTAIL.n326 B 0.009241f
C360 VTAIL.n327 B 0.039514f
C361 VTAIL.n328 B 0.026313f
C362 VTAIL.n329 B 0.237867f
C363 VTAIL.n330 B 0.024055f
C364 VTAIL.n331 B 0.017196f
C365 VTAIL.n332 B 0.009241f
C366 VTAIL.n333 B 0.021841f
C367 VTAIL.n334 B 0.009784f
C368 VTAIL.n335 B 0.017196f
C369 VTAIL.n336 B 0.009241f
C370 VTAIL.n337 B 0.021841f
C371 VTAIL.n338 B 0.009784f
C372 VTAIL.n339 B 0.017196f
C373 VTAIL.n340 B 0.009512f
C374 VTAIL.n341 B 0.021841f
C375 VTAIL.n342 B 0.009241f
C376 VTAIL.n343 B 0.009784f
C377 VTAIL.n344 B 0.017196f
C378 VTAIL.n345 B 0.009241f
C379 VTAIL.n346 B 0.021841f
C380 VTAIL.n347 B 0.009784f
C381 VTAIL.n348 B 0.017196f
C382 VTAIL.n349 B 0.009241f
C383 VTAIL.n350 B 0.016381f
C384 VTAIL.n351 B 0.01544f
C385 VTAIL.t7 B 0.036899f
C386 VTAIL.n352 B 0.12471f
C387 VTAIL.n353 B 0.875937f
C388 VTAIL.n354 B 0.009241f
C389 VTAIL.n355 B 0.009784f
C390 VTAIL.n356 B 0.021841f
C391 VTAIL.n357 B 0.021841f
C392 VTAIL.n358 B 0.009784f
C393 VTAIL.n359 B 0.009241f
C394 VTAIL.n360 B 0.017196f
C395 VTAIL.n361 B 0.017196f
C396 VTAIL.n362 B 0.009241f
C397 VTAIL.n363 B 0.009784f
C398 VTAIL.n364 B 0.021841f
C399 VTAIL.n365 B 0.021841f
C400 VTAIL.n366 B 0.009784f
C401 VTAIL.n367 B 0.009241f
C402 VTAIL.n368 B 0.017196f
C403 VTAIL.n369 B 0.017196f
C404 VTAIL.n370 B 0.009241f
C405 VTAIL.n371 B 0.009784f
C406 VTAIL.n372 B 0.021841f
C407 VTAIL.n373 B 0.021841f
C408 VTAIL.n374 B 0.021841f
C409 VTAIL.n375 B 0.009512f
C410 VTAIL.n376 B 0.009241f
C411 VTAIL.n377 B 0.017196f
C412 VTAIL.n378 B 0.017196f
C413 VTAIL.n379 B 0.009241f
C414 VTAIL.n380 B 0.009784f
C415 VTAIL.n381 B 0.021841f
C416 VTAIL.n382 B 0.021841f
C417 VTAIL.n383 B 0.009784f
C418 VTAIL.n384 B 0.009241f
C419 VTAIL.n385 B 0.017196f
C420 VTAIL.n386 B 0.017196f
C421 VTAIL.n387 B 0.009241f
C422 VTAIL.n388 B 0.009784f
C423 VTAIL.n389 B 0.021841f
C424 VTAIL.n390 B 0.047077f
C425 VTAIL.n391 B 0.009784f
C426 VTAIL.n392 B 0.009241f
C427 VTAIL.n393 B 0.039514f
C428 VTAIL.n394 B 0.026313f
C429 VTAIL.n395 B 0.237867f
C430 VTAIL.n396 B 0.024055f
C431 VTAIL.n397 B 0.017196f
C432 VTAIL.n398 B 0.009241f
C433 VTAIL.n399 B 0.021841f
C434 VTAIL.n400 B 0.009784f
C435 VTAIL.n401 B 0.017196f
C436 VTAIL.n402 B 0.009241f
C437 VTAIL.n403 B 0.021841f
C438 VTAIL.n404 B 0.009784f
C439 VTAIL.n405 B 0.017196f
C440 VTAIL.n406 B 0.009512f
C441 VTAIL.n407 B 0.021841f
C442 VTAIL.n408 B 0.009241f
C443 VTAIL.n409 B 0.009784f
C444 VTAIL.n410 B 0.017196f
C445 VTAIL.n411 B 0.009241f
C446 VTAIL.n412 B 0.021841f
C447 VTAIL.n413 B 0.009784f
C448 VTAIL.n414 B 0.017196f
C449 VTAIL.n415 B 0.009241f
C450 VTAIL.n416 B 0.016381f
C451 VTAIL.n417 B 0.01544f
C452 VTAIL.t6 B 0.036899f
C453 VTAIL.n418 B 0.12471f
C454 VTAIL.n419 B 0.875937f
C455 VTAIL.n420 B 0.009241f
C456 VTAIL.n421 B 0.009784f
C457 VTAIL.n422 B 0.021841f
C458 VTAIL.n423 B 0.021841f
C459 VTAIL.n424 B 0.009784f
C460 VTAIL.n425 B 0.009241f
C461 VTAIL.n426 B 0.017196f
C462 VTAIL.n427 B 0.017196f
C463 VTAIL.n428 B 0.009241f
C464 VTAIL.n429 B 0.009784f
C465 VTAIL.n430 B 0.021841f
C466 VTAIL.n431 B 0.021841f
C467 VTAIL.n432 B 0.009784f
C468 VTAIL.n433 B 0.009241f
C469 VTAIL.n434 B 0.017196f
C470 VTAIL.n435 B 0.017196f
C471 VTAIL.n436 B 0.009241f
C472 VTAIL.n437 B 0.009784f
C473 VTAIL.n438 B 0.021841f
C474 VTAIL.n439 B 0.021841f
C475 VTAIL.n440 B 0.021841f
C476 VTAIL.n441 B 0.009512f
C477 VTAIL.n442 B 0.009241f
C478 VTAIL.n443 B 0.017196f
C479 VTAIL.n444 B 0.017196f
C480 VTAIL.n445 B 0.009241f
C481 VTAIL.n446 B 0.009784f
C482 VTAIL.n447 B 0.021841f
C483 VTAIL.n448 B 0.021841f
C484 VTAIL.n449 B 0.009784f
C485 VTAIL.n450 B 0.009241f
C486 VTAIL.n451 B 0.017196f
C487 VTAIL.n452 B 0.017196f
C488 VTAIL.n453 B 0.009241f
C489 VTAIL.n454 B 0.009784f
C490 VTAIL.n455 B 0.021841f
C491 VTAIL.n456 B 0.047077f
C492 VTAIL.n457 B 0.009784f
C493 VTAIL.n458 B 0.009241f
C494 VTAIL.n459 B 0.039514f
C495 VTAIL.n460 B 0.026313f
C496 VTAIL.n461 B 1.22117f
C497 VTAIL.n462 B 0.024055f
C498 VTAIL.n463 B 0.017196f
C499 VTAIL.n464 B 0.009241f
C500 VTAIL.n465 B 0.021841f
C501 VTAIL.n466 B 0.009784f
C502 VTAIL.n467 B 0.017196f
C503 VTAIL.n468 B 0.009241f
C504 VTAIL.n469 B 0.021841f
C505 VTAIL.n470 B 0.009784f
C506 VTAIL.n471 B 0.017196f
C507 VTAIL.n472 B 0.009512f
C508 VTAIL.n473 B 0.021841f
C509 VTAIL.n474 B 0.009784f
C510 VTAIL.n475 B 0.017196f
C511 VTAIL.n476 B 0.009241f
C512 VTAIL.n477 B 0.021841f
C513 VTAIL.n478 B 0.009784f
C514 VTAIL.n479 B 0.017196f
C515 VTAIL.n480 B 0.009241f
C516 VTAIL.n481 B 0.016381f
C517 VTAIL.n482 B 0.01544f
C518 VTAIL.t3 B 0.036899f
C519 VTAIL.n483 B 0.12471f
C520 VTAIL.n484 B 0.875937f
C521 VTAIL.n485 B 0.009241f
C522 VTAIL.n486 B 0.009784f
C523 VTAIL.n487 B 0.021841f
C524 VTAIL.n488 B 0.021841f
C525 VTAIL.n489 B 0.009784f
C526 VTAIL.n490 B 0.009241f
C527 VTAIL.n491 B 0.017196f
C528 VTAIL.n492 B 0.017196f
C529 VTAIL.n493 B 0.009241f
C530 VTAIL.n494 B 0.009784f
C531 VTAIL.n495 B 0.021841f
C532 VTAIL.n496 B 0.021841f
C533 VTAIL.n497 B 0.009784f
C534 VTAIL.n498 B 0.009241f
C535 VTAIL.n499 B 0.017196f
C536 VTAIL.n500 B 0.017196f
C537 VTAIL.n501 B 0.009241f
C538 VTAIL.n502 B 0.009241f
C539 VTAIL.n503 B 0.009784f
C540 VTAIL.n504 B 0.021841f
C541 VTAIL.n505 B 0.021841f
C542 VTAIL.n506 B 0.021841f
C543 VTAIL.n507 B 0.009512f
C544 VTAIL.n508 B 0.009241f
C545 VTAIL.n509 B 0.017196f
C546 VTAIL.n510 B 0.017196f
C547 VTAIL.n511 B 0.009241f
C548 VTAIL.n512 B 0.009784f
C549 VTAIL.n513 B 0.021841f
C550 VTAIL.n514 B 0.021841f
C551 VTAIL.n515 B 0.009784f
C552 VTAIL.n516 B 0.009241f
C553 VTAIL.n517 B 0.017196f
C554 VTAIL.n518 B 0.017196f
C555 VTAIL.n519 B 0.009241f
C556 VTAIL.n520 B 0.009784f
C557 VTAIL.n521 B 0.021841f
C558 VTAIL.n522 B 0.047077f
C559 VTAIL.n523 B 0.009784f
C560 VTAIL.n524 B 0.009241f
C561 VTAIL.n525 B 0.039514f
C562 VTAIL.n526 B 0.026313f
C563 VTAIL.n527 B 1.11931f
C564 VDD1.t2 B 0.265646f
C565 VDD1.t3 B 0.265646f
C566 VDD1.n0 B 2.36845f
C567 VDD1.t1 B 0.265646f
C568 VDD1.t0 B 0.265646f
C569 VDD1.n1 B 3.16376f
C570 VP.t3 B 2.55467f
C571 VP.n0 B 0.971178f
C572 VP.n1 B 0.02037f
C573 VP.n2 B 0.040485f
C574 VP.n3 B 0.02037f
C575 VP.n4 B 0.037964f
C576 VP.t0 B 2.88041f
C577 VP.t1 B 2.86808f
C578 VP.n5 B 3.05073f
C579 VP.n6 B 1.24334f
C580 VP.t2 B 2.55467f
C581 VP.n7 B 0.971178f
C582 VP.n8 B 0.021657f
C583 VP.n9 B 0.032876f
C584 VP.n10 B 0.02037f
C585 VP.n11 B 0.02037f
C586 VP.n12 B 0.037964f
C587 VP.n13 B 0.040485f
C588 VP.n14 B 0.016467f
C589 VP.n15 B 0.02037f
C590 VP.n16 B 0.02037f
C591 VP.n17 B 0.02037f
C592 VP.n18 B 0.037964f
C593 VP.n19 B 0.037964f
C594 VP.n20 B 0.021657f
C595 VP.n21 B 0.032876f
C596 VP.n22 B 0.062397f
.ends

