* NGSPICE file created from diff_pair_sample_0933.ext - technology: sky130A

.subckt diff_pair_sample_0933 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=1.4274 ps=8.1 w=3.66 l=2.86
X1 VTAIL.t4 VN.t0 VDD2.t5 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=0.6039 ps=3.99 w=3.66 l=2.86
X2 VDD2.t4 VN.t1 VTAIL.t5 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0.6039 ps=3.99 w=3.66 l=2.86
X3 VTAIL.t3 VN.t2 VDD2.t3 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=0.6039 ps=3.99 w=3.66 l=2.86
X4 VTAIL.t8 VP.t1 VDD1.t4 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=0.6039 ps=3.99 w=3.66 l=2.86
X5 VDD1.t3 VP.t2 VTAIL.t10 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=1.4274 ps=8.1 w=3.66 l=2.86
X6 VDD2.t2 VN.t3 VTAIL.t0 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=1.4274 ps=8.1 w=3.66 l=2.86
X7 VTAIL.t9 VP.t3 VDD1.t2 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=0.6039 ps=3.99 w=3.66 l=2.86
X8 VDD2.t1 VN.t4 VTAIL.t1 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0.6039 ps=3.99 w=3.66 l=2.86
X9 B.t11 B.t9 B.t10 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0 ps=0 w=3.66 l=2.86
X10 B.t8 B.t6 B.t7 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0 ps=0 w=3.66 l=2.86
X11 VDD1.t1 VP.t4 VTAIL.t11 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0.6039 ps=3.99 w=3.66 l=2.86
X12 VDD2.t0 VN.t5 VTAIL.t2 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=0.6039 pd=3.99 as=1.4274 ps=8.1 w=3.66 l=2.86
X13 B.t5 B.t3 B.t4 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0 ps=0 w=3.66 l=2.86
X14 B.t2 B.t0 B.t1 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0 ps=0 w=3.66 l=2.86
X15 VDD1.t0 VP.t5 VTAIL.t6 w_n3522_n1700# sky130_fd_pr__pfet_01v8 ad=1.4274 pd=8.1 as=0.6039 ps=3.99 w=3.66 l=2.86
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n41 VP.n1 161.3
R8 VP.n40 VP.n39 161.3
R9 VP.n38 VP.n2 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n35 VP.n3 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n24 VP.n23 68.6047
R19 VP.n44 VP.n0 68.6047
R20 VP.n22 VP.n7 68.6047
R21 VP.n11 VP.t4 62.6986
R22 VP.n12 VP.n11 61.6686
R23 VP.n29 VP.n28 55.593
R24 VP.n40 VP.n2 55.593
R25 VP.n18 VP.n9 55.593
R26 VP.n24 VP.n22 43.4882
R27 VP.n23 VP.t5 30.8418
R28 VP.n34 VP.t3 30.8418
R29 VP.n0 VP.t2 30.8418
R30 VP.n7 VP.t0 30.8418
R31 VP.n12 VP.t1 30.8418
R32 VP.n28 VP.n27 25.5611
R33 VP.n41 VP.n40 25.5611
R34 VP.n19 VP.n18 25.5611
R35 VP.n27 VP.n6 24.5923
R36 VP.n29 VP.n4 24.5923
R37 VP.n33 VP.n4 24.5923
R38 VP.n36 VP.n35 24.5923
R39 VP.n36 VP.n2 24.5923
R40 VP.n42 VP.n41 24.5923
R41 VP.n20 VP.n19 24.5923
R42 VP.n14 VP.n13 24.5923
R43 VP.n14 VP.n9 24.5923
R44 VP.n23 VP.n6 21.6413
R45 VP.n42 VP.n0 21.6413
R46 VP.n20 VP.n7 21.6413
R47 VP.n34 VP.n33 12.2964
R48 VP.n35 VP.n34 12.2964
R49 VP.n13 VP.n12 12.2964
R50 VP.n11 VP.n10 5.42191
R51 VP.n22 VP.n21 0.354861
R52 VP.n25 VP.n24 0.354861
R53 VP.n44 VP.n43 0.354861
R54 VP VP.n44 0.267071
R55 VP.n15 VP.n10 0.189894
R56 VP.n16 VP.n15 0.189894
R57 VP.n17 VP.n16 0.189894
R58 VP.n17 VP.n8 0.189894
R59 VP.n21 VP.n8 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n5 0.189894
R62 VP.n30 VP.n5 0.189894
R63 VP.n31 VP.n30 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n32 VP.n3 0.189894
R66 VP.n37 VP.n3 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n39 VP.n38 0.189894
R69 VP.n39 VP.n1 0.189894
R70 VP.n43 VP.n1 0.189894
R71 VTAIL.n7 VTAIL.t0 115.602
R72 VTAIL.n11 VTAIL.t2 115.602
R73 VTAIL.n2 VTAIL.t10 115.602
R74 VTAIL.n10 VTAIL.t7 115.602
R75 VTAIL.n9 VTAIL.n8 106.721
R76 VTAIL.n6 VTAIL.n5 106.721
R77 VTAIL.n1 VTAIL.n0 106.721
R78 VTAIL.n4 VTAIL.n3 106.721
R79 VTAIL.n6 VTAIL.n4 21.0221
R80 VTAIL.n11 VTAIL.n10 18.2721
R81 VTAIL.n0 VTAIL.t5 8.88165
R82 VTAIL.n0 VTAIL.t3 8.88165
R83 VTAIL.n3 VTAIL.t6 8.88165
R84 VTAIL.n3 VTAIL.t9 8.88165
R85 VTAIL.n8 VTAIL.t11 8.88165
R86 VTAIL.n8 VTAIL.t8 8.88165
R87 VTAIL.n5 VTAIL.t1 8.88165
R88 VTAIL.n5 VTAIL.t4 8.88165
R89 VTAIL.n7 VTAIL.n6 2.7505
R90 VTAIL.n10 VTAIL.n9 2.7505
R91 VTAIL.n4 VTAIL.n2 2.7505
R92 VTAIL VTAIL.n11 2.00481
R93 VTAIL.n9 VTAIL.n7 1.84533
R94 VTAIL.n2 VTAIL.n1 1.84533
R95 VTAIL VTAIL.n1 0.74619
R96 VDD1 VDD1.t1 134.4
R97 VDD1.n1 VDD1.t0 134.287
R98 VDD1.n1 VDD1.n0 124.031
R99 VDD1.n3 VDD1.n2 123.4
R100 VDD1.n3 VDD1.n1 37.766
R101 VDD1.n2 VDD1.t4 8.88165
R102 VDD1.n2 VDD1.t5 8.88165
R103 VDD1.n0 VDD1.t2 8.88165
R104 VDD1.n0 VDD1.t3 8.88165
R105 VDD1 VDD1.n3 0.62981
R106 VN.n30 VN.n29 161.3
R107 VN.n28 VN.n17 161.3
R108 VN.n27 VN.n26 161.3
R109 VN.n25 VN.n18 161.3
R110 VN.n24 VN.n23 161.3
R111 VN.n22 VN.n19 161.3
R112 VN.n14 VN.n13 161.3
R113 VN.n12 VN.n1 161.3
R114 VN.n11 VN.n10 161.3
R115 VN.n9 VN.n2 161.3
R116 VN.n8 VN.n7 161.3
R117 VN.n6 VN.n3 161.3
R118 VN.n15 VN.n0 68.6047
R119 VN.n31 VN.n16 68.6047
R120 VN.n20 VN.t3 62.6988
R121 VN.n4 VN.t1 62.6988
R122 VN.n5 VN.n4 61.6686
R123 VN.n21 VN.n20 61.6686
R124 VN.n11 VN.n2 55.593
R125 VN.n27 VN.n18 55.593
R126 VN VN.n31 43.6534
R127 VN.n5 VN.t2 30.8418
R128 VN.n0 VN.t5 30.8418
R129 VN.n21 VN.t0 30.8418
R130 VN.n16 VN.t4 30.8418
R131 VN.n12 VN.n11 25.5611
R132 VN.n28 VN.n27 25.5611
R133 VN.n7 VN.n6 24.5923
R134 VN.n7 VN.n2 24.5923
R135 VN.n13 VN.n12 24.5923
R136 VN.n23 VN.n18 24.5923
R137 VN.n23 VN.n22 24.5923
R138 VN.n29 VN.n28 24.5923
R139 VN.n13 VN.n0 21.6413
R140 VN.n29 VN.n16 21.6413
R141 VN.n6 VN.n5 12.2964
R142 VN.n22 VN.n21 12.2964
R143 VN.n20 VN.n19 5.42195
R144 VN.n4 VN.n3 5.42195
R145 VN.n31 VN.n30 0.354861
R146 VN.n15 VN.n14 0.354861
R147 VN VN.n15 0.267071
R148 VN.n30 VN.n17 0.189894
R149 VN.n26 VN.n17 0.189894
R150 VN.n26 VN.n25 0.189894
R151 VN.n25 VN.n24 0.189894
R152 VN.n24 VN.n19 0.189894
R153 VN.n8 VN.n3 0.189894
R154 VN.n9 VN.n8 0.189894
R155 VN.n10 VN.n9 0.189894
R156 VN.n10 VN.n1 0.189894
R157 VN.n14 VN.n1 0.189894
R158 VDD2.n1 VDD2.t4 134.287
R159 VDD2.n2 VDD2.t1 132.28
R160 VDD2.n1 VDD2.n0 124.031
R161 VDD2 VDD2.n3 124.028
R162 VDD2.n2 VDD2.n1 35.808
R163 VDD2.n3 VDD2.t5 8.88165
R164 VDD2.n3 VDD2.t2 8.88165
R165 VDD2.n0 VDD2.t3 8.88165
R166 VDD2.n0 VDD2.t0 8.88165
R167 VDD2 VDD2.n2 2.12119
R168 B.n278 B.n97 585
R169 B.n277 B.n276 585
R170 B.n275 B.n98 585
R171 B.n274 B.n273 585
R172 B.n272 B.n99 585
R173 B.n271 B.n270 585
R174 B.n269 B.n100 585
R175 B.n268 B.n267 585
R176 B.n266 B.n101 585
R177 B.n265 B.n264 585
R178 B.n263 B.n102 585
R179 B.n262 B.n261 585
R180 B.n260 B.n103 585
R181 B.n259 B.n258 585
R182 B.n257 B.n104 585
R183 B.n256 B.n255 585
R184 B.n254 B.n105 585
R185 B.n252 B.n251 585
R186 B.n250 B.n108 585
R187 B.n249 B.n248 585
R188 B.n247 B.n109 585
R189 B.n246 B.n245 585
R190 B.n244 B.n110 585
R191 B.n243 B.n242 585
R192 B.n241 B.n111 585
R193 B.n240 B.n239 585
R194 B.n238 B.n112 585
R195 B.n237 B.n236 585
R196 B.n232 B.n113 585
R197 B.n231 B.n230 585
R198 B.n229 B.n114 585
R199 B.n228 B.n227 585
R200 B.n226 B.n115 585
R201 B.n225 B.n224 585
R202 B.n223 B.n116 585
R203 B.n222 B.n221 585
R204 B.n220 B.n117 585
R205 B.n219 B.n218 585
R206 B.n217 B.n118 585
R207 B.n216 B.n215 585
R208 B.n214 B.n119 585
R209 B.n213 B.n212 585
R210 B.n211 B.n120 585
R211 B.n210 B.n209 585
R212 B.n280 B.n279 585
R213 B.n281 B.n96 585
R214 B.n283 B.n282 585
R215 B.n284 B.n95 585
R216 B.n286 B.n285 585
R217 B.n287 B.n94 585
R218 B.n289 B.n288 585
R219 B.n290 B.n93 585
R220 B.n292 B.n291 585
R221 B.n293 B.n92 585
R222 B.n295 B.n294 585
R223 B.n296 B.n91 585
R224 B.n298 B.n297 585
R225 B.n299 B.n90 585
R226 B.n301 B.n300 585
R227 B.n302 B.n89 585
R228 B.n304 B.n303 585
R229 B.n305 B.n88 585
R230 B.n307 B.n306 585
R231 B.n308 B.n87 585
R232 B.n310 B.n309 585
R233 B.n311 B.n86 585
R234 B.n313 B.n312 585
R235 B.n314 B.n85 585
R236 B.n316 B.n315 585
R237 B.n317 B.n84 585
R238 B.n319 B.n318 585
R239 B.n320 B.n83 585
R240 B.n322 B.n321 585
R241 B.n323 B.n82 585
R242 B.n325 B.n324 585
R243 B.n326 B.n81 585
R244 B.n328 B.n327 585
R245 B.n329 B.n80 585
R246 B.n331 B.n330 585
R247 B.n332 B.n79 585
R248 B.n334 B.n333 585
R249 B.n335 B.n78 585
R250 B.n337 B.n336 585
R251 B.n338 B.n77 585
R252 B.n340 B.n339 585
R253 B.n341 B.n76 585
R254 B.n343 B.n342 585
R255 B.n344 B.n75 585
R256 B.n346 B.n345 585
R257 B.n347 B.n74 585
R258 B.n349 B.n348 585
R259 B.n350 B.n73 585
R260 B.n352 B.n351 585
R261 B.n353 B.n72 585
R262 B.n355 B.n354 585
R263 B.n356 B.n71 585
R264 B.n358 B.n357 585
R265 B.n359 B.n70 585
R266 B.n361 B.n360 585
R267 B.n362 B.n69 585
R268 B.n364 B.n363 585
R269 B.n365 B.n68 585
R270 B.n367 B.n366 585
R271 B.n368 B.n67 585
R272 B.n370 B.n369 585
R273 B.n371 B.n66 585
R274 B.n373 B.n372 585
R275 B.n374 B.n65 585
R276 B.n376 B.n375 585
R277 B.n377 B.n64 585
R278 B.n379 B.n378 585
R279 B.n380 B.n63 585
R280 B.n382 B.n381 585
R281 B.n383 B.n62 585
R282 B.n385 B.n384 585
R283 B.n386 B.n61 585
R284 B.n388 B.n387 585
R285 B.n389 B.n60 585
R286 B.n391 B.n390 585
R287 B.n392 B.n59 585
R288 B.n394 B.n393 585
R289 B.n395 B.n58 585
R290 B.n397 B.n396 585
R291 B.n398 B.n57 585
R292 B.n400 B.n399 585
R293 B.n401 B.n56 585
R294 B.n403 B.n402 585
R295 B.n404 B.n55 585
R296 B.n406 B.n405 585
R297 B.n407 B.n54 585
R298 B.n409 B.n408 585
R299 B.n410 B.n53 585
R300 B.n412 B.n411 585
R301 B.n413 B.n52 585
R302 B.n415 B.n414 585
R303 B.n416 B.n51 585
R304 B.n484 B.n483 585
R305 B.n482 B.n25 585
R306 B.n481 B.n480 585
R307 B.n479 B.n26 585
R308 B.n478 B.n477 585
R309 B.n476 B.n27 585
R310 B.n475 B.n474 585
R311 B.n473 B.n28 585
R312 B.n472 B.n471 585
R313 B.n470 B.n29 585
R314 B.n469 B.n468 585
R315 B.n467 B.n30 585
R316 B.n466 B.n465 585
R317 B.n464 B.n31 585
R318 B.n463 B.n462 585
R319 B.n461 B.n32 585
R320 B.n460 B.n459 585
R321 B.n457 B.n33 585
R322 B.n456 B.n455 585
R323 B.n454 B.n36 585
R324 B.n453 B.n452 585
R325 B.n451 B.n37 585
R326 B.n450 B.n449 585
R327 B.n448 B.n38 585
R328 B.n447 B.n446 585
R329 B.n445 B.n39 585
R330 B.n444 B.n443 585
R331 B.n442 B.n441 585
R332 B.n440 B.n43 585
R333 B.n439 B.n438 585
R334 B.n437 B.n44 585
R335 B.n436 B.n435 585
R336 B.n434 B.n45 585
R337 B.n433 B.n432 585
R338 B.n431 B.n46 585
R339 B.n430 B.n429 585
R340 B.n428 B.n47 585
R341 B.n427 B.n426 585
R342 B.n425 B.n48 585
R343 B.n424 B.n423 585
R344 B.n422 B.n49 585
R345 B.n421 B.n420 585
R346 B.n419 B.n50 585
R347 B.n418 B.n417 585
R348 B.n485 B.n24 585
R349 B.n487 B.n486 585
R350 B.n488 B.n23 585
R351 B.n490 B.n489 585
R352 B.n491 B.n22 585
R353 B.n493 B.n492 585
R354 B.n494 B.n21 585
R355 B.n496 B.n495 585
R356 B.n497 B.n20 585
R357 B.n499 B.n498 585
R358 B.n500 B.n19 585
R359 B.n502 B.n501 585
R360 B.n503 B.n18 585
R361 B.n505 B.n504 585
R362 B.n506 B.n17 585
R363 B.n508 B.n507 585
R364 B.n509 B.n16 585
R365 B.n511 B.n510 585
R366 B.n512 B.n15 585
R367 B.n514 B.n513 585
R368 B.n515 B.n14 585
R369 B.n517 B.n516 585
R370 B.n518 B.n13 585
R371 B.n520 B.n519 585
R372 B.n521 B.n12 585
R373 B.n523 B.n522 585
R374 B.n524 B.n11 585
R375 B.n526 B.n525 585
R376 B.n527 B.n10 585
R377 B.n529 B.n528 585
R378 B.n530 B.n9 585
R379 B.n532 B.n531 585
R380 B.n533 B.n8 585
R381 B.n535 B.n534 585
R382 B.n536 B.n7 585
R383 B.n538 B.n537 585
R384 B.n539 B.n6 585
R385 B.n541 B.n540 585
R386 B.n542 B.n5 585
R387 B.n544 B.n543 585
R388 B.n545 B.n4 585
R389 B.n547 B.n546 585
R390 B.n548 B.n3 585
R391 B.n550 B.n549 585
R392 B.n551 B.n0 585
R393 B.n2 B.n1 585
R394 B.n144 B.n143 585
R395 B.n145 B.n142 585
R396 B.n147 B.n146 585
R397 B.n148 B.n141 585
R398 B.n150 B.n149 585
R399 B.n151 B.n140 585
R400 B.n153 B.n152 585
R401 B.n154 B.n139 585
R402 B.n156 B.n155 585
R403 B.n157 B.n138 585
R404 B.n159 B.n158 585
R405 B.n160 B.n137 585
R406 B.n162 B.n161 585
R407 B.n163 B.n136 585
R408 B.n165 B.n164 585
R409 B.n166 B.n135 585
R410 B.n168 B.n167 585
R411 B.n169 B.n134 585
R412 B.n171 B.n170 585
R413 B.n172 B.n133 585
R414 B.n174 B.n173 585
R415 B.n175 B.n132 585
R416 B.n177 B.n176 585
R417 B.n178 B.n131 585
R418 B.n180 B.n179 585
R419 B.n181 B.n130 585
R420 B.n183 B.n182 585
R421 B.n184 B.n129 585
R422 B.n186 B.n185 585
R423 B.n187 B.n128 585
R424 B.n189 B.n188 585
R425 B.n190 B.n127 585
R426 B.n192 B.n191 585
R427 B.n193 B.n126 585
R428 B.n195 B.n194 585
R429 B.n196 B.n125 585
R430 B.n198 B.n197 585
R431 B.n199 B.n124 585
R432 B.n201 B.n200 585
R433 B.n202 B.n123 585
R434 B.n204 B.n203 585
R435 B.n205 B.n122 585
R436 B.n207 B.n206 585
R437 B.n208 B.n121 585
R438 B.n210 B.n121 502.111
R439 B.n280 B.n97 502.111
R440 B.n418 B.n51 502.111
R441 B.n485 B.n484 502.111
R442 B.n553 B.n552 256.663
R443 B.n233 B.t6 239.25
R444 B.n106 B.t0 239.25
R445 B.n40 B.t3 239.25
R446 B.n34 B.t9 239.25
R447 B.n552 B.n551 235.042
R448 B.n552 B.n2 235.042
R449 B.n106 B.t1 192.858
R450 B.n40 B.t5 192.858
R451 B.n233 B.t7 192.857
R452 B.n34 B.t11 192.857
R453 B.n211 B.n210 163.367
R454 B.n212 B.n211 163.367
R455 B.n212 B.n119 163.367
R456 B.n216 B.n119 163.367
R457 B.n217 B.n216 163.367
R458 B.n218 B.n217 163.367
R459 B.n218 B.n117 163.367
R460 B.n222 B.n117 163.367
R461 B.n223 B.n222 163.367
R462 B.n224 B.n223 163.367
R463 B.n224 B.n115 163.367
R464 B.n228 B.n115 163.367
R465 B.n229 B.n228 163.367
R466 B.n230 B.n229 163.367
R467 B.n230 B.n113 163.367
R468 B.n237 B.n113 163.367
R469 B.n238 B.n237 163.367
R470 B.n239 B.n238 163.367
R471 B.n239 B.n111 163.367
R472 B.n243 B.n111 163.367
R473 B.n244 B.n243 163.367
R474 B.n245 B.n244 163.367
R475 B.n245 B.n109 163.367
R476 B.n249 B.n109 163.367
R477 B.n250 B.n249 163.367
R478 B.n251 B.n250 163.367
R479 B.n251 B.n105 163.367
R480 B.n256 B.n105 163.367
R481 B.n257 B.n256 163.367
R482 B.n258 B.n257 163.367
R483 B.n258 B.n103 163.367
R484 B.n262 B.n103 163.367
R485 B.n263 B.n262 163.367
R486 B.n264 B.n263 163.367
R487 B.n264 B.n101 163.367
R488 B.n268 B.n101 163.367
R489 B.n269 B.n268 163.367
R490 B.n270 B.n269 163.367
R491 B.n270 B.n99 163.367
R492 B.n274 B.n99 163.367
R493 B.n275 B.n274 163.367
R494 B.n276 B.n275 163.367
R495 B.n276 B.n97 163.367
R496 B.n414 B.n51 163.367
R497 B.n414 B.n413 163.367
R498 B.n413 B.n412 163.367
R499 B.n412 B.n53 163.367
R500 B.n408 B.n53 163.367
R501 B.n408 B.n407 163.367
R502 B.n407 B.n406 163.367
R503 B.n406 B.n55 163.367
R504 B.n402 B.n55 163.367
R505 B.n402 B.n401 163.367
R506 B.n401 B.n400 163.367
R507 B.n400 B.n57 163.367
R508 B.n396 B.n57 163.367
R509 B.n396 B.n395 163.367
R510 B.n395 B.n394 163.367
R511 B.n394 B.n59 163.367
R512 B.n390 B.n59 163.367
R513 B.n390 B.n389 163.367
R514 B.n389 B.n388 163.367
R515 B.n388 B.n61 163.367
R516 B.n384 B.n61 163.367
R517 B.n384 B.n383 163.367
R518 B.n383 B.n382 163.367
R519 B.n382 B.n63 163.367
R520 B.n378 B.n63 163.367
R521 B.n378 B.n377 163.367
R522 B.n377 B.n376 163.367
R523 B.n376 B.n65 163.367
R524 B.n372 B.n65 163.367
R525 B.n372 B.n371 163.367
R526 B.n371 B.n370 163.367
R527 B.n370 B.n67 163.367
R528 B.n366 B.n67 163.367
R529 B.n366 B.n365 163.367
R530 B.n365 B.n364 163.367
R531 B.n364 B.n69 163.367
R532 B.n360 B.n69 163.367
R533 B.n360 B.n359 163.367
R534 B.n359 B.n358 163.367
R535 B.n358 B.n71 163.367
R536 B.n354 B.n71 163.367
R537 B.n354 B.n353 163.367
R538 B.n353 B.n352 163.367
R539 B.n352 B.n73 163.367
R540 B.n348 B.n73 163.367
R541 B.n348 B.n347 163.367
R542 B.n347 B.n346 163.367
R543 B.n346 B.n75 163.367
R544 B.n342 B.n75 163.367
R545 B.n342 B.n341 163.367
R546 B.n341 B.n340 163.367
R547 B.n340 B.n77 163.367
R548 B.n336 B.n77 163.367
R549 B.n336 B.n335 163.367
R550 B.n335 B.n334 163.367
R551 B.n334 B.n79 163.367
R552 B.n330 B.n79 163.367
R553 B.n330 B.n329 163.367
R554 B.n329 B.n328 163.367
R555 B.n328 B.n81 163.367
R556 B.n324 B.n81 163.367
R557 B.n324 B.n323 163.367
R558 B.n323 B.n322 163.367
R559 B.n322 B.n83 163.367
R560 B.n318 B.n83 163.367
R561 B.n318 B.n317 163.367
R562 B.n317 B.n316 163.367
R563 B.n316 B.n85 163.367
R564 B.n312 B.n85 163.367
R565 B.n312 B.n311 163.367
R566 B.n311 B.n310 163.367
R567 B.n310 B.n87 163.367
R568 B.n306 B.n87 163.367
R569 B.n306 B.n305 163.367
R570 B.n305 B.n304 163.367
R571 B.n304 B.n89 163.367
R572 B.n300 B.n89 163.367
R573 B.n300 B.n299 163.367
R574 B.n299 B.n298 163.367
R575 B.n298 B.n91 163.367
R576 B.n294 B.n91 163.367
R577 B.n294 B.n293 163.367
R578 B.n293 B.n292 163.367
R579 B.n292 B.n93 163.367
R580 B.n288 B.n93 163.367
R581 B.n288 B.n287 163.367
R582 B.n287 B.n286 163.367
R583 B.n286 B.n95 163.367
R584 B.n282 B.n95 163.367
R585 B.n282 B.n281 163.367
R586 B.n281 B.n280 163.367
R587 B.n484 B.n25 163.367
R588 B.n480 B.n25 163.367
R589 B.n480 B.n479 163.367
R590 B.n479 B.n478 163.367
R591 B.n478 B.n27 163.367
R592 B.n474 B.n27 163.367
R593 B.n474 B.n473 163.367
R594 B.n473 B.n472 163.367
R595 B.n472 B.n29 163.367
R596 B.n468 B.n29 163.367
R597 B.n468 B.n467 163.367
R598 B.n467 B.n466 163.367
R599 B.n466 B.n31 163.367
R600 B.n462 B.n31 163.367
R601 B.n462 B.n461 163.367
R602 B.n461 B.n460 163.367
R603 B.n460 B.n33 163.367
R604 B.n455 B.n33 163.367
R605 B.n455 B.n454 163.367
R606 B.n454 B.n453 163.367
R607 B.n453 B.n37 163.367
R608 B.n449 B.n37 163.367
R609 B.n449 B.n448 163.367
R610 B.n448 B.n447 163.367
R611 B.n447 B.n39 163.367
R612 B.n443 B.n39 163.367
R613 B.n443 B.n442 163.367
R614 B.n442 B.n43 163.367
R615 B.n438 B.n43 163.367
R616 B.n438 B.n437 163.367
R617 B.n437 B.n436 163.367
R618 B.n436 B.n45 163.367
R619 B.n432 B.n45 163.367
R620 B.n432 B.n431 163.367
R621 B.n431 B.n430 163.367
R622 B.n430 B.n47 163.367
R623 B.n426 B.n47 163.367
R624 B.n426 B.n425 163.367
R625 B.n425 B.n424 163.367
R626 B.n424 B.n49 163.367
R627 B.n420 B.n49 163.367
R628 B.n420 B.n419 163.367
R629 B.n419 B.n418 163.367
R630 B.n486 B.n485 163.367
R631 B.n486 B.n23 163.367
R632 B.n490 B.n23 163.367
R633 B.n491 B.n490 163.367
R634 B.n492 B.n491 163.367
R635 B.n492 B.n21 163.367
R636 B.n496 B.n21 163.367
R637 B.n497 B.n496 163.367
R638 B.n498 B.n497 163.367
R639 B.n498 B.n19 163.367
R640 B.n502 B.n19 163.367
R641 B.n503 B.n502 163.367
R642 B.n504 B.n503 163.367
R643 B.n504 B.n17 163.367
R644 B.n508 B.n17 163.367
R645 B.n509 B.n508 163.367
R646 B.n510 B.n509 163.367
R647 B.n510 B.n15 163.367
R648 B.n514 B.n15 163.367
R649 B.n515 B.n514 163.367
R650 B.n516 B.n515 163.367
R651 B.n516 B.n13 163.367
R652 B.n520 B.n13 163.367
R653 B.n521 B.n520 163.367
R654 B.n522 B.n521 163.367
R655 B.n522 B.n11 163.367
R656 B.n526 B.n11 163.367
R657 B.n527 B.n526 163.367
R658 B.n528 B.n527 163.367
R659 B.n528 B.n9 163.367
R660 B.n532 B.n9 163.367
R661 B.n533 B.n532 163.367
R662 B.n534 B.n533 163.367
R663 B.n534 B.n7 163.367
R664 B.n538 B.n7 163.367
R665 B.n539 B.n538 163.367
R666 B.n540 B.n539 163.367
R667 B.n540 B.n5 163.367
R668 B.n544 B.n5 163.367
R669 B.n545 B.n544 163.367
R670 B.n546 B.n545 163.367
R671 B.n546 B.n3 163.367
R672 B.n550 B.n3 163.367
R673 B.n551 B.n550 163.367
R674 B.n144 B.n2 163.367
R675 B.n145 B.n144 163.367
R676 B.n146 B.n145 163.367
R677 B.n146 B.n141 163.367
R678 B.n150 B.n141 163.367
R679 B.n151 B.n150 163.367
R680 B.n152 B.n151 163.367
R681 B.n152 B.n139 163.367
R682 B.n156 B.n139 163.367
R683 B.n157 B.n156 163.367
R684 B.n158 B.n157 163.367
R685 B.n158 B.n137 163.367
R686 B.n162 B.n137 163.367
R687 B.n163 B.n162 163.367
R688 B.n164 B.n163 163.367
R689 B.n164 B.n135 163.367
R690 B.n168 B.n135 163.367
R691 B.n169 B.n168 163.367
R692 B.n170 B.n169 163.367
R693 B.n170 B.n133 163.367
R694 B.n174 B.n133 163.367
R695 B.n175 B.n174 163.367
R696 B.n176 B.n175 163.367
R697 B.n176 B.n131 163.367
R698 B.n180 B.n131 163.367
R699 B.n181 B.n180 163.367
R700 B.n182 B.n181 163.367
R701 B.n182 B.n129 163.367
R702 B.n186 B.n129 163.367
R703 B.n187 B.n186 163.367
R704 B.n188 B.n187 163.367
R705 B.n188 B.n127 163.367
R706 B.n192 B.n127 163.367
R707 B.n193 B.n192 163.367
R708 B.n194 B.n193 163.367
R709 B.n194 B.n125 163.367
R710 B.n198 B.n125 163.367
R711 B.n199 B.n198 163.367
R712 B.n200 B.n199 163.367
R713 B.n200 B.n123 163.367
R714 B.n204 B.n123 163.367
R715 B.n205 B.n204 163.367
R716 B.n206 B.n205 163.367
R717 B.n206 B.n121 163.367
R718 B.n107 B.t2 130.993
R719 B.n41 B.t4 130.993
R720 B.n234 B.t8 130.989
R721 B.n35 B.t10 130.989
R722 B.n234 B.n233 61.8672
R723 B.n107 B.n106 61.8672
R724 B.n41 B.n40 61.8672
R725 B.n35 B.n34 61.8672
R726 B.n235 B.n234 59.5399
R727 B.n253 B.n107 59.5399
R728 B.n42 B.n41 59.5399
R729 B.n458 B.n35 59.5399
R730 B.n483 B.n24 32.6249
R731 B.n417 B.n416 32.6249
R732 B.n279 B.n278 32.6249
R733 B.n209 B.n208 32.6249
R734 B B.n553 18.0485
R735 B.n487 B.n24 10.6151
R736 B.n488 B.n487 10.6151
R737 B.n489 B.n488 10.6151
R738 B.n489 B.n22 10.6151
R739 B.n493 B.n22 10.6151
R740 B.n494 B.n493 10.6151
R741 B.n495 B.n494 10.6151
R742 B.n495 B.n20 10.6151
R743 B.n499 B.n20 10.6151
R744 B.n500 B.n499 10.6151
R745 B.n501 B.n500 10.6151
R746 B.n501 B.n18 10.6151
R747 B.n505 B.n18 10.6151
R748 B.n506 B.n505 10.6151
R749 B.n507 B.n506 10.6151
R750 B.n507 B.n16 10.6151
R751 B.n511 B.n16 10.6151
R752 B.n512 B.n511 10.6151
R753 B.n513 B.n512 10.6151
R754 B.n513 B.n14 10.6151
R755 B.n517 B.n14 10.6151
R756 B.n518 B.n517 10.6151
R757 B.n519 B.n518 10.6151
R758 B.n519 B.n12 10.6151
R759 B.n523 B.n12 10.6151
R760 B.n524 B.n523 10.6151
R761 B.n525 B.n524 10.6151
R762 B.n525 B.n10 10.6151
R763 B.n529 B.n10 10.6151
R764 B.n530 B.n529 10.6151
R765 B.n531 B.n530 10.6151
R766 B.n531 B.n8 10.6151
R767 B.n535 B.n8 10.6151
R768 B.n536 B.n535 10.6151
R769 B.n537 B.n536 10.6151
R770 B.n537 B.n6 10.6151
R771 B.n541 B.n6 10.6151
R772 B.n542 B.n541 10.6151
R773 B.n543 B.n542 10.6151
R774 B.n543 B.n4 10.6151
R775 B.n547 B.n4 10.6151
R776 B.n548 B.n547 10.6151
R777 B.n549 B.n548 10.6151
R778 B.n549 B.n0 10.6151
R779 B.n483 B.n482 10.6151
R780 B.n482 B.n481 10.6151
R781 B.n481 B.n26 10.6151
R782 B.n477 B.n26 10.6151
R783 B.n477 B.n476 10.6151
R784 B.n476 B.n475 10.6151
R785 B.n475 B.n28 10.6151
R786 B.n471 B.n28 10.6151
R787 B.n471 B.n470 10.6151
R788 B.n470 B.n469 10.6151
R789 B.n469 B.n30 10.6151
R790 B.n465 B.n30 10.6151
R791 B.n465 B.n464 10.6151
R792 B.n464 B.n463 10.6151
R793 B.n463 B.n32 10.6151
R794 B.n459 B.n32 10.6151
R795 B.n457 B.n456 10.6151
R796 B.n456 B.n36 10.6151
R797 B.n452 B.n36 10.6151
R798 B.n452 B.n451 10.6151
R799 B.n451 B.n450 10.6151
R800 B.n450 B.n38 10.6151
R801 B.n446 B.n38 10.6151
R802 B.n446 B.n445 10.6151
R803 B.n445 B.n444 10.6151
R804 B.n441 B.n440 10.6151
R805 B.n440 B.n439 10.6151
R806 B.n439 B.n44 10.6151
R807 B.n435 B.n44 10.6151
R808 B.n435 B.n434 10.6151
R809 B.n434 B.n433 10.6151
R810 B.n433 B.n46 10.6151
R811 B.n429 B.n46 10.6151
R812 B.n429 B.n428 10.6151
R813 B.n428 B.n427 10.6151
R814 B.n427 B.n48 10.6151
R815 B.n423 B.n48 10.6151
R816 B.n423 B.n422 10.6151
R817 B.n422 B.n421 10.6151
R818 B.n421 B.n50 10.6151
R819 B.n417 B.n50 10.6151
R820 B.n416 B.n415 10.6151
R821 B.n415 B.n52 10.6151
R822 B.n411 B.n52 10.6151
R823 B.n411 B.n410 10.6151
R824 B.n410 B.n409 10.6151
R825 B.n409 B.n54 10.6151
R826 B.n405 B.n54 10.6151
R827 B.n405 B.n404 10.6151
R828 B.n404 B.n403 10.6151
R829 B.n403 B.n56 10.6151
R830 B.n399 B.n56 10.6151
R831 B.n399 B.n398 10.6151
R832 B.n398 B.n397 10.6151
R833 B.n397 B.n58 10.6151
R834 B.n393 B.n58 10.6151
R835 B.n393 B.n392 10.6151
R836 B.n392 B.n391 10.6151
R837 B.n391 B.n60 10.6151
R838 B.n387 B.n60 10.6151
R839 B.n387 B.n386 10.6151
R840 B.n386 B.n385 10.6151
R841 B.n385 B.n62 10.6151
R842 B.n381 B.n62 10.6151
R843 B.n381 B.n380 10.6151
R844 B.n380 B.n379 10.6151
R845 B.n379 B.n64 10.6151
R846 B.n375 B.n64 10.6151
R847 B.n375 B.n374 10.6151
R848 B.n374 B.n373 10.6151
R849 B.n373 B.n66 10.6151
R850 B.n369 B.n66 10.6151
R851 B.n369 B.n368 10.6151
R852 B.n368 B.n367 10.6151
R853 B.n367 B.n68 10.6151
R854 B.n363 B.n68 10.6151
R855 B.n363 B.n362 10.6151
R856 B.n362 B.n361 10.6151
R857 B.n361 B.n70 10.6151
R858 B.n357 B.n70 10.6151
R859 B.n357 B.n356 10.6151
R860 B.n356 B.n355 10.6151
R861 B.n355 B.n72 10.6151
R862 B.n351 B.n72 10.6151
R863 B.n351 B.n350 10.6151
R864 B.n350 B.n349 10.6151
R865 B.n349 B.n74 10.6151
R866 B.n345 B.n74 10.6151
R867 B.n345 B.n344 10.6151
R868 B.n344 B.n343 10.6151
R869 B.n343 B.n76 10.6151
R870 B.n339 B.n76 10.6151
R871 B.n339 B.n338 10.6151
R872 B.n338 B.n337 10.6151
R873 B.n337 B.n78 10.6151
R874 B.n333 B.n78 10.6151
R875 B.n333 B.n332 10.6151
R876 B.n332 B.n331 10.6151
R877 B.n331 B.n80 10.6151
R878 B.n327 B.n80 10.6151
R879 B.n327 B.n326 10.6151
R880 B.n326 B.n325 10.6151
R881 B.n325 B.n82 10.6151
R882 B.n321 B.n82 10.6151
R883 B.n321 B.n320 10.6151
R884 B.n320 B.n319 10.6151
R885 B.n319 B.n84 10.6151
R886 B.n315 B.n84 10.6151
R887 B.n315 B.n314 10.6151
R888 B.n314 B.n313 10.6151
R889 B.n313 B.n86 10.6151
R890 B.n309 B.n86 10.6151
R891 B.n309 B.n308 10.6151
R892 B.n308 B.n307 10.6151
R893 B.n307 B.n88 10.6151
R894 B.n303 B.n88 10.6151
R895 B.n303 B.n302 10.6151
R896 B.n302 B.n301 10.6151
R897 B.n301 B.n90 10.6151
R898 B.n297 B.n90 10.6151
R899 B.n297 B.n296 10.6151
R900 B.n296 B.n295 10.6151
R901 B.n295 B.n92 10.6151
R902 B.n291 B.n92 10.6151
R903 B.n291 B.n290 10.6151
R904 B.n290 B.n289 10.6151
R905 B.n289 B.n94 10.6151
R906 B.n285 B.n94 10.6151
R907 B.n285 B.n284 10.6151
R908 B.n284 B.n283 10.6151
R909 B.n283 B.n96 10.6151
R910 B.n279 B.n96 10.6151
R911 B.n143 B.n1 10.6151
R912 B.n143 B.n142 10.6151
R913 B.n147 B.n142 10.6151
R914 B.n148 B.n147 10.6151
R915 B.n149 B.n148 10.6151
R916 B.n149 B.n140 10.6151
R917 B.n153 B.n140 10.6151
R918 B.n154 B.n153 10.6151
R919 B.n155 B.n154 10.6151
R920 B.n155 B.n138 10.6151
R921 B.n159 B.n138 10.6151
R922 B.n160 B.n159 10.6151
R923 B.n161 B.n160 10.6151
R924 B.n161 B.n136 10.6151
R925 B.n165 B.n136 10.6151
R926 B.n166 B.n165 10.6151
R927 B.n167 B.n166 10.6151
R928 B.n167 B.n134 10.6151
R929 B.n171 B.n134 10.6151
R930 B.n172 B.n171 10.6151
R931 B.n173 B.n172 10.6151
R932 B.n173 B.n132 10.6151
R933 B.n177 B.n132 10.6151
R934 B.n178 B.n177 10.6151
R935 B.n179 B.n178 10.6151
R936 B.n179 B.n130 10.6151
R937 B.n183 B.n130 10.6151
R938 B.n184 B.n183 10.6151
R939 B.n185 B.n184 10.6151
R940 B.n185 B.n128 10.6151
R941 B.n189 B.n128 10.6151
R942 B.n190 B.n189 10.6151
R943 B.n191 B.n190 10.6151
R944 B.n191 B.n126 10.6151
R945 B.n195 B.n126 10.6151
R946 B.n196 B.n195 10.6151
R947 B.n197 B.n196 10.6151
R948 B.n197 B.n124 10.6151
R949 B.n201 B.n124 10.6151
R950 B.n202 B.n201 10.6151
R951 B.n203 B.n202 10.6151
R952 B.n203 B.n122 10.6151
R953 B.n207 B.n122 10.6151
R954 B.n208 B.n207 10.6151
R955 B.n209 B.n120 10.6151
R956 B.n213 B.n120 10.6151
R957 B.n214 B.n213 10.6151
R958 B.n215 B.n214 10.6151
R959 B.n215 B.n118 10.6151
R960 B.n219 B.n118 10.6151
R961 B.n220 B.n219 10.6151
R962 B.n221 B.n220 10.6151
R963 B.n221 B.n116 10.6151
R964 B.n225 B.n116 10.6151
R965 B.n226 B.n225 10.6151
R966 B.n227 B.n226 10.6151
R967 B.n227 B.n114 10.6151
R968 B.n231 B.n114 10.6151
R969 B.n232 B.n231 10.6151
R970 B.n236 B.n232 10.6151
R971 B.n240 B.n112 10.6151
R972 B.n241 B.n240 10.6151
R973 B.n242 B.n241 10.6151
R974 B.n242 B.n110 10.6151
R975 B.n246 B.n110 10.6151
R976 B.n247 B.n246 10.6151
R977 B.n248 B.n247 10.6151
R978 B.n248 B.n108 10.6151
R979 B.n252 B.n108 10.6151
R980 B.n255 B.n254 10.6151
R981 B.n255 B.n104 10.6151
R982 B.n259 B.n104 10.6151
R983 B.n260 B.n259 10.6151
R984 B.n261 B.n260 10.6151
R985 B.n261 B.n102 10.6151
R986 B.n265 B.n102 10.6151
R987 B.n266 B.n265 10.6151
R988 B.n267 B.n266 10.6151
R989 B.n267 B.n100 10.6151
R990 B.n271 B.n100 10.6151
R991 B.n272 B.n271 10.6151
R992 B.n273 B.n272 10.6151
R993 B.n273 B.n98 10.6151
R994 B.n277 B.n98 10.6151
R995 B.n278 B.n277 10.6151
R996 B.n459 B.n458 9.36635
R997 B.n441 B.n42 9.36635
R998 B.n236 B.n235 9.36635
R999 B.n254 B.n253 9.36635
R1000 B.n553 B.n0 8.11757
R1001 B.n553 B.n1 8.11757
R1002 B.n458 B.n457 1.24928
R1003 B.n444 B.n42 1.24928
R1004 B.n235 B.n112 1.24928
R1005 B.n253 B.n252 1.24928
C0 VDD1 VP 2.68494f
C1 VDD2 VTAIL 4.92179f
C2 VDD1 w_n3522_n1700# 1.77637f
C3 VN VDD1 0.156008f
C4 VDD1 B 1.49786f
C5 VP w_n3522_n1700# 7.03771f
C6 VN VP 5.63895f
C7 VDD2 VDD1 1.50788f
C8 VN w_n3522_n1700# 6.58298f
C9 B VP 1.90439f
C10 B w_n3522_n1700# 7.72091f
C11 VN B 1.1419f
C12 VTAIL VDD1 4.86718f
C13 VDD2 VP 0.485267f
C14 VDD2 w_n3522_n1700# 1.86932f
C15 VDD2 VN 2.3582f
C16 VTAIL VP 3.16927f
C17 VDD2 B 1.57837f
C18 VTAIL w_n3522_n1700# 1.82257f
C19 VTAIL VN 3.15512f
C20 VTAIL B 1.84988f
C21 VDD2 VSUBS 1.386413f
C22 VDD1 VSUBS 1.885157f
C23 VTAIL VSUBS 0.594167f
C24 VN VSUBS 5.927f
C25 VP VSUBS 2.622928f
C26 B VSUBS 3.944643f
C27 w_n3522_n1700# VSUBS 75.525795f
C28 B.n0 VSUBS 0.006332f
C29 B.n1 VSUBS 0.006332f
C30 B.n2 VSUBS 0.009365f
C31 B.n3 VSUBS 0.007176f
C32 B.n4 VSUBS 0.007176f
C33 B.n5 VSUBS 0.007176f
C34 B.n6 VSUBS 0.007176f
C35 B.n7 VSUBS 0.007176f
C36 B.n8 VSUBS 0.007176f
C37 B.n9 VSUBS 0.007176f
C38 B.n10 VSUBS 0.007176f
C39 B.n11 VSUBS 0.007176f
C40 B.n12 VSUBS 0.007176f
C41 B.n13 VSUBS 0.007176f
C42 B.n14 VSUBS 0.007176f
C43 B.n15 VSUBS 0.007176f
C44 B.n16 VSUBS 0.007176f
C45 B.n17 VSUBS 0.007176f
C46 B.n18 VSUBS 0.007176f
C47 B.n19 VSUBS 0.007176f
C48 B.n20 VSUBS 0.007176f
C49 B.n21 VSUBS 0.007176f
C50 B.n22 VSUBS 0.007176f
C51 B.n23 VSUBS 0.007176f
C52 B.n24 VSUBS 0.01619f
C53 B.n25 VSUBS 0.007176f
C54 B.n26 VSUBS 0.007176f
C55 B.n27 VSUBS 0.007176f
C56 B.n28 VSUBS 0.007176f
C57 B.n29 VSUBS 0.007176f
C58 B.n30 VSUBS 0.007176f
C59 B.n31 VSUBS 0.007176f
C60 B.n32 VSUBS 0.007176f
C61 B.n33 VSUBS 0.007176f
C62 B.t10 VSUBS 0.095754f
C63 B.t11 VSUBS 0.115164f
C64 B.t9 VSUBS 0.519724f
C65 B.n34 VSUBS 0.092955f
C66 B.n35 VSUBS 0.070742f
C67 B.n36 VSUBS 0.007176f
C68 B.n37 VSUBS 0.007176f
C69 B.n38 VSUBS 0.007176f
C70 B.n39 VSUBS 0.007176f
C71 B.t4 VSUBS 0.095754f
C72 B.t5 VSUBS 0.115164f
C73 B.t3 VSUBS 0.519724f
C74 B.n40 VSUBS 0.092955f
C75 B.n41 VSUBS 0.070742f
C76 B.n42 VSUBS 0.016627f
C77 B.n43 VSUBS 0.007176f
C78 B.n44 VSUBS 0.007176f
C79 B.n45 VSUBS 0.007176f
C80 B.n46 VSUBS 0.007176f
C81 B.n47 VSUBS 0.007176f
C82 B.n48 VSUBS 0.007176f
C83 B.n49 VSUBS 0.007176f
C84 B.n50 VSUBS 0.007176f
C85 B.n51 VSUBS 0.01619f
C86 B.n52 VSUBS 0.007176f
C87 B.n53 VSUBS 0.007176f
C88 B.n54 VSUBS 0.007176f
C89 B.n55 VSUBS 0.007176f
C90 B.n56 VSUBS 0.007176f
C91 B.n57 VSUBS 0.007176f
C92 B.n58 VSUBS 0.007176f
C93 B.n59 VSUBS 0.007176f
C94 B.n60 VSUBS 0.007176f
C95 B.n61 VSUBS 0.007176f
C96 B.n62 VSUBS 0.007176f
C97 B.n63 VSUBS 0.007176f
C98 B.n64 VSUBS 0.007176f
C99 B.n65 VSUBS 0.007176f
C100 B.n66 VSUBS 0.007176f
C101 B.n67 VSUBS 0.007176f
C102 B.n68 VSUBS 0.007176f
C103 B.n69 VSUBS 0.007176f
C104 B.n70 VSUBS 0.007176f
C105 B.n71 VSUBS 0.007176f
C106 B.n72 VSUBS 0.007176f
C107 B.n73 VSUBS 0.007176f
C108 B.n74 VSUBS 0.007176f
C109 B.n75 VSUBS 0.007176f
C110 B.n76 VSUBS 0.007176f
C111 B.n77 VSUBS 0.007176f
C112 B.n78 VSUBS 0.007176f
C113 B.n79 VSUBS 0.007176f
C114 B.n80 VSUBS 0.007176f
C115 B.n81 VSUBS 0.007176f
C116 B.n82 VSUBS 0.007176f
C117 B.n83 VSUBS 0.007176f
C118 B.n84 VSUBS 0.007176f
C119 B.n85 VSUBS 0.007176f
C120 B.n86 VSUBS 0.007176f
C121 B.n87 VSUBS 0.007176f
C122 B.n88 VSUBS 0.007176f
C123 B.n89 VSUBS 0.007176f
C124 B.n90 VSUBS 0.007176f
C125 B.n91 VSUBS 0.007176f
C126 B.n92 VSUBS 0.007176f
C127 B.n93 VSUBS 0.007176f
C128 B.n94 VSUBS 0.007176f
C129 B.n95 VSUBS 0.007176f
C130 B.n96 VSUBS 0.007176f
C131 B.n97 VSUBS 0.01737f
C132 B.n98 VSUBS 0.007176f
C133 B.n99 VSUBS 0.007176f
C134 B.n100 VSUBS 0.007176f
C135 B.n101 VSUBS 0.007176f
C136 B.n102 VSUBS 0.007176f
C137 B.n103 VSUBS 0.007176f
C138 B.n104 VSUBS 0.007176f
C139 B.n105 VSUBS 0.007176f
C140 B.t2 VSUBS 0.095754f
C141 B.t1 VSUBS 0.115164f
C142 B.t0 VSUBS 0.519724f
C143 B.n106 VSUBS 0.092955f
C144 B.n107 VSUBS 0.070742f
C145 B.n108 VSUBS 0.007176f
C146 B.n109 VSUBS 0.007176f
C147 B.n110 VSUBS 0.007176f
C148 B.n111 VSUBS 0.007176f
C149 B.n112 VSUBS 0.00401f
C150 B.n113 VSUBS 0.007176f
C151 B.n114 VSUBS 0.007176f
C152 B.n115 VSUBS 0.007176f
C153 B.n116 VSUBS 0.007176f
C154 B.n117 VSUBS 0.007176f
C155 B.n118 VSUBS 0.007176f
C156 B.n119 VSUBS 0.007176f
C157 B.n120 VSUBS 0.007176f
C158 B.n121 VSUBS 0.01619f
C159 B.n122 VSUBS 0.007176f
C160 B.n123 VSUBS 0.007176f
C161 B.n124 VSUBS 0.007176f
C162 B.n125 VSUBS 0.007176f
C163 B.n126 VSUBS 0.007176f
C164 B.n127 VSUBS 0.007176f
C165 B.n128 VSUBS 0.007176f
C166 B.n129 VSUBS 0.007176f
C167 B.n130 VSUBS 0.007176f
C168 B.n131 VSUBS 0.007176f
C169 B.n132 VSUBS 0.007176f
C170 B.n133 VSUBS 0.007176f
C171 B.n134 VSUBS 0.007176f
C172 B.n135 VSUBS 0.007176f
C173 B.n136 VSUBS 0.007176f
C174 B.n137 VSUBS 0.007176f
C175 B.n138 VSUBS 0.007176f
C176 B.n139 VSUBS 0.007176f
C177 B.n140 VSUBS 0.007176f
C178 B.n141 VSUBS 0.007176f
C179 B.n142 VSUBS 0.007176f
C180 B.n143 VSUBS 0.007176f
C181 B.n144 VSUBS 0.007176f
C182 B.n145 VSUBS 0.007176f
C183 B.n146 VSUBS 0.007176f
C184 B.n147 VSUBS 0.007176f
C185 B.n148 VSUBS 0.007176f
C186 B.n149 VSUBS 0.007176f
C187 B.n150 VSUBS 0.007176f
C188 B.n151 VSUBS 0.007176f
C189 B.n152 VSUBS 0.007176f
C190 B.n153 VSUBS 0.007176f
C191 B.n154 VSUBS 0.007176f
C192 B.n155 VSUBS 0.007176f
C193 B.n156 VSUBS 0.007176f
C194 B.n157 VSUBS 0.007176f
C195 B.n158 VSUBS 0.007176f
C196 B.n159 VSUBS 0.007176f
C197 B.n160 VSUBS 0.007176f
C198 B.n161 VSUBS 0.007176f
C199 B.n162 VSUBS 0.007176f
C200 B.n163 VSUBS 0.007176f
C201 B.n164 VSUBS 0.007176f
C202 B.n165 VSUBS 0.007176f
C203 B.n166 VSUBS 0.007176f
C204 B.n167 VSUBS 0.007176f
C205 B.n168 VSUBS 0.007176f
C206 B.n169 VSUBS 0.007176f
C207 B.n170 VSUBS 0.007176f
C208 B.n171 VSUBS 0.007176f
C209 B.n172 VSUBS 0.007176f
C210 B.n173 VSUBS 0.007176f
C211 B.n174 VSUBS 0.007176f
C212 B.n175 VSUBS 0.007176f
C213 B.n176 VSUBS 0.007176f
C214 B.n177 VSUBS 0.007176f
C215 B.n178 VSUBS 0.007176f
C216 B.n179 VSUBS 0.007176f
C217 B.n180 VSUBS 0.007176f
C218 B.n181 VSUBS 0.007176f
C219 B.n182 VSUBS 0.007176f
C220 B.n183 VSUBS 0.007176f
C221 B.n184 VSUBS 0.007176f
C222 B.n185 VSUBS 0.007176f
C223 B.n186 VSUBS 0.007176f
C224 B.n187 VSUBS 0.007176f
C225 B.n188 VSUBS 0.007176f
C226 B.n189 VSUBS 0.007176f
C227 B.n190 VSUBS 0.007176f
C228 B.n191 VSUBS 0.007176f
C229 B.n192 VSUBS 0.007176f
C230 B.n193 VSUBS 0.007176f
C231 B.n194 VSUBS 0.007176f
C232 B.n195 VSUBS 0.007176f
C233 B.n196 VSUBS 0.007176f
C234 B.n197 VSUBS 0.007176f
C235 B.n198 VSUBS 0.007176f
C236 B.n199 VSUBS 0.007176f
C237 B.n200 VSUBS 0.007176f
C238 B.n201 VSUBS 0.007176f
C239 B.n202 VSUBS 0.007176f
C240 B.n203 VSUBS 0.007176f
C241 B.n204 VSUBS 0.007176f
C242 B.n205 VSUBS 0.007176f
C243 B.n206 VSUBS 0.007176f
C244 B.n207 VSUBS 0.007176f
C245 B.n208 VSUBS 0.01619f
C246 B.n209 VSUBS 0.01737f
C247 B.n210 VSUBS 0.01737f
C248 B.n211 VSUBS 0.007176f
C249 B.n212 VSUBS 0.007176f
C250 B.n213 VSUBS 0.007176f
C251 B.n214 VSUBS 0.007176f
C252 B.n215 VSUBS 0.007176f
C253 B.n216 VSUBS 0.007176f
C254 B.n217 VSUBS 0.007176f
C255 B.n218 VSUBS 0.007176f
C256 B.n219 VSUBS 0.007176f
C257 B.n220 VSUBS 0.007176f
C258 B.n221 VSUBS 0.007176f
C259 B.n222 VSUBS 0.007176f
C260 B.n223 VSUBS 0.007176f
C261 B.n224 VSUBS 0.007176f
C262 B.n225 VSUBS 0.007176f
C263 B.n226 VSUBS 0.007176f
C264 B.n227 VSUBS 0.007176f
C265 B.n228 VSUBS 0.007176f
C266 B.n229 VSUBS 0.007176f
C267 B.n230 VSUBS 0.007176f
C268 B.n231 VSUBS 0.007176f
C269 B.n232 VSUBS 0.007176f
C270 B.t8 VSUBS 0.095754f
C271 B.t7 VSUBS 0.115164f
C272 B.t6 VSUBS 0.519724f
C273 B.n233 VSUBS 0.092955f
C274 B.n234 VSUBS 0.070742f
C275 B.n235 VSUBS 0.016627f
C276 B.n236 VSUBS 0.006754f
C277 B.n237 VSUBS 0.007176f
C278 B.n238 VSUBS 0.007176f
C279 B.n239 VSUBS 0.007176f
C280 B.n240 VSUBS 0.007176f
C281 B.n241 VSUBS 0.007176f
C282 B.n242 VSUBS 0.007176f
C283 B.n243 VSUBS 0.007176f
C284 B.n244 VSUBS 0.007176f
C285 B.n245 VSUBS 0.007176f
C286 B.n246 VSUBS 0.007176f
C287 B.n247 VSUBS 0.007176f
C288 B.n248 VSUBS 0.007176f
C289 B.n249 VSUBS 0.007176f
C290 B.n250 VSUBS 0.007176f
C291 B.n251 VSUBS 0.007176f
C292 B.n252 VSUBS 0.00401f
C293 B.n253 VSUBS 0.016627f
C294 B.n254 VSUBS 0.006754f
C295 B.n255 VSUBS 0.007176f
C296 B.n256 VSUBS 0.007176f
C297 B.n257 VSUBS 0.007176f
C298 B.n258 VSUBS 0.007176f
C299 B.n259 VSUBS 0.007176f
C300 B.n260 VSUBS 0.007176f
C301 B.n261 VSUBS 0.007176f
C302 B.n262 VSUBS 0.007176f
C303 B.n263 VSUBS 0.007176f
C304 B.n264 VSUBS 0.007176f
C305 B.n265 VSUBS 0.007176f
C306 B.n266 VSUBS 0.007176f
C307 B.n267 VSUBS 0.007176f
C308 B.n268 VSUBS 0.007176f
C309 B.n269 VSUBS 0.007176f
C310 B.n270 VSUBS 0.007176f
C311 B.n271 VSUBS 0.007176f
C312 B.n272 VSUBS 0.007176f
C313 B.n273 VSUBS 0.007176f
C314 B.n274 VSUBS 0.007176f
C315 B.n275 VSUBS 0.007176f
C316 B.n276 VSUBS 0.007176f
C317 B.n277 VSUBS 0.007176f
C318 B.n278 VSUBS 0.016521f
C319 B.n279 VSUBS 0.017039f
C320 B.n280 VSUBS 0.01619f
C321 B.n281 VSUBS 0.007176f
C322 B.n282 VSUBS 0.007176f
C323 B.n283 VSUBS 0.007176f
C324 B.n284 VSUBS 0.007176f
C325 B.n285 VSUBS 0.007176f
C326 B.n286 VSUBS 0.007176f
C327 B.n287 VSUBS 0.007176f
C328 B.n288 VSUBS 0.007176f
C329 B.n289 VSUBS 0.007176f
C330 B.n290 VSUBS 0.007176f
C331 B.n291 VSUBS 0.007176f
C332 B.n292 VSUBS 0.007176f
C333 B.n293 VSUBS 0.007176f
C334 B.n294 VSUBS 0.007176f
C335 B.n295 VSUBS 0.007176f
C336 B.n296 VSUBS 0.007176f
C337 B.n297 VSUBS 0.007176f
C338 B.n298 VSUBS 0.007176f
C339 B.n299 VSUBS 0.007176f
C340 B.n300 VSUBS 0.007176f
C341 B.n301 VSUBS 0.007176f
C342 B.n302 VSUBS 0.007176f
C343 B.n303 VSUBS 0.007176f
C344 B.n304 VSUBS 0.007176f
C345 B.n305 VSUBS 0.007176f
C346 B.n306 VSUBS 0.007176f
C347 B.n307 VSUBS 0.007176f
C348 B.n308 VSUBS 0.007176f
C349 B.n309 VSUBS 0.007176f
C350 B.n310 VSUBS 0.007176f
C351 B.n311 VSUBS 0.007176f
C352 B.n312 VSUBS 0.007176f
C353 B.n313 VSUBS 0.007176f
C354 B.n314 VSUBS 0.007176f
C355 B.n315 VSUBS 0.007176f
C356 B.n316 VSUBS 0.007176f
C357 B.n317 VSUBS 0.007176f
C358 B.n318 VSUBS 0.007176f
C359 B.n319 VSUBS 0.007176f
C360 B.n320 VSUBS 0.007176f
C361 B.n321 VSUBS 0.007176f
C362 B.n322 VSUBS 0.007176f
C363 B.n323 VSUBS 0.007176f
C364 B.n324 VSUBS 0.007176f
C365 B.n325 VSUBS 0.007176f
C366 B.n326 VSUBS 0.007176f
C367 B.n327 VSUBS 0.007176f
C368 B.n328 VSUBS 0.007176f
C369 B.n329 VSUBS 0.007176f
C370 B.n330 VSUBS 0.007176f
C371 B.n331 VSUBS 0.007176f
C372 B.n332 VSUBS 0.007176f
C373 B.n333 VSUBS 0.007176f
C374 B.n334 VSUBS 0.007176f
C375 B.n335 VSUBS 0.007176f
C376 B.n336 VSUBS 0.007176f
C377 B.n337 VSUBS 0.007176f
C378 B.n338 VSUBS 0.007176f
C379 B.n339 VSUBS 0.007176f
C380 B.n340 VSUBS 0.007176f
C381 B.n341 VSUBS 0.007176f
C382 B.n342 VSUBS 0.007176f
C383 B.n343 VSUBS 0.007176f
C384 B.n344 VSUBS 0.007176f
C385 B.n345 VSUBS 0.007176f
C386 B.n346 VSUBS 0.007176f
C387 B.n347 VSUBS 0.007176f
C388 B.n348 VSUBS 0.007176f
C389 B.n349 VSUBS 0.007176f
C390 B.n350 VSUBS 0.007176f
C391 B.n351 VSUBS 0.007176f
C392 B.n352 VSUBS 0.007176f
C393 B.n353 VSUBS 0.007176f
C394 B.n354 VSUBS 0.007176f
C395 B.n355 VSUBS 0.007176f
C396 B.n356 VSUBS 0.007176f
C397 B.n357 VSUBS 0.007176f
C398 B.n358 VSUBS 0.007176f
C399 B.n359 VSUBS 0.007176f
C400 B.n360 VSUBS 0.007176f
C401 B.n361 VSUBS 0.007176f
C402 B.n362 VSUBS 0.007176f
C403 B.n363 VSUBS 0.007176f
C404 B.n364 VSUBS 0.007176f
C405 B.n365 VSUBS 0.007176f
C406 B.n366 VSUBS 0.007176f
C407 B.n367 VSUBS 0.007176f
C408 B.n368 VSUBS 0.007176f
C409 B.n369 VSUBS 0.007176f
C410 B.n370 VSUBS 0.007176f
C411 B.n371 VSUBS 0.007176f
C412 B.n372 VSUBS 0.007176f
C413 B.n373 VSUBS 0.007176f
C414 B.n374 VSUBS 0.007176f
C415 B.n375 VSUBS 0.007176f
C416 B.n376 VSUBS 0.007176f
C417 B.n377 VSUBS 0.007176f
C418 B.n378 VSUBS 0.007176f
C419 B.n379 VSUBS 0.007176f
C420 B.n380 VSUBS 0.007176f
C421 B.n381 VSUBS 0.007176f
C422 B.n382 VSUBS 0.007176f
C423 B.n383 VSUBS 0.007176f
C424 B.n384 VSUBS 0.007176f
C425 B.n385 VSUBS 0.007176f
C426 B.n386 VSUBS 0.007176f
C427 B.n387 VSUBS 0.007176f
C428 B.n388 VSUBS 0.007176f
C429 B.n389 VSUBS 0.007176f
C430 B.n390 VSUBS 0.007176f
C431 B.n391 VSUBS 0.007176f
C432 B.n392 VSUBS 0.007176f
C433 B.n393 VSUBS 0.007176f
C434 B.n394 VSUBS 0.007176f
C435 B.n395 VSUBS 0.007176f
C436 B.n396 VSUBS 0.007176f
C437 B.n397 VSUBS 0.007176f
C438 B.n398 VSUBS 0.007176f
C439 B.n399 VSUBS 0.007176f
C440 B.n400 VSUBS 0.007176f
C441 B.n401 VSUBS 0.007176f
C442 B.n402 VSUBS 0.007176f
C443 B.n403 VSUBS 0.007176f
C444 B.n404 VSUBS 0.007176f
C445 B.n405 VSUBS 0.007176f
C446 B.n406 VSUBS 0.007176f
C447 B.n407 VSUBS 0.007176f
C448 B.n408 VSUBS 0.007176f
C449 B.n409 VSUBS 0.007176f
C450 B.n410 VSUBS 0.007176f
C451 B.n411 VSUBS 0.007176f
C452 B.n412 VSUBS 0.007176f
C453 B.n413 VSUBS 0.007176f
C454 B.n414 VSUBS 0.007176f
C455 B.n415 VSUBS 0.007176f
C456 B.n416 VSUBS 0.01619f
C457 B.n417 VSUBS 0.01737f
C458 B.n418 VSUBS 0.01737f
C459 B.n419 VSUBS 0.007176f
C460 B.n420 VSUBS 0.007176f
C461 B.n421 VSUBS 0.007176f
C462 B.n422 VSUBS 0.007176f
C463 B.n423 VSUBS 0.007176f
C464 B.n424 VSUBS 0.007176f
C465 B.n425 VSUBS 0.007176f
C466 B.n426 VSUBS 0.007176f
C467 B.n427 VSUBS 0.007176f
C468 B.n428 VSUBS 0.007176f
C469 B.n429 VSUBS 0.007176f
C470 B.n430 VSUBS 0.007176f
C471 B.n431 VSUBS 0.007176f
C472 B.n432 VSUBS 0.007176f
C473 B.n433 VSUBS 0.007176f
C474 B.n434 VSUBS 0.007176f
C475 B.n435 VSUBS 0.007176f
C476 B.n436 VSUBS 0.007176f
C477 B.n437 VSUBS 0.007176f
C478 B.n438 VSUBS 0.007176f
C479 B.n439 VSUBS 0.007176f
C480 B.n440 VSUBS 0.007176f
C481 B.n441 VSUBS 0.006754f
C482 B.n442 VSUBS 0.007176f
C483 B.n443 VSUBS 0.007176f
C484 B.n444 VSUBS 0.00401f
C485 B.n445 VSUBS 0.007176f
C486 B.n446 VSUBS 0.007176f
C487 B.n447 VSUBS 0.007176f
C488 B.n448 VSUBS 0.007176f
C489 B.n449 VSUBS 0.007176f
C490 B.n450 VSUBS 0.007176f
C491 B.n451 VSUBS 0.007176f
C492 B.n452 VSUBS 0.007176f
C493 B.n453 VSUBS 0.007176f
C494 B.n454 VSUBS 0.007176f
C495 B.n455 VSUBS 0.007176f
C496 B.n456 VSUBS 0.007176f
C497 B.n457 VSUBS 0.00401f
C498 B.n458 VSUBS 0.016627f
C499 B.n459 VSUBS 0.006754f
C500 B.n460 VSUBS 0.007176f
C501 B.n461 VSUBS 0.007176f
C502 B.n462 VSUBS 0.007176f
C503 B.n463 VSUBS 0.007176f
C504 B.n464 VSUBS 0.007176f
C505 B.n465 VSUBS 0.007176f
C506 B.n466 VSUBS 0.007176f
C507 B.n467 VSUBS 0.007176f
C508 B.n468 VSUBS 0.007176f
C509 B.n469 VSUBS 0.007176f
C510 B.n470 VSUBS 0.007176f
C511 B.n471 VSUBS 0.007176f
C512 B.n472 VSUBS 0.007176f
C513 B.n473 VSUBS 0.007176f
C514 B.n474 VSUBS 0.007176f
C515 B.n475 VSUBS 0.007176f
C516 B.n476 VSUBS 0.007176f
C517 B.n477 VSUBS 0.007176f
C518 B.n478 VSUBS 0.007176f
C519 B.n479 VSUBS 0.007176f
C520 B.n480 VSUBS 0.007176f
C521 B.n481 VSUBS 0.007176f
C522 B.n482 VSUBS 0.007176f
C523 B.n483 VSUBS 0.01737f
C524 B.n484 VSUBS 0.01737f
C525 B.n485 VSUBS 0.01619f
C526 B.n486 VSUBS 0.007176f
C527 B.n487 VSUBS 0.007176f
C528 B.n488 VSUBS 0.007176f
C529 B.n489 VSUBS 0.007176f
C530 B.n490 VSUBS 0.007176f
C531 B.n491 VSUBS 0.007176f
C532 B.n492 VSUBS 0.007176f
C533 B.n493 VSUBS 0.007176f
C534 B.n494 VSUBS 0.007176f
C535 B.n495 VSUBS 0.007176f
C536 B.n496 VSUBS 0.007176f
C537 B.n497 VSUBS 0.007176f
C538 B.n498 VSUBS 0.007176f
C539 B.n499 VSUBS 0.007176f
C540 B.n500 VSUBS 0.007176f
C541 B.n501 VSUBS 0.007176f
C542 B.n502 VSUBS 0.007176f
C543 B.n503 VSUBS 0.007176f
C544 B.n504 VSUBS 0.007176f
C545 B.n505 VSUBS 0.007176f
C546 B.n506 VSUBS 0.007176f
C547 B.n507 VSUBS 0.007176f
C548 B.n508 VSUBS 0.007176f
C549 B.n509 VSUBS 0.007176f
C550 B.n510 VSUBS 0.007176f
C551 B.n511 VSUBS 0.007176f
C552 B.n512 VSUBS 0.007176f
C553 B.n513 VSUBS 0.007176f
C554 B.n514 VSUBS 0.007176f
C555 B.n515 VSUBS 0.007176f
C556 B.n516 VSUBS 0.007176f
C557 B.n517 VSUBS 0.007176f
C558 B.n518 VSUBS 0.007176f
C559 B.n519 VSUBS 0.007176f
C560 B.n520 VSUBS 0.007176f
C561 B.n521 VSUBS 0.007176f
C562 B.n522 VSUBS 0.007176f
C563 B.n523 VSUBS 0.007176f
C564 B.n524 VSUBS 0.007176f
C565 B.n525 VSUBS 0.007176f
C566 B.n526 VSUBS 0.007176f
C567 B.n527 VSUBS 0.007176f
C568 B.n528 VSUBS 0.007176f
C569 B.n529 VSUBS 0.007176f
C570 B.n530 VSUBS 0.007176f
C571 B.n531 VSUBS 0.007176f
C572 B.n532 VSUBS 0.007176f
C573 B.n533 VSUBS 0.007176f
C574 B.n534 VSUBS 0.007176f
C575 B.n535 VSUBS 0.007176f
C576 B.n536 VSUBS 0.007176f
C577 B.n537 VSUBS 0.007176f
C578 B.n538 VSUBS 0.007176f
C579 B.n539 VSUBS 0.007176f
C580 B.n540 VSUBS 0.007176f
C581 B.n541 VSUBS 0.007176f
C582 B.n542 VSUBS 0.007176f
C583 B.n543 VSUBS 0.007176f
C584 B.n544 VSUBS 0.007176f
C585 B.n545 VSUBS 0.007176f
C586 B.n546 VSUBS 0.007176f
C587 B.n547 VSUBS 0.007176f
C588 B.n548 VSUBS 0.007176f
C589 B.n549 VSUBS 0.007176f
C590 B.n550 VSUBS 0.007176f
C591 B.n551 VSUBS 0.009365f
C592 B.n552 VSUBS 0.009976f
C593 B.n553 VSUBS 0.019838f
C594 VDD2.t4 VSUBS 0.515946f
C595 VDD2.t3 VSUBS 0.064452f
C596 VDD2.t0 VSUBS 0.064452f
C597 VDD2.n0 VSUBS 0.367646f
C598 VDD2.n1 VSUBS 2.46613f
C599 VDD2.t1 VSUBS 0.508617f
C600 VDD2.n2 VSUBS 2.06477f
C601 VDD2.t5 VSUBS 0.064452f
C602 VDD2.t2 VSUBS 0.064452f
C603 VDD2.n3 VSUBS 0.367627f
C604 VN.t5 VSUBS 1.16751f
C605 VN.n0 VSUBS 0.637584f
C606 VN.n1 VSUBS 0.043787f
C607 VN.n2 VSUBS 0.07494f
C608 VN.n3 VSUBS 0.465159f
C609 VN.t2 VSUBS 1.16751f
C610 VN.t1 VSUBS 1.55027f
C611 VN.n4 VSUBS 0.584626f
C612 VN.n5 VSUBS 0.603104f
C613 VN.n6 VSUBS 0.061156f
C614 VN.n7 VSUBS 0.081199f
C615 VN.n8 VSUBS 0.043787f
C616 VN.n9 VSUBS 0.043787f
C617 VN.n10 VSUBS 0.043787f
C618 VN.n11 VSUBS 0.050904f
C619 VN.n12 VSUBS 0.082657f
C620 VN.n13 VSUBS 0.076388f
C621 VN.n14 VSUBS 0.07066f
C622 VN.n15 VSUBS 0.086075f
C623 VN.t4 VSUBS 1.16751f
C624 VN.n16 VSUBS 0.637584f
C625 VN.n17 VSUBS 0.043787f
C626 VN.n18 VSUBS 0.07494f
C627 VN.n19 VSUBS 0.465159f
C628 VN.t0 VSUBS 1.16751f
C629 VN.t3 VSUBS 1.55027f
C630 VN.n20 VSUBS 0.584626f
C631 VN.n21 VSUBS 0.603104f
C632 VN.n22 VSUBS 0.061156f
C633 VN.n23 VSUBS 0.081199f
C634 VN.n24 VSUBS 0.043787f
C635 VN.n25 VSUBS 0.043787f
C636 VN.n26 VSUBS 0.043787f
C637 VN.n27 VSUBS 0.050904f
C638 VN.n28 VSUBS 0.082657f
C639 VN.n29 VSUBS 0.076388f
C640 VN.n30 VSUBS 0.07066f
C641 VN.n31 VSUBS 2.0211f
C642 VDD1.t1 VSUBS 0.531711f
C643 VDD1.t0 VSUBS 0.531161f
C644 VDD1.t2 VSUBS 0.066353f
C645 VDD1.t3 VSUBS 0.066353f
C646 VDD1.n0 VSUBS 0.378487f
C647 VDD1.n1 VSUBS 2.65094f
C648 VDD1.t4 VSUBS 0.066353f
C649 VDD1.t5 VSUBS 0.066353f
C650 VDD1.n2 VSUBS 0.37556f
C651 VDD1.n3 VSUBS 2.15844f
C652 VTAIL.t5 VSUBS 0.088879f
C653 VTAIL.t3 VSUBS 0.088879f
C654 VTAIL.n0 VSUBS 0.438202f
C655 VTAIL.n1 VSUBS 0.700435f
C656 VTAIL.t10 VSUBS 0.63514f
C657 VTAIL.n2 VSUBS 0.944361f
C658 VTAIL.t6 VSUBS 0.088879f
C659 VTAIL.t9 VSUBS 0.088879f
C660 VTAIL.n3 VSUBS 0.438202f
C661 VTAIL.n4 VSUBS 1.99069f
C662 VTAIL.t1 VSUBS 0.088879f
C663 VTAIL.t4 VSUBS 0.088879f
C664 VTAIL.n5 VSUBS 0.438204f
C665 VTAIL.n6 VSUBS 1.99069f
C666 VTAIL.t0 VSUBS 0.635143f
C667 VTAIL.n7 VSUBS 0.944358f
C668 VTAIL.t11 VSUBS 0.088879f
C669 VTAIL.t8 VSUBS 0.088879f
C670 VTAIL.n8 VSUBS 0.438204f
C671 VTAIL.n9 VSUBS 0.898899f
C672 VTAIL.t7 VSUBS 0.63514f
C673 VTAIL.n10 VSUBS 1.76385f
C674 VTAIL.t2 VSUBS 0.63514f
C675 VTAIL.n11 VSUBS 1.69001f
C676 VP.t2 VSUBS 1.21763f
C677 VP.n0 VSUBS 0.664957f
C678 VP.n1 VSUBS 0.045667f
C679 VP.n2 VSUBS 0.078157f
C680 VP.n3 VSUBS 0.045667f
C681 VP.t3 VSUBS 1.21763f
C682 VP.n4 VSUBS 0.084685f
C683 VP.n5 VSUBS 0.045667f
C684 VP.n6 VSUBS 0.079668f
C685 VP.t0 VSUBS 1.21763f
C686 VP.n7 VSUBS 0.664957f
C687 VP.n8 VSUBS 0.045667f
C688 VP.n9 VSUBS 0.078157f
C689 VP.n10 VSUBS 0.485131f
C690 VP.t1 VSUBS 1.21763f
C691 VP.t4 VSUBS 1.61683f
C692 VP.n11 VSUBS 0.609726f
C693 VP.n12 VSUBS 0.628997f
C694 VP.n13 VSUBS 0.063781f
C695 VP.n14 VSUBS 0.084685f
C696 VP.n15 VSUBS 0.045667f
C697 VP.n16 VSUBS 0.045667f
C698 VP.n17 VSUBS 0.045667f
C699 VP.n18 VSUBS 0.053089f
C700 VP.n19 VSUBS 0.086206f
C701 VP.n20 VSUBS 0.079668f
C702 VP.n21 VSUBS 0.073693f
C703 VP.n22 VSUBS 2.08822f
C704 VP.t5 VSUBS 1.21763f
C705 VP.n23 VSUBS 0.664957f
C706 VP.n24 VSUBS 2.12608f
C707 VP.n25 VSUBS 0.073693f
C708 VP.n26 VSUBS 0.045667f
C709 VP.n27 VSUBS 0.086206f
C710 VP.n28 VSUBS 0.053089f
C711 VP.n29 VSUBS 0.078157f
C712 VP.n30 VSUBS 0.045667f
C713 VP.n31 VSUBS 0.045667f
C714 VP.n32 VSUBS 0.045667f
C715 VP.n33 VSUBS 0.063781f
C716 VP.n34 VSUBS 0.488353f
C717 VP.n35 VSUBS 0.063781f
C718 VP.n36 VSUBS 0.084685f
C719 VP.n37 VSUBS 0.045667f
C720 VP.n38 VSUBS 0.045667f
C721 VP.n39 VSUBS 0.045667f
C722 VP.n40 VSUBS 0.053089f
C723 VP.n41 VSUBS 0.086206f
C724 VP.n42 VSUBS 0.079668f
C725 VP.n43 VSUBS 0.073693f
C726 VP.n44 VSUBS 0.08977f
.ends

