* NGSPICE file created from diff_pair_sample_0953.ext - technology: sky130A

.subckt diff_pair_sample_0953 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t9 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X1 VTAIL.t8 VP.t0 VDD1.t9 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X2 VDD1.t8 VP.t1 VTAIL.t3 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=1.5327 ps=8.64 w=3.93 l=1.25
X3 VDD2.t6 VN.t1 VTAIL.t18 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X4 B.t11 B.t9 B.t10 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0 ps=0 w=3.93 l=1.25
X5 VTAIL.t0 VP.t2 VDD1.t7 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X6 VTAIL.t17 VN.t2 VDD2.t1 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X7 VDD2.t0 VN.t3 VTAIL.t16 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0.64845 ps=4.26 w=3.93 l=1.25
X8 VDD2.t7 VN.t4 VTAIL.t15 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0.64845 ps=4.26 w=3.93 l=1.25
X9 B.t8 B.t6 B.t7 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0 ps=0 w=3.93 l=1.25
X10 VDD1.t6 VP.t3 VTAIL.t5 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X11 VDD2.t4 VN.t5 VTAIL.t14 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=1.5327 ps=8.64 w=3.93 l=1.25
X12 VTAIL.t13 VN.t6 VDD2.t3 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X13 VDD1.t5 VP.t4 VTAIL.t7 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0.64845 ps=4.26 w=3.93 l=1.25
X14 B.t5 B.t3 B.t4 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0 ps=0 w=3.93 l=1.25
X15 VDD1.t4 VP.t5 VTAIL.t4 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=1.5327 ps=8.64 w=3.93 l=1.25
X16 VTAIL.t12 VN.t7 VDD2.t2 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X17 VTAIL.t9 VP.t6 VDD1.t3 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X18 VDD1.t2 VP.t7 VTAIL.t6 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X19 B.t2 B.t0 B.t1 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0 ps=0 w=3.93 l=1.25
X20 VDD2.t8 VN.t8 VTAIL.t11 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X21 VTAIL.t1 VP.t8 VDD1.t1 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=0.64845 ps=4.26 w=3.93 l=1.25
X22 VDD1.t0 VP.t9 VTAIL.t2 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=1.5327 pd=8.64 as=0.64845 ps=4.26 w=3.93 l=1.25
X23 VDD2.t5 VN.t9 VTAIL.t10 w_n2866_n1754# sky130_fd_pr__pfet_01v8 ad=0.64845 pd=4.26 as=1.5327 ps=8.64 w=3.93 l=1.25
R0 VN.n41 VN.n22 161.3
R1 VN.n40 VN.n39 161.3
R2 VN.n38 VN.n37 161.3
R3 VN.n36 VN.n24 161.3
R4 VN.n35 VN.n34 161.3
R5 VN.n33 VN.n32 161.3
R6 VN.n31 VN.n26 161.3
R7 VN.n30 VN.n29 161.3
R8 VN.n19 VN.n0 161.3
R9 VN.n18 VN.n17 161.3
R10 VN.n16 VN.n15 161.3
R11 VN.n14 VN.n2 161.3
R12 VN.n13 VN.n12 161.3
R13 VN.n11 VN.n10 161.3
R14 VN.n9 VN.n4 161.3
R15 VN.n8 VN.n7 161.3
R16 VN.n6 VN.t4 128.577
R17 VN.n28 VN.t5 128.577
R18 VN.n20 VN.t9 107.391
R19 VN.n42 VN.t3 107.391
R20 VN.n43 VN.n42 80.6037
R21 VN.n21 VN.n20 80.6037
R22 VN.n5 VN.t6 75.7709
R23 VN.n3 VN.t8 75.7709
R24 VN.n1 VN.t7 75.7709
R25 VN.n27 VN.t2 75.7709
R26 VN.n25 VN.t1 75.7709
R27 VN.n23 VN.t0 75.7709
R28 VN.n9 VN.n8 44.3785
R29 VN.n15 VN.n14 44.3785
R30 VN.n31 VN.n30 44.3785
R31 VN.n37 VN.n36 44.3785
R32 VN.n20 VN.n19 41.6278
R33 VN.n42 VN.n41 41.6278
R34 VN.n6 VN.n5 40.893
R35 VN.n28 VN.n27 40.893
R36 VN VN.n43 40.1581
R37 VN.n10 VN.n9 36.6083
R38 VN.n14 VN.n13 36.6083
R39 VN.n32 VN.n31 36.6083
R40 VN.n36 VN.n35 36.6083
R41 VN.n19 VN.n18 28.8382
R42 VN.n41 VN.n40 28.8382
R43 VN.n29 VN.n28 28.8325
R44 VN.n7 VN.n6 28.8325
R45 VN.n8 VN.n5 16.1487
R46 VN.n15 VN.n1 16.1487
R47 VN.n30 VN.n27 16.1487
R48 VN.n37 VN.n23 16.1487
R49 VN.n10 VN.n3 12.234
R50 VN.n13 VN.n3 12.234
R51 VN.n35 VN.n25 12.234
R52 VN.n32 VN.n25 12.234
R53 VN.n18 VN.n1 8.31928
R54 VN.n40 VN.n23 8.31928
R55 VN.n43 VN.n22 0.285035
R56 VN.n21 VN.n0 0.285035
R57 VN.n39 VN.n22 0.189894
R58 VN.n39 VN.n38 0.189894
R59 VN.n38 VN.n24 0.189894
R60 VN.n34 VN.n24 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n26 0.189894
R63 VN.n29 VN.n26 0.189894
R64 VN.n7 VN.n4 0.189894
R65 VN.n11 VN.n4 0.189894
R66 VN.n12 VN.n11 0.189894
R67 VN.n12 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n17 VN.n0 0.189894
R71 VN VN.n21 0.146778
R72 VDD2.n37 VDD2.n23 756.745
R73 VDD2.n14 VDD2.n0 756.745
R74 VDD2.n38 VDD2.n37 585
R75 VDD2.n36 VDD2.n35 585
R76 VDD2.n27 VDD2.n26 585
R77 VDD2.n30 VDD2.n29 585
R78 VDD2.n7 VDD2.n6 585
R79 VDD2.n4 VDD2.n3 585
R80 VDD2.n13 VDD2.n12 585
R81 VDD2.n15 VDD2.n14 585
R82 VDD2.t0 VDD2.n28 330.707
R83 VDD2.t7 VDD2.n5 330.707
R84 VDD2.n37 VDD2.n36 171.744
R85 VDD2.n36 VDD2.n26 171.744
R86 VDD2.n29 VDD2.n26 171.744
R87 VDD2.n6 VDD2.n3 171.744
R88 VDD2.n13 VDD2.n3 171.744
R89 VDD2.n14 VDD2.n13 171.744
R90 VDD2.n22 VDD2.n21 116.279
R91 VDD2 VDD2.n45 116.276
R92 VDD2.n44 VDD2.n43 115.314
R93 VDD2.n20 VDD2.n19 115.314
R94 VDD2.n29 VDD2.t0 85.8723
R95 VDD2.n6 VDD2.t7 85.8723
R96 VDD2.n20 VDD2.n18 51.9717
R97 VDD2.n42 VDD2.n41 50.6096
R98 VDD2.n42 VDD2.n22 33.5731
R99 VDD2.n30 VDD2.n28 16.3201
R100 VDD2.n7 VDD2.n5 16.3201
R101 VDD2.n31 VDD2.n27 12.8005
R102 VDD2.n8 VDD2.n4 12.8005
R103 VDD2.n35 VDD2.n34 12.0247
R104 VDD2.n12 VDD2.n11 12.0247
R105 VDD2.n38 VDD2.n25 11.249
R106 VDD2.n15 VDD2.n2 11.249
R107 VDD2.n39 VDD2.n23 10.4732
R108 VDD2.n16 VDD2.n0 10.4732
R109 VDD2.n41 VDD2.n40 9.45567
R110 VDD2.n18 VDD2.n17 9.45567
R111 VDD2.n40 VDD2.n39 9.3005
R112 VDD2.n25 VDD2.n24 9.3005
R113 VDD2.n34 VDD2.n33 9.3005
R114 VDD2.n32 VDD2.n31 9.3005
R115 VDD2.n17 VDD2.n16 9.3005
R116 VDD2.n2 VDD2.n1 9.3005
R117 VDD2.n11 VDD2.n10 9.3005
R118 VDD2.n9 VDD2.n8 9.3005
R119 VDD2.n45 VDD2.t1 8.27149
R120 VDD2.n45 VDD2.t4 8.27149
R121 VDD2.n43 VDD2.t9 8.27149
R122 VDD2.n43 VDD2.t6 8.27149
R123 VDD2.n21 VDD2.t2 8.27149
R124 VDD2.n21 VDD2.t5 8.27149
R125 VDD2.n19 VDD2.t3 8.27149
R126 VDD2.n19 VDD2.t8 8.27149
R127 VDD2.n32 VDD2.n28 3.78097
R128 VDD2.n9 VDD2.n5 3.78097
R129 VDD2.n41 VDD2.n23 3.49141
R130 VDD2.n18 VDD2.n0 3.49141
R131 VDD2.n39 VDD2.n38 2.71565
R132 VDD2.n16 VDD2.n15 2.71565
R133 VDD2.n35 VDD2.n25 1.93989
R134 VDD2.n12 VDD2.n2 1.93989
R135 VDD2.n44 VDD2.n42 1.36257
R136 VDD2.n34 VDD2.n27 1.16414
R137 VDD2.n11 VDD2.n4 1.16414
R138 VDD2 VDD2.n44 0.399207
R139 VDD2.n31 VDD2.n30 0.388379
R140 VDD2.n8 VDD2.n7 0.388379
R141 VDD2.n22 VDD2.n20 0.285671
R142 VDD2.n40 VDD2.n24 0.155672
R143 VDD2.n33 VDD2.n24 0.155672
R144 VDD2.n33 VDD2.n32 0.155672
R145 VDD2.n10 VDD2.n9 0.155672
R146 VDD2.n10 VDD2.n1 0.155672
R147 VDD2.n17 VDD2.n1 0.155672
R148 VTAIL.n88 VTAIL.n74 756.745
R149 VTAIL.n16 VTAIL.n2 756.745
R150 VTAIL.n68 VTAIL.n54 756.745
R151 VTAIL.n44 VTAIL.n30 756.745
R152 VTAIL.n81 VTAIL.n80 585
R153 VTAIL.n78 VTAIL.n77 585
R154 VTAIL.n87 VTAIL.n86 585
R155 VTAIL.n89 VTAIL.n88 585
R156 VTAIL.n9 VTAIL.n8 585
R157 VTAIL.n6 VTAIL.n5 585
R158 VTAIL.n15 VTAIL.n14 585
R159 VTAIL.n17 VTAIL.n16 585
R160 VTAIL.n69 VTAIL.n68 585
R161 VTAIL.n67 VTAIL.n66 585
R162 VTAIL.n58 VTAIL.n57 585
R163 VTAIL.n61 VTAIL.n60 585
R164 VTAIL.n45 VTAIL.n44 585
R165 VTAIL.n43 VTAIL.n42 585
R166 VTAIL.n34 VTAIL.n33 585
R167 VTAIL.n37 VTAIL.n36 585
R168 VTAIL.t10 VTAIL.n79 330.707
R169 VTAIL.t4 VTAIL.n7 330.707
R170 VTAIL.t3 VTAIL.n59 330.707
R171 VTAIL.t14 VTAIL.n35 330.707
R172 VTAIL.n80 VTAIL.n77 171.744
R173 VTAIL.n87 VTAIL.n77 171.744
R174 VTAIL.n88 VTAIL.n87 171.744
R175 VTAIL.n8 VTAIL.n5 171.744
R176 VTAIL.n15 VTAIL.n5 171.744
R177 VTAIL.n16 VTAIL.n15 171.744
R178 VTAIL.n68 VTAIL.n67 171.744
R179 VTAIL.n67 VTAIL.n57 171.744
R180 VTAIL.n60 VTAIL.n57 171.744
R181 VTAIL.n44 VTAIL.n43 171.744
R182 VTAIL.n43 VTAIL.n33 171.744
R183 VTAIL.n36 VTAIL.n33 171.744
R184 VTAIL.n53 VTAIL.n52 98.635
R185 VTAIL.n51 VTAIL.n50 98.635
R186 VTAIL.n29 VTAIL.n28 98.635
R187 VTAIL.n27 VTAIL.n26 98.635
R188 VTAIL.n95 VTAIL.n94 98.6348
R189 VTAIL.n1 VTAIL.n0 98.6348
R190 VTAIL.n23 VTAIL.n22 98.6348
R191 VTAIL.n25 VTAIL.n24 98.6348
R192 VTAIL.n80 VTAIL.t10 85.8723
R193 VTAIL.n8 VTAIL.t4 85.8723
R194 VTAIL.n60 VTAIL.t3 85.8723
R195 VTAIL.n36 VTAIL.t14 85.8723
R196 VTAIL.n93 VTAIL.n92 33.9308
R197 VTAIL.n21 VTAIL.n20 33.9308
R198 VTAIL.n73 VTAIL.n72 33.9308
R199 VTAIL.n49 VTAIL.n48 33.9308
R200 VTAIL.n27 VTAIL.n25 18.4789
R201 VTAIL.n93 VTAIL.n73 17.1169
R202 VTAIL.n81 VTAIL.n79 16.3201
R203 VTAIL.n9 VTAIL.n7 16.3201
R204 VTAIL.n61 VTAIL.n59 16.3201
R205 VTAIL.n37 VTAIL.n35 16.3201
R206 VTAIL.n82 VTAIL.n78 12.8005
R207 VTAIL.n10 VTAIL.n6 12.8005
R208 VTAIL.n62 VTAIL.n58 12.8005
R209 VTAIL.n38 VTAIL.n34 12.8005
R210 VTAIL.n86 VTAIL.n85 12.0247
R211 VTAIL.n14 VTAIL.n13 12.0247
R212 VTAIL.n66 VTAIL.n65 12.0247
R213 VTAIL.n42 VTAIL.n41 12.0247
R214 VTAIL.n89 VTAIL.n76 11.249
R215 VTAIL.n17 VTAIL.n4 11.249
R216 VTAIL.n69 VTAIL.n56 11.249
R217 VTAIL.n45 VTAIL.n32 11.249
R218 VTAIL.n90 VTAIL.n74 10.4732
R219 VTAIL.n18 VTAIL.n2 10.4732
R220 VTAIL.n70 VTAIL.n54 10.4732
R221 VTAIL.n46 VTAIL.n30 10.4732
R222 VTAIL.n92 VTAIL.n91 9.45567
R223 VTAIL.n20 VTAIL.n19 9.45567
R224 VTAIL.n72 VTAIL.n71 9.45567
R225 VTAIL.n48 VTAIL.n47 9.45567
R226 VTAIL.n91 VTAIL.n90 9.3005
R227 VTAIL.n76 VTAIL.n75 9.3005
R228 VTAIL.n85 VTAIL.n84 9.3005
R229 VTAIL.n83 VTAIL.n82 9.3005
R230 VTAIL.n19 VTAIL.n18 9.3005
R231 VTAIL.n4 VTAIL.n3 9.3005
R232 VTAIL.n13 VTAIL.n12 9.3005
R233 VTAIL.n11 VTAIL.n10 9.3005
R234 VTAIL.n71 VTAIL.n70 9.3005
R235 VTAIL.n56 VTAIL.n55 9.3005
R236 VTAIL.n65 VTAIL.n64 9.3005
R237 VTAIL.n63 VTAIL.n62 9.3005
R238 VTAIL.n47 VTAIL.n46 9.3005
R239 VTAIL.n32 VTAIL.n31 9.3005
R240 VTAIL.n41 VTAIL.n40 9.3005
R241 VTAIL.n39 VTAIL.n38 9.3005
R242 VTAIL.n94 VTAIL.t11 8.27149
R243 VTAIL.n94 VTAIL.t12 8.27149
R244 VTAIL.n0 VTAIL.t15 8.27149
R245 VTAIL.n0 VTAIL.t13 8.27149
R246 VTAIL.n22 VTAIL.t6 8.27149
R247 VTAIL.n22 VTAIL.t8 8.27149
R248 VTAIL.n24 VTAIL.t2 8.27149
R249 VTAIL.n24 VTAIL.t1 8.27149
R250 VTAIL.n52 VTAIL.t5 8.27149
R251 VTAIL.n52 VTAIL.t0 8.27149
R252 VTAIL.n50 VTAIL.t7 8.27149
R253 VTAIL.n50 VTAIL.t9 8.27149
R254 VTAIL.n28 VTAIL.t18 8.27149
R255 VTAIL.n28 VTAIL.t17 8.27149
R256 VTAIL.n26 VTAIL.t16 8.27149
R257 VTAIL.n26 VTAIL.t19 8.27149
R258 VTAIL.n83 VTAIL.n79 3.78097
R259 VTAIL.n11 VTAIL.n7 3.78097
R260 VTAIL.n63 VTAIL.n59 3.78097
R261 VTAIL.n39 VTAIL.n35 3.78097
R262 VTAIL.n92 VTAIL.n74 3.49141
R263 VTAIL.n20 VTAIL.n2 3.49141
R264 VTAIL.n72 VTAIL.n54 3.49141
R265 VTAIL.n48 VTAIL.n30 3.49141
R266 VTAIL.n90 VTAIL.n89 2.71565
R267 VTAIL.n18 VTAIL.n17 2.71565
R268 VTAIL.n70 VTAIL.n69 2.71565
R269 VTAIL.n46 VTAIL.n45 2.71565
R270 VTAIL.n86 VTAIL.n76 1.93989
R271 VTAIL.n14 VTAIL.n4 1.93989
R272 VTAIL.n66 VTAIL.n56 1.93989
R273 VTAIL.n42 VTAIL.n32 1.93989
R274 VTAIL.n29 VTAIL.n27 1.36257
R275 VTAIL.n49 VTAIL.n29 1.36257
R276 VTAIL.n53 VTAIL.n51 1.36257
R277 VTAIL.n73 VTAIL.n53 1.36257
R278 VTAIL.n25 VTAIL.n23 1.36257
R279 VTAIL.n23 VTAIL.n21 1.36257
R280 VTAIL.n95 VTAIL.n93 1.36257
R281 VTAIL.n85 VTAIL.n78 1.16414
R282 VTAIL.n13 VTAIL.n6 1.16414
R283 VTAIL.n65 VTAIL.n58 1.16414
R284 VTAIL.n41 VTAIL.n34 1.16414
R285 VTAIL.n51 VTAIL.n49 1.15136
R286 VTAIL.n21 VTAIL.n1 1.15136
R287 VTAIL VTAIL.n1 1.08024
R288 VTAIL.n82 VTAIL.n81 0.388379
R289 VTAIL.n10 VTAIL.n9 0.388379
R290 VTAIL.n62 VTAIL.n61 0.388379
R291 VTAIL.n38 VTAIL.n37 0.388379
R292 VTAIL VTAIL.n95 0.282828
R293 VTAIL.n84 VTAIL.n83 0.155672
R294 VTAIL.n84 VTAIL.n75 0.155672
R295 VTAIL.n91 VTAIL.n75 0.155672
R296 VTAIL.n12 VTAIL.n11 0.155672
R297 VTAIL.n12 VTAIL.n3 0.155672
R298 VTAIL.n19 VTAIL.n3 0.155672
R299 VTAIL.n71 VTAIL.n55 0.155672
R300 VTAIL.n64 VTAIL.n55 0.155672
R301 VTAIL.n64 VTAIL.n63 0.155672
R302 VTAIL.n47 VTAIL.n31 0.155672
R303 VTAIL.n40 VTAIL.n31 0.155672
R304 VTAIL.n40 VTAIL.n39 0.155672
R305 VP.n15 VP.n14 161.3
R306 VP.n16 VP.n11 161.3
R307 VP.n18 VP.n17 161.3
R308 VP.n20 VP.n19 161.3
R309 VP.n21 VP.n9 161.3
R310 VP.n23 VP.n22 161.3
R311 VP.n25 VP.n24 161.3
R312 VP.n26 VP.n7 161.3
R313 VP.n46 VP.n0 161.3
R314 VP.n45 VP.n44 161.3
R315 VP.n43 VP.n42 161.3
R316 VP.n41 VP.n2 161.3
R317 VP.n40 VP.n39 161.3
R318 VP.n38 VP.n37 161.3
R319 VP.n36 VP.n4 161.3
R320 VP.n35 VP.n34 161.3
R321 VP.n33 VP.n32 161.3
R322 VP.n31 VP.n6 161.3
R323 VP.n13 VP.t4 128.577
R324 VP.n30 VP.t9 107.391
R325 VP.n47 VP.t5 107.391
R326 VP.n27 VP.t1 107.391
R327 VP.n28 VP.n27 80.6037
R328 VP.n48 VP.n47 80.6037
R329 VP.n30 VP.n29 80.6037
R330 VP.n5 VP.t8 75.7709
R331 VP.n3 VP.t7 75.7709
R332 VP.n1 VP.t0 75.7709
R333 VP.n8 VP.t2 75.7709
R334 VP.n10 VP.t3 75.7709
R335 VP.n12 VP.t6 75.7709
R336 VP.n36 VP.n35 44.3785
R337 VP.n42 VP.n41 44.3785
R338 VP.n22 VP.n21 44.3785
R339 VP.n16 VP.n15 44.3785
R340 VP.n31 VP.n30 41.6278
R341 VP.n47 VP.n46 41.6278
R342 VP.n27 VP.n26 41.6278
R343 VP.n13 VP.n12 40.893
R344 VP.n29 VP.n28 39.8726
R345 VP.n37 VP.n36 36.6083
R346 VP.n41 VP.n40 36.6083
R347 VP.n21 VP.n20 36.6083
R348 VP.n17 VP.n16 36.6083
R349 VP.n32 VP.n31 28.8382
R350 VP.n46 VP.n45 28.8382
R351 VP.n26 VP.n25 28.8382
R352 VP.n14 VP.n13 28.8325
R353 VP.n35 VP.n5 16.1487
R354 VP.n42 VP.n1 16.1487
R355 VP.n22 VP.n8 16.1487
R356 VP.n15 VP.n12 16.1487
R357 VP.n37 VP.n3 12.234
R358 VP.n40 VP.n3 12.234
R359 VP.n17 VP.n10 12.234
R360 VP.n20 VP.n10 12.234
R361 VP.n32 VP.n5 8.31928
R362 VP.n45 VP.n1 8.31928
R363 VP.n25 VP.n8 8.31928
R364 VP.n28 VP.n7 0.285035
R365 VP.n29 VP.n6 0.285035
R366 VP.n48 VP.n0 0.285035
R367 VP.n14 VP.n11 0.189894
R368 VP.n18 VP.n11 0.189894
R369 VP.n19 VP.n18 0.189894
R370 VP.n19 VP.n9 0.189894
R371 VP.n23 VP.n9 0.189894
R372 VP.n24 VP.n23 0.189894
R373 VP.n24 VP.n7 0.189894
R374 VP.n33 VP.n6 0.189894
R375 VP.n34 VP.n33 0.189894
R376 VP.n34 VP.n4 0.189894
R377 VP.n38 VP.n4 0.189894
R378 VP.n39 VP.n38 0.189894
R379 VP.n39 VP.n2 0.189894
R380 VP.n43 VP.n2 0.189894
R381 VP.n44 VP.n43 0.189894
R382 VP.n44 VP.n0 0.189894
R383 VP VP.n48 0.146778
R384 VDD1.n14 VDD1.n0 756.745
R385 VDD1.n35 VDD1.n21 756.745
R386 VDD1.n15 VDD1.n14 585
R387 VDD1.n13 VDD1.n12 585
R388 VDD1.n4 VDD1.n3 585
R389 VDD1.n7 VDD1.n6 585
R390 VDD1.n28 VDD1.n27 585
R391 VDD1.n25 VDD1.n24 585
R392 VDD1.n34 VDD1.n33 585
R393 VDD1.n36 VDD1.n35 585
R394 VDD1.t5 VDD1.n5 330.707
R395 VDD1.t0 VDD1.n26 330.707
R396 VDD1.n14 VDD1.n13 171.744
R397 VDD1.n13 VDD1.n3 171.744
R398 VDD1.n6 VDD1.n3 171.744
R399 VDD1.n27 VDD1.n24 171.744
R400 VDD1.n34 VDD1.n24 171.744
R401 VDD1.n35 VDD1.n34 171.744
R402 VDD1.n43 VDD1.n42 116.279
R403 VDD1.n20 VDD1.n19 115.314
R404 VDD1.n45 VDD1.n44 115.314
R405 VDD1.n41 VDD1.n40 115.314
R406 VDD1.n6 VDD1.t5 85.8723
R407 VDD1.n27 VDD1.t0 85.8723
R408 VDD1.n20 VDD1.n18 51.9717
R409 VDD1.n41 VDD1.n39 51.9717
R410 VDD1.n45 VDD1.n43 34.8371
R411 VDD1.n7 VDD1.n5 16.3201
R412 VDD1.n28 VDD1.n26 16.3201
R413 VDD1.n8 VDD1.n4 12.8005
R414 VDD1.n29 VDD1.n25 12.8005
R415 VDD1.n12 VDD1.n11 12.0247
R416 VDD1.n33 VDD1.n32 12.0247
R417 VDD1.n15 VDD1.n2 11.249
R418 VDD1.n36 VDD1.n23 11.249
R419 VDD1.n16 VDD1.n0 10.4732
R420 VDD1.n37 VDD1.n21 10.4732
R421 VDD1.n18 VDD1.n17 9.45567
R422 VDD1.n39 VDD1.n38 9.45567
R423 VDD1.n17 VDD1.n16 9.3005
R424 VDD1.n2 VDD1.n1 9.3005
R425 VDD1.n11 VDD1.n10 9.3005
R426 VDD1.n9 VDD1.n8 9.3005
R427 VDD1.n38 VDD1.n37 9.3005
R428 VDD1.n23 VDD1.n22 9.3005
R429 VDD1.n32 VDD1.n31 9.3005
R430 VDD1.n30 VDD1.n29 9.3005
R431 VDD1.n44 VDD1.t7 8.27149
R432 VDD1.n44 VDD1.t8 8.27149
R433 VDD1.n19 VDD1.t3 8.27149
R434 VDD1.n19 VDD1.t6 8.27149
R435 VDD1.n42 VDD1.t9 8.27149
R436 VDD1.n42 VDD1.t4 8.27149
R437 VDD1.n40 VDD1.t1 8.27149
R438 VDD1.n40 VDD1.t2 8.27149
R439 VDD1.n9 VDD1.n5 3.78097
R440 VDD1.n30 VDD1.n26 3.78097
R441 VDD1.n18 VDD1.n0 3.49141
R442 VDD1.n39 VDD1.n21 3.49141
R443 VDD1.n16 VDD1.n15 2.71565
R444 VDD1.n37 VDD1.n36 2.71565
R445 VDD1.n12 VDD1.n2 1.93989
R446 VDD1.n33 VDD1.n23 1.93989
R447 VDD1.n11 VDD1.n4 1.16414
R448 VDD1.n32 VDD1.n25 1.16414
R449 VDD1 VDD1.n45 0.963862
R450 VDD1 VDD1.n20 0.399207
R451 VDD1.n8 VDD1.n7 0.388379
R452 VDD1.n29 VDD1.n28 0.388379
R453 VDD1.n43 VDD1.n41 0.285671
R454 VDD1.n17 VDD1.n1 0.155672
R455 VDD1.n10 VDD1.n1 0.155672
R456 VDD1.n10 VDD1.n9 0.155672
R457 VDD1.n31 VDD1.n30 0.155672
R458 VDD1.n31 VDD1.n22 0.155672
R459 VDD1.n38 VDD1.n22 0.155672
R460 B.n359 B.n46 585
R461 B.n361 B.n360 585
R462 B.n362 B.n45 585
R463 B.n364 B.n363 585
R464 B.n365 B.n44 585
R465 B.n367 B.n366 585
R466 B.n368 B.n43 585
R467 B.n370 B.n369 585
R468 B.n371 B.n42 585
R469 B.n373 B.n372 585
R470 B.n374 B.n41 585
R471 B.n376 B.n375 585
R472 B.n377 B.n40 585
R473 B.n379 B.n378 585
R474 B.n380 B.n39 585
R475 B.n382 B.n381 585
R476 B.n383 B.n38 585
R477 B.n385 B.n384 585
R478 B.n387 B.n35 585
R479 B.n389 B.n388 585
R480 B.n390 B.n34 585
R481 B.n392 B.n391 585
R482 B.n393 B.n33 585
R483 B.n395 B.n394 585
R484 B.n396 B.n32 585
R485 B.n398 B.n397 585
R486 B.n399 B.n29 585
R487 B.n402 B.n401 585
R488 B.n403 B.n28 585
R489 B.n405 B.n404 585
R490 B.n406 B.n27 585
R491 B.n408 B.n407 585
R492 B.n409 B.n26 585
R493 B.n411 B.n410 585
R494 B.n412 B.n25 585
R495 B.n414 B.n413 585
R496 B.n415 B.n24 585
R497 B.n417 B.n416 585
R498 B.n418 B.n23 585
R499 B.n420 B.n419 585
R500 B.n421 B.n22 585
R501 B.n423 B.n422 585
R502 B.n424 B.n21 585
R503 B.n426 B.n425 585
R504 B.n427 B.n20 585
R505 B.n358 B.n357 585
R506 B.n356 B.n47 585
R507 B.n355 B.n354 585
R508 B.n353 B.n48 585
R509 B.n352 B.n351 585
R510 B.n350 B.n49 585
R511 B.n349 B.n348 585
R512 B.n347 B.n50 585
R513 B.n346 B.n345 585
R514 B.n344 B.n51 585
R515 B.n343 B.n342 585
R516 B.n341 B.n52 585
R517 B.n340 B.n339 585
R518 B.n338 B.n53 585
R519 B.n337 B.n336 585
R520 B.n335 B.n54 585
R521 B.n334 B.n333 585
R522 B.n332 B.n55 585
R523 B.n331 B.n330 585
R524 B.n329 B.n56 585
R525 B.n328 B.n327 585
R526 B.n326 B.n57 585
R527 B.n325 B.n324 585
R528 B.n323 B.n58 585
R529 B.n322 B.n321 585
R530 B.n320 B.n59 585
R531 B.n319 B.n318 585
R532 B.n317 B.n60 585
R533 B.n316 B.n315 585
R534 B.n314 B.n61 585
R535 B.n313 B.n312 585
R536 B.n311 B.n62 585
R537 B.n310 B.n309 585
R538 B.n308 B.n63 585
R539 B.n307 B.n306 585
R540 B.n305 B.n64 585
R541 B.n304 B.n303 585
R542 B.n302 B.n65 585
R543 B.n301 B.n300 585
R544 B.n299 B.n66 585
R545 B.n298 B.n297 585
R546 B.n296 B.n67 585
R547 B.n295 B.n294 585
R548 B.n293 B.n68 585
R549 B.n292 B.n291 585
R550 B.n290 B.n69 585
R551 B.n289 B.n288 585
R552 B.n287 B.n70 585
R553 B.n286 B.n285 585
R554 B.n284 B.n71 585
R555 B.n283 B.n282 585
R556 B.n281 B.n72 585
R557 B.n280 B.n279 585
R558 B.n278 B.n73 585
R559 B.n277 B.n276 585
R560 B.n275 B.n74 585
R561 B.n274 B.n273 585
R562 B.n272 B.n75 585
R563 B.n271 B.n270 585
R564 B.n269 B.n76 585
R565 B.n268 B.n267 585
R566 B.n266 B.n77 585
R567 B.n265 B.n264 585
R568 B.n263 B.n78 585
R569 B.n262 B.n261 585
R570 B.n260 B.n79 585
R571 B.n259 B.n258 585
R572 B.n257 B.n80 585
R573 B.n256 B.n255 585
R574 B.n254 B.n81 585
R575 B.n253 B.n252 585
R576 B.n251 B.n82 585
R577 B.n250 B.n249 585
R578 B.n181 B.n180 585
R579 B.n182 B.n109 585
R580 B.n184 B.n183 585
R581 B.n185 B.n108 585
R582 B.n187 B.n186 585
R583 B.n188 B.n107 585
R584 B.n190 B.n189 585
R585 B.n191 B.n106 585
R586 B.n193 B.n192 585
R587 B.n194 B.n105 585
R588 B.n196 B.n195 585
R589 B.n197 B.n104 585
R590 B.n199 B.n198 585
R591 B.n200 B.n103 585
R592 B.n202 B.n201 585
R593 B.n203 B.n102 585
R594 B.n205 B.n204 585
R595 B.n206 B.n99 585
R596 B.n209 B.n208 585
R597 B.n210 B.n98 585
R598 B.n212 B.n211 585
R599 B.n213 B.n97 585
R600 B.n215 B.n214 585
R601 B.n216 B.n96 585
R602 B.n218 B.n217 585
R603 B.n219 B.n95 585
R604 B.n221 B.n220 585
R605 B.n223 B.n222 585
R606 B.n224 B.n91 585
R607 B.n226 B.n225 585
R608 B.n227 B.n90 585
R609 B.n229 B.n228 585
R610 B.n230 B.n89 585
R611 B.n232 B.n231 585
R612 B.n233 B.n88 585
R613 B.n235 B.n234 585
R614 B.n236 B.n87 585
R615 B.n238 B.n237 585
R616 B.n239 B.n86 585
R617 B.n241 B.n240 585
R618 B.n242 B.n85 585
R619 B.n244 B.n243 585
R620 B.n245 B.n84 585
R621 B.n247 B.n246 585
R622 B.n248 B.n83 585
R623 B.n179 B.n110 585
R624 B.n178 B.n177 585
R625 B.n176 B.n111 585
R626 B.n175 B.n174 585
R627 B.n173 B.n112 585
R628 B.n172 B.n171 585
R629 B.n170 B.n113 585
R630 B.n169 B.n168 585
R631 B.n167 B.n114 585
R632 B.n166 B.n165 585
R633 B.n164 B.n115 585
R634 B.n163 B.n162 585
R635 B.n161 B.n116 585
R636 B.n160 B.n159 585
R637 B.n158 B.n117 585
R638 B.n157 B.n156 585
R639 B.n155 B.n118 585
R640 B.n154 B.n153 585
R641 B.n152 B.n119 585
R642 B.n151 B.n150 585
R643 B.n149 B.n120 585
R644 B.n148 B.n147 585
R645 B.n146 B.n121 585
R646 B.n145 B.n144 585
R647 B.n143 B.n122 585
R648 B.n142 B.n141 585
R649 B.n140 B.n123 585
R650 B.n139 B.n138 585
R651 B.n137 B.n124 585
R652 B.n136 B.n135 585
R653 B.n134 B.n125 585
R654 B.n133 B.n132 585
R655 B.n131 B.n126 585
R656 B.n130 B.n129 585
R657 B.n128 B.n127 585
R658 B.n2 B.n0 585
R659 B.n481 B.n1 585
R660 B.n480 B.n479 585
R661 B.n478 B.n3 585
R662 B.n477 B.n476 585
R663 B.n475 B.n4 585
R664 B.n474 B.n473 585
R665 B.n472 B.n5 585
R666 B.n471 B.n470 585
R667 B.n469 B.n6 585
R668 B.n468 B.n467 585
R669 B.n466 B.n7 585
R670 B.n465 B.n464 585
R671 B.n463 B.n8 585
R672 B.n462 B.n461 585
R673 B.n460 B.n9 585
R674 B.n459 B.n458 585
R675 B.n457 B.n10 585
R676 B.n456 B.n455 585
R677 B.n454 B.n11 585
R678 B.n453 B.n452 585
R679 B.n451 B.n12 585
R680 B.n450 B.n449 585
R681 B.n448 B.n13 585
R682 B.n447 B.n446 585
R683 B.n445 B.n14 585
R684 B.n444 B.n443 585
R685 B.n442 B.n15 585
R686 B.n441 B.n440 585
R687 B.n439 B.n16 585
R688 B.n438 B.n437 585
R689 B.n436 B.n17 585
R690 B.n435 B.n434 585
R691 B.n433 B.n18 585
R692 B.n432 B.n431 585
R693 B.n430 B.n19 585
R694 B.n429 B.n428 585
R695 B.n483 B.n482 585
R696 B.n180 B.n179 526.135
R697 B.n428 B.n427 526.135
R698 B.n250 B.n83 526.135
R699 B.n359 B.n358 526.135
R700 B.n92 B.t9 280.142
R701 B.n100 B.t0 280.142
R702 B.n30 B.t6 280.142
R703 B.n36 B.t3 280.142
R704 B.n92 B.t11 264.914
R705 B.n36 B.t4 264.914
R706 B.n100 B.t2 264.914
R707 B.n30 B.t7 264.914
R708 B.n93 B.t10 234.272
R709 B.n37 B.t5 234.272
R710 B.n101 B.t1 234.272
R711 B.n31 B.t8 234.272
R712 B.n179 B.n178 163.367
R713 B.n178 B.n111 163.367
R714 B.n174 B.n111 163.367
R715 B.n174 B.n173 163.367
R716 B.n173 B.n172 163.367
R717 B.n172 B.n113 163.367
R718 B.n168 B.n113 163.367
R719 B.n168 B.n167 163.367
R720 B.n167 B.n166 163.367
R721 B.n166 B.n115 163.367
R722 B.n162 B.n115 163.367
R723 B.n162 B.n161 163.367
R724 B.n161 B.n160 163.367
R725 B.n160 B.n117 163.367
R726 B.n156 B.n117 163.367
R727 B.n156 B.n155 163.367
R728 B.n155 B.n154 163.367
R729 B.n154 B.n119 163.367
R730 B.n150 B.n119 163.367
R731 B.n150 B.n149 163.367
R732 B.n149 B.n148 163.367
R733 B.n148 B.n121 163.367
R734 B.n144 B.n121 163.367
R735 B.n144 B.n143 163.367
R736 B.n143 B.n142 163.367
R737 B.n142 B.n123 163.367
R738 B.n138 B.n123 163.367
R739 B.n138 B.n137 163.367
R740 B.n137 B.n136 163.367
R741 B.n136 B.n125 163.367
R742 B.n132 B.n125 163.367
R743 B.n132 B.n131 163.367
R744 B.n131 B.n130 163.367
R745 B.n130 B.n127 163.367
R746 B.n127 B.n2 163.367
R747 B.n482 B.n2 163.367
R748 B.n482 B.n481 163.367
R749 B.n481 B.n480 163.367
R750 B.n480 B.n3 163.367
R751 B.n476 B.n3 163.367
R752 B.n476 B.n475 163.367
R753 B.n475 B.n474 163.367
R754 B.n474 B.n5 163.367
R755 B.n470 B.n5 163.367
R756 B.n470 B.n469 163.367
R757 B.n469 B.n468 163.367
R758 B.n468 B.n7 163.367
R759 B.n464 B.n7 163.367
R760 B.n464 B.n463 163.367
R761 B.n463 B.n462 163.367
R762 B.n462 B.n9 163.367
R763 B.n458 B.n9 163.367
R764 B.n458 B.n457 163.367
R765 B.n457 B.n456 163.367
R766 B.n456 B.n11 163.367
R767 B.n452 B.n11 163.367
R768 B.n452 B.n451 163.367
R769 B.n451 B.n450 163.367
R770 B.n450 B.n13 163.367
R771 B.n446 B.n13 163.367
R772 B.n446 B.n445 163.367
R773 B.n445 B.n444 163.367
R774 B.n444 B.n15 163.367
R775 B.n440 B.n15 163.367
R776 B.n440 B.n439 163.367
R777 B.n439 B.n438 163.367
R778 B.n438 B.n17 163.367
R779 B.n434 B.n17 163.367
R780 B.n434 B.n433 163.367
R781 B.n433 B.n432 163.367
R782 B.n432 B.n19 163.367
R783 B.n428 B.n19 163.367
R784 B.n180 B.n109 163.367
R785 B.n184 B.n109 163.367
R786 B.n185 B.n184 163.367
R787 B.n186 B.n185 163.367
R788 B.n186 B.n107 163.367
R789 B.n190 B.n107 163.367
R790 B.n191 B.n190 163.367
R791 B.n192 B.n191 163.367
R792 B.n192 B.n105 163.367
R793 B.n196 B.n105 163.367
R794 B.n197 B.n196 163.367
R795 B.n198 B.n197 163.367
R796 B.n198 B.n103 163.367
R797 B.n202 B.n103 163.367
R798 B.n203 B.n202 163.367
R799 B.n204 B.n203 163.367
R800 B.n204 B.n99 163.367
R801 B.n209 B.n99 163.367
R802 B.n210 B.n209 163.367
R803 B.n211 B.n210 163.367
R804 B.n211 B.n97 163.367
R805 B.n215 B.n97 163.367
R806 B.n216 B.n215 163.367
R807 B.n217 B.n216 163.367
R808 B.n217 B.n95 163.367
R809 B.n221 B.n95 163.367
R810 B.n222 B.n221 163.367
R811 B.n222 B.n91 163.367
R812 B.n226 B.n91 163.367
R813 B.n227 B.n226 163.367
R814 B.n228 B.n227 163.367
R815 B.n228 B.n89 163.367
R816 B.n232 B.n89 163.367
R817 B.n233 B.n232 163.367
R818 B.n234 B.n233 163.367
R819 B.n234 B.n87 163.367
R820 B.n238 B.n87 163.367
R821 B.n239 B.n238 163.367
R822 B.n240 B.n239 163.367
R823 B.n240 B.n85 163.367
R824 B.n244 B.n85 163.367
R825 B.n245 B.n244 163.367
R826 B.n246 B.n245 163.367
R827 B.n246 B.n83 163.367
R828 B.n251 B.n250 163.367
R829 B.n252 B.n251 163.367
R830 B.n252 B.n81 163.367
R831 B.n256 B.n81 163.367
R832 B.n257 B.n256 163.367
R833 B.n258 B.n257 163.367
R834 B.n258 B.n79 163.367
R835 B.n262 B.n79 163.367
R836 B.n263 B.n262 163.367
R837 B.n264 B.n263 163.367
R838 B.n264 B.n77 163.367
R839 B.n268 B.n77 163.367
R840 B.n269 B.n268 163.367
R841 B.n270 B.n269 163.367
R842 B.n270 B.n75 163.367
R843 B.n274 B.n75 163.367
R844 B.n275 B.n274 163.367
R845 B.n276 B.n275 163.367
R846 B.n276 B.n73 163.367
R847 B.n280 B.n73 163.367
R848 B.n281 B.n280 163.367
R849 B.n282 B.n281 163.367
R850 B.n282 B.n71 163.367
R851 B.n286 B.n71 163.367
R852 B.n287 B.n286 163.367
R853 B.n288 B.n287 163.367
R854 B.n288 B.n69 163.367
R855 B.n292 B.n69 163.367
R856 B.n293 B.n292 163.367
R857 B.n294 B.n293 163.367
R858 B.n294 B.n67 163.367
R859 B.n298 B.n67 163.367
R860 B.n299 B.n298 163.367
R861 B.n300 B.n299 163.367
R862 B.n300 B.n65 163.367
R863 B.n304 B.n65 163.367
R864 B.n305 B.n304 163.367
R865 B.n306 B.n305 163.367
R866 B.n306 B.n63 163.367
R867 B.n310 B.n63 163.367
R868 B.n311 B.n310 163.367
R869 B.n312 B.n311 163.367
R870 B.n312 B.n61 163.367
R871 B.n316 B.n61 163.367
R872 B.n317 B.n316 163.367
R873 B.n318 B.n317 163.367
R874 B.n318 B.n59 163.367
R875 B.n322 B.n59 163.367
R876 B.n323 B.n322 163.367
R877 B.n324 B.n323 163.367
R878 B.n324 B.n57 163.367
R879 B.n328 B.n57 163.367
R880 B.n329 B.n328 163.367
R881 B.n330 B.n329 163.367
R882 B.n330 B.n55 163.367
R883 B.n334 B.n55 163.367
R884 B.n335 B.n334 163.367
R885 B.n336 B.n335 163.367
R886 B.n336 B.n53 163.367
R887 B.n340 B.n53 163.367
R888 B.n341 B.n340 163.367
R889 B.n342 B.n341 163.367
R890 B.n342 B.n51 163.367
R891 B.n346 B.n51 163.367
R892 B.n347 B.n346 163.367
R893 B.n348 B.n347 163.367
R894 B.n348 B.n49 163.367
R895 B.n352 B.n49 163.367
R896 B.n353 B.n352 163.367
R897 B.n354 B.n353 163.367
R898 B.n354 B.n47 163.367
R899 B.n358 B.n47 163.367
R900 B.n427 B.n426 163.367
R901 B.n426 B.n21 163.367
R902 B.n422 B.n21 163.367
R903 B.n422 B.n421 163.367
R904 B.n421 B.n420 163.367
R905 B.n420 B.n23 163.367
R906 B.n416 B.n23 163.367
R907 B.n416 B.n415 163.367
R908 B.n415 B.n414 163.367
R909 B.n414 B.n25 163.367
R910 B.n410 B.n25 163.367
R911 B.n410 B.n409 163.367
R912 B.n409 B.n408 163.367
R913 B.n408 B.n27 163.367
R914 B.n404 B.n27 163.367
R915 B.n404 B.n403 163.367
R916 B.n403 B.n402 163.367
R917 B.n402 B.n29 163.367
R918 B.n397 B.n29 163.367
R919 B.n397 B.n396 163.367
R920 B.n396 B.n395 163.367
R921 B.n395 B.n33 163.367
R922 B.n391 B.n33 163.367
R923 B.n391 B.n390 163.367
R924 B.n390 B.n389 163.367
R925 B.n389 B.n35 163.367
R926 B.n384 B.n35 163.367
R927 B.n384 B.n383 163.367
R928 B.n383 B.n382 163.367
R929 B.n382 B.n39 163.367
R930 B.n378 B.n39 163.367
R931 B.n378 B.n377 163.367
R932 B.n377 B.n376 163.367
R933 B.n376 B.n41 163.367
R934 B.n372 B.n41 163.367
R935 B.n372 B.n371 163.367
R936 B.n371 B.n370 163.367
R937 B.n370 B.n43 163.367
R938 B.n366 B.n43 163.367
R939 B.n366 B.n365 163.367
R940 B.n365 B.n364 163.367
R941 B.n364 B.n45 163.367
R942 B.n360 B.n45 163.367
R943 B.n360 B.n359 163.367
R944 B.n94 B.n93 59.5399
R945 B.n207 B.n101 59.5399
R946 B.n400 B.n31 59.5399
R947 B.n386 B.n37 59.5399
R948 B.n429 B.n20 34.1859
R949 B.n357 B.n46 34.1859
R950 B.n249 B.n248 34.1859
R951 B.n181 B.n110 34.1859
R952 B.n93 B.n92 30.6429
R953 B.n101 B.n100 30.6429
R954 B.n31 B.n30 30.6429
R955 B.n37 B.n36 30.6429
R956 B B.n483 18.0485
R957 B.n425 B.n20 10.6151
R958 B.n425 B.n424 10.6151
R959 B.n424 B.n423 10.6151
R960 B.n423 B.n22 10.6151
R961 B.n419 B.n22 10.6151
R962 B.n419 B.n418 10.6151
R963 B.n418 B.n417 10.6151
R964 B.n417 B.n24 10.6151
R965 B.n413 B.n24 10.6151
R966 B.n413 B.n412 10.6151
R967 B.n412 B.n411 10.6151
R968 B.n411 B.n26 10.6151
R969 B.n407 B.n26 10.6151
R970 B.n407 B.n406 10.6151
R971 B.n406 B.n405 10.6151
R972 B.n405 B.n28 10.6151
R973 B.n401 B.n28 10.6151
R974 B.n399 B.n398 10.6151
R975 B.n398 B.n32 10.6151
R976 B.n394 B.n32 10.6151
R977 B.n394 B.n393 10.6151
R978 B.n393 B.n392 10.6151
R979 B.n392 B.n34 10.6151
R980 B.n388 B.n34 10.6151
R981 B.n388 B.n387 10.6151
R982 B.n385 B.n38 10.6151
R983 B.n381 B.n38 10.6151
R984 B.n381 B.n380 10.6151
R985 B.n380 B.n379 10.6151
R986 B.n379 B.n40 10.6151
R987 B.n375 B.n40 10.6151
R988 B.n375 B.n374 10.6151
R989 B.n374 B.n373 10.6151
R990 B.n373 B.n42 10.6151
R991 B.n369 B.n42 10.6151
R992 B.n369 B.n368 10.6151
R993 B.n368 B.n367 10.6151
R994 B.n367 B.n44 10.6151
R995 B.n363 B.n44 10.6151
R996 B.n363 B.n362 10.6151
R997 B.n362 B.n361 10.6151
R998 B.n361 B.n46 10.6151
R999 B.n249 B.n82 10.6151
R1000 B.n253 B.n82 10.6151
R1001 B.n254 B.n253 10.6151
R1002 B.n255 B.n254 10.6151
R1003 B.n255 B.n80 10.6151
R1004 B.n259 B.n80 10.6151
R1005 B.n260 B.n259 10.6151
R1006 B.n261 B.n260 10.6151
R1007 B.n261 B.n78 10.6151
R1008 B.n265 B.n78 10.6151
R1009 B.n266 B.n265 10.6151
R1010 B.n267 B.n266 10.6151
R1011 B.n267 B.n76 10.6151
R1012 B.n271 B.n76 10.6151
R1013 B.n272 B.n271 10.6151
R1014 B.n273 B.n272 10.6151
R1015 B.n273 B.n74 10.6151
R1016 B.n277 B.n74 10.6151
R1017 B.n278 B.n277 10.6151
R1018 B.n279 B.n278 10.6151
R1019 B.n279 B.n72 10.6151
R1020 B.n283 B.n72 10.6151
R1021 B.n284 B.n283 10.6151
R1022 B.n285 B.n284 10.6151
R1023 B.n285 B.n70 10.6151
R1024 B.n289 B.n70 10.6151
R1025 B.n290 B.n289 10.6151
R1026 B.n291 B.n290 10.6151
R1027 B.n291 B.n68 10.6151
R1028 B.n295 B.n68 10.6151
R1029 B.n296 B.n295 10.6151
R1030 B.n297 B.n296 10.6151
R1031 B.n297 B.n66 10.6151
R1032 B.n301 B.n66 10.6151
R1033 B.n302 B.n301 10.6151
R1034 B.n303 B.n302 10.6151
R1035 B.n303 B.n64 10.6151
R1036 B.n307 B.n64 10.6151
R1037 B.n308 B.n307 10.6151
R1038 B.n309 B.n308 10.6151
R1039 B.n309 B.n62 10.6151
R1040 B.n313 B.n62 10.6151
R1041 B.n314 B.n313 10.6151
R1042 B.n315 B.n314 10.6151
R1043 B.n315 B.n60 10.6151
R1044 B.n319 B.n60 10.6151
R1045 B.n320 B.n319 10.6151
R1046 B.n321 B.n320 10.6151
R1047 B.n321 B.n58 10.6151
R1048 B.n325 B.n58 10.6151
R1049 B.n326 B.n325 10.6151
R1050 B.n327 B.n326 10.6151
R1051 B.n327 B.n56 10.6151
R1052 B.n331 B.n56 10.6151
R1053 B.n332 B.n331 10.6151
R1054 B.n333 B.n332 10.6151
R1055 B.n333 B.n54 10.6151
R1056 B.n337 B.n54 10.6151
R1057 B.n338 B.n337 10.6151
R1058 B.n339 B.n338 10.6151
R1059 B.n339 B.n52 10.6151
R1060 B.n343 B.n52 10.6151
R1061 B.n344 B.n343 10.6151
R1062 B.n345 B.n344 10.6151
R1063 B.n345 B.n50 10.6151
R1064 B.n349 B.n50 10.6151
R1065 B.n350 B.n349 10.6151
R1066 B.n351 B.n350 10.6151
R1067 B.n351 B.n48 10.6151
R1068 B.n355 B.n48 10.6151
R1069 B.n356 B.n355 10.6151
R1070 B.n357 B.n356 10.6151
R1071 B.n182 B.n181 10.6151
R1072 B.n183 B.n182 10.6151
R1073 B.n183 B.n108 10.6151
R1074 B.n187 B.n108 10.6151
R1075 B.n188 B.n187 10.6151
R1076 B.n189 B.n188 10.6151
R1077 B.n189 B.n106 10.6151
R1078 B.n193 B.n106 10.6151
R1079 B.n194 B.n193 10.6151
R1080 B.n195 B.n194 10.6151
R1081 B.n195 B.n104 10.6151
R1082 B.n199 B.n104 10.6151
R1083 B.n200 B.n199 10.6151
R1084 B.n201 B.n200 10.6151
R1085 B.n201 B.n102 10.6151
R1086 B.n205 B.n102 10.6151
R1087 B.n206 B.n205 10.6151
R1088 B.n208 B.n98 10.6151
R1089 B.n212 B.n98 10.6151
R1090 B.n213 B.n212 10.6151
R1091 B.n214 B.n213 10.6151
R1092 B.n214 B.n96 10.6151
R1093 B.n218 B.n96 10.6151
R1094 B.n219 B.n218 10.6151
R1095 B.n220 B.n219 10.6151
R1096 B.n224 B.n223 10.6151
R1097 B.n225 B.n224 10.6151
R1098 B.n225 B.n90 10.6151
R1099 B.n229 B.n90 10.6151
R1100 B.n230 B.n229 10.6151
R1101 B.n231 B.n230 10.6151
R1102 B.n231 B.n88 10.6151
R1103 B.n235 B.n88 10.6151
R1104 B.n236 B.n235 10.6151
R1105 B.n237 B.n236 10.6151
R1106 B.n237 B.n86 10.6151
R1107 B.n241 B.n86 10.6151
R1108 B.n242 B.n241 10.6151
R1109 B.n243 B.n242 10.6151
R1110 B.n243 B.n84 10.6151
R1111 B.n247 B.n84 10.6151
R1112 B.n248 B.n247 10.6151
R1113 B.n177 B.n110 10.6151
R1114 B.n177 B.n176 10.6151
R1115 B.n176 B.n175 10.6151
R1116 B.n175 B.n112 10.6151
R1117 B.n171 B.n112 10.6151
R1118 B.n171 B.n170 10.6151
R1119 B.n170 B.n169 10.6151
R1120 B.n169 B.n114 10.6151
R1121 B.n165 B.n114 10.6151
R1122 B.n165 B.n164 10.6151
R1123 B.n164 B.n163 10.6151
R1124 B.n163 B.n116 10.6151
R1125 B.n159 B.n116 10.6151
R1126 B.n159 B.n158 10.6151
R1127 B.n158 B.n157 10.6151
R1128 B.n157 B.n118 10.6151
R1129 B.n153 B.n118 10.6151
R1130 B.n153 B.n152 10.6151
R1131 B.n152 B.n151 10.6151
R1132 B.n151 B.n120 10.6151
R1133 B.n147 B.n120 10.6151
R1134 B.n147 B.n146 10.6151
R1135 B.n146 B.n145 10.6151
R1136 B.n145 B.n122 10.6151
R1137 B.n141 B.n122 10.6151
R1138 B.n141 B.n140 10.6151
R1139 B.n140 B.n139 10.6151
R1140 B.n139 B.n124 10.6151
R1141 B.n135 B.n124 10.6151
R1142 B.n135 B.n134 10.6151
R1143 B.n134 B.n133 10.6151
R1144 B.n133 B.n126 10.6151
R1145 B.n129 B.n126 10.6151
R1146 B.n129 B.n128 10.6151
R1147 B.n128 B.n0 10.6151
R1148 B.n479 B.n1 10.6151
R1149 B.n479 B.n478 10.6151
R1150 B.n478 B.n477 10.6151
R1151 B.n477 B.n4 10.6151
R1152 B.n473 B.n4 10.6151
R1153 B.n473 B.n472 10.6151
R1154 B.n472 B.n471 10.6151
R1155 B.n471 B.n6 10.6151
R1156 B.n467 B.n6 10.6151
R1157 B.n467 B.n466 10.6151
R1158 B.n466 B.n465 10.6151
R1159 B.n465 B.n8 10.6151
R1160 B.n461 B.n8 10.6151
R1161 B.n461 B.n460 10.6151
R1162 B.n460 B.n459 10.6151
R1163 B.n459 B.n10 10.6151
R1164 B.n455 B.n10 10.6151
R1165 B.n455 B.n454 10.6151
R1166 B.n454 B.n453 10.6151
R1167 B.n453 B.n12 10.6151
R1168 B.n449 B.n12 10.6151
R1169 B.n449 B.n448 10.6151
R1170 B.n448 B.n447 10.6151
R1171 B.n447 B.n14 10.6151
R1172 B.n443 B.n14 10.6151
R1173 B.n443 B.n442 10.6151
R1174 B.n442 B.n441 10.6151
R1175 B.n441 B.n16 10.6151
R1176 B.n437 B.n16 10.6151
R1177 B.n437 B.n436 10.6151
R1178 B.n436 B.n435 10.6151
R1179 B.n435 B.n18 10.6151
R1180 B.n431 B.n18 10.6151
R1181 B.n431 B.n430 10.6151
R1182 B.n430 B.n429 10.6151
R1183 B.n400 B.n399 6.5566
R1184 B.n387 B.n386 6.5566
R1185 B.n208 B.n207 6.5566
R1186 B.n220 B.n94 6.5566
R1187 B.n401 B.n400 4.05904
R1188 B.n386 B.n385 4.05904
R1189 B.n207 B.n206 4.05904
R1190 B.n223 B.n94 4.05904
R1191 B.n483 B.n0 2.81026
R1192 B.n483 B.n1 2.81026
C0 VDD1 VP 3.42277f
C1 VDD2 B 1.39485f
C2 VTAIL VN 3.6975f
C3 VP w_n2866_n1754# 5.93083f
C4 VDD2 VP 0.415195f
C5 VDD1 VN 0.154455f
C6 VN w_n2866_n1754# 5.56283f
C7 VP B 1.47057f
C8 VDD2 VN 3.16456f
C9 VDD1 VTAIL 5.88755f
C10 VN B 0.857783f
C11 VTAIL w_n2866_n1754# 1.82797f
C12 VDD2 VTAIL 5.93053f
C13 VDD1 w_n2866_n1754# 1.68429f
C14 VTAIL B 1.47394f
C15 VN VP 4.91639f
C16 VDD2 VDD1 1.3092f
C17 VTAIL VP 3.71172f
C18 VDD1 B 1.32938f
C19 VDD2 w_n2866_n1754# 1.75733f
C20 B w_n2866_n1754# 6.02027f
C21 VDD2 VSUBS 1.161621f
C22 VDD1 VSUBS 1.115676f
C23 VTAIL VSUBS 0.446854f
C24 VN VSUBS 5.22665f
C25 VP VSUBS 2.067677f
C26 B VSUBS 2.854146f
C27 w_n2866_n1754# VSUBS 63.3157f
C28 B.n0 VSUBS 0.004524f
C29 B.n1 VSUBS 0.004524f
C30 B.n2 VSUBS 0.007154f
C31 B.n3 VSUBS 0.007154f
C32 B.n4 VSUBS 0.007154f
C33 B.n5 VSUBS 0.007154f
C34 B.n6 VSUBS 0.007154f
C35 B.n7 VSUBS 0.007154f
C36 B.n8 VSUBS 0.007154f
C37 B.n9 VSUBS 0.007154f
C38 B.n10 VSUBS 0.007154f
C39 B.n11 VSUBS 0.007154f
C40 B.n12 VSUBS 0.007154f
C41 B.n13 VSUBS 0.007154f
C42 B.n14 VSUBS 0.007154f
C43 B.n15 VSUBS 0.007154f
C44 B.n16 VSUBS 0.007154f
C45 B.n17 VSUBS 0.007154f
C46 B.n18 VSUBS 0.007154f
C47 B.n19 VSUBS 0.007154f
C48 B.n20 VSUBS 0.017521f
C49 B.n21 VSUBS 0.007154f
C50 B.n22 VSUBS 0.007154f
C51 B.n23 VSUBS 0.007154f
C52 B.n24 VSUBS 0.007154f
C53 B.n25 VSUBS 0.007154f
C54 B.n26 VSUBS 0.007154f
C55 B.n27 VSUBS 0.007154f
C56 B.n28 VSUBS 0.007154f
C57 B.n29 VSUBS 0.007154f
C58 B.t8 VSUBS 0.058121f
C59 B.t7 VSUBS 0.069782f
C60 B.t6 VSUBS 0.233601f
C61 B.n30 VSUBS 0.126648f
C62 B.n31 VSUBS 0.111024f
C63 B.n32 VSUBS 0.007154f
C64 B.n33 VSUBS 0.007154f
C65 B.n34 VSUBS 0.007154f
C66 B.n35 VSUBS 0.007154f
C67 B.t5 VSUBS 0.058122f
C68 B.t4 VSUBS 0.069783f
C69 B.t3 VSUBS 0.233601f
C70 B.n36 VSUBS 0.126648f
C71 B.n37 VSUBS 0.111023f
C72 B.n38 VSUBS 0.007154f
C73 B.n39 VSUBS 0.007154f
C74 B.n40 VSUBS 0.007154f
C75 B.n41 VSUBS 0.007154f
C76 B.n42 VSUBS 0.007154f
C77 B.n43 VSUBS 0.007154f
C78 B.n44 VSUBS 0.007154f
C79 B.n45 VSUBS 0.007154f
C80 B.n46 VSUBS 0.016713f
C81 B.n47 VSUBS 0.007154f
C82 B.n48 VSUBS 0.007154f
C83 B.n49 VSUBS 0.007154f
C84 B.n50 VSUBS 0.007154f
C85 B.n51 VSUBS 0.007154f
C86 B.n52 VSUBS 0.007154f
C87 B.n53 VSUBS 0.007154f
C88 B.n54 VSUBS 0.007154f
C89 B.n55 VSUBS 0.007154f
C90 B.n56 VSUBS 0.007154f
C91 B.n57 VSUBS 0.007154f
C92 B.n58 VSUBS 0.007154f
C93 B.n59 VSUBS 0.007154f
C94 B.n60 VSUBS 0.007154f
C95 B.n61 VSUBS 0.007154f
C96 B.n62 VSUBS 0.007154f
C97 B.n63 VSUBS 0.007154f
C98 B.n64 VSUBS 0.007154f
C99 B.n65 VSUBS 0.007154f
C100 B.n66 VSUBS 0.007154f
C101 B.n67 VSUBS 0.007154f
C102 B.n68 VSUBS 0.007154f
C103 B.n69 VSUBS 0.007154f
C104 B.n70 VSUBS 0.007154f
C105 B.n71 VSUBS 0.007154f
C106 B.n72 VSUBS 0.007154f
C107 B.n73 VSUBS 0.007154f
C108 B.n74 VSUBS 0.007154f
C109 B.n75 VSUBS 0.007154f
C110 B.n76 VSUBS 0.007154f
C111 B.n77 VSUBS 0.007154f
C112 B.n78 VSUBS 0.007154f
C113 B.n79 VSUBS 0.007154f
C114 B.n80 VSUBS 0.007154f
C115 B.n81 VSUBS 0.007154f
C116 B.n82 VSUBS 0.007154f
C117 B.n83 VSUBS 0.017521f
C118 B.n84 VSUBS 0.007154f
C119 B.n85 VSUBS 0.007154f
C120 B.n86 VSUBS 0.007154f
C121 B.n87 VSUBS 0.007154f
C122 B.n88 VSUBS 0.007154f
C123 B.n89 VSUBS 0.007154f
C124 B.n90 VSUBS 0.007154f
C125 B.n91 VSUBS 0.007154f
C126 B.t10 VSUBS 0.058122f
C127 B.t11 VSUBS 0.069783f
C128 B.t9 VSUBS 0.233601f
C129 B.n92 VSUBS 0.126648f
C130 B.n93 VSUBS 0.111023f
C131 B.n94 VSUBS 0.016576f
C132 B.n95 VSUBS 0.007154f
C133 B.n96 VSUBS 0.007154f
C134 B.n97 VSUBS 0.007154f
C135 B.n98 VSUBS 0.007154f
C136 B.n99 VSUBS 0.007154f
C137 B.t1 VSUBS 0.058121f
C138 B.t2 VSUBS 0.069782f
C139 B.t0 VSUBS 0.233601f
C140 B.n100 VSUBS 0.126648f
C141 B.n101 VSUBS 0.111024f
C142 B.n102 VSUBS 0.007154f
C143 B.n103 VSUBS 0.007154f
C144 B.n104 VSUBS 0.007154f
C145 B.n105 VSUBS 0.007154f
C146 B.n106 VSUBS 0.007154f
C147 B.n107 VSUBS 0.007154f
C148 B.n108 VSUBS 0.007154f
C149 B.n109 VSUBS 0.007154f
C150 B.n110 VSUBS 0.016989f
C151 B.n111 VSUBS 0.007154f
C152 B.n112 VSUBS 0.007154f
C153 B.n113 VSUBS 0.007154f
C154 B.n114 VSUBS 0.007154f
C155 B.n115 VSUBS 0.007154f
C156 B.n116 VSUBS 0.007154f
C157 B.n117 VSUBS 0.007154f
C158 B.n118 VSUBS 0.007154f
C159 B.n119 VSUBS 0.007154f
C160 B.n120 VSUBS 0.007154f
C161 B.n121 VSUBS 0.007154f
C162 B.n122 VSUBS 0.007154f
C163 B.n123 VSUBS 0.007154f
C164 B.n124 VSUBS 0.007154f
C165 B.n125 VSUBS 0.007154f
C166 B.n126 VSUBS 0.007154f
C167 B.n127 VSUBS 0.007154f
C168 B.n128 VSUBS 0.007154f
C169 B.n129 VSUBS 0.007154f
C170 B.n130 VSUBS 0.007154f
C171 B.n131 VSUBS 0.007154f
C172 B.n132 VSUBS 0.007154f
C173 B.n133 VSUBS 0.007154f
C174 B.n134 VSUBS 0.007154f
C175 B.n135 VSUBS 0.007154f
C176 B.n136 VSUBS 0.007154f
C177 B.n137 VSUBS 0.007154f
C178 B.n138 VSUBS 0.007154f
C179 B.n139 VSUBS 0.007154f
C180 B.n140 VSUBS 0.007154f
C181 B.n141 VSUBS 0.007154f
C182 B.n142 VSUBS 0.007154f
C183 B.n143 VSUBS 0.007154f
C184 B.n144 VSUBS 0.007154f
C185 B.n145 VSUBS 0.007154f
C186 B.n146 VSUBS 0.007154f
C187 B.n147 VSUBS 0.007154f
C188 B.n148 VSUBS 0.007154f
C189 B.n149 VSUBS 0.007154f
C190 B.n150 VSUBS 0.007154f
C191 B.n151 VSUBS 0.007154f
C192 B.n152 VSUBS 0.007154f
C193 B.n153 VSUBS 0.007154f
C194 B.n154 VSUBS 0.007154f
C195 B.n155 VSUBS 0.007154f
C196 B.n156 VSUBS 0.007154f
C197 B.n157 VSUBS 0.007154f
C198 B.n158 VSUBS 0.007154f
C199 B.n159 VSUBS 0.007154f
C200 B.n160 VSUBS 0.007154f
C201 B.n161 VSUBS 0.007154f
C202 B.n162 VSUBS 0.007154f
C203 B.n163 VSUBS 0.007154f
C204 B.n164 VSUBS 0.007154f
C205 B.n165 VSUBS 0.007154f
C206 B.n166 VSUBS 0.007154f
C207 B.n167 VSUBS 0.007154f
C208 B.n168 VSUBS 0.007154f
C209 B.n169 VSUBS 0.007154f
C210 B.n170 VSUBS 0.007154f
C211 B.n171 VSUBS 0.007154f
C212 B.n172 VSUBS 0.007154f
C213 B.n173 VSUBS 0.007154f
C214 B.n174 VSUBS 0.007154f
C215 B.n175 VSUBS 0.007154f
C216 B.n176 VSUBS 0.007154f
C217 B.n177 VSUBS 0.007154f
C218 B.n178 VSUBS 0.007154f
C219 B.n179 VSUBS 0.016989f
C220 B.n180 VSUBS 0.017521f
C221 B.n181 VSUBS 0.017521f
C222 B.n182 VSUBS 0.007154f
C223 B.n183 VSUBS 0.007154f
C224 B.n184 VSUBS 0.007154f
C225 B.n185 VSUBS 0.007154f
C226 B.n186 VSUBS 0.007154f
C227 B.n187 VSUBS 0.007154f
C228 B.n188 VSUBS 0.007154f
C229 B.n189 VSUBS 0.007154f
C230 B.n190 VSUBS 0.007154f
C231 B.n191 VSUBS 0.007154f
C232 B.n192 VSUBS 0.007154f
C233 B.n193 VSUBS 0.007154f
C234 B.n194 VSUBS 0.007154f
C235 B.n195 VSUBS 0.007154f
C236 B.n196 VSUBS 0.007154f
C237 B.n197 VSUBS 0.007154f
C238 B.n198 VSUBS 0.007154f
C239 B.n199 VSUBS 0.007154f
C240 B.n200 VSUBS 0.007154f
C241 B.n201 VSUBS 0.007154f
C242 B.n202 VSUBS 0.007154f
C243 B.n203 VSUBS 0.007154f
C244 B.n204 VSUBS 0.007154f
C245 B.n205 VSUBS 0.007154f
C246 B.n206 VSUBS 0.004945f
C247 B.n207 VSUBS 0.016576f
C248 B.n208 VSUBS 0.005787f
C249 B.n209 VSUBS 0.007154f
C250 B.n210 VSUBS 0.007154f
C251 B.n211 VSUBS 0.007154f
C252 B.n212 VSUBS 0.007154f
C253 B.n213 VSUBS 0.007154f
C254 B.n214 VSUBS 0.007154f
C255 B.n215 VSUBS 0.007154f
C256 B.n216 VSUBS 0.007154f
C257 B.n217 VSUBS 0.007154f
C258 B.n218 VSUBS 0.007154f
C259 B.n219 VSUBS 0.007154f
C260 B.n220 VSUBS 0.005787f
C261 B.n221 VSUBS 0.007154f
C262 B.n222 VSUBS 0.007154f
C263 B.n223 VSUBS 0.004945f
C264 B.n224 VSUBS 0.007154f
C265 B.n225 VSUBS 0.007154f
C266 B.n226 VSUBS 0.007154f
C267 B.n227 VSUBS 0.007154f
C268 B.n228 VSUBS 0.007154f
C269 B.n229 VSUBS 0.007154f
C270 B.n230 VSUBS 0.007154f
C271 B.n231 VSUBS 0.007154f
C272 B.n232 VSUBS 0.007154f
C273 B.n233 VSUBS 0.007154f
C274 B.n234 VSUBS 0.007154f
C275 B.n235 VSUBS 0.007154f
C276 B.n236 VSUBS 0.007154f
C277 B.n237 VSUBS 0.007154f
C278 B.n238 VSUBS 0.007154f
C279 B.n239 VSUBS 0.007154f
C280 B.n240 VSUBS 0.007154f
C281 B.n241 VSUBS 0.007154f
C282 B.n242 VSUBS 0.007154f
C283 B.n243 VSUBS 0.007154f
C284 B.n244 VSUBS 0.007154f
C285 B.n245 VSUBS 0.007154f
C286 B.n246 VSUBS 0.007154f
C287 B.n247 VSUBS 0.007154f
C288 B.n248 VSUBS 0.017521f
C289 B.n249 VSUBS 0.016989f
C290 B.n250 VSUBS 0.016989f
C291 B.n251 VSUBS 0.007154f
C292 B.n252 VSUBS 0.007154f
C293 B.n253 VSUBS 0.007154f
C294 B.n254 VSUBS 0.007154f
C295 B.n255 VSUBS 0.007154f
C296 B.n256 VSUBS 0.007154f
C297 B.n257 VSUBS 0.007154f
C298 B.n258 VSUBS 0.007154f
C299 B.n259 VSUBS 0.007154f
C300 B.n260 VSUBS 0.007154f
C301 B.n261 VSUBS 0.007154f
C302 B.n262 VSUBS 0.007154f
C303 B.n263 VSUBS 0.007154f
C304 B.n264 VSUBS 0.007154f
C305 B.n265 VSUBS 0.007154f
C306 B.n266 VSUBS 0.007154f
C307 B.n267 VSUBS 0.007154f
C308 B.n268 VSUBS 0.007154f
C309 B.n269 VSUBS 0.007154f
C310 B.n270 VSUBS 0.007154f
C311 B.n271 VSUBS 0.007154f
C312 B.n272 VSUBS 0.007154f
C313 B.n273 VSUBS 0.007154f
C314 B.n274 VSUBS 0.007154f
C315 B.n275 VSUBS 0.007154f
C316 B.n276 VSUBS 0.007154f
C317 B.n277 VSUBS 0.007154f
C318 B.n278 VSUBS 0.007154f
C319 B.n279 VSUBS 0.007154f
C320 B.n280 VSUBS 0.007154f
C321 B.n281 VSUBS 0.007154f
C322 B.n282 VSUBS 0.007154f
C323 B.n283 VSUBS 0.007154f
C324 B.n284 VSUBS 0.007154f
C325 B.n285 VSUBS 0.007154f
C326 B.n286 VSUBS 0.007154f
C327 B.n287 VSUBS 0.007154f
C328 B.n288 VSUBS 0.007154f
C329 B.n289 VSUBS 0.007154f
C330 B.n290 VSUBS 0.007154f
C331 B.n291 VSUBS 0.007154f
C332 B.n292 VSUBS 0.007154f
C333 B.n293 VSUBS 0.007154f
C334 B.n294 VSUBS 0.007154f
C335 B.n295 VSUBS 0.007154f
C336 B.n296 VSUBS 0.007154f
C337 B.n297 VSUBS 0.007154f
C338 B.n298 VSUBS 0.007154f
C339 B.n299 VSUBS 0.007154f
C340 B.n300 VSUBS 0.007154f
C341 B.n301 VSUBS 0.007154f
C342 B.n302 VSUBS 0.007154f
C343 B.n303 VSUBS 0.007154f
C344 B.n304 VSUBS 0.007154f
C345 B.n305 VSUBS 0.007154f
C346 B.n306 VSUBS 0.007154f
C347 B.n307 VSUBS 0.007154f
C348 B.n308 VSUBS 0.007154f
C349 B.n309 VSUBS 0.007154f
C350 B.n310 VSUBS 0.007154f
C351 B.n311 VSUBS 0.007154f
C352 B.n312 VSUBS 0.007154f
C353 B.n313 VSUBS 0.007154f
C354 B.n314 VSUBS 0.007154f
C355 B.n315 VSUBS 0.007154f
C356 B.n316 VSUBS 0.007154f
C357 B.n317 VSUBS 0.007154f
C358 B.n318 VSUBS 0.007154f
C359 B.n319 VSUBS 0.007154f
C360 B.n320 VSUBS 0.007154f
C361 B.n321 VSUBS 0.007154f
C362 B.n322 VSUBS 0.007154f
C363 B.n323 VSUBS 0.007154f
C364 B.n324 VSUBS 0.007154f
C365 B.n325 VSUBS 0.007154f
C366 B.n326 VSUBS 0.007154f
C367 B.n327 VSUBS 0.007154f
C368 B.n328 VSUBS 0.007154f
C369 B.n329 VSUBS 0.007154f
C370 B.n330 VSUBS 0.007154f
C371 B.n331 VSUBS 0.007154f
C372 B.n332 VSUBS 0.007154f
C373 B.n333 VSUBS 0.007154f
C374 B.n334 VSUBS 0.007154f
C375 B.n335 VSUBS 0.007154f
C376 B.n336 VSUBS 0.007154f
C377 B.n337 VSUBS 0.007154f
C378 B.n338 VSUBS 0.007154f
C379 B.n339 VSUBS 0.007154f
C380 B.n340 VSUBS 0.007154f
C381 B.n341 VSUBS 0.007154f
C382 B.n342 VSUBS 0.007154f
C383 B.n343 VSUBS 0.007154f
C384 B.n344 VSUBS 0.007154f
C385 B.n345 VSUBS 0.007154f
C386 B.n346 VSUBS 0.007154f
C387 B.n347 VSUBS 0.007154f
C388 B.n348 VSUBS 0.007154f
C389 B.n349 VSUBS 0.007154f
C390 B.n350 VSUBS 0.007154f
C391 B.n351 VSUBS 0.007154f
C392 B.n352 VSUBS 0.007154f
C393 B.n353 VSUBS 0.007154f
C394 B.n354 VSUBS 0.007154f
C395 B.n355 VSUBS 0.007154f
C396 B.n356 VSUBS 0.007154f
C397 B.n357 VSUBS 0.017796f
C398 B.n358 VSUBS 0.016989f
C399 B.n359 VSUBS 0.017521f
C400 B.n360 VSUBS 0.007154f
C401 B.n361 VSUBS 0.007154f
C402 B.n362 VSUBS 0.007154f
C403 B.n363 VSUBS 0.007154f
C404 B.n364 VSUBS 0.007154f
C405 B.n365 VSUBS 0.007154f
C406 B.n366 VSUBS 0.007154f
C407 B.n367 VSUBS 0.007154f
C408 B.n368 VSUBS 0.007154f
C409 B.n369 VSUBS 0.007154f
C410 B.n370 VSUBS 0.007154f
C411 B.n371 VSUBS 0.007154f
C412 B.n372 VSUBS 0.007154f
C413 B.n373 VSUBS 0.007154f
C414 B.n374 VSUBS 0.007154f
C415 B.n375 VSUBS 0.007154f
C416 B.n376 VSUBS 0.007154f
C417 B.n377 VSUBS 0.007154f
C418 B.n378 VSUBS 0.007154f
C419 B.n379 VSUBS 0.007154f
C420 B.n380 VSUBS 0.007154f
C421 B.n381 VSUBS 0.007154f
C422 B.n382 VSUBS 0.007154f
C423 B.n383 VSUBS 0.007154f
C424 B.n384 VSUBS 0.007154f
C425 B.n385 VSUBS 0.004945f
C426 B.n386 VSUBS 0.016576f
C427 B.n387 VSUBS 0.005787f
C428 B.n388 VSUBS 0.007154f
C429 B.n389 VSUBS 0.007154f
C430 B.n390 VSUBS 0.007154f
C431 B.n391 VSUBS 0.007154f
C432 B.n392 VSUBS 0.007154f
C433 B.n393 VSUBS 0.007154f
C434 B.n394 VSUBS 0.007154f
C435 B.n395 VSUBS 0.007154f
C436 B.n396 VSUBS 0.007154f
C437 B.n397 VSUBS 0.007154f
C438 B.n398 VSUBS 0.007154f
C439 B.n399 VSUBS 0.005787f
C440 B.n400 VSUBS 0.016576f
C441 B.n401 VSUBS 0.004945f
C442 B.n402 VSUBS 0.007154f
C443 B.n403 VSUBS 0.007154f
C444 B.n404 VSUBS 0.007154f
C445 B.n405 VSUBS 0.007154f
C446 B.n406 VSUBS 0.007154f
C447 B.n407 VSUBS 0.007154f
C448 B.n408 VSUBS 0.007154f
C449 B.n409 VSUBS 0.007154f
C450 B.n410 VSUBS 0.007154f
C451 B.n411 VSUBS 0.007154f
C452 B.n412 VSUBS 0.007154f
C453 B.n413 VSUBS 0.007154f
C454 B.n414 VSUBS 0.007154f
C455 B.n415 VSUBS 0.007154f
C456 B.n416 VSUBS 0.007154f
C457 B.n417 VSUBS 0.007154f
C458 B.n418 VSUBS 0.007154f
C459 B.n419 VSUBS 0.007154f
C460 B.n420 VSUBS 0.007154f
C461 B.n421 VSUBS 0.007154f
C462 B.n422 VSUBS 0.007154f
C463 B.n423 VSUBS 0.007154f
C464 B.n424 VSUBS 0.007154f
C465 B.n425 VSUBS 0.007154f
C466 B.n426 VSUBS 0.007154f
C467 B.n427 VSUBS 0.017521f
C468 B.n428 VSUBS 0.016989f
C469 B.n429 VSUBS 0.016989f
C470 B.n430 VSUBS 0.007154f
C471 B.n431 VSUBS 0.007154f
C472 B.n432 VSUBS 0.007154f
C473 B.n433 VSUBS 0.007154f
C474 B.n434 VSUBS 0.007154f
C475 B.n435 VSUBS 0.007154f
C476 B.n436 VSUBS 0.007154f
C477 B.n437 VSUBS 0.007154f
C478 B.n438 VSUBS 0.007154f
C479 B.n439 VSUBS 0.007154f
C480 B.n440 VSUBS 0.007154f
C481 B.n441 VSUBS 0.007154f
C482 B.n442 VSUBS 0.007154f
C483 B.n443 VSUBS 0.007154f
C484 B.n444 VSUBS 0.007154f
C485 B.n445 VSUBS 0.007154f
C486 B.n446 VSUBS 0.007154f
C487 B.n447 VSUBS 0.007154f
C488 B.n448 VSUBS 0.007154f
C489 B.n449 VSUBS 0.007154f
C490 B.n450 VSUBS 0.007154f
C491 B.n451 VSUBS 0.007154f
C492 B.n452 VSUBS 0.007154f
C493 B.n453 VSUBS 0.007154f
C494 B.n454 VSUBS 0.007154f
C495 B.n455 VSUBS 0.007154f
C496 B.n456 VSUBS 0.007154f
C497 B.n457 VSUBS 0.007154f
C498 B.n458 VSUBS 0.007154f
C499 B.n459 VSUBS 0.007154f
C500 B.n460 VSUBS 0.007154f
C501 B.n461 VSUBS 0.007154f
C502 B.n462 VSUBS 0.007154f
C503 B.n463 VSUBS 0.007154f
C504 B.n464 VSUBS 0.007154f
C505 B.n465 VSUBS 0.007154f
C506 B.n466 VSUBS 0.007154f
C507 B.n467 VSUBS 0.007154f
C508 B.n468 VSUBS 0.007154f
C509 B.n469 VSUBS 0.007154f
C510 B.n470 VSUBS 0.007154f
C511 B.n471 VSUBS 0.007154f
C512 B.n472 VSUBS 0.007154f
C513 B.n473 VSUBS 0.007154f
C514 B.n474 VSUBS 0.007154f
C515 B.n475 VSUBS 0.007154f
C516 B.n476 VSUBS 0.007154f
C517 B.n477 VSUBS 0.007154f
C518 B.n478 VSUBS 0.007154f
C519 B.n479 VSUBS 0.007154f
C520 B.n480 VSUBS 0.007154f
C521 B.n481 VSUBS 0.007154f
C522 B.n482 VSUBS 0.007154f
C523 B.n483 VSUBS 0.0162f
C524 VDD1.n0 VSUBS 0.025515f
C525 VDD1.n1 VSUBS 0.023583f
C526 VDD1.n2 VSUBS 0.012673f
C527 VDD1.n3 VSUBS 0.029954f
C528 VDD1.n4 VSUBS 0.013418f
C529 VDD1.n5 VSUBS 0.091204f
C530 VDD1.t5 VSUBS 0.066153f
C531 VDD1.n6 VSUBS 0.022465f
C532 VDD1.n7 VSUBS 0.01884f
C533 VDD1.n8 VSUBS 0.012673f
C534 VDD1.n9 VSUBS 0.316244f
C535 VDD1.n10 VSUBS 0.023583f
C536 VDD1.n11 VSUBS 0.012673f
C537 VDD1.n12 VSUBS 0.013418f
C538 VDD1.n13 VSUBS 0.029954f
C539 VDD1.n14 VSUBS 0.071157f
C540 VDD1.n15 VSUBS 0.013418f
C541 VDD1.n16 VSUBS 0.012673f
C542 VDD1.n17 VSUBS 0.057412f
C543 VDD1.n18 VSUBS 0.05602f
C544 VDD1.t3 VSUBS 0.073241f
C545 VDD1.t6 VSUBS 0.073241f
C546 VDD1.n19 VSUBS 0.425639f
C547 VDD1.n20 VSUBS 0.611705f
C548 VDD1.n21 VSUBS 0.025515f
C549 VDD1.n22 VSUBS 0.023583f
C550 VDD1.n23 VSUBS 0.012673f
C551 VDD1.n24 VSUBS 0.029954f
C552 VDD1.n25 VSUBS 0.013418f
C553 VDD1.n26 VSUBS 0.091204f
C554 VDD1.t0 VSUBS 0.066153f
C555 VDD1.n27 VSUBS 0.022465f
C556 VDD1.n28 VSUBS 0.01884f
C557 VDD1.n29 VSUBS 0.012673f
C558 VDD1.n30 VSUBS 0.316245f
C559 VDD1.n31 VSUBS 0.023583f
C560 VDD1.n32 VSUBS 0.012673f
C561 VDD1.n33 VSUBS 0.013418f
C562 VDD1.n34 VSUBS 0.029954f
C563 VDD1.n35 VSUBS 0.071157f
C564 VDD1.n36 VSUBS 0.013418f
C565 VDD1.n37 VSUBS 0.012673f
C566 VDD1.n38 VSUBS 0.057412f
C567 VDD1.n39 VSUBS 0.05602f
C568 VDD1.t1 VSUBS 0.073241f
C569 VDD1.t2 VSUBS 0.073241f
C570 VDD1.n40 VSUBS 0.425637f
C571 VDD1.n41 VSUBS 0.604997f
C572 VDD1.t9 VSUBS 0.073241f
C573 VDD1.t4 VSUBS 0.073241f
C574 VDD1.n42 VSUBS 0.429944f
C575 VDD1.n43 VSUBS 1.83798f
C576 VDD1.t7 VSUBS 0.073241f
C577 VDD1.t8 VSUBS 0.073241f
C578 VDD1.n44 VSUBS 0.425637f
C579 VDD1.n45 VSUBS 2.00297f
C580 VP.n0 VSUBS 0.073636f
C581 VP.t0 VSUBS 0.695284f
C582 VP.n1 VSUBS 0.304018f
C583 VP.n2 VSUBS 0.055184f
C584 VP.t7 VSUBS 0.695284f
C585 VP.n3 VSUBS 0.304018f
C586 VP.n4 VSUBS 0.055184f
C587 VP.t8 VSUBS 0.695284f
C588 VP.n5 VSUBS 0.304018f
C589 VP.n6 VSUBS 0.073636f
C590 VP.n7 VSUBS 0.073636f
C591 VP.t1 VSUBS 0.800962f
C592 VP.t2 VSUBS 0.695284f
C593 VP.n8 VSUBS 0.304018f
C594 VP.n9 VSUBS 0.055184f
C595 VP.t3 VSUBS 0.695284f
C596 VP.n10 VSUBS 0.304018f
C597 VP.n11 VSUBS 0.055184f
C598 VP.t6 VSUBS 0.695284f
C599 VP.n12 VSUBS 0.381999f
C600 VP.t4 VSUBS 0.871223f
C601 VP.n13 VSUBS 0.393231f
C602 VP.n14 VSUBS 0.292594f
C603 VP.n15 VSUBS 0.089681f
C604 VP.n16 VSUBS 0.045756f
C605 VP.n17 VSUBS 0.085876f
C606 VP.n18 VSUBS 0.055184f
C607 VP.n19 VSUBS 0.055184f
C608 VP.n20 VSUBS 0.085876f
C609 VP.n21 VSUBS 0.045756f
C610 VP.n22 VSUBS 0.089681f
C611 VP.n23 VSUBS 0.055184f
C612 VP.n24 VSUBS 0.055184f
C613 VP.n25 VSUBS 0.075643f
C614 VP.n26 VSUBS 0.049378f
C615 VP.n27 VSUBS 0.413734f
C616 VP.n28 VSUBS 2.10511f
C617 VP.n29 VSUBS 2.15486f
C618 VP.t9 VSUBS 0.800962f
C619 VP.n30 VSUBS 0.413734f
C620 VP.n31 VSUBS 0.049378f
C621 VP.n32 VSUBS 0.075643f
C622 VP.n33 VSUBS 0.055184f
C623 VP.n34 VSUBS 0.055184f
C624 VP.n35 VSUBS 0.089681f
C625 VP.n36 VSUBS 0.045756f
C626 VP.n37 VSUBS 0.085876f
C627 VP.n38 VSUBS 0.055184f
C628 VP.n39 VSUBS 0.055184f
C629 VP.n40 VSUBS 0.085876f
C630 VP.n41 VSUBS 0.045756f
C631 VP.n42 VSUBS 0.089681f
C632 VP.n43 VSUBS 0.055184f
C633 VP.n44 VSUBS 0.055184f
C634 VP.n45 VSUBS 0.075643f
C635 VP.n46 VSUBS 0.049378f
C636 VP.t5 VSUBS 0.800962f
C637 VP.n47 VSUBS 0.413734f
C638 VP.n48 VSUBS 0.051682f
C639 VTAIL.t15 VSUBS 0.090101f
C640 VTAIL.t13 VSUBS 0.090101f
C641 VTAIL.n0 VSUBS 0.455639f
C642 VTAIL.n1 VSUBS 0.6446f
C643 VTAIL.n2 VSUBS 0.031388f
C644 VTAIL.n3 VSUBS 0.029012f
C645 VTAIL.n4 VSUBS 0.01559f
C646 VTAIL.n5 VSUBS 0.036849f
C647 VTAIL.n6 VSUBS 0.016507f
C648 VTAIL.n7 VSUBS 0.112199f
C649 VTAIL.t4 VSUBS 0.081381f
C650 VTAIL.n8 VSUBS 0.027637f
C651 VTAIL.n9 VSUBS 0.023177f
C652 VTAIL.n10 VSUBS 0.01559f
C653 VTAIL.n11 VSUBS 0.389042f
C654 VTAIL.n12 VSUBS 0.029012f
C655 VTAIL.n13 VSUBS 0.01559f
C656 VTAIL.n14 VSUBS 0.016507f
C657 VTAIL.n15 VSUBS 0.036849f
C658 VTAIL.n16 VSUBS 0.087537f
C659 VTAIL.n17 VSUBS 0.016507f
C660 VTAIL.n18 VSUBS 0.01559f
C661 VTAIL.n19 VSUBS 0.070628f
C662 VTAIL.n20 VSUBS 0.044055f
C663 VTAIL.n21 VSUBS 0.261714f
C664 VTAIL.t6 VSUBS 0.090101f
C665 VTAIL.t8 VSUBS 0.090101f
C666 VTAIL.n22 VSUBS 0.455639f
C667 VTAIL.n23 VSUBS 0.690738f
C668 VTAIL.t2 VSUBS 0.090101f
C669 VTAIL.t1 VSUBS 0.090101f
C670 VTAIL.n24 VSUBS 0.455639f
C671 VTAIL.n25 VSUBS 1.52889f
C672 VTAIL.t16 VSUBS 0.090101f
C673 VTAIL.t19 VSUBS 0.090101f
C674 VTAIL.n26 VSUBS 0.455642f
C675 VTAIL.n27 VSUBS 1.52888f
C676 VTAIL.t18 VSUBS 0.090101f
C677 VTAIL.t17 VSUBS 0.090101f
C678 VTAIL.n28 VSUBS 0.455642f
C679 VTAIL.n29 VSUBS 0.690735f
C680 VTAIL.n30 VSUBS 0.031388f
C681 VTAIL.n31 VSUBS 0.029012f
C682 VTAIL.n32 VSUBS 0.01559f
C683 VTAIL.n33 VSUBS 0.036849f
C684 VTAIL.n34 VSUBS 0.016507f
C685 VTAIL.n35 VSUBS 0.112199f
C686 VTAIL.t14 VSUBS 0.081381f
C687 VTAIL.n36 VSUBS 0.027637f
C688 VTAIL.n37 VSUBS 0.023177f
C689 VTAIL.n38 VSUBS 0.01559f
C690 VTAIL.n39 VSUBS 0.389042f
C691 VTAIL.n40 VSUBS 0.029012f
C692 VTAIL.n41 VSUBS 0.01559f
C693 VTAIL.n42 VSUBS 0.016507f
C694 VTAIL.n43 VSUBS 0.036849f
C695 VTAIL.n44 VSUBS 0.087537f
C696 VTAIL.n45 VSUBS 0.016507f
C697 VTAIL.n46 VSUBS 0.01559f
C698 VTAIL.n47 VSUBS 0.070628f
C699 VTAIL.n48 VSUBS 0.044055f
C700 VTAIL.n49 VSUBS 0.261714f
C701 VTAIL.t7 VSUBS 0.090101f
C702 VTAIL.t9 VSUBS 0.090101f
C703 VTAIL.n50 VSUBS 0.455642f
C704 VTAIL.n51 VSUBS 0.67099f
C705 VTAIL.t5 VSUBS 0.090101f
C706 VTAIL.t0 VSUBS 0.090101f
C707 VTAIL.n52 VSUBS 0.455642f
C708 VTAIL.n53 VSUBS 0.690735f
C709 VTAIL.n54 VSUBS 0.031388f
C710 VTAIL.n55 VSUBS 0.029012f
C711 VTAIL.n56 VSUBS 0.01559f
C712 VTAIL.n57 VSUBS 0.036849f
C713 VTAIL.n58 VSUBS 0.016507f
C714 VTAIL.n59 VSUBS 0.112199f
C715 VTAIL.t3 VSUBS 0.081381f
C716 VTAIL.n60 VSUBS 0.027637f
C717 VTAIL.n61 VSUBS 0.023177f
C718 VTAIL.n62 VSUBS 0.01559f
C719 VTAIL.n63 VSUBS 0.389042f
C720 VTAIL.n64 VSUBS 0.029012f
C721 VTAIL.n65 VSUBS 0.01559f
C722 VTAIL.n66 VSUBS 0.016507f
C723 VTAIL.n67 VSUBS 0.036849f
C724 VTAIL.n68 VSUBS 0.087537f
C725 VTAIL.n69 VSUBS 0.016507f
C726 VTAIL.n70 VSUBS 0.01559f
C727 VTAIL.n71 VSUBS 0.070628f
C728 VTAIL.n72 VSUBS 0.044055f
C729 VTAIL.n73 VSUBS 0.992274f
C730 VTAIL.n74 VSUBS 0.031388f
C731 VTAIL.n75 VSUBS 0.029012f
C732 VTAIL.n76 VSUBS 0.01559f
C733 VTAIL.n77 VSUBS 0.036849f
C734 VTAIL.n78 VSUBS 0.016507f
C735 VTAIL.n79 VSUBS 0.112199f
C736 VTAIL.t10 VSUBS 0.081381f
C737 VTAIL.n80 VSUBS 0.027637f
C738 VTAIL.n81 VSUBS 0.023177f
C739 VTAIL.n82 VSUBS 0.01559f
C740 VTAIL.n83 VSUBS 0.389042f
C741 VTAIL.n84 VSUBS 0.029012f
C742 VTAIL.n85 VSUBS 0.01559f
C743 VTAIL.n86 VSUBS 0.016507f
C744 VTAIL.n87 VSUBS 0.036849f
C745 VTAIL.n88 VSUBS 0.087537f
C746 VTAIL.n89 VSUBS 0.016507f
C747 VTAIL.n90 VSUBS 0.01559f
C748 VTAIL.n91 VSUBS 0.070628f
C749 VTAIL.n92 VSUBS 0.044055f
C750 VTAIL.n93 VSUBS 0.992274f
C751 VTAIL.t11 VSUBS 0.090101f
C752 VTAIL.t12 VSUBS 0.090101f
C753 VTAIL.n94 VSUBS 0.455639f
C754 VTAIL.n95 VSUBS 0.589799f
C755 VDD2.n0 VSUBS 0.025202f
C756 VDD2.n1 VSUBS 0.023294f
C757 VDD2.n2 VSUBS 0.012517f
C758 VDD2.n3 VSUBS 0.029587f
C759 VDD2.n4 VSUBS 0.013254f
C760 VDD2.n5 VSUBS 0.090086f
C761 VDD2.t7 VSUBS 0.065342f
C762 VDD2.n6 VSUBS 0.02219f
C763 VDD2.n7 VSUBS 0.01861f
C764 VDD2.n8 VSUBS 0.012517f
C765 VDD2.n9 VSUBS 0.312369f
C766 VDD2.n10 VSUBS 0.023294f
C767 VDD2.n11 VSUBS 0.012517f
C768 VDD2.n12 VSUBS 0.013254f
C769 VDD2.n13 VSUBS 0.029587f
C770 VDD2.n14 VSUBS 0.070285f
C771 VDD2.n15 VSUBS 0.013254f
C772 VDD2.n16 VSUBS 0.012517f
C773 VDD2.n17 VSUBS 0.056708f
C774 VDD2.n18 VSUBS 0.055333f
C775 VDD2.t3 VSUBS 0.072344f
C776 VDD2.t8 VSUBS 0.072344f
C777 VDD2.n19 VSUBS 0.420421f
C778 VDD2.n20 VSUBS 0.597583f
C779 VDD2.t2 VSUBS 0.072344f
C780 VDD2.t5 VSUBS 0.072344f
C781 VDD2.n21 VSUBS 0.424675f
C782 VDD2.n22 VSUBS 1.73598f
C783 VDD2.n23 VSUBS 0.025202f
C784 VDD2.n24 VSUBS 0.023294f
C785 VDD2.n25 VSUBS 0.012517f
C786 VDD2.n26 VSUBS 0.029587f
C787 VDD2.n27 VSUBS 0.013254f
C788 VDD2.n28 VSUBS 0.090086f
C789 VDD2.t0 VSUBS 0.065342f
C790 VDD2.n29 VSUBS 0.02219f
C791 VDD2.n30 VSUBS 0.01861f
C792 VDD2.n31 VSUBS 0.012517f
C793 VDD2.n32 VSUBS 0.312369f
C794 VDD2.n33 VSUBS 0.023294f
C795 VDD2.n34 VSUBS 0.012517f
C796 VDD2.n35 VSUBS 0.013254f
C797 VDD2.n36 VSUBS 0.029587f
C798 VDD2.n37 VSUBS 0.070285f
C799 VDD2.n38 VSUBS 0.013254f
C800 VDD2.n39 VSUBS 0.012517f
C801 VDD2.n40 VSUBS 0.056708f
C802 VDD2.n41 VSUBS 0.051435f
C803 VDD2.n42 VSUBS 1.60945f
C804 VDD2.t9 VSUBS 0.072344f
C805 VDD2.t6 VSUBS 0.072344f
C806 VDD2.n43 VSUBS 0.420423f
C807 VDD2.n44 VSUBS 0.459375f
C808 VDD2.t1 VSUBS 0.072344f
C809 VDD2.t4 VSUBS 0.072344f
C810 VDD2.n45 VSUBS 0.424656f
C811 VN.n0 VSUBS 0.07127f
C812 VN.t7 VSUBS 0.672946f
C813 VN.n1 VSUBS 0.29425f
C814 VN.n2 VSUBS 0.053411f
C815 VN.t8 VSUBS 0.672946f
C816 VN.n3 VSUBS 0.29425f
C817 VN.n4 VSUBS 0.053411f
C818 VN.t6 VSUBS 0.672946f
C819 VN.n5 VSUBS 0.369726f
C820 VN.t4 VSUBS 0.843232f
C821 VN.n6 VSUBS 0.380598f
C822 VN.n7 VSUBS 0.283193f
C823 VN.n8 VSUBS 0.0868f
C824 VN.n9 VSUBS 0.044285f
C825 VN.n10 VSUBS 0.083117f
C826 VN.n11 VSUBS 0.053411f
C827 VN.n12 VSUBS 0.053411f
C828 VN.n13 VSUBS 0.083117f
C829 VN.n14 VSUBS 0.044285f
C830 VN.n15 VSUBS 0.0868f
C831 VN.n16 VSUBS 0.053411f
C832 VN.n17 VSUBS 0.053411f
C833 VN.n18 VSUBS 0.073213f
C834 VN.n19 VSUBS 0.047791f
C835 VN.t9 VSUBS 0.775229f
C836 VN.n20 VSUBS 0.400441f
C837 VN.n21 VSUBS 0.050021f
C838 VN.n22 VSUBS 0.07127f
C839 VN.t0 VSUBS 0.672946f
C840 VN.n23 VSUBS 0.29425f
C841 VN.n24 VSUBS 0.053411f
C842 VN.t1 VSUBS 0.672946f
C843 VN.n25 VSUBS 0.29425f
C844 VN.n26 VSUBS 0.053411f
C845 VN.t2 VSUBS 0.672946f
C846 VN.n27 VSUBS 0.369726f
C847 VN.t5 VSUBS 0.843232f
C848 VN.n28 VSUBS 0.380598f
C849 VN.n29 VSUBS 0.283193f
C850 VN.n30 VSUBS 0.0868f
C851 VN.n31 VSUBS 0.044285f
C852 VN.n32 VSUBS 0.083117f
C853 VN.n33 VSUBS 0.053411f
C854 VN.n34 VSUBS 0.053411f
C855 VN.n35 VSUBS 0.083117f
C856 VN.n36 VSUBS 0.044285f
C857 VN.n37 VSUBS 0.0868f
C858 VN.n38 VSUBS 0.053411f
C859 VN.n39 VSUBS 0.053411f
C860 VN.n40 VSUBS 0.073213f
C861 VN.n41 VSUBS 0.047791f
C862 VN.t3 VSUBS 0.775229f
C863 VN.n42 VSUBS 0.400441f
C864 VN.n43 VSUBS 2.06773f
.ends

