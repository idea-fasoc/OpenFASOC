* NGSPICE file created from diff_pair_sample_1182.ext - technology: sky130A

.subckt diff_pair_sample_1182 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=0 ps=0 w=16.09 l=2.69
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=6.2751 ps=32.96 w=16.09 l=2.69
X2 VDD2.t0 VN.t1 VTAIL.t2 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=6.2751 ps=32.96 w=16.09 l=2.69
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=6.2751 ps=32.96 w=16.09 l=2.69
X4 B.t8 B.t6 B.t7 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=0 ps=0 w=16.09 l=2.69
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=6.2751 ps=32.96 w=16.09 l=2.69
X6 B.t5 B.t3 B.t4 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=0 ps=0 w=16.09 l=2.69
X7 B.t2 B.t0 B.t1 w_n2178_n4186# sky130_fd_pr__pfet_01v8 ad=6.2751 pd=32.96 as=0 ps=0 w=16.09 l=2.69
R0 B.n475 B.n474 585
R1 B.n476 B.n77 585
R2 B.n478 B.n477 585
R3 B.n479 B.n76 585
R4 B.n481 B.n480 585
R5 B.n482 B.n75 585
R6 B.n484 B.n483 585
R7 B.n485 B.n74 585
R8 B.n487 B.n486 585
R9 B.n488 B.n73 585
R10 B.n490 B.n489 585
R11 B.n491 B.n72 585
R12 B.n493 B.n492 585
R13 B.n494 B.n71 585
R14 B.n496 B.n495 585
R15 B.n497 B.n70 585
R16 B.n499 B.n498 585
R17 B.n500 B.n69 585
R18 B.n502 B.n501 585
R19 B.n503 B.n68 585
R20 B.n505 B.n504 585
R21 B.n506 B.n67 585
R22 B.n508 B.n507 585
R23 B.n509 B.n66 585
R24 B.n511 B.n510 585
R25 B.n512 B.n65 585
R26 B.n514 B.n513 585
R27 B.n515 B.n64 585
R28 B.n517 B.n516 585
R29 B.n518 B.n63 585
R30 B.n520 B.n519 585
R31 B.n521 B.n62 585
R32 B.n523 B.n522 585
R33 B.n524 B.n61 585
R34 B.n526 B.n525 585
R35 B.n527 B.n60 585
R36 B.n529 B.n528 585
R37 B.n530 B.n59 585
R38 B.n532 B.n531 585
R39 B.n533 B.n58 585
R40 B.n535 B.n534 585
R41 B.n536 B.n57 585
R42 B.n538 B.n537 585
R43 B.n539 B.n56 585
R44 B.n541 B.n540 585
R45 B.n542 B.n55 585
R46 B.n544 B.n543 585
R47 B.n545 B.n54 585
R48 B.n547 B.n546 585
R49 B.n548 B.n53 585
R50 B.n550 B.n549 585
R51 B.n551 B.n52 585
R52 B.n553 B.n552 585
R53 B.n554 B.n49 585
R54 B.n557 B.n556 585
R55 B.n558 B.n48 585
R56 B.n560 B.n559 585
R57 B.n561 B.n47 585
R58 B.n563 B.n562 585
R59 B.n564 B.n46 585
R60 B.n566 B.n565 585
R61 B.n567 B.n45 585
R62 B.n569 B.n568 585
R63 B.n571 B.n570 585
R64 B.n572 B.n41 585
R65 B.n574 B.n573 585
R66 B.n575 B.n40 585
R67 B.n577 B.n576 585
R68 B.n578 B.n39 585
R69 B.n580 B.n579 585
R70 B.n581 B.n38 585
R71 B.n583 B.n582 585
R72 B.n584 B.n37 585
R73 B.n586 B.n585 585
R74 B.n587 B.n36 585
R75 B.n589 B.n588 585
R76 B.n590 B.n35 585
R77 B.n592 B.n591 585
R78 B.n593 B.n34 585
R79 B.n595 B.n594 585
R80 B.n596 B.n33 585
R81 B.n598 B.n597 585
R82 B.n599 B.n32 585
R83 B.n601 B.n600 585
R84 B.n602 B.n31 585
R85 B.n604 B.n603 585
R86 B.n605 B.n30 585
R87 B.n607 B.n606 585
R88 B.n608 B.n29 585
R89 B.n610 B.n609 585
R90 B.n611 B.n28 585
R91 B.n613 B.n612 585
R92 B.n614 B.n27 585
R93 B.n616 B.n615 585
R94 B.n617 B.n26 585
R95 B.n619 B.n618 585
R96 B.n620 B.n25 585
R97 B.n622 B.n621 585
R98 B.n623 B.n24 585
R99 B.n625 B.n624 585
R100 B.n626 B.n23 585
R101 B.n628 B.n627 585
R102 B.n629 B.n22 585
R103 B.n631 B.n630 585
R104 B.n632 B.n21 585
R105 B.n634 B.n633 585
R106 B.n635 B.n20 585
R107 B.n637 B.n636 585
R108 B.n638 B.n19 585
R109 B.n640 B.n639 585
R110 B.n641 B.n18 585
R111 B.n643 B.n642 585
R112 B.n644 B.n17 585
R113 B.n646 B.n645 585
R114 B.n647 B.n16 585
R115 B.n649 B.n648 585
R116 B.n650 B.n15 585
R117 B.n473 B.n78 585
R118 B.n472 B.n471 585
R119 B.n470 B.n79 585
R120 B.n469 B.n468 585
R121 B.n467 B.n80 585
R122 B.n466 B.n465 585
R123 B.n464 B.n81 585
R124 B.n463 B.n462 585
R125 B.n461 B.n82 585
R126 B.n460 B.n459 585
R127 B.n458 B.n83 585
R128 B.n457 B.n456 585
R129 B.n455 B.n84 585
R130 B.n454 B.n453 585
R131 B.n452 B.n85 585
R132 B.n451 B.n450 585
R133 B.n449 B.n86 585
R134 B.n448 B.n447 585
R135 B.n446 B.n87 585
R136 B.n445 B.n444 585
R137 B.n443 B.n88 585
R138 B.n442 B.n441 585
R139 B.n440 B.n89 585
R140 B.n439 B.n438 585
R141 B.n437 B.n90 585
R142 B.n436 B.n435 585
R143 B.n434 B.n91 585
R144 B.n433 B.n432 585
R145 B.n431 B.n92 585
R146 B.n430 B.n429 585
R147 B.n428 B.n93 585
R148 B.n427 B.n426 585
R149 B.n425 B.n94 585
R150 B.n424 B.n423 585
R151 B.n422 B.n95 585
R152 B.n421 B.n420 585
R153 B.n419 B.n96 585
R154 B.n418 B.n417 585
R155 B.n416 B.n97 585
R156 B.n415 B.n414 585
R157 B.n413 B.n98 585
R158 B.n412 B.n411 585
R159 B.n410 B.n99 585
R160 B.n409 B.n408 585
R161 B.n407 B.n100 585
R162 B.n406 B.n405 585
R163 B.n404 B.n101 585
R164 B.n403 B.n402 585
R165 B.n401 B.n102 585
R166 B.n400 B.n399 585
R167 B.n398 B.n103 585
R168 B.n397 B.n396 585
R169 B.n395 B.n104 585
R170 B.n218 B.n167 585
R171 B.n220 B.n219 585
R172 B.n221 B.n166 585
R173 B.n223 B.n222 585
R174 B.n224 B.n165 585
R175 B.n226 B.n225 585
R176 B.n227 B.n164 585
R177 B.n229 B.n228 585
R178 B.n230 B.n163 585
R179 B.n232 B.n231 585
R180 B.n233 B.n162 585
R181 B.n235 B.n234 585
R182 B.n236 B.n161 585
R183 B.n238 B.n237 585
R184 B.n239 B.n160 585
R185 B.n241 B.n240 585
R186 B.n242 B.n159 585
R187 B.n244 B.n243 585
R188 B.n245 B.n158 585
R189 B.n247 B.n246 585
R190 B.n248 B.n157 585
R191 B.n250 B.n249 585
R192 B.n251 B.n156 585
R193 B.n253 B.n252 585
R194 B.n254 B.n155 585
R195 B.n256 B.n255 585
R196 B.n257 B.n154 585
R197 B.n259 B.n258 585
R198 B.n260 B.n153 585
R199 B.n262 B.n261 585
R200 B.n263 B.n152 585
R201 B.n265 B.n264 585
R202 B.n266 B.n151 585
R203 B.n268 B.n267 585
R204 B.n269 B.n150 585
R205 B.n271 B.n270 585
R206 B.n272 B.n149 585
R207 B.n274 B.n273 585
R208 B.n275 B.n148 585
R209 B.n277 B.n276 585
R210 B.n278 B.n147 585
R211 B.n280 B.n279 585
R212 B.n281 B.n146 585
R213 B.n283 B.n282 585
R214 B.n284 B.n145 585
R215 B.n286 B.n285 585
R216 B.n287 B.n144 585
R217 B.n289 B.n288 585
R218 B.n290 B.n143 585
R219 B.n292 B.n291 585
R220 B.n293 B.n142 585
R221 B.n295 B.n294 585
R222 B.n296 B.n141 585
R223 B.n298 B.n297 585
R224 B.n300 B.n299 585
R225 B.n301 B.n137 585
R226 B.n303 B.n302 585
R227 B.n304 B.n136 585
R228 B.n306 B.n305 585
R229 B.n307 B.n135 585
R230 B.n309 B.n308 585
R231 B.n310 B.n134 585
R232 B.n312 B.n311 585
R233 B.n314 B.n131 585
R234 B.n316 B.n315 585
R235 B.n317 B.n130 585
R236 B.n319 B.n318 585
R237 B.n320 B.n129 585
R238 B.n322 B.n321 585
R239 B.n323 B.n128 585
R240 B.n325 B.n324 585
R241 B.n326 B.n127 585
R242 B.n328 B.n327 585
R243 B.n329 B.n126 585
R244 B.n331 B.n330 585
R245 B.n332 B.n125 585
R246 B.n334 B.n333 585
R247 B.n335 B.n124 585
R248 B.n337 B.n336 585
R249 B.n338 B.n123 585
R250 B.n340 B.n339 585
R251 B.n341 B.n122 585
R252 B.n343 B.n342 585
R253 B.n344 B.n121 585
R254 B.n346 B.n345 585
R255 B.n347 B.n120 585
R256 B.n349 B.n348 585
R257 B.n350 B.n119 585
R258 B.n352 B.n351 585
R259 B.n353 B.n118 585
R260 B.n355 B.n354 585
R261 B.n356 B.n117 585
R262 B.n358 B.n357 585
R263 B.n359 B.n116 585
R264 B.n361 B.n360 585
R265 B.n362 B.n115 585
R266 B.n364 B.n363 585
R267 B.n365 B.n114 585
R268 B.n367 B.n366 585
R269 B.n368 B.n113 585
R270 B.n370 B.n369 585
R271 B.n371 B.n112 585
R272 B.n373 B.n372 585
R273 B.n374 B.n111 585
R274 B.n376 B.n375 585
R275 B.n377 B.n110 585
R276 B.n379 B.n378 585
R277 B.n380 B.n109 585
R278 B.n382 B.n381 585
R279 B.n383 B.n108 585
R280 B.n385 B.n384 585
R281 B.n386 B.n107 585
R282 B.n388 B.n387 585
R283 B.n389 B.n106 585
R284 B.n391 B.n390 585
R285 B.n392 B.n105 585
R286 B.n394 B.n393 585
R287 B.n217 B.n216 585
R288 B.n215 B.n168 585
R289 B.n214 B.n213 585
R290 B.n212 B.n169 585
R291 B.n211 B.n210 585
R292 B.n209 B.n170 585
R293 B.n208 B.n207 585
R294 B.n206 B.n171 585
R295 B.n205 B.n204 585
R296 B.n203 B.n172 585
R297 B.n202 B.n201 585
R298 B.n200 B.n173 585
R299 B.n199 B.n198 585
R300 B.n197 B.n174 585
R301 B.n196 B.n195 585
R302 B.n194 B.n175 585
R303 B.n193 B.n192 585
R304 B.n191 B.n176 585
R305 B.n190 B.n189 585
R306 B.n188 B.n177 585
R307 B.n187 B.n186 585
R308 B.n185 B.n178 585
R309 B.n184 B.n183 585
R310 B.n182 B.n179 585
R311 B.n181 B.n180 585
R312 B.n2 B.n0 585
R313 B.n689 B.n1 585
R314 B.n688 B.n687 585
R315 B.n686 B.n3 585
R316 B.n685 B.n684 585
R317 B.n683 B.n4 585
R318 B.n682 B.n681 585
R319 B.n680 B.n5 585
R320 B.n679 B.n678 585
R321 B.n677 B.n6 585
R322 B.n676 B.n675 585
R323 B.n674 B.n7 585
R324 B.n673 B.n672 585
R325 B.n671 B.n8 585
R326 B.n670 B.n669 585
R327 B.n668 B.n9 585
R328 B.n667 B.n666 585
R329 B.n665 B.n10 585
R330 B.n664 B.n663 585
R331 B.n662 B.n11 585
R332 B.n661 B.n660 585
R333 B.n659 B.n12 585
R334 B.n658 B.n657 585
R335 B.n656 B.n13 585
R336 B.n655 B.n654 585
R337 B.n653 B.n14 585
R338 B.n652 B.n651 585
R339 B.n691 B.n690 585
R340 B.n132 B.t2 507.781
R341 B.n50 B.t7 507.781
R342 B.n138 B.t5 507.781
R343 B.n42 B.t10 507.781
R344 B.n216 B.n167 468.476
R345 B.n652 B.n15 468.476
R346 B.n395 B.n394 468.476
R347 B.n474 B.n473 468.476
R348 B.n133 B.t1 449.211
R349 B.n51 B.t8 449.211
R350 B.n139 B.t4 449.211
R351 B.n43 B.t11 449.211
R352 B.n132 B.t0 352.332
R353 B.n138 B.t3 352.332
R354 B.n42 B.t9 352.332
R355 B.n50 B.t6 352.332
R356 B.n216 B.n215 163.367
R357 B.n215 B.n214 163.367
R358 B.n214 B.n169 163.367
R359 B.n210 B.n169 163.367
R360 B.n210 B.n209 163.367
R361 B.n209 B.n208 163.367
R362 B.n208 B.n171 163.367
R363 B.n204 B.n171 163.367
R364 B.n204 B.n203 163.367
R365 B.n203 B.n202 163.367
R366 B.n202 B.n173 163.367
R367 B.n198 B.n173 163.367
R368 B.n198 B.n197 163.367
R369 B.n197 B.n196 163.367
R370 B.n196 B.n175 163.367
R371 B.n192 B.n175 163.367
R372 B.n192 B.n191 163.367
R373 B.n191 B.n190 163.367
R374 B.n190 B.n177 163.367
R375 B.n186 B.n177 163.367
R376 B.n186 B.n185 163.367
R377 B.n185 B.n184 163.367
R378 B.n184 B.n179 163.367
R379 B.n180 B.n179 163.367
R380 B.n180 B.n2 163.367
R381 B.n690 B.n2 163.367
R382 B.n690 B.n689 163.367
R383 B.n689 B.n688 163.367
R384 B.n688 B.n3 163.367
R385 B.n684 B.n3 163.367
R386 B.n684 B.n683 163.367
R387 B.n683 B.n682 163.367
R388 B.n682 B.n5 163.367
R389 B.n678 B.n5 163.367
R390 B.n678 B.n677 163.367
R391 B.n677 B.n676 163.367
R392 B.n676 B.n7 163.367
R393 B.n672 B.n7 163.367
R394 B.n672 B.n671 163.367
R395 B.n671 B.n670 163.367
R396 B.n670 B.n9 163.367
R397 B.n666 B.n9 163.367
R398 B.n666 B.n665 163.367
R399 B.n665 B.n664 163.367
R400 B.n664 B.n11 163.367
R401 B.n660 B.n11 163.367
R402 B.n660 B.n659 163.367
R403 B.n659 B.n658 163.367
R404 B.n658 B.n13 163.367
R405 B.n654 B.n13 163.367
R406 B.n654 B.n653 163.367
R407 B.n653 B.n652 163.367
R408 B.n220 B.n167 163.367
R409 B.n221 B.n220 163.367
R410 B.n222 B.n221 163.367
R411 B.n222 B.n165 163.367
R412 B.n226 B.n165 163.367
R413 B.n227 B.n226 163.367
R414 B.n228 B.n227 163.367
R415 B.n228 B.n163 163.367
R416 B.n232 B.n163 163.367
R417 B.n233 B.n232 163.367
R418 B.n234 B.n233 163.367
R419 B.n234 B.n161 163.367
R420 B.n238 B.n161 163.367
R421 B.n239 B.n238 163.367
R422 B.n240 B.n239 163.367
R423 B.n240 B.n159 163.367
R424 B.n244 B.n159 163.367
R425 B.n245 B.n244 163.367
R426 B.n246 B.n245 163.367
R427 B.n246 B.n157 163.367
R428 B.n250 B.n157 163.367
R429 B.n251 B.n250 163.367
R430 B.n252 B.n251 163.367
R431 B.n252 B.n155 163.367
R432 B.n256 B.n155 163.367
R433 B.n257 B.n256 163.367
R434 B.n258 B.n257 163.367
R435 B.n258 B.n153 163.367
R436 B.n262 B.n153 163.367
R437 B.n263 B.n262 163.367
R438 B.n264 B.n263 163.367
R439 B.n264 B.n151 163.367
R440 B.n268 B.n151 163.367
R441 B.n269 B.n268 163.367
R442 B.n270 B.n269 163.367
R443 B.n270 B.n149 163.367
R444 B.n274 B.n149 163.367
R445 B.n275 B.n274 163.367
R446 B.n276 B.n275 163.367
R447 B.n276 B.n147 163.367
R448 B.n280 B.n147 163.367
R449 B.n281 B.n280 163.367
R450 B.n282 B.n281 163.367
R451 B.n282 B.n145 163.367
R452 B.n286 B.n145 163.367
R453 B.n287 B.n286 163.367
R454 B.n288 B.n287 163.367
R455 B.n288 B.n143 163.367
R456 B.n292 B.n143 163.367
R457 B.n293 B.n292 163.367
R458 B.n294 B.n293 163.367
R459 B.n294 B.n141 163.367
R460 B.n298 B.n141 163.367
R461 B.n299 B.n298 163.367
R462 B.n299 B.n137 163.367
R463 B.n303 B.n137 163.367
R464 B.n304 B.n303 163.367
R465 B.n305 B.n304 163.367
R466 B.n305 B.n135 163.367
R467 B.n309 B.n135 163.367
R468 B.n310 B.n309 163.367
R469 B.n311 B.n310 163.367
R470 B.n311 B.n131 163.367
R471 B.n316 B.n131 163.367
R472 B.n317 B.n316 163.367
R473 B.n318 B.n317 163.367
R474 B.n318 B.n129 163.367
R475 B.n322 B.n129 163.367
R476 B.n323 B.n322 163.367
R477 B.n324 B.n323 163.367
R478 B.n324 B.n127 163.367
R479 B.n328 B.n127 163.367
R480 B.n329 B.n328 163.367
R481 B.n330 B.n329 163.367
R482 B.n330 B.n125 163.367
R483 B.n334 B.n125 163.367
R484 B.n335 B.n334 163.367
R485 B.n336 B.n335 163.367
R486 B.n336 B.n123 163.367
R487 B.n340 B.n123 163.367
R488 B.n341 B.n340 163.367
R489 B.n342 B.n341 163.367
R490 B.n342 B.n121 163.367
R491 B.n346 B.n121 163.367
R492 B.n347 B.n346 163.367
R493 B.n348 B.n347 163.367
R494 B.n348 B.n119 163.367
R495 B.n352 B.n119 163.367
R496 B.n353 B.n352 163.367
R497 B.n354 B.n353 163.367
R498 B.n354 B.n117 163.367
R499 B.n358 B.n117 163.367
R500 B.n359 B.n358 163.367
R501 B.n360 B.n359 163.367
R502 B.n360 B.n115 163.367
R503 B.n364 B.n115 163.367
R504 B.n365 B.n364 163.367
R505 B.n366 B.n365 163.367
R506 B.n366 B.n113 163.367
R507 B.n370 B.n113 163.367
R508 B.n371 B.n370 163.367
R509 B.n372 B.n371 163.367
R510 B.n372 B.n111 163.367
R511 B.n376 B.n111 163.367
R512 B.n377 B.n376 163.367
R513 B.n378 B.n377 163.367
R514 B.n378 B.n109 163.367
R515 B.n382 B.n109 163.367
R516 B.n383 B.n382 163.367
R517 B.n384 B.n383 163.367
R518 B.n384 B.n107 163.367
R519 B.n388 B.n107 163.367
R520 B.n389 B.n388 163.367
R521 B.n390 B.n389 163.367
R522 B.n390 B.n105 163.367
R523 B.n394 B.n105 163.367
R524 B.n396 B.n395 163.367
R525 B.n396 B.n103 163.367
R526 B.n400 B.n103 163.367
R527 B.n401 B.n400 163.367
R528 B.n402 B.n401 163.367
R529 B.n402 B.n101 163.367
R530 B.n406 B.n101 163.367
R531 B.n407 B.n406 163.367
R532 B.n408 B.n407 163.367
R533 B.n408 B.n99 163.367
R534 B.n412 B.n99 163.367
R535 B.n413 B.n412 163.367
R536 B.n414 B.n413 163.367
R537 B.n414 B.n97 163.367
R538 B.n418 B.n97 163.367
R539 B.n419 B.n418 163.367
R540 B.n420 B.n419 163.367
R541 B.n420 B.n95 163.367
R542 B.n424 B.n95 163.367
R543 B.n425 B.n424 163.367
R544 B.n426 B.n425 163.367
R545 B.n426 B.n93 163.367
R546 B.n430 B.n93 163.367
R547 B.n431 B.n430 163.367
R548 B.n432 B.n431 163.367
R549 B.n432 B.n91 163.367
R550 B.n436 B.n91 163.367
R551 B.n437 B.n436 163.367
R552 B.n438 B.n437 163.367
R553 B.n438 B.n89 163.367
R554 B.n442 B.n89 163.367
R555 B.n443 B.n442 163.367
R556 B.n444 B.n443 163.367
R557 B.n444 B.n87 163.367
R558 B.n448 B.n87 163.367
R559 B.n449 B.n448 163.367
R560 B.n450 B.n449 163.367
R561 B.n450 B.n85 163.367
R562 B.n454 B.n85 163.367
R563 B.n455 B.n454 163.367
R564 B.n456 B.n455 163.367
R565 B.n456 B.n83 163.367
R566 B.n460 B.n83 163.367
R567 B.n461 B.n460 163.367
R568 B.n462 B.n461 163.367
R569 B.n462 B.n81 163.367
R570 B.n466 B.n81 163.367
R571 B.n467 B.n466 163.367
R572 B.n468 B.n467 163.367
R573 B.n468 B.n79 163.367
R574 B.n472 B.n79 163.367
R575 B.n473 B.n472 163.367
R576 B.n648 B.n15 163.367
R577 B.n648 B.n647 163.367
R578 B.n647 B.n646 163.367
R579 B.n646 B.n17 163.367
R580 B.n642 B.n17 163.367
R581 B.n642 B.n641 163.367
R582 B.n641 B.n640 163.367
R583 B.n640 B.n19 163.367
R584 B.n636 B.n19 163.367
R585 B.n636 B.n635 163.367
R586 B.n635 B.n634 163.367
R587 B.n634 B.n21 163.367
R588 B.n630 B.n21 163.367
R589 B.n630 B.n629 163.367
R590 B.n629 B.n628 163.367
R591 B.n628 B.n23 163.367
R592 B.n624 B.n23 163.367
R593 B.n624 B.n623 163.367
R594 B.n623 B.n622 163.367
R595 B.n622 B.n25 163.367
R596 B.n618 B.n25 163.367
R597 B.n618 B.n617 163.367
R598 B.n617 B.n616 163.367
R599 B.n616 B.n27 163.367
R600 B.n612 B.n27 163.367
R601 B.n612 B.n611 163.367
R602 B.n611 B.n610 163.367
R603 B.n610 B.n29 163.367
R604 B.n606 B.n29 163.367
R605 B.n606 B.n605 163.367
R606 B.n605 B.n604 163.367
R607 B.n604 B.n31 163.367
R608 B.n600 B.n31 163.367
R609 B.n600 B.n599 163.367
R610 B.n599 B.n598 163.367
R611 B.n598 B.n33 163.367
R612 B.n594 B.n33 163.367
R613 B.n594 B.n593 163.367
R614 B.n593 B.n592 163.367
R615 B.n592 B.n35 163.367
R616 B.n588 B.n35 163.367
R617 B.n588 B.n587 163.367
R618 B.n587 B.n586 163.367
R619 B.n586 B.n37 163.367
R620 B.n582 B.n37 163.367
R621 B.n582 B.n581 163.367
R622 B.n581 B.n580 163.367
R623 B.n580 B.n39 163.367
R624 B.n576 B.n39 163.367
R625 B.n576 B.n575 163.367
R626 B.n575 B.n574 163.367
R627 B.n574 B.n41 163.367
R628 B.n570 B.n41 163.367
R629 B.n570 B.n569 163.367
R630 B.n569 B.n45 163.367
R631 B.n565 B.n45 163.367
R632 B.n565 B.n564 163.367
R633 B.n564 B.n563 163.367
R634 B.n563 B.n47 163.367
R635 B.n559 B.n47 163.367
R636 B.n559 B.n558 163.367
R637 B.n558 B.n557 163.367
R638 B.n557 B.n49 163.367
R639 B.n552 B.n49 163.367
R640 B.n552 B.n551 163.367
R641 B.n551 B.n550 163.367
R642 B.n550 B.n53 163.367
R643 B.n546 B.n53 163.367
R644 B.n546 B.n545 163.367
R645 B.n545 B.n544 163.367
R646 B.n544 B.n55 163.367
R647 B.n540 B.n55 163.367
R648 B.n540 B.n539 163.367
R649 B.n539 B.n538 163.367
R650 B.n538 B.n57 163.367
R651 B.n534 B.n57 163.367
R652 B.n534 B.n533 163.367
R653 B.n533 B.n532 163.367
R654 B.n532 B.n59 163.367
R655 B.n528 B.n59 163.367
R656 B.n528 B.n527 163.367
R657 B.n527 B.n526 163.367
R658 B.n526 B.n61 163.367
R659 B.n522 B.n61 163.367
R660 B.n522 B.n521 163.367
R661 B.n521 B.n520 163.367
R662 B.n520 B.n63 163.367
R663 B.n516 B.n63 163.367
R664 B.n516 B.n515 163.367
R665 B.n515 B.n514 163.367
R666 B.n514 B.n65 163.367
R667 B.n510 B.n65 163.367
R668 B.n510 B.n509 163.367
R669 B.n509 B.n508 163.367
R670 B.n508 B.n67 163.367
R671 B.n504 B.n67 163.367
R672 B.n504 B.n503 163.367
R673 B.n503 B.n502 163.367
R674 B.n502 B.n69 163.367
R675 B.n498 B.n69 163.367
R676 B.n498 B.n497 163.367
R677 B.n497 B.n496 163.367
R678 B.n496 B.n71 163.367
R679 B.n492 B.n71 163.367
R680 B.n492 B.n491 163.367
R681 B.n491 B.n490 163.367
R682 B.n490 B.n73 163.367
R683 B.n486 B.n73 163.367
R684 B.n486 B.n485 163.367
R685 B.n485 B.n484 163.367
R686 B.n484 B.n75 163.367
R687 B.n480 B.n75 163.367
R688 B.n480 B.n479 163.367
R689 B.n479 B.n478 163.367
R690 B.n478 B.n77 163.367
R691 B.n474 B.n77 163.367
R692 B.n313 B.n133 59.5399
R693 B.n140 B.n139 59.5399
R694 B.n44 B.n43 59.5399
R695 B.n555 B.n51 59.5399
R696 B.n133 B.n132 58.5702
R697 B.n139 B.n138 58.5702
R698 B.n43 B.n42 58.5702
R699 B.n51 B.n50 58.5702
R700 B.n651 B.n650 30.4395
R701 B.n475 B.n78 30.4395
R702 B.n393 B.n104 30.4395
R703 B.n218 B.n217 30.4395
R704 B B.n691 18.0485
R705 B.n650 B.n649 10.6151
R706 B.n649 B.n16 10.6151
R707 B.n645 B.n16 10.6151
R708 B.n645 B.n644 10.6151
R709 B.n644 B.n643 10.6151
R710 B.n643 B.n18 10.6151
R711 B.n639 B.n18 10.6151
R712 B.n639 B.n638 10.6151
R713 B.n638 B.n637 10.6151
R714 B.n637 B.n20 10.6151
R715 B.n633 B.n20 10.6151
R716 B.n633 B.n632 10.6151
R717 B.n632 B.n631 10.6151
R718 B.n631 B.n22 10.6151
R719 B.n627 B.n22 10.6151
R720 B.n627 B.n626 10.6151
R721 B.n626 B.n625 10.6151
R722 B.n625 B.n24 10.6151
R723 B.n621 B.n24 10.6151
R724 B.n621 B.n620 10.6151
R725 B.n620 B.n619 10.6151
R726 B.n619 B.n26 10.6151
R727 B.n615 B.n26 10.6151
R728 B.n615 B.n614 10.6151
R729 B.n614 B.n613 10.6151
R730 B.n613 B.n28 10.6151
R731 B.n609 B.n28 10.6151
R732 B.n609 B.n608 10.6151
R733 B.n608 B.n607 10.6151
R734 B.n607 B.n30 10.6151
R735 B.n603 B.n30 10.6151
R736 B.n603 B.n602 10.6151
R737 B.n602 B.n601 10.6151
R738 B.n601 B.n32 10.6151
R739 B.n597 B.n32 10.6151
R740 B.n597 B.n596 10.6151
R741 B.n596 B.n595 10.6151
R742 B.n595 B.n34 10.6151
R743 B.n591 B.n34 10.6151
R744 B.n591 B.n590 10.6151
R745 B.n590 B.n589 10.6151
R746 B.n589 B.n36 10.6151
R747 B.n585 B.n36 10.6151
R748 B.n585 B.n584 10.6151
R749 B.n584 B.n583 10.6151
R750 B.n583 B.n38 10.6151
R751 B.n579 B.n38 10.6151
R752 B.n579 B.n578 10.6151
R753 B.n578 B.n577 10.6151
R754 B.n577 B.n40 10.6151
R755 B.n573 B.n40 10.6151
R756 B.n573 B.n572 10.6151
R757 B.n572 B.n571 10.6151
R758 B.n568 B.n567 10.6151
R759 B.n567 B.n566 10.6151
R760 B.n566 B.n46 10.6151
R761 B.n562 B.n46 10.6151
R762 B.n562 B.n561 10.6151
R763 B.n561 B.n560 10.6151
R764 B.n560 B.n48 10.6151
R765 B.n556 B.n48 10.6151
R766 B.n554 B.n553 10.6151
R767 B.n553 B.n52 10.6151
R768 B.n549 B.n52 10.6151
R769 B.n549 B.n548 10.6151
R770 B.n548 B.n547 10.6151
R771 B.n547 B.n54 10.6151
R772 B.n543 B.n54 10.6151
R773 B.n543 B.n542 10.6151
R774 B.n542 B.n541 10.6151
R775 B.n541 B.n56 10.6151
R776 B.n537 B.n56 10.6151
R777 B.n537 B.n536 10.6151
R778 B.n536 B.n535 10.6151
R779 B.n535 B.n58 10.6151
R780 B.n531 B.n58 10.6151
R781 B.n531 B.n530 10.6151
R782 B.n530 B.n529 10.6151
R783 B.n529 B.n60 10.6151
R784 B.n525 B.n60 10.6151
R785 B.n525 B.n524 10.6151
R786 B.n524 B.n523 10.6151
R787 B.n523 B.n62 10.6151
R788 B.n519 B.n62 10.6151
R789 B.n519 B.n518 10.6151
R790 B.n518 B.n517 10.6151
R791 B.n517 B.n64 10.6151
R792 B.n513 B.n64 10.6151
R793 B.n513 B.n512 10.6151
R794 B.n512 B.n511 10.6151
R795 B.n511 B.n66 10.6151
R796 B.n507 B.n66 10.6151
R797 B.n507 B.n506 10.6151
R798 B.n506 B.n505 10.6151
R799 B.n505 B.n68 10.6151
R800 B.n501 B.n68 10.6151
R801 B.n501 B.n500 10.6151
R802 B.n500 B.n499 10.6151
R803 B.n499 B.n70 10.6151
R804 B.n495 B.n70 10.6151
R805 B.n495 B.n494 10.6151
R806 B.n494 B.n493 10.6151
R807 B.n493 B.n72 10.6151
R808 B.n489 B.n72 10.6151
R809 B.n489 B.n488 10.6151
R810 B.n488 B.n487 10.6151
R811 B.n487 B.n74 10.6151
R812 B.n483 B.n74 10.6151
R813 B.n483 B.n482 10.6151
R814 B.n482 B.n481 10.6151
R815 B.n481 B.n76 10.6151
R816 B.n477 B.n76 10.6151
R817 B.n477 B.n476 10.6151
R818 B.n476 B.n475 10.6151
R819 B.n397 B.n104 10.6151
R820 B.n398 B.n397 10.6151
R821 B.n399 B.n398 10.6151
R822 B.n399 B.n102 10.6151
R823 B.n403 B.n102 10.6151
R824 B.n404 B.n403 10.6151
R825 B.n405 B.n404 10.6151
R826 B.n405 B.n100 10.6151
R827 B.n409 B.n100 10.6151
R828 B.n410 B.n409 10.6151
R829 B.n411 B.n410 10.6151
R830 B.n411 B.n98 10.6151
R831 B.n415 B.n98 10.6151
R832 B.n416 B.n415 10.6151
R833 B.n417 B.n416 10.6151
R834 B.n417 B.n96 10.6151
R835 B.n421 B.n96 10.6151
R836 B.n422 B.n421 10.6151
R837 B.n423 B.n422 10.6151
R838 B.n423 B.n94 10.6151
R839 B.n427 B.n94 10.6151
R840 B.n428 B.n427 10.6151
R841 B.n429 B.n428 10.6151
R842 B.n429 B.n92 10.6151
R843 B.n433 B.n92 10.6151
R844 B.n434 B.n433 10.6151
R845 B.n435 B.n434 10.6151
R846 B.n435 B.n90 10.6151
R847 B.n439 B.n90 10.6151
R848 B.n440 B.n439 10.6151
R849 B.n441 B.n440 10.6151
R850 B.n441 B.n88 10.6151
R851 B.n445 B.n88 10.6151
R852 B.n446 B.n445 10.6151
R853 B.n447 B.n446 10.6151
R854 B.n447 B.n86 10.6151
R855 B.n451 B.n86 10.6151
R856 B.n452 B.n451 10.6151
R857 B.n453 B.n452 10.6151
R858 B.n453 B.n84 10.6151
R859 B.n457 B.n84 10.6151
R860 B.n458 B.n457 10.6151
R861 B.n459 B.n458 10.6151
R862 B.n459 B.n82 10.6151
R863 B.n463 B.n82 10.6151
R864 B.n464 B.n463 10.6151
R865 B.n465 B.n464 10.6151
R866 B.n465 B.n80 10.6151
R867 B.n469 B.n80 10.6151
R868 B.n470 B.n469 10.6151
R869 B.n471 B.n470 10.6151
R870 B.n471 B.n78 10.6151
R871 B.n219 B.n218 10.6151
R872 B.n219 B.n166 10.6151
R873 B.n223 B.n166 10.6151
R874 B.n224 B.n223 10.6151
R875 B.n225 B.n224 10.6151
R876 B.n225 B.n164 10.6151
R877 B.n229 B.n164 10.6151
R878 B.n230 B.n229 10.6151
R879 B.n231 B.n230 10.6151
R880 B.n231 B.n162 10.6151
R881 B.n235 B.n162 10.6151
R882 B.n236 B.n235 10.6151
R883 B.n237 B.n236 10.6151
R884 B.n237 B.n160 10.6151
R885 B.n241 B.n160 10.6151
R886 B.n242 B.n241 10.6151
R887 B.n243 B.n242 10.6151
R888 B.n243 B.n158 10.6151
R889 B.n247 B.n158 10.6151
R890 B.n248 B.n247 10.6151
R891 B.n249 B.n248 10.6151
R892 B.n249 B.n156 10.6151
R893 B.n253 B.n156 10.6151
R894 B.n254 B.n253 10.6151
R895 B.n255 B.n254 10.6151
R896 B.n255 B.n154 10.6151
R897 B.n259 B.n154 10.6151
R898 B.n260 B.n259 10.6151
R899 B.n261 B.n260 10.6151
R900 B.n261 B.n152 10.6151
R901 B.n265 B.n152 10.6151
R902 B.n266 B.n265 10.6151
R903 B.n267 B.n266 10.6151
R904 B.n267 B.n150 10.6151
R905 B.n271 B.n150 10.6151
R906 B.n272 B.n271 10.6151
R907 B.n273 B.n272 10.6151
R908 B.n273 B.n148 10.6151
R909 B.n277 B.n148 10.6151
R910 B.n278 B.n277 10.6151
R911 B.n279 B.n278 10.6151
R912 B.n279 B.n146 10.6151
R913 B.n283 B.n146 10.6151
R914 B.n284 B.n283 10.6151
R915 B.n285 B.n284 10.6151
R916 B.n285 B.n144 10.6151
R917 B.n289 B.n144 10.6151
R918 B.n290 B.n289 10.6151
R919 B.n291 B.n290 10.6151
R920 B.n291 B.n142 10.6151
R921 B.n295 B.n142 10.6151
R922 B.n296 B.n295 10.6151
R923 B.n297 B.n296 10.6151
R924 B.n301 B.n300 10.6151
R925 B.n302 B.n301 10.6151
R926 B.n302 B.n136 10.6151
R927 B.n306 B.n136 10.6151
R928 B.n307 B.n306 10.6151
R929 B.n308 B.n307 10.6151
R930 B.n308 B.n134 10.6151
R931 B.n312 B.n134 10.6151
R932 B.n315 B.n314 10.6151
R933 B.n315 B.n130 10.6151
R934 B.n319 B.n130 10.6151
R935 B.n320 B.n319 10.6151
R936 B.n321 B.n320 10.6151
R937 B.n321 B.n128 10.6151
R938 B.n325 B.n128 10.6151
R939 B.n326 B.n325 10.6151
R940 B.n327 B.n326 10.6151
R941 B.n327 B.n126 10.6151
R942 B.n331 B.n126 10.6151
R943 B.n332 B.n331 10.6151
R944 B.n333 B.n332 10.6151
R945 B.n333 B.n124 10.6151
R946 B.n337 B.n124 10.6151
R947 B.n338 B.n337 10.6151
R948 B.n339 B.n338 10.6151
R949 B.n339 B.n122 10.6151
R950 B.n343 B.n122 10.6151
R951 B.n344 B.n343 10.6151
R952 B.n345 B.n344 10.6151
R953 B.n345 B.n120 10.6151
R954 B.n349 B.n120 10.6151
R955 B.n350 B.n349 10.6151
R956 B.n351 B.n350 10.6151
R957 B.n351 B.n118 10.6151
R958 B.n355 B.n118 10.6151
R959 B.n356 B.n355 10.6151
R960 B.n357 B.n356 10.6151
R961 B.n357 B.n116 10.6151
R962 B.n361 B.n116 10.6151
R963 B.n362 B.n361 10.6151
R964 B.n363 B.n362 10.6151
R965 B.n363 B.n114 10.6151
R966 B.n367 B.n114 10.6151
R967 B.n368 B.n367 10.6151
R968 B.n369 B.n368 10.6151
R969 B.n369 B.n112 10.6151
R970 B.n373 B.n112 10.6151
R971 B.n374 B.n373 10.6151
R972 B.n375 B.n374 10.6151
R973 B.n375 B.n110 10.6151
R974 B.n379 B.n110 10.6151
R975 B.n380 B.n379 10.6151
R976 B.n381 B.n380 10.6151
R977 B.n381 B.n108 10.6151
R978 B.n385 B.n108 10.6151
R979 B.n386 B.n385 10.6151
R980 B.n387 B.n386 10.6151
R981 B.n387 B.n106 10.6151
R982 B.n391 B.n106 10.6151
R983 B.n392 B.n391 10.6151
R984 B.n393 B.n392 10.6151
R985 B.n217 B.n168 10.6151
R986 B.n213 B.n168 10.6151
R987 B.n213 B.n212 10.6151
R988 B.n212 B.n211 10.6151
R989 B.n211 B.n170 10.6151
R990 B.n207 B.n170 10.6151
R991 B.n207 B.n206 10.6151
R992 B.n206 B.n205 10.6151
R993 B.n205 B.n172 10.6151
R994 B.n201 B.n172 10.6151
R995 B.n201 B.n200 10.6151
R996 B.n200 B.n199 10.6151
R997 B.n199 B.n174 10.6151
R998 B.n195 B.n174 10.6151
R999 B.n195 B.n194 10.6151
R1000 B.n194 B.n193 10.6151
R1001 B.n193 B.n176 10.6151
R1002 B.n189 B.n176 10.6151
R1003 B.n189 B.n188 10.6151
R1004 B.n188 B.n187 10.6151
R1005 B.n187 B.n178 10.6151
R1006 B.n183 B.n178 10.6151
R1007 B.n183 B.n182 10.6151
R1008 B.n182 B.n181 10.6151
R1009 B.n181 B.n0 10.6151
R1010 B.n687 B.n1 10.6151
R1011 B.n687 B.n686 10.6151
R1012 B.n686 B.n685 10.6151
R1013 B.n685 B.n4 10.6151
R1014 B.n681 B.n4 10.6151
R1015 B.n681 B.n680 10.6151
R1016 B.n680 B.n679 10.6151
R1017 B.n679 B.n6 10.6151
R1018 B.n675 B.n6 10.6151
R1019 B.n675 B.n674 10.6151
R1020 B.n674 B.n673 10.6151
R1021 B.n673 B.n8 10.6151
R1022 B.n669 B.n8 10.6151
R1023 B.n669 B.n668 10.6151
R1024 B.n668 B.n667 10.6151
R1025 B.n667 B.n10 10.6151
R1026 B.n663 B.n10 10.6151
R1027 B.n663 B.n662 10.6151
R1028 B.n662 B.n661 10.6151
R1029 B.n661 B.n12 10.6151
R1030 B.n657 B.n12 10.6151
R1031 B.n657 B.n656 10.6151
R1032 B.n656 B.n655 10.6151
R1033 B.n655 B.n14 10.6151
R1034 B.n651 B.n14 10.6151
R1035 B.n568 B.n44 6.5566
R1036 B.n556 B.n555 6.5566
R1037 B.n300 B.n140 6.5566
R1038 B.n313 B.n312 6.5566
R1039 B.n571 B.n44 4.05904
R1040 B.n555 B.n554 4.05904
R1041 B.n297 B.n140 4.05904
R1042 B.n314 B.n313 4.05904
R1043 B.n691 B.n0 2.81026
R1044 B.n691 B.n1 2.81026
R1045 VN VN.t0 233.244
R1046 VN VN.t1 185.679
R1047 VTAIL.n354 VTAIL.n270 756.745
R1048 VTAIL.n84 VTAIL.n0 756.745
R1049 VTAIL.n264 VTAIL.n180 756.745
R1050 VTAIL.n174 VTAIL.n90 756.745
R1051 VTAIL.n298 VTAIL.n297 585
R1052 VTAIL.n303 VTAIL.n302 585
R1053 VTAIL.n305 VTAIL.n304 585
R1054 VTAIL.n294 VTAIL.n293 585
R1055 VTAIL.n311 VTAIL.n310 585
R1056 VTAIL.n313 VTAIL.n312 585
R1057 VTAIL.n290 VTAIL.n289 585
R1058 VTAIL.n319 VTAIL.n318 585
R1059 VTAIL.n321 VTAIL.n320 585
R1060 VTAIL.n286 VTAIL.n285 585
R1061 VTAIL.n327 VTAIL.n326 585
R1062 VTAIL.n329 VTAIL.n328 585
R1063 VTAIL.n282 VTAIL.n281 585
R1064 VTAIL.n335 VTAIL.n334 585
R1065 VTAIL.n337 VTAIL.n336 585
R1066 VTAIL.n278 VTAIL.n277 585
R1067 VTAIL.n344 VTAIL.n343 585
R1068 VTAIL.n345 VTAIL.n276 585
R1069 VTAIL.n347 VTAIL.n346 585
R1070 VTAIL.n274 VTAIL.n273 585
R1071 VTAIL.n353 VTAIL.n352 585
R1072 VTAIL.n355 VTAIL.n354 585
R1073 VTAIL.n28 VTAIL.n27 585
R1074 VTAIL.n33 VTAIL.n32 585
R1075 VTAIL.n35 VTAIL.n34 585
R1076 VTAIL.n24 VTAIL.n23 585
R1077 VTAIL.n41 VTAIL.n40 585
R1078 VTAIL.n43 VTAIL.n42 585
R1079 VTAIL.n20 VTAIL.n19 585
R1080 VTAIL.n49 VTAIL.n48 585
R1081 VTAIL.n51 VTAIL.n50 585
R1082 VTAIL.n16 VTAIL.n15 585
R1083 VTAIL.n57 VTAIL.n56 585
R1084 VTAIL.n59 VTAIL.n58 585
R1085 VTAIL.n12 VTAIL.n11 585
R1086 VTAIL.n65 VTAIL.n64 585
R1087 VTAIL.n67 VTAIL.n66 585
R1088 VTAIL.n8 VTAIL.n7 585
R1089 VTAIL.n74 VTAIL.n73 585
R1090 VTAIL.n75 VTAIL.n6 585
R1091 VTAIL.n77 VTAIL.n76 585
R1092 VTAIL.n4 VTAIL.n3 585
R1093 VTAIL.n83 VTAIL.n82 585
R1094 VTAIL.n85 VTAIL.n84 585
R1095 VTAIL.n265 VTAIL.n264 585
R1096 VTAIL.n263 VTAIL.n262 585
R1097 VTAIL.n184 VTAIL.n183 585
R1098 VTAIL.n257 VTAIL.n256 585
R1099 VTAIL.n255 VTAIL.n186 585
R1100 VTAIL.n254 VTAIL.n253 585
R1101 VTAIL.n189 VTAIL.n187 585
R1102 VTAIL.n248 VTAIL.n247 585
R1103 VTAIL.n246 VTAIL.n245 585
R1104 VTAIL.n193 VTAIL.n192 585
R1105 VTAIL.n240 VTAIL.n239 585
R1106 VTAIL.n238 VTAIL.n237 585
R1107 VTAIL.n197 VTAIL.n196 585
R1108 VTAIL.n232 VTAIL.n231 585
R1109 VTAIL.n230 VTAIL.n229 585
R1110 VTAIL.n201 VTAIL.n200 585
R1111 VTAIL.n224 VTAIL.n223 585
R1112 VTAIL.n222 VTAIL.n221 585
R1113 VTAIL.n205 VTAIL.n204 585
R1114 VTAIL.n216 VTAIL.n215 585
R1115 VTAIL.n214 VTAIL.n213 585
R1116 VTAIL.n209 VTAIL.n208 585
R1117 VTAIL.n175 VTAIL.n174 585
R1118 VTAIL.n173 VTAIL.n172 585
R1119 VTAIL.n94 VTAIL.n93 585
R1120 VTAIL.n167 VTAIL.n166 585
R1121 VTAIL.n165 VTAIL.n96 585
R1122 VTAIL.n164 VTAIL.n163 585
R1123 VTAIL.n99 VTAIL.n97 585
R1124 VTAIL.n158 VTAIL.n157 585
R1125 VTAIL.n156 VTAIL.n155 585
R1126 VTAIL.n103 VTAIL.n102 585
R1127 VTAIL.n150 VTAIL.n149 585
R1128 VTAIL.n148 VTAIL.n147 585
R1129 VTAIL.n107 VTAIL.n106 585
R1130 VTAIL.n142 VTAIL.n141 585
R1131 VTAIL.n140 VTAIL.n139 585
R1132 VTAIL.n111 VTAIL.n110 585
R1133 VTAIL.n134 VTAIL.n133 585
R1134 VTAIL.n132 VTAIL.n131 585
R1135 VTAIL.n115 VTAIL.n114 585
R1136 VTAIL.n126 VTAIL.n125 585
R1137 VTAIL.n124 VTAIL.n123 585
R1138 VTAIL.n119 VTAIL.n118 585
R1139 VTAIL.n299 VTAIL.t2 327.466
R1140 VTAIL.n29 VTAIL.t0 327.466
R1141 VTAIL.n210 VTAIL.t1 327.466
R1142 VTAIL.n120 VTAIL.t3 327.466
R1143 VTAIL.n303 VTAIL.n297 171.744
R1144 VTAIL.n304 VTAIL.n303 171.744
R1145 VTAIL.n304 VTAIL.n293 171.744
R1146 VTAIL.n311 VTAIL.n293 171.744
R1147 VTAIL.n312 VTAIL.n311 171.744
R1148 VTAIL.n312 VTAIL.n289 171.744
R1149 VTAIL.n319 VTAIL.n289 171.744
R1150 VTAIL.n320 VTAIL.n319 171.744
R1151 VTAIL.n320 VTAIL.n285 171.744
R1152 VTAIL.n327 VTAIL.n285 171.744
R1153 VTAIL.n328 VTAIL.n327 171.744
R1154 VTAIL.n328 VTAIL.n281 171.744
R1155 VTAIL.n335 VTAIL.n281 171.744
R1156 VTAIL.n336 VTAIL.n335 171.744
R1157 VTAIL.n336 VTAIL.n277 171.744
R1158 VTAIL.n344 VTAIL.n277 171.744
R1159 VTAIL.n345 VTAIL.n344 171.744
R1160 VTAIL.n346 VTAIL.n345 171.744
R1161 VTAIL.n346 VTAIL.n273 171.744
R1162 VTAIL.n353 VTAIL.n273 171.744
R1163 VTAIL.n354 VTAIL.n353 171.744
R1164 VTAIL.n33 VTAIL.n27 171.744
R1165 VTAIL.n34 VTAIL.n33 171.744
R1166 VTAIL.n34 VTAIL.n23 171.744
R1167 VTAIL.n41 VTAIL.n23 171.744
R1168 VTAIL.n42 VTAIL.n41 171.744
R1169 VTAIL.n42 VTAIL.n19 171.744
R1170 VTAIL.n49 VTAIL.n19 171.744
R1171 VTAIL.n50 VTAIL.n49 171.744
R1172 VTAIL.n50 VTAIL.n15 171.744
R1173 VTAIL.n57 VTAIL.n15 171.744
R1174 VTAIL.n58 VTAIL.n57 171.744
R1175 VTAIL.n58 VTAIL.n11 171.744
R1176 VTAIL.n65 VTAIL.n11 171.744
R1177 VTAIL.n66 VTAIL.n65 171.744
R1178 VTAIL.n66 VTAIL.n7 171.744
R1179 VTAIL.n74 VTAIL.n7 171.744
R1180 VTAIL.n75 VTAIL.n74 171.744
R1181 VTAIL.n76 VTAIL.n75 171.744
R1182 VTAIL.n76 VTAIL.n3 171.744
R1183 VTAIL.n83 VTAIL.n3 171.744
R1184 VTAIL.n84 VTAIL.n83 171.744
R1185 VTAIL.n264 VTAIL.n263 171.744
R1186 VTAIL.n263 VTAIL.n183 171.744
R1187 VTAIL.n256 VTAIL.n183 171.744
R1188 VTAIL.n256 VTAIL.n255 171.744
R1189 VTAIL.n255 VTAIL.n254 171.744
R1190 VTAIL.n254 VTAIL.n187 171.744
R1191 VTAIL.n247 VTAIL.n187 171.744
R1192 VTAIL.n247 VTAIL.n246 171.744
R1193 VTAIL.n246 VTAIL.n192 171.744
R1194 VTAIL.n239 VTAIL.n192 171.744
R1195 VTAIL.n239 VTAIL.n238 171.744
R1196 VTAIL.n238 VTAIL.n196 171.744
R1197 VTAIL.n231 VTAIL.n196 171.744
R1198 VTAIL.n231 VTAIL.n230 171.744
R1199 VTAIL.n230 VTAIL.n200 171.744
R1200 VTAIL.n223 VTAIL.n200 171.744
R1201 VTAIL.n223 VTAIL.n222 171.744
R1202 VTAIL.n222 VTAIL.n204 171.744
R1203 VTAIL.n215 VTAIL.n204 171.744
R1204 VTAIL.n215 VTAIL.n214 171.744
R1205 VTAIL.n214 VTAIL.n208 171.744
R1206 VTAIL.n174 VTAIL.n173 171.744
R1207 VTAIL.n173 VTAIL.n93 171.744
R1208 VTAIL.n166 VTAIL.n93 171.744
R1209 VTAIL.n166 VTAIL.n165 171.744
R1210 VTAIL.n165 VTAIL.n164 171.744
R1211 VTAIL.n164 VTAIL.n97 171.744
R1212 VTAIL.n157 VTAIL.n97 171.744
R1213 VTAIL.n157 VTAIL.n156 171.744
R1214 VTAIL.n156 VTAIL.n102 171.744
R1215 VTAIL.n149 VTAIL.n102 171.744
R1216 VTAIL.n149 VTAIL.n148 171.744
R1217 VTAIL.n148 VTAIL.n106 171.744
R1218 VTAIL.n141 VTAIL.n106 171.744
R1219 VTAIL.n141 VTAIL.n140 171.744
R1220 VTAIL.n140 VTAIL.n110 171.744
R1221 VTAIL.n133 VTAIL.n110 171.744
R1222 VTAIL.n133 VTAIL.n132 171.744
R1223 VTAIL.n132 VTAIL.n114 171.744
R1224 VTAIL.n125 VTAIL.n114 171.744
R1225 VTAIL.n125 VTAIL.n124 171.744
R1226 VTAIL.n124 VTAIL.n118 171.744
R1227 VTAIL.t2 VTAIL.n297 85.8723
R1228 VTAIL.t0 VTAIL.n27 85.8723
R1229 VTAIL.t1 VTAIL.n208 85.8723
R1230 VTAIL.t3 VTAIL.n118 85.8723
R1231 VTAIL.n359 VTAIL.n358 32.3793
R1232 VTAIL.n89 VTAIL.n88 32.3793
R1233 VTAIL.n269 VTAIL.n268 32.3793
R1234 VTAIL.n179 VTAIL.n178 32.3793
R1235 VTAIL.n179 VTAIL.n89 31.4445
R1236 VTAIL.n359 VTAIL.n269 28.841
R1237 VTAIL.n299 VTAIL.n298 16.3895
R1238 VTAIL.n29 VTAIL.n28 16.3895
R1239 VTAIL.n210 VTAIL.n209 16.3895
R1240 VTAIL.n120 VTAIL.n119 16.3895
R1241 VTAIL.n347 VTAIL.n276 13.1884
R1242 VTAIL.n77 VTAIL.n6 13.1884
R1243 VTAIL.n257 VTAIL.n186 13.1884
R1244 VTAIL.n167 VTAIL.n96 13.1884
R1245 VTAIL.n302 VTAIL.n301 12.8005
R1246 VTAIL.n343 VTAIL.n342 12.8005
R1247 VTAIL.n348 VTAIL.n274 12.8005
R1248 VTAIL.n32 VTAIL.n31 12.8005
R1249 VTAIL.n73 VTAIL.n72 12.8005
R1250 VTAIL.n78 VTAIL.n4 12.8005
R1251 VTAIL.n258 VTAIL.n184 12.8005
R1252 VTAIL.n253 VTAIL.n188 12.8005
R1253 VTAIL.n213 VTAIL.n212 12.8005
R1254 VTAIL.n168 VTAIL.n94 12.8005
R1255 VTAIL.n163 VTAIL.n98 12.8005
R1256 VTAIL.n123 VTAIL.n122 12.8005
R1257 VTAIL.n305 VTAIL.n296 12.0247
R1258 VTAIL.n341 VTAIL.n278 12.0247
R1259 VTAIL.n352 VTAIL.n351 12.0247
R1260 VTAIL.n35 VTAIL.n26 12.0247
R1261 VTAIL.n71 VTAIL.n8 12.0247
R1262 VTAIL.n82 VTAIL.n81 12.0247
R1263 VTAIL.n262 VTAIL.n261 12.0247
R1264 VTAIL.n252 VTAIL.n189 12.0247
R1265 VTAIL.n216 VTAIL.n207 12.0247
R1266 VTAIL.n172 VTAIL.n171 12.0247
R1267 VTAIL.n162 VTAIL.n99 12.0247
R1268 VTAIL.n126 VTAIL.n117 12.0247
R1269 VTAIL.n306 VTAIL.n294 11.249
R1270 VTAIL.n338 VTAIL.n337 11.249
R1271 VTAIL.n355 VTAIL.n272 11.249
R1272 VTAIL.n36 VTAIL.n24 11.249
R1273 VTAIL.n68 VTAIL.n67 11.249
R1274 VTAIL.n85 VTAIL.n2 11.249
R1275 VTAIL.n265 VTAIL.n182 11.249
R1276 VTAIL.n249 VTAIL.n248 11.249
R1277 VTAIL.n217 VTAIL.n205 11.249
R1278 VTAIL.n175 VTAIL.n92 11.249
R1279 VTAIL.n159 VTAIL.n158 11.249
R1280 VTAIL.n127 VTAIL.n115 11.249
R1281 VTAIL.n310 VTAIL.n309 10.4732
R1282 VTAIL.n334 VTAIL.n280 10.4732
R1283 VTAIL.n356 VTAIL.n270 10.4732
R1284 VTAIL.n40 VTAIL.n39 10.4732
R1285 VTAIL.n64 VTAIL.n10 10.4732
R1286 VTAIL.n86 VTAIL.n0 10.4732
R1287 VTAIL.n266 VTAIL.n180 10.4732
R1288 VTAIL.n245 VTAIL.n191 10.4732
R1289 VTAIL.n221 VTAIL.n220 10.4732
R1290 VTAIL.n176 VTAIL.n90 10.4732
R1291 VTAIL.n155 VTAIL.n101 10.4732
R1292 VTAIL.n131 VTAIL.n130 10.4732
R1293 VTAIL.n313 VTAIL.n292 9.69747
R1294 VTAIL.n333 VTAIL.n282 9.69747
R1295 VTAIL.n43 VTAIL.n22 9.69747
R1296 VTAIL.n63 VTAIL.n12 9.69747
R1297 VTAIL.n244 VTAIL.n193 9.69747
R1298 VTAIL.n224 VTAIL.n203 9.69747
R1299 VTAIL.n154 VTAIL.n103 9.69747
R1300 VTAIL.n134 VTAIL.n113 9.69747
R1301 VTAIL.n358 VTAIL.n357 9.45567
R1302 VTAIL.n88 VTAIL.n87 9.45567
R1303 VTAIL.n268 VTAIL.n267 9.45567
R1304 VTAIL.n178 VTAIL.n177 9.45567
R1305 VTAIL.n357 VTAIL.n356 9.3005
R1306 VTAIL.n272 VTAIL.n271 9.3005
R1307 VTAIL.n351 VTAIL.n350 9.3005
R1308 VTAIL.n349 VTAIL.n348 9.3005
R1309 VTAIL.n288 VTAIL.n287 9.3005
R1310 VTAIL.n317 VTAIL.n316 9.3005
R1311 VTAIL.n315 VTAIL.n314 9.3005
R1312 VTAIL.n292 VTAIL.n291 9.3005
R1313 VTAIL.n309 VTAIL.n308 9.3005
R1314 VTAIL.n307 VTAIL.n306 9.3005
R1315 VTAIL.n296 VTAIL.n295 9.3005
R1316 VTAIL.n301 VTAIL.n300 9.3005
R1317 VTAIL.n323 VTAIL.n322 9.3005
R1318 VTAIL.n325 VTAIL.n324 9.3005
R1319 VTAIL.n284 VTAIL.n283 9.3005
R1320 VTAIL.n331 VTAIL.n330 9.3005
R1321 VTAIL.n333 VTAIL.n332 9.3005
R1322 VTAIL.n280 VTAIL.n279 9.3005
R1323 VTAIL.n339 VTAIL.n338 9.3005
R1324 VTAIL.n341 VTAIL.n340 9.3005
R1325 VTAIL.n342 VTAIL.n275 9.3005
R1326 VTAIL.n87 VTAIL.n86 9.3005
R1327 VTAIL.n2 VTAIL.n1 9.3005
R1328 VTAIL.n81 VTAIL.n80 9.3005
R1329 VTAIL.n79 VTAIL.n78 9.3005
R1330 VTAIL.n18 VTAIL.n17 9.3005
R1331 VTAIL.n47 VTAIL.n46 9.3005
R1332 VTAIL.n45 VTAIL.n44 9.3005
R1333 VTAIL.n22 VTAIL.n21 9.3005
R1334 VTAIL.n39 VTAIL.n38 9.3005
R1335 VTAIL.n37 VTAIL.n36 9.3005
R1336 VTAIL.n26 VTAIL.n25 9.3005
R1337 VTAIL.n31 VTAIL.n30 9.3005
R1338 VTAIL.n53 VTAIL.n52 9.3005
R1339 VTAIL.n55 VTAIL.n54 9.3005
R1340 VTAIL.n14 VTAIL.n13 9.3005
R1341 VTAIL.n61 VTAIL.n60 9.3005
R1342 VTAIL.n63 VTAIL.n62 9.3005
R1343 VTAIL.n10 VTAIL.n9 9.3005
R1344 VTAIL.n69 VTAIL.n68 9.3005
R1345 VTAIL.n71 VTAIL.n70 9.3005
R1346 VTAIL.n72 VTAIL.n5 9.3005
R1347 VTAIL.n236 VTAIL.n235 9.3005
R1348 VTAIL.n195 VTAIL.n194 9.3005
R1349 VTAIL.n242 VTAIL.n241 9.3005
R1350 VTAIL.n244 VTAIL.n243 9.3005
R1351 VTAIL.n191 VTAIL.n190 9.3005
R1352 VTAIL.n250 VTAIL.n249 9.3005
R1353 VTAIL.n252 VTAIL.n251 9.3005
R1354 VTAIL.n188 VTAIL.n185 9.3005
R1355 VTAIL.n267 VTAIL.n266 9.3005
R1356 VTAIL.n182 VTAIL.n181 9.3005
R1357 VTAIL.n261 VTAIL.n260 9.3005
R1358 VTAIL.n259 VTAIL.n258 9.3005
R1359 VTAIL.n234 VTAIL.n233 9.3005
R1360 VTAIL.n199 VTAIL.n198 9.3005
R1361 VTAIL.n228 VTAIL.n227 9.3005
R1362 VTAIL.n226 VTAIL.n225 9.3005
R1363 VTAIL.n203 VTAIL.n202 9.3005
R1364 VTAIL.n220 VTAIL.n219 9.3005
R1365 VTAIL.n218 VTAIL.n217 9.3005
R1366 VTAIL.n207 VTAIL.n206 9.3005
R1367 VTAIL.n212 VTAIL.n211 9.3005
R1368 VTAIL.n146 VTAIL.n145 9.3005
R1369 VTAIL.n105 VTAIL.n104 9.3005
R1370 VTAIL.n152 VTAIL.n151 9.3005
R1371 VTAIL.n154 VTAIL.n153 9.3005
R1372 VTAIL.n101 VTAIL.n100 9.3005
R1373 VTAIL.n160 VTAIL.n159 9.3005
R1374 VTAIL.n162 VTAIL.n161 9.3005
R1375 VTAIL.n98 VTAIL.n95 9.3005
R1376 VTAIL.n177 VTAIL.n176 9.3005
R1377 VTAIL.n92 VTAIL.n91 9.3005
R1378 VTAIL.n171 VTAIL.n170 9.3005
R1379 VTAIL.n169 VTAIL.n168 9.3005
R1380 VTAIL.n144 VTAIL.n143 9.3005
R1381 VTAIL.n109 VTAIL.n108 9.3005
R1382 VTAIL.n138 VTAIL.n137 9.3005
R1383 VTAIL.n136 VTAIL.n135 9.3005
R1384 VTAIL.n113 VTAIL.n112 9.3005
R1385 VTAIL.n130 VTAIL.n129 9.3005
R1386 VTAIL.n128 VTAIL.n127 9.3005
R1387 VTAIL.n117 VTAIL.n116 9.3005
R1388 VTAIL.n122 VTAIL.n121 9.3005
R1389 VTAIL.n314 VTAIL.n290 8.92171
R1390 VTAIL.n330 VTAIL.n329 8.92171
R1391 VTAIL.n44 VTAIL.n20 8.92171
R1392 VTAIL.n60 VTAIL.n59 8.92171
R1393 VTAIL.n241 VTAIL.n240 8.92171
R1394 VTAIL.n225 VTAIL.n201 8.92171
R1395 VTAIL.n151 VTAIL.n150 8.92171
R1396 VTAIL.n135 VTAIL.n111 8.92171
R1397 VTAIL.n318 VTAIL.n317 8.14595
R1398 VTAIL.n326 VTAIL.n284 8.14595
R1399 VTAIL.n48 VTAIL.n47 8.14595
R1400 VTAIL.n56 VTAIL.n14 8.14595
R1401 VTAIL.n237 VTAIL.n195 8.14595
R1402 VTAIL.n229 VTAIL.n228 8.14595
R1403 VTAIL.n147 VTAIL.n105 8.14595
R1404 VTAIL.n139 VTAIL.n138 8.14595
R1405 VTAIL.n321 VTAIL.n288 7.3702
R1406 VTAIL.n325 VTAIL.n286 7.3702
R1407 VTAIL.n51 VTAIL.n18 7.3702
R1408 VTAIL.n55 VTAIL.n16 7.3702
R1409 VTAIL.n236 VTAIL.n197 7.3702
R1410 VTAIL.n232 VTAIL.n199 7.3702
R1411 VTAIL.n146 VTAIL.n107 7.3702
R1412 VTAIL.n142 VTAIL.n109 7.3702
R1413 VTAIL.n322 VTAIL.n321 6.59444
R1414 VTAIL.n322 VTAIL.n286 6.59444
R1415 VTAIL.n52 VTAIL.n51 6.59444
R1416 VTAIL.n52 VTAIL.n16 6.59444
R1417 VTAIL.n233 VTAIL.n197 6.59444
R1418 VTAIL.n233 VTAIL.n232 6.59444
R1419 VTAIL.n143 VTAIL.n107 6.59444
R1420 VTAIL.n143 VTAIL.n142 6.59444
R1421 VTAIL.n318 VTAIL.n288 5.81868
R1422 VTAIL.n326 VTAIL.n325 5.81868
R1423 VTAIL.n48 VTAIL.n18 5.81868
R1424 VTAIL.n56 VTAIL.n55 5.81868
R1425 VTAIL.n237 VTAIL.n236 5.81868
R1426 VTAIL.n229 VTAIL.n199 5.81868
R1427 VTAIL.n147 VTAIL.n146 5.81868
R1428 VTAIL.n139 VTAIL.n109 5.81868
R1429 VTAIL.n317 VTAIL.n290 5.04292
R1430 VTAIL.n329 VTAIL.n284 5.04292
R1431 VTAIL.n47 VTAIL.n20 5.04292
R1432 VTAIL.n59 VTAIL.n14 5.04292
R1433 VTAIL.n240 VTAIL.n195 5.04292
R1434 VTAIL.n228 VTAIL.n201 5.04292
R1435 VTAIL.n150 VTAIL.n105 5.04292
R1436 VTAIL.n138 VTAIL.n111 5.04292
R1437 VTAIL.n314 VTAIL.n313 4.26717
R1438 VTAIL.n330 VTAIL.n282 4.26717
R1439 VTAIL.n44 VTAIL.n43 4.26717
R1440 VTAIL.n60 VTAIL.n12 4.26717
R1441 VTAIL.n241 VTAIL.n193 4.26717
R1442 VTAIL.n225 VTAIL.n224 4.26717
R1443 VTAIL.n151 VTAIL.n103 4.26717
R1444 VTAIL.n135 VTAIL.n134 4.26717
R1445 VTAIL.n300 VTAIL.n299 3.70982
R1446 VTAIL.n30 VTAIL.n29 3.70982
R1447 VTAIL.n211 VTAIL.n210 3.70982
R1448 VTAIL.n121 VTAIL.n120 3.70982
R1449 VTAIL.n310 VTAIL.n292 3.49141
R1450 VTAIL.n334 VTAIL.n333 3.49141
R1451 VTAIL.n358 VTAIL.n270 3.49141
R1452 VTAIL.n40 VTAIL.n22 3.49141
R1453 VTAIL.n64 VTAIL.n63 3.49141
R1454 VTAIL.n88 VTAIL.n0 3.49141
R1455 VTAIL.n268 VTAIL.n180 3.49141
R1456 VTAIL.n245 VTAIL.n244 3.49141
R1457 VTAIL.n221 VTAIL.n203 3.49141
R1458 VTAIL.n178 VTAIL.n90 3.49141
R1459 VTAIL.n155 VTAIL.n154 3.49141
R1460 VTAIL.n131 VTAIL.n113 3.49141
R1461 VTAIL.n309 VTAIL.n294 2.71565
R1462 VTAIL.n337 VTAIL.n280 2.71565
R1463 VTAIL.n356 VTAIL.n355 2.71565
R1464 VTAIL.n39 VTAIL.n24 2.71565
R1465 VTAIL.n67 VTAIL.n10 2.71565
R1466 VTAIL.n86 VTAIL.n85 2.71565
R1467 VTAIL.n266 VTAIL.n265 2.71565
R1468 VTAIL.n248 VTAIL.n191 2.71565
R1469 VTAIL.n220 VTAIL.n205 2.71565
R1470 VTAIL.n176 VTAIL.n175 2.71565
R1471 VTAIL.n158 VTAIL.n101 2.71565
R1472 VTAIL.n130 VTAIL.n115 2.71565
R1473 VTAIL.n306 VTAIL.n305 1.93989
R1474 VTAIL.n338 VTAIL.n278 1.93989
R1475 VTAIL.n352 VTAIL.n272 1.93989
R1476 VTAIL.n36 VTAIL.n35 1.93989
R1477 VTAIL.n68 VTAIL.n8 1.93989
R1478 VTAIL.n82 VTAIL.n2 1.93989
R1479 VTAIL.n262 VTAIL.n182 1.93989
R1480 VTAIL.n249 VTAIL.n189 1.93989
R1481 VTAIL.n217 VTAIL.n216 1.93989
R1482 VTAIL.n172 VTAIL.n92 1.93989
R1483 VTAIL.n159 VTAIL.n99 1.93989
R1484 VTAIL.n127 VTAIL.n126 1.93989
R1485 VTAIL.n269 VTAIL.n179 1.77205
R1486 VTAIL VTAIL.n89 1.17938
R1487 VTAIL.n302 VTAIL.n296 1.16414
R1488 VTAIL.n343 VTAIL.n341 1.16414
R1489 VTAIL.n351 VTAIL.n274 1.16414
R1490 VTAIL.n32 VTAIL.n26 1.16414
R1491 VTAIL.n73 VTAIL.n71 1.16414
R1492 VTAIL.n81 VTAIL.n4 1.16414
R1493 VTAIL.n261 VTAIL.n184 1.16414
R1494 VTAIL.n253 VTAIL.n252 1.16414
R1495 VTAIL.n213 VTAIL.n207 1.16414
R1496 VTAIL.n171 VTAIL.n94 1.16414
R1497 VTAIL.n163 VTAIL.n162 1.16414
R1498 VTAIL.n123 VTAIL.n117 1.16414
R1499 VTAIL VTAIL.n359 0.593172
R1500 VTAIL.n301 VTAIL.n298 0.388379
R1501 VTAIL.n342 VTAIL.n276 0.388379
R1502 VTAIL.n348 VTAIL.n347 0.388379
R1503 VTAIL.n31 VTAIL.n28 0.388379
R1504 VTAIL.n72 VTAIL.n6 0.388379
R1505 VTAIL.n78 VTAIL.n77 0.388379
R1506 VTAIL.n258 VTAIL.n257 0.388379
R1507 VTAIL.n188 VTAIL.n186 0.388379
R1508 VTAIL.n212 VTAIL.n209 0.388379
R1509 VTAIL.n168 VTAIL.n167 0.388379
R1510 VTAIL.n98 VTAIL.n96 0.388379
R1511 VTAIL.n122 VTAIL.n119 0.388379
R1512 VTAIL.n300 VTAIL.n295 0.155672
R1513 VTAIL.n307 VTAIL.n295 0.155672
R1514 VTAIL.n308 VTAIL.n307 0.155672
R1515 VTAIL.n308 VTAIL.n291 0.155672
R1516 VTAIL.n315 VTAIL.n291 0.155672
R1517 VTAIL.n316 VTAIL.n315 0.155672
R1518 VTAIL.n316 VTAIL.n287 0.155672
R1519 VTAIL.n323 VTAIL.n287 0.155672
R1520 VTAIL.n324 VTAIL.n323 0.155672
R1521 VTAIL.n324 VTAIL.n283 0.155672
R1522 VTAIL.n331 VTAIL.n283 0.155672
R1523 VTAIL.n332 VTAIL.n331 0.155672
R1524 VTAIL.n332 VTAIL.n279 0.155672
R1525 VTAIL.n339 VTAIL.n279 0.155672
R1526 VTAIL.n340 VTAIL.n339 0.155672
R1527 VTAIL.n340 VTAIL.n275 0.155672
R1528 VTAIL.n349 VTAIL.n275 0.155672
R1529 VTAIL.n350 VTAIL.n349 0.155672
R1530 VTAIL.n350 VTAIL.n271 0.155672
R1531 VTAIL.n357 VTAIL.n271 0.155672
R1532 VTAIL.n30 VTAIL.n25 0.155672
R1533 VTAIL.n37 VTAIL.n25 0.155672
R1534 VTAIL.n38 VTAIL.n37 0.155672
R1535 VTAIL.n38 VTAIL.n21 0.155672
R1536 VTAIL.n45 VTAIL.n21 0.155672
R1537 VTAIL.n46 VTAIL.n45 0.155672
R1538 VTAIL.n46 VTAIL.n17 0.155672
R1539 VTAIL.n53 VTAIL.n17 0.155672
R1540 VTAIL.n54 VTAIL.n53 0.155672
R1541 VTAIL.n54 VTAIL.n13 0.155672
R1542 VTAIL.n61 VTAIL.n13 0.155672
R1543 VTAIL.n62 VTAIL.n61 0.155672
R1544 VTAIL.n62 VTAIL.n9 0.155672
R1545 VTAIL.n69 VTAIL.n9 0.155672
R1546 VTAIL.n70 VTAIL.n69 0.155672
R1547 VTAIL.n70 VTAIL.n5 0.155672
R1548 VTAIL.n79 VTAIL.n5 0.155672
R1549 VTAIL.n80 VTAIL.n79 0.155672
R1550 VTAIL.n80 VTAIL.n1 0.155672
R1551 VTAIL.n87 VTAIL.n1 0.155672
R1552 VTAIL.n267 VTAIL.n181 0.155672
R1553 VTAIL.n260 VTAIL.n181 0.155672
R1554 VTAIL.n260 VTAIL.n259 0.155672
R1555 VTAIL.n259 VTAIL.n185 0.155672
R1556 VTAIL.n251 VTAIL.n185 0.155672
R1557 VTAIL.n251 VTAIL.n250 0.155672
R1558 VTAIL.n250 VTAIL.n190 0.155672
R1559 VTAIL.n243 VTAIL.n190 0.155672
R1560 VTAIL.n243 VTAIL.n242 0.155672
R1561 VTAIL.n242 VTAIL.n194 0.155672
R1562 VTAIL.n235 VTAIL.n194 0.155672
R1563 VTAIL.n235 VTAIL.n234 0.155672
R1564 VTAIL.n234 VTAIL.n198 0.155672
R1565 VTAIL.n227 VTAIL.n198 0.155672
R1566 VTAIL.n227 VTAIL.n226 0.155672
R1567 VTAIL.n226 VTAIL.n202 0.155672
R1568 VTAIL.n219 VTAIL.n202 0.155672
R1569 VTAIL.n219 VTAIL.n218 0.155672
R1570 VTAIL.n218 VTAIL.n206 0.155672
R1571 VTAIL.n211 VTAIL.n206 0.155672
R1572 VTAIL.n177 VTAIL.n91 0.155672
R1573 VTAIL.n170 VTAIL.n91 0.155672
R1574 VTAIL.n170 VTAIL.n169 0.155672
R1575 VTAIL.n169 VTAIL.n95 0.155672
R1576 VTAIL.n161 VTAIL.n95 0.155672
R1577 VTAIL.n161 VTAIL.n160 0.155672
R1578 VTAIL.n160 VTAIL.n100 0.155672
R1579 VTAIL.n153 VTAIL.n100 0.155672
R1580 VTAIL.n153 VTAIL.n152 0.155672
R1581 VTAIL.n152 VTAIL.n104 0.155672
R1582 VTAIL.n145 VTAIL.n104 0.155672
R1583 VTAIL.n145 VTAIL.n144 0.155672
R1584 VTAIL.n144 VTAIL.n108 0.155672
R1585 VTAIL.n137 VTAIL.n108 0.155672
R1586 VTAIL.n137 VTAIL.n136 0.155672
R1587 VTAIL.n136 VTAIL.n112 0.155672
R1588 VTAIL.n129 VTAIL.n112 0.155672
R1589 VTAIL.n129 VTAIL.n128 0.155672
R1590 VTAIL.n128 VTAIL.n116 0.155672
R1591 VTAIL.n121 VTAIL.n116 0.155672
R1592 VDD2.n173 VDD2.n89 756.745
R1593 VDD2.n84 VDD2.n0 756.745
R1594 VDD2.n174 VDD2.n173 585
R1595 VDD2.n172 VDD2.n171 585
R1596 VDD2.n93 VDD2.n92 585
R1597 VDD2.n166 VDD2.n165 585
R1598 VDD2.n164 VDD2.n95 585
R1599 VDD2.n163 VDD2.n162 585
R1600 VDD2.n98 VDD2.n96 585
R1601 VDD2.n157 VDD2.n156 585
R1602 VDD2.n155 VDD2.n154 585
R1603 VDD2.n102 VDD2.n101 585
R1604 VDD2.n149 VDD2.n148 585
R1605 VDD2.n147 VDD2.n146 585
R1606 VDD2.n106 VDD2.n105 585
R1607 VDD2.n141 VDD2.n140 585
R1608 VDD2.n139 VDD2.n138 585
R1609 VDD2.n110 VDD2.n109 585
R1610 VDD2.n133 VDD2.n132 585
R1611 VDD2.n131 VDD2.n130 585
R1612 VDD2.n114 VDD2.n113 585
R1613 VDD2.n125 VDD2.n124 585
R1614 VDD2.n123 VDD2.n122 585
R1615 VDD2.n118 VDD2.n117 585
R1616 VDD2.n28 VDD2.n27 585
R1617 VDD2.n33 VDD2.n32 585
R1618 VDD2.n35 VDD2.n34 585
R1619 VDD2.n24 VDD2.n23 585
R1620 VDD2.n41 VDD2.n40 585
R1621 VDD2.n43 VDD2.n42 585
R1622 VDD2.n20 VDD2.n19 585
R1623 VDD2.n49 VDD2.n48 585
R1624 VDD2.n51 VDD2.n50 585
R1625 VDD2.n16 VDD2.n15 585
R1626 VDD2.n57 VDD2.n56 585
R1627 VDD2.n59 VDD2.n58 585
R1628 VDD2.n12 VDD2.n11 585
R1629 VDD2.n65 VDD2.n64 585
R1630 VDD2.n67 VDD2.n66 585
R1631 VDD2.n8 VDD2.n7 585
R1632 VDD2.n74 VDD2.n73 585
R1633 VDD2.n75 VDD2.n6 585
R1634 VDD2.n77 VDD2.n76 585
R1635 VDD2.n4 VDD2.n3 585
R1636 VDD2.n83 VDD2.n82 585
R1637 VDD2.n85 VDD2.n84 585
R1638 VDD2.n119 VDD2.t1 327.466
R1639 VDD2.n29 VDD2.t0 327.466
R1640 VDD2.n173 VDD2.n172 171.744
R1641 VDD2.n172 VDD2.n92 171.744
R1642 VDD2.n165 VDD2.n92 171.744
R1643 VDD2.n165 VDD2.n164 171.744
R1644 VDD2.n164 VDD2.n163 171.744
R1645 VDD2.n163 VDD2.n96 171.744
R1646 VDD2.n156 VDD2.n96 171.744
R1647 VDD2.n156 VDD2.n155 171.744
R1648 VDD2.n155 VDD2.n101 171.744
R1649 VDD2.n148 VDD2.n101 171.744
R1650 VDD2.n148 VDD2.n147 171.744
R1651 VDD2.n147 VDD2.n105 171.744
R1652 VDD2.n140 VDD2.n105 171.744
R1653 VDD2.n140 VDD2.n139 171.744
R1654 VDD2.n139 VDD2.n109 171.744
R1655 VDD2.n132 VDD2.n109 171.744
R1656 VDD2.n132 VDD2.n131 171.744
R1657 VDD2.n131 VDD2.n113 171.744
R1658 VDD2.n124 VDD2.n113 171.744
R1659 VDD2.n124 VDD2.n123 171.744
R1660 VDD2.n123 VDD2.n117 171.744
R1661 VDD2.n33 VDD2.n27 171.744
R1662 VDD2.n34 VDD2.n33 171.744
R1663 VDD2.n34 VDD2.n23 171.744
R1664 VDD2.n41 VDD2.n23 171.744
R1665 VDD2.n42 VDD2.n41 171.744
R1666 VDD2.n42 VDD2.n19 171.744
R1667 VDD2.n49 VDD2.n19 171.744
R1668 VDD2.n50 VDD2.n49 171.744
R1669 VDD2.n50 VDD2.n15 171.744
R1670 VDD2.n57 VDD2.n15 171.744
R1671 VDD2.n58 VDD2.n57 171.744
R1672 VDD2.n58 VDD2.n11 171.744
R1673 VDD2.n65 VDD2.n11 171.744
R1674 VDD2.n66 VDD2.n65 171.744
R1675 VDD2.n66 VDD2.n7 171.744
R1676 VDD2.n74 VDD2.n7 171.744
R1677 VDD2.n75 VDD2.n74 171.744
R1678 VDD2.n76 VDD2.n75 171.744
R1679 VDD2.n76 VDD2.n3 171.744
R1680 VDD2.n83 VDD2.n3 171.744
R1681 VDD2.n84 VDD2.n83 171.744
R1682 VDD2.n178 VDD2.n88 91.7951
R1683 VDD2.t1 VDD2.n117 85.8723
R1684 VDD2.t0 VDD2.n27 85.8723
R1685 VDD2.n178 VDD2.n177 49.0581
R1686 VDD2.n119 VDD2.n118 16.3895
R1687 VDD2.n29 VDD2.n28 16.3895
R1688 VDD2.n166 VDD2.n95 13.1884
R1689 VDD2.n77 VDD2.n6 13.1884
R1690 VDD2.n167 VDD2.n93 12.8005
R1691 VDD2.n162 VDD2.n97 12.8005
R1692 VDD2.n122 VDD2.n121 12.8005
R1693 VDD2.n32 VDD2.n31 12.8005
R1694 VDD2.n73 VDD2.n72 12.8005
R1695 VDD2.n78 VDD2.n4 12.8005
R1696 VDD2.n171 VDD2.n170 12.0247
R1697 VDD2.n161 VDD2.n98 12.0247
R1698 VDD2.n125 VDD2.n116 12.0247
R1699 VDD2.n35 VDD2.n26 12.0247
R1700 VDD2.n71 VDD2.n8 12.0247
R1701 VDD2.n82 VDD2.n81 12.0247
R1702 VDD2.n174 VDD2.n91 11.249
R1703 VDD2.n158 VDD2.n157 11.249
R1704 VDD2.n126 VDD2.n114 11.249
R1705 VDD2.n36 VDD2.n24 11.249
R1706 VDD2.n68 VDD2.n67 11.249
R1707 VDD2.n85 VDD2.n2 11.249
R1708 VDD2.n175 VDD2.n89 10.4732
R1709 VDD2.n154 VDD2.n100 10.4732
R1710 VDD2.n130 VDD2.n129 10.4732
R1711 VDD2.n40 VDD2.n39 10.4732
R1712 VDD2.n64 VDD2.n10 10.4732
R1713 VDD2.n86 VDD2.n0 10.4732
R1714 VDD2.n153 VDD2.n102 9.69747
R1715 VDD2.n133 VDD2.n112 9.69747
R1716 VDD2.n43 VDD2.n22 9.69747
R1717 VDD2.n63 VDD2.n12 9.69747
R1718 VDD2.n177 VDD2.n176 9.45567
R1719 VDD2.n88 VDD2.n87 9.45567
R1720 VDD2.n145 VDD2.n144 9.3005
R1721 VDD2.n104 VDD2.n103 9.3005
R1722 VDD2.n151 VDD2.n150 9.3005
R1723 VDD2.n153 VDD2.n152 9.3005
R1724 VDD2.n100 VDD2.n99 9.3005
R1725 VDD2.n159 VDD2.n158 9.3005
R1726 VDD2.n161 VDD2.n160 9.3005
R1727 VDD2.n97 VDD2.n94 9.3005
R1728 VDD2.n176 VDD2.n175 9.3005
R1729 VDD2.n91 VDD2.n90 9.3005
R1730 VDD2.n170 VDD2.n169 9.3005
R1731 VDD2.n168 VDD2.n167 9.3005
R1732 VDD2.n143 VDD2.n142 9.3005
R1733 VDD2.n108 VDD2.n107 9.3005
R1734 VDD2.n137 VDD2.n136 9.3005
R1735 VDD2.n135 VDD2.n134 9.3005
R1736 VDD2.n112 VDD2.n111 9.3005
R1737 VDD2.n129 VDD2.n128 9.3005
R1738 VDD2.n127 VDD2.n126 9.3005
R1739 VDD2.n116 VDD2.n115 9.3005
R1740 VDD2.n121 VDD2.n120 9.3005
R1741 VDD2.n87 VDD2.n86 9.3005
R1742 VDD2.n2 VDD2.n1 9.3005
R1743 VDD2.n81 VDD2.n80 9.3005
R1744 VDD2.n79 VDD2.n78 9.3005
R1745 VDD2.n18 VDD2.n17 9.3005
R1746 VDD2.n47 VDD2.n46 9.3005
R1747 VDD2.n45 VDD2.n44 9.3005
R1748 VDD2.n22 VDD2.n21 9.3005
R1749 VDD2.n39 VDD2.n38 9.3005
R1750 VDD2.n37 VDD2.n36 9.3005
R1751 VDD2.n26 VDD2.n25 9.3005
R1752 VDD2.n31 VDD2.n30 9.3005
R1753 VDD2.n53 VDD2.n52 9.3005
R1754 VDD2.n55 VDD2.n54 9.3005
R1755 VDD2.n14 VDD2.n13 9.3005
R1756 VDD2.n61 VDD2.n60 9.3005
R1757 VDD2.n63 VDD2.n62 9.3005
R1758 VDD2.n10 VDD2.n9 9.3005
R1759 VDD2.n69 VDD2.n68 9.3005
R1760 VDD2.n71 VDD2.n70 9.3005
R1761 VDD2.n72 VDD2.n5 9.3005
R1762 VDD2.n150 VDD2.n149 8.92171
R1763 VDD2.n134 VDD2.n110 8.92171
R1764 VDD2.n44 VDD2.n20 8.92171
R1765 VDD2.n60 VDD2.n59 8.92171
R1766 VDD2.n146 VDD2.n104 8.14595
R1767 VDD2.n138 VDD2.n137 8.14595
R1768 VDD2.n48 VDD2.n47 8.14595
R1769 VDD2.n56 VDD2.n14 8.14595
R1770 VDD2.n145 VDD2.n106 7.3702
R1771 VDD2.n141 VDD2.n108 7.3702
R1772 VDD2.n51 VDD2.n18 7.3702
R1773 VDD2.n55 VDD2.n16 7.3702
R1774 VDD2.n142 VDD2.n106 6.59444
R1775 VDD2.n142 VDD2.n141 6.59444
R1776 VDD2.n52 VDD2.n51 6.59444
R1777 VDD2.n52 VDD2.n16 6.59444
R1778 VDD2.n146 VDD2.n145 5.81868
R1779 VDD2.n138 VDD2.n108 5.81868
R1780 VDD2.n48 VDD2.n18 5.81868
R1781 VDD2.n56 VDD2.n55 5.81868
R1782 VDD2.n149 VDD2.n104 5.04292
R1783 VDD2.n137 VDD2.n110 5.04292
R1784 VDD2.n47 VDD2.n20 5.04292
R1785 VDD2.n59 VDD2.n14 5.04292
R1786 VDD2.n150 VDD2.n102 4.26717
R1787 VDD2.n134 VDD2.n133 4.26717
R1788 VDD2.n44 VDD2.n43 4.26717
R1789 VDD2.n60 VDD2.n12 4.26717
R1790 VDD2.n120 VDD2.n119 3.70982
R1791 VDD2.n30 VDD2.n29 3.70982
R1792 VDD2.n177 VDD2.n89 3.49141
R1793 VDD2.n154 VDD2.n153 3.49141
R1794 VDD2.n130 VDD2.n112 3.49141
R1795 VDD2.n40 VDD2.n22 3.49141
R1796 VDD2.n64 VDD2.n63 3.49141
R1797 VDD2.n88 VDD2.n0 3.49141
R1798 VDD2.n175 VDD2.n174 2.71565
R1799 VDD2.n157 VDD2.n100 2.71565
R1800 VDD2.n129 VDD2.n114 2.71565
R1801 VDD2.n39 VDD2.n24 2.71565
R1802 VDD2.n67 VDD2.n10 2.71565
R1803 VDD2.n86 VDD2.n85 2.71565
R1804 VDD2.n171 VDD2.n91 1.93989
R1805 VDD2.n158 VDD2.n98 1.93989
R1806 VDD2.n126 VDD2.n125 1.93989
R1807 VDD2.n36 VDD2.n35 1.93989
R1808 VDD2.n68 VDD2.n8 1.93989
R1809 VDD2.n82 VDD2.n2 1.93989
R1810 VDD2.n170 VDD2.n93 1.16414
R1811 VDD2.n162 VDD2.n161 1.16414
R1812 VDD2.n122 VDD2.n116 1.16414
R1813 VDD2.n32 VDD2.n26 1.16414
R1814 VDD2.n73 VDD2.n71 1.16414
R1815 VDD2.n81 VDD2.n4 1.16414
R1816 VDD2 VDD2.n178 0.709552
R1817 VDD2.n167 VDD2.n166 0.388379
R1818 VDD2.n97 VDD2.n95 0.388379
R1819 VDD2.n121 VDD2.n118 0.388379
R1820 VDD2.n31 VDD2.n28 0.388379
R1821 VDD2.n72 VDD2.n6 0.388379
R1822 VDD2.n78 VDD2.n77 0.388379
R1823 VDD2.n176 VDD2.n90 0.155672
R1824 VDD2.n169 VDD2.n90 0.155672
R1825 VDD2.n169 VDD2.n168 0.155672
R1826 VDD2.n168 VDD2.n94 0.155672
R1827 VDD2.n160 VDD2.n94 0.155672
R1828 VDD2.n160 VDD2.n159 0.155672
R1829 VDD2.n159 VDD2.n99 0.155672
R1830 VDD2.n152 VDD2.n99 0.155672
R1831 VDD2.n152 VDD2.n151 0.155672
R1832 VDD2.n151 VDD2.n103 0.155672
R1833 VDD2.n144 VDD2.n103 0.155672
R1834 VDD2.n144 VDD2.n143 0.155672
R1835 VDD2.n143 VDD2.n107 0.155672
R1836 VDD2.n136 VDD2.n107 0.155672
R1837 VDD2.n136 VDD2.n135 0.155672
R1838 VDD2.n135 VDD2.n111 0.155672
R1839 VDD2.n128 VDD2.n111 0.155672
R1840 VDD2.n128 VDD2.n127 0.155672
R1841 VDD2.n127 VDD2.n115 0.155672
R1842 VDD2.n120 VDD2.n115 0.155672
R1843 VDD2.n30 VDD2.n25 0.155672
R1844 VDD2.n37 VDD2.n25 0.155672
R1845 VDD2.n38 VDD2.n37 0.155672
R1846 VDD2.n38 VDD2.n21 0.155672
R1847 VDD2.n45 VDD2.n21 0.155672
R1848 VDD2.n46 VDD2.n45 0.155672
R1849 VDD2.n46 VDD2.n17 0.155672
R1850 VDD2.n53 VDD2.n17 0.155672
R1851 VDD2.n54 VDD2.n53 0.155672
R1852 VDD2.n54 VDD2.n13 0.155672
R1853 VDD2.n61 VDD2.n13 0.155672
R1854 VDD2.n62 VDD2.n61 0.155672
R1855 VDD2.n62 VDD2.n9 0.155672
R1856 VDD2.n69 VDD2.n9 0.155672
R1857 VDD2.n70 VDD2.n69 0.155672
R1858 VDD2.n70 VDD2.n5 0.155672
R1859 VDD2.n79 VDD2.n5 0.155672
R1860 VDD2.n80 VDD2.n79 0.155672
R1861 VDD2.n80 VDD2.n1 0.155672
R1862 VDD2.n87 VDD2.n1 0.155672
R1863 VP.n0 VP.t0 233.243
R1864 VP.n0 VP.t1 185.249
R1865 VP VP.n0 0.431811
R1866 VDD1.n84 VDD1.n0 756.745
R1867 VDD1.n173 VDD1.n89 756.745
R1868 VDD1.n85 VDD1.n84 585
R1869 VDD1.n83 VDD1.n82 585
R1870 VDD1.n4 VDD1.n3 585
R1871 VDD1.n77 VDD1.n76 585
R1872 VDD1.n75 VDD1.n6 585
R1873 VDD1.n74 VDD1.n73 585
R1874 VDD1.n9 VDD1.n7 585
R1875 VDD1.n68 VDD1.n67 585
R1876 VDD1.n66 VDD1.n65 585
R1877 VDD1.n13 VDD1.n12 585
R1878 VDD1.n60 VDD1.n59 585
R1879 VDD1.n58 VDD1.n57 585
R1880 VDD1.n17 VDD1.n16 585
R1881 VDD1.n52 VDD1.n51 585
R1882 VDD1.n50 VDD1.n49 585
R1883 VDD1.n21 VDD1.n20 585
R1884 VDD1.n44 VDD1.n43 585
R1885 VDD1.n42 VDD1.n41 585
R1886 VDD1.n25 VDD1.n24 585
R1887 VDD1.n36 VDD1.n35 585
R1888 VDD1.n34 VDD1.n33 585
R1889 VDD1.n29 VDD1.n28 585
R1890 VDD1.n117 VDD1.n116 585
R1891 VDD1.n122 VDD1.n121 585
R1892 VDD1.n124 VDD1.n123 585
R1893 VDD1.n113 VDD1.n112 585
R1894 VDD1.n130 VDD1.n129 585
R1895 VDD1.n132 VDD1.n131 585
R1896 VDD1.n109 VDD1.n108 585
R1897 VDD1.n138 VDD1.n137 585
R1898 VDD1.n140 VDD1.n139 585
R1899 VDD1.n105 VDD1.n104 585
R1900 VDD1.n146 VDD1.n145 585
R1901 VDD1.n148 VDD1.n147 585
R1902 VDD1.n101 VDD1.n100 585
R1903 VDD1.n154 VDD1.n153 585
R1904 VDD1.n156 VDD1.n155 585
R1905 VDD1.n97 VDD1.n96 585
R1906 VDD1.n163 VDD1.n162 585
R1907 VDD1.n164 VDD1.n95 585
R1908 VDD1.n166 VDD1.n165 585
R1909 VDD1.n93 VDD1.n92 585
R1910 VDD1.n172 VDD1.n171 585
R1911 VDD1.n174 VDD1.n173 585
R1912 VDD1.n30 VDD1.t1 327.466
R1913 VDD1.n118 VDD1.t0 327.466
R1914 VDD1.n84 VDD1.n83 171.744
R1915 VDD1.n83 VDD1.n3 171.744
R1916 VDD1.n76 VDD1.n3 171.744
R1917 VDD1.n76 VDD1.n75 171.744
R1918 VDD1.n75 VDD1.n74 171.744
R1919 VDD1.n74 VDD1.n7 171.744
R1920 VDD1.n67 VDD1.n7 171.744
R1921 VDD1.n67 VDD1.n66 171.744
R1922 VDD1.n66 VDD1.n12 171.744
R1923 VDD1.n59 VDD1.n12 171.744
R1924 VDD1.n59 VDD1.n58 171.744
R1925 VDD1.n58 VDD1.n16 171.744
R1926 VDD1.n51 VDD1.n16 171.744
R1927 VDD1.n51 VDD1.n50 171.744
R1928 VDD1.n50 VDD1.n20 171.744
R1929 VDD1.n43 VDD1.n20 171.744
R1930 VDD1.n43 VDD1.n42 171.744
R1931 VDD1.n42 VDD1.n24 171.744
R1932 VDD1.n35 VDD1.n24 171.744
R1933 VDD1.n35 VDD1.n34 171.744
R1934 VDD1.n34 VDD1.n28 171.744
R1935 VDD1.n122 VDD1.n116 171.744
R1936 VDD1.n123 VDD1.n122 171.744
R1937 VDD1.n123 VDD1.n112 171.744
R1938 VDD1.n130 VDD1.n112 171.744
R1939 VDD1.n131 VDD1.n130 171.744
R1940 VDD1.n131 VDD1.n108 171.744
R1941 VDD1.n138 VDD1.n108 171.744
R1942 VDD1.n139 VDD1.n138 171.744
R1943 VDD1.n139 VDD1.n104 171.744
R1944 VDD1.n146 VDD1.n104 171.744
R1945 VDD1.n147 VDD1.n146 171.744
R1946 VDD1.n147 VDD1.n100 171.744
R1947 VDD1.n154 VDD1.n100 171.744
R1948 VDD1.n155 VDD1.n154 171.744
R1949 VDD1.n155 VDD1.n96 171.744
R1950 VDD1.n163 VDD1.n96 171.744
R1951 VDD1.n164 VDD1.n163 171.744
R1952 VDD1.n165 VDD1.n164 171.744
R1953 VDD1.n165 VDD1.n92 171.744
R1954 VDD1.n172 VDD1.n92 171.744
R1955 VDD1.n173 VDD1.n172 171.744
R1956 VDD1 VDD1.n177 92.9708
R1957 VDD1.t1 VDD1.n28 85.8723
R1958 VDD1.t0 VDD1.n116 85.8723
R1959 VDD1 VDD1.n88 49.7671
R1960 VDD1.n30 VDD1.n29 16.3895
R1961 VDD1.n118 VDD1.n117 16.3895
R1962 VDD1.n77 VDD1.n6 13.1884
R1963 VDD1.n166 VDD1.n95 13.1884
R1964 VDD1.n78 VDD1.n4 12.8005
R1965 VDD1.n73 VDD1.n8 12.8005
R1966 VDD1.n33 VDD1.n32 12.8005
R1967 VDD1.n121 VDD1.n120 12.8005
R1968 VDD1.n162 VDD1.n161 12.8005
R1969 VDD1.n167 VDD1.n93 12.8005
R1970 VDD1.n82 VDD1.n81 12.0247
R1971 VDD1.n72 VDD1.n9 12.0247
R1972 VDD1.n36 VDD1.n27 12.0247
R1973 VDD1.n124 VDD1.n115 12.0247
R1974 VDD1.n160 VDD1.n97 12.0247
R1975 VDD1.n171 VDD1.n170 12.0247
R1976 VDD1.n85 VDD1.n2 11.249
R1977 VDD1.n69 VDD1.n68 11.249
R1978 VDD1.n37 VDD1.n25 11.249
R1979 VDD1.n125 VDD1.n113 11.249
R1980 VDD1.n157 VDD1.n156 11.249
R1981 VDD1.n174 VDD1.n91 11.249
R1982 VDD1.n86 VDD1.n0 10.4732
R1983 VDD1.n65 VDD1.n11 10.4732
R1984 VDD1.n41 VDD1.n40 10.4732
R1985 VDD1.n129 VDD1.n128 10.4732
R1986 VDD1.n153 VDD1.n99 10.4732
R1987 VDD1.n175 VDD1.n89 10.4732
R1988 VDD1.n64 VDD1.n13 9.69747
R1989 VDD1.n44 VDD1.n23 9.69747
R1990 VDD1.n132 VDD1.n111 9.69747
R1991 VDD1.n152 VDD1.n101 9.69747
R1992 VDD1.n88 VDD1.n87 9.45567
R1993 VDD1.n177 VDD1.n176 9.45567
R1994 VDD1.n56 VDD1.n55 9.3005
R1995 VDD1.n15 VDD1.n14 9.3005
R1996 VDD1.n62 VDD1.n61 9.3005
R1997 VDD1.n64 VDD1.n63 9.3005
R1998 VDD1.n11 VDD1.n10 9.3005
R1999 VDD1.n70 VDD1.n69 9.3005
R2000 VDD1.n72 VDD1.n71 9.3005
R2001 VDD1.n8 VDD1.n5 9.3005
R2002 VDD1.n87 VDD1.n86 9.3005
R2003 VDD1.n2 VDD1.n1 9.3005
R2004 VDD1.n81 VDD1.n80 9.3005
R2005 VDD1.n79 VDD1.n78 9.3005
R2006 VDD1.n54 VDD1.n53 9.3005
R2007 VDD1.n19 VDD1.n18 9.3005
R2008 VDD1.n48 VDD1.n47 9.3005
R2009 VDD1.n46 VDD1.n45 9.3005
R2010 VDD1.n23 VDD1.n22 9.3005
R2011 VDD1.n40 VDD1.n39 9.3005
R2012 VDD1.n38 VDD1.n37 9.3005
R2013 VDD1.n27 VDD1.n26 9.3005
R2014 VDD1.n32 VDD1.n31 9.3005
R2015 VDD1.n176 VDD1.n175 9.3005
R2016 VDD1.n91 VDD1.n90 9.3005
R2017 VDD1.n170 VDD1.n169 9.3005
R2018 VDD1.n168 VDD1.n167 9.3005
R2019 VDD1.n107 VDD1.n106 9.3005
R2020 VDD1.n136 VDD1.n135 9.3005
R2021 VDD1.n134 VDD1.n133 9.3005
R2022 VDD1.n111 VDD1.n110 9.3005
R2023 VDD1.n128 VDD1.n127 9.3005
R2024 VDD1.n126 VDD1.n125 9.3005
R2025 VDD1.n115 VDD1.n114 9.3005
R2026 VDD1.n120 VDD1.n119 9.3005
R2027 VDD1.n142 VDD1.n141 9.3005
R2028 VDD1.n144 VDD1.n143 9.3005
R2029 VDD1.n103 VDD1.n102 9.3005
R2030 VDD1.n150 VDD1.n149 9.3005
R2031 VDD1.n152 VDD1.n151 9.3005
R2032 VDD1.n99 VDD1.n98 9.3005
R2033 VDD1.n158 VDD1.n157 9.3005
R2034 VDD1.n160 VDD1.n159 9.3005
R2035 VDD1.n161 VDD1.n94 9.3005
R2036 VDD1.n61 VDD1.n60 8.92171
R2037 VDD1.n45 VDD1.n21 8.92171
R2038 VDD1.n133 VDD1.n109 8.92171
R2039 VDD1.n149 VDD1.n148 8.92171
R2040 VDD1.n57 VDD1.n15 8.14595
R2041 VDD1.n49 VDD1.n48 8.14595
R2042 VDD1.n137 VDD1.n136 8.14595
R2043 VDD1.n145 VDD1.n103 8.14595
R2044 VDD1.n56 VDD1.n17 7.3702
R2045 VDD1.n52 VDD1.n19 7.3702
R2046 VDD1.n140 VDD1.n107 7.3702
R2047 VDD1.n144 VDD1.n105 7.3702
R2048 VDD1.n53 VDD1.n17 6.59444
R2049 VDD1.n53 VDD1.n52 6.59444
R2050 VDD1.n141 VDD1.n140 6.59444
R2051 VDD1.n141 VDD1.n105 6.59444
R2052 VDD1.n57 VDD1.n56 5.81868
R2053 VDD1.n49 VDD1.n19 5.81868
R2054 VDD1.n137 VDD1.n107 5.81868
R2055 VDD1.n145 VDD1.n144 5.81868
R2056 VDD1.n60 VDD1.n15 5.04292
R2057 VDD1.n48 VDD1.n21 5.04292
R2058 VDD1.n136 VDD1.n109 5.04292
R2059 VDD1.n148 VDD1.n103 5.04292
R2060 VDD1.n61 VDD1.n13 4.26717
R2061 VDD1.n45 VDD1.n44 4.26717
R2062 VDD1.n133 VDD1.n132 4.26717
R2063 VDD1.n149 VDD1.n101 4.26717
R2064 VDD1.n31 VDD1.n30 3.70982
R2065 VDD1.n119 VDD1.n118 3.70982
R2066 VDD1.n88 VDD1.n0 3.49141
R2067 VDD1.n65 VDD1.n64 3.49141
R2068 VDD1.n41 VDD1.n23 3.49141
R2069 VDD1.n129 VDD1.n111 3.49141
R2070 VDD1.n153 VDD1.n152 3.49141
R2071 VDD1.n177 VDD1.n89 3.49141
R2072 VDD1.n86 VDD1.n85 2.71565
R2073 VDD1.n68 VDD1.n11 2.71565
R2074 VDD1.n40 VDD1.n25 2.71565
R2075 VDD1.n128 VDD1.n113 2.71565
R2076 VDD1.n156 VDD1.n99 2.71565
R2077 VDD1.n175 VDD1.n174 2.71565
R2078 VDD1.n82 VDD1.n2 1.93989
R2079 VDD1.n69 VDD1.n9 1.93989
R2080 VDD1.n37 VDD1.n36 1.93989
R2081 VDD1.n125 VDD1.n124 1.93989
R2082 VDD1.n157 VDD1.n97 1.93989
R2083 VDD1.n171 VDD1.n91 1.93989
R2084 VDD1.n81 VDD1.n4 1.16414
R2085 VDD1.n73 VDD1.n72 1.16414
R2086 VDD1.n33 VDD1.n27 1.16414
R2087 VDD1.n121 VDD1.n115 1.16414
R2088 VDD1.n162 VDD1.n160 1.16414
R2089 VDD1.n170 VDD1.n93 1.16414
R2090 VDD1.n78 VDD1.n77 0.388379
R2091 VDD1.n8 VDD1.n6 0.388379
R2092 VDD1.n32 VDD1.n29 0.388379
R2093 VDD1.n120 VDD1.n117 0.388379
R2094 VDD1.n161 VDD1.n95 0.388379
R2095 VDD1.n167 VDD1.n166 0.388379
R2096 VDD1.n87 VDD1.n1 0.155672
R2097 VDD1.n80 VDD1.n1 0.155672
R2098 VDD1.n80 VDD1.n79 0.155672
R2099 VDD1.n79 VDD1.n5 0.155672
R2100 VDD1.n71 VDD1.n5 0.155672
R2101 VDD1.n71 VDD1.n70 0.155672
R2102 VDD1.n70 VDD1.n10 0.155672
R2103 VDD1.n63 VDD1.n10 0.155672
R2104 VDD1.n63 VDD1.n62 0.155672
R2105 VDD1.n62 VDD1.n14 0.155672
R2106 VDD1.n55 VDD1.n14 0.155672
R2107 VDD1.n55 VDD1.n54 0.155672
R2108 VDD1.n54 VDD1.n18 0.155672
R2109 VDD1.n47 VDD1.n18 0.155672
R2110 VDD1.n47 VDD1.n46 0.155672
R2111 VDD1.n46 VDD1.n22 0.155672
R2112 VDD1.n39 VDD1.n22 0.155672
R2113 VDD1.n39 VDD1.n38 0.155672
R2114 VDD1.n38 VDD1.n26 0.155672
R2115 VDD1.n31 VDD1.n26 0.155672
R2116 VDD1.n119 VDD1.n114 0.155672
R2117 VDD1.n126 VDD1.n114 0.155672
R2118 VDD1.n127 VDD1.n126 0.155672
R2119 VDD1.n127 VDD1.n110 0.155672
R2120 VDD1.n134 VDD1.n110 0.155672
R2121 VDD1.n135 VDD1.n134 0.155672
R2122 VDD1.n135 VDD1.n106 0.155672
R2123 VDD1.n142 VDD1.n106 0.155672
R2124 VDD1.n143 VDD1.n142 0.155672
R2125 VDD1.n143 VDD1.n102 0.155672
R2126 VDD1.n150 VDD1.n102 0.155672
R2127 VDD1.n151 VDD1.n150 0.155672
R2128 VDD1.n151 VDD1.n98 0.155672
R2129 VDD1.n158 VDD1.n98 0.155672
R2130 VDD1.n159 VDD1.n158 0.155672
R2131 VDD1.n159 VDD1.n94 0.155672
R2132 VDD1.n168 VDD1.n94 0.155672
R2133 VDD1.n169 VDD1.n168 0.155672
R2134 VDD1.n169 VDD1.n90 0.155672
R2135 VDD1.n176 VDD1.n90 0.155672
C0 w_n2178_n4186# B 10.052701f
C1 VDD1 VN 0.148163f
C2 VDD1 VDD2 0.685926f
C3 VDD1 B 2.04161f
C4 w_n2178_n4186# VTAIL 3.3127f
C5 VN VP 6.25868f
C6 VP VDD2 0.337162f
C7 VP B 1.5699f
C8 VDD1 VTAIL 6.15448f
C9 VP VTAIL 3.16546f
C10 VDD1 w_n2178_n4186# 2.07473f
C11 VN VDD2 3.66189f
C12 VN B 1.11311f
C13 B VDD2 2.07249f
C14 VP w_n2178_n4186# 3.38331f
C15 VN VTAIL 3.15112f
C16 VDD2 VTAIL 6.20487f
C17 B VTAIL 4.61525f
C18 VDD1 VP 3.84771f
C19 VN w_n2178_n4186# 3.10568f
C20 w_n2178_n4186# VDD2 2.10172f
C21 VDD2 VSUBS 1.077301f
C22 VDD1 VSUBS 5.34646f
C23 VTAIL VSUBS 1.170942f
C24 VN VSUBS 8.80534f
C25 VP VSUBS 1.86423f
C26 B VSUBS 4.322153f
C27 w_n2178_n4186# VSUBS 0.111679p
C28 VDD1.n0 VSUBS 0.029761f
C29 VDD1.n1 VSUBS 0.028398f
C30 VDD1.n2 VSUBS 0.01526f
C31 VDD1.n3 VSUBS 0.036069f
C32 VDD1.n4 VSUBS 0.016158f
C33 VDD1.n5 VSUBS 0.028398f
C34 VDD1.n6 VSUBS 0.015709f
C35 VDD1.n7 VSUBS 0.036069f
C36 VDD1.n8 VSUBS 0.01526f
C37 VDD1.n9 VSUBS 0.016158f
C38 VDD1.n10 VSUBS 0.028398f
C39 VDD1.n11 VSUBS 0.01526f
C40 VDD1.n12 VSUBS 0.036069f
C41 VDD1.n13 VSUBS 0.016158f
C42 VDD1.n14 VSUBS 0.028398f
C43 VDD1.n15 VSUBS 0.01526f
C44 VDD1.n16 VSUBS 0.036069f
C45 VDD1.n17 VSUBS 0.016158f
C46 VDD1.n18 VSUBS 0.028398f
C47 VDD1.n19 VSUBS 0.01526f
C48 VDD1.n20 VSUBS 0.036069f
C49 VDD1.n21 VSUBS 0.016158f
C50 VDD1.n22 VSUBS 0.028398f
C51 VDD1.n23 VSUBS 0.01526f
C52 VDD1.n24 VSUBS 0.036069f
C53 VDD1.n25 VSUBS 0.016158f
C54 VDD1.n26 VSUBS 0.028398f
C55 VDD1.n27 VSUBS 0.01526f
C56 VDD1.n28 VSUBS 0.027052f
C57 VDD1.n29 VSUBS 0.022945f
C58 VDD1.t1 VSUBS 0.077293f
C59 VDD1.n30 VSUBS 0.209313f
C60 VDD1.n31 VSUBS 1.95381f
C61 VDD1.n32 VSUBS 0.01526f
C62 VDD1.n33 VSUBS 0.016158f
C63 VDD1.n34 VSUBS 0.036069f
C64 VDD1.n35 VSUBS 0.036069f
C65 VDD1.n36 VSUBS 0.016158f
C66 VDD1.n37 VSUBS 0.01526f
C67 VDD1.n38 VSUBS 0.028398f
C68 VDD1.n39 VSUBS 0.028398f
C69 VDD1.n40 VSUBS 0.01526f
C70 VDD1.n41 VSUBS 0.016158f
C71 VDD1.n42 VSUBS 0.036069f
C72 VDD1.n43 VSUBS 0.036069f
C73 VDD1.n44 VSUBS 0.016158f
C74 VDD1.n45 VSUBS 0.01526f
C75 VDD1.n46 VSUBS 0.028398f
C76 VDD1.n47 VSUBS 0.028398f
C77 VDD1.n48 VSUBS 0.01526f
C78 VDD1.n49 VSUBS 0.016158f
C79 VDD1.n50 VSUBS 0.036069f
C80 VDD1.n51 VSUBS 0.036069f
C81 VDD1.n52 VSUBS 0.016158f
C82 VDD1.n53 VSUBS 0.01526f
C83 VDD1.n54 VSUBS 0.028398f
C84 VDD1.n55 VSUBS 0.028398f
C85 VDD1.n56 VSUBS 0.01526f
C86 VDD1.n57 VSUBS 0.016158f
C87 VDD1.n58 VSUBS 0.036069f
C88 VDD1.n59 VSUBS 0.036069f
C89 VDD1.n60 VSUBS 0.016158f
C90 VDD1.n61 VSUBS 0.01526f
C91 VDD1.n62 VSUBS 0.028398f
C92 VDD1.n63 VSUBS 0.028398f
C93 VDD1.n64 VSUBS 0.01526f
C94 VDD1.n65 VSUBS 0.016158f
C95 VDD1.n66 VSUBS 0.036069f
C96 VDD1.n67 VSUBS 0.036069f
C97 VDD1.n68 VSUBS 0.016158f
C98 VDD1.n69 VSUBS 0.01526f
C99 VDD1.n70 VSUBS 0.028398f
C100 VDD1.n71 VSUBS 0.028398f
C101 VDD1.n72 VSUBS 0.01526f
C102 VDD1.n73 VSUBS 0.016158f
C103 VDD1.n74 VSUBS 0.036069f
C104 VDD1.n75 VSUBS 0.036069f
C105 VDD1.n76 VSUBS 0.036069f
C106 VDD1.n77 VSUBS 0.015709f
C107 VDD1.n78 VSUBS 0.01526f
C108 VDD1.n79 VSUBS 0.028398f
C109 VDD1.n80 VSUBS 0.028398f
C110 VDD1.n81 VSUBS 0.01526f
C111 VDD1.n82 VSUBS 0.016158f
C112 VDD1.n83 VSUBS 0.036069f
C113 VDD1.n84 VSUBS 0.082404f
C114 VDD1.n85 VSUBS 0.016158f
C115 VDD1.n86 VSUBS 0.01526f
C116 VDD1.n87 VSUBS 0.066029f
C117 VDD1.n88 VSUBS 0.062546f
C118 VDD1.n89 VSUBS 0.029761f
C119 VDD1.n90 VSUBS 0.028398f
C120 VDD1.n91 VSUBS 0.01526f
C121 VDD1.n92 VSUBS 0.036069f
C122 VDD1.n93 VSUBS 0.016158f
C123 VDD1.n94 VSUBS 0.028398f
C124 VDD1.n95 VSUBS 0.015709f
C125 VDD1.n96 VSUBS 0.036069f
C126 VDD1.n97 VSUBS 0.016158f
C127 VDD1.n98 VSUBS 0.028398f
C128 VDD1.n99 VSUBS 0.01526f
C129 VDD1.n100 VSUBS 0.036069f
C130 VDD1.n101 VSUBS 0.016158f
C131 VDD1.n102 VSUBS 0.028398f
C132 VDD1.n103 VSUBS 0.01526f
C133 VDD1.n104 VSUBS 0.036069f
C134 VDD1.n105 VSUBS 0.016158f
C135 VDD1.n106 VSUBS 0.028398f
C136 VDD1.n107 VSUBS 0.01526f
C137 VDD1.n108 VSUBS 0.036069f
C138 VDD1.n109 VSUBS 0.016158f
C139 VDD1.n110 VSUBS 0.028398f
C140 VDD1.n111 VSUBS 0.01526f
C141 VDD1.n112 VSUBS 0.036069f
C142 VDD1.n113 VSUBS 0.016158f
C143 VDD1.n114 VSUBS 0.028398f
C144 VDD1.n115 VSUBS 0.01526f
C145 VDD1.n116 VSUBS 0.027052f
C146 VDD1.n117 VSUBS 0.022945f
C147 VDD1.t0 VSUBS 0.077293f
C148 VDD1.n118 VSUBS 0.209313f
C149 VDD1.n119 VSUBS 1.95381f
C150 VDD1.n120 VSUBS 0.01526f
C151 VDD1.n121 VSUBS 0.016158f
C152 VDD1.n122 VSUBS 0.036069f
C153 VDD1.n123 VSUBS 0.036069f
C154 VDD1.n124 VSUBS 0.016158f
C155 VDD1.n125 VSUBS 0.01526f
C156 VDD1.n126 VSUBS 0.028398f
C157 VDD1.n127 VSUBS 0.028398f
C158 VDD1.n128 VSUBS 0.01526f
C159 VDD1.n129 VSUBS 0.016158f
C160 VDD1.n130 VSUBS 0.036069f
C161 VDD1.n131 VSUBS 0.036069f
C162 VDD1.n132 VSUBS 0.016158f
C163 VDD1.n133 VSUBS 0.01526f
C164 VDD1.n134 VSUBS 0.028398f
C165 VDD1.n135 VSUBS 0.028398f
C166 VDD1.n136 VSUBS 0.01526f
C167 VDD1.n137 VSUBS 0.016158f
C168 VDD1.n138 VSUBS 0.036069f
C169 VDD1.n139 VSUBS 0.036069f
C170 VDD1.n140 VSUBS 0.016158f
C171 VDD1.n141 VSUBS 0.01526f
C172 VDD1.n142 VSUBS 0.028398f
C173 VDD1.n143 VSUBS 0.028398f
C174 VDD1.n144 VSUBS 0.01526f
C175 VDD1.n145 VSUBS 0.016158f
C176 VDD1.n146 VSUBS 0.036069f
C177 VDD1.n147 VSUBS 0.036069f
C178 VDD1.n148 VSUBS 0.016158f
C179 VDD1.n149 VSUBS 0.01526f
C180 VDD1.n150 VSUBS 0.028398f
C181 VDD1.n151 VSUBS 0.028398f
C182 VDD1.n152 VSUBS 0.01526f
C183 VDD1.n153 VSUBS 0.016158f
C184 VDD1.n154 VSUBS 0.036069f
C185 VDD1.n155 VSUBS 0.036069f
C186 VDD1.n156 VSUBS 0.016158f
C187 VDD1.n157 VSUBS 0.01526f
C188 VDD1.n158 VSUBS 0.028398f
C189 VDD1.n159 VSUBS 0.028398f
C190 VDD1.n160 VSUBS 0.01526f
C191 VDD1.n161 VSUBS 0.01526f
C192 VDD1.n162 VSUBS 0.016158f
C193 VDD1.n163 VSUBS 0.036069f
C194 VDD1.n164 VSUBS 0.036069f
C195 VDD1.n165 VSUBS 0.036069f
C196 VDD1.n166 VSUBS 0.015709f
C197 VDD1.n167 VSUBS 0.01526f
C198 VDD1.n168 VSUBS 0.028398f
C199 VDD1.n169 VSUBS 0.028398f
C200 VDD1.n170 VSUBS 0.01526f
C201 VDD1.n171 VSUBS 0.016158f
C202 VDD1.n172 VSUBS 0.036069f
C203 VDD1.n173 VSUBS 0.082404f
C204 VDD1.n174 VSUBS 0.016158f
C205 VDD1.n175 VSUBS 0.01526f
C206 VDD1.n176 VSUBS 0.066029f
C207 VDD1.n177 VSUBS 1.06884f
C208 VP.t1 VSUBS 4.83555f
C209 VP.t0 VSUBS 5.55584f
C210 VP.n0 VSUBS 6.20948f
C211 VDD2.n0 VSUBS 0.029984f
C212 VDD2.n1 VSUBS 0.028611f
C213 VDD2.n2 VSUBS 0.015374f
C214 VDD2.n3 VSUBS 0.036339f
C215 VDD2.n4 VSUBS 0.016279f
C216 VDD2.n5 VSUBS 0.028611f
C217 VDD2.n6 VSUBS 0.015826f
C218 VDD2.n7 VSUBS 0.036339f
C219 VDD2.n8 VSUBS 0.016279f
C220 VDD2.n9 VSUBS 0.028611f
C221 VDD2.n10 VSUBS 0.015374f
C222 VDD2.n11 VSUBS 0.036339f
C223 VDD2.n12 VSUBS 0.016279f
C224 VDD2.n13 VSUBS 0.028611f
C225 VDD2.n14 VSUBS 0.015374f
C226 VDD2.n15 VSUBS 0.036339f
C227 VDD2.n16 VSUBS 0.016279f
C228 VDD2.n17 VSUBS 0.028611f
C229 VDD2.n18 VSUBS 0.015374f
C230 VDD2.n19 VSUBS 0.036339f
C231 VDD2.n20 VSUBS 0.016279f
C232 VDD2.n21 VSUBS 0.028611f
C233 VDD2.n22 VSUBS 0.015374f
C234 VDD2.n23 VSUBS 0.036339f
C235 VDD2.n24 VSUBS 0.016279f
C236 VDD2.n25 VSUBS 0.028611f
C237 VDD2.n26 VSUBS 0.015374f
C238 VDD2.n27 VSUBS 0.027254f
C239 VDD2.n28 VSUBS 0.023117f
C240 VDD2.t0 VSUBS 0.077873f
C241 VDD2.n29 VSUBS 0.210882f
C242 VDD2.n30 VSUBS 1.96845f
C243 VDD2.n31 VSUBS 0.015374f
C244 VDD2.n32 VSUBS 0.016279f
C245 VDD2.n33 VSUBS 0.036339f
C246 VDD2.n34 VSUBS 0.036339f
C247 VDD2.n35 VSUBS 0.016279f
C248 VDD2.n36 VSUBS 0.015374f
C249 VDD2.n37 VSUBS 0.028611f
C250 VDD2.n38 VSUBS 0.028611f
C251 VDD2.n39 VSUBS 0.015374f
C252 VDD2.n40 VSUBS 0.016279f
C253 VDD2.n41 VSUBS 0.036339f
C254 VDD2.n42 VSUBS 0.036339f
C255 VDD2.n43 VSUBS 0.016279f
C256 VDD2.n44 VSUBS 0.015374f
C257 VDD2.n45 VSUBS 0.028611f
C258 VDD2.n46 VSUBS 0.028611f
C259 VDD2.n47 VSUBS 0.015374f
C260 VDD2.n48 VSUBS 0.016279f
C261 VDD2.n49 VSUBS 0.036339f
C262 VDD2.n50 VSUBS 0.036339f
C263 VDD2.n51 VSUBS 0.016279f
C264 VDD2.n52 VSUBS 0.015374f
C265 VDD2.n53 VSUBS 0.028611f
C266 VDD2.n54 VSUBS 0.028611f
C267 VDD2.n55 VSUBS 0.015374f
C268 VDD2.n56 VSUBS 0.016279f
C269 VDD2.n57 VSUBS 0.036339f
C270 VDD2.n58 VSUBS 0.036339f
C271 VDD2.n59 VSUBS 0.016279f
C272 VDD2.n60 VSUBS 0.015374f
C273 VDD2.n61 VSUBS 0.028611f
C274 VDD2.n62 VSUBS 0.028611f
C275 VDD2.n63 VSUBS 0.015374f
C276 VDD2.n64 VSUBS 0.016279f
C277 VDD2.n65 VSUBS 0.036339f
C278 VDD2.n66 VSUBS 0.036339f
C279 VDD2.n67 VSUBS 0.016279f
C280 VDD2.n68 VSUBS 0.015374f
C281 VDD2.n69 VSUBS 0.028611f
C282 VDD2.n70 VSUBS 0.028611f
C283 VDD2.n71 VSUBS 0.015374f
C284 VDD2.n72 VSUBS 0.015374f
C285 VDD2.n73 VSUBS 0.016279f
C286 VDD2.n74 VSUBS 0.036339f
C287 VDD2.n75 VSUBS 0.036339f
C288 VDD2.n76 VSUBS 0.036339f
C289 VDD2.n77 VSUBS 0.015826f
C290 VDD2.n78 VSUBS 0.015374f
C291 VDD2.n79 VSUBS 0.028611f
C292 VDD2.n80 VSUBS 0.028611f
C293 VDD2.n81 VSUBS 0.015374f
C294 VDD2.n82 VSUBS 0.016279f
C295 VDD2.n83 VSUBS 0.036339f
C296 VDD2.n84 VSUBS 0.083022f
C297 VDD2.n85 VSUBS 0.016279f
C298 VDD2.n86 VSUBS 0.015374f
C299 VDD2.n87 VSUBS 0.066524f
C300 VDD2.n88 VSUBS 1.01608f
C301 VDD2.n89 VSUBS 0.029984f
C302 VDD2.n90 VSUBS 0.028611f
C303 VDD2.n91 VSUBS 0.015374f
C304 VDD2.n92 VSUBS 0.036339f
C305 VDD2.n93 VSUBS 0.016279f
C306 VDD2.n94 VSUBS 0.028611f
C307 VDD2.n95 VSUBS 0.015826f
C308 VDD2.n96 VSUBS 0.036339f
C309 VDD2.n97 VSUBS 0.015374f
C310 VDD2.n98 VSUBS 0.016279f
C311 VDD2.n99 VSUBS 0.028611f
C312 VDD2.n100 VSUBS 0.015374f
C313 VDD2.n101 VSUBS 0.036339f
C314 VDD2.n102 VSUBS 0.016279f
C315 VDD2.n103 VSUBS 0.028611f
C316 VDD2.n104 VSUBS 0.015374f
C317 VDD2.n105 VSUBS 0.036339f
C318 VDD2.n106 VSUBS 0.016279f
C319 VDD2.n107 VSUBS 0.028611f
C320 VDD2.n108 VSUBS 0.015374f
C321 VDD2.n109 VSUBS 0.036339f
C322 VDD2.n110 VSUBS 0.016279f
C323 VDD2.n111 VSUBS 0.028611f
C324 VDD2.n112 VSUBS 0.015374f
C325 VDD2.n113 VSUBS 0.036339f
C326 VDD2.n114 VSUBS 0.016279f
C327 VDD2.n115 VSUBS 0.028611f
C328 VDD2.n116 VSUBS 0.015374f
C329 VDD2.n117 VSUBS 0.027254f
C330 VDD2.n118 VSUBS 0.023117f
C331 VDD2.t1 VSUBS 0.077873f
C332 VDD2.n119 VSUBS 0.210882f
C333 VDD2.n120 VSUBS 1.96845f
C334 VDD2.n121 VSUBS 0.015374f
C335 VDD2.n122 VSUBS 0.016279f
C336 VDD2.n123 VSUBS 0.036339f
C337 VDD2.n124 VSUBS 0.036339f
C338 VDD2.n125 VSUBS 0.016279f
C339 VDD2.n126 VSUBS 0.015374f
C340 VDD2.n127 VSUBS 0.028611f
C341 VDD2.n128 VSUBS 0.028611f
C342 VDD2.n129 VSUBS 0.015374f
C343 VDD2.n130 VSUBS 0.016279f
C344 VDD2.n131 VSUBS 0.036339f
C345 VDD2.n132 VSUBS 0.036339f
C346 VDD2.n133 VSUBS 0.016279f
C347 VDD2.n134 VSUBS 0.015374f
C348 VDD2.n135 VSUBS 0.028611f
C349 VDD2.n136 VSUBS 0.028611f
C350 VDD2.n137 VSUBS 0.015374f
C351 VDD2.n138 VSUBS 0.016279f
C352 VDD2.n139 VSUBS 0.036339f
C353 VDD2.n140 VSUBS 0.036339f
C354 VDD2.n141 VSUBS 0.016279f
C355 VDD2.n142 VSUBS 0.015374f
C356 VDD2.n143 VSUBS 0.028611f
C357 VDD2.n144 VSUBS 0.028611f
C358 VDD2.n145 VSUBS 0.015374f
C359 VDD2.n146 VSUBS 0.016279f
C360 VDD2.n147 VSUBS 0.036339f
C361 VDD2.n148 VSUBS 0.036339f
C362 VDD2.n149 VSUBS 0.016279f
C363 VDD2.n150 VSUBS 0.015374f
C364 VDD2.n151 VSUBS 0.028611f
C365 VDD2.n152 VSUBS 0.028611f
C366 VDD2.n153 VSUBS 0.015374f
C367 VDD2.n154 VSUBS 0.016279f
C368 VDD2.n155 VSUBS 0.036339f
C369 VDD2.n156 VSUBS 0.036339f
C370 VDD2.n157 VSUBS 0.016279f
C371 VDD2.n158 VSUBS 0.015374f
C372 VDD2.n159 VSUBS 0.028611f
C373 VDD2.n160 VSUBS 0.028611f
C374 VDD2.n161 VSUBS 0.015374f
C375 VDD2.n162 VSUBS 0.016279f
C376 VDD2.n163 VSUBS 0.036339f
C377 VDD2.n164 VSUBS 0.036339f
C378 VDD2.n165 VSUBS 0.036339f
C379 VDD2.n166 VSUBS 0.015826f
C380 VDD2.n167 VSUBS 0.015374f
C381 VDD2.n168 VSUBS 0.028611f
C382 VDD2.n169 VSUBS 0.028611f
C383 VDD2.n170 VSUBS 0.015374f
C384 VDD2.n171 VSUBS 0.016279f
C385 VDD2.n172 VSUBS 0.036339f
C386 VDD2.n173 VSUBS 0.083022f
C387 VDD2.n174 VSUBS 0.016279f
C388 VDD2.n175 VSUBS 0.015374f
C389 VDD2.n176 VSUBS 0.066524f
C390 VDD2.n177 VSUBS 0.061295f
C391 VDD2.n178 VSUBS 3.99383f
C392 VTAIL.n0 VSUBS 0.029969f
C393 VTAIL.n1 VSUBS 0.028597f
C394 VTAIL.n2 VSUBS 0.015367f
C395 VTAIL.n3 VSUBS 0.036322f
C396 VTAIL.n4 VSUBS 0.016271f
C397 VTAIL.n5 VSUBS 0.028597f
C398 VTAIL.n6 VSUBS 0.015819f
C399 VTAIL.n7 VSUBS 0.036322f
C400 VTAIL.n8 VSUBS 0.016271f
C401 VTAIL.n9 VSUBS 0.028597f
C402 VTAIL.n10 VSUBS 0.015367f
C403 VTAIL.n11 VSUBS 0.036322f
C404 VTAIL.n12 VSUBS 0.016271f
C405 VTAIL.n13 VSUBS 0.028597f
C406 VTAIL.n14 VSUBS 0.015367f
C407 VTAIL.n15 VSUBS 0.036322f
C408 VTAIL.n16 VSUBS 0.016271f
C409 VTAIL.n17 VSUBS 0.028597f
C410 VTAIL.n18 VSUBS 0.015367f
C411 VTAIL.n19 VSUBS 0.036322f
C412 VTAIL.n20 VSUBS 0.016271f
C413 VTAIL.n21 VSUBS 0.028597f
C414 VTAIL.n22 VSUBS 0.015367f
C415 VTAIL.n23 VSUBS 0.036322f
C416 VTAIL.n24 VSUBS 0.016271f
C417 VTAIL.n25 VSUBS 0.028597f
C418 VTAIL.n26 VSUBS 0.015367f
C419 VTAIL.n27 VSUBS 0.027241f
C420 VTAIL.n28 VSUBS 0.023106f
C421 VTAIL.t0 VSUBS 0.077835f
C422 VTAIL.n29 VSUBS 0.210779f
C423 VTAIL.n30 VSUBS 1.96749f
C424 VTAIL.n31 VSUBS 0.015367f
C425 VTAIL.n32 VSUBS 0.016271f
C426 VTAIL.n33 VSUBS 0.036322f
C427 VTAIL.n34 VSUBS 0.036322f
C428 VTAIL.n35 VSUBS 0.016271f
C429 VTAIL.n36 VSUBS 0.015367f
C430 VTAIL.n37 VSUBS 0.028597f
C431 VTAIL.n38 VSUBS 0.028597f
C432 VTAIL.n39 VSUBS 0.015367f
C433 VTAIL.n40 VSUBS 0.016271f
C434 VTAIL.n41 VSUBS 0.036322f
C435 VTAIL.n42 VSUBS 0.036322f
C436 VTAIL.n43 VSUBS 0.016271f
C437 VTAIL.n44 VSUBS 0.015367f
C438 VTAIL.n45 VSUBS 0.028597f
C439 VTAIL.n46 VSUBS 0.028597f
C440 VTAIL.n47 VSUBS 0.015367f
C441 VTAIL.n48 VSUBS 0.016271f
C442 VTAIL.n49 VSUBS 0.036322f
C443 VTAIL.n50 VSUBS 0.036322f
C444 VTAIL.n51 VSUBS 0.016271f
C445 VTAIL.n52 VSUBS 0.015367f
C446 VTAIL.n53 VSUBS 0.028597f
C447 VTAIL.n54 VSUBS 0.028597f
C448 VTAIL.n55 VSUBS 0.015367f
C449 VTAIL.n56 VSUBS 0.016271f
C450 VTAIL.n57 VSUBS 0.036322f
C451 VTAIL.n58 VSUBS 0.036322f
C452 VTAIL.n59 VSUBS 0.016271f
C453 VTAIL.n60 VSUBS 0.015367f
C454 VTAIL.n61 VSUBS 0.028597f
C455 VTAIL.n62 VSUBS 0.028597f
C456 VTAIL.n63 VSUBS 0.015367f
C457 VTAIL.n64 VSUBS 0.016271f
C458 VTAIL.n65 VSUBS 0.036322f
C459 VTAIL.n66 VSUBS 0.036322f
C460 VTAIL.n67 VSUBS 0.016271f
C461 VTAIL.n68 VSUBS 0.015367f
C462 VTAIL.n69 VSUBS 0.028597f
C463 VTAIL.n70 VSUBS 0.028597f
C464 VTAIL.n71 VSUBS 0.015367f
C465 VTAIL.n72 VSUBS 0.015367f
C466 VTAIL.n73 VSUBS 0.016271f
C467 VTAIL.n74 VSUBS 0.036322f
C468 VTAIL.n75 VSUBS 0.036322f
C469 VTAIL.n76 VSUBS 0.036322f
C470 VTAIL.n77 VSUBS 0.015819f
C471 VTAIL.n78 VSUBS 0.015367f
C472 VTAIL.n79 VSUBS 0.028597f
C473 VTAIL.n80 VSUBS 0.028597f
C474 VTAIL.n81 VSUBS 0.015367f
C475 VTAIL.n82 VSUBS 0.016271f
C476 VTAIL.n83 VSUBS 0.036322f
C477 VTAIL.n84 VSUBS 0.082981f
C478 VTAIL.n85 VSUBS 0.016271f
C479 VTAIL.n86 VSUBS 0.015367f
C480 VTAIL.n87 VSUBS 0.066492f
C481 VTAIL.n88 VSUBS 0.041523f
C482 VTAIL.n89 VSUBS 2.27966f
C483 VTAIL.n90 VSUBS 0.029969f
C484 VTAIL.n91 VSUBS 0.028597f
C485 VTAIL.n92 VSUBS 0.015367f
C486 VTAIL.n93 VSUBS 0.036322f
C487 VTAIL.n94 VSUBS 0.016271f
C488 VTAIL.n95 VSUBS 0.028597f
C489 VTAIL.n96 VSUBS 0.015819f
C490 VTAIL.n97 VSUBS 0.036322f
C491 VTAIL.n98 VSUBS 0.015367f
C492 VTAIL.n99 VSUBS 0.016271f
C493 VTAIL.n100 VSUBS 0.028597f
C494 VTAIL.n101 VSUBS 0.015367f
C495 VTAIL.n102 VSUBS 0.036322f
C496 VTAIL.n103 VSUBS 0.016271f
C497 VTAIL.n104 VSUBS 0.028597f
C498 VTAIL.n105 VSUBS 0.015367f
C499 VTAIL.n106 VSUBS 0.036322f
C500 VTAIL.n107 VSUBS 0.016271f
C501 VTAIL.n108 VSUBS 0.028597f
C502 VTAIL.n109 VSUBS 0.015367f
C503 VTAIL.n110 VSUBS 0.036322f
C504 VTAIL.n111 VSUBS 0.016271f
C505 VTAIL.n112 VSUBS 0.028597f
C506 VTAIL.n113 VSUBS 0.015367f
C507 VTAIL.n114 VSUBS 0.036322f
C508 VTAIL.n115 VSUBS 0.016271f
C509 VTAIL.n116 VSUBS 0.028597f
C510 VTAIL.n117 VSUBS 0.015367f
C511 VTAIL.n118 VSUBS 0.027241f
C512 VTAIL.n119 VSUBS 0.023106f
C513 VTAIL.t3 VSUBS 0.077835f
C514 VTAIL.n120 VSUBS 0.210779f
C515 VTAIL.n121 VSUBS 1.96749f
C516 VTAIL.n122 VSUBS 0.015367f
C517 VTAIL.n123 VSUBS 0.016271f
C518 VTAIL.n124 VSUBS 0.036322f
C519 VTAIL.n125 VSUBS 0.036322f
C520 VTAIL.n126 VSUBS 0.016271f
C521 VTAIL.n127 VSUBS 0.015367f
C522 VTAIL.n128 VSUBS 0.028597f
C523 VTAIL.n129 VSUBS 0.028597f
C524 VTAIL.n130 VSUBS 0.015367f
C525 VTAIL.n131 VSUBS 0.016271f
C526 VTAIL.n132 VSUBS 0.036322f
C527 VTAIL.n133 VSUBS 0.036322f
C528 VTAIL.n134 VSUBS 0.016271f
C529 VTAIL.n135 VSUBS 0.015367f
C530 VTAIL.n136 VSUBS 0.028597f
C531 VTAIL.n137 VSUBS 0.028597f
C532 VTAIL.n138 VSUBS 0.015367f
C533 VTAIL.n139 VSUBS 0.016271f
C534 VTAIL.n140 VSUBS 0.036322f
C535 VTAIL.n141 VSUBS 0.036322f
C536 VTAIL.n142 VSUBS 0.016271f
C537 VTAIL.n143 VSUBS 0.015367f
C538 VTAIL.n144 VSUBS 0.028597f
C539 VTAIL.n145 VSUBS 0.028597f
C540 VTAIL.n146 VSUBS 0.015367f
C541 VTAIL.n147 VSUBS 0.016271f
C542 VTAIL.n148 VSUBS 0.036322f
C543 VTAIL.n149 VSUBS 0.036322f
C544 VTAIL.n150 VSUBS 0.016271f
C545 VTAIL.n151 VSUBS 0.015367f
C546 VTAIL.n152 VSUBS 0.028597f
C547 VTAIL.n153 VSUBS 0.028597f
C548 VTAIL.n154 VSUBS 0.015367f
C549 VTAIL.n155 VSUBS 0.016271f
C550 VTAIL.n156 VSUBS 0.036322f
C551 VTAIL.n157 VSUBS 0.036322f
C552 VTAIL.n158 VSUBS 0.016271f
C553 VTAIL.n159 VSUBS 0.015367f
C554 VTAIL.n160 VSUBS 0.028597f
C555 VTAIL.n161 VSUBS 0.028597f
C556 VTAIL.n162 VSUBS 0.015367f
C557 VTAIL.n163 VSUBS 0.016271f
C558 VTAIL.n164 VSUBS 0.036322f
C559 VTAIL.n165 VSUBS 0.036322f
C560 VTAIL.n166 VSUBS 0.036322f
C561 VTAIL.n167 VSUBS 0.015819f
C562 VTAIL.n168 VSUBS 0.015367f
C563 VTAIL.n169 VSUBS 0.028597f
C564 VTAIL.n170 VSUBS 0.028597f
C565 VTAIL.n171 VSUBS 0.015367f
C566 VTAIL.n172 VSUBS 0.016271f
C567 VTAIL.n173 VSUBS 0.036322f
C568 VTAIL.n174 VSUBS 0.082981f
C569 VTAIL.n175 VSUBS 0.016271f
C570 VTAIL.n176 VSUBS 0.015367f
C571 VTAIL.n177 VSUBS 0.066492f
C572 VTAIL.n178 VSUBS 0.041523f
C573 VTAIL.n179 VSUBS 2.33427f
C574 VTAIL.n180 VSUBS 0.029969f
C575 VTAIL.n181 VSUBS 0.028597f
C576 VTAIL.n182 VSUBS 0.015367f
C577 VTAIL.n183 VSUBS 0.036322f
C578 VTAIL.n184 VSUBS 0.016271f
C579 VTAIL.n185 VSUBS 0.028597f
C580 VTAIL.n186 VSUBS 0.015819f
C581 VTAIL.n187 VSUBS 0.036322f
C582 VTAIL.n188 VSUBS 0.015367f
C583 VTAIL.n189 VSUBS 0.016271f
C584 VTAIL.n190 VSUBS 0.028597f
C585 VTAIL.n191 VSUBS 0.015367f
C586 VTAIL.n192 VSUBS 0.036322f
C587 VTAIL.n193 VSUBS 0.016271f
C588 VTAIL.n194 VSUBS 0.028597f
C589 VTAIL.n195 VSUBS 0.015367f
C590 VTAIL.n196 VSUBS 0.036322f
C591 VTAIL.n197 VSUBS 0.016271f
C592 VTAIL.n198 VSUBS 0.028597f
C593 VTAIL.n199 VSUBS 0.015367f
C594 VTAIL.n200 VSUBS 0.036322f
C595 VTAIL.n201 VSUBS 0.016271f
C596 VTAIL.n202 VSUBS 0.028597f
C597 VTAIL.n203 VSUBS 0.015367f
C598 VTAIL.n204 VSUBS 0.036322f
C599 VTAIL.n205 VSUBS 0.016271f
C600 VTAIL.n206 VSUBS 0.028597f
C601 VTAIL.n207 VSUBS 0.015367f
C602 VTAIL.n208 VSUBS 0.027241f
C603 VTAIL.n209 VSUBS 0.023106f
C604 VTAIL.t1 VSUBS 0.077835f
C605 VTAIL.n210 VSUBS 0.210779f
C606 VTAIL.n211 VSUBS 1.96749f
C607 VTAIL.n212 VSUBS 0.015367f
C608 VTAIL.n213 VSUBS 0.016271f
C609 VTAIL.n214 VSUBS 0.036322f
C610 VTAIL.n215 VSUBS 0.036322f
C611 VTAIL.n216 VSUBS 0.016271f
C612 VTAIL.n217 VSUBS 0.015367f
C613 VTAIL.n218 VSUBS 0.028597f
C614 VTAIL.n219 VSUBS 0.028597f
C615 VTAIL.n220 VSUBS 0.015367f
C616 VTAIL.n221 VSUBS 0.016271f
C617 VTAIL.n222 VSUBS 0.036322f
C618 VTAIL.n223 VSUBS 0.036322f
C619 VTAIL.n224 VSUBS 0.016271f
C620 VTAIL.n225 VSUBS 0.015367f
C621 VTAIL.n226 VSUBS 0.028597f
C622 VTAIL.n227 VSUBS 0.028597f
C623 VTAIL.n228 VSUBS 0.015367f
C624 VTAIL.n229 VSUBS 0.016271f
C625 VTAIL.n230 VSUBS 0.036322f
C626 VTAIL.n231 VSUBS 0.036322f
C627 VTAIL.n232 VSUBS 0.016271f
C628 VTAIL.n233 VSUBS 0.015367f
C629 VTAIL.n234 VSUBS 0.028597f
C630 VTAIL.n235 VSUBS 0.028597f
C631 VTAIL.n236 VSUBS 0.015367f
C632 VTAIL.n237 VSUBS 0.016271f
C633 VTAIL.n238 VSUBS 0.036322f
C634 VTAIL.n239 VSUBS 0.036322f
C635 VTAIL.n240 VSUBS 0.016271f
C636 VTAIL.n241 VSUBS 0.015367f
C637 VTAIL.n242 VSUBS 0.028597f
C638 VTAIL.n243 VSUBS 0.028597f
C639 VTAIL.n244 VSUBS 0.015367f
C640 VTAIL.n245 VSUBS 0.016271f
C641 VTAIL.n246 VSUBS 0.036322f
C642 VTAIL.n247 VSUBS 0.036322f
C643 VTAIL.n248 VSUBS 0.016271f
C644 VTAIL.n249 VSUBS 0.015367f
C645 VTAIL.n250 VSUBS 0.028597f
C646 VTAIL.n251 VSUBS 0.028597f
C647 VTAIL.n252 VSUBS 0.015367f
C648 VTAIL.n253 VSUBS 0.016271f
C649 VTAIL.n254 VSUBS 0.036322f
C650 VTAIL.n255 VSUBS 0.036322f
C651 VTAIL.n256 VSUBS 0.036322f
C652 VTAIL.n257 VSUBS 0.015819f
C653 VTAIL.n258 VSUBS 0.015367f
C654 VTAIL.n259 VSUBS 0.028597f
C655 VTAIL.n260 VSUBS 0.028597f
C656 VTAIL.n261 VSUBS 0.015367f
C657 VTAIL.n262 VSUBS 0.016271f
C658 VTAIL.n263 VSUBS 0.036322f
C659 VTAIL.n264 VSUBS 0.082981f
C660 VTAIL.n265 VSUBS 0.016271f
C661 VTAIL.n266 VSUBS 0.015367f
C662 VTAIL.n267 VSUBS 0.066492f
C663 VTAIL.n268 VSUBS 0.041523f
C664 VTAIL.n269 VSUBS 2.09437f
C665 VTAIL.n270 VSUBS 0.029969f
C666 VTAIL.n271 VSUBS 0.028597f
C667 VTAIL.n272 VSUBS 0.015367f
C668 VTAIL.n273 VSUBS 0.036322f
C669 VTAIL.n274 VSUBS 0.016271f
C670 VTAIL.n275 VSUBS 0.028597f
C671 VTAIL.n276 VSUBS 0.015819f
C672 VTAIL.n277 VSUBS 0.036322f
C673 VTAIL.n278 VSUBS 0.016271f
C674 VTAIL.n279 VSUBS 0.028597f
C675 VTAIL.n280 VSUBS 0.015367f
C676 VTAIL.n281 VSUBS 0.036322f
C677 VTAIL.n282 VSUBS 0.016271f
C678 VTAIL.n283 VSUBS 0.028597f
C679 VTAIL.n284 VSUBS 0.015367f
C680 VTAIL.n285 VSUBS 0.036322f
C681 VTAIL.n286 VSUBS 0.016271f
C682 VTAIL.n287 VSUBS 0.028597f
C683 VTAIL.n288 VSUBS 0.015367f
C684 VTAIL.n289 VSUBS 0.036322f
C685 VTAIL.n290 VSUBS 0.016271f
C686 VTAIL.n291 VSUBS 0.028597f
C687 VTAIL.n292 VSUBS 0.015367f
C688 VTAIL.n293 VSUBS 0.036322f
C689 VTAIL.n294 VSUBS 0.016271f
C690 VTAIL.n295 VSUBS 0.028597f
C691 VTAIL.n296 VSUBS 0.015367f
C692 VTAIL.n297 VSUBS 0.027241f
C693 VTAIL.n298 VSUBS 0.023106f
C694 VTAIL.t2 VSUBS 0.077835f
C695 VTAIL.n299 VSUBS 0.210779f
C696 VTAIL.n300 VSUBS 1.96749f
C697 VTAIL.n301 VSUBS 0.015367f
C698 VTAIL.n302 VSUBS 0.016271f
C699 VTAIL.n303 VSUBS 0.036322f
C700 VTAIL.n304 VSUBS 0.036322f
C701 VTAIL.n305 VSUBS 0.016271f
C702 VTAIL.n306 VSUBS 0.015367f
C703 VTAIL.n307 VSUBS 0.028597f
C704 VTAIL.n308 VSUBS 0.028597f
C705 VTAIL.n309 VSUBS 0.015367f
C706 VTAIL.n310 VSUBS 0.016271f
C707 VTAIL.n311 VSUBS 0.036322f
C708 VTAIL.n312 VSUBS 0.036322f
C709 VTAIL.n313 VSUBS 0.016271f
C710 VTAIL.n314 VSUBS 0.015367f
C711 VTAIL.n315 VSUBS 0.028597f
C712 VTAIL.n316 VSUBS 0.028597f
C713 VTAIL.n317 VSUBS 0.015367f
C714 VTAIL.n318 VSUBS 0.016271f
C715 VTAIL.n319 VSUBS 0.036322f
C716 VTAIL.n320 VSUBS 0.036322f
C717 VTAIL.n321 VSUBS 0.016271f
C718 VTAIL.n322 VSUBS 0.015367f
C719 VTAIL.n323 VSUBS 0.028597f
C720 VTAIL.n324 VSUBS 0.028597f
C721 VTAIL.n325 VSUBS 0.015367f
C722 VTAIL.n326 VSUBS 0.016271f
C723 VTAIL.n327 VSUBS 0.036322f
C724 VTAIL.n328 VSUBS 0.036322f
C725 VTAIL.n329 VSUBS 0.016271f
C726 VTAIL.n330 VSUBS 0.015367f
C727 VTAIL.n331 VSUBS 0.028597f
C728 VTAIL.n332 VSUBS 0.028597f
C729 VTAIL.n333 VSUBS 0.015367f
C730 VTAIL.n334 VSUBS 0.016271f
C731 VTAIL.n335 VSUBS 0.036322f
C732 VTAIL.n336 VSUBS 0.036322f
C733 VTAIL.n337 VSUBS 0.016271f
C734 VTAIL.n338 VSUBS 0.015367f
C735 VTAIL.n339 VSUBS 0.028597f
C736 VTAIL.n340 VSUBS 0.028597f
C737 VTAIL.n341 VSUBS 0.015367f
C738 VTAIL.n342 VSUBS 0.015367f
C739 VTAIL.n343 VSUBS 0.016271f
C740 VTAIL.n344 VSUBS 0.036322f
C741 VTAIL.n345 VSUBS 0.036322f
C742 VTAIL.n346 VSUBS 0.036322f
C743 VTAIL.n347 VSUBS 0.015819f
C744 VTAIL.n348 VSUBS 0.015367f
C745 VTAIL.n349 VSUBS 0.028597f
C746 VTAIL.n350 VSUBS 0.028597f
C747 VTAIL.n351 VSUBS 0.015367f
C748 VTAIL.n352 VSUBS 0.016271f
C749 VTAIL.n353 VSUBS 0.036322f
C750 VTAIL.n354 VSUBS 0.082981f
C751 VTAIL.n355 VSUBS 0.016271f
C752 VTAIL.n356 VSUBS 0.015367f
C753 VTAIL.n357 VSUBS 0.066492f
C754 VTAIL.n358 VSUBS 0.041523f
C755 VTAIL.n359 VSUBS 1.98574f
C756 VN.t1 VSUBS 4.708509f
C757 VN.t0 VSUBS 5.40752f
C758 B.n0 VSUBS 0.004468f
C759 B.n1 VSUBS 0.004468f
C760 B.n2 VSUBS 0.007065f
C761 B.n3 VSUBS 0.007065f
C762 B.n4 VSUBS 0.007065f
C763 B.n5 VSUBS 0.007065f
C764 B.n6 VSUBS 0.007065f
C765 B.n7 VSUBS 0.007065f
C766 B.n8 VSUBS 0.007065f
C767 B.n9 VSUBS 0.007065f
C768 B.n10 VSUBS 0.007065f
C769 B.n11 VSUBS 0.007065f
C770 B.n12 VSUBS 0.007065f
C771 B.n13 VSUBS 0.007065f
C772 B.n14 VSUBS 0.007065f
C773 B.n15 VSUBS 0.016175f
C774 B.n16 VSUBS 0.007065f
C775 B.n17 VSUBS 0.007065f
C776 B.n18 VSUBS 0.007065f
C777 B.n19 VSUBS 0.007065f
C778 B.n20 VSUBS 0.007065f
C779 B.n21 VSUBS 0.007065f
C780 B.n22 VSUBS 0.007065f
C781 B.n23 VSUBS 0.007065f
C782 B.n24 VSUBS 0.007065f
C783 B.n25 VSUBS 0.007065f
C784 B.n26 VSUBS 0.007065f
C785 B.n27 VSUBS 0.007065f
C786 B.n28 VSUBS 0.007065f
C787 B.n29 VSUBS 0.007065f
C788 B.n30 VSUBS 0.007065f
C789 B.n31 VSUBS 0.007065f
C790 B.n32 VSUBS 0.007065f
C791 B.n33 VSUBS 0.007065f
C792 B.n34 VSUBS 0.007065f
C793 B.n35 VSUBS 0.007065f
C794 B.n36 VSUBS 0.007065f
C795 B.n37 VSUBS 0.007065f
C796 B.n38 VSUBS 0.007065f
C797 B.n39 VSUBS 0.007065f
C798 B.n40 VSUBS 0.007065f
C799 B.n41 VSUBS 0.007065f
C800 B.t11 VSUBS 0.308061f
C801 B.t10 VSUBS 0.34251f
C802 B.t9 VSUBS 1.95736f
C803 B.n42 VSUBS 0.531312f
C804 B.n43 VSUBS 0.308743f
C805 B.n44 VSUBS 0.016369f
C806 B.n45 VSUBS 0.007065f
C807 B.n46 VSUBS 0.007065f
C808 B.n47 VSUBS 0.007065f
C809 B.n48 VSUBS 0.007065f
C810 B.n49 VSUBS 0.007065f
C811 B.t8 VSUBS 0.308064f
C812 B.t7 VSUBS 0.342513f
C813 B.t6 VSUBS 1.95736f
C814 B.n50 VSUBS 0.531309f
C815 B.n51 VSUBS 0.308739f
C816 B.n52 VSUBS 0.007065f
C817 B.n53 VSUBS 0.007065f
C818 B.n54 VSUBS 0.007065f
C819 B.n55 VSUBS 0.007065f
C820 B.n56 VSUBS 0.007065f
C821 B.n57 VSUBS 0.007065f
C822 B.n58 VSUBS 0.007065f
C823 B.n59 VSUBS 0.007065f
C824 B.n60 VSUBS 0.007065f
C825 B.n61 VSUBS 0.007065f
C826 B.n62 VSUBS 0.007065f
C827 B.n63 VSUBS 0.007065f
C828 B.n64 VSUBS 0.007065f
C829 B.n65 VSUBS 0.007065f
C830 B.n66 VSUBS 0.007065f
C831 B.n67 VSUBS 0.007065f
C832 B.n68 VSUBS 0.007065f
C833 B.n69 VSUBS 0.007065f
C834 B.n70 VSUBS 0.007065f
C835 B.n71 VSUBS 0.007065f
C836 B.n72 VSUBS 0.007065f
C837 B.n73 VSUBS 0.007065f
C838 B.n74 VSUBS 0.007065f
C839 B.n75 VSUBS 0.007065f
C840 B.n76 VSUBS 0.007065f
C841 B.n77 VSUBS 0.007065f
C842 B.n78 VSUBS 0.016306f
C843 B.n79 VSUBS 0.007065f
C844 B.n80 VSUBS 0.007065f
C845 B.n81 VSUBS 0.007065f
C846 B.n82 VSUBS 0.007065f
C847 B.n83 VSUBS 0.007065f
C848 B.n84 VSUBS 0.007065f
C849 B.n85 VSUBS 0.007065f
C850 B.n86 VSUBS 0.007065f
C851 B.n87 VSUBS 0.007065f
C852 B.n88 VSUBS 0.007065f
C853 B.n89 VSUBS 0.007065f
C854 B.n90 VSUBS 0.007065f
C855 B.n91 VSUBS 0.007065f
C856 B.n92 VSUBS 0.007065f
C857 B.n93 VSUBS 0.007065f
C858 B.n94 VSUBS 0.007065f
C859 B.n95 VSUBS 0.007065f
C860 B.n96 VSUBS 0.007065f
C861 B.n97 VSUBS 0.007065f
C862 B.n98 VSUBS 0.007065f
C863 B.n99 VSUBS 0.007065f
C864 B.n100 VSUBS 0.007065f
C865 B.n101 VSUBS 0.007065f
C866 B.n102 VSUBS 0.007065f
C867 B.n103 VSUBS 0.007065f
C868 B.n104 VSUBS 0.015411f
C869 B.n105 VSUBS 0.007065f
C870 B.n106 VSUBS 0.007065f
C871 B.n107 VSUBS 0.007065f
C872 B.n108 VSUBS 0.007065f
C873 B.n109 VSUBS 0.007065f
C874 B.n110 VSUBS 0.007065f
C875 B.n111 VSUBS 0.007065f
C876 B.n112 VSUBS 0.007065f
C877 B.n113 VSUBS 0.007065f
C878 B.n114 VSUBS 0.007065f
C879 B.n115 VSUBS 0.007065f
C880 B.n116 VSUBS 0.007065f
C881 B.n117 VSUBS 0.007065f
C882 B.n118 VSUBS 0.007065f
C883 B.n119 VSUBS 0.007065f
C884 B.n120 VSUBS 0.007065f
C885 B.n121 VSUBS 0.007065f
C886 B.n122 VSUBS 0.007065f
C887 B.n123 VSUBS 0.007065f
C888 B.n124 VSUBS 0.007065f
C889 B.n125 VSUBS 0.007065f
C890 B.n126 VSUBS 0.007065f
C891 B.n127 VSUBS 0.007065f
C892 B.n128 VSUBS 0.007065f
C893 B.n129 VSUBS 0.007065f
C894 B.n130 VSUBS 0.007065f
C895 B.n131 VSUBS 0.007065f
C896 B.t1 VSUBS 0.308064f
C897 B.t2 VSUBS 0.342513f
C898 B.t0 VSUBS 1.95736f
C899 B.n132 VSUBS 0.531309f
C900 B.n133 VSUBS 0.308739f
C901 B.n134 VSUBS 0.007065f
C902 B.n135 VSUBS 0.007065f
C903 B.n136 VSUBS 0.007065f
C904 B.n137 VSUBS 0.007065f
C905 B.t4 VSUBS 0.308061f
C906 B.t5 VSUBS 0.34251f
C907 B.t3 VSUBS 1.95736f
C908 B.n138 VSUBS 0.531312f
C909 B.n139 VSUBS 0.308743f
C910 B.n140 VSUBS 0.016369f
C911 B.n141 VSUBS 0.007065f
C912 B.n142 VSUBS 0.007065f
C913 B.n143 VSUBS 0.007065f
C914 B.n144 VSUBS 0.007065f
C915 B.n145 VSUBS 0.007065f
C916 B.n146 VSUBS 0.007065f
C917 B.n147 VSUBS 0.007065f
C918 B.n148 VSUBS 0.007065f
C919 B.n149 VSUBS 0.007065f
C920 B.n150 VSUBS 0.007065f
C921 B.n151 VSUBS 0.007065f
C922 B.n152 VSUBS 0.007065f
C923 B.n153 VSUBS 0.007065f
C924 B.n154 VSUBS 0.007065f
C925 B.n155 VSUBS 0.007065f
C926 B.n156 VSUBS 0.007065f
C927 B.n157 VSUBS 0.007065f
C928 B.n158 VSUBS 0.007065f
C929 B.n159 VSUBS 0.007065f
C930 B.n160 VSUBS 0.007065f
C931 B.n161 VSUBS 0.007065f
C932 B.n162 VSUBS 0.007065f
C933 B.n163 VSUBS 0.007065f
C934 B.n164 VSUBS 0.007065f
C935 B.n165 VSUBS 0.007065f
C936 B.n166 VSUBS 0.007065f
C937 B.n167 VSUBS 0.016175f
C938 B.n168 VSUBS 0.007065f
C939 B.n169 VSUBS 0.007065f
C940 B.n170 VSUBS 0.007065f
C941 B.n171 VSUBS 0.007065f
C942 B.n172 VSUBS 0.007065f
C943 B.n173 VSUBS 0.007065f
C944 B.n174 VSUBS 0.007065f
C945 B.n175 VSUBS 0.007065f
C946 B.n176 VSUBS 0.007065f
C947 B.n177 VSUBS 0.007065f
C948 B.n178 VSUBS 0.007065f
C949 B.n179 VSUBS 0.007065f
C950 B.n180 VSUBS 0.007065f
C951 B.n181 VSUBS 0.007065f
C952 B.n182 VSUBS 0.007065f
C953 B.n183 VSUBS 0.007065f
C954 B.n184 VSUBS 0.007065f
C955 B.n185 VSUBS 0.007065f
C956 B.n186 VSUBS 0.007065f
C957 B.n187 VSUBS 0.007065f
C958 B.n188 VSUBS 0.007065f
C959 B.n189 VSUBS 0.007065f
C960 B.n190 VSUBS 0.007065f
C961 B.n191 VSUBS 0.007065f
C962 B.n192 VSUBS 0.007065f
C963 B.n193 VSUBS 0.007065f
C964 B.n194 VSUBS 0.007065f
C965 B.n195 VSUBS 0.007065f
C966 B.n196 VSUBS 0.007065f
C967 B.n197 VSUBS 0.007065f
C968 B.n198 VSUBS 0.007065f
C969 B.n199 VSUBS 0.007065f
C970 B.n200 VSUBS 0.007065f
C971 B.n201 VSUBS 0.007065f
C972 B.n202 VSUBS 0.007065f
C973 B.n203 VSUBS 0.007065f
C974 B.n204 VSUBS 0.007065f
C975 B.n205 VSUBS 0.007065f
C976 B.n206 VSUBS 0.007065f
C977 B.n207 VSUBS 0.007065f
C978 B.n208 VSUBS 0.007065f
C979 B.n209 VSUBS 0.007065f
C980 B.n210 VSUBS 0.007065f
C981 B.n211 VSUBS 0.007065f
C982 B.n212 VSUBS 0.007065f
C983 B.n213 VSUBS 0.007065f
C984 B.n214 VSUBS 0.007065f
C985 B.n215 VSUBS 0.007065f
C986 B.n216 VSUBS 0.015411f
C987 B.n217 VSUBS 0.015411f
C988 B.n218 VSUBS 0.016175f
C989 B.n219 VSUBS 0.007065f
C990 B.n220 VSUBS 0.007065f
C991 B.n221 VSUBS 0.007065f
C992 B.n222 VSUBS 0.007065f
C993 B.n223 VSUBS 0.007065f
C994 B.n224 VSUBS 0.007065f
C995 B.n225 VSUBS 0.007065f
C996 B.n226 VSUBS 0.007065f
C997 B.n227 VSUBS 0.007065f
C998 B.n228 VSUBS 0.007065f
C999 B.n229 VSUBS 0.007065f
C1000 B.n230 VSUBS 0.007065f
C1001 B.n231 VSUBS 0.007065f
C1002 B.n232 VSUBS 0.007065f
C1003 B.n233 VSUBS 0.007065f
C1004 B.n234 VSUBS 0.007065f
C1005 B.n235 VSUBS 0.007065f
C1006 B.n236 VSUBS 0.007065f
C1007 B.n237 VSUBS 0.007065f
C1008 B.n238 VSUBS 0.007065f
C1009 B.n239 VSUBS 0.007065f
C1010 B.n240 VSUBS 0.007065f
C1011 B.n241 VSUBS 0.007065f
C1012 B.n242 VSUBS 0.007065f
C1013 B.n243 VSUBS 0.007065f
C1014 B.n244 VSUBS 0.007065f
C1015 B.n245 VSUBS 0.007065f
C1016 B.n246 VSUBS 0.007065f
C1017 B.n247 VSUBS 0.007065f
C1018 B.n248 VSUBS 0.007065f
C1019 B.n249 VSUBS 0.007065f
C1020 B.n250 VSUBS 0.007065f
C1021 B.n251 VSUBS 0.007065f
C1022 B.n252 VSUBS 0.007065f
C1023 B.n253 VSUBS 0.007065f
C1024 B.n254 VSUBS 0.007065f
C1025 B.n255 VSUBS 0.007065f
C1026 B.n256 VSUBS 0.007065f
C1027 B.n257 VSUBS 0.007065f
C1028 B.n258 VSUBS 0.007065f
C1029 B.n259 VSUBS 0.007065f
C1030 B.n260 VSUBS 0.007065f
C1031 B.n261 VSUBS 0.007065f
C1032 B.n262 VSUBS 0.007065f
C1033 B.n263 VSUBS 0.007065f
C1034 B.n264 VSUBS 0.007065f
C1035 B.n265 VSUBS 0.007065f
C1036 B.n266 VSUBS 0.007065f
C1037 B.n267 VSUBS 0.007065f
C1038 B.n268 VSUBS 0.007065f
C1039 B.n269 VSUBS 0.007065f
C1040 B.n270 VSUBS 0.007065f
C1041 B.n271 VSUBS 0.007065f
C1042 B.n272 VSUBS 0.007065f
C1043 B.n273 VSUBS 0.007065f
C1044 B.n274 VSUBS 0.007065f
C1045 B.n275 VSUBS 0.007065f
C1046 B.n276 VSUBS 0.007065f
C1047 B.n277 VSUBS 0.007065f
C1048 B.n278 VSUBS 0.007065f
C1049 B.n279 VSUBS 0.007065f
C1050 B.n280 VSUBS 0.007065f
C1051 B.n281 VSUBS 0.007065f
C1052 B.n282 VSUBS 0.007065f
C1053 B.n283 VSUBS 0.007065f
C1054 B.n284 VSUBS 0.007065f
C1055 B.n285 VSUBS 0.007065f
C1056 B.n286 VSUBS 0.007065f
C1057 B.n287 VSUBS 0.007065f
C1058 B.n288 VSUBS 0.007065f
C1059 B.n289 VSUBS 0.007065f
C1060 B.n290 VSUBS 0.007065f
C1061 B.n291 VSUBS 0.007065f
C1062 B.n292 VSUBS 0.007065f
C1063 B.n293 VSUBS 0.007065f
C1064 B.n294 VSUBS 0.007065f
C1065 B.n295 VSUBS 0.007065f
C1066 B.n296 VSUBS 0.007065f
C1067 B.n297 VSUBS 0.004883f
C1068 B.n298 VSUBS 0.007065f
C1069 B.n299 VSUBS 0.007065f
C1070 B.n300 VSUBS 0.005715f
C1071 B.n301 VSUBS 0.007065f
C1072 B.n302 VSUBS 0.007065f
C1073 B.n303 VSUBS 0.007065f
C1074 B.n304 VSUBS 0.007065f
C1075 B.n305 VSUBS 0.007065f
C1076 B.n306 VSUBS 0.007065f
C1077 B.n307 VSUBS 0.007065f
C1078 B.n308 VSUBS 0.007065f
C1079 B.n309 VSUBS 0.007065f
C1080 B.n310 VSUBS 0.007065f
C1081 B.n311 VSUBS 0.007065f
C1082 B.n312 VSUBS 0.005715f
C1083 B.n313 VSUBS 0.016369f
C1084 B.n314 VSUBS 0.004883f
C1085 B.n315 VSUBS 0.007065f
C1086 B.n316 VSUBS 0.007065f
C1087 B.n317 VSUBS 0.007065f
C1088 B.n318 VSUBS 0.007065f
C1089 B.n319 VSUBS 0.007065f
C1090 B.n320 VSUBS 0.007065f
C1091 B.n321 VSUBS 0.007065f
C1092 B.n322 VSUBS 0.007065f
C1093 B.n323 VSUBS 0.007065f
C1094 B.n324 VSUBS 0.007065f
C1095 B.n325 VSUBS 0.007065f
C1096 B.n326 VSUBS 0.007065f
C1097 B.n327 VSUBS 0.007065f
C1098 B.n328 VSUBS 0.007065f
C1099 B.n329 VSUBS 0.007065f
C1100 B.n330 VSUBS 0.007065f
C1101 B.n331 VSUBS 0.007065f
C1102 B.n332 VSUBS 0.007065f
C1103 B.n333 VSUBS 0.007065f
C1104 B.n334 VSUBS 0.007065f
C1105 B.n335 VSUBS 0.007065f
C1106 B.n336 VSUBS 0.007065f
C1107 B.n337 VSUBS 0.007065f
C1108 B.n338 VSUBS 0.007065f
C1109 B.n339 VSUBS 0.007065f
C1110 B.n340 VSUBS 0.007065f
C1111 B.n341 VSUBS 0.007065f
C1112 B.n342 VSUBS 0.007065f
C1113 B.n343 VSUBS 0.007065f
C1114 B.n344 VSUBS 0.007065f
C1115 B.n345 VSUBS 0.007065f
C1116 B.n346 VSUBS 0.007065f
C1117 B.n347 VSUBS 0.007065f
C1118 B.n348 VSUBS 0.007065f
C1119 B.n349 VSUBS 0.007065f
C1120 B.n350 VSUBS 0.007065f
C1121 B.n351 VSUBS 0.007065f
C1122 B.n352 VSUBS 0.007065f
C1123 B.n353 VSUBS 0.007065f
C1124 B.n354 VSUBS 0.007065f
C1125 B.n355 VSUBS 0.007065f
C1126 B.n356 VSUBS 0.007065f
C1127 B.n357 VSUBS 0.007065f
C1128 B.n358 VSUBS 0.007065f
C1129 B.n359 VSUBS 0.007065f
C1130 B.n360 VSUBS 0.007065f
C1131 B.n361 VSUBS 0.007065f
C1132 B.n362 VSUBS 0.007065f
C1133 B.n363 VSUBS 0.007065f
C1134 B.n364 VSUBS 0.007065f
C1135 B.n365 VSUBS 0.007065f
C1136 B.n366 VSUBS 0.007065f
C1137 B.n367 VSUBS 0.007065f
C1138 B.n368 VSUBS 0.007065f
C1139 B.n369 VSUBS 0.007065f
C1140 B.n370 VSUBS 0.007065f
C1141 B.n371 VSUBS 0.007065f
C1142 B.n372 VSUBS 0.007065f
C1143 B.n373 VSUBS 0.007065f
C1144 B.n374 VSUBS 0.007065f
C1145 B.n375 VSUBS 0.007065f
C1146 B.n376 VSUBS 0.007065f
C1147 B.n377 VSUBS 0.007065f
C1148 B.n378 VSUBS 0.007065f
C1149 B.n379 VSUBS 0.007065f
C1150 B.n380 VSUBS 0.007065f
C1151 B.n381 VSUBS 0.007065f
C1152 B.n382 VSUBS 0.007065f
C1153 B.n383 VSUBS 0.007065f
C1154 B.n384 VSUBS 0.007065f
C1155 B.n385 VSUBS 0.007065f
C1156 B.n386 VSUBS 0.007065f
C1157 B.n387 VSUBS 0.007065f
C1158 B.n388 VSUBS 0.007065f
C1159 B.n389 VSUBS 0.007065f
C1160 B.n390 VSUBS 0.007065f
C1161 B.n391 VSUBS 0.007065f
C1162 B.n392 VSUBS 0.007065f
C1163 B.n393 VSUBS 0.016175f
C1164 B.n394 VSUBS 0.016175f
C1165 B.n395 VSUBS 0.015411f
C1166 B.n396 VSUBS 0.007065f
C1167 B.n397 VSUBS 0.007065f
C1168 B.n398 VSUBS 0.007065f
C1169 B.n399 VSUBS 0.007065f
C1170 B.n400 VSUBS 0.007065f
C1171 B.n401 VSUBS 0.007065f
C1172 B.n402 VSUBS 0.007065f
C1173 B.n403 VSUBS 0.007065f
C1174 B.n404 VSUBS 0.007065f
C1175 B.n405 VSUBS 0.007065f
C1176 B.n406 VSUBS 0.007065f
C1177 B.n407 VSUBS 0.007065f
C1178 B.n408 VSUBS 0.007065f
C1179 B.n409 VSUBS 0.007065f
C1180 B.n410 VSUBS 0.007065f
C1181 B.n411 VSUBS 0.007065f
C1182 B.n412 VSUBS 0.007065f
C1183 B.n413 VSUBS 0.007065f
C1184 B.n414 VSUBS 0.007065f
C1185 B.n415 VSUBS 0.007065f
C1186 B.n416 VSUBS 0.007065f
C1187 B.n417 VSUBS 0.007065f
C1188 B.n418 VSUBS 0.007065f
C1189 B.n419 VSUBS 0.007065f
C1190 B.n420 VSUBS 0.007065f
C1191 B.n421 VSUBS 0.007065f
C1192 B.n422 VSUBS 0.007065f
C1193 B.n423 VSUBS 0.007065f
C1194 B.n424 VSUBS 0.007065f
C1195 B.n425 VSUBS 0.007065f
C1196 B.n426 VSUBS 0.007065f
C1197 B.n427 VSUBS 0.007065f
C1198 B.n428 VSUBS 0.007065f
C1199 B.n429 VSUBS 0.007065f
C1200 B.n430 VSUBS 0.007065f
C1201 B.n431 VSUBS 0.007065f
C1202 B.n432 VSUBS 0.007065f
C1203 B.n433 VSUBS 0.007065f
C1204 B.n434 VSUBS 0.007065f
C1205 B.n435 VSUBS 0.007065f
C1206 B.n436 VSUBS 0.007065f
C1207 B.n437 VSUBS 0.007065f
C1208 B.n438 VSUBS 0.007065f
C1209 B.n439 VSUBS 0.007065f
C1210 B.n440 VSUBS 0.007065f
C1211 B.n441 VSUBS 0.007065f
C1212 B.n442 VSUBS 0.007065f
C1213 B.n443 VSUBS 0.007065f
C1214 B.n444 VSUBS 0.007065f
C1215 B.n445 VSUBS 0.007065f
C1216 B.n446 VSUBS 0.007065f
C1217 B.n447 VSUBS 0.007065f
C1218 B.n448 VSUBS 0.007065f
C1219 B.n449 VSUBS 0.007065f
C1220 B.n450 VSUBS 0.007065f
C1221 B.n451 VSUBS 0.007065f
C1222 B.n452 VSUBS 0.007065f
C1223 B.n453 VSUBS 0.007065f
C1224 B.n454 VSUBS 0.007065f
C1225 B.n455 VSUBS 0.007065f
C1226 B.n456 VSUBS 0.007065f
C1227 B.n457 VSUBS 0.007065f
C1228 B.n458 VSUBS 0.007065f
C1229 B.n459 VSUBS 0.007065f
C1230 B.n460 VSUBS 0.007065f
C1231 B.n461 VSUBS 0.007065f
C1232 B.n462 VSUBS 0.007065f
C1233 B.n463 VSUBS 0.007065f
C1234 B.n464 VSUBS 0.007065f
C1235 B.n465 VSUBS 0.007065f
C1236 B.n466 VSUBS 0.007065f
C1237 B.n467 VSUBS 0.007065f
C1238 B.n468 VSUBS 0.007065f
C1239 B.n469 VSUBS 0.007065f
C1240 B.n470 VSUBS 0.007065f
C1241 B.n471 VSUBS 0.007065f
C1242 B.n472 VSUBS 0.007065f
C1243 B.n473 VSUBS 0.015411f
C1244 B.n474 VSUBS 0.016175f
C1245 B.n475 VSUBS 0.01528f
C1246 B.n476 VSUBS 0.007065f
C1247 B.n477 VSUBS 0.007065f
C1248 B.n478 VSUBS 0.007065f
C1249 B.n479 VSUBS 0.007065f
C1250 B.n480 VSUBS 0.007065f
C1251 B.n481 VSUBS 0.007065f
C1252 B.n482 VSUBS 0.007065f
C1253 B.n483 VSUBS 0.007065f
C1254 B.n484 VSUBS 0.007065f
C1255 B.n485 VSUBS 0.007065f
C1256 B.n486 VSUBS 0.007065f
C1257 B.n487 VSUBS 0.007065f
C1258 B.n488 VSUBS 0.007065f
C1259 B.n489 VSUBS 0.007065f
C1260 B.n490 VSUBS 0.007065f
C1261 B.n491 VSUBS 0.007065f
C1262 B.n492 VSUBS 0.007065f
C1263 B.n493 VSUBS 0.007065f
C1264 B.n494 VSUBS 0.007065f
C1265 B.n495 VSUBS 0.007065f
C1266 B.n496 VSUBS 0.007065f
C1267 B.n497 VSUBS 0.007065f
C1268 B.n498 VSUBS 0.007065f
C1269 B.n499 VSUBS 0.007065f
C1270 B.n500 VSUBS 0.007065f
C1271 B.n501 VSUBS 0.007065f
C1272 B.n502 VSUBS 0.007065f
C1273 B.n503 VSUBS 0.007065f
C1274 B.n504 VSUBS 0.007065f
C1275 B.n505 VSUBS 0.007065f
C1276 B.n506 VSUBS 0.007065f
C1277 B.n507 VSUBS 0.007065f
C1278 B.n508 VSUBS 0.007065f
C1279 B.n509 VSUBS 0.007065f
C1280 B.n510 VSUBS 0.007065f
C1281 B.n511 VSUBS 0.007065f
C1282 B.n512 VSUBS 0.007065f
C1283 B.n513 VSUBS 0.007065f
C1284 B.n514 VSUBS 0.007065f
C1285 B.n515 VSUBS 0.007065f
C1286 B.n516 VSUBS 0.007065f
C1287 B.n517 VSUBS 0.007065f
C1288 B.n518 VSUBS 0.007065f
C1289 B.n519 VSUBS 0.007065f
C1290 B.n520 VSUBS 0.007065f
C1291 B.n521 VSUBS 0.007065f
C1292 B.n522 VSUBS 0.007065f
C1293 B.n523 VSUBS 0.007065f
C1294 B.n524 VSUBS 0.007065f
C1295 B.n525 VSUBS 0.007065f
C1296 B.n526 VSUBS 0.007065f
C1297 B.n527 VSUBS 0.007065f
C1298 B.n528 VSUBS 0.007065f
C1299 B.n529 VSUBS 0.007065f
C1300 B.n530 VSUBS 0.007065f
C1301 B.n531 VSUBS 0.007065f
C1302 B.n532 VSUBS 0.007065f
C1303 B.n533 VSUBS 0.007065f
C1304 B.n534 VSUBS 0.007065f
C1305 B.n535 VSUBS 0.007065f
C1306 B.n536 VSUBS 0.007065f
C1307 B.n537 VSUBS 0.007065f
C1308 B.n538 VSUBS 0.007065f
C1309 B.n539 VSUBS 0.007065f
C1310 B.n540 VSUBS 0.007065f
C1311 B.n541 VSUBS 0.007065f
C1312 B.n542 VSUBS 0.007065f
C1313 B.n543 VSUBS 0.007065f
C1314 B.n544 VSUBS 0.007065f
C1315 B.n545 VSUBS 0.007065f
C1316 B.n546 VSUBS 0.007065f
C1317 B.n547 VSUBS 0.007065f
C1318 B.n548 VSUBS 0.007065f
C1319 B.n549 VSUBS 0.007065f
C1320 B.n550 VSUBS 0.007065f
C1321 B.n551 VSUBS 0.007065f
C1322 B.n552 VSUBS 0.007065f
C1323 B.n553 VSUBS 0.007065f
C1324 B.n554 VSUBS 0.004883f
C1325 B.n555 VSUBS 0.016369f
C1326 B.n556 VSUBS 0.005715f
C1327 B.n557 VSUBS 0.007065f
C1328 B.n558 VSUBS 0.007065f
C1329 B.n559 VSUBS 0.007065f
C1330 B.n560 VSUBS 0.007065f
C1331 B.n561 VSUBS 0.007065f
C1332 B.n562 VSUBS 0.007065f
C1333 B.n563 VSUBS 0.007065f
C1334 B.n564 VSUBS 0.007065f
C1335 B.n565 VSUBS 0.007065f
C1336 B.n566 VSUBS 0.007065f
C1337 B.n567 VSUBS 0.007065f
C1338 B.n568 VSUBS 0.005715f
C1339 B.n569 VSUBS 0.007065f
C1340 B.n570 VSUBS 0.007065f
C1341 B.n571 VSUBS 0.004883f
C1342 B.n572 VSUBS 0.007065f
C1343 B.n573 VSUBS 0.007065f
C1344 B.n574 VSUBS 0.007065f
C1345 B.n575 VSUBS 0.007065f
C1346 B.n576 VSUBS 0.007065f
C1347 B.n577 VSUBS 0.007065f
C1348 B.n578 VSUBS 0.007065f
C1349 B.n579 VSUBS 0.007065f
C1350 B.n580 VSUBS 0.007065f
C1351 B.n581 VSUBS 0.007065f
C1352 B.n582 VSUBS 0.007065f
C1353 B.n583 VSUBS 0.007065f
C1354 B.n584 VSUBS 0.007065f
C1355 B.n585 VSUBS 0.007065f
C1356 B.n586 VSUBS 0.007065f
C1357 B.n587 VSUBS 0.007065f
C1358 B.n588 VSUBS 0.007065f
C1359 B.n589 VSUBS 0.007065f
C1360 B.n590 VSUBS 0.007065f
C1361 B.n591 VSUBS 0.007065f
C1362 B.n592 VSUBS 0.007065f
C1363 B.n593 VSUBS 0.007065f
C1364 B.n594 VSUBS 0.007065f
C1365 B.n595 VSUBS 0.007065f
C1366 B.n596 VSUBS 0.007065f
C1367 B.n597 VSUBS 0.007065f
C1368 B.n598 VSUBS 0.007065f
C1369 B.n599 VSUBS 0.007065f
C1370 B.n600 VSUBS 0.007065f
C1371 B.n601 VSUBS 0.007065f
C1372 B.n602 VSUBS 0.007065f
C1373 B.n603 VSUBS 0.007065f
C1374 B.n604 VSUBS 0.007065f
C1375 B.n605 VSUBS 0.007065f
C1376 B.n606 VSUBS 0.007065f
C1377 B.n607 VSUBS 0.007065f
C1378 B.n608 VSUBS 0.007065f
C1379 B.n609 VSUBS 0.007065f
C1380 B.n610 VSUBS 0.007065f
C1381 B.n611 VSUBS 0.007065f
C1382 B.n612 VSUBS 0.007065f
C1383 B.n613 VSUBS 0.007065f
C1384 B.n614 VSUBS 0.007065f
C1385 B.n615 VSUBS 0.007065f
C1386 B.n616 VSUBS 0.007065f
C1387 B.n617 VSUBS 0.007065f
C1388 B.n618 VSUBS 0.007065f
C1389 B.n619 VSUBS 0.007065f
C1390 B.n620 VSUBS 0.007065f
C1391 B.n621 VSUBS 0.007065f
C1392 B.n622 VSUBS 0.007065f
C1393 B.n623 VSUBS 0.007065f
C1394 B.n624 VSUBS 0.007065f
C1395 B.n625 VSUBS 0.007065f
C1396 B.n626 VSUBS 0.007065f
C1397 B.n627 VSUBS 0.007065f
C1398 B.n628 VSUBS 0.007065f
C1399 B.n629 VSUBS 0.007065f
C1400 B.n630 VSUBS 0.007065f
C1401 B.n631 VSUBS 0.007065f
C1402 B.n632 VSUBS 0.007065f
C1403 B.n633 VSUBS 0.007065f
C1404 B.n634 VSUBS 0.007065f
C1405 B.n635 VSUBS 0.007065f
C1406 B.n636 VSUBS 0.007065f
C1407 B.n637 VSUBS 0.007065f
C1408 B.n638 VSUBS 0.007065f
C1409 B.n639 VSUBS 0.007065f
C1410 B.n640 VSUBS 0.007065f
C1411 B.n641 VSUBS 0.007065f
C1412 B.n642 VSUBS 0.007065f
C1413 B.n643 VSUBS 0.007065f
C1414 B.n644 VSUBS 0.007065f
C1415 B.n645 VSUBS 0.007065f
C1416 B.n646 VSUBS 0.007065f
C1417 B.n647 VSUBS 0.007065f
C1418 B.n648 VSUBS 0.007065f
C1419 B.n649 VSUBS 0.007065f
C1420 B.n650 VSUBS 0.016175f
C1421 B.n651 VSUBS 0.015411f
C1422 B.n652 VSUBS 0.015411f
C1423 B.n653 VSUBS 0.007065f
C1424 B.n654 VSUBS 0.007065f
C1425 B.n655 VSUBS 0.007065f
C1426 B.n656 VSUBS 0.007065f
C1427 B.n657 VSUBS 0.007065f
C1428 B.n658 VSUBS 0.007065f
C1429 B.n659 VSUBS 0.007065f
C1430 B.n660 VSUBS 0.007065f
C1431 B.n661 VSUBS 0.007065f
C1432 B.n662 VSUBS 0.007065f
C1433 B.n663 VSUBS 0.007065f
C1434 B.n664 VSUBS 0.007065f
C1435 B.n665 VSUBS 0.007065f
C1436 B.n666 VSUBS 0.007065f
C1437 B.n667 VSUBS 0.007065f
C1438 B.n668 VSUBS 0.007065f
C1439 B.n669 VSUBS 0.007065f
C1440 B.n670 VSUBS 0.007065f
C1441 B.n671 VSUBS 0.007065f
C1442 B.n672 VSUBS 0.007065f
C1443 B.n673 VSUBS 0.007065f
C1444 B.n674 VSUBS 0.007065f
C1445 B.n675 VSUBS 0.007065f
C1446 B.n676 VSUBS 0.007065f
C1447 B.n677 VSUBS 0.007065f
C1448 B.n678 VSUBS 0.007065f
C1449 B.n679 VSUBS 0.007065f
C1450 B.n680 VSUBS 0.007065f
C1451 B.n681 VSUBS 0.007065f
C1452 B.n682 VSUBS 0.007065f
C1453 B.n683 VSUBS 0.007065f
C1454 B.n684 VSUBS 0.007065f
C1455 B.n685 VSUBS 0.007065f
C1456 B.n686 VSUBS 0.007065f
C1457 B.n687 VSUBS 0.007065f
C1458 B.n688 VSUBS 0.007065f
C1459 B.n689 VSUBS 0.007065f
C1460 B.n690 VSUBS 0.007065f
C1461 B.n691 VSUBS 0.015998f
.ends

