* NGSPICE file created from diff_pair_sample_1279.ext - technology: sky130A

.subckt diff_pair_sample_1279 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=0 ps=0 w=11.81 l=1.46
X1 VTAIL.t19 VN.t0 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X2 VDD2.t4 VN.t1 VTAIL.t18 B.t9 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=1.94865 ps=12.14 w=11.81 l=1.46
X3 VDD1.t9 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X4 VTAIL.t2 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X5 VDD1.t7 VP.t2 VTAIL.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=1.94865 ps=12.14 w=11.81 l=1.46
X6 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=0 ps=0 w=11.81 l=1.46
X7 VTAIL.t17 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X8 VTAIL.t1 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X9 VDD2.t9 VN.t3 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X10 VDD2.t0 VN.t4 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=1.94865 ps=12.14 w=11.81 l=1.46
X11 VTAIL.t8 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X12 VDD1.t4 VP.t5 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=4.6059 ps=24.4 w=11.81 l=1.46
X13 VDD2.t3 VN.t5 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=4.6059 ps=24.4 w=11.81 l=1.46
X14 VDD2.t7 VN.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X15 VDD1.t3 VP.t6 VTAIL.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=4.6059 ps=24.4 w=11.81 l=1.46
X16 VDD2.t8 VN.t7 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=4.6059 ps=24.4 w=11.81 l=1.46
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=0 ps=0 w=11.81 l=1.46
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=0 ps=0 w=11.81 l=1.46
X19 VDD1.t2 VP.t7 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X20 VTAIL.t11 VN.t8 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X21 VTAIL.t10 VN.t9 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X22 VTAIL.t4 VP.t8 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.94865 pd=12.14 as=1.94865 ps=12.14 w=11.81 l=1.46
X23 VDD1.t0 VP.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=4.6059 pd=24.4 as=1.94865 ps=12.14 w=11.81 l=1.46
R0 B.n784 B.n783 585
R1 B.n303 B.n119 585
R2 B.n302 B.n301 585
R3 B.n300 B.n299 585
R4 B.n298 B.n297 585
R5 B.n296 B.n295 585
R6 B.n294 B.n293 585
R7 B.n292 B.n291 585
R8 B.n290 B.n289 585
R9 B.n288 B.n287 585
R10 B.n286 B.n285 585
R11 B.n284 B.n283 585
R12 B.n282 B.n281 585
R13 B.n280 B.n279 585
R14 B.n278 B.n277 585
R15 B.n276 B.n275 585
R16 B.n274 B.n273 585
R17 B.n272 B.n271 585
R18 B.n270 B.n269 585
R19 B.n268 B.n267 585
R20 B.n266 B.n265 585
R21 B.n264 B.n263 585
R22 B.n262 B.n261 585
R23 B.n260 B.n259 585
R24 B.n258 B.n257 585
R25 B.n256 B.n255 585
R26 B.n254 B.n253 585
R27 B.n252 B.n251 585
R28 B.n250 B.n249 585
R29 B.n248 B.n247 585
R30 B.n246 B.n245 585
R31 B.n244 B.n243 585
R32 B.n242 B.n241 585
R33 B.n240 B.n239 585
R34 B.n238 B.n237 585
R35 B.n236 B.n235 585
R36 B.n234 B.n233 585
R37 B.n232 B.n231 585
R38 B.n230 B.n229 585
R39 B.n228 B.n227 585
R40 B.n226 B.n225 585
R41 B.n223 B.n222 585
R42 B.n221 B.n220 585
R43 B.n219 B.n218 585
R44 B.n217 B.n216 585
R45 B.n215 B.n214 585
R46 B.n213 B.n212 585
R47 B.n211 B.n210 585
R48 B.n209 B.n208 585
R49 B.n207 B.n206 585
R50 B.n205 B.n204 585
R51 B.n202 B.n201 585
R52 B.n200 B.n199 585
R53 B.n198 B.n197 585
R54 B.n196 B.n195 585
R55 B.n194 B.n193 585
R56 B.n192 B.n191 585
R57 B.n190 B.n189 585
R58 B.n188 B.n187 585
R59 B.n186 B.n185 585
R60 B.n184 B.n183 585
R61 B.n182 B.n181 585
R62 B.n180 B.n179 585
R63 B.n178 B.n177 585
R64 B.n176 B.n175 585
R65 B.n174 B.n173 585
R66 B.n172 B.n171 585
R67 B.n170 B.n169 585
R68 B.n168 B.n167 585
R69 B.n166 B.n165 585
R70 B.n164 B.n163 585
R71 B.n162 B.n161 585
R72 B.n160 B.n159 585
R73 B.n158 B.n157 585
R74 B.n156 B.n155 585
R75 B.n154 B.n153 585
R76 B.n152 B.n151 585
R77 B.n150 B.n149 585
R78 B.n148 B.n147 585
R79 B.n146 B.n145 585
R80 B.n144 B.n143 585
R81 B.n142 B.n141 585
R82 B.n140 B.n139 585
R83 B.n138 B.n137 585
R84 B.n136 B.n135 585
R85 B.n134 B.n133 585
R86 B.n132 B.n131 585
R87 B.n130 B.n129 585
R88 B.n128 B.n127 585
R89 B.n126 B.n125 585
R90 B.n74 B.n73 585
R91 B.n789 B.n788 585
R92 B.n782 B.n120 585
R93 B.n120 B.n71 585
R94 B.n781 B.n70 585
R95 B.n793 B.n70 585
R96 B.n780 B.n69 585
R97 B.n794 B.n69 585
R98 B.n779 B.n68 585
R99 B.n795 B.n68 585
R100 B.n778 B.n777 585
R101 B.n777 B.n64 585
R102 B.n776 B.n63 585
R103 B.n801 B.n63 585
R104 B.n775 B.n62 585
R105 B.n802 B.n62 585
R106 B.n774 B.n61 585
R107 B.n803 B.n61 585
R108 B.n773 B.n772 585
R109 B.n772 B.n57 585
R110 B.n771 B.n56 585
R111 B.n809 B.n56 585
R112 B.n770 B.n55 585
R113 B.n810 B.n55 585
R114 B.n769 B.n54 585
R115 B.n811 B.n54 585
R116 B.n768 B.n767 585
R117 B.n767 B.n50 585
R118 B.n766 B.n49 585
R119 B.n817 B.n49 585
R120 B.n765 B.n48 585
R121 B.n818 B.n48 585
R122 B.n764 B.n47 585
R123 B.n819 B.n47 585
R124 B.n763 B.n762 585
R125 B.n762 B.n43 585
R126 B.n761 B.n42 585
R127 B.n825 B.n42 585
R128 B.n760 B.n41 585
R129 B.n826 B.n41 585
R130 B.n759 B.n40 585
R131 B.n827 B.n40 585
R132 B.n758 B.n757 585
R133 B.n757 B.n36 585
R134 B.n756 B.n35 585
R135 B.n833 B.n35 585
R136 B.n755 B.n34 585
R137 B.n834 B.n34 585
R138 B.n754 B.n33 585
R139 B.n835 B.n33 585
R140 B.n753 B.n752 585
R141 B.n752 B.n32 585
R142 B.n751 B.n28 585
R143 B.n841 B.n28 585
R144 B.n750 B.n27 585
R145 B.n842 B.n27 585
R146 B.n749 B.n26 585
R147 B.n843 B.n26 585
R148 B.n748 B.n747 585
R149 B.n747 B.n22 585
R150 B.n746 B.n21 585
R151 B.n849 B.n21 585
R152 B.n745 B.n20 585
R153 B.t2 B.n20 585
R154 B.n744 B.n19 585
R155 B.n850 B.n19 585
R156 B.n743 B.n742 585
R157 B.n742 B.n15 585
R158 B.n741 B.n14 585
R159 B.n856 B.n14 585
R160 B.n740 B.n13 585
R161 B.n857 B.n13 585
R162 B.n739 B.n12 585
R163 B.n858 B.n12 585
R164 B.n738 B.n737 585
R165 B.n737 B.n736 585
R166 B.n735 B.n734 585
R167 B.n735 B.n8 585
R168 B.n733 B.n7 585
R169 B.n865 B.n7 585
R170 B.n732 B.n6 585
R171 B.n866 B.n6 585
R172 B.n731 B.n5 585
R173 B.n867 B.n5 585
R174 B.n730 B.n729 585
R175 B.n729 B.n4 585
R176 B.n728 B.n304 585
R177 B.n728 B.n727 585
R178 B.n718 B.n305 585
R179 B.n306 B.n305 585
R180 B.n720 B.n719 585
R181 B.n721 B.n720 585
R182 B.n717 B.n311 585
R183 B.n311 B.n310 585
R184 B.n716 B.n715 585
R185 B.n715 B.n714 585
R186 B.n313 B.n312 585
R187 B.n314 B.n313 585
R188 B.n707 B.n706 585
R189 B.n708 B.n707 585
R190 B.n705 B.n318 585
R191 B.n318 B.t3 585
R192 B.n704 B.n703 585
R193 B.n703 B.n702 585
R194 B.n320 B.n319 585
R195 B.n321 B.n320 585
R196 B.n695 B.n694 585
R197 B.n696 B.n695 585
R198 B.n693 B.n326 585
R199 B.n326 B.n325 585
R200 B.n692 B.n691 585
R201 B.n691 B.n690 585
R202 B.n328 B.n327 585
R203 B.n683 B.n328 585
R204 B.n682 B.n681 585
R205 B.n684 B.n682 585
R206 B.n680 B.n333 585
R207 B.n333 B.n332 585
R208 B.n679 B.n678 585
R209 B.n678 B.n677 585
R210 B.n335 B.n334 585
R211 B.n336 B.n335 585
R212 B.n670 B.n669 585
R213 B.n671 B.n670 585
R214 B.n668 B.n341 585
R215 B.n341 B.n340 585
R216 B.n667 B.n666 585
R217 B.n666 B.n665 585
R218 B.n343 B.n342 585
R219 B.n344 B.n343 585
R220 B.n658 B.n657 585
R221 B.n659 B.n658 585
R222 B.n656 B.n348 585
R223 B.n352 B.n348 585
R224 B.n655 B.n654 585
R225 B.n654 B.n653 585
R226 B.n350 B.n349 585
R227 B.n351 B.n350 585
R228 B.n646 B.n645 585
R229 B.n647 B.n646 585
R230 B.n644 B.n357 585
R231 B.n357 B.n356 585
R232 B.n643 B.n642 585
R233 B.n642 B.n641 585
R234 B.n359 B.n358 585
R235 B.n360 B.n359 585
R236 B.n634 B.n633 585
R237 B.n635 B.n634 585
R238 B.n632 B.n365 585
R239 B.n365 B.n364 585
R240 B.n631 B.n630 585
R241 B.n630 B.n629 585
R242 B.n367 B.n366 585
R243 B.n368 B.n367 585
R244 B.n622 B.n621 585
R245 B.n623 B.n622 585
R246 B.n620 B.n373 585
R247 B.n373 B.n372 585
R248 B.n619 B.n618 585
R249 B.n618 B.n617 585
R250 B.n375 B.n374 585
R251 B.n376 B.n375 585
R252 B.n613 B.n612 585
R253 B.n379 B.n378 585
R254 B.n609 B.n608 585
R255 B.n610 B.n609 585
R256 B.n607 B.n425 585
R257 B.n606 B.n605 585
R258 B.n604 B.n603 585
R259 B.n602 B.n601 585
R260 B.n600 B.n599 585
R261 B.n598 B.n597 585
R262 B.n596 B.n595 585
R263 B.n594 B.n593 585
R264 B.n592 B.n591 585
R265 B.n590 B.n589 585
R266 B.n588 B.n587 585
R267 B.n586 B.n585 585
R268 B.n584 B.n583 585
R269 B.n582 B.n581 585
R270 B.n580 B.n579 585
R271 B.n578 B.n577 585
R272 B.n576 B.n575 585
R273 B.n574 B.n573 585
R274 B.n572 B.n571 585
R275 B.n570 B.n569 585
R276 B.n568 B.n567 585
R277 B.n566 B.n565 585
R278 B.n564 B.n563 585
R279 B.n562 B.n561 585
R280 B.n560 B.n559 585
R281 B.n558 B.n557 585
R282 B.n556 B.n555 585
R283 B.n554 B.n553 585
R284 B.n552 B.n551 585
R285 B.n550 B.n549 585
R286 B.n548 B.n547 585
R287 B.n546 B.n545 585
R288 B.n544 B.n543 585
R289 B.n542 B.n541 585
R290 B.n540 B.n539 585
R291 B.n538 B.n537 585
R292 B.n536 B.n535 585
R293 B.n534 B.n533 585
R294 B.n532 B.n531 585
R295 B.n530 B.n529 585
R296 B.n528 B.n527 585
R297 B.n526 B.n525 585
R298 B.n524 B.n523 585
R299 B.n522 B.n521 585
R300 B.n520 B.n519 585
R301 B.n518 B.n517 585
R302 B.n516 B.n515 585
R303 B.n514 B.n513 585
R304 B.n512 B.n511 585
R305 B.n510 B.n509 585
R306 B.n508 B.n507 585
R307 B.n506 B.n505 585
R308 B.n504 B.n503 585
R309 B.n502 B.n501 585
R310 B.n500 B.n499 585
R311 B.n498 B.n497 585
R312 B.n496 B.n495 585
R313 B.n494 B.n493 585
R314 B.n492 B.n491 585
R315 B.n490 B.n489 585
R316 B.n488 B.n487 585
R317 B.n486 B.n485 585
R318 B.n484 B.n483 585
R319 B.n482 B.n481 585
R320 B.n480 B.n479 585
R321 B.n478 B.n477 585
R322 B.n476 B.n475 585
R323 B.n474 B.n473 585
R324 B.n472 B.n471 585
R325 B.n470 B.n469 585
R326 B.n468 B.n467 585
R327 B.n466 B.n465 585
R328 B.n464 B.n463 585
R329 B.n462 B.n461 585
R330 B.n460 B.n459 585
R331 B.n458 B.n457 585
R332 B.n456 B.n455 585
R333 B.n454 B.n453 585
R334 B.n452 B.n451 585
R335 B.n450 B.n449 585
R336 B.n448 B.n447 585
R337 B.n446 B.n445 585
R338 B.n444 B.n443 585
R339 B.n442 B.n441 585
R340 B.n440 B.n439 585
R341 B.n438 B.n437 585
R342 B.n436 B.n435 585
R343 B.n434 B.n433 585
R344 B.n432 B.n424 585
R345 B.n610 B.n424 585
R346 B.n614 B.n377 585
R347 B.n377 B.n376 585
R348 B.n616 B.n615 585
R349 B.n617 B.n616 585
R350 B.n371 B.n370 585
R351 B.n372 B.n371 585
R352 B.n625 B.n624 585
R353 B.n624 B.n623 585
R354 B.n626 B.n369 585
R355 B.n369 B.n368 585
R356 B.n628 B.n627 585
R357 B.n629 B.n628 585
R358 B.n363 B.n362 585
R359 B.n364 B.n363 585
R360 B.n637 B.n636 585
R361 B.n636 B.n635 585
R362 B.n638 B.n361 585
R363 B.n361 B.n360 585
R364 B.n640 B.n639 585
R365 B.n641 B.n640 585
R366 B.n355 B.n354 585
R367 B.n356 B.n355 585
R368 B.n649 B.n648 585
R369 B.n648 B.n647 585
R370 B.n650 B.n353 585
R371 B.n353 B.n351 585
R372 B.n652 B.n651 585
R373 B.n653 B.n652 585
R374 B.n347 B.n346 585
R375 B.n352 B.n347 585
R376 B.n661 B.n660 585
R377 B.n660 B.n659 585
R378 B.n662 B.n345 585
R379 B.n345 B.n344 585
R380 B.n664 B.n663 585
R381 B.n665 B.n664 585
R382 B.n339 B.n338 585
R383 B.n340 B.n339 585
R384 B.n673 B.n672 585
R385 B.n672 B.n671 585
R386 B.n674 B.n337 585
R387 B.n337 B.n336 585
R388 B.n676 B.n675 585
R389 B.n677 B.n676 585
R390 B.n331 B.n330 585
R391 B.n332 B.n331 585
R392 B.n686 B.n685 585
R393 B.n685 B.n684 585
R394 B.n687 B.n329 585
R395 B.n683 B.n329 585
R396 B.n689 B.n688 585
R397 B.n690 B.n689 585
R398 B.n324 B.n323 585
R399 B.n325 B.n324 585
R400 B.n698 B.n697 585
R401 B.n697 B.n696 585
R402 B.n699 B.n322 585
R403 B.n322 B.n321 585
R404 B.n701 B.n700 585
R405 B.n702 B.n701 585
R406 B.n317 B.n316 585
R407 B.t3 B.n317 585
R408 B.n710 B.n709 585
R409 B.n709 B.n708 585
R410 B.n711 B.n315 585
R411 B.n315 B.n314 585
R412 B.n713 B.n712 585
R413 B.n714 B.n713 585
R414 B.n309 B.n308 585
R415 B.n310 B.n309 585
R416 B.n723 B.n722 585
R417 B.n722 B.n721 585
R418 B.n724 B.n307 585
R419 B.n307 B.n306 585
R420 B.n726 B.n725 585
R421 B.n727 B.n726 585
R422 B.n3 B.n0 585
R423 B.n4 B.n3 585
R424 B.n864 B.n1 585
R425 B.n865 B.n864 585
R426 B.n863 B.n862 585
R427 B.n863 B.n8 585
R428 B.n861 B.n9 585
R429 B.n736 B.n9 585
R430 B.n860 B.n859 585
R431 B.n859 B.n858 585
R432 B.n11 B.n10 585
R433 B.n857 B.n11 585
R434 B.n855 B.n854 585
R435 B.n856 B.n855 585
R436 B.n853 B.n16 585
R437 B.n16 B.n15 585
R438 B.n852 B.n851 585
R439 B.n851 B.n850 585
R440 B.n18 B.n17 585
R441 B.t2 B.n18 585
R442 B.n848 B.n847 585
R443 B.n849 B.n848 585
R444 B.n846 B.n23 585
R445 B.n23 B.n22 585
R446 B.n845 B.n844 585
R447 B.n844 B.n843 585
R448 B.n25 B.n24 585
R449 B.n842 B.n25 585
R450 B.n840 B.n839 585
R451 B.n841 B.n840 585
R452 B.n838 B.n29 585
R453 B.n32 B.n29 585
R454 B.n837 B.n836 585
R455 B.n836 B.n835 585
R456 B.n31 B.n30 585
R457 B.n834 B.n31 585
R458 B.n832 B.n831 585
R459 B.n833 B.n832 585
R460 B.n830 B.n37 585
R461 B.n37 B.n36 585
R462 B.n829 B.n828 585
R463 B.n828 B.n827 585
R464 B.n39 B.n38 585
R465 B.n826 B.n39 585
R466 B.n824 B.n823 585
R467 B.n825 B.n824 585
R468 B.n822 B.n44 585
R469 B.n44 B.n43 585
R470 B.n821 B.n820 585
R471 B.n820 B.n819 585
R472 B.n46 B.n45 585
R473 B.n818 B.n46 585
R474 B.n816 B.n815 585
R475 B.n817 B.n816 585
R476 B.n814 B.n51 585
R477 B.n51 B.n50 585
R478 B.n813 B.n812 585
R479 B.n812 B.n811 585
R480 B.n53 B.n52 585
R481 B.n810 B.n53 585
R482 B.n808 B.n807 585
R483 B.n809 B.n808 585
R484 B.n806 B.n58 585
R485 B.n58 B.n57 585
R486 B.n805 B.n804 585
R487 B.n804 B.n803 585
R488 B.n60 B.n59 585
R489 B.n802 B.n60 585
R490 B.n800 B.n799 585
R491 B.n801 B.n800 585
R492 B.n798 B.n65 585
R493 B.n65 B.n64 585
R494 B.n797 B.n796 585
R495 B.n796 B.n795 585
R496 B.n67 B.n66 585
R497 B.n794 B.n67 585
R498 B.n792 B.n791 585
R499 B.n793 B.n792 585
R500 B.n790 B.n72 585
R501 B.n72 B.n71 585
R502 B.n868 B.n867 585
R503 B.n866 B.n2 585
R504 B.n788 B.n72 506.916
R505 B.n784 B.n120 506.916
R506 B.n424 B.n375 506.916
R507 B.n612 B.n377 506.916
R508 B.n123 B.t18 400.233
R509 B.n121 B.t14 400.233
R510 B.n429 B.t21 400.233
R511 B.n426 B.t10 400.233
R512 B.n786 B.n785 256.663
R513 B.n786 B.n118 256.663
R514 B.n786 B.n117 256.663
R515 B.n786 B.n116 256.663
R516 B.n786 B.n115 256.663
R517 B.n786 B.n114 256.663
R518 B.n786 B.n113 256.663
R519 B.n786 B.n112 256.663
R520 B.n786 B.n111 256.663
R521 B.n786 B.n110 256.663
R522 B.n786 B.n109 256.663
R523 B.n786 B.n108 256.663
R524 B.n786 B.n107 256.663
R525 B.n786 B.n106 256.663
R526 B.n786 B.n105 256.663
R527 B.n786 B.n104 256.663
R528 B.n786 B.n103 256.663
R529 B.n786 B.n102 256.663
R530 B.n786 B.n101 256.663
R531 B.n786 B.n100 256.663
R532 B.n786 B.n99 256.663
R533 B.n786 B.n98 256.663
R534 B.n786 B.n97 256.663
R535 B.n786 B.n96 256.663
R536 B.n786 B.n95 256.663
R537 B.n786 B.n94 256.663
R538 B.n786 B.n93 256.663
R539 B.n786 B.n92 256.663
R540 B.n786 B.n91 256.663
R541 B.n786 B.n90 256.663
R542 B.n786 B.n89 256.663
R543 B.n786 B.n88 256.663
R544 B.n786 B.n87 256.663
R545 B.n786 B.n86 256.663
R546 B.n786 B.n85 256.663
R547 B.n786 B.n84 256.663
R548 B.n786 B.n83 256.663
R549 B.n786 B.n82 256.663
R550 B.n786 B.n81 256.663
R551 B.n786 B.n80 256.663
R552 B.n786 B.n79 256.663
R553 B.n786 B.n78 256.663
R554 B.n786 B.n77 256.663
R555 B.n786 B.n76 256.663
R556 B.n786 B.n75 256.663
R557 B.n787 B.n786 256.663
R558 B.n611 B.n610 256.663
R559 B.n610 B.n380 256.663
R560 B.n610 B.n381 256.663
R561 B.n610 B.n382 256.663
R562 B.n610 B.n383 256.663
R563 B.n610 B.n384 256.663
R564 B.n610 B.n385 256.663
R565 B.n610 B.n386 256.663
R566 B.n610 B.n387 256.663
R567 B.n610 B.n388 256.663
R568 B.n610 B.n389 256.663
R569 B.n610 B.n390 256.663
R570 B.n610 B.n391 256.663
R571 B.n610 B.n392 256.663
R572 B.n610 B.n393 256.663
R573 B.n610 B.n394 256.663
R574 B.n610 B.n395 256.663
R575 B.n610 B.n396 256.663
R576 B.n610 B.n397 256.663
R577 B.n610 B.n398 256.663
R578 B.n610 B.n399 256.663
R579 B.n610 B.n400 256.663
R580 B.n610 B.n401 256.663
R581 B.n610 B.n402 256.663
R582 B.n610 B.n403 256.663
R583 B.n610 B.n404 256.663
R584 B.n610 B.n405 256.663
R585 B.n610 B.n406 256.663
R586 B.n610 B.n407 256.663
R587 B.n610 B.n408 256.663
R588 B.n610 B.n409 256.663
R589 B.n610 B.n410 256.663
R590 B.n610 B.n411 256.663
R591 B.n610 B.n412 256.663
R592 B.n610 B.n413 256.663
R593 B.n610 B.n414 256.663
R594 B.n610 B.n415 256.663
R595 B.n610 B.n416 256.663
R596 B.n610 B.n417 256.663
R597 B.n610 B.n418 256.663
R598 B.n610 B.n419 256.663
R599 B.n610 B.n420 256.663
R600 B.n610 B.n421 256.663
R601 B.n610 B.n422 256.663
R602 B.n610 B.n423 256.663
R603 B.n870 B.n869 256.663
R604 B.n125 B.n74 163.367
R605 B.n129 B.n128 163.367
R606 B.n133 B.n132 163.367
R607 B.n137 B.n136 163.367
R608 B.n141 B.n140 163.367
R609 B.n145 B.n144 163.367
R610 B.n149 B.n148 163.367
R611 B.n153 B.n152 163.367
R612 B.n157 B.n156 163.367
R613 B.n161 B.n160 163.367
R614 B.n165 B.n164 163.367
R615 B.n169 B.n168 163.367
R616 B.n173 B.n172 163.367
R617 B.n177 B.n176 163.367
R618 B.n181 B.n180 163.367
R619 B.n185 B.n184 163.367
R620 B.n189 B.n188 163.367
R621 B.n193 B.n192 163.367
R622 B.n197 B.n196 163.367
R623 B.n201 B.n200 163.367
R624 B.n206 B.n205 163.367
R625 B.n210 B.n209 163.367
R626 B.n214 B.n213 163.367
R627 B.n218 B.n217 163.367
R628 B.n222 B.n221 163.367
R629 B.n227 B.n226 163.367
R630 B.n231 B.n230 163.367
R631 B.n235 B.n234 163.367
R632 B.n239 B.n238 163.367
R633 B.n243 B.n242 163.367
R634 B.n247 B.n246 163.367
R635 B.n251 B.n250 163.367
R636 B.n255 B.n254 163.367
R637 B.n259 B.n258 163.367
R638 B.n263 B.n262 163.367
R639 B.n267 B.n266 163.367
R640 B.n271 B.n270 163.367
R641 B.n275 B.n274 163.367
R642 B.n279 B.n278 163.367
R643 B.n283 B.n282 163.367
R644 B.n287 B.n286 163.367
R645 B.n291 B.n290 163.367
R646 B.n295 B.n294 163.367
R647 B.n299 B.n298 163.367
R648 B.n301 B.n119 163.367
R649 B.n618 B.n375 163.367
R650 B.n618 B.n373 163.367
R651 B.n622 B.n373 163.367
R652 B.n622 B.n367 163.367
R653 B.n630 B.n367 163.367
R654 B.n630 B.n365 163.367
R655 B.n634 B.n365 163.367
R656 B.n634 B.n359 163.367
R657 B.n642 B.n359 163.367
R658 B.n642 B.n357 163.367
R659 B.n646 B.n357 163.367
R660 B.n646 B.n350 163.367
R661 B.n654 B.n350 163.367
R662 B.n654 B.n348 163.367
R663 B.n658 B.n348 163.367
R664 B.n658 B.n343 163.367
R665 B.n666 B.n343 163.367
R666 B.n666 B.n341 163.367
R667 B.n670 B.n341 163.367
R668 B.n670 B.n335 163.367
R669 B.n678 B.n335 163.367
R670 B.n678 B.n333 163.367
R671 B.n682 B.n333 163.367
R672 B.n682 B.n328 163.367
R673 B.n691 B.n328 163.367
R674 B.n691 B.n326 163.367
R675 B.n695 B.n326 163.367
R676 B.n695 B.n320 163.367
R677 B.n703 B.n320 163.367
R678 B.n703 B.n318 163.367
R679 B.n707 B.n318 163.367
R680 B.n707 B.n313 163.367
R681 B.n715 B.n313 163.367
R682 B.n715 B.n311 163.367
R683 B.n720 B.n311 163.367
R684 B.n720 B.n305 163.367
R685 B.n728 B.n305 163.367
R686 B.n729 B.n728 163.367
R687 B.n729 B.n5 163.367
R688 B.n6 B.n5 163.367
R689 B.n7 B.n6 163.367
R690 B.n735 B.n7 163.367
R691 B.n737 B.n735 163.367
R692 B.n737 B.n12 163.367
R693 B.n13 B.n12 163.367
R694 B.n14 B.n13 163.367
R695 B.n742 B.n14 163.367
R696 B.n742 B.n19 163.367
R697 B.n20 B.n19 163.367
R698 B.n21 B.n20 163.367
R699 B.n747 B.n21 163.367
R700 B.n747 B.n26 163.367
R701 B.n27 B.n26 163.367
R702 B.n28 B.n27 163.367
R703 B.n752 B.n28 163.367
R704 B.n752 B.n33 163.367
R705 B.n34 B.n33 163.367
R706 B.n35 B.n34 163.367
R707 B.n757 B.n35 163.367
R708 B.n757 B.n40 163.367
R709 B.n41 B.n40 163.367
R710 B.n42 B.n41 163.367
R711 B.n762 B.n42 163.367
R712 B.n762 B.n47 163.367
R713 B.n48 B.n47 163.367
R714 B.n49 B.n48 163.367
R715 B.n767 B.n49 163.367
R716 B.n767 B.n54 163.367
R717 B.n55 B.n54 163.367
R718 B.n56 B.n55 163.367
R719 B.n772 B.n56 163.367
R720 B.n772 B.n61 163.367
R721 B.n62 B.n61 163.367
R722 B.n63 B.n62 163.367
R723 B.n777 B.n63 163.367
R724 B.n777 B.n68 163.367
R725 B.n69 B.n68 163.367
R726 B.n70 B.n69 163.367
R727 B.n120 B.n70 163.367
R728 B.n609 B.n379 163.367
R729 B.n609 B.n425 163.367
R730 B.n605 B.n604 163.367
R731 B.n601 B.n600 163.367
R732 B.n597 B.n596 163.367
R733 B.n593 B.n592 163.367
R734 B.n589 B.n588 163.367
R735 B.n585 B.n584 163.367
R736 B.n581 B.n580 163.367
R737 B.n577 B.n576 163.367
R738 B.n573 B.n572 163.367
R739 B.n569 B.n568 163.367
R740 B.n565 B.n564 163.367
R741 B.n561 B.n560 163.367
R742 B.n557 B.n556 163.367
R743 B.n553 B.n552 163.367
R744 B.n549 B.n548 163.367
R745 B.n545 B.n544 163.367
R746 B.n541 B.n540 163.367
R747 B.n537 B.n536 163.367
R748 B.n533 B.n532 163.367
R749 B.n529 B.n528 163.367
R750 B.n525 B.n524 163.367
R751 B.n521 B.n520 163.367
R752 B.n517 B.n516 163.367
R753 B.n513 B.n512 163.367
R754 B.n509 B.n508 163.367
R755 B.n505 B.n504 163.367
R756 B.n501 B.n500 163.367
R757 B.n497 B.n496 163.367
R758 B.n493 B.n492 163.367
R759 B.n489 B.n488 163.367
R760 B.n485 B.n484 163.367
R761 B.n481 B.n480 163.367
R762 B.n477 B.n476 163.367
R763 B.n473 B.n472 163.367
R764 B.n469 B.n468 163.367
R765 B.n465 B.n464 163.367
R766 B.n461 B.n460 163.367
R767 B.n457 B.n456 163.367
R768 B.n453 B.n452 163.367
R769 B.n449 B.n448 163.367
R770 B.n445 B.n444 163.367
R771 B.n441 B.n440 163.367
R772 B.n437 B.n436 163.367
R773 B.n433 B.n424 163.367
R774 B.n616 B.n377 163.367
R775 B.n616 B.n371 163.367
R776 B.n624 B.n371 163.367
R777 B.n624 B.n369 163.367
R778 B.n628 B.n369 163.367
R779 B.n628 B.n363 163.367
R780 B.n636 B.n363 163.367
R781 B.n636 B.n361 163.367
R782 B.n640 B.n361 163.367
R783 B.n640 B.n355 163.367
R784 B.n648 B.n355 163.367
R785 B.n648 B.n353 163.367
R786 B.n652 B.n353 163.367
R787 B.n652 B.n347 163.367
R788 B.n660 B.n347 163.367
R789 B.n660 B.n345 163.367
R790 B.n664 B.n345 163.367
R791 B.n664 B.n339 163.367
R792 B.n672 B.n339 163.367
R793 B.n672 B.n337 163.367
R794 B.n676 B.n337 163.367
R795 B.n676 B.n331 163.367
R796 B.n685 B.n331 163.367
R797 B.n685 B.n329 163.367
R798 B.n689 B.n329 163.367
R799 B.n689 B.n324 163.367
R800 B.n697 B.n324 163.367
R801 B.n697 B.n322 163.367
R802 B.n701 B.n322 163.367
R803 B.n701 B.n317 163.367
R804 B.n709 B.n317 163.367
R805 B.n709 B.n315 163.367
R806 B.n713 B.n315 163.367
R807 B.n713 B.n309 163.367
R808 B.n722 B.n309 163.367
R809 B.n722 B.n307 163.367
R810 B.n726 B.n307 163.367
R811 B.n726 B.n3 163.367
R812 B.n868 B.n3 163.367
R813 B.n864 B.n2 163.367
R814 B.n864 B.n863 163.367
R815 B.n863 B.n9 163.367
R816 B.n859 B.n9 163.367
R817 B.n859 B.n11 163.367
R818 B.n855 B.n11 163.367
R819 B.n855 B.n16 163.367
R820 B.n851 B.n16 163.367
R821 B.n851 B.n18 163.367
R822 B.n848 B.n18 163.367
R823 B.n848 B.n23 163.367
R824 B.n844 B.n23 163.367
R825 B.n844 B.n25 163.367
R826 B.n840 B.n25 163.367
R827 B.n840 B.n29 163.367
R828 B.n836 B.n29 163.367
R829 B.n836 B.n31 163.367
R830 B.n832 B.n31 163.367
R831 B.n832 B.n37 163.367
R832 B.n828 B.n37 163.367
R833 B.n828 B.n39 163.367
R834 B.n824 B.n39 163.367
R835 B.n824 B.n44 163.367
R836 B.n820 B.n44 163.367
R837 B.n820 B.n46 163.367
R838 B.n816 B.n46 163.367
R839 B.n816 B.n51 163.367
R840 B.n812 B.n51 163.367
R841 B.n812 B.n53 163.367
R842 B.n808 B.n53 163.367
R843 B.n808 B.n58 163.367
R844 B.n804 B.n58 163.367
R845 B.n804 B.n60 163.367
R846 B.n800 B.n60 163.367
R847 B.n800 B.n65 163.367
R848 B.n796 B.n65 163.367
R849 B.n796 B.n67 163.367
R850 B.n792 B.n67 163.367
R851 B.n792 B.n72 163.367
R852 B.n121 B.t16 107.379
R853 B.n429 B.t23 107.379
R854 B.n123 B.t19 107.365
R855 B.n426 B.t13 107.365
R856 B.n610 B.n376 88.2065
R857 B.n786 B.n71 88.2065
R858 B.n122 B.t17 72.6644
R859 B.n430 B.t22 72.6644
R860 B.n124 B.t20 72.6497
R861 B.n427 B.t12 72.6497
R862 B.n788 B.n787 71.676
R863 B.n125 B.n75 71.676
R864 B.n129 B.n76 71.676
R865 B.n133 B.n77 71.676
R866 B.n137 B.n78 71.676
R867 B.n141 B.n79 71.676
R868 B.n145 B.n80 71.676
R869 B.n149 B.n81 71.676
R870 B.n153 B.n82 71.676
R871 B.n157 B.n83 71.676
R872 B.n161 B.n84 71.676
R873 B.n165 B.n85 71.676
R874 B.n169 B.n86 71.676
R875 B.n173 B.n87 71.676
R876 B.n177 B.n88 71.676
R877 B.n181 B.n89 71.676
R878 B.n185 B.n90 71.676
R879 B.n189 B.n91 71.676
R880 B.n193 B.n92 71.676
R881 B.n197 B.n93 71.676
R882 B.n201 B.n94 71.676
R883 B.n206 B.n95 71.676
R884 B.n210 B.n96 71.676
R885 B.n214 B.n97 71.676
R886 B.n218 B.n98 71.676
R887 B.n222 B.n99 71.676
R888 B.n227 B.n100 71.676
R889 B.n231 B.n101 71.676
R890 B.n235 B.n102 71.676
R891 B.n239 B.n103 71.676
R892 B.n243 B.n104 71.676
R893 B.n247 B.n105 71.676
R894 B.n251 B.n106 71.676
R895 B.n255 B.n107 71.676
R896 B.n259 B.n108 71.676
R897 B.n263 B.n109 71.676
R898 B.n267 B.n110 71.676
R899 B.n271 B.n111 71.676
R900 B.n275 B.n112 71.676
R901 B.n279 B.n113 71.676
R902 B.n283 B.n114 71.676
R903 B.n287 B.n115 71.676
R904 B.n291 B.n116 71.676
R905 B.n295 B.n117 71.676
R906 B.n299 B.n118 71.676
R907 B.n785 B.n119 71.676
R908 B.n785 B.n784 71.676
R909 B.n301 B.n118 71.676
R910 B.n298 B.n117 71.676
R911 B.n294 B.n116 71.676
R912 B.n290 B.n115 71.676
R913 B.n286 B.n114 71.676
R914 B.n282 B.n113 71.676
R915 B.n278 B.n112 71.676
R916 B.n274 B.n111 71.676
R917 B.n270 B.n110 71.676
R918 B.n266 B.n109 71.676
R919 B.n262 B.n108 71.676
R920 B.n258 B.n107 71.676
R921 B.n254 B.n106 71.676
R922 B.n250 B.n105 71.676
R923 B.n246 B.n104 71.676
R924 B.n242 B.n103 71.676
R925 B.n238 B.n102 71.676
R926 B.n234 B.n101 71.676
R927 B.n230 B.n100 71.676
R928 B.n226 B.n99 71.676
R929 B.n221 B.n98 71.676
R930 B.n217 B.n97 71.676
R931 B.n213 B.n96 71.676
R932 B.n209 B.n95 71.676
R933 B.n205 B.n94 71.676
R934 B.n200 B.n93 71.676
R935 B.n196 B.n92 71.676
R936 B.n192 B.n91 71.676
R937 B.n188 B.n90 71.676
R938 B.n184 B.n89 71.676
R939 B.n180 B.n88 71.676
R940 B.n176 B.n87 71.676
R941 B.n172 B.n86 71.676
R942 B.n168 B.n85 71.676
R943 B.n164 B.n84 71.676
R944 B.n160 B.n83 71.676
R945 B.n156 B.n82 71.676
R946 B.n152 B.n81 71.676
R947 B.n148 B.n80 71.676
R948 B.n144 B.n79 71.676
R949 B.n140 B.n78 71.676
R950 B.n136 B.n77 71.676
R951 B.n132 B.n76 71.676
R952 B.n128 B.n75 71.676
R953 B.n787 B.n74 71.676
R954 B.n612 B.n611 71.676
R955 B.n425 B.n380 71.676
R956 B.n604 B.n381 71.676
R957 B.n600 B.n382 71.676
R958 B.n596 B.n383 71.676
R959 B.n592 B.n384 71.676
R960 B.n588 B.n385 71.676
R961 B.n584 B.n386 71.676
R962 B.n580 B.n387 71.676
R963 B.n576 B.n388 71.676
R964 B.n572 B.n389 71.676
R965 B.n568 B.n390 71.676
R966 B.n564 B.n391 71.676
R967 B.n560 B.n392 71.676
R968 B.n556 B.n393 71.676
R969 B.n552 B.n394 71.676
R970 B.n548 B.n395 71.676
R971 B.n544 B.n396 71.676
R972 B.n540 B.n397 71.676
R973 B.n536 B.n398 71.676
R974 B.n532 B.n399 71.676
R975 B.n528 B.n400 71.676
R976 B.n524 B.n401 71.676
R977 B.n520 B.n402 71.676
R978 B.n516 B.n403 71.676
R979 B.n512 B.n404 71.676
R980 B.n508 B.n405 71.676
R981 B.n504 B.n406 71.676
R982 B.n500 B.n407 71.676
R983 B.n496 B.n408 71.676
R984 B.n492 B.n409 71.676
R985 B.n488 B.n410 71.676
R986 B.n484 B.n411 71.676
R987 B.n480 B.n412 71.676
R988 B.n476 B.n413 71.676
R989 B.n472 B.n414 71.676
R990 B.n468 B.n415 71.676
R991 B.n464 B.n416 71.676
R992 B.n460 B.n417 71.676
R993 B.n456 B.n418 71.676
R994 B.n452 B.n419 71.676
R995 B.n448 B.n420 71.676
R996 B.n444 B.n421 71.676
R997 B.n440 B.n422 71.676
R998 B.n436 B.n423 71.676
R999 B.n611 B.n379 71.676
R1000 B.n605 B.n380 71.676
R1001 B.n601 B.n381 71.676
R1002 B.n597 B.n382 71.676
R1003 B.n593 B.n383 71.676
R1004 B.n589 B.n384 71.676
R1005 B.n585 B.n385 71.676
R1006 B.n581 B.n386 71.676
R1007 B.n577 B.n387 71.676
R1008 B.n573 B.n388 71.676
R1009 B.n569 B.n389 71.676
R1010 B.n565 B.n390 71.676
R1011 B.n561 B.n391 71.676
R1012 B.n557 B.n392 71.676
R1013 B.n553 B.n393 71.676
R1014 B.n549 B.n394 71.676
R1015 B.n545 B.n395 71.676
R1016 B.n541 B.n396 71.676
R1017 B.n537 B.n397 71.676
R1018 B.n533 B.n398 71.676
R1019 B.n529 B.n399 71.676
R1020 B.n525 B.n400 71.676
R1021 B.n521 B.n401 71.676
R1022 B.n517 B.n402 71.676
R1023 B.n513 B.n403 71.676
R1024 B.n509 B.n404 71.676
R1025 B.n505 B.n405 71.676
R1026 B.n501 B.n406 71.676
R1027 B.n497 B.n407 71.676
R1028 B.n493 B.n408 71.676
R1029 B.n489 B.n409 71.676
R1030 B.n485 B.n410 71.676
R1031 B.n481 B.n411 71.676
R1032 B.n477 B.n412 71.676
R1033 B.n473 B.n413 71.676
R1034 B.n469 B.n414 71.676
R1035 B.n465 B.n415 71.676
R1036 B.n461 B.n416 71.676
R1037 B.n457 B.n417 71.676
R1038 B.n453 B.n418 71.676
R1039 B.n449 B.n419 71.676
R1040 B.n445 B.n420 71.676
R1041 B.n441 B.n421 71.676
R1042 B.n437 B.n422 71.676
R1043 B.n433 B.n423 71.676
R1044 B.n869 B.n868 71.676
R1045 B.n869 B.n2 71.676
R1046 B.n203 B.n124 59.5399
R1047 B.n224 B.n122 59.5399
R1048 B.n431 B.n430 59.5399
R1049 B.n428 B.n427 59.5399
R1050 B.n617 B.n376 43.7816
R1051 B.n617 B.n372 43.7816
R1052 B.n623 B.n372 43.7816
R1053 B.n623 B.n368 43.7816
R1054 B.n629 B.n368 43.7816
R1055 B.n635 B.n364 43.7816
R1056 B.n635 B.n360 43.7816
R1057 B.n641 B.n360 43.7816
R1058 B.n641 B.n356 43.7816
R1059 B.n647 B.n356 43.7816
R1060 B.n647 B.n351 43.7816
R1061 B.n653 B.n351 43.7816
R1062 B.n653 B.n352 43.7816
R1063 B.n659 B.n344 43.7816
R1064 B.n665 B.n344 43.7816
R1065 B.n665 B.n340 43.7816
R1066 B.n671 B.n340 43.7816
R1067 B.n677 B.n336 43.7816
R1068 B.n677 B.n332 43.7816
R1069 B.n684 B.n332 43.7816
R1070 B.n684 B.n683 43.7816
R1071 B.n690 B.n325 43.7816
R1072 B.n696 B.n325 43.7816
R1073 B.n696 B.n321 43.7816
R1074 B.n702 B.n321 43.7816
R1075 B.n702 B.t3 43.7816
R1076 B.n708 B.t3 43.7816
R1077 B.n708 B.n314 43.7816
R1078 B.n714 B.n314 43.7816
R1079 B.n714 B.n310 43.7816
R1080 B.n721 B.n310 43.7816
R1081 B.n727 B.n306 43.7816
R1082 B.n727 B.n4 43.7816
R1083 B.n867 B.n4 43.7816
R1084 B.n867 B.n866 43.7816
R1085 B.n866 B.n865 43.7816
R1086 B.n865 B.n8 43.7816
R1087 B.n736 B.n8 43.7816
R1088 B.n858 B.n857 43.7816
R1089 B.n857 B.n856 43.7816
R1090 B.n856 B.n15 43.7816
R1091 B.n850 B.n15 43.7816
R1092 B.n850 B.t2 43.7816
R1093 B.t2 B.n849 43.7816
R1094 B.n849 B.n22 43.7816
R1095 B.n843 B.n22 43.7816
R1096 B.n843 B.n842 43.7816
R1097 B.n842 B.n841 43.7816
R1098 B.n835 B.n32 43.7816
R1099 B.n835 B.n834 43.7816
R1100 B.n834 B.n833 43.7816
R1101 B.n833 B.n36 43.7816
R1102 B.n827 B.n826 43.7816
R1103 B.n826 B.n825 43.7816
R1104 B.n825 B.n43 43.7816
R1105 B.n819 B.n43 43.7816
R1106 B.n818 B.n817 43.7816
R1107 B.n817 B.n50 43.7816
R1108 B.n811 B.n50 43.7816
R1109 B.n811 B.n810 43.7816
R1110 B.n810 B.n809 43.7816
R1111 B.n809 B.n57 43.7816
R1112 B.n803 B.n57 43.7816
R1113 B.n803 B.n802 43.7816
R1114 B.n801 B.n64 43.7816
R1115 B.n795 B.n64 43.7816
R1116 B.n795 B.n794 43.7816
R1117 B.n794 B.n793 43.7816
R1118 B.n793 B.n71 43.7816
R1119 B.n659 B.t9 34.7678
R1120 B.n819 B.t4 34.7678
R1121 B.n124 B.n123 34.7157
R1122 B.n122 B.n121 34.7157
R1123 B.n430 B.n429 34.7157
R1124 B.n427 B.n426 34.7157
R1125 B.n614 B.n613 32.9371
R1126 B.n432 B.n374 32.9371
R1127 B.n783 B.n782 32.9371
R1128 B.n790 B.n789 32.9371
R1129 B.n629 B.t11 32.1925
R1130 B.n683 B.t1 32.1925
R1131 B.t7 B.n306 32.1925
R1132 B.n736 B.t8 32.1925
R1133 B.n32 B.t6 32.1925
R1134 B.t15 B.n801 32.1925
R1135 B.t0 B.n336 23.1787
R1136 B.t5 B.n36 23.1787
R1137 B.n671 B.t0 20.6034
R1138 B.n827 B.t5 20.6034
R1139 B B.n870 18.0485
R1140 B.t11 B.n364 11.5896
R1141 B.n690 B.t1 11.5896
R1142 B.n721 B.t7 11.5896
R1143 B.n858 B.t8 11.5896
R1144 B.n841 B.t6 11.5896
R1145 B.n802 B.t15 11.5896
R1146 B.n615 B.n614 10.6151
R1147 B.n615 B.n370 10.6151
R1148 B.n625 B.n370 10.6151
R1149 B.n626 B.n625 10.6151
R1150 B.n627 B.n626 10.6151
R1151 B.n627 B.n362 10.6151
R1152 B.n637 B.n362 10.6151
R1153 B.n638 B.n637 10.6151
R1154 B.n639 B.n638 10.6151
R1155 B.n639 B.n354 10.6151
R1156 B.n649 B.n354 10.6151
R1157 B.n650 B.n649 10.6151
R1158 B.n651 B.n650 10.6151
R1159 B.n651 B.n346 10.6151
R1160 B.n661 B.n346 10.6151
R1161 B.n662 B.n661 10.6151
R1162 B.n663 B.n662 10.6151
R1163 B.n663 B.n338 10.6151
R1164 B.n673 B.n338 10.6151
R1165 B.n674 B.n673 10.6151
R1166 B.n675 B.n674 10.6151
R1167 B.n675 B.n330 10.6151
R1168 B.n686 B.n330 10.6151
R1169 B.n687 B.n686 10.6151
R1170 B.n688 B.n687 10.6151
R1171 B.n688 B.n323 10.6151
R1172 B.n698 B.n323 10.6151
R1173 B.n699 B.n698 10.6151
R1174 B.n700 B.n699 10.6151
R1175 B.n700 B.n316 10.6151
R1176 B.n710 B.n316 10.6151
R1177 B.n711 B.n710 10.6151
R1178 B.n712 B.n711 10.6151
R1179 B.n712 B.n308 10.6151
R1180 B.n723 B.n308 10.6151
R1181 B.n724 B.n723 10.6151
R1182 B.n725 B.n724 10.6151
R1183 B.n725 B.n0 10.6151
R1184 B.n613 B.n378 10.6151
R1185 B.n608 B.n378 10.6151
R1186 B.n608 B.n607 10.6151
R1187 B.n607 B.n606 10.6151
R1188 B.n606 B.n603 10.6151
R1189 B.n603 B.n602 10.6151
R1190 B.n602 B.n599 10.6151
R1191 B.n599 B.n598 10.6151
R1192 B.n598 B.n595 10.6151
R1193 B.n595 B.n594 10.6151
R1194 B.n594 B.n591 10.6151
R1195 B.n591 B.n590 10.6151
R1196 B.n590 B.n587 10.6151
R1197 B.n587 B.n586 10.6151
R1198 B.n586 B.n583 10.6151
R1199 B.n583 B.n582 10.6151
R1200 B.n582 B.n579 10.6151
R1201 B.n579 B.n578 10.6151
R1202 B.n578 B.n575 10.6151
R1203 B.n575 B.n574 10.6151
R1204 B.n574 B.n571 10.6151
R1205 B.n571 B.n570 10.6151
R1206 B.n570 B.n567 10.6151
R1207 B.n567 B.n566 10.6151
R1208 B.n566 B.n563 10.6151
R1209 B.n563 B.n562 10.6151
R1210 B.n562 B.n559 10.6151
R1211 B.n559 B.n558 10.6151
R1212 B.n558 B.n555 10.6151
R1213 B.n555 B.n554 10.6151
R1214 B.n554 B.n551 10.6151
R1215 B.n551 B.n550 10.6151
R1216 B.n550 B.n547 10.6151
R1217 B.n547 B.n546 10.6151
R1218 B.n546 B.n543 10.6151
R1219 B.n543 B.n542 10.6151
R1220 B.n542 B.n539 10.6151
R1221 B.n539 B.n538 10.6151
R1222 B.n538 B.n535 10.6151
R1223 B.n535 B.n534 10.6151
R1224 B.n531 B.n530 10.6151
R1225 B.n530 B.n527 10.6151
R1226 B.n527 B.n526 10.6151
R1227 B.n526 B.n523 10.6151
R1228 B.n523 B.n522 10.6151
R1229 B.n522 B.n519 10.6151
R1230 B.n519 B.n518 10.6151
R1231 B.n518 B.n515 10.6151
R1232 B.n515 B.n514 10.6151
R1233 B.n511 B.n510 10.6151
R1234 B.n510 B.n507 10.6151
R1235 B.n507 B.n506 10.6151
R1236 B.n506 B.n503 10.6151
R1237 B.n503 B.n502 10.6151
R1238 B.n502 B.n499 10.6151
R1239 B.n499 B.n498 10.6151
R1240 B.n498 B.n495 10.6151
R1241 B.n495 B.n494 10.6151
R1242 B.n494 B.n491 10.6151
R1243 B.n491 B.n490 10.6151
R1244 B.n490 B.n487 10.6151
R1245 B.n487 B.n486 10.6151
R1246 B.n486 B.n483 10.6151
R1247 B.n483 B.n482 10.6151
R1248 B.n482 B.n479 10.6151
R1249 B.n479 B.n478 10.6151
R1250 B.n478 B.n475 10.6151
R1251 B.n475 B.n474 10.6151
R1252 B.n474 B.n471 10.6151
R1253 B.n471 B.n470 10.6151
R1254 B.n470 B.n467 10.6151
R1255 B.n467 B.n466 10.6151
R1256 B.n466 B.n463 10.6151
R1257 B.n463 B.n462 10.6151
R1258 B.n462 B.n459 10.6151
R1259 B.n459 B.n458 10.6151
R1260 B.n458 B.n455 10.6151
R1261 B.n455 B.n454 10.6151
R1262 B.n454 B.n451 10.6151
R1263 B.n451 B.n450 10.6151
R1264 B.n450 B.n447 10.6151
R1265 B.n447 B.n446 10.6151
R1266 B.n446 B.n443 10.6151
R1267 B.n443 B.n442 10.6151
R1268 B.n442 B.n439 10.6151
R1269 B.n439 B.n438 10.6151
R1270 B.n438 B.n435 10.6151
R1271 B.n435 B.n434 10.6151
R1272 B.n434 B.n432 10.6151
R1273 B.n619 B.n374 10.6151
R1274 B.n620 B.n619 10.6151
R1275 B.n621 B.n620 10.6151
R1276 B.n621 B.n366 10.6151
R1277 B.n631 B.n366 10.6151
R1278 B.n632 B.n631 10.6151
R1279 B.n633 B.n632 10.6151
R1280 B.n633 B.n358 10.6151
R1281 B.n643 B.n358 10.6151
R1282 B.n644 B.n643 10.6151
R1283 B.n645 B.n644 10.6151
R1284 B.n645 B.n349 10.6151
R1285 B.n655 B.n349 10.6151
R1286 B.n656 B.n655 10.6151
R1287 B.n657 B.n656 10.6151
R1288 B.n657 B.n342 10.6151
R1289 B.n667 B.n342 10.6151
R1290 B.n668 B.n667 10.6151
R1291 B.n669 B.n668 10.6151
R1292 B.n669 B.n334 10.6151
R1293 B.n679 B.n334 10.6151
R1294 B.n680 B.n679 10.6151
R1295 B.n681 B.n680 10.6151
R1296 B.n681 B.n327 10.6151
R1297 B.n692 B.n327 10.6151
R1298 B.n693 B.n692 10.6151
R1299 B.n694 B.n693 10.6151
R1300 B.n694 B.n319 10.6151
R1301 B.n704 B.n319 10.6151
R1302 B.n705 B.n704 10.6151
R1303 B.n706 B.n705 10.6151
R1304 B.n706 B.n312 10.6151
R1305 B.n716 B.n312 10.6151
R1306 B.n717 B.n716 10.6151
R1307 B.n719 B.n717 10.6151
R1308 B.n719 B.n718 10.6151
R1309 B.n718 B.n304 10.6151
R1310 B.n730 B.n304 10.6151
R1311 B.n731 B.n730 10.6151
R1312 B.n732 B.n731 10.6151
R1313 B.n733 B.n732 10.6151
R1314 B.n734 B.n733 10.6151
R1315 B.n738 B.n734 10.6151
R1316 B.n739 B.n738 10.6151
R1317 B.n740 B.n739 10.6151
R1318 B.n741 B.n740 10.6151
R1319 B.n743 B.n741 10.6151
R1320 B.n744 B.n743 10.6151
R1321 B.n745 B.n744 10.6151
R1322 B.n746 B.n745 10.6151
R1323 B.n748 B.n746 10.6151
R1324 B.n749 B.n748 10.6151
R1325 B.n750 B.n749 10.6151
R1326 B.n751 B.n750 10.6151
R1327 B.n753 B.n751 10.6151
R1328 B.n754 B.n753 10.6151
R1329 B.n755 B.n754 10.6151
R1330 B.n756 B.n755 10.6151
R1331 B.n758 B.n756 10.6151
R1332 B.n759 B.n758 10.6151
R1333 B.n760 B.n759 10.6151
R1334 B.n761 B.n760 10.6151
R1335 B.n763 B.n761 10.6151
R1336 B.n764 B.n763 10.6151
R1337 B.n765 B.n764 10.6151
R1338 B.n766 B.n765 10.6151
R1339 B.n768 B.n766 10.6151
R1340 B.n769 B.n768 10.6151
R1341 B.n770 B.n769 10.6151
R1342 B.n771 B.n770 10.6151
R1343 B.n773 B.n771 10.6151
R1344 B.n774 B.n773 10.6151
R1345 B.n775 B.n774 10.6151
R1346 B.n776 B.n775 10.6151
R1347 B.n778 B.n776 10.6151
R1348 B.n779 B.n778 10.6151
R1349 B.n780 B.n779 10.6151
R1350 B.n781 B.n780 10.6151
R1351 B.n782 B.n781 10.6151
R1352 B.n862 B.n1 10.6151
R1353 B.n862 B.n861 10.6151
R1354 B.n861 B.n860 10.6151
R1355 B.n860 B.n10 10.6151
R1356 B.n854 B.n10 10.6151
R1357 B.n854 B.n853 10.6151
R1358 B.n853 B.n852 10.6151
R1359 B.n852 B.n17 10.6151
R1360 B.n847 B.n17 10.6151
R1361 B.n847 B.n846 10.6151
R1362 B.n846 B.n845 10.6151
R1363 B.n845 B.n24 10.6151
R1364 B.n839 B.n24 10.6151
R1365 B.n839 B.n838 10.6151
R1366 B.n838 B.n837 10.6151
R1367 B.n837 B.n30 10.6151
R1368 B.n831 B.n30 10.6151
R1369 B.n831 B.n830 10.6151
R1370 B.n830 B.n829 10.6151
R1371 B.n829 B.n38 10.6151
R1372 B.n823 B.n38 10.6151
R1373 B.n823 B.n822 10.6151
R1374 B.n822 B.n821 10.6151
R1375 B.n821 B.n45 10.6151
R1376 B.n815 B.n45 10.6151
R1377 B.n815 B.n814 10.6151
R1378 B.n814 B.n813 10.6151
R1379 B.n813 B.n52 10.6151
R1380 B.n807 B.n52 10.6151
R1381 B.n807 B.n806 10.6151
R1382 B.n806 B.n805 10.6151
R1383 B.n805 B.n59 10.6151
R1384 B.n799 B.n59 10.6151
R1385 B.n799 B.n798 10.6151
R1386 B.n798 B.n797 10.6151
R1387 B.n797 B.n66 10.6151
R1388 B.n791 B.n66 10.6151
R1389 B.n791 B.n790 10.6151
R1390 B.n789 B.n73 10.6151
R1391 B.n126 B.n73 10.6151
R1392 B.n127 B.n126 10.6151
R1393 B.n130 B.n127 10.6151
R1394 B.n131 B.n130 10.6151
R1395 B.n134 B.n131 10.6151
R1396 B.n135 B.n134 10.6151
R1397 B.n138 B.n135 10.6151
R1398 B.n139 B.n138 10.6151
R1399 B.n142 B.n139 10.6151
R1400 B.n143 B.n142 10.6151
R1401 B.n146 B.n143 10.6151
R1402 B.n147 B.n146 10.6151
R1403 B.n150 B.n147 10.6151
R1404 B.n151 B.n150 10.6151
R1405 B.n154 B.n151 10.6151
R1406 B.n155 B.n154 10.6151
R1407 B.n158 B.n155 10.6151
R1408 B.n159 B.n158 10.6151
R1409 B.n162 B.n159 10.6151
R1410 B.n163 B.n162 10.6151
R1411 B.n166 B.n163 10.6151
R1412 B.n167 B.n166 10.6151
R1413 B.n170 B.n167 10.6151
R1414 B.n171 B.n170 10.6151
R1415 B.n174 B.n171 10.6151
R1416 B.n175 B.n174 10.6151
R1417 B.n178 B.n175 10.6151
R1418 B.n179 B.n178 10.6151
R1419 B.n182 B.n179 10.6151
R1420 B.n183 B.n182 10.6151
R1421 B.n186 B.n183 10.6151
R1422 B.n187 B.n186 10.6151
R1423 B.n190 B.n187 10.6151
R1424 B.n191 B.n190 10.6151
R1425 B.n194 B.n191 10.6151
R1426 B.n195 B.n194 10.6151
R1427 B.n198 B.n195 10.6151
R1428 B.n199 B.n198 10.6151
R1429 B.n202 B.n199 10.6151
R1430 B.n207 B.n204 10.6151
R1431 B.n208 B.n207 10.6151
R1432 B.n211 B.n208 10.6151
R1433 B.n212 B.n211 10.6151
R1434 B.n215 B.n212 10.6151
R1435 B.n216 B.n215 10.6151
R1436 B.n219 B.n216 10.6151
R1437 B.n220 B.n219 10.6151
R1438 B.n223 B.n220 10.6151
R1439 B.n228 B.n225 10.6151
R1440 B.n229 B.n228 10.6151
R1441 B.n232 B.n229 10.6151
R1442 B.n233 B.n232 10.6151
R1443 B.n236 B.n233 10.6151
R1444 B.n237 B.n236 10.6151
R1445 B.n240 B.n237 10.6151
R1446 B.n241 B.n240 10.6151
R1447 B.n244 B.n241 10.6151
R1448 B.n245 B.n244 10.6151
R1449 B.n248 B.n245 10.6151
R1450 B.n249 B.n248 10.6151
R1451 B.n252 B.n249 10.6151
R1452 B.n253 B.n252 10.6151
R1453 B.n256 B.n253 10.6151
R1454 B.n257 B.n256 10.6151
R1455 B.n260 B.n257 10.6151
R1456 B.n261 B.n260 10.6151
R1457 B.n264 B.n261 10.6151
R1458 B.n265 B.n264 10.6151
R1459 B.n268 B.n265 10.6151
R1460 B.n269 B.n268 10.6151
R1461 B.n272 B.n269 10.6151
R1462 B.n273 B.n272 10.6151
R1463 B.n276 B.n273 10.6151
R1464 B.n277 B.n276 10.6151
R1465 B.n280 B.n277 10.6151
R1466 B.n281 B.n280 10.6151
R1467 B.n284 B.n281 10.6151
R1468 B.n285 B.n284 10.6151
R1469 B.n288 B.n285 10.6151
R1470 B.n289 B.n288 10.6151
R1471 B.n292 B.n289 10.6151
R1472 B.n293 B.n292 10.6151
R1473 B.n296 B.n293 10.6151
R1474 B.n297 B.n296 10.6151
R1475 B.n300 B.n297 10.6151
R1476 B.n302 B.n300 10.6151
R1477 B.n303 B.n302 10.6151
R1478 B.n783 B.n303 10.6151
R1479 B.n534 B.n428 9.36635
R1480 B.n511 B.n431 9.36635
R1481 B.n203 B.n202 9.36635
R1482 B.n225 B.n224 9.36635
R1483 B.n352 B.t9 9.01425
R1484 B.t4 B.n818 9.01425
R1485 B.n870 B.n0 8.11757
R1486 B.n870 B.n1 8.11757
R1487 B.n531 B.n428 1.24928
R1488 B.n514 B.n431 1.24928
R1489 B.n204 B.n203 1.24928
R1490 B.n224 B.n223 1.24928
R1491 VN.n7 VN.t4 225.363
R1492 VN.n34 VN.t5 225.363
R1493 VN.n12 VN.t6 194.946
R1494 VN.n6 VN.t2 194.946
R1495 VN.n18 VN.t9 194.946
R1496 VN.n25 VN.t7 194.946
R1497 VN.n39 VN.t3 194.946
R1498 VN.n33 VN.t0 194.946
R1499 VN.n45 VN.t8 194.946
R1500 VN.n52 VN.t1 194.946
R1501 VN.n26 VN.n25 181.852
R1502 VN.n53 VN.n52 181.852
R1503 VN.n51 VN.n27 161.3
R1504 VN.n50 VN.n49 161.3
R1505 VN.n48 VN.n28 161.3
R1506 VN.n47 VN.n46 161.3
R1507 VN.n44 VN.n29 161.3
R1508 VN.n43 VN.n42 161.3
R1509 VN.n41 VN.n30 161.3
R1510 VN.n40 VN.n39 161.3
R1511 VN.n38 VN.n31 161.3
R1512 VN.n37 VN.n36 161.3
R1513 VN.n35 VN.n32 161.3
R1514 VN.n24 VN.n0 161.3
R1515 VN.n23 VN.n22 161.3
R1516 VN.n21 VN.n1 161.3
R1517 VN.n20 VN.n19 161.3
R1518 VN.n17 VN.n2 161.3
R1519 VN.n16 VN.n15 161.3
R1520 VN.n14 VN.n3 161.3
R1521 VN.n13 VN.n12 161.3
R1522 VN.n11 VN.n4 161.3
R1523 VN.n10 VN.n9 161.3
R1524 VN.n8 VN.n5 161.3
R1525 VN.n23 VN.n1 56.5193
R1526 VN.n50 VN.n28 56.5193
R1527 VN.n7 VN.n6 51.5804
R1528 VN.n34 VN.n33 51.5804
R1529 VN.n11 VN.n10 50.6917
R1530 VN.n16 VN.n3 50.6917
R1531 VN.n38 VN.n37 50.6917
R1532 VN.n43 VN.n30 50.6917
R1533 VN VN.n53 46.9759
R1534 VN.n10 VN.n5 30.2951
R1535 VN.n17 VN.n16 30.2951
R1536 VN.n37 VN.n32 30.2951
R1537 VN.n44 VN.n43 30.2951
R1538 VN.n12 VN.n11 24.4675
R1539 VN.n12 VN.n3 24.4675
R1540 VN.n19 VN.n1 24.4675
R1541 VN.n24 VN.n23 24.4675
R1542 VN.n39 VN.n30 24.4675
R1543 VN.n39 VN.n38 24.4675
R1544 VN.n46 VN.n28 24.4675
R1545 VN.n51 VN.n50 24.4675
R1546 VN.n35 VN.n34 18.3855
R1547 VN.n8 VN.n7 18.3855
R1548 VN.n6 VN.n5 14.1914
R1549 VN.n18 VN.n17 14.1914
R1550 VN.n33 VN.n32 14.1914
R1551 VN.n45 VN.n44 14.1914
R1552 VN.n19 VN.n18 10.2766
R1553 VN.n46 VN.n45 10.2766
R1554 VN.n25 VN.n24 3.91522
R1555 VN.n52 VN.n51 3.91522
R1556 VN.n53 VN.n27 0.189894
R1557 VN.n49 VN.n27 0.189894
R1558 VN.n49 VN.n48 0.189894
R1559 VN.n48 VN.n47 0.189894
R1560 VN.n47 VN.n29 0.189894
R1561 VN.n42 VN.n29 0.189894
R1562 VN.n42 VN.n41 0.189894
R1563 VN.n41 VN.n40 0.189894
R1564 VN.n40 VN.n31 0.189894
R1565 VN.n36 VN.n31 0.189894
R1566 VN.n36 VN.n35 0.189894
R1567 VN.n9 VN.n8 0.189894
R1568 VN.n9 VN.n4 0.189894
R1569 VN.n13 VN.n4 0.189894
R1570 VN.n14 VN.n13 0.189894
R1571 VN.n15 VN.n14 0.189894
R1572 VN.n15 VN.n2 0.189894
R1573 VN.n20 VN.n2 0.189894
R1574 VN.n21 VN.n20 0.189894
R1575 VN.n22 VN.n21 0.189894
R1576 VN.n22 VN.n0 0.189894
R1577 VN.n26 VN.n0 0.189894
R1578 VN VN.n26 0.0516364
R1579 VDD2.n1 VDD2.t0 66.1691
R1580 VDD2.n4 VDD2.t4 64.6263
R1581 VDD2.n3 VDD2.n2 64.0515
R1582 VDD2 VDD2.n7 64.0487
R1583 VDD2.n6 VDD2.n5 62.9497
R1584 VDD2.n1 VDD2.n0 62.9495
R1585 VDD2.n4 VDD2.n3 41.2261
R1586 VDD2.n7 VDD2.t2 1.67705
R1587 VDD2.n7 VDD2.t3 1.67705
R1588 VDD2.n5 VDD2.t6 1.67705
R1589 VDD2.n5 VDD2.t9 1.67705
R1590 VDD2.n2 VDD2.t5 1.67705
R1591 VDD2.n2 VDD2.t8 1.67705
R1592 VDD2.n0 VDD2.t1 1.67705
R1593 VDD2.n0 VDD2.t7 1.67705
R1594 VDD2.n6 VDD2.n4 1.5436
R1595 VDD2 VDD2.n6 0.444466
R1596 VDD2.n3 VDD2.n1 0.33093
R1597 VTAIL.n11 VTAIL.t14 47.9475
R1598 VTAIL.n17 VTAIL.t12 47.9473
R1599 VTAIL.n2 VTAIL.t6 47.9473
R1600 VTAIL.n16 VTAIL.t0 47.9473
R1601 VTAIL.n15 VTAIL.n14 46.2709
R1602 VTAIL.n13 VTAIL.n12 46.2709
R1603 VTAIL.n10 VTAIL.n9 46.2709
R1604 VTAIL.n8 VTAIL.n7 46.2709
R1605 VTAIL.n19 VTAIL.n18 46.2707
R1606 VTAIL.n1 VTAIL.n0 46.2707
R1607 VTAIL.n4 VTAIL.n3 46.2707
R1608 VTAIL.n6 VTAIL.n5 46.2707
R1609 VTAIL.n8 VTAIL.n6 25.6341
R1610 VTAIL.n17 VTAIL.n16 24.091
R1611 VTAIL.n18 VTAIL.t13 1.67705
R1612 VTAIL.n18 VTAIL.t10 1.67705
R1613 VTAIL.n0 VTAIL.t15 1.67705
R1614 VTAIL.n0 VTAIL.t17 1.67705
R1615 VTAIL.n3 VTAIL.t3 1.67705
R1616 VTAIL.n3 VTAIL.t4 1.67705
R1617 VTAIL.n5 VTAIL.t9 1.67705
R1618 VTAIL.n5 VTAIL.t2 1.67705
R1619 VTAIL.n14 VTAIL.t5 1.67705
R1620 VTAIL.n14 VTAIL.t1 1.67705
R1621 VTAIL.n12 VTAIL.t7 1.67705
R1622 VTAIL.n12 VTAIL.t8 1.67705
R1623 VTAIL.n9 VTAIL.t16 1.67705
R1624 VTAIL.n9 VTAIL.t19 1.67705
R1625 VTAIL.n7 VTAIL.t18 1.67705
R1626 VTAIL.n7 VTAIL.t11 1.67705
R1627 VTAIL.n10 VTAIL.n8 1.5436
R1628 VTAIL.n11 VTAIL.n10 1.5436
R1629 VTAIL.n15 VTAIL.n13 1.5436
R1630 VTAIL.n16 VTAIL.n15 1.5436
R1631 VTAIL.n6 VTAIL.n4 1.5436
R1632 VTAIL.n4 VTAIL.n2 1.5436
R1633 VTAIL.n19 VTAIL.n17 1.5436
R1634 VTAIL.n13 VTAIL.n11 1.24188
R1635 VTAIL.n2 VTAIL.n1 1.24188
R1636 VTAIL VTAIL.n1 1.21602
R1637 VTAIL VTAIL.n19 0.328086
R1638 VP.n15 VP.t2 225.363
R1639 VP.n48 VP.t0 194.946
R1640 VP.n35 VP.t9 194.946
R1641 VP.n41 VP.t1 194.946
R1642 VP.n54 VP.t8 194.946
R1643 VP.n61 VP.t6 194.946
R1644 VP.n20 VP.t7 194.946
R1645 VP.n33 VP.t5 194.946
R1646 VP.n26 VP.t3 194.946
R1647 VP.n14 VP.t4 194.946
R1648 VP.n36 VP.n35 181.852
R1649 VP.n62 VP.n61 181.852
R1650 VP.n34 VP.n33 181.852
R1651 VP.n16 VP.n13 161.3
R1652 VP.n18 VP.n17 161.3
R1653 VP.n19 VP.n12 161.3
R1654 VP.n21 VP.n20 161.3
R1655 VP.n22 VP.n11 161.3
R1656 VP.n24 VP.n23 161.3
R1657 VP.n25 VP.n10 161.3
R1658 VP.n28 VP.n27 161.3
R1659 VP.n29 VP.n9 161.3
R1660 VP.n31 VP.n30 161.3
R1661 VP.n32 VP.n8 161.3
R1662 VP.n60 VP.n0 161.3
R1663 VP.n59 VP.n58 161.3
R1664 VP.n57 VP.n1 161.3
R1665 VP.n56 VP.n55 161.3
R1666 VP.n53 VP.n2 161.3
R1667 VP.n52 VP.n51 161.3
R1668 VP.n50 VP.n3 161.3
R1669 VP.n49 VP.n48 161.3
R1670 VP.n47 VP.n4 161.3
R1671 VP.n46 VP.n45 161.3
R1672 VP.n44 VP.n5 161.3
R1673 VP.n43 VP.n42 161.3
R1674 VP.n40 VP.n6 161.3
R1675 VP.n39 VP.n38 161.3
R1676 VP.n37 VP.n7 161.3
R1677 VP.n40 VP.n39 56.5193
R1678 VP.n59 VP.n1 56.5193
R1679 VP.n31 VP.n9 56.5193
R1680 VP.n15 VP.n14 51.5804
R1681 VP.n47 VP.n46 50.6917
R1682 VP.n52 VP.n3 50.6917
R1683 VP.n24 VP.n11 50.6917
R1684 VP.n19 VP.n18 50.6917
R1685 VP.n36 VP.n34 46.5952
R1686 VP.n46 VP.n5 30.2951
R1687 VP.n53 VP.n52 30.2951
R1688 VP.n25 VP.n24 30.2951
R1689 VP.n18 VP.n13 30.2951
R1690 VP.n39 VP.n7 24.4675
R1691 VP.n42 VP.n40 24.4675
R1692 VP.n48 VP.n47 24.4675
R1693 VP.n48 VP.n3 24.4675
R1694 VP.n55 VP.n1 24.4675
R1695 VP.n60 VP.n59 24.4675
R1696 VP.n32 VP.n31 24.4675
R1697 VP.n27 VP.n9 24.4675
R1698 VP.n20 VP.n19 24.4675
R1699 VP.n20 VP.n11 24.4675
R1700 VP.n16 VP.n15 18.3855
R1701 VP.n41 VP.n5 14.1914
R1702 VP.n54 VP.n53 14.1914
R1703 VP.n26 VP.n25 14.1914
R1704 VP.n14 VP.n13 14.1914
R1705 VP.n42 VP.n41 10.2766
R1706 VP.n55 VP.n54 10.2766
R1707 VP.n27 VP.n26 10.2766
R1708 VP.n35 VP.n7 3.91522
R1709 VP.n61 VP.n60 3.91522
R1710 VP.n33 VP.n32 3.91522
R1711 VP.n17 VP.n16 0.189894
R1712 VP.n17 VP.n12 0.189894
R1713 VP.n21 VP.n12 0.189894
R1714 VP.n22 VP.n21 0.189894
R1715 VP.n23 VP.n22 0.189894
R1716 VP.n23 VP.n10 0.189894
R1717 VP.n28 VP.n10 0.189894
R1718 VP.n29 VP.n28 0.189894
R1719 VP.n30 VP.n29 0.189894
R1720 VP.n30 VP.n8 0.189894
R1721 VP.n34 VP.n8 0.189894
R1722 VP.n37 VP.n36 0.189894
R1723 VP.n38 VP.n37 0.189894
R1724 VP.n38 VP.n6 0.189894
R1725 VP.n43 VP.n6 0.189894
R1726 VP.n44 VP.n43 0.189894
R1727 VP.n45 VP.n44 0.189894
R1728 VP.n45 VP.n4 0.189894
R1729 VP.n49 VP.n4 0.189894
R1730 VP.n50 VP.n49 0.189894
R1731 VP.n51 VP.n50 0.189894
R1732 VP.n51 VP.n2 0.189894
R1733 VP.n56 VP.n2 0.189894
R1734 VP.n57 VP.n56 0.189894
R1735 VP.n58 VP.n57 0.189894
R1736 VP.n58 VP.n0 0.189894
R1737 VP.n62 VP.n0 0.189894
R1738 VP VP.n62 0.0516364
R1739 VDD1.n1 VDD1.t7 66.1694
R1740 VDD1.n3 VDD1.t0 66.1691
R1741 VDD1.n5 VDD1.n4 64.0515
R1742 VDD1.n1 VDD1.n0 62.9497
R1743 VDD1.n7 VDD1.n6 62.9495
R1744 VDD1.n3 VDD1.n2 62.9495
R1745 VDD1.n7 VDD1.n5 42.5806
R1746 VDD1.n6 VDD1.t6 1.67705
R1747 VDD1.n6 VDD1.t4 1.67705
R1748 VDD1.n0 VDD1.t5 1.67705
R1749 VDD1.n0 VDD1.t2 1.67705
R1750 VDD1.n4 VDD1.t1 1.67705
R1751 VDD1.n4 VDD1.t3 1.67705
R1752 VDD1.n2 VDD1.t8 1.67705
R1753 VDD1.n2 VDD1.t9 1.67705
R1754 VDD1 VDD1.n7 1.09964
R1755 VDD1 VDD1.n1 0.444466
R1756 VDD1.n5 VDD1.n3 0.33093
C0 VP VN 6.68707f
C1 VDD2 VN 9.03568f
C2 VN VTAIL 9.210481f
C3 VDD2 VP 0.438278f
C4 VP VTAIL 9.2249f
C5 VDD2 VTAIL 10.9128f
C6 VN VDD1 0.150779f
C7 VP VDD1 9.31913f
C8 VDD2 VDD1 1.43344f
C9 VDD1 VTAIL 10.871201f
C10 VDD2 B 5.841194f
C11 VDD1 B 5.811207f
C12 VTAIL B 7.193978f
C13 VN B 12.80041f
C14 VP B 11.153502f
C15 VDD1.t7 B 2.41751f
C16 VDD1.t5 B 0.212109f
C17 VDD1.t2 B 0.212109f
C18 VDD1.n0 B 1.88896f
C19 VDD1.n1 B 0.691856f
C20 VDD1.t0 B 2.4175f
C21 VDD1.t8 B 0.212109f
C22 VDD1.t9 B 0.212109f
C23 VDD1.n2 B 1.88895f
C24 VDD1.n3 B 0.685144f
C25 VDD1.t1 B 0.212109f
C26 VDD1.t3 B 0.212109f
C27 VDD1.n4 B 1.89567f
C28 VDD1.n5 B 2.17338f
C29 VDD1.t6 B 0.212109f
C30 VDD1.t4 B 0.212109f
C31 VDD1.n6 B 1.88895f
C32 VDD1.n7 B 2.4422f
C33 VP.n0 B 0.030771f
C34 VP.t6 B 1.44493f
C35 VP.n1 B 0.039349f
C36 VP.n2 B 0.030771f
C37 VP.t8 B 1.44493f
C38 VP.n3 B 0.056177f
C39 VP.n4 B 0.030771f
C40 VP.t0 B 1.44493f
C41 VP.n5 B 0.049597f
C42 VP.n6 B 0.030771f
C43 VP.n7 B 0.033566f
C44 VP.n8 B 0.030771f
C45 VP.t5 B 1.44493f
C46 VP.n9 B 0.039349f
C47 VP.n10 B 0.030771f
C48 VP.t3 B 1.44493f
C49 VP.n11 B 0.056177f
C50 VP.n12 B 0.030771f
C51 VP.t7 B 1.44493f
C52 VP.n13 B 0.049597f
C53 VP.t2 B 1.53113f
C54 VP.t4 B 1.44493f
C55 VP.n14 B 0.582169f
C56 VP.n15 B 0.599845f
C57 VP.n16 B 0.190533f
C58 VP.n17 B 0.030771f
C59 VP.n18 B 0.029529f
C60 VP.n19 B 0.056177f
C61 VP.n20 B 0.552983f
C62 VP.n21 B 0.030771f
C63 VP.n22 B 0.030771f
C64 VP.n23 B 0.030771f
C65 VP.n24 B 0.029529f
C66 VP.n25 B 0.049597f
C67 VP.n26 B 0.523947f
C68 VP.n27 B 0.040927f
C69 VP.n28 B 0.030771f
C70 VP.n29 B 0.030771f
C71 VP.n30 B 0.030771f
C72 VP.n31 B 0.050496f
C73 VP.n32 B 0.033566f
C74 VP.n33 B 0.576824f
C75 VP.n34 B 1.50831f
C76 VP.t9 B 1.44493f
C77 VP.n35 B 0.576824f
C78 VP.n36 B 1.53205f
C79 VP.n37 B 0.030771f
C80 VP.n38 B 0.030771f
C81 VP.n39 B 0.050496f
C82 VP.n40 B 0.039349f
C83 VP.t1 B 1.44493f
C84 VP.n41 B 0.523947f
C85 VP.n42 B 0.040927f
C86 VP.n43 B 0.030771f
C87 VP.n44 B 0.030771f
C88 VP.n45 B 0.030771f
C89 VP.n46 B 0.029529f
C90 VP.n47 B 0.056177f
C91 VP.n48 B 0.552983f
C92 VP.n49 B 0.030771f
C93 VP.n50 B 0.030771f
C94 VP.n51 B 0.030771f
C95 VP.n52 B 0.029529f
C96 VP.n53 B 0.049597f
C97 VP.n54 B 0.523947f
C98 VP.n55 B 0.040927f
C99 VP.n56 B 0.030771f
C100 VP.n57 B 0.030771f
C101 VP.n58 B 0.030771f
C102 VP.n59 B 0.050496f
C103 VP.n60 B 0.033566f
C104 VP.n61 B 0.576824f
C105 VP.n62 B 0.030584f
C106 VTAIL.t15 B 0.228496f
C107 VTAIL.t17 B 0.228496f
C108 VTAIL.n0 B 1.96391f
C109 VTAIL.n1 B 0.433115f
C110 VTAIL.t6 B 2.5046f
C111 VTAIL.n2 B 0.541431f
C112 VTAIL.t3 B 0.228496f
C113 VTAIL.t4 B 0.228496f
C114 VTAIL.n3 B 1.96391f
C115 VTAIL.n4 B 0.482762f
C116 VTAIL.t9 B 0.228496f
C117 VTAIL.t2 B 0.228496f
C118 VTAIL.n5 B 1.96391f
C119 VTAIL.n6 B 1.74028f
C120 VTAIL.t18 B 0.228496f
C121 VTAIL.t11 B 0.228496f
C122 VTAIL.n7 B 1.96391f
C123 VTAIL.n8 B 1.74027f
C124 VTAIL.t16 B 0.228496f
C125 VTAIL.t19 B 0.228496f
C126 VTAIL.n9 B 1.96391f
C127 VTAIL.n10 B 0.482756f
C128 VTAIL.t14 B 2.50461f
C129 VTAIL.n11 B 0.541425f
C130 VTAIL.t7 B 0.228496f
C131 VTAIL.t8 B 0.228496f
C132 VTAIL.n12 B 1.96391f
C133 VTAIL.n13 B 0.458953f
C134 VTAIL.t5 B 0.228496f
C135 VTAIL.t1 B 0.228496f
C136 VTAIL.n14 B 1.96391f
C137 VTAIL.n15 B 0.482756f
C138 VTAIL.t0 B 2.5046f
C139 VTAIL.n16 B 1.70101f
C140 VTAIL.t12 B 2.5046f
C141 VTAIL.n17 B 1.70101f
C142 VTAIL.t13 B 0.228496f
C143 VTAIL.t10 B 0.228496f
C144 VTAIL.n18 B 1.96391f
C145 VTAIL.n19 B 0.386868f
C146 VDD2.t0 B 2.39154f
C147 VDD2.t1 B 0.209831f
C148 VDD2.t7 B 0.209831f
C149 VDD2.n0 B 1.86867f
C150 VDD2.n1 B 0.677785f
C151 VDD2.t5 B 0.209831f
C152 VDD2.t8 B 0.209831f
C153 VDD2.n2 B 1.87531f
C154 VDD2.n3 B 2.06429f
C155 VDD2.t4 B 2.38306f
C156 VDD2.n4 B 2.39691f
C157 VDD2.t6 B 0.209831f
C158 VDD2.t9 B 0.209831f
C159 VDD2.n5 B 1.86867f
C160 VDD2.n6 B 0.329069f
C161 VDD2.t2 B 0.209831f
C162 VDD2.t3 B 0.209831f
C163 VDD2.n7 B 1.87528f
C164 VN.n0 B 0.030352f
C165 VN.t7 B 1.42529f
C166 VN.n1 B 0.038814f
C167 VN.n2 B 0.030352f
C168 VN.t9 B 1.42529f
C169 VN.n3 B 0.055413f
C170 VN.n4 B 0.030352f
C171 VN.t6 B 1.42529f
C172 VN.n5 B 0.048922f
C173 VN.t4 B 1.51031f
C174 VN.t2 B 1.42529f
C175 VN.n6 B 0.574253f
C176 VN.n7 B 0.591688f
C177 VN.n8 B 0.187942f
C178 VN.n9 B 0.030352f
C179 VN.n10 B 0.029127f
C180 VN.n11 B 0.055413f
C181 VN.n12 B 0.545463f
C182 VN.n13 B 0.030352f
C183 VN.n14 B 0.030352f
C184 VN.n15 B 0.030352f
C185 VN.n16 B 0.029127f
C186 VN.n17 B 0.048922f
C187 VN.n18 B 0.516823f
C188 VN.n19 B 0.040371f
C189 VN.n20 B 0.030352f
C190 VN.n21 B 0.030352f
C191 VN.n22 B 0.030352f
C192 VN.n23 B 0.049809f
C193 VN.n24 B 0.033109f
C194 VN.n25 B 0.56898f
C195 VN.n26 B 0.030168f
C196 VN.n27 B 0.030352f
C197 VN.t1 B 1.42529f
C198 VN.n28 B 0.038814f
C199 VN.n29 B 0.030352f
C200 VN.t8 B 1.42529f
C201 VN.n30 B 0.055413f
C202 VN.n31 B 0.030352f
C203 VN.t3 B 1.42529f
C204 VN.n32 B 0.048922f
C205 VN.t5 B 1.51031f
C206 VN.t0 B 1.42529f
C207 VN.n33 B 0.574253f
C208 VN.n34 B 0.591688f
C209 VN.n35 B 0.187942f
C210 VN.n36 B 0.030352f
C211 VN.n37 B 0.029127f
C212 VN.n38 B 0.055413f
C213 VN.n39 B 0.545463f
C214 VN.n40 B 0.030352f
C215 VN.n41 B 0.030352f
C216 VN.n42 B 0.030352f
C217 VN.n43 B 0.029127f
C218 VN.n44 B 0.048922f
C219 VN.n45 B 0.516823f
C220 VN.n46 B 0.040371f
C221 VN.n47 B 0.030352f
C222 VN.n48 B 0.030352f
C223 VN.n49 B 0.030352f
C224 VN.n50 B 0.049809f
C225 VN.n51 B 0.033109f
C226 VN.n52 B 0.56898f
C227 VN.n53 B 1.5076f
.ends

