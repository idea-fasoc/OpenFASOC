* NGSPICE file created from diff_pair_sample_1600.ext - technology: sky130A

.subckt diff_pair_sample_1600 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t8 VN.t0 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=1.5972 ps=10.01 w=9.68 l=0.2
X1 VDD2.t0 VN.t1 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=1.5972 ps=10.01 w=9.68 l=0.2
X2 VTAIL.t11 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=1.5972 ps=10.01 w=9.68 l=0.2
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=0 ps=0 w=9.68 l=0.2
X4 VTAIL.t6 VN.t2 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=1.5972 ps=10.01 w=9.68 l=0.2
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=0 ps=0 w=9.68 l=0.2
X6 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=1.5972 ps=10.01 w=9.68 l=0.2
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=0 ps=0 w=9.68 l=0.2
X8 VDD1.t3 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=1.5972 ps=10.01 w=9.68 l=0.2
X9 VDD1.t2 VP.t3 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=3.7752 ps=20.14 w=9.68 l=0.2
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=0 ps=0 w=9.68 l=0.2
X11 VDD2.t4 VN.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=3.7752 ps=20.14 w=9.68 l=0.2
X12 VTAIL.t9 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=1.5972 ps=10.01 w=9.68 l=0.2
X13 VDD2.t3 VN.t4 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=3.7752 ps=20.14 w=9.68 l=0.2
X14 VDD2.t5 VN.t5 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.7752 pd=20.14 as=1.5972 ps=10.01 w=9.68 l=0.2
X15 VDD1.t0 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5972 pd=10.01 as=3.7752 ps=20.14 w=9.68 l=0.2
R0 VN.n2 VN.t4 1363.99
R1 VN.n0 VN.t5 1363.99
R2 VN.n6 VN.t1 1363.99
R3 VN.n4 VN.t3 1363.99
R4 VN.n1 VN.t0 1323.09
R5 VN.n5 VN.t2 1323.09
R6 VN.n7 VN.n4 161.489
R7 VN.n3 VN.n0 161.489
R8 VN.n3 VN.n2 161.3
R9 VN.n7 VN.n6 161.3
R10 VN VN.n7 37.9304
R11 VN.n1 VN.n0 36.5157
R12 VN.n2 VN.n1 36.5157
R13 VN.n6 VN.n5 36.5157
R14 VN.n5 VN.n4 36.5157
R15 VN VN.n3 0.0516364
R16 VDD2.n1 VDD2.t5 66.6962
R17 VDD2.n2 VDD2.t0 66.409
R18 VDD2.n1 VDD2.n0 64.4223
R19 VDD2 VDD2.n3 64.4195
R20 VDD2.n2 VDD2.n1 33.545
R21 VDD2.n3 VDD2.t1 2.04595
R22 VDD2.n3 VDD2.t4 2.04595
R23 VDD2.n0 VDD2.t2 2.04595
R24 VDD2.n0 VDD2.t3 2.04595
R25 VDD2 VDD2.n2 0.401362
R26 VTAIL.n7 VTAIL.t5 49.7302
R27 VTAIL.n11 VTAIL.t4 49.7301
R28 VTAIL.n2 VTAIL.t10 49.7301
R29 VTAIL.n10 VTAIL.t2 49.7301
R30 VTAIL.n9 VTAIL.n8 47.6848
R31 VTAIL.n6 VTAIL.n5 47.6848
R32 VTAIL.n1 VTAIL.n0 47.6846
R33 VTAIL.n4 VTAIL.n3 47.6846
R34 VTAIL.n6 VTAIL.n4 21.6255
R35 VTAIL.n11 VTAIL.n10 21.1686
R36 VTAIL.n0 VTAIL.t3 2.04595
R37 VTAIL.n0 VTAIL.t8 2.04595
R38 VTAIL.n3 VTAIL.t1 2.04595
R39 VTAIL.n3 VTAIL.t9 2.04595
R40 VTAIL.n8 VTAIL.t0 2.04595
R41 VTAIL.n8 VTAIL.t11 2.04595
R42 VTAIL.n5 VTAIL.t7 2.04595
R43 VTAIL.n5 VTAIL.t6 2.04595
R44 VTAIL.n9 VTAIL.n7 0.698776
R45 VTAIL.n2 VTAIL.n1 0.698776
R46 VTAIL.n7 VTAIL.n6 0.457397
R47 VTAIL.n10 VTAIL.n9 0.457397
R48 VTAIL.n4 VTAIL.n2 0.457397
R49 VTAIL VTAIL.n11 0.284983
R50 VTAIL VTAIL.n1 0.172914
R51 B.n75 B.t10 1402.79
R52 B.n72 B.t17 1402.79
R53 B.n282 B.t6 1402.79
R54 B.n276 B.t14 1402.79
R55 B.n521 B.n520 585
R56 B.n522 B.n521 585
R57 B.n230 B.n71 585
R58 B.n229 B.n228 585
R59 B.n227 B.n226 585
R60 B.n225 B.n224 585
R61 B.n223 B.n222 585
R62 B.n221 B.n220 585
R63 B.n219 B.n218 585
R64 B.n217 B.n216 585
R65 B.n215 B.n214 585
R66 B.n213 B.n212 585
R67 B.n211 B.n210 585
R68 B.n209 B.n208 585
R69 B.n207 B.n206 585
R70 B.n205 B.n204 585
R71 B.n203 B.n202 585
R72 B.n201 B.n200 585
R73 B.n199 B.n198 585
R74 B.n197 B.n196 585
R75 B.n195 B.n194 585
R76 B.n193 B.n192 585
R77 B.n191 B.n190 585
R78 B.n189 B.n188 585
R79 B.n187 B.n186 585
R80 B.n185 B.n184 585
R81 B.n183 B.n182 585
R82 B.n181 B.n180 585
R83 B.n179 B.n178 585
R84 B.n177 B.n176 585
R85 B.n175 B.n174 585
R86 B.n173 B.n172 585
R87 B.n171 B.n170 585
R88 B.n169 B.n168 585
R89 B.n167 B.n166 585
R90 B.n165 B.n164 585
R91 B.n163 B.n162 585
R92 B.n161 B.n160 585
R93 B.n159 B.n158 585
R94 B.n157 B.n156 585
R95 B.n155 B.n154 585
R96 B.n153 B.n152 585
R97 B.n151 B.n150 585
R98 B.n149 B.n148 585
R99 B.n147 B.n146 585
R100 B.n144 B.n143 585
R101 B.n142 B.n141 585
R102 B.n140 B.n139 585
R103 B.n138 B.n137 585
R104 B.n136 B.n135 585
R105 B.n134 B.n133 585
R106 B.n132 B.n131 585
R107 B.n130 B.n129 585
R108 B.n128 B.n127 585
R109 B.n126 B.n125 585
R110 B.n124 B.n123 585
R111 B.n122 B.n121 585
R112 B.n120 B.n119 585
R113 B.n118 B.n117 585
R114 B.n116 B.n115 585
R115 B.n114 B.n113 585
R116 B.n112 B.n111 585
R117 B.n110 B.n109 585
R118 B.n108 B.n107 585
R119 B.n106 B.n105 585
R120 B.n104 B.n103 585
R121 B.n102 B.n101 585
R122 B.n100 B.n99 585
R123 B.n98 B.n97 585
R124 B.n96 B.n95 585
R125 B.n94 B.n93 585
R126 B.n92 B.n91 585
R127 B.n90 B.n89 585
R128 B.n88 B.n87 585
R129 B.n86 B.n85 585
R130 B.n84 B.n83 585
R131 B.n82 B.n81 585
R132 B.n80 B.n79 585
R133 B.n78 B.n77 585
R134 B.n30 B.n29 585
R135 B.n519 B.n31 585
R136 B.n523 B.n31 585
R137 B.n518 B.n517 585
R138 B.n517 B.n27 585
R139 B.n516 B.n26 585
R140 B.n529 B.n26 585
R141 B.n515 B.n25 585
R142 B.n530 B.n25 585
R143 B.n514 B.n24 585
R144 B.n531 B.n24 585
R145 B.n513 B.n512 585
R146 B.n512 B.n20 585
R147 B.n511 B.n19 585
R148 B.n537 B.n19 585
R149 B.n510 B.n18 585
R150 B.n538 B.n18 585
R151 B.n509 B.n17 585
R152 B.n539 B.n17 585
R153 B.n508 B.n507 585
R154 B.n507 B.t2 585
R155 B.n506 B.n12 585
R156 B.n545 B.n12 585
R157 B.n505 B.n11 585
R158 B.n546 B.n11 585
R159 B.n504 B.n10 585
R160 B.n547 B.n10 585
R161 B.n503 B.n7 585
R162 B.n550 B.n7 585
R163 B.n502 B.n6 585
R164 B.n551 B.n6 585
R165 B.n501 B.n5 585
R166 B.n552 B.n5 585
R167 B.n500 B.n499 585
R168 B.n499 B.n4 585
R169 B.n498 B.n231 585
R170 B.n498 B.n497 585
R171 B.n488 B.n232 585
R172 B.n233 B.n232 585
R173 B.n490 B.n489 585
R174 B.n491 B.n490 585
R175 B.n487 B.n237 585
R176 B.n237 B.t1 585
R177 B.n486 B.n485 585
R178 B.n485 B.n484 585
R179 B.n239 B.n238 585
R180 B.n240 B.n239 585
R181 B.n477 B.n476 585
R182 B.n478 B.n477 585
R183 B.n475 B.n245 585
R184 B.n245 B.n244 585
R185 B.n474 B.n473 585
R186 B.n473 B.n472 585
R187 B.n247 B.n246 585
R188 B.n248 B.n247 585
R189 B.n465 B.n464 585
R190 B.n466 B.n465 585
R191 B.n463 B.n253 585
R192 B.n253 B.n252 585
R193 B.n462 B.n461 585
R194 B.n461 B.n460 585
R195 B.n457 B.n257 585
R196 B.n456 B.n455 585
R197 B.n453 B.n258 585
R198 B.n453 B.n256 585
R199 B.n452 B.n451 585
R200 B.n450 B.n449 585
R201 B.n448 B.n260 585
R202 B.n446 B.n445 585
R203 B.n444 B.n261 585
R204 B.n443 B.n442 585
R205 B.n440 B.n262 585
R206 B.n438 B.n437 585
R207 B.n436 B.n263 585
R208 B.n435 B.n434 585
R209 B.n432 B.n264 585
R210 B.n430 B.n429 585
R211 B.n428 B.n265 585
R212 B.n427 B.n426 585
R213 B.n424 B.n266 585
R214 B.n422 B.n421 585
R215 B.n420 B.n267 585
R216 B.n419 B.n418 585
R217 B.n416 B.n268 585
R218 B.n414 B.n413 585
R219 B.n412 B.n269 585
R220 B.n411 B.n410 585
R221 B.n408 B.n270 585
R222 B.n406 B.n405 585
R223 B.n404 B.n271 585
R224 B.n403 B.n402 585
R225 B.n400 B.n272 585
R226 B.n398 B.n397 585
R227 B.n396 B.n273 585
R228 B.n395 B.n394 585
R229 B.n392 B.n274 585
R230 B.n390 B.n389 585
R231 B.n387 B.n275 585
R232 B.n386 B.n385 585
R233 B.n383 B.n278 585
R234 B.n381 B.n380 585
R235 B.n379 B.n279 585
R236 B.n378 B.n377 585
R237 B.n375 B.n280 585
R238 B.n373 B.n372 585
R239 B.n371 B.n281 585
R240 B.n369 B.n368 585
R241 B.n366 B.n284 585
R242 B.n364 B.n363 585
R243 B.n362 B.n285 585
R244 B.n361 B.n360 585
R245 B.n358 B.n286 585
R246 B.n356 B.n355 585
R247 B.n354 B.n287 585
R248 B.n353 B.n352 585
R249 B.n350 B.n288 585
R250 B.n348 B.n347 585
R251 B.n346 B.n289 585
R252 B.n345 B.n344 585
R253 B.n342 B.n290 585
R254 B.n340 B.n339 585
R255 B.n338 B.n291 585
R256 B.n337 B.n336 585
R257 B.n334 B.n292 585
R258 B.n332 B.n331 585
R259 B.n330 B.n293 585
R260 B.n329 B.n328 585
R261 B.n326 B.n294 585
R262 B.n324 B.n323 585
R263 B.n322 B.n295 585
R264 B.n321 B.n320 585
R265 B.n318 B.n296 585
R266 B.n316 B.n315 585
R267 B.n314 B.n297 585
R268 B.n313 B.n312 585
R269 B.n310 B.n298 585
R270 B.n308 B.n307 585
R271 B.n306 B.n299 585
R272 B.n305 B.n304 585
R273 B.n302 B.n300 585
R274 B.n255 B.n254 585
R275 B.n459 B.n458 585
R276 B.n460 B.n459 585
R277 B.n251 B.n250 585
R278 B.n252 B.n251 585
R279 B.n468 B.n467 585
R280 B.n467 B.n466 585
R281 B.n469 B.n249 585
R282 B.n249 B.n248 585
R283 B.n471 B.n470 585
R284 B.n472 B.n471 585
R285 B.n243 B.n242 585
R286 B.n244 B.n243 585
R287 B.n480 B.n479 585
R288 B.n479 B.n478 585
R289 B.n481 B.n241 585
R290 B.n241 B.n240 585
R291 B.n483 B.n482 585
R292 B.n484 B.n483 585
R293 B.n236 B.n235 585
R294 B.t1 B.n236 585
R295 B.n493 B.n492 585
R296 B.n492 B.n491 585
R297 B.n494 B.n234 585
R298 B.n234 B.n233 585
R299 B.n496 B.n495 585
R300 B.n497 B.n496 585
R301 B.n3 B.n0 585
R302 B.n4 B.n3 585
R303 B.n549 B.n1 585
R304 B.n550 B.n549 585
R305 B.n548 B.n9 585
R306 B.n548 B.n547 585
R307 B.n14 B.n8 585
R308 B.n546 B.n8 585
R309 B.n544 B.n543 585
R310 B.n545 B.n544 585
R311 B.n542 B.n13 585
R312 B.n13 B.t2 585
R313 B.n541 B.n540 585
R314 B.n540 B.n539 585
R315 B.n16 B.n15 585
R316 B.n538 B.n16 585
R317 B.n536 B.n535 585
R318 B.n537 B.n536 585
R319 B.n534 B.n21 585
R320 B.n21 B.n20 585
R321 B.n533 B.n532 585
R322 B.n532 B.n531 585
R323 B.n23 B.n22 585
R324 B.n530 B.n23 585
R325 B.n528 B.n527 585
R326 B.n529 B.n528 585
R327 B.n526 B.n28 585
R328 B.n28 B.n27 585
R329 B.n525 B.n524 585
R330 B.n524 B.n523 585
R331 B.n553 B.n552 585
R332 B.n551 B.n2 585
R333 B.n524 B.n30 487.695
R334 B.n521 B.n31 487.695
R335 B.n461 B.n255 487.695
R336 B.n459 B.n257 487.695
R337 B.n522 B.n70 256.663
R338 B.n522 B.n69 256.663
R339 B.n522 B.n68 256.663
R340 B.n522 B.n67 256.663
R341 B.n522 B.n66 256.663
R342 B.n522 B.n65 256.663
R343 B.n522 B.n64 256.663
R344 B.n522 B.n63 256.663
R345 B.n522 B.n62 256.663
R346 B.n522 B.n61 256.663
R347 B.n522 B.n60 256.663
R348 B.n522 B.n59 256.663
R349 B.n522 B.n58 256.663
R350 B.n522 B.n57 256.663
R351 B.n522 B.n56 256.663
R352 B.n522 B.n55 256.663
R353 B.n522 B.n54 256.663
R354 B.n522 B.n53 256.663
R355 B.n522 B.n52 256.663
R356 B.n522 B.n51 256.663
R357 B.n522 B.n50 256.663
R358 B.n522 B.n49 256.663
R359 B.n522 B.n48 256.663
R360 B.n522 B.n47 256.663
R361 B.n522 B.n46 256.663
R362 B.n522 B.n45 256.663
R363 B.n522 B.n44 256.663
R364 B.n522 B.n43 256.663
R365 B.n522 B.n42 256.663
R366 B.n522 B.n41 256.663
R367 B.n522 B.n40 256.663
R368 B.n522 B.n39 256.663
R369 B.n522 B.n38 256.663
R370 B.n522 B.n37 256.663
R371 B.n522 B.n36 256.663
R372 B.n522 B.n35 256.663
R373 B.n522 B.n34 256.663
R374 B.n522 B.n33 256.663
R375 B.n522 B.n32 256.663
R376 B.n454 B.n256 256.663
R377 B.n259 B.n256 256.663
R378 B.n447 B.n256 256.663
R379 B.n441 B.n256 256.663
R380 B.n439 B.n256 256.663
R381 B.n433 B.n256 256.663
R382 B.n431 B.n256 256.663
R383 B.n425 B.n256 256.663
R384 B.n423 B.n256 256.663
R385 B.n417 B.n256 256.663
R386 B.n415 B.n256 256.663
R387 B.n409 B.n256 256.663
R388 B.n407 B.n256 256.663
R389 B.n401 B.n256 256.663
R390 B.n399 B.n256 256.663
R391 B.n393 B.n256 256.663
R392 B.n391 B.n256 256.663
R393 B.n384 B.n256 256.663
R394 B.n382 B.n256 256.663
R395 B.n376 B.n256 256.663
R396 B.n374 B.n256 256.663
R397 B.n367 B.n256 256.663
R398 B.n365 B.n256 256.663
R399 B.n359 B.n256 256.663
R400 B.n357 B.n256 256.663
R401 B.n351 B.n256 256.663
R402 B.n349 B.n256 256.663
R403 B.n343 B.n256 256.663
R404 B.n341 B.n256 256.663
R405 B.n335 B.n256 256.663
R406 B.n333 B.n256 256.663
R407 B.n327 B.n256 256.663
R408 B.n325 B.n256 256.663
R409 B.n319 B.n256 256.663
R410 B.n317 B.n256 256.663
R411 B.n311 B.n256 256.663
R412 B.n309 B.n256 256.663
R413 B.n303 B.n256 256.663
R414 B.n301 B.n256 256.663
R415 B.n555 B.n554 256.663
R416 B.n79 B.n78 163.367
R417 B.n83 B.n82 163.367
R418 B.n87 B.n86 163.367
R419 B.n91 B.n90 163.367
R420 B.n95 B.n94 163.367
R421 B.n99 B.n98 163.367
R422 B.n103 B.n102 163.367
R423 B.n107 B.n106 163.367
R424 B.n111 B.n110 163.367
R425 B.n115 B.n114 163.367
R426 B.n119 B.n118 163.367
R427 B.n123 B.n122 163.367
R428 B.n127 B.n126 163.367
R429 B.n131 B.n130 163.367
R430 B.n135 B.n134 163.367
R431 B.n139 B.n138 163.367
R432 B.n143 B.n142 163.367
R433 B.n148 B.n147 163.367
R434 B.n152 B.n151 163.367
R435 B.n156 B.n155 163.367
R436 B.n160 B.n159 163.367
R437 B.n164 B.n163 163.367
R438 B.n168 B.n167 163.367
R439 B.n172 B.n171 163.367
R440 B.n176 B.n175 163.367
R441 B.n180 B.n179 163.367
R442 B.n184 B.n183 163.367
R443 B.n188 B.n187 163.367
R444 B.n192 B.n191 163.367
R445 B.n196 B.n195 163.367
R446 B.n200 B.n199 163.367
R447 B.n204 B.n203 163.367
R448 B.n208 B.n207 163.367
R449 B.n212 B.n211 163.367
R450 B.n216 B.n215 163.367
R451 B.n220 B.n219 163.367
R452 B.n224 B.n223 163.367
R453 B.n228 B.n227 163.367
R454 B.n521 B.n71 163.367
R455 B.n461 B.n253 163.367
R456 B.n465 B.n253 163.367
R457 B.n465 B.n247 163.367
R458 B.n473 B.n247 163.367
R459 B.n473 B.n245 163.367
R460 B.n477 B.n245 163.367
R461 B.n477 B.n239 163.367
R462 B.n485 B.n239 163.367
R463 B.n485 B.n237 163.367
R464 B.n490 B.n237 163.367
R465 B.n490 B.n232 163.367
R466 B.n498 B.n232 163.367
R467 B.n499 B.n498 163.367
R468 B.n499 B.n5 163.367
R469 B.n6 B.n5 163.367
R470 B.n7 B.n6 163.367
R471 B.n10 B.n7 163.367
R472 B.n11 B.n10 163.367
R473 B.n12 B.n11 163.367
R474 B.n507 B.n12 163.367
R475 B.n507 B.n17 163.367
R476 B.n18 B.n17 163.367
R477 B.n19 B.n18 163.367
R478 B.n512 B.n19 163.367
R479 B.n512 B.n24 163.367
R480 B.n25 B.n24 163.367
R481 B.n26 B.n25 163.367
R482 B.n517 B.n26 163.367
R483 B.n517 B.n31 163.367
R484 B.n455 B.n453 163.367
R485 B.n453 B.n452 163.367
R486 B.n449 B.n448 163.367
R487 B.n446 B.n261 163.367
R488 B.n442 B.n440 163.367
R489 B.n438 B.n263 163.367
R490 B.n434 B.n432 163.367
R491 B.n430 B.n265 163.367
R492 B.n426 B.n424 163.367
R493 B.n422 B.n267 163.367
R494 B.n418 B.n416 163.367
R495 B.n414 B.n269 163.367
R496 B.n410 B.n408 163.367
R497 B.n406 B.n271 163.367
R498 B.n402 B.n400 163.367
R499 B.n398 B.n273 163.367
R500 B.n394 B.n392 163.367
R501 B.n390 B.n275 163.367
R502 B.n385 B.n383 163.367
R503 B.n381 B.n279 163.367
R504 B.n377 B.n375 163.367
R505 B.n373 B.n281 163.367
R506 B.n368 B.n366 163.367
R507 B.n364 B.n285 163.367
R508 B.n360 B.n358 163.367
R509 B.n356 B.n287 163.367
R510 B.n352 B.n350 163.367
R511 B.n348 B.n289 163.367
R512 B.n344 B.n342 163.367
R513 B.n340 B.n291 163.367
R514 B.n336 B.n334 163.367
R515 B.n332 B.n293 163.367
R516 B.n328 B.n326 163.367
R517 B.n324 B.n295 163.367
R518 B.n320 B.n318 163.367
R519 B.n316 B.n297 163.367
R520 B.n312 B.n310 163.367
R521 B.n308 B.n299 163.367
R522 B.n304 B.n302 163.367
R523 B.n459 B.n251 163.367
R524 B.n467 B.n251 163.367
R525 B.n467 B.n249 163.367
R526 B.n471 B.n249 163.367
R527 B.n471 B.n243 163.367
R528 B.n479 B.n243 163.367
R529 B.n479 B.n241 163.367
R530 B.n483 B.n241 163.367
R531 B.n483 B.n236 163.367
R532 B.n492 B.n236 163.367
R533 B.n492 B.n234 163.367
R534 B.n496 B.n234 163.367
R535 B.n496 B.n3 163.367
R536 B.n553 B.n3 163.367
R537 B.n549 B.n2 163.367
R538 B.n549 B.n548 163.367
R539 B.n548 B.n8 163.367
R540 B.n544 B.n8 163.367
R541 B.n544 B.n13 163.367
R542 B.n540 B.n13 163.367
R543 B.n540 B.n16 163.367
R544 B.n536 B.n16 163.367
R545 B.n536 B.n21 163.367
R546 B.n532 B.n21 163.367
R547 B.n532 B.n23 163.367
R548 B.n528 B.n23 163.367
R549 B.n528 B.n28 163.367
R550 B.n524 B.n28 163.367
R551 B.n460 B.n256 83.1165
R552 B.n523 B.n522 83.1165
R553 B.n72 B.t18 81.5637
R554 B.n282 B.t9 81.5637
R555 B.n75 B.t12 81.552
R556 B.n276 B.t16 81.552
R557 B.n32 B.n30 71.676
R558 B.n79 B.n33 71.676
R559 B.n83 B.n34 71.676
R560 B.n87 B.n35 71.676
R561 B.n91 B.n36 71.676
R562 B.n95 B.n37 71.676
R563 B.n99 B.n38 71.676
R564 B.n103 B.n39 71.676
R565 B.n107 B.n40 71.676
R566 B.n111 B.n41 71.676
R567 B.n115 B.n42 71.676
R568 B.n119 B.n43 71.676
R569 B.n123 B.n44 71.676
R570 B.n127 B.n45 71.676
R571 B.n131 B.n46 71.676
R572 B.n135 B.n47 71.676
R573 B.n139 B.n48 71.676
R574 B.n143 B.n49 71.676
R575 B.n148 B.n50 71.676
R576 B.n152 B.n51 71.676
R577 B.n156 B.n52 71.676
R578 B.n160 B.n53 71.676
R579 B.n164 B.n54 71.676
R580 B.n168 B.n55 71.676
R581 B.n172 B.n56 71.676
R582 B.n176 B.n57 71.676
R583 B.n180 B.n58 71.676
R584 B.n184 B.n59 71.676
R585 B.n188 B.n60 71.676
R586 B.n192 B.n61 71.676
R587 B.n196 B.n62 71.676
R588 B.n200 B.n63 71.676
R589 B.n204 B.n64 71.676
R590 B.n208 B.n65 71.676
R591 B.n212 B.n66 71.676
R592 B.n216 B.n67 71.676
R593 B.n220 B.n68 71.676
R594 B.n224 B.n69 71.676
R595 B.n228 B.n70 71.676
R596 B.n71 B.n70 71.676
R597 B.n227 B.n69 71.676
R598 B.n223 B.n68 71.676
R599 B.n219 B.n67 71.676
R600 B.n215 B.n66 71.676
R601 B.n211 B.n65 71.676
R602 B.n207 B.n64 71.676
R603 B.n203 B.n63 71.676
R604 B.n199 B.n62 71.676
R605 B.n195 B.n61 71.676
R606 B.n191 B.n60 71.676
R607 B.n187 B.n59 71.676
R608 B.n183 B.n58 71.676
R609 B.n179 B.n57 71.676
R610 B.n175 B.n56 71.676
R611 B.n171 B.n55 71.676
R612 B.n167 B.n54 71.676
R613 B.n163 B.n53 71.676
R614 B.n159 B.n52 71.676
R615 B.n155 B.n51 71.676
R616 B.n151 B.n50 71.676
R617 B.n147 B.n49 71.676
R618 B.n142 B.n48 71.676
R619 B.n138 B.n47 71.676
R620 B.n134 B.n46 71.676
R621 B.n130 B.n45 71.676
R622 B.n126 B.n44 71.676
R623 B.n122 B.n43 71.676
R624 B.n118 B.n42 71.676
R625 B.n114 B.n41 71.676
R626 B.n110 B.n40 71.676
R627 B.n106 B.n39 71.676
R628 B.n102 B.n38 71.676
R629 B.n98 B.n37 71.676
R630 B.n94 B.n36 71.676
R631 B.n90 B.n35 71.676
R632 B.n86 B.n34 71.676
R633 B.n82 B.n33 71.676
R634 B.n78 B.n32 71.676
R635 B.n454 B.n257 71.676
R636 B.n452 B.n259 71.676
R637 B.n448 B.n447 71.676
R638 B.n441 B.n261 71.676
R639 B.n440 B.n439 71.676
R640 B.n433 B.n263 71.676
R641 B.n432 B.n431 71.676
R642 B.n425 B.n265 71.676
R643 B.n424 B.n423 71.676
R644 B.n417 B.n267 71.676
R645 B.n416 B.n415 71.676
R646 B.n409 B.n269 71.676
R647 B.n408 B.n407 71.676
R648 B.n401 B.n271 71.676
R649 B.n400 B.n399 71.676
R650 B.n393 B.n273 71.676
R651 B.n392 B.n391 71.676
R652 B.n384 B.n275 71.676
R653 B.n383 B.n382 71.676
R654 B.n376 B.n279 71.676
R655 B.n375 B.n374 71.676
R656 B.n367 B.n281 71.676
R657 B.n366 B.n365 71.676
R658 B.n359 B.n285 71.676
R659 B.n358 B.n357 71.676
R660 B.n351 B.n287 71.676
R661 B.n350 B.n349 71.676
R662 B.n343 B.n289 71.676
R663 B.n342 B.n341 71.676
R664 B.n335 B.n291 71.676
R665 B.n334 B.n333 71.676
R666 B.n327 B.n293 71.676
R667 B.n326 B.n325 71.676
R668 B.n319 B.n295 71.676
R669 B.n318 B.n317 71.676
R670 B.n311 B.n297 71.676
R671 B.n310 B.n309 71.676
R672 B.n303 B.n299 71.676
R673 B.n302 B.n301 71.676
R674 B.n455 B.n454 71.676
R675 B.n449 B.n259 71.676
R676 B.n447 B.n446 71.676
R677 B.n442 B.n441 71.676
R678 B.n439 B.n438 71.676
R679 B.n434 B.n433 71.676
R680 B.n431 B.n430 71.676
R681 B.n426 B.n425 71.676
R682 B.n423 B.n422 71.676
R683 B.n418 B.n417 71.676
R684 B.n415 B.n414 71.676
R685 B.n410 B.n409 71.676
R686 B.n407 B.n406 71.676
R687 B.n402 B.n401 71.676
R688 B.n399 B.n398 71.676
R689 B.n394 B.n393 71.676
R690 B.n391 B.n390 71.676
R691 B.n385 B.n384 71.676
R692 B.n382 B.n381 71.676
R693 B.n377 B.n376 71.676
R694 B.n374 B.n373 71.676
R695 B.n368 B.n367 71.676
R696 B.n365 B.n364 71.676
R697 B.n360 B.n359 71.676
R698 B.n357 B.n356 71.676
R699 B.n352 B.n351 71.676
R700 B.n349 B.n348 71.676
R701 B.n344 B.n343 71.676
R702 B.n341 B.n340 71.676
R703 B.n336 B.n335 71.676
R704 B.n333 B.n332 71.676
R705 B.n328 B.n327 71.676
R706 B.n325 B.n324 71.676
R707 B.n320 B.n319 71.676
R708 B.n317 B.n316 71.676
R709 B.n312 B.n311 71.676
R710 B.n309 B.n308 71.676
R711 B.n304 B.n303 71.676
R712 B.n301 B.n255 71.676
R713 B.n554 B.n553 71.676
R714 B.n554 B.n2 71.676
R715 B.n73 B.t19 71.2849
R716 B.n283 B.t8 71.2849
R717 B.n76 B.t13 71.2732
R718 B.n277 B.t15 71.2732
R719 B.n145 B.n76 59.5399
R720 B.n74 B.n73 59.5399
R721 B.n370 B.n283 59.5399
R722 B.n388 B.n277 59.5399
R723 B.n460 B.n252 50.0172
R724 B.n466 B.n252 50.0172
R725 B.n466 B.n248 50.0172
R726 B.n472 B.n248 50.0172
R727 B.n478 B.n244 50.0172
R728 B.n478 B.n240 50.0172
R729 B.n484 B.n240 50.0172
R730 B.n484 B.t1 50.0172
R731 B.n491 B.t1 50.0172
R732 B.n497 B.n233 50.0172
R733 B.n552 B.n4 50.0172
R734 B.n552 B.n551 50.0172
R735 B.n551 B.n550 50.0172
R736 B.n547 B.n546 50.0172
R737 B.n545 B.t2 50.0172
R738 B.n539 B.t2 50.0172
R739 B.n539 B.n538 50.0172
R740 B.n538 B.n537 50.0172
R741 B.n537 B.n20 50.0172
R742 B.n531 B.n530 50.0172
R743 B.n530 B.n529 50.0172
R744 B.n529 B.n27 50.0172
R745 B.n523 B.n27 50.0172
R746 B.t3 B.n4 44.1329
R747 B.n550 B.t0 44.1329
R748 B.t7 B.n244 38.2486
R749 B.t11 B.n20 38.2486
R750 B.n458 B.n457 31.6883
R751 B.n462 B.n254 31.6883
R752 B.n520 B.n519 31.6883
R753 B.n525 B.n29 31.6883
R754 B.n491 B.t4 27.951
R755 B.t5 B.n545 27.951
R756 B.t4 B.n233 22.0667
R757 B.n546 B.t5 22.0667
R758 B B.n555 18.0485
R759 B.n472 B.t7 11.7691
R760 B.n531 B.t11 11.7691
R761 B.n458 B.n250 10.6151
R762 B.n468 B.n250 10.6151
R763 B.n469 B.n468 10.6151
R764 B.n470 B.n469 10.6151
R765 B.n470 B.n242 10.6151
R766 B.n480 B.n242 10.6151
R767 B.n481 B.n480 10.6151
R768 B.n482 B.n481 10.6151
R769 B.n482 B.n235 10.6151
R770 B.n493 B.n235 10.6151
R771 B.n494 B.n493 10.6151
R772 B.n495 B.n494 10.6151
R773 B.n495 B.n0 10.6151
R774 B.n457 B.n456 10.6151
R775 B.n456 B.n258 10.6151
R776 B.n451 B.n258 10.6151
R777 B.n451 B.n450 10.6151
R778 B.n450 B.n260 10.6151
R779 B.n445 B.n260 10.6151
R780 B.n445 B.n444 10.6151
R781 B.n444 B.n443 10.6151
R782 B.n443 B.n262 10.6151
R783 B.n437 B.n262 10.6151
R784 B.n437 B.n436 10.6151
R785 B.n436 B.n435 10.6151
R786 B.n435 B.n264 10.6151
R787 B.n429 B.n264 10.6151
R788 B.n429 B.n428 10.6151
R789 B.n428 B.n427 10.6151
R790 B.n427 B.n266 10.6151
R791 B.n421 B.n266 10.6151
R792 B.n421 B.n420 10.6151
R793 B.n420 B.n419 10.6151
R794 B.n419 B.n268 10.6151
R795 B.n413 B.n268 10.6151
R796 B.n413 B.n412 10.6151
R797 B.n412 B.n411 10.6151
R798 B.n411 B.n270 10.6151
R799 B.n405 B.n270 10.6151
R800 B.n405 B.n404 10.6151
R801 B.n404 B.n403 10.6151
R802 B.n403 B.n272 10.6151
R803 B.n397 B.n272 10.6151
R804 B.n397 B.n396 10.6151
R805 B.n396 B.n395 10.6151
R806 B.n395 B.n274 10.6151
R807 B.n389 B.n274 10.6151
R808 B.n387 B.n386 10.6151
R809 B.n386 B.n278 10.6151
R810 B.n380 B.n278 10.6151
R811 B.n380 B.n379 10.6151
R812 B.n379 B.n378 10.6151
R813 B.n378 B.n280 10.6151
R814 B.n372 B.n280 10.6151
R815 B.n372 B.n371 10.6151
R816 B.n369 B.n284 10.6151
R817 B.n363 B.n284 10.6151
R818 B.n363 B.n362 10.6151
R819 B.n362 B.n361 10.6151
R820 B.n361 B.n286 10.6151
R821 B.n355 B.n286 10.6151
R822 B.n355 B.n354 10.6151
R823 B.n354 B.n353 10.6151
R824 B.n353 B.n288 10.6151
R825 B.n347 B.n288 10.6151
R826 B.n347 B.n346 10.6151
R827 B.n346 B.n345 10.6151
R828 B.n345 B.n290 10.6151
R829 B.n339 B.n290 10.6151
R830 B.n339 B.n338 10.6151
R831 B.n338 B.n337 10.6151
R832 B.n337 B.n292 10.6151
R833 B.n331 B.n292 10.6151
R834 B.n331 B.n330 10.6151
R835 B.n330 B.n329 10.6151
R836 B.n329 B.n294 10.6151
R837 B.n323 B.n294 10.6151
R838 B.n323 B.n322 10.6151
R839 B.n322 B.n321 10.6151
R840 B.n321 B.n296 10.6151
R841 B.n315 B.n296 10.6151
R842 B.n315 B.n314 10.6151
R843 B.n314 B.n313 10.6151
R844 B.n313 B.n298 10.6151
R845 B.n307 B.n298 10.6151
R846 B.n307 B.n306 10.6151
R847 B.n306 B.n305 10.6151
R848 B.n305 B.n300 10.6151
R849 B.n300 B.n254 10.6151
R850 B.n463 B.n462 10.6151
R851 B.n464 B.n463 10.6151
R852 B.n464 B.n246 10.6151
R853 B.n474 B.n246 10.6151
R854 B.n475 B.n474 10.6151
R855 B.n476 B.n475 10.6151
R856 B.n476 B.n238 10.6151
R857 B.n486 B.n238 10.6151
R858 B.n487 B.n486 10.6151
R859 B.n489 B.n487 10.6151
R860 B.n489 B.n488 10.6151
R861 B.n488 B.n231 10.6151
R862 B.n500 B.n231 10.6151
R863 B.n501 B.n500 10.6151
R864 B.n502 B.n501 10.6151
R865 B.n503 B.n502 10.6151
R866 B.n504 B.n503 10.6151
R867 B.n505 B.n504 10.6151
R868 B.n506 B.n505 10.6151
R869 B.n508 B.n506 10.6151
R870 B.n509 B.n508 10.6151
R871 B.n510 B.n509 10.6151
R872 B.n511 B.n510 10.6151
R873 B.n513 B.n511 10.6151
R874 B.n514 B.n513 10.6151
R875 B.n515 B.n514 10.6151
R876 B.n516 B.n515 10.6151
R877 B.n518 B.n516 10.6151
R878 B.n519 B.n518 10.6151
R879 B.n9 B.n1 10.6151
R880 B.n14 B.n9 10.6151
R881 B.n543 B.n14 10.6151
R882 B.n543 B.n542 10.6151
R883 B.n542 B.n541 10.6151
R884 B.n541 B.n15 10.6151
R885 B.n535 B.n15 10.6151
R886 B.n535 B.n534 10.6151
R887 B.n534 B.n533 10.6151
R888 B.n533 B.n22 10.6151
R889 B.n527 B.n22 10.6151
R890 B.n527 B.n526 10.6151
R891 B.n526 B.n525 10.6151
R892 B.n77 B.n29 10.6151
R893 B.n80 B.n77 10.6151
R894 B.n81 B.n80 10.6151
R895 B.n84 B.n81 10.6151
R896 B.n85 B.n84 10.6151
R897 B.n88 B.n85 10.6151
R898 B.n89 B.n88 10.6151
R899 B.n92 B.n89 10.6151
R900 B.n93 B.n92 10.6151
R901 B.n96 B.n93 10.6151
R902 B.n97 B.n96 10.6151
R903 B.n100 B.n97 10.6151
R904 B.n101 B.n100 10.6151
R905 B.n104 B.n101 10.6151
R906 B.n105 B.n104 10.6151
R907 B.n108 B.n105 10.6151
R908 B.n109 B.n108 10.6151
R909 B.n112 B.n109 10.6151
R910 B.n113 B.n112 10.6151
R911 B.n116 B.n113 10.6151
R912 B.n117 B.n116 10.6151
R913 B.n120 B.n117 10.6151
R914 B.n121 B.n120 10.6151
R915 B.n124 B.n121 10.6151
R916 B.n125 B.n124 10.6151
R917 B.n128 B.n125 10.6151
R918 B.n129 B.n128 10.6151
R919 B.n132 B.n129 10.6151
R920 B.n133 B.n132 10.6151
R921 B.n136 B.n133 10.6151
R922 B.n137 B.n136 10.6151
R923 B.n140 B.n137 10.6151
R924 B.n141 B.n140 10.6151
R925 B.n144 B.n141 10.6151
R926 B.n149 B.n146 10.6151
R927 B.n150 B.n149 10.6151
R928 B.n153 B.n150 10.6151
R929 B.n154 B.n153 10.6151
R930 B.n157 B.n154 10.6151
R931 B.n158 B.n157 10.6151
R932 B.n161 B.n158 10.6151
R933 B.n162 B.n161 10.6151
R934 B.n166 B.n165 10.6151
R935 B.n169 B.n166 10.6151
R936 B.n170 B.n169 10.6151
R937 B.n173 B.n170 10.6151
R938 B.n174 B.n173 10.6151
R939 B.n177 B.n174 10.6151
R940 B.n178 B.n177 10.6151
R941 B.n181 B.n178 10.6151
R942 B.n182 B.n181 10.6151
R943 B.n185 B.n182 10.6151
R944 B.n186 B.n185 10.6151
R945 B.n189 B.n186 10.6151
R946 B.n190 B.n189 10.6151
R947 B.n193 B.n190 10.6151
R948 B.n194 B.n193 10.6151
R949 B.n197 B.n194 10.6151
R950 B.n198 B.n197 10.6151
R951 B.n201 B.n198 10.6151
R952 B.n202 B.n201 10.6151
R953 B.n205 B.n202 10.6151
R954 B.n206 B.n205 10.6151
R955 B.n209 B.n206 10.6151
R956 B.n210 B.n209 10.6151
R957 B.n213 B.n210 10.6151
R958 B.n214 B.n213 10.6151
R959 B.n217 B.n214 10.6151
R960 B.n218 B.n217 10.6151
R961 B.n221 B.n218 10.6151
R962 B.n222 B.n221 10.6151
R963 B.n225 B.n222 10.6151
R964 B.n226 B.n225 10.6151
R965 B.n229 B.n226 10.6151
R966 B.n230 B.n229 10.6151
R967 B.n520 B.n230 10.6151
R968 B.n76 B.n75 10.2793
R969 B.n73 B.n72 10.2793
R970 B.n283 B.n282 10.2793
R971 B.n277 B.n276 10.2793
R972 B.n555 B.n0 8.11757
R973 B.n555 B.n1 8.11757
R974 B.n388 B.n387 6.5566
R975 B.n371 B.n370 6.5566
R976 B.n146 B.n145 6.5566
R977 B.n162 B.n74 6.5566
R978 B.n497 B.t3 5.88482
R979 B.n547 B.t0 5.88482
R980 B.n389 B.n388 4.05904
R981 B.n370 B.n369 4.05904
R982 B.n145 B.n144 4.05904
R983 B.n165 B.n74 4.05904
R984 VP.n7 VP.t3 1363.99
R985 VP.n5 VP.t2 1363.99
R986 VP.n0 VP.t1 1363.99
R987 VP.n2 VP.t5 1363.99
R988 VP.n6 VP.t4 1323.09
R989 VP.n1 VP.t0 1323.09
R990 VP.n3 VP.n0 161.489
R991 VP.n8 VP.n7 161.3
R992 VP.n3 VP.n2 161.3
R993 VP.n5 VP.n4 161.3
R994 VP.n4 VP.n3 37.5497
R995 VP.n6 VP.n5 36.5157
R996 VP.n7 VP.n6 36.5157
R997 VP.n1 VP.n0 36.5157
R998 VP.n2 VP.n1 36.5157
R999 VP.n8 VP.n4 0.189894
R1000 VP VP.n8 0.0516364
R1001 VDD1 VDD1.t4 66.8099
R1002 VDD1.n1 VDD1.t3 66.6962
R1003 VDD1.n1 VDD1.n0 64.4223
R1004 VDD1.n3 VDD1.n2 64.3635
R1005 VDD1.n3 VDD1.n1 34.3565
R1006 VDD1.n2 VDD1.t5 2.04595
R1007 VDD1.n2 VDD1.t0 2.04595
R1008 VDD1.n0 VDD1.t1 2.04595
R1009 VDD1.n0 VDD1.t2 2.04595
R1010 VDD1 VDD1.n3 0.0565345
C0 VN VP 4.16402f
C1 VP VDD1 1.9007f
C2 VDD2 VP 0.255214f
C3 VTAIL VN 1.38225f
C4 VTAIL VDD1 13.4097f
C5 VTAIL VDD2 13.4397f
C6 VTAIL VP 1.39692f
C7 VN VDD1 0.147569f
C8 VDD2 VN 1.79734f
C9 VDD2 VDD1 0.534787f
C10 VDD2 B 3.679815f
C11 VDD1 B 3.875849f
C12 VTAIL B 5.116941f
C13 VN B 5.38596f
C14 VP B 4.090747f
C15 VDD1.t4 B 2.30433f
C16 VDD1.t3 B 2.30373f
C17 VDD1.t1 B 0.205665f
C18 VDD1.t2 B 0.205665f
C19 VDD1.n0 B 1.80833f
C20 VDD1.n1 B 1.91528f
C21 VDD1.t5 B 0.205665f
C22 VDD1.t0 B 0.205665f
C23 VDD1.n2 B 1.80807f
C24 VDD1.n3 B 2.07054f
C25 VP.t1 B 0.194901f
C26 VP.n0 B 0.092274f
C27 VP.t0 B 0.19243f
C28 VP.n1 B 0.082836f
C29 VP.t5 B 0.194901f
C30 VP.n2 B 0.092227f
C31 VP.n3 B 1.23358f
C32 VP.n4 B 1.2266f
C33 VP.t4 B 0.19243f
C34 VP.t2 B 0.194901f
C35 VP.n5 B 0.092227f
C36 VP.n6 B 0.082836f
C37 VP.t3 B 0.194901f
C38 VP.n7 B 0.092227f
C39 VP.n8 B 0.027205f
C40 VTAIL.t3 B 0.220931f
C41 VTAIL.t8 B 0.220931f
C42 VTAIL.n0 B 1.86257f
C43 VTAIL.n1 B 0.354886f
C44 VTAIL.t10 B 2.3728f
C45 VTAIL.n2 B 0.473673f
C46 VTAIL.t1 B 0.220931f
C47 VTAIL.t9 B 0.220931f
C48 VTAIL.n3 B 1.86257f
C49 VTAIL.n4 B 1.57035f
C50 VTAIL.t7 B 0.220931f
C51 VTAIL.t6 B 0.220931f
C52 VTAIL.n5 B 1.86258f
C53 VTAIL.n6 B 1.57035f
C54 VTAIL.t5 B 2.37282f
C55 VTAIL.n7 B 0.473657f
C56 VTAIL.t0 B 0.220931f
C57 VTAIL.t11 B 0.220931f
C58 VTAIL.n8 B 1.86258f
C59 VTAIL.n9 B 0.381356f
C60 VTAIL.t2 B 2.3728f
C61 VTAIL.n10 B 1.62014f
C62 VTAIL.t4 B 2.3728f
C63 VTAIL.n11 B 1.6041f
C64 VDD2.t5 B 2.32093f
C65 VDD2.t2 B 0.2072f
C66 VDD2.t3 B 0.2072f
C67 VDD2.n0 B 1.82183f
C68 VDD2.n1 B 1.85878f
C69 VDD2.t0 B 2.31954f
C70 VDD2.n2 B 2.11409f
C71 VDD2.t1 B 0.2072f
C72 VDD2.t4 B 0.2072f
C73 VDD2.n3 B 1.82181f
C74 VN.t5 B 0.192637f
C75 VN.n0 B 0.091203f
C76 VN.t0 B 0.190195f
C77 VN.n1 B 0.081873f
C78 VN.t4 B 0.192637f
C79 VN.n2 B 0.091155f
C80 VN.n3 B 0.0671f
C81 VN.t3 B 0.192637f
C82 VN.n4 B 0.091203f
C83 VN.t1 B 0.192637f
C84 VN.t2 B 0.190195f
C85 VN.n5 B 0.081873f
C86 VN.n6 B 0.091155f
C87 VN.n7 B 1.2422f
.ends

