* NGSPICE file created from diff_pair_sample_0176.ext - technology: sky130A

.subckt diff_pair_sample_0176 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=3.4905 ps=18.68 w=8.95 l=3.68
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=0 ps=0 w=8.95 l=3.68
X2 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=3.4905 ps=18.68 w=8.95 l=3.68
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=0 ps=0 w=8.95 l=3.68
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=0 ps=0 w=8.95 l=3.68
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=3.4905 ps=18.68 w=8.95 l=3.68
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=3.4905 ps=18.68 w=8.95 l=3.68
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4905 pd=18.68 as=0 ps=0 w=8.95 l=3.68
R0 VP.n0 VP.t1 138.861
R1 VP.n0 VP.t0 93.6504
R2 VP VP.n0 0.621237
R3 VTAIL.n1 VTAIL.t0 50.1014
R4 VTAIL.n3 VTAIL.t1 50.1011
R5 VTAIL.n0 VTAIL.t2 50.1011
R6 VTAIL.n2 VTAIL.t3 50.1011
R7 VTAIL.n1 VTAIL.n0 26.9962
R8 VTAIL.n3 VTAIL.n2 23.5393
R9 VTAIL.n2 VTAIL.n1 2.19878
R10 VTAIL VTAIL.n0 1.39274
R11 VTAIL VTAIL.n3 0.806535
R12 VDD1 VDD1.t1 106.457
R13 VDD1 VDD1.t0 67.7023
R14 B.n634 B.n633 585
R15 B.n635 B.n634 585
R16 B.n247 B.n97 585
R17 B.n246 B.n245 585
R18 B.n244 B.n243 585
R19 B.n242 B.n241 585
R20 B.n240 B.n239 585
R21 B.n238 B.n237 585
R22 B.n236 B.n235 585
R23 B.n234 B.n233 585
R24 B.n232 B.n231 585
R25 B.n230 B.n229 585
R26 B.n228 B.n227 585
R27 B.n226 B.n225 585
R28 B.n224 B.n223 585
R29 B.n222 B.n221 585
R30 B.n220 B.n219 585
R31 B.n218 B.n217 585
R32 B.n216 B.n215 585
R33 B.n214 B.n213 585
R34 B.n212 B.n211 585
R35 B.n210 B.n209 585
R36 B.n208 B.n207 585
R37 B.n206 B.n205 585
R38 B.n204 B.n203 585
R39 B.n202 B.n201 585
R40 B.n200 B.n199 585
R41 B.n198 B.n197 585
R42 B.n196 B.n195 585
R43 B.n194 B.n193 585
R44 B.n192 B.n191 585
R45 B.n190 B.n189 585
R46 B.n188 B.n187 585
R47 B.n186 B.n185 585
R48 B.n184 B.n183 585
R49 B.n182 B.n181 585
R50 B.n180 B.n179 585
R51 B.n178 B.n177 585
R52 B.n176 B.n175 585
R53 B.n174 B.n173 585
R54 B.n172 B.n171 585
R55 B.n170 B.n169 585
R56 B.n168 B.n167 585
R57 B.n165 B.n164 585
R58 B.n163 B.n162 585
R59 B.n161 B.n160 585
R60 B.n159 B.n158 585
R61 B.n157 B.n156 585
R62 B.n155 B.n154 585
R63 B.n153 B.n152 585
R64 B.n151 B.n150 585
R65 B.n149 B.n148 585
R66 B.n147 B.n146 585
R67 B.n145 B.n144 585
R68 B.n143 B.n142 585
R69 B.n141 B.n140 585
R70 B.n139 B.n138 585
R71 B.n137 B.n136 585
R72 B.n135 B.n134 585
R73 B.n133 B.n132 585
R74 B.n131 B.n130 585
R75 B.n129 B.n128 585
R76 B.n127 B.n126 585
R77 B.n125 B.n124 585
R78 B.n123 B.n122 585
R79 B.n121 B.n120 585
R80 B.n119 B.n118 585
R81 B.n117 B.n116 585
R82 B.n115 B.n114 585
R83 B.n113 B.n112 585
R84 B.n111 B.n110 585
R85 B.n109 B.n108 585
R86 B.n107 B.n106 585
R87 B.n105 B.n104 585
R88 B.n60 B.n59 585
R89 B.n638 B.n637 585
R90 B.n632 B.n98 585
R91 B.n98 B.n57 585
R92 B.n631 B.n56 585
R93 B.n642 B.n56 585
R94 B.n630 B.n55 585
R95 B.n643 B.n55 585
R96 B.n629 B.n54 585
R97 B.n644 B.n54 585
R98 B.n628 B.n627 585
R99 B.n627 B.n50 585
R100 B.n626 B.n49 585
R101 B.n650 B.n49 585
R102 B.n625 B.n48 585
R103 B.n651 B.n48 585
R104 B.n624 B.n47 585
R105 B.n652 B.n47 585
R106 B.n623 B.n622 585
R107 B.n622 B.n43 585
R108 B.n621 B.n42 585
R109 B.t3 B.n42 585
R110 B.n620 B.n41 585
R111 B.n658 B.n41 585
R112 B.n619 B.n40 585
R113 B.n659 B.n40 585
R114 B.n618 B.n617 585
R115 B.n617 B.n36 585
R116 B.n616 B.n35 585
R117 B.n665 B.n35 585
R118 B.n615 B.n34 585
R119 B.n666 B.n34 585
R120 B.n614 B.n33 585
R121 B.n667 B.n33 585
R122 B.n613 B.n612 585
R123 B.n612 B.n29 585
R124 B.n611 B.n28 585
R125 B.n673 B.n28 585
R126 B.n610 B.n27 585
R127 B.n674 B.n27 585
R128 B.n609 B.n26 585
R129 B.n675 B.n26 585
R130 B.n608 B.n607 585
R131 B.n607 B.n22 585
R132 B.n606 B.n21 585
R133 B.n681 B.n21 585
R134 B.n605 B.n20 585
R135 B.n682 B.n20 585
R136 B.n604 B.n19 585
R137 B.n683 B.n19 585
R138 B.n603 B.n602 585
R139 B.n602 B.t1 585
R140 B.n601 B.n15 585
R141 B.n689 B.n15 585
R142 B.n600 B.n14 585
R143 B.n690 B.n14 585
R144 B.n599 B.n13 585
R145 B.n691 B.n13 585
R146 B.n598 B.n597 585
R147 B.n597 B.n12 585
R148 B.n596 B.n595 585
R149 B.n596 B.n8 585
R150 B.n594 B.n7 585
R151 B.n698 B.n7 585
R152 B.n593 B.n6 585
R153 B.n699 B.n6 585
R154 B.n592 B.n5 585
R155 B.n700 B.n5 585
R156 B.n591 B.n590 585
R157 B.n590 B.n4 585
R158 B.n589 B.n248 585
R159 B.n589 B.n588 585
R160 B.n579 B.n249 585
R161 B.n250 B.n249 585
R162 B.n581 B.n580 585
R163 B.n582 B.n581 585
R164 B.n578 B.n255 585
R165 B.n255 B.n254 585
R166 B.n577 B.n576 585
R167 B.n576 B.n575 585
R168 B.n257 B.n256 585
R169 B.t0 B.n257 585
R170 B.n568 B.n567 585
R171 B.n569 B.n568 585
R172 B.n566 B.n262 585
R173 B.n262 B.n261 585
R174 B.n565 B.n564 585
R175 B.n564 B.n563 585
R176 B.n264 B.n263 585
R177 B.n265 B.n264 585
R178 B.n556 B.n555 585
R179 B.n557 B.n556 585
R180 B.n554 B.n270 585
R181 B.n270 B.n269 585
R182 B.n553 B.n552 585
R183 B.n552 B.n551 585
R184 B.n272 B.n271 585
R185 B.n273 B.n272 585
R186 B.n544 B.n543 585
R187 B.n545 B.n544 585
R188 B.n542 B.n278 585
R189 B.n278 B.n277 585
R190 B.n541 B.n540 585
R191 B.n540 B.n539 585
R192 B.n280 B.n279 585
R193 B.n281 B.n280 585
R194 B.n532 B.n531 585
R195 B.n533 B.n532 585
R196 B.n530 B.n286 585
R197 B.n286 B.n285 585
R198 B.n529 B.n528 585
R199 B.n528 B.t7 585
R200 B.n288 B.n287 585
R201 B.n289 B.n288 585
R202 B.n521 B.n520 585
R203 B.n522 B.n521 585
R204 B.n519 B.n294 585
R205 B.n294 B.n293 585
R206 B.n518 B.n517 585
R207 B.n517 B.n516 585
R208 B.n296 B.n295 585
R209 B.n297 B.n296 585
R210 B.n509 B.n508 585
R211 B.n510 B.n509 585
R212 B.n507 B.n302 585
R213 B.n302 B.n301 585
R214 B.n506 B.n505 585
R215 B.n505 B.n504 585
R216 B.n304 B.n303 585
R217 B.n305 B.n304 585
R218 B.n500 B.n499 585
R219 B.n308 B.n307 585
R220 B.n496 B.n495 585
R221 B.n497 B.n496 585
R222 B.n494 B.n345 585
R223 B.n493 B.n492 585
R224 B.n491 B.n490 585
R225 B.n489 B.n488 585
R226 B.n487 B.n486 585
R227 B.n485 B.n484 585
R228 B.n483 B.n482 585
R229 B.n481 B.n480 585
R230 B.n479 B.n478 585
R231 B.n477 B.n476 585
R232 B.n475 B.n474 585
R233 B.n473 B.n472 585
R234 B.n471 B.n470 585
R235 B.n469 B.n468 585
R236 B.n467 B.n466 585
R237 B.n465 B.n464 585
R238 B.n463 B.n462 585
R239 B.n461 B.n460 585
R240 B.n459 B.n458 585
R241 B.n457 B.n456 585
R242 B.n455 B.n454 585
R243 B.n453 B.n452 585
R244 B.n451 B.n450 585
R245 B.n449 B.n448 585
R246 B.n447 B.n446 585
R247 B.n445 B.n444 585
R248 B.n443 B.n442 585
R249 B.n441 B.n440 585
R250 B.n439 B.n438 585
R251 B.n437 B.n436 585
R252 B.n435 B.n434 585
R253 B.n433 B.n432 585
R254 B.n431 B.n430 585
R255 B.n429 B.n428 585
R256 B.n427 B.n426 585
R257 B.n425 B.n424 585
R258 B.n423 B.n422 585
R259 B.n421 B.n420 585
R260 B.n419 B.n418 585
R261 B.n416 B.n415 585
R262 B.n414 B.n413 585
R263 B.n412 B.n411 585
R264 B.n410 B.n409 585
R265 B.n408 B.n407 585
R266 B.n406 B.n405 585
R267 B.n404 B.n403 585
R268 B.n402 B.n401 585
R269 B.n400 B.n399 585
R270 B.n398 B.n397 585
R271 B.n396 B.n395 585
R272 B.n394 B.n393 585
R273 B.n392 B.n391 585
R274 B.n390 B.n389 585
R275 B.n388 B.n387 585
R276 B.n386 B.n385 585
R277 B.n384 B.n383 585
R278 B.n382 B.n381 585
R279 B.n380 B.n379 585
R280 B.n378 B.n377 585
R281 B.n376 B.n375 585
R282 B.n374 B.n373 585
R283 B.n372 B.n371 585
R284 B.n370 B.n369 585
R285 B.n368 B.n367 585
R286 B.n366 B.n365 585
R287 B.n364 B.n363 585
R288 B.n362 B.n361 585
R289 B.n360 B.n359 585
R290 B.n358 B.n357 585
R291 B.n356 B.n355 585
R292 B.n354 B.n353 585
R293 B.n352 B.n351 585
R294 B.n501 B.n306 585
R295 B.n306 B.n305 585
R296 B.n503 B.n502 585
R297 B.n504 B.n503 585
R298 B.n300 B.n299 585
R299 B.n301 B.n300 585
R300 B.n512 B.n511 585
R301 B.n511 B.n510 585
R302 B.n513 B.n298 585
R303 B.n298 B.n297 585
R304 B.n515 B.n514 585
R305 B.n516 B.n515 585
R306 B.n292 B.n291 585
R307 B.n293 B.n292 585
R308 B.n524 B.n523 585
R309 B.n523 B.n522 585
R310 B.n525 B.n290 585
R311 B.n290 B.n289 585
R312 B.n527 B.n526 585
R313 B.t7 B.n527 585
R314 B.n284 B.n283 585
R315 B.n285 B.n284 585
R316 B.n535 B.n534 585
R317 B.n534 B.n533 585
R318 B.n536 B.n282 585
R319 B.n282 B.n281 585
R320 B.n538 B.n537 585
R321 B.n539 B.n538 585
R322 B.n276 B.n275 585
R323 B.n277 B.n276 585
R324 B.n547 B.n546 585
R325 B.n546 B.n545 585
R326 B.n548 B.n274 585
R327 B.n274 B.n273 585
R328 B.n550 B.n549 585
R329 B.n551 B.n550 585
R330 B.n268 B.n267 585
R331 B.n269 B.n268 585
R332 B.n559 B.n558 585
R333 B.n558 B.n557 585
R334 B.n560 B.n266 585
R335 B.n266 B.n265 585
R336 B.n562 B.n561 585
R337 B.n563 B.n562 585
R338 B.n260 B.n259 585
R339 B.n261 B.n260 585
R340 B.n571 B.n570 585
R341 B.n570 B.n569 585
R342 B.n572 B.n258 585
R343 B.n258 B.t0 585
R344 B.n574 B.n573 585
R345 B.n575 B.n574 585
R346 B.n253 B.n252 585
R347 B.n254 B.n253 585
R348 B.n584 B.n583 585
R349 B.n583 B.n582 585
R350 B.n585 B.n251 585
R351 B.n251 B.n250 585
R352 B.n587 B.n586 585
R353 B.n588 B.n587 585
R354 B.n3 B.n0 585
R355 B.n4 B.n3 585
R356 B.n697 B.n1 585
R357 B.n698 B.n697 585
R358 B.n696 B.n695 585
R359 B.n696 B.n8 585
R360 B.n694 B.n9 585
R361 B.n12 B.n9 585
R362 B.n693 B.n692 585
R363 B.n692 B.n691 585
R364 B.n11 B.n10 585
R365 B.n690 B.n11 585
R366 B.n688 B.n687 585
R367 B.n689 B.n688 585
R368 B.n686 B.n16 585
R369 B.n16 B.t1 585
R370 B.n685 B.n684 585
R371 B.n684 B.n683 585
R372 B.n18 B.n17 585
R373 B.n682 B.n18 585
R374 B.n680 B.n679 585
R375 B.n681 B.n680 585
R376 B.n678 B.n23 585
R377 B.n23 B.n22 585
R378 B.n677 B.n676 585
R379 B.n676 B.n675 585
R380 B.n25 B.n24 585
R381 B.n674 B.n25 585
R382 B.n672 B.n671 585
R383 B.n673 B.n672 585
R384 B.n670 B.n30 585
R385 B.n30 B.n29 585
R386 B.n669 B.n668 585
R387 B.n668 B.n667 585
R388 B.n32 B.n31 585
R389 B.n666 B.n32 585
R390 B.n664 B.n663 585
R391 B.n665 B.n664 585
R392 B.n662 B.n37 585
R393 B.n37 B.n36 585
R394 B.n661 B.n660 585
R395 B.n660 B.n659 585
R396 B.n39 B.n38 585
R397 B.n658 B.n39 585
R398 B.n657 B.n656 585
R399 B.t3 B.n657 585
R400 B.n655 B.n44 585
R401 B.n44 B.n43 585
R402 B.n654 B.n653 585
R403 B.n653 B.n652 585
R404 B.n46 B.n45 585
R405 B.n651 B.n46 585
R406 B.n649 B.n648 585
R407 B.n650 B.n649 585
R408 B.n647 B.n51 585
R409 B.n51 B.n50 585
R410 B.n646 B.n645 585
R411 B.n645 B.n644 585
R412 B.n53 B.n52 585
R413 B.n643 B.n53 585
R414 B.n641 B.n640 585
R415 B.n642 B.n641 585
R416 B.n639 B.n58 585
R417 B.n58 B.n57 585
R418 B.n701 B.n700 585
R419 B.n699 B.n2 585
R420 B.n637 B.n58 521.33
R421 B.n634 B.n98 521.33
R422 B.n351 B.n304 521.33
R423 B.n499 B.n306 521.33
R424 B.n102 B.t13 267.861
R425 B.n99 B.t2 267.861
R426 B.n349 B.t6 267.861
R427 B.n346 B.t10 267.861
R428 B.n635 B.n96 256.663
R429 B.n635 B.n95 256.663
R430 B.n635 B.n94 256.663
R431 B.n635 B.n93 256.663
R432 B.n635 B.n92 256.663
R433 B.n635 B.n91 256.663
R434 B.n635 B.n90 256.663
R435 B.n635 B.n89 256.663
R436 B.n635 B.n88 256.663
R437 B.n635 B.n87 256.663
R438 B.n635 B.n86 256.663
R439 B.n635 B.n85 256.663
R440 B.n635 B.n84 256.663
R441 B.n635 B.n83 256.663
R442 B.n635 B.n82 256.663
R443 B.n635 B.n81 256.663
R444 B.n635 B.n80 256.663
R445 B.n635 B.n79 256.663
R446 B.n635 B.n78 256.663
R447 B.n635 B.n77 256.663
R448 B.n635 B.n76 256.663
R449 B.n635 B.n75 256.663
R450 B.n635 B.n74 256.663
R451 B.n635 B.n73 256.663
R452 B.n635 B.n72 256.663
R453 B.n635 B.n71 256.663
R454 B.n635 B.n70 256.663
R455 B.n635 B.n69 256.663
R456 B.n635 B.n68 256.663
R457 B.n635 B.n67 256.663
R458 B.n635 B.n66 256.663
R459 B.n635 B.n65 256.663
R460 B.n635 B.n64 256.663
R461 B.n635 B.n63 256.663
R462 B.n635 B.n62 256.663
R463 B.n635 B.n61 256.663
R464 B.n636 B.n635 256.663
R465 B.n498 B.n497 256.663
R466 B.n497 B.n309 256.663
R467 B.n497 B.n310 256.663
R468 B.n497 B.n311 256.663
R469 B.n497 B.n312 256.663
R470 B.n497 B.n313 256.663
R471 B.n497 B.n314 256.663
R472 B.n497 B.n315 256.663
R473 B.n497 B.n316 256.663
R474 B.n497 B.n317 256.663
R475 B.n497 B.n318 256.663
R476 B.n497 B.n319 256.663
R477 B.n497 B.n320 256.663
R478 B.n497 B.n321 256.663
R479 B.n497 B.n322 256.663
R480 B.n497 B.n323 256.663
R481 B.n497 B.n324 256.663
R482 B.n497 B.n325 256.663
R483 B.n497 B.n326 256.663
R484 B.n497 B.n327 256.663
R485 B.n497 B.n328 256.663
R486 B.n497 B.n329 256.663
R487 B.n497 B.n330 256.663
R488 B.n497 B.n331 256.663
R489 B.n497 B.n332 256.663
R490 B.n497 B.n333 256.663
R491 B.n497 B.n334 256.663
R492 B.n497 B.n335 256.663
R493 B.n497 B.n336 256.663
R494 B.n497 B.n337 256.663
R495 B.n497 B.n338 256.663
R496 B.n497 B.n339 256.663
R497 B.n497 B.n340 256.663
R498 B.n497 B.n341 256.663
R499 B.n497 B.n342 256.663
R500 B.n497 B.n343 256.663
R501 B.n497 B.n344 256.663
R502 B.n703 B.n702 256.663
R503 B.n104 B.n60 163.367
R504 B.n108 B.n107 163.367
R505 B.n112 B.n111 163.367
R506 B.n116 B.n115 163.367
R507 B.n120 B.n119 163.367
R508 B.n124 B.n123 163.367
R509 B.n128 B.n127 163.367
R510 B.n132 B.n131 163.367
R511 B.n136 B.n135 163.367
R512 B.n140 B.n139 163.367
R513 B.n144 B.n143 163.367
R514 B.n148 B.n147 163.367
R515 B.n152 B.n151 163.367
R516 B.n156 B.n155 163.367
R517 B.n160 B.n159 163.367
R518 B.n164 B.n163 163.367
R519 B.n169 B.n168 163.367
R520 B.n173 B.n172 163.367
R521 B.n177 B.n176 163.367
R522 B.n181 B.n180 163.367
R523 B.n185 B.n184 163.367
R524 B.n189 B.n188 163.367
R525 B.n193 B.n192 163.367
R526 B.n197 B.n196 163.367
R527 B.n201 B.n200 163.367
R528 B.n205 B.n204 163.367
R529 B.n209 B.n208 163.367
R530 B.n213 B.n212 163.367
R531 B.n217 B.n216 163.367
R532 B.n221 B.n220 163.367
R533 B.n225 B.n224 163.367
R534 B.n229 B.n228 163.367
R535 B.n233 B.n232 163.367
R536 B.n237 B.n236 163.367
R537 B.n241 B.n240 163.367
R538 B.n245 B.n244 163.367
R539 B.n634 B.n97 163.367
R540 B.n505 B.n304 163.367
R541 B.n505 B.n302 163.367
R542 B.n509 B.n302 163.367
R543 B.n509 B.n296 163.367
R544 B.n517 B.n296 163.367
R545 B.n517 B.n294 163.367
R546 B.n521 B.n294 163.367
R547 B.n521 B.n288 163.367
R548 B.n528 B.n288 163.367
R549 B.n528 B.n286 163.367
R550 B.n532 B.n286 163.367
R551 B.n532 B.n280 163.367
R552 B.n540 B.n280 163.367
R553 B.n540 B.n278 163.367
R554 B.n544 B.n278 163.367
R555 B.n544 B.n272 163.367
R556 B.n552 B.n272 163.367
R557 B.n552 B.n270 163.367
R558 B.n556 B.n270 163.367
R559 B.n556 B.n264 163.367
R560 B.n564 B.n264 163.367
R561 B.n564 B.n262 163.367
R562 B.n568 B.n262 163.367
R563 B.n568 B.n257 163.367
R564 B.n576 B.n257 163.367
R565 B.n576 B.n255 163.367
R566 B.n581 B.n255 163.367
R567 B.n581 B.n249 163.367
R568 B.n589 B.n249 163.367
R569 B.n590 B.n589 163.367
R570 B.n590 B.n5 163.367
R571 B.n6 B.n5 163.367
R572 B.n7 B.n6 163.367
R573 B.n596 B.n7 163.367
R574 B.n597 B.n596 163.367
R575 B.n597 B.n13 163.367
R576 B.n14 B.n13 163.367
R577 B.n15 B.n14 163.367
R578 B.n602 B.n15 163.367
R579 B.n602 B.n19 163.367
R580 B.n20 B.n19 163.367
R581 B.n21 B.n20 163.367
R582 B.n607 B.n21 163.367
R583 B.n607 B.n26 163.367
R584 B.n27 B.n26 163.367
R585 B.n28 B.n27 163.367
R586 B.n612 B.n28 163.367
R587 B.n612 B.n33 163.367
R588 B.n34 B.n33 163.367
R589 B.n35 B.n34 163.367
R590 B.n617 B.n35 163.367
R591 B.n617 B.n40 163.367
R592 B.n41 B.n40 163.367
R593 B.n42 B.n41 163.367
R594 B.n622 B.n42 163.367
R595 B.n622 B.n47 163.367
R596 B.n48 B.n47 163.367
R597 B.n49 B.n48 163.367
R598 B.n627 B.n49 163.367
R599 B.n627 B.n54 163.367
R600 B.n55 B.n54 163.367
R601 B.n56 B.n55 163.367
R602 B.n98 B.n56 163.367
R603 B.n496 B.n308 163.367
R604 B.n496 B.n345 163.367
R605 B.n492 B.n491 163.367
R606 B.n488 B.n487 163.367
R607 B.n484 B.n483 163.367
R608 B.n480 B.n479 163.367
R609 B.n476 B.n475 163.367
R610 B.n472 B.n471 163.367
R611 B.n468 B.n467 163.367
R612 B.n464 B.n463 163.367
R613 B.n460 B.n459 163.367
R614 B.n456 B.n455 163.367
R615 B.n452 B.n451 163.367
R616 B.n448 B.n447 163.367
R617 B.n444 B.n443 163.367
R618 B.n440 B.n439 163.367
R619 B.n436 B.n435 163.367
R620 B.n432 B.n431 163.367
R621 B.n428 B.n427 163.367
R622 B.n424 B.n423 163.367
R623 B.n420 B.n419 163.367
R624 B.n415 B.n414 163.367
R625 B.n411 B.n410 163.367
R626 B.n407 B.n406 163.367
R627 B.n403 B.n402 163.367
R628 B.n399 B.n398 163.367
R629 B.n395 B.n394 163.367
R630 B.n391 B.n390 163.367
R631 B.n387 B.n386 163.367
R632 B.n383 B.n382 163.367
R633 B.n379 B.n378 163.367
R634 B.n375 B.n374 163.367
R635 B.n371 B.n370 163.367
R636 B.n367 B.n366 163.367
R637 B.n363 B.n362 163.367
R638 B.n359 B.n358 163.367
R639 B.n355 B.n354 163.367
R640 B.n503 B.n306 163.367
R641 B.n503 B.n300 163.367
R642 B.n511 B.n300 163.367
R643 B.n511 B.n298 163.367
R644 B.n515 B.n298 163.367
R645 B.n515 B.n292 163.367
R646 B.n523 B.n292 163.367
R647 B.n523 B.n290 163.367
R648 B.n527 B.n290 163.367
R649 B.n527 B.n284 163.367
R650 B.n534 B.n284 163.367
R651 B.n534 B.n282 163.367
R652 B.n538 B.n282 163.367
R653 B.n538 B.n276 163.367
R654 B.n546 B.n276 163.367
R655 B.n546 B.n274 163.367
R656 B.n550 B.n274 163.367
R657 B.n550 B.n268 163.367
R658 B.n558 B.n268 163.367
R659 B.n558 B.n266 163.367
R660 B.n562 B.n266 163.367
R661 B.n562 B.n260 163.367
R662 B.n570 B.n260 163.367
R663 B.n570 B.n258 163.367
R664 B.n574 B.n258 163.367
R665 B.n574 B.n253 163.367
R666 B.n583 B.n253 163.367
R667 B.n583 B.n251 163.367
R668 B.n587 B.n251 163.367
R669 B.n587 B.n3 163.367
R670 B.n701 B.n3 163.367
R671 B.n697 B.n2 163.367
R672 B.n697 B.n696 163.367
R673 B.n696 B.n9 163.367
R674 B.n692 B.n9 163.367
R675 B.n692 B.n11 163.367
R676 B.n688 B.n11 163.367
R677 B.n688 B.n16 163.367
R678 B.n684 B.n16 163.367
R679 B.n684 B.n18 163.367
R680 B.n680 B.n18 163.367
R681 B.n680 B.n23 163.367
R682 B.n676 B.n23 163.367
R683 B.n676 B.n25 163.367
R684 B.n672 B.n25 163.367
R685 B.n672 B.n30 163.367
R686 B.n668 B.n30 163.367
R687 B.n668 B.n32 163.367
R688 B.n664 B.n32 163.367
R689 B.n664 B.n37 163.367
R690 B.n660 B.n37 163.367
R691 B.n660 B.n39 163.367
R692 B.n657 B.n39 163.367
R693 B.n657 B.n44 163.367
R694 B.n653 B.n44 163.367
R695 B.n653 B.n46 163.367
R696 B.n649 B.n46 163.367
R697 B.n649 B.n51 163.367
R698 B.n645 B.n51 163.367
R699 B.n645 B.n53 163.367
R700 B.n641 B.n53 163.367
R701 B.n641 B.n58 163.367
R702 B.n99 B.t4 148.25
R703 B.n349 B.t9 148.25
R704 B.n102 B.t14 148.24
R705 B.n346 B.t12 148.24
R706 B.n497 B.n305 105.941
R707 B.n635 B.n57 105.941
R708 B.n103 B.n102 77.7702
R709 B.n100 B.n99 77.7702
R710 B.n350 B.n349 77.7702
R711 B.n347 B.n346 77.7702
R712 B.n637 B.n636 71.676
R713 B.n104 B.n61 71.676
R714 B.n108 B.n62 71.676
R715 B.n112 B.n63 71.676
R716 B.n116 B.n64 71.676
R717 B.n120 B.n65 71.676
R718 B.n124 B.n66 71.676
R719 B.n128 B.n67 71.676
R720 B.n132 B.n68 71.676
R721 B.n136 B.n69 71.676
R722 B.n140 B.n70 71.676
R723 B.n144 B.n71 71.676
R724 B.n148 B.n72 71.676
R725 B.n152 B.n73 71.676
R726 B.n156 B.n74 71.676
R727 B.n160 B.n75 71.676
R728 B.n164 B.n76 71.676
R729 B.n169 B.n77 71.676
R730 B.n173 B.n78 71.676
R731 B.n177 B.n79 71.676
R732 B.n181 B.n80 71.676
R733 B.n185 B.n81 71.676
R734 B.n189 B.n82 71.676
R735 B.n193 B.n83 71.676
R736 B.n197 B.n84 71.676
R737 B.n201 B.n85 71.676
R738 B.n205 B.n86 71.676
R739 B.n209 B.n87 71.676
R740 B.n213 B.n88 71.676
R741 B.n217 B.n89 71.676
R742 B.n221 B.n90 71.676
R743 B.n225 B.n91 71.676
R744 B.n229 B.n92 71.676
R745 B.n233 B.n93 71.676
R746 B.n237 B.n94 71.676
R747 B.n241 B.n95 71.676
R748 B.n245 B.n96 71.676
R749 B.n97 B.n96 71.676
R750 B.n244 B.n95 71.676
R751 B.n240 B.n94 71.676
R752 B.n236 B.n93 71.676
R753 B.n232 B.n92 71.676
R754 B.n228 B.n91 71.676
R755 B.n224 B.n90 71.676
R756 B.n220 B.n89 71.676
R757 B.n216 B.n88 71.676
R758 B.n212 B.n87 71.676
R759 B.n208 B.n86 71.676
R760 B.n204 B.n85 71.676
R761 B.n200 B.n84 71.676
R762 B.n196 B.n83 71.676
R763 B.n192 B.n82 71.676
R764 B.n188 B.n81 71.676
R765 B.n184 B.n80 71.676
R766 B.n180 B.n79 71.676
R767 B.n176 B.n78 71.676
R768 B.n172 B.n77 71.676
R769 B.n168 B.n76 71.676
R770 B.n163 B.n75 71.676
R771 B.n159 B.n74 71.676
R772 B.n155 B.n73 71.676
R773 B.n151 B.n72 71.676
R774 B.n147 B.n71 71.676
R775 B.n143 B.n70 71.676
R776 B.n139 B.n69 71.676
R777 B.n135 B.n68 71.676
R778 B.n131 B.n67 71.676
R779 B.n127 B.n66 71.676
R780 B.n123 B.n65 71.676
R781 B.n119 B.n64 71.676
R782 B.n115 B.n63 71.676
R783 B.n111 B.n62 71.676
R784 B.n107 B.n61 71.676
R785 B.n636 B.n60 71.676
R786 B.n499 B.n498 71.676
R787 B.n345 B.n309 71.676
R788 B.n491 B.n310 71.676
R789 B.n487 B.n311 71.676
R790 B.n483 B.n312 71.676
R791 B.n479 B.n313 71.676
R792 B.n475 B.n314 71.676
R793 B.n471 B.n315 71.676
R794 B.n467 B.n316 71.676
R795 B.n463 B.n317 71.676
R796 B.n459 B.n318 71.676
R797 B.n455 B.n319 71.676
R798 B.n451 B.n320 71.676
R799 B.n447 B.n321 71.676
R800 B.n443 B.n322 71.676
R801 B.n439 B.n323 71.676
R802 B.n435 B.n324 71.676
R803 B.n431 B.n325 71.676
R804 B.n427 B.n326 71.676
R805 B.n423 B.n327 71.676
R806 B.n419 B.n328 71.676
R807 B.n414 B.n329 71.676
R808 B.n410 B.n330 71.676
R809 B.n406 B.n331 71.676
R810 B.n402 B.n332 71.676
R811 B.n398 B.n333 71.676
R812 B.n394 B.n334 71.676
R813 B.n390 B.n335 71.676
R814 B.n386 B.n336 71.676
R815 B.n382 B.n337 71.676
R816 B.n378 B.n338 71.676
R817 B.n374 B.n339 71.676
R818 B.n370 B.n340 71.676
R819 B.n366 B.n341 71.676
R820 B.n362 B.n342 71.676
R821 B.n358 B.n343 71.676
R822 B.n354 B.n344 71.676
R823 B.n498 B.n308 71.676
R824 B.n492 B.n309 71.676
R825 B.n488 B.n310 71.676
R826 B.n484 B.n311 71.676
R827 B.n480 B.n312 71.676
R828 B.n476 B.n313 71.676
R829 B.n472 B.n314 71.676
R830 B.n468 B.n315 71.676
R831 B.n464 B.n316 71.676
R832 B.n460 B.n317 71.676
R833 B.n456 B.n318 71.676
R834 B.n452 B.n319 71.676
R835 B.n448 B.n320 71.676
R836 B.n444 B.n321 71.676
R837 B.n440 B.n322 71.676
R838 B.n436 B.n323 71.676
R839 B.n432 B.n324 71.676
R840 B.n428 B.n325 71.676
R841 B.n424 B.n326 71.676
R842 B.n420 B.n327 71.676
R843 B.n415 B.n328 71.676
R844 B.n411 B.n329 71.676
R845 B.n407 B.n330 71.676
R846 B.n403 B.n331 71.676
R847 B.n399 B.n332 71.676
R848 B.n395 B.n333 71.676
R849 B.n391 B.n334 71.676
R850 B.n387 B.n335 71.676
R851 B.n383 B.n336 71.676
R852 B.n379 B.n337 71.676
R853 B.n375 B.n338 71.676
R854 B.n371 B.n339 71.676
R855 B.n367 B.n340 71.676
R856 B.n363 B.n341 71.676
R857 B.n359 B.n342 71.676
R858 B.n355 B.n343 71.676
R859 B.n351 B.n344 71.676
R860 B.n702 B.n701 71.676
R861 B.n702 B.n2 71.676
R862 B.n100 B.t5 70.4812
R863 B.n350 B.t8 70.4812
R864 B.n103 B.t15 70.4704
R865 B.n347 B.t11 70.4704
R866 B.n166 B.n103 59.5399
R867 B.n101 B.n100 59.5399
R868 B.n417 B.n350 59.5399
R869 B.n348 B.n347 59.5399
R870 B.n504 B.n305 52.584
R871 B.n504 B.n301 52.584
R872 B.n510 B.n301 52.584
R873 B.n510 B.n297 52.584
R874 B.n516 B.n297 52.584
R875 B.n516 B.n293 52.584
R876 B.n522 B.n293 52.584
R877 B.n522 B.n289 52.584
R878 B.t7 B.n289 52.584
R879 B.t7 B.n285 52.584
R880 B.n533 B.n285 52.584
R881 B.n533 B.n281 52.584
R882 B.n539 B.n281 52.584
R883 B.n539 B.n277 52.584
R884 B.n545 B.n277 52.584
R885 B.n545 B.n273 52.584
R886 B.n551 B.n273 52.584
R887 B.n551 B.n269 52.584
R888 B.n557 B.n269 52.584
R889 B.n557 B.n265 52.584
R890 B.n563 B.n265 52.584
R891 B.n563 B.n261 52.584
R892 B.n569 B.n261 52.584
R893 B.n569 B.t0 52.584
R894 B.n575 B.t0 52.584
R895 B.n575 B.n254 52.584
R896 B.n582 B.n254 52.584
R897 B.n582 B.n250 52.584
R898 B.n588 B.n250 52.584
R899 B.n588 B.n4 52.584
R900 B.n700 B.n4 52.584
R901 B.n700 B.n699 52.584
R902 B.n699 B.n698 52.584
R903 B.n698 B.n8 52.584
R904 B.n12 B.n8 52.584
R905 B.n691 B.n12 52.584
R906 B.n691 B.n690 52.584
R907 B.n690 B.n689 52.584
R908 B.n689 B.t1 52.584
R909 B.n683 B.t1 52.584
R910 B.n683 B.n682 52.584
R911 B.n682 B.n681 52.584
R912 B.n681 B.n22 52.584
R913 B.n675 B.n22 52.584
R914 B.n675 B.n674 52.584
R915 B.n674 B.n673 52.584
R916 B.n673 B.n29 52.584
R917 B.n667 B.n29 52.584
R918 B.n667 B.n666 52.584
R919 B.n666 B.n665 52.584
R920 B.n665 B.n36 52.584
R921 B.n659 B.n36 52.584
R922 B.n659 B.n658 52.584
R923 B.n658 B.t3 52.584
R924 B.t3 B.n43 52.584
R925 B.n652 B.n43 52.584
R926 B.n652 B.n651 52.584
R927 B.n651 B.n650 52.584
R928 B.n650 B.n50 52.584
R929 B.n644 B.n50 52.584
R930 B.n644 B.n643 52.584
R931 B.n643 B.n642 52.584
R932 B.n642 B.n57 52.584
R933 B.n501 B.n500 33.8737
R934 B.n352 B.n303 33.8737
R935 B.n633 B.n632 33.8737
R936 B.n639 B.n638 33.8737
R937 B B.n703 18.0485
R938 B.n502 B.n501 10.6151
R939 B.n502 B.n299 10.6151
R940 B.n512 B.n299 10.6151
R941 B.n513 B.n512 10.6151
R942 B.n514 B.n513 10.6151
R943 B.n514 B.n291 10.6151
R944 B.n524 B.n291 10.6151
R945 B.n525 B.n524 10.6151
R946 B.n526 B.n525 10.6151
R947 B.n526 B.n283 10.6151
R948 B.n535 B.n283 10.6151
R949 B.n536 B.n535 10.6151
R950 B.n537 B.n536 10.6151
R951 B.n537 B.n275 10.6151
R952 B.n547 B.n275 10.6151
R953 B.n548 B.n547 10.6151
R954 B.n549 B.n548 10.6151
R955 B.n549 B.n267 10.6151
R956 B.n559 B.n267 10.6151
R957 B.n560 B.n559 10.6151
R958 B.n561 B.n560 10.6151
R959 B.n561 B.n259 10.6151
R960 B.n571 B.n259 10.6151
R961 B.n572 B.n571 10.6151
R962 B.n573 B.n572 10.6151
R963 B.n573 B.n252 10.6151
R964 B.n584 B.n252 10.6151
R965 B.n585 B.n584 10.6151
R966 B.n586 B.n585 10.6151
R967 B.n586 B.n0 10.6151
R968 B.n500 B.n307 10.6151
R969 B.n495 B.n307 10.6151
R970 B.n495 B.n494 10.6151
R971 B.n494 B.n493 10.6151
R972 B.n493 B.n490 10.6151
R973 B.n490 B.n489 10.6151
R974 B.n489 B.n486 10.6151
R975 B.n486 B.n485 10.6151
R976 B.n485 B.n482 10.6151
R977 B.n482 B.n481 10.6151
R978 B.n481 B.n478 10.6151
R979 B.n478 B.n477 10.6151
R980 B.n477 B.n474 10.6151
R981 B.n474 B.n473 10.6151
R982 B.n473 B.n470 10.6151
R983 B.n470 B.n469 10.6151
R984 B.n469 B.n466 10.6151
R985 B.n466 B.n465 10.6151
R986 B.n465 B.n462 10.6151
R987 B.n462 B.n461 10.6151
R988 B.n461 B.n458 10.6151
R989 B.n458 B.n457 10.6151
R990 B.n457 B.n454 10.6151
R991 B.n454 B.n453 10.6151
R992 B.n453 B.n450 10.6151
R993 B.n450 B.n449 10.6151
R994 B.n449 B.n446 10.6151
R995 B.n446 B.n445 10.6151
R996 B.n445 B.n442 10.6151
R997 B.n442 B.n441 10.6151
R998 B.n441 B.n438 10.6151
R999 B.n438 B.n437 10.6151
R1000 B.n434 B.n433 10.6151
R1001 B.n433 B.n430 10.6151
R1002 B.n430 B.n429 10.6151
R1003 B.n429 B.n426 10.6151
R1004 B.n426 B.n425 10.6151
R1005 B.n425 B.n422 10.6151
R1006 B.n422 B.n421 10.6151
R1007 B.n421 B.n418 10.6151
R1008 B.n416 B.n413 10.6151
R1009 B.n413 B.n412 10.6151
R1010 B.n412 B.n409 10.6151
R1011 B.n409 B.n408 10.6151
R1012 B.n408 B.n405 10.6151
R1013 B.n405 B.n404 10.6151
R1014 B.n404 B.n401 10.6151
R1015 B.n401 B.n400 10.6151
R1016 B.n400 B.n397 10.6151
R1017 B.n397 B.n396 10.6151
R1018 B.n396 B.n393 10.6151
R1019 B.n393 B.n392 10.6151
R1020 B.n392 B.n389 10.6151
R1021 B.n389 B.n388 10.6151
R1022 B.n388 B.n385 10.6151
R1023 B.n385 B.n384 10.6151
R1024 B.n384 B.n381 10.6151
R1025 B.n381 B.n380 10.6151
R1026 B.n380 B.n377 10.6151
R1027 B.n377 B.n376 10.6151
R1028 B.n376 B.n373 10.6151
R1029 B.n373 B.n372 10.6151
R1030 B.n372 B.n369 10.6151
R1031 B.n369 B.n368 10.6151
R1032 B.n368 B.n365 10.6151
R1033 B.n365 B.n364 10.6151
R1034 B.n364 B.n361 10.6151
R1035 B.n361 B.n360 10.6151
R1036 B.n360 B.n357 10.6151
R1037 B.n357 B.n356 10.6151
R1038 B.n356 B.n353 10.6151
R1039 B.n353 B.n352 10.6151
R1040 B.n506 B.n303 10.6151
R1041 B.n507 B.n506 10.6151
R1042 B.n508 B.n507 10.6151
R1043 B.n508 B.n295 10.6151
R1044 B.n518 B.n295 10.6151
R1045 B.n519 B.n518 10.6151
R1046 B.n520 B.n519 10.6151
R1047 B.n520 B.n287 10.6151
R1048 B.n529 B.n287 10.6151
R1049 B.n530 B.n529 10.6151
R1050 B.n531 B.n530 10.6151
R1051 B.n531 B.n279 10.6151
R1052 B.n541 B.n279 10.6151
R1053 B.n542 B.n541 10.6151
R1054 B.n543 B.n542 10.6151
R1055 B.n543 B.n271 10.6151
R1056 B.n553 B.n271 10.6151
R1057 B.n554 B.n553 10.6151
R1058 B.n555 B.n554 10.6151
R1059 B.n555 B.n263 10.6151
R1060 B.n565 B.n263 10.6151
R1061 B.n566 B.n565 10.6151
R1062 B.n567 B.n566 10.6151
R1063 B.n567 B.n256 10.6151
R1064 B.n577 B.n256 10.6151
R1065 B.n578 B.n577 10.6151
R1066 B.n580 B.n578 10.6151
R1067 B.n580 B.n579 10.6151
R1068 B.n579 B.n248 10.6151
R1069 B.n591 B.n248 10.6151
R1070 B.n592 B.n591 10.6151
R1071 B.n593 B.n592 10.6151
R1072 B.n594 B.n593 10.6151
R1073 B.n595 B.n594 10.6151
R1074 B.n598 B.n595 10.6151
R1075 B.n599 B.n598 10.6151
R1076 B.n600 B.n599 10.6151
R1077 B.n601 B.n600 10.6151
R1078 B.n603 B.n601 10.6151
R1079 B.n604 B.n603 10.6151
R1080 B.n605 B.n604 10.6151
R1081 B.n606 B.n605 10.6151
R1082 B.n608 B.n606 10.6151
R1083 B.n609 B.n608 10.6151
R1084 B.n610 B.n609 10.6151
R1085 B.n611 B.n610 10.6151
R1086 B.n613 B.n611 10.6151
R1087 B.n614 B.n613 10.6151
R1088 B.n615 B.n614 10.6151
R1089 B.n616 B.n615 10.6151
R1090 B.n618 B.n616 10.6151
R1091 B.n619 B.n618 10.6151
R1092 B.n620 B.n619 10.6151
R1093 B.n621 B.n620 10.6151
R1094 B.n623 B.n621 10.6151
R1095 B.n624 B.n623 10.6151
R1096 B.n625 B.n624 10.6151
R1097 B.n626 B.n625 10.6151
R1098 B.n628 B.n626 10.6151
R1099 B.n629 B.n628 10.6151
R1100 B.n630 B.n629 10.6151
R1101 B.n631 B.n630 10.6151
R1102 B.n632 B.n631 10.6151
R1103 B.n695 B.n1 10.6151
R1104 B.n695 B.n694 10.6151
R1105 B.n694 B.n693 10.6151
R1106 B.n693 B.n10 10.6151
R1107 B.n687 B.n10 10.6151
R1108 B.n687 B.n686 10.6151
R1109 B.n686 B.n685 10.6151
R1110 B.n685 B.n17 10.6151
R1111 B.n679 B.n17 10.6151
R1112 B.n679 B.n678 10.6151
R1113 B.n678 B.n677 10.6151
R1114 B.n677 B.n24 10.6151
R1115 B.n671 B.n24 10.6151
R1116 B.n671 B.n670 10.6151
R1117 B.n670 B.n669 10.6151
R1118 B.n669 B.n31 10.6151
R1119 B.n663 B.n31 10.6151
R1120 B.n663 B.n662 10.6151
R1121 B.n662 B.n661 10.6151
R1122 B.n661 B.n38 10.6151
R1123 B.n656 B.n38 10.6151
R1124 B.n656 B.n655 10.6151
R1125 B.n655 B.n654 10.6151
R1126 B.n654 B.n45 10.6151
R1127 B.n648 B.n45 10.6151
R1128 B.n648 B.n647 10.6151
R1129 B.n647 B.n646 10.6151
R1130 B.n646 B.n52 10.6151
R1131 B.n640 B.n52 10.6151
R1132 B.n640 B.n639 10.6151
R1133 B.n638 B.n59 10.6151
R1134 B.n105 B.n59 10.6151
R1135 B.n106 B.n105 10.6151
R1136 B.n109 B.n106 10.6151
R1137 B.n110 B.n109 10.6151
R1138 B.n113 B.n110 10.6151
R1139 B.n114 B.n113 10.6151
R1140 B.n117 B.n114 10.6151
R1141 B.n118 B.n117 10.6151
R1142 B.n121 B.n118 10.6151
R1143 B.n122 B.n121 10.6151
R1144 B.n125 B.n122 10.6151
R1145 B.n126 B.n125 10.6151
R1146 B.n129 B.n126 10.6151
R1147 B.n130 B.n129 10.6151
R1148 B.n133 B.n130 10.6151
R1149 B.n134 B.n133 10.6151
R1150 B.n137 B.n134 10.6151
R1151 B.n138 B.n137 10.6151
R1152 B.n141 B.n138 10.6151
R1153 B.n142 B.n141 10.6151
R1154 B.n145 B.n142 10.6151
R1155 B.n146 B.n145 10.6151
R1156 B.n149 B.n146 10.6151
R1157 B.n150 B.n149 10.6151
R1158 B.n153 B.n150 10.6151
R1159 B.n154 B.n153 10.6151
R1160 B.n157 B.n154 10.6151
R1161 B.n158 B.n157 10.6151
R1162 B.n161 B.n158 10.6151
R1163 B.n162 B.n161 10.6151
R1164 B.n165 B.n162 10.6151
R1165 B.n170 B.n167 10.6151
R1166 B.n171 B.n170 10.6151
R1167 B.n174 B.n171 10.6151
R1168 B.n175 B.n174 10.6151
R1169 B.n178 B.n175 10.6151
R1170 B.n179 B.n178 10.6151
R1171 B.n182 B.n179 10.6151
R1172 B.n183 B.n182 10.6151
R1173 B.n187 B.n186 10.6151
R1174 B.n190 B.n187 10.6151
R1175 B.n191 B.n190 10.6151
R1176 B.n194 B.n191 10.6151
R1177 B.n195 B.n194 10.6151
R1178 B.n198 B.n195 10.6151
R1179 B.n199 B.n198 10.6151
R1180 B.n202 B.n199 10.6151
R1181 B.n203 B.n202 10.6151
R1182 B.n206 B.n203 10.6151
R1183 B.n207 B.n206 10.6151
R1184 B.n210 B.n207 10.6151
R1185 B.n211 B.n210 10.6151
R1186 B.n214 B.n211 10.6151
R1187 B.n215 B.n214 10.6151
R1188 B.n218 B.n215 10.6151
R1189 B.n219 B.n218 10.6151
R1190 B.n222 B.n219 10.6151
R1191 B.n223 B.n222 10.6151
R1192 B.n226 B.n223 10.6151
R1193 B.n227 B.n226 10.6151
R1194 B.n230 B.n227 10.6151
R1195 B.n231 B.n230 10.6151
R1196 B.n234 B.n231 10.6151
R1197 B.n235 B.n234 10.6151
R1198 B.n238 B.n235 10.6151
R1199 B.n239 B.n238 10.6151
R1200 B.n242 B.n239 10.6151
R1201 B.n243 B.n242 10.6151
R1202 B.n246 B.n243 10.6151
R1203 B.n247 B.n246 10.6151
R1204 B.n633 B.n247 10.6151
R1205 B.n703 B.n0 8.11757
R1206 B.n703 B.n1 8.11757
R1207 B.n434 B.n348 6.5566
R1208 B.n418 B.n417 6.5566
R1209 B.n167 B.n166 6.5566
R1210 B.n183 B.n101 6.5566
R1211 B.n437 B.n348 4.05904
R1212 B.n417 B.n416 4.05904
R1213 B.n166 B.n165 4.05904
R1214 B.n186 B.n101 4.05904
R1215 VN VN.t1 138.673
R1216 VN VN.t0 94.2711
R1217 VDD2.n0 VDD2.t1 105.069
R1218 VDD2.n0 VDD2.t0 66.7799
R1219 VDD2 VDD2.n0 0.922914
C0 VDD2 VN 2.23523f
C1 VP VTAIL 2.12843f
C2 VDD1 VP 2.46315f
C3 VP VN 5.40181f
C4 VDD2 VP 0.378083f
C5 VDD1 VTAIL 4.52061f
C6 VN VTAIL 2.11405f
C7 VDD2 VTAIL 4.57984f
C8 VDD1 VN 0.148618f
C9 VDD2 VDD1 0.792503f
C10 VDD2 B 4.281538f
C11 VDD1 B 7.44561f
C12 VTAIL B 6.618596f
C13 VN B 11.156651f
C14 VP B 7.552954f
C15 VDD2.t1 B 2.14427f
C16 VDD2.t0 B 1.63354f
C17 VDD2.n0 B 2.84419f
C18 VN.t0 B 2.72057f
C19 VN.t1 B 3.399f
C20 VDD1.t0 B 1.66682f
C21 VDD1.t1 B 2.2247f
C22 VTAIL.t2 B 1.66723f
C23 VTAIL.n0 B 1.72365f
C24 VTAIL.t0 B 1.66723f
C25 VTAIL.n1 B 1.78122f
C26 VTAIL.t3 B 1.66723f
C27 VTAIL.n2 B 1.53432f
C28 VTAIL.t1 B 1.66723f
C29 VTAIL.n3 B 1.43488f
C30 VP.t1 B 3.51921f
C31 VP.t0 B 2.80955f
C32 VP.n0 B 3.56026f
.ends

