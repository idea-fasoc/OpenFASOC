* NGSPICE file created from diff_pair_sample_1634.ext - technology: sky130A

.subckt diff_pair_sample_1634 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=3.0228 ps=18.65 w=18.32 l=3.96
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=0 ps=0 w=18.32 l=3.96
X2 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0228 pd=18.65 as=7.1448 ps=37.42 w=18.32 l=3.96
X3 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=3.0228 ps=18.65 w=18.32 l=3.96
X4 VDD2.t3 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0228 pd=18.65 as=7.1448 ps=37.42 w=18.32 l=3.96
X5 VDD2.t0 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0228 pd=18.65 as=7.1448 ps=37.42 w=18.32 l=3.96
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=0 ps=0 w=18.32 l=3.96
X7 VTAIL.t4 VN.t3 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=3.0228 ps=18.65 w=18.32 l=3.96
X8 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=3.0228 ps=18.65 w=18.32 l=3.96
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=0 ps=0 w=18.32 l=3.96
X10 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0228 pd=18.65 as=7.1448 ps=37.42 w=18.32 l=3.96
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1448 pd=37.42 as=0 ps=0 w=18.32 l=3.96
R0 VN.n0 VN.t0 145.382
R1 VN.n1 VN.t2 145.382
R2 VN.n0 VN.t1 143.946
R3 VN.n1 VN.t3 143.946
R4 VN VN.n1 57.1655
R5 VN VN.n0 1.75264
R6 VDD2.n2 VDD2.n0 112.802
R7 VDD2.n2 VDD2.n1 62.1996
R8 VDD2.n1 VDD2.t1 1.08129
R9 VDD2.n1 VDD2.t0 1.08129
R10 VDD2.n0 VDD2.t2 1.08129
R11 VDD2.n0 VDD2.t3 1.08129
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n810 VTAIL.n714 289.615
R14 VTAIL.n96 VTAIL.n0 289.615
R15 VTAIL.n198 VTAIL.n102 289.615
R16 VTAIL.n300 VTAIL.n204 289.615
R17 VTAIL.n708 VTAIL.n612 289.615
R18 VTAIL.n606 VTAIL.n510 289.615
R19 VTAIL.n504 VTAIL.n408 289.615
R20 VTAIL.n402 VTAIL.n306 289.615
R21 VTAIL.n746 VTAIL.n745 185
R22 VTAIL.n751 VTAIL.n750 185
R23 VTAIL.n753 VTAIL.n752 185
R24 VTAIL.n742 VTAIL.n741 185
R25 VTAIL.n759 VTAIL.n758 185
R26 VTAIL.n761 VTAIL.n760 185
R27 VTAIL.n738 VTAIL.n737 185
R28 VTAIL.n767 VTAIL.n766 185
R29 VTAIL.n769 VTAIL.n768 185
R30 VTAIL.n734 VTAIL.n733 185
R31 VTAIL.n775 VTAIL.n774 185
R32 VTAIL.n777 VTAIL.n776 185
R33 VTAIL.n730 VTAIL.n729 185
R34 VTAIL.n783 VTAIL.n782 185
R35 VTAIL.n785 VTAIL.n784 185
R36 VTAIL.n726 VTAIL.n725 185
R37 VTAIL.n792 VTAIL.n791 185
R38 VTAIL.n793 VTAIL.n724 185
R39 VTAIL.n795 VTAIL.n794 185
R40 VTAIL.n722 VTAIL.n721 185
R41 VTAIL.n801 VTAIL.n800 185
R42 VTAIL.n803 VTAIL.n802 185
R43 VTAIL.n718 VTAIL.n717 185
R44 VTAIL.n809 VTAIL.n808 185
R45 VTAIL.n811 VTAIL.n810 185
R46 VTAIL.n32 VTAIL.n31 185
R47 VTAIL.n37 VTAIL.n36 185
R48 VTAIL.n39 VTAIL.n38 185
R49 VTAIL.n28 VTAIL.n27 185
R50 VTAIL.n45 VTAIL.n44 185
R51 VTAIL.n47 VTAIL.n46 185
R52 VTAIL.n24 VTAIL.n23 185
R53 VTAIL.n53 VTAIL.n52 185
R54 VTAIL.n55 VTAIL.n54 185
R55 VTAIL.n20 VTAIL.n19 185
R56 VTAIL.n61 VTAIL.n60 185
R57 VTAIL.n63 VTAIL.n62 185
R58 VTAIL.n16 VTAIL.n15 185
R59 VTAIL.n69 VTAIL.n68 185
R60 VTAIL.n71 VTAIL.n70 185
R61 VTAIL.n12 VTAIL.n11 185
R62 VTAIL.n78 VTAIL.n77 185
R63 VTAIL.n79 VTAIL.n10 185
R64 VTAIL.n81 VTAIL.n80 185
R65 VTAIL.n8 VTAIL.n7 185
R66 VTAIL.n87 VTAIL.n86 185
R67 VTAIL.n89 VTAIL.n88 185
R68 VTAIL.n4 VTAIL.n3 185
R69 VTAIL.n95 VTAIL.n94 185
R70 VTAIL.n97 VTAIL.n96 185
R71 VTAIL.n134 VTAIL.n133 185
R72 VTAIL.n139 VTAIL.n138 185
R73 VTAIL.n141 VTAIL.n140 185
R74 VTAIL.n130 VTAIL.n129 185
R75 VTAIL.n147 VTAIL.n146 185
R76 VTAIL.n149 VTAIL.n148 185
R77 VTAIL.n126 VTAIL.n125 185
R78 VTAIL.n155 VTAIL.n154 185
R79 VTAIL.n157 VTAIL.n156 185
R80 VTAIL.n122 VTAIL.n121 185
R81 VTAIL.n163 VTAIL.n162 185
R82 VTAIL.n165 VTAIL.n164 185
R83 VTAIL.n118 VTAIL.n117 185
R84 VTAIL.n171 VTAIL.n170 185
R85 VTAIL.n173 VTAIL.n172 185
R86 VTAIL.n114 VTAIL.n113 185
R87 VTAIL.n180 VTAIL.n179 185
R88 VTAIL.n181 VTAIL.n112 185
R89 VTAIL.n183 VTAIL.n182 185
R90 VTAIL.n110 VTAIL.n109 185
R91 VTAIL.n189 VTAIL.n188 185
R92 VTAIL.n191 VTAIL.n190 185
R93 VTAIL.n106 VTAIL.n105 185
R94 VTAIL.n197 VTAIL.n196 185
R95 VTAIL.n199 VTAIL.n198 185
R96 VTAIL.n236 VTAIL.n235 185
R97 VTAIL.n241 VTAIL.n240 185
R98 VTAIL.n243 VTAIL.n242 185
R99 VTAIL.n232 VTAIL.n231 185
R100 VTAIL.n249 VTAIL.n248 185
R101 VTAIL.n251 VTAIL.n250 185
R102 VTAIL.n228 VTAIL.n227 185
R103 VTAIL.n257 VTAIL.n256 185
R104 VTAIL.n259 VTAIL.n258 185
R105 VTAIL.n224 VTAIL.n223 185
R106 VTAIL.n265 VTAIL.n264 185
R107 VTAIL.n267 VTAIL.n266 185
R108 VTAIL.n220 VTAIL.n219 185
R109 VTAIL.n273 VTAIL.n272 185
R110 VTAIL.n275 VTAIL.n274 185
R111 VTAIL.n216 VTAIL.n215 185
R112 VTAIL.n282 VTAIL.n281 185
R113 VTAIL.n283 VTAIL.n214 185
R114 VTAIL.n285 VTAIL.n284 185
R115 VTAIL.n212 VTAIL.n211 185
R116 VTAIL.n291 VTAIL.n290 185
R117 VTAIL.n293 VTAIL.n292 185
R118 VTAIL.n208 VTAIL.n207 185
R119 VTAIL.n299 VTAIL.n298 185
R120 VTAIL.n301 VTAIL.n300 185
R121 VTAIL.n709 VTAIL.n708 185
R122 VTAIL.n707 VTAIL.n706 185
R123 VTAIL.n616 VTAIL.n615 185
R124 VTAIL.n701 VTAIL.n700 185
R125 VTAIL.n699 VTAIL.n698 185
R126 VTAIL.n620 VTAIL.n619 185
R127 VTAIL.n693 VTAIL.n692 185
R128 VTAIL.n691 VTAIL.n622 185
R129 VTAIL.n690 VTAIL.n689 185
R130 VTAIL.n625 VTAIL.n623 185
R131 VTAIL.n684 VTAIL.n683 185
R132 VTAIL.n682 VTAIL.n681 185
R133 VTAIL.n629 VTAIL.n628 185
R134 VTAIL.n676 VTAIL.n675 185
R135 VTAIL.n674 VTAIL.n673 185
R136 VTAIL.n633 VTAIL.n632 185
R137 VTAIL.n668 VTAIL.n667 185
R138 VTAIL.n666 VTAIL.n665 185
R139 VTAIL.n637 VTAIL.n636 185
R140 VTAIL.n660 VTAIL.n659 185
R141 VTAIL.n658 VTAIL.n657 185
R142 VTAIL.n641 VTAIL.n640 185
R143 VTAIL.n652 VTAIL.n651 185
R144 VTAIL.n650 VTAIL.n649 185
R145 VTAIL.n645 VTAIL.n644 185
R146 VTAIL.n607 VTAIL.n606 185
R147 VTAIL.n605 VTAIL.n604 185
R148 VTAIL.n514 VTAIL.n513 185
R149 VTAIL.n599 VTAIL.n598 185
R150 VTAIL.n597 VTAIL.n596 185
R151 VTAIL.n518 VTAIL.n517 185
R152 VTAIL.n591 VTAIL.n590 185
R153 VTAIL.n589 VTAIL.n520 185
R154 VTAIL.n588 VTAIL.n587 185
R155 VTAIL.n523 VTAIL.n521 185
R156 VTAIL.n582 VTAIL.n581 185
R157 VTAIL.n580 VTAIL.n579 185
R158 VTAIL.n527 VTAIL.n526 185
R159 VTAIL.n574 VTAIL.n573 185
R160 VTAIL.n572 VTAIL.n571 185
R161 VTAIL.n531 VTAIL.n530 185
R162 VTAIL.n566 VTAIL.n565 185
R163 VTAIL.n564 VTAIL.n563 185
R164 VTAIL.n535 VTAIL.n534 185
R165 VTAIL.n558 VTAIL.n557 185
R166 VTAIL.n556 VTAIL.n555 185
R167 VTAIL.n539 VTAIL.n538 185
R168 VTAIL.n550 VTAIL.n549 185
R169 VTAIL.n548 VTAIL.n547 185
R170 VTAIL.n543 VTAIL.n542 185
R171 VTAIL.n505 VTAIL.n504 185
R172 VTAIL.n503 VTAIL.n502 185
R173 VTAIL.n412 VTAIL.n411 185
R174 VTAIL.n497 VTAIL.n496 185
R175 VTAIL.n495 VTAIL.n494 185
R176 VTAIL.n416 VTAIL.n415 185
R177 VTAIL.n489 VTAIL.n488 185
R178 VTAIL.n487 VTAIL.n418 185
R179 VTAIL.n486 VTAIL.n485 185
R180 VTAIL.n421 VTAIL.n419 185
R181 VTAIL.n480 VTAIL.n479 185
R182 VTAIL.n478 VTAIL.n477 185
R183 VTAIL.n425 VTAIL.n424 185
R184 VTAIL.n472 VTAIL.n471 185
R185 VTAIL.n470 VTAIL.n469 185
R186 VTAIL.n429 VTAIL.n428 185
R187 VTAIL.n464 VTAIL.n463 185
R188 VTAIL.n462 VTAIL.n461 185
R189 VTAIL.n433 VTAIL.n432 185
R190 VTAIL.n456 VTAIL.n455 185
R191 VTAIL.n454 VTAIL.n453 185
R192 VTAIL.n437 VTAIL.n436 185
R193 VTAIL.n448 VTAIL.n447 185
R194 VTAIL.n446 VTAIL.n445 185
R195 VTAIL.n441 VTAIL.n440 185
R196 VTAIL.n403 VTAIL.n402 185
R197 VTAIL.n401 VTAIL.n400 185
R198 VTAIL.n310 VTAIL.n309 185
R199 VTAIL.n395 VTAIL.n394 185
R200 VTAIL.n393 VTAIL.n392 185
R201 VTAIL.n314 VTAIL.n313 185
R202 VTAIL.n387 VTAIL.n386 185
R203 VTAIL.n385 VTAIL.n316 185
R204 VTAIL.n384 VTAIL.n383 185
R205 VTAIL.n319 VTAIL.n317 185
R206 VTAIL.n378 VTAIL.n377 185
R207 VTAIL.n376 VTAIL.n375 185
R208 VTAIL.n323 VTAIL.n322 185
R209 VTAIL.n370 VTAIL.n369 185
R210 VTAIL.n368 VTAIL.n367 185
R211 VTAIL.n327 VTAIL.n326 185
R212 VTAIL.n362 VTAIL.n361 185
R213 VTAIL.n360 VTAIL.n359 185
R214 VTAIL.n331 VTAIL.n330 185
R215 VTAIL.n354 VTAIL.n353 185
R216 VTAIL.n352 VTAIL.n351 185
R217 VTAIL.n335 VTAIL.n334 185
R218 VTAIL.n346 VTAIL.n345 185
R219 VTAIL.n344 VTAIL.n343 185
R220 VTAIL.n339 VTAIL.n338 185
R221 VTAIL.n747 VTAIL.t6 147.659
R222 VTAIL.n33 VTAIL.t7 147.659
R223 VTAIL.n135 VTAIL.t1 147.659
R224 VTAIL.n237 VTAIL.t2 147.659
R225 VTAIL.n646 VTAIL.t3 147.659
R226 VTAIL.n544 VTAIL.t0 147.659
R227 VTAIL.n442 VTAIL.t5 147.659
R228 VTAIL.n340 VTAIL.t4 147.659
R229 VTAIL.n751 VTAIL.n745 104.615
R230 VTAIL.n752 VTAIL.n751 104.615
R231 VTAIL.n752 VTAIL.n741 104.615
R232 VTAIL.n759 VTAIL.n741 104.615
R233 VTAIL.n760 VTAIL.n759 104.615
R234 VTAIL.n760 VTAIL.n737 104.615
R235 VTAIL.n767 VTAIL.n737 104.615
R236 VTAIL.n768 VTAIL.n767 104.615
R237 VTAIL.n768 VTAIL.n733 104.615
R238 VTAIL.n775 VTAIL.n733 104.615
R239 VTAIL.n776 VTAIL.n775 104.615
R240 VTAIL.n776 VTAIL.n729 104.615
R241 VTAIL.n783 VTAIL.n729 104.615
R242 VTAIL.n784 VTAIL.n783 104.615
R243 VTAIL.n784 VTAIL.n725 104.615
R244 VTAIL.n792 VTAIL.n725 104.615
R245 VTAIL.n793 VTAIL.n792 104.615
R246 VTAIL.n794 VTAIL.n793 104.615
R247 VTAIL.n794 VTAIL.n721 104.615
R248 VTAIL.n801 VTAIL.n721 104.615
R249 VTAIL.n802 VTAIL.n801 104.615
R250 VTAIL.n802 VTAIL.n717 104.615
R251 VTAIL.n809 VTAIL.n717 104.615
R252 VTAIL.n810 VTAIL.n809 104.615
R253 VTAIL.n37 VTAIL.n31 104.615
R254 VTAIL.n38 VTAIL.n37 104.615
R255 VTAIL.n38 VTAIL.n27 104.615
R256 VTAIL.n45 VTAIL.n27 104.615
R257 VTAIL.n46 VTAIL.n45 104.615
R258 VTAIL.n46 VTAIL.n23 104.615
R259 VTAIL.n53 VTAIL.n23 104.615
R260 VTAIL.n54 VTAIL.n53 104.615
R261 VTAIL.n54 VTAIL.n19 104.615
R262 VTAIL.n61 VTAIL.n19 104.615
R263 VTAIL.n62 VTAIL.n61 104.615
R264 VTAIL.n62 VTAIL.n15 104.615
R265 VTAIL.n69 VTAIL.n15 104.615
R266 VTAIL.n70 VTAIL.n69 104.615
R267 VTAIL.n70 VTAIL.n11 104.615
R268 VTAIL.n78 VTAIL.n11 104.615
R269 VTAIL.n79 VTAIL.n78 104.615
R270 VTAIL.n80 VTAIL.n79 104.615
R271 VTAIL.n80 VTAIL.n7 104.615
R272 VTAIL.n87 VTAIL.n7 104.615
R273 VTAIL.n88 VTAIL.n87 104.615
R274 VTAIL.n88 VTAIL.n3 104.615
R275 VTAIL.n95 VTAIL.n3 104.615
R276 VTAIL.n96 VTAIL.n95 104.615
R277 VTAIL.n139 VTAIL.n133 104.615
R278 VTAIL.n140 VTAIL.n139 104.615
R279 VTAIL.n140 VTAIL.n129 104.615
R280 VTAIL.n147 VTAIL.n129 104.615
R281 VTAIL.n148 VTAIL.n147 104.615
R282 VTAIL.n148 VTAIL.n125 104.615
R283 VTAIL.n155 VTAIL.n125 104.615
R284 VTAIL.n156 VTAIL.n155 104.615
R285 VTAIL.n156 VTAIL.n121 104.615
R286 VTAIL.n163 VTAIL.n121 104.615
R287 VTAIL.n164 VTAIL.n163 104.615
R288 VTAIL.n164 VTAIL.n117 104.615
R289 VTAIL.n171 VTAIL.n117 104.615
R290 VTAIL.n172 VTAIL.n171 104.615
R291 VTAIL.n172 VTAIL.n113 104.615
R292 VTAIL.n180 VTAIL.n113 104.615
R293 VTAIL.n181 VTAIL.n180 104.615
R294 VTAIL.n182 VTAIL.n181 104.615
R295 VTAIL.n182 VTAIL.n109 104.615
R296 VTAIL.n189 VTAIL.n109 104.615
R297 VTAIL.n190 VTAIL.n189 104.615
R298 VTAIL.n190 VTAIL.n105 104.615
R299 VTAIL.n197 VTAIL.n105 104.615
R300 VTAIL.n198 VTAIL.n197 104.615
R301 VTAIL.n241 VTAIL.n235 104.615
R302 VTAIL.n242 VTAIL.n241 104.615
R303 VTAIL.n242 VTAIL.n231 104.615
R304 VTAIL.n249 VTAIL.n231 104.615
R305 VTAIL.n250 VTAIL.n249 104.615
R306 VTAIL.n250 VTAIL.n227 104.615
R307 VTAIL.n257 VTAIL.n227 104.615
R308 VTAIL.n258 VTAIL.n257 104.615
R309 VTAIL.n258 VTAIL.n223 104.615
R310 VTAIL.n265 VTAIL.n223 104.615
R311 VTAIL.n266 VTAIL.n265 104.615
R312 VTAIL.n266 VTAIL.n219 104.615
R313 VTAIL.n273 VTAIL.n219 104.615
R314 VTAIL.n274 VTAIL.n273 104.615
R315 VTAIL.n274 VTAIL.n215 104.615
R316 VTAIL.n282 VTAIL.n215 104.615
R317 VTAIL.n283 VTAIL.n282 104.615
R318 VTAIL.n284 VTAIL.n283 104.615
R319 VTAIL.n284 VTAIL.n211 104.615
R320 VTAIL.n291 VTAIL.n211 104.615
R321 VTAIL.n292 VTAIL.n291 104.615
R322 VTAIL.n292 VTAIL.n207 104.615
R323 VTAIL.n299 VTAIL.n207 104.615
R324 VTAIL.n300 VTAIL.n299 104.615
R325 VTAIL.n708 VTAIL.n707 104.615
R326 VTAIL.n707 VTAIL.n615 104.615
R327 VTAIL.n700 VTAIL.n615 104.615
R328 VTAIL.n700 VTAIL.n699 104.615
R329 VTAIL.n699 VTAIL.n619 104.615
R330 VTAIL.n692 VTAIL.n619 104.615
R331 VTAIL.n692 VTAIL.n691 104.615
R332 VTAIL.n691 VTAIL.n690 104.615
R333 VTAIL.n690 VTAIL.n623 104.615
R334 VTAIL.n683 VTAIL.n623 104.615
R335 VTAIL.n683 VTAIL.n682 104.615
R336 VTAIL.n682 VTAIL.n628 104.615
R337 VTAIL.n675 VTAIL.n628 104.615
R338 VTAIL.n675 VTAIL.n674 104.615
R339 VTAIL.n674 VTAIL.n632 104.615
R340 VTAIL.n667 VTAIL.n632 104.615
R341 VTAIL.n667 VTAIL.n666 104.615
R342 VTAIL.n666 VTAIL.n636 104.615
R343 VTAIL.n659 VTAIL.n636 104.615
R344 VTAIL.n659 VTAIL.n658 104.615
R345 VTAIL.n658 VTAIL.n640 104.615
R346 VTAIL.n651 VTAIL.n640 104.615
R347 VTAIL.n651 VTAIL.n650 104.615
R348 VTAIL.n650 VTAIL.n644 104.615
R349 VTAIL.n606 VTAIL.n605 104.615
R350 VTAIL.n605 VTAIL.n513 104.615
R351 VTAIL.n598 VTAIL.n513 104.615
R352 VTAIL.n598 VTAIL.n597 104.615
R353 VTAIL.n597 VTAIL.n517 104.615
R354 VTAIL.n590 VTAIL.n517 104.615
R355 VTAIL.n590 VTAIL.n589 104.615
R356 VTAIL.n589 VTAIL.n588 104.615
R357 VTAIL.n588 VTAIL.n521 104.615
R358 VTAIL.n581 VTAIL.n521 104.615
R359 VTAIL.n581 VTAIL.n580 104.615
R360 VTAIL.n580 VTAIL.n526 104.615
R361 VTAIL.n573 VTAIL.n526 104.615
R362 VTAIL.n573 VTAIL.n572 104.615
R363 VTAIL.n572 VTAIL.n530 104.615
R364 VTAIL.n565 VTAIL.n530 104.615
R365 VTAIL.n565 VTAIL.n564 104.615
R366 VTAIL.n564 VTAIL.n534 104.615
R367 VTAIL.n557 VTAIL.n534 104.615
R368 VTAIL.n557 VTAIL.n556 104.615
R369 VTAIL.n556 VTAIL.n538 104.615
R370 VTAIL.n549 VTAIL.n538 104.615
R371 VTAIL.n549 VTAIL.n548 104.615
R372 VTAIL.n548 VTAIL.n542 104.615
R373 VTAIL.n504 VTAIL.n503 104.615
R374 VTAIL.n503 VTAIL.n411 104.615
R375 VTAIL.n496 VTAIL.n411 104.615
R376 VTAIL.n496 VTAIL.n495 104.615
R377 VTAIL.n495 VTAIL.n415 104.615
R378 VTAIL.n488 VTAIL.n415 104.615
R379 VTAIL.n488 VTAIL.n487 104.615
R380 VTAIL.n487 VTAIL.n486 104.615
R381 VTAIL.n486 VTAIL.n419 104.615
R382 VTAIL.n479 VTAIL.n419 104.615
R383 VTAIL.n479 VTAIL.n478 104.615
R384 VTAIL.n478 VTAIL.n424 104.615
R385 VTAIL.n471 VTAIL.n424 104.615
R386 VTAIL.n471 VTAIL.n470 104.615
R387 VTAIL.n470 VTAIL.n428 104.615
R388 VTAIL.n463 VTAIL.n428 104.615
R389 VTAIL.n463 VTAIL.n462 104.615
R390 VTAIL.n462 VTAIL.n432 104.615
R391 VTAIL.n455 VTAIL.n432 104.615
R392 VTAIL.n455 VTAIL.n454 104.615
R393 VTAIL.n454 VTAIL.n436 104.615
R394 VTAIL.n447 VTAIL.n436 104.615
R395 VTAIL.n447 VTAIL.n446 104.615
R396 VTAIL.n446 VTAIL.n440 104.615
R397 VTAIL.n402 VTAIL.n401 104.615
R398 VTAIL.n401 VTAIL.n309 104.615
R399 VTAIL.n394 VTAIL.n309 104.615
R400 VTAIL.n394 VTAIL.n393 104.615
R401 VTAIL.n393 VTAIL.n313 104.615
R402 VTAIL.n386 VTAIL.n313 104.615
R403 VTAIL.n386 VTAIL.n385 104.615
R404 VTAIL.n385 VTAIL.n384 104.615
R405 VTAIL.n384 VTAIL.n317 104.615
R406 VTAIL.n377 VTAIL.n317 104.615
R407 VTAIL.n377 VTAIL.n376 104.615
R408 VTAIL.n376 VTAIL.n322 104.615
R409 VTAIL.n369 VTAIL.n322 104.615
R410 VTAIL.n369 VTAIL.n368 104.615
R411 VTAIL.n368 VTAIL.n326 104.615
R412 VTAIL.n361 VTAIL.n326 104.615
R413 VTAIL.n361 VTAIL.n360 104.615
R414 VTAIL.n360 VTAIL.n330 104.615
R415 VTAIL.n353 VTAIL.n330 104.615
R416 VTAIL.n353 VTAIL.n352 104.615
R417 VTAIL.n352 VTAIL.n334 104.615
R418 VTAIL.n345 VTAIL.n334 104.615
R419 VTAIL.n345 VTAIL.n344 104.615
R420 VTAIL.n344 VTAIL.n338 104.615
R421 VTAIL.t6 VTAIL.n745 52.3082
R422 VTAIL.t7 VTAIL.n31 52.3082
R423 VTAIL.t1 VTAIL.n133 52.3082
R424 VTAIL.t2 VTAIL.n235 52.3082
R425 VTAIL.t3 VTAIL.n644 52.3082
R426 VTAIL.t0 VTAIL.n542 52.3082
R427 VTAIL.t5 VTAIL.n440 52.3082
R428 VTAIL.t4 VTAIL.n338 52.3082
R429 VTAIL.n815 VTAIL.n814 33.7369
R430 VTAIL.n101 VTAIL.n100 33.7369
R431 VTAIL.n203 VTAIL.n202 33.7369
R432 VTAIL.n305 VTAIL.n304 33.7369
R433 VTAIL.n713 VTAIL.n712 33.7369
R434 VTAIL.n611 VTAIL.n610 33.7369
R435 VTAIL.n509 VTAIL.n508 33.7369
R436 VTAIL.n407 VTAIL.n406 33.7369
R437 VTAIL.n815 VTAIL.n713 31.8583
R438 VTAIL.n407 VTAIL.n305 31.8583
R439 VTAIL.n747 VTAIL.n746 15.6677
R440 VTAIL.n33 VTAIL.n32 15.6677
R441 VTAIL.n135 VTAIL.n134 15.6677
R442 VTAIL.n237 VTAIL.n236 15.6677
R443 VTAIL.n646 VTAIL.n645 15.6677
R444 VTAIL.n544 VTAIL.n543 15.6677
R445 VTAIL.n442 VTAIL.n441 15.6677
R446 VTAIL.n340 VTAIL.n339 15.6677
R447 VTAIL.n795 VTAIL.n724 13.1884
R448 VTAIL.n81 VTAIL.n10 13.1884
R449 VTAIL.n183 VTAIL.n112 13.1884
R450 VTAIL.n285 VTAIL.n214 13.1884
R451 VTAIL.n693 VTAIL.n622 13.1884
R452 VTAIL.n591 VTAIL.n520 13.1884
R453 VTAIL.n489 VTAIL.n418 13.1884
R454 VTAIL.n387 VTAIL.n316 13.1884
R455 VTAIL.n750 VTAIL.n749 12.8005
R456 VTAIL.n791 VTAIL.n790 12.8005
R457 VTAIL.n796 VTAIL.n722 12.8005
R458 VTAIL.n36 VTAIL.n35 12.8005
R459 VTAIL.n77 VTAIL.n76 12.8005
R460 VTAIL.n82 VTAIL.n8 12.8005
R461 VTAIL.n138 VTAIL.n137 12.8005
R462 VTAIL.n179 VTAIL.n178 12.8005
R463 VTAIL.n184 VTAIL.n110 12.8005
R464 VTAIL.n240 VTAIL.n239 12.8005
R465 VTAIL.n281 VTAIL.n280 12.8005
R466 VTAIL.n286 VTAIL.n212 12.8005
R467 VTAIL.n694 VTAIL.n620 12.8005
R468 VTAIL.n689 VTAIL.n624 12.8005
R469 VTAIL.n649 VTAIL.n648 12.8005
R470 VTAIL.n592 VTAIL.n518 12.8005
R471 VTAIL.n587 VTAIL.n522 12.8005
R472 VTAIL.n547 VTAIL.n546 12.8005
R473 VTAIL.n490 VTAIL.n416 12.8005
R474 VTAIL.n485 VTAIL.n420 12.8005
R475 VTAIL.n445 VTAIL.n444 12.8005
R476 VTAIL.n388 VTAIL.n314 12.8005
R477 VTAIL.n383 VTAIL.n318 12.8005
R478 VTAIL.n343 VTAIL.n342 12.8005
R479 VTAIL.n753 VTAIL.n744 12.0247
R480 VTAIL.n789 VTAIL.n726 12.0247
R481 VTAIL.n800 VTAIL.n799 12.0247
R482 VTAIL.n39 VTAIL.n30 12.0247
R483 VTAIL.n75 VTAIL.n12 12.0247
R484 VTAIL.n86 VTAIL.n85 12.0247
R485 VTAIL.n141 VTAIL.n132 12.0247
R486 VTAIL.n177 VTAIL.n114 12.0247
R487 VTAIL.n188 VTAIL.n187 12.0247
R488 VTAIL.n243 VTAIL.n234 12.0247
R489 VTAIL.n279 VTAIL.n216 12.0247
R490 VTAIL.n290 VTAIL.n289 12.0247
R491 VTAIL.n698 VTAIL.n697 12.0247
R492 VTAIL.n688 VTAIL.n625 12.0247
R493 VTAIL.n652 VTAIL.n643 12.0247
R494 VTAIL.n596 VTAIL.n595 12.0247
R495 VTAIL.n586 VTAIL.n523 12.0247
R496 VTAIL.n550 VTAIL.n541 12.0247
R497 VTAIL.n494 VTAIL.n493 12.0247
R498 VTAIL.n484 VTAIL.n421 12.0247
R499 VTAIL.n448 VTAIL.n439 12.0247
R500 VTAIL.n392 VTAIL.n391 12.0247
R501 VTAIL.n382 VTAIL.n319 12.0247
R502 VTAIL.n346 VTAIL.n337 12.0247
R503 VTAIL.n754 VTAIL.n742 11.249
R504 VTAIL.n786 VTAIL.n785 11.249
R505 VTAIL.n803 VTAIL.n720 11.249
R506 VTAIL.n40 VTAIL.n28 11.249
R507 VTAIL.n72 VTAIL.n71 11.249
R508 VTAIL.n89 VTAIL.n6 11.249
R509 VTAIL.n142 VTAIL.n130 11.249
R510 VTAIL.n174 VTAIL.n173 11.249
R511 VTAIL.n191 VTAIL.n108 11.249
R512 VTAIL.n244 VTAIL.n232 11.249
R513 VTAIL.n276 VTAIL.n275 11.249
R514 VTAIL.n293 VTAIL.n210 11.249
R515 VTAIL.n701 VTAIL.n618 11.249
R516 VTAIL.n685 VTAIL.n684 11.249
R517 VTAIL.n653 VTAIL.n641 11.249
R518 VTAIL.n599 VTAIL.n516 11.249
R519 VTAIL.n583 VTAIL.n582 11.249
R520 VTAIL.n551 VTAIL.n539 11.249
R521 VTAIL.n497 VTAIL.n414 11.249
R522 VTAIL.n481 VTAIL.n480 11.249
R523 VTAIL.n449 VTAIL.n437 11.249
R524 VTAIL.n395 VTAIL.n312 11.249
R525 VTAIL.n379 VTAIL.n378 11.249
R526 VTAIL.n347 VTAIL.n335 11.249
R527 VTAIL.n758 VTAIL.n757 10.4732
R528 VTAIL.n782 VTAIL.n728 10.4732
R529 VTAIL.n804 VTAIL.n718 10.4732
R530 VTAIL.n44 VTAIL.n43 10.4732
R531 VTAIL.n68 VTAIL.n14 10.4732
R532 VTAIL.n90 VTAIL.n4 10.4732
R533 VTAIL.n146 VTAIL.n145 10.4732
R534 VTAIL.n170 VTAIL.n116 10.4732
R535 VTAIL.n192 VTAIL.n106 10.4732
R536 VTAIL.n248 VTAIL.n247 10.4732
R537 VTAIL.n272 VTAIL.n218 10.4732
R538 VTAIL.n294 VTAIL.n208 10.4732
R539 VTAIL.n702 VTAIL.n616 10.4732
R540 VTAIL.n681 VTAIL.n627 10.4732
R541 VTAIL.n657 VTAIL.n656 10.4732
R542 VTAIL.n600 VTAIL.n514 10.4732
R543 VTAIL.n579 VTAIL.n525 10.4732
R544 VTAIL.n555 VTAIL.n554 10.4732
R545 VTAIL.n498 VTAIL.n412 10.4732
R546 VTAIL.n477 VTAIL.n423 10.4732
R547 VTAIL.n453 VTAIL.n452 10.4732
R548 VTAIL.n396 VTAIL.n310 10.4732
R549 VTAIL.n375 VTAIL.n321 10.4732
R550 VTAIL.n351 VTAIL.n350 10.4732
R551 VTAIL.n761 VTAIL.n740 9.69747
R552 VTAIL.n781 VTAIL.n730 9.69747
R553 VTAIL.n808 VTAIL.n807 9.69747
R554 VTAIL.n47 VTAIL.n26 9.69747
R555 VTAIL.n67 VTAIL.n16 9.69747
R556 VTAIL.n94 VTAIL.n93 9.69747
R557 VTAIL.n149 VTAIL.n128 9.69747
R558 VTAIL.n169 VTAIL.n118 9.69747
R559 VTAIL.n196 VTAIL.n195 9.69747
R560 VTAIL.n251 VTAIL.n230 9.69747
R561 VTAIL.n271 VTAIL.n220 9.69747
R562 VTAIL.n298 VTAIL.n297 9.69747
R563 VTAIL.n706 VTAIL.n705 9.69747
R564 VTAIL.n680 VTAIL.n629 9.69747
R565 VTAIL.n660 VTAIL.n639 9.69747
R566 VTAIL.n604 VTAIL.n603 9.69747
R567 VTAIL.n578 VTAIL.n527 9.69747
R568 VTAIL.n558 VTAIL.n537 9.69747
R569 VTAIL.n502 VTAIL.n501 9.69747
R570 VTAIL.n476 VTAIL.n425 9.69747
R571 VTAIL.n456 VTAIL.n435 9.69747
R572 VTAIL.n400 VTAIL.n399 9.69747
R573 VTAIL.n374 VTAIL.n323 9.69747
R574 VTAIL.n354 VTAIL.n333 9.69747
R575 VTAIL.n814 VTAIL.n813 9.45567
R576 VTAIL.n100 VTAIL.n99 9.45567
R577 VTAIL.n202 VTAIL.n201 9.45567
R578 VTAIL.n304 VTAIL.n303 9.45567
R579 VTAIL.n712 VTAIL.n711 9.45567
R580 VTAIL.n610 VTAIL.n609 9.45567
R581 VTAIL.n508 VTAIL.n507 9.45567
R582 VTAIL.n406 VTAIL.n405 9.45567
R583 VTAIL.n813 VTAIL.n812 9.3005
R584 VTAIL.n716 VTAIL.n715 9.3005
R585 VTAIL.n807 VTAIL.n806 9.3005
R586 VTAIL.n805 VTAIL.n804 9.3005
R587 VTAIL.n720 VTAIL.n719 9.3005
R588 VTAIL.n799 VTAIL.n798 9.3005
R589 VTAIL.n797 VTAIL.n796 9.3005
R590 VTAIL.n736 VTAIL.n735 9.3005
R591 VTAIL.n765 VTAIL.n764 9.3005
R592 VTAIL.n763 VTAIL.n762 9.3005
R593 VTAIL.n740 VTAIL.n739 9.3005
R594 VTAIL.n757 VTAIL.n756 9.3005
R595 VTAIL.n755 VTAIL.n754 9.3005
R596 VTAIL.n744 VTAIL.n743 9.3005
R597 VTAIL.n749 VTAIL.n748 9.3005
R598 VTAIL.n771 VTAIL.n770 9.3005
R599 VTAIL.n773 VTAIL.n772 9.3005
R600 VTAIL.n732 VTAIL.n731 9.3005
R601 VTAIL.n779 VTAIL.n778 9.3005
R602 VTAIL.n781 VTAIL.n780 9.3005
R603 VTAIL.n728 VTAIL.n727 9.3005
R604 VTAIL.n787 VTAIL.n786 9.3005
R605 VTAIL.n789 VTAIL.n788 9.3005
R606 VTAIL.n790 VTAIL.n723 9.3005
R607 VTAIL.n99 VTAIL.n98 9.3005
R608 VTAIL.n2 VTAIL.n1 9.3005
R609 VTAIL.n93 VTAIL.n92 9.3005
R610 VTAIL.n91 VTAIL.n90 9.3005
R611 VTAIL.n6 VTAIL.n5 9.3005
R612 VTAIL.n85 VTAIL.n84 9.3005
R613 VTAIL.n83 VTAIL.n82 9.3005
R614 VTAIL.n22 VTAIL.n21 9.3005
R615 VTAIL.n51 VTAIL.n50 9.3005
R616 VTAIL.n49 VTAIL.n48 9.3005
R617 VTAIL.n26 VTAIL.n25 9.3005
R618 VTAIL.n43 VTAIL.n42 9.3005
R619 VTAIL.n41 VTAIL.n40 9.3005
R620 VTAIL.n30 VTAIL.n29 9.3005
R621 VTAIL.n35 VTAIL.n34 9.3005
R622 VTAIL.n57 VTAIL.n56 9.3005
R623 VTAIL.n59 VTAIL.n58 9.3005
R624 VTAIL.n18 VTAIL.n17 9.3005
R625 VTAIL.n65 VTAIL.n64 9.3005
R626 VTAIL.n67 VTAIL.n66 9.3005
R627 VTAIL.n14 VTAIL.n13 9.3005
R628 VTAIL.n73 VTAIL.n72 9.3005
R629 VTAIL.n75 VTAIL.n74 9.3005
R630 VTAIL.n76 VTAIL.n9 9.3005
R631 VTAIL.n201 VTAIL.n200 9.3005
R632 VTAIL.n104 VTAIL.n103 9.3005
R633 VTAIL.n195 VTAIL.n194 9.3005
R634 VTAIL.n193 VTAIL.n192 9.3005
R635 VTAIL.n108 VTAIL.n107 9.3005
R636 VTAIL.n187 VTAIL.n186 9.3005
R637 VTAIL.n185 VTAIL.n184 9.3005
R638 VTAIL.n124 VTAIL.n123 9.3005
R639 VTAIL.n153 VTAIL.n152 9.3005
R640 VTAIL.n151 VTAIL.n150 9.3005
R641 VTAIL.n128 VTAIL.n127 9.3005
R642 VTAIL.n145 VTAIL.n144 9.3005
R643 VTAIL.n143 VTAIL.n142 9.3005
R644 VTAIL.n132 VTAIL.n131 9.3005
R645 VTAIL.n137 VTAIL.n136 9.3005
R646 VTAIL.n159 VTAIL.n158 9.3005
R647 VTAIL.n161 VTAIL.n160 9.3005
R648 VTAIL.n120 VTAIL.n119 9.3005
R649 VTAIL.n167 VTAIL.n166 9.3005
R650 VTAIL.n169 VTAIL.n168 9.3005
R651 VTAIL.n116 VTAIL.n115 9.3005
R652 VTAIL.n175 VTAIL.n174 9.3005
R653 VTAIL.n177 VTAIL.n176 9.3005
R654 VTAIL.n178 VTAIL.n111 9.3005
R655 VTAIL.n303 VTAIL.n302 9.3005
R656 VTAIL.n206 VTAIL.n205 9.3005
R657 VTAIL.n297 VTAIL.n296 9.3005
R658 VTAIL.n295 VTAIL.n294 9.3005
R659 VTAIL.n210 VTAIL.n209 9.3005
R660 VTAIL.n289 VTAIL.n288 9.3005
R661 VTAIL.n287 VTAIL.n286 9.3005
R662 VTAIL.n226 VTAIL.n225 9.3005
R663 VTAIL.n255 VTAIL.n254 9.3005
R664 VTAIL.n253 VTAIL.n252 9.3005
R665 VTAIL.n230 VTAIL.n229 9.3005
R666 VTAIL.n247 VTAIL.n246 9.3005
R667 VTAIL.n245 VTAIL.n244 9.3005
R668 VTAIL.n234 VTAIL.n233 9.3005
R669 VTAIL.n239 VTAIL.n238 9.3005
R670 VTAIL.n261 VTAIL.n260 9.3005
R671 VTAIL.n263 VTAIL.n262 9.3005
R672 VTAIL.n222 VTAIL.n221 9.3005
R673 VTAIL.n269 VTAIL.n268 9.3005
R674 VTAIL.n271 VTAIL.n270 9.3005
R675 VTAIL.n218 VTAIL.n217 9.3005
R676 VTAIL.n277 VTAIL.n276 9.3005
R677 VTAIL.n279 VTAIL.n278 9.3005
R678 VTAIL.n280 VTAIL.n213 9.3005
R679 VTAIL.n672 VTAIL.n671 9.3005
R680 VTAIL.n631 VTAIL.n630 9.3005
R681 VTAIL.n678 VTAIL.n677 9.3005
R682 VTAIL.n680 VTAIL.n679 9.3005
R683 VTAIL.n627 VTAIL.n626 9.3005
R684 VTAIL.n686 VTAIL.n685 9.3005
R685 VTAIL.n688 VTAIL.n687 9.3005
R686 VTAIL.n624 VTAIL.n621 9.3005
R687 VTAIL.n711 VTAIL.n710 9.3005
R688 VTAIL.n614 VTAIL.n613 9.3005
R689 VTAIL.n705 VTAIL.n704 9.3005
R690 VTAIL.n703 VTAIL.n702 9.3005
R691 VTAIL.n618 VTAIL.n617 9.3005
R692 VTAIL.n697 VTAIL.n696 9.3005
R693 VTAIL.n695 VTAIL.n694 9.3005
R694 VTAIL.n670 VTAIL.n669 9.3005
R695 VTAIL.n635 VTAIL.n634 9.3005
R696 VTAIL.n664 VTAIL.n663 9.3005
R697 VTAIL.n662 VTAIL.n661 9.3005
R698 VTAIL.n639 VTAIL.n638 9.3005
R699 VTAIL.n656 VTAIL.n655 9.3005
R700 VTAIL.n654 VTAIL.n653 9.3005
R701 VTAIL.n643 VTAIL.n642 9.3005
R702 VTAIL.n648 VTAIL.n647 9.3005
R703 VTAIL.n570 VTAIL.n569 9.3005
R704 VTAIL.n529 VTAIL.n528 9.3005
R705 VTAIL.n576 VTAIL.n575 9.3005
R706 VTAIL.n578 VTAIL.n577 9.3005
R707 VTAIL.n525 VTAIL.n524 9.3005
R708 VTAIL.n584 VTAIL.n583 9.3005
R709 VTAIL.n586 VTAIL.n585 9.3005
R710 VTAIL.n522 VTAIL.n519 9.3005
R711 VTAIL.n609 VTAIL.n608 9.3005
R712 VTAIL.n512 VTAIL.n511 9.3005
R713 VTAIL.n603 VTAIL.n602 9.3005
R714 VTAIL.n601 VTAIL.n600 9.3005
R715 VTAIL.n516 VTAIL.n515 9.3005
R716 VTAIL.n595 VTAIL.n594 9.3005
R717 VTAIL.n593 VTAIL.n592 9.3005
R718 VTAIL.n568 VTAIL.n567 9.3005
R719 VTAIL.n533 VTAIL.n532 9.3005
R720 VTAIL.n562 VTAIL.n561 9.3005
R721 VTAIL.n560 VTAIL.n559 9.3005
R722 VTAIL.n537 VTAIL.n536 9.3005
R723 VTAIL.n554 VTAIL.n553 9.3005
R724 VTAIL.n552 VTAIL.n551 9.3005
R725 VTAIL.n541 VTAIL.n540 9.3005
R726 VTAIL.n546 VTAIL.n545 9.3005
R727 VTAIL.n468 VTAIL.n467 9.3005
R728 VTAIL.n427 VTAIL.n426 9.3005
R729 VTAIL.n474 VTAIL.n473 9.3005
R730 VTAIL.n476 VTAIL.n475 9.3005
R731 VTAIL.n423 VTAIL.n422 9.3005
R732 VTAIL.n482 VTAIL.n481 9.3005
R733 VTAIL.n484 VTAIL.n483 9.3005
R734 VTAIL.n420 VTAIL.n417 9.3005
R735 VTAIL.n507 VTAIL.n506 9.3005
R736 VTAIL.n410 VTAIL.n409 9.3005
R737 VTAIL.n501 VTAIL.n500 9.3005
R738 VTAIL.n499 VTAIL.n498 9.3005
R739 VTAIL.n414 VTAIL.n413 9.3005
R740 VTAIL.n493 VTAIL.n492 9.3005
R741 VTAIL.n491 VTAIL.n490 9.3005
R742 VTAIL.n466 VTAIL.n465 9.3005
R743 VTAIL.n431 VTAIL.n430 9.3005
R744 VTAIL.n460 VTAIL.n459 9.3005
R745 VTAIL.n458 VTAIL.n457 9.3005
R746 VTAIL.n435 VTAIL.n434 9.3005
R747 VTAIL.n452 VTAIL.n451 9.3005
R748 VTAIL.n450 VTAIL.n449 9.3005
R749 VTAIL.n439 VTAIL.n438 9.3005
R750 VTAIL.n444 VTAIL.n443 9.3005
R751 VTAIL.n366 VTAIL.n365 9.3005
R752 VTAIL.n325 VTAIL.n324 9.3005
R753 VTAIL.n372 VTAIL.n371 9.3005
R754 VTAIL.n374 VTAIL.n373 9.3005
R755 VTAIL.n321 VTAIL.n320 9.3005
R756 VTAIL.n380 VTAIL.n379 9.3005
R757 VTAIL.n382 VTAIL.n381 9.3005
R758 VTAIL.n318 VTAIL.n315 9.3005
R759 VTAIL.n405 VTAIL.n404 9.3005
R760 VTAIL.n308 VTAIL.n307 9.3005
R761 VTAIL.n399 VTAIL.n398 9.3005
R762 VTAIL.n397 VTAIL.n396 9.3005
R763 VTAIL.n312 VTAIL.n311 9.3005
R764 VTAIL.n391 VTAIL.n390 9.3005
R765 VTAIL.n389 VTAIL.n388 9.3005
R766 VTAIL.n364 VTAIL.n363 9.3005
R767 VTAIL.n329 VTAIL.n328 9.3005
R768 VTAIL.n358 VTAIL.n357 9.3005
R769 VTAIL.n356 VTAIL.n355 9.3005
R770 VTAIL.n333 VTAIL.n332 9.3005
R771 VTAIL.n350 VTAIL.n349 9.3005
R772 VTAIL.n348 VTAIL.n347 9.3005
R773 VTAIL.n337 VTAIL.n336 9.3005
R774 VTAIL.n342 VTAIL.n341 9.3005
R775 VTAIL.n762 VTAIL.n738 8.92171
R776 VTAIL.n778 VTAIL.n777 8.92171
R777 VTAIL.n811 VTAIL.n716 8.92171
R778 VTAIL.n48 VTAIL.n24 8.92171
R779 VTAIL.n64 VTAIL.n63 8.92171
R780 VTAIL.n97 VTAIL.n2 8.92171
R781 VTAIL.n150 VTAIL.n126 8.92171
R782 VTAIL.n166 VTAIL.n165 8.92171
R783 VTAIL.n199 VTAIL.n104 8.92171
R784 VTAIL.n252 VTAIL.n228 8.92171
R785 VTAIL.n268 VTAIL.n267 8.92171
R786 VTAIL.n301 VTAIL.n206 8.92171
R787 VTAIL.n709 VTAIL.n614 8.92171
R788 VTAIL.n677 VTAIL.n676 8.92171
R789 VTAIL.n661 VTAIL.n637 8.92171
R790 VTAIL.n607 VTAIL.n512 8.92171
R791 VTAIL.n575 VTAIL.n574 8.92171
R792 VTAIL.n559 VTAIL.n535 8.92171
R793 VTAIL.n505 VTAIL.n410 8.92171
R794 VTAIL.n473 VTAIL.n472 8.92171
R795 VTAIL.n457 VTAIL.n433 8.92171
R796 VTAIL.n403 VTAIL.n308 8.92171
R797 VTAIL.n371 VTAIL.n370 8.92171
R798 VTAIL.n355 VTAIL.n331 8.92171
R799 VTAIL.n766 VTAIL.n765 8.14595
R800 VTAIL.n774 VTAIL.n732 8.14595
R801 VTAIL.n812 VTAIL.n714 8.14595
R802 VTAIL.n52 VTAIL.n51 8.14595
R803 VTAIL.n60 VTAIL.n18 8.14595
R804 VTAIL.n98 VTAIL.n0 8.14595
R805 VTAIL.n154 VTAIL.n153 8.14595
R806 VTAIL.n162 VTAIL.n120 8.14595
R807 VTAIL.n200 VTAIL.n102 8.14595
R808 VTAIL.n256 VTAIL.n255 8.14595
R809 VTAIL.n264 VTAIL.n222 8.14595
R810 VTAIL.n302 VTAIL.n204 8.14595
R811 VTAIL.n710 VTAIL.n612 8.14595
R812 VTAIL.n673 VTAIL.n631 8.14595
R813 VTAIL.n665 VTAIL.n664 8.14595
R814 VTAIL.n608 VTAIL.n510 8.14595
R815 VTAIL.n571 VTAIL.n529 8.14595
R816 VTAIL.n563 VTAIL.n562 8.14595
R817 VTAIL.n506 VTAIL.n408 8.14595
R818 VTAIL.n469 VTAIL.n427 8.14595
R819 VTAIL.n461 VTAIL.n460 8.14595
R820 VTAIL.n404 VTAIL.n306 8.14595
R821 VTAIL.n367 VTAIL.n325 8.14595
R822 VTAIL.n359 VTAIL.n358 8.14595
R823 VTAIL.n769 VTAIL.n736 7.3702
R824 VTAIL.n773 VTAIL.n734 7.3702
R825 VTAIL.n55 VTAIL.n22 7.3702
R826 VTAIL.n59 VTAIL.n20 7.3702
R827 VTAIL.n157 VTAIL.n124 7.3702
R828 VTAIL.n161 VTAIL.n122 7.3702
R829 VTAIL.n259 VTAIL.n226 7.3702
R830 VTAIL.n263 VTAIL.n224 7.3702
R831 VTAIL.n672 VTAIL.n633 7.3702
R832 VTAIL.n668 VTAIL.n635 7.3702
R833 VTAIL.n570 VTAIL.n531 7.3702
R834 VTAIL.n566 VTAIL.n533 7.3702
R835 VTAIL.n468 VTAIL.n429 7.3702
R836 VTAIL.n464 VTAIL.n431 7.3702
R837 VTAIL.n366 VTAIL.n327 7.3702
R838 VTAIL.n362 VTAIL.n329 7.3702
R839 VTAIL.n770 VTAIL.n769 6.59444
R840 VTAIL.n770 VTAIL.n734 6.59444
R841 VTAIL.n56 VTAIL.n55 6.59444
R842 VTAIL.n56 VTAIL.n20 6.59444
R843 VTAIL.n158 VTAIL.n157 6.59444
R844 VTAIL.n158 VTAIL.n122 6.59444
R845 VTAIL.n260 VTAIL.n259 6.59444
R846 VTAIL.n260 VTAIL.n224 6.59444
R847 VTAIL.n669 VTAIL.n633 6.59444
R848 VTAIL.n669 VTAIL.n668 6.59444
R849 VTAIL.n567 VTAIL.n531 6.59444
R850 VTAIL.n567 VTAIL.n566 6.59444
R851 VTAIL.n465 VTAIL.n429 6.59444
R852 VTAIL.n465 VTAIL.n464 6.59444
R853 VTAIL.n363 VTAIL.n327 6.59444
R854 VTAIL.n363 VTAIL.n362 6.59444
R855 VTAIL.n766 VTAIL.n736 5.81868
R856 VTAIL.n774 VTAIL.n773 5.81868
R857 VTAIL.n814 VTAIL.n714 5.81868
R858 VTAIL.n52 VTAIL.n22 5.81868
R859 VTAIL.n60 VTAIL.n59 5.81868
R860 VTAIL.n100 VTAIL.n0 5.81868
R861 VTAIL.n154 VTAIL.n124 5.81868
R862 VTAIL.n162 VTAIL.n161 5.81868
R863 VTAIL.n202 VTAIL.n102 5.81868
R864 VTAIL.n256 VTAIL.n226 5.81868
R865 VTAIL.n264 VTAIL.n263 5.81868
R866 VTAIL.n304 VTAIL.n204 5.81868
R867 VTAIL.n712 VTAIL.n612 5.81868
R868 VTAIL.n673 VTAIL.n672 5.81868
R869 VTAIL.n665 VTAIL.n635 5.81868
R870 VTAIL.n610 VTAIL.n510 5.81868
R871 VTAIL.n571 VTAIL.n570 5.81868
R872 VTAIL.n563 VTAIL.n533 5.81868
R873 VTAIL.n508 VTAIL.n408 5.81868
R874 VTAIL.n469 VTAIL.n468 5.81868
R875 VTAIL.n461 VTAIL.n431 5.81868
R876 VTAIL.n406 VTAIL.n306 5.81868
R877 VTAIL.n367 VTAIL.n366 5.81868
R878 VTAIL.n359 VTAIL.n329 5.81868
R879 VTAIL.n765 VTAIL.n738 5.04292
R880 VTAIL.n777 VTAIL.n732 5.04292
R881 VTAIL.n812 VTAIL.n811 5.04292
R882 VTAIL.n51 VTAIL.n24 5.04292
R883 VTAIL.n63 VTAIL.n18 5.04292
R884 VTAIL.n98 VTAIL.n97 5.04292
R885 VTAIL.n153 VTAIL.n126 5.04292
R886 VTAIL.n165 VTAIL.n120 5.04292
R887 VTAIL.n200 VTAIL.n199 5.04292
R888 VTAIL.n255 VTAIL.n228 5.04292
R889 VTAIL.n267 VTAIL.n222 5.04292
R890 VTAIL.n302 VTAIL.n301 5.04292
R891 VTAIL.n710 VTAIL.n709 5.04292
R892 VTAIL.n676 VTAIL.n631 5.04292
R893 VTAIL.n664 VTAIL.n637 5.04292
R894 VTAIL.n608 VTAIL.n607 5.04292
R895 VTAIL.n574 VTAIL.n529 5.04292
R896 VTAIL.n562 VTAIL.n535 5.04292
R897 VTAIL.n506 VTAIL.n505 5.04292
R898 VTAIL.n472 VTAIL.n427 5.04292
R899 VTAIL.n460 VTAIL.n433 5.04292
R900 VTAIL.n404 VTAIL.n403 5.04292
R901 VTAIL.n370 VTAIL.n325 5.04292
R902 VTAIL.n358 VTAIL.n331 5.04292
R903 VTAIL.n748 VTAIL.n747 4.38563
R904 VTAIL.n34 VTAIL.n33 4.38563
R905 VTAIL.n136 VTAIL.n135 4.38563
R906 VTAIL.n238 VTAIL.n237 4.38563
R907 VTAIL.n647 VTAIL.n646 4.38563
R908 VTAIL.n545 VTAIL.n544 4.38563
R909 VTAIL.n443 VTAIL.n442 4.38563
R910 VTAIL.n341 VTAIL.n340 4.38563
R911 VTAIL.n762 VTAIL.n761 4.26717
R912 VTAIL.n778 VTAIL.n730 4.26717
R913 VTAIL.n808 VTAIL.n716 4.26717
R914 VTAIL.n48 VTAIL.n47 4.26717
R915 VTAIL.n64 VTAIL.n16 4.26717
R916 VTAIL.n94 VTAIL.n2 4.26717
R917 VTAIL.n150 VTAIL.n149 4.26717
R918 VTAIL.n166 VTAIL.n118 4.26717
R919 VTAIL.n196 VTAIL.n104 4.26717
R920 VTAIL.n252 VTAIL.n251 4.26717
R921 VTAIL.n268 VTAIL.n220 4.26717
R922 VTAIL.n298 VTAIL.n206 4.26717
R923 VTAIL.n706 VTAIL.n614 4.26717
R924 VTAIL.n677 VTAIL.n629 4.26717
R925 VTAIL.n661 VTAIL.n660 4.26717
R926 VTAIL.n604 VTAIL.n512 4.26717
R927 VTAIL.n575 VTAIL.n527 4.26717
R928 VTAIL.n559 VTAIL.n558 4.26717
R929 VTAIL.n502 VTAIL.n410 4.26717
R930 VTAIL.n473 VTAIL.n425 4.26717
R931 VTAIL.n457 VTAIL.n456 4.26717
R932 VTAIL.n400 VTAIL.n308 4.26717
R933 VTAIL.n371 VTAIL.n323 4.26717
R934 VTAIL.n355 VTAIL.n354 4.26717
R935 VTAIL.n509 VTAIL.n407 3.69878
R936 VTAIL.n713 VTAIL.n611 3.69878
R937 VTAIL.n305 VTAIL.n203 3.69878
R938 VTAIL.n758 VTAIL.n740 3.49141
R939 VTAIL.n782 VTAIL.n781 3.49141
R940 VTAIL.n807 VTAIL.n718 3.49141
R941 VTAIL.n44 VTAIL.n26 3.49141
R942 VTAIL.n68 VTAIL.n67 3.49141
R943 VTAIL.n93 VTAIL.n4 3.49141
R944 VTAIL.n146 VTAIL.n128 3.49141
R945 VTAIL.n170 VTAIL.n169 3.49141
R946 VTAIL.n195 VTAIL.n106 3.49141
R947 VTAIL.n248 VTAIL.n230 3.49141
R948 VTAIL.n272 VTAIL.n271 3.49141
R949 VTAIL.n297 VTAIL.n208 3.49141
R950 VTAIL.n705 VTAIL.n616 3.49141
R951 VTAIL.n681 VTAIL.n680 3.49141
R952 VTAIL.n657 VTAIL.n639 3.49141
R953 VTAIL.n603 VTAIL.n514 3.49141
R954 VTAIL.n579 VTAIL.n578 3.49141
R955 VTAIL.n555 VTAIL.n537 3.49141
R956 VTAIL.n501 VTAIL.n412 3.49141
R957 VTAIL.n477 VTAIL.n476 3.49141
R958 VTAIL.n453 VTAIL.n435 3.49141
R959 VTAIL.n399 VTAIL.n310 3.49141
R960 VTAIL.n375 VTAIL.n374 3.49141
R961 VTAIL.n351 VTAIL.n333 3.49141
R962 VTAIL.n757 VTAIL.n742 2.71565
R963 VTAIL.n785 VTAIL.n728 2.71565
R964 VTAIL.n804 VTAIL.n803 2.71565
R965 VTAIL.n43 VTAIL.n28 2.71565
R966 VTAIL.n71 VTAIL.n14 2.71565
R967 VTAIL.n90 VTAIL.n89 2.71565
R968 VTAIL.n145 VTAIL.n130 2.71565
R969 VTAIL.n173 VTAIL.n116 2.71565
R970 VTAIL.n192 VTAIL.n191 2.71565
R971 VTAIL.n247 VTAIL.n232 2.71565
R972 VTAIL.n275 VTAIL.n218 2.71565
R973 VTAIL.n294 VTAIL.n293 2.71565
R974 VTAIL.n702 VTAIL.n701 2.71565
R975 VTAIL.n684 VTAIL.n627 2.71565
R976 VTAIL.n656 VTAIL.n641 2.71565
R977 VTAIL.n600 VTAIL.n599 2.71565
R978 VTAIL.n582 VTAIL.n525 2.71565
R979 VTAIL.n554 VTAIL.n539 2.71565
R980 VTAIL.n498 VTAIL.n497 2.71565
R981 VTAIL.n480 VTAIL.n423 2.71565
R982 VTAIL.n452 VTAIL.n437 2.71565
R983 VTAIL.n396 VTAIL.n395 2.71565
R984 VTAIL.n378 VTAIL.n321 2.71565
R985 VTAIL.n350 VTAIL.n335 2.71565
R986 VTAIL.n754 VTAIL.n753 1.93989
R987 VTAIL.n786 VTAIL.n726 1.93989
R988 VTAIL.n800 VTAIL.n720 1.93989
R989 VTAIL.n40 VTAIL.n39 1.93989
R990 VTAIL.n72 VTAIL.n12 1.93989
R991 VTAIL.n86 VTAIL.n6 1.93989
R992 VTAIL.n142 VTAIL.n141 1.93989
R993 VTAIL.n174 VTAIL.n114 1.93989
R994 VTAIL.n188 VTAIL.n108 1.93989
R995 VTAIL.n244 VTAIL.n243 1.93989
R996 VTAIL.n276 VTAIL.n216 1.93989
R997 VTAIL.n290 VTAIL.n210 1.93989
R998 VTAIL.n698 VTAIL.n618 1.93989
R999 VTAIL.n685 VTAIL.n625 1.93989
R1000 VTAIL.n653 VTAIL.n652 1.93989
R1001 VTAIL.n596 VTAIL.n516 1.93989
R1002 VTAIL.n583 VTAIL.n523 1.93989
R1003 VTAIL.n551 VTAIL.n550 1.93989
R1004 VTAIL.n494 VTAIL.n414 1.93989
R1005 VTAIL.n481 VTAIL.n421 1.93989
R1006 VTAIL.n449 VTAIL.n448 1.93989
R1007 VTAIL.n392 VTAIL.n312 1.93989
R1008 VTAIL.n379 VTAIL.n319 1.93989
R1009 VTAIL.n347 VTAIL.n346 1.93989
R1010 VTAIL VTAIL.n101 1.90783
R1011 VTAIL VTAIL.n815 1.79145
R1012 VTAIL.n750 VTAIL.n744 1.16414
R1013 VTAIL.n791 VTAIL.n789 1.16414
R1014 VTAIL.n799 VTAIL.n722 1.16414
R1015 VTAIL.n36 VTAIL.n30 1.16414
R1016 VTAIL.n77 VTAIL.n75 1.16414
R1017 VTAIL.n85 VTAIL.n8 1.16414
R1018 VTAIL.n138 VTAIL.n132 1.16414
R1019 VTAIL.n179 VTAIL.n177 1.16414
R1020 VTAIL.n187 VTAIL.n110 1.16414
R1021 VTAIL.n240 VTAIL.n234 1.16414
R1022 VTAIL.n281 VTAIL.n279 1.16414
R1023 VTAIL.n289 VTAIL.n212 1.16414
R1024 VTAIL.n697 VTAIL.n620 1.16414
R1025 VTAIL.n689 VTAIL.n688 1.16414
R1026 VTAIL.n649 VTAIL.n643 1.16414
R1027 VTAIL.n595 VTAIL.n518 1.16414
R1028 VTAIL.n587 VTAIL.n586 1.16414
R1029 VTAIL.n547 VTAIL.n541 1.16414
R1030 VTAIL.n493 VTAIL.n416 1.16414
R1031 VTAIL.n485 VTAIL.n484 1.16414
R1032 VTAIL.n445 VTAIL.n439 1.16414
R1033 VTAIL.n391 VTAIL.n314 1.16414
R1034 VTAIL.n383 VTAIL.n382 1.16414
R1035 VTAIL.n343 VTAIL.n337 1.16414
R1036 VTAIL.n611 VTAIL.n509 0.470328
R1037 VTAIL.n203 VTAIL.n101 0.470328
R1038 VTAIL.n749 VTAIL.n746 0.388379
R1039 VTAIL.n790 VTAIL.n724 0.388379
R1040 VTAIL.n796 VTAIL.n795 0.388379
R1041 VTAIL.n35 VTAIL.n32 0.388379
R1042 VTAIL.n76 VTAIL.n10 0.388379
R1043 VTAIL.n82 VTAIL.n81 0.388379
R1044 VTAIL.n137 VTAIL.n134 0.388379
R1045 VTAIL.n178 VTAIL.n112 0.388379
R1046 VTAIL.n184 VTAIL.n183 0.388379
R1047 VTAIL.n239 VTAIL.n236 0.388379
R1048 VTAIL.n280 VTAIL.n214 0.388379
R1049 VTAIL.n286 VTAIL.n285 0.388379
R1050 VTAIL.n694 VTAIL.n693 0.388379
R1051 VTAIL.n624 VTAIL.n622 0.388379
R1052 VTAIL.n648 VTAIL.n645 0.388379
R1053 VTAIL.n592 VTAIL.n591 0.388379
R1054 VTAIL.n522 VTAIL.n520 0.388379
R1055 VTAIL.n546 VTAIL.n543 0.388379
R1056 VTAIL.n490 VTAIL.n489 0.388379
R1057 VTAIL.n420 VTAIL.n418 0.388379
R1058 VTAIL.n444 VTAIL.n441 0.388379
R1059 VTAIL.n388 VTAIL.n387 0.388379
R1060 VTAIL.n318 VTAIL.n316 0.388379
R1061 VTAIL.n342 VTAIL.n339 0.388379
R1062 VTAIL.n748 VTAIL.n743 0.155672
R1063 VTAIL.n755 VTAIL.n743 0.155672
R1064 VTAIL.n756 VTAIL.n755 0.155672
R1065 VTAIL.n756 VTAIL.n739 0.155672
R1066 VTAIL.n763 VTAIL.n739 0.155672
R1067 VTAIL.n764 VTAIL.n763 0.155672
R1068 VTAIL.n764 VTAIL.n735 0.155672
R1069 VTAIL.n771 VTAIL.n735 0.155672
R1070 VTAIL.n772 VTAIL.n771 0.155672
R1071 VTAIL.n772 VTAIL.n731 0.155672
R1072 VTAIL.n779 VTAIL.n731 0.155672
R1073 VTAIL.n780 VTAIL.n779 0.155672
R1074 VTAIL.n780 VTAIL.n727 0.155672
R1075 VTAIL.n787 VTAIL.n727 0.155672
R1076 VTAIL.n788 VTAIL.n787 0.155672
R1077 VTAIL.n788 VTAIL.n723 0.155672
R1078 VTAIL.n797 VTAIL.n723 0.155672
R1079 VTAIL.n798 VTAIL.n797 0.155672
R1080 VTAIL.n798 VTAIL.n719 0.155672
R1081 VTAIL.n805 VTAIL.n719 0.155672
R1082 VTAIL.n806 VTAIL.n805 0.155672
R1083 VTAIL.n806 VTAIL.n715 0.155672
R1084 VTAIL.n813 VTAIL.n715 0.155672
R1085 VTAIL.n34 VTAIL.n29 0.155672
R1086 VTAIL.n41 VTAIL.n29 0.155672
R1087 VTAIL.n42 VTAIL.n41 0.155672
R1088 VTAIL.n42 VTAIL.n25 0.155672
R1089 VTAIL.n49 VTAIL.n25 0.155672
R1090 VTAIL.n50 VTAIL.n49 0.155672
R1091 VTAIL.n50 VTAIL.n21 0.155672
R1092 VTAIL.n57 VTAIL.n21 0.155672
R1093 VTAIL.n58 VTAIL.n57 0.155672
R1094 VTAIL.n58 VTAIL.n17 0.155672
R1095 VTAIL.n65 VTAIL.n17 0.155672
R1096 VTAIL.n66 VTAIL.n65 0.155672
R1097 VTAIL.n66 VTAIL.n13 0.155672
R1098 VTAIL.n73 VTAIL.n13 0.155672
R1099 VTAIL.n74 VTAIL.n73 0.155672
R1100 VTAIL.n74 VTAIL.n9 0.155672
R1101 VTAIL.n83 VTAIL.n9 0.155672
R1102 VTAIL.n84 VTAIL.n83 0.155672
R1103 VTAIL.n84 VTAIL.n5 0.155672
R1104 VTAIL.n91 VTAIL.n5 0.155672
R1105 VTAIL.n92 VTAIL.n91 0.155672
R1106 VTAIL.n92 VTAIL.n1 0.155672
R1107 VTAIL.n99 VTAIL.n1 0.155672
R1108 VTAIL.n136 VTAIL.n131 0.155672
R1109 VTAIL.n143 VTAIL.n131 0.155672
R1110 VTAIL.n144 VTAIL.n143 0.155672
R1111 VTAIL.n144 VTAIL.n127 0.155672
R1112 VTAIL.n151 VTAIL.n127 0.155672
R1113 VTAIL.n152 VTAIL.n151 0.155672
R1114 VTAIL.n152 VTAIL.n123 0.155672
R1115 VTAIL.n159 VTAIL.n123 0.155672
R1116 VTAIL.n160 VTAIL.n159 0.155672
R1117 VTAIL.n160 VTAIL.n119 0.155672
R1118 VTAIL.n167 VTAIL.n119 0.155672
R1119 VTAIL.n168 VTAIL.n167 0.155672
R1120 VTAIL.n168 VTAIL.n115 0.155672
R1121 VTAIL.n175 VTAIL.n115 0.155672
R1122 VTAIL.n176 VTAIL.n175 0.155672
R1123 VTAIL.n176 VTAIL.n111 0.155672
R1124 VTAIL.n185 VTAIL.n111 0.155672
R1125 VTAIL.n186 VTAIL.n185 0.155672
R1126 VTAIL.n186 VTAIL.n107 0.155672
R1127 VTAIL.n193 VTAIL.n107 0.155672
R1128 VTAIL.n194 VTAIL.n193 0.155672
R1129 VTAIL.n194 VTAIL.n103 0.155672
R1130 VTAIL.n201 VTAIL.n103 0.155672
R1131 VTAIL.n238 VTAIL.n233 0.155672
R1132 VTAIL.n245 VTAIL.n233 0.155672
R1133 VTAIL.n246 VTAIL.n245 0.155672
R1134 VTAIL.n246 VTAIL.n229 0.155672
R1135 VTAIL.n253 VTAIL.n229 0.155672
R1136 VTAIL.n254 VTAIL.n253 0.155672
R1137 VTAIL.n254 VTAIL.n225 0.155672
R1138 VTAIL.n261 VTAIL.n225 0.155672
R1139 VTAIL.n262 VTAIL.n261 0.155672
R1140 VTAIL.n262 VTAIL.n221 0.155672
R1141 VTAIL.n269 VTAIL.n221 0.155672
R1142 VTAIL.n270 VTAIL.n269 0.155672
R1143 VTAIL.n270 VTAIL.n217 0.155672
R1144 VTAIL.n277 VTAIL.n217 0.155672
R1145 VTAIL.n278 VTAIL.n277 0.155672
R1146 VTAIL.n278 VTAIL.n213 0.155672
R1147 VTAIL.n287 VTAIL.n213 0.155672
R1148 VTAIL.n288 VTAIL.n287 0.155672
R1149 VTAIL.n288 VTAIL.n209 0.155672
R1150 VTAIL.n295 VTAIL.n209 0.155672
R1151 VTAIL.n296 VTAIL.n295 0.155672
R1152 VTAIL.n296 VTAIL.n205 0.155672
R1153 VTAIL.n303 VTAIL.n205 0.155672
R1154 VTAIL.n711 VTAIL.n613 0.155672
R1155 VTAIL.n704 VTAIL.n613 0.155672
R1156 VTAIL.n704 VTAIL.n703 0.155672
R1157 VTAIL.n703 VTAIL.n617 0.155672
R1158 VTAIL.n696 VTAIL.n617 0.155672
R1159 VTAIL.n696 VTAIL.n695 0.155672
R1160 VTAIL.n695 VTAIL.n621 0.155672
R1161 VTAIL.n687 VTAIL.n621 0.155672
R1162 VTAIL.n687 VTAIL.n686 0.155672
R1163 VTAIL.n686 VTAIL.n626 0.155672
R1164 VTAIL.n679 VTAIL.n626 0.155672
R1165 VTAIL.n679 VTAIL.n678 0.155672
R1166 VTAIL.n678 VTAIL.n630 0.155672
R1167 VTAIL.n671 VTAIL.n630 0.155672
R1168 VTAIL.n671 VTAIL.n670 0.155672
R1169 VTAIL.n670 VTAIL.n634 0.155672
R1170 VTAIL.n663 VTAIL.n634 0.155672
R1171 VTAIL.n663 VTAIL.n662 0.155672
R1172 VTAIL.n662 VTAIL.n638 0.155672
R1173 VTAIL.n655 VTAIL.n638 0.155672
R1174 VTAIL.n655 VTAIL.n654 0.155672
R1175 VTAIL.n654 VTAIL.n642 0.155672
R1176 VTAIL.n647 VTAIL.n642 0.155672
R1177 VTAIL.n609 VTAIL.n511 0.155672
R1178 VTAIL.n602 VTAIL.n511 0.155672
R1179 VTAIL.n602 VTAIL.n601 0.155672
R1180 VTAIL.n601 VTAIL.n515 0.155672
R1181 VTAIL.n594 VTAIL.n515 0.155672
R1182 VTAIL.n594 VTAIL.n593 0.155672
R1183 VTAIL.n593 VTAIL.n519 0.155672
R1184 VTAIL.n585 VTAIL.n519 0.155672
R1185 VTAIL.n585 VTAIL.n584 0.155672
R1186 VTAIL.n584 VTAIL.n524 0.155672
R1187 VTAIL.n577 VTAIL.n524 0.155672
R1188 VTAIL.n577 VTAIL.n576 0.155672
R1189 VTAIL.n576 VTAIL.n528 0.155672
R1190 VTAIL.n569 VTAIL.n528 0.155672
R1191 VTAIL.n569 VTAIL.n568 0.155672
R1192 VTAIL.n568 VTAIL.n532 0.155672
R1193 VTAIL.n561 VTAIL.n532 0.155672
R1194 VTAIL.n561 VTAIL.n560 0.155672
R1195 VTAIL.n560 VTAIL.n536 0.155672
R1196 VTAIL.n553 VTAIL.n536 0.155672
R1197 VTAIL.n553 VTAIL.n552 0.155672
R1198 VTAIL.n552 VTAIL.n540 0.155672
R1199 VTAIL.n545 VTAIL.n540 0.155672
R1200 VTAIL.n507 VTAIL.n409 0.155672
R1201 VTAIL.n500 VTAIL.n409 0.155672
R1202 VTAIL.n500 VTAIL.n499 0.155672
R1203 VTAIL.n499 VTAIL.n413 0.155672
R1204 VTAIL.n492 VTAIL.n413 0.155672
R1205 VTAIL.n492 VTAIL.n491 0.155672
R1206 VTAIL.n491 VTAIL.n417 0.155672
R1207 VTAIL.n483 VTAIL.n417 0.155672
R1208 VTAIL.n483 VTAIL.n482 0.155672
R1209 VTAIL.n482 VTAIL.n422 0.155672
R1210 VTAIL.n475 VTAIL.n422 0.155672
R1211 VTAIL.n475 VTAIL.n474 0.155672
R1212 VTAIL.n474 VTAIL.n426 0.155672
R1213 VTAIL.n467 VTAIL.n426 0.155672
R1214 VTAIL.n467 VTAIL.n466 0.155672
R1215 VTAIL.n466 VTAIL.n430 0.155672
R1216 VTAIL.n459 VTAIL.n430 0.155672
R1217 VTAIL.n459 VTAIL.n458 0.155672
R1218 VTAIL.n458 VTAIL.n434 0.155672
R1219 VTAIL.n451 VTAIL.n434 0.155672
R1220 VTAIL.n451 VTAIL.n450 0.155672
R1221 VTAIL.n450 VTAIL.n438 0.155672
R1222 VTAIL.n443 VTAIL.n438 0.155672
R1223 VTAIL.n405 VTAIL.n307 0.155672
R1224 VTAIL.n398 VTAIL.n307 0.155672
R1225 VTAIL.n398 VTAIL.n397 0.155672
R1226 VTAIL.n397 VTAIL.n311 0.155672
R1227 VTAIL.n390 VTAIL.n311 0.155672
R1228 VTAIL.n390 VTAIL.n389 0.155672
R1229 VTAIL.n389 VTAIL.n315 0.155672
R1230 VTAIL.n381 VTAIL.n315 0.155672
R1231 VTAIL.n381 VTAIL.n380 0.155672
R1232 VTAIL.n380 VTAIL.n320 0.155672
R1233 VTAIL.n373 VTAIL.n320 0.155672
R1234 VTAIL.n373 VTAIL.n372 0.155672
R1235 VTAIL.n372 VTAIL.n324 0.155672
R1236 VTAIL.n365 VTAIL.n324 0.155672
R1237 VTAIL.n365 VTAIL.n364 0.155672
R1238 VTAIL.n364 VTAIL.n328 0.155672
R1239 VTAIL.n357 VTAIL.n328 0.155672
R1240 VTAIL.n357 VTAIL.n356 0.155672
R1241 VTAIL.n356 VTAIL.n332 0.155672
R1242 VTAIL.n349 VTAIL.n332 0.155672
R1243 VTAIL.n349 VTAIL.n348 0.155672
R1244 VTAIL.n348 VTAIL.n336 0.155672
R1245 VTAIL.n341 VTAIL.n336 0.155672
R1246 B.n773 B.n772 585
R1247 B.n775 B.n155 585
R1248 B.n778 B.n777 585
R1249 B.n779 B.n154 585
R1250 B.n781 B.n780 585
R1251 B.n783 B.n153 585
R1252 B.n786 B.n785 585
R1253 B.n787 B.n152 585
R1254 B.n789 B.n788 585
R1255 B.n791 B.n151 585
R1256 B.n794 B.n793 585
R1257 B.n795 B.n150 585
R1258 B.n797 B.n796 585
R1259 B.n799 B.n149 585
R1260 B.n802 B.n801 585
R1261 B.n803 B.n148 585
R1262 B.n805 B.n804 585
R1263 B.n807 B.n147 585
R1264 B.n810 B.n809 585
R1265 B.n811 B.n146 585
R1266 B.n813 B.n812 585
R1267 B.n815 B.n145 585
R1268 B.n818 B.n817 585
R1269 B.n819 B.n144 585
R1270 B.n821 B.n820 585
R1271 B.n823 B.n143 585
R1272 B.n826 B.n825 585
R1273 B.n827 B.n142 585
R1274 B.n829 B.n828 585
R1275 B.n831 B.n141 585
R1276 B.n834 B.n833 585
R1277 B.n835 B.n140 585
R1278 B.n837 B.n836 585
R1279 B.n839 B.n139 585
R1280 B.n842 B.n841 585
R1281 B.n843 B.n138 585
R1282 B.n845 B.n844 585
R1283 B.n847 B.n137 585
R1284 B.n850 B.n849 585
R1285 B.n851 B.n136 585
R1286 B.n853 B.n852 585
R1287 B.n855 B.n135 585
R1288 B.n858 B.n857 585
R1289 B.n859 B.n134 585
R1290 B.n861 B.n860 585
R1291 B.n863 B.n133 585
R1292 B.n866 B.n865 585
R1293 B.n867 B.n132 585
R1294 B.n869 B.n868 585
R1295 B.n871 B.n131 585
R1296 B.n874 B.n873 585
R1297 B.n875 B.n130 585
R1298 B.n877 B.n876 585
R1299 B.n879 B.n129 585
R1300 B.n882 B.n881 585
R1301 B.n883 B.n128 585
R1302 B.n885 B.n884 585
R1303 B.n887 B.n127 585
R1304 B.n889 B.n888 585
R1305 B.n891 B.n890 585
R1306 B.n894 B.n893 585
R1307 B.n895 B.n122 585
R1308 B.n897 B.n896 585
R1309 B.n899 B.n121 585
R1310 B.n902 B.n901 585
R1311 B.n903 B.n120 585
R1312 B.n905 B.n904 585
R1313 B.n907 B.n119 585
R1314 B.n910 B.n909 585
R1315 B.n911 B.n116 585
R1316 B.n914 B.n913 585
R1317 B.n916 B.n115 585
R1318 B.n919 B.n918 585
R1319 B.n920 B.n114 585
R1320 B.n922 B.n921 585
R1321 B.n924 B.n113 585
R1322 B.n927 B.n926 585
R1323 B.n928 B.n112 585
R1324 B.n930 B.n929 585
R1325 B.n932 B.n111 585
R1326 B.n935 B.n934 585
R1327 B.n936 B.n110 585
R1328 B.n938 B.n937 585
R1329 B.n940 B.n109 585
R1330 B.n943 B.n942 585
R1331 B.n944 B.n108 585
R1332 B.n946 B.n945 585
R1333 B.n948 B.n107 585
R1334 B.n951 B.n950 585
R1335 B.n952 B.n106 585
R1336 B.n954 B.n953 585
R1337 B.n956 B.n105 585
R1338 B.n959 B.n958 585
R1339 B.n960 B.n104 585
R1340 B.n962 B.n961 585
R1341 B.n964 B.n103 585
R1342 B.n967 B.n966 585
R1343 B.n968 B.n102 585
R1344 B.n970 B.n969 585
R1345 B.n972 B.n101 585
R1346 B.n975 B.n974 585
R1347 B.n976 B.n100 585
R1348 B.n978 B.n977 585
R1349 B.n980 B.n99 585
R1350 B.n983 B.n982 585
R1351 B.n984 B.n98 585
R1352 B.n986 B.n985 585
R1353 B.n988 B.n97 585
R1354 B.n991 B.n990 585
R1355 B.n992 B.n96 585
R1356 B.n994 B.n993 585
R1357 B.n996 B.n95 585
R1358 B.n999 B.n998 585
R1359 B.n1000 B.n94 585
R1360 B.n1002 B.n1001 585
R1361 B.n1004 B.n93 585
R1362 B.n1007 B.n1006 585
R1363 B.n1008 B.n92 585
R1364 B.n1010 B.n1009 585
R1365 B.n1012 B.n91 585
R1366 B.n1015 B.n1014 585
R1367 B.n1016 B.n90 585
R1368 B.n1018 B.n1017 585
R1369 B.n1020 B.n89 585
R1370 B.n1023 B.n1022 585
R1371 B.n1024 B.n88 585
R1372 B.n1026 B.n1025 585
R1373 B.n1028 B.n87 585
R1374 B.n1031 B.n1030 585
R1375 B.n1032 B.n86 585
R1376 B.n771 B.n84 585
R1377 B.n1035 B.n84 585
R1378 B.n770 B.n83 585
R1379 B.n1036 B.n83 585
R1380 B.n769 B.n82 585
R1381 B.n1037 B.n82 585
R1382 B.n768 B.n767 585
R1383 B.n767 B.n78 585
R1384 B.n766 B.n77 585
R1385 B.n1043 B.n77 585
R1386 B.n765 B.n76 585
R1387 B.n1044 B.n76 585
R1388 B.n764 B.n75 585
R1389 B.n1045 B.n75 585
R1390 B.n763 B.n762 585
R1391 B.n762 B.n71 585
R1392 B.n761 B.n70 585
R1393 B.n1051 B.n70 585
R1394 B.n760 B.n69 585
R1395 B.n1052 B.n69 585
R1396 B.n759 B.n68 585
R1397 B.n1053 B.n68 585
R1398 B.n758 B.n757 585
R1399 B.n757 B.n64 585
R1400 B.n756 B.n63 585
R1401 B.n1059 B.n63 585
R1402 B.n755 B.n62 585
R1403 B.n1060 B.n62 585
R1404 B.n754 B.n61 585
R1405 B.n1061 B.n61 585
R1406 B.n753 B.n752 585
R1407 B.n752 B.n57 585
R1408 B.n751 B.n56 585
R1409 B.n1067 B.n56 585
R1410 B.n750 B.n55 585
R1411 B.n1068 B.n55 585
R1412 B.n749 B.n54 585
R1413 B.n1069 B.n54 585
R1414 B.n748 B.n747 585
R1415 B.n747 B.n50 585
R1416 B.n746 B.n49 585
R1417 B.n1075 B.n49 585
R1418 B.n745 B.n48 585
R1419 B.n1076 B.n48 585
R1420 B.n744 B.n47 585
R1421 B.n1077 B.n47 585
R1422 B.n743 B.n742 585
R1423 B.n742 B.n43 585
R1424 B.n741 B.n42 585
R1425 B.n1083 B.n42 585
R1426 B.n740 B.n41 585
R1427 B.n1084 B.n41 585
R1428 B.n739 B.n40 585
R1429 B.n1085 B.n40 585
R1430 B.n738 B.n737 585
R1431 B.n737 B.n36 585
R1432 B.n736 B.n35 585
R1433 B.n1091 B.n35 585
R1434 B.n735 B.n34 585
R1435 B.n1092 B.n34 585
R1436 B.n734 B.n33 585
R1437 B.n1093 B.n33 585
R1438 B.n733 B.n732 585
R1439 B.n732 B.n29 585
R1440 B.n731 B.n28 585
R1441 B.n1099 B.n28 585
R1442 B.n730 B.n27 585
R1443 B.n1100 B.n27 585
R1444 B.n729 B.n26 585
R1445 B.n1101 B.n26 585
R1446 B.n728 B.n727 585
R1447 B.n727 B.n22 585
R1448 B.n726 B.n21 585
R1449 B.n1107 B.n21 585
R1450 B.n725 B.n20 585
R1451 B.n1108 B.n20 585
R1452 B.n724 B.n19 585
R1453 B.n1109 B.n19 585
R1454 B.n723 B.n722 585
R1455 B.n722 B.n15 585
R1456 B.n721 B.n14 585
R1457 B.n1115 B.n14 585
R1458 B.n720 B.n13 585
R1459 B.n1116 B.n13 585
R1460 B.n719 B.n12 585
R1461 B.n1117 B.n12 585
R1462 B.n718 B.n717 585
R1463 B.n717 B.n8 585
R1464 B.n716 B.n7 585
R1465 B.n1123 B.n7 585
R1466 B.n715 B.n6 585
R1467 B.n1124 B.n6 585
R1468 B.n714 B.n5 585
R1469 B.n1125 B.n5 585
R1470 B.n713 B.n712 585
R1471 B.n712 B.n4 585
R1472 B.n711 B.n156 585
R1473 B.n711 B.n710 585
R1474 B.n701 B.n157 585
R1475 B.n158 B.n157 585
R1476 B.n703 B.n702 585
R1477 B.n704 B.n703 585
R1478 B.n700 B.n163 585
R1479 B.n163 B.n162 585
R1480 B.n699 B.n698 585
R1481 B.n698 B.n697 585
R1482 B.n165 B.n164 585
R1483 B.n166 B.n165 585
R1484 B.n690 B.n689 585
R1485 B.n691 B.n690 585
R1486 B.n688 B.n171 585
R1487 B.n171 B.n170 585
R1488 B.n687 B.n686 585
R1489 B.n686 B.n685 585
R1490 B.n173 B.n172 585
R1491 B.n174 B.n173 585
R1492 B.n678 B.n677 585
R1493 B.n679 B.n678 585
R1494 B.n676 B.n179 585
R1495 B.n179 B.n178 585
R1496 B.n675 B.n674 585
R1497 B.n674 B.n673 585
R1498 B.n181 B.n180 585
R1499 B.n182 B.n181 585
R1500 B.n666 B.n665 585
R1501 B.n667 B.n666 585
R1502 B.n664 B.n187 585
R1503 B.n187 B.n186 585
R1504 B.n663 B.n662 585
R1505 B.n662 B.n661 585
R1506 B.n189 B.n188 585
R1507 B.n190 B.n189 585
R1508 B.n654 B.n653 585
R1509 B.n655 B.n654 585
R1510 B.n652 B.n194 585
R1511 B.n198 B.n194 585
R1512 B.n651 B.n650 585
R1513 B.n650 B.n649 585
R1514 B.n196 B.n195 585
R1515 B.n197 B.n196 585
R1516 B.n642 B.n641 585
R1517 B.n643 B.n642 585
R1518 B.n640 B.n203 585
R1519 B.n203 B.n202 585
R1520 B.n639 B.n638 585
R1521 B.n638 B.n637 585
R1522 B.n205 B.n204 585
R1523 B.n206 B.n205 585
R1524 B.n630 B.n629 585
R1525 B.n631 B.n630 585
R1526 B.n628 B.n211 585
R1527 B.n211 B.n210 585
R1528 B.n627 B.n626 585
R1529 B.n626 B.n625 585
R1530 B.n213 B.n212 585
R1531 B.n214 B.n213 585
R1532 B.n618 B.n617 585
R1533 B.n619 B.n618 585
R1534 B.n616 B.n219 585
R1535 B.n219 B.n218 585
R1536 B.n615 B.n614 585
R1537 B.n614 B.n613 585
R1538 B.n221 B.n220 585
R1539 B.n222 B.n221 585
R1540 B.n606 B.n605 585
R1541 B.n607 B.n606 585
R1542 B.n604 B.n226 585
R1543 B.n230 B.n226 585
R1544 B.n603 B.n602 585
R1545 B.n602 B.n601 585
R1546 B.n228 B.n227 585
R1547 B.n229 B.n228 585
R1548 B.n594 B.n593 585
R1549 B.n595 B.n594 585
R1550 B.n592 B.n235 585
R1551 B.n235 B.n234 585
R1552 B.n591 B.n590 585
R1553 B.n590 B.n589 585
R1554 B.n237 B.n236 585
R1555 B.n238 B.n237 585
R1556 B.n582 B.n581 585
R1557 B.n583 B.n582 585
R1558 B.n580 B.n243 585
R1559 B.n243 B.n242 585
R1560 B.n579 B.n578 585
R1561 B.n578 B.n577 585
R1562 B.n574 B.n247 585
R1563 B.n573 B.n572 585
R1564 B.n570 B.n248 585
R1565 B.n570 B.n246 585
R1566 B.n569 B.n568 585
R1567 B.n567 B.n566 585
R1568 B.n565 B.n250 585
R1569 B.n563 B.n562 585
R1570 B.n561 B.n251 585
R1571 B.n560 B.n559 585
R1572 B.n557 B.n252 585
R1573 B.n555 B.n554 585
R1574 B.n553 B.n253 585
R1575 B.n552 B.n551 585
R1576 B.n549 B.n254 585
R1577 B.n547 B.n546 585
R1578 B.n545 B.n255 585
R1579 B.n544 B.n543 585
R1580 B.n541 B.n256 585
R1581 B.n539 B.n538 585
R1582 B.n537 B.n257 585
R1583 B.n536 B.n535 585
R1584 B.n533 B.n258 585
R1585 B.n531 B.n530 585
R1586 B.n529 B.n259 585
R1587 B.n528 B.n527 585
R1588 B.n525 B.n260 585
R1589 B.n523 B.n522 585
R1590 B.n521 B.n261 585
R1591 B.n520 B.n519 585
R1592 B.n517 B.n262 585
R1593 B.n515 B.n514 585
R1594 B.n513 B.n263 585
R1595 B.n512 B.n511 585
R1596 B.n509 B.n264 585
R1597 B.n507 B.n506 585
R1598 B.n505 B.n265 585
R1599 B.n504 B.n503 585
R1600 B.n501 B.n266 585
R1601 B.n499 B.n498 585
R1602 B.n497 B.n267 585
R1603 B.n496 B.n495 585
R1604 B.n493 B.n268 585
R1605 B.n491 B.n490 585
R1606 B.n489 B.n269 585
R1607 B.n488 B.n487 585
R1608 B.n485 B.n270 585
R1609 B.n483 B.n482 585
R1610 B.n481 B.n271 585
R1611 B.n480 B.n479 585
R1612 B.n477 B.n272 585
R1613 B.n475 B.n474 585
R1614 B.n473 B.n273 585
R1615 B.n472 B.n471 585
R1616 B.n469 B.n274 585
R1617 B.n467 B.n466 585
R1618 B.n465 B.n275 585
R1619 B.n464 B.n463 585
R1620 B.n461 B.n276 585
R1621 B.n459 B.n458 585
R1622 B.n457 B.n277 585
R1623 B.n455 B.n454 585
R1624 B.n452 B.n280 585
R1625 B.n450 B.n449 585
R1626 B.n448 B.n281 585
R1627 B.n447 B.n446 585
R1628 B.n444 B.n282 585
R1629 B.n442 B.n441 585
R1630 B.n440 B.n283 585
R1631 B.n439 B.n438 585
R1632 B.n436 B.n284 585
R1633 B.n434 B.n433 585
R1634 B.n432 B.n285 585
R1635 B.n431 B.n430 585
R1636 B.n428 B.n289 585
R1637 B.n426 B.n425 585
R1638 B.n424 B.n290 585
R1639 B.n423 B.n422 585
R1640 B.n420 B.n291 585
R1641 B.n418 B.n417 585
R1642 B.n416 B.n292 585
R1643 B.n415 B.n414 585
R1644 B.n412 B.n293 585
R1645 B.n410 B.n409 585
R1646 B.n408 B.n294 585
R1647 B.n407 B.n406 585
R1648 B.n404 B.n295 585
R1649 B.n402 B.n401 585
R1650 B.n400 B.n296 585
R1651 B.n399 B.n398 585
R1652 B.n396 B.n297 585
R1653 B.n394 B.n393 585
R1654 B.n392 B.n298 585
R1655 B.n391 B.n390 585
R1656 B.n388 B.n299 585
R1657 B.n386 B.n385 585
R1658 B.n384 B.n300 585
R1659 B.n383 B.n382 585
R1660 B.n380 B.n301 585
R1661 B.n378 B.n377 585
R1662 B.n376 B.n302 585
R1663 B.n375 B.n374 585
R1664 B.n372 B.n303 585
R1665 B.n370 B.n369 585
R1666 B.n368 B.n304 585
R1667 B.n367 B.n366 585
R1668 B.n364 B.n305 585
R1669 B.n362 B.n361 585
R1670 B.n360 B.n306 585
R1671 B.n359 B.n358 585
R1672 B.n356 B.n307 585
R1673 B.n354 B.n353 585
R1674 B.n352 B.n308 585
R1675 B.n351 B.n350 585
R1676 B.n348 B.n309 585
R1677 B.n346 B.n345 585
R1678 B.n344 B.n310 585
R1679 B.n343 B.n342 585
R1680 B.n340 B.n311 585
R1681 B.n338 B.n337 585
R1682 B.n336 B.n312 585
R1683 B.n335 B.n334 585
R1684 B.n332 B.n313 585
R1685 B.n330 B.n329 585
R1686 B.n328 B.n314 585
R1687 B.n327 B.n326 585
R1688 B.n324 B.n315 585
R1689 B.n322 B.n321 585
R1690 B.n320 B.n316 585
R1691 B.n319 B.n318 585
R1692 B.n245 B.n244 585
R1693 B.n246 B.n245 585
R1694 B.n576 B.n575 585
R1695 B.n577 B.n576 585
R1696 B.n241 B.n240 585
R1697 B.n242 B.n241 585
R1698 B.n585 B.n584 585
R1699 B.n584 B.n583 585
R1700 B.n586 B.n239 585
R1701 B.n239 B.n238 585
R1702 B.n588 B.n587 585
R1703 B.n589 B.n588 585
R1704 B.n233 B.n232 585
R1705 B.n234 B.n233 585
R1706 B.n597 B.n596 585
R1707 B.n596 B.n595 585
R1708 B.n598 B.n231 585
R1709 B.n231 B.n229 585
R1710 B.n600 B.n599 585
R1711 B.n601 B.n600 585
R1712 B.n225 B.n224 585
R1713 B.n230 B.n225 585
R1714 B.n609 B.n608 585
R1715 B.n608 B.n607 585
R1716 B.n610 B.n223 585
R1717 B.n223 B.n222 585
R1718 B.n612 B.n611 585
R1719 B.n613 B.n612 585
R1720 B.n217 B.n216 585
R1721 B.n218 B.n217 585
R1722 B.n621 B.n620 585
R1723 B.n620 B.n619 585
R1724 B.n622 B.n215 585
R1725 B.n215 B.n214 585
R1726 B.n624 B.n623 585
R1727 B.n625 B.n624 585
R1728 B.n209 B.n208 585
R1729 B.n210 B.n209 585
R1730 B.n633 B.n632 585
R1731 B.n632 B.n631 585
R1732 B.n634 B.n207 585
R1733 B.n207 B.n206 585
R1734 B.n636 B.n635 585
R1735 B.n637 B.n636 585
R1736 B.n201 B.n200 585
R1737 B.n202 B.n201 585
R1738 B.n645 B.n644 585
R1739 B.n644 B.n643 585
R1740 B.n646 B.n199 585
R1741 B.n199 B.n197 585
R1742 B.n648 B.n647 585
R1743 B.n649 B.n648 585
R1744 B.n193 B.n192 585
R1745 B.n198 B.n193 585
R1746 B.n657 B.n656 585
R1747 B.n656 B.n655 585
R1748 B.n658 B.n191 585
R1749 B.n191 B.n190 585
R1750 B.n660 B.n659 585
R1751 B.n661 B.n660 585
R1752 B.n185 B.n184 585
R1753 B.n186 B.n185 585
R1754 B.n669 B.n668 585
R1755 B.n668 B.n667 585
R1756 B.n670 B.n183 585
R1757 B.n183 B.n182 585
R1758 B.n672 B.n671 585
R1759 B.n673 B.n672 585
R1760 B.n177 B.n176 585
R1761 B.n178 B.n177 585
R1762 B.n681 B.n680 585
R1763 B.n680 B.n679 585
R1764 B.n682 B.n175 585
R1765 B.n175 B.n174 585
R1766 B.n684 B.n683 585
R1767 B.n685 B.n684 585
R1768 B.n169 B.n168 585
R1769 B.n170 B.n169 585
R1770 B.n693 B.n692 585
R1771 B.n692 B.n691 585
R1772 B.n694 B.n167 585
R1773 B.n167 B.n166 585
R1774 B.n696 B.n695 585
R1775 B.n697 B.n696 585
R1776 B.n161 B.n160 585
R1777 B.n162 B.n161 585
R1778 B.n706 B.n705 585
R1779 B.n705 B.n704 585
R1780 B.n707 B.n159 585
R1781 B.n159 B.n158 585
R1782 B.n709 B.n708 585
R1783 B.n710 B.n709 585
R1784 B.n2 B.n0 585
R1785 B.n4 B.n2 585
R1786 B.n3 B.n1 585
R1787 B.n1124 B.n3 585
R1788 B.n1122 B.n1121 585
R1789 B.n1123 B.n1122 585
R1790 B.n1120 B.n9 585
R1791 B.n9 B.n8 585
R1792 B.n1119 B.n1118 585
R1793 B.n1118 B.n1117 585
R1794 B.n11 B.n10 585
R1795 B.n1116 B.n11 585
R1796 B.n1114 B.n1113 585
R1797 B.n1115 B.n1114 585
R1798 B.n1112 B.n16 585
R1799 B.n16 B.n15 585
R1800 B.n1111 B.n1110 585
R1801 B.n1110 B.n1109 585
R1802 B.n18 B.n17 585
R1803 B.n1108 B.n18 585
R1804 B.n1106 B.n1105 585
R1805 B.n1107 B.n1106 585
R1806 B.n1104 B.n23 585
R1807 B.n23 B.n22 585
R1808 B.n1103 B.n1102 585
R1809 B.n1102 B.n1101 585
R1810 B.n25 B.n24 585
R1811 B.n1100 B.n25 585
R1812 B.n1098 B.n1097 585
R1813 B.n1099 B.n1098 585
R1814 B.n1096 B.n30 585
R1815 B.n30 B.n29 585
R1816 B.n1095 B.n1094 585
R1817 B.n1094 B.n1093 585
R1818 B.n32 B.n31 585
R1819 B.n1092 B.n32 585
R1820 B.n1090 B.n1089 585
R1821 B.n1091 B.n1090 585
R1822 B.n1088 B.n37 585
R1823 B.n37 B.n36 585
R1824 B.n1087 B.n1086 585
R1825 B.n1086 B.n1085 585
R1826 B.n39 B.n38 585
R1827 B.n1084 B.n39 585
R1828 B.n1082 B.n1081 585
R1829 B.n1083 B.n1082 585
R1830 B.n1080 B.n44 585
R1831 B.n44 B.n43 585
R1832 B.n1079 B.n1078 585
R1833 B.n1078 B.n1077 585
R1834 B.n46 B.n45 585
R1835 B.n1076 B.n46 585
R1836 B.n1074 B.n1073 585
R1837 B.n1075 B.n1074 585
R1838 B.n1072 B.n51 585
R1839 B.n51 B.n50 585
R1840 B.n1071 B.n1070 585
R1841 B.n1070 B.n1069 585
R1842 B.n53 B.n52 585
R1843 B.n1068 B.n53 585
R1844 B.n1066 B.n1065 585
R1845 B.n1067 B.n1066 585
R1846 B.n1064 B.n58 585
R1847 B.n58 B.n57 585
R1848 B.n1063 B.n1062 585
R1849 B.n1062 B.n1061 585
R1850 B.n60 B.n59 585
R1851 B.n1060 B.n60 585
R1852 B.n1058 B.n1057 585
R1853 B.n1059 B.n1058 585
R1854 B.n1056 B.n65 585
R1855 B.n65 B.n64 585
R1856 B.n1055 B.n1054 585
R1857 B.n1054 B.n1053 585
R1858 B.n67 B.n66 585
R1859 B.n1052 B.n67 585
R1860 B.n1050 B.n1049 585
R1861 B.n1051 B.n1050 585
R1862 B.n1048 B.n72 585
R1863 B.n72 B.n71 585
R1864 B.n1047 B.n1046 585
R1865 B.n1046 B.n1045 585
R1866 B.n74 B.n73 585
R1867 B.n1044 B.n74 585
R1868 B.n1042 B.n1041 585
R1869 B.n1043 B.n1042 585
R1870 B.n1040 B.n79 585
R1871 B.n79 B.n78 585
R1872 B.n1039 B.n1038 585
R1873 B.n1038 B.n1037 585
R1874 B.n81 B.n80 585
R1875 B.n1036 B.n81 585
R1876 B.n1034 B.n1033 585
R1877 B.n1035 B.n1034 585
R1878 B.n1127 B.n1126 585
R1879 B.n1126 B.n1125 585
R1880 B.n576 B.n247 492.5
R1881 B.n1034 B.n86 492.5
R1882 B.n578 B.n245 492.5
R1883 B.n773 B.n84 492.5
R1884 B.n286 B.t7 474.498
R1885 B.n278 B.t10 474.498
R1886 B.n117 B.t13 474.498
R1887 B.n123 B.t16 474.498
R1888 B.n287 B.t6 391.298
R1889 B.n124 B.t17 391.298
R1890 B.n279 B.t9 391.298
R1891 B.n118 B.t14 391.298
R1892 B.n286 B.t4 320.957
R1893 B.n278 B.t8 320.957
R1894 B.n117 B.t11 320.957
R1895 B.n123 B.t15 320.957
R1896 B.n774 B.n85 256.663
R1897 B.n776 B.n85 256.663
R1898 B.n782 B.n85 256.663
R1899 B.n784 B.n85 256.663
R1900 B.n790 B.n85 256.663
R1901 B.n792 B.n85 256.663
R1902 B.n798 B.n85 256.663
R1903 B.n800 B.n85 256.663
R1904 B.n806 B.n85 256.663
R1905 B.n808 B.n85 256.663
R1906 B.n814 B.n85 256.663
R1907 B.n816 B.n85 256.663
R1908 B.n822 B.n85 256.663
R1909 B.n824 B.n85 256.663
R1910 B.n830 B.n85 256.663
R1911 B.n832 B.n85 256.663
R1912 B.n838 B.n85 256.663
R1913 B.n840 B.n85 256.663
R1914 B.n846 B.n85 256.663
R1915 B.n848 B.n85 256.663
R1916 B.n854 B.n85 256.663
R1917 B.n856 B.n85 256.663
R1918 B.n862 B.n85 256.663
R1919 B.n864 B.n85 256.663
R1920 B.n870 B.n85 256.663
R1921 B.n872 B.n85 256.663
R1922 B.n878 B.n85 256.663
R1923 B.n880 B.n85 256.663
R1924 B.n886 B.n85 256.663
R1925 B.n126 B.n85 256.663
R1926 B.n892 B.n85 256.663
R1927 B.n898 B.n85 256.663
R1928 B.n900 B.n85 256.663
R1929 B.n906 B.n85 256.663
R1930 B.n908 B.n85 256.663
R1931 B.n915 B.n85 256.663
R1932 B.n917 B.n85 256.663
R1933 B.n923 B.n85 256.663
R1934 B.n925 B.n85 256.663
R1935 B.n931 B.n85 256.663
R1936 B.n933 B.n85 256.663
R1937 B.n939 B.n85 256.663
R1938 B.n941 B.n85 256.663
R1939 B.n947 B.n85 256.663
R1940 B.n949 B.n85 256.663
R1941 B.n955 B.n85 256.663
R1942 B.n957 B.n85 256.663
R1943 B.n963 B.n85 256.663
R1944 B.n965 B.n85 256.663
R1945 B.n971 B.n85 256.663
R1946 B.n973 B.n85 256.663
R1947 B.n979 B.n85 256.663
R1948 B.n981 B.n85 256.663
R1949 B.n987 B.n85 256.663
R1950 B.n989 B.n85 256.663
R1951 B.n995 B.n85 256.663
R1952 B.n997 B.n85 256.663
R1953 B.n1003 B.n85 256.663
R1954 B.n1005 B.n85 256.663
R1955 B.n1011 B.n85 256.663
R1956 B.n1013 B.n85 256.663
R1957 B.n1019 B.n85 256.663
R1958 B.n1021 B.n85 256.663
R1959 B.n1027 B.n85 256.663
R1960 B.n1029 B.n85 256.663
R1961 B.n571 B.n246 256.663
R1962 B.n249 B.n246 256.663
R1963 B.n564 B.n246 256.663
R1964 B.n558 B.n246 256.663
R1965 B.n556 B.n246 256.663
R1966 B.n550 B.n246 256.663
R1967 B.n548 B.n246 256.663
R1968 B.n542 B.n246 256.663
R1969 B.n540 B.n246 256.663
R1970 B.n534 B.n246 256.663
R1971 B.n532 B.n246 256.663
R1972 B.n526 B.n246 256.663
R1973 B.n524 B.n246 256.663
R1974 B.n518 B.n246 256.663
R1975 B.n516 B.n246 256.663
R1976 B.n510 B.n246 256.663
R1977 B.n508 B.n246 256.663
R1978 B.n502 B.n246 256.663
R1979 B.n500 B.n246 256.663
R1980 B.n494 B.n246 256.663
R1981 B.n492 B.n246 256.663
R1982 B.n486 B.n246 256.663
R1983 B.n484 B.n246 256.663
R1984 B.n478 B.n246 256.663
R1985 B.n476 B.n246 256.663
R1986 B.n470 B.n246 256.663
R1987 B.n468 B.n246 256.663
R1988 B.n462 B.n246 256.663
R1989 B.n460 B.n246 256.663
R1990 B.n453 B.n246 256.663
R1991 B.n451 B.n246 256.663
R1992 B.n445 B.n246 256.663
R1993 B.n443 B.n246 256.663
R1994 B.n437 B.n246 256.663
R1995 B.n435 B.n246 256.663
R1996 B.n429 B.n246 256.663
R1997 B.n427 B.n246 256.663
R1998 B.n421 B.n246 256.663
R1999 B.n419 B.n246 256.663
R2000 B.n413 B.n246 256.663
R2001 B.n411 B.n246 256.663
R2002 B.n405 B.n246 256.663
R2003 B.n403 B.n246 256.663
R2004 B.n397 B.n246 256.663
R2005 B.n395 B.n246 256.663
R2006 B.n389 B.n246 256.663
R2007 B.n387 B.n246 256.663
R2008 B.n381 B.n246 256.663
R2009 B.n379 B.n246 256.663
R2010 B.n373 B.n246 256.663
R2011 B.n371 B.n246 256.663
R2012 B.n365 B.n246 256.663
R2013 B.n363 B.n246 256.663
R2014 B.n357 B.n246 256.663
R2015 B.n355 B.n246 256.663
R2016 B.n349 B.n246 256.663
R2017 B.n347 B.n246 256.663
R2018 B.n341 B.n246 256.663
R2019 B.n339 B.n246 256.663
R2020 B.n333 B.n246 256.663
R2021 B.n331 B.n246 256.663
R2022 B.n325 B.n246 256.663
R2023 B.n323 B.n246 256.663
R2024 B.n317 B.n246 256.663
R2025 B.n576 B.n241 163.367
R2026 B.n584 B.n241 163.367
R2027 B.n584 B.n239 163.367
R2028 B.n588 B.n239 163.367
R2029 B.n588 B.n233 163.367
R2030 B.n596 B.n233 163.367
R2031 B.n596 B.n231 163.367
R2032 B.n600 B.n231 163.367
R2033 B.n600 B.n225 163.367
R2034 B.n608 B.n225 163.367
R2035 B.n608 B.n223 163.367
R2036 B.n612 B.n223 163.367
R2037 B.n612 B.n217 163.367
R2038 B.n620 B.n217 163.367
R2039 B.n620 B.n215 163.367
R2040 B.n624 B.n215 163.367
R2041 B.n624 B.n209 163.367
R2042 B.n632 B.n209 163.367
R2043 B.n632 B.n207 163.367
R2044 B.n636 B.n207 163.367
R2045 B.n636 B.n201 163.367
R2046 B.n644 B.n201 163.367
R2047 B.n644 B.n199 163.367
R2048 B.n648 B.n199 163.367
R2049 B.n648 B.n193 163.367
R2050 B.n656 B.n193 163.367
R2051 B.n656 B.n191 163.367
R2052 B.n660 B.n191 163.367
R2053 B.n660 B.n185 163.367
R2054 B.n668 B.n185 163.367
R2055 B.n668 B.n183 163.367
R2056 B.n672 B.n183 163.367
R2057 B.n672 B.n177 163.367
R2058 B.n680 B.n177 163.367
R2059 B.n680 B.n175 163.367
R2060 B.n684 B.n175 163.367
R2061 B.n684 B.n169 163.367
R2062 B.n692 B.n169 163.367
R2063 B.n692 B.n167 163.367
R2064 B.n696 B.n167 163.367
R2065 B.n696 B.n161 163.367
R2066 B.n705 B.n161 163.367
R2067 B.n705 B.n159 163.367
R2068 B.n709 B.n159 163.367
R2069 B.n709 B.n2 163.367
R2070 B.n1126 B.n2 163.367
R2071 B.n1126 B.n3 163.367
R2072 B.n1122 B.n3 163.367
R2073 B.n1122 B.n9 163.367
R2074 B.n1118 B.n9 163.367
R2075 B.n1118 B.n11 163.367
R2076 B.n1114 B.n11 163.367
R2077 B.n1114 B.n16 163.367
R2078 B.n1110 B.n16 163.367
R2079 B.n1110 B.n18 163.367
R2080 B.n1106 B.n18 163.367
R2081 B.n1106 B.n23 163.367
R2082 B.n1102 B.n23 163.367
R2083 B.n1102 B.n25 163.367
R2084 B.n1098 B.n25 163.367
R2085 B.n1098 B.n30 163.367
R2086 B.n1094 B.n30 163.367
R2087 B.n1094 B.n32 163.367
R2088 B.n1090 B.n32 163.367
R2089 B.n1090 B.n37 163.367
R2090 B.n1086 B.n37 163.367
R2091 B.n1086 B.n39 163.367
R2092 B.n1082 B.n39 163.367
R2093 B.n1082 B.n44 163.367
R2094 B.n1078 B.n44 163.367
R2095 B.n1078 B.n46 163.367
R2096 B.n1074 B.n46 163.367
R2097 B.n1074 B.n51 163.367
R2098 B.n1070 B.n51 163.367
R2099 B.n1070 B.n53 163.367
R2100 B.n1066 B.n53 163.367
R2101 B.n1066 B.n58 163.367
R2102 B.n1062 B.n58 163.367
R2103 B.n1062 B.n60 163.367
R2104 B.n1058 B.n60 163.367
R2105 B.n1058 B.n65 163.367
R2106 B.n1054 B.n65 163.367
R2107 B.n1054 B.n67 163.367
R2108 B.n1050 B.n67 163.367
R2109 B.n1050 B.n72 163.367
R2110 B.n1046 B.n72 163.367
R2111 B.n1046 B.n74 163.367
R2112 B.n1042 B.n74 163.367
R2113 B.n1042 B.n79 163.367
R2114 B.n1038 B.n79 163.367
R2115 B.n1038 B.n81 163.367
R2116 B.n1034 B.n81 163.367
R2117 B.n572 B.n570 163.367
R2118 B.n570 B.n569 163.367
R2119 B.n566 B.n565 163.367
R2120 B.n563 B.n251 163.367
R2121 B.n559 B.n557 163.367
R2122 B.n555 B.n253 163.367
R2123 B.n551 B.n549 163.367
R2124 B.n547 B.n255 163.367
R2125 B.n543 B.n541 163.367
R2126 B.n539 B.n257 163.367
R2127 B.n535 B.n533 163.367
R2128 B.n531 B.n259 163.367
R2129 B.n527 B.n525 163.367
R2130 B.n523 B.n261 163.367
R2131 B.n519 B.n517 163.367
R2132 B.n515 B.n263 163.367
R2133 B.n511 B.n509 163.367
R2134 B.n507 B.n265 163.367
R2135 B.n503 B.n501 163.367
R2136 B.n499 B.n267 163.367
R2137 B.n495 B.n493 163.367
R2138 B.n491 B.n269 163.367
R2139 B.n487 B.n485 163.367
R2140 B.n483 B.n271 163.367
R2141 B.n479 B.n477 163.367
R2142 B.n475 B.n273 163.367
R2143 B.n471 B.n469 163.367
R2144 B.n467 B.n275 163.367
R2145 B.n463 B.n461 163.367
R2146 B.n459 B.n277 163.367
R2147 B.n454 B.n452 163.367
R2148 B.n450 B.n281 163.367
R2149 B.n446 B.n444 163.367
R2150 B.n442 B.n283 163.367
R2151 B.n438 B.n436 163.367
R2152 B.n434 B.n285 163.367
R2153 B.n430 B.n428 163.367
R2154 B.n426 B.n290 163.367
R2155 B.n422 B.n420 163.367
R2156 B.n418 B.n292 163.367
R2157 B.n414 B.n412 163.367
R2158 B.n410 B.n294 163.367
R2159 B.n406 B.n404 163.367
R2160 B.n402 B.n296 163.367
R2161 B.n398 B.n396 163.367
R2162 B.n394 B.n298 163.367
R2163 B.n390 B.n388 163.367
R2164 B.n386 B.n300 163.367
R2165 B.n382 B.n380 163.367
R2166 B.n378 B.n302 163.367
R2167 B.n374 B.n372 163.367
R2168 B.n370 B.n304 163.367
R2169 B.n366 B.n364 163.367
R2170 B.n362 B.n306 163.367
R2171 B.n358 B.n356 163.367
R2172 B.n354 B.n308 163.367
R2173 B.n350 B.n348 163.367
R2174 B.n346 B.n310 163.367
R2175 B.n342 B.n340 163.367
R2176 B.n338 B.n312 163.367
R2177 B.n334 B.n332 163.367
R2178 B.n330 B.n314 163.367
R2179 B.n326 B.n324 163.367
R2180 B.n322 B.n316 163.367
R2181 B.n318 B.n245 163.367
R2182 B.n578 B.n243 163.367
R2183 B.n582 B.n243 163.367
R2184 B.n582 B.n237 163.367
R2185 B.n590 B.n237 163.367
R2186 B.n590 B.n235 163.367
R2187 B.n594 B.n235 163.367
R2188 B.n594 B.n228 163.367
R2189 B.n602 B.n228 163.367
R2190 B.n602 B.n226 163.367
R2191 B.n606 B.n226 163.367
R2192 B.n606 B.n221 163.367
R2193 B.n614 B.n221 163.367
R2194 B.n614 B.n219 163.367
R2195 B.n618 B.n219 163.367
R2196 B.n618 B.n213 163.367
R2197 B.n626 B.n213 163.367
R2198 B.n626 B.n211 163.367
R2199 B.n630 B.n211 163.367
R2200 B.n630 B.n205 163.367
R2201 B.n638 B.n205 163.367
R2202 B.n638 B.n203 163.367
R2203 B.n642 B.n203 163.367
R2204 B.n642 B.n196 163.367
R2205 B.n650 B.n196 163.367
R2206 B.n650 B.n194 163.367
R2207 B.n654 B.n194 163.367
R2208 B.n654 B.n189 163.367
R2209 B.n662 B.n189 163.367
R2210 B.n662 B.n187 163.367
R2211 B.n666 B.n187 163.367
R2212 B.n666 B.n181 163.367
R2213 B.n674 B.n181 163.367
R2214 B.n674 B.n179 163.367
R2215 B.n678 B.n179 163.367
R2216 B.n678 B.n173 163.367
R2217 B.n686 B.n173 163.367
R2218 B.n686 B.n171 163.367
R2219 B.n690 B.n171 163.367
R2220 B.n690 B.n165 163.367
R2221 B.n698 B.n165 163.367
R2222 B.n698 B.n163 163.367
R2223 B.n703 B.n163 163.367
R2224 B.n703 B.n157 163.367
R2225 B.n711 B.n157 163.367
R2226 B.n712 B.n711 163.367
R2227 B.n712 B.n5 163.367
R2228 B.n6 B.n5 163.367
R2229 B.n7 B.n6 163.367
R2230 B.n717 B.n7 163.367
R2231 B.n717 B.n12 163.367
R2232 B.n13 B.n12 163.367
R2233 B.n14 B.n13 163.367
R2234 B.n722 B.n14 163.367
R2235 B.n722 B.n19 163.367
R2236 B.n20 B.n19 163.367
R2237 B.n21 B.n20 163.367
R2238 B.n727 B.n21 163.367
R2239 B.n727 B.n26 163.367
R2240 B.n27 B.n26 163.367
R2241 B.n28 B.n27 163.367
R2242 B.n732 B.n28 163.367
R2243 B.n732 B.n33 163.367
R2244 B.n34 B.n33 163.367
R2245 B.n35 B.n34 163.367
R2246 B.n737 B.n35 163.367
R2247 B.n737 B.n40 163.367
R2248 B.n41 B.n40 163.367
R2249 B.n42 B.n41 163.367
R2250 B.n742 B.n42 163.367
R2251 B.n742 B.n47 163.367
R2252 B.n48 B.n47 163.367
R2253 B.n49 B.n48 163.367
R2254 B.n747 B.n49 163.367
R2255 B.n747 B.n54 163.367
R2256 B.n55 B.n54 163.367
R2257 B.n56 B.n55 163.367
R2258 B.n752 B.n56 163.367
R2259 B.n752 B.n61 163.367
R2260 B.n62 B.n61 163.367
R2261 B.n63 B.n62 163.367
R2262 B.n757 B.n63 163.367
R2263 B.n757 B.n68 163.367
R2264 B.n69 B.n68 163.367
R2265 B.n70 B.n69 163.367
R2266 B.n762 B.n70 163.367
R2267 B.n762 B.n75 163.367
R2268 B.n76 B.n75 163.367
R2269 B.n77 B.n76 163.367
R2270 B.n767 B.n77 163.367
R2271 B.n767 B.n82 163.367
R2272 B.n83 B.n82 163.367
R2273 B.n84 B.n83 163.367
R2274 B.n1030 B.n1028 163.367
R2275 B.n1026 B.n88 163.367
R2276 B.n1022 B.n1020 163.367
R2277 B.n1018 B.n90 163.367
R2278 B.n1014 B.n1012 163.367
R2279 B.n1010 B.n92 163.367
R2280 B.n1006 B.n1004 163.367
R2281 B.n1002 B.n94 163.367
R2282 B.n998 B.n996 163.367
R2283 B.n994 B.n96 163.367
R2284 B.n990 B.n988 163.367
R2285 B.n986 B.n98 163.367
R2286 B.n982 B.n980 163.367
R2287 B.n978 B.n100 163.367
R2288 B.n974 B.n972 163.367
R2289 B.n970 B.n102 163.367
R2290 B.n966 B.n964 163.367
R2291 B.n962 B.n104 163.367
R2292 B.n958 B.n956 163.367
R2293 B.n954 B.n106 163.367
R2294 B.n950 B.n948 163.367
R2295 B.n946 B.n108 163.367
R2296 B.n942 B.n940 163.367
R2297 B.n938 B.n110 163.367
R2298 B.n934 B.n932 163.367
R2299 B.n930 B.n112 163.367
R2300 B.n926 B.n924 163.367
R2301 B.n922 B.n114 163.367
R2302 B.n918 B.n916 163.367
R2303 B.n914 B.n116 163.367
R2304 B.n909 B.n907 163.367
R2305 B.n905 B.n120 163.367
R2306 B.n901 B.n899 163.367
R2307 B.n897 B.n122 163.367
R2308 B.n893 B.n891 163.367
R2309 B.n888 B.n887 163.367
R2310 B.n885 B.n128 163.367
R2311 B.n881 B.n879 163.367
R2312 B.n877 B.n130 163.367
R2313 B.n873 B.n871 163.367
R2314 B.n869 B.n132 163.367
R2315 B.n865 B.n863 163.367
R2316 B.n861 B.n134 163.367
R2317 B.n857 B.n855 163.367
R2318 B.n853 B.n136 163.367
R2319 B.n849 B.n847 163.367
R2320 B.n845 B.n138 163.367
R2321 B.n841 B.n839 163.367
R2322 B.n837 B.n140 163.367
R2323 B.n833 B.n831 163.367
R2324 B.n829 B.n142 163.367
R2325 B.n825 B.n823 163.367
R2326 B.n821 B.n144 163.367
R2327 B.n817 B.n815 163.367
R2328 B.n813 B.n146 163.367
R2329 B.n809 B.n807 163.367
R2330 B.n805 B.n148 163.367
R2331 B.n801 B.n799 163.367
R2332 B.n797 B.n150 163.367
R2333 B.n793 B.n791 163.367
R2334 B.n789 B.n152 163.367
R2335 B.n785 B.n783 163.367
R2336 B.n781 B.n154 163.367
R2337 B.n777 B.n775 163.367
R2338 B.n287 B.n286 83.2005
R2339 B.n279 B.n278 83.2005
R2340 B.n118 B.n117 83.2005
R2341 B.n124 B.n123 83.2005
R2342 B.n571 B.n247 71.676
R2343 B.n569 B.n249 71.676
R2344 B.n565 B.n564 71.676
R2345 B.n558 B.n251 71.676
R2346 B.n557 B.n556 71.676
R2347 B.n550 B.n253 71.676
R2348 B.n549 B.n548 71.676
R2349 B.n542 B.n255 71.676
R2350 B.n541 B.n540 71.676
R2351 B.n534 B.n257 71.676
R2352 B.n533 B.n532 71.676
R2353 B.n526 B.n259 71.676
R2354 B.n525 B.n524 71.676
R2355 B.n518 B.n261 71.676
R2356 B.n517 B.n516 71.676
R2357 B.n510 B.n263 71.676
R2358 B.n509 B.n508 71.676
R2359 B.n502 B.n265 71.676
R2360 B.n501 B.n500 71.676
R2361 B.n494 B.n267 71.676
R2362 B.n493 B.n492 71.676
R2363 B.n486 B.n269 71.676
R2364 B.n485 B.n484 71.676
R2365 B.n478 B.n271 71.676
R2366 B.n477 B.n476 71.676
R2367 B.n470 B.n273 71.676
R2368 B.n469 B.n468 71.676
R2369 B.n462 B.n275 71.676
R2370 B.n461 B.n460 71.676
R2371 B.n453 B.n277 71.676
R2372 B.n452 B.n451 71.676
R2373 B.n445 B.n281 71.676
R2374 B.n444 B.n443 71.676
R2375 B.n437 B.n283 71.676
R2376 B.n436 B.n435 71.676
R2377 B.n429 B.n285 71.676
R2378 B.n428 B.n427 71.676
R2379 B.n421 B.n290 71.676
R2380 B.n420 B.n419 71.676
R2381 B.n413 B.n292 71.676
R2382 B.n412 B.n411 71.676
R2383 B.n405 B.n294 71.676
R2384 B.n404 B.n403 71.676
R2385 B.n397 B.n296 71.676
R2386 B.n396 B.n395 71.676
R2387 B.n389 B.n298 71.676
R2388 B.n388 B.n387 71.676
R2389 B.n381 B.n300 71.676
R2390 B.n380 B.n379 71.676
R2391 B.n373 B.n302 71.676
R2392 B.n372 B.n371 71.676
R2393 B.n365 B.n304 71.676
R2394 B.n364 B.n363 71.676
R2395 B.n357 B.n306 71.676
R2396 B.n356 B.n355 71.676
R2397 B.n349 B.n308 71.676
R2398 B.n348 B.n347 71.676
R2399 B.n341 B.n310 71.676
R2400 B.n340 B.n339 71.676
R2401 B.n333 B.n312 71.676
R2402 B.n332 B.n331 71.676
R2403 B.n325 B.n314 71.676
R2404 B.n324 B.n323 71.676
R2405 B.n317 B.n316 71.676
R2406 B.n1029 B.n86 71.676
R2407 B.n1028 B.n1027 71.676
R2408 B.n1021 B.n88 71.676
R2409 B.n1020 B.n1019 71.676
R2410 B.n1013 B.n90 71.676
R2411 B.n1012 B.n1011 71.676
R2412 B.n1005 B.n92 71.676
R2413 B.n1004 B.n1003 71.676
R2414 B.n997 B.n94 71.676
R2415 B.n996 B.n995 71.676
R2416 B.n989 B.n96 71.676
R2417 B.n988 B.n987 71.676
R2418 B.n981 B.n98 71.676
R2419 B.n980 B.n979 71.676
R2420 B.n973 B.n100 71.676
R2421 B.n972 B.n971 71.676
R2422 B.n965 B.n102 71.676
R2423 B.n964 B.n963 71.676
R2424 B.n957 B.n104 71.676
R2425 B.n956 B.n955 71.676
R2426 B.n949 B.n106 71.676
R2427 B.n948 B.n947 71.676
R2428 B.n941 B.n108 71.676
R2429 B.n940 B.n939 71.676
R2430 B.n933 B.n110 71.676
R2431 B.n932 B.n931 71.676
R2432 B.n925 B.n112 71.676
R2433 B.n924 B.n923 71.676
R2434 B.n917 B.n114 71.676
R2435 B.n916 B.n915 71.676
R2436 B.n908 B.n116 71.676
R2437 B.n907 B.n906 71.676
R2438 B.n900 B.n120 71.676
R2439 B.n899 B.n898 71.676
R2440 B.n892 B.n122 71.676
R2441 B.n891 B.n126 71.676
R2442 B.n887 B.n886 71.676
R2443 B.n880 B.n128 71.676
R2444 B.n879 B.n878 71.676
R2445 B.n872 B.n130 71.676
R2446 B.n871 B.n870 71.676
R2447 B.n864 B.n132 71.676
R2448 B.n863 B.n862 71.676
R2449 B.n856 B.n134 71.676
R2450 B.n855 B.n854 71.676
R2451 B.n848 B.n136 71.676
R2452 B.n847 B.n846 71.676
R2453 B.n840 B.n138 71.676
R2454 B.n839 B.n838 71.676
R2455 B.n832 B.n140 71.676
R2456 B.n831 B.n830 71.676
R2457 B.n824 B.n142 71.676
R2458 B.n823 B.n822 71.676
R2459 B.n816 B.n144 71.676
R2460 B.n815 B.n814 71.676
R2461 B.n808 B.n146 71.676
R2462 B.n807 B.n806 71.676
R2463 B.n800 B.n148 71.676
R2464 B.n799 B.n798 71.676
R2465 B.n792 B.n150 71.676
R2466 B.n791 B.n790 71.676
R2467 B.n784 B.n152 71.676
R2468 B.n783 B.n782 71.676
R2469 B.n776 B.n154 71.676
R2470 B.n775 B.n774 71.676
R2471 B.n774 B.n773 71.676
R2472 B.n777 B.n776 71.676
R2473 B.n782 B.n781 71.676
R2474 B.n785 B.n784 71.676
R2475 B.n790 B.n789 71.676
R2476 B.n793 B.n792 71.676
R2477 B.n798 B.n797 71.676
R2478 B.n801 B.n800 71.676
R2479 B.n806 B.n805 71.676
R2480 B.n809 B.n808 71.676
R2481 B.n814 B.n813 71.676
R2482 B.n817 B.n816 71.676
R2483 B.n822 B.n821 71.676
R2484 B.n825 B.n824 71.676
R2485 B.n830 B.n829 71.676
R2486 B.n833 B.n832 71.676
R2487 B.n838 B.n837 71.676
R2488 B.n841 B.n840 71.676
R2489 B.n846 B.n845 71.676
R2490 B.n849 B.n848 71.676
R2491 B.n854 B.n853 71.676
R2492 B.n857 B.n856 71.676
R2493 B.n862 B.n861 71.676
R2494 B.n865 B.n864 71.676
R2495 B.n870 B.n869 71.676
R2496 B.n873 B.n872 71.676
R2497 B.n878 B.n877 71.676
R2498 B.n881 B.n880 71.676
R2499 B.n886 B.n885 71.676
R2500 B.n888 B.n126 71.676
R2501 B.n893 B.n892 71.676
R2502 B.n898 B.n897 71.676
R2503 B.n901 B.n900 71.676
R2504 B.n906 B.n905 71.676
R2505 B.n909 B.n908 71.676
R2506 B.n915 B.n914 71.676
R2507 B.n918 B.n917 71.676
R2508 B.n923 B.n922 71.676
R2509 B.n926 B.n925 71.676
R2510 B.n931 B.n930 71.676
R2511 B.n934 B.n933 71.676
R2512 B.n939 B.n938 71.676
R2513 B.n942 B.n941 71.676
R2514 B.n947 B.n946 71.676
R2515 B.n950 B.n949 71.676
R2516 B.n955 B.n954 71.676
R2517 B.n958 B.n957 71.676
R2518 B.n963 B.n962 71.676
R2519 B.n966 B.n965 71.676
R2520 B.n971 B.n970 71.676
R2521 B.n974 B.n973 71.676
R2522 B.n979 B.n978 71.676
R2523 B.n982 B.n981 71.676
R2524 B.n987 B.n986 71.676
R2525 B.n990 B.n989 71.676
R2526 B.n995 B.n994 71.676
R2527 B.n998 B.n997 71.676
R2528 B.n1003 B.n1002 71.676
R2529 B.n1006 B.n1005 71.676
R2530 B.n1011 B.n1010 71.676
R2531 B.n1014 B.n1013 71.676
R2532 B.n1019 B.n1018 71.676
R2533 B.n1022 B.n1021 71.676
R2534 B.n1027 B.n1026 71.676
R2535 B.n1030 B.n1029 71.676
R2536 B.n572 B.n571 71.676
R2537 B.n566 B.n249 71.676
R2538 B.n564 B.n563 71.676
R2539 B.n559 B.n558 71.676
R2540 B.n556 B.n555 71.676
R2541 B.n551 B.n550 71.676
R2542 B.n548 B.n547 71.676
R2543 B.n543 B.n542 71.676
R2544 B.n540 B.n539 71.676
R2545 B.n535 B.n534 71.676
R2546 B.n532 B.n531 71.676
R2547 B.n527 B.n526 71.676
R2548 B.n524 B.n523 71.676
R2549 B.n519 B.n518 71.676
R2550 B.n516 B.n515 71.676
R2551 B.n511 B.n510 71.676
R2552 B.n508 B.n507 71.676
R2553 B.n503 B.n502 71.676
R2554 B.n500 B.n499 71.676
R2555 B.n495 B.n494 71.676
R2556 B.n492 B.n491 71.676
R2557 B.n487 B.n486 71.676
R2558 B.n484 B.n483 71.676
R2559 B.n479 B.n478 71.676
R2560 B.n476 B.n475 71.676
R2561 B.n471 B.n470 71.676
R2562 B.n468 B.n467 71.676
R2563 B.n463 B.n462 71.676
R2564 B.n460 B.n459 71.676
R2565 B.n454 B.n453 71.676
R2566 B.n451 B.n450 71.676
R2567 B.n446 B.n445 71.676
R2568 B.n443 B.n442 71.676
R2569 B.n438 B.n437 71.676
R2570 B.n435 B.n434 71.676
R2571 B.n430 B.n429 71.676
R2572 B.n427 B.n426 71.676
R2573 B.n422 B.n421 71.676
R2574 B.n419 B.n418 71.676
R2575 B.n414 B.n413 71.676
R2576 B.n411 B.n410 71.676
R2577 B.n406 B.n405 71.676
R2578 B.n403 B.n402 71.676
R2579 B.n398 B.n397 71.676
R2580 B.n395 B.n394 71.676
R2581 B.n390 B.n389 71.676
R2582 B.n387 B.n386 71.676
R2583 B.n382 B.n381 71.676
R2584 B.n379 B.n378 71.676
R2585 B.n374 B.n373 71.676
R2586 B.n371 B.n370 71.676
R2587 B.n366 B.n365 71.676
R2588 B.n363 B.n362 71.676
R2589 B.n358 B.n357 71.676
R2590 B.n355 B.n354 71.676
R2591 B.n350 B.n349 71.676
R2592 B.n347 B.n346 71.676
R2593 B.n342 B.n341 71.676
R2594 B.n339 B.n338 71.676
R2595 B.n334 B.n333 71.676
R2596 B.n331 B.n330 71.676
R2597 B.n326 B.n325 71.676
R2598 B.n323 B.n322 71.676
R2599 B.n318 B.n317 71.676
R2600 B.n288 B.n287 59.5399
R2601 B.n456 B.n279 59.5399
R2602 B.n912 B.n118 59.5399
R2603 B.n125 B.n124 59.5399
R2604 B.n577 B.n246 56.4108
R2605 B.n1035 B.n85 56.4108
R2606 B.n1033 B.n1032 32.0005
R2607 B.n772 B.n771 32.0005
R2608 B.n579 B.n244 32.0005
R2609 B.n575 B.n574 32.0005
R2610 B.n577 B.n242 31.7021
R2611 B.n583 B.n242 31.7021
R2612 B.n583 B.n238 31.7021
R2613 B.n589 B.n238 31.7021
R2614 B.n589 B.n234 31.7021
R2615 B.n595 B.n234 31.7021
R2616 B.n595 B.n229 31.7021
R2617 B.n601 B.n229 31.7021
R2618 B.n601 B.n230 31.7021
R2619 B.n607 B.n222 31.7021
R2620 B.n613 B.n222 31.7021
R2621 B.n613 B.n218 31.7021
R2622 B.n619 B.n218 31.7021
R2623 B.n619 B.n214 31.7021
R2624 B.n625 B.n214 31.7021
R2625 B.n625 B.n210 31.7021
R2626 B.n631 B.n210 31.7021
R2627 B.n631 B.n206 31.7021
R2628 B.n637 B.n206 31.7021
R2629 B.n637 B.n202 31.7021
R2630 B.n643 B.n202 31.7021
R2631 B.n643 B.n197 31.7021
R2632 B.n649 B.n197 31.7021
R2633 B.n649 B.n198 31.7021
R2634 B.n655 B.n190 31.7021
R2635 B.n661 B.n190 31.7021
R2636 B.n661 B.n186 31.7021
R2637 B.n667 B.n186 31.7021
R2638 B.n667 B.n182 31.7021
R2639 B.n673 B.n182 31.7021
R2640 B.n673 B.n178 31.7021
R2641 B.n679 B.n178 31.7021
R2642 B.n679 B.n174 31.7021
R2643 B.n685 B.n174 31.7021
R2644 B.n685 B.n170 31.7021
R2645 B.n691 B.n170 31.7021
R2646 B.n697 B.n166 31.7021
R2647 B.n697 B.n162 31.7021
R2648 B.n704 B.n162 31.7021
R2649 B.n704 B.n158 31.7021
R2650 B.n710 B.n158 31.7021
R2651 B.n710 B.n4 31.7021
R2652 B.n1125 B.n4 31.7021
R2653 B.n1125 B.n1124 31.7021
R2654 B.n1124 B.n1123 31.7021
R2655 B.n1123 B.n8 31.7021
R2656 B.n1117 B.n8 31.7021
R2657 B.n1117 B.n1116 31.7021
R2658 B.n1116 B.n1115 31.7021
R2659 B.n1115 B.n15 31.7021
R2660 B.n1109 B.n1108 31.7021
R2661 B.n1108 B.n1107 31.7021
R2662 B.n1107 B.n22 31.7021
R2663 B.n1101 B.n22 31.7021
R2664 B.n1101 B.n1100 31.7021
R2665 B.n1100 B.n1099 31.7021
R2666 B.n1099 B.n29 31.7021
R2667 B.n1093 B.n29 31.7021
R2668 B.n1093 B.n1092 31.7021
R2669 B.n1092 B.n1091 31.7021
R2670 B.n1091 B.n36 31.7021
R2671 B.n1085 B.n36 31.7021
R2672 B.n1084 B.n1083 31.7021
R2673 B.n1083 B.n43 31.7021
R2674 B.n1077 B.n43 31.7021
R2675 B.n1077 B.n1076 31.7021
R2676 B.n1076 B.n1075 31.7021
R2677 B.n1075 B.n50 31.7021
R2678 B.n1069 B.n50 31.7021
R2679 B.n1069 B.n1068 31.7021
R2680 B.n1068 B.n1067 31.7021
R2681 B.n1067 B.n57 31.7021
R2682 B.n1061 B.n57 31.7021
R2683 B.n1061 B.n1060 31.7021
R2684 B.n1060 B.n1059 31.7021
R2685 B.n1059 B.n64 31.7021
R2686 B.n1053 B.n64 31.7021
R2687 B.n1052 B.n1051 31.7021
R2688 B.n1051 B.n71 31.7021
R2689 B.n1045 B.n71 31.7021
R2690 B.n1045 B.n1044 31.7021
R2691 B.n1044 B.n1043 31.7021
R2692 B.n1043 B.n78 31.7021
R2693 B.n1037 B.n78 31.7021
R2694 B.n1037 B.n1036 31.7021
R2695 B.n1036 B.n1035 31.7021
R2696 B.t1 B.n166 28.9049
R2697 B.t0 B.n15 28.9049
R2698 B.n230 B.t5 20.5133
R2699 B.t12 B.n1052 20.5133
R2700 B B.n1127 18.0485
R2701 B.n655 B.t2 16.7837
R2702 B.n1085 B.t3 16.7837
R2703 B.n198 B.t2 14.9189
R2704 B.t3 B.n1084 14.9189
R2705 B.n607 B.t5 11.1893
R2706 B.n1053 B.t12 11.1893
R2707 B.n1032 B.n1031 10.6151
R2708 B.n1031 B.n87 10.6151
R2709 B.n1025 B.n87 10.6151
R2710 B.n1025 B.n1024 10.6151
R2711 B.n1024 B.n1023 10.6151
R2712 B.n1023 B.n89 10.6151
R2713 B.n1017 B.n89 10.6151
R2714 B.n1017 B.n1016 10.6151
R2715 B.n1016 B.n1015 10.6151
R2716 B.n1015 B.n91 10.6151
R2717 B.n1009 B.n91 10.6151
R2718 B.n1009 B.n1008 10.6151
R2719 B.n1008 B.n1007 10.6151
R2720 B.n1007 B.n93 10.6151
R2721 B.n1001 B.n93 10.6151
R2722 B.n1001 B.n1000 10.6151
R2723 B.n1000 B.n999 10.6151
R2724 B.n999 B.n95 10.6151
R2725 B.n993 B.n95 10.6151
R2726 B.n993 B.n992 10.6151
R2727 B.n992 B.n991 10.6151
R2728 B.n991 B.n97 10.6151
R2729 B.n985 B.n97 10.6151
R2730 B.n985 B.n984 10.6151
R2731 B.n984 B.n983 10.6151
R2732 B.n983 B.n99 10.6151
R2733 B.n977 B.n99 10.6151
R2734 B.n977 B.n976 10.6151
R2735 B.n976 B.n975 10.6151
R2736 B.n975 B.n101 10.6151
R2737 B.n969 B.n101 10.6151
R2738 B.n969 B.n968 10.6151
R2739 B.n968 B.n967 10.6151
R2740 B.n967 B.n103 10.6151
R2741 B.n961 B.n103 10.6151
R2742 B.n961 B.n960 10.6151
R2743 B.n960 B.n959 10.6151
R2744 B.n959 B.n105 10.6151
R2745 B.n953 B.n105 10.6151
R2746 B.n953 B.n952 10.6151
R2747 B.n952 B.n951 10.6151
R2748 B.n951 B.n107 10.6151
R2749 B.n945 B.n107 10.6151
R2750 B.n945 B.n944 10.6151
R2751 B.n944 B.n943 10.6151
R2752 B.n943 B.n109 10.6151
R2753 B.n937 B.n109 10.6151
R2754 B.n937 B.n936 10.6151
R2755 B.n936 B.n935 10.6151
R2756 B.n935 B.n111 10.6151
R2757 B.n929 B.n111 10.6151
R2758 B.n929 B.n928 10.6151
R2759 B.n928 B.n927 10.6151
R2760 B.n927 B.n113 10.6151
R2761 B.n921 B.n113 10.6151
R2762 B.n921 B.n920 10.6151
R2763 B.n920 B.n919 10.6151
R2764 B.n919 B.n115 10.6151
R2765 B.n913 B.n115 10.6151
R2766 B.n911 B.n910 10.6151
R2767 B.n910 B.n119 10.6151
R2768 B.n904 B.n119 10.6151
R2769 B.n904 B.n903 10.6151
R2770 B.n903 B.n902 10.6151
R2771 B.n902 B.n121 10.6151
R2772 B.n896 B.n121 10.6151
R2773 B.n896 B.n895 10.6151
R2774 B.n895 B.n894 10.6151
R2775 B.n890 B.n889 10.6151
R2776 B.n889 B.n127 10.6151
R2777 B.n884 B.n127 10.6151
R2778 B.n884 B.n883 10.6151
R2779 B.n883 B.n882 10.6151
R2780 B.n882 B.n129 10.6151
R2781 B.n876 B.n129 10.6151
R2782 B.n876 B.n875 10.6151
R2783 B.n875 B.n874 10.6151
R2784 B.n874 B.n131 10.6151
R2785 B.n868 B.n131 10.6151
R2786 B.n868 B.n867 10.6151
R2787 B.n867 B.n866 10.6151
R2788 B.n866 B.n133 10.6151
R2789 B.n860 B.n133 10.6151
R2790 B.n860 B.n859 10.6151
R2791 B.n859 B.n858 10.6151
R2792 B.n858 B.n135 10.6151
R2793 B.n852 B.n135 10.6151
R2794 B.n852 B.n851 10.6151
R2795 B.n851 B.n850 10.6151
R2796 B.n850 B.n137 10.6151
R2797 B.n844 B.n137 10.6151
R2798 B.n844 B.n843 10.6151
R2799 B.n843 B.n842 10.6151
R2800 B.n842 B.n139 10.6151
R2801 B.n836 B.n139 10.6151
R2802 B.n836 B.n835 10.6151
R2803 B.n835 B.n834 10.6151
R2804 B.n834 B.n141 10.6151
R2805 B.n828 B.n141 10.6151
R2806 B.n828 B.n827 10.6151
R2807 B.n827 B.n826 10.6151
R2808 B.n826 B.n143 10.6151
R2809 B.n820 B.n143 10.6151
R2810 B.n820 B.n819 10.6151
R2811 B.n819 B.n818 10.6151
R2812 B.n818 B.n145 10.6151
R2813 B.n812 B.n145 10.6151
R2814 B.n812 B.n811 10.6151
R2815 B.n811 B.n810 10.6151
R2816 B.n810 B.n147 10.6151
R2817 B.n804 B.n147 10.6151
R2818 B.n804 B.n803 10.6151
R2819 B.n803 B.n802 10.6151
R2820 B.n802 B.n149 10.6151
R2821 B.n796 B.n149 10.6151
R2822 B.n796 B.n795 10.6151
R2823 B.n795 B.n794 10.6151
R2824 B.n794 B.n151 10.6151
R2825 B.n788 B.n151 10.6151
R2826 B.n788 B.n787 10.6151
R2827 B.n787 B.n786 10.6151
R2828 B.n786 B.n153 10.6151
R2829 B.n780 B.n153 10.6151
R2830 B.n780 B.n779 10.6151
R2831 B.n779 B.n778 10.6151
R2832 B.n778 B.n155 10.6151
R2833 B.n772 B.n155 10.6151
R2834 B.n580 B.n579 10.6151
R2835 B.n581 B.n580 10.6151
R2836 B.n581 B.n236 10.6151
R2837 B.n591 B.n236 10.6151
R2838 B.n592 B.n591 10.6151
R2839 B.n593 B.n592 10.6151
R2840 B.n593 B.n227 10.6151
R2841 B.n603 B.n227 10.6151
R2842 B.n604 B.n603 10.6151
R2843 B.n605 B.n604 10.6151
R2844 B.n605 B.n220 10.6151
R2845 B.n615 B.n220 10.6151
R2846 B.n616 B.n615 10.6151
R2847 B.n617 B.n616 10.6151
R2848 B.n617 B.n212 10.6151
R2849 B.n627 B.n212 10.6151
R2850 B.n628 B.n627 10.6151
R2851 B.n629 B.n628 10.6151
R2852 B.n629 B.n204 10.6151
R2853 B.n639 B.n204 10.6151
R2854 B.n640 B.n639 10.6151
R2855 B.n641 B.n640 10.6151
R2856 B.n641 B.n195 10.6151
R2857 B.n651 B.n195 10.6151
R2858 B.n652 B.n651 10.6151
R2859 B.n653 B.n652 10.6151
R2860 B.n653 B.n188 10.6151
R2861 B.n663 B.n188 10.6151
R2862 B.n664 B.n663 10.6151
R2863 B.n665 B.n664 10.6151
R2864 B.n665 B.n180 10.6151
R2865 B.n675 B.n180 10.6151
R2866 B.n676 B.n675 10.6151
R2867 B.n677 B.n676 10.6151
R2868 B.n677 B.n172 10.6151
R2869 B.n687 B.n172 10.6151
R2870 B.n688 B.n687 10.6151
R2871 B.n689 B.n688 10.6151
R2872 B.n689 B.n164 10.6151
R2873 B.n699 B.n164 10.6151
R2874 B.n700 B.n699 10.6151
R2875 B.n702 B.n700 10.6151
R2876 B.n702 B.n701 10.6151
R2877 B.n701 B.n156 10.6151
R2878 B.n713 B.n156 10.6151
R2879 B.n714 B.n713 10.6151
R2880 B.n715 B.n714 10.6151
R2881 B.n716 B.n715 10.6151
R2882 B.n718 B.n716 10.6151
R2883 B.n719 B.n718 10.6151
R2884 B.n720 B.n719 10.6151
R2885 B.n721 B.n720 10.6151
R2886 B.n723 B.n721 10.6151
R2887 B.n724 B.n723 10.6151
R2888 B.n725 B.n724 10.6151
R2889 B.n726 B.n725 10.6151
R2890 B.n728 B.n726 10.6151
R2891 B.n729 B.n728 10.6151
R2892 B.n730 B.n729 10.6151
R2893 B.n731 B.n730 10.6151
R2894 B.n733 B.n731 10.6151
R2895 B.n734 B.n733 10.6151
R2896 B.n735 B.n734 10.6151
R2897 B.n736 B.n735 10.6151
R2898 B.n738 B.n736 10.6151
R2899 B.n739 B.n738 10.6151
R2900 B.n740 B.n739 10.6151
R2901 B.n741 B.n740 10.6151
R2902 B.n743 B.n741 10.6151
R2903 B.n744 B.n743 10.6151
R2904 B.n745 B.n744 10.6151
R2905 B.n746 B.n745 10.6151
R2906 B.n748 B.n746 10.6151
R2907 B.n749 B.n748 10.6151
R2908 B.n750 B.n749 10.6151
R2909 B.n751 B.n750 10.6151
R2910 B.n753 B.n751 10.6151
R2911 B.n754 B.n753 10.6151
R2912 B.n755 B.n754 10.6151
R2913 B.n756 B.n755 10.6151
R2914 B.n758 B.n756 10.6151
R2915 B.n759 B.n758 10.6151
R2916 B.n760 B.n759 10.6151
R2917 B.n761 B.n760 10.6151
R2918 B.n763 B.n761 10.6151
R2919 B.n764 B.n763 10.6151
R2920 B.n765 B.n764 10.6151
R2921 B.n766 B.n765 10.6151
R2922 B.n768 B.n766 10.6151
R2923 B.n769 B.n768 10.6151
R2924 B.n770 B.n769 10.6151
R2925 B.n771 B.n770 10.6151
R2926 B.n574 B.n573 10.6151
R2927 B.n573 B.n248 10.6151
R2928 B.n568 B.n248 10.6151
R2929 B.n568 B.n567 10.6151
R2930 B.n567 B.n250 10.6151
R2931 B.n562 B.n250 10.6151
R2932 B.n562 B.n561 10.6151
R2933 B.n561 B.n560 10.6151
R2934 B.n560 B.n252 10.6151
R2935 B.n554 B.n252 10.6151
R2936 B.n554 B.n553 10.6151
R2937 B.n553 B.n552 10.6151
R2938 B.n552 B.n254 10.6151
R2939 B.n546 B.n254 10.6151
R2940 B.n546 B.n545 10.6151
R2941 B.n545 B.n544 10.6151
R2942 B.n544 B.n256 10.6151
R2943 B.n538 B.n256 10.6151
R2944 B.n538 B.n537 10.6151
R2945 B.n537 B.n536 10.6151
R2946 B.n536 B.n258 10.6151
R2947 B.n530 B.n258 10.6151
R2948 B.n530 B.n529 10.6151
R2949 B.n529 B.n528 10.6151
R2950 B.n528 B.n260 10.6151
R2951 B.n522 B.n260 10.6151
R2952 B.n522 B.n521 10.6151
R2953 B.n521 B.n520 10.6151
R2954 B.n520 B.n262 10.6151
R2955 B.n514 B.n262 10.6151
R2956 B.n514 B.n513 10.6151
R2957 B.n513 B.n512 10.6151
R2958 B.n512 B.n264 10.6151
R2959 B.n506 B.n264 10.6151
R2960 B.n506 B.n505 10.6151
R2961 B.n505 B.n504 10.6151
R2962 B.n504 B.n266 10.6151
R2963 B.n498 B.n266 10.6151
R2964 B.n498 B.n497 10.6151
R2965 B.n497 B.n496 10.6151
R2966 B.n496 B.n268 10.6151
R2967 B.n490 B.n268 10.6151
R2968 B.n490 B.n489 10.6151
R2969 B.n489 B.n488 10.6151
R2970 B.n488 B.n270 10.6151
R2971 B.n482 B.n270 10.6151
R2972 B.n482 B.n481 10.6151
R2973 B.n481 B.n480 10.6151
R2974 B.n480 B.n272 10.6151
R2975 B.n474 B.n272 10.6151
R2976 B.n474 B.n473 10.6151
R2977 B.n473 B.n472 10.6151
R2978 B.n472 B.n274 10.6151
R2979 B.n466 B.n274 10.6151
R2980 B.n466 B.n465 10.6151
R2981 B.n465 B.n464 10.6151
R2982 B.n464 B.n276 10.6151
R2983 B.n458 B.n276 10.6151
R2984 B.n458 B.n457 10.6151
R2985 B.n455 B.n280 10.6151
R2986 B.n449 B.n280 10.6151
R2987 B.n449 B.n448 10.6151
R2988 B.n448 B.n447 10.6151
R2989 B.n447 B.n282 10.6151
R2990 B.n441 B.n282 10.6151
R2991 B.n441 B.n440 10.6151
R2992 B.n440 B.n439 10.6151
R2993 B.n439 B.n284 10.6151
R2994 B.n433 B.n432 10.6151
R2995 B.n432 B.n431 10.6151
R2996 B.n431 B.n289 10.6151
R2997 B.n425 B.n289 10.6151
R2998 B.n425 B.n424 10.6151
R2999 B.n424 B.n423 10.6151
R3000 B.n423 B.n291 10.6151
R3001 B.n417 B.n291 10.6151
R3002 B.n417 B.n416 10.6151
R3003 B.n416 B.n415 10.6151
R3004 B.n415 B.n293 10.6151
R3005 B.n409 B.n293 10.6151
R3006 B.n409 B.n408 10.6151
R3007 B.n408 B.n407 10.6151
R3008 B.n407 B.n295 10.6151
R3009 B.n401 B.n295 10.6151
R3010 B.n401 B.n400 10.6151
R3011 B.n400 B.n399 10.6151
R3012 B.n399 B.n297 10.6151
R3013 B.n393 B.n297 10.6151
R3014 B.n393 B.n392 10.6151
R3015 B.n392 B.n391 10.6151
R3016 B.n391 B.n299 10.6151
R3017 B.n385 B.n299 10.6151
R3018 B.n385 B.n384 10.6151
R3019 B.n384 B.n383 10.6151
R3020 B.n383 B.n301 10.6151
R3021 B.n377 B.n301 10.6151
R3022 B.n377 B.n376 10.6151
R3023 B.n376 B.n375 10.6151
R3024 B.n375 B.n303 10.6151
R3025 B.n369 B.n303 10.6151
R3026 B.n369 B.n368 10.6151
R3027 B.n368 B.n367 10.6151
R3028 B.n367 B.n305 10.6151
R3029 B.n361 B.n305 10.6151
R3030 B.n361 B.n360 10.6151
R3031 B.n360 B.n359 10.6151
R3032 B.n359 B.n307 10.6151
R3033 B.n353 B.n307 10.6151
R3034 B.n353 B.n352 10.6151
R3035 B.n352 B.n351 10.6151
R3036 B.n351 B.n309 10.6151
R3037 B.n345 B.n309 10.6151
R3038 B.n345 B.n344 10.6151
R3039 B.n344 B.n343 10.6151
R3040 B.n343 B.n311 10.6151
R3041 B.n337 B.n311 10.6151
R3042 B.n337 B.n336 10.6151
R3043 B.n336 B.n335 10.6151
R3044 B.n335 B.n313 10.6151
R3045 B.n329 B.n313 10.6151
R3046 B.n329 B.n328 10.6151
R3047 B.n328 B.n327 10.6151
R3048 B.n327 B.n315 10.6151
R3049 B.n321 B.n315 10.6151
R3050 B.n321 B.n320 10.6151
R3051 B.n320 B.n319 10.6151
R3052 B.n319 B.n244 10.6151
R3053 B.n575 B.n240 10.6151
R3054 B.n585 B.n240 10.6151
R3055 B.n586 B.n585 10.6151
R3056 B.n587 B.n586 10.6151
R3057 B.n587 B.n232 10.6151
R3058 B.n597 B.n232 10.6151
R3059 B.n598 B.n597 10.6151
R3060 B.n599 B.n598 10.6151
R3061 B.n599 B.n224 10.6151
R3062 B.n609 B.n224 10.6151
R3063 B.n610 B.n609 10.6151
R3064 B.n611 B.n610 10.6151
R3065 B.n611 B.n216 10.6151
R3066 B.n621 B.n216 10.6151
R3067 B.n622 B.n621 10.6151
R3068 B.n623 B.n622 10.6151
R3069 B.n623 B.n208 10.6151
R3070 B.n633 B.n208 10.6151
R3071 B.n634 B.n633 10.6151
R3072 B.n635 B.n634 10.6151
R3073 B.n635 B.n200 10.6151
R3074 B.n645 B.n200 10.6151
R3075 B.n646 B.n645 10.6151
R3076 B.n647 B.n646 10.6151
R3077 B.n647 B.n192 10.6151
R3078 B.n657 B.n192 10.6151
R3079 B.n658 B.n657 10.6151
R3080 B.n659 B.n658 10.6151
R3081 B.n659 B.n184 10.6151
R3082 B.n669 B.n184 10.6151
R3083 B.n670 B.n669 10.6151
R3084 B.n671 B.n670 10.6151
R3085 B.n671 B.n176 10.6151
R3086 B.n681 B.n176 10.6151
R3087 B.n682 B.n681 10.6151
R3088 B.n683 B.n682 10.6151
R3089 B.n683 B.n168 10.6151
R3090 B.n693 B.n168 10.6151
R3091 B.n694 B.n693 10.6151
R3092 B.n695 B.n694 10.6151
R3093 B.n695 B.n160 10.6151
R3094 B.n706 B.n160 10.6151
R3095 B.n707 B.n706 10.6151
R3096 B.n708 B.n707 10.6151
R3097 B.n708 B.n0 10.6151
R3098 B.n1121 B.n1 10.6151
R3099 B.n1121 B.n1120 10.6151
R3100 B.n1120 B.n1119 10.6151
R3101 B.n1119 B.n10 10.6151
R3102 B.n1113 B.n10 10.6151
R3103 B.n1113 B.n1112 10.6151
R3104 B.n1112 B.n1111 10.6151
R3105 B.n1111 B.n17 10.6151
R3106 B.n1105 B.n17 10.6151
R3107 B.n1105 B.n1104 10.6151
R3108 B.n1104 B.n1103 10.6151
R3109 B.n1103 B.n24 10.6151
R3110 B.n1097 B.n24 10.6151
R3111 B.n1097 B.n1096 10.6151
R3112 B.n1096 B.n1095 10.6151
R3113 B.n1095 B.n31 10.6151
R3114 B.n1089 B.n31 10.6151
R3115 B.n1089 B.n1088 10.6151
R3116 B.n1088 B.n1087 10.6151
R3117 B.n1087 B.n38 10.6151
R3118 B.n1081 B.n38 10.6151
R3119 B.n1081 B.n1080 10.6151
R3120 B.n1080 B.n1079 10.6151
R3121 B.n1079 B.n45 10.6151
R3122 B.n1073 B.n45 10.6151
R3123 B.n1073 B.n1072 10.6151
R3124 B.n1072 B.n1071 10.6151
R3125 B.n1071 B.n52 10.6151
R3126 B.n1065 B.n52 10.6151
R3127 B.n1065 B.n1064 10.6151
R3128 B.n1064 B.n1063 10.6151
R3129 B.n1063 B.n59 10.6151
R3130 B.n1057 B.n59 10.6151
R3131 B.n1057 B.n1056 10.6151
R3132 B.n1056 B.n1055 10.6151
R3133 B.n1055 B.n66 10.6151
R3134 B.n1049 B.n66 10.6151
R3135 B.n1049 B.n1048 10.6151
R3136 B.n1048 B.n1047 10.6151
R3137 B.n1047 B.n73 10.6151
R3138 B.n1041 B.n73 10.6151
R3139 B.n1041 B.n1040 10.6151
R3140 B.n1040 B.n1039 10.6151
R3141 B.n1039 B.n80 10.6151
R3142 B.n1033 B.n80 10.6151
R3143 B.n913 B.n912 9.36635
R3144 B.n890 B.n125 9.36635
R3145 B.n457 B.n456 9.36635
R3146 B.n433 B.n288 9.36635
R3147 B.n1127 B.n0 2.81026
R3148 B.n1127 B.n1 2.81026
R3149 B.n691 B.t1 2.7977
R3150 B.n1109 B.t0 2.7977
R3151 B.n912 B.n911 1.24928
R3152 B.n894 B.n125 1.24928
R3153 B.n456 B.n455 1.24928
R3154 B.n288 B.n284 1.24928
R3155 VP.n18 VP.n0 161.3
R3156 VP.n17 VP.n16 161.3
R3157 VP.n15 VP.n1 161.3
R3158 VP.n14 VP.n13 161.3
R3159 VP.n12 VP.n2 161.3
R3160 VP.n11 VP.n10 161.3
R3161 VP.n9 VP.n3 161.3
R3162 VP.n8 VP.n7 161.3
R3163 VP.n4 VP.t2 145.382
R3164 VP.n4 VP.t0 143.946
R3165 VP.n6 VP.t1 111.493
R3166 VP.n19 VP.t3 111.493
R3167 VP.n6 VP.n5 62.9523
R3168 VP.n20 VP.n19 62.9523
R3169 VP.n5 VP.n4 57.1277
R3170 VP.n13 VP.n12 56.5617
R3171 VP.n7 VP.n3 24.5923
R3172 VP.n11 VP.n3 24.5923
R3173 VP.n12 VP.n11 24.5923
R3174 VP.n13 VP.n1 24.5923
R3175 VP.n17 VP.n1 24.5923
R3176 VP.n18 VP.n17 24.5923
R3177 VP.n7 VP.n6 19.4281
R3178 VP.n19 VP.n18 19.4281
R3179 VP.n8 VP.n5 0.417304
R3180 VP.n20 VP.n0 0.417304
R3181 VP VP.n20 0.394524
R3182 VP.n9 VP.n8 0.189894
R3183 VP.n10 VP.n9 0.189894
R3184 VP.n10 VP.n2 0.189894
R3185 VP.n14 VP.n2 0.189894
R3186 VP.n15 VP.n14 0.189894
R3187 VP.n16 VP.n15 0.189894
R3188 VP.n16 VP.n0 0.189894
R3189 VDD1 VDD1.n1 113.328
R3190 VDD1 VDD1.n0 62.2578
R3191 VDD1.n0 VDD1.t1 1.08129
R3192 VDD1.n0 VDD1.t3 1.08129
R3193 VDD1.n1 VDD1.t2 1.08129
R3194 VDD1.n1 VDD1.t0 1.08129
C0 VP VN 8.33989f
C1 VP VDD2 0.481336f
C2 VP VTAIL 7.37065f
C3 VN VDD1 0.150721f
C4 VDD1 VDD2 1.36149f
C5 VN VDD2 7.545939f
C6 VTAIL VDD1 7.10823f
C7 VN VTAIL 7.35654f
C8 VTAIL VDD2 7.17155f
C9 VP VDD1 7.87547f
C10 VDD2 B 5.021659f
C11 VDD1 B 10.28737f
C12 VTAIL B 14.66905f
C13 VN B 13.82583f
C14 VP B 12.270749f
C15 VDD1.t1 B 0.392536f
C16 VDD1.t3 B 0.392536f
C17 VDD1.n0 B 3.58073f
C18 VDD1.t2 B 0.392536f
C19 VDD1.t0 B 0.392536f
C20 VDD1.n1 B 4.60596f
C21 VP.n0 B 0.034525f
C22 VP.t3 B 3.66486f
C23 VP.n1 B 0.034047f
C24 VP.n2 B 0.01836f
C25 VP.n3 B 0.034047f
C26 VP.t0 B 3.98083f
C27 VP.t2 B 3.99417f
C28 VP.n4 B 3.78422f
C29 VP.n5 B 1.28905f
C30 VP.t1 B 3.66486f
C31 VP.n6 B 1.33971f
C32 VP.n7 B 0.030517f
C33 VP.n8 B 0.034525f
C34 VP.n9 B 0.01836f
C35 VP.n10 B 0.01836f
C36 VP.n11 B 0.034047f
C37 VP.n12 B 0.026689f
C38 VP.n13 B 0.026689f
C39 VP.n14 B 0.01836f
C40 VP.n15 B 0.01836f
C41 VP.n16 B 0.01836f
C42 VP.n17 B 0.034047f
C43 VP.n18 B 0.030517f
C44 VP.n19 B 1.33971f
C45 VP.n20 B 0.059226f
C46 VTAIL.n0 B 0.023155f
C47 VTAIL.n1 B 0.015864f
C48 VTAIL.n2 B 0.008525f
C49 VTAIL.n3 B 0.02015f
C50 VTAIL.n4 B 0.009026f
C51 VTAIL.n5 B 0.015864f
C52 VTAIL.n6 B 0.008525f
C53 VTAIL.n7 B 0.02015f
C54 VTAIL.n8 B 0.009026f
C55 VTAIL.n9 B 0.015864f
C56 VTAIL.n10 B 0.008776f
C57 VTAIL.n11 B 0.02015f
C58 VTAIL.n12 B 0.009026f
C59 VTAIL.n13 B 0.015864f
C60 VTAIL.n14 B 0.008525f
C61 VTAIL.n15 B 0.02015f
C62 VTAIL.n16 B 0.009026f
C63 VTAIL.n17 B 0.015864f
C64 VTAIL.n18 B 0.008525f
C65 VTAIL.n19 B 0.02015f
C66 VTAIL.n20 B 0.009026f
C67 VTAIL.n21 B 0.015864f
C68 VTAIL.n22 B 0.008525f
C69 VTAIL.n23 B 0.02015f
C70 VTAIL.n24 B 0.009026f
C71 VTAIL.n25 B 0.015864f
C72 VTAIL.n26 B 0.008525f
C73 VTAIL.n27 B 0.02015f
C74 VTAIL.n28 B 0.009026f
C75 VTAIL.n29 B 0.015864f
C76 VTAIL.n30 B 0.008525f
C77 VTAIL.n31 B 0.015112f
C78 VTAIL.n32 B 0.011903f
C79 VTAIL.t7 B 0.033405f
C80 VTAIL.n33 B 0.116676f
C81 VTAIL.n34 B 1.27354f
C82 VTAIL.n35 B 0.008525f
C83 VTAIL.n36 B 0.009026f
C84 VTAIL.n37 B 0.02015f
C85 VTAIL.n38 B 0.02015f
C86 VTAIL.n39 B 0.009026f
C87 VTAIL.n40 B 0.008525f
C88 VTAIL.n41 B 0.015864f
C89 VTAIL.n42 B 0.015864f
C90 VTAIL.n43 B 0.008525f
C91 VTAIL.n44 B 0.009026f
C92 VTAIL.n45 B 0.02015f
C93 VTAIL.n46 B 0.02015f
C94 VTAIL.n47 B 0.009026f
C95 VTAIL.n48 B 0.008525f
C96 VTAIL.n49 B 0.015864f
C97 VTAIL.n50 B 0.015864f
C98 VTAIL.n51 B 0.008525f
C99 VTAIL.n52 B 0.009026f
C100 VTAIL.n53 B 0.02015f
C101 VTAIL.n54 B 0.02015f
C102 VTAIL.n55 B 0.009026f
C103 VTAIL.n56 B 0.008525f
C104 VTAIL.n57 B 0.015864f
C105 VTAIL.n58 B 0.015864f
C106 VTAIL.n59 B 0.008525f
C107 VTAIL.n60 B 0.009026f
C108 VTAIL.n61 B 0.02015f
C109 VTAIL.n62 B 0.02015f
C110 VTAIL.n63 B 0.009026f
C111 VTAIL.n64 B 0.008525f
C112 VTAIL.n65 B 0.015864f
C113 VTAIL.n66 B 0.015864f
C114 VTAIL.n67 B 0.008525f
C115 VTAIL.n68 B 0.009026f
C116 VTAIL.n69 B 0.02015f
C117 VTAIL.n70 B 0.02015f
C118 VTAIL.n71 B 0.009026f
C119 VTAIL.n72 B 0.008525f
C120 VTAIL.n73 B 0.015864f
C121 VTAIL.n74 B 0.015864f
C122 VTAIL.n75 B 0.008525f
C123 VTAIL.n76 B 0.008525f
C124 VTAIL.n77 B 0.009026f
C125 VTAIL.n78 B 0.02015f
C126 VTAIL.n79 B 0.02015f
C127 VTAIL.n80 B 0.02015f
C128 VTAIL.n81 B 0.008776f
C129 VTAIL.n82 B 0.008525f
C130 VTAIL.n83 B 0.015864f
C131 VTAIL.n84 B 0.015864f
C132 VTAIL.n85 B 0.008525f
C133 VTAIL.n86 B 0.009026f
C134 VTAIL.n87 B 0.02015f
C135 VTAIL.n88 B 0.02015f
C136 VTAIL.n89 B 0.009026f
C137 VTAIL.n90 B 0.008525f
C138 VTAIL.n91 B 0.015864f
C139 VTAIL.n92 B 0.015864f
C140 VTAIL.n93 B 0.008525f
C141 VTAIL.n94 B 0.009026f
C142 VTAIL.n95 B 0.02015f
C143 VTAIL.n96 B 0.045135f
C144 VTAIL.n97 B 0.009026f
C145 VTAIL.n98 B 0.008525f
C146 VTAIL.n99 B 0.038403f
C147 VTAIL.n100 B 0.025462f
C148 VTAIL.n101 B 0.136046f
C149 VTAIL.n102 B 0.023155f
C150 VTAIL.n103 B 0.015864f
C151 VTAIL.n104 B 0.008525f
C152 VTAIL.n105 B 0.02015f
C153 VTAIL.n106 B 0.009026f
C154 VTAIL.n107 B 0.015864f
C155 VTAIL.n108 B 0.008525f
C156 VTAIL.n109 B 0.02015f
C157 VTAIL.n110 B 0.009026f
C158 VTAIL.n111 B 0.015864f
C159 VTAIL.n112 B 0.008776f
C160 VTAIL.n113 B 0.02015f
C161 VTAIL.n114 B 0.009026f
C162 VTAIL.n115 B 0.015864f
C163 VTAIL.n116 B 0.008525f
C164 VTAIL.n117 B 0.02015f
C165 VTAIL.n118 B 0.009026f
C166 VTAIL.n119 B 0.015864f
C167 VTAIL.n120 B 0.008525f
C168 VTAIL.n121 B 0.02015f
C169 VTAIL.n122 B 0.009026f
C170 VTAIL.n123 B 0.015864f
C171 VTAIL.n124 B 0.008525f
C172 VTAIL.n125 B 0.02015f
C173 VTAIL.n126 B 0.009026f
C174 VTAIL.n127 B 0.015864f
C175 VTAIL.n128 B 0.008525f
C176 VTAIL.n129 B 0.02015f
C177 VTAIL.n130 B 0.009026f
C178 VTAIL.n131 B 0.015864f
C179 VTAIL.n132 B 0.008525f
C180 VTAIL.n133 B 0.015112f
C181 VTAIL.n134 B 0.011903f
C182 VTAIL.t1 B 0.033405f
C183 VTAIL.n135 B 0.116676f
C184 VTAIL.n136 B 1.27354f
C185 VTAIL.n137 B 0.008525f
C186 VTAIL.n138 B 0.009026f
C187 VTAIL.n139 B 0.02015f
C188 VTAIL.n140 B 0.02015f
C189 VTAIL.n141 B 0.009026f
C190 VTAIL.n142 B 0.008525f
C191 VTAIL.n143 B 0.015864f
C192 VTAIL.n144 B 0.015864f
C193 VTAIL.n145 B 0.008525f
C194 VTAIL.n146 B 0.009026f
C195 VTAIL.n147 B 0.02015f
C196 VTAIL.n148 B 0.02015f
C197 VTAIL.n149 B 0.009026f
C198 VTAIL.n150 B 0.008525f
C199 VTAIL.n151 B 0.015864f
C200 VTAIL.n152 B 0.015864f
C201 VTAIL.n153 B 0.008525f
C202 VTAIL.n154 B 0.009026f
C203 VTAIL.n155 B 0.02015f
C204 VTAIL.n156 B 0.02015f
C205 VTAIL.n157 B 0.009026f
C206 VTAIL.n158 B 0.008525f
C207 VTAIL.n159 B 0.015864f
C208 VTAIL.n160 B 0.015864f
C209 VTAIL.n161 B 0.008525f
C210 VTAIL.n162 B 0.009026f
C211 VTAIL.n163 B 0.02015f
C212 VTAIL.n164 B 0.02015f
C213 VTAIL.n165 B 0.009026f
C214 VTAIL.n166 B 0.008525f
C215 VTAIL.n167 B 0.015864f
C216 VTAIL.n168 B 0.015864f
C217 VTAIL.n169 B 0.008525f
C218 VTAIL.n170 B 0.009026f
C219 VTAIL.n171 B 0.02015f
C220 VTAIL.n172 B 0.02015f
C221 VTAIL.n173 B 0.009026f
C222 VTAIL.n174 B 0.008525f
C223 VTAIL.n175 B 0.015864f
C224 VTAIL.n176 B 0.015864f
C225 VTAIL.n177 B 0.008525f
C226 VTAIL.n178 B 0.008525f
C227 VTAIL.n179 B 0.009026f
C228 VTAIL.n180 B 0.02015f
C229 VTAIL.n181 B 0.02015f
C230 VTAIL.n182 B 0.02015f
C231 VTAIL.n183 B 0.008776f
C232 VTAIL.n184 B 0.008525f
C233 VTAIL.n185 B 0.015864f
C234 VTAIL.n186 B 0.015864f
C235 VTAIL.n187 B 0.008525f
C236 VTAIL.n188 B 0.009026f
C237 VTAIL.n189 B 0.02015f
C238 VTAIL.n190 B 0.02015f
C239 VTAIL.n191 B 0.009026f
C240 VTAIL.n192 B 0.008525f
C241 VTAIL.n193 B 0.015864f
C242 VTAIL.n194 B 0.015864f
C243 VTAIL.n195 B 0.008525f
C244 VTAIL.n196 B 0.009026f
C245 VTAIL.n197 B 0.02015f
C246 VTAIL.n198 B 0.045135f
C247 VTAIL.n199 B 0.009026f
C248 VTAIL.n200 B 0.008525f
C249 VTAIL.n201 B 0.038403f
C250 VTAIL.n202 B 0.025462f
C251 VTAIL.n203 B 0.227596f
C252 VTAIL.n204 B 0.023155f
C253 VTAIL.n205 B 0.015864f
C254 VTAIL.n206 B 0.008525f
C255 VTAIL.n207 B 0.02015f
C256 VTAIL.n208 B 0.009026f
C257 VTAIL.n209 B 0.015864f
C258 VTAIL.n210 B 0.008525f
C259 VTAIL.n211 B 0.02015f
C260 VTAIL.n212 B 0.009026f
C261 VTAIL.n213 B 0.015864f
C262 VTAIL.n214 B 0.008776f
C263 VTAIL.n215 B 0.02015f
C264 VTAIL.n216 B 0.009026f
C265 VTAIL.n217 B 0.015864f
C266 VTAIL.n218 B 0.008525f
C267 VTAIL.n219 B 0.02015f
C268 VTAIL.n220 B 0.009026f
C269 VTAIL.n221 B 0.015864f
C270 VTAIL.n222 B 0.008525f
C271 VTAIL.n223 B 0.02015f
C272 VTAIL.n224 B 0.009026f
C273 VTAIL.n225 B 0.015864f
C274 VTAIL.n226 B 0.008525f
C275 VTAIL.n227 B 0.02015f
C276 VTAIL.n228 B 0.009026f
C277 VTAIL.n229 B 0.015864f
C278 VTAIL.n230 B 0.008525f
C279 VTAIL.n231 B 0.02015f
C280 VTAIL.n232 B 0.009026f
C281 VTAIL.n233 B 0.015864f
C282 VTAIL.n234 B 0.008525f
C283 VTAIL.n235 B 0.015112f
C284 VTAIL.n236 B 0.011903f
C285 VTAIL.t2 B 0.033405f
C286 VTAIL.n237 B 0.116676f
C287 VTAIL.n238 B 1.27354f
C288 VTAIL.n239 B 0.008525f
C289 VTAIL.n240 B 0.009026f
C290 VTAIL.n241 B 0.02015f
C291 VTAIL.n242 B 0.02015f
C292 VTAIL.n243 B 0.009026f
C293 VTAIL.n244 B 0.008525f
C294 VTAIL.n245 B 0.015864f
C295 VTAIL.n246 B 0.015864f
C296 VTAIL.n247 B 0.008525f
C297 VTAIL.n248 B 0.009026f
C298 VTAIL.n249 B 0.02015f
C299 VTAIL.n250 B 0.02015f
C300 VTAIL.n251 B 0.009026f
C301 VTAIL.n252 B 0.008525f
C302 VTAIL.n253 B 0.015864f
C303 VTAIL.n254 B 0.015864f
C304 VTAIL.n255 B 0.008525f
C305 VTAIL.n256 B 0.009026f
C306 VTAIL.n257 B 0.02015f
C307 VTAIL.n258 B 0.02015f
C308 VTAIL.n259 B 0.009026f
C309 VTAIL.n260 B 0.008525f
C310 VTAIL.n261 B 0.015864f
C311 VTAIL.n262 B 0.015864f
C312 VTAIL.n263 B 0.008525f
C313 VTAIL.n264 B 0.009026f
C314 VTAIL.n265 B 0.02015f
C315 VTAIL.n266 B 0.02015f
C316 VTAIL.n267 B 0.009026f
C317 VTAIL.n268 B 0.008525f
C318 VTAIL.n269 B 0.015864f
C319 VTAIL.n270 B 0.015864f
C320 VTAIL.n271 B 0.008525f
C321 VTAIL.n272 B 0.009026f
C322 VTAIL.n273 B 0.02015f
C323 VTAIL.n274 B 0.02015f
C324 VTAIL.n275 B 0.009026f
C325 VTAIL.n276 B 0.008525f
C326 VTAIL.n277 B 0.015864f
C327 VTAIL.n278 B 0.015864f
C328 VTAIL.n279 B 0.008525f
C329 VTAIL.n280 B 0.008525f
C330 VTAIL.n281 B 0.009026f
C331 VTAIL.n282 B 0.02015f
C332 VTAIL.n283 B 0.02015f
C333 VTAIL.n284 B 0.02015f
C334 VTAIL.n285 B 0.008776f
C335 VTAIL.n286 B 0.008525f
C336 VTAIL.n287 B 0.015864f
C337 VTAIL.n288 B 0.015864f
C338 VTAIL.n289 B 0.008525f
C339 VTAIL.n290 B 0.009026f
C340 VTAIL.n291 B 0.02015f
C341 VTAIL.n292 B 0.02015f
C342 VTAIL.n293 B 0.009026f
C343 VTAIL.n294 B 0.008525f
C344 VTAIL.n295 B 0.015864f
C345 VTAIL.n296 B 0.015864f
C346 VTAIL.n297 B 0.008525f
C347 VTAIL.n298 B 0.009026f
C348 VTAIL.n299 B 0.02015f
C349 VTAIL.n300 B 0.045135f
C350 VTAIL.n301 B 0.009026f
C351 VTAIL.n302 B 0.008525f
C352 VTAIL.n303 B 0.038403f
C353 VTAIL.n304 B 0.025462f
C354 VTAIL.n305 B 1.41545f
C355 VTAIL.n306 B 0.023155f
C356 VTAIL.n307 B 0.015864f
C357 VTAIL.n308 B 0.008525f
C358 VTAIL.n309 B 0.02015f
C359 VTAIL.n310 B 0.009026f
C360 VTAIL.n311 B 0.015864f
C361 VTAIL.n312 B 0.008525f
C362 VTAIL.n313 B 0.02015f
C363 VTAIL.n314 B 0.009026f
C364 VTAIL.n315 B 0.015864f
C365 VTAIL.n316 B 0.008776f
C366 VTAIL.n317 B 0.02015f
C367 VTAIL.n318 B 0.008525f
C368 VTAIL.n319 B 0.009026f
C369 VTAIL.n320 B 0.015864f
C370 VTAIL.n321 B 0.008525f
C371 VTAIL.n322 B 0.02015f
C372 VTAIL.n323 B 0.009026f
C373 VTAIL.n324 B 0.015864f
C374 VTAIL.n325 B 0.008525f
C375 VTAIL.n326 B 0.02015f
C376 VTAIL.n327 B 0.009026f
C377 VTAIL.n328 B 0.015864f
C378 VTAIL.n329 B 0.008525f
C379 VTAIL.n330 B 0.02015f
C380 VTAIL.n331 B 0.009026f
C381 VTAIL.n332 B 0.015864f
C382 VTAIL.n333 B 0.008525f
C383 VTAIL.n334 B 0.02015f
C384 VTAIL.n335 B 0.009026f
C385 VTAIL.n336 B 0.015864f
C386 VTAIL.n337 B 0.008525f
C387 VTAIL.n338 B 0.015112f
C388 VTAIL.n339 B 0.011903f
C389 VTAIL.t4 B 0.033405f
C390 VTAIL.n340 B 0.116676f
C391 VTAIL.n341 B 1.27354f
C392 VTAIL.n342 B 0.008525f
C393 VTAIL.n343 B 0.009026f
C394 VTAIL.n344 B 0.02015f
C395 VTAIL.n345 B 0.02015f
C396 VTAIL.n346 B 0.009026f
C397 VTAIL.n347 B 0.008525f
C398 VTAIL.n348 B 0.015864f
C399 VTAIL.n349 B 0.015864f
C400 VTAIL.n350 B 0.008525f
C401 VTAIL.n351 B 0.009026f
C402 VTAIL.n352 B 0.02015f
C403 VTAIL.n353 B 0.02015f
C404 VTAIL.n354 B 0.009026f
C405 VTAIL.n355 B 0.008525f
C406 VTAIL.n356 B 0.015864f
C407 VTAIL.n357 B 0.015864f
C408 VTAIL.n358 B 0.008525f
C409 VTAIL.n359 B 0.009026f
C410 VTAIL.n360 B 0.02015f
C411 VTAIL.n361 B 0.02015f
C412 VTAIL.n362 B 0.009026f
C413 VTAIL.n363 B 0.008525f
C414 VTAIL.n364 B 0.015864f
C415 VTAIL.n365 B 0.015864f
C416 VTAIL.n366 B 0.008525f
C417 VTAIL.n367 B 0.009026f
C418 VTAIL.n368 B 0.02015f
C419 VTAIL.n369 B 0.02015f
C420 VTAIL.n370 B 0.009026f
C421 VTAIL.n371 B 0.008525f
C422 VTAIL.n372 B 0.015864f
C423 VTAIL.n373 B 0.015864f
C424 VTAIL.n374 B 0.008525f
C425 VTAIL.n375 B 0.009026f
C426 VTAIL.n376 B 0.02015f
C427 VTAIL.n377 B 0.02015f
C428 VTAIL.n378 B 0.009026f
C429 VTAIL.n379 B 0.008525f
C430 VTAIL.n380 B 0.015864f
C431 VTAIL.n381 B 0.015864f
C432 VTAIL.n382 B 0.008525f
C433 VTAIL.n383 B 0.009026f
C434 VTAIL.n384 B 0.02015f
C435 VTAIL.n385 B 0.02015f
C436 VTAIL.n386 B 0.02015f
C437 VTAIL.n387 B 0.008776f
C438 VTAIL.n388 B 0.008525f
C439 VTAIL.n389 B 0.015864f
C440 VTAIL.n390 B 0.015864f
C441 VTAIL.n391 B 0.008525f
C442 VTAIL.n392 B 0.009026f
C443 VTAIL.n393 B 0.02015f
C444 VTAIL.n394 B 0.02015f
C445 VTAIL.n395 B 0.009026f
C446 VTAIL.n396 B 0.008525f
C447 VTAIL.n397 B 0.015864f
C448 VTAIL.n398 B 0.015864f
C449 VTAIL.n399 B 0.008525f
C450 VTAIL.n400 B 0.009026f
C451 VTAIL.n401 B 0.02015f
C452 VTAIL.n402 B 0.045135f
C453 VTAIL.n403 B 0.009026f
C454 VTAIL.n404 B 0.008525f
C455 VTAIL.n405 B 0.038403f
C456 VTAIL.n406 B 0.025462f
C457 VTAIL.n407 B 1.41545f
C458 VTAIL.n408 B 0.023155f
C459 VTAIL.n409 B 0.015864f
C460 VTAIL.n410 B 0.008525f
C461 VTAIL.n411 B 0.02015f
C462 VTAIL.n412 B 0.009026f
C463 VTAIL.n413 B 0.015864f
C464 VTAIL.n414 B 0.008525f
C465 VTAIL.n415 B 0.02015f
C466 VTAIL.n416 B 0.009026f
C467 VTAIL.n417 B 0.015864f
C468 VTAIL.n418 B 0.008776f
C469 VTAIL.n419 B 0.02015f
C470 VTAIL.n420 B 0.008525f
C471 VTAIL.n421 B 0.009026f
C472 VTAIL.n422 B 0.015864f
C473 VTAIL.n423 B 0.008525f
C474 VTAIL.n424 B 0.02015f
C475 VTAIL.n425 B 0.009026f
C476 VTAIL.n426 B 0.015864f
C477 VTAIL.n427 B 0.008525f
C478 VTAIL.n428 B 0.02015f
C479 VTAIL.n429 B 0.009026f
C480 VTAIL.n430 B 0.015864f
C481 VTAIL.n431 B 0.008525f
C482 VTAIL.n432 B 0.02015f
C483 VTAIL.n433 B 0.009026f
C484 VTAIL.n434 B 0.015864f
C485 VTAIL.n435 B 0.008525f
C486 VTAIL.n436 B 0.02015f
C487 VTAIL.n437 B 0.009026f
C488 VTAIL.n438 B 0.015864f
C489 VTAIL.n439 B 0.008525f
C490 VTAIL.n440 B 0.015112f
C491 VTAIL.n441 B 0.011903f
C492 VTAIL.t5 B 0.033405f
C493 VTAIL.n442 B 0.116676f
C494 VTAIL.n443 B 1.27354f
C495 VTAIL.n444 B 0.008525f
C496 VTAIL.n445 B 0.009026f
C497 VTAIL.n446 B 0.02015f
C498 VTAIL.n447 B 0.02015f
C499 VTAIL.n448 B 0.009026f
C500 VTAIL.n449 B 0.008525f
C501 VTAIL.n450 B 0.015864f
C502 VTAIL.n451 B 0.015864f
C503 VTAIL.n452 B 0.008525f
C504 VTAIL.n453 B 0.009026f
C505 VTAIL.n454 B 0.02015f
C506 VTAIL.n455 B 0.02015f
C507 VTAIL.n456 B 0.009026f
C508 VTAIL.n457 B 0.008525f
C509 VTAIL.n458 B 0.015864f
C510 VTAIL.n459 B 0.015864f
C511 VTAIL.n460 B 0.008525f
C512 VTAIL.n461 B 0.009026f
C513 VTAIL.n462 B 0.02015f
C514 VTAIL.n463 B 0.02015f
C515 VTAIL.n464 B 0.009026f
C516 VTAIL.n465 B 0.008525f
C517 VTAIL.n466 B 0.015864f
C518 VTAIL.n467 B 0.015864f
C519 VTAIL.n468 B 0.008525f
C520 VTAIL.n469 B 0.009026f
C521 VTAIL.n470 B 0.02015f
C522 VTAIL.n471 B 0.02015f
C523 VTAIL.n472 B 0.009026f
C524 VTAIL.n473 B 0.008525f
C525 VTAIL.n474 B 0.015864f
C526 VTAIL.n475 B 0.015864f
C527 VTAIL.n476 B 0.008525f
C528 VTAIL.n477 B 0.009026f
C529 VTAIL.n478 B 0.02015f
C530 VTAIL.n479 B 0.02015f
C531 VTAIL.n480 B 0.009026f
C532 VTAIL.n481 B 0.008525f
C533 VTAIL.n482 B 0.015864f
C534 VTAIL.n483 B 0.015864f
C535 VTAIL.n484 B 0.008525f
C536 VTAIL.n485 B 0.009026f
C537 VTAIL.n486 B 0.02015f
C538 VTAIL.n487 B 0.02015f
C539 VTAIL.n488 B 0.02015f
C540 VTAIL.n489 B 0.008776f
C541 VTAIL.n490 B 0.008525f
C542 VTAIL.n491 B 0.015864f
C543 VTAIL.n492 B 0.015864f
C544 VTAIL.n493 B 0.008525f
C545 VTAIL.n494 B 0.009026f
C546 VTAIL.n495 B 0.02015f
C547 VTAIL.n496 B 0.02015f
C548 VTAIL.n497 B 0.009026f
C549 VTAIL.n498 B 0.008525f
C550 VTAIL.n499 B 0.015864f
C551 VTAIL.n500 B 0.015864f
C552 VTAIL.n501 B 0.008525f
C553 VTAIL.n502 B 0.009026f
C554 VTAIL.n503 B 0.02015f
C555 VTAIL.n504 B 0.045135f
C556 VTAIL.n505 B 0.009026f
C557 VTAIL.n506 B 0.008525f
C558 VTAIL.n507 B 0.038403f
C559 VTAIL.n508 B 0.025462f
C560 VTAIL.n509 B 0.227596f
C561 VTAIL.n510 B 0.023155f
C562 VTAIL.n511 B 0.015864f
C563 VTAIL.n512 B 0.008525f
C564 VTAIL.n513 B 0.02015f
C565 VTAIL.n514 B 0.009026f
C566 VTAIL.n515 B 0.015864f
C567 VTAIL.n516 B 0.008525f
C568 VTAIL.n517 B 0.02015f
C569 VTAIL.n518 B 0.009026f
C570 VTAIL.n519 B 0.015864f
C571 VTAIL.n520 B 0.008776f
C572 VTAIL.n521 B 0.02015f
C573 VTAIL.n522 B 0.008525f
C574 VTAIL.n523 B 0.009026f
C575 VTAIL.n524 B 0.015864f
C576 VTAIL.n525 B 0.008525f
C577 VTAIL.n526 B 0.02015f
C578 VTAIL.n527 B 0.009026f
C579 VTAIL.n528 B 0.015864f
C580 VTAIL.n529 B 0.008525f
C581 VTAIL.n530 B 0.02015f
C582 VTAIL.n531 B 0.009026f
C583 VTAIL.n532 B 0.015864f
C584 VTAIL.n533 B 0.008525f
C585 VTAIL.n534 B 0.02015f
C586 VTAIL.n535 B 0.009026f
C587 VTAIL.n536 B 0.015864f
C588 VTAIL.n537 B 0.008525f
C589 VTAIL.n538 B 0.02015f
C590 VTAIL.n539 B 0.009026f
C591 VTAIL.n540 B 0.015864f
C592 VTAIL.n541 B 0.008525f
C593 VTAIL.n542 B 0.015112f
C594 VTAIL.n543 B 0.011903f
C595 VTAIL.t0 B 0.033405f
C596 VTAIL.n544 B 0.116676f
C597 VTAIL.n545 B 1.27354f
C598 VTAIL.n546 B 0.008525f
C599 VTAIL.n547 B 0.009026f
C600 VTAIL.n548 B 0.02015f
C601 VTAIL.n549 B 0.02015f
C602 VTAIL.n550 B 0.009026f
C603 VTAIL.n551 B 0.008525f
C604 VTAIL.n552 B 0.015864f
C605 VTAIL.n553 B 0.015864f
C606 VTAIL.n554 B 0.008525f
C607 VTAIL.n555 B 0.009026f
C608 VTAIL.n556 B 0.02015f
C609 VTAIL.n557 B 0.02015f
C610 VTAIL.n558 B 0.009026f
C611 VTAIL.n559 B 0.008525f
C612 VTAIL.n560 B 0.015864f
C613 VTAIL.n561 B 0.015864f
C614 VTAIL.n562 B 0.008525f
C615 VTAIL.n563 B 0.009026f
C616 VTAIL.n564 B 0.02015f
C617 VTAIL.n565 B 0.02015f
C618 VTAIL.n566 B 0.009026f
C619 VTAIL.n567 B 0.008525f
C620 VTAIL.n568 B 0.015864f
C621 VTAIL.n569 B 0.015864f
C622 VTAIL.n570 B 0.008525f
C623 VTAIL.n571 B 0.009026f
C624 VTAIL.n572 B 0.02015f
C625 VTAIL.n573 B 0.02015f
C626 VTAIL.n574 B 0.009026f
C627 VTAIL.n575 B 0.008525f
C628 VTAIL.n576 B 0.015864f
C629 VTAIL.n577 B 0.015864f
C630 VTAIL.n578 B 0.008525f
C631 VTAIL.n579 B 0.009026f
C632 VTAIL.n580 B 0.02015f
C633 VTAIL.n581 B 0.02015f
C634 VTAIL.n582 B 0.009026f
C635 VTAIL.n583 B 0.008525f
C636 VTAIL.n584 B 0.015864f
C637 VTAIL.n585 B 0.015864f
C638 VTAIL.n586 B 0.008525f
C639 VTAIL.n587 B 0.009026f
C640 VTAIL.n588 B 0.02015f
C641 VTAIL.n589 B 0.02015f
C642 VTAIL.n590 B 0.02015f
C643 VTAIL.n591 B 0.008776f
C644 VTAIL.n592 B 0.008525f
C645 VTAIL.n593 B 0.015864f
C646 VTAIL.n594 B 0.015864f
C647 VTAIL.n595 B 0.008525f
C648 VTAIL.n596 B 0.009026f
C649 VTAIL.n597 B 0.02015f
C650 VTAIL.n598 B 0.02015f
C651 VTAIL.n599 B 0.009026f
C652 VTAIL.n600 B 0.008525f
C653 VTAIL.n601 B 0.015864f
C654 VTAIL.n602 B 0.015864f
C655 VTAIL.n603 B 0.008525f
C656 VTAIL.n604 B 0.009026f
C657 VTAIL.n605 B 0.02015f
C658 VTAIL.n606 B 0.045135f
C659 VTAIL.n607 B 0.009026f
C660 VTAIL.n608 B 0.008525f
C661 VTAIL.n609 B 0.038403f
C662 VTAIL.n610 B 0.025462f
C663 VTAIL.n611 B 0.227596f
C664 VTAIL.n612 B 0.023155f
C665 VTAIL.n613 B 0.015864f
C666 VTAIL.n614 B 0.008525f
C667 VTAIL.n615 B 0.02015f
C668 VTAIL.n616 B 0.009026f
C669 VTAIL.n617 B 0.015864f
C670 VTAIL.n618 B 0.008525f
C671 VTAIL.n619 B 0.02015f
C672 VTAIL.n620 B 0.009026f
C673 VTAIL.n621 B 0.015864f
C674 VTAIL.n622 B 0.008776f
C675 VTAIL.n623 B 0.02015f
C676 VTAIL.n624 B 0.008525f
C677 VTAIL.n625 B 0.009026f
C678 VTAIL.n626 B 0.015864f
C679 VTAIL.n627 B 0.008525f
C680 VTAIL.n628 B 0.02015f
C681 VTAIL.n629 B 0.009026f
C682 VTAIL.n630 B 0.015864f
C683 VTAIL.n631 B 0.008525f
C684 VTAIL.n632 B 0.02015f
C685 VTAIL.n633 B 0.009026f
C686 VTAIL.n634 B 0.015864f
C687 VTAIL.n635 B 0.008525f
C688 VTAIL.n636 B 0.02015f
C689 VTAIL.n637 B 0.009026f
C690 VTAIL.n638 B 0.015864f
C691 VTAIL.n639 B 0.008525f
C692 VTAIL.n640 B 0.02015f
C693 VTAIL.n641 B 0.009026f
C694 VTAIL.n642 B 0.015864f
C695 VTAIL.n643 B 0.008525f
C696 VTAIL.n644 B 0.015112f
C697 VTAIL.n645 B 0.011903f
C698 VTAIL.t3 B 0.033405f
C699 VTAIL.n646 B 0.116676f
C700 VTAIL.n647 B 1.27354f
C701 VTAIL.n648 B 0.008525f
C702 VTAIL.n649 B 0.009026f
C703 VTAIL.n650 B 0.02015f
C704 VTAIL.n651 B 0.02015f
C705 VTAIL.n652 B 0.009026f
C706 VTAIL.n653 B 0.008525f
C707 VTAIL.n654 B 0.015864f
C708 VTAIL.n655 B 0.015864f
C709 VTAIL.n656 B 0.008525f
C710 VTAIL.n657 B 0.009026f
C711 VTAIL.n658 B 0.02015f
C712 VTAIL.n659 B 0.02015f
C713 VTAIL.n660 B 0.009026f
C714 VTAIL.n661 B 0.008525f
C715 VTAIL.n662 B 0.015864f
C716 VTAIL.n663 B 0.015864f
C717 VTAIL.n664 B 0.008525f
C718 VTAIL.n665 B 0.009026f
C719 VTAIL.n666 B 0.02015f
C720 VTAIL.n667 B 0.02015f
C721 VTAIL.n668 B 0.009026f
C722 VTAIL.n669 B 0.008525f
C723 VTAIL.n670 B 0.015864f
C724 VTAIL.n671 B 0.015864f
C725 VTAIL.n672 B 0.008525f
C726 VTAIL.n673 B 0.009026f
C727 VTAIL.n674 B 0.02015f
C728 VTAIL.n675 B 0.02015f
C729 VTAIL.n676 B 0.009026f
C730 VTAIL.n677 B 0.008525f
C731 VTAIL.n678 B 0.015864f
C732 VTAIL.n679 B 0.015864f
C733 VTAIL.n680 B 0.008525f
C734 VTAIL.n681 B 0.009026f
C735 VTAIL.n682 B 0.02015f
C736 VTAIL.n683 B 0.02015f
C737 VTAIL.n684 B 0.009026f
C738 VTAIL.n685 B 0.008525f
C739 VTAIL.n686 B 0.015864f
C740 VTAIL.n687 B 0.015864f
C741 VTAIL.n688 B 0.008525f
C742 VTAIL.n689 B 0.009026f
C743 VTAIL.n690 B 0.02015f
C744 VTAIL.n691 B 0.02015f
C745 VTAIL.n692 B 0.02015f
C746 VTAIL.n693 B 0.008776f
C747 VTAIL.n694 B 0.008525f
C748 VTAIL.n695 B 0.015864f
C749 VTAIL.n696 B 0.015864f
C750 VTAIL.n697 B 0.008525f
C751 VTAIL.n698 B 0.009026f
C752 VTAIL.n699 B 0.02015f
C753 VTAIL.n700 B 0.02015f
C754 VTAIL.n701 B 0.009026f
C755 VTAIL.n702 B 0.008525f
C756 VTAIL.n703 B 0.015864f
C757 VTAIL.n704 B 0.015864f
C758 VTAIL.n705 B 0.008525f
C759 VTAIL.n706 B 0.009026f
C760 VTAIL.n707 B 0.02015f
C761 VTAIL.n708 B 0.045135f
C762 VTAIL.n709 B 0.009026f
C763 VTAIL.n710 B 0.008525f
C764 VTAIL.n711 B 0.038403f
C765 VTAIL.n712 B 0.025462f
C766 VTAIL.n713 B 1.41545f
C767 VTAIL.n714 B 0.023155f
C768 VTAIL.n715 B 0.015864f
C769 VTAIL.n716 B 0.008525f
C770 VTAIL.n717 B 0.02015f
C771 VTAIL.n718 B 0.009026f
C772 VTAIL.n719 B 0.015864f
C773 VTAIL.n720 B 0.008525f
C774 VTAIL.n721 B 0.02015f
C775 VTAIL.n722 B 0.009026f
C776 VTAIL.n723 B 0.015864f
C777 VTAIL.n724 B 0.008776f
C778 VTAIL.n725 B 0.02015f
C779 VTAIL.n726 B 0.009026f
C780 VTAIL.n727 B 0.015864f
C781 VTAIL.n728 B 0.008525f
C782 VTAIL.n729 B 0.02015f
C783 VTAIL.n730 B 0.009026f
C784 VTAIL.n731 B 0.015864f
C785 VTAIL.n732 B 0.008525f
C786 VTAIL.n733 B 0.02015f
C787 VTAIL.n734 B 0.009026f
C788 VTAIL.n735 B 0.015864f
C789 VTAIL.n736 B 0.008525f
C790 VTAIL.n737 B 0.02015f
C791 VTAIL.n738 B 0.009026f
C792 VTAIL.n739 B 0.015864f
C793 VTAIL.n740 B 0.008525f
C794 VTAIL.n741 B 0.02015f
C795 VTAIL.n742 B 0.009026f
C796 VTAIL.n743 B 0.015864f
C797 VTAIL.n744 B 0.008525f
C798 VTAIL.n745 B 0.015112f
C799 VTAIL.n746 B 0.011903f
C800 VTAIL.t6 B 0.033405f
C801 VTAIL.n747 B 0.116676f
C802 VTAIL.n748 B 1.27354f
C803 VTAIL.n749 B 0.008525f
C804 VTAIL.n750 B 0.009026f
C805 VTAIL.n751 B 0.02015f
C806 VTAIL.n752 B 0.02015f
C807 VTAIL.n753 B 0.009026f
C808 VTAIL.n754 B 0.008525f
C809 VTAIL.n755 B 0.015864f
C810 VTAIL.n756 B 0.015864f
C811 VTAIL.n757 B 0.008525f
C812 VTAIL.n758 B 0.009026f
C813 VTAIL.n759 B 0.02015f
C814 VTAIL.n760 B 0.02015f
C815 VTAIL.n761 B 0.009026f
C816 VTAIL.n762 B 0.008525f
C817 VTAIL.n763 B 0.015864f
C818 VTAIL.n764 B 0.015864f
C819 VTAIL.n765 B 0.008525f
C820 VTAIL.n766 B 0.009026f
C821 VTAIL.n767 B 0.02015f
C822 VTAIL.n768 B 0.02015f
C823 VTAIL.n769 B 0.009026f
C824 VTAIL.n770 B 0.008525f
C825 VTAIL.n771 B 0.015864f
C826 VTAIL.n772 B 0.015864f
C827 VTAIL.n773 B 0.008525f
C828 VTAIL.n774 B 0.009026f
C829 VTAIL.n775 B 0.02015f
C830 VTAIL.n776 B 0.02015f
C831 VTAIL.n777 B 0.009026f
C832 VTAIL.n778 B 0.008525f
C833 VTAIL.n779 B 0.015864f
C834 VTAIL.n780 B 0.015864f
C835 VTAIL.n781 B 0.008525f
C836 VTAIL.n782 B 0.009026f
C837 VTAIL.n783 B 0.02015f
C838 VTAIL.n784 B 0.02015f
C839 VTAIL.n785 B 0.009026f
C840 VTAIL.n786 B 0.008525f
C841 VTAIL.n787 B 0.015864f
C842 VTAIL.n788 B 0.015864f
C843 VTAIL.n789 B 0.008525f
C844 VTAIL.n790 B 0.008525f
C845 VTAIL.n791 B 0.009026f
C846 VTAIL.n792 B 0.02015f
C847 VTAIL.n793 B 0.02015f
C848 VTAIL.n794 B 0.02015f
C849 VTAIL.n795 B 0.008776f
C850 VTAIL.n796 B 0.008525f
C851 VTAIL.n797 B 0.015864f
C852 VTAIL.n798 B 0.015864f
C853 VTAIL.n799 B 0.008525f
C854 VTAIL.n800 B 0.009026f
C855 VTAIL.n801 B 0.02015f
C856 VTAIL.n802 B 0.02015f
C857 VTAIL.n803 B 0.009026f
C858 VTAIL.n804 B 0.008525f
C859 VTAIL.n805 B 0.015864f
C860 VTAIL.n806 B 0.015864f
C861 VTAIL.n807 B 0.008525f
C862 VTAIL.n808 B 0.009026f
C863 VTAIL.n809 B 0.02015f
C864 VTAIL.n810 B 0.045135f
C865 VTAIL.n811 B 0.009026f
C866 VTAIL.n812 B 0.008525f
C867 VTAIL.n813 B 0.038403f
C868 VTAIL.n814 B 0.025462f
C869 VTAIL.n815 B 1.31795f
C870 VDD2.t2 B 0.387271f
C871 VDD2.t3 B 0.387271f
C872 VDD2.n0 B 4.51512f
C873 VDD2.t1 B 0.387271f
C874 VDD2.t0 B 0.387271f
C875 VDD2.n1 B 3.53218f
C876 VDD2.n2 B 4.77908f
C877 VN.t0 B 3.92219f
C878 VN.t1 B 3.90909f
C879 VN.n0 B 2.37364f
C880 VN.t2 B 3.92219f
C881 VN.t3 B 3.90909f
C882 VN.n1 B 3.72028f
.ends

