* NGSPICE file created from diff_pair_sample_1786.ext - technology: sky130A

.subckt diff_pair_sample_1786 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X1 VDD1.t6 VP.t1 VTAIL.t11 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=6.2049 ps=32.6 w=15.91 l=3.32
X2 VDD2.t7 VN.t0 VTAIL.t4 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X3 VTAIL.t5 VN.t1 VDD2.t6 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X4 VTAIL.t10 VP.t2 VDD1.t5 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X5 B.t11 B.t9 B.t10 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=0 ps=0 w=15.91 l=3.32
X6 VDD2.t5 VN.t2 VTAIL.t6 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=6.2049 ps=32.6 w=15.91 l=3.32
X7 VTAIL.t12 VP.t3 VDD1.t4 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=2.62515 ps=16.24 w=15.91 l=3.32
X8 B.t8 B.t6 B.t7 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=0 ps=0 w=15.91 l=3.32
X9 VDD1.t3 VP.t4 VTAIL.t15 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=6.2049 ps=32.6 w=15.91 l=3.32
X10 VTAIL.t7 VN.t3 VDD2.t4 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X11 VDD2.t3 VN.t4 VTAIL.t3 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X12 B.t5 B.t3 B.t4 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=0 ps=0 w=15.91 l=3.32
X13 VDD2.t2 VN.t5 VTAIL.t2 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=6.2049 ps=32.6 w=15.91 l=3.32
X14 VTAIL.t13 VP.t5 VDD1.t2 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X15 VTAIL.t8 VP.t6 VDD1.t1 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=2.62515 ps=16.24 w=15.91 l=3.32
X16 VTAIL.t1 VN.t6 VDD2.t1 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=2.62515 ps=16.24 w=15.91 l=3.32
X17 VDD1.t0 VP.t7 VTAIL.t9 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=2.62515 pd=16.24 as=2.62515 ps=16.24 w=15.91 l=3.32
X18 B.t2 B.t0 B.t1 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=0 ps=0 w=15.91 l=3.32
X19 VTAIL.t0 VN.t7 VDD2.t0 w_n4620_n4150# sky130_fd_pr__pfet_01v8 ad=6.2049 pd=32.6 as=2.62515 ps=16.24 w=15.91 l=3.32
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n23 VP.t6 147.798
R38 VP.n12 VP.t3 115.492
R39 VP.n58 VP.t7 115.492
R40 VP.n4 VP.t2 115.492
R41 VP.n0 VP.t4 115.492
R42 VP.n13 VP.t1 115.492
R43 VP.n17 VP.t5 115.492
R44 VP.n22 VP.t0 115.492
R45 VP.n48 VP.n12 79.0572
R46 VP.n84 VP.n0 79.0572
R47 VP.n47 VP.n13 79.0572
R48 VP.n23 VP.n22 70.9133
R49 VP.n48 VP.n47 57.2872
R50 VP.n65 VP.n6 56.5193
R51 VP.n28 VP.n19 56.5193
R52 VP.n56 VP.n10 50.2061
R53 VP.n76 VP.n2 50.2061
R54 VP.n39 VP.n15 50.2061
R55 VP.n52 VP.n10 30.7807
R56 VP.n80 VP.n2 30.7807
R57 VP.n43 VP.n15 30.7807
R58 VP.n51 VP.n50 24.4675
R59 VP.n52 VP.n51 24.4675
R60 VP.n57 VP.n56 24.4675
R61 VP.n59 VP.n57 24.4675
R62 VP.n63 VP.n8 24.4675
R63 VP.n64 VP.n63 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n69 VP.n6 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n71 VP.n70 24.4675
R68 VP.n75 VP.n74 24.4675
R69 VP.n76 VP.n75 24.4675
R70 VP.n81 VP.n80 24.4675
R71 VP.n82 VP.n81 24.4675
R72 VP.n44 VP.n43 24.4675
R73 VP.n45 VP.n44 24.4675
R74 VP.n32 VP.n19 24.4675
R75 VP.n33 VP.n32 24.4675
R76 VP.n34 VP.n33 24.4675
R77 VP.n38 VP.n37 24.4675
R78 VP.n39 VP.n38 24.4675
R79 VP.n26 VP.n21 24.4675
R80 VP.n27 VP.n26 24.4675
R81 VP.n28 VP.n27 24.4675
R82 VP.n59 VP.n58 20.7975
R83 VP.n74 VP.n4 20.7975
R84 VP.n37 VP.n17 20.7975
R85 VP.n50 VP.n12 11.0107
R86 VP.n82 VP.n0 11.0107
R87 VP.n45 VP.n13 11.0107
R88 VP.n24 VP.n23 4.35326
R89 VP.n58 VP.n8 3.67055
R90 VP.n71 VP.n4 3.67055
R91 VP.n34 VP.n17 3.67055
R92 VP.n22 VP.n21 3.67055
R93 VP.n47 VP.n46 0.354971
R94 VP.n49 VP.n48 0.354971
R95 VP.n84 VP.n83 0.354971
R96 VP VP.n84 0.26696
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VTAIL.n11 VTAIL.t8 59.0728
R133 VTAIL.n10 VTAIL.t6 59.0728
R134 VTAIL.n7 VTAIL.t1 59.0728
R135 VTAIL.n15 VTAIL.t2 59.0727
R136 VTAIL.n2 VTAIL.t0 59.0727
R137 VTAIL.n3 VTAIL.t15 59.0727
R138 VTAIL.n6 VTAIL.t12 59.0727
R139 VTAIL.n14 VTAIL.t11 59.0727
R140 VTAIL.n13 VTAIL.n12 57.0298
R141 VTAIL.n9 VTAIL.n8 57.0298
R142 VTAIL.n1 VTAIL.n0 57.0296
R143 VTAIL.n5 VTAIL.n4 57.0296
R144 VTAIL.n15 VTAIL.n14 29.2289
R145 VTAIL.n7 VTAIL.n6 29.2289
R146 VTAIL.n9 VTAIL.n7 3.14705
R147 VTAIL.n10 VTAIL.n9 3.14705
R148 VTAIL.n13 VTAIL.n11 3.14705
R149 VTAIL.n14 VTAIL.n13 3.14705
R150 VTAIL.n6 VTAIL.n5 3.14705
R151 VTAIL.n5 VTAIL.n3 3.14705
R152 VTAIL.n2 VTAIL.n1 3.14705
R153 VTAIL VTAIL.n15 3.08886
R154 VTAIL.n0 VTAIL.t3 2.04355
R155 VTAIL.n0 VTAIL.t5 2.04355
R156 VTAIL.n4 VTAIL.t9 2.04355
R157 VTAIL.n4 VTAIL.t10 2.04355
R158 VTAIL.n12 VTAIL.t14 2.04355
R159 VTAIL.n12 VTAIL.t13 2.04355
R160 VTAIL.n8 VTAIL.t4 2.04355
R161 VTAIL.n8 VTAIL.t7 2.04355
R162 VTAIL.n11 VTAIL.n10 0.470328
R163 VTAIL.n3 VTAIL.n2 0.470328
R164 VTAIL VTAIL.n1 0.0586897
R165 VDD1 VDD1.n0 75.3401
R166 VDD1.n3 VDD1.n2 75.2263
R167 VDD1.n3 VDD1.n1 75.2263
R168 VDD1.n5 VDD1.n4 73.7084
R169 VDD1.n5 VDD1.n3 52.1733
R170 VDD1.n4 VDD1.t2 2.04355
R171 VDD1.n4 VDD1.t6 2.04355
R172 VDD1.n0 VDD1.t1 2.04355
R173 VDD1.n0 VDD1.t7 2.04355
R174 VDD1.n2 VDD1.t5 2.04355
R175 VDD1.n2 VDD1.t3 2.04355
R176 VDD1.n1 VDD1.t4 2.04355
R177 VDD1.n1 VDD1.t0 2.04355
R178 VDD1 VDD1.n5 1.51559
R179 VN.n68 VN.n67 161.3
R180 VN.n66 VN.n36 161.3
R181 VN.n65 VN.n64 161.3
R182 VN.n63 VN.n37 161.3
R183 VN.n62 VN.n61 161.3
R184 VN.n60 VN.n38 161.3
R185 VN.n59 VN.n58 161.3
R186 VN.n57 VN.n56 161.3
R187 VN.n55 VN.n40 161.3
R188 VN.n54 VN.n53 161.3
R189 VN.n52 VN.n41 161.3
R190 VN.n51 VN.n50 161.3
R191 VN.n49 VN.n42 161.3
R192 VN.n48 VN.n47 161.3
R193 VN.n46 VN.n43 161.3
R194 VN.n33 VN.n32 161.3
R195 VN.n31 VN.n1 161.3
R196 VN.n30 VN.n29 161.3
R197 VN.n28 VN.n2 161.3
R198 VN.n27 VN.n26 161.3
R199 VN.n25 VN.n3 161.3
R200 VN.n24 VN.n23 161.3
R201 VN.n22 VN.n21 161.3
R202 VN.n20 VN.n5 161.3
R203 VN.n19 VN.n18 161.3
R204 VN.n17 VN.n6 161.3
R205 VN.n16 VN.n15 161.3
R206 VN.n14 VN.n7 161.3
R207 VN.n13 VN.n12 161.3
R208 VN.n11 VN.n8 161.3
R209 VN.n45 VN.t2 147.798
R210 VN.n10 VN.t7 147.798
R211 VN.n9 VN.t4 115.492
R212 VN.n4 VN.t1 115.492
R213 VN.n0 VN.t5 115.492
R214 VN.n44 VN.t3 115.492
R215 VN.n39 VN.t0 115.492
R216 VN.n35 VN.t6 115.492
R217 VN.n34 VN.n0 79.0572
R218 VN.n69 VN.n35 79.0572
R219 VN.n45 VN.n44 70.9133
R220 VN.n10 VN.n9 70.9133
R221 VN VN.n69 57.4526
R222 VN.n15 VN.n6 56.5193
R223 VN.n50 VN.n41 56.5193
R224 VN.n26 VN.n2 50.2061
R225 VN.n61 VN.n37 50.2061
R226 VN.n30 VN.n2 30.7807
R227 VN.n65 VN.n37 30.7807
R228 VN.n13 VN.n8 24.4675
R229 VN.n14 VN.n13 24.4675
R230 VN.n15 VN.n14 24.4675
R231 VN.n19 VN.n6 24.4675
R232 VN.n20 VN.n19 24.4675
R233 VN.n21 VN.n20 24.4675
R234 VN.n25 VN.n24 24.4675
R235 VN.n26 VN.n25 24.4675
R236 VN.n31 VN.n30 24.4675
R237 VN.n32 VN.n31 24.4675
R238 VN.n50 VN.n49 24.4675
R239 VN.n49 VN.n48 24.4675
R240 VN.n48 VN.n43 24.4675
R241 VN.n61 VN.n60 24.4675
R242 VN.n60 VN.n59 24.4675
R243 VN.n56 VN.n55 24.4675
R244 VN.n55 VN.n54 24.4675
R245 VN.n54 VN.n41 24.4675
R246 VN.n67 VN.n66 24.4675
R247 VN.n66 VN.n65 24.4675
R248 VN.n24 VN.n4 20.7975
R249 VN.n59 VN.n39 20.7975
R250 VN.n32 VN.n0 11.0107
R251 VN.n67 VN.n35 11.0107
R252 VN.n46 VN.n45 4.35328
R253 VN.n11 VN.n10 4.35328
R254 VN.n9 VN.n8 3.67055
R255 VN.n21 VN.n4 3.67055
R256 VN.n44 VN.n43 3.67055
R257 VN.n56 VN.n39 3.67055
R258 VN.n69 VN.n68 0.354971
R259 VN.n34 VN.n33 0.354971
R260 VN VN.n34 0.26696
R261 VN.n68 VN.n36 0.189894
R262 VN.n64 VN.n36 0.189894
R263 VN.n64 VN.n63 0.189894
R264 VN.n63 VN.n62 0.189894
R265 VN.n62 VN.n38 0.189894
R266 VN.n58 VN.n38 0.189894
R267 VN.n58 VN.n57 0.189894
R268 VN.n57 VN.n40 0.189894
R269 VN.n53 VN.n40 0.189894
R270 VN.n53 VN.n52 0.189894
R271 VN.n52 VN.n51 0.189894
R272 VN.n51 VN.n42 0.189894
R273 VN.n47 VN.n42 0.189894
R274 VN.n47 VN.n46 0.189894
R275 VN.n12 VN.n11 0.189894
R276 VN.n12 VN.n7 0.189894
R277 VN.n16 VN.n7 0.189894
R278 VN.n17 VN.n16 0.189894
R279 VN.n18 VN.n17 0.189894
R280 VN.n18 VN.n5 0.189894
R281 VN.n22 VN.n5 0.189894
R282 VN.n23 VN.n22 0.189894
R283 VN.n23 VN.n3 0.189894
R284 VN.n27 VN.n3 0.189894
R285 VN.n28 VN.n27 0.189894
R286 VN.n29 VN.n28 0.189894
R287 VN.n29 VN.n1 0.189894
R288 VN.n33 VN.n1 0.189894
R289 VDD2.n2 VDD2.n1 75.2263
R290 VDD2.n2 VDD2.n0 75.2263
R291 VDD2 VDD2.n5 75.2235
R292 VDD2.n4 VDD2.n3 73.7086
R293 VDD2.n4 VDD2.n2 51.5903
R294 VDD2.n5 VDD2.t4 2.04355
R295 VDD2.n5 VDD2.t5 2.04355
R296 VDD2.n3 VDD2.t1 2.04355
R297 VDD2.n3 VDD2.t7 2.04355
R298 VDD2.n1 VDD2.t6 2.04355
R299 VDD2.n1 VDD2.t2 2.04355
R300 VDD2.n0 VDD2.t0 2.04355
R301 VDD2.n0 VDD2.t3 2.04355
R302 VDD2 VDD2.n4 1.63197
R303 B.n707 B.n706 585
R304 B.n708 B.n95 585
R305 B.n710 B.n709 585
R306 B.n711 B.n94 585
R307 B.n713 B.n712 585
R308 B.n714 B.n93 585
R309 B.n716 B.n715 585
R310 B.n717 B.n92 585
R311 B.n719 B.n718 585
R312 B.n720 B.n91 585
R313 B.n722 B.n721 585
R314 B.n723 B.n90 585
R315 B.n725 B.n724 585
R316 B.n726 B.n89 585
R317 B.n728 B.n727 585
R318 B.n729 B.n88 585
R319 B.n731 B.n730 585
R320 B.n732 B.n87 585
R321 B.n734 B.n733 585
R322 B.n735 B.n86 585
R323 B.n737 B.n736 585
R324 B.n738 B.n85 585
R325 B.n740 B.n739 585
R326 B.n741 B.n84 585
R327 B.n743 B.n742 585
R328 B.n744 B.n83 585
R329 B.n746 B.n745 585
R330 B.n747 B.n82 585
R331 B.n749 B.n748 585
R332 B.n750 B.n81 585
R333 B.n752 B.n751 585
R334 B.n753 B.n80 585
R335 B.n755 B.n754 585
R336 B.n756 B.n79 585
R337 B.n758 B.n757 585
R338 B.n759 B.n78 585
R339 B.n761 B.n760 585
R340 B.n762 B.n77 585
R341 B.n764 B.n763 585
R342 B.n765 B.n76 585
R343 B.n767 B.n766 585
R344 B.n768 B.n75 585
R345 B.n770 B.n769 585
R346 B.n771 B.n74 585
R347 B.n773 B.n772 585
R348 B.n774 B.n73 585
R349 B.n776 B.n775 585
R350 B.n777 B.n72 585
R351 B.n779 B.n778 585
R352 B.n780 B.n71 585
R353 B.n782 B.n781 585
R354 B.n783 B.n67 585
R355 B.n785 B.n784 585
R356 B.n786 B.n66 585
R357 B.n788 B.n787 585
R358 B.n789 B.n65 585
R359 B.n791 B.n790 585
R360 B.n792 B.n64 585
R361 B.n794 B.n793 585
R362 B.n795 B.n63 585
R363 B.n797 B.n796 585
R364 B.n798 B.n62 585
R365 B.n800 B.n799 585
R366 B.n802 B.n59 585
R367 B.n804 B.n803 585
R368 B.n805 B.n58 585
R369 B.n807 B.n806 585
R370 B.n808 B.n57 585
R371 B.n810 B.n809 585
R372 B.n811 B.n56 585
R373 B.n813 B.n812 585
R374 B.n814 B.n55 585
R375 B.n816 B.n815 585
R376 B.n817 B.n54 585
R377 B.n819 B.n818 585
R378 B.n820 B.n53 585
R379 B.n822 B.n821 585
R380 B.n823 B.n52 585
R381 B.n825 B.n824 585
R382 B.n826 B.n51 585
R383 B.n828 B.n827 585
R384 B.n829 B.n50 585
R385 B.n831 B.n830 585
R386 B.n832 B.n49 585
R387 B.n834 B.n833 585
R388 B.n835 B.n48 585
R389 B.n837 B.n836 585
R390 B.n838 B.n47 585
R391 B.n840 B.n839 585
R392 B.n841 B.n46 585
R393 B.n843 B.n842 585
R394 B.n844 B.n45 585
R395 B.n846 B.n845 585
R396 B.n847 B.n44 585
R397 B.n849 B.n848 585
R398 B.n850 B.n43 585
R399 B.n852 B.n851 585
R400 B.n853 B.n42 585
R401 B.n855 B.n854 585
R402 B.n856 B.n41 585
R403 B.n858 B.n857 585
R404 B.n859 B.n40 585
R405 B.n861 B.n860 585
R406 B.n862 B.n39 585
R407 B.n864 B.n863 585
R408 B.n865 B.n38 585
R409 B.n867 B.n866 585
R410 B.n868 B.n37 585
R411 B.n870 B.n869 585
R412 B.n871 B.n36 585
R413 B.n873 B.n872 585
R414 B.n874 B.n35 585
R415 B.n876 B.n875 585
R416 B.n877 B.n34 585
R417 B.n879 B.n878 585
R418 B.n880 B.n33 585
R419 B.n705 B.n96 585
R420 B.n704 B.n703 585
R421 B.n702 B.n97 585
R422 B.n701 B.n700 585
R423 B.n699 B.n98 585
R424 B.n698 B.n697 585
R425 B.n696 B.n99 585
R426 B.n695 B.n694 585
R427 B.n693 B.n100 585
R428 B.n692 B.n691 585
R429 B.n690 B.n101 585
R430 B.n689 B.n688 585
R431 B.n687 B.n102 585
R432 B.n686 B.n685 585
R433 B.n684 B.n103 585
R434 B.n683 B.n682 585
R435 B.n681 B.n104 585
R436 B.n680 B.n679 585
R437 B.n678 B.n105 585
R438 B.n677 B.n676 585
R439 B.n675 B.n106 585
R440 B.n674 B.n673 585
R441 B.n672 B.n107 585
R442 B.n671 B.n670 585
R443 B.n669 B.n108 585
R444 B.n668 B.n667 585
R445 B.n666 B.n109 585
R446 B.n665 B.n664 585
R447 B.n663 B.n110 585
R448 B.n662 B.n661 585
R449 B.n660 B.n111 585
R450 B.n659 B.n658 585
R451 B.n657 B.n112 585
R452 B.n656 B.n655 585
R453 B.n654 B.n113 585
R454 B.n653 B.n652 585
R455 B.n651 B.n114 585
R456 B.n650 B.n649 585
R457 B.n648 B.n115 585
R458 B.n647 B.n646 585
R459 B.n645 B.n116 585
R460 B.n644 B.n643 585
R461 B.n642 B.n117 585
R462 B.n641 B.n640 585
R463 B.n639 B.n118 585
R464 B.n638 B.n637 585
R465 B.n636 B.n119 585
R466 B.n635 B.n634 585
R467 B.n633 B.n120 585
R468 B.n632 B.n631 585
R469 B.n630 B.n121 585
R470 B.n629 B.n628 585
R471 B.n627 B.n122 585
R472 B.n626 B.n625 585
R473 B.n624 B.n123 585
R474 B.n623 B.n622 585
R475 B.n621 B.n124 585
R476 B.n620 B.n619 585
R477 B.n618 B.n125 585
R478 B.n617 B.n616 585
R479 B.n615 B.n126 585
R480 B.n614 B.n613 585
R481 B.n612 B.n127 585
R482 B.n611 B.n610 585
R483 B.n609 B.n128 585
R484 B.n608 B.n607 585
R485 B.n606 B.n129 585
R486 B.n605 B.n604 585
R487 B.n603 B.n130 585
R488 B.n602 B.n601 585
R489 B.n600 B.n131 585
R490 B.n599 B.n598 585
R491 B.n597 B.n132 585
R492 B.n596 B.n595 585
R493 B.n594 B.n133 585
R494 B.n593 B.n592 585
R495 B.n591 B.n134 585
R496 B.n590 B.n589 585
R497 B.n588 B.n135 585
R498 B.n587 B.n586 585
R499 B.n585 B.n136 585
R500 B.n584 B.n583 585
R501 B.n582 B.n137 585
R502 B.n581 B.n580 585
R503 B.n579 B.n138 585
R504 B.n578 B.n577 585
R505 B.n576 B.n139 585
R506 B.n575 B.n574 585
R507 B.n573 B.n140 585
R508 B.n572 B.n571 585
R509 B.n570 B.n141 585
R510 B.n569 B.n568 585
R511 B.n567 B.n142 585
R512 B.n566 B.n565 585
R513 B.n564 B.n143 585
R514 B.n563 B.n562 585
R515 B.n561 B.n144 585
R516 B.n560 B.n559 585
R517 B.n558 B.n145 585
R518 B.n557 B.n556 585
R519 B.n555 B.n146 585
R520 B.n554 B.n553 585
R521 B.n552 B.n147 585
R522 B.n551 B.n550 585
R523 B.n549 B.n148 585
R524 B.n548 B.n547 585
R525 B.n546 B.n149 585
R526 B.n545 B.n544 585
R527 B.n543 B.n150 585
R528 B.n542 B.n541 585
R529 B.n540 B.n151 585
R530 B.n539 B.n538 585
R531 B.n537 B.n152 585
R532 B.n536 B.n535 585
R533 B.n534 B.n153 585
R534 B.n533 B.n532 585
R535 B.n531 B.n154 585
R536 B.n530 B.n529 585
R537 B.n528 B.n155 585
R538 B.n527 B.n526 585
R539 B.n525 B.n156 585
R540 B.n524 B.n523 585
R541 B.n522 B.n157 585
R542 B.n521 B.n520 585
R543 B.n519 B.n158 585
R544 B.n344 B.n343 585
R545 B.n345 B.n220 585
R546 B.n347 B.n346 585
R547 B.n348 B.n219 585
R548 B.n350 B.n349 585
R549 B.n351 B.n218 585
R550 B.n353 B.n352 585
R551 B.n354 B.n217 585
R552 B.n356 B.n355 585
R553 B.n357 B.n216 585
R554 B.n359 B.n358 585
R555 B.n360 B.n215 585
R556 B.n362 B.n361 585
R557 B.n363 B.n214 585
R558 B.n365 B.n364 585
R559 B.n366 B.n213 585
R560 B.n368 B.n367 585
R561 B.n369 B.n212 585
R562 B.n371 B.n370 585
R563 B.n372 B.n211 585
R564 B.n374 B.n373 585
R565 B.n375 B.n210 585
R566 B.n377 B.n376 585
R567 B.n378 B.n209 585
R568 B.n380 B.n379 585
R569 B.n381 B.n208 585
R570 B.n383 B.n382 585
R571 B.n384 B.n207 585
R572 B.n386 B.n385 585
R573 B.n387 B.n206 585
R574 B.n389 B.n388 585
R575 B.n390 B.n205 585
R576 B.n392 B.n391 585
R577 B.n393 B.n204 585
R578 B.n395 B.n394 585
R579 B.n396 B.n203 585
R580 B.n398 B.n397 585
R581 B.n399 B.n202 585
R582 B.n401 B.n400 585
R583 B.n402 B.n201 585
R584 B.n404 B.n403 585
R585 B.n405 B.n200 585
R586 B.n407 B.n406 585
R587 B.n408 B.n199 585
R588 B.n410 B.n409 585
R589 B.n411 B.n198 585
R590 B.n413 B.n412 585
R591 B.n414 B.n197 585
R592 B.n416 B.n415 585
R593 B.n417 B.n196 585
R594 B.n419 B.n418 585
R595 B.n420 B.n195 585
R596 B.n422 B.n421 585
R597 B.n424 B.n192 585
R598 B.n426 B.n425 585
R599 B.n427 B.n191 585
R600 B.n429 B.n428 585
R601 B.n430 B.n190 585
R602 B.n432 B.n431 585
R603 B.n433 B.n189 585
R604 B.n435 B.n434 585
R605 B.n436 B.n188 585
R606 B.n438 B.n437 585
R607 B.n440 B.n439 585
R608 B.n441 B.n184 585
R609 B.n443 B.n442 585
R610 B.n444 B.n183 585
R611 B.n446 B.n445 585
R612 B.n447 B.n182 585
R613 B.n449 B.n448 585
R614 B.n450 B.n181 585
R615 B.n452 B.n451 585
R616 B.n453 B.n180 585
R617 B.n455 B.n454 585
R618 B.n456 B.n179 585
R619 B.n458 B.n457 585
R620 B.n459 B.n178 585
R621 B.n461 B.n460 585
R622 B.n462 B.n177 585
R623 B.n464 B.n463 585
R624 B.n465 B.n176 585
R625 B.n467 B.n466 585
R626 B.n468 B.n175 585
R627 B.n470 B.n469 585
R628 B.n471 B.n174 585
R629 B.n473 B.n472 585
R630 B.n474 B.n173 585
R631 B.n476 B.n475 585
R632 B.n477 B.n172 585
R633 B.n479 B.n478 585
R634 B.n480 B.n171 585
R635 B.n482 B.n481 585
R636 B.n483 B.n170 585
R637 B.n485 B.n484 585
R638 B.n486 B.n169 585
R639 B.n488 B.n487 585
R640 B.n489 B.n168 585
R641 B.n491 B.n490 585
R642 B.n492 B.n167 585
R643 B.n494 B.n493 585
R644 B.n495 B.n166 585
R645 B.n497 B.n496 585
R646 B.n498 B.n165 585
R647 B.n500 B.n499 585
R648 B.n501 B.n164 585
R649 B.n503 B.n502 585
R650 B.n504 B.n163 585
R651 B.n506 B.n505 585
R652 B.n507 B.n162 585
R653 B.n509 B.n508 585
R654 B.n510 B.n161 585
R655 B.n512 B.n511 585
R656 B.n513 B.n160 585
R657 B.n515 B.n514 585
R658 B.n516 B.n159 585
R659 B.n518 B.n517 585
R660 B.n342 B.n221 585
R661 B.n341 B.n340 585
R662 B.n339 B.n222 585
R663 B.n338 B.n337 585
R664 B.n336 B.n223 585
R665 B.n335 B.n334 585
R666 B.n333 B.n224 585
R667 B.n332 B.n331 585
R668 B.n330 B.n225 585
R669 B.n329 B.n328 585
R670 B.n327 B.n226 585
R671 B.n326 B.n325 585
R672 B.n324 B.n227 585
R673 B.n323 B.n322 585
R674 B.n321 B.n228 585
R675 B.n320 B.n319 585
R676 B.n318 B.n229 585
R677 B.n317 B.n316 585
R678 B.n315 B.n230 585
R679 B.n314 B.n313 585
R680 B.n312 B.n231 585
R681 B.n311 B.n310 585
R682 B.n309 B.n232 585
R683 B.n308 B.n307 585
R684 B.n306 B.n233 585
R685 B.n305 B.n304 585
R686 B.n303 B.n234 585
R687 B.n302 B.n301 585
R688 B.n300 B.n235 585
R689 B.n299 B.n298 585
R690 B.n297 B.n236 585
R691 B.n296 B.n295 585
R692 B.n294 B.n237 585
R693 B.n293 B.n292 585
R694 B.n291 B.n238 585
R695 B.n290 B.n289 585
R696 B.n288 B.n239 585
R697 B.n287 B.n286 585
R698 B.n285 B.n240 585
R699 B.n284 B.n283 585
R700 B.n282 B.n241 585
R701 B.n281 B.n280 585
R702 B.n279 B.n242 585
R703 B.n278 B.n277 585
R704 B.n276 B.n243 585
R705 B.n275 B.n274 585
R706 B.n273 B.n244 585
R707 B.n272 B.n271 585
R708 B.n270 B.n245 585
R709 B.n269 B.n268 585
R710 B.n267 B.n246 585
R711 B.n266 B.n265 585
R712 B.n264 B.n247 585
R713 B.n263 B.n262 585
R714 B.n261 B.n248 585
R715 B.n260 B.n259 585
R716 B.n258 B.n249 585
R717 B.n257 B.n256 585
R718 B.n255 B.n250 585
R719 B.n254 B.n253 585
R720 B.n252 B.n251 585
R721 B.n2 B.n0 585
R722 B.n973 B.n1 585
R723 B.n972 B.n971 585
R724 B.n970 B.n3 585
R725 B.n969 B.n968 585
R726 B.n967 B.n4 585
R727 B.n966 B.n965 585
R728 B.n964 B.n5 585
R729 B.n963 B.n962 585
R730 B.n961 B.n6 585
R731 B.n960 B.n959 585
R732 B.n958 B.n7 585
R733 B.n957 B.n956 585
R734 B.n955 B.n8 585
R735 B.n954 B.n953 585
R736 B.n952 B.n9 585
R737 B.n951 B.n950 585
R738 B.n949 B.n10 585
R739 B.n948 B.n947 585
R740 B.n946 B.n11 585
R741 B.n945 B.n944 585
R742 B.n943 B.n12 585
R743 B.n942 B.n941 585
R744 B.n940 B.n13 585
R745 B.n939 B.n938 585
R746 B.n937 B.n14 585
R747 B.n936 B.n935 585
R748 B.n934 B.n15 585
R749 B.n933 B.n932 585
R750 B.n931 B.n16 585
R751 B.n930 B.n929 585
R752 B.n928 B.n17 585
R753 B.n927 B.n926 585
R754 B.n925 B.n18 585
R755 B.n924 B.n923 585
R756 B.n922 B.n19 585
R757 B.n921 B.n920 585
R758 B.n919 B.n20 585
R759 B.n918 B.n917 585
R760 B.n916 B.n21 585
R761 B.n915 B.n914 585
R762 B.n913 B.n22 585
R763 B.n912 B.n911 585
R764 B.n910 B.n23 585
R765 B.n909 B.n908 585
R766 B.n907 B.n24 585
R767 B.n906 B.n905 585
R768 B.n904 B.n25 585
R769 B.n903 B.n902 585
R770 B.n901 B.n26 585
R771 B.n900 B.n899 585
R772 B.n898 B.n27 585
R773 B.n897 B.n896 585
R774 B.n895 B.n28 585
R775 B.n894 B.n893 585
R776 B.n892 B.n29 585
R777 B.n891 B.n890 585
R778 B.n889 B.n30 585
R779 B.n888 B.n887 585
R780 B.n886 B.n31 585
R781 B.n885 B.n884 585
R782 B.n883 B.n32 585
R783 B.n882 B.n881 585
R784 B.n975 B.n974 585
R785 B.n343 B.n342 449.257
R786 B.n882 B.n33 449.257
R787 B.n517 B.n158 449.257
R788 B.n707 B.n96 449.257
R789 B.n185 B.t0 324.416
R790 B.n193 B.t9 324.416
R791 B.n60 B.t3 324.416
R792 B.n68 B.t6 324.416
R793 B.n185 B.t2 182.463
R794 B.n68 B.t7 182.463
R795 B.n193 B.t11 182.442
R796 B.n60 B.t4 182.442
R797 B.n342 B.n341 163.367
R798 B.n341 B.n222 163.367
R799 B.n337 B.n222 163.367
R800 B.n337 B.n336 163.367
R801 B.n336 B.n335 163.367
R802 B.n335 B.n224 163.367
R803 B.n331 B.n224 163.367
R804 B.n331 B.n330 163.367
R805 B.n330 B.n329 163.367
R806 B.n329 B.n226 163.367
R807 B.n325 B.n226 163.367
R808 B.n325 B.n324 163.367
R809 B.n324 B.n323 163.367
R810 B.n323 B.n228 163.367
R811 B.n319 B.n228 163.367
R812 B.n319 B.n318 163.367
R813 B.n318 B.n317 163.367
R814 B.n317 B.n230 163.367
R815 B.n313 B.n230 163.367
R816 B.n313 B.n312 163.367
R817 B.n312 B.n311 163.367
R818 B.n311 B.n232 163.367
R819 B.n307 B.n232 163.367
R820 B.n307 B.n306 163.367
R821 B.n306 B.n305 163.367
R822 B.n305 B.n234 163.367
R823 B.n301 B.n234 163.367
R824 B.n301 B.n300 163.367
R825 B.n300 B.n299 163.367
R826 B.n299 B.n236 163.367
R827 B.n295 B.n236 163.367
R828 B.n295 B.n294 163.367
R829 B.n294 B.n293 163.367
R830 B.n293 B.n238 163.367
R831 B.n289 B.n238 163.367
R832 B.n289 B.n288 163.367
R833 B.n288 B.n287 163.367
R834 B.n287 B.n240 163.367
R835 B.n283 B.n240 163.367
R836 B.n283 B.n282 163.367
R837 B.n282 B.n281 163.367
R838 B.n281 B.n242 163.367
R839 B.n277 B.n242 163.367
R840 B.n277 B.n276 163.367
R841 B.n276 B.n275 163.367
R842 B.n275 B.n244 163.367
R843 B.n271 B.n244 163.367
R844 B.n271 B.n270 163.367
R845 B.n270 B.n269 163.367
R846 B.n269 B.n246 163.367
R847 B.n265 B.n246 163.367
R848 B.n265 B.n264 163.367
R849 B.n264 B.n263 163.367
R850 B.n263 B.n248 163.367
R851 B.n259 B.n248 163.367
R852 B.n259 B.n258 163.367
R853 B.n258 B.n257 163.367
R854 B.n257 B.n250 163.367
R855 B.n253 B.n250 163.367
R856 B.n253 B.n252 163.367
R857 B.n252 B.n2 163.367
R858 B.n974 B.n2 163.367
R859 B.n974 B.n973 163.367
R860 B.n973 B.n972 163.367
R861 B.n972 B.n3 163.367
R862 B.n968 B.n3 163.367
R863 B.n968 B.n967 163.367
R864 B.n967 B.n966 163.367
R865 B.n966 B.n5 163.367
R866 B.n962 B.n5 163.367
R867 B.n962 B.n961 163.367
R868 B.n961 B.n960 163.367
R869 B.n960 B.n7 163.367
R870 B.n956 B.n7 163.367
R871 B.n956 B.n955 163.367
R872 B.n955 B.n954 163.367
R873 B.n954 B.n9 163.367
R874 B.n950 B.n9 163.367
R875 B.n950 B.n949 163.367
R876 B.n949 B.n948 163.367
R877 B.n948 B.n11 163.367
R878 B.n944 B.n11 163.367
R879 B.n944 B.n943 163.367
R880 B.n943 B.n942 163.367
R881 B.n942 B.n13 163.367
R882 B.n938 B.n13 163.367
R883 B.n938 B.n937 163.367
R884 B.n937 B.n936 163.367
R885 B.n936 B.n15 163.367
R886 B.n932 B.n15 163.367
R887 B.n932 B.n931 163.367
R888 B.n931 B.n930 163.367
R889 B.n930 B.n17 163.367
R890 B.n926 B.n17 163.367
R891 B.n926 B.n925 163.367
R892 B.n925 B.n924 163.367
R893 B.n924 B.n19 163.367
R894 B.n920 B.n19 163.367
R895 B.n920 B.n919 163.367
R896 B.n919 B.n918 163.367
R897 B.n918 B.n21 163.367
R898 B.n914 B.n21 163.367
R899 B.n914 B.n913 163.367
R900 B.n913 B.n912 163.367
R901 B.n912 B.n23 163.367
R902 B.n908 B.n23 163.367
R903 B.n908 B.n907 163.367
R904 B.n907 B.n906 163.367
R905 B.n906 B.n25 163.367
R906 B.n902 B.n25 163.367
R907 B.n902 B.n901 163.367
R908 B.n901 B.n900 163.367
R909 B.n900 B.n27 163.367
R910 B.n896 B.n27 163.367
R911 B.n896 B.n895 163.367
R912 B.n895 B.n894 163.367
R913 B.n894 B.n29 163.367
R914 B.n890 B.n29 163.367
R915 B.n890 B.n889 163.367
R916 B.n889 B.n888 163.367
R917 B.n888 B.n31 163.367
R918 B.n884 B.n31 163.367
R919 B.n884 B.n883 163.367
R920 B.n883 B.n882 163.367
R921 B.n343 B.n220 163.367
R922 B.n347 B.n220 163.367
R923 B.n348 B.n347 163.367
R924 B.n349 B.n348 163.367
R925 B.n349 B.n218 163.367
R926 B.n353 B.n218 163.367
R927 B.n354 B.n353 163.367
R928 B.n355 B.n354 163.367
R929 B.n355 B.n216 163.367
R930 B.n359 B.n216 163.367
R931 B.n360 B.n359 163.367
R932 B.n361 B.n360 163.367
R933 B.n361 B.n214 163.367
R934 B.n365 B.n214 163.367
R935 B.n366 B.n365 163.367
R936 B.n367 B.n366 163.367
R937 B.n367 B.n212 163.367
R938 B.n371 B.n212 163.367
R939 B.n372 B.n371 163.367
R940 B.n373 B.n372 163.367
R941 B.n373 B.n210 163.367
R942 B.n377 B.n210 163.367
R943 B.n378 B.n377 163.367
R944 B.n379 B.n378 163.367
R945 B.n379 B.n208 163.367
R946 B.n383 B.n208 163.367
R947 B.n384 B.n383 163.367
R948 B.n385 B.n384 163.367
R949 B.n385 B.n206 163.367
R950 B.n389 B.n206 163.367
R951 B.n390 B.n389 163.367
R952 B.n391 B.n390 163.367
R953 B.n391 B.n204 163.367
R954 B.n395 B.n204 163.367
R955 B.n396 B.n395 163.367
R956 B.n397 B.n396 163.367
R957 B.n397 B.n202 163.367
R958 B.n401 B.n202 163.367
R959 B.n402 B.n401 163.367
R960 B.n403 B.n402 163.367
R961 B.n403 B.n200 163.367
R962 B.n407 B.n200 163.367
R963 B.n408 B.n407 163.367
R964 B.n409 B.n408 163.367
R965 B.n409 B.n198 163.367
R966 B.n413 B.n198 163.367
R967 B.n414 B.n413 163.367
R968 B.n415 B.n414 163.367
R969 B.n415 B.n196 163.367
R970 B.n419 B.n196 163.367
R971 B.n420 B.n419 163.367
R972 B.n421 B.n420 163.367
R973 B.n421 B.n192 163.367
R974 B.n426 B.n192 163.367
R975 B.n427 B.n426 163.367
R976 B.n428 B.n427 163.367
R977 B.n428 B.n190 163.367
R978 B.n432 B.n190 163.367
R979 B.n433 B.n432 163.367
R980 B.n434 B.n433 163.367
R981 B.n434 B.n188 163.367
R982 B.n438 B.n188 163.367
R983 B.n439 B.n438 163.367
R984 B.n439 B.n184 163.367
R985 B.n443 B.n184 163.367
R986 B.n444 B.n443 163.367
R987 B.n445 B.n444 163.367
R988 B.n445 B.n182 163.367
R989 B.n449 B.n182 163.367
R990 B.n450 B.n449 163.367
R991 B.n451 B.n450 163.367
R992 B.n451 B.n180 163.367
R993 B.n455 B.n180 163.367
R994 B.n456 B.n455 163.367
R995 B.n457 B.n456 163.367
R996 B.n457 B.n178 163.367
R997 B.n461 B.n178 163.367
R998 B.n462 B.n461 163.367
R999 B.n463 B.n462 163.367
R1000 B.n463 B.n176 163.367
R1001 B.n467 B.n176 163.367
R1002 B.n468 B.n467 163.367
R1003 B.n469 B.n468 163.367
R1004 B.n469 B.n174 163.367
R1005 B.n473 B.n174 163.367
R1006 B.n474 B.n473 163.367
R1007 B.n475 B.n474 163.367
R1008 B.n475 B.n172 163.367
R1009 B.n479 B.n172 163.367
R1010 B.n480 B.n479 163.367
R1011 B.n481 B.n480 163.367
R1012 B.n481 B.n170 163.367
R1013 B.n485 B.n170 163.367
R1014 B.n486 B.n485 163.367
R1015 B.n487 B.n486 163.367
R1016 B.n487 B.n168 163.367
R1017 B.n491 B.n168 163.367
R1018 B.n492 B.n491 163.367
R1019 B.n493 B.n492 163.367
R1020 B.n493 B.n166 163.367
R1021 B.n497 B.n166 163.367
R1022 B.n498 B.n497 163.367
R1023 B.n499 B.n498 163.367
R1024 B.n499 B.n164 163.367
R1025 B.n503 B.n164 163.367
R1026 B.n504 B.n503 163.367
R1027 B.n505 B.n504 163.367
R1028 B.n505 B.n162 163.367
R1029 B.n509 B.n162 163.367
R1030 B.n510 B.n509 163.367
R1031 B.n511 B.n510 163.367
R1032 B.n511 B.n160 163.367
R1033 B.n515 B.n160 163.367
R1034 B.n516 B.n515 163.367
R1035 B.n517 B.n516 163.367
R1036 B.n521 B.n158 163.367
R1037 B.n522 B.n521 163.367
R1038 B.n523 B.n522 163.367
R1039 B.n523 B.n156 163.367
R1040 B.n527 B.n156 163.367
R1041 B.n528 B.n527 163.367
R1042 B.n529 B.n528 163.367
R1043 B.n529 B.n154 163.367
R1044 B.n533 B.n154 163.367
R1045 B.n534 B.n533 163.367
R1046 B.n535 B.n534 163.367
R1047 B.n535 B.n152 163.367
R1048 B.n539 B.n152 163.367
R1049 B.n540 B.n539 163.367
R1050 B.n541 B.n540 163.367
R1051 B.n541 B.n150 163.367
R1052 B.n545 B.n150 163.367
R1053 B.n546 B.n545 163.367
R1054 B.n547 B.n546 163.367
R1055 B.n547 B.n148 163.367
R1056 B.n551 B.n148 163.367
R1057 B.n552 B.n551 163.367
R1058 B.n553 B.n552 163.367
R1059 B.n553 B.n146 163.367
R1060 B.n557 B.n146 163.367
R1061 B.n558 B.n557 163.367
R1062 B.n559 B.n558 163.367
R1063 B.n559 B.n144 163.367
R1064 B.n563 B.n144 163.367
R1065 B.n564 B.n563 163.367
R1066 B.n565 B.n564 163.367
R1067 B.n565 B.n142 163.367
R1068 B.n569 B.n142 163.367
R1069 B.n570 B.n569 163.367
R1070 B.n571 B.n570 163.367
R1071 B.n571 B.n140 163.367
R1072 B.n575 B.n140 163.367
R1073 B.n576 B.n575 163.367
R1074 B.n577 B.n576 163.367
R1075 B.n577 B.n138 163.367
R1076 B.n581 B.n138 163.367
R1077 B.n582 B.n581 163.367
R1078 B.n583 B.n582 163.367
R1079 B.n583 B.n136 163.367
R1080 B.n587 B.n136 163.367
R1081 B.n588 B.n587 163.367
R1082 B.n589 B.n588 163.367
R1083 B.n589 B.n134 163.367
R1084 B.n593 B.n134 163.367
R1085 B.n594 B.n593 163.367
R1086 B.n595 B.n594 163.367
R1087 B.n595 B.n132 163.367
R1088 B.n599 B.n132 163.367
R1089 B.n600 B.n599 163.367
R1090 B.n601 B.n600 163.367
R1091 B.n601 B.n130 163.367
R1092 B.n605 B.n130 163.367
R1093 B.n606 B.n605 163.367
R1094 B.n607 B.n606 163.367
R1095 B.n607 B.n128 163.367
R1096 B.n611 B.n128 163.367
R1097 B.n612 B.n611 163.367
R1098 B.n613 B.n612 163.367
R1099 B.n613 B.n126 163.367
R1100 B.n617 B.n126 163.367
R1101 B.n618 B.n617 163.367
R1102 B.n619 B.n618 163.367
R1103 B.n619 B.n124 163.367
R1104 B.n623 B.n124 163.367
R1105 B.n624 B.n623 163.367
R1106 B.n625 B.n624 163.367
R1107 B.n625 B.n122 163.367
R1108 B.n629 B.n122 163.367
R1109 B.n630 B.n629 163.367
R1110 B.n631 B.n630 163.367
R1111 B.n631 B.n120 163.367
R1112 B.n635 B.n120 163.367
R1113 B.n636 B.n635 163.367
R1114 B.n637 B.n636 163.367
R1115 B.n637 B.n118 163.367
R1116 B.n641 B.n118 163.367
R1117 B.n642 B.n641 163.367
R1118 B.n643 B.n642 163.367
R1119 B.n643 B.n116 163.367
R1120 B.n647 B.n116 163.367
R1121 B.n648 B.n647 163.367
R1122 B.n649 B.n648 163.367
R1123 B.n649 B.n114 163.367
R1124 B.n653 B.n114 163.367
R1125 B.n654 B.n653 163.367
R1126 B.n655 B.n654 163.367
R1127 B.n655 B.n112 163.367
R1128 B.n659 B.n112 163.367
R1129 B.n660 B.n659 163.367
R1130 B.n661 B.n660 163.367
R1131 B.n661 B.n110 163.367
R1132 B.n665 B.n110 163.367
R1133 B.n666 B.n665 163.367
R1134 B.n667 B.n666 163.367
R1135 B.n667 B.n108 163.367
R1136 B.n671 B.n108 163.367
R1137 B.n672 B.n671 163.367
R1138 B.n673 B.n672 163.367
R1139 B.n673 B.n106 163.367
R1140 B.n677 B.n106 163.367
R1141 B.n678 B.n677 163.367
R1142 B.n679 B.n678 163.367
R1143 B.n679 B.n104 163.367
R1144 B.n683 B.n104 163.367
R1145 B.n684 B.n683 163.367
R1146 B.n685 B.n684 163.367
R1147 B.n685 B.n102 163.367
R1148 B.n689 B.n102 163.367
R1149 B.n690 B.n689 163.367
R1150 B.n691 B.n690 163.367
R1151 B.n691 B.n100 163.367
R1152 B.n695 B.n100 163.367
R1153 B.n696 B.n695 163.367
R1154 B.n697 B.n696 163.367
R1155 B.n697 B.n98 163.367
R1156 B.n701 B.n98 163.367
R1157 B.n702 B.n701 163.367
R1158 B.n703 B.n702 163.367
R1159 B.n703 B.n96 163.367
R1160 B.n878 B.n33 163.367
R1161 B.n878 B.n877 163.367
R1162 B.n877 B.n876 163.367
R1163 B.n876 B.n35 163.367
R1164 B.n872 B.n35 163.367
R1165 B.n872 B.n871 163.367
R1166 B.n871 B.n870 163.367
R1167 B.n870 B.n37 163.367
R1168 B.n866 B.n37 163.367
R1169 B.n866 B.n865 163.367
R1170 B.n865 B.n864 163.367
R1171 B.n864 B.n39 163.367
R1172 B.n860 B.n39 163.367
R1173 B.n860 B.n859 163.367
R1174 B.n859 B.n858 163.367
R1175 B.n858 B.n41 163.367
R1176 B.n854 B.n41 163.367
R1177 B.n854 B.n853 163.367
R1178 B.n853 B.n852 163.367
R1179 B.n852 B.n43 163.367
R1180 B.n848 B.n43 163.367
R1181 B.n848 B.n847 163.367
R1182 B.n847 B.n846 163.367
R1183 B.n846 B.n45 163.367
R1184 B.n842 B.n45 163.367
R1185 B.n842 B.n841 163.367
R1186 B.n841 B.n840 163.367
R1187 B.n840 B.n47 163.367
R1188 B.n836 B.n47 163.367
R1189 B.n836 B.n835 163.367
R1190 B.n835 B.n834 163.367
R1191 B.n834 B.n49 163.367
R1192 B.n830 B.n49 163.367
R1193 B.n830 B.n829 163.367
R1194 B.n829 B.n828 163.367
R1195 B.n828 B.n51 163.367
R1196 B.n824 B.n51 163.367
R1197 B.n824 B.n823 163.367
R1198 B.n823 B.n822 163.367
R1199 B.n822 B.n53 163.367
R1200 B.n818 B.n53 163.367
R1201 B.n818 B.n817 163.367
R1202 B.n817 B.n816 163.367
R1203 B.n816 B.n55 163.367
R1204 B.n812 B.n55 163.367
R1205 B.n812 B.n811 163.367
R1206 B.n811 B.n810 163.367
R1207 B.n810 B.n57 163.367
R1208 B.n806 B.n57 163.367
R1209 B.n806 B.n805 163.367
R1210 B.n805 B.n804 163.367
R1211 B.n804 B.n59 163.367
R1212 B.n799 B.n59 163.367
R1213 B.n799 B.n798 163.367
R1214 B.n798 B.n797 163.367
R1215 B.n797 B.n63 163.367
R1216 B.n793 B.n63 163.367
R1217 B.n793 B.n792 163.367
R1218 B.n792 B.n791 163.367
R1219 B.n791 B.n65 163.367
R1220 B.n787 B.n65 163.367
R1221 B.n787 B.n786 163.367
R1222 B.n786 B.n785 163.367
R1223 B.n785 B.n67 163.367
R1224 B.n781 B.n67 163.367
R1225 B.n781 B.n780 163.367
R1226 B.n780 B.n779 163.367
R1227 B.n779 B.n72 163.367
R1228 B.n775 B.n72 163.367
R1229 B.n775 B.n774 163.367
R1230 B.n774 B.n773 163.367
R1231 B.n773 B.n74 163.367
R1232 B.n769 B.n74 163.367
R1233 B.n769 B.n768 163.367
R1234 B.n768 B.n767 163.367
R1235 B.n767 B.n76 163.367
R1236 B.n763 B.n76 163.367
R1237 B.n763 B.n762 163.367
R1238 B.n762 B.n761 163.367
R1239 B.n761 B.n78 163.367
R1240 B.n757 B.n78 163.367
R1241 B.n757 B.n756 163.367
R1242 B.n756 B.n755 163.367
R1243 B.n755 B.n80 163.367
R1244 B.n751 B.n80 163.367
R1245 B.n751 B.n750 163.367
R1246 B.n750 B.n749 163.367
R1247 B.n749 B.n82 163.367
R1248 B.n745 B.n82 163.367
R1249 B.n745 B.n744 163.367
R1250 B.n744 B.n743 163.367
R1251 B.n743 B.n84 163.367
R1252 B.n739 B.n84 163.367
R1253 B.n739 B.n738 163.367
R1254 B.n738 B.n737 163.367
R1255 B.n737 B.n86 163.367
R1256 B.n733 B.n86 163.367
R1257 B.n733 B.n732 163.367
R1258 B.n732 B.n731 163.367
R1259 B.n731 B.n88 163.367
R1260 B.n727 B.n88 163.367
R1261 B.n727 B.n726 163.367
R1262 B.n726 B.n725 163.367
R1263 B.n725 B.n90 163.367
R1264 B.n721 B.n90 163.367
R1265 B.n721 B.n720 163.367
R1266 B.n720 B.n719 163.367
R1267 B.n719 B.n92 163.367
R1268 B.n715 B.n92 163.367
R1269 B.n715 B.n714 163.367
R1270 B.n714 B.n713 163.367
R1271 B.n713 B.n94 163.367
R1272 B.n709 B.n94 163.367
R1273 B.n709 B.n708 163.367
R1274 B.n708 B.n707 163.367
R1275 B.n186 B.t1 111.674
R1276 B.n69 B.t8 111.674
R1277 B.n194 B.t10 111.654
R1278 B.n61 B.t5 111.654
R1279 B.n186 B.n185 70.7884
R1280 B.n194 B.n193 70.7884
R1281 B.n61 B.n60 70.7884
R1282 B.n69 B.n68 70.7884
R1283 B.n187 B.n186 59.5399
R1284 B.n423 B.n194 59.5399
R1285 B.n801 B.n61 59.5399
R1286 B.n70 B.n69 59.5399
R1287 B.n881 B.n880 29.1907
R1288 B.n519 B.n518 29.1907
R1289 B.n344 B.n221 29.1907
R1290 B.n706 B.n705 29.1907
R1291 B B.n975 18.0485
R1292 B.n880 B.n879 10.6151
R1293 B.n879 B.n34 10.6151
R1294 B.n875 B.n34 10.6151
R1295 B.n875 B.n874 10.6151
R1296 B.n874 B.n873 10.6151
R1297 B.n873 B.n36 10.6151
R1298 B.n869 B.n36 10.6151
R1299 B.n869 B.n868 10.6151
R1300 B.n868 B.n867 10.6151
R1301 B.n867 B.n38 10.6151
R1302 B.n863 B.n38 10.6151
R1303 B.n863 B.n862 10.6151
R1304 B.n862 B.n861 10.6151
R1305 B.n861 B.n40 10.6151
R1306 B.n857 B.n40 10.6151
R1307 B.n857 B.n856 10.6151
R1308 B.n856 B.n855 10.6151
R1309 B.n855 B.n42 10.6151
R1310 B.n851 B.n42 10.6151
R1311 B.n851 B.n850 10.6151
R1312 B.n850 B.n849 10.6151
R1313 B.n849 B.n44 10.6151
R1314 B.n845 B.n44 10.6151
R1315 B.n845 B.n844 10.6151
R1316 B.n844 B.n843 10.6151
R1317 B.n843 B.n46 10.6151
R1318 B.n839 B.n46 10.6151
R1319 B.n839 B.n838 10.6151
R1320 B.n838 B.n837 10.6151
R1321 B.n837 B.n48 10.6151
R1322 B.n833 B.n48 10.6151
R1323 B.n833 B.n832 10.6151
R1324 B.n832 B.n831 10.6151
R1325 B.n831 B.n50 10.6151
R1326 B.n827 B.n50 10.6151
R1327 B.n827 B.n826 10.6151
R1328 B.n826 B.n825 10.6151
R1329 B.n825 B.n52 10.6151
R1330 B.n821 B.n52 10.6151
R1331 B.n821 B.n820 10.6151
R1332 B.n820 B.n819 10.6151
R1333 B.n819 B.n54 10.6151
R1334 B.n815 B.n54 10.6151
R1335 B.n815 B.n814 10.6151
R1336 B.n814 B.n813 10.6151
R1337 B.n813 B.n56 10.6151
R1338 B.n809 B.n56 10.6151
R1339 B.n809 B.n808 10.6151
R1340 B.n808 B.n807 10.6151
R1341 B.n807 B.n58 10.6151
R1342 B.n803 B.n58 10.6151
R1343 B.n803 B.n802 10.6151
R1344 B.n800 B.n62 10.6151
R1345 B.n796 B.n62 10.6151
R1346 B.n796 B.n795 10.6151
R1347 B.n795 B.n794 10.6151
R1348 B.n794 B.n64 10.6151
R1349 B.n790 B.n64 10.6151
R1350 B.n790 B.n789 10.6151
R1351 B.n789 B.n788 10.6151
R1352 B.n788 B.n66 10.6151
R1353 B.n784 B.n783 10.6151
R1354 B.n783 B.n782 10.6151
R1355 B.n782 B.n71 10.6151
R1356 B.n778 B.n71 10.6151
R1357 B.n778 B.n777 10.6151
R1358 B.n777 B.n776 10.6151
R1359 B.n776 B.n73 10.6151
R1360 B.n772 B.n73 10.6151
R1361 B.n772 B.n771 10.6151
R1362 B.n771 B.n770 10.6151
R1363 B.n770 B.n75 10.6151
R1364 B.n766 B.n75 10.6151
R1365 B.n766 B.n765 10.6151
R1366 B.n765 B.n764 10.6151
R1367 B.n764 B.n77 10.6151
R1368 B.n760 B.n77 10.6151
R1369 B.n760 B.n759 10.6151
R1370 B.n759 B.n758 10.6151
R1371 B.n758 B.n79 10.6151
R1372 B.n754 B.n79 10.6151
R1373 B.n754 B.n753 10.6151
R1374 B.n753 B.n752 10.6151
R1375 B.n752 B.n81 10.6151
R1376 B.n748 B.n81 10.6151
R1377 B.n748 B.n747 10.6151
R1378 B.n747 B.n746 10.6151
R1379 B.n746 B.n83 10.6151
R1380 B.n742 B.n83 10.6151
R1381 B.n742 B.n741 10.6151
R1382 B.n741 B.n740 10.6151
R1383 B.n740 B.n85 10.6151
R1384 B.n736 B.n85 10.6151
R1385 B.n736 B.n735 10.6151
R1386 B.n735 B.n734 10.6151
R1387 B.n734 B.n87 10.6151
R1388 B.n730 B.n87 10.6151
R1389 B.n730 B.n729 10.6151
R1390 B.n729 B.n728 10.6151
R1391 B.n728 B.n89 10.6151
R1392 B.n724 B.n89 10.6151
R1393 B.n724 B.n723 10.6151
R1394 B.n723 B.n722 10.6151
R1395 B.n722 B.n91 10.6151
R1396 B.n718 B.n91 10.6151
R1397 B.n718 B.n717 10.6151
R1398 B.n717 B.n716 10.6151
R1399 B.n716 B.n93 10.6151
R1400 B.n712 B.n93 10.6151
R1401 B.n712 B.n711 10.6151
R1402 B.n711 B.n710 10.6151
R1403 B.n710 B.n95 10.6151
R1404 B.n706 B.n95 10.6151
R1405 B.n520 B.n519 10.6151
R1406 B.n520 B.n157 10.6151
R1407 B.n524 B.n157 10.6151
R1408 B.n525 B.n524 10.6151
R1409 B.n526 B.n525 10.6151
R1410 B.n526 B.n155 10.6151
R1411 B.n530 B.n155 10.6151
R1412 B.n531 B.n530 10.6151
R1413 B.n532 B.n531 10.6151
R1414 B.n532 B.n153 10.6151
R1415 B.n536 B.n153 10.6151
R1416 B.n537 B.n536 10.6151
R1417 B.n538 B.n537 10.6151
R1418 B.n538 B.n151 10.6151
R1419 B.n542 B.n151 10.6151
R1420 B.n543 B.n542 10.6151
R1421 B.n544 B.n543 10.6151
R1422 B.n544 B.n149 10.6151
R1423 B.n548 B.n149 10.6151
R1424 B.n549 B.n548 10.6151
R1425 B.n550 B.n549 10.6151
R1426 B.n550 B.n147 10.6151
R1427 B.n554 B.n147 10.6151
R1428 B.n555 B.n554 10.6151
R1429 B.n556 B.n555 10.6151
R1430 B.n556 B.n145 10.6151
R1431 B.n560 B.n145 10.6151
R1432 B.n561 B.n560 10.6151
R1433 B.n562 B.n561 10.6151
R1434 B.n562 B.n143 10.6151
R1435 B.n566 B.n143 10.6151
R1436 B.n567 B.n566 10.6151
R1437 B.n568 B.n567 10.6151
R1438 B.n568 B.n141 10.6151
R1439 B.n572 B.n141 10.6151
R1440 B.n573 B.n572 10.6151
R1441 B.n574 B.n573 10.6151
R1442 B.n574 B.n139 10.6151
R1443 B.n578 B.n139 10.6151
R1444 B.n579 B.n578 10.6151
R1445 B.n580 B.n579 10.6151
R1446 B.n580 B.n137 10.6151
R1447 B.n584 B.n137 10.6151
R1448 B.n585 B.n584 10.6151
R1449 B.n586 B.n585 10.6151
R1450 B.n586 B.n135 10.6151
R1451 B.n590 B.n135 10.6151
R1452 B.n591 B.n590 10.6151
R1453 B.n592 B.n591 10.6151
R1454 B.n592 B.n133 10.6151
R1455 B.n596 B.n133 10.6151
R1456 B.n597 B.n596 10.6151
R1457 B.n598 B.n597 10.6151
R1458 B.n598 B.n131 10.6151
R1459 B.n602 B.n131 10.6151
R1460 B.n603 B.n602 10.6151
R1461 B.n604 B.n603 10.6151
R1462 B.n604 B.n129 10.6151
R1463 B.n608 B.n129 10.6151
R1464 B.n609 B.n608 10.6151
R1465 B.n610 B.n609 10.6151
R1466 B.n610 B.n127 10.6151
R1467 B.n614 B.n127 10.6151
R1468 B.n615 B.n614 10.6151
R1469 B.n616 B.n615 10.6151
R1470 B.n616 B.n125 10.6151
R1471 B.n620 B.n125 10.6151
R1472 B.n621 B.n620 10.6151
R1473 B.n622 B.n621 10.6151
R1474 B.n622 B.n123 10.6151
R1475 B.n626 B.n123 10.6151
R1476 B.n627 B.n626 10.6151
R1477 B.n628 B.n627 10.6151
R1478 B.n628 B.n121 10.6151
R1479 B.n632 B.n121 10.6151
R1480 B.n633 B.n632 10.6151
R1481 B.n634 B.n633 10.6151
R1482 B.n634 B.n119 10.6151
R1483 B.n638 B.n119 10.6151
R1484 B.n639 B.n638 10.6151
R1485 B.n640 B.n639 10.6151
R1486 B.n640 B.n117 10.6151
R1487 B.n644 B.n117 10.6151
R1488 B.n645 B.n644 10.6151
R1489 B.n646 B.n645 10.6151
R1490 B.n646 B.n115 10.6151
R1491 B.n650 B.n115 10.6151
R1492 B.n651 B.n650 10.6151
R1493 B.n652 B.n651 10.6151
R1494 B.n652 B.n113 10.6151
R1495 B.n656 B.n113 10.6151
R1496 B.n657 B.n656 10.6151
R1497 B.n658 B.n657 10.6151
R1498 B.n658 B.n111 10.6151
R1499 B.n662 B.n111 10.6151
R1500 B.n663 B.n662 10.6151
R1501 B.n664 B.n663 10.6151
R1502 B.n664 B.n109 10.6151
R1503 B.n668 B.n109 10.6151
R1504 B.n669 B.n668 10.6151
R1505 B.n670 B.n669 10.6151
R1506 B.n670 B.n107 10.6151
R1507 B.n674 B.n107 10.6151
R1508 B.n675 B.n674 10.6151
R1509 B.n676 B.n675 10.6151
R1510 B.n676 B.n105 10.6151
R1511 B.n680 B.n105 10.6151
R1512 B.n681 B.n680 10.6151
R1513 B.n682 B.n681 10.6151
R1514 B.n682 B.n103 10.6151
R1515 B.n686 B.n103 10.6151
R1516 B.n687 B.n686 10.6151
R1517 B.n688 B.n687 10.6151
R1518 B.n688 B.n101 10.6151
R1519 B.n692 B.n101 10.6151
R1520 B.n693 B.n692 10.6151
R1521 B.n694 B.n693 10.6151
R1522 B.n694 B.n99 10.6151
R1523 B.n698 B.n99 10.6151
R1524 B.n699 B.n698 10.6151
R1525 B.n700 B.n699 10.6151
R1526 B.n700 B.n97 10.6151
R1527 B.n704 B.n97 10.6151
R1528 B.n705 B.n704 10.6151
R1529 B.n345 B.n344 10.6151
R1530 B.n346 B.n345 10.6151
R1531 B.n346 B.n219 10.6151
R1532 B.n350 B.n219 10.6151
R1533 B.n351 B.n350 10.6151
R1534 B.n352 B.n351 10.6151
R1535 B.n352 B.n217 10.6151
R1536 B.n356 B.n217 10.6151
R1537 B.n357 B.n356 10.6151
R1538 B.n358 B.n357 10.6151
R1539 B.n358 B.n215 10.6151
R1540 B.n362 B.n215 10.6151
R1541 B.n363 B.n362 10.6151
R1542 B.n364 B.n363 10.6151
R1543 B.n364 B.n213 10.6151
R1544 B.n368 B.n213 10.6151
R1545 B.n369 B.n368 10.6151
R1546 B.n370 B.n369 10.6151
R1547 B.n370 B.n211 10.6151
R1548 B.n374 B.n211 10.6151
R1549 B.n375 B.n374 10.6151
R1550 B.n376 B.n375 10.6151
R1551 B.n376 B.n209 10.6151
R1552 B.n380 B.n209 10.6151
R1553 B.n381 B.n380 10.6151
R1554 B.n382 B.n381 10.6151
R1555 B.n382 B.n207 10.6151
R1556 B.n386 B.n207 10.6151
R1557 B.n387 B.n386 10.6151
R1558 B.n388 B.n387 10.6151
R1559 B.n388 B.n205 10.6151
R1560 B.n392 B.n205 10.6151
R1561 B.n393 B.n392 10.6151
R1562 B.n394 B.n393 10.6151
R1563 B.n394 B.n203 10.6151
R1564 B.n398 B.n203 10.6151
R1565 B.n399 B.n398 10.6151
R1566 B.n400 B.n399 10.6151
R1567 B.n400 B.n201 10.6151
R1568 B.n404 B.n201 10.6151
R1569 B.n405 B.n404 10.6151
R1570 B.n406 B.n405 10.6151
R1571 B.n406 B.n199 10.6151
R1572 B.n410 B.n199 10.6151
R1573 B.n411 B.n410 10.6151
R1574 B.n412 B.n411 10.6151
R1575 B.n412 B.n197 10.6151
R1576 B.n416 B.n197 10.6151
R1577 B.n417 B.n416 10.6151
R1578 B.n418 B.n417 10.6151
R1579 B.n418 B.n195 10.6151
R1580 B.n422 B.n195 10.6151
R1581 B.n425 B.n424 10.6151
R1582 B.n425 B.n191 10.6151
R1583 B.n429 B.n191 10.6151
R1584 B.n430 B.n429 10.6151
R1585 B.n431 B.n430 10.6151
R1586 B.n431 B.n189 10.6151
R1587 B.n435 B.n189 10.6151
R1588 B.n436 B.n435 10.6151
R1589 B.n437 B.n436 10.6151
R1590 B.n441 B.n440 10.6151
R1591 B.n442 B.n441 10.6151
R1592 B.n442 B.n183 10.6151
R1593 B.n446 B.n183 10.6151
R1594 B.n447 B.n446 10.6151
R1595 B.n448 B.n447 10.6151
R1596 B.n448 B.n181 10.6151
R1597 B.n452 B.n181 10.6151
R1598 B.n453 B.n452 10.6151
R1599 B.n454 B.n453 10.6151
R1600 B.n454 B.n179 10.6151
R1601 B.n458 B.n179 10.6151
R1602 B.n459 B.n458 10.6151
R1603 B.n460 B.n459 10.6151
R1604 B.n460 B.n177 10.6151
R1605 B.n464 B.n177 10.6151
R1606 B.n465 B.n464 10.6151
R1607 B.n466 B.n465 10.6151
R1608 B.n466 B.n175 10.6151
R1609 B.n470 B.n175 10.6151
R1610 B.n471 B.n470 10.6151
R1611 B.n472 B.n471 10.6151
R1612 B.n472 B.n173 10.6151
R1613 B.n476 B.n173 10.6151
R1614 B.n477 B.n476 10.6151
R1615 B.n478 B.n477 10.6151
R1616 B.n478 B.n171 10.6151
R1617 B.n482 B.n171 10.6151
R1618 B.n483 B.n482 10.6151
R1619 B.n484 B.n483 10.6151
R1620 B.n484 B.n169 10.6151
R1621 B.n488 B.n169 10.6151
R1622 B.n489 B.n488 10.6151
R1623 B.n490 B.n489 10.6151
R1624 B.n490 B.n167 10.6151
R1625 B.n494 B.n167 10.6151
R1626 B.n495 B.n494 10.6151
R1627 B.n496 B.n495 10.6151
R1628 B.n496 B.n165 10.6151
R1629 B.n500 B.n165 10.6151
R1630 B.n501 B.n500 10.6151
R1631 B.n502 B.n501 10.6151
R1632 B.n502 B.n163 10.6151
R1633 B.n506 B.n163 10.6151
R1634 B.n507 B.n506 10.6151
R1635 B.n508 B.n507 10.6151
R1636 B.n508 B.n161 10.6151
R1637 B.n512 B.n161 10.6151
R1638 B.n513 B.n512 10.6151
R1639 B.n514 B.n513 10.6151
R1640 B.n514 B.n159 10.6151
R1641 B.n518 B.n159 10.6151
R1642 B.n340 B.n221 10.6151
R1643 B.n340 B.n339 10.6151
R1644 B.n339 B.n338 10.6151
R1645 B.n338 B.n223 10.6151
R1646 B.n334 B.n223 10.6151
R1647 B.n334 B.n333 10.6151
R1648 B.n333 B.n332 10.6151
R1649 B.n332 B.n225 10.6151
R1650 B.n328 B.n225 10.6151
R1651 B.n328 B.n327 10.6151
R1652 B.n327 B.n326 10.6151
R1653 B.n326 B.n227 10.6151
R1654 B.n322 B.n227 10.6151
R1655 B.n322 B.n321 10.6151
R1656 B.n321 B.n320 10.6151
R1657 B.n320 B.n229 10.6151
R1658 B.n316 B.n229 10.6151
R1659 B.n316 B.n315 10.6151
R1660 B.n315 B.n314 10.6151
R1661 B.n314 B.n231 10.6151
R1662 B.n310 B.n231 10.6151
R1663 B.n310 B.n309 10.6151
R1664 B.n309 B.n308 10.6151
R1665 B.n308 B.n233 10.6151
R1666 B.n304 B.n233 10.6151
R1667 B.n304 B.n303 10.6151
R1668 B.n303 B.n302 10.6151
R1669 B.n302 B.n235 10.6151
R1670 B.n298 B.n235 10.6151
R1671 B.n298 B.n297 10.6151
R1672 B.n297 B.n296 10.6151
R1673 B.n296 B.n237 10.6151
R1674 B.n292 B.n237 10.6151
R1675 B.n292 B.n291 10.6151
R1676 B.n291 B.n290 10.6151
R1677 B.n290 B.n239 10.6151
R1678 B.n286 B.n239 10.6151
R1679 B.n286 B.n285 10.6151
R1680 B.n285 B.n284 10.6151
R1681 B.n284 B.n241 10.6151
R1682 B.n280 B.n241 10.6151
R1683 B.n280 B.n279 10.6151
R1684 B.n279 B.n278 10.6151
R1685 B.n278 B.n243 10.6151
R1686 B.n274 B.n243 10.6151
R1687 B.n274 B.n273 10.6151
R1688 B.n273 B.n272 10.6151
R1689 B.n272 B.n245 10.6151
R1690 B.n268 B.n245 10.6151
R1691 B.n268 B.n267 10.6151
R1692 B.n267 B.n266 10.6151
R1693 B.n266 B.n247 10.6151
R1694 B.n262 B.n247 10.6151
R1695 B.n262 B.n261 10.6151
R1696 B.n261 B.n260 10.6151
R1697 B.n260 B.n249 10.6151
R1698 B.n256 B.n249 10.6151
R1699 B.n256 B.n255 10.6151
R1700 B.n255 B.n254 10.6151
R1701 B.n254 B.n251 10.6151
R1702 B.n251 B.n0 10.6151
R1703 B.n971 B.n1 10.6151
R1704 B.n971 B.n970 10.6151
R1705 B.n970 B.n969 10.6151
R1706 B.n969 B.n4 10.6151
R1707 B.n965 B.n4 10.6151
R1708 B.n965 B.n964 10.6151
R1709 B.n964 B.n963 10.6151
R1710 B.n963 B.n6 10.6151
R1711 B.n959 B.n6 10.6151
R1712 B.n959 B.n958 10.6151
R1713 B.n958 B.n957 10.6151
R1714 B.n957 B.n8 10.6151
R1715 B.n953 B.n8 10.6151
R1716 B.n953 B.n952 10.6151
R1717 B.n952 B.n951 10.6151
R1718 B.n951 B.n10 10.6151
R1719 B.n947 B.n10 10.6151
R1720 B.n947 B.n946 10.6151
R1721 B.n946 B.n945 10.6151
R1722 B.n945 B.n12 10.6151
R1723 B.n941 B.n12 10.6151
R1724 B.n941 B.n940 10.6151
R1725 B.n940 B.n939 10.6151
R1726 B.n939 B.n14 10.6151
R1727 B.n935 B.n14 10.6151
R1728 B.n935 B.n934 10.6151
R1729 B.n934 B.n933 10.6151
R1730 B.n933 B.n16 10.6151
R1731 B.n929 B.n16 10.6151
R1732 B.n929 B.n928 10.6151
R1733 B.n928 B.n927 10.6151
R1734 B.n927 B.n18 10.6151
R1735 B.n923 B.n18 10.6151
R1736 B.n923 B.n922 10.6151
R1737 B.n922 B.n921 10.6151
R1738 B.n921 B.n20 10.6151
R1739 B.n917 B.n20 10.6151
R1740 B.n917 B.n916 10.6151
R1741 B.n916 B.n915 10.6151
R1742 B.n915 B.n22 10.6151
R1743 B.n911 B.n22 10.6151
R1744 B.n911 B.n910 10.6151
R1745 B.n910 B.n909 10.6151
R1746 B.n909 B.n24 10.6151
R1747 B.n905 B.n24 10.6151
R1748 B.n905 B.n904 10.6151
R1749 B.n904 B.n903 10.6151
R1750 B.n903 B.n26 10.6151
R1751 B.n899 B.n26 10.6151
R1752 B.n899 B.n898 10.6151
R1753 B.n898 B.n897 10.6151
R1754 B.n897 B.n28 10.6151
R1755 B.n893 B.n28 10.6151
R1756 B.n893 B.n892 10.6151
R1757 B.n892 B.n891 10.6151
R1758 B.n891 B.n30 10.6151
R1759 B.n887 B.n30 10.6151
R1760 B.n887 B.n886 10.6151
R1761 B.n886 B.n885 10.6151
R1762 B.n885 B.n32 10.6151
R1763 B.n881 B.n32 10.6151
R1764 B.n802 B.n801 9.36635
R1765 B.n784 B.n70 9.36635
R1766 B.n423 B.n422 9.36635
R1767 B.n440 B.n187 9.36635
R1768 B.n975 B.n0 2.81026
R1769 B.n975 B.n1 2.81026
R1770 B.n801 B.n800 1.24928
R1771 B.n70 B.n66 1.24928
R1772 B.n424 B.n423 1.24928
R1773 B.n437 B.n187 1.24928
C0 VDD2 VN 11.8829f
C1 VDD1 VDD2 2.14903f
C2 VDD2 B 2.09291f
C3 VDD2 VP 0.59617f
C4 VDD2 w_n4620_n4150# 2.43497f
C5 VN VTAIL 12.334599f
C6 VDD1 VTAIL 9.49239f
C7 VTAIL B 6.61975f
C8 VP VTAIL 12.348701f
C9 VDD1 VN 0.152913f
C10 VN B 1.43875f
C11 w_n4620_n4150# VTAIL 5.13769f
C12 VP VN 9.27046f
C13 VDD1 B 1.97423f
C14 VDD1 VP 12.324401f
C15 VP B 2.45157f
C16 VN w_n4620_n4150# 9.68204f
C17 VDD1 w_n4620_n4150# 2.29006f
C18 w_n4620_n4150# B 12.3137f
C19 VP w_n4620_n4150# 10.2839f
C20 VDD2 VTAIL 9.55164f
C21 VDD2 VSUBS 2.38442f
C22 VDD1 VSUBS 3.05292f
C23 VTAIL VSUBS 1.633521f
C24 VN VSUBS 7.82802f
C25 VP VSUBS 4.469206f
C26 B VSUBS 6.137279f
C27 w_n4620_n4150# VSUBS 0.234899p
C28 B.n0 VSUBS 0.00462f
C29 B.n1 VSUBS 0.00462f
C30 B.n2 VSUBS 0.007307f
C31 B.n3 VSUBS 0.007307f
C32 B.n4 VSUBS 0.007307f
C33 B.n5 VSUBS 0.007307f
C34 B.n6 VSUBS 0.007307f
C35 B.n7 VSUBS 0.007307f
C36 B.n8 VSUBS 0.007307f
C37 B.n9 VSUBS 0.007307f
C38 B.n10 VSUBS 0.007307f
C39 B.n11 VSUBS 0.007307f
C40 B.n12 VSUBS 0.007307f
C41 B.n13 VSUBS 0.007307f
C42 B.n14 VSUBS 0.007307f
C43 B.n15 VSUBS 0.007307f
C44 B.n16 VSUBS 0.007307f
C45 B.n17 VSUBS 0.007307f
C46 B.n18 VSUBS 0.007307f
C47 B.n19 VSUBS 0.007307f
C48 B.n20 VSUBS 0.007307f
C49 B.n21 VSUBS 0.007307f
C50 B.n22 VSUBS 0.007307f
C51 B.n23 VSUBS 0.007307f
C52 B.n24 VSUBS 0.007307f
C53 B.n25 VSUBS 0.007307f
C54 B.n26 VSUBS 0.007307f
C55 B.n27 VSUBS 0.007307f
C56 B.n28 VSUBS 0.007307f
C57 B.n29 VSUBS 0.007307f
C58 B.n30 VSUBS 0.007307f
C59 B.n31 VSUBS 0.007307f
C60 B.n32 VSUBS 0.007307f
C61 B.n33 VSUBS 0.016268f
C62 B.n34 VSUBS 0.007307f
C63 B.n35 VSUBS 0.007307f
C64 B.n36 VSUBS 0.007307f
C65 B.n37 VSUBS 0.007307f
C66 B.n38 VSUBS 0.007307f
C67 B.n39 VSUBS 0.007307f
C68 B.n40 VSUBS 0.007307f
C69 B.n41 VSUBS 0.007307f
C70 B.n42 VSUBS 0.007307f
C71 B.n43 VSUBS 0.007307f
C72 B.n44 VSUBS 0.007307f
C73 B.n45 VSUBS 0.007307f
C74 B.n46 VSUBS 0.007307f
C75 B.n47 VSUBS 0.007307f
C76 B.n48 VSUBS 0.007307f
C77 B.n49 VSUBS 0.007307f
C78 B.n50 VSUBS 0.007307f
C79 B.n51 VSUBS 0.007307f
C80 B.n52 VSUBS 0.007307f
C81 B.n53 VSUBS 0.007307f
C82 B.n54 VSUBS 0.007307f
C83 B.n55 VSUBS 0.007307f
C84 B.n56 VSUBS 0.007307f
C85 B.n57 VSUBS 0.007307f
C86 B.n58 VSUBS 0.007307f
C87 B.n59 VSUBS 0.007307f
C88 B.t5 VSUBS 0.55554f
C89 B.t4 VSUBS 0.581867f
C90 B.t3 VSUBS 2.50889f
C91 B.n60 VSUBS 0.338564f
C92 B.n61 VSUBS 0.078275f
C93 B.n62 VSUBS 0.007307f
C94 B.n63 VSUBS 0.007307f
C95 B.n64 VSUBS 0.007307f
C96 B.n65 VSUBS 0.007307f
C97 B.n66 VSUBS 0.004083f
C98 B.n67 VSUBS 0.007307f
C99 B.t8 VSUBS 0.555523f
C100 B.t7 VSUBS 0.581854f
C101 B.t6 VSUBS 2.50889f
C102 B.n68 VSUBS 0.338577f
C103 B.n69 VSUBS 0.078291f
C104 B.n70 VSUBS 0.016929f
C105 B.n71 VSUBS 0.007307f
C106 B.n72 VSUBS 0.007307f
C107 B.n73 VSUBS 0.007307f
C108 B.n74 VSUBS 0.007307f
C109 B.n75 VSUBS 0.007307f
C110 B.n76 VSUBS 0.007307f
C111 B.n77 VSUBS 0.007307f
C112 B.n78 VSUBS 0.007307f
C113 B.n79 VSUBS 0.007307f
C114 B.n80 VSUBS 0.007307f
C115 B.n81 VSUBS 0.007307f
C116 B.n82 VSUBS 0.007307f
C117 B.n83 VSUBS 0.007307f
C118 B.n84 VSUBS 0.007307f
C119 B.n85 VSUBS 0.007307f
C120 B.n86 VSUBS 0.007307f
C121 B.n87 VSUBS 0.007307f
C122 B.n88 VSUBS 0.007307f
C123 B.n89 VSUBS 0.007307f
C124 B.n90 VSUBS 0.007307f
C125 B.n91 VSUBS 0.007307f
C126 B.n92 VSUBS 0.007307f
C127 B.n93 VSUBS 0.007307f
C128 B.n94 VSUBS 0.007307f
C129 B.n95 VSUBS 0.007307f
C130 B.n96 VSUBS 0.015538f
C131 B.n97 VSUBS 0.007307f
C132 B.n98 VSUBS 0.007307f
C133 B.n99 VSUBS 0.007307f
C134 B.n100 VSUBS 0.007307f
C135 B.n101 VSUBS 0.007307f
C136 B.n102 VSUBS 0.007307f
C137 B.n103 VSUBS 0.007307f
C138 B.n104 VSUBS 0.007307f
C139 B.n105 VSUBS 0.007307f
C140 B.n106 VSUBS 0.007307f
C141 B.n107 VSUBS 0.007307f
C142 B.n108 VSUBS 0.007307f
C143 B.n109 VSUBS 0.007307f
C144 B.n110 VSUBS 0.007307f
C145 B.n111 VSUBS 0.007307f
C146 B.n112 VSUBS 0.007307f
C147 B.n113 VSUBS 0.007307f
C148 B.n114 VSUBS 0.007307f
C149 B.n115 VSUBS 0.007307f
C150 B.n116 VSUBS 0.007307f
C151 B.n117 VSUBS 0.007307f
C152 B.n118 VSUBS 0.007307f
C153 B.n119 VSUBS 0.007307f
C154 B.n120 VSUBS 0.007307f
C155 B.n121 VSUBS 0.007307f
C156 B.n122 VSUBS 0.007307f
C157 B.n123 VSUBS 0.007307f
C158 B.n124 VSUBS 0.007307f
C159 B.n125 VSUBS 0.007307f
C160 B.n126 VSUBS 0.007307f
C161 B.n127 VSUBS 0.007307f
C162 B.n128 VSUBS 0.007307f
C163 B.n129 VSUBS 0.007307f
C164 B.n130 VSUBS 0.007307f
C165 B.n131 VSUBS 0.007307f
C166 B.n132 VSUBS 0.007307f
C167 B.n133 VSUBS 0.007307f
C168 B.n134 VSUBS 0.007307f
C169 B.n135 VSUBS 0.007307f
C170 B.n136 VSUBS 0.007307f
C171 B.n137 VSUBS 0.007307f
C172 B.n138 VSUBS 0.007307f
C173 B.n139 VSUBS 0.007307f
C174 B.n140 VSUBS 0.007307f
C175 B.n141 VSUBS 0.007307f
C176 B.n142 VSUBS 0.007307f
C177 B.n143 VSUBS 0.007307f
C178 B.n144 VSUBS 0.007307f
C179 B.n145 VSUBS 0.007307f
C180 B.n146 VSUBS 0.007307f
C181 B.n147 VSUBS 0.007307f
C182 B.n148 VSUBS 0.007307f
C183 B.n149 VSUBS 0.007307f
C184 B.n150 VSUBS 0.007307f
C185 B.n151 VSUBS 0.007307f
C186 B.n152 VSUBS 0.007307f
C187 B.n153 VSUBS 0.007307f
C188 B.n154 VSUBS 0.007307f
C189 B.n155 VSUBS 0.007307f
C190 B.n156 VSUBS 0.007307f
C191 B.n157 VSUBS 0.007307f
C192 B.n158 VSUBS 0.015538f
C193 B.n159 VSUBS 0.007307f
C194 B.n160 VSUBS 0.007307f
C195 B.n161 VSUBS 0.007307f
C196 B.n162 VSUBS 0.007307f
C197 B.n163 VSUBS 0.007307f
C198 B.n164 VSUBS 0.007307f
C199 B.n165 VSUBS 0.007307f
C200 B.n166 VSUBS 0.007307f
C201 B.n167 VSUBS 0.007307f
C202 B.n168 VSUBS 0.007307f
C203 B.n169 VSUBS 0.007307f
C204 B.n170 VSUBS 0.007307f
C205 B.n171 VSUBS 0.007307f
C206 B.n172 VSUBS 0.007307f
C207 B.n173 VSUBS 0.007307f
C208 B.n174 VSUBS 0.007307f
C209 B.n175 VSUBS 0.007307f
C210 B.n176 VSUBS 0.007307f
C211 B.n177 VSUBS 0.007307f
C212 B.n178 VSUBS 0.007307f
C213 B.n179 VSUBS 0.007307f
C214 B.n180 VSUBS 0.007307f
C215 B.n181 VSUBS 0.007307f
C216 B.n182 VSUBS 0.007307f
C217 B.n183 VSUBS 0.007307f
C218 B.n184 VSUBS 0.007307f
C219 B.t1 VSUBS 0.555523f
C220 B.t2 VSUBS 0.581854f
C221 B.t0 VSUBS 2.50889f
C222 B.n185 VSUBS 0.338577f
C223 B.n186 VSUBS 0.078291f
C224 B.n187 VSUBS 0.016929f
C225 B.n188 VSUBS 0.007307f
C226 B.n189 VSUBS 0.007307f
C227 B.n190 VSUBS 0.007307f
C228 B.n191 VSUBS 0.007307f
C229 B.n192 VSUBS 0.007307f
C230 B.t10 VSUBS 0.55554f
C231 B.t11 VSUBS 0.581867f
C232 B.t9 VSUBS 2.50889f
C233 B.n193 VSUBS 0.338564f
C234 B.n194 VSUBS 0.078275f
C235 B.n195 VSUBS 0.007307f
C236 B.n196 VSUBS 0.007307f
C237 B.n197 VSUBS 0.007307f
C238 B.n198 VSUBS 0.007307f
C239 B.n199 VSUBS 0.007307f
C240 B.n200 VSUBS 0.007307f
C241 B.n201 VSUBS 0.007307f
C242 B.n202 VSUBS 0.007307f
C243 B.n203 VSUBS 0.007307f
C244 B.n204 VSUBS 0.007307f
C245 B.n205 VSUBS 0.007307f
C246 B.n206 VSUBS 0.007307f
C247 B.n207 VSUBS 0.007307f
C248 B.n208 VSUBS 0.007307f
C249 B.n209 VSUBS 0.007307f
C250 B.n210 VSUBS 0.007307f
C251 B.n211 VSUBS 0.007307f
C252 B.n212 VSUBS 0.007307f
C253 B.n213 VSUBS 0.007307f
C254 B.n214 VSUBS 0.007307f
C255 B.n215 VSUBS 0.007307f
C256 B.n216 VSUBS 0.007307f
C257 B.n217 VSUBS 0.007307f
C258 B.n218 VSUBS 0.007307f
C259 B.n219 VSUBS 0.007307f
C260 B.n220 VSUBS 0.007307f
C261 B.n221 VSUBS 0.015538f
C262 B.n222 VSUBS 0.007307f
C263 B.n223 VSUBS 0.007307f
C264 B.n224 VSUBS 0.007307f
C265 B.n225 VSUBS 0.007307f
C266 B.n226 VSUBS 0.007307f
C267 B.n227 VSUBS 0.007307f
C268 B.n228 VSUBS 0.007307f
C269 B.n229 VSUBS 0.007307f
C270 B.n230 VSUBS 0.007307f
C271 B.n231 VSUBS 0.007307f
C272 B.n232 VSUBS 0.007307f
C273 B.n233 VSUBS 0.007307f
C274 B.n234 VSUBS 0.007307f
C275 B.n235 VSUBS 0.007307f
C276 B.n236 VSUBS 0.007307f
C277 B.n237 VSUBS 0.007307f
C278 B.n238 VSUBS 0.007307f
C279 B.n239 VSUBS 0.007307f
C280 B.n240 VSUBS 0.007307f
C281 B.n241 VSUBS 0.007307f
C282 B.n242 VSUBS 0.007307f
C283 B.n243 VSUBS 0.007307f
C284 B.n244 VSUBS 0.007307f
C285 B.n245 VSUBS 0.007307f
C286 B.n246 VSUBS 0.007307f
C287 B.n247 VSUBS 0.007307f
C288 B.n248 VSUBS 0.007307f
C289 B.n249 VSUBS 0.007307f
C290 B.n250 VSUBS 0.007307f
C291 B.n251 VSUBS 0.007307f
C292 B.n252 VSUBS 0.007307f
C293 B.n253 VSUBS 0.007307f
C294 B.n254 VSUBS 0.007307f
C295 B.n255 VSUBS 0.007307f
C296 B.n256 VSUBS 0.007307f
C297 B.n257 VSUBS 0.007307f
C298 B.n258 VSUBS 0.007307f
C299 B.n259 VSUBS 0.007307f
C300 B.n260 VSUBS 0.007307f
C301 B.n261 VSUBS 0.007307f
C302 B.n262 VSUBS 0.007307f
C303 B.n263 VSUBS 0.007307f
C304 B.n264 VSUBS 0.007307f
C305 B.n265 VSUBS 0.007307f
C306 B.n266 VSUBS 0.007307f
C307 B.n267 VSUBS 0.007307f
C308 B.n268 VSUBS 0.007307f
C309 B.n269 VSUBS 0.007307f
C310 B.n270 VSUBS 0.007307f
C311 B.n271 VSUBS 0.007307f
C312 B.n272 VSUBS 0.007307f
C313 B.n273 VSUBS 0.007307f
C314 B.n274 VSUBS 0.007307f
C315 B.n275 VSUBS 0.007307f
C316 B.n276 VSUBS 0.007307f
C317 B.n277 VSUBS 0.007307f
C318 B.n278 VSUBS 0.007307f
C319 B.n279 VSUBS 0.007307f
C320 B.n280 VSUBS 0.007307f
C321 B.n281 VSUBS 0.007307f
C322 B.n282 VSUBS 0.007307f
C323 B.n283 VSUBS 0.007307f
C324 B.n284 VSUBS 0.007307f
C325 B.n285 VSUBS 0.007307f
C326 B.n286 VSUBS 0.007307f
C327 B.n287 VSUBS 0.007307f
C328 B.n288 VSUBS 0.007307f
C329 B.n289 VSUBS 0.007307f
C330 B.n290 VSUBS 0.007307f
C331 B.n291 VSUBS 0.007307f
C332 B.n292 VSUBS 0.007307f
C333 B.n293 VSUBS 0.007307f
C334 B.n294 VSUBS 0.007307f
C335 B.n295 VSUBS 0.007307f
C336 B.n296 VSUBS 0.007307f
C337 B.n297 VSUBS 0.007307f
C338 B.n298 VSUBS 0.007307f
C339 B.n299 VSUBS 0.007307f
C340 B.n300 VSUBS 0.007307f
C341 B.n301 VSUBS 0.007307f
C342 B.n302 VSUBS 0.007307f
C343 B.n303 VSUBS 0.007307f
C344 B.n304 VSUBS 0.007307f
C345 B.n305 VSUBS 0.007307f
C346 B.n306 VSUBS 0.007307f
C347 B.n307 VSUBS 0.007307f
C348 B.n308 VSUBS 0.007307f
C349 B.n309 VSUBS 0.007307f
C350 B.n310 VSUBS 0.007307f
C351 B.n311 VSUBS 0.007307f
C352 B.n312 VSUBS 0.007307f
C353 B.n313 VSUBS 0.007307f
C354 B.n314 VSUBS 0.007307f
C355 B.n315 VSUBS 0.007307f
C356 B.n316 VSUBS 0.007307f
C357 B.n317 VSUBS 0.007307f
C358 B.n318 VSUBS 0.007307f
C359 B.n319 VSUBS 0.007307f
C360 B.n320 VSUBS 0.007307f
C361 B.n321 VSUBS 0.007307f
C362 B.n322 VSUBS 0.007307f
C363 B.n323 VSUBS 0.007307f
C364 B.n324 VSUBS 0.007307f
C365 B.n325 VSUBS 0.007307f
C366 B.n326 VSUBS 0.007307f
C367 B.n327 VSUBS 0.007307f
C368 B.n328 VSUBS 0.007307f
C369 B.n329 VSUBS 0.007307f
C370 B.n330 VSUBS 0.007307f
C371 B.n331 VSUBS 0.007307f
C372 B.n332 VSUBS 0.007307f
C373 B.n333 VSUBS 0.007307f
C374 B.n334 VSUBS 0.007307f
C375 B.n335 VSUBS 0.007307f
C376 B.n336 VSUBS 0.007307f
C377 B.n337 VSUBS 0.007307f
C378 B.n338 VSUBS 0.007307f
C379 B.n339 VSUBS 0.007307f
C380 B.n340 VSUBS 0.007307f
C381 B.n341 VSUBS 0.007307f
C382 B.n342 VSUBS 0.015538f
C383 B.n343 VSUBS 0.016268f
C384 B.n344 VSUBS 0.016268f
C385 B.n345 VSUBS 0.007307f
C386 B.n346 VSUBS 0.007307f
C387 B.n347 VSUBS 0.007307f
C388 B.n348 VSUBS 0.007307f
C389 B.n349 VSUBS 0.007307f
C390 B.n350 VSUBS 0.007307f
C391 B.n351 VSUBS 0.007307f
C392 B.n352 VSUBS 0.007307f
C393 B.n353 VSUBS 0.007307f
C394 B.n354 VSUBS 0.007307f
C395 B.n355 VSUBS 0.007307f
C396 B.n356 VSUBS 0.007307f
C397 B.n357 VSUBS 0.007307f
C398 B.n358 VSUBS 0.007307f
C399 B.n359 VSUBS 0.007307f
C400 B.n360 VSUBS 0.007307f
C401 B.n361 VSUBS 0.007307f
C402 B.n362 VSUBS 0.007307f
C403 B.n363 VSUBS 0.007307f
C404 B.n364 VSUBS 0.007307f
C405 B.n365 VSUBS 0.007307f
C406 B.n366 VSUBS 0.007307f
C407 B.n367 VSUBS 0.007307f
C408 B.n368 VSUBS 0.007307f
C409 B.n369 VSUBS 0.007307f
C410 B.n370 VSUBS 0.007307f
C411 B.n371 VSUBS 0.007307f
C412 B.n372 VSUBS 0.007307f
C413 B.n373 VSUBS 0.007307f
C414 B.n374 VSUBS 0.007307f
C415 B.n375 VSUBS 0.007307f
C416 B.n376 VSUBS 0.007307f
C417 B.n377 VSUBS 0.007307f
C418 B.n378 VSUBS 0.007307f
C419 B.n379 VSUBS 0.007307f
C420 B.n380 VSUBS 0.007307f
C421 B.n381 VSUBS 0.007307f
C422 B.n382 VSUBS 0.007307f
C423 B.n383 VSUBS 0.007307f
C424 B.n384 VSUBS 0.007307f
C425 B.n385 VSUBS 0.007307f
C426 B.n386 VSUBS 0.007307f
C427 B.n387 VSUBS 0.007307f
C428 B.n388 VSUBS 0.007307f
C429 B.n389 VSUBS 0.007307f
C430 B.n390 VSUBS 0.007307f
C431 B.n391 VSUBS 0.007307f
C432 B.n392 VSUBS 0.007307f
C433 B.n393 VSUBS 0.007307f
C434 B.n394 VSUBS 0.007307f
C435 B.n395 VSUBS 0.007307f
C436 B.n396 VSUBS 0.007307f
C437 B.n397 VSUBS 0.007307f
C438 B.n398 VSUBS 0.007307f
C439 B.n399 VSUBS 0.007307f
C440 B.n400 VSUBS 0.007307f
C441 B.n401 VSUBS 0.007307f
C442 B.n402 VSUBS 0.007307f
C443 B.n403 VSUBS 0.007307f
C444 B.n404 VSUBS 0.007307f
C445 B.n405 VSUBS 0.007307f
C446 B.n406 VSUBS 0.007307f
C447 B.n407 VSUBS 0.007307f
C448 B.n408 VSUBS 0.007307f
C449 B.n409 VSUBS 0.007307f
C450 B.n410 VSUBS 0.007307f
C451 B.n411 VSUBS 0.007307f
C452 B.n412 VSUBS 0.007307f
C453 B.n413 VSUBS 0.007307f
C454 B.n414 VSUBS 0.007307f
C455 B.n415 VSUBS 0.007307f
C456 B.n416 VSUBS 0.007307f
C457 B.n417 VSUBS 0.007307f
C458 B.n418 VSUBS 0.007307f
C459 B.n419 VSUBS 0.007307f
C460 B.n420 VSUBS 0.007307f
C461 B.n421 VSUBS 0.007307f
C462 B.n422 VSUBS 0.006877f
C463 B.n423 VSUBS 0.016929f
C464 B.n424 VSUBS 0.004083f
C465 B.n425 VSUBS 0.007307f
C466 B.n426 VSUBS 0.007307f
C467 B.n427 VSUBS 0.007307f
C468 B.n428 VSUBS 0.007307f
C469 B.n429 VSUBS 0.007307f
C470 B.n430 VSUBS 0.007307f
C471 B.n431 VSUBS 0.007307f
C472 B.n432 VSUBS 0.007307f
C473 B.n433 VSUBS 0.007307f
C474 B.n434 VSUBS 0.007307f
C475 B.n435 VSUBS 0.007307f
C476 B.n436 VSUBS 0.007307f
C477 B.n437 VSUBS 0.004083f
C478 B.n438 VSUBS 0.007307f
C479 B.n439 VSUBS 0.007307f
C480 B.n440 VSUBS 0.006877f
C481 B.n441 VSUBS 0.007307f
C482 B.n442 VSUBS 0.007307f
C483 B.n443 VSUBS 0.007307f
C484 B.n444 VSUBS 0.007307f
C485 B.n445 VSUBS 0.007307f
C486 B.n446 VSUBS 0.007307f
C487 B.n447 VSUBS 0.007307f
C488 B.n448 VSUBS 0.007307f
C489 B.n449 VSUBS 0.007307f
C490 B.n450 VSUBS 0.007307f
C491 B.n451 VSUBS 0.007307f
C492 B.n452 VSUBS 0.007307f
C493 B.n453 VSUBS 0.007307f
C494 B.n454 VSUBS 0.007307f
C495 B.n455 VSUBS 0.007307f
C496 B.n456 VSUBS 0.007307f
C497 B.n457 VSUBS 0.007307f
C498 B.n458 VSUBS 0.007307f
C499 B.n459 VSUBS 0.007307f
C500 B.n460 VSUBS 0.007307f
C501 B.n461 VSUBS 0.007307f
C502 B.n462 VSUBS 0.007307f
C503 B.n463 VSUBS 0.007307f
C504 B.n464 VSUBS 0.007307f
C505 B.n465 VSUBS 0.007307f
C506 B.n466 VSUBS 0.007307f
C507 B.n467 VSUBS 0.007307f
C508 B.n468 VSUBS 0.007307f
C509 B.n469 VSUBS 0.007307f
C510 B.n470 VSUBS 0.007307f
C511 B.n471 VSUBS 0.007307f
C512 B.n472 VSUBS 0.007307f
C513 B.n473 VSUBS 0.007307f
C514 B.n474 VSUBS 0.007307f
C515 B.n475 VSUBS 0.007307f
C516 B.n476 VSUBS 0.007307f
C517 B.n477 VSUBS 0.007307f
C518 B.n478 VSUBS 0.007307f
C519 B.n479 VSUBS 0.007307f
C520 B.n480 VSUBS 0.007307f
C521 B.n481 VSUBS 0.007307f
C522 B.n482 VSUBS 0.007307f
C523 B.n483 VSUBS 0.007307f
C524 B.n484 VSUBS 0.007307f
C525 B.n485 VSUBS 0.007307f
C526 B.n486 VSUBS 0.007307f
C527 B.n487 VSUBS 0.007307f
C528 B.n488 VSUBS 0.007307f
C529 B.n489 VSUBS 0.007307f
C530 B.n490 VSUBS 0.007307f
C531 B.n491 VSUBS 0.007307f
C532 B.n492 VSUBS 0.007307f
C533 B.n493 VSUBS 0.007307f
C534 B.n494 VSUBS 0.007307f
C535 B.n495 VSUBS 0.007307f
C536 B.n496 VSUBS 0.007307f
C537 B.n497 VSUBS 0.007307f
C538 B.n498 VSUBS 0.007307f
C539 B.n499 VSUBS 0.007307f
C540 B.n500 VSUBS 0.007307f
C541 B.n501 VSUBS 0.007307f
C542 B.n502 VSUBS 0.007307f
C543 B.n503 VSUBS 0.007307f
C544 B.n504 VSUBS 0.007307f
C545 B.n505 VSUBS 0.007307f
C546 B.n506 VSUBS 0.007307f
C547 B.n507 VSUBS 0.007307f
C548 B.n508 VSUBS 0.007307f
C549 B.n509 VSUBS 0.007307f
C550 B.n510 VSUBS 0.007307f
C551 B.n511 VSUBS 0.007307f
C552 B.n512 VSUBS 0.007307f
C553 B.n513 VSUBS 0.007307f
C554 B.n514 VSUBS 0.007307f
C555 B.n515 VSUBS 0.007307f
C556 B.n516 VSUBS 0.007307f
C557 B.n517 VSUBS 0.016268f
C558 B.n518 VSUBS 0.016268f
C559 B.n519 VSUBS 0.015538f
C560 B.n520 VSUBS 0.007307f
C561 B.n521 VSUBS 0.007307f
C562 B.n522 VSUBS 0.007307f
C563 B.n523 VSUBS 0.007307f
C564 B.n524 VSUBS 0.007307f
C565 B.n525 VSUBS 0.007307f
C566 B.n526 VSUBS 0.007307f
C567 B.n527 VSUBS 0.007307f
C568 B.n528 VSUBS 0.007307f
C569 B.n529 VSUBS 0.007307f
C570 B.n530 VSUBS 0.007307f
C571 B.n531 VSUBS 0.007307f
C572 B.n532 VSUBS 0.007307f
C573 B.n533 VSUBS 0.007307f
C574 B.n534 VSUBS 0.007307f
C575 B.n535 VSUBS 0.007307f
C576 B.n536 VSUBS 0.007307f
C577 B.n537 VSUBS 0.007307f
C578 B.n538 VSUBS 0.007307f
C579 B.n539 VSUBS 0.007307f
C580 B.n540 VSUBS 0.007307f
C581 B.n541 VSUBS 0.007307f
C582 B.n542 VSUBS 0.007307f
C583 B.n543 VSUBS 0.007307f
C584 B.n544 VSUBS 0.007307f
C585 B.n545 VSUBS 0.007307f
C586 B.n546 VSUBS 0.007307f
C587 B.n547 VSUBS 0.007307f
C588 B.n548 VSUBS 0.007307f
C589 B.n549 VSUBS 0.007307f
C590 B.n550 VSUBS 0.007307f
C591 B.n551 VSUBS 0.007307f
C592 B.n552 VSUBS 0.007307f
C593 B.n553 VSUBS 0.007307f
C594 B.n554 VSUBS 0.007307f
C595 B.n555 VSUBS 0.007307f
C596 B.n556 VSUBS 0.007307f
C597 B.n557 VSUBS 0.007307f
C598 B.n558 VSUBS 0.007307f
C599 B.n559 VSUBS 0.007307f
C600 B.n560 VSUBS 0.007307f
C601 B.n561 VSUBS 0.007307f
C602 B.n562 VSUBS 0.007307f
C603 B.n563 VSUBS 0.007307f
C604 B.n564 VSUBS 0.007307f
C605 B.n565 VSUBS 0.007307f
C606 B.n566 VSUBS 0.007307f
C607 B.n567 VSUBS 0.007307f
C608 B.n568 VSUBS 0.007307f
C609 B.n569 VSUBS 0.007307f
C610 B.n570 VSUBS 0.007307f
C611 B.n571 VSUBS 0.007307f
C612 B.n572 VSUBS 0.007307f
C613 B.n573 VSUBS 0.007307f
C614 B.n574 VSUBS 0.007307f
C615 B.n575 VSUBS 0.007307f
C616 B.n576 VSUBS 0.007307f
C617 B.n577 VSUBS 0.007307f
C618 B.n578 VSUBS 0.007307f
C619 B.n579 VSUBS 0.007307f
C620 B.n580 VSUBS 0.007307f
C621 B.n581 VSUBS 0.007307f
C622 B.n582 VSUBS 0.007307f
C623 B.n583 VSUBS 0.007307f
C624 B.n584 VSUBS 0.007307f
C625 B.n585 VSUBS 0.007307f
C626 B.n586 VSUBS 0.007307f
C627 B.n587 VSUBS 0.007307f
C628 B.n588 VSUBS 0.007307f
C629 B.n589 VSUBS 0.007307f
C630 B.n590 VSUBS 0.007307f
C631 B.n591 VSUBS 0.007307f
C632 B.n592 VSUBS 0.007307f
C633 B.n593 VSUBS 0.007307f
C634 B.n594 VSUBS 0.007307f
C635 B.n595 VSUBS 0.007307f
C636 B.n596 VSUBS 0.007307f
C637 B.n597 VSUBS 0.007307f
C638 B.n598 VSUBS 0.007307f
C639 B.n599 VSUBS 0.007307f
C640 B.n600 VSUBS 0.007307f
C641 B.n601 VSUBS 0.007307f
C642 B.n602 VSUBS 0.007307f
C643 B.n603 VSUBS 0.007307f
C644 B.n604 VSUBS 0.007307f
C645 B.n605 VSUBS 0.007307f
C646 B.n606 VSUBS 0.007307f
C647 B.n607 VSUBS 0.007307f
C648 B.n608 VSUBS 0.007307f
C649 B.n609 VSUBS 0.007307f
C650 B.n610 VSUBS 0.007307f
C651 B.n611 VSUBS 0.007307f
C652 B.n612 VSUBS 0.007307f
C653 B.n613 VSUBS 0.007307f
C654 B.n614 VSUBS 0.007307f
C655 B.n615 VSUBS 0.007307f
C656 B.n616 VSUBS 0.007307f
C657 B.n617 VSUBS 0.007307f
C658 B.n618 VSUBS 0.007307f
C659 B.n619 VSUBS 0.007307f
C660 B.n620 VSUBS 0.007307f
C661 B.n621 VSUBS 0.007307f
C662 B.n622 VSUBS 0.007307f
C663 B.n623 VSUBS 0.007307f
C664 B.n624 VSUBS 0.007307f
C665 B.n625 VSUBS 0.007307f
C666 B.n626 VSUBS 0.007307f
C667 B.n627 VSUBS 0.007307f
C668 B.n628 VSUBS 0.007307f
C669 B.n629 VSUBS 0.007307f
C670 B.n630 VSUBS 0.007307f
C671 B.n631 VSUBS 0.007307f
C672 B.n632 VSUBS 0.007307f
C673 B.n633 VSUBS 0.007307f
C674 B.n634 VSUBS 0.007307f
C675 B.n635 VSUBS 0.007307f
C676 B.n636 VSUBS 0.007307f
C677 B.n637 VSUBS 0.007307f
C678 B.n638 VSUBS 0.007307f
C679 B.n639 VSUBS 0.007307f
C680 B.n640 VSUBS 0.007307f
C681 B.n641 VSUBS 0.007307f
C682 B.n642 VSUBS 0.007307f
C683 B.n643 VSUBS 0.007307f
C684 B.n644 VSUBS 0.007307f
C685 B.n645 VSUBS 0.007307f
C686 B.n646 VSUBS 0.007307f
C687 B.n647 VSUBS 0.007307f
C688 B.n648 VSUBS 0.007307f
C689 B.n649 VSUBS 0.007307f
C690 B.n650 VSUBS 0.007307f
C691 B.n651 VSUBS 0.007307f
C692 B.n652 VSUBS 0.007307f
C693 B.n653 VSUBS 0.007307f
C694 B.n654 VSUBS 0.007307f
C695 B.n655 VSUBS 0.007307f
C696 B.n656 VSUBS 0.007307f
C697 B.n657 VSUBS 0.007307f
C698 B.n658 VSUBS 0.007307f
C699 B.n659 VSUBS 0.007307f
C700 B.n660 VSUBS 0.007307f
C701 B.n661 VSUBS 0.007307f
C702 B.n662 VSUBS 0.007307f
C703 B.n663 VSUBS 0.007307f
C704 B.n664 VSUBS 0.007307f
C705 B.n665 VSUBS 0.007307f
C706 B.n666 VSUBS 0.007307f
C707 B.n667 VSUBS 0.007307f
C708 B.n668 VSUBS 0.007307f
C709 B.n669 VSUBS 0.007307f
C710 B.n670 VSUBS 0.007307f
C711 B.n671 VSUBS 0.007307f
C712 B.n672 VSUBS 0.007307f
C713 B.n673 VSUBS 0.007307f
C714 B.n674 VSUBS 0.007307f
C715 B.n675 VSUBS 0.007307f
C716 B.n676 VSUBS 0.007307f
C717 B.n677 VSUBS 0.007307f
C718 B.n678 VSUBS 0.007307f
C719 B.n679 VSUBS 0.007307f
C720 B.n680 VSUBS 0.007307f
C721 B.n681 VSUBS 0.007307f
C722 B.n682 VSUBS 0.007307f
C723 B.n683 VSUBS 0.007307f
C724 B.n684 VSUBS 0.007307f
C725 B.n685 VSUBS 0.007307f
C726 B.n686 VSUBS 0.007307f
C727 B.n687 VSUBS 0.007307f
C728 B.n688 VSUBS 0.007307f
C729 B.n689 VSUBS 0.007307f
C730 B.n690 VSUBS 0.007307f
C731 B.n691 VSUBS 0.007307f
C732 B.n692 VSUBS 0.007307f
C733 B.n693 VSUBS 0.007307f
C734 B.n694 VSUBS 0.007307f
C735 B.n695 VSUBS 0.007307f
C736 B.n696 VSUBS 0.007307f
C737 B.n697 VSUBS 0.007307f
C738 B.n698 VSUBS 0.007307f
C739 B.n699 VSUBS 0.007307f
C740 B.n700 VSUBS 0.007307f
C741 B.n701 VSUBS 0.007307f
C742 B.n702 VSUBS 0.007307f
C743 B.n703 VSUBS 0.007307f
C744 B.n704 VSUBS 0.007307f
C745 B.n705 VSUBS 0.016504f
C746 B.n706 VSUBS 0.015302f
C747 B.n707 VSUBS 0.016268f
C748 B.n708 VSUBS 0.007307f
C749 B.n709 VSUBS 0.007307f
C750 B.n710 VSUBS 0.007307f
C751 B.n711 VSUBS 0.007307f
C752 B.n712 VSUBS 0.007307f
C753 B.n713 VSUBS 0.007307f
C754 B.n714 VSUBS 0.007307f
C755 B.n715 VSUBS 0.007307f
C756 B.n716 VSUBS 0.007307f
C757 B.n717 VSUBS 0.007307f
C758 B.n718 VSUBS 0.007307f
C759 B.n719 VSUBS 0.007307f
C760 B.n720 VSUBS 0.007307f
C761 B.n721 VSUBS 0.007307f
C762 B.n722 VSUBS 0.007307f
C763 B.n723 VSUBS 0.007307f
C764 B.n724 VSUBS 0.007307f
C765 B.n725 VSUBS 0.007307f
C766 B.n726 VSUBS 0.007307f
C767 B.n727 VSUBS 0.007307f
C768 B.n728 VSUBS 0.007307f
C769 B.n729 VSUBS 0.007307f
C770 B.n730 VSUBS 0.007307f
C771 B.n731 VSUBS 0.007307f
C772 B.n732 VSUBS 0.007307f
C773 B.n733 VSUBS 0.007307f
C774 B.n734 VSUBS 0.007307f
C775 B.n735 VSUBS 0.007307f
C776 B.n736 VSUBS 0.007307f
C777 B.n737 VSUBS 0.007307f
C778 B.n738 VSUBS 0.007307f
C779 B.n739 VSUBS 0.007307f
C780 B.n740 VSUBS 0.007307f
C781 B.n741 VSUBS 0.007307f
C782 B.n742 VSUBS 0.007307f
C783 B.n743 VSUBS 0.007307f
C784 B.n744 VSUBS 0.007307f
C785 B.n745 VSUBS 0.007307f
C786 B.n746 VSUBS 0.007307f
C787 B.n747 VSUBS 0.007307f
C788 B.n748 VSUBS 0.007307f
C789 B.n749 VSUBS 0.007307f
C790 B.n750 VSUBS 0.007307f
C791 B.n751 VSUBS 0.007307f
C792 B.n752 VSUBS 0.007307f
C793 B.n753 VSUBS 0.007307f
C794 B.n754 VSUBS 0.007307f
C795 B.n755 VSUBS 0.007307f
C796 B.n756 VSUBS 0.007307f
C797 B.n757 VSUBS 0.007307f
C798 B.n758 VSUBS 0.007307f
C799 B.n759 VSUBS 0.007307f
C800 B.n760 VSUBS 0.007307f
C801 B.n761 VSUBS 0.007307f
C802 B.n762 VSUBS 0.007307f
C803 B.n763 VSUBS 0.007307f
C804 B.n764 VSUBS 0.007307f
C805 B.n765 VSUBS 0.007307f
C806 B.n766 VSUBS 0.007307f
C807 B.n767 VSUBS 0.007307f
C808 B.n768 VSUBS 0.007307f
C809 B.n769 VSUBS 0.007307f
C810 B.n770 VSUBS 0.007307f
C811 B.n771 VSUBS 0.007307f
C812 B.n772 VSUBS 0.007307f
C813 B.n773 VSUBS 0.007307f
C814 B.n774 VSUBS 0.007307f
C815 B.n775 VSUBS 0.007307f
C816 B.n776 VSUBS 0.007307f
C817 B.n777 VSUBS 0.007307f
C818 B.n778 VSUBS 0.007307f
C819 B.n779 VSUBS 0.007307f
C820 B.n780 VSUBS 0.007307f
C821 B.n781 VSUBS 0.007307f
C822 B.n782 VSUBS 0.007307f
C823 B.n783 VSUBS 0.007307f
C824 B.n784 VSUBS 0.006877f
C825 B.n785 VSUBS 0.007307f
C826 B.n786 VSUBS 0.007307f
C827 B.n787 VSUBS 0.007307f
C828 B.n788 VSUBS 0.007307f
C829 B.n789 VSUBS 0.007307f
C830 B.n790 VSUBS 0.007307f
C831 B.n791 VSUBS 0.007307f
C832 B.n792 VSUBS 0.007307f
C833 B.n793 VSUBS 0.007307f
C834 B.n794 VSUBS 0.007307f
C835 B.n795 VSUBS 0.007307f
C836 B.n796 VSUBS 0.007307f
C837 B.n797 VSUBS 0.007307f
C838 B.n798 VSUBS 0.007307f
C839 B.n799 VSUBS 0.007307f
C840 B.n800 VSUBS 0.004083f
C841 B.n801 VSUBS 0.016929f
C842 B.n802 VSUBS 0.006877f
C843 B.n803 VSUBS 0.007307f
C844 B.n804 VSUBS 0.007307f
C845 B.n805 VSUBS 0.007307f
C846 B.n806 VSUBS 0.007307f
C847 B.n807 VSUBS 0.007307f
C848 B.n808 VSUBS 0.007307f
C849 B.n809 VSUBS 0.007307f
C850 B.n810 VSUBS 0.007307f
C851 B.n811 VSUBS 0.007307f
C852 B.n812 VSUBS 0.007307f
C853 B.n813 VSUBS 0.007307f
C854 B.n814 VSUBS 0.007307f
C855 B.n815 VSUBS 0.007307f
C856 B.n816 VSUBS 0.007307f
C857 B.n817 VSUBS 0.007307f
C858 B.n818 VSUBS 0.007307f
C859 B.n819 VSUBS 0.007307f
C860 B.n820 VSUBS 0.007307f
C861 B.n821 VSUBS 0.007307f
C862 B.n822 VSUBS 0.007307f
C863 B.n823 VSUBS 0.007307f
C864 B.n824 VSUBS 0.007307f
C865 B.n825 VSUBS 0.007307f
C866 B.n826 VSUBS 0.007307f
C867 B.n827 VSUBS 0.007307f
C868 B.n828 VSUBS 0.007307f
C869 B.n829 VSUBS 0.007307f
C870 B.n830 VSUBS 0.007307f
C871 B.n831 VSUBS 0.007307f
C872 B.n832 VSUBS 0.007307f
C873 B.n833 VSUBS 0.007307f
C874 B.n834 VSUBS 0.007307f
C875 B.n835 VSUBS 0.007307f
C876 B.n836 VSUBS 0.007307f
C877 B.n837 VSUBS 0.007307f
C878 B.n838 VSUBS 0.007307f
C879 B.n839 VSUBS 0.007307f
C880 B.n840 VSUBS 0.007307f
C881 B.n841 VSUBS 0.007307f
C882 B.n842 VSUBS 0.007307f
C883 B.n843 VSUBS 0.007307f
C884 B.n844 VSUBS 0.007307f
C885 B.n845 VSUBS 0.007307f
C886 B.n846 VSUBS 0.007307f
C887 B.n847 VSUBS 0.007307f
C888 B.n848 VSUBS 0.007307f
C889 B.n849 VSUBS 0.007307f
C890 B.n850 VSUBS 0.007307f
C891 B.n851 VSUBS 0.007307f
C892 B.n852 VSUBS 0.007307f
C893 B.n853 VSUBS 0.007307f
C894 B.n854 VSUBS 0.007307f
C895 B.n855 VSUBS 0.007307f
C896 B.n856 VSUBS 0.007307f
C897 B.n857 VSUBS 0.007307f
C898 B.n858 VSUBS 0.007307f
C899 B.n859 VSUBS 0.007307f
C900 B.n860 VSUBS 0.007307f
C901 B.n861 VSUBS 0.007307f
C902 B.n862 VSUBS 0.007307f
C903 B.n863 VSUBS 0.007307f
C904 B.n864 VSUBS 0.007307f
C905 B.n865 VSUBS 0.007307f
C906 B.n866 VSUBS 0.007307f
C907 B.n867 VSUBS 0.007307f
C908 B.n868 VSUBS 0.007307f
C909 B.n869 VSUBS 0.007307f
C910 B.n870 VSUBS 0.007307f
C911 B.n871 VSUBS 0.007307f
C912 B.n872 VSUBS 0.007307f
C913 B.n873 VSUBS 0.007307f
C914 B.n874 VSUBS 0.007307f
C915 B.n875 VSUBS 0.007307f
C916 B.n876 VSUBS 0.007307f
C917 B.n877 VSUBS 0.007307f
C918 B.n878 VSUBS 0.007307f
C919 B.n879 VSUBS 0.007307f
C920 B.n880 VSUBS 0.016268f
C921 B.n881 VSUBS 0.015538f
C922 B.n882 VSUBS 0.015538f
C923 B.n883 VSUBS 0.007307f
C924 B.n884 VSUBS 0.007307f
C925 B.n885 VSUBS 0.007307f
C926 B.n886 VSUBS 0.007307f
C927 B.n887 VSUBS 0.007307f
C928 B.n888 VSUBS 0.007307f
C929 B.n889 VSUBS 0.007307f
C930 B.n890 VSUBS 0.007307f
C931 B.n891 VSUBS 0.007307f
C932 B.n892 VSUBS 0.007307f
C933 B.n893 VSUBS 0.007307f
C934 B.n894 VSUBS 0.007307f
C935 B.n895 VSUBS 0.007307f
C936 B.n896 VSUBS 0.007307f
C937 B.n897 VSUBS 0.007307f
C938 B.n898 VSUBS 0.007307f
C939 B.n899 VSUBS 0.007307f
C940 B.n900 VSUBS 0.007307f
C941 B.n901 VSUBS 0.007307f
C942 B.n902 VSUBS 0.007307f
C943 B.n903 VSUBS 0.007307f
C944 B.n904 VSUBS 0.007307f
C945 B.n905 VSUBS 0.007307f
C946 B.n906 VSUBS 0.007307f
C947 B.n907 VSUBS 0.007307f
C948 B.n908 VSUBS 0.007307f
C949 B.n909 VSUBS 0.007307f
C950 B.n910 VSUBS 0.007307f
C951 B.n911 VSUBS 0.007307f
C952 B.n912 VSUBS 0.007307f
C953 B.n913 VSUBS 0.007307f
C954 B.n914 VSUBS 0.007307f
C955 B.n915 VSUBS 0.007307f
C956 B.n916 VSUBS 0.007307f
C957 B.n917 VSUBS 0.007307f
C958 B.n918 VSUBS 0.007307f
C959 B.n919 VSUBS 0.007307f
C960 B.n920 VSUBS 0.007307f
C961 B.n921 VSUBS 0.007307f
C962 B.n922 VSUBS 0.007307f
C963 B.n923 VSUBS 0.007307f
C964 B.n924 VSUBS 0.007307f
C965 B.n925 VSUBS 0.007307f
C966 B.n926 VSUBS 0.007307f
C967 B.n927 VSUBS 0.007307f
C968 B.n928 VSUBS 0.007307f
C969 B.n929 VSUBS 0.007307f
C970 B.n930 VSUBS 0.007307f
C971 B.n931 VSUBS 0.007307f
C972 B.n932 VSUBS 0.007307f
C973 B.n933 VSUBS 0.007307f
C974 B.n934 VSUBS 0.007307f
C975 B.n935 VSUBS 0.007307f
C976 B.n936 VSUBS 0.007307f
C977 B.n937 VSUBS 0.007307f
C978 B.n938 VSUBS 0.007307f
C979 B.n939 VSUBS 0.007307f
C980 B.n940 VSUBS 0.007307f
C981 B.n941 VSUBS 0.007307f
C982 B.n942 VSUBS 0.007307f
C983 B.n943 VSUBS 0.007307f
C984 B.n944 VSUBS 0.007307f
C985 B.n945 VSUBS 0.007307f
C986 B.n946 VSUBS 0.007307f
C987 B.n947 VSUBS 0.007307f
C988 B.n948 VSUBS 0.007307f
C989 B.n949 VSUBS 0.007307f
C990 B.n950 VSUBS 0.007307f
C991 B.n951 VSUBS 0.007307f
C992 B.n952 VSUBS 0.007307f
C993 B.n953 VSUBS 0.007307f
C994 B.n954 VSUBS 0.007307f
C995 B.n955 VSUBS 0.007307f
C996 B.n956 VSUBS 0.007307f
C997 B.n957 VSUBS 0.007307f
C998 B.n958 VSUBS 0.007307f
C999 B.n959 VSUBS 0.007307f
C1000 B.n960 VSUBS 0.007307f
C1001 B.n961 VSUBS 0.007307f
C1002 B.n962 VSUBS 0.007307f
C1003 B.n963 VSUBS 0.007307f
C1004 B.n964 VSUBS 0.007307f
C1005 B.n965 VSUBS 0.007307f
C1006 B.n966 VSUBS 0.007307f
C1007 B.n967 VSUBS 0.007307f
C1008 B.n968 VSUBS 0.007307f
C1009 B.n969 VSUBS 0.007307f
C1010 B.n970 VSUBS 0.007307f
C1011 B.n971 VSUBS 0.007307f
C1012 B.n972 VSUBS 0.007307f
C1013 B.n973 VSUBS 0.007307f
C1014 B.n974 VSUBS 0.007307f
C1015 B.n975 VSUBS 0.016545f
C1016 VDD2.t0 VSUBS 0.397504f
C1017 VDD2.t3 VSUBS 0.397504f
C1018 VDD2.n0 VSUBS 3.29074f
C1019 VDD2.t6 VSUBS 0.397504f
C1020 VDD2.t2 VSUBS 0.397504f
C1021 VDD2.n1 VSUBS 3.29074f
C1022 VDD2.n2 VSUBS 5.64447f
C1023 VDD2.t1 VSUBS 0.397504f
C1024 VDD2.t7 VSUBS 0.397504f
C1025 VDD2.n3 VSUBS 3.2689f
C1026 VDD2.n4 VSUBS 4.75415f
C1027 VDD2.t4 VSUBS 0.397504f
C1028 VDD2.t5 VSUBS 0.397504f
C1029 VDD2.n5 VSUBS 3.29067f
C1030 VN.t5 VSUBS 3.39677f
C1031 VN.n0 VSUBS 1.26554f
C1032 VN.n1 VSUBS 0.023438f
C1033 VN.n2 VSUBS 0.022141f
C1034 VN.n3 VSUBS 0.023438f
C1035 VN.t1 VSUBS 3.39677f
C1036 VN.n4 VSUBS 1.17805f
C1037 VN.n5 VSUBS 0.023438f
C1038 VN.n6 VSUBS 0.034215f
C1039 VN.n7 VSUBS 0.023438f
C1040 VN.n8 VSUBS 0.02535f
C1041 VN.t4 VSUBS 3.39677f
C1042 VN.n9 VSUBS 1.25007f
C1043 VN.t7 VSUBS 3.69034f
C1044 VN.n10 VSUBS 1.20149f
C1045 VN.n11 VSUBS 0.277408f
C1046 VN.n12 VSUBS 0.023438f
C1047 VN.n13 VSUBS 0.043682f
C1048 VN.n14 VSUBS 0.043682f
C1049 VN.n15 VSUBS 0.034215f
C1050 VN.n16 VSUBS 0.023438f
C1051 VN.n17 VSUBS 0.023438f
C1052 VN.n18 VSUBS 0.023438f
C1053 VN.n19 VSUBS 0.043682f
C1054 VN.n20 VSUBS 0.043682f
C1055 VN.n21 VSUBS 0.02535f
C1056 VN.n22 VSUBS 0.023438f
C1057 VN.n23 VSUBS 0.023438f
C1058 VN.n24 VSUBS 0.040446f
C1059 VN.n25 VSUBS 0.043682f
C1060 VN.n26 VSUBS 0.043016f
C1061 VN.n27 VSUBS 0.023438f
C1062 VN.n28 VSUBS 0.023438f
C1063 VN.n29 VSUBS 0.023438f
C1064 VN.n30 VSUBS 0.046954f
C1065 VN.n31 VSUBS 0.043682f
C1066 VN.n32 VSUBS 0.031819f
C1067 VN.n33 VSUBS 0.037828f
C1068 VN.n34 VSUBS 0.060142f
C1069 VN.t6 VSUBS 3.39677f
C1070 VN.n35 VSUBS 1.26554f
C1071 VN.n36 VSUBS 0.023438f
C1072 VN.n37 VSUBS 0.022141f
C1073 VN.n38 VSUBS 0.023438f
C1074 VN.t0 VSUBS 3.39677f
C1075 VN.n39 VSUBS 1.17805f
C1076 VN.n40 VSUBS 0.023438f
C1077 VN.n41 VSUBS 0.034215f
C1078 VN.n42 VSUBS 0.023438f
C1079 VN.n43 VSUBS 0.02535f
C1080 VN.t2 VSUBS 3.69034f
C1081 VN.t3 VSUBS 3.39677f
C1082 VN.n44 VSUBS 1.25007f
C1083 VN.n45 VSUBS 1.20149f
C1084 VN.n46 VSUBS 0.277408f
C1085 VN.n47 VSUBS 0.023438f
C1086 VN.n48 VSUBS 0.043682f
C1087 VN.n49 VSUBS 0.043682f
C1088 VN.n50 VSUBS 0.034215f
C1089 VN.n51 VSUBS 0.023438f
C1090 VN.n52 VSUBS 0.023438f
C1091 VN.n53 VSUBS 0.023438f
C1092 VN.n54 VSUBS 0.043682f
C1093 VN.n55 VSUBS 0.043682f
C1094 VN.n56 VSUBS 0.02535f
C1095 VN.n57 VSUBS 0.023438f
C1096 VN.n58 VSUBS 0.023438f
C1097 VN.n59 VSUBS 0.040446f
C1098 VN.n60 VSUBS 0.043682f
C1099 VN.n61 VSUBS 0.043016f
C1100 VN.n62 VSUBS 0.023438f
C1101 VN.n63 VSUBS 0.023438f
C1102 VN.n64 VSUBS 0.023438f
C1103 VN.n65 VSUBS 0.046954f
C1104 VN.n66 VSUBS 0.043682f
C1105 VN.n67 VSUBS 0.031819f
C1106 VN.n68 VSUBS 0.037828f
C1107 VN.n69 VSUBS 1.62402f
C1108 VDD1.t1 VSUBS 0.369093f
C1109 VDD1.t7 VSUBS 0.369093f
C1110 VDD1.n0 VSUBS 3.05724f
C1111 VDD1.t4 VSUBS 0.369093f
C1112 VDD1.t0 VSUBS 0.369093f
C1113 VDD1.n1 VSUBS 3.05553f
C1114 VDD1.t5 VSUBS 0.369093f
C1115 VDD1.t3 VSUBS 0.369093f
C1116 VDD1.n2 VSUBS 3.05553f
C1117 VDD1.n3 VSUBS 5.30157f
C1118 VDD1.t2 VSUBS 0.369093f
C1119 VDD1.t6 VSUBS 0.369093f
C1120 VDD1.n4 VSUBS 3.03525f
C1121 VDD1.n5 VSUBS 4.45126f
C1122 VTAIL.t3 VSUBS 0.307566f
C1123 VTAIL.t5 VSUBS 0.307566f
C1124 VTAIL.n0 VSUBS 2.39627f
C1125 VTAIL.n1 VSUBS 0.811887f
C1126 VTAIL.t0 VSUBS 3.13382f
C1127 VTAIL.n2 VSUBS 0.945594f
C1128 VTAIL.t15 VSUBS 3.13382f
C1129 VTAIL.n3 VSUBS 0.945594f
C1130 VTAIL.t9 VSUBS 0.307566f
C1131 VTAIL.t10 VSUBS 0.307566f
C1132 VTAIL.n4 VSUBS 2.39627f
C1133 VTAIL.n5 VSUBS 1.05533f
C1134 VTAIL.t12 VSUBS 3.13382f
C1135 VTAIL.n6 VSUBS 2.57004f
C1136 VTAIL.t1 VSUBS 3.13385f
C1137 VTAIL.n7 VSUBS 2.57001f
C1138 VTAIL.t4 VSUBS 0.307566f
C1139 VTAIL.t7 VSUBS 0.307566f
C1140 VTAIL.n8 VSUBS 2.39627f
C1141 VTAIL.n9 VSUBS 1.05533f
C1142 VTAIL.t6 VSUBS 3.13385f
C1143 VTAIL.n10 VSUBS 0.945571f
C1144 VTAIL.t8 VSUBS 3.13385f
C1145 VTAIL.n11 VSUBS 0.945571f
C1146 VTAIL.t14 VSUBS 0.307566f
C1147 VTAIL.t13 VSUBS 0.307566f
C1148 VTAIL.n12 VSUBS 2.39627f
C1149 VTAIL.n13 VSUBS 1.05533f
C1150 VTAIL.t11 VSUBS 3.13382f
C1151 VTAIL.n14 VSUBS 2.57004f
C1152 VTAIL.t2 VSUBS 3.13382f
C1153 VTAIL.n15 VSUBS 2.56545f
C1154 VP.t4 VSUBS 3.67477f
C1155 VP.n0 VSUBS 1.36912f
C1156 VP.n1 VSUBS 0.025356f
C1157 VP.n2 VSUBS 0.023953f
C1158 VP.n3 VSUBS 0.025356f
C1159 VP.t2 VSUBS 3.67477f
C1160 VP.n4 VSUBS 1.27447f
C1161 VP.n5 VSUBS 0.025356f
C1162 VP.n6 VSUBS 0.037015f
C1163 VP.n7 VSUBS 0.025356f
C1164 VP.n8 VSUBS 0.027424f
C1165 VP.n9 VSUBS 0.025356f
C1166 VP.n10 VSUBS 0.023953f
C1167 VP.n11 VSUBS 0.025356f
C1168 VP.t3 VSUBS 3.67477f
C1169 VP.n12 VSUBS 1.36912f
C1170 VP.t1 VSUBS 3.67477f
C1171 VP.n13 VSUBS 1.36912f
C1172 VP.n14 VSUBS 0.025356f
C1173 VP.n15 VSUBS 0.023953f
C1174 VP.n16 VSUBS 0.025356f
C1175 VP.t5 VSUBS 3.67477f
C1176 VP.n17 VSUBS 1.27447f
C1177 VP.n18 VSUBS 0.025356f
C1178 VP.n19 VSUBS 0.037015f
C1179 VP.n20 VSUBS 0.025356f
C1180 VP.n21 VSUBS 0.027424f
C1181 VP.t6 VSUBS 3.99237f
C1182 VP.t0 VSUBS 3.67477f
C1183 VP.n22 VSUBS 1.35238f
C1184 VP.n23 VSUBS 1.29982f
C1185 VP.n24 VSUBS 0.300112f
C1186 VP.n25 VSUBS 0.025356f
C1187 VP.n26 VSUBS 0.047257f
C1188 VP.n27 VSUBS 0.047257f
C1189 VP.n28 VSUBS 0.037015f
C1190 VP.n29 VSUBS 0.025356f
C1191 VP.n30 VSUBS 0.025356f
C1192 VP.n31 VSUBS 0.025356f
C1193 VP.n32 VSUBS 0.047257f
C1194 VP.n33 VSUBS 0.047257f
C1195 VP.n34 VSUBS 0.027424f
C1196 VP.n35 VSUBS 0.025356f
C1197 VP.n36 VSUBS 0.025356f
C1198 VP.n37 VSUBS 0.043756f
C1199 VP.n38 VSUBS 0.047257f
C1200 VP.n39 VSUBS 0.046537f
C1201 VP.n40 VSUBS 0.025356f
C1202 VP.n41 VSUBS 0.025356f
C1203 VP.n42 VSUBS 0.025356f
C1204 VP.n43 VSUBS 0.050796f
C1205 VP.n44 VSUBS 0.047257f
C1206 VP.n45 VSUBS 0.034424f
C1207 VP.n46 VSUBS 0.040924f
C1208 VP.n47 VSUBS 1.74701f
C1209 VP.n48 VSUBS 1.76292f
C1210 VP.n49 VSUBS 0.040924f
C1211 VP.n50 VSUBS 0.034424f
C1212 VP.n51 VSUBS 0.047257f
C1213 VP.n52 VSUBS 0.050796f
C1214 VP.n53 VSUBS 0.025356f
C1215 VP.n54 VSUBS 0.025356f
C1216 VP.n55 VSUBS 0.025356f
C1217 VP.n56 VSUBS 0.046537f
C1218 VP.n57 VSUBS 0.047257f
C1219 VP.t7 VSUBS 3.67477f
C1220 VP.n58 VSUBS 1.27447f
C1221 VP.n59 VSUBS 0.043756f
C1222 VP.n60 VSUBS 0.025356f
C1223 VP.n61 VSUBS 0.025356f
C1224 VP.n62 VSUBS 0.025356f
C1225 VP.n63 VSUBS 0.047257f
C1226 VP.n64 VSUBS 0.047257f
C1227 VP.n65 VSUBS 0.037015f
C1228 VP.n66 VSUBS 0.025356f
C1229 VP.n67 VSUBS 0.025356f
C1230 VP.n68 VSUBS 0.025356f
C1231 VP.n69 VSUBS 0.047257f
C1232 VP.n70 VSUBS 0.047257f
C1233 VP.n71 VSUBS 0.027424f
C1234 VP.n72 VSUBS 0.025356f
C1235 VP.n73 VSUBS 0.025356f
C1236 VP.n74 VSUBS 0.043756f
C1237 VP.n75 VSUBS 0.047257f
C1238 VP.n76 VSUBS 0.046537f
C1239 VP.n77 VSUBS 0.025356f
C1240 VP.n78 VSUBS 0.025356f
C1241 VP.n79 VSUBS 0.025356f
C1242 VP.n80 VSUBS 0.050796f
C1243 VP.n81 VSUBS 0.047257f
C1244 VP.n82 VSUBS 0.034424f
C1245 VP.n83 VSUBS 0.040924f
C1246 VP.n84 VSUBS 0.065064f
.ends

