* NGSPICE file created from diff_pair_sample_1798.ext - technology: sky130A

.subckt diff_pair_sample_1798 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=3.9624 ps=21.1 w=10.16 l=1.31
X1 VTAIL.t12 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=1.6764 ps=10.49 w=10.16 l=1.31
X2 VDD1.t7 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X3 VTAIL.t1 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X4 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=0 ps=0 w=10.16 l=1.31
X5 VTAIL.t11 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=0 ps=0 w=10.16 l=1.31
X7 VTAIL.t8 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X8 VDD2.t3 VN.t4 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X9 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=3.9624 ps=21.1 w=10.16 l=1.31
X10 VDD2.t2 VN.t5 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=3.9624 ps=21.1 w=10.16 l=1.31
X11 VDD2.t1 VN.t6 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X12 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=0 ps=0 w=10.16 l=1.31
X13 VTAIL.t5 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=1.6764 ps=10.49 w=10.16 l=1.31
X14 VDD1.t3 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=3.9624 ps=21.1 w=10.16 l=1.31
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=0 ps=0 w=10.16 l=1.31
X16 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X17 VTAIL.t15 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=1.6764 ps=10.49 w=10.16 l=1.31
X18 VDD1.t1 VP.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6764 pd=10.49 as=1.6764 ps=10.49 w=10.16 l=1.31
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.9624 pd=21.1 as=1.6764 ps=10.49 w=10.16 l=1.31
R0 VN.n5 VN.t1 214.504
R1 VN.n25 VN.t5 214.504
R2 VN.n4 VN.t4 186.913
R3 VN.n10 VN.t2 186.913
R4 VN.n17 VN.t0 186.913
R5 VN.n24 VN.t3 186.913
R6 VN.n22 VN.t6 186.913
R7 VN.n36 VN.t7 186.913
R8 VN.n18 VN.n17 175.564
R9 VN.n37 VN.n36 175.564
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n29 VN.n21 161.3
R15 VN.n28 VN.n27 161.3
R16 VN.n26 VN.n23 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n5 VN.n4 62.2212
R25 VN.n25 VN.n24 62.2212
R26 VN.n9 VN.n8 56.5617
R27 VN.n29 VN.n28 56.5617
R28 VN.n15 VN.n1 51.2335
R29 VN.n34 VN.n20 51.2335
R30 VN VN.n37 43.7297
R31 VN.n16 VN.n15 29.9206
R32 VN.n35 VN.n34 29.9206
R33 VN.n26 VN.n25 27.6221
R34 VN.n6 VN.n5 27.6221
R35 VN.n8 VN.n3 24.5923
R36 VN.n11 VN.n9 24.5923
R37 VN.n28 VN.n23 24.5923
R38 VN.n30 VN.n29 24.5923
R39 VN.n10 VN.n1 21.1495
R40 VN.n22 VN.n20 21.1495
R41 VN.n17 VN.n16 10.3291
R42 VN.n36 VN.n35 10.3291
R43 VN.n4 VN.n3 3.44336
R44 VN.n11 VN.n10 3.44336
R45 VN.n24 VN.n23 3.44336
R46 VN.n30 VN.n22 3.44336
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n27 VN.n21 0.189894
R53 VN.n27 VN.n26 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VTAIL.n434 VTAIL.n386 289.615
R63 VTAIL.n50 VTAIL.n2 289.615
R64 VTAIL.n104 VTAIL.n56 289.615
R65 VTAIL.n160 VTAIL.n112 289.615
R66 VTAIL.n380 VTAIL.n332 289.615
R67 VTAIL.n324 VTAIL.n276 289.615
R68 VTAIL.n270 VTAIL.n222 289.615
R69 VTAIL.n214 VTAIL.n166 289.615
R70 VTAIL.n402 VTAIL.n401 185
R71 VTAIL.n407 VTAIL.n406 185
R72 VTAIL.n409 VTAIL.n408 185
R73 VTAIL.n398 VTAIL.n397 185
R74 VTAIL.n415 VTAIL.n414 185
R75 VTAIL.n417 VTAIL.n416 185
R76 VTAIL.n394 VTAIL.n393 185
R77 VTAIL.n424 VTAIL.n423 185
R78 VTAIL.n425 VTAIL.n392 185
R79 VTAIL.n427 VTAIL.n426 185
R80 VTAIL.n390 VTAIL.n389 185
R81 VTAIL.n433 VTAIL.n432 185
R82 VTAIL.n435 VTAIL.n434 185
R83 VTAIL.n18 VTAIL.n17 185
R84 VTAIL.n23 VTAIL.n22 185
R85 VTAIL.n25 VTAIL.n24 185
R86 VTAIL.n14 VTAIL.n13 185
R87 VTAIL.n31 VTAIL.n30 185
R88 VTAIL.n33 VTAIL.n32 185
R89 VTAIL.n10 VTAIL.n9 185
R90 VTAIL.n40 VTAIL.n39 185
R91 VTAIL.n41 VTAIL.n8 185
R92 VTAIL.n43 VTAIL.n42 185
R93 VTAIL.n6 VTAIL.n5 185
R94 VTAIL.n49 VTAIL.n48 185
R95 VTAIL.n51 VTAIL.n50 185
R96 VTAIL.n72 VTAIL.n71 185
R97 VTAIL.n77 VTAIL.n76 185
R98 VTAIL.n79 VTAIL.n78 185
R99 VTAIL.n68 VTAIL.n67 185
R100 VTAIL.n85 VTAIL.n84 185
R101 VTAIL.n87 VTAIL.n86 185
R102 VTAIL.n64 VTAIL.n63 185
R103 VTAIL.n94 VTAIL.n93 185
R104 VTAIL.n95 VTAIL.n62 185
R105 VTAIL.n97 VTAIL.n96 185
R106 VTAIL.n60 VTAIL.n59 185
R107 VTAIL.n103 VTAIL.n102 185
R108 VTAIL.n105 VTAIL.n104 185
R109 VTAIL.n128 VTAIL.n127 185
R110 VTAIL.n133 VTAIL.n132 185
R111 VTAIL.n135 VTAIL.n134 185
R112 VTAIL.n124 VTAIL.n123 185
R113 VTAIL.n141 VTAIL.n140 185
R114 VTAIL.n143 VTAIL.n142 185
R115 VTAIL.n120 VTAIL.n119 185
R116 VTAIL.n150 VTAIL.n149 185
R117 VTAIL.n151 VTAIL.n118 185
R118 VTAIL.n153 VTAIL.n152 185
R119 VTAIL.n116 VTAIL.n115 185
R120 VTAIL.n159 VTAIL.n158 185
R121 VTAIL.n161 VTAIL.n160 185
R122 VTAIL.n381 VTAIL.n380 185
R123 VTAIL.n379 VTAIL.n378 185
R124 VTAIL.n336 VTAIL.n335 185
R125 VTAIL.n373 VTAIL.n372 185
R126 VTAIL.n371 VTAIL.n338 185
R127 VTAIL.n370 VTAIL.n369 185
R128 VTAIL.n341 VTAIL.n339 185
R129 VTAIL.n364 VTAIL.n363 185
R130 VTAIL.n362 VTAIL.n361 185
R131 VTAIL.n345 VTAIL.n344 185
R132 VTAIL.n356 VTAIL.n355 185
R133 VTAIL.n354 VTAIL.n353 185
R134 VTAIL.n349 VTAIL.n348 185
R135 VTAIL.n325 VTAIL.n324 185
R136 VTAIL.n323 VTAIL.n322 185
R137 VTAIL.n280 VTAIL.n279 185
R138 VTAIL.n317 VTAIL.n316 185
R139 VTAIL.n315 VTAIL.n282 185
R140 VTAIL.n314 VTAIL.n313 185
R141 VTAIL.n285 VTAIL.n283 185
R142 VTAIL.n308 VTAIL.n307 185
R143 VTAIL.n306 VTAIL.n305 185
R144 VTAIL.n289 VTAIL.n288 185
R145 VTAIL.n300 VTAIL.n299 185
R146 VTAIL.n298 VTAIL.n297 185
R147 VTAIL.n293 VTAIL.n292 185
R148 VTAIL.n271 VTAIL.n270 185
R149 VTAIL.n269 VTAIL.n268 185
R150 VTAIL.n226 VTAIL.n225 185
R151 VTAIL.n263 VTAIL.n262 185
R152 VTAIL.n261 VTAIL.n228 185
R153 VTAIL.n260 VTAIL.n259 185
R154 VTAIL.n231 VTAIL.n229 185
R155 VTAIL.n254 VTAIL.n253 185
R156 VTAIL.n252 VTAIL.n251 185
R157 VTAIL.n235 VTAIL.n234 185
R158 VTAIL.n246 VTAIL.n245 185
R159 VTAIL.n244 VTAIL.n243 185
R160 VTAIL.n239 VTAIL.n238 185
R161 VTAIL.n215 VTAIL.n214 185
R162 VTAIL.n213 VTAIL.n212 185
R163 VTAIL.n170 VTAIL.n169 185
R164 VTAIL.n207 VTAIL.n206 185
R165 VTAIL.n205 VTAIL.n172 185
R166 VTAIL.n204 VTAIL.n203 185
R167 VTAIL.n175 VTAIL.n173 185
R168 VTAIL.n198 VTAIL.n197 185
R169 VTAIL.n196 VTAIL.n195 185
R170 VTAIL.n179 VTAIL.n178 185
R171 VTAIL.n190 VTAIL.n189 185
R172 VTAIL.n188 VTAIL.n187 185
R173 VTAIL.n183 VTAIL.n182 185
R174 VTAIL.n403 VTAIL.t9 149.524
R175 VTAIL.n19 VTAIL.t12 149.524
R176 VTAIL.n73 VTAIL.t6 149.524
R177 VTAIL.n129 VTAIL.t5 149.524
R178 VTAIL.n350 VTAIL.t3 149.524
R179 VTAIL.n294 VTAIL.t0 149.524
R180 VTAIL.n240 VTAIL.t13 149.524
R181 VTAIL.n184 VTAIL.t15 149.524
R182 VTAIL.n407 VTAIL.n401 104.615
R183 VTAIL.n408 VTAIL.n407 104.615
R184 VTAIL.n408 VTAIL.n397 104.615
R185 VTAIL.n415 VTAIL.n397 104.615
R186 VTAIL.n416 VTAIL.n415 104.615
R187 VTAIL.n416 VTAIL.n393 104.615
R188 VTAIL.n424 VTAIL.n393 104.615
R189 VTAIL.n425 VTAIL.n424 104.615
R190 VTAIL.n426 VTAIL.n425 104.615
R191 VTAIL.n426 VTAIL.n389 104.615
R192 VTAIL.n433 VTAIL.n389 104.615
R193 VTAIL.n434 VTAIL.n433 104.615
R194 VTAIL.n23 VTAIL.n17 104.615
R195 VTAIL.n24 VTAIL.n23 104.615
R196 VTAIL.n24 VTAIL.n13 104.615
R197 VTAIL.n31 VTAIL.n13 104.615
R198 VTAIL.n32 VTAIL.n31 104.615
R199 VTAIL.n32 VTAIL.n9 104.615
R200 VTAIL.n40 VTAIL.n9 104.615
R201 VTAIL.n41 VTAIL.n40 104.615
R202 VTAIL.n42 VTAIL.n41 104.615
R203 VTAIL.n42 VTAIL.n5 104.615
R204 VTAIL.n49 VTAIL.n5 104.615
R205 VTAIL.n50 VTAIL.n49 104.615
R206 VTAIL.n77 VTAIL.n71 104.615
R207 VTAIL.n78 VTAIL.n77 104.615
R208 VTAIL.n78 VTAIL.n67 104.615
R209 VTAIL.n85 VTAIL.n67 104.615
R210 VTAIL.n86 VTAIL.n85 104.615
R211 VTAIL.n86 VTAIL.n63 104.615
R212 VTAIL.n94 VTAIL.n63 104.615
R213 VTAIL.n95 VTAIL.n94 104.615
R214 VTAIL.n96 VTAIL.n95 104.615
R215 VTAIL.n96 VTAIL.n59 104.615
R216 VTAIL.n103 VTAIL.n59 104.615
R217 VTAIL.n104 VTAIL.n103 104.615
R218 VTAIL.n133 VTAIL.n127 104.615
R219 VTAIL.n134 VTAIL.n133 104.615
R220 VTAIL.n134 VTAIL.n123 104.615
R221 VTAIL.n141 VTAIL.n123 104.615
R222 VTAIL.n142 VTAIL.n141 104.615
R223 VTAIL.n142 VTAIL.n119 104.615
R224 VTAIL.n150 VTAIL.n119 104.615
R225 VTAIL.n151 VTAIL.n150 104.615
R226 VTAIL.n152 VTAIL.n151 104.615
R227 VTAIL.n152 VTAIL.n115 104.615
R228 VTAIL.n159 VTAIL.n115 104.615
R229 VTAIL.n160 VTAIL.n159 104.615
R230 VTAIL.n380 VTAIL.n379 104.615
R231 VTAIL.n379 VTAIL.n335 104.615
R232 VTAIL.n372 VTAIL.n335 104.615
R233 VTAIL.n372 VTAIL.n371 104.615
R234 VTAIL.n371 VTAIL.n370 104.615
R235 VTAIL.n370 VTAIL.n339 104.615
R236 VTAIL.n363 VTAIL.n339 104.615
R237 VTAIL.n363 VTAIL.n362 104.615
R238 VTAIL.n362 VTAIL.n344 104.615
R239 VTAIL.n355 VTAIL.n344 104.615
R240 VTAIL.n355 VTAIL.n354 104.615
R241 VTAIL.n354 VTAIL.n348 104.615
R242 VTAIL.n324 VTAIL.n323 104.615
R243 VTAIL.n323 VTAIL.n279 104.615
R244 VTAIL.n316 VTAIL.n279 104.615
R245 VTAIL.n316 VTAIL.n315 104.615
R246 VTAIL.n315 VTAIL.n314 104.615
R247 VTAIL.n314 VTAIL.n283 104.615
R248 VTAIL.n307 VTAIL.n283 104.615
R249 VTAIL.n307 VTAIL.n306 104.615
R250 VTAIL.n306 VTAIL.n288 104.615
R251 VTAIL.n299 VTAIL.n288 104.615
R252 VTAIL.n299 VTAIL.n298 104.615
R253 VTAIL.n298 VTAIL.n292 104.615
R254 VTAIL.n270 VTAIL.n269 104.615
R255 VTAIL.n269 VTAIL.n225 104.615
R256 VTAIL.n262 VTAIL.n225 104.615
R257 VTAIL.n262 VTAIL.n261 104.615
R258 VTAIL.n261 VTAIL.n260 104.615
R259 VTAIL.n260 VTAIL.n229 104.615
R260 VTAIL.n253 VTAIL.n229 104.615
R261 VTAIL.n253 VTAIL.n252 104.615
R262 VTAIL.n252 VTAIL.n234 104.615
R263 VTAIL.n245 VTAIL.n234 104.615
R264 VTAIL.n245 VTAIL.n244 104.615
R265 VTAIL.n244 VTAIL.n238 104.615
R266 VTAIL.n214 VTAIL.n213 104.615
R267 VTAIL.n213 VTAIL.n169 104.615
R268 VTAIL.n206 VTAIL.n169 104.615
R269 VTAIL.n206 VTAIL.n205 104.615
R270 VTAIL.n205 VTAIL.n204 104.615
R271 VTAIL.n204 VTAIL.n173 104.615
R272 VTAIL.n197 VTAIL.n173 104.615
R273 VTAIL.n197 VTAIL.n196 104.615
R274 VTAIL.n196 VTAIL.n178 104.615
R275 VTAIL.n189 VTAIL.n178 104.615
R276 VTAIL.n189 VTAIL.n188 104.615
R277 VTAIL.n188 VTAIL.n182 104.615
R278 VTAIL.t9 VTAIL.n401 52.3082
R279 VTAIL.t12 VTAIL.n17 52.3082
R280 VTAIL.t6 VTAIL.n71 52.3082
R281 VTAIL.t5 VTAIL.n127 52.3082
R282 VTAIL.t3 VTAIL.n348 52.3082
R283 VTAIL.t0 VTAIL.n292 52.3082
R284 VTAIL.t13 VTAIL.n238 52.3082
R285 VTAIL.t15 VTAIL.n182 52.3082
R286 VTAIL.n331 VTAIL.n330 49.8403
R287 VTAIL.n221 VTAIL.n220 49.8403
R288 VTAIL.n1 VTAIL.n0 49.8402
R289 VTAIL.n111 VTAIL.n110 49.8402
R290 VTAIL.n439 VTAIL.n438 36.0641
R291 VTAIL.n55 VTAIL.n54 36.0641
R292 VTAIL.n109 VTAIL.n108 36.0641
R293 VTAIL.n165 VTAIL.n164 36.0641
R294 VTAIL.n385 VTAIL.n384 36.0641
R295 VTAIL.n329 VTAIL.n328 36.0641
R296 VTAIL.n275 VTAIL.n274 36.0641
R297 VTAIL.n219 VTAIL.n218 36.0641
R298 VTAIL.n439 VTAIL.n385 22.5393
R299 VTAIL.n219 VTAIL.n165 22.5393
R300 VTAIL.n427 VTAIL.n392 13.1884
R301 VTAIL.n43 VTAIL.n8 13.1884
R302 VTAIL.n97 VTAIL.n62 13.1884
R303 VTAIL.n153 VTAIL.n118 13.1884
R304 VTAIL.n373 VTAIL.n338 13.1884
R305 VTAIL.n317 VTAIL.n282 13.1884
R306 VTAIL.n263 VTAIL.n228 13.1884
R307 VTAIL.n207 VTAIL.n172 13.1884
R308 VTAIL.n423 VTAIL.n422 12.8005
R309 VTAIL.n428 VTAIL.n390 12.8005
R310 VTAIL.n39 VTAIL.n38 12.8005
R311 VTAIL.n44 VTAIL.n6 12.8005
R312 VTAIL.n93 VTAIL.n92 12.8005
R313 VTAIL.n98 VTAIL.n60 12.8005
R314 VTAIL.n149 VTAIL.n148 12.8005
R315 VTAIL.n154 VTAIL.n116 12.8005
R316 VTAIL.n374 VTAIL.n336 12.8005
R317 VTAIL.n369 VTAIL.n340 12.8005
R318 VTAIL.n318 VTAIL.n280 12.8005
R319 VTAIL.n313 VTAIL.n284 12.8005
R320 VTAIL.n264 VTAIL.n226 12.8005
R321 VTAIL.n259 VTAIL.n230 12.8005
R322 VTAIL.n208 VTAIL.n170 12.8005
R323 VTAIL.n203 VTAIL.n174 12.8005
R324 VTAIL.n421 VTAIL.n394 12.0247
R325 VTAIL.n432 VTAIL.n431 12.0247
R326 VTAIL.n37 VTAIL.n10 12.0247
R327 VTAIL.n48 VTAIL.n47 12.0247
R328 VTAIL.n91 VTAIL.n64 12.0247
R329 VTAIL.n102 VTAIL.n101 12.0247
R330 VTAIL.n147 VTAIL.n120 12.0247
R331 VTAIL.n158 VTAIL.n157 12.0247
R332 VTAIL.n378 VTAIL.n377 12.0247
R333 VTAIL.n368 VTAIL.n341 12.0247
R334 VTAIL.n322 VTAIL.n321 12.0247
R335 VTAIL.n312 VTAIL.n285 12.0247
R336 VTAIL.n268 VTAIL.n267 12.0247
R337 VTAIL.n258 VTAIL.n231 12.0247
R338 VTAIL.n212 VTAIL.n211 12.0247
R339 VTAIL.n202 VTAIL.n175 12.0247
R340 VTAIL.n418 VTAIL.n417 11.249
R341 VTAIL.n435 VTAIL.n388 11.249
R342 VTAIL.n34 VTAIL.n33 11.249
R343 VTAIL.n51 VTAIL.n4 11.249
R344 VTAIL.n88 VTAIL.n87 11.249
R345 VTAIL.n105 VTAIL.n58 11.249
R346 VTAIL.n144 VTAIL.n143 11.249
R347 VTAIL.n161 VTAIL.n114 11.249
R348 VTAIL.n381 VTAIL.n334 11.249
R349 VTAIL.n365 VTAIL.n364 11.249
R350 VTAIL.n325 VTAIL.n278 11.249
R351 VTAIL.n309 VTAIL.n308 11.249
R352 VTAIL.n271 VTAIL.n224 11.249
R353 VTAIL.n255 VTAIL.n254 11.249
R354 VTAIL.n215 VTAIL.n168 11.249
R355 VTAIL.n199 VTAIL.n198 11.249
R356 VTAIL.n414 VTAIL.n396 10.4732
R357 VTAIL.n436 VTAIL.n386 10.4732
R358 VTAIL.n30 VTAIL.n12 10.4732
R359 VTAIL.n52 VTAIL.n2 10.4732
R360 VTAIL.n84 VTAIL.n66 10.4732
R361 VTAIL.n106 VTAIL.n56 10.4732
R362 VTAIL.n140 VTAIL.n122 10.4732
R363 VTAIL.n162 VTAIL.n112 10.4732
R364 VTAIL.n382 VTAIL.n332 10.4732
R365 VTAIL.n361 VTAIL.n343 10.4732
R366 VTAIL.n326 VTAIL.n276 10.4732
R367 VTAIL.n305 VTAIL.n287 10.4732
R368 VTAIL.n272 VTAIL.n222 10.4732
R369 VTAIL.n251 VTAIL.n233 10.4732
R370 VTAIL.n216 VTAIL.n166 10.4732
R371 VTAIL.n195 VTAIL.n177 10.4732
R372 VTAIL.n403 VTAIL.n402 10.2747
R373 VTAIL.n19 VTAIL.n18 10.2747
R374 VTAIL.n73 VTAIL.n72 10.2747
R375 VTAIL.n129 VTAIL.n128 10.2747
R376 VTAIL.n350 VTAIL.n349 10.2747
R377 VTAIL.n294 VTAIL.n293 10.2747
R378 VTAIL.n240 VTAIL.n239 10.2747
R379 VTAIL.n184 VTAIL.n183 10.2747
R380 VTAIL.n413 VTAIL.n398 9.69747
R381 VTAIL.n29 VTAIL.n14 9.69747
R382 VTAIL.n83 VTAIL.n68 9.69747
R383 VTAIL.n139 VTAIL.n124 9.69747
R384 VTAIL.n360 VTAIL.n345 9.69747
R385 VTAIL.n304 VTAIL.n289 9.69747
R386 VTAIL.n250 VTAIL.n235 9.69747
R387 VTAIL.n194 VTAIL.n179 9.69747
R388 VTAIL.n438 VTAIL.n437 9.45567
R389 VTAIL.n54 VTAIL.n53 9.45567
R390 VTAIL.n108 VTAIL.n107 9.45567
R391 VTAIL.n164 VTAIL.n163 9.45567
R392 VTAIL.n384 VTAIL.n383 9.45567
R393 VTAIL.n328 VTAIL.n327 9.45567
R394 VTAIL.n274 VTAIL.n273 9.45567
R395 VTAIL.n218 VTAIL.n217 9.45567
R396 VTAIL.n437 VTAIL.n436 9.3005
R397 VTAIL.n388 VTAIL.n387 9.3005
R398 VTAIL.n431 VTAIL.n430 9.3005
R399 VTAIL.n429 VTAIL.n428 9.3005
R400 VTAIL.n405 VTAIL.n404 9.3005
R401 VTAIL.n400 VTAIL.n399 9.3005
R402 VTAIL.n411 VTAIL.n410 9.3005
R403 VTAIL.n413 VTAIL.n412 9.3005
R404 VTAIL.n396 VTAIL.n395 9.3005
R405 VTAIL.n419 VTAIL.n418 9.3005
R406 VTAIL.n421 VTAIL.n420 9.3005
R407 VTAIL.n422 VTAIL.n391 9.3005
R408 VTAIL.n53 VTAIL.n52 9.3005
R409 VTAIL.n4 VTAIL.n3 9.3005
R410 VTAIL.n47 VTAIL.n46 9.3005
R411 VTAIL.n45 VTAIL.n44 9.3005
R412 VTAIL.n21 VTAIL.n20 9.3005
R413 VTAIL.n16 VTAIL.n15 9.3005
R414 VTAIL.n27 VTAIL.n26 9.3005
R415 VTAIL.n29 VTAIL.n28 9.3005
R416 VTAIL.n12 VTAIL.n11 9.3005
R417 VTAIL.n35 VTAIL.n34 9.3005
R418 VTAIL.n37 VTAIL.n36 9.3005
R419 VTAIL.n38 VTAIL.n7 9.3005
R420 VTAIL.n107 VTAIL.n106 9.3005
R421 VTAIL.n58 VTAIL.n57 9.3005
R422 VTAIL.n101 VTAIL.n100 9.3005
R423 VTAIL.n99 VTAIL.n98 9.3005
R424 VTAIL.n75 VTAIL.n74 9.3005
R425 VTAIL.n70 VTAIL.n69 9.3005
R426 VTAIL.n81 VTAIL.n80 9.3005
R427 VTAIL.n83 VTAIL.n82 9.3005
R428 VTAIL.n66 VTAIL.n65 9.3005
R429 VTAIL.n89 VTAIL.n88 9.3005
R430 VTAIL.n91 VTAIL.n90 9.3005
R431 VTAIL.n92 VTAIL.n61 9.3005
R432 VTAIL.n163 VTAIL.n162 9.3005
R433 VTAIL.n114 VTAIL.n113 9.3005
R434 VTAIL.n157 VTAIL.n156 9.3005
R435 VTAIL.n155 VTAIL.n154 9.3005
R436 VTAIL.n131 VTAIL.n130 9.3005
R437 VTAIL.n126 VTAIL.n125 9.3005
R438 VTAIL.n137 VTAIL.n136 9.3005
R439 VTAIL.n139 VTAIL.n138 9.3005
R440 VTAIL.n122 VTAIL.n121 9.3005
R441 VTAIL.n145 VTAIL.n144 9.3005
R442 VTAIL.n147 VTAIL.n146 9.3005
R443 VTAIL.n148 VTAIL.n117 9.3005
R444 VTAIL.n352 VTAIL.n351 9.3005
R445 VTAIL.n347 VTAIL.n346 9.3005
R446 VTAIL.n358 VTAIL.n357 9.3005
R447 VTAIL.n360 VTAIL.n359 9.3005
R448 VTAIL.n343 VTAIL.n342 9.3005
R449 VTAIL.n366 VTAIL.n365 9.3005
R450 VTAIL.n368 VTAIL.n367 9.3005
R451 VTAIL.n340 VTAIL.n337 9.3005
R452 VTAIL.n383 VTAIL.n382 9.3005
R453 VTAIL.n334 VTAIL.n333 9.3005
R454 VTAIL.n377 VTAIL.n376 9.3005
R455 VTAIL.n375 VTAIL.n374 9.3005
R456 VTAIL.n296 VTAIL.n295 9.3005
R457 VTAIL.n291 VTAIL.n290 9.3005
R458 VTAIL.n302 VTAIL.n301 9.3005
R459 VTAIL.n304 VTAIL.n303 9.3005
R460 VTAIL.n287 VTAIL.n286 9.3005
R461 VTAIL.n310 VTAIL.n309 9.3005
R462 VTAIL.n312 VTAIL.n311 9.3005
R463 VTAIL.n284 VTAIL.n281 9.3005
R464 VTAIL.n327 VTAIL.n326 9.3005
R465 VTAIL.n278 VTAIL.n277 9.3005
R466 VTAIL.n321 VTAIL.n320 9.3005
R467 VTAIL.n319 VTAIL.n318 9.3005
R468 VTAIL.n242 VTAIL.n241 9.3005
R469 VTAIL.n237 VTAIL.n236 9.3005
R470 VTAIL.n248 VTAIL.n247 9.3005
R471 VTAIL.n250 VTAIL.n249 9.3005
R472 VTAIL.n233 VTAIL.n232 9.3005
R473 VTAIL.n256 VTAIL.n255 9.3005
R474 VTAIL.n258 VTAIL.n257 9.3005
R475 VTAIL.n230 VTAIL.n227 9.3005
R476 VTAIL.n273 VTAIL.n272 9.3005
R477 VTAIL.n224 VTAIL.n223 9.3005
R478 VTAIL.n267 VTAIL.n266 9.3005
R479 VTAIL.n265 VTAIL.n264 9.3005
R480 VTAIL.n186 VTAIL.n185 9.3005
R481 VTAIL.n181 VTAIL.n180 9.3005
R482 VTAIL.n192 VTAIL.n191 9.3005
R483 VTAIL.n194 VTAIL.n193 9.3005
R484 VTAIL.n177 VTAIL.n176 9.3005
R485 VTAIL.n200 VTAIL.n199 9.3005
R486 VTAIL.n202 VTAIL.n201 9.3005
R487 VTAIL.n174 VTAIL.n171 9.3005
R488 VTAIL.n217 VTAIL.n216 9.3005
R489 VTAIL.n168 VTAIL.n167 9.3005
R490 VTAIL.n211 VTAIL.n210 9.3005
R491 VTAIL.n209 VTAIL.n208 9.3005
R492 VTAIL.n410 VTAIL.n409 8.92171
R493 VTAIL.n26 VTAIL.n25 8.92171
R494 VTAIL.n80 VTAIL.n79 8.92171
R495 VTAIL.n136 VTAIL.n135 8.92171
R496 VTAIL.n357 VTAIL.n356 8.92171
R497 VTAIL.n301 VTAIL.n300 8.92171
R498 VTAIL.n247 VTAIL.n246 8.92171
R499 VTAIL.n191 VTAIL.n190 8.92171
R500 VTAIL.n406 VTAIL.n400 8.14595
R501 VTAIL.n22 VTAIL.n16 8.14595
R502 VTAIL.n76 VTAIL.n70 8.14595
R503 VTAIL.n132 VTAIL.n126 8.14595
R504 VTAIL.n353 VTAIL.n347 8.14595
R505 VTAIL.n297 VTAIL.n291 8.14595
R506 VTAIL.n243 VTAIL.n237 8.14595
R507 VTAIL.n187 VTAIL.n181 8.14595
R508 VTAIL.n405 VTAIL.n402 7.3702
R509 VTAIL.n21 VTAIL.n18 7.3702
R510 VTAIL.n75 VTAIL.n72 7.3702
R511 VTAIL.n131 VTAIL.n128 7.3702
R512 VTAIL.n352 VTAIL.n349 7.3702
R513 VTAIL.n296 VTAIL.n293 7.3702
R514 VTAIL.n242 VTAIL.n239 7.3702
R515 VTAIL.n186 VTAIL.n183 7.3702
R516 VTAIL.n406 VTAIL.n405 5.81868
R517 VTAIL.n22 VTAIL.n21 5.81868
R518 VTAIL.n76 VTAIL.n75 5.81868
R519 VTAIL.n132 VTAIL.n131 5.81868
R520 VTAIL.n353 VTAIL.n352 5.81868
R521 VTAIL.n297 VTAIL.n296 5.81868
R522 VTAIL.n243 VTAIL.n242 5.81868
R523 VTAIL.n187 VTAIL.n186 5.81868
R524 VTAIL.n409 VTAIL.n400 5.04292
R525 VTAIL.n25 VTAIL.n16 5.04292
R526 VTAIL.n79 VTAIL.n70 5.04292
R527 VTAIL.n135 VTAIL.n126 5.04292
R528 VTAIL.n356 VTAIL.n347 5.04292
R529 VTAIL.n300 VTAIL.n291 5.04292
R530 VTAIL.n246 VTAIL.n237 5.04292
R531 VTAIL.n190 VTAIL.n181 5.04292
R532 VTAIL.n410 VTAIL.n398 4.26717
R533 VTAIL.n26 VTAIL.n14 4.26717
R534 VTAIL.n80 VTAIL.n68 4.26717
R535 VTAIL.n136 VTAIL.n124 4.26717
R536 VTAIL.n357 VTAIL.n345 4.26717
R537 VTAIL.n301 VTAIL.n289 4.26717
R538 VTAIL.n247 VTAIL.n235 4.26717
R539 VTAIL.n191 VTAIL.n179 4.26717
R540 VTAIL.n414 VTAIL.n413 3.49141
R541 VTAIL.n438 VTAIL.n386 3.49141
R542 VTAIL.n30 VTAIL.n29 3.49141
R543 VTAIL.n54 VTAIL.n2 3.49141
R544 VTAIL.n84 VTAIL.n83 3.49141
R545 VTAIL.n108 VTAIL.n56 3.49141
R546 VTAIL.n140 VTAIL.n139 3.49141
R547 VTAIL.n164 VTAIL.n112 3.49141
R548 VTAIL.n384 VTAIL.n332 3.49141
R549 VTAIL.n361 VTAIL.n360 3.49141
R550 VTAIL.n328 VTAIL.n276 3.49141
R551 VTAIL.n305 VTAIL.n304 3.49141
R552 VTAIL.n274 VTAIL.n222 3.49141
R553 VTAIL.n251 VTAIL.n250 3.49141
R554 VTAIL.n218 VTAIL.n166 3.49141
R555 VTAIL.n195 VTAIL.n194 3.49141
R556 VTAIL.n404 VTAIL.n403 2.84303
R557 VTAIL.n20 VTAIL.n19 2.84303
R558 VTAIL.n74 VTAIL.n73 2.84303
R559 VTAIL.n130 VTAIL.n129 2.84303
R560 VTAIL.n351 VTAIL.n350 2.84303
R561 VTAIL.n295 VTAIL.n294 2.84303
R562 VTAIL.n241 VTAIL.n240 2.84303
R563 VTAIL.n185 VTAIL.n184 2.84303
R564 VTAIL.n417 VTAIL.n396 2.71565
R565 VTAIL.n436 VTAIL.n435 2.71565
R566 VTAIL.n33 VTAIL.n12 2.71565
R567 VTAIL.n52 VTAIL.n51 2.71565
R568 VTAIL.n87 VTAIL.n66 2.71565
R569 VTAIL.n106 VTAIL.n105 2.71565
R570 VTAIL.n143 VTAIL.n122 2.71565
R571 VTAIL.n162 VTAIL.n161 2.71565
R572 VTAIL.n382 VTAIL.n381 2.71565
R573 VTAIL.n364 VTAIL.n343 2.71565
R574 VTAIL.n326 VTAIL.n325 2.71565
R575 VTAIL.n308 VTAIL.n287 2.71565
R576 VTAIL.n272 VTAIL.n271 2.71565
R577 VTAIL.n254 VTAIL.n233 2.71565
R578 VTAIL.n216 VTAIL.n215 2.71565
R579 VTAIL.n198 VTAIL.n177 2.71565
R580 VTAIL.n0 VTAIL.t14 1.94932
R581 VTAIL.n0 VTAIL.t11 1.94932
R582 VTAIL.n110 VTAIL.t7 1.94932
R583 VTAIL.n110 VTAIL.t1 1.94932
R584 VTAIL.n330 VTAIL.t2 1.94932
R585 VTAIL.n330 VTAIL.t4 1.94932
R586 VTAIL.n220 VTAIL.t10 1.94932
R587 VTAIL.n220 VTAIL.t8 1.94932
R588 VTAIL.n418 VTAIL.n394 1.93989
R589 VTAIL.n432 VTAIL.n388 1.93989
R590 VTAIL.n34 VTAIL.n10 1.93989
R591 VTAIL.n48 VTAIL.n4 1.93989
R592 VTAIL.n88 VTAIL.n64 1.93989
R593 VTAIL.n102 VTAIL.n58 1.93989
R594 VTAIL.n144 VTAIL.n120 1.93989
R595 VTAIL.n158 VTAIL.n114 1.93989
R596 VTAIL.n378 VTAIL.n334 1.93989
R597 VTAIL.n365 VTAIL.n341 1.93989
R598 VTAIL.n322 VTAIL.n278 1.93989
R599 VTAIL.n309 VTAIL.n285 1.93989
R600 VTAIL.n268 VTAIL.n224 1.93989
R601 VTAIL.n255 VTAIL.n231 1.93989
R602 VTAIL.n212 VTAIL.n168 1.93989
R603 VTAIL.n199 VTAIL.n175 1.93989
R604 VTAIL.n221 VTAIL.n219 1.41429
R605 VTAIL.n275 VTAIL.n221 1.41429
R606 VTAIL.n331 VTAIL.n329 1.41429
R607 VTAIL.n385 VTAIL.n331 1.41429
R608 VTAIL.n165 VTAIL.n111 1.41429
R609 VTAIL.n111 VTAIL.n109 1.41429
R610 VTAIL.n55 VTAIL.n1 1.41429
R611 VTAIL VTAIL.n439 1.3561
R612 VTAIL.n423 VTAIL.n421 1.16414
R613 VTAIL.n431 VTAIL.n390 1.16414
R614 VTAIL.n39 VTAIL.n37 1.16414
R615 VTAIL.n47 VTAIL.n6 1.16414
R616 VTAIL.n93 VTAIL.n91 1.16414
R617 VTAIL.n101 VTAIL.n60 1.16414
R618 VTAIL.n149 VTAIL.n147 1.16414
R619 VTAIL.n157 VTAIL.n116 1.16414
R620 VTAIL.n377 VTAIL.n336 1.16414
R621 VTAIL.n369 VTAIL.n368 1.16414
R622 VTAIL.n321 VTAIL.n280 1.16414
R623 VTAIL.n313 VTAIL.n312 1.16414
R624 VTAIL.n267 VTAIL.n226 1.16414
R625 VTAIL.n259 VTAIL.n258 1.16414
R626 VTAIL.n211 VTAIL.n170 1.16414
R627 VTAIL.n203 VTAIL.n202 1.16414
R628 VTAIL.n329 VTAIL.n275 0.470328
R629 VTAIL.n109 VTAIL.n55 0.470328
R630 VTAIL.n422 VTAIL.n392 0.388379
R631 VTAIL.n428 VTAIL.n427 0.388379
R632 VTAIL.n38 VTAIL.n8 0.388379
R633 VTAIL.n44 VTAIL.n43 0.388379
R634 VTAIL.n92 VTAIL.n62 0.388379
R635 VTAIL.n98 VTAIL.n97 0.388379
R636 VTAIL.n148 VTAIL.n118 0.388379
R637 VTAIL.n154 VTAIL.n153 0.388379
R638 VTAIL.n374 VTAIL.n373 0.388379
R639 VTAIL.n340 VTAIL.n338 0.388379
R640 VTAIL.n318 VTAIL.n317 0.388379
R641 VTAIL.n284 VTAIL.n282 0.388379
R642 VTAIL.n264 VTAIL.n263 0.388379
R643 VTAIL.n230 VTAIL.n228 0.388379
R644 VTAIL.n208 VTAIL.n207 0.388379
R645 VTAIL.n174 VTAIL.n172 0.388379
R646 VTAIL.n404 VTAIL.n399 0.155672
R647 VTAIL.n411 VTAIL.n399 0.155672
R648 VTAIL.n412 VTAIL.n411 0.155672
R649 VTAIL.n412 VTAIL.n395 0.155672
R650 VTAIL.n419 VTAIL.n395 0.155672
R651 VTAIL.n420 VTAIL.n419 0.155672
R652 VTAIL.n420 VTAIL.n391 0.155672
R653 VTAIL.n429 VTAIL.n391 0.155672
R654 VTAIL.n430 VTAIL.n429 0.155672
R655 VTAIL.n430 VTAIL.n387 0.155672
R656 VTAIL.n437 VTAIL.n387 0.155672
R657 VTAIL.n20 VTAIL.n15 0.155672
R658 VTAIL.n27 VTAIL.n15 0.155672
R659 VTAIL.n28 VTAIL.n27 0.155672
R660 VTAIL.n28 VTAIL.n11 0.155672
R661 VTAIL.n35 VTAIL.n11 0.155672
R662 VTAIL.n36 VTAIL.n35 0.155672
R663 VTAIL.n36 VTAIL.n7 0.155672
R664 VTAIL.n45 VTAIL.n7 0.155672
R665 VTAIL.n46 VTAIL.n45 0.155672
R666 VTAIL.n46 VTAIL.n3 0.155672
R667 VTAIL.n53 VTAIL.n3 0.155672
R668 VTAIL.n74 VTAIL.n69 0.155672
R669 VTAIL.n81 VTAIL.n69 0.155672
R670 VTAIL.n82 VTAIL.n81 0.155672
R671 VTAIL.n82 VTAIL.n65 0.155672
R672 VTAIL.n89 VTAIL.n65 0.155672
R673 VTAIL.n90 VTAIL.n89 0.155672
R674 VTAIL.n90 VTAIL.n61 0.155672
R675 VTAIL.n99 VTAIL.n61 0.155672
R676 VTAIL.n100 VTAIL.n99 0.155672
R677 VTAIL.n100 VTAIL.n57 0.155672
R678 VTAIL.n107 VTAIL.n57 0.155672
R679 VTAIL.n130 VTAIL.n125 0.155672
R680 VTAIL.n137 VTAIL.n125 0.155672
R681 VTAIL.n138 VTAIL.n137 0.155672
R682 VTAIL.n138 VTAIL.n121 0.155672
R683 VTAIL.n145 VTAIL.n121 0.155672
R684 VTAIL.n146 VTAIL.n145 0.155672
R685 VTAIL.n146 VTAIL.n117 0.155672
R686 VTAIL.n155 VTAIL.n117 0.155672
R687 VTAIL.n156 VTAIL.n155 0.155672
R688 VTAIL.n156 VTAIL.n113 0.155672
R689 VTAIL.n163 VTAIL.n113 0.155672
R690 VTAIL.n383 VTAIL.n333 0.155672
R691 VTAIL.n376 VTAIL.n333 0.155672
R692 VTAIL.n376 VTAIL.n375 0.155672
R693 VTAIL.n375 VTAIL.n337 0.155672
R694 VTAIL.n367 VTAIL.n337 0.155672
R695 VTAIL.n367 VTAIL.n366 0.155672
R696 VTAIL.n366 VTAIL.n342 0.155672
R697 VTAIL.n359 VTAIL.n342 0.155672
R698 VTAIL.n359 VTAIL.n358 0.155672
R699 VTAIL.n358 VTAIL.n346 0.155672
R700 VTAIL.n351 VTAIL.n346 0.155672
R701 VTAIL.n327 VTAIL.n277 0.155672
R702 VTAIL.n320 VTAIL.n277 0.155672
R703 VTAIL.n320 VTAIL.n319 0.155672
R704 VTAIL.n319 VTAIL.n281 0.155672
R705 VTAIL.n311 VTAIL.n281 0.155672
R706 VTAIL.n311 VTAIL.n310 0.155672
R707 VTAIL.n310 VTAIL.n286 0.155672
R708 VTAIL.n303 VTAIL.n286 0.155672
R709 VTAIL.n303 VTAIL.n302 0.155672
R710 VTAIL.n302 VTAIL.n290 0.155672
R711 VTAIL.n295 VTAIL.n290 0.155672
R712 VTAIL.n273 VTAIL.n223 0.155672
R713 VTAIL.n266 VTAIL.n223 0.155672
R714 VTAIL.n266 VTAIL.n265 0.155672
R715 VTAIL.n265 VTAIL.n227 0.155672
R716 VTAIL.n257 VTAIL.n227 0.155672
R717 VTAIL.n257 VTAIL.n256 0.155672
R718 VTAIL.n256 VTAIL.n232 0.155672
R719 VTAIL.n249 VTAIL.n232 0.155672
R720 VTAIL.n249 VTAIL.n248 0.155672
R721 VTAIL.n248 VTAIL.n236 0.155672
R722 VTAIL.n241 VTAIL.n236 0.155672
R723 VTAIL.n217 VTAIL.n167 0.155672
R724 VTAIL.n210 VTAIL.n167 0.155672
R725 VTAIL.n210 VTAIL.n209 0.155672
R726 VTAIL.n209 VTAIL.n171 0.155672
R727 VTAIL.n201 VTAIL.n171 0.155672
R728 VTAIL.n201 VTAIL.n200 0.155672
R729 VTAIL.n200 VTAIL.n176 0.155672
R730 VTAIL.n193 VTAIL.n176 0.155672
R731 VTAIL.n193 VTAIL.n192 0.155672
R732 VTAIL.n192 VTAIL.n180 0.155672
R733 VTAIL.n185 VTAIL.n180 0.155672
R734 VTAIL VTAIL.n1 0.0586897
R735 VDD2.n2 VDD2.n1 67.1705
R736 VDD2.n2 VDD2.n0 67.1705
R737 VDD2 VDD2.n5 67.1676
R738 VDD2.n4 VDD2.n3 66.5191
R739 VDD2.n4 VDD2.n2 38.836
R740 VDD2.n5 VDD2.t4 1.94932
R741 VDD2.n5 VDD2.t2 1.94932
R742 VDD2.n3 VDD2.t0 1.94932
R743 VDD2.n3 VDD2.t1 1.94932
R744 VDD2.n1 VDD2.t5 1.94932
R745 VDD2.n1 VDD2.t7 1.94932
R746 VDD2.n0 VDD2.t6 1.94932
R747 VDD2.n0 VDD2.t3 1.94932
R748 VDD2 VDD2.n4 0.765586
R749 B.n678 B.n677 585
R750 B.n267 B.n102 585
R751 B.n266 B.n265 585
R752 B.n264 B.n263 585
R753 B.n262 B.n261 585
R754 B.n260 B.n259 585
R755 B.n258 B.n257 585
R756 B.n256 B.n255 585
R757 B.n254 B.n253 585
R758 B.n252 B.n251 585
R759 B.n250 B.n249 585
R760 B.n248 B.n247 585
R761 B.n246 B.n245 585
R762 B.n244 B.n243 585
R763 B.n242 B.n241 585
R764 B.n240 B.n239 585
R765 B.n238 B.n237 585
R766 B.n236 B.n235 585
R767 B.n234 B.n233 585
R768 B.n232 B.n231 585
R769 B.n230 B.n229 585
R770 B.n228 B.n227 585
R771 B.n226 B.n225 585
R772 B.n224 B.n223 585
R773 B.n222 B.n221 585
R774 B.n220 B.n219 585
R775 B.n218 B.n217 585
R776 B.n216 B.n215 585
R777 B.n214 B.n213 585
R778 B.n212 B.n211 585
R779 B.n210 B.n209 585
R780 B.n208 B.n207 585
R781 B.n206 B.n205 585
R782 B.n204 B.n203 585
R783 B.n202 B.n201 585
R784 B.n200 B.n199 585
R785 B.n198 B.n197 585
R786 B.n196 B.n195 585
R787 B.n194 B.n193 585
R788 B.n192 B.n191 585
R789 B.n190 B.n189 585
R790 B.n188 B.n187 585
R791 B.n186 B.n185 585
R792 B.n184 B.n183 585
R793 B.n182 B.n181 585
R794 B.n180 B.n179 585
R795 B.n178 B.n177 585
R796 B.n176 B.n175 585
R797 B.n174 B.n173 585
R798 B.n172 B.n171 585
R799 B.n170 B.n169 585
R800 B.n168 B.n167 585
R801 B.n166 B.n165 585
R802 B.n164 B.n163 585
R803 B.n162 B.n161 585
R804 B.n160 B.n159 585
R805 B.n158 B.n157 585
R806 B.n156 B.n155 585
R807 B.n154 B.n153 585
R808 B.n152 B.n151 585
R809 B.n150 B.n149 585
R810 B.n148 B.n147 585
R811 B.n146 B.n145 585
R812 B.n144 B.n143 585
R813 B.n142 B.n141 585
R814 B.n140 B.n139 585
R815 B.n138 B.n137 585
R816 B.n136 B.n135 585
R817 B.n134 B.n133 585
R818 B.n132 B.n131 585
R819 B.n130 B.n129 585
R820 B.n128 B.n127 585
R821 B.n126 B.n125 585
R822 B.n124 B.n123 585
R823 B.n122 B.n121 585
R824 B.n120 B.n119 585
R825 B.n118 B.n117 585
R826 B.n116 B.n115 585
R827 B.n114 B.n113 585
R828 B.n112 B.n111 585
R829 B.n110 B.n109 585
R830 B.n60 B.n59 585
R831 B.n676 B.n61 585
R832 B.n681 B.n61 585
R833 B.n675 B.n674 585
R834 B.n674 B.n57 585
R835 B.n673 B.n56 585
R836 B.n687 B.n56 585
R837 B.n672 B.n55 585
R838 B.n688 B.n55 585
R839 B.n671 B.n54 585
R840 B.n689 B.n54 585
R841 B.n670 B.n669 585
R842 B.n669 B.n53 585
R843 B.n668 B.n49 585
R844 B.n695 B.n49 585
R845 B.n667 B.n48 585
R846 B.n696 B.n48 585
R847 B.n666 B.n47 585
R848 B.n697 B.n47 585
R849 B.n665 B.n664 585
R850 B.n664 B.n43 585
R851 B.n663 B.n42 585
R852 B.n703 B.n42 585
R853 B.n662 B.n41 585
R854 B.n704 B.n41 585
R855 B.n661 B.n40 585
R856 B.n705 B.n40 585
R857 B.n660 B.n659 585
R858 B.n659 B.n39 585
R859 B.n658 B.n35 585
R860 B.n711 B.n35 585
R861 B.n657 B.n34 585
R862 B.n712 B.n34 585
R863 B.n656 B.n33 585
R864 B.n713 B.n33 585
R865 B.n655 B.n654 585
R866 B.n654 B.n29 585
R867 B.n653 B.n28 585
R868 B.n719 B.n28 585
R869 B.n652 B.n27 585
R870 B.n720 B.n27 585
R871 B.n651 B.n26 585
R872 B.n721 B.n26 585
R873 B.n650 B.n649 585
R874 B.n649 B.n22 585
R875 B.n648 B.n21 585
R876 B.n727 B.n21 585
R877 B.n647 B.n20 585
R878 B.n728 B.n20 585
R879 B.n646 B.n19 585
R880 B.n729 B.n19 585
R881 B.n645 B.n644 585
R882 B.n644 B.n15 585
R883 B.n643 B.n14 585
R884 B.n735 B.n14 585
R885 B.n642 B.n13 585
R886 B.n736 B.n13 585
R887 B.n641 B.n12 585
R888 B.n737 B.n12 585
R889 B.n640 B.n639 585
R890 B.n639 B.n8 585
R891 B.n638 B.n7 585
R892 B.n743 B.n7 585
R893 B.n637 B.n6 585
R894 B.n744 B.n6 585
R895 B.n636 B.n5 585
R896 B.n745 B.n5 585
R897 B.n635 B.n634 585
R898 B.n634 B.n4 585
R899 B.n633 B.n268 585
R900 B.n633 B.n632 585
R901 B.n623 B.n269 585
R902 B.n270 B.n269 585
R903 B.n625 B.n624 585
R904 B.n626 B.n625 585
R905 B.n622 B.n274 585
R906 B.n278 B.n274 585
R907 B.n621 B.n620 585
R908 B.n620 B.n619 585
R909 B.n276 B.n275 585
R910 B.n277 B.n276 585
R911 B.n612 B.n611 585
R912 B.n613 B.n612 585
R913 B.n610 B.n282 585
R914 B.n286 B.n282 585
R915 B.n609 B.n608 585
R916 B.n608 B.n607 585
R917 B.n284 B.n283 585
R918 B.n285 B.n284 585
R919 B.n600 B.n599 585
R920 B.n601 B.n600 585
R921 B.n598 B.n291 585
R922 B.n291 B.n290 585
R923 B.n597 B.n596 585
R924 B.n596 B.n595 585
R925 B.n293 B.n292 585
R926 B.n294 B.n293 585
R927 B.n588 B.n587 585
R928 B.n589 B.n588 585
R929 B.n586 B.n299 585
R930 B.n299 B.n298 585
R931 B.n585 B.n584 585
R932 B.n584 B.n583 585
R933 B.n301 B.n300 585
R934 B.n576 B.n301 585
R935 B.n575 B.n574 585
R936 B.n577 B.n575 585
R937 B.n573 B.n306 585
R938 B.n306 B.n305 585
R939 B.n572 B.n571 585
R940 B.n571 B.n570 585
R941 B.n308 B.n307 585
R942 B.n309 B.n308 585
R943 B.n563 B.n562 585
R944 B.n564 B.n563 585
R945 B.n561 B.n314 585
R946 B.n314 B.n313 585
R947 B.n560 B.n559 585
R948 B.n559 B.n558 585
R949 B.n316 B.n315 585
R950 B.n551 B.n316 585
R951 B.n550 B.n549 585
R952 B.n552 B.n550 585
R953 B.n548 B.n321 585
R954 B.n321 B.n320 585
R955 B.n547 B.n546 585
R956 B.n546 B.n545 585
R957 B.n323 B.n322 585
R958 B.n324 B.n323 585
R959 B.n538 B.n537 585
R960 B.n539 B.n538 585
R961 B.n327 B.n326 585
R962 B.n374 B.n372 585
R963 B.n375 B.n371 585
R964 B.n375 B.n328 585
R965 B.n378 B.n377 585
R966 B.n379 B.n370 585
R967 B.n381 B.n380 585
R968 B.n383 B.n369 585
R969 B.n386 B.n385 585
R970 B.n387 B.n368 585
R971 B.n389 B.n388 585
R972 B.n391 B.n367 585
R973 B.n394 B.n393 585
R974 B.n395 B.n366 585
R975 B.n397 B.n396 585
R976 B.n399 B.n365 585
R977 B.n402 B.n401 585
R978 B.n403 B.n364 585
R979 B.n405 B.n404 585
R980 B.n407 B.n363 585
R981 B.n410 B.n409 585
R982 B.n411 B.n362 585
R983 B.n413 B.n412 585
R984 B.n415 B.n361 585
R985 B.n418 B.n417 585
R986 B.n419 B.n360 585
R987 B.n421 B.n420 585
R988 B.n423 B.n359 585
R989 B.n426 B.n425 585
R990 B.n427 B.n358 585
R991 B.n429 B.n428 585
R992 B.n431 B.n357 585
R993 B.n434 B.n433 585
R994 B.n435 B.n356 585
R995 B.n437 B.n436 585
R996 B.n439 B.n355 585
R997 B.n442 B.n441 585
R998 B.n444 B.n352 585
R999 B.n446 B.n445 585
R1000 B.n448 B.n351 585
R1001 B.n451 B.n450 585
R1002 B.n452 B.n350 585
R1003 B.n454 B.n453 585
R1004 B.n456 B.n349 585
R1005 B.n459 B.n458 585
R1006 B.n460 B.n348 585
R1007 B.n465 B.n464 585
R1008 B.n467 B.n347 585
R1009 B.n470 B.n469 585
R1010 B.n471 B.n346 585
R1011 B.n473 B.n472 585
R1012 B.n475 B.n345 585
R1013 B.n478 B.n477 585
R1014 B.n479 B.n344 585
R1015 B.n481 B.n480 585
R1016 B.n483 B.n343 585
R1017 B.n486 B.n485 585
R1018 B.n487 B.n342 585
R1019 B.n489 B.n488 585
R1020 B.n491 B.n341 585
R1021 B.n494 B.n493 585
R1022 B.n495 B.n340 585
R1023 B.n497 B.n496 585
R1024 B.n499 B.n339 585
R1025 B.n502 B.n501 585
R1026 B.n503 B.n338 585
R1027 B.n505 B.n504 585
R1028 B.n507 B.n337 585
R1029 B.n510 B.n509 585
R1030 B.n511 B.n336 585
R1031 B.n513 B.n512 585
R1032 B.n515 B.n335 585
R1033 B.n518 B.n517 585
R1034 B.n519 B.n334 585
R1035 B.n521 B.n520 585
R1036 B.n523 B.n333 585
R1037 B.n526 B.n525 585
R1038 B.n527 B.n332 585
R1039 B.n529 B.n528 585
R1040 B.n531 B.n331 585
R1041 B.n532 B.n330 585
R1042 B.n535 B.n534 585
R1043 B.n536 B.n329 585
R1044 B.n329 B.n328 585
R1045 B.n541 B.n540 585
R1046 B.n540 B.n539 585
R1047 B.n542 B.n325 585
R1048 B.n325 B.n324 585
R1049 B.n544 B.n543 585
R1050 B.n545 B.n544 585
R1051 B.n319 B.n318 585
R1052 B.n320 B.n319 585
R1053 B.n554 B.n553 585
R1054 B.n553 B.n552 585
R1055 B.n555 B.n317 585
R1056 B.n551 B.n317 585
R1057 B.n557 B.n556 585
R1058 B.n558 B.n557 585
R1059 B.n312 B.n311 585
R1060 B.n313 B.n312 585
R1061 B.n566 B.n565 585
R1062 B.n565 B.n564 585
R1063 B.n567 B.n310 585
R1064 B.n310 B.n309 585
R1065 B.n569 B.n568 585
R1066 B.n570 B.n569 585
R1067 B.n304 B.n303 585
R1068 B.n305 B.n304 585
R1069 B.n579 B.n578 585
R1070 B.n578 B.n577 585
R1071 B.n580 B.n302 585
R1072 B.n576 B.n302 585
R1073 B.n582 B.n581 585
R1074 B.n583 B.n582 585
R1075 B.n297 B.n296 585
R1076 B.n298 B.n297 585
R1077 B.n591 B.n590 585
R1078 B.n590 B.n589 585
R1079 B.n592 B.n295 585
R1080 B.n295 B.n294 585
R1081 B.n594 B.n593 585
R1082 B.n595 B.n594 585
R1083 B.n289 B.n288 585
R1084 B.n290 B.n289 585
R1085 B.n603 B.n602 585
R1086 B.n602 B.n601 585
R1087 B.n604 B.n287 585
R1088 B.n287 B.n285 585
R1089 B.n606 B.n605 585
R1090 B.n607 B.n606 585
R1091 B.n281 B.n280 585
R1092 B.n286 B.n281 585
R1093 B.n615 B.n614 585
R1094 B.n614 B.n613 585
R1095 B.n616 B.n279 585
R1096 B.n279 B.n277 585
R1097 B.n618 B.n617 585
R1098 B.n619 B.n618 585
R1099 B.n273 B.n272 585
R1100 B.n278 B.n273 585
R1101 B.n628 B.n627 585
R1102 B.n627 B.n626 585
R1103 B.n629 B.n271 585
R1104 B.n271 B.n270 585
R1105 B.n631 B.n630 585
R1106 B.n632 B.n631 585
R1107 B.n2 B.n0 585
R1108 B.n4 B.n2 585
R1109 B.n3 B.n1 585
R1110 B.n744 B.n3 585
R1111 B.n742 B.n741 585
R1112 B.n743 B.n742 585
R1113 B.n740 B.n9 585
R1114 B.n9 B.n8 585
R1115 B.n739 B.n738 585
R1116 B.n738 B.n737 585
R1117 B.n11 B.n10 585
R1118 B.n736 B.n11 585
R1119 B.n734 B.n733 585
R1120 B.n735 B.n734 585
R1121 B.n732 B.n16 585
R1122 B.n16 B.n15 585
R1123 B.n731 B.n730 585
R1124 B.n730 B.n729 585
R1125 B.n18 B.n17 585
R1126 B.n728 B.n18 585
R1127 B.n726 B.n725 585
R1128 B.n727 B.n726 585
R1129 B.n724 B.n23 585
R1130 B.n23 B.n22 585
R1131 B.n723 B.n722 585
R1132 B.n722 B.n721 585
R1133 B.n25 B.n24 585
R1134 B.n720 B.n25 585
R1135 B.n718 B.n717 585
R1136 B.n719 B.n718 585
R1137 B.n716 B.n30 585
R1138 B.n30 B.n29 585
R1139 B.n715 B.n714 585
R1140 B.n714 B.n713 585
R1141 B.n32 B.n31 585
R1142 B.n712 B.n32 585
R1143 B.n710 B.n709 585
R1144 B.n711 B.n710 585
R1145 B.n708 B.n36 585
R1146 B.n39 B.n36 585
R1147 B.n707 B.n706 585
R1148 B.n706 B.n705 585
R1149 B.n38 B.n37 585
R1150 B.n704 B.n38 585
R1151 B.n702 B.n701 585
R1152 B.n703 B.n702 585
R1153 B.n700 B.n44 585
R1154 B.n44 B.n43 585
R1155 B.n699 B.n698 585
R1156 B.n698 B.n697 585
R1157 B.n46 B.n45 585
R1158 B.n696 B.n46 585
R1159 B.n694 B.n693 585
R1160 B.n695 B.n694 585
R1161 B.n692 B.n50 585
R1162 B.n53 B.n50 585
R1163 B.n691 B.n690 585
R1164 B.n690 B.n689 585
R1165 B.n52 B.n51 585
R1166 B.n688 B.n52 585
R1167 B.n686 B.n685 585
R1168 B.n687 B.n686 585
R1169 B.n684 B.n58 585
R1170 B.n58 B.n57 585
R1171 B.n683 B.n682 585
R1172 B.n682 B.n681 585
R1173 B.n747 B.n746 585
R1174 B.n746 B.n745 585
R1175 B.n540 B.n327 535.745
R1176 B.n682 B.n60 535.745
R1177 B.n538 B.n329 535.745
R1178 B.n678 B.n61 535.745
R1179 B.n461 B.t19 391.568
R1180 B.n353 B.t15 391.568
R1181 B.n106 B.t12 391.568
R1182 B.n103 B.t8 391.568
R1183 B.n461 B.t21 282.557
R1184 B.n103 B.t10 282.557
R1185 B.n353 B.t18 282.557
R1186 B.n106 B.t13 282.557
R1187 B.n680 B.n679 256.663
R1188 B.n680 B.n101 256.663
R1189 B.n680 B.n100 256.663
R1190 B.n680 B.n99 256.663
R1191 B.n680 B.n98 256.663
R1192 B.n680 B.n97 256.663
R1193 B.n680 B.n96 256.663
R1194 B.n680 B.n95 256.663
R1195 B.n680 B.n94 256.663
R1196 B.n680 B.n93 256.663
R1197 B.n680 B.n92 256.663
R1198 B.n680 B.n91 256.663
R1199 B.n680 B.n90 256.663
R1200 B.n680 B.n89 256.663
R1201 B.n680 B.n88 256.663
R1202 B.n680 B.n87 256.663
R1203 B.n680 B.n86 256.663
R1204 B.n680 B.n85 256.663
R1205 B.n680 B.n84 256.663
R1206 B.n680 B.n83 256.663
R1207 B.n680 B.n82 256.663
R1208 B.n680 B.n81 256.663
R1209 B.n680 B.n80 256.663
R1210 B.n680 B.n79 256.663
R1211 B.n680 B.n78 256.663
R1212 B.n680 B.n77 256.663
R1213 B.n680 B.n76 256.663
R1214 B.n680 B.n75 256.663
R1215 B.n680 B.n74 256.663
R1216 B.n680 B.n73 256.663
R1217 B.n680 B.n72 256.663
R1218 B.n680 B.n71 256.663
R1219 B.n680 B.n70 256.663
R1220 B.n680 B.n69 256.663
R1221 B.n680 B.n68 256.663
R1222 B.n680 B.n67 256.663
R1223 B.n680 B.n66 256.663
R1224 B.n680 B.n65 256.663
R1225 B.n680 B.n64 256.663
R1226 B.n680 B.n63 256.663
R1227 B.n680 B.n62 256.663
R1228 B.n373 B.n328 256.663
R1229 B.n376 B.n328 256.663
R1230 B.n382 B.n328 256.663
R1231 B.n384 B.n328 256.663
R1232 B.n390 B.n328 256.663
R1233 B.n392 B.n328 256.663
R1234 B.n398 B.n328 256.663
R1235 B.n400 B.n328 256.663
R1236 B.n406 B.n328 256.663
R1237 B.n408 B.n328 256.663
R1238 B.n414 B.n328 256.663
R1239 B.n416 B.n328 256.663
R1240 B.n422 B.n328 256.663
R1241 B.n424 B.n328 256.663
R1242 B.n430 B.n328 256.663
R1243 B.n432 B.n328 256.663
R1244 B.n438 B.n328 256.663
R1245 B.n440 B.n328 256.663
R1246 B.n447 B.n328 256.663
R1247 B.n449 B.n328 256.663
R1248 B.n455 B.n328 256.663
R1249 B.n457 B.n328 256.663
R1250 B.n466 B.n328 256.663
R1251 B.n468 B.n328 256.663
R1252 B.n474 B.n328 256.663
R1253 B.n476 B.n328 256.663
R1254 B.n482 B.n328 256.663
R1255 B.n484 B.n328 256.663
R1256 B.n490 B.n328 256.663
R1257 B.n492 B.n328 256.663
R1258 B.n498 B.n328 256.663
R1259 B.n500 B.n328 256.663
R1260 B.n506 B.n328 256.663
R1261 B.n508 B.n328 256.663
R1262 B.n514 B.n328 256.663
R1263 B.n516 B.n328 256.663
R1264 B.n522 B.n328 256.663
R1265 B.n524 B.n328 256.663
R1266 B.n530 B.n328 256.663
R1267 B.n533 B.n328 256.663
R1268 B.n462 B.t20 250.75
R1269 B.n104 B.t11 250.75
R1270 B.n354 B.t17 250.75
R1271 B.n107 B.t14 250.75
R1272 B.n540 B.n325 163.367
R1273 B.n544 B.n325 163.367
R1274 B.n544 B.n319 163.367
R1275 B.n553 B.n319 163.367
R1276 B.n553 B.n317 163.367
R1277 B.n557 B.n317 163.367
R1278 B.n557 B.n312 163.367
R1279 B.n565 B.n312 163.367
R1280 B.n565 B.n310 163.367
R1281 B.n569 B.n310 163.367
R1282 B.n569 B.n304 163.367
R1283 B.n578 B.n304 163.367
R1284 B.n578 B.n302 163.367
R1285 B.n582 B.n302 163.367
R1286 B.n582 B.n297 163.367
R1287 B.n590 B.n297 163.367
R1288 B.n590 B.n295 163.367
R1289 B.n594 B.n295 163.367
R1290 B.n594 B.n289 163.367
R1291 B.n602 B.n289 163.367
R1292 B.n602 B.n287 163.367
R1293 B.n606 B.n287 163.367
R1294 B.n606 B.n281 163.367
R1295 B.n614 B.n281 163.367
R1296 B.n614 B.n279 163.367
R1297 B.n618 B.n279 163.367
R1298 B.n618 B.n273 163.367
R1299 B.n627 B.n273 163.367
R1300 B.n627 B.n271 163.367
R1301 B.n631 B.n271 163.367
R1302 B.n631 B.n2 163.367
R1303 B.n746 B.n2 163.367
R1304 B.n746 B.n3 163.367
R1305 B.n742 B.n3 163.367
R1306 B.n742 B.n9 163.367
R1307 B.n738 B.n9 163.367
R1308 B.n738 B.n11 163.367
R1309 B.n734 B.n11 163.367
R1310 B.n734 B.n16 163.367
R1311 B.n730 B.n16 163.367
R1312 B.n730 B.n18 163.367
R1313 B.n726 B.n18 163.367
R1314 B.n726 B.n23 163.367
R1315 B.n722 B.n23 163.367
R1316 B.n722 B.n25 163.367
R1317 B.n718 B.n25 163.367
R1318 B.n718 B.n30 163.367
R1319 B.n714 B.n30 163.367
R1320 B.n714 B.n32 163.367
R1321 B.n710 B.n32 163.367
R1322 B.n710 B.n36 163.367
R1323 B.n706 B.n36 163.367
R1324 B.n706 B.n38 163.367
R1325 B.n702 B.n38 163.367
R1326 B.n702 B.n44 163.367
R1327 B.n698 B.n44 163.367
R1328 B.n698 B.n46 163.367
R1329 B.n694 B.n46 163.367
R1330 B.n694 B.n50 163.367
R1331 B.n690 B.n50 163.367
R1332 B.n690 B.n52 163.367
R1333 B.n686 B.n52 163.367
R1334 B.n686 B.n58 163.367
R1335 B.n682 B.n58 163.367
R1336 B.n375 B.n374 163.367
R1337 B.n377 B.n375 163.367
R1338 B.n381 B.n370 163.367
R1339 B.n385 B.n383 163.367
R1340 B.n389 B.n368 163.367
R1341 B.n393 B.n391 163.367
R1342 B.n397 B.n366 163.367
R1343 B.n401 B.n399 163.367
R1344 B.n405 B.n364 163.367
R1345 B.n409 B.n407 163.367
R1346 B.n413 B.n362 163.367
R1347 B.n417 B.n415 163.367
R1348 B.n421 B.n360 163.367
R1349 B.n425 B.n423 163.367
R1350 B.n429 B.n358 163.367
R1351 B.n433 B.n431 163.367
R1352 B.n437 B.n356 163.367
R1353 B.n441 B.n439 163.367
R1354 B.n446 B.n352 163.367
R1355 B.n450 B.n448 163.367
R1356 B.n454 B.n350 163.367
R1357 B.n458 B.n456 163.367
R1358 B.n465 B.n348 163.367
R1359 B.n469 B.n467 163.367
R1360 B.n473 B.n346 163.367
R1361 B.n477 B.n475 163.367
R1362 B.n481 B.n344 163.367
R1363 B.n485 B.n483 163.367
R1364 B.n489 B.n342 163.367
R1365 B.n493 B.n491 163.367
R1366 B.n497 B.n340 163.367
R1367 B.n501 B.n499 163.367
R1368 B.n505 B.n338 163.367
R1369 B.n509 B.n507 163.367
R1370 B.n513 B.n336 163.367
R1371 B.n517 B.n515 163.367
R1372 B.n521 B.n334 163.367
R1373 B.n525 B.n523 163.367
R1374 B.n529 B.n332 163.367
R1375 B.n532 B.n531 163.367
R1376 B.n534 B.n329 163.367
R1377 B.n538 B.n323 163.367
R1378 B.n546 B.n323 163.367
R1379 B.n546 B.n321 163.367
R1380 B.n550 B.n321 163.367
R1381 B.n550 B.n316 163.367
R1382 B.n559 B.n316 163.367
R1383 B.n559 B.n314 163.367
R1384 B.n563 B.n314 163.367
R1385 B.n563 B.n308 163.367
R1386 B.n571 B.n308 163.367
R1387 B.n571 B.n306 163.367
R1388 B.n575 B.n306 163.367
R1389 B.n575 B.n301 163.367
R1390 B.n584 B.n301 163.367
R1391 B.n584 B.n299 163.367
R1392 B.n588 B.n299 163.367
R1393 B.n588 B.n293 163.367
R1394 B.n596 B.n293 163.367
R1395 B.n596 B.n291 163.367
R1396 B.n600 B.n291 163.367
R1397 B.n600 B.n284 163.367
R1398 B.n608 B.n284 163.367
R1399 B.n608 B.n282 163.367
R1400 B.n612 B.n282 163.367
R1401 B.n612 B.n276 163.367
R1402 B.n620 B.n276 163.367
R1403 B.n620 B.n274 163.367
R1404 B.n625 B.n274 163.367
R1405 B.n625 B.n269 163.367
R1406 B.n633 B.n269 163.367
R1407 B.n634 B.n633 163.367
R1408 B.n634 B.n5 163.367
R1409 B.n6 B.n5 163.367
R1410 B.n7 B.n6 163.367
R1411 B.n639 B.n7 163.367
R1412 B.n639 B.n12 163.367
R1413 B.n13 B.n12 163.367
R1414 B.n14 B.n13 163.367
R1415 B.n644 B.n14 163.367
R1416 B.n644 B.n19 163.367
R1417 B.n20 B.n19 163.367
R1418 B.n21 B.n20 163.367
R1419 B.n649 B.n21 163.367
R1420 B.n649 B.n26 163.367
R1421 B.n27 B.n26 163.367
R1422 B.n28 B.n27 163.367
R1423 B.n654 B.n28 163.367
R1424 B.n654 B.n33 163.367
R1425 B.n34 B.n33 163.367
R1426 B.n35 B.n34 163.367
R1427 B.n659 B.n35 163.367
R1428 B.n659 B.n40 163.367
R1429 B.n41 B.n40 163.367
R1430 B.n42 B.n41 163.367
R1431 B.n664 B.n42 163.367
R1432 B.n664 B.n47 163.367
R1433 B.n48 B.n47 163.367
R1434 B.n49 B.n48 163.367
R1435 B.n669 B.n49 163.367
R1436 B.n669 B.n54 163.367
R1437 B.n55 B.n54 163.367
R1438 B.n56 B.n55 163.367
R1439 B.n674 B.n56 163.367
R1440 B.n674 B.n61 163.367
R1441 B.n111 B.n110 163.367
R1442 B.n115 B.n114 163.367
R1443 B.n119 B.n118 163.367
R1444 B.n123 B.n122 163.367
R1445 B.n127 B.n126 163.367
R1446 B.n131 B.n130 163.367
R1447 B.n135 B.n134 163.367
R1448 B.n139 B.n138 163.367
R1449 B.n143 B.n142 163.367
R1450 B.n147 B.n146 163.367
R1451 B.n151 B.n150 163.367
R1452 B.n155 B.n154 163.367
R1453 B.n159 B.n158 163.367
R1454 B.n163 B.n162 163.367
R1455 B.n167 B.n166 163.367
R1456 B.n171 B.n170 163.367
R1457 B.n175 B.n174 163.367
R1458 B.n179 B.n178 163.367
R1459 B.n183 B.n182 163.367
R1460 B.n187 B.n186 163.367
R1461 B.n191 B.n190 163.367
R1462 B.n195 B.n194 163.367
R1463 B.n199 B.n198 163.367
R1464 B.n203 B.n202 163.367
R1465 B.n207 B.n206 163.367
R1466 B.n211 B.n210 163.367
R1467 B.n215 B.n214 163.367
R1468 B.n219 B.n218 163.367
R1469 B.n223 B.n222 163.367
R1470 B.n227 B.n226 163.367
R1471 B.n231 B.n230 163.367
R1472 B.n235 B.n234 163.367
R1473 B.n239 B.n238 163.367
R1474 B.n243 B.n242 163.367
R1475 B.n247 B.n246 163.367
R1476 B.n251 B.n250 163.367
R1477 B.n255 B.n254 163.367
R1478 B.n259 B.n258 163.367
R1479 B.n263 B.n262 163.367
R1480 B.n265 B.n102 163.367
R1481 B.n539 B.n328 99.0611
R1482 B.n681 B.n680 99.0611
R1483 B.n373 B.n327 71.676
R1484 B.n377 B.n376 71.676
R1485 B.n382 B.n381 71.676
R1486 B.n385 B.n384 71.676
R1487 B.n390 B.n389 71.676
R1488 B.n393 B.n392 71.676
R1489 B.n398 B.n397 71.676
R1490 B.n401 B.n400 71.676
R1491 B.n406 B.n405 71.676
R1492 B.n409 B.n408 71.676
R1493 B.n414 B.n413 71.676
R1494 B.n417 B.n416 71.676
R1495 B.n422 B.n421 71.676
R1496 B.n425 B.n424 71.676
R1497 B.n430 B.n429 71.676
R1498 B.n433 B.n432 71.676
R1499 B.n438 B.n437 71.676
R1500 B.n441 B.n440 71.676
R1501 B.n447 B.n446 71.676
R1502 B.n450 B.n449 71.676
R1503 B.n455 B.n454 71.676
R1504 B.n458 B.n457 71.676
R1505 B.n466 B.n465 71.676
R1506 B.n469 B.n468 71.676
R1507 B.n474 B.n473 71.676
R1508 B.n477 B.n476 71.676
R1509 B.n482 B.n481 71.676
R1510 B.n485 B.n484 71.676
R1511 B.n490 B.n489 71.676
R1512 B.n493 B.n492 71.676
R1513 B.n498 B.n497 71.676
R1514 B.n501 B.n500 71.676
R1515 B.n506 B.n505 71.676
R1516 B.n509 B.n508 71.676
R1517 B.n514 B.n513 71.676
R1518 B.n517 B.n516 71.676
R1519 B.n522 B.n521 71.676
R1520 B.n525 B.n524 71.676
R1521 B.n530 B.n529 71.676
R1522 B.n533 B.n532 71.676
R1523 B.n62 B.n60 71.676
R1524 B.n111 B.n63 71.676
R1525 B.n115 B.n64 71.676
R1526 B.n119 B.n65 71.676
R1527 B.n123 B.n66 71.676
R1528 B.n127 B.n67 71.676
R1529 B.n131 B.n68 71.676
R1530 B.n135 B.n69 71.676
R1531 B.n139 B.n70 71.676
R1532 B.n143 B.n71 71.676
R1533 B.n147 B.n72 71.676
R1534 B.n151 B.n73 71.676
R1535 B.n155 B.n74 71.676
R1536 B.n159 B.n75 71.676
R1537 B.n163 B.n76 71.676
R1538 B.n167 B.n77 71.676
R1539 B.n171 B.n78 71.676
R1540 B.n175 B.n79 71.676
R1541 B.n179 B.n80 71.676
R1542 B.n183 B.n81 71.676
R1543 B.n187 B.n82 71.676
R1544 B.n191 B.n83 71.676
R1545 B.n195 B.n84 71.676
R1546 B.n199 B.n85 71.676
R1547 B.n203 B.n86 71.676
R1548 B.n207 B.n87 71.676
R1549 B.n211 B.n88 71.676
R1550 B.n215 B.n89 71.676
R1551 B.n219 B.n90 71.676
R1552 B.n223 B.n91 71.676
R1553 B.n227 B.n92 71.676
R1554 B.n231 B.n93 71.676
R1555 B.n235 B.n94 71.676
R1556 B.n239 B.n95 71.676
R1557 B.n243 B.n96 71.676
R1558 B.n247 B.n97 71.676
R1559 B.n251 B.n98 71.676
R1560 B.n255 B.n99 71.676
R1561 B.n259 B.n100 71.676
R1562 B.n263 B.n101 71.676
R1563 B.n679 B.n102 71.676
R1564 B.n679 B.n678 71.676
R1565 B.n265 B.n101 71.676
R1566 B.n262 B.n100 71.676
R1567 B.n258 B.n99 71.676
R1568 B.n254 B.n98 71.676
R1569 B.n250 B.n97 71.676
R1570 B.n246 B.n96 71.676
R1571 B.n242 B.n95 71.676
R1572 B.n238 B.n94 71.676
R1573 B.n234 B.n93 71.676
R1574 B.n230 B.n92 71.676
R1575 B.n226 B.n91 71.676
R1576 B.n222 B.n90 71.676
R1577 B.n218 B.n89 71.676
R1578 B.n214 B.n88 71.676
R1579 B.n210 B.n87 71.676
R1580 B.n206 B.n86 71.676
R1581 B.n202 B.n85 71.676
R1582 B.n198 B.n84 71.676
R1583 B.n194 B.n83 71.676
R1584 B.n190 B.n82 71.676
R1585 B.n186 B.n81 71.676
R1586 B.n182 B.n80 71.676
R1587 B.n178 B.n79 71.676
R1588 B.n174 B.n78 71.676
R1589 B.n170 B.n77 71.676
R1590 B.n166 B.n76 71.676
R1591 B.n162 B.n75 71.676
R1592 B.n158 B.n74 71.676
R1593 B.n154 B.n73 71.676
R1594 B.n150 B.n72 71.676
R1595 B.n146 B.n71 71.676
R1596 B.n142 B.n70 71.676
R1597 B.n138 B.n69 71.676
R1598 B.n134 B.n68 71.676
R1599 B.n130 B.n67 71.676
R1600 B.n126 B.n66 71.676
R1601 B.n122 B.n65 71.676
R1602 B.n118 B.n64 71.676
R1603 B.n114 B.n63 71.676
R1604 B.n110 B.n62 71.676
R1605 B.n374 B.n373 71.676
R1606 B.n376 B.n370 71.676
R1607 B.n383 B.n382 71.676
R1608 B.n384 B.n368 71.676
R1609 B.n391 B.n390 71.676
R1610 B.n392 B.n366 71.676
R1611 B.n399 B.n398 71.676
R1612 B.n400 B.n364 71.676
R1613 B.n407 B.n406 71.676
R1614 B.n408 B.n362 71.676
R1615 B.n415 B.n414 71.676
R1616 B.n416 B.n360 71.676
R1617 B.n423 B.n422 71.676
R1618 B.n424 B.n358 71.676
R1619 B.n431 B.n430 71.676
R1620 B.n432 B.n356 71.676
R1621 B.n439 B.n438 71.676
R1622 B.n440 B.n352 71.676
R1623 B.n448 B.n447 71.676
R1624 B.n449 B.n350 71.676
R1625 B.n456 B.n455 71.676
R1626 B.n457 B.n348 71.676
R1627 B.n467 B.n466 71.676
R1628 B.n468 B.n346 71.676
R1629 B.n475 B.n474 71.676
R1630 B.n476 B.n344 71.676
R1631 B.n483 B.n482 71.676
R1632 B.n484 B.n342 71.676
R1633 B.n491 B.n490 71.676
R1634 B.n492 B.n340 71.676
R1635 B.n499 B.n498 71.676
R1636 B.n500 B.n338 71.676
R1637 B.n507 B.n506 71.676
R1638 B.n508 B.n336 71.676
R1639 B.n515 B.n514 71.676
R1640 B.n516 B.n334 71.676
R1641 B.n523 B.n522 71.676
R1642 B.n524 B.n332 71.676
R1643 B.n531 B.n530 71.676
R1644 B.n534 B.n533 71.676
R1645 B.n463 B.n462 59.5399
R1646 B.n443 B.n354 59.5399
R1647 B.n108 B.n107 59.5399
R1648 B.n105 B.n104 59.5399
R1649 B.n539 B.n324 48.4618
R1650 B.n545 B.n324 48.4618
R1651 B.n545 B.n320 48.4618
R1652 B.n552 B.n320 48.4618
R1653 B.n552 B.n551 48.4618
R1654 B.n558 B.n313 48.4618
R1655 B.n564 B.n313 48.4618
R1656 B.n564 B.n309 48.4618
R1657 B.n570 B.n309 48.4618
R1658 B.n570 B.n305 48.4618
R1659 B.n577 B.n305 48.4618
R1660 B.n577 B.n576 48.4618
R1661 B.n583 B.n298 48.4618
R1662 B.n589 B.n298 48.4618
R1663 B.n589 B.n294 48.4618
R1664 B.n595 B.n294 48.4618
R1665 B.n601 B.n290 48.4618
R1666 B.n601 B.n285 48.4618
R1667 B.n607 B.n285 48.4618
R1668 B.n607 B.n286 48.4618
R1669 B.n613 B.n277 48.4618
R1670 B.n619 B.n277 48.4618
R1671 B.n619 B.n278 48.4618
R1672 B.n626 B.n270 48.4618
R1673 B.n632 B.n270 48.4618
R1674 B.n632 B.n4 48.4618
R1675 B.n745 B.n4 48.4618
R1676 B.n745 B.n744 48.4618
R1677 B.n744 B.n743 48.4618
R1678 B.n743 B.n8 48.4618
R1679 B.n737 B.n8 48.4618
R1680 B.n736 B.n735 48.4618
R1681 B.n735 B.n15 48.4618
R1682 B.n729 B.n15 48.4618
R1683 B.n728 B.n727 48.4618
R1684 B.n727 B.n22 48.4618
R1685 B.n721 B.n22 48.4618
R1686 B.n721 B.n720 48.4618
R1687 B.n719 B.n29 48.4618
R1688 B.n713 B.n29 48.4618
R1689 B.n713 B.n712 48.4618
R1690 B.n712 B.n711 48.4618
R1691 B.n705 B.n39 48.4618
R1692 B.n705 B.n704 48.4618
R1693 B.n704 B.n703 48.4618
R1694 B.n703 B.n43 48.4618
R1695 B.n697 B.n43 48.4618
R1696 B.n697 B.n696 48.4618
R1697 B.n696 B.n695 48.4618
R1698 B.n689 B.n53 48.4618
R1699 B.n689 B.n688 48.4618
R1700 B.n688 B.n687 48.4618
R1701 B.n687 B.n57 48.4618
R1702 B.n681 B.n57 48.4618
R1703 B.n278 B.t6 47.7491
R1704 B.t0 B.n736 47.7491
R1705 B.n613 B.t1 40.6225
R1706 B.n729 B.t2 40.6225
R1707 B.n683 B.n59 34.8103
R1708 B.n677 B.n676 34.8103
R1709 B.n537 B.n536 34.8103
R1710 B.n541 B.n326 34.8103
R1711 B.t7 B.n290 32.0705
R1712 B.n720 B.t4 32.0705
R1713 B.n462 B.n461 31.8066
R1714 B.n354 B.n353 31.8066
R1715 B.n107 B.n106 31.8066
R1716 B.n104 B.n103 31.8066
R1717 B.n558 B.t16 24.9438
R1718 B.n576 B.t5 24.9438
R1719 B.n39 B.t3 24.9438
R1720 B.n695 B.t9 24.9438
R1721 B.n551 B.t16 23.5185
R1722 B.n583 B.t5 23.5185
R1723 B.n711 B.t3 23.5185
R1724 B.n53 B.t9 23.5185
R1725 B B.n747 18.0485
R1726 B.n595 B.t7 16.3918
R1727 B.t4 B.n719 16.3918
R1728 B.n109 B.n59 10.6151
R1729 B.n112 B.n109 10.6151
R1730 B.n113 B.n112 10.6151
R1731 B.n116 B.n113 10.6151
R1732 B.n117 B.n116 10.6151
R1733 B.n120 B.n117 10.6151
R1734 B.n121 B.n120 10.6151
R1735 B.n124 B.n121 10.6151
R1736 B.n125 B.n124 10.6151
R1737 B.n128 B.n125 10.6151
R1738 B.n129 B.n128 10.6151
R1739 B.n132 B.n129 10.6151
R1740 B.n133 B.n132 10.6151
R1741 B.n136 B.n133 10.6151
R1742 B.n137 B.n136 10.6151
R1743 B.n140 B.n137 10.6151
R1744 B.n141 B.n140 10.6151
R1745 B.n144 B.n141 10.6151
R1746 B.n145 B.n144 10.6151
R1747 B.n148 B.n145 10.6151
R1748 B.n149 B.n148 10.6151
R1749 B.n152 B.n149 10.6151
R1750 B.n153 B.n152 10.6151
R1751 B.n156 B.n153 10.6151
R1752 B.n157 B.n156 10.6151
R1753 B.n160 B.n157 10.6151
R1754 B.n161 B.n160 10.6151
R1755 B.n164 B.n161 10.6151
R1756 B.n165 B.n164 10.6151
R1757 B.n168 B.n165 10.6151
R1758 B.n169 B.n168 10.6151
R1759 B.n172 B.n169 10.6151
R1760 B.n173 B.n172 10.6151
R1761 B.n176 B.n173 10.6151
R1762 B.n177 B.n176 10.6151
R1763 B.n181 B.n180 10.6151
R1764 B.n184 B.n181 10.6151
R1765 B.n185 B.n184 10.6151
R1766 B.n188 B.n185 10.6151
R1767 B.n189 B.n188 10.6151
R1768 B.n192 B.n189 10.6151
R1769 B.n193 B.n192 10.6151
R1770 B.n196 B.n193 10.6151
R1771 B.n197 B.n196 10.6151
R1772 B.n201 B.n200 10.6151
R1773 B.n204 B.n201 10.6151
R1774 B.n205 B.n204 10.6151
R1775 B.n208 B.n205 10.6151
R1776 B.n209 B.n208 10.6151
R1777 B.n212 B.n209 10.6151
R1778 B.n213 B.n212 10.6151
R1779 B.n216 B.n213 10.6151
R1780 B.n217 B.n216 10.6151
R1781 B.n220 B.n217 10.6151
R1782 B.n221 B.n220 10.6151
R1783 B.n224 B.n221 10.6151
R1784 B.n225 B.n224 10.6151
R1785 B.n228 B.n225 10.6151
R1786 B.n229 B.n228 10.6151
R1787 B.n232 B.n229 10.6151
R1788 B.n233 B.n232 10.6151
R1789 B.n236 B.n233 10.6151
R1790 B.n237 B.n236 10.6151
R1791 B.n240 B.n237 10.6151
R1792 B.n241 B.n240 10.6151
R1793 B.n244 B.n241 10.6151
R1794 B.n245 B.n244 10.6151
R1795 B.n248 B.n245 10.6151
R1796 B.n249 B.n248 10.6151
R1797 B.n252 B.n249 10.6151
R1798 B.n253 B.n252 10.6151
R1799 B.n256 B.n253 10.6151
R1800 B.n257 B.n256 10.6151
R1801 B.n260 B.n257 10.6151
R1802 B.n261 B.n260 10.6151
R1803 B.n264 B.n261 10.6151
R1804 B.n266 B.n264 10.6151
R1805 B.n267 B.n266 10.6151
R1806 B.n677 B.n267 10.6151
R1807 B.n537 B.n322 10.6151
R1808 B.n547 B.n322 10.6151
R1809 B.n548 B.n547 10.6151
R1810 B.n549 B.n548 10.6151
R1811 B.n549 B.n315 10.6151
R1812 B.n560 B.n315 10.6151
R1813 B.n561 B.n560 10.6151
R1814 B.n562 B.n561 10.6151
R1815 B.n562 B.n307 10.6151
R1816 B.n572 B.n307 10.6151
R1817 B.n573 B.n572 10.6151
R1818 B.n574 B.n573 10.6151
R1819 B.n574 B.n300 10.6151
R1820 B.n585 B.n300 10.6151
R1821 B.n586 B.n585 10.6151
R1822 B.n587 B.n586 10.6151
R1823 B.n587 B.n292 10.6151
R1824 B.n597 B.n292 10.6151
R1825 B.n598 B.n597 10.6151
R1826 B.n599 B.n598 10.6151
R1827 B.n599 B.n283 10.6151
R1828 B.n609 B.n283 10.6151
R1829 B.n610 B.n609 10.6151
R1830 B.n611 B.n610 10.6151
R1831 B.n611 B.n275 10.6151
R1832 B.n621 B.n275 10.6151
R1833 B.n622 B.n621 10.6151
R1834 B.n624 B.n622 10.6151
R1835 B.n624 B.n623 10.6151
R1836 B.n623 B.n268 10.6151
R1837 B.n635 B.n268 10.6151
R1838 B.n636 B.n635 10.6151
R1839 B.n637 B.n636 10.6151
R1840 B.n638 B.n637 10.6151
R1841 B.n640 B.n638 10.6151
R1842 B.n641 B.n640 10.6151
R1843 B.n642 B.n641 10.6151
R1844 B.n643 B.n642 10.6151
R1845 B.n645 B.n643 10.6151
R1846 B.n646 B.n645 10.6151
R1847 B.n647 B.n646 10.6151
R1848 B.n648 B.n647 10.6151
R1849 B.n650 B.n648 10.6151
R1850 B.n651 B.n650 10.6151
R1851 B.n652 B.n651 10.6151
R1852 B.n653 B.n652 10.6151
R1853 B.n655 B.n653 10.6151
R1854 B.n656 B.n655 10.6151
R1855 B.n657 B.n656 10.6151
R1856 B.n658 B.n657 10.6151
R1857 B.n660 B.n658 10.6151
R1858 B.n661 B.n660 10.6151
R1859 B.n662 B.n661 10.6151
R1860 B.n663 B.n662 10.6151
R1861 B.n665 B.n663 10.6151
R1862 B.n666 B.n665 10.6151
R1863 B.n667 B.n666 10.6151
R1864 B.n668 B.n667 10.6151
R1865 B.n670 B.n668 10.6151
R1866 B.n671 B.n670 10.6151
R1867 B.n672 B.n671 10.6151
R1868 B.n673 B.n672 10.6151
R1869 B.n675 B.n673 10.6151
R1870 B.n676 B.n675 10.6151
R1871 B.n372 B.n326 10.6151
R1872 B.n372 B.n371 10.6151
R1873 B.n378 B.n371 10.6151
R1874 B.n379 B.n378 10.6151
R1875 B.n380 B.n379 10.6151
R1876 B.n380 B.n369 10.6151
R1877 B.n386 B.n369 10.6151
R1878 B.n387 B.n386 10.6151
R1879 B.n388 B.n387 10.6151
R1880 B.n388 B.n367 10.6151
R1881 B.n394 B.n367 10.6151
R1882 B.n395 B.n394 10.6151
R1883 B.n396 B.n395 10.6151
R1884 B.n396 B.n365 10.6151
R1885 B.n402 B.n365 10.6151
R1886 B.n403 B.n402 10.6151
R1887 B.n404 B.n403 10.6151
R1888 B.n404 B.n363 10.6151
R1889 B.n410 B.n363 10.6151
R1890 B.n411 B.n410 10.6151
R1891 B.n412 B.n411 10.6151
R1892 B.n412 B.n361 10.6151
R1893 B.n418 B.n361 10.6151
R1894 B.n419 B.n418 10.6151
R1895 B.n420 B.n419 10.6151
R1896 B.n420 B.n359 10.6151
R1897 B.n426 B.n359 10.6151
R1898 B.n427 B.n426 10.6151
R1899 B.n428 B.n427 10.6151
R1900 B.n428 B.n357 10.6151
R1901 B.n434 B.n357 10.6151
R1902 B.n435 B.n434 10.6151
R1903 B.n436 B.n435 10.6151
R1904 B.n436 B.n355 10.6151
R1905 B.n442 B.n355 10.6151
R1906 B.n445 B.n444 10.6151
R1907 B.n445 B.n351 10.6151
R1908 B.n451 B.n351 10.6151
R1909 B.n452 B.n451 10.6151
R1910 B.n453 B.n452 10.6151
R1911 B.n453 B.n349 10.6151
R1912 B.n459 B.n349 10.6151
R1913 B.n460 B.n459 10.6151
R1914 B.n464 B.n460 10.6151
R1915 B.n470 B.n347 10.6151
R1916 B.n471 B.n470 10.6151
R1917 B.n472 B.n471 10.6151
R1918 B.n472 B.n345 10.6151
R1919 B.n478 B.n345 10.6151
R1920 B.n479 B.n478 10.6151
R1921 B.n480 B.n479 10.6151
R1922 B.n480 B.n343 10.6151
R1923 B.n486 B.n343 10.6151
R1924 B.n487 B.n486 10.6151
R1925 B.n488 B.n487 10.6151
R1926 B.n488 B.n341 10.6151
R1927 B.n494 B.n341 10.6151
R1928 B.n495 B.n494 10.6151
R1929 B.n496 B.n495 10.6151
R1930 B.n496 B.n339 10.6151
R1931 B.n502 B.n339 10.6151
R1932 B.n503 B.n502 10.6151
R1933 B.n504 B.n503 10.6151
R1934 B.n504 B.n337 10.6151
R1935 B.n510 B.n337 10.6151
R1936 B.n511 B.n510 10.6151
R1937 B.n512 B.n511 10.6151
R1938 B.n512 B.n335 10.6151
R1939 B.n518 B.n335 10.6151
R1940 B.n519 B.n518 10.6151
R1941 B.n520 B.n519 10.6151
R1942 B.n520 B.n333 10.6151
R1943 B.n526 B.n333 10.6151
R1944 B.n527 B.n526 10.6151
R1945 B.n528 B.n527 10.6151
R1946 B.n528 B.n331 10.6151
R1947 B.n331 B.n330 10.6151
R1948 B.n535 B.n330 10.6151
R1949 B.n536 B.n535 10.6151
R1950 B.n542 B.n541 10.6151
R1951 B.n543 B.n542 10.6151
R1952 B.n543 B.n318 10.6151
R1953 B.n554 B.n318 10.6151
R1954 B.n555 B.n554 10.6151
R1955 B.n556 B.n555 10.6151
R1956 B.n556 B.n311 10.6151
R1957 B.n566 B.n311 10.6151
R1958 B.n567 B.n566 10.6151
R1959 B.n568 B.n567 10.6151
R1960 B.n568 B.n303 10.6151
R1961 B.n579 B.n303 10.6151
R1962 B.n580 B.n579 10.6151
R1963 B.n581 B.n580 10.6151
R1964 B.n581 B.n296 10.6151
R1965 B.n591 B.n296 10.6151
R1966 B.n592 B.n591 10.6151
R1967 B.n593 B.n592 10.6151
R1968 B.n593 B.n288 10.6151
R1969 B.n603 B.n288 10.6151
R1970 B.n604 B.n603 10.6151
R1971 B.n605 B.n604 10.6151
R1972 B.n605 B.n280 10.6151
R1973 B.n615 B.n280 10.6151
R1974 B.n616 B.n615 10.6151
R1975 B.n617 B.n616 10.6151
R1976 B.n617 B.n272 10.6151
R1977 B.n628 B.n272 10.6151
R1978 B.n629 B.n628 10.6151
R1979 B.n630 B.n629 10.6151
R1980 B.n630 B.n0 10.6151
R1981 B.n741 B.n1 10.6151
R1982 B.n741 B.n740 10.6151
R1983 B.n740 B.n739 10.6151
R1984 B.n739 B.n10 10.6151
R1985 B.n733 B.n10 10.6151
R1986 B.n733 B.n732 10.6151
R1987 B.n732 B.n731 10.6151
R1988 B.n731 B.n17 10.6151
R1989 B.n725 B.n17 10.6151
R1990 B.n725 B.n724 10.6151
R1991 B.n724 B.n723 10.6151
R1992 B.n723 B.n24 10.6151
R1993 B.n717 B.n24 10.6151
R1994 B.n717 B.n716 10.6151
R1995 B.n716 B.n715 10.6151
R1996 B.n715 B.n31 10.6151
R1997 B.n709 B.n31 10.6151
R1998 B.n709 B.n708 10.6151
R1999 B.n708 B.n707 10.6151
R2000 B.n707 B.n37 10.6151
R2001 B.n701 B.n37 10.6151
R2002 B.n701 B.n700 10.6151
R2003 B.n700 B.n699 10.6151
R2004 B.n699 B.n45 10.6151
R2005 B.n693 B.n45 10.6151
R2006 B.n693 B.n692 10.6151
R2007 B.n692 B.n691 10.6151
R2008 B.n691 B.n51 10.6151
R2009 B.n685 B.n51 10.6151
R2010 B.n685 B.n684 10.6151
R2011 B.n684 B.n683 10.6151
R2012 B.n177 B.n108 9.36635
R2013 B.n200 B.n105 9.36635
R2014 B.n443 B.n442 9.36635
R2015 B.n463 B.n347 9.36635
R2016 B.n286 B.t1 7.83983
R2017 B.t2 B.n728 7.83983
R2018 B.n747 B.n0 2.81026
R2019 B.n747 B.n1 2.81026
R2020 B.n180 B.n108 1.24928
R2021 B.n197 B.n105 1.24928
R2022 B.n444 B.n443 1.24928
R2023 B.n464 B.n463 1.24928
R2024 B.n626 B.t6 0.713166
R2025 B.n737 B.t0 0.713166
R2026 VP.n11 VP.t7 214.504
R2027 VP.n5 VP.t3 186.913
R2028 VP.n29 VP.t0 186.913
R2029 VP.n36 VP.t1 186.913
R2030 VP.n43 VP.t2 186.913
R2031 VP.n23 VP.t4 186.913
R2032 VP.n16 VP.t5 186.913
R2033 VP.n10 VP.t6 186.913
R2034 VP.n25 VP.n5 175.564
R2035 VP.n44 VP.n43 175.564
R2036 VP.n24 VP.n23 175.564
R2037 VP.n12 VP.n9 161.3
R2038 VP.n14 VP.n13 161.3
R2039 VP.n15 VP.n8 161.3
R2040 VP.n18 VP.n17 161.3
R2041 VP.n19 VP.n7 161.3
R2042 VP.n21 VP.n20 161.3
R2043 VP.n22 VP.n6 161.3
R2044 VP.n42 VP.n0 161.3
R2045 VP.n41 VP.n40 161.3
R2046 VP.n39 VP.n1 161.3
R2047 VP.n38 VP.n37 161.3
R2048 VP.n35 VP.n2 161.3
R2049 VP.n34 VP.n33 161.3
R2050 VP.n32 VP.n3 161.3
R2051 VP.n31 VP.n30 161.3
R2052 VP.n28 VP.n4 161.3
R2053 VP.n27 VP.n26 161.3
R2054 VP.n11 VP.n10 62.2212
R2055 VP.n35 VP.n34 56.5617
R2056 VP.n15 VP.n14 56.5617
R2057 VP.n30 VP.n28 51.2335
R2058 VP.n41 VP.n1 51.2335
R2059 VP.n21 VP.n7 51.2335
R2060 VP.n25 VP.n24 43.349
R2061 VP.n28 VP.n27 29.9206
R2062 VP.n42 VP.n41 29.9206
R2063 VP.n22 VP.n21 29.9206
R2064 VP.n12 VP.n11 27.6221
R2065 VP.n34 VP.n3 24.5923
R2066 VP.n37 VP.n35 24.5923
R2067 VP.n17 VP.n15 24.5923
R2068 VP.n14 VP.n9 24.5923
R2069 VP.n30 VP.n29 21.1495
R2070 VP.n36 VP.n1 21.1495
R2071 VP.n16 VP.n7 21.1495
R2072 VP.n27 VP.n5 10.3291
R2073 VP.n43 VP.n42 10.3291
R2074 VP.n23 VP.n22 10.3291
R2075 VP.n29 VP.n3 3.44336
R2076 VP.n37 VP.n36 3.44336
R2077 VP.n17 VP.n16 3.44336
R2078 VP.n10 VP.n9 3.44336
R2079 VP.n13 VP.n12 0.189894
R2080 VP.n13 VP.n8 0.189894
R2081 VP.n18 VP.n8 0.189894
R2082 VP.n19 VP.n18 0.189894
R2083 VP.n20 VP.n19 0.189894
R2084 VP.n20 VP.n6 0.189894
R2085 VP.n24 VP.n6 0.189894
R2086 VP.n26 VP.n25 0.189894
R2087 VP.n26 VP.n4 0.189894
R2088 VP.n31 VP.n4 0.189894
R2089 VP.n32 VP.n31 0.189894
R2090 VP.n33 VP.n32 0.189894
R2091 VP.n33 VP.n2 0.189894
R2092 VP.n38 VP.n2 0.189894
R2093 VP.n39 VP.n38 0.189894
R2094 VP.n40 VP.n39 0.189894
R2095 VP.n40 VP.n0 0.189894
R2096 VP.n44 VP.n0 0.189894
R2097 VP VP.n44 0.0516364
R2098 VDD1 VDD1.n0 67.2842
R2099 VDD1.n3 VDD1.n2 67.1705
R2100 VDD1.n3 VDD1.n1 67.1705
R2101 VDD1.n5 VDD1.n4 66.5189
R2102 VDD1.n5 VDD1.n3 39.419
R2103 VDD1.n4 VDD1.t2 1.94932
R2104 VDD1.n4 VDD1.t3 1.94932
R2105 VDD1.n0 VDD1.t0 1.94932
R2106 VDD1.n0 VDD1.t1 1.94932
R2107 VDD1.n2 VDD1.t6 1.94932
R2108 VDD1.n2 VDD1.t5 1.94932
R2109 VDD1.n1 VDD1.t4 1.94932
R2110 VDD1.n1 VDD1.t7 1.94932
R2111 VDD1 VDD1.n5 0.649207
C0 VN VDD1 0.149579f
C1 VN VDD2 6.18474f
C2 VN VTAIL 6.23578f
C3 VP VDD1 6.417f
C4 VP VDD2 0.382584f
C5 VTAIL VP 6.24988f
C6 VN VP 5.74269f
C7 VDD1 VDD2 1.13131f
C8 VTAIL VDD1 7.83704f
C9 VTAIL VDD2 7.882811f
C10 VDD2 B 3.931486f
C11 VDD1 B 4.227607f
C12 VTAIL B 8.430452f
C13 VN B 10.500951f
C14 VP B 8.895383f
C15 VDD1.t0 B 0.2029f
C16 VDD1.t1 B 0.2029f
C17 VDD1.n0 B 1.79611f
C18 VDD1.t4 B 0.2029f
C19 VDD1.t7 B 0.2029f
C20 VDD1.n1 B 1.79537f
C21 VDD1.t6 B 0.2029f
C22 VDD1.t5 B 0.2029f
C23 VDD1.n2 B 1.79537f
C24 VDD1.n3 B 2.48612f
C25 VDD1.t2 B 0.2029f
C26 VDD1.t3 B 0.2029f
C27 VDD1.n4 B 1.79165f
C28 VDD1.n5 B 2.41063f
C29 VP.n0 B 0.033918f
C30 VP.t2 B 1.22362f
C31 VP.n1 B 0.056936f
C32 VP.n2 B 0.033918f
C33 VP.n3 B 0.036194f
C34 VP.n4 B 0.033918f
C35 VP.t3 B 1.22362f
C36 VP.n5 B 0.511688f
C37 VP.n6 B 0.033918f
C38 VP.t4 B 1.22362f
C39 VP.n7 B 0.056936f
C40 VP.n8 B 0.033918f
C41 VP.n9 B 0.036194f
C42 VP.t7 B 1.29552f
C43 VP.t6 B 1.22362f
C44 VP.n10 B 0.497762f
C45 VP.n11 B 0.535597f
C46 VP.n12 B 0.177945f
C47 VP.n13 B 0.033918f
C48 VP.n14 B 0.049305f
C49 VP.n15 B 0.049305f
C50 VP.t5 B 1.22362f
C51 VP.n16 B 0.452759f
C52 VP.n17 B 0.036194f
C53 VP.n18 B 0.033918f
C54 VP.n19 B 0.033918f
C55 VP.n20 B 0.033918f
C56 VP.n21 B 0.033014f
C57 VP.n22 B 0.049201f
C58 VP.n23 B 0.511688f
C59 VP.n24 B 1.48012f
C60 VP.n25 B 1.50832f
C61 VP.n26 B 0.033918f
C62 VP.n27 B 0.049201f
C63 VP.n28 B 0.033014f
C64 VP.t0 B 1.22362f
C65 VP.n29 B 0.452759f
C66 VP.n30 B 0.056936f
C67 VP.n31 B 0.033918f
C68 VP.n32 B 0.033918f
C69 VP.n33 B 0.033918f
C70 VP.n34 B 0.049305f
C71 VP.n35 B 0.049305f
C72 VP.t1 B 1.22362f
C73 VP.n36 B 0.452759f
C74 VP.n37 B 0.036194f
C75 VP.n38 B 0.033918f
C76 VP.n39 B 0.033918f
C77 VP.n40 B 0.033918f
C78 VP.n41 B 0.033014f
C79 VP.n42 B 0.049201f
C80 VP.n43 B 0.511688f
C81 VP.n44 B 0.031496f
C82 VDD2.t6 B 0.202804f
C83 VDD2.t3 B 0.202804f
C84 VDD2.n0 B 1.79452f
C85 VDD2.t5 B 0.202804f
C86 VDD2.t7 B 0.202804f
C87 VDD2.n1 B 1.79452f
C88 VDD2.n2 B 2.43143f
C89 VDD2.t0 B 0.202804f
C90 VDD2.t1 B 0.202804f
C91 VDD2.n3 B 1.79082f
C92 VDD2.n4 B 2.37918f
C93 VDD2.t4 B 0.202804f
C94 VDD2.t2 B 0.202804f
C95 VDD2.n5 B 1.79449f
C96 VTAIL.t14 B 0.157245f
C97 VTAIL.t11 B 0.157245f
C98 VTAIL.n0 B 1.33704f
C99 VTAIL.n1 B 0.27528f
C100 VTAIL.n2 B 0.028586f
C101 VTAIL.n3 B 0.019585f
C102 VTAIL.n4 B 0.010524f
C103 VTAIL.n5 B 0.024875f
C104 VTAIL.n6 B 0.011143f
C105 VTAIL.n7 B 0.019585f
C106 VTAIL.n8 B 0.010834f
C107 VTAIL.n9 B 0.024875f
C108 VTAIL.n10 B 0.011143f
C109 VTAIL.n11 B 0.019585f
C110 VTAIL.n12 B 0.010524f
C111 VTAIL.n13 B 0.024875f
C112 VTAIL.n14 B 0.011143f
C113 VTAIL.n15 B 0.019585f
C114 VTAIL.n16 B 0.010524f
C115 VTAIL.n17 B 0.018657f
C116 VTAIL.n18 B 0.017585f
C117 VTAIL.t12 B 0.041821f
C118 VTAIL.n19 B 0.127376f
C119 VTAIL.n20 B 0.827749f
C120 VTAIL.n21 B 0.010524f
C121 VTAIL.n22 B 0.011143f
C122 VTAIL.n23 B 0.024875f
C123 VTAIL.n24 B 0.024875f
C124 VTAIL.n25 B 0.011143f
C125 VTAIL.n26 B 0.010524f
C126 VTAIL.n27 B 0.019585f
C127 VTAIL.n28 B 0.019585f
C128 VTAIL.n29 B 0.010524f
C129 VTAIL.n30 B 0.011143f
C130 VTAIL.n31 B 0.024875f
C131 VTAIL.n32 B 0.024875f
C132 VTAIL.n33 B 0.011143f
C133 VTAIL.n34 B 0.010524f
C134 VTAIL.n35 B 0.019585f
C135 VTAIL.n36 B 0.019585f
C136 VTAIL.n37 B 0.010524f
C137 VTAIL.n38 B 0.010524f
C138 VTAIL.n39 B 0.011143f
C139 VTAIL.n40 B 0.024875f
C140 VTAIL.n41 B 0.024875f
C141 VTAIL.n42 B 0.024875f
C142 VTAIL.n43 B 0.010834f
C143 VTAIL.n44 B 0.010524f
C144 VTAIL.n45 B 0.019585f
C145 VTAIL.n46 B 0.019585f
C146 VTAIL.n47 B 0.010524f
C147 VTAIL.n48 B 0.011143f
C148 VTAIL.n49 B 0.024875f
C149 VTAIL.n50 B 0.055721f
C150 VTAIL.n51 B 0.011143f
C151 VTAIL.n52 B 0.010524f
C152 VTAIL.n53 B 0.050621f
C153 VTAIL.n54 B 0.031526f
C154 VTAIL.n55 B 0.138627f
C155 VTAIL.n56 B 0.028586f
C156 VTAIL.n57 B 0.019585f
C157 VTAIL.n58 B 0.010524f
C158 VTAIL.n59 B 0.024875f
C159 VTAIL.n60 B 0.011143f
C160 VTAIL.n61 B 0.019585f
C161 VTAIL.n62 B 0.010834f
C162 VTAIL.n63 B 0.024875f
C163 VTAIL.n64 B 0.011143f
C164 VTAIL.n65 B 0.019585f
C165 VTAIL.n66 B 0.010524f
C166 VTAIL.n67 B 0.024875f
C167 VTAIL.n68 B 0.011143f
C168 VTAIL.n69 B 0.019585f
C169 VTAIL.n70 B 0.010524f
C170 VTAIL.n71 B 0.018657f
C171 VTAIL.n72 B 0.017585f
C172 VTAIL.t6 B 0.041821f
C173 VTAIL.n73 B 0.127376f
C174 VTAIL.n74 B 0.827749f
C175 VTAIL.n75 B 0.010524f
C176 VTAIL.n76 B 0.011143f
C177 VTAIL.n77 B 0.024875f
C178 VTAIL.n78 B 0.024875f
C179 VTAIL.n79 B 0.011143f
C180 VTAIL.n80 B 0.010524f
C181 VTAIL.n81 B 0.019585f
C182 VTAIL.n82 B 0.019585f
C183 VTAIL.n83 B 0.010524f
C184 VTAIL.n84 B 0.011143f
C185 VTAIL.n85 B 0.024875f
C186 VTAIL.n86 B 0.024875f
C187 VTAIL.n87 B 0.011143f
C188 VTAIL.n88 B 0.010524f
C189 VTAIL.n89 B 0.019585f
C190 VTAIL.n90 B 0.019585f
C191 VTAIL.n91 B 0.010524f
C192 VTAIL.n92 B 0.010524f
C193 VTAIL.n93 B 0.011143f
C194 VTAIL.n94 B 0.024875f
C195 VTAIL.n95 B 0.024875f
C196 VTAIL.n96 B 0.024875f
C197 VTAIL.n97 B 0.010834f
C198 VTAIL.n98 B 0.010524f
C199 VTAIL.n99 B 0.019585f
C200 VTAIL.n100 B 0.019585f
C201 VTAIL.n101 B 0.010524f
C202 VTAIL.n102 B 0.011143f
C203 VTAIL.n103 B 0.024875f
C204 VTAIL.n104 B 0.055721f
C205 VTAIL.n105 B 0.011143f
C206 VTAIL.n106 B 0.010524f
C207 VTAIL.n107 B 0.050621f
C208 VTAIL.n108 B 0.031526f
C209 VTAIL.n109 B 0.138627f
C210 VTAIL.t7 B 0.157245f
C211 VTAIL.t1 B 0.157245f
C212 VTAIL.n110 B 1.33704f
C213 VTAIL.n111 B 0.36083f
C214 VTAIL.n112 B 0.028586f
C215 VTAIL.n113 B 0.019585f
C216 VTAIL.n114 B 0.010524f
C217 VTAIL.n115 B 0.024875f
C218 VTAIL.n116 B 0.011143f
C219 VTAIL.n117 B 0.019585f
C220 VTAIL.n118 B 0.010834f
C221 VTAIL.n119 B 0.024875f
C222 VTAIL.n120 B 0.011143f
C223 VTAIL.n121 B 0.019585f
C224 VTAIL.n122 B 0.010524f
C225 VTAIL.n123 B 0.024875f
C226 VTAIL.n124 B 0.011143f
C227 VTAIL.n125 B 0.019585f
C228 VTAIL.n126 B 0.010524f
C229 VTAIL.n127 B 0.018657f
C230 VTAIL.n128 B 0.017585f
C231 VTAIL.t5 B 0.041821f
C232 VTAIL.n129 B 0.127376f
C233 VTAIL.n130 B 0.827749f
C234 VTAIL.n131 B 0.010524f
C235 VTAIL.n132 B 0.011143f
C236 VTAIL.n133 B 0.024875f
C237 VTAIL.n134 B 0.024875f
C238 VTAIL.n135 B 0.011143f
C239 VTAIL.n136 B 0.010524f
C240 VTAIL.n137 B 0.019585f
C241 VTAIL.n138 B 0.019585f
C242 VTAIL.n139 B 0.010524f
C243 VTAIL.n140 B 0.011143f
C244 VTAIL.n141 B 0.024875f
C245 VTAIL.n142 B 0.024875f
C246 VTAIL.n143 B 0.011143f
C247 VTAIL.n144 B 0.010524f
C248 VTAIL.n145 B 0.019585f
C249 VTAIL.n146 B 0.019585f
C250 VTAIL.n147 B 0.010524f
C251 VTAIL.n148 B 0.010524f
C252 VTAIL.n149 B 0.011143f
C253 VTAIL.n150 B 0.024875f
C254 VTAIL.n151 B 0.024875f
C255 VTAIL.n152 B 0.024875f
C256 VTAIL.n153 B 0.010834f
C257 VTAIL.n154 B 0.010524f
C258 VTAIL.n155 B 0.019585f
C259 VTAIL.n156 B 0.019585f
C260 VTAIL.n157 B 0.010524f
C261 VTAIL.n158 B 0.011143f
C262 VTAIL.n159 B 0.024875f
C263 VTAIL.n160 B 0.055721f
C264 VTAIL.n161 B 0.011143f
C265 VTAIL.n162 B 0.010524f
C266 VTAIL.n163 B 0.050621f
C267 VTAIL.n164 B 0.031526f
C268 VTAIL.n165 B 1.01698f
C269 VTAIL.n166 B 0.028586f
C270 VTAIL.n167 B 0.019585f
C271 VTAIL.n168 B 0.010524f
C272 VTAIL.n169 B 0.024875f
C273 VTAIL.n170 B 0.011143f
C274 VTAIL.n171 B 0.019585f
C275 VTAIL.n172 B 0.010834f
C276 VTAIL.n173 B 0.024875f
C277 VTAIL.n174 B 0.010524f
C278 VTAIL.n175 B 0.011143f
C279 VTAIL.n176 B 0.019585f
C280 VTAIL.n177 B 0.010524f
C281 VTAIL.n178 B 0.024875f
C282 VTAIL.n179 B 0.011143f
C283 VTAIL.n180 B 0.019585f
C284 VTAIL.n181 B 0.010524f
C285 VTAIL.n182 B 0.018657f
C286 VTAIL.n183 B 0.017585f
C287 VTAIL.t15 B 0.041821f
C288 VTAIL.n184 B 0.127376f
C289 VTAIL.n185 B 0.827749f
C290 VTAIL.n186 B 0.010524f
C291 VTAIL.n187 B 0.011143f
C292 VTAIL.n188 B 0.024875f
C293 VTAIL.n189 B 0.024875f
C294 VTAIL.n190 B 0.011143f
C295 VTAIL.n191 B 0.010524f
C296 VTAIL.n192 B 0.019585f
C297 VTAIL.n193 B 0.019585f
C298 VTAIL.n194 B 0.010524f
C299 VTAIL.n195 B 0.011143f
C300 VTAIL.n196 B 0.024875f
C301 VTAIL.n197 B 0.024875f
C302 VTAIL.n198 B 0.011143f
C303 VTAIL.n199 B 0.010524f
C304 VTAIL.n200 B 0.019585f
C305 VTAIL.n201 B 0.019585f
C306 VTAIL.n202 B 0.010524f
C307 VTAIL.n203 B 0.011143f
C308 VTAIL.n204 B 0.024875f
C309 VTAIL.n205 B 0.024875f
C310 VTAIL.n206 B 0.024875f
C311 VTAIL.n207 B 0.010834f
C312 VTAIL.n208 B 0.010524f
C313 VTAIL.n209 B 0.019585f
C314 VTAIL.n210 B 0.019585f
C315 VTAIL.n211 B 0.010524f
C316 VTAIL.n212 B 0.011143f
C317 VTAIL.n213 B 0.024875f
C318 VTAIL.n214 B 0.055721f
C319 VTAIL.n215 B 0.011143f
C320 VTAIL.n216 B 0.010524f
C321 VTAIL.n217 B 0.050621f
C322 VTAIL.n218 B 0.031526f
C323 VTAIL.n219 B 1.01698f
C324 VTAIL.t10 B 0.157245f
C325 VTAIL.t8 B 0.157245f
C326 VTAIL.n220 B 1.33704f
C327 VTAIL.n221 B 0.360822f
C328 VTAIL.n222 B 0.028586f
C329 VTAIL.n223 B 0.019585f
C330 VTAIL.n224 B 0.010524f
C331 VTAIL.n225 B 0.024875f
C332 VTAIL.n226 B 0.011143f
C333 VTAIL.n227 B 0.019585f
C334 VTAIL.n228 B 0.010834f
C335 VTAIL.n229 B 0.024875f
C336 VTAIL.n230 B 0.010524f
C337 VTAIL.n231 B 0.011143f
C338 VTAIL.n232 B 0.019585f
C339 VTAIL.n233 B 0.010524f
C340 VTAIL.n234 B 0.024875f
C341 VTAIL.n235 B 0.011143f
C342 VTAIL.n236 B 0.019585f
C343 VTAIL.n237 B 0.010524f
C344 VTAIL.n238 B 0.018657f
C345 VTAIL.n239 B 0.017585f
C346 VTAIL.t13 B 0.041821f
C347 VTAIL.n240 B 0.127376f
C348 VTAIL.n241 B 0.827749f
C349 VTAIL.n242 B 0.010524f
C350 VTAIL.n243 B 0.011143f
C351 VTAIL.n244 B 0.024875f
C352 VTAIL.n245 B 0.024875f
C353 VTAIL.n246 B 0.011143f
C354 VTAIL.n247 B 0.010524f
C355 VTAIL.n248 B 0.019585f
C356 VTAIL.n249 B 0.019585f
C357 VTAIL.n250 B 0.010524f
C358 VTAIL.n251 B 0.011143f
C359 VTAIL.n252 B 0.024875f
C360 VTAIL.n253 B 0.024875f
C361 VTAIL.n254 B 0.011143f
C362 VTAIL.n255 B 0.010524f
C363 VTAIL.n256 B 0.019585f
C364 VTAIL.n257 B 0.019585f
C365 VTAIL.n258 B 0.010524f
C366 VTAIL.n259 B 0.011143f
C367 VTAIL.n260 B 0.024875f
C368 VTAIL.n261 B 0.024875f
C369 VTAIL.n262 B 0.024875f
C370 VTAIL.n263 B 0.010834f
C371 VTAIL.n264 B 0.010524f
C372 VTAIL.n265 B 0.019585f
C373 VTAIL.n266 B 0.019585f
C374 VTAIL.n267 B 0.010524f
C375 VTAIL.n268 B 0.011143f
C376 VTAIL.n269 B 0.024875f
C377 VTAIL.n270 B 0.055721f
C378 VTAIL.n271 B 0.011143f
C379 VTAIL.n272 B 0.010524f
C380 VTAIL.n273 B 0.050621f
C381 VTAIL.n274 B 0.031526f
C382 VTAIL.n275 B 0.138627f
C383 VTAIL.n276 B 0.028586f
C384 VTAIL.n277 B 0.019585f
C385 VTAIL.n278 B 0.010524f
C386 VTAIL.n279 B 0.024875f
C387 VTAIL.n280 B 0.011143f
C388 VTAIL.n281 B 0.019585f
C389 VTAIL.n282 B 0.010834f
C390 VTAIL.n283 B 0.024875f
C391 VTAIL.n284 B 0.010524f
C392 VTAIL.n285 B 0.011143f
C393 VTAIL.n286 B 0.019585f
C394 VTAIL.n287 B 0.010524f
C395 VTAIL.n288 B 0.024875f
C396 VTAIL.n289 B 0.011143f
C397 VTAIL.n290 B 0.019585f
C398 VTAIL.n291 B 0.010524f
C399 VTAIL.n292 B 0.018657f
C400 VTAIL.n293 B 0.017585f
C401 VTAIL.t0 B 0.041821f
C402 VTAIL.n294 B 0.127376f
C403 VTAIL.n295 B 0.827749f
C404 VTAIL.n296 B 0.010524f
C405 VTAIL.n297 B 0.011143f
C406 VTAIL.n298 B 0.024875f
C407 VTAIL.n299 B 0.024875f
C408 VTAIL.n300 B 0.011143f
C409 VTAIL.n301 B 0.010524f
C410 VTAIL.n302 B 0.019585f
C411 VTAIL.n303 B 0.019585f
C412 VTAIL.n304 B 0.010524f
C413 VTAIL.n305 B 0.011143f
C414 VTAIL.n306 B 0.024875f
C415 VTAIL.n307 B 0.024875f
C416 VTAIL.n308 B 0.011143f
C417 VTAIL.n309 B 0.010524f
C418 VTAIL.n310 B 0.019585f
C419 VTAIL.n311 B 0.019585f
C420 VTAIL.n312 B 0.010524f
C421 VTAIL.n313 B 0.011143f
C422 VTAIL.n314 B 0.024875f
C423 VTAIL.n315 B 0.024875f
C424 VTAIL.n316 B 0.024875f
C425 VTAIL.n317 B 0.010834f
C426 VTAIL.n318 B 0.010524f
C427 VTAIL.n319 B 0.019585f
C428 VTAIL.n320 B 0.019585f
C429 VTAIL.n321 B 0.010524f
C430 VTAIL.n322 B 0.011143f
C431 VTAIL.n323 B 0.024875f
C432 VTAIL.n324 B 0.055721f
C433 VTAIL.n325 B 0.011143f
C434 VTAIL.n326 B 0.010524f
C435 VTAIL.n327 B 0.050621f
C436 VTAIL.n328 B 0.031526f
C437 VTAIL.n329 B 0.138627f
C438 VTAIL.t2 B 0.157245f
C439 VTAIL.t4 B 0.157245f
C440 VTAIL.n330 B 1.33704f
C441 VTAIL.n331 B 0.360822f
C442 VTAIL.n332 B 0.028586f
C443 VTAIL.n333 B 0.019585f
C444 VTAIL.n334 B 0.010524f
C445 VTAIL.n335 B 0.024875f
C446 VTAIL.n336 B 0.011143f
C447 VTAIL.n337 B 0.019585f
C448 VTAIL.n338 B 0.010834f
C449 VTAIL.n339 B 0.024875f
C450 VTAIL.n340 B 0.010524f
C451 VTAIL.n341 B 0.011143f
C452 VTAIL.n342 B 0.019585f
C453 VTAIL.n343 B 0.010524f
C454 VTAIL.n344 B 0.024875f
C455 VTAIL.n345 B 0.011143f
C456 VTAIL.n346 B 0.019585f
C457 VTAIL.n347 B 0.010524f
C458 VTAIL.n348 B 0.018657f
C459 VTAIL.n349 B 0.017585f
C460 VTAIL.t3 B 0.041821f
C461 VTAIL.n350 B 0.127376f
C462 VTAIL.n351 B 0.827749f
C463 VTAIL.n352 B 0.010524f
C464 VTAIL.n353 B 0.011143f
C465 VTAIL.n354 B 0.024875f
C466 VTAIL.n355 B 0.024875f
C467 VTAIL.n356 B 0.011143f
C468 VTAIL.n357 B 0.010524f
C469 VTAIL.n358 B 0.019585f
C470 VTAIL.n359 B 0.019585f
C471 VTAIL.n360 B 0.010524f
C472 VTAIL.n361 B 0.011143f
C473 VTAIL.n362 B 0.024875f
C474 VTAIL.n363 B 0.024875f
C475 VTAIL.n364 B 0.011143f
C476 VTAIL.n365 B 0.010524f
C477 VTAIL.n366 B 0.019585f
C478 VTAIL.n367 B 0.019585f
C479 VTAIL.n368 B 0.010524f
C480 VTAIL.n369 B 0.011143f
C481 VTAIL.n370 B 0.024875f
C482 VTAIL.n371 B 0.024875f
C483 VTAIL.n372 B 0.024875f
C484 VTAIL.n373 B 0.010834f
C485 VTAIL.n374 B 0.010524f
C486 VTAIL.n375 B 0.019585f
C487 VTAIL.n376 B 0.019585f
C488 VTAIL.n377 B 0.010524f
C489 VTAIL.n378 B 0.011143f
C490 VTAIL.n379 B 0.024875f
C491 VTAIL.n380 B 0.055721f
C492 VTAIL.n381 B 0.011143f
C493 VTAIL.n382 B 0.010524f
C494 VTAIL.n383 B 0.050621f
C495 VTAIL.n384 B 0.031526f
C496 VTAIL.n385 B 1.01698f
C497 VTAIL.n386 B 0.028586f
C498 VTAIL.n387 B 0.019585f
C499 VTAIL.n388 B 0.010524f
C500 VTAIL.n389 B 0.024875f
C501 VTAIL.n390 B 0.011143f
C502 VTAIL.n391 B 0.019585f
C503 VTAIL.n392 B 0.010834f
C504 VTAIL.n393 B 0.024875f
C505 VTAIL.n394 B 0.011143f
C506 VTAIL.n395 B 0.019585f
C507 VTAIL.n396 B 0.010524f
C508 VTAIL.n397 B 0.024875f
C509 VTAIL.n398 B 0.011143f
C510 VTAIL.n399 B 0.019585f
C511 VTAIL.n400 B 0.010524f
C512 VTAIL.n401 B 0.018657f
C513 VTAIL.n402 B 0.017585f
C514 VTAIL.t9 B 0.041821f
C515 VTAIL.n403 B 0.127376f
C516 VTAIL.n404 B 0.827749f
C517 VTAIL.n405 B 0.010524f
C518 VTAIL.n406 B 0.011143f
C519 VTAIL.n407 B 0.024875f
C520 VTAIL.n408 B 0.024875f
C521 VTAIL.n409 B 0.011143f
C522 VTAIL.n410 B 0.010524f
C523 VTAIL.n411 B 0.019585f
C524 VTAIL.n412 B 0.019585f
C525 VTAIL.n413 B 0.010524f
C526 VTAIL.n414 B 0.011143f
C527 VTAIL.n415 B 0.024875f
C528 VTAIL.n416 B 0.024875f
C529 VTAIL.n417 B 0.011143f
C530 VTAIL.n418 B 0.010524f
C531 VTAIL.n419 B 0.019585f
C532 VTAIL.n420 B 0.019585f
C533 VTAIL.n421 B 0.010524f
C534 VTAIL.n422 B 0.010524f
C535 VTAIL.n423 B 0.011143f
C536 VTAIL.n424 B 0.024875f
C537 VTAIL.n425 B 0.024875f
C538 VTAIL.n426 B 0.024875f
C539 VTAIL.n427 B 0.010834f
C540 VTAIL.n428 B 0.010524f
C541 VTAIL.n429 B 0.019585f
C542 VTAIL.n430 B 0.019585f
C543 VTAIL.n431 B 0.010524f
C544 VTAIL.n432 B 0.011143f
C545 VTAIL.n433 B 0.024875f
C546 VTAIL.n434 B 0.055721f
C547 VTAIL.n435 B 0.011143f
C548 VTAIL.n436 B 0.010524f
C549 VTAIL.n437 B 0.050621f
C550 VTAIL.n438 B 0.031526f
C551 VTAIL.n439 B 1.01331f
C552 VN.n0 B 0.03346f
C553 VN.t0 B 1.2071f
C554 VN.n1 B 0.056167f
C555 VN.n2 B 0.03346f
C556 VN.n3 B 0.035705f
C557 VN.t1 B 1.27803f
C558 VN.t4 B 1.2071f
C559 VN.n4 B 0.491043f
C560 VN.n5 B 0.528367f
C561 VN.n6 B 0.175542f
C562 VN.n7 B 0.03346f
C563 VN.n8 B 0.048639f
C564 VN.n9 B 0.048639f
C565 VN.t2 B 1.2071f
C566 VN.n10 B 0.446647f
C567 VN.n11 B 0.035705f
C568 VN.n12 B 0.03346f
C569 VN.n13 B 0.03346f
C570 VN.n14 B 0.03346f
C571 VN.n15 B 0.032568f
C572 VN.n16 B 0.048537f
C573 VN.n17 B 0.50478f
C574 VN.n18 B 0.031071f
C575 VN.n19 B 0.03346f
C576 VN.t7 B 1.2071f
C577 VN.n20 B 0.056167f
C578 VN.n21 B 0.03346f
C579 VN.t6 B 1.2071f
C580 VN.n22 B 0.446647f
C581 VN.n23 B 0.035705f
C582 VN.t5 B 1.27803f
C583 VN.t3 B 1.2071f
C584 VN.n24 B 0.491043f
C585 VN.n25 B 0.528367f
C586 VN.n26 B 0.175542f
C587 VN.n27 B 0.03346f
C588 VN.n28 B 0.048639f
C589 VN.n29 B 0.048639f
C590 VN.n30 B 0.035705f
C591 VN.n31 B 0.03346f
C592 VN.n32 B 0.03346f
C593 VN.n33 B 0.03346f
C594 VN.n34 B 0.032568f
C595 VN.n35 B 0.048537f
C596 VN.n36 B 0.50478f
C597 VN.n37 B 1.48206f
.ends

