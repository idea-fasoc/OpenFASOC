* NGSPICE file created from diff_pair_sample_0100.ext - technology: sky130A

.subckt diff_pair_sample_0100 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=6.1074 ps=32.1 w=15.66 l=1.45
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=0 ps=0 w=15.66 l=1.45
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=0 ps=0 w=15.66 l=1.45
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=0 ps=0 w=15.66 l=1.45
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=0 ps=0 w=15.66 l=1.45
X5 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=6.1074 ps=32.1 w=15.66 l=1.45
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=6.1074 ps=32.1 w=15.66 l=1.45
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1074 pd=32.1 as=6.1074 ps=32.1 w=15.66 l=1.45
R0 VP.n0 VP.t1 412.356
R1 VP.n0 VP.t0 367.976
R2 VP VP.n0 0.146778
R3 VTAIL.n1 VTAIL.t1 44.2302
R4 VTAIL.n3 VTAIL.t0 44.2301
R5 VTAIL.n0 VTAIL.t3 44.2301
R6 VTAIL.n2 VTAIL.t2 44.2301
R7 VTAIL.n1 VTAIL.n0 28.9358
R8 VTAIL.n3 VTAIL.n2 27.4014
R9 VTAIL.n2 VTAIL.n1 1.23757
R10 VTAIL VTAIL.n0 0.912138
R11 VTAIL VTAIL.n3 0.325931
R12 VDD1 VDD1.t1 102.046
R13 VDD1 VDD1.t0 61.3507
R14 B.n504 B.n503 585
R15 B.n506 B.n98 585
R16 B.n509 B.n508 585
R17 B.n510 B.n97 585
R18 B.n512 B.n511 585
R19 B.n514 B.n96 585
R20 B.n517 B.n516 585
R21 B.n518 B.n95 585
R22 B.n520 B.n519 585
R23 B.n522 B.n94 585
R24 B.n525 B.n524 585
R25 B.n526 B.n93 585
R26 B.n528 B.n527 585
R27 B.n530 B.n92 585
R28 B.n533 B.n532 585
R29 B.n534 B.n91 585
R30 B.n536 B.n535 585
R31 B.n538 B.n90 585
R32 B.n541 B.n540 585
R33 B.n542 B.n89 585
R34 B.n544 B.n543 585
R35 B.n546 B.n88 585
R36 B.n549 B.n548 585
R37 B.n550 B.n87 585
R38 B.n552 B.n551 585
R39 B.n554 B.n86 585
R40 B.n557 B.n556 585
R41 B.n558 B.n85 585
R42 B.n560 B.n559 585
R43 B.n562 B.n84 585
R44 B.n565 B.n564 585
R45 B.n566 B.n83 585
R46 B.n568 B.n567 585
R47 B.n570 B.n82 585
R48 B.n573 B.n572 585
R49 B.n574 B.n81 585
R50 B.n576 B.n575 585
R51 B.n578 B.n80 585
R52 B.n581 B.n580 585
R53 B.n582 B.n79 585
R54 B.n584 B.n583 585
R55 B.n586 B.n78 585
R56 B.n589 B.n588 585
R57 B.n590 B.n77 585
R58 B.n592 B.n591 585
R59 B.n594 B.n76 585
R60 B.n597 B.n596 585
R61 B.n598 B.n75 585
R62 B.n600 B.n599 585
R63 B.n602 B.n74 585
R64 B.n604 B.n603 585
R65 B.n606 B.n605 585
R66 B.n609 B.n608 585
R67 B.n610 B.n69 585
R68 B.n612 B.n611 585
R69 B.n614 B.n68 585
R70 B.n617 B.n616 585
R71 B.n618 B.n67 585
R72 B.n620 B.n619 585
R73 B.n622 B.n66 585
R74 B.n625 B.n624 585
R75 B.n626 B.n63 585
R76 B.n629 B.n628 585
R77 B.n631 B.n62 585
R78 B.n634 B.n633 585
R79 B.n635 B.n61 585
R80 B.n637 B.n636 585
R81 B.n639 B.n60 585
R82 B.n642 B.n641 585
R83 B.n643 B.n59 585
R84 B.n645 B.n644 585
R85 B.n647 B.n58 585
R86 B.n650 B.n649 585
R87 B.n651 B.n57 585
R88 B.n653 B.n652 585
R89 B.n655 B.n56 585
R90 B.n658 B.n657 585
R91 B.n659 B.n55 585
R92 B.n661 B.n660 585
R93 B.n663 B.n54 585
R94 B.n666 B.n665 585
R95 B.n667 B.n53 585
R96 B.n669 B.n668 585
R97 B.n671 B.n52 585
R98 B.n674 B.n673 585
R99 B.n675 B.n51 585
R100 B.n677 B.n676 585
R101 B.n679 B.n50 585
R102 B.n682 B.n681 585
R103 B.n683 B.n49 585
R104 B.n685 B.n684 585
R105 B.n687 B.n48 585
R106 B.n690 B.n689 585
R107 B.n691 B.n47 585
R108 B.n693 B.n692 585
R109 B.n695 B.n46 585
R110 B.n698 B.n697 585
R111 B.n699 B.n45 585
R112 B.n701 B.n700 585
R113 B.n703 B.n44 585
R114 B.n706 B.n705 585
R115 B.n707 B.n43 585
R116 B.n709 B.n708 585
R117 B.n711 B.n42 585
R118 B.n714 B.n713 585
R119 B.n715 B.n41 585
R120 B.n717 B.n716 585
R121 B.n719 B.n40 585
R122 B.n722 B.n721 585
R123 B.n723 B.n39 585
R124 B.n725 B.n724 585
R125 B.n727 B.n38 585
R126 B.n730 B.n729 585
R127 B.n731 B.n37 585
R128 B.n502 B.n35 585
R129 B.n734 B.n35 585
R130 B.n501 B.n34 585
R131 B.n735 B.n34 585
R132 B.n500 B.n33 585
R133 B.n736 B.n33 585
R134 B.n499 B.n498 585
R135 B.n498 B.n29 585
R136 B.n497 B.n28 585
R137 B.n742 B.n28 585
R138 B.n496 B.n27 585
R139 B.n743 B.n27 585
R140 B.n495 B.n26 585
R141 B.n744 B.n26 585
R142 B.n494 B.n493 585
R143 B.n493 B.n22 585
R144 B.n492 B.n21 585
R145 B.n750 B.n21 585
R146 B.n491 B.n20 585
R147 B.n751 B.n20 585
R148 B.n490 B.n19 585
R149 B.n752 B.n19 585
R150 B.n489 B.n488 585
R151 B.n488 B.n15 585
R152 B.n487 B.n14 585
R153 B.n758 B.n14 585
R154 B.n486 B.n13 585
R155 B.n759 B.n13 585
R156 B.n485 B.n12 585
R157 B.n760 B.n12 585
R158 B.n484 B.n483 585
R159 B.n483 B.n482 585
R160 B.n481 B.n480 585
R161 B.n481 B.n8 585
R162 B.n479 B.n7 585
R163 B.n767 B.n7 585
R164 B.n478 B.n6 585
R165 B.n768 B.n6 585
R166 B.n477 B.n5 585
R167 B.n769 B.n5 585
R168 B.n476 B.n475 585
R169 B.n475 B.n4 585
R170 B.n474 B.n99 585
R171 B.n474 B.n473 585
R172 B.n464 B.n100 585
R173 B.n101 B.n100 585
R174 B.n466 B.n465 585
R175 B.n467 B.n466 585
R176 B.n463 B.n106 585
R177 B.n106 B.n105 585
R178 B.n462 B.n461 585
R179 B.n461 B.n460 585
R180 B.n108 B.n107 585
R181 B.n109 B.n108 585
R182 B.n453 B.n452 585
R183 B.n454 B.n453 585
R184 B.n451 B.n114 585
R185 B.n114 B.n113 585
R186 B.n450 B.n449 585
R187 B.n449 B.n448 585
R188 B.n116 B.n115 585
R189 B.n117 B.n116 585
R190 B.n441 B.n440 585
R191 B.n442 B.n441 585
R192 B.n439 B.n121 585
R193 B.n125 B.n121 585
R194 B.n438 B.n437 585
R195 B.n437 B.n436 585
R196 B.n123 B.n122 585
R197 B.n124 B.n123 585
R198 B.n429 B.n428 585
R199 B.n430 B.n429 585
R200 B.n427 B.n130 585
R201 B.n130 B.n129 585
R202 B.n426 B.n425 585
R203 B.n425 B.n424 585
R204 B.n421 B.n134 585
R205 B.n420 B.n419 585
R206 B.n417 B.n135 585
R207 B.n417 B.n133 585
R208 B.n416 B.n415 585
R209 B.n414 B.n413 585
R210 B.n412 B.n137 585
R211 B.n410 B.n409 585
R212 B.n408 B.n138 585
R213 B.n407 B.n406 585
R214 B.n404 B.n139 585
R215 B.n402 B.n401 585
R216 B.n400 B.n140 585
R217 B.n399 B.n398 585
R218 B.n396 B.n141 585
R219 B.n394 B.n393 585
R220 B.n392 B.n142 585
R221 B.n391 B.n390 585
R222 B.n388 B.n143 585
R223 B.n386 B.n385 585
R224 B.n384 B.n144 585
R225 B.n383 B.n382 585
R226 B.n380 B.n145 585
R227 B.n378 B.n377 585
R228 B.n376 B.n146 585
R229 B.n375 B.n374 585
R230 B.n372 B.n147 585
R231 B.n370 B.n369 585
R232 B.n368 B.n148 585
R233 B.n367 B.n366 585
R234 B.n364 B.n149 585
R235 B.n362 B.n361 585
R236 B.n360 B.n150 585
R237 B.n359 B.n358 585
R238 B.n356 B.n151 585
R239 B.n354 B.n353 585
R240 B.n352 B.n152 585
R241 B.n351 B.n350 585
R242 B.n348 B.n153 585
R243 B.n346 B.n345 585
R244 B.n344 B.n154 585
R245 B.n343 B.n342 585
R246 B.n340 B.n155 585
R247 B.n338 B.n337 585
R248 B.n336 B.n156 585
R249 B.n335 B.n334 585
R250 B.n332 B.n157 585
R251 B.n330 B.n329 585
R252 B.n328 B.n158 585
R253 B.n327 B.n326 585
R254 B.n324 B.n159 585
R255 B.n322 B.n321 585
R256 B.n320 B.n160 585
R257 B.n318 B.n317 585
R258 B.n315 B.n163 585
R259 B.n313 B.n312 585
R260 B.n311 B.n164 585
R261 B.n310 B.n309 585
R262 B.n307 B.n165 585
R263 B.n305 B.n304 585
R264 B.n303 B.n166 585
R265 B.n302 B.n301 585
R266 B.n299 B.n167 585
R267 B.n297 B.n296 585
R268 B.n295 B.n168 585
R269 B.n294 B.n293 585
R270 B.n291 B.n172 585
R271 B.n289 B.n288 585
R272 B.n287 B.n173 585
R273 B.n286 B.n285 585
R274 B.n283 B.n174 585
R275 B.n281 B.n280 585
R276 B.n279 B.n175 585
R277 B.n278 B.n277 585
R278 B.n275 B.n176 585
R279 B.n273 B.n272 585
R280 B.n271 B.n177 585
R281 B.n270 B.n269 585
R282 B.n267 B.n178 585
R283 B.n265 B.n264 585
R284 B.n263 B.n179 585
R285 B.n262 B.n261 585
R286 B.n259 B.n180 585
R287 B.n257 B.n256 585
R288 B.n255 B.n181 585
R289 B.n254 B.n253 585
R290 B.n251 B.n182 585
R291 B.n249 B.n248 585
R292 B.n247 B.n183 585
R293 B.n246 B.n245 585
R294 B.n243 B.n184 585
R295 B.n241 B.n240 585
R296 B.n239 B.n185 585
R297 B.n238 B.n237 585
R298 B.n235 B.n186 585
R299 B.n233 B.n232 585
R300 B.n231 B.n187 585
R301 B.n230 B.n229 585
R302 B.n227 B.n188 585
R303 B.n225 B.n224 585
R304 B.n223 B.n189 585
R305 B.n222 B.n221 585
R306 B.n219 B.n190 585
R307 B.n217 B.n216 585
R308 B.n215 B.n191 585
R309 B.n214 B.n213 585
R310 B.n211 B.n192 585
R311 B.n209 B.n208 585
R312 B.n207 B.n193 585
R313 B.n206 B.n205 585
R314 B.n203 B.n194 585
R315 B.n201 B.n200 585
R316 B.n199 B.n195 585
R317 B.n198 B.n197 585
R318 B.n132 B.n131 585
R319 B.n133 B.n132 585
R320 B.n423 B.n422 585
R321 B.n424 B.n423 585
R322 B.n128 B.n127 585
R323 B.n129 B.n128 585
R324 B.n432 B.n431 585
R325 B.n431 B.n430 585
R326 B.n433 B.n126 585
R327 B.n126 B.n124 585
R328 B.n435 B.n434 585
R329 B.n436 B.n435 585
R330 B.n120 B.n119 585
R331 B.n125 B.n120 585
R332 B.n444 B.n443 585
R333 B.n443 B.n442 585
R334 B.n445 B.n118 585
R335 B.n118 B.n117 585
R336 B.n447 B.n446 585
R337 B.n448 B.n447 585
R338 B.n112 B.n111 585
R339 B.n113 B.n112 585
R340 B.n456 B.n455 585
R341 B.n455 B.n454 585
R342 B.n457 B.n110 585
R343 B.n110 B.n109 585
R344 B.n459 B.n458 585
R345 B.n460 B.n459 585
R346 B.n104 B.n103 585
R347 B.n105 B.n104 585
R348 B.n469 B.n468 585
R349 B.n468 B.n467 585
R350 B.n470 B.n102 585
R351 B.n102 B.n101 585
R352 B.n472 B.n471 585
R353 B.n473 B.n472 585
R354 B.n3 B.n0 585
R355 B.n4 B.n3 585
R356 B.n766 B.n1 585
R357 B.n767 B.n766 585
R358 B.n765 B.n764 585
R359 B.n765 B.n8 585
R360 B.n763 B.n9 585
R361 B.n482 B.n9 585
R362 B.n762 B.n761 585
R363 B.n761 B.n760 585
R364 B.n11 B.n10 585
R365 B.n759 B.n11 585
R366 B.n757 B.n756 585
R367 B.n758 B.n757 585
R368 B.n755 B.n16 585
R369 B.n16 B.n15 585
R370 B.n754 B.n753 585
R371 B.n753 B.n752 585
R372 B.n18 B.n17 585
R373 B.n751 B.n18 585
R374 B.n749 B.n748 585
R375 B.n750 B.n749 585
R376 B.n747 B.n23 585
R377 B.n23 B.n22 585
R378 B.n746 B.n745 585
R379 B.n745 B.n744 585
R380 B.n25 B.n24 585
R381 B.n743 B.n25 585
R382 B.n741 B.n740 585
R383 B.n742 B.n741 585
R384 B.n739 B.n30 585
R385 B.n30 B.n29 585
R386 B.n738 B.n737 585
R387 B.n737 B.n736 585
R388 B.n32 B.n31 585
R389 B.n735 B.n32 585
R390 B.n733 B.n732 585
R391 B.n734 B.n733 585
R392 B.n770 B.n769 585
R393 B.n768 B.n2 585
R394 B.n733 B.n37 540.549
R395 B.n504 B.n35 540.549
R396 B.n425 B.n132 540.549
R397 B.n423 B.n134 540.549
R398 B.n64 B.t6 465.529
R399 B.n70 B.t2 465.529
R400 B.n169 B.t13 465.529
R401 B.n161 B.t9 465.529
R402 B.n505 B.n36 256.663
R403 B.n507 B.n36 256.663
R404 B.n513 B.n36 256.663
R405 B.n515 B.n36 256.663
R406 B.n521 B.n36 256.663
R407 B.n523 B.n36 256.663
R408 B.n529 B.n36 256.663
R409 B.n531 B.n36 256.663
R410 B.n537 B.n36 256.663
R411 B.n539 B.n36 256.663
R412 B.n545 B.n36 256.663
R413 B.n547 B.n36 256.663
R414 B.n553 B.n36 256.663
R415 B.n555 B.n36 256.663
R416 B.n561 B.n36 256.663
R417 B.n563 B.n36 256.663
R418 B.n569 B.n36 256.663
R419 B.n571 B.n36 256.663
R420 B.n577 B.n36 256.663
R421 B.n579 B.n36 256.663
R422 B.n585 B.n36 256.663
R423 B.n587 B.n36 256.663
R424 B.n593 B.n36 256.663
R425 B.n595 B.n36 256.663
R426 B.n601 B.n36 256.663
R427 B.n73 B.n36 256.663
R428 B.n607 B.n36 256.663
R429 B.n613 B.n36 256.663
R430 B.n615 B.n36 256.663
R431 B.n621 B.n36 256.663
R432 B.n623 B.n36 256.663
R433 B.n630 B.n36 256.663
R434 B.n632 B.n36 256.663
R435 B.n638 B.n36 256.663
R436 B.n640 B.n36 256.663
R437 B.n646 B.n36 256.663
R438 B.n648 B.n36 256.663
R439 B.n654 B.n36 256.663
R440 B.n656 B.n36 256.663
R441 B.n662 B.n36 256.663
R442 B.n664 B.n36 256.663
R443 B.n670 B.n36 256.663
R444 B.n672 B.n36 256.663
R445 B.n678 B.n36 256.663
R446 B.n680 B.n36 256.663
R447 B.n686 B.n36 256.663
R448 B.n688 B.n36 256.663
R449 B.n694 B.n36 256.663
R450 B.n696 B.n36 256.663
R451 B.n702 B.n36 256.663
R452 B.n704 B.n36 256.663
R453 B.n710 B.n36 256.663
R454 B.n712 B.n36 256.663
R455 B.n718 B.n36 256.663
R456 B.n720 B.n36 256.663
R457 B.n726 B.n36 256.663
R458 B.n728 B.n36 256.663
R459 B.n418 B.n133 256.663
R460 B.n136 B.n133 256.663
R461 B.n411 B.n133 256.663
R462 B.n405 B.n133 256.663
R463 B.n403 B.n133 256.663
R464 B.n397 B.n133 256.663
R465 B.n395 B.n133 256.663
R466 B.n389 B.n133 256.663
R467 B.n387 B.n133 256.663
R468 B.n381 B.n133 256.663
R469 B.n379 B.n133 256.663
R470 B.n373 B.n133 256.663
R471 B.n371 B.n133 256.663
R472 B.n365 B.n133 256.663
R473 B.n363 B.n133 256.663
R474 B.n357 B.n133 256.663
R475 B.n355 B.n133 256.663
R476 B.n349 B.n133 256.663
R477 B.n347 B.n133 256.663
R478 B.n341 B.n133 256.663
R479 B.n339 B.n133 256.663
R480 B.n333 B.n133 256.663
R481 B.n331 B.n133 256.663
R482 B.n325 B.n133 256.663
R483 B.n323 B.n133 256.663
R484 B.n316 B.n133 256.663
R485 B.n314 B.n133 256.663
R486 B.n308 B.n133 256.663
R487 B.n306 B.n133 256.663
R488 B.n300 B.n133 256.663
R489 B.n298 B.n133 256.663
R490 B.n292 B.n133 256.663
R491 B.n290 B.n133 256.663
R492 B.n284 B.n133 256.663
R493 B.n282 B.n133 256.663
R494 B.n276 B.n133 256.663
R495 B.n274 B.n133 256.663
R496 B.n268 B.n133 256.663
R497 B.n266 B.n133 256.663
R498 B.n260 B.n133 256.663
R499 B.n258 B.n133 256.663
R500 B.n252 B.n133 256.663
R501 B.n250 B.n133 256.663
R502 B.n244 B.n133 256.663
R503 B.n242 B.n133 256.663
R504 B.n236 B.n133 256.663
R505 B.n234 B.n133 256.663
R506 B.n228 B.n133 256.663
R507 B.n226 B.n133 256.663
R508 B.n220 B.n133 256.663
R509 B.n218 B.n133 256.663
R510 B.n212 B.n133 256.663
R511 B.n210 B.n133 256.663
R512 B.n204 B.n133 256.663
R513 B.n202 B.n133 256.663
R514 B.n196 B.n133 256.663
R515 B.n772 B.n771 256.663
R516 B.n729 B.n727 163.367
R517 B.n725 B.n39 163.367
R518 B.n721 B.n719 163.367
R519 B.n717 B.n41 163.367
R520 B.n713 B.n711 163.367
R521 B.n709 B.n43 163.367
R522 B.n705 B.n703 163.367
R523 B.n701 B.n45 163.367
R524 B.n697 B.n695 163.367
R525 B.n693 B.n47 163.367
R526 B.n689 B.n687 163.367
R527 B.n685 B.n49 163.367
R528 B.n681 B.n679 163.367
R529 B.n677 B.n51 163.367
R530 B.n673 B.n671 163.367
R531 B.n669 B.n53 163.367
R532 B.n665 B.n663 163.367
R533 B.n661 B.n55 163.367
R534 B.n657 B.n655 163.367
R535 B.n653 B.n57 163.367
R536 B.n649 B.n647 163.367
R537 B.n645 B.n59 163.367
R538 B.n641 B.n639 163.367
R539 B.n637 B.n61 163.367
R540 B.n633 B.n631 163.367
R541 B.n629 B.n63 163.367
R542 B.n624 B.n622 163.367
R543 B.n620 B.n67 163.367
R544 B.n616 B.n614 163.367
R545 B.n612 B.n69 163.367
R546 B.n608 B.n606 163.367
R547 B.n603 B.n602 163.367
R548 B.n600 B.n75 163.367
R549 B.n596 B.n594 163.367
R550 B.n592 B.n77 163.367
R551 B.n588 B.n586 163.367
R552 B.n584 B.n79 163.367
R553 B.n580 B.n578 163.367
R554 B.n576 B.n81 163.367
R555 B.n572 B.n570 163.367
R556 B.n568 B.n83 163.367
R557 B.n564 B.n562 163.367
R558 B.n560 B.n85 163.367
R559 B.n556 B.n554 163.367
R560 B.n552 B.n87 163.367
R561 B.n548 B.n546 163.367
R562 B.n544 B.n89 163.367
R563 B.n540 B.n538 163.367
R564 B.n536 B.n91 163.367
R565 B.n532 B.n530 163.367
R566 B.n528 B.n93 163.367
R567 B.n524 B.n522 163.367
R568 B.n520 B.n95 163.367
R569 B.n516 B.n514 163.367
R570 B.n512 B.n97 163.367
R571 B.n508 B.n506 163.367
R572 B.n425 B.n130 163.367
R573 B.n429 B.n130 163.367
R574 B.n429 B.n123 163.367
R575 B.n437 B.n123 163.367
R576 B.n437 B.n121 163.367
R577 B.n441 B.n121 163.367
R578 B.n441 B.n116 163.367
R579 B.n449 B.n116 163.367
R580 B.n449 B.n114 163.367
R581 B.n453 B.n114 163.367
R582 B.n453 B.n108 163.367
R583 B.n461 B.n108 163.367
R584 B.n461 B.n106 163.367
R585 B.n466 B.n106 163.367
R586 B.n466 B.n100 163.367
R587 B.n474 B.n100 163.367
R588 B.n475 B.n474 163.367
R589 B.n475 B.n5 163.367
R590 B.n6 B.n5 163.367
R591 B.n7 B.n6 163.367
R592 B.n481 B.n7 163.367
R593 B.n483 B.n481 163.367
R594 B.n483 B.n12 163.367
R595 B.n13 B.n12 163.367
R596 B.n14 B.n13 163.367
R597 B.n488 B.n14 163.367
R598 B.n488 B.n19 163.367
R599 B.n20 B.n19 163.367
R600 B.n21 B.n20 163.367
R601 B.n493 B.n21 163.367
R602 B.n493 B.n26 163.367
R603 B.n27 B.n26 163.367
R604 B.n28 B.n27 163.367
R605 B.n498 B.n28 163.367
R606 B.n498 B.n33 163.367
R607 B.n34 B.n33 163.367
R608 B.n35 B.n34 163.367
R609 B.n419 B.n417 163.367
R610 B.n417 B.n416 163.367
R611 B.n413 B.n412 163.367
R612 B.n410 B.n138 163.367
R613 B.n406 B.n404 163.367
R614 B.n402 B.n140 163.367
R615 B.n398 B.n396 163.367
R616 B.n394 B.n142 163.367
R617 B.n390 B.n388 163.367
R618 B.n386 B.n144 163.367
R619 B.n382 B.n380 163.367
R620 B.n378 B.n146 163.367
R621 B.n374 B.n372 163.367
R622 B.n370 B.n148 163.367
R623 B.n366 B.n364 163.367
R624 B.n362 B.n150 163.367
R625 B.n358 B.n356 163.367
R626 B.n354 B.n152 163.367
R627 B.n350 B.n348 163.367
R628 B.n346 B.n154 163.367
R629 B.n342 B.n340 163.367
R630 B.n338 B.n156 163.367
R631 B.n334 B.n332 163.367
R632 B.n330 B.n158 163.367
R633 B.n326 B.n324 163.367
R634 B.n322 B.n160 163.367
R635 B.n317 B.n315 163.367
R636 B.n313 B.n164 163.367
R637 B.n309 B.n307 163.367
R638 B.n305 B.n166 163.367
R639 B.n301 B.n299 163.367
R640 B.n297 B.n168 163.367
R641 B.n293 B.n291 163.367
R642 B.n289 B.n173 163.367
R643 B.n285 B.n283 163.367
R644 B.n281 B.n175 163.367
R645 B.n277 B.n275 163.367
R646 B.n273 B.n177 163.367
R647 B.n269 B.n267 163.367
R648 B.n265 B.n179 163.367
R649 B.n261 B.n259 163.367
R650 B.n257 B.n181 163.367
R651 B.n253 B.n251 163.367
R652 B.n249 B.n183 163.367
R653 B.n245 B.n243 163.367
R654 B.n241 B.n185 163.367
R655 B.n237 B.n235 163.367
R656 B.n233 B.n187 163.367
R657 B.n229 B.n227 163.367
R658 B.n225 B.n189 163.367
R659 B.n221 B.n219 163.367
R660 B.n217 B.n191 163.367
R661 B.n213 B.n211 163.367
R662 B.n209 B.n193 163.367
R663 B.n205 B.n203 163.367
R664 B.n201 B.n195 163.367
R665 B.n197 B.n132 163.367
R666 B.n423 B.n128 163.367
R667 B.n431 B.n128 163.367
R668 B.n431 B.n126 163.367
R669 B.n435 B.n126 163.367
R670 B.n435 B.n120 163.367
R671 B.n443 B.n120 163.367
R672 B.n443 B.n118 163.367
R673 B.n447 B.n118 163.367
R674 B.n447 B.n112 163.367
R675 B.n455 B.n112 163.367
R676 B.n455 B.n110 163.367
R677 B.n459 B.n110 163.367
R678 B.n459 B.n104 163.367
R679 B.n468 B.n104 163.367
R680 B.n468 B.n102 163.367
R681 B.n472 B.n102 163.367
R682 B.n472 B.n3 163.367
R683 B.n770 B.n3 163.367
R684 B.n766 B.n2 163.367
R685 B.n766 B.n765 163.367
R686 B.n765 B.n9 163.367
R687 B.n761 B.n9 163.367
R688 B.n761 B.n11 163.367
R689 B.n757 B.n11 163.367
R690 B.n757 B.n16 163.367
R691 B.n753 B.n16 163.367
R692 B.n753 B.n18 163.367
R693 B.n749 B.n18 163.367
R694 B.n749 B.n23 163.367
R695 B.n745 B.n23 163.367
R696 B.n745 B.n25 163.367
R697 B.n741 B.n25 163.367
R698 B.n741 B.n30 163.367
R699 B.n737 B.n30 163.367
R700 B.n737 B.n32 163.367
R701 B.n733 B.n32 163.367
R702 B.n70 B.t4 102.319
R703 B.n169 B.t15 102.319
R704 B.n64 B.t7 102.299
R705 B.n161 B.t12 102.299
R706 B.n728 B.n37 71.676
R707 B.n727 B.n726 71.676
R708 B.n720 B.n39 71.676
R709 B.n719 B.n718 71.676
R710 B.n712 B.n41 71.676
R711 B.n711 B.n710 71.676
R712 B.n704 B.n43 71.676
R713 B.n703 B.n702 71.676
R714 B.n696 B.n45 71.676
R715 B.n695 B.n694 71.676
R716 B.n688 B.n47 71.676
R717 B.n687 B.n686 71.676
R718 B.n680 B.n49 71.676
R719 B.n679 B.n678 71.676
R720 B.n672 B.n51 71.676
R721 B.n671 B.n670 71.676
R722 B.n664 B.n53 71.676
R723 B.n663 B.n662 71.676
R724 B.n656 B.n55 71.676
R725 B.n655 B.n654 71.676
R726 B.n648 B.n57 71.676
R727 B.n647 B.n646 71.676
R728 B.n640 B.n59 71.676
R729 B.n639 B.n638 71.676
R730 B.n632 B.n61 71.676
R731 B.n631 B.n630 71.676
R732 B.n623 B.n63 71.676
R733 B.n622 B.n621 71.676
R734 B.n615 B.n67 71.676
R735 B.n614 B.n613 71.676
R736 B.n607 B.n69 71.676
R737 B.n606 B.n73 71.676
R738 B.n602 B.n601 71.676
R739 B.n595 B.n75 71.676
R740 B.n594 B.n593 71.676
R741 B.n587 B.n77 71.676
R742 B.n586 B.n585 71.676
R743 B.n579 B.n79 71.676
R744 B.n578 B.n577 71.676
R745 B.n571 B.n81 71.676
R746 B.n570 B.n569 71.676
R747 B.n563 B.n83 71.676
R748 B.n562 B.n561 71.676
R749 B.n555 B.n85 71.676
R750 B.n554 B.n553 71.676
R751 B.n547 B.n87 71.676
R752 B.n546 B.n545 71.676
R753 B.n539 B.n89 71.676
R754 B.n538 B.n537 71.676
R755 B.n531 B.n91 71.676
R756 B.n530 B.n529 71.676
R757 B.n523 B.n93 71.676
R758 B.n522 B.n521 71.676
R759 B.n515 B.n95 71.676
R760 B.n514 B.n513 71.676
R761 B.n507 B.n97 71.676
R762 B.n506 B.n505 71.676
R763 B.n505 B.n504 71.676
R764 B.n508 B.n507 71.676
R765 B.n513 B.n512 71.676
R766 B.n516 B.n515 71.676
R767 B.n521 B.n520 71.676
R768 B.n524 B.n523 71.676
R769 B.n529 B.n528 71.676
R770 B.n532 B.n531 71.676
R771 B.n537 B.n536 71.676
R772 B.n540 B.n539 71.676
R773 B.n545 B.n544 71.676
R774 B.n548 B.n547 71.676
R775 B.n553 B.n552 71.676
R776 B.n556 B.n555 71.676
R777 B.n561 B.n560 71.676
R778 B.n564 B.n563 71.676
R779 B.n569 B.n568 71.676
R780 B.n572 B.n571 71.676
R781 B.n577 B.n576 71.676
R782 B.n580 B.n579 71.676
R783 B.n585 B.n584 71.676
R784 B.n588 B.n587 71.676
R785 B.n593 B.n592 71.676
R786 B.n596 B.n595 71.676
R787 B.n601 B.n600 71.676
R788 B.n603 B.n73 71.676
R789 B.n608 B.n607 71.676
R790 B.n613 B.n612 71.676
R791 B.n616 B.n615 71.676
R792 B.n621 B.n620 71.676
R793 B.n624 B.n623 71.676
R794 B.n630 B.n629 71.676
R795 B.n633 B.n632 71.676
R796 B.n638 B.n637 71.676
R797 B.n641 B.n640 71.676
R798 B.n646 B.n645 71.676
R799 B.n649 B.n648 71.676
R800 B.n654 B.n653 71.676
R801 B.n657 B.n656 71.676
R802 B.n662 B.n661 71.676
R803 B.n665 B.n664 71.676
R804 B.n670 B.n669 71.676
R805 B.n673 B.n672 71.676
R806 B.n678 B.n677 71.676
R807 B.n681 B.n680 71.676
R808 B.n686 B.n685 71.676
R809 B.n689 B.n688 71.676
R810 B.n694 B.n693 71.676
R811 B.n697 B.n696 71.676
R812 B.n702 B.n701 71.676
R813 B.n705 B.n704 71.676
R814 B.n710 B.n709 71.676
R815 B.n713 B.n712 71.676
R816 B.n718 B.n717 71.676
R817 B.n721 B.n720 71.676
R818 B.n726 B.n725 71.676
R819 B.n729 B.n728 71.676
R820 B.n418 B.n134 71.676
R821 B.n416 B.n136 71.676
R822 B.n412 B.n411 71.676
R823 B.n405 B.n138 71.676
R824 B.n404 B.n403 71.676
R825 B.n397 B.n140 71.676
R826 B.n396 B.n395 71.676
R827 B.n389 B.n142 71.676
R828 B.n388 B.n387 71.676
R829 B.n381 B.n144 71.676
R830 B.n380 B.n379 71.676
R831 B.n373 B.n146 71.676
R832 B.n372 B.n371 71.676
R833 B.n365 B.n148 71.676
R834 B.n364 B.n363 71.676
R835 B.n357 B.n150 71.676
R836 B.n356 B.n355 71.676
R837 B.n349 B.n152 71.676
R838 B.n348 B.n347 71.676
R839 B.n341 B.n154 71.676
R840 B.n340 B.n339 71.676
R841 B.n333 B.n156 71.676
R842 B.n332 B.n331 71.676
R843 B.n325 B.n158 71.676
R844 B.n324 B.n323 71.676
R845 B.n316 B.n160 71.676
R846 B.n315 B.n314 71.676
R847 B.n308 B.n164 71.676
R848 B.n307 B.n306 71.676
R849 B.n300 B.n166 71.676
R850 B.n299 B.n298 71.676
R851 B.n292 B.n168 71.676
R852 B.n291 B.n290 71.676
R853 B.n284 B.n173 71.676
R854 B.n283 B.n282 71.676
R855 B.n276 B.n175 71.676
R856 B.n275 B.n274 71.676
R857 B.n268 B.n177 71.676
R858 B.n267 B.n266 71.676
R859 B.n260 B.n179 71.676
R860 B.n259 B.n258 71.676
R861 B.n252 B.n181 71.676
R862 B.n251 B.n250 71.676
R863 B.n244 B.n183 71.676
R864 B.n243 B.n242 71.676
R865 B.n236 B.n185 71.676
R866 B.n235 B.n234 71.676
R867 B.n228 B.n187 71.676
R868 B.n227 B.n226 71.676
R869 B.n220 B.n189 71.676
R870 B.n219 B.n218 71.676
R871 B.n212 B.n191 71.676
R872 B.n211 B.n210 71.676
R873 B.n204 B.n193 71.676
R874 B.n203 B.n202 71.676
R875 B.n196 B.n195 71.676
R876 B.n419 B.n418 71.676
R877 B.n413 B.n136 71.676
R878 B.n411 B.n410 71.676
R879 B.n406 B.n405 71.676
R880 B.n403 B.n402 71.676
R881 B.n398 B.n397 71.676
R882 B.n395 B.n394 71.676
R883 B.n390 B.n389 71.676
R884 B.n387 B.n386 71.676
R885 B.n382 B.n381 71.676
R886 B.n379 B.n378 71.676
R887 B.n374 B.n373 71.676
R888 B.n371 B.n370 71.676
R889 B.n366 B.n365 71.676
R890 B.n363 B.n362 71.676
R891 B.n358 B.n357 71.676
R892 B.n355 B.n354 71.676
R893 B.n350 B.n349 71.676
R894 B.n347 B.n346 71.676
R895 B.n342 B.n341 71.676
R896 B.n339 B.n338 71.676
R897 B.n334 B.n333 71.676
R898 B.n331 B.n330 71.676
R899 B.n326 B.n325 71.676
R900 B.n323 B.n322 71.676
R901 B.n317 B.n316 71.676
R902 B.n314 B.n313 71.676
R903 B.n309 B.n308 71.676
R904 B.n306 B.n305 71.676
R905 B.n301 B.n300 71.676
R906 B.n298 B.n297 71.676
R907 B.n293 B.n292 71.676
R908 B.n290 B.n289 71.676
R909 B.n285 B.n284 71.676
R910 B.n282 B.n281 71.676
R911 B.n277 B.n276 71.676
R912 B.n274 B.n273 71.676
R913 B.n269 B.n268 71.676
R914 B.n266 B.n265 71.676
R915 B.n261 B.n260 71.676
R916 B.n258 B.n257 71.676
R917 B.n253 B.n252 71.676
R918 B.n250 B.n249 71.676
R919 B.n245 B.n244 71.676
R920 B.n242 B.n241 71.676
R921 B.n237 B.n236 71.676
R922 B.n234 B.n233 71.676
R923 B.n229 B.n228 71.676
R924 B.n226 B.n225 71.676
R925 B.n221 B.n220 71.676
R926 B.n218 B.n217 71.676
R927 B.n213 B.n212 71.676
R928 B.n210 B.n209 71.676
R929 B.n205 B.n204 71.676
R930 B.n202 B.n201 71.676
R931 B.n197 B.n196 71.676
R932 B.n771 B.n770 71.676
R933 B.n771 B.n2 71.676
R934 B.n71 B.t5 67.7976
R935 B.n170 B.t14 67.7976
R936 B.n424 B.n133 67.7817
R937 B.n734 B.n36 67.7817
R938 B.n65 B.t8 67.7769
R939 B.n162 B.t11 67.7769
R940 B.n627 B.n65 59.5399
R941 B.n72 B.n71 59.5399
R942 B.n171 B.n170 59.5399
R943 B.n319 B.n162 59.5399
R944 B.n424 B.n129 35.7301
R945 B.n430 B.n129 35.7301
R946 B.n430 B.n124 35.7301
R947 B.n436 B.n124 35.7301
R948 B.n436 B.n125 35.7301
R949 B.n442 B.n117 35.7301
R950 B.n448 B.n117 35.7301
R951 B.n448 B.n113 35.7301
R952 B.n454 B.n113 35.7301
R953 B.n454 B.n109 35.7301
R954 B.n460 B.n109 35.7301
R955 B.n460 B.n105 35.7301
R956 B.n467 B.n105 35.7301
R957 B.n473 B.n101 35.7301
R958 B.n473 B.n4 35.7301
R959 B.n769 B.n4 35.7301
R960 B.n769 B.n768 35.7301
R961 B.n768 B.n767 35.7301
R962 B.n767 B.n8 35.7301
R963 B.n482 B.n8 35.7301
R964 B.n760 B.n759 35.7301
R965 B.n759 B.n758 35.7301
R966 B.n758 B.n15 35.7301
R967 B.n752 B.n15 35.7301
R968 B.n752 B.n751 35.7301
R969 B.n751 B.n750 35.7301
R970 B.n750 B.n22 35.7301
R971 B.n744 B.n22 35.7301
R972 B.n743 B.n742 35.7301
R973 B.n742 B.n29 35.7301
R974 B.n736 B.n29 35.7301
R975 B.n736 B.n735 35.7301
R976 B.n735 B.n734 35.7301
R977 B.n422 B.n421 35.1225
R978 B.n426 B.n131 35.1225
R979 B.n732 B.n731 35.1225
R980 B.n503 B.n502 35.1224
R981 B.n65 B.n64 34.5217
R982 B.n71 B.n70 34.5217
R983 B.n170 B.n169 34.5217
R984 B.n162 B.n161 34.5217
R985 B.n125 B.t10 29.9503
R986 B.t3 B.n743 29.9503
R987 B.t1 B.n101 25.7469
R988 B.n482 B.t0 25.7469
R989 B B.n772 18.0485
R990 B.n422 B.n127 10.6151
R991 B.n432 B.n127 10.6151
R992 B.n433 B.n432 10.6151
R993 B.n434 B.n433 10.6151
R994 B.n434 B.n119 10.6151
R995 B.n444 B.n119 10.6151
R996 B.n445 B.n444 10.6151
R997 B.n446 B.n445 10.6151
R998 B.n446 B.n111 10.6151
R999 B.n456 B.n111 10.6151
R1000 B.n457 B.n456 10.6151
R1001 B.n458 B.n457 10.6151
R1002 B.n458 B.n103 10.6151
R1003 B.n469 B.n103 10.6151
R1004 B.n470 B.n469 10.6151
R1005 B.n471 B.n470 10.6151
R1006 B.n471 B.n0 10.6151
R1007 B.n421 B.n420 10.6151
R1008 B.n420 B.n135 10.6151
R1009 B.n415 B.n135 10.6151
R1010 B.n415 B.n414 10.6151
R1011 B.n414 B.n137 10.6151
R1012 B.n409 B.n137 10.6151
R1013 B.n409 B.n408 10.6151
R1014 B.n408 B.n407 10.6151
R1015 B.n407 B.n139 10.6151
R1016 B.n401 B.n139 10.6151
R1017 B.n401 B.n400 10.6151
R1018 B.n400 B.n399 10.6151
R1019 B.n399 B.n141 10.6151
R1020 B.n393 B.n141 10.6151
R1021 B.n393 B.n392 10.6151
R1022 B.n392 B.n391 10.6151
R1023 B.n391 B.n143 10.6151
R1024 B.n385 B.n143 10.6151
R1025 B.n385 B.n384 10.6151
R1026 B.n384 B.n383 10.6151
R1027 B.n383 B.n145 10.6151
R1028 B.n377 B.n145 10.6151
R1029 B.n377 B.n376 10.6151
R1030 B.n376 B.n375 10.6151
R1031 B.n375 B.n147 10.6151
R1032 B.n369 B.n147 10.6151
R1033 B.n369 B.n368 10.6151
R1034 B.n368 B.n367 10.6151
R1035 B.n367 B.n149 10.6151
R1036 B.n361 B.n149 10.6151
R1037 B.n361 B.n360 10.6151
R1038 B.n360 B.n359 10.6151
R1039 B.n359 B.n151 10.6151
R1040 B.n353 B.n151 10.6151
R1041 B.n353 B.n352 10.6151
R1042 B.n352 B.n351 10.6151
R1043 B.n351 B.n153 10.6151
R1044 B.n345 B.n153 10.6151
R1045 B.n345 B.n344 10.6151
R1046 B.n344 B.n343 10.6151
R1047 B.n343 B.n155 10.6151
R1048 B.n337 B.n155 10.6151
R1049 B.n337 B.n336 10.6151
R1050 B.n336 B.n335 10.6151
R1051 B.n335 B.n157 10.6151
R1052 B.n329 B.n157 10.6151
R1053 B.n329 B.n328 10.6151
R1054 B.n328 B.n327 10.6151
R1055 B.n327 B.n159 10.6151
R1056 B.n321 B.n159 10.6151
R1057 B.n321 B.n320 10.6151
R1058 B.n318 B.n163 10.6151
R1059 B.n312 B.n163 10.6151
R1060 B.n312 B.n311 10.6151
R1061 B.n311 B.n310 10.6151
R1062 B.n310 B.n165 10.6151
R1063 B.n304 B.n165 10.6151
R1064 B.n304 B.n303 10.6151
R1065 B.n303 B.n302 10.6151
R1066 B.n302 B.n167 10.6151
R1067 B.n296 B.n295 10.6151
R1068 B.n295 B.n294 10.6151
R1069 B.n294 B.n172 10.6151
R1070 B.n288 B.n172 10.6151
R1071 B.n288 B.n287 10.6151
R1072 B.n287 B.n286 10.6151
R1073 B.n286 B.n174 10.6151
R1074 B.n280 B.n174 10.6151
R1075 B.n280 B.n279 10.6151
R1076 B.n279 B.n278 10.6151
R1077 B.n278 B.n176 10.6151
R1078 B.n272 B.n176 10.6151
R1079 B.n272 B.n271 10.6151
R1080 B.n271 B.n270 10.6151
R1081 B.n270 B.n178 10.6151
R1082 B.n264 B.n178 10.6151
R1083 B.n264 B.n263 10.6151
R1084 B.n263 B.n262 10.6151
R1085 B.n262 B.n180 10.6151
R1086 B.n256 B.n180 10.6151
R1087 B.n256 B.n255 10.6151
R1088 B.n255 B.n254 10.6151
R1089 B.n254 B.n182 10.6151
R1090 B.n248 B.n182 10.6151
R1091 B.n248 B.n247 10.6151
R1092 B.n247 B.n246 10.6151
R1093 B.n246 B.n184 10.6151
R1094 B.n240 B.n184 10.6151
R1095 B.n240 B.n239 10.6151
R1096 B.n239 B.n238 10.6151
R1097 B.n238 B.n186 10.6151
R1098 B.n232 B.n186 10.6151
R1099 B.n232 B.n231 10.6151
R1100 B.n231 B.n230 10.6151
R1101 B.n230 B.n188 10.6151
R1102 B.n224 B.n188 10.6151
R1103 B.n224 B.n223 10.6151
R1104 B.n223 B.n222 10.6151
R1105 B.n222 B.n190 10.6151
R1106 B.n216 B.n190 10.6151
R1107 B.n216 B.n215 10.6151
R1108 B.n215 B.n214 10.6151
R1109 B.n214 B.n192 10.6151
R1110 B.n208 B.n192 10.6151
R1111 B.n208 B.n207 10.6151
R1112 B.n207 B.n206 10.6151
R1113 B.n206 B.n194 10.6151
R1114 B.n200 B.n194 10.6151
R1115 B.n200 B.n199 10.6151
R1116 B.n199 B.n198 10.6151
R1117 B.n198 B.n131 10.6151
R1118 B.n427 B.n426 10.6151
R1119 B.n428 B.n427 10.6151
R1120 B.n428 B.n122 10.6151
R1121 B.n438 B.n122 10.6151
R1122 B.n439 B.n438 10.6151
R1123 B.n440 B.n439 10.6151
R1124 B.n440 B.n115 10.6151
R1125 B.n450 B.n115 10.6151
R1126 B.n451 B.n450 10.6151
R1127 B.n452 B.n451 10.6151
R1128 B.n452 B.n107 10.6151
R1129 B.n462 B.n107 10.6151
R1130 B.n463 B.n462 10.6151
R1131 B.n465 B.n463 10.6151
R1132 B.n465 B.n464 10.6151
R1133 B.n464 B.n99 10.6151
R1134 B.n476 B.n99 10.6151
R1135 B.n477 B.n476 10.6151
R1136 B.n478 B.n477 10.6151
R1137 B.n479 B.n478 10.6151
R1138 B.n480 B.n479 10.6151
R1139 B.n484 B.n480 10.6151
R1140 B.n485 B.n484 10.6151
R1141 B.n486 B.n485 10.6151
R1142 B.n487 B.n486 10.6151
R1143 B.n489 B.n487 10.6151
R1144 B.n490 B.n489 10.6151
R1145 B.n491 B.n490 10.6151
R1146 B.n492 B.n491 10.6151
R1147 B.n494 B.n492 10.6151
R1148 B.n495 B.n494 10.6151
R1149 B.n496 B.n495 10.6151
R1150 B.n497 B.n496 10.6151
R1151 B.n499 B.n497 10.6151
R1152 B.n500 B.n499 10.6151
R1153 B.n501 B.n500 10.6151
R1154 B.n502 B.n501 10.6151
R1155 B.n764 B.n1 10.6151
R1156 B.n764 B.n763 10.6151
R1157 B.n763 B.n762 10.6151
R1158 B.n762 B.n10 10.6151
R1159 B.n756 B.n10 10.6151
R1160 B.n756 B.n755 10.6151
R1161 B.n755 B.n754 10.6151
R1162 B.n754 B.n17 10.6151
R1163 B.n748 B.n17 10.6151
R1164 B.n748 B.n747 10.6151
R1165 B.n747 B.n746 10.6151
R1166 B.n746 B.n24 10.6151
R1167 B.n740 B.n24 10.6151
R1168 B.n740 B.n739 10.6151
R1169 B.n739 B.n738 10.6151
R1170 B.n738 B.n31 10.6151
R1171 B.n732 B.n31 10.6151
R1172 B.n731 B.n730 10.6151
R1173 B.n730 B.n38 10.6151
R1174 B.n724 B.n38 10.6151
R1175 B.n724 B.n723 10.6151
R1176 B.n723 B.n722 10.6151
R1177 B.n722 B.n40 10.6151
R1178 B.n716 B.n40 10.6151
R1179 B.n716 B.n715 10.6151
R1180 B.n715 B.n714 10.6151
R1181 B.n714 B.n42 10.6151
R1182 B.n708 B.n42 10.6151
R1183 B.n708 B.n707 10.6151
R1184 B.n707 B.n706 10.6151
R1185 B.n706 B.n44 10.6151
R1186 B.n700 B.n44 10.6151
R1187 B.n700 B.n699 10.6151
R1188 B.n699 B.n698 10.6151
R1189 B.n698 B.n46 10.6151
R1190 B.n692 B.n46 10.6151
R1191 B.n692 B.n691 10.6151
R1192 B.n691 B.n690 10.6151
R1193 B.n690 B.n48 10.6151
R1194 B.n684 B.n48 10.6151
R1195 B.n684 B.n683 10.6151
R1196 B.n683 B.n682 10.6151
R1197 B.n682 B.n50 10.6151
R1198 B.n676 B.n50 10.6151
R1199 B.n676 B.n675 10.6151
R1200 B.n675 B.n674 10.6151
R1201 B.n674 B.n52 10.6151
R1202 B.n668 B.n52 10.6151
R1203 B.n668 B.n667 10.6151
R1204 B.n667 B.n666 10.6151
R1205 B.n666 B.n54 10.6151
R1206 B.n660 B.n54 10.6151
R1207 B.n660 B.n659 10.6151
R1208 B.n659 B.n658 10.6151
R1209 B.n658 B.n56 10.6151
R1210 B.n652 B.n56 10.6151
R1211 B.n652 B.n651 10.6151
R1212 B.n651 B.n650 10.6151
R1213 B.n650 B.n58 10.6151
R1214 B.n644 B.n58 10.6151
R1215 B.n644 B.n643 10.6151
R1216 B.n643 B.n642 10.6151
R1217 B.n642 B.n60 10.6151
R1218 B.n636 B.n60 10.6151
R1219 B.n636 B.n635 10.6151
R1220 B.n635 B.n634 10.6151
R1221 B.n634 B.n62 10.6151
R1222 B.n628 B.n62 10.6151
R1223 B.n626 B.n625 10.6151
R1224 B.n625 B.n66 10.6151
R1225 B.n619 B.n66 10.6151
R1226 B.n619 B.n618 10.6151
R1227 B.n618 B.n617 10.6151
R1228 B.n617 B.n68 10.6151
R1229 B.n611 B.n68 10.6151
R1230 B.n611 B.n610 10.6151
R1231 B.n610 B.n609 10.6151
R1232 B.n605 B.n604 10.6151
R1233 B.n604 B.n74 10.6151
R1234 B.n599 B.n74 10.6151
R1235 B.n599 B.n598 10.6151
R1236 B.n598 B.n597 10.6151
R1237 B.n597 B.n76 10.6151
R1238 B.n591 B.n76 10.6151
R1239 B.n591 B.n590 10.6151
R1240 B.n590 B.n589 10.6151
R1241 B.n589 B.n78 10.6151
R1242 B.n583 B.n78 10.6151
R1243 B.n583 B.n582 10.6151
R1244 B.n582 B.n581 10.6151
R1245 B.n581 B.n80 10.6151
R1246 B.n575 B.n80 10.6151
R1247 B.n575 B.n574 10.6151
R1248 B.n574 B.n573 10.6151
R1249 B.n573 B.n82 10.6151
R1250 B.n567 B.n82 10.6151
R1251 B.n567 B.n566 10.6151
R1252 B.n566 B.n565 10.6151
R1253 B.n565 B.n84 10.6151
R1254 B.n559 B.n84 10.6151
R1255 B.n559 B.n558 10.6151
R1256 B.n558 B.n557 10.6151
R1257 B.n557 B.n86 10.6151
R1258 B.n551 B.n86 10.6151
R1259 B.n551 B.n550 10.6151
R1260 B.n550 B.n549 10.6151
R1261 B.n549 B.n88 10.6151
R1262 B.n543 B.n88 10.6151
R1263 B.n543 B.n542 10.6151
R1264 B.n542 B.n541 10.6151
R1265 B.n541 B.n90 10.6151
R1266 B.n535 B.n90 10.6151
R1267 B.n535 B.n534 10.6151
R1268 B.n534 B.n533 10.6151
R1269 B.n533 B.n92 10.6151
R1270 B.n527 B.n92 10.6151
R1271 B.n527 B.n526 10.6151
R1272 B.n526 B.n525 10.6151
R1273 B.n525 B.n94 10.6151
R1274 B.n519 B.n94 10.6151
R1275 B.n519 B.n518 10.6151
R1276 B.n518 B.n517 10.6151
R1277 B.n517 B.n96 10.6151
R1278 B.n511 B.n96 10.6151
R1279 B.n511 B.n510 10.6151
R1280 B.n510 B.n509 10.6151
R1281 B.n509 B.n98 10.6151
R1282 B.n503 B.n98 10.6151
R1283 B.n467 B.t1 9.98378
R1284 B.n760 B.t0 9.98378
R1285 B.n320 B.n319 9.36635
R1286 B.n296 B.n171 9.36635
R1287 B.n628 B.n627 9.36635
R1288 B.n605 B.n72 9.36635
R1289 B.n772 B.n0 8.11757
R1290 B.n772 B.n1 8.11757
R1291 B.n442 B.t10 5.78029
R1292 B.n744 B.t3 5.78029
R1293 B.n319 B.n318 1.24928
R1294 B.n171 B.n167 1.24928
R1295 B.n627 B.n626 1.24928
R1296 B.n609 B.n72 1.24928
R1297 VN VN.t1 412.64
R1298 VN VN.t0 368.122
R1299 VDD2.n0 VDD2.t1 101.138
R1300 VDD2.n0 VDD2.t0 60.9089
R1301 VDD2 VDD2.n0 0.44231
C0 VP VDD1 3.29359f
C1 VDD1 VN 0.147929f
C2 VP VN 5.58958f
C3 VTAIL VDD1 6.1726f
C4 VTAIL VP 2.61075f
C5 VTAIL VN 2.59623f
C6 VDD2 VDD1 0.541302f
C7 VDD2 VP 0.285657f
C8 VDD2 VN 3.16018f
C9 VDD2 VTAIL 6.21233f
C10 VDD2 B 4.684463f
C11 VDD1 B 7.8503f
C12 VTAIL B 8.194579f
C13 VN B 10.522981f
C14 VP B 5.206395f
C15 VDD2.t1 B 3.47868f
C16 VDD2.t0 B 2.8807f
C17 VDD2.n0 B 2.96158f
C18 VN.t0 B 2.9247f
C19 VN.t1 B 3.22229f
C20 VDD1.t0 B 2.89036f
C21 VDD1.t1 B 3.51944f
C22 VTAIL.t3 B 2.76329f
C23 VTAIL.n0 B 1.66503f
C24 VTAIL.t1 B 2.76331f
C25 VTAIL.n1 B 1.68587f
C26 VTAIL.t2 B 2.76329f
C27 VTAIL.n2 B 1.58752f
C28 VTAIL.t0 B 2.76329f
C29 VTAIL.n3 B 1.52909f
C30 VP.t1 B 3.26317f
C31 VP.t0 B 2.96532f
C32 VP.n0 B 5.22876f
.ends

