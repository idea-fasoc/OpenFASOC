* NGSPICE file created from diff_pair_sample_0507.ext - technology: sky130A

.subckt diff_pair_sample_0507 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0 ps=0 w=4.68 l=1.38
X1 VTAIL.t7 VP.t0 VDD1.t1 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0.7722 ps=5.01 w=4.68 l=1.38
X2 VTAIL.t1 VN.t0 VDD2.t3 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0.7722 ps=5.01 w=4.68 l=1.38
X3 VDD2.t2 VN.t1 VTAIL.t2 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=0.7722 pd=5.01 as=1.8252 ps=10.14 w=4.68 l=1.38
X4 VDD1.t3 VP.t1 VTAIL.t6 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=0.7722 pd=5.01 as=1.8252 ps=10.14 w=4.68 l=1.38
X5 VDD2.t1 VN.t2 VTAIL.t0 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=0.7722 pd=5.01 as=1.8252 ps=10.14 w=4.68 l=1.38
X6 VTAIL.t5 VP.t2 VDD1.t2 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0.7722 ps=5.01 w=4.68 l=1.38
X7 VDD1.t0 VP.t3 VTAIL.t4 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=0.7722 pd=5.01 as=1.8252 ps=10.14 w=4.68 l=1.38
X8 B.t8 B.t6 B.t7 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0 ps=0 w=4.68 l=1.38
X9 B.t5 B.t3 B.t4 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0 ps=0 w=4.68 l=1.38
X10 VTAIL.t3 VN.t3 VDD2.t0 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0.7722 ps=5.01 w=4.68 l=1.38
X11 B.t2 B.t0 B.t1 w_n1996_n1904# sky130_fd_pr__pfet_01v8 ad=1.8252 pd=10.14 as=0 ps=0 w=4.68 l=1.38
R0 B.n288 B.n43 585
R1 B.n290 B.n289 585
R2 B.n291 B.n42 585
R3 B.n293 B.n292 585
R4 B.n294 B.n41 585
R5 B.n296 B.n295 585
R6 B.n297 B.n40 585
R7 B.n299 B.n298 585
R8 B.n300 B.n39 585
R9 B.n302 B.n301 585
R10 B.n303 B.n38 585
R11 B.n305 B.n304 585
R12 B.n306 B.n37 585
R13 B.n308 B.n307 585
R14 B.n309 B.n36 585
R15 B.n311 B.n310 585
R16 B.n312 B.n35 585
R17 B.n314 B.n313 585
R18 B.n315 B.n31 585
R19 B.n317 B.n316 585
R20 B.n318 B.n30 585
R21 B.n320 B.n319 585
R22 B.n321 B.n29 585
R23 B.n323 B.n322 585
R24 B.n324 B.n28 585
R25 B.n326 B.n325 585
R26 B.n327 B.n27 585
R27 B.n329 B.n328 585
R28 B.n330 B.n26 585
R29 B.n332 B.n331 585
R30 B.n334 B.n23 585
R31 B.n336 B.n335 585
R32 B.n337 B.n22 585
R33 B.n339 B.n338 585
R34 B.n340 B.n21 585
R35 B.n342 B.n341 585
R36 B.n343 B.n20 585
R37 B.n345 B.n344 585
R38 B.n346 B.n19 585
R39 B.n348 B.n347 585
R40 B.n349 B.n18 585
R41 B.n351 B.n350 585
R42 B.n352 B.n17 585
R43 B.n354 B.n353 585
R44 B.n355 B.n16 585
R45 B.n357 B.n356 585
R46 B.n358 B.n15 585
R47 B.n360 B.n359 585
R48 B.n361 B.n14 585
R49 B.n363 B.n362 585
R50 B.n287 B.n286 585
R51 B.n285 B.n44 585
R52 B.n284 B.n283 585
R53 B.n282 B.n45 585
R54 B.n281 B.n280 585
R55 B.n279 B.n46 585
R56 B.n278 B.n277 585
R57 B.n276 B.n47 585
R58 B.n275 B.n274 585
R59 B.n273 B.n48 585
R60 B.n272 B.n271 585
R61 B.n270 B.n49 585
R62 B.n269 B.n268 585
R63 B.n267 B.n50 585
R64 B.n266 B.n265 585
R65 B.n264 B.n51 585
R66 B.n263 B.n262 585
R67 B.n261 B.n52 585
R68 B.n260 B.n259 585
R69 B.n258 B.n53 585
R70 B.n257 B.n256 585
R71 B.n255 B.n54 585
R72 B.n254 B.n253 585
R73 B.n252 B.n55 585
R74 B.n251 B.n250 585
R75 B.n249 B.n56 585
R76 B.n248 B.n247 585
R77 B.n246 B.n57 585
R78 B.n245 B.n244 585
R79 B.n243 B.n58 585
R80 B.n242 B.n241 585
R81 B.n240 B.n59 585
R82 B.n239 B.n238 585
R83 B.n237 B.n60 585
R84 B.n236 B.n235 585
R85 B.n234 B.n61 585
R86 B.n233 B.n232 585
R87 B.n231 B.n62 585
R88 B.n230 B.n229 585
R89 B.n228 B.n63 585
R90 B.n227 B.n226 585
R91 B.n225 B.n64 585
R92 B.n224 B.n223 585
R93 B.n222 B.n65 585
R94 B.n221 B.n220 585
R95 B.n219 B.n66 585
R96 B.n218 B.n217 585
R97 B.n141 B.n96 585
R98 B.n143 B.n142 585
R99 B.n144 B.n95 585
R100 B.n146 B.n145 585
R101 B.n147 B.n94 585
R102 B.n149 B.n148 585
R103 B.n150 B.n93 585
R104 B.n152 B.n151 585
R105 B.n153 B.n92 585
R106 B.n155 B.n154 585
R107 B.n156 B.n91 585
R108 B.n158 B.n157 585
R109 B.n159 B.n90 585
R110 B.n161 B.n160 585
R111 B.n162 B.n89 585
R112 B.n164 B.n163 585
R113 B.n165 B.n88 585
R114 B.n167 B.n166 585
R115 B.n168 B.n87 585
R116 B.n170 B.n169 585
R117 B.n172 B.n84 585
R118 B.n174 B.n173 585
R119 B.n175 B.n83 585
R120 B.n177 B.n176 585
R121 B.n178 B.n82 585
R122 B.n180 B.n179 585
R123 B.n181 B.n81 585
R124 B.n183 B.n182 585
R125 B.n184 B.n80 585
R126 B.n186 B.n185 585
R127 B.n188 B.n187 585
R128 B.n189 B.n76 585
R129 B.n191 B.n190 585
R130 B.n192 B.n75 585
R131 B.n194 B.n193 585
R132 B.n195 B.n74 585
R133 B.n197 B.n196 585
R134 B.n198 B.n73 585
R135 B.n200 B.n199 585
R136 B.n201 B.n72 585
R137 B.n203 B.n202 585
R138 B.n204 B.n71 585
R139 B.n206 B.n205 585
R140 B.n207 B.n70 585
R141 B.n209 B.n208 585
R142 B.n210 B.n69 585
R143 B.n212 B.n211 585
R144 B.n213 B.n68 585
R145 B.n215 B.n214 585
R146 B.n216 B.n67 585
R147 B.n140 B.n139 585
R148 B.n138 B.n97 585
R149 B.n137 B.n136 585
R150 B.n135 B.n98 585
R151 B.n134 B.n133 585
R152 B.n132 B.n99 585
R153 B.n131 B.n130 585
R154 B.n129 B.n100 585
R155 B.n128 B.n127 585
R156 B.n126 B.n101 585
R157 B.n125 B.n124 585
R158 B.n123 B.n102 585
R159 B.n122 B.n121 585
R160 B.n120 B.n103 585
R161 B.n119 B.n118 585
R162 B.n117 B.n104 585
R163 B.n116 B.n115 585
R164 B.n114 B.n105 585
R165 B.n113 B.n112 585
R166 B.n111 B.n106 585
R167 B.n110 B.n109 585
R168 B.n108 B.n107 585
R169 B.n2 B.n0 585
R170 B.n397 B.n1 585
R171 B.n396 B.n395 585
R172 B.n394 B.n3 585
R173 B.n393 B.n392 585
R174 B.n391 B.n4 585
R175 B.n390 B.n389 585
R176 B.n388 B.n5 585
R177 B.n387 B.n386 585
R178 B.n385 B.n6 585
R179 B.n384 B.n383 585
R180 B.n382 B.n7 585
R181 B.n381 B.n380 585
R182 B.n379 B.n8 585
R183 B.n378 B.n377 585
R184 B.n376 B.n9 585
R185 B.n375 B.n374 585
R186 B.n373 B.n10 585
R187 B.n372 B.n371 585
R188 B.n370 B.n11 585
R189 B.n369 B.n368 585
R190 B.n367 B.n12 585
R191 B.n366 B.n365 585
R192 B.n364 B.n13 585
R193 B.n399 B.n398 585
R194 B.n139 B.n96 511.721
R195 B.n362 B.n13 511.721
R196 B.n217 B.n216 511.721
R197 B.n288 B.n287 511.721
R198 B.n77 B.t6 286.693
R199 B.n85 B.t9 286.693
R200 B.n24 B.t3 286.693
R201 B.n32 B.t0 286.693
R202 B.n77 B.t8 279.06
R203 B.n32 B.t1 279.06
R204 B.n85 B.t11 279.06
R205 B.n24 B.t4 279.06
R206 B.n78 B.t7 245.897
R207 B.n33 B.t2 245.897
R208 B.n86 B.t10 245.897
R209 B.n25 B.t5 245.897
R210 B.n139 B.n138 163.367
R211 B.n138 B.n137 163.367
R212 B.n137 B.n98 163.367
R213 B.n133 B.n98 163.367
R214 B.n133 B.n132 163.367
R215 B.n132 B.n131 163.367
R216 B.n131 B.n100 163.367
R217 B.n127 B.n100 163.367
R218 B.n127 B.n126 163.367
R219 B.n126 B.n125 163.367
R220 B.n125 B.n102 163.367
R221 B.n121 B.n102 163.367
R222 B.n121 B.n120 163.367
R223 B.n120 B.n119 163.367
R224 B.n119 B.n104 163.367
R225 B.n115 B.n104 163.367
R226 B.n115 B.n114 163.367
R227 B.n114 B.n113 163.367
R228 B.n113 B.n106 163.367
R229 B.n109 B.n106 163.367
R230 B.n109 B.n108 163.367
R231 B.n108 B.n2 163.367
R232 B.n398 B.n2 163.367
R233 B.n398 B.n397 163.367
R234 B.n397 B.n396 163.367
R235 B.n396 B.n3 163.367
R236 B.n392 B.n3 163.367
R237 B.n392 B.n391 163.367
R238 B.n391 B.n390 163.367
R239 B.n390 B.n5 163.367
R240 B.n386 B.n5 163.367
R241 B.n386 B.n385 163.367
R242 B.n385 B.n384 163.367
R243 B.n384 B.n7 163.367
R244 B.n380 B.n7 163.367
R245 B.n380 B.n379 163.367
R246 B.n379 B.n378 163.367
R247 B.n378 B.n9 163.367
R248 B.n374 B.n9 163.367
R249 B.n374 B.n373 163.367
R250 B.n373 B.n372 163.367
R251 B.n372 B.n11 163.367
R252 B.n368 B.n11 163.367
R253 B.n368 B.n367 163.367
R254 B.n367 B.n366 163.367
R255 B.n366 B.n13 163.367
R256 B.n143 B.n96 163.367
R257 B.n144 B.n143 163.367
R258 B.n145 B.n144 163.367
R259 B.n145 B.n94 163.367
R260 B.n149 B.n94 163.367
R261 B.n150 B.n149 163.367
R262 B.n151 B.n150 163.367
R263 B.n151 B.n92 163.367
R264 B.n155 B.n92 163.367
R265 B.n156 B.n155 163.367
R266 B.n157 B.n156 163.367
R267 B.n157 B.n90 163.367
R268 B.n161 B.n90 163.367
R269 B.n162 B.n161 163.367
R270 B.n163 B.n162 163.367
R271 B.n163 B.n88 163.367
R272 B.n167 B.n88 163.367
R273 B.n168 B.n167 163.367
R274 B.n169 B.n168 163.367
R275 B.n169 B.n84 163.367
R276 B.n174 B.n84 163.367
R277 B.n175 B.n174 163.367
R278 B.n176 B.n175 163.367
R279 B.n176 B.n82 163.367
R280 B.n180 B.n82 163.367
R281 B.n181 B.n180 163.367
R282 B.n182 B.n181 163.367
R283 B.n182 B.n80 163.367
R284 B.n186 B.n80 163.367
R285 B.n187 B.n186 163.367
R286 B.n187 B.n76 163.367
R287 B.n191 B.n76 163.367
R288 B.n192 B.n191 163.367
R289 B.n193 B.n192 163.367
R290 B.n193 B.n74 163.367
R291 B.n197 B.n74 163.367
R292 B.n198 B.n197 163.367
R293 B.n199 B.n198 163.367
R294 B.n199 B.n72 163.367
R295 B.n203 B.n72 163.367
R296 B.n204 B.n203 163.367
R297 B.n205 B.n204 163.367
R298 B.n205 B.n70 163.367
R299 B.n209 B.n70 163.367
R300 B.n210 B.n209 163.367
R301 B.n211 B.n210 163.367
R302 B.n211 B.n68 163.367
R303 B.n215 B.n68 163.367
R304 B.n216 B.n215 163.367
R305 B.n217 B.n66 163.367
R306 B.n221 B.n66 163.367
R307 B.n222 B.n221 163.367
R308 B.n223 B.n222 163.367
R309 B.n223 B.n64 163.367
R310 B.n227 B.n64 163.367
R311 B.n228 B.n227 163.367
R312 B.n229 B.n228 163.367
R313 B.n229 B.n62 163.367
R314 B.n233 B.n62 163.367
R315 B.n234 B.n233 163.367
R316 B.n235 B.n234 163.367
R317 B.n235 B.n60 163.367
R318 B.n239 B.n60 163.367
R319 B.n240 B.n239 163.367
R320 B.n241 B.n240 163.367
R321 B.n241 B.n58 163.367
R322 B.n245 B.n58 163.367
R323 B.n246 B.n245 163.367
R324 B.n247 B.n246 163.367
R325 B.n247 B.n56 163.367
R326 B.n251 B.n56 163.367
R327 B.n252 B.n251 163.367
R328 B.n253 B.n252 163.367
R329 B.n253 B.n54 163.367
R330 B.n257 B.n54 163.367
R331 B.n258 B.n257 163.367
R332 B.n259 B.n258 163.367
R333 B.n259 B.n52 163.367
R334 B.n263 B.n52 163.367
R335 B.n264 B.n263 163.367
R336 B.n265 B.n264 163.367
R337 B.n265 B.n50 163.367
R338 B.n269 B.n50 163.367
R339 B.n270 B.n269 163.367
R340 B.n271 B.n270 163.367
R341 B.n271 B.n48 163.367
R342 B.n275 B.n48 163.367
R343 B.n276 B.n275 163.367
R344 B.n277 B.n276 163.367
R345 B.n277 B.n46 163.367
R346 B.n281 B.n46 163.367
R347 B.n282 B.n281 163.367
R348 B.n283 B.n282 163.367
R349 B.n283 B.n44 163.367
R350 B.n287 B.n44 163.367
R351 B.n362 B.n361 163.367
R352 B.n361 B.n360 163.367
R353 B.n360 B.n15 163.367
R354 B.n356 B.n15 163.367
R355 B.n356 B.n355 163.367
R356 B.n355 B.n354 163.367
R357 B.n354 B.n17 163.367
R358 B.n350 B.n17 163.367
R359 B.n350 B.n349 163.367
R360 B.n349 B.n348 163.367
R361 B.n348 B.n19 163.367
R362 B.n344 B.n19 163.367
R363 B.n344 B.n343 163.367
R364 B.n343 B.n342 163.367
R365 B.n342 B.n21 163.367
R366 B.n338 B.n21 163.367
R367 B.n338 B.n337 163.367
R368 B.n337 B.n336 163.367
R369 B.n336 B.n23 163.367
R370 B.n331 B.n23 163.367
R371 B.n331 B.n330 163.367
R372 B.n330 B.n329 163.367
R373 B.n329 B.n27 163.367
R374 B.n325 B.n27 163.367
R375 B.n325 B.n324 163.367
R376 B.n324 B.n323 163.367
R377 B.n323 B.n29 163.367
R378 B.n319 B.n29 163.367
R379 B.n319 B.n318 163.367
R380 B.n318 B.n317 163.367
R381 B.n317 B.n31 163.367
R382 B.n313 B.n31 163.367
R383 B.n313 B.n312 163.367
R384 B.n312 B.n311 163.367
R385 B.n311 B.n36 163.367
R386 B.n307 B.n36 163.367
R387 B.n307 B.n306 163.367
R388 B.n306 B.n305 163.367
R389 B.n305 B.n38 163.367
R390 B.n301 B.n38 163.367
R391 B.n301 B.n300 163.367
R392 B.n300 B.n299 163.367
R393 B.n299 B.n40 163.367
R394 B.n295 B.n40 163.367
R395 B.n295 B.n294 163.367
R396 B.n294 B.n293 163.367
R397 B.n293 B.n42 163.367
R398 B.n289 B.n42 163.367
R399 B.n289 B.n288 163.367
R400 B.n79 B.n78 59.5399
R401 B.n171 B.n86 59.5399
R402 B.n333 B.n25 59.5399
R403 B.n34 B.n33 59.5399
R404 B.n364 B.n363 33.2493
R405 B.n286 B.n43 33.2493
R406 B.n218 B.n67 33.2493
R407 B.n141 B.n140 33.2493
R408 B.n78 B.n77 33.1641
R409 B.n86 B.n85 33.1641
R410 B.n25 B.n24 33.1641
R411 B.n33 B.n32 33.1641
R412 B B.n399 18.0485
R413 B.n363 B.n14 10.6151
R414 B.n359 B.n14 10.6151
R415 B.n359 B.n358 10.6151
R416 B.n358 B.n357 10.6151
R417 B.n357 B.n16 10.6151
R418 B.n353 B.n16 10.6151
R419 B.n353 B.n352 10.6151
R420 B.n352 B.n351 10.6151
R421 B.n351 B.n18 10.6151
R422 B.n347 B.n18 10.6151
R423 B.n347 B.n346 10.6151
R424 B.n346 B.n345 10.6151
R425 B.n345 B.n20 10.6151
R426 B.n341 B.n20 10.6151
R427 B.n341 B.n340 10.6151
R428 B.n340 B.n339 10.6151
R429 B.n339 B.n22 10.6151
R430 B.n335 B.n22 10.6151
R431 B.n335 B.n334 10.6151
R432 B.n332 B.n26 10.6151
R433 B.n328 B.n26 10.6151
R434 B.n328 B.n327 10.6151
R435 B.n327 B.n326 10.6151
R436 B.n326 B.n28 10.6151
R437 B.n322 B.n28 10.6151
R438 B.n322 B.n321 10.6151
R439 B.n321 B.n320 10.6151
R440 B.n320 B.n30 10.6151
R441 B.n316 B.n315 10.6151
R442 B.n315 B.n314 10.6151
R443 B.n314 B.n35 10.6151
R444 B.n310 B.n35 10.6151
R445 B.n310 B.n309 10.6151
R446 B.n309 B.n308 10.6151
R447 B.n308 B.n37 10.6151
R448 B.n304 B.n37 10.6151
R449 B.n304 B.n303 10.6151
R450 B.n303 B.n302 10.6151
R451 B.n302 B.n39 10.6151
R452 B.n298 B.n39 10.6151
R453 B.n298 B.n297 10.6151
R454 B.n297 B.n296 10.6151
R455 B.n296 B.n41 10.6151
R456 B.n292 B.n41 10.6151
R457 B.n292 B.n291 10.6151
R458 B.n291 B.n290 10.6151
R459 B.n290 B.n43 10.6151
R460 B.n219 B.n218 10.6151
R461 B.n220 B.n219 10.6151
R462 B.n220 B.n65 10.6151
R463 B.n224 B.n65 10.6151
R464 B.n225 B.n224 10.6151
R465 B.n226 B.n225 10.6151
R466 B.n226 B.n63 10.6151
R467 B.n230 B.n63 10.6151
R468 B.n231 B.n230 10.6151
R469 B.n232 B.n231 10.6151
R470 B.n232 B.n61 10.6151
R471 B.n236 B.n61 10.6151
R472 B.n237 B.n236 10.6151
R473 B.n238 B.n237 10.6151
R474 B.n238 B.n59 10.6151
R475 B.n242 B.n59 10.6151
R476 B.n243 B.n242 10.6151
R477 B.n244 B.n243 10.6151
R478 B.n244 B.n57 10.6151
R479 B.n248 B.n57 10.6151
R480 B.n249 B.n248 10.6151
R481 B.n250 B.n249 10.6151
R482 B.n250 B.n55 10.6151
R483 B.n254 B.n55 10.6151
R484 B.n255 B.n254 10.6151
R485 B.n256 B.n255 10.6151
R486 B.n256 B.n53 10.6151
R487 B.n260 B.n53 10.6151
R488 B.n261 B.n260 10.6151
R489 B.n262 B.n261 10.6151
R490 B.n262 B.n51 10.6151
R491 B.n266 B.n51 10.6151
R492 B.n267 B.n266 10.6151
R493 B.n268 B.n267 10.6151
R494 B.n268 B.n49 10.6151
R495 B.n272 B.n49 10.6151
R496 B.n273 B.n272 10.6151
R497 B.n274 B.n273 10.6151
R498 B.n274 B.n47 10.6151
R499 B.n278 B.n47 10.6151
R500 B.n279 B.n278 10.6151
R501 B.n280 B.n279 10.6151
R502 B.n280 B.n45 10.6151
R503 B.n284 B.n45 10.6151
R504 B.n285 B.n284 10.6151
R505 B.n286 B.n285 10.6151
R506 B.n142 B.n141 10.6151
R507 B.n142 B.n95 10.6151
R508 B.n146 B.n95 10.6151
R509 B.n147 B.n146 10.6151
R510 B.n148 B.n147 10.6151
R511 B.n148 B.n93 10.6151
R512 B.n152 B.n93 10.6151
R513 B.n153 B.n152 10.6151
R514 B.n154 B.n153 10.6151
R515 B.n154 B.n91 10.6151
R516 B.n158 B.n91 10.6151
R517 B.n159 B.n158 10.6151
R518 B.n160 B.n159 10.6151
R519 B.n160 B.n89 10.6151
R520 B.n164 B.n89 10.6151
R521 B.n165 B.n164 10.6151
R522 B.n166 B.n165 10.6151
R523 B.n166 B.n87 10.6151
R524 B.n170 B.n87 10.6151
R525 B.n173 B.n172 10.6151
R526 B.n173 B.n83 10.6151
R527 B.n177 B.n83 10.6151
R528 B.n178 B.n177 10.6151
R529 B.n179 B.n178 10.6151
R530 B.n179 B.n81 10.6151
R531 B.n183 B.n81 10.6151
R532 B.n184 B.n183 10.6151
R533 B.n185 B.n184 10.6151
R534 B.n189 B.n188 10.6151
R535 B.n190 B.n189 10.6151
R536 B.n190 B.n75 10.6151
R537 B.n194 B.n75 10.6151
R538 B.n195 B.n194 10.6151
R539 B.n196 B.n195 10.6151
R540 B.n196 B.n73 10.6151
R541 B.n200 B.n73 10.6151
R542 B.n201 B.n200 10.6151
R543 B.n202 B.n201 10.6151
R544 B.n202 B.n71 10.6151
R545 B.n206 B.n71 10.6151
R546 B.n207 B.n206 10.6151
R547 B.n208 B.n207 10.6151
R548 B.n208 B.n69 10.6151
R549 B.n212 B.n69 10.6151
R550 B.n213 B.n212 10.6151
R551 B.n214 B.n213 10.6151
R552 B.n214 B.n67 10.6151
R553 B.n140 B.n97 10.6151
R554 B.n136 B.n97 10.6151
R555 B.n136 B.n135 10.6151
R556 B.n135 B.n134 10.6151
R557 B.n134 B.n99 10.6151
R558 B.n130 B.n99 10.6151
R559 B.n130 B.n129 10.6151
R560 B.n129 B.n128 10.6151
R561 B.n128 B.n101 10.6151
R562 B.n124 B.n101 10.6151
R563 B.n124 B.n123 10.6151
R564 B.n123 B.n122 10.6151
R565 B.n122 B.n103 10.6151
R566 B.n118 B.n103 10.6151
R567 B.n118 B.n117 10.6151
R568 B.n117 B.n116 10.6151
R569 B.n116 B.n105 10.6151
R570 B.n112 B.n105 10.6151
R571 B.n112 B.n111 10.6151
R572 B.n111 B.n110 10.6151
R573 B.n110 B.n107 10.6151
R574 B.n107 B.n0 10.6151
R575 B.n395 B.n1 10.6151
R576 B.n395 B.n394 10.6151
R577 B.n394 B.n393 10.6151
R578 B.n393 B.n4 10.6151
R579 B.n389 B.n4 10.6151
R580 B.n389 B.n388 10.6151
R581 B.n388 B.n387 10.6151
R582 B.n387 B.n6 10.6151
R583 B.n383 B.n6 10.6151
R584 B.n383 B.n382 10.6151
R585 B.n382 B.n381 10.6151
R586 B.n381 B.n8 10.6151
R587 B.n377 B.n8 10.6151
R588 B.n377 B.n376 10.6151
R589 B.n376 B.n375 10.6151
R590 B.n375 B.n10 10.6151
R591 B.n371 B.n10 10.6151
R592 B.n371 B.n370 10.6151
R593 B.n370 B.n369 10.6151
R594 B.n369 B.n12 10.6151
R595 B.n365 B.n12 10.6151
R596 B.n365 B.n364 10.6151
R597 B.n334 B.n333 9.36635
R598 B.n316 B.n34 9.36635
R599 B.n171 B.n170 9.36635
R600 B.n188 B.n79 9.36635
R601 B.n399 B.n0 2.81026
R602 B.n399 B.n1 2.81026
R603 B.n333 B.n332 1.24928
R604 B.n34 B.n30 1.24928
R605 B.n172 B.n171 1.24928
R606 B.n185 B.n79 1.24928
R607 VP.n4 VP.n3 168.433
R608 VP.n10 VP.n9 168.433
R609 VP.n8 VP.n0 161.3
R610 VP.n7 VP.n6 161.3
R611 VP.n5 VP.n1 161.3
R612 VP.n2 VP.t0 120.371
R613 VP.n2 VP.t3 120.138
R614 VP.n3 VP.t2 81.7309
R615 VP.n9 VP.t1 81.7309
R616 VP.n4 VP.n2 54.5735
R617 VP.n7 VP.n1 40.577
R618 VP.n8 VP.n7 40.577
R619 VP.n3 VP.n1 17.4607
R620 VP.n9 VP.n8 17.4607
R621 VP.n5 VP.n4 0.189894
R622 VP.n6 VP.n5 0.189894
R623 VP.n6 VP.n0 0.189894
R624 VP.n10 VP.n0 0.189894
R625 VP VP.n10 0.0516364
R626 VDD1 VDD1.n1 139.103
R627 VDD1 VDD1.n0 106.466
R628 VDD1.n0 VDD1.t1 6.94601
R629 VDD1.n0 VDD1.t0 6.94601
R630 VDD1.n1 VDD1.t2 6.94601
R631 VDD1.n1 VDD1.t3 6.94601
R632 VTAIL.n186 VTAIL.n168 756.745
R633 VTAIL.n18 VTAIL.n0 756.745
R634 VTAIL.n42 VTAIL.n24 756.745
R635 VTAIL.n66 VTAIL.n48 756.745
R636 VTAIL.n162 VTAIL.n144 756.745
R637 VTAIL.n138 VTAIL.n120 756.745
R638 VTAIL.n114 VTAIL.n96 756.745
R639 VTAIL.n90 VTAIL.n72 756.745
R640 VTAIL.n177 VTAIL.n176 585
R641 VTAIL.n179 VTAIL.n178 585
R642 VTAIL.n172 VTAIL.n171 585
R643 VTAIL.n185 VTAIL.n184 585
R644 VTAIL.n187 VTAIL.n186 585
R645 VTAIL.n9 VTAIL.n8 585
R646 VTAIL.n11 VTAIL.n10 585
R647 VTAIL.n4 VTAIL.n3 585
R648 VTAIL.n17 VTAIL.n16 585
R649 VTAIL.n19 VTAIL.n18 585
R650 VTAIL.n33 VTAIL.n32 585
R651 VTAIL.n35 VTAIL.n34 585
R652 VTAIL.n28 VTAIL.n27 585
R653 VTAIL.n41 VTAIL.n40 585
R654 VTAIL.n43 VTAIL.n42 585
R655 VTAIL.n57 VTAIL.n56 585
R656 VTAIL.n59 VTAIL.n58 585
R657 VTAIL.n52 VTAIL.n51 585
R658 VTAIL.n65 VTAIL.n64 585
R659 VTAIL.n67 VTAIL.n66 585
R660 VTAIL.n163 VTAIL.n162 585
R661 VTAIL.n161 VTAIL.n160 585
R662 VTAIL.n148 VTAIL.n147 585
R663 VTAIL.n155 VTAIL.n154 585
R664 VTAIL.n153 VTAIL.n152 585
R665 VTAIL.n139 VTAIL.n138 585
R666 VTAIL.n137 VTAIL.n136 585
R667 VTAIL.n124 VTAIL.n123 585
R668 VTAIL.n131 VTAIL.n130 585
R669 VTAIL.n129 VTAIL.n128 585
R670 VTAIL.n115 VTAIL.n114 585
R671 VTAIL.n113 VTAIL.n112 585
R672 VTAIL.n100 VTAIL.n99 585
R673 VTAIL.n107 VTAIL.n106 585
R674 VTAIL.n105 VTAIL.n104 585
R675 VTAIL.n91 VTAIL.n90 585
R676 VTAIL.n89 VTAIL.n88 585
R677 VTAIL.n76 VTAIL.n75 585
R678 VTAIL.n83 VTAIL.n82 585
R679 VTAIL.n81 VTAIL.n80 585
R680 VTAIL.n175 VTAIL.t0 328.587
R681 VTAIL.n7 VTAIL.t1 328.587
R682 VTAIL.n31 VTAIL.t6 328.587
R683 VTAIL.n55 VTAIL.t5 328.587
R684 VTAIL.n151 VTAIL.t4 328.587
R685 VTAIL.n127 VTAIL.t7 328.587
R686 VTAIL.n103 VTAIL.t2 328.587
R687 VTAIL.n79 VTAIL.t3 328.587
R688 VTAIL.n178 VTAIL.n177 171.744
R689 VTAIL.n178 VTAIL.n171 171.744
R690 VTAIL.n185 VTAIL.n171 171.744
R691 VTAIL.n186 VTAIL.n185 171.744
R692 VTAIL.n10 VTAIL.n9 171.744
R693 VTAIL.n10 VTAIL.n3 171.744
R694 VTAIL.n17 VTAIL.n3 171.744
R695 VTAIL.n18 VTAIL.n17 171.744
R696 VTAIL.n34 VTAIL.n33 171.744
R697 VTAIL.n34 VTAIL.n27 171.744
R698 VTAIL.n41 VTAIL.n27 171.744
R699 VTAIL.n42 VTAIL.n41 171.744
R700 VTAIL.n58 VTAIL.n57 171.744
R701 VTAIL.n58 VTAIL.n51 171.744
R702 VTAIL.n65 VTAIL.n51 171.744
R703 VTAIL.n66 VTAIL.n65 171.744
R704 VTAIL.n162 VTAIL.n161 171.744
R705 VTAIL.n161 VTAIL.n147 171.744
R706 VTAIL.n154 VTAIL.n147 171.744
R707 VTAIL.n154 VTAIL.n153 171.744
R708 VTAIL.n138 VTAIL.n137 171.744
R709 VTAIL.n137 VTAIL.n123 171.744
R710 VTAIL.n130 VTAIL.n123 171.744
R711 VTAIL.n130 VTAIL.n129 171.744
R712 VTAIL.n114 VTAIL.n113 171.744
R713 VTAIL.n113 VTAIL.n99 171.744
R714 VTAIL.n106 VTAIL.n99 171.744
R715 VTAIL.n106 VTAIL.n105 171.744
R716 VTAIL.n90 VTAIL.n89 171.744
R717 VTAIL.n89 VTAIL.n75 171.744
R718 VTAIL.n82 VTAIL.n75 171.744
R719 VTAIL.n82 VTAIL.n81 171.744
R720 VTAIL.n177 VTAIL.t0 85.8723
R721 VTAIL.n9 VTAIL.t1 85.8723
R722 VTAIL.n33 VTAIL.t6 85.8723
R723 VTAIL.n57 VTAIL.t5 85.8723
R724 VTAIL.n153 VTAIL.t4 85.8723
R725 VTAIL.n129 VTAIL.t7 85.8723
R726 VTAIL.n105 VTAIL.t2 85.8723
R727 VTAIL.n81 VTAIL.t3 85.8723
R728 VTAIL.n191 VTAIL.n190 34.5126
R729 VTAIL.n23 VTAIL.n22 34.5126
R730 VTAIL.n47 VTAIL.n46 34.5126
R731 VTAIL.n71 VTAIL.n70 34.5126
R732 VTAIL.n167 VTAIL.n166 34.5126
R733 VTAIL.n143 VTAIL.n142 34.5126
R734 VTAIL.n119 VTAIL.n118 34.5126
R735 VTAIL.n95 VTAIL.n94 34.5126
R736 VTAIL.n191 VTAIL.n167 17.8755
R737 VTAIL.n95 VTAIL.n71 17.8755
R738 VTAIL.n176 VTAIL.n175 16.3651
R739 VTAIL.n8 VTAIL.n7 16.3651
R740 VTAIL.n32 VTAIL.n31 16.3651
R741 VTAIL.n56 VTAIL.n55 16.3651
R742 VTAIL.n152 VTAIL.n151 16.3651
R743 VTAIL.n128 VTAIL.n127 16.3651
R744 VTAIL.n104 VTAIL.n103 16.3651
R745 VTAIL.n80 VTAIL.n79 16.3651
R746 VTAIL.n179 VTAIL.n174 12.8005
R747 VTAIL.n11 VTAIL.n6 12.8005
R748 VTAIL.n35 VTAIL.n30 12.8005
R749 VTAIL.n59 VTAIL.n54 12.8005
R750 VTAIL.n155 VTAIL.n150 12.8005
R751 VTAIL.n131 VTAIL.n126 12.8005
R752 VTAIL.n107 VTAIL.n102 12.8005
R753 VTAIL.n83 VTAIL.n78 12.8005
R754 VTAIL.n180 VTAIL.n172 12.0247
R755 VTAIL.n12 VTAIL.n4 12.0247
R756 VTAIL.n36 VTAIL.n28 12.0247
R757 VTAIL.n60 VTAIL.n52 12.0247
R758 VTAIL.n156 VTAIL.n148 12.0247
R759 VTAIL.n132 VTAIL.n124 12.0247
R760 VTAIL.n108 VTAIL.n100 12.0247
R761 VTAIL.n84 VTAIL.n76 12.0247
R762 VTAIL.n184 VTAIL.n183 11.249
R763 VTAIL.n16 VTAIL.n15 11.249
R764 VTAIL.n40 VTAIL.n39 11.249
R765 VTAIL.n64 VTAIL.n63 11.249
R766 VTAIL.n160 VTAIL.n159 11.249
R767 VTAIL.n136 VTAIL.n135 11.249
R768 VTAIL.n112 VTAIL.n111 11.249
R769 VTAIL.n88 VTAIL.n87 11.249
R770 VTAIL.n187 VTAIL.n170 10.4732
R771 VTAIL.n19 VTAIL.n2 10.4732
R772 VTAIL.n43 VTAIL.n26 10.4732
R773 VTAIL.n67 VTAIL.n50 10.4732
R774 VTAIL.n163 VTAIL.n146 10.4732
R775 VTAIL.n139 VTAIL.n122 10.4732
R776 VTAIL.n115 VTAIL.n98 10.4732
R777 VTAIL.n91 VTAIL.n74 10.4732
R778 VTAIL.n188 VTAIL.n168 9.69747
R779 VTAIL.n20 VTAIL.n0 9.69747
R780 VTAIL.n44 VTAIL.n24 9.69747
R781 VTAIL.n68 VTAIL.n48 9.69747
R782 VTAIL.n164 VTAIL.n144 9.69747
R783 VTAIL.n140 VTAIL.n120 9.69747
R784 VTAIL.n116 VTAIL.n96 9.69747
R785 VTAIL.n92 VTAIL.n72 9.69747
R786 VTAIL.n190 VTAIL.n189 9.45567
R787 VTAIL.n22 VTAIL.n21 9.45567
R788 VTAIL.n46 VTAIL.n45 9.45567
R789 VTAIL.n70 VTAIL.n69 9.45567
R790 VTAIL.n166 VTAIL.n165 9.45567
R791 VTAIL.n142 VTAIL.n141 9.45567
R792 VTAIL.n118 VTAIL.n117 9.45567
R793 VTAIL.n94 VTAIL.n93 9.45567
R794 VTAIL.n189 VTAIL.n188 9.3005
R795 VTAIL.n170 VTAIL.n169 9.3005
R796 VTAIL.n183 VTAIL.n182 9.3005
R797 VTAIL.n181 VTAIL.n180 9.3005
R798 VTAIL.n174 VTAIL.n173 9.3005
R799 VTAIL.n21 VTAIL.n20 9.3005
R800 VTAIL.n2 VTAIL.n1 9.3005
R801 VTAIL.n15 VTAIL.n14 9.3005
R802 VTAIL.n13 VTAIL.n12 9.3005
R803 VTAIL.n6 VTAIL.n5 9.3005
R804 VTAIL.n45 VTAIL.n44 9.3005
R805 VTAIL.n26 VTAIL.n25 9.3005
R806 VTAIL.n39 VTAIL.n38 9.3005
R807 VTAIL.n37 VTAIL.n36 9.3005
R808 VTAIL.n30 VTAIL.n29 9.3005
R809 VTAIL.n69 VTAIL.n68 9.3005
R810 VTAIL.n50 VTAIL.n49 9.3005
R811 VTAIL.n63 VTAIL.n62 9.3005
R812 VTAIL.n61 VTAIL.n60 9.3005
R813 VTAIL.n54 VTAIL.n53 9.3005
R814 VTAIL.n165 VTAIL.n164 9.3005
R815 VTAIL.n146 VTAIL.n145 9.3005
R816 VTAIL.n159 VTAIL.n158 9.3005
R817 VTAIL.n157 VTAIL.n156 9.3005
R818 VTAIL.n150 VTAIL.n149 9.3005
R819 VTAIL.n141 VTAIL.n140 9.3005
R820 VTAIL.n122 VTAIL.n121 9.3005
R821 VTAIL.n135 VTAIL.n134 9.3005
R822 VTAIL.n133 VTAIL.n132 9.3005
R823 VTAIL.n126 VTAIL.n125 9.3005
R824 VTAIL.n117 VTAIL.n116 9.3005
R825 VTAIL.n98 VTAIL.n97 9.3005
R826 VTAIL.n111 VTAIL.n110 9.3005
R827 VTAIL.n109 VTAIL.n108 9.3005
R828 VTAIL.n102 VTAIL.n101 9.3005
R829 VTAIL.n93 VTAIL.n92 9.3005
R830 VTAIL.n74 VTAIL.n73 9.3005
R831 VTAIL.n87 VTAIL.n86 9.3005
R832 VTAIL.n85 VTAIL.n84 9.3005
R833 VTAIL.n78 VTAIL.n77 9.3005
R834 VTAIL.n190 VTAIL.n168 4.26717
R835 VTAIL.n22 VTAIL.n0 4.26717
R836 VTAIL.n46 VTAIL.n24 4.26717
R837 VTAIL.n70 VTAIL.n48 4.26717
R838 VTAIL.n166 VTAIL.n144 4.26717
R839 VTAIL.n142 VTAIL.n120 4.26717
R840 VTAIL.n118 VTAIL.n96 4.26717
R841 VTAIL.n94 VTAIL.n72 4.26717
R842 VTAIL.n175 VTAIL.n173 3.73474
R843 VTAIL.n7 VTAIL.n5 3.73474
R844 VTAIL.n31 VTAIL.n29 3.73474
R845 VTAIL.n55 VTAIL.n53 3.73474
R846 VTAIL.n151 VTAIL.n149 3.73474
R847 VTAIL.n127 VTAIL.n125 3.73474
R848 VTAIL.n103 VTAIL.n101 3.73474
R849 VTAIL.n79 VTAIL.n77 3.73474
R850 VTAIL.n188 VTAIL.n187 3.49141
R851 VTAIL.n20 VTAIL.n19 3.49141
R852 VTAIL.n44 VTAIL.n43 3.49141
R853 VTAIL.n68 VTAIL.n67 3.49141
R854 VTAIL.n164 VTAIL.n163 3.49141
R855 VTAIL.n140 VTAIL.n139 3.49141
R856 VTAIL.n116 VTAIL.n115 3.49141
R857 VTAIL.n92 VTAIL.n91 3.49141
R858 VTAIL.n184 VTAIL.n170 2.71565
R859 VTAIL.n16 VTAIL.n2 2.71565
R860 VTAIL.n40 VTAIL.n26 2.71565
R861 VTAIL.n64 VTAIL.n50 2.71565
R862 VTAIL.n160 VTAIL.n146 2.71565
R863 VTAIL.n136 VTAIL.n122 2.71565
R864 VTAIL.n112 VTAIL.n98 2.71565
R865 VTAIL.n88 VTAIL.n74 2.71565
R866 VTAIL.n183 VTAIL.n172 1.93989
R867 VTAIL.n15 VTAIL.n4 1.93989
R868 VTAIL.n39 VTAIL.n28 1.93989
R869 VTAIL.n63 VTAIL.n52 1.93989
R870 VTAIL.n159 VTAIL.n148 1.93989
R871 VTAIL.n135 VTAIL.n124 1.93989
R872 VTAIL.n111 VTAIL.n100 1.93989
R873 VTAIL.n87 VTAIL.n76 1.93989
R874 VTAIL.n119 VTAIL.n95 1.47464
R875 VTAIL.n167 VTAIL.n143 1.47464
R876 VTAIL.n71 VTAIL.n47 1.47464
R877 VTAIL.n180 VTAIL.n179 1.16414
R878 VTAIL.n12 VTAIL.n11 1.16414
R879 VTAIL.n36 VTAIL.n35 1.16414
R880 VTAIL.n60 VTAIL.n59 1.16414
R881 VTAIL.n156 VTAIL.n155 1.16414
R882 VTAIL.n132 VTAIL.n131 1.16414
R883 VTAIL.n108 VTAIL.n107 1.16414
R884 VTAIL.n84 VTAIL.n83 1.16414
R885 VTAIL VTAIL.n23 0.795759
R886 VTAIL VTAIL.n191 0.679379
R887 VTAIL.n143 VTAIL.n119 0.470328
R888 VTAIL.n47 VTAIL.n23 0.470328
R889 VTAIL.n176 VTAIL.n174 0.388379
R890 VTAIL.n8 VTAIL.n6 0.388379
R891 VTAIL.n32 VTAIL.n30 0.388379
R892 VTAIL.n56 VTAIL.n54 0.388379
R893 VTAIL.n152 VTAIL.n150 0.388379
R894 VTAIL.n128 VTAIL.n126 0.388379
R895 VTAIL.n104 VTAIL.n102 0.388379
R896 VTAIL.n80 VTAIL.n78 0.388379
R897 VTAIL.n181 VTAIL.n173 0.155672
R898 VTAIL.n182 VTAIL.n181 0.155672
R899 VTAIL.n182 VTAIL.n169 0.155672
R900 VTAIL.n189 VTAIL.n169 0.155672
R901 VTAIL.n13 VTAIL.n5 0.155672
R902 VTAIL.n14 VTAIL.n13 0.155672
R903 VTAIL.n14 VTAIL.n1 0.155672
R904 VTAIL.n21 VTAIL.n1 0.155672
R905 VTAIL.n37 VTAIL.n29 0.155672
R906 VTAIL.n38 VTAIL.n37 0.155672
R907 VTAIL.n38 VTAIL.n25 0.155672
R908 VTAIL.n45 VTAIL.n25 0.155672
R909 VTAIL.n61 VTAIL.n53 0.155672
R910 VTAIL.n62 VTAIL.n61 0.155672
R911 VTAIL.n62 VTAIL.n49 0.155672
R912 VTAIL.n69 VTAIL.n49 0.155672
R913 VTAIL.n165 VTAIL.n145 0.155672
R914 VTAIL.n158 VTAIL.n145 0.155672
R915 VTAIL.n158 VTAIL.n157 0.155672
R916 VTAIL.n157 VTAIL.n149 0.155672
R917 VTAIL.n141 VTAIL.n121 0.155672
R918 VTAIL.n134 VTAIL.n121 0.155672
R919 VTAIL.n134 VTAIL.n133 0.155672
R920 VTAIL.n133 VTAIL.n125 0.155672
R921 VTAIL.n117 VTAIL.n97 0.155672
R922 VTAIL.n110 VTAIL.n97 0.155672
R923 VTAIL.n110 VTAIL.n109 0.155672
R924 VTAIL.n109 VTAIL.n101 0.155672
R925 VTAIL.n93 VTAIL.n73 0.155672
R926 VTAIL.n86 VTAIL.n73 0.155672
R927 VTAIL.n86 VTAIL.n85 0.155672
R928 VTAIL.n85 VTAIL.n77 0.155672
R929 VN.n0 VN.t0 120.371
R930 VN.n1 VN.t1 120.371
R931 VN.n0 VN.t2 120.138
R932 VN.n1 VN.t3 120.138
R933 VN VN.n1 54.9541
R934 VN VN.n0 17.564
R935 VDD2.n2 VDD2.n0 138.578
R936 VDD2.n2 VDD2.n1 106.406
R937 VDD2.n1 VDD2.t0 6.94601
R938 VDD2.n1 VDD2.t2 6.94601
R939 VDD2.n0 VDD2.t3 6.94601
R940 VDD2.n0 VDD2.t1 6.94601
R941 VDD2 VDD2.n2 0.0586897
C0 VDD2 VTAIL 3.36237f
C1 VDD2 VP 0.321052f
C2 VN VTAIL 1.88594f
C3 VN VP 3.94986f
C4 VDD1 VTAIL 3.31634f
C5 VDD1 VP 1.95097f
C6 VTAIL w_n1996_n1904# 2.26078f
C7 B VTAIL 2.1101f
C8 VP w_n1996_n1904# 3.25765f
C9 B VP 1.21012f
C10 VDD2 VN 1.78265f
C11 VDD2 VDD1 0.728177f
C12 VDD2 w_n1996_n1904# 1.03922f
C13 VDD2 B 0.88175f
C14 VDD1 VN 0.151958f
C15 VN w_n1996_n1904# 3.00423f
C16 B VN 0.795197f
C17 VDD1 w_n1996_n1904# 1.01056f
C18 VDD1 B 0.849423f
C19 B w_n1996_n1904# 5.69691f
C20 VP VTAIL 1.90004f
C21 VDD2 VSUBS 0.534507f
C22 VDD1 VSUBS 2.783171f
C23 VTAIL VSUBS 0.494918f
C24 VN VSUBS 3.89814f
C25 VP VSUBS 1.262747f
C26 B VSUBS 2.486744f
C27 w_n1996_n1904# VSUBS 47.6884f
C28 VDD2.t3 VSUBS 0.066295f
C29 VDD2.t1 VSUBS 0.066295f
C30 VDD2.n0 VSUBS 0.610321f
C31 VDD2.t0 VSUBS 0.066295f
C32 VDD2.t2 VSUBS 0.066295f
C33 VDD2.n1 VSUBS 0.408707f
C34 VDD2.n2 VSUBS 2.02678f
C35 VN.t0 VSUBS 0.734305f
C36 VN.t2 VSUBS 0.733547f
C37 VN.n0 VSUBS 0.571806f
C38 VN.t1 VSUBS 0.734305f
C39 VN.t3 VSUBS 0.733547f
C40 VN.n1 VSUBS 1.51949f
C41 VTAIL.n0 VSUBS 0.022803f
C42 VTAIL.n1 VSUBS 0.020514f
C43 VTAIL.n2 VSUBS 0.011024f
C44 VTAIL.n3 VSUBS 0.026056f
C45 VTAIL.n4 VSUBS 0.011672f
C46 VTAIL.n5 VSUBS 0.345671f
C47 VTAIL.n6 VSUBS 0.011024f
C48 VTAIL.t1 VSUBS 0.056967f
C49 VTAIL.n7 VSUBS 0.083637f
C50 VTAIL.n8 VSUBS 0.016507f
C51 VTAIL.n9 VSUBS 0.019542f
C52 VTAIL.n10 VSUBS 0.026056f
C53 VTAIL.n11 VSUBS 0.011672f
C54 VTAIL.n12 VSUBS 0.011024f
C55 VTAIL.n13 VSUBS 0.020514f
C56 VTAIL.n14 VSUBS 0.020514f
C57 VTAIL.n15 VSUBS 0.011024f
C58 VTAIL.n16 VSUBS 0.011672f
C59 VTAIL.n17 VSUBS 0.026056f
C60 VTAIL.n18 VSUBS 0.063971f
C61 VTAIL.n19 VSUBS 0.011672f
C62 VTAIL.n20 VSUBS 0.011024f
C63 VTAIL.n21 VSUBS 0.050781f
C64 VTAIL.n22 VSUBS 0.03231f
C65 VTAIL.n23 VSUBS 0.103047f
C66 VTAIL.n24 VSUBS 0.022803f
C67 VTAIL.n25 VSUBS 0.020514f
C68 VTAIL.n26 VSUBS 0.011024f
C69 VTAIL.n27 VSUBS 0.026056f
C70 VTAIL.n28 VSUBS 0.011672f
C71 VTAIL.n29 VSUBS 0.345671f
C72 VTAIL.n30 VSUBS 0.011024f
C73 VTAIL.t6 VSUBS 0.056967f
C74 VTAIL.n31 VSUBS 0.083637f
C75 VTAIL.n32 VSUBS 0.016507f
C76 VTAIL.n33 VSUBS 0.019542f
C77 VTAIL.n34 VSUBS 0.026056f
C78 VTAIL.n35 VSUBS 0.011672f
C79 VTAIL.n36 VSUBS 0.011024f
C80 VTAIL.n37 VSUBS 0.020514f
C81 VTAIL.n38 VSUBS 0.020514f
C82 VTAIL.n39 VSUBS 0.011024f
C83 VTAIL.n40 VSUBS 0.011672f
C84 VTAIL.n41 VSUBS 0.026056f
C85 VTAIL.n42 VSUBS 0.063971f
C86 VTAIL.n43 VSUBS 0.011672f
C87 VTAIL.n44 VSUBS 0.011024f
C88 VTAIL.n45 VSUBS 0.050781f
C89 VTAIL.n46 VSUBS 0.03231f
C90 VTAIL.n47 VSUBS 0.147923f
C91 VTAIL.n48 VSUBS 0.022803f
C92 VTAIL.n49 VSUBS 0.020514f
C93 VTAIL.n50 VSUBS 0.011024f
C94 VTAIL.n51 VSUBS 0.026056f
C95 VTAIL.n52 VSUBS 0.011672f
C96 VTAIL.n53 VSUBS 0.345671f
C97 VTAIL.n54 VSUBS 0.011024f
C98 VTAIL.t5 VSUBS 0.056967f
C99 VTAIL.n55 VSUBS 0.083637f
C100 VTAIL.n56 VSUBS 0.016507f
C101 VTAIL.n57 VSUBS 0.019542f
C102 VTAIL.n58 VSUBS 0.026056f
C103 VTAIL.n59 VSUBS 0.011672f
C104 VTAIL.n60 VSUBS 0.011024f
C105 VTAIL.n61 VSUBS 0.020514f
C106 VTAIL.n62 VSUBS 0.020514f
C107 VTAIL.n63 VSUBS 0.011024f
C108 VTAIL.n64 VSUBS 0.011672f
C109 VTAIL.n65 VSUBS 0.026056f
C110 VTAIL.n66 VSUBS 0.063971f
C111 VTAIL.n67 VSUBS 0.011672f
C112 VTAIL.n68 VSUBS 0.011024f
C113 VTAIL.n69 VSUBS 0.050781f
C114 VTAIL.n70 VSUBS 0.03231f
C115 VTAIL.n71 VSUBS 0.759664f
C116 VTAIL.n72 VSUBS 0.022803f
C117 VTAIL.n73 VSUBS 0.020514f
C118 VTAIL.n74 VSUBS 0.011024f
C119 VTAIL.n75 VSUBS 0.026056f
C120 VTAIL.n76 VSUBS 0.011672f
C121 VTAIL.n77 VSUBS 0.345671f
C122 VTAIL.n78 VSUBS 0.011024f
C123 VTAIL.t3 VSUBS 0.056967f
C124 VTAIL.n79 VSUBS 0.083637f
C125 VTAIL.n80 VSUBS 0.016507f
C126 VTAIL.n81 VSUBS 0.019542f
C127 VTAIL.n82 VSUBS 0.026056f
C128 VTAIL.n83 VSUBS 0.011672f
C129 VTAIL.n84 VSUBS 0.011024f
C130 VTAIL.n85 VSUBS 0.020514f
C131 VTAIL.n86 VSUBS 0.020514f
C132 VTAIL.n87 VSUBS 0.011024f
C133 VTAIL.n88 VSUBS 0.011672f
C134 VTAIL.n89 VSUBS 0.026056f
C135 VTAIL.n90 VSUBS 0.063971f
C136 VTAIL.n91 VSUBS 0.011672f
C137 VTAIL.n92 VSUBS 0.011024f
C138 VTAIL.n93 VSUBS 0.050781f
C139 VTAIL.n94 VSUBS 0.03231f
C140 VTAIL.n95 VSUBS 0.759664f
C141 VTAIL.n96 VSUBS 0.022803f
C142 VTAIL.n97 VSUBS 0.020514f
C143 VTAIL.n98 VSUBS 0.011024f
C144 VTAIL.n99 VSUBS 0.026056f
C145 VTAIL.n100 VSUBS 0.011672f
C146 VTAIL.n101 VSUBS 0.345671f
C147 VTAIL.n102 VSUBS 0.011024f
C148 VTAIL.t2 VSUBS 0.056967f
C149 VTAIL.n103 VSUBS 0.083637f
C150 VTAIL.n104 VSUBS 0.016507f
C151 VTAIL.n105 VSUBS 0.019542f
C152 VTAIL.n106 VSUBS 0.026056f
C153 VTAIL.n107 VSUBS 0.011672f
C154 VTAIL.n108 VSUBS 0.011024f
C155 VTAIL.n109 VSUBS 0.020514f
C156 VTAIL.n110 VSUBS 0.020514f
C157 VTAIL.n111 VSUBS 0.011024f
C158 VTAIL.n112 VSUBS 0.011672f
C159 VTAIL.n113 VSUBS 0.026056f
C160 VTAIL.n114 VSUBS 0.063971f
C161 VTAIL.n115 VSUBS 0.011672f
C162 VTAIL.n116 VSUBS 0.011024f
C163 VTAIL.n117 VSUBS 0.050781f
C164 VTAIL.n118 VSUBS 0.03231f
C165 VTAIL.n119 VSUBS 0.147923f
C166 VTAIL.n120 VSUBS 0.022803f
C167 VTAIL.n121 VSUBS 0.020514f
C168 VTAIL.n122 VSUBS 0.011024f
C169 VTAIL.n123 VSUBS 0.026056f
C170 VTAIL.n124 VSUBS 0.011672f
C171 VTAIL.n125 VSUBS 0.345671f
C172 VTAIL.n126 VSUBS 0.011024f
C173 VTAIL.t7 VSUBS 0.056967f
C174 VTAIL.n127 VSUBS 0.083637f
C175 VTAIL.n128 VSUBS 0.016507f
C176 VTAIL.n129 VSUBS 0.019542f
C177 VTAIL.n130 VSUBS 0.026056f
C178 VTAIL.n131 VSUBS 0.011672f
C179 VTAIL.n132 VSUBS 0.011024f
C180 VTAIL.n133 VSUBS 0.020514f
C181 VTAIL.n134 VSUBS 0.020514f
C182 VTAIL.n135 VSUBS 0.011024f
C183 VTAIL.n136 VSUBS 0.011672f
C184 VTAIL.n137 VSUBS 0.026056f
C185 VTAIL.n138 VSUBS 0.063971f
C186 VTAIL.n139 VSUBS 0.011672f
C187 VTAIL.n140 VSUBS 0.011024f
C188 VTAIL.n141 VSUBS 0.050781f
C189 VTAIL.n142 VSUBS 0.03231f
C190 VTAIL.n143 VSUBS 0.147923f
C191 VTAIL.n144 VSUBS 0.022803f
C192 VTAIL.n145 VSUBS 0.020514f
C193 VTAIL.n146 VSUBS 0.011024f
C194 VTAIL.n147 VSUBS 0.026056f
C195 VTAIL.n148 VSUBS 0.011672f
C196 VTAIL.n149 VSUBS 0.345671f
C197 VTAIL.n150 VSUBS 0.011024f
C198 VTAIL.t4 VSUBS 0.056967f
C199 VTAIL.n151 VSUBS 0.083637f
C200 VTAIL.n152 VSUBS 0.016507f
C201 VTAIL.n153 VSUBS 0.019542f
C202 VTAIL.n154 VSUBS 0.026056f
C203 VTAIL.n155 VSUBS 0.011672f
C204 VTAIL.n156 VSUBS 0.011024f
C205 VTAIL.n157 VSUBS 0.020514f
C206 VTAIL.n158 VSUBS 0.020514f
C207 VTAIL.n159 VSUBS 0.011024f
C208 VTAIL.n160 VSUBS 0.011672f
C209 VTAIL.n161 VSUBS 0.026056f
C210 VTAIL.n162 VSUBS 0.063971f
C211 VTAIL.n163 VSUBS 0.011672f
C212 VTAIL.n164 VSUBS 0.011024f
C213 VTAIL.n165 VSUBS 0.050781f
C214 VTAIL.n166 VSUBS 0.03231f
C215 VTAIL.n167 VSUBS 0.759664f
C216 VTAIL.n168 VSUBS 0.022803f
C217 VTAIL.n169 VSUBS 0.020514f
C218 VTAIL.n170 VSUBS 0.011024f
C219 VTAIL.n171 VSUBS 0.026056f
C220 VTAIL.n172 VSUBS 0.011672f
C221 VTAIL.n173 VSUBS 0.345671f
C222 VTAIL.n174 VSUBS 0.011024f
C223 VTAIL.t0 VSUBS 0.056967f
C224 VTAIL.n175 VSUBS 0.083637f
C225 VTAIL.n176 VSUBS 0.016507f
C226 VTAIL.n177 VSUBS 0.019542f
C227 VTAIL.n178 VSUBS 0.026056f
C228 VTAIL.n179 VSUBS 0.011672f
C229 VTAIL.n180 VSUBS 0.011024f
C230 VTAIL.n181 VSUBS 0.020514f
C231 VTAIL.n182 VSUBS 0.020514f
C232 VTAIL.n183 VSUBS 0.011024f
C233 VTAIL.n184 VSUBS 0.011672f
C234 VTAIL.n185 VSUBS 0.026056f
C235 VTAIL.n186 VSUBS 0.063971f
C236 VTAIL.n187 VSUBS 0.011672f
C237 VTAIL.n188 VSUBS 0.011024f
C238 VTAIL.n189 VSUBS 0.050781f
C239 VTAIL.n190 VSUBS 0.03231f
C240 VTAIL.n191 VSUBS 0.707095f
C241 VDD1.t1 VSUBS 0.063116f
C242 VDD1.t0 VSUBS 0.063116f
C243 VDD1.n0 VSUBS 0.389298f
C244 VDD1.t2 VSUBS 0.063116f
C245 VDD1.t3 VSUBS 0.063116f
C246 VDD1.n1 VSUBS 0.591651f
C247 VP.n0 VSUBS 0.038157f
C248 VP.t1 VSUBS 0.641427f
C249 VP.n1 VSUBS 0.065307f
C250 VP.t0 VSUBS 0.771939f
C251 VP.t3 VSUBS 0.771142f
C252 VP.n2 VSUBS 1.57696f
C253 VP.t2 VSUBS 0.641427f
C254 VP.n3 VSUBS 0.348622f
C255 VP.n4 VSUBS 1.76823f
C256 VP.n5 VSUBS 0.038157f
C257 VP.n6 VSUBS 0.038157f
C258 VP.n7 VSUBS 0.030818f
C259 VP.n8 VSUBS 0.065307f
C260 VP.n9 VSUBS 0.348622f
C261 VP.n10 VSUBS 0.033261f
C262 B.n0 VSUBS 0.005939f
C263 B.n1 VSUBS 0.005939f
C264 B.n2 VSUBS 0.009392f
C265 B.n3 VSUBS 0.009392f
C266 B.n4 VSUBS 0.009392f
C267 B.n5 VSUBS 0.009392f
C268 B.n6 VSUBS 0.009392f
C269 B.n7 VSUBS 0.009392f
C270 B.n8 VSUBS 0.009392f
C271 B.n9 VSUBS 0.009392f
C272 B.n10 VSUBS 0.009392f
C273 B.n11 VSUBS 0.009392f
C274 B.n12 VSUBS 0.009392f
C275 B.n13 VSUBS 0.021425f
C276 B.n14 VSUBS 0.009392f
C277 B.n15 VSUBS 0.009392f
C278 B.n16 VSUBS 0.009392f
C279 B.n17 VSUBS 0.009392f
C280 B.n18 VSUBS 0.009392f
C281 B.n19 VSUBS 0.009392f
C282 B.n20 VSUBS 0.009392f
C283 B.n21 VSUBS 0.009392f
C284 B.n22 VSUBS 0.009392f
C285 B.n23 VSUBS 0.009392f
C286 B.t5 VSUBS 0.091206f
C287 B.t4 VSUBS 0.109572f
C288 B.t3 VSUBS 0.401117f
C289 B.n24 VSUBS 0.196521f
C290 B.n25 VSUBS 0.167937f
C291 B.n26 VSUBS 0.009392f
C292 B.n27 VSUBS 0.009392f
C293 B.n28 VSUBS 0.009392f
C294 B.n29 VSUBS 0.009392f
C295 B.n30 VSUBS 0.005248f
C296 B.n31 VSUBS 0.009392f
C297 B.t2 VSUBS 0.091208f
C298 B.t1 VSUBS 0.109574f
C299 B.t0 VSUBS 0.401117f
C300 B.n32 VSUBS 0.19652f
C301 B.n33 VSUBS 0.167936f
C302 B.n34 VSUBS 0.02176f
C303 B.n35 VSUBS 0.009392f
C304 B.n36 VSUBS 0.009392f
C305 B.n37 VSUBS 0.009392f
C306 B.n38 VSUBS 0.009392f
C307 B.n39 VSUBS 0.009392f
C308 B.n40 VSUBS 0.009392f
C309 B.n41 VSUBS 0.009392f
C310 B.n42 VSUBS 0.009392f
C311 B.n43 VSUBS 0.021957f
C312 B.n44 VSUBS 0.009392f
C313 B.n45 VSUBS 0.009392f
C314 B.n46 VSUBS 0.009392f
C315 B.n47 VSUBS 0.009392f
C316 B.n48 VSUBS 0.009392f
C317 B.n49 VSUBS 0.009392f
C318 B.n50 VSUBS 0.009392f
C319 B.n51 VSUBS 0.009392f
C320 B.n52 VSUBS 0.009392f
C321 B.n53 VSUBS 0.009392f
C322 B.n54 VSUBS 0.009392f
C323 B.n55 VSUBS 0.009392f
C324 B.n56 VSUBS 0.009392f
C325 B.n57 VSUBS 0.009392f
C326 B.n58 VSUBS 0.009392f
C327 B.n59 VSUBS 0.009392f
C328 B.n60 VSUBS 0.009392f
C329 B.n61 VSUBS 0.009392f
C330 B.n62 VSUBS 0.009392f
C331 B.n63 VSUBS 0.009392f
C332 B.n64 VSUBS 0.009392f
C333 B.n65 VSUBS 0.009392f
C334 B.n66 VSUBS 0.009392f
C335 B.n67 VSUBS 0.023047f
C336 B.n68 VSUBS 0.009392f
C337 B.n69 VSUBS 0.009392f
C338 B.n70 VSUBS 0.009392f
C339 B.n71 VSUBS 0.009392f
C340 B.n72 VSUBS 0.009392f
C341 B.n73 VSUBS 0.009392f
C342 B.n74 VSUBS 0.009392f
C343 B.n75 VSUBS 0.009392f
C344 B.n76 VSUBS 0.009392f
C345 B.t7 VSUBS 0.091208f
C346 B.t8 VSUBS 0.109574f
C347 B.t6 VSUBS 0.401117f
C348 B.n77 VSUBS 0.19652f
C349 B.n78 VSUBS 0.167936f
C350 B.n79 VSUBS 0.02176f
C351 B.n80 VSUBS 0.009392f
C352 B.n81 VSUBS 0.009392f
C353 B.n82 VSUBS 0.009392f
C354 B.n83 VSUBS 0.009392f
C355 B.n84 VSUBS 0.009392f
C356 B.t10 VSUBS 0.091206f
C357 B.t11 VSUBS 0.109572f
C358 B.t9 VSUBS 0.401117f
C359 B.n85 VSUBS 0.196521f
C360 B.n86 VSUBS 0.167937f
C361 B.n87 VSUBS 0.009392f
C362 B.n88 VSUBS 0.009392f
C363 B.n89 VSUBS 0.009392f
C364 B.n90 VSUBS 0.009392f
C365 B.n91 VSUBS 0.009392f
C366 B.n92 VSUBS 0.009392f
C367 B.n93 VSUBS 0.009392f
C368 B.n94 VSUBS 0.009392f
C369 B.n95 VSUBS 0.009392f
C370 B.n96 VSUBS 0.023047f
C371 B.n97 VSUBS 0.009392f
C372 B.n98 VSUBS 0.009392f
C373 B.n99 VSUBS 0.009392f
C374 B.n100 VSUBS 0.009392f
C375 B.n101 VSUBS 0.009392f
C376 B.n102 VSUBS 0.009392f
C377 B.n103 VSUBS 0.009392f
C378 B.n104 VSUBS 0.009392f
C379 B.n105 VSUBS 0.009392f
C380 B.n106 VSUBS 0.009392f
C381 B.n107 VSUBS 0.009392f
C382 B.n108 VSUBS 0.009392f
C383 B.n109 VSUBS 0.009392f
C384 B.n110 VSUBS 0.009392f
C385 B.n111 VSUBS 0.009392f
C386 B.n112 VSUBS 0.009392f
C387 B.n113 VSUBS 0.009392f
C388 B.n114 VSUBS 0.009392f
C389 B.n115 VSUBS 0.009392f
C390 B.n116 VSUBS 0.009392f
C391 B.n117 VSUBS 0.009392f
C392 B.n118 VSUBS 0.009392f
C393 B.n119 VSUBS 0.009392f
C394 B.n120 VSUBS 0.009392f
C395 B.n121 VSUBS 0.009392f
C396 B.n122 VSUBS 0.009392f
C397 B.n123 VSUBS 0.009392f
C398 B.n124 VSUBS 0.009392f
C399 B.n125 VSUBS 0.009392f
C400 B.n126 VSUBS 0.009392f
C401 B.n127 VSUBS 0.009392f
C402 B.n128 VSUBS 0.009392f
C403 B.n129 VSUBS 0.009392f
C404 B.n130 VSUBS 0.009392f
C405 B.n131 VSUBS 0.009392f
C406 B.n132 VSUBS 0.009392f
C407 B.n133 VSUBS 0.009392f
C408 B.n134 VSUBS 0.009392f
C409 B.n135 VSUBS 0.009392f
C410 B.n136 VSUBS 0.009392f
C411 B.n137 VSUBS 0.009392f
C412 B.n138 VSUBS 0.009392f
C413 B.n139 VSUBS 0.021425f
C414 B.n140 VSUBS 0.021425f
C415 B.n141 VSUBS 0.023047f
C416 B.n142 VSUBS 0.009392f
C417 B.n143 VSUBS 0.009392f
C418 B.n144 VSUBS 0.009392f
C419 B.n145 VSUBS 0.009392f
C420 B.n146 VSUBS 0.009392f
C421 B.n147 VSUBS 0.009392f
C422 B.n148 VSUBS 0.009392f
C423 B.n149 VSUBS 0.009392f
C424 B.n150 VSUBS 0.009392f
C425 B.n151 VSUBS 0.009392f
C426 B.n152 VSUBS 0.009392f
C427 B.n153 VSUBS 0.009392f
C428 B.n154 VSUBS 0.009392f
C429 B.n155 VSUBS 0.009392f
C430 B.n156 VSUBS 0.009392f
C431 B.n157 VSUBS 0.009392f
C432 B.n158 VSUBS 0.009392f
C433 B.n159 VSUBS 0.009392f
C434 B.n160 VSUBS 0.009392f
C435 B.n161 VSUBS 0.009392f
C436 B.n162 VSUBS 0.009392f
C437 B.n163 VSUBS 0.009392f
C438 B.n164 VSUBS 0.009392f
C439 B.n165 VSUBS 0.009392f
C440 B.n166 VSUBS 0.009392f
C441 B.n167 VSUBS 0.009392f
C442 B.n168 VSUBS 0.009392f
C443 B.n169 VSUBS 0.009392f
C444 B.n170 VSUBS 0.008839f
C445 B.n171 VSUBS 0.02176f
C446 B.n172 VSUBS 0.005248f
C447 B.n173 VSUBS 0.009392f
C448 B.n174 VSUBS 0.009392f
C449 B.n175 VSUBS 0.009392f
C450 B.n176 VSUBS 0.009392f
C451 B.n177 VSUBS 0.009392f
C452 B.n178 VSUBS 0.009392f
C453 B.n179 VSUBS 0.009392f
C454 B.n180 VSUBS 0.009392f
C455 B.n181 VSUBS 0.009392f
C456 B.n182 VSUBS 0.009392f
C457 B.n183 VSUBS 0.009392f
C458 B.n184 VSUBS 0.009392f
C459 B.n185 VSUBS 0.005248f
C460 B.n186 VSUBS 0.009392f
C461 B.n187 VSUBS 0.009392f
C462 B.n188 VSUBS 0.008839f
C463 B.n189 VSUBS 0.009392f
C464 B.n190 VSUBS 0.009392f
C465 B.n191 VSUBS 0.009392f
C466 B.n192 VSUBS 0.009392f
C467 B.n193 VSUBS 0.009392f
C468 B.n194 VSUBS 0.009392f
C469 B.n195 VSUBS 0.009392f
C470 B.n196 VSUBS 0.009392f
C471 B.n197 VSUBS 0.009392f
C472 B.n198 VSUBS 0.009392f
C473 B.n199 VSUBS 0.009392f
C474 B.n200 VSUBS 0.009392f
C475 B.n201 VSUBS 0.009392f
C476 B.n202 VSUBS 0.009392f
C477 B.n203 VSUBS 0.009392f
C478 B.n204 VSUBS 0.009392f
C479 B.n205 VSUBS 0.009392f
C480 B.n206 VSUBS 0.009392f
C481 B.n207 VSUBS 0.009392f
C482 B.n208 VSUBS 0.009392f
C483 B.n209 VSUBS 0.009392f
C484 B.n210 VSUBS 0.009392f
C485 B.n211 VSUBS 0.009392f
C486 B.n212 VSUBS 0.009392f
C487 B.n213 VSUBS 0.009392f
C488 B.n214 VSUBS 0.009392f
C489 B.n215 VSUBS 0.009392f
C490 B.n216 VSUBS 0.023047f
C491 B.n217 VSUBS 0.021425f
C492 B.n218 VSUBS 0.021425f
C493 B.n219 VSUBS 0.009392f
C494 B.n220 VSUBS 0.009392f
C495 B.n221 VSUBS 0.009392f
C496 B.n222 VSUBS 0.009392f
C497 B.n223 VSUBS 0.009392f
C498 B.n224 VSUBS 0.009392f
C499 B.n225 VSUBS 0.009392f
C500 B.n226 VSUBS 0.009392f
C501 B.n227 VSUBS 0.009392f
C502 B.n228 VSUBS 0.009392f
C503 B.n229 VSUBS 0.009392f
C504 B.n230 VSUBS 0.009392f
C505 B.n231 VSUBS 0.009392f
C506 B.n232 VSUBS 0.009392f
C507 B.n233 VSUBS 0.009392f
C508 B.n234 VSUBS 0.009392f
C509 B.n235 VSUBS 0.009392f
C510 B.n236 VSUBS 0.009392f
C511 B.n237 VSUBS 0.009392f
C512 B.n238 VSUBS 0.009392f
C513 B.n239 VSUBS 0.009392f
C514 B.n240 VSUBS 0.009392f
C515 B.n241 VSUBS 0.009392f
C516 B.n242 VSUBS 0.009392f
C517 B.n243 VSUBS 0.009392f
C518 B.n244 VSUBS 0.009392f
C519 B.n245 VSUBS 0.009392f
C520 B.n246 VSUBS 0.009392f
C521 B.n247 VSUBS 0.009392f
C522 B.n248 VSUBS 0.009392f
C523 B.n249 VSUBS 0.009392f
C524 B.n250 VSUBS 0.009392f
C525 B.n251 VSUBS 0.009392f
C526 B.n252 VSUBS 0.009392f
C527 B.n253 VSUBS 0.009392f
C528 B.n254 VSUBS 0.009392f
C529 B.n255 VSUBS 0.009392f
C530 B.n256 VSUBS 0.009392f
C531 B.n257 VSUBS 0.009392f
C532 B.n258 VSUBS 0.009392f
C533 B.n259 VSUBS 0.009392f
C534 B.n260 VSUBS 0.009392f
C535 B.n261 VSUBS 0.009392f
C536 B.n262 VSUBS 0.009392f
C537 B.n263 VSUBS 0.009392f
C538 B.n264 VSUBS 0.009392f
C539 B.n265 VSUBS 0.009392f
C540 B.n266 VSUBS 0.009392f
C541 B.n267 VSUBS 0.009392f
C542 B.n268 VSUBS 0.009392f
C543 B.n269 VSUBS 0.009392f
C544 B.n270 VSUBS 0.009392f
C545 B.n271 VSUBS 0.009392f
C546 B.n272 VSUBS 0.009392f
C547 B.n273 VSUBS 0.009392f
C548 B.n274 VSUBS 0.009392f
C549 B.n275 VSUBS 0.009392f
C550 B.n276 VSUBS 0.009392f
C551 B.n277 VSUBS 0.009392f
C552 B.n278 VSUBS 0.009392f
C553 B.n279 VSUBS 0.009392f
C554 B.n280 VSUBS 0.009392f
C555 B.n281 VSUBS 0.009392f
C556 B.n282 VSUBS 0.009392f
C557 B.n283 VSUBS 0.009392f
C558 B.n284 VSUBS 0.009392f
C559 B.n285 VSUBS 0.009392f
C560 B.n286 VSUBS 0.022515f
C561 B.n287 VSUBS 0.021425f
C562 B.n288 VSUBS 0.023047f
C563 B.n289 VSUBS 0.009392f
C564 B.n290 VSUBS 0.009392f
C565 B.n291 VSUBS 0.009392f
C566 B.n292 VSUBS 0.009392f
C567 B.n293 VSUBS 0.009392f
C568 B.n294 VSUBS 0.009392f
C569 B.n295 VSUBS 0.009392f
C570 B.n296 VSUBS 0.009392f
C571 B.n297 VSUBS 0.009392f
C572 B.n298 VSUBS 0.009392f
C573 B.n299 VSUBS 0.009392f
C574 B.n300 VSUBS 0.009392f
C575 B.n301 VSUBS 0.009392f
C576 B.n302 VSUBS 0.009392f
C577 B.n303 VSUBS 0.009392f
C578 B.n304 VSUBS 0.009392f
C579 B.n305 VSUBS 0.009392f
C580 B.n306 VSUBS 0.009392f
C581 B.n307 VSUBS 0.009392f
C582 B.n308 VSUBS 0.009392f
C583 B.n309 VSUBS 0.009392f
C584 B.n310 VSUBS 0.009392f
C585 B.n311 VSUBS 0.009392f
C586 B.n312 VSUBS 0.009392f
C587 B.n313 VSUBS 0.009392f
C588 B.n314 VSUBS 0.009392f
C589 B.n315 VSUBS 0.009392f
C590 B.n316 VSUBS 0.008839f
C591 B.n317 VSUBS 0.009392f
C592 B.n318 VSUBS 0.009392f
C593 B.n319 VSUBS 0.009392f
C594 B.n320 VSUBS 0.009392f
C595 B.n321 VSUBS 0.009392f
C596 B.n322 VSUBS 0.009392f
C597 B.n323 VSUBS 0.009392f
C598 B.n324 VSUBS 0.009392f
C599 B.n325 VSUBS 0.009392f
C600 B.n326 VSUBS 0.009392f
C601 B.n327 VSUBS 0.009392f
C602 B.n328 VSUBS 0.009392f
C603 B.n329 VSUBS 0.009392f
C604 B.n330 VSUBS 0.009392f
C605 B.n331 VSUBS 0.009392f
C606 B.n332 VSUBS 0.005248f
C607 B.n333 VSUBS 0.02176f
C608 B.n334 VSUBS 0.008839f
C609 B.n335 VSUBS 0.009392f
C610 B.n336 VSUBS 0.009392f
C611 B.n337 VSUBS 0.009392f
C612 B.n338 VSUBS 0.009392f
C613 B.n339 VSUBS 0.009392f
C614 B.n340 VSUBS 0.009392f
C615 B.n341 VSUBS 0.009392f
C616 B.n342 VSUBS 0.009392f
C617 B.n343 VSUBS 0.009392f
C618 B.n344 VSUBS 0.009392f
C619 B.n345 VSUBS 0.009392f
C620 B.n346 VSUBS 0.009392f
C621 B.n347 VSUBS 0.009392f
C622 B.n348 VSUBS 0.009392f
C623 B.n349 VSUBS 0.009392f
C624 B.n350 VSUBS 0.009392f
C625 B.n351 VSUBS 0.009392f
C626 B.n352 VSUBS 0.009392f
C627 B.n353 VSUBS 0.009392f
C628 B.n354 VSUBS 0.009392f
C629 B.n355 VSUBS 0.009392f
C630 B.n356 VSUBS 0.009392f
C631 B.n357 VSUBS 0.009392f
C632 B.n358 VSUBS 0.009392f
C633 B.n359 VSUBS 0.009392f
C634 B.n360 VSUBS 0.009392f
C635 B.n361 VSUBS 0.009392f
C636 B.n362 VSUBS 0.023047f
C637 B.n363 VSUBS 0.023047f
C638 B.n364 VSUBS 0.021425f
C639 B.n365 VSUBS 0.009392f
C640 B.n366 VSUBS 0.009392f
C641 B.n367 VSUBS 0.009392f
C642 B.n368 VSUBS 0.009392f
C643 B.n369 VSUBS 0.009392f
C644 B.n370 VSUBS 0.009392f
C645 B.n371 VSUBS 0.009392f
C646 B.n372 VSUBS 0.009392f
C647 B.n373 VSUBS 0.009392f
C648 B.n374 VSUBS 0.009392f
C649 B.n375 VSUBS 0.009392f
C650 B.n376 VSUBS 0.009392f
C651 B.n377 VSUBS 0.009392f
C652 B.n378 VSUBS 0.009392f
C653 B.n379 VSUBS 0.009392f
C654 B.n380 VSUBS 0.009392f
C655 B.n381 VSUBS 0.009392f
C656 B.n382 VSUBS 0.009392f
C657 B.n383 VSUBS 0.009392f
C658 B.n384 VSUBS 0.009392f
C659 B.n385 VSUBS 0.009392f
C660 B.n386 VSUBS 0.009392f
C661 B.n387 VSUBS 0.009392f
C662 B.n388 VSUBS 0.009392f
C663 B.n389 VSUBS 0.009392f
C664 B.n390 VSUBS 0.009392f
C665 B.n391 VSUBS 0.009392f
C666 B.n392 VSUBS 0.009392f
C667 B.n393 VSUBS 0.009392f
C668 B.n394 VSUBS 0.009392f
C669 B.n395 VSUBS 0.009392f
C670 B.n396 VSUBS 0.009392f
C671 B.n397 VSUBS 0.009392f
C672 B.n398 VSUBS 0.009392f
C673 B.n399 VSUBS 0.021266f
.ends

