* NGSPICE file created from diff_pair_sample_1322.ext - technology: sky130A

.subckt diff_pair_sample_1322 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=0 ps=0 w=15.54 l=0.87
X1 VTAIL.t10 VP.t0 VDD1.t1 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=2.5641 ps=15.87 w=15.54 l=0.87
X2 VDD1.t0 VP.t1 VTAIL.t9 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=2.5641 ps=15.87 w=15.54 l=0.87
X3 VDD1.t5 VP.t2 VTAIL.t8 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=6.0606 ps=31.86 w=15.54 l=0.87
X4 VDD1.t4 VP.t3 VTAIL.t7 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=2.5641 ps=15.87 w=15.54 l=0.87
X5 VDD2.t5 VN.t0 VTAIL.t1 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=6.0606 ps=31.86 w=15.54 l=0.87
X6 VDD2.t4 VN.t1 VTAIL.t0 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=2.5641 ps=15.87 w=15.54 l=0.87
X7 B.t8 B.t6 B.t7 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=0 ps=0 w=15.54 l=0.87
X8 VTAIL.t6 VP.t4 VDD1.t3 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=2.5641 ps=15.87 w=15.54 l=0.87
X9 VDD2.t3 VN.t2 VTAIL.t4 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=6.0606 ps=31.86 w=15.54 l=0.87
X10 B.t5 B.t3 B.t4 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=0 ps=0 w=15.54 l=0.87
X11 VTAIL.t2 VN.t3 VDD2.t2 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=2.5641 ps=15.87 w=15.54 l=0.87
X12 VTAIL.t3 VN.t4 VDD2.t1 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=2.5641 ps=15.87 w=15.54 l=0.87
X13 VDD1.t2 VP.t5 VTAIL.t5 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=2.5641 pd=15.87 as=6.0606 ps=31.86 w=15.54 l=0.87
X14 B.t2 B.t0 B.t1 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=0 ps=0 w=15.54 l=0.87
X15 VDD2.t0 VN.t5 VTAIL.t11 w_n1930_n4076# sky130_fd_pr__pfet_01v8 ad=6.0606 pd=31.86 as=2.5641 ps=15.87 w=15.54 l=0.87
R0 B.n124 B.t0 632.433
R1 B.n130 B.t6 632.433
R2 B.n40 B.t9 632.433
R3 B.n46 B.t3 632.433
R4 B.n441 B.n74 585
R5 B.n443 B.n442 585
R6 B.n444 B.n73 585
R7 B.n446 B.n445 585
R8 B.n447 B.n72 585
R9 B.n449 B.n448 585
R10 B.n450 B.n71 585
R11 B.n452 B.n451 585
R12 B.n453 B.n70 585
R13 B.n455 B.n454 585
R14 B.n456 B.n69 585
R15 B.n458 B.n457 585
R16 B.n459 B.n68 585
R17 B.n461 B.n460 585
R18 B.n462 B.n67 585
R19 B.n464 B.n463 585
R20 B.n465 B.n66 585
R21 B.n467 B.n466 585
R22 B.n468 B.n65 585
R23 B.n470 B.n469 585
R24 B.n471 B.n64 585
R25 B.n473 B.n472 585
R26 B.n474 B.n63 585
R27 B.n476 B.n475 585
R28 B.n477 B.n62 585
R29 B.n479 B.n478 585
R30 B.n480 B.n61 585
R31 B.n482 B.n481 585
R32 B.n483 B.n60 585
R33 B.n485 B.n484 585
R34 B.n486 B.n59 585
R35 B.n488 B.n487 585
R36 B.n489 B.n58 585
R37 B.n491 B.n490 585
R38 B.n492 B.n57 585
R39 B.n494 B.n493 585
R40 B.n495 B.n56 585
R41 B.n497 B.n496 585
R42 B.n498 B.n55 585
R43 B.n500 B.n499 585
R44 B.n501 B.n54 585
R45 B.n503 B.n502 585
R46 B.n504 B.n53 585
R47 B.n506 B.n505 585
R48 B.n507 B.n52 585
R49 B.n509 B.n508 585
R50 B.n510 B.n51 585
R51 B.n512 B.n511 585
R52 B.n513 B.n50 585
R53 B.n515 B.n514 585
R54 B.n516 B.n49 585
R55 B.n518 B.n517 585
R56 B.n520 B.n519 585
R57 B.n521 B.n45 585
R58 B.n523 B.n522 585
R59 B.n524 B.n44 585
R60 B.n526 B.n525 585
R61 B.n527 B.n43 585
R62 B.n529 B.n528 585
R63 B.n530 B.n42 585
R64 B.n532 B.n531 585
R65 B.n533 B.n39 585
R66 B.n536 B.n535 585
R67 B.n537 B.n38 585
R68 B.n539 B.n538 585
R69 B.n540 B.n37 585
R70 B.n542 B.n541 585
R71 B.n543 B.n36 585
R72 B.n545 B.n544 585
R73 B.n546 B.n35 585
R74 B.n548 B.n547 585
R75 B.n549 B.n34 585
R76 B.n551 B.n550 585
R77 B.n552 B.n33 585
R78 B.n554 B.n553 585
R79 B.n555 B.n32 585
R80 B.n557 B.n556 585
R81 B.n558 B.n31 585
R82 B.n560 B.n559 585
R83 B.n561 B.n30 585
R84 B.n563 B.n562 585
R85 B.n564 B.n29 585
R86 B.n566 B.n565 585
R87 B.n567 B.n28 585
R88 B.n569 B.n568 585
R89 B.n570 B.n27 585
R90 B.n572 B.n571 585
R91 B.n573 B.n26 585
R92 B.n575 B.n574 585
R93 B.n576 B.n25 585
R94 B.n578 B.n577 585
R95 B.n579 B.n24 585
R96 B.n581 B.n580 585
R97 B.n582 B.n23 585
R98 B.n584 B.n583 585
R99 B.n585 B.n22 585
R100 B.n587 B.n586 585
R101 B.n588 B.n21 585
R102 B.n590 B.n589 585
R103 B.n591 B.n20 585
R104 B.n593 B.n592 585
R105 B.n594 B.n19 585
R106 B.n596 B.n595 585
R107 B.n597 B.n18 585
R108 B.n599 B.n598 585
R109 B.n600 B.n17 585
R110 B.n602 B.n601 585
R111 B.n603 B.n16 585
R112 B.n605 B.n604 585
R113 B.n606 B.n15 585
R114 B.n608 B.n607 585
R115 B.n609 B.n14 585
R116 B.n611 B.n610 585
R117 B.n612 B.n13 585
R118 B.n440 B.n439 585
R119 B.n438 B.n75 585
R120 B.n437 B.n436 585
R121 B.n435 B.n76 585
R122 B.n434 B.n433 585
R123 B.n432 B.n77 585
R124 B.n431 B.n430 585
R125 B.n429 B.n78 585
R126 B.n428 B.n427 585
R127 B.n426 B.n79 585
R128 B.n425 B.n424 585
R129 B.n423 B.n80 585
R130 B.n422 B.n421 585
R131 B.n420 B.n81 585
R132 B.n419 B.n418 585
R133 B.n417 B.n82 585
R134 B.n416 B.n415 585
R135 B.n414 B.n83 585
R136 B.n413 B.n412 585
R137 B.n411 B.n84 585
R138 B.n410 B.n409 585
R139 B.n408 B.n85 585
R140 B.n407 B.n406 585
R141 B.n405 B.n86 585
R142 B.n404 B.n403 585
R143 B.n402 B.n87 585
R144 B.n401 B.n400 585
R145 B.n399 B.n88 585
R146 B.n398 B.n397 585
R147 B.n396 B.n89 585
R148 B.n395 B.n394 585
R149 B.n393 B.n90 585
R150 B.n392 B.n391 585
R151 B.n390 B.n91 585
R152 B.n389 B.n388 585
R153 B.n387 B.n92 585
R154 B.n386 B.n385 585
R155 B.n384 B.n93 585
R156 B.n383 B.n382 585
R157 B.n381 B.n94 585
R158 B.n380 B.n379 585
R159 B.n378 B.n95 585
R160 B.n377 B.n376 585
R161 B.n375 B.n96 585
R162 B.n374 B.n373 585
R163 B.n201 B.n158 585
R164 B.n203 B.n202 585
R165 B.n204 B.n157 585
R166 B.n206 B.n205 585
R167 B.n207 B.n156 585
R168 B.n209 B.n208 585
R169 B.n210 B.n155 585
R170 B.n212 B.n211 585
R171 B.n213 B.n154 585
R172 B.n215 B.n214 585
R173 B.n216 B.n153 585
R174 B.n218 B.n217 585
R175 B.n219 B.n152 585
R176 B.n221 B.n220 585
R177 B.n222 B.n151 585
R178 B.n224 B.n223 585
R179 B.n225 B.n150 585
R180 B.n227 B.n226 585
R181 B.n228 B.n149 585
R182 B.n230 B.n229 585
R183 B.n231 B.n148 585
R184 B.n233 B.n232 585
R185 B.n234 B.n147 585
R186 B.n236 B.n235 585
R187 B.n237 B.n146 585
R188 B.n239 B.n238 585
R189 B.n240 B.n145 585
R190 B.n242 B.n241 585
R191 B.n243 B.n144 585
R192 B.n245 B.n244 585
R193 B.n246 B.n143 585
R194 B.n248 B.n247 585
R195 B.n249 B.n142 585
R196 B.n251 B.n250 585
R197 B.n252 B.n141 585
R198 B.n254 B.n253 585
R199 B.n255 B.n140 585
R200 B.n257 B.n256 585
R201 B.n258 B.n139 585
R202 B.n260 B.n259 585
R203 B.n261 B.n138 585
R204 B.n263 B.n262 585
R205 B.n264 B.n137 585
R206 B.n266 B.n265 585
R207 B.n267 B.n136 585
R208 B.n269 B.n268 585
R209 B.n270 B.n135 585
R210 B.n272 B.n271 585
R211 B.n273 B.n134 585
R212 B.n275 B.n274 585
R213 B.n276 B.n133 585
R214 B.n278 B.n277 585
R215 B.n280 B.n279 585
R216 B.n281 B.n129 585
R217 B.n283 B.n282 585
R218 B.n284 B.n128 585
R219 B.n286 B.n285 585
R220 B.n287 B.n127 585
R221 B.n289 B.n288 585
R222 B.n290 B.n126 585
R223 B.n292 B.n291 585
R224 B.n293 B.n123 585
R225 B.n296 B.n295 585
R226 B.n297 B.n122 585
R227 B.n299 B.n298 585
R228 B.n300 B.n121 585
R229 B.n302 B.n301 585
R230 B.n303 B.n120 585
R231 B.n305 B.n304 585
R232 B.n306 B.n119 585
R233 B.n308 B.n307 585
R234 B.n309 B.n118 585
R235 B.n311 B.n310 585
R236 B.n312 B.n117 585
R237 B.n314 B.n313 585
R238 B.n315 B.n116 585
R239 B.n317 B.n316 585
R240 B.n318 B.n115 585
R241 B.n320 B.n319 585
R242 B.n321 B.n114 585
R243 B.n323 B.n322 585
R244 B.n324 B.n113 585
R245 B.n326 B.n325 585
R246 B.n327 B.n112 585
R247 B.n329 B.n328 585
R248 B.n330 B.n111 585
R249 B.n332 B.n331 585
R250 B.n333 B.n110 585
R251 B.n335 B.n334 585
R252 B.n336 B.n109 585
R253 B.n338 B.n337 585
R254 B.n339 B.n108 585
R255 B.n341 B.n340 585
R256 B.n342 B.n107 585
R257 B.n344 B.n343 585
R258 B.n345 B.n106 585
R259 B.n347 B.n346 585
R260 B.n348 B.n105 585
R261 B.n350 B.n349 585
R262 B.n351 B.n104 585
R263 B.n353 B.n352 585
R264 B.n354 B.n103 585
R265 B.n356 B.n355 585
R266 B.n357 B.n102 585
R267 B.n359 B.n358 585
R268 B.n360 B.n101 585
R269 B.n362 B.n361 585
R270 B.n363 B.n100 585
R271 B.n365 B.n364 585
R272 B.n366 B.n99 585
R273 B.n368 B.n367 585
R274 B.n369 B.n98 585
R275 B.n371 B.n370 585
R276 B.n372 B.n97 585
R277 B.n200 B.n199 585
R278 B.n198 B.n159 585
R279 B.n197 B.n196 585
R280 B.n195 B.n160 585
R281 B.n194 B.n193 585
R282 B.n192 B.n161 585
R283 B.n191 B.n190 585
R284 B.n189 B.n162 585
R285 B.n188 B.n187 585
R286 B.n186 B.n163 585
R287 B.n185 B.n184 585
R288 B.n183 B.n164 585
R289 B.n182 B.n181 585
R290 B.n180 B.n165 585
R291 B.n179 B.n178 585
R292 B.n177 B.n166 585
R293 B.n176 B.n175 585
R294 B.n174 B.n167 585
R295 B.n173 B.n172 585
R296 B.n171 B.n168 585
R297 B.n170 B.n169 585
R298 B.n2 B.n0 585
R299 B.n645 B.n1 585
R300 B.n644 B.n643 585
R301 B.n642 B.n3 585
R302 B.n641 B.n640 585
R303 B.n639 B.n4 585
R304 B.n638 B.n637 585
R305 B.n636 B.n5 585
R306 B.n635 B.n634 585
R307 B.n633 B.n6 585
R308 B.n632 B.n631 585
R309 B.n630 B.n7 585
R310 B.n629 B.n628 585
R311 B.n627 B.n8 585
R312 B.n626 B.n625 585
R313 B.n624 B.n9 585
R314 B.n623 B.n622 585
R315 B.n621 B.n10 585
R316 B.n620 B.n619 585
R317 B.n618 B.n11 585
R318 B.n617 B.n616 585
R319 B.n615 B.n12 585
R320 B.n614 B.n613 585
R321 B.n647 B.n646 585
R322 B.n201 B.n200 506.916
R323 B.n614 B.n13 506.916
R324 B.n374 B.n97 506.916
R325 B.n441 B.n440 506.916
R326 B.n124 B.t2 462.757
R327 B.n46 B.t4 462.757
R328 B.n130 B.t8 462.757
R329 B.n40 B.t10 462.757
R330 B.n125 B.t1 439.483
R331 B.n47 B.t5 439.483
R332 B.n131 B.t7 439.483
R333 B.n41 B.t11 439.483
R334 B.n200 B.n159 163.367
R335 B.n196 B.n159 163.367
R336 B.n196 B.n195 163.367
R337 B.n195 B.n194 163.367
R338 B.n194 B.n161 163.367
R339 B.n190 B.n161 163.367
R340 B.n190 B.n189 163.367
R341 B.n189 B.n188 163.367
R342 B.n188 B.n163 163.367
R343 B.n184 B.n163 163.367
R344 B.n184 B.n183 163.367
R345 B.n183 B.n182 163.367
R346 B.n182 B.n165 163.367
R347 B.n178 B.n165 163.367
R348 B.n178 B.n177 163.367
R349 B.n177 B.n176 163.367
R350 B.n176 B.n167 163.367
R351 B.n172 B.n167 163.367
R352 B.n172 B.n171 163.367
R353 B.n171 B.n170 163.367
R354 B.n170 B.n2 163.367
R355 B.n646 B.n2 163.367
R356 B.n646 B.n645 163.367
R357 B.n645 B.n644 163.367
R358 B.n644 B.n3 163.367
R359 B.n640 B.n3 163.367
R360 B.n640 B.n639 163.367
R361 B.n639 B.n638 163.367
R362 B.n638 B.n5 163.367
R363 B.n634 B.n5 163.367
R364 B.n634 B.n633 163.367
R365 B.n633 B.n632 163.367
R366 B.n632 B.n7 163.367
R367 B.n628 B.n7 163.367
R368 B.n628 B.n627 163.367
R369 B.n627 B.n626 163.367
R370 B.n626 B.n9 163.367
R371 B.n622 B.n9 163.367
R372 B.n622 B.n621 163.367
R373 B.n621 B.n620 163.367
R374 B.n620 B.n11 163.367
R375 B.n616 B.n11 163.367
R376 B.n616 B.n615 163.367
R377 B.n615 B.n614 163.367
R378 B.n202 B.n201 163.367
R379 B.n202 B.n157 163.367
R380 B.n206 B.n157 163.367
R381 B.n207 B.n206 163.367
R382 B.n208 B.n207 163.367
R383 B.n208 B.n155 163.367
R384 B.n212 B.n155 163.367
R385 B.n213 B.n212 163.367
R386 B.n214 B.n213 163.367
R387 B.n214 B.n153 163.367
R388 B.n218 B.n153 163.367
R389 B.n219 B.n218 163.367
R390 B.n220 B.n219 163.367
R391 B.n220 B.n151 163.367
R392 B.n224 B.n151 163.367
R393 B.n225 B.n224 163.367
R394 B.n226 B.n225 163.367
R395 B.n226 B.n149 163.367
R396 B.n230 B.n149 163.367
R397 B.n231 B.n230 163.367
R398 B.n232 B.n231 163.367
R399 B.n232 B.n147 163.367
R400 B.n236 B.n147 163.367
R401 B.n237 B.n236 163.367
R402 B.n238 B.n237 163.367
R403 B.n238 B.n145 163.367
R404 B.n242 B.n145 163.367
R405 B.n243 B.n242 163.367
R406 B.n244 B.n243 163.367
R407 B.n244 B.n143 163.367
R408 B.n248 B.n143 163.367
R409 B.n249 B.n248 163.367
R410 B.n250 B.n249 163.367
R411 B.n250 B.n141 163.367
R412 B.n254 B.n141 163.367
R413 B.n255 B.n254 163.367
R414 B.n256 B.n255 163.367
R415 B.n256 B.n139 163.367
R416 B.n260 B.n139 163.367
R417 B.n261 B.n260 163.367
R418 B.n262 B.n261 163.367
R419 B.n262 B.n137 163.367
R420 B.n266 B.n137 163.367
R421 B.n267 B.n266 163.367
R422 B.n268 B.n267 163.367
R423 B.n268 B.n135 163.367
R424 B.n272 B.n135 163.367
R425 B.n273 B.n272 163.367
R426 B.n274 B.n273 163.367
R427 B.n274 B.n133 163.367
R428 B.n278 B.n133 163.367
R429 B.n279 B.n278 163.367
R430 B.n279 B.n129 163.367
R431 B.n283 B.n129 163.367
R432 B.n284 B.n283 163.367
R433 B.n285 B.n284 163.367
R434 B.n285 B.n127 163.367
R435 B.n289 B.n127 163.367
R436 B.n290 B.n289 163.367
R437 B.n291 B.n290 163.367
R438 B.n291 B.n123 163.367
R439 B.n296 B.n123 163.367
R440 B.n297 B.n296 163.367
R441 B.n298 B.n297 163.367
R442 B.n298 B.n121 163.367
R443 B.n302 B.n121 163.367
R444 B.n303 B.n302 163.367
R445 B.n304 B.n303 163.367
R446 B.n304 B.n119 163.367
R447 B.n308 B.n119 163.367
R448 B.n309 B.n308 163.367
R449 B.n310 B.n309 163.367
R450 B.n310 B.n117 163.367
R451 B.n314 B.n117 163.367
R452 B.n315 B.n314 163.367
R453 B.n316 B.n315 163.367
R454 B.n316 B.n115 163.367
R455 B.n320 B.n115 163.367
R456 B.n321 B.n320 163.367
R457 B.n322 B.n321 163.367
R458 B.n322 B.n113 163.367
R459 B.n326 B.n113 163.367
R460 B.n327 B.n326 163.367
R461 B.n328 B.n327 163.367
R462 B.n328 B.n111 163.367
R463 B.n332 B.n111 163.367
R464 B.n333 B.n332 163.367
R465 B.n334 B.n333 163.367
R466 B.n334 B.n109 163.367
R467 B.n338 B.n109 163.367
R468 B.n339 B.n338 163.367
R469 B.n340 B.n339 163.367
R470 B.n340 B.n107 163.367
R471 B.n344 B.n107 163.367
R472 B.n345 B.n344 163.367
R473 B.n346 B.n345 163.367
R474 B.n346 B.n105 163.367
R475 B.n350 B.n105 163.367
R476 B.n351 B.n350 163.367
R477 B.n352 B.n351 163.367
R478 B.n352 B.n103 163.367
R479 B.n356 B.n103 163.367
R480 B.n357 B.n356 163.367
R481 B.n358 B.n357 163.367
R482 B.n358 B.n101 163.367
R483 B.n362 B.n101 163.367
R484 B.n363 B.n362 163.367
R485 B.n364 B.n363 163.367
R486 B.n364 B.n99 163.367
R487 B.n368 B.n99 163.367
R488 B.n369 B.n368 163.367
R489 B.n370 B.n369 163.367
R490 B.n370 B.n97 163.367
R491 B.n375 B.n374 163.367
R492 B.n376 B.n375 163.367
R493 B.n376 B.n95 163.367
R494 B.n380 B.n95 163.367
R495 B.n381 B.n380 163.367
R496 B.n382 B.n381 163.367
R497 B.n382 B.n93 163.367
R498 B.n386 B.n93 163.367
R499 B.n387 B.n386 163.367
R500 B.n388 B.n387 163.367
R501 B.n388 B.n91 163.367
R502 B.n392 B.n91 163.367
R503 B.n393 B.n392 163.367
R504 B.n394 B.n393 163.367
R505 B.n394 B.n89 163.367
R506 B.n398 B.n89 163.367
R507 B.n399 B.n398 163.367
R508 B.n400 B.n399 163.367
R509 B.n400 B.n87 163.367
R510 B.n404 B.n87 163.367
R511 B.n405 B.n404 163.367
R512 B.n406 B.n405 163.367
R513 B.n406 B.n85 163.367
R514 B.n410 B.n85 163.367
R515 B.n411 B.n410 163.367
R516 B.n412 B.n411 163.367
R517 B.n412 B.n83 163.367
R518 B.n416 B.n83 163.367
R519 B.n417 B.n416 163.367
R520 B.n418 B.n417 163.367
R521 B.n418 B.n81 163.367
R522 B.n422 B.n81 163.367
R523 B.n423 B.n422 163.367
R524 B.n424 B.n423 163.367
R525 B.n424 B.n79 163.367
R526 B.n428 B.n79 163.367
R527 B.n429 B.n428 163.367
R528 B.n430 B.n429 163.367
R529 B.n430 B.n77 163.367
R530 B.n434 B.n77 163.367
R531 B.n435 B.n434 163.367
R532 B.n436 B.n435 163.367
R533 B.n436 B.n75 163.367
R534 B.n440 B.n75 163.367
R535 B.n610 B.n13 163.367
R536 B.n610 B.n609 163.367
R537 B.n609 B.n608 163.367
R538 B.n608 B.n15 163.367
R539 B.n604 B.n15 163.367
R540 B.n604 B.n603 163.367
R541 B.n603 B.n602 163.367
R542 B.n602 B.n17 163.367
R543 B.n598 B.n17 163.367
R544 B.n598 B.n597 163.367
R545 B.n597 B.n596 163.367
R546 B.n596 B.n19 163.367
R547 B.n592 B.n19 163.367
R548 B.n592 B.n591 163.367
R549 B.n591 B.n590 163.367
R550 B.n590 B.n21 163.367
R551 B.n586 B.n21 163.367
R552 B.n586 B.n585 163.367
R553 B.n585 B.n584 163.367
R554 B.n584 B.n23 163.367
R555 B.n580 B.n23 163.367
R556 B.n580 B.n579 163.367
R557 B.n579 B.n578 163.367
R558 B.n578 B.n25 163.367
R559 B.n574 B.n25 163.367
R560 B.n574 B.n573 163.367
R561 B.n573 B.n572 163.367
R562 B.n572 B.n27 163.367
R563 B.n568 B.n27 163.367
R564 B.n568 B.n567 163.367
R565 B.n567 B.n566 163.367
R566 B.n566 B.n29 163.367
R567 B.n562 B.n29 163.367
R568 B.n562 B.n561 163.367
R569 B.n561 B.n560 163.367
R570 B.n560 B.n31 163.367
R571 B.n556 B.n31 163.367
R572 B.n556 B.n555 163.367
R573 B.n555 B.n554 163.367
R574 B.n554 B.n33 163.367
R575 B.n550 B.n33 163.367
R576 B.n550 B.n549 163.367
R577 B.n549 B.n548 163.367
R578 B.n548 B.n35 163.367
R579 B.n544 B.n35 163.367
R580 B.n544 B.n543 163.367
R581 B.n543 B.n542 163.367
R582 B.n542 B.n37 163.367
R583 B.n538 B.n37 163.367
R584 B.n538 B.n537 163.367
R585 B.n537 B.n536 163.367
R586 B.n536 B.n39 163.367
R587 B.n531 B.n39 163.367
R588 B.n531 B.n530 163.367
R589 B.n530 B.n529 163.367
R590 B.n529 B.n43 163.367
R591 B.n525 B.n43 163.367
R592 B.n525 B.n524 163.367
R593 B.n524 B.n523 163.367
R594 B.n523 B.n45 163.367
R595 B.n519 B.n45 163.367
R596 B.n519 B.n518 163.367
R597 B.n518 B.n49 163.367
R598 B.n514 B.n49 163.367
R599 B.n514 B.n513 163.367
R600 B.n513 B.n512 163.367
R601 B.n512 B.n51 163.367
R602 B.n508 B.n51 163.367
R603 B.n508 B.n507 163.367
R604 B.n507 B.n506 163.367
R605 B.n506 B.n53 163.367
R606 B.n502 B.n53 163.367
R607 B.n502 B.n501 163.367
R608 B.n501 B.n500 163.367
R609 B.n500 B.n55 163.367
R610 B.n496 B.n55 163.367
R611 B.n496 B.n495 163.367
R612 B.n495 B.n494 163.367
R613 B.n494 B.n57 163.367
R614 B.n490 B.n57 163.367
R615 B.n490 B.n489 163.367
R616 B.n489 B.n488 163.367
R617 B.n488 B.n59 163.367
R618 B.n484 B.n59 163.367
R619 B.n484 B.n483 163.367
R620 B.n483 B.n482 163.367
R621 B.n482 B.n61 163.367
R622 B.n478 B.n61 163.367
R623 B.n478 B.n477 163.367
R624 B.n477 B.n476 163.367
R625 B.n476 B.n63 163.367
R626 B.n472 B.n63 163.367
R627 B.n472 B.n471 163.367
R628 B.n471 B.n470 163.367
R629 B.n470 B.n65 163.367
R630 B.n466 B.n65 163.367
R631 B.n466 B.n465 163.367
R632 B.n465 B.n464 163.367
R633 B.n464 B.n67 163.367
R634 B.n460 B.n67 163.367
R635 B.n460 B.n459 163.367
R636 B.n459 B.n458 163.367
R637 B.n458 B.n69 163.367
R638 B.n454 B.n69 163.367
R639 B.n454 B.n453 163.367
R640 B.n453 B.n452 163.367
R641 B.n452 B.n71 163.367
R642 B.n448 B.n71 163.367
R643 B.n448 B.n447 163.367
R644 B.n447 B.n446 163.367
R645 B.n446 B.n73 163.367
R646 B.n442 B.n73 163.367
R647 B.n442 B.n441 163.367
R648 B.n294 B.n125 59.5399
R649 B.n132 B.n131 59.5399
R650 B.n534 B.n41 59.5399
R651 B.n48 B.n47 59.5399
R652 B.n613 B.n612 32.9371
R653 B.n439 B.n74 32.9371
R654 B.n373 B.n372 32.9371
R655 B.n199 B.n158 32.9371
R656 B.n125 B.n124 23.2732
R657 B.n131 B.n130 23.2732
R658 B.n41 B.n40 23.2732
R659 B.n47 B.n46 23.2732
R660 B B.n647 18.0485
R661 B.n612 B.n611 10.6151
R662 B.n611 B.n14 10.6151
R663 B.n607 B.n14 10.6151
R664 B.n607 B.n606 10.6151
R665 B.n606 B.n605 10.6151
R666 B.n605 B.n16 10.6151
R667 B.n601 B.n16 10.6151
R668 B.n601 B.n600 10.6151
R669 B.n600 B.n599 10.6151
R670 B.n599 B.n18 10.6151
R671 B.n595 B.n18 10.6151
R672 B.n595 B.n594 10.6151
R673 B.n594 B.n593 10.6151
R674 B.n593 B.n20 10.6151
R675 B.n589 B.n20 10.6151
R676 B.n589 B.n588 10.6151
R677 B.n588 B.n587 10.6151
R678 B.n587 B.n22 10.6151
R679 B.n583 B.n22 10.6151
R680 B.n583 B.n582 10.6151
R681 B.n582 B.n581 10.6151
R682 B.n581 B.n24 10.6151
R683 B.n577 B.n24 10.6151
R684 B.n577 B.n576 10.6151
R685 B.n576 B.n575 10.6151
R686 B.n575 B.n26 10.6151
R687 B.n571 B.n26 10.6151
R688 B.n571 B.n570 10.6151
R689 B.n570 B.n569 10.6151
R690 B.n569 B.n28 10.6151
R691 B.n565 B.n28 10.6151
R692 B.n565 B.n564 10.6151
R693 B.n564 B.n563 10.6151
R694 B.n563 B.n30 10.6151
R695 B.n559 B.n30 10.6151
R696 B.n559 B.n558 10.6151
R697 B.n558 B.n557 10.6151
R698 B.n557 B.n32 10.6151
R699 B.n553 B.n32 10.6151
R700 B.n553 B.n552 10.6151
R701 B.n552 B.n551 10.6151
R702 B.n551 B.n34 10.6151
R703 B.n547 B.n34 10.6151
R704 B.n547 B.n546 10.6151
R705 B.n546 B.n545 10.6151
R706 B.n545 B.n36 10.6151
R707 B.n541 B.n36 10.6151
R708 B.n541 B.n540 10.6151
R709 B.n540 B.n539 10.6151
R710 B.n539 B.n38 10.6151
R711 B.n535 B.n38 10.6151
R712 B.n533 B.n532 10.6151
R713 B.n532 B.n42 10.6151
R714 B.n528 B.n42 10.6151
R715 B.n528 B.n527 10.6151
R716 B.n527 B.n526 10.6151
R717 B.n526 B.n44 10.6151
R718 B.n522 B.n44 10.6151
R719 B.n522 B.n521 10.6151
R720 B.n521 B.n520 10.6151
R721 B.n517 B.n516 10.6151
R722 B.n516 B.n515 10.6151
R723 B.n515 B.n50 10.6151
R724 B.n511 B.n50 10.6151
R725 B.n511 B.n510 10.6151
R726 B.n510 B.n509 10.6151
R727 B.n509 B.n52 10.6151
R728 B.n505 B.n52 10.6151
R729 B.n505 B.n504 10.6151
R730 B.n504 B.n503 10.6151
R731 B.n503 B.n54 10.6151
R732 B.n499 B.n54 10.6151
R733 B.n499 B.n498 10.6151
R734 B.n498 B.n497 10.6151
R735 B.n497 B.n56 10.6151
R736 B.n493 B.n56 10.6151
R737 B.n493 B.n492 10.6151
R738 B.n492 B.n491 10.6151
R739 B.n491 B.n58 10.6151
R740 B.n487 B.n58 10.6151
R741 B.n487 B.n486 10.6151
R742 B.n486 B.n485 10.6151
R743 B.n485 B.n60 10.6151
R744 B.n481 B.n60 10.6151
R745 B.n481 B.n480 10.6151
R746 B.n480 B.n479 10.6151
R747 B.n479 B.n62 10.6151
R748 B.n475 B.n62 10.6151
R749 B.n475 B.n474 10.6151
R750 B.n474 B.n473 10.6151
R751 B.n473 B.n64 10.6151
R752 B.n469 B.n64 10.6151
R753 B.n469 B.n468 10.6151
R754 B.n468 B.n467 10.6151
R755 B.n467 B.n66 10.6151
R756 B.n463 B.n66 10.6151
R757 B.n463 B.n462 10.6151
R758 B.n462 B.n461 10.6151
R759 B.n461 B.n68 10.6151
R760 B.n457 B.n68 10.6151
R761 B.n457 B.n456 10.6151
R762 B.n456 B.n455 10.6151
R763 B.n455 B.n70 10.6151
R764 B.n451 B.n70 10.6151
R765 B.n451 B.n450 10.6151
R766 B.n450 B.n449 10.6151
R767 B.n449 B.n72 10.6151
R768 B.n445 B.n72 10.6151
R769 B.n445 B.n444 10.6151
R770 B.n444 B.n443 10.6151
R771 B.n443 B.n74 10.6151
R772 B.n373 B.n96 10.6151
R773 B.n377 B.n96 10.6151
R774 B.n378 B.n377 10.6151
R775 B.n379 B.n378 10.6151
R776 B.n379 B.n94 10.6151
R777 B.n383 B.n94 10.6151
R778 B.n384 B.n383 10.6151
R779 B.n385 B.n384 10.6151
R780 B.n385 B.n92 10.6151
R781 B.n389 B.n92 10.6151
R782 B.n390 B.n389 10.6151
R783 B.n391 B.n390 10.6151
R784 B.n391 B.n90 10.6151
R785 B.n395 B.n90 10.6151
R786 B.n396 B.n395 10.6151
R787 B.n397 B.n396 10.6151
R788 B.n397 B.n88 10.6151
R789 B.n401 B.n88 10.6151
R790 B.n402 B.n401 10.6151
R791 B.n403 B.n402 10.6151
R792 B.n403 B.n86 10.6151
R793 B.n407 B.n86 10.6151
R794 B.n408 B.n407 10.6151
R795 B.n409 B.n408 10.6151
R796 B.n409 B.n84 10.6151
R797 B.n413 B.n84 10.6151
R798 B.n414 B.n413 10.6151
R799 B.n415 B.n414 10.6151
R800 B.n415 B.n82 10.6151
R801 B.n419 B.n82 10.6151
R802 B.n420 B.n419 10.6151
R803 B.n421 B.n420 10.6151
R804 B.n421 B.n80 10.6151
R805 B.n425 B.n80 10.6151
R806 B.n426 B.n425 10.6151
R807 B.n427 B.n426 10.6151
R808 B.n427 B.n78 10.6151
R809 B.n431 B.n78 10.6151
R810 B.n432 B.n431 10.6151
R811 B.n433 B.n432 10.6151
R812 B.n433 B.n76 10.6151
R813 B.n437 B.n76 10.6151
R814 B.n438 B.n437 10.6151
R815 B.n439 B.n438 10.6151
R816 B.n203 B.n158 10.6151
R817 B.n204 B.n203 10.6151
R818 B.n205 B.n204 10.6151
R819 B.n205 B.n156 10.6151
R820 B.n209 B.n156 10.6151
R821 B.n210 B.n209 10.6151
R822 B.n211 B.n210 10.6151
R823 B.n211 B.n154 10.6151
R824 B.n215 B.n154 10.6151
R825 B.n216 B.n215 10.6151
R826 B.n217 B.n216 10.6151
R827 B.n217 B.n152 10.6151
R828 B.n221 B.n152 10.6151
R829 B.n222 B.n221 10.6151
R830 B.n223 B.n222 10.6151
R831 B.n223 B.n150 10.6151
R832 B.n227 B.n150 10.6151
R833 B.n228 B.n227 10.6151
R834 B.n229 B.n228 10.6151
R835 B.n229 B.n148 10.6151
R836 B.n233 B.n148 10.6151
R837 B.n234 B.n233 10.6151
R838 B.n235 B.n234 10.6151
R839 B.n235 B.n146 10.6151
R840 B.n239 B.n146 10.6151
R841 B.n240 B.n239 10.6151
R842 B.n241 B.n240 10.6151
R843 B.n241 B.n144 10.6151
R844 B.n245 B.n144 10.6151
R845 B.n246 B.n245 10.6151
R846 B.n247 B.n246 10.6151
R847 B.n247 B.n142 10.6151
R848 B.n251 B.n142 10.6151
R849 B.n252 B.n251 10.6151
R850 B.n253 B.n252 10.6151
R851 B.n253 B.n140 10.6151
R852 B.n257 B.n140 10.6151
R853 B.n258 B.n257 10.6151
R854 B.n259 B.n258 10.6151
R855 B.n259 B.n138 10.6151
R856 B.n263 B.n138 10.6151
R857 B.n264 B.n263 10.6151
R858 B.n265 B.n264 10.6151
R859 B.n265 B.n136 10.6151
R860 B.n269 B.n136 10.6151
R861 B.n270 B.n269 10.6151
R862 B.n271 B.n270 10.6151
R863 B.n271 B.n134 10.6151
R864 B.n275 B.n134 10.6151
R865 B.n276 B.n275 10.6151
R866 B.n277 B.n276 10.6151
R867 B.n281 B.n280 10.6151
R868 B.n282 B.n281 10.6151
R869 B.n282 B.n128 10.6151
R870 B.n286 B.n128 10.6151
R871 B.n287 B.n286 10.6151
R872 B.n288 B.n287 10.6151
R873 B.n288 B.n126 10.6151
R874 B.n292 B.n126 10.6151
R875 B.n293 B.n292 10.6151
R876 B.n295 B.n122 10.6151
R877 B.n299 B.n122 10.6151
R878 B.n300 B.n299 10.6151
R879 B.n301 B.n300 10.6151
R880 B.n301 B.n120 10.6151
R881 B.n305 B.n120 10.6151
R882 B.n306 B.n305 10.6151
R883 B.n307 B.n306 10.6151
R884 B.n307 B.n118 10.6151
R885 B.n311 B.n118 10.6151
R886 B.n312 B.n311 10.6151
R887 B.n313 B.n312 10.6151
R888 B.n313 B.n116 10.6151
R889 B.n317 B.n116 10.6151
R890 B.n318 B.n317 10.6151
R891 B.n319 B.n318 10.6151
R892 B.n319 B.n114 10.6151
R893 B.n323 B.n114 10.6151
R894 B.n324 B.n323 10.6151
R895 B.n325 B.n324 10.6151
R896 B.n325 B.n112 10.6151
R897 B.n329 B.n112 10.6151
R898 B.n330 B.n329 10.6151
R899 B.n331 B.n330 10.6151
R900 B.n331 B.n110 10.6151
R901 B.n335 B.n110 10.6151
R902 B.n336 B.n335 10.6151
R903 B.n337 B.n336 10.6151
R904 B.n337 B.n108 10.6151
R905 B.n341 B.n108 10.6151
R906 B.n342 B.n341 10.6151
R907 B.n343 B.n342 10.6151
R908 B.n343 B.n106 10.6151
R909 B.n347 B.n106 10.6151
R910 B.n348 B.n347 10.6151
R911 B.n349 B.n348 10.6151
R912 B.n349 B.n104 10.6151
R913 B.n353 B.n104 10.6151
R914 B.n354 B.n353 10.6151
R915 B.n355 B.n354 10.6151
R916 B.n355 B.n102 10.6151
R917 B.n359 B.n102 10.6151
R918 B.n360 B.n359 10.6151
R919 B.n361 B.n360 10.6151
R920 B.n361 B.n100 10.6151
R921 B.n365 B.n100 10.6151
R922 B.n366 B.n365 10.6151
R923 B.n367 B.n366 10.6151
R924 B.n367 B.n98 10.6151
R925 B.n371 B.n98 10.6151
R926 B.n372 B.n371 10.6151
R927 B.n199 B.n198 10.6151
R928 B.n198 B.n197 10.6151
R929 B.n197 B.n160 10.6151
R930 B.n193 B.n160 10.6151
R931 B.n193 B.n192 10.6151
R932 B.n192 B.n191 10.6151
R933 B.n191 B.n162 10.6151
R934 B.n187 B.n162 10.6151
R935 B.n187 B.n186 10.6151
R936 B.n186 B.n185 10.6151
R937 B.n185 B.n164 10.6151
R938 B.n181 B.n164 10.6151
R939 B.n181 B.n180 10.6151
R940 B.n180 B.n179 10.6151
R941 B.n179 B.n166 10.6151
R942 B.n175 B.n166 10.6151
R943 B.n175 B.n174 10.6151
R944 B.n174 B.n173 10.6151
R945 B.n173 B.n168 10.6151
R946 B.n169 B.n168 10.6151
R947 B.n169 B.n0 10.6151
R948 B.n643 B.n1 10.6151
R949 B.n643 B.n642 10.6151
R950 B.n642 B.n641 10.6151
R951 B.n641 B.n4 10.6151
R952 B.n637 B.n4 10.6151
R953 B.n637 B.n636 10.6151
R954 B.n636 B.n635 10.6151
R955 B.n635 B.n6 10.6151
R956 B.n631 B.n6 10.6151
R957 B.n631 B.n630 10.6151
R958 B.n630 B.n629 10.6151
R959 B.n629 B.n8 10.6151
R960 B.n625 B.n8 10.6151
R961 B.n625 B.n624 10.6151
R962 B.n624 B.n623 10.6151
R963 B.n623 B.n10 10.6151
R964 B.n619 B.n10 10.6151
R965 B.n619 B.n618 10.6151
R966 B.n618 B.n617 10.6151
R967 B.n617 B.n12 10.6151
R968 B.n613 B.n12 10.6151
R969 B.n535 B.n534 9.36635
R970 B.n517 B.n48 9.36635
R971 B.n277 B.n132 9.36635
R972 B.n295 B.n294 9.36635
R973 B.n647 B.n0 2.81026
R974 B.n647 B.n1 2.81026
R975 B.n534 B.n533 1.24928
R976 B.n520 B.n48 1.24928
R977 B.n280 B.n132 1.24928
R978 B.n294 B.n293 1.24928
R979 VP.n5 VP.t1 491.878
R980 VP.n12 VP.t3 475.63
R981 VP.n19 VP.t2 475.63
R982 VP.n9 VP.t5 475.63
R983 VP.n1 VP.t0 430.476
R984 VP.n4 VP.t4 430.476
R985 VP.n20 VP.n19 161.3
R986 VP.n7 VP.n6 161.3
R987 VP.n8 VP.n3 161.3
R988 VP.n10 VP.n9 161.3
R989 VP.n18 VP.n0 161.3
R990 VP.n17 VP.n16 161.3
R991 VP.n15 VP.n14 161.3
R992 VP.n13 VP.n2 161.3
R993 VP.n12 VP.n11 161.3
R994 VP.n14 VP.n13 55.1086
R995 VP.n18 VP.n17 55.1086
R996 VP.n8 VP.n7 55.1086
R997 VP.n11 VP.n10 44.5308
R998 VP.n6 VP.n5 43.7016
R999 VP.n5 VP.n4 42.7308
R1000 VP.n14 VP.n1 12.2964
R1001 VP.n17 VP.n1 12.2964
R1002 VP.n7 VP.n4 12.2964
R1003 VP.n13 VP.n12 2.19141
R1004 VP.n19 VP.n18 2.19141
R1005 VP.n9 VP.n8 2.19141
R1006 VP.n6 VP.n3 0.189894
R1007 VP.n10 VP.n3 0.189894
R1008 VP.n11 VP.n2 0.189894
R1009 VP.n15 VP.n2 0.189894
R1010 VP.n16 VP.n15 0.189894
R1011 VP.n16 VP.n0 0.189894
R1012 VP.n20 VP.n0 0.189894
R1013 VP VP.n20 0.0516364
R1014 VDD1.n80 VDD1.n0 756.745
R1015 VDD1.n165 VDD1.n85 756.745
R1016 VDD1.n81 VDD1.n80 585
R1017 VDD1.n79 VDD1.n78 585
R1018 VDD1.n4 VDD1.n3 585
R1019 VDD1.n8 VDD1.n6 585
R1020 VDD1.n73 VDD1.n72 585
R1021 VDD1.n71 VDD1.n70 585
R1022 VDD1.n10 VDD1.n9 585
R1023 VDD1.n65 VDD1.n64 585
R1024 VDD1.n63 VDD1.n62 585
R1025 VDD1.n14 VDD1.n13 585
R1026 VDD1.n57 VDD1.n56 585
R1027 VDD1.n55 VDD1.n54 585
R1028 VDD1.n18 VDD1.n17 585
R1029 VDD1.n49 VDD1.n48 585
R1030 VDD1.n47 VDD1.n46 585
R1031 VDD1.n22 VDD1.n21 585
R1032 VDD1.n41 VDD1.n40 585
R1033 VDD1.n39 VDD1.n38 585
R1034 VDD1.n26 VDD1.n25 585
R1035 VDD1.n33 VDD1.n32 585
R1036 VDD1.n31 VDD1.n30 585
R1037 VDD1.n114 VDD1.n113 585
R1038 VDD1.n116 VDD1.n115 585
R1039 VDD1.n109 VDD1.n108 585
R1040 VDD1.n122 VDD1.n121 585
R1041 VDD1.n124 VDD1.n123 585
R1042 VDD1.n105 VDD1.n104 585
R1043 VDD1.n130 VDD1.n129 585
R1044 VDD1.n132 VDD1.n131 585
R1045 VDD1.n101 VDD1.n100 585
R1046 VDD1.n138 VDD1.n137 585
R1047 VDD1.n140 VDD1.n139 585
R1048 VDD1.n97 VDD1.n96 585
R1049 VDD1.n146 VDD1.n145 585
R1050 VDD1.n148 VDD1.n147 585
R1051 VDD1.n93 VDD1.n92 585
R1052 VDD1.n155 VDD1.n154 585
R1053 VDD1.n156 VDD1.n91 585
R1054 VDD1.n158 VDD1.n157 585
R1055 VDD1.n89 VDD1.n88 585
R1056 VDD1.n164 VDD1.n163 585
R1057 VDD1.n166 VDD1.n165 585
R1058 VDD1.n29 VDD1.t0 327.466
R1059 VDD1.n112 VDD1.t4 327.466
R1060 VDD1.n80 VDD1.n79 171.744
R1061 VDD1.n79 VDD1.n3 171.744
R1062 VDD1.n8 VDD1.n3 171.744
R1063 VDD1.n72 VDD1.n8 171.744
R1064 VDD1.n72 VDD1.n71 171.744
R1065 VDD1.n71 VDD1.n9 171.744
R1066 VDD1.n64 VDD1.n9 171.744
R1067 VDD1.n64 VDD1.n63 171.744
R1068 VDD1.n63 VDD1.n13 171.744
R1069 VDD1.n56 VDD1.n13 171.744
R1070 VDD1.n56 VDD1.n55 171.744
R1071 VDD1.n55 VDD1.n17 171.744
R1072 VDD1.n48 VDD1.n17 171.744
R1073 VDD1.n48 VDD1.n47 171.744
R1074 VDD1.n47 VDD1.n21 171.744
R1075 VDD1.n40 VDD1.n21 171.744
R1076 VDD1.n40 VDD1.n39 171.744
R1077 VDD1.n39 VDD1.n25 171.744
R1078 VDD1.n32 VDD1.n25 171.744
R1079 VDD1.n32 VDD1.n31 171.744
R1080 VDD1.n115 VDD1.n114 171.744
R1081 VDD1.n115 VDD1.n108 171.744
R1082 VDD1.n122 VDD1.n108 171.744
R1083 VDD1.n123 VDD1.n122 171.744
R1084 VDD1.n123 VDD1.n104 171.744
R1085 VDD1.n130 VDD1.n104 171.744
R1086 VDD1.n131 VDD1.n130 171.744
R1087 VDD1.n131 VDD1.n100 171.744
R1088 VDD1.n138 VDD1.n100 171.744
R1089 VDD1.n139 VDD1.n138 171.744
R1090 VDD1.n139 VDD1.n96 171.744
R1091 VDD1.n146 VDD1.n96 171.744
R1092 VDD1.n147 VDD1.n146 171.744
R1093 VDD1.n147 VDD1.n92 171.744
R1094 VDD1.n155 VDD1.n92 171.744
R1095 VDD1.n156 VDD1.n155 171.744
R1096 VDD1.n157 VDD1.n156 171.744
R1097 VDD1.n157 VDD1.n88 171.744
R1098 VDD1.n164 VDD1.n88 171.744
R1099 VDD1.n165 VDD1.n164 171.744
R1100 VDD1.n31 VDD1.t0 85.8723
R1101 VDD1.n114 VDD1.t4 85.8723
R1102 VDD1.n171 VDD1.n170 73.9521
R1103 VDD1.n173 VDD1.n172 73.7489
R1104 VDD1 VDD1.n84 53.1891
R1105 VDD1.n171 VDD1.n169 53.0756
R1106 VDD1.n173 VDD1.n171 41.5742
R1107 VDD1.n30 VDD1.n29 16.3895
R1108 VDD1.n113 VDD1.n112 16.3895
R1109 VDD1.n6 VDD1.n4 13.1884
R1110 VDD1.n158 VDD1.n89 13.1884
R1111 VDD1.n78 VDD1.n77 12.8005
R1112 VDD1.n74 VDD1.n73 12.8005
R1113 VDD1.n33 VDD1.n28 12.8005
R1114 VDD1.n116 VDD1.n111 12.8005
R1115 VDD1.n159 VDD1.n91 12.8005
R1116 VDD1.n163 VDD1.n162 12.8005
R1117 VDD1.n81 VDD1.n2 12.0247
R1118 VDD1.n70 VDD1.n7 12.0247
R1119 VDD1.n34 VDD1.n26 12.0247
R1120 VDD1.n117 VDD1.n109 12.0247
R1121 VDD1.n154 VDD1.n153 12.0247
R1122 VDD1.n166 VDD1.n87 12.0247
R1123 VDD1.n82 VDD1.n0 11.249
R1124 VDD1.n69 VDD1.n10 11.249
R1125 VDD1.n38 VDD1.n37 11.249
R1126 VDD1.n121 VDD1.n120 11.249
R1127 VDD1.n152 VDD1.n93 11.249
R1128 VDD1.n167 VDD1.n85 11.249
R1129 VDD1.n66 VDD1.n65 10.4732
R1130 VDD1.n41 VDD1.n24 10.4732
R1131 VDD1.n124 VDD1.n107 10.4732
R1132 VDD1.n149 VDD1.n148 10.4732
R1133 VDD1.n62 VDD1.n12 9.69747
R1134 VDD1.n42 VDD1.n22 9.69747
R1135 VDD1.n125 VDD1.n105 9.69747
R1136 VDD1.n145 VDD1.n95 9.69747
R1137 VDD1.n84 VDD1.n83 9.45567
R1138 VDD1.n169 VDD1.n168 9.45567
R1139 VDD1.n16 VDD1.n15 9.3005
R1140 VDD1.n59 VDD1.n58 9.3005
R1141 VDD1.n61 VDD1.n60 9.3005
R1142 VDD1.n12 VDD1.n11 9.3005
R1143 VDD1.n67 VDD1.n66 9.3005
R1144 VDD1.n69 VDD1.n68 9.3005
R1145 VDD1.n7 VDD1.n5 9.3005
R1146 VDD1.n75 VDD1.n74 9.3005
R1147 VDD1.n83 VDD1.n82 9.3005
R1148 VDD1.n2 VDD1.n1 9.3005
R1149 VDD1.n77 VDD1.n76 9.3005
R1150 VDD1.n53 VDD1.n52 9.3005
R1151 VDD1.n51 VDD1.n50 9.3005
R1152 VDD1.n20 VDD1.n19 9.3005
R1153 VDD1.n45 VDD1.n44 9.3005
R1154 VDD1.n43 VDD1.n42 9.3005
R1155 VDD1.n24 VDD1.n23 9.3005
R1156 VDD1.n37 VDD1.n36 9.3005
R1157 VDD1.n35 VDD1.n34 9.3005
R1158 VDD1.n28 VDD1.n27 9.3005
R1159 VDD1.n168 VDD1.n167 9.3005
R1160 VDD1.n87 VDD1.n86 9.3005
R1161 VDD1.n162 VDD1.n161 9.3005
R1162 VDD1.n134 VDD1.n133 9.3005
R1163 VDD1.n103 VDD1.n102 9.3005
R1164 VDD1.n128 VDD1.n127 9.3005
R1165 VDD1.n126 VDD1.n125 9.3005
R1166 VDD1.n107 VDD1.n106 9.3005
R1167 VDD1.n120 VDD1.n119 9.3005
R1168 VDD1.n118 VDD1.n117 9.3005
R1169 VDD1.n111 VDD1.n110 9.3005
R1170 VDD1.n136 VDD1.n135 9.3005
R1171 VDD1.n99 VDD1.n98 9.3005
R1172 VDD1.n142 VDD1.n141 9.3005
R1173 VDD1.n144 VDD1.n143 9.3005
R1174 VDD1.n95 VDD1.n94 9.3005
R1175 VDD1.n150 VDD1.n149 9.3005
R1176 VDD1.n152 VDD1.n151 9.3005
R1177 VDD1.n153 VDD1.n90 9.3005
R1178 VDD1.n160 VDD1.n159 9.3005
R1179 VDD1.n61 VDD1.n14 8.92171
R1180 VDD1.n46 VDD1.n45 8.92171
R1181 VDD1.n129 VDD1.n128 8.92171
R1182 VDD1.n144 VDD1.n97 8.92171
R1183 VDD1.n58 VDD1.n57 8.14595
R1184 VDD1.n49 VDD1.n20 8.14595
R1185 VDD1.n132 VDD1.n103 8.14595
R1186 VDD1.n141 VDD1.n140 8.14595
R1187 VDD1.n54 VDD1.n16 7.3702
R1188 VDD1.n50 VDD1.n18 7.3702
R1189 VDD1.n133 VDD1.n101 7.3702
R1190 VDD1.n137 VDD1.n99 7.3702
R1191 VDD1.n54 VDD1.n53 6.59444
R1192 VDD1.n53 VDD1.n18 6.59444
R1193 VDD1.n136 VDD1.n101 6.59444
R1194 VDD1.n137 VDD1.n136 6.59444
R1195 VDD1.n57 VDD1.n16 5.81868
R1196 VDD1.n50 VDD1.n49 5.81868
R1197 VDD1.n133 VDD1.n132 5.81868
R1198 VDD1.n140 VDD1.n99 5.81868
R1199 VDD1.n58 VDD1.n14 5.04292
R1200 VDD1.n46 VDD1.n20 5.04292
R1201 VDD1.n129 VDD1.n103 5.04292
R1202 VDD1.n141 VDD1.n97 5.04292
R1203 VDD1.n62 VDD1.n61 4.26717
R1204 VDD1.n45 VDD1.n22 4.26717
R1205 VDD1.n128 VDD1.n105 4.26717
R1206 VDD1.n145 VDD1.n144 4.26717
R1207 VDD1.n29 VDD1.n27 3.70982
R1208 VDD1.n112 VDD1.n110 3.70982
R1209 VDD1.n65 VDD1.n12 3.49141
R1210 VDD1.n42 VDD1.n41 3.49141
R1211 VDD1.n125 VDD1.n124 3.49141
R1212 VDD1.n148 VDD1.n95 3.49141
R1213 VDD1.n84 VDD1.n0 2.71565
R1214 VDD1.n66 VDD1.n10 2.71565
R1215 VDD1.n38 VDD1.n24 2.71565
R1216 VDD1.n121 VDD1.n107 2.71565
R1217 VDD1.n149 VDD1.n93 2.71565
R1218 VDD1.n169 VDD1.n85 2.71565
R1219 VDD1.n172 VDD1.t3 2.0922
R1220 VDD1.n172 VDD1.t2 2.0922
R1221 VDD1.n170 VDD1.t1 2.0922
R1222 VDD1.n170 VDD1.t5 2.0922
R1223 VDD1.n82 VDD1.n81 1.93989
R1224 VDD1.n70 VDD1.n69 1.93989
R1225 VDD1.n37 VDD1.n26 1.93989
R1226 VDD1.n120 VDD1.n109 1.93989
R1227 VDD1.n154 VDD1.n152 1.93989
R1228 VDD1.n167 VDD1.n166 1.93989
R1229 VDD1.n78 VDD1.n2 1.16414
R1230 VDD1.n73 VDD1.n7 1.16414
R1231 VDD1.n34 VDD1.n33 1.16414
R1232 VDD1.n117 VDD1.n116 1.16414
R1233 VDD1.n153 VDD1.n91 1.16414
R1234 VDD1.n163 VDD1.n87 1.16414
R1235 VDD1.n77 VDD1.n4 0.388379
R1236 VDD1.n74 VDD1.n6 0.388379
R1237 VDD1.n30 VDD1.n28 0.388379
R1238 VDD1.n113 VDD1.n111 0.388379
R1239 VDD1.n159 VDD1.n158 0.388379
R1240 VDD1.n162 VDD1.n89 0.388379
R1241 VDD1 VDD1.n173 0.200931
R1242 VDD1.n83 VDD1.n1 0.155672
R1243 VDD1.n76 VDD1.n1 0.155672
R1244 VDD1.n76 VDD1.n75 0.155672
R1245 VDD1.n75 VDD1.n5 0.155672
R1246 VDD1.n68 VDD1.n5 0.155672
R1247 VDD1.n68 VDD1.n67 0.155672
R1248 VDD1.n67 VDD1.n11 0.155672
R1249 VDD1.n60 VDD1.n11 0.155672
R1250 VDD1.n60 VDD1.n59 0.155672
R1251 VDD1.n59 VDD1.n15 0.155672
R1252 VDD1.n52 VDD1.n15 0.155672
R1253 VDD1.n52 VDD1.n51 0.155672
R1254 VDD1.n51 VDD1.n19 0.155672
R1255 VDD1.n44 VDD1.n19 0.155672
R1256 VDD1.n44 VDD1.n43 0.155672
R1257 VDD1.n43 VDD1.n23 0.155672
R1258 VDD1.n36 VDD1.n23 0.155672
R1259 VDD1.n36 VDD1.n35 0.155672
R1260 VDD1.n35 VDD1.n27 0.155672
R1261 VDD1.n118 VDD1.n110 0.155672
R1262 VDD1.n119 VDD1.n118 0.155672
R1263 VDD1.n119 VDD1.n106 0.155672
R1264 VDD1.n126 VDD1.n106 0.155672
R1265 VDD1.n127 VDD1.n126 0.155672
R1266 VDD1.n127 VDD1.n102 0.155672
R1267 VDD1.n134 VDD1.n102 0.155672
R1268 VDD1.n135 VDD1.n134 0.155672
R1269 VDD1.n135 VDD1.n98 0.155672
R1270 VDD1.n142 VDD1.n98 0.155672
R1271 VDD1.n143 VDD1.n142 0.155672
R1272 VDD1.n143 VDD1.n94 0.155672
R1273 VDD1.n150 VDD1.n94 0.155672
R1274 VDD1.n151 VDD1.n150 0.155672
R1275 VDD1.n151 VDD1.n90 0.155672
R1276 VDD1.n160 VDD1.n90 0.155672
R1277 VDD1.n161 VDD1.n160 0.155672
R1278 VDD1.n161 VDD1.n86 0.155672
R1279 VDD1.n168 VDD1.n86 0.155672
R1280 VTAIL.n346 VTAIL.n266 756.745
R1281 VTAIL.n82 VTAIL.n2 756.745
R1282 VTAIL.n260 VTAIL.n180 756.745
R1283 VTAIL.n172 VTAIL.n92 756.745
R1284 VTAIL.n295 VTAIL.n294 585
R1285 VTAIL.n297 VTAIL.n296 585
R1286 VTAIL.n290 VTAIL.n289 585
R1287 VTAIL.n303 VTAIL.n302 585
R1288 VTAIL.n305 VTAIL.n304 585
R1289 VTAIL.n286 VTAIL.n285 585
R1290 VTAIL.n311 VTAIL.n310 585
R1291 VTAIL.n313 VTAIL.n312 585
R1292 VTAIL.n282 VTAIL.n281 585
R1293 VTAIL.n319 VTAIL.n318 585
R1294 VTAIL.n321 VTAIL.n320 585
R1295 VTAIL.n278 VTAIL.n277 585
R1296 VTAIL.n327 VTAIL.n326 585
R1297 VTAIL.n329 VTAIL.n328 585
R1298 VTAIL.n274 VTAIL.n273 585
R1299 VTAIL.n336 VTAIL.n335 585
R1300 VTAIL.n337 VTAIL.n272 585
R1301 VTAIL.n339 VTAIL.n338 585
R1302 VTAIL.n270 VTAIL.n269 585
R1303 VTAIL.n345 VTAIL.n344 585
R1304 VTAIL.n347 VTAIL.n346 585
R1305 VTAIL.n31 VTAIL.n30 585
R1306 VTAIL.n33 VTAIL.n32 585
R1307 VTAIL.n26 VTAIL.n25 585
R1308 VTAIL.n39 VTAIL.n38 585
R1309 VTAIL.n41 VTAIL.n40 585
R1310 VTAIL.n22 VTAIL.n21 585
R1311 VTAIL.n47 VTAIL.n46 585
R1312 VTAIL.n49 VTAIL.n48 585
R1313 VTAIL.n18 VTAIL.n17 585
R1314 VTAIL.n55 VTAIL.n54 585
R1315 VTAIL.n57 VTAIL.n56 585
R1316 VTAIL.n14 VTAIL.n13 585
R1317 VTAIL.n63 VTAIL.n62 585
R1318 VTAIL.n65 VTAIL.n64 585
R1319 VTAIL.n10 VTAIL.n9 585
R1320 VTAIL.n72 VTAIL.n71 585
R1321 VTAIL.n73 VTAIL.n8 585
R1322 VTAIL.n75 VTAIL.n74 585
R1323 VTAIL.n6 VTAIL.n5 585
R1324 VTAIL.n81 VTAIL.n80 585
R1325 VTAIL.n83 VTAIL.n82 585
R1326 VTAIL.n261 VTAIL.n260 585
R1327 VTAIL.n259 VTAIL.n258 585
R1328 VTAIL.n184 VTAIL.n183 585
R1329 VTAIL.n188 VTAIL.n186 585
R1330 VTAIL.n253 VTAIL.n252 585
R1331 VTAIL.n251 VTAIL.n250 585
R1332 VTAIL.n190 VTAIL.n189 585
R1333 VTAIL.n245 VTAIL.n244 585
R1334 VTAIL.n243 VTAIL.n242 585
R1335 VTAIL.n194 VTAIL.n193 585
R1336 VTAIL.n237 VTAIL.n236 585
R1337 VTAIL.n235 VTAIL.n234 585
R1338 VTAIL.n198 VTAIL.n197 585
R1339 VTAIL.n229 VTAIL.n228 585
R1340 VTAIL.n227 VTAIL.n226 585
R1341 VTAIL.n202 VTAIL.n201 585
R1342 VTAIL.n221 VTAIL.n220 585
R1343 VTAIL.n219 VTAIL.n218 585
R1344 VTAIL.n206 VTAIL.n205 585
R1345 VTAIL.n213 VTAIL.n212 585
R1346 VTAIL.n211 VTAIL.n210 585
R1347 VTAIL.n173 VTAIL.n172 585
R1348 VTAIL.n171 VTAIL.n170 585
R1349 VTAIL.n96 VTAIL.n95 585
R1350 VTAIL.n100 VTAIL.n98 585
R1351 VTAIL.n165 VTAIL.n164 585
R1352 VTAIL.n163 VTAIL.n162 585
R1353 VTAIL.n102 VTAIL.n101 585
R1354 VTAIL.n157 VTAIL.n156 585
R1355 VTAIL.n155 VTAIL.n154 585
R1356 VTAIL.n106 VTAIL.n105 585
R1357 VTAIL.n149 VTAIL.n148 585
R1358 VTAIL.n147 VTAIL.n146 585
R1359 VTAIL.n110 VTAIL.n109 585
R1360 VTAIL.n141 VTAIL.n140 585
R1361 VTAIL.n139 VTAIL.n138 585
R1362 VTAIL.n114 VTAIL.n113 585
R1363 VTAIL.n133 VTAIL.n132 585
R1364 VTAIL.n131 VTAIL.n130 585
R1365 VTAIL.n118 VTAIL.n117 585
R1366 VTAIL.n125 VTAIL.n124 585
R1367 VTAIL.n123 VTAIL.n122 585
R1368 VTAIL.n293 VTAIL.t4 327.466
R1369 VTAIL.n29 VTAIL.t8 327.466
R1370 VTAIL.n209 VTAIL.t5 327.466
R1371 VTAIL.n121 VTAIL.t1 327.466
R1372 VTAIL.n296 VTAIL.n295 171.744
R1373 VTAIL.n296 VTAIL.n289 171.744
R1374 VTAIL.n303 VTAIL.n289 171.744
R1375 VTAIL.n304 VTAIL.n303 171.744
R1376 VTAIL.n304 VTAIL.n285 171.744
R1377 VTAIL.n311 VTAIL.n285 171.744
R1378 VTAIL.n312 VTAIL.n311 171.744
R1379 VTAIL.n312 VTAIL.n281 171.744
R1380 VTAIL.n319 VTAIL.n281 171.744
R1381 VTAIL.n320 VTAIL.n319 171.744
R1382 VTAIL.n320 VTAIL.n277 171.744
R1383 VTAIL.n327 VTAIL.n277 171.744
R1384 VTAIL.n328 VTAIL.n327 171.744
R1385 VTAIL.n328 VTAIL.n273 171.744
R1386 VTAIL.n336 VTAIL.n273 171.744
R1387 VTAIL.n337 VTAIL.n336 171.744
R1388 VTAIL.n338 VTAIL.n337 171.744
R1389 VTAIL.n338 VTAIL.n269 171.744
R1390 VTAIL.n345 VTAIL.n269 171.744
R1391 VTAIL.n346 VTAIL.n345 171.744
R1392 VTAIL.n32 VTAIL.n31 171.744
R1393 VTAIL.n32 VTAIL.n25 171.744
R1394 VTAIL.n39 VTAIL.n25 171.744
R1395 VTAIL.n40 VTAIL.n39 171.744
R1396 VTAIL.n40 VTAIL.n21 171.744
R1397 VTAIL.n47 VTAIL.n21 171.744
R1398 VTAIL.n48 VTAIL.n47 171.744
R1399 VTAIL.n48 VTAIL.n17 171.744
R1400 VTAIL.n55 VTAIL.n17 171.744
R1401 VTAIL.n56 VTAIL.n55 171.744
R1402 VTAIL.n56 VTAIL.n13 171.744
R1403 VTAIL.n63 VTAIL.n13 171.744
R1404 VTAIL.n64 VTAIL.n63 171.744
R1405 VTAIL.n64 VTAIL.n9 171.744
R1406 VTAIL.n72 VTAIL.n9 171.744
R1407 VTAIL.n73 VTAIL.n72 171.744
R1408 VTAIL.n74 VTAIL.n73 171.744
R1409 VTAIL.n74 VTAIL.n5 171.744
R1410 VTAIL.n81 VTAIL.n5 171.744
R1411 VTAIL.n82 VTAIL.n81 171.744
R1412 VTAIL.n260 VTAIL.n259 171.744
R1413 VTAIL.n259 VTAIL.n183 171.744
R1414 VTAIL.n188 VTAIL.n183 171.744
R1415 VTAIL.n252 VTAIL.n188 171.744
R1416 VTAIL.n252 VTAIL.n251 171.744
R1417 VTAIL.n251 VTAIL.n189 171.744
R1418 VTAIL.n244 VTAIL.n189 171.744
R1419 VTAIL.n244 VTAIL.n243 171.744
R1420 VTAIL.n243 VTAIL.n193 171.744
R1421 VTAIL.n236 VTAIL.n193 171.744
R1422 VTAIL.n236 VTAIL.n235 171.744
R1423 VTAIL.n235 VTAIL.n197 171.744
R1424 VTAIL.n228 VTAIL.n197 171.744
R1425 VTAIL.n228 VTAIL.n227 171.744
R1426 VTAIL.n227 VTAIL.n201 171.744
R1427 VTAIL.n220 VTAIL.n201 171.744
R1428 VTAIL.n220 VTAIL.n219 171.744
R1429 VTAIL.n219 VTAIL.n205 171.744
R1430 VTAIL.n212 VTAIL.n205 171.744
R1431 VTAIL.n212 VTAIL.n211 171.744
R1432 VTAIL.n172 VTAIL.n171 171.744
R1433 VTAIL.n171 VTAIL.n95 171.744
R1434 VTAIL.n100 VTAIL.n95 171.744
R1435 VTAIL.n164 VTAIL.n100 171.744
R1436 VTAIL.n164 VTAIL.n163 171.744
R1437 VTAIL.n163 VTAIL.n101 171.744
R1438 VTAIL.n156 VTAIL.n101 171.744
R1439 VTAIL.n156 VTAIL.n155 171.744
R1440 VTAIL.n155 VTAIL.n105 171.744
R1441 VTAIL.n148 VTAIL.n105 171.744
R1442 VTAIL.n148 VTAIL.n147 171.744
R1443 VTAIL.n147 VTAIL.n109 171.744
R1444 VTAIL.n140 VTAIL.n109 171.744
R1445 VTAIL.n140 VTAIL.n139 171.744
R1446 VTAIL.n139 VTAIL.n113 171.744
R1447 VTAIL.n132 VTAIL.n113 171.744
R1448 VTAIL.n132 VTAIL.n131 171.744
R1449 VTAIL.n131 VTAIL.n117 171.744
R1450 VTAIL.n124 VTAIL.n117 171.744
R1451 VTAIL.n124 VTAIL.n123 171.744
R1452 VTAIL.n295 VTAIL.t4 85.8723
R1453 VTAIL.n31 VTAIL.t8 85.8723
R1454 VTAIL.n211 VTAIL.t5 85.8723
R1455 VTAIL.n123 VTAIL.t1 85.8723
R1456 VTAIL.n179 VTAIL.n178 57.0703
R1457 VTAIL.n91 VTAIL.n90 57.0703
R1458 VTAIL.n1 VTAIL.n0 57.0701
R1459 VTAIL.n89 VTAIL.n88 57.0701
R1460 VTAIL.n351 VTAIL.n350 35.6763
R1461 VTAIL.n87 VTAIL.n86 35.6763
R1462 VTAIL.n265 VTAIL.n264 35.6763
R1463 VTAIL.n177 VTAIL.n176 35.6763
R1464 VTAIL.n91 VTAIL.n89 27.8324
R1465 VTAIL.n351 VTAIL.n265 26.7979
R1466 VTAIL.n294 VTAIL.n293 16.3895
R1467 VTAIL.n30 VTAIL.n29 16.3895
R1468 VTAIL.n210 VTAIL.n209 16.3895
R1469 VTAIL.n122 VTAIL.n121 16.3895
R1470 VTAIL.n339 VTAIL.n270 13.1884
R1471 VTAIL.n75 VTAIL.n6 13.1884
R1472 VTAIL.n186 VTAIL.n184 13.1884
R1473 VTAIL.n98 VTAIL.n96 13.1884
R1474 VTAIL.n297 VTAIL.n292 12.8005
R1475 VTAIL.n340 VTAIL.n272 12.8005
R1476 VTAIL.n344 VTAIL.n343 12.8005
R1477 VTAIL.n33 VTAIL.n28 12.8005
R1478 VTAIL.n76 VTAIL.n8 12.8005
R1479 VTAIL.n80 VTAIL.n79 12.8005
R1480 VTAIL.n258 VTAIL.n257 12.8005
R1481 VTAIL.n254 VTAIL.n253 12.8005
R1482 VTAIL.n213 VTAIL.n208 12.8005
R1483 VTAIL.n170 VTAIL.n169 12.8005
R1484 VTAIL.n166 VTAIL.n165 12.8005
R1485 VTAIL.n125 VTAIL.n120 12.8005
R1486 VTAIL.n298 VTAIL.n290 12.0247
R1487 VTAIL.n335 VTAIL.n334 12.0247
R1488 VTAIL.n347 VTAIL.n268 12.0247
R1489 VTAIL.n34 VTAIL.n26 12.0247
R1490 VTAIL.n71 VTAIL.n70 12.0247
R1491 VTAIL.n83 VTAIL.n4 12.0247
R1492 VTAIL.n261 VTAIL.n182 12.0247
R1493 VTAIL.n250 VTAIL.n187 12.0247
R1494 VTAIL.n214 VTAIL.n206 12.0247
R1495 VTAIL.n173 VTAIL.n94 12.0247
R1496 VTAIL.n162 VTAIL.n99 12.0247
R1497 VTAIL.n126 VTAIL.n118 12.0247
R1498 VTAIL.n302 VTAIL.n301 11.249
R1499 VTAIL.n333 VTAIL.n274 11.249
R1500 VTAIL.n348 VTAIL.n266 11.249
R1501 VTAIL.n38 VTAIL.n37 11.249
R1502 VTAIL.n69 VTAIL.n10 11.249
R1503 VTAIL.n84 VTAIL.n2 11.249
R1504 VTAIL.n262 VTAIL.n180 11.249
R1505 VTAIL.n249 VTAIL.n190 11.249
R1506 VTAIL.n218 VTAIL.n217 11.249
R1507 VTAIL.n174 VTAIL.n92 11.249
R1508 VTAIL.n161 VTAIL.n102 11.249
R1509 VTAIL.n130 VTAIL.n129 11.249
R1510 VTAIL.n305 VTAIL.n288 10.4732
R1511 VTAIL.n330 VTAIL.n329 10.4732
R1512 VTAIL.n41 VTAIL.n24 10.4732
R1513 VTAIL.n66 VTAIL.n65 10.4732
R1514 VTAIL.n246 VTAIL.n245 10.4732
R1515 VTAIL.n221 VTAIL.n204 10.4732
R1516 VTAIL.n158 VTAIL.n157 10.4732
R1517 VTAIL.n133 VTAIL.n116 10.4732
R1518 VTAIL.n306 VTAIL.n286 9.69747
R1519 VTAIL.n326 VTAIL.n276 9.69747
R1520 VTAIL.n42 VTAIL.n22 9.69747
R1521 VTAIL.n62 VTAIL.n12 9.69747
R1522 VTAIL.n242 VTAIL.n192 9.69747
R1523 VTAIL.n222 VTAIL.n202 9.69747
R1524 VTAIL.n154 VTAIL.n104 9.69747
R1525 VTAIL.n134 VTAIL.n114 9.69747
R1526 VTAIL.n350 VTAIL.n349 9.45567
R1527 VTAIL.n86 VTAIL.n85 9.45567
R1528 VTAIL.n264 VTAIL.n263 9.45567
R1529 VTAIL.n176 VTAIL.n175 9.45567
R1530 VTAIL.n349 VTAIL.n348 9.3005
R1531 VTAIL.n268 VTAIL.n267 9.3005
R1532 VTAIL.n343 VTAIL.n342 9.3005
R1533 VTAIL.n315 VTAIL.n314 9.3005
R1534 VTAIL.n284 VTAIL.n283 9.3005
R1535 VTAIL.n309 VTAIL.n308 9.3005
R1536 VTAIL.n307 VTAIL.n306 9.3005
R1537 VTAIL.n288 VTAIL.n287 9.3005
R1538 VTAIL.n301 VTAIL.n300 9.3005
R1539 VTAIL.n299 VTAIL.n298 9.3005
R1540 VTAIL.n292 VTAIL.n291 9.3005
R1541 VTAIL.n317 VTAIL.n316 9.3005
R1542 VTAIL.n280 VTAIL.n279 9.3005
R1543 VTAIL.n323 VTAIL.n322 9.3005
R1544 VTAIL.n325 VTAIL.n324 9.3005
R1545 VTAIL.n276 VTAIL.n275 9.3005
R1546 VTAIL.n331 VTAIL.n330 9.3005
R1547 VTAIL.n333 VTAIL.n332 9.3005
R1548 VTAIL.n334 VTAIL.n271 9.3005
R1549 VTAIL.n341 VTAIL.n340 9.3005
R1550 VTAIL.n85 VTAIL.n84 9.3005
R1551 VTAIL.n4 VTAIL.n3 9.3005
R1552 VTAIL.n79 VTAIL.n78 9.3005
R1553 VTAIL.n51 VTAIL.n50 9.3005
R1554 VTAIL.n20 VTAIL.n19 9.3005
R1555 VTAIL.n45 VTAIL.n44 9.3005
R1556 VTAIL.n43 VTAIL.n42 9.3005
R1557 VTAIL.n24 VTAIL.n23 9.3005
R1558 VTAIL.n37 VTAIL.n36 9.3005
R1559 VTAIL.n35 VTAIL.n34 9.3005
R1560 VTAIL.n28 VTAIL.n27 9.3005
R1561 VTAIL.n53 VTAIL.n52 9.3005
R1562 VTAIL.n16 VTAIL.n15 9.3005
R1563 VTAIL.n59 VTAIL.n58 9.3005
R1564 VTAIL.n61 VTAIL.n60 9.3005
R1565 VTAIL.n12 VTAIL.n11 9.3005
R1566 VTAIL.n67 VTAIL.n66 9.3005
R1567 VTAIL.n69 VTAIL.n68 9.3005
R1568 VTAIL.n70 VTAIL.n7 9.3005
R1569 VTAIL.n77 VTAIL.n76 9.3005
R1570 VTAIL.n196 VTAIL.n195 9.3005
R1571 VTAIL.n239 VTAIL.n238 9.3005
R1572 VTAIL.n241 VTAIL.n240 9.3005
R1573 VTAIL.n192 VTAIL.n191 9.3005
R1574 VTAIL.n247 VTAIL.n246 9.3005
R1575 VTAIL.n249 VTAIL.n248 9.3005
R1576 VTAIL.n187 VTAIL.n185 9.3005
R1577 VTAIL.n255 VTAIL.n254 9.3005
R1578 VTAIL.n263 VTAIL.n262 9.3005
R1579 VTAIL.n182 VTAIL.n181 9.3005
R1580 VTAIL.n257 VTAIL.n256 9.3005
R1581 VTAIL.n233 VTAIL.n232 9.3005
R1582 VTAIL.n231 VTAIL.n230 9.3005
R1583 VTAIL.n200 VTAIL.n199 9.3005
R1584 VTAIL.n225 VTAIL.n224 9.3005
R1585 VTAIL.n223 VTAIL.n222 9.3005
R1586 VTAIL.n204 VTAIL.n203 9.3005
R1587 VTAIL.n217 VTAIL.n216 9.3005
R1588 VTAIL.n215 VTAIL.n214 9.3005
R1589 VTAIL.n208 VTAIL.n207 9.3005
R1590 VTAIL.n108 VTAIL.n107 9.3005
R1591 VTAIL.n151 VTAIL.n150 9.3005
R1592 VTAIL.n153 VTAIL.n152 9.3005
R1593 VTAIL.n104 VTAIL.n103 9.3005
R1594 VTAIL.n159 VTAIL.n158 9.3005
R1595 VTAIL.n161 VTAIL.n160 9.3005
R1596 VTAIL.n99 VTAIL.n97 9.3005
R1597 VTAIL.n167 VTAIL.n166 9.3005
R1598 VTAIL.n175 VTAIL.n174 9.3005
R1599 VTAIL.n94 VTAIL.n93 9.3005
R1600 VTAIL.n169 VTAIL.n168 9.3005
R1601 VTAIL.n145 VTAIL.n144 9.3005
R1602 VTAIL.n143 VTAIL.n142 9.3005
R1603 VTAIL.n112 VTAIL.n111 9.3005
R1604 VTAIL.n137 VTAIL.n136 9.3005
R1605 VTAIL.n135 VTAIL.n134 9.3005
R1606 VTAIL.n116 VTAIL.n115 9.3005
R1607 VTAIL.n129 VTAIL.n128 9.3005
R1608 VTAIL.n127 VTAIL.n126 9.3005
R1609 VTAIL.n120 VTAIL.n119 9.3005
R1610 VTAIL.n310 VTAIL.n309 8.92171
R1611 VTAIL.n325 VTAIL.n278 8.92171
R1612 VTAIL.n46 VTAIL.n45 8.92171
R1613 VTAIL.n61 VTAIL.n14 8.92171
R1614 VTAIL.n241 VTAIL.n194 8.92171
R1615 VTAIL.n226 VTAIL.n225 8.92171
R1616 VTAIL.n153 VTAIL.n106 8.92171
R1617 VTAIL.n138 VTAIL.n137 8.92171
R1618 VTAIL.n313 VTAIL.n284 8.14595
R1619 VTAIL.n322 VTAIL.n321 8.14595
R1620 VTAIL.n49 VTAIL.n20 8.14595
R1621 VTAIL.n58 VTAIL.n57 8.14595
R1622 VTAIL.n238 VTAIL.n237 8.14595
R1623 VTAIL.n229 VTAIL.n200 8.14595
R1624 VTAIL.n150 VTAIL.n149 8.14595
R1625 VTAIL.n141 VTAIL.n112 8.14595
R1626 VTAIL.n314 VTAIL.n282 7.3702
R1627 VTAIL.n318 VTAIL.n280 7.3702
R1628 VTAIL.n50 VTAIL.n18 7.3702
R1629 VTAIL.n54 VTAIL.n16 7.3702
R1630 VTAIL.n234 VTAIL.n196 7.3702
R1631 VTAIL.n230 VTAIL.n198 7.3702
R1632 VTAIL.n146 VTAIL.n108 7.3702
R1633 VTAIL.n142 VTAIL.n110 7.3702
R1634 VTAIL.n317 VTAIL.n282 6.59444
R1635 VTAIL.n318 VTAIL.n317 6.59444
R1636 VTAIL.n53 VTAIL.n18 6.59444
R1637 VTAIL.n54 VTAIL.n53 6.59444
R1638 VTAIL.n234 VTAIL.n233 6.59444
R1639 VTAIL.n233 VTAIL.n198 6.59444
R1640 VTAIL.n146 VTAIL.n145 6.59444
R1641 VTAIL.n145 VTAIL.n110 6.59444
R1642 VTAIL.n314 VTAIL.n313 5.81868
R1643 VTAIL.n321 VTAIL.n280 5.81868
R1644 VTAIL.n50 VTAIL.n49 5.81868
R1645 VTAIL.n57 VTAIL.n16 5.81868
R1646 VTAIL.n237 VTAIL.n196 5.81868
R1647 VTAIL.n230 VTAIL.n229 5.81868
R1648 VTAIL.n149 VTAIL.n108 5.81868
R1649 VTAIL.n142 VTAIL.n141 5.81868
R1650 VTAIL.n310 VTAIL.n284 5.04292
R1651 VTAIL.n322 VTAIL.n278 5.04292
R1652 VTAIL.n46 VTAIL.n20 5.04292
R1653 VTAIL.n58 VTAIL.n14 5.04292
R1654 VTAIL.n238 VTAIL.n194 5.04292
R1655 VTAIL.n226 VTAIL.n200 5.04292
R1656 VTAIL.n150 VTAIL.n106 5.04292
R1657 VTAIL.n138 VTAIL.n112 5.04292
R1658 VTAIL.n309 VTAIL.n286 4.26717
R1659 VTAIL.n326 VTAIL.n325 4.26717
R1660 VTAIL.n45 VTAIL.n22 4.26717
R1661 VTAIL.n62 VTAIL.n61 4.26717
R1662 VTAIL.n242 VTAIL.n241 4.26717
R1663 VTAIL.n225 VTAIL.n202 4.26717
R1664 VTAIL.n154 VTAIL.n153 4.26717
R1665 VTAIL.n137 VTAIL.n114 4.26717
R1666 VTAIL.n293 VTAIL.n291 3.70982
R1667 VTAIL.n29 VTAIL.n27 3.70982
R1668 VTAIL.n209 VTAIL.n207 3.70982
R1669 VTAIL.n121 VTAIL.n119 3.70982
R1670 VTAIL.n306 VTAIL.n305 3.49141
R1671 VTAIL.n329 VTAIL.n276 3.49141
R1672 VTAIL.n42 VTAIL.n41 3.49141
R1673 VTAIL.n65 VTAIL.n12 3.49141
R1674 VTAIL.n245 VTAIL.n192 3.49141
R1675 VTAIL.n222 VTAIL.n221 3.49141
R1676 VTAIL.n157 VTAIL.n104 3.49141
R1677 VTAIL.n134 VTAIL.n133 3.49141
R1678 VTAIL.n302 VTAIL.n288 2.71565
R1679 VTAIL.n330 VTAIL.n274 2.71565
R1680 VTAIL.n350 VTAIL.n266 2.71565
R1681 VTAIL.n38 VTAIL.n24 2.71565
R1682 VTAIL.n66 VTAIL.n10 2.71565
R1683 VTAIL.n86 VTAIL.n2 2.71565
R1684 VTAIL.n264 VTAIL.n180 2.71565
R1685 VTAIL.n246 VTAIL.n190 2.71565
R1686 VTAIL.n218 VTAIL.n204 2.71565
R1687 VTAIL.n176 VTAIL.n92 2.71565
R1688 VTAIL.n158 VTAIL.n102 2.71565
R1689 VTAIL.n130 VTAIL.n116 2.71565
R1690 VTAIL.n0 VTAIL.t11 2.0922
R1691 VTAIL.n0 VTAIL.t3 2.0922
R1692 VTAIL.n88 VTAIL.t7 2.0922
R1693 VTAIL.n88 VTAIL.t10 2.0922
R1694 VTAIL.n178 VTAIL.t9 2.0922
R1695 VTAIL.n178 VTAIL.t6 2.0922
R1696 VTAIL.n90 VTAIL.t0 2.0922
R1697 VTAIL.n90 VTAIL.t2 2.0922
R1698 VTAIL.n301 VTAIL.n290 1.93989
R1699 VTAIL.n335 VTAIL.n333 1.93989
R1700 VTAIL.n348 VTAIL.n347 1.93989
R1701 VTAIL.n37 VTAIL.n26 1.93989
R1702 VTAIL.n71 VTAIL.n69 1.93989
R1703 VTAIL.n84 VTAIL.n83 1.93989
R1704 VTAIL.n262 VTAIL.n261 1.93989
R1705 VTAIL.n250 VTAIL.n249 1.93989
R1706 VTAIL.n217 VTAIL.n206 1.93989
R1707 VTAIL.n174 VTAIL.n173 1.93989
R1708 VTAIL.n162 VTAIL.n161 1.93989
R1709 VTAIL.n129 VTAIL.n118 1.93989
R1710 VTAIL.n298 VTAIL.n297 1.16414
R1711 VTAIL.n334 VTAIL.n272 1.16414
R1712 VTAIL.n344 VTAIL.n268 1.16414
R1713 VTAIL.n34 VTAIL.n33 1.16414
R1714 VTAIL.n70 VTAIL.n8 1.16414
R1715 VTAIL.n80 VTAIL.n4 1.16414
R1716 VTAIL.n258 VTAIL.n182 1.16414
R1717 VTAIL.n253 VTAIL.n187 1.16414
R1718 VTAIL.n214 VTAIL.n213 1.16414
R1719 VTAIL.n170 VTAIL.n94 1.16414
R1720 VTAIL.n165 VTAIL.n99 1.16414
R1721 VTAIL.n126 VTAIL.n125 1.16414
R1722 VTAIL.n177 VTAIL.n91 1.03498
R1723 VTAIL.n265 VTAIL.n179 1.03498
R1724 VTAIL.n89 VTAIL.n87 1.03498
R1725 VTAIL.n179 VTAIL.n177 0.987569
R1726 VTAIL.n87 VTAIL.n1 0.987569
R1727 VTAIL VTAIL.n351 0.718172
R1728 VTAIL.n294 VTAIL.n292 0.388379
R1729 VTAIL.n340 VTAIL.n339 0.388379
R1730 VTAIL.n343 VTAIL.n270 0.388379
R1731 VTAIL.n30 VTAIL.n28 0.388379
R1732 VTAIL.n76 VTAIL.n75 0.388379
R1733 VTAIL.n79 VTAIL.n6 0.388379
R1734 VTAIL.n257 VTAIL.n184 0.388379
R1735 VTAIL.n254 VTAIL.n186 0.388379
R1736 VTAIL.n210 VTAIL.n208 0.388379
R1737 VTAIL.n169 VTAIL.n96 0.388379
R1738 VTAIL.n166 VTAIL.n98 0.388379
R1739 VTAIL.n122 VTAIL.n120 0.388379
R1740 VTAIL VTAIL.n1 0.31731
R1741 VTAIL.n299 VTAIL.n291 0.155672
R1742 VTAIL.n300 VTAIL.n299 0.155672
R1743 VTAIL.n300 VTAIL.n287 0.155672
R1744 VTAIL.n307 VTAIL.n287 0.155672
R1745 VTAIL.n308 VTAIL.n307 0.155672
R1746 VTAIL.n308 VTAIL.n283 0.155672
R1747 VTAIL.n315 VTAIL.n283 0.155672
R1748 VTAIL.n316 VTAIL.n315 0.155672
R1749 VTAIL.n316 VTAIL.n279 0.155672
R1750 VTAIL.n323 VTAIL.n279 0.155672
R1751 VTAIL.n324 VTAIL.n323 0.155672
R1752 VTAIL.n324 VTAIL.n275 0.155672
R1753 VTAIL.n331 VTAIL.n275 0.155672
R1754 VTAIL.n332 VTAIL.n331 0.155672
R1755 VTAIL.n332 VTAIL.n271 0.155672
R1756 VTAIL.n341 VTAIL.n271 0.155672
R1757 VTAIL.n342 VTAIL.n341 0.155672
R1758 VTAIL.n342 VTAIL.n267 0.155672
R1759 VTAIL.n349 VTAIL.n267 0.155672
R1760 VTAIL.n35 VTAIL.n27 0.155672
R1761 VTAIL.n36 VTAIL.n35 0.155672
R1762 VTAIL.n36 VTAIL.n23 0.155672
R1763 VTAIL.n43 VTAIL.n23 0.155672
R1764 VTAIL.n44 VTAIL.n43 0.155672
R1765 VTAIL.n44 VTAIL.n19 0.155672
R1766 VTAIL.n51 VTAIL.n19 0.155672
R1767 VTAIL.n52 VTAIL.n51 0.155672
R1768 VTAIL.n52 VTAIL.n15 0.155672
R1769 VTAIL.n59 VTAIL.n15 0.155672
R1770 VTAIL.n60 VTAIL.n59 0.155672
R1771 VTAIL.n60 VTAIL.n11 0.155672
R1772 VTAIL.n67 VTAIL.n11 0.155672
R1773 VTAIL.n68 VTAIL.n67 0.155672
R1774 VTAIL.n68 VTAIL.n7 0.155672
R1775 VTAIL.n77 VTAIL.n7 0.155672
R1776 VTAIL.n78 VTAIL.n77 0.155672
R1777 VTAIL.n78 VTAIL.n3 0.155672
R1778 VTAIL.n85 VTAIL.n3 0.155672
R1779 VTAIL.n263 VTAIL.n181 0.155672
R1780 VTAIL.n256 VTAIL.n181 0.155672
R1781 VTAIL.n256 VTAIL.n255 0.155672
R1782 VTAIL.n255 VTAIL.n185 0.155672
R1783 VTAIL.n248 VTAIL.n185 0.155672
R1784 VTAIL.n248 VTAIL.n247 0.155672
R1785 VTAIL.n247 VTAIL.n191 0.155672
R1786 VTAIL.n240 VTAIL.n191 0.155672
R1787 VTAIL.n240 VTAIL.n239 0.155672
R1788 VTAIL.n239 VTAIL.n195 0.155672
R1789 VTAIL.n232 VTAIL.n195 0.155672
R1790 VTAIL.n232 VTAIL.n231 0.155672
R1791 VTAIL.n231 VTAIL.n199 0.155672
R1792 VTAIL.n224 VTAIL.n199 0.155672
R1793 VTAIL.n224 VTAIL.n223 0.155672
R1794 VTAIL.n223 VTAIL.n203 0.155672
R1795 VTAIL.n216 VTAIL.n203 0.155672
R1796 VTAIL.n216 VTAIL.n215 0.155672
R1797 VTAIL.n215 VTAIL.n207 0.155672
R1798 VTAIL.n175 VTAIL.n93 0.155672
R1799 VTAIL.n168 VTAIL.n93 0.155672
R1800 VTAIL.n168 VTAIL.n167 0.155672
R1801 VTAIL.n167 VTAIL.n97 0.155672
R1802 VTAIL.n160 VTAIL.n97 0.155672
R1803 VTAIL.n160 VTAIL.n159 0.155672
R1804 VTAIL.n159 VTAIL.n103 0.155672
R1805 VTAIL.n152 VTAIL.n103 0.155672
R1806 VTAIL.n152 VTAIL.n151 0.155672
R1807 VTAIL.n151 VTAIL.n107 0.155672
R1808 VTAIL.n144 VTAIL.n107 0.155672
R1809 VTAIL.n144 VTAIL.n143 0.155672
R1810 VTAIL.n143 VTAIL.n111 0.155672
R1811 VTAIL.n136 VTAIL.n111 0.155672
R1812 VTAIL.n136 VTAIL.n135 0.155672
R1813 VTAIL.n135 VTAIL.n115 0.155672
R1814 VTAIL.n128 VTAIL.n115 0.155672
R1815 VTAIL.n128 VTAIL.n127 0.155672
R1816 VTAIL.n127 VTAIL.n119 0.155672
R1817 VN.n2 VN.t5 491.878
R1818 VN.n10 VN.t0 491.878
R1819 VN.n6 VN.t2 475.63
R1820 VN.n14 VN.t1 475.63
R1821 VN.n1 VN.t4 430.476
R1822 VN.n9 VN.t3 430.476
R1823 VN.n7 VN.n6 161.3
R1824 VN.n15 VN.n14 161.3
R1825 VN.n13 VN.n8 161.3
R1826 VN.n12 VN.n11 161.3
R1827 VN.n5 VN.n0 161.3
R1828 VN.n4 VN.n3 161.3
R1829 VN.n5 VN.n4 55.1086
R1830 VN.n13 VN.n12 55.1086
R1831 VN VN.n15 44.9115
R1832 VN.n11 VN.n10 43.7016
R1833 VN.n3 VN.n2 43.7016
R1834 VN.n2 VN.n1 42.7308
R1835 VN.n10 VN.n9 42.7308
R1836 VN.n4 VN.n1 12.2964
R1837 VN.n12 VN.n9 12.2964
R1838 VN.n6 VN.n5 2.19141
R1839 VN.n14 VN.n13 2.19141
R1840 VN.n15 VN.n8 0.189894
R1841 VN.n11 VN.n8 0.189894
R1842 VN.n3 VN.n0 0.189894
R1843 VN.n7 VN.n0 0.189894
R1844 VN VN.n7 0.0516364
R1845 VDD2.n167 VDD2.n87 756.745
R1846 VDD2.n80 VDD2.n0 756.745
R1847 VDD2.n168 VDD2.n167 585
R1848 VDD2.n166 VDD2.n165 585
R1849 VDD2.n91 VDD2.n90 585
R1850 VDD2.n95 VDD2.n93 585
R1851 VDD2.n160 VDD2.n159 585
R1852 VDD2.n158 VDD2.n157 585
R1853 VDD2.n97 VDD2.n96 585
R1854 VDD2.n152 VDD2.n151 585
R1855 VDD2.n150 VDD2.n149 585
R1856 VDD2.n101 VDD2.n100 585
R1857 VDD2.n144 VDD2.n143 585
R1858 VDD2.n142 VDD2.n141 585
R1859 VDD2.n105 VDD2.n104 585
R1860 VDD2.n136 VDD2.n135 585
R1861 VDD2.n134 VDD2.n133 585
R1862 VDD2.n109 VDD2.n108 585
R1863 VDD2.n128 VDD2.n127 585
R1864 VDD2.n126 VDD2.n125 585
R1865 VDD2.n113 VDD2.n112 585
R1866 VDD2.n120 VDD2.n119 585
R1867 VDD2.n118 VDD2.n117 585
R1868 VDD2.n29 VDD2.n28 585
R1869 VDD2.n31 VDD2.n30 585
R1870 VDD2.n24 VDD2.n23 585
R1871 VDD2.n37 VDD2.n36 585
R1872 VDD2.n39 VDD2.n38 585
R1873 VDD2.n20 VDD2.n19 585
R1874 VDD2.n45 VDD2.n44 585
R1875 VDD2.n47 VDD2.n46 585
R1876 VDD2.n16 VDD2.n15 585
R1877 VDD2.n53 VDD2.n52 585
R1878 VDD2.n55 VDD2.n54 585
R1879 VDD2.n12 VDD2.n11 585
R1880 VDD2.n61 VDD2.n60 585
R1881 VDD2.n63 VDD2.n62 585
R1882 VDD2.n8 VDD2.n7 585
R1883 VDD2.n70 VDD2.n69 585
R1884 VDD2.n71 VDD2.n6 585
R1885 VDD2.n73 VDD2.n72 585
R1886 VDD2.n4 VDD2.n3 585
R1887 VDD2.n79 VDD2.n78 585
R1888 VDD2.n81 VDD2.n80 585
R1889 VDD2.n116 VDD2.t4 327.466
R1890 VDD2.n27 VDD2.t0 327.466
R1891 VDD2.n167 VDD2.n166 171.744
R1892 VDD2.n166 VDD2.n90 171.744
R1893 VDD2.n95 VDD2.n90 171.744
R1894 VDD2.n159 VDD2.n95 171.744
R1895 VDD2.n159 VDD2.n158 171.744
R1896 VDD2.n158 VDD2.n96 171.744
R1897 VDD2.n151 VDD2.n96 171.744
R1898 VDD2.n151 VDD2.n150 171.744
R1899 VDD2.n150 VDD2.n100 171.744
R1900 VDD2.n143 VDD2.n100 171.744
R1901 VDD2.n143 VDD2.n142 171.744
R1902 VDD2.n142 VDD2.n104 171.744
R1903 VDD2.n135 VDD2.n104 171.744
R1904 VDD2.n135 VDD2.n134 171.744
R1905 VDD2.n134 VDD2.n108 171.744
R1906 VDD2.n127 VDD2.n108 171.744
R1907 VDD2.n127 VDD2.n126 171.744
R1908 VDD2.n126 VDD2.n112 171.744
R1909 VDD2.n119 VDD2.n112 171.744
R1910 VDD2.n119 VDD2.n118 171.744
R1911 VDD2.n30 VDD2.n29 171.744
R1912 VDD2.n30 VDD2.n23 171.744
R1913 VDD2.n37 VDD2.n23 171.744
R1914 VDD2.n38 VDD2.n37 171.744
R1915 VDD2.n38 VDD2.n19 171.744
R1916 VDD2.n45 VDD2.n19 171.744
R1917 VDD2.n46 VDD2.n45 171.744
R1918 VDD2.n46 VDD2.n15 171.744
R1919 VDD2.n53 VDD2.n15 171.744
R1920 VDD2.n54 VDD2.n53 171.744
R1921 VDD2.n54 VDD2.n11 171.744
R1922 VDD2.n61 VDD2.n11 171.744
R1923 VDD2.n62 VDD2.n61 171.744
R1924 VDD2.n62 VDD2.n7 171.744
R1925 VDD2.n70 VDD2.n7 171.744
R1926 VDD2.n71 VDD2.n70 171.744
R1927 VDD2.n72 VDD2.n71 171.744
R1928 VDD2.n72 VDD2.n3 171.744
R1929 VDD2.n79 VDD2.n3 171.744
R1930 VDD2.n80 VDD2.n79 171.744
R1931 VDD2.n118 VDD2.t4 85.8723
R1932 VDD2.n29 VDD2.t0 85.8723
R1933 VDD2.n86 VDD2.n85 73.9521
R1934 VDD2 VDD2.n173 73.9493
R1935 VDD2.n86 VDD2.n84 53.0756
R1936 VDD2.n172 VDD2.n171 52.355
R1937 VDD2.n172 VDD2.n86 40.4739
R1938 VDD2.n117 VDD2.n116 16.3895
R1939 VDD2.n28 VDD2.n27 16.3895
R1940 VDD2.n93 VDD2.n91 13.1884
R1941 VDD2.n73 VDD2.n4 13.1884
R1942 VDD2.n165 VDD2.n164 12.8005
R1943 VDD2.n161 VDD2.n160 12.8005
R1944 VDD2.n120 VDD2.n115 12.8005
R1945 VDD2.n31 VDD2.n26 12.8005
R1946 VDD2.n74 VDD2.n6 12.8005
R1947 VDD2.n78 VDD2.n77 12.8005
R1948 VDD2.n168 VDD2.n89 12.0247
R1949 VDD2.n157 VDD2.n94 12.0247
R1950 VDD2.n121 VDD2.n113 12.0247
R1951 VDD2.n32 VDD2.n24 12.0247
R1952 VDD2.n69 VDD2.n68 12.0247
R1953 VDD2.n81 VDD2.n2 12.0247
R1954 VDD2.n169 VDD2.n87 11.249
R1955 VDD2.n156 VDD2.n97 11.249
R1956 VDD2.n125 VDD2.n124 11.249
R1957 VDD2.n36 VDD2.n35 11.249
R1958 VDD2.n67 VDD2.n8 11.249
R1959 VDD2.n82 VDD2.n0 11.249
R1960 VDD2.n153 VDD2.n152 10.4732
R1961 VDD2.n128 VDD2.n111 10.4732
R1962 VDD2.n39 VDD2.n22 10.4732
R1963 VDD2.n64 VDD2.n63 10.4732
R1964 VDD2.n149 VDD2.n99 9.69747
R1965 VDD2.n129 VDD2.n109 9.69747
R1966 VDD2.n40 VDD2.n20 9.69747
R1967 VDD2.n60 VDD2.n10 9.69747
R1968 VDD2.n171 VDD2.n170 9.45567
R1969 VDD2.n84 VDD2.n83 9.45567
R1970 VDD2.n103 VDD2.n102 9.3005
R1971 VDD2.n146 VDD2.n145 9.3005
R1972 VDD2.n148 VDD2.n147 9.3005
R1973 VDD2.n99 VDD2.n98 9.3005
R1974 VDD2.n154 VDD2.n153 9.3005
R1975 VDD2.n156 VDD2.n155 9.3005
R1976 VDD2.n94 VDD2.n92 9.3005
R1977 VDD2.n162 VDD2.n161 9.3005
R1978 VDD2.n170 VDD2.n169 9.3005
R1979 VDD2.n89 VDD2.n88 9.3005
R1980 VDD2.n164 VDD2.n163 9.3005
R1981 VDD2.n140 VDD2.n139 9.3005
R1982 VDD2.n138 VDD2.n137 9.3005
R1983 VDD2.n107 VDD2.n106 9.3005
R1984 VDD2.n132 VDD2.n131 9.3005
R1985 VDD2.n130 VDD2.n129 9.3005
R1986 VDD2.n111 VDD2.n110 9.3005
R1987 VDD2.n124 VDD2.n123 9.3005
R1988 VDD2.n122 VDD2.n121 9.3005
R1989 VDD2.n115 VDD2.n114 9.3005
R1990 VDD2.n83 VDD2.n82 9.3005
R1991 VDD2.n2 VDD2.n1 9.3005
R1992 VDD2.n77 VDD2.n76 9.3005
R1993 VDD2.n49 VDD2.n48 9.3005
R1994 VDD2.n18 VDD2.n17 9.3005
R1995 VDD2.n43 VDD2.n42 9.3005
R1996 VDD2.n41 VDD2.n40 9.3005
R1997 VDD2.n22 VDD2.n21 9.3005
R1998 VDD2.n35 VDD2.n34 9.3005
R1999 VDD2.n33 VDD2.n32 9.3005
R2000 VDD2.n26 VDD2.n25 9.3005
R2001 VDD2.n51 VDD2.n50 9.3005
R2002 VDD2.n14 VDD2.n13 9.3005
R2003 VDD2.n57 VDD2.n56 9.3005
R2004 VDD2.n59 VDD2.n58 9.3005
R2005 VDD2.n10 VDD2.n9 9.3005
R2006 VDD2.n65 VDD2.n64 9.3005
R2007 VDD2.n67 VDD2.n66 9.3005
R2008 VDD2.n68 VDD2.n5 9.3005
R2009 VDD2.n75 VDD2.n74 9.3005
R2010 VDD2.n148 VDD2.n101 8.92171
R2011 VDD2.n133 VDD2.n132 8.92171
R2012 VDD2.n44 VDD2.n43 8.92171
R2013 VDD2.n59 VDD2.n12 8.92171
R2014 VDD2.n145 VDD2.n144 8.14595
R2015 VDD2.n136 VDD2.n107 8.14595
R2016 VDD2.n47 VDD2.n18 8.14595
R2017 VDD2.n56 VDD2.n55 8.14595
R2018 VDD2.n141 VDD2.n103 7.3702
R2019 VDD2.n137 VDD2.n105 7.3702
R2020 VDD2.n48 VDD2.n16 7.3702
R2021 VDD2.n52 VDD2.n14 7.3702
R2022 VDD2.n141 VDD2.n140 6.59444
R2023 VDD2.n140 VDD2.n105 6.59444
R2024 VDD2.n51 VDD2.n16 6.59444
R2025 VDD2.n52 VDD2.n51 6.59444
R2026 VDD2.n144 VDD2.n103 5.81868
R2027 VDD2.n137 VDD2.n136 5.81868
R2028 VDD2.n48 VDD2.n47 5.81868
R2029 VDD2.n55 VDD2.n14 5.81868
R2030 VDD2.n145 VDD2.n101 5.04292
R2031 VDD2.n133 VDD2.n107 5.04292
R2032 VDD2.n44 VDD2.n18 5.04292
R2033 VDD2.n56 VDD2.n12 5.04292
R2034 VDD2.n149 VDD2.n148 4.26717
R2035 VDD2.n132 VDD2.n109 4.26717
R2036 VDD2.n43 VDD2.n20 4.26717
R2037 VDD2.n60 VDD2.n59 4.26717
R2038 VDD2.n116 VDD2.n114 3.70982
R2039 VDD2.n27 VDD2.n25 3.70982
R2040 VDD2.n152 VDD2.n99 3.49141
R2041 VDD2.n129 VDD2.n128 3.49141
R2042 VDD2.n40 VDD2.n39 3.49141
R2043 VDD2.n63 VDD2.n10 3.49141
R2044 VDD2.n171 VDD2.n87 2.71565
R2045 VDD2.n153 VDD2.n97 2.71565
R2046 VDD2.n125 VDD2.n111 2.71565
R2047 VDD2.n36 VDD2.n22 2.71565
R2048 VDD2.n64 VDD2.n8 2.71565
R2049 VDD2.n84 VDD2.n0 2.71565
R2050 VDD2.n173 VDD2.t2 2.0922
R2051 VDD2.n173 VDD2.t5 2.0922
R2052 VDD2.n85 VDD2.t1 2.0922
R2053 VDD2.n85 VDD2.t3 2.0922
R2054 VDD2.n169 VDD2.n168 1.93989
R2055 VDD2.n157 VDD2.n156 1.93989
R2056 VDD2.n124 VDD2.n113 1.93989
R2057 VDD2.n35 VDD2.n24 1.93989
R2058 VDD2.n69 VDD2.n67 1.93989
R2059 VDD2.n82 VDD2.n81 1.93989
R2060 VDD2.n165 VDD2.n89 1.16414
R2061 VDD2.n160 VDD2.n94 1.16414
R2062 VDD2.n121 VDD2.n120 1.16414
R2063 VDD2.n32 VDD2.n31 1.16414
R2064 VDD2.n68 VDD2.n6 1.16414
R2065 VDD2.n78 VDD2.n2 1.16414
R2066 VDD2 VDD2.n172 0.834552
R2067 VDD2.n164 VDD2.n91 0.388379
R2068 VDD2.n161 VDD2.n93 0.388379
R2069 VDD2.n117 VDD2.n115 0.388379
R2070 VDD2.n28 VDD2.n26 0.388379
R2071 VDD2.n74 VDD2.n73 0.388379
R2072 VDD2.n77 VDD2.n4 0.388379
R2073 VDD2.n170 VDD2.n88 0.155672
R2074 VDD2.n163 VDD2.n88 0.155672
R2075 VDD2.n163 VDD2.n162 0.155672
R2076 VDD2.n162 VDD2.n92 0.155672
R2077 VDD2.n155 VDD2.n92 0.155672
R2078 VDD2.n155 VDD2.n154 0.155672
R2079 VDD2.n154 VDD2.n98 0.155672
R2080 VDD2.n147 VDD2.n98 0.155672
R2081 VDD2.n147 VDD2.n146 0.155672
R2082 VDD2.n146 VDD2.n102 0.155672
R2083 VDD2.n139 VDD2.n102 0.155672
R2084 VDD2.n139 VDD2.n138 0.155672
R2085 VDD2.n138 VDD2.n106 0.155672
R2086 VDD2.n131 VDD2.n106 0.155672
R2087 VDD2.n131 VDD2.n130 0.155672
R2088 VDD2.n130 VDD2.n110 0.155672
R2089 VDD2.n123 VDD2.n110 0.155672
R2090 VDD2.n123 VDD2.n122 0.155672
R2091 VDD2.n122 VDD2.n114 0.155672
R2092 VDD2.n33 VDD2.n25 0.155672
R2093 VDD2.n34 VDD2.n33 0.155672
R2094 VDD2.n34 VDD2.n21 0.155672
R2095 VDD2.n41 VDD2.n21 0.155672
R2096 VDD2.n42 VDD2.n41 0.155672
R2097 VDD2.n42 VDD2.n17 0.155672
R2098 VDD2.n49 VDD2.n17 0.155672
R2099 VDD2.n50 VDD2.n49 0.155672
R2100 VDD2.n50 VDD2.n13 0.155672
R2101 VDD2.n57 VDD2.n13 0.155672
R2102 VDD2.n58 VDD2.n57 0.155672
R2103 VDD2.n58 VDD2.n9 0.155672
R2104 VDD2.n65 VDD2.n9 0.155672
R2105 VDD2.n66 VDD2.n65 0.155672
R2106 VDD2.n66 VDD2.n5 0.155672
R2107 VDD2.n75 VDD2.n5 0.155672
R2108 VDD2.n76 VDD2.n75 0.155672
R2109 VDD2.n76 VDD2.n1 0.155672
R2110 VDD2.n83 VDD2.n1 0.155672
C0 VTAIL VDD2 11.359501f
C1 VDD1 VN 0.148731f
C2 VDD2 w_n1930_n4076# 2.1462f
C3 VTAIL VP 5.7193f
C4 VTAIL B 3.47092f
C5 VP w_n1930_n4076# 3.54739f
C6 VDD1 VDD2 0.773654f
C7 B w_n1930_n4076# 8.2803f
C8 VN VDD2 6.11333f
C9 VDD1 VP 6.27198f
C10 VP VN 5.89974f
C11 VDD1 B 1.87217f
C12 B VN 0.844465f
C13 VTAIL w_n1930_n4076# 3.48569f
C14 VP VDD2 0.312824f
C15 B VDD2 1.90514f
C16 VDD1 VTAIL 11.3254f
C17 VTAIL VN 5.70461f
C18 VDD1 w_n1930_n4076# 2.11663f
C19 VN w_n1930_n4076# 3.30269f
C20 B VP 1.24431f
C21 VDD2 VSUBS 1.518311f
C22 VDD1 VSUBS 1.326086f
C23 VTAIL VSUBS 0.9212f
C24 VN VSUBS 4.7616f
C25 VP VSUBS 1.726719f
C26 B VSUBS 3.21971f
C27 w_n1930_n4076# VSUBS 96.41511f
C28 VDD2.n0 VSUBS 0.028058f
C29 VDD2.n1 VSUBS 0.025436f
C30 VDD2.n2 VSUBS 0.013668f
C31 VDD2.n3 VSUBS 0.032307f
C32 VDD2.n4 VSUBS 0.01407f
C33 VDD2.n5 VSUBS 0.025436f
C34 VDD2.n6 VSUBS 0.014472f
C35 VDD2.n7 VSUBS 0.032307f
C36 VDD2.n8 VSUBS 0.014472f
C37 VDD2.n9 VSUBS 0.025436f
C38 VDD2.n10 VSUBS 0.013668f
C39 VDD2.n11 VSUBS 0.032307f
C40 VDD2.n12 VSUBS 0.014472f
C41 VDD2.n13 VSUBS 0.025436f
C42 VDD2.n14 VSUBS 0.013668f
C43 VDD2.n15 VSUBS 0.032307f
C44 VDD2.n16 VSUBS 0.014472f
C45 VDD2.n17 VSUBS 0.025436f
C46 VDD2.n18 VSUBS 0.013668f
C47 VDD2.n19 VSUBS 0.032307f
C48 VDD2.n20 VSUBS 0.014472f
C49 VDD2.n21 VSUBS 0.025436f
C50 VDD2.n22 VSUBS 0.013668f
C51 VDD2.n23 VSUBS 0.032307f
C52 VDD2.n24 VSUBS 0.014472f
C53 VDD2.n25 VSUBS 1.68652f
C54 VDD2.n26 VSUBS 0.013668f
C55 VDD2.t0 VSUBS 0.069197f
C56 VDD2.n27 VSUBS 0.183355f
C57 VDD2.n28 VSUBS 0.020552f
C58 VDD2.n29 VSUBS 0.02423f
C59 VDD2.n30 VSUBS 0.032307f
C60 VDD2.n31 VSUBS 0.014472f
C61 VDD2.n32 VSUBS 0.013668f
C62 VDD2.n33 VSUBS 0.025436f
C63 VDD2.n34 VSUBS 0.025436f
C64 VDD2.n35 VSUBS 0.013668f
C65 VDD2.n36 VSUBS 0.014472f
C66 VDD2.n37 VSUBS 0.032307f
C67 VDD2.n38 VSUBS 0.032307f
C68 VDD2.n39 VSUBS 0.014472f
C69 VDD2.n40 VSUBS 0.013668f
C70 VDD2.n41 VSUBS 0.025436f
C71 VDD2.n42 VSUBS 0.025436f
C72 VDD2.n43 VSUBS 0.013668f
C73 VDD2.n44 VSUBS 0.014472f
C74 VDD2.n45 VSUBS 0.032307f
C75 VDD2.n46 VSUBS 0.032307f
C76 VDD2.n47 VSUBS 0.014472f
C77 VDD2.n48 VSUBS 0.013668f
C78 VDD2.n49 VSUBS 0.025436f
C79 VDD2.n50 VSUBS 0.025436f
C80 VDD2.n51 VSUBS 0.013668f
C81 VDD2.n52 VSUBS 0.014472f
C82 VDD2.n53 VSUBS 0.032307f
C83 VDD2.n54 VSUBS 0.032307f
C84 VDD2.n55 VSUBS 0.014472f
C85 VDD2.n56 VSUBS 0.013668f
C86 VDD2.n57 VSUBS 0.025436f
C87 VDD2.n58 VSUBS 0.025436f
C88 VDD2.n59 VSUBS 0.013668f
C89 VDD2.n60 VSUBS 0.014472f
C90 VDD2.n61 VSUBS 0.032307f
C91 VDD2.n62 VSUBS 0.032307f
C92 VDD2.n63 VSUBS 0.014472f
C93 VDD2.n64 VSUBS 0.013668f
C94 VDD2.n65 VSUBS 0.025436f
C95 VDD2.n66 VSUBS 0.025436f
C96 VDD2.n67 VSUBS 0.013668f
C97 VDD2.n68 VSUBS 0.013668f
C98 VDD2.n69 VSUBS 0.014472f
C99 VDD2.n70 VSUBS 0.032307f
C100 VDD2.n71 VSUBS 0.032307f
C101 VDD2.n72 VSUBS 0.032307f
C102 VDD2.n73 VSUBS 0.01407f
C103 VDD2.n74 VSUBS 0.013668f
C104 VDD2.n75 VSUBS 0.025436f
C105 VDD2.n76 VSUBS 0.025436f
C106 VDD2.n77 VSUBS 0.013668f
C107 VDD2.n78 VSUBS 0.014472f
C108 VDD2.n79 VSUBS 0.032307f
C109 VDD2.n80 VSUBS 0.078584f
C110 VDD2.n81 VSUBS 0.014472f
C111 VDD2.n82 VSUBS 0.013668f
C112 VDD2.n83 VSUBS 0.065049f
C113 VDD2.n84 VSUBS 0.058765f
C114 VDD2.t1 VSUBS 0.312362f
C115 VDD2.t3 VSUBS 0.312362f
C116 VDD2.n85 VSUBS 2.56174f
C117 VDD2.n86 VSUBS 2.45218f
C118 VDD2.n87 VSUBS 0.028058f
C119 VDD2.n88 VSUBS 0.025436f
C120 VDD2.n89 VSUBS 0.013668f
C121 VDD2.n90 VSUBS 0.032307f
C122 VDD2.n91 VSUBS 0.01407f
C123 VDD2.n92 VSUBS 0.025436f
C124 VDD2.n93 VSUBS 0.01407f
C125 VDD2.n94 VSUBS 0.013668f
C126 VDD2.n95 VSUBS 0.032307f
C127 VDD2.n96 VSUBS 0.032307f
C128 VDD2.n97 VSUBS 0.014472f
C129 VDD2.n98 VSUBS 0.025436f
C130 VDD2.n99 VSUBS 0.013668f
C131 VDD2.n100 VSUBS 0.032307f
C132 VDD2.n101 VSUBS 0.014472f
C133 VDD2.n102 VSUBS 0.025436f
C134 VDD2.n103 VSUBS 0.013668f
C135 VDD2.n104 VSUBS 0.032307f
C136 VDD2.n105 VSUBS 0.014472f
C137 VDD2.n106 VSUBS 0.025436f
C138 VDD2.n107 VSUBS 0.013668f
C139 VDD2.n108 VSUBS 0.032307f
C140 VDD2.n109 VSUBS 0.014472f
C141 VDD2.n110 VSUBS 0.025436f
C142 VDD2.n111 VSUBS 0.013668f
C143 VDD2.n112 VSUBS 0.032307f
C144 VDD2.n113 VSUBS 0.014472f
C145 VDD2.n114 VSUBS 1.68652f
C146 VDD2.n115 VSUBS 0.013668f
C147 VDD2.t4 VSUBS 0.069197f
C148 VDD2.n116 VSUBS 0.183355f
C149 VDD2.n117 VSUBS 0.020552f
C150 VDD2.n118 VSUBS 0.02423f
C151 VDD2.n119 VSUBS 0.032307f
C152 VDD2.n120 VSUBS 0.014472f
C153 VDD2.n121 VSUBS 0.013668f
C154 VDD2.n122 VSUBS 0.025436f
C155 VDD2.n123 VSUBS 0.025436f
C156 VDD2.n124 VSUBS 0.013668f
C157 VDD2.n125 VSUBS 0.014472f
C158 VDD2.n126 VSUBS 0.032307f
C159 VDD2.n127 VSUBS 0.032307f
C160 VDD2.n128 VSUBS 0.014472f
C161 VDD2.n129 VSUBS 0.013668f
C162 VDD2.n130 VSUBS 0.025436f
C163 VDD2.n131 VSUBS 0.025436f
C164 VDD2.n132 VSUBS 0.013668f
C165 VDD2.n133 VSUBS 0.014472f
C166 VDD2.n134 VSUBS 0.032307f
C167 VDD2.n135 VSUBS 0.032307f
C168 VDD2.n136 VSUBS 0.014472f
C169 VDD2.n137 VSUBS 0.013668f
C170 VDD2.n138 VSUBS 0.025436f
C171 VDD2.n139 VSUBS 0.025436f
C172 VDD2.n140 VSUBS 0.013668f
C173 VDD2.n141 VSUBS 0.014472f
C174 VDD2.n142 VSUBS 0.032307f
C175 VDD2.n143 VSUBS 0.032307f
C176 VDD2.n144 VSUBS 0.014472f
C177 VDD2.n145 VSUBS 0.013668f
C178 VDD2.n146 VSUBS 0.025436f
C179 VDD2.n147 VSUBS 0.025436f
C180 VDD2.n148 VSUBS 0.013668f
C181 VDD2.n149 VSUBS 0.014472f
C182 VDD2.n150 VSUBS 0.032307f
C183 VDD2.n151 VSUBS 0.032307f
C184 VDD2.n152 VSUBS 0.014472f
C185 VDD2.n153 VSUBS 0.013668f
C186 VDD2.n154 VSUBS 0.025436f
C187 VDD2.n155 VSUBS 0.025436f
C188 VDD2.n156 VSUBS 0.013668f
C189 VDD2.n157 VSUBS 0.014472f
C190 VDD2.n158 VSUBS 0.032307f
C191 VDD2.n159 VSUBS 0.032307f
C192 VDD2.n160 VSUBS 0.014472f
C193 VDD2.n161 VSUBS 0.013668f
C194 VDD2.n162 VSUBS 0.025436f
C195 VDD2.n163 VSUBS 0.025436f
C196 VDD2.n164 VSUBS 0.013668f
C197 VDD2.n165 VSUBS 0.014472f
C198 VDD2.n166 VSUBS 0.032307f
C199 VDD2.n167 VSUBS 0.078584f
C200 VDD2.n168 VSUBS 0.014472f
C201 VDD2.n169 VSUBS 0.013668f
C202 VDD2.n170 VSUBS 0.065049f
C203 VDD2.n171 VSUBS 0.057239f
C204 VDD2.n172 VSUBS 2.40899f
C205 VDD2.t2 VSUBS 0.312362f
C206 VDD2.t5 VSUBS 0.312362f
C207 VDD2.n173 VSUBS 2.56171f
C208 VN.n0 VSUBS 0.049687f
C209 VN.t4 VSUBS 1.8422f
C210 VN.n1 VSUBS 0.717993f
C211 VN.t5 VSUBS 1.93234f
C212 VN.n2 VSUBS 0.731823f
C213 VN.n3 VSUBS 0.206017f
C214 VN.n4 VSUBS 0.062847f
C215 VN.n5 VSUBS 0.015647f
C216 VN.t2 VSUBS 1.90802f
C217 VN.n6 VSUBS 0.721626f
C218 VN.n7 VSUBS 0.038506f
C219 VN.n8 VSUBS 0.049687f
C220 VN.t3 VSUBS 1.8422f
C221 VN.n9 VSUBS 0.717993f
C222 VN.t0 VSUBS 1.93234f
C223 VN.n10 VSUBS 0.731823f
C224 VN.n11 VSUBS 0.206017f
C225 VN.n12 VSUBS 0.062847f
C226 VN.n13 VSUBS 0.015647f
C227 VN.t1 VSUBS 1.90802f
C228 VN.n14 VSUBS 0.721626f
C229 VN.n15 VSUBS 2.28926f
C230 VTAIL.t11 VSUBS 0.345019f
C231 VTAIL.t3 VSUBS 0.345019f
C232 VTAIL.n0 VSUBS 2.67542f
C233 VTAIL.n1 VSUBS 0.758827f
C234 VTAIL.n2 VSUBS 0.030992f
C235 VTAIL.n3 VSUBS 0.028096f
C236 VTAIL.n4 VSUBS 0.015097f
C237 VTAIL.n5 VSUBS 0.035685f
C238 VTAIL.n6 VSUBS 0.015541f
C239 VTAIL.n7 VSUBS 0.028096f
C240 VTAIL.n8 VSUBS 0.015985f
C241 VTAIL.n9 VSUBS 0.035685f
C242 VTAIL.n10 VSUBS 0.015985f
C243 VTAIL.n11 VSUBS 0.028096f
C244 VTAIL.n12 VSUBS 0.015097f
C245 VTAIL.n13 VSUBS 0.035685f
C246 VTAIL.n14 VSUBS 0.015985f
C247 VTAIL.n15 VSUBS 0.028096f
C248 VTAIL.n16 VSUBS 0.015097f
C249 VTAIL.n17 VSUBS 0.035685f
C250 VTAIL.n18 VSUBS 0.015985f
C251 VTAIL.n19 VSUBS 0.028096f
C252 VTAIL.n20 VSUBS 0.015097f
C253 VTAIL.n21 VSUBS 0.035685f
C254 VTAIL.n22 VSUBS 0.015985f
C255 VTAIL.n23 VSUBS 0.028096f
C256 VTAIL.n24 VSUBS 0.015097f
C257 VTAIL.n25 VSUBS 0.035685f
C258 VTAIL.n26 VSUBS 0.015985f
C259 VTAIL.n27 VSUBS 1.86284f
C260 VTAIL.n28 VSUBS 0.015097f
C261 VTAIL.t8 VSUBS 0.076432f
C262 VTAIL.n29 VSUBS 0.202525f
C263 VTAIL.n30 VSUBS 0.022701f
C264 VTAIL.n31 VSUBS 0.026764f
C265 VTAIL.n32 VSUBS 0.035685f
C266 VTAIL.n33 VSUBS 0.015985f
C267 VTAIL.n34 VSUBS 0.015097f
C268 VTAIL.n35 VSUBS 0.028096f
C269 VTAIL.n36 VSUBS 0.028096f
C270 VTAIL.n37 VSUBS 0.015097f
C271 VTAIL.n38 VSUBS 0.015985f
C272 VTAIL.n39 VSUBS 0.035685f
C273 VTAIL.n40 VSUBS 0.035685f
C274 VTAIL.n41 VSUBS 0.015985f
C275 VTAIL.n42 VSUBS 0.015097f
C276 VTAIL.n43 VSUBS 0.028096f
C277 VTAIL.n44 VSUBS 0.028096f
C278 VTAIL.n45 VSUBS 0.015097f
C279 VTAIL.n46 VSUBS 0.015985f
C280 VTAIL.n47 VSUBS 0.035685f
C281 VTAIL.n48 VSUBS 0.035685f
C282 VTAIL.n49 VSUBS 0.015985f
C283 VTAIL.n50 VSUBS 0.015097f
C284 VTAIL.n51 VSUBS 0.028096f
C285 VTAIL.n52 VSUBS 0.028096f
C286 VTAIL.n53 VSUBS 0.015097f
C287 VTAIL.n54 VSUBS 0.015985f
C288 VTAIL.n55 VSUBS 0.035685f
C289 VTAIL.n56 VSUBS 0.035685f
C290 VTAIL.n57 VSUBS 0.015985f
C291 VTAIL.n58 VSUBS 0.015097f
C292 VTAIL.n59 VSUBS 0.028096f
C293 VTAIL.n60 VSUBS 0.028096f
C294 VTAIL.n61 VSUBS 0.015097f
C295 VTAIL.n62 VSUBS 0.015985f
C296 VTAIL.n63 VSUBS 0.035685f
C297 VTAIL.n64 VSUBS 0.035685f
C298 VTAIL.n65 VSUBS 0.015985f
C299 VTAIL.n66 VSUBS 0.015097f
C300 VTAIL.n67 VSUBS 0.028096f
C301 VTAIL.n68 VSUBS 0.028096f
C302 VTAIL.n69 VSUBS 0.015097f
C303 VTAIL.n70 VSUBS 0.015097f
C304 VTAIL.n71 VSUBS 0.015985f
C305 VTAIL.n72 VSUBS 0.035685f
C306 VTAIL.n73 VSUBS 0.035685f
C307 VTAIL.n74 VSUBS 0.035685f
C308 VTAIL.n75 VSUBS 0.015541f
C309 VTAIL.n76 VSUBS 0.015097f
C310 VTAIL.n77 VSUBS 0.028096f
C311 VTAIL.n78 VSUBS 0.028096f
C312 VTAIL.n79 VSUBS 0.015097f
C313 VTAIL.n80 VSUBS 0.015985f
C314 VTAIL.n81 VSUBS 0.035685f
C315 VTAIL.n82 VSUBS 0.0868f
C316 VTAIL.n83 VSUBS 0.015985f
C317 VTAIL.n84 VSUBS 0.015097f
C318 VTAIL.n85 VSUBS 0.07185f
C319 VTAIL.n86 VSUBS 0.043872f
C320 VTAIL.n87 VSUBS 0.210916f
C321 VTAIL.t7 VSUBS 0.345019f
C322 VTAIL.t10 VSUBS 0.345019f
C323 VTAIL.n88 VSUBS 2.67542f
C324 VTAIL.n89 VSUBS 2.51618f
C325 VTAIL.t0 VSUBS 0.345019f
C326 VTAIL.t2 VSUBS 0.345019f
C327 VTAIL.n90 VSUBS 2.67544f
C328 VTAIL.n91 VSUBS 2.51617f
C329 VTAIL.n92 VSUBS 0.030992f
C330 VTAIL.n93 VSUBS 0.028096f
C331 VTAIL.n94 VSUBS 0.015097f
C332 VTAIL.n95 VSUBS 0.035685f
C333 VTAIL.n96 VSUBS 0.015541f
C334 VTAIL.n97 VSUBS 0.028096f
C335 VTAIL.n98 VSUBS 0.015541f
C336 VTAIL.n99 VSUBS 0.015097f
C337 VTAIL.n100 VSUBS 0.035685f
C338 VTAIL.n101 VSUBS 0.035685f
C339 VTAIL.n102 VSUBS 0.015985f
C340 VTAIL.n103 VSUBS 0.028096f
C341 VTAIL.n104 VSUBS 0.015097f
C342 VTAIL.n105 VSUBS 0.035685f
C343 VTAIL.n106 VSUBS 0.015985f
C344 VTAIL.n107 VSUBS 0.028096f
C345 VTAIL.n108 VSUBS 0.015097f
C346 VTAIL.n109 VSUBS 0.035685f
C347 VTAIL.n110 VSUBS 0.015985f
C348 VTAIL.n111 VSUBS 0.028096f
C349 VTAIL.n112 VSUBS 0.015097f
C350 VTAIL.n113 VSUBS 0.035685f
C351 VTAIL.n114 VSUBS 0.015985f
C352 VTAIL.n115 VSUBS 0.028096f
C353 VTAIL.n116 VSUBS 0.015097f
C354 VTAIL.n117 VSUBS 0.035685f
C355 VTAIL.n118 VSUBS 0.015985f
C356 VTAIL.n119 VSUBS 1.86284f
C357 VTAIL.n120 VSUBS 0.015097f
C358 VTAIL.t1 VSUBS 0.076432f
C359 VTAIL.n121 VSUBS 0.202525f
C360 VTAIL.n122 VSUBS 0.022701f
C361 VTAIL.n123 VSUBS 0.026764f
C362 VTAIL.n124 VSUBS 0.035685f
C363 VTAIL.n125 VSUBS 0.015985f
C364 VTAIL.n126 VSUBS 0.015097f
C365 VTAIL.n127 VSUBS 0.028096f
C366 VTAIL.n128 VSUBS 0.028096f
C367 VTAIL.n129 VSUBS 0.015097f
C368 VTAIL.n130 VSUBS 0.015985f
C369 VTAIL.n131 VSUBS 0.035685f
C370 VTAIL.n132 VSUBS 0.035685f
C371 VTAIL.n133 VSUBS 0.015985f
C372 VTAIL.n134 VSUBS 0.015097f
C373 VTAIL.n135 VSUBS 0.028096f
C374 VTAIL.n136 VSUBS 0.028096f
C375 VTAIL.n137 VSUBS 0.015097f
C376 VTAIL.n138 VSUBS 0.015985f
C377 VTAIL.n139 VSUBS 0.035685f
C378 VTAIL.n140 VSUBS 0.035685f
C379 VTAIL.n141 VSUBS 0.015985f
C380 VTAIL.n142 VSUBS 0.015097f
C381 VTAIL.n143 VSUBS 0.028096f
C382 VTAIL.n144 VSUBS 0.028096f
C383 VTAIL.n145 VSUBS 0.015097f
C384 VTAIL.n146 VSUBS 0.015985f
C385 VTAIL.n147 VSUBS 0.035685f
C386 VTAIL.n148 VSUBS 0.035685f
C387 VTAIL.n149 VSUBS 0.015985f
C388 VTAIL.n150 VSUBS 0.015097f
C389 VTAIL.n151 VSUBS 0.028096f
C390 VTAIL.n152 VSUBS 0.028096f
C391 VTAIL.n153 VSUBS 0.015097f
C392 VTAIL.n154 VSUBS 0.015985f
C393 VTAIL.n155 VSUBS 0.035685f
C394 VTAIL.n156 VSUBS 0.035685f
C395 VTAIL.n157 VSUBS 0.015985f
C396 VTAIL.n158 VSUBS 0.015097f
C397 VTAIL.n159 VSUBS 0.028096f
C398 VTAIL.n160 VSUBS 0.028096f
C399 VTAIL.n161 VSUBS 0.015097f
C400 VTAIL.n162 VSUBS 0.015985f
C401 VTAIL.n163 VSUBS 0.035685f
C402 VTAIL.n164 VSUBS 0.035685f
C403 VTAIL.n165 VSUBS 0.015985f
C404 VTAIL.n166 VSUBS 0.015097f
C405 VTAIL.n167 VSUBS 0.028096f
C406 VTAIL.n168 VSUBS 0.028096f
C407 VTAIL.n169 VSUBS 0.015097f
C408 VTAIL.n170 VSUBS 0.015985f
C409 VTAIL.n171 VSUBS 0.035685f
C410 VTAIL.n172 VSUBS 0.0868f
C411 VTAIL.n173 VSUBS 0.015985f
C412 VTAIL.n174 VSUBS 0.015097f
C413 VTAIL.n175 VSUBS 0.07185f
C414 VTAIL.n176 VSUBS 0.043872f
C415 VTAIL.n177 VSUBS 0.210916f
C416 VTAIL.t9 VSUBS 0.345019f
C417 VTAIL.t6 VSUBS 0.345019f
C418 VTAIL.n178 VSUBS 2.67544f
C419 VTAIL.n179 VSUBS 0.823782f
C420 VTAIL.n180 VSUBS 0.030992f
C421 VTAIL.n181 VSUBS 0.028096f
C422 VTAIL.n182 VSUBS 0.015097f
C423 VTAIL.n183 VSUBS 0.035685f
C424 VTAIL.n184 VSUBS 0.015541f
C425 VTAIL.n185 VSUBS 0.028096f
C426 VTAIL.n186 VSUBS 0.015541f
C427 VTAIL.n187 VSUBS 0.015097f
C428 VTAIL.n188 VSUBS 0.035685f
C429 VTAIL.n189 VSUBS 0.035685f
C430 VTAIL.n190 VSUBS 0.015985f
C431 VTAIL.n191 VSUBS 0.028096f
C432 VTAIL.n192 VSUBS 0.015097f
C433 VTAIL.n193 VSUBS 0.035685f
C434 VTAIL.n194 VSUBS 0.015985f
C435 VTAIL.n195 VSUBS 0.028096f
C436 VTAIL.n196 VSUBS 0.015097f
C437 VTAIL.n197 VSUBS 0.035685f
C438 VTAIL.n198 VSUBS 0.015985f
C439 VTAIL.n199 VSUBS 0.028096f
C440 VTAIL.n200 VSUBS 0.015097f
C441 VTAIL.n201 VSUBS 0.035685f
C442 VTAIL.n202 VSUBS 0.015985f
C443 VTAIL.n203 VSUBS 0.028096f
C444 VTAIL.n204 VSUBS 0.015097f
C445 VTAIL.n205 VSUBS 0.035685f
C446 VTAIL.n206 VSUBS 0.015985f
C447 VTAIL.n207 VSUBS 1.86284f
C448 VTAIL.n208 VSUBS 0.015097f
C449 VTAIL.t5 VSUBS 0.076432f
C450 VTAIL.n209 VSUBS 0.202525f
C451 VTAIL.n210 VSUBS 0.022701f
C452 VTAIL.n211 VSUBS 0.026764f
C453 VTAIL.n212 VSUBS 0.035685f
C454 VTAIL.n213 VSUBS 0.015985f
C455 VTAIL.n214 VSUBS 0.015097f
C456 VTAIL.n215 VSUBS 0.028096f
C457 VTAIL.n216 VSUBS 0.028096f
C458 VTAIL.n217 VSUBS 0.015097f
C459 VTAIL.n218 VSUBS 0.015985f
C460 VTAIL.n219 VSUBS 0.035685f
C461 VTAIL.n220 VSUBS 0.035685f
C462 VTAIL.n221 VSUBS 0.015985f
C463 VTAIL.n222 VSUBS 0.015097f
C464 VTAIL.n223 VSUBS 0.028096f
C465 VTAIL.n224 VSUBS 0.028096f
C466 VTAIL.n225 VSUBS 0.015097f
C467 VTAIL.n226 VSUBS 0.015985f
C468 VTAIL.n227 VSUBS 0.035685f
C469 VTAIL.n228 VSUBS 0.035685f
C470 VTAIL.n229 VSUBS 0.015985f
C471 VTAIL.n230 VSUBS 0.015097f
C472 VTAIL.n231 VSUBS 0.028096f
C473 VTAIL.n232 VSUBS 0.028096f
C474 VTAIL.n233 VSUBS 0.015097f
C475 VTAIL.n234 VSUBS 0.015985f
C476 VTAIL.n235 VSUBS 0.035685f
C477 VTAIL.n236 VSUBS 0.035685f
C478 VTAIL.n237 VSUBS 0.015985f
C479 VTAIL.n238 VSUBS 0.015097f
C480 VTAIL.n239 VSUBS 0.028096f
C481 VTAIL.n240 VSUBS 0.028096f
C482 VTAIL.n241 VSUBS 0.015097f
C483 VTAIL.n242 VSUBS 0.015985f
C484 VTAIL.n243 VSUBS 0.035685f
C485 VTAIL.n244 VSUBS 0.035685f
C486 VTAIL.n245 VSUBS 0.015985f
C487 VTAIL.n246 VSUBS 0.015097f
C488 VTAIL.n247 VSUBS 0.028096f
C489 VTAIL.n248 VSUBS 0.028096f
C490 VTAIL.n249 VSUBS 0.015097f
C491 VTAIL.n250 VSUBS 0.015985f
C492 VTAIL.n251 VSUBS 0.035685f
C493 VTAIL.n252 VSUBS 0.035685f
C494 VTAIL.n253 VSUBS 0.015985f
C495 VTAIL.n254 VSUBS 0.015097f
C496 VTAIL.n255 VSUBS 0.028096f
C497 VTAIL.n256 VSUBS 0.028096f
C498 VTAIL.n257 VSUBS 0.015097f
C499 VTAIL.n258 VSUBS 0.015985f
C500 VTAIL.n259 VSUBS 0.035685f
C501 VTAIL.n260 VSUBS 0.0868f
C502 VTAIL.n261 VSUBS 0.015985f
C503 VTAIL.n262 VSUBS 0.015097f
C504 VTAIL.n263 VSUBS 0.07185f
C505 VTAIL.n264 VSUBS 0.043872f
C506 VTAIL.n265 VSUBS 1.80965f
C507 VTAIL.n266 VSUBS 0.030992f
C508 VTAIL.n267 VSUBS 0.028096f
C509 VTAIL.n268 VSUBS 0.015097f
C510 VTAIL.n269 VSUBS 0.035685f
C511 VTAIL.n270 VSUBS 0.015541f
C512 VTAIL.n271 VSUBS 0.028096f
C513 VTAIL.n272 VSUBS 0.015985f
C514 VTAIL.n273 VSUBS 0.035685f
C515 VTAIL.n274 VSUBS 0.015985f
C516 VTAIL.n275 VSUBS 0.028096f
C517 VTAIL.n276 VSUBS 0.015097f
C518 VTAIL.n277 VSUBS 0.035685f
C519 VTAIL.n278 VSUBS 0.015985f
C520 VTAIL.n279 VSUBS 0.028096f
C521 VTAIL.n280 VSUBS 0.015097f
C522 VTAIL.n281 VSUBS 0.035685f
C523 VTAIL.n282 VSUBS 0.015985f
C524 VTAIL.n283 VSUBS 0.028096f
C525 VTAIL.n284 VSUBS 0.015097f
C526 VTAIL.n285 VSUBS 0.035685f
C527 VTAIL.n286 VSUBS 0.015985f
C528 VTAIL.n287 VSUBS 0.028096f
C529 VTAIL.n288 VSUBS 0.015097f
C530 VTAIL.n289 VSUBS 0.035685f
C531 VTAIL.n290 VSUBS 0.015985f
C532 VTAIL.n291 VSUBS 1.86284f
C533 VTAIL.n292 VSUBS 0.015097f
C534 VTAIL.t4 VSUBS 0.076432f
C535 VTAIL.n293 VSUBS 0.202525f
C536 VTAIL.n294 VSUBS 0.022701f
C537 VTAIL.n295 VSUBS 0.026764f
C538 VTAIL.n296 VSUBS 0.035685f
C539 VTAIL.n297 VSUBS 0.015985f
C540 VTAIL.n298 VSUBS 0.015097f
C541 VTAIL.n299 VSUBS 0.028096f
C542 VTAIL.n300 VSUBS 0.028096f
C543 VTAIL.n301 VSUBS 0.015097f
C544 VTAIL.n302 VSUBS 0.015985f
C545 VTAIL.n303 VSUBS 0.035685f
C546 VTAIL.n304 VSUBS 0.035685f
C547 VTAIL.n305 VSUBS 0.015985f
C548 VTAIL.n306 VSUBS 0.015097f
C549 VTAIL.n307 VSUBS 0.028096f
C550 VTAIL.n308 VSUBS 0.028096f
C551 VTAIL.n309 VSUBS 0.015097f
C552 VTAIL.n310 VSUBS 0.015985f
C553 VTAIL.n311 VSUBS 0.035685f
C554 VTAIL.n312 VSUBS 0.035685f
C555 VTAIL.n313 VSUBS 0.015985f
C556 VTAIL.n314 VSUBS 0.015097f
C557 VTAIL.n315 VSUBS 0.028096f
C558 VTAIL.n316 VSUBS 0.028096f
C559 VTAIL.n317 VSUBS 0.015097f
C560 VTAIL.n318 VSUBS 0.015985f
C561 VTAIL.n319 VSUBS 0.035685f
C562 VTAIL.n320 VSUBS 0.035685f
C563 VTAIL.n321 VSUBS 0.015985f
C564 VTAIL.n322 VSUBS 0.015097f
C565 VTAIL.n323 VSUBS 0.028096f
C566 VTAIL.n324 VSUBS 0.028096f
C567 VTAIL.n325 VSUBS 0.015097f
C568 VTAIL.n326 VSUBS 0.015985f
C569 VTAIL.n327 VSUBS 0.035685f
C570 VTAIL.n328 VSUBS 0.035685f
C571 VTAIL.n329 VSUBS 0.015985f
C572 VTAIL.n330 VSUBS 0.015097f
C573 VTAIL.n331 VSUBS 0.028096f
C574 VTAIL.n332 VSUBS 0.028096f
C575 VTAIL.n333 VSUBS 0.015097f
C576 VTAIL.n334 VSUBS 0.015097f
C577 VTAIL.n335 VSUBS 0.015985f
C578 VTAIL.n336 VSUBS 0.035685f
C579 VTAIL.n337 VSUBS 0.035685f
C580 VTAIL.n338 VSUBS 0.035685f
C581 VTAIL.n339 VSUBS 0.015541f
C582 VTAIL.n340 VSUBS 0.015097f
C583 VTAIL.n341 VSUBS 0.028096f
C584 VTAIL.n342 VSUBS 0.028096f
C585 VTAIL.n343 VSUBS 0.015097f
C586 VTAIL.n344 VSUBS 0.015985f
C587 VTAIL.n345 VSUBS 0.035685f
C588 VTAIL.n346 VSUBS 0.0868f
C589 VTAIL.n347 VSUBS 0.015985f
C590 VTAIL.n348 VSUBS 0.015097f
C591 VTAIL.n349 VSUBS 0.07185f
C592 VTAIL.n350 VSUBS 0.043872f
C593 VTAIL.n351 VSUBS 1.78097f
C594 VDD1.n0 VSUBS 0.028067f
C595 VDD1.n1 VSUBS 0.025444f
C596 VDD1.n2 VSUBS 0.013673f
C597 VDD1.n3 VSUBS 0.032317f
C598 VDD1.n4 VSUBS 0.014075f
C599 VDD1.n5 VSUBS 0.025444f
C600 VDD1.n6 VSUBS 0.014075f
C601 VDD1.n7 VSUBS 0.013673f
C602 VDD1.n8 VSUBS 0.032317f
C603 VDD1.n9 VSUBS 0.032317f
C604 VDD1.n10 VSUBS 0.014477f
C605 VDD1.n11 VSUBS 0.025444f
C606 VDD1.n12 VSUBS 0.013673f
C607 VDD1.n13 VSUBS 0.032317f
C608 VDD1.n14 VSUBS 0.014477f
C609 VDD1.n15 VSUBS 0.025444f
C610 VDD1.n16 VSUBS 0.013673f
C611 VDD1.n17 VSUBS 0.032317f
C612 VDD1.n18 VSUBS 0.014477f
C613 VDD1.n19 VSUBS 0.025444f
C614 VDD1.n20 VSUBS 0.013673f
C615 VDD1.n21 VSUBS 0.032317f
C616 VDD1.n22 VSUBS 0.014477f
C617 VDD1.n23 VSUBS 0.025444f
C618 VDD1.n24 VSUBS 0.013673f
C619 VDD1.n25 VSUBS 0.032317f
C620 VDD1.n26 VSUBS 0.014477f
C621 VDD1.n27 VSUBS 1.68703f
C622 VDD1.n28 VSUBS 0.013673f
C623 VDD1.t0 VSUBS 0.069218f
C624 VDD1.n29 VSUBS 0.183412f
C625 VDD1.n30 VSUBS 0.020559f
C626 VDD1.n31 VSUBS 0.024238f
C627 VDD1.n32 VSUBS 0.032317f
C628 VDD1.n33 VSUBS 0.014477f
C629 VDD1.n34 VSUBS 0.013673f
C630 VDD1.n35 VSUBS 0.025444f
C631 VDD1.n36 VSUBS 0.025444f
C632 VDD1.n37 VSUBS 0.013673f
C633 VDD1.n38 VSUBS 0.014477f
C634 VDD1.n39 VSUBS 0.032317f
C635 VDD1.n40 VSUBS 0.032317f
C636 VDD1.n41 VSUBS 0.014477f
C637 VDD1.n42 VSUBS 0.013673f
C638 VDD1.n43 VSUBS 0.025444f
C639 VDD1.n44 VSUBS 0.025444f
C640 VDD1.n45 VSUBS 0.013673f
C641 VDD1.n46 VSUBS 0.014477f
C642 VDD1.n47 VSUBS 0.032317f
C643 VDD1.n48 VSUBS 0.032317f
C644 VDD1.n49 VSUBS 0.014477f
C645 VDD1.n50 VSUBS 0.013673f
C646 VDD1.n51 VSUBS 0.025444f
C647 VDD1.n52 VSUBS 0.025444f
C648 VDD1.n53 VSUBS 0.013673f
C649 VDD1.n54 VSUBS 0.014477f
C650 VDD1.n55 VSUBS 0.032317f
C651 VDD1.n56 VSUBS 0.032317f
C652 VDD1.n57 VSUBS 0.014477f
C653 VDD1.n58 VSUBS 0.013673f
C654 VDD1.n59 VSUBS 0.025444f
C655 VDD1.n60 VSUBS 0.025444f
C656 VDD1.n61 VSUBS 0.013673f
C657 VDD1.n62 VSUBS 0.014477f
C658 VDD1.n63 VSUBS 0.032317f
C659 VDD1.n64 VSUBS 0.032317f
C660 VDD1.n65 VSUBS 0.014477f
C661 VDD1.n66 VSUBS 0.013673f
C662 VDD1.n67 VSUBS 0.025444f
C663 VDD1.n68 VSUBS 0.025444f
C664 VDD1.n69 VSUBS 0.013673f
C665 VDD1.n70 VSUBS 0.014477f
C666 VDD1.n71 VSUBS 0.032317f
C667 VDD1.n72 VSUBS 0.032317f
C668 VDD1.n73 VSUBS 0.014477f
C669 VDD1.n74 VSUBS 0.013673f
C670 VDD1.n75 VSUBS 0.025444f
C671 VDD1.n76 VSUBS 0.025444f
C672 VDD1.n77 VSUBS 0.013673f
C673 VDD1.n78 VSUBS 0.014477f
C674 VDD1.n79 VSUBS 0.032317f
C675 VDD1.n80 VSUBS 0.078608f
C676 VDD1.n81 VSUBS 0.014477f
C677 VDD1.n82 VSUBS 0.013673f
C678 VDD1.n83 VSUBS 0.06507f
C679 VDD1.n84 VSUBS 0.059153f
C680 VDD1.n85 VSUBS 0.028067f
C681 VDD1.n86 VSUBS 0.025444f
C682 VDD1.n87 VSUBS 0.013673f
C683 VDD1.n88 VSUBS 0.032317f
C684 VDD1.n89 VSUBS 0.014075f
C685 VDD1.n90 VSUBS 0.025444f
C686 VDD1.n91 VSUBS 0.014477f
C687 VDD1.n92 VSUBS 0.032317f
C688 VDD1.n93 VSUBS 0.014477f
C689 VDD1.n94 VSUBS 0.025444f
C690 VDD1.n95 VSUBS 0.013673f
C691 VDD1.n96 VSUBS 0.032317f
C692 VDD1.n97 VSUBS 0.014477f
C693 VDD1.n98 VSUBS 0.025444f
C694 VDD1.n99 VSUBS 0.013673f
C695 VDD1.n100 VSUBS 0.032317f
C696 VDD1.n101 VSUBS 0.014477f
C697 VDD1.n102 VSUBS 0.025444f
C698 VDD1.n103 VSUBS 0.013673f
C699 VDD1.n104 VSUBS 0.032317f
C700 VDD1.n105 VSUBS 0.014477f
C701 VDD1.n106 VSUBS 0.025444f
C702 VDD1.n107 VSUBS 0.013673f
C703 VDD1.n108 VSUBS 0.032317f
C704 VDD1.n109 VSUBS 0.014477f
C705 VDD1.n110 VSUBS 1.68703f
C706 VDD1.n111 VSUBS 0.013673f
C707 VDD1.t4 VSUBS 0.069218f
C708 VDD1.n112 VSUBS 0.183412f
C709 VDD1.n113 VSUBS 0.020559f
C710 VDD1.n114 VSUBS 0.024238f
C711 VDD1.n115 VSUBS 0.032317f
C712 VDD1.n116 VSUBS 0.014477f
C713 VDD1.n117 VSUBS 0.013673f
C714 VDD1.n118 VSUBS 0.025444f
C715 VDD1.n119 VSUBS 0.025444f
C716 VDD1.n120 VSUBS 0.013673f
C717 VDD1.n121 VSUBS 0.014477f
C718 VDD1.n122 VSUBS 0.032317f
C719 VDD1.n123 VSUBS 0.032317f
C720 VDD1.n124 VSUBS 0.014477f
C721 VDD1.n125 VSUBS 0.013673f
C722 VDD1.n126 VSUBS 0.025444f
C723 VDD1.n127 VSUBS 0.025444f
C724 VDD1.n128 VSUBS 0.013673f
C725 VDD1.n129 VSUBS 0.014477f
C726 VDD1.n130 VSUBS 0.032317f
C727 VDD1.n131 VSUBS 0.032317f
C728 VDD1.n132 VSUBS 0.014477f
C729 VDD1.n133 VSUBS 0.013673f
C730 VDD1.n134 VSUBS 0.025444f
C731 VDD1.n135 VSUBS 0.025444f
C732 VDD1.n136 VSUBS 0.013673f
C733 VDD1.n137 VSUBS 0.014477f
C734 VDD1.n138 VSUBS 0.032317f
C735 VDD1.n139 VSUBS 0.032317f
C736 VDD1.n140 VSUBS 0.014477f
C737 VDD1.n141 VSUBS 0.013673f
C738 VDD1.n142 VSUBS 0.025444f
C739 VDD1.n143 VSUBS 0.025444f
C740 VDD1.n144 VSUBS 0.013673f
C741 VDD1.n145 VSUBS 0.014477f
C742 VDD1.n146 VSUBS 0.032317f
C743 VDD1.n147 VSUBS 0.032317f
C744 VDD1.n148 VSUBS 0.014477f
C745 VDD1.n149 VSUBS 0.013673f
C746 VDD1.n150 VSUBS 0.025444f
C747 VDD1.n151 VSUBS 0.025444f
C748 VDD1.n152 VSUBS 0.013673f
C749 VDD1.n153 VSUBS 0.013673f
C750 VDD1.n154 VSUBS 0.014477f
C751 VDD1.n155 VSUBS 0.032317f
C752 VDD1.n156 VSUBS 0.032317f
C753 VDD1.n157 VSUBS 0.032317f
C754 VDD1.n158 VSUBS 0.014075f
C755 VDD1.n159 VSUBS 0.013673f
C756 VDD1.n160 VSUBS 0.025444f
C757 VDD1.n161 VSUBS 0.025444f
C758 VDD1.n162 VSUBS 0.013673f
C759 VDD1.n163 VSUBS 0.014477f
C760 VDD1.n164 VSUBS 0.032317f
C761 VDD1.n165 VSUBS 0.078608f
C762 VDD1.n166 VSUBS 0.014477f
C763 VDD1.n167 VSUBS 0.013673f
C764 VDD1.n168 VSUBS 0.06507f
C765 VDD1.n169 VSUBS 0.058783f
C766 VDD1.t1 VSUBS 0.312458f
C767 VDD1.t5 VSUBS 0.312458f
C768 VDD1.n170 VSUBS 2.56253f
C769 VDD1.n171 VSUBS 2.53667f
C770 VDD1.t3 VSUBS 0.312458f
C771 VDD1.t2 VSUBS 0.312458f
C772 VDD1.n172 VSUBS 2.5609f
C773 VDD1.n173 VSUBS 2.88744f
C774 VP.n0 VSUBS 0.050802f
C775 VP.t0 VSUBS 1.88356f
C776 VP.n1 VSUBS 0.688123f
C777 VP.n2 VSUBS 0.050802f
C778 VP.n3 VSUBS 0.050802f
C779 VP.t5 VSUBS 1.95085f
C780 VP.t4 VSUBS 1.88356f
C781 VP.n4 VSUBS 0.734111f
C782 VP.t1 VSUBS 1.97572f
C783 VP.n5 VSUBS 0.748251f
C784 VP.n6 VSUBS 0.210642f
C785 VP.n7 VSUBS 0.064258f
C786 VP.n8 VSUBS 0.015998f
C787 VP.n9 VSUBS 0.737826f
C788 VP.n10 VSUBS 2.30741f
C789 VP.n11 VSUBS 2.34854f
C790 VP.t3 VSUBS 1.95085f
C791 VP.n12 VSUBS 0.737826f
C792 VP.n13 VSUBS 0.015998f
C793 VP.n14 VSUBS 0.064258f
C794 VP.n15 VSUBS 0.050802f
C795 VP.n16 VSUBS 0.050802f
C796 VP.n17 VSUBS 0.064258f
C797 VP.n18 VSUBS 0.015998f
C798 VP.t2 VSUBS 1.95085f
C799 VP.n19 VSUBS 0.737826f
C800 VP.n20 VSUBS 0.03937f
C801 B.n0 VSUBS 0.004326f
C802 B.n1 VSUBS 0.004326f
C803 B.n2 VSUBS 0.006841f
C804 B.n3 VSUBS 0.006841f
C805 B.n4 VSUBS 0.006841f
C806 B.n5 VSUBS 0.006841f
C807 B.n6 VSUBS 0.006841f
C808 B.n7 VSUBS 0.006841f
C809 B.n8 VSUBS 0.006841f
C810 B.n9 VSUBS 0.006841f
C811 B.n10 VSUBS 0.006841f
C812 B.n11 VSUBS 0.006841f
C813 B.n12 VSUBS 0.006841f
C814 B.n13 VSUBS 0.016752f
C815 B.n14 VSUBS 0.006841f
C816 B.n15 VSUBS 0.006841f
C817 B.n16 VSUBS 0.006841f
C818 B.n17 VSUBS 0.006841f
C819 B.n18 VSUBS 0.006841f
C820 B.n19 VSUBS 0.006841f
C821 B.n20 VSUBS 0.006841f
C822 B.n21 VSUBS 0.006841f
C823 B.n22 VSUBS 0.006841f
C824 B.n23 VSUBS 0.006841f
C825 B.n24 VSUBS 0.006841f
C826 B.n25 VSUBS 0.006841f
C827 B.n26 VSUBS 0.006841f
C828 B.n27 VSUBS 0.006841f
C829 B.n28 VSUBS 0.006841f
C830 B.n29 VSUBS 0.006841f
C831 B.n30 VSUBS 0.006841f
C832 B.n31 VSUBS 0.006841f
C833 B.n32 VSUBS 0.006841f
C834 B.n33 VSUBS 0.006841f
C835 B.n34 VSUBS 0.006841f
C836 B.n35 VSUBS 0.006841f
C837 B.n36 VSUBS 0.006841f
C838 B.n37 VSUBS 0.006841f
C839 B.n38 VSUBS 0.006841f
C840 B.n39 VSUBS 0.006841f
C841 B.t11 VSUBS 0.285778f
C842 B.t10 VSUBS 0.299604f
C843 B.t9 VSUBS 0.544586f
C844 B.n40 VSUBS 0.395072f
C845 B.n41 VSUBS 0.28467f
C846 B.n42 VSUBS 0.006841f
C847 B.n43 VSUBS 0.006841f
C848 B.n44 VSUBS 0.006841f
C849 B.n45 VSUBS 0.006841f
C850 B.t5 VSUBS 0.285781f
C851 B.t4 VSUBS 0.299607f
C852 B.t3 VSUBS 0.544586f
C853 B.n46 VSUBS 0.395069f
C854 B.n47 VSUBS 0.284667f
C855 B.n48 VSUBS 0.015851f
C856 B.n49 VSUBS 0.006841f
C857 B.n50 VSUBS 0.006841f
C858 B.n51 VSUBS 0.006841f
C859 B.n52 VSUBS 0.006841f
C860 B.n53 VSUBS 0.006841f
C861 B.n54 VSUBS 0.006841f
C862 B.n55 VSUBS 0.006841f
C863 B.n56 VSUBS 0.006841f
C864 B.n57 VSUBS 0.006841f
C865 B.n58 VSUBS 0.006841f
C866 B.n59 VSUBS 0.006841f
C867 B.n60 VSUBS 0.006841f
C868 B.n61 VSUBS 0.006841f
C869 B.n62 VSUBS 0.006841f
C870 B.n63 VSUBS 0.006841f
C871 B.n64 VSUBS 0.006841f
C872 B.n65 VSUBS 0.006841f
C873 B.n66 VSUBS 0.006841f
C874 B.n67 VSUBS 0.006841f
C875 B.n68 VSUBS 0.006841f
C876 B.n69 VSUBS 0.006841f
C877 B.n70 VSUBS 0.006841f
C878 B.n71 VSUBS 0.006841f
C879 B.n72 VSUBS 0.006841f
C880 B.n73 VSUBS 0.006841f
C881 B.n74 VSUBS 0.015951f
C882 B.n75 VSUBS 0.006841f
C883 B.n76 VSUBS 0.006841f
C884 B.n77 VSUBS 0.006841f
C885 B.n78 VSUBS 0.006841f
C886 B.n79 VSUBS 0.006841f
C887 B.n80 VSUBS 0.006841f
C888 B.n81 VSUBS 0.006841f
C889 B.n82 VSUBS 0.006841f
C890 B.n83 VSUBS 0.006841f
C891 B.n84 VSUBS 0.006841f
C892 B.n85 VSUBS 0.006841f
C893 B.n86 VSUBS 0.006841f
C894 B.n87 VSUBS 0.006841f
C895 B.n88 VSUBS 0.006841f
C896 B.n89 VSUBS 0.006841f
C897 B.n90 VSUBS 0.006841f
C898 B.n91 VSUBS 0.006841f
C899 B.n92 VSUBS 0.006841f
C900 B.n93 VSUBS 0.006841f
C901 B.n94 VSUBS 0.006841f
C902 B.n95 VSUBS 0.006841f
C903 B.n96 VSUBS 0.006841f
C904 B.n97 VSUBS 0.016752f
C905 B.n98 VSUBS 0.006841f
C906 B.n99 VSUBS 0.006841f
C907 B.n100 VSUBS 0.006841f
C908 B.n101 VSUBS 0.006841f
C909 B.n102 VSUBS 0.006841f
C910 B.n103 VSUBS 0.006841f
C911 B.n104 VSUBS 0.006841f
C912 B.n105 VSUBS 0.006841f
C913 B.n106 VSUBS 0.006841f
C914 B.n107 VSUBS 0.006841f
C915 B.n108 VSUBS 0.006841f
C916 B.n109 VSUBS 0.006841f
C917 B.n110 VSUBS 0.006841f
C918 B.n111 VSUBS 0.006841f
C919 B.n112 VSUBS 0.006841f
C920 B.n113 VSUBS 0.006841f
C921 B.n114 VSUBS 0.006841f
C922 B.n115 VSUBS 0.006841f
C923 B.n116 VSUBS 0.006841f
C924 B.n117 VSUBS 0.006841f
C925 B.n118 VSUBS 0.006841f
C926 B.n119 VSUBS 0.006841f
C927 B.n120 VSUBS 0.006841f
C928 B.n121 VSUBS 0.006841f
C929 B.n122 VSUBS 0.006841f
C930 B.n123 VSUBS 0.006841f
C931 B.t1 VSUBS 0.285781f
C932 B.t2 VSUBS 0.299607f
C933 B.t0 VSUBS 0.544586f
C934 B.n124 VSUBS 0.395069f
C935 B.n125 VSUBS 0.284667f
C936 B.n126 VSUBS 0.006841f
C937 B.n127 VSUBS 0.006841f
C938 B.n128 VSUBS 0.006841f
C939 B.n129 VSUBS 0.006841f
C940 B.t7 VSUBS 0.285778f
C941 B.t8 VSUBS 0.299604f
C942 B.t6 VSUBS 0.544586f
C943 B.n130 VSUBS 0.395072f
C944 B.n131 VSUBS 0.28467f
C945 B.n132 VSUBS 0.015851f
C946 B.n133 VSUBS 0.006841f
C947 B.n134 VSUBS 0.006841f
C948 B.n135 VSUBS 0.006841f
C949 B.n136 VSUBS 0.006841f
C950 B.n137 VSUBS 0.006841f
C951 B.n138 VSUBS 0.006841f
C952 B.n139 VSUBS 0.006841f
C953 B.n140 VSUBS 0.006841f
C954 B.n141 VSUBS 0.006841f
C955 B.n142 VSUBS 0.006841f
C956 B.n143 VSUBS 0.006841f
C957 B.n144 VSUBS 0.006841f
C958 B.n145 VSUBS 0.006841f
C959 B.n146 VSUBS 0.006841f
C960 B.n147 VSUBS 0.006841f
C961 B.n148 VSUBS 0.006841f
C962 B.n149 VSUBS 0.006841f
C963 B.n150 VSUBS 0.006841f
C964 B.n151 VSUBS 0.006841f
C965 B.n152 VSUBS 0.006841f
C966 B.n153 VSUBS 0.006841f
C967 B.n154 VSUBS 0.006841f
C968 B.n155 VSUBS 0.006841f
C969 B.n156 VSUBS 0.006841f
C970 B.n157 VSUBS 0.006841f
C971 B.n158 VSUBS 0.016752f
C972 B.n159 VSUBS 0.006841f
C973 B.n160 VSUBS 0.006841f
C974 B.n161 VSUBS 0.006841f
C975 B.n162 VSUBS 0.006841f
C976 B.n163 VSUBS 0.006841f
C977 B.n164 VSUBS 0.006841f
C978 B.n165 VSUBS 0.006841f
C979 B.n166 VSUBS 0.006841f
C980 B.n167 VSUBS 0.006841f
C981 B.n168 VSUBS 0.006841f
C982 B.n169 VSUBS 0.006841f
C983 B.n170 VSUBS 0.006841f
C984 B.n171 VSUBS 0.006841f
C985 B.n172 VSUBS 0.006841f
C986 B.n173 VSUBS 0.006841f
C987 B.n174 VSUBS 0.006841f
C988 B.n175 VSUBS 0.006841f
C989 B.n176 VSUBS 0.006841f
C990 B.n177 VSUBS 0.006841f
C991 B.n178 VSUBS 0.006841f
C992 B.n179 VSUBS 0.006841f
C993 B.n180 VSUBS 0.006841f
C994 B.n181 VSUBS 0.006841f
C995 B.n182 VSUBS 0.006841f
C996 B.n183 VSUBS 0.006841f
C997 B.n184 VSUBS 0.006841f
C998 B.n185 VSUBS 0.006841f
C999 B.n186 VSUBS 0.006841f
C1000 B.n187 VSUBS 0.006841f
C1001 B.n188 VSUBS 0.006841f
C1002 B.n189 VSUBS 0.006841f
C1003 B.n190 VSUBS 0.006841f
C1004 B.n191 VSUBS 0.006841f
C1005 B.n192 VSUBS 0.006841f
C1006 B.n193 VSUBS 0.006841f
C1007 B.n194 VSUBS 0.006841f
C1008 B.n195 VSUBS 0.006841f
C1009 B.n196 VSUBS 0.006841f
C1010 B.n197 VSUBS 0.006841f
C1011 B.n198 VSUBS 0.006841f
C1012 B.n199 VSUBS 0.015442f
C1013 B.n200 VSUBS 0.015442f
C1014 B.n201 VSUBS 0.016752f
C1015 B.n202 VSUBS 0.006841f
C1016 B.n203 VSUBS 0.006841f
C1017 B.n204 VSUBS 0.006841f
C1018 B.n205 VSUBS 0.006841f
C1019 B.n206 VSUBS 0.006841f
C1020 B.n207 VSUBS 0.006841f
C1021 B.n208 VSUBS 0.006841f
C1022 B.n209 VSUBS 0.006841f
C1023 B.n210 VSUBS 0.006841f
C1024 B.n211 VSUBS 0.006841f
C1025 B.n212 VSUBS 0.006841f
C1026 B.n213 VSUBS 0.006841f
C1027 B.n214 VSUBS 0.006841f
C1028 B.n215 VSUBS 0.006841f
C1029 B.n216 VSUBS 0.006841f
C1030 B.n217 VSUBS 0.006841f
C1031 B.n218 VSUBS 0.006841f
C1032 B.n219 VSUBS 0.006841f
C1033 B.n220 VSUBS 0.006841f
C1034 B.n221 VSUBS 0.006841f
C1035 B.n222 VSUBS 0.006841f
C1036 B.n223 VSUBS 0.006841f
C1037 B.n224 VSUBS 0.006841f
C1038 B.n225 VSUBS 0.006841f
C1039 B.n226 VSUBS 0.006841f
C1040 B.n227 VSUBS 0.006841f
C1041 B.n228 VSUBS 0.006841f
C1042 B.n229 VSUBS 0.006841f
C1043 B.n230 VSUBS 0.006841f
C1044 B.n231 VSUBS 0.006841f
C1045 B.n232 VSUBS 0.006841f
C1046 B.n233 VSUBS 0.006841f
C1047 B.n234 VSUBS 0.006841f
C1048 B.n235 VSUBS 0.006841f
C1049 B.n236 VSUBS 0.006841f
C1050 B.n237 VSUBS 0.006841f
C1051 B.n238 VSUBS 0.006841f
C1052 B.n239 VSUBS 0.006841f
C1053 B.n240 VSUBS 0.006841f
C1054 B.n241 VSUBS 0.006841f
C1055 B.n242 VSUBS 0.006841f
C1056 B.n243 VSUBS 0.006841f
C1057 B.n244 VSUBS 0.006841f
C1058 B.n245 VSUBS 0.006841f
C1059 B.n246 VSUBS 0.006841f
C1060 B.n247 VSUBS 0.006841f
C1061 B.n248 VSUBS 0.006841f
C1062 B.n249 VSUBS 0.006841f
C1063 B.n250 VSUBS 0.006841f
C1064 B.n251 VSUBS 0.006841f
C1065 B.n252 VSUBS 0.006841f
C1066 B.n253 VSUBS 0.006841f
C1067 B.n254 VSUBS 0.006841f
C1068 B.n255 VSUBS 0.006841f
C1069 B.n256 VSUBS 0.006841f
C1070 B.n257 VSUBS 0.006841f
C1071 B.n258 VSUBS 0.006841f
C1072 B.n259 VSUBS 0.006841f
C1073 B.n260 VSUBS 0.006841f
C1074 B.n261 VSUBS 0.006841f
C1075 B.n262 VSUBS 0.006841f
C1076 B.n263 VSUBS 0.006841f
C1077 B.n264 VSUBS 0.006841f
C1078 B.n265 VSUBS 0.006841f
C1079 B.n266 VSUBS 0.006841f
C1080 B.n267 VSUBS 0.006841f
C1081 B.n268 VSUBS 0.006841f
C1082 B.n269 VSUBS 0.006841f
C1083 B.n270 VSUBS 0.006841f
C1084 B.n271 VSUBS 0.006841f
C1085 B.n272 VSUBS 0.006841f
C1086 B.n273 VSUBS 0.006841f
C1087 B.n274 VSUBS 0.006841f
C1088 B.n275 VSUBS 0.006841f
C1089 B.n276 VSUBS 0.006841f
C1090 B.n277 VSUBS 0.006439f
C1091 B.n278 VSUBS 0.006841f
C1092 B.n279 VSUBS 0.006841f
C1093 B.n280 VSUBS 0.003823f
C1094 B.n281 VSUBS 0.006841f
C1095 B.n282 VSUBS 0.006841f
C1096 B.n283 VSUBS 0.006841f
C1097 B.n284 VSUBS 0.006841f
C1098 B.n285 VSUBS 0.006841f
C1099 B.n286 VSUBS 0.006841f
C1100 B.n287 VSUBS 0.006841f
C1101 B.n288 VSUBS 0.006841f
C1102 B.n289 VSUBS 0.006841f
C1103 B.n290 VSUBS 0.006841f
C1104 B.n291 VSUBS 0.006841f
C1105 B.n292 VSUBS 0.006841f
C1106 B.n293 VSUBS 0.003823f
C1107 B.n294 VSUBS 0.015851f
C1108 B.n295 VSUBS 0.006439f
C1109 B.n296 VSUBS 0.006841f
C1110 B.n297 VSUBS 0.006841f
C1111 B.n298 VSUBS 0.006841f
C1112 B.n299 VSUBS 0.006841f
C1113 B.n300 VSUBS 0.006841f
C1114 B.n301 VSUBS 0.006841f
C1115 B.n302 VSUBS 0.006841f
C1116 B.n303 VSUBS 0.006841f
C1117 B.n304 VSUBS 0.006841f
C1118 B.n305 VSUBS 0.006841f
C1119 B.n306 VSUBS 0.006841f
C1120 B.n307 VSUBS 0.006841f
C1121 B.n308 VSUBS 0.006841f
C1122 B.n309 VSUBS 0.006841f
C1123 B.n310 VSUBS 0.006841f
C1124 B.n311 VSUBS 0.006841f
C1125 B.n312 VSUBS 0.006841f
C1126 B.n313 VSUBS 0.006841f
C1127 B.n314 VSUBS 0.006841f
C1128 B.n315 VSUBS 0.006841f
C1129 B.n316 VSUBS 0.006841f
C1130 B.n317 VSUBS 0.006841f
C1131 B.n318 VSUBS 0.006841f
C1132 B.n319 VSUBS 0.006841f
C1133 B.n320 VSUBS 0.006841f
C1134 B.n321 VSUBS 0.006841f
C1135 B.n322 VSUBS 0.006841f
C1136 B.n323 VSUBS 0.006841f
C1137 B.n324 VSUBS 0.006841f
C1138 B.n325 VSUBS 0.006841f
C1139 B.n326 VSUBS 0.006841f
C1140 B.n327 VSUBS 0.006841f
C1141 B.n328 VSUBS 0.006841f
C1142 B.n329 VSUBS 0.006841f
C1143 B.n330 VSUBS 0.006841f
C1144 B.n331 VSUBS 0.006841f
C1145 B.n332 VSUBS 0.006841f
C1146 B.n333 VSUBS 0.006841f
C1147 B.n334 VSUBS 0.006841f
C1148 B.n335 VSUBS 0.006841f
C1149 B.n336 VSUBS 0.006841f
C1150 B.n337 VSUBS 0.006841f
C1151 B.n338 VSUBS 0.006841f
C1152 B.n339 VSUBS 0.006841f
C1153 B.n340 VSUBS 0.006841f
C1154 B.n341 VSUBS 0.006841f
C1155 B.n342 VSUBS 0.006841f
C1156 B.n343 VSUBS 0.006841f
C1157 B.n344 VSUBS 0.006841f
C1158 B.n345 VSUBS 0.006841f
C1159 B.n346 VSUBS 0.006841f
C1160 B.n347 VSUBS 0.006841f
C1161 B.n348 VSUBS 0.006841f
C1162 B.n349 VSUBS 0.006841f
C1163 B.n350 VSUBS 0.006841f
C1164 B.n351 VSUBS 0.006841f
C1165 B.n352 VSUBS 0.006841f
C1166 B.n353 VSUBS 0.006841f
C1167 B.n354 VSUBS 0.006841f
C1168 B.n355 VSUBS 0.006841f
C1169 B.n356 VSUBS 0.006841f
C1170 B.n357 VSUBS 0.006841f
C1171 B.n358 VSUBS 0.006841f
C1172 B.n359 VSUBS 0.006841f
C1173 B.n360 VSUBS 0.006841f
C1174 B.n361 VSUBS 0.006841f
C1175 B.n362 VSUBS 0.006841f
C1176 B.n363 VSUBS 0.006841f
C1177 B.n364 VSUBS 0.006841f
C1178 B.n365 VSUBS 0.006841f
C1179 B.n366 VSUBS 0.006841f
C1180 B.n367 VSUBS 0.006841f
C1181 B.n368 VSUBS 0.006841f
C1182 B.n369 VSUBS 0.006841f
C1183 B.n370 VSUBS 0.006841f
C1184 B.n371 VSUBS 0.006841f
C1185 B.n372 VSUBS 0.016752f
C1186 B.n373 VSUBS 0.015442f
C1187 B.n374 VSUBS 0.015442f
C1188 B.n375 VSUBS 0.006841f
C1189 B.n376 VSUBS 0.006841f
C1190 B.n377 VSUBS 0.006841f
C1191 B.n378 VSUBS 0.006841f
C1192 B.n379 VSUBS 0.006841f
C1193 B.n380 VSUBS 0.006841f
C1194 B.n381 VSUBS 0.006841f
C1195 B.n382 VSUBS 0.006841f
C1196 B.n383 VSUBS 0.006841f
C1197 B.n384 VSUBS 0.006841f
C1198 B.n385 VSUBS 0.006841f
C1199 B.n386 VSUBS 0.006841f
C1200 B.n387 VSUBS 0.006841f
C1201 B.n388 VSUBS 0.006841f
C1202 B.n389 VSUBS 0.006841f
C1203 B.n390 VSUBS 0.006841f
C1204 B.n391 VSUBS 0.006841f
C1205 B.n392 VSUBS 0.006841f
C1206 B.n393 VSUBS 0.006841f
C1207 B.n394 VSUBS 0.006841f
C1208 B.n395 VSUBS 0.006841f
C1209 B.n396 VSUBS 0.006841f
C1210 B.n397 VSUBS 0.006841f
C1211 B.n398 VSUBS 0.006841f
C1212 B.n399 VSUBS 0.006841f
C1213 B.n400 VSUBS 0.006841f
C1214 B.n401 VSUBS 0.006841f
C1215 B.n402 VSUBS 0.006841f
C1216 B.n403 VSUBS 0.006841f
C1217 B.n404 VSUBS 0.006841f
C1218 B.n405 VSUBS 0.006841f
C1219 B.n406 VSUBS 0.006841f
C1220 B.n407 VSUBS 0.006841f
C1221 B.n408 VSUBS 0.006841f
C1222 B.n409 VSUBS 0.006841f
C1223 B.n410 VSUBS 0.006841f
C1224 B.n411 VSUBS 0.006841f
C1225 B.n412 VSUBS 0.006841f
C1226 B.n413 VSUBS 0.006841f
C1227 B.n414 VSUBS 0.006841f
C1228 B.n415 VSUBS 0.006841f
C1229 B.n416 VSUBS 0.006841f
C1230 B.n417 VSUBS 0.006841f
C1231 B.n418 VSUBS 0.006841f
C1232 B.n419 VSUBS 0.006841f
C1233 B.n420 VSUBS 0.006841f
C1234 B.n421 VSUBS 0.006841f
C1235 B.n422 VSUBS 0.006841f
C1236 B.n423 VSUBS 0.006841f
C1237 B.n424 VSUBS 0.006841f
C1238 B.n425 VSUBS 0.006841f
C1239 B.n426 VSUBS 0.006841f
C1240 B.n427 VSUBS 0.006841f
C1241 B.n428 VSUBS 0.006841f
C1242 B.n429 VSUBS 0.006841f
C1243 B.n430 VSUBS 0.006841f
C1244 B.n431 VSUBS 0.006841f
C1245 B.n432 VSUBS 0.006841f
C1246 B.n433 VSUBS 0.006841f
C1247 B.n434 VSUBS 0.006841f
C1248 B.n435 VSUBS 0.006841f
C1249 B.n436 VSUBS 0.006841f
C1250 B.n437 VSUBS 0.006841f
C1251 B.n438 VSUBS 0.006841f
C1252 B.n439 VSUBS 0.016244f
C1253 B.n440 VSUBS 0.015442f
C1254 B.n441 VSUBS 0.016752f
C1255 B.n442 VSUBS 0.006841f
C1256 B.n443 VSUBS 0.006841f
C1257 B.n444 VSUBS 0.006841f
C1258 B.n445 VSUBS 0.006841f
C1259 B.n446 VSUBS 0.006841f
C1260 B.n447 VSUBS 0.006841f
C1261 B.n448 VSUBS 0.006841f
C1262 B.n449 VSUBS 0.006841f
C1263 B.n450 VSUBS 0.006841f
C1264 B.n451 VSUBS 0.006841f
C1265 B.n452 VSUBS 0.006841f
C1266 B.n453 VSUBS 0.006841f
C1267 B.n454 VSUBS 0.006841f
C1268 B.n455 VSUBS 0.006841f
C1269 B.n456 VSUBS 0.006841f
C1270 B.n457 VSUBS 0.006841f
C1271 B.n458 VSUBS 0.006841f
C1272 B.n459 VSUBS 0.006841f
C1273 B.n460 VSUBS 0.006841f
C1274 B.n461 VSUBS 0.006841f
C1275 B.n462 VSUBS 0.006841f
C1276 B.n463 VSUBS 0.006841f
C1277 B.n464 VSUBS 0.006841f
C1278 B.n465 VSUBS 0.006841f
C1279 B.n466 VSUBS 0.006841f
C1280 B.n467 VSUBS 0.006841f
C1281 B.n468 VSUBS 0.006841f
C1282 B.n469 VSUBS 0.006841f
C1283 B.n470 VSUBS 0.006841f
C1284 B.n471 VSUBS 0.006841f
C1285 B.n472 VSUBS 0.006841f
C1286 B.n473 VSUBS 0.006841f
C1287 B.n474 VSUBS 0.006841f
C1288 B.n475 VSUBS 0.006841f
C1289 B.n476 VSUBS 0.006841f
C1290 B.n477 VSUBS 0.006841f
C1291 B.n478 VSUBS 0.006841f
C1292 B.n479 VSUBS 0.006841f
C1293 B.n480 VSUBS 0.006841f
C1294 B.n481 VSUBS 0.006841f
C1295 B.n482 VSUBS 0.006841f
C1296 B.n483 VSUBS 0.006841f
C1297 B.n484 VSUBS 0.006841f
C1298 B.n485 VSUBS 0.006841f
C1299 B.n486 VSUBS 0.006841f
C1300 B.n487 VSUBS 0.006841f
C1301 B.n488 VSUBS 0.006841f
C1302 B.n489 VSUBS 0.006841f
C1303 B.n490 VSUBS 0.006841f
C1304 B.n491 VSUBS 0.006841f
C1305 B.n492 VSUBS 0.006841f
C1306 B.n493 VSUBS 0.006841f
C1307 B.n494 VSUBS 0.006841f
C1308 B.n495 VSUBS 0.006841f
C1309 B.n496 VSUBS 0.006841f
C1310 B.n497 VSUBS 0.006841f
C1311 B.n498 VSUBS 0.006841f
C1312 B.n499 VSUBS 0.006841f
C1313 B.n500 VSUBS 0.006841f
C1314 B.n501 VSUBS 0.006841f
C1315 B.n502 VSUBS 0.006841f
C1316 B.n503 VSUBS 0.006841f
C1317 B.n504 VSUBS 0.006841f
C1318 B.n505 VSUBS 0.006841f
C1319 B.n506 VSUBS 0.006841f
C1320 B.n507 VSUBS 0.006841f
C1321 B.n508 VSUBS 0.006841f
C1322 B.n509 VSUBS 0.006841f
C1323 B.n510 VSUBS 0.006841f
C1324 B.n511 VSUBS 0.006841f
C1325 B.n512 VSUBS 0.006841f
C1326 B.n513 VSUBS 0.006841f
C1327 B.n514 VSUBS 0.006841f
C1328 B.n515 VSUBS 0.006841f
C1329 B.n516 VSUBS 0.006841f
C1330 B.n517 VSUBS 0.006439f
C1331 B.n518 VSUBS 0.006841f
C1332 B.n519 VSUBS 0.006841f
C1333 B.n520 VSUBS 0.003823f
C1334 B.n521 VSUBS 0.006841f
C1335 B.n522 VSUBS 0.006841f
C1336 B.n523 VSUBS 0.006841f
C1337 B.n524 VSUBS 0.006841f
C1338 B.n525 VSUBS 0.006841f
C1339 B.n526 VSUBS 0.006841f
C1340 B.n527 VSUBS 0.006841f
C1341 B.n528 VSUBS 0.006841f
C1342 B.n529 VSUBS 0.006841f
C1343 B.n530 VSUBS 0.006841f
C1344 B.n531 VSUBS 0.006841f
C1345 B.n532 VSUBS 0.006841f
C1346 B.n533 VSUBS 0.003823f
C1347 B.n534 VSUBS 0.015851f
C1348 B.n535 VSUBS 0.006439f
C1349 B.n536 VSUBS 0.006841f
C1350 B.n537 VSUBS 0.006841f
C1351 B.n538 VSUBS 0.006841f
C1352 B.n539 VSUBS 0.006841f
C1353 B.n540 VSUBS 0.006841f
C1354 B.n541 VSUBS 0.006841f
C1355 B.n542 VSUBS 0.006841f
C1356 B.n543 VSUBS 0.006841f
C1357 B.n544 VSUBS 0.006841f
C1358 B.n545 VSUBS 0.006841f
C1359 B.n546 VSUBS 0.006841f
C1360 B.n547 VSUBS 0.006841f
C1361 B.n548 VSUBS 0.006841f
C1362 B.n549 VSUBS 0.006841f
C1363 B.n550 VSUBS 0.006841f
C1364 B.n551 VSUBS 0.006841f
C1365 B.n552 VSUBS 0.006841f
C1366 B.n553 VSUBS 0.006841f
C1367 B.n554 VSUBS 0.006841f
C1368 B.n555 VSUBS 0.006841f
C1369 B.n556 VSUBS 0.006841f
C1370 B.n557 VSUBS 0.006841f
C1371 B.n558 VSUBS 0.006841f
C1372 B.n559 VSUBS 0.006841f
C1373 B.n560 VSUBS 0.006841f
C1374 B.n561 VSUBS 0.006841f
C1375 B.n562 VSUBS 0.006841f
C1376 B.n563 VSUBS 0.006841f
C1377 B.n564 VSUBS 0.006841f
C1378 B.n565 VSUBS 0.006841f
C1379 B.n566 VSUBS 0.006841f
C1380 B.n567 VSUBS 0.006841f
C1381 B.n568 VSUBS 0.006841f
C1382 B.n569 VSUBS 0.006841f
C1383 B.n570 VSUBS 0.006841f
C1384 B.n571 VSUBS 0.006841f
C1385 B.n572 VSUBS 0.006841f
C1386 B.n573 VSUBS 0.006841f
C1387 B.n574 VSUBS 0.006841f
C1388 B.n575 VSUBS 0.006841f
C1389 B.n576 VSUBS 0.006841f
C1390 B.n577 VSUBS 0.006841f
C1391 B.n578 VSUBS 0.006841f
C1392 B.n579 VSUBS 0.006841f
C1393 B.n580 VSUBS 0.006841f
C1394 B.n581 VSUBS 0.006841f
C1395 B.n582 VSUBS 0.006841f
C1396 B.n583 VSUBS 0.006841f
C1397 B.n584 VSUBS 0.006841f
C1398 B.n585 VSUBS 0.006841f
C1399 B.n586 VSUBS 0.006841f
C1400 B.n587 VSUBS 0.006841f
C1401 B.n588 VSUBS 0.006841f
C1402 B.n589 VSUBS 0.006841f
C1403 B.n590 VSUBS 0.006841f
C1404 B.n591 VSUBS 0.006841f
C1405 B.n592 VSUBS 0.006841f
C1406 B.n593 VSUBS 0.006841f
C1407 B.n594 VSUBS 0.006841f
C1408 B.n595 VSUBS 0.006841f
C1409 B.n596 VSUBS 0.006841f
C1410 B.n597 VSUBS 0.006841f
C1411 B.n598 VSUBS 0.006841f
C1412 B.n599 VSUBS 0.006841f
C1413 B.n600 VSUBS 0.006841f
C1414 B.n601 VSUBS 0.006841f
C1415 B.n602 VSUBS 0.006841f
C1416 B.n603 VSUBS 0.006841f
C1417 B.n604 VSUBS 0.006841f
C1418 B.n605 VSUBS 0.006841f
C1419 B.n606 VSUBS 0.006841f
C1420 B.n607 VSUBS 0.006841f
C1421 B.n608 VSUBS 0.006841f
C1422 B.n609 VSUBS 0.006841f
C1423 B.n610 VSUBS 0.006841f
C1424 B.n611 VSUBS 0.006841f
C1425 B.n612 VSUBS 0.016752f
C1426 B.n613 VSUBS 0.015442f
C1427 B.n614 VSUBS 0.015442f
C1428 B.n615 VSUBS 0.006841f
C1429 B.n616 VSUBS 0.006841f
C1430 B.n617 VSUBS 0.006841f
C1431 B.n618 VSUBS 0.006841f
C1432 B.n619 VSUBS 0.006841f
C1433 B.n620 VSUBS 0.006841f
C1434 B.n621 VSUBS 0.006841f
C1435 B.n622 VSUBS 0.006841f
C1436 B.n623 VSUBS 0.006841f
C1437 B.n624 VSUBS 0.006841f
C1438 B.n625 VSUBS 0.006841f
C1439 B.n626 VSUBS 0.006841f
C1440 B.n627 VSUBS 0.006841f
C1441 B.n628 VSUBS 0.006841f
C1442 B.n629 VSUBS 0.006841f
C1443 B.n630 VSUBS 0.006841f
C1444 B.n631 VSUBS 0.006841f
C1445 B.n632 VSUBS 0.006841f
C1446 B.n633 VSUBS 0.006841f
C1447 B.n634 VSUBS 0.006841f
C1448 B.n635 VSUBS 0.006841f
C1449 B.n636 VSUBS 0.006841f
C1450 B.n637 VSUBS 0.006841f
C1451 B.n638 VSUBS 0.006841f
C1452 B.n639 VSUBS 0.006841f
C1453 B.n640 VSUBS 0.006841f
C1454 B.n641 VSUBS 0.006841f
C1455 B.n642 VSUBS 0.006841f
C1456 B.n643 VSUBS 0.006841f
C1457 B.n644 VSUBS 0.006841f
C1458 B.n645 VSUBS 0.006841f
C1459 B.n646 VSUBS 0.006841f
C1460 B.n647 VSUBS 0.015491f
.ends

