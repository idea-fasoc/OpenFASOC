* NGSPICE file created from diff_pair_sample_1194.ext - technology: sky130A

.subckt diff_pair_sample_1194 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X1 B.t11 B.t9 B.t10 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0 ps=0 w=1.18 l=2.8
X2 B.t8 B.t6 B.t7 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0 ps=0 w=1.18 l=2.8
X3 VTAIL.t9 VN.t1 VDD2.t6 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X4 VDD1.t7 VP.t0 VTAIL.t4 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X5 VDD2.t5 VN.t2 VTAIL.t10 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.4602 ps=3.14 w=1.18 l=2.8
X6 VTAIL.t0 VP.t1 VDD1.t6 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0.1947 ps=1.51 w=1.18 l=2.8
X7 VDD2.t4 VN.t3 VTAIL.t14 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.4602 ps=3.14 w=1.18 l=2.8
X8 VTAIL.t12 VN.t4 VDD2.t3 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0.1947 ps=1.51 w=1.18 l=2.8
X9 VDD1.t5 VP.t2 VTAIL.t1 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.4602 ps=3.14 w=1.18 l=2.8
X10 B.t5 B.t3 B.t4 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0 ps=0 w=1.18 l=2.8
X11 VDD1.t4 VP.t3 VTAIL.t7 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.4602 ps=3.14 w=1.18 l=2.8
X12 VTAIL.t6 VP.t4 VDD1.t3 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0.1947 ps=1.51 w=1.18 l=2.8
X13 VTAIL.t15 VN.t5 VDD2.t2 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X14 VDD1.t2 VP.t5 VTAIL.t3 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X15 B.t2 B.t0 B.t1 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0 ps=0 w=1.18 l=2.8
X16 VTAIL.t11 VN.t6 VDD2.t1 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.4602 pd=3.14 as=0.1947 ps=1.51 w=1.18 l=2.8
X17 VDD2.t0 VN.t7 VTAIL.t13 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X18 VTAIL.t2 VP.t6 VDD1.t1 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
X19 VTAIL.t5 VP.t7 VDD1.t0 w_n4100_n1204# sky130_fd_pr__pfet_01v8 ad=0.1947 pd=1.51 as=0.1947 ps=1.51 w=1.18 l=2.8
R0 VN.n56 VN.n55 161.3
R1 VN.n54 VN.n30 161.3
R2 VN.n53 VN.n52 161.3
R3 VN.n51 VN.n31 161.3
R4 VN.n50 VN.n49 161.3
R5 VN.n48 VN.n32 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n27 VN.n26 161.3
R13 VN.n25 VN.n1 161.3
R14 VN.n24 VN.n23 161.3
R15 VN.n22 VN.n2 161.3
R16 VN.n21 VN.n20 161.3
R17 VN.n19 VN.n3 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n28 VN.n0 68.3588
R25 VN.n57 VN.n29 68.3588
R26 VN.n8 VN.n7 58.3801
R27 VN.n37 VN.n36 58.3801
R28 VN.n13 VN.n12 56.5617
R29 VN.n42 VN.n41 56.5617
R30 VN.n24 VN.n2 52.2023
R31 VN.n53 VN.n31 52.2023
R32 VN VN.n57 43.8996
R33 VN.n37 VN.t3 42.1188
R34 VN.n8 VN.t4 42.1188
R35 VN.n25 VN.n24 28.9518
R36 VN.n54 VN.n53 28.9518
R37 VN.n11 VN.n6 24.5923
R38 VN.n12 VN.n11 24.5923
R39 VN.n13 VN.n4 24.5923
R40 VN.n17 VN.n4 24.5923
R41 VN.n20 VN.n19 24.5923
R42 VN.n20 VN.n2 24.5923
R43 VN.n26 VN.n25 24.5923
R44 VN.n41 VN.n40 24.5923
R45 VN.n40 VN.n35 24.5923
R46 VN.n49 VN.n31 24.5923
R47 VN.n49 VN.n48 24.5923
R48 VN.n46 VN.n33 24.5923
R49 VN.n42 VN.n33 24.5923
R50 VN.n55 VN.n54 24.5923
R51 VN.n26 VN.n0 21.8872
R52 VN.n55 VN.n29 21.8872
R53 VN.n7 VN.n6 15.4934
R54 VN.n18 VN.n17 15.4934
R55 VN.n36 VN.n35 15.4934
R56 VN.n47 VN.n46 15.4934
R57 VN.n7 VN.t7 10.1569
R58 VN.n18 VN.t5 10.1569
R59 VN.n0 VN.t2 10.1569
R60 VN.n36 VN.t1 10.1569
R61 VN.n47 VN.t0 10.1569
R62 VN.n29 VN.t6 10.1569
R63 VN.n19 VN.n18 9.09948
R64 VN.n48 VN.n47 9.09948
R65 VN.n38 VN.n37 5.39044
R66 VN.n9 VN.n8 5.39044
R67 VN.n57 VN.n56 0.354861
R68 VN.n28 VN.n27 0.354861
R69 VN VN.n28 0.267071
R70 VN.n56 VN.n30 0.189894
R71 VN.n52 VN.n30 0.189894
R72 VN.n52 VN.n51 0.189894
R73 VN.n51 VN.n50 0.189894
R74 VN.n50 VN.n32 0.189894
R75 VN.n45 VN.n32 0.189894
R76 VN.n45 VN.n44 0.189894
R77 VN.n44 VN.n43 0.189894
R78 VN.n43 VN.n34 0.189894
R79 VN.n39 VN.n34 0.189894
R80 VN.n39 VN.n38 0.189894
R81 VN.n10 VN.n9 0.189894
R82 VN.n10 VN.n5 0.189894
R83 VN.n14 VN.n5 0.189894
R84 VN.n15 VN.n14 0.189894
R85 VN.n16 VN.n15 0.189894
R86 VN.n16 VN.n3 0.189894
R87 VN.n21 VN.n3 0.189894
R88 VN.n22 VN.n21 0.189894
R89 VN.n23 VN.n22 0.189894
R90 VN.n23 VN.n1 0.189894
R91 VN.n27 VN.n1 0.189894
R92 VTAIL.n15 VTAIL.t10 374.075
R93 VTAIL.n2 VTAIL.t12 374.075
R94 VTAIL.n3 VTAIL.t7 374.075
R95 VTAIL.n6 VTAIL.t0 374.075
R96 VTAIL.n14 VTAIL.t1 374.075
R97 VTAIL.n11 VTAIL.t6 374.075
R98 VTAIL.n10 VTAIL.t14 374.075
R99 VTAIL.n7 VTAIL.t11 374.075
R100 VTAIL.n1 VTAIL.n0 331.137
R101 VTAIL.n5 VTAIL.n4 331.137
R102 VTAIL.n13 VTAIL.n12 331.135
R103 VTAIL.n9 VTAIL.n8 331.135
R104 VTAIL.n0 VTAIL.t13 27.5471
R105 VTAIL.n0 VTAIL.t15 27.5471
R106 VTAIL.n4 VTAIL.t3 27.5471
R107 VTAIL.n4 VTAIL.t2 27.5471
R108 VTAIL.n12 VTAIL.t4 27.5471
R109 VTAIL.n12 VTAIL.t5 27.5471
R110 VTAIL.n8 VTAIL.t8 27.5471
R111 VTAIL.n8 VTAIL.t9 27.5471
R112 VTAIL.n15 VTAIL.n14 16.0824
R113 VTAIL.n7 VTAIL.n6 16.0824
R114 VTAIL.n9 VTAIL.n7 2.69878
R115 VTAIL.n10 VTAIL.n9 2.69878
R116 VTAIL.n13 VTAIL.n11 2.69878
R117 VTAIL.n14 VTAIL.n13 2.69878
R118 VTAIL.n6 VTAIL.n5 2.69878
R119 VTAIL.n5 VTAIL.n3 2.69878
R120 VTAIL.n2 VTAIL.n1 2.69878
R121 VTAIL VTAIL.n15 2.64059
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 349.11
R126 VDD2.n2 VDD2.n0 349.11
R127 VDD2 VDD2.n5 349.106
R128 VDD2.n4 VDD2.n3 347.815
R129 VDD2.n4 VDD2.n2 36.8748
R130 VDD2.n5 VDD2.t6 27.5471
R131 VDD2.n5 VDD2.t4 27.5471
R132 VDD2.n3 VDD2.t1 27.5471
R133 VDD2.n3 VDD2.t7 27.5471
R134 VDD2.n1 VDD2.t2 27.5471
R135 VDD2.n1 VDD2.t5 27.5471
R136 VDD2.n0 VDD2.t3 27.5471
R137 VDD2.n0 VDD2.t0 27.5471
R138 VDD2 VDD2.n4 1.40783
R139 B.n437 B.n436 585
R140 B.n438 B.n47 585
R141 B.n440 B.n439 585
R142 B.n441 B.n46 585
R143 B.n443 B.n442 585
R144 B.n444 B.n45 585
R145 B.n446 B.n445 585
R146 B.n447 B.n44 585
R147 B.n449 B.n448 585
R148 B.n450 B.n41 585
R149 B.n453 B.n452 585
R150 B.n454 B.n40 585
R151 B.n456 B.n455 585
R152 B.n457 B.n39 585
R153 B.n459 B.n458 585
R154 B.n460 B.n38 585
R155 B.n462 B.n461 585
R156 B.n463 B.n37 585
R157 B.n465 B.n464 585
R158 B.n467 B.n466 585
R159 B.n468 B.n33 585
R160 B.n470 B.n469 585
R161 B.n471 B.n32 585
R162 B.n473 B.n472 585
R163 B.n474 B.n31 585
R164 B.n476 B.n475 585
R165 B.n477 B.n30 585
R166 B.n479 B.n478 585
R167 B.n480 B.n29 585
R168 B.n435 B.n48 585
R169 B.n434 B.n433 585
R170 B.n432 B.n49 585
R171 B.n431 B.n430 585
R172 B.n429 B.n50 585
R173 B.n428 B.n427 585
R174 B.n426 B.n51 585
R175 B.n425 B.n424 585
R176 B.n423 B.n52 585
R177 B.n422 B.n421 585
R178 B.n420 B.n53 585
R179 B.n419 B.n418 585
R180 B.n417 B.n54 585
R181 B.n416 B.n415 585
R182 B.n414 B.n55 585
R183 B.n413 B.n412 585
R184 B.n411 B.n56 585
R185 B.n410 B.n409 585
R186 B.n408 B.n57 585
R187 B.n407 B.n406 585
R188 B.n405 B.n58 585
R189 B.n404 B.n403 585
R190 B.n402 B.n59 585
R191 B.n401 B.n400 585
R192 B.n399 B.n60 585
R193 B.n398 B.n397 585
R194 B.n396 B.n61 585
R195 B.n395 B.n394 585
R196 B.n393 B.n62 585
R197 B.n392 B.n391 585
R198 B.n390 B.n63 585
R199 B.n389 B.n388 585
R200 B.n387 B.n64 585
R201 B.n386 B.n385 585
R202 B.n384 B.n65 585
R203 B.n383 B.n382 585
R204 B.n381 B.n66 585
R205 B.n380 B.n379 585
R206 B.n378 B.n67 585
R207 B.n377 B.n376 585
R208 B.n375 B.n68 585
R209 B.n374 B.n373 585
R210 B.n372 B.n69 585
R211 B.n371 B.n370 585
R212 B.n369 B.n70 585
R213 B.n368 B.n367 585
R214 B.n366 B.n71 585
R215 B.n365 B.n364 585
R216 B.n363 B.n72 585
R217 B.n362 B.n361 585
R218 B.n360 B.n73 585
R219 B.n359 B.n358 585
R220 B.n357 B.n74 585
R221 B.n356 B.n355 585
R222 B.n354 B.n75 585
R223 B.n353 B.n352 585
R224 B.n351 B.n76 585
R225 B.n350 B.n349 585
R226 B.n348 B.n77 585
R227 B.n347 B.n346 585
R228 B.n345 B.n78 585
R229 B.n344 B.n343 585
R230 B.n342 B.n79 585
R231 B.n341 B.n340 585
R232 B.n339 B.n80 585
R233 B.n338 B.n337 585
R234 B.n336 B.n81 585
R235 B.n335 B.n334 585
R236 B.n333 B.n82 585
R237 B.n332 B.n331 585
R238 B.n330 B.n83 585
R239 B.n329 B.n328 585
R240 B.n327 B.n84 585
R241 B.n326 B.n325 585
R242 B.n324 B.n85 585
R243 B.n323 B.n322 585
R244 B.n321 B.n86 585
R245 B.n320 B.n319 585
R246 B.n318 B.n87 585
R247 B.n317 B.n316 585
R248 B.n315 B.n88 585
R249 B.n314 B.n313 585
R250 B.n312 B.n89 585
R251 B.n311 B.n310 585
R252 B.n309 B.n90 585
R253 B.n308 B.n307 585
R254 B.n306 B.n91 585
R255 B.n305 B.n304 585
R256 B.n303 B.n92 585
R257 B.n302 B.n301 585
R258 B.n300 B.n93 585
R259 B.n299 B.n298 585
R260 B.n297 B.n94 585
R261 B.n296 B.n295 585
R262 B.n294 B.n95 585
R263 B.n293 B.n292 585
R264 B.n291 B.n96 585
R265 B.n290 B.n289 585
R266 B.n288 B.n97 585
R267 B.n287 B.n286 585
R268 B.n285 B.n98 585
R269 B.n284 B.n283 585
R270 B.n282 B.n99 585
R271 B.n281 B.n280 585
R272 B.n279 B.n100 585
R273 B.n278 B.n277 585
R274 B.n276 B.n101 585
R275 B.n275 B.n274 585
R276 B.n273 B.n102 585
R277 B.n228 B.n121 585
R278 B.n230 B.n229 585
R279 B.n231 B.n120 585
R280 B.n233 B.n232 585
R281 B.n234 B.n119 585
R282 B.n236 B.n235 585
R283 B.n237 B.n118 585
R284 B.n239 B.n238 585
R285 B.n240 B.n117 585
R286 B.n242 B.n241 585
R287 B.n244 B.n243 585
R288 B.n245 B.n113 585
R289 B.n247 B.n246 585
R290 B.n248 B.n112 585
R291 B.n250 B.n249 585
R292 B.n251 B.n111 585
R293 B.n253 B.n252 585
R294 B.n254 B.n110 585
R295 B.n256 B.n255 585
R296 B.n258 B.n107 585
R297 B.n260 B.n259 585
R298 B.n261 B.n106 585
R299 B.n263 B.n262 585
R300 B.n264 B.n105 585
R301 B.n266 B.n265 585
R302 B.n267 B.n104 585
R303 B.n269 B.n268 585
R304 B.n270 B.n103 585
R305 B.n272 B.n271 585
R306 B.n227 B.n226 585
R307 B.n225 B.n122 585
R308 B.n224 B.n223 585
R309 B.n222 B.n123 585
R310 B.n221 B.n220 585
R311 B.n219 B.n124 585
R312 B.n218 B.n217 585
R313 B.n216 B.n125 585
R314 B.n215 B.n214 585
R315 B.n213 B.n126 585
R316 B.n212 B.n211 585
R317 B.n210 B.n127 585
R318 B.n209 B.n208 585
R319 B.n207 B.n128 585
R320 B.n206 B.n205 585
R321 B.n204 B.n129 585
R322 B.n203 B.n202 585
R323 B.n201 B.n130 585
R324 B.n200 B.n199 585
R325 B.n198 B.n131 585
R326 B.n197 B.n196 585
R327 B.n195 B.n132 585
R328 B.n194 B.n193 585
R329 B.n192 B.n133 585
R330 B.n191 B.n190 585
R331 B.n189 B.n134 585
R332 B.n188 B.n187 585
R333 B.n186 B.n135 585
R334 B.n185 B.n184 585
R335 B.n183 B.n136 585
R336 B.n182 B.n181 585
R337 B.n180 B.n137 585
R338 B.n179 B.n178 585
R339 B.n177 B.n138 585
R340 B.n176 B.n175 585
R341 B.n174 B.n139 585
R342 B.n173 B.n172 585
R343 B.n171 B.n140 585
R344 B.n170 B.n169 585
R345 B.n168 B.n141 585
R346 B.n167 B.n166 585
R347 B.n165 B.n142 585
R348 B.n164 B.n163 585
R349 B.n162 B.n143 585
R350 B.n161 B.n160 585
R351 B.n159 B.n144 585
R352 B.n158 B.n157 585
R353 B.n156 B.n145 585
R354 B.n155 B.n154 585
R355 B.n153 B.n146 585
R356 B.n152 B.n151 585
R357 B.n150 B.n147 585
R358 B.n149 B.n148 585
R359 B.n2 B.n0 585
R360 B.n561 B.n1 585
R361 B.n560 B.n559 585
R362 B.n558 B.n3 585
R363 B.n557 B.n556 585
R364 B.n555 B.n4 585
R365 B.n554 B.n553 585
R366 B.n552 B.n5 585
R367 B.n551 B.n550 585
R368 B.n549 B.n6 585
R369 B.n548 B.n547 585
R370 B.n546 B.n7 585
R371 B.n545 B.n544 585
R372 B.n543 B.n8 585
R373 B.n542 B.n541 585
R374 B.n540 B.n9 585
R375 B.n539 B.n538 585
R376 B.n537 B.n10 585
R377 B.n536 B.n535 585
R378 B.n534 B.n11 585
R379 B.n533 B.n532 585
R380 B.n531 B.n12 585
R381 B.n530 B.n529 585
R382 B.n528 B.n13 585
R383 B.n527 B.n526 585
R384 B.n525 B.n14 585
R385 B.n524 B.n523 585
R386 B.n522 B.n15 585
R387 B.n521 B.n520 585
R388 B.n519 B.n16 585
R389 B.n518 B.n517 585
R390 B.n516 B.n17 585
R391 B.n515 B.n514 585
R392 B.n513 B.n18 585
R393 B.n512 B.n511 585
R394 B.n510 B.n19 585
R395 B.n509 B.n508 585
R396 B.n507 B.n20 585
R397 B.n506 B.n505 585
R398 B.n504 B.n21 585
R399 B.n503 B.n502 585
R400 B.n501 B.n22 585
R401 B.n500 B.n499 585
R402 B.n498 B.n23 585
R403 B.n497 B.n496 585
R404 B.n495 B.n24 585
R405 B.n494 B.n493 585
R406 B.n492 B.n25 585
R407 B.n491 B.n490 585
R408 B.n489 B.n26 585
R409 B.n488 B.n487 585
R410 B.n486 B.n27 585
R411 B.n485 B.n484 585
R412 B.n483 B.n28 585
R413 B.n482 B.n481 585
R414 B.n563 B.n562 585
R415 B.n226 B.n121 535.745
R416 B.n482 B.n29 535.745
R417 B.n273 B.n272 535.745
R418 B.n436 B.n435 535.745
R419 B.n108 B.t8 425.394
R420 B.n114 B.t11 425.394
R421 B.n34 B.t1 425.394
R422 B.n42 B.t4 425.394
R423 B.n109 B.t7 364.69
R424 B.n115 B.t10 364.69
R425 B.n35 B.t2 364.69
R426 B.n43 B.t5 364.69
R427 B.n108 B.t6 209.06
R428 B.n114 B.t9 209.06
R429 B.n34 B.t0 209.06
R430 B.n42 B.t3 209.06
R431 B.n226 B.n225 163.367
R432 B.n225 B.n224 163.367
R433 B.n224 B.n123 163.367
R434 B.n220 B.n123 163.367
R435 B.n220 B.n219 163.367
R436 B.n219 B.n218 163.367
R437 B.n218 B.n125 163.367
R438 B.n214 B.n125 163.367
R439 B.n214 B.n213 163.367
R440 B.n213 B.n212 163.367
R441 B.n212 B.n127 163.367
R442 B.n208 B.n127 163.367
R443 B.n208 B.n207 163.367
R444 B.n207 B.n206 163.367
R445 B.n206 B.n129 163.367
R446 B.n202 B.n129 163.367
R447 B.n202 B.n201 163.367
R448 B.n201 B.n200 163.367
R449 B.n200 B.n131 163.367
R450 B.n196 B.n131 163.367
R451 B.n196 B.n195 163.367
R452 B.n195 B.n194 163.367
R453 B.n194 B.n133 163.367
R454 B.n190 B.n133 163.367
R455 B.n190 B.n189 163.367
R456 B.n189 B.n188 163.367
R457 B.n188 B.n135 163.367
R458 B.n184 B.n135 163.367
R459 B.n184 B.n183 163.367
R460 B.n183 B.n182 163.367
R461 B.n182 B.n137 163.367
R462 B.n178 B.n137 163.367
R463 B.n178 B.n177 163.367
R464 B.n177 B.n176 163.367
R465 B.n176 B.n139 163.367
R466 B.n172 B.n139 163.367
R467 B.n172 B.n171 163.367
R468 B.n171 B.n170 163.367
R469 B.n170 B.n141 163.367
R470 B.n166 B.n141 163.367
R471 B.n166 B.n165 163.367
R472 B.n165 B.n164 163.367
R473 B.n164 B.n143 163.367
R474 B.n160 B.n143 163.367
R475 B.n160 B.n159 163.367
R476 B.n159 B.n158 163.367
R477 B.n158 B.n145 163.367
R478 B.n154 B.n145 163.367
R479 B.n154 B.n153 163.367
R480 B.n153 B.n152 163.367
R481 B.n152 B.n147 163.367
R482 B.n148 B.n147 163.367
R483 B.n148 B.n2 163.367
R484 B.n562 B.n2 163.367
R485 B.n562 B.n561 163.367
R486 B.n561 B.n560 163.367
R487 B.n560 B.n3 163.367
R488 B.n556 B.n3 163.367
R489 B.n556 B.n555 163.367
R490 B.n555 B.n554 163.367
R491 B.n554 B.n5 163.367
R492 B.n550 B.n5 163.367
R493 B.n550 B.n549 163.367
R494 B.n549 B.n548 163.367
R495 B.n548 B.n7 163.367
R496 B.n544 B.n7 163.367
R497 B.n544 B.n543 163.367
R498 B.n543 B.n542 163.367
R499 B.n542 B.n9 163.367
R500 B.n538 B.n9 163.367
R501 B.n538 B.n537 163.367
R502 B.n537 B.n536 163.367
R503 B.n536 B.n11 163.367
R504 B.n532 B.n11 163.367
R505 B.n532 B.n531 163.367
R506 B.n531 B.n530 163.367
R507 B.n530 B.n13 163.367
R508 B.n526 B.n13 163.367
R509 B.n526 B.n525 163.367
R510 B.n525 B.n524 163.367
R511 B.n524 B.n15 163.367
R512 B.n520 B.n15 163.367
R513 B.n520 B.n519 163.367
R514 B.n519 B.n518 163.367
R515 B.n518 B.n17 163.367
R516 B.n514 B.n17 163.367
R517 B.n514 B.n513 163.367
R518 B.n513 B.n512 163.367
R519 B.n512 B.n19 163.367
R520 B.n508 B.n19 163.367
R521 B.n508 B.n507 163.367
R522 B.n507 B.n506 163.367
R523 B.n506 B.n21 163.367
R524 B.n502 B.n21 163.367
R525 B.n502 B.n501 163.367
R526 B.n501 B.n500 163.367
R527 B.n500 B.n23 163.367
R528 B.n496 B.n23 163.367
R529 B.n496 B.n495 163.367
R530 B.n495 B.n494 163.367
R531 B.n494 B.n25 163.367
R532 B.n490 B.n25 163.367
R533 B.n490 B.n489 163.367
R534 B.n489 B.n488 163.367
R535 B.n488 B.n27 163.367
R536 B.n484 B.n27 163.367
R537 B.n484 B.n483 163.367
R538 B.n483 B.n482 163.367
R539 B.n230 B.n121 163.367
R540 B.n231 B.n230 163.367
R541 B.n232 B.n231 163.367
R542 B.n232 B.n119 163.367
R543 B.n236 B.n119 163.367
R544 B.n237 B.n236 163.367
R545 B.n238 B.n237 163.367
R546 B.n238 B.n117 163.367
R547 B.n242 B.n117 163.367
R548 B.n243 B.n242 163.367
R549 B.n243 B.n113 163.367
R550 B.n247 B.n113 163.367
R551 B.n248 B.n247 163.367
R552 B.n249 B.n248 163.367
R553 B.n249 B.n111 163.367
R554 B.n253 B.n111 163.367
R555 B.n254 B.n253 163.367
R556 B.n255 B.n254 163.367
R557 B.n255 B.n107 163.367
R558 B.n260 B.n107 163.367
R559 B.n261 B.n260 163.367
R560 B.n262 B.n261 163.367
R561 B.n262 B.n105 163.367
R562 B.n266 B.n105 163.367
R563 B.n267 B.n266 163.367
R564 B.n268 B.n267 163.367
R565 B.n268 B.n103 163.367
R566 B.n272 B.n103 163.367
R567 B.n274 B.n273 163.367
R568 B.n274 B.n101 163.367
R569 B.n278 B.n101 163.367
R570 B.n279 B.n278 163.367
R571 B.n280 B.n279 163.367
R572 B.n280 B.n99 163.367
R573 B.n284 B.n99 163.367
R574 B.n285 B.n284 163.367
R575 B.n286 B.n285 163.367
R576 B.n286 B.n97 163.367
R577 B.n290 B.n97 163.367
R578 B.n291 B.n290 163.367
R579 B.n292 B.n291 163.367
R580 B.n292 B.n95 163.367
R581 B.n296 B.n95 163.367
R582 B.n297 B.n296 163.367
R583 B.n298 B.n297 163.367
R584 B.n298 B.n93 163.367
R585 B.n302 B.n93 163.367
R586 B.n303 B.n302 163.367
R587 B.n304 B.n303 163.367
R588 B.n304 B.n91 163.367
R589 B.n308 B.n91 163.367
R590 B.n309 B.n308 163.367
R591 B.n310 B.n309 163.367
R592 B.n310 B.n89 163.367
R593 B.n314 B.n89 163.367
R594 B.n315 B.n314 163.367
R595 B.n316 B.n315 163.367
R596 B.n316 B.n87 163.367
R597 B.n320 B.n87 163.367
R598 B.n321 B.n320 163.367
R599 B.n322 B.n321 163.367
R600 B.n322 B.n85 163.367
R601 B.n326 B.n85 163.367
R602 B.n327 B.n326 163.367
R603 B.n328 B.n327 163.367
R604 B.n328 B.n83 163.367
R605 B.n332 B.n83 163.367
R606 B.n333 B.n332 163.367
R607 B.n334 B.n333 163.367
R608 B.n334 B.n81 163.367
R609 B.n338 B.n81 163.367
R610 B.n339 B.n338 163.367
R611 B.n340 B.n339 163.367
R612 B.n340 B.n79 163.367
R613 B.n344 B.n79 163.367
R614 B.n345 B.n344 163.367
R615 B.n346 B.n345 163.367
R616 B.n346 B.n77 163.367
R617 B.n350 B.n77 163.367
R618 B.n351 B.n350 163.367
R619 B.n352 B.n351 163.367
R620 B.n352 B.n75 163.367
R621 B.n356 B.n75 163.367
R622 B.n357 B.n356 163.367
R623 B.n358 B.n357 163.367
R624 B.n358 B.n73 163.367
R625 B.n362 B.n73 163.367
R626 B.n363 B.n362 163.367
R627 B.n364 B.n363 163.367
R628 B.n364 B.n71 163.367
R629 B.n368 B.n71 163.367
R630 B.n369 B.n368 163.367
R631 B.n370 B.n369 163.367
R632 B.n370 B.n69 163.367
R633 B.n374 B.n69 163.367
R634 B.n375 B.n374 163.367
R635 B.n376 B.n375 163.367
R636 B.n376 B.n67 163.367
R637 B.n380 B.n67 163.367
R638 B.n381 B.n380 163.367
R639 B.n382 B.n381 163.367
R640 B.n382 B.n65 163.367
R641 B.n386 B.n65 163.367
R642 B.n387 B.n386 163.367
R643 B.n388 B.n387 163.367
R644 B.n388 B.n63 163.367
R645 B.n392 B.n63 163.367
R646 B.n393 B.n392 163.367
R647 B.n394 B.n393 163.367
R648 B.n394 B.n61 163.367
R649 B.n398 B.n61 163.367
R650 B.n399 B.n398 163.367
R651 B.n400 B.n399 163.367
R652 B.n400 B.n59 163.367
R653 B.n404 B.n59 163.367
R654 B.n405 B.n404 163.367
R655 B.n406 B.n405 163.367
R656 B.n406 B.n57 163.367
R657 B.n410 B.n57 163.367
R658 B.n411 B.n410 163.367
R659 B.n412 B.n411 163.367
R660 B.n412 B.n55 163.367
R661 B.n416 B.n55 163.367
R662 B.n417 B.n416 163.367
R663 B.n418 B.n417 163.367
R664 B.n418 B.n53 163.367
R665 B.n422 B.n53 163.367
R666 B.n423 B.n422 163.367
R667 B.n424 B.n423 163.367
R668 B.n424 B.n51 163.367
R669 B.n428 B.n51 163.367
R670 B.n429 B.n428 163.367
R671 B.n430 B.n429 163.367
R672 B.n430 B.n49 163.367
R673 B.n434 B.n49 163.367
R674 B.n435 B.n434 163.367
R675 B.n478 B.n29 163.367
R676 B.n478 B.n477 163.367
R677 B.n477 B.n476 163.367
R678 B.n476 B.n31 163.367
R679 B.n472 B.n31 163.367
R680 B.n472 B.n471 163.367
R681 B.n471 B.n470 163.367
R682 B.n470 B.n33 163.367
R683 B.n466 B.n33 163.367
R684 B.n466 B.n465 163.367
R685 B.n465 B.n37 163.367
R686 B.n461 B.n37 163.367
R687 B.n461 B.n460 163.367
R688 B.n460 B.n459 163.367
R689 B.n459 B.n39 163.367
R690 B.n455 B.n39 163.367
R691 B.n455 B.n454 163.367
R692 B.n454 B.n453 163.367
R693 B.n453 B.n41 163.367
R694 B.n448 B.n41 163.367
R695 B.n448 B.n447 163.367
R696 B.n447 B.n446 163.367
R697 B.n446 B.n45 163.367
R698 B.n442 B.n45 163.367
R699 B.n442 B.n441 163.367
R700 B.n441 B.n440 163.367
R701 B.n440 B.n47 163.367
R702 B.n436 B.n47 163.367
R703 B.n109 B.n108 60.7035
R704 B.n115 B.n114 60.7035
R705 B.n35 B.n34 60.7035
R706 B.n43 B.n42 60.7035
R707 B.n257 B.n109 59.5399
R708 B.n116 B.n115 59.5399
R709 B.n36 B.n35 59.5399
R710 B.n451 B.n43 59.5399
R711 B.n481 B.n480 34.8103
R712 B.n437 B.n48 34.8103
R713 B.n271 B.n102 34.8103
R714 B.n228 B.n227 34.8103
R715 B B.n563 18.0485
R716 B.n480 B.n479 10.6151
R717 B.n479 B.n30 10.6151
R718 B.n475 B.n30 10.6151
R719 B.n475 B.n474 10.6151
R720 B.n474 B.n473 10.6151
R721 B.n473 B.n32 10.6151
R722 B.n469 B.n32 10.6151
R723 B.n469 B.n468 10.6151
R724 B.n468 B.n467 10.6151
R725 B.n464 B.n463 10.6151
R726 B.n463 B.n462 10.6151
R727 B.n462 B.n38 10.6151
R728 B.n458 B.n38 10.6151
R729 B.n458 B.n457 10.6151
R730 B.n457 B.n456 10.6151
R731 B.n456 B.n40 10.6151
R732 B.n452 B.n40 10.6151
R733 B.n450 B.n449 10.6151
R734 B.n449 B.n44 10.6151
R735 B.n445 B.n44 10.6151
R736 B.n445 B.n444 10.6151
R737 B.n444 B.n443 10.6151
R738 B.n443 B.n46 10.6151
R739 B.n439 B.n46 10.6151
R740 B.n439 B.n438 10.6151
R741 B.n438 B.n437 10.6151
R742 B.n275 B.n102 10.6151
R743 B.n276 B.n275 10.6151
R744 B.n277 B.n276 10.6151
R745 B.n277 B.n100 10.6151
R746 B.n281 B.n100 10.6151
R747 B.n282 B.n281 10.6151
R748 B.n283 B.n282 10.6151
R749 B.n283 B.n98 10.6151
R750 B.n287 B.n98 10.6151
R751 B.n288 B.n287 10.6151
R752 B.n289 B.n288 10.6151
R753 B.n289 B.n96 10.6151
R754 B.n293 B.n96 10.6151
R755 B.n294 B.n293 10.6151
R756 B.n295 B.n294 10.6151
R757 B.n295 B.n94 10.6151
R758 B.n299 B.n94 10.6151
R759 B.n300 B.n299 10.6151
R760 B.n301 B.n300 10.6151
R761 B.n301 B.n92 10.6151
R762 B.n305 B.n92 10.6151
R763 B.n306 B.n305 10.6151
R764 B.n307 B.n306 10.6151
R765 B.n307 B.n90 10.6151
R766 B.n311 B.n90 10.6151
R767 B.n312 B.n311 10.6151
R768 B.n313 B.n312 10.6151
R769 B.n313 B.n88 10.6151
R770 B.n317 B.n88 10.6151
R771 B.n318 B.n317 10.6151
R772 B.n319 B.n318 10.6151
R773 B.n319 B.n86 10.6151
R774 B.n323 B.n86 10.6151
R775 B.n324 B.n323 10.6151
R776 B.n325 B.n324 10.6151
R777 B.n325 B.n84 10.6151
R778 B.n329 B.n84 10.6151
R779 B.n330 B.n329 10.6151
R780 B.n331 B.n330 10.6151
R781 B.n331 B.n82 10.6151
R782 B.n335 B.n82 10.6151
R783 B.n336 B.n335 10.6151
R784 B.n337 B.n336 10.6151
R785 B.n337 B.n80 10.6151
R786 B.n341 B.n80 10.6151
R787 B.n342 B.n341 10.6151
R788 B.n343 B.n342 10.6151
R789 B.n343 B.n78 10.6151
R790 B.n347 B.n78 10.6151
R791 B.n348 B.n347 10.6151
R792 B.n349 B.n348 10.6151
R793 B.n349 B.n76 10.6151
R794 B.n353 B.n76 10.6151
R795 B.n354 B.n353 10.6151
R796 B.n355 B.n354 10.6151
R797 B.n355 B.n74 10.6151
R798 B.n359 B.n74 10.6151
R799 B.n360 B.n359 10.6151
R800 B.n361 B.n360 10.6151
R801 B.n361 B.n72 10.6151
R802 B.n365 B.n72 10.6151
R803 B.n366 B.n365 10.6151
R804 B.n367 B.n366 10.6151
R805 B.n367 B.n70 10.6151
R806 B.n371 B.n70 10.6151
R807 B.n372 B.n371 10.6151
R808 B.n373 B.n372 10.6151
R809 B.n373 B.n68 10.6151
R810 B.n377 B.n68 10.6151
R811 B.n378 B.n377 10.6151
R812 B.n379 B.n378 10.6151
R813 B.n379 B.n66 10.6151
R814 B.n383 B.n66 10.6151
R815 B.n384 B.n383 10.6151
R816 B.n385 B.n384 10.6151
R817 B.n385 B.n64 10.6151
R818 B.n389 B.n64 10.6151
R819 B.n390 B.n389 10.6151
R820 B.n391 B.n390 10.6151
R821 B.n391 B.n62 10.6151
R822 B.n395 B.n62 10.6151
R823 B.n396 B.n395 10.6151
R824 B.n397 B.n396 10.6151
R825 B.n397 B.n60 10.6151
R826 B.n401 B.n60 10.6151
R827 B.n402 B.n401 10.6151
R828 B.n403 B.n402 10.6151
R829 B.n403 B.n58 10.6151
R830 B.n407 B.n58 10.6151
R831 B.n408 B.n407 10.6151
R832 B.n409 B.n408 10.6151
R833 B.n409 B.n56 10.6151
R834 B.n413 B.n56 10.6151
R835 B.n414 B.n413 10.6151
R836 B.n415 B.n414 10.6151
R837 B.n415 B.n54 10.6151
R838 B.n419 B.n54 10.6151
R839 B.n420 B.n419 10.6151
R840 B.n421 B.n420 10.6151
R841 B.n421 B.n52 10.6151
R842 B.n425 B.n52 10.6151
R843 B.n426 B.n425 10.6151
R844 B.n427 B.n426 10.6151
R845 B.n427 B.n50 10.6151
R846 B.n431 B.n50 10.6151
R847 B.n432 B.n431 10.6151
R848 B.n433 B.n432 10.6151
R849 B.n433 B.n48 10.6151
R850 B.n229 B.n228 10.6151
R851 B.n229 B.n120 10.6151
R852 B.n233 B.n120 10.6151
R853 B.n234 B.n233 10.6151
R854 B.n235 B.n234 10.6151
R855 B.n235 B.n118 10.6151
R856 B.n239 B.n118 10.6151
R857 B.n240 B.n239 10.6151
R858 B.n241 B.n240 10.6151
R859 B.n245 B.n244 10.6151
R860 B.n246 B.n245 10.6151
R861 B.n246 B.n112 10.6151
R862 B.n250 B.n112 10.6151
R863 B.n251 B.n250 10.6151
R864 B.n252 B.n251 10.6151
R865 B.n252 B.n110 10.6151
R866 B.n256 B.n110 10.6151
R867 B.n259 B.n258 10.6151
R868 B.n259 B.n106 10.6151
R869 B.n263 B.n106 10.6151
R870 B.n264 B.n263 10.6151
R871 B.n265 B.n264 10.6151
R872 B.n265 B.n104 10.6151
R873 B.n269 B.n104 10.6151
R874 B.n270 B.n269 10.6151
R875 B.n271 B.n270 10.6151
R876 B.n227 B.n122 10.6151
R877 B.n223 B.n122 10.6151
R878 B.n223 B.n222 10.6151
R879 B.n222 B.n221 10.6151
R880 B.n221 B.n124 10.6151
R881 B.n217 B.n124 10.6151
R882 B.n217 B.n216 10.6151
R883 B.n216 B.n215 10.6151
R884 B.n215 B.n126 10.6151
R885 B.n211 B.n126 10.6151
R886 B.n211 B.n210 10.6151
R887 B.n210 B.n209 10.6151
R888 B.n209 B.n128 10.6151
R889 B.n205 B.n128 10.6151
R890 B.n205 B.n204 10.6151
R891 B.n204 B.n203 10.6151
R892 B.n203 B.n130 10.6151
R893 B.n199 B.n130 10.6151
R894 B.n199 B.n198 10.6151
R895 B.n198 B.n197 10.6151
R896 B.n197 B.n132 10.6151
R897 B.n193 B.n132 10.6151
R898 B.n193 B.n192 10.6151
R899 B.n192 B.n191 10.6151
R900 B.n191 B.n134 10.6151
R901 B.n187 B.n134 10.6151
R902 B.n187 B.n186 10.6151
R903 B.n186 B.n185 10.6151
R904 B.n185 B.n136 10.6151
R905 B.n181 B.n136 10.6151
R906 B.n181 B.n180 10.6151
R907 B.n180 B.n179 10.6151
R908 B.n179 B.n138 10.6151
R909 B.n175 B.n138 10.6151
R910 B.n175 B.n174 10.6151
R911 B.n174 B.n173 10.6151
R912 B.n173 B.n140 10.6151
R913 B.n169 B.n140 10.6151
R914 B.n169 B.n168 10.6151
R915 B.n168 B.n167 10.6151
R916 B.n167 B.n142 10.6151
R917 B.n163 B.n142 10.6151
R918 B.n163 B.n162 10.6151
R919 B.n162 B.n161 10.6151
R920 B.n161 B.n144 10.6151
R921 B.n157 B.n144 10.6151
R922 B.n157 B.n156 10.6151
R923 B.n156 B.n155 10.6151
R924 B.n155 B.n146 10.6151
R925 B.n151 B.n146 10.6151
R926 B.n151 B.n150 10.6151
R927 B.n150 B.n149 10.6151
R928 B.n149 B.n0 10.6151
R929 B.n559 B.n1 10.6151
R930 B.n559 B.n558 10.6151
R931 B.n558 B.n557 10.6151
R932 B.n557 B.n4 10.6151
R933 B.n553 B.n4 10.6151
R934 B.n553 B.n552 10.6151
R935 B.n552 B.n551 10.6151
R936 B.n551 B.n6 10.6151
R937 B.n547 B.n6 10.6151
R938 B.n547 B.n546 10.6151
R939 B.n546 B.n545 10.6151
R940 B.n545 B.n8 10.6151
R941 B.n541 B.n8 10.6151
R942 B.n541 B.n540 10.6151
R943 B.n540 B.n539 10.6151
R944 B.n539 B.n10 10.6151
R945 B.n535 B.n10 10.6151
R946 B.n535 B.n534 10.6151
R947 B.n534 B.n533 10.6151
R948 B.n533 B.n12 10.6151
R949 B.n529 B.n12 10.6151
R950 B.n529 B.n528 10.6151
R951 B.n528 B.n527 10.6151
R952 B.n527 B.n14 10.6151
R953 B.n523 B.n14 10.6151
R954 B.n523 B.n522 10.6151
R955 B.n522 B.n521 10.6151
R956 B.n521 B.n16 10.6151
R957 B.n517 B.n16 10.6151
R958 B.n517 B.n516 10.6151
R959 B.n516 B.n515 10.6151
R960 B.n515 B.n18 10.6151
R961 B.n511 B.n18 10.6151
R962 B.n511 B.n510 10.6151
R963 B.n510 B.n509 10.6151
R964 B.n509 B.n20 10.6151
R965 B.n505 B.n20 10.6151
R966 B.n505 B.n504 10.6151
R967 B.n504 B.n503 10.6151
R968 B.n503 B.n22 10.6151
R969 B.n499 B.n22 10.6151
R970 B.n499 B.n498 10.6151
R971 B.n498 B.n497 10.6151
R972 B.n497 B.n24 10.6151
R973 B.n493 B.n24 10.6151
R974 B.n493 B.n492 10.6151
R975 B.n492 B.n491 10.6151
R976 B.n491 B.n26 10.6151
R977 B.n487 B.n26 10.6151
R978 B.n487 B.n486 10.6151
R979 B.n486 B.n485 10.6151
R980 B.n485 B.n28 10.6151
R981 B.n481 B.n28 10.6151
R982 B.n464 B.n36 6.5566
R983 B.n452 B.n451 6.5566
R984 B.n244 B.n116 6.5566
R985 B.n257 B.n256 6.5566
R986 B.n467 B.n36 4.05904
R987 B.n451 B.n450 4.05904
R988 B.n241 B.n116 4.05904
R989 B.n258 B.n257 4.05904
R990 B.n563 B.n0 2.81026
R991 B.n563 B.n1 2.81026
R992 VP.n19 VP.n16 161.3
R993 VP.n21 VP.n20 161.3
R994 VP.n22 VP.n15 161.3
R995 VP.n24 VP.n23 161.3
R996 VP.n25 VP.n14 161.3
R997 VP.n27 VP.n26 161.3
R998 VP.n29 VP.n13 161.3
R999 VP.n31 VP.n30 161.3
R1000 VP.n32 VP.n12 161.3
R1001 VP.n34 VP.n33 161.3
R1002 VP.n35 VP.n11 161.3
R1003 VP.n37 VP.n36 161.3
R1004 VP.n69 VP.n68 161.3
R1005 VP.n67 VP.n1 161.3
R1006 VP.n66 VP.n65 161.3
R1007 VP.n64 VP.n2 161.3
R1008 VP.n63 VP.n62 161.3
R1009 VP.n61 VP.n3 161.3
R1010 VP.n59 VP.n58 161.3
R1011 VP.n57 VP.n4 161.3
R1012 VP.n56 VP.n55 161.3
R1013 VP.n54 VP.n5 161.3
R1014 VP.n53 VP.n52 161.3
R1015 VP.n51 VP.n6 161.3
R1016 VP.n50 VP.n49 161.3
R1017 VP.n47 VP.n7 161.3
R1018 VP.n46 VP.n45 161.3
R1019 VP.n44 VP.n8 161.3
R1020 VP.n43 VP.n42 161.3
R1021 VP.n41 VP.n9 161.3
R1022 VP.n40 VP.n39 68.3588
R1023 VP.n70 VP.n0 68.3588
R1024 VP.n38 VP.n10 68.3588
R1025 VP.n18 VP.n17 58.3802
R1026 VP.n55 VP.n54 56.5617
R1027 VP.n23 VP.n22 56.5617
R1028 VP.n46 VP.n8 52.2023
R1029 VP.n66 VP.n2 52.2023
R1030 VP.n34 VP.n12 52.2023
R1031 VP.n39 VP.n38 43.7344
R1032 VP.n18 VP.t4 42.1185
R1033 VP.n42 VP.n8 28.9518
R1034 VP.n67 VP.n66 28.9518
R1035 VP.n35 VP.n34 28.9518
R1036 VP.n42 VP.n41 24.5923
R1037 VP.n47 VP.n46 24.5923
R1038 VP.n49 VP.n47 24.5923
R1039 VP.n53 VP.n6 24.5923
R1040 VP.n54 VP.n53 24.5923
R1041 VP.n55 VP.n4 24.5923
R1042 VP.n59 VP.n4 24.5923
R1043 VP.n62 VP.n61 24.5923
R1044 VP.n62 VP.n2 24.5923
R1045 VP.n68 VP.n67 24.5923
R1046 VP.n36 VP.n35 24.5923
R1047 VP.n23 VP.n14 24.5923
R1048 VP.n27 VP.n14 24.5923
R1049 VP.n30 VP.n29 24.5923
R1050 VP.n30 VP.n12 24.5923
R1051 VP.n21 VP.n16 24.5923
R1052 VP.n22 VP.n21 24.5923
R1053 VP.n41 VP.n40 21.8872
R1054 VP.n68 VP.n0 21.8872
R1055 VP.n36 VP.n10 21.8872
R1056 VP.n48 VP.n6 15.4934
R1057 VP.n60 VP.n59 15.4934
R1058 VP.n28 VP.n27 15.4934
R1059 VP.n17 VP.n16 15.4934
R1060 VP.n40 VP.t1 10.1569
R1061 VP.n48 VP.t5 10.1569
R1062 VP.n60 VP.t6 10.1569
R1063 VP.n0 VP.t3 10.1569
R1064 VP.n10 VP.t2 10.1569
R1065 VP.n28 VP.t7 10.1569
R1066 VP.n17 VP.t0 10.1569
R1067 VP.n49 VP.n48 9.09948
R1068 VP.n61 VP.n60 9.09948
R1069 VP.n29 VP.n28 9.09948
R1070 VP.n19 VP.n18 5.3904
R1071 VP.n38 VP.n37 0.354861
R1072 VP.n39 VP.n9 0.354861
R1073 VP.n70 VP.n69 0.354861
R1074 VP VP.n70 0.267071
R1075 VP.n20 VP.n19 0.189894
R1076 VP.n20 VP.n15 0.189894
R1077 VP.n24 VP.n15 0.189894
R1078 VP.n25 VP.n24 0.189894
R1079 VP.n26 VP.n25 0.189894
R1080 VP.n26 VP.n13 0.189894
R1081 VP.n31 VP.n13 0.189894
R1082 VP.n32 VP.n31 0.189894
R1083 VP.n33 VP.n32 0.189894
R1084 VP.n33 VP.n11 0.189894
R1085 VP.n37 VP.n11 0.189894
R1086 VP.n43 VP.n9 0.189894
R1087 VP.n44 VP.n43 0.189894
R1088 VP.n45 VP.n44 0.189894
R1089 VP.n45 VP.n7 0.189894
R1090 VP.n50 VP.n7 0.189894
R1091 VP.n51 VP.n50 0.189894
R1092 VP.n52 VP.n51 0.189894
R1093 VP.n52 VP.n5 0.189894
R1094 VP.n56 VP.n5 0.189894
R1095 VP.n57 VP.n56 0.189894
R1096 VP.n58 VP.n57 0.189894
R1097 VP.n58 VP.n3 0.189894
R1098 VP.n63 VP.n3 0.189894
R1099 VP.n64 VP.n63 0.189894
R1100 VP.n65 VP.n64 0.189894
R1101 VP.n65 VP.n1 0.189894
R1102 VP.n69 VP.n1 0.189894
R1103 VDD1 VDD1.n0 349.221
R1104 VDD1.n3 VDD1.n2 349.11
R1105 VDD1.n3 VDD1.n1 349.11
R1106 VDD1.n5 VDD1.n4 347.815
R1107 VDD1.n5 VDD1.n3 37.4578
R1108 VDD1.n4 VDD1.t0 27.5471
R1109 VDD1.n4 VDD1.t5 27.5471
R1110 VDD1.n0 VDD1.t3 27.5471
R1111 VDD1.n0 VDD1.t7 27.5471
R1112 VDD1.n2 VDD1.t1 27.5471
R1113 VDD1.n2 VDD1.t4 27.5471
R1114 VDD1.n1 VDD1.t6 27.5471
R1115 VDD1.n1 VDD1.t2 27.5471
R1116 VDD1 VDD1.n5 1.29145
C0 VDD2 w_n4100_n1204# 1.84292f
C1 B VP 2.01728f
C2 B VTAIL 1.32318f
C3 VTAIL VP 2.63424f
C4 VDD1 B 1.41735f
C5 B VN 1.12411f
C6 VDD1 VP 1.67427f
C7 VP VN 5.9103f
C8 VDD1 VTAIL 4.62564f
C9 VTAIL VN 2.62013f
C10 VDD1 VN 0.159207f
C11 B w_n4100_n1204# 7.467471f
C12 w_n4100_n1204# VP 8.75076f
C13 w_n4100_n1204# VTAIL 1.74253f
C14 VDD1 w_n4100_n1204# 1.72083f
C15 w_n4100_n1204# VN 8.22506f
C16 VDD2 B 1.52026f
C17 VDD2 VP 0.549895f
C18 VDD2 VTAIL 4.6814f
C19 VDD1 VDD2 1.88113f
C20 VDD2 VN 1.28737f
C21 VDD2 VSUBS 1.172165f
C22 VDD1 VSUBS 1.824597f
C23 VTAIL VSUBS 0.55195f
C24 VN VSUBS 7.24516f
C25 VP VSUBS 3.174228f
C26 B VSUBS 4.046648f
C27 w_n4100_n1204# VSUBS 63.517197f
C28 VDD1.t3 VSUBS 0.017064f
C29 VDD1.t7 VSUBS 0.017064f
C30 VDD1.n0 VSUBS 0.058455f
C31 VDD1.t6 VSUBS 0.017064f
C32 VDD1.t2 VSUBS 0.017064f
C33 VDD1.n1 VSUBS 0.058302f
C34 VDD1.t1 VSUBS 0.017064f
C35 VDD1.t4 VSUBS 0.017064f
C36 VDD1.n2 VSUBS 0.058302f
C37 VDD1.n3 VSUBS 2.05588f
C38 VDD1.t0 VSUBS 0.017064f
C39 VDD1.t5 VSUBS 0.017064f
C40 VDD1.n4 VSUBS 0.056837f
C41 VDD1.n5 VSUBS 1.61667f
C42 VP.t3 VSUBS 0.431261f
C43 VP.n0 VSUBS 0.507286f
C44 VP.n1 VSUBS 0.064913f
C45 VP.n2 VSUBS 0.115974f
C46 VP.n3 VSUBS 0.064913f
C47 VP.t6 VSUBS 0.431261f
C48 VP.n4 VSUBS 0.120374f
C49 VP.n5 VSUBS 0.064913f
C50 VP.n6 VSUBS 0.098387f
C51 VP.n7 VSUBS 0.064913f
C52 VP.n8 VSUBS 0.065409f
C53 VP.n9 VSUBS 0.104751f
C54 VP.t1 VSUBS 0.431261f
C55 VP.t2 VSUBS 0.431261f
C56 VP.n10 VSUBS 0.507286f
C57 VP.n11 VSUBS 0.064913f
C58 VP.n12 VSUBS 0.115974f
C59 VP.n13 VSUBS 0.064913f
C60 VP.t7 VSUBS 0.431261f
C61 VP.n14 VSUBS 0.120374f
C62 VP.n15 VSUBS 0.064913f
C63 VP.n16 VSUBS 0.098387f
C64 VP.t4 VSUBS 0.945907f
C65 VP.t0 VSUBS 0.431261f
C66 VP.n17 VSUBS 0.465237f
C67 VP.n18 VSUBS 0.468808f
C68 VP.n19 VSUBS 0.68465f
C69 VP.n20 VSUBS 0.064913f
C70 VP.n21 VSUBS 0.120374f
C71 VP.n22 VSUBS 0.09436f
C72 VP.n23 VSUBS 0.09436f
C73 VP.n24 VSUBS 0.064913f
C74 VP.n25 VSUBS 0.064913f
C75 VP.n26 VSUBS 0.064913f
C76 VP.n27 VSUBS 0.098387f
C77 VP.n28 VSUBS 0.259775f
C78 VP.n29 VSUBS 0.082936f
C79 VP.n30 VSUBS 0.120374f
C80 VP.n31 VSUBS 0.064913f
C81 VP.n32 VSUBS 0.064913f
C82 VP.n33 VSUBS 0.064913f
C83 VP.n34 VSUBS 0.065409f
C84 VP.n35 VSUBS 0.127712f
C85 VP.n36 VSUBS 0.113838f
C86 VP.n37 VSUBS 0.104751f
C87 VP.n38 VSUBS 2.99144f
C88 VP.n39 VSUBS 3.04494f
C89 VP.n40 VSUBS 0.507286f
C90 VP.n41 VSUBS 0.113838f
C91 VP.n42 VSUBS 0.127712f
C92 VP.n43 VSUBS 0.064913f
C93 VP.n44 VSUBS 0.064913f
C94 VP.n45 VSUBS 0.064913f
C95 VP.n46 VSUBS 0.115974f
C96 VP.n47 VSUBS 0.120374f
C97 VP.t5 VSUBS 0.431261f
C98 VP.n48 VSUBS 0.259775f
C99 VP.n49 VSUBS 0.082936f
C100 VP.n50 VSUBS 0.064913f
C101 VP.n51 VSUBS 0.064913f
C102 VP.n52 VSUBS 0.064913f
C103 VP.n53 VSUBS 0.120374f
C104 VP.n54 VSUBS 0.09436f
C105 VP.n55 VSUBS 0.09436f
C106 VP.n56 VSUBS 0.064913f
C107 VP.n57 VSUBS 0.064913f
C108 VP.n58 VSUBS 0.064913f
C109 VP.n59 VSUBS 0.098387f
C110 VP.n60 VSUBS 0.259775f
C111 VP.n61 VSUBS 0.082936f
C112 VP.n62 VSUBS 0.120374f
C113 VP.n63 VSUBS 0.064913f
C114 VP.n64 VSUBS 0.064913f
C115 VP.n65 VSUBS 0.064913f
C116 VP.n66 VSUBS 0.065409f
C117 VP.n67 VSUBS 0.127712f
C118 VP.n68 VSUBS 0.113838f
C119 VP.n69 VSUBS 0.104751f
C120 VP.n70 VSUBS 0.125711f
C121 B.n0 VSUBS 0.007761f
C122 B.n1 VSUBS 0.007761f
C123 B.n2 VSUBS 0.012274f
C124 B.n3 VSUBS 0.012274f
C125 B.n4 VSUBS 0.012274f
C126 B.n5 VSUBS 0.012274f
C127 B.n6 VSUBS 0.012274f
C128 B.n7 VSUBS 0.012274f
C129 B.n8 VSUBS 0.012274f
C130 B.n9 VSUBS 0.012274f
C131 B.n10 VSUBS 0.012274f
C132 B.n11 VSUBS 0.012274f
C133 B.n12 VSUBS 0.012274f
C134 B.n13 VSUBS 0.012274f
C135 B.n14 VSUBS 0.012274f
C136 B.n15 VSUBS 0.012274f
C137 B.n16 VSUBS 0.012274f
C138 B.n17 VSUBS 0.012274f
C139 B.n18 VSUBS 0.012274f
C140 B.n19 VSUBS 0.012274f
C141 B.n20 VSUBS 0.012274f
C142 B.n21 VSUBS 0.012274f
C143 B.n22 VSUBS 0.012274f
C144 B.n23 VSUBS 0.012274f
C145 B.n24 VSUBS 0.012274f
C146 B.n25 VSUBS 0.012274f
C147 B.n26 VSUBS 0.012274f
C148 B.n27 VSUBS 0.012274f
C149 B.n28 VSUBS 0.012274f
C150 B.n29 VSUBS 0.030676f
C151 B.n30 VSUBS 0.012274f
C152 B.n31 VSUBS 0.012274f
C153 B.n32 VSUBS 0.012274f
C154 B.n33 VSUBS 0.012274f
C155 B.t2 VSUBS 0.03901f
C156 B.t1 VSUBS 0.049083f
C157 B.t0 VSUBS 0.29293f
C158 B.n34 VSUBS 0.113552f
C159 B.n35 VSUBS 0.088094f
C160 B.n36 VSUBS 0.028437f
C161 B.n37 VSUBS 0.012274f
C162 B.n38 VSUBS 0.012274f
C163 B.n39 VSUBS 0.012274f
C164 B.n40 VSUBS 0.012274f
C165 B.n41 VSUBS 0.012274f
C166 B.t5 VSUBS 0.03901f
C167 B.t4 VSUBS 0.049083f
C168 B.t3 VSUBS 0.29293f
C169 B.n42 VSUBS 0.113552f
C170 B.n43 VSUBS 0.088094f
C171 B.n44 VSUBS 0.012274f
C172 B.n45 VSUBS 0.012274f
C173 B.n46 VSUBS 0.012274f
C174 B.n47 VSUBS 0.012274f
C175 B.n48 VSUBS 0.030609f
C176 B.n49 VSUBS 0.012274f
C177 B.n50 VSUBS 0.012274f
C178 B.n51 VSUBS 0.012274f
C179 B.n52 VSUBS 0.012274f
C180 B.n53 VSUBS 0.012274f
C181 B.n54 VSUBS 0.012274f
C182 B.n55 VSUBS 0.012274f
C183 B.n56 VSUBS 0.012274f
C184 B.n57 VSUBS 0.012274f
C185 B.n58 VSUBS 0.012274f
C186 B.n59 VSUBS 0.012274f
C187 B.n60 VSUBS 0.012274f
C188 B.n61 VSUBS 0.012274f
C189 B.n62 VSUBS 0.012274f
C190 B.n63 VSUBS 0.012274f
C191 B.n64 VSUBS 0.012274f
C192 B.n65 VSUBS 0.012274f
C193 B.n66 VSUBS 0.012274f
C194 B.n67 VSUBS 0.012274f
C195 B.n68 VSUBS 0.012274f
C196 B.n69 VSUBS 0.012274f
C197 B.n70 VSUBS 0.012274f
C198 B.n71 VSUBS 0.012274f
C199 B.n72 VSUBS 0.012274f
C200 B.n73 VSUBS 0.012274f
C201 B.n74 VSUBS 0.012274f
C202 B.n75 VSUBS 0.012274f
C203 B.n76 VSUBS 0.012274f
C204 B.n77 VSUBS 0.012274f
C205 B.n78 VSUBS 0.012274f
C206 B.n79 VSUBS 0.012274f
C207 B.n80 VSUBS 0.012274f
C208 B.n81 VSUBS 0.012274f
C209 B.n82 VSUBS 0.012274f
C210 B.n83 VSUBS 0.012274f
C211 B.n84 VSUBS 0.012274f
C212 B.n85 VSUBS 0.012274f
C213 B.n86 VSUBS 0.012274f
C214 B.n87 VSUBS 0.012274f
C215 B.n88 VSUBS 0.012274f
C216 B.n89 VSUBS 0.012274f
C217 B.n90 VSUBS 0.012274f
C218 B.n91 VSUBS 0.012274f
C219 B.n92 VSUBS 0.012274f
C220 B.n93 VSUBS 0.012274f
C221 B.n94 VSUBS 0.012274f
C222 B.n95 VSUBS 0.012274f
C223 B.n96 VSUBS 0.012274f
C224 B.n97 VSUBS 0.012274f
C225 B.n98 VSUBS 0.012274f
C226 B.n99 VSUBS 0.012274f
C227 B.n100 VSUBS 0.012274f
C228 B.n101 VSUBS 0.012274f
C229 B.n102 VSUBS 0.029249f
C230 B.n103 VSUBS 0.012274f
C231 B.n104 VSUBS 0.012274f
C232 B.n105 VSUBS 0.012274f
C233 B.n106 VSUBS 0.012274f
C234 B.n107 VSUBS 0.012274f
C235 B.t7 VSUBS 0.03901f
C236 B.t8 VSUBS 0.049083f
C237 B.t6 VSUBS 0.29293f
C238 B.n108 VSUBS 0.113552f
C239 B.n109 VSUBS 0.088094f
C240 B.n110 VSUBS 0.012274f
C241 B.n111 VSUBS 0.012274f
C242 B.n112 VSUBS 0.012274f
C243 B.n113 VSUBS 0.012274f
C244 B.t10 VSUBS 0.03901f
C245 B.t11 VSUBS 0.049083f
C246 B.t9 VSUBS 0.29293f
C247 B.n114 VSUBS 0.113552f
C248 B.n115 VSUBS 0.088094f
C249 B.n116 VSUBS 0.028437f
C250 B.n117 VSUBS 0.012274f
C251 B.n118 VSUBS 0.012274f
C252 B.n119 VSUBS 0.012274f
C253 B.n120 VSUBS 0.012274f
C254 B.n121 VSUBS 0.030676f
C255 B.n122 VSUBS 0.012274f
C256 B.n123 VSUBS 0.012274f
C257 B.n124 VSUBS 0.012274f
C258 B.n125 VSUBS 0.012274f
C259 B.n126 VSUBS 0.012274f
C260 B.n127 VSUBS 0.012274f
C261 B.n128 VSUBS 0.012274f
C262 B.n129 VSUBS 0.012274f
C263 B.n130 VSUBS 0.012274f
C264 B.n131 VSUBS 0.012274f
C265 B.n132 VSUBS 0.012274f
C266 B.n133 VSUBS 0.012274f
C267 B.n134 VSUBS 0.012274f
C268 B.n135 VSUBS 0.012274f
C269 B.n136 VSUBS 0.012274f
C270 B.n137 VSUBS 0.012274f
C271 B.n138 VSUBS 0.012274f
C272 B.n139 VSUBS 0.012274f
C273 B.n140 VSUBS 0.012274f
C274 B.n141 VSUBS 0.012274f
C275 B.n142 VSUBS 0.012274f
C276 B.n143 VSUBS 0.012274f
C277 B.n144 VSUBS 0.012274f
C278 B.n145 VSUBS 0.012274f
C279 B.n146 VSUBS 0.012274f
C280 B.n147 VSUBS 0.012274f
C281 B.n148 VSUBS 0.012274f
C282 B.n149 VSUBS 0.012274f
C283 B.n150 VSUBS 0.012274f
C284 B.n151 VSUBS 0.012274f
C285 B.n152 VSUBS 0.012274f
C286 B.n153 VSUBS 0.012274f
C287 B.n154 VSUBS 0.012274f
C288 B.n155 VSUBS 0.012274f
C289 B.n156 VSUBS 0.012274f
C290 B.n157 VSUBS 0.012274f
C291 B.n158 VSUBS 0.012274f
C292 B.n159 VSUBS 0.012274f
C293 B.n160 VSUBS 0.012274f
C294 B.n161 VSUBS 0.012274f
C295 B.n162 VSUBS 0.012274f
C296 B.n163 VSUBS 0.012274f
C297 B.n164 VSUBS 0.012274f
C298 B.n165 VSUBS 0.012274f
C299 B.n166 VSUBS 0.012274f
C300 B.n167 VSUBS 0.012274f
C301 B.n168 VSUBS 0.012274f
C302 B.n169 VSUBS 0.012274f
C303 B.n170 VSUBS 0.012274f
C304 B.n171 VSUBS 0.012274f
C305 B.n172 VSUBS 0.012274f
C306 B.n173 VSUBS 0.012274f
C307 B.n174 VSUBS 0.012274f
C308 B.n175 VSUBS 0.012274f
C309 B.n176 VSUBS 0.012274f
C310 B.n177 VSUBS 0.012274f
C311 B.n178 VSUBS 0.012274f
C312 B.n179 VSUBS 0.012274f
C313 B.n180 VSUBS 0.012274f
C314 B.n181 VSUBS 0.012274f
C315 B.n182 VSUBS 0.012274f
C316 B.n183 VSUBS 0.012274f
C317 B.n184 VSUBS 0.012274f
C318 B.n185 VSUBS 0.012274f
C319 B.n186 VSUBS 0.012274f
C320 B.n187 VSUBS 0.012274f
C321 B.n188 VSUBS 0.012274f
C322 B.n189 VSUBS 0.012274f
C323 B.n190 VSUBS 0.012274f
C324 B.n191 VSUBS 0.012274f
C325 B.n192 VSUBS 0.012274f
C326 B.n193 VSUBS 0.012274f
C327 B.n194 VSUBS 0.012274f
C328 B.n195 VSUBS 0.012274f
C329 B.n196 VSUBS 0.012274f
C330 B.n197 VSUBS 0.012274f
C331 B.n198 VSUBS 0.012274f
C332 B.n199 VSUBS 0.012274f
C333 B.n200 VSUBS 0.012274f
C334 B.n201 VSUBS 0.012274f
C335 B.n202 VSUBS 0.012274f
C336 B.n203 VSUBS 0.012274f
C337 B.n204 VSUBS 0.012274f
C338 B.n205 VSUBS 0.012274f
C339 B.n206 VSUBS 0.012274f
C340 B.n207 VSUBS 0.012274f
C341 B.n208 VSUBS 0.012274f
C342 B.n209 VSUBS 0.012274f
C343 B.n210 VSUBS 0.012274f
C344 B.n211 VSUBS 0.012274f
C345 B.n212 VSUBS 0.012274f
C346 B.n213 VSUBS 0.012274f
C347 B.n214 VSUBS 0.012274f
C348 B.n215 VSUBS 0.012274f
C349 B.n216 VSUBS 0.012274f
C350 B.n217 VSUBS 0.012274f
C351 B.n218 VSUBS 0.012274f
C352 B.n219 VSUBS 0.012274f
C353 B.n220 VSUBS 0.012274f
C354 B.n221 VSUBS 0.012274f
C355 B.n222 VSUBS 0.012274f
C356 B.n223 VSUBS 0.012274f
C357 B.n224 VSUBS 0.012274f
C358 B.n225 VSUBS 0.012274f
C359 B.n226 VSUBS 0.029249f
C360 B.n227 VSUBS 0.029249f
C361 B.n228 VSUBS 0.030676f
C362 B.n229 VSUBS 0.012274f
C363 B.n230 VSUBS 0.012274f
C364 B.n231 VSUBS 0.012274f
C365 B.n232 VSUBS 0.012274f
C366 B.n233 VSUBS 0.012274f
C367 B.n234 VSUBS 0.012274f
C368 B.n235 VSUBS 0.012274f
C369 B.n236 VSUBS 0.012274f
C370 B.n237 VSUBS 0.012274f
C371 B.n238 VSUBS 0.012274f
C372 B.n239 VSUBS 0.012274f
C373 B.n240 VSUBS 0.012274f
C374 B.n241 VSUBS 0.008483f
C375 B.n242 VSUBS 0.012274f
C376 B.n243 VSUBS 0.012274f
C377 B.n244 VSUBS 0.009927f
C378 B.n245 VSUBS 0.012274f
C379 B.n246 VSUBS 0.012274f
C380 B.n247 VSUBS 0.012274f
C381 B.n248 VSUBS 0.012274f
C382 B.n249 VSUBS 0.012274f
C383 B.n250 VSUBS 0.012274f
C384 B.n251 VSUBS 0.012274f
C385 B.n252 VSUBS 0.012274f
C386 B.n253 VSUBS 0.012274f
C387 B.n254 VSUBS 0.012274f
C388 B.n255 VSUBS 0.012274f
C389 B.n256 VSUBS 0.009927f
C390 B.n257 VSUBS 0.028437f
C391 B.n258 VSUBS 0.008483f
C392 B.n259 VSUBS 0.012274f
C393 B.n260 VSUBS 0.012274f
C394 B.n261 VSUBS 0.012274f
C395 B.n262 VSUBS 0.012274f
C396 B.n263 VSUBS 0.012274f
C397 B.n264 VSUBS 0.012274f
C398 B.n265 VSUBS 0.012274f
C399 B.n266 VSUBS 0.012274f
C400 B.n267 VSUBS 0.012274f
C401 B.n268 VSUBS 0.012274f
C402 B.n269 VSUBS 0.012274f
C403 B.n270 VSUBS 0.012274f
C404 B.n271 VSUBS 0.030676f
C405 B.n272 VSUBS 0.030676f
C406 B.n273 VSUBS 0.029249f
C407 B.n274 VSUBS 0.012274f
C408 B.n275 VSUBS 0.012274f
C409 B.n276 VSUBS 0.012274f
C410 B.n277 VSUBS 0.012274f
C411 B.n278 VSUBS 0.012274f
C412 B.n279 VSUBS 0.012274f
C413 B.n280 VSUBS 0.012274f
C414 B.n281 VSUBS 0.012274f
C415 B.n282 VSUBS 0.012274f
C416 B.n283 VSUBS 0.012274f
C417 B.n284 VSUBS 0.012274f
C418 B.n285 VSUBS 0.012274f
C419 B.n286 VSUBS 0.012274f
C420 B.n287 VSUBS 0.012274f
C421 B.n288 VSUBS 0.012274f
C422 B.n289 VSUBS 0.012274f
C423 B.n290 VSUBS 0.012274f
C424 B.n291 VSUBS 0.012274f
C425 B.n292 VSUBS 0.012274f
C426 B.n293 VSUBS 0.012274f
C427 B.n294 VSUBS 0.012274f
C428 B.n295 VSUBS 0.012274f
C429 B.n296 VSUBS 0.012274f
C430 B.n297 VSUBS 0.012274f
C431 B.n298 VSUBS 0.012274f
C432 B.n299 VSUBS 0.012274f
C433 B.n300 VSUBS 0.012274f
C434 B.n301 VSUBS 0.012274f
C435 B.n302 VSUBS 0.012274f
C436 B.n303 VSUBS 0.012274f
C437 B.n304 VSUBS 0.012274f
C438 B.n305 VSUBS 0.012274f
C439 B.n306 VSUBS 0.012274f
C440 B.n307 VSUBS 0.012274f
C441 B.n308 VSUBS 0.012274f
C442 B.n309 VSUBS 0.012274f
C443 B.n310 VSUBS 0.012274f
C444 B.n311 VSUBS 0.012274f
C445 B.n312 VSUBS 0.012274f
C446 B.n313 VSUBS 0.012274f
C447 B.n314 VSUBS 0.012274f
C448 B.n315 VSUBS 0.012274f
C449 B.n316 VSUBS 0.012274f
C450 B.n317 VSUBS 0.012274f
C451 B.n318 VSUBS 0.012274f
C452 B.n319 VSUBS 0.012274f
C453 B.n320 VSUBS 0.012274f
C454 B.n321 VSUBS 0.012274f
C455 B.n322 VSUBS 0.012274f
C456 B.n323 VSUBS 0.012274f
C457 B.n324 VSUBS 0.012274f
C458 B.n325 VSUBS 0.012274f
C459 B.n326 VSUBS 0.012274f
C460 B.n327 VSUBS 0.012274f
C461 B.n328 VSUBS 0.012274f
C462 B.n329 VSUBS 0.012274f
C463 B.n330 VSUBS 0.012274f
C464 B.n331 VSUBS 0.012274f
C465 B.n332 VSUBS 0.012274f
C466 B.n333 VSUBS 0.012274f
C467 B.n334 VSUBS 0.012274f
C468 B.n335 VSUBS 0.012274f
C469 B.n336 VSUBS 0.012274f
C470 B.n337 VSUBS 0.012274f
C471 B.n338 VSUBS 0.012274f
C472 B.n339 VSUBS 0.012274f
C473 B.n340 VSUBS 0.012274f
C474 B.n341 VSUBS 0.012274f
C475 B.n342 VSUBS 0.012274f
C476 B.n343 VSUBS 0.012274f
C477 B.n344 VSUBS 0.012274f
C478 B.n345 VSUBS 0.012274f
C479 B.n346 VSUBS 0.012274f
C480 B.n347 VSUBS 0.012274f
C481 B.n348 VSUBS 0.012274f
C482 B.n349 VSUBS 0.012274f
C483 B.n350 VSUBS 0.012274f
C484 B.n351 VSUBS 0.012274f
C485 B.n352 VSUBS 0.012274f
C486 B.n353 VSUBS 0.012274f
C487 B.n354 VSUBS 0.012274f
C488 B.n355 VSUBS 0.012274f
C489 B.n356 VSUBS 0.012274f
C490 B.n357 VSUBS 0.012274f
C491 B.n358 VSUBS 0.012274f
C492 B.n359 VSUBS 0.012274f
C493 B.n360 VSUBS 0.012274f
C494 B.n361 VSUBS 0.012274f
C495 B.n362 VSUBS 0.012274f
C496 B.n363 VSUBS 0.012274f
C497 B.n364 VSUBS 0.012274f
C498 B.n365 VSUBS 0.012274f
C499 B.n366 VSUBS 0.012274f
C500 B.n367 VSUBS 0.012274f
C501 B.n368 VSUBS 0.012274f
C502 B.n369 VSUBS 0.012274f
C503 B.n370 VSUBS 0.012274f
C504 B.n371 VSUBS 0.012274f
C505 B.n372 VSUBS 0.012274f
C506 B.n373 VSUBS 0.012274f
C507 B.n374 VSUBS 0.012274f
C508 B.n375 VSUBS 0.012274f
C509 B.n376 VSUBS 0.012274f
C510 B.n377 VSUBS 0.012274f
C511 B.n378 VSUBS 0.012274f
C512 B.n379 VSUBS 0.012274f
C513 B.n380 VSUBS 0.012274f
C514 B.n381 VSUBS 0.012274f
C515 B.n382 VSUBS 0.012274f
C516 B.n383 VSUBS 0.012274f
C517 B.n384 VSUBS 0.012274f
C518 B.n385 VSUBS 0.012274f
C519 B.n386 VSUBS 0.012274f
C520 B.n387 VSUBS 0.012274f
C521 B.n388 VSUBS 0.012274f
C522 B.n389 VSUBS 0.012274f
C523 B.n390 VSUBS 0.012274f
C524 B.n391 VSUBS 0.012274f
C525 B.n392 VSUBS 0.012274f
C526 B.n393 VSUBS 0.012274f
C527 B.n394 VSUBS 0.012274f
C528 B.n395 VSUBS 0.012274f
C529 B.n396 VSUBS 0.012274f
C530 B.n397 VSUBS 0.012274f
C531 B.n398 VSUBS 0.012274f
C532 B.n399 VSUBS 0.012274f
C533 B.n400 VSUBS 0.012274f
C534 B.n401 VSUBS 0.012274f
C535 B.n402 VSUBS 0.012274f
C536 B.n403 VSUBS 0.012274f
C537 B.n404 VSUBS 0.012274f
C538 B.n405 VSUBS 0.012274f
C539 B.n406 VSUBS 0.012274f
C540 B.n407 VSUBS 0.012274f
C541 B.n408 VSUBS 0.012274f
C542 B.n409 VSUBS 0.012274f
C543 B.n410 VSUBS 0.012274f
C544 B.n411 VSUBS 0.012274f
C545 B.n412 VSUBS 0.012274f
C546 B.n413 VSUBS 0.012274f
C547 B.n414 VSUBS 0.012274f
C548 B.n415 VSUBS 0.012274f
C549 B.n416 VSUBS 0.012274f
C550 B.n417 VSUBS 0.012274f
C551 B.n418 VSUBS 0.012274f
C552 B.n419 VSUBS 0.012274f
C553 B.n420 VSUBS 0.012274f
C554 B.n421 VSUBS 0.012274f
C555 B.n422 VSUBS 0.012274f
C556 B.n423 VSUBS 0.012274f
C557 B.n424 VSUBS 0.012274f
C558 B.n425 VSUBS 0.012274f
C559 B.n426 VSUBS 0.012274f
C560 B.n427 VSUBS 0.012274f
C561 B.n428 VSUBS 0.012274f
C562 B.n429 VSUBS 0.012274f
C563 B.n430 VSUBS 0.012274f
C564 B.n431 VSUBS 0.012274f
C565 B.n432 VSUBS 0.012274f
C566 B.n433 VSUBS 0.012274f
C567 B.n434 VSUBS 0.012274f
C568 B.n435 VSUBS 0.029249f
C569 B.n436 VSUBS 0.030676f
C570 B.n437 VSUBS 0.029315f
C571 B.n438 VSUBS 0.012274f
C572 B.n439 VSUBS 0.012274f
C573 B.n440 VSUBS 0.012274f
C574 B.n441 VSUBS 0.012274f
C575 B.n442 VSUBS 0.012274f
C576 B.n443 VSUBS 0.012274f
C577 B.n444 VSUBS 0.012274f
C578 B.n445 VSUBS 0.012274f
C579 B.n446 VSUBS 0.012274f
C580 B.n447 VSUBS 0.012274f
C581 B.n448 VSUBS 0.012274f
C582 B.n449 VSUBS 0.012274f
C583 B.n450 VSUBS 0.008483f
C584 B.n451 VSUBS 0.028437f
C585 B.n452 VSUBS 0.009927f
C586 B.n453 VSUBS 0.012274f
C587 B.n454 VSUBS 0.012274f
C588 B.n455 VSUBS 0.012274f
C589 B.n456 VSUBS 0.012274f
C590 B.n457 VSUBS 0.012274f
C591 B.n458 VSUBS 0.012274f
C592 B.n459 VSUBS 0.012274f
C593 B.n460 VSUBS 0.012274f
C594 B.n461 VSUBS 0.012274f
C595 B.n462 VSUBS 0.012274f
C596 B.n463 VSUBS 0.012274f
C597 B.n464 VSUBS 0.009927f
C598 B.n465 VSUBS 0.012274f
C599 B.n466 VSUBS 0.012274f
C600 B.n467 VSUBS 0.008483f
C601 B.n468 VSUBS 0.012274f
C602 B.n469 VSUBS 0.012274f
C603 B.n470 VSUBS 0.012274f
C604 B.n471 VSUBS 0.012274f
C605 B.n472 VSUBS 0.012274f
C606 B.n473 VSUBS 0.012274f
C607 B.n474 VSUBS 0.012274f
C608 B.n475 VSUBS 0.012274f
C609 B.n476 VSUBS 0.012274f
C610 B.n477 VSUBS 0.012274f
C611 B.n478 VSUBS 0.012274f
C612 B.n479 VSUBS 0.012274f
C613 B.n480 VSUBS 0.030676f
C614 B.n481 VSUBS 0.029249f
C615 B.n482 VSUBS 0.029249f
C616 B.n483 VSUBS 0.012274f
C617 B.n484 VSUBS 0.012274f
C618 B.n485 VSUBS 0.012274f
C619 B.n486 VSUBS 0.012274f
C620 B.n487 VSUBS 0.012274f
C621 B.n488 VSUBS 0.012274f
C622 B.n489 VSUBS 0.012274f
C623 B.n490 VSUBS 0.012274f
C624 B.n491 VSUBS 0.012274f
C625 B.n492 VSUBS 0.012274f
C626 B.n493 VSUBS 0.012274f
C627 B.n494 VSUBS 0.012274f
C628 B.n495 VSUBS 0.012274f
C629 B.n496 VSUBS 0.012274f
C630 B.n497 VSUBS 0.012274f
C631 B.n498 VSUBS 0.012274f
C632 B.n499 VSUBS 0.012274f
C633 B.n500 VSUBS 0.012274f
C634 B.n501 VSUBS 0.012274f
C635 B.n502 VSUBS 0.012274f
C636 B.n503 VSUBS 0.012274f
C637 B.n504 VSUBS 0.012274f
C638 B.n505 VSUBS 0.012274f
C639 B.n506 VSUBS 0.012274f
C640 B.n507 VSUBS 0.012274f
C641 B.n508 VSUBS 0.012274f
C642 B.n509 VSUBS 0.012274f
C643 B.n510 VSUBS 0.012274f
C644 B.n511 VSUBS 0.012274f
C645 B.n512 VSUBS 0.012274f
C646 B.n513 VSUBS 0.012274f
C647 B.n514 VSUBS 0.012274f
C648 B.n515 VSUBS 0.012274f
C649 B.n516 VSUBS 0.012274f
C650 B.n517 VSUBS 0.012274f
C651 B.n518 VSUBS 0.012274f
C652 B.n519 VSUBS 0.012274f
C653 B.n520 VSUBS 0.012274f
C654 B.n521 VSUBS 0.012274f
C655 B.n522 VSUBS 0.012274f
C656 B.n523 VSUBS 0.012274f
C657 B.n524 VSUBS 0.012274f
C658 B.n525 VSUBS 0.012274f
C659 B.n526 VSUBS 0.012274f
C660 B.n527 VSUBS 0.012274f
C661 B.n528 VSUBS 0.012274f
C662 B.n529 VSUBS 0.012274f
C663 B.n530 VSUBS 0.012274f
C664 B.n531 VSUBS 0.012274f
C665 B.n532 VSUBS 0.012274f
C666 B.n533 VSUBS 0.012274f
C667 B.n534 VSUBS 0.012274f
C668 B.n535 VSUBS 0.012274f
C669 B.n536 VSUBS 0.012274f
C670 B.n537 VSUBS 0.012274f
C671 B.n538 VSUBS 0.012274f
C672 B.n539 VSUBS 0.012274f
C673 B.n540 VSUBS 0.012274f
C674 B.n541 VSUBS 0.012274f
C675 B.n542 VSUBS 0.012274f
C676 B.n543 VSUBS 0.012274f
C677 B.n544 VSUBS 0.012274f
C678 B.n545 VSUBS 0.012274f
C679 B.n546 VSUBS 0.012274f
C680 B.n547 VSUBS 0.012274f
C681 B.n548 VSUBS 0.012274f
C682 B.n549 VSUBS 0.012274f
C683 B.n550 VSUBS 0.012274f
C684 B.n551 VSUBS 0.012274f
C685 B.n552 VSUBS 0.012274f
C686 B.n553 VSUBS 0.012274f
C687 B.n554 VSUBS 0.012274f
C688 B.n555 VSUBS 0.012274f
C689 B.n556 VSUBS 0.012274f
C690 B.n557 VSUBS 0.012274f
C691 B.n558 VSUBS 0.012274f
C692 B.n559 VSUBS 0.012274f
C693 B.n560 VSUBS 0.012274f
C694 B.n561 VSUBS 0.012274f
C695 B.n562 VSUBS 0.012274f
C696 B.n563 VSUBS 0.027792f
C697 VDD2.t3 VSUBS 0.017695f
C698 VDD2.t0 VSUBS 0.017695f
C699 VDD2.n0 VSUBS 0.060457f
C700 VDD2.t2 VSUBS 0.017695f
C701 VDD2.t5 VSUBS 0.017695f
C702 VDD2.n1 VSUBS 0.060457f
C703 VDD2.n2 VSUBS 2.0923f
C704 VDD2.t1 VSUBS 0.017695f
C705 VDD2.t7 VSUBS 0.017695f
C706 VDD2.n3 VSUBS 0.058939f
C707 VDD2.n4 VSUBS 1.65307f
C708 VDD2.t6 VSUBS 0.017695f
C709 VDD2.t4 VSUBS 0.017695f
C710 VDD2.n5 VSUBS 0.060452f
C711 VTAIL.t13 VSUBS 0.034153f
C712 VTAIL.t15 VSUBS 0.034153f
C713 VTAIL.n0 VSUBS 0.098775f
C714 VTAIL.n1 VSUBS 0.594922f
C715 VTAIL.t12 VSUBS 0.172562f
C716 VTAIL.n2 VSUBS 0.662861f
C717 VTAIL.t7 VSUBS 0.172562f
C718 VTAIL.n3 VSUBS 0.662861f
C719 VTAIL.t3 VSUBS 0.034153f
C720 VTAIL.t2 VSUBS 0.034153f
C721 VTAIL.n4 VSUBS 0.098775f
C722 VTAIL.n5 VSUBS 0.9065f
C723 VTAIL.t0 VSUBS 0.172562f
C724 VTAIL.n6 VSUBS 1.54343f
C725 VTAIL.t11 VSUBS 0.172562f
C726 VTAIL.n7 VSUBS 1.54344f
C727 VTAIL.t8 VSUBS 0.034153f
C728 VTAIL.t9 VSUBS 0.034153f
C729 VTAIL.n8 VSUBS 0.098775f
C730 VTAIL.n9 VSUBS 0.9065f
C731 VTAIL.t14 VSUBS 0.172562f
C732 VTAIL.n10 VSUBS 0.662861f
C733 VTAIL.t6 VSUBS 0.172562f
C734 VTAIL.n11 VSUBS 0.662861f
C735 VTAIL.t4 VSUBS 0.034153f
C736 VTAIL.t5 VSUBS 0.034153f
C737 VTAIL.n12 VSUBS 0.098775f
C738 VTAIL.n13 VSUBS 0.9065f
C739 VTAIL.t1 VSUBS 0.172562f
C740 VTAIL.n14 VSUBS 1.54343f
C741 VTAIL.t10 VSUBS 0.172562f
C742 VTAIL.n15 VSUBS 1.53657f
C743 VN.t2 VSUBS 0.371408f
C744 VN.n0 VSUBS 0.436881f
C745 VN.n1 VSUBS 0.055904f
C746 VN.n2 VSUBS 0.099878f
C747 VN.n3 VSUBS 0.055904f
C748 VN.t5 VSUBS 0.371408f
C749 VN.n4 VSUBS 0.103668f
C750 VN.n5 VSUBS 0.055904f
C751 VN.n6 VSUBS 0.084732f
C752 VN.t7 VSUBS 0.371408f
C753 VN.n7 VSUBS 0.400668f
C754 VN.t4 VSUBS 0.81463f
C755 VN.n8 VSUBS 0.403743f
C756 VN.n9 VSUBS 0.589628f
C757 VN.n10 VSUBS 0.055904f
C758 VN.n11 VSUBS 0.103668f
C759 VN.n12 VSUBS 0.081265f
C760 VN.n13 VSUBS 0.081265f
C761 VN.n14 VSUBS 0.055904f
C762 VN.n15 VSUBS 0.055904f
C763 VN.n16 VSUBS 0.055904f
C764 VN.n17 VSUBS 0.084732f
C765 VN.n18 VSUBS 0.223722f
C766 VN.n19 VSUBS 0.071426f
C767 VN.n20 VSUBS 0.103668f
C768 VN.n21 VSUBS 0.055904f
C769 VN.n22 VSUBS 0.055904f
C770 VN.n23 VSUBS 0.055904f
C771 VN.n24 VSUBS 0.056331f
C772 VN.n25 VSUBS 0.109987f
C773 VN.n26 VSUBS 0.098038f
C774 VN.n27 VSUBS 0.090213f
C775 VN.n28 VSUBS 0.108264f
C776 VN.t6 VSUBS 0.371408f
C777 VN.n29 VSUBS 0.436881f
C778 VN.n30 VSUBS 0.055904f
C779 VN.n31 VSUBS 0.099878f
C780 VN.n32 VSUBS 0.055904f
C781 VN.t0 VSUBS 0.371408f
C782 VN.n33 VSUBS 0.103668f
C783 VN.n34 VSUBS 0.055904f
C784 VN.n35 VSUBS 0.084732f
C785 VN.t3 VSUBS 0.81463f
C786 VN.t1 VSUBS 0.371408f
C787 VN.n36 VSUBS 0.400668f
C788 VN.n37 VSUBS 0.403742f
C789 VN.n38 VSUBS 0.589628f
C790 VN.n39 VSUBS 0.055904f
C791 VN.n40 VSUBS 0.103668f
C792 VN.n41 VSUBS 0.081265f
C793 VN.n42 VSUBS 0.081265f
C794 VN.n43 VSUBS 0.055904f
C795 VN.n44 VSUBS 0.055904f
C796 VN.n45 VSUBS 0.055904f
C797 VN.n46 VSUBS 0.084732f
C798 VN.n47 VSUBS 0.223722f
C799 VN.n48 VSUBS 0.071426f
C800 VN.n49 VSUBS 0.103668f
C801 VN.n50 VSUBS 0.055904f
C802 VN.n51 VSUBS 0.055904f
C803 VN.n52 VSUBS 0.055904f
C804 VN.n53 VSUBS 0.056331f
C805 VN.n54 VSUBS 0.109987f
C806 VN.n55 VSUBS 0.098038f
C807 VN.n56 VSUBS 0.090213f
C808 VN.n57 VSUBS 2.60028f
.ends

