* NGSPICE file created from diff_pair_sample_0359.ext - technology: sky130A

.subckt diff_pair_sample_0359 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.91555 pd=18 as=6.8913 ps=36.12 w=17.67 l=4
X1 VTAIL.t5 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=2.91555 ps=18 w=17.67 l=4
X2 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=2.91555 ps=18 w=17.67 l=4
X3 VTAIL.t4 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=2.91555 ps=18 w=17.67 l=4
X4 VDD1.t0 VP.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.91555 pd=18 as=6.8913 ps=36.12 w=17.67 l=4
X5 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=0 ps=0 w=17.67 l=4
X6 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=0 ps=0 w=17.67 l=4
X7 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=2.91555 ps=18 w=17.67 l=4
X8 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.91555 pd=18 as=6.8913 ps=36.12 w=17.67 l=4
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=0 ps=0 w=17.67 l=4
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8913 pd=36.12 as=0 ps=0 w=17.67 l=4
X11 VDD2.t0 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.91555 pd=18 as=6.8913 ps=36.12 w=17.67 l=4
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n4 VP.t1 140.243
R9 VP.n4 VP.t3 138.797
R10 VP.n6 VP.t2 106.463
R11 VP.n19 VP.t0 106.463
R12 VP.n6 VP.n5 61.8742
R13 VP.n20 VP.n19 61.8742
R14 VP.n5 VP.n4 56.7559
R15 VP.n13 VP.n12 56.5193
R16 VP.n7 VP.n3 24.4675
R17 VP.n11 VP.n3 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n13 VP.n1 24.4675
R20 VP.n17 VP.n1 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n7 VP.n6 20.3081
R23 VP.n19 VP.n18 20.3081
R24 VP.n8 VP.n5 0.417535
R25 VP.n20 VP.n0 0.417535
R26 VP VP.n20 0.394291
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VTAIL.n778 VTAIL.n686 289.615
R35 VTAIL.n92 VTAIL.n0 289.615
R36 VTAIL.n190 VTAIL.n98 289.615
R37 VTAIL.n288 VTAIL.n196 289.615
R38 VTAIL.n680 VTAIL.n588 289.615
R39 VTAIL.n582 VTAIL.n490 289.615
R40 VTAIL.n484 VTAIL.n392 289.615
R41 VTAIL.n386 VTAIL.n294 289.615
R42 VTAIL.n719 VTAIL.n718 185
R43 VTAIL.n721 VTAIL.n720 185
R44 VTAIL.n714 VTAIL.n713 185
R45 VTAIL.n727 VTAIL.n726 185
R46 VTAIL.n729 VTAIL.n728 185
R47 VTAIL.n710 VTAIL.n709 185
R48 VTAIL.n735 VTAIL.n734 185
R49 VTAIL.n737 VTAIL.n736 185
R50 VTAIL.n706 VTAIL.n705 185
R51 VTAIL.n743 VTAIL.n742 185
R52 VTAIL.n745 VTAIL.n744 185
R53 VTAIL.n702 VTAIL.n701 185
R54 VTAIL.n751 VTAIL.n750 185
R55 VTAIL.n753 VTAIL.n752 185
R56 VTAIL.n698 VTAIL.n697 185
R57 VTAIL.n760 VTAIL.n759 185
R58 VTAIL.n761 VTAIL.n696 185
R59 VTAIL.n763 VTAIL.n762 185
R60 VTAIL.n694 VTAIL.n693 185
R61 VTAIL.n769 VTAIL.n768 185
R62 VTAIL.n771 VTAIL.n770 185
R63 VTAIL.n690 VTAIL.n689 185
R64 VTAIL.n777 VTAIL.n776 185
R65 VTAIL.n779 VTAIL.n778 185
R66 VTAIL.n33 VTAIL.n32 185
R67 VTAIL.n35 VTAIL.n34 185
R68 VTAIL.n28 VTAIL.n27 185
R69 VTAIL.n41 VTAIL.n40 185
R70 VTAIL.n43 VTAIL.n42 185
R71 VTAIL.n24 VTAIL.n23 185
R72 VTAIL.n49 VTAIL.n48 185
R73 VTAIL.n51 VTAIL.n50 185
R74 VTAIL.n20 VTAIL.n19 185
R75 VTAIL.n57 VTAIL.n56 185
R76 VTAIL.n59 VTAIL.n58 185
R77 VTAIL.n16 VTAIL.n15 185
R78 VTAIL.n65 VTAIL.n64 185
R79 VTAIL.n67 VTAIL.n66 185
R80 VTAIL.n12 VTAIL.n11 185
R81 VTAIL.n74 VTAIL.n73 185
R82 VTAIL.n75 VTAIL.n10 185
R83 VTAIL.n77 VTAIL.n76 185
R84 VTAIL.n8 VTAIL.n7 185
R85 VTAIL.n83 VTAIL.n82 185
R86 VTAIL.n85 VTAIL.n84 185
R87 VTAIL.n4 VTAIL.n3 185
R88 VTAIL.n91 VTAIL.n90 185
R89 VTAIL.n93 VTAIL.n92 185
R90 VTAIL.n131 VTAIL.n130 185
R91 VTAIL.n133 VTAIL.n132 185
R92 VTAIL.n126 VTAIL.n125 185
R93 VTAIL.n139 VTAIL.n138 185
R94 VTAIL.n141 VTAIL.n140 185
R95 VTAIL.n122 VTAIL.n121 185
R96 VTAIL.n147 VTAIL.n146 185
R97 VTAIL.n149 VTAIL.n148 185
R98 VTAIL.n118 VTAIL.n117 185
R99 VTAIL.n155 VTAIL.n154 185
R100 VTAIL.n157 VTAIL.n156 185
R101 VTAIL.n114 VTAIL.n113 185
R102 VTAIL.n163 VTAIL.n162 185
R103 VTAIL.n165 VTAIL.n164 185
R104 VTAIL.n110 VTAIL.n109 185
R105 VTAIL.n172 VTAIL.n171 185
R106 VTAIL.n173 VTAIL.n108 185
R107 VTAIL.n175 VTAIL.n174 185
R108 VTAIL.n106 VTAIL.n105 185
R109 VTAIL.n181 VTAIL.n180 185
R110 VTAIL.n183 VTAIL.n182 185
R111 VTAIL.n102 VTAIL.n101 185
R112 VTAIL.n189 VTAIL.n188 185
R113 VTAIL.n191 VTAIL.n190 185
R114 VTAIL.n229 VTAIL.n228 185
R115 VTAIL.n231 VTAIL.n230 185
R116 VTAIL.n224 VTAIL.n223 185
R117 VTAIL.n237 VTAIL.n236 185
R118 VTAIL.n239 VTAIL.n238 185
R119 VTAIL.n220 VTAIL.n219 185
R120 VTAIL.n245 VTAIL.n244 185
R121 VTAIL.n247 VTAIL.n246 185
R122 VTAIL.n216 VTAIL.n215 185
R123 VTAIL.n253 VTAIL.n252 185
R124 VTAIL.n255 VTAIL.n254 185
R125 VTAIL.n212 VTAIL.n211 185
R126 VTAIL.n261 VTAIL.n260 185
R127 VTAIL.n263 VTAIL.n262 185
R128 VTAIL.n208 VTAIL.n207 185
R129 VTAIL.n270 VTAIL.n269 185
R130 VTAIL.n271 VTAIL.n206 185
R131 VTAIL.n273 VTAIL.n272 185
R132 VTAIL.n204 VTAIL.n203 185
R133 VTAIL.n279 VTAIL.n278 185
R134 VTAIL.n281 VTAIL.n280 185
R135 VTAIL.n200 VTAIL.n199 185
R136 VTAIL.n287 VTAIL.n286 185
R137 VTAIL.n289 VTAIL.n288 185
R138 VTAIL.n681 VTAIL.n680 185
R139 VTAIL.n679 VTAIL.n678 185
R140 VTAIL.n592 VTAIL.n591 185
R141 VTAIL.n673 VTAIL.n672 185
R142 VTAIL.n671 VTAIL.n670 185
R143 VTAIL.n596 VTAIL.n595 185
R144 VTAIL.n600 VTAIL.n598 185
R145 VTAIL.n665 VTAIL.n664 185
R146 VTAIL.n663 VTAIL.n662 185
R147 VTAIL.n602 VTAIL.n601 185
R148 VTAIL.n657 VTAIL.n656 185
R149 VTAIL.n655 VTAIL.n654 185
R150 VTAIL.n606 VTAIL.n605 185
R151 VTAIL.n649 VTAIL.n648 185
R152 VTAIL.n647 VTAIL.n646 185
R153 VTAIL.n610 VTAIL.n609 185
R154 VTAIL.n641 VTAIL.n640 185
R155 VTAIL.n639 VTAIL.n638 185
R156 VTAIL.n614 VTAIL.n613 185
R157 VTAIL.n633 VTAIL.n632 185
R158 VTAIL.n631 VTAIL.n630 185
R159 VTAIL.n618 VTAIL.n617 185
R160 VTAIL.n625 VTAIL.n624 185
R161 VTAIL.n623 VTAIL.n622 185
R162 VTAIL.n583 VTAIL.n582 185
R163 VTAIL.n581 VTAIL.n580 185
R164 VTAIL.n494 VTAIL.n493 185
R165 VTAIL.n575 VTAIL.n574 185
R166 VTAIL.n573 VTAIL.n572 185
R167 VTAIL.n498 VTAIL.n497 185
R168 VTAIL.n502 VTAIL.n500 185
R169 VTAIL.n567 VTAIL.n566 185
R170 VTAIL.n565 VTAIL.n564 185
R171 VTAIL.n504 VTAIL.n503 185
R172 VTAIL.n559 VTAIL.n558 185
R173 VTAIL.n557 VTAIL.n556 185
R174 VTAIL.n508 VTAIL.n507 185
R175 VTAIL.n551 VTAIL.n550 185
R176 VTAIL.n549 VTAIL.n548 185
R177 VTAIL.n512 VTAIL.n511 185
R178 VTAIL.n543 VTAIL.n542 185
R179 VTAIL.n541 VTAIL.n540 185
R180 VTAIL.n516 VTAIL.n515 185
R181 VTAIL.n535 VTAIL.n534 185
R182 VTAIL.n533 VTAIL.n532 185
R183 VTAIL.n520 VTAIL.n519 185
R184 VTAIL.n527 VTAIL.n526 185
R185 VTAIL.n525 VTAIL.n524 185
R186 VTAIL.n485 VTAIL.n484 185
R187 VTAIL.n483 VTAIL.n482 185
R188 VTAIL.n396 VTAIL.n395 185
R189 VTAIL.n477 VTAIL.n476 185
R190 VTAIL.n475 VTAIL.n474 185
R191 VTAIL.n400 VTAIL.n399 185
R192 VTAIL.n404 VTAIL.n402 185
R193 VTAIL.n469 VTAIL.n468 185
R194 VTAIL.n467 VTAIL.n466 185
R195 VTAIL.n406 VTAIL.n405 185
R196 VTAIL.n461 VTAIL.n460 185
R197 VTAIL.n459 VTAIL.n458 185
R198 VTAIL.n410 VTAIL.n409 185
R199 VTAIL.n453 VTAIL.n452 185
R200 VTAIL.n451 VTAIL.n450 185
R201 VTAIL.n414 VTAIL.n413 185
R202 VTAIL.n445 VTAIL.n444 185
R203 VTAIL.n443 VTAIL.n442 185
R204 VTAIL.n418 VTAIL.n417 185
R205 VTAIL.n437 VTAIL.n436 185
R206 VTAIL.n435 VTAIL.n434 185
R207 VTAIL.n422 VTAIL.n421 185
R208 VTAIL.n429 VTAIL.n428 185
R209 VTAIL.n427 VTAIL.n426 185
R210 VTAIL.n387 VTAIL.n386 185
R211 VTAIL.n385 VTAIL.n384 185
R212 VTAIL.n298 VTAIL.n297 185
R213 VTAIL.n379 VTAIL.n378 185
R214 VTAIL.n377 VTAIL.n376 185
R215 VTAIL.n302 VTAIL.n301 185
R216 VTAIL.n306 VTAIL.n304 185
R217 VTAIL.n371 VTAIL.n370 185
R218 VTAIL.n369 VTAIL.n368 185
R219 VTAIL.n308 VTAIL.n307 185
R220 VTAIL.n363 VTAIL.n362 185
R221 VTAIL.n361 VTAIL.n360 185
R222 VTAIL.n312 VTAIL.n311 185
R223 VTAIL.n355 VTAIL.n354 185
R224 VTAIL.n353 VTAIL.n352 185
R225 VTAIL.n316 VTAIL.n315 185
R226 VTAIL.n347 VTAIL.n346 185
R227 VTAIL.n345 VTAIL.n344 185
R228 VTAIL.n320 VTAIL.n319 185
R229 VTAIL.n339 VTAIL.n338 185
R230 VTAIL.n337 VTAIL.n336 185
R231 VTAIL.n324 VTAIL.n323 185
R232 VTAIL.n331 VTAIL.n330 185
R233 VTAIL.n329 VTAIL.n328 185
R234 VTAIL.n717 VTAIL.t3 147.659
R235 VTAIL.n31 VTAIL.t2 147.659
R236 VTAIL.n129 VTAIL.t6 147.659
R237 VTAIL.n227 VTAIL.t4 147.659
R238 VTAIL.n621 VTAIL.t7 147.659
R239 VTAIL.n523 VTAIL.t5 147.659
R240 VTAIL.n425 VTAIL.t0 147.659
R241 VTAIL.n327 VTAIL.t1 147.659
R242 VTAIL.n720 VTAIL.n719 104.615
R243 VTAIL.n720 VTAIL.n713 104.615
R244 VTAIL.n727 VTAIL.n713 104.615
R245 VTAIL.n728 VTAIL.n727 104.615
R246 VTAIL.n728 VTAIL.n709 104.615
R247 VTAIL.n735 VTAIL.n709 104.615
R248 VTAIL.n736 VTAIL.n735 104.615
R249 VTAIL.n736 VTAIL.n705 104.615
R250 VTAIL.n743 VTAIL.n705 104.615
R251 VTAIL.n744 VTAIL.n743 104.615
R252 VTAIL.n744 VTAIL.n701 104.615
R253 VTAIL.n751 VTAIL.n701 104.615
R254 VTAIL.n752 VTAIL.n751 104.615
R255 VTAIL.n752 VTAIL.n697 104.615
R256 VTAIL.n760 VTAIL.n697 104.615
R257 VTAIL.n761 VTAIL.n760 104.615
R258 VTAIL.n762 VTAIL.n761 104.615
R259 VTAIL.n762 VTAIL.n693 104.615
R260 VTAIL.n769 VTAIL.n693 104.615
R261 VTAIL.n770 VTAIL.n769 104.615
R262 VTAIL.n770 VTAIL.n689 104.615
R263 VTAIL.n777 VTAIL.n689 104.615
R264 VTAIL.n778 VTAIL.n777 104.615
R265 VTAIL.n34 VTAIL.n33 104.615
R266 VTAIL.n34 VTAIL.n27 104.615
R267 VTAIL.n41 VTAIL.n27 104.615
R268 VTAIL.n42 VTAIL.n41 104.615
R269 VTAIL.n42 VTAIL.n23 104.615
R270 VTAIL.n49 VTAIL.n23 104.615
R271 VTAIL.n50 VTAIL.n49 104.615
R272 VTAIL.n50 VTAIL.n19 104.615
R273 VTAIL.n57 VTAIL.n19 104.615
R274 VTAIL.n58 VTAIL.n57 104.615
R275 VTAIL.n58 VTAIL.n15 104.615
R276 VTAIL.n65 VTAIL.n15 104.615
R277 VTAIL.n66 VTAIL.n65 104.615
R278 VTAIL.n66 VTAIL.n11 104.615
R279 VTAIL.n74 VTAIL.n11 104.615
R280 VTAIL.n75 VTAIL.n74 104.615
R281 VTAIL.n76 VTAIL.n75 104.615
R282 VTAIL.n76 VTAIL.n7 104.615
R283 VTAIL.n83 VTAIL.n7 104.615
R284 VTAIL.n84 VTAIL.n83 104.615
R285 VTAIL.n84 VTAIL.n3 104.615
R286 VTAIL.n91 VTAIL.n3 104.615
R287 VTAIL.n92 VTAIL.n91 104.615
R288 VTAIL.n132 VTAIL.n131 104.615
R289 VTAIL.n132 VTAIL.n125 104.615
R290 VTAIL.n139 VTAIL.n125 104.615
R291 VTAIL.n140 VTAIL.n139 104.615
R292 VTAIL.n140 VTAIL.n121 104.615
R293 VTAIL.n147 VTAIL.n121 104.615
R294 VTAIL.n148 VTAIL.n147 104.615
R295 VTAIL.n148 VTAIL.n117 104.615
R296 VTAIL.n155 VTAIL.n117 104.615
R297 VTAIL.n156 VTAIL.n155 104.615
R298 VTAIL.n156 VTAIL.n113 104.615
R299 VTAIL.n163 VTAIL.n113 104.615
R300 VTAIL.n164 VTAIL.n163 104.615
R301 VTAIL.n164 VTAIL.n109 104.615
R302 VTAIL.n172 VTAIL.n109 104.615
R303 VTAIL.n173 VTAIL.n172 104.615
R304 VTAIL.n174 VTAIL.n173 104.615
R305 VTAIL.n174 VTAIL.n105 104.615
R306 VTAIL.n181 VTAIL.n105 104.615
R307 VTAIL.n182 VTAIL.n181 104.615
R308 VTAIL.n182 VTAIL.n101 104.615
R309 VTAIL.n189 VTAIL.n101 104.615
R310 VTAIL.n190 VTAIL.n189 104.615
R311 VTAIL.n230 VTAIL.n229 104.615
R312 VTAIL.n230 VTAIL.n223 104.615
R313 VTAIL.n237 VTAIL.n223 104.615
R314 VTAIL.n238 VTAIL.n237 104.615
R315 VTAIL.n238 VTAIL.n219 104.615
R316 VTAIL.n245 VTAIL.n219 104.615
R317 VTAIL.n246 VTAIL.n245 104.615
R318 VTAIL.n246 VTAIL.n215 104.615
R319 VTAIL.n253 VTAIL.n215 104.615
R320 VTAIL.n254 VTAIL.n253 104.615
R321 VTAIL.n254 VTAIL.n211 104.615
R322 VTAIL.n261 VTAIL.n211 104.615
R323 VTAIL.n262 VTAIL.n261 104.615
R324 VTAIL.n262 VTAIL.n207 104.615
R325 VTAIL.n270 VTAIL.n207 104.615
R326 VTAIL.n271 VTAIL.n270 104.615
R327 VTAIL.n272 VTAIL.n271 104.615
R328 VTAIL.n272 VTAIL.n203 104.615
R329 VTAIL.n279 VTAIL.n203 104.615
R330 VTAIL.n280 VTAIL.n279 104.615
R331 VTAIL.n280 VTAIL.n199 104.615
R332 VTAIL.n287 VTAIL.n199 104.615
R333 VTAIL.n288 VTAIL.n287 104.615
R334 VTAIL.n680 VTAIL.n679 104.615
R335 VTAIL.n679 VTAIL.n591 104.615
R336 VTAIL.n672 VTAIL.n591 104.615
R337 VTAIL.n672 VTAIL.n671 104.615
R338 VTAIL.n671 VTAIL.n595 104.615
R339 VTAIL.n600 VTAIL.n595 104.615
R340 VTAIL.n664 VTAIL.n600 104.615
R341 VTAIL.n664 VTAIL.n663 104.615
R342 VTAIL.n663 VTAIL.n601 104.615
R343 VTAIL.n656 VTAIL.n601 104.615
R344 VTAIL.n656 VTAIL.n655 104.615
R345 VTAIL.n655 VTAIL.n605 104.615
R346 VTAIL.n648 VTAIL.n605 104.615
R347 VTAIL.n648 VTAIL.n647 104.615
R348 VTAIL.n647 VTAIL.n609 104.615
R349 VTAIL.n640 VTAIL.n609 104.615
R350 VTAIL.n640 VTAIL.n639 104.615
R351 VTAIL.n639 VTAIL.n613 104.615
R352 VTAIL.n632 VTAIL.n613 104.615
R353 VTAIL.n632 VTAIL.n631 104.615
R354 VTAIL.n631 VTAIL.n617 104.615
R355 VTAIL.n624 VTAIL.n617 104.615
R356 VTAIL.n624 VTAIL.n623 104.615
R357 VTAIL.n582 VTAIL.n581 104.615
R358 VTAIL.n581 VTAIL.n493 104.615
R359 VTAIL.n574 VTAIL.n493 104.615
R360 VTAIL.n574 VTAIL.n573 104.615
R361 VTAIL.n573 VTAIL.n497 104.615
R362 VTAIL.n502 VTAIL.n497 104.615
R363 VTAIL.n566 VTAIL.n502 104.615
R364 VTAIL.n566 VTAIL.n565 104.615
R365 VTAIL.n565 VTAIL.n503 104.615
R366 VTAIL.n558 VTAIL.n503 104.615
R367 VTAIL.n558 VTAIL.n557 104.615
R368 VTAIL.n557 VTAIL.n507 104.615
R369 VTAIL.n550 VTAIL.n507 104.615
R370 VTAIL.n550 VTAIL.n549 104.615
R371 VTAIL.n549 VTAIL.n511 104.615
R372 VTAIL.n542 VTAIL.n511 104.615
R373 VTAIL.n542 VTAIL.n541 104.615
R374 VTAIL.n541 VTAIL.n515 104.615
R375 VTAIL.n534 VTAIL.n515 104.615
R376 VTAIL.n534 VTAIL.n533 104.615
R377 VTAIL.n533 VTAIL.n519 104.615
R378 VTAIL.n526 VTAIL.n519 104.615
R379 VTAIL.n526 VTAIL.n525 104.615
R380 VTAIL.n484 VTAIL.n483 104.615
R381 VTAIL.n483 VTAIL.n395 104.615
R382 VTAIL.n476 VTAIL.n395 104.615
R383 VTAIL.n476 VTAIL.n475 104.615
R384 VTAIL.n475 VTAIL.n399 104.615
R385 VTAIL.n404 VTAIL.n399 104.615
R386 VTAIL.n468 VTAIL.n404 104.615
R387 VTAIL.n468 VTAIL.n467 104.615
R388 VTAIL.n467 VTAIL.n405 104.615
R389 VTAIL.n460 VTAIL.n405 104.615
R390 VTAIL.n460 VTAIL.n459 104.615
R391 VTAIL.n459 VTAIL.n409 104.615
R392 VTAIL.n452 VTAIL.n409 104.615
R393 VTAIL.n452 VTAIL.n451 104.615
R394 VTAIL.n451 VTAIL.n413 104.615
R395 VTAIL.n444 VTAIL.n413 104.615
R396 VTAIL.n444 VTAIL.n443 104.615
R397 VTAIL.n443 VTAIL.n417 104.615
R398 VTAIL.n436 VTAIL.n417 104.615
R399 VTAIL.n436 VTAIL.n435 104.615
R400 VTAIL.n435 VTAIL.n421 104.615
R401 VTAIL.n428 VTAIL.n421 104.615
R402 VTAIL.n428 VTAIL.n427 104.615
R403 VTAIL.n386 VTAIL.n385 104.615
R404 VTAIL.n385 VTAIL.n297 104.615
R405 VTAIL.n378 VTAIL.n297 104.615
R406 VTAIL.n378 VTAIL.n377 104.615
R407 VTAIL.n377 VTAIL.n301 104.615
R408 VTAIL.n306 VTAIL.n301 104.615
R409 VTAIL.n370 VTAIL.n306 104.615
R410 VTAIL.n370 VTAIL.n369 104.615
R411 VTAIL.n369 VTAIL.n307 104.615
R412 VTAIL.n362 VTAIL.n307 104.615
R413 VTAIL.n362 VTAIL.n361 104.615
R414 VTAIL.n361 VTAIL.n311 104.615
R415 VTAIL.n354 VTAIL.n311 104.615
R416 VTAIL.n354 VTAIL.n353 104.615
R417 VTAIL.n353 VTAIL.n315 104.615
R418 VTAIL.n346 VTAIL.n315 104.615
R419 VTAIL.n346 VTAIL.n345 104.615
R420 VTAIL.n345 VTAIL.n319 104.615
R421 VTAIL.n338 VTAIL.n319 104.615
R422 VTAIL.n338 VTAIL.n337 104.615
R423 VTAIL.n337 VTAIL.n323 104.615
R424 VTAIL.n330 VTAIL.n323 104.615
R425 VTAIL.n330 VTAIL.n329 104.615
R426 VTAIL.n719 VTAIL.t3 52.3082
R427 VTAIL.n33 VTAIL.t2 52.3082
R428 VTAIL.n131 VTAIL.t6 52.3082
R429 VTAIL.n229 VTAIL.t4 52.3082
R430 VTAIL.n623 VTAIL.t7 52.3082
R431 VTAIL.n525 VTAIL.t5 52.3082
R432 VTAIL.n427 VTAIL.t0 52.3082
R433 VTAIL.n329 VTAIL.t1 52.3082
R434 VTAIL.n783 VTAIL.n782 35.0944
R435 VTAIL.n97 VTAIL.n96 35.0944
R436 VTAIL.n195 VTAIL.n194 35.0944
R437 VTAIL.n293 VTAIL.n292 35.0944
R438 VTAIL.n685 VTAIL.n684 35.0944
R439 VTAIL.n587 VTAIL.n586 35.0944
R440 VTAIL.n489 VTAIL.n488 35.0944
R441 VTAIL.n391 VTAIL.n390 35.0944
R442 VTAIL.n783 VTAIL.n685 31.3324
R443 VTAIL.n391 VTAIL.n293 31.3324
R444 VTAIL.n718 VTAIL.n717 15.6677
R445 VTAIL.n32 VTAIL.n31 15.6677
R446 VTAIL.n130 VTAIL.n129 15.6677
R447 VTAIL.n228 VTAIL.n227 15.6677
R448 VTAIL.n622 VTAIL.n621 15.6677
R449 VTAIL.n524 VTAIL.n523 15.6677
R450 VTAIL.n426 VTAIL.n425 15.6677
R451 VTAIL.n328 VTAIL.n327 15.6677
R452 VTAIL.n763 VTAIL.n694 13.1884
R453 VTAIL.n77 VTAIL.n8 13.1884
R454 VTAIL.n175 VTAIL.n106 13.1884
R455 VTAIL.n273 VTAIL.n204 13.1884
R456 VTAIL.n598 VTAIL.n596 13.1884
R457 VTAIL.n500 VTAIL.n498 13.1884
R458 VTAIL.n402 VTAIL.n400 13.1884
R459 VTAIL.n304 VTAIL.n302 13.1884
R460 VTAIL.n721 VTAIL.n716 12.8005
R461 VTAIL.n764 VTAIL.n696 12.8005
R462 VTAIL.n768 VTAIL.n767 12.8005
R463 VTAIL.n35 VTAIL.n30 12.8005
R464 VTAIL.n78 VTAIL.n10 12.8005
R465 VTAIL.n82 VTAIL.n81 12.8005
R466 VTAIL.n133 VTAIL.n128 12.8005
R467 VTAIL.n176 VTAIL.n108 12.8005
R468 VTAIL.n180 VTAIL.n179 12.8005
R469 VTAIL.n231 VTAIL.n226 12.8005
R470 VTAIL.n274 VTAIL.n206 12.8005
R471 VTAIL.n278 VTAIL.n277 12.8005
R472 VTAIL.n670 VTAIL.n669 12.8005
R473 VTAIL.n666 VTAIL.n665 12.8005
R474 VTAIL.n625 VTAIL.n620 12.8005
R475 VTAIL.n572 VTAIL.n571 12.8005
R476 VTAIL.n568 VTAIL.n567 12.8005
R477 VTAIL.n527 VTAIL.n522 12.8005
R478 VTAIL.n474 VTAIL.n473 12.8005
R479 VTAIL.n470 VTAIL.n469 12.8005
R480 VTAIL.n429 VTAIL.n424 12.8005
R481 VTAIL.n376 VTAIL.n375 12.8005
R482 VTAIL.n372 VTAIL.n371 12.8005
R483 VTAIL.n331 VTAIL.n326 12.8005
R484 VTAIL.n722 VTAIL.n714 12.0247
R485 VTAIL.n759 VTAIL.n758 12.0247
R486 VTAIL.n771 VTAIL.n692 12.0247
R487 VTAIL.n36 VTAIL.n28 12.0247
R488 VTAIL.n73 VTAIL.n72 12.0247
R489 VTAIL.n85 VTAIL.n6 12.0247
R490 VTAIL.n134 VTAIL.n126 12.0247
R491 VTAIL.n171 VTAIL.n170 12.0247
R492 VTAIL.n183 VTAIL.n104 12.0247
R493 VTAIL.n232 VTAIL.n224 12.0247
R494 VTAIL.n269 VTAIL.n268 12.0247
R495 VTAIL.n281 VTAIL.n202 12.0247
R496 VTAIL.n673 VTAIL.n594 12.0247
R497 VTAIL.n662 VTAIL.n599 12.0247
R498 VTAIL.n626 VTAIL.n618 12.0247
R499 VTAIL.n575 VTAIL.n496 12.0247
R500 VTAIL.n564 VTAIL.n501 12.0247
R501 VTAIL.n528 VTAIL.n520 12.0247
R502 VTAIL.n477 VTAIL.n398 12.0247
R503 VTAIL.n466 VTAIL.n403 12.0247
R504 VTAIL.n430 VTAIL.n422 12.0247
R505 VTAIL.n379 VTAIL.n300 12.0247
R506 VTAIL.n368 VTAIL.n305 12.0247
R507 VTAIL.n332 VTAIL.n324 12.0247
R508 VTAIL.n726 VTAIL.n725 11.249
R509 VTAIL.n757 VTAIL.n698 11.249
R510 VTAIL.n772 VTAIL.n690 11.249
R511 VTAIL.n40 VTAIL.n39 11.249
R512 VTAIL.n71 VTAIL.n12 11.249
R513 VTAIL.n86 VTAIL.n4 11.249
R514 VTAIL.n138 VTAIL.n137 11.249
R515 VTAIL.n169 VTAIL.n110 11.249
R516 VTAIL.n184 VTAIL.n102 11.249
R517 VTAIL.n236 VTAIL.n235 11.249
R518 VTAIL.n267 VTAIL.n208 11.249
R519 VTAIL.n282 VTAIL.n200 11.249
R520 VTAIL.n674 VTAIL.n592 11.249
R521 VTAIL.n661 VTAIL.n602 11.249
R522 VTAIL.n630 VTAIL.n629 11.249
R523 VTAIL.n576 VTAIL.n494 11.249
R524 VTAIL.n563 VTAIL.n504 11.249
R525 VTAIL.n532 VTAIL.n531 11.249
R526 VTAIL.n478 VTAIL.n396 11.249
R527 VTAIL.n465 VTAIL.n406 11.249
R528 VTAIL.n434 VTAIL.n433 11.249
R529 VTAIL.n380 VTAIL.n298 11.249
R530 VTAIL.n367 VTAIL.n308 11.249
R531 VTAIL.n336 VTAIL.n335 11.249
R532 VTAIL.n729 VTAIL.n712 10.4732
R533 VTAIL.n754 VTAIL.n753 10.4732
R534 VTAIL.n776 VTAIL.n775 10.4732
R535 VTAIL.n43 VTAIL.n26 10.4732
R536 VTAIL.n68 VTAIL.n67 10.4732
R537 VTAIL.n90 VTAIL.n89 10.4732
R538 VTAIL.n141 VTAIL.n124 10.4732
R539 VTAIL.n166 VTAIL.n165 10.4732
R540 VTAIL.n188 VTAIL.n187 10.4732
R541 VTAIL.n239 VTAIL.n222 10.4732
R542 VTAIL.n264 VTAIL.n263 10.4732
R543 VTAIL.n286 VTAIL.n285 10.4732
R544 VTAIL.n678 VTAIL.n677 10.4732
R545 VTAIL.n658 VTAIL.n657 10.4732
R546 VTAIL.n633 VTAIL.n616 10.4732
R547 VTAIL.n580 VTAIL.n579 10.4732
R548 VTAIL.n560 VTAIL.n559 10.4732
R549 VTAIL.n535 VTAIL.n518 10.4732
R550 VTAIL.n482 VTAIL.n481 10.4732
R551 VTAIL.n462 VTAIL.n461 10.4732
R552 VTAIL.n437 VTAIL.n420 10.4732
R553 VTAIL.n384 VTAIL.n383 10.4732
R554 VTAIL.n364 VTAIL.n363 10.4732
R555 VTAIL.n339 VTAIL.n322 10.4732
R556 VTAIL.n730 VTAIL.n710 9.69747
R557 VTAIL.n750 VTAIL.n700 9.69747
R558 VTAIL.n779 VTAIL.n688 9.69747
R559 VTAIL.n44 VTAIL.n24 9.69747
R560 VTAIL.n64 VTAIL.n14 9.69747
R561 VTAIL.n93 VTAIL.n2 9.69747
R562 VTAIL.n142 VTAIL.n122 9.69747
R563 VTAIL.n162 VTAIL.n112 9.69747
R564 VTAIL.n191 VTAIL.n100 9.69747
R565 VTAIL.n240 VTAIL.n220 9.69747
R566 VTAIL.n260 VTAIL.n210 9.69747
R567 VTAIL.n289 VTAIL.n198 9.69747
R568 VTAIL.n681 VTAIL.n590 9.69747
R569 VTAIL.n654 VTAIL.n604 9.69747
R570 VTAIL.n634 VTAIL.n614 9.69747
R571 VTAIL.n583 VTAIL.n492 9.69747
R572 VTAIL.n556 VTAIL.n506 9.69747
R573 VTAIL.n536 VTAIL.n516 9.69747
R574 VTAIL.n485 VTAIL.n394 9.69747
R575 VTAIL.n458 VTAIL.n408 9.69747
R576 VTAIL.n438 VTAIL.n418 9.69747
R577 VTAIL.n387 VTAIL.n296 9.69747
R578 VTAIL.n360 VTAIL.n310 9.69747
R579 VTAIL.n340 VTAIL.n320 9.69747
R580 VTAIL.n782 VTAIL.n781 9.45567
R581 VTAIL.n96 VTAIL.n95 9.45567
R582 VTAIL.n194 VTAIL.n193 9.45567
R583 VTAIL.n292 VTAIL.n291 9.45567
R584 VTAIL.n684 VTAIL.n683 9.45567
R585 VTAIL.n586 VTAIL.n585 9.45567
R586 VTAIL.n488 VTAIL.n487 9.45567
R587 VTAIL.n390 VTAIL.n389 9.45567
R588 VTAIL.n781 VTAIL.n780 9.3005
R589 VTAIL.n688 VTAIL.n687 9.3005
R590 VTAIL.n775 VTAIL.n774 9.3005
R591 VTAIL.n773 VTAIL.n772 9.3005
R592 VTAIL.n692 VTAIL.n691 9.3005
R593 VTAIL.n767 VTAIL.n766 9.3005
R594 VTAIL.n739 VTAIL.n738 9.3005
R595 VTAIL.n708 VTAIL.n707 9.3005
R596 VTAIL.n733 VTAIL.n732 9.3005
R597 VTAIL.n731 VTAIL.n730 9.3005
R598 VTAIL.n712 VTAIL.n711 9.3005
R599 VTAIL.n725 VTAIL.n724 9.3005
R600 VTAIL.n723 VTAIL.n722 9.3005
R601 VTAIL.n716 VTAIL.n715 9.3005
R602 VTAIL.n741 VTAIL.n740 9.3005
R603 VTAIL.n704 VTAIL.n703 9.3005
R604 VTAIL.n747 VTAIL.n746 9.3005
R605 VTAIL.n749 VTAIL.n748 9.3005
R606 VTAIL.n700 VTAIL.n699 9.3005
R607 VTAIL.n755 VTAIL.n754 9.3005
R608 VTAIL.n757 VTAIL.n756 9.3005
R609 VTAIL.n758 VTAIL.n695 9.3005
R610 VTAIL.n765 VTAIL.n764 9.3005
R611 VTAIL.n95 VTAIL.n94 9.3005
R612 VTAIL.n2 VTAIL.n1 9.3005
R613 VTAIL.n89 VTAIL.n88 9.3005
R614 VTAIL.n87 VTAIL.n86 9.3005
R615 VTAIL.n6 VTAIL.n5 9.3005
R616 VTAIL.n81 VTAIL.n80 9.3005
R617 VTAIL.n53 VTAIL.n52 9.3005
R618 VTAIL.n22 VTAIL.n21 9.3005
R619 VTAIL.n47 VTAIL.n46 9.3005
R620 VTAIL.n45 VTAIL.n44 9.3005
R621 VTAIL.n26 VTAIL.n25 9.3005
R622 VTAIL.n39 VTAIL.n38 9.3005
R623 VTAIL.n37 VTAIL.n36 9.3005
R624 VTAIL.n30 VTAIL.n29 9.3005
R625 VTAIL.n55 VTAIL.n54 9.3005
R626 VTAIL.n18 VTAIL.n17 9.3005
R627 VTAIL.n61 VTAIL.n60 9.3005
R628 VTAIL.n63 VTAIL.n62 9.3005
R629 VTAIL.n14 VTAIL.n13 9.3005
R630 VTAIL.n69 VTAIL.n68 9.3005
R631 VTAIL.n71 VTAIL.n70 9.3005
R632 VTAIL.n72 VTAIL.n9 9.3005
R633 VTAIL.n79 VTAIL.n78 9.3005
R634 VTAIL.n193 VTAIL.n192 9.3005
R635 VTAIL.n100 VTAIL.n99 9.3005
R636 VTAIL.n187 VTAIL.n186 9.3005
R637 VTAIL.n185 VTAIL.n184 9.3005
R638 VTAIL.n104 VTAIL.n103 9.3005
R639 VTAIL.n179 VTAIL.n178 9.3005
R640 VTAIL.n151 VTAIL.n150 9.3005
R641 VTAIL.n120 VTAIL.n119 9.3005
R642 VTAIL.n145 VTAIL.n144 9.3005
R643 VTAIL.n143 VTAIL.n142 9.3005
R644 VTAIL.n124 VTAIL.n123 9.3005
R645 VTAIL.n137 VTAIL.n136 9.3005
R646 VTAIL.n135 VTAIL.n134 9.3005
R647 VTAIL.n128 VTAIL.n127 9.3005
R648 VTAIL.n153 VTAIL.n152 9.3005
R649 VTAIL.n116 VTAIL.n115 9.3005
R650 VTAIL.n159 VTAIL.n158 9.3005
R651 VTAIL.n161 VTAIL.n160 9.3005
R652 VTAIL.n112 VTAIL.n111 9.3005
R653 VTAIL.n167 VTAIL.n166 9.3005
R654 VTAIL.n169 VTAIL.n168 9.3005
R655 VTAIL.n170 VTAIL.n107 9.3005
R656 VTAIL.n177 VTAIL.n176 9.3005
R657 VTAIL.n291 VTAIL.n290 9.3005
R658 VTAIL.n198 VTAIL.n197 9.3005
R659 VTAIL.n285 VTAIL.n284 9.3005
R660 VTAIL.n283 VTAIL.n282 9.3005
R661 VTAIL.n202 VTAIL.n201 9.3005
R662 VTAIL.n277 VTAIL.n276 9.3005
R663 VTAIL.n249 VTAIL.n248 9.3005
R664 VTAIL.n218 VTAIL.n217 9.3005
R665 VTAIL.n243 VTAIL.n242 9.3005
R666 VTAIL.n241 VTAIL.n240 9.3005
R667 VTAIL.n222 VTAIL.n221 9.3005
R668 VTAIL.n235 VTAIL.n234 9.3005
R669 VTAIL.n233 VTAIL.n232 9.3005
R670 VTAIL.n226 VTAIL.n225 9.3005
R671 VTAIL.n251 VTAIL.n250 9.3005
R672 VTAIL.n214 VTAIL.n213 9.3005
R673 VTAIL.n257 VTAIL.n256 9.3005
R674 VTAIL.n259 VTAIL.n258 9.3005
R675 VTAIL.n210 VTAIL.n209 9.3005
R676 VTAIL.n265 VTAIL.n264 9.3005
R677 VTAIL.n267 VTAIL.n266 9.3005
R678 VTAIL.n268 VTAIL.n205 9.3005
R679 VTAIL.n275 VTAIL.n274 9.3005
R680 VTAIL.n608 VTAIL.n607 9.3005
R681 VTAIL.n651 VTAIL.n650 9.3005
R682 VTAIL.n653 VTAIL.n652 9.3005
R683 VTAIL.n604 VTAIL.n603 9.3005
R684 VTAIL.n659 VTAIL.n658 9.3005
R685 VTAIL.n661 VTAIL.n660 9.3005
R686 VTAIL.n599 VTAIL.n597 9.3005
R687 VTAIL.n667 VTAIL.n666 9.3005
R688 VTAIL.n683 VTAIL.n682 9.3005
R689 VTAIL.n590 VTAIL.n589 9.3005
R690 VTAIL.n677 VTAIL.n676 9.3005
R691 VTAIL.n675 VTAIL.n674 9.3005
R692 VTAIL.n594 VTAIL.n593 9.3005
R693 VTAIL.n669 VTAIL.n668 9.3005
R694 VTAIL.n645 VTAIL.n644 9.3005
R695 VTAIL.n643 VTAIL.n642 9.3005
R696 VTAIL.n612 VTAIL.n611 9.3005
R697 VTAIL.n637 VTAIL.n636 9.3005
R698 VTAIL.n635 VTAIL.n634 9.3005
R699 VTAIL.n616 VTAIL.n615 9.3005
R700 VTAIL.n629 VTAIL.n628 9.3005
R701 VTAIL.n627 VTAIL.n626 9.3005
R702 VTAIL.n620 VTAIL.n619 9.3005
R703 VTAIL.n510 VTAIL.n509 9.3005
R704 VTAIL.n553 VTAIL.n552 9.3005
R705 VTAIL.n555 VTAIL.n554 9.3005
R706 VTAIL.n506 VTAIL.n505 9.3005
R707 VTAIL.n561 VTAIL.n560 9.3005
R708 VTAIL.n563 VTAIL.n562 9.3005
R709 VTAIL.n501 VTAIL.n499 9.3005
R710 VTAIL.n569 VTAIL.n568 9.3005
R711 VTAIL.n585 VTAIL.n584 9.3005
R712 VTAIL.n492 VTAIL.n491 9.3005
R713 VTAIL.n579 VTAIL.n578 9.3005
R714 VTAIL.n577 VTAIL.n576 9.3005
R715 VTAIL.n496 VTAIL.n495 9.3005
R716 VTAIL.n571 VTAIL.n570 9.3005
R717 VTAIL.n547 VTAIL.n546 9.3005
R718 VTAIL.n545 VTAIL.n544 9.3005
R719 VTAIL.n514 VTAIL.n513 9.3005
R720 VTAIL.n539 VTAIL.n538 9.3005
R721 VTAIL.n537 VTAIL.n536 9.3005
R722 VTAIL.n518 VTAIL.n517 9.3005
R723 VTAIL.n531 VTAIL.n530 9.3005
R724 VTAIL.n529 VTAIL.n528 9.3005
R725 VTAIL.n522 VTAIL.n521 9.3005
R726 VTAIL.n412 VTAIL.n411 9.3005
R727 VTAIL.n455 VTAIL.n454 9.3005
R728 VTAIL.n457 VTAIL.n456 9.3005
R729 VTAIL.n408 VTAIL.n407 9.3005
R730 VTAIL.n463 VTAIL.n462 9.3005
R731 VTAIL.n465 VTAIL.n464 9.3005
R732 VTAIL.n403 VTAIL.n401 9.3005
R733 VTAIL.n471 VTAIL.n470 9.3005
R734 VTAIL.n487 VTAIL.n486 9.3005
R735 VTAIL.n394 VTAIL.n393 9.3005
R736 VTAIL.n481 VTAIL.n480 9.3005
R737 VTAIL.n479 VTAIL.n478 9.3005
R738 VTAIL.n398 VTAIL.n397 9.3005
R739 VTAIL.n473 VTAIL.n472 9.3005
R740 VTAIL.n449 VTAIL.n448 9.3005
R741 VTAIL.n447 VTAIL.n446 9.3005
R742 VTAIL.n416 VTAIL.n415 9.3005
R743 VTAIL.n441 VTAIL.n440 9.3005
R744 VTAIL.n439 VTAIL.n438 9.3005
R745 VTAIL.n420 VTAIL.n419 9.3005
R746 VTAIL.n433 VTAIL.n432 9.3005
R747 VTAIL.n431 VTAIL.n430 9.3005
R748 VTAIL.n424 VTAIL.n423 9.3005
R749 VTAIL.n314 VTAIL.n313 9.3005
R750 VTAIL.n357 VTAIL.n356 9.3005
R751 VTAIL.n359 VTAIL.n358 9.3005
R752 VTAIL.n310 VTAIL.n309 9.3005
R753 VTAIL.n365 VTAIL.n364 9.3005
R754 VTAIL.n367 VTAIL.n366 9.3005
R755 VTAIL.n305 VTAIL.n303 9.3005
R756 VTAIL.n373 VTAIL.n372 9.3005
R757 VTAIL.n389 VTAIL.n388 9.3005
R758 VTAIL.n296 VTAIL.n295 9.3005
R759 VTAIL.n383 VTAIL.n382 9.3005
R760 VTAIL.n381 VTAIL.n380 9.3005
R761 VTAIL.n300 VTAIL.n299 9.3005
R762 VTAIL.n375 VTAIL.n374 9.3005
R763 VTAIL.n351 VTAIL.n350 9.3005
R764 VTAIL.n349 VTAIL.n348 9.3005
R765 VTAIL.n318 VTAIL.n317 9.3005
R766 VTAIL.n343 VTAIL.n342 9.3005
R767 VTAIL.n341 VTAIL.n340 9.3005
R768 VTAIL.n322 VTAIL.n321 9.3005
R769 VTAIL.n335 VTAIL.n334 9.3005
R770 VTAIL.n333 VTAIL.n332 9.3005
R771 VTAIL.n326 VTAIL.n325 9.3005
R772 VTAIL.n734 VTAIL.n733 8.92171
R773 VTAIL.n749 VTAIL.n702 8.92171
R774 VTAIL.n780 VTAIL.n686 8.92171
R775 VTAIL.n48 VTAIL.n47 8.92171
R776 VTAIL.n63 VTAIL.n16 8.92171
R777 VTAIL.n94 VTAIL.n0 8.92171
R778 VTAIL.n146 VTAIL.n145 8.92171
R779 VTAIL.n161 VTAIL.n114 8.92171
R780 VTAIL.n192 VTAIL.n98 8.92171
R781 VTAIL.n244 VTAIL.n243 8.92171
R782 VTAIL.n259 VTAIL.n212 8.92171
R783 VTAIL.n290 VTAIL.n196 8.92171
R784 VTAIL.n682 VTAIL.n588 8.92171
R785 VTAIL.n653 VTAIL.n606 8.92171
R786 VTAIL.n638 VTAIL.n637 8.92171
R787 VTAIL.n584 VTAIL.n490 8.92171
R788 VTAIL.n555 VTAIL.n508 8.92171
R789 VTAIL.n540 VTAIL.n539 8.92171
R790 VTAIL.n486 VTAIL.n392 8.92171
R791 VTAIL.n457 VTAIL.n410 8.92171
R792 VTAIL.n442 VTAIL.n441 8.92171
R793 VTAIL.n388 VTAIL.n294 8.92171
R794 VTAIL.n359 VTAIL.n312 8.92171
R795 VTAIL.n344 VTAIL.n343 8.92171
R796 VTAIL.n737 VTAIL.n708 8.14595
R797 VTAIL.n746 VTAIL.n745 8.14595
R798 VTAIL.n51 VTAIL.n22 8.14595
R799 VTAIL.n60 VTAIL.n59 8.14595
R800 VTAIL.n149 VTAIL.n120 8.14595
R801 VTAIL.n158 VTAIL.n157 8.14595
R802 VTAIL.n247 VTAIL.n218 8.14595
R803 VTAIL.n256 VTAIL.n255 8.14595
R804 VTAIL.n650 VTAIL.n649 8.14595
R805 VTAIL.n641 VTAIL.n612 8.14595
R806 VTAIL.n552 VTAIL.n551 8.14595
R807 VTAIL.n543 VTAIL.n514 8.14595
R808 VTAIL.n454 VTAIL.n453 8.14595
R809 VTAIL.n445 VTAIL.n416 8.14595
R810 VTAIL.n356 VTAIL.n355 8.14595
R811 VTAIL.n347 VTAIL.n318 8.14595
R812 VTAIL.n738 VTAIL.n706 7.3702
R813 VTAIL.n742 VTAIL.n704 7.3702
R814 VTAIL.n52 VTAIL.n20 7.3702
R815 VTAIL.n56 VTAIL.n18 7.3702
R816 VTAIL.n150 VTAIL.n118 7.3702
R817 VTAIL.n154 VTAIL.n116 7.3702
R818 VTAIL.n248 VTAIL.n216 7.3702
R819 VTAIL.n252 VTAIL.n214 7.3702
R820 VTAIL.n646 VTAIL.n608 7.3702
R821 VTAIL.n642 VTAIL.n610 7.3702
R822 VTAIL.n548 VTAIL.n510 7.3702
R823 VTAIL.n544 VTAIL.n512 7.3702
R824 VTAIL.n450 VTAIL.n412 7.3702
R825 VTAIL.n446 VTAIL.n414 7.3702
R826 VTAIL.n352 VTAIL.n314 7.3702
R827 VTAIL.n348 VTAIL.n316 7.3702
R828 VTAIL.n741 VTAIL.n706 6.59444
R829 VTAIL.n742 VTAIL.n741 6.59444
R830 VTAIL.n55 VTAIL.n20 6.59444
R831 VTAIL.n56 VTAIL.n55 6.59444
R832 VTAIL.n153 VTAIL.n118 6.59444
R833 VTAIL.n154 VTAIL.n153 6.59444
R834 VTAIL.n251 VTAIL.n216 6.59444
R835 VTAIL.n252 VTAIL.n251 6.59444
R836 VTAIL.n646 VTAIL.n645 6.59444
R837 VTAIL.n645 VTAIL.n610 6.59444
R838 VTAIL.n548 VTAIL.n547 6.59444
R839 VTAIL.n547 VTAIL.n512 6.59444
R840 VTAIL.n450 VTAIL.n449 6.59444
R841 VTAIL.n449 VTAIL.n414 6.59444
R842 VTAIL.n352 VTAIL.n351 6.59444
R843 VTAIL.n351 VTAIL.n316 6.59444
R844 VTAIL.n738 VTAIL.n737 5.81868
R845 VTAIL.n745 VTAIL.n704 5.81868
R846 VTAIL.n52 VTAIL.n51 5.81868
R847 VTAIL.n59 VTAIL.n18 5.81868
R848 VTAIL.n150 VTAIL.n149 5.81868
R849 VTAIL.n157 VTAIL.n116 5.81868
R850 VTAIL.n248 VTAIL.n247 5.81868
R851 VTAIL.n255 VTAIL.n214 5.81868
R852 VTAIL.n649 VTAIL.n608 5.81868
R853 VTAIL.n642 VTAIL.n641 5.81868
R854 VTAIL.n551 VTAIL.n510 5.81868
R855 VTAIL.n544 VTAIL.n543 5.81868
R856 VTAIL.n453 VTAIL.n412 5.81868
R857 VTAIL.n446 VTAIL.n445 5.81868
R858 VTAIL.n355 VTAIL.n314 5.81868
R859 VTAIL.n348 VTAIL.n347 5.81868
R860 VTAIL.n734 VTAIL.n708 5.04292
R861 VTAIL.n746 VTAIL.n702 5.04292
R862 VTAIL.n782 VTAIL.n686 5.04292
R863 VTAIL.n48 VTAIL.n22 5.04292
R864 VTAIL.n60 VTAIL.n16 5.04292
R865 VTAIL.n96 VTAIL.n0 5.04292
R866 VTAIL.n146 VTAIL.n120 5.04292
R867 VTAIL.n158 VTAIL.n114 5.04292
R868 VTAIL.n194 VTAIL.n98 5.04292
R869 VTAIL.n244 VTAIL.n218 5.04292
R870 VTAIL.n256 VTAIL.n212 5.04292
R871 VTAIL.n292 VTAIL.n196 5.04292
R872 VTAIL.n684 VTAIL.n588 5.04292
R873 VTAIL.n650 VTAIL.n606 5.04292
R874 VTAIL.n638 VTAIL.n612 5.04292
R875 VTAIL.n586 VTAIL.n490 5.04292
R876 VTAIL.n552 VTAIL.n508 5.04292
R877 VTAIL.n540 VTAIL.n514 5.04292
R878 VTAIL.n488 VTAIL.n392 5.04292
R879 VTAIL.n454 VTAIL.n410 5.04292
R880 VTAIL.n442 VTAIL.n416 5.04292
R881 VTAIL.n390 VTAIL.n294 5.04292
R882 VTAIL.n356 VTAIL.n312 5.04292
R883 VTAIL.n344 VTAIL.n318 5.04292
R884 VTAIL.n717 VTAIL.n715 4.38563
R885 VTAIL.n31 VTAIL.n29 4.38563
R886 VTAIL.n129 VTAIL.n127 4.38563
R887 VTAIL.n227 VTAIL.n225 4.38563
R888 VTAIL.n621 VTAIL.n619 4.38563
R889 VTAIL.n523 VTAIL.n521 4.38563
R890 VTAIL.n425 VTAIL.n423 4.38563
R891 VTAIL.n327 VTAIL.n325 4.38563
R892 VTAIL.n733 VTAIL.n710 4.26717
R893 VTAIL.n750 VTAIL.n749 4.26717
R894 VTAIL.n780 VTAIL.n779 4.26717
R895 VTAIL.n47 VTAIL.n24 4.26717
R896 VTAIL.n64 VTAIL.n63 4.26717
R897 VTAIL.n94 VTAIL.n93 4.26717
R898 VTAIL.n145 VTAIL.n122 4.26717
R899 VTAIL.n162 VTAIL.n161 4.26717
R900 VTAIL.n192 VTAIL.n191 4.26717
R901 VTAIL.n243 VTAIL.n220 4.26717
R902 VTAIL.n260 VTAIL.n259 4.26717
R903 VTAIL.n290 VTAIL.n289 4.26717
R904 VTAIL.n682 VTAIL.n681 4.26717
R905 VTAIL.n654 VTAIL.n653 4.26717
R906 VTAIL.n637 VTAIL.n614 4.26717
R907 VTAIL.n584 VTAIL.n583 4.26717
R908 VTAIL.n556 VTAIL.n555 4.26717
R909 VTAIL.n539 VTAIL.n516 4.26717
R910 VTAIL.n486 VTAIL.n485 4.26717
R911 VTAIL.n458 VTAIL.n457 4.26717
R912 VTAIL.n441 VTAIL.n418 4.26717
R913 VTAIL.n388 VTAIL.n387 4.26717
R914 VTAIL.n360 VTAIL.n359 4.26717
R915 VTAIL.n343 VTAIL.n320 4.26717
R916 VTAIL.n489 VTAIL.n391 3.73326
R917 VTAIL.n685 VTAIL.n587 3.73326
R918 VTAIL.n293 VTAIL.n195 3.73326
R919 VTAIL.n730 VTAIL.n729 3.49141
R920 VTAIL.n753 VTAIL.n700 3.49141
R921 VTAIL.n776 VTAIL.n688 3.49141
R922 VTAIL.n44 VTAIL.n43 3.49141
R923 VTAIL.n67 VTAIL.n14 3.49141
R924 VTAIL.n90 VTAIL.n2 3.49141
R925 VTAIL.n142 VTAIL.n141 3.49141
R926 VTAIL.n165 VTAIL.n112 3.49141
R927 VTAIL.n188 VTAIL.n100 3.49141
R928 VTAIL.n240 VTAIL.n239 3.49141
R929 VTAIL.n263 VTAIL.n210 3.49141
R930 VTAIL.n286 VTAIL.n198 3.49141
R931 VTAIL.n678 VTAIL.n590 3.49141
R932 VTAIL.n657 VTAIL.n604 3.49141
R933 VTAIL.n634 VTAIL.n633 3.49141
R934 VTAIL.n580 VTAIL.n492 3.49141
R935 VTAIL.n559 VTAIL.n506 3.49141
R936 VTAIL.n536 VTAIL.n535 3.49141
R937 VTAIL.n482 VTAIL.n394 3.49141
R938 VTAIL.n461 VTAIL.n408 3.49141
R939 VTAIL.n438 VTAIL.n437 3.49141
R940 VTAIL.n384 VTAIL.n296 3.49141
R941 VTAIL.n363 VTAIL.n310 3.49141
R942 VTAIL.n340 VTAIL.n339 3.49141
R943 VTAIL.n726 VTAIL.n712 2.71565
R944 VTAIL.n754 VTAIL.n698 2.71565
R945 VTAIL.n775 VTAIL.n690 2.71565
R946 VTAIL.n40 VTAIL.n26 2.71565
R947 VTAIL.n68 VTAIL.n12 2.71565
R948 VTAIL.n89 VTAIL.n4 2.71565
R949 VTAIL.n138 VTAIL.n124 2.71565
R950 VTAIL.n166 VTAIL.n110 2.71565
R951 VTAIL.n187 VTAIL.n102 2.71565
R952 VTAIL.n236 VTAIL.n222 2.71565
R953 VTAIL.n264 VTAIL.n208 2.71565
R954 VTAIL.n285 VTAIL.n200 2.71565
R955 VTAIL.n677 VTAIL.n592 2.71565
R956 VTAIL.n658 VTAIL.n602 2.71565
R957 VTAIL.n630 VTAIL.n616 2.71565
R958 VTAIL.n579 VTAIL.n494 2.71565
R959 VTAIL.n560 VTAIL.n504 2.71565
R960 VTAIL.n532 VTAIL.n518 2.71565
R961 VTAIL.n481 VTAIL.n396 2.71565
R962 VTAIL.n462 VTAIL.n406 2.71565
R963 VTAIL.n434 VTAIL.n420 2.71565
R964 VTAIL.n383 VTAIL.n298 2.71565
R965 VTAIL.n364 VTAIL.n308 2.71565
R966 VTAIL.n336 VTAIL.n322 2.71565
R967 VTAIL.n725 VTAIL.n714 1.93989
R968 VTAIL.n759 VTAIL.n757 1.93989
R969 VTAIL.n772 VTAIL.n771 1.93989
R970 VTAIL.n39 VTAIL.n28 1.93989
R971 VTAIL.n73 VTAIL.n71 1.93989
R972 VTAIL.n86 VTAIL.n85 1.93989
R973 VTAIL.n137 VTAIL.n126 1.93989
R974 VTAIL.n171 VTAIL.n169 1.93989
R975 VTAIL.n184 VTAIL.n183 1.93989
R976 VTAIL.n235 VTAIL.n224 1.93989
R977 VTAIL.n269 VTAIL.n267 1.93989
R978 VTAIL.n282 VTAIL.n281 1.93989
R979 VTAIL.n674 VTAIL.n673 1.93989
R980 VTAIL.n662 VTAIL.n661 1.93989
R981 VTAIL.n629 VTAIL.n618 1.93989
R982 VTAIL.n576 VTAIL.n575 1.93989
R983 VTAIL.n564 VTAIL.n563 1.93989
R984 VTAIL.n531 VTAIL.n520 1.93989
R985 VTAIL.n478 VTAIL.n477 1.93989
R986 VTAIL.n466 VTAIL.n465 1.93989
R987 VTAIL.n433 VTAIL.n422 1.93989
R988 VTAIL.n380 VTAIL.n379 1.93989
R989 VTAIL.n368 VTAIL.n367 1.93989
R990 VTAIL.n335 VTAIL.n324 1.93989
R991 VTAIL VTAIL.n97 1.92507
R992 VTAIL VTAIL.n783 1.80869
R993 VTAIL.n722 VTAIL.n721 1.16414
R994 VTAIL.n758 VTAIL.n696 1.16414
R995 VTAIL.n768 VTAIL.n692 1.16414
R996 VTAIL.n36 VTAIL.n35 1.16414
R997 VTAIL.n72 VTAIL.n10 1.16414
R998 VTAIL.n82 VTAIL.n6 1.16414
R999 VTAIL.n134 VTAIL.n133 1.16414
R1000 VTAIL.n170 VTAIL.n108 1.16414
R1001 VTAIL.n180 VTAIL.n104 1.16414
R1002 VTAIL.n232 VTAIL.n231 1.16414
R1003 VTAIL.n268 VTAIL.n206 1.16414
R1004 VTAIL.n278 VTAIL.n202 1.16414
R1005 VTAIL.n670 VTAIL.n594 1.16414
R1006 VTAIL.n665 VTAIL.n599 1.16414
R1007 VTAIL.n626 VTAIL.n625 1.16414
R1008 VTAIL.n572 VTAIL.n496 1.16414
R1009 VTAIL.n567 VTAIL.n501 1.16414
R1010 VTAIL.n528 VTAIL.n527 1.16414
R1011 VTAIL.n474 VTAIL.n398 1.16414
R1012 VTAIL.n469 VTAIL.n403 1.16414
R1013 VTAIL.n430 VTAIL.n429 1.16414
R1014 VTAIL.n376 VTAIL.n300 1.16414
R1015 VTAIL.n371 VTAIL.n305 1.16414
R1016 VTAIL.n332 VTAIL.n331 1.16414
R1017 VTAIL.n587 VTAIL.n489 0.470328
R1018 VTAIL.n195 VTAIL.n97 0.470328
R1019 VTAIL.n718 VTAIL.n716 0.388379
R1020 VTAIL.n764 VTAIL.n763 0.388379
R1021 VTAIL.n767 VTAIL.n694 0.388379
R1022 VTAIL.n32 VTAIL.n30 0.388379
R1023 VTAIL.n78 VTAIL.n77 0.388379
R1024 VTAIL.n81 VTAIL.n8 0.388379
R1025 VTAIL.n130 VTAIL.n128 0.388379
R1026 VTAIL.n176 VTAIL.n175 0.388379
R1027 VTAIL.n179 VTAIL.n106 0.388379
R1028 VTAIL.n228 VTAIL.n226 0.388379
R1029 VTAIL.n274 VTAIL.n273 0.388379
R1030 VTAIL.n277 VTAIL.n204 0.388379
R1031 VTAIL.n669 VTAIL.n596 0.388379
R1032 VTAIL.n666 VTAIL.n598 0.388379
R1033 VTAIL.n622 VTAIL.n620 0.388379
R1034 VTAIL.n571 VTAIL.n498 0.388379
R1035 VTAIL.n568 VTAIL.n500 0.388379
R1036 VTAIL.n524 VTAIL.n522 0.388379
R1037 VTAIL.n473 VTAIL.n400 0.388379
R1038 VTAIL.n470 VTAIL.n402 0.388379
R1039 VTAIL.n426 VTAIL.n424 0.388379
R1040 VTAIL.n375 VTAIL.n302 0.388379
R1041 VTAIL.n372 VTAIL.n304 0.388379
R1042 VTAIL.n328 VTAIL.n326 0.388379
R1043 VTAIL.n723 VTAIL.n715 0.155672
R1044 VTAIL.n724 VTAIL.n723 0.155672
R1045 VTAIL.n724 VTAIL.n711 0.155672
R1046 VTAIL.n731 VTAIL.n711 0.155672
R1047 VTAIL.n732 VTAIL.n731 0.155672
R1048 VTAIL.n732 VTAIL.n707 0.155672
R1049 VTAIL.n739 VTAIL.n707 0.155672
R1050 VTAIL.n740 VTAIL.n739 0.155672
R1051 VTAIL.n740 VTAIL.n703 0.155672
R1052 VTAIL.n747 VTAIL.n703 0.155672
R1053 VTAIL.n748 VTAIL.n747 0.155672
R1054 VTAIL.n748 VTAIL.n699 0.155672
R1055 VTAIL.n755 VTAIL.n699 0.155672
R1056 VTAIL.n756 VTAIL.n755 0.155672
R1057 VTAIL.n756 VTAIL.n695 0.155672
R1058 VTAIL.n765 VTAIL.n695 0.155672
R1059 VTAIL.n766 VTAIL.n765 0.155672
R1060 VTAIL.n766 VTAIL.n691 0.155672
R1061 VTAIL.n773 VTAIL.n691 0.155672
R1062 VTAIL.n774 VTAIL.n773 0.155672
R1063 VTAIL.n774 VTAIL.n687 0.155672
R1064 VTAIL.n781 VTAIL.n687 0.155672
R1065 VTAIL.n37 VTAIL.n29 0.155672
R1066 VTAIL.n38 VTAIL.n37 0.155672
R1067 VTAIL.n38 VTAIL.n25 0.155672
R1068 VTAIL.n45 VTAIL.n25 0.155672
R1069 VTAIL.n46 VTAIL.n45 0.155672
R1070 VTAIL.n46 VTAIL.n21 0.155672
R1071 VTAIL.n53 VTAIL.n21 0.155672
R1072 VTAIL.n54 VTAIL.n53 0.155672
R1073 VTAIL.n54 VTAIL.n17 0.155672
R1074 VTAIL.n61 VTAIL.n17 0.155672
R1075 VTAIL.n62 VTAIL.n61 0.155672
R1076 VTAIL.n62 VTAIL.n13 0.155672
R1077 VTAIL.n69 VTAIL.n13 0.155672
R1078 VTAIL.n70 VTAIL.n69 0.155672
R1079 VTAIL.n70 VTAIL.n9 0.155672
R1080 VTAIL.n79 VTAIL.n9 0.155672
R1081 VTAIL.n80 VTAIL.n79 0.155672
R1082 VTAIL.n80 VTAIL.n5 0.155672
R1083 VTAIL.n87 VTAIL.n5 0.155672
R1084 VTAIL.n88 VTAIL.n87 0.155672
R1085 VTAIL.n88 VTAIL.n1 0.155672
R1086 VTAIL.n95 VTAIL.n1 0.155672
R1087 VTAIL.n135 VTAIL.n127 0.155672
R1088 VTAIL.n136 VTAIL.n135 0.155672
R1089 VTAIL.n136 VTAIL.n123 0.155672
R1090 VTAIL.n143 VTAIL.n123 0.155672
R1091 VTAIL.n144 VTAIL.n143 0.155672
R1092 VTAIL.n144 VTAIL.n119 0.155672
R1093 VTAIL.n151 VTAIL.n119 0.155672
R1094 VTAIL.n152 VTAIL.n151 0.155672
R1095 VTAIL.n152 VTAIL.n115 0.155672
R1096 VTAIL.n159 VTAIL.n115 0.155672
R1097 VTAIL.n160 VTAIL.n159 0.155672
R1098 VTAIL.n160 VTAIL.n111 0.155672
R1099 VTAIL.n167 VTAIL.n111 0.155672
R1100 VTAIL.n168 VTAIL.n167 0.155672
R1101 VTAIL.n168 VTAIL.n107 0.155672
R1102 VTAIL.n177 VTAIL.n107 0.155672
R1103 VTAIL.n178 VTAIL.n177 0.155672
R1104 VTAIL.n178 VTAIL.n103 0.155672
R1105 VTAIL.n185 VTAIL.n103 0.155672
R1106 VTAIL.n186 VTAIL.n185 0.155672
R1107 VTAIL.n186 VTAIL.n99 0.155672
R1108 VTAIL.n193 VTAIL.n99 0.155672
R1109 VTAIL.n233 VTAIL.n225 0.155672
R1110 VTAIL.n234 VTAIL.n233 0.155672
R1111 VTAIL.n234 VTAIL.n221 0.155672
R1112 VTAIL.n241 VTAIL.n221 0.155672
R1113 VTAIL.n242 VTAIL.n241 0.155672
R1114 VTAIL.n242 VTAIL.n217 0.155672
R1115 VTAIL.n249 VTAIL.n217 0.155672
R1116 VTAIL.n250 VTAIL.n249 0.155672
R1117 VTAIL.n250 VTAIL.n213 0.155672
R1118 VTAIL.n257 VTAIL.n213 0.155672
R1119 VTAIL.n258 VTAIL.n257 0.155672
R1120 VTAIL.n258 VTAIL.n209 0.155672
R1121 VTAIL.n265 VTAIL.n209 0.155672
R1122 VTAIL.n266 VTAIL.n265 0.155672
R1123 VTAIL.n266 VTAIL.n205 0.155672
R1124 VTAIL.n275 VTAIL.n205 0.155672
R1125 VTAIL.n276 VTAIL.n275 0.155672
R1126 VTAIL.n276 VTAIL.n201 0.155672
R1127 VTAIL.n283 VTAIL.n201 0.155672
R1128 VTAIL.n284 VTAIL.n283 0.155672
R1129 VTAIL.n284 VTAIL.n197 0.155672
R1130 VTAIL.n291 VTAIL.n197 0.155672
R1131 VTAIL.n683 VTAIL.n589 0.155672
R1132 VTAIL.n676 VTAIL.n589 0.155672
R1133 VTAIL.n676 VTAIL.n675 0.155672
R1134 VTAIL.n675 VTAIL.n593 0.155672
R1135 VTAIL.n668 VTAIL.n593 0.155672
R1136 VTAIL.n668 VTAIL.n667 0.155672
R1137 VTAIL.n667 VTAIL.n597 0.155672
R1138 VTAIL.n660 VTAIL.n597 0.155672
R1139 VTAIL.n660 VTAIL.n659 0.155672
R1140 VTAIL.n659 VTAIL.n603 0.155672
R1141 VTAIL.n652 VTAIL.n603 0.155672
R1142 VTAIL.n652 VTAIL.n651 0.155672
R1143 VTAIL.n651 VTAIL.n607 0.155672
R1144 VTAIL.n644 VTAIL.n607 0.155672
R1145 VTAIL.n644 VTAIL.n643 0.155672
R1146 VTAIL.n643 VTAIL.n611 0.155672
R1147 VTAIL.n636 VTAIL.n611 0.155672
R1148 VTAIL.n636 VTAIL.n635 0.155672
R1149 VTAIL.n635 VTAIL.n615 0.155672
R1150 VTAIL.n628 VTAIL.n615 0.155672
R1151 VTAIL.n628 VTAIL.n627 0.155672
R1152 VTAIL.n627 VTAIL.n619 0.155672
R1153 VTAIL.n585 VTAIL.n491 0.155672
R1154 VTAIL.n578 VTAIL.n491 0.155672
R1155 VTAIL.n578 VTAIL.n577 0.155672
R1156 VTAIL.n577 VTAIL.n495 0.155672
R1157 VTAIL.n570 VTAIL.n495 0.155672
R1158 VTAIL.n570 VTAIL.n569 0.155672
R1159 VTAIL.n569 VTAIL.n499 0.155672
R1160 VTAIL.n562 VTAIL.n499 0.155672
R1161 VTAIL.n562 VTAIL.n561 0.155672
R1162 VTAIL.n561 VTAIL.n505 0.155672
R1163 VTAIL.n554 VTAIL.n505 0.155672
R1164 VTAIL.n554 VTAIL.n553 0.155672
R1165 VTAIL.n553 VTAIL.n509 0.155672
R1166 VTAIL.n546 VTAIL.n509 0.155672
R1167 VTAIL.n546 VTAIL.n545 0.155672
R1168 VTAIL.n545 VTAIL.n513 0.155672
R1169 VTAIL.n538 VTAIL.n513 0.155672
R1170 VTAIL.n538 VTAIL.n537 0.155672
R1171 VTAIL.n537 VTAIL.n517 0.155672
R1172 VTAIL.n530 VTAIL.n517 0.155672
R1173 VTAIL.n530 VTAIL.n529 0.155672
R1174 VTAIL.n529 VTAIL.n521 0.155672
R1175 VTAIL.n487 VTAIL.n393 0.155672
R1176 VTAIL.n480 VTAIL.n393 0.155672
R1177 VTAIL.n480 VTAIL.n479 0.155672
R1178 VTAIL.n479 VTAIL.n397 0.155672
R1179 VTAIL.n472 VTAIL.n397 0.155672
R1180 VTAIL.n472 VTAIL.n471 0.155672
R1181 VTAIL.n471 VTAIL.n401 0.155672
R1182 VTAIL.n464 VTAIL.n401 0.155672
R1183 VTAIL.n464 VTAIL.n463 0.155672
R1184 VTAIL.n463 VTAIL.n407 0.155672
R1185 VTAIL.n456 VTAIL.n407 0.155672
R1186 VTAIL.n456 VTAIL.n455 0.155672
R1187 VTAIL.n455 VTAIL.n411 0.155672
R1188 VTAIL.n448 VTAIL.n411 0.155672
R1189 VTAIL.n448 VTAIL.n447 0.155672
R1190 VTAIL.n447 VTAIL.n415 0.155672
R1191 VTAIL.n440 VTAIL.n415 0.155672
R1192 VTAIL.n440 VTAIL.n439 0.155672
R1193 VTAIL.n439 VTAIL.n419 0.155672
R1194 VTAIL.n432 VTAIL.n419 0.155672
R1195 VTAIL.n432 VTAIL.n431 0.155672
R1196 VTAIL.n431 VTAIL.n423 0.155672
R1197 VTAIL.n389 VTAIL.n295 0.155672
R1198 VTAIL.n382 VTAIL.n295 0.155672
R1199 VTAIL.n382 VTAIL.n381 0.155672
R1200 VTAIL.n381 VTAIL.n299 0.155672
R1201 VTAIL.n374 VTAIL.n299 0.155672
R1202 VTAIL.n374 VTAIL.n373 0.155672
R1203 VTAIL.n373 VTAIL.n303 0.155672
R1204 VTAIL.n366 VTAIL.n303 0.155672
R1205 VTAIL.n366 VTAIL.n365 0.155672
R1206 VTAIL.n365 VTAIL.n309 0.155672
R1207 VTAIL.n358 VTAIL.n309 0.155672
R1208 VTAIL.n358 VTAIL.n357 0.155672
R1209 VTAIL.n357 VTAIL.n313 0.155672
R1210 VTAIL.n350 VTAIL.n313 0.155672
R1211 VTAIL.n350 VTAIL.n349 0.155672
R1212 VTAIL.n349 VTAIL.n317 0.155672
R1213 VTAIL.n342 VTAIL.n317 0.155672
R1214 VTAIL.n342 VTAIL.n341 0.155672
R1215 VTAIL.n341 VTAIL.n321 0.155672
R1216 VTAIL.n334 VTAIL.n321 0.155672
R1217 VTAIL.n334 VTAIL.n333 0.155672
R1218 VTAIL.n333 VTAIL.n325 0.155672
R1219 VDD1 VDD1.n1 114.261
R1220 VDD1 VDD1.n0 63.6492
R1221 VDD1.n0 VDD1.t2 1.12104
R1222 VDD1.n0 VDD1.t0 1.12104
R1223 VDD1.n1 VDD1.t1 1.12104
R1224 VDD1.n1 VDD1.t3 1.12104
R1225 B.n766 B.n765 585
R1226 B.n767 B.n155 585
R1227 B.n769 B.n768 585
R1228 B.n771 B.n154 585
R1229 B.n774 B.n773 585
R1230 B.n775 B.n153 585
R1231 B.n777 B.n776 585
R1232 B.n779 B.n152 585
R1233 B.n782 B.n781 585
R1234 B.n783 B.n151 585
R1235 B.n785 B.n784 585
R1236 B.n787 B.n150 585
R1237 B.n790 B.n789 585
R1238 B.n791 B.n149 585
R1239 B.n793 B.n792 585
R1240 B.n795 B.n148 585
R1241 B.n798 B.n797 585
R1242 B.n799 B.n147 585
R1243 B.n801 B.n800 585
R1244 B.n803 B.n146 585
R1245 B.n806 B.n805 585
R1246 B.n807 B.n145 585
R1247 B.n809 B.n808 585
R1248 B.n811 B.n144 585
R1249 B.n814 B.n813 585
R1250 B.n815 B.n143 585
R1251 B.n817 B.n816 585
R1252 B.n819 B.n142 585
R1253 B.n822 B.n821 585
R1254 B.n823 B.n141 585
R1255 B.n825 B.n824 585
R1256 B.n827 B.n140 585
R1257 B.n830 B.n829 585
R1258 B.n831 B.n139 585
R1259 B.n833 B.n832 585
R1260 B.n835 B.n138 585
R1261 B.n838 B.n837 585
R1262 B.n839 B.n137 585
R1263 B.n841 B.n840 585
R1264 B.n843 B.n136 585
R1265 B.n846 B.n845 585
R1266 B.n847 B.n135 585
R1267 B.n849 B.n848 585
R1268 B.n851 B.n134 585
R1269 B.n854 B.n853 585
R1270 B.n855 B.n133 585
R1271 B.n857 B.n856 585
R1272 B.n859 B.n132 585
R1273 B.n862 B.n861 585
R1274 B.n863 B.n131 585
R1275 B.n865 B.n864 585
R1276 B.n867 B.n130 585
R1277 B.n870 B.n869 585
R1278 B.n871 B.n129 585
R1279 B.n873 B.n872 585
R1280 B.n875 B.n128 585
R1281 B.n877 B.n876 585
R1282 B.n879 B.n878 585
R1283 B.n882 B.n881 585
R1284 B.n883 B.n123 585
R1285 B.n885 B.n884 585
R1286 B.n887 B.n122 585
R1287 B.n890 B.n889 585
R1288 B.n891 B.n121 585
R1289 B.n893 B.n892 585
R1290 B.n895 B.n120 585
R1291 B.n897 B.n896 585
R1292 B.n899 B.n898 585
R1293 B.n902 B.n901 585
R1294 B.n903 B.n115 585
R1295 B.n905 B.n904 585
R1296 B.n907 B.n114 585
R1297 B.n910 B.n909 585
R1298 B.n911 B.n113 585
R1299 B.n913 B.n912 585
R1300 B.n915 B.n112 585
R1301 B.n918 B.n917 585
R1302 B.n919 B.n111 585
R1303 B.n921 B.n920 585
R1304 B.n923 B.n110 585
R1305 B.n926 B.n925 585
R1306 B.n927 B.n109 585
R1307 B.n929 B.n928 585
R1308 B.n931 B.n108 585
R1309 B.n934 B.n933 585
R1310 B.n935 B.n107 585
R1311 B.n937 B.n936 585
R1312 B.n939 B.n106 585
R1313 B.n942 B.n941 585
R1314 B.n943 B.n105 585
R1315 B.n945 B.n944 585
R1316 B.n947 B.n104 585
R1317 B.n950 B.n949 585
R1318 B.n951 B.n103 585
R1319 B.n953 B.n952 585
R1320 B.n955 B.n102 585
R1321 B.n958 B.n957 585
R1322 B.n959 B.n101 585
R1323 B.n961 B.n960 585
R1324 B.n963 B.n100 585
R1325 B.n966 B.n965 585
R1326 B.n967 B.n99 585
R1327 B.n969 B.n968 585
R1328 B.n971 B.n98 585
R1329 B.n974 B.n973 585
R1330 B.n975 B.n97 585
R1331 B.n977 B.n976 585
R1332 B.n979 B.n96 585
R1333 B.n982 B.n981 585
R1334 B.n983 B.n95 585
R1335 B.n985 B.n984 585
R1336 B.n987 B.n94 585
R1337 B.n990 B.n989 585
R1338 B.n991 B.n93 585
R1339 B.n993 B.n992 585
R1340 B.n995 B.n92 585
R1341 B.n998 B.n997 585
R1342 B.n999 B.n91 585
R1343 B.n1001 B.n1000 585
R1344 B.n1003 B.n90 585
R1345 B.n1006 B.n1005 585
R1346 B.n1007 B.n89 585
R1347 B.n1009 B.n1008 585
R1348 B.n1011 B.n88 585
R1349 B.n1014 B.n1013 585
R1350 B.n1015 B.n87 585
R1351 B.n763 B.n85 585
R1352 B.n1018 B.n85 585
R1353 B.n762 B.n84 585
R1354 B.n1019 B.n84 585
R1355 B.n761 B.n83 585
R1356 B.n1020 B.n83 585
R1357 B.n760 B.n759 585
R1358 B.n759 B.n79 585
R1359 B.n758 B.n78 585
R1360 B.n1026 B.n78 585
R1361 B.n757 B.n77 585
R1362 B.n1027 B.n77 585
R1363 B.n756 B.n76 585
R1364 B.n1028 B.n76 585
R1365 B.n755 B.n754 585
R1366 B.n754 B.n72 585
R1367 B.n753 B.n71 585
R1368 B.n1034 B.n71 585
R1369 B.n752 B.n70 585
R1370 B.n1035 B.n70 585
R1371 B.n751 B.n69 585
R1372 B.n1036 B.n69 585
R1373 B.n750 B.n749 585
R1374 B.n749 B.n65 585
R1375 B.n748 B.n64 585
R1376 B.n1042 B.n64 585
R1377 B.n747 B.n63 585
R1378 B.n1043 B.n63 585
R1379 B.n746 B.n62 585
R1380 B.n1044 B.n62 585
R1381 B.n745 B.n744 585
R1382 B.n744 B.n58 585
R1383 B.n743 B.n57 585
R1384 B.n1050 B.n57 585
R1385 B.n742 B.n56 585
R1386 B.n1051 B.n56 585
R1387 B.n741 B.n55 585
R1388 B.n1052 B.n55 585
R1389 B.n740 B.n739 585
R1390 B.n739 B.n51 585
R1391 B.n738 B.n50 585
R1392 B.n1058 B.n50 585
R1393 B.n737 B.n49 585
R1394 B.n1059 B.n49 585
R1395 B.n736 B.n48 585
R1396 B.n1060 B.n48 585
R1397 B.n735 B.n734 585
R1398 B.n734 B.n44 585
R1399 B.n733 B.n43 585
R1400 B.n1066 B.n43 585
R1401 B.n732 B.n42 585
R1402 B.n1067 B.n42 585
R1403 B.n731 B.n41 585
R1404 B.n1068 B.n41 585
R1405 B.n730 B.n729 585
R1406 B.n729 B.n37 585
R1407 B.n728 B.n36 585
R1408 B.n1074 B.n36 585
R1409 B.n727 B.n35 585
R1410 B.n1075 B.n35 585
R1411 B.n726 B.n34 585
R1412 B.n1076 B.n34 585
R1413 B.n725 B.n724 585
R1414 B.n724 B.n30 585
R1415 B.n723 B.n29 585
R1416 B.n1082 B.n29 585
R1417 B.n722 B.n28 585
R1418 B.n1083 B.n28 585
R1419 B.n721 B.n27 585
R1420 B.n1084 B.n27 585
R1421 B.n720 B.n719 585
R1422 B.n719 B.n23 585
R1423 B.n718 B.n22 585
R1424 B.n1090 B.n22 585
R1425 B.n717 B.n21 585
R1426 B.n1091 B.n21 585
R1427 B.n716 B.n20 585
R1428 B.n1092 B.n20 585
R1429 B.n715 B.n714 585
R1430 B.n714 B.n16 585
R1431 B.n713 B.n15 585
R1432 B.n1098 B.n15 585
R1433 B.n712 B.n14 585
R1434 B.n1099 B.n14 585
R1435 B.n711 B.n13 585
R1436 B.n1100 B.n13 585
R1437 B.n710 B.n709 585
R1438 B.n709 B.n12 585
R1439 B.n708 B.n707 585
R1440 B.n708 B.n8 585
R1441 B.n706 B.n7 585
R1442 B.n1107 B.n7 585
R1443 B.n705 B.n6 585
R1444 B.n1108 B.n6 585
R1445 B.n704 B.n5 585
R1446 B.n1109 B.n5 585
R1447 B.n703 B.n702 585
R1448 B.n702 B.n4 585
R1449 B.n701 B.n156 585
R1450 B.n701 B.n700 585
R1451 B.n691 B.n157 585
R1452 B.n158 B.n157 585
R1453 B.n693 B.n692 585
R1454 B.n694 B.n693 585
R1455 B.n690 B.n163 585
R1456 B.n163 B.n162 585
R1457 B.n689 B.n688 585
R1458 B.n688 B.n687 585
R1459 B.n165 B.n164 585
R1460 B.n166 B.n165 585
R1461 B.n680 B.n679 585
R1462 B.n681 B.n680 585
R1463 B.n678 B.n171 585
R1464 B.n171 B.n170 585
R1465 B.n677 B.n676 585
R1466 B.n676 B.n675 585
R1467 B.n173 B.n172 585
R1468 B.n174 B.n173 585
R1469 B.n668 B.n667 585
R1470 B.n669 B.n668 585
R1471 B.n666 B.n179 585
R1472 B.n179 B.n178 585
R1473 B.n665 B.n664 585
R1474 B.n664 B.n663 585
R1475 B.n181 B.n180 585
R1476 B.n182 B.n181 585
R1477 B.n656 B.n655 585
R1478 B.n657 B.n656 585
R1479 B.n654 B.n187 585
R1480 B.n187 B.n186 585
R1481 B.n653 B.n652 585
R1482 B.n652 B.n651 585
R1483 B.n189 B.n188 585
R1484 B.n190 B.n189 585
R1485 B.n644 B.n643 585
R1486 B.n645 B.n644 585
R1487 B.n642 B.n194 585
R1488 B.n198 B.n194 585
R1489 B.n641 B.n640 585
R1490 B.n640 B.n639 585
R1491 B.n196 B.n195 585
R1492 B.n197 B.n196 585
R1493 B.n632 B.n631 585
R1494 B.n633 B.n632 585
R1495 B.n630 B.n203 585
R1496 B.n203 B.n202 585
R1497 B.n629 B.n628 585
R1498 B.n628 B.n627 585
R1499 B.n205 B.n204 585
R1500 B.n206 B.n205 585
R1501 B.n620 B.n619 585
R1502 B.n621 B.n620 585
R1503 B.n618 B.n211 585
R1504 B.n211 B.n210 585
R1505 B.n617 B.n616 585
R1506 B.n616 B.n615 585
R1507 B.n213 B.n212 585
R1508 B.n214 B.n213 585
R1509 B.n608 B.n607 585
R1510 B.n609 B.n608 585
R1511 B.n606 B.n219 585
R1512 B.n219 B.n218 585
R1513 B.n605 B.n604 585
R1514 B.n604 B.n603 585
R1515 B.n221 B.n220 585
R1516 B.n222 B.n221 585
R1517 B.n596 B.n595 585
R1518 B.n597 B.n596 585
R1519 B.n594 B.n226 585
R1520 B.n230 B.n226 585
R1521 B.n593 B.n592 585
R1522 B.n592 B.n591 585
R1523 B.n228 B.n227 585
R1524 B.n229 B.n228 585
R1525 B.n584 B.n583 585
R1526 B.n585 B.n584 585
R1527 B.n582 B.n235 585
R1528 B.n235 B.n234 585
R1529 B.n581 B.n580 585
R1530 B.n580 B.n579 585
R1531 B.n237 B.n236 585
R1532 B.n238 B.n237 585
R1533 B.n572 B.n571 585
R1534 B.n573 B.n572 585
R1535 B.n570 B.n243 585
R1536 B.n243 B.n242 585
R1537 B.n569 B.n568 585
R1538 B.n568 B.n567 585
R1539 B.n564 B.n247 585
R1540 B.n563 B.n562 585
R1541 B.n560 B.n248 585
R1542 B.n560 B.n246 585
R1543 B.n559 B.n558 585
R1544 B.n557 B.n556 585
R1545 B.n555 B.n250 585
R1546 B.n553 B.n552 585
R1547 B.n551 B.n251 585
R1548 B.n550 B.n549 585
R1549 B.n547 B.n252 585
R1550 B.n545 B.n544 585
R1551 B.n543 B.n253 585
R1552 B.n542 B.n541 585
R1553 B.n539 B.n254 585
R1554 B.n537 B.n536 585
R1555 B.n535 B.n255 585
R1556 B.n534 B.n533 585
R1557 B.n531 B.n256 585
R1558 B.n529 B.n528 585
R1559 B.n527 B.n257 585
R1560 B.n526 B.n525 585
R1561 B.n523 B.n258 585
R1562 B.n521 B.n520 585
R1563 B.n519 B.n259 585
R1564 B.n518 B.n517 585
R1565 B.n515 B.n260 585
R1566 B.n513 B.n512 585
R1567 B.n511 B.n261 585
R1568 B.n510 B.n509 585
R1569 B.n507 B.n262 585
R1570 B.n505 B.n504 585
R1571 B.n503 B.n263 585
R1572 B.n502 B.n501 585
R1573 B.n499 B.n264 585
R1574 B.n497 B.n496 585
R1575 B.n495 B.n265 585
R1576 B.n494 B.n493 585
R1577 B.n491 B.n266 585
R1578 B.n489 B.n488 585
R1579 B.n487 B.n267 585
R1580 B.n486 B.n485 585
R1581 B.n483 B.n268 585
R1582 B.n481 B.n480 585
R1583 B.n479 B.n269 585
R1584 B.n478 B.n477 585
R1585 B.n475 B.n270 585
R1586 B.n473 B.n472 585
R1587 B.n471 B.n271 585
R1588 B.n470 B.n469 585
R1589 B.n467 B.n272 585
R1590 B.n465 B.n464 585
R1591 B.n463 B.n273 585
R1592 B.n462 B.n461 585
R1593 B.n459 B.n274 585
R1594 B.n457 B.n456 585
R1595 B.n455 B.n275 585
R1596 B.n454 B.n453 585
R1597 B.n451 B.n276 585
R1598 B.n449 B.n448 585
R1599 B.n447 B.n277 585
R1600 B.n446 B.n445 585
R1601 B.n443 B.n281 585
R1602 B.n441 B.n440 585
R1603 B.n439 B.n282 585
R1604 B.n438 B.n437 585
R1605 B.n435 B.n283 585
R1606 B.n433 B.n432 585
R1607 B.n431 B.n284 585
R1608 B.n429 B.n428 585
R1609 B.n426 B.n287 585
R1610 B.n424 B.n423 585
R1611 B.n422 B.n288 585
R1612 B.n421 B.n420 585
R1613 B.n418 B.n289 585
R1614 B.n416 B.n415 585
R1615 B.n414 B.n290 585
R1616 B.n413 B.n412 585
R1617 B.n410 B.n291 585
R1618 B.n408 B.n407 585
R1619 B.n406 B.n292 585
R1620 B.n405 B.n404 585
R1621 B.n402 B.n293 585
R1622 B.n400 B.n399 585
R1623 B.n398 B.n294 585
R1624 B.n397 B.n396 585
R1625 B.n394 B.n295 585
R1626 B.n392 B.n391 585
R1627 B.n390 B.n296 585
R1628 B.n389 B.n388 585
R1629 B.n386 B.n297 585
R1630 B.n384 B.n383 585
R1631 B.n382 B.n298 585
R1632 B.n381 B.n380 585
R1633 B.n378 B.n299 585
R1634 B.n376 B.n375 585
R1635 B.n374 B.n300 585
R1636 B.n373 B.n372 585
R1637 B.n370 B.n301 585
R1638 B.n368 B.n367 585
R1639 B.n366 B.n302 585
R1640 B.n365 B.n364 585
R1641 B.n362 B.n303 585
R1642 B.n360 B.n359 585
R1643 B.n358 B.n304 585
R1644 B.n357 B.n356 585
R1645 B.n354 B.n305 585
R1646 B.n352 B.n351 585
R1647 B.n350 B.n306 585
R1648 B.n349 B.n348 585
R1649 B.n346 B.n307 585
R1650 B.n344 B.n343 585
R1651 B.n342 B.n308 585
R1652 B.n341 B.n340 585
R1653 B.n338 B.n309 585
R1654 B.n336 B.n335 585
R1655 B.n334 B.n310 585
R1656 B.n333 B.n332 585
R1657 B.n330 B.n311 585
R1658 B.n328 B.n327 585
R1659 B.n326 B.n312 585
R1660 B.n325 B.n324 585
R1661 B.n322 B.n313 585
R1662 B.n320 B.n319 585
R1663 B.n318 B.n314 585
R1664 B.n317 B.n316 585
R1665 B.n245 B.n244 585
R1666 B.n246 B.n245 585
R1667 B.n566 B.n565 585
R1668 B.n567 B.n566 585
R1669 B.n241 B.n240 585
R1670 B.n242 B.n241 585
R1671 B.n575 B.n574 585
R1672 B.n574 B.n573 585
R1673 B.n576 B.n239 585
R1674 B.n239 B.n238 585
R1675 B.n578 B.n577 585
R1676 B.n579 B.n578 585
R1677 B.n233 B.n232 585
R1678 B.n234 B.n233 585
R1679 B.n587 B.n586 585
R1680 B.n586 B.n585 585
R1681 B.n588 B.n231 585
R1682 B.n231 B.n229 585
R1683 B.n590 B.n589 585
R1684 B.n591 B.n590 585
R1685 B.n225 B.n224 585
R1686 B.n230 B.n225 585
R1687 B.n599 B.n598 585
R1688 B.n598 B.n597 585
R1689 B.n600 B.n223 585
R1690 B.n223 B.n222 585
R1691 B.n602 B.n601 585
R1692 B.n603 B.n602 585
R1693 B.n217 B.n216 585
R1694 B.n218 B.n217 585
R1695 B.n611 B.n610 585
R1696 B.n610 B.n609 585
R1697 B.n612 B.n215 585
R1698 B.n215 B.n214 585
R1699 B.n614 B.n613 585
R1700 B.n615 B.n614 585
R1701 B.n209 B.n208 585
R1702 B.n210 B.n209 585
R1703 B.n623 B.n622 585
R1704 B.n622 B.n621 585
R1705 B.n624 B.n207 585
R1706 B.n207 B.n206 585
R1707 B.n626 B.n625 585
R1708 B.n627 B.n626 585
R1709 B.n201 B.n200 585
R1710 B.n202 B.n201 585
R1711 B.n635 B.n634 585
R1712 B.n634 B.n633 585
R1713 B.n636 B.n199 585
R1714 B.n199 B.n197 585
R1715 B.n638 B.n637 585
R1716 B.n639 B.n638 585
R1717 B.n193 B.n192 585
R1718 B.n198 B.n193 585
R1719 B.n647 B.n646 585
R1720 B.n646 B.n645 585
R1721 B.n648 B.n191 585
R1722 B.n191 B.n190 585
R1723 B.n650 B.n649 585
R1724 B.n651 B.n650 585
R1725 B.n185 B.n184 585
R1726 B.n186 B.n185 585
R1727 B.n659 B.n658 585
R1728 B.n658 B.n657 585
R1729 B.n660 B.n183 585
R1730 B.n183 B.n182 585
R1731 B.n662 B.n661 585
R1732 B.n663 B.n662 585
R1733 B.n177 B.n176 585
R1734 B.n178 B.n177 585
R1735 B.n671 B.n670 585
R1736 B.n670 B.n669 585
R1737 B.n672 B.n175 585
R1738 B.n175 B.n174 585
R1739 B.n674 B.n673 585
R1740 B.n675 B.n674 585
R1741 B.n169 B.n168 585
R1742 B.n170 B.n169 585
R1743 B.n683 B.n682 585
R1744 B.n682 B.n681 585
R1745 B.n684 B.n167 585
R1746 B.n167 B.n166 585
R1747 B.n686 B.n685 585
R1748 B.n687 B.n686 585
R1749 B.n161 B.n160 585
R1750 B.n162 B.n161 585
R1751 B.n696 B.n695 585
R1752 B.n695 B.n694 585
R1753 B.n697 B.n159 585
R1754 B.n159 B.n158 585
R1755 B.n699 B.n698 585
R1756 B.n700 B.n699 585
R1757 B.n3 B.n0 585
R1758 B.n4 B.n3 585
R1759 B.n1106 B.n1 585
R1760 B.n1107 B.n1106 585
R1761 B.n1105 B.n1104 585
R1762 B.n1105 B.n8 585
R1763 B.n1103 B.n9 585
R1764 B.n12 B.n9 585
R1765 B.n1102 B.n1101 585
R1766 B.n1101 B.n1100 585
R1767 B.n11 B.n10 585
R1768 B.n1099 B.n11 585
R1769 B.n1097 B.n1096 585
R1770 B.n1098 B.n1097 585
R1771 B.n1095 B.n17 585
R1772 B.n17 B.n16 585
R1773 B.n1094 B.n1093 585
R1774 B.n1093 B.n1092 585
R1775 B.n19 B.n18 585
R1776 B.n1091 B.n19 585
R1777 B.n1089 B.n1088 585
R1778 B.n1090 B.n1089 585
R1779 B.n1087 B.n24 585
R1780 B.n24 B.n23 585
R1781 B.n1086 B.n1085 585
R1782 B.n1085 B.n1084 585
R1783 B.n26 B.n25 585
R1784 B.n1083 B.n26 585
R1785 B.n1081 B.n1080 585
R1786 B.n1082 B.n1081 585
R1787 B.n1079 B.n31 585
R1788 B.n31 B.n30 585
R1789 B.n1078 B.n1077 585
R1790 B.n1077 B.n1076 585
R1791 B.n33 B.n32 585
R1792 B.n1075 B.n33 585
R1793 B.n1073 B.n1072 585
R1794 B.n1074 B.n1073 585
R1795 B.n1071 B.n38 585
R1796 B.n38 B.n37 585
R1797 B.n1070 B.n1069 585
R1798 B.n1069 B.n1068 585
R1799 B.n40 B.n39 585
R1800 B.n1067 B.n40 585
R1801 B.n1065 B.n1064 585
R1802 B.n1066 B.n1065 585
R1803 B.n1063 B.n45 585
R1804 B.n45 B.n44 585
R1805 B.n1062 B.n1061 585
R1806 B.n1061 B.n1060 585
R1807 B.n47 B.n46 585
R1808 B.n1059 B.n47 585
R1809 B.n1057 B.n1056 585
R1810 B.n1058 B.n1057 585
R1811 B.n1055 B.n52 585
R1812 B.n52 B.n51 585
R1813 B.n1054 B.n1053 585
R1814 B.n1053 B.n1052 585
R1815 B.n54 B.n53 585
R1816 B.n1051 B.n54 585
R1817 B.n1049 B.n1048 585
R1818 B.n1050 B.n1049 585
R1819 B.n1047 B.n59 585
R1820 B.n59 B.n58 585
R1821 B.n1046 B.n1045 585
R1822 B.n1045 B.n1044 585
R1823 B.n61 B.n60 585
R1824 B.n1043 B.n61 585
R1825 B.n1041 B.n1040 585
R1826 B.n1042 B.n1041 585
R1827 B.n1039 B.n66 585
R1828 B.n66 B.n65 585
R1829 B.n1038 B.n1037 585
R1830 B.n1037 B.n1036 585
R1831 B.n68 B.n67 585
R1832 B.n1035 B.n68 585
R1833 B.n1033 B.n1032 585
R1834 B.n1034 B.n1033 585
R1835 B.n1031 B.n73 585
R1836 B.n73 B.n72 585
R1837 B.n1030 B.n1029 585
R1838 B.n1029 B.n1028 585
R1839 B.n75 B.n74 585
R1840 B.n1027 B.n75 585
R1841 B.n1025 B.n1024 585
R1842 B.n1026 B.n1025 585
R1843 B.n1023 B.n80 585
R1844 B.n80 B.n79 585
R1845 B.n1022 B.n1021 585
R1846 B.n1021 B.n1020 585
R1847 B.n82 B.n81 585
R1848 B.n1019 B.n82 585
R1849 B.n1017 B.n1016 585
R1850 B.n1018 B.n1017 585
R1851 B.n1110 B.n1109 585
R1852 B.n1108 B.n2 585
R1853 B.n1017 B.n87 482.89
R1854 B.n765 B.n85 482.89
R1855 B.n568 B.n245 482.89
R1856 B.n566 B.n247 482.89
R1857 B.n116 B.t6 464.144
R1858 B.n278 B.t17 464.144
R1859 B.n124 B.t13 464.144
R1860 B.n285 B.t11 464.144
R1861 B.n125 B.t14 380.168
R1862 B.n286 B.t10 380.168
R1863 B.n117 B.t7 380.168
R1864 B.n279 B.t16 380.168
R1865 B.n116 B.t4 315.954
R1866 B.n124 B.t12 315.954
R1867 B.n285 B.t8 315.954
R1868 B.n278 B.t15 315.954
R1869 B.n764 B.n86 256.663
R1870 B.n770 B.n86 256.663
R1871 B.n772 B.n86 256.663
R1872 B.n778 B.n86 256.663
R1873 B.n780 B.n86 256.663
R1874 B.n786 B.n86 256.663
R1875 B.n788 B.n86 256.663
R1876 B.n794 B.n86 256.663
R1877 B.n796 B.n86 256.663
R1878 B.n802 B.n86 256.663
R1879 B.n804 B.n86 256.663
R1880 B.n810 B.n86 256.663
R1881 B.n812 B.n86 256.663
R1882 B.n818 B.n86 256.663
R1883 B.n820 B.n86 256.663
R1884 B.n826 B.n86 256.663
R1885 B.n828 B.n86 256.663
R1886 B.n834 B.n86 256.663
R1887 B.n836 B.n86 256.663
R1888 B.n842 B.n86 256.663
R1889 B.n844 B.n86 256.663
R1890 B.n850 B.n86 256.663
R1891 B.n852 B.n86 256.663
R1892 B.n858 B.n86 256.663
R1893 B.n860 B.n86 256.663
R1894 B.n866 B.n86 256.663
R1895 B.n868 B.n86 256.663
R1896 B.n874 B.n86 256.663
R1897 B.n127 B.n86 256.663
R1898 B.n880 B.n86 256.663
R1899 B.n886 B.n86 256.663
R1900 B.n888 B.n86 256.663
R1901 B.n894 B.n86 256.663
R1902 B.n119 B.n86 256.663
R1903 B.n900 B.n86 256.663
R1904 B.n906 B.n86 256.663
R1905 B.n908 B.n86 256.663
R1906 B.n914 B.n86 256.663
R1907 B.n916 B.n86 256.663
R1908 B.n922 B.n86 256.663
R1909 B.n924 B.n86 256.663
R1910 B.n930 B.n86 256.663
R1911 B.n932 B.n86 256.663
R1912 B.n938 B.n86 256.663
R1913 B.n940 B.n86 256.663
R1914 B.n946 B.n86 256.663
R1915 B.n948 B.n86 256.663
R1916 B.n954 B.n86 256.663
R1917 B.n956 B.n86 256.663
R1918 B.n962 B.n86 256.663
R1919 B.n964 B.n86 256.663
R1920 B.n970 B.n86 256.663
R1921 B.n972 B.n86 256.663
R1922 B.n978 B.n86 256.663
R1923 B.n980 B.n86 256.663
R1924 B.n986 B.n86 256.663
R1925 B.n988 B.n86 256.663
R1926 B.n994 B.n86 256.663
R1927 B.n996 B.n86 256.663
R1928 B.n1002 B.n86 256.663
R1929 B.n1004 B.n86 256.663
R1930 B.n1010 B.n86 256.663
R1931 B.n1012 B.n86 256.663
R1932 B.n561 B.n246 256.663
R1933 B.n249 B.n246 256.663
R1934 B.n554 B.n246 256.663
R1935 B.n548 B.n246 256.663
R1936 B.n546 B.n246 256.663
R1937 B.n540 B.n246 256.663
R1938 B.n538 B.n246 256.663
R1939 B.n532 B.n246 256.663
R1940 B.n530 B.n246 256.663
R1941 B.n524 B.n246 256.663
R1942 B.n522 B.n246 256.663
R1943 B.n516 B.n246 256.663
R1944 B.n514 B.n246 256.663
R1945 B.n508 B.n246 256.663
R1946 B.n506 B.n246 256.663
R1947 B.n500 B.n246 256.663
R1948 B.n498 B.n246 256.663
R1949 B.n492 B.n246 256.663
R1950 B.n490 B.n246 256.663
R1951 B.n484 B.n246 256.663
R1952 B.n482 B.n246 256.663
R1953 B.n476 B.n246 256.663
R1954 B.n474 B.n246 256.663
R1955 B.n468 B.n246 256.663
R1956 B.n466 B.n246 256.663
R1957 B.n460 B.n246 256.663
R1958 B.n458 B.n246 256.663
R1959 B.n452 B.n246 256.663
R1960 B.n450 B.n246 256.663
R1961 B.n444 B.n246 256.663
R1962 B.n442 B.n246 256.663
R1963 B.n436 B.n246 256.663
R1964 B.n434 B.n246 256.663
R1965 B.n427 B.n246 256.663
R1966 B.n425 B.n246 256.663
R1967 B.n419 B.n246 256.663
R1968 B.n417 B.n246 256.663
R1969 B.n411 B.n246 256.663
R1970 B.n409 B.n246 256.663
R1971 B.n403 B.n246 256.663
R1972 B.n401 B.n246 256.663
R1973 B.n395 B.n246 256.663
R1974 B.n393 B.n246 256.663
R1975 B.n387 B.n246 256.663
R1976 B.n385 B.n246 256.663
R1977 B.n379 B.n246 256.663
R1978 B.n377 B.n246 256.663
R1979 B.n371 B.n246 256.663
R1980 B.n369 B.n246 256.663
R1981 B.n363 B.n246 256.663
R1982 B.n361 B.n246 256.663
R1983 B.n355 B.n246 256.663
R1984 B.n353 B.n246 256.663
R1985 B.n347 B.n246 256.663
R1986 B.n345 B.n246 256.663
R1987 B.n339 B.n246 256.663
R1988 B.n337 B.n246 256.663
R1989 B.n331 B.n246 256.663
R1990 B.n329 B.n246 256.663
R1991 B.n323 B.n246 256.663
R1992 B.n321 B.n246 256.663
R1993 B.n315 B.n246 256.663
R1994 B.n1112 B.n1111 256.663
R1995 B.n1013 B.n1011 163.367
R1996 B.n1009 B.n89 163.367
R1997 B.n1005 B.n1003 163.367
R1998 B.n1001 B.n91 163.367
R1999 B.n997 B.n995 163.367
R2000 B.n993 B.n93 163.367
R2001 B.n989 B.n987 163.367
R2002 B.n985 B.n95 163.367
R2003 B.n981 B.n979 163.367
R2004 B.n977 B.n97 163.367
R2005 B.n973 B.n971 163.367
R2006 B.n969 B.n99 163.367
R2007 B.n965 B.n963 163.367
R2008 B.n961 B.n101 163.367
R2009 B.n957 B.n955 163.367
R2010 B.n953 B.n103 163.367
R2011 B.n949 B.n947 163.367
R2012 B.n945 B.n105 163.367
R2013 B.n941 B.n939 163.367
R2014 B.n937 B.n107 163.367
R2015 B.n933 B.n931 163.367
R2016 B.n929 B.n109 163.367
R2017 B.n925 B.n923 163.367
R2018 B.n921 B.n111 163.367
R2019 B.n917 B.n915 163.367
R2020 B.n913 B.n113 163.367
R2021 B.n909 B.n907 163.367
R2022 B.n905 B.n115 163.367
R2023 B.n901 B.n899 163.367
R2024 B.n896 B.n895 163.367
R2025 B.n893 B.n121 163.367
R2026 B.n889 B.n887 163.367
R2027 B.n885 B.n123 163.367
R2028 B.n881 B.n879 163.367
R2029 B.n876 B.n875 163.367
R2030 B.n873 B.n129 163.367
R2031 B.n869 B.n867 163.367
R2032 B.n865 B.n131 163.367
R2033 B.n861 B.n859 163.367
R2034 B.n857 B.n133 163.367
R2035 B.n853 B.n851 163.367
R2036 B.n849 B.n135 163.367
R2037 B.n845 B.n843 163.367
R2038 B.n841 B.n137 163.367
R2039 B.n837 B.n835 163.367
R2040 B.n833 B.n139 163.367
R2041 B.n829 B.n827 163.367
R2042 B.n825 B.n141 163.367
R2043 B.n821 B.n819 163.367
R2044 B.n817 B.n143 163.367
R2045 B.n813 B.n811 163.367
R2046 B.n809 B.n145 163.367
R2047 B.n805 B.n803 163.367
R2048 B.n801 B.n147 163.367
R2049 B.n797 B.n795 163.367
R2050 B.n793 B.n149 163.367
R2051 B.n789 B.n787 163.367
R2052 B.n785 B.n151 163.367
R2053 B.n781 B.n779 163.367
R2054 B.n777 B.n153 163.367
R2055 B.n773 B.n771 163.367
R2056 B.n769 B.n155 163.367
R2057 B.n568 B.n243 163.367
R2058 B.n572 B.n243 163.367
R2059 B.n572 B.n237 163.367
R2060 B.n580 B.n237 163.367
R2061 B.n580 B.n235 163.367
R2062 B.n584 B.n235 163.367
R2063 B.n584 B.n228 163.367
R2064 B.n592 B.n228 163.367
R2065 B.n592 B.n226 163.367
R2066 B.n596 B.n226 163.367
R2067 B.n596 B.n221 163.367
R2068 B.n604 B.n221 163.367
R2069 B.n604 B.n219 163.367
R2070 B.n608 B.n219 163.367
R2071 B.n608 B.n213 163.367
R2072 B.n616 B.n213 163.367
R2073 B.n616 B.n211 163.367
R2074 B.n620 B.n211 163.367
R2075 B.n620 B.n205 163.367
R2076 B.n628 B.n205 163.367
R2077 B.n628 B.n203 163.367
R2078 B.n632 B.n203 163.367
R2079 B.n632 B.n196 163.367
R2080 B.n640 B.n196 163.367
R2081 B.n640 B.n194 163.367
R2082 B.n644 B.n194 163.367
R2083 B.n644 B.n189 163.367
R2084 B.n652 B.n189 163.367
R2085 B.n652 B.n187 163.367
R2086 B.n656 B.n187 163.367
R2087 B.n656 B.n181 163.367
R2088 B.n664 B.n181 163.367
R2089 B.n664 B.n179 163.367
R2090 B.n668 B.n179 163.367
R2091 B.n668 B.n173 163.367
R2092 B.n676 B.n173 163.367
R2093 B.n676 B.n171 163.367
R2094 B.n680 B.n171 163.367
R2095 B.n680 B.n165 163.367
R2096 B.n688 B.n165 163.367
R2097 B.n688 B.n163 163.367
R2098 B.n693 B.n163 163.367
R2099 B.n693 B.n157 163.367
R2100 B.n701 B.n157 163.367
R2101 B.n702 B.n701 163.367
R2102 B.n702 B.n5 163.367
R2103 B.n6 B.n5 163.367
R2104 B.n7 B.n6 163.367
R2105 B.n708 B.n7 163.367
R2106 B.n709 B.n708 163.367
R2107 B.n709 B.n13 163.367
R2108 B.n14 B.n13 163.367
R2109 B.n15 B.n14 163.367
R2110 B.n714 B.n15 163.367
R2111 B.n714 B.n20 163.367
R2112 B.n21 B.n20 163.367
R2113 B.n22 B.n21 163.367
R2114 B.n719 B.n22 163.367
R2115 B.n719 B.n27 163.367
R2116 B.n28 B.n27 163.367
R2117 B.n29 B.n28 163.367
R2118 B.n724 B.n29 163.367
R2119 B.n724 B.n34 163.367
R2120 B.n35 B.n34 163.367
R2121 B.n36 B.n35 163.367
R2122 B.n729 B.n36 163.367
R2123 B.n729 B.n41 163.367
R2124 B.n42 B.n41 163.367
R2125 B.n43 B.n42 163.367
R2126 B.n734 B.n43 163.367
R2127 B.n734 B.n48 163.367
R2128 B.n49 B.n48 163.367
R2129 B.n50 B.n49 163.367
R2130 B.n739 B.n50 163.367
R2131 B.n739 B.n55 163.367
R2132 B.n56 B.n55 163.367
R2133 B.n57 B.n56 163.367
R2134 B.n744 B.n57 163.367
R2135 B.n744 B.n62 163.367
R2136 B.n63 B.n62 163.367
R2137 B.n64 B.n63 163.367
R2138 B.n749 B.n64 163.367
R2139 B.n749 B.n69 163.367
R2140 B.n70 B.n69 163.367
R2141 B.n71 B.n70 163.367
R2142 B.n754 B.n71 163.367
R2143 B.n754 B.n76 163.367
R2144 B.n77 B.n76 163.367
R2145 B.n78 B.n77 163.367
R2146 B.n759 B.n78 163.367
R2147 B.n759 B.n83 163.367
R2148 B.n84 B.n83 163.367
R2149 B.n85 B.n84 163.367
R2150 B.n562 B.n560 163.367
R2151 B.n560 B.n559 163.367
R2152 B.n556 B.n555 163.367
R2153 B.n553 B.n251 163.367
R2154 B.n549 B.n547 163.367
R2155 B.n545 B.n253 163.367
R2156 B.n541 B.n539 163.367
R2157 B.n537 B.n255 163.367
R2158 B.n533 B.n531 163.367
R2159 B.n529 B.n257 163.367
R2160 B.n525 B.n523 163.367
R2161 B.n521 B.n259 163.367
R2162 B.n517 B.n515 163.367
R2163 B.n513 B.n261 163.367
R2164 B.n509 B.n507 163.367
R2165 B.n505 B.n263 163.367
R2166 B.n501 B.n499 163.367
R2167 B.n497 B.n265 163.367
R2168 B.n493 B.n491 163.367
R2169 B.n489 B.n267 163.367
R2170 B.n485 B.n483 163.367
R2171 B.n481 B.n269 163.367
R2172 B.n477 B.n475 163.367
R2173 B.n473 B.n271 163.367
R2174 B.n469 B.n467 163.367
R2175 B.n465 B.n273 163.367
R2176 B.n461 B.n459 163.367
R2177 B.n457 B.n275 163.367
R2178 B.n453 B.n451 163.367
R2179 B.n449 B.n277 163.367
R2180 B.n445 B.n443 163.367
R2181 B.n441 B.n282 163.367
R2182 B.n437 B.n435 163.367
R2183 B.n433 B.n284 163.367
R2184 B.n428 B.n426 163.367
R2185 B.n424 B.n288 163.367
R2186 B.n420 B.n418 163.367
R2187 B.n416 B.n290 163.367
R2188 B.n412 B.n410 163.367
R2189 B.n408 B.n292 163.367
R2190 B.n404 B.n402 163.367
R2191 B.n400 B.n294 163.367
R2192 B.n396 B.n394 163.367
R2193 B.n392 B.n296 163.367
R2194 B.n388 B.n386 163.367
R2195 B.n384 B.n298 163.367
R2196 B.n380 B.n378 163.367
R2197 B.n376 B.n300 163.367
R2198 B.n372 B.n370 163.367
R2199 B.n368 B.n302 163.367
R2200 B.n364 B.n362 163.367
R2201 B.n360 B.n304 163.367
R2202 B.n356 B.n354 163.367
R2203 B.n352 B.n306 163.367
R2204 B.n348 B.n346 163.367
R2205 B.n344 B.n308 163.367
R2206 B.n340 B.n338 163.367
R2207 B.n336 B.n310 163.367
R2208 B.n332 B.n330 163.367
R2209 B.n328 B.n312 163.367
R2210 B.n324 B.n322 163.367
R2211 B.n320 B.n314 163.367
R2212 B.n316 B.n245 163.367
R2213 B.n566 B.n241 163.367
R2214 B.n574 B.n241 163.367
R2215 B.n574 B.n239 163.367
R2216 B.n578 B.n239 163.367
R2217 B.n578 B.n233 163.367
R2218 B.n586 B.n233 163.367
R2219 B.n586 B.n231 163.367
R2220 B.n590 B.n231 163.367
R2221 B.n590 B.n225 163.367
R2222 B.n598 B.n225 163.367
R2223 B.n598 B.n223 163.367
R2224 B.n602 B.n223 163.367
R2225 B.n602 B.n217 163.367
R2226 B.n610 B.n217 163.367
R2227 B.n610 B.n215 163.367
R2228 B.n614 B.n215 163.367
R2229 B.n614 B.n209 163.367
R2230 B.n622 B.n209 163.367
R2231 B.n622 B.n207 163.367
R2232 B.n626 B.n207 163.367
R2233 B.n626 B.n201 163.367
R2234 B.n634 B.n201 163.367
R2235 B.n634 B.n199 163.367
R2236 B.n638 B.n199 163.367
R2237 B.n638 B.n193 163.367
R2238 B.n646 B.n193 163.367
R2239 B.n646 B.n191 163.367
R2240 B.n650 B.n191 163.367
R2241 B.n650 B.n185 163.367
R2242 B.n658 B.n185 163.367
R2243 B.n658 B.n183 163.367
R2244 B.n662 B.n183 163.367
R2245 B.n662 B.n177 163.367
R2246 B.n670 B.n177 163.367
R2247 B.n670 B.n175 163.367
R2248 B.n674 B.n175 163.367
R2249 B.n674 B.n169 163.367
R2250 B.n682 B.n169 163.367
R2251 B.n682 B.n167 163.367
R2252 B.n686 B.n167 163.367
R2253 B.n686 B.n161 163.367
R2254 B.n695 B.n161 163.367
R2255 B.n695 B.n159 163.367
R2256 B.n699 B.n159 163.367
R2257 B.n699 B.n3 163.367
R2258 B.n1110 B.n3 163.367
R2259 B.n1106 B.n2 163.367
R2260 B.n1106 B.n1105 163.367
R2261 B.n1105 B.n9 163.367
R2262 B.n1101 B.n9 163.367
R2263 B.n1101 B.n11 163.367
R2264 B.n1097 B.n11 163.367
R2265 B.n1097 B.n17 163.367
R2266 B.n1093 B.n17 163.367
R2267 B.n1093 B.n19 163.367
R2268 B.n1089 B.n19 163.367
R2269 B.n1089 B.n24 163.367
R2270 B.n1085 B.n24 163.367
R2271 B.n1085 B.n26 163.367
R2272 B.n1081 B.n26 163.367
R2273 B.n1081 B.n31 163.367
R2274 B.n1077 B.n31 163.367
R2275 B.n1077 B.n33 163.367
R2276 B.n1073 B.n33 163.367
R2277 B.n1073 B.n38 163.367
R2278 B.n1069 B.n38 163.367
R2279 B.n1069 B.n40 163.367
R2280 B.n1065 B.n40 163.367
R2281 B.n1065 B.n45 163.367
R2282 B.n1061 B.n45 163.367
R2283 B.n1061 B.n47 163.367
R2284 B.n1057 B.n47 163.367
R2285 B.n1057 B.n52 163.367
R2286 B.n1053 B.n52 163.367
R2287 B.n1053 B.n54 163.367
R2288 B.n1049 B.n54 163.367
R2289 B.n1049 B.n59 163.367
R2290 B.n1045 B.n59 163.367
R2291 B.n1045 B.n61 163.367
R2292 B.n1041 B.n61 163.367
R2293 B.n1041 B.n66 163.367
R2294 B.n1037 B.n66 163.367
R2295 B.n1037 B.n68 163.367
R2296 B.n1033 B.n68 163.367
R2297 B.n1033 B.n73 163.367
R2298 B.n1029 B.n73 163.367
R2299 B.n1029 B.n75 163.367
R2300 B.n1025 B.n75 163.367
R2301 B.n1025 B.n80 163.367
R2302 B.n1021 B.n80 163.367
R2303 B.n1021 B.n82 163.367
R2304 B.n1017 B.n82 163.367
R2305 B.n117 B.n116 83.9763
R2306 B.n125 B.n124 83.9763
R2307 B.n286 B.n285 83.9763
R2308 B.n279 B.n278 83.9763
R2309 B.n1012 B.n87 71.676
R2310 B.n1011 B.n1010 71.676
R2311 B.n1004 B.n89 71.676
R2312 B.n1003 B.n1002 71.676
R2313 B.n996 B.n91 71.676
R2314 B.n995 B.n994 71.676
R2315 B.n988 B.n93 71.676
R2316 B.n987 B.n986 71.676
R2317 B.n980 B.n95 71.676
R2318 B.n979 B.n978 71.676
R2319 B.n972 B.n97 71.676
R2320 B.n971 B.n970 71.676
R2321 B.n964 B.n99 71.676
R2322 B.n963 B.n962 71.676
R2323 B.n956 B.n101 71.676
R2324 B.n955 B.n954 71.676
R2325 B.n948 B.n103 71.676
R2326 B.n947 B.n946 71.676
R2327 B.n940 B.n105 71.676
R2328 B.n939 B.n938 71.676
R2329 B.n932 B.n107 71.676
R2330 B.n931 B.n930 71.676
R2331 B.n924 B.n109 71.676
R2332 B.n923 B.n922 71.676
R2333 B.n916 B.n111 71.676
R2334 B.n915 B.n914 71.676
R2335 B.n908 B.n113 71.676
R2336 B.n907 B.n906 71.676
R2337 B.n900 B.n115 71.676
R2338 B.n899 B.n119 71.676
R2339 B.n895 B.n894 71.676
R2340 B.n888 B.n121 71.676
R2341 B.n887 B.n886 71.676
R2342 B.n880 B.n123 71.676
R2343 B.n879 B.n127 71.676
R2344 B.n875 B.n874 71.676
R2345 B.n868 B.n129 71.676
R2346 B.n867 B.n866 71.676
R2347 B.n860 B.n131 71.676
R2348 B.n859 B.n858 71.676
R2349 B.n852 B.n133 71.676
R2350 B.n851 B.n850 71.676
R2351 B.n844 B.n135 71.676
R2352 B.n843 B.n842 71.676
R2353 B.n836 B.n137 71.676
R2354 B.n835 B.n834 71.676
R2355 B.n828 B.n139 71.676
R2356 B.n827 B.n826 71.676
R2357 B.n820 B.n141 71.676
R2358 B.n819 B.n818 71.676
R2359 B.n812 B.n143 71.676
R2360 B.n811 B.n810 71.676
R2361 B.n804 B.n145 71.676
R2362 B.n803 B.n802 71.676
R2363 B.n796 B.n147 71.676
R2364 B.n795 B.n794 71.676
R2365 B.n788 B.n149 71.676
R2366 B.n787 B.n786 71.676
R2367 B.n780 B.n151 71.676
R2368 B.n779 B.n778 71.676
R2369 B.n772 B.n153 71.676
R2370 B.n771 B.n770 71.676
R2371 B.n764 B.n155 71.676
R2372 B.n765 B.n764 71.676
R2373 B.n770 B.n769 71.676
R2374 B.n773 B.n772 71.676
R2375 B.n778 B.n777 71.676
R2376 B.n781 B.n780 71.676
R2377 B.n786 B.n785 71.676
R2378 B.n789 B.n788 71.676
R2379 B.n794 B.n793 71.676
R2380 B.n797 B.n796 71.676
R2381 B.n802 B.n801 71.676
R2382 B.n805 B.n804 71.676
R2383 B.n810 B.n809 71.676
R2384 B.n813 B.n812 71.676
R2385 B.n818 B.n817 71.676
R2386 B.n821 B.n820 71.676
R2387 B.n826 B.n825 71.676
R2388 B.n829 B.n828 71.676
R2389 B.n834 B.n833 71.676
R2390 B.n837 B.n836 71.676
R2391 B.n842 B.n841 71.676
R2392 B.n845 B.n844 71.676
R2393 B.n850 B.n849 71.676
R2394 B.n853 B.n852 71.676
R2395 B.n858 B.n857 71.676
R2396 B.n861 B.n860 71.676
R2397 B.n866 B.n865 71.676
R2398 B.n869 B.n868 71.676
R2399 B.n874 B.n873 71.676
R2400 B.n876 B.n127 71.676
R2401 B.n881 B.n880 71.676
R2402 B.n886 B.n885 71.676
R2403 B.n889 B.n888 71.676
R2404 B.n894 B.n893 71.676
R2405 B.n896 B.n119 71.676
R2406 B.n901 B.n900 71.676
R2407 B.n906 B.n905 71.676
R2408 B.n909 B.n908 71.676
R2409 B.n914 B.n913 71.676
R2410 B.n917 B.n916 71.676
R2411 B.n922 B.n921 71.676
R2412 B.n925 B.n924 71.676
R2413 B.n930 B.n929 71.676
R2414 B.n933 B.n932 71.676
R2415 B.n938 B.n937 71.676
R2416 B.n941 B.n940 71.676
R2417 B.n946 B.n945 71.676
R2418 B.n949 B.n948 71.676
R2419 B.n954 B.n953 71.676
R2420 B.n957 B.n956 71.676
R2421 B.n962 B.n961 71.676
R2422 B.n965 B.n964 71.676
R2423 B.n970 B.n969 71.676
R2424 B.n973 B.n972 71.676
R2425 B.n978 B.n977 71.676
R2426 B.n981 B.n980 71.676
R2427 B.n986 B.n985 71.676
R2428 B.n989 B.n988 71.676
R2429 B.n994 B.n993 71.676
R2430 B.n997 B.n996 71.676
R2431 B.n1002 B.n1001 71.676
R2432 B.n1005 B.n1004 71.676
R2433 B.n1010 B.n1009 71.676
R2434 B.n1013 B.n1012 71.676
R2435 B.n561 B.n247 71.676
R2436 B.n559 B.n249 71.676
R2437 B.n555 B.n554 71.676
R2438 B.n548 B.n251 71.676
R2439 B.n547 B.n546 71.676
R2440 B.n540 B.n253 71.676
R2441 B.n539 B.n538 71.676
R2442 B.n532 B.n255 71.676
R2443 B.n531 B.n530 71.676
R2444 B.n524 B.n257 71.676
R2445 B.n523 B.n522 71.676
R2446 B.n516 B.n259 71.676
R2447 B.n515 B.n514 71.676
R2448 B.n508 B.n261 71.676
R2449 B.n507 B.n506 71.676
R2450 B.n500 B.n263 71.676
R2451 B.n499 B.n498 71.676
R2452 B.n492 B.n265 71.676
R2453 B.n491 B.n490 71.676
R2454 B.n484 B.n267 71.676
R2455 B.n483 B.n482 71.676
R2456 B.n476 B.n269 71.676
R2457 B.n475 B.n474 71.676
R2458 B.n468 B.n271 71.676
R2459 B.n467 B.n466 71.676
R2460 B.n460 B.n273 71.676
R2461 B.n459 B.n458 71.676
R2462 B.n452 B.n275 71.676
R2463 B.n451 B.n450 71.676
R2464 B.n444 B.n277 71.676
R2465 B.n443 B.n442 71.676
R2466 B.n436 B.n282 71.676
R2467 B.n435 B.n434 71.676
R2468 B.n427 B.n284 71.676
R2469 B.n426 B.n425 71.676
R2470 B.n419 B.n288 71.676
R2471 B.n418 B.n417 71.676
R2472 B.n411 B.n290 71.676
R2473 B.n410 B.n409 71.676
R2474 B.n403 B.n292 71.676
R2475 B.n402 B.n401 71.676
R2476 B.n395 B.n294 71.676
R2477 B.n394 B.n393 71.676
R2478 B.n387 B.n296 71.676
R2479 B.n386 B.n385 71.676
R2480 B.n379 B.n298 71.676
R2481 B.n378 B.n377 71.676
R2482 B.n371 B.n300 71.676
R2483 B.n370 B.n369 71.676
R2484 B.n363 B.n302 71.676
R2485 B.n362 B.n361 71.676
R2486 B.n355 B.n304 71.676
R2487 B.n354 B.n353 71.676
R2488 B.n347 B.n306 71.676
R2489 B.n346 B.n345 71.676
R2490 B.n339 B.n308 71.676
R2491 B.n338 B.n337 71.676
R2492 B.n331 B.n310 71.676
R2493 B.n330 B.n329 71.676
R2494 B.n323 B.n312 71.676
R2495 B.n322 B.n321 71.676
R2496 B.n315 B.n314 71.676
R2497 B.n562 B.n561 71.676
R2498 B.n556 B.n249 71.676
R2499 B.n554 B.n553 71.676
R2500 B.n549 B.n548 71.676
R2501 B.n546 B.n545 71.676
R2502 B.n541 B.n540 71.676
R2503 B.n538 B.n537 71.676
R2504 B.n533 B.n532 71.676
R2505 B.n530 B.n529 71.676
R2506 B.n525 B.n524 71.676
R2507 B.n522 B.n521 71.676
R2508 B.n517 B.n516 71.676
R2509 B.n514 B.n513 71.676
R2510 B.n509 B.n508 71.676
R2511 B.n506 B.n505 71.676
R2512 B.n501 B.n500 71.676
R2513 B.n498 B.n497 71.676
R2514 B.n493 B.n492 71.676
R2515 B.n490 B.n489 71.676
R2516 B.n485 B.n484 71.676
R2517 B.n482 B.n481 71.676
R2518 B.n477 B.n476 71.676
R2519 B.n474 B.n473 71.676
R2520 B.n469 B.n468 71.676
R2521 B.n466 B.n465 71.676
R2522 B.n461 B.n460 71.676
R2523 B.n458 B.n457 71.676
R2524 B.n453 B.n452 71.676
R2525 B.n450 B.n449 71.676
R2526 B.n445 B.n444 71.676
R2527 B.n442 B.n441 71.676
R2528 B.n437 B.n436 71.676
R2529 B.n434 B.n433 71.676
R2530 B.n428 B.n427 71.676
R2531 B.n425 B.n424 71.676
R2532 B.n420 B.n419 71.676
R2533 B.n417 B.n416 71.676
R2534 B.n412 B.n411 71.676
R2535 B.n409 B.n408 71.676
R2536 B.n404 B.n403 71.676
R2537 B.n401 B.n400 71.676
R2538 B.n396 B.n395 71.676
R2539 B.n393 B.n392 71.676
R2540 B.n388 B.n387 71.676
R2541 B.n385 B.n384 71.676
R2542 B.n380 B.n379 71.676
R2543 B.n377 B.n376 71.676
R2544 B.n372 B.n371 71.676
R2545 B.n369 B.n368 71.676
R2546 B.n364 B.n363 71.676
R2547 B.n361 B.n360 71.676
R2548 B.n356 B.n355 71.676
R2549 B.n353 B.n352 71.676
R2550 B.n348 B.n347 71.676
R2551 B.n345 B.n344 71.676
R2552 B.n340 B.n339 71.676
R2553 B.n337 B.n336 71.676
R2554 B.n332 B.n331 71.676
R2555 B.n329 B.n328 71.676
R2556 B.n324 B.n323 71.676
R2557 B.n321 B.n320 71.676
R2558 B.n316 B.n315 71.676
R2559 B.n1111 B.n1110 71.676
R2560 B.n1111 B.n2 71.676
R2561 B.n118 B.n117 59.5399
R2562 B.n126 B.n125 59.5399
R2563 B.n430 B.n286 59.5399
R2564 B.n280 B.n279 59.5399
R2565 B.n567 B.n246 53.2147
R2566 B.n1018 B.n86 53.2147
R2567 B.n567 B.n242 32.6002
R2568 B.n573 B.n242 32.6002
R2569 B.n573 B.n238 32.6002
R2570 B.n579 B.n238 32.6002
R2571 B.n579 B.n234 32.6002
R2572 B.n585 B.n234 32.6002
R2573 B.n585 B.n229 32.6002
R2574 B.n591 B.n229 32.6002
R2575 B.n591 B.n230 32.6002
R2576 B.n597 B.n222 32.6002
R2577 B.n603 B.n222 32.6002
R2578 B.n603 B.n218 32.6002
R2579 B.n609 B.n218 32.6002
R2580 B.n609 B.n214 32.6002
R2581 B.n615 B.n214 32.6002
R2582 B.n615 B.n210 32.6002
R2583 B.n621 B.n210 32.6002
R2584 B.n621 B.n206 32.6002
R2585 B.n627 B.n206 32.6002
R2586 B.n627 B.n202 32.6002
R2587 B.n633 B.n202 32.6002
R2588 B.n633 B.n197 32.6002
R2589 B.n639 B.n197 32.6002
R2590 B.n639 B.n198 32.6002
R2591 B.n645 B.n190 32.6002
R2592 B.n651 B.n190 32.6002
R2593 B.n651 B.n186 32.6002
R2594 B.n657 B.n186 32.6002
R2595 B.n657 B.n182 32.6002
R2596 B.n663 B.n182 32.6002
R2597 B.n663 B.n178 32.6002
R2598 B.n669 B.n178 32.6002
R2599 B.n669 B.n174 32.6002
R2600 B.n675 B.n174 32.6002
R2601 B.n675 B.n170 32.6002
R2602 B.n681 B.n170 32.6002
R2603 B.n687 B.n166 32.6002
R2604 B.n687 B.n162 32.6002
R2605 B.n694 B.n162 32.6002
R2606 B.n694 B.n158 32.6002
R2607 B.n700 B.n158 32.6002
R2608 B.n700 B.n4 32.6002
R2609 B.n1109 B.n4 32.6002
R2610 B.n1109 B.n1108 32.6002
R2611 B.n1108 B.n1107 32.6002
R2612 B.n1107 B.n8 32.6002
R2613 B.n12 B.n8 32.6002
R2614 B.n1100 B.n12 32.6002
R2615 B.n1100 B.n1099 32.6002
R2616 B.n1099 B.n1098 32.6002
R2617 B.n1098 B.n16 32.6002
R2618 B.n1092 B.n1091 32.6002
R2619 B.n1091 B.n1090 32.6002
R2620 B.n1090 B.n23 32.6002
R2621 B.n1084 B.n23 32.6002
R2622 B.n1084 B.n1083 32.6002
R2623 B.n1083 B.n1082 32.6002
R2624 B.n1082 B.n30 32.6002
R2625 B.n1076 B.n30 32.6002
R2626 B.n1076 B.n1075 32.6002
R2627 B.n1075 B.n1074 32.6002
R2628 B.n1074 B.n37 32.6002
R2629 B.n1068 B.n37 32.6002
R2630 B.n1067 B.n1066 32.6002
R2631 B.n1066 B.n44 32.6002
R2632 B.n1060 B.n44 32.6002
R2633 B.n1060 B.n1059 32.6002
R2634 B.n1059 B.n1058 32.6002
R2635 B.n1058 B.n51 32.6002
R2636 B.n1052 B.n51 32.6002
R2637 B.n1052 B.n1051 32.6002
R2638 B.n1051 B.n1050 32.6002
R2639 B.n1050 B.n58 32.6002
R2640 B.n1044 B.n58 32.6002
R2641 B.n1044 B.n1043 32.6002
R2642 B.n1043 B.n1042 32.6002
R2643 B.n1042 B.n65 32.6002
R2644 B.n1036 B.n65 32.6002
R2645 B.n1035 B.n1034 32.6002
R2646 B.n1034 B.n72 32.6002
R2647 B.n1028 B.n72 32.6002
R2648 B.n1028 B.n1027 32.6002
R2649 B.n1027 B.n1026 32.6002
R2650 B.n1026 B.n79 32.6002
R2651 B.n1020 B.n79 32.6002
R2652 B.n1020 B.n1019 32.6002
R2653 B.n1019 B.n1018 32.6002
R2654 B.n565 B.n564 31.3761
R2655 B.n569 B.n244 31.3761
R2656 B.n766 B.n763 31.3761
R2657 B.n1016 B.n1015 31.3761
R2658 B.n230 B.t9 27.8061
R2659 B.t5 B.n1035 27.8061
R2660 B.n198 B.t1 25.8885
R2661 B.t3 B.n1067 25.8885
R2662 B B.n1112 18.0485
R2663 B.n681 B.t0 17.2592
R2664 B.n1092 B.t2 17.2592
R2665 B.t0 B.n166 15.3415
R2666 B.t2 B.n16 15.3415
R2667 B.n565 B.n240 10.6151
R2668 B.n575 B.n240 10.6151
R2669 B.n576 B.n575 10.6151
R2670 B.n577 B.n576 10.6151
R2671 B.n577 B.n232 10.6151
R2672 B.n587 B.n232 10.6151
R2673 B.n588 B.n587 10.6151
R2674 B.n589 B.n588 10.6151
R2675 B.n589 B.n224 10.6151
R2676 B.n599 B.n224 10.6151
R2677 B.n600 B.n599 10.6151
R2678 B.n601 B.n600 10.6151
R2679 B.n601 B.n216 10.6151
R2680 B.n611 B.n216 10.6151
R2681 B.n612 B.n611 10.6151
R2682 B.n613 B.n612 10.6151
R2683 B.n613 B.n208 10.6151
R2684 B.n623 B.n208 10.6151
R2685 B.n624 B.n623 10.6151
R2686 B.n625 B.n624 10.6151
R2687 B.n625 B.n200 10.6151
R2688 B.n635 B.n200 10.6151
R2689 B.n636 B.n635 10.6151
R2690 B.n637 B.n636 10.6151
R2691 B.n637 B.n192 10.6151
R2692 B.n647 B.n192 10.6151
R2693 B.n648 B.n647 10.6151
R2694 B.n649 B.n648 10.6151
R2695 B.n649 B.n184 10.6151
R2696 B.n659 B.n184 10.6151
R2697 B.n660 B.n659 10.6151
R2698 B.n661 B.n660 10.6151
R2699 B.n661 B.n176 10.6151
R2700 B.n671 B.n176 10.6151
R2701 B.n672 B.n671 10.6151
R2702 B.n673 B.n672 10.6151
R2703 B.n673 B.n168 10.6151
R2704 B.n683 B.n168 10.6151
R2705 B.n684 B.n683 10.6151
R2706 B.n685 B.n684 10.6151
R2707 B.n685 B.n160 10.6151
R2708 B.n696 B.n160 10.6151
R2709 B.n697 B.n696 10.6151
R2710 B.n698 B.n697 10.6151
R2711 B.n698 B.n0 10.6151
R2712 B.n564 B.n563 10.6151
R2713 B.n563 B.n248 10.6151
R2714 B.n558 B.n248 10.6151
R2715 B.n558 B.n557 10.6151
R2716 B.n557 B.n250 10.6151
R2717 B.n552 B.n250 10.6151
R2718 B.n552 B.n551 10.6151
R2719 B.n551 B.n550 10.6151
R2720 B.n550 B.n252 10.6151
R2721 B.n544 B.n252 10.6151
R2722 B.n544 B.n543 10.6151
R2723 B.n543 B.n542 10.6151
R2724 B.n542 B.n254 10.6151
R2725 B.n536 B.n254 10.6151
R2726 B.n536 B.n535 10.6151
R2727 B.n535 B.n534 10.6151
R2728 B.n534 B.n256 10.6151
R2729 B.n528 B.n256 10.6151
R2730 B.n528 B.n527 10.6151
R2731 B.n527 B.n526 10.6151
R2732 B.n526 B.n258 10.6151
R2733 B.n520 B.n258 10.6151
R2734 B.n520 B.n519 10.6151
R2735 B.n519 B.n518 10.6151
R2736 B.n518 B.n260 10.6151
R2737 B.n512 B.n260 10.6151
R2738 B.n512 B.n511 10.6151
R2739 B.n511 B.n510 10.6151
R2740 B.n510 B.n262 10.6151
R2741 B.n504 B.n262 10.6151
R2742 B.n504 B.n503 10.6151
R2743 B.n503 B.n502 10.6151
R2744 B.n502 B.n264 10.6151
R2745 B.n496 B.n264 10.6151
R2746 B.n496 B.n495 10.6151
R2747 B.n495 B.n494 10.6151
R2748 B.n494 B.n266 10.6151
R2749 B.n488 B.n266 10.6151
R2750 B.n488 B.n487 10.6151
R2751 B.n487 B.n486 10.6151
R2752 B.n486 B.n268 10.6151
R2753 B.n480 B.n268 10.6151
R2754 B.n480 B.n479 10.6151
R2755 B.n479 B.n478 10.6151
R2756 B.n478 B.n270 10.6151
R2757 B.n472 B.n270 10.6151
R2758 B.n472 B.n471 10.6151
R2759 B.n471 B.n470 10.6151
R2760 B.n470 B.n272 10.6151
R2761 B.n464 B.n272 10.6151
R2762 B.n464 B.n463 10.6151
R2763 B.n463 B.n462 10.6151
R2764 B.n462 B.n274 10.6151
R2765 B.n456 B.n274 10.6151
R2766 B.n456 B.n455 10.6151
R2767 B.n455 B.n454 10.6151
R2768 B.n454 B.n276 10.6151
R2769 B.n448 B.n447 10.6151
R2770 B.n447 B.n446 10.6151
R2771 B.n446 B.n281 10.6151
R2772 B.n440 B.n281 10.6151
R2773 B.n440 B.n439 10.6151
R2774 B.n439 B.n438 10.6151
R2775 B.n438 B.n283 10.6151
R2776 B.n432 B.n283 10.6151
R2777 B.n432 B.n431 10.6151
R2778 B.n429 B.n287 10.6151
R2779 B.n423 B.n287 10.6151
R2780 B.n423 B.n422 10.6151
R2781 B.n422 B.n421 10.6151
R2782 B.n421 B.n289 10.6151
R2783 B.n415 B.n289 10.6151
R2784 B.n415 B.n414 10.6151
R2785 B.n414 B.n413 10.6151
R2786 B.n413 B.n291 10.6151
R2787 B.n407 B.n291 10.6151
R2788 B.n407 B.n406 10.6151
R2789 B.n406 B.n405 10.6151
R2790 B.n405 B.n293 10.6151
R2791 B.n399 B.n293 10.6151
R2792 B.n399 B.n398 10.6151
R2793 B.n398 B.n397 10.6151
R2794 B.n397 B.n295 10.6151
R2795 B.n391 B.n295 10.6151
R2796 B.n391 B.n390 10.6151
R2797 B.n390 B.n389 10.6151
R2798 B.n389 B.n297 10.6151
R2799 B.n383 B.n297 10.6151
R2800 B.n383 B.n382 10.6151
R2801 B.n382 B.n381 10.6151
R2802 B.n381 B.n299 10.6151
R2803 B.n375 B.n299 10.6151
R2804 B.n375 B.n374 10.6151
R2805 B.n374 B.n373 10.6151
R2806 B.n373 B.n301 10.6151
R2807 B.n367 B.n301 10.6151
R2808 B.n367 B.n366 10.6151
R2809 B.n366 B.n365 10.6151
R2810 B.n365 B.n303 10.6151
R2811 B.n359 B.n303 10.6151
R2812 B.n359 B.n358 10.6151
R2813 B.n358 B.n357 10.6151
R2814 B.n357 B.n305 10.6151
R2815 B.n351 B.n305 10.6151
R2816 B.n351 B.n350 10.6151
R2817 B.n350 B.n349 10.6151
R2818 B.n349 B.n307 10.6151
R2819 B.n343 B.n307 10.6151
R2820 B.n343 B.n342 10.6151
R2821 B.n342 B.n341 10.6151
R2822 B.n341 B.n309 10.6151
R2823 B.n335 B.n309 10.6151
R2824 B.n335 B.n334 10.6151
R2825 B.n334 B.n333 10.6151
R2826 B.n333 B.n311 10.6151
R2827 B.n327 B.n311 10.6151
R2828 B.n327 B.n326 10.6151
R2829 B.n326 B.n325 10.6151
R2830 B.n325 B.n313 10.6151
R2831 B.n319 B.n313 10.6151
R2832 B.n319 B.n318 10.6151
R2833 B.n318 B.n317 10.6151
R2834 B.n317 B.n244 10.6151
R2835 B.n570 B.n569 10.6151
R2836 B.n571 B.n570 10.6151
R2837 B.n571 B.n236 10.6151
R2838 B.n581 B.n236 10.6151
R2839 B.n582 B.n581 10.6151
R2840 B.n583 B.n582 10.6151
R2841 B.n583 B.n227 10.6151
R2842 B.n593 B.n227 10.6151
R2843 B.n594 B.n593 10.6151
R2844 B.n595 B.n594 10.6151
R2845 B.n595 B.n220 10.6151
R2846 B.n605 B.n220 10.6151
R2847 B.n606 B.n605 10.6151
R2848 B.n607 B.n606 10.6151
R2849 B.n607 B.n212 10.6151
R2850 B.n617 B.n212 10.6151
R2851 B.n618 B.n617 10.6151
R2852 B.n619 B.n618 10.6151
R2853 B.n619 B.n204 10.6151
R2854 B.n629 B.n204 10.6151
R2855 B.n630 B.n629 10.6151
R2856 B.n631 B.n630 10.6151
R2857 B.n631 B.n195 10.6151
R2858 B.n641 B.n195 10.6151
R2859 B.n642 B.n641 10.6151
R2860 B.n643 B.n642 10.6151
R2861 B.n643 B.n188 10.6151
R2862 B.n653 B.n188 10.6151
R2863 B.n654 B.n653 10.6151
R2864 B.n655 B.n654 10.6151
R2865 B.n655 B.n180 10.6151
R2866 B.n665 B.n180 10.6151
R2867 B.n666 B.n665 10.6151
R2868 B.n667 B.n666 10.6151
R2869 B.n667 B.n172 10.6151
R2870 B.n677 B.n172 10.6151
R2871 B.n678 B.n677 10.6151
R2872 B.n679 B.n678 10.6151
R2873 B.n679 B.n164 10.6151
R2874 B.n689 B.n164 10.6151
R2875 B.n690 B.n689 10.6151
R2876 B.n692 B.n690 10.6151
R2877 B.n692 B.n691 10.6151
R2878 B.n691 B.n156 10.6151
R2879 B.n703 B.n156 10.6151
R2880 B.n704 B.n703 10.6151
R2881 B.n705 B.n704 10.6151
R2882 B.n706 B.n705 10.6151
R2883 B.n707 B.n706 10.6151
R2884 B.n710 B.n707 10.6151
R2885 B.n711 B.n710 10.6151
R2886 B.n712 B.n711 10.6151
R2887 B.n713 B.n712 10.6151
R2888 B.n715 B.n713 10.6151
R2889 B.n716 B.n715 10.6151
R2890 B.n717 B.n716 10.6151
R2891 B.n718 B.n717 10.6151
R2892 B.n720 B.n718 10.6151
R2893 B.n721 B.n720 10.6151
R2894 B.n722 B.n721 10.6151
R2895 B.n723 B.n722 10.6151
R2896 B.n725 B.n723 10.6151
R2897 B.n726 B.n725 10.6151
R2898 B.n727 B.n726 10.6151
R2899 B.n728 B.n727 10.6151
R2900 B.n730 B.n728 10.6151
R2901 B.n731 B.n730 10.6151
R2902 B.n732 B.n731 10.6151
R2903 B.n733 B.n732 10.6151
R2904 B.n735 B.n733 10.6151
R2905 B.n736 B.n735 10.6151
R2906 B.n737 B.n736 10.6151
R2907 B.n738 B.n737 10.6151
R2908 B.n740 B.n738 10.6151
R2909 B.n741 B.n740 10.6151
R2910 B.n742 B.n741 10.6151
R2911 B.n743 B.n742 10.6151
R2912 B.n745 B.n743 10.6151
R2913 B.n746 B.n745 10.6151
R2914 B.n747 B.n746 10.6151
R2915 B.n748 B.n747 10.6151
R2916 B.n750 B.n748 10.6151
R2917 B.n751 B.n750 10.6151
R2918 B.n752 B.n751 10.6151
R2919 B.n753 B.n752 10.6151
R2920 B.n755 B.n753 10.6151
R2921 B.n756 B.n755 10.6151
R2922 B.n757 B.n756 10.6151
R2923 B.n758 B.n757 10.6151
R2924 B.n760 B.n758 10.6151
R2925 B.n761 B.n760 10.6151
R2926 B.n762 B.n761 10.6151
R2927 B.n763 B.n762 10.6151
R2928 B.n1104 B.n1 10.6151
R2929 B.n1104 B.n1103 10.6151
R2930 B.n1103 B.n1102 10.6151
R2931 B.n1102 B.n10 10.6151
R2932 B.n1096 B.n10 10.6151
R2933 B.n1096 B.n1095 10.6151
R2934 B.n1095 B.n1094 10.6151
R2935 B.n1094 B.n18 10.6151
R2936 B.n1088 B.n18 10.6151
R2937 B.n1088 B.n1087 10.6151
R2938 B.n1087 B.n1086 10.6151
R2939 B.n1086 B.n25 10.6151
R2940 B.n1080 B.n25 10.6151
R2941 B.n1080 B.n1079 10.6151
R2942 B.n1079 B.n1078 10.6151
R2943 B.n1078 B.n32 10.6151
R2944 B.n1072 B.n32 10.6151
R2945 B.n1072 B.n1071 10.6151
R2946 B.n1071 B.n1070 10.6151
R2947 B.n1070 B.n39 10.6151
R2948 B.n1064 B.n39 10.6151
R2949 B.n1064 B.n1063 10.6151
R2950 B.n1063 B.n1062 10.6151
R2951 B.n1062 B.n46 10.6151
R2952 B.n1056 B.n46 10.6151
R2953 B.n1056 B.n1055 10.6151
R2954 B.n1055 B.n1054 10.6151
R2955 B.n1054 B.n53 10.6151
R2956 B.n1048 B.n53 10.6151
R2957 B.n1048 B.n1047 10.6151
R2958 B.n1047 B.n1046 10.6151
R2959 B.n1046 B.n60 10.6151
R2960 B.n1040 B.n60 10.6151
R2961 B.n1040 B.n1039 10.6151
R2962 B.n1039 B.n1038 10.6151
R2963 B.n1038 B.n67 10.6151
R2964 B.n1032 B.n67 10.6151
R2965 B.n1032 B.n1031 10.6151
R2966 B.n1031 B.n1030 10.6151
R2967 B.n1030 B.n74 10.6151
R2968 B.n1024 B.n74 10.6151
R2969 B.n1024 B.n1023 10.6151
R2970 B.n1023 B.n1022 10.6151
R2971 B.n1022 B.n81 10.6151
R2972 B.n1016 B.n81 10.6151
R2973 B.n1015 B.n1014 10.6151
R2974 B.n1014 B.n88 10.6151
R2975 B.n1008 B.n88 10.6151
R2976 B.n1008 B.n1007 10.6151
R2977 B.n1007 B.n1006 10.6151
R2978 B.n1006 B.n90 10.6151
R2979 B.n1000 B.n90 10.6151
R2980 B.n1000 B.n999 10.6151
R2981 B.n999 B.n998 10.6151
R2982 B.n998 B.n92 10.6151
R2983 B.n992 B.n92 10.6151
R2984 B.n992 B.n991 10.6151
R2985 B.n991 B.n990 10.6151
R2986 B.n990 B.n94 10.6151
R2987 B.n984 B.n94 10.6151
R2988 B.n984 B.n983 10.6151
R2989 B.n983 B.n982 10.6151
R2990 B.n982 B.n96 10.6151
R2991 B.n976 B.n96 10.6151
R2992 B.n976 B.n975 10.6151
R2993 B.n975 B.n974 10.6151
R2994 B.n974 B.n98 10.6151
R2995 B.n968 B.n98 10.6151
R2996 B.n968 B.n967 10.6151
R2997 B.n967 B.n966 10.6151
R2998 B.n966 B.n100 10.6151
R2999 B.n960 B.n100 10.6151
R3000 B.n960 B.n959 10.6151
R3001 B.n959 B.n958 10.6151
R3002 B.n958 B.n102 10.6151
R3003 B.n952 B.n102 10.6151
R3004 B.n952 B.n951 10.6151
R3005 B.n951 B.n950 10.6151
R3006 B.n950 B.n104 10.6151
R3007 B.n944 B.n104 10.6151
R3008 B.n944 B.n943 10.6151
R3009 B.n943 B.n942 10.6151
R3010 B.n942 B.n106 10.6151
R3011 B.n936 B.n106 10.6151
R3012 B.n936 B.n935 10.6151
R3013 B.n935 B.n934 10.6151
R3014 B.n934 B.n108 10.6151
R3015 B.n928 B.n108 10.6151
R3016 B.n928 B.n927 10.6151
R3017 B.n927 B.n926 10.6151
R3018 B.n926 B.n110 10.6151
R3019 B.n920 B.n110 10.6151
R3020 B.n920 B.n919 10.6151
R3021 B.n919 B.n918 10.6151
R3022 B.n918 B.n112 10.6151
R3023 B.n912 B.n112 10.6151
R3024 B.n912 B.n911 10.6151
R3025 B.n911 B.n910 10.6151
R3026 B.n910 B.n114 10.6151
R3027 B.n904 B.n114 10.6151
R3028 B.n904 B.n903 10.6151
R3029 B.n903 B.n902 10.6151
R3030 B.n898 B.n897 10.6151
R3031 B.n897 B.n120 10.6151
R3032 B.n892 B.n120 10.6151
R3033 B.n892 B.n891 10.6151
R3034 B.n891 B.n890 10.6151
R3035 B.n890 B.n122 10.6151
R3036 B.n884 B.n122 10.6151
R3037 B.n884 B.n883 10.6151
R3038 B.n883 B.n882 10.6151
R3039 B.n878 B.n877 10.6151
R3040 B.n877 B.n128 10.6151
R3041 B.n872 B.n128 10.6151
R3042 B.n872 B.n871 10.6151
R3043 B.n871 B.n870 10.6151
R3044 B.n870 B.n130 10.6151
R3045 B.n864 B.n130 10.6151
R3046 B.n864 B.n863 10.6151
R3047 B.n863 B.n862 10.6151
R3048 B.n862 B.n132 10.6151
R3049 B.n856 B.n132 10.6151
R3050 B.n856 B.n855 10.6151
R3051 B.n855 B.n854 10.6151
R3052 B.n854 B.n134 10.6151
R3053 B.n848 B.n134 10.6151
R3054 B.n848 B.n847 10.6151
R3055 B.n847 B.n846 10.6151
R3056 B.n846 B.n136 10.6151
R3057 B.n840 B.n136 10.6151
R3058 B.n840 B.n839 10.6151
R3059 B.n839 B.n838 10.6151
R3060 B.n838 B.n138 10.6151
R3061 B.n832 B.n138 10.6151
R3062 B.n832 B.n831 10.6151
R3063 B.n831 B.n830 10.6151
R3064 B.n830 B.n140 10.6151
R3065 B.n824 B.n140 10.6151
R3066 B.n824 B.n823 10.6151
R3067 B.n823 B.n822 10.6151
R3068 B.n822 B.n142 10.6151
R3069 B.n816 B.n142 10.6151
R3070 B.n816 B.n815 10.6151
R3071 B.n815 B.n814 10.6151
R3072 B.n814 B.n144 10.6151
R3073 B.n808 B.n144 10.6151
R3074 B.n808 B.n807 10.6151
R3075 B.n807 B.n806 10.6151
R3076 B.n806 B.n146 10.6151
R3077 B.n800 B.n146 10.6151
R3078 B.n800 B.n799 10.6151
R3079 B.n799 B.n798 10.6151
R3080 B.n798 B.n148 10.6151
R3081 B.n792 B.n148 10.6151
R3082 B.n792 B.n791 10.6151
R3083 B.n791 B.n790 10.6151
R3084 B.n790 B.n150 10.6151
R3085 B.n784 B.n150 10.6151
R3086 B.n784 B.n783 10.6151
R3087 B.n783 B.n782 10.6151
R3088 B.n782 B.n152 10.6151
R3089 B.n776 B.n152 10.6151
R3090 B.n776 B.n775 10.6151
R3091 B.n775 B.n774 10.6151
R3092 B.n774 B.n154 10.6151
R3093 B.n768 B.n154 10.6151
R3094 B.n768 B.n767 10.6151
R3095 B.n767 B.n766 10.6151
R3096 B.n280 B.n276 9.36635
R3097 B.n430 B.n429 9.36635
R3098 B.n902 B.n118 9.36635
R3099 B.n878 B.n126 9.36635
R3100 B.n1112 B.n0 8.11757
R3101 B.n1112 B.n1 8.11757
R3102 B.n645 B.t1 6.7122
R3103 B.n1068 B.t3 6.7122
R3104 B.n597 B.t9 4.79457
R3105 B.n1036 B.t5 4.79457
R3106 B.n448 B.n280 1.24928
R3107 B.n431 B.n430 1.24928
R3108 B.n898 B.n118 1.24928
R3109 B.n882 B.n126 1.24928
R3110 VN.n0 VN.t1 140.243
R3111 VN.n1 VN.t2 140.243
R3112 VN.n0 VN.t3 138.797
R3113 VN.n1 VN.t0 138.797
R3114 VN VN.n1 56.7939
R3115 VN VN.n0 1.72194
R3116 VDD2.n2 VDD2.n0 113.737
R3117 VDD2.n2 VDD2.n1 63.5911
R3118 VDD2.n1 VDD2.t3 1.12104
R3119 VDD2.n1 VDD2.t1 1.12104
R3120 VDD2.n0 VDD2.t2 1.12104
R3121 VDD2.n0 VDD2.t0 1.12104
R3122 VDD2 VDD2.n2 0.0586897
C0 VDD1 VDD2 1.37192f
C1 VP VN 8.252191f
C2 VP VTAIL 7.1602f
C3 VN VTAIL 7.14609f
C4 VP VDD1 7.63071f
C5 VP VDD2 0.483549f
C6 VDD1 VN 0.150424f
C7 VDD2 VN 7.29868f
C8 VDD1 VTAIL 6.98678f
C9 VDD2 VTAIL 7.05037f
C10 VDD2 B 4.994799f
C11 VDD1 B 10.20857f
C12 VTAIL B 14.29391f
C13 VN B 13.854899f
C14 VP B 12.311513f
C15 VDD2.t2 B 0.376095f
C16 VDD2.t0 B 0.376095f
C17 VDD2.n0 B 4.38014f
C18 VDD2.t3 B 0.376095f
C19 VDD2.t1 B 0.376095f
C20 VDD2.n1 B 3.4271f
C21 VDD2.n2 B 4.75862f
C22 VN.t1 B 3.83243f
C23 VN.t3 B 3.81905f
C24 VN.n0 B 2.31341f
C25 VN.t2 B 3.83243f
C26 VN.t0 B 3.81905f
C27 VN.n1 B 3.65083f
C28 VDD1.t2 B 0.378702f
C29 VDD1.t0 B 0.378702f
C30 VDD1.n0 B 3.45137f
C31 VDD1.t1 B 0.378702f
C32 VDD1.t3 B 0.378702f
C33 VDD1.n1 B 4.4395f
C34 VTAIL.n0 B 0.023636f
C35 VTAIL.n1 B 0.015972f
C36 VTAIL.n2 B 0.008583f
C37 VTAIL.n3 B 0.020286f
C38 VTAIL.n4 B 0.009088f
C39 VTAIL.n5 B 0.015972f
C40 VTAIL.n6 B 0.008583f
C41 VTAIL.n7 B 0.020286f
C42 VTAIL.n8 B 0.008835f
C43 VTAIL.n9 B 0.015972f
C44 VTAIL.n10 B 0.009088f
C45 VTAIL.n11 B 0.020286f
C46 VTAIL.n12 B 0.009088f
C47 VTAIL.n13 B 0.015972f
C48 VTAIL.n14 B 0.008583f
C49 VTAIL.n15 B 0.020286f
C50 VTAIL.n16 B 0.009088f
C51 VTAIL.n17 B 0.015972f
C52 VTAIL.n18 B 0.008583f
C53 VTAIL.n19 B 0.020286f
C54 VTAIL.n20 B 0.009088f
C55 VTAIL.n21 B 0.015972f
C56 VTAIL.n22 B 0.008583f
C57 VTAIL.n23 B 0.020286f
C58 VTAIL.n24 B 0.009088f
C59 VTAIL.n25 B 0.015972f
C60 VTAIL.n26 B 0.008583f
C61 VTAIL.n27 B 0.020286f
C62 VTAIL.n28 B 0.009088f
C63 VTAIL.n29 B 1.23461f
C64 VTAIL.n30 B 0.008583f
C65 VTAIL.t2 B 0.033596f
C66 VTAIL.n31 B 0.114865f
C67 VTAIL.n32 B 0.011984f
C68 VTAIL.n33 B 0.015215f
C69 VTAIL.n34 B 0.020286f
C70 VTAIL.n35 B 0.009088f
C71 VTAIL.n36 B 0.008583f
C72 VTAIL.n37 B 0.015972f
C73 VTAIL.n38 B 0.015972f
C74 VTAIL.n39 B 0.008583f
C75 VTAIL.n40 B 0.009088f
C76 VTAIL.n41 B 0.020286f
C77 VTAIL.n42 B 0.020286f
C78 VTAIL.n43 B 0.009088f
C79 VTAIL.n44 B 0.008583f
C80 VTAIL.n45 B 0.015972f
C81 VTAIL.n46 B 0.015972f
C82 VTAIL.n47 B 0.008583f
C83 VTAIL.n48 B 0.009088f
C84 VTAIL.n49 B 0.020286f
C85 VTAIL.n50 B 0.020286f
C86 VTAIL.n51 B 0.009088f
C87 VTAIL.n52 B 0.008583f
C88 VTAIL.n53 B 0.015972f
C89 VTAIL.n54 B 0.015972f
C90 VTAIL.n55 B 0.008583f
C91 VTAIL.n56 B 0.009088f
C92 VTAIL.n57 B 0.020286f
C93 VTAIL.n58 B 0.020286f
C94 VTAIL.n59 B 0.009088f
C95 VTAIL.n60 B 0.008583f
C96 VTAIL.n61 B 0.015972f
C97 VTAIL.n62 B 0.015972f
C98 VTAIL.n63 B 0.008583f
C99 VTAIL.n64 B 0.009088f
C100 VTAIL.n65 B 0.020286f
C101 VTAIL.n66 B 0.020286f
C102 VTAIL.n67 B 0.009088f
C103 VTAIL.n68 B 0.008583f
C104 VTAIL.n69 B 0.015972f
C105 VTAIL.n70 B 0.015972f
C106 VTAIL.n71 B 0.008583f
C107 VTAIL.n72 B 0.008583f
C108 VTAIL.n73 B 0.009088f
C109 VTAIL.n74 B 0.020286f
C110 VTAIL.n75 B 0.020286f
C111 VTAIL.n76 B 0.020286f
C112 VTAIL.n77 B 0.008835f
C113 VTAIL.n78 B 0.008583f
C114 VTAIL.n79 B 0.015972f
C115 VTAIL.n80 B 0.015972f
C116 VTAIL.n81 B 0.008583f
C117 VTAIL.n82 B 0.009088f
C118 VTAIL.n83 B 0.020286f
C119 VTAIL.n84 B 0.020286f
C120 VTAIL.n85 B 0.009088f
C121 VTAIL.n86 B 0.008583f
C122 VTAIL.n87 B 0.015972f
C123 VTAIL.n88 B 0.015972f
C124 VTAIL.n89 B 0.008583f
C125 VTAIL.n90 B 0.009088f
C126 VTAIL.n91 B 0.020286f
C127 VTAIL.n92 B 0.046013f
C128 VTAIL.n93 B 0.009088f
C129 VTAIL.n94 B 0.008583f
C130 VTAIL.n95 B 0.040192f
C131 VTAIL.n96 B 0.026058f
C132 VTAIL.n97 B 0.138721f
C133 VTAIL.n98 B 0.023636f
C134 VTAIL.n99 B 0.015972f
C135 VTAIL.n100 B 0.008583f
C136 VTAIL.n101 B 0.020286f
C137 VTAIL.n102 B 0.009088f
C138 VTAIL.n103 B 0.015972f
C139 VTAIL.n104 B 0.008583f
C140 VTAIL.n105 B 0.020286f
C141 VTAIL.n106 B 0.008835f
C142 VTAIL.n107 B 0.015972f
C143 VTAIL.n108 B 0.009088f
C144 VTAIL.n109 B 0.020286f
C145 VTAIL.n110 B 0.009088f
C146 VTAIL.n111 B 0.015972f
C147 VTAIL.n112 B 0.008583f
C148 VTAIL.n113 B 0.020286f
C149 VTAIL.n114 B 0.009088f
C150 VTAIL.n115 B 0.015972f
C151 VTAIL.n116 B 0.008583f
C152 VTAIL.n117 B 0.020286f
C153 VTAIL.n118 B 0.009088f
C154 VTAIL.n119 B 0.015972f
C155 VTAIL.n120 B 0.008583f
C156 VTAIL.n121 B 0.020286f
C157 VTAIL.n122 B 0.009088f
C158 VTAIL.n123 B 0.015972f
C159 VTAIL.n124 B 0.008583f
C160 VTAIL.n125 B 0.020286f
C161 VTAIL.n126 B 0.009088f
C162 VTAIL.n127 B 1.23461f
C163 VTAIL.n128 B 0.008583f
C164 VTAIL.t6 B 0.033596f
C165 VTAIL.n129 B 0.114865f
C166 VTAIL.n130 B 0.011984f
C167 VTAIL.n131 B 0.015215f
C168 VTAIL.n132 B 0.020286f
C169 VTAIL.n133 B 0.009088f
C170 VTAIL.n134 B 0.008583f
C171 VTAIL.n135 B 0.015972f
C172 VTAIL.n136 B 0.015972f
C173 VTAIL.n137 B 0.008583f
C174 VTAIL.n138 B 0.009088f
C175 VTAIL.n139 B 0.020286f
C176 VTAIL.n140 B 0.020286f
C177 VTAIL.n141 B 0.009088f
C178 VTAIL.n142 B 0.008583f
C179 VTAIL.n143 B 0.015972f
C180 VTAIL.n144 B 0.015972f
C181 VTAIL.n145 B 0.008583f
C182 VTAIL.n146 B 0.009088f
C183 VTAIL.n147 B 0.020286f
C184 VTAIL.n148 B 0.020286f
C185 VTAIL.n149 B 0.009088f
C186 VTAIL.n150 B 0.008583f
C187 VTAIL.n151 B 0.015972f
C188 VTAIL.n152 B 0.015972f
C189 VTAIL.n153 B 0.008583f
C190 VTAIL.n154 B 0.009088f
C191 VTAIL.n155 B 0.020286f
C192 VTAIL.n156 B 0.020286f
C193 VTAIL.n157 B 0.009088f
C194 VTAIL.n158 B 0.008583f
C195 VTAIL.n159 B 0.015972f
C196 VTAIL.n160 B 0.015972f
C197 VTAIL.n161 B 0.008583f
C198 VTAIL.n162 B 0.009088f
C199 VTAIL.n163 B 0.020286f
C200 VTAIL.n164 B 0.020286f
C201 VTAIL.n165 B 0.009088f
C202 VTAIL.n166 B 0.008583f
C203 VTAIL.n167 B 0.015972f
C204 VTAIL.n168 B 0.015972f
C205 VTAIL.n169 B 0.008583f
C206 VTAIL.n170 B 0.008583f
C207 VTAIL.n171 B 0.009088f
C208 VTAIL.n172 B 0.020286f
C209 VTAIL.n173 B 0.020286f
C210 VTAIL.n174 B 0.020286f
C211 VTAIL.n175 B 0.008835f
C212 VTAIL.n176 B 0.008583f
C213 VTAIL.n177 B 0.015972f
C214 VTAIL.n178 B 0.015972f
C215 VTAIL.n179 B 0.008583f
C216 VTAIL.n180 B 0.009088f
C217 VTAIL.n181 B 0.020286f
C218 VTAIL.n182 B 0.020286f
C219 VTAIL.n183 B 0.009088f
C220 VTAIL.n184 B 0.008583f
C221 VTAIL.n185 B 0.015972f
C222 VTAIL.n186 B 0.015972f
C223 VTAIL.n187 B 0.008583f
C224 VTAIL.n188 B 0.009088f
C225 VTAIL.n189 B 0.020286f
C226 VTAIL.n190 B 0.046013f
C227 VTAIL.n191 B 0.009088f
C228 VTAIL.n192 B 0.008583f
C229 VTAIL.n193 B 0.040192f
C230 VTAIL.n194 B 0.026058f
C231 VTAIL.n195 B 0.231781f
C232 VTAIL.n196 B 0.023636f
C233 VTAIL.n197 B 0.015972f
C234 VTAIL.n198 B 0.008583f
C235 VTAIL.n199 B 0.020286f
C236 VTAIL.n200 B 0.009088f
C237 VTAIL.n201 B 0.015972f
C238 VTAIL.n202 B 0.008583f
C239 VTAIL.n203 B 0.020286f
C240 VTAIL.n204 B 0.008835f
C241 VTAIL.n205 B 0.015972f
C242 VTAIL.n206 B 0.009088f
C243 VTAIL.n207 B 0.020286f
C244 VTAIL.n208 B 0.009088f
C245 VTAIL.n209 B 0.015972f
C246 VTAIL.n210 B 0.008583f
C247 VTAIL.n211 B 0.020286f
C248 VTAIL.n212 B 0.009088f
C249 VTAIL.n213 B 0.015972f
C250 VTAIL.n214 B 0.008583f
C251 VTAIL.n215 B 0.020286f
C252 VTAIL.n216 B 0.009088f
C253 VTAIL.n217 B 0.015972f
C254 VTAIL.n218 B 0.008583f
C255 VTAIL.n219 B 0.020286f
C256 VTAIL.n220 B 0.009088f
C257 VTAIL.n221 B 0.015972f
C258 VTAIL.n222 B 0.008583f
C259 VTAIL.n223 B 0.020286f
C260 VTAIL.n224 B 0.009088f
C261 VTAIL.n225 B 1.23461f
C262 VTAIL.n226 B 0.008583f
C263 VTAIL.t4 B 0.033596f
C264 VTAIL.n227 B 0.114865f
C265 VTAIL.n228 B 0.011984f
C266 VTAIL.n229 B 0.015215f
C267 VTAIL.n230 B 0.020286f
C268 VTAIL.n231 B 0.009088f
C269 VTAIL.n232 B 0.008583f
C270 VTAIL.n233 B 0.015972f
C271 VTAIL.n234 B 0.015972f
C272 VTAIL.n235 B 0.008583f
C273 VTAIL.n236 B 0.009088f
C274 VTAIL.n237 B 0.020286f
C275 VTAIL.n238 B 0.020286f
C276 VTAIL.n239 B 0.009088f
C277 VTAIL.n240 B 0.008583f
C278 VTAIL.n241 B 0.015972f
C279 VTAIL.n242 B 0.015972f
C280 VTAIL.n243 B 0.008583f
C281 VTAIL.n244 B 0.009088f
C282 VTAIL.n245 B 0.020286f
C283 VTAIL.n246 B 0.020286f
C284 VTAIL.n247 B 0.009088f
C285 VTAIL.n248 B 0.008583f
C286 VTAIL.n249 B 0.015972f
C287 VTAIL.n250 B 0.015972f
C288 VTAIL.n251 B 0.008583f
C289 VTAIL.n252 B 0.009088f
C290 VTAIL.n253 B 0.020286f
C291 VTAIL.n254 B 0.020286f
C292 VTAIL.n255 B 0.009088f
C293 VTAIL.n256 B 0.008583f
C294 VTAIL.n257 B 0.015972f
C295 VTAIL.n258 B 0.015972f
C296 VTAIL.n259 B 0.008583f
C297 VTAIL.n260 B 0.009088f
C298 VTAIL.n261 B 0.020286f
C299 VTAIL.n262 B 0.020286f
C300 VTAIL.n263 B 0.009088f
C301 VTAIL.n264 B 0.008583f
C302 VTAIL.n265 B 0.015972f
C303 VTAIL.n266 B 0.015972f
C304 VTAIL.n267 B 0.008583f
C305 VTAIL.n268 B 0.008583f
C306 VTAIL.n269 B 0.009088f
C307 VTAIL.n270 B 0.020286f
C308 VTAIL.n271 B 0.020286f
C309 VTAIL.n272 B 0.020286f
C310 VTAIL.n273 B 0.008835f
C311 VTAIL.n274 B 0.008583f
C312 VTAIL.n275 B 0.015972f
C313 VTAIL.n276 B 0.015972f
C314 VTAIL.n277 B 0.008583f
C315 VTAIL.n278 B 0.009088f
C316 VTAIL.n279 B 0.020286f
C317 VTAIL.n280 B 0.020286f
C318 VTAIL.n281 B 0.009088f
C319 VTAIL.n282 B 0.008583f
C320 VTAIL.n283 B 0.015972f
C321 VTAIL.n284 B 0.015972f
C322 VTAIL.n285 B 0.008583f
C323 VTAIL.n286 B 0.009088f
C324 VTAIL.n287 B 0.020286f
C325 VTAIL.n288 B 0.046013f
C326 VTAIL.n289 B 0.009088f
C327 VTAIL.n290 B 0.008583f
C328 VTAIL.n291 B 0.040192f
C329 VTAIL.n292 B 0.026058f
C330 VTAIL.n293 B 1.40063f
C331 VTAIL.n294 B 0.023636f
C332 VTAIL.n295 B 0.015972f
C333 VTAIL.n296 B 0.008583f
C334 VTAIL.n297 B 0.020286f
C335 VTAIL.n298 B 0.009088f
C336 VTAIL.n299 B 0.015972f
C337 VTAIL.n300 B 0.008583f
C338 VTAIL.n301 B 0.020286f
C339 VTAIL.n302 B 0.008835f
C340 VTAIL.n303 B 0.015972f
C341 VTAIL.n304 B 0.008835f
C342 VTAIL.n305 B 0.008583f
C343 VTAIL.n306 B 0.020286f
C344 VTAIL.n307 B 0.020286f
C345 VTAIL.n308 B 0.009088f
C346 VTAIL.n309 B 0.015972f
C347 VTAIL.n310 B 0.008583f
C348 VTAIL.n311 B 0.020286f
C349 VTAIL.n312 B 0.009088f
C350 VTAIL.n313 B 0.015972f
C351 VTAIL.n314 B 0.008583f
C352 VTAIL.n315 B 0.020286f
C353 VTAIL.n316 B 0.009088f
C354 VTAIL.n317 B 0.015972f
C355 VTAIL.n318 B 0.008583f
C356 VTAIL.n319 B 0.020286f
C357 VTAIL.n320 B 0.009088f
C358 VTAIL.n321 B 0.015972f
C359 VTAIL.n322 B 0.008583f
C360 VTAIL.n323 B 0.020286f
C361 VTAIL.n324 B 0.009088f
C362 VTAIL.n325 B 1.23461f
C363 VTAIL.n326 B 0.008583f
C364 VTAIL.t1 B 0.033596f
C365 VTAIL.n327 B 0.114865f
C366 VTAIL.n328 B 0.011984f
C367 VTAIL.n329 B 0.015215f
C368 VTAIL.n330 B 0.020286f
C369 VTAIL.n331 B 0.009088f
C370 VTAIL.n332 B 0.008583f
C371 VTAIL.n333 B 0.015972f
C372 VTAIL.n334 B 0.015972f
C373 VTAIL.n335 B 0.008583f
C374 VTAIL.n336 B 0.009088f
C375 VTAIL.n337 B 0.020286f
C376 VTAIL.n338 B 0.020286f
C377 VTAIL.n339 B 0.009088f
C378 VTAIL.n340 B 0.008583f
C379 VTAIL.n341 B 0.015972f
C380 VTAIL.n342 B 0.015972f
C381 VTAIL.n343 B 0.008583f
C382 VTAIL.n344 B 0.009088f
C383 VTAIL.n345 B 0.020286f
C384 VTAIL.n346 B 0.020286f
C385 VTAIL.n347 B 0.009088f
C386 VTAIL.n348 B 0.008583f
C387 VTAIL.n349 B 0.015972f
C388 VTAIL.n350 B 0.015972f
C389 VTAIL.n351 B 0.008583f
C390 VTAIL.n352 B 0.009088f
C391 VTAIL.n353 B 0.020286f
C392 VTAIL.n354 B 0.020286f
C393 VTAIL.n355 B 0.009088f
C394 VTAIL.n356 B 0.008583f
C395 VTAIL.n357 B 0.015972f
C396 VTAIL.n358 B 0.015972f
C397 VTAIL.n359 B 0.008583f
C398 VTAIL.n360 B 0.009088f
C399 VTAIL.n361 B 0.020286f
C400 VTAIL.n362 B 0.020286f
C401 VTAIL.n363 B 0.009088f
C402 VTAIL.n364 B 0.008583f
C403 VTAIL.n365 B 0.015972f
C404 VTAIL.n366 B 0.015972f
C405 VTAIL.n367 B 0.008583f
C406 VTAIL.n368 B 0.009088f
C407 VTAIL.n369 B 0.020286f
C408 VTAIL.n370 B 0.020286f
C409 VTAIL.n371 B 0.009088f
C410 VTAIL.n372 B 0.008583f
C411 VTAIL.n373 B 0.015972f
C412 VTAIL.n374 B 0.015972f
C413 VTAIL.n375 B 0.008583f
C414 VTAIL.n376 B 0.009088f
C415 VTAIL.n377 B 0.020286f
C416 VTAIL.n378 B 0.020286f
C417 VTAIL.n379 B 0.009088f
C418 VTAIL.n380 B 0.008583f
C419 VTAIL.n381 B 0.015972f
C420 VTAIL.n382 B 0.015972f
C421 VTAIL.n383 B 0.008583f
C422 VTAIL.n384 B 0.009088f
C423 VTAIL.n385 B 0.020286f
C424 VTAIL.n386 B 0.046013f
C425 VTAIL.n387 B 0.009088f
C426 VTAIL.n388 B 0.008583f
C427 VTAIL.n389 B 0.040192f
C428 VTAIL.n390 B 0.026058f
C429 VTAIL.n391 B 1.40063f
C430 VTAIL.n392 B 0.023636f
C431 VTAIL.n393 B 0.015972f
C432 VTAIL.n394 B 0.008583f
C433 VTAIL.n395 B 0.020286f
C434 VTAIL.n396 B 0.009088f
C435 VTAIL.n397 B 0.015972f
C436 VTAIL.n398 B 0.008583f
C437 VTAIL.n399 B 0.020286f
C438 VTAIL.n400 B 0.008835f
C439 VTAIL.n401 B 0.015972f
C440 VTAIL.n402 B 0.008835f
C441 VTAIL.n403 B 0.008583f
C442 VTAIL.n404 B 0.020286f
C443 VTAIL.n405 B 0.020286f
C444 VTAIL.n406 B 0.009088f
C445 VTAIL.n407 B 0.015972f
C446 VTAIL.n408 B 0.008583f
C447 VTAIL.n409 B 0.020286f
C448 VTAIL.n410 B 0.009088f
C449 VTAIL.n411 B 0.015972f
C450 VTAIL.n412 B 0.008583f
C451 VTAIL.n413 B 0.020286f
C452 VTAIL.n414 B 0.009088f
C453 VTAIL.n415 B 0.015972f
C454 VTAIL.n416 B 0.008583f
C455 VTAIL.n417 B 0.020286f
C456 VTAIL.n418 B 0.009088f
C457 VTAIL.n419 B 0.015972f
C458 VTAIL.n420 B 0.008583f
C459 VTAIL.n421 B 0.020286f
C460 VTAIL.n422 B 0.009088f
C461 VTAIL.n423 B 1.23461f
C462 VTAIL.n424 B 0.008583f
C463 VTAIL.t0 B 0.033596f
C464 VTAIL.n425 B 0.114865f
C465 VTAIL.n426 B 0.011984f
C466 VTAIL.n427 B 0.015215f
C467 VTAIL.n428 B 0.020286f
C468 VTAIL.n429 B 0.009088f
C469 VTAIL.n430 B 0.008583f
C470 VTAIL.n431 B 0.015972f
C471 VTAIL.n432 B 0.015972f
C472 VTAIL.n433 B 0.008583f
C473 VTAIL.n434 B 0.009088f
C474 VTAIL.n435 B 0.020286f
C475 VTAIL.n436 B 0.020286f
C476 VTAIL.n437 B 0.009088f
C477 VTAIL.n438 B 0.008583f
C478 VTAIL.n439 B 0.015972f
C479 VTAIL.n440 B 0.015972f
C480 VTAIL.n441 B 0.008583f
C481 VTAIL.n442 B 0.009088f
C482 VTAIL.n443 B 0.020286f
C483 VTAIL.n444 B 0.020286f
C484 VTAIL.n445 B 0.009088f
C485 VTAIL.n446 B 0.008583f
C486 VTAIL.n447 B 0.015972f
C487 VTAIL.n448 B 0.015972f
C488 VTAIL.n449 B 0.008583f
C489 VTAIL.n450 B 0.009088f
C490 VTAIL.n451 B 0.020286f
C491 VTAIL.n452 B 0.020286f
C492 VTAIL.n453 B 0.009088f
C493 VTAIL.n454 B 0.008583f
C494 VTAIL.n455 B 0.015972f
C495 VTAIL.n456 B 0.015972f
C496 VTAIL.n457 B 0.008583f
C497 VTAIL.n458 B 0.009088f
C498 VTAIL.n459 B 0.020286f
C499 VTAIL.n460 B 0.020286f
C500 VTAIL.n461 B 0.009088f
C501 VTAIL.n462 B 0.008583f
C502 VTAIL.n463 B 0.015972f
C503 VTAIL.n464 B 0.015972f
C504 VTAIL.n465 B 0.008583f
C505 VTAIL.n466 B 0.009088f
C506 VTAIL.n467 B 0.020286f
C507 VTAIL.n468 B 0.020286f
C508 VTAIL.n469 B 0.009088f
C509 VTAIL.n470 B 0.008583f
C510 VTAIL.n471 B 0.015972f
C511 VTAIL.n472 B 0.015972f
C512 VTAIL.n473 B 0.008583f
C513 VTAIL.n474 B 0.009088f
C514 VTAIL.n475 B 0.020286f
C515 VTAIL.n476 B 0.020286f
C516 VTAIL.n477 B 0.009088f
C517 VTAIL.n478 B 0.008583f
C518 VTAIL.n479 B 0.015972f
C519 VTAIL.n480 B 0.015972f
C520 VTAIL.n481 B 0.008583f
C521 VTAIL.n482 B 0.009088f
C522 VTAIL.n483 B 0.020286f
C523 VTAIL.n484 B 0.046013f
C524 VTAIL.n485 B 0.009088f
C525 VTAIL.n486 B 0.008583f
C526 VTAIL.n487 B 0.040192f
C527 VTAIL.n488 B 0.026058f
C528 VTAIL.n489 B 0.231781f
C529 VTAIL.n490 B 0.023636f
C530 VTAIL.n491 B 0.015972f
C531 VTAIL.n492 B 0.008583f
C532 VTAIL.n493 B 0.020286f
C533 VTAIL.n494 B 0.009088f
C534 VTAIL.n495 B 0.015972f
C535 VTAIL.n496 B 0.008583f
C536 VTAIL.n497 B 0.020286f
C537 VTAIL.n498 B 0.008835f
C538 VTAIL.n499 B 0.015972f
C539 VTAIL.n500 B 0.008835f
C540 VTAIL.n501 B 0.008583f
C541 VTAIL.n502 B 0.020286f
C542 VTAIL.n503 B 0.020286f
C543 VTAIL.n504 B 0.009088f
C544 VTAIL.n505 B 0.015972f
C545 VTAIL.n506 B 0.008583f
C546 VTAIL.n507 B 0.020286f
C547 VTAIL.n508 B 0.009088f
C548 VTAIL.n509 B 0.015972f
C549 VTAIL.n510 B 0.008583f
C550 VTAIL.n511 B 0.020286f
C551 VTAIL.n512 B 0.009088f
C552 VTAIL.n513 B 0.015972f
C553 VTAIL.n514 B 0.008583f
C554 VTAIL.n515 B 0.020286f
C555 VTAIL.n516 B 0.009088f
C556 VTAIL.n517 B 0.015972f
C557 VTAIL.n518 B 0.008583f
C558 VTAIL.n519 B 0.020286f
C559 VTAIL.n520 B 0.009088f
C560 VTAIL.n521 B 1.23461f
C561 VTAIL.n522 B 0.008583f
C562 VTAIL.t5 B 0.033596f
C563 VTAIL.n523 B 0.114865f
C564 VTAIL.n524 B 0.011984f
C565 VTAIL.n525 B 0.015215f
C566 VTAIL.n526 B 0.020286f
C567 VTAIL.n527 B 0.009088f
C568 VTAIL.n528 B 0.008583f
C569 VTAIL.n529 B 0.015972f
C570 VTAIL.n530 B 0.015972f
C571 VTAIL.n531 B 0.008583f
C572 VTAIL.n532 B 0.009088f
C573 VTAIL.n533 B 0.020286f
C574 VTAIL.n534 B 0.020286f
C575 VTAIL.n535 B 0.009088f
C576 VTAIL.n536 B 0.008583f
C577 VTAIL.n537 B 0.015972f
C578 VTAIL.n538 B 0.015972f
C579 VTAIL.n539 B 0.008583f
C580 VTAIL.n540 B 0.009088f
C581 VTAIL.n541 B 0.020286f
C582 VTAIL.n542 B 0.020286f
C583 VTAIL.n543 B 0.009088f
C584 VTAIL.n544 B 0.008583f
C585 VTAIL.n545 B 0.015972f
C586 VTAIL.n546 B 0.015972f
C587 VTAIL.n547 B 0.008583f
C588 VTAIL.n548 B 0.009088f
C589 VTAIL.n549 B 0.020286f
C590 VTAIL.n550 B 0.020286f
C591 VTAIL.n551 B 0.009088f
C592 VTAIL.n552 B 0.008583f
C593 VTAIL.n553 B 0.015972f
C594 VTAIL.n554 B 0.015972f
C595 VTAIL.n555 B 0.008583f
C596 VTAIL.n556 B 0.009088f
C597 VTAIL.n557 B 0.020286f
C598 VTAIL.n558 B 0.020286f
C599 VTAIL.n559 B 0.009088f
C600 VTAIL.n560 B 0.008583f
C601 VTAIL.n561 B 0.015972f
C602 VTAIL.n562 B 0.015972f
C603 VTAIL.n563 B 0.008583f
C604 VTAIL.n564 B 0.009088f
C605 VTAIL.n565 B 0.020286f
C606 VTAIL.n566 B 0.020286f
C607 VTAIL.n567 B 0.009088f
C608 VTAIL.n568 B 0.008583f
C609 VTAIL.n569 B 0.015972f
C610 VTAIL.n570 B 0.015972f
C611 VTAIL.n571 B 0.008583f
C612 VTAIL.n572 B 0.009088f
C613 VTAIL.n573 B 0.020286f
C614 VTAIL.n574 B 0.020286f
C615 VTAIL.n575 B 0.009088f
C616 VTAIL.n576 B 0.008583f
C617 VTAIL.n577 B 0.015972f
C618 VTAIL.n578 B 0.015972f
C619 VTAIL.n579 B 0.008583f
C620 VTAIL.n580 B 0.009088f
C621 VTAIL.n581 B 0.020286f
C622 VTAIL.n582 B 0.046013f
C623 VTAIL.n583 B 0.009088f
C624 VTAIL.n584 B 0.008583f
C625 VTAIL.n585 B 0.040192f
C626 VTAIL.n586 B 0.026058f
C627 VTAIL.n587 B 0.231781f
C628 VTAIL.n588 B 0.023636f
C629 VTAIL.n589 B 0.015972f
C630 VTAIL.n590 B 0.008583f
C631 VTAIL.n591 B 0.020286f
C632 VTAIL.n592 B 0.009088f
C633 VTAIL.n593 B 0.015972f
C634 VTAIL.n594 B 0.008583f
C635 VTAIL.n595 B 0.020286f
C636 VTAIL.n596 B 0.008835f
C637 VTAIL.n597 B 0.015972f
C638 VTAIL.n598 B 0.008835f
C639 VTAIL.n599 B 0.008583f
C640 VTAIL.n600 B 0.020286f
C641 VTAIL.n601 B 0.020286f
C642 VTAIL.n602 B 0.009088f
C643 VTAIL.n603 B 0.015972f
C644 VTAIL.n604 B 0.008583f
C645 VTAIL.n605 B 0.020286f
C646 VTAIL.n606 B 0.009088f
C647 VTAIL.n607 B 0.015972f
C648 VTAIL.n608 B 0.008583f
C649 VTAIL.n609 B 0.020286f
C650 VTAIL.n610 B 0.009088f
C651 VTAIL.n611 B 0.015972f
C652 VTAIL.n612 B 0.008583f
C653 VTAIL.n613 B 0.020286f
C654 VTAIL.n614 B 0.009088f
C655 VTAIL.n615 B 0.015972f
C656 VTAIL.n616 B 0.008583f
C657 VTAIL.n617 B 0.020286f
C658 VTAIL.n618 B 0.009088f
C659 VTAIL.n619 B 1.23461f
C660 VTAIL.n620 B 0.008583f
C661 VTAIL.t7 B 0.033596f
C662 VTAIL.n621 B 0.114865f
C663 VTAIL.n622 B 0.011984f
C664 VTAIL.n623 B 0.015215f
C665 VTAIL.n624 B 0.020286f
C666 VTAIL.n625 B 0.009088f
C667 VTAIL.n626 B 0.008583f
C668 VTAIL.n627 B 0.015972f
C669 VTAIL.n628 B 0.015972f
C670 VTAIL.n629 B 0.008583f
C671 VTAIL.n630 B 0.009088f
C672 VTAIL.n631 B 0.020286f
C673 VTAIL.n632 B 0.020286f
C674 VTAIL.n633 B 0.009088f
C675 VTAIL.n634 B 0.008583f
C676 VTAIL.n635 B 0.015972f
C677 VTAIL.n636 B 0.015972f
C678 VTAIL.n637 B 0.008583f
C679 VTAIL.n638 B 0.009088f
C680 VTAIL.n639 B 0.020286f
C681 VTAIL.n640 B 0.020286f
C682 VTAIL.n641 B 0.009088f
C683 VTAIL.n642 B 0.008583f
C684 VTAIL.n643 B 0.015972f
C685 VTAIL.n644 B 0.015972f
C686 VTAIL.n645 B 0.008583f
C687 VTAIL.n646 B 0.009088f
C688 VTAIL.n647 B 0.020286f
C689 VTAIL.n648 B 0.020286f
C690 VTAIL.n649 B 0.009088f
C691 VTAIL.n650 B 0.008583f
C692 VTAIL.n651 B 0.015972f
C693 VTAIL.n652 B 0.015972f
C694 VTAIL.n653 B 0.008583f
C695 VTAIL.n654 B 0.009088f
C696 VTAIL.n655 B 0.020286f
C697 VTAIL.n656 B 0.020286f
C698 VTAIL.n657 B 0.009088f
C699 VTAIL.n658 B 0.008583f
C700 VTAIL.n659 B 0.015972f
C701 VTAIL.n660 B 0.015972f
C702 VTAIL.n661 B 0.008583f
C703 VTAIL.n662 B 0.009088f
C704 VTAIL.n663 B 0.020286f
C705 VTAIL.n664 B 0.020286f
C706 VTAIL.n665 B 0.009088f
C707 VTAIL.n666 B 0.008583f
C708 VTAIL.n667 B 0.015972f
C709 VTAIL.n668 B 0.015972f
C710 VTAIL.n669 B 0.008583f
C711 VTAIL.n670 B 0.009088f
C712 VTAIL.n671 B 0.020286f
C713 VTAIL.n672 B 0.020286f
C714 VTAIL.n673 B 0.009088f
C715 VTAIL.n674 B 0.008583f
C716 VTAIL.n675 B 0.015972f
C717 VTAIL.n676 B 0.015972f
C718 VTAIL.n677 B 0.008583f
C719 VTAIL.n678 B 0.009088f
C720 VTAIL.n679 B 0.020286f
C721 VTAIL.n680 B 0.046013f
C722 VTAIL.n681 B 0.009088f
C723 VTAIL.n682 B 0.008583f
C724 VTAIL.n683 B 0.040192f
C725 VTAIL.n684 B 0.026058f
C726 VTAIL.n685 B 1.40063f
C727 VTAIL.n686 B 0.023636f
C728 VTAIL.n687 B 0.015972f
C729 VTAIL.n688 B 0.008583f
C730 VTAIL.n689 B 0.020286f
C731 VTAIL.n690 B 0.009088f
C732 VTAIL.n691 B 0.015972f
C733 VTAIL.n692 B 0.008583f
C734 VTAIL.n693 B 0.020286f
C735 VTAIL.n694 B 0.008835f
C736 VTAIL.n695 B 0.015972f
C737 VTAIL.n696 B 0.009088f
C738 VTAIL.n697 B 0.020286f
C739 VTAIL.n698 B 0.009088f
C740 VTAIL.n699 B 0.015972f
C741 VTAIL.n700 B 0.008583f
C742 VTAIL.n701 B 0.020286f
C743 VTAIL.n702 B 0.009088f
C744 VTAIL.n703 B 0.015972f
C745 VTAIL.n704 B 0.008583f
C746 VTAIL.n705 B 0.020286f
C747 VTAIL.n706 B 0.009088f
C748 VTAIL.n707 B 0.015972f
C749 VTAIL.n708 B 0.008583f
C750 VTAIL.n709 B 0.020286f
C751 VTAIL.n710 B 0.009088f
C752 VTAIL.n711 B 0.015972f
C753 VTAIL.n712 B 0.008583f
C754 VTAIL.n713 B 0.020286f
C755 VTAIL.n714 B 0.009088f
C756 VTAIL.n715 B 1.23461f
C757 VTAIL.n716 B 0.008583f
C758 VTAIL.t3 B 0.033596f
C759 VTAIL.n717 B 0.114865f
C760 VTAIL.n718 B 0.011984f
C761 VTAIL.n719 B 0.015215f
C762 VTAIL.n720 B 0.020286f
C763 VTAIL.n721 B 0.009088f
C764 VTAIL.n722 B 0.008583f
C765 VTAIL.n723 B 0.015972f
C766 VTAIL.n724 B 0.015972f
C767 VTAIL.n725 B 0.008583f
C768 VTAIL.n726 B 0.009088f
C769 VTAIL.n727 B 0.020286f
C770 VTAIL.n728 B 0.020286f
C771 VTAIL.n729 B 0.009088f
C772 VTAIL.n730 B 0.008583f
C773 VTAIL.n731 B 0.015972f
C774 VTAIL.n732 B 0.015972f
C775 VTAIL.n733 B 0.008583f
C776 VTAIL.n734 B 0.009088f
C777 VTAIL.n735 B 0.020286f
C778 VTAIL.n736 B 0.020286f
C779 VTAIL.n737 B 0.009088f
C780 VTAIL.n738 B 0.008583f
C781 VTAIL.n739 B 0.015972f
C782 VTAIL.n740 B 0.015972f
C783 VTAIL.n741 B 0.008583f
C784 VTAIL.n742 B 0.009088f
C785 VTAIL.n743 B 0.020286f
C786 VTAIL.n744 B 0.020286f
C787 VTAIL.n745 B 0.009088f
C788 VTAIL.n746 B 0.008583f
C789 VTAIL.n747 B 0.015972f
C790 VTAIL.n748 B 0.015972f
C791 VTAIL.n749 B 0.008583f
C792 VTAIL.n750 B 0.009088f
C793 VTAIL.n751 B 0.020286f
C794 VTAIL.n752 B 0.020286f
C795 VTAIL.n753 B 0.009088f
C796 VTAIL.n754 B 0.008583f
C797 VTAIL.n755 B 0.015972f
C798 VTAIL.n756 B 0.015972f
C799 VTAIL.n757 B 0.008583f
C800 VTAIL.n758 B 0.008583f
C801 VTAIL.n759 B 0.009088f
C802 VTAIL.n760 B 0.020286f
C803 VTAIL.n761 B 0.020286f
C804 VTAIL.n762 B 0.020286f
C805 VTAIL.n763 B 0.008835f
C806 VTAIL.n764 B 0.008583f
C807 VTAIL.n765 B 0.015972f
C808 VTAIL.n766 B 0.015972f
C809 VTAIL.n767 B 0.008583f
C810 VTAIL.n768 B 0.009088f
C811 VTAIL.n769 B 0.020286f
C812 VTAIL.n770 B 0.020286f
C813 VTAIL.n771 B 0.009088f
C814 VTAIL.n772 B 0.008583f
C815 VTAIL.n773 B 0.015972f
C816 VTAIL.n774 B 0.015972f
C817 VTAIL.n775 B 0.008583f
C818 VTAIL.n776 B 0.009088f
C819 VTAIL.n777 B 0.020286f
C820 VTAIL.n778 B 0.046013f
C821 VTAIL.n779 B 0.009088f
C822 VTAIL.n780 B 0.008583f
C823 VTAIL.n781 B 0.040192f
C824 VTAIL.n782 B 0.026058f
C825 VTAIL.n783 B 1.30158f
C826 VP.n0 B 0.034561f
C827 VP.t0 B 3.5708f
C828 VP.n1 B 0.034244f
C829 VP.n2 B 0.018374f
C830 VP.n3 B 0.034244f
C831 VP.t3 B 3.8907f
C832 VP.t1 B 3.90432f
C833 VP.n4 B 3.71495f
C834 VP.n5 B 1.27934f
C835 VP.t2 B 3.5708f
C836 VP.n6 B 1.31117f
C837 VP.n7 B 0.031369f
C838 VP.n8 B 0.034561f
C839 VP.n9 B 0.018374f
C840 VP.n10 B 0.018374f
C841 VP.n11 B 0.034244f
C842 VP.n12 B 0.026823f
C843 VP.n13 B 0.026823f
C844 VP.n14 B 0.018374f
C845 VP.n15 B 0.018374f
C846 VP.n16 B 0.018374f
C847 VP.n17 B 0.034244f
C848 VP.n18 B 0.031369f
C849 VP.n19 B 1.31117f
C850 VP.n20 B 0.058726f
.ends

