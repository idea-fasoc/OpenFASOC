* NGSPICE file created from diff_pair_sample_1667.ext - technology: sky130A

.subckt diff_pair_sample_1667 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0 ps=0 w=3.23 l=1.61
X1 VDD2.t9 VN.t0 VTAIL.t16 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=1.2597 ps=7.24 w=3.23 l=1.61
X2 VDD1.t9 VP.t0 VTAIL.t4 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=1.2597 ps=7.24 w=3.23 l=1.61
X3 VDD2.t8 VN.t1 VTAIL.t10 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0.53295 ps=3.56 w=3.23 l=1.61
X4 VTAIL.t13 VN.t2 VDD2.t7 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X5 VDD2.t6 VN.t3 VTAIL.t12 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X6 VDD1.t8 VP.t1 VTAIL.t19 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X7 VDD1.t7 VP.t2 VTAIL.t5 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0.53295 ps=3.56 w=3.23 l=1.61
X8 B.t8 B.t6 B.t7 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0 ps=0 w=3.23 l=1.61
X9 VTAIL.t2 VP.t3 VDD1.t6 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X10 B.t5 B.t3 B.t4 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0 ps=0 w=3.23 l=1.61
X11 VDD2.t5 VN.t4 VTAIL.t14 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=1.2597 ps=7.24 w=3.23 l=1.61
X12 B.t2 B.t0 B.t1 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0 ps=0 w=3.23 l=1.61
X13 VTAIL.t9 VN.t5 VDD2.t4 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X14 VTAIL.t0 VP.t4 VDD1.t5 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X15 VTAIL.t1 VP.t5 VDD1.t4 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X16 VDD1.t3 VP.t6 VTAIL.t6 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X17 VTAIL.t15 VN.t6 VDD2.t3 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X18 VTAIL.t17 VN.t7 VDD2.t2 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X19 VDD1.t2 VP.t7 VTAIL.t3 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0.53295 ps=3.56 w=3.23 l=1.61
X20 VDD1.t1 VP.t8 VTAIL.t7 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=1.2597 ps=7.24 w=3.23 l=1.61
X21 VDD2.t1 VN.t8 VTAIL.t11 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X22 VTAIL.t8 VP.t9 VDD1.t0 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=0.53295 pd=3.56 as=0.53295 ps=3.56 w=3.23 l=1.61
X23 VDD2.t0 VN.t9 VTAIL.t18 w_n3298_n1614# sky130_fd_pr__pfet_01v8 ad=1.2597 pd=7.24 as=0.53295 ps=3.56 w=3.23 l=1.61
R0 B.n260 B.n259 585
R1 B.n258 B.n91 585
R2 B.n257 B.n256 585
R3 B.n255 B.n92 585
R4 B.n254 B.n253 585
R5 B.n252 B.n93 585
R6 B.n251 B.n250 585
R7 B.n249 B.n94 585
R8 B.n248 B.n247 585
R9 B.n246 B.n95 585
R10 B.n245 B.n244 585
R11 B.n243 B.n96 585
R12 B.n242 B.n241 585
R13 B.n240 B.n97 585
R14 B.n239 B.n238 585
R15 B.n237 B.n98 585
R16 B.n236 B.n235 585
R17 B.n231 B.n99 585
R18 B.n230 B.n229 585
R19 B.n228 B.n100 585
R20 B.n227 B.n226 585
R21 B.n225 B.n101 585
R22 B.n224 B.n223 585
R23 B.n222 B.n102 585
R24 B.n221 B.n220 585
R25 B.n218 B.n103 585
R26 B.n217 B.n216 585
R27 B.n215 B.n106 585
R28 B.n214 B.n213 585
R29 B.n212 B.n107 585
R30 B.n211 B.n210 585
R31 B.n209 B.n108 585
R32 B.n208 B.n207 585
R33 B.n206 B.n109 585
R34 B.n205 B.n204 585
R35 B.n203 B.n110 585
R36 B.n202 B.n201 585
R37 B.n200 B.n111 585
R38 B.n199 B.n198 585
R39 B.n197 B.n112 585
R40 B.n196 B.n195 585
R41 B.n261 B.n90 585
R42 B.n263 B.n262 585
R43 B.n264 B.n89 585
R44 B.n266 B.n265 585
R45 B.n267 B.n88 585
R46 B.n269 B.n268 585
R47 B.n270 B.n87 585
R48 B.n272 B.n271 585
R49 B.n273 B.n86 585
R50 B.n275 B.n274 585
R51 B.n276 B.n85 585
R52 B.n278 B.n277 585
R53 B.n279 B.n84 585
R54 B.n281 B.n280 585
R55 B.n282 B.n83 585
R56 B.n284 B.n283 585
R57 B.n285 B.n82 585
R58 B.n287 B.n286 585
R59 B.n288 B.n81 585
R60 B.n290 B.n289 585
R61 B.n291 B.n80 585
R62 B.n293 B.n292 585
R63 B.n294 B.n79 585
R64 B.n296 B.n295 585
R65 B.n297 B.n78 585
R66 B.n299 B.n298 585
R67 B.n300 B.n77 585
R68 B.n302 B.n301 585
R69 B.n303 B.n76 585
R70 B.n305 B.n304 585
R71 B.n306 B.n75 585
R72 B.n308 B.n307 585
R73 B.n309 B.n74 585
R74 B.n311 B.n310 585
R75 B.n312 B.n73 585
R76 B.n314 B.n313 585
R77 B.n315 B.n72 585
R78 B.n317 B.n316 585
R79 B.n318 B.n71 585
R80 B.n320 B.n319 585
R81 B.n321 B.n70 585
R82 B.n323 B.n322 585
R83 B.n324 B.n69 585
R84 B.n326 B.n325 585
R85 B.n327 B.n68 585
R86 B.n329 B.n328 585
R87 B.n330 B.n67 585
R88 B.n332 B.n331 585
R89 B.n333 B.n66 585
R90 B.n335 B.n334 585
R91 B.n336 B.n65 585
R92 B.n338 B.n337 585
R93 B.n339 B.n64 585
R94 B.n341 B.n340 585
R95 B.n342 B.n63 585
R96 B.n344 B.n343 585
R97 B.n345 B.n62 585
R98 B.n347 B.n346 585
R99 B.n348 B.n61 585
R100 B.n350 B.n349 585
R101 B.n351 B.n60 585
R102 B.n353 B.n352 585
R103 B.n354 B.n59 585
R104 B.n356 B.n355 585
R105 B.n357 B.n58 585
R106 B.n359 B.n358 585
R107 B.n360 B.n57 585
R108 B.n362 B.n361 585
R109 B.n363 B.n56 585
R110 B.n365 B.n364 585
R111 B.n366 B.n55 585
R112 B.n368 B.n367 585
R113 B.n369 B.n54 585
R114 B.n371 B.n370 585
R115 B.n372 B.n53 585
R116 B.n374 B.n373 585
R117 B.n375 B.n52 585
R118 B.n377 B.n376 585
R119 B.n378 B.n51 585
R120 B.n380 B.n379 585
R121 B.n381 B.n50 585
R122 B.n383 B.n382 585
R123 B.n384 B.n49 585
R124 B.n386 B.n385 585
R125 B.n387 B.n48 585
R126 B.n389 B.n388 585
R127 B.n452 B.n23 585
R128 B.n451 B.n450 585
R129 B.n449 B.n24 585
R130 B.n448 B.n447 585
R131 B.n446 B.n25 585
R132 B.n445 B.n444 585
R133 B.n443 B.n26 585
R134 B.n442 B.n441 585
R135 B.n440 B.n27 585
R136 B.n439 B.n438 585
R137 B.n437 B.n28 585
R138 B.n436 B.n435 585
R139 B.n434 B.n29 585
R140 B.n433 B.n432 585
R141 B.n431 B.n30 585
R142 B.n430 B.n429 585
R143 B.n427 B.n31 585
R144 B.n426 B.n425 585
R145 B.n424 B.n34 585
R146 B.n423 B.n422 585
R147 B.n421 B.n35 585
R148 B.n420 B.n419 585
R149 B.n418 B.n36 585
R150 B.n417 B.n416 585
R151 B.n415 B.n37 585
R152 B.n413 B.n412 585
R153 B.n411 B.n40 585
R154 B.n410 B.n409 585
R155 B.n408 B.n41 585
R156 B.n407 B.n406 585
R157 B.n405 B.n42 585
R158 B.n404 B.n403 585
R159 B.n402 B.n43 585
R160 B.n401 B.n400 585
R161 B.n399 B.n44 585
R162 B.n398 B.n397 585
R163 B.n396 B.n45 585
R164 B.n395 B.n394 585
R165 B.n393 B.n46 585
R166 B.n392 B.n391 585
R167 B.n390 B.n47 585
R168 B.n454 B.n453 585
R169 B.n455 B.n22 585
R170 B.n457 B.n456 585
R171 B.n458 B.n21 585
R172 B.n460 B.n459 585
R173 B.n461 B.n20 585
R174 B.n463 B.n462 585
R175 B.n464 B.n19 585
R176 B.n466 B.n465 585
R177 B.n467 B.n18 585
R178 B.n469 B.n468 585
R179 B.n470 B.n17 585
R180 B.n472 B.n471 585
R181 B.n473 B.n16 585
R182 B.n475 B.n474 585
R183 B.n476 B.n15 585
R184 B.n478 B.n477 585
R185 B.n479 B.n14 585
R186 B.n481 B.n480 585
R187 B.n482 B.n13 585
R188 B.n484 B.n483 585
R189 B.n485 B.n12 585
R190 B.n487 B.n486 585
R191 B.n488 B.n11 585
R192 B.n490 B.n489 585
R193 B.n491 B.n10 585
R194 B.n493 B.n492 585
R195 B.n494 B.n9 585
R196 B.n496 B.n495 585
R197 B.n497 B.n8 585
R198 B.n499 B.n498 585
R199 B.n500 B.n7 585
R200 B.n502 B.n501 585
R201 B.n503 B.n6 585
R202 B.n505 B.n504 585
R203 B.n506 B.n5 585
R204 B.n508 B.n507 585
R205 B.n509 B.n4 585
R206 B.n511 B.n510 585
R207 B.n512 B.n3 585
R208 B.n514 B.n513 585
R209 B.n515 B.n0 585
R210 B.n2 B.n1 585
R211 B.n134 B.n133 585
R212 B.n136 B.n135 585
R213 B.n137 B.n132 585
R214 B.n139 B.n138 585
R215 B.n140 B.n131 585
R216 B.n142 B.n141 585
R217 B.n143 B.n130 585
R218 B.n145 B.n144 585
R219 B.n146 B.n129 585
R220 B.n148 B.n147 585
R221 B.n149 B.n128 585
R222 B.n151 B.n150 585
R223 B.n152 B.n127 585
R224 B.n154 B.n153 585
R225 B.n155 B.n126 585
R226 B.n157 B.n156 585
R227 B.n158 B.n125 585
R228 B.n160 B.n159 585
R229 B.n161 B.n124 585
R230 B.n163 B.n162 585
R231 B.n164 B.n123 585
R232 B.n166 B.n165 585
R233 B.n167 B.n122 585
R234 B.n169 B.n168 585
R235 B.n170 B.n121 585
R236 B.n172 B.n171 585
R237 B.n173 B.n120 585
R238 B.n175 B.n174 585
R239 B.n176 B.n119 585
R240 B.n178 B.n177 585
R241 B.n179 B.n118 585
R242 B.n181 B.n180 585
R243 B.n182 B.n117 585
R244 B.n184 B.n183 585
R245 B.n185 B.n116 585
R246 B.n187 B.n186 585
R247 B.n188 B.n115 585
R248 B.n190 B.n189 585
R249 B.n191 B.n114 585
R250 B.n193 B.n192 585
R251 B.n194 B.n113 585
R252 B.n196 B.n113 492.5
R253 B.n261 B.n260 492.5
R254 B.n388 B.n47 492.5
R255 B.n454 B.n23 492.5
R256 B.n232 B.t1 263.767
R257 B.n38 B.t8 263.767
R258 B.n104 B.t10 263.767
R259 B.n32 B.t5 263.767
R260 B.n517 B.n516 256.663
R261 B.n104 B.t9 254.178
R262 B.n232 B.t0 254.178
R263 B.n38 B.t6 254.178
R264 B.n32 B.t3 254.178
R265 B.n516 B.n515 235.042
R266 B.n516 B.n2 235.042
R267 B.n233 B.t2 226.143
R268 B.n39 B.t7 226.143
R269 B.n105 B.t11 226.143
R270 B.n33 B.t4 226.143
R271 B.n197 B.n196 163.367
R272 B.n198 B.n197 163.367
R273 B.n198 B.n111 163.367
R274 B.n202 B.n111 163.367
R275 B.n203 B.n202 163.367
R276 B.n204 B.n203 163.367
R277 B.n204 B.n109 163.367
R278 B.n208 B.n109 163.367
R279 B.n209 B.n208 163.367
R280 B.n210 B.n209 163.367
R281 B.n210 B.n107 163.367
R282 B.n214 B.n107 163.367
R283 B.n215 B.n214 163.367
R284 B.n216 B.n215 163.367
R285 B.n216 B.n103 163.367
R286 B.n221 B.n103 163.367
R287 B.n222 B.n221 163.367
R288 B.n223 B.n222 163.367
R289 B.n223 B.n101 163.367
R290 B.n227 B.n101 163.367
R291 B.n228 B.n227 163.367
R292 B.n229 B.n228 163.367
R293 B.n229 B.n99 163.367
R294 B.n236 B.n99 163.367
R295 B.n237 B.n236 163.367
R296 B.n238 B.n237 163.367
R297 B.n238 B.n97 163.367
R298 B.n242 B.n97 163.367
R299 B.n243 B.n242 163.367
R300 B.n244 B.n243 163.367
R301 B.n244 B.n95 163.367
R302 B.n248 B.n95 163.367
R303 B.n249 B.n248 163.367
R304 B.n250 B.n249 163.367
R305 B.n250 B.n93 163.367
R306 B.n254 B.n93 163.367
R307 B.n255 B.n254 163.367
R308 B.n256 B.n255 163.367
R309 B.n256 B.n91 163.367
R310 B.n260 B.n91 163.367
R311 B.n388 B.n387 163.367
R312 B.n387 B.n386 163.367
R313 B.n386 B.n49 163.367
R314 B.n382 B.n49 163.367
R315 B.n382 B.n381 163.367
R316 B.n381 B.n380 163.367
R317 B.n380 B.n51 163.367
R318 B.n376 B.n51 163.367
R319 B.n376 B.n375 163.367
R320 B.n375 B.n374 163.367
R321 B.n374 B.n53 163.367
R322 B.n370 B.n53 163.367
R323 B.n370 B.n369 163.367
R324 B.n369 B.n368 163.367
R325 B.n368 B.n55 163.367
R326 B.n364 B.n55 163.367
R327 B.n364 B.n363 163.367
R328 B.n363 B.n362 163.367
R329 B.n362 B.n57 163.367
R330 B.n358 B.n57 163.367
R331 B.n358 B.n357 163.367
R332 B.n357 B.n356 163.367
R333 B.n356 B.n59 163.367
R334 B.n352 B.n59 163.367
R335 B.n352 B.n351 163.367
R336 B.n351 B.n350 163.367
R337 B.n350 B.n61 163.367
R338 B.n346 B.n61 163.367
R339 B.n346 B.n345 163.367
R340 B.n345 B.n344 163.367
R341 B.n344 B.n63 163.367
R342 B.n340 B.n63 163.367
R343 B.n340 B.n339 163.367
R344 B.n339 B.n338 163.367
R345 B.n338 B.n65 163.367
R346 B.n334 B.n65 163.367
R347 B.n334 B.n333 163.367
R348 B.n333 B.n332 163.367
R349 B.n332 B.n67 163.367
R350 B.n328 B.n67 163.367
R351 B.n328 B.n327 163.367
R352 B.n327 B.n326 163.367
R353 B.n326 B.n69 163.367
R354 B.n322 B.n69 163.367
R355 B.n322 B.n321 163.367
R356 B.n321 B.n320 163.367
R357 B.n320 B.n71 163.367
R358 B.n316 B.n71 163.367
R359 B.n316 B.n315 163.367
R360 B.n315 B.n314 163.367
R361 B.n314 B.n73 163.367
R362 B.n310 B.n73 163.367
R363 B.n310 B.n309 163.367
R364 B.n309 B.n308 163.367
R365 B.n308 B.n75 163.367
R366 B.n304 B.n75 163.367
R367 B.n304 B.n303 163.367
R368 B.n303 B.n302 163.367
R369 B.n302 B.n77 163.367
R370 B.n298 B.n77 163.367
R371 B.n298 B.n297 163.367
R372 B.n297 B.n296 163.367
R373 B.n296 B.n79 163.367
R374 B.n292 B.n79 163.367
R375 B.n292 B.n291 163.367
R376 B.n291 B.n290 163.367
R377 B.n290 B.n81 163.367
R378 B.n286 B.n81 163.367
R379 B.n286 B.n285 163.367
R380 B.n285 B.n284 163.367
R381 B.n284 B.n83 163.367
R382 B.n280 B.n83 163.367
R383 B.n280 B.n279 163.367
R384 B.n279 B.n278 163.367
R385 B.n278 B.n85 163.367
R386 B.n274 B.n85 163.367
R387 B.n274 B.n273 163.367
R388 B.n273 B.n272 163.367
R389 B.n272 B.n87 163.367
R390 B.n268 B.n87 163.367
R391 B.n268 B.n267 163.367
R392 B.n267 B.n266 163.367
R393 B.n266 B.n89 163.367
R394 B.n262 B.n89 163.367
R395 B.n262 B.n261 163.367
R396 B.n450 B.n23 163.367
R397 B.n450 B.n449 163.367
R398 B.n449 B.n448 163.367
R399 B.n448 B.n25 163.367
R400 B.n444 B.n25 163.367
R401 B.n444 B.n443 163.367
R402 B.n443 B.n442 163.367
R403 B.n442 B.n27 163.367
R404 B.n438 B.n27 163.367
R405 B.n438 B.n437 163.367
R406 B.n437 B.n436 163.367
R407 B.n436 B.n29 163.367
R408 B.n432 B.n29 163.367
R409 B.n432 B.n431 163.367
R410 B.n431 B.n430 163.367
R411 B.n430 B.n31 163.367
R412 B.n425 B.n31 163.367
R413 B.n425 B.n424 163.367
R414 B.n424 B.n423 163.367
R415 B.n423 B.n35 163.367
R416 B.n419 B.n35 163.367
R417 B.n419 B.n418 163.367
R418 B.n418 B.n417 163.367
R419 B.n417 B.n37 163.367
R420 B.n412 B.n37 163.367
R421 B.n412 B.n411 163.367
R422 B.n411 B.n410 163.367
R423 B.n410 B.n41 163.367
R424 B.n406 B.n41 163.367
R425 B.n406 B.n405 163.367
R426 B.n405 B.n404 163.367
R427 B.n404 B.n43 163.367
R428 B.n400 B.n43 163.367
R429 B.n400 B.n399 163.367
R430 B.n399 B.n398 163.367
R431 B.n398 B.n45 163.367
R432 B.n394 B.n45 163.367
R433 B.n394 B.n393 163.367
R434 B.n393 B.n392 163.367
R435 B.n392 B.n47 163.367
R436 B.n455 B.n454 163.367
R437 B.n456 B.n455 163.367
R438 B.n456 B.n21 163.367
R439 B.n460 B.n21 163.367
R440 B.n461 B.n460 163.367
R441 B.n462 B.n461 163.367
R442 B.n462 B.n19 163.367
R443 B.n466 B.n19 163.367
R444 B.n467 B.n466 163.367
R445 B.n468 B.n467 163.367
R446 B.n468 B.n17 163.367
R447 B.n472 B.n17 163.367
R448 B.n473 B.n472 163.367
R449 B.n474 B.n473 163.367
R450 B.n474 B.n15 163.367
R451 B.n478 B.n15 163.367
R452 B.n479 B.n478 163.367
R453 B.n480 B.n479 163.367
R454 B.n480 B.n13 163.367
R455 B.n484 B.n13 163.367
R456 B.n485 B.n484 163.367
R457 B.n486 B.n485 163.367
R458 B.n486 B.n11 163.367
R459 B.n490 B.n11 163.367
R460 B.n491 B.n490 163.367
R461 B.n492 B.n491 163.367
R462 B.n492 B.n9 163.367
R463 B.n496 B.n9 163.367
R464 B.n497 B.n496 163.367
R465 B.n498 B.n497 163.367
R466 B.n498 B.n7 163.367
R467 B.n502 B.n7 163.367
R468 B.n503 B.n502 163.367
R469 B.n504 B.n503 163.367
R470 B.n504 B.n5 163.367
R471 B.n508 B.n5 163.367
R472 B.n509 B.n508 163.367
R473 B.n510 B.n509 163.367
R474 B.n510 B.n3 163.367
R475 B.n514 B.n3 163.367
R476 B.n515 B.n514 163.367
R477 B.n133 B.n2 163.367
R478 B.n136 B.n133 163.367
R479 B.n137 B.n136 163.367
R480 B.n138 B.n137 163.367
R481 B.n138 B.n131 163.367
R482 B.n142 B.n131 163.367
R483 B.n143 B.n142 163.367
R484 B.n144 B.n143 163.367
R485 B.n144 B.n129 163.367
R486 B.n148 B.n129 163.367
R487 B.n149 B.n148 163.367
R488 B.n150 B.n149 163.367
R489 B.n150 B.n127 163.367
R490 B.n154 B.n127 163.367
R491 B.n155 B.n154 163.367
R492 B.n156 B.n155 163.367
R493 B.n156 B.n125 163.367
R494 B.n160 B.n125 163.367
R495 B.n161 B.n160 163.367
R496 B.n162 B.n161 163.367
R497 B.n162 B.n123 163.367
R498 B.n166 B.n123 163.367
R499 B.n167 B.n166 163.367
R500 B.n168 B.n167 163.367
R501 B.n168 B.n121 163.367
R502 B.n172 B.n121 163.367
R503 B.n173 B.n172 163.367
R504 B.n174 B.n173 163.367
R505 B.n174 B.n119 163.367
R506 B.n178 B.n119 163.367
R507 B.n179 B.n178 163.367
R508 B.n180 B.n179 163.367
R509 B.n180 B.n117 163.367
R510 B.n184 B.n117 163.367
R511 B.n185 B.n184 163.367
R512 B.n186 B.n185 163.367
R513 B.n186 B.n115 163.367
R514 B.n190 B.n115 163.367
R515 B.n191 B.n190 163.367
R516 B.n192 B.n191 163.367
R517 B.n192 B.n113 163.367
R518 B.n219 B.n105 59.5399
R519 B.n234 B.n233 59.5399
R520 B.n414 B.n39 59.5399
R521 B.n428 B.n33 59.5399
R522 B.n105 B.n104 37.6247
R523 B.n233 B.n232 37.6247
R524 B.n39 B.n38 37.6247
R525 B.n33 B.n32 37.6247
R526 B.n453 B.n452 32.0005
R527 B.n390 B.n389 32.0005
R528 B.n259 B.n90 32.0005
R529 B.n195 B.n194 32.0005
R530 B B.n517 18.0485
R531 B.n453 B.n22 10.6151
R532 B.n457 B.n22 10.6151
R533 B.n458 B.n457 10.6151
R534 B.n459 B.n458 10.6151
R535 B.n459 B.n20 10.6151
R536 B.n463 B.n20 10.6151
R537 B.n464 B.n463 10.6151
R538 B.n465 B.n464 10.6151
R539 B.n465 B.n18 10.6151
R540 B.n469 B.n18 10.6151
R541 B.n470 B.n469 10.6151
R542 B.n471 B.n470 10.6151
R543 B.n471 B.n16 10.6151
R544 B.n475 B.n16 10.6151
R545 B.n476 B.n475 10.6151
R546 B.n477 B.n476 10.6151
R547 B.n477 B.n14 10.6151
R548 B.n481 B.n14 10.6151
R549 B.n482 B.n481 10.6151
R550 B.n483 B.n482 10.6151
R551 B.n483 B.n12 10.6151
R552 B.n487 B.n12 10.6151
R553 B.n488 B.n487 10.6151
R554 B.n489 B.n488 10.6151
R555 B.n489 B.n10 10.6151
R556 B.n493 B.n10 10.6151
R557 B.n494 B.n493 10.6151
R558 B.n495 B.n494 10.6151
R559 B.n495 B.n8 10.6151
R560 B.n499 B.n8 10.6151
R561 B.n500 B.n499 10.6151
R562 B.n501 B.n500 10.6151
R563 B.n501 B.n6 10.6151
R564 B.n505 B.n6 10.6151
R565 B.n506 B.n505 10.6151
R566 B.n507 B.n506 10.6151
R567 B.n507 B.n4 10.6151
R568 B.n511 B.n4 10.6151
R569 B.n512 B.n511 10.6151
R570 B.n513 B.n512 10.6151
R571 B.n513 B.n0 10.6151
R572 B.n452 B.n451 10.6151
R573 B.n451 B.n24 10.6151
R574 B.n447 B.n24 10.6151
R575 B.n447 B.n446 10.6151
R576 B.n446 B.n445 10.6151
R577 B.n445 B.n26 10.6151
R578 B.n441 B.n26 10.6151
R579 B.n441 B.n440 10.6151
R580 B.n440 B.n439 10.6151
R581 B.n439 B.n28 10.6151
R582 B.n435 B.n28 10.6151
R583 B.n435 B.n434 10.6151
R584 B.n434 B.n433 10.6151
R585 B.n433 B.n30 10.6151
R586 B.n429 B.n30 10.6151
R587 B.n427 B.n426 10.6151
R588 B.n426 B.n34 10.6151
R589 B.n422 B.n34 10.6151
R590 B.n422 B.n421 10.6151
R591 B.n421 B.n420 10.6151
R592 B.n420 B.n36 10.6151
R593 B.n416 B.n36 10.6151
R594 B.n416 B.n415 10.6151
R595 B.n413 B.n40 10.6151
R596 B.n409 B.n40 10.6151
R597 B.n409 B.n408 10.6151
R598 B.n408 B.n407 10.6151
R599 B.n407 B.n42 10.6151
R600 B.n403 B.n42 10.6151
R601 B.n403 B.n402 10.6151
R602 B.n402 B.n401 10.6151
R603 B.n401 B.n44 10.6151
R604 B.n397 B.n44 10.6151
R605 B.n397 B.n396 10.6151
R606 B.n396 B.n395 10.6151
R607 B.n395 B.n46 10.6151
R608 B.n391 B.n46 10.6151
R609 B.n391 B.n390 10.6151
R610 B.n389 B.n48 10.6151
R611 B.n385 B.n48 10.6151
R612 B.n385 B.n384 10.6151
R613 B.n384 B.n383 10.6151
R614 B.n383 B.n50 10.6151
R615 B.n379 B.n50 10.6151
R616 B.n379 B.n378 10.6151
R617 B.n378 B.n377 10.6151
R618 B.n377 B.n52 10.6151
R619 B.n373 B.n52 10.6151
R620 B.n373 B.n372 10.6151
R621 B.n372 B.n371 10.6151
R622 B.n371 B.n54 10.6151
R623 B.n367 B.n54 10.6151
R624 B.n367 B.n366 10.6151
R625 B.n366 B.n365 10.6151
R626 B.n365 B.n56 10.6151
R627 B.n361 B.n56 10.6151
R628 B.n361 B.n360 10.6151
R629 B.n360 B.n359 10.6151
R630 B.n359 B.n58 10.6151
R631 B.n355 B.n58 10.6151
R632 B.n355 B.n354 10.6151
R633 B.n354 B.n353 10.6151
R634 B.n353 B.n60 10.6151
R635 B.n349 B.n60 10.6151
R636 B.n349 B.n348 10.6151
R637 B.n348 B.n347 10.6151
R638 B.n347 B.n62 10.6151
R639 B.n343 B.n62 10.6151
R640 B.n343 B.n342 10.6151
R641 B.n342 B.n341 10.6151
R642 B.n341 B.n64 10.6151
R643 B.n337 B.n64 10.6151
R644 B.n337 B.n336 10.6151
R645 B.n336 B.n335 10.6151
R646 B.n335 B.n66 10.6151
R647 B.n331 B.n66 10.6151
R648 B.n331 B.n330 10.6151
R649 B.n330 B.n329 10.6151
R650 B.n329 B.n68 10.6151
R651 B.n325 B.n68 10.6151
R652 B.n325 B.n324 10.6151
R653 B.n324 B.n323 10.6151
R654 B.n323 B.n70 10.6151
R655 B.n319 B.n70 10.6151
R656 B.n319 B.n318 10.6151
R657 B.n318 B.n317 10.6151
R658 B.n317 B.n72 10.6151
R659 B.n313 B.n72 10.6151
R660 B.n313 B.n312 10.6151
R661 B.n312 B.n311 10.6151
R662 B.n311 B.n74 10.6151
R663 B.n307 B.n74 10.6151
R664 B.n307 B.n306 10.6151
R665 B.n306 B.n305 10.6151
R666 B.n305 B.n76 10.6151
R667 B.n301 B.n76 10.6151
R668 B.n301 B.n300 10.6151
R669 B.n300 B.n299 10.6151
R670 B.n299 B.n78 10.6151
R671 B.n295 B.n78 10.6151
R672 B.n295 B.n294 10.6151
R673 B.n294 B.n293 10.6151
R674 B.n293 B.n80 10.6151
R675 B.n289 B.n80 10.6151
R676 B.n289 B.n288 10.6151
R677 B.n288 B.n287 10.6151
R678 B.n287 B.n82 10.6151
R679 B.n283 B.n82 10.6151
R680 B.n283 B.n282 10.6151
R681 B.n282 B.n281 10.6151
R682 B.n281 B.n84 10.6151
R683 B.n277 B.n84 10.6151
R684 B.n277 B.n276 10.6151
R685 B.n276 B.n275 10.6151
R686 B.n275 B.n86 10.6151
R687 B.n271 B.n86 10.6151
R688 B.n271 B.n270 10.6151
R689 B.n270 B.n269 10.6151
R690 B.n269 B.n88 10.6151
R691 B.n265 B.n88 10.6151
R692 B.n265 B.n264 10.6151
R693 B.n264 B.n263 10.6151
R694 B.n263 B.n90 10.6151
R695 B.n134 B.n1 10.6151
R696 B.n135 B.n134 10.6151
R697 B.n135 B.n132 10.6151
R698 B.n139 B.n132 10.6151
R699 B.n140 B.n139 10.6151
R700 B.n141 B.n140 10.6151
R701 B.n141 B.n130 10.6151
R702 B.n145 B.n130 10.6151
R703 B.n146 B.n145 10.6151
R704 B.n147 B.n146 10.6151
R705 B.n147 B.n128 10.6151
R706 B.n151 B.n128 10.6151
R707 B.n152 B.n151 10.6151
R708 B.n153 B.n152 10.6151
R709 B.n153 B.n126 10.6151
R710 B.n157 B.n126 10.6151
R711 B.n158 B.n157 10.6151
R712 B.n159 B.n158 10.6151
R713 B.n159 B.n124 10.6151
R714 B.n163 B.n124 10.6151
R715 B.n164 B.n163 10.6151
R716 B.n165 B.n164 10.6151
R717 B.n165 B.n122 10.6151
R718 B.n169 B.n122 10.6151
R719 B.n170 B.n169 10.6151
R720 B.n171 B.n170 10.6151
R721 B.n171 B.n120 10.6151
R722 B.n175 B.n120 10.6151
R723 B.n176 B.n175 10.6151
R724 B.n177 B.n176 10.6151
R725 B.n177 B.n118 10.6151
R726 B.n181 B.n118 10.6151
R727 B.n182 B.n181 10.6151
R728 B.n183 B.n182 10.6151
R729 B.n183 B.n116 10.6151
R730 B.n187 B.n116 10.6151
R731 B.n188 B.n187 10.6151
R732 B.n189 B.n188 10.6151
R733 B.n189 B.n114 10.6151
R734 B.n193 B.n114 10.6151
R735 B.n194 B.n193 10.6151
R736 B.n195 B.n112 10.6151
R737 B.n199 B.n112 10.6151
R738 B.n200 B.n199 10.6151
R739 B.n201 B.n200 10.6151
R740 B.n201 B.n110 10.6151
R741 B.n205 B.n110 10.6151
R742 B.n206 B.n205 10.6151
R743 B.n207 B.n206 10.6151
R744 B.n207 B.n108 10.6151
R745 B.n211 B.n108 10.6151
R746 B.n212 B.n211 10.6151
R747 B.n213 B.n212 10.6151
R748 B.n213 B.n106 10.6151
R749 B.n217 B.n106 10.6151
R750 B.n218 B.n217 10.6151
R751 B.n220 B.n102 10.6151
R752 B.n224 B.n102 10.6151
R753 B.n225 B.n224 10.6151
R754 B.n226 B.n225 10.6151
R755 B.n226 B.n100 10.6151
R756 B.n230 B.n100 10.6151
R757 B.n231 B.n230 10.6151
R758 B.n235 B.n231 10.6151
R759 B.n239 B.n98 10.6151
R760 B.n240 B.n239 10.6151
R761 B.n241 B.n240 10.6151
R762 B.n241 B.n96 10.6151
R763 B.n245 B.n96 10.6151
R764 B.n246 B.n245 10.6151
R765 B.n247 B.n246 10.6151
R766 B.n247 B.n94 10.6151
R767 B.n251 B.n94 10.6151
R768 B.n252 B.n251 10.6151
R769 B.n253 B.n252 10.6151
R770 B.n253 B.n92 10.6151
R771 B.n257 B.n92 10.6151
R772 B.n258 B.n257 10.6151
R773 B.n259 B.n258 10.6151
R774 B.n517 B.n0 8.11757
R775 B.n517 B.n1 8.11757
R776 B.n428 B.n427 6.5566
R777 B.n415 B.n414 6.5566
R778 B.n220 B.n219 6.5566
R779 B.n235 B.n234 6.5566
R780 B.n429 B.n428 4.05904
R781 B.n414 B.n413 4.05904
R782 B.n219 B.n218 4.05904
R783 B.n234 B.n98 4.05904
R784 VN.n29 VN.n28 179.406
R785 VN.n59 VN.n58 179.406
R786 VN.n57 VN.n30 161.3
R787 VN.n56 VN.n55 161.3
R788 VN.n54 VN.n31 161.3
R789 VN.n53 VN.n52 161.3
R790 VN.n50 VN.n32 161.3
R791 VN.n49 VN.n48 161.3
R792 VN.n47 VN.n33 161.3
R793 VN.n46 VN.n45 161.3
R794 VN.n43 VN.n34 161.3
R795 VN.n42 VN.n41 161.3
R796 VN.n40 VN.n35 161.3
R797 VN.n39 VN.n38 161.3
R798 VN.n27 VN.n0 161.3
R799 VN.n26 VN.n25 161.3
R800 VN.n24 VN.n1 161.3
R801 VN.n23 VN.n22 161.3
R802 VN.n20 VN.n2 161.3
R803 VN.n19 VN.n18 161.3
R804 VN.n17 VN.n3 161.3
R805 VN.n16 VN.n15 161.3
R806 VN.n13 VN.n4 161.3
R807 VN.n12 VN.n11 161.3
R808 VN.n10 VN.n5 161.3
R809 VN.n9 VN.n8 161.3
R810 VN.n6 VN.t9 80.1055
R811 VN.n36 VN.t4 80.1055
R812 VN.n7 VN.n6 56.8385
R813 VN.n37 VN.n36 56.8385
R814 VN.n12 VN.n5 56.5193
R815 VN.n19 VN.n3 56.5193
R816 VN.n42 VN.n35 56.5193
R817 VN.n49 VN.n33 56.5193
R818 VN.n26 VN.n1 56.0336
R819 VN.n56 VN.n31 56.0336
R820 VN.n7 VN.t5 48.3502
R821 VN.n14 VN.t3 48.3502
R822 VN.n21 VN.t6 48.3502
R823 VN.n28 VN.t0 48.3502
R824 VN.n37 VN.t2 48.3502
R825 VN.n44 VN.t8 48.3502
R826 VN.n51 VN.t7 48.3502
R827 VN.n58 VN.t1 48.3502
R828 VN VN.n59 41.366
R829 VN.n22 VN.n1 24.9531
R830 VN.n52 VN.n31 24.9531
R831 VN.n8 VN.n5 24.4675
R832 VN.n13 VN.n12 24.4675
R833 VN.n15 VN.n3 24.4675
R834 VN.n20 VN.n19 24.4675
R835 VN.n27 VN.n26 24.4675
R836 VN.n38 VN.n35 24.4675
R837 VN.n45 VN.n33 24.4675
R838 VN.n43 VN.n42 24.4675
R839 VN.n50 VN.n49 24.4675
R840 VN.n57 VN.n56 24.4675
R841 VN.n39 VN.n36 18.1515
R842 VN.n9 VN.n6 18.1515
R843 VN.n22 VN.n21 15.17
R844 VN.n52 VN.n51 15.17
R845 VN.n14 VN.n13 12.234
R846 VN.n15 VN.n14 12.234
R847 VN.n45 VN.n44 12.234
R848 VN.n44 VN.n43 12.234
R849 VN.n8 VN.n7 9.29796
R850 VN.n21 VN.n20 9.29796
R851 VN.n38 VN.n37 9.29796
R852 VN.n51 VN.n50 9.29796
R853 VN.n28 VN.n27 6.36192
R854 VN.n58 VN.n57 6.36192
R855 VN.n59 VN.n30 0.189894
R856 VN.n55 VN.n30 0.189894
R857 VN.n55 VN.n54 0.189894
R858 VN.n54 VN.n53 0.189894
R859 VN.n53 VN.n32 0.189894
R860 VN.n48 VN.n32 0.189894
R861 VN.n48 VN.n47 0.189894
R862 VN.n47 VN.n46 0.189894
R863 VN.n46 VN.n34 0.189894
R864 VN.n41 VN.n34 0.189894
R865 VN.n41 VN.n40 0.189894
R866 VN.n40 VN.n39 0.189894
R867 VN.n10 VN.n9 0.189894
R868 VN.n11 VN.n10 0.189894
R869 VN.n11 VN.n4 0.189894
R870 VN.n16 VN.n4 0.189894
R871 VN.n17 VN.n16 0.189894
R872 VN.n18 VN.n17 0.189894
R873 VN.n18 VN.n2 0.189894
R874 VN.n23 VN.n2 0.189894
R875 VN.n24 VN.n23 0.189894
R876 VN.n25 VN.n24 0.189894
R877 VN.n25 VN.n0 0.189894
R878 VN.n29 VN.n0 0.189894
R879 VN VN.n29 0.0516364
R880 VTAIL.n72 VTAIL.n62 756.745
R881 VTAIL.n12 VTAIL.n2 756.745
R882 VTAIL.n56 VTAIL.n46 756.745
R883 VTAIL.n36 VTAIL.n26 756.745
R884 VTAIL.n66 VTAIL.n65 585
R885 VTAIL.n71 VTAIL.n70 585
R886 VTAIL.n73 VTAIL.n72 585
R887 VTAIL.n6 VTAIL.n5 585
R888 VTAIL.n11 VTAIL.n10 585
R889 VTAIL.n13 VTAIL.n12 585
R890 VTAIL.n57 VTAIL.n56 585
R891 VTAIL.n55 VTAIL.n54 585
R892 VTAIL.n50 VTAIL.n49 585
R893 VTAIL.n37 VTAIL.n36 585
R894 VTAIL.n35 VTAIL.n34 585
R895 VTAIL.n30 VTAIL.n29 585
R896 VTAIL.n67 VTAIL.t16 336.901
R897 VTAIL.n7 VTAIL.t4 336.901
R898 VTAIL.n51 VTAIL.t7 336.901
R899 VTAIL.n31 VTAIL.t14 336.901
R900 VTAIL.n71 VTAIL.n65 171.744
R901 VTAIL.n72 VTAIL.n71 171.744
R902 VTAIL.n11 VTAIL.n5 171.744
R903 VTAIL.n12 VTAIL.n11 171.744
R904 VTAIL.n56 VTAIL.n55 171.744
R905 VTAIL.n55 VTAIL.n49 171.744
R906 VTAIL.n36 VTAIL.n35 171.744
R907 VTAIL.n35 VTAIL.n29 171.744
R908 VTAIL.n45 VTAIL.n44 113.305
R909 VTAIL.n43 VTAIL.n42 113.305
R910 VTAIL.n25 VTAIL.n24 113.305
R911 VTAIL.n23 VTAIL.n22 113.305
R912 VTAIL.n79 VTAIL.n78 113.305
R913 VTAIL.n1 VTAIL.n0 113.305
R914 VTAIL.n19 VTAIL.n18 113.305
R915 VTAIL.n21 VTAIL.n20 113.305
R916 VTAIL.t16 VTAIL.n65 85.8723
R917 VTAIL.t4 VTAIL.n5 85.8723
R918 VTAIL.t7 VTAIL.n49 85.8723
R919 VTAIL.t14 VTAIL.n29 85.8723
R920 VTAIL.n77 VTAIL.n76 34.3187
R921 VTAIL.n17 VTAIL.n16 34.3187
R922 VTAIL.n61 VTAIL.n60 34.3187
R923 VTAIL.n41 VTAIL.n40 34.3187
R924 VTAIL.n23 VTAIL.n21 18.4962
R925 VTAIL.n77 VTAIL.n61 16.8238
R926 VTAIL.n67 VTAIL.n66 16.193
R927 VTAIL.n7 VTAIL.n6 16.193
R928 VTAIL.n51 VTAIL.n50 16.193
R929 VTAIL.n31 VTAIL.n30 16.193
R930 VTAIL.n70 VTAIL.n69 12.8005
R931 VTAIL.n10 VTAIL.n9 12.8005
R932 VTAIL.n54 VTAIL.n53 12.8005
R933 VTAIL.n34 VTAIL.n33 12.8005
R934 VTAIL.n73 VTAIL.n64 12.0247
R935 VTAIL.n13 VTAIL.n4 12.0247
R936 VTAIL.n57 VTAIL.n48 12.0247
R937 VTAIL.n37 VTAIL.n28 12.0247
R938 VTAIL.n74 VTAIL.n62 11.249
R939 VTAIL.n14 VTAIL.n2 11.249
R940 VTAIL.n58 VTAIL.n46 11.249
R941 VTAIL.n38 VTAIL.n26 11.249
R942 VTAIL.n78 VTAIL.t12 10.064
R943 VTAIL.n78 VTAIL.t15 10.064
R944 VTAIL.n0 VTAIL.t18 10.064
R945 VTAIL.n0 VTAIL.t9 10.064
R946 VTAIL.n18 VTAIL.t19 10.064
R947 VTAIL.n18 VTAIL.t0 10.064
R948 VTAIL.n20 VTAIL.t3 10.064
R949 VTAIL.n20 VTAIL.t1 10.064
R950 VTAIL.n44 VTAIL.t6 10.064
R951 VTAIL.n44 VTAIL.t2 10.064
R952 VTAIL.n42 VTAIL.t5 10.064
R953 VTAIL.n42 VTAIL.t8 10.064
R954 VTAIL.n24 VTAIL.t11 10.064
R955 VTAIL.n24 VTAIL.t13 10.064
R956 VTAIL.n22 VTAIL.t10 10.064
R957 VTAIL.n22 VTAIL.t17 10.064
R958 VTAIL.n76 VTAIL.n75 9.45567
R959 VTAIL.n16 VTAIL.n15 9.45567
R960 VTAIL.n60 VTAIL.n59 9.45567
R961 VTAIL.n40 VTAIL.n39 9.45567
R962 VTAIL.n75 VTAIL.n74 9.3005
R963 VTAIL.n64 VTAIL.n63 9.3005
R964 VTAIL.n69 VTAIL.n68 9.3005
R965 VTAIL.n15 VTAIL.n14 9.3005
R966 VTAIL.n4 VTAIL.n3 9.3005
R967 VTAIL.n9 VTAIL.n8 9.3005
R968 VTAIL.n59 VTAIL.n58 9.3005
R969 VTAIL.n48 VTAIL.n47 9.3005
R970 VTAIL.n53 VTAIL.n52 9.3005
R971 VTAIL.n39 VTAIL.n38 9.3005
R972 VTAIL.n28 VTAIL.n27 9.3005
R973 VTAIL.n33 VTAIL.n32 9.3005
R974 VTAIL.n52 VTAIL.n51 3.91276
R975 VTAIL.n32 VTAIL.n31 3.91276
R976 VTAIL.n68 VTAIL.n67 3.91276
R977 VTAIL.n8 VTAIL.n7 3.91276
R978 VTAIL.n76 VTAIL.n62 2.71565
R979 VTAIL.n16 VTAIL.n2 2.71565
R980 VTAIL.n60 VTAIL.n46 2.71565
R981 VTAIL.n40 VTAIL.n26 2.71565
R982 VTAIL.n74 VTAIL.n73 1.93989
R983 VTAIL.n14 VTAIL.n13 1.93989
R984 VTAIL.n58 VTAIL.n57 1.93989
R985 VTAIL.n38 VTAIL.n37 1.93989
R986 VTAIL.n25 VTAIL.n23 1.67291
R987 VTAIL.n41 VTAIL.n25 1.67291
R988 VTAIL.n45 VTAIL.n43 1.67291
R989 VTAIL.n61 VTAIL.n45 1.67291
R990 VTAIL.n21 VTAIL.n19 1.67291
R991 VTAIL.n19 VTAIL.n17 1.67291
R992 VTAIL.n79 VTAIL.n77 1.67291
R993 VTAIL VTAIL.n1 1.313
R994 VTAIL.n43 VTAIL.n41 1.30653
R995 VTAIL.n17 VTAIL.n1 1.30653
R996 VTAIL.n70 VTAIL.n64 1.16414
R997 VTAIL.n10 VTAIL.n4 1.16414
R998 VTAIL.n54 VTAIL.n48 1.16414
R999 VTAIL.n34 VTAIL.n28 1.16414
R1000 VTAIL.n69 VTAIL.n66 0.388379
R1001 VTAIL.n9 VTAIL.n6 0.388379
R1002 VTAIL.n53 VTAIL.n50 0.388379
R1003 VTAIL.n33 VTAIL.n30 0.388379
R1004 VTAIL VTAIL.n79 0.360414
R1005 VTAIL.n68 VTAIL.n63 0.155672
R1006 VTAIL.n75 VTAIL.n63 0.155672
R1007 VTAIL.n8 VTAIL.n3 0.155672
R1008 VTAIL.n15 VTAIL.n3 0.155672
R1009 VTAIL.n59 VTAIL.n47 0.155672
R1010 VTAIL.n52 VTAIL.n47 0.155672
R1011 VTAIL.n39 VTAIL.n27 0.155672
R1012 VTAIL.n32 VTAIL.n27 0.155672
R1013 VDD2.n29 VDD2.n19 756.745
R1014 VDD2.n10 VDD2.n0 756.745
R1015 VDD2.n30 VDD2.n29 585
R1016 VDD2.n28 VDD2.n27 585
R1017 VDD2.n23 VDD2.n22 585
R1018 VDD2.n4 VDD2.n3 585
R1019 VDD2.n9 VDD2.n8 585
R1020 VDD2.n11 VDD2.n10 585
R1021 VDD2.n24 VDD2.t8 336.901
R1022 VDD2.n5 VDD2.t0 336.901
R1023 VDD2.n29 VDD2.n28 171.744
R1024 VDD2.n28 VDD2.n22 171.744
R1025 VDD2.n9 VDD2.n3 171.744
R1026 VDD2.n10 VDD2.n9 171.744
R1027 VDD2.n18 VDD2.n17 131.184
R1028 VDD2 VDD2.n37 131.18
R1029 VDD2.n36 VDD2.n35 129.984
R1030 VDD2.n16 VDD2.n15 129.984
R1031 VDD2.t8 VDD2.n22 85.8723
R1032 VDD2.t0 VDD2.n3 85.8723
R1033 VDD2.n16 VDD2.n14 52.6699
R1034 VDD2.n34 VDD2.n33 50.9975
R1035 VDD2.n34 VDD2.n18 34.4437
R1036 VDD2.n24 VDD2.n23 16.193
R1037 VDD2.n5 VDD2.n4 16.193
R1038 VDD2.n27 VDD2.n26 12.8005
R1039 VDD2.n8 VDD2.n7 12.8005
R1040 VDD2.n30 VDD2.n21 12.0247
R1041 VDD2.n11 VDD2.n2 12.0247
R1042 VDD2.n31 VDD2.n19 11.249
R1043 VDD2.n12 VDD2.n0 11.249
R1044 VDD2.n37 VDD2.t7 10.064
R1045 VDD2.n37 VDD2.t5 10.064
R1046 VDD2.n35 VDD2.t2 10.064
R1047 VDD2.n35 VDD2.t1 10.064
R1048 VDD2.n17 VDD2.t3 10.064
R1049 VDD2.n17 VDD2.t9 10.064
R1050 VDD2.n15 VDD2.t4 10.064
R1051 VDD2.n15 VDD2.t6 10.064
R1052 VDD2.n33 VDD2.n32 9.45567
R1053 VDD2.n14 VDD2.n13 9.45567
R1054 VDD2.n32 VDD2.n31 9.3005
R1055 VDD2.n21 VDD2.n20 9.3005
R1056 VDD2.n26 VDD2.n25 9.3005
R1057 VDD2.n13 VDD2.n12 9.3005
R1058 VDD2.n2 VDD2.n1 9.3005
R1059 VDD2.n7 VDD2.n6 9.3005
R1060 VDD2.n25 VDD2.n24 3.91276
R1061 VDD2.n6 VDD2.n5 3.91276
R1062 VDD2.n33 VDD2.n19 2.71565
R1063 VDD2.n14 VDD2.n0 2.71565
R1064 VDD2.n31 VDD2.n30 1.93989
R1065 VDD2.n12 VDD2.n11 1.93989
R1066 VDD2.n36 VDD2.n34 1.67291
R1067 VDD2.n27 VDD2.n21 1.16414
R1068 VDD2.n8 VDD2.n2 1.16414
R1069 VDD2 VDD2.n36 0.476793
R1070 VDD2.n26 VDD2.n23 0.388379
R1071 VDD2.n7 VDD2.n4 0.388379
R1072 VDD2.n18 VDD2.n16 0.363257
R1073 VDD2.n32 VDD2.n20 0.155672
R1074 VDD2.n25 VDD2.n20 0.155672
R1075 VDD2.n6 VDD2.n1 0.155672
R1076 VDD2.n13 VDD2.n1 0.155672
R1077 VP.n39 VP.n38 179.406
R1078 VP.n68 VP.n67 179.406
R1079 VP.n37 VP.n36 179.406
R1080 VP.n17 VP.n16 161.3
R1081 VP.n18 VP.n13 161.3
R1082 VP.n20 VP.n19 161.3
R1083 VP.n21 VP.n12 161.3
R1084 VP.n24 VP.n23 161.3
R1085 VP.n25 VP.n11 161.3
R1086 VP.n27 VP.n26 161.3
R1087 VP.n28 VP.n10 161.3
R1088 VP.n31 VP.n30 161.3
R1089 VP.n32 VP.n9 161.3
R1090 VP.n34 VP.n33 161.3
R1091 VP.n35 VP.n8 161.3
R1092 VP.n66 VP.n0 161.3
R1093 VP.n65 VP.n64 161.3
R1094 VP.n63 VP.n1 161.3
R1095 VP.n62 VP.n61 161.3
R1096 VP.n59 VP.n2 161.3
R1097 VP.n58 VP.n57 161.3
R1098 VP.n56 VP.n3 161.3
R1099 VP.n55 VP.n54 161.3
R1100 VP.n52 VP.n4 161.3
R1101 VP.n51 VP.n50 161.3
R1102 VP.n49 VP.n5 161.3
R1103 VP.n48 VP.n47 161.3
R1104 VP.n45 VP.n6 161.3
R1105 VP.n44 VP.n43 161.3
R1106 VP.n42 VP.n7 161.3
R1107 VP.n41 VP.n40 161.3
R1108 VP.n14 VP.t2 80.1055
R1109 VP.n15 VP.n14 56.8385
R1110 VP.n51 VP.n5 56.5193
R1111 VP.n58 VP.n3 56.5193
R1112 VP.n27 VP.n11 56.5193
R1113 VP.n20 VP.n13 56.5193
R1114 VP.n44 VP.n7 56.0336
R1115 VP.n65 VP.n1 56.0336
R1116 VP.n34 VP.n9 56.0336
R1117 VP.n39 VP.t7 48.3502
R1118 VP.n46 VP.t5 48.3502
R1119 VP.n53 VP.t1 48.3502
R1120 VP.n60 VP.t4 48.3502
R1121 VP.n67 VP.t0 48.3502
R1122 VP.n36 VP.t8 48.3502
R1123 VP.n29 VP.t3 48.3502
R1124 VP.n22 VP.t6 48.3502
R1125 VP.n15 VP.t9 48.3502
R1126 VP.n38 VP.n37 40.9853
R1127 VP.n45 VP.n44 24.9531
R1128 VP.n61 VP.n1 24.9531
R1129 VP.n30 VP.n9 24.9531
R1130 VP.n40 VP.n7 24.4675
R1131 VP.n47 VP.n5 24.4675
R1132 VP.n52 VP.n51 24.4675
R1133 VP.n54 VP.n3 24.4675
R1134 VP.n59 VP.n58 24.4675
R1135 VP.n66 VP.n65 24.4675
R1136 VP.n35 VP.n34 24.4675
R1137 VP.n28 VP.n27 24.4675
R1138 VP.n21 VP.n20 24.4675
R1139 VP.n23 VP.n11 24.4675
R1140 VP.n16 VP.n13 24.4675
R1141 VP.n17 VP.n14 18.1515
R1142 VP.n46 VP.n45 15.17
R1143 VP.n61 VP.n60 15.17
R1144 VP.n30 VP.n29 15.17
R1145 VP.n53 VP.n52 12.234
R1146 VP.n54 VP.n53 12.234
R1147 VP.n22 VP.n21 12.234
R1148 VP.n23 VP.n22 12.234
R1149 VP.n47 VP.n46 9.29796
R1150 VP.n60 VP.n59 9.29796
R1151 VP.n29 VP.n28 9.29796
R1152 VP.n16 VP.n15 9.29796
R1153 VP.n40 VP.n39 6.36192
R1154 VP.n67 VP.n66 6.36192
R1155 VP.n36 VP.n35 6.36192
R1156 VP.n18 VP.n17 0.189894
R1157 VP.n19 VP.n18 0.189894
R1158 VP.n19 VP.n12 0.189894
R1159 VP.n24 VP.n12 0.189894
R1160 VP.n25 VP.n24 0.189894
R1161 VP.n26 VP.n25 0.189894
R1162 VP.n26 VP.n10 0.189894
R1163 VP.n31 VP.n10 0.189894
R1164 VP.n32 VP.n31 0.189894
R1165 VP.n33 VP.n32 0.189894
R1166 VP.n33 VP.n8 0.189894
R1167 VP.n37 VP.n8 0.189894
R1168 VP.n41 VP.n38 0.189894
R1169 VP.n42 VP.n41 0.189894
R1170 VP.n43 VP.n42 0.189894
R1171 VP.n43 VP.n6 0.189894
R1172 VP.n48 VP.n6 0.189894
R1173 VP.n49 VP.n48 0.189894
R1174 VP.n50 VP.n49 0.189894
R1175 VP.n50 VP.n4 0.189894
R1176 VP.n55 VP.n4 0.189894
R1177 VP.n56 VP.n55 0.189894
R1178 VP.n57 VP.n56 0.189894
R1179 VP.n57 VP.n2 0.189894
R1180 VP.n62 VP.n2 0.189894
R1181 VP.n63 VP.n62 0.189894
R1182 VP.n64 VP.n63 0.189894
R1183 VP.n64 VP.n0 0.189894
R1184 VP.n68 VP.n0 0.189894
R1185 VP VP.n68 0.0516364
R1186 VDD1.n10 VDD1.n0 756.745
R1187 VDD1.n27 VDD1.n17 756.745
R1188 VDD1.n11 VDD1.n10 585
R1189 VDD1.n9 VDD1.n8 585
R1190 VDD1.n4 VDD1.n3 585
R1191 VDD1.n21 VDD1.n20 585
R1192 VDD1.n26 VDD1.n25 585
R1193 VDD1.n28 VDD1.n27 585
R1194 VDD1.n5 VDD1.t7 336.901
R1195 VDD1.n22 VDD1.t2 336.901
R1196 VDD1.n10 VDD1.n9 171.744
R1197 VDD1.n9 VDD1.n3 171.744
R1198 VDD1.n26 VDD1.n20 171.744
R1199 VDD1.n27 VDD1.n26 171.744
R1200 VDD1.n35 VDD1.n34 131.184
R1201 VDD1.n16 VDD1.n15 129.984
R1202 VDD1.n37 VDD1.n36 129.984
R1203 VDD1.n33 VDD1.n32 129.984
R1204 VDD1.t7 VDD1.n3 85.8723
R1205 VDD1.t2 VDD1.n20 85.8723
R1206 VDD1.n16 VDD1.n14 52.6699
R1207 VDD1.n33 VDD1.n31 52.6699
R1208 VDD1.n37 VDD1.n35 35.863
R1209 VDD1.n5 VDD1.n4 16.193
R1210 VDD1.n22 VDD1.n21 16.193
R1211 VDD1.n8 VDD1.n7 12.8005
R1212 VDD1.n25 VDD1.n24 12.8005
R1213 VDD1.n11 VDD1.n2 12.0247
R1214 VDD1.n28 VDD1.n19 12.0247
R1215 VDD1.n12 VDD1.n0 11.249
R1216 VDD1.n29 VDD1.n17 11.249
R1217 VDD1.n36 VDD1.t6 10.064
R1218 VDD1.n36 VDD1.t1 10.064
R1219 VDD1.n15 VDD1.t0 10.064
R1220 VDD1.n15 VDD1.t3 10.064
R1221 VDD1.n34 VDD1.t5 10.064
R1222 VDD1.n34 VDD1.t9 10.064
R1223 VDD1.n32 VDD1.t4 10.064
R1224 VDD1.n32 VDD1.t8 10.064
R1225 VDD1.n14 VDD1.n13 9.45567
R1226 VDD1.n31 VDD1.n30 9.45567
R1227 VDD1.n13 VDD1.n12 9.3005
R1228 VDD1.n2 VDD1.n1 9.3005
R1229 VDD1.n7 VDD1.n6 9.3005
R1230 VDD1.n30 VDD1.n29 9.3005
R1231 VDD1.n19 VDD1.n18 9.3005
R1232 VDD1.n24 VDD1.n23 9.3005
R1233 VDD1.n6 VDD1.n5 3.91276
R1234 VDD1.n23 VDD1.n22 3.91276
R1235 VDD1.n14 VDD1.n0 2.71565
R1236 VDD1.n31 VDD1.n17 2.71565
R1237 VDD1.n12 VDD1.n11 1.93989
R1238 VDD1.n29 VDD1.n28 1.93989
R1239 VDD1 VDD1.n37 1.19662
R1240 VDD1.n8 VDD1.n2 1.16414
R1241 VDD1.n25 VDD1.n19 1.16414
R1242 VDD1 VDD1.n16 0.476793
R1243 VDD1.n7 VDD1.n4 0.388379
R1244 VDD1.n24 VDD1.n21 0.388379
R1245 VDD1.n35 VDD1.n33 0.363257
R1246 VDD1.n13 VDD1.n1 0.155672
R1247 VDD1.n6 VDD1.n1 0.155672
R1248 VDD1.n23 VDD1.n18 0.155672
R1249 VDD1.n30 VDD1.n18 0.155672
C0 w_n3298_n1614# VDD1 1.78589f
C1 VDD1 VN 0.156182f
C2 B VDD2 1.4931f
C3 w_n3298_n1614# VN 6.58854f
C4 VDD1 VTAIL 5.54639f
C5 VP VDD1 3.20126f
C6 w_n3298_n1614# VTAIL 1.78962f
C7 VN VTAIL 3.6643f
C8 w_n3298_n1614# VP 7.0129f
C9 VDD2 VDD1 1.52999f
C10 VP VN 5.32168f
C11 B VDD1 1.41359f
C12 w_n3298_n1614# VDD2 1.87763f
C13 VP VTAIL 3.67849f
C14 VDD2 VN 2.89799f
C15 B w_n3298_n1614# 6.43666f
C16 B VN 0.945114f
C17 VDD2 VTAIL 5.59231f
C18 VP VDD2 0.462188f
C19 B VTAIL 1.43725f
C20 B VP 1.65618f
C21 VDD2 VSUBS 1.233828f
C22 VDD1 VSUBS 1.253824f
C23 VTAIL VSUBS 0.466499f
C24 VN VSUBS 5.79668f
C25 VP VSUBS 2.425778f
C26 B VSUBS 3.199646f
C27 w_n3298_n1614# VSUBS 67.318794f
C28 VDD1.n0 VSUBS 0.025176f
C29 VDD1.n1 VSUBS 0.023455f
C30 VDD1.n2 VSUBS 0.012603f
C31 VDD1.n3 VSUBS 0.022342f
C32 VDD1.n4 VSUBS 0.018391f
C33 VDD1.t7 VSUBS 0.066722f
C34 VDD1.n5 VSUBS 0.085756f
C35 VDD1.n6 VSUBS 0.239461f
C36 VDD1.n7 VSUBS 0.012603f
C37 VDD1.n8 VSUBS 0.013345f
C38 VDD1.n9 VSUBS 0.02979f
C39 VDD1.n10 VSUBS 0.070091f
C40 VDD1.n11 VSUBS 0.013345f
C41 VDD1.n12 VSUBS 0.012603f
C42 VDD1.n13 VSUBS 0.057738f
C43 VDD1.n14 VSUBS 0.056944f
C44 VDD1.t0 VSUBS 0.059866f
C45 VDD1.t3 VSUBS 0.059866f
C46 VDD1.n15 VSUBS 0.323746f
C47 VDD1.n16 VSUBS 0.636025f
C48 VDD1.n17 VSUBS 0.025176f
C49 VDD1.n18 VSUBS 0.023455f
C50 VDD1.n19 VSUBS 0.012603f
C51 VDD1.n20 VSUBS 0.022342f
C52 VDD1.n21 VSUBS 0.018391f
C53 VDD1.t2 VSUBS 0.066722f
C54 VDD1.n22 VSUBS 0.085756f
C55 VDD1.n23 VSUBS 0.239461f
C56 VDD1.n24 VSUBS 0.012603f
C57 VDD1.n25 VSUBS 0.013345f
C58 VDD1.n26 VSUBS 0.02979f
C59 VDD1.n27 VSUBS 0.070091f
C60 VDD1.n28 VSUBS 0.013345f
C61 VDD1.n29 VSUBS 0.012603f
C62 VDD1.n30 VSUBS 0.057738f
C63 VDD1.n31 VSUBS 0.056944f
C64 VDD1.t4 VSUBS 0.059866f
C65 VDD1.t8 VSUBS 0.059866f
C66 VDD1.n32 VSUBS 0.323745f
C67 VDD1.n33 VSUBS 0.628944f
C68 VDD1.t5 VSUBS 0.059866f
C69 VDD1.t9 VSUBS 0.059866f
C70 VDD1.n34 VSUBS 0.328611f
C71 VDD1.n35 VSUBS 1.951f
C72 VDD1.t6 VSUBS 0.059866f
C73 VDD1.t1 VSUBS 0.059866f
C74 VDD1.n36 VSUBS 0.323745f
C75 VDD1.n37 VSUBS 2.05813f
C76 VP.n0 VSUBS 0.053752f
C77 VP.t0 VSUBS 0.702525f
C78 VP.n1 VSUBS 0.064179f
C79 VP.n2 VSUBS 0.053752f
C80 VP.t4 VSUBS 0.702525f
C81 VP.n3 VSUBS 0.073975f
C82 VP.n4 VSUBS 0.053752f
C83 VP.t1 VSUBS 0.702525f
C84 VP.n5 VSUBS 0.082962f
C85 VP.n6 VSUBS 0.053752f
C86 VP.t5 VSUBS 0.702525f
C87 VP.n7 VSUBS 0.091817f
C88 VP.n8 VSUBS 0.053752f
C89 VP.t8 VSUBS 0.702525f
C90 VP.n9 VSUBS 0.064179f
C91 VP.n10 VSUBS 0.053752f
C92 VP.t3 VSUBS 0.702525f
C93 VP.n11 VSUBS 0.073975f
C94 VP.n12 VSUBS 0.053752f
C95 VP.t6 VSUBS 0.702525f
C96 VP.n13 VSUBS 0.082962f
C97 VP.t2 VSUBS 0.912571f
C98 VP.n14 VSUBS 0.419801f
C99 VP.t9 VSUBS 0.702525f
C100 VP.n15 VSUBS 0.410347f
C101 VP.n16 VSUBS 0.069516f
C102 VP.n17 VSUBS 0.341571f
C103 VP.n18 VSUBS 0.053752f
C104 VP.n19 VSUBS 0.053752f
C105 VP.n20 VSUBS 0.073975f
C106 VP.n21 VSUBS 0.075451f
C107 VP.n22 VSUBS 0.310582f
C108 VP.n23 VSUBS 0.075451f
C109 VP.n24 VSUBS 0.053752f
C110 VP.n25 VSUBS 0.053752f
C111 VP.n26 VSUBS 0.053752f
C112 VP.n27 VSUBS 0.082962f
C113 VP.n28 VSUBS 0.069516f
C114 VP.n29 VSUBS 0.310582f
C115 VP.n30 VSUBS 0.082327f
C116 VP.n31 VSUBS 0.053752f
C117 VP.n32 VSUBS 0.053752f
C118 VP.n33 VSUBS 0.053752f
C119 VP.n34 VSUBS 0.091817f
C120 VP.n35 VSUBS 0.063581f
C121 VP.n36 VSUBS 0.421998f
C122 VP.n37 VSUBS 2.14189f
C123 VP.n38 VSUBS 2.18903f
C124 VP.t7 VSUBS 0.702525f
C125 VP.n39 VSUBS 0.421998f
C126 VP.n40 VSUBS 0.063581f
C127 VP.n41 VSUBS 0.053752f
C128 VP.n42 VSUBS 0.053752f
C129 VP.n43 VSUBS 0.053752f
C130 VP.n44 VSUBS 0.064179f
C131 VP.n45 VSUBS 0.082327f
C132 VP.n46 VSUBS 0.310582f
C133 VP.n47 VSUBS 0.069516f
C134 VP.n48 VSUBS 0.053752f
C135 VP.n49 VSUBS 0.053752f
C136 VP.n50 VSUBS 0.053752f
C137 VP.n51 VSUBS 0.073975f
C138 VP.n52 VSUBS 0.075451f
C139 VP.n53 VSUBS 0.310582f
C140 VP.n54 VSUBS 0.075451f
C141 VP.n55 VSUBS 0.053752f
C142 VP.n56 VSUBS 0.053752f
C143 VP.n57 VSUBS 0.053752f
C144 VP.n58 VSUBS 0.082962f
C145 VP.n59 VSUBS 0.069516f
C146 VP.n60 VSUBS 0.310582f
C147 VP.n61 VSUBS 0.082327f
C148 VP.n62 VSUBS 0.053752f
C149 VP.n63 VSUBS 0.053752f
C150 VP.n64 VSUBS 0.053752f
C151 VP.n65 VSUBS 0.091817f
C152 VP.n66 VSUBS 0.063581f
C153 VP.n67 VSUBS 0.421998f
C154 VP.n68 VSUBS 0.054162f
C155 VDD2.n0 VSUBS 0.024845f
C156 VDD2.n1 VSUBS 0.023146f
C157 VDD2.n2 VSUBS 0.012438f
C158 VDD2.n3 VSUBS 0.022048f
C159 VDD2.n4 VSUBS 0.018149f
C160 VDD2.t0 VSUBS 0.065844f
C161 VDD2.n5 VSUBS 0.084627f
C162 VDD2.n6 VSUBS 0.236309f
C163 VDD2.n7 VSUBS 0.012438f
C164 VDD2.n8 VSUBS 0.013169f
C165 VDD2.n9 VSUBS 0.029398f
C166 VDD2.n10 VSUBS 0.069168f
C167 VDD2.n11 VSUBS 0.013169f
C168 VDD2.n12 VSUBS 0.012438f
C169 VDD2.n13 VSUBS 0.056979f
C170 VDD2.n14 VSUBS 0.056194f
C171 VDD2.t4 VSUBS 0.059078f
C172 VDD2.t6 VSUBS 0.059078f
C173 VDD2.n15 VSUBS 0.319484f
C174 VDD2.n16 VSUBS 0.620666f
C175 VDD2.t3 VSUBS 0.059078f
C176 VDD2.t9 VSUBS 0.059078f
C177 VDD2.n17 VSUBS 0.324286f
C178 VDD2.n18 VSUBS 1.83927f
C179 VDD2.n19 VSUBS 0.024845f
C180 VDD2.n20 VSUBS 0.023146f
C181 VDD2.n21 VSUBS 0.012438f
C182 VDD2.n22 VSUBS 0.022048f
C183 VDD2.n23 VSUBS 0.018149f
C184 VDD2.t8 VSUBS 0.065844f
C185 VDD2.n24 VSUBS 0.084627f
C186 VDD2.n25 VSUBS 0.236309f
C187 VDD2.n26 VSUBS 0.012438f
C188 VDD2.n27 VSUBS 0.013169f
C189 VDD2.n28 VSUBS 0.029398f
C190 VDD2.n29 VSUBS 0.069168f
C191 VDD2.n30 VSUBS 0.013169f
C192 VDD2.n31 VSUBS 0.012438f
C193 VDD2.n32 VSUBS 0.056979f
C194 VDD2.n33 VSUBS 0.050755f
C195 VDD2.n34 VSUBS 1.67808f
C196 VDD2.t2 VSUBS 0.059078f
C197 VDD2.t1 VSUBS 0.059078f
C198 VDD2.n35 VSUBS 0.319485f
C199 VDD2.n36 VSUBS 0.461801f
C200 VDD2.t7 VSUBS 0.059078f
C201 VDD2.t5 VSUBS 0.059078f
C202 VDD2.n37 VSUBS 0.324269f
C203 VTAIL.t18 VSUBS 0.078705f
C204 VTAIL.t9 VSUBS 0.078705f
C205 VTAIL.n0 VSUBS 0.36735f
C206 VTAIL.n1 VSUBS 0.678263f
C207 VTAIL.n2 VSUBS 0.033099f
C208 VTAIL.n3 VSUBS 0.030835f
C209 VTAIL.n4 VSUBS 0.016569f
C210 VTAIL.n5 VSUBS 0.029373f
C211 VTAIL.n6 VSUBS 0.024179f
C212 VTAIL.t4 VSUBS 0.087718f
C213 VTAIL.n7 VSUBS 0.112742f
C214 VTAIL.n8 VSUBS 0.314815f
C215 VTAIL.n9 VSUBS 0.016569f
C216 VTAIL.n10 VSUBS 0.017544f
C217 VTAIL.n11 VSUBS 0.039164f
C218 VTAIL.n12 VSUBS 0.092147f
C219 VTAIL.n13 VSUBS 0.017544f
C220 VTAIL.n14 VSUBS 0.016569f
C221 VTAIL.n15 VSUBS 0.075908f
C222 VTAIL.n16 VSUBS 0.04636f
C223 VTAIL.n17 VSUBS 0.324887f
C224 VTAIL.t19 VSUBS 0.078705f
C225 VTAIL.t0 VSUBS 0.078705f
C226 VTAIL.n18 VSUBS 0.36735f
C227 VTAIL.n19 VSUBS 0.750426f
C228 VTAIL.t3 VSUBS 0.078705f
C229 VTAIL.t1 VSUBS 0.078705f
C230 VTAIL.n20 VSUBS 0.36735f
C231 VTAIL.n21 VSUBS 1.61211f
C232 VTAIL.t10 VSUBS 0.078705f
C233 VTAIL.t17 VSUBS 0.078705f
C234 VTAIL.n22 VSUBS 0.367352f
C235 VTAIL.n23 VSUBS 1.61211f
C236 VTAIL.t11 VSUBS 0.078705f
C237 VTAIL.t13 VSUBS 0.078705f
C238 VTAIL.n24 VSUBS 0.367352f
C239 VTAIL.n25 VSUBS 0.750424f
C240 VTAIL.n26 VSUBS 0.033099f
C241 VTAIL.n27 VSUBS 0.030835f
C242 VTAIL.n28 VSUBS 0.016569f
C243 VTAIL.n29 VSUBS 0.029373f
C244 VTAIL.n30 VSUBS 0.024179f
C245 VTAIL.t14 VSUBS 0.087718f
C246 VTAIL.n31 VSUBS 0.112742f
C247 VTAIL.n32 VSUBS 0.314815f
C248 VTAIL.n33 VSUBS 0.016569f
C249 VTAIL.n34 VSUBS 0.017544f
C250 VTAIL.n35 VSUBS 0.039164f
C251 VTAIL.n36 VSUBS 0.092147f
C252 VTAIL.n37 VSUBS 0.017544f
C253 VTAIL.n38 VSUBS 0.016569f
C254 VTAIL.n39 VSUBS 0.075908f
C255 VTAIL.n40 VSUBS 0.04636f
C256 VTAIL.n41 VSUBS 0.324887f
C257 VTAIL.t5 VSUBS 0.078705f
C258 VTAIL.t8 VSUBS 0.078705f
C259 VTAIL.n42 VSUBS 0.367352f
C260 VTAIL.n43 VSUBS 0.714021f
C261 VTAIL.t6 VSUBS 0.078705f
C262 VTAIL.t2 VSUBS 0.078705f
C263 VTAIL.n44 VSUBS 0.367352f
C264 VTAIL.n45 VSUBS 0.750424f
C265 VTAIL.n46 VSUBS 0.033099f
C266 VTAIL.n47 VSUBS 0.030835f
C267 VTAIL.n48 VSUBS 0.016569f
C268 VTAIL.n49 VSUBS 0.029373f
C269 VTAIL.n50 VSUBS 0.024179f
C270 VTAIL.t7 VSUBS 0.087718f
C271 VTAIL.n51 VSUBS 0.112742f
C272 VTAIL.n52 VSUBS 0.314815f
C273 VTAIL.n53 VSUBS 0.016569f
C274 VTAIL.n54 VSUBS 0.017544f
C275 VTAIL.n55 VSUBS 0.039164f
C276 VTAIL.n56 VSUBS 0.092147f
C277 VTAIL.n57 VSUBS 0.017544f
C278 VTAIL.n58 VSUBS 0.016569f
C279 VTAIL.n59 VSUBS 0.075908f
C280 VTAIL.n60 VSUBS 0.04636f
C281 VTAIL.n61 VSUBS 1.05681f
C282 VTAIL.n62 VSUBS 0.033099f
C283 VTAIL.n63 VSUBS 0.030835f
C284 VTAIL.n64 VSUBS 0.016569f
C285 VTAIL.n65 VSUBS 0.029373f
C286 VTAIL.n66 VSUBS 0.024179f
C287 VTAIL.t16 VSUBS 0.087718f
C288 VTAIL.n67 VSUBS 0.112742f
C289 VTAIL.n68 VSUBS 0.314815f
C290 VTAIL.n69 VSUBS 0.016569f
C291 VTAIL.n70 VSUBS 0.017544f
C292 VTAIL.n71 VSUBS 0.039164f
C293 VTAIL.n72 VSUBS 0.092147f
C294 VTAIL.n73 VSUBS 0.017544f
C295 VTAIL.n74 VSUBS 0.016569f
C296 VTAIL.n75 VSUBS 0.075908f
C297 VTAIL.n76 VSUBS 0.04636f
C298 VTAIL.n77 VSUBS 1.05681f
C299 VTAIL.t12 VSUBS 0.078705f
C300 VTAIL.t15 VSUBS 0.078705f
C301 VTAIL.n78 VSUBS 0.36735f
C302 VTAIL.n79 VSUBS 0.620019f
C303 VN.n0 VSUBS 0.05159f
C304 VN.t0 VSUBS 0.674259f
C305 VN.n1 VSUBS 0.061597f
C306 VN.n2 VSUBS 0.05159f
C307 VN.t6 VSUBS 0.674259f
C308 VN.n3 VSUBS 0.070999f
C309 VN.n4 VSUBS 0.05159f
C310 VN.t3 VSUBS 0.674259f
C311 VN.n5 VSUBS 0.079624f
C312 VN.t9 VSUBS 0.875854f
C313 VN.n6 VSUBS 0.40291f
C314 VN.t5 VSUBS 0.674259f
C315 VN.n7 VSUBS 0.393837f
C316 VN.n8 VSUBS 0.066719f
C317 VN.n9 VSUBS 0.327828f
C318 VN.n10 VSUBS 0.05159f
C319 VN.n11 VSUBS 0.05159f
C320 VN.n12 VSUBS 0.070999f
C321 VN.n13 VSUBS 0.072415f
C322 VN.n14 VSUBS 0.298086f
C323 VN.n15 VSUBS 0.072415f
C324 VN.n16 VSUBS 0.05159f
C325 VN.n17 VSUBS 0.05159f
C326 VN.n18 VSUBS 0.05159f
C327 VN.n19 VSUBS 0.079624f
C328 VN.n20 VSUBS 0.066719f
C329 VN.n21 VSUBS 0.298086f
C330 VN.n22 VSUBS 0.079014f
C331 VN.n23 VSUBS 0.05159f
C332 VN.n24 VSUBS 0.05159f
C333 VN.n25 VSUBS 0.05159f
C334 VN.n26 VSUBS 0.088123f
C335 VN.n27 VSUBS 0.061022f
C336 VN.n28 VSUBS 0.405018f
C337 VN.n29 VSUBS 0.051983f
C338 VN.n30 VSUBS 0.05159f
C339 VN.t1 VSUBS 0.674259f
C340 VN.n31 VSUBS 0.061597f
C341 VN.n32 VSUBS 0.05159f
C342 VN.t7 VSUBS 0.674259f
C343 VN.n33 VSUBS 0.070999f
C344 VN.n34 VSUBS 0.05159f
C345 VN.t8 VSUBS 0.674259f
C346 VN.n35 VSUBS 0.079624f
C347 VN.t4 VSUBS 0.875854f
C348 VN.n36 VSUBS 0.40291f
C349 VN.t2 VSUBS 0.674259f
C350 VN.n37 VSUBS 0.393837f
C351 VN.n38 VSUBS 0.066719f
C352 VN.n39 VSUBS 0.327828f
C353 VN.n40 VSUBS 0.05159f
C354 VN.n41 VSUBS 0.05159f
C355 VN.n42 VSUBS 0.070999f
C356 VN.n43 VSUBS 0.072415f
C357 VN.n44 VSUBS 0.298086f
C358 VN.n45 VSUBS 0.072415f
C359 VN.n46 VSUBS 0.05159f
C360 VN.n47 VSUBS 0.05159f
C361 VN.n48 VSUBS 0.05159f
C362 VN.n49 VSUBS 0.079624f
C363 VN.n50 VSUBS 0.066719f
C364 VN.n51 VSUBS 0.298086f
C365 VN.n52 VSUBS 0.079014f
C366 VN.n53 VSUBS 0.05159f
C367 VN.n54 VSUBS 0.05159f
C368 VN.n55 VSUBS 0.05159f
C369 VN.n56 VSUBS 0.088123f
C370 VN.n57 VSUBS 0.061022f
C371 VN.n58 VSUBS 0.405018f
C372 VN.n59 VSUBS 2.08963f
C373 B.n0 VSUBS 0.006599f
C374 B.n1 VSUBS 0.006599f
C375 B.n2 VSUBS 0.00976f
C376 B.n3 VSUBS 0.007479f
C377 B.n4 VSUBS 0.007479f
C378 B.n5 VSUBS 0.007479f
C379 B.n6 VSUBS 0.007479f
C380 B.n7 VSUBS 0.007479f
C381 B.n8 VSUBS 0.007479f
C382 B.n9 VSUBS 0.007479f
C383 B.n10 VSUBS 0.007479f
C384 B.n11 VSUBS 0.007479f
C385 B.n12 VSUBS 0.007479f
C386 B.n13 VSUBS 0.007479f
C387 B.n14 VSUBS 0.007479f
C388 B.n15 VSUBS 0.007479f
C389 B.n16 VSUBS 0.007479f
C390 B.n17 VSUBS 0.007479f
C391 B.n18 VSUBS 0.007479f
C392 B.n19 VSUBS 0.007479f
C393 B.n20 VSUBS 0.007479f
C394 B.n21 VSUBS 0.007479f
C395 B.n22 VSUBS 0.007479f
C396 B.n23 VSUBS 0.017498f
C397 B.n24 VSUBS 0.007479f
C398 B.n25 VSUBS 0.007479f
C399 B.n26 VSUBS 0.007479f
C400 B.n27 VSUBS 0.007479f
C401 B.n28 VSUBS 0.007479f
C402 B.n29 VSUBS 0.007479f
C403 B.n30 VSUBS 0.007479f
C404 B.n31 VSUBS 0.007479f
C405 B.t4 VSUBS 0.050891f
C406 B.t5 VSUBS 0.063702f
C407 B.t3 VSUBS 0.264832f
C408 B.n32 VSUBS 0.114184f
C409 B.n33 VSUBS 0.10048f
C410 B.n34 VSUBS 0.007479f
C411 B.n35 VSUBS 0.007479f
C412 B.n36 VSUBS 0.007479f
C413 B.n37 VSUBS 0.007479f
C414 B.t7 VSUBS 0.050891f
C415 B.t8 VSUBS 0.063702f
C416 B.t6 VSUBS 0.264832f
C417 B.n38 VSUBS 0.114183f
C418 B.n39 VSUBS 0.100479f
C419 B.n40 VSUBS 0.007479f
C420 B.n41 VSUBS 0.007479f
C421 B.n42 VSUBS 0.007479f
C422 B.n43 VSUBS 0.007479f
C423 B.n44 VSUBS 0.007479f
C424 B.n45 VSUBS 0.007479f
C425 B.n46 VSUBS 0.007479f
C426 B.n47 VSUBS 0.017498f
C427 B.n48 VSUBS 0.007479f
C428 B.n49 VSUBS 0.007479f
C429 B.n50 VSUBS 0.007479f
C430 B.n51 VSUBS 0.007479f
C431 B.n52 VSUBS 0.007479f
C432 B.n53 VSUBS 0.007479f
C433 B.n54 VSUBS 0.007479f
C434 B.n55 VSUBS 0.007479f
C435 B.n56 VSUBS 0.007479f
C436 B.n57 VSUBS 0.007479f
C437 B.n58 VSUBS 0.007479f
C438 B.n59 VSUBS 0.007479f
C439 B.n60 VSUBS 0.007479f
C440 B.n61 VSUBS 0.007479f
C441 B.n62 VSUBS 0.007479f
C442 B.n63 VSUBS 0.007479f
C443 B.n64 VSUBS 0.007479f
C444 B.n65 VSUBS 0.007479f
C445 B.n66 VSUBS 0.007479f
C446 B.n67 VSUBS 0.007479f
C447 B.n68 VSUBS 0.007479f
C448 B.n69 VSUBS 0.007479f
C449 B.n70 VSUBS 0.007479f
C450 B.n71 VSUBS 0.007479f
C451 B.n72 VSUBS 0.007479f
C452 B.n73 VSUBS 0.007479f
C453 B.n74 VSUBS 0.007479f
C454 B.n75 VSUBS 0.007479f
C455 B.n76 VSUBS 0.007479f
C456 B.n77 VSUBS 0.007479f
C457 B.n78 VSUBS 0.007479f
C458 B.n79 VSUBS 0.007479f
C459 B.n80 VSUBS 0.007479f
C460 B.n81 VSUBS 0.007479f
C461 B.n82 VSUBS 0.007479f
C462 B.n83 VSUBS 0.007479f
C463 B.n84 VSUBS 0.007479f
C464 B.n85 VSUBS 0.007479f
C465 B.n86 VSUBS 0.007479f
C466 B.n87 VSUBS 0.007479f
C467 B.n88 VSUBS 0.007479f
C468 B.n89 VSUBS 0.007479f
C469 B.n90 VSUBS 0.017938f
C470 B.n91 VSUBS 0.007479f
C471 B.n92 VSUBS 0.007479f
C472 B.n93 VSUBS 0.007479f
C473 B.n94 VSUBS 0.007479f
C474 B.n95 VSUBS 0.007479f
C475 B.n96 VSUBS 0.007479f
C476 B.n97 VSUBS 0.007479f
C477 B.n98 VSUBS 0.005169f
C478 B.n99 VSUBS 0.007479f
C479 B.n100 VSUBS 0.007479f
C480 B.n101 VSUBS 0.007479f
C481 B.n102 VSUBS 0.007479f
C482 B.n103 VSUBS 0.007479f
C483 B.t11 VSUBS 0.050891f
C484 B.t10 VSUBS 0.063702f
C485 B.t9 VSUBS 0.264832f
C486 B.n104 VSUBS 0.114184f
C487 B.n105 VSUBS 0.10048f
C488 B.n106 VSUBS 0.007479f
C489 B.n107 VSUBS 0.007479f
C490 B.n108 VSUBS 0.007479f
C491 B.n109 VSUBS 0.007479f
C492 B.n110 VSUBS 0.007479f
C493 B.n111 VSUBS 0.007479f
C494 B.n112 VSUBS 0.007479f
C495 B.n113 VSUBS 0.017036f
C496 B.n114 VSUBS 0.007479f
C497 B.n115 VSUBS 0.007479f
C498 B.n116 VSUBS 0.007479f
C499 B.n117 VSUBS 0.007479f
C500 B.n118 VSUBS 0.007479f
C501 B.n119 VSUBS 0.007479f
C502 B.n120 VSUBS 0.007479f
C503 B.n121 VSUBS 0.007479f
C504 B.n122 VSUBS 0.007479f
C505 B.n123 VSUBS 0.007479f
C506 B.n124 VSUBS 0.007479f
C507 B.n125 VSUBS 0.007479f
C508 B.n126 VSUBS 0.007479f
C509 B.n127 VSUBS 0.007479f
C510 B.n128 VSUBS 0.007479f
C511 B.n129 VSUBS 0.007479f
C512 B.n130 VSUBS 0.007479f
C513 B.n131 VSUBS 0.007479f
C514 B.n132 VSUBS 0.007479f
C515 B.n133 VSUBS 0.007479f
C516 B.n134 VSUBS 0.007479f
C517 B.n135 VSUBS 0.007479f
C518 B.n136 VSUBS 0.007479f
C519 B.n137 VSUBS 0.007479f
C520 B.n138 VSUBS 0.007479f
C521 B.n139 VSUBS 0.007479f
C522 B.n140 VSUBS 0.007479f
C523 B.n141 VSUBS 0.007479f
C524 B.n142 VSUBS 0.007479f
C525 B.n143 VSUBS 0.007479f
C526 B.n144 VSUBS 0.007479f
C527 B.n145 VSUBS 0.007479f
C528 B.n146 VSUBS 0.007479f
C529 B.n147 VSUBS 0.007479f
C530 B.n148 VSUBS 0.007479f
C531 B.n149 VSUBS 0.007479f
C532 B.n150 VSUBS 0.007479f
C533 B.n151 VSUBS 0.007479f
C534 B.n152 VSUBS 0.007479f
C535 B.n153 VSUBS 0.007479f
C536 B.n154 VSUBS 0.007479f
C537 B.n155 VSUBS 0.007479f
C538 B.n156 VSUBS 0.007479f
C539 B.n157 VSUBS 0.007479f
C540 B.n158 VSUBS 0.007479f
C541 B.n159 VSUBS 0.007479f
C542 B.n160 VSUBS 0.007479f
C543 B.n161 VSUBS 0.007479f
C544 B.n162 VSUBS 0.007479f
C545 B.n163 VSUBS 0.007479f
C546 B.n164 VSUBS 0.007479f
C547 B.n165 VSUBS 0.007479f
C548 B.n166 VSUBS 0.007479f
C549 B.n167 VSUBS 0.007479f
C550 B.n168 VSUBS 0.007479f
C551 B.n169 VSUBS 0.007479f
C552 B.n170 VSUBS 0.007479f
C553 B.n171 VSUBS 0.007479f
C554 B.n172 VSUBS 0.007479f
C555 B.n173 VSUBS 0.007479f
C556 B.n174 VSUBS 0.007479f
C557 B.n175 VSUBS 0.007479f
C558 B.n176 VSUBS 0.007479f
C559 B.n177 VSUBS 0.007479f
C560 B.n178 VSUBS 0.007479f
C561 B.n179 VSUBS 0.007479f
C562 B.n180 VSUBS 0.007479f
C563 B.n181 VSUBS 0.007479f
C564 B.n182 VSUBS 0.007479f
C565 B.n183 VSUBS 0.007479f
C566 B.n184 VSUBS 0.007479f
C567 B.n185 VSUBS 0.007479f
C568 B.n186 VSUBS 0.007479f
C569 B.n187 VSUBS 0.007479f
C570 B.n188 VSUBS 0.007479f
C571 B.n189 VSUBS 0.007479f
C572 B.n190 VSUBS 0.007479f
C573 B.n191 VSUBS 0.007479f
C574 B.n192 VSUBS 0.007479f
C575 B.n193 VSUBS 0.007479f
C576 B.n194 VSUBS 0.017036f
C577 B.n195 VSUBS 0.017498f
C578 B.n196 VSUBS 0.017498f
C579 B.n197 VSUBS 0.007479f
C580 B.n198 VSUBS 0.007479f
C581 B.n199 VSUBS 0.007479f
C582 B.n200 VSUBS 0.007479f
C583 B.n201 VSUBS 0.007479f
C584 B.n202 VSUBS 0.007479f
C585 B.n203 VSUBS 0.007479f
C586 B.n204 VSUBS 0.007479f
C587 B.n205 VSUBS 0.007479f
C588 B.n206 VSUBS 0.007479f
C589 B.n207 VSUBS 0.007479f
C590 B.n208 VSUBS 0.007479f
C591 B.n209 VSUBS 0.007479f
C592 B.n210 VSUBS 0.007479f
C593 B.n211 VSUBS 0.007479f
C594 B.n212 VSUBS 0.007479f
C595 B.n213 VSUBS 0.007479f
C596 B.n214 VSUBS 0.007479f
C597 B.n215 VSUBS 0.007479f
C598 B.n216 VSUBS 0.007479f
C599 B.n217 VSUBS 0.007479f
C600 B.n218 VSUBS 0.005169f
C601 B.n219 VSUBS 0.017328f
C602 B.n220 VSUBS 0.006049f
C603 B.n221 VSUBS 0.007479f
C604 B.n222 VSUBS 0.007479f
C605 B.n223 VSUBS 0.007479f
C606 B.n224 VSUBS 0.007479f
C607 B.n225 VSUBS 0.007479f
C608 B.n226 VSUBS 0.007479f
C609 B.n227 VSUBS 0.007479f
C610 B.n228 VSUBS 0.007479f
C611 B.n229 VSUBS 0.007479f
C612 B.n230 VSUBS 0.007479f
C613 B.n231 VSUBS 0.007479f
C614 B.t2 VSUBS 0.050891f
C615 B.t1 VSUBS 0.063702f
C616 B.t0 VSUBS 0.264832f
C617 B.n232 VSUBS 0.114183f
C618 B.n233 VSUBS 0.100479f
C619 B.n234 VSUBS 0.017328f
C620 B.n235 VSUBS 0.006049f
C621 B.n236 VSUBS 0.007479f
C622 B.n237 VSUBS 0.007479f
C623 B.n238 VSUBS 0.007479f
C624 B.n239 VSUBS 0.007479f
C625 B.n240 VSUBS 0.007479f
C626 B.n241 VSUBS 0.007479f
C627 B.n242 VSUBS 0.007479f
C628 B.n243 VSUBS 0.007479f
C629 B.n244 VSUBS 0.007479f
C630 B.n245 VSUBS 0.007479f
C631 B.n246 VSUBS 0.007479f
C632 B.n247 VSUBS 0.007479f
C633 B.n248 VSUBS 0.007479f
C634 B.n249 VSUBS 0.007479f
C635 B.n250 VSUBS 0.007479f
C636 B.n251 VSUBS 0.007479f
C637 B.n252 VSUBS 0.007479f
C638 B.n253 VSUBS 0.007479f
C639 B.n254 VSUBS 0.007479f
C640 B.n255 VSUBS 0.007479f
C641 B.n256 VSUBS 0.007479f
C642 B.n257 VSUBS 0.007479f
C643 B.n258 VSUBS 0.007479f
C644 B.n259 VSUBS 0.016596f
C645 B.n260 VSUBS 0.017498f
C646 B.n261 VSUBS 0.017036f
C647 B.n262 VSUBS 0.007479f
C648 B.n263 VSUBS 0.007479f
C649 B.n264 VSUBS 0.007479f
C650 B.n265 VSUBS 0.007479f
C651 B.n266 VSUBS 0.007479f
C652 B.n267 VSUBS 0.007479f
C653 B.n268 VSUBS 0.007479f
C654 B.n269 VSUBS 0.007479f
C655 B.n270 VSUBS 0.007479f
C656 B.n271 VSUBS 0.007479f
C657 B.n272 VSUBS 0.007479f
C658 B.n273 VSUBS 0.007479f
C659 B.n274 VSUBS 0.007479f
C660 B.n275 VSUBS 0.007479f
C661 B.n276 VSUBS 0.007479f
C662 B.n277 VSUBS 0.007479f
C663 B.n278 VSUBS 0.007479f
C664 B.n279 VSUBS 0.007479f
C665 B.n280 VSUBS 0.007479f
C666 B.n281 VSUBS 0.007479f
C667 B.n282 VSUBS 0.007479f
C668 B.n283 VSUBS 0.007479f
C669 B.n284 VSUBS 0.007479f
C670 B.n285 VSUBS 0.007479f
C671 B.n286 VSUBS 0.007479f
C672 B.n287 VSUBS 0.007479f
C673 B.n288 VSUBS 0.007479f
C674 B.n289 VSUBS 0.007479f
C675 B.n290 VSUBS 0.007479f
C676 B.n291 VSUBS 0.007479f
C677 B.n292 VSUBS 0.007479f
C678 B.n293 VSUBS 0.007479f
C679 B.n294 VSUBS 0.007479f
C680 B.n295 VSUBS 0.007479f
C681 B.n296 VSUBS 0.007479f
C682 B.n297 VSUBS 0.007479f
C683 B.n298 VSUBS 0.007479f
C684 B.n299 VSUBS 0.007479f
C685 B.n300 VSUBS 0.007479f
C686 B.n301 VSUBS 0.007479f
C687 B.n302 VSUBS 0.007479f
C688 B.n303 VSUBS 0.007479f
C689 B.n304 VSUBS 0.007479f
C690 B.n305 VSUBS 0.007479f
C691 B.n306 VSUBS 0.007479f
C692 B.n307 VSUBS 0.007479f
C693 B.n308 VSUBS 0.007479f
C694 B.n309 VSUBS 0.007479f
C695 B.n310 VSUBS 0.007479f
C696 B.n311 VSUBS 0.007479f
C697 B.n312 VSUBS 0.007479f
C698 B.n313 VSUBS 0.007479f
C699 B.n314 VSUBS 0.007479f
C700 B.n315 VSUBS 0.007479f
C701 B.n316 VSUBS 0.007479f
C702 B.n317 VSUBS 0.007479f
C703 B.n318 VSUBS 0.007479f
C704 B.n319 VSUBS 0.007479f
C705 B.n320 VSUBS 0.007479f
C706 B.n321 VSUBS 0.007479f
C707 B.n322 VSUBS 0.007479f
C708 B.n323 VSUBS 0.007479f
C709 B.n324 VSUBS 0.007479f
C710 B.n325 VSUBS 0.007479f
C711 B.n326 VSUBS 0.007479f
C712 B.n327 VSUBS 0.007479f
C713 B.n328 VSUBS 0.007479f
C714 B.n329 VSUBS 0.007479f
C715 B.n330 VSUBS 0.007479f
C716 B.n331 VSUBS 0.007479f
C717 B.n332 VSUBS 0.007479f
C718 B.n333 VSUBS 0.007479f
C719 B.n334 VSUBS 0.007479f
C720 B.n335 VSUBS 0.007479f
C721 B.n336 VSUBS 0.007479f
C722 B.n337 VSUBS 0.007479f
C723 B.n338 VSUBS 0.007479f
C724 B.n339 VSUBS 0.007479f
C725 B.n340 VSUBS 0.007479f
C726 B.n341 VSUBS 0.007479f
C727 B.n342 VSUBS 0.007479f
C728 B.n343 VSUBS 0.007479f
C729 B.n344 VSUBS 0.007479f
C730 B.n345 VSUBS 0.007479f
C731 B.n346 VSUBS 0.007479f
C732 B.n347 VSUBS 0.007479f
C733 B.n348 VSUBS 0.007479f
C734 B.n349 VSUBS 0.007479f
C735 B.n350 VSUBS 0.007479f
C736 B.n351 VSUBS 0.007479f
C737 B.n352 VSUBS 0.007479f
C738 B.n353 VSUBS 0.007479f
C739 B.n354 VSUBS 0.007479f
C740 B.n355 VSUBS 0.007479f
C741 B.n356 VSUBS 0.007479f
C742 B.n357 VSUBS 0.007479f
C743 B.n358 VSUBS 0.007479f
C744 B.n359 VSUBS 0.007479f
C745 B.n360 VSUBS 0.007479f
C746 B.n361 VSUBS 0.007479f
C747 B.n362 VSUBS 0.007479f
C748 B.n363 VSUBS 0.007479f
C749 B.n364 VSUBS 0.007479f
C750 B.n365 VSUBS 0.007479f
C751 B.n366 VSUBS 0.007479f
C752 B.n367 VSUBS 0.007479f
C753 B.n368 VSUBS 0.007479f
C754 B.n369 VSUBS 0.007479f
C755 B.n370 VSUBS 0.007479f
C756 B.n371 VSUBS 0.007479f
C757 B.n372 VSUBS 0.007479f
C758 B.n373 VSUBS 0.007479f
C759 B.n374 VSUBS 0.007479f
C760 B.n375 VSUBS 0.007479f
C761 B.n376 VSUBS 0.007479f
C762 B.n377 VSUBS 0.007479f
C763 B.n378 VSUBS 0.007479f
C764 B.n379 VSUBS 0.007479f
C765 B.n380 VSUBS 0.007479f
C766 B.n381 VSUBS 0.007479f
C767 B.n382 VSUBS 0.007479f
C768 B.n383 VSUBS 0.007479f
C769 B.n384 VSUBS 0.007479f
C770 B.n385 VSUBS 0.007479f
C771 B.n386 VSUBS 0.007479f
C772 B.n387 VSUBS 0.007479f
C773 B.n388 VSUBS 0.017036f
C774 B.n389 VSUBS 0.017036f
C775 B.n390 VSUBS 0.017498f
C776 B.n391 VSUBS 0.007479f
C777 B.n392 VSUBS 0.007479f
C778 B.n393 VSUBS 0.007479f
C779 B.n394 VSUBS 0.007479f
C780 B.n395 VSUBS 0.007479f
C781 B.n396 VSUBS 0.007479f
C782 B.n397 VSUBS 0.007479f
C783 B.n398 VSUBS 0.007479f
C784 B.n399 VSUBS 0.007479f
C785 B.n400 VSUBS 0.007479f
C786 B.n401 VSUBS 0.007479f
C787 B.n402 VSUBS 0.007479f
C788 B.n403 VSUBS 0.007479f
C789 B.n404 VSUBS 0.007479f
C790 B.n405 VSUBS 0.007479f
C791 B.n406 VSUBS 0.007479f
C792 B.n407 VSUBS 0.007479f
C793 B.n408 VSUBS 0.007479f
C794 B.n409 VSUBS 0.007479f
C795 B.n410 VSUBS 0.007479f
C796 B.n411 VSUBS 0.007479f
C797 B.n412 VSUBS 0.007479f
C798 B.n413 VSUBS 0.005169f
C799 B.n414 VSUBS 0.017328f
C800 B.n415 VSUBS 0.006049f
C801 B.n416 VSUBS 0.007479f
C802 B.n417 VSUBS 0.007479f
C803 B.n418 VSUBS 0.007479f
C804 B.n419 VSUBS 0.007479f
C805 B.n420 VSUBS 0.007479f
C806 B.n421 VSUBS 0.007479f
C807 B.n422 VSUBS 0.007479f
C808 B.n423 VSUBS 0.007479f
C809 B.n424 VSUBS 0.007479f
C810 B.n425 VSUBS 0.007479f
C811 B.n426 VSUBS 0.007479f
C812 B.n427 VSUBS 0.006049f
C813 B.n428 VSUBS 0.017328f
C814 B.n429 VSUBS 0.005169f
C815 B.n430 VSUBS 0.007479f
C816 B.n431 VSUBS 0.007479f
C817 B.n432 VSUBS 0.007479f
C818 B.n433 VSUBS 0.007479f
C819 B.n434 VSUBS 0.007479f
C820 B.n435 VSUBS 0.007479f
C821 B.n436 VSUBS 0.007479f
C822 B.n437 VSUBS 0.007479f
C823 B.n438 VSUBS 0.007479f
C824 B.n439 VSUBS 0.007479f
C825 B.n440 VSUBS 0.007479f
C826 B.n441 VSUBS 0.007479f
C827 B.n442 VSUBS 0.007479f
C828 B.n443 VSUBS 0.007479f
C829 B.n444 VSUBS 0.007479f
C830 B.n445 VSUBS 0.007479f
C831 B.n446 VSUBS 0.007479f
C832 B.n447 VSUBS 0.007479f
C833 B.n448 VSUBS 0.007479f
C834 B.n449 VSUBS 0.007479f
C835 B.n450 VSUBS 0.007479f
C836 B.n451 VSUBS 0.007479f
C837 B.n452 VSUBS 0.017498f
C838 B.n453 VSUBS 0.017036f
C839 B.n454 VSUBS 0.017036f
C840 B.n455 VSUBS 0.007479f
C841 B.n456 VSUBS 0.007479f
C842 B.n457 VSUBS 0.007479f
C843 B.n458 VSUBS 0.007479f
C844 B.n459 VSUBS 0.007479f
C845 B.n460 VSUBS 0.007479f
C846 B.n461 VSUBS 0.007479f
C847 B.n462 VSUBS 0.007479f
C848 B.n463 VSUBS 0.007479f
C849 B.n464 VSUBS 0.007479f
C850 B.n465 VSUBS 0.007479f
C851 B.n466 VSUBS 0.007479f
C852 B.n467 VSUBS 0.007479f
C853 B.n468 VSUBS 0.007479f
C854 B.n469 VSUBS 0.007479f
C855 B.n470 VSUBS 0.007479f
C856 B.n471 VSUBS 0.007479f
C857 B.n472 VSUBS 0.007479f
C858 B.n473 VSUBS 0.007479f
C859 B.n474 VSUBS 0.007479f
C860 B.n475 VSUBS 0.007479f
C861 B.n476 VSUBS 0.007479f
C862 B.n477 VSUBS 0.007479f
C863 B.n478 VSUBS 0.007479f
C864 B.n479 VSUBS 0.007479f
C865 B.n480 VSUBS 0.007479f
C866 B.n481 VSUBS 0.007479f
C867 B.n482 VSUBS 0.007479f
C868 B.n483 VSUBS 0.007479f
C869 B.n484 VSUBS 0.007479f
C870 B.n485 VSUBS 0.007479f
C871 B.n486 VSUBS 0.007479f
C872 B.n487 VSUBS 0.007479f
C873 B.n488 VSUBS 0.007479f
C874 B.n489 VSUBS 0.007479f
C875 B.n490 VSUBS 0.007479f
C876 B.n491 VSUBS 0.007479f
C877 B.n492 VSUBS 0.007479f
C878 B.n493 VSUBS 0.007479f
C879 B.n494 VSUBS 0.007479f
C880 B.n495 VSUBS 0.007479f
C881 B.n496 VSUBS 0.007479f
C882 B.n497 VSUBS 0.007479f
C883 B.n498 VSUBS 0.007479f
C884 B.n499 VSUBS 0.007479f
C885 B.n500 VSUBS 0.007479f
C886 B.n501 VSUBS 0.007479f
C887 B.n502 VSUBS 0.007479f
C888 B.n503 VSUBS 0.007479f
C889 B.n504 VSUBS 0.007479f
C890 B.n505 VSUBS 0.007479f
C891 B.n506 VSUBS 0.007479f
C892 B.n507 VSUBS 0.007479f
C893 B.n508 VSUBS 0.007479f
C894 B.n509 VSUBS 0.007479f
C895 B.n510 VSUBS 0.007479f
C896 B.n511 VSUBS 0.007479f
C897 B.n512 VSUBS 0.007479f
C898 B.n513 VSUBS 0.007479f
C899 B.n514 VSUBS 0.007479f
C900 B.n515 VSUBS 0.00976f
C901 B.n516 VSUBS 0.010396f
C902 B.n517 VSUBS 0.020674f
.ends

