* NGSPICE file created from diff_pair_sample_0516.ext - technology: sky130A

.subckt diff_pair_sample_0516 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X1 VDD1.t5 VP.t1 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X2 VTAIL.t13 VP.t2 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0.1617 ps=1.31 w=0.98 l=1.34
X3 VTAIL.t0 VN.t0 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0.1617 ps=1.31 w=0.98 l=1.34
X4 VDD2.t6 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.3822 ps=2.74 w=0.98 l=1.34
X5 VDD1.t1 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.3822 ps=2.74 w=0.98 l=1.34
X6 VTAIL.t11 VP.t4 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0.1617 ps=1.31 w=0.98 l=1.34
X7 VDD1.t3 VP.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.3822 ps=2.74 w=0.98 l=1.34
X8 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X9 VTAIL.t9 VP.t6 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X10 VDD2.t4 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.3822 ps=2.74 w=0.98 l=1.34
X11 VTAIL.t4 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X12 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0 ps=0 w=0.98 l=1.34
X13 VTAIL.t6 VN.t5 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X14 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0.1617 ps=1.31 w=0.98 l=1.34
X15 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0 ps=0 w=0.98 l=1.34
X16 VDD1.t7 VP.t7 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X17 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0 ps=0 w=0.98 l=1.34
X18 VDD2.t0 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=1.34
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0 ps=0 w=0.98 l=1.34
R0 VP.n25 VP.n5 173.228
R1 VP.n44 VP.n43 173.228
R2 VP.n24 VP.n23 173.228
R3 VP.n12 VP.n9 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n15 VP.n8 161.3
R6 VP.n18 VP.n17 161.3
R7 VP.n19 VP.n7 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n22 VP.n6 161.3
R10 VP.n42 VP.n0 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n39 VP.n1 161.3
R13 VP.n38 VP.n37 161.3
R14 VP.n35 VP.n2 161.3
R15 VP.n34 VP.n33 161.3
R16 VP.n32 VP.n3 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n28 VP.n4 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n11 VP.n10 60.9506
R21 VP.n35 VP.n34 56.4773
R22 VP.n15 VP.n14 56.4773
R23 VP.n30 VP.n28 48.2005
R24 VP.n41 VP.n1 48.2005
R25 VP.n21 VP.n7 48.2005
R26 VP.n11 VP.t2 46.6677
R27 VP.n25 VP.n24 36.5763
R28 VP.n28 VP.n27 32.6207
R29 VP.n42 VP.n41 32.6207
R30 VP.n22 VP.n21 32.6207
R31 VP.n12 VP.n11 27.2319
R32 VP.n34 VP.n3 24.3439
R33 VP.n37 VP.n35 24.3439
R34 VP.n17 VP.n15 24.3439
R35 VP.n14 VP.n9 24.3439
R36 VP.n30 VP.n29 20.2056
R37 VP.n36 VP.n1 20.2056
R38 VP.n16 VP.n7 20.2056
R39 VP.n5 VP.t4 17.6259
R40 VP.n29 VP.t7 17.6259
R41 VP.n36 VP.t6 17.6259
R42 VP.n43 VP.t3 17.6259
R43 VP.n23 VP.t5 17.6259
R44 VP.n16 VP.t0 17.6259
R45 VP.n10 VP.t1 17.6259
R46 VP.n27 VP.n5 12.4157
R47 VP.n43 VP.n42 12.4157
R48 VP.n23 VP.n22 12.4157
R49 VP.n29 VP.n3 4.13888
R50 VP.n37 VP.n36 4.13888
R51 VP.n17 VP.n16 4.13888
R52 VP.n10 VP.n9 4.13888
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VDD1 VDD1.n0 240.524
R73 VDD1.n3 VDD1.n2 240.409
R74 VDD1.n3 VDD1.n1 240.409
R75 VDD1.n5 VDD1.n4 239.745
R76 VDD1.n5 VDD1.n3 31.6216
R77 VDD1.n4 VDD1.t4 20.2046
R78 VDD1.n4 VDD1.t3 20.2046
R79 VDD1.n0 VDD1.t6 20.2046
R80 VDD1.n0 VDD1.t5 20.2046
R81 VDD1.n2 VDD1.t0 20.2046
R82 VDD1.n2 VDD1.t1 20.2046
R83 VDD1.n1 VDD1.t2 20.2046
R84 VDD1.n1 VDD1.t7 20.2046
R85 VDD1 VDD1.n5 0.662138
R86 VTAIL.n14 VTAIL.t10 243.27
R87 VTAIL.n11 VTAIL.t13 243.27
R88 VTAIL.n10 VTAIL.t2 243.27
R89 VTAIL.n7 VTAIL.t0 243.27
R90 VTAIL.n15 VTAIL.t5 243.269
R91 VTAIL.n2 VTAIL.t1 243.269
R92 VTAIL.n3 VTAIL.t12 243.269
R93 VTAIL.n6 VTAIL.t11 243.269
R94 VTAIL.n13 VTAIL.n12 223.066
R95 VTAIL.n9 VTAIL.n8 223.066
R96 VTAIL.n1 VTAIL.n0 223.065
R97 VTAIL.n5 VTAIL.n4 223.065
R98 VTAIL.n0 VTAIL.t7 20.2046
R99 VTAIL.n0 VTAIL.t6 20.2046
R100 VTAIL.n4 VTAIL.t8 20.2046
R101 VTAIL.n4 VTAIL.t9 20.2046
R102 VTAIL.n12 VTAIL.t14 20.2046
R103 VTAIL.n12 VTAIL.t15 20.2046
R104 VTAIL.n8 VTAIL.t3 20.2046
R105 VTAIL.n8 VTAIL.t4 20.2046
R106 VTAIL.n15 VTAIL.n14 14.6514
R107 VTAIL.n7 VTAIL.n6 14.6514
R108 VTAIL.n9 VTAIL.n7 1.44016
R109 VTAIL.n10 VTAIL.n9 1.44016
R110 VTAIL.n13 VTAIL.n11 1.44016
R111 VTAIL.n14 VTAIL.n13 1.44016
R112 VTAIL.n6 VTAIL.n5 1.44016
R113 VTAIL.n5 VTAIL.n3 1.44016
R114 VTAIL.n2 VTAIL.n1 1.44016
R115 VTAIL VTAIL.n15 1.38197
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 B.n411 B.n410 585
R120 B.n132 B.n75 585
R121 B.n131 B.n130 585
R122 B.n129 B.n128 585
R123 B.n127 B.n126 585
R124 B.n125 B.n124 585
R125 B.n123 B.n122 585
R126 B.n121 B.n120 585
R127 B.n119 B.n118 585
R128 B.n116 B.n115 585
R129 B.n114 B.n113 585
R130 B.n112 B.n111 585
R131 B.n110 B.n109 585
R132 B.n108 B.n107 585
R133 B.n106 B.n105 585
R134 B.n104 B.n103 585
R135 B.n102 B.n101 585
R136 B.n100 B.n99 585
R137 B.n98 B.n97 585
R138 B.n95 B.n94 585
R139 B.n93 B.n92 585
R140 B.n91 B.n90 585
R141 B.n89 B.n88 585
R142 B.n87 B.n86 585
R143 B.n85 B.n84 585
R144 B.n83 B.n82 585
R145 B.n81 B.n80 585
R146 B.n60 B.n59 585
R147 B.n409 B.n61 585
R148 B.n414 B.n61 585
R149 B.n408 B.n407 585
R150 B.n407 B.n57 585
R151 B.n406 B.n56 585
R152 B.n420 B.n56 585
R153 B.n405 B.n55 585
R154 B.n421 B.n55 585
R155 B.n404 B.n54 585
R156 B.n422 B.n54 585
R157 B.n403 B.n402 585
R158 B.n402 B.n53 585
R159 B.n401 B.n49 585
R160 B.n428 B.n49 585
R161 B.n400 B.n48 585
R162 B.n429 B.n48 585
R163 B.n399 B.n47 585
R164 B.n430 B.n47 585
R165 B.n398 B.n397 585
R166 B.n397 B.n43 585
R167 B.n396 B.n42 585
R168 B.n436 B.n42 585
R169 B.n395 B.n41 585
R170 B.n437 B.n41 585
R171 B.n394 B.n40 585
R172 B.n438 B.n40 585
R173 B.n393 B.n392 585
R174 B.n392 B.n39 585
R175 B.n391 B.n35 585
R176 B.n444 B.n35 585
R177 B.n390 B.n34 585
R178 B.n445 B.n34 585
R179 B.n389 B.n33 585
R180 B.n446 B.n33 585
R181 B.n388 B.n387 585
R182 B.n387 B.n29 585
R183 B.n386 B.n28 585
R184 B.n452 B.n28 585
R185 B.n385 B.n27 585
R186 B.n453 B.n27 585
R187 B.n384 B.n26 585
R188 B.n454 B.n26 585
R189 B.n383 B.n382 585
R190 B.n382 B.n22 585
R191 B.n381 B.n21 585
R192 B.n460 B.n21 585
R193 B.n380 B.n20 585
R194 B.n461 B.n20 585
R195 B.n379 B.n19 585
R196 B.n462 B.n19 585
R197 B.n378 B.n377 585
R198 B.n377 B.n15 585
R199 B.n376 B.n14 585
R200 B.n468 B.n14 585
R201 B.n375 B.n13 585
R202 B.n469 B.n13 585
R203 B.n374 B.n12 585
R204 B.n470 B.n12 585
R205 B.n373 B.n372 585
R206 B.n372 B.n371 585
R207 B.n370 B.n369 585
R208 B.n370 B.n8 585
R209 B.n368 B.n7 585
R210 B.n477 B.n7 585
R211 B.n367 B.n6 585
R212 B.n478 B.n6 585
R213 B.n366 B.n5 585
R214 B.n479 B.n5 585
R215 B.n365 B.n364 585
R216 B.n364 B.n4 585
R217 B.n363 B.n133 585
R218 B.n363 B.n362 585
R219 B.n353 B.n134 585
R220 B.n135 B.n134 585
R221 B.n355 B.n354 585
R222 B.n356 B.n355 585
R223 B.n352 B.n140 585
R224 B.n140 B.n139 585
R225 B.n351 B.n350 585
R226 B.n350 B.n349 585
R227 B.n142 B.n141 585
R228 B.n143 B.n142 585
R229 B.n342 B.n341 585
R230 B.n343 B.n342 585
R231 B.n340 B.n147 585
R232 B.n151 B.n147 585
R233 B.n339 B.n338 585
R234 B.n338 B.n337 585
R235 B.n149 B.n148 585
R236 B.n150 B.n149 585
R237 B.n330 B.n329 585
R238 B.n331 B.n330 585
R239 B.n328 B.n156 585
R240 B.n156 B.n155 585
R241 B.n327 B.n326 585
R242 B.n326 B.n325 585
R243 B.n158 B.n157 585
R244 B.n159 B.n158 585
R245 B.n318 B.n317 585
R246 B.n319 B.n318 585
R247 B.n316 B.n164 585
R248 B.n164 B.n163 585
R249 B.n315 B.n314 585
R250 B.n314 B.n313 585
R251 B.n166 B.n165 585
R252 B.n306 B.n166 585
R253 B.n305 B.n304 585
R254 B.n307 B.n305 585
R255 B.n303 B.n171 585
R256 B.n171 B.n170 585
R257 B.n302 B.n301 585
R258 B.n301 B.n300 585
R259 B.n173 B.n172 585
R260 B.n174 B.n173 585
R261 B.n293 B.n292 585
R262 B.n294 B.n293 585
R263 B.n291 B.n179 585
R264 B.n179 B.n178 585
R265 B.n290 B.n289 585
R266 B.n289 B.n288 585
R267 B.n181 B.n180 585
R268 B.n281 B.n181 585
R269 B.n280 B.n279 585
R270 B.n282 B.n280 585
R271 B.n278 B.n186 585
R272 B.n186 B.n185 585
R273 B.n277 B.n276 585
R274 B.n276 B.n275 585
R275 B.n188 B.n187 585
R276 B.n189 B.n188 585
R277 B.n268 B.n267 585
R278 B.n269 B.n268 585
R279 B.n192 B.n191 585
R280 B.n215 B.n214 585
R281 B.n216 B.n212 585
R282 B.n212 B.n193 585
R283 B.n218 B.n217 585
R284 B.n220 B.n211 585
R285 B.n223 B.n222 585
R286 B.n224 B.n210 585
R287 B.n226 B.n225 585
R288 B.n228 B.n209 585
R289 B.n231 B.n230 585
R290 B.n232 B.n205 585
R291 B.n234 B.n233 585
R292 B.n236 B.n204 585
R293 B.n239 B.n238 585
R294 B.n240 B.n203 585
R295 B.n242 B.n241 585
R296 B.n244 B.n202 585
R297 B.n247 B.n246 585
R298 B.n248 B.n199 585
R299 B.n251 B.n250 585
R300 B.n253 B.n198 585
R301 B.n256 B.n255 585
R302 B.n257 B.n197 585
R303 B.n259 B.n258 585
R304 B.n261 B.n196 585
R305 B.n262 B.n195 585
R306 B.n265 B.n264 585
R307 B.n266 B.n194 585
R308 B.n194 B.n193 585
R309 B.n271 B.n270 585
R310 B.n270 B.n269 585
R311 B.n272 B.n190 585
R312 B.n190 B.n189 585
R313 B.n274 B.n273 585
R314 B.n275 B.n274 585
R315 B.n184 B.n183 585
R316 B.n185 B.n184 585
R317 B.n284 B.n283 585
R318 B.n283 B.n282 585
R319 B.n285 B.n182 585
R320 B.n281 B.n182 585
R321 B.n287 B.n286 585
R322 B.n288 B.n287 585
R323 B.n177 B.n176 585
R324 B.n178 B.n177 585
R325 B.n296 B.n295 585
R326 B.n295 B.n294 585
R327 B.n297 B.n175 585
R328 B.n175 B.n174 585
R329 B.n299 B.n298 585
R330 B.n300 B.n299 585
R331 B.n169 B.n168 585
R332 B.n170 B.n169 585
R333 B.n309 B.n308 585
R334 B.n308 B.n307 585
R335 B.n310 B.n167 585
R336 B.n306 B.n167 585
R337 B.n312 B.n311 585
R338 B.n313 B.n312 585
R339 B.n162 B.n161 585
R340 B.n163 B.n162 585
R341 B.n321 B.n320 585
R342 B.n320 B.n319 585
R343 B.n322 B.n160 585
R344 B.n160 B.n159 585
R345 B.n324 B.n323 585
R346 B.n325 B.n324 585
R347 B.n154 B.n153 585
R348 B.n155 B.n154 585
R349 B.n333 B.n332 585
R350 B.n332 B.n331 585
R351 B.n334 B.n152 585
R352 B.n152 B.n150 585
R353 B.n336 B.n335 585
R354 B.n337 B.n336 585
R355 B.n146 B.n145 585
R356 B.n151 B.n146 585
R357 B.n345 B.n344 585
R358 B.n344 B.n343 585
R359 B.n346 B.n144 585
R360 B.n144 B.n143 585
R361 B.n348 B.n347 585
R362 B.n349 B.n348 585
R363 B.n138 B.n137 585
R364 B.n139 B.n138 585
R365 B.n358 B.n357 585
R366 B.n357 B.n356 585
R367 B.n359 B.n136 585
R368 B.n136 B.n135 585
R369 B.n361 B.n360 585
R370 B.n362 B.n361 585
R371 B.n3 B.n0 585
R372 B.n4 B.n3 585
R373 B.n476 B.n1 585
R374 B.n477 B.n476 585
R375 B.n475 B.n474 585
R376 B.n475 B.n8 585
R377 B.n473 B.n9 585
R378 B.n371 B.n9 585
R379 B.n472 B.n471 585
R380 B.n471 B.n470 585
R381 B.n11 B.n10 585
R382 B.n469 B.n11 585
R383 B.n467 B.n466 585
R384 B.n468 B.n467 585
R385 B.n465 B.n16 585
R386 B.n16 B.n15 585
R387 B.n464 B.n463 585
R388 B.n463 B.n462 585
R389 B.n18 B.n17 585
R390 B.n461 B.n18 585
R391 B.n459 B.n458 585
R392 B.n460 B.n459 585
R393 B.n457 B.n23 585
R394 B.n23 B.n22 585
R395 B.n456 B.n455 585
R396 B.n455 B.n454 585
R397 B.n25 B.n24 585
R398 B.n453 B.n25 585
R399 B.n451 B.n450 585
R400 B.n452 B.n451 585
R401 B.n449 B.n30 585
R402 B.n30 B.n29 585
R403 B.n448 B.n447 585
R404 B.n447 B.n446 585
R405 B.n32 B.n31 585
R406 B.n445 B.n32 585
R407 B.n443 B.n442 585
R408 B.n444 B.n443 585
R409 B.n441 B.n36 585
R410 B.n39 B.n36 585
R411 B.n440 B.n439 585
R412 B.n439 B.n438 585
R413 B.n38 B.n37 585
R414 B.n437 B.n38 585
R415 B.n435 B.n434 585
R416 B.n436 B.n435 585
R417 B.n433 B.n44 585
R418 B.n44 B.n43 585
R419 B.n432 B.n431 585
R420 B.n431 B.n430 585
R421 B.n46 B.n45 585
R422 B.n429 B.n46 585
R423 B.n427 B.n426 585
R424 B.n428 B.n427 585
R425 B.n425 B.n50 585
R426 B.n53 B.n50 585
R427 B.n424 B.n423 585
R428 B.n423 B.n422 585
R429 B.n52 B.n51 585
R430 B.n421 B.n52 585
R431 B.n419 B.n418 585
R432 B.n420 B.n419 585
R433 B.n417 B.n58 585
R434 B.n58 B.n57 585
R435 B.n416 B.n415 585
R436 B.n415 B.n414 585
R437 B.n480 B.n479 585
R438 B.n478 B.n2 585
R439 B.n415 B.n60 526.135
R440 B.n411 B.n61 526.135
R441 B.n268 B.n194 526.135
R442 B.n270 B.n192 526.135
R443 B.n78 B.t17 266.296
R444 B.n76 B.t14 266.296
R445 B.n200 B.t11 266.296
R446 B.n206 B.t21 266.296
R447 B.n413 B.n412 256.663
R448 B.n413 B.n74 256.663
R449 B.n413 B.n73 256.663
R450 B.n413 B.n72 256.663
R451 B.n413 B.n71 256.663
R452 B.n413 B.n70 256.663
R453 B.n413 B.n69 256.663
R454 B.n413 B.n68 256.663
R455 B.n413 B.n67 256.663
R456 B.n413 B.n66 256.663
R457 B.n413 B.n65 256.663
R458 B.n413 B.n64 256.663
R459 B.n413 B.n63 256.663
R460 B.n413 B.n62 256.663
R461 B.n213 B.n193 256.663
R462 B.n219 B.n193 256.663
R463 B.n221 B.n193 256.663
R464 B.n227 B.n193 256.663
R465 B.n229 B.n193 256.663
R466 B.n235 B.n193 256.663
R467 B.n237 B.n193 256.663
R468 B.n243 B.n193 256.663
R469 B.n245 B.n193 256.663
R470 B.n252 B.n193 256.663
R471 B.n254 B.n193 256.663
R472 B.n260 B.n193 256.663
R473 B.n263 B.n193 256.663
R474 B.n482 B.n481 256.663
R475 B.n269 B.n193 237.411
R476 B.n414 B.n413 237.411
R477 B.n79 B.t18 233.907
R478 B.n77 B.t15 233.907
R479 B.n201 B.t10 233.907
R480 B.n207 B.t20 233.907
R481 B.n78 B.t16 222.416
R482 B.n76 B.t12 222.416
R483 B.n200 B.t8 222.416
R484 B.n206 B.t19 222.416
R485 B.n82 B.n81 163.367
R486 B.n86 B.n85 163.367
R487 B.n90 B.n89 163.367
R488 B.n94 B.n93 163.367
R489 B.n99 B.n98 163.367
R490 B.n103 B.n102 163.367
R491 B.n107 B.n106 163.367
R492 B.n111 B.n110 163.367
R493 B.n115 B.n114 163.367
R494 B.n120 B.n119 163.367
R495 B.n124 B.n123 163.367
R496 B.n128 B.n127 163.367
R497 B.n130 B.n75 163.367
R498 B.n268 B.n188 163.367
R499 B.n276 B.n188 163.367
R500 B.n276 B.n186 163.367
R501 B.n280 B.n186 163.367
R502 B.n280 B.n181 163.367
R503 B.n289 B.n181 163.367
R504 B.n289 B.n179 163.367
R505 B.n293 B.n179 163.367
R506 B.n293 B.n173 163.367
R507 B.n301 B.n173 163.367
R508 B.n301 B.n171 163.367
R509 B.n305 B.n171 163.367
R510 B.n305 B.n166 163.367
R511 B.n314 B.n166 163.367
R512 B.n314 B.n164 163.367
R513 B.n318 B.n164 163.367
R514 B.n318 B.n158 163.367
R515 B.n326 B.n158 163.367
R516 B.n326 B.n156 163.367
R517 B.n330 B.n156 163.367
R518 B.n330 B.n149 163.367
R519 B.n338 B.n149 163.367
R520 B.n338 B.n147 163.367
R521 B.n342 B.n147 163.367
R522 B.n342 B.n142 163.367
R523 B.n350 B.n142 163.367
R524 B.n350 B.n140 163.367
R525 B.n355 B.n140 163.367
R526 B.n355 B.n134 163.367
R527 B.n363 B.n134 163.367
R528 B.n364 B.n363 163.367
R529 B.n364 B.n5 163.367
R530 B.n6 B.n5 163.367
R531 B.n7 B.n6 163.367
R532 B.n370 B.n7 163.367
R533 B.n372 B.n370 163.367
R534 B.n372 B.n12 163.367
R535 B.n13 B.n12 163.367
R536 B.n14 B.n13 163.367
R537 B.n377 B.n14 163.367
R538 B.n377 B.n19 163.367
R539 B.n20 B.n19 163.367
R540 B.n21 B.n20 163.367
R541 B.n382 B.n21 163.367
R542 B.n382 B.n26 163.367
R543 B.n27 B.n26 163.367
R544 B.n28 B.n27 163.367
R545 B.n387 B.n28 163.367
R546 B.n387 B.n33 163.367
R547 B.n34 B.n33 163.367
R548 B.n35 B.n34 163.367
R549 B.n392 B.n35 163.367
R550 B.n392 B.n40 163.367
R551 B.n41 B.n40 163.367
R552 B.n42 B.n41 163.367
R553 B.n397 B.n42 163.367
R554 B.n397 B.n47 163.367
R555 B.n48 B.n47 163.367
R556 B.n49 B.n48 163.367
R557 B.n402 B.n49 163.367
R558 B.n402 B.n54 163.367
R559 B.n55 B.n54 163.367
R560 B.n56 B.n55 163.367
R561 B.n407 B.n56 163.367
R562 B.n407 B.n61 163.367
R563 B.n214 B.n212 163.367
R564 B.n218 B.n212 163.367
R565 B.n222 B.n220 163.367
R566 B.n226 B.n210 163.367
R567 B.n230 B.n228 163.367
R568 B.n234 B.n205 163.367
R569 B.n238 B.n236 163.367
R570 B.n242 B.n203 163.367
R571 B.n246 B.n244 163.367
R572 B.n251 B.n199 163.367
R573 B.n255 B.n253 163.367
R574 B.n259 B.n197 163.367
R575 B.n262 B.n261 163.367
R576 B.n264 B.n194 163.367
R577 B.n270 B.n190 163.367
R578 B.n274 B.n190 163.367
R579 B.n274 B.n184 163.367
R580 B.n283 B.n184 163.367
R581 B.n283 B.n182 163.367
R582 B.n287 B.n182 163.367
R583 B.n287 B.n177 163.367
R584 B.n295 B.n177 163.367
R585 B.n295 B.n175 163.367
R586 B.n299 B.n175 163.367
R587 B.n299 B.n169 163.367
R588 B.n308 B.n169 163.367
R589 B.n308 B.n167 163.367
R590 B.n312 B.n167 163.367
R591 B.n312 B.n162 163.367
R592 B.n320 B.n162 163.367
R593 B.n320 B.n160 163.367
R594 B.n324 B.n160 163.367
R595 B.n324 B.n154 163.367
R596 B.n332 B.n154 163.367
R597 B.n332 B.n152 163.367
R598 B.n336 B.n152 163.367
R599 B.n336 B.n146 163.367
R600 B.n344 B.n146 163.367
R601 B.n344 B.n144 163.367
R602 B.n348 B.n144 163.367
R603 B.n348 B.n138 163.367
R604 B.n357 B.n138 163.367
R605 B.n357 B.n136 163.367
R606 B.n361 B.n136 163.367
R607 B.n361 B.n3 163.367
R608 B.n480 B.n3 163.367
R609 B.n476 B.n2 163.367
R610 B.n476 B.n475 163.367
R611 B.n475 B.n9 163.367
R612 B.n471 B.n9 163.367
R613 B.n471 B.n11 163.367
R614 B.n467 B.n11 163.367
R615 B.n467 B.n16 163.367
R616 B.n463 B.n16 163.367
R617 B.n463 B.n18 163.367
R618 B.n459 B.n18 163.367
R619 B.n459 B.n23 163.367
R620 B.n455 B.n23 163.367
R621 B.n455 B.n25 163.367
R622 B.n451 B.n25 163.367
R623 B.n451 B.n30 163.367
R624 B.n447 B.n30 163.367
R625 B.n447 B.n32 163.367
R626 B.n443 B.n32 163.367
R627 B.n443 B.n36 163.367
R628 B.n439 B.n36 163.367
R629 B.n439 B.n38 163.367
R630 B.n435 B.n38 163.367
R631 B.n435 B.n44 163.367
R632 B.n431 B.n44 163.367
R633 B.n431 B.n46 163.367
R634 B.n427 B.n46 163.367
R635 B.n427 B.n50 163.367
R636 B.n423 B.n50 163.367
R637 B.n423 B.n52 163.367
R638 B.n419 B.n52 163.367
R639 B.n419 B.n58 163.367
R640 B.n415 B.n58 163.367
R641 B.n269 B.n189 119.585
R642 B.n275 B.n189 119.585
R643 B.n275 B.n185 119.585
R644 B.n282 B.n185 119.585
R645 B.n282 B.n281 119.585
R646 B.n288 B.n178 119.585
R647 B.n294 B.n178 119.585
R648 B.n294 B.n174 119.585
R649 B.n300 B.n174 119.585
R650 B.n300 B.n170 119.585
R651 B.n307 B.n170 119.585
R652 B.n307 B.n306 119.585
R653 B.n313 B.n163 119.585
R654 B.n319 B.n163 119.585
R655 B.n319 B.n159 119.585
R656 B.n325 B.n159 119.585
R657 B.n331 B.n155 119.585
R658 B.n331 B.n150 119.585
R659 B.n337 B.n150 119.585
R660 B.n337 B.n151 119.585
R661 B.n343 B.n143 119.585
R662 B.n349 B.n143 119.585
R663 B.n349 B.n139 119.585
R664 B.n356 B.n139 119.585
R665 B.n362 B.n135 119.585
R666 B.n362 B.n4 119.585
R667 B.n479 B.n4 119.585
R668 B.n479 B.n478 119.585
R669 B.n478 B.n477 119.585
R670 B.n477 B.n8 119.585
R671 B.n371 B.n8 119.585
R672 B.n470 B.n469 119.585
R673 B.n469 B.n468 119.585
R674 B.n468 B.n15 119.585
R675 B.n462 B.n15 119.585
R676 B.n461 B.n460 119.585
R677 B.n460 B.n22 119.585
R678 B.n454 B.n22 119.585
R679 B.n454 B.n453 119.585
R680 B.n452 B.n29 119.585
R681 B.n446 B.n29 119.585
R682 B.n446 B.n445 119.585
R683 B.n445 B.n444 119.585
R684 B.n438 B.n39 119.585
R685 B.n438 B.n437 119.585
R686 B.n437 B.n436 119.585
R687 B.n436 B.n43 119.585
R688 B.n430 B.n43 119.585
R689 B.n430 B.n429 119.585
R690 B.n429 B.n428 119.585
R691 B.n422 B.n53 119.585
R692 B.n422 B.n421 119.585
R693 B.n421 B.n420 119.585
R694 B.n420 B.n57 119.585
R695 B.n414 B.n57 119.585
R696 B.n306 B.t0 84.413
R697 B.n39 B.t5 84.413
R698 B.n325 B.t3 73.8614
R699 B.t6 B.n452 73.8614
R700 B.n62 B.n60 71.676
R701 B.n82 B.n63 71.676
R702 B.n86 B.n64 71.676
R703 B.n90 B.n65 71.676
R704 B.n94 B.n66 71.676
R705 B.n99 B.n67 71.676
R706 B.n103 B.n68 71.676
R707 B.n107 B.n69 71.676
R708 B.n111 B.n70 71.676
R709 B.n115 B.n71 71.676
R710 B.n120 B.n72 71.676
R711 B.n124 B.n73 71.676
R712 B.n128 B.n74 71.676
R713 B.n412 B.n75 71.676
R714 B.n412 B.n411 71.676
R715 B.n130 B.n74 71.676
R716 B.n127 B.n73 71.676
R717 B.n123 B.n72 71.676
R718 B.n119 B.n71 71.676
R719 B.n114 B.n70 71.676
R720 B.n110 B.n69 71.676
R721 B.n106 B.n68 71.676
R722 B.n102 B.n67 71.676
R723 B.n98 B.n66 71.676
R724 B.n93 B.n65 71.676
R725 B.n89 B.n64 71.676
R726 B.n85 B.n63 71.676
R727 B.n81 B.n62 71.676
R728 B.n213 B.n192 71.676
R729 B.n219 B.n218 71.676
R730 B.n222 B.n221 71.676
R731 B.n227 B.n226 71.676
R732 B.n230 B.n229 71.676
R733 B.n235 B.n234 71.676
R734 B.n238 B.n237 71.676
R735 B.n243 B.n242 71.676
R736 B.n246 B.n245 71.676
R737 B.n252 B.n251 71.676
R738 B.n255 B.n254 71.676
R739 B.n260 B.n259 71.676
R740 B.n263 B.n262 71.676
R741 B.n214 B.n213 71.676
R742 B.n220 B.n219 71.676
R743 B.n221 B.n210 71.676
R744 B.n228 B.n227 71.676
R745 B.n229 B.n205 71.676
R746 B.n236 B.n235 71.676
R747 B.n237 B.n203 71.676
R748 B.n244 B.n243 71.676
R749 B.n245 B.n199 71.676
R750 B.n253 B.n252 71.676
R751 B.n254 B.n197 71.676
R752 B.n261 B.n260 71.676
R753 B.n264 B.n263 71.676
R754 B.n481 B.n480 71.676
R755 B.n481 B.n2 71.676
R756 B.n281 B.t9 70.3442
R757 B.n53 B.t13 70.3442
R758 B.t2 B.n135 66.827
R759 B.n371 B.t1 66.827
R760 B.n151 B.t4 63.3099
R761 B.t7 B.n461 63.3099
R762 B.n96 B.n79 59.5399
R763 B.n117 B.n77 59.5399
R764 B.n249 B.n201 59.5399
R765 B.n208 B.n207 59.5399
R766 B.n343 B.t4 56.2755
R767 B.n462 B.t7 56.2755
R768 B.n356 B.t2 52.7583
R769 B.n470 B.t1 52.7583
R770 B.n288 B.t9 49.2411
R771 B.n428 B.t13 49.2411
R772 B.t3 B.n155 45.7239
R773 B.n453 B.t6 45.7239
R774 B.n313 B.t0 35.1724
R775 B.n444 B.t5 35.1724
R776 B.n271 B.n191 34.1859
R777 B.n267 B.n266 34.1859
R778 B.n410 B.n409 34.1859
R779 B.n416 B.n59 34.1859
R780 B.n79 B.n78 32.3884
R781 B.n77 B.n76 32.3884
R782 B.n201 B.n200 32.3884
R783 B.n207 B.n206 32.3884
R784 B B.n482 18.0485
R785 B.n272 B.n271 10.6151
R786 B.n273 B.n272 10.6151
R787 B.n273 B.n183 10.6151
R788 B.n284 B.n183 10.6151
R789 B.n285 B.n284 10.6151
R790 B.n286 B.n285 10.6151
R791 B.n286 B.n176 10.6151
R792 B.n296 B.n176 10.6151
R793 B.n297 B.n296 10.6151
R794 B.n298 B.n297 10.6151
R795 B.n298 B.n168 10.6151
R796 B.n309 B.n168 10.6151
R797 B.n310 B.n309 10.6151
R798 B.n311 B.n310 10.6151
R799 B.n311 B.n161 10.6151
R800 B.n321 B.n161 10.6151
R801 B.n322 B.n321 10.6151
R802 B.n323 B.n322 10.6151
R803 B.n323 B.n153 10.6151
R804 B.n333 B.n153 10.6151
R805 B.n334 B.n333 10.6151
R806 B.n335 B.n334 10.6151
R807 B.n335 B.n145 10.6151
R808 B.n345 B.n145 10.6151
R809 B.n346 B.n345 10.6151
R810 B.n347 B.n346 10.6151
R811 B.n347 B.n137 10.6151
R812 B.n358 B.n137 10.6151
R813 B.n359 B.n358 10.6151
R814 B.n360 B.n359 10.6151
R815 B.n360 B.n0 10.6151
R816 B.n215 B.n191 10.6151
R817 B.n216 B.n215 10.6151
R818 B.n217 B.n216 10.6151
R819 B.n217 B.n211 10.6151
R820 B.n223 B.n211 10.6151
R821 B.n224 B.n223 10.6151
R822 B.n225 B.n224 10.6151
R823 B.n225 B.n209 10.6151
R824 B.n232 B.n231 10.6151
R825 B.n233 B.n232 10.6151
R826 B.n233 B.n204 10.6151
R827 B.n239 B.n204 10.6151
R828 B.n240 B.n239 10.6151
R829 B.n241 B.n240 10.6151
R830 B.n241 B.n202 10.6151
R831 B.n247 B.n202 10.6151
R832 B.n248 B.n247 10.6151
R833 B.n250 B.n198 10.6151
R834 B.n256 B.n198 10.6151
R835 B.n257 B.n256 10.6151
R836 B.n258 B.n257 10.6151
R837 B.n258 B.n196 10.6151
R838 B.n196 B.n195 10.6151
R839 B.n265 B.n195 10.6151
R840 B.n266 B.n265 10.6151
R841 B.n267 B.n187 10.6151
R842 B.n277 B.n187 10.6151
R843 B.n278 B.n277 10.6151
R844 B.n279 B.n278 10.6151
R845 B.n279 B.n180 10.6151
R846 B.n290 B.n180 10.6151
R847 B.n291 B.n290 10.6151
R848 B.n292 B.n291 10.6151
R849 B.n292 B.n172 10.6151
R850 B.n302 B.n172 10.6151
R851 B.n303 B.n302 10.6151
R852 B.n304 B.n303 10.6151
R853 B.n304 B.n165 10.6151
R854 B.n315 B.n165 10.6151
R855 B.n316 B.n315 10.6151
R856 B.n317 B.n316 10.6151
R857 B.n317 B.n157 10.6151
R858 B.n327 B.n157 10.6151
R859 B.n328 B.n327 10.6151
R860 B.n329 B.n328 10.6151
R861 B.n329 B.n148 10.6151
R862 B.n339 B.n148 10.6151
R863 B.n340 B.n339 10.6151
R864 B.n341 B.n340 10.6151
R865 B.n341 B.n141 10.6151
R866 B.n351 B.n141 10.6151
R867 B.n352 B.n351 10.6151
R868 B.n354 B.n352 10.6151
R869 B.n354 B.n353 10.6151
R870 B.n353 B.n133 10.6151
R871 B.n365 B.n133 10.6151
R872 B.n366 B.n365 10.6151
R873 B.n367 B.n366 10.6151
R874 B.n368 B.n367 10.6151
R875 B.n369 B.n368 10.6151
R876 B.n373 B.n369 10.6151
R877 B.n374 B.n373 10.6151
R878 B.n375 B.n374 10.6151
R879 B.n376 B.n375 10.6151
R880 B.n378 B.n376 10.6151
R881 B.n379 B.n378 10.6151
R882 B.n380 B.n379 10.6151
R883 B.n381 B.n380 10.6151
R884 B.n383 B.n381 10.6151
R885 B.n384 B.n383 10.6151
R886 B.n385 B.n384 10.6151
R887 B.n386 B.n385 10.6151
R888 B.n388 B.n386 10.6151
R889 B.n389 B.n388 10.6151
R890 B.n390 B.n389 10.6151
R891 B.n391 B.n390 10.6151
R892 B.n393 B.n391 10.6151
R893 B.n394 B.n393 10.6151
R894 B.n395 B.n394 10.6151
R895 B.n396 B.n395 10.6151
R896 B.n398 B.n396 10.6151
R897 B.n399 B.n398 10.6151
R898 B.n400 B.n399 10.6151
R899 B.n401 B.n400 10.6151
R900 B.n403 B.n401 10.6151
R901 B.n404 B.n403 10.6151
R902 B.n405 B.n404 10.6151
R903 B.n406 B.n405 10.6151
R904 B.n408 B.n406 10.6151
R905 B.n409 B.n408 10.6151
R906 B.n474 B.n1 10.6151
R907 B.n474 B.n473 10.6151
R908 B.n473 B.n472 10.6151
R909 B.n472 B.n10 10.6151
R910 B.n466 B.n10 10.6151
R911 B.n466 B.n465 10.6151
R912 B.n465 B.n464 10.6151
R913 B.n464 B.n17 10.6151
R914 B.n458 B.n17 10.6151
R915 B.n458 B.n457 10.6151
R916 B.n457 B.n456 10.6151
R917 B.n456 B.n24 10.6151
R918 B.n450 B.n24 10.6151
R919 B.n450 B.n449 10.6151
R920 B.n449 B.n448 10.6151
R921 B.n448 B.n31 10.6151
R922 B.n442 B.n31 10.6151
R923 B.n442 B.n441 10.6151
R924 B.n441 B.n440 10.6151
R925 B.n440 B.n37 10.6151
R926 B.n434 B.n37 10.6151
R927 B.n434 B.n433 10.6151
R928 B.n433 B.n432 10.6151
R929 B.n432 B.n45 10.6151
R930 B.n426 B.n45 10.6151
R931 B.n426 B.n425 10.6151
R932 B.n425 B.n424 10.6151
R933 B.n424 B.n51 10.6151
R934 B.n418 B.n51 10.6151
R935 B.n418 B.n417 10.6151
R936 B.n417 B.n416 10.6151
R937 B.n80 B.n59 10.6151
R938 B.n83 B.n80 10.6151
R939 B.n84 B.n83 10.6151
R940 B.n87 B.n84 10.6151
R941 B.n88 B.n87 10.6151
R942 B.n91 B.n88 10.6151
R943 B.n92 B.n91 10.6151
R944 B.n95 B.n92 10.6151
R945 B.n100 B.n97 10.6151
R946 B.n101 B.n100 10.6151
R947 B.n104 B.n101 10.6151
R948 B.n105 B.n104 10.6151
R949 B.n108 B.n105 10.6151
R950 B.n109 B.n108 10.6151
R951 B.n112 B.n109 10.6151
R952 B.n113 B.n112 10.6151
R953 B.n116 B.n113 10.6151
R954 B.n121 B.n118 10.6151
R955 B.n122 B.n121 10.6151
R956 B.n125 B.n122 10.6151
R957 B.n126 B.n125 10.6151
R958 B.n129 B.n126 10.6151
R959 B.n131 B.n129 10.6151
R960 B.n132 B.n131 10.6151
R961 B.n410 B.n132 10.6151
R962 B.n209 B.n208 9.36635
R963 B.n250 B.n249 9.36635
R964 B.n96 B.n95 9.36635
R965 B.n118 B.n117 9.36635
R966 B.n482 B.n0 8.11757
R967 B.n482 B.n1 8.11757
R968 B.n231 B.n208 1.24928
R969 B.n249 B.n248 1.24928
R970 B.n97 B.n96 1.24928
R971 B.n117 B.n116 1.24928
R972 VN.n18 VN.n17 173.228
R973 VN.n37 VN.n36 173.228
R974 VN.n35 VN.n19 161.3
R975 VN.n34 VN.n33 161.3
R976 VN.n32 VN.n20 161.3
R977 VN.n31 VN.n30 161.3
R978 VN.n29 VN.n21 161.3
R979 VN.n28 VN.n27 161.3
R980 VN.n26 VN.n23 161.3
R981 VN.n16 VN.n0 161.3
R982 VN.n15 VN.n14 161.3
R983 VN.n13 VN.n1 161.3
R984 VN.n12 VN.n11 161.3
R985 VN.n9 VN.n2 161.3
R986 VN.n8 VN.n7 161.3
R987 VN.n6 VN.n3 161.3
R988 VN.n5 VN.n4 60.9506
R989 VN.n25 VN.n24 60.9506
R990 VN.n9 VN.n8 56.4773
R991 VN.n29 VN.n28 56.4773
R992 VN.n15 VN.n1 48.2005
R993 VN.n34 VN.n20 48.2005
R994 VN.n5 VN.t6 46.6677
R995 VN.n25 VN.t3 46.6677
R996 VN VN.n37 36.9569
R997 VN.n16 VN.n15 32.6207
R998 VN.n35 VN.n34 32.6207
R999 VN.n26 VN.n25 27.2319
R1000 VN.n6 VN.n5 27.2319
R1001 VN.n8 VN.n3 24.3439
R1002 VN.n11 VN.n9 24.3439
R1003 VN.n28 VN.n23 24.3439
R1004 VN.n30 VN.n29 24.3439
R1005 VN.n10 VN.n1 20.2056
R1006 VN.n22 VN.n20 20.2056
R1007 VN.n4 VN.t2 17.6259
R1008 VN.n10 VN.t5 17.6259
R1009 VN.n17 VN.t1 17.6259
R1010 VN.n24 VN.t4 17.6259
R1011 VN.n22 VN.t7 17.6259
R1012 VN.n36 VN.t0 17.6259
R1013 VN.n17 VN.n16 12.4157
R1014 VN.n36 VN.n35 12.4157
R1015 VN.n4 VN.n3 4.13888
R1016 VN.n11 VN.n10 4.13888
R1017 VN.n24 VN.n23 4.13888
R1018 VN.n30 VN.n22 4.13888
R1019 VN.n37 VN.n19 0.189894
R1020 VN.n33 VN.n19 0.189894
R1021 VN.n33 VN.n32 0.189894
R1022 VN.n32 VN.n31 0.189894
R1023 VN.n31 VN.n21 0.189894
R1024 VN.n27 VN.n21 0.189894
R1025 VN.n27 VN.n26 0.189894
R1026 VN.n7 VN.n6 0.189894
R1027 VN.n7 VN.n2 0.189894
R1028 VN.n12 VN.n2 0.189894
R1029 VN.n13 VN.n12 0.189894
R1030 VN.n14 VN.n13 0.189894
R1031 VN.n14 VN.n0 0.189894
R1032 VN.n18 VN.n0 0.189894
R1033 VN VN.n18 0.0516364
R1034 VDD2.n2 VDD2.n1 240.409
R1035 VDD2.n2 VDD2.n0 240.409
R1036 VDD2 VDD2.n5 240.406
R1037 VDD2.n4 VDD2.n3 239.745
R1038 VDD2.n4 VDD2.n2 31.0386
R1039 VDD2.n5 VDD2.t3 20.2046
R1040 VDD2.n5 VDD2.t4 20.2046
R1041 VDD2.n3 VDD2.t7 20.2046
R1042 VDD2.n3 VDD2.t0 20.2046
R1043 VDD2.n1 VDD2.t2 20.2046
R1044 VDD2.n1 VDD2.t6 20.2046
R1045 VDD2.n0 VDD2.t1 20.2046
R1046 VDD2.n0 VDD2.t5 20.2046
R1047 VDD2 VDD2.n4 0.778517
C0 VDD2 VDD1 1.14586f
C1 VTAIL VP 1.66307f
C2 VTAIL VDD1 3.23752f
C3 VTAIL VDD2 3.28349f
C4 VN VP 4.09475f
C5 VN VDD1 0.156004f
C6 VN VDD2 0.985075f
C7 VP VDD1 1.22022f
C8 VDD2 VP 0.393592f
C9 VN VTAIL 1.64896f
C10 VDD2 B 3.088926f
C11 VDD1 B 3.368651f
C12 VTAIL B 2.729537f
C13 VN B 9.163063f
C14 VP B 8.17011f
C15 VDD2.t1 B 0.014654f
C16 VDD2.t5 B 0.014654f
C17 VDD2.n0 B 0.057658f
C18 VDD2.t2 B 0.014654f
C19 VDD2.t6 B 0.014654f
C20 VDD2.n1 B 0.057658f
C21 VDD2.n2 B 1.38657f
C22 VDD2.t7 B 0.014654f
C23 VDD2.t0 B 0.014654f
C24 VDD2.n3 B 0.056919f
C25 VDD2.n4 B 1.21286f
C26 VDD2.t3 B 0.014654f
C27 VDD2.t4 B 0.014654f
C28 VDD2.n5 B 0.057653f
C29 VN.n0 B 0.025388f
C30 VN.t1 B 0.061653f
C31 VN.n1 B 0.043795f
C32 VN.n2 B 0.025388f
C33 VN.n3 B 0.028066f
C34 VN.t6 B 0.147569f
C35 VN.t2 B 0.061653f
C36 VN.n4 B 0.089936f
C37 VN.n5 B 0.089622f
C38 VN.n6 B 0.134712f
C39 VN.n7 B 0.025388f
C40 VN.n8 B 0.037223f
C41 VN.n9 B 0.037223f
C42 VN.t5 B 0.061653f
C43 VN.n10 B 0.054624f
C44 VN.n11 B 0.028066f
C45 VN.n12 B 0.025388f
C46 VN.n13 B 0.025388f
C47 VN.n14 B 0.025388f
C48 VN.n15 B 0.022728f
C49 VN.n16 B 0.039981f
C50 VN.n17 B 0.103057f
C51 VN.n18 B 0.023257f
C52 VN.n19 B 0.025388f
C53 VN.t0 B 0.061653f
C54 VN.n20 B 0.043795f
C55 VN.n21 B 0.025388f
C56 VN.t7 B 0.061653f
C57 VN.n22 B 0.054624f
C58 VN.n23 B 0.028066f
C59 VN.t3 B 0.147569f
C60 VN.t4 B 0.061653f
C61 VN.n24 B 0.089936f
C62 VN.n25 B 0.089622f
C63 VN.n26 B 0.134712f
C64 VN.n27 B 0.025388f
C65 VN.n28 B 0.037223f
C66 VN.n29 B 0.037223f
C67 VN.n30 B 0.028066f
C68 VN.n31 B 0.025388f
C69 VN.n32 B 0.025388f
C70 VN.n33 B 0.025388f
C71 VN.n34 B 0.022728f
C72 VN.n35 B 0.039981f
C73 VN.n36 B 0.103057f
C74 VN.n37 B 0.842642f
C75 VTAIL.t7 B 0.01737f
C76 VTAIL.t6 B 0.01737f
C77 VTAIL.n0 B 0.056206f
C78 VTAIL.n1 B 0.24391f
C79 VTAIL.t1 B 0.096419f
C80 VTAIL.n2 B 0.28082f
C81 VTAIL.t12 B 0.096419f
C82 VTAIL.n3 B 0.28082f
C83 VTAIL.t8 B 0.01737f
C84 VTAIL.t9 B 0.01737f
C85 VTAIL.n4 B 0.056206f
C86 VTAIL.n5 B 0.343751f
C87 VTAIL.t11 B 0.096419f
C88 VTAIL.n6 B 0.716645f
C89 VTAIL.t0 B 0.096419f
C90 VTAIL.n7 B 0.716645f
C91 VTAIL.t3 B 0.01737f
C92 VTAIL.t4 B 0.01737f
C93 VTAIL.n8 B 0.056206f
C94 VTAIL.n9 B 0.343751f
C95 VTAIL.t2 B 0.096419f
C96 VTAIL.n10 B 0.280819f
C97 VTAIL.t13 B 0.096419f
C98 VTAIL.n11 B 0.280819f
C99 VTAIL.t14 B 0.01737f
C100 VTAIL.t15 B 0.01737f
C101 VTAIL.n12 B 0.056206f
C102 VTAIL.n13 B 0.343751f
C103 VTAIL.t10 B 0.096419f
C104 VTAIL.n14 B 0.716645f
C105 VTAIL.t5 B 0.096419f
C106 VTAIL.n15 B 0.71244f
C107 VDD1.t6 B 0.013915f
C108 VDD1.t5 B 0.013915f
C109 VDD1.n0 B 0.05489f
C110 VDD1.t2 B 0.013915f
C111 VDD1.t7 B 0.013915f
C112 VDD1.n1 B 0.054751f
C113 VDD1.t0 B 0.013915f
C114 VDD1.t1 B 0.013915f
C115 VDD1.n2 B 0.054751f
C116 VDD1.n3 B 1.3548f
C117 VDD1.t4 B 0.013915f
C118 VDD1.t3 B 0.013915f
C119 VDD1.n4 B 0.05405f
C120 VDD1.n5 B 1.1732f
C121 VP.n0 B 0.025611f
C122 VP.t3 B 0.062195f
C123 VP.n1 B 0.04418f
C124 VP.n2 B 0.025611f
C125 VP.n3 B 0.028313f
C126 VP.n4 B 0.025611f
C127 VP.t4 B 0.062195f
C128 VP.n5 B 0.103962f
C129 VP.n6 B 0.025611f
C130 VP.t5 B 0.062195f
C131 VP.n7 B 0.04418f
C132 VP.n8 B 0.025611f
C133 VP.n9 B 0.028313f
C134 VP.t2 B 0.148865f
C135 VP.t1 B 0.062195f
C136 VP.n10 B 0.090726f
C137 VP.n11 B 0.090409f
C138 VP.n12 B 0.135895f
C139 VP.n13 B 0.025611f
C140 VP.n14 B 0.03755f
C141 VP.n15 B 0.03755f
C142 VP.t0 B 0.062195f
C143 VP.n16 B 0.055103f
C144 VP.n17 B 0.028313f
C145 VP.n18 B 0.025611f
C146 VP.n19 B 0.025611f
C147 VP.n20 B 0.025611f
C148 VP.n21 B 0.022928f
C149 VP.n22 B 0.040332f
C150 VP.n23 B 0.103962f
C151 VP.n24 B 0.833073f
C152 VP.n25 B 0.858171f
C153 VP.n26 B 0.025611f
C154 VP.n27 B 0.040332f
C155 VP.n28 B 0.022928f
C156 VP.t7 B 0.062195f
C157 VP.n29 B 0.055103f
C158 VP.n30 B 0.04418f
C159 VP.n31 B 0.025611f
C160 VP.n32 B 0.025611f
C161 VP.n33 B 0.025611f
C162 VP.n34 B 0.03755f
C163 VP.n35 B 0.03755f
C164 VP.t6 B 0.062195f
C165 VP.n36 B 0.055103f
C166 VP.n37 B 0.028313f
C167 VP.n38 B 0.025611f
C168 VP.n39 B 0.025611f
C169 VP.n40 B 0.025611f
C170 VP.n41 B 0.022928f
C171 VP.n42 B 0.040332f
C172 VP.n43 B 0.103962f
C173 VP.n44 B 0.023461f
.ends

