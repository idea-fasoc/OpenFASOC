* NGSPICE file created from diff_pair_sample_1539.ext - technology: sky130A

.subckt diff_pair_sample_1539 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X1 VDD1.t7 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.34
X2 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X3 VTAIL.t7 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X4 VTAIL.t14 VN.t1 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.34
X5 VDD1.t4 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.34
X6 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.34
X7 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.34
X8 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.34
X9 VDD2.t6 VN.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.34
X10 VTAIL.t12 VN.t3 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X11 VTAIL.t11 VN.t4 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.34
X12 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X13 VDD2.t4 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.34
X14 VDD2.t3 VN.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.34
X16 VDD2.t1 VN.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X17 VTAIL.t6 VP.t6 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.34
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.34
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.34
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n56 161.3
R8 VN.n55 VN.n40 161.3
R9 VN.n54 VN.n53 161.3
R10 VN.n52 VN.n41 161.3
R11 VN.n51 VN.n50 161.3
R12 VN.n49 VN.n42 161.3
R13 VN.n48 VN.n47 161.3
R14 VN.n46 VN.n43 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n21 161.3
R23 VN.n20 VN.n5 161.3
R24 VN.n19 VN.n18 161.3
R25 VN.n17 VN.n6 161.3
R26 VN.n16 VN.n15 161.3
R27 VN.n14 VN.n7 161.3
R28 VN.n13 VN.n12 161.3
R29 VN.n11 VN.n8 161.3
R30 VN.n45 VN.t5 112.716
R31 VN.n10 VN.t4 112.716
R32 VN.n9 VN.t7 80.1655
R33 VN.n4 VN.t0 80.1655
R34 VN.n0 VN.t2 80.1655
R35 VN.n44 VN.t3 80.1655
R36 VN.n39 VN.t6 80.1655
R37 VN.n35 VN.t1 80.1655
R38 VN.n34 VN.n0 77.5892
R39 VN.n69 VN.n35 77.5892
R40 VN.n10 VN.n9 70.4248
R41 VN.n45 VN.n44 70.4248
R42 VN.n15 VN.n6 56.5193
R43 VN.n50 VN.n41 56.5193
R44 VN VN.n69 53.9374
R45 VN.n26 VN.n2 48.2635
R46 VN.n61 VN.n37 48.2635
R47 VN.n30 VN.n2 32.7233
R48 VN.n65 VN.n37 32.7233
R49 VN.n13 VN.n8 24.4675
R50 VN.n14 VN.n13 24.4675
R51 VN.n15 VN.n14 24.4675
R52 VN.n19 VN.n6 24.4675
R53 VN.n20 VN.n19 24.4675
R54 VN.n21 VN.n20 24.4675
R55 VN.n25 VN.n24 24.4675
R56 VN.n26 VN.n25 24.4675
R57 VN.n31 VN.n30 24.4675
R58 VN.n32 VN.n31 24.4675
R59 VN.n50 VN.n49 24.4675
R60 VN.n49 VN.n48 24.4675
R61 VN.n48 VN.n43 24.4675
R62 VN.n61 VN.n60 24.4675
R63 VN.n60 VN.n59 24.4675
R64 VN.n56 VN.n55 24.4675
R65 VN.n55 VN.n54 24.4675
R66 VN.n54 VN.n41 24.4675
R67 VN.n67 VN.n66 24.4675
R68 VN.n66 VN.n65 24.4675
R69 VN.n24 VN.n4 20.3081
R70 VN.n59 VN.n39 20.3081
R71 VN.n32 VN.n0 12.4787
R72 VN.n67 VN.n35 12.4787
R73 VN.n46 VN.n45 4.27761
R74 VN.n11 VN.n10 4.27761
R75 VN.n9 VN.n8 4.15989
R76 VN.n21 VN.n4 4.15989
R77 VN.n44 VN.n43 4.15989
R78 VN.n56 VN.n39 4.15989
R79 VN.n69 VN.n68 0.354971
R80 VN.n34 VN.n33 0.354971
R81 VN VN.n34 0.26696
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n40 0.189894
R90 VN.n53 VN.n40 0.189894
R91 VN.n53 VN.n52 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n42 0.189894
R94 VN.n47 VN.n42 0.189894
R95 VN.n47 VN.n46 0.189894
R96 VN.n12 VN.n11 0.189894
R97 VN.n12 VN.n7 0.189894
R98 VN.n16 VN.n7 0.189894
R99 VN.n17 VN.n16 0.189894
R100 VN.n18 VN.n17 0.189894
R101 VN.n18 VN.n5 0.189894
R102 VN.n22 VN.n5 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VDD2.n2 VDD2.n1 65.093
R111 VDD2.n2 VDD2.n0 65.093
R112 VDD2 VDD2.n5 65.0903
R113 VDD2.n4 VDD2.n3 63.5667
R114 VDD2.n4 VDD2.n2 47.5299
R115 VDD2.n5 VDD2.t2 1.78268
R116 VDD2.n5 VDD2.t4 1.78268
R117 VDD2.n3 VDD2.t7 1.78268
R118 VDD2.n3 VDD2.t3 1.78268
R119 VDD2.n1 VDD2.t5 1.78268
R120 VDD2.n1 VDD2.t6 1.78268
R121 VDD2.n0 VDD2.t0 1.78268
R122 VDD2.n0 VDD2.t1 1.78268
R123 VDD2 VDD2.n4 1.64059
R124 VTAIL.n11 VTAIL.t0 48.67
R125 VTAIL.n10 VTAIL.t10 48.67
R126 VTAIL.n7 VTAIL.t14 48.67
R127 VTAIL.n15 VTAIL.t13 48.6699
R128 VTAIL.n2 VTAIL.t11 48.6699
R129 VTAIL.n3 VTAIL.t4 48.6699
R130 VTAIL.n6 VTAIL.t1 48.6699
R131 VTAIL.n14 VTAIL.t3 48.6699
R132 VTAIL.n13 VTAIL.n12 46.8879
R133 VTAIL.n9 VTAIL.n8 46.8879
R134 VTAIL.n1 VTAIL.n0 46.8877
R135 VTAIL.n5 VTAIL.n4 46.8877
R136 VTAIL.n15 VTAIL.n14 25.1083
R137 VTAIL.n7 VTAIL.n6 25.1083
R138 VTAIL.n9 VTAIL.n7 3.16429
R139 VTAIL.n10 VTAIL.n9 3.16429
R140 VTAIL.n13 VTAIL.n11 3.16429
R141 VTAIL.n14 VTAIL.n13 3.16429
R142 VTAIL.n6 VTAIL.n5 3.16429
R143 VTAIL.n5 VTAIL.n3 3.16429
R144 VTAIL.n2 VTAIL.n1 3.16429
R145 VTAIL VTAIL.n15 3.1061
R146 VTAIL.n0 VTAIL.t8 1.78268
R147 VTAIL.n0 VTAIL.t15 1.78268
R148 VTAIL.n4 VTAIL.t5 1.78268
R149 VTAIL.n4 VTAIL.t6 1.78268
R150 VTAIL.n12 VTAIL.t2 1.78268
R151 VTAIL.n12 VTAIL.t7 1.78268
R152 VTAIL.n8 VTAIL.t9 1.78268
R153 VTAIL.n8 VTAIL.t12 1.78268
R154 VTAIL.n11 VTAIL.n10 0.470328
R155 VTAIL.n3 VTAIL.n2 0.470328
R156 VTAIL VTAIL.n1 0.0586897
R157 B.n773 B.n772 585
R158 B.n775 B.n161 585
R159 B.n778 B.n777 585
R160 B.n779 B.n160 585
R161 B.n781 B.n780 585
R162 B.n783 B.n159 585
R163 B.n786 B.n785 585
R164 B.n787 B.n158 585
R165 B.n789 B.n788 585
R166 B.n791 B.n157 585
R167 B.n794 B.n793 585
R168 B.n795 B.n156 585
R169 B.n797 B.n796 585
R170 B.n799 B.n155 585
R171 B.n802 B.n801 585
R172 B.n803 B.n154 585
R173 B.n805 B.n804 585
R174 B.n807 B.n153 585
R175 B.n810 B.n809 585
R176 B.n811 B.n152 585
R177 B.n813 B.n812 585
R178 B.n815 B.n151 585
R179 B.n818 B.n817 585
R180 B.n819 B.n150 585
R181 B.n821 B.n820 585
R182 B.n823 B.n149 585
R183 B.n826 B.n825 585
R184 B.n827 B.n148 585
R185 B.n829 B.n828 585
R186 B.n831 B.n147 585
R187 B.n834 B.n833 585
R188 B.n835 B.n146 585
R189 B.n837 B.n836 585
R190 B.n839 B.n145 585
R191 B.n842 B.n841 585
R192 B.n843 B.n144 585
R193 B.n845 B.n844 585
R194 B.n847 B.n143 585
R195 B.n850 B.n849 585
R196 B.n852 B.n140 585
R197 B.n854 B.n853 585
R198 B.n856 B.n139 585
R199 B.n859 B.n858 585
R200 B.n860 B.n138 585
R201 B.n862 B.n861 585
R202 B.n864 B.n137 585
R203 B.n867 B.n866 585
R204 B.n868 B.n133 585
R205 B.n870 B.n869 585
R206 B.n872 B.n132 585
R207 B.n875 B.n874 585
R208 B.n876 B.n131 585
R209 B.n878 B.n877 585
R210 B.n880 B.n130 585
R211 B.n883 B.n882 585
R212 B.n884 B.n129 585
R213 B.n886 B.n885 585
R214 B.n888 B.n128 585
R215 B.n891 B.n890 585
R216 B.n892 B.n127 585
R217 B.n894 B.n893 585
R218 B.n896 B.n126 585
R219 B.n899 B.n898 585
R220 B.n900 B.n125 585
R221 B.n902 B.n901 585
R222 B.n904 B.n124 585
R223 B.n907 B.n906 585
R224 B.n908 B.n123 585
R225 B.n910 B.n909 585
R226 B.n912 B.n122 585
R227 B.n915 B.n914 585
R228 B.n916 B.n121 585
R229 B.n918 B.n917 585
R230 B.n920 B.n120 585
R231 B.n923 B.n922 585
R232 B.n924 B.n119 585
R233 B.n926 B.n925 585
R234 B.n928 B.n118 585
R235 B.n931 B.n930 585
R236 B.n932 B.n117 585
R237 B.n934 B.n933 585
R238 B.n936 B.n116 585
R239 B.n939 B.n938 585
R240 B.n940 B.n115 585
R241 B.n942 B.n941 585
R242 B.n944 B.n114 585
R243 B.n947 B.n946 585
R244 B.n948 B.n113 585
R245 B.n771 B.n111 585
R246 B.n951 B.n111 585
R247 B.n770 B.n110 585
R248 B.n952 B.n110 585
R249 B.n769 B.n109 585
R250 B.n953 B.n109 585
R251 B.n768 B.n767 585
R252 B.n767 B.n105 585
R253 B.n766 B.n104 585
R254 B.n959 B.n104 585
R255 B.n765 B.n103 585
R256 B.n960 B.n103 585
R257 B.n764 B.n102 585
R258 B.n961 B.n102 585
R259 B.n763 B.n762 585
R260 B.n762 B.n98 585
R261 B.n761 B.n97 585
R262 B.n967 B.n97 585
R263 B.n760 B.n96 585
R264 B.n968 B.n96 585
R265 B.n759 B.n95 585
R266 B.n969 B.n95 585
R267 B.n758 B.n757 585
R268 B.n757 B.n91 585
R269 B.n756 B.n90 585
R270 B.n975 B.n90 585
R271 B.n755 B.n89 585
R272 B.n976 B.n89 585
R273 B.n754 B.n88 585
R274 B.n977 B.n88 585
R275 B.n753 B.n752 585
R276 B.n752 B.n84 585
R277 B.n751 B.n83 585
R278 B.n983 B.n83 585
R279 B.n750 B.n82 585
R280 B.n984 B.n82 585
R281 B.n749 B.n81 585
R282 B.n985 B.n81 585
R283 B.n748 B.n747 585
R284 B.n747 B.n77 585
R285 B.n746 B.n76 585
R286 B.n991 B.n76 585
R287 B.n745 B.n75 585
R288 B.n992 B.n75 585
R289 B.n744 B.n74 585
R290 B.n993 B.n74 585
R291 B.n743 B.n742 585
R292 B.n742 B.n70 585
R293 B.n741 B.n69 585
R294 B.n999 B.n69 585
R295 B.n740 B.n68 585
R296 B.n1000 B.n68 585
R297 B.n739 B.n67 585
R298 B.n1001 B.n67 585
R299 B.n738 B.n737 585
R300 B.n737 B.n63 585
R301 B.n736 B.n62 585
R302 B.n1007 B.n62 585
R303 B.n735 B.n61 585
R304 B.n1008 B.n61 585
R305 B.n734 B.n60 585
R306 B.n1009 B.n60 585
R307 B.n733 B.n732 585
R308 B.n732 B.n56 585
R309 B.n731 B.n55 585
R310 B.n1015 B.n55 585
R311 B.n730 B.n54 585
R312 B.n1016 B.n54 585
R313 B.n729 B.n53 585
R314 B.n1017 B.n53 585
R315 B.n728 B.n727 585
R316 B.n727 B.n49 585
R317 B.n726 B.n48 585
R318 B.n1023 B.n48 585
R319 B.n725 B.n47 585
R320 B.n1024 B.n47 585
R321 B.n724 B.n46 585
R322 B.n1025 B.n46 585
R323 B.n723 B.n722 585
R324 B.n722 B.n42 585
R325 B.n721 B.n41 585
R326 B.n1031 B.n41 585
R327 B.n720 B.n40 585
R328 B.n1032 B.n40 585
R329 B.n719 B.n39 585
R330 B.n1033 B.n39 585
R331 B.n718 B.n717 585
R332 B.n717 B.n35 585
R333 B.n716 B.n34 585
R334 B.n1039 B.n34 585
R335 B.n715 B.n33 585
R336 B.n1040 B.n33 585
R337 B.n714 B.n32 585
R338 B.n1041 B.n32 585
R339 B.n713 B.n712 585
R340 B.n712 B.n28 585
R341 B.n711 B.n27 585
R342 B.n1047 B.n27 585
R343 B.n710 B.n26 585
R344 B.n1048 B.n26 585
R345 B.n709 B.n25 585
R346 B.n1049 B.n25 585
R347 B.n708 B.n707 585
R348 B.n707 B.n21 585
R349 B.n706 B.n20 585
R350 B.n1055 B.n20 585
R351 B.n705 B.n19 585
R352 B.n1056 B.n19 585
R353 B.n704 B.n18 585
R354 B.n1057 B.n18 585
R355 B.n703 B.n702 585
R356 B.n702 B.t0 585
R357 B.n701 B.n14 585
R358 B.n1063 B.n14 585
R359 B.n700 B.n13 585
R360 B.n1064 B.n13 585
R361 B.n699 B.n12 585
R362 B.n1065 B.n12 585
R363 B.n698 B.n697 585
R364 B.n697 B.n8 585
R365 B.n696 B.n7 585
R366 B.n1071 B.n7 585
R367 B.n695 B.n6 585
R368 B.n1072 B.n6 585
R369 B.n694 B.n5 585
R370 B.n1073 B.n5 585
R371 B.n693 B.n692 585
R372 B.n692 B.n4 585
R373 B.n691 B.n162 585
R374 B.n691 B.n690 585
R375 B.n681 B.n163 585
R376 B.n164 B.n163 585
R377 B.n683 B.n682 585
R378 B.n684 B.n683 585
R379 B.n680 B.n169 585
R380 B.n169 B.n168 585
R381 B.n679 B.n678 585
R382 B.n678 B.n677 585
R383 B.n171 B.n170 585
R384 B.t4 B.n171 585
R385 B.n670 B.n669 585
R386 B.n671 B.n670 585
R387 B.n668 B.n176 585
R388 B.n176 B.n175 585
R389 B.n667 B.n666 585
R390 B.n666 B.n665 585
R391 B.n178 B.n177 585
R392 B.n179 B.n178 585
R393 B.n658 B.n657 585
R394 B.n659 B.n658 585
R395 B.n656 B.n184 585
R396 B.n184 B.n183 585
R397 B.n655 B.n654 585
R398 B.n654 B.n653 585
R399 B.n186 B.n185 585
R400 B.n187 B.n186 585
R401 B.n646 B.n645 585
R402 B.n647 B.n646 585
R403 B.n644 B.n192 585
R404 B.n192 B.n191 585
R405 B.n643 B.n642 585
R406 B.n642 B.n641 585
R407 B.n194 B.n193 585
R408 B.n195 B.n194 585
R409 B.n634 B.n633 585
R410 B.n635 B.n634 585
R411 B.n632 B.n200 585
R412 B.n200 B.n199 585
R413 B.n631 B.n630 585
R414 B.n630 B.n629 585
R415 B.n202 B.n201 585
R416 B.n203 B.n202 585
R417 B.n622 B.n621 585
R418 B.n623 B.n622 585
R419 B.n620 B.n208 585
R420 B.n208 B.n207 585
R421 B.n619 B.n618 585
R422 B.n618 B.n617 585
R423 B.n210 B.n209 585
R424 B.n211 B.n210 585
R425 B.n610 B.n609 585
R426 B.n611 B.n610 585
R427 B.n608 B.n215 585
R428 B.n219 B.n215 585
R429 B.n607 B.n606 585
R430 B.n606 B.n605 585
R431 B.n217 B.n216 585
R432 B.n218 B.n217 585
R433 B.n598 B.n597 585
R434 B.n599 B.n598 585
R435 B.n596 B.n224 585
R436 B.n224 B.n223 585
R437 B.n595 B.n594 585
R438 B.n594 B.n593 585
R439 B.n226 B.n225 585
R440 B.n227 B.n226 585
R441 B.n586 B.n585 585
R442 B.n587 B.n586 585
R443 B.n584 B.n232 585
R444 B.n232 B.n231 585
R445 B.n583 B.n582 585
R446 B.n582 B.n581 585
R447 B.n234 B.n233 585
R448 B.n235 B.n234 585
R449 B.n574 B.n573 585
R450 B.n575 B.n574 585
R451 B.n572 B.n240 585
R452 B.n240 B.n239 585
R453 B.n571 B.n570 585
R454 B.n570 B.n569 585
R455 B.n242 B.n241 585
R456 B.n243 B.n242 585
R457 B.n562 B.n561 585
R458 B.n563 B.n562 585
R459 B.n560 B.n248 585
R460 B.n248 B.n247 585
R461 B.n559 B.n558 585
R462 B.n558 B.n557 585
R463 B.n250 B.n249 585
R464 B.n251 B.n250 585
R465 B.n550 B.n549 585
R466 B.n551 B.n550 585
R467 B.n548 B.n256 585
R468 B.n256 B.n255 585
R469 B.n547 B.n546 585
R470 B.n546 B.n545 585
R471 B.n258 B.n257 585
R472 B.n259 B.n258 585
R473 B.n538 B.n537 585
R474 B.n539 B.n538 585
R475 B.n536 B.n264 585
R476 B.n264 B.n263 585
R477 B.n535 B.n534 585
R478 B.n534 B.n533 585
R479 B.n266 B.n265 585
R480 B.n267 B.n266 585
R481 B.n526 B.n525 585
R482 B.n527 B.n526 585
R483 B.n524 B.n272 585
R484 B.n272 B.n271 585
R485 B.n523 B.n522 585
R486 B.n522 B.n521 585
R487 B.n274 B.n273 585
R488 B.n275 B.n274 585
R489 B.n514 B.n513 585
R490 B.n515 B.n514 585
R491 B.n512 B.n280 585
R492 B.n280 B.n279 585
R493 B.n511 B.n510 585
R494 B.n510 B.n509 585
R495 B.n506 B.n284 585
R496 B.n505 B.n504 585
R497 B.n502 B.n285 585
R498 B.n502 B.n283 585
R499 B.n501 B.n500 585
R500 B.n499 B.n498 585
R501 B.n497 B.n287 585
R502 B.n495 B.n494 585
R503 B.n493 B.n288 585
R504 B.n492 B.n491 585
R505 B.n489 B.n289 585
R506 B.n487 B.n486 585
R507 B.n485 B.n290 585
R508 B.n484 B.n483 585
R509 B.n481 B.n291 585
R510 B.n479 B.n478 585
R511 B.n477 B.n292 585
R512 B.n476 B.n475 585
R513 B.n473 B.n293 585
R514 B.n471 B.n470 585
R515 B.n469 B.n294 585
R516 B.n468 B.n467 585
R517 B.n465 B.n295 585
R518 B.n463 B.n462 585
R519 B.n461 B.n296 585
R520 B.n460 B.n459 585
R521 B.n457 B.n297 585
R522 B.n455 B.n454 585
R523 B.n453 B.n298 585
R524 B.n452 B.n451 585
R525 B.n449 B.n299 585
R526 B.n447 B.n446 585
R527 B.n445 B.n300 585
R528 B.n444 B.n443 585
R529 B.n441 B.n301 585
R530 B.n439 B.n438 585
R531 B.n437 B.n302 585
R532 B.n436 B.n435 585
R533 B.n433 B.n303 585
R534 B.n431 B.n430 585
R535 B.n428 B.n304 585
R536 B.n427 B.n426 585
R537 B.n424 B.n307 585
R538 B.n422 B.n421 585
R539 B.n420 B.n308 585
R540 B.n419 B.n418 585
R541 B.n416 B.n309 585
R542 B.n414 B.n413 585
R543 B.n412 B.n310 585
R544 B.n411 B.n410 585
R545 B.n408 B.n407 585
R546 B.n406 B.n405 585
R547 B.n404 B.n315 585
R548 B.n402 B.n401 585
R549 B.n400 B.n316 585
R550 B.n399 B.n398 585
R551 B.n396 B.n317 585
R552 B.n394 B.n393 585
R553 B.n392 B.n318 585
R554 B.n391 B.n390 585
R555 B.n388 B.n319 585
R556 B.n386 B.n385 585
R557 B.n384 B.n320 585
R558 B.n383 B.n382 585
R559 B.n380 B.n321 585
R560 B.n378 B.n377 585
R561 B.n376 B.n322 585
R562 B.n375 B.n374 585
R563 B.n372 B.n323 585
R564 B.n370 B.n369 585
R565 B.n368 B.n324 585
R566 B.n367 B.n366 585
R567 B.n364 B.n325 585
R568 B.n362 B.n361 585
R569 B.n360 B.n326 585
R570 B.n359 B.n358 585
R571 B.n356 B.n327 585
R572 B.n354 B.n353 585
R573 B.n352 B.n328 585
R574 B.n351 B.n350 585
R575 B.n348 B.n329 585
R576 B.n346 B.n345 585
R577 B.n344 B.n330 585
R578 B.n343 B.n342 585
R579 B.n340 B.n331 585
R580 B.n338 B.n337 585
R581 B.n336 B.n332 585
R582 B.n335 B.n334 585
R583 B.n282 B.n281 585
R584 B.n283 B.n282 585
R585 B.n508 B.n507 585
R586 B.n509 B.n508 585
R587 B.n278 B.n277 585
R588 B.n279 B.n278 585
R589 B.n517 B.n516 585
R590 B.n516 B.n515 585
R591 B.n518 B.n276 585
R592 B.n276 B.n275 585
R593 B.n520 B.n519 585
R594 B.n521 B.n520 585
R595 B.n270 B.n269 585
R596 B.n271 B.n270 585
R597 B.n529 B.n528 585
R598 B.n528 B.n527 585
R599 B.n530 B.n268 585
R600 B.n268 B.n267 585
R601 B.n532 B.n531 585
R602 B.n533 B.n532 585
R603 B.n262 B.n261 585
R604 B.n263 B.n262 585
R605 B.n541 B.n540 585
R606 B.n540 B.n539 585
R607 B.n542 B.n260 585
R608 B.n260 B.n259 585
R609 B.n544 B.n543 585
R610 B.n545 B.n544 585
R611 B.n254 B.n253 585
R612 B.n255 B.n254 585
R613 B.n553 B.n552 585
R614 B.n552 B.n551 585
R615 B.n554 B.n252 585
R616 B.n252 B.n251 585
R617 B.n556 B.n555 585
R618 B.n557 B.n556 585
R619 B.n246 B.n245 585
R620 B.n247 B.n246 585
R621 B.n565 B.n564 585
R622 B.n564 B.n563 585
R623 B.n566 B.n244 585
R624 B.n244 B.n243 585
R625 B.n568 B.n567 585
R626 B.n569 B.n568 585
R627 B.n238 B.n237 585
R628 B.n239 B.n238 585
R629 B.n577 B.n576 585
R630 B.n576 B.n575 585
R631 B.n578 B.n236 585
R632 B.n236 B.n235 585
R633 B.n580 B.n579 585
R634 B.n581 B.n580 585
R635 B.n230 B.n229 585
R636 B.n231 B.n230 585
R637 B.n589 B.n588 585
R638 B.n588 B.n587 585
R639 B.n590 B.n228 585
R640 B.n228 B.n227 585
R641 B.n592 B.n591 585
R642 B.n593 B.n592 585
R643 B.n222 B.n221 585
R644 B.n223 B.n222 585
R645 B.n601 B.n600 585
R646 B.n600 B.n599 585
R647 B.n602 B.n220 585
R648 B.n220 B.n218 585
R649 B.n604 B.n603 585
R650 B.n605 B.n604 585
R651 B.n214 B.n213 585
R652 B.n219 B.n214 585
R653 B.n613 B.n612 585
R654 B.n612 B.n611 585
R655 B.n614 B.n212 585
R656 B.n212 B.n211 585
R657 B.n616 B.n615 585
R658 B.n617 B.n616 585
R659 B.n206 B.n205 585
R660 B.n207 B.n206 585
R661 B.n625 B.n624 585
R662 B.n624 B.n623 585
R663 B.n626 B.n204 585
R664 B.n204 B.n203 585
R665 B.n628 B.n627 585
R666 B.n629 B.n628 585
R667 B.n198 B.n197 585
R668 B.n199 B.n198 585
R669 B.n637 B.n636 585
R670 B.n636 B.n635 585
R671 B.n638 B.n196 585
R672 B.n196 B.n195 585
R673 B.n640 B.n639 585
R674 B.n641 B.n640 585
R675 B.n190 B.n189 585
R676 B.n191 B.n190 585
R677 B.n649 B.n648 585
R678 B.n648 B.n647 585
R679 B.n650 B.n188 585
R680 B.n188 B.n187 585
R681 B.n652 B.n651 585
R682 B.n653 B.n652 585
R683 B.n182 B.n181 585
R684 B.n183 B.n182 585
R685 B.n661 B.n660 585
R686 B.n660 B.n659 585
R687 B.n662 B.n180 585
R688 B.n180 B.n179 585
R689 B.n664 B.n663 585
R690 B.n665 B.n664 585
R691 B.n174 B.n173 585
R692 B.n175 B.n174 585
R693 B.n673 B.n672 585
R694 B.n672 B.n671 585
R695 B.n674 B.n172 585
R696 B.n172 B.t4 585
R697 B.n676 B.n675 585
R698 B.n677 B.n676 585
R699 B.n167 B.n166 585
R700 B.n168 B.n167 585
R701 B.n686 B.n685 585
R702 B.n685 B.n684 585
R703 B.n687 B.n165 585
R704 B.n165 B.n164 585
R705 B.n689 B.n688 585
R706 B.n690 B.n689 585
R707 B.n2 B.n0 585
R708 B.n4 B.n2 585
R709 B.n3 B.n1 585
R710 B.n1072 B.n3 585
R711 B.n1070 B.n1069 585
R712 B.n1071 B.n1070 585
R713 B.n1068 B.n9 585
R714 B.n9 B.n8 585
R715 B.n1067 B.n1066 585
R716 B.n1066 B.n1065 585
R717 B.n11 B.n10 585
R718 B.n1064 B.n11 585
R719 B.n1062 B.n1061 585
R720 B.n1063 B.n1062 585
R721 B.n1060 B.n15 585
R722 B.n15 B.t0 585
R723 B.n1059 B.n1058 585
R724 B.n1058 B.n1057 585
R725 B.n17 B.n16 585
R726 B.n1056 B.n17 585
R727 B.n1054 B.n1053 585
R728 B.n1055 B.n1054 585
R729 B.n1052 B.n22 585
R730 B.n22 B.n21 585
R731 B.n1051 B.n1050 585
R732 B.n1050 B.n1049 585
R733 B.n24 B.n23 585
R734 B.n1048 B.n24 585
R735 B.n1046 B.n1045 585
R736 B.n1047 B.n1046 585
R737 B.n1044 B.n29 585
R738 B.n29 B.n28 585
R739 B.n1043 B.n1042 585
R740 B.n1042 B.n1041 585
R741 B.n31 B.n30 585
R742 B.n1040 B.n31 585
R743 B.n1038 B.n1037 585
R744 B.n1039 B.n1038 585
R745 B.n1036 B.n36 585
R746 B.n36 B.n35 585
R747 B.n1035 B.n1034 585
R748 B.n1034 B.n1033 585
R749 B.n38 B.n37 585
R750 B.n1032 B.n38 585
R751 B.n1030 B.n1029 585
R752 B.n1031 B.n1030 585
R753 B.n1028 B.n43 585
R754 B.n43 B.n42 585
R755 B.n1027 B.n1026 585
R756 B.n1026 B.n1025 585
R757 B.n45 B.n44 585
R758 B.n1024 B.n45 585
R759 B.n1022 B.n1021 585
R760 B.n1023 B.n1022 585
R761 B.n1020 B.n50 585
R762 B.n50 B.n49 585
R763 B.n1019 B.n1018 585
R764 B.n1018 B.n1017 585
R765 B.n52 B.n51 585
R766 B.n1016 B.n52 585
R767 B.n1014 B.n1013 585
R768 B.n1015 B.n1014 585
R769 B.n1012 B.n57 585
R770 B.n57 B.n56 585
R771 B.n1011 B.n1010 585
R772 B.n1010 B.n1009 585
R773 B.n59 B.n58 585
R774 B.n1008 B.n59 585
R775 B.n1006 B.n1005 585
R776 B.n1007 B.n1006 585
R777 B.n1004 B.n64 585
R778 B.n64 B.n63 585
R779 B.n1003 B.n1002 585
R780 B.n1002 B.n1001 585
R781 B.n66 B.n65 585
R782 B.n1000 B.n66 585
R783 B.n998 B.n997 585
R784 B.n999 B.n998 585
R785 B.n996 B.n71 585
R786 B.n71 B.n70 585
R787 B.n995 B.n994 585
R788 B.n994 B.n993 585
R789 B.n73 B.n72 585
R790 B.n992 B.n73 585
R791 B.n990 B.n989 585
R792 B.n991 B.n990 585
R793 B.n988 B.n78 585
R794 B.n78 B.n77 585
R795 B.n987 B.n986 585
R796 B.n986 B.n985 585
R797 B.n80 B.n79 585
R798 B.n984 B.n80 585
R799 B.n982 B.n981 585
R800 B.n983 B.n982 585
R801 B.n980 B.n85 585
R802 B.n85 B.n84 585
R803 B.n979 B.n978 585
R804 B.n978 B.n977 585
R805 B.n87 B.n86 585
R806 B.n976 B.n87 585
R807 B.n974 B.n973 585
R808 B.n975 B.n974 585
R809 B.n972 B.n92 585
R810 B.n92 B.n91 585
R811 B.n971 B.n970 585
R812 B.n970 B.n969 585
R813 B.n94 B.n93 585
R814 B.n968 B.n94 585
R815 B.n966 B.n965 585
R816 B.n967 B.n966 585
R817 B.n964 B.n99 585
R818 B.n99 B.n98 585
R819 B.n963 B.n962 585
R820 B.n962 B.n961 585
R821 B.n101 B.n100 585
R822 B.n960 B.n101 585
R823 B.n958 B.n957 585
R824 B.n959 B.n958 585
R825 B.n956 B.n106 585
R826 B.n106 B.n105 585
R827 B.n955 B.n954 585
R828 B.n954 B.n953 585
R829 B.n108 B.n107 585
R830 B.n952 B.n108 585
R831 B.n950 B.n949 585
R832 B.n951 B.n950 585
R833 B.n1075 B.n1074 585
R834 B.n1074 B.n1073 585
R835 B.n508 B.n284 478.086
R836 B.n950 B.n113 478.086
R837 B.n510 B.n282 478.086
R838 B.n773 B.n111 478.086
R839 B.n311 B.t12 289.11
R840 B.n305 B.t19 289.11
R841 B.n134 B.t16 289.11
R842 B.n141 B.t8 289.11
R843 B.n774 B.n112 256.663
R844 B.n776 B.n112 256.663
R845 B.n782 B.n112 256.663
R846 B.n784 B.n112 256.663
R847 B.n790 B.n112 256.663
R848 B.n792 B.n112 256.663
R849 B.n798 B.n112 256.663
R850 B.n800 B.n112 256.663
R851 B.n806 B.n112 256.663
R852 B.n808 B.n112 256.663
R853 B.n814 B.n112 256.663
R854 B.n816 B.n112 256.663
R855 B.n822 B.n112 256.663
R856 B.n824 B.n112 256.663
R857 B.n830 B.n112 256.663
R858 B.n832 B.n112 256.663
R859 B.n838 B.n112 256.663
R860 B.n840 B.n112 256.663
R861 B.n846 B.n112 256.663
R862 B.n848 B.n112 256.663
R863 B.n855 B.n112 256.663
R864 B.n857 B.n112 256.663
R865 B.n863 B.n112 256.663
R866 B.n865 B.n112 256.663
R867 B.n871 B.n112 256.663
R868 B.n873 B.n112 256.663
R869 B.n879 B.n112 256.663
R870 B.n881 B.n112 256.663
R871 B.n887 B.n112 256.663
R872 B.n889 B.n112 256.663
R873 B.n895 B.n112 256.663
R874 B.n897 B.n112 256.663
R875 B.n903 B.n112 256.663
R876 B.n905 B.n112 256.663
R877 B.n911 B.n112 256.663
R878 B.n913 B.n112 256.663
R879 B.n919 B.n112 256.663
R880 B.n921 B.n112 256.663
R881 B.n927 B.n112 256.663
R882 B.n929 B.n112 256.663
R883 B.n935 B.n112 256.663
R884 B.n937 B.n112 256.663
R885 B.n943 B.n112 256.663
R886 B.n945 B.n112 256.663
R887 B.n503 B.n283 256.663
R888 B.n286 B.n283 256.663
R889 B.n496 B.n283 256.663
R890 B.n490 B.n283 256.663
R891 B.n488 B.n283 256.663
R892 B.n482 B.n283 256.663
R893 B.n480 B.n283 256.663
R894 B.n474 B.n283 256.663
R895 B.n472 B.n283 256.663
R896 B.n466 B.n283 256.663
R897 B.n464 B.n283 256.663
R898 B.n458 B.n283 256.663
R899 B.n456 B.n283 256.663
R900 B.n450 B.n283 256.663
R901 B.n448 B.n283 256.663
R902 B.n442 B.n283 256.663
R903 B.n440 B.n283 256.663
R904 B.n434 B.n283 256.663
R905 B.n432 B.n283 256.663
R906 B.n425 B.n283 256.663
R907 B.n423 B.n283 256.663
R908 B.n417 B.n283 256.663
R909 B.n415 B.n283 256.663
R910 B.n409 B.n283 256.663
R911 B.n314 B.n283 256.663
R912 B.n403 B.n283 256.663
R913 B.n397 B.n283 256.663
R914 B.n395 B.n283 256.663
R915 B.n389 B.n283 256.663
R916 B.n387 B.n283 256.663
R917 B.n381 B.n283 256.663
R918 B.n379 B.n283 256.663
R919 B.n373 B.n283 256.663
R920 B.n371 B.n283 256.663
R921 B.n365 B.n283 256.663
R922 B.n363 B.n283 256.663
R923 B.n357 B.n283 256.663
R924 B.n355 B.n283 256.663
R925 B.n349 B.n283 256.663
R926 B.n347 B.n283 256.663
R927 B.n341 B.n283 256.663
R928 B.n339 B.n283 256.663
R929 B.n333 B.n283 256.663
R930 B.n508 B.n278 163.367
R931 B.n516 B.n278 163.367
R932 B.n516 B.n276 163.367
R933 B.n520 B.n276 163.367
R934 B.n520 B.n270 163.367
R935 B.n528 B.n270 163.367
R936 B.n528 B.n268 163.367
R937 B.n532 B.n268 163.367
R938 B.n532 B.n262 163.367
R939 B.n540 B.n262 163.367
R940 B.n540 B.n260 163.367
R941 B.n544 B.n260 163.367
R942 B.n544 B.n254 163.367
R943 B.n552 B.n254 163.367
R944 B.n552 B.n252 163.367
R945 B.n556 B.n252 163.367
R946 B.n556 B.n246 163.367
R947 B.n564 B.n246 163.367
R948 B.n564 B.n244 163.367
R949 B.n568 B.n244 163.367
R950 B.n568 B.n238 163.367
R951 B.n576 B.n238 163.367
R952 B.n576 B.n236 163.367
R953 B.n580 B.n236 163.367
R954 B.n580 B.n230 163.367
R955 B.n588 B.n230 163.367
R956 B.n588 B.n228 163.367
R957 B.n592 B.n228 163.367
R958 B.n592 B.n222 163.367
R959 B.n600 B.n222 163.367
R960 B.n600 B.n220 163.367
R961 B.n604 B.n220 163.367
R962 B.n604 B.n214 163.367
R963 B.n612 B.n214 163.367
R964 B.n612 B.n212 163.367
R965 B.n616 B.n212 163.367
R966 B.n616 B.n206 163.367
R967 B.n624 B.n206 163.367
R968 B.n624 B.n204 163.367
R969 B.n628 B.n204 163.367
R970 B.n628 B.n198 163.367
R971 B.n636 B.n198 163.367
R972 B.n636 B.n196 163.367
R973 B.n640 B.n196 163.367
R974 B.n640 B.n190 163.367
R975 B.n648 B.n190 163.367
R976 B.n648 B.n188 163.367
R977 B.n652 B.n188 163.367
R978 B.n652 B.n182 163.367
R979 B.n660 B.n182 163.367
R980 B.n660 B.n180 163.367
R981 B.n664 B.n180 163.367
R982 B.n664 B.n174 163.367
R983 B.n672 B.n174 163.367
R984 B.n672 B.n172 163.367
R985 B.n676 B.n172 163.367
R986 B.n676 B.n167 163.367
R987 B.n685 B.n167 163.367
R988 B.n685 B.n165 163.367
R989 B.n689 B.n165 163.367
R990 B.n689 B.n2 163.367
R991 B.n1074 B.n2 163.367
R992 B.n1074 B.n3 163.367
R993 B.n1070 B.n3 163.367
R994 B.n1070 B.n9 163.367
R995 B.n1066 B.n9 163.367
R996 B.n1066 B.n11 163.367
R997 B.n1062 B.n11 163.367
R998 B.n1062 B.n15 163.367
R999 B.n1058 B.n15 163.367
R1000 B.n1058 B.n17 163.367
R1001 B.n1054 B.n17 163.367
R1002 B.n1054 B.n22 163.367
R1003 B.n1050 B.n22 163.367
R1004 B.n1050 B.n24 163.367
R1005 B.n1046 B.n24 163.367
R1006 B.n1046 B.n29 163.367
R1007 B.n1042 B.n29 163.367
R1008 B.n1042 B.n31 163.367
R1009 B.n1038 B.n31 163.367
R1010 B.n1038 B.n36 163.367
R1011 B.n1034 B.n36 163.367
R1012 B.n1034 B.n38 163.367
R1013 B.n1030 B.n38 163.367
R1014 B.n1030 B.n43 163.367
R1015 B.n1026 B.n43 163.367
R1016 B.n1026 B.n45 163.367
R1017 B.n1022 B.n45 163.367
R1018 B.n1022 B.n50 163.367
R1019 B.n1018 B.n50 163.367
R1020 B.n1018 B.n52 163.367
R1021 B.n1014 B.n52 163.367
R1022 B.n1014 B.n57 163.367
R1023 B.n1010 B.n57 163.367
R1024 B.n1010 B.n59 163.367
R1025 B.n1006 B.n59 163.367
R1026 B.n1006 B.n64 163.367
R1027 B.n1002 B.n64 163.367
R1028 B.n1002 B.n66 163.367
R1029 B.n998 B.n66 163.367
R1030 B.n998 B.n71 163.367
R1031 B.n994 B.n71 163.367
R1032 B.n994 B.n73 163.367
R1033 B.n990 B.n73 163.367
R1034 B.n990 B.n78 163.367
R1035 B.n986 B.n78 163.367
R1036 B.n986 B.n80 163.367
R1037 B.n982 B.n80 163.367
R1038 B.n982 B.n85 163.367
R1039 B.n978 B.n85 163.367
R1040 B.n978 B.n87 163.367
R1041 B.n974 B.n87 163.367
R1042 B.n974 B.n92 163.367
R1043 B.n970 B.n92 163.367
R1044 B.n970 B.n94 163.367
R1045 B.n966 B.n94 163.367
R1046 B.n966 B.n99 163.367
R1047 B.n962 B.n99 163.367
R1048 B.n962 B.n101 163.367
R1049 B.n958 B.n101 163.367
R1050 B.n958 B.n106 163.367
R1051 B.n954 B.n106 163.367
R1052 B.n954 B.n108 163.367
R1053 B.n950 B.n108 163.367
R1054 B.n504 B.n502 163.367
R1055 B.n502 B.n501 163.367
R1056 B.n498 B.n497 163.367
R1057 B.n495 B.n288 163.367
R1058 B.n491 B.n489 163.367
R1059 B.n487 B.n290 163.367
R1060 B.n483 B.n481 163.367
R1061 B.n479 B.n292 163.367
R1062 B.n475 B.n473 163.367
R1063 B.n471 B.n294 163.367
R1064 B.n467 B.n465 163.367
R1065 B.n463 B.n296 163.367
R1066 B.n459 B.n457 163.367
R1067 B.n455 B.n298 163.367
R1068 B.n451 B.n449 163.367
R1069 B.n447 B.n300 163.367
R1070 B.n443 B.n441 163.367
R1071 B.n439 B.n302 163.367
R1072 B.n435 B.n433 163.367
R1073 B.n431 B.n304 163.367
R1074 B.n426 B.n424 163.367
R1075 B.n422 B.n308 163.367
R1076 B.n418 B.n416 163.367
R1077 B.n414 B.n310 163.367
R1078 B.n410 B.n408 163.367
R1079 B.n405 B.n404 163.367
R1080 B.n402 B.n316 163.367
R1081 B.n398 B.n396 163.367
R1082 B.n394 B.n318 163.367
R1083 B.n390 B.n388 163.367
R1084 B.n386 B.n320 163.367
R1085 B.n382 B.n380 163.367
R1086 B.n378 B.n322 163.367
R1087 B.n374 B.n372 163.367
R1088 B.n370 B.n324 163.367
R1089 B.n366 B.n364 163.367
R1090 B.n362 B.n326 163.367
R1091 B.n358 B.n356 163.367
R1092 B.n354 B.n328 163.367
R1093 B.n350 B.n348 163.367
R1094 B.n346 B.n330 163.367
R1095 B.n342 B.n340 163.367
R1096 B.n338 B.n332 163.367
R1097 B.n334 B.n282 163.367
R1098 B.n510 B.n280 163.367
R1099 B.n514 B.n280 163.367
R1100 B.n514 B.n274 163.367
R1101 B.n522 B.n274 163.367
R1102 B.n522 B.n272 163.367
R1103 B.n526 B.n272 163.367
R1104 B.n526 B.n266 163.367
R1105 B.n534 B.n266 163.367
R1106 B.n534 B.n264 163.367
R1107 B.n538 B.n264 163.367
R1108 B.n538 B.n258 163.367
R1109 B.n546 B.n258 163.367
R1110 B.n546 B.n256 163.367
R1111 B.n550 B.n256 163.367
R1112 B.n550 B.n250 163.367
R1113 B.n558 B.n250 163.367
R1114 B.n558 B.n248 163.367
R1115 B.n562 B.n248 163.367
R1116 B.n562 B.n242 163.367
R1117 B.n570 B.n242 163.367
R1118 B.n570 B.n240 163.367
R1119 B.n574 B.n240 163.367
R1120 B.n574 B.n234 163.367
R1121 B.n582 B.n234 163.367
R1122 B.n582 B.n232 163.367
R1123 B.n586 B.n232 163.367
R1124 B.n586 B.n226 163.367
R1125 B.n594 B.n226 163.367
R1126 B.n594 B.n224 163.367
R1127 B.n598 B.n224 163.367
R1128 B.n598 B.n217 163.367
R1129 B.n606 B.n217 163.367
R1130 B.n606 B.n215 163.367
R1131 B.n610 B.n215 163.367
R1132 B.n610 B.n210 163.367
R1133 B.n618 B.n210 163.367
R1134 B.n618 B.n208 163.367
R1135 B.n622 B.n208 163.367
R1136 B.n622 B.n202 163.367
R1137 B.n630 B.n202 163.367
R1138 B.n630 B.n200 163.367
R1139 B.n634 B.n200 163.367
R1140 B.n634 B.n194 163.367
R1141 B.n642 B.n194 163.367
R1142 B.n642 B.n192 163.367
R1143 B.n646 B.n192 163.367
R1144 B.n646 B.n186 163.367
R1145 B.n654 B.n186 163.367
R1146 B.n654 B.n184 163.367
R1147 B.n658 B.n184 163.367
R1148 B.n658 B.n178 163.367
R1149 B.n666 B.n178 163.367
R1150 B.n666 B.n176 163.367
R1151 B.n670 B.n176 163.367
R1152 B.n670 B.n171 163.367
R1153 B.n678 B.n171 163.367
R1154 B.n678 B.n169 163.367
R1155 B.n683 B.n169 163.367
R1156 B.n683 B.n163 163.367
R1157 B.n691 B.n163 163.367
R1158 B.n692 B.n691 163.367
R1159 B.n692 B.n5 163.367
R1160 B.n6 B.n5 163.367
R1161 B.n7 B.n6 163.367
R1162 B.n697 B.n7 163.367
R1163 B.n697 B.n12 163.367
R1164 B.n13 B.n12 163.367
R1165 B.n14 B.n13 163.367
R1166 B.n702 B.n14 163.367
R1167 B.n702 B.n18 163.367
R1168 B.n19 B.n18 163.367
R1169 B.n20 B.n19 163.367
R1170 B.n707 B.n20 163.367
R1171 B.n707 B.n25 163.367
R1172 B.n26 B.n25 163.367
R1173 B.n27 B.n26 163.367
R1174 B.n712 B.n27 163.367
R1175 B.n712 B.n32 163.367
R1176 B.n33 B.n32 163.367
R1177 B.n34 B.n33 163.367
R1178 B.n717 B.n34 163.367
R1179 B.n717 B.n39 163.367
R1180 B.n40 B.n39 163.367
R1181 B.n41 B.n40 163.367
R1182 B.n722 B.n41 163.367
R1183 B.n722 B.n46 163.367
R1184 B.n47 B.n46 163.367
R1185 B.n48 B.n47 163.367
R1186 B.n727 B.n48 163.367
R1187 B.n727 B.n53 163.367
R1188 B.n54 B.n53 163.367
R1189 B.n55 B.n54 163.367
R1190 B.n732 B.n55 163.367
R1191 B.n732 B.n60 163.367
R1192 B.n61 B.n60 163.367
R1193 B.n62 B.n61 163.367
R1194 B.n737 B.n62 163.367
R1195 B.n737 B.n67 163.367
R1196 B.n68 B.n67 163.367
R1197 B.n69 B.n68 163.367
R1198 B.n742 B.n69 163.367
R1199 B.n742 B.n74 163.367
R1200 B.n75 B.n74 163.367
R1201 B.n76 B.n75 163.367
R1202 B.n747 B.n76 163.367
R1203 B.n747 B.n81 163.367
R1204 B.n82 B.n81 163.367
R1205 B.n83 B.n82 163.367
R1206 B.n752 B.n83 163.367
R1207 B.n752 B.n88 163.367
R1208 B.n89 B.n88 163.367
R1209 B.n90 B.n89 163.367
R1210 B.n757 B.n90 163.367
R1211 B.n757 B.n95 163.367
R1212 B.n96 B.n95 163.367
R1213 B.n97 B.n96 163.367
R1214 B.n762 B.n97 163.367
R1215 B.n762 B.n102 163.367
R1216 B.n103 B.n102 163.367
R1217 B.n104 B.n103 163.367
R1218 B.n767 B.n104 163.367
R1219 B.n767 B.n109 163.367
R1220 B.n110 B.n109 163.367
R1221 B.n111 B.n110 163.367
R1222 B.n946 B.n944 163.367
R1223 B.n942 B.n115 163.367
R1224 B.n938 B.n936 163.367
R1225 B.n934 B.n117 163.367
R1226 B.n930 B.n928 163.367
R1227 B.n926 B.n119 163.367
R1228 B.n922 B.n920 163.367
R1229 B.n918 B.n121 163.367
R1230 B.n914 B.n912 163.367
R1231 B.n910 B.n123 163.367
R1232 B.n906 B.n904 163.367
R1233 B.n902 B.n125 163.367
R1234 B.n898 B.n896 163.367
R1235 B.n894 B.n127 163.367
R1236 B.n890 B.n888 163.367
R1237 B.n886 B.n129 163.367
R1238 B.n882 B.n880 163.367
R1239 B.n878 B.n131 163.367
R1240 B.n874 B.n872 163.367
R1241 B.n870 B.n133 163.367
R1242 B.n866 B.n864 163.367
R1243 B.n862 B.n138 163.367
R1244 B.n858 B.n856 163.367
R1245 B.n854 B.n140 163.367
R1246 B.n849 B.n847 163.367
R1247 B.n845 B.n144 163.367
R1248 B.n841 B.n839 163.367
R1249 B.n837 B.n146 163.367
R1250 B.n833 B.n831 163.367
R1251 B.n829 B.n148 163.367
R1252 B.n825 B.n823 163.367
R1253 B.n821 B.n150 163.367
R1254 B.n817 B.n815 163.367
R1255 B.n813 B.n152 163.367
R1256 B.n809 B.n807 163.367
R1257 B.n805 B.n154 163.367
R1258 B.n801 B.n799 163.367
R1259 B.n797 B.n156 163.367
R1260 B.n793 B.n791 163.367
R1261 B.n789 B.n158 163.367
R1262 B.n785 B.n783 163.367
R1263 B.n781 B.n160 163.367
R1264 B.n777 B.n775 163.367
R1265 B.n311 B.t15 143.556
R1266 B.n141 B.t10 143.556
R1267 B.n305 B.t21 143.543
R1268 B.n134 B.t17 143.543
R1269 B.n509 B.n283 86.6041
R1270 B.n951 B.n112 86.6041
R1271 B.n312 B.t14 72.3812
R1272 B.n142 B.t11 72.3812
R1273 B.n306 B.t20 72.3675
R1274 B.n135 B.t18 72.3675
R1275 B.n503 B.n284 71.676
R1276 B.n501 B.n286 71.676
R1277 B.n497 B.n496 71.676
R1278 B.n490 B.n288 71.676
R1279 B.n489 B.n488 71.676
R1280 B.n482 B.n290 71.676
R1281 B.n481 B.n480 71.676
R1282 B.n474 B.n292 71.676
R1283 B.n473 B.n472 71.676
R1284 B.n466 B.n294 71.676
R1285 B.n465 B.n464 71.676
R1286 B.n458 B.n296 71.676
R1287 B.n457 B.n456 71.676
R1288 B.n450 B.n298 71.676
R1289 B.n449 B.n448 71.676
R1290 B.n442 B.n300 71.676
R1291 B.n441 B.n440 71.676
R1292 B.n434 B.n302 71.676
R1293 B.n433 B.n432 71.676
R1294 B.n425 B.n304 71.676
R1295 B.n424 B.n423 71.676
R1296 B.n417 B.n308 71.676
R1297 B.n416 B.n415 71.676
R1298 B.n409 B.n310 71.676
R1299 B.n408 B.n314 71.676
R1300 B.n404 B.n403 71.676
R1301 B.n397 B.n316 71.676
R1302 B.n396 B.n395 71.676
R1303 B.n389 B.n318 71.676
R1304 B.n388 B.n387 71.676
R1305 B.n381 B.n320 71.676
R1306 B.n380 B.n379 71.676
R1307 B.n373 B.n322 71.676
R1308 B.n372 B.n371 71.676
R1309 B.n365 B.n324 71.676
R1310 B.n364 B.n363 71.676
R1311 B.n357 B.n326 71.676
R1312 B.n356 B.n355 71.676
R1313 B.n349 B.n328 71.676
R1314 B.n348 B.n347 71.676
R1315 B.n341 B.n330 71.676
R1316 B.n340 B.n339 71.676
R1317 B.n333 B.n332 71.676
R1318 B.n945 B.n113 71.676
R1319 B.n944 B.n943 71.676
R1320 B.n937 B.n115 71.676
R1321 B.n936 B.n935 71.676
R1322 B.n929 B.n117 71.676
R1323 B.n928 B.n927 71.676
R1324 B.n921 B.n119 71.676
R1325 B.n920 B.n919 71.676
R1326 B.n913 B.n121 71.676
R1327 B.n912 B.n911 71.676
R1328 B.n905 B.n123 71.676
R1329 B.n904 B.n903 71.676
R1330 B.n897 B.n125 71.676
R1331 B.n896 B.n895 71.676
R1332 B.n889 B.n127 71.676
R1333 B.n888 B.n887 71.676
R1334 B.n881 B.n129 71.676
R1335 B.n880 B.n879 71.676
R1336 B.n873 B.n131 71.676
R1337 B.n872 B.n871 71.676
R1338 B.n865 B.n133 71.676
R1339 B.n864 B.n863 71.676
R1340 B.n857 B.n138 71.676
R1341 B.n856 B.n855 71.676
R1342 B.n848 B.n140 71.676
R1343 B.n847 B.n846 71.676
R1344 B.n840 B.n144 71.676
R1345 B.n839 B.n838 71.676
R1346 B.n832 B.n146 71.676
R1347 B.n831 B.n830 71.676
R1348 B.n824 B.n148 71.676
R1349 B.n823 B.n822 71.676
R1350 B.n816 B.n150 71.676
R1351 B.n815 B.n814 71.676
R1352 B.n808 B.n152 71.676
R1353 B.n807 B.n806 71.676
R1354 B.n800 B.n154 71.676
R1355 B.n799 B.n798 71.676
R1356 B.n792 B.n156 71.676
R1357 B.n791 B.n790 71.676
R1358 B.n784 B.n158 71.676
R1359 B.n783 B.n782 71.676
R1360 B.n776 B.n160 71.676
R1361 B.n775 B.n774 71.676
R1362 B.n774 B.n773 71.676
R1363 B.n777 B.n776 71.676
R1364 B.n782 B.n781 71.676
R1365 B.n785 B.n784 71.676
R1366 B.n790 B.n789 71.676
R1367 B.n793 B.n792 71.676
R1368 B.n798 B.n797 71.676
R1369 B.n801 B.n800 71.676
R1370 B.n806 B.n805 71.676
R1371 B.n809 B.n808 71.676
R1372 B.n814 B.n813 71.676
R1373 B.n817 B.n816 71.676
R1374 B.n822 B.n821 71.676
R1375 B.n825 B.n824 71.676
R1376 B.n830 B.n829 71.676
R1377 B.n833 B.n832 71.676
R1378 B.n838 B.n837 71.676
R1379 B.n841 B.n840 71.676
R1380 B.n846 B.n845 71.676
R1381 B.n849 B.n848 71.676
R1382 B.n855 B.n854 71.676
R1383 B.n858 B.n857 71.676
R1384 B.n863 B.n862 71.676
R1385 B.n866 B.n865 71.676
R1386 B.n871 B.n870 71.676
R1387 B.n874 B.n873 71.676
R1388 B.n879 B.n878 71.676
R1389 B.n882 B.n881 71.676
R1390 B.n887 B.n886 71.676
R1391 B.n890 B.n889 71.676
R1392 B.n895 B.n894 71.676
R1393 B.n898 B.n897 71.676
R1394 B.n903 B.n902 71.676
R1395 B.n906 B.n905 71.676
R1396 B.n911 B.n910 71.676
R1397 B.n914 B.n913 71.676
R1398 B.n919 B.n918 71.676
R1399 B.n922 B.n921 71.676
R1400 B.n927 B.n926 71.676
R1401 B.n930 B.n929 71.676
R1402 B.n935 B.n934 71.676
R1403 B.n938 B.n937 71.676
R1404 B.n943 B.n942 71.676
R1405 B.n946 B.n945 71.676
R1406 B.n504 B.n503 71.676
R1407 B.n498 B.n286 71.676
R1408 B.n496 B.n495 71.676
R1409 B.n491 B.n490 71.676
R1410 B.n488 B.n487 71.676
R1411 B.n483 B.n482 71.676
R1412 B.n480 B.n479 71.676
R1413 B.n475 B.n474 71.676
R1414 B.n472 B.n471 71.676
R1415 B.n467 B.n466 71.676
R1416 B.n464 B.n463 71.676
R1417 B.n459 B.n458 71.676
R1418 B.n456 B.n455 71.676
R1419 B.n451 B.n450 71.676
R1420 B.n448 B.n447 71.676
R1421 B.n443 B.n442 71.676
R1422 B.n440 B.n439 71.676
R1423 B.n435 B.n434 71.676
R1424 B.n432 B.n431 71.676
R1425 B.n426 B.n425 71.676
R1426 B.n423 B.n422 71.676
R1427 B.n418 B.n417 71.676
R1428 B.n415 B.n414 71.676
R1429 B.n410 B.n409 71.676
R1430 B.n405 B.n314 71.676
R1431 B.n403 B.n402 71.676
R1432 B.n398 B.n397 71.676
R1433 B.n395 B.n394 71.676
R1434 B.n390 B.n389 71.676
R1435 B.n387 B.n386 71.676
R1436 B.n382 B.n381 71.676
R1437 B.n379 B.n378 71.676
R1438 B.n374 B.n373 71.676
R1439 B.n371 B.n370 71.676
R1440 B.n366 B.n365 71.676
R1441 B.n363 B.n362 71.676
R1442 B.n358 B.n357 71.676
R1443 B.n355 B.n354 71.676
R1444 B.n350 B.n349 71.676
R1445 B.n347 B.n346 71.676
R1446 B.n342 B.n341 71.676
R1447 B.n339 B.n338 71.676
R1448 B.n334 B.n333 71.676
R1449 B.n312 B.n311 71.1763
R1450 B.n306 B.n305 71.1763
R1451 B.n135 B.n134 71.1763
R1452 B.n142 B.n141 71.1763
R1453 B.n313 B.n312 59.5399
R1454 B.n429 B.n306 59.5399
R1455 B.n136 B.n135 59.5399
R1456 B.n851 B.n142 59.5399
R1457 B.n509 B.n279 45.652
R1458 B.n515 B.n279 45.652
R1459 B.n515 B.n275 45.652
R1460 B.n521 B.n275 45.652
R1461 B.n521 B.n271 45.652
R1462 B.n527 B.n271 45.652
R1463 B.n527 B.n267 45.652
R1464 B.n533 B.n267 45.652
R1465 B.n539 B.n263 45.652
R1466 B.n539 B.n259 45.652
R1467 B.n545 B.n259 45.652
R1468 B.n545 B.n255 45.652
R1469 B.n551 B.n255 45.652
R1470 B.n551 B.n251 45.652
R1471 B.n557 B.n251 45.652
R1472 B.n557 B.n247 45.652
R1473 B.n563 B.n247 45.652
R1474 B.n563 B.n243 45.652
R1475 B.n569 B.n243 45.652
R1476 B.n569 B.n239 45.652
R1477 B.n575 B.n239 45.652
R1478 B.n581 B.n235 45.652
R1479 B.n581 B.n231 45.652
R1480 B.n587 B.n231 45.652
R1481 B.n587 B.n227 45.652
R1482 B.n593 B.n227 45.652
R1483 B.n593 B.n223 45.652
R1484 B.n599 B.n223 45.652
R1485 B.n599 B.n218 45.652
R1486 B.n605 B.n218 45.652
R1487 B.n605 B.n219 45.652
R1488 B.n611 B.n211 45.652
R1489 B.n617 B.n211 45.652
R1490 B.n617 B.n207 45.652
R1491 B.n623 B.n207 45.652
R1492 B.n623 B.n203 45.652
R1493 B.n629 B.n203 45.652
R1494 B.n629 B.n199 45.652
R1495 B.n635 B.n199 45.652
R1496 B.n635 B.n195 45.652
R1497 B.n641 B.n195 45.652
R1498 B.n647 B.n191 45.652
R1499 B.n647 B.n187 45.652
R1500 B.n653 B.n187 45.652
R1501 B.n653 B.n183 45.652
R1502 B.n659 B.n183 45.652
R1503 B.n659 B.n179 45.652
R1504 B.n665 B.n179 45.652
R1505 B.n665 B.n175 45.652
R1506 B.n671 B.n175 45.652
R1507 B.n671 B.t4 45.652
R1508 B.n677 B.t4 45.652
R1509 B.n677 B.n168 45.652
R1510 B.n684 B.n168 45.652
R1511 B.n684 B.n164 45.652
R1512 B.n690 B.n164 45.652
R1513 B.n690 B.n4 45.652
R1514 B.n1073 B.n4 45.652
R1515 B.n1073 B.n1072 45.652
R1516 B.n1072 B.n1071 45.652
R1517 B.n1071 B.n8 45.652
R1518 B.n1065 B.n8 45.652
R1519 B.n1065 B.n1064 45.652
R1520 B.n1064 B.n1063 45.652
R1521 B.n1063 B.t0 45.652
R1522 B.n1057 B.t0 45.652
R1523 B.n1057 B.n1056 45.652
R1524 B.n1056 B.n1055 45.652
R1525 B.n1055 B.n21 45.652
R1526 B.n1049 B.n21 45.652
R1527 B.n1049 B.n1048 45.652
R1528 B.n1048 B.n1047 45.652
R1529 B.n1047 B.n28 45.652
R1530 B.n1041 B.n28 45.652
R1531 B.n1041 B.n1040 45.652
R1532 B.n1039 B.n35 45.652
R1533 B.n1033 B.n35 45.652
R1534 B.n1033 B.n1032 45.652
R1535 B.n1032 B.n1031 45.652
R1536 B.n1031 B.n42 45.652
R1537 B.n1025 B.n42 45.652
R1538 B.n1025 B.n1024 45.652
R1539 B.n1024 B.n1023 45.652
R1540 B.n1023 B.n49 45.652
R1541 B.n1017 B.n49 45.652
R1542 B.n1016 B.n1015 45.652
R1543 B.n1015 B.n56 45.652
R1544 B.n1009 B.n56 45.652
R1545 B.n1009 B.n1008 45.652
R1546 B.n1008 B.n1007 45.652
R1547 B.n1007 B.n63 45.652
R1548 B.n1001 B.n63 45.652
R1549 B.n1001 B.n1000 45.652
R1550 B.n1000 B.n999 45.652
R1551 B.n999 B.n70 45.652
R1552 B.n993 B.n992 45.652
R1553 B.n992 B.n991 45.652
R1554 B.n991 B.n77 45.652
R1555 B.n985 B.n77 45.652
R1556 B.n985 B.n984 45.652
R1557 B.n984 B.n983 45.652
R1558 B.n983 B.n84 45.652
R1559 B.n977 B.n84 45.652
R1560 B.n977 B.n976 45.652
R1561 B.n976 B.n975 45.652
R1562 B.n975 B.n91 45.652
R1563 B.n969 B.n91 45.652
R1564 B.n969 B.n968 45.652
R1565 B.n967 B.n98 45.652
R1566 B.n961 B.n98 45.652
R1567 B.n961 B.n960 45.652
R1568 B.n960 B.n959 45.652
R1569 B.n959 B.n105 45.652
R1570 B.n953 B.n105 45.652
R1571 B.n953 B.n952 45.652
R1572 B.n952 B.n951 45.652
R1573 B.t6 B.n191 36.2532
R1574 B.n1040 B.t2 36.2532
R1575 B.n949 B.n948 31.0639
R1576 B.n772 B.n771 31.0639
R1577 B.n511 B.n281 31.0639
R1578 B.n507 B.n506 31.0639
R1579 B.n533 B.t13 28.197
R1580 B.n575 B.t1 28.197
R1581 B.n993 B.t3 28.197
R1582 B.t9 B.n967 28.197
R1583 B.n611 B.t5 26.8543
R1584 B.n1017 B.t7 26.8543
R1585 B.n219 B.t5 18.7982
R1586 B.t7 B.n1016 18.7982
R1587 B B.n1075 18.0485
R1588 B.t13 B.n263 17.4555
R1589 B.t1 B.n235 17.4555
R1590 B.t3 B.n70 17.4555
R1591 B.n968 B.t9 17.4555
R1592 B.n948 B.n947 10.6151
R1593 B.n947 B.n114 10.6151
R1594 B.n941 B.n114 10.6151
R1595 B.n941 B.n940 10.6151
R1596 B.n940 B.n939 10.6151
R1597 B.n939 B.n116 10.6151
R1598 B.n933 B.n116 10.6151
R1599 B.n933 B.n932 10.6151
R1600 B.n932 B.n931 10.6151
R1601 B.n931 B.n118 10.6151
R1602 B.n925 B.n118 10.6151
R1603 B.n925 B.n924 10.6151
R1604 B.n924 B.n923 10.6151
R1605 B.n923 B.n120 10.6151
R1606 B.n917 B.n120 10.6151
R1607 B.n917 B.n916 10.6151
R1608 B.n916 B.n915 10.6151
R1609 B.n915 B.n122 10.6151
R1610 B.n909 B.n122 10.6151
R1611 B.n909 B.n908 10.6151
R1612 B.n908 B.n907 10.6151
R1613 B.n907 B.n124 10.6151
R1614 B.n901 B.n124 10.6151
R1615 B.n901 B.n900 10.6151
R1616 B.n900 B.n899 10.6151
R1617 B.n899 B.n126 10.6151
R1618 B.n893 B.n126 10.6151
R1619 B.n893 B.n892 10.6151
R1620 B.n892 B.n891 10.6151
R1621 B.n891 B.n128 10.6151
R1622 B.n885 B.n128 10.6151
R1623 B.n885 B.n884 10.6151
R1624 B.n884 B.n883 10.6151
R1625 B.n883 B.n130 10.6151
R1626 B.n877 B.n130 10.6151
R1627 B.n877 B.n876 10.6151
R1628 B.n876 B.n875 10.6151
R1629 B.n875 B.n132 10.6151
R1630 B.n869 B.n868 10.6151
R1631 B.n868 B.n867 10.6151
R1632 B.n867 B.n137 10.6151
R1633 B.n861 B.n137 10.6151
R1634 B.n861 B.n860 10.6151
R1635 B.n860 B.n859 10.6151
R1636 B.n859 B.n139 10.6151
R1637 B.n853 B.n139 10.6151
R1638 B.n853 B.n852 10.6151
R1639 B.n850 B.n143 10.6151
R1640 B.n844 B.n143 10.6151
R1641 B.n844 B.n843 10.6151
R1642 B.n843 B.n842 10.6151
R1643 B.n842 B.n145 10.6151
R1644 B.n836 B.n145 10.6151
R1645 B.n836 B.n835 10.6151
R1646 B.n835 B.n834 10.6151
R1647 B.n834 B.n147 10.6151
R1648 B.n828 B.n147 10.6151
R1649 B.n828 B.n827 10.6151
R1650 B.n827 B.n826 10.6151
R1651 B.n826 B.n149 10.6151
R1652 B.n820 B.n149 10.6151
R1653 B.n820 B.n819 10.6151
R1654 B.n819 B.n818 10.6151
R1655 B.n818 B.n151 10.6151
R1656 B.n812 B.n151 10.6151
R1657 B.n812 B.n811 10.6151
R1658 B.n811 B.n810 10.6151
R1659 B.n810 B.n153 10.6151
R1660 B.n804 B.n153 10.6151
R1661 B.n804 B.n803 10.6151
R1662 B.n803 B.n802 10.6151
R1663 B.n802 B.n155 10.6151
R1664 B.n796 B.n155 10.6151
R1665 B.n796 B.n795 10.6151
R1666 B.n795 B.n794 10.6151
R1667 B.n794 B.n157 10.6151
R1668 B.n788 B.n157 10.6151
R1669 B.n788 B.n787 10.6151
R1670 B.n787 B.n786 10.6151
R1671 B.n786 B.n159 10.6151
R1672 B.n780 B.n159 10.6151
R1673 B.n780 B.n779 10.6151
R1674 B.n779 B.n778 10.6151
R1675 B.n778 B.n161 10.6151
R1676 B.n772 B.n161 10.6151
R1677 B.n512 B.n511 10.6151
R1678 B.n513 B.n512 10.6151
R1679 B.n513 B.n273 10.6151
R1680 B.n523 B.n273 10.6151
R1681 B.n524 B.n523 10.6151
R1682 B.n525 B.n524 10.6151
R1683 B.n525 B.n265 10.6151
R1684 B.n535 B.n265 10.6151
R1685 B.n536 B.n535 10.6151
R1686 B.n537 B.n536 10.6151
R1687 B.n537 B.n257 10.6151
R1688 B.n547 B.n257 10.6151
R1689 B.n548 B.n547 10.6151
R1690 B.n549 B.n548 10.6151
R1691 B.n549 B.n249 10.6151
R1692 B.n559 B.n249 10.6151
R1693 B.n560 B.n559 10.6151
R1694 B.n561 B.n560 10.6151
R1695 B.n561 B.n241 10.6151
R1696 B.n571 B.n241 10.6151
R1697 B.n572 B.n571 10.6151
R1698 B.n573 B.n572 10.6151
R1699 B.n573 B.n233 10.6151
R1700 B.n583 B.n233 10.6151
R1701 B.n584 B.n583 10.6151
R1702 B.n585 B.n584 10.6151
R1703 B.n585 B.n225 10.6151
R1704 B.n595 B.n225 10.6151
R1705 B.n596 B.n595 10.6151
R1706 B.n597 B.n596 10.6151
R1707 B.n597 B.n216 10.6151
R1708 B.n607 B.n216 10.6151
R1709 B.n608 B.n607 10.6151
R1710 B.n609 B.n608 10.6151
R1711 B.n609 B.n209 10.6151
R1712 B.n619 B.n209 10.6151
R1713 B.n620 B.n619 10.6151
R1714 B.n621 B.n620 10.6151
R1715 B.n621 B.n201 10.6151
R1716 B.n631 B.n201 10.6151
R1717 B.n632 B.n631 10.6151
R1718 B.n633 B.n632 10.6151
R1719 B.n633 B.n193 10.6151
R1720 B.n643 B.n193 10.6151
R1721 B.n644 B.n643 10.6151
R1722 B.n645 B.n644 10.6151
R1723 B.n645 B.n185 10.6151
R1724 B.n655 B.n185 10.6151
R1725 B.n656 B.n655 10.6151
R1726 B.n657 B.n656 10.6151
R1727 B.n657 B.n177 10.6151
R1728 B.n667 B.n177 10.6151
R1729 B.n668 B.n667 10.6151
R1730 B.n669 B.n668 10.6151
R1731 B.n669 B.n170 10.6151
R1732 B.n679 B.n170 10.6151
R1733 B.n680 B.n679 10.6151
R1734 B.n682 B.n680 10.6151
R1735 B.n682 B.n681 10.6151
R1736 B.n681 B.n162 10.6151
R1737 B.n693 B.n162 10.6151
R1738 B.n694 B.n693 10.6151
R1739 B.n695 B.n694 10.6151
R1740 B.n696 B.n695 10.6151
R1741 B.n698 B.n696 10.6151
R1742 B.n699 B.n698 10.6151
R1743 B.n700 B.n699 10.6151
R1744 B.n701 B.n700 10.6151
R1745 B.n703 B.n701 10.6151
R1746 B.n704 B.n703 10.6151
R1747 B.n705 B.n704 10.6151
R1748 B.n706 B.n705 10.6151
R1749 B.n708 B.n706 10.6151
R1750 B.n709 B.n708 10.6151
R1751 B.n710 B.n709 10.6151
R1752 B.n711 B.n710 10.6151
R1753 B.n713 B.n711 10.6151
R1754 B.n714 B.n713 10.6151
R1755 B.n715 B.n714 10.6151
R1756 B.n716 B.n715 10.6151
R1757 B.n718 B.n716 10.6151
R1758 B.n719 B.n718 10.6151
R1759 B.n720 B.n719 10.6151
R1760 B.n721 B.n720 10.6151
R1761 B.n723 B.n721 10.6151
R1762 B.n724 B.n723 10.6151
R1763 B.n725 B.n724 10.6151
R1764 B.n726 B.n725 10.6151
R1765 B.n728 B.n726 10.6151
R1766 B.n729 B.n728 10.6151
R1767 B.n730 B.n729 10.6151
R1768 B.n731 B.n730 10.6151
R1769 B.n733 B.n731 10.6151
R1770 B.n734 B.n733 10.6151
R1771 B.n735 B.n734 10.6151
R1772 B.n736 B.n735 10.6151
R1773 B.n738 B.n736 10.6151
R1774 B.n739 B.n738 10.6151
R1775 B.n740 B.n739 10.6151
R1776 B.n741 B.n740 10.6151
R1777 B.n743 B.n741 10.6151
R1778 B.n744 B.n743 10.6151
R1779 B.n745 B.n744 10.6151
R1780 B.n746 B.n745 10.6151
R1781 B.n748 B.n746 10.6151
R1782 B.n749 B.n748 10.6151
R1783 B.n750 B.n749 10.6151
R1784 B.n751 B.n750 10.6151
R1785 B.n753 B.n751 10.6151
R1786 B.n754 B.n753 10.6151
R1787 B.n755 B.n754 10.6151
R1788 B.n756 B.n755 10.6151
R1789 B.n758 B.n756 10.6151
R1790 B.n759 B.n758 10.6151
R1791 B.n760 B.n759 10.6151
R1792 B.n761 B.n760 10.6151
R1793 B.n763 B.n761 10.6151
R1794 B.n764 B.n763 10.6151
R1795 B.n765 B.n764 10.6151
R1796 B.n766 B.n765 10.6151
R1797 B.n768 B.n766 10.6151
R1798 B.n769 B.n768 10.6151
R1799 B.n770 B.n769 10.6151
R1800 B.n771 B.n770 10.6151
R1801 B.n506 B.n505 10.6151
R1802 B.n505 B.n285 10.6151
R1803 B.n500 B.n285 10.6151
R1804 B.n500 B.n499 10.6151
R1805 B.n499 B.n287 10.6151
R1806 B.n494 B.n287 10.6151
R1807 B.n494 B.n493 10.6151
R1808 B.n493 B.n492 10.6151
R1809 B.n492 B.n289 10.6151
R1810 B.n486 B.n289 10.6151
R1811 B.n486 B.n485 10.6151
R1812 B.n485 B.n484 10.6151
R1813 B.n484 B.n291 10.6151
R1814 B.n478 B.n291 10.6151
R1815 B.n478 B.n477 10.6151
R1816 B.n477 B.n476 10.6151
R1817 B.n476 B.n293 10.6151
R1818 B.n470 B.n293 10.6151
R1819 B.n470 B.n469 10.6151
R1820 B.n469 B.n468 10.6151
R1821 B.n468 B.n295 10.6151
R1822 B.n462 B.n295 10.6151
R1823 B.n462 B.n461 10.6151
R1824 B.n461 B.n460 10.6151
R1825 B.n460 B.n297 10.6151
R1826 B.n454 B.n297 10.6151
R1827 B.n454 B.n453 10.6151
R1828 B.n453 B.n452 10.6151
R1829 B.n452 B.n299 10.6151
R1830 B.n446 B.n299 10.6151
R1831 B.n446 B.n445 10.6151
R1832 B.n445 B.n444 10.6151
R1833 B.n444 B.n301 10.6151
R1834 B.n438 B.n301 10.6151
R1835 B.n438 B.n437 10.6151
R1836 B.n437 B.n436 10.6151
R1837 B.n436 B.n303 10.6151
R1838 B.n430 B.n303 10.6151
R1839 B.n428 B.n427 10.6151
R1840 B.n427 B.n307 10.6151
R1841 B.n421 B.n307 10.6151
R1842 B.n421 B.n420 10.6151
R1843 B.n420 B.n419 10.6151
R1844 B.n419 B.n309 10.6151
R1845 B.n413 B.n309 10.6151
R1846 B.n413 B.n412 10.6151
R1847 B.n412 B.n411 10.6151
R1848 B.n407 B.n406 10.6151
R1849 B.n406 B.n315 10.6151
R1850 B.n401 B.n315 10.6151
R1851 B.n401 B.n400 10.6151
R1852 B.n400 B.n399 10.6151
R1853 B.n399 B.n317 10.6151
R1854 B.n393 B.n317 10.6151
R1855 B.n393 B.n392 10.6151
R1856 B.n392 B.n391 10.6151
R1857 B.n391 B.n319 10.6151
R1858 B.n385 B.n319 10.6151
R1859 B.n385 B.n384 10.6151
R1860 B.n384 B.n383 10.6151
R1861 B.n383 B.n321 10.6151
R1862 B.n377 B.n321 10.6151
R1863 B.n377 B.n376 10.6151
R1864 B.n376 B.n375 10.6151
R1865 B.n375 B.n323 10.6151
R1866 B.n369 B.n323 10.6151
R1867 B.n369 B.n368 10.6151
R1868 B.n368 B.n367 10.6151
R1869 B.n367 B.n325 10.6151
R1870 B.n361 B.n325 10.6151
R1871 B.n361 B.n360 10.6151
R1872 B.n360 B.n359 10.6151
R1873 B.n359 B.n327 10.6151
R1874 B.n353 B.n327 10.6151
R1875 B.n353 B.n352 10.6151
R1876 B.n352 B.n351 10.6151
R1877 B.n351 B.n329 10.6151
R1878 B.n345 B.n329 10.6151
R1879 B.n345 B.n344 10.6151
R1880 B.n344 B.n343 10.6151
R1881 B.n343 B.n331 10.6151
R1882 B.n337 B.n331 10.6151
R1883 B.n337 B.n336 10.6151
R1884 B.n336 B.n335 10.6151
R1885 B.n335 B.n281 10.6151
R1886 B.n507 B.n277 10.6151
R1887 B.n517 B.n277 10.6151
R1888 B.n518 B.n517 10.6151
R1889 B.n519 B.n518 10.6151
R1890 B.n519 B.n269 10.6151
R1891 B.n529 B.n269 10.6151
R1892 B.n530 B.n529 10.6151
R1893 B.n531 B.n530 10.6151
R1894 B.n531 B.n261 10.6151
R1895 B.n541 B.n261 10.6151
R1896 B.n542 B.n541 10.6151
R1897 B.n543 B.n542 10.6151
R1898 B.n543 B.n253 10.6151
R1899 B.n553 B.n253 10.6151
R1900 B.n554 B.n553 10.6151
R1901 B.n555 B.n554 10.6151
R1902 B.n555 B.n245 10.6151
R1903 B.n565 B.n245 10.6151
R1904 B.n566 B.n565 10.6151
R1905 B.n567 B.n566 10.6151
R1906 B.n567 B.n237 10.6151
R1907 B.n577 B.n237 10.6151
R1908 B.n578 B.n577 10.6151
R1909 B.n579 B.n578 10.6151
R1910 B.n579 B.n229 10.6151
R1911 B.n589 B.n229 10.6151
R1912 B.n590 B.n589 10.6151
R1913 B.n591 B.n590 10.6151
R1914 B.n591 B.n221 10.6151
R1915 B.n601 B.n221 10.6151
R1916 B.n602 B.n601 10.6151
R1917 B.n603 B.n602 10.6151
R1918 B.n603 B.n213 10.6151
R1919 B.n613 B.n213 10.6151
R1920 B.n614 B.n613 10.6151
R1921 B.n615 B.n614 10.6151
R1922 B.n615 B.n205 10.6151
R1923 B.n625 B.n205 10.6151
R1924 B.n626 B.n625 10.6151
R1925 B.n627 B.n626 10.6151
R1926 B.n627 B.n197 10.6151
R1927 B.n637 B.n197 10.6151
R1928 B.n638 B.n637 10.6151
R1929 B.n639 B.n638 10.6151
R1930 B.n639 B.n189 10.6151
R1931 B.n649 B.n189 10.6151
R1932 B.n650 B.n649 10.6151
R1933 B.n651 B.n650 10.6151
R1934 B.n651 B.n181 10.6151
R1935 B.n661 B.n181 10.6151
R1936 B.n662 B.n661 10.6151
R1937 B.n663 B.n662 10.6151
R1938 B.n663 B.n173 10.6151
R1939 B.n673 B.n173 10.6151
R1940 B.n674 B.n673 10.6151
R1941 B.n675 B.n674 10.6151
R1942 B.n675 B.n166 10.6151
R1943 B.n686 B.n166 10.6151
R1944 B.n687 B.n686 10.6151
R1945 B.n688 B.n687 10.6151
R1946 B.n688 B.n0 10.6151
R1947 B.n1069 B.n1 10.6151
R1948 B.n1069 B.n1068 10.6151
R1949 B.n1068 B.n1067 10.6151
R1950 B.n1067 B.n10 10.6151
R1951 B.n1061 B.n10 10.6151
R1952 B.n1061 B.n1060 10.6151
R1953 B.n1060 B.n1059 10.6151
R1954 B.n1059 B.n16 10.6151
R1955 B.n1053 B.n16 10.6151
R1956 B.n1053 B.n1052 10.6151
R1957 B.n1052 B.n1051 10.6151
R1958 B.n1051 B.n23 10.6151
R1959 B.n1045 B.n23 10.6151
R1960 B.n1045 B.n1044 10.6151
R1961 B.n1044 B.n1043 10.6151
R1962 B.n1043 B.n30 10.6151
R1963 B.n1037 B.n30 10.6151
R1964 B.n1037 B.n1036 10.6151
R1965 B.n1036 B.n1035 10.6151
R1966 B.n1035 B.n37 10.6151
R1967 B.n1029 B.n37 10.6151
R1968 B.n1029 B.n1028 10.6151
R1969 B.n1028 B.n1027 10.6151
R1970 B.n1027 B.n44 10.6151
R1971 B.n1021 B.n44 10.6151
R1972 B.n1021 B.n1020 10.6151
R1973 B.n1020 B.n1019 10.6151
R1974 B.n1019 B.n51 10.6151
R1975 B.n1013 B.n51 10.6151
R1976 B.n1013 B.n1012 10.6151
R1977 B.n1012 B.n1011 10.6151
R1978 B.n1011 B.n58 10.6151
R1979 B.n1005 B.n58 10.6151
R1980 B.n1005 B.n1004 10.6151
R1981 B.n1004 B.n1003 10.6151
R1982 B.n1003 B.n65 10.6151
R1983 B.n997 B.n65 10.6151
R1984 B.n997 B.n996 10.6151
R1985 B.n996 B.n995 10.6151
R1986 B.n995 B.n72 10.6151
R1987 B.n989 B.n72 10.6151
R1988 B.n989 B.n988 10.6151
R1989 B.n988 B.n987 10.6151
R1990 B.n987 B.n79 10.6151
R1991 B.n981 B.n79 10.6151
R1992 B.n981 B.n980 10.6151
R1993 B.n980 B.n979 10.6151
R1994 B.n979 B.n86 10.6151
R1995 B.n973 B.n86 10.6151
R1996 B.n973 B.n972 10.6151
R1997 B.n972 B.n971 10.6151
R1998 B.n971 B.n93 10.6151
R1999 B.n965 B.n93 10.6151
R2000 B.n965 B.n964 10.6151
R2001 B.n964 B.n963 10.6151
R2002 B.n963 B.n100 10.6151
R2003 B.n957 B.n100 10.6151
R2004 B.n957 B.n956 10.6151
R2005 B.n956 B.n955 10.6151
R2006 B.n955 B.n107 10.6151
R2007 B.n949 B.n107 10.6151
R2008 B.n641 B.t6 9.39934
R2009 B.t2 B.n1039 9.39934
R2010 B.n136 B.n132 9.36635
R2011 B.n851 B.n850 9.36635
R2012 B.n430 B.n429 9.36635
R2013 B.n407 B.n313 9.36635
R2014 B.n1075 B.n0 2.81026
R2015 B.n1075 B.n1 2.81026
R2016 B.n869 B.n136 1.24928
R2017 B.n852 B.n851 1.24928
R2018 B.n429 B.n428 1.24928
R2019 B.n411 B.n313 1.24928
R2020 VP.n24 VP.n21 161.3
R2021 VP.n26 VP.n25 161.3
R2022 VP.n27 VP.n20 161.3
R2023 VP.n29 VP.n28 161.3
R2024 VP.n30 VP.n19 161.3
R2025 VP.n32 VP.n31 161.3
R2026 VP.n33 VP.n18 161.3
R2027 VP.n35 VP.n34 161.3
R2028 VP.n37 VP.n36 161.3
R2029 VP.n38 VP.n16 161.3
R2030 VP.n40 VP.n39 161.3
R2031 VP.n41 VP.n15 161.3
R2032 VP.n43 VP.n42 161.3
R2033 VP.n44 VP.n14 161.3
R2034 VP.n46 VP.n45 161.3
R2035 VP.n83 VP.n82 161.3
R2036 VP.n81 VP.n1 161.3
R2037 VP.n80 VP.n79 161.3
R2038 VP.n78 VP.n2 161.3
R2039 VP.n77 VP.n76 161.3
R2040 VP.n75 VP.n3 161.3
R2041 VP.n74 VP.n73 161.3
R2042 VP.n72 VP.n71 161.3
R2043 VP.n70 VP.n5 161.3
R2044 VP.n69 VP.n68 161.3
R2045 VP.n67 VP.n6 161.3
R2046 VP.n66 VP.n65 161.3
R2047 VP.n64 VP.n7 161.3
R2048 VP.n63 VP.n62 161.3
R2049 VP.n61 VP.n8 161.3
R2050 VP.n60 VP.n59 161.3
R2051 VP.n57 VP.n9 161.3
R2052 VP.n56 VP.n55 161.3
R2053 VP.n54 VP.n10 161.3
R2054 VP.n53 VP.n52 161.3
R2055 VP.n51 VP.n11 161.3
R2056 VP.n50 VP.n49 161.3
R2057 VP.n23 VP.t7 112.716
R2058 VP.n12 VP.t4 80.1655
R2059 VP.n58 VP.t1 80.1655
R2060 VP.n4 VP.t6 80.1655
R2061 VP.n0 VP.t3 80.1655
R2062 VP.n13 VP.t0 80.1655
R2063 VP.n17 VP.t2 80.1655
R2064 VP.n22 VP.t5 80.1655
R2065 VP.n48 VP.n12 77.5892
R2066 VP.n84 VP.n0 77.5892
R2067 VP.n47 VP.n13 77.5892
R2068 VP.n23 VP.n22 70.4248
R2069 VP.n65 VP.n6 56.5193
R2070 VP.n28 VP.n19 56.5193
R2071 VP.n48 VP.n47 53.7721
R2072 VP.n56 VP.n10 48.2635
R2073 VP.n76 VP.n2 48.2635
R2074 VP.n39 VP.n15 48.2635
R2075 VP.n52 VP.n10 32.7233
R2076 VP.n80 VP.n2 32.7233
R2077 VP.n43 VP.n15 32.7233
R2078 VP.n51 VP.n50 24.4675
R2079 VP.n52 VP.n51 24.4675
R2080 VP.n57 VP.n56 24.4675
R2081 VP.n59 VP.n57 24.4675
R2082 VP.n63 VP.n8 24.4675
R2083 VP.n64 VP.n63 24.4675
R2084 VP.n65 VP.n64 24.4675
R2085 VP.n69 VP.n6 24.4675
R2086 VP.n70 VP.n69 24.4675
R2087 VP.n71 VP.n70 24.4675
R2088 VP.n75 VP.n74 24.4675
R2089 VP.n76 VP.n75 24.4675
R2090 VP.n81 VP.n80 24.4675
R2091 VP.n82 VP.n81 24.4675
R2092 VP.n44 VP.n43 24.4675
R2093 VP.n45 VP.n44 24.4675
R2094 VP.n32 VP.n19 24.4675
R2095 VP.n33 VP.n32 24.4675
R2096 VP.n34 VP.n33 24.4675
R2097 VP.n38 VP.n37 24.4675
R2098 VP.n39 VP.n38 24.4675
R2099 VP.n26 VP.n21 24.4675
R2100 VP.n27 VP.n26 24.4675
R2101 VP.n28 VP.n27 24.4675
R2102 VP.n59 VP.n58 20.3081
R2103 VP.n74 VP.n4 20.3081
R2104 VP.n37 VP.n17 20.3081
R2105 VP.n50 VP.n12 12.4787
R2106 VP.n82 VP.n0 12.4787
R2107 VP.n45 VP.n13 12.4787
R2108 VP.n24 VP.n23 4.27758
R2109 VP.n58 VP.n8 4.15989
R2110 VP.n71 VP.n4 4.15989
R2111 VP.n34 VP.n17 4.15989
R2112 VP.n22 VP.n21 4.15989
R2113 VP.n47 VP.n46 0.354971
R2114 VP.n49 VP.n48 0.354971
R2115 VP.n84 VP.n83 0.354971
R2116 VP VP.n84 0.26696
R2117 VP.n25 VP.n24 0.189894
R2118 VP.n25 VP.n20 0.189894
R2119 VP.n29 VP.n20 0.189894
R2120 VP.n30 VP.n29 0.189894
R2121 VP.n31 VP.n30 0.189894
R2122 VP.n31 VP.n18 0.189894
R2123 VP.n35 VP.n18 0.189894
R2124 VP.n36 VP.n35 0.189894
R2125 VP.n36 VP.n16 0.189894
R2126 VP.n40 VP.n16 0.189894
R2127 VP.n41 VP.n40 0.189894
R2128 VP.n42 VP.n41 0.189894
R2129 VP.n42 VP.n14 0.189894
R2130 VP.n46 VP.n14 0.189894
R2131 VP.n49 VP.n11 0.189894
R2132 VP.n53 VP.n11 0.189894
R2133 VP.n54 VP.n53 0.189894
R2134 VP.n55 VP.n54 0.189894
R2135 VP.n55 VP.n9 0.189894
R2136 VP.n60 VP.n9 0.189894
R2137 VP.n61 VP.n60 0.189894
R2138 VP.n62 VP.n61 0.189894
R2139 VP.n62 VP.n7 0.189894
R2140 VP.n66 VP.n7 0.189894
R2141 VP.n67 VP.n66 0.189894
R2142 VP.n68 VP.n67 0.189894
R2143 VP.n68 VP.n5 0.189894
R2144 VP.n72 VP.n5 0.189894
R2145 VP.n73 VP.n72 0.189894
R2146 VP.n73 VP.n3 0.189894
R2147 VP.n77 VP.n3 0.189894
R2148 VP.n78 VP.n77 0.189894
R2149 VP.n79 VP.n78 0.189894
R2150 VP.n79 VP.n1 0.189894
R2151 VP.n83 VP.n1 0.189894
R2152 VDD1 VDD1.n0 65.2068
R2153 VDD1.n3 VDD1.n2 65.093
R2154 VDD1.n3 VDD1.n1 65.093
R2155 VDD1.n5 VDD1.n4 63.5665
R2156 VDD1.n5 VDD1.n3 48.113
R2157 VDD1.n4 VDD1.t5 1.78268
R2158 VDD1.n4 VDD1.t7 1.78268
R2159 VDD1.n0 VDD1.t0 1.78268
R2160 VDD1.n0 VDD1.t2 1.78268
R2161 VDD1.n2 VDD1.t1 1.78268
R2162 VDD1.n2 VDD1.t4 1.78268
R2163 VDD1.n1 VDD1.t3 1.78268
R2164 VDD1.n1 VDD1.t6 1.78268
R2165 VDD1 VDD1.n5 1.52421
C0 VDD1 VN 0.152879f
C1 VP VN 8.40473f
C2 VTAIL VN 9.126901f
C3 VDD2 VN 8.44736f
C4 VP VDD1 8.890941f
C5 VTAIL VDD1 8.08239f
C6 VP VTAIL 9.14101f
C7 VDD2 VDD1 2.15897f
C8 VP VDD2 0.598228f
C9 VDD2 VTAIL 8.141769f
C10 VDD2 B 6.082298f
C11 VDD1 B 6.606905f
C12 VTAIL B 10.454473f
C13 VN B 18.290218f
C14 VP B 16.94458f
C15 VDD1.t0 B 0.243602f
C16 VDD1.t2 B 0.243602f
C17 VDD1.n0 B 2.17837f
C18 VDD1.t3 B 0.243602f
C19 VDD1.t6 B 0.243602f
C20 VDD1.n1 B 2.17701f
C21 VDD1.t1 B 0.243602f
C22 VDD1.t4 B 0.243602f
C23 VDD1.n2 B 2.17701f
C24 VDD1.n3 B 4.10611f
C25 VDD1.t5 B 0.243602f
C26 VDD1.t7 B 0.243602f
C27 VDD1.n4 B 2.16157f
C28 VDD1.n5 B 3.51744f
C29 VP.t3 B 1.95645f
C30 VP.n0 B 0.764665f
C31 VP.n1 B 0.019395f
C32 VP.n2 B 0.017335f
C33 VP.n3 B 0.019395f
C34 VP.t6 B 1.95645f
C35 VP.n4 B 0.690168f
C36 VP.n5 B 0.019395f
C37 VP.n6 B 0.028314f
C38 VP.n7 B 0.019395f
C39 VP.n8 B 0.021335f
C40 VP.n9 B 0.019395f
C41 VP.n10 B 0.017335f
C42 VP.n11 B 0.019395f
C43 VP.t4 B 1.95645f
C44 VP.n12 B 0.764665f
C45 VP.t0 B 1.95645f
C46 VP.n13 B 0.764665f
C47 VP.n14 B 0.019395f
C48 VP.n15 B 0.017335f
C49 VP.n16 B 0.019395f
C50 VP.t2 B 1.95645f
C51 VP.n17 B 0.690168f
C52 VP.n18 B 0.019395f
C53 VP.n19 B 0.028314f
C54 VP.n20 B 0.019395f
C55 VP.n21 B 0.021335f
C56 VP.t7 B 2.19561f
C57 VP.t5 B 1.95645f
C58 VP.n22 B 0.750221f
C59 VP.n23 B 0.716247f
C60 VP.n24 B 0.229669f
C61 VP.n25 B 0.019395f
C62 VP.n26 B 0.036148f
C63 VP.n27 B 0.036148f
C64 VP.n28 B 0.028314f
C65 VP.n29 B 0.019395f
C66 VP.n30 B 0.019395f
C67 VP.n31 B 0.019395f
C68 VP.n32 B 0.036148f
C69 VP.n33 B 0.036148f
C70 VP.n34 B 0.021335f
C71 VP.n35 B 0.019395f
C72 VP.n36 B 0.019395f
C73 VP.n37 B 0.033113f
C74 VP.n38 B 0.036148f
C75 VP.n39 B 0.036323f
C76 VP.n40 B 0.019395f
C77 VP.n41 B 0.019395f
C78 VP.n42 B 0.019395f
C79 VP.n43 B 0.039118f
C80 VP.n44 B 0.036148f
C81 VP.n45 B 0.027402f
C82 VP.n46 B 0.031304f
C83 VP.n47 B 1.22466f
C84 VP.n48 B 1.23762f
C85 VP.n49 B 0.031304f
C86 VP.n50 B 0.027402f
C87 VP.n51 B 0.036148f
C88 VP.n52 B 0.039118f
C89 VP.n53 B 0.019395f
C90 VP.n54 B 0.019395f
C91 VP.n55 B 0.019395f
C92 VP.n56 B 0.036323f
C93 VP.n57 B 0.036148f
C94 VP.t1 B 1.95645f
C95 VP.n58 B 0.690168f
C96 VP.n59 B 0.033113f
C97 VP.n60 B 0.019395f
C98 VP.n61 B 0.019395f
C99 VP.n62 B 0.019395f
C100 VP.n63 B 0.036148f
C101 VP.n64 B 0.036148f
C102 VP.n65 B 0.028314f
C103 VP.n66 B 0.019395f
C104 VP.n67 B 0.019395f
C105 VP.n68 B 0.019395f
C106 VP.n69 B 0.036148f
C107 VP.n70 B 0.036148f
C108 VP.n71 B 0.021335f
C109 VP.n72 B 0.019395f
C110 VP.n73 B 0.019395f
C111 VP.n74 B 0.033113f
C112 VP.n75 B 0.036148f
C113 VP.n76 B 0.036323f
C114 VP.n77 B 0.019395f
C115 VP.n78 B 0.019395f
C116 VP.n79 B 0.019395f
C117 VP.n80 B 0.039118f
C118 VP.n81 B 0.036148f
C119 VP.n82 B 0.027402f
C120 VP.n83 B 0.031304f
C121 VP.n84 B 0.048919f
C122 VTAIL.t8 B 0.18126f
C123 VTAIL.t15 B 0.18126f
C124 VTAIL.n0 B 1.54972f
C125 VTAIL.n1 B 0.413809f
C126 VTAIL.t11 B 1.97585f
C127 VTAIL.n2 B 0.509409f
C128 VTAIL.t4 B 1.97585f
C129 VTAIL.n3 B 0.509409f
C130 VTAIL.t5 B 0.18126f
C131 VTAIL.t6 B 0.18126f
C132 VTAIL.n4 B 1.54972f
C133 VTAIL.n5 B 0.620411f
C134 VTAIL.t1 B 1.97585f
C135 VTAIL.n6 B 1.60623f
C136 VTAIL.t14 B 1.97586f
C137 VTAIL.n7 B 1.60622f
C138 VTAIL.t9 B 0.18126f
C139 VTAIL.t12 B 0.18126f
C140 VTAIL.n8 B 1.54973f
C141 VTAIL.n9 B 0.620406f
C142 VTAIL.t10 B 1.97586f
C143 VTAIL.n10 B 0.509397f
C144 VTAIL.t0 B 1.97586f
C145 VTAIL.n11 B 0.509397f
C146 VTAIL.t2 B 0.18126f
C147 VTAIL.t7 B 0.18126f
C148 VTAIL.n12 B 1.54973f
C149 VTAIL.n13 B 0.620406f
C150 VTAIL.t3 B 1.97585f
C151 VTAIL.n14 B 1.60623f
C152 VTAIL.t13 B 1.97585f
C153 VTAIL.n15 B 1.60236f
C154 VDD2.t0 B 0.238531f
C155 VDD2.t1 B 0.238531f
C156 VDD2.n0 B 2.13169f
C157 VDD2.t5 B 0.238531f
C158 VDD2.t6 B 0.238531f
C159 VDD2.n1 B 2.13169f
C160 VDD2.n2 B 3.96444f
C161 VDD2.t7 B 0.238531f
C162 VDD2.t3 B 0.238531f
C163 VDD2.n3 B 2.11659f
C164 VDD2.n4 B 3.41025f
C165 VDD2.t2 B 0.238531f
C166 VDD2.t4 B 0.238531f
C167 VDD2.n5 B 2.13165f
C168 VN.t2 B 1.91742f
C169 VN.n0 B 0.749409f
C170 VN.n1 B 0.019008f
C171 VN.n2 B 0.016989f
C172 VN.n3 B 0.019008f
C173 VN.t0 B 1.91742f
C174 VN.n4 B 0.676398f
C175 VN.n5 B 0.019008f
C176 VN.n6 B 0.027749f
C177 VN.n7 B 0.019008f
C178 VN.n8 B 0.020909f
C179 VN.t7 B 1.91742f
C180 VN.n9 B 0.735253f
C181 VN.t4 B 2.1518f
C182 VN.n10 B 0.701956f
C183 VN.n11 B 0.225086f
C184 VN.n12 B 0.019008f
C185 VN.n13 B 0.035427f
C186 VN.n14 B 0.035427f
C187 VN.n15 B 0.027749f
C188 VN.n16 B 0.019008f
C189 VN.n17 B 0.019008f
C190 VN.n18 B 0.019008f
C191 VN.n19 B 0.035427f
C192 VN.n20 B 0.035427f
C193 VN.n21 B 0.020909f
C194 VN.n22 B 0.019008f
C195 VN.n23 B 0.019008f
C196 VN.n24 B 0.032453f
C197 VN.n25 B 0.035427f
C198 VN.n26 B 0.035598f
C199 VN.n27 B 0.019008f
C200 VN.n28 B 0.019008f
C201 VN.n29 B 0.019008f
C202 VN.n30 B 0.038338f
C203 VN.n31 B 0.035427f
C204 VN.n32 B 0.026856f
C205 VN.n33 B 0.030679f
C206 VN.n34 B 0.047943f
C207 VN.t1 B 1.91742f
C208 VN.n35 B 0.749409f
C209 VN.n36 B 0.019008f
C210 VN.n37 B 0.016989f
C211 VN.n38 B 0.019008f
C212 VN.t6 B 1.91742f
C213 VN.n39 B 0.676398f
C214 VN.n40 B 0.019008f
C215 VN.n41 B 0.027749f
C216 VN.n42 B 0.019008f
C217 VN.n43 B 0.020909f
C218 VN.t5 B 2.1518f
C219 VN.t3 B 1.91742f
C220 VN.n44 B 0.735253f
C221 VN.n45 B 0.701956f
C222 VN.n46 B 0.225086f
C223 VN.n47 B 0.019008f
C224 VN.n48 B 0.035427f
C225 VN.n49 B 0.035427f
C226 VN.n50 B 0.027749f
C227 VN.n51 B 0.019008f
C228 VN.n52 B 0.019008f
C229 VN.n53 B 0.019008f
C230 VN.n54 B 0.035427f
C231 VN.n55 B 0.035427f
C232 VN.n56 B 0.020909f
C233 VN.n57 B 0.019008f
C234 VN.n58 B 0.019008f
C235 VN.n59 B 0.032453f
C236 VN.n60 B 0.035427f
C237 VN.n61 B 0.035598f
C238 VN.n62 B 0.019008f
C239 VN.n63 B 0.019008f
C240 VN.n64 B 0.019008f
C241 VN.n65 B 0.038338f
C242 VN.n66 B 0.035427f
C243 VN.n67 B 0.026856f
C244 VN.n68 B 0.030679f
C245 VN.n69 B 1.20781f
.ends

