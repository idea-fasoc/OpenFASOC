* NGSPICE file created from diff_pair_sample_0902.ext - technology: sky130A

.subckt diff_pair_sample_0902 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.17 as=1.1076 ps=6.46 w=2.84 l=2.78
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0 ps=0 w=2.84 l=2.78
X2 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0.4686 ps=3.17 w=2.84 l=2.78
X3 VDD1.t2 VP.t1 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.17 as=1.1076 ps=6.46 w=2.84 l=2.78
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0 ps=0 w=2.84 l=2.78
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0 ps=0 w=2.84 l=2.78
X6 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.17 as=1.1076 ps=6.46 w=2.84 l=2.78
X7 VTAIL.t1 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0.4686 ps=3.17 w=2.84 l=2.78
X8 VDD2.t0 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.17 as=1.1076 ps=6.46 w=2.84 l=2.78
X9 VTAIL.t6 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0.4686 ps=3.17 w=2.84 l=2.78
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0 ps=0 w=2.84 l=2.78
X11 VTAIL.t5 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1076 pd=6.46 as=0.4686 ps=3.17 w=2.84 l=2.78
R0 VP.n16 VP.n0 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n13 VP.n1 161.3
R3 VP.n12 VP.n11 161.3
R4 VP.n10 VP.n2 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n3 161.3
R7 VP.n6 VP.n5 108.204
R8 VP.n18 VP.n17 108.204
R9 VP.n4 VP.t2 59.4693
R10 VP.n4 VP.t0 58.5833
R11 VP.n6 VP.n4 43.409
R12 VP.n11 VP.n10 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n5 VP.t3 24.6206
R15 VP.n17 VP.t1 24.6206
R16 VP.n9 VP.n3 24.5923
R17 VP.n10 VP.n9 24.5923
R18 VP.n15 VP.n1 24.5923
R19 VP.n16 VP.n15 24.5923
R20 VP.n5 VP.n3 2.7056
R21 VP.n17 VP.n16 2.7056
R22 VP.n7 VP.n6 0.278335
R23 VP.n18 VP.n0 0.278335
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153485
R31 VTAIL.n5 VTAIL.t6 72.6731
R32 VTAIL.n4 VTAIL.t0 72.6731
R33 VTAIL.n3 VTAIL.t1 72.6731
R34 VTAIL.n7 VTAIL.t2 72.6729
R35 VTAIL.n0 VTAIL.t3 72.6729
R36 VTAIL.n1 VTAIL.t4 72.6729
R37 VTAIL.n2 VTAIL.t5 72.6729
R38 VTAIL.n6 VTAIL.t7 72.6729
R39 VTAIL.n7 VTAIL.n6 17.4962
R40 VTAIL.n3 VTAIL.n2 17.4962
R41 VTAIL.n4 VTAIL.n3 2.68153
R42 VTAIL.n6 VTAIL.n5 2.68153
R43 VTAIL.n2 VTAIL.n1 2.68153
R44 VTAIL VTAIL.n0 1.39921
R45 VTAIL VTAIL.n7 1.28283
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 VDD1 VDD1.n1 117.111
R49 VDD1 VDD1.n0 82.4382
R50 VDD1.n0 VDD1.t1 6.97233
R51 VDD1.n0 VDD1.t3 6.97233
R52 VDD1.n1 VDD1.t0 6.97233
R53 VDD1.n1 VDD1.t2 6.97233
R54 B.n489 B.n488 585
R55 B.n490 B.n489 585
R56 B.n165 B.n87 585
R57 B.n164 B.n163 585
R58 B.n162 B.n161 585
R59 B.n160 B.n159 585
R60 B.n158 B.n157 585
R61 B.n156 B.n155 585
R62 B.n154 B.n153 585
R63 B.n152 B.n151 585
R64 B.n150 B.n149 585
R65 B.n148 B.n147 585
R66 B.n146 B.n145 585
R67 B.n144 B.n143 585
R68 B.n142 B.n141 585
R69 B.n140 B.n139 585
R70 B.n138 B.n137 585
R71 B.n136 B.n135 585
R72 B.n134 B.n133 585
R73 B.n132 B.n131 585
R74 B.n130 B.n129 585
R75 B.n128 B.n127 585
R76 B.n126 B.n125 585
R77 B.n124 B.n123 585
R78 B.n122 B.n121 585
R79 B.n119 B.n118 585
R80 B.n117 B.n116 585
R81 B.n115 B.n114 585
R82 B.n113 B.n112 585
R83 B.n111 B.n110 585
R84 B.n109 B.n108 585
R85 B.n107 B.n106 585
R86 B.n105 B.n104 585
R87 B.n103 B.n102 585
R88 B.n101 B.n100 585
R89 B.n99 B.n98 585
R90 B.n97 B.n96 585
R91 B.n95 B.n94 585
R92 B.n68 B.n67 585
R93 B.n493 B.n492 585
R94 B.n487 B.n88 585
R95 B.n88 B.n65 585
R96 B.n486 B.n64 585
R97 B.n497 B.n64 585
R98 B.n485 B.n63 585
R99 B.n498 B.n63 585
R100 B.n484 B.n62 585
R101 B.n499 B.n62 585
R102 B.n483 B.n482 585
R103 B.n482 B.n58 585
R104 B.n481 B.n57 585
R105 B.n505 B.n57 585
R106 B.n480 B.n56 585
R107 B.n506 B.n56 585
R108 B.n479 B.n55 585
R109 B.n507 B.n55 585
R110 B.n478 B.n477 585
R111 B.n477 B.n51 585
R112 B.n476 B.n50 585
R113 B.n513 B.n50 585
R114 B.n475 B.n49 585
R115 B.n514 B.n49 585
R116 B.n474 B.n48 585
R117 B.n515 B.n48 585
R118 B.n473 B.n472 585
R119 B.n472 B.n44 585
R120 B.n471 B.n43 585
R121 B.n521 B.n43 585
R122 B.n470 B.n42 585
R123 B.n522 B.n42 585
R124 B.n469 B.n41 585
R125 B.n523 B.n41 585
R126 B.n468 B.n467 585
R127 B.n467 B.n37 585
R128 B.n466 B.n36 585
R129 B.n529 B.n36 585
R130 B.n465 B.n35 585
R131 B.n530 B.n35 585
R132 B.n464 B.n34 585
R133 B.n531 B.n34 585
R134 B.n463 B.n462 585
R135 B.n462 B.n33 585
R136 B.n461 B.n29 585
R137 B.n537 B.n29 585
R138 B.n460 B.n28 585
R139 B.n538 B.n28 585
R140 B.n459 B.n27 585
R141 B.n539 B.n27 585
R142 B.n458 B.n457 585
R143 B.n457 B.n23 585
R144 B.n456 B.n22 585
R145 B.n545 B.n22 585
R146 B.n455 B.n21 585
R147 B.n546 B.n21 585
R148 B.n454 B.n20 585
R149 B.n547 B.n20 585
R150 B.n453 B.n452 585
R151 B.n452 B.n16 585
R152 B.n451 B.n15 585
R153 B.n553 B.n15 585
R154 B.n450 B.n14 585
R155 B.n554 B.n14 585
R156 B.n449 B.n13 585
R157 B.n555 B.n13 585
R158 B.n448 B.n447 585
R159 B.n447 B.n12 585
R160 B.n446 B.n445 585
R161 B.n446 B.n8 585
R162 B.n444 B.n7 585
R163 B.n562 B.n7 585
R164 B.n443 B.n6 585
R165 B.n563 B.n6 585
R166 B.n442 B.n5 585
R167 B.n564 B.n5 585
R168 B.n441 B.n440 585
R169 B.n440 B.n4 585
R170 B.n439 B.n166 585
R171 B.n439 B.n438 585
R172 B.n429 B.n167 585
R173 B.n168 B.n167 585
R174 B.n431 B.n430 585
R175 B.n432 B.n431 585
R176 B.n428 B.n173 585
R177 B.n173 B.n172 585
R178 B.n427 B.n426 585
R179 B.n426 B.n425 585
R180 B.n175 B.n174 585
R181 B.n176 B.n175 585
R182 B.n418 B.n417 585
R183 B.n419 B.n418 585
R184 B.n416 B.n181 585
R185 B.n181 B.n180 585
R186 B.n415 B.n414 585
R187 B.n414 B.n413 585
R188 B.n183 B.n182 585
R189 B.n184 B.n183 585
R190 B.n406 B.n405 585
R191 B.n407 B.n406 585
R192 B.n404 B.n189 585
R193 B.n189 B.n188 585
R194 B.n403 B.n402 585
R195 B.n402 B.n401 585
R196 B.n191 B.n190 585
R197 B.n394 B.n191 585
R198 B.n393 B.n392 585
R199 B.n395 B.n393 585
R200 B.n391 B.n196 585
R201 B.n196 B.n195 585
R202 B.n390 B.n389 585
R203 B.n389 B.n388 585
R204 B.n198 B.n197 585
R205 B.n199 B.n198 585
R206 B.n381 B.n380 585
R207 B.n382 B.n381 585
R208 B.n379 B.n204 585
R209 B.n204 B.n203 585
R210 B.n378 B.n377 585
R211 B.n377 B.n376 585
R212 B.n206 B.n205 585
R213 B.n207 B.n206 585
R214 B.n369 B.n368 585
R215 B.n370 B.n369 585
R216 B.n367 B.n212 585
R217 B.n212 B.n211 585
R218 B.n366 B.n365 585
R219 B.n365 B.n364 585
R220 B.n214 B.n213 585
R221 B.n215 B.n214 585
R222 B.n357 B.n356 585
R223 B.n358 B.n357 585
R224 B.n355 B.n220 585
R225 B.n220 B.n219 585
R226 B.n354 B.n353 585
R227 B.n353 B.n352 585
R228 B.n222 B.n221 585
R229 B.n223 B.n222 585
R230 B.n345 B.n344 585
R231 B.n346 B.n345 585
R232 B.n343 B.n228 585
R233 B.n228 B.n227 585
R234 B.n342 B.n341 585
R235 B.n341 B.n340 585
R236 B.n230 B.n229 585
R237 B.n231 B.n230 585
R238 B.n336 B.n335 585
R239 B.n234 B.n233 585
R240 B.n332 B.n331 585
R241 B.n333 B.n332 585
R242 B.n330 B.n253 585
R243 B.n329 B.n328 585
R244 B.n327 B.n326 585
R245 B.n325 B.n324 585
R246 B.n323 B.n322 585
R247 B.n321 B.n320 585
R248 B.n319 B.n318 585
R249 B.n317 B.n316 585
R250 B.n315 B.n314 585
R251 B.n313 B.n312 585
R252 B.n311 B.n310 585
R253 B.n309 B.n308 585
R254 B.n307 B.n306 585
R255 B.n305 B.n304 585
R256 B.n303 B.n302 585
R257 B.n301 B.n300 585
R258 B.n299 B.n298 585
R259 B.n297 B.n296 585
R260 B.n295 B.n294 585
R261 B.n293 B.n292 585
R262 B.n291 B.n290 585
R263 B.n288 B.n287 585
R264 B.n286 B.n285 585
R265 B.n284 B.n283 585
R266 B.n282 B.n281 585
R267 B.n280 B.n279 585
R268 B.n278 B.n277 585
R269 B.n276 B.n275 585
R270 B.n274 B.n273 585
R271 B.n272 B.n271 585
R272 B.n270 B.n269 585
R273 B.n268 B.n267 585
R274 B.n266 B.n265 585
R275 B.n264 B.n263 585
R276 B.n262 B.n261 585
R277 B.n260 B.n259 585
R278 B.n337 B.n232 585
R279 B.n232 B.n231 585
R280 B.n339 B.n338 585
R281 B.n340 B.n339 585
R282 B.n226 B.n225 585
R283 B.n227 B.n226 585
R284 B.n348 B.n347 585
R285 B.n347 B.n346 585
R286 B.n349 B.n224 585
R287 B.n224 B.n223 585
R288 B.n351 B.n350 585
R289 B.n352 B.n351 585
R290 B.n218 B.n217 585
R291 B.n219 B.n218 585
R292 B.n360 B.n359 585
R293 B.n359 B.n358 585
R294 B.n361 B.n216 585
R295 B.n216 B.n215 585
R296 B.n363 B.n362 585
R297 B.n364 B.n363 585
R298 B.n210 B.n209 585
R299 B.n211 B.n210 585
R300 B.n372 B.n371 585
R301 B.n371 B.n370 585
R302 B.n373 B.n208 585
R303 B.n208 B.n207 585
R304 B.n375 B.n374 585
R305 B.n376 B.n375 585
R306 B.n202 B.n201 585
R307 B.n203 B.n202 585
R308 B.n384 B.n383 585
R309 B.n383 B.n382 585
R310 B.n385 B.n200 585
R311 B.n200 B.n199 585
R312 B.n387 B.n386 585
R313 B.n388 B.n387 585
R314 B.n194 B.n193 585
R315 B.n195 B.n194 585
R316 B.n397 B.n396 585
R317 B.n396 B.n395 585
R318 B.n398 B.n192 585
R319 B.n394 B.n192 585
R320 B.n400 B.n399 585
R321 B.n401 B.n400 585
R322 B.n187 B.n186 585
R323 B.n188 B.n187 585
R324 B.n409 B.n408 585
R325 B.n408 B.n407 585
R326 B.n410 B.n185 585
R327 B.n185 B.n184 585
R328 B.n412 B.n411 585
R329 B.n413 B.n412 585
R330 B.n179 B.n178 585
R331 B.n180 B.n179 585
R332 B.n421 B.n420 585
R333 B.n420 B.n419 585
R334 B.n422 B.n177 585
R335 B.n177 B.n176 585
R336 B.n424 B.n423 585
R337 B.n425 B.n424 585
R338 B.n171 B.n170 585
R339 B.n172 B.n171 585
R340 B.n434 B.n433 585
R341 B.n433 B.n432 585
R342 B.n435 B.n169 585
R343 B.n169 B.n168 585
R344 B.n437 B.n436 585
R345 B.n438 B.n437 585
R346 B.n3 B.n0 585
R347 B.n4 B.n3 585
R348 B.n561 B.n1 585
R349 B.n562 B.n561 585
R350 B.n560 B.n559 585
R351 B.n560 B.n8 585
R352 B.n558 B.n9 585
R353 B.n12 B.n9 585
R354 B.n557 B.n556 585
R355 B.n556 B.n555 585
R356 B.n11 B.n10 585
R357 B.n554 B.n11 585
R358 B.n552 B.n551 585
R359 B.n553 B.n552 585
R360 B.n550 B.n17 585
R361 B.n17 B.n16 585
R362 B.n549 B.n548 585
R363 B.n548 B.n547 585
R364 B.n19 B.n18 585
R365 B.n546 B.n19 585
R366 B.n544 B.n543 585
R367 B.n545 B.n544 585
R368 B.n542 B.n24 585
R369 B.n24 B.n23 585
R370 B.n541 B.n540 585
R371 B.n540 B.n539 585
R372 B.n26 B.n25 585
R373 B.n538 B.n26 585
R374 B.n536 B.n535 585
R375 B.n537 B.n536 585
R376 B.n534 B.n30 585
R377 B.n33 B.n30 585
R378 B.n533 B.n532 585
R379 B.n532 B.n531 585
R380 B.n32 B.n31 585
R381 B.n530 B.n32 585
R382 B.n528 B.n527 585
R383 B.n529 B.n528 585
R384 B.n526 B.n38 585
R385 B.n38 B.n37 585
R386 B.n525 B.n524 585
R387 B.n524 B.n523 585
R388 B.n40 B.n39 585
R389 B.n522 B.n40 585
R390 B.n520 B.n519 585
R391 B.n521 B.n520 585
R392 B.n518 B.n45 585
R393 B.n45 B.n44 585
R394 B.n517 B.n516 585
R395 B.n516 B.n515 585
R396 B.n47 B.n46 585
R397 B.n514 B.n47 585
R398 B.n512 B.n511 585
R399 B.n513 B.n512 585
R400 B.n510 B.n52 585
R401 B.n52 B.n51 585
R402 B.n509 B.n508 585
R403 B.n508 B.n507 585
R404 B.n54 B.n53 585
R405 B.n506 B.n54 585
R406 B.n504 B.n503 585
R407 B.n505 B.n504 585
R408 B.n502 B.n59 585
R409 B.n59 B.n58 585
R410 B.n501 B.n500 585
R411 B.n500 B.n499 585
R412 B.n61 B.n60 585
R413 B.n498 B.n61 585
R414 B.n496 B.n495 585
R415 B.n497 B.n496 585
R416 B.n494 B.n66 585
R417 B.n66 B.n65 585
R418 B.n565 B.n564 585
R419 B.n563 B.n2 585
R420 B.n492 B.n66 502.111
R421 B.n489 B.n88 502.111
R422 B.n259 B.n230 502.111
R423 B.n335 B.n232 502.111
R424 B.n490 B.n86 256.663
R425 B.n490 B.n85 256.663
R426 B.n490 B.n84 256.663
R427 B.n490 B.n83 256.663
R428 B.n490 B.n82 256.663
R429 B.n490 B.n81 256.663
R430 B.n490 B.n80 256.663
R431 B.n490 B.n79 256.663
R432 B.n490 B.n78 256.663
R433 B.n490 B.n77 256.663
R434 B.n490 B.n76 256.663
R435 B.n490 B.n75 256.663
R436 B.n490 B.n74 256.663
R437 B.n490 B.n73 256.663
R438 B.n490 B.n72 256.663
R439 B.n490 B.n71 256.663
R440 B.n490 B.n70 256.663
R441 B.n490 B.n69 256.663
R442 B.n491 B.n490 256.663
R443 B.n334 B.n333 256.663
R444 B.n333 B.n235 256.663
R445 B.n333 B.n236 256.663
R446 B.n333 B.n237 256.663
R447 B.n333 B.n238 256.663
R448 B.n333 B.n239 256.663
R449 B.n333 B.n240 256.663
R450 B.n333 B.n241 256.663
R451 B.n333 B.n242 256.663
R452 B.n333 B.n243 256.663
R453 B.n333 B.n244 256.663
R454 B.n333 B.n245 256.663
R455 B.n333 B.n246 256.663
R456 B.n333 B.n247 256.663
R457 B.n333 B.n248 256.663
R458 B.n333 B.n249 256.663
R459 B.n333 B.n250 256.663
R460 B.n333 B.n251 256.663
R461 B.n333 B.n252 256.663
R462 B.n567 B.n566 256.663
R463 B.n92 B.t15 232.923
R464 B.n89 B.t4 232.923
R465 B.n257 B.t12 232.923
R466 B.n254 B.t8 232.923
R467 B.n333 B.n231 172.15
R468 B.n490 B.n65 172.15
R469 B.n94 B.n68 163.367
R470 B.n98 B.n97 163.367
R471 B.n102 B.n101 163.367
R472 B.n106 B.n105 163.367
R473 B.n110 B.n109 163.367
R474 B.n114 B.n113 163.367
R475 B.n118 B.n117 163.367
R476 B.n123 B.n122 163.367
R477 B.n127 B.n126 163.367
R478 B.n131 B.n130 163.367
R479 B.n135 B.n134 163.367
R480 B.n139 B.n138 163.367
R481 B.n143 B.n142 163.367
R482 B.n147 B.n146 163.367
R483 B.n151 B.n150 163.367
R484 B.n155 B.n154 163.367
R485 B.n159 B.n158 163.367
R486 B.n163 B.n162 163.367
R487 B.n489 B.n87 163.367
R488 B.n341 B.n230 163.367
R489 B.n341 B.n228 163.367
R490 B.n345 B.n228 163.367
R491 B.n345 B.n222 163.367
R492 B.n353 B.n222 163.367
R493 B.n353 B.n220 163.367
R494 B.n357 B.n220 163.367
R495 B.n357 B.n214 163.367
R496 B.n365 B.n214 163.367
R497 B.n365 B.n212 163.367
R498 B.n369 B.n212 163.367
R499 B.n369 B.n206 163.367
R500 B.n377 B.n206 163.367
R501 B.n377 B.n204 163.367
R502 B.n381 B.n204 163.367
R503 B.n381 B.n198 163.367
R504 B.n389 B.n198 163.367
R505 B.n389 B.n196 163.367
R506 B.n393 B.n196 163.367
R507 B.n393 B.n191 163.367
R508 B.n402 B.n191 163.367
R509 B.n402 B.n189 163.367
R510 B.n406 B.n189 163.367
R511 B.n406 B.n183 163.367
R512 B.n414 B.n183 163.367
R513 B.n414 B.n181 163.367
R514 B.n418 B.n181 163.367
R515 B.n418 B.n175 163.367
R516 B.n426 B.n175 163.367
R517 B.n426 B.n173 163.367
R518 B.n431 B.n173 163.367
R519 B.n431 B.n167 163.367
R520 B.n439 B.n167 163.367
R521 B.n440 B.n439 163.367
R522 B.n440 B.n5 163.367
R523 B.n6 B.n5 163.367
R524 B.n7 B.n6 163.367
R525 B.n446 B.n7 163.367
R526 B.n447 B.n446 163.367
R527 B.n447 B.n13 163.367
R528 B.n14 B.n13 163.367
R529 B.n15 B.n14 163.367
R530 B.n452 B.n15 163.367
R531 B.n452 B.n20 163.367
R532 B.n21 B.n20 163.367
R533 B.n22 B.n21 163.367
R534 B.n457 B.n22 163.367
R535 B.n457 B.n27 163.367
R536 B.n28 B.n27 163.367
R537 B.n29 B.n28 163.367
R538 B.n462 B.n29 163.367
R539 B.n462 B.n34 163.367
R540 B.n35 B.n34 163.367
R541 B.n36 B.n35 163.367
R542 B.n467 B.n36 163.367
R543 B.n467 B.n41 163.367
R544 B.n42 B.n41 163.367
R545 B.n43 B.n42 163.367
R546 B.n472 B.n43 163.367
R547 B.n472 B.n48 163.367
R548 B.n49 B.n48 163.367
R549 B.n50 B.n49 163.367
R550 B.n477 B.n50 163.367
R551 B.n477 B.n55 163.367
R552 B.n56 B.n55 163.367
R553 B.n57 B.n56 163.367
R554 B.n482 B.n57 163.367
R555 B.n482 B.n62 163.367
R556 B.n63 B.n62 163.367
R557 B.n64 B.n63 163.367
R558 B.n88 B.n64 163.367
R559 B.n332 B.n234 163.367
R560 B.n332 B.n253 163.367
R561 B.n328 B.n327 163.367
R562 B.n324 B.n323 163.367
R563 B.n320 B.n319 163.367
R564 B.n316 B.n315 163.367
R565 B.n312 B.n311 163.367
R566 B.n308 B.n307 163.367
R567 B.n304 B.n303 163.367
R568 B.n300 B.n299 163.367
R569 B.n296 B.n295 163.367
R570 B.n292 B.n291 163.367
R571 B.n287 B.n286 163.367
R572 B.n283 B.n282 163.367
R573 B.n279 B.n278 163.367
R574 B.n275 B.n274 163.367
R575 B.n271 B.n270 163.367
R576 B.n267 B.n266 163.367
R577 B.n263 B.n262 163.367
R578 B.n339 B.n232 163.367
R579 B.n339 B.n226 163.367
R580 B.n347 B.n226 163.367
R581 B.n347 B.n224 163.367
R582 B.n351 B.n224 163.367
R583 B.n351 B.n218 163.367
R584 B.n359 B.n218 163.367
R585 B.n359 B.n216 163.367
R586 B.n363 B.n216 163.367
R587 B.n363 B.n210 163.367
R588 B.n371 B.n210 163.367
R589 B.n371 B.n208 163.367
R590 B.n375 B.n208 163.367
R591 B.n375 B.n202 163.367
R592 B.n383 B.n202 163.367
R593 B.n383 B.n200 163.367
R594 B.n387 B.n200 163.367
R595 B.n387 B.n194 163.367
R596 B.n396 B.n194 163.367
R597 B.n396 B.n192 163.367
R598 B.n400 B.n192 163.367
R599 B.n400 B.n187 163.367
R600 B.n408 B.n187 163.367
R601 B.n408 B.n185 163.367
R602 B.n412 B.n185 163.367
R603 B.n412 B.n179 163.367
R604 B.n420 B.n179 163.367
R605 B.n420 B.n177 163.367
R606 B.n424 B.n177 163.367
R607 B.n424 B.n171 163.367
R608 B.n433 B.n171 163.367
R609 B.n433 B.n169 163.367
R610 B.n437 B.n169 163.367
R611 B.n437 B.n3 163.367
R612 B.n565 B.n3 163.367
R613 B.n561 B.n2 163.367
R614 B.n561 B.n560 163.367
R615 B.n560 B.n9 163.367
R616 B.n556 B.n9 163.367
R617 B.n556 B.n11 163.367
R618 B.n552 B.n11 163.367
R619 B.n552 B.n17 163.367
R620 B.n548 B.n17 163.367
R621 B.n548 B.n19 163.367
R622 B.n544 B.n19 163.367
R623 B.n544 B.n24 163.367
R624 B.n540 B.n24 163.367
R625 B.n540 B.n26 163.367
R626 B.n536 B.n26 163.367
R627 B.n536 B.n30 163.367
R628 B.n532 B.n30 163.367
R629 B.n532 B.n32 163.367
R630 B.n528 B.n32 163.367
R631 B.n528 B.n38 163.367
R632 B.n524 B.n38 163.367
R633 B.n524 B.n40 163.367
R634 B.n520 B.n40 163.367
R635 B.n520 B.n45 163.367
R636 B.n516 B.n45 163.367
R637 B.n516 B.n47 163.367
R638 B.n512 B.n47 163.367
R639 B.n512 B.n52 163.367
R640 B.n508 B.n52 163.367
R641 B.n508 B.n54 163.367
R642 B.n504 B.n54 163.367
R643 B.n504 B.n59 163.367
R644 B.n500 B.n59 163.367
R645 B.n500 B.n61 163.367
R646 B.n496 B.n61 163.367
R647 B.n496 B.n66 163.367
R648 B.n89 B.t6 138.198
R649 B.n257 B.t14 138.198
R650 B.n92 B.t16 138.196
R651 B.n254 B.t11 138.196
R652 B.n340 B.n231 92.1755
R653 B.n340 B.n227 92.1755
R654 B.n346 B.n227 92.1755
R655 B.n346 B.n223 92.1755
R656 B.n352 B.n223 92.1755
R657 B.n352 B.n219 92.1755
R658 B.n358 B.n219 92.1755
R659 B.n364 B.n215 92.1755
R660 B.n364 B.n211 92.1755
R661 B.n370 B.n211 92.1755
R662 B.n370 B.n207 92.1755
R663 B.n376 B.n207 92.1755
R664 B.n376 B.n203 92.1755
R665 B.n382 B.n203 92.1755
R666 B.n382 B.n199 92.1755
R667 B.n388 B.n199 92.1755
R668 B.n388 B.n195 92.1755
R669 B.n395 B.n195 92.1755
R670 B.n395 B.n394 92.1755
R671 B.n401 B.n188 92.1755
R672 B.n407 B.n188 92.1755
R673 B.n407 B.n184 92.1755
R674 B.n413 B.n184 92.1755
R675 B.n413 B.n180 92.1755
R676 B.n419 B.n180 92.1755
R677 B.n419 B.n176 92.1755
R678 B.n425 B.n176 92.1755
R679 B.n432 B.n172 92.1755
R680 B.n432 B.n168 92.1755
R681 B.n438 B.n168 92.1755
R682 B.n438 B.n4 92.1755
R683 B.n564 B.n4 92.1755
R684 B.n564 B.n563 92.1755
R685 B.n563 B.n562 92.1755
R686 B.n562 B.n8 92.1755
R687 B.n12 B.n8 92.1755
R688 B.n555 B.n12 92.1755
R689 B.n555 B.n554 92.1755
R690 B.n553 B.n16 92.1755
R691 B.n547 B.n16 92.1755
R692 B.n547 B.n546 92.1755
R693 B.n546 B.n545 92.1755
R694 B.n545 B.n23 92.1755
R695 B.n539 B.n23 92.1755
R696 B.n539 B.n538 92.1755
R697 B.n538 B.n537 92.1755
R698 B.n531 B.n33 92.1755
R699 B.n531 B.n530 92.1755
R700 B.n530 B.n529 92.1755
R701 B.n529 B.n37 92.1755
R702 B.n523 B.n37 92.1755
R703 B.n523 B.n522 92.1755
R704 B.n522 B.n521 92.1755
R705 B.n521 B.n44 92.1755
R706 B.n515 B.n44 92.1755
R707 B.n515 B.n514 92.1755
R708 B.n514 B.n513 92.1755
R709 B.n513 B.n51 92.1755
R710 B.n507 B.n506 92.1755
R711 B.n506 B.n505 92.1755
R712 B.n505 B.n58 92.1755
R713 B.n499 B.n58 92.1755
R714 B.n499 B.n498 92.1755
R715 B.n498 B.n497 92.1755
R716 B.n497 B.n65 92.1755
R717 B.n90 B.t7 77.8836
R718 B.n258 B.t13 77.8836
R719 B.n93 B.t17 77.8818
R720 B.n255 B.t10 77.8818
R721 B.n358 B.t9 75.9093
R722 B.n401 B.t1 75.9093
R723 B.n537 B.t2 75.9093
R724 B.n507 B.t5 75.9093
R725 B.n492 B.n491 71.676
R726 B.n94 B.n69 71.676
R727 B.n98 B.n70 71.676
R728 B.n102 B.n71 71.676
R729 B.n106 B.n72 71.676
R730 B.n110 B.n73 71.676
R731 B.n114 B.n74 71.676
R732 B.n118 B.n75 71.676
R733 B.n123 B.n76 71.676
R734 B.n127 B.n77 71.676
R735 B.n131 B.n78 71.676
R736 B.n135 B.n79 71.676
R737 B.n139 B.n80 71.676
R738 B.n143 B.n81 71.676
R739 B.n147 B.n82 71.676
R740 B.n151 B.n83 71.676
R741 B.n155 B.n84 71.676
R742 B.n159 B.n85 71.676
R743 B.n163 B.n86 71.676
R744 B.n87 B.n86 71.676
R745 B.n162 B.n85 71.676
R746 B.n158 B.n84 71.676
R747 B.n154 B.n83 71.676
R748 B.n150 B.n82 71.676
R749 B.n146 B.n81 71.676
R750 B.n142 B.n80 71.676
R751 B.n138 B.n79 71.676
R752 B.n134 B.n78 71.676
R753 B.n130 B.n77 71.676
R754 B.n126 B.n76 71.676
R755 B.n122 B.n75 71.676
R756 B.n117 B.n74 71.676
R757 B.n113 B.n73 71.676
R758 B.n109 B.n72 71.676
R759 B.n105 B.n71 71.676
R760 B.n101 B.n70 71.676
R761 B.n97 B.n69 71.676
R762 B.n491 B.n68 71.676
R763 B.n335 B.n334 71.676
R764 B.n253 B.n235 71.676
R765 B.n327 B.n236 71.676
R766 B.n323 B.n237 71.676
R767 B.n319 B.n238 71.676
R768 B.n315 B.n239 71.676
R769 B.n311 B.n240 71.676
R770 B.n307 B.n241 71.676
R771 B.n303 B.n242 71.676
R772 B.n299 B.n243 71.676
R773 B.n295 B.n244 71.676
R774 B.n291 B.n245 71.676
R775 B.n286 B.n246 71.676
R776 B.n282 B.n247 71.676
R777 B.n278 B.n248 71.676
R778 B.n274 B.n249 71.676
R779 B.n270 B.n250 71.676
R780 B.n266 B.n251 71.676
R781 B.n262 B.n252 71.676
R782 B.n334 B.n234 71.676
R783 B.n328 B.n235 71.676
R784 B.n324 B.n236 71.676
R785 B.n320 B.n237 71.676
R786 B.n316 B.n238 71.676
R787 B.n312 B.n239 71.676
R788 B.n308 B.n240 71.676
R789 B.n304 B.n241 71.676
R790 B.n300 B.n242 71.676
R791 B.n296 B.n243 71.676
R792 B.n292 B.n244 71.676
R793 B.n287 B.n245 71.676
R794 B.n283 B.n246 71.676
R795 B.n279 B.n247 71.676
R796 B.n275 B.n248 71.676
R797 B.n271 B.n249 71.676
R798 B.n267 B.n250 71.676
R799 B.n263 B.n251 71.676
R800 B.n259 B.n252 71.676
R801 B.n566 B.n565 71.676
R802 B.n566 B.n2 71.676
R803 B.t0 B.n172 62.3542
R804 B.n554 B.t3 62.3542
R805 B.n93 B.n92 60.3157
R806 B.n90 B.n89 60.3157
R807 B.n258 B.n257 60.3157
R808 B.n255 B.n254 60.3157
R809 B.n120 B.n93 59.5399
R810 B.n91 B.n90 59.5399
R811 B.n289 B.n258 59.5399
R812 B.n256 B.n255 59.5399
R813 B.n337 B.n336 32.6249
R814 B.n260 B.n229 32.6249
R815 B.n488 B.n487 32.6249
R816 B.n494 B.n493 32.6249
R817 B.n425 B.t0 29.8218
R818 B.t3 B.n553 29.8218
R819 B B.n567 18.0485
R820 B.t9 B.n215 16.2667
R821 B.n394 B.t1 16.2667
R822 B.n33 B.t2 16.2667
R823 B.t5 B.n51 16.2667
R824 B.n338 B.n337 10.6151
R825 B.n338 B.n225 10.6151
R826 B.n348 B.n225 10.6151
R827 B.n349 B.n348 10.6151
R828 B.n350 B.n349 10.6151
R829 B.n350 B.n217 10.6151
R830 B.n360 B.n217 10.6151
R831 B.n361 B.n360 10.6151
R832 B.n362 B.n361 10.6151
R833 B.n362 B.n209 10.6151
R834 B.n372 B.n209 10.6151
R835 B.n373 B.n372 10.6151
R836 B.n374 B.n373 10.6151
R837 B.n374 B.n201 10.6151
R838 B.n384 B.n201 10.6151
R839 B.n385 B.n384 10.6151
R840 B.n386 B.n385 10.6151
R841 B.n386 B.n193 10.6151
R842 B.n397 B.n193 10.6151
R843 B.n398 B.n397 10.6151
R844 B.n399 B.n398 10.6151
R845 B.n399 B.n186 10.6151
R846 B.n409 B.n186 10.6151
R847 B.n410 B.n409 10.6151
R848 B.n411 B.n410 10.6151
R849 B.n411 B.n178 10.6151
R850 B.n421 B.n178 10.6151
R851 B.n422 B.n421 10.6151
R852 B.n423 B.n422 10.6151
R853 B.n423 B.n170 10.6151
R854 B.n434 B.n170 10.6151
R855 B.n435 B.n434 10.6151
R856 B.n436 B.n435 10.6151
R857 B.n436 B.n0 10.6151
R858 B.n336 B.n233 10.6151
R859 B.n331 B.n233 10.6151
R860 B.n331 B.n330 10.6151
R861 B.n330 B.n329 10.6151
R862 B.n329 B.n326 10.6151
R863 B.n326 B.n325 10.6151
R864 B.n325 B.n322 10.6151
R865 B.n322 B.n321 10.6151
R866 B.n321 B.n318 10.6151
R867 B.n318 B.n317 10.6151
R868 B.n317 B.n314 10.6151
R869 B.n314 B.n313 10.6151
R870 B.n313 B.n310 10.6151
R871 B.n310 B.n309 10.6151
R872 B.n306 B.n305 10.6151
R873 B.n305 B.n302 10.6151
R874 B.n302 B.n301 10.6151
R875 B.n301 B.n298 10.6151
R876 B.n298 B.n297 10.6151
R877 B.n297 B.n294 10.6151
R878 B.n294 B.n293 10.6151
R879 B.n293 B.n290 10.6151
R880 B.n288 B.n285 10.6151
R881 B.n285 B.n284 10.6151
R882 B.n284 B.n281 10.6151
R883 B.n281 B.n280 10.6151
R884 B.n280 B.n277 10.6151
R885 B.n277 B.n276 10.6151
R886 B.n276 B.n273 10.6151
R887 B.n273 B.n272 10.6151
R888 B.n272 B.n269 10.6151
R889 B.n269 B.n268 10.6151
R890 B.n268 B.n265 10.6151
R891 B.n265 B.n264 10.6151
R892 B.n264 B.n261 10.6151
R893 B.n261 B.n260 10.6151
R894 B.n342 B.n229 10.6151
R895 B.n343 B.n342 10.6151
R896 B.n344 B.n343 10.6151
R897 B.n344 B.n221 10.6151
R898 B.n354 B.n221 10.6151
R899 B.n355 B.n354 10.6151
R900 B.n356 B.n355 10.6151
R901 B.n356 B.n213 10.6151
R902 B.n366 B.n213 10.6151
R903 B.n367 B.n366 10.6151
R904 B.n368 B.n367 10.6151
R905 B.n368 B.n205 10.6151
R906 B.n378 B.n205 10.6151
R907 B.n379 B.n378 10.6151
R908 B.n380 B.n379 10.6151
R909 B.n380 B.n197 10.6151
R910 B.n390 B.n197 10.6151
R911 B.n391 B.n390 10.6151
R912 B.n392 B.n391 10.6151
R913 B.n392 B.n190 10.6151
R914 B.n403 B.n190 10.6151
R915 B.n404 B.n403 10.6151
R916 B.n405 B.n404 10.6151
R917 B.n405 B.n182 10.6151
R918 B.n415 B.n182 10.6151
R919 B.n416 B.n415 10.6151
R920 B.n417 B.n416 10.6151
R921 B.n417 B.n174 10.6151
R922 B.n427 B.n174 10.6151
R923 B.n428 B.n427 10.6151
R924 B.n430 B.n428 10.6151
R925 B.n430 B.n429 10.6151
R926 B.n429 B.n166 10.6151
R927 B.n441 B.n166 10.6151
R928 B.n442 B.n441 10.6151
R929 B.n443 B.n442 10.6151
R930 B.n444 B.n443 10.6151
R931 B.n445 B.n444 10.6151
R932 B.n448 B.n445 10.6151
R933 B.n449 B.n448 10.6151
R934 B.n450 B.n449 10.6151
R935 B.n451 B.n450 10.6151
R936 B.n453 B.n451 10.6151
R937 B.n454 B.n453 10.6151
R938 B.n455 B.n454 10.6151
R939 B.n456 B.n455 10.6151
R940 B.n458 B.n456 10.6151
R941 B.n459 B.n458 10.6151
R942 B.n460 B.n459 10.6151
R943 B.n461 B.n460 10.6151
R944 B.n463 B.n461 10.6151
R945 B.n464 B.n463 10.6151
R946 B.n465 B.n464 10.6151
R947 B.n466 B.n465 10.6151
R948 B.n468 B.n466 10.6151
R949 B.n469 B.n468 10.6151
R950 B.n470 B.n469 10.6151
R951 B.n471 B.n470 10.6151
R952 B.n473 B.n471 10.6151
R953 B.n474 B.n473 10.6151
R954 B.n475 B.n474 10.6151
R955 B.n476 B.n475 10.6151
R956 B.n478 B.n476 10.6151
R957 B.n479 B.n478 10.6151
R958 B.n480 B.n479 10.6151
R959 B.n481 B.n480 10.6151
R960 B.n483 B.n481 10.6151
R961 B.n484 B.n483 10.6151
R962 B.n485 B.n484 10.6151
R963 B.n486 B.n485 10.6151
R964 B.n487 B.n486 10.6151
R965 B.n559 B.n1 10.6151
R966 B.n559 B.n558 10.6151
R967 B.n558 B.n557 10.6151
R968 B.n557 B.n10 10.6151
R969 B.n551 B.n10 10.6151
R970 B.n551 B.n550 10.6151
R971 B.n550 B.n549 10.6151
R972 B.n549 B.n18 10.6151
R973 B.n543 B.n18 10.6151
R974 B.n543 B.n542 10.6151
R975 B.n542 B.n541 10.6151
R976 B.n541 B.n25 10.6151
R977 B.n535 B.n25 10.6151
R978 B.n535 B.n534 10.6151
R979 B.n534 B.n533 10.6151
R980 B.n533 B.n31 10.6151
R981 B.n527 B.n31 10.6151
R982 B.n527 B.n526 10.6151
R983 B.n526 B.n525 10.6151
R984 B.n525 B.n39 10.6151
R985 B.n519 B.n39 10.6151
R986 B.n519 B.n518 10.6151
R987 B.n518 B.n517 10.6151
R988 B.n517 B.n46 10.6151
R989 B.n511 B.n46 10.6151
R990 B.n511 B.n510 10.6151
R991 B.n510 B.n509 10.6151
R992 B.n509 B.n53 10.6151
R993 B.n503 B.n53 10.6151
R994 B.n503 B.n502 10.6151
R995 B.n502 B.n501 10.6151
R996 B.n501 B.n60 10.6151
R997 B.n495 B.n60 10.6151
R998 B.n495 B.n494 10.6151
R999 B.n493 B.n67 10.6151
R1000 B.n95 B.n67 10.6151
R1001 B.n96 B.n95 10.6151
R1002 B.n99 B.n96 10.6151
R1003 B.n100 B.n99 10.6151
R1004 B.n103 B.n100 10.6151
R1005 B.n104 B.n103 10.6151
R1006 B.n107 B.n104 10.6151
R1007 B.n108 B.n107 10.6151
R1008 B.n111 B.n108 10.6151
R1009 B.n112 B.n111 10.6151
R1010 B.n115 B.n112 10.6151
R1011 B.n116 B.n115 10.6151
R1012 B.n119 B.n116 10.6151
R1013 B.n124 B.n121 10.6151
R1014 B.n125 B.n124 10.6151
R1015 B.n128 B.n125 10.6151
R1016 B.n129 B.n128 10.6151
R1017 B.n132 B.n129 10.6151
R1018 B.n133 B.n132 10.6151
R1019 B.n136 B.n133 10.6151
R1020 B.n137 B.n136 10.6151
R1021 B.n141 B.n140 10.6151
R1022 B.n144 B.n141 10.6151
R1023 B.n145 B.n144 10.6151
R1024 B.n148 B.n145 10.6151
R1025 B.n149 B.n148 10.6151
R1026 B.n152 B.n149 10.6151
R1027 B.n153 B.n152 10.6151
R1028 B.n156 B.n153 10.6151
R1029 B.n157 B.n156 10.6151
R1030 B.n160 B.n157 10.6151
R1031 B.n161 B.n160 10.6151
R1032 B.n164 B.n161 10.6151
R1033 B.n165 B.n164 10.6151
R1034 B.n488 B.n165 10.6151
R1035 B.n567 B.n0 8.11757
R1036 B.n567 B.n1 8.11757
R1037 B.n306 B.n256 6.5566
R1038 B.n290 B.n289 6.5566
R1039 B.n121 B.n120 6.5566
R1040 B.n137 B.n91 6.5566
R1041 B.n309 B.n256 4.05904
R1042 B.n289 B.n288 4.05904
R1043 B.n120 B.n119 4.05904
R1044 B.n140 B.n91 4.05904
R1045 VN.n0 VN.t0 59.4693
R1046 VN.n1 VN.t1 59.4693
R1047 VN.n0 VN.t3 58.5833
R1048 VN.n1 VN.t2 58.5833
R1049 VN VN.n1 43.6879
R1050 VN VN.n0 3.525
R1051 VDD2.n2 VDD2.n0 116.587
R1052 VDD2.n2 VDD2.n1 82.38
R1053 VDD2.n1 VDD2.t1 6.97233
R1054 VDD2.n1 VDD2.t2 6.97233
R1055 VDD2.n0 VDD2.t3 6.97233
R1056 VDD2.n0 VDD2.t0 6.97233
R1057 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 1.91432f
C1 VDD2 VTAIL 3.37129f
C2 VP VDD1 1.64599f
C3 VDD1 VTAIL 3.31587f
C4 VP VTAIL 1.92843f
C5 VN VDD2 1.39027f
C6 VN VDD1 0.154356f
C7 VDD2 VDD1 1.06463f
C8 VN VP 4.62748f
C9 VP VDD2 0.411614f
C10 VDD2 B 3.092804f
C11 VDD1 B 5.4365f
C12 VTAIL B 4.274913f
C13 VN B 9.621389f
C14 VP B 8.479405f
C15 VDD2.t3 B 0.046132f
C16 VDD2.t0 B 0.046132f
C17 VDD2.n0 B 0.577436f
C18 VDD2.t1 B 0.046132f
C19 VDD2.t2 B 0.046132f
C20 VDD2.n1 B 0.338165f
C21 VDD2.n2 B 2.11787f
C22 VN.t0 B 0.526667f
C23 VN.t3 B 0.522535f
C24 VN.n0 B 0.326352f
C25 VN.t1 B 0.526667f
C26 VN.t2 B 0.522535f
C27 VN.n1 B 1.16856f
C28 VDD1.t1 B 0.043797f
C29 VDD1.t3 B 0.043797f
C30 VDD1.n0 B 0.32128f
C31 VDD1.t0 B 0.043797f
C32 VDD1.t2 B 0.043797f
C33 VDD1.n1 B 0.562357f
C34 VTAIL.t3 B 0.298911f
C35 VTAIL.n0 B 0.247962f
C36 VTAIL.t4 B 0.298911f
C37 VTAIL.n1 B 0.313117f
C38 VTAIL.t5 B 0.298911f
C39 VTAIL.n2 B 0.764061f
C40 VTAIL.t1 B 0.298912f
C41 VTAIL.n3 B 0.76406f
C42 VTAIL.t0 B 0.298912f
C43 VTAIL.n4 B 0.313116f
C44 VTAIL.t6 B 0.298912f
C45 VTAIL.n5 B 0.313116f
C46 VTAIL.t7 B 0.298911f
C47 VTAIL.n6 B 0.764061f
C48 VTAIL.t2 B 0.298911f
C49 VTAIL.n7 B 0.692993f
C50 VP.n0 B 0.024601f
C51 VP.t1 B 0.364427f
C52 VP.n1 B 0.036893f
C53 VP.n2 B 0.018661f
C54 VP.n3 B 0.0194f
C55 VP.t0 B 0.525515f
C56 VP.t2 B 0.52967f
C57 VP.n4 B 1.16515f
C58 VP.t3 B 0.364427f
C59 VP.n5 B 0.213995f
C60 VP.n6 B 0.826204f
C61 VP.n7 B 0.024601f
C62 VP.n8 B 0.018661f
C63 VP.n9 B 0.034605f
C64 VP.n10 B 0.036893f
C65 VP.n11 B 0.015072f
C66 VP.n12 B 0.018661f
C67 VP.n13 B 0.018661f
C68 VP.n14 B 0.018661f
C69 VP.n15 B 0.034605f
C70 VP.n16 B 0.0194f
C71 VP.n17 B 0.213995f
C72 VP.n18 B 0.034706f
.ends

