* NGSPICE file created from diff_pair_sample_0508.ext - technology: sky130A

.subckt diff_pair_sample_0508 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=1.2639 ps=7.99 w=7.66 l=3.45
X1 VTAIL.t11 VP.t1 VDD1.t8 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X2 VDD1.t7 VP.t2 VTAIL.t12 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=2.9874 ps=16.1 w=7.66 l=3.45
X3 VTAIL.t8 VN.t0 VDD2.t9 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X4 VDD2.t8 VN.t1 VTAIL.t5 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X5 VDD2.t7 VN.t2 VTAIL.t3 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=2.9874 ps=16.1 w=7.66 l=3.45
X6 VTAIL.t9 VN.t3 VDD2.t6 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X7 VTAIL.t15 VP.t3 VDD1.t6 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X8 VDD2.t5 VN.t4 VTAIL.t2 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=1.2639 ps=7.99 w=7.66 l=3.45
X9 VTAIL.t14 VP.t4 VDD1.t5 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X10 B.t11 B.t9 B.t10 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=0 ps=0 w=7.66 l=3.45
X11 B.t8 B.t6 B.t7 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=0 ps=0 w=7.66 l=3.45
X12 VDD2.t4 VN.t5 VTAIL.t1 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=2.9874 ps=16.1 w=7.66 l=3.45
X13 B.t5 B.t3 B.t4 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=0 ps=0 w=7.66 l=3.45
X14 VDD1.t4 VP.t5 VTAIL.t19 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=1.2639 ps=7.99 w=7.66 l=3.45
X15 VDD2.t3 VN.t6 VTAIL.t7 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X16 VDD1.t3 VP.t6 VTAIL.t13 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X17 B.t2 B.t0 B.t1 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=0 ps=0 w=7.66 l=3.45
X18 VTAIL.t6 VN.t7 VDD2.t2 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X19 VDD1.t2 VP.t7 VTAIL.t18 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X20 VTAIL.t4 VN.t8 VDD2.t1 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X21 VDD2.t0 VN.t9 VTAIL.t0 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=2.9874 pd=16.1 as=1.2639 ps=7.99 w=7.66 l=3.45
X22 VTAIL.t10 VP.t8 VDD1.t1 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=1.2639 ps=7.99 w=7.66 l=3.45
X23 VDD1.t0 VP.t9 VTAIL.t17 w_n5506_n2500# sky130_fd_pr__pfet_01v8 ad=1.2639 pd=7.99 as=2.9874 ps=16.1 w=7.66 l=3.45
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n20 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n19 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n18 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n117 VP.n116 161.3
R24 VP.n115 VP.n1 161.3
R25 VP.n114 VP.n113 161.3
R26 VP.n112 VP.n2 161.3
R27 VP.n111 VP.n110 161.3
R28 VP.n109 VP.n3 161.3
R29 VP.n108 VP.n107 161.3
R30 VP.n106 VP.n105 161.3
R31 VP.n104 VP.n5 161.3
R32 VP.n103 VP.n102 161.3
R33 VP.n101 VP.n6 161.3
R34 VP.n100 VP.n99 161.3
R35 VP.n98 VP.n7 161.3
R36 VP.n97 VP.n96 161.3
R37 VP.n95 VP.n8 161.3
R38 VP.n94 VP.n93 161.3
R39 VP.n91 VP.n9 161.3
R40 VP.n90 VP.n89 161.3
R41 VP.n88 VP.n10 161.3
R42 VP.n87 VP.n86 161.3
R43 VP.n85 VP.n11 161.3
R44 VP.n84 VP.n83 161.3
R45 VP.n82 VP.n12 161.3
R46 VP.n81 VP.n80 161.3
R47 VP.n78 VP.n13 161.3
R48 VP.n77 VP.n76 161.3
R49 VP.n75 VP.n14 161.3
R50 VP.n74 VP.n73 161.3
R51 VP.n72 VP.n15 161.3
R52 VP.n71 VP.n70 161.3
R53 VP.n31 VP.t5 86.4515
R54 VP.n69 VP.n16 74.9986
R55 VP.n118 VP.n0 74.9986
R56 VP.n68 VP.n17 74.9986
R57 VP.n31 VP.n30 73.4663
R58 VP.n69 VP.n68 54.6056
R59 VP.n86 VP.n10 54.1398
R60 VP.n99 VP.n6 54.1398
R61 VP.n49 VP.n23 54.1398
R62 VP.n36 VP.n27 54.1398
R63 VP.n16 VP.t0 53.5095
R64 VP.n79 VP.t8 53.5095
R65 VP.n92 VP.t6 53.5095
R66 VP.n4 VP.t4 53.5095
R67 VP.n0 VP.t9 53.5095
R68 VP.n17 VP.t2 53.5095
R69 VP.n21 VP.t3 53.5095
R70 VP.n42 VP.t7 53.5095
R71 VP.n30 VP.t1 53.5095
R72 VP.n77 VP.n14 48.3272
R73 VP.n110 VP.n2 48.3272
R74 VP.n60 VP.n19 48.3272
R75 VP.n73 VP.n14 32.8269
R76 VP.n114 VP.n2 32.8269
R77 VP.n64 VP.n19 32.8269
R78 VP.n90 VP.n10 27.0143
R79 VP.n99 VP.n98 27.0143
R80 VP.n49 VP.n48 27.0143
R81 VP.n40 VP.n27 27.0143
R82 VP.n72 VP.n71 24.5923
R83 VP.n73 VP.n72 24.5923
R84 VP.n78 VP.n77 24.5923
R85 VP.n80 VP.n78 24.5923
R86 VP.n84 VP.n12 24.5923
R87 VP.n85 VP.n84 24.5923
R88 VP.n86 VP.n85 24.5923
R89 VP.n91 VP.n90 24.5923
R90 VP.n93 VP.n91 24.5923
R91 VP.n97 VP.n8 24.5923
R92 VP.n98 VP.n97 24.5923
R93 VP.n103 VP.n6 24.5923
R94 VP.n104 VP.n103 24.5923
R95 VP.n105 VP.n104 24.5923
R96 VP.n109 VP.n108 24.5923
R97 VP.n110 VP.n109 24.5923
R98 VP.n115 VP.n114 24.5923
R99 VP.n116 VP.n115 24.5923
R100 VP.n65 VP.n64 24.5923
R101 VP.n66 VP.n65 24.5923
R102 VP.n53 VP.n23 24.5923
R103 VP.n54 VP.n53 24.5923
R104 VP.n55 VP.n54 24.5923
R105 VP.n59 VP.n58 24.5923
R106 VP.n60 VP.n59 24.5923
R107 VP.n41 VP.n40 24.5923
R108 VP.n43 VP.n41 24.5923
R109 VP.n47 VP.n25 24.5923
R110 VP.n48 VP.n47 24.5923
R111 VP.n34 VP.n29 24.5923
R112 VP.n35 VP.n34 24.5923
R113 VP.n36 VP.n35 24.5923
R114 VP.n80 VP.n79 23.1168
R115 VP.n108 VP.n4 23.1168
R116 VP.n58 VP.n21 23.1168
R117 VP.n71 VP.n16 15.2474
R118 VP.n116 VP.n0 15.2474
R119 VP.n66 VP.n17 15.2474
R120 VP.n93 VP.n92 12.2964
R121 VP.n92 VP.n8 12.2964
R122 VP.n43 VP.n42 12.2964
R123 VP.n42 VP.n25 12.2964
R124 VP.n32 VP.n31 4.13276
R125 VP.n79 VP.n12 1.47601
R126 VP.n105 VP.n4 1.47601
R127 VP.n55 VP.n21 1.47601
R128 VP.n30 VP.n29 1.47601
R129 VP.n68 VP.n67 0.354861
R130 VP.n70 VP.n69 0.354861
R131 VP.n118 VP.n117 0.354861
R132 VP VP.n118 0.267071
R133 VP.n33 VP.n32 0.189894
R134 VP.n33 VP.n28 0.189894
R135 VP.n37 VP.n28 0.189894
R136 VP.n38 VP.n37 0.189894
R137 VP.n39 VP.n38 0.189894
R138 VP.n39 VP.n26 0.189894
R139 VP.n44 VP.n26 0.189894
R140 VP.n45 VP.n44 0.189894
R141 VP.n46 VP.n45 0.189894
R142 VP.n46 VP.n24 0.189894
R143 VP.n50 VP.n24 0.189894
R144 VP.n51 VP.n50 0.189894
R145 VP.n52 VP.n51 0.189894
R146 VP.n52 VP.n22 0.189894
R147 VP.n56 VP.n22 0.189894
R148 VP.n57 VP.n56 0.189894
R149 VP.n57 VP.n20 0.189894
R150 VP.n61 VP.n20 0.189894
R151 VP.n62 VP.n61 0.189894
R152 VP.n63 VP.n62 0.189894
R153 VP.n63 VP.n18 0.189894
R154 VP.n67 VP.n18 0.189894
R155 VP.n70 VP.n15 0.189894
R156 VP.n74 VP.n15 0.189894
R157 VP.n75 VP.n74 0.189894
R158 VP.n76 VP.n75 0.189894
R159 VP.n76 VP.n13 0.189894
R160 VP.n81 VP.n13 0.189894
R161 VP.n82 VP.n81 0.189894
R162 VP.n83 VP.n82 0.189894
R163 VP.n83 VP.n11 0.189894
R164 VP.n87 VP.n11 0.189894
R165 VP.n88 VP.n87 0.189894
R166 VP.n89 VP.n88 0.189894
R167 VP.n89 VP.n9 0.189894
R168 VP.n94 VP.n9 0.189894
R169 VP.n95 VP.n94 0.189894
R170 VP.n96 VP.n95 0.189894
R171 VP.n96 VP.n7 0.189894
R172 VP.n100 VP.n7 0.189894
R173 VP.n101 VP.n100 0.189894
R174 VP.n102 VP.n101 0.189894
R175 VP.n102 VP.n5 0.189894
R176 VP.n106 VP.n5 0.189894
R177 VP.n107 VP.n106 0.189894
R178 VP.n107 VP.n3 0.189894
R179 VP.n111 VP.n3 0.189894
R180 VP.n112 VP.n111 0.189894
R181 VP.n113 VP.n112 0.189894
R182 VP.n113 VP.n1 0.189894
R183 VP.n117 VP.n1 0.189894
R184 VTAIL.n11 VTAIL.t1 75.3715
R185 VTAIL.n17 VTAIL.t3 75.3713
R186 VTAIL.n2 VTAIL.t17 75.3713
R187 VTAIL.n16 VTAIL.t12 75.3713
R188 VTAIL.n15 VTAIL.n14 71.128
R189 VTAIL.n13 VTAIL.n12 71.128
R190 VTAIL.n10 VTAIL.n9 71.128
R191 VTAIL.n8 VTAIL.n7 71.128
R192 VTAIL.n19 VTAIL.n18 71.1278
R193 VTAIL.n1 VTAIL.n0 71.1278
R194 VTAIL.n4 VTAIL.n3 71.1278
R195 VTAIL.n6 VTAIL.n5 71.1278
R196 VTAIL.n8 VTAIL.n6 25.4876
R197 VTAIL.n17 VTAIL.n16 22.2289
R198 VTAIL.n18 VTAIL.t7 4.24397
R199 VTAIL.n18 VTAIL.t6 4.24397
R200 VTAIL.n0 VTAIL.t0 4.24397
R201 VTAIL.n0 VTAIL.t9 4.24397
R202 VTAIL.n3 VTAIL.t13 4.24397
R203 VTAIL.n3 VTAIL.t14 4.24397
R204 VTAIL.n5 VTAIL.t16 4.24397
R205 VTAIL.n5 VTAIL.t10 4.24397
R206 VTAIL.n14 VTAIL.t18 4.24397
R207 VTAIL.n14 VTAIL.t15 4.24397
R208 VTAIL.n12 VTAIL.t19 4.24397
R209 VTAIL.n12 VTAIL.t11 4.24397
R210 VTAIL.n9 VTAIL.t5 4.24397
R211 VTAIL.n9 VTAIL.t8 4.24397
R212 VTAIL.n7 VTAIL.t2 4.24397
R213 VTAIL.n7 VTAIL.t4 4.24397
R214 VTAIL.n10 VTAIL.n8 3.25912
R215 VTAIL.n11 VTAIL.n10 3.25912
R216 VTAIL.n15 VTAIL.n13 3.25912
R217 VTAIL.n16 VTAIL.n15 3.25912
R218 VTAIL.n6 VTAIL.n4 3.25912
R219 VTAIL.n4 VTAIL.n2 3.25912
R220 VTAIL.n19 VTAIL.n17 3.25912
R221 VTAIL VTAIL.n1 2.50266
R222 VTAIL.n13 VTAIL.n11 2.09964
R223 VTAIL.n2 VTAIL.n1 2.09964
R224 VTAIL VTAIL.n19 0.756965
R225 VDD1.n1 VDD1.t4 95.3089
R226 VDD1.n3 VDD1.t9 95.3087
R227 VDD1.n5 VDD1.n4 90.1952
R228 VDD1.n1 VDD1.n0 87.8068
R229 VDD1.n7 VDD1.n6 87.8066
R230 VDD1.n3 VDD1.n2 87.8066
R231 VDD1.n7 VDD1.n5 48.0095
R232 VDD1.n6 VDD1.t6 4.24397
R233 VDD1.n6 VDD1.t7 4.24397
R234 VDD1.n0 VDD1.t8 4.24397
R235 VDD1.n0 VDD1.t2 4.24397
R236 VDD1.n4 VDD1.t5 4.24397
R237 VDD1.n4 VDD1.t0 4.24397
R238 VDD1.n2 VDD1.t1 4.24397
R239 VDD1.n2 VDD1.t3 4.24397
R240 VDD1 VDD1.n7 2.38628
R241 VDD1 VDD1.n1 0.873345
R242 VDD1.n5 VDD1.n3 0.759809
R243 VN.n102 VN.n101 161.3
R244 VN.n100 VN.n53 161.3
R245 VN.n99 VN.n98 161.3
R246 VN.n97 VN.n54 161.3
R247 VN.n96 VN.n95 161.3
R248 VN.n94 VN.n55 161.3
R249 VN.n93 VN.n92 161.3
R250 VN.n91 VN.n90 161.3
R251 VN.n89 VN.n57 161.3
R252 VN.n88 VN.n87 161.3
R253 VN.n86 VN.n58 161.3
R254 VN.n85 VN.n84 161.3
R255 VN.n83 VN.n59 161.3
R256 VN.n82 VN.n81 161.3
R257 VN.n80 VN.n60 161.3
R258 VN.n79 VN.n78 161.3
R259 VN.n77 VN.n61 161.3
R260 VN.n76 VN.n75 161.3
R261 VN.n74 VN.n63 161.3
R262 VN.n73 VN.n72 161.3
R263 VN.n71 VN.n64 161.3
R264 VN.n70 VN.n69 161.3
R265 VN.n68 VN.n65 161.3
R266 VN.n50 VN.n49 161.3
R267 VN.n48 VN.n1 161.3
R268 VN.n47 VN.n46 161.3
R269 VN.n45 VN.n2 161.3
R270 VN.n44 VN.n43 161.3
R271 VN.n42 VN.n3 161.3
R272 VN.n41 VN.n40 161.3
R273 VN.n39 VN.n38 161.3
R274 VN.n37 VN.n5 161.3
R275 VN.n36 VN.n35 161.3
R276 VN.n34 VN.n6 161.3
R277 VN.n33 VN.n32 161.3
R278 VN.n31 VN.n7 161.3
R279 VN.n30 VN.n29 161.3
R280 VN.n28 VN.n8 161.3
R281 VN.n27 VN.n26 161.3
R282 VN.n24 VN.n9 161.3
R283 VN.n23 VN.n22 161.3
R284 VN.n21 VN.n10 161.3
R285 VN.n20 VN.n19 161.3
R286 VN.n18 VN.n11 161.3
R287 VN.n17 VN.n16 161.3
R288 VN.n15 VN.n12 161.3
R289 VN.n67 VN.t5 86.4517
R290 VN.n14 VN.t9 86.4517
R291 VN.n51 VN.n0 74.9986
R292 VN.n103 VN.n52 74.9986
R293 VN.n14 VN.n13 73.4663
R294 VN.n67 VN.n66 73.4663
R295 VN VN.n103 54.7709
R296 VN.n19 VN.n10 54.1398
R297 VN.n32 VN.n6 54.1398
R298 VN.n72 VN.n63 54.1398
R299 VN.n84 VN.n58 54.1398
R300 VN.n13 VN.t3 53.5095
R301 VN.n25 VN.t6 53.5095
R302 VN.n4 VN.t7 53.5095
R303 VN.n0 VN.t2 53.5095
R304 VN.n66 VN.t0 53.5095
R305 VN.n62 VN.t1 53.5095
R306 VN.n56 VN.t8 53.5095
R307 VN.n52 VN.t4 53.5095
R308 VN.n43 VN.n2 48.3272
R309 VN.n95 VN.n54 48.3272
R310 VN.n47 VN.n2 32.8269
R311 VN.n99 VN.n54 32.8269
R312 VN.n23 VN.n10 27.0143
R313 VN.n32 VN.n31 27.0143
R314 VN.n76 VN.n63 27.0143
R315 VN.n84 VN.n83 27.0143
R316 VN.n17 VN.n12 24.5923
R317 VN.n18 VN.n17 24.5923
R318 VN.n19 VN.n18 24.5923
R319 VN.n24 VN.n23 24.5923
R320 VN.n26 VN.n24 24.5923
R321 VN.n30 VN.n8 24.5923
R322 VN.n31 VN.n30 24.5923
R323 VN.n36 VN.n6 24.5923
R324 VN.n37 VN.n36 24.5923
R325 VN.n38 VN.n37 24.5923
R326 VN.n42 VN.n41 24.5923
R327 VN.n43 VN.n42 24.5923
R328 VN.n48 VN.n47 24.5923
R329 VN.n49 VN.n48 24.5923
R330 VN.n72 VN.n71 24.5923
R331 VN.n71 VN.n70 24.5923
R332 VN.n70 VN.n65 24.5923
R333 VN.n83 VN.n82 24.5923
R334 VN.n82 VN.n60 24.5923
R335 VN.n78 VN.n77 24.5923
R336 VN.n77 VN.n76 24.5923
R337 VN.n95 VN.n94 24.5923
R338 VN.n94 VN.n93 24.5923
R339 VN.n90 VN.n89 24.5923
R340 VN.n89 VN.n88 24.5923
R341 VN.n88 VN.n58 24.5923
R342 VN.n101 VN.n100 24.5923
R343 VN.n100 VN.n99 24.5923
R344 VN.n41 VN.n4 23.1168
R345 VN.n93 VN.n56 23.1168
R346 VN.n49 VN.n0 15.2474
R347 VN.n101 VN.n52 15.2474
R348 VN.n26 VN.n25 12.2964
R349 VN.n25 VN.n8 12.2964
R350 VN.n62 VN.n60 12.2964
R351 VN.n78 VN.n62 12.2964
R352 VN.n68 VN.n67 4.13278
R353 VN.n15 VN.n14 4.13278
R354 VN.n13 VN.n12 1.47601
R355 VN.n38 VN.n4 1.47601
R356 VN.n66 VN.n65 1.47601
R357 VN.n90 VN.n56 1.47601
R358 VN.n103 VN.n102 0.354861
R359 VN.n51 VN.n50 0.354861
R360 VN VN.n51 0.267071
R361 VN.n102 VN.n53 0.189894
R362 VN.n98 VN.n53 0.189894
R363 VN.n98 VN.n97 0.189894
R364 VN.n97 VN.n96 0.189894
R365 VN.n96 VN.n55 0.189894
R366 VN.n92 VN.n55 0.189894
R367 VN.n92 VN.n91 0.189894
R368 VN.n91 VN.n57 0.189894
R369 VN.n87 VN.n57 0.189894
R370 VN.n87 VN.n86 0.189894
R371 VN.n86 VN.n85 0.189894
R372 VN.n85 VN.n59 0.189894
R373 VN.n81 VN.n59 0.189894
R374 VN.n81 VN.n80 0.189894
R375 VN.n80 VN.n79 0.189894
R376 VN.n79 VN.n61 0.189894
R377 VN.n75 VN.n61 0.189894
R378 VN.n75 VN.n74 0.189894
R379 VN.n74 VN.n73 0.189894
R380 VN.n73 VN.n64 0.189894
R381 VN.n69 VN.n64 0.189894
R382 VN.n69 VN.n68 0.189894
R383 VN.n16 VN.n15 0.189894
R384 VN.n16 VN.n11 0.189894
R385 VN.n20 VN.n11 0.189894
R386 VN.n21 VN.n20 0.189894
R387 VN.n22 VN.n21 0.189894
R388 VN.n22 VN.n9 0.189894
R389 VN.n27 VN.n9 0.189894
R390 VN.n28 VN.n27 0.189894
R391 VN.n29 VN.n28 0.189894
R392 VN.n29 VN.n7 0.189894
R393 VN.n33 VN.n7 0.189894
R394 VN.n34 VN.n33 0.189894
R395 VN.n35 VN.n34 0.189894
R396 VN.n35 VN.n5 0.189894
R397 VN.n39 VN.n5 0.189894
R398 VN.n40 VN.n39 0.189894
R399 VN.n40 VN.n3 0.189894
R400 VN.n44 VN.n3 0.189894
R401 VN.n45 VN.n44 0.189894
R402 VN.n46 VN.n45 0.189894
R403 VN.n46 VN.n1 0.189894
R404 VN.n50 VN.n1 0.189894
R405 VDD2.n1 VDD2.t0 95.3087
R406 VDD2.n4 VDD2.t5 92.0503
R407 VDD2.n3 VDD2.n2 90.1952
R408 VDD2 VDD2.n7 90.1924
R409 VDD2.n6 VDD2.n5 87.8068
R410 VDD2.n1 VDD2.n0 87.8066
R411 VDD2.n4 VDD2.n3 45.7972
R412 VDD2.n7 VDD2.t9 4.24397
R413 VDD2.n7 VDD2.t4 4.24397
R414 VDD2.n5 VDD2.t1 4.24397
R415 VDD2.n5 VDD2.t8 4.24397
R416 VDD2.n2 VDD2.t2 4.24397
R417 VDD2.n2 VDD2.t7 4.24397
R418 VDD2.n0 VDD2.t6 4.24397
R419 VDD2.n0 VDD2.t3 4.24397
R420 VDD2.n6 VDD2.n4 3.25912
R421 VDD2 VDD2.n6 0.873345
R422 VDD2.n3 VDD2.n1 0.759809
R423 B.n668 B.n77 585
R424 B.n670 B.n669 585
R425 B.n671 B.n76 585
R426 B.n673 B.n672 585
R427 B.n674 B.n75 585
R428 B.n676 B.n675 585
R429 B.n677 B.n74 585
R430 B.n679 B.n678 585
R431 B.n680 B.n73 585
R432 B.n682 B.n681 585
R433 B.n683 B.n72 585
R434 B.n685 B.n684 585
R435 B.n686 B.n71 585
R436 B.n688 B.n687 585
R437 B.n689 B.n70 585
R438 B.n691 B.n690 585
R439 B.n692 B.n69 585
R440 B.n694 B.n693 585
R441 B.n695 B.n68 585
R442 B.n697 B.n696 585
R443 B.n698 B.n67 585
R444 B.n700 B.n699 585
R445 B.n701 B.n66 585
R446 B.n703 B.n702 585
R447 B.n704 B.n65 585
R448 B.n706 B.n705 585
R449 B.n707 B.n64 585
R450 B.n709 B.n708 585
R451 B.n710 B.n61 585
R452 B.n713 B.n712 585
R453 B.n714 B.n60 585
R454 B.n716 B.n715 585
R455 B.n717 B.n59 585
R456 B.n719 B.n718 585
R457 B.n720 B.n58 585
R458 B.n722 B.n721 585
R459 B.n723 B.n57 585
R460 B.n725 B.n724 585
R461 B.n727 B.n726 585
R462 B.n728 B.n53 585
R463 B.n730 B.n729 585
R464 B.n731 B.n52 585
R465 B.n733 B.n732 585
R466 B.n734 B.n51 585
R467 B.n736 B.n735 585
R468 B.n737 B.n50 585
R469 B.n739 B.n738 585
R470 B.n740 B.n49 585
R471 B.n742 B.n741 585
R472 B.n743 B.n48 585
R473 B.n745 B.n744 585
R474 B.n746 B.n47 585
R475 B.n748 B.n747 585
R476 B.n749 B.n46 585
R477 B.n751 B.n750 585
R478 B.n752 B.n45 585
R479 B.n754 B.n753 585
R480 B.n755 B.n44 585
R481 B.n757 B.n756 585
R482 B.n758 B.n43 585
R483 B.n760 B.n759 585
R484 B.n761 B.n42 585
R485 B.n763 B.n762 585
R486 B.n764 B.n41 585
R487 B.n766 B.n765 585
R488 B.n767 B.n40 585
R489 B.n769 B.n768 585
R490 B.n667 B.n666 585
R491 B.n665 B.n78 585
R492 B.n664 B.n663 585
R493 B.n662 B.n79 585
R494 B.n661 B.n660 585
R495 B.n659 B.n80 585
R496 B.n658 B.n657 585
R497 B.n656 B.n81 585
R498 B.n655 B.n654 585
R499 B.n653 B.n82 585
R500 B.n652 B.n651 585
R501 B.n650 B.n83 585
R502 B.n649 B.n648 585
R503 B.n647 B.n84 585
R504 B.n646 B.n645 585
R505 B.n644 B.n85 585
R506 B.n643 B.n642 585
R507 B.n641 B.n86 585
R508 B.n640 B.n639 585
R509 B.n638 B.n87 585
R510 B.n637 B.n636 585
R511 B.n635 B.n88 585
R512 B.n634 B.n633 585
R513 B.n632 B.n89 585
R514 B.n631 B.n630 585
R515 B.n629 B.n90 585
R516 B.n628 B.n627 585
R517 B.n626 B.n91 585
R518 B.n625 B.n624 585
R519 B.n623 B.n92 585
R520 B.n622 B.n621 585
R521 B.n620 B.n93 585
R522 B.n619 B.n618 585
R523 B.n617 B.n94 585
R524 B.n616 B.n615 585
R525 B.n614 B.n95 585
R526 B.n613 B.n612 585
R527 B.n611 B.n96 585
R528 B.n610 B.n609 585
R529 B.n608 B.n97 585
R530 B.n607 B.n606 585
R531 B.n605 B.n98 585
R532 B.n604 B.n603 585
R533 B.n602 B.n99 585
R534 B.n601 B.n600 585
R535 B.n599 B.n100 585
R536 B.n598 B.n597 585
R537 B.n596 B.n101 585
R538 B.n595 B.n594 585
R539 B.n593 B.n102 585
R540 B.n592 B.n591 585
R541 B.n590 B.n103 585
R542 B.n589 B.n588 585
R543 B.n587 B.n104 585
R544 B.n586 B.n585 585
R545 B.n584 B.n105 585
R546 B.n583 B.n582 585
R547 B.n581 B.n106 585
R548 B.n580 B.n579 585
R549 B.n578 B.n107 585
R550 B.n577 B.n576 585
R551 B.n575 B.n108 585
R552 B.n574 B.n573 585
R553 B.n572 B.n109 585
R554 B.n571 B.n570 585
R555 B.n569 B.n110 585
R556 B.n568 B.n567 585
R557 B.n566 B.n111 585
R558 B.n565 B.n564 585
R559 B.n563 B.n112 585
R560 B.n562 B.n561 585
R561 B.n560 B.n113 585
R562 B.n559 B.n558 585
R563 B.n557 B.n114 585
R564 B.n556 B.n555 585
R565 B.n554 B.n115 585
R566 B.n553 B.n552 585
R567 B.n551 B.n116 585
R568 B.n550 B.n549 585
R569 B.n548 B.n117 585
R570 B.n547 B.n546 585
R571 B.n545 B.n118 585
R572 B.n544 B.n543 585
R573 B.n542 B.n119 585
R574 B.n541 B.n540 585
R575 B.n539 B.n120 585
R576 B.n538 B.n537 585
R577 B.n536 B.n121 585
R578 B.n535 B.n534 585
R579 B.n533 B.n122 585
R580 B.n532 B.n531 585
R581 B.n530 B.n123 585
R582 B.n529 B.n528 585
R583 B.n527 B.n124 585
R584 B.n526 B.n525 585
R585 B.n524 B.n125 585
R586 B.n523 B.n522 585
R587 B.n521 B.n126 585
R588 B.n520 B.n519 585
R589 B.n518 B.n127 585
R590 B.n517 B.n516 585
R591 B.n515 B.n128 585
R592 B.n514 B.n513 585
R593 B.n512 B.n129 585
R594 B.n511 B.n510 585
R595 B.n509 B.n130 585
R596 B.n508 B.n507 585
R597 B.n506 B.n131 585
R598 B.n505 B.n504 585
R599 B.n503 B.n132 585
R600 B.n502 B.n501 585
R601 B.n500 B.n133 585
R602 B.n499 B.n498 585
R603 B.n497 B.n134 585
R604 B.n496 B.n495 585
R605 B.n494 B.n135 585
R606 B.n493 B.n492 585
R607 B.n491 B.n136 585
R608 B.n490 B.n489 585
R609 B.n488 B.n137 585
R610 B.n487 B.n486 585
R611 B.n485 B.n138 585
R612 B.n484 B.n483 585
R613 B.n482 B.n139 585
R614 B.n481 B.n480 585
R615 B.n479 B.n140 585
R616 B.n478 B.n477 585
R617 B.n476 B.n141 585
R618 B.n475 B.n474 585
R619 B.n473 B.n142 585
R620 B.n472 B.n471 585
R621 B.n470 B.n143 585
R622 B.n469 B.n468 585
R623 B.n467 B.n144 585
R624 B.n466 B.n465 585
R625 B.n464 B.n145 585
R626 B.n463 B.n462 585
R627 B.n461 B.n146 585
R628 B.n460 B.n459 585
R629 B.n458 B.n147 585
R630 B.n457 B.n456 585
R631 B.n455 B.n148 585
R632 B.n454 B.n453 585
R633 B.n452 B.n149 585
R634 B.n451 B.n450 585
R635 B.n449 B.n150 585
R636 B.n448 B.n447 585
R637 B.n446 B.n151 585
R638 B.n445 B.n444 585
R639 B.n443 B.n152 585
R640 B.n442 B.n441 585
R641 B.n340 B.n339 585
R642 B.n341 B.n190 585
R643 B.n343 B.n342 585
R644 B.n344 B.n189 585
R645 B.n346 B.n345 585
R646 B.n347 B.n188 585
R647 B.n349 B.n348 585
R648 B.n350 B.n187 585
R649 B.n352 B.n351 585
R650 B.n353 B.n186 585
R651 B.n355 B.n354 585
R652 B.n356 B.n185 585
R653 B.n358 B.n357 585
R654 B.n359 B.n184 585
R655 B.n361 B.n360 585
R656 B.n362 B.n183 585
R657 B.n364 B.n363 585
R658 B.n365 B.n182 585
R659 B.n367 B.n366 585
R660 B.n368 B.n181 585
R661 B.n370 B.n369 585
R662 B.n371 B.n180 585
R663 B.n373 B.n372 585
R664 B.n374 B.n179 585
R665 B.n376 B.n375 585
R666 B.n377 B.n178 585
R667 B.n379 B.n378 585
R668 B.n380 B.n177 585
R669 B.n382 B.n381 585
R670 B.n384 B.n383 585
R671 B.n385 B.n173 585
R672 B.n387 B.n386 585
R673 B.n388 B.n172 585
R674 B.n390 B.n389 585
R675 B.n391 B.n171 585
R676 B.n393 B.n392 585
R677 B.n394 B.n170 585
R678 B.n396 B.n395 585
R679 B.n398 B.n167 585
R680 B.n400 B.n399 585
R681 B.n401 B.n166 585
R682 B.n403 B.n402 585
R683 B.n404 B.n165 585
R684 B.n406 B.n405 585
R685 B.n407 B.n164 585
R686 B.n409 B.n408 585
R687 B.n410 B.n163 585
R688 B.n412 B.n411 585
R689 B.n413 B.n162 585
R690 B.n415 B.n414 585
R691 B.n416 B.n161 585
R692 B.n418 B.n417 585
R693 B.n419 B.n160 585
R694 B.n421 B.n420 585
R695 B.n422 B.n159 585
R696 B.n424 B.n423 585
R697 B.n425 B.n158 585
R698 B.n427 B.n426 585
R699 B.n428 B.n157 585
R700 B.n430 B.n429 585
R701 B.n431 B.n156 585
R702 B.n433 B.n432 585
R703 B.n434 B.n155 585
R704 B.n436 B.n435 585
R705 B.n437 B.n154 585
R706 B.n439 B.n438 585
R707 B.n440 B.n153 585
R708 B.n338 B.n191 585
R709 B.n337 B.n336 585
R710 B.n335 B.n192 585
R711 B.n334 B.n333 585
R712 B.n332 B.n193 585
R713 B.n331 B.n330 585
R714 B.n329 B.n194 585
R715 B.n328 B.n327 585
R716 B.n326 B.n195 585
R717 B.n325 B.n324 585
R718 B.n323 B.n196 585
R719 B.n322 B.n321 585
R720 B.n320 B.n197 585
R721 B.n319 B.n318 585
R722 B.n317 B.n198 585
R723 B.n316 B.n315 585
R724 B.n314 B.n199 585
R725 B.n313 B.n312 585
R726 B.n311 B.n200 585
R727 B.n310 B.n309 585
R728 B.n308 B.n201 585
R729 B.n307 B.n306 585
R730 B.n305 B.n202 585
R731 B.n304 B.n303 585
R732 B.n302 B.n203 585
R733 B.n301 B.n300 585
R734 B.n299 B.n204 585
R735 B.n298 B.n297 585
R736 B.n296 B.n205 585
R737 B.n295 B.n294 585
R738 B.n293 B.n206 585
R739 B.n292 B.n291 585
R740 B.n290 B.n207 585
R741 B.n289 B.n288 585
R742 B.n287 B.n208 585
R743 B.n286 B.n285 585
R744 B.n284 B.n209 585
R745 B.n283 B.n282 585
R746 B.n281 B.n210 585
R747 B.n280 B.n279 585
R748 B.n278 B.n211 585
R749 B.n277 B.n276 585
R750 B.n275 B.n212 585
R751 B.n274 B.n273 585
R752 B.n272 B.n213 585
R753 B.n271 B.n270 585
R754 B.n269 B.n214 585
R755 B.n268 B.n267 585
R756 B.n266 B.n215 585
R757 B.n265 B.n264 585
R758 B.n263 B.n216 585
R759 B.n262 B.n261 585
R760 B.n260 B.n217 585
R761 B.n259 B.n258 585
R762 B.n257 B.n218 585
R763 B.n256 B.n255 585
R764 B.n254 B.n219 585
R765 B.n253 B.n252 585
R766 B.n251 B.n220 585
R767 B.n250 B.n249 585
R768 B.n248 B.n221 585
R769 B.n247 B.n246 585
R770 B.n245 B.n222 585
R771 B.n244 B.n243 585
R772 B.n242 B.n223 585
R773 B.n241 B.n240 585
R774 B.n239 B.n224 585
R775 B.n238 B.n237 585
R776 B.n236 B.n225 585
R777 B.n235 B.n234 585
R778 B.n233 B.n226 585
R779 B.n232 B.n231 585
R780 B.n230 B.n227 585
R781 B.n229 B.n228 585
R782 B.n2 B.n0 585
R783 B.n881 B.n1 585
R784 B.n880 B.n879 585
R785 B.n878 B.n3 585
R786 B.n877 B.n876 585
R787 B.n875 B.n4 585
R788 B.n874 B.n873 585
R789 B.n872 B.n5 585
R790 B.n871 B.n870 585
R791 B.n869 B.n6 585
R792 B.n868 B.n867 585
R793 B.n866 B.n7 585
R794 B.n865 B.n864 585
R795 B.n863 B.n8 585
R796 B.n862 B.n861 585
R797 B.n860 B.n9 585
R798 B.n859 B.n858 585
R799 B.n857 B.n10 585
R800 B.n856 B.n855 585
R801 B.n854 B.n11 585
R802 B.n853 B.n852 585
R803 B.n851 B.n12 585
R804 B.n850 B.n849 585
R805 B.n848 B.n13 585
R806 B.n847 B.n846 585
R807 B.n845 B.n14 585
R808 B.n844 B.n843 585
R809 B.n842 B.n15 585
R810 B.n841 B.n840 585
R811 B.n839 B.n16 585
R812 B.n838 B.n837 585
R813 B.n836 B.n17 585
R814 B.n835 B.n834 585
R815 B.n833 B.n18 585
R816 B.n832 B.n831 585
R817 B.n830 B.n19 585
R818 B.n829 B.n828 585
R819 B.n827 B.n20 585
R820 B.n826 B.n825 585
R821 B.n824 B.n21 585
R822 B.n823 B.n822 585
R823 B.n821 B.n22 585
R824 B.n820 B.n819 585
R825 B.n818 B.n23 585
R826 B.n817 B.n816 585
R827 B.n815 B.n24 585
R828 B.n814 B.n813 585
R829 B.n812 B.n25 585
R830 B.n811 B.n810 585
R831 B.n809 B.n26 585
R832 B.n808 B.n807 585
R833 B.n806 B.n27 585
R834 B.n805 B.n804 585
R835 B.n803 B.n28 585
R836 B.n802 B.n801 585
R837 B.n800 B.n29 585
R838 B.n799 B.n798 585
R839 B.n797 B.n30 585
R840 B.n796 B.n795 585
R841 B.n794 B.n31 585
R842 B.n793 B.n792 585
R843 B.n791 B.n32 585
R844 B.n790 B.n789 585
R845 B.n788 B.n33 585
R846 B.n787 B.n786 585
R847 B.n785 B.n34 585
R848 B.n784 B.n783 585
R849 B.n782 B.n35 585
R850 B.n781 B.n780 585
R851 B.n779 B.n36 585
R852 B.n778 B.n777 585
R853 B.n776 B.n37 585
R854 B.n775 B.n774 585
R855 B.n773 B.n38 585
R856 B.n772 B.n771 585
R857 B.n770 B.n39 585
R858 B.n883 B.n882 585
R859 B.n340 B.n191 492.5
R860 B.n768 B.n39 492.5
R861 B.n442 B.n153 492.5
R862 B.n666 B.n77 492.5
R863 B.n168 B.t6 262.558
R864 B.n174 B.t3 262.558
R865 B.n54 B.t9 262.558
R866 B.n62 B.t0 262.558
R867 B.n168 B.t8 185.75
R868 B.n62 B.t1 185.75
R869 B.n174 B.t5 185.743
R870 B.n54 B.t10 185.743
R871 B.n336 B.n191 163.367
R872 B.n336 B.n335 163.367
R873 B.n335 B.n334 163.367
R874 B.n334 B.n193 163.367
R875 B.n330 B.n193 163.367
R876 B.n330 B.n329 163.367
R877 B.n329 B.n328 163.367
R878 B.n328 B.n195 163.367
R879 B.n324 B.n195 163.367
R880 B.n324 B.n323 163.367
R881 B.n323 B.n322 163.367
R882 B.n322 B.n197 163.367
R883 B.n318 B.n197 163.367
R884 B.n318 B.n317 163.367
R885 B.n317 B.n316 163.367
R886 B.n316 B.n199 163.367
R887 B.n312 B.n199 163.367
R888 B.n312 B.n311 163.367
R889 B.n311 B.n310 163.367
R890 B.n310 B.n201 163.367
R891 B.n306 B.n201 163.367
R892 B.n306 B.n305 163.367
R893 B.n305 B.n304 163.367
R894 B.n304 B.n203 163.367
R895 B.n300 B.n203 163.367
R896 B.n300 B.n299 163.367
R897 B.n299 B.n298 163.367
R898 B.n298 B.n205 163.367
R899 B.n294 B.n205 163.367
R900 B.n294 B.n293 163.367
R901 B.n293 B.n292 163.367
R902 B.n292 B.n207 163.367
R903 B.n288 B.n207 163.367
R904 B.n288 B.n287 163.367
R905 B.n287 B.n286 163.367
R906 B.n286 B.n209 163.367
R907 B.n282 B.n209 163.367
R908 B.n282 B.n281 163.367
R909 B.n281 B.n280 163.367
R910 B.n280 B.n211 163.367
R911 B.n276 B.n211 163.367
R912 B.n276 B.n275 163.367
R913 B.n275 B.n274 163.367
R914 B.n274 B.n213 163.367
R915 B.n270 B.n213 163.367
R916 B.n270 B.n269 163.367
R917 B.n269 B.n268 163.367
R918 B.n268 B.n215 163.367
R919 B.n264 B.n215 163.367
R920 B.n264 B.n263 163.367
R921 B.n263 B.n262 163.367
R922 B.n262 B.n217 163.367
R923 B.n258 B.n217 163.367
R924 B.n258 B.n257 163.367
R925 B.n257 B.n256 163.367
R926 B.n256 B.n219 163.367
R927 B.n252 B.n219 163.367
R928 B.n252 B.n251 163.367
R929 B.n251 B.n250 163.367
R930 B.n250 B.n221 163.367
R931 B.n246 B.n221 163.367
R932 B.n246 B.n245 163.367
R933 B.n245 B.n244 163.367
R934 B.n244 B.n223 163.367
R935 B.n240 B.n223 163.367
R936 B.n240 B.n239 163.367
R937 B.n239 B.n238 163.367
R938 B.n238 B.n225 163.367
R939 B.n234 B.n225 163.367
R940 B.n234 B.n233 163.367
R941 B.n233 B.n232 163.367
R942 B.n232 B.n227 163.367
R943 B.n228 B.n227 163.367
R944 B.n228 B.n2 163.367
R945 B.n882 B.n2 163.367
R946 B.n882 B.n881 163.367
R947 B.n881 B.n880 163.367
R948 B.n880 B.n3 163.367
R949 B.n876 B.n3 163.367
R950 B.n876 B.n875 163.367
R951 B.n875 B.n874 163.367
R952 B.n874 B.n5 163.367
R953 B.n870 B.n5 163.367
R954 B.n870 B.n869 163.367
R955 B.n869 B.n868 163.367
R956 B.n868 B.n7 163.367
R957 B.n864 B.n7 163.367
R958 B.n864 B.n863 163.367
R959 B.n863 B.n862 163.367
R960 B.n862 B.n9 163.367
R961 B.n858 B.n9 163.367
R962 B.n858 B.n857 163.367
R963 B.n857 B.n856 163.367
R964 B.n856 B.n11 163.367
R965 B.n852 B.n11 163.367
R966 B.n852 B.n851 163.367
R967 B.n851 B.n850 163.367
R968 B.n850 B.n13 163.367
R969 B.n846 B.n13 163.367
R970 B.n846 B.n845 163.367
R971 B.n845 B.n844 163.367
R972 B.n844 B.n15 163.367
R973 B.n840 B.n15 163.367
R974 B.n840 B.n839 163.367
R975 B.n839 B.n838 163.367
R976 B.n838 B.n17 163.367
R977 B.n834 B.n17 163.367
R978 B.n834 B.n833 163.367
R979 B.n833 B.n832 163.367
R980 B.n832 B.n19 163.367
R981 B.n828 B.n19 163.367
R982 B.n828 B.n827 163.367
R983 B.n827 B.n826 163.367
R984 B.n826 B.n21 163.367
R985 B.n822 B.n21 163.367
R986 B.n822 B.n821 163.367
R987 B.n821 B.n820 163.367
R988 B.n820 B.n23 163.367
R989 B.n816 B.n23 163.367
R990 B.n816 B.n815 163.367
R991 B.n815 B.n814 163.367
R992 B.n814 B.n25 163.367
R993 B.n810 B.n25 163.367
R994 B.n810 B.n809 163.367
R995 B.n809 B.n808 163.367
R996 B.n808 B.n27 163.367
R997 B.n804 B.n27 163.367
R998 B.n804 B.n803 163.367
R999 B.n803 B.n802 163.367
R1000 B.n802 B.n29 163.367
R1001 B.n798 B.n29 163.367
R1002 B.n798 B.n797 163.367
R1003 B.n797 B.n796 163.367
R1004 B.n796 B.n31 163.367
R1005 B.n792 B.n31 163.367
R1006 B.n792 B.n791 163.367
R1007 B.n791 B.n790 163.367
R1008 B.n790 B.n33 163.367
R1009 B.n786 B.n33 163.367
R1010 B.n786 B.n785 163.367
R1011 B.n785 B.n784 163.367
R1012 B.n784 B.n35 163.367
R1013 B.n780 B.n35 163.367
R1014 B.n780 B.n779 163.367
R1015 B.n779 B.n778 163.367
R1016 B.n778 B.n37 163.367
R1017 B.n774 B.n37 163.367
R1018 B.n774 B.n773 163.367
R1019 B.n773 B.n772 163.367
R1020 B.n772 B.n39 163.367
R1021 B.n341 B.n340 163.367
R1022 B.n342 B.n341 163.367
R1023 B.n342 B.n189 163.367
R1024 B.n346 B.n189 163.367
R1025 B.n347 B.n346 163.367
R1026 B.n348 B.n347 163.367
R1027 B.n348 B.n187 163.367
R1028 B.n352 B.n187 163.367
R1029 B.n353 B.n352 163.367
R1030 B.n354 B.n353 163.367
R1031 B.n354 B.n185 163.367
R1032 B.n358 B.n185 163.367
R1033 B.n359 B.n358 163.367
R1034 B.n360 B.n359 163.367
R1035 B.n360 B.n183 163.367
R1036 B.n364 B.n183 163.367
R1037 B.n365 B.n364 163.367
R1038 B.n366 B.n365 163.367
R1039 B.n366 B.n181 163.367
R1040 B.n370 B.n181 163.367
R1041 B.n371 B.n370 163.367
R1042 B.n372 B.n371 163.367
R1043 B.n372 B.n179 163.367
R1044 B.n376 B.n179 163.367
R1045 B.n377 B.n376 163.367
R1046 B.n378 B.n377 163.367
R1047 B.n378 B.n177 163.367
R1048 B.n382 B.n177 163.367
R1049 B.n383 B.n382 163.367
R1050 B.n383 B.n173 163.367
R1051 B.n387 B.n173 163.367
R1052 B.n388 B.n387 163.367
R1053 B.n389 B.n388 163.367
R1054 B.n389 B.n171 163.367
R1055 B.n393 B.n171 163.367
R1056 B.n394 B.n393 163.367
R1057 B.n395 B.n394 163.367
R1058 B.n395 B.n167 163.367
R1059 B.n400 B.n167 163.367
R1060 B.n401 B.n400 163.367
R1061 B.n402 B.n401 163.367
R1062 B.n402 B.n165 163.367
R1063 B.n406 B.n165 163.367
R1064 B.n407 B.n406 163.367
R1065 B.n408 B.n407 163.367
R1066 B.n408 B.n163 163.367
R1067 B.n412 B.n163 163.367
R1068 B.n413 B.n412 163.367
R1069 B.n414 B.n413 163.367
R1070 B.n414 B.n161 163.367
R1071 B.n418 B.n161 163.367
R1072 B.n419 B.n418 163.367
R1073 B.n420 B.n419 163.367
R1074 B.n420 B.n159 163.367
R1075 B.n424 B.n159 163.367
R1076 B.n425 B.n424 163.367
R1077 B.n426 B.n425 163.367
R1078 B.n426 B.n157 163.367
R1079 B.n430 B.n157 163.367
R1080 B.n431 B.n430 163.367
R1081 B.n432 B.n431 163.367
R1082 B.n432 B.n155 163.367
R1083 B.n436 B.n155 163.367
R1084 B.n437 B.n436 163.367
R1085 B.n438 B.n437 163.367
R1086 B.n438 B.n153 163.367
R1087 B.n443 B.n442 163.367
R1088 B.n444 B.n443 163.367
R1089 B.n444 B.n151 163.367
R1090 B.n448 B.n151 163.367
R1091 B.n449 B.n448 163.367
R1092 B.n450 B.n449 163.367
R1093 B.n450 B.n149 163.367
R1094 B.n454 B.n149 163.367
R1095 B.n455 B.n454 163.367
R1096 B.n456 B.n455 163.367
R1097 B.n456 B.n147 163.367
R1098 B.n460 B.n147 163.367
R1099 B.n461 B.n460 163.367
R1100 B.n462 B.n461 163.367
R1101 B.n462 B.n145 163.367
R1102 B.n466 B.n145 163.367
R1103 B.n467 B.n466 163.367
R1104 B.n468 B.n467 163.367
R1105 B.n468 B.n143 163.367
R1106 B.n472 B.n143 163.367
R1107 B.n473 B.n472 163.367
R1108 B.n474 B.n473 163.367
R1109 B.n474 B.n141 163.367
R1110 B.n478 B.n141 163.367
R1111 B.n479 B.n478 163.367
R1112 B.n480 B.n479 163.367
R1113 B.n480 B.n139 163.367
R1114 B.n484 B.n139 163.367
R1115 B.n485 B.n484 163.367
R1116 B.n486 B.n485 163.367
R1117 B.n486 B.n137 163.367
R1118 B.n490 B.n137 163.367
R1119 B.n491 B.n490 163.367
R1120 B.n492 B.n491 163.367
R1121 B.n492 B.n135 163.367
R1122 B.n496 B.n135 163.367
R1123 B.n497 B.n496 163.367
R1124 B.n498 B.n497 163.367
R1125 B.n498 B.n133 163.367
R1126 B.n502 B.n133 163.367
R1127 B.n503 B.n502 163.367
R1128 B.n504 B.n503 163.367
R1129 B.n504 B.n131 163.367
R1130 B.n508 B.n131 163.367
R1131 B.n509 B.n508 163.367
R1132 B.n510 B.n509 163.367
R1133 B.n510 B.n129 163.367
R1134 B.n514 B.n129 163.367
R1135 B.n515 B.n514 163.367
R1136 B.n516 B.n515 163.367
R1137 B.n516 B.n127 163.367
R1138 B.n520 B.n127 163.367
R1139 B.n521 B.n520 163.367
R1140 B.n522 B.n521 163.367
R1141 B.n522 B.n125 163.367
R1142 B.n526 B.n125 163.367
R1143 B.n527 B.n526 163.367
R1144 B.n528 B.n527 163.367
R1145 B.n528 B.n123 163.367
R1146 B.n532 B.n123 163.367
R1147 B.n533 B.n532 163.367
R1148 B.n534 B.n533 163.367
R1149 B.n534 B.n121 163.367
R1150 B.n538 B.n121 163.367
R1151 B.n539 B.n538 163.367
R1152 B.n540 B.n539 163.367
R1153 B.n540 B.n119 163.367
R1154 B.n544 B.n119 163.367
R1155 B.n545 B.n544 163.367
R1156 B.n546 B.n545 163.367
R1157 B.n546 B.n117 163.367
R1158 B.n550 B.n117 163.367
R1159 B.n551 B.n550 163.367
R1160 B.n552 B.n551 163.367
R1161 B.n552 B.n115 163.367
R1162 B.n556 B.n115 163.367
R1163 B.n557 B.n556 163.367
R1164 B.n558 B.n557 163.367
R1165 B.n558 B.n113 163.367
R1166 B.n562 B.n113 163.367
R1167 B.n563 B.n562 163.367
R1168 B.n564 B.n563 163.367
R1169 B.n564 B.n111 163.367
R1170 B.n568 B.n111 163.367
R1171 B.n569 B.n568 163.367
R1172 B.n570 B.n569 163.367
R1173 B.n570 B.n109 163.367
R1174 B.n574 B.n109 163.367
R1175 B.n575 B.n574 163.367
R1176 B.n576 B.n575 163.367
R1177 B.n576 B.n107 163.367
R1178 B.n580 B.n107 163.367
R1179 B.n581 B.n580 163.367
R1180 B.n582 B.n581 163.367
R1181 B.n582 B.n105 163.367
R1182 B.n586 B.n105 163.367
R1183 B.n587 B.n586 163.367
R1184 B.n588 B.n587 163.367
R1185 B.n588 B.n103 163.367
R1186 B.n592 B.n103 163.367
R1187 B.n593 B.n592 163.367
R1188 B.n594 B.n593 163.367
R1189 B.n594 B.n101 163.367
R1190 B.n598 B.n101 163.367
R1191 B.n599 B.n598 163.367
R1192 B.n600 B.n599 163.367
R1193 B.n600 B.n99 163.367
R1194 B.n604 B.n99 163.367
R1195 B.n605 B.n604 163.367
R1196 B.n606 B.n605 163.367
R1197 B.n606 B.n97 163.367
R1198 B.n610 B.n97 163.367
R1199 B.n611 B.n610 163.367
R1200 B.n612 B.n611 163.367
R1201 B.n612 B.n95 163.367
R1202 B.n616 B.n95 163.367
R1203 B.n617 B.n616 163.367
R1204 B.n618 B.n617 163.367
R1205 B.n618 B.n93 163.367
R1206 B.n622 B.n93 163.367
R1207 B.n623 B.n622 163.367
R1208 B.n624 B.n623 163.367
R1209 B.n624 B.n91 163.367
R1210 B.n628 B.n91 163.367
R1211 B.n629 B.n628 163.367
R1212 B.n630 B.n629 163.367
R1213 B.n630 B.n89 163.367
R1214 B.n634 B.n89 163.367
R1215 B.n635 B.n634 163.367
R1216 B.n636 B.n635 163.367
R1217 B.n636 B.n87 163.367
R1218 B.n640 B.n87 163.367
R1219 B.n641 B.n640 163.367
R1220 B.n642 B.n641 163.367
R1221 B.n642 B.n85 163.367
R1222 B.n646 B.n85 163.367
R1223 B.n647 B.n646 163.367
R1224 B.n648 B.n647 163.367
R1225 B.n648 B.n83 163.367
R1226 B.n652 B.n83 163.367
R1227 B.n653 B.n652 163.367
R1228 B.n654 B.n653 163.367
R1229 B.n654 B.n81 163.367
R1230 B.n658 B.n81 163.367
R1231 B.n659 B.n658 163.367
R1232 B.n660 B.n659 163.367
R1233 B.n660 B.n79 163.367
R1234 B.n664 B.n79 163.367
R1235 B.n665 B.n664 163.367
R1236 B.n666 B.n665 163.367
R1237 B.n768 B.n767 163.367
R1238 B.n767 B.n766 163.367
R1239 B.n766 B.n41 163.367
R1240 B.n762 B.n41 163.367
R1241 B.n762 B.n761 163.367
R1242 B.n761 B.n760 163.367
R1243 B.n760 B.n43 163.367
R1244 B.n756 B.n43 163.367
R1245 B.n756 B.n755 163.367
R1246 B.n755 B.n754 163.367
R1247 B.n754 B.n45 163.367
R1248 B.n750 B.n45 163.367
R1249 B.n750 B.n749 163.367
R1250 B.n749 B.n748 163.367
R1251 B.n748 B.n47 163.367
R1252 B.n744 B.n47 163.367
R1253 B.n744 B.n743 163.367
R1254 B.n743 B.n742 163.367
R1255 B.n742 B.n49 163.367
R1256 B.n738 B.n49 163.367
R1257 B.n738 B.n737 163.367
R1258 B.n737 B.n736 163.367
R1259 B.n736 B.n51 163.367
R1260 B.n732 B.n51 163.367
R1261 B.n732 B.n731 163.367
R1262 B.n731 B.n730 163.367
R1263 B.n730 B.n53 163.367
R1264 B.n726 B.n53 163.367
R1265 B.n726 B.n725 163.367
R1266 B.n725 B.n57 163.367
R1267 B.n721 B.n57 163.367
R1268 B.n721 B.n720 163.367
R1269 B.n720 B.n719 163.367
R1270 B.n719 B.n59 163.367
R1271 B.n715 B.n59 163.367
R1272 B.n715 B.n714 163.367
R1273 B.n714 B.n713 163.367
R1274 B.n713 B.n61 163.367
R1275 B.n708 B.n61 163.367
R1276 B.n708 B.n707 163.367
R1277 B.n707 B.n706 163.367
R1278 B.n706 B.n65 163.367
R1279 B.n702 B.n65 163.367
R1280 B.n702 B.n701 163.367
R1281 B.n701 B.n700 163.367
R1282 B.n700 B.n67 163.367
R1283 B.n696 B.n67 163.367
R1284 B.n696 B.n695 163.367
R1285 B.n695 B.n694 163.367
R1286 B.n694 B.n69 163.367
R1287 B.n690 B.n69 163.367
R1288 B.n690 B.n689 163.367
R1289 B.n689 B.n688 163.367
R1290 B.n688 B.n71 163.367
R1291 B.n684 B.n71 163.367
R1292 B.n684 B.n683 163.367
R1293 B.n683 B.n682 163.367
R1294 B.n682 B.n73 163.367
R1295 B.n678 B.n73 163.367
R1296 B.n678 B.n677 163.367
R1297 B.n677 B.n676 163.367
R1298 B.n676 B.n75 163.367
R1299 B.n672 B.n75 163.367
R1300 B.n672 B.n671 163.367
R1301 B.n671 B.n670 163.367
R1302 B.n670 B.n77 163.367
R1303 B.n169 B.t7 112.442
R1304 B.n63 B.t2 112.442
R1305 B.n175 B.t4 112.433
R1306 B.n55 B.t11 112.433
R1307 B.n169 B.n168 73.3096
R1308 B.n175 B.n174 73.3096
R1309 B.n55 B.n54 73.3096
R1310 B.n63 B.n62 73.3096
R1311 B.n397 B.n169 59.5399
R1312 B.n176 B.n175 59.5399
R1313 B.n56 B.n55 59.5399
R1314 B.n711 B.n63 59.5399
R1315 B.n770 B.n769 32.0005
R1316 B.n668 B.n667 32.0005
R1317 B.n441 B.n440 32.0005
R1318 B.n339 B.n338 32.0005
R1319 B B.n883 18.0485
R1320 B.n769 B.n40 10.6151
R1321 B.n765 B.n40 10.6151
R1322 B.n765 B.n764 10.6151
R1323 B.n764 B.n763 10.6151
R1324 B.n763 B.n42 10.6151
R1325 B.n759 B.n42 10.6151
R1326 B.n759 B.n758 10.6151
R1327 B.n758 B.n757 10.6151
R1328 B.n757 B.n44 10.6151
R1329 B.n753 B.n44 10.6151
R1330 B.n753 B.n752 10.6151
R1331 B.n752 B.n751 10.6151
R1332 B.n751 B.n46 10.6151
R1333 B.n747 B.n46 10.6151
R1334 B.n747 B.n746 10.6151
R1335 B.n746 B.n745 10.6151
R1336 B.n745 B.n48 10.6151
R1337 B.n741 B.n48 10.6151
R1338 B.n741 B.n740 10.6151
R1339 B.n740 B.n739 10.6151
R1340 B.n739 B.n50 10.6151
R1341 B.n735 B.n50 10.6151
R1342 B.n735 B.n734 10.6151
R1343 B.n734 B.n733 10.6151
R1344 B.n733 B.n52 10.6151
R1345 B.n729 B.n52 10.6151
R1346 B.n729 B.n728 10.6151
R1347 B.n728 B.n727 10.6151
R1348 B.n724 B.n723 10.6151
R1349 B.n723 B.n722 10.6151
R1350 B.n722 B.n58 10.6151
R1351 B.n718 B.n58 10.6151
R1352 B.n718 B.n717 10.6151
R1353 B.n717 B.n716 10.6151
R1354 B.n716 B.n60 10.6151
R1355 B.n712 B.n60 10.6151
R1356 B.n710 B.n709 10.6151
R1357 B.n709 B.n64 10.6151
R1358 B.n705 B.n64 10.6151
R1359 B.n705 B.n704 10.6151
R1360 B.n704 B.n703 10.6151
R1361 B.n703 B.n66 10.6151
R1362 B.n699 B.n66 10.6151
R1363 B.n699 B.n698 10.6151
R1364 B.n698 B.n697 10.6151
R1365 B.n697 B.n68 10.6151
R1366 B.n693 B.n68 10.6151
R1367 B.n693 B.n692 10.6151
R1368 B.n692 B.n691 10.6151
R1369 B.n691 B.n70 10.6151
R1370 B.n687 B.n70 10.6151
R1371 B.n687 B.n686 10.6151
R1372 B.n686 B.n685 10.6151
R1373 B.n685 B.n72 10.6151
R1374 B.n681 B.n72 10.6151
R1375 B.n681 B.n680 10.6151
R1376 B.n680 B.n679 10.6151
R1377 B.n679 B.n74 10.6151
R1378 B.n675 B.n74 10.6151
R1379 B.n675 B.n674 10.6151
R1380 B.n674 B.n673 10.6151
R1381 B.n673 B.n76 10.6151
R1382 B.n669 B.n76 10.6151
R1383 B.n669 B.n668 10.6151
R1384 B.n441 B.n152 10.6151
R1385 B.n445 B.n152 10.6151
R1386 B.n446 B.n445 10.6151
R1387 B.n447 B.n446 10.6151
R1388 B.n447 B.n150 10.6151
R1389 B.n451 B.n150 10.6151
R1390 B.n452 B.n451 10.6151
R1391 B.n453 B.n452 10.6151
R1392 B.n453 B.n148 10.6151
R1393 B.n457 B.n148 10.6151
R1394 B.n458 B.n457 10.6151
R1395 B.n459 B.n458 10.6151
R1396 B.n459 B.n146 10.6151
R1397 B.n463 B.n146 10.6151
R1398 B.n464 B.n463 10.6151
R1399 B.n465 B.n464 10.6151
R1400 B.n465 B.n144 10.6151
R1401 B.n469 B.n144 10.6151
R1402 B.n470 B.n469 10.6151
R1403 B.n471 B.n470 10.6151
R1404 B.n471 B.n142 10.6151
R1405 B.n475 B.n142 10.6151
R1406 B.n476 B.n475 10.6151
R1407 B.n477 B.n476 10.6151
R1408 B.n477 B.n140 10.6151
R1409 B.n481 B.n140 10.6151
R1410 B.n482 B.n481 10.6151
R1411 B.n483 B.n482 10.6151
R1412 B.n483 B.n138 10.6151
R1413 B.n487 B.n138 10.6151
R1414 B.n488 B.n487 10.6151
R1415 B.n489 B.n488 10.6151
R1416 B.n489 B.n136 10.6151
R1417 B.n493 B.n136 10.6151
R1418 B.n494 B.n493 10.6151
R1419 B.n495 B.n494 10.6151
R1420 B.n495 B.n134 10.6151
R1421 B.n499 B.n134 10.6151
R1422 B.n500 B.n499 10.6151
R1423 B.n501 B.n500 10.6151
R1424 B.n501 B.n132 10.6151
R1425 B.n505 B.n132 10.6151
R1426 B.n506 B.n505 10.6151
R1427 B.n507 B.n506 10.6151
R1428 B.n507 B.n130 10.6151
R1429 B.n511 B.n130 10.6151
R1430 B.n512 B.n511 10.6151
R1431 B.n513 B.n512 10.6151
R1432 B.n513 B.n128 10.6151
R1433 B.n517 B.n128 10.6151
R1434 B.n518 B.n517 10.6151
R1435 B.n519 B.n518 10.6151
R1436 B.n519 B.n126 10.6151
R1437 B.n523 B.n126 10.6151
R1438 B.n524 B.n523 10.6151
R1439 B.n525 B.n524 10.6151
R1440 B.n525 B.n124 10.6151
R1441 B.n529 B.n124 10.6151
R1442 B.n530 B.n529 10.6151
R1443 B.n531 B.n530 10.6151
R1444 B.n531 B.n122 10.6151
R1445 B.n535 B.n122 10.6151
R1446 B.n536 B.n535 10.6151
R1447 B.n537 B.n536 10.6151
R1448 B.n537 B.n120 10.6151
R1449 B.n541 B.n120 10.6151
R1450 B.n542 B.n541 10.6151
R1451 B.n543 B.n542 10.6151
R1452 B.n543 B.n118 10.6151
R1453 B.n547 B.n118 10.6151
R1454 B.n548 B.n547 10.6151
R1455 B.n549 B.n548 10.6151
R1456 B.n549 B.n116 10.6151
R1457 B.n553 B.n116 10.6151
R1458 B.n554 B.n553 10.6151
R1459 B.n555 B.n554 10.6151
R1460 B.n555 B.n114 10.6151
R1461 B.n559 B.n114 10.6151
R1462 B.n560 B.n559 10.6151
R1463 B.n561 B.n560 10.6151
R1464 B.n561 B.n112 10.6151
R1465 B.n565 B.n112 10.6151
R1466 B.n566 B.n565 10.6151
R1467 B.n567 B.n566 10.6151
R1468 B.n567 B.n110 10.6151
R1469 B.n571 B.n110 10.6151
R1470 B.n572 B.n571 10.6151
R1471 B.n573 B.n572 10.6151
R1472 B.n573 B.n108 10.6151
R1473 B.n577 B.n108 10.6151
R1474 B.n578 B.n577 10.6151
R1475 B.n579 B.n578 10.6151
R1476 B.n579 B.n106 10.6151
R1477 B.n583 B.n106 10.6151
R1478 B.n584 B.n583 10.6151
R1479 B.n585 B.n584 10.6151
R1480 B.n585 B.n104 10.6151
R1481 B.n589 B.n104 10.6151
R1482 B.n590 B.n589 10.6151
R1483 B.n591 B.n590 10.6151
R1484 B.n591 B.n102 10.6151
R1485 B.n595 B.n102 10.6151
R1486 B.n596 B.n595 10.6151
R1487 B.n597 B.n596 10.6151
R1488 B.n597 B.n100 10.6151
R1489 B.n601 B.n100 10.6151
R1490 B.n602 B.n601 10.6151
R1491 B.n603 B.n602 10.6151
R1492 B.n603 B.n98 10.6151
R1493 B.n607 B.n98 10.6151
R1494 B.n608 B.n607 10.6151
R1495 B.n609 B.n608 10.6151
R1496 B.n609 B.n96 10.6151
R1497 B.n613 B.n96 10.6151
R1498 B.n614 B.n613 10.6151
R1499 B.n615 B.n614 10.6151
R1500 B.n615 B.n94 10.6151
R1501 B.n619 B.n94 10.6151
R1502 B.n620 B.n619 10.6151
R1503 B.n621 B.n620 10.6151
R1504 B.n621 B.n92 10.6151
R1505 B.n625 B.n92 10.6151
R1506 B.n626 B.n625 10.6151
R1507 B.n627 B.n626 10.6151
R1508 B.n627 B.n90 10.6151
R1509 B.n631 B.n90 10.6151
R1510 B.n632 B.n631 10.6151
R1511 B.n633 B.n632 10.6151
R1512 B.n633 B.n88 10.6151
R1513 B.n637 B.n88 10.6151
R1514 B.n638 B.n637 10.6151
R1515 B.n639 B.n638 10.6151
R1516 B.n639 B.n86 10.6151
R1517 B.n643 B.n86 10.6151
R1518 B.n644 B.n643 10.6151
R1519 B.n645 B.n644 10.6151
R1520 B.n645 B.n84 10.6151
R1521 B.n649 B.n84 10.6151
R1522 B.n650 B.n649 10.6151
R1523 B.n651 B.n650 10.6151
R1524 B.n651 B.n82 10.6151
R1525 B.n655 B.n82 10.6151
R1526 B.n656 B.n655 10.6151
R1527 B.n657 B.n656 10.6151
R1528 B.n657 B.n80 10.6151
R1529 B.n661 B.n80 10.6151
R1530 B.n662 B.n661 10.6151
R1531 B.n663 B.n662 10.6151
R1532 B.n663 B.n78 10.6151
R1533 B.n667 B.n78 10.6151
R1534 B.n339 B.n190 10.6151
R1535 B.n343 B.n190 10.6151
R1536 B.n344 B.n343 10.6151
R1537 B.n345 B.n344 10.6151
R1538 B.n345 B.n188 10.6151
R1539 B.n349 B.n188 10.6151
R1540 B.n350 B.n349 10.6151
R1541 B.n351 B.n350 10.6151
R1542 B.n351 B.n186 10.6151
R1543 B.n355 B.n186 10.6151
R1544 B.n356 B.n355 10.6151
R1545 B.n357 B.n356 10.6151
R1546 B.n357 B.n184 10.6151
R1547 B.n361 B.n184 10.6151
R1548 B.n362 B.n361 10.6151
R1549 B.n363 B.n362 10.6151
R1550 B.n363 B.n182 10.6151
R1551 B.n367 B.n182 10.6151
R1552 B.n368 B.n367 10.6151
R1553 B.n369 B.n368 10.6151
R1554 B.n369 B.n180 10.6151
R1555 B.n373 B.n180 10.6151
R1556 B.n374 B.n373 10.6151
R1557 B.n375 B.n374 10.6151
R1558 B.n375 B.n178 10.6151
R1559 B.n379 B.n178 10.6151
R1560 B.n380 B.n379 10.6151
R1561 B.n381 B.n380 10.6151
R1562 B.n385 B.n384 10.6151
R1563 B.n386 B.n385 10.6151
R1564 B.n386 B.n172 10.6151
R1565 B.n390 B.n172 10.6151
R1566 B.n391 B.n390 10.6151
R1567 B.n392 B.n391 10.6151
R1568 B.n392 B.n170 10.6151
R1569 B.n396 B.n170 10.6151
R1570 B.n399 B.n398 10.6151
R1571 B.n399 B.n166 10.6151
R1572 B.n403 B.n166 10.6151
R1573 B.n404 B.n403 10.6151
R1574 B.n405 B.n404 10.6151
R1575 B.n405 B.n164 10.6151
R1576 B.n409 B.n164 10.6151
R1577 B.n410 B.n409 10.6151
R1578 B.n411 B.n410 10.6151
R1579 B.n411 B.n162 10.6151
R1580 B.n415 B.n162 10.6151
R1581 B.n416 B.n415 10.6151
R1582 B.n417 B.n416 10.6151
R1583 B.n417 B.n160 10.6151
R1584 B.n421 B.n160 10.6151
R1585 B.n422 B.n421 10.6151
R1586 B.n423 B.n422 10.6151
R1587 B.n423 B.n158 10.6151
R1588 B.n427 B.n158 10.6151
R1589 B.n428 B.n427 10.6151
R1590 B.n429 B.n428 10.6151
R1591 B.n429 B.n156 10.6151
R1592 B.n433 B.n156 10.6151
R1593 B.n434 B.n433 10.6151
R1594 B.n435 B.n434 10.6151
R1595 B.n435 B.n154 10.6151
R1596 B.n439 B.n154 10.6151
R1597 B.n440 B.n439 10.6151
R1598 B.n338 B.n337 10.6151
R1599 B.n337 B.n192 10.6151
R1600 B.n333 B.n192 10.6151
R1601 B.n333 B.n332 10.6151
R1602 B.n332 B.n331 10.6151
R1603 B.n331 B.n194 10.6151
R1604 B.n327 B.n194 10.6151
R1605 B.n327 B.n326 10.6151
R1606 B.n326 B.n325 10.6151
R1607 B.n325 B.n196 10.6151
R1608 B.n321 B.n196 10.6151
R1609 B.n321 B.n320 10.6151
R1610 B.n320 B.n319 10.6151
R1611 B.n319 B.n198 10.6151
R1612 B.n315 B.n198 10.6151
R1613 B.n315 B.n314 10.6151
R1614 B.n314 B.n313 10.6151
R1615 B.n313 B.n200 10.6151
R1616 B.n309 B.n200 10.6151
R1617 B.n309 B.n308 10.6151
R1618 B.n308 B.n307 10.6151
R1619 B.n307 B.n202 10.6151
R1620 B.n303 B.n202 10.6151
R1621 B.n303 B.n302 10.6151
R1622 B.n302 B.n301 10.6151
R1623 B.n301 B.n204 10.6151
R1624 B.n297 B.n204 10.6151
R1625 B.n297 B.n296 10.6151
R1626 B.n296 B.n295 10.6151
R1627 B.n295 B.n206 10.6151
R1628 B.n291 B.n206 10.6151
R1629 B.n291 B.n290 10.6151
R1630 B.n290 B.n289 10.6151
R1631 B.n289 B.n208 10.6151
R1632 B.n285 B.n208 10.6151
R1633 B.n285 B.n284 10.6151
R1634 B.n284 B.n283 10.6151
R1635 B.n283 B.n210 10.6151
R1636 B.n279 B.n210 10.6151
R1637 B.n279 B.n278 10.6151
R1638 B.n278 B.n277 10.6151
R1639 B.n277 B.n212 10.6151
R1640 B.n273 B.n212 10.6151
R1641 B.n273 B.n272 10.6151
R1642 B.n272 B.n271 10.6151
R1643 B.n271 B.n214 10.6151
R1644 B.n267 B.n214 10.6151
R1645 B.n267 B.n266 10.6151
R1646 B.n266 B.n265 10.6151
R1647 B.n265 B.n216 10.6151
R1648 B.n261 B.n216 10.6151
R1649 B.n261 B.n260 10.6151
R1650 B.n260 B.n259 10.6151
R1651 B.n259 B.n218 10.6151
R1652 B.n255 B.n218 10.6151
R1653 B.n255 B.n254 10.6151
R1654 B.n254 B.n253 10.6151
R1655 B.n253 B.n220 10.6151
R1656 B.n249 B.n220 10.6151
R1657 B.n249 B.n248 10.6151
R1658 B.n248 B.n247 10.6151
R1659 B.n247 B.n222 10.6151
R1660 B.n243 B.n222 10.6151
R1661 B.n243 B.n242 10.6151
R1662 B.n242 B.n241 10.6151
R1663 B.n241 B.n224 10.6151
R1664 B.n237 B.n224 10.6151
R1665 B.n237 B.n236 10.6151
R1666 B.n236 B.n235 10.6151
R1667 B.n235 B.n226 10.6151
R1668 B.n231 B.n226 10.6151
R1669 B.n231 B.n230 10.6151
R1670 B.n230 B.n229 10.6151
R1671 B.n229 B.n0 10.6151
R1672 B.n879 B.n1 10.6151
R1673 B.n879 B.n878 10.6151
R1674 B.n878 B.n877 10.6151
R1675 B.n877 B.n4 10.6151
R1676 B.n873 B.n4 10.6151
R1677 B.n873 B.n872 10.6151
R1678 B.n872 B.n871 10.6151
R1679 B.n871 B.n6 10.6151
R1680 B.n867 B.n6 10.6151
R1681 B.n867 B.n866 10.6151
R1682 B.n866 B.n865 10.6151
R1683 B.n865 B.n8 10.6151
R1684 B.n861 B.n8 10.6151
R1685 B.n861 B.n860 10.6151
R1686 B.n860 B.n859 10.6151
R1687 B.n859 B.n10 10.6151
R1688 B.n855 B.n10 10.6151
R1689 B.n855 B.n854 10.6151
R1690 B.n854 B.n853 10.6151
R1691 B.n853 B.n12 10.6151
R1692 B.n849 B.n12 10.6151
R1693 B.n849 B.n848 10.6151
R1694 B.n848 B.n847 10.6151
R1695 B.n847 B.n14 10.6151
R1696 B.n843 B.n14 10.6151
R1697 B.n843 B.n842 10.6151
R1698 B.n842 B.n841 10.6151
R1699 B.n841 B.n16 10.6151
R1700 B.n837 B.n16 10.6151
R1701 B.n837 B.n836 10.6151
R1702 B.n836 B.n835 10.6151
R1703 B.n835 B.n18 10.6151
R1704 B.n831 B.n18 10.6151
R1705 B.n831 B.n830 10.6151
R1706 B.n830 B.n829 10.6151
R1707 B.n829 B.n20 10.6151
R1708 B.n825 B.n20 10.6151
R1709 B.n825 B.n824 10.6151
R1710 B.n824 B.n823 10.6151
R1711 B.n823 B.n22 10.6151
R1712 B.n819 B.n22 10.6151
R1713 B.n819 B.n818 10.6151
R1714 B.n818 B.n817 10.6151
R1715 B.n817 B.n24 10.6151
R1716 B.n813 B.n24 10.6151
R1717 B.n813 B.n812 10.6151
R1718 B.n812 B.n811 10.6151
R1719 B.n811 B.n26 10.6151
R1720 B.n807 B.n26 10.6151
R1721 B.n807 B.n806 10.6151
R1722 B.n806 B.n805 10.6151
R1723 B.n805 B.n28 10.6151
R1724 B.n801 B.n28 10.6151
R1725 B.n801 B.n800 10.6151
R1726 B.n800 B.n799 10.6151
R1727 B.n799 B.n30 10.6151
R1728 B.n795 B.n30 10.6151
R1729 B.n795 B.n794 10.6151
R1730 B.n794 B.n793 10.6151
R1731 B.n793 B.n32 10.6151
R1732 B.n789 B.n32 10.6151
R1733 B.n789 B.n788 10.6151
R1734 B.n788 B.n787 10.6151
R1735 B.n787 B.n34 10.6151
R1736 B.n783 B.n34 10.6151
R1737 B.n783 B.n782 10.6151
R1738 B.n782 B.n781 10.6151
R1739 B.n781 B.n36 10.6151
R1740 B.n777 B.n36 10.6151
R1741 B.n777 B.n776 10.6151
R1742 B.n776 B.n775 10.6151
R1743 B.n775 B.n38 10.6151
R1744 B.n771 B.n38 10.6151
R1745 B.n771 B.n770 10.6151
R1746 B.n724 B.n56 6.5566
R1747 B.n712 B.n711 6.5566
R1748 B.n384 B.n176 6.5566
R1749 B.n397 B.n396 6.5566
R1750 B.n727 B.n56 4.05904
R1751 B.n711 B.n710 4.05904
R1752 B.n381 B.n176 4.05904
R1753 B.n398 B.n397 4.05904
R1754 B.n883 B.n0 2.81026
R1755 B.n883 B.n1 2.81026
C0 VTAIL VDD2 9.076071f
C1 VTAIL B 3.03779f
C2 VDD2 w_n5506_n2500# 3.00118f
C3 VN VDD2 7.35244f
C4 w_n5506_n2500# B 10.759f
C5 VN B 1.45314f
C6 VTAIL w_n5506_n2500# 2.74257f
C7 VN VTAIL 8.56312f
C8 VP VDD1 7.88556f
C9 VN w_n5506_n2500# 11.932799f
C10 VP VDD2 0.692053f
C11 VP B 2.66767f
C12 VDD2 VDD1 2.72746f
C13 VTAIL VP 8.577299f
C14 VDD1 B 2.46242f
C15 VP w_n5506_n2500# 12.6523f
C16 VN VP 8.83781f
C17 VTAIL VDD1 9.017941f
C18 VDD1 w_n5506_n2500# 2.81345f
C19 VN VDD1 0.155598f
C20 VDD2 B 2.61344f
C21 VDD2 VSUBS 2.424349f
C22 VDD1 VSUBS 2.215378f
C23 VTAIL VSUBS 1.374189f
C24 VN VSUBS 9.093731f
C25 VP VSUBS 5.177292f
C26 B VSUBS 6.055258f
C27 w_n5506_n2500# VSUBS 0.170928p
C28 B.n0 VSUBS 0.006731f
C29 B.n1 VSUBS 0.006731f
C30 B.n2 VSUBS 0.010644f
C31 B.n3 VSUBS 0.010644f
C32 B.n4 VSUBS 0.010644f
C33 B.n5 VSUBS 0.010644f
C34 B.n6 VSUBS 0.010644f
C35 B.n7 VSUBS 0.010644f
C36 B.n8 VSUBS 0.010644f
C37 B.n9 VSUBS 0.010644f
C38 B.n10 VSUBS 0.010644f
C39 B.n11 VSUBS 0.010644f
C40 B.n12 VSUBS 0.010644f
C41 B.n13 VSUBS 0.010644f
C42 B.n14 VSUBS 0.010644f
C43 B.n15 VSUBS 0.010644f
C44 B.n16 VSUBS 0.010644f
C45 B.n17 VSUBS 0.010644f
C46 B.n18 VSUBS 0.010644f
C47 B.n19 VSUBS 0.010644f
C48 B.n20 VSUBS 0.010644f
C49 B.n21 VSUBS 0.010644f
C50 B.n22 VSUBS 0.010644f
C51 B.n23 VSUBS 0.010644f
C52 B.n24 VSUBS 0.010644f
C53 B.n25 VSUBS 0.010644f
C54 B.n26 VSUBS 0.010644f
C55 B.n27 VSUBS 0.010644f
C56 B.n28 VSUBS 0.010644f
C57 B.n29 VSUBS 0.010644f
C58 B.n30 VSUBS 0.010644f
C59 B.n31 VSUBS 0.010644f
C60 B.n32 VSUBS 0.010644f
C61 B.n33 VSUBS 0.010644f
C62 B.n34 VSUBS 0.010644f
C63 B.n35 VSUBS 0.010644f
C64 B.n36 VSUBS 0.010644f
C65 B.n37 VSUBS 0.010644f
C66 B.n38 VSUBS 0.010644f
C67 B.n39 VSUBS 0.024309f
C68 B.n40 VSUBS 0.010644f
C69 B.n41 VSUBS 0.010644f
C70 B.n42 VSUBS 0.010644f
C71 B.n43 VSUBS 0.010644f
C72 B.n44 VSUBS 0.010644f
C73 B.n45 VSUBS 0.010644f
C74 B.n46 VSUBS 0.010644f
C75 B.n47 VSUBS 0.010644f
C76 B.n48 VSUBS 0.010644f
C77 B.n49 VSUBS 0.010644f
C78 B.n50 VSUBS 0.010644f
C79 B.n51 VSUBS 0.010644f
C80 B.n52 VSUBS 0.010644f
C81 B.n53 VSUBS 0.010644f
C82 B.t11 VSUBS 0.356731f
C83 B.t10 VSUBS 0.395669f
C84 B.t9 VSUBS 1.90543f
C85 B.n54 VSUBS 0.228091f
C86 B.n55 VSUBS 0.113839f
C87 B.n56 VSUBS 0.024661f
C88 B.n57 VSUBS 0.010644f
C89 B.n58 VSUBS 0.010644f
C90 B.n59 VSUBS 0.010644f
C91 B.n60 VSUBS 0.010644f
C92 B.n61 VSUBS 0.010644f
C93 B.t2 VSUBS 0.356728f
C94 B.t1 VSUBS 0.395666f
C95 B.t0 VSUBS 1.90543f
C96 B.n62 VSUBS 0.228095f
C97 B.n63 VSUBS 0.113841f
C98 B.n64 VSUBS 0.010644f
C99 B.n65 VSUBS 0.010644f
C100 B.n66 VSUBS 0.010644f
C101 B.n67 VSUBS 0.010644f
C102 B.n68 VSUBS 0.010644f
C103 B.n69 VSUBS 0.010644f
C104 B.n70 VSUBS 0.010644f
C105 B.n71 VSUBS 0.010644f
C106 B.n72 VSUBS 0.010644f
C107 B.n73 VSUBS 0.010644f
C108 B.n74 VSUBS 0.010644f
C109 B.n75 VSUBS 0.010644f
C110 B.n76 VSUBS 0.010644f
C111 B.n77 VSUBS 0.024841f
C112 B.n78 VSUBS 0.010644f
C113 B.n79 VSUBS 0.010644f
C114 B.n80 VSUBS 0.010644f
C115 B.n81 VSUBS 0.010644f
C116 B.n82 VSUBS 0.010644f
C117 B.n83 VSUBS 0.010644f
C118 B.n84 VSUBS 0.010644f
C119 B.n85 VSUBS 0.010644f
C120 B.n86 VSUBS 0.010644f
C121 B.n87 VSUBS 0.010644f
C122 B.n88 VSUBS 0.010644f
C123 B.n89 VSUBS 0.010644f
C124 B.n90 VSUBS 0.010644f
C125 B.n91 VSUBS 0.010644f
C126 B.n92 VSUBS 0.010644f
C127 B.n93 VSUBS 0.010644f
C128 B.n94 VSUBS 0.010644f
C129 B.n95 VSUBS 0.010644f
C130 B.n96 VSUBS 0.010644f
C131 B.n97 VSUBS 0.010644f
C132 B.n98 VSUBS 0.010644f
C133 B.n99 VSUBS 0.010644f
C134 B.n100 VSUBS 0.010644f
C135 B.n101 VSUBS 0.010644f
C136 B.n102 VSUBS 0.010644f
C137 B.n103 VSUBS 0.010644f
C138 B.n104 VSUBS 0.010644f
C139 B.n105 VSUBS 0.010644f
C140 B.n106 VSUBS 0.010644f
C141 B.n107 VSUBS 0.010644f
C142 B.n108 VSUBS 0.010644f
C143 B.n109 VSUBS 0.010644f
C144 B.n110 VSUBS 0.010644f
C145 B.n111 VSUBS 0.010644f
C146 B.n112 VSUBS 0.010644f
C147 B.n113 VSUBS 0.010644f
C148 B.n114 VSUBS 0.010644f
C149 B.n115 VSUBS 0.010644f
C150 B.n116 VSUBS 0.010644f
C151 B.n117 VSUBS 0.010644f
C152 B.n118 VSUBS 0.010644f
C153 B.n119 VSUBS 0.010644f
C154 B.n120 VSUBS 0.010644f
C155 B.n121 VSUBS 0.010644f
C156 B.n122 VSUBS 0.010644f
C157 B.n123 VSUBS 0.010644f
C158 B.n124 VSUBS 0.010644f
C159 B.n125 VSUBS 0.010644f
C160 B.n126 VSUBS 0.010644f
C161 B.n127 VSUBS 0.010644f
C162 B.n128 VSUBS 0.010644f
C163 B.n129 VSUBS 0.010644f
C164 B.n130 VSUBS 0.010644f
C165 B.n131 VSUBS 0.010644f
C166 B.n132 VSUBS 0.010644f
C167 B.n133 VSUBS 0.010644f
C168 B.n134 VSUBS 0.010644f
C169 B.n135 VSUBS 0.010644f
C170 B.n136 VSUBS 0.010644f
C171 B.n137 VSUBS 0.010644f
C172 B.n138 VSUBS 0.010644f
C173 B.n139 VSUBS 0.010644f
C174 B.n140 VSUBS 0.010644f
C175 B.n141 VSUBS 0.010644f
C176 B.n142 VSUBS 0.010644f
C177 B.n143 VSUBS 0.010644f
C178 B.n144 VSUBS 0.010644f
C179 B.n145 VSUBS 0.010644f
C180 B.n146 VSUBS 0.010644f
C181 B.n147 VSUBS 0.010644f
C182 B.n148 VSUBS 0.010644f
C183 B.n149 VSUBS 0.010644f
C184 B.n150 VSUBS 0.010644f
C185 B.n151 VSUBS 0.010644f
C186 B.n152 VSUBS 0.010644f
C187 B.n153 VSUBS 0.024841f
C188 B.n154 VSUBS 0.010644f
C189 B.n155 VSUBS 0.010644f
C190 B.n156 VSUBS 0.010644f
C191 B.n157 VSUBS 0.010644f
C192 B.n158 VSUBS 0.010644f
C193 B.n159 VSUBS 0.010644f
C194 B.n160 VSUBS 0.010644f
C195 B.n161 VSUBS 0.010644f
C196 B.n162 VSUBS 0.010644f
C197 B.n163 VSUBS 0.010644f
C198 B.n164 VSUBS 0.010644f
C199 B.n165 VSUBS 0.010644f
C200 B.n166 VSUBS 0.010644f
C201 B.n167 VSUBS 0.010644f
C202 B.t7 VSUBS 0.356728f
C203 B.t8 VSUBS 0.395666f
C204 B.t6 VSUBS 1.90543f
C205 B.n168 VSUBS 0.228095f
C206 B.n169 VSUBS 0.113841f
C207 B.n170 VSUBS 0.010644f
C208 B.n171 VSUBS 0.010644f
C209 B.n172 VSUBS 0.010644f
C210 B.n173 VSUBS 0.010644f
C211 B.t4 VSUBS 0.356731f
C212 B.t5 VSUBS 0.395669f
C213 B.t3 VSUBS 1.90543f
C214 B.n174 VSUBS 0.228091f
C215 B.n175 VSUBS 0.113839f
C216 B.n176 VSUBS 0.024661f
C217 B.n177 VSUBS 0.010644f
C218 B.n178 VSUBS 0.010644f
C219 B.n179 VSUBS 0.010644f
C220 B.n180 VSUBS 0.010644f
C221 B.n181 VSUBS 0.010644f
C222 B.n182 VSUBS 0.010644f
C223 B.n183 VSUBS 0.010644f
C224 B.n184 VSUBS 0.010644f
C225 B.n185 VSUBS 0.010644f
C226 B.n186 VSUBS 0.010644f
C227 B.n187 VSUBS 0.010644f
C228 B.n188 VSUBS 0.010644f
C229 B.n189 VSUBS 0.010644f
C230 B.n190 VSUBS 0.010644f
C231 B.n191 VSUBS 0.024309f
C232 B.n192 VSUBS 0.010644f
C233 B.n193 VSUBS 0.010644f
C234 B.n194 VSUBS 0.010644f
C235 B.n195 VSUBS 0.010644f
C236 B.n196 VSUBS 0.010644f
C237 B.n197 VSUBS 0.010644f
C238 B.n198 VSUBS 0.010644f
C239 B.n199 VSUBS 0.010644f
C240 B.n200 VSUBS 0.010644f
C241 B.n201 VSUBS 0.010644f
C242 B.n202 VSUBS 0.010644f
C243 B.n203 VSUBS 0.010644f
C244 B.n204 VSUBS 0.010644f
C245 B.n205 VSUBS 0.010644f
C246 B.n206 VSUBS 0.010644f
C247 B.n207 VSUBS 0.010644f
C248 B.n208 VSUBS 0.010644f
C249 B.n209 VSUBS 0.010644f
C250 B.n210 VSUBS 0.010644f
C251 B.n211 VSUBS 0.010644f
C252 B.n212 VSUBS 0.010644f
C253 B.n213 VSUBS 0.010644f
C254 B.n214 VSUBS 0.010644f
C255 B.n215 VSUBS 0.010644f
C256 B.n216 VSUBS 0.010644f
C257 B.n217 VSUBS 0.010644f
C258 B.n218 VSUBS 0.010644f
C259 B.n219 VSUBS 0.010644f
C260 B.n220 VSUBS 0.010644f
C261 B.n221 VSUBS 0.010644f
C262 B.n222 VSUBS 0.010644f
C263 B.n223 VSUBS 0.010644f
C264 B.n224 VSUBS 0.010644f
C265 B.n225 VSUBS 0.010644f
C266 B.n226 VSUBS 0.010644f
C267 B.n227 VSUBS 0.010644f
C268 B.n228 VSUBS 0.010644f
C269 B.n229 VSUBS 0.010644f
C270 B.n230 VSUBS 0.010644f
C271 B.n231 VSUBS 0.010644f
C272 B.n232 VSUBS 0.010644f
C273 B.n233 VSUBS 0.010644f
C274 B.n234 VSUBS 0.010644f
C275 B.n235 VSUBS 0.010644f
C276 B.n236 VSUBS 0.010644f
C277 B.n237 VSUBS 0.010644f
C278 B.n238 VSUBS 0.010644f
C279 B.n239 VSUBS 0.010644f
C280 B.n240 VSUBS 0.010644f
C281 B.n241 VSUBS 0.010644f
C282 B.n242 VSUBS 0.010644f
C283 B.n243 VSUBS 0.010644f
C284 B.n244 VSUBS 0.010644f
C285 B.n245 VSUBS 0.010644f
C286 B.n246 VSUBS 0.010644f
C287 B.n247 VSUBS 0.010644f
C288 B.n248 VSUBS 0.010644f
C289 B.n249 VSUBS 0.010644f
C290 B.n250 VSUBS 0.010644f
C291 B.n251 VSUBS 0.010644f
C292 B.n252 VSUBS 0.010644f
C293 B.n253 VSUBS 0.010644f
C294 B.n254 VSUBS 0.010644f
C295 B.n255 VSUBS 0.010644f
C296 B.n256 VSUBS 0.010644f
C297 B.n257 VSUBS 0.010644f
C298 B.n258 VSUBS 0.010644f
C299 B.n259 VSUBS 0.010644f
C300 B.n260 VSUBS 0.010644f
C301 B.n261 VSUBS 0.010644f
C302 B.n262 VSUBS 0.010644f
C303 B.n263 VSUBS 0.010644f
C304 B.n264 VSUBS 0.010644f
C305 B.n265 VSUBS 0.010644f
C306 B.n266 VSUBS 0.010644f
C307 B.n267 VSUBS 0.010644f
C308 B.n268 VSUBS 0.010644f
C309 B.n269 VSUBS 0.010644f
C310 B.n270 VSUBS 0.010644f
C311 B.n271 VSUBS 0.010644f
C312 B.n272 VSUBS 0.010644f
C313 B.n273 VSUBS 0.010644f
C314 B.n274 VSUBS 0.010644f
C315 B.n275 VSUBS 0.010644f
C316 B.n276 VSUBS 0.010644f
C317 B.n277 VSUBS 0.010644f
C318 B.n278 VSUBS 0.010644f
C319 B.n279 VSUBS 0.010644f
C320 B.n280 VSUBS 0.010644f
C321 B.n281 VSUBS 0.010644f
C322 B.n282 VSUBS 0.010644f
C323 B.n283 VSUBS 0.010644f
C324 B.n284 VSUBS 0.010644f
C325 B.n285 VSUBS 0.010644f
C326 B.n286 VSUBS 0.010644f
C327 B.n287 VSUBS 0.010644f
C328 B.n288 VSUBS 0.010644f
C329 B.n289 VSUBS 0.010644f
C330 B.n290 VSUBS 0.010644f
C331 B.n291 VSUBS 0.010644f
C332 B.n292 VSUBS 0.010644f
C333 B.n293 VSUBS 0.010644f
C334 B.n294 VSUBS 0.010644f
C335 B.n295 VSUBS 0.010644f
C336 B.n296 VSUBS 0.010644f
C337 B.n297 VSUBS 0.010644f
C338 B.n298 VSUBS 0.010644f
C339 B.n299 VSUBS 0.010644f
C340 B.n300 VSUBS 0.010644f
C341 B.n301 VSUBS 0.010644f
C342 B.n302 VSUBS 0.010644f
C343 B.n303 VSUBS 0.010644f
C344 B.n304 VSUBS 0.010644f
C345 B.n305 VSUBS 0.010644f
C346 B.n306 VSUBS 0.010644f
C347 B.n307 VSUBS 0.010644f
C348 B.n308 VSUBS 0.010644f
C349 B.n309 VSUBS 0.010644f
C350 B.n310 VSUBS 0.010644f
C351 B.n311 VSUBS 0.010644f
C352 B.n312 VSUBS 0.010644f
C353 B.n313 VSUBS 0.010644f
C354 B.n314 VSUBS 0.010644f
C355 B.n315 VSUBS 0.010644f
C356 B.n316 VSUBS 0.010644f
C357 B.n317 VSUBS 0.010644f
C358 B.n318 VSUBS 0.010644f
C359 B.n319 VSUBS 0.010644f
C360 B.n320 VSUBS 0.010644f
C361 B.n321 VSUBS 0.010644f
C362 B.n322 VSUBS 0.010644f
C363 B.n323 VSUBS 0.010644f
C364 B.n324 VSUBS 0.010644f
C365 B.n325 VSUBS 0.010644f
C366 B.n326 VSUBS 0.010644f
C367 B.n327 VSUBS 0.010644f
C368 B.n328 VSUBS 0.010644f
C369 B.n329 VSUBS 0.010644f
C370 B.n330 VSUBS 0.010644f
C371 B.n331 VSUBS 0.010644f
C372 B.n332 VSUBS 0.010644f
C373 B.n333 VSUBS 0.010644f
C374 B.n334 VSUBS 0.010644f
C375 B.n335 VSUBS 0.010644f
C376 B.n336 VSUBS 0.010644f
C377 B.n337 VSUBS 0.010644f
C378 B.n338 VSUBS 0.024309f
C379 B.n339 VSUBS 0.024841f
C380 B.n340 VSUBS 0.024841f
C381 B.n341 VSUBS 0.010644f
C382 B.n342 VSUBS 0.010644f
C383 B.n343 VSUBS 0.010644f
C384 B.n344 VSUBS 0.010644f
C385 B.n345 VSUBS 0.010644f
C386 B.n346 VSUBS 0.010644f
C387 B.n347 VSUBS 0.010644f
C388 B.n348 VSUBS 0.010644f
C389 B.n349 VSUBS 0.010644f
C390 B.n350 VSUBS 0.010644f
C391 B.n351 VSUBS 0.010644f
C392 B.n352 VSUBS 0.010644f
C393 B.n353 VSUBS 0.010644f
C394 B.n354 VSUBS 0.010644f
C395 B.n355 VSUBS 0.010644f
C396 B.n356 VSUBS 0.010644f
C397 B.n357 VSUBS 0.010644f
C398 B.n358 VSUBS 0.010644f
C399 B.n359 VSUBS 0.010644f
C400 B.n360 VSUBS 0.010644f
C401 B.n361 VSUBS 0.010644f
C402 B.n362 VSUBS 0.010644f
C403 B.n363 VSUBS 0.010644f
C404 B.n364 VSUBS 0.010644f
C405 B.n365 VSUBS 0.010644f
C406 B.n366 VSUBS 0.010644f
C407 B.n367 VSUBS 0.010644f
C408 B.n368 VSUBS 0.010644f
C409 B.n369 VSUBS 0.010644f
C410 B.n370 VSUBS 0.010644f
C411 B.n371 VSUBS 0.010644f
C412 B.n372 VSUBS 0.010644f
C413 B.n373 VSUBS 0.010644f
C414 B.n374 VSUBS 0.010644f
C415 B.n375 VSUBS 0.010644f
C416 B.n376 VSUBS 0.010644f
C417 B.n377 VSUBS 0.010644f
C418 B.n378 VSUBS 0.010644f
C419 B.n379 VSUBS 0.010644f
C420 B.n380 VSUBS 0.010644f
C421 B.n381 VSUBS 0.007357f
C422 B.n382 VSUBS 0.010644f
C423 B.n383 VSUBS 0.010644f
C424 B.n384 VSUBS 0.008609f
C425 B.n385 VSUBS 0.010644f
C426 B.n386 VSUBS 0.010644f
C427 B.n387 VSUBS 0.010644f
C428 B.n388 VSUBS 0.010644f
C429 B.n389 VSUBS 0.010644f
C430 B.n390 VSUBS 0.010644f
C431 B.n391 VSUBS 0.010644f
C432 B.n392 VSUBS 0.010644f
C433 B.n393 VSUBS 0.010644f
C434 B.n394 VSUBS 0.010644f
C435 B.n395 VSUBS 0.010644f
C436 B.n396 VSUBS 0.008609f
C437 B.n397 VSUBS 0.024661f
C438 B.n398 VSUBS 0.007357f
C439 B.n399 VSUBS 0.010644f
C440 B.n400 VSUBS 0.010644f
C441 B.n401 VSUBS 0.010644f
C442 B.n402 VSUBS 0.010644f
C443 B.n403 VSUBS 0.010644f
C444 B.n404 VSUBS 0.010644f
C445 B.n405 VSUBS 0.010644f
C446 B.n406 VSUBS 0.010644f
C447 B.n407 VSUBS 0.010644f
C448 B.n408 VSUBS 0.010644f
C449 B.n409 VSUBS 0.010644f
C450 B.n410 VSUBS 0.010644f
C451 B.n411 VSUBS 0.010644f
C452 B.n412 VSUBS 0.010644f
C453 B.n413 VSUBS 0.010644f
C454 B.n414 VSUBS 0.010644f
C455 B.n415 VSUBS 0.010644f
C456 B.n416 VSUBS 0.010644f
C457 B.n417 VSUBS 0.010644f
C458 B.n418 VSUBS 0.010644f
C459 B.n419 VSUBS 0.010644f
C460 B.n420 VSUBS 0.010644f
C461 B.n421 VSUBS 0.010644f
C462 B.n422 VSUBS 0.010644f
C463 B.n423 VSUBS 0.010644f
C464 B.n424 VSUBS 0.010644f
C465 B.n425 VSUBS 0.010644f
C466 B.n426 VSUBS 0.010644f
C467 B.n427 VSUBS 0.010644f
C468 B.n428 VSUBS 0.010644f
C469 B.n429 VSUBS 0.010644f
C470 B.n430 VSUBS 0.010644f
C471 B.n431 VSUBS 0.010644f
C472 B.n432 VSUBS 0.010644f
C473 B.n433 VSUBS 0.010644f
C474 B.n434 VSUBS 0.010644f
C475 B.n435 VSUBS 0.010644f
C476 B.n436 VSUBS 0.010644f
C477 B.n437 VSUBS 0.010644f
C478 B.n438 VSUBS 0.010644f
C479 B.n439 VSUBS 0.010644f
C480 B.n440 VSUBS 0.024841f
C481 B.n441 VSUBS 0.024309f
C482 B.n442 VSUBS 0.024309f
C483 B.n443 VSUBS 0.010644f
C484 B.n444 VSUBS 0.010644f
C485 B.n445 VSUBS 0.010644f
C486 B.n446 VSUBS 0.010644f
C487 B.n447 VSUBS 0.010644f
C488 B.n448 VSUBS 0.010644f
C489 B.n449 VSUBS 0.010644f
C490 B.n450 VSUBS 0.010644f
C491 B.n451 VSUBS 0.010644f
C492 B.n452 VSUBS 0.010644f
C493 B.n453 VSUBS 0.010644f
C494 B.n454 VSUBS 0.010644f
C495 B.n455 VSUBS 0.010644f
C496 B.n456 VSUBS 0.010644f
C497 B.n457 VSUBS 0.010644f
C498 B.n458 VSUBS 0.010644f
C499 B.n459 VSUBS 0.010644f
C500 B.n460 VSUBS 0.010644f
C501 B.n461 VSUBS 0.010644f
C502 B.n462 VSUBS 0.010644f
C503 B.n463 VSUBS 0.010644f
C504 B.n464 VSUBS 0.010644f
C505 B.n465 VSUBS 0.010644f
C506 B.n466 VSUBS 0.010644f
C507 B.n467 VSUBS 0.010644f
C508 B.n468 VSUBS 0.010644f
C509 B.n469 VSUBS 0.010644f
C510 B.n470 VSUBS 0.010644f
C511 B.n471 VSUBS 0.010644f
C512 B.n472 VSUBS 0.010644f
C513 B.n473 VSUBS 0.010644f
C514 B.n474 VSUBS 0.010644f
C515 B.n475 VSUBS 0.010644f
C516 B.n476 VSUBS 0.010644f
C517 B.n477 VSUBS 0.010644f
C518 B.n478 VSUBS 0.010644f
C519 B.n479 VSUBS 0.010644f
C520 B.n480 VSUBS 0.010644f
C521 B.n481 VSUBS 0.010644f
C522 B.n482 VSUBS 0.010644f
C523 B.n483 VSUBS 0.010644f
C524 B.n484 VSUBS 0.010644f
C525 B.n485 VSUBS 0.010644f
C526 B.n486 VSUBS 0.010644f
C527 B.n487 VSUBS 0.010644f
C528 B.n488 VSUBS 0.010644f
C529 B.n489 VSUBS 0.010644f
C530 B.n490 VSUBS 0.010644f
C531 B.n491 VSUBS 0.010644f
C532 B.n492 VSUBS 0.010644f
C533 B.n493 VSUBS 0.010644f
C534 B.n494 VSUBS 0.010644f
C535 B.n495 VSUBS 0.010644f
C536 B.n496 VSUBS 0.010644f
C537 B.n497 VSUBS 0.010644f
C538 B.n498 VSUBS 0.010644f
C539 B.n499 VSUBS 0.010644f
C540 B.n500 VSUBS 0.010644f
C541 B.n501 VSUBS 0.010644f
C542 B.n502 VSUBS 0.010644f
C543 B.n503 VSUBS 0.010644f
C544 B.n504 VSUBS 0.010644f
C545 B.n505 VSUBS 0.010644f
C546 B.n506 VSUBS 0.010644f
C547 B.n507 VSUBS 0.010644f
C548 B.n508 VSUBS 0.010644f
C549 B.n509 VSUBS 0.010644f
C550 B.n510 VSUBS 0.010644f
C551 B.n511 VSUBS 0.010644f
C552 B.n512 VSUBS 0.010644f
C553 B.n513 VSUBS 0.010644f
C554 B.n514 VSUBS 0.010644f
C555 B.n515 VSUBS 0.010644f
C556 B.n516 VSUBS 0.010644f
C557 B.n517 VSUBS 0.010644f
C558 B.n518 VSUBS 0.010644f
C559 B.n519 VSUBS 0.010644f
C560 B.n520 VSUBS 0.010644f
C561 B.n521 VSUBS 0.010644f
C562 B.n522 VSUBS 0.010644f
C563 B.n523 VSUBS 0.010644f
C564 B.n524 VSUBS 0.010644f
C565 B.n525 VSUBS 0.010644f
C566 B.n526 VSUBS 0.010644f
C567 B.n527 VSUBS 0.010644f
C568 B.n528 VSUBS 0.010644f
C569 B.n529 VSUBS 0.010644f
C570 B.n530 VSUBS 0.010644f
C571 B.n531 VSUBS 0.010644f
C572 B.n532 VSUBS 0.010644f
C573 B.n533 VSUBS 0.010644f
C574 B.n534 VSUBS 0.010644f
C575 B.n535 VSUBS 0.010644f
C576 B.n536 VSUBS 0.010644f
C577 B.n537 VSUBS 0.010644f
C578 B.n538 VSUBS 0.010644f
C579 B.n539 VSUBS 0.010644f
C580 B.n540 VSUBS 0.010644f
C581 B.n541 VSUBS 0.010644f
C582 B.n542 VSUBS 0.010644f
C583 B.n543 VSUBS 0.010644f
C584 B.n544 VSUBS 0.010644f
C585 B.n545 VSUBS 0.010644f
C586 B.n546 VSUBS 0.010644f
C587 B.n547 VSUBS 0.010644f
C588 B.n548 VSUBS 0.010644f
C589 B.n549 VSUBS 0.010644f
C590 B.n550 VSUBS 0.010644f
C591 B.n551 VSUBS 0.010644f
C592 B.n552 VSUBS 0.010644f
C593 B.n553 VSUBS 0.010644f
C594 B.n554 VSUBS 0.010644f
C595 B.n555 VSUBS 0.010644f
C596 B.n556 VSUBS 0.010644f
C597 B.n557 VSUBS 0.010644f
C598 B.n558 VSUBS 0.010644f
C599 B.n559 VSUBS 0.010644f
C600 B.n560 VSUBS 0.010644f
C601 B.n561 VSUBS 0.010644f
C602 B.n562 VSUBS 0.010644f
C603 B.n563 VSUBS 0.010644f
C604 B.n564 VSUBS 0.010644f
C605 B.n565 VSUBS 0.010644f
C606 B.n566 VSUBS 0.010644f
C607 B.n567 VSUBS 0.010644f
C608 B.n568 VSUBS 0.010644f
C609 B.n569 VSUBS 0.010644f
C610 B.n570 VSUBS 0.010644f
C611 B.n571 VSUBS 0.010644f
C612 B.n572 VSUBS 0.010644f
C613 B.n573 VSUBS 0.010644f
C614 B.n574 VSUBS 0.010644f
C615 B.n575 VSUBS 0.010644f
C616 B.n576 VSUBS 0.010644f
C617 B.n577 VSUBS 0.010644f
C618 B.n578 VSUBS 0.010644f
C619 B.n579 VSUBS 0.010644f
C620 B.n580 VSUBS 0.010644f
C621 B.n581 VSUBS 0.010644f
C622 B.n582 VSUBS 0.010644f
C623 B.n583 VSUBS 0.010644f
C624 B.n584 VSUBS 0.010644f
C625 B.n585 VSUBS 0.010644f
C626 B.n586 VSUBS 0.010644f
C627 B.n587 VSUBS 0.010644f
C628 B.n588 VSUBS 0.010644f
C629 B.n589 VSUBS 0.010644f
C630 B.n590 VSUBS 0.010644f
C631 B.n591 VSUBS 0.010644f
C632 B.n592 VSUBS 0.010644f
C633 B.n593 VSUBS 0.010644f
C634 B.n594 VSUBS 0.010644f
C635 B.n595 VSUBS 0.010644f
C636 B.n596 VSUBS 0.010644f
C637 B.n597 VSUBS 0.010644f
C638 B.n598 VSUBS 0.010644f
C639 B.n599 VSUBS 0.010644f
C640 B.n600 VSUBS 0.010644f
C641 B.n601 VSUBS 0.010644f
C642 B.n602 VSUBS 0.010644f
C643 B.n603 VSUBS 0.010644f
C644 B.n604 VSUBS 0.010644f
C645 B.n605 VSUBS 0.010644f
C646 B.n606 VSUBS 0.010644f
C647 B.n607 VSUBS 0.010644f
C648 B.n608 VSUBS 0.010644f
C649 B.n609 VSUBS 0.010644f
C650 B.n610 VSUBS 0.010644f
C651 B.n611 VSUBS 0.010644f
C652 B.n612 VSUBS 0.010644f
C653 B.n613 VSUBS 0.010644f
C654 B.n614 VSUBS 0.010644f
C655 B.n615 VSUBS 0.010644f
C656 B.n616 VSUBS 0.010644f
C657 B.n617 VSUBS 0.010644f
C658 B.n618 VSUBS 0.010644f
C659 B.n619 VSUBS 0.010644f
C660 B.n620 VSUBS 0.010644f
C661 B.n621 VSUBS 0.010644f
C662 B.n622 VSUBS 0.010644f
C663 B.n623 VSUBS 0.010644f
C664 B.n624 VSUBS 0.010644f
C665 B.n625 VSUBS 0.010644f
C666 B.n626 VSUBS 0.010644f
C667 B.n627 VSUBS 0.010644f
C668 B.n628 VSUBS 0.010644f
C669 B.n629 VSUBS 0.010644f
C670 B.n630 VSUBS 0.010644f
C671 B.n631 VSUBS 0.010644f
C672 B.n632 VSUBS 0.010644f
C673 B.n633 VSUBS 0.010644f
C674 B.n634 VSUBS 0.010644f
C675 B.n635 VSUBS 0.010644f
C676 B.n636 VSUBS 0.010644f
C677 B.n637 VSUBS 0.010644f
C678 B.n638 VSUBS 0.010644f
C679 B.n639 VSUBS 0.010644f
C680 B.n640 VSUBS 0.010644f
C681 B.n641 VSUBS 0.010644f
C682 B.n642 VSUBS 0.010644f
C683 B.n643 VSUBS 0.010644f
C684 B.n644 VSUBS 0.010644f
C685 B.n645 VSUBS 0.010644f
C686 B.n646 VSUBS 0.010644f
C687 B.n647 VSUBS 0.010644f
C688 B.n648 VSUBS 0.010644f
C689 B.n649 VSUBS 0.010644f
C690 B.n650 VSUBS 0.010644f
C691 B.n651 VSUBS 0.010644f
C692 B.n652 VSUBS 0.010644f
C693 B.n653 VSUBS 0.010644f
C694 B.n654 VSUBS 0.010644f
C695 B.n655 VSUBS 0.010644f
C696 B.n656 VSUBS 0.010644f
C697 B.n657 VSUBS 0.010644f
C698 B.n658 VSUBS 0.010644f
C699 B.n659 VSUBS 0.010644f
C700 B.n660 VSUBS 0.010644f
C701 B.n661 VSUBS 0.010644f
C702 B.n662 VSUBS 0.010644f
C703 B.n663 VSUBS 0.010644f
C704 B.n664 VSUBS 0.010644f
C705 B.n665 VSUBS 0.010644f
C706 B.n666 VSUBS 0.024309f
C707 B.n667 VSUBS 0.025593f
C708 B.n668 VSUBS 0.023558f
C709 B.n669 VSUBS 0.010644f
C710 B.n670 VSUBS 0.010644f
C711 B.n671 VSUBS 0.010644f
C712 B.n672 VSUBS 0.010644f
C713 B.n673 VSUBS 0.010644f
C714 B.n674 VSUBS 0.010644f
C715 B.n675 VSUBS 0.010644f
C716 B.n676 VSUBS 0.010644f
C717 B.n677 VSUBS 0.010644f
C718 B.n678 VSUBS 0.010644f
C719 B.n679 VSUBS 0.010644f
C720 B.n680 VSUBS 0.010644f
C721 B.n681 VSUBS 0.010644f
C722 B.n682 VSUBS 0.010644f
C723 B.n683 VSUBS 0.010644f
C724 B.n684 VSUBS 0.010644f
C725 B.n685 VSUBS 0.010644f
C726 B.n686 VSUBS 0.010644f
C727 B.n687 VSUBS 0.010644f
C728 B.n688 VSUBS 0.010644f
C729 B.n689 VSUBS 0.010644f
C730 B.n690 VSUBS 0.010644f
C731 B.n691 VSUBS 0.010644f
C732 B.n692 VSUBS 0.010644f
C733 B.n693 VSUBS 0.010644f
C734 B.n694 VSUBS 0.010644f
C735 B.n695 VSUBS 0.010644f
C736 B.n696 VSUBS 0.010644f
C737 B.n697 VSUBS 0.010644f
C738 B.n698 VSUBS 0.010644f
C739 B.n699 VSUBS 0.010644f
C740 B.n700 VSUBS 0.010644f
C741 B.n701 VSUBS 0.010644f
C742 B.n702 VSUBS 0.010644f
C743 B.n703 VSUBS 0.010644f
C744 B.n704 VSUBS 0.010644f
C745 B.n705 VSUBS 0.010644f
C746 B.n706 VSUBS 0.010644f
C747 B.n707 VSUBS 0.010644f
C748 B.n708 VSUBS 0.010644f
C749 B.n709 VSUBS 0.010644f
C750 B.n710 VSUBS 0.007357f
C751 B.n711 VSUBS 0.024661f
C752 B.n712 VSUBS 0.008609f
C753 B.n713 VSUBS 0.010644f
C754 B.n714 VSUBS 0.010644f
C755 B.n715 VSUBS 0.010644f
C756 B.n716 VSUBS 0.010644f
C757 B.n717 VSUBS 0.010644f
C758 B.n718 VSUBS 0.010644f
C759 B.n719 VSUBS 0.010644f
C760 B.n720 VSUBS 0.010644f
C761 B.n721 VSUBS 0.010644f
C762 B.n722 VSUBS 0.010644f
C763 B.n723 VSUBS 0.010644f
C764 B.n724 VSUBS 0.008609f
C765 B.n725 VSUBS 0.010644f
C766 B.n726 VSUBS 0.010644f
C767 B.n727 VSUBS 0.007357f
C768 B.n728 VSUBS 0.010644f
C769 B.n729 VSUBS 0.010644f
C770 B.n730 VSUBS 0.010644f
C771 B.n731 VSUBS 0.010644f
C772 B.n732 VSUBS 0.010644f
C773 B.n733 VSUBS 0.010644f
C774 B.n734 VSUBS 0.010644f
C775 B.n735 VSUBS 0.010644f
C776 B.n736 VSUBS 0.010644f
C777 B.n737 VSUBS 0.010644f
C778 B.n738 VSUBS 0.010644f
C779 B.n739 VSUBS 0.010644f
C780 B.n740 VSUBS 0.010644f
C781 B.n741 VSUBS 0.010644f
C782 B.n742 VSUBS 0.010644f
C783 B.n743 VSUBS 0.010644f
C784 B.n744 VSUBS 0.010644f
C785 B.n745 VSUBS 0.010644f
C786 B.n746 VSUBS 0.010644f
C787 B.n747 VSUBS 0.010644f
C788 B.n748 VSUBS 0.010644f
C789 B.n749 VSUBS 0.010644f
C790 B.n750 VSUBS 0.010644f
C791 B.n751 VSUBS 0.010644f
C792 B.n752 VSUBS 0.010644f
C793 B.n753 VSUBS 0.010644f
C794 B.n754 VSUBS 0.010644f
C795 B.n755 VSUBS 0.010644f
C796 B.n756 VSUBS 0.010644f
C797 B.n757 VSUBS 0.010644f
C798 B.n758 VSUBS 0.010644f
C799 B.n759 VSUBS 0.010644f
C800 B.n760 VSUBS 0.010644f
C801 B.n761 VSUBS 0.010644f
C802 B.n762 VSUBS 0.010644f
C803 B.n763 VSUBS 0.010644f
C804 B.n764 VSUBS 0.010644f
C805 B.n765 VSUBS 0.010644f
C806 B.n766 VSUBS 0.010644f
C807 B.n767 VSUBS 0.010644f
C808 B.n768 VSUBS 0.024841f
C809 B.n769 VSUBS 0.024841f
C810 B.n770 VSUBS 0.024309f
C811 B.n771 VSUBS 0.010644f
C812 B.n772 VSUBS 0.010644f
C813 B.n773 VSUBS 0.010644f
C814 B.n774 VSUBS 0.010644f
C815 B.n775 VSUBS 0.010644f
C816 B.n776 VSUBS 0.010644f
C817 B.n777 VSUBS 0.010644f
C818 B.n778 VSUBS 0.010644f
C819 B.n779 VSUBS 0.010644f
C820 B.n780 VSUBS 0.010644f
C821 B.n781 VSUBS 0.010644f
C822 B.n782 VSUBS 0.010644f
C823 B.n783 VSUBS 0.010644f
C824 B.n784 VSUBS 0.010644f
C825 B.n785 VSUBS 0.010644f
C826 B.n786 VSUBS 0.010644f
C827 B.n787 VSUBS 0.010644f
C828 B.n788 VSUBS 0.010644f
C829 B.n789 VSUBS 0.010644f
C830 B.n790 VSUBS 0.010644f
C831 B.n791 VSUBS 0.010644f
C832 B.n792 VSUBS 0.010644f
C833 B.n793 VSUBS 0.010644f
C834 B.n794 VSUBS 0.010644f
C835 B.n795 VSUBS 0.010644f
C836 B.n796 VSUBS 0.010644f
C837 B.n797 VSUBS 0.010644f
C838 B.n798 VSUBS 0.010644f
C839 B.n799 VSUBS 0.010644f
C840 B.n800 VSUBS 0.010644f
C841 B.n801 VSUBS 0.010644f
C842 B.n802 VSUBS 0.010644f
C843 B.n803 VSUBS 0.010644f
C844 B.n804 VSUBS 0.010644f
C845 B.n805 VSUBS 0.010644f
C846 B.n806 VSUBS 0.010644f
C847 B.n807 VSUBS 0.010644f
C848 B.n808 VSUBS 0.010644f
C849 B.n809 VSUBS 0.010644f
C850 B.n810 VSUBS 0.010644f
C851 B.n811 VSUBS 0.010644f
C852 B.n812 VSUBS 0.010644f
C853 B.n813 VSUBS 0.010644f
C854 B.n814 VSUBS 0.010644f
C855 B.n815 VSUBS 0.010644f
C856 B.n816 VSUBS 0.010644f
C857 B.n817 VSUBS 0.010644f
C858 B.n818 VSUBS 0.010644f
C859 B.n819 VSUBS 0.010644f
C860 B.n820 VSUBS 0.010644f
C861 B.n821 VSUBS 0.010644f
C862 B.n822 VSUBS 0.010644f
C863 B.n823 VSUBS 0.010644f
C864 B.n824 VSUBS 0.010644f
C865 B.n825 VSUBS 0.010644f
C866 B.n826 VSUBS 0.010644f
C867 B.n827 VSUBS 0.010644f
C868 B.n828 VSUBS 0.010644f
C869 B.n829 VSUBS 0.010644f
C870 B.n830 VSUBS 0.010644f
C871 B.n831 VSUBS 0.010644f
C872 B.n832 VSUBS 0.010644f
C873 B.n833 VSUBS 0.010644f
C874 B.n834 VSUBS 0.010644f
C875 B.n835 VSUBS 0.010644f
C876 B.n836 VSUBS 0.010644f
C877 B.n837 VSUBS 0.010644f
C878 B.n838 VSUBS 0.010644f
C879 B.n839 VSUBS 0.010644f
C880 B.n840 VSUBS 0.010644f
C881 B.n841 VSUBS 0.010644f
C882 B.n842 VSUBS 0.010644f
C883 B.n843 VSUBS 0.010644f
C884 B.n844 VSUBS 0.010644f
C885 B.n845 VSUBS 0.010644f
C886 B.n846 VSUBS 0.010644f
C887 B.n847 VSUBS 0.010644f
C888 B.n848 VSUBS 0.010644f
C889 B.n849 VSUBS 0.010644f
C890 B.n850 VSUBS 0.010644f
C891 B.n851 VSUBS 0.010644f
C892 B.n852 VSUBS 0.010644f
C893 B.n853 VSUBS 0.010644f
C894 B.n854 VSUBS 0.010644f
C895 B.n855 VSUBS 0.010644f
C896 B.n856 VSUBS 0.010644f
C897 B.n857 VSUBS 0.010644f
C898 B.n858 VSUBS 0.010644f
C899 B.n859 VSUBS 0.010644f
C900 B.n860 VSUBS 0.010644f
C901 B.n861 VSUBS 0.010644f
C902 B.n862 VSUBS 0.010644f
C903 B.n863 VSUBS 0.010644f
C904 B.n864 VSUBS 0.010644f
C905 B.n865 VSUBS 0.010644f
C906 B.n866 VSUBS 0.010644f
C907 B.n867 VSUBS 0.010644f
C908 B.n868 VSUBS 0.010644f
C909 B.n869 VSUBS 0.010644f
C910 B.n870 VSUBS 0.010644f
C911 B.n871 VSUBS 0.010644f
C912 B.n872 VSUBS 0.010644f
C913 B.n873 VSUBS 0.010644f
C914 B.n874 VSUBS 0.010644f
C915 B.n875 VSUBS 0.010644f
C916 B.n876 VSUBS 0.010644f
C917 B.n877 VSUBS 0.010644f
C918 B.n878 VSUBS 0.010644f
C919 B.n879 VSUBS 0.010644f
C920 B.n880 VSUBS 0.010644f
C921 B.n881 VSUBS 0.010644f
C922 B.n882 VSUBS 0.010644f
C923 B.n883 VSUBS 0.024102f
C924 VDD2.t0 VSUBS 1.96843f
C925 VDD2.t6 VSUBS 0.203282f
C926 VDD2.t3 VSUBS 0.203282f
C927 VDD2.n0 VSUBS 1.46326f
C928 VDD2.n1 VSUBS 1.96408f
C929 VDD2.t2 VSUBS 0.203282f
C930 VDD2.t7 VSUBS 0.203282f
C931 VDD2.n2 VSUBS 1.49455f
C932 VDD2.n3 VSUBS 4.419509f
C933 VDD2.t5 VSUBS 1.93403f
C934 VDD2.n4 VSUBS 4.46647f
C935 VDD2.t1 VSUBS 0.203282f
C936 VDD2.t8 VSUBS 0.203282f
C937 VDD2.n5 VSUBS 1.46327f
C938 VDD2.n6 VSUBS 1.00351f
C939 VDD2.t9 VSUBS 0.203282f
C940 VDD2.t4 VSUBS 0.203282f
C941 VDD2.n7 VSUBS 1.4945f
C942 VN.t2 VSUBS 2.02839f
C943 VN.n0 VSUBS 0.850596f
C944 VN.n1 VSUBS 0.028634f
C945 VN.n2 VSUBS 0.025552f
C946 VN.n3 VSUBS 0.028634f
C947 VN.t7 VSUBS 2.02839f
C948 VN.n4 VSUBS 0.733107f
C949 VN.n5 VSUBS 0.028634f
C950 VN.n6 VSUBS 0.049952f
C951 VN.n7 VSUBS 0.028634f
C952 VN.n8 VSUBS 0.039993f
C953 VN.n9 VSUBS 0.028634f
C954 VN.n10 VSUBS 0.031181f
C955 VN.n11 VSUBS 0.028634f
C956 VN.n12 VSUBS 0.028459f
C957 VN.t3 VSUBS 2.02839f
C958 VN.n13 VSUBS 0.820369f
C959 VN.t9 VSUBS 2.38746f
C960 VN.n14 VSUBS 0.780492f
C961 VN.n15 VSUBS 0.341468f
C962 VN.n16 VSUBS 0.028634f
C963 VN.n17 VSUBS 0.0531f
C964 VN.n18 VSUBS 0.0531f
C965 VN.n19 VSUBS 0.049952f
C966 VN.n20 VSUBS 0.028634f
C967 VN.n21 VSUBS 0.028634f
C968 VN.n22 VSUBS 0.028634f
C969 VN.n23 VSUBS 0.055215f
C970 VN.n24 VSUBS 0.0531f
C971 VN.t6 VSUBS 2.02839f
C972 VN.n25 VSUBS 0.733107f
C973 VN.n26 VSUBS 0.039993f
C974 VN.n27 VSUBS 0.028634f
C975 VN.n28 VSUBS 0.028634f
C976 VN.n29 VSUBS 0.028634f
C977 VN.n30 VSUBS 0.0531f
C978 VN.n31 VSUBS 0.055215f
C979 VN.n32 VSUBS 0.031181f
C980 VN.n33 VSUBS 0.028634f
C981 VN.n34 VSUBS 0.028634f
C982 VN.n35 VSUBS 0.028634f
C983 VN.n36 VSUBS 0.0531f
C984 VN.n37 VSUBS 0.0531f
C985 VN.n38 VSUBS 0.028459f
C986 VN.n39 VSUBS 0.028634f
C987 VN.n40 VSUBS 0.028634f
C988 VN.n41 VSUBS 0.051527f
C989 VN.n42 VSUBS 0.0531f
C990 VN.n43 VSUBS 0.053357f
C991 VN.n44 VSUBS 0.028634f
C992 VN.n45 VSUBS 0.028634f
C993 VN.n46 VSUBS 0.028634f
C994 VN.n47 VSUBS 0.05744f
C995 VN.n48 VSUBS 0.0531f
C996 VN.n49 VSUBS 0.043138f
C997 VN.n50 VSUBS 0.046208f
C998 VN.n51 VSUBS 0.070384f
C999 VN.t4 VSUBS 2.02839f
C1000 VN.n52 VSUBS 0.850596f
C1001 VN.n53 VSUBS 0.028634f
C1002 VN.n54 VSUBS 0.025552f
C1003 VN.n55 VSUBS 0.028634f
C1004 VN.t8 VSUBS 2.02839f
C1005 VN.n56 VSUBS 0.733107f
C1006 VN.n57 VSUBS 0.028634f
C1007 VN.n58 VSUBS 0.049952f
C1008 VN.n59 VSUBS 0.028634f
C1009 VN.n60 VSUBS 0.039993f
C1010 VN.n61 VSUBS 0.028634f
C1011 VN.t1 VSUBS 2.02839f
C1012 VN.n62 VSUBS 0.733107f
C1013 VN.n63 VSUBS 0.031181f
C1014 VN.n64 VSUBS 0.028634f
C1015 VN.n65 VSUBS 0.028459f
C1016 VN.t5 VSUBS 2.38746f
C1017 VN.t0 VSUBS 2.02839f
C1018 VN.n66 VSUBS 0.820369f
C1019 VN.n67 VSUBS 0.780492f
C1020 VN.n68 VSUBS 0.341468f
C1021 VN.n69 VSUBS 0.028634f
C1022 VN.n70 VSUBS 0.0531f
C1023 VN.n71 VSUBS 0.0531f
C1024 VN.n72 VSUBS 0.049952f
C1025 VN.n73 VSUBS 0.028634f
C1026 VN.n74 VSUBS 0.028634f
C1027 VN.n75 VSUBS 0.028634f
C1028 VN.n76 VSUBS 0.055215f
C1029 VN.n77 VSUBS 0.0531f
C1030 VN.n78 VSUBS 0.039993f
C1031 VN.n79 VSUBS 0.028634f
C1032 VN.n80 VSUBS 0.028634f
C1033 VN.n81 VSUBS 0.028634f
C1034 VN.n82 VSUBS 0.0531f
C1035 VN.n83 VSUBS 0.055215f
C1036 VN.n84 VSUBS 0.031181f
C1037 VN.n85 VSUBS 0.028634f
C1038 VN.n86 VSUBS 0.028634f
C1039 VN.n87 VSUBS 0.028634f
C1040 VN.n88 VSUBS 0.0531f
C1041 VN.n89 VSUBS 0.0531f
C1042 VN.n90 VSUBS 0.028459f
C1043 VN.n91 VSUBS 0.028634f
C1044 VN.n92 VSUBS 0.028634f
C1045 VN.n93 VSUBS 0.051527f
C1046 VN.n94 VSUBS 0.0531f
C1047 VN.n95 VSUBS 0.053357f
C1048 VN.n96 VSUBS 0.028634f
C1049 VN.n97 VSUBS 0.028634f
C1050 VN.n98 VSUBS 0.028634f
C1051 VN.n99 VSUBS 0.05744f
C1052 VN.n100 VSUBS 0.0531f
C1053 VN.n101 VSUBS 0.043138f
C1054 VN.n102 VSUBS 0.046208f
C1055 VN.n103 VSUBS 1.85867f
C1056 VDD1.t4 VSUBS 1.96653f
C1057 VDD1.t8 VSUBS 0.203086f
C1058 VDD1.t2 VSUBS 0.203086f
C1059 VDD1.n0 VSUBS 1.46186f
C1060 VDD1.n1 VSUBS 1.97343f
C1061 VDD1.t9 VSUBS 1.96653f
C1062 VDD1.t1 VSUBS 0.203086f
C1063 VDD1.t3 VSUBS 0.203086f
C1064 VDD1.n2 VSUBS 1.46185f
C1065 VDD1.n3 VSUBS 1.96219f
C1066 VDD1.t5 VSUBS 0.203086f
C1067 VDD1.t0 VSUBS 0.203086f
C1068 VDD1.n4 VSUBS 1.49311f
C1069 VDD1.n5 VSUBS 4.60932f
C1070 VDD1.t6 VSUBS 0.203086f
C1071 VDD1.t7 VSUBS 0.203086f
C1072 VDD1.n6 VSUBS 1.46185f
C1073 VDD1.n7 VSUBS 4.56637f
C1074 VTAIL.t0 VSUBS 0.19607f
C1075 VTAIL.t9 VSUBS 0.19607f
C1076 VTAIL.n0 VSUBS 1.28694f
C1077 VTAIL.n1 VSUBS 1.09733f
C1078 VTAIL.t17 VSUBS 1.73016f
C1079 VTAIL.n2 VSUBS 1.26781f
C1080 VTAIL.t13 VSUBS 0.19607f
C1081 VTAIL.t14 VSUBS 0.19607f
C1082 VTAIL.n3 VSUBS 1.28694f
C1083 VTAIL.n4 VSUBS 1.2973f
C1084 VTAIL.t16 VSUBS 0.19607f
C1085 VTAIL.t10 VSUBS 0.19607f
C1086 VTAIL.n5 VSUBS 1.28694f
C1087 VTAIL.n6 VSUBS 2.76662f
C1088 VTAIL.t2 VSUBS 0.19607f
C1089 VTAIL.t4 VSUBS 0.19607f
C1090 VTAIL.n7 VSUBS 1.28695f
C1091 VTAIL.n8 VSUBS 2.76662f
C1092 VTAIL.t5 VSUBS 0.19607f
C1093 VTAIL.t8 VSUBS 0.19607f
C1094 VTAIL.n9 VSUBS 1.28695f
C1095 VTAIL.n10 VSUBS 1.2973f
C1096 VTAIL.t1 VSUBS 1.73016f
C1097 VTAIL.n11 VSUBS 1.2678f
C1098 VTAIL.t19 VSUBS 0.19607f
C1099 VTAIL.t11 VSUBS 0.19607f
C1100 VTAIL.n12 VSUBS 1.28695f
C1101 VTAIL.n13 VSUBS 1.17628f
C1102 VTAIL.t18 VSUBS 0.19607f
C1103 VTAIL.t15 VSUBS 0.19607f
C1104 VTAIL.n14 VSUBS 1.28695f
C1105 VTAIL.n15 VSUBS 1.2973f
C1106 VTAIL.t12 VSUBS 1.73016f
C1107 VTAIL.n16 VSUBS 2.51804f
C1108 VTAIL.t3 VSUBS 1.73016f
C1109 VTAIL.n17 VSUBS 2.51804f
C1110 VTAIL.t7 VSUBS 0.19607f
C1111 VTAIL.t6 VSUBS 0.19607f
C1112 VTAIL.n18 VSUBS 1.28694f
C1113 VTAIL.n19 VSUBS 1.03615f
C1114 VP.t9 VSUBS 2.25194f
C1115 VP.n0 VSUBS 0.94434f
C1116 VP.n1 VSUBS 0.03179f
C1117 VP.n2 VSUBS 0.028368f
C1118 VP.n3 VSUBS 0.03179f
C1119 VP.t4 VSUBS 2.25194f
C1120 VP.n4 VSUBS 0.813902f
C1121 VP.n5 VSUBS 0.03179f
C1122 VP.n6 VSUBS 0.055457f
C1123 VP.n7 VSUBS 0.03179f
C1124 VP.n8 VSUBS 0.0444f
C1125 VP.n9 VSUBS 0.03179f
C1126 VP.n10 VSUBS 0.034618f
C1127 VP.n11 VSUBS 0.03179f
C1128 VP.n12 VSUBS 0.031595f
C1129 VP.n13 VSUBS 0.03179f
C1130 VP.n14 VSUBS 0.028368f
C1131 VP.n15 VSUBS 0.03179f
C1132 VP.t0 VSUBS 2.25194f
C1133 VP.n16 VSUBS 0.94434f
C1134 VP.t2 VSUBS 2.25194f
C1135 VP.n17 VSUBS 0.94434f
C1136 VP.n18 VSUBS 0.03179f
C1137 VP.n19 VSUBS 0.028368f
C1138 VP.n20 VSUBS 0.03179f
C1139 VP.t3 VSUBS 2.25194f
C1140 VP.n21 VSUBS 0.813902f
C1141 VP.n22 VSUBS 0.03179f
C1142 VP.n23 VSUBS 0.055457f
C1143 VP.n24 VSUBS 0.03179f
C1144 VP.n25 VSUBS 0.0444f
C1145 VP.n26 VSUBS 0.03179f
C1146 VP.n27 VSUBS 0.034618f
C1147 VP.n28 VSUBS 0.03179f
C1148 VP.n29 VSUBS 0.031595f
C1149 VP.t5 VSUBS 2.65058f
C1150 VP.t1 VSUBS 2.25194f
C1151 VP.n30 VSUBS 0.910782f
C1152 VP.n31 VSUBS 0.866511f
C1153 VP.n32 VSUBS 0.379102f
C1154 VP.n33 VSUBS 0.03179f
C1155 VP.n34 VSUBS 0.058952f
C1156 VP.n35 VSUBS 0.058952f
C1157 VP.n36 VSUBS 0.055457f
C1158 VP.n37 VSUBS 0.03179f
C1159 VP.n38 VSUBS 0.03179f
C1160 VP.n39 VSUBS 0.03179f
C1161 VP.n40 VSUBS 0.0613f
C1162 VP.n41 VSUBS 0.058952f
C1163 VP.t7 VSUBS 2.25194f
C1164 VP.n42 VSUBS 0.813902f
C1165 VP.n43 VSUBS 0.0444f
C1166 VP.n44 VSUBS 0.03179f
C1167 VP.n45 VSUBS 0.03179f
C1168 VP.n46 VSUBS 0.03179f
C1169 VP.n47 VSUBS 0.058952f
C1170 VP.n48 VSUBS 0.0613f
C1171 VP.n49 VSUBS 0.034618f
C1172 VP.n50 VSUBS 0.03179f
C1173 VP.n51 VSUBS 0.03179f
C1174 VP.n52 VSUBS 0.03179f
C1175 VP.n53 VSUBS 0.058952f
C1176 VP.n54 VSUBS 0.058952f
C1177 VP.n55 VSUBS 0.031595f
C1178 VP.n56 VSUBS 0.03179f
C1179 VP.n57 VSUBS 0.03179f
C1180 VP.n58 VSUBS 0.057206f
C1181 VP.n59 VSUBS 0.058952f
C1182 VP.n60 VSUBS 0.059238f
C1183 VP.n61 VSUBS 0.03179f
C1184 VP.n62 VSUBS 0.03179f
C1185 VP.n63 VSUBS 0.03179f
C1186 VP.n64 VSUBS 0.06377f
C1187 VP.n65 VSUBS 0.058952f
C1188 VP.n66 VSUBS 0.047893f
C1189 VP.n67 VSUBS 0.0513f
C1190 VP.n68 VSUBS 2.05089f
C1191 VP.n69 VSUBS 2.07188f
C1192 VP.n70 VSUBS 0.0513f
C1193 VP.n71 VSUBS 0.047893f
C1194 VP.n72 VSUBS 0.058952f
C1195 VP.n73 VSUBS 0.06377f
C1196 VP.n74 VSUBS 0.03179f
C1197 VP.n75 VSUBS 0.03179f
C1198 VP.n76 VSUBS 0.03179f
C1199 VP.n77 VSUBS 0.059238f
C1200 VP.n78 VSUBS 0.058952f
C1201 VP.t8 VSUBS 2.25194f
C1202 VP.n79 VSUBS 0.813902f
C1203 VP.n80 VSUBS 0.057206f
C1204 VP.n81 VSUBS 0.03179f
C1205 VP.n82 VSUBS 0.03179f
C1206 VP.n83 VSUBS 0.03179f
C1207 VP.n84 VSUBS 0.058952f
C1208 VP.n85 VSUBS 0.058952f
C1209 VP.n86 VSUBS 0.055457f
C1210 VP.n87 VSUBS 0.03179f
C1211 VP.n88 VSUBS 0.03179f
C1212 VP.n89 VSUBS 0.03179f
C1213 VP.n90 VSUBS 0.0613f
C1214 VP.n91 VSUBS 0.058952f
C1215 VP.t6 VSUBS 2.25194f
C1216 VP.n92 VSUBS 0.813902f
C1217 VP.n93 VSUBS 0.0444f
C1218 VP.n94 VSUBS 0.03179f
C1219 VP.n95 VSUBS 0.03179f
C1220 VP.n96 VSUBS 0.03179f
C1221 VP.n97 VSUBS 0.058952f
C1222 VP.n98 VSUBS 0.0613f
C1223 VP.n99 VSUBS 0.034618f
C1224 VP.n100 VSUBS 0.03179f
C1225 VP.n101 VSUBS 0.03179f
C1226 VP.n102 VSUBS 0.03179f
C1227 VP.n103 VSUBS 0.058952f
C1228 VP.n104 VSUBS 0.058952f
C1229 VP.n105 VSUBS 0.031595f
C1230 VP.n106 VSUBS 0.03179f
C1231 VP.n107 VSUBS 0.03179f
C1232 VP.n108 VSUBS 0.057206f
C1233 VP.n109 VSUBS 0.058952f
C1234 VP.n110 VSUBS 0.059238f
C1235 VP.n111 VSUBS 0.03179f
C1236 VP.n112 VSUBS 0.03179f
C1237 VP.n113 VSUBS 0.03179f
C1238 VP.n114 VSUBS 0.06377f
C1239 VP.n115 VSUBS 0.058952f
C1240 VP.n116 VSUBS 0.047893f
C1241 VP.n117 VSUBS 0.0513f
C1242 VP.n118 VSUBS 0.078141f
.ends

