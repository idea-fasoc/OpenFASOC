* NGSPICE file created from diff_pair_sample_0834.ext - technology: sky130A

.subckt diff_pair_sample_0834 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X1 VTAIL.t5 VN.t0 VDD2.t7 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=1.50315 ps=9.44 w=9.11 l=3.99
X2 VTAIL.t14 VP.t1 VDD1.t3 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X3 B.t11 B.t9 B.t10 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=0 ps=0 w=9.11 l=3.99
X4 B.t8 B.t6 B.t7 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=0 ps=0 w=9.11 l=3.99
X5 VDD2.t6 VN.t1 VTAIL.t2 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X6 B.t5 B.t3 B.t4 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=0 ps=0 w=9.11 l=3.99
X7 VTAIL.t13 VP.t2 VDD1.t6 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=1.50315 ps=9.44 w=9.11 l=3.99
X8 VDD1.t5 VP.t3 VTAIL.t12 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=3.5529 ps=19 w=9.11 l=3.99
X9 VDD2.t5 VN.t2 VTAIL.t4 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=3.5529 ps=19 w=9.11 l=3.99
X10 B.t2 B.t0 B.t1 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=0 ps=0 w=9.11 l=3.99
X11 VDD2.t4 VN.t3 VTAIL.t6 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X12 VDD1.t1 VP.t4 VTAIL.t11 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X13 VDD1.t7 VP.t5 VTAIL.t10 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X14 VDD2.t3 VN.t4 VTAIL.t7 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=3.5529 ps=19 w=9.11 l=3.99
X15 VTAIL.t0 VN.t5 VDD2.t2 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
X16 VTAIL.t9 VP.t6 VDD1.t4 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=1.50315 ps=9.44 w=9.11 l=3.99
X17 VTAIL.t3 VN.t6 VDD2.t1 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=3.5529 pd=19 as=1.50315 ps=9.44 w=9.11 l=3.99
X18 VDD1.t2 VP.t7 VTAIL.t8 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=3.5529 ps=19 w=9.11 l=3.99
X19 VTAIL.t1 VN.t7 VDD2.t0 w_n5290_n2790# sky130_fd_pr__pfet_01v8 ad=1.50315 pd=9.44 as=1.50315 ps=9.44 w=9.11 l=3.99
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n13 161.3
R17 VP.n92 VP.n0 161.3
R18 VP.n91 VP.n90 161.3
R19 VP.n89 VP.n1 161.3
R20 VP.n88 VP.n87 161.3
R21 VP.n86 VP.n2 161.3
R22 VP.n85 VP.n84 161.3
R23 VP.n83 VP.n3 161.3
R24 VP.n82 VP.n81 161.3
R25 VP.n79 VP.n4 161.3
R26 VP.n78 VP.n77 161.3
R27 VP.n76 VP.n5 161.3
R28 VP.n75 VP.n74 161.3
R29 VP.n73 VP.n6 161.3
R30 VP.n72 VP.n71 161.3
R31 VP.n70 VP.n7 161.3
R32 VP.n69 VP.n68 161.3
R33 VP.n67 VP.n8 161.3
R34 VP.n65 VP.n64 161.3
R35 VP.n63 VP.n9 161.3
R36 VP.n62 VP.n61 161.3
R37 VP.n60 VP.n10 161.3
R38 VP.n59 VP.n58 161.3
R39 VP.n57 VP.n11 161.3
R40 VP.n56 VP.n55 161.3
R41 VP.n54 VP.n12 161.3
R42 VP.n22 VP.t6 87.0715
R43 VP.n23 VP.n22 67.3497
R44 VP.n53 VP.n52 58.6935
R45 VP.n94 VP.n93 58.6935
R46 VP.n51 VP.n50 58.6935
R47 VP.n60 VP.n59 56.5193
R48 VP.n44 VP.n43 56.5193
R49 VP.n87 VP.n86 56.5193
R50 VP.n52 VP.n51 55.504
R51 VP.n53 VP.t2 55.0258
R52 VP.n66 VP.t4 55.0258
R53 VP.n80 VP.t1 55.0258
R54 VP.n93 VP.t3 55.0258
R55 VP.n50 VP.t7 55.0258
R56 VP.n37 VP.t0 55.0258
R57 VP.n23 VP.t5 55.0258
R58 VP.n73 VP.n72 40.4934
R59 VP.n74 VP.n73 40.4934
R60 VP.n31 VP.n30 40.4934
R61 VP.n30 VP.n29 40.4934
R62 VP.n55 VP.n54 24.4675
R63 VP.n55 VP.n11 24.4675
R64 VP.n59 VP.n11 24.4675
R65 VP.n61 VP.n60 24.4675
R66 VP.n61 VP.n9 24.4675
R67 VP.n65 VP.n9 24.4675
R68 VP.n68 VP.n67 24.4675
R69 VP.n68 VP.n7 24.4675
R70 VP.n72 VP.n7 24.4675
R71 VP.n74 VP.n5 24.4675
R72 VP.n78 VP.n5 24.4675
R73 VP.n79 VP.n78 24.4675
R74 VP.n81 VP.n3 24.4675
R75 VP.n85 VP.n3 24.4675
R76 VP.n86 VP.n85 24.4675
R77 VP.n87 VP.n1 24.4675
R78 VP.n91 VP.n1 24.4675
R79 VP.n92 VP.n91 24.4675
R80 VP.n44 VP.n14 24.4675
R81 VP.n48 VP.n14 24.4675
R82 VP.n49 VP.n48 24.4675
R83 VP.n31 VP.n18 24.4675
R84 VP.n35 VP.n18 24.4675
R85 VP.n36 VP.n35 24.4675
R86 VP.n38 VP.n16 24.4675
R87 VP.n42 VP.n16 24.4675
R88 VP.n43 VP.n42 24.4675
R89 VP.n25 VP.n24 24.4675
R90 VP.n25 VP.n20 24.4675
R91 VP.n29 VP.n20 24.4675
R92 VP.n54 VP.n53 23.4888
R93 VP.n93 VP.n92 23.4888
R94 VP.n50 VP.n49 23.4888
R95 VP.n66 VP.n65 16.6381
R96 VP.n81 VP.n80 16.6381
R97 VP.n38 VP.n37 16.6381
R98 VP.n67 VP.n66 7.82994
R99 VP.n80 VP.n79 7.82994
R100 VP.n37 VP.n36 7.82994
R101 VP.n24 VP.n23 7.82994
R102 VP.n22 VP.n21 2.57369
R103 VP.n51 VP.n13 0.417535
R104 VP.n52 VP.n12 0.417535
R105 VP.n94 VP.n0 0.417535
R106 VP VP.n94 0.394291
R107 VP.n26 VP.n21 0.189894
R108 VP.n27 VP.n26 0.189894
R109 VP.n28 VP.n27 0.189894
R110 VP.n28 VP.n19 0.189894
R111 VP.n32 VP.n19 0.189894
R112 VP.n33 VP.n32 0.189894
R113 VP.n34 VP.n33 0.189894
R114 VP.n34 VP.n17 0.189894
R115 VP.n39 VP.n17 0.189894
R116 VP.n40 VP.n39 0.189894
R117 VP.n41 VP.n40 0.189894
R118 VP.n41 VP.n15 0.189894
R119 VP.n45 VP.n15 0.189894
R120 VP.n46 VP.n45 0.189894
R121 VP.n47 VP.n46 0.189894
R122 VP.n47 VP.n13 0.189894
R123 VP.n56 VP.n12 0.189894
R124 VP.n57 VP.n56 0.189894
R125 VP.n58 VP.n57 0.189894
R126 VP.n58 VP.n10 0.189894
R127 VP.n62 VP.n10 0.189894
R128 VP.n63 VP.n62 0.189894
R129 VP.n64 VP.n63 0.189894
R130 VP.n64 VP.n8 0.189894
R131 VP.n69 VP.n8 0.189894
R132 VP.n70 VP.n69 0.189894
R133 VP.n71 VP.n70 0.189894
R134 VP.n71 VP.n6 0.189894
R135 VP.n75 VP.n6 0.189894
R136 VP.n76 VP.n75 0.189894
R137 VP.n77 VP.n76 0.189894
R138 VP.n77 VP.n4 0.189894
R139 VP.n82 VP.n4 0.189894
R140 VP.n83 VP.n82 0.189894
R141 VP.n84 VP.n83 0.189894
R142 VP.n84 VP.n2 0.189894
R143 VP.n88 VP.n2 0.189894
R144 VP.n89 VP.n88 0.189894
R145 VP.n90 VP.n89 0.189894
R146 VP.n90 VP.n0 0.189894
R147 VDD1 VDD1.n0 85.7864
R148 VDD1.n3 VDD1.n2 85.6726
R149 VDD1.n3 VDD1.n1 85.6726
R150 VDD1.n5 VDD1.n4 83.866
R151 VDD1.n5 VDD1.n3 48.9104
R152 VDD1.n4 VDD1.t0 3.56856
R153 VDD1.n4 VDD1.t2 3.56856
R154 VDD1.n0 VDD1.t4 3.56856
R155 VDD1.n0 VDD1.t7 3.56856
R156 VDD1.n2 VDD1.t3 3.56856
R157 VDD1.n2 VDD1.t5 3.56856
R158 VDD1.n1 VDD1.t6 3.56856
R159 VDD1.n1 VDD1.t1 3.56856
R160 VDD1 VDD1.n5 1.80438
R161 VTAIL.n11 VTAIL.t9 70.7554
R162 VTAIL.n10 VTAIL.t4 70.7554
R163 VTAIL.n7 VTAIL.t5 70.7554
R164 VTAIL.n15 VTAIL.t7 70.7551
R165 VTAIL.n2 VTAIL.t3 70.7551
R166 VTAIL.n3 VTAIL.t12 70.7551
R167 VTAIL.n6 VTAIL.t13 70.7551
R168 VTAIL.n14 VTAIL.t8 70.7551
R169 VTAIL.n13 VTAIL.n12 67.1874
R170 VTAIL.n9 VTAIL.n8 67.1874
R171 VTAIL.n1 VTAIL.n0 67.1871
R172 VTAIL.n5 VTAIL.n4 67.1871
R173 VTAIL.n15 VTAIL.n14 23.9445
R174 VTAIL.n7 VTAIL.n6 23.9445
R175 VTAIL.n9 VTAIL.n7 3.72464
R176 VTAIL.n10 VTAIL.n9 3.72464
R177 VTAIL.n13 VTAIL.n11 3.72464
R178 VTAIL.n14 VTAIL.n13 3.72464
R179 VTAIL.n6 VTAIL.n5 3.72464
R180 VTAIL.n5 VTAIL.n3 3.72464
R181 VTAIL.n2 VTAIL.n1 3.72464
R182 VTAIL VTAIL.n15 3.66645
R183 VTAIL.n0 VTAIL.t6 3.56856
R184 VTAIL.n0 VTAIL.t1 3.56856
R185 VTAIL.n4 VTAIL.t11 3.56856
R186 VTAIL.n4 VTAIL.t14 3.56856
R187 VTAIL.n12 VTAIL.t10 3.56856
R188 VTAIL.n12 VTAIL.t15 3.56856
R189 VTAIL.n8 VTAIL.t2 3.56856
R190 VTAIL.n8 VTAIL.t0 3.56856
R191 VTAIL.n11 VTAIL.n10 0.470328
R192 VTAIL.n3 VTAIL.n2 0.470328
R193 VTAIL VTAIL.n1 0.0586897
R194 VN.n75 VN.n39 161.3
R195 VN.n74 VN.n73 161.3
R196 VN.n72 VN.n40 161.3
R197 VN.n71 VN.n70 161.3
R198 VN.n69 VN.n41 161.3
R199 VN.n68 VN.n67 161.3
R200 VN.n66 VN.n42 161.3
R201 VN.n65 VN.n64 161.3
R202 VN.n62 VN.n43 161.3
R203 VN.n61 VN.n60 161.3
R204 VN.n59 VN.n44 161.3
R205 VN.n58 VN.n57 161.3
R206 VN.n56 VN.n45 161.3
R207 VN.n55 VN.n54 161.3
R208 VN.n53 VN.n46 161.3
R209 VN.n52 VN.n51 161.3
R210 VN.n50 VN.n47 161.3
R211 VN.n36 VN.n0 161.3
R212 VN.n35 VN.n34 161.3
R213 VN.n33 VN.n1 161.3
R214 VN.n32 VN.n31 161.3
R215 VN.n30 VN.n2 161.3
R216 VN.n29 VN.n28 161.3
R217 VN.n27 VN.n3 161.3
R218 VN.n26 VN.n25 161.3
R219 VN.n23 VN.n4 161.3
R220 VN.n22 VN.n21 161.3
R221 VN.n20 VN.n5 161.3
R222 VN.n19 VN.n18 161.3
R223 VN.n17 VN.n6 161.3
R224 VN.n16 VN.n15 161.3
R225 VN.n14 VN.n7 161.3
R226 VN.n13 VN.n12 161.3
R227 VN.n11 VN.n8 161.3
R228 VN.n9 VN.t6 87.072
R229 VN.n48 VN.t2 87.072
R230 VN.n10 VN.n9 67.3496
R231 VN.n49 VN.n48 67.3496
R232 VN.n38 VN.n37 58.6935
R233 VN.n77 VN.n76 58.6935
R234 VN.n31 VN.n30 56.5193
R235 VN.n70 VN.n69 56.5193
R236 VN VN.n77 55.542
R237 VN.n10 VN.t3 55.0258
R238 VN.n24 VN.t7 55.0258
R239 VN.n37 VN.t4 55.0258
R240 VN.n49 VN.t5 55.0258
R241 VN.n63 VN.t1 55.0258
R242 VN.n76 VN.t0 55.0258
R243 VN.n17 VN.n16 40.4934
R244 VN.n18 VN.n17 40.4934
R245 VN.n56 VN.n55 40.4934
R246 VN.n57 VN.n56 40.4934
R247 VN.n12 VN.n11 24.4675
R248 VN.n12 VN.n7 24.4675
R249 VN.n16 VN.n7 24.4675
R250 VN.n18 VN.n5 24.4675
R251 VN.n22 VN.n5 24.4675
R252 VN.n23 VN.n22 24.4675
R253 VN.n25 VN.n3 24.4675
R254 VN.n29 VN.n3 24.4675
R255 VN.n30 VN.n29 24.4675
R256 VN.n31 VN.n1 24.4675
R257 VN.n35 VN.n1 24.4675
R258 VN.n36 VN.n35 24.4675
R259 VN.n55 VN.n46 24.4675
R260 VN.n51 VN.n46 24.4675
R261 VN.n51 VN.n50 24.4675
R262 VN.n69 VN.n68 24.4675
R263 VN.n68 VN.n42 24.4675
R264 VN.n64 VN.n42 24.4675
R265 VN.n62 VN.n61 24.4675
R266 VN.n61 VN.n44 24.4675
R267 VN.n57 VN.n44 24.4675
R268 VN.n75 VN.n74 24.4675
R269 VN.n74 VN.n40 24.4675
R270 VN.n70 VN.n40 24.4675
R271 VN.n37 VN.n36 23.4888
R272 VN.n76 VN.n75 23.4888
R273 VN.n25 VN.n24 16.6381
R274 VN.n64 VN.n63 16.6381
R275 VN.n11 VN.n10 7.82994
R276 VN.n24 VN.n23 7.82994
R277 VN.n50 VN.n49 7.82994
R278 VN.n63 VN.n62 7.82994
R279 VN.n48 VN.n47 2.57372
R280 VN.n9 VN.n8 2.57372
R281 VN.n77 VN.n39 0.417535
R282 VN.n38 VN.n0 0.417535
R283 VN VN.n38 0.394291
R284 VN.n73 VN.n39 0.189894
R285 VN.n73 VN.n72 0.189894
R286 VN.n72 VN.n71 0.189894
R287 VN.n71 VN.n41 0.189894
R288 VN.n67 VN.n41 0.189894
R289 VN.n67 VN.n66 0.189894
R290 VN.n66 VN.n65 0.189894
R291 VN.n65 VN.n43 0.189894
R292 VN.n60 VN.n43 0.189894
R293 VN.n60 VN.n59 0.189894
R294 VN.n59 VN.n58 0.189894
R295 VN.n58 VN.n45 0.189894
R296 VN.n54 VN.n45 0.189894
R297 VN.n54 VN.n53 0.189894
R298 VN.n53 VN.n52 0.189894
R299 VN.n52 VN.n47 0.189894
R300 VN.n13 VN.n8 0.189894
R301 VN.n14 VN.n13 0.189894
R302 VN.n15 VN.n14 0.189894
R303 VN.n15 VN.n6 0.189894
R304 VN.n19 VN.n6 0.189894
R305 VN.n20 VN.n19 0.189894
R306 VN.n21 VN.n20 0.189894
R307 VN.n21 VN.n4 0.189894
R308 VN.n26 VN.n4 0.189894
R309 VN.n27 VN.n26 0.189894
R310 VN.n28 VN.n27 0.189894
R311 VN.n28 VN.n2 0.189894
R312 VN.n32 VN.n2 0.189894
R313 VN.n33 VN.n32 0.189894
R314 VN.n34 VN.n33 0.189894
R315 VN.n34 VN.n0 0.189894
R316 VDD2.n2 VDD2.n1 85.6726
R317 VDD2.n2 VDD2.n0 85.6726
R318 VDD2 VDD2.n5 85.6698
R319 VDD2.n4 VDD2.n3 83.8661
R320 VDD2.n4 VDD2.n2 48.3274
R321 VDD2.n5 VDD2.t2 3.56856
R322 VDD2.n5 VDD2.t5 3.56856
R323 VDD2.n3 VDD2.t7 3.56856
R324 VDD2.n3 VDD2.t6 3.56856
R325 VDD2.n1 VDD2.t0 3.56856
R326 VDD2.n1 VDD2.t3 3.56856
R327 VDD2.n0 VDD2.t1 3.56856
R328 VDD2.n0 VDD2.t4 3.56856
R329 VDD2 VDD2.n4 1.92076
R330 B.n449 B.n152 585
R331 B.n448 B.n447 585
R332 B.n446 B.n153 585
R333 B.n445 B.n444 585
R334 B.n443 B.n154 585
R335 B.n442 B.n441 585
R336 B.n440 B.n155 585
R337 B.n439 B.n438 585
R338 B.n437 B.n156 585
R339 B.n436 B.n435 585
R340 B.n434 B.n157 585
R341 B.n433 B.n432 585
R342 B.n431 B.n158 585
R343 B.n430 B.n429 585
R344 B.n428 B.n159 585
R345 B.n427 B.n426 585
R346 B.n425 B.n160 585
R347 B.n424 B.n423 585
R348 B.n422 B.n161 585
R349 B.n421 B.n420 585
R350 B.n419 B.n162 585
R351 B.n418 B.n417 585
R352 B.n416 B.n163 585
R353 B.n415 B.n414 585
R354 B.n413 B.n164 585
R355 B.n412 B.n411 585
R356 B.n410 B.n165 585
R357 B.n409 B.n408 585
R358 B.n407 B.n166 585
R359 B.n406 B.n405 585
R360 B.n404 B.n167 585
R361 B.n403 B.n402 585
R362 B.n401 B.n168 585
R363 B.n400 B.n399 585
R364 B.n395 B.n169 585
R365 B.n394 B.n393 585
R366 B.n392 B.n170 585
R367 B.n391 B.n390 585
R368 B.n389 B.n171 585
R369 B.n388 B.n387 585
R370 B.n386 B.n172 585
R371 B.n385 B.n384 585
R372 B.n383 B.n173 585
R373 B.n381 B.n380 585
R374 B.n379 B.n176 585
R375 B.n378 B.n377 585
R376 B.n376 B.n177 585
R377 B.n375 B.n374 585
R378 B.n373 B.n178 585
R379 B.n372 B.n371 585
R380 B.n370 B.n179 585
R381 B.n369 B.n368 585
R382 B.n367 B.n180 585
R383 B.n366 B.n365 585
R384 B.n364 B.n181 585
R385 B.n363 B.n362 585
R386 B.n361 B.n182 585
R387 B.n360 B.n359 585
R388 B.n358 B.n183 585
R389 B.n357 B.n356 585
R390 B.n355 B.n184 585
R391 B.n354 B.n353 585
R392 B.n352 B.n185 585
R393 B.n351 B.n350 585
R394 B.n349 B.n186 585
R395 B.n348 B.n347 585
R396 B.n346 B.n187 585
R397 B.n345 B.n344 585
R398 B.n343 B.n188 585
R399 B.n342 B.n341 585
R400 B.n340 B.n189 585
R401 B.n339 B.n338 585
R402 B.n337 B.n190 585
R403 B.n336 B.n335 585
R404 B.n334 B.n191 585
R405 B.n333 B.n332 585
R406 B.n451 B.n450 585
R407 B.n452 B.n151 585
R408 B.n454 B.n453 585
R409 B.n455 B.n150 585
R410 B.n457 B.n456 585
R411 B.n458 B.n149 585
R412 B.n460 B.n459 585
R413 B.n461 B.n148 585
R414 B.n463 B.n462 585
R415 B.n464 B.n147 585
R416 B.n466 B.n465 585
R417 B.n467 B.n146 585
R418 B.n469 B.n468 585
R419 B.n470 B.n145 585
R420 B.n472 B.n471 585
R421 B.n473 B.n144 585
R422 B.n475 B.n474 585
R423 B.n476 B.n143 585
R424 B.n478 B.n477 585
R425 B.n479 B.n142 585
R426 B.n481 B.n480 585
R427 B.n482 B.n141 585
R428 B.n484 B.n483 585
R429 B.n485 B.n140 585
R430 B.n487 B.n486 585
R431 B.n488 B.n139 585
R432 B.n490 B.n489 585
R433 B.n491 B.n138 585
R434 B.n493 B.n492 585
R435 B.n494 B.n137 585
R436 B.n496 B.n495 585
R437 B.n497 B.n136 585
R438 B.n499 B.n498 585
R439 B.n500 B.n135 585
R440 B.n502 B.n501 585
R441 B.n503 B.n134 585
R442 B.n505 B.n504 585
R443 B.n506 B.n133 585
R444 B.n508 B.n507 585
R445 B.n509 B.n132 585
R446 B.n511 B.n510 585
R447 B.n512 B.n131 585
R448 B.n514 B.n513 585
R449 B.n515 B.n130 585
R450 B.n517 B.n516 585
R451 B.n518 B.n129 585
R452 B.n520 B.n519 585
R453 B.n521 B.n128 585
R454 B.n523 B.n522 585
R455 B.n524 B.n127 585
R456 B.n526 B.n525 585
R457 B.n527 B.n126 585
R458 B.n529 B.n528 585
R459 B.n530 B.n125 585
R460 B.n532 B.n531 585
R461 B.n533 B.n124 585
R462 B.n535 B.n534 585
R463 B.n536 B.n123 585
R464 B.n538 B.n537 585
R465 B.n539 B.n122 585
R466 B.n541 B.n540 585
R467 B.n542 B.n121 585
R468 B.n544 B.n543 585
R469 B.n545 B.n120 585
R470 B.n547 B.n546 585
R471 B.n548 B.n119 585
R472 B.n550 B.n549 585
R473 B.n551 B.n118 585
R474 B.n553 B.n552 585
R475 B.n554 B.n117 585
R476 B.n556 B.n555 585
R477 B.n557 B.n116 585
R478 B.n559 B.n558 585
R479 B.n560 B.n115 585
R480 B.n562 B.n561 585
R481 B.n563 B.n114 585
R482 B.n565 B.n564 585
R483 B.n566 B.n113 585
R484 B.n568 B.n567 585
R485 B.n569 B.n112 585
R486 B.n571 B.n570 585
R487 B.n572 B.n111 585
R488 B.n574 B.n573 585
R489 B.n575 B.n110 585
R490 B.n577 B.n576 585
R491 B.n578 B.n109 585
R492 B.n580 B.n579 585
R493 B.n581 B.n108 585
R494 B.n583 B.n582 585
R495 B.n584 B.n107 585
R496 B.n586 B.n585 585
R497 B.n587 B.n106 585
R498 B.n589 B.n588 585
R499 B.n590 B.n105 585
R500 B.n592 B.n591 585
R501 B.n593 B.n104 585
R502 B.n595 B.n594 585
R503 B.n596 B.n103 585
R504 B.n598 B.n597 585
R505 B.n599 B.n102 585
R506 B.n601 B.n600 585
R507 B.n602 B.n101 585
R508 B.n604 B.n603 585
R509 B.n605 B.n100 585
R510 B.n607 B.n606 585
R511 B.n608 B.n99 585
R512 B.n610 B.n609 585
R513 B.n611 B.n98 585
R514 B.n613 B.n612 585
R515 B.n614 B.n97 585
R516 B.n616 B.n615 585
R517 B.n617 B.n96 585
R518 B.n619 B.n618 585
R519 B.n620 B.n95 585
R520 B.n622 B.n621 585
R521 B.n623 B.n94 585
R522 B.n625 B.n624 585
R523 B.n626 B.n93 585
R524 B.n628 B.n627 585
R525 B.n629 B.n92 585
R526 B.n631 B.n630 585
R527 B.n632 B.n91 585
R528 B.n634 B.n633 585
R529 B.n635 B.n90 585
R530 B.n637 B.n636 585
R531 B.n638 B.n89 585
R532 B.n640 B.n639 585
R533 B.n641 B.n88 585
R534 B.n643 B.n642 585
R535 B.n644 B.n87 585
R536 B.n646 B.n645 585
R537 B.n647 B.n86 585
R538 B.n649 B.n648 585
R539 B.n650 B.n85 585
R540 B.n652 B.n651 585
R541 B.n653 B.n84 585
R542 B.n655 B.n654 585
R543 B.n656 B.n83 585
R544 B.n658 B.n657 585
R545 B.n659 B.n82 585
R546 B.n661 B.n660 585
R547 B.n662 B.n81 585
R548 B.n664 B.n663 585
R549 B.n665 B.n80 585
R550 B.n781 B.n780 585
R551 B.n779 B.n38 585
R552 B.n778 B.n777 585
R553 B.n776 B.n39 585
R554 B.n775 B.n774 585
R555 B.n773 B.n40 585
R556 B.n772 B.n771 585
R557 B.n770 B.n41 585
R558 B.n769 B.n768 585
R559 B.n767 B.n42 585
R560 B.n766 B.n765 585
R561 B.n764 B.n43 585
R562 B.n763 B.n762 585
R563 B.n761 B.n44 585
R564 B.n760 B.n759 585
R565 B.n758 B.n45 585
R566 B.n757 B.n756 585
R567 B.n755 B.n46 585
R568 B.n754 B.n753 585
R569 B.n752 B.n47 585
R570 B.n751 B.n750 585
R571 B.n749 B.n48 585
R572 B.n748 B.n747 585
R573 B.n746 B.n49 585
R574 B.n745 B.n744 585
R575 B.n743 B.n50 585
R576 B.n742 B.n741 585
R577 B.n740 B.n51 585
R578 B.n739 B.n738 585
R579 B.n737 B.n52 585
R580 B.n736 B.n735 585
R581 B.n734 B.n53 585
R582 B.n733 B.n732 585
R583 B.n731 B.n730 585
R584 B.n729 B.n57 585
R585 B.n728 B.n727 585
R586 B.n726 B.n58 585
R587 B.n725 B.n724 585
R588 B.n723 B.n59 585
R589 B.n722 B.n721 585
R590 B.n720 B.n60 585
R591 B.n719 B.n718 585
R592 B.n717 B.n61 585
R593 B.n715 B.n714 585
R594 B.n713 B.n64 585
R595 B.n712 B.n711 585
R596 B.n710 B.n65 585
R597 B.n709 B.n708 585
R598 B.n707 B.n66 585
R599 B.n706 B.n705 585
R600 B.n704 B.n67 585
R601 B.n703 B.n702 585
R602 B.n701 B.n68 585
R603 B.n700 B.n699 585
R604 B.n698 B.n69 585
R605 B.n697 B.n696 585
R606 B.n695 B.n70 585
R607 B.n694 B.n693 585
R608 B.n692 B.n71 585
R609 B.n691 B.n690 585
R610 B.n689 B.n72 585
R611 B.n688 B.n687 585
R612 B.n686 B.n73 585
R613 B.n685 B.n684 585
R614 B.n683 B.n74 585
R615 B.n682 B.n681 585
R616 B.n680 B.n75 585
R617 B.n679 B.n678 585
R618 B.n677 B.n76 585
R619 B.n676 B.n675 585
R620 B.n674 B.n77 585
R621 B.n673 B.n672 585
R622 B.n671 B.n78 585
R623 B.n670 B.n669 585
R624 B.n668 B.n79 585
R625 B.n667 B.n666 585
R626 B.n782 B.n37 585
R627 B.n784 B.n783 585
R628 B.n785 B.n36 585
R629 B.n787 B.n786 585
R630 B.n788 B.n35 585
R631 B.n790 B.n789 585
R632 B.n791 B.n34 585
R633 B.n793 B.n792 585
R634 B.n794 B.n33 585
R635 B.n796 B.n795 585
R636 B.n797 B.n32 585
R637 B.n799 B.n798 585
R638 B.n800 B.n31 585
R639 B.n802 B.n801 585
R640 B.n803 B.n30 585
R641 B.n805 B.n804 585
R642 B.n806 B.n29 585
R643 B.n808 B.n807 585
R644 B.n809 B.n28 585
R645 B.n811 B.n810 585
R646 B.n812 B.n27 585
R647 B.n814 B.n813 585
R648 B.n815 B.n26 585
R649 B.n817 B.n816 585
R650 B.n818 B.n25 585
R651 B.n820 B.n819 585
R652 B.n821 B.n24 585
R653 B.n823 B.n822 585
R654 B.n824 B.n23 585
R655 B.n826 B.n825 585
R656 B.n827 B.n22 585
R657 B.n829 B.n828 585
R658 B.n830 B.n21 585
R659 B.n832 B.n831 585
R660 B.n833 B.n20 585
R661 B.n835 B.n834 585
R662 B.n836 B.n19 585
R663 B.n838 B.n837 585
R664 B.n839 B.n18 585
R665 B.n841 B.n840 585
R666 B.n842 B.n17 585
R667 B.n844 B.n843 585
R668 B.n845 B.n16 585
R669 B.n847 B.n846 585
R670 B.n848 B.n15 585
R671 B.n850 B.n849 585
R672 B.n851 B.n14 585
R673 B.n853 B.n852 585
R674 B.n854 B.n13 585
R675 B.n856 B.n855 585
R676 B.n857 B.n12 585
R677 B.n859 B.n858 585
R678 B.n860 B.n11 585
R679 B.n862 B.n861 585
R680 B.n863 B.n10 585
R681 B.n865 B.n864 585
R682 B.n866 B.n9 585
R683 B.n868 B.n867 585
R684 B.n869 B.n8 585
R685 B.n871 B.n870 585
R686 B.n872 B.n7 585
R687 B.n874 B.n873 585
R688 B.n875 B.n6 585
R689 B.n877 B.n876 585
R690 B.n878 B.n5 585
R691 B.n880 B.n879 585
R692 B.n881 B.n4 585
R693 B.n883 B.n882 585
R694 B.n884 B.n3 585
R695 B.n886 B.n885 585
R696 B.n887 B.n0 585
R697 B.n2 B.n1 585
R698 B.n228 B.n227 585
R699 B.n229 B.n226 585
R700 B.n231 B.n230 585
R701 B.n232 B.n225 585
R702 B.n234 B.n233 585
R703 B.n235 B.n224 585
R704 B.n237 B.n236 585
R705 B.n238 B.n223 585
R706 B.n240 B.n239 585
R707 B.n241 B.n222 585
R708 B.n243 B.n242 585
R709 B.n244 B.n221 585
R710 B.n246 B.n245 585
R711 B.n247 B.n220 585
R712 B.n249 B.n248 585
R713 B.n250 B.n219 585
R714 B.n252 B.n251 585
R715 B.n253 B.n218 585
R716 B.n255 B.n254 585
R717 B.n256 B.n217 585
R718 B.n258 B.n257 585
R719 B.n259 B.n216 585
R720 B.n261 B.n260 585
R721 B.n262 B.n215 585
R722 B.n264 B.n263 585
R723 B.n265 B.n214 585
R724 B.n267 B.n266 585
R725 B.n268 B.n213 585
R726 B.n270 B.n269 585
R727 B.n271 B.n212 585
R728 B.n273 B.n272 585
R729 B.n274 B.n211 585
R730 B.n276 B.n275 585
R731 B.n277 B.n210 585
R732 B.n279 B.n278 585
R733 B.n280 B.n209 585
R734 B.n282 B.n281 585
R735 B.n283 B.n208 585
R736 B.n285 B.n284 585
R737 B.n286 B.n207 585
R738 B.n288 B.n287 585
R739 B.n289 B.n206 585
R740 B.n291 B.n290 585
R741 B.n292 B.n205 585
R742 B.n294 B.n293 585
R743 B.n295 B.n204 585
R744 B.n297 B.n296 585
R745 B.n298 B.n203 585
R746 B.n300 B.n299 585
R747 B.n301 B.n202 585
R748 B.n303 B.n302 585
R749 B.n304 B.n201 585
R750 B.n306 B.n305 585
R751 B.n307 B.n200 585
R752 B.n309 B.n308 585
R753 B.n310 B.n199 585
R754 B.n312 B.n311 585
R755 B.n313 B.n198 585
R756 B.n315 B.n314 585
R757 B.n316 B.n197 585
R758 B.n318 B.n317 585
R759 B.n319 B.n196 585
R760 B.n321 B.n320 585
R761 B.n322 B.n195 585
R762 B.n324 B.n323 585
R763 B.n325 B.n194 585
R764 B.n327 B.n326 585
R765 B.n328 B.n193 585
R766 B.n330 B.n329 585
R767 B.n331 B.n192 585
R768 B.n332 B.n331 506.916
R769 B.n450 B.n449 506.916
R770 B.n666 B.n665 506.916
R771 B.n780 B.n37 506.916
R772 B.n174 B.t6 264.51
R773 B.n396 B.t3 264.51
R774 B.n62 B.t9 264.51
R775 B.n54 B.t0 264.51
R776 B.n889 B.n888 256.663
R777 B.n888 B.n887 235.042
R778 B.n888 B.n2 235.042
R779 B.n396 B.t4 197.069
R780 B.n62 B.t11 197.069
R781 B.n174 B.t7 197.059
R782 B.n54 B.t2 197.059
R783 B.n332 B.n191 163.367
R784 B.n336 B.n191 163.367
R785 B.n337 B.n336 163.367
R786 B.n338 B.n337 163.367
R787 B.n338 B.n189 163.367
R788 B.n342 B.n189 163.367
R789 B.n343 B.n342 163.367
R790 B.n344 B.n343 163.367
R791 B.n344 B.n187 163.367
R792 B.n348 B.n187 163.367
R793 B.n349 B.n348 163.367
R794 B.n350 B.n349 163.367
R795 B.n350 B.n185 163.367
R796 B.n354 B.n185 163.367
R797 B.n355 B.n354 163.367
R798 B.n356 B.n355 163.367
R799 B.n356 B.n183 163.367
R800 B.n360 B.n183 163.367
R801 B.n361 B.n360 163.367
R802 B.n362 B.n361 163.367
R803 B.n362 B.n181 163.367
R804 B.n366 B.n181 163.367
R805 B.n367 B.n366 163.367
R806 B.n368 B.n367 163.367
R807 B.n368 B.n179 163.367
R808 B.n372 B.n179 163.367
R809 B.n373 B.n372 163.367
R810 B.n374 B.n373 163.367
R811 B.n374 B.n177 163.367
R812 B.n378 B.n177 163.367
R813 B.n379 B.n378 163.367
R814 B.n380 B.n379 163.367
R815 B.n380 B.n173 163.367
R816 B.n385 B.n173 163.367
R817 B.n386 B.n385 163.367
R818 B.n387 B.n386 163.367
R819 B.n387 B.n171 163.367
R820 B.n391 B.n171 163.367
R821 B.n392 B.n391 163.367
R822 B.n393 B.n392 163.367
R823 B.n393 B.n169 163.367
R824 B.n400 B.n169 163.367
R825 B.n401 B.n400 163.367
R826 B.n402 B.n401 163.367
R827 B.n402 B.n167 163.367
R828 B.n406 B.n167 163.367
R829 B.n407 B.n406 163.367
R830 B.n408 B.n407 163.367
R831 B.n408 B.n165 163.367
R832 B.n412 B.n165 163.367
R833 B.n413 B.n412 163.367
R834 B.n414 B.n413 163.367
R835 B.n414 B.n163 163.367
R836 B.n418 B.n163 163.367
R837 B.n419 B.n418 163.367
R838 B.n420 B.n419 163.367
R839 B.n420 B.n161 163.367
R840 B.n424 B.n161 163.367
R841 B.n425 B.n424 163.367
R842 B.n426 B.n425 163.367
R843 B.n426 B.n159 163.367
R844 B.n430 B.n159 163.367
R845 B.n431 B.n430 163.367
R846 B.n432 B.n431 163.367
R847 B.n432 B.n157 163.367
R848 B.n436 B.n157 163.367
R849 B.n437 B.n436 163.367
R850 B.n438 B.n437 163.367
R851 B.n438 B.n155 163.367
R852 B.n442 B.n155 163.367
R853 B.n443 B.n442 163.367
R854 B.n444 B.n443 163.367
R855 B.n444 B.n153 163.367
R856 B.n448 B.n153 163.367
R857 B.n449 B.n448 163.367
R858 B.n665 B.n664 163.367
R859 B.n664 B.n81 163.367
R860 B.n660 B.n81 163.367
R861 B.n660 B.n659 163.367
R862 B.n659 B.n658 163.367
R863 B.n658 B.n83 163.367
R864 B.n654 B.n83 163.367
R865 B.n654 B.n653 163.367
R866 B.n653 B.n652 163.367
R867 B.n652 B.n85 163.367
R868 B.n648 B.n85 163.367
R869 B.n648 B.n647 163.367
R870 B.n647 B.n646 163.367
R871 B.n646 B.n87 163.367
R872 B.n642 B.n87 163.367
R873 B.n642 B.n641 163.367
R874 B.n641 B.n640 163.367
R875 B.n640 B.n89 163.367
R876 B.n636 B.n89 163.367
R877 B.n636 B.n635 163.367
R878 B.n635 B.n634 163.367
R879 B.n634 B.n91 163.367
R880 B.n630 B.n91 163.367
R881 B.n630 B.n629 163.367
R882 B.n629 B.n628 163.367
R883 B.n628 B.n93 163.367
R884 B.n624 B.n93 163.367
R885 B.n624 B.n623 163.367
R886 B.n623 B.n622 163.367
R887 B.n622 B.n95 163.367
R888 B.n618 B.n95 163.367
R889 B.n618 B.n617 163.367
R890 B.n617 B.n616 163.367
R891 B.n616 B.n97 163.367
R892 B.n612 B.n97 163.367
R893 B.n612 B.n611 163.367
R894 B.n611 B.n610 163.367
R895 B.n610 B.n99 163.367
R896 B.n606 B.n99 163.367
R897 B.n606 B.n605 163.367
R898 B.n605 B.n604 163.367
R899 B.n604 B.n101 163.367
R900 B.n600 B.n101 163.367
R901 B.n600 B.n599 163.367
R902 B.n599 B.n598 163.367
R903 B.n598 B.n103 163.367
R904 B.n594 B.n103 163.367
R905 B.n594 B.n593 163.367
R906 B.n593 B.n592 163.367
R907 B.n592 B.n105 163.367
R908 B.n588 B.n105 163.367
R909 B.n588 B.n587 163.367
R910 B.n587 B.n586 163.367
R911 B.n586 B.n107 163.367
R912 B.n582 B.n107 163.367
R913 B.n582 B.n581 163.367
R914 B.n581 B.n580 163.367
R915 B.n580 B.n109 163.367
R916 B.n576 B.n109 163.367
R917 B.n576 B.n575 163.367
R918 B.n575 B.n574 163.367
R919 B.n574 B.n111 163.367
R920 B.n570 B.n111 163.367
R921 B.n570 B.n569 163.367
R922 B.n569 B.n568 163.367
R923 B.n568 B.n113 163.367
R924 B.n564 B.n113 163.367
R925 B.n564 B.n563 163.367
R926 B.n563 B.n562 163.367
R927 B.n562 B.n115 163.367
R928 B.n558 B.n115 163.367
R929 B.n558 B.n557 163.367
R930 B.n557 B.n556 163.367
R931 B.n556 B.n117 163.367
R932 B.n552 B.n117 163.367
R933 B.n552 B.n551 163.367
R934 B.n551 B.n550 163.367
R935 B.n550 B.n119 163.367
R936 B.n546 B.n119 163.367
R937 B.n546 B.n545 163.367
R938 B.n545 B.n544 163.367
R939 B.n544 B.n121 163.367
R940 B.n540 B.n121 163.367
R941 B.n540 B.n539 163.367
R942 B.n539 B.n538 163.367
R943 B.n538 B.n123 163.367
R944 B.n534 B.n123 163.367
R945 B.n534 B.n533 163.367
R946 B.n533 B.n532 163.367
R947 B.n532 B.n125 163.367
R948 B.n528 B.n125 163.367
R949 B.n528 B.n527 163.367
R950 B.n527 B.n526 163.367
R951 B.n526 B.n127 163.367
R952 B.n522 B.n127 163.367
R953 B.n522 B.n521 163.367
R954 B.n521 B.n520 163.367
R955 B.n520 B.n129 163.367
R956 B.n516 B.n129 163.367
R957 B.n516 B.n515 163.367
R958 B.n515 B.n514 163.367
R959 B.n514 B.n131 163.367
R960 B.n510 B.n131 163.367
R961 B.n510 B.n509 163.367
R962 B.n509 B.n508 163.367
R963 B.n508 B.n133 163.367
R964 B.n504 B.n133 163.367
R965 B.n504 B.n503 163.367
R966 B.n503 B.n502 163.367
R967 B.n502 B.n135 163.367
R968 B.n498 B.n135 163.367
R969 B.n498 B.n497 163.367
R970 B.n497 B.n496 163.367
R971 B.n496 B.n137 163.367
R972 B.n492 B.n137 163.367
R973 B.n492 B.n491 163.367
R974 B.n491 B.n490 163.367
R975 B.n490 B.n139 163.367
R976 B.n486 B.n139 163.367
R977 B.n486 B.n485 163.367
R978 B.n485 B.n484 163.367
R979 B.n484 B.n141 163.367
R980 B.n480 B.n141 163.367
R981 B.n480 B.n479 163.367
R982 B.n479 B.n478 163.367
R983 B.n478 B.n143 163.367
R984 B.n474 B.n143 163.367
R985 B.n474 B.n473 163.367
R986 B.n473 B.n472 163.367
R987 B.n472 B.n145 163.367
R988 B.n468 B.n145 163.367
R989 B.n468 B.n467 163.367
R990 B.n467 B.n466 163.367
R991 B.n466 B.n147 163.367
R992 B.n462 B.n147 163.367
R993 B.n462 B.n461 163.367
R994 B.n461 B.n460 163.367
R995 B.n460 B.n149 163.367
R996 B.n456 B.n149 163.367
R997 B.n456 B.n455 163.367
R998 B.n455 B.n454 163.367
R999 B.n454 B.n151 163.367
R1000 B.n450 B.n151 163.367
R1001 B.n780 B.n779 163.367
R1002 B.n779 B.n778 163.367
R1003 B.n778 B.n39 163.367
R1004 B.n774 B.n39 163.367
R1005 B.n774 B.n773 163.367
R1006 B.n773 B.n772 163.367
R1007 B.n772 B.n41 163.367
R1008 B.n768 B.n41 163.367
R1009 B.n768 B.n767 163.367
R1010 B.n767 B.n766 163.367
R1011 B.n766 B.n43 163.367
R1012 B.n762 B.n43 163.367
R1013 B.n762 B.n761 163.367
R1014 B.n761 B.n760 163.367
R1015 B.n760 B.n45 163.367
R1016 B.n756 B.n45 163.367
R1017 B.n756 B.n755 163.367
R1018 B.n755 B.n754 163.367
R1019 B.n754 B.n47 163.367
R1020 B.n750 B.n47 163.367
R1021 B.n750 B.n749 163.367
R1022 B.n749 B.n748 163.367
R1023 B.n748 B.n49 163.367
R1024 B.n744 B.n49 163.367
R1025 B.n744 B.n743 163.367
R1026 B.n743 B.n742 163.367
R1027 B.n742 B.n51 163.367
R1028 B.n738 B.n51 163.367
R1029 B.n738 B.n737 163.367
R1030 B.n737 B.n736 163.367
R1031 B.n736 B.n53 163.367
R1032 B.n732 B.n53 163.367
R1033 B.n732 B.n731 163.367
R1034 B.n731 B.n57 163.367
R1035 B.n727 B.n57 163.367
R1036 B.n727 B.n726 163.367
R1037 B.n726 B.n725 163.367
R1038 B.n725 B.n59 163.367
R1039 B.n721 B.n59 163.367
R1040 B.n721 B.n720 163.367
R1041 B.n720 B.n719 163.367
R1042 B.n719 B.n61 163.367
R1043 B.n714 B.n61 163.367
R1044 B.n714 B.n713 163.367
R1045 B.n713 B.n712 163.367
R1046 B.n712 B.n65 163.367
R1047 B.n708 B.n65 163.367
R1048 B.n708 B.n707 163.367
R1049 B.n707 B.n706 163.367
R1050 B.n706 B.n67 163.367
R1051 B.n702 B.n67 163.367
R1052 B.n702 B.n701 163.367
R1053 B.n701 B.n700 163.367
R1054 B.n700 B.n69 163.367
R1055 B.n696 B.n69 163.367
R1056 B.n696 B.n695 163.367
R1057 B.n695 B.n694 163.367
R1058 B.n694 B.n71 163.367
R1059 B.n690 B.n71 163.367
R1060 B.n690 B.n689 163.367
R1061 B.n689 B.n688 163.367
R1062 B.n688 B.n73 163.367
R1063 B.n684 B.n73 163.367
R1064 B.n684 B.n683 163.367
R1065 B.n683 B.n682 163.367
R1066 B.n682 B.n75 163.367
R1067 B.n678 B.n75 163.367
R1068 B.n678 B.n677 163.367
R1069 B.n677 B.n676 163.367
R1070 B.n676 B.n77 163.367
R1071 B.n672 B.n77 163.367
R1072 B.n672 B.n671 163.367
R1073 B.n671 B.n670 163.367
R1074 B.n670 B.n79 163.367
R1075 B.n666 B.n79 163.367
R1076 B.n784 B.n37 163.367
R1077 B.n785 B.n784 163.367
R1078 B.n786 B.n785 163.367
R1079 B.n786 B.n35 163.367
R1080 B.n790 B.n35 163.367
R1081 B.n791 B.n790 163.367
R1082 B.n792 B.n791 163.367
R1083 B.n792 B.n33 163.367
R1084 B.n796 B.n33 163.367
R1085 B.n797 B.n796 163.367
R1086 B.n798 B.n797 163.367
R1087 B.n798 B.n31 163.367
R1088 B.n802 B.n31 163.367
R1089 B.n803 B.n802 163.367
R1090 B.n804 B.n803 163.367
R1091 B.n804 B.n29 163.367
R1092 B.n808 B.n29 163.367
R1093 B.n809 B.n808 163.367
R1094 B.n810 B.n809 163.367
R1095 B.n810 B.n27 163.367
R1096 B.n814 B.n27 163.367
R1097 B.n815 B.n814 163.367
R1098 B.n816 B.n815 163.367
R1099 B.n816 B.n25 163.367
R1100 B.n820 B.n25 163.367
R1101 B.n821 B.n820 163.367
R1102 B.n822 B.n821 163.367
R1103 B.n822 B.n23 163.367
R1104 B.n826 B.n23 163.367
R1105 B.n827 B.n826 163.367
R1106 B.n828 B.n827 163.367
R1107 B.n828 B.n21 163.367
R1108 B.n832 B.n21 163.367
R1109 B.n833 B.n832 163.367
R1110 B.n834 B.n833 163.367
R1111 B.n834 B.n19 163.367
R1112 B.n838 B.n19 163.367
R1113 B.n839 B.n838 163.367
R1114 B.n840 B.n839 163.367
R1115 B.n840 B.n17 163.367
R1116 B.n844 B.n17 163.367
R1117 B.n845 B.n844 163.367
R1118 B.n846 B.n845 163.367
R1119 B.n846 B.n15 163.367
R1120 B.n850 B.n15 163.367
R1121 B.n851 B.n850 163.367
R1122 B.n852 B.n851 163.367
R1123 B.n852 B.n13 163.367
R1124 B.n856 B.n13 163.367
R1125 B.n857 B.n856 163.367
R1126 B.n858 B.n857 163.367
R1127 B.n858 B.n11 163.367
R1128 B.n862 B.n11 163.367
R1129 B.n863 B.n862 163.367
R1130 B.n864 B.n863 163.367
R1131 B.n864 B.n9 163.367
R1132 B.n868 B.n9 163.367
R1133 B.n869 B.n868 163.367
R1134 B.n870 B.n869 163.367
R1135 B.n870 B.n7 163.367
R1136 B.n874 B.n7 163.367
R1137 B.n875 B.n874 163.367
R1138 B.n876 B.n875 163.367
R1139 B.n876 B.n5 163.367
R1140 B.n880 B.n5 163.367
R1141 B.n881 B.n880 163.367
R1142 B.n882 B.n881 163.367
R1143 B.n882 B.n3 163.367
R1144 B.n886 B.n3 163.367
R1145 B.n887 B.n886 163.367
R1146 B.n228 B.n2 163.367
R1147 B.n229 B.n228 163.367
R1148 B.n230 B.n229 163.367
R1149 B.n230 B.n225 163.367
R1150 B.n234 B.n225 163.367
R1151 B.n235 B.n234 163.367
R1152 B.n236 B.n235 163.367
R1153 B.n236 B.n223 163.367
R1154 B.n240 B.n223 163.367
R1155 B.n241 B.n240 163.367
R1156 B.n242 B.n241 163.367
R1157 B.n242 B.n221 163.367
R1158 B.n246 B.n221 163.367
R1159 B.n247 B.n246 163.367
R1160 B.n248 B.n247 163.367
R1161 B.n248 B.n219 163.367
R1162 B.n252 B.n219 163.367
R1163 B.n253 B.n252 163.367
R1164 B.n254 B.n253 163.367
R1165 B.n254 B.n217 163.367
R1166 B.n258 B.n217 163.367
R1167 B.n259 B.n258 163.367
R1168 B.n260 B.n259 163.367
R1169 B.n260 B.n215 163.367
R1170 B.n264 B.n215 163.367
R1171 B.n265 B.n264 163.367
R1172 B.n266 B.n265 163.367
R1173 B.n266 B.n213 163.367
R1174 B.n270 B.n213 163.367
R1175 B.n271 B.n270 163.367
R1176 B.n272 B.n271 163.367
R1177 B.n272 B.n211 163.367
R1178 B.n276 B.n211 163.367
R1179 B.n277 B.n276 163.367
R1180 B.n278 B.n277 163.367
R1181 B.n278 B.n209 163.367
R1182 B.n282 B.n209 163.367
R1183 B.n283 B.n282 163.367
R1184 B.n284 B.n283 163.367
R1185 B.n284 B.n207 163.367
R1186 B.n288 B.n207 163.367
R1187 B.n289 B.n288 163.367
R1188 B.n290 B.n289 163.367
R1189 B.n290 B.n205 163.367
R1190 B.n294 B.n205 163.367
R1191 B.n295 B.n294 163.367
R1192 B.n296 B.n295 163.367
R1193 B.n296 B.n203 163.367
R1194 B.n300 B.n203 163.367
R1195 B.n301 B.n300 163.367
R1196 B.n302 B.n301 163.367
R1197 B.n302 B.n201 163.367
R1198 B.n306 B.n201 163.367
R1199 B.n307 B.n306 163.367
R1200 B.n308 B.n307 163.367
R1201 B.n308 B.n199 163.367
R1202 B.n312 B.n199 163.367
R1203 B.n313 B.n312 163.367
R1204 B.n314 B.n313 163.367
R1205 B.n314 B.n197 163.367
R1206 B.n318 B.n197 163.367
R1207 B.n319 B.n318 163.367
R1208 B.n320 B.n319 163.367
R1209 B.n320 B.n195 163.367
R1210 B.n324 B.n195 163.367
R1211 B.n325 B.n324 163.367
R1212 B.n326 B.n325 163.367
R1213 B.n326 B.n193 163.367
R1214 B.n330 B.n193 163.367
R1215 B.n331 B.n330 163.367
R1216 B.n397 B.t5 113.287
R1217 B.n63 B.t10 113.287
R1218 B.n175 B.t8 113.276
R1219 B.n55 B.t1 113.276
R1220 B.n175 B.n174 83.7823
R1221 B.n397 B.n396 83.7823
R1222 B.n63 B.n62 83.7823
R1223 B.n55 B.n54 83.7823
R1224 B.n382 B.n175 59.5399
R1225 B.n398 B.n397 59.5399
R1226 B.n716 B.n63 59.5399
R1227 B.n56 B.n55 59.5399
R1228 B.n782 B.n781 32.9371
R1229 B.n667 B.n80 32.9371
R1230 B.n451 B.n152 32.9371
R1231 B.n333 B.n192 32.9371
R1232 B B.n889 18.0485
R1233 B.n783 B.n782 10.6151
R1234 B.n783 B.n36 10.6151
R1235 B.n787 B.n36 10.6151
R1236 B.n788 B.n787 10.6151
R1237 B.n789 B.n788 10.6151
R1238 B.n789 B.n34 10.6151
R1239 B.n793 B.n34 10.6151
R1240 B.n794 B.n793 10.6151
R1241 B.n795 B.n794 10.6151
R1242 B.n795 B.n32 10.6151
R1243 B.n799 B.n32 10.6151
R1244 B.n800 B.n799 10.6151
R1245 B.n801 B.n800 10.6151
R1246 B.n801 B.n30 10.6151
R1247 B.n805 B.n30 10.6151
R1248 B.n806 B.n805 10.6151
R1249 B.n807 B.n806 10.6151
R1250 B.n807 B.n28 10.6151
R1251 B.n811 B.n28 10.6151
R1252 B.n812 B.n811 10.6151
R1253 B.n813 B.n812 10.6151
R1254 B.n813 B.n26 10.6151
R1255 B.n817 B.n26 10.6151
R1256 B.n818 B.n817 10.6151
R1257 B.n819 B.n818 10.6151
R1258 B.n819 B.n24 10.6151
R1259 B.n823 B.n24 10.6151
R1260 B.n824 B.n823 10.6151
R1261 B.n825 B.n824 10.6151
R1262 B.n825 B.n22 10.6151
R1263 B.n829 B.n22 10.6151
R1264 B.n830 B.n829 10.6151
R1265 B.n831 B.n830 10.6151
R1266 B.n831 B.n20 10.6151
R1267 B.n835 B.n20 10.6151
R1268 B.n836 B.n835 10.6151
R1269 B.n837 B.n836 10.6151
R1270 B.n837 B.n18 10.6151
R1271 B.n841 B.n18 10.6151
R1272 B.n842 B.n841 10.6151
R1273 B.n843 B.n842 10.6151
R1274 B.n843 B.n16 10.6151
R1275 B.n847 B.n16 10.6151
R1276 B.n848 B.n847 10.6151
R1277 B.n849 B.n848 10.6151
R1278 B.n849 B.n14 10.6151
R1279 B.n853 B.n14 10.6151
R1280 B.n854 B.n853 10.6151
R1281 B.n855 B.n854 10.6151
R1282 B.n855 B.n12 10.6151
R1283 B.n859 B.n12 10.6151
R1284 B.n860 B.n859 10.6151
R1285 B.n861 B.n860 10.6151
R1286 B.n861 B.n10 10.6151
R1287 B.n865 B.n10 10.6151
R1288 B.n866 B.n865 10.6151
R1289 B.n867 B.n866 10.6151
R1290 B.n867 B.n8 10.6151
R1291 B.n871 B.n8 10.6151
R1292 B.n872 B.n871 10.6151
R1293 B.n873 B.n872 10.6151
R1294 B.n873 B.n6 10.6151
R1295 B.n877 B.n6 10.6151
R1296 B.n878 B.n877 10.6151
R1297 B.n879 B.n878 10.6151
R1298 B.n879 B.n4 10.6151
R1299 B.n883 B.n4 10.6151
R1300 B.n884 B.n883 10.6151
R1301 B.n885 B.n884 10.6151
R1302 B.n885 B.n0 10.6151
R1303 B.n781 B.n38 10.6151
R1304 B.n777 B.n38 10.6151
R1305 B.n777 B.n776 10.6151
R1306 B.n776 B.n775 10.6151
R1307 B.n775 B.n40 10.6151
R1308 B.n771 B.n40 10.6151
R1309 B.n771 B.n770 10.6151
R1310 B.n770 B.n769 10.6151
R1311 B.n769 B.n42 10.6151
R1312 B.n765 B.n42 10.6151
R1313 B.n765 B.n764 10.6151
R1314 B.n764 B.n763 10.6151
R1315 B.n763 B.n44 10.6151
R1316 B.n759 B.n44 10.6151
R1317 B.n759 B.n758 10.6151
R1318 B.n758 B.n757 10.6151
R1319 B.n757 B.n46 10.6151
R1320 B.n753 B.n46 10.6151
R1321 B.n753 B.n752 10.6151
R1322 B.n752 B.n751 10.6151
R1323 B.n751 B.n48 10.6151
R1324 B.n747 B.n48 10.6151
R1325 B.n747 B.n746 10.6151
R1326 B.n746 B.n745 10.6151
R1327 B.n745 B.n50 10.6151
R1328 B.n741 B.n50 10.6151
R1329 B.n741 B.n740 10.6151
R1330 B.n740 B.n739 10.6151
R1331 B.n739 B.n52 10.6151
R1332 B.n735 B.n52 10.6151
R1333 B.n735 B.n734 10.6151
R1334 B.n734 B.n733 10.6151
R1335 B.n730 B.n729 10.6151
R1336 B.n729 B.n728 10.6151
R1337 B.n728 B.n58 10.6151
R1338 B.n724 B.n58 10.6151
R1339 B.n724 B.n723 10.6151
R1340 B.n723 B.n722 10.6151
R1341 B.n722 B.n60 10.6151
R1342 B.n718 B.n60 10.6151
R1343 B.n718 B.n717 10.6151
R1344 B.n715 B.n64 10.6151
R1345 B.n711 B.n64 10.6151
R1346 B.n711 B.n710 10.6151
R1347 B.n710 B.n709 10.6151
R1348 B.n709 B.n66 10.6151
R1349 B.n705 B.n66 10.6151
R1350 B.n705 B.n704 10.6151
R1351 B.n704 B.n703 10.6151
R1352 B.n703 B.n68 10.6151
R1353 B.n699 B.n68 10.6151
R1354 B.n699 B.n698 10.6151
R1355 B.n698 B.n697 10.6151
R1356 B.n697 B.n70 10.6151
R1357 B.n693 B.n70 10.6151
R1358 B.n693 B.n692 10.6151
R1359 B.n692 B.n691 10.6151
R1360 B.n691 B.n72 10.6151
R1361 B.n687 B.n72 10.6151
R1362 B.n687 B.n686 10.6151
R1363 B.n686 B.n685 10.6151
R1364 B.n685 B.n74 10.6151
R1365 B.n681 B.n74 10.6151
R1366 B.n681 B.n680 10.6151
R1367 B.n680 B.n679 10.6151
R1368 B.n679 B.n76 10.6151
R1369 B.n675 B.n76 10.6151
R1370 B.n675 B.n674 10.6151
R1371 B.n674 B.n673 10.6151
R1372 B.n673 B.n78 10.6151
R1373 B.n669 B.n78 10.6151
R1374 B.n669 B.n668 10.6151
R1375 B.n668 B.n667 10.6151
R1376 B.n663 B.n80 10.6151
R1377 B.n663 B.n662 10.6151
R1378 B.n662 B.n661 10.6151
R1379 B.n661 B.n82 10.6151
R1380 B.n657 B.n82 10.6151
R1381 B.n657 B.n656 10.6151
R1382 B.n656 B.n655 10.6151
R1383 B.n655 B.n84 10.6151
R1384 B.n651 B.n84 10.6151
R1385 B.n651 B.n650 10.6151
R1386 B.n650 B.n649 10.6151
R1387 B.n649 B.n86 10.6151
R1388 B.n645 B.n86 10.6151
R1389 B.n645 B.n644 10.6151
R1390 B.n644 B.n643 10.6151
R1391 B.n643 B.n88 10.6151
R1392 B.n639 B.n88 10.6151
R1393 B.n639 B.n638 10.6151
R1394 B.n638 B.n637 10.6151
R1395 B.n637 B.n90 10.6151
R1396 B.n633 B.n90 10.6151
R1397 B.n633 B.n632 10.6151
R1398 B.n632 B.n631 10.6151
R1399 B.n631 B.n92 10.6151
R1400 B.n627 B.n92 10.6151
R1401 B.n627 B.n626 10.6151
R1402 B.n626 B.n625 10.6151
R1403 B.n625 B.n94 10.6151
R1404 B.n621 B.n94 10.6151
R1405 B.n621 B.n620 10.6151
R1406 B.n620 B.n619 10.6151
R1407 B.n619 B.n96 10.6151
R1408 B.n615 B.n96 10.6151
R1409 B.n615 B.n614 10.6151
R1410 B.n614 B.n613 10.6151
R1411 B.n613 B.n98 10.6151
R1412 B.n609 B.n98 10.6151
R1413 B.n609 B.n608 10.6151
R1414 B.n608 B.n607 10.6151
R1415 B.n607 B.n100 10.6151
R1416 B.n603 B.n100 10.6151
R1417 B.n603 B.n602 10.6151
R1418 B.n602 B.n601 10.6151
R1419 B.n601 B.n102 10.6151
R1420 B.n597 B.n102 10.6151
R1421 B.n597 B.n596 10.6151
R1422 B.n596 B.n595 10.6151
R1423 B.n595 B.n104 10.6151
R1424 B.n591 B.n104 10.6151
R1425 B.n591 B.n590 10.6151
R1426 B.n590 B.n589 10.6151
R1427 B.n589 B.n106 10.6151
R1428 B.n585 B.n106 10.6151
R1429 B.n585 B.n584 10.6151
R1430 B.n584 B.n583 10.6151
R1431 B.n583 B.n108 10.6151
R1432 B.n579 B.n108 10.6151
R1433 B.n579 B.n578 10.6151
R1434 B.n578 B.n577 10.6151
R1435 B.n577 B.n110 10.6151
R1436 B.n573 B.n110 10.6151
R1437 B.n573 B.n572 10.6151
R1438 B.n572 B.n571 10.6151
R1439 B.n571 B.n112 10.6151
R1440 B.n567 B.n112 10.6151
R1441 B.n567 B.n566 10.6151
R1442 B.n566 B.n565 10.6151
R1443 B.n565 B.n114 10.6151
R1444 B.n561 B.n114 10.6151
R1445 B.n561 B.n560 10.6151
R1446 B.n560 B.n559 10.6151
R1447 B.n559 B.n116 10.6151
R1448 B.n555 B.n116 10.6151
R1449 B.n555 B.n554 10.6151
R1450 B.n554 B.n553 10.6151
R1451 B.n553 B.n118 10.6151
R1452 B.n549 B.n118 10.6151
R1453 B.n549 B.n548 10.6151
R1454 B.n548 B.n547 10.6151
R1455 B.n547 B.n120 10.6151
R1456 B.n543 B.n120 10.6151
R1457 B.n543 B.n542 10.6151
R1458 B.n542 B.n541 10.6151
R1459 B.n541 B.n122 10.6151
R1460 B.n537 B.n122 10.6151
R1461 B.n537 B.n536 10.6151
R1462 B.n536 B.n535 10.6151
R1463 B.n535 B.n124 10.6151
R1464 B.n531 B.n124 10.6151
R1465 B.n531 B.n530 10.6151
R1466 B.n530 B.n529 10.6151
R1467 B.n529 B.n126 10.6151
R1468 B.n525 B.n126 10.6151
R1469 B.n525 B.n524 10.6151
R1470 B.n524 B.n523 10.6151
R1471 B.n523 B.n128 10.6151
R1472 B.n519 B.n128 10.6151
R1473 B.n519 B.n518 10.6151
R1474 B.n518 B.n517 10.6151
R1475 B.n517 B.n130 10.6151
R1476 B.n513 B.n130 10.6151
R1477 B.n513 B.n512 10.6151
R1478 B.n512 B.n511 10.6151
R1479 B.n511 B.n132 10.6151
R1480 B.n507 B.n132 10.6151
R1481 B.n507 B.n506 10.6151
R1482 B.n506 B.n505 10.6151
R1483 B.n505 B.n134 10.6151
R1484 B.n501 B.n134 10.6151
R1485 B.n501 B.n500 10.6151
R1486 B.n500 B.n499 10.6151
R1487 B.n499 B.n136 10.6151
R1488 B.n495 B.n136 10.6151
R1489 B.n495 B.n494 10.6151
R1490 B.n494 B.n493 10.6151
R1491 B.n493 B.n138 10.6151
R1492 B.n489 B.n138 10.6151
R1493 B.n489 B.n488 10.6151
R1494 B.n488 B.n487 10.6151
R1495 B.n487 B.n140 10.6151
R1496 B.n483 B.n140 10.6151
R1497 B.n483 B.n482 10.6151
R1498 B.n482 B.n481 10.6151
R1499 B.n481 B.n142 10.6151
R1500 B.n477 B.n142 10.6151
R1501 B.n477 B.n476 10.6151
R1502 B.n476 B.n475 10.6151
R1503 B.n475 B.n144 10.6151
R1504 B.n471 B.n144 10.6151
R1505 B.n471 B.n470 10.6151
R1506 B.n470 B.n469 10.6151
R1507 B.n469 B.n146 10.6151
R1508 B.n465 B.n146 10.6151
R1509 B.n465 B.n464 10.6151
R1510 B.n464 B.n463 10.6151
R1511 B.n463 B.n148 10.6151
R1512 B.n459 B.n148 10.6151
R1513 B.n459 B.n458 10.6151
R1514 B.n458 B.n457 10.6151
R1515 B.n457 B.n150 10.6151
R1516 B.n453 B.n150 10.6151
R1517 B.n453 B.n452 10.6151
R1518 B.n452 B.n451 10.6151
R1519 B.n227 B.n1 10.6151
R1520 B.n227 B.n226 10.6151
R1521 B.n231 B.n226 10.6151
R1522 B.n232 B.n231 10.6151
R1523 B.n233 B.n232 10.6151
R1524 B.n233 B.n224 10.6151
R1525 B.n237 B.n224 10.6151
R1526 B.n238 B.n237 10.6151
R1527 B.n239 B.n238 10.6151
R1528 B.n239 B.n222 10.6151
R1529 B.n243 B.n222 10.6151
R1530 B.n244 B.n243 10.6151
R1531 B.n245 B.n244 10.6151
R1532 B.n245 B.n220 10.6151
R1533 B.n249 B.n220 10.6151
R1534 B.n250 B.n249 10.6151
R1535 B.n251 B.n250 10.6151
R1536 B.n251 B.n218 10.6151
R1537 B.n255 B.n218 10.6151
R1538 B.n256 B.n255 10.6151
R1539 B.n257 B.n256 10.6151
R1540 B.n257 B.n216 10.6151
R1541 B.n261 B.n216 10.6151
R1542 B.n262 B.n261 10.6151
R1543 B.n263 B.n262 10.6151
R1544 B.n263 B.n214 10.6151
R1545 B.n267 B.n214 10.6151
R1546 B.n268 B.n267 10.6151
R1547 B.n269 B.n268 10.6151
R1548 B.n269 B.n212 10.6151
R1549 B.n273 B.n212 10.6151
R1550 B.n274 B.n273 10.6151
R1551 B.n275 B.n274 10.6151
R1552 B.n275 B.n210 10.6151
R1553 B.n279 B.n210 10.6151
R1554 B.n280 B.n279 10.6151
R1555 B.n281 B.n280 10.6151
R1556 B.n281 B.n208 10.6151
R1557 B.n285 B.n208 10.6151
R1558 B.n286 B.n285 10.6151
R1559 B.n287 B.n286 10.6151
R1560 B.n287 B.n206 10.6151
R1561 B.n291 B.n206 10.6151
R1562 B.n292 B.n291 10.6151
R1563 B.n293 B.n292 10.6151
R1564 B.n293 B.n204 10.6151
R1565 B.n297 B.n204 10.6151
R1566 B.n298 B.n297 10.6151
R1567 B.n299 B.n298 10.6151
R1568 B.n299 B.n202 10.6151
R1569 B.n303 B.n202 10.6151
R1570 B.n304 B.n303 10.6151
R1571 B.n305 B.n304 10.6151
R1572 B.n305 B.n200 10.6151
R1573 B.n309 B.n200 10.6151
R1574 B.n310 B.n309 10.6151
R1575 B.n311 B.n310 10.6151
R1576 B.n311 B.n198 10.6151
R1577 B.n315 B.n198 10.6151
R1578 B.n316 B.n315 10.6151
R1579 B.n317 B.n316 10.6151
R1580 B.n317 B.n196 10.6151
R1581 B.n321 B.n196 10.6151
R1582 B.n322 B.n321 10.6151
R1583 B.n323 B.n322 10.6151
R1584 B.n323 B.n194 10.6151
R1585 B.n327 B.n194 10.6151
R1586 B.n328 B.n327 10.6151
R1587 B.n329 B.n328 10.6151
R1588 B.n329 B.n192 10.6151
R1589 B.n334 B.n333 10.6151
R1590 B.n335 B.n334 10.6151
R1591 B.n335 B.n190 10.6151
R1592 B.n339 B.n190 10.6151
R1593 B.n340 B.n339 10.6151
R1594 B.n341 B.n340 10.6151
R1595 B.n341 B.n188 10.6151
R1596 B.n345 B.n188 10.6151
R1597 B.n346 B.n345 10.6151
R1598 B.n347 B.n346 10.6151
R1599 B.n347 B.n186 10.6151
R1600 B.n351 B.n186 10.6151
R1601 B.n352 B.n351 10.6151
R1602 B.n353 B.n352 10.6151
R1603 B.n353 B.n184 10.6151
R1604 B.n357 B.n184 10.6151
R1605 B.n358 B.n357 10.6151
R1606 B.n359 B.n358 10.6151
R1607 B.n359 B.n182 10.6151
R1608 B.n363 B.n182 10.6151
R1609 B.n364 B.n363 10.6151
R1610 B.n365 B.n364 10.6151
R1611 B.n365 B.n180 10.6151
R1612 B.n369 B.n180 10.6151
R1613 B.n370 B.n369 10.6151
R1614 B.n371 B.n370 10.6151
R1615 B.n371 B.n178 10.6151
R1616 B.n375 B.n178 10.6151
R1617 B.n376 B.n375 10.6151
R1618 B.n377 B.n376 10.6151
R1619 B.n377 B.n176 10.6151
R1620 B.n381 B.n176 10.6151
R1621 B.n384 B.n383 10.6151
R1622 B.n384 B.n172 10.6151
R1623 B.n388 B.n172 10.6151
R1624 B.n389 B.n388 10.6151
R1625 B.n390 B.n389 10.6151
R1626 B.n390 B.n170 10.6151
R1627 B.n394 B.n170 10.6151
R1628 B.n395 B.n394 10.6151
R1629 B.n399 B.n395 10.6151
R1630 B.n403 B.n168 10.6151
R1631 B.n404 B.n403 10.6151
R1632 B.n405 B.n404 10.6151
R1633 B.n405 B.n166 10.6151
R1634 B.n409 B.n166 10.6151
R1635 B.n410 B.n409 10.6151
R1636 B.n411 B.n410 10.6151
R1637 B.n411 B.n164 10.6151
R1638 B.n415 B.n164 10.6151
R1639 B.n416 B.n415 10.6151
R1640 B.n417 B.n416 10.6151
R1641 B.n417 B.n162 10.6151
R1642 B.n421 B.n162 10.6151
R1643 B.n422 B.n421 10.6151
R1644 B.n423 B.n422 10.6151
R1645 B.n423 B.n160 10.6151
R1646 B.n427 B.n160 10.6151
R1647 B.n428 B.n427 10.6151
R1648 B.n429 B.n428 10.6151
R1649 B.n429 B.n158 10.6151
R1650 B.n433 B.n158 10.6151
R1651 B.n434 B.n433 10.6151
R1652 B.n435 B.n434 10.6151
R1653 B.n435 B.n156 10.6151
R1654 B.n439 B.n156 10.6151
R1655 B.n440 B.n439 10.6151
R1656 B.n441 B.n440 10.6151
R1657 B.n441 B.n154 10.6151
R1658 B.n445 B.n154 10.6151
R1659 B.n446 B.n445 10.6151
R1660 B.n447 B.n446 10.6151
R1661 B.n447 B.n152 10.6151
R1662 B.n733 B.n56 9.36635
R1663 B.n716 B.n715 9.36635
R1664 B.n382 B.n381 9.36635
R1665 B.n398 B.n168 9.36635
R1666 B.n889 B.n0 8.11757
R1667 B.n889 B.n1 8.11757
R1668 B.n730 B.n56 1.24928
R1669 B.n717 B.n716 1.24928
R1670 B.n383 B.n382 1.24928
R1671 B.n399 B.n398 1.24928
C0 B VN 1.51479f
C1 w_n5290_n2790# B 11.432599f
C2 w_n5290_n2790# VN 11.0985f
C3 VDD2 B 2.13613f
C4 VTAIL VP 8.209929f
C5 VDD2 VN 7.184811f
C6 w_n5290_n2790# VDD2 2.49825f
C7 VDD1 VTAIL 7.9426f
C8 VDD1 VP 7.69605f
C9 VTAIL B 4.53317f
C10 VTAIL VN 8.195829f
C11 w_n5290_n2790# VTAIL 3.7012f
C12 VDD2 VTAIL 8.00634f
C13 B VP 2.6803f
C14 VN VP 8.828059f
C15 w_n5290_n2790# VP 11.7894f
C16 VDD1 B 1.99637f
C17 VDD2 VP 0.667736f
C18 VDD1 VN 0.154396f
C19 VDD1 w_n5290_n2790# 2.32523f
C20 VDD1 VDD2 2.5005f
C21 VDD2 VSUBS 2.56144f
C22 VDD1 VSUBS 3.29891f
C23 VTAIL VSUBS 1.490417f
C24 VN VSUBS 8.620719f
C25 VP VSUBS 4.933962f
C26 B VSUBS 6.308521f
C27 w_n5290_n2790# VSUBS 0.182632p
C28 B.n0 VSUBS 0.007649f
C29 B.n1 VSUBS 0.007649f
C30 B.n2 VSUBS 0.011313f
C31 B.n3 VSUBS 0.008669f
C32 B.n4 VSUBS 0.008669f
C33 B.n5 VSUBS 0.008669f
C34 B.n6 VSUBS 0.008669f
C35 B.n7 VSUBS 0.008669f
C36 B.n8 VSUBS 0.008669f
C37 B.n9 VSUBS 0.008669f
C38 B.n10 VSUBS 0.008669f
C39 B.n11 VSUBS 0.008669f
C40 B.n12 VSUBS 0.008669f
C41 B.n13 VSUBS 0.008669f
C42 B.n14 VSUBS 0.008669f
C43 B.n15 VSUBS 0.008669f
C44 B.n16 VSUBS 0.008669f
C45 B.n17 VSUBS 0.008669f
C46 B.n18 VSUBS 0.008669f
C47 B.n19 VSUBS 0.008669f
C48 B.n20 VSUBS 0.008669f
C49 B.n21 VSUBS 0.008669f
C50 B.n22 VSUBS 0.008669f
C51 B.n23 VSUBS 0.008669f
C52 B.n24 VSUBS 0.008669f
C53 B.n25 VSUBS 0.008669f
C54 B.n26 VSUBS 0.008669f
C55 B.n27 VSUBS 0.008669f
C56 B.n28 VSUBS 0.008669f
C57 B.n29 VSUBS 0.008669f
C58 B.n30 VSUBS 0.008669f
C59 B.n31 VSUBS 0.008669f
C60 B.n32 VSUBS 0.008669f
C61 B.n33 VSUBS 0.008669f
C62 B.n34 VSUBS 0.008669f
C63 B.n35 VSUBS 0.008669f
C64 B.n36 VSUBS 0.008669f
C65 B.n37 VSUBS 0.019717f
C66 B.n38 VSUBS 0.008669f
C67 B.n39 VSUBS 0.008669f
C68 B.n40 VSUBS 0.008669f
C69 B.n41 VSUBS 0.008669f
C70 B.n42 VSUBS 0.008669f
C71 B.n43 VSUBS 0.008669f
C72 B.n44 VSUBS 0.008669f
C73 B.n45 VSUBS 0.008669f
C74 B.n46 VSUBS 0.008669f
C75 B.n47 VSUBS 0.008669f
C76 B.n48 VSUBS 0.008669f
C77 B.n49 VSUBS 0.008669f
C78 B.n50 VSUBS 0.008669f
C79 B.n51 VSUBS 0.008669f
C80 B.n52 VSUBS 0.008669f
C81 B.n53 VSUBS 0.008669f
C82 B.t1 VSUBS 0.355194f
C83 B.t2 VSUBS 0.390655f
C84 B.t0 VSUBS 2.13299f
C85 B.n54 VSUBS 0.22659f
C86 B.n55 VSUBS 0.095769f
C87 B.n56 VSUBS 0.020086f
C88 B.n57 VSUBS 0.008669f
C89 B.n58 VSUBS 0.008669f
C90 B.n59 VSUBS 0.008669f
C91 B.n60 VSUBS 0.008669f
C92 B.n61 VSUBS 0.008669f
C93 B.t10 VSUBS 0.35519f
C94 B.t11 VSUBS 0.39065f
C95 B.t9 VSUBS 2.13299f
C96 B.n62 VSUBS 0.226594f
C97 B.n63 VSUBS 0.095773f
C98 B.n64 VSUBS 0.008669f
C99 B.n65 VSUBS 0.008669f
C100 B.n66 VSUBS 0.008669f
C101 B.n67 VSUBS 0.008669f
C102 B.n68 VSUBS 0.008669f
C103 B.n69 VSUBS 0.008669f
C104 B.n70 VSUBS 0.008669f
C105 B.n71 VSUBS 0.008669f
C106 B.n72 VSUBS 0.008669f
C107 B.n73 VSUBS 0.008669f
C108 B.n74 VSUBS 0.008669f
C109 B.n75 VSUBS 0.008669f
C110 B.n76 VSUBS 0.008669f
C111 B.n77 VSUBS 0.008669f
C112 B.n78 VSUBS 0.008669f
C113 B.n79 VSUBS 0.008669f
C114 B.n80 VSUBS 0.019717f
C115 B.n81 VSUBS 0.008669f
C116 B.n82 VSUBS 0.008669f
C117 B.n83 VSUBS 0.008669f
C118 B.n84 VSUBS 0.008669f
C119 B.n85 VSUBS 0.008669f
C120 B.n86 VSUBS 0.008669f
C121 B.n87 VSUBS 0.008669f
C122 B.n88 VSUBS 0.008669f
C123 B.n89 VSUBS 0.008669f
C124 B.n90 VSUBS 0.008669f
C125 B.n91 VSUBS 0.008669f
C126 B.n92 VSUBS 0.008669f
C127 B.n93 VSUBS 0.008669f
C128 B.n94 VSUBS 0.008669f
C129 B.n95 VSUBS 0.008669f
C130 B.n96 VSUBS 0.008669f
C131 B.n97 VSUBS 0.008669f
C132 B.n98 VSUBS 0.008669f
C133 B.n99 VSUBS 0.008669f
C134 B.n100 VSUBS 0.008669f
C135 B.n101 VSUBS 0.008669f
C136 B.n102 VSUBS 0.008669f
C137 B.n103 VSUBS 0.008669f
C138 B.n104 VSUBS 0.008669f
C139 B.n105 VSUBS 0.008669f
C140 B.n106 VSUBS 0.008669f
C141 B.n107 VSUBS 0.008669f
C142 B.n108 VSUBS 0.008669f
C143 B.n109 VSUBS 0.008669f
C144 B.n110 VSUBS 0.008669f
C145 B.n111 VSUBS 0.008669f
C146 B.n112 VSUBS 0.008669f
C147 B.n113 VSUBS 0.008669f
C148 B.n114 VSUBS 0.008669f
C149 B.n115 VSUBS 0.008669f
C150 B.n116 VSUBS 0.008669f
C151 B.n117 VSUBS 0.008669f
C152 B.n118 VSUBS 0.008669f
C153 B.n119 VSUBS 0.008669f
C154 B.n120 VSUBS 0.008669f
C155 B.n121 VSUBS 0.008669f
C156 B.n122 VSUBS 0.008669f
C157 B.n123 VSUBS 0.008669f
C158 B.n124 VSUBS 0.008669f
C159 B.n125 VSUBS 0.008669f
C160 B.n126 VSUBS 0.008669f
C161 B.n127 VSUBS 0.008669f
C162 B.n128 VSUBS 0.008669f
C163 B.n129 VSUBS 0.008669f
C164 B.n130 VSUBS 0.008669f
C165 B.n131 VSUBS 0.008669f
C166 B.n132 VSUBS 0.008669f
C167 B.n133 VSUBS 0.008669f
C168 B.n134 VSUBS 0.008669f
C169 B.n135 VSUBS 0.008669f
C170 B.n136 VSUBS 0.008669f
C171 B.n137 VSUBS 0.008669f
C172 B.n138 VSUBS 0.008669f
C173 B.n139 VSUBS 0.008669f
C174 B.n140 VSUBS 0.008669f
C175 B.n141 VSUBS 0.008669f
C176 B.n142 VSUBS 0.008669f
C177 B.n143 VSUBS 0.008669f
C178 B.n144 VSUBS 0.008669f
C179 B.n145 VSUBS 0.008669f
C180 B.n146 VSUBS 0.008669f
C181 B.n147 VSUBS 0.008669f
C182 B.n148 VSUBS 0.008669f
C183 B.n149 VSUBS 0.008669f
C184 B.n150 VSUBS 0.008669f
C185 B.n151 VSUBS 0.008669f
C186 B.n152 VSUBS 0.020064f
C187 B.n153 VSUBS 0.008669f
C188 B.n154 VSUBS 0.008669f
C189 B.n155 VSUBS 0.008669f
C190 B.n156 VSUBS 0.008669f
C191 B.n157 VSUBS 0.008669f
C192 B.n158 VSUBS 0.008669f
C193 B.n159 VSUBS 0.008669f
C194 B.n160 VSUBS 0.008669f
C195 B.n161 VSUBS 0.008669f
C196 B.n162 VSUBS 0.008669f
C197 B.n163 VSUBS 0.008669f
C198 B.n164 VSUBS 0.008669f
C199 B.n165 VSUBS 0.008669f
C200 B.n166 VSUBS 0.008669f
C201 B.n167 VSUBS 0.008669f
C202 B.n168 VSUBS 0.008159f
C203 B.n169 VSUBS 0.008669f
C204 B.n170 VSUBS 0.008669f
C205 B.n171 VSUBS 0.008669f
C206 B.n172 VSUBS 0.008669f
C207 B.n173 VSUBS 0.008669f
C208 B.t8 VSUBS 0.355194f
C209 B.t7 VSUBS 0.390655f
C210 B.t6 VSUBS 2.13299f
C211 B.n174 VSUBS 0.22659f
C212 B.n175 VSUBS 0.095769f
C213 B.n176 VSUBS 0.008669f
C214 B.n177 VSUBS 0.008669f
C215 B.n178 VSUBS 0.008669f
C216 B.n179 VSUBS 0.008669f
C217 B.n180 VSUBS 0.008669f
C218 B.n181 VSUBS 0.008669f
C219 B.n182 VSUBS 0.008669f
C220 B.n183 VSUBS 0.008669f
C221 B.n184 VSUBS 0.008669f
C222 B.n185 VSUBS 0.008669f
C223 B.n186 VSUBS 0.008669f
C224 B.n187 VSUBS 0.008669f
C225 B.n188 VSUBS 0.008669f
C226 B.n189 VSUBS 0.008669f
C227 B.n190 VSUBS 0.008669f
C228 B.n191 VSUBS 0.008669f
C229 B.n192 VSUBS 0.019717f
C230 B.n193 VSUBS 0.008669f
C231 B.n194 VSUBS 0.008669f
C232 B.n195 VSUBS 0.008669f
C233 B.n196 VSUBS 0.008669f
C234 B.n197 VSUBS 0.008669f
C235 B.n198 VSUBS 0.008669f
C236 B.n199 VSUBS 0.008669f
C237 B.n200 VSUBS 0.008669f
C238 B.n201 VSUBS 0.008669f
C239 B.n202 VSUBS 0.008669f
C240 B.n203 VSUBS 0.008669f
C241 B.n204 VSUBS 0.008669f
C242 B.n205 VSUBS 0.008669f
C243 B.n206 VSUBS 0.008669f
C244 B.n207 VSUBS 0.008669f
C245 B.n208 VSUBS 0.008669f
C246 B.n209 VSUBS 0.008669f
C247 B.n210 VSUBS 0.008669f
C248 B.n211 VSUBS 0.008669f
C249 B.n212 VSUBS 0.008669f
C250 B.n213 VSUBS 0.008669f
C251 B.n214 VSUBS 0.008669f
C252 B.n215 VSUBS 0.008669f
C253 B.n216 VSUBS 0.008669f
C254 B.n217 VSUBS 0.008669f
C255 B.n218 VSUBS 0.008669f
C256 B.n219 VSUBS 0.008669f
C257 B.n220 VSUBS 0.008669f
C258 B.n221 VSUBS 0.008669f
C259 B.n222 VSUBS 0.008669f
C260 B.n223 VSUBS 0.008669f
C261 B.n224 VSUBS 0.008669f
C262 B.n225 VSUBS 0.008669f
C263 B.n226 VSUBS 0.008669f
C264 B.n227 VSUBS 0.008669f
C265 B.n228 VSUBS 0.008669f
C266 B.n229 VSUBS 0.008669f
C267 B.n230 VSUBS 0.008669f
C268 B.n231 VSUBS 0.008669f
C269 B.n232 VSUBS 0.008669f
C270 B.n233 VSUBS 0.008669f
C271 B.n234 VSUBS 0.008669f
C272 B.n235 VSUBS 0.008669f
C273 B.n236 VSUBS 0.008669f
C274 B.n237 VSUBS 0.008669f
C275 B.n238 VSUBS 0.008669f
C276 B.n239 VSUBS 0.008669f
C277 B.n240 VSUBS 0.008669f
C278 B.n241 VSUBS 0.008669f
C279 B.n242 VSUBS 0.008669f
C280 B.n243 VSUBS 0.008669f
C281 B.n244 VSUBS 0.008669f
C282 B.n245 VSUBS 0.008669f
C283 B.n246 VSUBS 0.008669f
C284 B.n247 VSUBS 0.008669f
C285 B.n248 VSUBS 0.008669f
C286 B.n249 VSUBS 0.008669f
C287 B.n250 VSUBS 0.008669f
C288 B.n251 VSUBS 0.008669f
C289 B.n252 VSUBS 0.008669f
C290 B.n253 VSUBS 0.008669f
C291 B.n254 VSUBS 0.008669f
C292 B.n255 VSUBS 0.008669f
C293 B.n256 VSUBS 0.008669f
C294 B.n257 VSUBS 0.008669f
C295 B.n258 VSUBS 0.008669f
C296 B.n259 VSUBS 0.008669f
C297 B.n260 VSUBS 0.008669f
C298 B.n261 VSUBS 0.008669f
C299 B.n262 VSUBS 0.008669f
C300 B.n263 VSUBS 0.008669f
C301 B.n264 VSUBS 0.008669f
C302 B.n265 VSUBS 0.008669f
C303 B.n266 VSUBS 0.008669f
C304 B.n267 VSUBS 0.008669f
C305 B.n268 VSUBS 0.008669f
C306 B.n269 VSUBS 0.008669f
C307 B.n270 VSUBS 0.008669f
C308 B.n271 VSUBS 0.008669f
C309 B.n272 VSUBS 0.008669f
C310 B.n273 VSUBS 0.008669f
C311 B.n274 VSUBS 0.008669f
C312 B.n275 VSUBS 0.008669f
C313 B.n276 VSUBS 0.008669f
C314 B.n277 VSUBS 0.008669f
C315 B.n278 VSUBS 0.008669f
C316 B.n279 VSUBS 0.008669f
C317 B.n280 VSUBS 0.008669f
C318 B.n281 VSUBS 0.008669f
C319 B.n282 VSUBS 0.008669f
C320 B.n283 VSUBS 0.008669f
C321 B.n284 VSUBS 0.008669f
C322 B.n285 VSUBS 0.008669f
C323 B.n286 VSUBS 0.008669f
C324 B.n287 VSUBS 0.008669f
C325 B.n288 VSUBS 0.008669f
C326 B.n289 VSUBS 0.008669f
C327 B.n290 VSUBS 0.008669f
C328 B.n291 VSUBS 0.008669f
C329 B.n292 VSUBS 0.008669f
C330 B.n293 VSUBS 0.008669f
C331 B.n294 VSUBS 0.008669f
C332 B.n295 VSUBS 0.008669f
C333 B.n296 VSUBS 0.008669f
C334 B.n297 VSUBS 0.008669f
C335 B.n298 VSUBS 0.008669f
C336 B.n299 VSUBS 0.008669f
C337 B.n300 VSUBS 0.008669f
C338 B.n301 VSUBS 0.008669f
C339 B.n302 VSUBS 0.008669f
C340 B.n303 VSUBS 0.008669f
C341 B.n304 VSUBS 0.008669f
C342 B.n305 VSUBS 0.008669f
C343 B.n306 VSUBS 0.008669f
C344 B.n307 VSUBS 0.008669f
C345 B.n308 VSUBS 0.008669f
C346 B.n309 VSUBS 0.008669f
C347 B.n310 VSUBS 0.008669f
C348 B.n311 VSUBS 0.008669f
C349 B.n312 VSUBS 0.008669f
C350 B.n313 VSUBS 0.008669f
C351 B.n314 VSUBS 0.008669f
C352 B.n315 VSUBS 0.008669f
C353 B.n316 VSUBS 0.008669f
C354 B.n317 VSUBS 0.008669f
C355 B.n318 VSUBS 0.008669f
C356 B.n319 VSUBS 0.008669f
C357 B.n320 VSUBS 0.008669f
C358 B.n321 VSUBS 0.008669f
C359 B.n322 VSUBS 0.008669f
C360 B.n323 VSUBS 0.008669f
C361 B.n324 VSUBS 0.008669f
C362 B.n325 VSUBS 0.008669f
C363 B.n326 VSUBS 0.008669f
C364 B.n327 VSUBS 0.008669f
C365 B.n328 VSUBS 0.008669f
C366 B.n329 VSUBS 0.008669f
C367 B.n330 VSUBS 0.008669f
C368 B.n331 VSUBS 0.019717f
C369 B.n332 VSUBS 0.02108f
C370 B.n333 VSUBS 0.02108f
C371 B.n334 VSUBS 0.008669f
C372 B.n335 VSUBS 0.008669f
C373 B.n336 VSUBS 0.008669f
C374 B.n337 VSUBS 0.008669f
C375 B.n338 VSUBS 0.008669f
C376 B.n339 VSUBS 0.008669f
C377 B.n340 VSUBS 0.008669f
C378 B.n341 VSUBS 0.008669f
C379 B.n342 VSUBS 0.008669f
C380 B.n343 VSUBS 0.008669f
C381 B.n344 VSUBS 0.008669f
C382 B.n345 VSUBS 0.008669f
C383 B.n346 VSUBS 0.008669f
C384 B.n347 VSUBS 0.008669f
C385 B.n348 VSUBS 0.008669f
C386 B.n349 VSUBS 0.008669f
C387 B.n350 VSUBS 0.008669f
C388 B.n351 VSUBS 0.008669f
C389 B.n352 VSUBS 0.008669f
C390 B.n353 VSUBS 0.008669f
C391 B.n354 VSUBS 0.008669f
C392 B.n355 VSUBS 0.008669f
C393 B.n356 VSUBS 0.008669f
C394 B.n357 VSUBS 0.008669f
C395 B.n358 VSUBS 0.008669f
C396 B.n359 VSUBS 0.008669f
C397 B.n360 VSUBS 0.008669f
C398 B.n361 VSUBS 0.008669f
C399 B.n362 VSUBS 0.008669f
C400 B.n363 VSUBS 0.008669f
C401 B.n364 VSUBS 0.008669f
C402 B.n365 VSUBS 0.008669f
C403 B.n366 VSUBS 0.008669f
C404 B.n367 VSUBS 0.008669f
C405 B.n368 VSUBS 0.008669f
C406 B.n369 VSUBS 0.008669f
C407 B.n370 VSUBS 0.008669f
C408 B.n371 VSUBS 0.008669f
C409 B.n372 VSUBS 0.008669f
C410 B.n373 VSUBS 0.008669f
C411 B.n374 VSUBS 0.008669f
C412 B.n375 VSUBS 0.008669f
C413 B.n376 VSUBS 0.008669f
C414 B.n377 VSUBS 0.008669f
C415 B.n378 VSUBS 0.008669f
C416 B.n379 VSUBS 0.008669f
C417 B.n380 VSUBS 0.008669f
C418 B.n381 VSUBS 0.008159f
C419 B.n382 VSUBS 0.020086f
C420 B.n383 VSUBS 0.004845f
C421 B.n384 VSUBS 0.008669f
C422 B.n385 VSUBS 0.008669f
C423 B.n386 VSUBS 0.008669f
C424 B.n387 VSUBS 0.008669f
C425 B.n388 VSUBS 0.008669f
C426 B.n389 VSUBS 0.008669f
C427 B.n390 VSUBS 0.008669f
C428 B.n391 VSUBS 0.008669f
C429 B.n392 VSUBS 0.008669f
C430 B.n393 VSUBS 0.008669f
C431 B.n394 VSUBS 0.008669f
C432 B.n395 VSUBS 0.008669f
C433 B.t5 VSUBS 0.35519f
C434 B.t4 VSUBS 0.39065f
C435 B.t3 VSUBS 2.13299f
C436 B.n396 VSUBS 0.226594f
C437 B.n397 VSUBS 0.095773f
C438 B.n398 VSUBS 0.020086f
C439 B.n399 VSUBS 0.004845f
C440 B.n400 VSUBS 0.008669f
C441 B.n401 VSUBS 0.008669f
C442 B.n402 VSUBS 0.008669f
C443 B.n403 VSUBS 0.008669f
C444 B.n404 VSUBS 0.008669f
C445 B.n405 VSUBS 0.008669f
C446 B.n406 VSUBS 0.008669f
C447 B.n407 VSUBS 0.008669f
C448 B.n408 VSUBS 0.008669f
C449 B.n409 VSUBS 0.008669f
C450 B.n410 VSUBS 0.008669f
C451 B.n411 VSUBS 0.008669f
C452 B.n412 VSUBS 0.008669f
C453 B.n413 VSUBS 0.008669f
C454 B.n414 VSUBS 0.008669f
C455 B.n415 VSUBS 0.008669f
C456 B.n416 VSUBS 0.008669f
C457 B.n417 VSUBS 0.008669f
C458 B.n418 VSUBS 0.008669f
C459 B.n419 VSUBS 0.008669f
C460 B.n420 VSUBS 0.008669f
C461 B.n421 VSUBS 0.008669f
C462 B.n422 VSUBS 0.008669f
C463 B.n423 VSUBS 0.008669f
C464 B.n424 VSUBS 0.008669f
C465 B.n425 VSUBS 0.008669f
C466 B.n426 VSUBS 0.008669f
C467 B.n427 VSUBS 0.008669f
C468 B.n428 VSUBS 0.008669f
C469 B.n429 VSUBS 0.008669f
C470 B.n430 VSUBS 0.008669f
C471 B.n431 VSUBS 0.008669f
C472 B.n432 VSUBS 0.008669f
C473 B.n433 VSUBS 0.008669f
C474 B.n434 VSUBS 0.008669f
C475 B.n435 VSUBS 0.008669f
C476 B.n436 VSUBS 0.008669f
C477 B.n437 VSUBS 0.008669f
C478 B.n438 VSUBS 0.008669f
C479 B.n439 VSUBS 0.008669f
C480 B.n440 VSUBS 0.008669f
C481 B.n441 VSUBS 0.008669f
C482 B.n442 VSUBS 0.008669f
C483 B.n443 VSUBS 0.008669f
C484 B.n444 VSUBS 0.008669f
C485 B.n445 VSUBS 0.008669f
C486 B.n446 VSUBS 0.008669f
C487 B.n447 VSUBS 0.008669f
C488 B.n448 VSUBS 0.008669f
C489 B.n449 VSUBS 0.02108f
C490 B.n450 VSUBS 0.019717f
C491 B.n451 VSUBS 0.020733f
C492 B.n452 VSUBS 0.008669f
C493 B.n453 VSUBS 0.008669f
C494 B.n454 VSUBS 0.008669f
C495 B.n455 VSUBS 0.008669f
C496 B.n456 VSUBS 0.008669f
C497 B.n457 VSUBS 0.008669f
C498 B.n458 VSUBS 0.008669f
C499 B.n459 VSUBS 0.008669f
C500 B.n460 VSUBS 0.008669f
C501 B.n461 VSUBS 0.008669f
C502 B.n462 VSUBS 0.008669f
C503 B.n463 VSUBS 0.008669f
C504 B.n464 VSUBS 0.008669f
C505 B.n465 VSUBS 0.008669f
C506 B.n466 VSUBS 0.008669f
C507 B.n467 VSUBS 0.008669f
C508 B.n468 VSUBS 0.008669f
C509 B.n469 VSUBS 0.008669f
C510 B.n470 VSUBS 0.008669f
C511 B.n471 VSUBS 0.008669f
C512 B.n472 VSUBS 0.008669f
C513 B.n473 VSUBS 0.008669f
C514 B.n474 VSUBS 0.008669f
C515 B.n475 VSUBS 0.008669f
C516 B.n476 VSUBS 0.008669f
C517 B.n477 VSUBS 0.008669f
C518 B.n478 VSUBS 0.008669f
C519 B.n479 VSUBS 0.008669f
C520 B.n480 VSUBS 0.008669f
C521 B.n481 VSUBS 0.008669f
C522 B.n482 VSUBS 0.008669f
C523 B.n483 VSUBS 0.008669f
C524 B.n484 VSUBS 0.008669f
C525 B.n485 VSUBS 0.008669f
C526 B.n486 VSUBS 0.008669f
C527 B.n487 VSUBS 0.008669f
C528 B.n488 VSUBS 0.008669f
C529 B.n489 VSUBS 0.008669f
C530 B.n490 VSUBS 0.008669f
C531 B.n491 VSUBS 0.008669f
C532 B.n492 VSUBS 0.008669f
C533 B.n493 VSUBS 0.008669f
C534 B.n494 VSUBS 0.008669f
C535 B.n495 VSUBS 0.008669f
C536 B.n496 VSUBS 0.008669f
C537 B.n497 VSUBS 0.008669f
C538 B.n498 VSUBS 0.008669f
C539 B.n499 VSUBS 0.008669f
C540 B.n500 VSUBS 0.008669f
C541 B.n501 VSUBS 0.008669f
C542 B.n502 VSUBS 0.008669f
C543 B.n503 VSUBS 0.008669f
C544 B.n504 VSUBS 0.008669f
C545 B.n505 VSUBS 0.008669f
C546 B.n506 VSUBS 0.008669f
C547 B.n507 VSUBS 0.008669f
C548 B.n508 VSUBS 0.008669f
C549 B.n509 VSUBS 0.008669f
C550 B.n510 VSUBS 0.008669f
C551 B.n511 VSUBS 0.008669f
C552 B.n512 VSUBS 0.008669f
C553 B.n513 VSUBS 0.008669f
C554 B.n514 VSUBS 0.008669f
C555 B.n515 VSUBS 0.008669f
C556 B.n516 VSUBS 0.008669f
C557 B.n517 VSUBS 0.008669f
C558 B.n518 VSUBS 0.008669f
C559 B.n519 VSUBS 0.008669f
C560 B.n520 VSUBS 0.008669f
C561 B.n521 VSUBS 0.008669f
C562 B.n522 VSUBS 0.008669f
C563 B.n523 VSUBS 0.008669f
C564 B.n524 VSUBS 0.008669f
C565 B.n525 VSUBS 0.008669f
C566 B.n526 VSUBS 0.008669f
C567 B.n527 VSUBS 0.008669f
C568 B.n528 VSUBS 0.008669f
C569 B.n529 VSUBS 0.008669f
C570 B.n530 VSUBS 0.008669f
C571 B.n531 VSUBS 0.008669f
C572 B.n532 VSUBS 0.008669f
C573 B.n533 VSUBS 0.008669f
C574 B.n534 VSUBS 0.008669f
C575 B.n535 VSUBS 0.008669f
C576 B.n536 VSUBS 0.008669f
C577 B.n537 VSUBS 0.008669f
C578 B.n538 VSUBS 0.008669f
C579 B.n539 VSUBS 0.008669f
C580 B.n540 VSUBS 0.008669f
C581 B.n541 VSUBS 0.008669f
C582 B.n542 VSUBS 0.008669f
C583 B.n543 VSUBS 0.008669f
C584 B.n544 VSUBS 0.008669f
C585 B.n545 VSUBS 0.008669f
C586 B.n546 VSUBS 0.008669f
C587 B.n547 VSUBS 0.008669f
C588 B.n548 VSUBS 0.008669f
C589 B.n549 VSUBS 0.008669f
C590 B.n550 VSUBS 0.008669f
C591 B.n551 VSUBS 0.008669f
C592 B.n552 VSUBS 0.008669f
C593 B.n553 VSUBS 0.008669f
C594 B.n554 VSUBS 0.008669f
C595 B.n555 VSUBS 0.008669f
C596 B.n556 VSUBS 0.008669f
C597 B.n557 VSUBS 0.008669f
C598 B.n558 VSUBS 0.008669f
C599 B.n559 VSUBS 0.008669f
C600 B.n560 VSUBS 0.008669f
C601 B.n561 VSUBS 0.008669f
C602 B.n562 VSUBS 0.008669f
C603 B.n563 VSUBS 0.008669f
C604 B.n564 VSUBS 0.008669f
C605 B.n565 VSUBS 0.008669f
C606 B.n566 VSUBS 0.008669f
C607 B.n567 VSUBS 0.008669f
C608 B.n568 VSUBS 0.008669f
C609 B.n569 VSUBS 0.008669f
C610 B.n570 VSUBS 0.008669f
C611 B.n571 VSUBS 0.008669f
C612 B.n572 VSUBS 0.008669f
C613 B.n573 VSUBS 0.008669f
C614 B.n574 VSUBS 0.008669f
C615 B.n575 VSUBS 0.008669f
C616 B.n576 VSUBS 0.008669f
C617 B.n577 VSUBS 0.008669f
C618 B.n578 VSUBS 0.008669f
C619 B.n579 VSUBS 0.008669f
C620 B.n580 VSUBS 0.008669f
C621 B.n581 VSUBS 0.008669f
C622 B.n582 VSUBS 0.008669f
C623 B.n583 VSUBS 0.008669f
C624 B.n584 VSUBS 0.008669f
C625 B.n585 VSUBS 0.008669f
C626 B.n586 VSUBS 0.008669f
C627 B.n587 VSUBS 0.008669f
C628 B.n588 VSUBS 0.008669f
C629 B.n589 VSUBS 0.008669f
C630 B.n590 VSUBS 0.008669f
C631 B.n591 VSUBS 0.008669f
C632 B.n592 VSUBS 0.008669f
C633 B.n593 VSUBS 0.008669f
C634 B.n594 VSUBS 0.008669f
C635 B.n595 VSUBS 0.008669f
C636 B.n596 VSUBS 0.008669f
C637 B.n597 VSUBS 0.008669f
C638 B.n598 VSUBS 0.008669f
C639 B.n599 VSUBS 0.008669f
C640 B.n600 VSUBS 0.008669f
C641 B.n601 VSUBS 0.008669f
C642 B.n602 VSUBS 0.008669f
C643 B.n603 VSUBS 0.008669f
C644 B.n604 VSUBS 0.008669f
C645 B.n605 VSUBS 0.008669f
C646 B.n606 VSUBS 0.008669f
C647 B.n607 VSUBS 0.008669f
C648 B.n608 VSUBS 0.008669f
C649 B.n609 VSUBS 0.008669f
C650 B.n610 VSUBS 0.008669f
C651 B.n611 VSUBS 0.008669f
C652 B.n612 VSUBS 0.008669f
C653 B.n613 VSUBS 0.008669f
C654 B.n614 VSUBS 0.008669f
C655 B.n615 VSUBS 0.008669f
C656 B.n616 VSUBS 0.008669f
C657 B.n617 VSUBS 0.008669f
C658 B.n618 VSUBS 0.008669f
C659 B.n619 VSUBS 0.008669f
C660 B.n620 VSUBS 0.008669f
C661 B.n621 VSUBS 0.008669f
C662 B.n622 VSUBS 0.008669f
C663 B.n623 VSUBS 0.008669f
C664 B.n624 VSUBS 0.008669f
C665 B.n625 VSUBS 0.008669f
C666 B.n626 VSUBS 0.008669f
C667 B.n627 VSUBS 0.008669f
C668 B.n628 VSUBS 0.008669f
C669 B.n629 VSUBS 0.008669f
C670 B.n630 VSUBS 0.008669f
C671 B.n631 VSUBS 0.008669f
C672 B.n632 VSUBS 0.008669f
C673 B.n633 VSUBS 0.008669f
C674 B.n634 VSUBS 0.008669f
C675 B.n635 VSUBS 0.008669f
C676 B.n636 VSUBS 0.008669f
C677 B.n637 VSUBS 0.008669f
C678 B.n638 VSUBS 0.008669f
C679 B.n639 VSUBS 0.008669f
C680 B.n640 VSUBS 0.008669f
C681 B.n641 VSUBS 0.008669f
C682 B.n642 VSUBS 0.008669f
C683 B.n643 VSUBS 0.008669f
C684 B.n644 VSUBS 0.008669f
C685 B.n645 VSUBS 0.008669f
C686 B.n646 VSUBS 0.008669f
C687 B.n647 VSUBS 0.008669f
C688 B.n648 VSUBS 0.008669f
C689 B.n649 VSUBS 0.008669f
C690 B.n650 VSUBS 0.008669f
C691 B.n651 VSUBS 0.008669f
C692 B.n652 VSUBS 0.008669f
C693 B.n653 VSUBS 0.008669f
C694 B.n654 VSUBS 0.008669f
C695 B.n655 VSUBS 0.008669f
C696 B.n656 VSUBS 0.008669f
C697 B.n657 VSUBS 0.008669f
C698 B.n658 VSUBS 0.008669f
C699 B.n659 VSUBS 0.008669f
C700 B.n660 VSUBS 0.008669f
C701 B.n661 VSUBS 0.008669f
C702 B.n662 VSUBS 0.008669f
C703 B.n663 VSUBS 0.008669f
C704 B.n664 VSUBS 0.008669f
C705 B.n665 VSUBS 0.019717f
C706 B.n666 VSUBS 0.02108f
C707 B.n667 VSUBS 0.02108f
C708 B.n668 VSUBS 0.008669f
C709 B.n669 VSUBS 0.008669f
C710 B.n670 VSUBS 0.008669f
C711 B.n671 VSUBS 0.008669f
C712 B.n672 VSUBS 0.008669f
C713 B.n673 VSUBS 0.008669f
C714 B.n674 VSUBS 0.008669f
C715 B.n675 VSUBS 0.008669f
C716 B.n676 VSUBS 0.008669f
C717 B.n677 VSUBS 0.008669f
C718 B.n678 VSUBS 0.008669f
C719 B.n679 VSUBS 0.008669f
C720 B.n680 VSUBS 0.008669f
C721 B.n681 VSUBS 0.008669f
C722 B.n682 VSUBS 0.008669f
C723 B.n683 VSUBS 0.008669f
C724 B.n684 VSUBS 0.008669f
C725 B.n685 VSUBS 0.008669f
C726 B.n686 VSUBS 0.008669f
C727 B.n687 VSUBS 0.008669f
C728 B.n688 VSUBS 0.008669f
C729 B.n689 VSUBS 0.008669f
C730 B.n690 VSUBS 0.008669f
C731 B.n691 VSUBS 0.008669f
C732 B.n692 VSUBS 0.008669f
C733 B.n693 VSUBS 0.008669f
C734 B.n694 VSUBS 0.008669f
C735 B.n695 VSUBS 0.008669f
C736 B.n696 VSUBS 0.008669f
C737 B.n697 VSUBS 0.008669f
C738 B.n698 VSUBS 0.008669f
C739 B.n699 VSUBS 0.008669f
C740 B.n700 VSUBS 0.008669f
C741 B.n701 VSUBS 0.008669f
C742 B.n702 VSUBS 0.008669f
C743 B.n703 VSUBS 0.008669f
C744 B.n704 VSUBS 0.008669f
C745 B.n705 VSUBS 0.008669f
C746 B.n706 VSUBS 0.008669f
C747 B.n707 VSUBS 0.008669f
C748 B.n708 VSUBS 0.008669f
C749 B.n709 VSUBS 0.008669f
C750 B.n710 VSUBS 0.008669f
C751 B.n711 VSUBS 0.008669f
C752 B.n712 VSUBS 0.008669f
C753 B.n713 VSUBS 0.008669f
C754 B.n714 VSUBS 0.008669f
C755 B.n715 VSUBS 0.008159f
C756 B.n716 VSUBS 0.020086f
C757 B.n717 VSUBS 0.004845f
C758 B.n718 VSUBS 0.008669f
C759 B.n719 VSUBS 0.008669f
C760 B.n720 VSUBS 0.008669f
C761 B.n721 VSUBS 0.008669f
C762 B.n722 VSUBS 0.008669f
C763 B.n723 VSUBS 0.008669f
C764 B.n724 VSUBS 0.008669f
C765 B.n725 VSUBS 0.008669f
C766 B.n726 VSUBS 0.008669f
C767 B.n727 VSUBS 0.008669f
C768 B.n728 VSUBS 0.008669f
C769 B.n729 VSUBS 0.008669f
C770 B.n730 VSUBS 0.004845f
C771 B.n731 VSUBS 0.008669f
C772 B.n732 VSUBS 0.008669f
C773 B.n733 VSUBS 0.008159f
C774 B.n734 VSUBS 0.008669f
C775 B.n735 VSUBS 0.008669f
C776 B.n736 VSUBS 0.008669f
C777 B.n737 VSUBS 0.008669f
C778 B.n738 VSUBS 0.008669f
C779 B.n739 VSUBS 0.008669f
C780 B.n740 VSUBS 0.008669f
C781 B.n741 VSUBS 0.008669f
C782 B.n742 VSUBS 0.008669f
C783 B.n743 VSUBS 0.008669f
C784 B.n744 VSUBS 0.008669f
C785 B.n745 VSUBS 0.008669f
C786 B.n746 VSUBS 0.008669f
C787 B.n747 VSUBS 0.008669f
C788 B.n748 VSUBS 0.008669f
C789 B.n749 VSUBS 0.008669f
C790 B.n750 VSUBS 0.008669f
C791 B.n751 VSUBS 0.008669f
C792 B.n752 VSUBS 0.008669f
C793 B.n753 VSUBS 0.008669f
C794 B.n754 VSUBS 0.008669f
C795 B.n755 VSUBS 0.008669f
C796 B.n756 VSUBS 0.008669f
C797 B.n757 VSUBS 0.008669f
C798 B.n758 VSUBS 0.008669f
C799 B.n759 VSUBS 0.008669f
C800 B.n760 VSUBS 0.008669f
C801 B.n761 VSUBS 0.008669f
C802 B.n762 VSUBS 0.008669f
C803 B.n763 VSUBS 0.008669f
C804 B.n764 VSUBS 0.008669f
C805 B.n765 VSUBS 0.008669f
C806 B.n766 VSUBS 0.008669f
C807 B.n767 VSUBS 0.008669f
C808 B.n768 VSUBS 0.008669f
C809 B.n769 VSUBS 0.008669f
C810 B.n770 VSUBS 0.008669f
C811 B.n771 VSUBS 0.008669f
C812 B.n772 VSUBS 0.008669f
C813 B.n773 VSUBS 0.008669f
C814 B.n774 VSUBS 0.008669f
C815 B.n775 VSUBS 0.008669f
C816 B.n776 VSUBS 0.008669f
C817 B.n777 VSUBS 0.008669f
C818 B.n778 VSUBS 0.008669f
C819 B.n779 VSUBS 0.008669f
C820 B.n780 VSUBS 0.02108f
C821 B.n781 VSUBS 0.02108f
C822 B.n782 VSUBS 0.019717f
C823 B.n783 VSUBS 0.008669f
C824 B.n784 VSUBS 0.008669f
C825 B.n785 VSUBS 0.008669f
C826 B.n786 VSUBS 0.008669f
C827 B.n787 VSUBS 0.008669f
C828 B.n788 VSUBS 0.008669f
C829 B.n789 VSUBS 0.008669f
C830 B.n790 VSUBS 0.008669f
C831 B.n791 VSUBS 0.008669f
C832 B.n792 VSUBS 0.008669f
C833 B.n793 VSUBS 0.008669f
C834 B.n794 VSUBS 0.008669f
C835 B.n795 VSUBS 0.008669f
C836 B.n796 VSUBS 0.008669f
C837 B.n797 VSUBS 0.008669f
C838 B.n798 VSUBS 0.008669f
C839 B.n799 VSUBS 0.008669f
C840 B.n800 VSUBS 0.008669f
C841 B.n801 VSUBS 0.008669f
C842 B.n802 VSUBS 0.008669f
C843 B.n803 VSUBS 0.008669f
C844 B.n804 VSUBS 0.008669f
C845 B.n805 VSUBS 0.008669f
C846 B.n806 VSUBS 0.008669f
C847 B.n807 VSUBS 0.008669f
C848 B.n808 VSUBS 0.008669f
C849 B.n809 VSUBS 0.008669f
C850 B.n810 VSUBS 0.008669f
C851 B.n811 VSUBS 0.008669f
C852 B.n812 VSUBS 0.008669f
C853 B.n813 VSUBS 0.008669f
C854 B.n814 VSUBS 0.008669f
C855 B.n815 VSUBS 0.008669f
C856 B.n816 VSUBS 0.008669f
C857 B.n817 VSUBS 0.008669f
C858 B.n818 VSUBS 0.008669f
C859 B.n819 VSUBS 0.008669f
C860 B.n820 VSUBS 0.008669f
C861 B.n821 VSUBS 0.008669f
C862 B.n822 VSUBS 0.008669f
C863 B.n823 VSUBS 0.008669f
C864 B.n824 VSUBS 0.008669f
C865 B.n825 VSUBS 0.008669f
C866 B.n826 VSUBS 0.008669f
C867 B.n827 VSUBS 0.008669f
C868 B.n828 VSUBS 0.008669f
C869 B.n829 VSUBS 0.008669f
C870 B.n830 VSUBS 0.008669f
C871 B.n831 VSUBS 0.008669f
C872 B.n832 VSUBS 0.008669f
C873 B.n833 VSUBS 0.008669f
C874 B.n834 VSUBS 0.008669f
C875 B.n835 VSUBS 0.008669f
C876 B.n836 VSUBS 0.008669f
C877 B.n837 VSUBS 0.008669f
C878 B.n838 VSUBS 0.008669f
C879 B.n839 VSUBS 0.008669f
C880 B.n840 VSUBS 0.008669f
C881 B.n841 VSUBS 0.008669f
C882 B.n842 VSUBS 0.008669f
C883 B.n843 VSUBS 0.008669f
C884 B.n844 VSUBS 0.008669f
C885 B.n845 VSUBS 0.008669f
C886 B.n846 VSUBS 0.008669f
C887 B.n847 VSUBS 0.008669f
C888 B.n848 VSUBS 0.008669f
C889 B.n849 VSUBS 0.008669f
C890 B.n850 VSUBS 0.008669f
C891 B.n851 VSUBS 0.008669f
C892 B.n852 VSUBS 0.008669f
C893 B.n853 VSUBS 0.008669f
C894 B.n854 VSUBS 0.008669f
C895 B.n855 VSUBS 0.008669f
C896 B.n856 VSUBS 0.008669f
C897 B.n857 VSUBS 0.008669f
C898 B.n858 VSUBS 0.008669f
C899 B.n859 VSUBS 0.008669f
C900 B.n860 VSUBS 0.008669f
C901 B.n861 VSUBS 0.008669f
C902 B.n862 VSUBS 0.008669f
C903 B.n863 VSUBS 0.008669f
C904 B.n864 VSUBS 0.008669f
C905 B.n865 VSUBS 0.008669f
C906 B.n866 VSUBS 0.008669f
C907 B.n867 VSUBS 0.008669f
C908 B.n868 VSUBS 0.008669f
C909 B.n869 VSUBS 0.008669f
C910 B.n870 VSUBS 0.008669f
C911 B.n871 VSUBS 0.008669f
C912 B.n872 VSUBS 0.008669f
C913 B.n873 VSUBS 0.008669f
C914 B.n874 VSUBS 0.008669f
C915 B.n875 VSUBS 0.008669f
C916 B.n876 VSUBS 0.008669f
C917 B.n877 VSUBS 0.008669f
C918 B.n878 VSUBS 0.008669f
C919 B.n879 VSUBS 0.008669f
C920 B.n880 VSUBS 0.008669f
C921 B.n881 VSUBS 0.008669f
C922 B.n882 VSUBS 0.008669f
C923 B.n883 VSUBS 0.008669f
C924 B.n884 VSUBS 0.008669f
C925 B.n885 VSUBS 0.008669f
C926 B.n886 VSUBS 0.008669f
C927 B.n887 VSUBS 0.011313f
C928 B.n888 VSUBS 0.012051f
C929 B.n889 VSUBS 0.023965f
C930 VDD2.t1 VSUBS 0.25351f
C931 VDD2.t4 VSUBS 0.25351f
C932 VDD2.n0 VSUBS 1.92092f
C933 VDD2.t0 VSUBS 0.25351f
C934 VDD2.t3 VSUBS 0.25351f
C935 VDD2.n1 VSUBS 1.92092f
C936 VDD2.n2 VSUBS 6.1263f
C937 VDD2.t7 VSUBS 0.25351f
C938 VDD2.t6 VSUBS 0.25351f
C939 VDD2.n3 VSUBS 1.89457f
C940 VDD2.n4 VSUBS 4.8434f
C941 VDD2.t2 VSUBS 0.25351f
C942 VDD2.t5 VSUBS 0.25351f
C943 VDD2.n5 VSUBS 1.92086f
C944 VN.n0 VSUBS 0.04849f
C945 VN.t4 VSUBS 2.52993f
C946 VN.n1 VSUBS 0.048046f
C947 VN.n2 VSUBS 0.025779f
C948 VN.n3 VSUBS 0.048046f
C949 VN.n4 VSUBS 0.025779f
C950 VN.t7 VSUBS 2.52993f
C951 VN.n5 VSUBS 0.048046f
C952 VN.n6 VSUBS 0.025779f
C953 VN.n7 VSUBS 0.048046f
C954 VN.n8 VSUBS 0.340658f
C955 VN.t3 VSUBS 2.52993f
C956 VN.t6 VSUBS 2.93752f
C957 VN.n9 VSUBS 0.948596f
C958 VN.n10 VSUBS 0.989316f
C959 VN.n11 VSUBS 0.031916f
C960 VN.n12 VSUBS 0.048046f
C961 VN.n13 VSUBS 0.025779f
C962 VN.n14 VSUBS 0.025779f
C963 VN.n15 VSUBS 0.025779f
C964 VN.n16 VSUBS 0.051236f
C965 VN.n17 VSUBS 0.02084f
C966 VN.n18 VSUBS 0.051236f
C967 VN.n19 VSUBS 0.025779f
C968 VN.n20 VSUBS 0.025779f
C969 VN.n21 VSUBS 0.025779f
C970 VN.n22 VSUBS 0.048046f
C971 VN.n23 VSUBS 0.031916f
C972 VN.n24 VSUBS 0.89906f
C973 VN.n25 VSUBS 0.040455f
C974 VN.n26 VSUBS 0.025779f
C975 VN.n27 VSUBS 0.025779f
C976 VN.n28 VSUBS 0.025779f
C977 VN.n29 VSUBS 0.048046f
C978 VN.n30 VSUBS 0.042661f
C979 VN.n31 VSUBS 0.032604f
C980 VN.n32 VSUBS 0.025779f
C981 VN.n33 VSUBS 0.025779f
C982 VN.n34 VSUBS 0.025779f
C983 VN.n35 VSUBS 0.048046f
C984 VN.n36 VSUBS 0.047097f
C985 VN.n37 VSUBS 1.01875f
C986 VN.n38 VSUBS 0.077452f
C987 VN.n39 VSUBS 0.04849f
C988 VN.t0 VSUBS 2.52993f
C989 VN.n40 VSUBS 0.048046f
C990 VN.n41 VSUBS 0.025779f
C991 VN.n42 VSUBS 0.048046f
C992 VN.n43 VSUBS 0.025779f
C993 VN.t1 VSUBS 2.52993f
C994 VN.n44 VSUBS 0.048046f
C995 VN.n45 VSUBS 0.025779f
C996 VN.n46 VSUBS 0.048046f
C997 VN.n47 VSUBS 0.340658f
C998 VN.t5 VSUBS 2.52993f
C999 VN.t2 VSUBS 2.93752f
C1000 VN.n48 VSUBS 0.948596f
C1001 VN.n49 VSUBS 0.989316f
C1002 VN.n50 VSUBS 0.031916f
C1003 VN.n51 VSUBS 0.048046f
C1004 VN.n52 VSUBS 0.025779f
C1005 VN.n53 VSUBS 0.025779f
C1006 VN.n54 VSUBS 0.025779f
C1007 VN.n55 VSUBS 0.051236f
C1008 VN.n56 VSUBS 0.02084f
C1009 VN.n57 VSUBS 0.051236f
C1010 VN.n58 VSUBS 0.025779f
C1011 VN.n59 VSUBS 0.025779f
C1012 VN.n60 VSUBS 0.025779f
C1013 VN.n61 VSUBS 0.048046f
C1014 VN.n62 VSUBS 0.031916f
C1015 VN.n63 VSUBS 0.89906f
C1016 VN.n64 VSUBS 0.040455f
C1017 VN.n65 VSUBS 0.025779f
C1018 VN.n66 VSUBS 0.025779f
C1019 VN.n67 VSUBS 0.025779f
C1020 VN.n68 VSUBS 0.048046f
C1021 VN.n69 VSUBS 0.042661f
C1022 VN.n70 VSUBS 0.032604f
C1023 VN.n71 VSUBS 0.025779f
C1024 VN.n72 VSUBS 0.025779f
C1025 VN.n73 VSUBS 0.025779f
C1026 VN.n74 VSUBS 0.048046f
C1027 VN.n75 VSUBS 0.047097f
C1028 VN.n76 VSUBS 1.01875f
C1029 VN.n77 VSUBS 1.73654f
C1030 VTAIL.t6 VSUBS 0.20073f
C1031 VTAIL.t1 VSUBS 0.20073f
C1032 VTAIL.n0 VSUBS 1.38209f
C1033 VTAIL.n1 VSUBS 0.900771f
C1034 VTAIL.t3 VSUBS 1.84235f
C1035 VTAIL.n2 VSUBS 1.02494f
C1036 VTAIL.t12 VSUBS 1.84235f
C1037 VTAIL.n3 VSUBS 1.02494f
C1038 VTAIL.t11 VSUBS 0.20073f
C1039 VTAIL.t14 VSUBS 0.20073f
C1040 VTAIL.n4 VSUBS 1.38209f
C1041 VTAIL.n5 VSUBS 1.23014f
C1042 VTAIL.t13 VSUBS 1.84235f
C1043 VTAIL.n6 VSUBS 2.40168f
C1044 VTAIL.t5 VSUBS 1.84236f
C1045 VTAIL.n7 VSUBS 2.40167f
C1046 VTAIL.t2 VSUBS 0.20073f
C1047 VTAIL.t0 VSUBS 0.20073f
C1048 VTAIL.n8 VSUBS 1.38209f
C1049 VTAIL.n9 VSUBS 1.23014f
C1050 VTAIL.t4 VSUBS 1.84236f
C1051 VTAIL.n10 VSUBS 1.02493f
C1052 VTAIL.t9 VSUBS 1.84236f
C1053 VTAIL.n11 VSUBS 1.02493f
C1054 VTAIL.t10 VSUBS 0.20073f
C1055 VTAIL.t15 VSUBS 0.20073f
C1056 VTAIL.n12 VSUBS 1.38209f
C1057 VTAIL.n13 VSUBS 1.23014f
C1058 VTAIL.t8 VSUBS 1.84235f
C1059 VTAIL.n14 VSUBS 2.40168f
C1060 VTAIL.t7 VSUBS 1.84235f
C1061 VTAIL.n15 VSUBS 2.39645f
C1062 VDD1.t4 VSUBS 0.230566f
C1063 VDD1.t7 VSUBS 0.230566f
C1064 VDD1.n0 VSUBS 1.74879f
C1065 VDD1.t6 VSUBS 0.230566f
C1066 VDD1.t1 VSUBS 0.230566f
C1067 VDD1.n1 VSUBS 1.74706f
C1068 VDD1.t3 VSUBS 0.230566f
C1069 VDD1.t5 VSUBS 0.230566f
C1070 VDD1.n2 VSUBS 1.74706f
C1071 VDD1.n3 VSUBS 5.63774f
C1072 VDD1.t0 VSUBS 0.230566f
C1073 VDD1.t2 VSUBS 0.230566f
C1074 VDD1.n4 VSUBS 1.72309f
C1075 VDD1.n5 VSUBS 4.44542f
C1076 VP.n0 VSUBS 0.053903f
C1077 VP.t3 VSUBS 2.81233f
C1078 VP.n1 VSUBS 0.053409f
C1079 VP.n2 VSUBS 0.028657f
C1080 VP.n3 VSUBS 0.053409f
C1081 VP.n4 VSUBS 0.028657f
C1082 VP.t1 VSUBS 2.81233f
C1083 VP.n5 VSUBS 0.053409f
C1084 VP.n6 VSUBS 0.028657f
C1085 VP.n7 VSUBS 0.053409f
C1086 VP.n8 VSUBS 0.028657f
C1087 VP.t4 VSUBS 2.81233f
C1088 VP.n9 VSUBS 0.053409f
C1089 VP.n10 VSUBS 0.028657f
C1090 VP.n11 VSUBS 0.053409f
C1091 VP.n12 VSUBS 0.053903f
C1092 VP.t2 VSUBS 2.81233f
C1093 VP.n13 VSUBS 0.053903f
C1094 VP.t7 VSUBS 2.81233f
C1095 VP.n14 VSUBS 0.053409f
C1096 VP.n15 VSUBS 0.028657f
C1097 VP.n16 VSUBS 0.053409f
C1098 VP.n17 VSUBS 0.028657f
C1099 VP.t0 VSUBS 2.81233f
C1100 VP.n18 VSUBS 0.053409f
C1101 VP.n19 VSUBS 0.028657f
C1102 VP.n20 VSUBS 0.053409f
C1103 VP.n21 VSUBS 0.378684f
C1104 VP.t5 VSUBS 2.81233f
C1105 VP.t6 VSUBS 3.26541f
C1106 VP.n22 VSUBS 1.05448f
C1107 VP.n23 VSUBS 1.09975f
C1108 VP.n24 VSUBS 0.035478f
C1109 VP.n25 VSUBS 0.053409f
C1110 VP.n26 VSUBS 0.028657f
C1111 VP.n27 VSUBS 0.028657f
C1112 VP.n28 VSUBS 0.028657f
C1113 VP.n29 VSUBS 0.056955f
C1114 VP.n30 VSUBS 0.023166f
C1115 VP.n31 VSUBS 0.056955f
C1116 VP.n32 VSUBS 0.028657f
C1117 VP.n33 VSUBS 0.028657f
C1118 VP.n34 VSUBS 0.028657f
C1119 VP.n35 VSUBS 0.053409f
C1120 VP.n36 VSUBS 0.035478f
C1121 VP.n37 VSUBS 0.999416f
C1122 VP.n38 VSUBS 0.044971f
C1123 VP.n39 VSUBS 0.028657f
C1124 VP.n40 VSUBS 0.028657f
C1125 VP.n41 VSUBS 0.028657f
C1126 VP.n42 VSUBS 0.053409f
C1127 VP.n43 VSUBS 0.047423f
C1128 VP.n44 VSUBS 0.036244f
C1129 VP.n45 VSUBS 0.028657f
C1130 VP.n46 VSUBS 0.028657f
C1131 VP.n47 VSUBS 0.028657f
C1132 VP.n48 VSUBS 0.053409f
C1133 VP.n49 VSUBS 0.052354f
C1134 VP.n50 VSUBS 1.13247f
C1135 VP.n51 VSUBS 1.92347f
C1136 VP.n52 VSUBS 1.94203f
C1137 VP.n53 VSUBS 1.13247f
C1138 VP.n54 VSUBS 0.052354f
C1139 VP.n55 VSUBS 0.053409f
C1140 VP.n56 VSUBS 0.028657f
C1141 VP.n57 VSUBS 0.028657f
C1142 VP.n58 VSUBS 0.028657f
C1143 VP.n59 VSUBS 0.036244f
C1144 VP.n60 VSUBS 0.047423f
C1145 VP.n61 VSUBS 0.053409f
C1146 VP.n62 VSUBS 0.028657f
C1147 VP.n63 VSUBS 0.028657f
C1148 VP.n64 VSUBS 0.028657f
C1149 VP.n65 VSUBS 0.044971f
C1150 VP.n66 VSUBS 0.999416f
C1151 VP.n67 VSUBS 0.035478f
C1152 VP.n68 VSUBS 0.053409f
C1153 VP.n69 VSUBS 0.028657f
C1154 VP.n70 VSUBS 0.028657f
C1155 VP.n71 VSUBS 0.028657f
C1156 VP.n72 VSUBS 0.056955f
C1157 VP.n73 VSUBS 0.023166f
C1158 VP.n74 VSUBS 0.056955f
C1159 VP.n75 VSUBS 0.028657f
C1160 VP.n76 VSUBS 0.028657f
C1161 VP.n77 VSUBS 0.028657f
C1162 VP.n78 VSUBS 0.053409f
C1163 VP.n79 VSUBS 0.035478f
C1164 VP.n80 VSUBS 0.999416f
C1165 VP.n81 VSUBS 0.044971f
C1166 VP.n82 VSUBS 0.028657f
C1167 VP.n83 VSUBS 0.028657f
C1168 VP.n84 VSUBS 0.028657f
C1169 VP.n85 VSUBS 0.053409f
C1170 VP.n86 VSUBS 0.047423f
C1171 VP.n87 VSUBS 0.036244f
C1172 VP.n88 VSUBS 0.028657f
C1173 VP.n89 VSUBS 0.028657f
C1174 VP.n90 VSUBS 0.028657f
C1175 VP.n91 VSUBS 0.053409f
C1176 VP.n92 VSUBS 0.052354f
C1177 VP.n93 VSUBS 1.13247f
C1178 VP.n94 VSUBS 0.086098f
.ends

