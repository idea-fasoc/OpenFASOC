* NGSPICE file created from diff_pair_sample_0566.ext - technology: sky130A

.subckt diff_pair_sample_0566 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=1.55
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=3.8727 ps=20.64 w=9.93 l=1.55
X2 B.t8 B.t6 B.t7 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=1.55
X3 B.t5 B.t3 B.t4 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=1.55
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=3.8727 ps=20.64 w=9.93 l=1.55
X5 B.t2 B.t0 B.t1 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=1.55
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=3.8727 ps=20.64 w=9.93 l=1.55
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n1722_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=3.8727 ps=20.64 w=9.93 l=1.55
R0 B.n339 B.n56 585
R1 B.n341 B.n340 585
R2 B.n342 B.n55 585
R3 B.n344 B.n343 585
R4 B.n345 B.n54 585
R5 B.n347 B.n346 585
R6 B.n348 B.n53 585
R7 B.n350 B.n349 585
R8 B.n351 B.n52 585
R9 B.n353 B.n352 585
R10 B.n354 B.n51 585
R11 B.n356 B.n355 585
R12 B.n357 B.n50 585
R13 B.n359 B.n358 585
R14 B.n360 B.n49 585
R15 B.n362 B.n361 585
R16 B.n363 B.n48 585
R17 B.n365 B.n364 585
R18 B.n366 B.n47 585
R19 B.n368 B.n367 585
R20 B.n369 B.n46 585
R21 B.n371 B.n370 585
R22 B.n372 B.n45 585
R23 B.n374 B.n373 585
R24 B.n375 B.n44 585
R25 B.n377 B.n376 585
R26 B.n378 B.n43 585
R27 B.n380 B.n379 585
R28 B.n381 B.n42 585
R29 B.n383 B.n382 585
R30 B.n384 B.n41 585
R31 B.n386 B.n385 585
R32 B.n387 B.n40 585
R33 B.n389 B.n388 585
R34 B.n390 B.n39 585
R35 B.n392 B.n391 585
R36 B.n394 B.n393 585
R37 B.n395 B.n35 585
R38 B.n397 B.n396 585
R39 B.n398 B.n34 585
R40 B.n400 B.n399 585
R41 B.n401 B.n33 585
R42 B.n403 B.n402 585
R43 B.n404 B.n32 585
R44 B.n406 B.n405 585
R45 B.n408 B.n29 585
R46 B.n410 B.n409 585
R47 B.n411 B.n28 585
R48 B.n413 B.n412 585
R49 B.n414 B.n27 585
R50 B.n416 B.n415 585
R51 B.n417 B.n26 585
R52 B.n419 B.n418 585
R53 B.n420 B.n25 585
R54 B.n422 B.n421 585
R55 B.n423 B.n24 585
R56 B.n425 B.n424 585
R57 B.n426 B.n23 585
R58 B.n428 B.n427 585
R59 B.n429 B.n22 585
R60 B.n431 B.n430 585
R61 B.n432 B.n21 585
R62 B.n434 B.n433 585
R63 B.n435 B.n20 585
R64 B.n437 B.n436 585
R65 B.n438 B.n19 585
R66 B.n440 B.n439 585
R67 B.n441 B.n18 585
R68 B.n443 B.n442 585
R69 B.n444 B.n17 585
R70 B.n446 B.n445 585
R71 B.n447 B.n16 585
R72 B.n449 B.n448 585
R73 B.n450 B.n15 585
R74 B.n452 B.n451 585
R75 B.n453 B.n14 585
R76 B.n455 B.n454 585
R77 B.n456 B.n13 585
R78 B.n458 B.n457 585
R79 B.n459 B.n12 585
R80 B.n461 B.n460 585
R81 B.n338 B.n337 585
R82 B.n336 B.n57 585
R83 B.n335 B.n334 585
R84 B.n333 B.n58 585
R85 B.n332 B.n331 585
R86 B.n330 B.n59 585
R87 B.n329 B.n328 585
R88 B.n327 B.n60 585
R89 B.n326 B.n325 585
R90 B.n324 B.n61 585
R91 B.n323 B.n322 585
R92 B.n321 B.n62 585
R93 B.n320 B.n319 585
R94 B.n318 B.n63 585
R95 B.n317 B.n316 585
R96 B.n315 B.n64 585
R97 B.n314 B.n313 585
R98 B.n312 B.n65 585
R99 B.n311 B.n310 585
R100 B.n309 B.n66 585
R101 B.n308 B.n307 585
R102 B.n306 B.n67 585
R103 B.n305 B.n304 585
R104 B.n303 B.n68 585
R105 B.n302 B.n301 585
R106 B.n300 B.n69 585
R107 B.n299 B.n298 585
R108 B.n297 B.n70 585
R109 B.n296 B.n295 585
R110 B.n294 B.n71 585
R111 B.n293 B.n292 585
R112 B.n291 B.n72 585
R113 B.n290 B.n289 585
R114 B.n288 B.n73 585
R115 B.n287 B.n286 585
R116 B.n285 B.n74 585
R117 B.n284 B.n283 585
R118 B.n282 B.n75 585
R119 B.n281 B.n280 585
R120 B.n158 B.n157 585
R121 B.n159 B.n120 585
R122 B.n161 B.n160 585
R123 B.n162 B.n119 585
R124 B.n164 B.n163 585
R125 B.n165 B.n118 585
R126 B.n167 B.n166 585
R127 B.n168 B.n117 585
R128 B.n170 B.n169 585
R129 B.n171 B.n116 585
R130 B.n173 B.n172 585
R131 B.n174 B.n115 585
R132 B.n176 B.n175 585
R133 B.n177 B.n114 585
R134 B.n179 B.n178 585
R135 B.n180 B.n113 585
R136 B.n182 B.n181 585
R137 B.n183 B.n112 585
R138 B.n185 B.n184 585
R139 B.n186 B.n111 585
R140 B.n188 B.n187 585
R141 B.n189 B.n110 585
R142 B.n191 B.n190 585
R143 B.n192 B.n109 585
R144 B.n194 B.n193 585
R145 B.n195 B.n108 585
R146 B.n197 B.n196 585
R147 B.n198 B.n107 585
R148 B.n200 B.n199 585
R149 B.n201 B.n106 585
R150 B.n203 B.n202 585
R151 B.n204 B.n105 585
R152 B.n206 B.n205 585
R153 B.n207 B.n104 585
R154 B.n209 B.n208 585
R155 B.n210 B.n101 585
R156 B.n213 B.n212 585
R157 B.n214 B.n100 585
R158 B.n216 B.n215 585
R159 B.n217 B.n99 585
R160 B.n219 B.n218 585
R161 B.n220 B.n98 585
R162 B.n222 B.n221 585
R163 B.n223 B.n97 585
R164 B.n225 B.n224 585
R165 B.n227 B.n226 585
R166 B.n228 B.n93 585
R167 B.n230 B.n229 585
R168 B.n231 B.n92 585
R169 B.n233 B.n232 585
R170 B.n234 B.n91 585
R171 B.n236 B.n235 585
R172 B.n237 B.n90 585
R173 B.n239 B.n238 585
R174 B.n240 B.n89 585
R175 B.n242 B.n241 585
R176 B.n243 B.n88 585
R177 B.n245 B.n244 585
R178 B.n246 B.n87 585
R179 B.n248 B.n247 585
R180 B.n249 B.n86 585
R181 B.n251 B.n250 585
R182 B.n252 B.n85 585
R183 B.n254 B.n253 585
R184 B.n255 B.n84 585
R185 B.n257 B.n256 585
R186 B.n258 B.n83 585
R187 B.n260 B.n259 585
R188 B.n261 B.n82 585
R189 B.n263 B.n262 585
R190 B.n264 B.n81 585
R191 B.n266 B.n265 585
R192 B.n267 B.n80 585
R193 B.n269 B.n268 585
R194 B.n270 B.n79 585
R195 B.n272 B.n271 585
R196 B.n273 B.n78 585
R197 B.n275 B.n274 585
R198 B.n276 B.n77 585
R199 B.n278 B.n277 585
R200 B.n279 B.n76 585
R201 B.n156 B.n121 585
R202 B.n155 B.n154 585
R203 B.n153 B.n122 585
R204 B.n152 B.n151 585
R205 B.n150 B.n123 585
R206 B.n149 B.n148 585
R207 B.n147 B.n124 585
R208 B.n146 B.n145 585
R209 B.n144 B.n125 585
R210 B.n143 B.n142 585
R211 B.n141 B.n126 585
R212 B.n140 B.n139 585
R213 B.n138 B.n127 585
R214 B.n137 B.n136 585
R215 B.n135 B.n128 585
R216 B.n134 B.n133 585
R217 B.n132 B.n129 585
R218 B.n131 B.n130 585
R219 B.n2 B.n0 585
R220 B.n489 B.n1 585
R221 B.n488 B.n487 585
R222 B.n486 B.n3 585
R223 B.n485 B.n484 585
R224 B.n483 B.n4 585
R225 B.n482 B.n481 585
R226 B.n480 B.n5 585
R227 B.n479 B.n478 585
R228 B.n477 B.n6 585
R229 B.n476 B.n475 585
R230 B.n474 B.n7 585
R231 B.n473 B.n472 585
R232 B.n471 B.n8 585
R233 B.n470 B.n469 585
R234 B.n468 B.n9 585
R235 B.n467 B.n466 585
R236 B.n465 B.n10 585
R237 B.n464 B.n463 585
R238 B.n462 B.n11 585
R239 B.n491 B.n490 585
R240 B.n158 B.n121 497.305
R241 B.n460 B.n11 497.305
R242 B.n280 B.n279 497.305
R243 B.n339 B.n338 497.305
R244 B.n94 B.t5 374.68
R245 B.n36 B.t10 374.68
R246 B.n102 B.t2 374.68
R247 B.n30 B.t7 374.68
R248 B.n94 B.t3 360.017
R249 B.n102 B.t0 360.017
R250 B.n30 B.t6 360.017
R251 B.n36 B.t9 360.017
R252 B.n95 B.t4 338.219
R253 B.n37 B.t11 338.219
R254 B.n103 B.t1 338.219
R255 B.n31 B.t8 338.219
R256 B.n154 B.n121 163.367
R257 B.n154 B.n153 163.367
R258 B.n153 B.n152 163.367
R259 B.n152 B.n123 163.367
R260 B.n148 B.n123 163.367
R261 B.n148 B.n147 163.367
R262 B.n147 B.n146 163.367
R263 B.n146 B.n125 163.367
R264 B.n142 B.n125 163.367
R265 B.n142 B.n141 163.367
R266 B.n141 B.n140 163.367
R267 B.n140 B.n127 163.367
R268 B.n136 B.n127 163.367
R269 B.n136 B.n135 163.367
R270 B.n135 B.n134 163.367
R271 B.n134 B.n129 163.367
R272 B.n130 B.n129 163.367
R273 B.n130 B.n2 163.367
R274 B.n490 B.n2 163.367
R275 B.n490 B.n489 163.367
R276 B.n489 B.n488 163.367
R277 B.n488 B.n3 163.367
R278 B.n484 B.n3 163.367
R279 B.n484 B.n483 163.367
R280 B.n483 B.n482 163.367
R281 B.n482 B.n5 163.367
R282 B.n478 B.n5 163.367
R283 B.n478 B.n477 163.367
R284 B.n477 B.n476 163.367
R285 B.n476 B.n7 163.367
R286 B.n472 B.n7 163.367
R287 B.n472 B.n471 163.367
R288 B.n471 B.n470 163.367
R289 B.n470 B.n9 163.367
R290 B.n466 B.n9 163.367
R291 B.n466 B.n465 163.367
R292 B.n465 B.n464 163.367
R293 B.n464 B.n11 163.367
R294 B.n159 B.n158 163.367
R295 B.n160 B.n159 163.367
R296 B.n160 B.n119 163.367
R297 B.n164 B.n119 163.367
R298 B.n165 B.n164 163.367
R299 B.n166 B.n165 163.367
R300 B.n166 B.n117 163.367
R301 B.n170 B.n117 163.367
R302 B.n171 B.n170 163.367
R303 B.n172 B.n171 163.367
R304 B.n172 B.n115 163.367
R305 B.n176 B.n115 163.367
R306 B.n177 B.n176 163.367
R307 B.n178 B.n177 163.367
R308 B.n178 B.n113 163.367
R309 B.n182 B.n113 163.367
R310 B.n183 B.n182 163.367
R311 B.n184 B.n183 163.367
R312 B.n184 B.n111 163.367
R313 B.n188 B.n111 163.367
R314 B.n189 B.n188 163.367
R315 B.n190 B.n189 163.367
R316 B.n190 B.n109 163.367
R317 B.n194 B.n109 163.367
R318 B.n195 B.n194 163.367
R319 B.n196 B.n195 163.367
R320 B.n196 B.n107 163.367
R321 B.n200 B.n107 163.367
R322 B.n201 B.n200 163.367
R323 B.n202 B.n201 163.367
R324 B.n202 B.n105 163.367
R325 B.n206 B.n105 163.367
R326 B.n207 B.n206 163.367
R327 B.n208 B.n207 163.367
R328 B.n208 B.n101 163.367
R329 B.n213 B.n101 163.367
R330 B.n214 B.n213 163.367
R331 B.n215 B.n214 163.367
R332 B.n215 B.n99 163.367
R333 B.n219 B.n99 163.367
R334 B.n220 B.n219 163.367
R335 B.n221 B.n220 163.367
R336 B.n221 B.n97 163.367
R337 B.n225 B.n97 163.367
R338 B.n226 B.n225 163.367
R339 B.n226 B.n93 163.367
R340 B.n230 B.n93 163.367
R341 B.n231 B.n230 163.367
R342 B.n232 B.n231 163.367
R343 B.n232 B.n91 163.367
R344 B.n236 B.n91 163.367
R345 B.n237 B.n236 163.367
R346 B.n238 B.n237 163.367
R347 B.n238 B.n89 163.367
R348 B.n242 B.n89 163.367
R349 B.n243 B.n242 163.367
R350 B.n244 B.n243 163.367
R351 B.n244 B.n87 163.367
R352 B.n248 B.n87 163.367
R353 B.n249 B.n248 163.367
R354 B.n250 B.n249 163.367
R355 B.n250 B.n85 163.367
R356 B.n254 B.n85 163.367
R357 B.n255 B.n254 163.367
R358 B.n256 B.n255 163.367
R359 B.n256 B.n83 163.367
R360 B.n260 B.n83 163.367
R361 B.n261 B.n260 163.367
R362 B.n262 B.n261 163.367
R363 B.n262 B.n81 163.367
R364 B.n266 B.n81 163.367
R365 B.n267 B.n266 163.367
R366 B.n268 B.n267 163.367
R367 B.n268 B.n79 163.367
R368 B.n272 B.n79 163.367
R369 B.n273 B.n272 163.367
R370 B.n274 B.n273 163.367
R371 B.n274 B.n77 163.367
R372 B.n278 B.n77 163.367
R373 B.n279 B.n278 163.367
R374 B.n280 B.n75 163.367
R375 B.n284 B.n75 163.367
R376 B.n285 B.n284 163.367
R377 B.n286 B.n285 163.367
R378 B.n286 B.n73 163.367
R379 B.n290 B.n73 163.367
R380 B.n291 B.n290 163.367
R381 B.n292 B.n291 163.367
R382 B.n292 B.n71 163.367
R383 B.n296 B.n71 163.367
R384 B.n297 B.n296 163.367
R385 B.n298 B.n297 163.367
R386 B.n298 B.n69 163.367
R387 B.n302 B.n69 163.367
R388 B.n303 B.n302 163.367
R389 B.n304 B.n303 163.367
R390 B.n304 B.n67 163.367
R391 B.n308 B.n67 163.367
R392 B.n309 B.n308 163.367
R393 B.n310 B.n309 163.367
R394 B.n310 B.n65 163.367
R395 B.n314 B.n65 163.367
R396 B.n315 B.n314 163.367
R397 B.n316 B.n315 163.367
R398 B.n316 B.n63 163.367
R399 B.n320 B.n63 163.367
R400 B.n321 B.n320 163.367
R401 B.n322 B.n321 163.367
R402 B.n322 B.n61 163.367
R403 B.n326 B.n61 163.367
R404 B.n327 B.n326 163.367
R405 B.n328 B.n327 163.367
R406 B.n328 B.n59 163.367
R407 B.n332 B.n59 163.367
R408 B.n333 B.n332 163.367
R409 B.n334 B.n333 163.367
R410 B.n334 B.n57 163.367
R411 B.n338 B.n57 163.367
R412 B.n460 B.n459 163.367
R413 B.n459 B.n458 163.367
R414 B.n458 B.n13 163.367
R415 B.n454 B.n13 163.367
R416 B.n454 B.n453 163.367
R417 B.n453 B.n452 163.367
R418 B.n452 B.n15 163.367
R419 B.n448 B.n15 163.367
R420 B.n448 B.n447 163.367
R421 B.n447 B.n446 163.367
R422 B.n446 B.n17 163.367
R423 B.n442 B.n17 163.367
R424 B.n442 B.n441 163.367
R425 B.n441 B.n440 163.367
R426 B.n440 B.n19 163.367
R427 B.n436 B.n19 163.367
R428 B.n436 B.n435 163.367
R429 B.n435 B.n434 163.367
R430 B.n434 B.n21 163.367
R431 B.n430 B.n21 163.367
R432 B.n430 B.n429 163.367
R433 B.n429 B.n428 163.367
R434 B.n428 B.n23 163.367
R435 B.n424 B.n23 163.367
R436 B.n424 B.n423 163.367
R437 B.n423 B.n422 163.367
R438 B.n422 B.n25 163.367
R439 B.n418 B.n25 163.367
R440 B.n418 B.n417 163.367
R441 B.n417 B.n416 163.367
R442 B.n416 B.n27 163.367
R443 B.n412 B.n27 163.367
R444 B.n412 B.n411 163.367
R445 B.n411 B.n410 163.367
R446 B.n410 B.n29 163.367
R447 B.n405 B.n29 163.367
R448 B.n405 B.n404 163.367
R449 B.n404 B.n403 163.367
R450 B.n403 B.n33 163.367
R451 B.n399 B.n33 163.367
R452 B.n399 B.n398 163.367
R453 B.n398 B.n397 163.367
R454 B.n397 B.n35 163.367
R455 B.n393 B.n35 163.367
R456 B.n393 B.n392 163.367
R457 B.n392 B.n39 163.367
R458 B.n388 B.n39 163.367
R459 B.n388 B.n387 163.367
R460 B.n387 B.n386 163.367
R461 B.n386 B.n41 163.367
R462 B.n382 B.n41 163.367
R463 B.n382 B.n381 163.367
R464 B.n381 B.n380 163.367
R465 B.n380 B.n43 163.367
R466 B.n376 B.n43 163.367
R467 B.n376 B.n375 163.367
R468 B.n375 B.n374 163.367
R469 B.n374 B.n45 163.367
R470 B.n370 B.n45 163.367
R471 B.n370 B.n369 163.367
R472 B.n369 B.n368 163.367
R473 B.n368 B.n47 163.367
R474 B.n364 B.n47 163.367
R475 B.n364 B.n363 163.367
R476 B.n363 B.n362 163.367
R477 B.n362 B.n49 163.367
R478 B.n358 B.n49 163.367
R479 B.n358 B.n357 163.367
R480 B.n357 B.n356 163.367
R481 B.n356 B.n51 163.367
R482 B.n352 B.n51 163.367
R483 B.n352 B.n351 163.367
R484 B.n351 B.n350 163.367
R485 B.n350 B.n53 163.367
R486 B.n346 B.n53 163.367
R487 B.n346 B.n345 163.367
R488 B.n345 B.n344 163.367
R489 B.n344 B.n55 163.367
R490 B.n340 B.n55 163.367
R491 B.n340 B.n339 163.367
R492 B.n96 B.n95 59.5399
R493 B.n211 B.n103 59.5399
R494 B.n407 B.n31 59.5399
R495 B.n38 B.n37 59.5399
R496 B.n95 B.n94 36.4611
R497 B.n103 B.n102 36.4611
R498 B.n31 B.n30 36.4611
R499 B.n37 B.n36 36.4611
R500 B.n462 B.n461 32.3127
R501 B.n337 B.n56 32.3127
R502 B.n281 B.n76 32.3127
R503 B.n157 B.n156 32.3127
R504 B B.n491 18.0485
R505 B.n461 B.n12 10.6151
R506 B.n457 B.n12 10.6151
R507 B.n457 B.n456 10.6151
R508 B.n456 B.n455 10.6151
R509 B.n455 B.n14 10.6151
R510 B.n451 B.n14 10.6151
R511 B.n451 B.n450 10.6151
R512 B.n450 B.n449 10.6151
R513 B.n449 B.n16 10.6151
R514 B.n445 B.n16 10.6151
R515 B.n445 B.n444 10.6151
R516 B.n444 B.n443 10.6151
R517 B.n443 B.n18 10.6151
R518 B.n439 B.n18 10.6151
R519 B.n439 B.n438 10.6151
R520 B.n438 B.n437 10.6151
R521 B.n437 B.n20 10.6151
R522 B.n433 B.n20 10.6151
R523 B.n433 B.n432 10.6151
R524 B.n432 B.n431 10.6151
R525 B.n431 B.n22 10.6151
R526 B.n427 B.n22 10.6151
R527 B.n427 B.n426 10.6151
R528 B.n426 B.n425 10.6151
R529 B.n425 B.n24 10.6151
R530 B.n421 B.n24 10.6151
R531 B.n421 B.n420 10.6151
R532 B.n420 B.n419 10.6151
R533 B.n419 B.n26 10.6151
R534 B.n415 B.n26 10.6151
R535 B.n415 B.n414 10.6151
R536 B.n414 B.n413 10.6151
R537 B.n413 B.n28 10.6151
R538 B.n409 B.n28 10.6151
R539 B.n409 B.n408 10.6151
R540 B.n406 B.n32 10.6151
R541 B.n402 B.n32 10.6151
R542 B.n402 B.n401 10.6151
R543 B.n401 B.n400 10.6151
R544 B.n400 B.n34 10.6151
R545 B.n396 B.n34 10.6151
R546 B.n396 B.n395 10.6151
R547 B.n395 B.n394 10.6151
R548 B.n391 B.n390 10.6151
R549 B.n390 B.n389 10.6151
R550 B.n389 B.n40 10.6151
R551 B.n385 B.n40 10.6151
R552 B.n385 B.n384 10.6151
R553 B.n384 B.n383 10.6151
R554 B.n383 B.n42 10.6151
R555 B.n379 B.n42 10.6151
R556 B.n379 B.n378 10.6151
R557 B.n378 B.n377 10.6151
R558 B.n377 B.n44 10.6151
R559 B.n373 B.n44 10.6151
R560 B.n373 B.n372 10.6151
R561 B.n372 B.n371 10.6151
R562 B.n371 B.n46 10.6151
R563 B.n367 B.n46 10.6151
R564 B.n367 B.n366 10.6151
R565 B.n366 B.n365 10.6151
R566 B.n365 B.n48 10.6151
R567 B.n361 B.n48 10.6151
R568 B.n361 B.n360 10.6151
R569 B.n360 B.n359 10.6151
R570 B.n359 B.n50 10.6151
R571 B.n355 B.n50 10.6151
R572 B.n355 B.n354 10.6151
R573 B.n354 B.n353 10.6151
R574 B.n353 B.n52 10.6151
R575 B.n349 B.n52 10.6151
R576 B.n349 B.n348 10.6151
R577 B.n348 B.n347 10.6151
R578 B.n347 B.n54 10.6151
R579 B.n343 B.n54 10.6151
R580 B.n343 B.n342 10.6151
R581 B.n342 B.n341 10.6151
R582 B.n341 B.n56 10.6151
R583 B.n282 B.n281 10.6151
R584 B.n283 B.n282 10.6151
R585 B.n283 B.n74 10.6151
R586 B.n287 B.n74 10.6151
R587 B.n288 B.n287 10.6151
R588 B.n289 B.n288 10.6151
R589 B.n289 B.n72 10.6151
R590 B.n293 B.n72 10.6151
R591 B.n294 B.n293 10.6151
R592 B.n295 B.n294 10.6151
R593 B.n295 B.n70 10.6151
R594 B.n299 B.n70 10.6151
R595 B.n300 B.n299 10.6151
R596 B.n301 B.n300 10.6151
R597 B.n301 B.n68 10.6151
R598 B.n305 B.n68 10.6151
R599 B.n306 B.n305 10.6151
R600 B.n307 B.n306 10.6151
R601 B.n307 B.n66 10.6151
R602 B.n311 B.n66 10.6151
R603 B.n312 B.n311 10.6151
R604 B.n313 B.n312 10.6151
R605 B.n313 B.n64 10.6151
R606 B.n317 B.n64 10.6151
R607 B.n318 B.n317 10.6151
R608 B.n319 B.n318 10.6151
R609 B.n319 B.n62 10.6151
R610 B.n323 B.n62 10.6151
R611 B.n324 B.n323 10.6151
R612 B.n325 B.n324 10.6151
R613 B.n325 B.n60 10.6151
R614 B.n329 B.n60 10.6151
R615 B.n330 B.n329 10.6151
R616 B.n331 B.n330 10.6151
R617 B.n331 B.n58 10.6151
R618 B.n335 B.n58 10.6151
R619 B.n336 B.n335 10.6151
R620 B.n337 B.n336 10.6151
R621 B.n157 B.n120 10.6151
R622 B.n161 B.n120 10.6151
R623 B.n162 B.n161 10.6151
R624 B.n163 B.n162 10.6151
R625 B.n163 B.n118 10.6151
R626 B.n167 B.n118 10.6151
R627 B.n168 B.n167 10.6151
R628 B.n169 B.n168 10.6151
R629 B.n169 B.n116 10.6151
R630 B.n173 B.n116 10.6151
R631 B.n174 B.n173 10.6151
R632 B.n175 B.n174 10.6151
R633 B.n175 B.n114 10.6151
R634 B.n179 B.n114 10.6151
R635 B.n180 B.n179 10.6151
R636 B.n181 B.n180 10.6151
R637 B.n181 B.n112 10.6151
R638 B.n185 B.n112 10.6151
R639 B.n186 B.n185 10.6151
R640 B.n187 B.n186 10.6151
R641 B.n187 B.n110 10.6151
R642 B.n191 B.n110 10.6151
R643 B.n192 B.n191 10.6151
R644 B.n193 B.n192 10.6151
R645 B.n193 B.n108 10.6151
R646 B.n197 B.n108 10.6151
R647 B.n198 B.n197 10.6151
R648 B.n199 B.n198 10.6151
R649 B.n199 B.n106 10.6151
R650 B.n203 B.n106 10.6151
R651 B.n204 B.n203 10.6151
R652 B.n205 B.n204 10.6151
R653 B.n205 B.n104 10.6151
R654 B.n209 B.n104 10.6151
R655 B.n210 B.n209 10.6151
R656 B.n212 B.n100 10.6151
R657 B.n216 B.n100 10.6151
R658 B.n217 B.n216 10.6151
R659 B.n218 B.n217 10.6151
R660 B.n218 B.n98 10.6151
R661 B.n222 B.n98 10.6151
R662 B.n223 B.n222 10.6151
R663 B.n224 B.n223 10.6151
R664 B.n228 B.n227 10.6151
R665 B.n229 B.n228 10.6151
R666 B.n229 B.n92 10.6151
R667 B.n233 B.n92 10.6151
R668 B.n234 B.n233 10.6151
R669 B.n235 B.n234 10.6151
R670 B.n235 B.n90 10.6151
R671 B.n239 B.n90 10.6151
R672 B.n240 B.n239 10.6151
R673 B.n241 B.n240 10.6151
R674 B.n241 B.n88 10.6151
R675 B.n245 B.n88 10.6151
R676 B.n246 B.n245 10.6151
R677 B.n247 B.n246 10.6151
R678 B.n247 B.n86 10.6151
R679 B.n251 B.n86 10.6151
R680 B.n252 B.n251 10.6151
R681 B.n253 B.n252 10.6151
R682 B.n253 B.n84 10.6151
R683 B.n257 B.n84 10.6151
R684 B.n258 B.n257 10.6151
R685 B.n259 B.n258 10.6151
R686 B.n259 B.n82 10.6151
R687 B.n263 B.n82 10.6151
R688 B.n264 B.n263 10.6151
R689 B.n265 B.n264 10.6151
R690 B.n265 B.n80 10.6151
R691 B.n269 B.n80 10.6151
R692 B.n270 B.n269 10.6151
R693 B.n271 B.n270 10.6151
R694 B.n271 B.n78 10.6151
R695 B.n275 B.n78 10.6151
R696 B.n276 B.n275 10.6151
R697 B.n277 B.n276 10.6151
R698 B.n277 B.n76 10.6151
R699 B.n156 B.n155 10.6151
R700 B.n155 B.n122 10.6151
R701 B.n151 B.n122 10.6151
R702 B.n151 B.n150 10.6151
R703 B.n150 B.n149 10.6151
R704 B.n149 B.n124 10.6151
R705 B.n145 B.n124 10.6151
R706 B.n145 B.n144 10.6151
R707 B.n144 B.n143 10.6151
R708 B.n143 B.n126 10.6151
R709 B.n139 B.n126 10.6151
R710 B.n139 B.n138 10.6151
R711 B.n138 B.n137 10.6151
R712 B.n137 B.n128 10.6151
R713 B.n133 B.n128 10.6151
R714 B.n133 B.n132 10.6151
R715 B.n132 B.n131 10.6151
R716 B.n131 B.n0 10.6151
R717 B.n487 B.n1 10.6151
R718 B.n487 B.n486 10.6151
R719 B.n486 B.n485 10.6151
R720 B.n485 B.n4 10.6151
R721 B.n481 B.n4 10.6151
R722 B.n481 B.n480 10.6151
R723 B.n480 B.n479 10.6151
R724 B.n479 B.n6 10.6151
R725 B.n475 B.n6 10.6151
R726 B.n475 B.n474 10.6151
R727 B.n474 B.n473 10.6151
R728 B.n473 B.n8 10.6151
R729 B.n469 B.n8 10.6151
R730 B.n469 B.n468 10.6151
R731 B.n468 B.n467 10.6151
R732 B.n467 B.n10 10.6151
R733 B.n463 B.n10 10.6151
R734 B.n463 B.n462 10.6151
R735 B.n407 B.n406 6.5566
R736 B.n394 B.n38 6.5566
R737 B.n212 B.n211 6.5566
R738 B.n224 B.n96 6.5566
R739 B.n408 B.n407 4.05904
R740 B.n391 B.n38 4.05904
R741 B.n211 B.n210 4.05904
R742 B.n227 B.n96 4.05904
R743 B.n491 B.n0 2.81026
R744 B.n491 B.n1 2.81026
R745 VP.n0 VP.t0 300.803
R746 VP.n0 VP.t1 260.498
R747 VP VP.n0 0.146778
R748 VTAIL.n210 VTAIL.n162 756.745
R749 VTAIL.n48 VTAIL.n0 756.745
R750 VTAIL.n156 VTAIL.n108 756.745
R751 VTAIL.n102 VTAIL.n54 756.745
R752 VTAIL.n178 VTAIL.n177 585
R753 VTAIL.n183 VTAIL.n182 585
R754 VTAIL.n185 VTAIL.n184 585
R755 VTAIL.n174 VTAIL.n173 585
R756 VTAIL.n191 VTAIL.n190 585
R757 VTAIL.n193 VTAIL.n192 585
R758 VTAIL.n170 VTAIL.n169 585
R759 VTAIL.n200 VTAIL.n199 585
R760 VTAIL.n201 VTAIL.n168 585
R761 VTAIL.n203 VTAIL.n202 585
R762 VTAIL.n166 VTAIL.n165 585
R763 VTAIL.n209 VTAIL.n208 585
R764 VTAIL.n211 VTAIL.n210 585
R765 VTAIL.n16 VTAIL.n15 585
R766 VTAIL.n21 VTAIL.n20 585
R767 VTAIL.n23 VTAIL.n22 585
R768 VTAIL.n12 VTAIL.n11 585
R769 VTAIL.n29 VTAIL.n28 585
R770 VTAIL.n31 VTAIL.n30 585
R771 VTAIL.n8 VTAIL.n7 585
R772 VTAIL.n38 VTAIL.n37 585
R773 VTAIL.n39 VTAIL.n6 585
R774 VTAIL.n41 VTAIL.n40 585
R775 VTAIL.n4 VTAIL.n3 585
R776 VTAIL.n47 VTAIL.n46 585
R777 VTAIL.n49 VTAIL.n48 585
R778 VTAIL.n157 VTAIL.n156 585
R779 VTAIL.n155 VTAIL.n154 585
R780 VTAIL.n112 VTAIL.n111 585
R781 VTAIL.n149 VTAIL.n148 585
R782 VTAIL.n147 VTAIL.n114 585
R783 VTAIL.n146 VTAIL.n145 585
R784 VTAIL.n117 VTAIL.n115 585
R785 VTAIL.n140 VTAIL.n139 585
R786 VTAIL.n138 VTAIL.n137 585
R787 VTAIL.n121 VTAIL.n120 585
R788 VTAIL.n132 VTAIL.n131 585
R789 VTAIL.n130 VTAIL.n129 585
R790 VTAIL.n125 VTAIL.n124 585
R791 VTAIL.n103 VTAIL.n102 585
R792 VTAIL.n101 VTAIL.n100 585
R793 VTAIL.n58 VTAIL.n57 585
R794 VTAIL.n95 VTAIL.n94 585
R795 VTAIL.n93 VTAIL.n60 585
R796 VTAIL.n92 VTAIL.n91 585
R797 VTAIL.n63 VTAIL.n61 585
R798 VTAIL.n86 VTAIL.n85 585
R799 VTAIL.n84 VTAIL.n83 585
R800 VTAIL.n67 VTAIL.n66 585
R801 VTAIL.n78 VTAIL.n77 585
R802 VTAIL.n76 VTAIL.n75 585
R803 VTAIL.n71 VTAIL.n70 585
R804 VTAIL.n179 VTAIL.t0 329.038
R805 VTAIL.n17 VTAIL.t3 329.038
R806 VTAIL.n126 VTAIL.t2 329.038
R807 VTAIL.n72 VTAIL.t1 329.038
R808 VTAIL.n183 VTAIL.n177 171.744
R809 VTAIL.n184 VTAIL.n183 171.744
R810 VTAIL.n184 VTAIL.n173 171.744
R811 VTAIL.n191 VTAIL.n173 171.744
R812 VTAIL.n192 VTAIL.n191 171.744
R813 VTAIL.n192 VTAIL.n169 171.744
R814 VTAIL.n200 VTAIL.n169 171.744
R815 VTAIL.n201 VTAIL.n200 171.744
R816 VTAIL.n202 VTAIL.n201 171.744
R817 VTAIL.n202 VTAIL.n165 171.744
R818 VTAIL.n209 VTAIL.n165 171.744
R819 VTAIL.n210 VTAIL.n209 171.744
R820 VTAIL.n21 VTAIL.n15 171.744
R821 VTAIL.n22 VTAIL.n21 171.744
R822 VTAIL.n22 VTAIL.n11 171.744
R823 VTAIL.n29 VTAIL.n11 171.744
R824 VTAIL.n30 VTAIL.n29 171.744
R825 VTAIL.n30 VTAIL.n7 171.744
R826 VTAIL.n38 VTAIL.n7 171.744
R827 VTAIL.n39 VTAIL.n38 171.744
R828 VTAIL.n40 VTAIL.n39 171.744
R829 VTAIL.n40 VTAIL.n3 171.744
R830 VTAIL.n47 VTAIL.n3 171.744
R831 VTAIL.n48 VTAIL.n47 171.744
R832 VTAIL.n156 VTAIL.n155 171.744
R833 VTAIL.n155 VTAIL.n111 171.744
R834 VTAIL.n148 VTAIL.n111 171.744
R835 VTAIL.n148 VTAIL.n147 171.744
R836 VTAIL.n147 VTAIL.n146 171.744
R837 VTAIL.n146 VTAIL.n115 171.744
R838 VTAIL.n139 VTAIL.n115 171.744
R839 VTAIL.n139 VTAIL.n138 171.744
R840 VTAIL.n138 VTAIL.n120 171.744
R841 VTAIL.n131 VTAIL.n120 171.744
R842 VTAIL.n131 VTAIL.n130 171.744
R843 VTAIL.n130 VTAIL.n124 171.744
R844 VTAIL.n102 VTAIL.n101 171.744
R845 VTAIL.n101 VTAIL.n57 171.744
R846 VTAIL.n94 VTAIL.n57 171.744
R847 VTAIL.n94 VTAIL.n93 171.744
R848 VTAIL.n93 VTAIL.n92 171.744
R849 VTAIL.n92 VTAIL.n61 171.744
R850 VTAIL.n85 VTAIL.n61 171.744
R851 VTAIL.n85 VTAIL.n84 171.744
R852 VTAIL.n84 VTAIL.n66 171.744
R853 VTAIL.n77 VTAIL.n66 171.744
R854 VTAIL.n77 VTAIL.n76 171.744
R855 VTAIL.n76 VTAIL.n70 171.744
R856 VTAIL.t0 VTAIL.n177 85.8723
R857 VTAIL.t3 VTAIL.n15 85.8723
R858 VTAIL.t2 VTAIL.n124 85.8723
R859 VTAIL.t1 VTAIL.n70 85.8723
R860 VTAIL.n215 VTAIL.n214 31.6035
R861 VTAIL.n53 VTAIL.n52 31.6035
R862 VTAIL.n161 VTAIL.n160 31.6035
R863 VTAIL.n107 VTAIL.n106 31.6035
R864 VTAIL.n107 VTAIL.n53 24.1686
R865 VTAIL.n215 VTAIL.n161 22.5479
R866 VTAIL.n203 VTAIL.n168 13.1884
R867 VTAIL.n41 VTAIL.n6 13.1884
R868 VTAIL.n149 VTAIL.n114 13.1884
R869 VTAIL.n95 VTAIL.n60 13.1884
R870 VTAIL.n199 VTAIL.n198 12.8005
R871 VTAIL.n204 VTAIL.n166 12.8005
R872 VTAIL.n37 VTAIL.n36 12.8005
R873 VTAIL.n42 VTAIL.n4 12.8005
R874 VTAIL.n150 VTAIL.n112 12.8005
R875 VTAIL.n145 VTAIL.n116 12.8005
R876 VTAIL.n96 VTAIL.n58 12.8005
R877 VTAIL.n91 VTAIL.n62 12.8005
R878 VTAIL.n197 VTAIL.n170 12.0247
R879 VTAIL.n208 VTAIL.n207 12.0247
R880 VTAIL.n35 VTAIL.n8 12.0247
R881 VTAIL.n46 VTAIL.n45 12.0247
R882 VTAIL.n154 VTAIL.n153 12.0247
R883 VTAIL.n144 VTAIL.n117 12.0247
R884 VTAIL.n100 VTAIL.n99 12.0247
R885 VTAIL.n90 VTAIL.n63 12.0247
R886 VTAIL.n194 VTAIL.n193 11.249
R887 VTAIL.n211 VTAIL.n164 11.249
R888 VTAIL.n32 VTAIL.n31 11.249
R889 VTAIL.n49 VTAIL.n2 11.249
R890 VTAIL.n157 VTAIL.n110 11.249
R891 VTAIL.n141 VTAIL.n140 11.249
R892 VTAIL.n103 VTAIL.n56 11.249
R893 VTAIL.n87 VTAIL.n86 11.249
R894 VTAIL.n179 VTAIL.n178 10.7239
R895 VTAIL.n17 VTAIL.n16 10.7239
R896 VTAIL.n126 VTAIL.n125 10.7239
R897 VTAIL.n72 VTAIL.n71 10.7239
R898 VTAIL.n190 VTAIL.n172 10.4732
R899 VTAIL.n212 VTAIL.n162 10.4732
R900 VTAIL.n28 VTAIL.n10 10.4732
R901 VTAIL.n50 VTAIL.n0 10.4732
R902 VTAIL.n158 VTAIL.n108 10.4732
R903 VTAIL.n137 VTAIL.n119 10.4732
R904 VTAIL.n104 VTAIL.n54 10.4732
R905 VTAIL.n83 VTAIL.n65 10.4732
R906 VTAIL.n189 VTAIL.n174 9.69747
R907 VTAIL.n27 VTAIL.n12 9.69747
R908 VTAIL.n136 VTAIL.n121 9.69747
R909 VTAIL.n82 VTAIL.n67 9.69747
R910 VTAIL.n214 VTAIL.n213 9.45567
R911 VTAIL.n52 VTAIL.n51 9.45567
R912 VTAIL.n160 VTAIL.n159 9.45567
R913 VTAIL.n106 VTAIL.n105 9.45567
R914 VTAIL.n213 VTAIL.n212 9.3005
R915 VTAIL.n164 VTAIL.n163 9.3005
R916 VTAIL.n207 VTAIL.n206 9.3005
R917 VTAIL.n205 VTAIL.n204 9.3005
R918 VTAIL.n181 VTAIL.n180 9.3005
R919 VTAIL.n176 VTAIL.n175 9.3005
R920 VTAIL.n187 VTAIL.n186 9.3005
R921 VTAIL.n189 VTAIL.n188 9.3005
R922 VTAIL.n172 VTAIL.n171 9.3005
R923 VTAIL.n195 VTAIL.n194 9.3005
R924 VTAIL.n197 VTAIL.n196 9.3005
R925 VTAIL.n198 VTAIL.n167 9.3005
R926 VTAIL.n51 VTAIL.n50 9.3005
R927 VTAIL.n2 VTAIL.n1 9.3005
R928 VTAIL.n45 VTAIL.n44 9.3005
R929 VTAIL.n43 VTAIL.n42 9.3005
R930 VTAIL.n19 VTAIL.n18 9.3005
R931 VTAIL.n14 VTAIL.n13 9.3005
R932 VTAIL.n25 VTAIL.n24 9.3005
R933 VTAIL.n27 VTAIL.n26 9.3005
R934 VTAIL.n10 VTAIL.n9 9.3005
R935 VTAIL.n33 VTAIL.n32 9.3005
R936 VTAIL.n35 VTAIL.n34 9.3005
R937 VTAIL.n36 VTAIL.n5 9.3005
R938 VTAIL.n128 VTAIL.n127 9.3005
R939 VTAIL.n123 VTAIL.n122 9.3005
R940 VTAIL.n134 VTAIL.n133 9.3005
R941 VTAIL.n136 VTAIL.n135 9.3005
R942 VTAIL.n119 VTAIL.n118 9.3005
R943 VTAIL.n142 VTAIL.n141 9.3005
R944 VTAIL.n144 VTAIL.n143 9.3005
R945 VTAIL.n116 VTAIL.n113 9.3005
R946 VTAIL.n159 VTAIL.n158 9.3005
R947 VTAIL.n110 VTAIL.n109 9.3005
R948 VTAIL.n153 VTAIL.n152 9.3005
R949 VTAIL.n151 VTAIL.n150 9.3005
R950 VTAIL.n74 VTAIL.n73 9.3005
R951 VTAIL.n69 VTAIL.n68 9.3005
R952 VTAIL.n80 VTAIL.n79 9.3005
R953 VTAIL.n82 VTAIL.n81 9.3005
R954 VTAIL.n65 VTAIL.n64 9.3005
R955 VTAIL.n88 VTAIL.n87 9.3005
R956 VTAIL.n90 VTAIL.n89 9.3005
R957 VTAIL.n62 VTAIL.n59 9.3005
R958 VTAIL.n105 VTAIL.n104 9.3005
R959 VTAIL.n56 VTAIL.n55 9.3005
R960 VTAIL.n99 VTAIL.n98 9.3005
R961 VTAIL.n97 VTAIL.n96 9.3005
R962 VTAIL.n186 VTAIL.n185 8.92171
R963 VTAIL.n24 VTAIL.n23 8.92171
R964 VTAIL.n133 VTAIL.n132 8.92171
R965 VTAIL.n79 VTAIL.n78 8.92171
R966 VTAIL.n182 VTAIL.n176 8.14595
R967 VTAIL.n20 VTAIL.n14 8.14595
R968 VTAIL.n129 VTAIL.n123 8.14595
R969 VTAIL.n75 VTAIL.n69 8.14595
R970 VTAIL.n181 VTAIL.n178 7.3702
R971 VTAIL.n19 VTAIL.n16 7.3702
R972 VTAIL.n128 VTAIL.n125 7.3702
R973 VTAIL.n74 VTAIL.n71 7.3702
R974 VTAIL.n182 VTAIL.n181 5.81868
R975 VTAIL.n20 VTAIL.n19 5.81868
R976 VTAIL.n129 VTAIL.n128 5.81868
R977 VTAIL.n75 VTAIL.n74 5.81868
R978 VTAIL.n185 VTAIL.n176 5.04292
R979 VTAIL.n23 VTAIL.n14 5.04292
R980 VTAIL.n132 VTAIL.n123 5.04292
R981 VTAIL.n78 VTAIL.n69 5.04292
R982 VTAIL.n186 VTAIL.n174 4.26717
R983 VTAIL.n24 VTAIL.n12 4.26717
R984 VTAIL.n133 VTAIL.n121 4.26717
R985 VTAIL.n79 VTAIL.n67 4.26717
R986 VTAIL.n190 VTAIL.n189 3.49141
R987 VTAIL.n214 VTAIL.n162 3.49141
R988 VTAIL.n28 VTAIL.n27 3.49141
R989 VTAIL.n52 VTAIL.n0 3.49141
R990 VTAIL.n160 VTAIL.n108 3.49141
R991 VTAIL.n137 VTAIL.n136 3.49141
R992 VTAIL.n106 VTAIL.n54 3.49141
R993 VTAIL.n83 VTAIL.n82 3.49141
R994 VTAIL.n193 VTAIL.n172 2.71565
R995 VTAIL.n212 VTAIL.n211 2.71565
R996 VTAIL.n31 VTAIL.n10 2.71565
R997 VTAIL.n50 VTAIL.n49 2.71565
R998 VTAIL.n158 VTAIL.n157 2.71565
R999 VTAIL.n140 VTAIL.n119 2.71565
R1000 VTAIL.n104 VTAIL.n103 2.71565
R1001 VTAIL.n86 VTAIL.n65 2.71565
R1002 VTAIL.n180 VTAIL.n179 2.41283
R1003 VTAIL.n18 VTAIL.n17 2.41283
R1004 VTAIL.n127 VTAIL.n126 2.41283
R1005 VTAIL.n73 VTAIL.n72 2.41283
R1006 VTAIL.n194 VTAIL.n170 1.93989
R1007 VTAIL.n208 VTAIL.n164 1.93989
R1008 VTAIL.n32 VTAIL.n8 1.93989
R1009 VTAIL.n46 VTAIL.n2 1.93989
R1010 VTAIL.n154 VTAIL.n110 1.93989
R1011 VTAIL.n141 VTAIL.n117 1.93989
R1012 VTAIL.n100 VTAIL.n56 1.93989
R1013 VTAIL.n87 VTAIL.n63 1.93989
R1014 VTAIL.n161 VTAIL.n107 1.28067
R1015 VTAIL.n199 VTAIL.n197 1.16414
R1016 VTAIL.n207 VTAIL.n166 1.16414
R1017 VTAIL.n37 VTAIL.n35 1.16414
R1018 VTAIL.n45 VTAIL.n4 1.16414
R1019 VTAIL.n153 VTAIL.n112 1.16414
R1020 VTAIL.n145 VTAIL.n144 1.16414
R1021 VTAIL.n99 VTAIL.n58 1.16414
R1022 VTAIL.n91 VTAIL.n90 1.16414
R1023 VTAIL VTAIL.n53 0.93369
R1024 VTAIL.n198 VTAIL.n168 0.388379
R1025 VTAIL.n204 VTAIL.n203 0.388379
R1026 VTAIL.n36 VTAIL.n6 0.388379
R1027 VTAIL.n42 VTAIL.n41 0.388379
R1028 VTAIL.n150 VTAIL.n149 0.388379
R1029 VTAIL.n116 VTAIL.n114 0.388379
R1030 VTAIL.n96 VTAIL.n95 0.388379
R1031 VTAIL.n62 VTAIL.n60 0.388379
R1032 VTAIL VTAIL.n215 0.347483
R1033 VTAIL.n180 VTAIL.n175 0.155672
R1034 VTAIL.n187 VTAIL.n175 0.155672
R1035 VTAIL.n188 VTAIL.n187 0.155672
R1036 VTAIL.n188 VTAIL.n171 0.155672
R1037 VTAIL.n195 VTAIL.n171 0.155672
R1038 VTAIL.n196 VTAIL.n195 0.155672
R1039 VTAIL.n196 VTAIL.n167 0.155672
R1040 VTAIL.n205 VTAIL.n167 0.155672
R1041 VTAIL.n206 VTAIL.n205 0.155672
R1042 VTAIL.n206 VTAIL.n163 0.155672
R1043 VTAIL.n213 VTAIL.n163 0.155672
R1044 VTAIL.n18 VTAIL.n13 0.155672
R1045 VTAIL.n25 VTAIL.n13 0.155672
R1046 VTAIL.n26 VTAIL.n25 0.155672
R1047 VTAIL.n26 VTAIL.n9 0.155672
R1048 VTAIL.n33 VTAIL.n9 0.155672
R1049 VTAIL.n34 VTAIL.n33 0.155672
R1050 VTAIL.n34 VTAIL.n5 0.155672
R1051 VTAIL.n43 VTAIL.n5 0.155672
R1052 VTAIL.n44 VTAIL.n43 0.155672
R1053 VTAIL.n44 VTAIL.n1 0.155672
R1054 VTAIL.n51 VTAIL.n1 0.155672
R1055 VTAIL.n159 VTAIL.n109 0.155672
R1056 VTAIL.n152 VTAIL.n109 0.155672
R1057 VTAIL.n152 VTAIL.n151 0.155672
R1058 VTAIL.n151 VTAIL.n113 0.155672
R1059 VTAIL.n143 VTAIL.n113 0.155672
R1060 VTAIL.n143 VTAIL.n142 0.155672
R1061 VTAIL.n142 VTAIL.n118 0.155672
R1062 VTAIL.n135 VTAIL.n118 0.155672
R1063 VTAIL.n135 VTAIL.n134 0.155672
R1064 VTAIL.n134 VTAIL.n122 0.155672
R1065 VTAIL.n127 VTAIL.n122 0.155672
R1066 VTAIL.n105 VTAIL.n55 0.155672
R1067 VTAIL.n98 VTAIL.n55 0.155672
R1068 VTAIL.n98 VTAIL.n97 0.155672
R1069 VTAIL.n97 VTAIL.n59 0.155672
R1070 VTAIL.n89 VTAIL.n59 0.155672
R1071 VTAIL.n89 VTAIL.n88 0.155672
R1072 VTAIL.n88 VTAIL.n64 0.155672
R1073 VTAIL.n81 VTAIL.n64 0.155672
R1074 VTAIL.n81 VTAIL.n80 0.155672
R1075 VTAIL.n80 VTAIL.n68 0.155672
R1076 VTAIL.n73 VTAIL.n68 0.155672
R1077 VDD1.n48 VDD1.n0 756.745
R1078 VDD1.n101 VDD1.n53 756.745
R1079 VDD1.n49 VDD1.n48 585
R1080 VDD1.n47 VDD1.n46 585
R1081 VDD1.n4 VDD1.n3 585
R1082 VDD1.n41 VDD1.n40 585
R1083 VDD1.n39 VDD1.n6 585
R1084 VDD1.n38 VDD1.n37 585
R1085 VDD1.n9 VDD1.n7 585
R1086 VDD1.n32 VDD1.n31 585
R1087 VDD1.n30 VDD1.n29 585
R1088 VDD1.n13 VDD1.n12 585
R1089 VDD1.n24 VDD1.n23 585
R1090 VDD1.n22 VDD1.n21 585
R1091 VDD1.n17 VDD1.n16 585
R1092 VDD1.n69 VDD1.n68 585
R1093 VDD1.n74 VDD1.n73 585
R1094 VDD1.n76 VDD1.n75 585
R1095 VDD1.n65 VDD1.n64 585
R1096 VDD1.n82 VDD1.n81 585
R1097 VDD1.n84 VDD1.n83 585
R1098 VDD1.n61 VDD1.n60 585
R1099 VDD1.n91 VDD1.n90 585
R1100 VDD1.n92 VDD1.n59 585
R1101 VDD1.n94 VDD1.n93 585
R1102 VDD1.n57 VDD1.n56 585
R1103 VDD1.n100 VDD1.n99 585
R1104 VDD1.n102 VDD1.n101 585
R1105 VDD1.n70 VDD1.t0 329.038
R1106 VDD1.n18 VDD1.t1 329.038
R1107 VDD1.n48 VDD1.n47 171.744
R1108 VDD1.n47 VDD1.n3 171.744
R1109 VDD1.n40 VDD1.n3 171.744
R1110 VDD1.n40 VDD1.n39 171.744
R1111 VDD1.n39 VDD1.n38 171.744
R1112 VDD1.n38 VDD1.n7 171.744
R1113 VDD1.n31 VDD1.n7 171.744
R1114 VDD1.n31 VDD1.n30 171.744
R1115 VDD1.n30 VDD1.n12 171.744
R1116 VDD1.n23 VDD1.n12 171.744
R1117 VDD1.n23 VDD1.n22 171.744
R1118 VDD1.n22 VDD1.n16 171.744
R1119 VDD1.n74 VDD1.n68 171.744
R1120 VDD1.n75 VDD1.n74 171.744
R1121 VDD1.n75 VDD1.n64 171.744
R1122 VDD1.n82 VDD1.n64 171.744
R1123 VDD1.n83 VDD1.n82 171.744
R1124 VDD1.n83 VDD1.n60 171.744
R1125 VDD1.n91 VDD1.n60 171.744
R1126 VDD1.n92 VDD1.n91 171.744
R1127 VDD1.n93 VDD1.n92 171.744
R1128 VDD1.n93 VDD1.n56 171.744
R1129 VDD1.n100 VDD1.n56 171.744
R1130 VDD1.n101 VDD1.n100 171.744
R1131 VDD1.t1 VDD1.n16 85.8723
R1132 VDD1.t0 VDD1.n68 85.8723
R1133 VDD1 VDD1.n105 84.6735
R1134 VDD1 VDD1.n52 48.7457
R1135 VDD1.n41 VDD1.n6 13.1884
R1136 VDD1.n94 VDD1.n59 13.1884
R1137 VDD1.n42 VDD1.n4 12.8005
R1138 VDD1.n37 VDD1.n8 12.8005
R1139 VDD1.n90 VDD1.n89 12.8005
R1140 VDD1.n95 VDD1.n57 12.8005
R1141 VDD1.n46 VDD1.n45 12.0247
R1142 VDD1.n36 VDD1.n9 12.0247
R1143 VDD1.n88 VDD1.n61 12.0247
R1144 VDD1.n99 VDD1.n98 12.0247
R1145 VDD1.n49 VDD1.n2 11.249
R1146 VDD1.n33 VDD1.n32 11.249
R1147 VDD1.n85 VDD1.n84 11.249
R1148 VDD1.n102 VDD1.n55 11.249
R1149 VDD1.n18 VDD1.n17 10.7239
R1150 VDD1.n70 VDD1.n69 10.7239
R1151 VDD1.n50 VDD1.n0 10.4732
R1152 VDD1.n29 VDD1.n11 10.4732
R1153 VDD1.n81 VDD1.n63 10.4732
R1154 VDD1.n103 VDD1.n53 10.4732
R1155 VDD1.n28 VDD1.n13 9.69747
R1156 VDD1.n80 VDD1.n65 9.69747
R1157 VDD1.n52 VDD1.n51 9.45567
R1158 VDD1.n105 VDD1.n104 9.45567
R1159 VDD1.n20 VDD1.n19 9.3005
R1160 VDD1.n15 VDD1.n14 9.3005
R1161 VDD1.n26 VDD1.n25 9.3005
R1162 VDD1.n28 VDD1.n27 9.3005
R1163 VDD1.n11 VDD1.n10 9.3005
R1164 VDD1.n34 VDD1.n33 9.3005
R1165 VDD1.n36 VDD1.n35 9.3005
R1166 VDD1.n8 VDD1.n5 9.3005
R1167 VDD1.n51 VDD1.n50 9.3005
R1168 VDD1.n2 VDD1.n1 9.3005
R1169 VDD1.n45 VDD1.n44 9.3005
R1170 VDD1.n43 VDD1.n42 9.3005
R1171 VDD1.n104 VDD1.n103 9.3005
R1172 VDD1.n55 VDD1.n54 9.3005
R1173 VDD1.n98 VDD1.n97 9.3005
R1174 VDD1.n96 VDD1.n95 9.3005
R1175 VDD1.n72 VDD1.n71 9.3005
R1176 VDD1.n67 VDD1.n66 9.3005
R1177 VDD1.n78 VDD1.n77 9.3005
R1178 VDD1.n80 VDD1.n79 9.3005
R1179 VDD1.n63 VDD1.n62 9.3005
R1180 VDD1.n86 VDD1.n85 9.3005
R1181 VDD1.n88 VDD1.n87 9.3005
R1182 VDD1.n89 VDD1.n58 9.3005
R1183 VDD1.n25 VDD1.n24 8.92171
R1184 VDD1.n77 VDD1.n76 8.92171
R1185 VDD1.n21 VDD1.n15 8.14595
R1186 VDD1.n73 VDD1.n67 8.14595
R1187 VDD1.n20 VDD1.n17 7.3702
R1188 VDD1.n72 VDD1.n69 7.3702
R1189 VDD1.n21 VDD1.n20 5.81868
R1190 VDD1.n73 VDD1.n72 5.81868
R1191 VDD1.n24 VDD1.n15 5.04292
R1192 VDD1.n76 VDD1.n67 5.04292
R1193 VDD1.n25 VDD1.n13 4.26717
R1194 VDD1.n77 VDD1.n65 4.26717
R1195 VDD1.n52 VDD1.n0 3.49141
R1196 VDD1.n29 VDD1.n28 3.49141
R1197 VDD1.n81 VDD1.n80 3.49141
R1198 VDD1.n105 VDD1.n53 3.49141
R1199 VDD1.n50 VDD1.n49 2.71565
R1200 VDD1.n32 VDD1.n11 2.71565
R1201 VDD1.n84 VDD1.n63 2.71565
R1202 VDD1.n103 VDD1.n102 2.71565
R1203 VDD1.n19 VDD1.n18 2.41283
R1204 VDD1.n71 VDD1.n70 2.41283
R1205 VDD1.n46 VDD1.n2 1.93989
R1206 VDD1.n33 VDD1.n9 1.93989
R1207 VDD1.n85 VDD1.n61 1.93989
R1208 VDD1.n99 VDD1.n55 1.93989
R1209 VDD1.n45 VDD1.n4 1.16414
R1210 VDD1.n37 VDD1.n36 1.16414
R1211 VDD1.n90 VDD1.n88 1.16414
R1212 VDD1.n98 VDD1.n57 1.16414
R1213 VDD1.n42 VDD1.n41 0.388379
R1214 VDD1.n8 VDD1.n6 0.388379
R1215 VDD1.n89 VDD1.n59 0.388379
R1216 VDD1.n95 VDD1.n94 0.388379
R1217 VDD1.n51 VDD1.n1 0.155672
R1218 VDD1.n44 VDD1.n1 0.155672
R1219 VDD1.n44 VDD1.n43 0.155672
R1220 VDD1.n43 VDD1.n5 0.155672
R1221 VDD1.n35 VDD1.n5 0.155672
R1222 VDD1.n35 VDD1.n34 0.155672
R1223 VDD1.n34 VDD1.n10 0.155672
R1224 VDD1.n27 VDD1.n10 0.155672
R1225 VDD1.n27 VDD1.n26 0.155672
R1226 VDD1.n26 VDD1.n14 0.155672
R1227 VDD1.n19 VDD1.n14 0.155672
R1228 VDD1.n71 VDD1.n66 0.155672
R1229 VDD1.n78 VDD1.n66 0.155672
R1230 VDD1.n79 VDD1.n78 0.155672
R1231 VDD1.n79 VDD1.n62 0.155672
R1232 VDD1.n86 VDD1.n62 0.155672
R1233 VDD1.n87 VDD1.n86 0.155672
R1234 VDD1.n87 VDD1.n58 0.155672
R1235 VDD1.n96 VDD1.n58 0.155672
R1236 VDD1.n97 VDD1.n96 0.155672
R1237 VDD1.n97 VDD1.n54 0.155672
R1238 VDD1.n104 VDD1.n54 0.155672
R1239 VN VN.t0 301.087
R1240 VN VN.t1 260.644
R1241 VDD2.n101 VDD2.n53 756.745
R1242 VDD2.n48 VDD2.n0 756.745
R1243 VDD2.n102 VDD2.n101 585
R1244 VDD2.n100 VDD2.n99 585
R1245 VDD2.n57 VDD2.n56 585
R1246 VDD2.n94 VDD2.n93 585
R1247 VDD2.n92 VDD2.n59 585
R1248 VDD2.n91 VDD2.n90 585
R1249 VDD2.n62 VDD2.n60 585
R1250 VDD2.n85 VDD2.n84 585
R1251 VDD2.n83 VDD2.n82 585
R1252 VDD2.n66 VDD2.n65 585
R1253 VDD2.n77 VDD2.n76 585
R1254 VDD2.n75 VDD2.n74 585
R1255 VDD2.n70 VDD2.n69 585
R1256 VDD2.n16 VDD2.n15 585
R1257 VDD2.n21 VDD2.n20 585
R1258 VDD2.n23 VDD2.n22 585
R1259 VDD2.n12 VDD2.n11 585
R1260 VDD2.n29 VDD2.n28 585
R1261 VDD2.n31 VDD2.n30 585
R1262 VDD2.n8 VDD2.n7 585
R1263 VDD2.n38 VDD2.n37 585
R1264 VDD2.n39 VDD2.n6 585
R1265 VDD2.n41 VDD2.n40 585
R1266 VDD2.n4 VDD2.n3 585
R1267 VDD2.n47 VDD2.n46 585
R1268 VDD2.n49 VDD2.n48 585
R1269 VDD2.n17 VDD2.t0 329.038
R1270 VDD2.n71 VDD2.t1 329.038
R1271 VDD2.n101 VDD2.n100 171.744
R1272 VDD2.n100 VDD2.n56 171.744
R1273 VDD2.n93 VDD2.n56 171.744
R1274 VDD2.n93 VDD2.n92 171.744
R1275 VDD2.n92 VDD2.n91 171.744
R1276 VDD2.n91 VDD2.n60 171.744
R1277 VDD2.n84 VDD2.n60 171.744
R1278 VDD2.n84 VDD2.n83 171.744
R1279 VDD2.n83 VDD2.n65 171.744
R1280 VDD2.n76 VDD2.n65 171.744
R1281 VDD2.n76 VDD2.n75 171.744
R1282 VDD2.n75 VDD2.n69 171.744
R1283 VDD2.n21 VDD2.n15 171.744
R1284 VDD2.n22 VDD2.n21 171.744
R1285 VDD2.n22 VDD2.n11 171.744
R1286 VDD2.n29 VDD2.n11 171.744
R1287 VDD2.n30 VDD2.n29 171.744
R1288 VDD2.n30 VDD2.n7 171.744
R1289 VDD2.n38 VDD2.n7 171.744
R1290 VDD2.n39 VDD2.n38 171.744
R1291 VDD2.n40 VDD2.n39 171.744
R1292 VDD2.n40 VDD2.n3 171.744
R1293 VDD2.n47 VDD2.n3 171.744
R1294 VDD2.n48 VDD2.n47 171.744
R1295 VDD2.t1 VDD2.n69 85.8723
R1296 VDD2.t0 VDD2.n15 85.8723
R1297 VDD2.n106 VDD2.n52 83.7435
R1298 VDD2.n106 VDD2.n105 48.2823
R1299 VDD2.n94 VDD2.n59 13.1884
R1300 VDD2.n41 VDD2.n6 13.1884
R1301 VDD2.n95 VDD2.n57 12.8005
R1302 VDD2.n90 VDD2.n61 12.8005
R1303 VDD2.n37 VDD2.n36 12.8005
R1304 VDD2.n42 VDD2.n4 12.8005
R1305 VDD2.n99 VDD2.n98 12.0247
R1306 VDD2.n89 VDD2.n62 12.0247
R1307 VDD2.n35 VDD2.n8 12.0247
R1308 VDD2.n46 VDD2.n45 12.0247
R1309 VDD2.n102 VDD2.n55 11.249
R1310 VDD2.n86 VDD2.n85 11.249
R1311 VDD2.n32 VDD2.n31 11.249
R1312 VDD2.n49 VDD2.n2 11.249
R1313 VDD2.n71 VDD2.n70 10.7239
R1314 VDD2.n17 VDD2.n16 10.7239
R1315 VDD2.n103 VDD2.n53 10.4732
R1316 VDD2.n82 VDD2.n64 10.4732
R1317 VDD2.n28 VDD2.n10 10.4732
R1318 VDD2.n50 VDD2.n0 10.4732
R1319 VDD2.n81 VDD2.n66 9.69747
R1320 VDD2.n27 VDD2.n12 9.69747
R1321 VDD2.n105 VDD2.n104 9.45567
R1322 VDD2.n52 VDD2.n51 9.45567
R1323 VDD2.n73 VDD2.n72 9.3005
R1324 VDD2.n68 VDD2.n67 9.3005
R1325 VDD2.n79 VDD2.n78 9.3005
R1326 VDD2.n81 VDD2.n80 9.3005
R1327 VDD2.n64 VDD2.n63 9.3005
R1328 VDD2.n87 VDD2.n86 9.3005
R1329 VDD2.n89 VDD2.n88 9.3005
R1330 VDD2.n61 VDD2.n58 9.3005
R1331 VDD2.n104 VDD2.n103 9.3005
R1332 VDD2.n55 VDD2.n54 9.3005
R1333 VDD2.n98 VDD2.n97 9.3005
R1334 VDD2.n96 VDD2.n95 9.3005
R1335 VDD2.n51 VDD2.n50 9.3005
R1336 VDD2.n2 VDD2.n1 9.3005
R1337 VDD2.n45 VDD2.n44 9.3005
R1338 VDD2.n43 VDD2.n42 9.3005
R1339 VDD2.n19 VDD2.n18 9.3005
R1340 VDD2.n14 VDD2.n13 9.3005
R1341 VDD2.n25 VDD2.n24 9.3005
R1342 VDD2.n27 VDD2.n26 9.3005
R1343 VDD2.n10 VDD2.n9 9.3005
R1344 VDD2.n33 VDD2.n32 9.3005
R1345 VDD2.n35 VDD2.n34 9.3005
R1346 VDD2.n36 VDD2.n5 9.3005
R1347 VDD2.n78 VDD2.n77 8.92171
R1348 VDD2.n24 VDD2.n23 8.92171
R1349 VDD2.n74 VDD2.n68 8.14595
R1350 VDD2.n20 VDD2.n14 8.14595
R1351 VDD2.n73 VDD2.n70 7.3702
R1352 VDD2.n19 VDD2.n16 7.3702
R1353 VDD2.n74 VDD2.n73 5.81868
R1354 VDD2.n20 VDD2.n19 5.81868
R1355 VDD2.n77 VDD2.n68 5.04292
R1356 VDD2.n23 VDD2.n14 5.04292
R1357 VDD2.n78 VDD2.n66 4.26717
R1358 VDD2.n24 VDD2.n12 4.26717
R1359 VDD2.n105 VDD2.n53 3.49141
R1360 VDD2.n82 VDD2.n81 3.49141
R1361 VDD2.n28 VDD2.n27 3.49141
R1362 VDD2.n52 VDD2.n0 3.49141
R1363 VDD2.n103 VDD2.n102 2.71565
R1364 VDD2.n85 VDD2.n64 2.71565
R1365 VDD2.n31 VDD2.n10 2.71565
R1366 VDD2.n50 VDD2.n49 2.71565
R1367 VDD2.n72 VDD2.n71 2.41283
R1368 VDD2.n18 VDD2.n17 2.41283
R1369 VDD2.n99 VDD2.n55 1.93989
R1370 VDD2.n86 VDD2.n62 1.93989
R1371 VDD2.n32 VDD2.n8 1.93989
R1372 VDD2.n46 VDD2.n2 1.93989
R1373 VDD2.n98 VDD2.n57 1.16414
R1374 VDD2.n90 VDD2.n89 1.16414
R1375 VDD2.n37 VDD2.n35 1.16414
R1376 VDD2.n45 VDD2.n4 1.16414
R1377 VDD2 VDD2.n106 0.463862
R1378 VDD2.n95 VDD2.n94 0.388379
R1379 VDD2.n61 VDD2.n59 0.388379
R1380 VDD2.n36 VDD2.n6 0.388379
R1381 VDD2.n42 VDD2.n41 0.388379
R1382 VDD2.n104 VDD2.n54 0.155672
R1383 VDD2.n97 VDD2.n54 0.155672
R1384 VDD2.n97 VDD2.n96 0.155672
R1385 VDD2.n96 VDD2.n58 0.155672
R1386 VDD2.n88 VDD2.n58 0.155672
R1387 VDD2.n88 VDD2.n87 0.155672
R1388 VDD2.n87 VDD2.n63 0.155672
R1389 VDD2.n80 VDD2.n63 0.155672
R1390 VDD2.n80 VDD2.n79 0.155672
R1391 VDD2.n79 VDD2.n67 0.155672
R1392 VDD2.n72 VDD2.n67 0.155672
R1393 VDD2.n18 VDD2.n13 0.155672
R1394 VDD2.n25 VDD2.n13 0.155672
R1395 VDD2.n26 VDD2.n25 0.155672
R1396 VDD2.n26 VDD2.n9 0.155672
R1397 VDD2.n33 VDD2.n9 0.155672
R1398 VDD2.n34 VDD2.n33 0.155672
R1399 VDD2.n34 VDD2.n5 0.155672
R1400 VDD2.n43 VDD2.n5 0.155672
R1401 VDD2.n44 VDD2.n43 0.155672
R1402 VDD2.n44 VDD2.n1 0.155672
R1403 VDD2.n51 VDD2.n1 0.155672
C0 VP VN 4.57627f
C1 VP w_n1722_n2954# 2.45661f
C2 VTAIL VP 1.82485f
C3 VDD2 VP 0.28885f
C4 B VN 0.848123f
C5 VDD1 VN 0.147641f
C6 B w_n1722_n2954# 7.09352f
C7 w_n1722_n2954# VDD1 1.51655f
C8 B VTAIL 2.76048f
C9 B VDD2 1.41879f
C10 VDD2 VDD1 0.551419f
C11 VTAIL VDD1 4.44601f
C12 w_n1722_n2954# VN 2.23953f
C13 B VP 1.20081f
C14 VP VDD1 2.26324f
C15 VDD2 VN 2.1248f
C16 VTAIL VN 1.81049f
C17 VTAIL w_n1722_n2954# 2.47926f
C18 VDD2 w_n1722_n2954# 1.5299f
C19 VTAIL VDD2 4.48875f
C20 B VDD1 1.39798f
C21 VDD2 VSUBS 0.740381f
C22 VDD1 VSUBS 3.122201f
C23 VTAIL VSUBS 0.784528f
C24 VN VSUBS 6.20167f
C25 VP VSUBS 1.283502f
C26 B VSUBS 2.942392f
C27 w_n1722_n2954# VSUBS 62.8392f
C28 VDD2.n0 VSUBS 0.020928f
C29 VDD2.n1 VSUBS 0.020298f
C30 VDD2.n2 VSUBS 0.010907f
C31 VDD2.n3 VSUBS 0.025781f
C32 VDD2.n4 VSUBS 0.011549f
C33 VDD2.n5 VSUBS 0.020298f
C34 VDD2.n6 VSUBS 0.011228f
C35 VDD2.n7 VSUBS 0.025781f
C36 VDD2.n8 VSUBS 0.011549f
C37 VDD2.n9 VSUBS 0.020298f
C38 VDD2.n10 VSUBS 0.010907f
C39 VDD2.n11 VSUBS 0.025781f
C40 VDD2.n12 VSUBS 0.011549f
C41 VDD2.n13 VSUBS 0.020298f
C42 VDD2.n14 VSUBS 0.010907f
C43 VDD2.n15 VSUBS 0.019336f
C44 VDD2.n16 VSUBS 0.019394f
C45 VDD2.t0 VSUBS 0.055425f
C46 VDD2.n17 VSUBS 0.14087f
C47 VDD2.n18 VSUBS 0.813178f
C48 VDD2.n19 VSUBS 0.010907f
C49 VDD2.n20 VSUBS 0.011549f
C50 VDD2.n21 VSUBS 0.025781f
C51 VDD2.n22 VSUBS 0.025781f
C52 VDD2.n23 VSUBS 0.011549f
C53 VDD2.n24 VSUBS 0.010907f
C54 VDD2.n25 VSUBS 0.020298f
C55 VDD2.n26 VSUBS 0.020298f
C56 VDD2.n27 VSUBS 0.010907f
C57 VDD2.n28 VSUBS 0.011549f
C58 VDD2.n29 VSUBS 0.025781f
C59 VDD2.n30 VSUBS 0.025781f
C60 VDD2.n31 VSUBS 0.011549f
C61 VDD2.n32 VSUBS 0.010907f
C62 VDD2.n33 VSUBS 0.020298f
C63 VDD2.n34 VSUBS 0.020298f
C64 VDD2.n35 VSUBS 0.010907f
C65 VDD2.n36 VSUBS 0.010907f
C66 VDD2.n37 VSUBS 0.011549f
C67 VDD2.n38 VSUBS 0.025781f
C68 VDD2.n39 VSUBS 0.025781f
C69 VDD2.n40 VSUBS 0.025781f
C70 VDD2.n41 VSUBS 0.011228f
C71 VDD2.n42 VSUBS 0.010907f
C72 VDD2.n43 VSUBS 0.020298f
C73 VDD2.n44 VSUBS 0.020298f
C74 VDD2.n45 VSUBS 0.010907f
C75 VDD2.n46 VSUBS 0.011549f
C76 VDD2.n47 VSUBS 0.025781f
C77 VDD2.n48 VSUBS 0.057727f
C78 VDD2.n49 VSUBS 0.011549f
C79 VDD2.n50 VSUBS 0.010907f
C80 VDD2.n51 VSUBS 0.046086f
C81 VDD2.n52 VSUBS 0.485676f
C82 VDD2.n53 VSUBS 0.020928f
C83 VDD2.n54 VSUBS 0.020298f
C84 VDD2.n55 VSUBS 0.010907f
C85 VDD2.n56 VSUBS 0.025781f
C86 VDD2.n57 VSUBS 0.011549f
C87 VDD2.n58 VSUBS 0.020298f
C88 VDD2.n59 VSUBS 0.011228f
C89 VDD2.n60 VSUBS 0.025781f
C90 VDD2.n61 VSUBS 0.010907f
C91 VDD2.n62 VSUBS 0.011549f
C92 VDD2.n63 VSUBS 0.020298f
C93 VDD2.n64 VSUBS 0.010907f
C94 VDD2.n65 VSUBS 0.025781f
C95 VDD2.n66 VSUBS 0.011549f
C96 VDD2.n67 VSUBS 0.020298f
C97 VDD2.n68 VSUBS 0.010907f
C98 VDD2.n69 VSUBS 0.019336f
C99 VDD2.n70 VSUBS 0.019394f
C100 VDD2.t1 VSUBS 0.055425f
C101 VDD2.n71 VSUBS 0.14087f
C102 VDD2.n72 VSUBS 0.813178f
C103 VDD2.n73 VSUBS 0.010907f
C104 VDD2.n74 VSUBS 0.011549f
C105 VDD2.n75 VSUBS 0.025781f
C106 VDD2.n76 VSUBS 0.025781f
C107 VDD2.n77 VSUBS 0.011549f
C108 VDD2.n78 VSUBS 0.010907f
C109 VDD2.n79 VSUBS 0.020298f
C110 VDD2.n80 VSUBS 0.020298f
C111 VDD2.n81 VSUBS 0.010907f
C112 VDD2.n82 VSUBS 0.011549f
C113 VDD2.n83 VSUBS 0.025781f
C114 VDD2.n84 VSUBS 0.025781f
C115 VDD2.n85 VSUBS 0.011549f
C116 VDD2.n86 VSUBS 0.010907f
C117 VDD2.n87 VSUBS 0.020298f
C118 VDD2.n88 VSUBS 0.020298f
C119 VDD2.n89 VSUBS 0.010907f
C120 VDD2.n90 VSUBS 0.011549f
C121 VDD2.n91 VSUBS 0.025781f
C122 VDD2.n92 VSUBS 0.025781f
C123 VDD2.n93 VSUBS 0.025781f
C124 VDD2.n94 VSUBS 0.011228f
C125 VDD2.n95 VSUBS 0.010907f
C126 VDD2.n96 VSUBS 0.020298f
C127 VDD2.n97 VSUBS 0.020298f
C128 VDD2.n98 VSUBS 0.010907f
C129 VDD2.n99 VSUBS 0.011549f
C130 VDD2.n100 VSUBS 0.025781f
C131 VDD2.n101 VSUBS 0.057727f
C132 VDD2.n102 VSUBS 0.011549f
C133 VDD2.n103 VSUBS 0.010907f
C134 VDD2.n104 VSUBS 0.046086f
C135 VDD2.n105 VSUBS 0.042819f
C136 VDD2.n106 VSUBS 2.13095f
C137 VN.t1 VSUBS 2.15188f
C138 VN.t0 VSUBS 2.45798f
C139 VDD1.n0 VSUBS 0.021006f
C140 VDD1.n1 VSUBS 0.020374f
C141 VDD1.n2 VSUBS 0.010948f
C142 VDD1.n3 VSUBS 0.025877f
C143 VDD1.n4 VSUBS 0.011592f
C144 VDD1.n5 VSUBS 0.020374f
C145 VDD1.n6 VSUBS 0.01127f
C146 VDD1.n7 VSUBS 0.025877f
C147 VDD1.n8 VSUBS 0.010948f
C148 VDD1.n9 VSUBS 0.011592f
C149 VDD1.n10 VSUBS 0.020374f
C150 VDD1.n11 VSUBS 0.010948f
C151 VDD1.n12 VSUBS 0.025877f
C152 VDD1.n13 VSUBS 0.011592f
C153 VDD1.n14 VSUBS 0.020374f
C154 VDD1.n15 VSUBS 0.010948f
C155 VDD1.n16 VSUBS 0.019408f
C156 VDD1.n17 VSUBS 0.019466f
C157 VDD1.t1 VSUBS 0.055632f
C158 VDD1.n18 VSUBS 0.141398f
C159 VDD1.n19 VSUBS 0.816227f
C160 VDD1.n20 VSUBS 0.010948f
C161 VDD1.n21 VSUBS 0.011592f
C162 VDD1.n22 VSUBS 0.025877f
C163 VDD1.n23 VSUBS 0.025877f
C164 VDD1.n24 VSUBS 0.011592f
C165 VDD1.n25 VSUBS 0.010948f
C166 VDD1.n26 VSUBS 0.020374f
C167 VDD1.n27 VSUBS 0.020374f
C168 VDD1.n28 VSUBS 0.010948f
C169 VDD1.n29 VSUBS 0.011592f
C170 VDD1.n30 VSUBS 0.025877f
C171 VDD1.n31 VSUBS 0.025877f
C172 VDD1.n32 VSUBS 0.011592f
C173 VDD1.n33 VSUBS 0.010948f
C174 VDD1.n34 VSUBS 0.020374f
C175 VDD1.n35 VSUBS 0.020374f
C176 VDD1.n36 VSUBS 0.010948f
C177 VDD1.n37 VSUBS 0.011592f
C178 VDD1.n38 VSUBS 0.025877f
C179 VDD1.n39 VSUBS 0.025877f
C180 VDD1.n40 VSUBS 0.025877f
C181 VDD1.n41 VSUBS 0.01127f
C182 VDD1.n42 VSUBS 0.010948f
C183 VDD1.n43 VSUBS 0.020374f
C184 VDD1.n44 VSUBS 0.020374f
C185 VDD1.n45 VSUBS 0.010948f
C186 VDD1.n46 VSUBS 0.011592f
C187 VDD1.n47 VSUBS 0.025877f
C188 VDD1.n48 VSUBS 0.057943f
C189 VDD1.n49 VSUBS 0.011592f
C190 VDD1.n50 VSUBS 0.010948f
C191 VDD1.n51 VSUBS 0.046259f
C192 VDD1.n52 VSUBS 0.043637f
C193 VDD1.n53 VSUBS 0.021006f
C194 VDD1.n54 VSUBS 0.020374f
C195 VDD1.n55 VSUBS 0.010948f
C196 VDD1.n56 VSUBS 0.025877f
C197 VDD1.n57 VSUBS 0.011592f
C198 VDD1.n58 VSUBS 0.020374f
C199 VDD1.n59 VSUBS 0.01127f
C200 VDD1.n60 VSUBS 0.025877f
C201 VDD1.n61 VSUBS 0.011592f
C202 VDD1.n62 VSUBS 0.020374f
C203 VDD1.n63 VSUBS 0.010948f
C204 VDD1.n64 VSUBS 0.025877f
C205 VDD1.n65 VSUBS 0.011592f
C206 VDD1.n66 VSUBS 0.020374f
C207 VDD1.n67 VSUBS 0.010948f
C208 VDD1.n68 VSUBS 0.019408f
C209 VDD1.n69 VSUBS 0.019466f
C210 VDD1.t0 VSUBS 0.055632f
C211 VDD1.n70 VSUBS 0.141398f
C212 VDD1.n71 VSUBS 0.816227f
C213 VDD1.n72 VSUBS 0.010948f
C214 VDD1.n73 VSUBS 0.011592f
C215 VDD1.n74 VSUBS 0.025877f
C216 VDD1.n75 VSUBS 0.025877f
C217 VDD1.n76 VSUBS 0.011592f
C218 VDD1.n77 VSUBS 0.010948f
C219 VDD1.n78 VSUBS 0.020374f
C220 VDD1.n79 VSUBS 0.020374f
C221 VDD1.n80 VSUBS 0.010948f
C222 VDD1.n81 VSUBS 0.011592f
C223 VDD1.n82 VSUBS 0.025877f
C224 VDD1.n83 VSUBS 0.025877f
C225 VDD1.n84 VSUBS 0.011592f
C226 VDD1.n85 VSUBS 0.010948f
C227 VDD1.n86 VSUBS 0.020374f
C228 VDD1.n87 VSUBS 0.020374f
C229 VDD1.n88 VSUBS 0.010948f
C230 VDD1.n89 VSUBS 0.010948f
C231 VDD1.n90 VSUBS 0.011592f
C232 VDD1.n91 VSUBS 0.025877f
C233 VDD1.n92 VSUBS 0.025877f
C234 VDD1.n93 VSUBS 0.025877f
C235 VDD1.n94 VSUBS 0.01127f
C236 VDD1.n95 VSUBS 0.010948f
C237 VDD1.n96 VSUBS 0.020374f
C238 VDD1.n97 VSUBS 0.020374f
C239 VDD1.n98 VSUBS 0.010948f
C240 VDD1.n99 VSUBS 0.011592f
C241 VDD1.n100 VSUBS 0.025877f
C242 VDD1.n101 VSUBS 0.057943f
C243 VDD1.n102 VSUBS 0.011592f
C244 VDD1.n103 VSUBS 0.010948f
C245 VDD1.n104 VSUBS 0.046259f
C246 VDD1.n105 VSUBS 0.519137f
C247 VTAIL.n0 VSUBS 0.02434f
C248 VTAIL.n1 VSUBS 0.023607f
C249 VTAIL.n2 VSUBS 0.012686f
C250 VTAIL.n3 VSUBS 0.029984f
C251 VTAIL.n4 VSUBS 0.013432f
C252 VTAIL.n5 VSUBS 0.023607f
C253 VTAIL.n6 VSUBS 0.013059f
C254 VTAIL.n7 VSUBS 0.029984f
C255 VTAIL.n8 VSUBS 0.013432f
C256 VTAIL.n9 VSUBS 0.023607f
C257 VTAIL.n10 VSUBS 0.012686f
C258 VTAIL.n11 VSUBS 0.029984f
C259 VTAIL.n12 VSUBS 0.013432f
C260 VTAIL.n13 VSUBS 0.023607f
C261 VTAIL.n14 VSUBS 0.012686f
C262 VTAIL.n15 VSUBS 0.022488f
C263 VTAIL.n16 VSUBS 0.022556f
C264 VTAIL.t3 VSUBS 0.064461f
C265 VTAIL.n17 VSUBS 0.163838f
C266 VTAIL.n18 VSUBS 0.94576f
C267 VTAIL.n19 VSUBS 0.012686f
C268 VTAIL.n20 VSUBS 0.013432f
C269 VTAIL.n21 VSUBS 0.029984f
C270 VTAIL.n22 VSUBS 0.029984f
C271 VTAIL.n23 VSUBS 0.013432f
C272 VTAIL.n24 VSUBS 0.012686f
C273 VTAIL.n25 VSUBS 0.023607f
C274 VTAIL.n26 VSUBS 0.023607f
C275 VTAIL.n27 VSUBS 0.012686f
C276 VTAIL.n28 VSUBS 0.013432f
C277 VTAIL.n29 VSUBS 0.029984f
C278 VTAIL.n30 VSUBS 0.029984f
C279 VTAIL.n31 VSUBS 0.013432f
C280 VTAIL.n32 VSUBS 0.012686f
C281 VTAIL.n33 VSUBS 0.023607f
C282 VTAIL.n34 VSUBS 0.023607f
C283 VTAIL.n35 VSUBS 0.012686f
C284 VTAIL.n36 VSUBS 0.012686f
C285 VTAIL.n37 VSUBS 0.013432f
C286 VTAIL.n38 VSUBS 0.029984f
C287 VTAIL.n39 VSUBS 0.029984f
C288 VTAIL.n40 VSUBS 0.029984f
C289 VTAIL.n41 VSUBS 0.013059f
C290 VTAIL.n42 VSUBS 0.012686f
C291 VTAIL.n43 VSUBS 0.023607f
C292 VTAIL.n44 VSUBS 0.023607f
C293 VTAIL.n45 VSUBS 0.012686f
C294 VTAIL.n46 VSUBS 0.013432f
C295 VTAIL.n47 VSUBS 0.029984f
C296 VTAIL.n48 VSUBS 0.067139f
C297 VTAIL.n49 VSUBS 0.013432f
C298 VTAIL.n50 VSUBS 0.012686f
C299 VTAIL.n51 VSUBS 0.0536f
C300 VTAIL.n52 VSUBS 0.033492f
C301 VTAIL.n53 VSUBS 1.30902f
C302 VTAIL.n54 VSUBS 0.02434f
C303 VTAIL.n55 VSUBS 0.023607f
C304 VTAIL.n56 VSUBS 0.012686f
C305 VTAIL.n57 VSUBS 0.029984f
C306 VTAIL.n58 VSUBS 0.013432f
C307 VTAIL.n59 VSUBS 0.023607f
C308 VTAIL.n60 VSUBS 0.013059f
C309 VTAIL.n61 VSUBS 0.029984f
C310 VTAIL.n62 VSUBS 0.012686f
C311 VTAIL.n63 VSUBS 0.013432f
C312 VTAIL.n64 VSUBS 0.023607f
C313 VTAIL.n65 VSUBS 0.012686f
C314 VTAIL.n66 VSUBS 0.029984f
C315 VTAIL.n67 VSUBS 0.013432f
C316 VTAIL.n68 VSUBS 0.023607f
C317 VTAIL.n69 VSUBS 0.012686f
C318 VTAIL.n70 VSUBS 0.022488f
C319 VTAIL.n71 VSUBS 0.022556f
C320 VTAIL.t1 VSUBS 0.064461f
C321 VTAIL.n72 VSUBS 0.163838f
C322 VTAIL.n73 VSUBS 0.94576f
C323 VTAIL.n74 VSUBS 0.012686f
C324 VTAIL.n75 VSUBS 0.013432f
C325 VTAIL.n76 VSUBS 0.029984f
C326 VTAIL.n77 VSUBS 0.029984f
C327 VTAIL.n78 VSUBS 0.013432f
C328 VTAIL.n79 VSUBS 0.012686f
C329 VTAIL.n80 VSUBS 0.023607f
C330 VTAIL.n81 VSUBS 0.023607f
C331 VTAIL.n82 VSUBS 0.012686f
C332 VTAIL.n83 VSUBS 0.013432f
C333 VTAIL.n84 VSUBS 0.029984f
C334 VTAIL.n85 VSUBS 0.029984f
C335 VTAIL.n86 VSUBS 0.013432f
C336 VTAIL.n87 VSUBS 0.012686f
C337 VTAIL.n88 VSUBS 0.023607f
C338 VTAIL.n89 VSUBS 0.023607f
C339 VTAIL.n90 VSUBS 0.012686f
C340 VTAIL.n91 VSUBS 0.013432f
C341 VTAIL.n92 VSUBS 0.029984f
C342 VTAIL.n93 VSUBS 0.029984f
C343 VTAIL.n94 VSUBS 0.029984f
C344 VTAIL.n95 VSUBS 0.013059f
C345 VTAIL.n96 VSUBS 0.012686f
C346 VTAIL.n97 VSUBS 0.023607f
C347 VTAIL.n98 VSUBS 0.023607f
C348 VTAIL.n99 VSUBS 0.012686f
C349 VTAIL.n100 VSUBS 0.013432f
C350 VTAIL.n101 VSUBS 0.029984f
C351 VTAIL.n102 VSUBS 0.067139f
C352 VTAIL.n103 VSUBS 0.013432f
C353 VTAIL.n104 VSUBS 0.012686f
C354 VTAIL.n105 VSUBS 0.0536f
C355 VTAIL.n106 VSUBS 0.033492f
C356 VTAIL.n107 VSUBS 1.33541f
C357 VTAIL.n108 VSUBS 0.02434f
C358 VTAIL.n109 VSUBS 0.023607f
C359 VTAIL.n110 VSUBS 0.012686f
C360 VTAIL.n111 VSUBS 0.029984f
C361 VTAIL.n112 VSUBS 0.013432f
C362 VTAIL.n113 VSUBS 0.023607f
C363 VTAIL.n114 VSUBS 0.013059f
C364 VTAIL.n115 VSUBS 0.029984f
C365 VTAIL.n116 VSUBS 0.012686f
C366 VTAIL.n117 VSUBS 0.013432f
C367 VTAIL.n118 VSUBS 0.023607f
C368 VTAIL.n119 VSUBS 0.012686f
C369 VTAIL.n120 VSUBS 0.029984f
C370 VTAIL.n121 VSUBS 0.013432f
C371 VTAIL.n122 VSUBS 0.023607f
C372 VTAIL.n123 VSUBS 0.012686f
C373 VTAIL.n124 VSUBS 0.022488f
C374 VTAIL.n125 VSUBS 0.022556f
C375 VTAIL.t2 VSUBS 0.064461f
C376 VTAIL.n126 VSUBS 0.163838f
C377 VTAIL.n127 VSUBS 0.94576f
C378 VTAIL.n128 VSUBS 0.012686f
C379 VTAIL.n129 VSUBS 0.013432f
C380 VTAIL.n130 VSUBS 0.029984f
C381 VTAIL.n131 VSUBS 0.029984f
C382 VTAIL.n132 VSUBS 0.013432f
C383 VTAIL.n133 VSUBS 0.012686f
C384 VTAIL.n134 VSUBS 0.023607f
C385 VTAIL.n135 VSUBS 0.023607f
C386 VTAIL.n136 VSUBS 0.012686f
C387 VTAIL.n137 VSUBS 0.013432f
C388 VTAIL.n138 VSUBS 0.029984f
C389 VTAIL.n139 VSUBS 0.029984f
C390 VTAIL.n140 VSUBS 0.013432f
C391 VTAIL.n141 VSUBS 0.012686f
C392 VTAIL.n142 VSUBS 0.023607f
C393 VTAIL.n143 VSUBS 0.023607f
C394 VTAIL.n144 VSUBS 0.012686f
C395 VTAIL.n145 VSUBS 0.013432f
C396 VTAIL.n146 VSUBS 0.029984f
C397 VTAIL.n147 VSUBS 0.029984f
C398 VTAIL.n148 VSUBS 0.029984f
C399 VTAIL.n149 VSUBS 0.013059f
C400 VTAIL.n150 VSUBS 0.012686f
C401 VTAIL.n151 VSUBS 0.023607f
C402 VTAIL.n152 VSUBS 0.023607f
C403 VTAIL.n153 VSUBS 0.012686f
C404 VTAIL.n154 VSUBS 0.013432f
C405 VTAIL.n155 VSUBS 0.029984f
C406 VTAIL.n156 VSUBS 0.067139f
C407 VTAIL.n157 VSUBS 0.013432f
C408 VTAIL.n158 VSUBS 0.012686f
C409 VTAIL.n159 VSUBS 0.0536f
C410 VTAIL.n160 VSUBS 0.033492f
C411 VTAIL.n161 VSUBS 1.21213f
C412 VTAIL.n162 VSUBS 0.02434f
C413 VTAIL.n163 VSUBS 0.023607f
C414 VTAIL.n164 VSUBS 0.012686f
C415 VTAIL.n165 VSUBS 0.029984f
C416 VTAIL.n166 VSUBS 0.013432f
C417 VTAIL.n167 VSUBS 0.023607f
C418 VTAIL.n168 VSUBS 0.013059f
C419 VTAIL.n169 VSUBS 0.029984f
C420 VTAIL.n170 VSUBS 0.013432f
C421 VTAIL.n171 VSUBS 0.023607f
C422 VTAIL.n172 VSUBS 0.012686f
C423 VTAIL.n173 VSUBS 0.029984f
C424 VTAIL.n174 VSUBS 0.013432f
C425 VTAIL.n175 VSUBS 0.023607f
C426 VTAIL.n176 VSUBS 0.012686f
C427 VTAIL.n177 VSUBS 0.022488f
C428 VTAIL.n178 VSUBS 0.022556f
C429 VTAIL.t0 VSUBS 0.064461f
C430 VTAIL.n179 VSUBS 0.163838f
C431 VTAIL.n180 VSUBS 0.94576f
C432 VTAIL.n181 VSUBS 0.012686f
C433 VTAIL.n182 VSUBS 0.013432f
C434 VTAIL.n183 VSUBS 0.029984f
C435 VTAIL.n184 VSUBS 0.029984f
C436 VTAIL.n185 VSUBS 0.013432f
C437 VTAIL.n186 VSUBS 0.012686f
C438 VTAIL.n187 VSUBS 0.023607f
C439 VTAIL.n188 VSUBS 0.023607f
C440 VTAIL.n189 VSUBS 0.012686f
C441 VTAIL.n190 VSUBS 0.013432f
C442 VTAIL.n191 VSUBS 0.029984f
C443 VTAIL.n192 VSUBS 0.029984f
C444 VTAIL.n193 VSUBS 0.013432f
C445 VTAIL.n194 VSUBS 0.012686f
C446 VTAIL.n195 VSUBS 0.023607f
C447 VTAIL.n196 VSUBS 0.023607f
C448 VTAIL.n197 VSUBS 0.012686f
C449 VTAIL.n198 VSUBS 0.012686f
C450 VTAIL.n199 VSUBS 0.013432f
C451 VTAIL.n200 VSUBS 0.029984f
C452 VTAIL.n201 VSUBS 0.029984f
C453 VTAIL.n202 VSUBS 0.029984f
C454 VTAIL.n203 VSUBS 0.013059f
C455 VTAIL.n204 VSUBS 0.012686f
C456 VTAIL.n205 VSUBS 0.023607f
C457 VTAIL.n206 VSUBS 0.023607f
C458 VTAIL.n207 VSUBS 0.012686f
C459 VTAIL.n208 VSUBS 0.013432f
C460 VTAIL.n209 VSUBS 0.029984f
C461 VTAIL.n210 VSUBS 0.067139f
C462 VTAIL.n211 VSUBS 0.013432f
C463 VTAIL.n212 VSUBS 0.012686f
C464 VTAIL.n213 VSUBS 0.0536f
C465 VTAIL.n214 VSUBS 0.033492f
C466 VTAIL.n215 VSUBS 1.14114f
C467 VP.t0 VSUBS 2.60851f
C468 VP.t1 VSUBS 2.2881f
C469 VP.n0 VSUBS 4.45407f
C470 B.n0 VSUBS 0.004482f
C471 B.n1 VSUBS 0.004482f
C472 B.n2 VSUBS 0.007088f
C473 B.n3 VSUBS 0.007088f
C474 B.n4 VSUBS 0.007088f
C475 B.n5 VSUBS 0.007088f
C476 B.n6 VSUBS 0.007088f
C477 B.n7 VSUBS 0.007088f
C478 B.n8 VSUBS 0.007088f
C479 B.n9 VSUBS 0.007088f
C480 B.n10 VSUBS 0.007088f
C481 B.n11 VSUBS 0.015819f
C482 B.n12 VSUBS 0.007088f
C483 B.n13 VSUBS 0.007088f
C484 B.n14 VSUBS 0.007088f
C485 B.n15 VSUBS 0.007088f
C486 B.n16 VSUBS 0.007088f
C487 B.n17 VSUBS 0.007088f
C488 B.n18 VSUBS 0.007088f
C489 B.n19 VSUBS 0.007088f
C490 B.n20 VSUBS 0.007088f
C491 B.n21 VSUBS 0.007088f
C492 B.n22 VSUBS 0.007088f
C493 B.n23 VSUBS 0.007088f
C494 B.n24 VSUBS 0.007088f
C495 B.n25 VSUBS 0.007088f
C496 B.n26 VSUBS 0.007088f
C497 B.n27 VSUBS 0.007088f
C498 B.n28 VSUBS 0.007088f
C499 B.n29 VSUBS 0.007088f
C500 B.t8 VSUBS 0.167984f
C501 B.t7 VSUBS 0.188459f
C502 B.t6 VSUBS 0.692426f
C503 B.n30 VSUBS 0.301446f
C504 B.n31 VSUBS 0.220519f
C505 B.n32 VSUBS 0.007088f
C506 B.n33 VSUBS 0.007088f
C507 B.n34 VSUBS 0.007088f
C508 B.n35 VSUBS 0.007088f
C509 B.t11 VSUBS 0.167986f
C510 B.t10 VSUBS 0.188461f
C511 B.t9 VSUBS 0.692426f
C512 B.n36 VSUBS 0.301443f
C513 B.n37 VSUBS 0.220516f
C514 B.n38 VSUBS 0.016423f
C515 B.n39 VSUBS 0.007088f
C516 B.n40 VSUBS 0.007088f
C517 B.n41 VSUBS 0.007088f
C518 B.n42 VSUBS 0.007088f
C519 B.n43 VSUBS 0.007088f
C520 B.n44 VSUBS 0.007088f
C521 B.n45 VSUBS 0.007088f
C522 B.n46 VSUBS 0.007088f
C523 B.n47 VSUBS 0.007088f
C524 B.n48 VSUBS 0.007088f
C525 B.n49 VSUBS 0.007088f
C526 B.n50 VSUBS 0.007088f
C527 B.n51 VSUBS 0.007088f
C528 B.n52 VSUBS 0.007088f
C529 B.n53 VSUBS 0.007088f
C530 B.n54 VSUBS 0.007088f
C531 B.n55 VSUBS 0.007088f
C532 B.n56 VSUBS 0.016274f
C533 B.n57 VSUBS 0.007088f
C534 B.n58 VSUBS 0.007088f
C535 B.n59 VSUBS 0.007088f
C536 B.n60 VSUBS 0.007088f
C537 B.n61 VSUBS 0.007088f
C538 B.n62 VSUBS 0.007088f
C539 B.n63 VSUBS 0.007088f
C540 B.n64 VSUBS 0.007088f
C541 B.n65 VSUBS 0.007088f
C542 B.n66 VSUBS 0.007088f
C543 B.n67 VSUBS 0.007088f
C544 B.n68 VSUBS 0.007088f
C545 B.n69 VSUBS 0.007088f
C546 B.n70 VSUBS 0.007088f
C547 B.n71 VSUBS 0.007088f
C548 B.n72 VSUBS 0.007088f
C549 B.n73 VSUBS 0.007088f
C550 B.n74 VSUBS 0.007088f
C551 B.n75 VSUBS 0.007088f
C552 B.n76 VSUBS 0.01712f
C553 B.n77 VSUBS 0.007088f
C554 B.n78 VSUBS 0.007088f
C555 B.n79 VSUBS 0.007088f
C556 B.n80 VSUBS 0.007088f
C557 B.n81 VSUBS 0.007088f
C558 B.n82 VSUBS 0.007088f
C559 B.n83 VSUBS 0.007088f
C560 B.n84 VSUBS 0.007088f
C561 B.n85 VSUBS 0.007088f
C562 B.n86 VSUBS 0.007088f
C563 B.n87 VSUBS 0.007088f
C564 B.n88 VSUBS 0.007088f
C565 B.n89 VSUBS 0.007088f
C566 B.n90 VSUBS 0.007088f
C567 B.n91 VSUBS 0.007088f
C568 B.n92 VSUBS 0.007088f
C569 B.n93 VSUBS 0.007088f
C570 B.t4 VSUBS 0.167986f
C571 B.t5 VSUBS 0.188461f
C572 B.t3 VSUBS 0.692426f
C573 B.n94 VSUBS 0.301443f
C574 B.n95 VSUBS 0.220516f
C575 B.n96 VSUBS 0.016423f
C576 B.n97 VSUBS 0.007088f
C577 B.n98 VSUBS 0.007088f
C578 B.n99 VSUBS 0.007088f
C579 B.n100 VSUBS 0.007088f
C580 B.n101 VSUBS 0.007088f
C581 B.t1 VSUBS 0.167984f
C582 B.t2 VSUBS 0.188459f
C583 B.t0 VSUBS 0.692426f
C584 B.n102 VSUBS 0.301446f
C585 B.n103 VSUBS 0.220519f
C586 B.n104 VSUBS 0.007088f
C587 B.n105 VSUBS 0.007088f
C588 B.n106 VSUBS 0.007088f
C589 B.n107 VSUBS 0.007088f
C590 B.n108 VSUBS 0.007088f
C591 B.n109 VSUBS 0.007088f
C592 B.n110 VSUBS 0.007088f
C593 B.n111 VSUBS 0.007088f
C594 B.n112 VSUBS 0.007088f
C595 B.n113 VSUBS 0.007088f
C596 B.n114 VSUBS 0.007088f
C597 B.n115 VSUBS 0.007088f
C598 B.n116 VSUBS 0.007088f
C599 B.n117 VSUBS 0.007088f
C600 B.n118 VSUBS 0.007088f
C601 B.n119 VSUBS 0.007088f
C602 B.n120 VSUBS 0.007088f
C603 B.n121 VSUBS 0.015819f
C604 B.n122 VSUBS 0.007088f
C605 B.n123 VSUBS 0.007088f
C606 B.n124 VSUBS 0.007088f
C607 B.n125 VSUBS 0.007088f
C608 B.n126 VSUBS 0.007088f
C609 B.n127 VSUBS 0.007088f
C610 B.n128 VSUBS 0.007088f
C611 B.n129 VSUBS 0.007088f
C612 B.n130 VSUBS 0.007088f
C613 B.n131 VSUBS 0.007088f
C614 B.n132 VSUBS 0.007088f
C615 B.n133 VSUBS 0.007088f
C616 B.n134 VSUBS 0.007088f
C617 B.n135 VSUBS 0.007088f
C618 B.n136 VSUBS 0.007088f
C619 B.n137 VSUBS 0.007088f
C620 B.n138 VSUBS 0.007088f
C621 B.n139 VSUBS 0.007088f
C622 B.n140 VSUBS 0.007088f
C623 B.n141 VSUBS 0.007088f
C624 B.n142 VSUBS 0.007088f
C625 B.n143 VSUBS 0.007088f
C626 B.n144 VSUBS 0.007088f
C627 B.n145 VSUBS 0.007088f
C628 B.n146 VSUBS 0.007088f
C629 B.n147 VSUBS 0.007088f
C630 B.n148 VSUBS 0.007088f
C631 B.n149 VSUBS 0.007088f
C632 B.n150 VSUBS 0.007088f
C633 B.n151 VSUBS 0.007088f
C634 B.n152 VSUBS 0.007088f
C635 B.n153 VSUBS 0.007088f
C636 B.n154 VSUBS 0.007088f
C637 B.n155 VSUBS 0.007088f
C638 B.n156 VSUBS 0.015819f
C639 B.n157 VSUBS 0.01712f
C640 B.n158 VSUBS 0.01712f
C641 B.n159 VSUBS 0.007088f
C642 B.n160 VSUBS 0.007088f
C643 B.n161 VSUBS 0.007088f
C644 B.n162 VSUBS 0.007088f
C645 B.n163 VSUBS 0.007088f
C646 B.n164 VSUBS 0.007088f
C647 B.n165 VSUBS 0.007088f
C648 B.n166 VSUBS 0.007088f
C649 B.n167 VSUBS 0.007088f
C650 B.n168 VSUBS 0.007088f
C651 B.n169 VSUBS 0.007088f
C652 B.n170 VSUBS 0.007088f
C653 B.n171 VSUBS 0.007088f
C654 B.n172 VSUBS 0.007088f
C655 B.n173 VSUBS 0.007088f
C656 B.n174 VSUBS 0.007088f
C657 B.n175 VSUBS 0.007088f
C658 B.n176 VSUBS 0.007088f
C659 B.n177 VSUBS 0.007088f
C660 B.n178 VSUBS 0.007088f
C661 B.n179 VSUBS 0.007088f
C662 B.n180 VSUBS 0.007088f
C663 B.n181 VSUBS 0.007088f
C664 B.n182 VSUBS 0.007088f
C665 B.n183 VSUBS 0.007088f
C666 B.n184 VSUBS 0.007088f
C667 B.n185 VSUBS 0.007088f
C668 B.n186 VSUBS 0.007088f
C669 B.n187 VSUBS 0.007088f
C670 B.n188 VSUBS 0.007088f
C671 B.n189 VSUBS 0.007088f
C672 B.n190 VSUBS 0.007088f
C673 B.n191 VSUBS 0.007088f
C674 B.n192 VSUBS 0.007088f
C675 B.n193 VSUBS 0.007088f
C676 B.n194 VSUBS 0.007088f
C677 B.n195 VSUBS 0.007088f
C678 B.n196 VSUBS 0.007088f
C679 B.n197 VSUBS 0.007088f
C680 B.n198 VSUBS 0.007088f
C681 B.n199 VSUBS 0.007088f
C682 B.n200 VSUBS 0.007088f
C683 B.n201 VSUBS 0.007088f
C684 B.n202 VSUBS 0.007088f
C685 B.n203 VSUBS 0.007088f
C686 B.n204 VSUBS 0.007088f
C687 B.n205 VSUBS 0.007088f
C688 B.n206 VSUBS 0.007088f
C689 B.n207 VSUBS 0.007088f
C690 B.n208 VSUBS 0.007088f
C691 B.n209 VSUBS 0.007088f
C692 B.n210 VSUBS 0.004899f
C693 B.n211 VSUBS 0.016423f
C694 B.n212 VSUBS 0.005733f
C695 B.n213 VSUBS 0.007088f
C696 B.n214 VSUBS 0.007088f
C697 B.n215 VSUBS 0.007088f
C698 B.n216 VSUBS 0.007088f
C699 B.n217 VSUBS 0.007088f
C700 B.n218 VSUBS 0.007088f
C701 B.n219 VSUBS 0.007088f
C702 B.n220 VSUBS 0.007088f
C703 B.n221 VSUBS 0.007088f
C704 B.n222 VSUBS 0.007088f
C705 B.n223 VSUBS 0.007088f
C706 B.n224 VSUBS 0.005733f
C707 B.n225 VSUBS 0.007088f
C708 B.n226 VSUBS 0.007088f
C709 B.n227 VSUBS 0.004899f
C710 B.n228 VSUBS 0.007088f
C711 B.n229 VSUBS 0.007088f
C712 B.n230 VSUBS 0.007088f
C713 B.n231 VSUBS 0.007088f
C714 B.n232 VSUBS 0.007088f
C715 B.n233 VSUBS 0.007088f
C716 B.n234 VSUBS 0.007088f
C717 B.n235 VSUBS 0.007088f
C718 B.n236 VSUBS 0.007088f
C719 B.n237 VSUBS 0.007088f
C720 B.n238 VSUBS 0.007088f
C721 B.n239 VSUBS 0.007088f
C722 B.n240 VSUBS 0.007088f
C723 B.n241 VSUBS 0.007088f
C724 B.n242 VSUBS 0.007088f
C725 B.n243 VSUBS 0.007088f
C726 B.n244 VSUBS 0.007088f
C727 B.n245 VSUBS 0.007088f
C728 B.n246 VSUBS 0.007088f
C729 B.n247 VSUBS 0.007088f
C730 B.n248 VSUBS 0.007088f
C731 B.n249 VSUBS 0.007088f
C732 B.n250 VSUBS 0.007088f
C733 B.n251 VSUBS 0.007088f
C734 B.n252 VSUBS 0.007088f
C735 B.n253 VSUBS 0.007088f
C736 B.n254 VSUBS 0.007088f
C737 B.n255 VSUBS 0.007088f
C738 B.n256 VSUBS 0.007088f
C739 B.n257 VSUBS 0.007088f
C740 B.n258 VSUBS 0.007088f
C741 B.n259 VSUBS 0.007088f
C742 B.n260 VSUBS 0.007088f
C743 B.n261 VSUBS 0.007088f
C744 B.n262 VSUBS 0.007088f
C745 B.n263 VSUBS 0.007088f
C746 B.n264 VSUBS 0.007088f
C747 B.n265 VSUBS 0.007088f
C748 B.n266 VSUBS 0.007088f
C749 B.n267 VSUBS 0.007088f
C750 B.n268 VSUBS 0.007088f
C751 B.n269 VSUBS 0.007088f
C752 B.n270 VSUBS 0.007088f
C753 B.n271 VSUBS 0.007088f
C754 B.n272 VSUBS 0.007088f
C755 B.n273 VSUBS 0.007088f
C756 B.n274 VSUBS 0.007088f
C757 B.n275 VSUBS 0.007088f
C758 B.n276 VSUBS 0.007088f
C759 B.n277 VSUBS 0.007088f
C760 B.n278 VSUBS 0.007088f
C761 B.n279 VSUBS 0.01712f
C762 B.n280 VSUBS 0.015819f
C763 B.n281 VSUBS 0.015819f
C764 B.n282 VSUBS 0.007088f
C765 B.n283 VSUBS 0.007088f
C766 B.n284 VSUBS 0.007088f
C767 B.n285 VSUBS 0.007088f
C768 B.n286 VSUBS 0.007088f
C769 B.n287 VSUBS 0.007088f
C770 B.n288 VSUBS 0.007088f
C771 B.n289 VSUBS 0.007088f
C772 B.n290 VSUBS 0.007088f
C773 B.n291 VSUBS 0.007088f
C774 B.n292 VSUBS 0.007088f
C775 B.n293 VSUBS 0.007088f
C776 B.n294 VSUBS 0.007088f
C777 B.n295 VSUBS 0.007088f
C778 B.n296 VSUBS 0.007088f
C779 B.n297 VSUBS 0.007088f
C780 B.n298 VSUBS 0.007088f
C781 B.n299 VSUBS 0.007088f
C782 B.n300 VSUBS 0.007088f
C783 B.n301 VSUBS 0.007088f
C784 B.n302 VSUBS 0.007088f
C785 B.n303 VSUBS 0.007088f
C786 B.n304 VSUBS 0.007088f
C787 B.n305 VSUBS 0.007088f
C788 B.n306 VSUBS 0.007088f
C789 B.n307 VSUBS 0.007088f
C790 B.n308 VSUBS 0.007088f
C791 B.n309 VSUBS 0.007088f
C792 B.n310 VSUBS 0.007088f
C793 B.n311 VSUBS 0.007088f
C794 B.n312 VSUBS 0.007088f
C795 B.n313 VSUBS 0.007088f
C796 B.n314 VSUBS 0.007088f
C797 B.n315 VSUBS 0.007088f
C798 B.n316 VSUBS 0.007088f
C799 B.n317 VSUBS 0.007088f
C800 B.n318 VSUBS 0.007088f
C801 B.n319 VSUBS 0.007088f
C802 B.n320 VSUBS 0.007088f
C803 B.n321 VSUBS 0.007088f
C804 B.n322 VSUBS 0.007088f
C805 B.n323 VSUBS 0.007088f
C806 B.n324 VSUBS 0.007088f
C807 B.n325 VSUBS 0.007088f
C808 B.n326 VSUBS 0.007088f
C809 B.n327 VSUBS 0.007088f
C810 B.n328 VSUBS 0.007088f
C811 B.n329 VSUBS 0.007088f
C812 B.n330 VSUBS 0.007088f
C813 B.n331 VSUBS 0.007088f
C814 B.n332 VSUBS 0.007088f
C815 B.n333 VSUBS 0.007088f
C816 B.n334 VSUBS 0.007088f
C817 B.n335 VSUBS 0.007088f
C818 B.n336 VSUBS 0.007088f
C819 B.n337 VSUBS 0.016666f
C820 B.n338 VSUBS 0.015819f
C821 B.n339 VSUBS 0.01712f
C822 B.n340 VSUBS 0.007088f
C823 B.n341 VSUBS 0.007088f
C824 B.n342 VSUBS 0.007088f
C825 B.n343 VSUBS 0.007088f
C826 B.n344 VSUBS 0.007088f
C827 B.n345 VSUBS 0.007088f
C828 B.n346 VSUBS 0.007088f
C829 B.n347 VSUBS 0.007088f
C830 B.n348 VSUBS 0.007088f
C831 B.n349 VSUBS 0.007088f
C832 B.n350 VSUBS 0.007088f
C833 B.n351 VSUBS 0.007088f
C834 B.n352 VSUBS 0.007088f
C835 B.n353 VSUBS 0.007088f
C836 B.n354 VSUBS 0.007088f
C837 B.n355 VSUBS 0.007088f
C838 B.n356 VSUBS 0.007088f
C839 B.n357 VSUBS 0.007088f
C840 B.n358 VSUBS 0.007088f
C841 B.n359 VSUBS 0.007088f
C842 B.n360 VSUBS 0.007088f
C843 B.n361 VSUBS 0.007088f
C844 B.n362 VSUBS 0.007088f
C845 B.n363 VSUBS 0.007088f
C846 B.n364 VSUBS 0.007088f
C847 B.n365 VSUBS 0.007088f
C848 B.n366 VSUBS 0.007088f
C849 B.n367 VSUBS 0.007088f
C850 B.n368 VSUBS 0.007088f
C851 B.n369 VSUBS 0.007088f
C852 B.n370 VSUBS 0.007088f
C853 B.n371 VSUBS 0.007088f
C854 B.n372 VSUBS 0.007088f
C855 B.n373 VSUBS 0.007088f
C856 B.n374 VSUBS 0.007088f
C857 B.n375 VSUBS 0.007088f
C858 B.n376 VSUBS 0.007088f
C859 B.n377 VSUBS 0.007088f
C860 B.n378 VSUBS 0.007088f
C861 B.n379 VSUBS 0.007088f
C862 B.n380 VSUBS 0.007088f
C863 B.n381 VSUBS 0.007088f
C864 B.n382 VSUBS 0.007088f
C865 B.n383 VSUBS 0.007088f
C866 B.n384 VSUBS 0.007088f
C867 B.n385 VSUBS 0.007088f
C868 B.n386 VSUBS 0.007088f
C869 B.n387 VSUBS 0.007088f
C870 B.n388 VSUBS 0.007088f
C871 B.n389 VSUBS 0.007088f
C872 B.n390 VSUBS 0.007088f
C873 B.n391 VSUBS 0.004899f
C874 B.n392 VSUBS 0.007088f
C875 B.n393 VSUBS 0.007088f
C876 B.n394 VSUBS 0.005733f
C877 B.n395 VSUBS 0.007088f
C878 B.n396 VSUBS 0.007088f
C879 B.n397 VSUBS 0.007088f
C880 B.n398 VSUBS 0.007088f
C881 B.n399 VSUBS 0.007088f
C882 B.n400 VSUBS 0.007088f
C883 B.n401 VSUBS 0.007088f
C884 B.n402 VSUBS 0.007088f
C885 B.n403 VSUBS 0.007088f
C886 B.n404 VSUBS 0.007088f
C887 B.n405 VSUBS 0.007088f
C888 B.n406 VSUBS 0.005733f
C889 B.n407 VSUBS 0.016423f
C890 B.n408 VSUBS 0.004899f
C891 B.n409 VSUBS 0.007088f
C892 B.n410 VSUBS 0.007088f
C893 B.n411 VSUBS 0.007088f
C894 B.n412 VSUBS 0.007088f
C895 B.n413 VSUBS 0.007088f
C896 B.n414 VSUBS 0.007088f
C897 B.n415 VSUBS 0.007088f
C898 B.n416 VSUBS 0.007088f
C899 B.n417 VSUBS 0.007088f
C900 B.n418 VSUBS 0.007088f
C901 B.n419 VSUBS 0.007088f
C902 B.n420 VSUBS 0.007088f
C903 B.n421 VSUBS 0.007088f
C904 B.n422 VSUBS 0.007088f
C905 B.n423 VSUBS 0.007088f
C906 B.n424 VSUBS 0.007088f
C907 B.n425 VSUBS 0.007088f
C908 B.n426 VSUBS 0.007088f
C909 B.n427 VSUBS 0.007088f
C910 B.n428 VSUBS 0.007088f
C911 B.n429 VSUBS 0.007088f
C912 B.n430 VSUBS 0.007088f
C913 B.n431 VSUBS 0.007088f
C914 B.n432 VSUBS 0.007088f
C915 B.n433 VSUBS 0.007088f
C916 B.n434 VSUBS 0.007088f
C917 B.n435 VSUBS 0.007088f
C918 B.n436 VSUBS 0.007088f
C919 B.n437 VSUBS 0.007088f
C920 B.n438 VSUBS 0.007088f
C921 B.n439 VSUBS 0.007088f
C922 B.n440 VSUBS 0.007088f
C923 B.n441 VSUBS 0.007088f
C924 B.n442 VSUBS 0.007088f
C925 B.n443 VSUBS 0.007088f
C926 B.n444 VSUBS 0.007088f
C927 B.n445 VSUBS 0.007088f
C928 B.n446 VSUBS 0.007088f
C929 B.n447 VSUBS 0.007088f
C930 B.n448 VSUBS 0.007088f
C931 B.n449 VSUBS 0.007088f
C932 B.n450 VSUBS 0.007088f
C933 B.n451 VSUBS 0.007088f
C934 B.n452 VSUBS 0.007088f
C935 B.n453 VSUBS 0.007088f
C936 B.n454 VSUBS 0.007088f
C937 B.n455 VSUBS 0.007088f
C938 B.n456 VSUBS 0.007088f
C939 B.n457 VSUBS 0.007088f
C940 B.n458 VSUBS 0.007088f
C941 B.n459 VSUBS 0.007088f
C942 B.n460 VSUBS 0.01712f
C943 B.n461 VSUBS 0.01712f
C944 B.n462 VSUBS 0.015819f
C945 B.n463 VSUBS 0.007088f
C946 B.n464 VSUBS 0.007088f
C947 B.n465 VSUBS 0.007088f
C948 B.n466 VSUBS 0.007088f
C949 B.n467 VSUBS 0.007088f
C950 B.n468 VSUBS 0.007088f
C951 B.n469 VSUBS 0.007088f
C952 B.n470 VSUBS 0.007088f
C953 B.n471 VSUBS 0.007088f
C954 B.n472 VSUBS 0.007088f
C955 B.n473 VSUBS 0.007088f
C956 B.n474 VSUBS 0.007088f
C957 B.n475 VSUBS 0.007088f
C958 B.n476 VSUBS 0.007088f
C959 B.n477 VSUBS 0.007088f
C960 B.n478 VSUBS 0.007088f
C961 B.n479 VSUBS 0.007088f
C962 B.n480 VSUBS 0.007088f
C963 B.n481 VSUBS 0.007088f
C964 B.n482 VSUBS 0.007088f
C965 B.n483 VSUBS 0.007088f
C966 B.n484 VSUBS 0.007088f
C967 B.n485 VSUBS 0.007088f
C968 B.n486 VSUBS 0.007088f
C969 B.n487 VSUBS 0.007088f
C970 B.n488 VSUBS 0.007088f
C971 B.n489 VSUBS 0.007088f
C972 B.n490 VSUBS 0.007088f
C973 B.n491 VSUBS 0.01605f
.ends

