* NGSPICE file created from diff_pair_sample_0956.ext - technology: sky130A

.subckt diff_pair_sample_0956 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.39745 pd=14.86 as=5.6667 ps=29.84 w=14.53 l=1.54
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=0 ps=0 w=14.53 l=1.54
X2 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=2.39745 ps=14.86 w=14.53 l=1.54
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=0 ps=0 w=14.53 l=1.54
X4 VTAIL.t4 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=2.39745 ps=14.86 w=14.53 l=1.54
X5 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.39745 pd=14.86 as=5.6667 ps=29.84 w=14.53 l=1.54
X6 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.39745 pd=14.86 as=5.6667 ps=29.84 w=14.53 l=1.54
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=0 ps=0 w=14.53 l=1.54
X8 VDD2.t1 VN.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.39745 pd=14.86 as=5.6667 ps=29.84 w=14.53 l=1.54
X9 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=2.39745 ps=14.86 w=14.53 l=1.54
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=0 ps=0 w=14.53 l=1.54
X11 VTAIL.t7 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=5.6667 pd=29.84 as=2.39745 ps=14.86 w=14.53 l=1.54
R0 VN.n0 VN.t1 264.325
R1 VN.n1 VN.t2 264.325
R2 VN.n0 VN.t0 264.005
R3 VN.n1 VN.t3 264.005
R4 VN VN.n1 58.1922
R5 VN VN.n0 12.9232
R6 VTAIL.n5 VTAIL.t3 43.9231
R7 VTAIL.n4 VTAIL.t6 43.9231
R8 VTAIL.n3 VTAIL.t7 43.9231
R9 VTAIL.n6 VTAIL.t0 43.923
R10 VTAIL.n7 VTAIL.t5 43.9228
R11 VTAIL.n0 VTAIL.t4 43.9228
R12 VTAIL.n1 VTAIL.t1 43.9228
R13 VTAIL.n2 VTAIL.t2 43.9228
R14 VTAIL.n7 VTAIL.n6 26.5048
R15 VTAIL.n3 VTAIL.n2 26.5048
R16 VTAIL.n4 VTAIL.n3 1.61257
R17 VTAIL.n6 VTAIL.n5 1.61257
R18 VTAIL.n2 VTAIL.n1 1.61257
R19 VTAIL VTAIL.n0 0.864724
R20 VTAIL VTAIL.n7 0.748345
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 100.316
R24 VDD2.n2 VDD2.n1 59.2392
R25 VDD2.n1 VDD2.t0 1.3632
R26 VDD2.n1 VDD2.t1 1.3632
R27 VDD2.n0 VDD2.t2 1.3632
R28 VDD2.n0 VDD2.t3 1.3632
R29 VDD2 VDD2.n2 0.0586897
R30 B.n747 B.n746 585
R31 B.n318 B.n101 585
R32 B.n317 B.n316 585
R33 B.n315 B.n314 585
R34 B.n313 B.n312 585
R35 B.n311 B.n310 585
R36 B.n309 B.n308 585
R37 B.n307 B.n306 585
R38 B.n305 B.n304 585
R39 B.n303 B.n302 585
R40 B.n301 B.n300 585
R41 B.n299 B.n298 585
R42 B.n297 B.n296 585
R43 B.n295 B.n294 585
R44 B.n293 B.n292 585
R45 B.n291 B.n290 585
R46 B.n289 B.n288 585
R47 B.n287 B.n286 585
R48 B.n285 B.n284 585
R49 B.n283 B.n282 585
R50 B.n281 B.n280 585
R51 B.n279 B.n278 585
R52 B.n277 B.n276 585
R53 B.n275 B.n274 585
R54 B.n273 B.n272 585
R55 B.n271 B.n270 585
R56 B.n269 B.n268 585
R57 B.n267 B.n266 585
R58 B.n265 B.n264 585
R59 B.n263 B.n262 585
R60 B.n261 B.n260 585
R61 B.n259 B.n258 585
R62 B.n257 B.n256 585
R63 B.n255 B.n254 585
R64 B.n253 B.n252 585
R65 B.n251 B.n250 585
R66 B.n249 B.n248 585
R67 B.n247 B.n246 585
R68 B.n245 B.n244 585
R69 B.n243 B.n242 585
R70 B.n241 B.n240 585
R71 B.n239 B.n238 585
R72 B.n237 B.n236 585
R73 B.n235 B.n234 585
R74 B.n233 B.n232 585
R75 B.n231 B.n230 585
R76 B.n229 B.n228 585
R77 B.n227 B.n226 585
R78 B.n225 B.n224 585
R79 B.n222 B.n221 585
R80 B.n220 B.n219 585
R81 B.n218 B.n217 585
R82 B.n216 B.n215 585
R83 B.n214 B.n213 585
R84 B.n212 B.n211 585
R85 B.n210 B.n209 585
R86 B.n208 B.n207 585
R87 B.n206 B.n205 585
R88 B.n204 B.n203 585
R89 B.n201 B.n200 585
R90 B.n199 B.n198 585
R91 B.n197 B.n196 585
R92 B.n195 B.n194 585
R93 B.n193 B.n192 585
R94 B.n191 B.n190 585
R95 B.n189 B.n188 585
R96 B.n187 B.n186 585
R97 B.n185 B.n184 585
R98 B.n183 B.n182 585
R99 B.n181 B.n180 585
R100 B.n179 B.n178 585
R101 B.n177 B.n176 585
R102 B.n175 B.n174 585
R103 B.n173 B.n172 585
R104 B.n171 B.n170 585
R105 B.n169 B.n168 585
R106 B.n167 B.n166 585
R107 B.n165 B.n164 585
R108 B.n163 B.n162 585
R109 B.n161 B.n160 585
R110 B.n159 B.n158 585
R111 B.n157 B.n156 585
R112 B.n155 B.n154 585
R113 B.n153 B.n152 585
R114 B.n151 B.n150 585
R115 B.n149 B.n148 585
R116 B.n147 B.n146 585
R117 B.n145 B.n144 585
R118 B.n143 B.n142 585
R119 B.n141 B.n140 585
R120 B.n139 B.n138 585
R121 B.n137 B.n136 585
R122 B.n135 B.n134 585
R123 B.n133 B.n132 585
R124 B.n131 B.n130 585
R125 B.n129 B.n128 585
R126 B.n127 B.n126 585
R127 B.n125 B.n124 585
R128 B.n123 B.n122 585
R129 B.n121 B.n120 585
R130 B.n119 B.n118 585
R131 B.n117 B.n116 585
R132 B.n115 B.n114 585
R133 B.n113 B.n112 585
R134 B.n111 B.n110 585
R135 B.n109 B.n108 585
R136 B.n107 B.n106 585
R137 B.n46 B.n45 585
R138 B.n745 B.n47 585
R139 B.n750 B.n47 585
R140 B.n744 B.n743 585
R141 B.n743 B.n43 585
R142 B.n742 B.n42 585
R143 B.n756 B.n42 585
R144 B.n741 B.n41 585
R145 B.n757 B.n41 585
R146 B.n740 B.n40 585
R147 B.n758 B.n40 585
R148 B.n739 B.n738 585
R149 B.n738 B.n39 585
R150 B.n737 B.n35 585
R151 B.n764 B.n35 585
R152 B.n736 B.n34 585
R153 B.n765 B.n34 585
R154 B.n735 B.n33 585
R155 B.n766 B.n33 585
R156 B.n734 B.n733 585
R157 B.n733 B.n29 585
R158 B.n732 B.n28 585
R159 B.n772 B.n28 585
R160 B.n731 B.n27 585
R161 B.n773 B.n27 585
R162 B.n730 B.n26 585
R163 B.n774 B.n26 585
R164 B.n729 B.n728 585
R165 B.n728 B.n22 585
R166 B.n727 B.n21 585
R167 B.n780 B.n21 585
R168 B.n726 B.n20 585
R169 B.n781 B.n20 585
R170 B.n725 B.n19 585
R171 B.n782 B.n19 585
R172 B.n724 B.n723 585
R173 B.n723 B.n15 585
R174 B.n722 B.n14 585
R175 B.n788 B.n14 585
R176 B.n721 B.n13 585
R177 B.n789 B.n13 585
R178 B.n720 B.n12 585
R179 B.n790 B.n12 585
R180 B.n719 B.n718 585
R181 B.n718 B.n717 585
R182 B.n716 B.n715 585
R183 B.n716 B.n8 585
R184 B.n714 B.n7 585
R185 B.n797 B.n7 585
R186 B.n713 B.n6 585
R187 B.n798 B.n6 585
R188 B.n712 B.n5 585
R189 B.n799 B.n5 585
R190 B.n711 B.n710 585
R191 B.n710 B.n4 585
R192 B.n709 B.n319 585
R193 B.n709 B.n708 585
R194 B.n699 B.n320 585
R195 B.n321 B.n320 585
R196 B.n701 B.n700 585
R197 B.n702 B.n701 585
R198 B.n698 B.n326 585
R199 B.n326 B.n325 585
R200 B.n697 B.n696 585
R201 B.n696 B.n695 585
R202 B.n328 B.n327 585
R203 B.n329 B.n328 585
R204 B.n688 B.n687 585
R205 B.n689 B.n688 585
R206 B.n686 B.n334 585
R207 B.n334 B.n333 585
R208 B.n685 B.n684 585
R209 B.n684 B.n683 585
R210 B.n336 B.n335 585
R211 B.n337 B.n336 585
R212 B.n676 B.n675 585
R213 B.n677 B.n676 585
R214 B.n674 B.n342 585
R215 B.n342 B.n341 585
R216 B.n673 B.n672 585
R217 B.n672 B.n671 585
R218 B.n344 B.n343 585
R219 B.n345 B.n344 585
R220 B.n664 B.n663 585
R221 B.n665 B.n664 585
R222 B.n662 B.n350 585
R223 B.n350 B.n349 585
R224 B.n661 B.n660 585
R225 B.n660 B.n659 585
R226 B.n352 B.n351 585
R227 B.n652 B.n352 585
R228 B.n651 B.n650 585
R229 B.n653 B.n651 585
R230 B.n649 B.n357 585
R231 B.n357 B.n356 585
R232 B.n648 B.n647 585
R233 B.n647 B.n646 585
R234 B.n359 B.n358 585
R235 B.n360 B.n359 585
R236 B.n639 B.n638 585
R237 B.n640 B.n639 585
R238 B.n363 B.n362 585
R239 B.n426 B.n425 585
R240 B.n427 B.n423 585
R241 B.n423 B.n364 585
R242 B.n429 B.n428 585
R243 B.n431 B.n422 585
R244 B.n434 B.n433 585
R245 B.n435 B.n421 585
R246 B.n437 B.n436 585
R247 B.n439 B.n420 585
R248 B.n442 B.n441 585
R249 B.n443 B.n419 585
R250 B.n445 B.n444 585
R251 B.n447 B.n418 585
R252 B.n450 B.n449 585
R253 B.n451 B.n417 585
R254 B.n453 B.n452 585
R255 B.n455 B.n416 585
R256 B.n458 B.n457 585
R257 B.n459 B.n415 585
R258 B.n461 B.n460 585
R259 B.n463 B.n414 585
R260 B.n466 B.n465 585
R261 B.n467 B.n413 585
R262 B.n469 B.n468 585
R263 B.n471 B.n412 585
R264 B.n474 B.n473 585
R265 B.n475 B.n411 585
R266 B.n477 B.n476 585
R267 B.n479 B.n410 585
R268 B.n482 B.n481 585
R269 B.n483 B.n409 585
R270 B.n485 B.n484 585
R271 B.n487 B.n408 585
R272 B.n490 B.n489 585
R273 B.n491 B.n407 585
R274 B.n493 B.n492 585
R275 B.n495 B.n406 585
R276 B.n498 B.n497 585
R277 B.n499 B.n405 585
R278 B.n501 B.n500 585
R279 B.n503 B.n404 585
R280 B.n506 B.n505 585
R281 B.n507 B.n403 585
R282 B.n509 B.n508 585
R283 B.n511 B.n402 585
R284 B.n514 B.n513 585
R285 B.n515 B.n401 585
R286 B.n517 B.n516 585
R287 B.n519 B.n400 585
R288 B.n522 B.n521 585
R289 B.n523 B.n396 585
R290 B.n525 B.n524 585
R291 B.n527 B.n395 585
R292 B.n530 B.n529 585
R293 B.n531 B.n394 585
R294 B.n533 B.n532 585
R295 B.n535 B.n393 585
R296 B.n538 B.n537 585
R297 B.n539 B.n390 585
R298 B.n542 B.n541 585
R299 B.n544 B.n389 585
R300 B.n547 B.n546 585
R301 B.n548 B.n388 585
R302 B.n550 B.n549 585
R303 B.n552 B.n387 585
R304 B.n555 B.n554 585
R305 B.n556 B.n386 585
R306 B.n558 B.n557 585
R307 B.n560 B.n385 585
R308 B.n563 B.n562 585
R309 B.n564 B.n384 585
R310 B.n566 B.n565 585
R311 B.n568 B.n383 585
R312 B.n571 B.n570 585
R313 B.n572 B.n382 585
R314 B.n574 B.n573 585
R315 B.n576 B.n381 585
R316 B.n579 B.n578 585
R317 B.n580 B.n380 585
R318 B.n582 B.n581 585
R319 B.n584 B.n379 585
R320 B.n587 B.n586 585
R321 B.n588 B.n378 585
R322 B.n590 B.n589 585
R323 B.n592 B.n377 585
R324 B.n595 B.n594 585
R325 B.n596 B.n376 585
R326 B.n598 B.n597 585
R327 B.n600 B.n375 585
R328 B.n603 B.n602 585
R329 B.n604 B.n374 585
R330 B.n606 B.n605 585
R331 B.n608 B.n373 585
R332 B.n611 B.n610 585
R333 B.n612 B.n372 585
R334 B.n614 B.n613 585
R335 B.n616 B.n371 585
R336 B.n619 B.n618 585
R337 B.n620 B.n370 585
R338 B.n622 B.n621 585
R339 B.n624 B.n369 585
R340 B.n627 B.n626 585
R341 B.n628 B.n368 585
R342 B.n630 B.n629 585
R343 B.n632 B.n367 585
R344 B.n633 B.n366 585
R345 B.n636 B.n635 585
R346 B.n637 B.n365 585
R347 B.n365 B.n364 585
R348 B.n642 B.n641 585
R349 B.n641 B.n640 585
R350 B.n643 B.n361 585
R351 B.n361 B.n360 585
R352 B.n645 B.n644 585
R353 B.n646 B.n645 585
R354 B.n355 B.n354 585
R355 B.n356 B.n355 585
R356 B.n655 B.n654 585
R357 B.n654 B.n653 585
R358 B.n656 B.n353 585
R359 B.n652 B.n353 585
R360 B.n658 B.n657 585
R361 B.n659 B.n658 585
R362 B.n348 B.n347 585
R363 B.n349 B.n348 585
R364 B.n667 B.n666 585
R365 B.n666 B.n665 585
R366 B.n668 B.n346 585
R367 B.n346 B.n345 585
R368 B.n670 B.n669 585
R369 B.n671 B.n670 585
R370 B.n340 B.n339 585
R371 B.n341 B.n340 585
R372 B.n679 B.n678 585
R373 B.n678 B.n677 585
R374 B.n680 B.n338 585
R375 B.n338 B.n337 585
R376 B.n682 B.n681 585
R377 B.n683 B.n682 585
R378 B.n332 B.n331 585
R379 B.n333 B.n332 585
R380 B.n691 B.n690 585
R381 B.n690 B.n689 585
R382 B.n692 B.n330 585
R383 B.n330 B.n329 585
R384 B.n694 B.n693 585
R385 B.n695 B.n694 585
R386 B.n324 B.n323 585
R387 B.n325 B.n324 585
R388 B.n704 B.n703 585
R389 B.n703 B.n702 585
R390 B.n705 B.n322 585
R391 B.n322 B.n321 585
R392 B.n707 B.n706 585
R393 B.n708 B.n707 585
R394 B.n3 B.n0 585
R395 B.n4 B.n3 585
R396 B.n796 B.n1 585
R397 B.n797 B.n796 585
R398 B.n795 B.n794 585
R399 B.n795 B.n8 585
R400 B.n793 B.n9 585
R401 B.n717 B.n9 585
R402 B.n792 B.n791 585
R403 B.n791 B.n790 585
R404 B.n11 B.n10 585
R405 B.n789 B.n11 585
R406 B.n787 B.n786 585
R407 B.n788 B.n787 585
R408 B.n785 B.n16 585
R409 B.n16 B.n15 585
R410 B.n784 B.n783 585
R411 B.n783 B.n782 585
R412 B.n18 B.n17 585
R413 B.n781 B.n18 585
R414 B.n779 B.n778 585
R415 B.n780 B.n779 585
R416 B.n777 B.n23 585
R417 B.n23 B.n22 585
R418 B.n776 B.n775 585
R419 B.n775 B.n774 585
R420 B.n25 B.n24 585
R421 B.n773 B.n25 585
R422 B.n771 B.n770 585
R423 B.n772 B.n771 585
R424 B.n769 B.n30 585
R425 B.n30 B.n29 585
R426 B.n768 B.n767 585
R427 B.n767 B.n766 585
R428 B.n32 B.n31 585
R429 B.n765 B.n32 585
R430 B.n763 B.n762 585
R431 B.n764 B.n763 585
R432 B.n761 B.n36 585
R433 B.n39 B.n36 585
R434 B.n760 B.n759 585
R435 B.n759 B.n758 585
R436 B.n38 B.n37 585
R437 B.n757 B.n38 585
R438 B.n755 B.n754 585
R439 B.n756 B.n755 585
R440 B.n753 B.n44 585
R441 B.n44 B.n43 585
R442 B.n752 B.n751 585
R443 B.n751 B.n750 585
R444 B.n800 B.n799 585
R445 B.n798 B.n2 585
R446 B.n751 B.n46 492.5
R447 B.n747 B.n47 492.5
R448 B.n639 B.n365 492.5
R449 B.n641 B.n363 492.5
R450 B.n104 B.t15 432.971
R451 B.n102 B.t11 432.971
R452 B.n391 B.t8 432.971
R453 B.n397 B.t4 432.971
R454 B.n749 B.n748 256.663
R455 B.n749 B.n100 256.663
R456 B.n749 B.n99 256.663
R457 B.n749 B.n98 256.663
R458 B.n749 B.n97 256.663
R459 B.n749 B.n96 256.663
R460 B.n749 B.n95 256.663
R461 B.n749 B.n94 256.663
R462 B.n749 B.n93 256.663
R463 B.n749 B.n92 256.663
R464 B.n749 B.n91 256.663
R465 B.n749 B.n90 256.663
R466 B.n749 B.n89 256.663
R467 B.n749 B.n88 256.663
R468 B.n749 B.n87 256.663
R469 B.n749 B.n86 256.663
R470 B.n749 B.n85 256.663
R471 B.n749 B.n84 256.663
R472 B.n749 B.n83 256.663
R473 B.n749 B.n82 256.663
R474 B.n749 B.n81 256.663
R475 B.n749 B.n80 256.663
R476 B.n749 B.n79 256.663
R477 B.n749 B.n78 256.663
R478 B.n749 B.n77 256.663
R479 B.n749 B.n76 256.663
R480 B.n749 B.n75 256.663
R481 B.n749 B.n74 256.663
R482 B.n749 B.n73 256.663
R483 B.n749 B.n72 256.663
R484 B.n749 B.n71 256.663
R485 B.n749 B.n70 256.663
R486 B.n749 B.n69 256.663
R487 B.n749 B.n68 256.663
R488 B.n749 B.n67 256.663
R489 B.n749 B.n66 256.663
R490 B.n749 B.n65 256.663
R491 B.n749 B.n64 256.663
R492 B.n749 B.n63 256.663
R493 B.n749 B.n62 256.663
R494 B.n749 B.n61 256.663
R495 B.n749 B.n60 256.663
R496 B.n749 B.n59 256.663
R497 B.n749 B.n58 256.663
R498 B.n749 B.n57 256.663
R499 B.n749 B.n56 256.663
R500 B.n749 B.n55 256.663
R501 B.n749 B.n54 256.663
R502 B.n749 B.n53 256.663
R503 B.n749 B.n52 256.663
R504 B.n749 B.n51 256.663
R505 B.n749 B.n50 256.663
R506 B.n749 B.n49 256.663
R507 B.n749 B.n48 256.663
R508 B.n424 B.n364 256.663
R509 B.n430 B.n364 256.663
R510 B.n432 B.n364 256.663
R511 B.n438 B.n364 256.663
R512 B.n440 B.n364 256.663
R513 B.n446 B.n364 256.663
R514 B.n448 B.n364 256.663
R515 B.n454 B.n364 256.663
R516 B.n456 B.n364 256.663
R517 B.n462 B.n364 256.663
R518 B.n464 B.n364 256.663
R519 B.n470 B.n364 256.663
R520 B.n472 B.n364 256.663
R521 B.n478 B.n364 256.663
R522 B.n480 B.n364 256.663
R523 B.n486 B.n364 256.663
R524 B.n488 B.n364 256.663
R525 B.n494 B.n364 256.663
R526 B.n496 B.n364 256.663
R527 B.n502 B.n364 256.663
R528 B.n504 B.n364 256.663
R529 B.n510 B.n364 256.663
R530 B.n512 B.n364 256.663
R531 B.n518 B.n364 256.663
R532 B.n520 B.n364 256.663
R533 B.n526 B.n364 256.663
R534 B.n528 B.n364 256.663
R535 B.n534 B.n364 256.663
R536 B.n536 B.n364 256.663
R537 B.n543 B.n364 256.663
R538 B.n545 B.n364 256.663
R539 B.n551 B.n364 256.663
R540 B.n553 B.n364 256.663
R541 B.n559 B.n364 256.663
R542 B.n561 B.n364 256.663
R543 B.n567 B.n364 256.663
R544 B.n569 B.n364 256.663
R545 B.n575 B.n364 256.663
R546 B.n577 B.n364 256.663
R547 B.n583 B.n364 256.663
R548 B.n585 B.n364 256.663
R549 B.n591 B.n364 256.663
R550 B.n593 B.n364 256.663
R551 B.n599 B.n364 256.663
R552 B.n601 B.n364 256.663
R553 B.n607 B.n364 256.663
R554 B.n609 B.n364 256.663
R555 B.n615 B.n364 256.663
R556 B.n617 B.n364 256.663
R557 B.n623 B.n364 256.663
R558 B.n625 B.n364 256.663
R559 B.n631 B.n364 256.663
R560 B.n634 B.n364 256.663
R561 B.n802 B.n801 256.663
R562 B.n108 B.n107 163.367
R563 B.n112 B.n111 163.367
R564 B.n116 B.n115 163.367
R565 B.n120 B.n119 163.367
R566 B.n124 B.n123 163.367
R567 B.n128 B.n127 163.367
R568 B.n132 B.n131 163.367
R569 B.n136 B.n135 163.367
R570 B.n140 B.n139 163.367
R571 B.n144 B.n143 163.367
R572 B.n148 B.n147 163.367
R573 B.n152 B.n151 163.367
R574 B.n156 B.n155 163.367
R575 B.n160 B.n159 163.367
R576 B.n164 B.n163 163.367
R577 B.n168 B.n167 163.367
R578 B.n172 B.n171 163.367
R579 B.n176 B.n175 163.367
R580 B.n180 B.n179 163.367
R581 B.n184 B.n183 163.367
R582 B.n188 B.n187 163.367
R583 B.n192 B.n191 163.367
R584 B.n196 B.n195 163.367
R585 B.n200 B.n199 163.367
R586 B.n205 B.n204 163.367
R587 B.n209 B.n208 163.367
R588 B.n213 B.n212 163.367
R589 B.n217 B.n216 163.367
R590 B.n221 B.n220 163.367
R591 B.n226 B.n225 163.367
R592 B.n230 B.n229 163.367
R593 B.n234 B.n233 163.367
R594 B.n238 B.n237 163.367
R595 B.n242 B.n241 163.367
R596 B.n246 B.n245 163.367
R597 B.n250 B.n249 163.367
R598 B.n254 B.n253 163.367
R599 B.n258 B.n257 163.367
R600 B.n262 B.n261 163.367
R601 B.n266 B.n265 163.367
R602 B.n270 B.n269 163.367
R603 B.n274 B.n273 163.367
R604 B.n278 B.n277 163.367
R605 B.n282 B.n281 163.367
R606 B.n286 B.n285 163.367
R607 B.n290 B.n289 163.367
R608 B.n294 B.n293 163.367
R609 B.n298 B.n297 163.367
R610 B.n302 B.n301 163.367
R611 B.n306 B.n305 163.367
R612 B.n310 B.n309 163.367
R613 B.n314 B.n313 163.367
R614 B.n316 B.n101 163.367
R615 B.n639 B.n359 163.367
R616 B.n647 B.n359 163.367
R617 B.n647 B.n357 163.367
R618 B.n651 B.n357 163.367
R619 B.n651 B.n352 163.367
R620 B.n660 B.n352 163.367
R621 B.n660 B.n350 163.367
R622 B.n664 B.n350 163.367
R623 B.n664 B.n344 163.367
R624 B.n672 B.n344 163.367
R625 B.n672 B.n342 163.367
R626 B.n676 B.n342 163.367
R627 B.n676 B.n336 163.367
R628 B.n684 B.n336 163.367
R629 B.n684 B.n334 163.367
R630 B.n688 B.n334 163.367
R631 B.n688 B.n328 163.367
R632 B.n696 B.n328 163.367
R633 B.n696 B.n326 163.367
R634 B.n701 B.n326 163.367
R635 B.n701 B.n320 163.367
R636 B.n709 B.n320 163.367
R637 B.n710 B.n709 163.367
R638 B.n710 B.n5 163.367
R639 B.n6 B.n5 163.367
R640 B.n7 B.n6 163.367
R641 B.n716 B.n7 163.367
R642 B.n718 B.n716 163.367
R643 B.n718 B.n12 163.367
R644 B.n13 B.n12 163.367
R645 B.n14 B.n13 163.367
R646 B.n723 B.n14 163.367
R647 B.n723 B.n19 163.367
R648 B.n20 B.n19 163.367
R649 B.n21 B.n20 163.367
R650 B.n728 B.n21 163.367
R651 B.n728 B.n26 163.367
R652 B.n27 B.n26 163.367
R653 B.n28 B.n27 163.367
R654 B.n733 B.n28 163.367
R655 B.n733 B.n33 163.367
R656 B.n34 B.n33 163.367
R657 B.n35 B.n34 163.367
R658 B.n738 B.n35 163.367
R659 B.n738 B.n40 163.367
R660 B.n41 B.n40 163.367
R661 B.n42 B.n41 163.367
R662 B.n743 B.n42 163.367
R663 B.n743 B.n47 163.367
R664 B.n425 B.n423 163.367
R665 B.n429 B.n423 163.367
R666 B.n433 B.n431 163.367
R667 B.n437 B.n421 163.367
R668 B.n441 B.n439 163.367
R669 B.n445 B.n419 163.367
R670 B.n449 B.n447 163.367
R671 B.n453 B.n417 163.367
R672 B.n457 B.n455 163.367
R673 B.n461 B.n415 163.367
R674 B.n465 B.n463 163.367
R675 B.n469 B.n413 163.367
R676 B.n473 B.n471 163.367
R677 B.n477 B.n411 163.367
R678 B.n481 B.n479 163.367
R679 B.n485 B.n409 163.367
R680 B.n489 B.n487 163.367
R681 B.n493 B.n407 163.367
R682 B.n497 B.n495 163.367
R683 B.n501 B.n405 163.367
R684 B.n505 B.n503 163.367
R685 B.n509 B.n403 163.367
R686 B.n513 B.n511 163.367
R687 B.n517 B.n401 163.367
R688 B.n521 B.n519 163.367
R689 B.n525 B.n396 163.367
R690 B.n529 B.n527 163.367
R691 B.n533 B.n394 163.367
R692 B.n537 B.n535 163.367
R693 B.n542 B.n390 163.367
R694 B.n546 B.n544 163.367
R695 B.n550 B.n388 163.367
R696 B.n554 B.n552 163.367
R697 B.n558 B.n386 163.367
R698 B.n562 B.n560 163.367
R699 B.n566 B.n384 163.367
R700 B.n570 B.n568 163.367
R701 B.n574 B.n382 163.367
R702 B.n578 B.n576 163.367
R703 B.n582 B.n380 163.367
R704 B.n586 B.n584 163.367
R705 B.n590 B.n378 163.367
R706 B.n594 B.n592 163.367
R707 B.n598 B.n376 163.367
R708 B.n602 B.n600 163.367
R709 B.n606 B.n374 163.367
R710 B.n610 B.n608 163.367
R711 B.n614 B.n372 163.367
R712 B.n618 B.n616 163.367
R713 B.n622 B.n370 163.367
R714 B.n626 B.n624 163.367
R715 B.n630 B.n368 163.367
R716 B.n633 B.n632 163.367
R717 B.n635 B.n365 163.367
R718 B.n641 B.n361 163.367
R719 B.n645 B.n361 163.367
R720 B.n645 B.n355 163.367
R721 B.n654 B.n355 163.367
R722 B.n654 B.n353 163.367
R723 B.n658 B.n353 163.367
R724 B.n658 B.n348 163.367
R725 B.n666 B.n348 163.367
R726 B.n666 B.n346 163.367
R727 B.n670 B.n346 163.367
R728 B.n670 B.n340 163.367
R729 B.n678 B.n340 163.367
R730 B.n678 B.n338 163.367
R731 B.n682 B.n338 163.367
R732 B.n682 B.n332 163.367
R733 B.n690 B.n332 163.367
R734 B.n690 B.n330 163.367
R735 B.n694 B.n330 163.367
R736 B.n694 B.n324 163.367
R737 B.n703 B.n324 163.367
R738 B.n703 B.n322 163.367
R739 B.n707 B.n322 163.367
R740 B.n707 B.n3 163.367
R741 B.n800 B.n3 163.367
R742 B.n796 B.n2 163.367
R743 B.n796 B.n795 163.367
R744 B.n795 B.n9 163.367
R745 B.n791 B.n9 163.367
R746 B.n791 B.n11 163.367
R747 B.n787 B.n11 163.367
R748 B.n787 B.n16 163.367
R749 B.n783 B.n16 163.367
R750 B.n783 B.n18 163.367
R751 B.n779 B.n18 163.367
R752 B.n779 B.n23 163.367
R753 B.n775 B.n23 163.367
R754 B.n775 B.n25 163.367
R755 B.n771 B.n25 163.367
R756 B.n771 B.n30 163.367
R757 B.n767 B.n30 163.367
R758 B.n767 B.n32 163.367
R759 B.n763 B.n32 163.367
R760 B.n763 B.n36 163.367
R761 B.n759 B.n36 163.367
R762 B.n759 B.n38 163.367
R763 B.n755 B.n38 163.367
R764 B.n755 B.n44 163.367
R765 B.n751 B.n44 163.367
R766 B.n102 B.t13 108.621
R767 B.n391 B.t10 108.621
R768 B.n104 B.t16 108.603
R769 B.n397 B.t7 108.603
R770 B.n640 B.n364 72.7599
R771 B.n750 B.n749 72.7599
R772 B.n103 B.t14 72.3546
R773 B.n392 B.t9 72.3546
R774 B.n105 B.t17 72.3358
R775 B.n398 B.t6 72.3358
R776 B.n48 B.n46 71.676
R777 B.n108 B.n49 71.676
R778 B.n112 B.n50 71.676
R779 B.n116 B.n51 71.676
R780 B.n120 B.n52 71.676
R781 B.n124 B.n53 71.676
R782 B.n128 B.n54 71.676
R783 B.n132 B.n55 71.676
R784 B.n136 B.n56 71.676
R785 B.n140 B.n57 71.676
R786 B.n144 B.n58 71.676
R787 B.n148 B.n59 71.676
R788 B.n152 B.n60 71.676
R789 B.n156 B.n61 71.676
R790 B.n160 B.n62 71.676
R791 B.n164 B.n63 71.676
R792 B.n168 B.n64 71.676
R793 B.n172 B.n65 71.676
R794 B.n176 B.n66 71.676
R795 B.n180 B.n67 71.676
R796 B.n184 B.n68 71.676
R797 B.n188 B.n69 71.676
R798 B.n192 B.n70 71.676
R799 B.n196 B.n71 71.676
R800 B.n200 B.n72 71.676
R801 B.n205 B.n73 71.676
R802 B.n209 B.n74 71.676
R803 B.n213 B.n75 71.676
R804 B.n217 B.n76 71.676
R805 B.n221 B.n77 71.676
R806 B.n226 B.n78 71.676
R807 B.n230 B.n79 71.676
R808 B.n234 B.n80 71.676
R809 B.n238 B.n81 71.676
R810 B.n242 B.n82 71.676
R811 B.n246 B.n83 71.676
R812 B.n250 B.n84 71.676
R813 B.n254 B.n85 71.676
R814 B.n258 B.n86 71.676
R815 B.n262 B.n87 71.676
R816 B.n266 B.n88 71.676
R817 B.n270 B.n89 71.676
R818 B.n274 B.n90 71.676
R819 B.n278 B.n91 71.676
R820 B.n282 B.n92 71.676
R821 B.n286 B.n93 71.676
R822 B.n290 B.n94 71.676
R823 B.n294 B.n95 71.676
R824 B.n298 B.n96 71.676
R825 B.n302 B.n97 71.676
R826 B.n306 B.n98 71.676
R827 B.n310 B.n99 71.676
R828 B.n314 B.n100 71.676
R829 B.n748 B.n101 71.676
R830 B.n748 B.n747 71.676
R831 B.n316 B.n100 71.676
R832 B.n313 B.n99 71.676
R833 B.n309 B.n98 71.676
R834 B.n305 B.n97 71.676
R835 B.n301 B.n96 71.676
R836 B.n297 B.n95 71.676
R837 B.n293 B.n94 71.676
R838 B.n289 B.n93 71.676
R839 B.n285 B.n92 71.676
R840 B.n281 B.n91 71.676
R841 B.n277 B.n90 71.676
R842 B.n273 B.n89 71.676
R843 B.n269 B.n88 71.676
R844 B.n265 B.n87 71.676
R845 B.n261 B.n86 71.676
R846 B.n257 B.n85 71.676
R847 B.n253 B.n84 71.676
R848 B.n249 B.n83 71.676
R849 B.n245 B.n82 71.676
R850 B.n241 B.n81 71.676
R851 B.n237 B.n80 71.676
R852 B.n233 B.n79 71.676
R853 B.n229 B.n78 71.676
R854 B.n225 B.n77 71.676
R855 B.n220 B.n76 71.676
R856 B.n216 B.n75 71.676
R857 B.n212 B.n74 71.676
R858 B.n208 B.n73 71.676
R859 B.n204 B.n72 71.676
R860 B.n199 B.n71 71.676
R861 B.n195 B.n70 71.676
R862 B.n191 B.n69 71.676
R863 B.n187 B.n68 71.676
R864 B.n183 B.n67 71.676
R865 B.n179 B.n66 71.676
R866 B.n175 B.n65 71.676
R867 B.n171 B.n64 71.676
R868 B.n167 B.n63 71.676
R869 B.n163 B.n62 71.676
R870 B.n159 B.n61 71.676
R871 B.n155 B.n60 71.676
R872 B.n151 B.n59 71.676
R873 B.n147 B.n58 71.676
R874 B.n143 B.n57 71.676
R875 B.n139 B.n56 71.676
R876 B.n135 B.n55 71.676
R877 B.n131 B.n54 71.676
R878 B.n127 B.n53 71.676
R879 B.n123 B.n52 71.676
R880 B.n119 B.n51 71.676
R881 B.n115 B.n50 71.676
R882 B.n111 B.n49 71.676
R883 B.n107 B.n48 71.676
R884 B.n424 B.n363 71.676
R885 B.n430 B.n429 71.676
R886 B.n433 B.n432 71.676
R887 B.n438 B.n437 71.676
R888 B.n441 B.n440 71.676
R889 B.n446 B.n445 71.676
R890 B.n449 B.n448 71.676
R891 B.n454 B.n453 71.676
R892 B.n457 B.n456 71.676
R893 B.n462 B.n461 71.676
R894 B.n465 B.n464 71.676
R895 B.n470 B.n469 71.676
R896 B.n473 B.n472 71.676
R897 B.n478 B.n477 71.676
R898 B.n481 B.n480 71.676
R899 B.n486 B.n485 71.676
R900 B.n489 B.n488 71.676
R901 B.n494 B.n493 71.676
R902 B.n497 B.n496 71.676
R903 B.n502 B.n501 71.676
R904 B.n505 B.n504 71.676
R905 B.n510 B.n509 71.676
R906 B.n513 B.n512 71.676
R907 B.n518 B.n517 71.676
R908 B.n521 B.n520 71.676
R909 B.n526 B.n525 71.676
R910 B.n529 B.n528 71.676
R911 B.n534 B.n533 71.676
R912 B.n537 B.n536 71.676
R913 B.n543 B.n542 71.676
R914 B.n546 B.n545 71.676
R915 B.n551 B.n550 71.676
R916 B.n554 B.n553 71.676
R917 B.n559 B.n558 71.676
R918 B.n562 B.n561 71.676
R919 B.n567 B.n566 71.676
R920 B.n570 B.n569 71.676
R921 B.n575 B.n574 71.676
R922 B.n578 B.n577 71.676
R923 B.n583 B.n582 71.676
R924 B.n586 B.n585 71.676
R925 B.n591 B.n590 71.676
R926 B.n594 B.n593 71.676
R927 B.n599 B.n598 71.676
R928 B.n602 B.n601 71.676
R929 B.n607 B.n606 71.676
R930 B.n610 B.n609 71.676
R931 B.n615 B.n614 71.676
R932 B.n618 B.n617 71.676
R933 B.n623 B.n622 71.676
R934 B.n626 B.n625 71.676
R935 B.n631 B.n630 71.676
R936 B.n634 B.n633 71.676
R937 B.n425 B.n424 71.676
R938 B.n431 B.n430 71.676
R939 B.n432 B.n421 71.676
R940 B.n439 B.n438 71.676
R941 B.n440 B.n419 71.676
R942 B.n447 B.n446 71.676
R943 B.n448 B.n417 71.676
R944 B.n455 B.n454 71.676
R945 B.n456 B.n415 71.676
R946 B.n463 B.n462 71.676
R947 B.n464 B.n413 71.676
R948 B.n471 B.n470 71.676
R949 B.n472 B.n411 71.676
R950 B.n479 B.n478 71.676
R951 B.n480 B.n409 71.676
R952 B.n487 B.n486 71.676
R953 B.n488 B.n407 71.676
R954 B.n495 B.n494 71.676
R955 B.n496 B.n405 71.676
R956 B.n503 B.n502 71.676
R957 B.n504 B.n403 71.676
R958 B.n511 B.n510 71.676
R959 B.n512 B.n401 71.676
R960 B.n519 B.n518 71.676
R961 B.n520 B.n396 71.676
R962 B.n527 B.n526 71.676
R963 B.n528 B.n394 71.676
R964 B.n535 B.n534 71.676
R965 B.n536 B.n390 71.676
R966 B.n544 B.n543 71.676
R967 B.n545 B.n388 71.676
R968 B.n552 B.n551 71.676
R969 B.n553 B.n386 71.676
R970 B.n560 B.n559 71.676
R971 B.n561 B.n384 71.676
R972 B.n568 B.n567 71.676
R973 B.n569 B.n382 71.676
R974 B.n576 B.n575 71.676
R975 B.n577 B.n380 71.676
R976 B.n584 B.n583 71.676
R977 B.n585 B.n378 71.676
R978 B.n592 B.n591 71.676
R979 B.n593 B.n376 71.676
R980 B.n600 B.n599 71.676
R981 B.n601 B.n374 71.676
R982 B.n608 B.n607 71.676
R983 B.n609 B.n372 71.676
R984 B.n616 B.n615 71.676
R985 B.n617 B.n370 71.676
R986 B.n624 B.n623 71.676
R987 B.n625 B.n368 71.676
R988 B.n632 B.n631 71.676
R989 B.n635 B.n634 71.676
R990 B.n801 B.n800 71.676
R991 B.n801 B.n2 71.676
R992 B.n202 B.n105 59.5399
R993 B.n223 B.n103 59.5399
R994 B.n540 B.n392 59.5399
R995 B.n399 B.n398 59.5399
R996 B.n640 B.n360 37.7687
R997 B.n646 B.n360 37.7687
R998 B.n646 B.n356 37.7687
R999 B.n653 B.n356 37.7687
R1000 B.n653 B.n652 37.7687
R1001 B.n659 B.n349 37.7687
R1002 B.n665 B.n349 37.7687
R1003 B.n665 B.n345 37.7687
R1004 B.n671 B.n345 37.7687
R1005 B.n671 B.n341 37.7687
R1006 B.n677 B.n341 37.7687
R1007 B.n677 B.n337 37.7687
R1008 B.n683 B.n337 37.7687
R1009 B.n689 B.n333 37.7687
R1010 B.n689 B.n329 37.7687
R1011 B.n695 B.n329 37.7687
R1012 B.n695 B.n325 37.7687
R1013 B.n702 B.n325 37.7687
R1014 B.n708 B.n321 37.7687
R1015 B.n708 B.n4 37.7687
R1016 B.n799 B.n4 37.7687
R1017 B.n799 B.n798 37.7687
R1018 B.n798 B.n797 37.7687
R1019 B.n797 B.n8 37.7687
R1020 B.n717 B.n8 37.7687
R1021 B.n790 B.n789 37.7687
R1022 B.n789 B.n788 37.7687
R1023 B.n788 B.n15 37.7687
R1024 B.n782 B.n15 37.7687
R1025 B.n782 B.n781 37.7687
R1026 B.n780 B.n22 37.7687
R1027 B.n774 B.n22 37.7687
R1028 B.n774 B.n773 37.7687
R1029 B.n773 B.n772 37.7687
R1030 B.n772 B.n29 37.7687
R1031 B.n766 B.n29 37.7687
R1032 B.n766 B.n765 37.7687
R1033 B.n765 B.n764 37.7687
R1034 B.n758 B.n39 37.7687
R1035 B.n758 B.n757 37.7687
R1036 B.n757 B.n756 37.7687
R1037 B.n756 B.n43 37.7687
R1038 B.n750 B.n43 37.7687
R1039 B.n105 B.n104 36.2672
R1040 B.n103 B.n102 36.2672
R1041 B.n392 B.n391 36.2672
R1042 B.n398 B.n397 36.2672
R1043 B.n652 B.t5 35.5471
R1044 B.n39 B.t12 35.5471
R1045 B.t1 B.n321 32.2146
R1046 B.n717 B.t3 32.2146
R1047 B.n642 B.n362 32.0005
R1048 B.n638 B.n637 32.0005
R1049 B.n746 B.n745 32.0005
R1050 B.n752 B.n45 32.0005
R1051 B.n683 B.t2 24.4388
R1052 B.t0 B.n780 24.4388
R1053 B B.n802 18.0485
R1054 B.t2 B.n333 13.3305
R1055 B.n781 B.t0 13.3305
R1056 B.n643 B.n642 10.6151
R1057 B.n644 B.n643 10.6151
R1058 B.n644 B.n354 10.6151
R1059 B.n655 B.n354 10.6151
R1060 B.n656 B.n655 10.6151
R1061 B.n657 B.n656 10.6151
R1062 B.n657 B.n347 10.6151
R1063 B.n667 B.n347 10.6151
R1064 B.n668 B.n667 10.6151
R1065 B.n669 B.n668 10.6151
R1066 B.n669 B.n339 10.6151
R1067 B.n679 B.n339 10.6151
R1068 B.n680 B.n679 10.6151
R1069 B.n681 B.n680 10.6151
R1070 B.n681 B.n331 10.6151
R1071 B.n691 B.n331 10.6151
R1072 B.n692 B.n691 10.6151
R1073 B.n693 B.n692 10.6151
R1074 B.n693 B.n323 10.6151
R1075 B.n704 B.n323 10.6151
R1076 B.n705 B.n704 10.6151
R1077 B.n706 B.n705 10.6151
R1078 B.n706 B.n0 10.6151
R1079 B.n426 B.n362 10.6151
R1080 B.n427 B.n426 10.6151
R1081 B.n428 B.n427 10.6151
R1082 B.n428 B.n422 10.6151
R1083 B.n434 B.n422 10.6151
R1084 B.n435 B.n434 10.6151
R1085 B.n436 B.n435 10.6151
R1086 B.n436 B.n420 10.6151
R1087 B.n442 B.n420 10.6151
R1088 B.n443 B.n442 10.6151
R1089 B.n444 B.n443 10.6151
R1090 B.n444 B.n418 10.6151
R1091 B.n450 B.n418 10.6151
R1092 B.n451 B.n450 10.6151
R1093 B.n452 B.n451 10.6151
R1094 B.n452 B.n416 10.6151
R1095 B.n458 B.n416 10.6151
R1096 B.n459 B.n458 10.6151
R1097 B.n460 B.n459 10.6151
R1098 B.n460 B.n414 10.6151
R1099 B.n466 B.n414 10.6151
R1100 B.n467 B.n466 10.6151
R1101 B.n468 B.n467 10.6151
R1102 B.n468 B.n412 10.6151
R1103 B.n474 B.n412 10.6151
R1104 B.n475 B.n474 10.6151
R1105 B.n476 B.n475 10.6151
R1106 B.n476 B.n410 10.6151
R1107 B.n482 B.n410 10.6151
R1108 B.n483 B.n482 10.6151
R1109 B.n484 B.n483 10.6151
R1110 B.n484 B.n408 10.6151
R1111 B.n490 B.n408 10.6151
R1112 B.n491 B.n490 10.6151
R1113 B.n492 B.n491 10.6151
R1114 B.n492 B.n406 10.6151
R1115 B.n498 B.n406 10.6151
R1116 B.n499 B.n498 10.6151
R1117 B.n500 B.n499 10.6151
R1118 B.n500 B.n404 10.6151
R1119 B.n506 B.n404 10.6151
R1120 B.n507 B.n506 10.6151
R1121 B.n508 B.n507 10.6151
R1122 B.n508 B.n402 10.6151
R1123 B.n514 B.n402 10.6151
R1124 B.n515 B.n514 10.6151
R1125 B.n516 B.n515 10.6151
R1126 B.n516 B.n400 10.6151
R1127 B.n523 B.n522 10.6151
R1128 B.n524 B.n523 10.6151
R1129 B.n524 B.n395 10.6151
R1130 B.n530 B.n395 10.6151
R1131 B.n531 B.n530 10.6151
R1132 B.n532 B.n531 10.6151
R1133 B.n532 B.n393 10.6151
R1134 B.n538 B.n393 10.6151
R1135 B.n539 B.n538 10.6151
R1136 B.n541 B.n389 10.6151
R1137 B.n547 B.n389 10.6151
R1138 B.n548 B.n547 10.6151
R1139 B.n549 B.n548 10.6151
R1140 B.n549 B.n387 10.6151
R1141 B.n555 B.n387 10.6151
R1142 B.n556 B.n555 10.6151
R1143 B.n557 B.n556 10.6151
R1144 B.n557 B.n385 10.6151
R1145 B.n563 B.n385 10.6151
R1146 B.n564 B.n563 10.6151
R1147 B.n565 B.n564 10.6151
R1148 B.n565 B.n383 10.6151
R1149 B.n571 B.n383 10.6151
R1150 B.n572 B.n571 10.6151
R1151 B.n573 B.n572 10.6151
R1152 B.n573 B.n381 10.6151
R1153 B.n579 B.n381 10.6151
R1154 B.n580 B.n579 10.6151
R1155 B.n581 B.n580 10.6151
R1156 B.n581 B.n379 10.6151
R1157 B.n587 B.n379 10.6151
R1158 B.n588 B.n587 10.6151
R1159 B.n589 B.n588 10.6151
R1160 B.n589 B.n377 10.6151
R1161 B.n595 B.n377 10.6151
R1162 B.n596 B.n595 10.6151
R1163 B.n597 B.n596 10.6151
R1164 B.n597 B.n375 10.6151
R1165 B.n603 B.n375 10.6151
R1166 B.n604 B.n603 10.6151
R1167 B.n605 B.n604 10.6151
R1168 B.n605 B.n373 10.6151
R1169 B.n611 B.n373 10.6151
R1170 B.n612 B.n611 10.6151
R1171 B.n613 B.n612 10.6151
R1172 B.n613 B.n371 10.6151
R1173 B.n619 B.n371 10.6151
R1174 B.n620 B.n619 10.6151
R1175 B.n621 B.n620 10.6151
R1176 B.n621 B.n369 10.6151
R1177 B.n627 B.n369 10.6151
R1178 B.n628 B.n627 10.6151
R1179 B.n629 B.n628 10.6151
R1180 B.n629 B.n367 10.6151
R1181 B.n367 B.n366 10.6151
R1182 B.n636 B.n366 10.6151
R1183 B.n637 B.n636 10.6151
R1184 B.n638 B.n358 10.6151
R1185 B.n648 B.n358 10.6151
R1186 B.n649 B.n648 10.6151
R1187 B.n650 B.n649 10.6151
R1188 B.n650 B.n351 10.6151
R1189 B.n661 B.n351 10.6151
R1190 B.n662 B.n661 10.6151
R1191 B.n663 B.n662 10.6151
R1192 B.n663 B.n343 10.6151
R1193 B.n673 B.n343 10.6151
R1194 B.n674 B.n673 10.6151
R1195 B.n675 B.n674 10.6151
R1196 B.n675 B.n335 10.6151
R1197 B.n685 B.n335 10.6151
R1198 B.n686 B.n685 10.6151
R1199 B.n687 B.n686 10.6151
R1200 B.n687 B.n327 10.6151
R1201 B.n697 B.n327 10.6151
R1202 B.n698 B.n697 10.6151
R1203 B.n700 B.n698 10.6151
R1204 B.n700 B.n699 10.6151
R1205 B.n699 B.n319 10.6151
R1206 B.n711 B.n319 10.6151
R1207 B.n712 B.n711 10.6151
R1208 B.n713 B.n712 10.6151
R1209 B.n714 B.n713 10.6151
R1210 B.n715 B.n714 10.6151
R1211 B.n719 B.n715 10.6151
R1212 B.n720 B.n719 10.6151
R1213 B.n721 B.n720 10.6151
R1214 B.n722 B.n721 10.6151
R1215 B.n724 B.n722 10.6151
R1216 B.n725 B.n724 10.6151
R1217 B.n726 B.n725 10.6151
R1218 B.n727 B.n726 10.6151
R1219 B.n729 B.n727 10.6151
R1220 B.n730 B.n729 10.6151
R1221 B.n731 B.n730 10.6151
R1222 B.n732 B.n731 10.6151
R1223 B.n734 B.n732 10.6151
R1224 B.n735 B.n734 10.6151
R1225 B.n736 B.n735 10.6151
R1226 B.n737 B.n736 10.6151
R1227 B.n739 B.n737 10.6151
R1228 B.n740 B.n739 10.6151
R1229 B.n741 B.n740 10.6151
R1230 B.n742 B.n741 10.6151
R1231 B.n744 B.n742 10.6151
R1232 B.n745 B.n744 10.6151
R1233 B.n794 B.n1 10.6151
R1234 B.n794 B.n793 10.6151
R1235 B.n793 B.n792 10.6151
R1236 B.n792 B.n10 10.6151
R1237 B.n786 B.n10 10.6151
R1238 B.n786 B.n785 10.6151
R1239 B.n785 B.n784 10.6151
R1240 B.n784 B.n17 10.6151
R1241 B.n778 B.n17 10.6151
R1242 B.n778 B.n777 10.6151
R1243 B.n777 B.n776 10.6151
R1244 B.n776 B.n24 10.6151
R1245 B.n770 B.n24 10.6151
R1246 B.n770 B.n769 10.6151
R1247 B.n769 B.n768 10.6151
R1248 B.n768 B.n31 10.6151
R1249 B.n762 B.n31 10.6151
R1250 B.n762 B.n761 10.6151
R1251 B.n761 B.n760 10.6151
R1252 B.n760 B.n37 10.6151
R1253 B.n754 B.n37 10.6151
R1254 B.n754 B.n753 10.6151
R1255 B.n753 B.n752 10.6151
R1256 B.n106 B.n45 10.6151
R1257 B.n109 B.n106 10.6151
R1258 B.n110 B.n109 10.6151
R1259 B.n113 B.n110 10.6151
R1260 B.n114 B.n113 10.6151
R1261 B.n117 B.n114 10.6151
R1262 B.n118 B.n117 10.6151
R1263 B.n121 B.n118 10.6151
R1264 B.n122 B.n121 10.6151
R1265 B.n125 B.n122 10.6151
R1266 B.n126 B.n125 10.6151
R1267 B.n129 B.n126 10.6151
R1268 B.n130 B.n129 10.6151
R1269 B.n133 B.n130 10.6151
R1270 B.n134 B.n133 10.6151
R1271 B.n137 B.n134 10.6151
R1272 B.n138 B.n137 10.6151
R1273 B.n141 B.n138 10.6151
R1274 B.n142 B.n141 10.6151
R1275 B.n145 B.n142 10.6151
R1276 B.n146 B.n145 10.6151
R1277 B.n149 B.n146 10.6151
R1278 B.n150 B.n149 10.6151
R1279 B.n153 B.n150 10.6151
R1280 B.n154 B.n153 10.6151
R1281 B.n157 B.n154 10.6151
R1282 B.n158 B.n157 10.6151
R1283 B.n161 B.n158 10.6151
R1284 B.n162 B.n161 10.6151
R1285 B.n165 B.n162 10.6151
R1286 B.n166 B.n165 10.6151
R1287 B.n169 B.n166 10.6151
R1288 B.n170 B.n169 10.6151
R1289 B.n173 B.n170 10.6151
R1290 B.n174 B.n173 10.6151
R1291 B.n177 B.n174 10.6151
R1292 B.n178 B.n177 10.6151
R1293 B.n181 B.n178 10.6151
R1294 B.n182 B.n181 10.6151
R1295 B.n185 B.n182 10.6151
R1296 B.n186 B.n185 10.6151
R1297 B.n189 B.n186 10.6151
R1298 B.n190 B.n189 10.6151
R1299 B.n193 B.n190 10.6151
R1300 B.n194 B.n193 10.6151
R1301 B.n197 B.n194 10.6151
R1302 B.n198 B.n197 10.6151
R1303 B.n201 B.n198 10.6151
R1304 B.n206 B.n203 10.6151
R1305 B.n207 B.n206 10.6151
R1306 B.n210 B.n207 10.6151
R1307 B.n211 B.n210 10.6151
R1308 B.n214 B.n211 10.6151
R1309 B.n215 B.n214 10.6151
R1310 B.n218 B.n215 10.6151
R1311 B.n219 B.n218 10.6151
R1312 B.n222 B.n219 10.6151
R1313 B.n227 B.n224 10.6151
R1314 B.n228 B.n227 10.6151
R1315 B.n231 B.n228 10.6151
R1316 B.n232 B.n231 10.6151
R1317 B.n235 B.n232 10.6151
R1318 B.n236 B.n235 10.6151
R1319 B.n239 B.n236 10.6151
R1320 B.n240 B.n239 10.6151
R1321 B.n243 B.n240 10.6151
R1322 B.n244 B.n243 10.6151
R1323 B.n247 B.n244 10.6151
R1324 B.n248 B.n247 10.6151
R1325 B.n251 B.n248 10.6151
R1326 B.n252 B.n251 10.6151
R1327 B.n255 B.n252 10.6151
R1328 B.n256 B.n255 10.6151
R1329 B.n259 B.n256 10.6151
R1330 B.n260 B.n259 10.6151
R1331 B.n263 B.n260 10.6151
R1332 B.n264 B.n263 10.6151
R1333 B.n267 B.n264 10.6151
R1334 B.n268 B.n267 10.6151
R1335 B.n271 B.n268 10.6151
R1336 B.n272 B.n271 10.6151
R1337 B.n275 B.n272 10.6151
R1338 B.n276 B.n275 10.6151
R1339 B.n279 B.n276 10.6151
R1340 B.n280 B.n279 10.6151
R1341 B.n283 B.n280 10.6151
R1342 B.n284 B.n283 10.6151
R1343 B.n287 B.n284 10.6151
R1344 B.n288 B.n287 10.6151
R1345 B.n291 B.n288 10.6151
R1346 B.n292 B.n291 10.6151
R1347 B.n295 B.n292 10.6151
R1348 B.n296 B.n295 10.6151
R1349 B.n299 B.n296 10.6151
R1350 B.n300 B.n299 10.6151
R1351 B.n303 B.n300 10.6151
R1352 B.n304 B.n303 10.6151
R1353 B.n307 B.n304 10.6151
R1354 B.n308 B.n307 10.6151
R1355 B.n311 B.n308 10.6151
R1356 B.n312 B.n311 10.6151
R1357 B.n315 B.n312 10.6151
R1358 B.n317 B.n315 10.6151
R1359 B.n318 B.n317 10.6151
R1360 B.n746 B.n318 10.6151
R1361 B.n400 B.n399 9.36635
R1362 B.n541 B.n540 9.36635
R1363 B.n202 B.n201 9.36635
R1364 B.n224 B.n223 9.36635
R1365 B.n802 B.n0 8.11757
R1366 B.n802 B.n1 8.11757
R1367 B.n702 B.t1 5.55465
R1368 B.n790 B.t3 5.55465
R1369 B.n659 B.t5 2.22216
R1370 B.n764 B.t12 2.22216
R1371 B.n522 B.n399 1.24928
R1372 B.n540 B.n539 1.24928
R1373 B.n203 B.n202 1.24928
R1374 B.n223 B.n222 1.24928
R1375 VP.n2 VP.t0 264.325
R1376 VP.n2 VP.t1 264.005
R1377 VP.n4 VP.t3 227.386
R1378 VP.n11 VP.t2 227.386
R1379 VP.n4 VP.n3 176.714
R1380 VP.n12 VP.n11 176.714
R1381 VP.n10 VP.n0 161.3
R1382 VP.n9 VP.n8 161.3
R1383 VP.n7 VP.n1 161.3
R1384 VP.n6 VP.n5 161.3
R1385 VP.n3 VP.n2 57.8115
R1386 VP.n9 VP.n1 56.5193
R1387 VP.n5 VP.n1 24.4675
R1388 VP.n10 VP.n9 24.4675
R1389 VP.n5 VP.n4 9.05329
R1390 VP.n11 VP.n10 9.05329
R1391 VP.n6 VP.n3 0.189894
R1392 VP.n7 VP.n6 0.189894
R1393 VP.n8 VP.n7 0.189894
R1394 VP.n8 VP.n0 0.189894
R1395 VP.n12 VP.n0 0.189894
R1396 VP VP.n12 0.0516364
R1397 VDD1 VDD1.n1 100.841
R1398 VDD1 VDD1.n0 59.2973
R1399 VDD1.n0 VDD1.t3 1.3632
R1400 VDD1.n0 VDD1.t2 1.3632
R1401 VDD1.n1 VDD1.t0 1.3632
R1402 VDD1.n1 VDD1.t1 1.3632
C0 VDD2 VDD1 0.769559f
C1 VP VDD1 5.21798f
C2 VDD2 VP 0.326974f
C3 VTAIL VN 4.69152f
C4 VN VDD1 0.148161f
C5 VTAIL VDD1 6.26451f
C6 VDD2 VN 5.03964f
C7 VDD2 VTAIL 6.31161f
C8 VN VP 5.89533f
C9 VTAIL VP 4.70563f
C10 VDD2 B 3.370049f
C11 VDD1 B 7.43082f
C12 VTAIL B 10.912781f
C13 VN B 9.15134f
C14 VP B 6.840808f
C15 VDD1.t3 B 0.307386f
C16 VDD1.t2 B 0.307386f
C17 VDD1.n0 B 2.76519f
C18 VDD1.t0 B 0.307386f
C19 VDD1.t1 B 0.307386f
C20 VDD1.n1 B 3.51931f
C21 VP.n0 B 0.034653f
C22 VP.t2 B 2.12321f
C23 VP.n1 B 0.050588f
C24 VP.t0 B 2.24887f
C25 VP.t1 B 2.24776f
C26 VP.n2 B 2.99113f
C27 VP.n3 B 2.03016f
C28 VP.t3 B 2.12321f
C29 VP.n4 B 0.828286f
C30 VP.n5 B 0.044495f
C31 VP.n6 B 0.034653f
C32 VP.n7 B 0.034653f
C33 VP.n8 B 0.034653f
C34 VP.n9 B 0.050588f
C35 VP.n10 B 0.044495f
C36 VP.n11 B 0.828286f
C37 VP.n12 B 0.03374f
C38 VDD2.t2 B 0.30466f
C39 VDD2.t3 B 0.30466f
C40 VDD2.n0 B 3.4608f
C41 VDD2.t0 B 0.30466f
C42 VDD2.t1 B 0.30466f
C43 VDD2.n1 B 2.74029f
C44 VDD2.n2 B 3.73673f
C45 VTAIL.t4 B 1.97954f
C46 VTAIL.n0 B 0.286119f
C47 VTAIL.t1 B 1.97954f
C48 VTAIL.n1 B 0.3235f
C49 VTAIL.t2 B 1.97954f
C50 VTAIL.n2 B 1.21743f
C51 VTAIL.t7 B 1.97954f
C52 VTAIL.n3 B 1.21742f
C53 VTAIL.t6 B 1.97954f
C54 VTAIL.n4 B 0.323495f
C55 VTAIL.t3 B 1.97954f
C56 VTAIL.n5 B 0.323495f
C57 VTAIL.t0 B 1.97955f
C58 VTAIL.n6 B 1.21742f
C59 VTAIL.t5 B 1.97954f
C60 VTAIL.n7 B 1.17423f
C61 VN.t1 B 2.21358f
C62 VN.t0 B 2.21249f
C63 VN.n0 B 1.576f
C64 VN.t2 B 2.21358f
C65 VN.t3 B 2.21249f
C66 VN.n1 B 2.96412f
.ends

