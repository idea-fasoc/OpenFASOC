* NGSPICE file created from diff_pair_sample_0005.ext - technology: sky130A

.subckt diff_pair_sample_0005 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t4 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.30525 ps=2.18 w=1.85 l=3.47
X1 VDD1.t5 VP.t0 VTAIL.t0 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0.30525 ps=2.18 w=1.85 l=3.47
X2 VDD2.t5 VN.t1 VTAIL.t10 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0.30525 ps=2.18 w=1.85 l=3.47
X3 VDD1.t4 VP.t1 VTAIL.t3 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0.30525 ps=2.18 w=1.85 l=3.47
X4 B.t11 B.t9 B.t10 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0 ps=0 w=1.85 l=3.47
X5 VDD2.t3 VN.t2 VTAIL.t9 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.7215 ps=4.48 w=1.85 l=3.47
X6 B.t8 B.t6 B.t7 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0 ps=0 w=1.85 l=3.47
X7 VTAIL.t2 VP.t2 VDD1.t3 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.30525 ps=2.18 w=1.85 l=3.47
X8 VDD2.t2 VN.t3 VTAIL.t8 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0.30525 ps=2.18 w=1.85 l=3.47
X9 B.t5 B.t3 B.t4 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0 ps=0 w=1.85 l=3.47
X10 VDD2.t1 VN.t4 VTAIL.t7 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.7215 ps=4.48 w=1.85 l=3.47
X11 VDD1.t2 VP.t3 VTAIL.t5 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.7215 ps=4.48 w=1.85 l=3.47
X12 B.t2 B.t0 B.t1 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.7215 pd=4.48 as=0 ps=0 w=1.85 l=3.47
X13 VDD1.t1 VP.t4 VTAIL.t1 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.7215 ps=4.48 w=1.85 l=3.47
X14 VTAIL.t4 VP.t5 VDD1.t0 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.30525 ps=2.18 w=1.85 l=3.47
X15 VTAIL.t6 VN.t5 VDD2.t0 w_n4010_n1338# sky130_fd_pr__pfet_01v8 ad=0.30525 pd=2.18 as=0.30525 ps=2.18 w=1.85 l=3.47
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n17 VN.n0 75.3872
R15 VN.n35 VN.n18 75.3872
R16 VN.n9 VN.n2 50.2061
R17 VN.n27 VN.n20 50.2061
R18 VN.n5 VN.n4 50.1968
R19 VN.n23 VN.n22 50.1968
R20 VN.n5 VN.t1 46.9277
R21 VN.n23 VN.t2 46.9277
R22 VN VN.n35 44.7177
R23 VN.n13 VN.n2 30.7807
R24 VN.n31 VN.n20 30.7807
R25 VN.n7 VN.n4 24.4675
R26 VN.n8 VN.n7 24.4675
R27 VN.n9 VN.n8 24.4675
R28 VN.n14 VN.n13 24.4675
R29 VN.n15 VN.n14 24.4675
R30 VN.n27 VN.n26 24.4675
R31 VN.n26 VN.n25 24.4675
R32 VN.n25 VN.n22 24.4675
R33 VN.n33 VN.n32 24.4675
R34 VN.n32 VN.n31 24.4675
R35 VN.n15 VN.n0 14.6807
R36 VN.n33 VN.n18 14.6807
R37 VN.n4 VN.t5 12.8492
R38 VN.n0 VN.t4 12.8492
R39 VN.n22 VN.t0 12.8492
R40 VN.n18 VN.t3 12.8492
R41 VN.n6 VN.n5 2.99386
R42 VN.n24 VN.n23 2.99386
R43 VN.n35 VN.n34 0.354971
R44 VN.n17 VN.n16 0.354971
R45 VN VN.n17 0.26696
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VDD2.n11 VDD2.n9 756.745
R59 VDD2.n2 VDD2.n0 756.745
R60 VDD2.n12 VDD2.n11 585
R61 VDD2.n3 VDD2.n2 585
R62 VDD2.t5 VDD2.n1 415.613
R63 VDD2.t2 VDD2.n10 415.613
R64 VDD2.n8 VDD2.n7 203.619
R65 VDD2 VDD2.n17 203.617
R66 VDD2.n11 VDD2.t2 85.8723
R67 VDD2.n2 VDD2.t5 85.8723
R68 VDD2.n8 VDD2.n6 54.5627
R69 VDD2.n16 VDD2.n15 52.1611
R70 VDD2.n16 VDD2.n8 35.9567
R71 VDD2.n17 VDD2.t4 17.5708
R72 VDD2.n17 VDD2.t3 17.5708
R73 VDD2.n7 VDD2.t0 17.5708
R74 VDD2.n7 VDD2.t1 17.5708
R75 VDD2.n12 VDD2.n10 14.9339
R76 VDD2.n3 VDD2.n1 14.9339
R77 VDD2.n13 VDD2.n9 12.8005
R78 VDD2.n4 VDD2.n0 12.8005
R79 VDD2.n15 VDD2.n14 9.45567
R80 VDD2.n6 VDD2.n5 9.45567
R81 VDD2.n14 VDD2.n13 9.3005
R82 VDD2.n5 VDD2.n4 9.3005
R83 VDD2.n14 VDD2.n10 5.44463
R84 VDD2.n5 VDD2.n1 5.44463
R85 VDD2 VDD2.n16 2.51559
R86 VDD2.n15 VDD2.n9 1.16414
R87 VDD2.n6 VDD2.n0 1.16414
R88 VDD2.n13 VDD2.n12 0.388379
R89 VDD2.n4 VDD2.n3 0.388379
R90 VTAIL.n34 VTAIL.n32 756.745
R91 VTAIL.n4 VTAIL.n2 756.745
R92 VTAIL.n26 VTAIL.n24 756.745
R93 VTAIL.n16 VTAIL.n14 756.745
R94 VTAIL.n35 VTAIL.n34 585
R95 VTAIL.n5 VTAIL.n4 585
R96 VTAIL.n27 VTAIL.n26 585
R97 VTAIL.n17 VTAIL.n16 585
R98 VTAIL.t7 VTAIL.n33 415.613
R99 VTAIL.t5 VTAIL.n3 415.613
R100 VTAIL.t1 VTAIL.n25 415.613
R101 VTAIL.t9 VTAIL.n15 415.613
R102 VTAIL.n23 VTAIL.n22 186.177
R103 VTAIL.n13 VTAIL.n12 186.177
R104 VTAIL.n1 VTAIL.n0 186.177
R105 VTAIL.n11 VTAIL.n10 186.177
R106 VTAIL.n34 VTAIL.t7 85.8723
R107 VTAIL.n4 VTAIL.t5 85.8723
R108 VTAIL.n26 VTAIL.t1 85.8723
R109 VTAIL.n16 VTAIL.t9 85.8723
R110 VTAIL.n39 VTAIL.n38 35.4823
R111 VTAIL.n9 VTAIL.n8 35.4823
R112 VTAIL.n31 VTAIL.n30 35.4823
R113 VTAIL.n21 VTAIL.n20 35.4823
R114 VTAIL.n13 VTAIL.n11 20.5134
R115 VTAIL.n0 VTAIL.t10 17.5708
R116 VTAIL.n0 VTAIL.t6 17.5708
R117 VTAIL.n10 VTAIL.t3 17.5708
R118 VTAIL.n10 VTAIL.t4 17.5708
R119 VTAIL.n22 VTAIL.t0 17.5708
R120 VTAIL.n22 VTAIL.t2 17.5708
R121 VTAIL.n12 VTAIL.t8 17.5708
R122 VTAIL.n12 VTAIL.t11 17.5708
R123 VTAIL.n39 VTAIL.n31 17.2376
R124 VTAIL.n35 VTAIL.n33 14.9339
R125 VTAIL.n5 VTAIL.n3 14.9339
R126 VTAIL.n27 VTAIL.n25 14.9339
R127 VTAIL.n17 VTAIL.n15 14.9339
R128 VTAIL.n36 VTAIL.n32 12.8005
R129 VTAIL.n6 VTAIL.n2 12.8005
R130 VTAIL.n28 VTAIL.n24 12.8005
R131 VTAIL.n18 VTAIL.n14 12.8005
R132 VTAIL.n38 VTAIL.n37 9.45567
R133 VTAIL.n8 VTAIL.n7 9.45567
R134 VTAIL.n30 VTAIL.n29 9.45567
R135 VTAIL.n20 VTAIL.n19 9.45567
R136 VTAIL.n37 VTAIL.n36 9.3005
R137 VTAIL.n7 VTAIL.n6 9.3005
R138 VTAIL.n29 VTAIL.n28 9.3005
R139 VTAIL.n19 VTAIL.n18 9.3005
R140 VTAIL.n37 VTAIL.n33 5.44463
R141 VTAIL.n7 VTAIL.n3 5.44463
R142 VTAIL.n29 VTAIL.n25 5.44463
R143 VTAIL.n19 VTAIL.n15 5.44463
R144 VTAIL.n21 VTAIL.n13 3.27636
R145 VTAIL.n31 VTAIL.n23 3.27636
R146 VTAIL.n11 VTAIL.n9 3.27636
R147 VTAIL VTAIL.n39 2.39921
R148 VTAIL.n23 VTAIL.n21 2.10826
R149 VTAIL.n9 VTAIL.n1 2.10826
R150 VTAIL.n38 VTAIL.n32 1.16414
R151 VTAIL.n8 VTAIL.n2 1.16414
R152 VTAIL.n30 VTAIL.n24 1.16414
R153 VTAIL.n20 VTAIL.n14 1.16414
R154 VTAIL VTAIL.n1 0.877655
R155 VTAIL.n36 VTAIL.n35 0.388379
R156 VTAIL.n6 VTAIL.n5 0.388379
R157 VTAIL.n28 VTAIL.n27 0.388379
R158 VTAIL.n18 VTAIL.n17 0.388379
R159 VP.n16 VP.n15 161.3
R160 VP.n17 VP.n12 161.3
R161 VP.n19 VP.n18 161.3
R162 VP.n20 VP.n11 161.3
R163 VP.n22 VP.n21 161.3
R164 VP.n23 VP.n10 161.3
R165 VP.n25 VP.n24 161.3
R166 VP.n50 VP.n49 161.3
R167 VP.n48 VP.n1 161.3
R168 VP.n47 VP.n46 161.3
R169 VP.n45 VP.n2 161.3
R170 VP.n44 VP.n43 161.3
R171 VP.n42 VP.n3 161.3
R172 VP.n41 VP.n40 161.3
R173 VP.n39 VP.n4 161.3
R174 VP.n38 VP.n37 161.3
R175 VP.n36 VP.n5 161.3
R176 VP.n35 VP.n34 161.3
R177 VP.n33 VP.n6 161.3
R178 VP.n32 VP.n31 161.3
R179 VP.n30 VP.n7 161.3
R180 VP.n29 VP.n28 161.3
R181 VP.n27 VP.n8 75.3872
R182 VP.n51 VP.n0 75.3872
R183 VP.n26 VP.n9 75.3872
R184 VP.n35 VP.n6 50.2061
R185 VP.n43 VP.n2 50.2061
R186 VP.n18 VP.n11 50.2061
R187 VP.n14 VP.n13 50.1968
R188 VP.n14 VP.t0 46.9275
R189 VP.n27 VP.n26 44.5524
R190 VP.n31 VP.n6 30.7807
R191 VP.n47 VP.n2 30.7807
R192 VP.n22 VP.n11 30.7807
R193 VP.n30 VP.n29 24.4675
R194 VP.n31 VP.n30 24.4675
R195 VP.n36 VP.n35 24.4675
R196 VP.n37 VP.n36 24.4675
R197 VP.n37 VP.n4 24.4675
R198 VP.n41 VP.n4 24.4675
R199 VP.n42 VP.n41 24.4675
R200 VP.n43 VP.n42 24.4675
R201 VP.n48 VP.n47 24.4675
R202 VP.n49 VP.n48 24.4675
R203 VP.n23 VP.n22 24.4675
R204 VP.n24 VP.n23 24.4675
R205 VP.n16 VP.n13 24.4675
R206 VP.n17 VP.n16 24.4675
R207 VP.n18 VP.n17 24.4675
R208 VP.n29 VP.n8 14.6807
R209 VP.n49 VP.n0 14.6807
R210 VP.n24 VP.n9 14.6807
R211 VP.n4 VP.t5 12.8492
R212 VP.n8 VP.t1 12.8492
R213 VP.n0 VP.t3 12.8492
R214 VP.n13 VP.t2 12.8492
R215 VP.n9 VP.t4 12.8492
R216 VP.n15 VP.n14 2.99384
R217 VP.n26 VP.n25 0.354971
R218 VP.n28 VP.n27 0.354971
R219 VP.n51 VP.n50 0.354971
R220 VP VP.n51 0.26696
R221 VP.n15 VP.n12 0.189894
R222 VP.n19 VP.n12 0.189894
R223 VP.n20 VP.n19 0.189894
R224 VP.n21 VP.n20 0.189894
R225 VP.n21 VP.n10 0.189894
R226 VP.n25 VP.n10 0.189894
R227 VP.n28 VP.n7 0.189894
R228 VP.n32 VP.n7 0.189894
R229 VP.n33 VP.n32 0.189894
R230 VP.n34 VP.n33 0.189894
R231 VP.n34 VP.n5 0.189894
R232 VP.n38 VP.n5 0.189894
R233 VP.n39 VP.n38 0.189894
R234 VP.n40 VP.n39 0.189894
R235 VP.n40 VP.n3 0.189894
R236 VP.n44 VP.n3 0.189894
R237 VP.n45 VP.n44 0.189894
R238 VP.n46 VP.n45 0.189894
R239 VP.n46 VP.n1 0.189894
R240 VP.n50 VP.n1 0.189894
R241 VDD1.n2 VDD1.n0 756.745
R242 VDD1.n9 VDD1.n7 756.745
R243 VDD1.n3 VDD1.n2 585
R244 VDD1.n10 VDD1.n9 585
R245 VDD1.t4 VDD1.n8 415.613
R246 VDD1.t5 VDD1.n1 415.613
R247 VDD1.n15 VDD1.n14 203.619
R248 VDD1.n17 VDD1.n16 202.856
R249 VDD1.n2 VDD1.t5 85.8723
R250 VDD1.n9 VDD1.t4 85.8723
R251 VDD1 VDD1.n6 54.6762
R252 VDD1.n15 VDD1.n13 54.5627
R253 VDD1.n17 VDD1.n15 38.1776
R254 VDD1.n16 VDD1.t3 17.5708
R255 VDD1.n16 VDD1.t1 17.5708
R256 VDD1.n14 VDD1.t0 17.5708
R257 VDD1.n14 VDD1.t2 17.5708
R258 VDD1.n3 VDD1.n1 14.9339
R259 VDD1.n10 VDD1.n8 14.9339
R260 VDD1.n4 VDD1.n0 12.8005
R261 VDD1.n11 VDD1.n7 12.8005
R262 VDD1.n6 VDD1.n5 9.45567
R263 VDD1.n13 VDD1.n12 9.45567
R264 VDD1.n5 VDD1.n4 9.3005
R265 VDD1.n12 VDD1.n11 9.3005
R266 VDD1.n5 VDD1.n1 5.44463
R267 VDD1.n12 VDD1.n8 5.44463
R268 VDD1.n6 VDD1.n0 1.16414
R269 VDD1.n13 VDD1.n7 1.16414
R270 VDD1 VDD1.n17 0.761276
R271 VDD1.n4 VDD1.n3 0.388379
R272 VDD1.n11 VDD1.n10 0.388379
R273 B.n441 B.n440 585
R274 B.n442 B.n49 585
R275 B.n444 B.n443 585
R276 B.n445 B.n48 585
R277 B.n447 B.n446 585
R278 B.n448 B.n47 585
R279 B.n450 B.n449 585
R280 B.n451 B.n46 585
R281 B.n453 B.n452 585
R282 B.n454 B.n45 585
R283 B.n456 B.n455 585
R284 B.n457 B.n42 585
R285 B.n460 B.n459 585
R286 B.n461 B.n41 585
R287 B.n463 B.n462 585
R288 B.n464 B.n40 585
R289 B.n466 B.n465 585
R290 B.n467 B.n39 585
R291 B.n469 B.n468 585
R292 B.n470 B.n35 585
R293 B.n472 B.n471 585
R294 B.n473 B.n34 585
R295 B.n475 B.n474 585
R296 B.n476 B.n33 585
R297 B.n478 B.n477 585
R298 B.n479 B.n32 585
R299 B.n481 B.n480 585
R300 B.n482 B.n31 585
R301 B.n484 B.n483 585
R302 B.n485 B.n30 585
R303 B.n487 B.n486 585
R304 B.n488 B.n29 585
R305 B.n490 B.n489 585
R306 B.n439 B.n50 585
R307 B.n438 B.n437 585
R308 B.n436 B.n51 585
R309 B.n435 B.n434 585
R310 B.n433 B.n52 585
R311 B.n432 B.n431 585
R312 B.n430 B.n53 585
R313 B.n429 B.n428 585
R314 B.n427 B.n54 585
R315 B.n426 B.n425 585
R316 B.n424 B.n55 585
R317 B.n423 B.n422 585
R318 B.n421 B.n56 585
R319 B.n420 B.n419 585
R320 B.n418 B.n57 585
R321 B.n417 B.n416 585
R322 B.n415 B.n58 585
R323 B.n414 B.n413 585
R324 B.n412 B.n59 585
R325 B.n411 B.n410 585
R326 B.n409 B.n60 585
R327 B.n408 B.n407 585
R328 B.n406 B.n61 585
R329 B.n405 B.n404 585
R330 B.n403 B.n62 585
R331 B.n402 B.n401 585
R332 B.n400 B.n63 585
R333 B.n399 B.n398 585
R334 B.n397 B.n64 585
R335 B.n396 B.n395 585
R336 B.n394 B.n65 585
R337 B.n393 B.n392 585
R338 B.n391 B.n66 585
R339 B.n390 B.n389 585
R340 B.n388 B.n67 585
R341 B.n387 B.n386 585
R342 B.n385 B.n68 585
R343 B.n384 B.n383 585
R344 B.n382 B.n69 585
R345 B.n381 B.n380 585
R346 B.n379 B.n70 585
R347 B.n378 B.n377 585
R348 B.n376 B.n71 585
R349 B.n375 B.n374 585
R350 B.n373 B.n72 585
R351 B.n372 B.n371 585
R352 B.n370 B.n73 585
R353 B.n369 B.n368 585
R354 B.n367 B.n74 585
R355 B.n366 B.n365 585
R356 B.n364 B.n75 585
R357 B.n363 B.n362 585
R358 B.n361 B.n76 585
R359 B.n360 B.n359 585
R360 B.n358 B.n77 585
R361 B.n357 B.n356 585
R362 B.n355 B.n78 585
R363 B.n354 B.n353 585
R364 B.n352 B.n79 585
R365 B.n351 B.n350 585
R366 B.n349 B.n80 585
R367 B.n348 B.n347 585
R368 B.n346 B.n81 585
R369 B.n345 B.n344 585
R370 B.n343 B.n82 585
R371 B.n342 B.n341 585
R372 B.n340 B.n83 585
R373 B.n339 B.n338 585
R374 B.n337 B.n84 585
R375 B.n336 B.n335 585
R376 B.n334 B.n85 585
R377 B.n333 B.n332 585
R378 B.n331 B.n86 585
R379 B.n330 B.n329 585
R380 B.n328 B.n87 585
R381 B.n327 B.n326 585
R382 B.n325 B.n88 585
R383 B.n324 B.n323 585
R384 B.n322 B.n89 585
R385 B.n321 B.n320 585
R386 B.n319 B.n90 585
R387 B.n318 B.n317 585
R388 B.n316 B.n91 585
R389 B.n315 B.n314 585
R390 B.n313 B.n92 585
R391 B.n312 B.n311 585
R392 B.n310 B.n93 585
R393 B.n309 B.n308 585
R394 B.n307 B.n94 585
R395 B.n306 B.n305 585
R396 B.n304 B.n95 585
R397 B.n303 B.n302 585
R398 B.n301 B.n96 585
R399 B.n300 B.n299 585
R400 B.n298 B.n97 585
R401 B.n297 B.n296 585
R402 B.n295 B.n98 585
R403 B.n294 B.n293 585
R404 B.n292 B.n99 585
R405 B.n291 B.n290 585
R406 B.n289 B.n100 585
R407 B.n288 B.n287 585
R408 B.n286 B.n101 585
R409 B.n285 B.n284 585
R410 B.n283 B.n102 585
R411 B.n282 B.n281 585
R412 B.n280 B.n103 585
R413 B.n227 B.n226 585
R414 B.n228 B.n121 585
R415 B.n230 B.n229 585
R416 B.n231 B.n120 585
R417 B.n233 B.n232 585
R418 B.n234 B.n119 585
R419 B.n236 B.n235 585
R420 B.n237 B.n118 585
R421 B.n239 B.n238 585
R422 B.n240 B.n117 585
R423 B.n242 B.n241 585
R424 B.n243 B.n114 585
R425 B.n246 B.n245 585
R426 B.n247 B.n113 585
R427 B.n249 B.n248 585
R428 B.n250 B.n112 585
R429 B.n252 B.n251 585
R430 B.n253 B.n111 585
R431 B.n255 B.n254 585
R432 B.n256 B.n110 585
R433 B.n261 B.n260 585
R434 B.n262 B.n109 585
R435 B.n264 B.n263 585
R436 B.n265 B.n108 585
R437 B.n267 B.n266 585
R438 B.n268 B.n107 585
R439 B.n270 B.n269 585
R440 B.n271 B.n106 585
R441 B.n273 B.n272 585
R442 B.n274 B.n105 585
R443 B.n276 B.n275 585
R444 B.n277 B.n104 585
R445 B.n279 B.n278 585
R446 B.n225 B.n122 585
R447 B.n224 B.n223 585
R448 B.n222 B.n123 585
R449 B.n221 B.n220 585
R450 B.n219 B.n124 585
R451 B.n218 B.n217 585
R452 B.n216 B.n125 585
R453 B.n215 B.n214 585
R454 B.n213 B.n126 585
R455 B.n212 B.n211 585
R456 B.n210 B.n127 585
R457 B.n209 B.n208 585
R458 B.n207 B.n128 585
R459 B.n206 B.n205 585
R460 B.n204 B.n129 585
R461 B.n203 B.n202 585
R462 B.n201 B.n130 585
R463 B.n200 B.n199 585
R464 B.n198 B.n131 585
R465 B.n197 B.n196 585
R466 B.n195 B.n132 585
R467 B.n194 B.n193 585
R468 B.n192 B.n133 585
R469 B.n191 B.n190 585
R470 B.n189 B.n134 585
R471 B.n188 B.n187 585
R472 B.n186 B.n135 585
R473 B.n185 B.n184 585
R474 B.n183 B.n136 585
R475 B.n182 B.n181 585
R476 B.n180 B.n137 585
R477 B.n179 B.n178 585
R478 B.n177 B.n138 585
R479 B.n176 B.n175 585
R480 B.n174 B.n139 585
R481 B.n173 B.n172 585
R482 B.n171 B.n140 585
R483 B.n170 B.n169 585
R484 B.n168 B.n141 585
R485 B.n167 B.n166 585
R486 B.n165 B.n142 585
R487 B.n164 B.n163 585
R488 B.n162 B.n143 585
R489 B.n161 B.n160 585
R490 B.n159 B.n144 585
R491 B.n158 B.n157 585
R492 B.n156 B.n145 585
R493 B.n155 B.n154 585
R494 B.n153 B.n146 585
R495 B.n152 B.n151 585
R496 B.n150 B.n147 585
R497 B.n149 B.n148 585
R498 B.n2 B.n0 585
R499 B.n569 B.n1 585
R500 B.n568 B.n567 585
R501 B.n566 B.n3 585
R502 B.n565 B.n564 585
R503 B.n563 B.n4 585
R504 B.n562 B.n561 585
R505 B.n560 B.n5 585
R506 B.n559 B.n558 585
R507 B.n557 B.n6 585
R508 B.n556 B.n555 585
R509 B.n554 B.n7 585
R510 B.n553 B.n552 585
R511 B.n551 B.n8 585
R512 B.n550 B.n549 585
R513 B.n548 B.n9 585
R514 B.n547 B.n546 585
R515 B.n545 B.n10 585
R516 B.n544 B.n543 585
R517 B.n542 B.n11 585
R518 B.n541 B.n540 585
R519 B.n539 B.n12 585
R520 B.n538 B.n537 585
R521 B.n536 B.n13 585
R522 B.n535 B.n534 585
R523 B.n533 B.n14 585
R524 B.n532 B.n531 585
R525 B.n530 B.n15 585
R526 B.n529 B.n528 585
R527 B.n527 B.n16 585
R528 B.n526 B.n525 585
R529 B.n524 B.n17 585
R530 B.n523 B.n522 585
R531 B.n521 B.n18 585
R532 B.n520 B.n519 585
R533 B.n518 B.n19 585
R534 B.n517 B.n516 585
R535 B.n515 B.n20 585
R536 B.n514 B.n513 585
R537 B.n512 B.n21 585
R538 B.n511 B.n510 585
R539 B.n509 B.n22 585
R540 B.n508 B.n507 585
R541 B.n506 B.n23 585
R542 B.n505 B.n504 585
R543 B.n503 B.n24 585
R544 B.n502 B.n501 585
R545 B.n500 B.n25 585
R546 B.n499 B.n498 585
R547 B.n497 B.n26 585
R548 B.n496 B.n495 585
R549 B.n494 B.n27 585
R550 B.n493 B.n492 585
R551 B.n491 B.n28 585
R552 B.n571 B.n570 585
R553 B.n227 B.n122 478.086
R554 B.n491 B.n490 478.086
R555 B.n280 B.n279 478.086
R556 B.n441 B.n50 478.086
R557 B.n257 B.t11 319.125
R558 B.n43 B.t4 319.125
R559 B.n115 B.t8 319.125
R560 B.n36 B.t1 319.125
R561 B.n258 B.t10 245.429
R562 B.n44 B.t5 245.429
R563 B.n116 B.t7 245.429
R564 B.n37 B.t2 245.429
R565 B.n257 B.t9 209.481
R566 B.n115 B.t6 209.481
R567 B.n36 B.t0 209.481
R568 B.n43 B.t3 209.481
R569 B.n223 B.n122 163.367
R570 B.n223 B.n222 163.367
R571 B.n222 B.n221 163.367
R572 B.n221 B.n124 163.367
R573 B.n217 B.n124 163.367
R574 B.n217 B.n216 163.367
R575 B.n216 B.n215 163.367
R576 B.n215 B.n126 163.367
R577 B.n211 B.n126 163.367
R578 B.n211 B.n210 163.367
R579 B.n210 B.n209 163.367
R580 B.n209 B.n128 163.367
R581 B.n205 B.n128 163.367
R582 B.n205 B.n204 163.367
R583 B.n204 B.n203 163.367
R584 B.n203 B.n130 163.367
R585 B.n199 B.n130 163.367
R586 B.n199 B.n198 163.367
R587 B.n198 B.n197 163.367
R588 B.n197 B.n132 163.367
R589 B.n193 B.n132 163.367
R590 B.n193 B.n192 163.367
R591 B.n192 B.n191 163.367
R592 B.n191 B.n134 163.367
R593 B.n187 B.n134 163.367
R594 B.n187 B.n186 163.367
R595 B.n186 B.n185 163.367
R596 B.n185 B.n136 163.367
R597 B.n181 B.n136 163.367
R598 B.n181 B.n180 163.367
R599 B.n180 B.n179 163.367
R600 B.n179 B.n138 163.367
R601 B.n175 B.n138 163.367
R602 B.n175 B.n174 163.367
R603 B.n174 B.n173 163.367
R604 B.n173 B.n140 163.367
R605 B.n169 B.n140 163.367
R606 B.n169 B.n168 163.367
R607 B.n168 B.n167 163.367
R608 B.n167 B.n142 163.367
R609 B.n163 B.n142 163.367
R610 B.n163 B.n162 163.367
R611 B.n162 B.n161 163.367
R612 B.n161 B.n144 163.367
R613 B.n157 B.n144 163.367
R614 B.n157 B.n156 163.367
R615 B.n156 B.n155 163.367
R616 B.n155 B.n146 163.367
R617 B.n151 B.n146 163.367
R618 B.n151 B.n150 163.367
R619 B.n150 B.n149 163.367
R620 B.n149 B.n2 163.367
R621 B.n570 B.n2 163.367
R622 B.n570 B.n569 163.367
R623 B.n569 B.n568 163.367
R624 B.n568 B.n3 163.367
R625 B.n564 B.n3 163.367
R626 B.n564 B.n563 163.367
R627 B.n563 B.n562 163.367
R628 B.n562 B.n5 163.367
R629 B.n558 B.n5 163.367
R630 B.n558 B.n557 163.367
R631 B.n557 B.n556 163.367
R632 B.n556 B.n7 163.367
R633 B.n552 B.n7 163.367
R634 B.n552 B.n551 163.367
R635 B.n551 B.n550 163.367
R636 B.n550 B.n9 163.367
R637 B.n546 B.n9 163.367
R638 B.n546 B.n545 163.367
R639 B.n545 B.n544 163.367
R640 B.n544 B.n11 163.367
R641 B.n540 B.n11 163.367
R642 B.n540 B.n539 163.367
R643 B.n539 B.n538 163.367
R644 B.n538 B.n13 163.367
R645 B.n534 B.n13 163.367
R646 B.n534 B.n533 163.367
R647 B.n533 B.n532 163.367
R648 B.n532 B.n15 163.367
R649 B.n528 B.n15 163.367
R650 B.n528 B.n527 163.367
R651 B.n527 B.n526 163.367
R652 B.n526 B.n17 163.367
R653 B.n522 B.n17 163.367
R654 B.n522 B.n521 163.367
R655 B.n521 B.n520 163.367
R656 B.n520 B.n19 163.367
R657 B.n516 B.n19 163.367
R658 B.n516 B.n515 163.367
R659 B.n515 B.n514 163.367
R660 B.n514 B.n21 163.367
R661 B.n510 B.n21 163.367
R662 B.n510 B.n509 163.367
R663 B.n509 B.n508 163.367
R664 B.n508 B.n23 163.367
R665 B.n504 B.n23 163.367
R666 B.n504 B.n503 163.367
R667 B.n503 B.n502 163.367
R668 B.n502 B.n25 163.367
R669 B.n498 B.n25 163.367
R670 B.n498 B.n497 163.367
R671 B.n497 B.n496 163.367
R672 B.n496 B.n27 163.367
R673 B.n492 B.n27 163.367
R674 B.n492 B.n491 163.367
R675 B.n228 B.n227 163.367
R676 B.n229 B.n228 163.367
R677 B.n229 B.n120 163.367
R678 B.n233 B.n120 163.367
R679 B.n234 B.n233 163.367
R680 B.n235 B.n234 163.367
R681 B.n235 B.n118 163.367
R682 B.n239 B.n118 163.367
R683 B.n240 B.n239 163.367
R684 B.n241 B.n240 163.367
R685 B.n241 B.n114 163.367
R686 B.n246 B.n114 163.367
R687 B.n247 B.n246 163.367
R688 B.n248 B.n247 163.367
R689 B.n248 B.n112 163.367
R690 B.n252 B.n112 163.367
R691 B.n253 B.n252 163.367
R692 B.n254 B.n253 163.367
R693 B.n254 B.n110 163.367
R694 B.n261 B.n110 163.367
R695 B.n262 B.n261 163.367
R696 B.n263 B.n262 163.367
R697 B.n263 B.n108 163.367
R698 B.n267 B.n108 163.367
R699 B.n268 B.n267 163.367
R700 B.n269 B.n268 163.367
R701 B.n269 B.n106 163.367
R702 B.n273 B.n106 163.367
R703 B.n274 B.n273 163.367
R704 B.n275 B.n274 163.367
R705 B.n275 B.n104 163.367
R706 B.n279 B.n104 163.367
R707 B.n281 B.n280 163.367
R708 B.n281 B.n102 163.367
R709 B.n285 B.n102 163.367
R710 B.n286 B.n285 163.367
R711 B.n287 B.n286 163.367
R712 B.n287 B.n100 163.367
R713 B.n291 B.n100 163.367
R714 B.n292 B.n291 163.367
R715 B.n293 B.n292 163.367
R716 B.n293 B.n98 163.367
R717 B.n297 B.n98 163.367
R718 B.n298 B.n297 163.367
R719 B.n299 B.n298 163.367
R720 B.n299 B.n96 163.367
R721 B.n303 B.n96 163.367
R722 B.n304 B.n303 163.367
R723 B.n305 B.n304 163.367
R724 B.n305 B.n94 163.367
R725 B.n309 B.n94 163.367
R726 B.n310 B.n309 163.367
R727 B.n311 B.n310 163.367
R728 B.n311 B.n92 163.367
R729 B.n315 B.n92 163.367
R730 B.n316 B.n315 163.367
R731 B.n317 B.n316 163.367
R732 B.n317 B.n90 163.367
R733 B.n321 B.n90 163.367
R734 B.n322 B.n321 163.367
R735 B.n323 B.n322 163.367
R736 B.n323 B.n88 163.367
R737 B.n327 B.n88 163.367
R738 B.n328 B.n327 163.367
R739 B.n329 B.n328 163.367
R740 B.n329 B.n86 163.367
R741 B.n333 B.n86 163.367
R742 B.n334 B.n333 163.367
R743 B.n335 B.n334 163.367
R744 B.n335 B.n84 163.367
R745 B.n339 B.n84 163.367
R746 B.n340 B.n339 163.367
R747 B.n341 B.n340 163.367
R748 B.n341 B.n82 163.367
R749 B.n345 B.n82 163.367
R750 B.n346 B.n345 163.367
R751 B.n347 B.n346 163.367
R752 B.n347 B.n80 163.367
R753 B.n351 B.n80 163.367
R754 B.n352 B.n351 163.367
R755 B.n353 B.n352 163.367
R756 B.n353 B.n78 163.367
R757 B.n357 B.n78 163.367
R758 B.n358 B.n357 163.367
R759 B.n359 B.n358 163.367
R760 B.n359 B.n76 163.367
R761 B.n363 B.n76 163.367
R762 B.n364 B.n363 163.367
R763 B.n365 B.n364 163.367
R764 B.n365 B.n74 163.367
R765 B.n369 B.n74 163.367
R766 B.n370 B.n369 163.367
R767 B.n371 B.n370 163.367
R768 B.n371 B.n72 163.367
R769 B.n375 B.n72 163.367
R770 B.n376 B.n375 163.367
R771 B.n377 B.n376 163.367
R772 B.n377 B.n70 163.367
R773 B.n381 B.n70 163.367
R774 B.n382 B.n381 163.367
R775 B.n383 B.n382 163.367
R776 B.n383 B.n68 163.367
R777 B.n387 B.n68 163.367
R778 B.n388 B.n387 163.367
R779 B.n389 B.n388 163.367
R780 B.n389 B.n66 163.367
R781 B.n393 B.n66 163.367
R782 B.n394 B.n393 163.367
R783 B.n395 B.n394 163.367
R784 B.n395 B.n64 163.367
R785 B.n399 B.n64 163.367
R786 B.n400 B.n399 163.367
R787 B.n401 B.n400 163.367
R788 B.n401 B.n62 163.367
R789 B.n405 B.n62 163.367
R790 B.n406 B.n405 163.367
R791 B.n407 B.n406 163.367
R792 B.n407 B.n60 163.367
R793 B.n411 B.n60 163.367
R794 B.n412 B.n411 163.367
R795 B.n413 B.n412 163.367
R796 B.n413 B.n58 163.367
R797 B.n417 B.n58 163.367
R798 B.n418 B.n417 163.367
R799 B.n419 B.n418 163.367
R800 B.n419 B.n56 163.367
R801 B.n423 B.n56 163.367
R802 B.n424 B.n423 163.367
R803 B.n425 B.n424 163.367
R804 B.n425 B.n54 163.367
R805 B.n429 B.n54 163.367
R806 B.n430 B.n429 163.367
R807 B.n431 B.n430 163.367
R808 B.n431 B.n52 163.367
R809 B.n435 B.n52 163.367
R810 B.n436 B.n435 163.367
R811 B.n437 B.n436 163.367
R812 B.n437 B.n50 163.367
R813 B.n490 B.n29 163.367
R814 B.n486 B.n29 163.367
R815 B.n486 B.n485 163.367
R816 B.n485 B.n484 163.367
R817 B.n484 B.n31 163.367
R818 B.n480 B.n31 163.367
R819 B.n480 B.n479 163.367
R820 B.n479 B.n478 163.367
R821 B.n478 B.n33 163.367
R822 B.n474 B.n33 163.367
R823 B.n474 B.n473 163.367
R824 B.n473 B.n472 163.367
R825 B.n472 B.n35 163.367
R826 B.n468 B.n35 163.367
R827 B.n468 B.n467 163.367
R828 B.n467 B.n466 163.367
R829 B.n466 B.n40 163.367
R830 B.n462 B.n40 163.367
R831 B.n462 B.n461 163.367
R832 B.n461 B.n460 163.367
R833 B.n460 B.n42 163.367
R834 B.n455 B.n42 163.367
R835 B.n455 B.n454 163.367
R836 B.n454 B.n453 163.367
R837 B.n453 B.n46 163.367
R838 B.n449 B.n46 163.367
R839 B.n449 B.n448 163.367
R840 B.n448 B.n447 163.367
R841 B.n447 B.n48 163.367
R842 B.n443 B.n48 163.367
R843 B.n443 B.n442 163.367
R844 B.n442 B.n441 163.367
R845 B.n258 B.n257 73.6975
R846 B.n116 B.n115 73.6975
R847 B.n37 B.n36 73.6975
R848 B.n44 B.n43 73.6975
R849 B.n259 B.n258 59.5399
R850 B.n244 B.n116 59.5399
R851 B.n38 B.n37 59.5399
R852 B.n458 B.n44 59.5399
R853 B.n489 B.n28 31.0639
R854 B.n440 B.n439 31.0639
R855 B.n278 B.n103 31.0639
R856 B.n226 B.n225 31.0639
R857 B B.n571 18.0485
R858 B.n489 B.n488 10.6151
R859 B.n488 B.n487 10.6151
R860 B.n487 B.n30 10.6151
R861 B.n483 B.n30 10.6151
R862 B.n483 B.n482 10.6151
R863 B.n482 B.n481 10.6151
R864 B.n481 B.n32 10.6151
R865 B.n477 B.n32 10.6151
R866 B.n477 B.n476 10.6151
R867 B.n476 B.n475 10.6151
R868 B.n475 B.n34 10.6151
R869 B.n471 B.n470 10.6151
R870 B.n470 B.n469 10.6151
R871 B.n469 B.n39 10.6151
R872 B.n465 B.n39 10.6151
R873 B.n465 B.n464 10.6151
R874 B.n464 B.n463 10.6151
R875 B.n463 B.n41 10.6151
R876 B.n459 B.n41 10.6151
R877 B.n457 B.n456 10.6151
R878 B.n456 B.n45 10.6151
R879 B.n452 B.n45 10.6151
R880 B.n452 B.n451 10.6151
R881 B.n451 B.n450 10.6151
R882 B.n450 B.n47 10.6151
R883 B.n446 B.n47 10.6151
R884 B.n446 B.n445 10.6151
R885 B.n445 B.n444 10.6151
R886 B.n444 B.n49 10.6151
R887 B.n440 B.n49 10.6151
R888 B.n282 B.n103 10.6151
R889 B.n283 B.n282 10.6151
R890 B.n284 B.n283 10.6151
R891 B.n284 B.n101 10.6151
R892 B.n288 B.n101 10.6151
R893 B.n289 B.n288 10.6151
R894 B.n290 B.n289 10.6151
R895 B.n290 B.n99 10.6151
R896 B.n294 B.n99 10.6151
R897 B.n295 B.n294 10.6151
R898 B.n296 B.n295 10.6151
R899 B.n296 B.n97 10.6151
R900 B.n300 B.n97 10.6151
R901 B.n301 B.n300 10.6151
R902 B.n302 B.n301 10.6151
R903 B.n302 B.n95 10.6151
R904 B.n306 B.n95 10.6151
R905 B.n307 B.n306 10.6151
R906 B.n308 B.n307 10.6151
R907 B.n308 B.n93 10.6151
R908 B.n312 B.n93 10.6151
R909 B.n313 B.n312 10.6151
R910 B.n314 B.n313 10.6151
R911 B.n314 B.n91 10.6151
R912 B.n318 B.n91 10.6151
R913 B.n319 B.n318 10.6151
R914 B.n320 B.n319 10.6151
R915 B.n320 B.n89 10.6151
R916 B.n324 B.n89 10.6151
R917 B.n325 B.n324 10.6151
R918 B.n326 B.n325 10.6151
R919 B.n326 B.n87 10.6151
R920 B.n330 B.n87 10.6151
R921 B.n331 B.n330 10.6151
R922 B.n332 B.n331 10.6151
R923 B.n332 B.n85 10.6151
R924 B.n336 B.n85 10.6151
R925 B.n337 B.n336 10.6151
R926 B.n338 B.n337 10.6151
R927 B.n338 B.n83 10.6151
R928 B.n342 B.n83 10.6151
R929 B.n343 B.n342 10.6151
R930 B.n344 B.n343 10.6151
R931 B.n344 B.n81 10.6151
R932 B.n348 B.n81 10.6151
R933 B.n349 B.n348 10.6151
R934 B.n350 B.n349 10.6151
R935 B.n350 B.n79 10.6151
R936 B.n354 B.n79 10.6151
R937 B.n355 B.n354 10.6151
R938 B.n356 B.n355 10.6151
R939 B.n356 B.n77 10.6151
R940 B.n360 B.n77 10.6151
R941 B.n361 B.n360 10.6151
R942 B.n362 B.n361 10.6151
R943 B.n362 B.n75 10.6151
R944 B.n366 B.n75 10.6151
R945 B.n367 B.n366 10.6151
R946 B.n368 B.n367 10.6151
R947 B.n368 B.n73 10.6151
R948 B.n372 B.n73 10.6151
R949 B.n373 B.n372 10.6151
R950 B.n374 B.n373 10.6151
R951 B.n374 B.n71 10.6151
R952 B.n378 B.n71 10.6151
R953 B.n379 B.n378 10.6151
R954 B.n380 B.n379 10.6151
R955 B.n380 B.n69 10.6151
R956 B.n384 B.n69 10.6151
R957 B.n385 B.n384 10.6151
R958 B.n386 B.n385 10.6151
R959 B.n386 B.n67 10.6151
R960 B.n390 B.n67 10.6151
R961 B.n391 B.n390 10.6151
R962 B.n392 B.n391 10.6151
R963 B.n392 B.n65 10.6151
R964 B.n396 B.n65 10.6151
R965 B.n397 B.n396 10.6151
R966 B.n398 B.n397 10.6151
R967 B.n398 B.n63 10.6151
R968 B.n402 B.n63 10.6151
R969 B.n403 B.n402 10.6151
R970 B.n404 B.n403 10.6151
R971 B.n404 B.n61 10.6151
R972 B.n408 B.n61 10.6151
R973 B.n409 B.n408 10.6151
R974 B.n410 B.n409 10.6151
R975 B.n410 B.n59 10.6151
R976 B.n414 B.n59 10.6151
R977 B.n415 B.n414 10.6151
R978 B.n416 B.n415 10.6151
R979 B.n416 B.n57 10.6151
R980 B.n420 B.n57 10.6151
R981 B.n421 B.n420 10.6151
R982 B.n422 B.n421 10.6151
R983 B.n422 B.n55 10.6151
R984 B.n426 B.n55 10.6151
R985 B.n427 B.n426 10.6151
R986 B.n428 B.n427 10.6151
R987 B.n428 B.n53 10.6151
R988 B.n432 B.n53 10.6151
R989 B.n433 B.n432 10.6151
R990 B.n434 B.n433 10.6151
R991 B.n434 B.n51 10.6151
R992 B.n438 B.n51 10.6151
R993 B.n439 B.n438 10.6151
R994 B.n226 B.n121 10.6151
R995 B.n230 B.n121 10.6151
R996 B.n231 B.n230 10.6151
R997 B.n232 B.n231 10.6151
R998 B.n232 B.n119 10.6151
R999 B.n236 B.n119 10.6151
R1000 B.n237 B.n236 10.6151
R1001 B.n238 B.n237 10.6151
R1002 B.n238 B.n117 10.6151
R1003 B.n242 B.n117 10.6151
R1004 B.n243 B.n242 10.6151
R1005 B.n245 B.n113 10.6151
R1006 B.n249 B.n113 10.6151
R1007 B.n250 B.n249 10.6151
R1008 B.n251 B.n250 10.6151
R1009 B.n251 B.n111 10.6151
R1010 B.n255 B.n111 10.6151
R1011 B.n256 B.n255 10.6151
R1012 B.n260 B.n256 10.6151
R1013 B.n264 B.n109 10.6151
R1014 B.n265 B.n264 10.6151
R1015 B.n266 B.n265 10.6151
R1016 B.n266 B.n107 10.6151
R1017 B.n270 B.n107 10.6151
R1018 B.n271 B.n270 10.6151
R1019 B.n272 B.n271 10.6151
R1020 B.n272 B.n105 10.6151
R1021 B.n276 B.n105 10.6151
R1022 B.n277 B.n276 10.6151
R1023 B.n278 B.n277 10.6151
R1024 B.n225 B.n224 10.6151
R1025 B.n224 B.n123 10.6151
R1026 B.n220 B.n123 10.6151
R1027 B.n220 B.n219 10.6151
R1028 B.n219 B.n218 10.6151
R1029 B.n218 B.n125 10.6151
R1030 B.n214 B.n125 10.6151
R1031 B.n214 B.n213 10.6151
R1032 B.n213 B.n212 10.6151
R1033 B.n212 B.n127 10.6151
R1034 B.n208 B.n127 10.6151
R1035 B.n208 B.n207 10.6151
R1036 B.n207 B.n206 10.6151
R1037 B.n206 B.n129 10.6151
R1038 B.n202 B.n129 10.6151
R1039 B.n202 B.n201 10.6151
R1040 B.n201 B.n200 10.6151
R1041 B.n200 B.n131 10.6151
R1042 B.n196 B.n131 10.6151
R1043 B.n196 B.n195 10.6151
R1044 B.n195 B.n194 10.6151
R1045 B.n194 B.n133 10.6151
R1046 B.n190 B.n133 10.6151
R1047 B.n190 B.n189 10.6151
R1048 B.n189 B.n188 10.6151
R1049 B.n188 B.n135 10.6151
R1050 B.n184 B.n135 10.6151
R1051 B.n184 B.n183 10.6151
R1052 B.n183 B.n182 10.6151
R1053 B.n182 B.n137 10.6151
R1054 B.n178 B.n137 10.6151
R1055 B.n178 B.n177 10.6151
R1056 B.n177 B.n176 10.6151
R1057 B.n176 B.n139 10.6151
R1058 B.n172 B.n139 10.6151
R1059 B.n172 B.n171 10.6151
R1060 B.n171 B.n170 10.6151
R1061 B.n170 B.n141 10.6151
R1062 B.n166 B.n141 10.6151
R1063 B.n166 B.n165 10.6151
R1064 B.n165 B.n164 10.6151
R1065 B.n164 B.n143 10.6151
R1066 B.n160 B.n143 10.6151
R1067 B.n160 B.n159 10.6151
R1068 B.n159 B.n158 10.6151
R1069 B.n158 B.n145 10.6151
R1070 B.n154 B.n145 10.6151
R1071 B.n154 B.n153 10.6151
R1072 B.n153 B.n152 10.6151
R1073 B.n152 B.n147 10.6151
R1074 B.n148 B.n147 10.6151
R1075 B.n148 B.n0 10.6151
R1076 B.n567 B.n1 10.6151
R1077 B.n567 B.n566 10.6151
R1078 B.n566 B.n565 10.6151
R1079 B.n565 B.n4 10.6151
R1080 B.n561 B.n4 10.6151
R1081 B.n561 B.n560 10.6151
R1082 B.n560 B.n559 10.6151
R1083 B.n559 B.n6 10.6151
R1084 B.n555 B.n6 10.6151
R1085 B.n555 B.n554 10.6151
R1086 B.n554 B.n553 10.6151
R1087 B.n553 B.n8 10.6151
R1088 B.n549 B.n8 10.6151
R1089 B.n549 B.n548 10.6151
R1090 B.n548 B.n547 10.6151
R1091 B.n547 B.n10 10.6151
R1092 B.n543 B.n10 10.6151
R1093 B.n543 B.n542 10.6151
R1094 B.n542 B.n541 10.6151
R1095 B.n541 B.n12 10.6151
R1096 B.n537 B.n12 10.6151
R1097 B.n537 B.n536 10.6151
R1098 B.n536 B.n535 10.6151
R1099 B.n535 B.n14 10.6151
R1100 B.n531 B.n14 10.6151
R1101 B.n531 B.n530 10.6151
R1102 B.n530 B.n529 10.6151
R1103 B.n529 B.n16 10.6151
R1104 B.n525 B.n16 10.6151
R1105 B.n525 B.n524 10.6151
R1106 B.n524 B.n523 10.6151
R1107 B.n523 B.n18 10.6151
R1108 B.n519 B.n18 10.6151
R1109 B.n519 B.n518 10.6151
R1110 B.n518 B.n517 10.6151
R1111 B.n517 B.n20 10.6151
R1112 B.n513 B.n20 10.6151
R1113 B.n513 B.n512 10.6151
R1114 B.n512 B.n511 10.6151
R1115 B.n511 B.n22 10.6151
R1116 B.n507 B.n22 10.6151
R1117 B.n507 B.n506 10.6151
R1118 B.n506 B.n505 10.6151
R1119 B.n505 B.n24 10.6151
R1120 B.n501 B.n24 10.6151
R1121 B.n501 B.n500 10.6151
R1122 B.n500 B.n499 10.6151
R1123 B.n499 B.n26 10.6151
R1124 B.n495 B.n26 10.6151
R1125 B.n495 B.n494 10.6151
R1126 B.n494 B.n493 10.6151
R1127 B.n493 B.n28 10.6151
R1128 B.n471 B.n38 6.5566
R1129 B.n459 B.n458 6.5566
R1130 B.n245 B.n244 6.5566
R1131 B.n260 B.n259 6.5566
R1132 B.n38 B.n34 4.05904
R1133 B.n458 B.n457 4.05904
R1134 B.n244 B.n243 4.05904
R1135 B.n259 B.n109 4.05904
R1136 B.n571 B.n0 2.81026
R1137 B.n571 B.n1 2.81026
C0 w_n4010_n1338# VDD1 1.80003f
C1 VDD1 VTAIL 4.68199f
C2 B w_n4010_n1338# 8.10208f
C3 VP VDD1 1.80936f
C4 VDD1 VN 0.15849f
C5 B VTAIL 1.49876f
C6 B VP 2.08478f
C7 B VN 1.21157f
C8 w_n4010_n1338# VTAIL 1.62112f
C9 VP w_n4010_n1338# 8.14054f
C10 w_n4010_n1338# VN 7.62477f
C11 VDD1 VDD2 1.74532f
C12 VP VTAIL 2.61583f
C13 VTAIL VN 2.6017f
C14 B VDD2 1.59822f
C15 VP VN 5.89854f
C16 w_n4010_n1338# VDD2 1.91215f
C17 VDD2 VTAIL 4.74115f
C18 VP VDD2 0.539274f
C19 VDD2 VN 1.43178f
C20 B VDD1 1.50279f
C21 VDD2 VSUBS 1.220427f
C22 VDD1 VSUBS 1.598405f
C23 VTAIL VSUBS 0.625187f
C24 VN VSUBS 6.75643f
C25 VP VSUBS 3.013931f
C26 B VSUBS 4.361547f
C27 w_n4010_n1338# VSUBS 68.57101f
C28 B.n0 VSUBS 0.007146f
C29 B.n1 VSUBS 0.007146f
C30 B.n2 VSUBS 0.0113f
C31 B.n3 VSUBS 0.0113f
C32 B.n4 VSUBS 0.0113f
C33 B.n5 VSUBS 0.0113f
C34 B.n6 VSUBS 0.0113f
C35 B.n7 VSUBS 0.0113f
C36 B.n8 VSUBS 0.0113f
C37 B.n9 VSUBS 0.0113f
C38 B.n10 VSUBS 0.0113f
C39 B.n11 VSUBS 0.0113f
C40 B.n12 VSUBS 0.0113f
C41 B.n13 VSUBS 0.0113f
C42 B.n14 VSUBS 0.0113f
C43 B.n15 VSUBS 0.0113f
C44 B.n16 VSUBS 0.0113f
C45 B.n17 VSUBS 0.0113f
C46 B.n18 VSUBS 0.0113f
C47 B.n19 VSUBS 0.0113f
C48 B.n20 VSUBS 0.0113f
C49 B.n21 VSUBS 0.0113f
C50 B.n22 VSUBS 0.0113f
C51 B.n23 VSUBS 0.0113f
C52 B.n24 VSUBS 0.0113f
C53 B.n25 VSUBS 0.0113f
C54 B.n26 VSUBS 0.0113f
C55 B.n27 VSUBS 0.0113f
C56 B.n28 VSUBS 0.025199f
C57 B.n29 VSUBS 0.0113f
C58 B.n30 VSUBS 0.0113f
C59 B.n31 VSUBS 0.0113f
C60 B.n32 VSUBS 0.0113f
C61 B.n33 VSUBS 0.0113f
C62 B.n34 VSUBS 0.007811f
C63 B.n35 VSUBS 0.0113f
C64 B.t2 VSUBS 0.050671f
C65 B.t1 VSUBS 0.072338f
C66 B.t0 VSUBS 0.521084f
C67 B.n36 VSUBS 0.131128f
C68 B.n37 VSUBS 0.109942f
C69 B.n38 VSUBS 0.026182f
C70 B.n39 VSUBS 0.0113f
C71 B.n40 VSUBS 0.0113f
C72 B.n41 VSUBS 0.0113f
C73 B.n42 VSUBS 0.0113f
C74 B.t5 VSUBS 0.050671f
C75 B.t4 VSUBS 0.072338f
C76 B.t3 VSUBS 0.521084f
C77 B.n43 VSUBS 0.131128f
C78 B.n44 VSUBS 0.109942f
C79 B.n45 VSUBS 0.0113f
C80 B.n46 VSUBS 0.0113f
C81 B.n47 VSUBS 0.0113f
C82 B.n48 VSUBS 0.0113f
C83 B.n49 VSUBS 0.0113f
C84 B.n50 VSUBS 0.025199f
C85 B.n51 VSUBS 0.0113f
C86 B.n52 VSUBS 0.0113f
C87 B.n53 VSUBS 0.0113f
C88 B.n54 VSUBS 0.0113f
C89 B.n55 VSUBS 0.0113f
C90 B.n56 VSUBS 0.0113f
C91 B.n57 VSUBS 0.0113f
C92 B.n58 VSUBS 0.0113f
C93 B.n59 VSUBS 0.0113f
C94 B.n60 VSUBS 0.0113f
C95 B.n61 VSUBS 0.0113f
C96 B.n62 VSUBS 0.0113f
C97 B.n63 VSUBS 0.0113f
C98 B.n64 VSUBS 0.0113f
C99 B.n65 VSUBS 0.0113f
C100 B.n66 VSUBS 0.0113f
C101 B.n67 VSUBS 0.0113f
C102 B.n68 VSUBS 0.0113f
C103 B.n69 VSUBS 0.0113f
C104 B.n70 VSUBS 0.0113f
C105 B.n71 VSUBS 0.0113f
C106 B.n72 VSUBS 0.0113f
C107 B.n73 VSUBS 0.0113f
C108 B.n74 VSUBS 0.0113f
C109 B.n75 VSUBS 0.0113f
C110 B.n76 VSUBS 0.0113f
C111 B.n77 VSUBS 0.0113f
C112 B.n78 VSUBS 0.0113f
C113 B.n79 VSUBS 0.0113f
C114 B.n80 VSUBS 0.0113f
C115 B.n81 VSUBS 0.0113f
C116 B.n82 VSUBS 0.0113f
C117 B.n83 VSUBS 0.0113f
C118 B.n84 VSUBS 0.0113f
C119 B.n85 VSUBS 0.0113f
C120 B.n86 VSUBS 0.0113f
C121 B.n87 VSUBS 0.0113f
C122 B.n88 VSUBS 0.0113f
C123 B.n89 VSUBS 0.0113f
C124 B.n90 VSUBS 0.0113f
C125 B.n91 VSUBS 0.0113f
C126 B.n92 VSUBS 0.0113f
C127 B.n93 VSUBS 0.0113f
C128 B.n94 VSUBS 0.0113f
C129 B.n95 VSUBS 0.0113f
C130 B.n96 VSUBS 0.0113f
C131 B.n97 VSUBS 0.0113f
C132 B.n98 VSUBS 0.0113f
C133 B.n99 VSUBS 0.0113f
C134 B.n100 VSUBS 0.0113f
C135 B.n101 VSUBS 0.0113f
C136 B.n102 VSUBS 0.0113f
C137 B.n103 VSUBS 0.025199f
C138 B.n104 VSUBS 0.0113f
C139 B.n105 VSUBS 0.0113f
C140 B.n106 VSUBS 0.0113f
C141 B.n107 VSUBS 0.0113f
C142 B.n108 VSUBS 0.0113f
C143 B.n109 VSUBS 0.007811f
C144 B.n110 VSUBS 0.0113f
C145 B.n111 VSUBS 0.0113f
C146 B.n112 VSUBS 0.0113f
C147 B.n113 VSUBS 0.0113f
C148 B.n114 VSUBS 0.0113f
C149 B.t7 VSUBS 0.050671f
C150 B.t8 VSUBS 0.072338f
C151 B.t6 VSUBS 0.521084f
C152 B.n115 VSUBS 0.131128f
C153 B.n116 VSUBS 0.109942f
C154 B.n117 VSUBS 0.0113f
C155 B.n118 VSUBS 0.0113f
C156 B.n119 VSUBS 0.0113f
C157 B.n120 VSUBS 0.0113f
C158 B.n121 VSUBS 0.0113f
C159 B.n122 VSUBS 0.025199f
C160 B.n123 VSUBS 0.0113f
C161 B.n124 VSUBS 0.0113f
C162 B.n125 VSUBS 0.0113f
C163 B.n126 VSUBS 0.0113f
C164 B.n127 VSUBS 0.0113f
C165 B.n128 VSUBS 0.0113f
C166 B.n129 VSUBS 0.0113f
C167 B.n130 VSUBS 0.0113f
C168 B.n131 VSUBS 0.0113f
C169 B.n132 VSUBS 0.0113f
C170 B.n133 VSUBS 0.0113f
C171 B.n134 VSUBS 0.0113f
C172 B.n135 VSUBS 0.0113f
C173 B.n136 VSUBS 0.0113f
C174 B.n137 VSUBS 0.0113f
C175 B.n138 VSUBS 0.0113f
C176 B.n139 VSUBS 0.0113f
C177 B.n140 VSUBS 0.0113f
C178 B.n141 VSUBS 0.0113f
C179 B.n142 VSUBS 0.0113f
C180 B.n143 VSUBS 0.0113f
C181 B.n144 VSUBS 0.0113f
C182 B.n145 VSUBS 0.0113f
C183 B.n146 VSUBS 0.0113f
C184 B.n147 VSUBS 0.0113f
C185 B.n148 VSUBS 0.0113f
C186 B.n149 VSUBS 0.0113f
C187 B.n150 VSUBS 0.0113f
C188 B.n151 VSUBS 0.0113f
C189 B.n152 VSUBS 0.0113f
C190 B.n153 VSUBS 0.0113f
C191 B.n154 VSUBS 0.0113f
C192 B.n155 VSUBS 0.0113f
C193 B.n156 VSUBS 0.0113f
C194 B.n157 VSUBS 0.0113f
C195 B.n158 VSUBS 0.0113f
C196 B.n159 VSUBS 0.0113f
C197 B.n160 VSUBS 0.0113f
C198 B.n161 VSUBS 0.0113f
C199 B.n162 VSUBS 0.0113f
C200 B.n163 VSUBS 0.0113f
C201 B.n164 VSUBS 0.0113f
C202 B.n165 VSUBS 0.0113f
C203 B.n166 VSUBS 0.0113f
C204 B.n167 VSUBS 0.0113f
C205 B.n168 VSUBS 0.0113f
C206 B.n169 VSUBS 0.0113f
C207 B.n170 VSUBS 0.0113f
C208 B.n171 VSUBS 0.0113f
C209 B.n172 VSUBS 0.0113f
C210 B.n173 VSUBS 0.0113f
C211 B.n174 VSUBS 0.0113f
C212 B.n175 VSUBS 0.0113f
C213 B.n176 VSUBS 0.0113f
C214 B.n177 VSUBS 0.0113f
C215 B.n178 VSUBS 0.0113f
C216 B.n179 VSUBS 0.0113f
C217 B.n180 VSUBS 0.0113f
C218 B.n181 VSUBS 0.0113f
C219 B.n182 VSUBS 0.0113f
C220 B.n183 VSUBS 0.0113f
C221 B.n184 VSUBS 0.0113f
C222 B.n185 VSUBS 0.0113f
C223 B.n186 VSUBS 0.0113f
C224 B.n187 VSUBS 0.0113f
C225 B.n188 VSUBS 0.0113f
C226 B.n189 VSUBS 0.0113f
C227 B.n190 VSUBS 0.0113f
C228 B.n191 VSUBS 0.0113f
C229 B.n192 VSUBS 0.0113f
C230 B.n193 VSUBS 0.0113f
C231 B.n194 VSUBS 0.0113f
C232 B.n195 VSUBS 0.0113f
C233 B.n196 VSUBS 0.0113f
C234 B.n197 VSUBS 0.0113f
C235 B.n198 VSUBS 0.0113f
C236 B.n199 VSUBS 0.0113f
C237 B.n200 VSUBS 0.0113f
C238 B.n201 VSUBS 0.0113f
C239 B.n202 VSUBS 0.0113f
C240 B.n203 VSUBS 0.0113f
C241 B.n204 VSUBS 0.0113f
C242 B.n205 VSUBS 0.0113f
C243 B.n206 VSUBS 0.0113f
C244 B.n207 VSUBS 0.0113f
C245 B.n208 VSUBS 0.0113f
C246 B.n209 VSUBS 0.0113f
C247 B.n210 VSUBS 0.0113f
C248 B.n211 VSUBS 0.0113f
C249 B.n212 VSUBS 0.0113f
C250 B.n213 VSUBS 0.0113f
C251 B.n214 VSUBS 0.0113f
C252 B.n215 VSUBS 0.0113f
C253 B.n216 VSUBS 0.0113f
C254 B.n217 VSUBS 0.0113f
C255 B.n218 VSUBS 0.0113f
C256 B.n219 VSUBS 0.0113f
C257 B.n220 VSUBS 0.0113f
C258 B.n221 VSUBS 0.0113f
C259 B.n222 VSUBS 0.0113f
C260 B.n223 VSUBS 0.0113f
C261 B.n224 VSUBS 0.0113f
C262 B.n225 VSUBS 0.025199f
C263 B.n226 VSUBS 0.025986f
C264 B.n227 VSUBS 0.025986f
C265 B.n228 VSUBS 0.0113f
C266 B.n229 VSUBS 0.0113f
C267 B.n230 VSUBS 0.0113f
C268 B.n231 VSUBS 0.0113f
C269 B.n232 VSUBS 0.0113f
C270 B.n233 VSUBS 0.0113f
C271 B.n234 VSUBS 0.0113f
C272 B.n235 VSUBS 0.0113f
C273 B.n236 VSUBS 0.0113f
C274 B.n237 VSUBS 0.0113f
C275 B.n238 VSUBS 0.0113f
C276 B.n239 VSUBS 0.0113f
C277 B.n240 VSUBS 0.0113f
C278 B.n241 VSUBS 0.0113f
C279 B.n242 VSUBS 0.0113f
C280 B.n243 VSUBS 0.007811f
C281 B.n244 VSUBS 0.026182f
C282 B.n245 VSUBS 0.00914f
C283 B.n246 VSUBS 0.0113f
C284 B.n247 VSUBS 0.0113f
C285 B.n248 VSUBS 0.0113f
C286 B.n249 VSUBS 0.0113f
C287 B.n250 VSUBS 0.0113f
C288 B.n251 VSUBS 0.0113f
C289 B.n252 VSUBS 0.0113f
C290 B.n253 VSUBS 0.0113f
C291 B.n254 VSUBS 0.0113f
C292 B.n255 VSUBS 0.0113f
C293 B.n256 VSUBS 0.0113f
C294 B.t10 VSUBS 0.050671f
C295 B.t11 VSUBS 0.072338f
C296 B.t9 VSUBS 0.521084f
C297 B.n257 VSUBS 0.131128f
C298 B.n258 VSUBS 0.109942f
C299 B.n259 VSUBS 0.026182f
C300 B.n260 VSUBS 0.00914f
C301 B.n261 VSUBS 0.0113f
C302 B.n262 VSUBS 0.0113f
C303 B.n263 VSUBS 0.0113f
C304 B.n264 VSUBS 0.0113f
C305 B.n265 VSUBS 0.0113f
C306 B.n266 VSUBS 0.0113f
C307 B.n267 VSUBS 0.0113f
C308 B.n268 VSUBS 0.0113f
C309 B.n269 VSUBS 0.0113f
C310 B.n270 VSUBS 0.0113f
C311 B.n271 VSUBS 0.0113f
C312 B.n272 VSUBS 0.0113f
C313 B.n273 VSUBS 0.0113f
C314 B.n274 VSUBS 0.0113f
C315 B.n275 VSUBS 0.0113f
C316 B.n276 VSUBS 0.0113f
C317 B.n277 VSUBS 0.0113f
C318 B.n278 VSUBS 0.025986f
C319 B.n279 VSUBS 0.025986f
C320 B.n280 VSUBS 0.025199f
C321 B.n281 VSUBS 0.0113f
C322 B.n282 VSUBS 0.0113f
C323 B.n283 VSUBS 0.0113f
C324 B.n284 VSUBS 0.0113f
C325 B.n285 VSUBS 0.0113f
C326 B.n286 VSUBS 0.0113f
C327 B.n287 VSUBS 0.0113f
C328 B.n288 VSUBS 0.0113f
C329 B.n289 VSUBS 0.0113f
C330 B.n290 VSUBS 0.0113f
C331 B.n291 VSUBS 0.0113f
C332 B.n292 VSUBS 0.0113f
C333 B.n293 VSUBS 0.0113f
C334 B.n294 VSUBS 0.0113f
C335 B.n295 VSUBS 0.0113f
C336 B.n296 VSUBS 0.0113f
C337 B.n297 VSUBS 0.0113f
C338 B.n298 VSUBS 0.0113f
C339 B.n299 VSUBS 0.0113f
C340 B.n300 VSUBS 0.0113f
C341 B.n301 VSUBS 0.0113f
C342 B.n302 VSUBS 0.0113f
C343 B.n303 VSUBS 0.0113f
C344 B.n304 VSUBS 0.0113f
C345 B.n305 VSUBS 0.0113f
C346 B.n306 VSUBS 0.0113f
C347 B.n307 VSUBS 0.0113f
C348 B.n308 VSUBS 0.0113f
C349 B.n309 VSUBS 0.0113f
C350 B.n310 VSUBS 0.0113f
C351 B.n311 VSUBS 0.0113f
C352 B.n312 VSUBS 0.0113f
C353 B.n313 VSUBS 0.0113f
C354 B.n314 VSUBS 0.0113f
C355 B.n315 VSUBS 0.0113f
C356 B.n316 VSUBS 0.0113f
C357 B.n317 VSUBS 0.0113f
C358 B.n318 VSUBS 0.0113f
C359 B.n319 VSUBS 0.0113f
C360 B.n320 VSUBS 0.0113f
C361 B.n321 VSUBS 0.0113f
C362 B.n322 VSUBS 0.0113f
C363 B.n323 VSUBS 0.0113f
C364 B.n324 VSUBS 0.0113f
C365 B.n325 VSUBS 0.0113f
C366 B.n326 VSUBS 0.0113f
C367 B.n327 VSUBS 0.0113f
C368 B.n328 VSUBS 0.0113f
C369 B.n329 VSUBS 0.0113f
C370 B.n330 VSUBS 0.0113f
C371 B.n331 VSUBS 0.0113f
C372 B.n332 VSUBS 0.0113f
C373 B.n333 VSUBS 0.0113f
C374 B.n334 VSUBS 0.0113f
C375 B.n335 VSUBS 0.0113f
C376 B.n336 VSUBS 0.0113f
C377 B.n337 VSUBS 0.0113f
C378 B.n338 VSUBS 0.0113f
C379 B.n339 VSUBS 0.0113f
C380 B.n340 VSUBS 0.0113f
C381 B.n341 VSUBS 0.0113f
C382 B.n342 VSUBS 0.0113f
C383 B.n343 VSUBS 0.0113f
C384 B.n344 VSUBS 0.0113f
C385 B.n345 VSUBS 0.0113f
C386 B.n346 VSUBS 0.0113f
C387 B.n347 VSUBS 0.0113f
C388 B.n348 VSUBS 0.0113f
C389 B.n349 VSUBS 0.0113f
C390 B.n350 VSUBS 0.0113f
C391 B.n351 VSUBS 0.0113f
C392 B.n352 VSUBS 0.0113f
C393 B.n353 VSUBS 0.0113f
C394 B.n354 VSUBS 0.0113f
C395 B.n355 VSUBS 0.0113f
C396 B.n356 VSUBS 0.0113f
C397 B.n357 VSUBS 0.0113f
C398 B.n358 VSUBS 0.0113f
C399 B.n359 VSUBS 0.0113f
C400 B.n360 VSUBS 0.0113f
C401 B.n361 VSUBS 0.0113f
C402 B.n362 VSUBS 0.0113f
C403 B.n363 VSUBS 0.0113f
C404 B.n364 VSUBS 0.0113f
C405 B.n365 VSUBS 0.0113f
C406 B.n366 VSUBS 0.0113f
C407 B.n367 VSUBS 0.0113f
C408 B.n368 VSUBS 0.0113f
C409 B.n369 VSUBS 0.0113f
C410 B.n370 VSUBS 0.0113f
C411 B.n371 VSUBS 0.0113f
C412 B.n372 VSUBS 0.0113f
C413 B.n373 VSUBS 0.0113f
C414 B.n374 VSUBS 0.0113f
C415 B.n375 VSUBS 0.0113f
C416 B.n376 VSUBS 0.0113f
C417 B.n377 VSUBS 0.0113f
C418 B.n378 VSUBS 0.0113f
C419 B.n379 VSUBS 0.0113f
C420 B.n380 VSUBS 0.0113f
C421 B.n381 VSUBS 0.0113f
C422 B.n382 VSUBS 0.0113f
C423 B.n383 VSUBS 0.0113f
C424 B.n384 VSUBS 0.0113f
C425 B.n385 VSUBS 0.0113f
C426 B.n386 VSUBS 0.0113f
C427 B.n387 VSUBS 0.0113f
C428 B.n388 VSUBS 0.0113f
C429 B.n389 VSUBS 0.0113f
C430 B.n390 VSUBS 0.0113f
C431 B.n391 VSUBS 0.0113f
C432 B.n392 VSUBS 0.0113f
C433 B.n393 VSUBS 0.0113f
C434 B.n394 VSUBS 0.0113f
C435 B.n395 VSUBS 0.0113f
C436 B.n396 VSUBS 0.0113f
C437 B.n397 VSUBS 0.0113f
C438 B.n398 VSUBS 0.0113f
C439 B.n399 VSUBS 0.0113f
C440 B.n400 VSUBS 0.0113f
C441 B.n401 VSUBS 0.0113f
C442 B.n402 VSUBS 0.0113f
C443 B.n403 VSUBS 0.0113f
C444 B.n404 VSUBS 0.0113f
C445 B.n405 VSUBS 0.0113f
C446 B.n406 VSUBS 0.0113f
C447 B.n407 VSUBS 0.0113f
C448 B.n408 VSUBS 0.0113f
C449 B.n409 VSUBS 0.0113f
C450 B.n410 VSUBS 0.0113f
C451 B.n411 VSUBS 0.0113f
C452 B.n412 VSUBS 0.0113f
C453 B.n413 VSUBS 0.0113f
C454 B.n414 VSUBS 0.0113f
C455 B.n415 VSUBS 0.0113f
C456 B.n416 VSUBS 0.0113f
C457 B.n417 VSUBS 0.0113f
C458 B.n418 VSUBS 0.0113f
C459 B.n419 VSUBS 0.0113f
C460 B.n420 VSUBS 0.0113f
C461 B.n421 VSUBS 0.0113f
C462 B.n422 VSUBS 0.0113f
C463 B.n423 VSUBS 0.0113f
C464 B.n424 VSUBS 0.0113f
C465 B.n425 VSUBS 0.0113f
C466 B.n426 VSUBS 0.0113f
C467 B.n427 VSUBS 0.0113f
C468 B.n428 VSUBS 0.0113f
C469 B.n429 VSUBS 0.0113f
C470 B.n430 VSUBS 0.0113f
C471 B.n431 VSUBS 0.0113f
C472 B.n432 VSUBS 0.0113f
C473 B.n433 VSUBS 0.0113f
C474 B.n434 VSUBS 0.0113f
C475 B.n435 VSUBS 0.0113f
C476 B.n436 VSUBS 0.0113f
C477 B.n437 VSUBS 0.0113f
C478 B.n438 VSUBS 0.0113f
C479 B.n439 VSUBS 0.026602f
C480 B.n440 VSUBS 0.024582f
C481 B.n441 VSUBS 0.025986f
C482 B.n442 VSUBS 0.0113f
C483 B.n443 VSUBS 0.0113f
C484 B.n444 VSUBS 0.0113f
C485 B.n445 VSUBS 0.0113f
C486 B.n446 VSUBS 0.0113f
C487 B.n447 VSUBS 0.0113f
C488 B.n448 VSUBS 0.0113f
C489 B.n449 VSUBS 0.0113f
C490 B.n450 VSUBS 0.0113f
C491 B.n451 VSUBS 0.0113f
C492 B.n452 VSUBS 0.0113f
C493 B.n453 VSUBS 0.0113f
C494 B.n454 VSUBS 0.0113f
C495 B.n455 VSUBS 0.0113f
C496 B.n456 VSUBS 0.0113f
C497 B.n457 VSUBS 0.007811f
C498 B.n458 VSUBS 0.026182f
C499 B.n459 VSUBS 0.00914f
C500 B.n460 VSUBS 0.0113f
C501 B.n461 VSUBS 0.0113f
C502 B.n462 VSUBS 0.0113f
C503 B.n463 VSUBS 0.0113f
C504 B.n464 VSUBS 0.0113f
C505 B.n465 VSUBS 0.0113f
C506 B.n466 VSUBS 0.0113f
C507 B.n467 VSUBS 0.0113f
C508 B.n468 VSUBS 0.0113f
C509 B.n469 VSUBS 0.0113f
C510 B.n470 VSUBS 0.0113f
C511 B.n471 VSUBS 0.00914f
C512 B.n472 VSUBS 0.0113f
C513 B.n473 VSUBS 0.0113f
C514 B.n474 VSUBS 0.0113f
C515 B.n475 VSUBS 0.0113f
C516 B.n476 VSUBS 0.0113f
C517 B.n477 VSUBS 0.0113f
C518 B.n478 VSUBS 0.0113f
C519 B.n479 VSUBS 0.0113f
C520 B.n480 VSUBS 0.0113f
C521 B.n481 VSUBS 0.0113f
C522 B.n482 VSUBS 0.0113f
C523 B.n483 VSUBS 0.0113f
C524 B.n484 VSUBS 0.0113f
C525 B.n485 VSUBS 0.0113f
C526 B.n486 VSUBS 0.0113f
C527 B.n487 VSUBS 0.0113f
C528 B.n488 VSUBS 0.0113f
C529 B.n489 VSUBS 0.025986f
C530 B.n490 VSUBS 0.025986f
C531 B.n491 VSUBS 0.025199f
C532 B.n492 VSUBS 0.0113f
C533 B.n493 VSUBS 0.0113f
C534 B.n494 VSUBS 0.0113f
C535 B.n495 VSUBS 0.0113f
C536 B.n496 VSUBS 0.0113f
C537 B.n497 VSUBS 0.0113f
C538 B.n498 VSUBS 0.0113f
C539 B.n499 VSUBS 0.0113f
C540 B.n500 VSUBS 0.0113f
C541 B.n501 VSUBS 0.0113f
C542 B.n502 VSUBS 0.0113f
C543 B.n503 VSUBS 0.0113f
C544 B.n504 VSUBS 0.0113f
C545 B.n505 VSUBS 0.0113f
C546 B.n506 VSUBS 0.0113f
C547 B.n507 VSUBS 0.0113f
C548 B.n508 VSUBS 0.0113f
C549 B.n509 VSUBS 0.0113f
C550 B.n510 VSUBS 0.0113f
C551 B.n511 VSUBS 0.0113f
C552 B.n512 VSUBS 0.0113f
C553 B.n513 VSUBS 0.0113f
C554 B.n514 VSUBS 0.0113f
C555 B.n515 VSUBS 0.0113f
C556 B.n516 VSUBS 0.0113f
C557 B.n517 VSUBS 0.0113f
C558 B.n518 VSUBS 0.0113f
C559 B.n519 VSUBS 0.0113f
C560 B.n520 VSUBS 0.0113f
C561 B.n521 VSUBS 0.0113f
C562 B.n522 VSUBS 0.0113f
C563 B.n523 VSUBS 0.0113f
C564 B.n524 VSUBS 0.0113f
C565 B.n525 VSUBS 0.0113f
C566 B.n526 VSUBS 0.0113f
C567 B.n527 VSUBS 0.0113f
C568 B.n528 VSUBS 0.0113f
C569 B.n529 VSUBS 0.0113f
C570 B.n530 VSUBS 0.0113f
C571 B.n531 VSUBS 0.0113f
C572 B.n532 VSUBS 0.0113f
C573 B.n533 VSUBS 0.0113f
C574 B.n534 VSUBS 0.0113f
C575 B.n535 VSUBS 0.0113f
C576 B.n536 VSUBS 0.0113f
C577 B.n537 VSUBS 0.0113f
C578 B.n538 VSUBS 0.0113f
C579 B.n539 VSUBS 0.0113f
C580 B.n540 VSUBS 0.0113f
C581 B.n541 VSUBS 0.0113f
C582 B.n542 VSUBS 0.0113f
C583 B.n543 VSUBS 0.0113f
C584 B.n544 VSUBS 0.0113f
C585 B.n545 VSUBS 0.0113f
C586 B.n546 VSUBS 0.0113f
C587 B.n547 VSUBS 0.0113f
C588 B.n548 VSUBS 0.0113f
C589 B.n549 VSUBS 0.0113f
C590 B.n550 VSUBS 0.0113f
C591 B.n551 VSUBS 0.0113f
C592 B.n552 VSUBS 0.0113f
C593 B.n553 VSUBS 0.0113f
C594 B.n554 VSUBS 0.0113f
C595 B.n555 VSUBS 0.0113f
C596 B.n556 VSUBS 0.0113f
C597 B.n557 VSUBS 0.0113f
C598 B.n558 VSUBS 0.0113f
C599 B.n559 VSUBS 0.0113f
C600 B.n560 VSUBS 0.0113f
C601 B.n561 VSUBS 0.0113f
C602 B.n562 VSUBS 0.0113f
C603 B.n563 VSUBS 0.0113f
C604 B.n564 VSUBS 0.0113f
C605 B.n565 VSUBS 0.0113f
C606 B.n566 VSUBS 0.0113f
C607 B.n567 VSUBS 0.0113f
C608 B.n568 VSUBS 0.0113f
C609 B.n569 VSUBS 0.0113f
C610 B.n570 VSUBS 0.0113f
C611 B.n571 VSUBS 0.025588f
C612 VDD1.n0 VSUBS 0.018238f
C613 VDD1.n1 VSUBS 0.048911f
C614 VDD1.t5 VSUBS 0.046938f
C615 VDD1.n2 VSUBS 0.045246f
C616 VDD1.n3 VSUBS 0.011553f
C617 VDD1.n4 VSUBS 0.009203f
C618 VDD1.n5 VSUBS 0.104329f
C619 VDD1.n6 VSUBS 0.045321f
C620 VDD1.n7 VSUBS 0.018238f
C621 VDD1.n8 VSUBS 0.048911f
C622 VDD1.t4 VSUBS 0.046938f
C623 VDD1.n9 VSUBS 0.045246f
C624 VDD1.n10 VSUBS 0.011553f
C625 VDD1.n11 VSUBS 0.009203f
C626 VDD1.n12 VSUBS 0.104329f
C627 VDD1.n13 VSUBS 0.044707f
C628 VDD1.t0 VSUBS 0.025037f
C629 VDD1.t2 VSUBS 0.025037f
C630 VDD1.n14 VSUBS 0.107675f
C631 VDD1.n15 VSUBS 1.80567f
C632 VDD1.t3 VSUBS 0.025037f
C633 VDD1.t1 VSUBS 0.025037f
C634 VDD1.n16 VSUBS 0.106153f
C635 VDD1.n17 VSUBS 1.57467f
C636 VP.t3 VSUBS 0.823948f
C637 VP.n0 VSUBS 0.616551f
C638 VP.n1 VSUBS 0.055865f
C639 VP.n2 VSUBS 0.052775f
C640 VP.n3 VSUBS 0.055865f
C641 VP.t5 VSUBS 0.823948f
C642 VP.n4 VSUBS 0.43913f
C643 VP.n5 VSUBS 0.055865f
C644 VP.n6 VSUBS 0.052775f
C645 VP.n7 VSUBS 0.055865f
C646 VP.t1 VSUBS 0.823948f
C647 VP.n8 VSUBS 0.616551f
C648 VP.t4 VSUBS 0.823948f
C649 VP.n9 VSUBS 0.616551f
C650 VP.n10 VSUBS 0.055865f
C651 VP.n11 VSUBS 0.052775f
C652 VP.n12 VSUBS 0.055865f
C653 VP.t2 VSUBS 0.823948f
C654 VP.n13 VSUBS 0.608768f
C655 VP.t0 VSUBS 1.41369f
C656 VP.n14 VSUBS 0.638171f
C657 VP.n15 VSUBS 0.682124f
C658 VP.n16 VSUBS 0.104118f
C659 VP.n17 VSUBS 0.104118f
C660 VP.n18 VSUBS 0.102532f
C661 VP.n19 VSUBS 0.055865f
C662 VP.n20 VSUBS 0.055865f
C663 VP.n21 VSUBS 0.055865f
C664 VP.n22 VSUBS 0.111917f
C665 VP.n23 VSUBS 0.104118f
C666 VP.n24 VSUBS 0.083557f
C667 VP.n25 VSUBS 0.090165f
C668 VP.n26 VSUBS 2.68764f
C669 VP.n27 VSUBS 2.73271f
C670 VP.n28 VSUBS 0.090165f
C671 VP.n29 VSUBS 0.083557f
C672 VP.n30 VSUBS 0.104118f
C673 VP.n31 VSUBS 0.111917f
C674 VP.n32 VSUBS 0.055865f
C675 VP.n33 VSUBS 0.055865f
C676 VP.n34 VSUBS 0.055865f
C677 VP.n35 VSUBS 0.102532f
C678 VP.n36 VSUBS 0.104118f
C679 VP.n37 VSUBS 0.104118f
C680 VP.n38 VSUBS 0.055865f
C681 VP.n39 VSUBS 0.055865f
C682 VP.n40 VSUBS 0.055865f
C683 VP.n41 VSUBS 0.104118f
C684 VP.n42 VSUBS 0.104118f
C685 VP.n43 VSUBS 0.102532f
C686 VP.n44 VSUBS 0.055865f
C687 VP.n45 VSUBS 0.055865f
C688 VP.n46 VSUBS 0.055865f
C689 VP.n47 VSUBS 0.111917f
C690 VP.n48 VSUBS 0.104118f
C691 VP.n49 VSUBS 0.083557f
C692 VP.n50 VSUBS 0.090165f
C693 VP.n51 VSUBS 0.139084f
C694 VTAIL.t10 VSUBS 0.053595f
C695 VTAIL.t6 VSUBS 0.053595f
C696 VTAIL.n0 VSUBS 0.194175f
C697 VTAIL.n1 VSUBS 0.711855f
C698 VTAIL.n2 VSUBS 0.039041f
C699 VTAIL.n3 VSUBS 0.104702f
C700 VTAIL.t5 VSUBS 0.100478f
C701 VTAIL.n4 VSUBS 0.096857f
C702 VTAIL.n5 VSUBS 0.02473f
C703 VTAIL.n6 VSUBS 0.0197f
C704 VTAIL.n7 VSUBS 0.223332f
C705 VTAIL.n8 VSUBS 0.054625f
C706 VTAIL.n9 VSUBS 0.672091f
C707 VTAIL.t3 VSUBS 0.053595f
C708 VTAIL.t4 VSUBS 0.053595f
C709 VTAIL.n10 VSUBS 0.194175f
C710 VTAIL.n11 VSUBS 2.20656f
C711 VTAIL.t8 VSUBS 0.053595f
C712 VTAIL.t11 VSUBS 0.053595f
C713 VTAIL.n12 VSUBS 0.194176f
C714 VTAIL.n13 VSUBS 2.20656f
C715 VTAIL.n14 VSUBS 0.039041f
C716 VTAIL.n15 VSUBS 0.104702f
C717 VTAIL.t9 VSUBS 0.100478f
C718 VTAIL.n16 VSUBS 0.096857f
C719 VTAIL.n17 VSUBS 0.02473f
C720 VTAIL.n18 VSUBS 0.0197f
C721 VTAIL.n19 VSUBS 0.223332f
C722 VTAIL.n20 VSUBS 0.054625f
C723 VTAIL.n21 VSUBS 0.672091f
C724 VTAIL.t0 VSUBS 0.053595f
C725 VTAIL.t2 VSUBS 0.053595f
C726 VTAIL.n22 VSUBS 0.194176f
C727 VTAIL.n23 VSUBS 0.995212f
C728 VTAIL.n24 VSUBS 0.039041f
C729 VTAIL.n25 VSUBS 0.104702f
C730 VTAIL.t1 VSUBS 0.100478f
C731 VTAIL.n26 VSUBS 0.096857f
C732 VTAIL.n27 VSUBS 0.02473f
C733 VTAIL.n28 VSUBS 0.0197f
C734 VTAIL.n29 VSUBS 0.223332f
C735 VTAIL.n30 VSUBS 0.054625f
C736 VTAIL.n31 VSUBS 1.49647f
C737 VTAIL.n32 VSUBS 0.039041f
C738 VTAIL.n33 VSUBS 0.104702f
C739 VTAIL.t7 VSUBS 0.100478f
C740 VTAIL.n34 VSUBS 0.096857f
C741 VTAIL.n35 VSUBS 0.02473f
C742 VTAIL.n36 VSUBS 0.0197f
C743 VTAIL.n37 VSUBS 0.223332f
C744 VTAIL.n38 VSUBS 0.054625f
C745 VTAIL.n39 VSUBS 1.39285f
C746 VDD2.n0 VSUBS 0.018487f
C747 VDD2.n1 VSUBS 0.049578f
C748 VDD2.t5 VSUBS 0.047578f
C749 VDD2.n2 VSUBS 0.045863f
C750 VDD2.n3 VSUBS 0.01171f
C751 VDD2.n4 VSUBS 0.009328f
C752 VDD2.n5 VSUBS 0.105752f
C753 VDD2.n6 VSUBS 0.045317f
C754 VDD2.t0 VSUBS 0.025378f
C755 VDD2.t1 VSUBS 0.025378f
C756 VDD2.n7 VSUBS 0.109144f
C757 VDD2.n8 VSUBS 1.73667f
C758 VDD2.n9 VSUBS 0.018487f
C759 VDD2.n10 VSUBS 0.049578f
C760 VDD2.t2 VSUBS 0.047578f
C761 VDD2.n11 VSUBS 0.045863f
C762 VDD2.n12 VSUBS 0.01171f
C763 VDD2.n13 VSUBS 0.009328f
C764 VDD2.n14 VSUBS 0.105752f
C765 VDD2.n15 VSUBS 0.037824f
C766 VDD2.n16 VSUBS 1.39126f
C767 VDD2.t4 VSUBS 0.025378f
C768 VDD2.t3 VSUBS 0.025378f
C769 VDD2.n17 VSUBS 0.109136f
C770 VN.t4 VSUBS 0.706422f
C771 VN.n0 VSUBS 0.528607f
C772 VN.n1 VSUBS 0.047897f
C773 VN.n2 VSUBS 0.045247f
C774 VN.n3 VSUBS 0.047897f
C775 VN.t5 VSUBS 0.706422f
C776 VN.n4 VSUBS 0.521934f
C777 VN.t1 VSUBS 1.21205f
C778 VN.n5 VSUBS 0.547143f
C779 VN.n6 VSUBS 0.584827f
C780 VN.n7 VSUBS 0.089267f
C781 VN.n8 VSUBS 0.089267f
C782 VN.n9 VSUBS 0.087908f
C783 VN.n10 VSUBS 0.047897f
C784 VN.n11 VSUBS 0.047897f
C785 VN.n12 VSUBS 0.047897f
C786 VN.n13 VSUBS 0.095953f
C787 VN.n14 VSUBS 0.089267f
C788 VN.n15 VSUBS 0.071638f
C789 VN.n16 VSUBS 0.077304f
C790 VN.n17 VSUBS 0.119245f
C791 VN.t3 VSUBS 0.706422f
C792 VN.n18 VSUBS 0.528607f
C793 VN.n19 VSUBS 0.047897f
C794 VN.n20 VSUBS 0.045247f
C795 VN.n21 VSUBS 0.047897f
C796 VN.t0 VSUBS 0.706422f
C797 VN.n22 VSUBS 0.521934f
C798 VN.t2 VSUBS 1.21205f
C799 VN.n23 VSUBS 0.547143f
C800 VN.n24 VSUBS 0.584827f
C801 VN.n25 VSUBS 0.089267f
C802 VN.n26 VSUBS 0.089267f
C803 VN.n27 VSUBS 0.087908f
C804 VN.n28 VSUBS 0.047897f
C805 VN.n29 VSUBS 0.047897f
C806 VN.n30 VSUBS 0.047897f
C807 VN.n31 VSUBS 0.095953f
C808 VN.n32 VSUBS 0.089267f
C809 VN.n33 VSUBS 0.071638f
C810 VN.n34 VSUBS 0.077304f
C811 VN.n35 VSUBS 2.32468f
.ends

