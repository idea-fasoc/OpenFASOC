* NGSPICE file created from diff_pair_sample_1236.ext - technology: sky130A

.subckt diff_pair_sample_1236 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=1.3101 ps=8.27 w=7.94 l=3.52
X1 B.t11 B.t9 B.t10 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=0 ps=0 w=7.94 l=3.52
X2 VDD1.t5 VP.t0 VTAIL.t5 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=3.0966 ps=16.66 w=7.94 l=3.52
X3 VTAIL.t7 VN.t1 VDD2.t4 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=1.3101 ps=8.27 w=7.94 l=3.52
X4 VDD2.t3 VN.t2 VTAIL.t8 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=1.3101 ps=8.27 w=7.94 l=3.52
X5 VDD1.t4 VP.t1 VTAIL.t1 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=1.3101 ps=8.27 w=7.94 l=3.52
X6 VTAIL.t0 VP.t2 VDD1.t3 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=1.3101 ps=8.27 w=7.94 l=3.52
X7 VDD2.t2 VN.t3 VTAIL.t9 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=3.0966 ps=16.66 w=7.94 l=3.52
X8 B.t8 B.t6 B.t7 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=0 ps=0 w=7.94 l=3.52
X9 B.t5 B.t3 B.t4 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=0 ps=0 w=7.94 l=3.52
X10 VDD2.t1 VN.t4 VTAIL.t6 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=3.0966 ps=16.66 w=7.94 l=3.52
X11 VDD1.t2 VP.t3 VTAIL.t4 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=3.0966 ps=16.66 w=7.94 l=3.52
X12 VTAIL.t2 VP.t4 VDD1.t1 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=1.3101 ps=8.27 w=7.94 l=3.52
X13 B.t2 B.t0 B.t1 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=0 ps=0 w=7.94 l=3.52
X14 VTAIL.t10 VN.t5 VDD2.t0 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=1.3101 pd=8.27 as=1.3101 ps=8.27 w=7.94 l=3.52
X15 VDD1.t0 VP.t5 VTAIL.t3 w_n4050_n2556# sky130_fd_pr__pfet_01v8 ad=3.0966 pd=16.66 as=1.3101 ps=8.27 w=7.94 l=3.52
R0 VN.n38 VN.n37 161.3
R1 VN.n36 VN.n21 161.3
R2 VN.n35 VN.n34 161.3
R3 VN.n33 VN.n22 161.3
R4 VN.n32 VN.n31 161.3
R5 VN.n30 VN.n23 161.3
R6 VN.n29 VN.n28 161.3
R7 VN.n27 VN.n24 161.3
R8 VN.n18 VN.n17 161.3
R9 VN.n16 VN.n1 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n2 161.3
R12 VN.n12 VN.n11 161.3
R13 VN.n10 VN.n3 161.3
R14 VN.n9 VN.n8 161.3
R15 VN.n7 VN.n4 161.3
R16 VN.n26 VN.t3 86.6956
R17 VN.n6 VN.t2 86.6956
R18 VN.n19 VN.n0 85.0223
R19 VN.n39 VN.n20 85.0223
R20 VN.n6 VN.n5 62.0355
R21 VN.n26 VN.n25 62.0355
R22 VN.n11 VN.n2 56.4773
R23 VN.n31 VN.n22 56.4773
R24 VN.n5 VN.t1 54.3624
R25 VN.n0 VN.t4 54.3624
R26 VN.n25 VN.t5 54.3624
R27 VN.n20 VN.t0 54.3624
R28 VN VN.n39 49.3881
R29 VN.n9 VN.n4 24.3439
R30 VN.n10 VN.n9 24.3439
R31 VN.n11 VN.n10 24.3439
R32 VN.n15 VN.n2 24.3439
R33 VN.n16 VN.n15 24.3439
R34 VN.n17 VN.n16 24.3439
R35 VN.n31 VN.n30 24.3439
R36 VN.n30 VN.n29 24.3439
R37 VN.n29 VN.n24 24.3439
R38 VN.n37 VN.n36 24.3439
R39 VN.n36 VN.n35 24.3439
R40 VN.n35 VN.n22 24.3439
R41 VN.n5 VN.n4 12.1722
R42 VN.n25 VN.n24 12.1722
R43 VN.n17 VN.n0 4.86919
R44 VN.n37 VN.n20 4.86919
R45 VN.n27 VN.n26 3.33651
R46 VN.n7 VN.n6 3.33651
R47 VN.n39 VN.n38 0.355081
R48 VN.n19 VN.n18 0.355081
R49 VN VN.n19 0.26685
R50 VN.n38 VN.n21 0.189894
R51 VN.n34 VN.n21 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n32 0.189894
R54 VN.n32 VN.n23 0.189894
R55 VN.n28 VN.n23 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n8 VN.n3 0.189894
R59 VN.n12 VN.n3 0.189894
R60 VN.n13 VN.n12 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n1 0.189894
R63 VN.n18 VN.n1 0.189894
R64 VTAIL.n170 VTAIL.n134 756.745
R65 VTAIL.n38 VTAIL.n2 756.745
R66 VTAIL.n128 VTAIL.n92 756.745
R67 VTAIL.n84 VTAIL.n48 756.745
R68 VTAIL.n146 VTAIL.n145 585
R69 VTAIL.n151 VTAIL.n150 585
R70 VTAIL.n153 VTAIL.n152 585
R71 VTAIL.n142 VTAIL.n141 585
R72 VTAIL.n159 VTAIL.n158 585
R73 VTAIL.n161 VTAIL.n160 585
R74 VTAIL.n138 VTAIL.n137 585
R75 VTAIL.n168 VTAIL.n167 585
R76 VTAIL.n169 VTAIL.n136 585
R77 VTAIL.n171 VTAIL.n170 585
R78 VTAIL.n14 VTAIL.n13 585
R79 VTAIL.n19 VTAIL.n18 585
R80 VTAIL.n21 VTAIL.n20 585
R81 VTAIL.n10 VTAIL.n9 585
R82 VTAIL.n27 VTAIL.n26 585
R83 VTAIL.n29 VTAIL.n28 585
R84 VTAIL.n6 VTAIL.n5 585
R85 VTAIL.n36 VTAIL.n35 585
R86 VTAIL.n37 VTAIL.n4 585
R87 VTAIL.n39 VTAIL.n38 585
R88 VTAIL.n129 VTAIL.n128 585
R89 VTAIL.n127 VTAIL.n94 585
R90 VTAIL.n126 VTAIL.n125 585
R91 VTAIL.n97 VTAIL.n95 585
R92 VTAIL.n120 VTAIL.n119 585
R93 VTAIL.n118 VTAIL.n117 585
R94 VTAIL.n101 VTAIL.n100 585
R95 VTAIL.n112 VTAIL.n111 585
R96 VTAIL.n110 VTAIL.n109 585
R97 VTAIL.n105 VTAIL.n104 585
R98 VTAIL.n85 VTAIL.n84 585
R99 VTAIL.n83 VTAIL.n50 585
R100 VTAIL.n82 VTAIL.n81 585
R101 VTAIL.n53 VTAIL.n51 585
R102 VTAIL.n76 VTAIL.n75 585
R103 VTAIL.n74 VTAIL.n73 585
R104 VTAIL.n57 VTAIL.n56 585
R105 VTAIL.n68 VTAIL.n67 585
R106 VTAIL.n66 VTAIL.n65 585
R107 VTAIL.n61 VTAIL.n60 585
R108 VTAIL.n147 VTAIL.t6 329.043
R109 VTAIL.n15 VTAIL.t4 329.043
R110 VTAIL.n106 VTAIL.t5 329.043
R111 VTAIL.n62 VTAIL.t9 329.043
R112 VTAIL.n151 VTAIL.n145 171.744
R113 VTAIL.n152 VTAIL.n151 171.744
R114 VTAIL.n152 VTAIL.n141 171.744
R115 VTAIL.n159 VTAIL.n141 171.744
R116 VTAIL.n160 VTAIL.n159 171.744
R117 VTAIL.n160 VTAIL.n137 171.744
R118 VTAIL.n168 VTAIL.n137 171.744
R119 VTAIL.n169 VTAIL.n168 171.744
R120 VTAIL.n170 VTAIL.n169 171.744
R121 VTAIL.n19 VTAIL.n13 171.744
R122 VTAIL.n20 VTAIL.n19 171.744
R123 VTAIL.n20 VTAIL.n9 171.744
R124 VTAIL.n27 VTAIL.n9 171.744
R125 VTAIL.n28 VTAIL.n27 171.744
R126 VTAIL.n28 VTAIL.n5 171.744
R127 VTAIL.n36 VTAIL.n5 171.744
R128 VTAIL.n37 VTAIL.n36 171.744
R129 VTAIL.n38 VTAIL.n37 171.744
R130 VTAIL.n128 VTAIL.n127 171.744
R131 VTAIL.n127 VTAIL.n126 171.744
R132 VTAIL.n126 VTAIL.n95 171.744
R133 VTAIL.n119 VTAIL.n95 171.744
R134 VTAIL.n119 VTAIL.n118 171.744
R135 VTAIL.n118 VTAIL.n100 171.744
R136 VTAIL.n111 VTAIL.n100 171.744
R137 VTAIL.n111 VTAIL.n110 171.744
R138 VTAIL.n110 VTAIL.n104 171.744
R139 VTAIL.n84 VTAIL.n83 171.744
R140 VTAIL.n83 VTAIL.n82 171.744
R141 VTAIL.n82 VTAIL.n51 171.744
R142 VTAIL.n75 VTAIL.n51 171.744
R143 VTAIL.n75 VTAIL.n74 171.744
R144 VTAIL.n74 VTAIL.n56 171.744
R145 VTAIL.n67 VTAIL.n56 171.744
R146 VTAIL.n67 VTAIL.n66 171.744
R147 VTAIL.n66 VTAIL.n60 171.744
R148 VTAIL.t6 VTAIL.n145 85.8723
R149 VTAIL.t4 VTAIL.n13 85.8723
R150 VTAIL.t5 VTAIL.n104 85.8723
R151 VTAIL.t9 VTAIL.n60 85.8723
R152 VTAIL.n91 VTAIL.n90 68.3956
R153 VTAIL.n47 VTAIL.n46 68.3956
R154 VTAIL.n1 VTAIL.n0 68.3954
R155 VTAIL.n45 VTAIL.n44 68.3954
R156 VTAIL.n175 VTAIL.n174 34.9005
R157 VTAIL.n43 VTAIL.n42 34.9005
R158 VTAIL.n133 VTAIL.n132 34.9005
R159 VTAIL.n89 VTAIL.n88 34.9005
R160 VTAIL.n47 VTAIL.n45 25.8496
R161 VTAIL.n175 VTAIL.n133 22.5307
R162 VTAIL.n171 VTAIL.n136 13.1884
R163 VTAIL.n39 VTAIL.n4 13.1884
R164 VTAIL.n129 VTAIL.n94 13.1884
R165 VTAIL.n85 VTAIL.n50 13.1884
R166 VTAIL.n167 VTAIL.n166 12.8005
R167 VTAIL.n172 VTAIL.n134 12.8005
R168 VTAIL.n35 VTAIL.n34 12.8005
R169 VTAIL.n40 VTAIL.n2 12.8005
R170 VTAIL.n130 VTAIL.n92 12.8005
R171 VTAIL.n125 VTAIL.n96 12.8005
R172 VTAIL.n86 VTAIL.n48 12.8005
R173 VTAIL.n81 VTAIL.n52 12.8005
R174 VTAIL.n165 VTAIL.n138 12.0247
R175 VTAIL.n33 VTAIL.n6 12.0247
R176 VTAIL.n124 VTAIL.n97 12.0247
R177 VTAIL.n80 VTAIL.n53 12.0247
R178 VTAIL.n162 VTAIL.n161 11.249
R179 VTAIL.n30 VTAIL.n29 11.249
R180 VTAIL.n121 VTAIL.n120 11.249
R181 VTAIL.n77 VTAIL.n76 11.249
R182 VTAIL.n147 VTAIL.n146 10.7238
R183 VTAIL.n15 VTAIL.n14 10.7238
R184 VTAIL.n106 VTAIL.n105 10.7238
R185 VTAIL.n62 VTAIL.n61 10.7238
R186 VTAIL.n158 VTAIL.n140 10.4732
R187 VTAIL.n26 VTAIL.n8 10.4732
R188 VTAIL.n117 VTAIL.n99 10.4732
R189 VTAIL.n73 VTAIL.n55 10.4732
R190 VTAIL.n157 VTAIL.n142 9.69747
R191 VTAIL.n25 VTAIL.n10 9.69747
R192 VTAIL.n116 VTAIL.n101 9.69747
R193 VTAIL.n72 VTAIL.n57 9.69747
R194 VTAIL.n174 VTAIL.n173 9.45567
R195 VTAIL.n42 VTAIL.n41 9.45567
R196 VTAIL.n132 VTAIL.n131 9.45567
R197 VTAIL.n88 VTAIL.n87 9.45567
R198 VTAIL.n173 VTAIL.n172 9.3005
R199 VTAIL.n149 VTAIL.n148 9.3005
R200 VTAIL.n144 VTAIL.n143 9.3005
R201 VTAIL.n155 VTAIL.n154 9.3005
R202 VTAIL.n157 VTAIL.n156 9.3005
R203 VTAIL.n140 VTAIL.n139 9.3005
R204 VTAIL.n163 VTAIL.n162 9.3005
R205 VTAIL.n165 VTAIL.n164 9.3005
R206 VTAIL.n166 VTAIL.n135 9.3005
R207 VTAIL.n41 VTAIL.n40 9.3005
R208 VTAIL.n17 VTAIL.n16 9.3005
R209 VTAIL.n12 VTAIL.n11 9.3005
R210 VTAIL.n23 VTAIL.n22 9.3005
R211 VTAIL.n25 VTAIL.n24 9.3005
R212 VTAIL.n8 VTAIL.n7 9.3005
R213 VTAIL.n31 VTAIL.n30 9.3005
R214 VTAIL.n33 VTAIL.n32 9.3005
R215 VTAIL.n34 VTAIL.n3 9.3005
R216 VTAIL.n108 VTAIL.n107 9.3005
R217 VTAIL.n103 VTAIL.n102 9.3005
R218 VTAIL.n114 VTAIL.n113 9.3005
R219 VTAIL.n116 VTAIL.n115 9.3005
R220 VTAIL.n99 VTAIL.n98 9.3005
R221 VTAIL.n122 VTAIL.n121 9.3005
R222 VTAIL.n124 VTAIL.n123 9.3005
R223 VTAIL.n96 VTAIL.n93 9.3005
R224 VTAIL.n131 VTAIL.n130 9.3005
R225 VTAIL.n64 VTAIL.n63 9.3005
R226 VTAIL.n59 VTAIL.n58 9.3005
R227 VTAIL.n70 VTAIL.n69 9.3005
R228 VTAIL.n72 VTAIL.n71 9.3005
R229 VTAIL.n55 VTAIL.n54 9.3005
R230 VTAIL.n78 VTAIL.n77 9.3005
R231 VTAIL.n80 VTAIL.n79 9.3005
R232 VTAIL.n52 VTAIL.n49 9.3005
R233 VTAIL.n87 VTAIL.n86 9.3005
R234 VTAIL.n154 VTAIL.n153 8.92171
R235 VTAIL.n22 VTAIL.n21 8.92171
R236 VTAIL.n113 VTAIL.n112 8.92171
R237 VTAIL.n69 VTAIL.n68 8.92171
R238 VTAIL.n150 VTAIL.n144 8.14595
R239 VTAIL.n18 VTAIL.n12 8.14595
R240 VTAIL.n109 VTAIL.n103 8.14595
R241 VTAIL.n65 VTAIL.n59 8.14595
R242 VTAIL.n149 VTAIL.n146 7.3702
R243 VTAIL.n17 VTAIL.n14 7.3702
R244 VTAIL.n108 VTAIL.n105 7.3702
R245 VTAIL.n64 VTAIL.n61 7.3702
R246 VTAIL.n150 VTAIL.n149 5.81868
R247 VTAIL.n18 VTAIL.n17 5.81868
R248 VTAIL.n109 VTAIL.n108 5.81868
R249 VTAIL.n65 VTAIL.n64 5.81868
R250 VTAIL.n153 VTAIL.n144 5.04292
R251 VTAIL.n21 VTAIL.n12 5.04292
R252 VTAIL.n112 VTAIL.n103 5.04292
R253 VTAIL.n68 VTAIL.n59 5.04292
R254 VTAIL.n154 VTAIL.n142 4.26717
R255 VTAIL.n22 VTAIL.n10 4.26717
R256 VTAIL.n113 VTAIL.n101 4.26717
R257 VTAIL.n69 VTAIL.n57 4.26717
R258 VTAIL.n0 VTAIL.t8 4.09433
R259 VTAIL.n0 VTAIL.t7 4.09433
R260 VTAIL.n44 VTAIL.t1 4.09433
R261 VTAIL.n44 VTAIL.t2 4.09433
R262 VTAIL.n90 VTAIL.t3 4.09433
R263 VTAIL.n90 VTAIL.t0 4.09433
R264 VTAIL.n46 VTAIL.t11 4.09433
R265 VTAIL.n46 VTAIL.t10 4.09433
R266 VTAIL.n158 VTAIL.n157 3.49141
R267 VTAIL.n26 VTAIL.n25 3.49141
R268 VTAIL.n117 VTAIL.n116 3.49141
R269 VTAIL.n73 VTAIL.n72 3.49141
R270 VTAIL.n89 VTAIL.n47 3.31947
R271 VTAIL.n133 VTAIL.n91 3.31947
R272 VTAIL.n45 VTAIL.n43 3.31947
R273 VTAIL.n161 VTAIL.n140 2.71565
R274 VTAIL.n29 VTAIL.n8 2.71565
R275 VTAIL.n120 VTAIL.n99 2.71565
R276 VTAIL.n76 VTAIL.n55 2.71565
R277 VTAIL VTAIL.n175 2.43153
R278 VTAIL.n148 VTAIL.n147 2.4129
R279 VTAIL.n16 VTAIL.n15 2.4129
R280 VTAIL.n107 VTAIL.n106 2.4129
R281 VTAIL.n63 VTAIL.n62 2.4129
R282 VTAIL.n91 VTAIL.n89 2.12981
R283 VTAIL.n43 VTAIL.n1 2.12981
R284 VTAIL.n162 VTAIL.n138 1.93989
R285 VTAIL.n30 VTAIL.n6 1.93989
R286 VTAIL.n121 VTAIL.n97 1.93989
R287 VTAIL.n77 VTAIL.n53 1.93989
R288 VTAIL.n167 VTAIL.n165 1.16414
R289 VTAIL.n174 VTAIL.n134 1.16414
R290 VTAIL.n35 VTAIL.n33 1.16414
R291 VTAIL.n42 VTAIL.n2 1.16414
R292 VTAIL.n132 VTAIL.n92 1.16414
R293 VTAIL.n125 VTAIL.n124 1.16414
R294 VTAIL.n88 VTAIL.n48 1.16414
R295 VTAIL.n81 VTAIL.n80 1.16414
R296 VTAIL VTAIL.n1 0.888431
R297 VTAIL.n166 VTAIL.n136 0.388379
R298 VTAIL.n172 VTAIL.n171 0.388379
R299 VTAIL.n34 VTAIL.n4 0.388379
R300 VTAIL.n40 VTAIL.n39 0.388379
R301 VTAIL.n130 VTAIL.n129 0.388379
R302 VTAIL.n96 VTAIL.n94 0.388379
R303 VTAIL.n86 VTAIL.n85 0.388379
R304 VTAIL.n52 VTAIL.n50 0.388379
R305 VTAIL.n148 VTAIL.n143 0.155672
R306 VTAIL.n155 VTAIL.n143 0.155672
R307 VTAIL.n156 VTAIL.n155 0.155672
R308 VTAIL.n156 VTAIL.n139 0.155672
R309 VTAIL.n163 VTAIL.n139 0.155672
R310 VTAIL.n164 VTAIL.n163 0.155672
R311 VTAIL.n164 VTAIL.n135 0.155672
R312 VTAIL.n173 VTAIL.n135 0.155672
R313 VTAIL.n16 VTAIL.n11 0.155672
R314 VTAIL.n23 VTAIL.n11 0.155672
R315 VTAIL.n24 VTAIL.n23 0.155672
R316 VTAIL.n24 VTAIL.n7 0.155672
R317 VTAIL.n31 VTAIL.n7 0.155672
R318 VTAIL.n32 VTAIL.n31 0.155672
R319 VTAIL.n32 VTAIL.n3 0.155672
R320 VTAIL.n41 VTAIL.n3 0.155672
R321 VTAIL.n131 VTAIL.n93 0.155672
R322 VTAIL.n123 VTAIL.n93 0.155672
R323 VTAIL.n123 VTAIL.n122 0.155672
R324 VTAIL.n122 VTAIL.n98 0.155672
R325 VTAIL.n115 VTAIL.n98 0.155672
R326 VTAIL.n115 VTAIL.n114 0.155672
R327 VTAIL.n114 VTAIL.n102 0.155672
R328 VTAIL.n107 VTAIL.n102 0.155672
R329 VTAIL.n87 VTAIL.n49 0.155672
R330 VTAIL.n79 VTAIL.n49 0.155672
R331 VTAIL.n79 VTAIL.n78 0.155672
R332 VTAIL.n78 VTAIL.n54 0.155672
R333 VTAIL.n71 VTAIL.n54 0.155672
R334 VTAIL.n71 VTAIL.n70 0.155672
R335 VTAIL.n70 VTAIL.n58 0.155672
R336 VTAIL.n63 VTAIL.n58 0.155672
R337 VDD2.n79 VDD2.n43 756.745
R338 VDD2.n36 VDD2.n0 756.745
R339 VDD2.n80 VDD2.n79 585
R340 VDD2.n78 VDD2.n45 585
R341 VDD2.n77 VDD2.n76 585
R342 VDD2.n48 VDD2.n46 585
R343 VDD2.n71 VDD2.n70 585
R344 VDD2.n69 VDD2.n68 585
R345 VDD2.n52 VDD2.n51 585
R346 VDD2.n63 VDD2.n62 585
R347 VDD2.n61 VDD2.n60 585
R348 VDD2.n56 VDD2.n55 585
R349 VDD2.n12 VDD2.n11 585
R350 VDD2.n17 VDD2.n16 585
R351 VDD2.n19 VDD2.n18 585
R352 VDD2.n8 VDD2.n7 585
R353 VDD2.n25 VDD2.n24 585
R354 VDD2.n27 VDD2.n26 585
R355 VDD2.n4 VDD2.n3 585
R356 VDD2.n34 VDD2.n33 585
R357 VDD2.n35 VDD2.n2 585
R358 VDD2.n37 VDD2.n36 585
R359 VDD2.n57 VDD2.t5 329.043
R360 VDD2.n13 VDD2.t3 329.043
R361 VDD2.n79 VDD2.n78 171.744
R362 VDD2.n78 VDD2.n77 171.744
R363 VDD2.n77 VDD2.n46 171.744
R364 VDD2.n70 VDD2.n46 171.744
R365 VDD2.n70 VDD2.n69 171.744
R366 VDD2.n69 VDD2.n51 171.744
R367 VDD2.n62 VDD2.n51 171.744
R368 VDD2.n62 VDD2.n61 171.744
R369 VDD2.n61 VDD2.n55 171.744
R370 VDD2.n17 VDD2.n11 171.744
R371 VDD2.n18 VDD2.n17 171.744
R372 VDD2.n18 VDD2.n7 171.744
R373 VDD2.n25 VDD2.n7 171.744
R374 VDD2.n26 VDD2.n25 171.744
R375 VDD2.n26 VDD2.n3 171.744
R376 VDD2.n34 VDD2.n3 171.744
R377 VDD2.n35 VDD2.n34 171.744
R378 VDD2.n36 VDD2.n35 171.744
R379 VDD2.t5 VDD2.n55 85.8723
R380 VDD2.t3 VDD2.n11 85.8723
R381 VDD2.n42 VDD2.n41 85.8486
R382 VDD2 VDD2.n85 85.8458
R383 VDD2.n42 VDD2.n40 54.0132
R384 VDD2.n84 VDD2.n83 51.5793
R385 VDD2.n84 VDD2.n42 41.3468
R386 VDD2.n80 VDD2.n45 13.1884
R387 VDD2.n37 VDD2.n2 13.1884
R388 VDD2.n81 VDD2.n43 12.8005
R389 VDD2.n76 VDD2.n47 12.8005
R390 VDD2.n33 VDD2.n32 12.8005
R391 VDD2.n38 VDD2.n0 12.8005
R392 VDD2.n75 VDD2.n48 12.0247
R393 VDD2.n31 VDD2.n4 12.0247
R394 VDD2.n72 VDD2.n71 11.249
R395 VDD2.n28 VDD2.n27 11.249
R396 VDD2.n57 VDD2.n56 10.7238
R397 VDD2.n13 VDD2.n12 10.7238
R398 VDD2.n68 VDD2.n50 10.4732
R399 VDD2.n24 VDD2.n6 10.4732
R400 VDD2.n67 VDD2.n52 9.69747
R401 VDD2.n23 VDD2.n8 9.69747
R402 VDD2.n83 VDD2.n82 9.45567
R403 VDD2.n40 VDD2.n39 9.45567
R404 VDD2.n59 VDD2.n58 9.3005
R405 VDD2.n54 VDD2.n53 9.3005
R406 VDD2.n65 VDD2.n64 9.3005
R407 VDD2.n67 VDD2.n66 9.3005
R408 VDD2.n50 VDD2.n49 9.3005
R409 VDD2.n73 VDD2.n72 9.3005
R410 VDD2.n75 VDD2.n74 9.3005
R411 VDD2.n47 VDD2.n44 9.3005
R412 VDD2.n82 VDD2.n81 9.3005
R413 VDD2.n39 VDD2.n38 9.3005
R414 VDD2.n15 VDD2.n14 9.3005
R415 VDD2.n10 VDD2.n9 9.3005
R416 VDD2.n21 VDD2.n20 9.3005
R417 VDD2.n23 VDD2.n22 9.3005
R418 VDD2.n6 VDD2.n5 9.3005
R419 VDD2.n29 VDD2.n28 9.3005
R420 VDD2.n31 VDD2.n30 9.3005
R421 VDD2.n32 VDD2.n1 9.3005
R422 VDD2.n64 VDD2.n63 8.92171
R423 VDD2.n20 VDD2.n19 8.92171
R424 VDD2.n60 VDD2.n54 8.14595
R425 VDD2.n16 VDD2.n10 8.14595
R426 VDD2.n59 VDD2.n56 7.3702
R427 VDD2.n15 VDD2.n12 7.3702
R428 VDD2.n60 VDD2.n59 5.81868
R429 VDD2.n16 VDD2.n15 5.81868
R430 VDD2.n63 VDD2.n54 5.04292
R431 VDD2.n19 VDD2.n10 5.04292
R432 VDD2.n64 VDD2.n52 4.26717
R433 VDD2.n20 VDD2.n8 4.26717
R434 VDD2.n85 VDD2.t0 4.09433
R435 VDD2.n85 VDD2.t2 4.09433
R436 VDD2.n41 VDD2.t4 4.09433
R437 VDD2.n41 VDD2.t1 4.09433
R438 VDD2.n68 VDD2.n67 3.49141
R439 VDD2.n24 VDD2.n23 3.49141
R440 VDD2.n71 VDD2.n50 2.71565
R441 VDD2.n27 VDD2.n6 2.71565
R442 VDD2 VDD2.n84 2.54791
R443 VDD2.n58 VDD2.n57 2.4129
R444 VDD2.n14 VDD2.n13 2.4129
R445 VDD2.n72 VDD2.n48 1.93989
R446 VDD2.n28 VDD2.n4 1.93989
R447 VDD2.n83 VDD2.n43 1.16414
R448 VDD2.n76 VDD2.n75 1.16414
R449 VDD2.n33 VDD2.n31 1.16414
R450 VDD2.n40 VDD2.n0 1.16414
R451 VDD2.n81 VDD2.n80 0.388379
R452 VDD2.n47 VDD2.n45 0.388379
R453 VDD2.n32 VDD2.n2 0.388379
R454 VDD2.n38 VDD2.n37 0.388379
R455 VDD2.n82 VDD2.n44 0.155672
R456 VDD2.n74 VDD2.n44 0.155672
R457 VDD2.n74 VDD2.n73 0.155672
R458 VDD2.n73 VDD2.n49 0.155672
R459 VDD2.n66 VDD2.n49 0.155672
R460 VDD2.n66 VDD2.n65 0.155672
R461 VDD2.n65 VDD2.n53 0.155672
R462 VDD2.n58 VDD2.n53 0.155672
R463 VDD2.n14 VDD2.n9 0.155672
R464 VDD2.n21 VDD2.n9 0.155672
R465 VDD2.n22 VDD2.n21 0.155672
R466 VDD2.n22 VDD2.n5 0.155672
R467 VDD2.n29 VDD2.n5 0.155672
R468 VDD2.n30 VDD2.n29 0.155672
R469 VDD2.n30 VDD2.n1 0.155672
R470 VDD2.n39 VDD2.n1 0.155672
R471 B.n369 B.n368 585
R472 B.n367 B.n122 585
R473 B.n366 B.n365 585
R474 B.n364 B.n123 585
R475 B.n363 B.n362 585
R476 B.n361 B.n124 585
R477 B.n360 B.n359 585
R478 B.n358 B.n125 585
R479 B.n357 B.n356 585
R480 B.n355 B.n126 585
R481 B.n354 B.n353 585
R482 B.n352 B.n127 585
R483 B.n351 B.n350 585
R484 B.n349 B.n128 585
R485 B.n348 B.n347 585
R486 B.n346 B.n129 585
R487 B.n345 B.n344 585
R488 B.n343 B.n130 585
R489 B.n342 B.n341 585
R490 B.n340 B.n131 585
R491 B.n339 B.n338 585
R492 B.n337 B.n132 585
R493 B.n336 B.n335 585
R494 B.n334 B.n133 585
R495 B.n333 B.n332 585
R496 B.n331 B.n134 585
R497 B.n330 B.n329 585
R498 B.n328 B.n135 585
R499 B.n327 B.n326 585
R500 B.n325 B.n136 585
R501 B.n324 B.n323 585
R502 B.n319 B.n137 585
R503 B.n318 B.n317 585
R504 B.n316 B.n138 585
R505 B.n315 B.n314 585
R506 B.n313 B.n139 585
R507 B.n312 B.n311 585
R508 B.n310 B.n140 585
R509 B.n309 B.n308 585
R510 B.n306 B.n141 585
R511 B.n305 B.n304 585
R512 B.n303 B.n144 585
R513 B.n302 B.n301 585
R514 B.n300 B.n145 585
R515 B.n299 B.n298 585
R516 B.n297 B.n146 585
R517 B.n296 B.n295 585
R518 B.n294 B.n147 585
R519 B.n293 B.n292 585
R520 B.n291 B.n148 585
R521 B.n290 B.n289 585
R522 B.n288 B.n149 585
R523 B.n287 B.n286 585
R524 B.n285 B.n150 585
R525 B.n284 B.n283 585
R526 B.n282 B.n151 585
R527 B.n281 B.n280 585
R528 B.n279 B.n152 585
R529 B.n278 B.n277 585
R530 B.n276 B.n153 585
R531 B.n275 B.n274 585
R532 B.n273 B.n154 585
R533 B.n272 B.n271 585
R534 B.n270 B.n155 585
R535 B.n269 B.n268 585
R536 B.n267 B.n156 585
R537 B.n266 B.n265 585
R538 B.n264 B.n157 585
R539 B.n263 B.n262 585
R540 B.n370 B.n121 585
R541 B.n372 B.n371 585
R542 B.n373 B.n120 585
R543 B.n375 B.n374 585
R544 B.n376 B.n119 585
R545 B.n378 B.n377 585
R546 B.n379 B.n118 585
R547 B.n381 B.n380 585
R548 B.n382 B.n117 585
R549 B.n384 B.n383 585
R550 B.n385 B.n116 585
R551 B.n387 B.n386 585
R552 B.n388 B.n115 585
R553 B.n390 B.n389 585
R554 B.n391 B.n114 585
R555 B.n393 B.n392 585
R556 B.n394 B.n113 585
R557 B.n396 B.n395 585
R558 B.n397 B.n112 585
R559 B.n399 B.n398 585
R560 B.n400 B.n111 585
R561 B.n402 B.n401 585
R562 B.n403 B.n110 585
R563 B.n405 B.n404 585
R564 B.n406 B.n109 585
R565 B.n408 B.n407 585
R566 B.n409 B.n108 585
R567 B.n411 B.n410 585
R568 B.n412 B.n107 585
R569 B.n414 B.n413 585
R570 B.n415 B.n106 585
R571 B.n417 B.n416 585
R572 B.n418 B.n105 585
R573 B.n420 B.n419 585
R574 B.n421 B.n104 585
R575 B.n423 B.n422 585
R576 B.n424 B.n103 585
R577 B.n426 B.n425 585
R578 B.n427 B.n102 585
R579 B.n429 B.n428 585
R580 B.n430 B.n101 585
R581 B.n432 B.n431 585
R582 B.n433 B.n100 585
R583 B.n435 B.n434 585
R584 B.n436 B.n99 585
R585 B.n438 B.n437 585
R586 B.n439 B.n98 585
R587 B.n441 B.n440 585
R588 B.n442 B.n97 585
R589 B.n444 B.n443 585
R590 B.n445 B.n96 585
R591 B.n447 B.n446 585
R592 B.n448 B.n95 585
R593 B.n450 B.n449 585
R594 B.n451 B.n94 585
R595 B.n453 B.n452 585
R596 B.n454 B.n93 585
R597 B.n456 B.n455 585
R598 B.n457 B.n92 585
R599 B.n459 B.n458 585
R600 B.n460 B.n91 585
R601 B.n462 B.n461 585
R602 B.n463 B.n90 585
R603 B.n465 B.n464 585
R604 B.n466 B.n89 585
R605 B.n468 B.n467 585
R606 B.n469 B.n88 585
R607 B.n471 B.n470 585
R608 B.n472 B.n87 585
R609 B.n474 B.n473 585
R610 B.n475 B.n86 585
R611 B.n477 B.n476 585
R612 B.n478 B.n85 585
R613 B.n480 B.n479 585
R614 B.n481 B.n84 585
R615 B.n483 B.n482 585
R616 B.n484 B.n83 585
R617 B.n486 B.n485 585
R618 B.n487 B.n82 585
R619 B.n489 B.n488 585
R620 B.n490 B.n81 585
R621 B.n492 B.n491 585
R622 B.n493 B.n80 585
R623 B.n495 B.n494 585
R624 B.n496 B.n79 585
R625 B.n498 B.n497 585
R626 B.n499 B.n78 585
R627 B.n501 B.n500 585
R628 B.n502 B.n77 585
R629 B.n504 B.n503 585
R630 B.n505 B.n76 585
R631 B.n507 B.n506 585
R632 B.n508 B.n75 585
R633 B.n510 B.n509 585
R634 B.n511 B.n74 585
R635 B.n513 B.n512 585
R636 B.n514 B.n73 585
R637 B.n516 B.n515 585
R638 B.n517 B.n72 585
R639 B.n519 B.n518 585
R640 B.n520 B.n71 585
R641 B.n522 B.n521 585
R642 B.n523 B.n70 585
R643 B.n525 B.n524 585
R644 B.n526 B.n69 585
R645 B.n528 B.n527 585
R646 B.n529 B.n68 585
R647 B.n531 B.n530 585
R648 B.n636 B.n635 585
R649 B.n634 B.n29 585
R650 B.n633 B.n632 585
R651 B.n631 B.n30 585
R652 B.n630 B.n629 585
R653 B.n628 B.n31 585
R654 B.n627 B.n626 585
R655 B.n625 B.n32 585
R656 B.n624 B.n623 585
R657 B.n622 B.n33 585
R658 B.n621 B.n620 585
R659 B.n619 B.n34 585
R660 B.n618 B.n617 585
R661 B.n616 B.n35 585
R662 B.n615 B.n614 585
R663 B.n613 B.n36 585
R664 B.n612 B.n611 585
R665 B.n610 B.n37 585
R666 B.n609 B.n608 585
R667 B.n607 B.n38 585
R668 B.n606 B.n605 585
R669 B.n604 B.n39 585
R670 B.n603 B.n602 585
R671 B.n601 B.n40 585
R672 B.n600 B.n599 585
R673 B.n598 B.n41 585
R674 B.n597 B.n596 585
R675 B.n595 B.n42 585
R676 B.n594 B.n593 585
R677 B.n592 B.n43 585
R678 B.n590 B.n589 585
R679 B.n588 B.n46 585
R680 B.n587 B.n586 585
R681 B.n585 B.n47 585
R682 B.n584 B.n583 585
R683 B.n582 B.n48 585
R684 B.n581 B.n580 585
R685 B.n579 B.n49 585
R686 B.n578 B.n577 585
R687 B.n576 B.n575 585
R688 B.n574 B.n53 585
R689 B.n573 B.n572 585
R690 B.n571 B.n54 585
R691 B.n570 B.n569 585
R692 B.n568 B.n55 585
R693 B.n567 B.n566 585
R694 B.n565 B.n56 585
R695 B.n564 B.n563 585
R696 B.n562 B.n57 585
R697 B.n561 B.n560 585
R698 B.n559 B.n58 585
R699 B.n558 B.n557 585
R700 B.n556 B.n59 585
R701 B.n555 B.n554 585
R702 B.n553 B.n60 585
R703 B.n552 B.n551 585
R704 B.n550 B.n61 585
R705 B.n549 B.n548 585
R706 B.n547 B.n62 585
R707 B.n546 B.n545 585
R708 B.n544 B.n63 585
R709 B.n543 B.n542 585
R710 B.n541 B.n64 585
R711 B.n540 B.n539 585
R712 B.n538 B.n65 585
R713 B.n537 B.n536 585
R714 B.n535 B.n66 585
R715 B.n534 B.n533 585
R716 B.n532 B.n67 585
R717 B.n637 B.n28 585
R718 B.n639 B.n638 585
R719 B.n640 B.n27 585
R720 B.n642 B.n641 585
R721 B.n643 B.n26 585
R722 B.n645 B.n644 585
R723 B.n646 B.n25 585
R724 B.n648 B.n647 585
R725 B.n649 B.n24 585
R726 B.n651 B.n650 585
R727 B.n652 B.n23 585
R728 B.n654 B.n653 585
R729 B.n655 B.n22 585
R730 B.n657 B.n656 585
R731 B.n658 B.n21 585
R732 B.n660 B.n659 585
R733 B.n661 B.n20 585
R734 B.n663 B.n662 585
R735 B.n664 B.n19 585
R736 B.n666 B.n665 585
R737 B.n667 B.n18 585
R738 B.n669 B.n668 585
R739 B.n670 B.n17 585
R740 B.n672 B.n671 585
R741 B.n673 B.n16 585
R742 B.n675 B.n674 585
R743 B.n676 B.n15 585
R744 B.n678 B.n677 585
R745 B.n679 B.n14 585
R746 B.n681 B.n680 585
R747 B.n682 B.n13 585
R748 B.n684 B.n683 585
R749 B.n685 B.n12 585
R750 B.n687 B.n686 585
R751 B.n688 B.n11 585
R752 B.n690 B.n689 585
R753 B.n691 B.n10 585
R754 B.n693 B.n692 585
R755 B.n694 B.n9 585
R756 B.n696 B.n695 585
R757 B.n697 B.n8 585
R758 B.n699 B.n698 585
R759 B.n700 B.n7 585
R760 B.n702 B.n701 585
R761 B.n703 B.n6 585
R762 B.n705 B.n704 585
R763 B.n706 B.n5 585
R764 B.n708 B.n707 585
R765 B.n709 B.n4 585
R766 B.n711 B.n710 585
R767 B.n712 B.n3 585
R768 B.n714 B.n713 585
R769 B.n715 B.n0 585
R770 B.n2 B.n1 585
R771 B.n185 B.n184 585
R772 B.n186 B.n183 585
R773 B.n188 B.n187 585
R774 B.n189 B.n182 585
R775 B.n191 B.n190 585
R776 B.n192 B.n181 585
R777 B.n194 B.n193 585
R778 B.n195 B.n180 585
R779 B.n197 B.n196 585
R780 B.n198 B.n179 585
R781 B.n200 B.n199 585
R782 B.n201 B.n178 585
R783 B.n203 B.n202 585
R784 B.n204 B.n177 585
R785 B.n206 B.n205 585
R786 B.n207 B.n176 585
R787 B.n209 B.n208 585
R788 B.n210 B.n175 585
R789 B.n212 B.n211 585
R790 B.n213 B.n174 585
R791 B.n215 B.n214 585
R792 B.n216 B.n173 585
R793 B.n218 B.n217 585
R794 B.n219 B.n172 585
R795 B.n221 B.n220 585
R796 B.n222 B.n171 585
R797 B.n224 B.n223 585
R798 B.n225 B.n170 585
R799 B.n227 B.n226 585
R800 B.n228 B.n169 585
R801 B.n230 B.n229 585
R802 B.n231 B.n168 585
R803 B.n233 B.n232 585
R804 B.n234 B.n167 585
R805 B.n236 B.n235 585
R806 B.n237 B.n166 585
R807 B.n239 B.n238 585
R808 B.n240 B.n165 585
R809 B.n242 B.n241 585
R810 B.n243 B.n164 585
R811 B.n245 B.n244 585
R812 B.n246 B.n163 585
R813 B.n248 B.n247 585
R814 B.n249 B.n162 585
R815 B.n251 B.n250 585
R816 B.n252 B.n161 585
R817 B.n254 B.n253 585
R818 B.n255 B.n160 585
R819 B.n257 B.n256 585
R820 B.n258 B.n159 585
R821 B.n260 B.n259 585
R822 B.n261 B.n158 585
R823 B.n262 B.n261 478.086
R824 B.n368 B.n121 478.086
R825 B.n530 B.n67 478.086
R826 B.n637 B.n636 478.086
R827 B.n320 B.t7 377.387
R828 B.n50 B.t11 377.387
R829 B.n142 B.t1 377.387
R830 B.n44 B.t5 377.387
R831 B.n321 B.t8 302.721
R832 B.n51 B.t10 302.721
R833 B.n143 B.t2 302.721
R834 B.n45 B.t4 302.721
R835 B.n320 B.t6 264.147
R836 B.n50 B.t9 264.147
R837 B.n142 B.t0 263.887
R838 B.n44 B.t3 263.887
R839 B.n717 B.n716 256.663
R840 B.n716 B.n715 235.042
R841 B.n716 B.n2 235.042
R842 B.n262 B.n157 163.367
R843 B.n266 B.n157 163.367
R844 B.n267 B.n266 163.367
R845 B.n268 B.n267 163.367
R846 B.n268 B.n155 163.367
R847 B.n272 B.n155 163.367
R848 B.n273 B.n272 163.367
R849 B.n274 B.n273 163.367
R850 B.n274 B.n153 163.367
R851 B.n278 B.n153 163.367
R852 B.n279 B.n278 163.367
R853 B.n280 B.n279 163.367
R854 B.n280 B.n151 163.367
R855 B.n284 B.n151 163.367
R856 B.n285 B.n284 163.367
R857 B.n286 B.n285 163.367
R858 B.n286 B.n149 163.367
R859 B.n290 B.n149 163.367
R860 B.n291 B.n290 163.367
R861 B.n292 B.n291 163.367
R862 B.n292 B.n147 163.367
R863 B.n296 B.n147 163.367
R864 B.n297 B.n296 163.367
R865 B.n298 B.n297 163.367
R866 B.n298 B.n145 163.367
R867 B.n302 B.n145 163.367
R868 B.n303 B.n302 163.367
R869 B.n304 B.n303 163.367
R870 B.n304 B.n141 163.367
R871 B.n309 B.n141 163.367
R872 B.n310 B.n309 163.367
R873 B.n311 B.n310 163.367
R874 B.n311 B.n139 163.367
R875 B.n315 B.n139 163.367
R876 B.n316 B.n315 163.367
R877 B.n317 B.n316 163.367
R878 B.n317 B.n137 163.367
R879 B.n324 B.n137 163.367
R880 B.n325 B.n324 163.367
R881 B.n326 B.n325 163.367
R882 B.n326 B.n135 163.367
R883 B.n330 B.n135 163.367
R884 B.n331 B.n330 163.367
R885 B.n332 B.n331 163.367
R886 B.n332 B.n133 163.367
R887 B.n336 B.n133 163.367
R888 B.n337 B.n336 163.367
R889 B.n338 B.n337 163.367
R890 B.n338 B.n131 163.367
R891 B.n342 B.n131 163.367
R892 B.n343 B.n342 163.367
R893 B.n344 B.n343 163.367
R894 B.n344 B.n129 163.367
R895 B.n348 B.n129 163.367
R896 B.n349 B.n348 163.367
R897 B.n350 B.n349 163.367
R898 B.n350 B.n127 163.367
R899 B.n354 B.n127 163.367
R900 B.n355 B.n354 163.367
R901 B.n356 B.n355 163.367
R902 B.n356 B.n125 163.367
R903 B.n360 B.n125 163.367
R904 B.n361 B.n360 163.367
R905 B.n362 B.n361 163.367
R906 B.n362 B.n123 163.367
R907 B.n366 B.n123 163.367
R908 B.n367 B.n366 163.367
R909 B.n368 B.n367 163.367
R910 B.n530 B.n529 163.367
R911 B.n529 B.n528 163.367
R912 B.n528 B.n69 163.367
R913 B.n524 B.n69 163.367
R914 B.n524 B.n523 163.367
R915 B.n523 B.n522 163.367
R916 B.n522 B.n71 163.367
R917 B.n518 B.n71 163.367
R918 B.n518 B.n517 163.367
R919 B.n517 B.n516 163.367
R920 B.n516 B.n73 163.367
R921 B.n512 B.n73 163.367
R922 B.n512 B.n511 163.367
R923 B.n511 B.n510 163.367
R924 B.n510 B.n75 163.367
R925 B.n506 B.n75 163.367
R926 B.n506 B.n505 163.367
R927 B.n505 B.n504 163.367
R928 B.n504 B.n77 163.367
R929 B.n500 B.n77 163.367
R930 B.n500 B.n499 163.367
R931 B.n499 B.n498 163.367
R932 B.n498 B.n79 163.367
R933 B.n494 B.n79 163.367
R934 B.n494 B.n493 163.367
R935 B.n493 B.n492 163.367
R936 B.n492 B.n81 163.367
R937 B.n488 B.n81 163.367
R938 B.n488 B.n487 163.367
R939 B.n487 B.n486 163.367
R940 B.n486 B.n83 163.367
R941 B.n482 B.n83 163.367
R942 B.n482 B.n481 163.367
R943 B.n481 B.n480 163.367
R944 B.n480 B.n85 163.367
R945 B.n476 B.n85 163.367
R946 B.n476 B.n475 163.367
R947 B.n475 B.n474 163.367
R948 B.n474 B.n87 163.367
R949 B.n470 B.n87 163.367
R950 B.n470 B.n469 163.367
R951 B.n469 B.n468 163.367
R952 B.n468 B.n89 163.367
R953 B.n464 B.n89 163.367
R954 B.n464 B.n463 163.367
R955 B.n463 B.n462 163.367
R956 B.n462 B.n91 163.367
R957 B.n458 B.n91 163.367
R958 B.n458 B.n457 163.367
R959 B.n457 B.n456 163.367
R960 B.n456 B.n93 163.367
R961 B.n452 B.n93 163.367
R962 B.n452 B.n451 163.367
R963 B.n451 B.n450 163.367
R964 B.n450 B.n95 163.367
R965 B.n446 B.n95 163.367
R966 B.n446 B.n445 163.367
R967 B.n445 B.n444 163.367
R968 B.n444 B.n97 163.367
R969 B.n440 B.n97 163.367
R970 B.n440 B.n439 163.367
R971 B.n439 B.n438 163.367
R972 B.n438 B.n99 163.367
R973 B.n434 B.n99 163.367
R974 B.n434 B.n433 163.367
R975 B.n433 B.n432 163.367
R976 B.n432 B.n101 163.367
R977 B.n428 B.n101 163.367
R978 B.n428 B.n427 163.367
R979 B.n427 B.n426 163.367
R980 B.n426 B.n103 163.367
R981 B.n422 B.n103 163.367
R982 B.n422 B.n421 163.367
R983 B.n421 B.n420 163.367
R984 B.n420 B.n105 163.367
R985 B.n416 B.n105 163.367
R986 B.n416 B.n415 163.367
R987 B.n415 B.n414 163.367
R988 B.n414 B.n107 163.367
R989 B.n410 B.n107 163.367
R990 B.n410 B.n409 163.367
R991 B.n409 B.n408 163.367
R992 B.n408 B.n109 163.367
R993 B.n404 B.n109 163.367
R994 B.n404 B.n403 163.367
R995 B.n403 B.n402 163.367
R996 B.n402 B.n111 163.367
R997 B.n398 B.n111 163.367
R998 B.n398 B.n397 163.367
R999 B.n397 B.n396 163.367
R1000 B.n396 B.n113 163.367
R1001 B.n392 B.n113 163.367
R1002 B.n392 B.n391 163.367
R1003 B.n391 B.n390 163.367
R1004 B.n390 B.n115 163.367
R1005 B.n386 B.n115 163.367
R1006 B.n386 B.n385 163.367
R1007 B.n385 B.n384 163.367
R1008 B.n384 B.n117 163.367
R1009 B.n380 B.n117 163.367
R1010 B.n380 B.n379 163.367
R1011 B.n379 B.n378 163.367
R1012 B.n378 B.n119 163.367
R1013 B.n374 B.n119 163.367
R1014 B.n374 B.n373 163.367
R1015 B.n373 B.n372 163.367
R1016 B.n372 B.n121 163.367
R1017 B.n636 B.n29 163.367
R1018 B.n632 B.n29 163.367
R1019 B.n632 B.n631 163.367
R1020 B.n631 B.n630 163.367
R1021 B.n630 B.n31 163.367
R1022 B.n626 B.n31 163.367
R1023 B.n626 B.n625 163.367
R1024 B.n625 B.n624 163.367
R1025 B.n624 B.n33 163.367
R1026 B.n620 B.n33 163.367
R1027 B.n620 B.n619 163.367
R1028 B.n619 B.n618 163.367
R1029 B.n618 B.n35 163.367
R1030 B.n614 B.n35 163.367
R1031 B.n614 B.n613 163.367
R1032 B.n613 B.n612 163.367
R1033 B.n612 B.n37 163.367
R1034 B.n608 B.n37 163.367
R1035 B.n608 B.n607 163.367
R1036 B.n607 B.n606 163.367
R1037 B.n606 B.n39 163.367
R1038 B.n602 B.n39 163.367
R1039 B.n602 B.n601 163.367
R1040 B.n601 B.n600 163.367
R1041 B.n600 B.n41 163.367
R1042 B.n596 B.n41 163.367
R1043 B.n596 B.n595 163.367
R1044 B.n595 B.n594 163.367
R1045 B.n594 B.n43 163.367
R1046 B.n589 B.n43 163.367
R1047 B.n589 B.n588 163.367
R1048 B.n588 B.n587 163.367
R1049 B.n587 B.n47 163.367
R1050 B.n583 B.n47 163.367
R1051 B.n583 B.n582 163.367
R1052 B.n582 B.n581 163.367
R1053 B.n581 B.n49 163.367
R1054 B.n577 B.n49 163.367
R1055 B.n577 B.n576 163.367
R1056 B.n576 B.n53 163.367
R1057 B.n572 B.n53 163.367
R1058 B.n572 B.n571 163.367
R1059 B.n571 B.n570 163.367
R1060 B.n570 B.n55 163.367
R1061 B.n566 B.n55 163.367
R1062 B.n566 B.n565 163.367
R1063 B.n565 B.n564 163.367
R1064 B.n564 B.n57 163.367
R1065 B.n560 B.n57 163.367
R1066 B.n560 B.n559 163.367
R1067 B.n559 B.n558 163.367
R1068 B.n558 B.n59 163.367
R1069 B.n554 B.n59 163.367
R1070 B.n554 B.n553 163.367
R1071 B.n553 B.n552 163.367
R1072 B.n552 B.n61 163.367
R1073 B.n548 B.n61 163.367
R1074 B.n548 B.n547 163.367
R1075 B.n547 B.n546 163.367
R1076 B.n546 B.n63 163.367
R1077 B.n542 B.n63 163.367
R1078 B.n542 B.n541 163.367
R1079 B.n541 B.n540 163.367
R1080 B.n540 B.n65 163.367
R1081 B.n536 B.n65 163.367
R1082 B.n536 B.n535 163.367
R1083 B.n535 B.n534 163.367
R1084 B.n534 B.n67 163.367
R1085 B.n638 B.n637 163.367
R1086 B.n638 B.n27 163.367
R1087 B.n642 B.n27 163.367
R1088 B.n643 B.n642 163.367
R1089 B.n644 B.n643 163.367
R1090 B.n644 B.n25 163.367
R1091 B.n648 B.n25 163.367
R1092 B.n649 B.n648 163.367
R1093 B.n650 B.n649 163.367
R1094 B.n650 B.n23 163.367
R1095 B.n654 B.n23 163.367
R1096 B.n655 B.n654 163.367
R1097 B.n656 B.n655 163.367
R1098 B.n656 B.n21 163.367
R1099 B.n660 B.n21 163.367
R1100 B.n661 B.n660 163.367
R1101 B.n662 B.n661 163.367
R1102 B.n662 B.n19 163.367
R1103 B.n666 B.n19 163.367
R1104 B.n667 B.n666 163.367
R1105 B.n668 B.n667 163.367
R1106 B.n668 B.n17 163.367
R1107 B.n672 B.n17 163.367
R1108 B.n673 B.n672 163.367
R1109 B.n674 B.n673 163.367
R1110 B.n674 B.n15 163.367
R1111 B.n678 B.n15 163.367
R1112 B.n679 B.n678 163.367
R1113 B.n680 B.n679 163.367
R1114 B.n680 B.n13 163.367
R1115 B.n684 B.n13 163.367
R1116 B.n685 B.n684 163.367
R1117 B.n686 B.n685 163.367
R1118 B.n686 B.n11 163.367
R1119 B.n690 B.n11 163.367
R1120 B.n691 B.n690 163.367
R1121 B.n692 B.n691 163.367
R1122 B.n692 B.n9 163.367
R1123 B.n696 B.n9 163.367
R1124 B.n697 B.n696 163.367
R1125 B.n698 B.n697 163.367
R1126 B.n698 B.n7 163.367
R1127 B.n702 B.n7 163.367
R1128 B.n703 B.n702 163.367
R1129 B.n704 B.n703 163.367
R1130 B.n704 B.n5 163.367
R1131 B.n708 B.n5 163.367
R1132 B.n709 B.n708 163.367
R1133 B.n710 B.n709 163.367
R1134 B.n710 B.n3 163.367
R1135 B.n714 B.n3 163.367
R1136 B.n715 B.n714 163.367
R1137 B.n184 B.n2 163.367
R1138 B.n184 B.n183 163.367
R1139 B.n188 B.n183 163.367
R1140 B.n189 B.n188 163.367
R1141 B.n190 B.n189 163.367
R1142 B.n190 B.n181 163.367
R1143 B.n194 B.n181 163.367
R1144 B.n195 B.n194 163.367
R1145 B.n196 B.n195 163.367
R1146 B.n196 B.n179 163.367
R1147 B.n200 B.n179 163.367
R1148 B.n201 B.n200 163.367
R1149 B.n202 B.n201 163.367
R1150 B.n202 B.n177 163.367
R1151 B.n206 B.n177 163.367
R1152 B.n207 B.n206 163.367
R1153 B.n208 B.n207 163.367
R1154 B.n208 B.n175 163.367
R1155 B.n212 B.n175 163.367
R1156 B.n213 B.n212 163.367
R1157 B.n214 B.n213 163.367
R1158 B.n214 B.n173 163.367
R1159 B.n218 B.n173 163.367
R1160 B.n219 B.n218 163.367
R1161 B.n220 B.n219 163.367
R1162 B.n220 B.n171 163.367
R1163 B.n224 B.n171 163.367
R1164 B.n225 B.n224 163.367
R1165 B.n226 B.n225 163.367
R1166 B.n226 B.n169 163.367
R1167 B.n230 B.n169 163.367
R1168 B.n231 B.n230 163.367
R1169 B.n232 B.n231 163.367
R1170 B.n232 B.n167 163.367
R1171 B.n236 B.n167 163.367
R1172 B.n237 B.n236 163.367
R1173 B.n238 B.n237 163.367
R1174 B.n238 B.n165 163.367
R1175 B.n242 B.n165 163.367
R1176 B.n243 B.n242 163.367
R1177 B.n244 B.n243 163.367
R1178 B.n244 B.n163 163.367
R1179 B.n248 B.n163 163.367
R1180 B.n249 B.n248 163.367
R1181 B.n250 B.n249 163.367
R1182 B.n250 B.n161 163.367
R1183 B.n254 B.n161 163.367
R1184 B.n255 B.n254 163.367
R1185 B.n256 B.n255 163.367
R1186 B.n256 B.n159 163.367
R1187 B.n260 B.n159 163.367
R1188 B.n261 B.n260 163.367
R1189 B.n143 B.n142 74.6672
R1190 B.n321 B.n320 74.6672
R1191 B.n51 B.n50 74.6672
R1192 B.n45 B.n44 74.6672
R1193 B.n307 B.n143 59.5399
R1194 B.n322 B.n321 59.5399
R1195 B.n52 B.n51 59.5399
R1196 B.n591 B.n45 59.5399
R1197 B.n635 B.n28 31.0639
R1198 B.n532 B.n531 31.0639
R1199 B.n370 B.n369 31.0639
R1200 B.n263 B.n158 31.0639
R1201 B B.n717 18.0485
R1202 B.n639 B.n28 10.6151
R1203 B.n640 B.n639 10.6151
R1204 B.n641 B.n640 10.6151
R1205 B.n641 B.n26 10.6151
R1206 B.n645 B.n26 10.6151
R1207 B.n646 B.n645 10.6151
R1208 B.n647 B.n646 10.6151
R1209 B.n647 B.n24 10.6151
R1210 B.n651 B.n24 10.6151
R1211 B.n652 B.n651 10.6151
R1212 B.n653 B.n652 10.6151
R1213 B.n653 B.n22 10.6151
R1214 B.n657 B.n22 10.6151
R1215 B.n658 B.n657 10.6151
R1216 B.n659 B.n658 10.6151
R1217 B.n659 B.n20 10.6151
R1218 B.n663 B.n20 10.6151
R1219 B.n664 B.n663 10.6151
R1220 B.n665 B.n664 10.6151
R1221 B.n665 B.n18 10.6151
R1222 B.n669 B.n18 10.6151
R1223 B.n670 B.n669 10.6151
R1224 B.n671 B.n670 10.6151
R1225 B.n671 B.n16 10.6151
R1226 B.n675 B.n16 10.6151
R1227 B.n676 B.n675 10.6151
R1228 B.n677 B.n676 10.6151
R1229 B.n677 B.n14 10.6151
R1230 B.n681 B.n14 10.6151
R1231 B.n682 B.n681 10.6151
R1232 B.n683 B.n682 10.6151
R1233 B.n683 B.n12 10.6151
R1234 B.n687 B.n12 10.6151
R1235 B.n688 B.n687 10.6151
R1236 B.n689 B.n688 10.6151
R1237 B.n689 B.n10 10.6151
R1238 B.n693 B.n10 10.6151
R1239 B.n694 B.n693 10.6151
R1240 B.n695 B.n694 10.6151
R1241 B.n695 B.n8 10.6151
R1242 B.n699 B.n8 10.6151
R1243 B.n700 B.n699 10.6151
R1244 B.n701 B.n700 10.6151
R1245 B.n701 B.n6 10.6151
R1246 B.n705 B.n6 10.6151
R1247 B.n706 B.n705 10.6151
R1248 B.n707 B.n706 10.6151
R1249 B.n707 B.n4 10.6151
R1250 B.n711 B.n4 10.6151
R1251 B.n712 B.n711 10.6151
R1252 B.n713 B.n712 10.6151
R1253 B.n713 B.n0 10.6151
R1254 B.n635 B.n634 10.6151
R1255 B.n634 B.n633 10.6151
R1256 B.n633 B.n30 10.6151
R1257 B.n629 B.n30 10.6151
R1258 B.n629 B.n628 10.6151
R1259 B.n628 B.n627 10.6151
R1260 B.n627 B.n32 10.6151
R1261 B.n623 B.n32 10.6151
R1262 B.n623 B.n622 10.6151
R1263 B.n622 B.n621 10.6151
R1264 B.n621 B.n34 10.6151
R1265 B.n617 B.n34 10.6151
R1266 B.n617 B.n616 10.6151
R1267 B.n616 B.n615 10.6151
R1268 B.n615 B.n36 10.6151
R1269 B.n611 B.n36 10.6151
R1270 B.n611 B.n610 10.6151
R1271 B.n610 B.n609 10.6151
R1272 B.n609 B.n38 10.6151
R1273 B.n605 B.n38 10.6151
R1274 B.n605 B.n604 10.6151
R1275 B.n604 B.n603 10.6151
R1276 B.n603 B.n40 10.6151
R1277 B.n599 B.n40 10.6151
R1278 B.n599 B.n598 10.6151
R1279 B.n598 B.n597 10.6151
R1280 B.n597 B.n42 10.6151
R1281 B.n593 B.n42 10.6151
R1282 B.n593 B.n592 10.6151
R1283 B.n590 B.n46 10.6151
R1284 B.n586 B.n46 10.6151
R1285 B.n586 B.n585 10.6151
R1286 B.n585 B.n584 10.6151
R1287 B.n584 B.n48 10.6151
R1288 B.n580 B.n48 10.6151
R1289 B.n580 B.n579 10.6151
R1290 B.n579 B.n578 10.6151
R1291 B.n575 B.n574 10.6151
R1292 B.n574 B.n573 10.6151
R1293 B.n573 B.n54 10.6151
R1294 B.n569 B.n54 10.6151
R1295 B.n569 B.n568 10.6151
R1296 B.n568 B.n567 10.6151
R1297 B.n567 B.n56 10.6151
R1298 B.n563 B.n56 10.6151
R1299 B.n563 B.n562 10.6151
R1300 B.n562 B.n561 10.6151
R1301 B.n561 B.n58 10.6151
R1302 B.n557 B.n58 10.6151
R1303 B.n557 B.n556 10.6151
R1304 B.n556 B.n555 10.6151
R1305 B.n555 B.n60 10.6151
R1306 B.n551 B.n60 10.6151
R1307 B.n551 B.n550 10.6151
R1308 B.n550 B.n549 10.6151
R1309 B.n549 B.n62 10.6151
R1310 B.n545 B.n62 10.6151
R1311 B.n545 B.n544 10.6151
R1312 B.n544 B.n543 10.6151
R1313 B.n543 B.n64 10.6151
R1314 B.n539 B.n64 10.6151
R1315 B.n539 B.n538 10.6151
R1316 B.n538 B.n537 10.6151
R1317 B.n537 B.n66 10.6151
R1318 B.n533 B.n66 10.6151
R1319 B.n533 B.n532 10.6151
R1320 B.n531 B.n68 10.6151
R1321 B.n527 B.n68 10.6151
R1322 B.n527 B.n526 10.6151
R1323 B.n526 B.n525 10.6151
R1324 B.n525 B.n70 10.6151
R1325 B.n521 B.n70 10.6151
R1326 B.n521 B.n520 10.6151
R1327 B.n520 B.n519 10.6151
R1328 B.n519 B.n72 10.6151
R1329 B.n515 B.n72 10.6151
R1330 B.n515 B.n514 10.6151
R1331 B.n514 B.n513 10.6151
R1332 B.n513 B.n74 10.6151
R1333 B.n509 B.n74 10.6151
R1334 B.n509 B.n508 10.6151
R1335 B.n508 B.n507 10.6151
R1336 B.n507 B.n76 10.6151
R1337 B.n503 B.n76 10.6151
R1338 B.n503 B.n502 10.6151
R1339 B.n502 B.n501 10.6151
R1340 B.n501 B.n78 10.6151
R1341 B.n497 B.n78 10.6151
R1342 B.n497 B.n496 10.6151
R1343 B.n496 B.n495 10.6151
R1344 B.n495 B.n80 10.6151
R1345 B.n491 B.n80 10.6151
R1346 B.n491 B.n490 10.6151
R1347 B.n490 B.n489 10.6151
R1348 B.n489 B.n82 10.6151
R1349 B.n485 B.n82 10.6151
R1350 B.n485 B.n484 10.6151
R1351 B.n484 B.n483 10.6151
R1352 B.n483 B.n84 10.6151
R1353 B.n479 B.n84 10.6151
R1354 B.n479 B.n478 10.6151
R1355 B.n478 B.n477 10.6151
R1356 B.n477 B.n86 10.6151
R1357 B.n473 B.n86 10.6151
R1358 B.n473 B.n472 10.6151
R1359 B.n472 B.n471 10.6151
R1360 B.n471 B.n88 10.6151
R1361 B.n467 B.n88 10.6151
R1362 B.n467 B.n466 10.6151
R1363 B.n466 B.n465 10.6151
R1364 B.n465 B.n90 10.6151
R1365 B.n461 B.n90 10.6151
R1366 B.n461 B.n460 10.6151
R1367 B.n460 B.n459 10.6151
R1368 B.n459 B.n92 10.6151
R1369 B.n455 B.n92 10.6151
R1370 B.n455 B.n454 10.6151
R1371 B.n454 B.n453 10.6151
R1372 B.n453 B.n94 10.6151
R1373 B.n449 B.n94 10.6151
R1374 B.n449 B.n448 10.6151
R1375 B.n448 B.n447 10.6151
R1376 B.n447 B.n96 10.6151
R1377 B.n443 B.n96 10.6151
R1378 B.n443 B.n442 10.6151
R1379 B.n442 B.n441 10.6151
R1380 B.n441 B.n98 10.6151
R1381 B.n437 B.n98 10.6151
R1382 B.n437 B.n436 10.6151
R1383 B.n436 B.n435 10.6151
R1384 B.n435 B.n100 10.6151
R1385 B.n431 B.n100 10.6151
R1386 B.n431 B.n430 10.6151
R1387 B.n430 B.n429 10.6151
R1388 B.n429 B.n102 10.6151
R1389 B.n425 B.n102 10.6151
R1390 B.n425 B.n424 10.6151
R1391 B.n424 B.n423 10.6151
R1392 B.n423 B.n104 10.6151
R1393 B.n419 B.n104 10.6151
R1394 B.n419 B.n418 10.6151
R1395 B.n418 B.n417 10.6151
R1396 B.n417 B.n106 10.6151
R1397 B.n413 B.n106 10.6151
R1398 B.n413 B.n412 10.6151
R1399 B.n412 B.n411 10.6151
R1400 B.n411 B.n108 10.6151
R1401 B.n407 B.n108 10.6151
R1402 B.n407 B.n406 10.6151
R1403 B.n406 B.n405 10.6151
R1404 B.n405 B.n110 10.6151
R1405 B.n401 B.n110 10.6151
R1406 B.n401 B.n400 10.6151
R1407 B.n400 B.n399 10.6151
R1408 B.n399 B.n112 10.6151
R1409 B.n395 B.n112 10.6151
R1410 B.n395 B.n394 10.6151
R1411 B.n394 B.n393 10.6151
R1412 B.n393 B.n114 10.6151
R1413 B.n389 B.n114 10.6151
R1414 B.n389 B.n388 10.6151
R1415 B.n388 B.n387 10.6151
R1416 B.n387 B.n116 10.6151
R1417 B.n383 B.n116 10.6151
R1418 B.n383 B.n382 10.6151
R1419 B.n382 B.n381 10.6151
R1420 B.n381 B.n118 10.6151
R1421 B.n377 B.n118 10.6151
R1422 B.n377 B.n376 10.6151
R1423 B.n376 B.n375 10.6151
R1424 B.n375 B.n120 10.6151
R1425 B.n371 B.n120 10.6151
R1426 B.n371 B.n370 10.6151
R1427 B.n185 B.n1 10.6151
R1428 B.n186 B.n185 10.6151
R1429 B.n187 B.n186 10.6151
R1430 B.n187 B.n182 10.6151
R1431 B.n191 B.n182 10.6151
R1432 B.n192 B.n191 10.6151
R1433 B.n193 B.n192 10.6151
R1434 B.n193 B.n180 10.6151
R1435 B.n197 B.n180 10.6151
R1436 B.n198 B.n197 10.6151
R1437 B.n199 B.n198 10.6151
R1438 B.n199 B.n178 10.6151
R1439 B.n203 B.n178 10.6151
R1440 B.n204 B.n203 10.6151
R1441 B.n205 B.n204 10.6151
R1442 B.n205 B.n176 10.6151
R1443 B.n209 B.n176 10.6151
R1444 B.n210 B.n209 10.6151
R1445 B.n211 B.n210 10.6151
R1446 B.n211 B.n174 10.6151
R1447 B.n215 B.n174 10.6151
R1448 B.n216 B.n215 10.6151
R1449 B.n217 B.n216 10.6151
R1450 B.n217 B.n172 10.6151
R1451 B.n221 B.n172 10.6151
R1452 B.n222 B.n221 10.6151
R1453 B.n223 B.n222 10.6151
R1454 B.n223 B.n170 10.6151
R1455 B.n227 B.n170 10.6151
R1456 B.n228 B.n227 10.6151
R1457 B.n229 B.n228 10.6151
R1458 B.n229 B.n168 10.6151
R1459 B.n233 B.n168 10.6151
R1460 B.n234 B.n233 10.6151
R1461 B.n235 B.n234 10.6151
R1462 B.n235 B.n166 10.6151
R1463 B.n239 B.n166 10.6151
R1464 B.n240 B.n239 10.6151
R1465 B.n241 B.n240 10.6151
R1466 B.n241 B.n164 10.6151
R1467 B.n245 B.n164 10.6151
R1468 B.n246 B.n245 10.6151
R1469 B.n247 B.n246 10.6151
R1470 B.n247 B.n162 10.6151
R1471 B.n251 B.n162 10.6151
R1472 B.n252 B.n251 10.6151
R1473 B.n253 B.n252 10.6151
R1474 B.n253 B.n160 10.6151
R1475 B.n257 B.n160 10.6151
R1476 B.n258 B.n257 10.6151
R1477 B.n259 B.n258 10.6151
R1478 B.n259 B.n158 10.6151
R1479 B.n264 B.n263 10.6151
R1480 B.n265 B.n264 10.6151
R1481 B.n265 B.n156 10.6151
R1482 B.n269 B.n156 10.6151
R1483 B.n270 B.n269 10.6151
R1484 B.n271 B.n270 10.6151
R1485 B.n271 B.n154 10.6151
R1486 B.n275 B.n154 10.6151
R1487 B.n276 B.n275 10.6151
R1488 B.n277 B.n276 10.6151
R1489 B.n277 B.n152 10.6151
R1490 B.n281 B.n152 10.6151
R1491 B.n282 B.n281 10.6151
R1492 B.n283 B.n282 10.6151
R1493 B.n283 B.n150 10.6151
R1494 B.n287 B.n150 10.6151
R1495 B.n288 B.n287 10.6151
R1496 B.n289 B.n288 10.6151
R1497 B.n289 B.n148 10.6151
R1498 B.n293 B.n148 10.6151
R1499 B.n294 B.n293 10.6151
R1500 B.n295 B.n294 10.6151
R1501 B.n295 B.n146 10.6151
R1502 B.n299 B.n146 10.6151
R1503 B.n300 B.n299 10.6151
R1504 B.n301 B.n300 10.6151
R1505 B.n301 B.n144 10.6151
R1506 B.n305 B.n144 10.6151
R1507 B.n306 B.n305 10.6151
R1508 B.n308 B.n140 10.6151
R1509 B.n312 B.n140 10.6151
R1510 B.n313 B.n312 10.6151
R1511 B.n314 B.n313 10.6151
R1512 B.n314 B.n138 10.6151
R1513 B.n318 B.n138 10.6151
R1514 B.n319 B.n318 10.6151
R1515 B.n323 B.n319 10.6151
R1516 B.n327 B.n136 10.6151
R1517 B.n328 B.n327 10.6151
R1518 B.n329 B.n328 10.6151
R1519 B.n329 B.n134 10.6151
R1520 B.n333 B.n134 10.6151
R1521 B.n334 B.n333 10.6151
R1522 B.n335 B.n334 10.6151
R1523 B.n335 B.n132 10.6151
R1524 B.n339 B.n132 10.6151
R1525 B.n340 B.n339 10.6151
R1526 B.n341 B.n340 10.6151
R1527 B.n341 B.n130 10.6151
R1528 B.n345 B.n130 10.6151
R1529 B.n346 B.n345 10.6151
R1530 B.n347 B.n346 10.6151
R1531 B.n347 B.n128 10.6151
R1532 B.n351 B.n128 10.6151
R1533 B.n352 B.n351 10.6151
R1534 B.n353 B.n352 10.6151
R1535 B.n353 B.n126 10.6151
R1536 B.n357 B.n126 10.6151
R1537 B.n358 B.n357 10.6151
R1538 B.n359 B.n358 10.6151
R1539 B.n359 B.n124 10.6151
R1540 B.n363 B.n124 10.6151
R1541 B.n364 B.n363 10.6151
R1542 B.n365 B.n364 10.6151
R1543 B.n365 B.n122 10.6151
R1544 B.n369 B.n122 10.6151
R1545 B.n717 B.n0 8.11757
R1546 B.n717 B.n1 8.11757
R1547 B.n591 B.n590 6.4005
R1548 B.n578 B.n52 6.4005
R1549 B.n308 B.n307 6.4005
R1550 B.n323 B.n322 6.4005
R1551 B.n592 B.n591 4.21513
R1552 B.n575 B.n52 4.21513
R1553 B.n307 B.n306 4.21513
R1554 B.n322 B.n136 4.21513
R1555 VP.n16 VP.n13 161.3
R1556 VP.n18 VP.n17 161.3
R1557 VP.n19 VP.n12 161.3
R1558 VP.n21 VP.n20 161.3
R1559 VP.n22 VP.n11 161.3
R1560 VP.n24 VP.n23 161.3
R1561 VP.n25 VP.n10 161.3
R1562 VP.n27 VP.n26 161.3
R1563 VP.n55 VP.n54 161.3
R1564 VP.n53 VP.n1 161.3
R1565 VP.n52 VP.n51 161.3
R1566 VP.n50 VP.n2 161.3
R1567 VP.n49 VP.n48 161.3
R1568 VP.n47 VP.n3 161.3
R1569 VP.n46 VP.n45 161.3
R1570 VP.n44 VP.n4 161.3
R1571 VP.n43 VP.n42 161.3
R1572 VP.n40 VP.n5 161.3
R1573 VP.n39 VP.n38 161.3
R1574 VP.n37 VP.n6 161.3
R1575 VP.n36 VP.n35 161.3
R1576 VP.n34 VP.n7 161.3
R1577 VP.n33 VP.n32 161.3
R1578 VP.n31 VP.n8 161.3
R1579 VP.n15 VP.t5 86.6954
R1580 VP.n30 VP.n29 85.0223
R1581 VP.n56 VP.n0 85.0223
R1582 VP.n28 VP.n9 85.0223
R1583 VP.n15 VP.n14 62.0356
R1584 VP.n35 VP.n6 56.4773
R1585 VP.n48 VP.n2 56.4773
R1586 VP.n20 VP.n11 56.4773
R1587 VP.n29 VP.t1 54.3624
R1588 VP.n41 VP.t4 54.3624
R1589 VP.n0 VP.t3 54.3624
R1590 VP.n9 VP.t0 54.3624
R1591 VP.n14 VP.t2 54.3624
R1592 VP.n30 VP.n28 49.2226
R1593 VP.n33 VP.n8 24.3439
R1594 VP.n34 VP.n33 24.3439
R1595 VP.n35 VP.n34 24.3439
R1596 VP.n39 VP.n6 24.3439
R1597 VP.n40 VP.n39 24.3439
R1598 VP.n42 VP.n40 24.3439
R1599 VP.n46 VP.n4 24.3439
R1600 VP.n47 VP.n46 24.3439
R1601 VP.n48 VP.n47 24.3439
R1602 VP.n52 VP.n2 24.3439
R1603 VP.n53 VP.n52 24.3439
R1604 VP.n54 VP.n53 24.3439
R1605 VP.n24 VP.n11 24.3439
R1606 VP.n25 VP.n24 24.3439
R1607 VP.n26 VP.n25 24.3439
R1608 VP.n18 VP.n13 24.3439
R1609 VP.n19 VP.n18 24.3439
R1610 VP.n20 VP.n19 24.3439
R1611 VP.n42 VP.n41 12.1722
R1612 VP.n41 VP.n4 12.1722
R1613 VP.n14 VP.n13 12.1722
R1614 VP.n29 VP.n8 4.86919
R1615 VP.n54 VP.n0 4.86919
R1616 VP.n26 VP.n9 4.86919
R1617 VP.n16 VP.n15 3.33649
R1618 VP.n28 VP.n27 0.355081
R1619 VP.n31 VP.n30 0.355081
R1620 VP.n56 VP.n55 0.355081
R1621 VP VP.n56 0.26685
R1622 VP.n17 VP.n16 0.189894
R1623 VP.n17 VP.n12 0.189894
R1624 VP.n21 VP.n12 0.189894
R1625 VP.n22 VP.n21 0.189894
R1626 VP.n23 VP.n22 0.189894
R1627 VP.n23 VP.n10 0.189894
R1628 VP.n27 VP.n10 0.189894
R1629 VP.n32 VP.n31 0.189894
R1630 VP.n32 VP.n7 0.189894
R1631 VP.n36 VP.n7 0.189894
R1632 VP.n37 VP.n36 0.189894
R1633 VP.n38 VP.n37 0.189894
R1634 VP.n38 VP.n5 0.189894
R1635 VP.n43 VP.n5 0.189894
R1636 VP.n44 VP.n43 0.189894
R1637 VP.n45 VP.n44 0.189894
R1638 VP.n45 VP.n3 0.189894
R1639 VP.n49 VP.n3 0.189894
R1640 VP.n50 VP.n49 0.189894
R1641 VP.n51 VP.n50 0.189894
R1642 VP.n51 VP.n1 0.189894
R1643 VP.n55 VP.n1 0.189894
R1644 VDD1.n36 VDD1.n0 756.745
R1645 VDD1.n77 VDD1.n41 756.745
R1646 VDD1.n37 VDD1.n36 585
R1647 VDD1.n35 VDD1.n2 585
R1648 VDD1.n34 VDD1.n33 585
R1649 VDD1.n5 VDD1.n3 585
R1650 VDD1.n28 VDD1.n27 585
R1651 VDD1.n26 VDD1.n25 585
R1652 VDD1.n9 VDD1.n8 585
R1653 VDD1.n20 VDD1.n19 585
R1654 VDD1.n18 VDD1.n17 585
R1655 VDD1.n13 VDD1.n12 585
R1656 VDD1.n53 VDD1.n52 585
R1657 VDD1.n58 VDD1.n57 585
R1658 VDD1.n60 VDD1.n59 585
R1659 VDD1.n49 VDD1.n48 585
R1660 VDD1.n66 VDD1.n65 585
R1661 VDD1.n68 VDD1.n67 585
R1662 VDD1.n45 VDD1.n44 585
R1663 VDD1.n75 VDD1.n74 585
R1664 VDD1.n76 VDD1.n43 585
R1665 VDD1.n78 VDD1.n77 585
R1666 VDD1.n14 VDD1.t0 329.043
R1667 VDD1.n54 VDD1.t4 329.043
R1668 VDD1.n36 VDD1.n35 171.744
R1669 VDD1.n35 VDD1.n34 171.744
R1670 VDD1.n34 VDD1.n3 171.744
R1671 VDD1.n27 VDD1.n3 171.744
R1672 VDD1.n27 VDD1.n26 171.744
R1673 VDD1.n26 VDD1.n8 171.744
R1674 VDD1.n19 VDD1.n8 171.744
R1675 VDD1.n19 VDD1.n18 171.744
R1676 VDD1.n18 VDD1.n12 171.744
R1677 VDD1.n58 VDD1.n52 171.744
R1678 VDD1.n59 VDD1.n58 171.744
R1679 VDD1.n59 VDD1.n48 171.744
R1680 VDD1.n66 VDD1.n48 171.744
R1681 VDD1.n67 VDD1.n66 171.744
R1682 VDD1.n67 VDD1.n44 171.744
R1683 VDD1.n75 VDD1.n44 171.744
R1684 VDD1.n76 VDD1.n75 171.744
R1685 VDD1.n77 VDD1.n76 171.744
R1686 VDD1.t0 VDD1.n12 85.8723
R1687 VDD1.t4 VDD1.n52 85.8723
R1688 VDD1.n83 VDD1.n82 85.8486
R1689 VDD1.n85 VDD1.n84 85.0742
R1690 VDD1 VDD1.n40 54.1267
R1691 VDD1.n83 VDD1.n81 54.0132
R1692 VDD1.n85 VDD1.n83 43.5892
R1693 VDD1.n37 VDD1.n2 13.1884
R1694 VDD1.n78 VDD1.n43 13.1884
R1695 VDD1.n38 VDD1.n0 12.8005
R1696 VDD1.n33 VDD1.n4 12.8005
R1697 VDD1.n74 VDD1.n73 12.8005
R1698 VDD1.n79 VDD1.n41 12.8005
R1699 VDD1.n32 VDD1.n5 12.0247
R1700 VDD1.n72 VDD1.n45 12.0247
R1701 VDD1.n29 VDD1.n28 11.249
R1702 VDD1.n69 VDD1.n68 11.249
R1703 VDD1.n14 VDD1.n13 10.7238
R1704 VDD1.n54 VDD1.n53 10.7238
R1705 VDD1.n25 VDD1.n7 10.4732
R1706 VDD1.n65 VDD1.n47 10.4732
R1707 VDD1.n24 VDD1.n9 9.69747
R1708 VDD1.n64 VDD1.n49 9.69747
R1709 VDD1.n40 VDD1.n39 9.45567
R1710 VDD1.n81 VDD1.n80 9.45567
R1711 VDD1.n16 VDD1.n15 9.3005
R1712 VDD1.n11 VDD1.n10 9.3005
R1713 VDD1.n22 VDD1.n21 9.3005
R1714 VDD1.n24 VDD1.n23 9.3005
R1715 VDD1.n7 VDD1.n6 9.3005
R1716 VDD1.n30 VDD1.n29 9.3005
R1717 VDD1.n32 VDD1.n31 9.3005
R1718 VDD1.n4 VDD1.n1 9.3005
R1719 VDD1.n39 VDD1.n38 9.3005
R1720 VDD1.n80 VDD1.n79 9.3005
R1721 VDD1.n56 VDD1.n55 9.3005
R1722 VDD1.n51 VDD1.n50 9.3005
R1723 VDD1.n62 VDD1.n61 9.3005
R1724 VDD1.n64 VDD1.n63 9.3005
R1725 VDD1.n47 VDD1.n46 9.3005
R1726 VDD1.n70 VDD1.n69 9.3005
R1727 VDD1.n72 VDD1.n71 9.3005
R1728 VDD1.n73 VDD1.n42 9.3005
R1729 VDD1.n21 VDD1.n20 8.92171
R1730 VDD1.n61 VDD1.n60 8.92171
R1731 VDD1.n17 VDD1.n11 8.14595
R1732 VDD1.n57 VDD1.n51 8.14595
R1733 VDD1.n16 VDD1.n13 7.3702
R1734 VDD1.n56 VDD1.n53 7.3702
R1735 VDD1.n17 VDD1.n16 5.81868
R1736 VDD1.n57 VDD1.n56 5.81868
R1737 VDD1.n20 VDD1.n11 5.04292
R1738 VDD1.n60 VDD1.n51 5.04292
R1739 VDD1.n21 VDD1.n9 4.26717
R1740 VDD1.n61 VDD1.n49 4.26717
R1741 VDD1.n84 VDD1.t3 4.09433
R1742 VDD1.n84 VDD1.t5 4.09433
R1743 VDD1.n82 VDD1.t1 4.09433
R1744 VDD1.n82 VDD1.t2 4.09433
R1745 VDD1.n25 VDD1.n24 3.49141
R1746 VDD1.n65 VDD1.n64 3.49141
R1747 VDD1.n28 VDD1.n7 2.71565
R1748 VDD1.n68 VDD1.n47 2.71565
R1749 VDD1.n15 VDD1.n14 2.4129
R1750 VDD1.n55 VDD1.n54 2.4129
R1751 VDD1.n29 VDD1.n5 1.93989
R1752 VDD1.n69 VDD1.n45 1.93989
R1753 VDD1.n40 VDD1.n0 1.16414
R1754 VDD1.n33 VDD1.n32 1.16414
R1755 VDD1.n74 VDD1.n72 1.16414
R1756 VDD1.n81 VDD1.n41 1.16414
R1757 VDD1 VDD1.n85 0.772052
R1758 VDD1.n38 VDD1.n37 0.388379
R1759 VDD1.n4 VDD1.n2 0.388379
R1760 VDD1.n73 VDD1.n43 0.388379
R1761 VDD1.n79 VDD1.n78 0.388379
R1762 VDD1.n39 VDD1.n1 0.155672
R1763 VDD1.n31 VDD1.n1 0.155672
R1764 VDD1.n31 VDD1.n30 0.155672
R1765 VDD1.n30 VDD1.n6 0.155672
R1766 VDD1.n23 VDD1.n6 0.155672
R1767 VDD1.n23 VDD1.n22 0.155672
R1768 VDD1.n22 VDD1.n10 0.155672
R1769 VDD1.n15 VDD1.n10 0.155672
R1770 VDD1.n55 VDD1.n50 0.155672
R1771 VDD1.n62 VDD1.n50 0.155672
R1772 VDD1.n63 VDD1.n62 0.155672
R1773 VDD1.n63 VDD1.n46 0.155672
R1774 VDD1.n70 VDD1.n46 0.155672
R1775 VDD1.n71 VDD1.n70 0.155672
R1776 VDD1.n71 VDD1.n42 0.155672
R1777 VDD1.n80 VDD1.n42 0.155672
C0 VN B 1.31465f
C1 VP VN 7.07924f
C2 VN VTAIL 5.38779f
C3 VP B 2.19778f
C4 VDD1 VN 0.151783f
C5 VN w_n4050_n2556# 7.8473f
C6 VTAIL B 3.08598f
C7 VDD1 B 2.00609f
C8 w_n4050_n2556# B 9.82483f
C9 VP VTAIL 5.40197f
C10 VP VDD1 5.19364f
C11 VP w_n4050_n2556# 8.373469f
C12 VDD1 VTAIL 6.70692f
C13 w_n4050_n2556# VTAIL 2.49906f
C14 VDD1 w_n4050_n2556# 2.23747f
C15 VDD2 VN 4.81207f
C16 VDD2 B 2.10225f
C17 VDD2 VP 0.535879f
C18 VDD2 VTAIL 6.7654f
C19 VDD2 VDD1 1.76624f
C20 VDD2 w_n4050_n2556# 2.35196f
C21 VDD2 VSUBS 2.048982f
C22 VDD1 VSUBS 2.061688f
C23 VTAIL VSUBS 1.234345f
C24 VN VSUBS 6.68109f
C25 VP VSUBS 3.507689f
C26 B VSUBS 5.20516f
C27 w_n4050_n2556# VSUBS 0.12845p
C28 VDD1.n0 VSUBS 0.031449f
C29 VDD1.n1 VSUBS 0.029888f
C30 VDD1.n2 VSUBS 0.016533f
C31 VDD1.n3 VSUBS 0.037961f
C32 VDD1.n4 VSUBS 0.016061f
C33 VDD1.n5 VSUBS 0.017005f
C34 VDD1.n6 VSUBS 0.029888f
C35 VDD1.n7 VSUBS 0.016061f
C36 VDD1.n8 VSUBS 0.037961f
C37 VDD1.n9 VSUBS 0.017005f
C38 VDD1.n10 VSUBS 0.029888f
C39 VDD1.n11 VSUBS 0.016061f
C40 VDD1.n12 VSUBS 0.028471f
C41 VDD1.n13 VSUBS 0.028556f
C42 VDD1.t0 VSUBS 0.081531f
C43 VDD1.n14 VSUBS 0.180635f
C44 VDD1.n15 VSUBS 0.936558f
C45 VDD1.n16 VSUBS 0.016061f
C46 VDD1.n17 VSUBS 0.017005f
C47 VDD1.n18 VSUBS 0.037961f
C48 VDD1.n19 VSUBS 0.037961f
C49 VDD1.n20 VSUBS 0.017005f
C50 VDD1.n21 VSUBS 0.016061f
C51 VDD1.n22 VSUBS 0.029888f
C52 VDD1.n23 VSUBS 0.029888f
C53 VDD1.n24 VSUBS 0.016061f
C54 VDD1.n25 VSUBS 0.017005f
C55 VDD1.n26 VSUBS 0.037961f
C56 VDD1.n27 VSUBS 0.037961f
C57 VDD1.n28 VSUBS 0.017005f
C58 VDD1.n29 VSUBS 0.016061f
C59 VDD1.n30 VSUBS 0.029888f
C60 VDD1.n31 VSUBS 0.029888f
C61 VDD1.n32 VSUBS 0.016061f
C62 VDD1.n33 VSUBS 0.017005f
C63 VDD1.n34 VSUBS 0.037961f
C64 VDD1.n35 VSUBS 0.037961f
C65 VDD1.n36 VSUBS 0.087159f
C66 VDD1.n37 VSUBS 0.016533f
C67 VDD1.n38 VSUBS 0.016061f
C68 VDD1.n39 VSUBS 0.074801f
C69 VDD1.n40 VSUBS 0.078796f
C70 VDD1.n41 VSUBS 0.031449f
C71 VDD1.n42 VSUBS 0.029888f
C72 VDD1.n43 VSUBS 0.016533f
C73 VDD1.n44 VSUBS 0.037961f
C74 VDD1.n45 VSUBS 0.017005f
C75 VDD1.n46 VSUBS 0.029888f
C76 VDD1.n47 VSUBS 0.016061f
C77 VDD1.n48 VSUBS 0.037961f
C78 VDD1.n49 VSUBS 0.017005f
C79 VDD1.n50 VSUBS 0.029888f
C80 VDD1.n51 VSUBS 0.016061f
C81 VDD1.n52 VSUBS 0.028471f
C82 VDD1.n53 VSUBS 0.028556f
C83 VDD1.t4 VSUBS 0.081531f
C84 VDD1.n54 VSUBS 0.180635f
C85 VDD1.n55 VSUBS 0.936557f
C86 VDD1.n56 VSUBS 0.016061f
C87 VDD1.n57 VSUBS 0.017005f
C88 VDD1.n58 VSUBS 0.037961f
C89 VDD1.n59 VSUBS 0.037961f
C90 VDD1.n60 VSUBS 0.017005f
C91 VDD1.n61 VSUBS 0.016061f
C92 VDD1.n62 VSUBS 0.029888f
C93 VDD1.n63 VSUBS 0.029888f
C94 VDD1.n64 VSUBS 0.016061f
C95 VDD1.n65 VSUBS 0.017005f
C96 VDD1.n66 VSUBS 0.037961f
C97 VDD1.n67 VSUBS 0.037961f
C98 VDD1.n68 VSUBS 0.017005f
C99 VDD1.n69 VSUBS 0.016061f
C100 VDD1.n70 VSUBS 0.029888f
C101 VDD1.n71 VSUBS 0.029888f
C102 VDD1.n72 VSUBS 0.016061f
C103 VDD1.n73 VSUBS 0.016061f
C104 VDD1.n74 VSUBS 0.017005f
C105 VDD1.n75 VSUBS 0.037961f
C106 VDD1.n76 VSUBS 0.037961f
C107 VDD1.n77 VSUBS 0.087159f
C108 VDD1.n78 VSUBS 0.016533f
C109 VDD1.n79 VSUBS 0.016061f
C110 VDD1.n80 VSUBS 0.074801f
C111 VDD1.n81 VSUBS 0.077703f
C112 VDD1.t1 VSUBS 0.187532f
C113 VDD1.t2 VSUBS 0.187532f
C114 VDD1.n82 VSUBS 1.36544f
C115 VDD1.n83 VSUBS 3.81125f
C116 VDD1.t3 VSUBS 0.187532f
C117 VDD1.t5 VSUBS 0.187532f
C118 VDD1.n84 VSUBS 1.35723f
C119 VDD1.n85 VSUBS 3.53063f
C120 VP.t3 VSUBS 2.54077f
C121 VP.n0 VSUBS 1.03879f
C122 VP.n1 VSUBS 0.03389f
C123 VP.n2 VSUBS 0.056821f
C124 VP.n3 VSUBS 0.03389f
C125 VP.n4 VSUBS 0.047808f
C126 VP.n5 VSUBS 0.03389f
C127 VP.n6 VSUBS 0.042555f
C128 VP.n7 VSUBS 0.03389f
C129 VP.n8 VSUBS 0.038405f
C130 VP.t0 VSUBS 2.54077f
C131 VP.n9 VSUBS 1.03879f
C132 VP.n10 VSUBS 0.03389f
C133 VP.n11 VSUBS 0.056821f
C134 VP.n12 VSUBS 0.03389f
C135 VP.n13 VSUBS 0.047808f
C136 VP.t5 VSUBS 2.97696f
C137 VP.t2 VSUBS 2.54077f
C138 VP.n14 VSUBS 1.03337f
C139 VP.n15 VSUBS 0.989189f
C140 VP.n16 VSUBS 0.422291f
C141 VP.n17 VSUBS 0.03389f
C142 VP.n18 VSUBS 0.063478f
C143 VP.n19 VSUBS 0.063478f
C144 VP.n20 VSUBS 0.042555f
C145 VP.n21 VSUBS 0.03389f
C146 VP.n22 VSUBS 0.03389f
C147 VP.n23 VSUBS 0.03389f
C148 VP.n24 VSUBS 0.063478f
C149 VP.n25 VSUBS 0.063478f
C150 VP.n26 VSUBS 0.038405f
C151 VP.n27 VSUBS 0.054706f
C152 VP.n28 VSUBS 1.89797f
C153 VP.t1 VSUBS 2.54077f
C154 VP.n29 VSUBS 1.03879f
C155 VP.n30 VSUBS 1.92265f
C156 VP.n31 VSUBS 0.054706f
C157 VP.n32 VSUBS 0.03389f
C158 VP.n33 VSUBS 0.063478f
C159 VP.n34 VSUBS 0.063478f
C160 VP.n35 VSUBS 0.056821f
C161 VP.n36 VSUBS 0.03389f
C162 VP.n37 VSUBS 0.03389f
C163 VP.n38 VSUBS 0.03389f
C164 VP.n39 VSUBS 0.063478f
C165 VP.n40 VSUBS 0.063478f
C166 VP.t4 VSUBS 2.54077f
C167 VP.n41 VSUBS 0.916153f
C168 VP.n42 VSUBS 0.047808f
C169 VP.n43 VSUBS 0.03389f
C170 VP.n44 VSUBS 0.03389f
C171 VP.n45 VSUBS 0.03389f
C172 VP.n46 VSUBS 0.063478f
C173 VP.n47 VSUBS 0.063478f
C174 VP.n48 VSUBS 0.042555f
C175 VP.n49 VSUBS 0.03389f
C176 VP.n50 VSUBS 0.03389f
C177 VP.n51 VSUBS 0.03389f
C178 VP.n52 VSUBS 0.063478f
C179 VP.n53 VSUBS 0.063478f
C180 VP.n54 VSUBS 0.038405f
C181 VP.n55 VSUBS 0.054706f
C182 VP.n56 VSUBS 0.097058f
C183 B.n0 VSUBS 0.008821f
C184 B.n1 VSUBS 0.008821f
C185 B.n2 VSUBS 0.013046f
C186 B.n3 VSUBS 0.009997f
C187 B.n4 VSUBS 0.009997f
C188 B.n5 VSUBS 0.009997f
C189 B.n6 VSUBS 0.009997f
C190 B.n7 VSUBS 0.009997f
C191 B.n8 VSUBS 0.009997f
C192 B.n9 VSUBS 0.009997f
C193 B.n10 VSUBS 0.009997f
C194 B.n11 VSUBS 0.009997f
C195 B.n12 VSUBS 0.009997f
C196 B.n13 VSUBS 0.009997f
C197 B.n14 VSUBS 0.009997f
C198 B.n15 VSUBS 0.009997f
C199 B.n16 VSUBS 0.009997f
C200 B.n17 VSUBS 0.009997f
C201 B.n18 VSUBS 0.009997f
C202 B.n19 VSUBS 0.009997f
C203 B.n20 VSUBS 0.009997f
C204 B.n21 VSUBS 0.009997f
C205 B.n22 VSUBS 0.009997f
C206 B.n23 VSUBS 0.009997f
C207 B.n24 VSUBS 0.009997f
C208 B.n25 VSUBS 0.009997f
C209 B.n26 VSUBS 0.009997f
C210 B.n27 VSUBS 0.009997f
C211 B.n28 VSUBS 0.02211f
C212 B.n29 VSUBS 0.009997f
C213 B.n30 VSUBS 0.009997f
C214 B.n31 VSUBS 0.009997f
C215 B.n32 VSUBS 0.009997f
C216 B.n33 VSUBS 0.009997f
C217 B.n34 VSUBS 0.009997f
C218 B.n35 VSUBS 0.009997f
C219 B.n36 VSUBS 0.009997f
C220 B.n37 VSUBS 0.009997f
C221 B.n38 VSUBS 0.009997f
C222 B.n39 VSUBS 0.009997f
C223 B.n40 VSUBS 0.009997f
C224 B.n41 VSUBS 0.009997f
C225 B.n42 VSUBS 0.009997f
C226 B.n43 VSUBS 0.009997f
C227 B.t4 VSUBS 0.179185f
C228 B.t5 VSUBS 0.23132f
C229 B.t3 VSUBS 1.89131f
C230 B.n44 VSUBS 0.377745f
C231 B.n45 VSUBS 0.277766f
C232 B.n46 VSUBS 0.009997f
C233 B.n47 VSUBS 0.009997f
C234 B.n48 VSUBS 0.009997f
C235 B.n49 VSUBS 0.009997f
C236 B.t10 VSUBS 0.179188f
C237 B.t11 VSUBS 0.231323f
C238 B.t9 VSUBS 1.89144f
C239 B.n50 VSUBS 0.377609f
C240 B.n51 VSUBS 0.277762f
C241 B.n52 VSUBS 0.023162f
C242 B.n53 VSUBS 0.009997f
C243 B.n54 VSUBS 0.009997f
C244 B.n55 VSUBS 0.009997f
C245 B.n56 VSUBS 0.009997f
C246 B.n57 VSUBS 0.009997f
C247 B.n58 VSUBS 0.009997f
C248 B.n59 VSUBS 0.009997f
C249 B.n60 VSUBS 0.009997f
C250 B.n61 VSUBS 0.009997f
C251 B.n62 VSUBS 0.009997f
C252 B.n63 VSUBS 0.009997f
C253 B.n64 VSUBS 0.009997f
C254 B.n65 VSUBS 0.009997f
C255 B.n66 VSUBS 0.009997f
C256 B.n67 VSUBS 0.02317f
C257 B.n68 VSUBS 0.009997f
C258 B.n69 VSUBS 0.009997f
C259 B.n70 VSUBS 0.009997f
C260 B.n71 VSUBS 0.009997f
C261 B.n72 VSUBS 0.009997f
C262 B.n73 VSUBS 0.009997f
C263 B.n74 VSUBS 0.009997f
C264 B.n75 VSUBS 0.009997f
C265 B.n76 VSUBS 0.009997f
C266 B.n77 VSUBS 0.009997f
C267 B.n78 VSUBS 0.009997f
C268 B.n79 VSUBS 0.009997f
C269 B.n80 VSUBS 0.009997f
C270 B.n81 VSUBS 0.009997f
C271 B.n82 VSUBS 0.009997f
C272 B.n83 VSUBS 0.009997f
C273 B.n84 VSUBS 0.009997f
C274 B.n85 VSUBS 0.009997f
C275 B.n86 VSUBS 0.009997f
C276 B.n87 VSUBS 0.009997f
C277 B.n88 VSUBS 0.009997f
C278 B.n89 VSUBS 0.009997f
C279 B.n90 VSUBS 0.009997f
C280 B.n91 VSUBS 0.009997f
C281 B.n92 VSUBS 0.009997f
C282 B.n93 VSUBS 0.009997f
C283 B.n94 VSUBS 0.009997f
C284 B.n95 VSUBS 0.009997f
C285 B.n96 VSUBS 0.009997f
C286 B.n97 VSUBS 0.009997f
C287 B.n98 VSUBS 0.009997f
C288 B.n99 VSUBS 0.009997f
C289 B.n100 VSUBS 0.009997f
C290 B.n101 VSUBS 0.009997f
C291 B.n102 VSUBS 0.009997f
C292 B.n103 VSUBS 0.009997f
C293 B.n104 VSUBS 0.009997f
C294 B.n105 VSUBS 0.009997f
C295 B.n106 VSUBS 0.009997f
C296 B.n107 VSUBS 0.009997f
C297 B.n108 VSUBS 0.009997f
C298 B.n109 VSUBS 0.009997f
C299 B.n110 VSUBS 0.009997f
C300 B.n111 VSUBS 0.009997f
C301 B.n112 VSUBS 0.009997f
C302 B.n113 VSUBS 0.009997f
C303 B.n114 VSUBS 0.009997f
C304 B.n115 VSUBS 0.009997f
C305 B.n116 VSUBS 0.009997f
C306 B.n117 VSUBS 0.009997f
C307 B.n118 VSUBS 0.009997f
C308 B.n119 VSUBS 0.009997f
C309 B.n120 VSUBS 0.009997f
C310 B.n121 VSUBS 0.02211f
C311 B.n122 VSUBS 0.009997f
C312 B.n123 VSUBS 0.009997f
C313 B.n124 VSUBS 0.009997f
C314 B.n125 VSUBS 0.009997f
C315 B.n126 VSUBS 0.009997f
C316 B.n127 VSUBS 0.009997f
C317 B.n128 VSUBS 0.009997f
C318 B.n129 VSUBS 0.009997f
C319 B.n130 VSUBS 0.009997f
C320 B.n131 VSUBS 0.009997f
C321 B.n132 VSUBS 0.009997f
C322 B.n133 VSUBS 0.009997f
C323 B.n134 VSUBS 0.009997f
C324 B.n135 VSUBS 0.009997f
C325 B.n136 VSUBS 0.006983f
C326 B.n137 VSUBS 0.009997f
C327 B.n138 VSUBS 0.009997f
C328 B.n139 VSUBS 0.009997f
C329 B.n140 VSUBS 0.009997f
C330 B.n141 VSUBS 0.009997f
C331 B.t2 VSUBS 0.179185f
C332 B.t1 VSUBS 0.23132f
C333 B.t0 VSUBS 1.89131f
C334 B.n142 VSUBS 0.377745f
C335 B.n143 VSUBS 0.277766f
C336 B.n144 VSUBS 0.009997f
C337 B.n145 VSUBS 0.009997f
C338 B.n146 VSUBS 0.009997f
C339 B.n147 VSUBS 0.009997f
C340 B.n148 VSUBS 0.009997f
C341 B.n149 VSUBS 0.009997f
C342 B.n150 VSUBS 0.009997f
C343 B.n151 VSUBS 0.009997f
C344 B.n152 VSUBS 0.009997f
C345 B.n153 VSUBS 0.009997f
C346 B.n154 VSUBS 0.009997f
C347 B.n155 VSUBS 0.009997f
C348 B.n156 VSUBS 0.009997f
C349 B.n157 VSUBS 0.009997f
C350 B.n158 VSUBS 0.02211f
C351 B.n159 VSUBS 0.009997f
C352 B.n160 VSUBS 0.009997f
C353 B.n161 VSUBS 0.009997f
C354 B.n162 VSUBS 0.009997f
C355 B.n163 VSUBS 0.009997f
C356 B.n164 VSUBS 0.009997f
C357 B.n165 VSUBS 0.009997f
C358 B.n166 VSUBS 0.009997f
C359 B.n167 VSUBS 0.009997f
C360 B.n168 VSUBS 0.009997f
C361 B.n169 VSUBS 0.009997f
C362 B.n170 VSUBS 0.009997f
C363 B.n171 VSUBS 0.009997f
C364 B.n172 VSUBS 0.009997f
C365 B.n173 VSUBS 0.009997f
C366 B.n174 VSUBS 0.009997f
C367 B.n175 VSUBS 0.009997f
C368 B.n176 VSUBS 0.009997f
C369 B.n177 VSUBS 0.009997f
C370 B.n178 VSUBS 0.009997f
C371 B.n179 VSUBS 0.009997f
C372 B.n180 VSUBS 0.009997f
C373 B.n181 VSUBS 0.009997f
C374 B.n182 VSUBS 0.009997f
C375 B.n183 VSUBS 0.009997f
C376 B.n184 VSUBS 0.009997f
C377 B.n185 VSUBS 0.009997f
C378 B.n186 VSUBS 0.009997f
C379 B.n187 VSUBS 0.009997f
C380 B.n188 VSUBS 0.009997f
C381 B.n189 VSUBS 0.009997f
C382 B.n190 VSUBS 0.009997f
C383 B.n191 VSUBS 0.009997f
C384 B.n192 VSUBS 0.009997f
C385 B.n193 VSUBS 0.009997f
C386 B.n194 VSUBS 0.009997f
C387 B.n195 VSUBS 0.009997f
C388 B.n196 VSUBS 0.009997f
C389 B.n197 VSUBS 0.009997f
C390 B.n198 VSUBS 0.009997f
C391 B.n199 VSUBS 0.009997f
C392 B.n200 VSUBS 0.009997f
C393 B.n201 VSUBS 0.009997f
C394 B.n202 VSUBS 0.009997f
C395 B.n203 VSUBS 0.009997f
C396 B.n204 VSUBS 0.009997f
C397 B.n205 VSUBS 0.009997f
C398 B.n206 VSUBS 0.009997f
C399 B.n207 VSUBS 0.009997f
C400 B.n208 VSUBS 0.009997f
C401 B.n209 VSUBS 0.009997f
C402 B.n210 VSUBS 0.009997f
C403 B.n211 VSUBS 0.009997f
C404 B.n212 VSUBS 0.009997f
C405 B.n213 VSUBS 0.009997f
C406 B.n214 VSUBS 0.009997f
C407 B.n215 VSUBS 0.009997f
C408 B.n216 VSUBS 0.009997f
C409 B.n217 VSUBS 0.009997f
C410 B.n218 VSUBS 0.009997f
C411 B.n219 VSUBS 0.009997f
C412 B.n220 VSUBS 0.009997f
C413 B.n221 VSUBS 0.009997f
C414 B.n222 VSUBS 0.009997f
C415 B.n223 VSUBS 0.009997f
C416 B.n224 VSUBS 0.009997f
C417 B.n225 VSUBS 0.009997f
C418 B.n226 VSUBS 0.009997f
C419 B.n227 VSUBS 0.009997f
C420 B.n228 VSUBS 0.009997f
C421 B.n229 VSUBS 0.009997f
C422 B.n230 VSUBS 0.009997f
C423 B.n231 VSUBS 0.009997f
C424 B.n232 VSUBS 0.009997f
C425 B.n233 VSUBS 0.009997f
C426 B.n234 VSUBS 0.009997f
C427 B.n235 VSUBS 0.009997f
C428 B.n236 VSUBS 0.009997f
C429 B.n237 VSUBS 0.009997f
C430 B.n238 VSUBS 0.009997f
C431 B.n239 VSUBS 0.009997f
C432 B.n240 VSUBS 0.009997f
C433 B.n241 VSUBS 0.009997f
C434 B.n242 VSUBS 0.009997f
C435 B.n243 VSUBS 0.009997f
C436 B.n244 VSUBS 0.009997f
C437 B.n245 VSUBS 0.009997f
C438 B.n246 VSUBS 0.009997f
C439 B.n247 VSUBS 0.009997f
C440 B.n248 VSUBS 0.009997f
C441 B.n249 VSUBS 0.009997f
C442 B.n250 VSUBS 0.009997f
C443 B.n251 VSUBS 0.009997f
C444 B.n252 VSUBS 0.009997f
C445 B.n253 VSUBS 0.009997f
C446 B.n254 VSUBS 0.009997f
C447 B.n255 VSUBS 0.009997f
C448 B.n256 VSUBS 0.009997f
C449 B.n257 VSUBS 0.009997f
C450 B.n258 VSUBS 0.009997f
C451 B.n259 VSUBS 0.009997f
C452 B.n260 VSUBS 0.009997f
C453 B.n261 VSUBS 0.02211f
C454 B.n262 VSUBS 0.02317f
C455 B.n263 VSUBS 0.02317f
C456 B.n264 VSUBS 0.009997f
C457 B.n265 VSUBS 0.009997f
C458 B.n266 VSUBS 0.009997f
C459 B.n267 VSUBS 0.009997f
C460 B.n268 VSUBS 0.009997f
C461 B.n269 VSUBS 0.009997f
C462 B.n270 VSUBS 0.009997f
C463 B.n271 VSUBS 0.009997f
C464 B.n272 VSUBS 0.009997f
C465 B.n273 VSUBS 0.009997f
C466 B.n274 VSUBS 0.009997f
C467 B.n275 VSUBS 0.009997f
C468 B.n276 VSUBS 0.009997f
C469 B.n277 VSUBS 0.009997f
C470 B.n278 VSUBS 0.009997f
C471 B.n279 VSUBS 0.009997f
C472 B.n280 VSUBS 0.009997f
C473 B.n281 VSUBS 0.009997f
C474 B.n282 VSUBS 0.009997f
C475 B.n283 VSUBS 0.009997f
C476 B.n284 VSUBS 0.009997f
C477 B.n285 VSUBS 0.009997f
C478 B.n286 VSUBS 0.009997f
C479 B.n287 VSUBS 0.009997f
C480 B.n288 VSUBS 0.009997f
C481 B.n289 VSUBS 0.009997f
C482 B.n290 VSUBS 0.009997f
C483 B.n291 VSUBS 0.009997f
C484 B.n292 VSUBS 0.009997f
C485 B.n293 VSUBS 0.009997f
C486 B.n294 VSUBS 0.009997f
C487 B.n295 VSUBS 0.009997f
C488 B.n296 VSUBS 0.009997f
C489 B.n297 VSUBS 0.009997f
C490 B.n298 VSUBS 0.009997f
C491 B.n299 VSUBS 0.009997f
C492 B.n300 VSUBS 0.009997f
C493 B.n301 VSUBS 0.009997f
C494 B.n302 VSUBS 0.009997f
C495 B.n303 VSUBS 0.009997f
C496 B.n304 VSUBS 0.009997f
C497 B.n305 VSUBS 0.009997f
C498 B.n306 VSUBS 0.006983f
C499 B.n307 VSUBS 0.023162f
C500 B.n308 VSUBS 0.008012f
C501 B.n309 VSUBS 0.009997f
C502 B.n310 VSUBS 0.009997f
C503 B.n311 VSUBS 0.009997f
C504 B.n312 VSUBS 0.009997f
C505 B.n313 VSUBS 0.009997f
C506 B.n314 VSUBS 0.009997f
C507 B.n315 VSUBS 0.009997f
C508 B.n316 VSUBS 0.009997f
C509 B.n317 VSUBS 0.009997f
C510 B.n318 VSUBS 0.009997f
C511 B.n319 VSUBS 0.009997f
C512 B.t8 VSUBS 0.179188f
C513 B.t7 VSUBS 0.231323f
C514 B.t6 VSUBS 1.89144f
C515 B.n320 VSUBS 0.377609f
C516 B.n321 VSUBS 0.277762f
C517 B.n322 VSUBS 0.023162f
C518 B.n323 VSUBS 0.008012f
C519 B.n324 VSUBS 0.009997f
C520 B.n325 VSUBS 0.009997f
C521 B.n326 VSUBS 0.009997f
C522 B.n327 VSUBS 0.009997f
C523 B.n328 VSUBS 0.009997f
C524 B.n329 VSUBS 0.009997f
C525 B.n330 VSUBS 0.009997f
C526 B.n331 VSUBS 0.009997f
C527 B.n332 VSUBS 0.009997f
C528 B.n333 VSUBS 0.009997f
C529 B.n334 VSUBS 0.009997f
C530 B.n335 VSUBS 0.009997f
C531 B.n336 VSUBS 0.009997f
C532 B.n337 VSUBS 0.009997f
C533 B.n338 VSUBS 0.009997f
C534 B.n339 VSUBS 0.009997f
C535 B.n340 VSUBS 0.009997f
C536 B.n341 VSUBS 0.009997f
C537 B.n342 VSUBS 0.009997f
C538 B.n343 VSUBS 0.009997f
C539 B.n344 VSUBS 0.009997f
C540 B.n345 VSUBS 0.009997f
C541 B.n346 VSUBS 0.009997f
C542 B.n347 VSUBS 0.009997f
C543 B.n348 VSUBS 0.009997f
C544 B.n349 VSUBS 0.009997f
C545 B.n350 VSUBS 0.009997f
C546 B.n351 VSUBS 0.009997f
C547 B.n352 VSUBS 0.009997f
C548 B.n353 VSUBS 0.009997f
C549 B.n354 VSUBS 0.009997f
C550 B.n355 VSUBS 0.009997f
C551 B.n356 VSUBS 0.009997f
C552 B.n357 VSUBS 0.009997f
C553 B.n358 VSUBS 0.009997f
C554 B.n359 VSUBS 0.009997f
C555 B.n360 VSUBS 0.009997f
C556 B.n361 VSUBS 0.009997f
C557 B.n362 VSUBS 0.009997f
C558 B.n363 VSUBS 0.009997f
C559 B.n364 VSUBS 0.009997f
C560 B.n365 VSUBS 0.009997f
C561 B.n366 VSUBS 0.009997f
C562 B.n367 VSUBS 0.009997f
C563 B.n368 VSUBS 0.02317f
C564 B.n369 VSUBS 0.021928f
C565 B.n370 VSUBS 0.023352f
C566 B.n371 VSUBS 0.009997f
C567 B.n372 VSUBS 0.009997f
C568 B.n373 VSUBS 0.009997f
C569 B.n374 VSUBS 0.009997f
C570 B.n375 VSUBS 0.009997f
C571 B.n376 VSUBS 0.009997f
C572 B.n377 VSUBS 0.009997f
C573 B.n378 VSUBS 0.009997f
C574 B.n379 VSUBS 0.009997f
C575 B.n380 VSUBS 0.009997f
C576 B.n381 VSUBS 0.009997f
C577 B.n382 VSUBS 0.009997f
C578 B.n383 VSUBS 0.009997f
C579 B.n384 VSUBS 0.009997f
C580 B.n385 VSUBS 0.009997f
C581 B.n386 VSUBS 0.009997f
C582 B.n387 VSUBS 0.009997f
C583 B.n388 VSUBS 0.009997f
C584 B.n389 VSUBS 0.009997f
C585 B.n390 VSUBS 0.009997f
C586 B.n391 VSUBS 0.009997f
C587 B.n392 VSUBS 0.009997f
C588 B.n393 VSUBS 0.009997f
C589 B.n394 VSUBS 0.009997f
C590 B.n395 VSUBS 0.009997f
C591 B.n396 VSUBS 0.009997f
C592 B.n397 VSUBS 0.009997f
C593 B.n398 VSUBS 0.009997f
C594 B.n399 VSUBS 0.009997f
C595 B.n400 VSUBS 0.009997f
C596 B.n401 VSUBS 0.009997f
C597 B.n402 VSUBS 0.009997f
C598 B.n403 VSUBS 0.009997f
C599 B.n404 VSUBS 0.009997f
C600 B.n405 VSUBS 0.009997f
C601 B.n406 VSUBS 0.009997f
C602 B.n407 VSUBS 0.009997f
C603 B.n408 VSUBS 0.009997f
C604 B.n409 VSUBS 0.009997f
C605 B.n410 VSUBS 0.009997f
C606 B.n411 VSUBS 0.009997f
C607 B.n412 VSUBS 0.009997f
C608 B.n413 VSUBS 0.009997f
C609 B.n414 VSUBS 0.009997f
C610 B.n415 VSUBS 0.009997f
C611 B.n416 VSUBS 0.009997f
C612 B.n417 VSUBS 0.009997f
C613 B.n418 VSUBS 0.009997f
C614 B.n419 VSUBS 0.009997f
C615 B.n420 VSUBS 0.009997f
C616 B.n421 VSUBS 0.009997f
C617 B.n422 VSUBS 0.009997f
C618 B.n423 VSUBS 0.009997f
C619 B.n424 VSUBS 0.009997f
C620 B.n425 VSUBS 0.009997f
C621 B.n426 VSUBS 0.009997f
C622 B.n427 VSUBS 0.009997f
C623 B.n428 VSUBS 0.009997f
C624 B.n429 VSUBS 0.009997f
C625 B.n430 VSUBS 0.009997f
C626 B.n431 VSUBS 0.009997f
C627 B.n432 VSUBS 0.009997f
C628 B.n433 VSUBS 0.009997f
C629 B.n434 VSUBS 0.009997f
C630 B.n435 VSUBS 0.009997f
C631 B.n436 VSUBS 0.009997f
C632 B.n437 VSUBS 0.009997f
C633 B.n438 VSUBS 0.009997f
C634 B.n439 VSUBS 0.009997f
C635 B.n440 VSUBS 0.009997f
C636 B.n441 VSUBS 0.009997f
C637 B.n442 VSUBS 0.009997f
C638 B.n443 VSUBS 0.009997f
C639 B.n444 VSUBS 0.009997f
C640 B.n445 VSUBS 0.009997f
C641 B.n446 VSUBS 0.009997f
C642 B.n447 VSUBS 0.009997f
C643 B.n448 VSUBS 0.009997f
C644 B.n449 VSUBS 0.009997f
C645 B.n450 VSUBS 0.009997f
C646 B.n451 VSUBS 0.009997f
C647 B.n452 VSUBS 0.009997f
C648 B.n453 VSUBS 0.009997f
C649 B.n454 VSUBS 0.009997f
C650 B.n455 VSUBS 0.009997f
C651 B.n456 VSUBS 0.009997f
C652 B.n457 VSUBS 0.009997f
C653 B.n458 VSUBS 0.009997f
C654 B.n459 VSUBS 0.009997f
C655 B.n460 VSUBS 0.009997f
C656 B.n461 VSUBS 0.009997f
C657 B.n462 VSUBS 0.009997f
C658 B.n463 VSUBS 0.009997f
C659 B.n464 VSUBS 0.009997f
C660 B.n465 VSUBS 0.009997f
C661 B.n466 VSUBS 0.009997f
C662 B.n467 VSUBS 0.009997f
C663 B.n468 VSUBS 0.009997f
C664 B.n469 VSUBS 0.009997f
C665 B.n470 VSUBS 0.009997f
C666 B.n471 VSUBS 0.009997f
C667 B.n472 VSUBS 0.009997f
C668 B.n473 VSUBS 0.009997f
C669 B.n474 VSUBS 0.009997f
C670 B.n475 VSUBS 0.009997f
C671 B.n476 VSUBS 0.009997f
C672 B.n477 VSUBS 0.009997f
C673 B.n478 VSUBS 0.009997f
C674 B.n479 VSUBS 0.009997f
C675 B.n480 VSUBS 0.009997f
C676 B.n481 VSUBS 0.009997f
C677 B.n482 VSUBS 0.009997f
C678 B.n483 VSUBS 0.009997f
C679 B.n484 VSUBS 0.009997f
C680 B.n485 VSUBS 0.009997f
C681 B.n486 VSUBS 0.009997f
C682 B.n487 VSUBS 0.009997f
C683 B.n488 VSUBS 0.009997f
C684 B.n489 VSUBS 0.009997f
C685 B.n490 VSUBS 0.009997f
C686 B.n491 VSUBS 0.009997f
C687 B.n492 VSUBS 0.009997f
C688 B.n493 VSUBS 0.009997f
C689 B.n494 VSUBS 0.009997f
C690 B.n495 VSUBS 0.009997f
C691 B.n496 VSUBS 0.009997f
C692 B.n497 VSUBS 0.009997f
C693 B.n498 VSUBS 0.009997f
C694 B.n499 VSUBS 0.009997f
C695 B.n500 VSUBS 0.009997f
C696 B.n501 VSUBS 0.009997f
C697 B.n502 VSUBS 0.009997f
C698 B.n503 VSUBS 0.009997f
C699 B.n504 VSUBS 0.009997f
C700 B.n505 VSUBS 0.009997f
C701 B.n506 VSUBS 0.009997f
C702 B.n507 VSUBS 0.009997f
C703 B.n508 VSUBS 0.009997f
C704 B.n509 VSUBS 0.009997f
C705 B.n510 VSUBS 0.009997f
C706 B.n511 VSUBS 0.009997f
C707 B.n512 VSUBS 0.009997f
C708 B.n513 VSUBS 0.009997f
C709 B.n514 VSUBS 0.009997f
C710 B.n515 VSUBS 0.009997f
C711 B.n516 VSUBS 0.009997f
C712 B.n517 VSUBS 0.009997f
C713 B.n518 VSUBS 0.009997f
C714 B.n519 VSUBS 0.009997f
C715 B.n520 VSUBS 0.009997f
C716 B.n521 VSUBS 0.009997f
C717 B.n522 VSUBS 0.009997f
C718 B.n523 VSUBS 0.009997f
C719 B.n524 VSUBS 0.009997f
C720 B.n525 VSUBS 0.009997f
C721 B.n526 VSUBS 0.009997f
C722 B.n527 VSUBS 0.009997f
C723 B.n528 VSUBS 0.009997f
C724 B.n529 VSUBS 0.009997f
C725 B.n530 VSUBS 0.02211f
C726 B.n531 VSUBS 0.02211f
C727 B.n532 VSUBS 0.02317f
C728 B.n533 VSUBS 0.009997f
C729 B.n534 VSUBS 0.009997f
C730 B.n535 VSUBS 0.009997f
C731 B.n536 VSUBS 0.009997f
C732 B.n537 VSUBS 0.009997f
C733 B.n538 VSUBS 0.009997f
C734 B.n539 VSUBS 0.009997f
C735 B.n540 VSUBS 0.009997f
C736 B.n541 VSUBS 0.009997f
C737 B.n542 VSUBS 0.009997f
C738 B.n543 VSUBS 0.009997f
C739 B.n544 VSUBS 0.009997f
C740 B.n545 VSUBS 0.009997f
C741 B.n546 VSUBS 0.009997f
C742 B.n547 VSUBS 0.009997f
C743 B.n548 VSUBS 0.009997f
C744 B.n549 VSUBS 0.009997f
C745 B.n550 VSUBS 0.009997f
C746 B.n551 VSUBS 0.009997f
C747 B.n552 VSUBS 0.009997f
C748 B.n553 VSUBS 0.009997f
C749 B.n554 VSUBS 0.009997f
C750 B.n555 VSUBS 0.009997f
C751 B.n556 VSUBS 0.009997f
C752 B.n557 VSUBS 0.009997f
C753 B.n558 VSUBS 0.009997f
C754 B.n559 VSUBS 0.009997f
C755 B.n560 VSUBS 0.009997f
C756 B.n561 VSUBS 0.009997f
C757 B.n562 VSUBS 0.009997f
C758 B.n563 VSUBS 0.009997f
C759 B.n564 VSUBS 0.009997f
C760 B.n565 VSUBS 0.009997f
C761 B.n566 VSUBS 0.009997f
C762 B.n567 VSUBS 0.009997f
C763 B.n568 VSUBS 0.009997f
C764 B.n569 VSUBS 0.009997f
C765 B.n570 VSUBS 0.009997f
C766 B.n571 VSUBS 0.009997f
C767 B.n572 VSUBS 0.009997f
C768 B.n573 VSUBS 0.009997f
C769 B.n574 VSUBS 0.009997f
C770 B.n575 VSUBS 0.006983f
C771 B.n576 VSUBS 0.009997f
C772 B.n577 VSUBS 0.009997f
C773 B.n578 VSUBS 0.008012f
C774 B.n579 VSUBS 0.009997f
C775 B.n580 VSUBS 0.009997f
C776 B.n581 VSUBS 0.009997f
C777 B.n582 VSUBS 0.009997f
C778 B.n583 VSUBS 0.009997f
C779 B.n584 VSUBS 0.009997f
C780 B.n585 VSUBS 0.009997f
C781 B.n586 VSUBS 0.009997f
C782 B.n587 VSUBS 0.009997f
C783 B.n588 VSUBS 0.009997f
C784 B.n589 VSUBS 0.009997f
C785 B.n590 VSUBS 0.008012f
C786 B.n591 VSUBS 0.023162f
C787 B.n592 VSUBS 0.006983f
C788 B.n593 VSUBS 0.009997f
C789 B.n594 VSUBS 0.009997f
C790 B.n595 VSUBS 0.009997f
C791 B.n596 VSUBS 0.009997f
C792 B.n597 VSUBS 0.009997f
C793 B.n598 VSUBS 0.009997f
C794 B.n599 VSUBS 0.009997f
C795 B.n600 VSUBS 0.009997f
C796 B.n601 VSUBS 0.009997f
C797 B.n602 VSUBS 0.009997f
C798 B.n603 VSUBS 0.009997f
C799 B.n604 VSUBS 0.009997f
C800 B.n605 VSUBS 0.009997f
C801 B.n606 VSUBS 0.009997f
C802 B.n607 VSUBS 0.009997f
C803 B.n608 VSUBS 0.009997f
C804 B.n609 VSUBS 0.009997f
C805 B.n610 VSUBS 0.009997f
C806 B.n611 VSUBS 0.009997f
C807 B.n612 VSUBS 0.009997f
C808 B.n613 VSUBS 0.009997f
C809 B.n614 VSUBS 0.009997f
C810 B.n615 VSUBS 0.009997f
C811 B.n616 VSUBS 0.009997f
C812 B.n617 VSUBS 0.009997f
C813 B.n618 VSUBS 0.009997f
C814 B.n619 VSUBS 0.009997f
C815 B.n620 VSUBS 0.009997f
C816 B.n621 VSUBS 0.009997f
C817 B.n622 VSUBS 0.009997f
C818 B.n623 VSUBS 0.009997f
C819 B.n624 VSUBS 0.009997f
C820 B.n625 VSUBS 0.009997f
C821 B.n626 VSUBS 0.009997f
C822 B.n627 VSUBS 0.009997f
C823 B.n628 VSUBS 0.009997f
C824 B.n629 VSUBS 0.009997f
C825 B.n630 VSUBS 0.009997f
C826 B.n631 VSUBS 0.009997f
C827 B.n632 VSUBS 0.009997f
C828 B.n633 VSUBS 0.009997f
C829 B.n634 VSUBS 0.009997f
C830 B.n635 VSUBS 0.02317f
C831 B.n636 VSUBS 0.02317f
C832 B.n637 VSUBS 0.02211f
C833 B.n638 VSUBS 0.009997f
C834 B.n639 VSUBS 0.009997f
C835 B.n640 VSUBS 0.009997f
C836 B.n641 VSUBS 0.009997f
C837 B.n642 VSUBS 0.009997f
C838 B.n643 VSUBS 0.009997f
C839 B.n644 VSUBS 0.009997f
C840 B.n645 VSUBS 0.009997f
C841 B.n646 VSUBS 0.009997f
C842 B.n647 VSUBS 0.009997f
C843 B.n648 VSUBS 0.009997f
C844 B.n649 VSUBS 0.009997f
C845 B.n650 VSUBS 0.009997f
C846 B.n651 VSUBS 0.009997f
C847 B.n652 VSUBS 0.009997f
C848 B.n653 VSUBS 0.009997f
C849 B.n654 VSUBS 0.009997f
C850 B.n655 VSUBS 0.009997f
C851 B.n656 VSUBS 0.009997f
C852 B.n657 VSUBS 0.009997f
C853 B.n658 VSUBS 0.009997f
C854 B.n659 VSUBS 0.009997f
C855 B.n660 VSUBS 0.009997f
C856 B.n661 VSUBS 0.009997f
C857 B.n662 VSUBS 0.009997f
C858 B.n663 VSUBS 0.009997f
C859 B.n664 VSUBS 0.009997f
C860 B.n665 VSUBS 0.009997f
C861 B.n666 VSUBS 0.009997f
C862 B.n667 VSUBS 0.009997f
C863 B.n668 VSUBS 0.009997f
C864 B.n669 VSUBS 0.009997f
C865 B.n670 VSUBS 0.009997f
C866 B.n671 VSUBS 0.009997f
C867 B.n672 VSUBS 0.009997f
C868 B.n673 VSUBS 0.009997f
C869 B.n674 VSUBS 0.009997f
C870 B.n675 VSUBS 0.009997f
C871 B.n676 VSUBS 0.009997f
C872 B.n677 VSUBS 0.009997f
C873 B.n678 VSUBS 0.009997f
C874 B.n679 VSUBS 0.009997f
C875 B.n680 VSUBS 0.009997f
C876 B.n681 VSUBS 0.009997f
C877 B.n682 VSUBS 0.009997f
C878 B.n683 VSUBS 0.009997f
C879 B.n684 VSUBS 0.009997f
C880 B.n685 VSUBS 0.009997f
C881 B.n686 VSUBS 0.009997f
C882 B.n687 VSUBS 0.009997f
C883 B.n688 VSUBS 0.009997f
C884 B.n689 VSUBS 0.009997f
C885 B.n690 VSUBS 0.009997f
C886 B.n691 VSUBS 0.009997f
C887 B.n692 VSUBS 0.009997f
C888 B.n693 VSUBS 0.009997f
C889 B.n694 VSUBS 0.009997f
C890 B.n695 VSUBS 0.009997f
C891 B.n696 VSUBS 0.009997f
C892 B.n697 VSUBS 0.009997f
C893 B.n698 VSUBS 0.009997f
C894 B.n699 VSUBS 0.009997f
C895 B.n700 VSUBS 0.009997f
C896 B.n701 VSUBS 0.009997f
C897 B.n702 VSUBS 0.009997f
C898 B.n703 VSUBS 0.009997f
C899 B.n704 VSUBS 0.009997f
C900 B.n705 VSUBS 0.009997f
C901 B.n706 VSUBS 0.009997f
C902 B.n707 VSUBS 0.009997f
C903 B.n708 VSUBS 0.009997f
C904 B.n709 VSUBS 0.009997f
C905 B.n710 VSUBS 0.009997f
C906 B.n711 VSUBS 0.009997f
C907 B.n712 VSUBS 0.009997f
C908 B.n713 VSUBS 0.009997f
C909 B.n714 VSUBS 0.009997f
C910 B.n715 VSUBS 0.013046f
C911 B.n716 VSUBS 0.013897f
C912 B.n717 VSUBS 0.027635f
C913 VDD2.n0 VSUBS 0.031666f
C914 VDD2.n1 VSUBS 0.030095f
C915 VDD2.n2 VSUBS 0.016647f
C916 VDD2.n3 VSUBS 0.038224f
C917 VDD2.n4 VSUBS 0.017123f
C918 VDD2.n5 VSUBS 0.030095f
C919 VDD2.n6 VSUBS 0.016171f
C920 VDD2.n7 VSUBS 0.038224f
C921 VDD2.n8 VSUBS 0.017123f
C922 VDD2.n9 VSUBS 0.030095f
C923 VDD2.n10 VSUBS 0.016171f
C924 VDD2.n11 VSUBS 0.028668f
C925 VDD2.n12 VSUBS 0.028753f
C926 VDD2.t3 VSUBS 0.082094f
C927 VDD2.n13 VSUBS 0.181882f
C928 VDD2.n14 VSUBS 0.943024f
C929 VDD2.n15 VSUBS 0.016171f
C930 VDD2.n16 VSUBS 0.017123f
C931 VDD2.n17 VSUBS 0.038224f
C932 VDD2.n18 VSUBS 0.038224f
C933 VDD2.n19 VSUBS 0.017123f
C934 VDD2.n20 VSUBS 0.016171f
C935 VDD2.n21 VSUBS 0.030095f
C936 VDD2.n22 VSUBS 0.030095f
C937 VDD2.n23 VSUBS 0.016171f
C938 VDD2.n24 VSUBS 0.017123f
C939 VDD2.n25 VSUBS 0.038224f
C940 VDD2.n26 VSUBS 0.038224f
C941 VDD2.n27 VSUBS 0.017123f
C942 VDD2.n28 VSUBS 0.016171f
C943 VDD2.n29 VSUBS 0.030095f
C944 VDD2.n30 VSUBS 0.030095f
C945 VDD2.n31 VSUBS 0.016171f
C946 VDD2.n32 VSUBS 0.016171f
C947 VDD2.n33 VSUBS 0.017123f
C948 VDD2.n34 VSUBS 0.038224f
C949 VDD2.n35 VSUBS 0.038224f
C950 VDD2.n36 VSUBS 0.087761f
C951 VDD2.n37 VSUBS 0.016647f
C952 VDD2.n38 VSUBS 0.016171f
C953 VDD2.n39 VSUBS 0.075318f
C954 VDD2.n40 VSUBS 0.078239f
C955 VDD2.t4 VSUBS 0.188826f
C956 VDD2.t1 VSUBS 0.188826f
C957 VDD2.n41 VSUBS 1.37487f
C958 VDD2.n42 VSUBS 3.66369f
C959 VDD2.n43 VSUBS 0.031666f
C960 VDD2.n44 VSUBS 0.030095f
C961 VDD2.n45 VSUBS 0.016647f
C962 VDD2.n46 VSUBS 0.038224f
C963 VDD2.n47 VSUBS 0.016171f
C964 VDD2.n48 VSUBS 0.017123f
C965 VDD2.n49 VSUBS 0.030095f
C966 VDD2.n50 VSUBS 0.016171f
C967 VDD2.n51 VSUBS 0.038224f
C968 VDD2.n52 VSUBS 0.017123f
C969 VDD2.n53 VSUBS 0.030095f
C970 VDD2.n54 VSUBS 0.016171f
C971 VDD2.n55 VSUBS 0.028668f
C972 VDD2.n56 VSUBS 0.028753f
C973 VDD2.t5 VSUBS 0.082094f
C974 VDD2.n57 VSUBS 0.181882f
C975 VDD2.n58 VSUBS 0.943024f
C976 VDD2.n59 VSUBS 0.016171f
C977 VDD2.n60 VSUBS 0.017123f
C978 VDD2.n61 VSUBS 0.038224f
C979 VDD2.n62 VSUBS 0.038224f
C980 VDD2.n63 VSUBS 0.017123f
C981 VDD2.n64 VSUBS 0.016171f
C982 VDD2.n65 VSUBS 0.030095f
C983 VDD2.n66 VSUBS 0.030095f
C984 VDD2.n67 VSUBS 0.016171f
C985 VDD2.n68 VSUBS 0.017123f
C986 VDD2.n69 VSUBS 0.038224f
C987 VDD2.n70 VSUBS 0.038224f
C988 VDD2.n71 VSUBS 0.017123f
C989 VDD2.n72 VSUBS 0.016171f
C990 VDD2.n73 VSUBS 0.030095f
C991 VDD2.n74 VSUBS 0.030095f
C992 VDD2.n75 VSUBS 0.016171f
C993 VDD2.n76 VSUBS 0.017123f
C994 VDD2.n77 VSUBS 0.038224f
C995 VDD2.n78 VSUBS 0.038224f
C996 VDD2.n79 VSUBS 0.087761f
C997 VDD2.n80 VSUBS 0.016647f
C998 VDD2.n81 VSUBS 0.016171f
C999 VDD2.n82 VSUBS 0.075318f
C1000 VDD2.n83 VSUBS 0.064831f
C1001 VDD2.n84 VSUBS 3.01052f
C1002 VDD2.t0 VSUBS 0.188826f
C1003 VDD2.t2 VSUBS 0.188826f
C1004 VDD2.n85 VSUBS 1.37483f
C1005 VTAIL.t8 VSUBS 0.202714f
C1006 VTAIL.t7 VSUBS 0.202714f
C1007 VTAIL.n0 VSUBS 1.33596f
C1008 VTAIL.n1 VSUBS 0.945299f
C1009 VTAIL.n2 VSUBS 0.033995f
C1010 VTAIL.n3 VSUBS 0.032308f
C1011 VTAIL.n4 VSUBS 0.017872f
C1012 VTAIL.n5 VSUBS 0.041035f
C1013 VTAIL.n6 VSUBS 0.018382f
C1014 VTAIL.n7 VSUBS 0.032308f
C1015 VTAIL.n8 VSUBS 0.017361f
C1016 VTAIL.n9 VSUBS 0.041035f
C1017 VTAIL.n10 VSUBS 0.018382f
C1018 VTAIL.n11 VSUBS 0.032308f
C1019 VTAIL.n12 VSUBS 0.017361f
C1020 VTAIL.n13 VSUBS 0.030776f
C1021 VTAIL.n14 VSUBS 0.030868f
C1022 VTAIL.t4 VSUBS 0.088132f
C1023 VTAIL.n15 VSUBS 0.195259f
C1024 VTAIL.n16 VSUBS 1.01238f
C1025 VTAIL.n17 VSUBS 0.017361f
C1026 VTAIL.n18 VSUBS 0.018382f
C1027 VTAIL.n19 VSUBS 0.041035f
C1028 VTAIL.n20 VSUBS 0.041035f
C1029 VTAIL.n21 VSUBS 0.018382f
C1030 VTAIL.n22 VSUBS 0.017361f
C1031 VTAIL.n23 VSUBS 0.032308f
C1032 VTAIL.n24 VSUBS 0.032308f
C1033 VTAIL.n25 VSUBS 0.017361f
C1034 VTAIL.n26 VSUBS 0.018382f
C1035 VTAIL.n27 VSUBS 0.041035f
C1036 VTAIL.n28 VSUBS 0.041035f
C1037 VTAIL.n29 VSUBS 0.018382f
C1038 VTAIL.n30 VSUBS 0.017361f
C1039 VTAIL.n31 VSUBS 0.032308f
C1040 VTAIL.n32 VSUBS 0.032308f
C1041 VTAIL.n33 VSUBS 0.017361f
C1042 VTAIL.n34 VSUBS 0.017361f
C1043 VTAIL.n35 VSUBS 0.018382f
C1044 VTAIL.n36 VSUBS 0.041035f
C1045 VTAIL.n37 VSUBS 0.041035f
C1046 VTAIL.n38 VSUBS 0.094216f
C1047 VTAIL.n39 VSUBS 0.017872f
C1048 VTAIL.n40 VSUBS 0.017361f
C1049 VTAIL.n41 VSUBS 0.080857f
C1050 VTAIL.n42 VSUBS 0.047336f
C1051 VTAIL.n43 VSUBS 0.598272f
C1052 VTAIL.t1 VSUBS 0.202714f
C1053 VTAIL.t2 VSUBS 0.202714f
C1054 VTAIL.n44 VSUBS 1.33596f
C1055 VTAIL.n45 VSUBS 2.81918f
C1056 VTAIL.t11 VSUBS 0.202714f
C1057 VTAIL.t10 VSUBS 0.202714f
C1058 VTAIL.n46 VSUBS 1.33597f
C1059 VTAIL.n47 VSUBS 2.81917f
C1060 VTAIL.n48 VSUBS 0.033995f
C1061 VTAIL.n49 VSUBS 0.032308f
C1062 VTAIL.n50 VSUBS 0.017872f
C1063 VTAIL.n51 VSUBS 0.041035f
C1064 VTAIL.n52 VSUBS 0.017361f
C1065 VTAIL.n53 VSUBS 0.018382f
C1066 VTAIL.n54 VSUBS 0.032308f
C1067 VTAIL.n55 VSUBS 0.017361f
C1068 VTAIL.n56 VSUBS 0.041035f
C1069 VTAIL.n57 VSUBS 0.018382f
C1070 VTAIL.n58 VSUBS 0.032308f
C1071 VTAIL.n59 VSUBS 0.017361f
C1072 VTAIL.n60 VSUBS 0.030776f
C1073 VTAIL.n61 VSUBS 0.030868f
C1074 VTAIL.t9 VSUBS 0.088132f
C1075 VTAIL.n62 VSUBS 0.195259f
C1076 VTAIL.n63 VSUBS 1.01238f
C1077 VTAIL.n64 VSUBS 0.017361f
C1078 VTAIL.n65 VSUBS 0.018382f
C1079 VTAIL.n66 VSUBS 0.041035f
C1080 VTAIL.n67 VSUBS 0.041035f
C1081 VTAIL.n68 VSUBS 0.018382f
C1082 VTAIL.n69 VSUBS 0.017361f
C1083 VTAIL.n70 VSUBS 0.032308f
C1084 VTAIL.n71 VSUBS 0.032308f
C1085 VTAIL.n72 VSUBS 0.017361f
C1086 VTAIL.n73 VSUBS 0.018382f
C1087 VTAIL.n74 VSUBS 0.041035f
C1088 VTAIL.n75 VSUBS 0.041035f
C1089 VTAIL.n76 VSUBS 0.018382f
C1090 VTAIL.n77 VSUBS 0.017361f
C1091 VTAIL.n78 VSUBS 0.032308f
C1092 VTAIL.n79 VSUBS 0.032308f
C1093 VTAIL.n80 VSUBS 0.017361f
C1094 VTAIL.n81 VSUBS 0.018382f
C1095 VTAIL.n82 VSUBS 0.041035f
C1096 VTAIL.n83 VSUBS 0.041035f
C1097 VTAIL.n84 VSUBS 0.094216f
C1098 VTAIL.n85 VSUBS 0.017872f
C1099 VTAIL.n86 VSUBS 0.017361f
C1100 VTAIL.n87 VSUBS 0.080857f
C1101 VTAIL.n88 VSUBS 0.047336f
C1102 VTAIL.n89 VSUBS 0.598272f
C1103 VTAIL.t3 VSUBS 0.202714f
C1104 VTAIL.t0 VSUBS 0.202714f
C1105 VTAIL.n90 VSUBS 1.33597f
C1106 VTAIL.n91 VSUBS 1.19837f
C1107 VTAIL.n92 VSUBS 0.033995f
C1108 VTAIL.n93 VSUBS 0.032308f
C1109 VTAIL.n94 VSUBS 0.017872f
C1110 VTAIL.n95 VSUBS 0.041035f
C1111 VTAIL.n96 VSUBS 0.017361f
C1112 VTAIL.n97 VSUBS 0.018382f
C1113 VTAIL.n98 VSUBS 0.032308f
C1114 VTAIL.n99 VSUBS 0.017361f
C1115 VTAIL.n100 VSUBS 0.041035f
C1116 VTAIL.n101 VSUBS 0.018382f
C1117 VTAIL.n102 VSUBS 0.032308f
C1118 VTAIL.n103 VSUBS 0.017361f
C1119 VTAIL.n104 VSUBS 0.030776f
C1120 VTAIL.n105 VSUBS 0.030868f
C1121 VTAIL.t5 VSUBS 0.088132f
C1122 VTAIL.n106 VSUBS 0.195259f
C1123 VTAIL.n107 VSUBS 1.01238f
C1124 VTAIL.n108 VSUBS 0.017361f
C1125 VTAIL.n109 VSUBS 0.018382f
C1126 VTAIL.n110 VSUBS 0.041035f
C1127 VTAIL.n111 VSUBS 0.041035f
C1128 VTAIL.n112 VSUBS 0.018382f
C1129 VTAIL.n113 VSUBS 0.017361f
C1130 VTAIL.n114 VSUBS 0.032308f
C1131 VTAIL.n115 VSUBS 0.032308f
C1132 VTAIL.n116 VSUBS 0.017361f
C1133 VTAIL.n117 VSUBS 0.018382f
C1134 VTAIL.n118 VSUBS 0.041035f
C1135 VTAIL.n119 VSUBS 0.041035f
C1136 VTAIL.n120 VSUBS 0.018382f
C1137 VTAIL.n121 VSUBS 0.017361f
C1138 VTAIL.n122 VSUBS 0.032308f
C1139 VTAIL.n123 VSUBS 0.032308f
C1140 VTAIL.n124 VSUBS 0.017361f
C1141 VTAIL.n125 VSUBS 0.018382f
C1142 VTAIL.n126 VSUBS 0.041035f
C1143 VTAIL.n127 VSUBS 0.041035f
C1144 VTAIL.n128 VSUBS 0.094216f
C1145 VTAIL.n129 VSUBS 0.017872f
C1146 VTAIL.n130 VSUBS 0.017361f
C1147 VTAIL.n131 VSUBS 0.080857f
C1148 VTAIL.n132 VSUBS 0.047336f
C1149 VTAIL.n133 VSUBS 1.87356f
C1150 VTAIL.n134 VSUBS 0.033995f
C1151 VTAIL.n135 VSUBS 0.032308f
C1152 VTAIL.n136 VSUBS 0.017872f
C1153 VTAIL.n137 VSUBS 0.041035f
C1154 VTAIL.n138 VSUBS 0.018382f
C1155 VTAIL.n139 VSUBS 0.032308f
C1156 VTAIL.n140 VSUBS 0.017361f
C1157 VTAIL.n141 VSUBS 0.041035f
C1158 VTAIL.n142 VSUBS 0.018382f
C1159 VTAIL.n143 VSUBS 0.032308f
C1160 VTAIL.n144 VSUBS 0.017361f
C1161 VTAIL.n145 VSUBS 0.030776f
C1162 VTAIL.n146 VSUBS 0.030868f
C1163 VTAIL.t6 VSUBS 0.088132f
C1164 VTAIL.n147 VSUBS 0.195259f
C1165 VTAIL.n148 VSUBS 1.01238f
C1166 VTAIL.n149 VSUBS 0.017361f
C1167 VTAIL.n150 VSUBS 0.018382f
C1168 VTAIL.n151 VSUBS 0.041035f
C1169 VTAIL.n152 VSUBS 0.041035f
C1170 VTAIL.n153 VSUBS 0.018382f
C1171 VTAIL.n154 VSUBS 0.017361f
C1172 VTAIL.n155 VSUBS 0.032308f
C1173 VTAIL.n156 VSUBS 0.032308f
C1174 VTAIL.n157 VSUBS 0.017361f
C1175 VTAIL.n158 VSUBS 0.018382f
C1176 VTAIL.n159 VSUBS 0.041035f
C1177 VTAIL.n160 VSUBS 0.041035f
C1178 VTAIL.n161 VSUBS 0.018382f
C1179 VTAIL.n162 VSUBS 0.017361f
C1180 VTAIL.n163 VSUBS 0.032308f
C1181 VTAIL.n164 VSUBS 0.032308f
C1182 VTAIL.n165 VSUBS 0.017361f
C1183 VTAIL.n166 VSUBS 0.017361f
C1184 VTAIL.n167 VSUBS 0.018382f
C1185 VTAIL.n168 VSUBS 0.041035f
C1186 VTAIL.n169 VSUBS 0.041035f
C1187 VTAIL.n170 VSUBS 0.094216f
C1188 VTAIL.n171 VSUBS 0.017872f
C1189 VTAIL.n172 VSUBS 0.017361f
C1190 VTAIL.n173 VSUBS 0.080857f
C1191 VTAIL.n174 VSUBS 0.047336f
C1192 VTAIL.n175 VSUBS 1.78112f
C1193 VN.t4 VSUBS 2.24969f
C1194 VN.n0 VSUBS 0.919784f
C1195 VN.n1 VSUBS 0.030007f
C1196 VN.n2 VSUBS 0.050311f
C1197 VN.n3 VSUBS 0.030007f
C1198 VN.n4 VSUBS 0.042331f
C1199 VN.t1 VSUBS 2.24969f
C1200 VN.n5 VSUBS 0.914982f
C1201 VN.t2 VSUBS 2.63591f
C1202 VN.n6 VSUBS 0.875862f
C1203 VN.n7 VSUBS 0.373911f
C1204 VN.n8 VSUBS 0.030007f
C1205 VN.n9 VSUBS 0.056206f
C1206 VN.n10 VSUBS 0.056206f
C1207 VN.n11 VSUBS 0.03768f
C1208 VN.n12 VSUBS 0.030007f
C1209 VN.n13 VSUBS 0.030007f
C1210 VN.n14 VSUBS 0.030007f
C1211 VN.n15 VSUBS 0.056206f
C1212 VN.n16 VSUBS 0.056206f
C1213 VN.n17 VSUBS 0.034005f
C1214 VN.n18 VSUBS 0.048439f
C1215 VN.n19 VSUBS 0.085938f
C1216 VN.t0 VSUBS 2.24969f
C1217 VN.n20 VSUBS 0.919784f
C1218 VN.n21 VSUBS 0.030007f
C1219 VN.n22 VSUBS 0.050311f
C1220 VN.n23 VSUBS 0.030007f
C1221 VN.n24 VSUBS 0.042331f
C1222 VN.t3 VSUBS 2.63591f
C1223 VN.t5 VSUBS 2.24969f
C1224 VN.n25 VSUBS 0.914982f
C1225 VN.n26 VSUBS 0.875862f
C1226 VN.n27 VSUBS 0.373911f
C1227 VN.n28 VSUBS 0.030007f
C1228 VN.n29 VSUBS 0.056206f
C1229 VN.n30 VSUBS 0.056206f
C1230 VN.n31 VSUBS 0.03768f
C1231 VN.n32 VSUBS 0.030007f
C1232 VN.n33 VSUBS 0.030007f
C1233 VN.n34 VSUBS 0.030007f
C1234 VN.n35 VSUBS 0.056206f
C1235 VN.n36 VSUBS 0.056206f
C1236 VN.n37 VSUBS 0.034005f
C1237 VN.n38 VSUBS 0.048439f
C1238 VN.n39 VSUBS 1.69289f
.ends

