* NGSPICE file created from diff_pair_sample_0478.ext - technology: sky130A

.subckt diff_pair_sample_0478 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=0.98
X1 VTAIL.t11 VN.t0 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=0.98
X2 VDD1.t4 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=0.98
X3 VDD1.t3 VP.t2 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=0.98
X4 VDD2.t4 VN.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=0.98
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=0.98
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=0.98
X7 VTAIL.t4 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=0.98
X8 VDD2.t3 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=0.98
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=0.98
X10 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=0.98
X11 VTAIL.t2 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=0.98
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=0.98
X13 VDD2.t0 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=0.98
X14 VDD1.t1 VP.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=0.98
X15 VTAIL.t9 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=0.98
R0 VP.n20 VP.n19 161.3
R1 VP.n7 VP.n6 161.3
R2 VP.n8 VP.n3 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n18 VP.n0 161.3
R5 VP.n17 VP.n16 161.3
R6 VP.n15 VP.n14 161.3
R7 VP.n13 VP.n2 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n5 VP.t2 109.773
R10 VP.n12 VP.t1 90.2525
R11 VP.n19 VP.t0 90.2525
R12 VP.n9 VP.t4 90.2525
R13 VP.n1 VP.t5 49.9219
R14 VP.n4 VP.t3 49.9219
R15 VP.n14 VP.n13 49.7204
R16 VP.n18 VP.n17 49.7204
R17 VP.n8 VP.n7 49.7204
R18 VP.n6 VP.n5 43.1531
R19 VP.n5 VP.n4 42.1911
R20 VP.n11 VP.n10 34.8376
R21 VP.n14 VP.n1 12.234
R22 VP.n17 VP.n1 12.234
R23 VP.n7 VP.n4 12.234
R24 VP.n13 VP.n12 10.2247
R25 VP.n19 VP.n18 10.2247
R26 VP.n9 VP.n8 10.2247
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VTAIL.n34 VTAIL.n32 289.615
R36 VTAIL.n4 VTAIL.n2 289.615
R37 VTAIL.n26 VTAIL.n24 289.615
R38 VTAIL.n16 VTAIL.n14 289.615
R39 VTAIL.n35 VTAIL.n34 185
R40 VTAIL.n5 VTAIL.n4 185
R41 VTAIL.n27 VTAIL.n26 185
R42 VTAIL.n17 VTAIL.n16 185
R43 VTAIL.t3 VTAIL.n33 167.117
R44 VTAIL.t8 VTAIL.n3 167.117
R45 VTAIL.t7 VTAIL.n25 167.117
R46 VTAIL.t1 VTAIL.n15 167.117
R47 VTAIL.n23 VTAIL.n22 84.6987
R48 VTAIL.n13 VTAIL.n12 84.6987
R49 VTAIL.n1 VTAIL.n0 84.6986
R50 VTAIL.n11 VTAIL.n10 84.6986
R51 VTAIL.n34 VTAIL.t3 52.3082
R52 VTAIL.n4 VTAIL.t8 52.3082
R53 VTAIL.n26 VTAIL.t7 52.3082
R54 VTAIL.n16 VTAIL.t1 52.3082
R55 VTAIL.n39 VTAIL.n38 31.9914
R56 VTAIL.n9 VTAIL.n8 31.9914
R57 VTAIL.n31 VTAIL.n30 31.9914
R58 VTAIL.n21 VTAIL.n20 31.9914
R59 VTAIL.n13 VTAIL.n11 16.3755
R60 VTAIL.n39 VTAIL.n31 15.2462
R61 VTAIL.n0 VTAIL.t0 9.75419
R62 VTAIL.n0 VTAIL.t2 9.75419
R63 VTAIL.n10 VTAIL.t5 9.75419
R64 VTAIL.n10 VTAIL.t9 9.75419
R65 VTAIL.n22 VTAIL.t6 9.75419
R66 VTAIL.n22 VTAIL.t4 9.75419
R67 VTAIL.n12 VTAIL.t10 9.75419
R68 VTAIL.n12 VTAIL.t11 9.75419
R69 VTAIL.n35 VTAIL.n33 9.71174
R70 VTAIL.n5 VTAIL.n3 9.71174
R71 VTAIL.n27 VTAIL.n25 9.71174
R72 VTAIL.n17 VTAIL.n15 9.71174
R73 VTAIL.n38 VTAIL.n37 9.45567
R74 VTAIL.n8 VTAIL.n7 9.45567
R75 VTAIL.n30 VTAIL.n29 9.45567
R76 VTAIL.n20 VTAIL.n19 9.45567
R77 VTAIL.n37 VTAIL.n36 9.3005
R78 VTAIL.n7 VTAIL.n6 9.3005
R79 VTAIL.n29 VTAIL.n28 9.3005
R80 VTAIL.n19 VTAIL.n18 9.3005
R81 VTAIL.n38 VTAIL.n32 8.14595
R82 VTAIL.n8 VTAIL.n2 8.14595
R83 VTAIL.n30 VTAIL.n24 8.14595
R84 VTAIL.n20 VTAIL.n14 8.14595
R85 VTAIL.n36 VTAIL.n35 7.3702
R86 VTAIL.n6 VTAIL.n5 7.3702
R87 VTAIL.n28 VTAIL.n27 7.3702
R88 VTAIL.n18 VTAIL.n17 7.3702
R89 VTAIL.n36 VTAIL.n32 5.81868
R90 VTAIL.n6 VTAIL.n2 5.81868
R91 VTAIL.n28 VTAIL.n24 5.81868
R92 VTAIL.n18 VTAIL.n14 5.81868
R93 VTAIL.n37 VTAIL.n33 3.44771
R94 VTAIL.n7 VTAIL.n3 3.44771
R95 VTAIL.n29 VTAIL.n25 3.44771
R96 VTAIL.n19 VTAIL.n15 3.44771
R97 VTAIL.n21 VTAIL.n13 1.12981
R98 VTAIL.n31 VTAIL.n23 1.12981
R99 VTAIL.n11 VTAIL.n9 1.12981
R100 VTAIL.n23 VTAIL.n21 1.03498
R101 VTAIL.n9 VTAIL.n1 1.03498
R102 VTAIL VTAIL.n39 0.789293
R103 VTAIL VTAIL.n1 0.341017
R104 VDD1.n2 VDD1.n0 289.615
R105 VDD1.n9 VDD1.n7 289.615
R106 VDD1.n3 VDD1.n2 185
R107 VDD1.n10 VDD1.n9 185
R108 VDD1.t3 VDD1.n1 167.117
R109 VDD1.t4 VDD1.n8 167.117
R110 VDD1.n15 VDD1.n14 101.605
R111 VDD1.n17 VDD1.n16 101.377
R112 VDD1.n2 VDD1.t3 52.3082
R113 VDD1.n9 VDD1.t4 52.3082
R114 VDD1 VDD1.n6 49.5754
R115 VDD1.n15 VDD1.n13 49.4618
R116 VDD1.n17 VDD1.n15 30.2832
R117 VDD1.n16 VDD1.t2 9.75419
R118 VDD1.n16 VDD1.t1 9.75419
R119 VDD1.n14 VDD1.t0 9.75419
R120 VDD1.n14 VDD1.t5 9.75419
R121 VDD1.n3 VDD1.n1 9.71174
R122 VDD1.n10 VDD1.n8 9.71174
R123 VDD1.n6 VDD1.n5 9.45567
R124 VDD1.n13 VDD1.n12 9.45567
R125 VDD1.n5 VDD1.n4 9.3005
R126 VDD1.n12 VDD1.n11 9.3005
R127 VDD1.n6 VDD1.n0 8.14595
R128 VDD1.n13 VDD1.n7 8.14595
R129 VDD1.n4 VDD1.n3 7.3702
R130 VDD1.n11 VDD1.n10 7.3702
R131 VDD1.n4 VDD1.n0 5.81868
R132 VDD1.n11 VDD1.n7 5.81868
R133 VDD1.n5 VDD1.n1 3.44771
R134 VDD1.n12 VDD1.n8 3.44771
R135 VDD1 VDD1.n17 0.224638
R136 B.n367 B.n366 585
R137 B.n130 B.n62 585
R138 B.n129 B.n128 585
R139 B.n127 B.n126 585
R140 B.n125 B.n124 585
R141 B.n123 B.n122 585
R142 B.n121 B.n120 585
R143 B.n119 B.n118 585
R144 B.n117 B.n116 585
R145 B.n115 B.n114 585
R146 B.n113 B.n112 585
R147 B.n111 B.n110 585
R148 B.n109 B.n108 585
R149 B.n107 B.n106 585
R150 B.n105 B.n104 585
R151 B.n103 B.n102 585
R152 B.n101 B.n100 585
R153 B.n99 B.n98 585
R154 B.n97 B.n96 585
R155 B.n95 B.n94 585
R156 B.n93 B.n92 585
R157 B.n91 B.n90 585
R158 B.n89 B.n88 585
R159 B.n87 B.n86 585
R160 B.n85 B.n84 585
R161 B.n83 B.n82 585
R162 B.n81 B.n80 585
R163 B.n79 B.n78 585
R164 B.n77 B.n76 585
R165 B.n75 B.n74 585
R166 B.n73 B.n72 585
R167 B.n71 B.n70 585
R168 B.n46 B.n45 585
R169 B.n372 B.n371 585
R170 B.n365 B.n63 585
R171 B.n63 B.n43 585
R172 B.n364 B.n42 585
R173 B.n376 B.n42 585
R174 B.n363 B.n41 585
R175 B.n377 B.n41 585
R176 B.n362 B.n40 585
R177 B.n378 B.n40 585
R178 B.n361 B.n360 585
R179 B.n360 B.n36 585
R180 B.n359 B.n35 585
R181 B.n384 B.n35 585
R182 B.n358 B.n34 585
R183 B.n385 B.n34 585
R184 B.n357 B.n33 585
R185 B.n386 B.n33 585
R186 B.n356 B.n355 585
R187 B.n355 B.n29 585
R188 B.n354 B.n28 585
R189 B.n392 B.n28 585
R190 B.n353 B.n27 585
R191 B.n393 B.n27 585
R192 B.n352 B.n26 585
R193 B.n394 B.n26 585
R194 B.n351 B.n350 585
R195 B.n350 B.n25 585
R196 B.n349 B.n21 585
R197 B.n400 B.n21 585
R198 B.n348 B.n20 585
R199 B.n401 B.n20 585
R200 B.n347 B.n19 585
R201 B.n402 B.n19 585
R202 B.n346 B.n345 585
R203 B.n345 B.n18 585
R204 B.n344 B.n14 585
R205 B.n408 B.n14 585
R206 B.n343 B.n13 585
R207 B.n409 B.n13 585
R208 B.n342 B.n12 585
R209 B.n410 B.n12 585
R210 B.n341 B.n340 585
R211 B.n340 B.n339 585
R212 B.n338 B.n337 585
R213 B.n338 B.n8 585
R214 B.n336 B.n7 585
R215 B.n417 B.n7 585
R216 B.n335 B.n6 585
R217 B.n418 B.n6 585
R218 B.n334 B.n5 585
R219 B.n419 B.n5 585
R220 B.n333 B.n332 585
R221 B.n332 B.n4 585
R222 B.n331 B.n131 585
R223 B.n331 B.n330 585
R224 B.n321 B.n132 585
R225 B.n133 B.n132 585
R226 B.n323 B.n322 585
R227 B.n324 B.n323 585
R228 B.n320 B.n138 585
R229 B.n138 B.n137 585
R230 B.n319 B.n318 585
R231 B.n318 B.n317 585
R232 B.n140 B.n139 585
R233 B.n310 B.n140 585
R234 B.n309 B.n308 585
R235 B.n311 B.n309 585
R236 B.n307 B.n145 585
R237 B.n145 B.n144 585
R238 B.n306 B.n305 585
R239 B.n305 B.n304 585
R240 B.n147 B.n146 585
R241 B.n297 B.n147 585
R242 B.n296 B.n295 585
R243 B.n298 B.n296 585
R244 B.n294 B.n152 585
R245 B.n152 B.n151 585
R246 B.n293 B.n292 585
R247 B.n292 B.n291 585
R248 B.n154 B.n153 585
R249 B.n155 B.n154 585
R250 B.n284 B.n283 585
R251 B.n285 B.n284 585
R252 B.n282 B.n160 585
R253 B.n160 B.n159 585
R254 B.n281 B.n280 585
R255 B.n280 B.n279 585
R256 B.n162 B.n161 585
R257 B.n163 B.n162 585
R258 B.n272 B.n271 585
R259 B.n273 B.n272 585
R260 B.n270 B.n168 585
R261 B.n168 B.n167 585
R262 B.n269 B.n268 585
R263 B.n268 B.n267 585
R264 B.n170 B.n169 585
R265 B.n171 B.n170 585
R266 B.n263 B.n262 585
R267 B.n174 B.n173 585
R268 B.n259 B.n258 585
R269 B.n260 B.n259 585
R270 B.n257 B.n191 585
R271 B.n256 B.n255 585
R272 B.n254 B.n253 585
R273 B.n252 B.n251 585
R274 B.n250 B.n249 585
R275 B.n248 B.n247 585
R276 B.n246 B.n245 585
R277 B.n244 B.n243 585
R278 B.n242 B.n241 585
R279 B.n239 B.n238 585
R280 B.n237 B.n236 585
R281 B.n235 B.n234 585
R282 B.n233 B.n232 585
R283 B.n231 B.n230 585
R284 B.n229 B.n228 585
R285 B.n227 B.n226 585
R286 B.n225 B.n224 585
R287 B.n223 B.n222 585
R288 B.n221 B.n220 585
R289 B.n218 B.n217 585
R290 B.n216 B.n215 585
R291 B.n214 B.n213 585
R292 B.n212 B.n211 585
R293 B.n210 B.n209 585
R294 B.n208 B.n207 585
R295 B.n206 B.n205 585
R296 B.n204 B.n203 585
R297 B.n202 B.n201 585
R298 B.n200 B.n199 585
R299 B.n198 B.n197 585
R300 B.n196 B.n190 585
R301 B.n260 B.n190 585
R302 B.n264 B.n172 585
R303 B.n172 B.n171 585
R304 B.n266 B.n265 585
R305 B.n267 B.n266 585
R306 B.n166 B.n165 585
R307 B.n167 B.n166 585
R308 B.n275 B.n274 585
R309 B.n274 B.n273 585
R310 B.n276 B.n164 585
R311 B.n164 B.n163 585
R312 B.n278 B.n277 585
R313 B.n279 B.n278 585
R314 B.n158 B.n157 585
R315 B.n159 B.n158 585
R316 B.n287 B.n286 585
R317 B.n286 B.n285 585
R318 B.n288 B.n156 585
R319 B.n156 B.n155 585
R320 B.n290 B.n289 585
R321 B.n291 B.n290 585
R322 B.n150 B.n149 585
R323 B.n151 B.n150 585
R324 B.n300 B.n299 585
R325 B.n299 B.n298 585
R326 B.n301 B.n148 585
R327 B.n297 B.n148 585
R328 B.n303 B.n302 585
R329 B.n304 B.n303 585
R330 B.n143 B.n142 585
R331 B.n144 B.n143 585
R332 B.n313 B.n312 585
R333 B.n312 B.n311 585
R334 B.n314 B.n141 585
R335 B.n310 B.n141 585
R336 B.n316 B.n315 585
R337 B.n317 B.n316 585
R338 B.n136 B.n135 585
R339 B.n137 B.n136 585
R340 B.n326 B.n325 585
R341 B.n325 B.n324 585
R342 B.n327 B.n134 585
R343 B.n134 B.n133 585
R344 B.n329 B.n328 585
R345 B.n330 B.n329 585
R346 B.n3 B.n0 585
R347 B.n4 B.n3 585
R348 B.n416 B.n1 585
R349 B.n417 B.n416 585
R350 B.n415 B.n414 585
R351 B.n415 B.n8 585
R352 B.n413 B.n9 585
R353 B.n339 B.n9 585
R354 B.n412 B.n411 585
R355 B.n411 B.n410 585
R356 B.n11 B.n10 585
R357 B.n409 B.n11 585
R358 B.n407 B.n406 585
R359 B.n408 B.n407 585
R360 B.n405 B.n15 585
R361 B.n18 B.n15 585
R362 B.n404 B.n403 585
R363 B.n403 B.n402 585
R364 B.n17 B.n16 585
R365 B.n401 B.n17 585
R366 B.n399 B.n398 585
R367 B.n400 B.n399 585
R368 B.n397 B.n22 585
R369 B.n25 B.n22 585
R370 B.n396 B.n395 585
R371 B.n395 B.n394 585
R372 B.n24 B.n23 585
R373 B.n393 B.n24 585
R374 B.n391 B.n390 585
R375 B.n392 B.n391 585
R376 B.n389 B.n30 585
R377 B.n30 B.n29 585
R378 B.n388 B.n387 585
R379 B.n387 B.n386 585
R380 B.n32 B.n31 585
R381 B.n385 B.n32 585
R382 B.n383 B.n382 585
R383 B.n384 B.n383 585
R384 B.n381 B.n37 585
R385 B.n37 B.n36 585
R386 B.n380 B.n379 585
R387 B.n379 B.n378 585
R388 B.n39 B.n38 585
R389 B.n377 B.n39 585
R390 B.n375 B.n374 585
R391 B.n376 B.n375 585
R392 B.n373 B.n44 585
R393 B.n44 B.n43 585
R394 B.n420 B.n419 585
R395 B.n418 B.n2 585
R396 B.n371 B.n44 516.524
R397 B.n367 B.n63 516.524
R398 B.n190 B.n170 516.524
R399 B.n262 B.n172 516.524
R400 B.n369 B.n368 256.663
R401 B.n369 B.n61 256.663
R402 B.n369 B.n60 256.663
R403 B.n369 B.n59 256.663
R404 B.n369 B.n58 256.663
R405 B.n369 B.n57 256.663
R406 B.n369 B.n56 256.663
R407 B.n369 B.n55 256.663
R408 B.n369 B.n54 256.663
R409 B.n369 B.n53 256.663
R410 B.n369 B.n52 256.663
R411 B.n369 B.n51 256.663
R412 B.n369 B.n50 256.663
R413 B.n369 B.n49 256.663
R414 B.n369 B.n48 256.663
R415 B.n369 B.n47 256.663
R416 B.n370 B.n369 256.663
R417 B.n261 B.n260 256.663
R418 B.n260 B.n175 256.663
R419 B.n260 B.n176 256.663
R420 B.n260 B.n177 256.663
R421 B.n260 B.n178 256.663
R422 B.n260 B.n179 256.663
R423 B.n260 B.n180 256.663
R424 B.n260 B.n181 256.663
R425 B.n260 B.n182 256.663
R426 B.n260 B.n183 256.663
R427 B.n260 B.n184 256.663
R428 B.n260 B.n185 256.663
R429 B.n260 B.n186 256.663
R430 B.n260 B.n187 256.663
R431 B.n260 B.n188 256.663
R432 B.n260 B.n189 256.663
R433 B.n422 B.n421 256.663
R434 B.n67 B.t6 252.709
R435 B.n64 B.t17 252.709
R436 B.n194 B.t10 252.709
R437 B.n192 B.t14 252.709
R438 B.n260 B.n171 188.227
R439 B.n369 B.n43 188.227
R440 B.n70 B.n46 163.367
R441 B.n74 B.n73 163.367
R442 B.n78 B.n77 163.367
R443 B.n82 B.n81 163.367
R444 B.n86 B.n85 163.367
R445 B.n90 B.n89 163.367
R446 B.n94 B.n93 163.367
R447 B.n98 B.n97 163.367
R448 B.n102 B.n101 163.367
R449 B.n106 B.n105 163.367
R450 B.n110 B.n109 163.367
R451 B.n114 B.n113 163.367
R452 B.n118 B.n117 163.367
R453 B.n122 B.n121 163.367
R454 B.n126 B.n125 163.367
R455 B.n128 B.n62 163.367
R456 B.n268 B.n170 163.367
R457 B.n268 B.n168 163.367
R458 B.n272 B.n168 163.367
R459 B.n272 B.n162 163.367
R460 B.n280 B.n162 163.367
R461 B.n280 B.n160 163.367
R462 B.n284 B.n160 163.367
R463 B.n284 B.n154 163.367
R464 B.n292 B.n154 163.367
R465 B.n292 B.n152 163.367
R466 B.n296 B.n152 163.367
R467 B.n296 B.n147 163.367
R468 B.n305 B.n147 163.367
R469 B.n305 B.n145 163.367
R470 B.n309 B.n145 163.367
R471 B.n309 B.n140 163.367
R472 B.n318 B.n140 163.367
R473 B.n318 B.n138 163.367
R474 B.n323 B.n138 163.367
R475 B.n323 B.n132 163.367
R476 B.n331 B.n132 163.367
R477 B.n332 B.n331 163.367
R478 B.n332 B.n5 163.367
R479 B.n6 B.n5 163.367
R480 B.n7 B.n6 163.367
R481 B.n338 B.n7 163.367
R482 B.n340 B.n338 163.367
R483 B.n340 B.n12 163.367
R484 B.n13 B.n12 163.367
R485 B.n14 B.n13 163.367
R486 B.n345 B.n14 163.367
R487 B.n345 B.n19 163.367
R488 B.n20 B.n19 163.367
R489 B.n21 B.n20 163.367
R490 B.n350 B.n21 163.367
R491 B.n350 B.n26 163.367
R492 B.n27 B.n26 163.367
R493 B.n28 B.n27 163.367
R494 B.n355 B.n28 163.367
R495 B.n355 B.n33 163.367
R496 B.n34 B.n33 163.367
R497 B.n35 B.n34 163.367
R498 B.n360 B.n35 163.367
R499 B.n360 B.n40 163.367
R500 B.n41 B.n40 163.367
R501 B.n42 B.n41 163.367
R502 B.n63 B.n42 163.367
R503 B.n259 B.n174 163.367
R504 B.n259 B.n191 163.367
R505 B.n255 B.n254 163.367
R506 B.n251 B.n250 163.367
R507 B.n247 B.n246 163.367
R508 B.n243 B.n242 163.367
R509 B.n238 B.n237 163.367
R510 B.n234 B.n233 163.367
R511 B.n230 B.n229 163.367
R512 B.n226 B.n225 163.367
R513 B.n222 B.n221 163.367
R514 B.n217 B.n216 163.367
R515 B.n213 B.n212 163.367
R516 B.n209 B.n208 163.367
R517 B.n205 B.n204 163.367
R518 B.n201 B.n200 163.367
R519 B.n197 B.n190 163.367
R520 B.n266 B.n172 163.367
R521 B.n266 B.n166 163.367
R522 B.n274 B.n166 163.367
R523 B.n274 B.n164 163.367
R524 B.n278 B.n164 163.367
R525 B.n278 B.n158 163.367
R526 B.n286 B.n158 163.367
R527 B.n286 B.n156 163.367
R528 B.n290 B.n156 163.367
R529 B.n290 B.n150 163.367
R530 B.n299 B.n150 163.367
R531 B.n299 B.n148 163.367
R532 B.n303 B.n148 163.367
R533 B.n303 B.n143 163.367
R534 B.n312 B.n143 163.367
R535 B.n312 B.n141 163.367
R536 B.n316 B.n141 163.367
R537 B.n316 B.n136 163.367
R538 B.n325 B.n136 163.367
R539 B.n325 B.n134 163.367
R540 B.n329 B.n134 163.367
R541 B.n329 B.n3 163.367
R542 B.n420 B.n3 163.367
R543 B.n416 B.n2 163.367
R544 B.n416 B.n415 163.367
R545 B.n415 B.n9 163.367
R546 B.n411 B.n9 163.367
R547 B.n411 B.n11 163.367
R548 B.n407 B.n11 163.367
R549 B.n407 B.n15 163.367
R550 B.n403 B.n15 163.367
R551 B.n403 B.n17 163.367
R552 B.n399 B.n17 163.367
R553 B.n399 B.n22 163.367
R554 B.n395 B.n22 163.367
R555 B.n395 B.n24 163.367
R556 B.n391 B.n24 163.367
R557 B.n391 B.n30 163.367
R558 B.n387 B.n30 163.367
R559 B.n387 B.n32 163.367
R560 B.n383 B.n32 163.367
R561 B.n383 B.n37 163.367
R562 B.n379 B.n37 163.367
R563 B.n379 B.n39 163.367
R564 B.n375 B.n39 163.367
R565 B.n375 B.n44 163.367
R566 B.n64 B.t18 149.006
R567 B.n194 B.t13 149.006
R568 B.n67 B.t8 149.006
R569 B.n192 B.t16 149.006
R570 B.n65 B.t19 123.6
R571 B.n195 B.t12 123.6
R572 B.n68 B.t9 123.6
R573 B.n193 B.t15 123.6
R574 B.n267 B.n171 102.397
R575 B.n267 B.n167 102.397
R576 B.n273 B.n167 102.397
R577 B.n273 B.n163 102.397
R578 B.n279 B.n163 102.397
R579 B.n285 B.n159 102.397
R580 B.n285 B.n155 102.397
R581 B.n291 B.n155 102.397
R582 B.n291 B.n151 102.397
R583 B.n298 B.n151 102.397
R584 B.n298 B.n297 102.397
R585 B.n304 B.n144 102.397
R586 B.n311 B.n144 102.397
R587 B.n311 B.n310 102.397
R588 B.n317 B.n137 102.397
R589 B.n324 B.n137 102.397
R590 B.n330 B.n133 102.397
R591 B.n330 B.n4 102.397
R592 B.n419 B.n4 102.397
R593 B.n419 B.n418 102.397
R594 B.n418 B.n417 102.397
R595 B.n417 B.n8 102.397
R596 B.n339 B.n8 102.397
R597 B.n410 B.n409 102.397
R598 B.n409 B.n408 102.397
R599 B.n402 B.n18 102.397
R600 B.n402 B.n401 102.397
R601 B.n401 B.n400 102.397
R602 B.n394 B.n25 102.397
R603 B.n394 B.n393 102.397
R604 B.n393 B.n392 102.397
R605 B.n392 B.n29 102.397
R606 B.n386 B.n29 102.397
R607 B.n386 B.n385 102.397
R608 B.n384 B.n36 102.397
R609 B.n378 B.n36 102.397
R610 B.n378 B.n377 102.397
R611 B.n377 B.n376 102.397
R612 B.n376 B.n43 102.397
R613 B.n324 B.t1 99.3845
R614 B.n410 B.t0 99.3845
R615 B.n317 B.t4 90.3496
R616 B.n408 B.t2 90.3496
R617 B.t11 B.n159 81.3147
R618 B.n385 B.t7 81.3147
R619 B.n304 B.t5 75.2914
R620 B.n400 B.t3 75.2914
R621 B.n371 B.n370 71.676
R622 B.n70 B.n47 71.676
R623 B.n74 B.n48 71.676
R624 B.n78 B.n49 71.676
R625 B.n82 B.n50 71.676
R626 B.n86 B.n51 71.676
R627 B.n90 B.n52 71.676
R628 B.n94 B.n53 71.676
R629 B.n98 B.n54 71.676
R630 B.n102 B.n55 71.676
R631 B.n106 B.n56 71.676
R632 B.n110 B.n57 71.676
R633 B.n114 B.n58 71.676
R634 B.n118 B.n59 71.676
R635 B.n122 B.n60 71.676
R636 B.n126 B.n61 71.676
R637 B.n368 B.n62 71.676
R638 B.n368 B.n367 71.676
R639 B.n128 B.n61 71.676
R640 B.n125 B.n60 71.676
R641 B.n121 B.n59 71.676
R642 B.n117 B.n58 71.676
R643 B.n113 B.n57 71.676
R644 B.n109 B.n56 71.676
R645 B.n105 B.n55 71.676
R646 B.n101 B.n54 71.676
R647 B.n97 B.n53 71.676
R648 B.n93 B.n52 71.676
R649 B.n89 B.n51 71.676
R650 B.n85 B.n50 71.676
R651 B.n81 B.n49 71.676
R652 B.n77 B.n48 71.676
R653 B.n73 B.n47 71.676
R654 B.n370 B.n46 71.676
R655 B.n262 B.n261 71.676
R656 B.n191 B.n175 71.676
R657 B.n254 B.n176 71.676
R658 B.n250 B.n177 71.676
R659 B.n246 B.n178 71.676
R660 B.n242 B.n179 71.676
R661 B.n237 B.n180 71.676
R662 B.n233 B.n181 71.676
R663 B.n229 B.n182 71.676
R664 B.n225 B.n183 71.676
R665 B.n221 B.n184 71.676
R666 B.n216 B.n185 71.676
R667 B.n212 B.n186 71.676
R668 B.n208 B.n187 71.676
R669 B.n204 B.n188 71.676
R670 B.n200 B.n189 71.676
R671 B.n261 B.n174 71.676
R672 B.n255 B.n175 71.676
R673 B.n251 B.n176 71.676
R674 B.n247 B.n177 71.676
R675 B.n243 B.n178 71.676
R676 B.n238 B.n179 71.676
R677 B.n234 B.n180 71.676
R678 B.n230 B.n181 71.676
R679 B.n226 B.n182 71.676
R680 B.n222 B.n183 71.676
R681 B.n217 B.n184 71.676
R682 B.n213 B.n185 71.676
R683 B.n209 B.n186 71.676
R684 B.n205 B.n187 71.676
R685 B.n201 B.n188 71.676
R686 B.n197 B.n189 71.676
R687 B.n421 B.n420 71.676
R688 B.n421 B.n2 71.676
R689 B.n69 B.n68 59.5399
R690 B.n66 B.n65 59.5399
R691 B.n219 B.n195 59.5399
R692 B.n240 B.n193 59.5399
R693 B.n264 B.n263 33.5615
R694 B.n196 B.n169 33.5615
R695 B.n366 B.n365 33.5615
R696 B.n373 B.n372 33.5615
R697 B.n297 B.t5 27.1052
R698 B.n25 B.t3 27.1052
R699 B.n68 B.n67 25.4066
R700 B.n65 B.n64 25.4066
R701 B.n195 B.n194 25.4066
R702 B.n193 B.n192 25.4066
R703 B.n279 B.t11 21.082
R704 B.t7 B.n384 21.082
R705 B B.n422 18.0485
R706 B.n310 B.t4 12.047
R707 B.n18 B.t2 12.047
R708 B.n265 B.n264 10.6151
R709 B.n265 B.n165 10.6151
R710 B.n275 B.n165 10.6151
R711 B.n276 B.n275 10.6151
R712 B.n277 B.n276 10.6151
R713 B.n277 B.n157 10.6151
R714 B.n287 B.n157 10.6151
R715 B.n288 B.n287 10.6151
R716 B.n289 B.n288 10.6151
R717 B.n289 B.n149 10.6151
R718 B.n300 B.n149 10.6151
R719 B.n301 B.n300 10.6151
R720 B.n302 B.n301 10.6151
R721 B.n302 B.n142 10.6151
R722 B.n313 B.n142 10.6151
R723 B.n314 B.n313 10.6151
R724 B.n315 B.n314 10.6151
R725 B.n315 B.n135 10.6151
R726 B.n326 B.n135 10.6151
R727 B.n327 B.n326 10.6151
R728 B.n328 B.n327 10.6151
R729 B.n328 B.n0 10.6151
R730 B.n263 B.n173 10.6151
R731 B.n258 B.n173 10.6151
R732 B.n258 B.n257 10.6151
R733 B.n257 B.n256 10.6151
R734 B.n256 B.n253 10.6151
R735 B.n253 B.n252 10.6151
R736 B.n252 B.n249 10.6151
R737 B.n249 B.n248 10.6151
R738 B.n248 B.n245 10.6151
R739 B.n245 B.n244 10.6151
R740 B.n244 B.n241 10.6151
R741 B.n239 B.n236 10.6151
R742 B.n236 B.n235 10.6151
R743 B.n235 B.n232 10.6151
R744 B.n232 B.n231 10.6151
R745 B.n231 B.n228 10.6151
R746 B.n228 B.n227 10.6151
R747 B.n227 B.n224 10.6151
R748 B.n224 B.n223 10.6151
R749 B.n223 B.n220 10.6151
R750 B.n218 B.n215 10.6151
R751 B.n215 B.n214 10.6151
R752 B.n214 B.n211 10.6151
R753 B.n211 B.n210 10.6151
R754 B.n210 B.n207 10.6151
R755 B.n207 B.n206 10.6151
R756 B.n206 B.n203 10.6151
R757 B.n203 B.n202 10.6151
R758 B.n202 B.n199 10.6151
R759 B.n199 B.n198 10.6151
R760 B.n198 B.n196 10.6151
R761 B.n269 B.n169 10.6151
R762 B.n270 B.n269 10.6151
R763 B.n271 B.n270 10.6151
R764 B.n271 B.n161 10.6151
R765 B.n281 B.n161 10.6151
R766 B.n282 B.n281 10.6151
R767 B.n283 B.n282 10.6151
R768 B.n283 B.n153 10.6151
R769 B.n293 B.n153 10.6151
R770 B.n294 B.n293 10.6151
R771 B.n295 B.n294 10.6151
R772 B.n295 B.n146 10.6151
R773 B.n306 B.n146 10.6151
R774 B.n307 B.n306 10.6151
R775 B.n308 B.n307 10.6151
R776 B.n308 B.n139 10.6151
R777 B.n319 B.n139 10.6151
R778 B.n320 B.n319 10.6151
R779 B.n322 B.n320 10.6151
R780 B.n322 B.n321 10.6151
R781 B.n321 B.n131 10.6151
R782 B.n333 B.n131 10.6151
R783 B.n334 B.n333 10.6151
R784 B.n335 B.n334 10.6151
R785 B.n336 B.n335 10.6151
R786 B.n337 B.n336 10.6151
R787 B.n341 B.n337 10.6151
R788 B.n342 B.n341 10.6151
R789 B.n343 B.n342 10.6151
R790 B.n344 B.n343 10.6151
R791 B.n346 B.n344 10.6151
R792 B.n347 B.n346 10.6151
R793 B.n348 B.n347 10.6151
R794 B.n349 B.n348 10.6151
R795 B.n351 B.n349 10.6151
R796 B.n352 B.n351 10.6151
R797 B.n353 B.n352 10.6151
R798 B.n354 B.n353 10.6151
R799 B.n356 B.n354 10.6151
R800 B.n357 B.n356 10.6151
R801 B.n358 B.n357 10.6151
R802 B.n359 B.n358 10.6151
R803 B.n361 B.n359 10.6151
R804 B.n362 B.n361 10.6151
R805 B.n363 B.n362 10.6151
R806 B.n364 B.n363 10.6151
R807 B.n365 B.n364 10.6151
R808 B.n414 B.n1 10.6151
R809 B.n414 B.n413 10.6151
R810 B.n413 B.n412 10.6151
R811 B.n412 B.n10 10.6151
R812 B.n406 B.n10 10.6151
R813 B.n406 B.n405 10.6151
R814 B.n405 B.n404 10.6151
R815 B.n404 B.n16 10.6151
R816 B.n398 B.n16 10.6151
R817 B.n398 B.n397 10.6151
R818 B.n397 B.n396 10.6151
R819 B.n396 B.n23 10.6151
R820 B.n390 B.n23 10.6151
R821 B.n390 B.n389 10.6151
R822 B.n389 B.n388 10.6151
R823 B.n388 B.n31 10.6151
R824 B.n382 B.n31 10.6151
R825 B.n382 B.n381 10.6151
R826 B.n381 B.n380 10.6151
R827 B.n380 B.n38 10.6151
R828 B.n374 B.n38 10.6151
R829 B.n374 B.n373 10.6151
R830 B.n372 B.n45 10.6151
R831 B.n71 B.n45 10.6151
R832 B.n72 B.n71 10.6151
R833 B.n75 B.n72 10.6151
R834 B.n76 B.n75 10.6151
R835 B.n79 B.n76 10.6151
R836 B.n80 B.n79 10.6151
R837 B.n83 B.n80 10.6151
R838 B.n84 B.n83 10.6151
R839 B.n87 B.n84 10.6151
R840 B.n88 B.n87 10.6151
R841 B.n92 B.n91 10.6151
R842 B.n95 B.n92 10.6151
R843 B.n96 B.n95 10.6151
R844 B.n99 B.n96 10.6151
R845 B.n100 B.n99 10.6151
R846 B.n103 B.n100 10.6151
R847 B.n104 B.n103 10.6151
R848 B.n107 B.n104 10.6151
R849 B.n108 B.n107 10.6151
R850 B.n112 B.n111 10.6151
R851 B.n115 B.n112 10.6151
R852 B.n116 B.n115 10.6151
R853 B.n119 B.n116 10.6151
R854 B.n120 B.n119 10.6151
R855 B.n123 B.n120 10.6151
R856 B.n124 B.n123 10.6151
R857 B.n127 B.n124 10.6151
R858 B.n129 B.n127 10.6151
R859 B.n130 B.n129 10.6151
R860 B.n366 B.n130 10.6151
R861 B.n241 B.n240 9.36635
R862 B.n219 B.n218 9.36635
R863 B.n88 B.n69 9.36635
R864 B.n111 B.n66 9.36635
R865 B.n422 B.n0 8.11757
R866 B.n422 B.n1 8.11757
R867 B.t1 B.n133 3.01214
R868 B.n339 B.t0 3.01214
R869 B.n240 B.n239 1.24928
R870 B.n220 B.n219 1.24928
R871 B.n91 B.n69 1.24928
R872 B.n108 B.n66 1.24928
R873 VN.n7 VN.n6 161.3
R874 VN.n15 VN.n14 161.3
R875 VN.n13 VN.n8 161.3
R876 VN.n12 VN.n11 161.3
R877 VN.n5 VN.n0 161.3
R878 VN.n4 VN.n3 161.3
R879 VN.n2 VN.t2 109.773
R880 VN.n10 VN.t3 109.773
R881 VN.n6 VN.t5 90.2525
R882 VN.n14 VN.t1 90.2525
R883 VN.n1 VN.t4 49.9219
R884 VN.n9 VN.t0 49.9219
R885 VN.n5 VN.n4 49.7204
R886 VN.n13 VN.n12 49.7204
R887 VN.n11 VN.n10 43.1531
R888 VN.n3 VN.n2 43.1531
R889 VN.n2 VN.n1 42.1911
R890 VN.n10 VN.n9 42.1911
R891 VN VN.n15 35.2183
R892 VN.n4 VN.n1 12.234
R893 VN.n12 VN.n9 12.234
R894 VN.n6 VN.n5 10.2247
R895 VN.n14 VN.n13 10.2247
R896 VN.n15 VN.n8 0.189894
R897 VN.n11 VN.n8 0.189894
R898 VN.n3 VN.n0 0.189894
R899 VN.n7 VN.n0 0.189894
R900 VN VN.n7 0.0516364
R901 VDD2.n11 VDD2.n9 289.615
R902 VDD2.n2 VDD2.n0 289.615
R903 VDD2.n12 VDD2.n11 185
R904 VDD2.n3 VDD2.n2 185
R905 VDD2.t4 VDD2.n10 167.117
R906 VDD2.t3 VDD2.n1 167.117
R907 VDD2.n8 VDD2.n7 101.605
R908 VDD2 VDD2.n17 101.602
R909 VDD2.n11 VDD2.t4 52.3082
R910 VDD2.n2 VDD2.t3 52.3082
R911 VDD2.n8 VDD2.n6 49.4618
R912 VDD2.n16 VDD2.n15 48.6702
R913 VDD2.n16 VDD2.n8 29.1356
R914 VDD2.n17 VDD2.t5 9.75419
R915 VDD2.n17 VDD2.t2 9.75419
R916 VDD2.n7 VDD2.t1 9.75419
R917 VDD2.n7 VDD2.t0 9.75419
R918 VDD2.n12 VDD2.n10 9.71174
R919 VDD2.n3 VDD2.n1 9.71174
R920 VDD2.n15 VDD2.n14 9.45567
R921 VDD2.n6 VDD2.n5 9.45567
R922 VDD2.n14 VDD2.n13 9.3005
R923 VDD2.n5 VDD2.n4 9.3005
R924 VDD2.n15 VDD2.n9 8.14595
R925 VDD2.n6 VDD2.n0 8.14595
R926 VDD2.n13 VDD2.n12 7.3702
R927 VDD2.n4 VDD2.n3 7.3702
R928 VDD2.n13 VDD2.n9 5.81868
R929 VDD2.n4 VDD2.n0 5.81868
R930 VDD2.n14 VDD2.n10 3.44771
R931 VDD2.n5 VDD2.n1 3.44771
R932 VDD2 VDD2.n16 0.905672
C0 VTAIL VN 1.43625f
C1 VDD2 VN 1.14409f
C2 VDD1 VTAIL 3.23213f
C3 VDD1 VDD2 0.810163f
C4 VTAIL VP 1.45043f
C5 VDD2 VP 0.326883f
C6 VTAIL VDD2 3.27383f
C7 VDD1 VN 0.154778f
C8 VP VN 3.50982f
C9 VDD1 VP 1.31428f
C10 VDD2 B 2.811093f
C11 VDD1 B 2.893592f
C12 VTAIL B 2.636957f
C13 VN B 6.671124f
C14 VP B 5.751659f
C15 VDD2.n0 B 0.025428f
C16 VDD2.n1 B 0.056144f
C17 VDD2.t3 B 0.042082f
C18 VDD2.n2 B 0.044047f
C19 VDD2.n3 B 0.014001f
C20 VDD2.n4 B 0.009234f
C21 VDD2.n5 B 0.124432f
C22 VDD2.n6 B 0.041027f
C23 VDD2.t1 B 0.027565f
C24 VDD2.t0 B 0.027565f
C25 VDD2.n7 B 0.173919f
C26 VDD2.n8 B 0.94843f
C27 VDD2.n9 B 0.025428f
C28 VDD2.n10 B 0.056144f
C29 VDD2.t4 B 0.042082f
C30 VDD2.n11 B 0.044047f
C31 VDD2.n12 B 0.014001f
C32 VDD2.n13 B 0.009234f
C33 VDD2.n14 B 0.124432f
C34 VDD2.n15 B 0.03979f
C35 VDD2.n16 B 0.905433f
C36 VDD2.t5 B 0.027565f
C37 VDD2.t2 B 0.027565f
C38 VDD2.n17 B 0.17391f
C39 VN.n0 B 0.025945f
C40 VN.t4 B 0.120899f
C41 VN.n1 B 0.098221f
C42 VN.t2 B 0.179632f
C43 VN.n2 B 0.104749f
C44 VN.n3 B 0.112806f
C45 VN.n4 B 0.035934f
C46 VN.n5 B 0.009577f
C47 VN.t5 B 0.159852f
C48 VN.n6 B 0.104576f
C49 VN.n7 B 0.020107f
C50 VN.n8 B 0.025945f
C51 VN.t0 B 0.120899f
C52 VN.n9 B 0.098221f
C53 VN.t3 B 0.179632f
C54 VN.n10 B 0.104749f
C55 VN.n11 B 0.112806f
C56 VN.n12 B 0.035934f
C57 VN.n13 B 0.009577f
C58 VN.t1 B 0.159852f
C59 VN.n14 B 0.104576f
C60 VN.n15 B 0.78344f
C61 VDD1.n0 B 0.024192f
C62 VDD1.n1 B 0.053416f
C63 VDD1.t3 B 0.040037f
C64 VDD1.n2 B 0.041906f
C65 VDD1.n3 B 0.01332f
C66 VDD1.n4 B 0.008785f
C67 VDD1.n5 B 0.118385f
C68 VDD1.n6 B 0.039299f
C69 VDD1.n7 B 0.024192f
C70 VDD1.n8 B 0.053416f
C71 VDD1.t4 B 0.040037f
C72 VDD1.n9 B 0.041906f
C73 VDD1.n10 B 0.01332f
C74 VDD1.n11 B 0.008785f
C75 VDD1.n12 B 0.118385f
C76 VDD1.n13 B 0.039033f
C77 VDD1.t0 B 0.026226f
C78 VDD1.t5 B 0.026226f
C79 VDD1.n14 B 0.165466f
C80 VDD1.n15 B 0.953003f
C81 VDD1.t2 B 0.026226f
C82 VDD1.t1 B 0.026226f
C83 VDD1.n16 B 0.165007f
C84 VDD1.n17 B 0.996124f
C85 VTAIL.t0 B 0.034402f
C86 VTAIL.t2 B 0.034402f
C87 VTAIL.n0 B 0.184672f
C88 VTAIL.n1 B 0.263103f
C89 VTAIL.n2 B 0.031735f
C90 VTAIL.n3 B 0.070069f
C91 VTAIL.t8 B 0.052519f
C92 VTAIL.n4 B 0.054971f
C93 VTAIL.n5 B 0.017473f
C94 VTAIL.n6 B 0.011524f
C95 VTAIL.n7 B 0.155293f
C96 VTAIL.n8 B 0.034849f
C97 VTAIL.n9 B 0.167672f
C98 VTAIL.t5 B 0.034402f
C99 VTAIL.t9 B 0.034402f
C100 VTAIL.n10 B 0.184672f
C101 VTAIL.n11 B 0.814437f
C102 VTAIL.t10 B 0.034402f
C103 VTAIL.t11 B 0.034402f
C104 VTAIL.n12 B 0.184673f
C105 VTAIL.n13 B 0.814436f
C106 VTAIL.n14 B 0.031735f
C107 VTAIL.n15 B 0.070069f
C108 VTAIL.t1 B 0.052519f
C109 VTAIL.n16 B 0.054971f
C110 VTAIL.n17 B 0.017473f
C111 VTAIL.n18 B 0.011524f
C112 VTAIL.n19 B 0.155293f
C113 VTAIL.n20 B 0.034849f
C114 VTAIL.n21 B 0.167672f
C115 VTAIL.t6 B 0.034402f
C116 VTAIL.t4 B 0.034402f
C117 VTAIL.n22 B 0.184673f
C118 VTAIL.n23 B 0.317608f
C119 VTAIL.n24 B 0.031735f
C120 VTAIL.n25 B 0.070069f
C121 VTAIL.t7 B 0.052519f
C122 VTAIL.n26 B 0.054971f
C123 VTAIL.n27 B 0.017473f
C124 VTAIL.n28 B 0.011524f
C125 VTAIL.n29 B 0.155293f
C126 VTAIL.n30 B 0.034849f
C127 VTAIL.n31 B 0.586463f
C128 VTAIL.n32 B 0.031735f
C129 VTAIL.n33 B 0.070069f
C130 VTAIL.t3 B 0.052519f
C131 VTAIL.n34 B 0.054971f
C132 VTAIL.n35 B 0.017473f
C133 VTAIL.n36 B 0.011524f
C134 VTAIL.n37 B 0.155293f
C135 VTAIL.n38 B 0.034849f
C136 VTAIL.n39 B 0.562933f
C137 VP.n0 B 0.026218f
C138 VP.t5 B 0.122172f
C139 VP.n1 B 0.07285f
C140 VP.n2 B 0.026218f
C141 VP.n3 B 0.026218f
C142 VP.t4 B 0.161536f
C143 VP.t3 B 0.122172f
C144 VP.n4 B 0.099255f
C145 VP.t2 B 0.181523f
C146 VP.n5 B 0.105852f
C147 VP.n6 B 0.113994f
C148 VP.n7 B 0.036312f
C149 VP.n8 B 0.009678f
C150 VP.n9 B 0.105677f
C151 VP.n10 B 0.774256f
C152 VP.n11 B 0.80131f
C153 VP.t1 B 0.161536f
C154 VP.n12 B 0.105677f
C155 VP.n13 B 0.009678f
C156 VP.n14 B 0.036312f
C157 VP.n15 B 0.026218f
C158 VP.n16 B 0.026218f
C159 VP.n17 B 0.036312f
C160 VP.n18 B 0.009678f
C161 VP.t0 B 0.161536f
C162 VP.n19 B 0.105677f
C163 VP.n20 B 0.020318f
.ends

