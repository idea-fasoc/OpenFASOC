* NGSPICE file created from diff_pair_sample_1764.ext - technology: sky130A

.subckt diff_pair_sample_1764 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X1 VTAIL.t6 VP.t0 VDD1.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X2 VTAIL.t18 VN.t1 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X3 VDD1.t8 VP.t1 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=2.6676 ps=14.46 w=6.84 l=1.92
X4 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X5 VTAIL.t3 VP.t3 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X6 VDD2.t7 VN.t2 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=1.1286 ps=7.17 w=6.84 l=1.92
X7 VDD1.t5 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=1.1286 ps=7.17 w=6.84 l=1.92
X8 VDD2.t6 VN.t3 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=1.1286 ps=7.17 w=6.84 l=1.92
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=0 ps=0 w=6.84 l=1.92
X10 VDD2.t5 VN.t4 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X11 VDD1.t4 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=1.1286 ps=7.17 w=6.84 l=1.92
X12 VTAIL.t9 VN.t5 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X13 VTAIL.t4 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X14 VDD2.t3 VN.t6 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=2.6676 ps=14.46 w=6.84 l=1.92
X15 VTAIL.t0 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X16 VDD2.t2 VN.t7 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=2.6676 ps=14.46 w=6.84 l=1.92
X17 VDD1.t1 VP.t8 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X18 VTAIL.t14 VN.t8 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
X19 VDD1.t0 VP.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=2.6676 ps=14.46 w=6.84 l=1.92
X20 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=0 ps=0 w=6.84 l=1.92
X21 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=0 ps=0 w=6.84 l=1.92
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.6676 pd=14.46 as=0 ps=0 w=6.84 l=1.92
X23 VTAIL.t13 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1286 pd=7.17 as=1.1286 ps=7.17 w=6.84 l=1.92
R0 VN.n59 VN.n31 161.3
R1 VN.n58 VN.n57 161.3
R2 VN.n56 VN.n32 161.3
R3 VN.n55 VN.n54 161.3
R4 VN.n52 VN.n33 161.3
R5 VN.n51 VN.n50 161.3
R6 VN.n49 VN.n34 161.3
R7 VN.n48 VN.n47 161.3
R8 VN.n46 VN.n35 161.3
R9 VN.n45 VN.n44 161.3
R10 VN.n43 VN.n36 161.3
R11 VN.n42 VN.n41 161.3
R12 VN.n40 VN.n37 161.3
R13 VN.n28 VN.n0 161.3
R14 VN.n27 VN.n26 161.3
R15 VN.n25 VN.n1 161.3
R16 VN.n24 VN.n23 161.3
R17 VN.n21 VN.n2 161.3
R18 VN.n20 VN.n19 161.3
R19 VN.n18 VN.n3 161.3
R20 VN.n17 VN.n16 161.3
R21 VN.n15 VN.n4 161.3
R22 VN.n14 VN.n13 161.3
R23 VN.n12 VN.n5 161.3
R24 VN.n11 VN.n10 161.3
R25 VN.n9 VN.n6 161.3
R26 VN.n7 VN.t3 117.356
R27 VN.n38 VN.t7 117.356
R28 VN.n30 VN.n29 86.3164
R29 VN.n61 VN.n60 86.3164
R30 VN.n29 VN.t6 85.8567
R31 VN.n15 VN.t4 85.8567
R32 VN.n8 VN.t8 85.8567
R33 VN.n22 VN.t9 85.8567
R34 VN.n60 VN.t2 85.8567
R35 VN.n46 VN.t0 85.8567
R36 VN.n39 VN.t1 85.8567
R37 VN.n53 VN.t5 85.8567
R38 VN.n8 VN.n7 58.0791
R39 VN.n39 VN.n38 58.0791
R40 VN.n10 VN.n5 52.6866
R41 VN.n20 VN.n3 52.6866
R42 VN.n27 VN.n1 52.6866
R43 VN.n41 VN.n36 52.6866
R44 VN.n51 VN.n34 52.6866
R45 VN.n58 VN.n32 52.6866
R46 VN VN.n61 45.8656
R47 VN.n14 VN.n5 28.4674
R48 VN.n16 VN.n3 28.4674
R49 VN.n28 VN.n27 28.4674
R50 VN.n45 VN.n36 28.4674
R51 VN.n47 VN.n34 28.4674
R52 VN.n59 VN.n58 28.4674
R53 VN.n10 VN.n9 24.5923
R54 VN.n15 VN.n14 24.5923
R55 VN.n16 VN.n15 24.5923
R56 VN.n21 VN.n20 24.5923
R57 VN.n23 VN.n1 24.5923
R58 VN.n29 VN.n28 24.5923
R59 VN.n41 VN.n40 24.5923
R60 VN.n47 VN.n46 24.5923
R61 VN.n46 VN.n45 24.5923
R62 VN.n54 VN.n32 24.5923
R63 VN.n52 VN.n51 24.5923
R64 VN.n60 VN.n59 24.5923
R65 VN.n38 VN.n37 12.6034
R66 VN.n7 VN.n6 12.6034
R67 VN.n9 VN.n8 12.2964
R68 VN.n22 VN.n21 12.2964
R69 VN.n23 VN.n22 12.2964
R70 VN.n40 VN.n39 12.2964
R71 VN.n54 VN.n53 12.2964
R72 VN.n53 VN.n52 12.2964
R73 VN.n61 VN.n31 0.278335
R74 VN.n30 VN.n0 0.278335
R75 VN.n57 VN.n31 0.189894
R76 VN.n57 VN.n56 0.189894
R77 VN.n56 VN.n55 0.189894
R78 VN.n55 VN.n33 0.189894
R79 VN.n50 VN.n33 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n48 0.189894
R82 VN.n48 VN.n35 0.189894
R83 VN.n44 VN.n35 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n42 0.189894
R86 VN.n42 VN.n37 0.189894
R87 VN.n11 VN.n6 0.189894
R88 VN.n12 VN.n11 0.189894
R89 VN.n13 VN.n12 0.189894
R90 VN.n13 VN.n4 0.189894
R91 VN.n17 VN.n4 0.189894
R92 VN.n18 VN.n17 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n19 VN.n2 0.189894
R95 VN.n24 VN.n2 0.189894
R96 VN.n25 VN.n24 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n26 VN.n0 0.189894
R99 VN VN.n30 0.153485
R100 VTAIL.n11 VTAIL.t16 53.5631
R101 VTAIL.n17 VTAIL.t12 53.563
R102 VTAIL.n2 VTAIL.t19 53.563
R103 VTAIL.n16 VTAIL.t7 53.563
R104 VTAIL.n15 VTAIL.n14 50.6684
R105 VTAIL.n13 VTAIL.n12 50.6684
R106 VTAIL.n10 VTAIL.n9 50.6684
R107 VTAIL.n8 VTAIL.n7 50.6684
R108 VTAIL.n19 VTAIL.n18 50.6673
R109 VTAIL.n1 VTAIL.n0 50.6673
R110 VTAIL.n4 VTAIL.n3 50.6673
R111 VTAIL.n6 VTAIL.n5 50.6673
R112 VTAIL.n8 VTAIL.n6 22.1427
R113 VTAIL.n17 VTAIL.n16 20.2031
R114 VTAIL.n18 VTAIL.t15 2.89524
R115 VTAIL.n18 VTAIL.t13 2.89524
R116 VTAIL.n0 VTAIL.t11 2.89524
R117 VTAIL.n0 VTAIL.t14 2.89524
R118 VTAIL.n3 VTAIL.t2 2.89524
R119 VTAIL.n3 VTAIL.t0 2.89524
R120 VTAIL.n5 VTAIL.t1 2.89524
R121 VTAIL.n5 VTAIL.t4 2.89524
R122 VTAIL.n14 VTAIL.t8 2.89524
R123 VTAIL.n14 VTAIL.t3 2.89524
R124 VTAIL.n12 VTAIL.t5 2.89524
R125 VTAIL.n12 VTAIL.t6 2.89524
R126 VTAIL.n9 VTAIL.t10 2.89524
R127 VTAIL.n9 VTAIL.t18 2.89524
R128 VTAIL.n7 VTAIL.t17 2.89524
R129 VTAIL.n7 VTAIL.t9 2.89524
R130 VTAIL.n10 VTAIL.n8 1.94016
R131 VTAIL.n11 VTAIL.n10 1.94016
R132 VTAIL.n15 VTAIL.n13 1.94016
R133 VTAIL.n16 VTAIL.n15 1.94016
R134 VTAIL.n6 VTAIL.n4 1.94016
R135 VTAIL.n4 VTAIL.n2 1.94016
R136 VTAIL.n19 VTAIL.n17 1.94016
R137 VTAIL VTAIL.n1 1.51343
R138 VTAIL.n13 VTAIL.n11 1.44016
R139 VTAIL.n2 VTAIL.n1 1.44016
R140 VTAIL VTAIL.n19 0.427224
R141 VDD2.n1 VDD2.t6 72.1815
R142 VDD2.n4 VDD2.t7 70.2419
R143 VDD2.n3 VDD2.n2 68.7455
R144 VDD2 VDD2.n7 68.7436
R145 VDD2.n6 VDD2.n5 67.3472
R146 VDD2.n1 VDD2.n0 67.3461
R147 VDD2.n4 VDD2.n3 38.8252
R148 VDD2.n7 VDD2.t8 2.89524
R149 VDD2.n7 VDD2.t2 2.89524
R150 VDD2.n5 VDD2.t4 2.89524
R151 VDD2.n5 VDD2.t9 2.89524
R152 VDD2.n2 VDD2.t0 2.89524
R153 VDD2.n2 VDD2.t3 2.89524
R154 VDD2.n0 VDD2.t1 2.89524
R155 VDD2.n0 VDD2.t5 2.89524
R156 VDD2.n6 VDD2.n4 1.94016
R157 VDD2 VDD2.n6 0.543603
R158 VDD2.n3 VDD2.n1 0.430068
R159 B.n706 B.n705 585
R160 B.n245 B.n120 585
R161 B.n244 B.n243 585
R162 B.n242 B.n241 585
R163 B.n240 B.n239 585
R164 B.n238 B.n237 585
R165 B.n236 B.n235 585
R166 B.n234 B.n233 585
R167 B.n232 B.n231 585
R168 B.n230 B.n229 585
R169 B.n228 B.n227 585
R170 B.n226 B.n225 585
R171 B.n224 B.n223 585
R172 B.n222 B.n221 585
R173 B.n220 B.n219 585
R174 B.n218 B.n217 585
R175 B.n216 B.n215 585
R176 B.n214 B.n213 585
R177 B.n212 B.n211 585
R178 B.n210 B.n209 585
R179 B.n208 B.n207 585
R180 B.n206 B.n205 585
R181 B.n204 B.n203 585
R182 B.n202 B.n201 585
R183 B.n200 B.n199 585
R184 B.n198 B.n197 585
R185 B.n196 B.n195 585
R186 B.n194 B.n193 585
R187 B.n192 B.n191 585
R188 B.n190 B.n189 585
R189 B.n188 B.n187 585
R190 B.n186 B.n185 585
R191 B.n184 B.n183 585
R192 B.n182 B.n181 585
R193 B.n180 B.n179 585
R194 B.n178 B.n177 585
R195 B.n176 B.n175 585
R196 B.n174 B.n173 585
R197 B.n172 B.n171 585
R198 B.n170 B.n169 585
R199 B.n168 B.n167 585
R200 B.n166 B.n165 585
R201 B.n164 B.n163 585
R202 B.n162 B.n161 585
R203 B.n160 B.n159 585
R204 B.n158 B.n157 585
R205 B.n156 B.n155 585
R206 B.n154 B.n153 585
R207 B.n152 B.n151 585
R208 B.n150 B.n149 585
R209 B.n148 B.n147 585
R210 B.n146 B.n145 585
R211 B.n144 B.n143 585
R212 B.n142 B.n141 585
R213 B.n140 B.n139 585
R214 B.n138 B.n137 585
R215 B.n136 B.n135 585
R216 B.n134 B.n133 585
R217 B.n132 B.n131 585
R218 B.n130 B.n129 585
R219 B.n128 B.n127 585
R220 B.n88 B.n87 585
R221 B.n704 B.n89 585
R222 B.n709 B.n89 585
R223 B.n703 B.n702 585
R224 B.n702 B.n85 585
R225 B.n701 B.n84 585
R226 B.n715 B.n84 585
R227 B.n700 B.n83 585
R228 B.n716 B.n83 585
R229 B.n699 B.n82 585
R230 B.n717 B.n82 585
R231 B.n698 B.n697 585
R232 B.n697 B.n78 585
R233 B.n696 B.n77 585
R234 B.n723 B.n77 585
R235 B.n695 B.n76 585
R236 B.n724 B.n76 585
R237 B.n694 B.n75 585
R238 B.n725 B.n75 585
R239 B.n693 B.n692 585
R240 B.n692 B.n71 585
R241 B.n691 B.n70 585
R242 B.n731 B.n70 585
R243 B.n690 B.n69 585
R244 B.n732 B.n69 585
R245 B.n689 B.n68 585
R246 B.n733 B.n68 585
R247 B.n688 B.n687 585
R248 B.n687 B.n64 585
R249 B.n686 B.n63 585
R250 B.n739 B.n63 585
R251 B.n685 B.n62 585
R252 B.n740 B.n62 585
R253 B.n684 B.n61 585
R254 B.n741 B.n61 585
R255 B.n683 B.n682 585
R256 B.n682 B.n57 585
R257 B.n681 B.n56 585
R258 B.n747 B.n56 585
R259 B.n680 B.n55 585
R260 B.n748 B.n55 585
R261 B.n679 B.n54 585
R262 B.n749 B.n54 585
R263 B.n678 B.n677 585
R264 B.n677 B.n50 585
R265 B.n676 B.n49 585
R266 B.n755 B.n49 585
R267 B.n675 B.n48 585
R268 B.n756 B.n48 585
R269 B.n674 B.n47 585
R270 B.n757 B.n47 585
R271 B.n673 B.n672 585
R272 B.n672 B.n43 585
R273 B.n671 B.n42 585
R274 B.n763 B.n42 585
R275 B.n670 B.n41 585
R276 B.n764 B.n41 585
R277 B.n669 B.n40 585
R278 B.n765 B.n40 585
R279 B.n668 B.n667 585
R280 B.n667 B.n39 585
R281 B.n666 B.n35 585
R282 B.n771 B.n35 585
R283 B.n665 B.n34 585
R284 B.n772 B.n34 585
R285 B.n664 B.n33 585
R286 B.n773 B.n33 585
R287 B.n663 B.n662 585
R288 B.n662 B.n29 585
R289 B.n661 B.n28 585
R290 B.n779 B.n28 585
R291 B.n660 B.n27 585
R292 B.n780 B.n27 585
R293 B.n659 B.n26 585
R294 B.n781 B.n26 585
R295 B.n658 B.n657 585
R296 B.n657 B.n22 585
R297 B.n656 B.n21 585
R298 B.n787 B.n21 585
R299 B.n655 B.n20 585
R300 B.n788 B.n20 585
R301 B.n654 B.n19 585
R302 B.n789 B.n19 585
R303 B.n653 B.n652 585
R304 B.n652 B.n15 585
R305 B.n651 B.n14 585
R306 B.n795 B.n14 585
R307 B.n650 B.n13 585
R308 B.n796 B.n13 585
R309 B.n649 B.n12 585
R310 B.n797 B.n12 585
R311 B.n648 B.n647 585
R312 B.n647 B.n8 585
R313 B.n646 B.n7 585
R314 B.n803 B.n7 585
R315 B.n645 B.n6 585
R316 B.n804 B.n6 585
R317 B.n644 B.n5 585
R318 B.n805 B.n5 585
R319 B.n643 B.n642 585
R320 B.n642 B.n4 585
R321 B.n641 B.n246 585
R322 B.n641 B.n640 585
R323 B.n631 B.n247 585
R324 B.n248 B.n247 585
R325 B.n633 B.n632 585
R326 B.n634 B.n633 585
R327 B.n630 B.n252 585
R328 B.n256 B.n252 585
R329 B.n629 B.n628 585
R330 B.n628 B.n627 585
R331 B.n254 B.n253 585
R332 B.n255 B.n254 585
R333 B.n620 B.n619 585
R334 B.n621 B.n620 585
R335 B.n618 B.n261 585
R336 B.n261 B.n260 585
R337 B.n617 B.n616 585
R338 B.n616 B.n615 585
R339 B.n263 B.n262 585
R340 B.n264 B.n263 585
R341 B.n608 B.n607 585
R342 B.n609 B.n608 585
R343 B.n606 B.n269 585
R344 B.n269 B.n268 585
R345 B.n605 B.n604 585
R346 B.n604 B.n603 585
R347 B.n271 B.n270 585
R348 B.n272 B.n271 585
R349 B.n596 B.n595 585
R350 B.n597 B.n596 585
R351 B.n594 B.n277 585
R352 B.n277 B.n276 585
R353 B.n593 B.n592 585
R354 B.n592 B.n591 585
R355 B.n279 B.n278 585
R356 B.n584 B.n279 585
R357 B.n583 B.n582 585
R358 B.n585 B.n583 585
R359 B.n581 B.n284 585
R360 B.n284 B.n283 585
R361 B.n580 B.n579 585
R362 B.n579 B.n578 585
R363 B.n286 B.n285 585
R364 B.n287 B.n286 585
R365 B.n571 B.n570 585
R366 B.n572 B.n571 585
R367 B.n569 B.n291 585
R368 B.n295 B.n291 585
R369 B.n568 B.n567 585
R370 B.n567 B.n566 585
R371 B.n293 B.n292 585
R372 B.n294 B.n293 585
R373 B.n559 B.n558 585
R374 B.n560 B.n559 585
R375 B.n557 B.n300 585
R376 B.n300 B.n299 585
R377 B.n556 B.n555 585
R378 B.n555 B.n554 585
R379 B.n302 B.n301 585
R380 B.n303 B.n302 585
R381 B.n547 B.n546 585
R382 B.n548 B.n547 585
R383 B.n545 B.n308 585
R384 B.n308 B.n307 585
R385 B.n544 B.n543 585
R386 B.n543 B.n542 585
R387 B.n310 B.n309 585
R388 B.n311 B.n310 585
R389 B.n535 B.n534 585
R390 B.n536 B.n535 585
R391 B.n533 B.n316 585
R392 B.n316 B.n315 585
R393 B.n532 B.n531 585
R394 B.n531 B.n530 585
R395 B.n318 B.n317 585
R396 B.n319 B.n318 585
R397 B.n523 B.n522 585
R398 B.n524 B.n523 585
R399 B.n521 B.n324 585
R400 B.n324 B.n323 585
R401 B.n520 B.n519 585
R402 B.n519 B.n518 585
R403 B.n326 B.n325 585
R404 B.n327 B.n326 585
R405 B.n511 B.n510 585
R406 B.n512 B.n511 585
R407 B.n509 B.n332 585
R408 B.n332 B.n331 585
R409 B.n508 B.n507 585
R410 B.n507 B.n506 585
R411 B.n334 B.n333 585
R412 B.n335 B.n334 585
R413 B.n499 B.n498 585
R414 B.n500 B.n499 585
R415 B.n338 B.n337 585
R416 B.n375 B.n373 585
R417 B.n376 B.n372 585
R418 B.n376 B.n339 585
R419 B.n379 B.n378 585
R420 B.n380 B.n371 585
R421 B.n382 B.n381 585
R422 B.n384 B.n370 585
R423 B.n387 B.n386 585
R424 B.n388 B.n369 585
R425 B.n390 B.n389 585
R426 B.n392 B.n368 585
R427 B.n395 B.n394 585
R428 B.n396 B.n367 585
R429 B.n398 B.n397 585
R430 B.n400 B.n366 585
R431 B.n403 B.n402 585
R432 B.n404 B.n365 585
R433 B.n406 B.n405 585
R434 B.n408 B.n364 585
R435 B.n411 B.n410 585
R436 B.n412 B.n363 585
R437 B.n414 B.n413 585
R438 B.n416 B.n362 585
R439 B.n419 B.n418 585
R440 B.n420 B.n361 585
R441 B.n425 B.n424 585
R442 B.n427 B.n360 585
R443 B.n430 B.n429 585
R444 B.n431 B.n359 585
R445 B.n433 B.n432 585
R446 B.n435 B.n358 585
R447 B.n438 B.n437 585
R448 B.n439 B.n357 585
R449 B.n441 B.n440 585
R450 B.n443 B.n356 585
R451 B.n446 B.n445 585
R452 B.n448 B.n353 585
R453 B.n450 B.n449 585
R454 B.n452 B.n352 585
R455 B.n455 B.n454 585
R456 B.n456 B.n351 585
R457 B.n458 B.n457 585
R458 B.n460 B.n350 585
R459 B.n463 B.n462 585
R460 B.n464 B.n349 585
R461 B.n466 B.n465 585
R462 B.n468 B.n348 585
R463 B.n471 B.n470 585
R464 B.n472 B.n347 585
R465 B.n474 B.n473 585
R466 B.n476 B.n346 585
R467 B.n479 B.n478 585
R468 B.n480 B.n345 585
R469 B.n482 B.n481 585
R470 B.n484 B.n344 585
R471 B.n487 B.n486 585
R472 B.n488 B.n343 585
R473 B.n490 B.n489 585
R474 B.n492 B.n342 585
R475 B.n493 B.n341 585
R476 B.n496 B.n495 585
R477 B.n497 B.n340 585
R478 B.n340 B.n339 585
R479 B.n502 B.n501 585
R480 B.n501 B.n500 585
R481 B.n503 B.n336 585
R482 B.n336 B.n335 585
R483 B.n505 B.n504 585
R484 B.n506 B.n505 585
R485 B.n330 B.n329 585
R486 B.n331 B.n330 585
R487 B.n514 B.n513 585
R488 B.n513 B.n512 585
R489 B.n515 B.n328 585
R490 B.n328 B.n327 585
R491 B.n517 B.n516 585
R492 B.n518 B.n517 585
R493 B.n322 B.n321 585
R494 B.n323 B.n322 585
R495 B.n526 B.n525 585
R496 B.n525 B.n524 585
R497 B.n527 B.n320 585
R498 B.n320 B.n319 585
R499 B.n529 B.n528 585
R500 B.n530 B.n529 585
R501 B.n314 B.n313 585
R502 B.n315 B.n314 585
R503 B.n538 B.n537 585
R504 B.n537 B.n536 585
R505 B.n539 B.n312 585
R506 B.n312 B.n311 585
R507 B.n541 B.n540 585
R508 B.n542 B.n541 585
R509 B.n306 B.n305 585
R510 B.n307 B.n306 585
R511 B.n550 B.n549 585
R512 B.n549 B.n548 585
R513 B.n551 B.n304 585
R514 B.n304 B.n303 585
R515 B.n553 B.n552 585
R516 B.n554 B.n553 585
R517 B.n298 B.n297 585
R518 B.n299 B.n298 585
R519 B.n562 B.n561 585
R520 B.n561 B.n560 585
R521 B.n563 B.n296 585
R522 B.n296 B.n294 585
R523 B.n565 B.n564 585
R524 B.n566 B.n565 585
R525 B.n290 B.n289 585
R526 B.n295 B.n290 585
R527 B.n574 B.n573 585
R528 B.n573 B.n572 585
R529 B.n575 B.n288 585
R530 B.n288 B.n287 585
R531 B.n577 B.n576 585
R532 B.n578 B.n577 585
R533 B.n282 B.n281 585
R534 B.n283 B.n282 585
R535 B.n587 B.n586 585
R536 B.n586 B.n585 585
R537 B.n588 B.n280 585
R538 B.n584 B.n280 585
R539 B.n590 B.n589 585
R540 B.n591 B.n590 585
R541 B.n275 B.n274 585
R542 B.n276 B.n275 585
R543 B.n599 B.n598 585
R544 B.n598 B.n597 585
R545 B.n600 B.n273 585
R546 B.n273 B.n272 585
R547 B.n602 B.n601 585
R548 B.n603 B.n602 585
R549 B.n267 B.n266 585
R550 B.n268 B.n267 585
R551 B.n611 B.n610 585
R552 B.n610 B.n609 585
R553 B.n612 B.n265 585
R554 B.n265 B.n264 585
R555 B.n614 B.n613 585
R556 B.n615 B.n614 585
R557 B.n259 B.n258 585
R558 B.n260 B.n259 585
R559 B.n623 B.n622 585
R560 B.n622 B.n621 585
R561 B.n624 B.n257 585
R562 B.n257 B.n255 585
R563 B.n626 B.n625 585
R564 B.n627 B.n626 585
R565 B.n251 B.n250 585
R566 B.n256 B.n251 585
R567 B.n636 B.n635 585
R568 B.n635 B.n634 585
R569 B.n637 B.n249 585
R570 B.n249 B.n248 585
R571 B.n639 B.n638 585
R572 B.n640 B.n639 585
R573 B.n2 B.n0 585
R574 B.n4 B.n2 585
R575 B.n3 B.n1 585
R576 B.n804 B.n3 585
R577 B.n802 B.n801 585
R578 B.n803 B.n802 585
R579 B.n800 B.n9 585
R580 B.n9 B.n8 585
R581 B.n799 B.n798 585
R582 B.n798 B.n797 585
R583 B.n11 B.n10 585
R584 B.n796 B.n11 585
R585 B.n794 B.n793 585
R586 B.n795 B.n794 585
R587 B.n792 B.n16 585
R588 B.n16 B.n15 585
R589 B.n791 B.n790 585
R590 B.n790 B.n789 585
R591 B.n18 B.n17 585
R592 B.n788 B.n18 585
R593 B.n786 B.n785 585
R594 B.n787 B.n786 585
R595 B.n784 B.n23 585
R596 B.n23 B.n22 585
R597 B.n783 B.n782 585
R598 B.n782 B.n781 585
R599 B.n25 B.n24 585
R600 B.n780 B.n25 585
R601 B.n778 B.n777 585
R602 B.n779 B.n778 585
R603 B.n776 B.n30 585
R604 B.n30 B.n29 585
R605 B.n775 B.n774 585
R606 B.n774 B.n773 585
R607 B.n32 B.n31 585
R608 B.n772 B.n32 585
R609 B.n770 B.n769 585
R610 B.n771 B.n770 585
R611 B.n768 B.n36 585
R612 B.n39 B.n36 585
R613 B.n767 B.n766 585
R614 B.n766 B.n765 585
R615 B.n38 B.n37 585
R616 B.n764 B.n38 585
R617 B.n762 B.n761 585
R618 B.n763 B.n762 585
R619 B.n760 B.n44 585
R620 B.n44 B.n43 585
R621 B.n759 B.n758 585
R622 B.n758 B.n757 585
R623 B.n46 B.n45 585
R624 B.n756 B.n46 585
R625 B.n754 B.n753 585
R626 B.n755 B.n754 585
R627 B.n752 B.n51 585
R628 B.n51 B.n50 585
R629 B.n751 B.n750 585
R630 B.n750 B.n749 585
R631 B.n53 B.n52 585
R632 B.n748 B.n53 585
R633 B.n746 B.n745 585
R634 B.n747 B.n746 585
R635 B.n744 B.n58 585
R636 B.n58 B.n57 585
R637 B.n743 B.n742 585
R638 B.n742 B.n741 585
R639 B.n60 B.n59 585
R640 B.n740 B.n60 585
R641 B.n738 B.n737 585
R642 B.n739 B.n738 585
R643 B.n736 B.n65 585
R644 B.n65 B.n64 585
R645 B.n735 B.n734 585
R646 B.n734 B.n733 585
R647 B.n67 B.n66 585
R648 B.n732 B.n67 585
R649 B.n730 B.n729 585
R650 B.n731 B.n730 585
R651 B.n728 B.n72 585
R652 B.n72 B.n71 585
R653 B.n727 B.n726 585
R654 B.n726 B.n725 585
R655 B.n74 B.n73 585
R656 B.n724 B.n74 585
R657 B.n722 B.n721 585
R658 B.n723 B.n722 585
R659 B.n720 B.n79 585
R660 B.n79 B.n78 585
R661 B.n719 B.n718 585
R662 B.n718 B.n717 585
R663 B.n81 B.n80 585
R664 B.n716 B.n81 585
R665 B.n714 B.n713 585
R666 B.n715 B.n714 585
R667 B.n712 B.n86 585
R668 B.n86 B.n85 585
R669 B.n711 B.n710 585
R670 B.n710 B.n709 585
R671 B.n807 B.n806 585
R672 B.n806 B.n805 585
R673 B.n501 B.n338 506.916
R674 B.n710 B.n88 506.916
R675 B.n499 B.n340 506.916
R676 B.n706 B.n89 506.916
R677 B.n354 B.t14 292.579
R678 B.n421 B.t21 292.579
R679 B.n124 B.t18 292.579
R680 B.n121 B.t10 292.579
R681 B.n708 B.n707 256.663
R682 B.n708 B.n119 256.663
R683 B.n708 B.n118 256.663
R684 B.n708 B.n117 256.663
R685 B.n708 B.n116 256.663
R686 B.n708 B.n115 256.663
R687 B.n708 B.n114 256.663
R688 B.n708 B.n113 256.663
R689 B.n708 B.n112 256.663
R690 B.n708 B.n111 256.663
R691 B.n708 B.n110 256.663
R692 B.n708 B.n109 256.663
R693 B.n708 B.n108 256.663
R694 B.n708 B.n107 256.663
R695 B.n708 B.n106 256.663
R696 B.n708 B.n105 256.663
R697 B.n708 B.n104 256.663
R698 B.n708 B.n103 256.663
R699 B.n708 B.n102 256.663
R700 B.n708 B.n101 256.663
R701 B.n708 B.n100 256.663
R702 B.n708 B.n99 256.663
R703 B.n708 B.n98 256.663
R704 B.n708 B.n97 256.663
R705 B.n708 B.n96 256.663
R706 B.n708 B.n95 256.663
R707 B.n708 B.n94 256.663
R708 B.n708 B.n93 256.663
R709 B.n708 B.n92 256.663
R710 B.n708 B.n91 256.663
R711 B.n708 B.n90 256.663
R712 B.n374 B.n339 256.663
R713 B.n377 B.n339 256.663
R714 B.n383 B.n339 256.663
R715 B.n385 B.n339 256.663
R716 B.n391 B.n339 256.663
R717 B.n393 B.n339 256.663
R718 B.n399 B.n339 256.663
R719 B.n401 B.n339 256.663
R720 B.n407 B.n339 256.663
R721 B.n409 B.n339 256.663
R722 B.n415 B.n339 256.663
R723 B.n417 B.n339 256.663
R724 B.n426 B.n339 256.663
R725 B.n428 B.n339 256.663
R726 B.n434 B.n339 256.663
R727 B.n436 B.n339 256.663
R728 B.n442 B.n339 256.663
R729 B.n444 B.n339 256.663
R730 B.n451 B.n339 256.663
R731 B.n453 B.n339 256.663
R732 B.n459 B.n339 256.663
R733 B.n461 B.n339 256.663
R734 B.n467 B.n339 256.663
R735 B.n469 B.n339 256.663
R736 B.n475 B.n339 256.663
R737 B.n477 B.n339 256.663
R738 B.n483 B.n339 256.663
R739 B.n485 B.n339 256.663
R740 B.n491 B.n339 256.663
R741 B.n494 B.n339 256.663
R742 B.n501 B.n336 163.367
R743 B.n505 B.n336 163.367
R744 B.n505 B.n330 163.367
R745 B.n513 B.n330 163.367
R746 B.n513 B.n328 163.367
R747 B.n517 B.n328 163.367
R748 B.n517 B.n322 163.367
R749 B.n525 B.n322 163.367
R750 B.n525 B.n320 163.367
R751 B.n529 B.n320 163.367
R752 B.n529 B.n314 163.367
R753 B.n537 B.n314 163.367
R754 B.n537 B.n312 163.367
R755 B.n541 B.n312 163.367
R756 B.n541 B.n306 163.367
R757 B.n549 B.n306 163.367
R758 B.n549 B.n304 163.367
R759 B.n553 B.n304 163.367
R760 B.n553 B.n298 163.367
R761 B.n561 B.n298 163.367
R762 B.n561 B.n296 163.367
R763 B.n565 B.n296 163.367
R764 B.n565 B.n290 163.367
R765 B.n573 B.n290 163.367
R766 B.n573 B.n288 163.367
R767 B.n577 B.n288 163.367
R768 B.n577 B.n282 163.367
R769 B.n586 B.n282 163.367
R770 B.n586 B.n280 163.367
R771 B.n590 B.n280 163.367
R772 B.n590 B.n275 163.367
R773 B.n598 B.n275 163.367
R774 B.n598 B.n273 163.367
R775 B.n602 B.n273 163.367
R776 B.n602 B.n267 163.367
R777 B.n610 B.n267 163.367
R778 B.n610 B.n265 163.367
R779 B.n614 B.n265 163.367
R780 B.n614 B.n259 163.367
R781 B.n622 B.n259 163.367
R782 B.n622 B.n257 163.367
R783 B.n626 B.n257 163.367
R784 B.n626 B.n251 163.367
R785 B.n635 B.n251 163.367
R786 B.n635 B.n249 163.367
R787 B.n639 B.n249 163.367
R788 B.n639 B.n2 163.367
R789 B.n806 B.n2 163.367
R790 B.n806 B.n3 163.367
R791 B.n802 B.n3 163.367
R792 B.n802 B.n9 163.367
R793 B.n798 B.n9 163.367
R794 B.n798 B.n11 163.367
R795 B.n794 B.n11 163.367
R796 B.n794 B.n16 163.367
R797 B.n790 B.n16 163.367
R798 B.n790 B.n18 163.367
R799 B.n786 B.n18 163.367
R800 B.n786 B.n23 163.367
R801 B.n782 B.n23 163.367
R802 B.n782 B.n25 163.367
R803 B.n778 B.n25 163.367
R804 B.n778 B.n30 163.367
R805 B.n774 B.n30 163.367
R806 B.n774 B.n32 163.367
R807 B.n770 B.n32 163.367
R808 B.n770 B.n36 163.367
R809 B.n766 B.n36 163.367
R810 B.n766 B.n38 163.367
R811 B.n762 B.n38 163.367
R812 B.n762 B.n44 163.367
R813 B.n758 B.n44 163.367
R814 B.n758 B.n46 163.367
R815 B.n754 B.n46 163.367
R816 B.n754 B.n51 163.367
R817 B.n750 B.n51 163.367
R818 B.n750 B.n53 163.367
R819 B.n746 B.n53 163.367
R820 B.n746 B.n58 163.367
R821 B.n742 B.n58 163.367
R822 B.n742 B.n60 163.367
R823 B.n738 B.n60 163.367
R824 B.n738 B.n65 163.367
R825 B.n734 B.n65 163.367
R826 B.n734 B.n67 163.367
R827 B.n730 B.n67 163.367
R828 B.n730 B.n72 163.367
R829 B.n726 B.n72 163.367
R830 B.n726 B.n74 163.367
R831 B.n722 B.n74 163.367
R832 B.n722 B.n79 163.367
R833 B.n718 B.n79 163.367
R834 B.n718 B.n81 163.367
R835 B.n714 B.n81 163.367
R836 B.n714 B.n86 163.367
R837 B.n710 B.n86 163.367
R838 B.n376 B.n375 163.367
R839 B.n378 B.n376 163.367
R840 B.n382 B.n371 163.367
R841 B.n386 B.n384 163.367
R842 B.n390 B.n369 163.367
R843 B.n394 B.n392 163.367
R844 B.n398 B.n367 163.367
R845 B.n402 B.n400 163.367
R846 B.n406 B.n365 163.367
R847 B.n410 B.n408 163.367
R848 B.n414 B.n363 163.367
R849 B.n418 B.n416 163.367
R850 B.n425 B.n361 163.367
R851 B.n429 B.n427 163.367
R852 B.n433 B.n359 163.367
R853 B.n437 B.n435 163.367
R854 B.n441 B.n357 163.367
R855 B.n445 B.n443 163.367
R856 B.n450 B.n353 163.367
R857 B.n454 B.n452 163.367
R858 B.n458 B.n351 163.367
R859 B.n462 B.n460 163.367
R860 B.n466 B.n349 163.367
R861 B.n470 B.n468 163.367
R862 B.n474 B.n347 163.367
R863 B.n478 B.n476 163.367
R864 B.n482 B.n345 163.367
R865 B.n486 B.n484 163.367
R866 B.n490 B.n343 163.367
R867 B.n493 B.n492 163.367
R868 B.n495 B.n340 163.367
R869 B.n499 B.n334 163.367
R870 B.n507 B.n334 163.367
R871 B.n507 B.n332 163.367
R872 B.n511 B.n332 163.367
R873 B.n511 B.n326 163.367
R874 B.n519 B.n326 163.367
R875 B.n519 B.n324 163.367
R876 B.n523 B.n324 163.367
R877 B.n523 B.n318 163.367
R878 B.n531 B.n318 163.367
R879 B.n531 B.n316 163.367
R880 B.n535 B.n316 163.367
R881 B.n535 B.n310 163.367
R882 B.n543 B.n310 163.367
R883 B.n543 B.n308 163.367
R884 B.n547 B.n308 163.367
R885 B.n547 B.n302 163.367
R886 B.n555 B.n302 163.367
R887 B.n555 B.n300 163.367
R888 B.n559 B.n300 163.367
R889 B.n559 B.n293 163.367
R890 B.n567 B.n293 163.367
R891 B.n567 B.n291 163.367
R892 B.n571 B.n291 163.367
R893 B.n571 B.n286 163.367
R894 B.n579 B.n286 163.367
R895 B.n579 B.n284 163.367
R896 B.n583 B.n284 163.367
R897 B.n583 B.n279 163.367
R898 B.n592 B.n279 163.367
R899 B.n592 B.n277 163.367
R900 B.n596 B.n277 163.367
R901 B.n596 B.n271 163.367
R902 B.n604 B.n271 163.367
R903 B.n604 B.n269 163.367
R904 B.n608 B.n269 163.367
R905 B.n608 B.n263 163.367
R906 B.n616 B.n263 163.367
R907 B.n616 B.n261 163.367
R908 B.n620 B.n261 163.367
R909 B.n620 B.n254 163.367
R910 B.n628 B.n254 163.367
R911 B.n628 B.n252 163.367
R912 B.n633 B.n252 163.367
R913 B.n633 B.n247 163.367
R914 B.n641 B.n247 163.367
R915 B.n642 B.n641 163.367
R916 B.n642 B.n5 163.367
R917 B.n6 B.n5 163.367
R918 B.n7 B.n6 163.367
R919 B.n647 B.n7 163.367
R920 B.n647 B.n12 163.367
R921 B.n13 B.n12 163.367
R922 B.n14 B.n13 163.367
R923 B.n652 B.n14 163.367
R924 B.n652 B.n19 163.367
R925 B.n20 B.n19 163.367
R926 B.n21 B.n20 163.367
R927 B.n657 B.n21 163.367
R928 B.n657 B.n26 163.367
R929 B.n27 B.n26 163.367
R930 B.n28 B.n27 163.367
R931 B.n662 B.n28 163.367
R932 B.n662 B.n33 163.367
R933 B.n34 B.n33 163.367
R934 B.n35 B.n34 163.367
R935 B.n667 B.n35 163.367
R936 B.n667 B.n40 163.367
R937 B.n41 B.n40 163.367
R938 B.n42 B.n41 163.367
R939 B.n672 B.n42 163.367
R940 B.n672 B.n47 163.367
R941 B.n48 B.n47 163.367
R942 B.n49 B.n48 163.367
R943 B.n677 B.n49 163.367
R944 B.n677 B.n54 163.367
R945 B.n55 B.n54 163.367
R946 B.n56 B.n55 163.367
R947 B.n682 B.n56 163.367
R948 B.n682 B.n61 163.367
R949 B.n62 B.n61 163.367
R950 B.n63 B.n62 163.367
R951 B.n687 B.n63 163.367
R952 B.n687 B.n68 163.367
R953 B.n69 B.n68 163.367
R954 B.n70 B.n69 163.367
R955 B.n692 B.n70 163.367
R956 B.n692 B.n75 163.367
R957 B.n76 B.n75 163.367
R958 B.n77 B.n76 163.367
R959 B.n697 B.n77 163.367
R960 B.n697 B.n82 163.367
R961 B.n83 B.n82 163.367
R962 B.n84 B.n83 163.367
R963 B.n702 B.n84 163.367
R964 B.n702 B.n89 163.367
R965 B.n129 B.n128 163.367
R966 B.n133 B.n132 163.367
R967 B.n137 B.n136 163.367
R968 B.n141 B.n140 163.367
R969 B.n145 B.n144 163.367
R970 B.n149 B.n148 163.367
R971 B.n153 B.n152 163.367
R972 B.n157 B.n156 163.367
R973 B.n161 B.n160 163.367
R974 B.n165 B.n164 163.367
R975 B.n169 B.n168 163.367
R976 B.n173 B.n172 163.367
R977 B.n177 B.n176 163.367
R978 B.n181 B.n180 163.367
R979 B.n185 B.n184 163.367
R980 B.n189 B.n188 163.367
R981 B.n193 B.n192 163.367
R982 B.n197 B.n196 163.367
R983 B.n201 B.n200 163.367
R984 B.n205 B.n204 163.367
R985 B.n209 B.n208 163.367
R986 B.n213 B.n212 163.367
R987 B.n217 B.n216 163.367
R988 B.n221 B.n220 163.367
R989 B.n225 B.n224 163.367
R990 B.n229 B.n228 163.367
R991 B.n233 B.n232 163.367
R992 B.n237 B.n236 163.367
R993 B.n241 B.n240 163.367
R994 B.n243 B.n120 163.367
R995 B.n354 B.t17 113.444
R996 B.n121 B.t12 113.444
R997 B.n421 B.t23 113.436
R998 B.n124 B.t19 113.436
R999 B.n500 B.n339 100.784
R1000 B.n709 B.n708 100.784
R1001 B.n374 B.n338 71.676
R1002 B.n378 B.n377 71.676
R1003 B.n383 B.n382 71.676
R1004 B.n386 B.n385 71.676
R1005 B.n391 B.n390 71.676
R1006 B.n394 B.n393 71.676
R1007 B.n399 B.n398 71.676
R1008 B.n402 B.n401 71.676
R1009 B.n407 B.n406 71.676
R1010 B.n410 B.n409 71.676
R1011 B.n415 B.n414 71.676
R1012 B.n418 B.n417 71.676
R1013 B.n426 B.n425 71.676
R1014 B.n429 B.n428 71.676
R1015 B.n434 B.n433 71.676
R1016 B.n437 B.n436 71.676
R1017 B.n442 B.n441 71.676
R1018 B.n445 B.n444 71.676
R1019 B.n451 B.n450 71.676
R1020 B.n454 B.n453 71.676
R1021 B.n459 B.n458 71.676
R1022 B.n462 B.n461 71.676
R1023 B.n467 B.n466 71.676
R1024 B.n470 B.n469 71.676
R1025 B.n475 B.n474 71.676
R1026 B.n478 B.n477 71.676
R1027 B.n483 B.n482 71.676
R1028 B.n486 B.n485 71.676
R1029 B.n491 B.n490 71.676
R1030 B.n494 B.n493 71.676
R1031 B.n90 B.n88 71.676
R1032 B.n129 B.n91 71.676
R1033 B.n133 B.n92 71.676
R1034 B.n137 B.n93 71.676
R1035 B.n141 B.n94 71.676
R1036 B.n145 B.n95 71.676
R1037 B.n149 B.n96 71.676
R1038 B.n153 B.n97 71.676
R1039 B.n157 B.n98 71.676
R1040 B.n161 B.n99 71.676
R1041 B.n165 B.n100 71.676
R1042 B.n169 B.n101 71.676
R1043 B.n173 B.n102 71.676
R1044 B.n177 B.n103 71.676
R1045 B.n181 B.n104 71.676
R1046 B.n185 B.n105 71.676
R1047 B.n189 B.n106 71.676
R1048 B.n193 B.n107 71.676
R1049 B.n197 B.n108 71.676
R1050 B.n201 B.n109 71.676
R1051 B.n205 B.n110 71.676
R1052 B.n209 B.n111 71.676
R1053 B.n213 B.n112 71.676
R1054 B.n217 B.n113 71.676
R1055 B.n221 B.n114 71.676
R1056 B.n225 B.n115 71.676
R1057 B.n229 B.n116 71.676
R1058 B.n233 B.n117 71.676
R1059 B.n237 B.n118 71.676
R1060 B.n241 B.n119 71.676
R1061 B.n707 B.n120 71.676
R1062 B.n707 B.n706 71.676
R1063 B.n243 B.n119 71.676
R1064 B.n240 B.n118 71.676
R1065 B.n236 B.n117 71.676
R1066 B.n232 B.n116 71.676
R1067 B.n228 B.n115 71.676
R1068 B.n224 B.n114 71.676
R1069 B.n220 B.n113 71.676
R1070 B.n216 B.n112 71.676
R1071 B.n212 B.n111 71.676
R1072 B.n208 B.n110 71.676
R1073 B.n204 B.n109 71.676
R1074 B.n200 B.n108 71.676
R1075 B.n196 B.n107 71.676
R1076 B.n192 B.n106 71.676
R1077 B.n188 B.n105 71.676
R1078 B.n184 B.n104 71.676
R1079 B.n180 B.n103 71.676
R1080 B.n176 B.n102 71.676
R1081 B.n172 B.n101 71.676
R1082 B.n168 B.n100 71.676
R1083 B.n164 B.n99 71.676
R1084 B.n160 B.n98 71.676
R1085 B.n156 B.n97 71.676
R1086 B.n152 B.n96 71.676
R1087 B.n148 B.n95 71.676
R1088 B.n144 B.n94 71.676
R1089 B.n140 B.n93 71.676
R1090 B.n136 B.n92 71.676
R1091 B.n132 B.n91 71.676
R1092 B.n128 B.n90 71.676
R1093 B.n375 B.n374 71.676
R1094 B.n377 B.n371 71.676
R1095 B.n384 B.n383 71.676
R1096 B.n385 B.n369 71.676
R1097 B.n392 B.n391 71.676
R1098 B.n393 B.n367 71.676
R1099 B.n400 B.n399 71.676
R1100 B.n401 B.n365 71.676
R1101 B.n408 B.n407 71.676
R1102 B.n409 B.n363 71.676
R1103 B.n416 B.n415 71.676
R1104 B.n417 B.n361 71.676
R1105 B.n427 B.n426 71.676
R1106 B.n428 B.n359 71.676
R1107 B.n435 B.n434 71.676
R1108 B.n436 B.n357 71.676
R1109 B.n443 B.n442 71.676
R1110 B.n444 B.n353 71.676
R1111 B.n452 B.n451 71.676
R1112 B.n453 B.n351 71.676
R1113 B.n460 B.n459 71.676
R1114 B.n461 B.n349 71.676
R1115 B.n468 B.n467 71.676
R1116 B.n469 B.n347 71.676
R1117 B.n476 B.n475 71.676
R1118 B.n477 B.n345 71.676
R1119 B.n484 B.n483 71.676
R1120 B.n485 B.n343 71.676
R1121 B.n492 B.n491 71.676
R1122 B.n495 B.n494 71.676
R1123 B.n355 B.t16 69.8069
R1124 B.n122 B.t13 69.8069
R1125 B.n422 B.t22 69.7992
R1126 B.n125 B.t20 69.7992
R1127 B.n500 B.n335 61.7421
R1128 B.n506 B.n335 61.7421
R1129 B.n506 B.n331 61.7421
R1130 B.n512 B.n331 61.7421
R1131 B.n512 B.n327 61.7421
R1132 B.n518 B.n327 61.7421
R1133 B.n524 B.n323 61.7421
R1134 B.n524 B.n319 61.7421
R1135 B.n530 B.n319 61.7421
R1136 B.n530 B.n315 61.7421
R1137 B.n536 B.n315 61.7421
R1138 B.n536 B.n311 61.7421
R1139 B.n542 B.n311 61.7421
R1140 B.n542 B.n307 61.7421
R1141 B.n548 B.n307 61.7421
R1142 B.n554 B.n303 61.7421
R1143 B.n554 B.n299 61.7421
R1144 B.n560 B.n299 61.7421
R1145 B.n560 B.n294 61.7421
R1146 B.n566 B.n294 61.7421
R1147 B.n566 B.n295 61.7421
R1148 B.n572 B.n287 61.7421
R1149 B.n578 B.n287 61.7421
R1150 B.n578 B.n283 61.7421
R1151 B.n585 B.n283 61.7421
R1152 B.n585 B.n584 61.7421
R1153 B.n591 B.n276 61.7421
R1154 B.n597 B.n276 61.7421
R1155 B.n597 B.n272 61.7421
R1156 B.n603 B.n272 61.7421
R1157 B.n603 B.n268 61.7421
R1158 B.n609 B.n268 61.7421
R1159 B.n615 B.n264 61.7421
R1160 B.n615 B.n260 61.7421
R1161 B.n621 B.n260 61.7421
R1162 B.n621 B.n255 61.7421
R1163 B.n627 B.n255 61.7421
R1164 B.n627 B.n256 61.7421
R1165 B.n634 B.n248 61.7421
R1166 B.n640 B.n248 61.7421
R1167 B.n640 B.n4 61.7421
R1168 B.n805 B.n4 61.7421
R1169 B.n805 B.n804 61.7421
R1170 B.n804 B.n803 61.7421
R1171 B.n803 B.n8 61.7421
R1172 B.n797 B.n8 61.7421
R1173 B.n796 B.n795 61.7421
R1174 B.n795 B.n15 61.7421
R1175 B.n789 B.n15 61.7421
R1176 B.n789 B.n788 61.7421
R1177 B.n788 B.n787 61.7421
R1178 B.n787 B.n22 61.7421
R1179 B.n781 B.n780 61.7421
R1180 B.n780 B.n779 61.7421
R1181 B.n779 B.n29 61.7421
R1182 B.n773 B.n29 61.7421
R1183 B.n773 B.n772 61.7421
R1184 B.n772 B.n771 61.7421
R1185 B.n765 B.n39 61.7421
R1186 B.n765 B.n764 61.7421
R1187 B.n764 B.n763 61.7421
R1188 B.n763 B.n43 61.7421
R1189 B.n757 B.n43 61.7421
R1190 B.n756 B.n755 61.7421
R1191 B.n755 B.n50 61.7421
R1192 B.n749 B.n50 61.7421
R1193 B.n749 B.n748 61.7421
R1194 B.n748 B.n747 61.7421
R1195 B.n747 B.n57 61.7421
R1196 B.n741 B.n740 61.7421
R1197 B.n740 B.n739 61.7421
R1198 B.n739 B.n64 61.7421
R1199 B.n733 B.n64 61.7421
R1200 B.n733 B.n732 61.7421
R1201 B.n732 B.n731 61.7421
R1202 B.n731 B.n71 61.7421
R1203 B.n725 B.n71 61.7421
R1204 B.n725 B.n724 61.7421
R1205 B.n723 B.n78 61.7421
R1206 B.n717 B.n78 61.7421
R1207 B.n717 B.n716 61.7421
R1208 B.n716 B.n715 61.7421
R1209 B.n715 B.n85 61.7421
R1210 B.n709 B.n85 61.7421
R1211 B.n447 B.n355 59.5399
R1212 B.n423 B.n422 59.5399
R1213 B.n126 B.n125 59.5399
R1214 B.n123 B.n122 59.5399
R1215 B.n634 B.t9 56.2943
R1216 B.n797 B.t5 56.2943
R1217 B.n584 B.t2 52.6625
R1218 B.n39 B.t8 52.6625
R1219 B.n518 B.t15 49.0306
R1220 B.t11 B.n723 49.0306
R1221 B.n572 B.t4 47.2147
R1222 B.n757 B.t3 47.2147
R1223 B.n355 B.n354 43.6369
R1224 B.n422 B.n421 43.6369
R1225 B.n125 B.n124 43.6369
R1226 B.n122 B.n121 43.6369
R1227 B.n548 B.t1 38.135
R1228 B.n741 B.t7 38.135
R1229 B.n711 B.n87 32.9371
R1230 B.n705 B.n704 32.9371
R1231 B.n498 B.n497 32.9371
R1232 B.n502 B.n337 32.9371
R1233 B.t0 B.n264 32.6873
R1234 B.t6 B.n22 32.6873
R1235 B.n609 B.t0 29.0554
R1236 B.n781 B.t6 29.0554
R1237 B.t1 B.n303 23.6076
R1238 B.t7 B.n57 23.6076
R1239 B B.n807 18.0485
R1240 B.n295 B.t4 14.5279
R1241 B.t3 B.n756 14.5279
R1242 B.t15 B.n323 12.712
R1243 B.n724 B.t11 12.712
R1244 B.n127 B.n87 10.6151
R1245 B.n130 B.n127 10.6151
R1246 B.n131 B.n130 10.6151
R1247 B.n134 B.n131 10.6151
R1248 B.n135 B.n134 10.6151
R1249 B.n138 B.n135 10.6151
R1250 B.n139 B.n138 10.6151
R1251 B.n142 B.n139 10.6151
R1252 B.n143 B.n142 10.6151
R1253 B.n146 B.n143 10.6151
R1254 B.n147 B.n146 10.6151
R1255 B.n150 B.n147 10.6151
R1256 B.n151 B.n150 10.6151
R1257 B.n154 B.n151 10.6151
R1258 B.n155 B.n154 10.6151
R1259 B.n158 B.n155 10.6151
R1260 B.n159 B.n158 10.6151
R1261 B.n162 B.n159 10.6151
R1262 B.n163 B.n162 10.6151
R1263 B.n166 B.n163 10.6151
R1264 B.n167 B.n166 10.6151
R1265 B.n170 B.n167 10.6151
R1266 B.n171 B.n170 10.6151
R1267 B.n174 B.n171 10.6151
R1268 B.n175 B.n174 10.6151
R1269 B.n179 B.n178 10.6151
R1270 B.n182 B.n179 10.6151
R1271 B.n183 B.n182 10.6151
R1272 B.n186 B.n183 10.6151
R1273 B.n187 B.n186 10.6151
R1274 B.n190 B.n187 10.6151
R1275 B.n191 B.n190 10.6151
R1276 B.n194 B.n191 10.6151
R1277 B.n195 B.n194 10.6151
R1278 B.n199 B.n198 10.6151
R1279 B.n202 B.n199 10.6151
R1280 B.n203 B.n202 10.6151
R1281 B.n206 B.n203 10.6151
R1282 B.n207 B.n206 10.6151
R1283 B.n210 B.n207 10.6151
R1284 B.n211 B.n210 10.6151
R1285 B.n214 B.n211 10.6151
R1286 B.n215 B.n214 10.6151
R1287 B.n218 B.n215 10.6151
R1288 B.n219 B.n218 10.6151
R1289 B.n222 B.n219 10.6151
R1290 B.n223 B.n222 10.6151
R1291 B.n226 B.n223 10.6151
R1292 B.n227 B.n226 10.6151
R1293 B.n230 B.n227 10.6151
R1294 B.n231 B.n230 10.6151
R1295 B.n234 B.n231 10.6151
R1296 B.n235 B.n234 10.6151
R1297 B.n238 B.n235 10.6151
R1298 B.n239 B.n238 10.6151
R1299 B.n242 B.n239 10.6151
R1300 B.n244 B.n242 10.6151
R1301 B.n245 B.n244 10.6151
R1302 B.n705 B.n245 10.6151
R1303 B.n498 B.n333 10.6151
R1304 B.n508 B.n333 10.6151
R1305 B.n509 B.n508 10.6151
R1306 B.n510 B.n509 10.6151
R1307 B.n510 B.n325 10.6151
R1308 B.n520 B.n325 10.6151
R1309 B.n521 B.n520 10.6151
R1310 B.n522 B.n521 10.6151
R1311 B.n522 B.n317 10.6151
R1312 B.n532 B.n317 10.6151
R1313 B.n533 B.n532 10.6151
R1314 B.n534 B.n533 10.6151
R1315 B.n534 B.n309 10.6151
R1316 B.n544 B.n309 10.6151
R1317 B.n545 B.n544 10.6151
R1318 B.n546 B.n545 10.6151
R1319 B.n546 B.n301 10.6151
R1320 B.n556 B.n301 10.6151
R1321 B.n557 B.n556 10.6151
R1322 B.n558 B.n557 10.6151
R1323 B.n558 B.n292 10.6151
R1324 B.n568 B.n292 10.6151
R1325 B.n569 B.n568 10.6151
R1326 B.n570 B.n569 10.6151
R1327 B.n570 B.n285 10.6151
R1328 B.n580 B.n285 10.6151
R1329 B.n581 B.n580 10.6151
R1330 B.n582 B.n581 10.6151
R1331 B.n582 B.n278 10.6151
R1332 B.n593 B.n278 10.6151
R1333 B.n594 B.n593 10.6151
R1334 B.n595 B.n594 10.6151
R1335 B.n595 B.n270 10.6151
R1336 B.n605 B.n270 10.6151
R1337 B.n606 B.n605 10.6151
R1338 B.n607 B.n606 10.6151
R1339 B.n607 B.n262 10.6151
R1340 B.n617 B.n262 10.6151
R1341 B.n618 B.n617 10.6151
R1342 B.n619 B.n618 10.6151
R1343 B.n619 B.n253 10.6151
R1344 B.n629 B.n253 10.6151
R1345 B.n630 B.n629 10.6151
R1346 B.n632 B.n630 10.6151
R1347 B.n632 B.n631 10.6151
R1348 B.n631 B.n246 10.6151
R1349 B.n643 B.n246 10.6151
R1350 B.n644 B.n643 10.6151
R1351 B.n645 B.n644 10.6151
R1352 B.n646 B.n645 10.6151
R1353 B.n648 B.n646 10.6151
R1354 B.n649 B.n648 10.6151
R1355 B.n650 B.n649 10.6151
R1356 B.n651 B.n650 10.6151
R1357 B.n653 B.n651 10.6151
R1358 B.n654 B.n653 10.6151
R1359 B.n655 B.n654 10.6151
R1360 B.n656 B.n655 10.6151
R1361 B.n658 B.n656 10.6151
R1362 B.n659 B.n658 10.6151
R1363 B.n660 B.n659 10.6151
R1364 B.n661 B.n660 10.6151
R1365 B.n663 B.n661 10.6151
R1366 B.n664 B.n663 10.6151
R1367 B.n665 B.n664 10.6151
R1368 B.n666 B.n665 10.6151
R1369 B.n668 B.n666 10.6151
R1370 B.n669 B.n668 10.6151
R1371 B.n670 B.n669 10.6151
R1372 B.n671 B.n670 10.6151
R1373 B.n673 B.n671 10.6151
R1374 B.n674 B.n673 10.6151
R1375 B.n675 B.n674 10.6151
R1376 B.n676 B.n675 10.6151
R1377 B.n678 B.n676 10.6151
R1378 B.n679 B.n678 10.6151
R1379 B.n680 B.n679 10.6151
R1380 B.n681 B.n680 10.6151
R1381 B.n683 B.n681 10.6151
R1382 B.n684 B.n683 10.6151
R1383 B.n685 B.n684 10.6151
R1384 B.n686 B.n685 10.6151
R1385 B.n688 B.n686 10.6151
R1386 B.n689 B.n688 10.6151
R1387 B.n690 B.n689 10.6151
R1388 B.n691 B.n690 10.6151
R1389 B.n693 B.n691 10.6151
R1390 B.n694 B.n693 10.6151
R1391 B.n695 B.n694 10.6151
R1392 B.n696 B.n695 10.6151
R1393 B.n698 B.n696 10.6151
R1394 B.n699 B.n698 10.6151
R1395 B.n700 B.n699 10.6151
R1396 B.n701 B.n700 10.6151
R1397 B.n703 B.n701 10.6151
R1398 B.n704 B.n703 10.6151
R1399 B.n373 B.n337 10.6151
R1400 B.n373 B.n372 10.6151
R1401 B.n379 B.n372 10.6151
R1402 B.n380 B.n379 10.6151
R1403 B.n381 B.n380 10.6151
R1404 B.n381 B.n370 10.6151
R1405 B.n387 B.n370 10.6151
R1406 B.n388 B.n387 10.6151
R1407 B.n389 B.n388 10.6151
R1408 B.n389 B.n368 10.6151
R1409 B.n395 B.n368 10.6151
R1410 B.n396 B.n395 10.6151
R1411 B.n397 B.n396 10.6151
R1412 B.n397 B.n366 10.6151
R1413 B.n403 B.n366 10.6151
R1414 B.n404 B.n403 10.6151
R1415 B.n405 B.n404 10.6151
R1416 B.n405 B.n364 10.6151
R1417 B.n411 B.n364 10.6151
R1418 B.n412 B.n411 10.6151
R1419 B.n413 B.n412 10.6151
R1420 B.n413 B.n362 10.6151
R1421 B.n419 B.n362 10.6151
R1422 B.n420 B.n419 10.6151
R1423 B.n424 B.n420 10.6151
R1424 B.n430 B.n360 10.6151
R1425 B.n431 B.n430 10.6151
R1426 B.n432 B.n431 10.6151
R1427 B.n432 B.n358 10.6151
R1428 B.n438 B.n358 10.6151
R1429 B.n439 B.n438 10.6151
R1430 B.n440 B.n439 10.6151
R1431 B.n440 B.n356 10.6151
R1432 B.n446 B.n356 10.6151
R1433 B.n449 B.n448 10.6151
R1434 B.n449 B.n352 10.6151
R1435 B.n455 B.n352 10.6151
R1436 B.n456 B.n455 10.6151
R1437 B.n457 B.n456 10.6151
R1438 B.n457 B.n350 10.6151
R1439 B.n463 B.n350 10.6151
R1440 B.n464 B.n463 10.6151
R1441 B.n465 B.n464 10.6151
R1442 B.n465 B.n348 10.6151
R1443 B.n471 B.n348 10.6151
R1444 B.n472 B.n471 10.6151
R1445 B.n473 B.n472 10.6151
R1446 B.n473 B.n346 10.6151
R1447 B.n479 B.n346 10.6151
R1448 B.n480 B.n479 10.6151
R1449 B.n481 B.n480 10.6151
R1450 B.n481 B.n344 10.6151
R1451 B.n487 B.n344 10.6151
R1452 B.n488 B.n487 10.6151
R1453 B.n489 B.n488 10.6151
R1454 B.n489 B.n342 10.6151
R1455 B.n342 B.n341 10.6151
R1456 B.n496 B.n341 10.6151
R1457 B.n497 B.n496 10.6151
R1458 B.n503 B.n502 10.6151
R1459 B.n504 B.n503 10.6151
R1460 B.n504 B.n329 10.6151
R1461 B.n514 B.n329 10.6151
R1462 B.n515 B.n514 10.6151
R1463 B.n516 B.n515 10.6151
R1464 B.n516 B.n321 10.6151
R1465 B.n526 B.n321 10.6151
R1466 B.n527 B.n526 10.6151
R1467 B.n528 B.n527 10.6151
R1468 B.n528 B.n313 10.6151
R1469 B.n538 B.n313 10.6151
R1470 B.n539 B.n538 10.6151
R1471 B.n540 B.n539 10.6151
R1472 B.n540 B.n305 10.6151
R1473 B.n550 B.n305 10.6151
R1474 B.n551 B.n550 10.6151
R1475 B.n552 B.n551 10.6151
R1476 B.n552 B.n297 10.6151
R1477 B.n562 B.n297 10.6151
R1478 B.n563 B.n562 10.6151
R1479 B.n564 B.n563 10.6151
R1480 B.n564 B.n289 10.6151
R1481 B.n574 B.n289 10.6151
R1482 B.n575 B.n574 10.6151
R1483 B.n576 B.n575 10.6151
R1484 B.n576 B.n281 10.6151
R1485 B.n587 B.n281 10.6151
R1486 B.n588 B.n587 10.6151
R1487 B.n589 B.n588 10.6151
R1488 B.n589 B.n274 10.6151
R1489 B.n599 B.n274 10.6151
R1490 B.n600 B.n599 10.6151
R1491 B.n601 B.n600 10.6151
R1492 B.n601 B.n266 10.6151
R1493 B.n611 B.n266 10.6151
R1494 B.n612 B.n611 10.6151
R1495 B.n613 B.n612 10.6151
R1496 B.n613 B.n258 10.6151
R1497 B.n623 B.n258 10.6151
R1498 B.n624 B.n623 10.6151
R1499 B.n625 B.n624 10.6151
R1500 B.n625 B.n250 10.6151
R1501 B.n636 B.n250 10.6151
R1502 B.n637 B.n636 10.6151
R1503 B.n638 B.n637 10.6151
R1504 B.n638 B.n0 10.6151
R1505 B.n801 B.n1 10.6151
R1506 B.n801 B.n800 10.6151
R1507 B.n800 B.n799 10.6151
R1508 B.n799 B.n10 10.6151
R1509 B.n793 B.n10 10.6151
R1510 B.n793 B.n792 10.6151
R1511 B.n792 B.n791 10.6151
R1512 B.n791 B.n17 10.6151
R1513 B.n785 B.n17 10.6151
R1514 B.n785 B.n784 10.6151
R1515 B.n784 B.n783 10.6151
R1516 B.n783 B.n24 10.6151
R1517 B.n777 B.n24 10.6151
R1518 B.n777 B.n776 10.6151
R1519 B.n776 B.n775 10.6151
R1520 B.n775 B.n31 10.6151
R1521 B.n769 B.n31 10.6151
R1522 B.n769 B.n768 10.6151
R1523 B.n768 B.n767 10.6151
R1524 B.n767 B.n37 10.6151
R1525 B.n761 B.n37 10.6151
R1526 B.n761 B.n760 10.6151
R1527 B.n760 B.n759 10.6151
R1528 B.n759 B.n45 10.6151
R1529 B.n753 B.n45 10.6151
R1530 B.n753 B.n752 10.6151
R1531 B.n752 B.n751 10.6151
R1532 B.n751 B.n52 10.6151
R1533 B.n745 B.n52 10.6151
R1534 B.n745 B.n744 10.6151
R1535 B.n744 B.n743 10.6151
R1536 B.n743 B.n59 10.6151
R1537 B.n737 B.n59 10.6151
R1538 B.n737 B.n736 10.6151
R1539 B.n736 B.n735 10.6151
R1540 B.n735 B.n66 10.6151
R1541 B.n729 B.n66 10.6151
R1542 B.n729 B.n728 10.6151
R1543 B.n728 B.n727 10.6151
R1544 B.n727 B.n73 10.6151
R1545 B.n721 B.n73 10.6151
R1546 B.n721 B.n720 10.6151
R1547 B.n720 B.n719 10.6151
R1548 B.n719 B.n80 10.6151
R1549 B.n713 B.n80 10.6151
R1550 B.n713 B.n712 10.6151
R1551 B.n712 B.n711 10.6151
R1552 B.n175 B.n126 9.36635
R1553 B.n198 B.n123 9.36635
R1554 B.n424 B.n423 9.36635
R1555 B.n448 B.n447 9.36635
R1556 B.n591 B.t2 9.08015
R1557 B.n771 B.t8 9.08015
R1558 B.n256 B.t9 5.44829
R1559 B.t5 B.n796 5.44829
R1560 B.n807 B.n0 2.81026
R1561 B.n807 B.n1 2.81026
R1562 B.n178 B.n126 1.24928
R1563 B.n195 B.n123 1.24928
R1564 B.n423 B.n360 1.24928
R1565 B.n447 B.n446 1.24928
R1566 VP.n18 VP.n15 161.3
R1567 VP.n20 VP.n19 161.3
R1568 VP.n21 VP.n14 161.3
R1569 VP.n23 VP.n22 161.3
R1570 VP.n24 VP.n13 161.3
R1571 VP.n26 VP.n25 161.3
R1572 VP.n27 VP.n12 161.3
R1573 VP.n29 VP.n28 161.3
R1574 VP.n30 VP.n11 161.3
R1575 VP.n33 VP.n32 161.3
R1576 VP.n34 VP.n10 161.3
R1577 VP.n36 VP.n35 161.3
R1578 VP.n37 VP.n9 161.3
R1579 VP.n68 VP.n0 161.3
R1580 VP.n67 VP.n66 161.3
R1581 VP.n65 VP.n1 161.3
R1582 VP.n64 VP.n63 161.3
R1583 VP.n61 VP.n2 161.3
R1584 VP.n60 VP.n59 161.3
R1585 VP.n58 VP.n3 161.3
R1586 VP.n57 VP.n56 161.3
R1587 VP.n55 VP.n4 161.3
R1588 VP.n54 VP.n53 161.3
R1589 VP.n52 VP.n5 161.3
R1590 VP.n51 VP.n50 161.3
R1591 VP.n49 VP.n6 161.3
R1592 VP.n47 VP.n46 161.3
R1593 VP.n45 VP.n7 161.3
R1594 VP.n44 VP.n43 161.3
R1595 VP.n42 VP.n8 161.3
R1596 VP.n16 VP.t5 117.356
R1597 VP.n41 VP.n40 86.3164
R1598 VP.n70 VP.n69 86.3164
R1599 VP.n39 VP.n38 86.3164
R1600 VP.n69 VP.t1 85.8567
R1601 VP.n55 VP.t2 85.8567
R1602 VP.n41 VP.t4 85.8567
R1603 VP.n48 VP.t6 85.8567
R1604 VP.n62 VP.t7 85.8567
R1605 VP.n24 VP.t8 85.8567
R1606 VP.n38 VP.t9 85.8567
R1607 VP.n31 VP.t3 85.8567
R1608 VP.n17 VP.t0 85.8567
R1609 VP.n17 VP.n16 58.0791
R1610 VP.n43 VP.n7 52.6866
R1611 VP.n50 VP.n5 52.6866
R1612 VP.n60 VP.n3 52.6866
R1613 VP.n67 VP.n1 52.6866
R1614 VP.n36 VP.n10 52.6866
R1615 VP.n29 VP.n12 52.6866
R1616 VP.n19 VP.n14 52.6866
R1617 VP.n40 VP.n39 45.5868
R1618 VP.n43 VP.n42 28.4674
R1619 VP.n54 VP.n5 28.4674
R1620 VP.n56 VP.n3 28.4674
R1621 VP.n68 VP.n67 28.4674
R1622 VP.n37 VP.n36 28.4674
R1623 VP.n25 VP.n12 28.4674
R1624 VP.n23 VP.n14 28.4674
R1625 VP.n42 VP.n41 24.5923
R1626 VP.n47 VP.n7 24.5923
R1627 VP.n50 VP.n49 24.5923
R1628 VP.n55 VP.n54 24.5923
R1629 VP.n56 VP.n55 24.5923
R1630 VP.n61 VP.n60 24.5923
R1631 VP.n63 VP.n1 24.5923
R1632 VP.n69 VP.n68 24.5923
R1633 VP.n38 VP.n37 24.5923
R1634 VP.n30 VP.n29 24.5923
R1635 VP.n32 VP.n10 24.5923
R1636 VP.n24 VP.n23 24.5923
R1637 VP.n25 VP.n24 24.5923
R1638 VP.n19 VP.n18 24.5923
R1639 VP.n16 VP.n15 12.6034
R1640 VP.n48 VP.n47 12.2964
R1641 VP.n49 VP.n48 12.2964
R1642 VP.n62 VP.n61 12.2964
R1643 VP.n63 VP.n62 12.2964
R1644 VP.n31 VP.n30 12.2964
R1645 VP.n32 VP.n31 12.2964
R1646 VP.n18 VP.n17 12.2964
R1647 VP.n39 VP.n9 0.278335
R1648 VP.n40 VP.n8 0.278335
R1649 VP.n70 VP.n0 0.278335
R1650 VP.n20 VP.n15 0.189894
R1651 VP.n21 VP.n20 0.189894
R1652 VP.n22 VP.n21 0.189894
R1653 VP.n22 VP.n13 0.189894
R1654 VP.n26 VP.n13 0.189894
R1655 VP.n27 VP.n26 0.189894
R1656 VP.n28 VP.n27 0.189894
R1657 VP.n28 VP.n11 0.189894
R1658 VP.n33 VP.n11 0.189894
R1659 VP.n34 VP.n33 0.189894
R1660 VP.n35 VP.n34 0.189894
R1661 VP.n35 VP.n9 0.189894
R1662 VP.n44 VP.n8 0.189894
R1663 VP.n45 VP.n44 0.189894
R1664 VP.n46 VP.n45 0.189894
R1665 VP.n46 VP.n6 0.189894
R1666 VP.n51 VP.n6 0.189894
R1667 VP.n52 VP.n51 0.189894
R1668 VP.n53 VP.n52 0.189894
R1669 VP.n53 VP.n4 0.189894
R1670 VP.n57 VP.n4 0.189894
R1671 VP.n58 VP.n57 0.189894
R1672 VP.n59 VP.n58 0.189894
R1673 VP.n59 VP.n2 0.189894
R1674 VP.n64 VP.n2 0.189894
R1675 VP.n65 VP.n64 0.189894
R1676 VP.n66 VP.n65 0.189894
R1677 VP.n66 VP.n0 0.189894
R1678 VP VP.n70 0.153485
R1679 VDD1.n1 VDD1.t4 72.1816
R1680 VDD1.n3 VDD1.t5 72.1815
R1681 VDD1.n5 VDD1.n4 68.7455
R1682 VDD1.n1 VDD1.n0 67.3472
R1683 VDD1.n7 VDD1.n6 67.3471
R1684 VDD1.n3 VDD1.n2 67.3461
R1685 VDD1.n7 VDD1.n5 40.3781
R1686 VDD1.n6 VDD1.t6 2.89524
R1687 VDD1.n6 VDD1.t0 2.89524
R1688 VDD1.n0 VDD1.t9 2.89524
R1689 VDD1.n0 VDD1.t1 2.89524
R1690 VDD1.n4 VDD1.t2 2.89524
R1691 VDD1.n4 VDD1.t8 2.89524
R1692 VDD1.n2 VDD1.t3 2.89524
R1693 VDD1.n2 VDD1.t7 2.89524
R1694 VDD1 VDD1.n7 1.39705
R1695 VDD1 VDD1.n1 0.543603
R1696 VDD1.n5 VDD1.n3 0.430068
C0 VN VTAIL 6.60993f
C1 VP VDD1 6.22283f
C2 VDD2 VDD1 1.73119f
C3 VP VDD2 0.496693f
C4 VN VDD1 0.152126f
C5 VDD1 VTAIL 7.70218f
C6 VN VP 6.43461f
C7 VP VTAIL 6.62418f
C8 VN VDD2 5.88107f
C9 VDD2 VTAIL 7.74924f
C10 VDD2 B 5.47356f
C11 VDD1 B 5.464736f
C12 VTAIL B 5.316459f
C13 VN B 14.34307f
C14 VP B 12.868841f
C15 VDD1.t4 B 1.34809f
C16 VDD1.t9 B 0.123364f
C17 VDD1.t1 B 0.123364f
C18 VDD1.n0 B 1.05357f
C19 VDD1.n1 B 0.733019f
C20 VDD1.t5 B 1.34808f
C21 VDD1.t3 B 0.123364f
C22 VDD1.t7 B 0.123364f
C23 VDD1.n2 B 1.05356f
C24 VDD1.n3 B 0.725914f
C25 VDD1.t2 B 0.123364f
C26 VDD1.t8 B 0.123364f
C27 VDD1.n4 B 1.06239f
C28 VDD1.n5 B 2.12759f
C29 VDD1.t6 B 0.123364f
C30 VDD1.t0 B 0.123364f
C31 VDD1.n6 B 1.05356f
C32 VDD1.n7 B 2.26466f
C33 VP.n0 B 0.037099f
C34 VP.t1 B 0.985237f
C35 VP.n1 B 0.049987f
C36 VP.n2 B 0.028141f
C37 VP.t7 B 0.985237f
C38 VP.n3 B 0.028882f
C39 VP.n4 B 0.028141f
C40 VP.t2 B 0.985237f
C41 VP.n5 B 0.028882f
C42 VP.n6 B 0.028141f
C43 VP.t6 B 0.985237f
C44 VP.n7 B 0.049987f
C45 VP.n8 B 0.037099f
C46 VP.t4 B 0.985237f
C47 VP.n9 B 0.037099f
C48 VP.t9 B 0.985237f
C49 VP.n10 B 0.049987f
C50 VP.n11 B 0.028141f
C51 VP.t3 B 0.985237f
C52 VP.n12 B 0.028882f
C53 VP.n13 B 0.028141f
C54 VP.t8 B 0.985237f
C55 VP.n14 B 0.028882f
C56 VP.n15 B 0.208436f
C57 VP.t0 B 0.985237f
C58 VP.t5 B 1.12185f
C59 VP.n16 B 0.438557f
C60 VP.n17 B 0.436221f
C61 VP.n18 B 0.039304f
C62 VP.n19 B 0.049987f
C63 VP.n20 B 0.028141f
C64 VP.n21 B 0.028141f
C65 VP.n22 B 0.028141f
C66 VP.n23 B 0.055131f
C67 VP.n24 B 0.397422f
C68 VP.n25 B 0.055131f
C69 VP.n26 B 0.028141f
C70 VP.n27 B 0.028141f
C71 VP.n28 B 0.028141f
C72 VP.n29 B 0.049987f
C73 VP.n30 B 0.039304f
C74 VP.n31 B 0.370999f
C75 VP.n32 B 0.039304f
C76 VP.n33 B 0.028141f
C77 VP.n34 B 0.028141f
C78 VP.n35 B 0.028141f
C79 VP.n36 B 0.028882f
C80 VP.n37 B 0.055131f
C81 VP.n38 B 0.461481f
C82 VP.n39 B 1.3464f
C83 VP.n40 B 1.36866f
C84 VP.n41 B 0.461481f
C85 VP.n42 B 0.055131f
C86 VP.n43 B 0.028882f
C87 VP.n44 B 0.028141f
C88 VP.n45 B 0.028141f
C89 VP.n46 B 0.028141f
C90 VP.n47 B 0.039304f
C91 VP.n48 B 0.370999f
C92 VP.n49 B 0.039304f
C93 VP.n50 B 0.049987f
C94 VP.n51 B 0.028141f
C95 VP.n52 B 0.028141f
C96 VP.n53 B 0.028141f
C97 VP.n54 B 0.055131f
C98 VP.n55 B 0.397422f
C99 VP.n56 B 0.055131f
C100 VP.n57 B 0.028141f
C101 VP.n58 B 0.028141f
C102 VP.n59 B 0.028141f
C103 VP.n60 B 0.049987f
C104 VP.n61 B 0.039304f
C105 VP.n62 B 0.370999f
C106 VP.n63 B 0.039304f
C107 VP.n64 B 0.028141f
C108 VP.n65 B 0.028141f
C109 VP.n66 B 0.028141f
C110 VP.n67 B 0.028882f
C111 VP.n68 B 0.055131f
C112 VP.n69 B 0.461481f
C113 VP.n70 B 0.029737f
C114 VDD2.t6 B 1.32704f
C115 VDD2.t1 B 0.121438f
C116 VDD2.t5 B 0.121438f
C117 VDD2.n0 B 1.03712f
C118 VDD2.n1 B 0.714581f
C119 VDD2.t0 B 0.121438f
C120 VDD2.t3 B 0.121438f
C121 VDD2.n2 B 1.0458f
C122 VDD2.n3 B 2.00128f
C123 VDD2.t7 B 1.31693f
C124 VDD2.n4 B 2.18969f
C125 VDD2.t4 B 0.121438f
C126 VDD2.t9 B 0.121438f
C127 VDD2.n5 B 1.03712f
C128 VDD2.n6 B 0.355286f
C129 VDD2.t8 B 0.121438f
C130 VDD2.t2 B 0.121438f
C131 VDD2.n7 B 1.04577f
C132 VTAIL.t11 B 0.145394f
C133 VTAIL.t14 B 0.145394f
C134 VTAIL.n0 B 1.1742f
C135 VTAIL.n1 B 0.497043f
C136 VTAIL.t19 B 1.49369f
C137 VTAIL.n2 B 0.611065f
C138 VTAIL.t2 B 0.145394f
C139 VTAIL.t0 B 0.145394f
C140 VTAIL.n3 B 1.1742f
C141 VTAIL.n4 B 0.577367f
C142 VTAIL.t1 B 0.145394f
C143 VTAIL.t4 B 0.145394f
C144 VTAIL.n5 B 1.1742f
C145 VTAIL.n6 B 1.62196f
C146 VTAIL.t17 B 0.145394f
C147 VTAIL.t9 B 0.145394f
C148 VTAIL.n7 B 1.17421f
C149 VTAIL.n8 B 1.62195f
C150 VTAIL.t10 B 0.145394f
C151 VTAIL.t18 B 0.145394f
C152 VTAIL.n9 B 1.17421f
C153 VTAIL.n10 B 0.577358f
C154 VTAIL.t16 B 1.49371f
C155 VTAIL.n11 B 0.611052f
C156 VTAIL.t5 B 0.145394f
C157 VTAIL.t6 B 0.145394f
C158 VTAIL.n12 B 1.17421f
C159 VTAIL.n13 B 0.534021f
C160 VTAIL.t8 B 0.145394f
C161 VTAIL.t3 B 0.145394f
C162 VTAIL.n14 B 1.17421f
C163 VTAIL.n15 B 0.577358f
C164 VTAIL.t7 B 1.49369f
C165 VTAIL.n16 B 1.53088f
C166 VTAIL.t12 B 1.49369f
C167 VTAIL.n17 B 1.53088f
C168 VTAIL.t15 B 0.145394f
C169 VTAIL.t13 B 0.145394f
C170 VTAIL.n18 B 1.1742f
C171 VTAIL.n19 B 0.446234f
C172 VN.n0 B 0.036444f
C173 VN.t6 B 0.967849f
C174 VN.n1 B 0.049105f
C175 VN.n2 B 0.027644f
C176 VN.t9 B 0.967849f
C177 VN.n3 B 0.028372f
C178 VN.n4 B 0.027644f
C179 VN.t4 B 0.967849f
C180 VN.n5 B 0.028372f
C181 VN.n6 B 0.204758f
C182 VN.t8 B 0.967849f
C183 VN.t3 B 1.10205f
C184 VN.n7 B 0.430817f
C185 VN.n8 B 0.428522f
C186 VN.n9 B 0.03861f
C187 VN.n10 B 0.049105f
C188 VN.n11 B 0.027644f
C189 VN.n12 B 0.027644f
C190 VN.n13 B 0.027644f
C191 VN.n14 B 0.054158f
C192 VN.n15 B 0.390408f
C193 VN.n16 B 0.054158f
C194 VN.n17 B 0.027644f
C195 VN.n18 B 0.027644f
C196 VN.n19 B 0.027644f
C197 VN.n20 B 0.049105f
C198 VN.n21 B 0.03861f
C199 VN.n22 B 0.364452f
C200 VN.n23 B 0.03861f
C201 VN.n24 B 0.027644f
C202 VN.n25 B 0.027644f
C203 VN.n26 B 0.027644f
C204 VN.n27 B 0.028372f
C205 VN.n28 B 0.054158f
C206 VN.n29 B 0.453336f
C207 VN.n30 B 0.029212f
C208 VN.n31 B 0.036444f
C209 VN.t2 B 0.967849f
C210 VN.n32 B 0.049105f
C211 VN.n33 B 0.027644f
C212 VN.t5 B 0.967849f
C213 VN.n34 B 0.028372f
C214 VN.n35 B 0.027644f
C215 VN.t0 B 0.967849f
C216 VN.n36 B 0.028372f
C217 VN.n37 B 0.204758f
C218 VN.t1 B 0.967849f
C219 VN.t7 B 1.10205f
C220 VN.n38 B 0.430817f
C221 VN.n39 B 0.428522f
C222 VN.n40 B 0.03861f
C223 VN.n41 B 0.049105f
C224 VN.n42 B 0.027644f
C225 VN.n43 B 0.027644f
C226 VN.n44 B 0.027644f
C227 VN.n45 B 0.054158f
C228 VN.n46 B 0.390408f
C229 VN.n47 B 0.054158f
C230 VN.n48 B 0.027644f
C231 VN.n49 B 0.027644f
C232 VN.n50 B 0.027644f
C233 VN.n51 B 0.049105f
C234 VN.n52 B 0.03861f
C235 VN.n53 B 0.364452f
C236 VN.n54 B 0.03861f
C237 VN.n55 B 0.027644f
C238 VN.n56 B 0.027644f
C239 VN.n57 B 0.027644f
C240 VN.n58 B 0.028372f
C241 VN.n59 B 0.054158f
C242 VN.n60 B 0.453336f
C243 VN.n61 B 1.33772f
.ends

