* NGSPICE file created from diff_pair_sample_1574.ext - technology: sky130A

.subckt diff_pair_sample_1574 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X1 VDD2.t9 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X2 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0 ps=0 w=0.72 l=3.7
X3 VDD1.t9 VP.t1 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.2808 ps=2.22 w=0.72 l=3.7
X4 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X5 VDD2.t7 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0.1188 ps=1.05 w=0.72 l=3.7
X6 VDD1.t1 VP.t2 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X7 VDD1.t6 VP.t3 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0.1188 ps=1.05 w=0.72 l=3.7
X8 VDD1.t2 VP.t4 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X9 VDD1.t4 VP.t5 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0.1188 ps=1.05 w=0.72 l=3.7
X10 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0 ps=0 w=0.72 l=3.7
X11 VTAIL.t5 VN.t3 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X12 VTAIL.t13 VP.t6 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X13 VDD1.t7 VP.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.2808 ps=2.22 w=0.72 l=3.7
X14 VTAIL.t11 VP.t8 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X15 VDD2.t5 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.2808 ps=2.22 w=0.72 l=3.7
X16 VDD2.t4 VN.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.2808 ps=2.22 w=0.72 l=3.7
X17 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0 ps=0 w=0.72 l=3.7
X18 VTAIL.t10 VP.t9 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X19 VDD2.t3 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0.1188 ps=1.05 w=0.72 l=3.7
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.2808 pd=2.22 as=0 ps=0 w=0.72 l=3.7
X21 VTAIL.t9 VN.t7 VDD2.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X22 VTAIL.t7 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
X23 VDD2.t0 VN.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1188 pd=1.05 as=0.1188 ps=1.05 w=0.72 l=3.7
R0 VP.n33 VP.n32 161.3
R1 VP.n34 VP.n29 161.3
R2 VP.n36 VP.n35 161.3
R3 VP.n37 VP.n28 161.3
R4 VP.n39 VP.n38 161.3
R5 VP.n40 VP.n27 161.3
R6 VP.n42 VP.n41 161.3
R7 VP.n43 VP.n26 161.3
R8 VP.n45 VP.n44 161.3
R9 VP.n46 VP.n25 161.3
R10 VP.n48 VP.n47 161.3
R11 VP.n49 VP.n24 161.3
R12 VP.n51 VP.n50 161.3
R13 VP.n52 VP.n23 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n22 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n21 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n20 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n19 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n68 VP.n18 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n125 VP.n124 161.3
R26 VP.n123 VP.n1 161.3
R27 VP.n122 VP.n121 161.3
R28 VP.n120 VP.n2 161.3
R29 VP.n119 VP.n118 161.3
R30 VP.n117 VP.n3 161.3
R31 VP.n116 VP.n115 161.3
R32 VP.n114 VP.n4 161.3
R33 VP.n113 VP.n112 161.3
R34 VP.n110 VP.n5 161.3
R35 VP.n109 VP.n108 161.3
R36 VP.n107 VP.n6 161.3
R37 VP.n106 VP.n105 161.3
R38 VP.n104 VP.n7 161.3
R39 VP.n103 VP.n102 161.3
R40 VP.n101 VP.n8 161.3
R41 VP.n100 VP.n99 161.3
R42 VP.n98 VP.n9 161.3
R43 VP.n97 VP.n96 161.3
R44 VP.n95 VP.n10 161.3
R45 VP.n94 VP.n93 161.3
R46 VP.n92 VP.n11 161.3
R47 VP.n91 VP.n90 161.3
R48 VP.n89 VP.n12 161.3
R49 VP.n88 VP.n87 161.3
R50 VP.n85 VP.n13 161.3
R51 VP.n84 VP.n83 161.3
R52 VP.n82 VP.n14 161.3
R53 VP.n81 VP.n80 161.3
R54 VP.n79 VP.n15 161.3
R55 VP.n78 VP.n77 161.3
R56 VP.n76 VP.n16 161.3
R57 VP.n75 VP.n74 161.3
R58 VP.n73 VP.n72 87.2945
R59 VP.n126 VP.n0 87.2945
R60 VP.n71 VP.n17 87.2945
R61 VP.n31 VP.n30 73.7076
R62 VP.n72 VP.n71 50.5791
R63 VP.n80 VP.n79 44.9365
R64 VP.n118 VP.n2 44.9365
R65 VP.n63 VP.n19 44.9365
R66 VP.n93 VP.n92 42.0302
R67 VP.n105 VP.n6 42.0302
R68 VP.n50 VP.n23 42.0302
R69 VP.n38 VP.n37 42.0302
R70 VP.n93 VP.n10 39.1239
R71 VP.n105 VP.n104 39.1239
R72 VP.n50 VP.n49 39.1239
R73 VP.n38 VP.n27 39.1239
R74 VP.n30 VP.t5 36.6421
R75 VP.n80 VP.n14 36.2176
R76 VP.n118 VP.n117 36.2176
R77 VP.n63 VP.n62 36.2176
R78 VP.n74 VP.n16 24.5923
R79 VP.n78 VP.n16 24.5923
R80 VP.n79 VP.n78 24.5923
R81 VP.n84 VP.n14 24.5923
R82 VP.n85 VP.n84 24.5923
R83 VP.n87 VP.n12 24.5923
R84 VP.n91 VP.n12 24.5923
R85 VP.n92 VP.n91 24.5923
R86 VP.n97 VP.n10 24.5923
R87 VP.n98 VP.n97 24.5923
R88 VP.n99 VP.n98 24.5923
R89 VP.n99 VP.n8 24.5923
R90 VP.n103 VP.n8 24.5923
R91 VP.n104 VP.n103 24.5923
R92 VP.n109 VP.n6 24.5923
R93 VP.n110 VP.n109 24.5923
R94 VP.n112 VP.n110 24.5923
R95 VP.n116 VP.n4 24.5923
R96 VP.n117 VP.n116 24.5923
R97 VP.n122 VP.n2 24.5923
R98 VP.n123 VP.n122 24.5923
R99 VP.n124 VP.n123 24.5923
R100 VP.n67 VP.n19 24.5923
R101 VP.n68 VP.n67 24.5923
R102 VP.n69 VP.n68 24.5923
R103 VP.n54 VP.n23 24.5923
R104 VP.n55 VP.n54 24.5923
R105 VP.n57 VP.n55 24.5923
R106 VP.n61 VP.n21 24.5923
R107 VP.n62 VP.n61 24.5923
R108 VP.n42 VP.n27 24.5923
R109 VP.n43 VP.n42 24.5923
R110 VP.n44 VP.n43 24.5923
R111 VP.n44 VP.n25 24.5923
R112 VP.n48 VP.n25 24.5923
R113 VP.n49 VP.n48 24.5923
R114 VP.n32 VP.n29 24.5923
R115 VP.n36 VP.n29 24.5923
R116 VP.n37 VP.n36 24.5923
R117 VP.n86 VP.n85 23.1168
R118 VP.n111 VP.n4 23.1168
R119 VP.n56 VP.n21 23.1168
R120 VP.n99 VP.t2 4.69023
R121 VP.n73 VP.t3 4.69023
R122 VP.n86 VP.t6 4.69023
R123 VP.n111 VP.t8 4.69023
R124 VP.n0 VP.t1 4.69023
R125 VP.n44 VP.t4 4.69023
R126 VP.n17 VP.t7 4.69023
R127 VP.n56 VP.t9 4.69023
R128 VP.n31 VP.t0 4.69023
R129 VP.n33 VP.n30 3.364
R130 VP.n74 VP.n73 2.95152
R131 VP.n124 VP.n0 2.95152
R132 VP.n69 VP.n17 2.95152
R133 VP.n87 VP.n86 1.47601
R134 VP.n112 VP.n111 1.47601
R135 VP.n57 VP.n56 1.47601
R136 VP.n32 VP.n31 1.47601
R137 VP.n71 VP.n70 0.354861
R138 VP.n75 VP.n72 0.354861
R139 VP.n126 VP.n125 0.354861
R140 VP VP.n126 0.267071
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n28 0.189894
R144 VP.n39 VP.n28 0.189894
R145 VP.n40 VP.n39 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n41 VP.n26 0.189894
R148 VP.n45 VP.n26 0.189894
R149 VP.n46 VP.n45 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n47 VP.n24 0.189894
R152 VP.n51 VP.n24 0.189894
R153 VP.n52 VP.n51 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n53 VP.n22 0.189894
R156 VP.n58 VP.n22 0.189894
R157 VP.n59 VP.n58 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n60 VP.n20 0.189894
R160 VP.n64 VP.n20 0.189894
R161 VP.n65 VP.n64 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n66 VP.n18 0.189894
R164 VP.n70 VP.n18 0.189894
R165 VP.n76 VP.n75 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n77 VP.n15 0.189894
R168 VP.n81 VP.n15 0.189894
R169 VP.n82 VP.n81 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n83 VP.n13 0.189894
R172 VP.n88 VP.n13 0.189894
R173 VP.n89 VP.n88 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n90 VP.n11 0.189894
R176 VP.n94 VP.n11 0.189894
R177 VP.n95 VP.n94 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n96 VP.n9 0.189894
R180 VP.n100 VP.n9 0.189894
R181 VP.n101 VP.n100 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n102 VP.n7 0.189894
R184 VP.n106 VP.n7 0.189894
R185 VP.n107 VP.n106 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n108 VP.n5 0.189894
R188 VP.n113 VP.n5 0.189894
R189 VP.n114 VP.n113 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n115 VP.n3 0.189894
R192 VP.n119 VP.n3 0.189894
R193 VP.n120 VP.n119 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n121 VP.n1 0.189894
R196 VP.n125 VP.n1 0.189894
R197 VDD1.n1 VDD1.t4 267.166
R198 VDD1.n3 VDD1.t6 267.166
R199 VDD1.n5 VDD1.n4 238.742
R200 VDD1.n7 VDD1.n6 236.191
R201 VDD1.n1 VDD1.n0 236.191
R202 VDD1.n3 VDD1.n2 236.191
R203 VDD1.n7 VDD1.n5 43.1582
R204 VDD1.n6 VDD1.t0 27.5005
R205 VDD1.n6 VDD1.t7 27.5005
R206 VDD1.n0 VDD1.t5 27.5005
R207 VDD1.n0 VDD1.t2 27.5005
R208 VDD1.n4 VDD1.t3 27.5005
R209 VDD1.n4 VDD1.t9 27.5005
R210 VDD1.n2 VDD1.t8 27.5005
R211 VDD1.n2 VDD1.t1 27.5005
R212 VDD1 VDD1.n7 2.54791
R213 VDD1 VDD1.n1 0.927224
R214 VDD1.n5 VDD1.n3 0.813688
R215 VTAIL.n17 VTAIL.t8 247.012
R216 VTAIL.n2 VTAIL.t18 247.012
R217 VTAIL.n16 VTAIL.t12 247.012
R218 VTAIL.n11 VTAIL.t6 247.012
R219 VTAIL.n19 VTAIL.n18 219.512
R220 VTAIL.n1 VTAIL.n0 219.512
R221 VTAIL.n4 VTAIL.n3 219.512
R222 VTAIL.n6 VTAIL.n5 219.512
R223 VTAIL.n15 VTAIL.n14 219.512
R224 VTAIL.n13 VTAIL.n12 219.512
R225 VTAIL.n10 VTAIL.n9 219.512
R226 VTAIL.n8 VTAIL.n7 219.512
R227 VTAIL.n18 VTAIL.t3 27.5005
R228 VTAIL.n18 VTAIL.t9 27.5005
R229 VTAIL.n0 VTAIL.t4 27.5005
R230 VTAIL.n0 VTAIL.t7 27.5005
R231 VTAIL.n3 VTAIL.t17 27.5005
R232 VTAIL.n3 VTAIL.t11 27.5005
R233 VTAIL.n5 VTAIL.t16 27.5005
R234 VTAIL.n5 VTAIL.t13 27.5005
R235 VTAIL.n14 VTAIL.t15 27.5005
R236 VTAIL.n14 VTAIL.t10 27.5005
R237 VTAIL.n12 VTAIL.t14 27.5005
R238 VTAIL.n12 VTAIL.t19 27.5005
R239 VTAIL.n9 VTAIL.t1 27.5005
R240 VTAIL.n9 VTAIL.t2 27.5005
R241 VTAIL.n7 VTAIL.t0 27.5005
R242 VTAIL.n7 VTAIL.t5 27.5005
R243 VTAIL.n8 VTAIL.n6 19.9358
R244 VTAIL.n17 VTAIL.n16 16.4617
R245 VTAIL.n10 VTAIL.n8 3.47464
R246 VTAIL.n11 VTAIL.n10 3.47464
R247 VTAIL.n15 VTAIL.n13 3.47464
R248 VTAIL.n16 VTAIL.n15 3.47464
R249 VTAIL.n6 VTAIL.n4 3.47464
R250 VTAIL.n4 VTAIL.n2 3.47464
R251 VTAIL.n19 VTAIL.n17 3.47464
R252 VTAIL VTAIL.n1 2.66429
R253 VTAIL.n13 VTAIL.n11 2.2074
R254 VTAIL.n2 VTAIL.n1 2.2074
R255 VTAIL VTAIL.n19 0.810845
R256 B.n771 B.n770 585
R257 B.n208 B.n156 585
R258 B.n207 B.n206 585
R259 B.n205 B.n204 585
R260 B.n203 B.n202 585
R261 B.n201 B.n200 585
R262 B.n199 B.n198 585
R263 B.n197 B.n196 585
R264 B.n195 B.n194 585
R265 B.n193 B.n192 585
R266 B.n191 B.n190 585
R267 B.n189 B.n188 585
R268 B.n187 B.n186 585
R269 B.n185 B.n184 585
R270 B.n183 B.n182 585
R271 B.n181 B.n180 585
R272 B.n179 B.n178 585
R273 B.n177 B.n176 585
R274 B.n175 B.n174 585
R275 B.n173 B.n172 585
R276 B.n171 B.n170 585
R277 B.n169 B.n168 585
R278 B.n167 B.n166 585
R279 B.n165 B.n164 585
R280 B.n144 B.n143 585
R281 B.n776 B.n775 585
R282 B.n769 B.n157 585
R283 B.n157 B.n141 585
R284 B.n768 B.n140 585
R285 B.n780 B.n140 585
R286 B.n767 B.n139 585
R287 B.n781 B.n139 585
R288 B.n766 B.n138 585
R289 B.n782 B.n138 585
R290 B.n765 B.n764 585
R291 B.n764 B.n134 585
R292 B.n763 B.n133 585
R293 B.n788 B.n133 585
R294 B.n762 B.n132 585
R295 B.n789 B.n132 585
R296 B.n761 B.n131 585
R297 B.n790 B.n131 585
R298 B.n760 B.n759 585
R299 B.n759 B.n127 585
R300 B.n758 B.n126 585
R301 B.t18 B.n126 585
R302 B.n757 B.n125 585
R303 B.n796 B.n125 585
R304 B.n756 B.n124 585
R305 B.n797 B.n124 585
R306 B.n755 B.n754 585
R307 B.n754 B.n120 585
R308 B.n753 B.n119 585
R309 B.n803 B.n119 585
R310 B.n752 B.n118 585
R311 B.n804 B.n118 585
R312 B.n751 B.n117 585
R313 B.n805 B.n117 585
R314 B.n750 B.n749 585
R315 B.n749 B.n113 585
R316 B.n748 B.n112 585
R317 B.n811 B.n112 585
R318 B.n747 B.n111 585
R319 B.n812 B.n111 585
R320 B.n746 B.n110 585
R321 B.n813 B.n110 585
R322 B.n745 B.n744 585
R323 B.n744 B.n106 585
R324 B.n743 B.n105 585
R325 B.n819 B.n105 585
R326 B.n742 B.n104 585
R327 B.n820 B.n104 585
R328 B.n741 B.n103 585
R329 B.n821 B.n103 585
R330 B.n740 B.n739 585
R331 B.n739 B.n102 585
R332 B.n738 B.n98 585
R333 B.n827 B.n98 585
R334 B.n737 B.n97 585
R335 B.n828 B.n97 585
R336 B.n736 B.n96 585
R337 B.n829 B.n96 585
R338 B.n735 B.n734 585
R339 B.n734 B.n92 585
R340 B.n733 B.n91 585
R341 B.n835 B.n91 585
R342 B.n732 B.n90 585
R343 B.n836 B.n90 585
R344 B.n731 B.n89 585
R345 B.n837 B.n89 585
R346 B.n730 B.n729 585
R347 B.n729 B.n85 585
R348 B.n728 B.n84 585
R349 B.n843 B.n84 585
R350 B.n727 B.n83 585
R351 B.n844 B.n83 585
R352 B.n726 B.n82 585
R353 B.n845 B.n82 585
R354 B.n725 B.n724 585
R355 B.n724 B.n78 585
R356 B.n723 B.n77 585
R357 B.n851 B.n77 585
R358 B.n722 B.n76 585
R359 B.n852 B.n76 585
R360 B.n721 B.n75 585
R361 B.n853 B.n75 585
R362 B.n720 B.n719 585
R363 B.n719 B.n71 585
R364 B.n718 B.n70 585
R365 B.n859 B.n70 585
R366 B.n717 B.n69 585
R367 B.n860 B.n69 585
R368 B.n716 B.n68 585
R369 B.n861 B.n68 585
R370 B.n715 B.n714 585
R371 B.n714 B.n64 585
R372 B.n713 B.n63 585
R373 B.n867 B.n63 585
R374 B.n712 B.n62 585
R375 B.n868 B.n62 585
R376 B.n711 B.n61 585
R377 B.n869 B.n61 585
R378 B.n710 B.n709 585
R379 B.n709 B.n57 585
R380 B.n708 B.n56 585
R381 B.n875 B.n56 585
R382 B.n707 B.n55 585
R383 B.n876 B.n55 585
R384 B.n706 B.n54 585
R385 B.n877 B.n54 585
R386 B.n705 B.n704 585
R387 B.n704 B.n50 585
R388 B.n703 B.n49 585
R389 B.n883 B.n49 585
R390 B.n702 B.n48 585
R391 B.n884 B.n48 585
R392 B.n701 B.n47 585
R393 B.n885 B.n47 585
R394 B.n700 B.n699 585
R395 B.n699 B.n43 585
R396 B.n698 B.n42 585
R397 B.n891 B.n42 585
R398 B.n697 B.n41 585
R399 B.n892 B.n41 585
R400 B.n696 B.n40 585
R401 B.n893 B.n40 585
R402 B.n695 B.n694 585
R403 B.n694 B.n36 585
R404 B.n693 B.n35 585
R405 B.n899 B.n35 585
R406 B.n692 B.n34 585
R407 B.n900 B.n34 585
R408 B.n691 B.n33 585
R409 B.n901 B.n33 585
R410 B.n690 B.n689 585
R411 B.n689 B.n29 585
R412 B.n688 B.n28 585
R413 B.n907 B.n28 585
R414 B.n687 B.n27 585
R415 B.n908 B.n27 585
R416 B.n686 B.n26 585
R417 B.n909 B.n26 585
R418 B.n685 B.n684 585
R419 B.n684 B.n22 585
R420 B.n683 B.n21 585
R421 B.n915 B.n21 585
R422 B.n682 B.n20 585
R423 B.n916 B.n20 585
R424 B.n681 B.n19 585
R425 B.n917 B.n19 585
R426 B.n680 B.n679 585
R427 B.n679 B.n15 585
R428 B.n678 B.n14 585
R429 B.n923 B.n14 585
R430 B.n677 B.n13 585
R431 B.n924 B.n13 585
R432 B.n676 B.n12 585
R433 B.n925 B.n12 585
R434 B.n675 B.n674 585
R435 B.n674 B.n8 585
R436 B.n673 B.n7 585
R437 B.n931 B.n7 585
R438 B.n672 B.n6 585
R439 B.n932 B.n6 585
R440 B.n671 B.n5 585
R441 B.n933 B.n5 585
R442 B.n670 B.n669 585
R443 B.n669 B.n4 585
R444 B.n668 B.n209 585
R445 B.n668 B.n667 585
R446 B.n658 B.n210 585
R447 B.n211 B.n210 585
R448 B.n660 B.n659 585
R449 B.n661 B.n660 585
R450 B.n657 B.n216 585
R451 B.n216 B.n215 585
R452 B.n656 B.n655 585
R453 B.n655 B.n654 585
R454 B.n218 B.n217 585
R455 B.n219 B.n218 585
R456 B.n647 B.n646 585
R457 B.n648 B.n647 585
R458 B.n645 B.n224 585
R459 B.n224 B.n223 585
R460 B.n644 B.n643 585
R461 B.n643 B.n642 585
R462 B.n226 B.n225 585
R463 B.n227 B.n226 585
R464 B.n635 B.n634 585
R465 B.n636 B.n635 585
R466 B.n633 B.n232 585
R467 B.n232 B.n231 585
R468 B.n632 B.n631 585
R469 B.n631 B.n630 585
R470 B.n234 B.n233 585
R471 B.n235 B.n234 585
R472 B.n623 B.n622 585
R473 B.n624 B.n623 585
R474 B.n621 B.n240 585
R475 B.n240 B.n239 585
R476 B.n620 B.n619 585
R477 B.n619 B.n618 585
R478 B.n242 B.n241 585
R479 B.n243 B.n242 585
R480 B.n611 B.n610 585
R481 B.n612 B.n611 585
R482 B.n609 B.n248 585
R483 B.n248 B.n247 585
R484 B.n608 B.n607 585
R485 B.n607 B.n606 585
R486 B.n250 B.n249 585
R487 B.n251 B.n250 585
R488 B.n599 B.n598 585
R489 B.n600 B.n599 585
R490 B.n597 B.n256 585
R491 B.n256 B.n255 585
R492 B.n596 B.n595 585
R493 B.n595 B.n594 585
R494 B.n258 B.n257 585
R495 B.n259 B.n258 585
R496 B.n587 B.n586 585
R497 B.n588 B.n587 585
R498 B.n585 B.n264 585
R499 B.n264 B.n263 585
R500 B.n584 B.n583 585
R501 B.n583 B.n582 585
R502 B.n266 B.n265 585
R503 B.n267 B.n266 585
R504 B.n575 B.n574 585
R505 B.n576 B.n575 585
R506 B.n573 B.n272 585
R507 B.n272 B.n271 585
R508 B.n572 B.n571 585
R509 B.n571 B.n570 585
R510 B.n274 B.n273 585
R511 B.n275 B.n274 585
R512 B.n563 B.n562 585
R513 B.n564 B.n563 585
R514 B.n561 B.n280 585
R515 B.n280 B.n279 585
R516 B.n560 B.n559 585
R517 B.n559 B.n558 585
R518 B.n282 B.n281 585
R519 B.n283 B.n282 585
R520 B.n551 B.n550 585
R521 B.n552 B.n551 585
R522 B.n549 B.n288 585
R523 B.n288 B.n287 585
R524 B.n548 B.n547 585
R525 B.n547 B.n546 585
R526 B.n290 B.n289 585
R527 B.n291 B.n290 585
R528 B.n539 B.n538 585
R529 B.n540 B.n539 585
R530 B.n537 B.n296 585
R531 B.n296 B.n295 585
R532 B.n536 B.n535 585
R533 B.n535 B.n534 585
R534 B.n298 B.n297 585
R535 B.n299 B.n298 585
R536 B.n527 B.n526 585
R537 B.n528 B.n527 585
R538 B.n525 B.n304 585
R539 B.n304 B.n303 585
R540 B.n524 B.n523 585
R541 B.n523 B.n522 585
R542 B.n306 B.n305 585
R543 B.n307 B.n306 585
R544 B.n515 B.n514 585
R545 B.n516 B.n515 585
R546 B.n513 B.n312 585
R547 B.n312 B.n311 585
R548 B.n512 B.n511 585
R549 B.n511 B.n510 585
R550 B.n314 B.n313 585
R551 B.n503 B.n314 585
R552 B.n502 B.n501 585
R553 B.n504 B.n502 585
R554 B.n500 B.n319 585
R555 B.n319 B.n318 585
R556 B.n499 B.n498 585
R557 B.n498 B.n497 585
R558 B.n321 B.n320 585
R559 B.n322 B.n321 585
R560 B.n490 B.n489 585
R561 B.n491 B.n490 585
R562 B.n488 B.n327 585
R563 B.n327 B.n326 585
R564 B.n487 B.n486 585
R565 B.n486 B.n485 585
R566 B.n329 B.n328 585
R567 B.n330 B.n329 585
R568 B.n478 B.n477 585
R569 B.n479 B.n478 585
R570 B.n476 B.n335 585
R571 B.n335 B.n334 585
R572 B.n475 B.n474 585
R573 B.n474 B.n473 585
R574 B.n337 B.n336 585
R575 B.n338 B.n337 585
R576 B.n466 B.n465 585
R577 B.n467 B.n466 585
R578 B.n464 B.n343 585
R579 B.n343 B.n342 585
R580 B.n463 B.n462 585
R581 B.n462 B.t11 585
R582 B.n345 B.n344 585
R583 B.n346 B.n345 585
R584 B.n455 B.n454 585
R585 B.n456 B.n455 585
R586 B.n453 B.n351 585
R587 B.n351 B.n350 585
R588 B.n452 B.n451 585
R589 B.n451 B.n450 585
R590 B.n353 B.n352 585
R591 B.n354 B.n353 585
R592 B.n443 B.n442 585
R593 B.n444 B.n443 585
R594 B.n441 B.n359 585
R595 B.n359 B.n358 585
R596 B.n440 B.n439 585
R597 B.n439 B.n438 585
R598 B.n361 B.n360 585
R599 B.n362 B.n361 585
R600 B.n434 B.n433 585
R601 B.n365 B.n364 585
R602 B.n430 B.n429 585
R603 B.n431 B.n430 585
R604 B.n428 B.n378 585
R605 B.n427 B.n426 585
R606 B.n425 B.n424 585
R607 B.n423 B.n422 585
R608 B.n421 B.n420 585
R609 B.n418 B.n417 585
R610 B.n416 B.n415 585
R611 B.n414 B.n413 585
R612 B.n412 B.n411 585
R613 B.n410 B.n409 585
R614 B.n408 B.n407 585
R615 B.n406 B.n405 585
R616 B.n404 B.n403 585
R617 B.n402 B.n401 585
R618 B.n400 B.n399 585
R619 B.n397 B.n396 585
R620 B.n395 B.n394 585
R621 B.n393 B.n392 585
R622 B.n391 B.n390 585
R623 B.n389 B.n388 585
R624 B.n387 B.n386 585
R625 B.n385 B.n384 585
R626 B.n383 B.n377 585
R627 B.n431 B.n377 585
R628 B.n435 B.n363 585
R629 B.n363 B.n362 585
R630 B.n437 B.n436 585
R631 B.n438 B.n437 585
R632 B.n357 B.n356 585
R633 B.n358 B.n357 585
R634 B.n446 B.n445 585
R635 B.n445 B.n444 585
R636 B.n447 B.n355 585
R637 B.n355 B.n354 585
R638 B.n449 B.n448 585
R639 B.n450 B.n449 585
R640 B.n349 B.n348 585
R641 B.n350 B.n349 585
R642 B.n458 B.n457 585
R643 B.n457 B.n456 585
R644 B.n459 B.n347 585
R645 B.n347 B.n346 585
R646 B.n461 B.n460 585
R647 B.t11 B.n461 585
R648 B.n341 B.n340 585
R649 B.n342 B.n341 585
R650 B.n469 B.n468 585
R651 B.n468 B.n467 585
R652 B.n470 B.n339 585
R653 B.n339 B.n338 585
R654 B.n472 B.n471 585
R655 B.n473 B.n472 585
R656 B.n333 B.n332 585
R657 B.n334 B.n333 585
R658 B.n481 B.n480 585
R659 B.n480 B.n479 585
R660 B.n482 B.n331 585
R661 B.n331 B.n330 585
R662 B.n484 B.n483 585
R663 B.n485 B.n484 585
R664 B.n325 B.n324 585
R665 B.n326 B.n325 585
R666 B.n493 B.n492 585
R667 B.n492 B.n491 585
R668 B.n494 B.n323 585
R669 B.n323 B.n322 585
R670 B.n496 B.n495 585
R671 B.n497 B.n496 585
R672 B.n317 B.n316 585
R673 B.n318 B.n317 585
R674 B.n506 B.n505 585
R675 B.n505 B.n504 585
R676 B.n507 B.n315 585
R677 B.n503 B.n315 585
R678 B.n509 B.n508 585
R679 B.n510 B.n509 585
R680 B.n310 B.n309 585
R681 B.n311 B.n310 585
R682 B.n518 B.n517 585
R683 B.n517 B.n516 585
R684 B.n519 B.n308 585
R685 B.n308 B.n307 585
R686 B.n521 B.n520 585
R687 B.n522 B.n521 585
R688 B.n302 B.n301 585
R689 B.n303 B.n302 585
R690 B.n530 B.n529 585
R691 B.n529 B.n528 585
R692 B.n531 B.n300 585
R693 B.n300 B.n299 585
R694 B.n533 B.n532 585
R695 B.n534 B.n533 585
R696 B.n294 B.n293 585
R697 B.n295 B.n294 585
R698 B.n542 B.n541 585
R699 B.n541 B.n540 585
R700 B.n543 B.n292 585
R701 B.n292 B.n291 585
R702 B.n545 B.n544 585
R703 B.n546 B.n545 585
R704 B.n286 B.n285 585
R705 B.n287 B.n286 585
R706 B.n554 B.n553 585
R707 B.n553 B.n552 585
R708 B.n555 B.n284 585
R709 B.n284 B.n283 585
R710 B.n557 B.n556 585
R711 B.n558 B.n557 585
R712 B.n278 B.n277 585
R713 B.n279 B.n278 585
R714 B.n566 B.n565 585
R715 B.n565 B.n564 585
R716 B.n567 B.n276 585
R717 B.n276 B.n275 585
R718 B.n569 B.n568 585
R719 B.n570 B.n569 585
R720 B.n270 B.n269 585
R721 B.n271 B.n270 585
R722 B.n578 B.n577 585
R723 B.n577 B.n576 585
R724 B.n579 B.n268 585
R725 B.n268 B.n267 585
R726 B.n581 B.n580 585
R727 B.n582 B.n581 585
R728 B.n262 B.n261 585
R729 B.n263 B.n262 585
R730 B.n590 B.n589 585
R731 B.n589 B.n588 585
R732 B.n591 B.n260 585
R733 B.n260 B.n259 585
R734 B.n593 B.n592 585
R735 B.n594 B.n593 585
R736 B.n254 B.n253 585
R737 B.n255 B.n254 585
R738 B.n602 B.n601 585
R739 B.n601 B.n600 585
R740 B.n603 B.n252 585
R741 B.n252 B.n251 585
R742 B.n605 B.n604 585
R743 B.n606 B.n605 585
R744 B.n246 B.n245 585
R745 B.n247 B.n246 585
R746 B.n614 B.n613 585
R747 B.n613 B.n612 585
R748 B.n615 B.n244 585
R749 B.n244 B.n243 585
R750 B.n617 B.n616 585
R751 B.n618 B.n617 585
R752 B.n238 B.n237 585
R753 B.n239 B.n238 585
R754 B.n626 B.n625 585
R755 B.n625 B.n624 585
R756 B.n627 B.n236 585
R757 B.n236 B.n235 585
R758 B.n629 B.n628 585
R759 B.n630 B.n629 585
R760 B.n230 B.n229 585
R761 B.n231 B.n230 585
R762 B.n638 B.n637 585
R763 B.n637 B.n636 585
R764 B.n639 B.n228 585
R765 B.n228 B.n227 585
R766 B.n641 B.n640 585
R767 B.n642 B.n641 585
R768 B.n222 B.n221 585
R769 B.n223 B.n222 585
R770 B.n650 B.n649 585
R771 B.n649 B.n648 585
R772 B.n651 B.n220 585
R773 B.n220 B.n219 585
R774 B.n653 B.n652 585
R775 B.n654 B.n653 585
R776 B.n214 B.n213 585
R777 B.n215 B.n214 585
R778 B.n663 B.n662 585
R779 B.n662 B.n661 585
R780 B.n664 B.n212 585
R781 B.n212 B.n211 585
R782 B.n666 B.n665 585
R783 B.n667 B.n666 585
R784 B.n2 B.n0 585
R785 B.n4 B.n2 585
R786 B.n3 B.n1 585
R787 B.n932 B.n3 585
R788 B.n930 B.n929 585
R789 B.n931 B.n930 585
R790 B.n928 B.n9 585
R791 B.n9 B.n8 585
R792 B.n927 B.n926 585
R793 B.n926 B.n925 585
R794 B.n11 B.n10 585
R795 B.n924 B.n11 585
R796 B.n922 B.n921 585
R797 B.n923 B.n922 585
R798 B.n920 B.n16 585
R799 B.n16 B.n15 585
R800 B.n919 B.n918 585
R801 B.n918 B.n917 585
R802 B.n18 B.n17 585
R803 B.n916 B.n18 585
R804 B.n914 B.n913 585
R805 B.n915 B.n914 585
R806 B.n912 B.n23 585
R807 B.n23 B.n22 585
R808 B.n911 B.n910 585
R809 B.n910 B.n909 585
R810 B.n25 B.n24 585
R811 B.n908 B.n25 585
R812 B.n906 B.n905 585
R813 B.n907 B.n906 585
R814 B.n904 B.n30 585
R815 B.n30 B.n29 585
R816 B.n903 B.n902 585
R817 B.n902 B.n901 585
R818 B.n32 B.n31 585
R819 B.n900 B.n32 585
R820 B.n898 B.n897 585
R821 B.n899 B.n898 585
R822 B.n896 B.n37 585
R823 B.n37 B.n36 585
R824 B.n895 B.n894 585
R825 B.n894 B.n893 585
R826 B.n39 B.n38 585
R827 B.n892 B.n39 585
R828 B.n890 B.n889 585
R829 B.n891 B.n890 585
R830 B.n888 B.n44 585
R831 B.n44 B.n43 585
R832 B.n887 B.n886 585
R833 B.n886 B.n885 585
R834 B.n46 B.n45 585
R835 B.n884 B.n46 585
R836 B.n882 B.n881 585
R837 B.n883 B.n882 585
R838 B.n880 B.n51 585
R839 B.n51 B.n50 585
R840 B.n879 B.n878 585
R841 B.n878 B.n877 585
R842 B.n53 B.n52 585
R843 B.n876 B.n53 585
R844 B.n874 B.n873 585
R845 B.n875 B.n874 585
R846 B.n872 B.n58 585
R847 B.n58 B.n57 585
R848 B.n871 B.n870 585
R849 B.n870 B.n869 585
R850 B.n60 B.n59 585
R851 B.n868 B.n60 585
R852 B.n866 B.n865 585
R853 B.n867 B.n866 585
R854 B.n864 B.n65 585
R855 B.n65 B.n64 585
R856 B.n863 B.n862 585
R857 B.n862 B.n861 585
R858 B.n67 B.n66 585
R859 B.n860 B.n67 585
R860 B.n858 B.n857 585
R861 B.n859 B.n858 585
R862 B.n856 B.n72 585
R863 B.n72 B.n71 585
R864 B.n855 B.n854 585
R865 B.n854 B.n853 585
R866 B.n74 B.n73 585
R867 B.n852 B.n74 585
R868 B.n850 B.n849 585
R869 B.n851 B.n850 585
R870 B.n848 B.n79 585
R871 B.n79 B.n78 585
R872 B.n847 B.n846 585
R873 B.n846 B.n845 585
R874 B.n81 B.n80 585
R875 B.n844 B.n81 585
R876 B.n842 B.n841 585
R877 B.n843 B.n842 585
R878 B.n840 B.n86 585
R879 B.n86 B.n85 585
R880 B.n839 B.n838 585
R881 B.n838 B.n837 585
R882 B.n88 B.n87 585
R883 B.n836 B.n88 585
R884 B.n834 B.n833 585
R885 B.n835 B.n834 585
R886 B.n832 B.n93 585
R887 B.n93 B.n92 585
R888 B.n831 B.n830 585
R889 B.n830 B.n829 585
R890 B.n95 B.n94 585
R891 B.n828 B.n95 585
R892 B.n826 B.n825 585
R893 B.n827 B.n826 585
R894 B.n824 B.n99 585
R895 B.n102 B.n99 585
R896 B.n823 B.n822 585
R897 B.n822 B.n821 585
R898 B.n101 B.n100 585
R899 B.n820 B.n101 585
R900 B.n818 B.n817 585
R901 B.n819 B.n818 585
R902 B.n816 B.n107 585
R903 B.n107 B.n106 585
R904 B.n815 B.n814 585
R905 B.n814 B.n813 585
R906 B.n109 B.n108 585
R907 B.n812 B.n109 585
R908 B.n810 B.n809 585
R909 B.n811 B.n810 585
R910 B.n808 B.n114 585
R911 B.n114 B.n113 585
R912 B.n807 B.n806 585
R913 B.n806 B.n805 585
R914 B.n116 B.n115 585
R915 B.n804 B.n116 585
R916 B.n802 B.n801 585
R917 B.n803 B.n802 585
R918 B.n800 B.n121 585
R919 B.n121 B.n120 585
R920 B.n799 B.n798 585
R921 B.n798 B.n797 585
R922 B.n123 B.n122 585
R923 B.n796 B.n123 585
R924 B.n795 B.n794 585
R925 B.t18 B.n795 585
R926 B.n793 B.n128 585
R927 B.n128 B.n127 585
R928 B.n792 B.n791 585
R929 B.n791 B.n790 585
R930 B.n130 B.n129 585
R931 B.n789 B.n130 585
R932 B.n787 B.n786 585
R933 B.n788 B.n787 585
R934 B.n785 B.n135 585
R935 B.n135 B.n134 585
R936 B.n784 B.n783 585
R937 B.n783 B.n782 585
R938 B.n137 B.n136 585
R939 B.n781 B.n137 585
R940 B.n779 B.n778 585
R941 B.n780 B.n779 585
R942 B.n777 B.n142 585
R943 B.n142 B.n141 585
R944 B.n935 B.n934 585
R945 B.n934 B.n933 585
R946 B.n433 B.n363 574.183
R947 B.n775 B.n142 574.183
R948 B.n377 B.n361 574.183
R949 B.n771 B.n157 574.183
R950 B.n381 B.t13 314.318
R951 B.n379 B.t16 314.318
R952 B.n161 B.t19 314.318
R953 B.n158 B.t22 314.318
R954 B.n773 B.n772 256.663
R955 B.n773 B.n155 256.663
R956 B.n773 B.n154 256.663
R957 B.n773 B.n153 256.663
R958 B.n773 B.n152 256.663
R959 B.n773 B.n151 256.663
R960 B.n773 B.n150 256.663
R961 B.n773 B.n149 256.663
R962 B.n773 B.n148 256.663
R963 B.n773 B.n147 256.663
R964 B.n773 B.n146 256.663
R965 B.n773 B.n145 256.663
R966 B.n774 B.n773 256.663
R967 B.n432 B.n431 256.663
R968 B.n431 B.n366 256.663
R969 B.n431 B.n367 256.663
R970 B.n431 B.n368 256.663
R971 B.n431 B.n369 256.663
R972 B.n431 B.n370 256.663
R973 B.n431 B.n371 256.663
R974 B.n431 B.n372 256.663
R975 B.n431 B.n373 256.663
R976 B.n431 B.n374 256.663
R977 B.n431 B.n375 256.663
R978 B.n431 B.n376 256.663
R979 B.n431 B.n362 255.047
R980 B.n773 B.n141 255.047
R981 B.n382 B.t12 236.161
R982 B.n380 B.t15 236.161
R983 B.n162 B.t20 236.161
R984 B.n159 B.t23 236.161
R985 B.n381 B.t10 210.113
R986 B.n379 B.t14 210.113
R987 B.n161 B.t17 210.113
R988 B.n158 B.t21 210.113
R989 B.n437 B.n363 163.367
R990 B.n437 B.n357 163.367
R991 B.n445 B.n357 163.367
R992 B.n445 B.n355 163.367
R993 B.n449 B.n355 163.367
R994 B.n449 B.n349 163.367
R995 B.n457 B.n349 163.367
R996 B.n457 B.n347 163.367
R997 B.n461 B.n347 163.367
R998 B.n461 B.n341 163.367
R999 B.n468 B.n341 163.367
R1000 B.n468 B.n339 163.367
R1001 B.n472 B.n339 163.367
R1002 B.n472 B.n333 163.367
R1003 B.n480 B.n333 163.367
R1004 B.n480 B.n331 163.367
R1005 B.n484 B.n331 163.367
R1006 B.n484 B.n325 163.367
R1007 B.n492 B.n325 163.367
R1008 B.n492 B.n323 163.367
R1009 B.n496 B.n323 163.367
R1010 B.n496 B.n317 163.367
R1011 B.n505 B.n317 163.367
R1012 B.n505 B.n315 163.367
R1013 B.n509 B.n315 163.367
R1014 B.n509 B.n310 163.367
R1015 B.n517 B.n310 163.367
R1016 B.n517 B.n308 163.367
R1017 B.n521 B.n308 163.367
R1018 B.n521 B.n302 163.367
R1019 B.n529 B.n302 163.367
R1020 B.n529 B.n300 163.367
R1021 B.n533 B.n300 163.367
R1022 B.n533 B.n294 163.367
R1023 B.n541 B.n294 163.367
R1024 B.n541 B.n292 163.367
R1025 B.n545 B.n292 163.367
R1026 B.n545 B.n286 163.367
R1027 B.n553 B.n286 163.367
R1028 B.n553 B.n284 163.367
R1029 B.n557 B.n284 163.367
R1030 B.n557 B.n278 163.367
R1031 B.n565 B.n278 163.367
R1032 B.n565 B.n276 163.367
R1033 B.n569 B.n276 163.367
R1034 B.n569 B.n270 163.367
R1035 B.n577 B.n270 163.367
R1036 B.n577 B.n268 163.367
R1037 B.n581 B.n268 163.367
R1038 B.n581 B.n262 163.367
R1039 B.n589 B.n262 163.367
R1040 B.n589 B.n260 163.367
R1041 B.n593 B.n260 163.367
R1042 B.n593 B.n254 163.367
R1043 B.n601 B.n254 163.367
R1044 B.n601 B.n252 163.367
R1045 B.n605 B.n252 163.367
R1046 B.n605 B.n246 163.367
R1047 B.n613 B.n246 163.367
R1048 B.n613 B.n244 163.367
R1049 B.n617 B.n244 163.367
R1050 B.n617 B.n238 163.367
R1051 B.n625 B.n238 163.367
R1052 B.n625 B.n236 163.367
R1053 B.n629 B.n236 163.367
R1054 B.n629 B.n230 163.367
R1055 B.n637 B.n230 163.367
R1056 B.n637 B.n228 163.367
R1057 B.n641 B.n228 163.367
R1058 B.n641 B.n222 163.367
R1059 B.n649 B.n222 163.367
R1060 B.n649 B.n220 163.367
R1061 B.n653 B.n220 163.367
R1062 B.n653 B.n214 163.367
R1063 B.n662 B.n214 163.367
R1064 B.n662 B.n212 163.367
R1065 B.n666 B.n212 163.367
R1066 B.n666 B.n2 163.367
R1067 B.n934 B.n2 163.367
R1068 B.n934 B.n3 163.367
R1069 B.n930 B.n3 163.367
R1070 B.n930 B.n9 163.367
R1071 B.n926 B.n9 163.367
R1072 B.n926 B.n11 163.367
R1073 B.n922 B.n11 163.367
R1074 B.n922 B.n16 163.367
R1075 B.n918 B.n16 163.367
R1076 B.n918 B.n18 163.367
R1077 B.n914 B.n18 163.367
R1078 B.n914 B.n23 163.367
R1079 B.n910 B.n23 163.367
R1080 B.n910 B.n25 163.367
R1081 B.n906 B.n25 163.367
R1082 B.n906 B.n30 163.367
R1083 B.n902 B.n30 163.367
R1084 B.n902 B.n32 163.367
R1085 B.n898 B.n32 163.367
R1086 B.n898 B.n37 163.367
R1087 B.n894 B.n37 163.367
R1088 B.n894 B.n39 163.367
R1089 B.n890 B.n39 163.367
R1090 B.n890 B.n44 163.367
R1091 B.n886 B.n44 163.367
R1092 B.n886 B.n46 163.367
R1093 B.n882 B.n46 163.367
R1094 B.n882 B.n51 163.367
R1095 B.n878 B.n51 163.367
R1096 B.n878 B.n53 163.367
R1097 B.n874 B.n53 163.367
R1098 B.n874 B.n58 163.367
R1099 B.n870 B.n58 163.367
R1100 B.n870 B.n60 163.367
R1101 B.n866 B.n60 163.367
R1102 B.n866 B.n65 163.367
R1103 B.n862 B.n65 163.367
R1104 B.n862 B.n67 163.367
R1105 B.n858 B.n67 163.367
R1106 B.n858 B.n72 163.367
R1107 B.n854 B.n72 163.367
R1108 B.n854 B.n74 163.367
R1109 B.n850 B.n74 163.367
R1110 B.n850 B.n79 163.367
R1111 B.n846 B.n79 163.367
R1112 B.n846 B.n81 163.367
R1113 B.n842 B.n81 163.367
R1114 B.n842 B.n86 163.367
R1115 B.n838 B.n86 163.367
R1116 B.n838 B.n88 163.367
R1117 B.n834 B.n88 163.367
R1118 B.n834 B.n93 163.367
R1119 B.n830 B.n93 163.367
R1120 B.n830 B.n95 163.367
R1121 B.n826 B.n95 163.367
R1122 B.n826 B.n99 163.367
R1123 B.n822 B.n99 163.367
R1124 B.n822 B.n101 163.367
R1125 B.n818 B.n101 163.367
R1126 B.n818 B.n107 163.367
R1127 B.n814 B.n107 163.367
R1128 B.n814 B.n109 163.367
R1129 B.n810 B.n109 163.367
R1130 B.n810 B.n114 163.367
R1131 B.n806 B.n114 163.367
R1132 B.n806 B.n116 163.367
R1133 B.n802 B.n116 163.367
R1134 B.n802 B.n121 163.367
R1135 B.n798 B.n121 163.367
R1136 B.n798 B.n123 163.367
R1137 B.n795 B.n123 163.367
R1138 B.n795 B.n128 163.367
R1139 B.n791 B.n128 163.367
R1140 B.n791 B.n130 163.367
R1141 B.n787 B.n130 163.367
R1142 B.n787 B.n135 163.367
R1143 B.n783 B.n135 163.367
R1144 B.n783 B.n137 163.367
R1145 B.n779 B.n137 163.367
R1146 B.n779 B.n142 163.367
R1147 B.n430 B.n365 163.367
R1148 B.n430 B.n378 163.367
R1149 B.n426 B.n425 163.367
R1150 B.n422 B.n421 163.367
R1151 B.n417 B.n416 163.367
R1152 B.n413 B.n412 163.367
R1153 B.n409 B.n408 163.367
R1154 B.n405 B.n404 163.367
R1155 B.n401 B.n400 163.367
R1156 B.n396 B.n395 163.367
R1157 B.n392 B.n391 163.367
R1158 B.n388 B.n387 163.367
R1159 B.n384 B.n377 163.367
R1160 B.n439 B.n361 163.367
R1161 B.n439 B.n359 163.367
R1162 B.n443 B.n359 163.367
R1163 B.n443 B.n353 163.367
R1164 B.n451 B.n353 163.367
R1165 B.n451 B.n351 163.367
R1166 B.n455 B.n351 163.367
R1167 B.n455 B.n345 163.367
R1168 B.n462 B.n345 163.367
R1169 B.n462 B.n343 163.367
R1170 B.n466 B.n343 163.367
R1171 B.n466 B.n337 163.367
R1172 B.n474 B.n337 163.367
R1173 B.n474 B.n335 163.367
R1174 B.n478 B.n335 163.367
R1175 B.n478 B.n329 163.367
R1176 B.n486 B.n329 163.367
R1177 B.n486 B.n327 163.367
R1178 B.n490 B.n327 163.367
R1179 B.n490 B.n321 163.367
R1180 B.n498 B.n321 163.367
R1181 B.n498 B.n319 163.367
R1182 B.n502 B.n319 163.367
R1183 B.n502 B.n314 163.367
R1184 B.n511 B.n314 163.367
R1185 B.n511 B.n312 163.367
R1186 B.n515 B.n312 163.367
R1187 B.n515 B.n306 163.367
R1188 B.n523 B.n306 163.367
R1189 B.n523 B.n304 163.367
R1190 B.n527 B.n304 163.367
R1191 B.n527 B.n298 163.367
R1192 B.n535 B.n298 163.367
R1193 B.n535 B.n296 163.367
R1194 B.n539 B.n296 163.367
R1195 B.n539 B.n290 163.367
R1196 B.n547 B.n290 163.367
R1197 B.n547 B.n288 163.367
R1198 B.n551 B.n288 163.367
R1199 B.n551 B.n282 163.367
R1200 B.n559 B.n282 163.367
R1201 B.n559 B.n280 163.367
R1202 B.n563 B.n280 163.367
R1203 B.n563 B.n274 163.367
R1204 B.n571 B.n274 163.367
R1205 B.n571 B.n272 163.367
R1206 B.n575 B.n272 163.367
R1207 B.n575 B.n266 163.367
R1208 B.n583 B.n266 163.367
R1209 B.n583 B.n264 163.367
R1210 B.n587 B.n264 163.367
R1211 B.n587 B.n258 163.367
R1212 B.n595 B.n258 163.367
R1213 B.n595 B.n256 163.367
R1214 B.n599 B.n256 163.367
R1215 B.n599 B.n250 163.367
R1216 B.n607 B.n250 163.367
R1217 B.n607 B.n248 163.367
R1218 B.n611 B.n248 163.367
R1219 B.n611 B.n242 163.367
R1220 B.n619 B.n242 163.367
R1221 B.n619 B.n240 163.367
R1222 B.n623 B.n240 163.367
R1223 B.n623 B.n234 163.367
R1224 B.n631 B.n234 163.367
R1225 B.n631 B.n232 163.367
R1226 B.n635 B.n232 163.367
R1227 B.n635 B.n226 163.367
R1228 B.n643 B.n226 163.367
R1229 B.n643 B.n224 163.367
R1230 B.n647 B.n224 163.367
R1231 B.n647 B.n218 163.367
R1232 B.n655 B.n218 163.367
R1233 B.n655 B.n216 163.367
R1234 B.n660 B.n216 163.367
R1235 B.n660 B.n210 163.367
R1236 B.n668 B.n210 163.367
R1237 B.n669 B.n668 163.367
R1238 B.n669 B.n5 163.367
R1239 B.n6 B.n5 163.367
R1240 B.n7 B.n6 163.367
R1241 B.n674 B.n7 163.367
R1242 B.n674 B.n12 163.367
R1243 B.n13 B.n12 163.367
R1244 B.n14 B.n13 163.367
R1245 B.n679 B.n14 163.367
R1246 B.n679 B.n19 163.367
R1247 B.n20 B.n19 163.367
R1248 B.n21 B.n20 163.367
R1249 B.n684 B.n21 163.367
R1250 B.n684 B.n26 163.367
R1251 B.n27 B.n26 163.367
R1252 B.n28 B.n27 163.367
R1253 B.n689 B.n28 163.367
R1254 B.n689 B.n33 163.367
R1255 B.n34 B.n33 163.367
R1256 B.n35 B.n34 163.367
R1257 B.n694 B.n35 163.367
R1258 B.n694 B.n40 163.367
R1259 B.n41 B.n40 163.367
R1260 B.n42 B.n41 163.367
R1261 B.n699 B.n42 163.367
R1262 B.n699 B.n47 163.367
R1263 B.n48 B.n47 163.367
R1264 B.n49 B.n48 163.367
R1265 B.n704 B.n49 163.367
R1266 B.n704 B.n54 163.367
R1267 B.n55 B.n54 163.367
R1268 B.n56 B.n55 163.367
R1269 B.n709 B.n56 163.367
R1270 B.n709 B.n61 163.367
R1271 B.n62 B.n61 163.367
R1272 B.n63 B.n62 163.367
R1273 B.n714 B.n63 163.367
R1274 B.n714 B.n68 163.367
R1275 B.n69 B.n68 163.367
R1276 B.n70 B.n69 163.367
R1277 B.n719 B.n70 163.367
R1278 B.n719 B.n75 163.367
R1279 B.n76 B.n75 163.367
R1280 B.n77 B.n76 163.367
R1281 B.n724 B.n77 163.367
R1282 B.n724 B.n82 163.367
R1283 B.n83 B.n82 163.367
R1284 B.n84 B.n83 163.367
R1285 B.n729 B.n84 163.367
R1286 B.n729 B.n89 163.367
R1287 B.n90 B.n89 163.367
R1288 B.n91 B.n90 163.367
R1289 B.n734 B.n91 163.367
R1290 B.n734 B.n96 163.367
R1291 B.n97 B.n96 163.367
R1292 B.n98 B.n97 163.367
R1293 B.n739 B.n98 163.367
R1294 B.n739 B.n103 163.367
R1295 B.n104 B.n103 163.367
R1296 B.n105 B.n104 163.367
R1297 B.n744 B.n105 163.367
R1298 B.n744 B.n110 163.367
R1299 B.n111 B.n110 163.367
R1300 B.n112 B.n111 163.367
R1301 B.n749 B.n112 163.367
R1302 B.n749 B.n117 163.367
R1303 B.n118 B.n117 163.367
R1304 B.n119 B.n118 163.367
R1305 B.n754 B.n119 163.367
R1306 B.n754 B.n124 163.367
R1307 B.n125 B.n124 163.367
R1308 B.n126 B.n125 163.367
R1309 B.n759 B.n126 163.367
R1310 B.n759 B.n131 163.367
R1311 B.n132 B.n131 163.367
R1312 B.n133 B.n132 163.367
R1313 B.n764 B.n133 163.367
R1314 B.n764 B.n138 163.367
R1315 B.n139 B.n138 163.367
R1316 B.n140 B.n139 163.367
R1317 B.n157 B.n140 163.367
R1318 B.n164 B.n144 163.367
R1319 B.n168 B.n167 163.367
R1320 B.n172 B.n171 163.367
R1321 B.n176 B.n175 163.367
R1322 B.n180 B.n179 163.367
R1323 B.n184 B.n183 163.367
R1324 B.n188 B.n187 163.367
R1325 B.n192 B.n191 163.367
R1326 B.n196 B.n195 163.367
R1327 B.n200 B.n199 163.367
R1328 B.n204 B.n203 163.367
R1329 B.n206 B.n156 163.367
R1330 B.n438 B.n362 124.772
R1331 B.n438 B.n358 124.772
R1332 B.n444 B.n358 124.772
R1333 B.n444 B.n354 124.772
R1334 B.n450 B.n354 124.772
R1335 B.n450 B.n350 124.772
R1336 B.n456 B.n350 124.772
R1337 B.n456 B.n346 124.772
R1338 B.t11 B.n346 124.772
R1339 B.t11 B.n342 124.772
R1340 B.n467 B.n342 124.772
R1341 B.n467 B.n338 124.772
R1342 B.n473 B.n338 124.772
R1343 B.n473 B.n334 124.772
R1344 B.n479 B.n334 124.772
R1345 B.n479 B.n330 124.772
R1346 B.n485 B.n330 124.772
R1347 B.n485 B.n326 124.772
R1348 B.n491 B.n326 124.772
R1349 B.n491 B.n322 124.772
R1350 B.n497 B.n322 124.772
R1351 B.n497 B.n318 124.772
R1352 B.n504 B.n318 124.772
R1353 B.n504 B.n503 124.772
R1354 B.n510 B.n311 124.772
R1355 B.n516 B.n311 124.772
R1356 B.n516 B.n307 124.772
R1357 B.n522 B.n307 124.772
R1358 B.n522 B.n303 124.772
R1359 B.n528 B.n303 124.772
R1360 B.n528 B.n299 124.772
R1361 B.n534 B.n299 124.772
R1362 B.n534 B.n295 124.772
R1363 B.n540 B.n295 124.772
R1364 B.n546 B.n291 124.772
R1365 B.n546 B.n287 124.772
R1366 B.n552 B.n287 124.772
R1367 B.n552 B.n283 124.772
R1368 B.n558 B.n283 124.772
R1369 B.n558 B.n279 124.772
R1370 B.n564 B.n279 124.772
R1371 B.n564 B.n275 124.772
R1372 B.n570 B.n275 124.772
R1373 B.n570 B.n271 124.772
R1374 B.n576 B.n271 124.772
R1375 B.n582 B.n267 124.772
R1376 B.n582 B.n263 124.772
R1377 B.n588 B.n263 124.772
R1378 B.n588 B.n259 124.772
R1379 B.n594 B.n259 124.772
R1380 B.n594 B.n255 124.772
R1381 B.n600 B.n255 124.772
R1382 B.n600 B.n251 124.772
R1383 B.n606 B.n251 124.772
R1384 B.n606 B.n247 124.772
R1385 B.n612 B.n247 124.772
R1386 B.n618 B.n243 124.772
R1387 B.n618 B.n239 124.772
R1388 B.n624 B.n239 124.772
R1389 B.n624 B.n235 124.772
R1390 B.n630 B.n235 124.772
R1391 B.n630 B.n231 124.772
R1392 B.n636 B.n231 124.772
R1393 B.n636 B.n227 124.772
R1394 B.n642 B.n227 124.772
R1395 B.n642 B.n223 124.772
R1396 B.n648 B.n223 124.772
R1397 B.n654 B.n219 124.772
R1398 B.n654 B.n215 124.772
R1399 B.n661 B.n215 124.772
R1400 B.n661 B.n211 124.772
R1401 B.n667 B.n211 124.772
R1402 B.n667 B.n4 124.772
R1403 B.n933 B.n4 124.772
R1404 B.n933 B.n932 124.772
R1405 B.n932 B.n931 124.772
R1406 B.n931 B.n8 124.772
R1407 B.n925 B.n8 124.772
R1408 B.n925 B.n924 124.772
R1409 B.n924 B.n923 124.772
R1410 B.n923 B.n15 124.772
R1411 B.n917 B.n916 124.772
R1412 B.n916 B.n915 124.772
R1413 B.n915 B.n22 124.772
R1414 B.n909 B.n22 124.772
R1415 B.n909 B.n908 124.772
R1416 B.n908 B.n907 124.772
R1417 B.n907 B.n29 124.772
R1418 B.n901 B.n29 124.772
R1419 B.n901 B.n900 124.772
R1420 B.n900 B.n899 124.772
R1421 B.n899 B.n36 124.772
R1422 B.n893 B.n892 124.772
R1423 B.n892 B.n891 124.772
R1424 B.n891 B.n43 124.772
R1425 B.n885 B.n43 124.772
R1426 B.n885 B.n884 124.772
R1427 B.n884 B.n883 124.772
R1428 B.n883 B.n50 124.772
R1429 B.n877 B.n50 124.772
R1430 B.n877 B.n876 124.772
R1431 B.n876 B.n875 124.772
R1432 B.n875 B.n57 124.772
R1433 B.n869 B.n868 124.772
R1434 B.n868 B.n867 124.772
R1435 B.n867 B.n64 124.772
R1436 B.n861 B.n64 124.772
R1437 B.n861 B.n860 124.772
R1438 B.n860 B.n859 124.772
R1439 B.n859 B.n71 124.772
R1440 B.n853 B.n71 124.772
R1441 B.n853 B.n852 124.772
R1442 B.n852 B.n851 124.772
R1443 B.n851 B.n78 124.772
R1444 B.n845 B.n844 124.772
R1445 B.n844 B.n843 124.772
R1446 B.n843 B.n85 124.772
R1447 B.n837 B.n85 124.772
R1448 B.n837 B.n836 124.772
R1449 B.n836 B.n835 124.772
R1450 B.n835 B.n92 124.772
R1451 B.n829 B.n92 124.772
R1452 B.n829 B.n828 124.772
R1453 B.n828 B.n827 124.772
R1454 B.n821 B.n102 124.772
R1455 B.n821 B.n820 124.772
R1456 B.n820 B.n819 124.772
R1457 B.n819 B.n106 124.772
R1458 B.n813 B.n106 124.772
R1459 B.n813 B.n812 124.772
R1460 B.n812 B.n811 124.772
R1461 B.n811 B.n113 124.772
R1462 B.n805 B.n113 124.772
R1463 B.n805 B.n804 124.772
R1464 B.n804 B.n803 124.772
R1465 B.n803 B.n120 124.772
R1466 B.n797 B.n120 124.772
R1467 B.n797 B.n796 124.772
R1468 B.n796 B.t18 124.772
R1469 B.t18 B.n127 124.772
R1470 B.n790 B.n127 124.772
R1471 B.n790 B.n789 124.772
R1472 B.n789 B.n788 124.772
R1473 B.n788 B.n134 124.772
R1474 B.n782 B.n134 124.772
R1475 B.n782 B.n781 124.772
R1476 B.n781 B.n780 124.772
R1477 B.n780 B.n141 124.772
R1478 B.n510 B.t0 117.431
R1479 B.n827 B.t8 117.431
R1480 B.n540 B.t5 113.761
R1481 B.n845 B.t9 113.761
R1482 B.n576 B.t1 95.4133
R1483 B.n869 B.t3 95.4133
R1484 B.n382 B.n381 78.1581
R1485 B.n380 B.n379 78.1581
R1486 B.n162 B.n161 78.1581
R1487 B.n159 B.n158 78.1581
R1488 B.n612 B.t2 77.0647
R1489 B.n893 B.t7 77.0647
R1490 B.n433 B.n432 71.676
R1491 B.n378 B.n366 71.676
R1492 B.n425 B.n367 71.676
R1493 B.n421 B.n368 71.676
R1494 B.n416 B.n369 71.676
R1495 B.n412 B.n370 71.676
R1496 B.n408 B.n371 71.676
R1497 B.n404 B.n372 71.676
R1498 B.n400 B.n373 71.676
R1499 B.n395 B.n374 71.676
R1500 B.n391 B.n375 71.676
R1501 B.n387 B.n376 71.676
R1502 B.n775 B.n774 71.676
R1503 B.n164 B.n145 71.676
R1504 B.n168 B.n146 71.676
R1505 B.n172 B.n147 71.676
R1506 B.n176 B.n148 71.676
R1507 B.n180 B.n149 71.676
R1508 B.n184 B.n150 71.676
R1509 B.n188 B.n151 71.676
R1510 B.n192 B.n152 71.676
R1511 B.n196 B.n153 71.676
R1512 B.n200 B.n154 71.676
R1513 B.n204 B.n155 71.676
R1514 B.n772 B.n156 71.676
R1515 B.n772 B.n771 71.676
R1516 B.n206 B.n155 71.676
R1517 B.n203 B.n154 71.676
R1518 B.n199 B.n153 71.676
R1519 B.n195 B.n152 71.676
R1520 B.n191 B.n151 71.676
R1521 B.n187 B.n150 71.676
R1522 B.n183 B.n149 71.676
R1523 B.n179 B.n148 71.676
R1524 B.n175 B.n147 71.676
R1525 B.n171 B.n146 71.676
R1526 B.n167 B.n145 71.676
R1527 B.n774 B.n144 71.676
R1528 B.n432 B.n365 71.676
R1529 B.n426 B.n366 71.676
R1530 B.n422 B.n367 71.676
R1531 B.n417 B.n368 71.676
R1532 B.n413 B.n369 71.676
R1533 B.n409 B.n370 71.676
R1534 B.n405 B.n371 71.676
R1535 B.n401 B.n372 71.676
R1536 B.n396 B.n373 71.676
R1537 B.n392 B.n374 71.676
R1538 B.n388 B.n375 71.676
R1539 B.n384 B.n376 71.676
R1540 B.t6 B.n219 66.0555
R1541 B.t4 B.n15 66.0555
R1542 B.n398 B.n382 59.5399
R1543 B.n419 B.n380 59.5399
R1544 B.n163 B.n162 59.5399
R1545 B.n160 B.n159 59.5399
R1546 B.n648 B.t6 58.7161
R1547 B.n917 B.t4 58.7161
R1548 B.t2 B.n243 47.7069
R1549 B.t7 B.n36 47.7069
R1550 B.n777 B.n776 37.3078
R1551 B.n770 B.n769 37.3078
R1552 B.n383 B.n360 37.3078
R1553 B.n435 B.n434 37.3078
R1554 B.t1 B.n267 29.3583
R1555 B.t3 B.n57 29.3583
R1556 B B.n935 18.0485
R1557 B.t5 B.n291 11.0097
R1558 B.t9 B.n78 11.0097
R1559 B.n776 B.n143 10.6151
R1560 B.n165 B.n143 10.6151
R1561 B.n166 B.n165 10.6151
R1562 B.n169 B.n166 10.6151
R1563 B.n170 B.n169 10.6151
R1564 B.n173 B.n170 10.6151
R1565 B.n174 B.n173 10.6151
R1566 B.n178 B.n177 10.6151
R1567 B.n181 B.n178 10.6151
R1568 B.n182 B.n181 10.6151
R1569 B.n185 B.n182 10.6151
R1570 B.n186 B.n185 10.6151
R1571 B.n189 B.n186 10.6151
R1572 B.n190 B.n189 10.6151
R1573 B.n193 B.n190 10.6151
R1574 B.n194 B.n193 10.6151
R1575 B.n198 B.n197 10.6151
R1576 B.n201 B.n198 10.6151
R1577 B.n202 B.n201 10.6151
R1578 B.n205 B.n202 10.6151
R1579 B.n207 B.n205 10.6151
R1580 B.n208 B.n207 10.6151
R1581 B.n770 B.n208 10.6151
R1582 B.n440 B.n360 10.6151
R1583 B.n441 B.n440 10.6151
R1584 B.n442 B.n441 10.6151
R1585 B.n442 B.n352 10.6151
R1586 B.n452 B.n352 10.6151
R1587 B.n453 B.n452 10.6151
R1588 B.n454 B.n453 10.6151
R1589 B.n454 B.n344 10.6151
R1590 B.n463 B.n344 10.6151
R1591 B.n464 B.n463 10.6151
R1592 B.n465 B.n464 10.6151
R1593 B.n465 B.n336 10.6151
R1594 B.n475 B.n336 10.6151
R1595 B.n476 B.n475 10.6151
R1596 B.n477 B.n476 10.6151
R1597 B.n477 B.n328 10.6151
R1598 B.n487 B.n328 10.6151
R1599 B.n488 B.n487 10.6151
R1600 B.n489 B.n488 10.6151
R1601 B.n489 B.n320 10.6151
R1602 B.n499 B.n320 10.6151
R1603 B.n500 B.n499 10.6151
R1604 B.n501 B.n500 10.6151
R1605 B.n501 B.n313 10.6151
R1606 B.n512 B.n313 10.6151
R1607 B.n513 B.n512 10.6151
R1608 B.n514 B.n513 10.6151
R1609 B.n514 B.n305 10.6151
R1610 B.n524 B.n305 10.6151
R1611 B.n525 B.n524 10.6151
R1612 B.n526 B.n525 10.6151
R1613 B.n526 B.n297 10.6151
R1614 B.n536 B.n297 10.6151
R1615 B.n537 B.n536 10.6151
R1616 B.n538 B.n537 10.6151
R1617 B.n538 B.n289 10.6151
R1618 B.n548 B.n289 10.6151
R1619 B.n549 B.n548 10.6151
R1620 B.n550 B.n549 10.6151
R1621 B.n550 B.n281 10.6151
R1622 B.n560 B.n281 10.6151
R1623 B.n561 B.n560 10.6151
R1624 B.n562 B.n561 10.6151
R1625 B.n562 B.n273 10.6151
R1626 B.n572 B.n273 10.6151
R1627 B.n573 B.n572 10.6151
R1628 B.n574 B.n573 10.6151
R1629 B.n574 B.n265 10.6151
R1630 B.n584 B.n265 10.6151
R1631 B.n585 B.n584 10.6151
R1632 B.n586 B.n585 10.6151
R1633 B.n586 B.n257 10.6151
R1634 B.n596 B.n257 10.6151
R1635 B.n597 B.n596 10.6151
R1636 B.n598 B.n597 10.6151
R1637 B.n598 B.n249 10.6151
R1638 B.n608 B.n249 10.6151
R1639 B.n609 B.n608 10.6151
R1640 B.n610 B.n609 10.6151
R1641 B.n610 B.n241 10.6151
R1642 B.n620 B.n241 10.6151
R1643 B.n621 B.n620 10.6151
R1644 B.n622 B.n621 10.6151
R1645 B.n622 B.n233 10.6151
R1646 B.n632 B.n233 10.6151
R1647 B.n633 B.n632 10.6151
R1648 B.n634 B.n633 10.6151
R1649 B.n634 B.n225 10.6151
R1650 B.n644 B.n225 10.6151
R1651 B.n645 B.n644 10.6151
R1652 B.n646 B.n645 10.6151
R1653 B.n646 B.n217 10.6151
R1654 B.n656 B.n217 10.6151
R1655 B.n657 B.n656 10.6151
R1656 B.n659 B.n657 10.6151
R1657 B.n659 B.n658 10.6151
R1658 B.n658 B.n209 10.6151
R1659 B.n670 B.n209 10.6151
R1660 B.n671 B.n670 10.6151
R1661 B.n672 B.n671 10.6151
R1662 B.n673 B.n672 10.6151
R1663 B.n675 B.n673 10.6151
R1664 B.n676 B.n675 10.6151
R1665 B.n677 B.n676 10.6151
R1666 B.n678 B.n677 10.6151
R1667 B.n680 B.n678 10.6151
R1668 B.n681 B.n680 10.6151
R1669 B.n682 B.n681 10.6151
R1670 B.n683 B.n682 10.6151
R1671 B.n685 B.n683 10.6151
R1672 B.n686 B.n685 10.6151
R1673 B.n687 B.n686 10.6151
R1674 B.n688 B.n687 10.6151
R1675 B.n690 B.n688 10.6151
R1676 B.n691 B.n690 10.6151
R1677 B.n692 B.n691 10.6151
R1678 B.n693 B.n692 10.6151
R1679 B.n695 B.n693 10.6151
R1680 B.n696 B.n695 10.6151
R1681 B.n697 B.n696 10.6151
R1682 B.n698 B.n697 10.6151
R1683 B.n700 B.n698 10.6151
R1684 B.n701 B.n700 10.6151
R1685 B.n702 B.n701 10.6151
R1686 B.n703 B.n702 10.6151
R1687 B.n705 B.n703 10.6151
R1688 B.n706 B.n705 10.6151
R1689 B.n707 B.n706 10.6151
R1690 B.n708 B.n707 10.6151
R1691 B.n710 B.n708 10.6151
R1692 B.n711 B.n710 10.6151
R1693 B.n712 B.n711 10.6151
R1694 B.n713 B.n712 10.6151
R1695 B.n715 B.n713 10.6151
R1696 B.n716 B.n715 10.6151
R1697 B.n717 B.n716 10.6151
R1698 B.n718 B.n717 10.6151
R1699 B.n720 B.n718 10.6151
R1700 B.n721 B.n720 10.6151
R1701 B.n722 B.n721 10.6151
R1702 B.n723 B.n722 10.6151
R1703 B.n725 B.n723 10.6151
R1704 B.n726 B.n725 10.6151
R1705 B.n727 B.n726 10.6151
R1706 B.n728 B.n727 10.6151
R1707 B.n730 B.n728 10.6151
R1708 B.n731 B.n730 10.6151
R1709 B.n732 B.n731 10.6151
R1710 B.n733 B.n732 10.6151
R1711 B.n735 B.n733 10.6151
R1712 B.n736 B.n735 10.6151
R1713 B.n737 B.n736 10.6151
R1714 B.n738 B.n737 10.6151
R1715 B.n740 B.n738 10.6151
R1716 B.n741 B.n740 10.6151
R1717 B.n742 B.n741 10.6151
R1718 B.n743 B.n742 10.6151
R1719 B.n745 B.n743 10.6151
R1720 B.n746 B.n745 10.6151
R1721 B.n747 B.n746 10.6151
R1722 B.n748 B.n747 10.6151
R1723 B.n750 B.n748 10.6151
R1724 B.n751 B.n750 10.6151
R1725 B.n752 B.n751 10.6151
R1726 B.n753 B.n752 10.6151
R1727 B.n755 B.n753 10.6151
R1728 B.n756 B.n755 10.6151
R1729 B.n757 B.n756 10.6151
R1730 B.n758 B.n757 10.6151
R1731 B.n760 B.n758 10.6151
R1732 B.n761 B.n760 10.6151
R1733 B.n762 B.n761 10.6151
R1734 B.n763 B.n762 10.6151
R1735 B.n765 B.n763 10.6151
R1736 B.n766 B.n765 10.6151
R1737 B.n767 B.n766 10.6151
R1738 B.n768 B.n767 10.6151
R1739 B.n769 B.n768 10.6151
R1740 B.n434 B.n364 10.6151
R1741 B.n429 B.n364 10.6151
R1742 B.n429 B.n428 10.6151
R1743 B.n428 B.n427 10.6151
R1744 B.n427 B.n424 10.6151
R1745 B.n424 B.n423 10.6151
R1746 B.n423 B.n420 10.6151
R1747 B.n418 B.n415 10.6151
R1748 B.n415 B.n414 10.6151
R1749 B.n414 B.n411 10.6151
R1750 B.n411 B.n410 10.6151
R1751 B.n410 B.n407 10.6151
R1752 B.n407 B.n406 10.6151
R1753 B.n406 B.n403 10.6151
R1754 B.n403 B.n402 10.6151
R1755 B.n402 B.n399 10.6151
R1756 B.n397 B.n394 10.6151
R1757 B.n394 B.n393 10.6151
R1758 B.n393 B.n390 10.6151
R1759 B.n390 B.n389 10.6151
R1760 B.n389 B.n386 10.6151
R1761 B.n386 B.n385 10.6151
R1762 B.n385 B.n383 10.6151
R1763 B.n436 B.n435 10.6151
R1764 B.n436 B.n356 10.6151
R1765 B.n446 B.n356 10.6151
R1766 B.n447 B.n446 10.6151
R1767 B.n448 B.n447 10.6151
R1768 B.n448 B.n348 10.6151
R1769 B.n458 B.n348 10.6151
R1770 B.n459 B.n458 10.6151
R1771 B.n460 B.n459 10.6151
R1772 B.n460 B.n340 10.6151
R1773 B.n469 B.n340 10.6151
R1774 B.n470 B.n469 10.6151
R1775 B.n471 B.n470 10.6151
R1776 B.n471 B.n332 10.6151
R1777 B.n481 B.n332 10.6151
R1778 B.n482 B.n481 10.6151
R1779 B.n483 B.n482 10.6151
R1780 B.n483 B.n324 10.6151
R1781 B.n493 B.n324 10.6151
R1782 B.n494 B.n493 10.6151
R1783 B.n495 B.n494 10.6151
R1784 B.n495 B.n316 10.6151
R1785 B.n506 B.n316 10.6151
R1786 B.n507 B.n506 10.6151
R1787 B.n508 B.n507 10.6151
R1788 B.n508 B.n309 10.6151
R1789 B.n518 B.n309 10.6151
R1790 B.n519 B.n518 10.6151
R1791 B.n520 B.n519 10.6151
R1792 B.n520 B.n301 10.6151
R1793 B.n530 B.n301 10.6151
R1794 B.n531 B.n530 10.6151
R1795 B.n532 B.n531 10.6151
R1796 B.n532 B.n293 10.6151
R1797 B.n542 B.n293 10.6151
R1798 B.n543 B.n542 10.6151
R1799 B.n544 B.n543 10.6151
R1800 B.n544 B.n285 10.6151
R1801 B.n554 B.n285 10.6151
R1802 B.n555 B.n554 10.6151
R1803 B.n556 B.n555 10.6151
R1804 B.n556 B.n277 10.6151
R1805 B.n566 B.n277 10.6151
R1806 B.n567 B.n566 10.6151
R1807 B.n568 B.n567 10.6151
R1808 B.n568 B.n269 10.6151
R1809 B.n578 B.n269 10.6151
R1810 B.n579 B.n578 10.6151
R1811 B.n580 B.n579 10.6151
R1812 B.n580 B.n261 10.6151
R1813 B.n590 B.n261 10.6151
R1814 B.n591 B.n590 10.6151
R1815 B.n592 B.n591 10.6151
R1816 B.n592 B.n253 10.6151
R1817 B.n602 B.n253 10.6151
R1818 B.n603 B.n602 10.6151
R1819 B.n604 B.n603 10.6151
R1820 B.n604 B.n245 10.6151
R1821 B.n614 B.n245 10.6151
R1822 B.n615 B.n614 10.6151
R1823 B.n616 B.n615 10.6151
R1824 B.n616 B.n237 10.6151
R1825 B.n626 B.n237 10.6151
R1826 B.n627 B.n626 10.6151
R1827 B.n628 B.n627 10.6151
R1828 B.n628 B.n229 10.6151
R1829 B.n638 B.n229 10.6151
R1830 B.n639 B.n638 10.6151
R1831 B.n640 B.n639 10.6151
R1832 B.n640 B.n221 10.6151
R1833 B.n650 B.n221 10.6151
R1834 B.n651 B.n650 10.6151
R1835 B.n652 B.n651 10.6151
R1836 B.n652 B.n213 10.6151
R1837 B.n663 B.n213 10.6151
R1838 B.n664 B.n663 10.6151
R1839 B.n665 B.n664 10.6151
R1840 B.n665 B.n0 10.6151
R1841 B.n929 B.n1 10.6151
R1842 B.n929 B.n928 10.6151
R1843 B.n928 B.n927 10.6151
R1844 B.n927 B.n10 10.6151
R1845 B.n921 B.n10 10.6151
R1846 B.n921 B.n920 10.6151
R1847 B.n920 B.n919 10.6151
R1848 B.n919 B.n17 10.6151
R1849 B.n913 B.n17 10.6151
R1850 B.n913 B.n912 10.6151
R1851 B.n912 B.n911 10.6151
R1852 B.n911 B.n24 10.6151
R1853 B.n905 B.n24 10.6151
R1854 B.n905 B.n904 10.6151
R1855 B.n904 B.n903 10.6151
R1856 B.n903 B.n31 10.6151
R1857 B.n897 B.n31 10.6151
R1858 B.n897 B.n896 10.6151
R1859 B.n896 B.n895 10.6151
R1860 B.n895 B.n38 10.6151
R1861 B.n889 B.n38 10.6151
R1862 B.n889 B.n888 10.6151
R1863 B.n888 B.n887 10.6151
R1864 B.n887 B.n45 10.6151
R1865 B.n881 B.n45 10.6151
R1866 B.n881 B.n880 10.6151
R1867 B.n880 B.n879 10.6151
R1868 B.n879 B.n52 10.6151
R1869 B.n873 B.n52 10.6151
R1870 B.n873 B.n872 10.6151
R1871 B.n872 B.n871 10.6151
R1872 B.n871 B.n59 10.6151
R1873 B.n865 B.n59 10.6151
R1874 B.n865 B.n864 10.6151
R1875 B.n864 B.n863 10.6151
R1876 B.n863 B.n66 10.6151
R1877 B.n857 B.n66 10.6151
R1878 B.n857 B.n856 10.6151
R1879 B.n856 B.n855 10.6151
R1880 B.n855 B.n73 10.6151
R1881 B.n849 B.n73 10.6151
R1882 B.n849 B.n848 10.6151
R1883 B.n848 B.n847 10.6151
R1884 B.n847 B.n80 10.6151
R1885 B.n841 B.n80 10.6151
R1886 B.n841 B.n840 10.6151
R1887 B.n840 B.n839 10.6151
R1888 B.n839 B.n87 10.6151
R1889 B.n833 B.n87 10.6151
R1890 B.n833 B.n832 10.6151
R1891 B.n832 B.n831 10.6151
R1892 B.n831 B.n94 10.6151
R1893 B.n825 B.n94 10.6151
R1894 B.n825 B.n824 10.6151
R1895 B.n824 B.n823 10.6151
R1896 B.n823 B.n100 10.6151
R1897 B.n817 B.n100 10.6151
R1898 B.n817 B.n816 10.6151
R1899 B.n816 B.n815 10.6151
R1900 B.n815 B.n108 10.6151
R1901 B.n809 B.n108 10.6151
R1902 B.n809 B.n808 10.6151
R1903 B.n808 B.n807 10.6151
R1904 B.n807 B.n115 10.6151
R1905 B.n801 B.n115 10.6151
R1906 B.n801 B.n800 10.6151
R1907 B.n800 B.n799 10.6151
R1908 B.n799 B.n122 10.6151
R1909 B.n794 B.n122 10.6151
R1910 B.n794 B.n793 10.6151
R1911 B.n793 B.n792 10.6151
R1912 B.n792 B.n129 10.6151
R1913 B.n786 B.n129 10.6151
R1914 B.n786 B.n785 10.6151
R1915 B.n785 B.n784 10.6151
R1916 B.n784 B.n136 10.6151
R1917 B.n778 B.n136 10.6151
R1918 B.n778 B.n777 10.6151
R1919 B.n174 B.n163 9.36635
R1920 B.n197 B.n160 9.36635
R1921 B.n420 B.n419 9.36635
R1922 B.n398 B.n397 9.36635
R1923 B.n503 B.t0 7.33995
R1924 B.n102 B.t8 7.33995
R1925 B.n935 B.n0 2.81026
R1926 B.n935 B.n1 2.81026
R1927 B.n177 B.n163 1.24928
R1928 B.n194 B.n160 1.24928
R1929 B.n419 B.n418 1.24928
R1930 B.n399 B.n398 1.24928
R1931 VN.n108 VN.n107 161.3
R1932 VN.n106 VN.n56 161.3
R1933 VN.n105 VN.n104 161.3
R1934 VN.n103 VN.n57 161.3
R1935 VN.n102 VN.n101 161.3
R1936 VN.n100 VN.n58 161.3
R1937 VN.n99 VN.n98 161.3
R1938 VN.n97 VN.n59 161.3
R1939 VN.n96 VN.n95 161.3
R1940 VN.n94 VN.n60 161.3
R1941 VN.n93 VN.n92 161.3
R1942 VN.n91 VN.n62 161.3
R1943 VN.n90 VN.n89 161.3
R1944 VN.n88 VN.n63 161.3
R1945 VN.n87 VN.n86 161.3
R1946 VN.n85 VN.n64 161.3
R1947 VN.n84 VN.n83 161.3
R1948 VN.n82 VN.n65 161.3
R1949 VN.n81 VN.n80 161.3
R1950 VN.n79 VN.n66 161.3
R1951 VN.n78 VN.n77 161.3
R1952 VN.n76 VN.n67 161.3
R1953 VN.n75 VN.n74 161.3
R1954 VN.n73 VN.n68 161.3
R1955 VN.n72 VN.n71 161.3
R1956 VN.n53 VN.n52 161.3
R1957 VN.n51 VN.n1 161.3
R1958 VN.n50 VN.n49 161.3
R1959 VN.n48 VN.n2 161.3
R1960 VN.n47 VN.n46 161.3
R1961 VN.n45 VN.n3 161.3
R1962 VN.n44 VN.n43 161.3
R1963 VN.n42 VN.n4 161.3
R1964 VN.n41 VN.n40 161.3
R1965 VN.n38 VN.n5 161.3
R1966 VN.n37 VN.n36 161.3
R1967 VN.n35 VN.n6 161.3
R1968 VN.n34 VN.n33 161.3
R1969 VN.n32 VN.n7 161.3
R1970 VN.n31 VN.n30 161.3
R1971 VN.n29 VN.n8 161.3
R1972 VN.n28 VN.n27 161.3
R1973 VN.n26 VN.n9 161.3
R1974 VN.n25 VN.n24 161.3
R1975 VN.n23 VN.n10 161.3
R1976 VN.n22 VN.n21 161.3
R1977 VN.n20 VN.n11 161.3
R1978 VN.n19 VN.n18 161.3
R1979 VN.n17 VN.n12 161.3
R1980 VN.n16 VN.n15 161.3
R1981 VN.n54 VN.n0 87.2945
R1982 VN.n109 VN.n55 87.2945
R1983 VN.n14 VN.n13 73.7075
R1984 VN.n70 VN.n69 73.7075
R1985 VN VN.n109 50.7443
R1986 VN.n46 VN.n2 44.9365
R1987 VN.n101 VN.n57 44.9365
R1988 VN.n21 VN.n20 42.0302
R1989 VN.n33 VN.n6 42.0302
R1990 VN.n77 VN.n76 42.0302
R1991 VN.n89 VN.n62 42.0302
R1992 VN.n21 VN.n10 39.1239
R1993 VN.n33 VN.n32 39.1239
R1994 VN.n77 VN.n66 39.1239
R1995 VN.n89 VN.n88 39.1239
R1996 VN.n69 VN.t4 36.6423
R1997 VN.n13 VN.t2 36.6423
R1998 VN.n46 VN.n45 36.2176
R1999 VN.n101 VN.n100 36.2176
R2000 VN.n15 VN.n12 24.5923
R2001 VN.n19 VN.n12 24.5923
R2002 VN.n20 VN.n19 24.5923
R2003 VN.n25 VN.n10 24.5923
R2004 VN.n26 VN.n25 24.5923
R2005 VN.n27 VN.n26 24.5923
R2006 VN.n27 VN.n8 24.5923
R2007 VN.n31 VN.n8 24.5923
R2008 VN.n32 VN.n31 24.5923
R2009 VN.n37 VN.n6 24.5923
R2010 VN.n38 VN.n37 24.5923
R2011 VN.n40 VN.n38 24.5923
R2012 VN.n44 VN.n4 24.5923
R2013 VN.n45 VN.n44 24.5923
R2014 VN.n50 VN.n2 24.5923
R2015 VN.n51 VN.n50 24.5923
R2016 VN.n52 VN.n51 24.5923
R2017 VN.n76 VN.n75 24.5923
R2018 VN.n75 VN.n68 24.5923
R2019 VN.n71 VN.n68 24.5923
R2020 VN.n88 VN.n87 24.5923
R2021 VN.n87 VN.n64 24.5923
R2022 VN.n83 VN.n64 24.5923
R2023 VN.n83 VN.n82 24.5923
R2024 VN.n82 VN.n81 24.5923
R2025 VN.n81 VN.n66 24.5923
R2026 VN.n100 VN.n99 24.5923
R2027 VN.n99 VN.n59 24.5923
R2028 VN.n95 VN.n94 24.5923
R2029 VN.n94 VN.n93 24.5923
R2030 VN.n93 VN.n62 24.5923
R2031 VN.n107 VN.n106 24.5923
R2032 VN.n106 VN.n105 24.5923
R2033 VN.n105 VN.n57 24.5923
R2034 VN.n39 VN.n4 23.1168
R2035 VN.n61 VN.n59 23.1168
R2036 VN.n27 VN.t9 4.69023
R2037 VN.n14 VN.t8 4.69023
R2038 VN.n39 VN.t7 4.69023
R2039 VN.n0 VN.t5 4.69023
R2040 VN.n83 VN.t0 4.69023
R2041 VN.n70 VN.t1 4.69023
R2042 VN.n61 VN.t3 4.69023
R2043 VN.n55 VN.t6 4.69023
R2044 VN.n72 VN.n69 3.36401
R2045 VN.n16 VN.n13 3.36401
R2046 VN.n52 VN.n0 2.95152
R2047 VN.n107 VN.n55 2.95152
R2048 VN.n15 VN.n14 1.47601
R2049 VN.n40 VN.n39 1.47601
R2050 VN.n71 VN.n70 1.47601
R2051 VN.n95 VN.n61 1.47601
R2052 VN.n109 VN.n108 0.354861
R2053 VN.n54 VN.n53 0.354861
R2054 VN VN.n54 0.267071
R2055 VN.n108 VN.n56 0.189894
R2056 VN.n104 VN.n56 0.189894
R2057 VN.n104 VN.n103 0.189894
R2058 VN.n103 VN.n102 0.189894
R2059 VN.n102 VN.n58 0.189894
R2060 VN.n98 VN.n58 0.189894
R2061 VN.n98 VN.n97 0.189894
R2062 VN.n97 VN.n96 0.189894
R2063 VN.n96 VN.n60 0.189894
R2064 VN.n92 VN.n60 0.189894
R2065 VN.n92 VN.n91 0.189894
R2066 VN.n91 VN.n90 0.189894
R2067 VN.n90 VN.n63 0.189894
R2068 VN.n86 VN.n63 0.189894
R2069 VN.n86 VN.n85 0.189894
R2070 VN.n85 VN.n84 0.189894
R2071 VN.n84 VN.n65 0.189894
R2072 VN.n80 VN.n65 0.189894
R2073 VN.n80 VN.n79 0.189894
R2074 VN.n79 VN.n78 0.189894
R2075 VN.n78 VN.n67 0.189894
R2076 VN.n74 VN.n67 0.189894
R2077 VN.n74 VN.n73 0.189894
R2078 VN.n73 VN.n72 0.189894
R2079 VN.n17 VN.n16 0.189894
R2080 VN.n18 VN.n17 0.189894
R2081 VN.n18 VN.n11 0.189894
R2082 VN.n22 VN.n11 0.189894
R2083 VN.n23 VN.n22 0.189894
R2084 VN.n24 VN.n23 0.189894
R2085 VN.n24 VN.n9 0.189894
R2086 VN.n28 VN.n9 0.189894
R2087 VN.n29 VN.n28 0.189894
R2088 VN.n30 VN.n29 0.189894
R2089 VN.n30 VN.n7 0.189894
R2090 VN.n34 VN.n7 0.189894
R2091 VN.n35 VN.n34 0.189894
R2092 VN.n36 VN.n35 0.189894
R2093 VN.n36 VN.n5 0.189894
R2094 VN.n41 VN.n5 0.189894
R2095 VN.n42 VN.n41 0.189894
R2096 VN.n43 VN.n42 0.189894
R2097 VN.n43 VN.n3 0.189894
R2098 VN.n47 VN.n3 0.189894
R2099 VN.n48 VN.n47 0.189894
R2100 VN.n49 VN.n48 0.189894
R2101 VN.n49 VN.n1 0.189894
R2102 VN.n53 VN.n1 0.189894
R2103 VDD2.n1 VDD2.t7 267.166
R2104 VDD2.n4 VDD2.t3 263.692
R2105 VDD2.n3 VDD2.n2 238.742
R2106 VDD2 VDD2.n7 238.738
R2107 VDD2.n6 VDD2.n5 236.191
R2108 VDD2.n1 VDD2.n0 236.191
R2109 VDD2.n4 VDD2.n3 40.8381
R2110 VDD2.n7 VDD2.t8 27.5005
R2111 VDD2.n7 VDD2.t5 27.5005
R2112 VDD2.n5 VDD2.t6 27.5005
R2113 VDD2.n5 VDD2.t9 27.5005
R2114 VDD2.n2 VDD2.t2 27.5005
R2115 VDD2.n2 VDD2.t4 27.5005
R2116 VDD2.n0 VDD2.t1 27.5005
R2117 VDD2.n0 VDD2.t0 27.5005
R2118 VDD2.n6 VDD2.n4 3.47464
R2119 VDD2 VDD2.n6 0.927224
R2120 VDD2.n3 VDD2.n1 0.813688
C0 VN VTAIL 3.54645f
C1 VDD2 VP 0.734721f
C2 VN VDD2 1.21955f
C3 VN VP 7.93492f
C4 VTAIL VDD1 6.514451f
C5 VDD2 VDD1 2.88799f
C6 VDD1 VP 1.78348f
C7 VDD2 VTAIL 6.57547f
C8 VN VDD1 0.164295f
C9 VTAIL VP 3.56058f
C10 VDD2 B 6.56543f
C11 VDD1 B 6.499499f
C12 VTAIL B 3.761964f
C13 VN B 22.725409f
C14 VP B 20.868464f
C15 VDD2.t7 B 0.090722f
C16 VDD2.t1 B 0.017864f
C17 VDD2.t0 B 0.017864f
C18 VDD2.n0 B 0.043919f
C19 VDD2.n1 B 0.961394f
C20 VDD2.t2 B 0.017864f
C21 VDD2.t4 B 0.017864f
C22 VDD2.n2 B 0.051426f
C23 VDD2.n3 B 3.35651f
C24 VDD2.t3 B 0.08484f
C25 VDD2.n4 B 3.10118f
C26 VDD2.t6 B 0.017864f
C27 VDD2.t9 B 0.017864f
C28 VDD2.n5 B 0.043919f
C29 VDD2.n6 B 0.525589f
C30 VDD2.t8 B 0.017864f
C31 VDD2.t5 B 0.017864f
C32 VDD2.n7 B 0.051412f
C33 VN.t5 B 0.116217f
C34 VN.n0 B 0.204092f
C35 VN.n1 B 0.028986f
C36 VN.n2 B 0.055674f
C37 VN.n3 B 0.028986f
C38 VN.n4 B 0.05216f
C39 VN.n5 B 0.028986f
C40 VN.n6 B 0.056835f
C41 VN.n7 B 0.028986f
C42 VN.n8 B 0.053752f
C43 VN.n9 B 0.028986f
C44 VN.t9 B 0.116217f
C45 VN.n10 B 0.057695f
C46 VN.n11 B 0.028986f
C47 VN.n12 B 0.053752f
C48 VN.t2 B 0.393351f
C49 VN.n13 B 0.272255f
C50 VN.t8 B 0.116217f
C51 VN.n14 B 0.190324f
C52 VN.n15 B 0.028808f
C53 VN.n16 B 0.368079f
C54 VN.n17 B 0.028986f
C55 VN.n18 B 0.028986f
C56 VN.n19 B 0.053752f
C57 VN.n20 B 0.056835f
C58 VN.n21 B 0.023494f
C59 VN.n22 B 0.028986f
C60 VN.n23 B 0.028986f
C61 VN.n24 B 0.028986f
C62 VN.n25 B 0.053752f
C63 VN.n26 B 0.053752f
C64 VN.n27 B 0.125887f
C65 VN.n28 B 0.028986f
C66 VN.n29 B 0.028986f
C67 VN.n30 B 0.028986f
C68 VN.n31 B 0.053752f
C69 VN.n32 B 0.057695f
C70 VN.n33 B 0.023494f
C71 VN.n34 B 0.028986f
C72 VN.n35 B 0.028986f
C73 VN.n36 B 0.028986f
C74 VN.n37 B 0.053752f
C75 VN.n38 B 0.053752f
C76 VN.t7 B 0.116217f
C77 VN.n39 B 0.098671f
C78 VN.n40 B 0.028808f
C79 VN.n41 B 0.028986f
C80 VN.n42 B 0.028986f
C81 VN.n43 B 0.028986f
C82 VN.n44 B 0.053752f
C83 VN.n45 B 0.058182f
C84 VN.n46 B 0.024168f
C85 VN.n47 B 0.028986f
C86 VN.n48 B 0.028986f
C87 VN.n49 B 0.028986f
C88 VN.n50 B 0.053752f
C89 VN.n51 B 0.053752f
C90 VN.n52 B 0.0304f
C91 VN.n53 B 0.046776f
C92 VN.n54 B 0.087267f
C93 VN.t6 B 0.116217f
C94 VN.n55 B 0.204092f
C95 VN.n56 B 0.028986f
C96 VN.n57 B 0.055674f
C97 VN.n58 B 0.028986f
C98 VN.n59 B 0.05216f
C99 VN.n60 B 0.028986f
C100 VN.t3 B 0.116217f
C101 VN.n61 B 0.098671f
C102 VN.n62 B 0.056835f
C103 VN.n63 B 0.028986f
C104 VN.n64 B 0.053752f
C105 VN.n65 B 0.028986f
C106 VN.t0 B 0.116217f
C107 VN.n66 B 0.057695f
C108 VN.n67 B 0.028986f
C109 VN.n68 B 0.053752f
C110 VN.t4 B 0.393351f
C111 VN.n69 B 0.272255f
C112 VN.t1 B 0.116217f
C113 VN.n70 B 0.190324f
C114 VN.n71 B 0.028808f
C115 VN.n72 B 0.368079f
C116 VN.n73 B 0.028986f
C117 VN.n74 B 0.028986f
C118 VN.n75 B 0.053752f
C119 VN.n76 B 0.056835f
C120 VN.n77 B 0.023494f
C121 VN.n78 B 0.028986f
C122 VN.n79 B 0.028986f
C123 VN.n80 B 0.028986f
C124 VN.n81 B 0.053752f
C125 VN.n82 B 0.053752f
C126 VN.n83 B 0.125887f
C127 VN.n84 B 0.028986f
C128 VN.n85 B 0.028986f
C129 VN.n86 B 0.028986f
C130 VN.n87 B 0.053752f
C131 VN.n88 B 0.057695f
C132 VN.n89 B 0.023494f
C133 VN.n90 B 0.028986f
C134 VN.n91 B 0.028986f
C135 VN.n92 B 0.028986f
C136 VN.n93 B 0.053752f
C137 VN.n94 B 0.053752f
C138 VN.n95 B 0.028808f
C139 VN.n96 B 0.028986f
C140 VN.n97 B 0.028986f
C141 VN.n98 B 0.028986f
C142 VN.n99 B 0.053752f
C143 VN.n100 B 0.058182f
C144 VN.n101 B 0.024168f
C145 VN.n102 B 0.028986f
C146 VN.n103 B 0.028986f
C147 VN.n104 B 0.028986f
C148 VN.n105 B 0.053752f
C149 VN.n106 B 0.053752f
C150 VN.n107 B 0.0304f
C151 VN.n108 B 0.046776f
C152 VN.n109 B 1.7046f
C153 VTAIL.t4 B 0.029965f
C154 VTAIL.t7 B 0.029965f
C155 VTAIL.n0 B 0.064189f
C156 VTAIL.n1 B 0.89924f
C157 VTAIL.t18 B 0.133002f
C158 VTAIL.n2 B 1.04966f
C159 VTAIL.t17 B 0.029965f
C160 VTAIL.t11 B 0.029965f
C161 VTAIL.n3 B 0.064189f
C162 VTAIL.n4 B 1.2518f
C163 VTAIL.t16 B 0.029965f
C164 VTAIL.t13 B 0.029965f
C165 VTAIL.n5 B 0.064189f
C166 VTAIL.n6 B 2.66208f
C167 VTAIL.t0 B 0.029965f
C168 VTAIL.t5 B 0.029965f
C169 VTAIL.n7 B 0.064189f
C170 VTAIL.n8 B 2.66208f
C171 VTAIL.t1 B 0.029965f
C172 VTAIL.t2 B 0.029965f
C173 VTAIL.n9 B 0.064189f
C174 VTAIL.n10 B 1.2518f
C175 VTAIL.t6 B 0.133002f
C176 VTAIL.n11 B 1.04966f
C177 VTAIL.t14 B 0.029965f
C178 VTAIL.t19 B 0.029965f
C179 VTAIL.n12 B 0.064189f
C180 VTAIL.n13 B 1.03675f
C181 VTAIL.t15 B 0.029965f
C182 VTAIL.t10 B 0.029965f
C183 VTAIL.n14 B 0.064189f
C184 VTAIL.n15 B 1.2518f
C185 VTAIL.t12 B 0.133002f
C186 VTAIL.n16 B 2.08543f
C187 VTAIL.t8 B 0.133002f
C188 VTAIL.n17 B 2.08543f
C189 VTAIL.t3 B 0.029965f
C190 VTAIL.t9 B 0.029965f
C191 VTAIL.n18 B 0.064189f
C192 VTAIL.n19 B 0.799762f
C193 VDD1.t4 B 0.088684f
C194 VDD1.t5 B 0.017463f
C195 VDD1.t2 B 0.017463f
C196 VDD1.n0 B 0.042933f
C197 VDD1.n1 B 0.950156f
C198 VDD1.t6 B 0.088684f
C199 VDD1.t8 B 0.017463f
C200 VDD1.t1 B 0.017463f
C201 VDD1.n2 B 0.042933f
C202 VDD1.n3 B 0.939802f
C203 VDD1.t3 B 0.017463f
C204 VDD1.t9 B 0.017463f
C205 VDD1.n4 B 0.050271f
C206 VDD1.n5 B 3.45708f
C207 VDD1.t0 B 0.017463f
C208 VDD1.t7 B 0.017463f
C209 VDD1.n6 B 0.042933f
C210 VDD1.n7 B 3.21325f
C211 VP.t1 B 0.117657f
C212 VP.n0 B 0.20662f
C213 VP.n1 B 0.029345f
C214 VP.n2 B 0.056364f
C215 VP.n3 B 0.029345f
C216 VP.n4 B 0.052806f
C217 VP.n5 B 0.029345f
C218 VP.n6 B 0.057539f
C219 VP.n7 B 0.029345f
C220 VP.n8 B 0.054418f
C221 VP.n9 B 0.029345f
C222 VP.t2 B 0.117657f
C223 VP.n10 B 0.05841f
C224 VP.n11 B 0.029345f
C225 VP.n12 B 0.054418f
C226 VP.n13 B 0.029345f
C227 VP.t6 B 0.117657f
C228 VP.n14 B 0.058902f
C229 VP.n15 B 0.029345f
C230 VP.n16 B 0.054418f
C231 VP.t7 B 0.117657f
C232 VP.n17 B 0.20662f
C233 VP.n18 B 0.029345f
C234 VP.n19 B 0.056364f
C235 VP.n20 B 0.029345f
C236 VP.n21 B 0.052806f
C237 VP.n22 B 0.029345f
C238 VP.n23 B 0.057539f
C239 VP.n24 B 0.029345f
C240 VP.n25 B 0.054418f
C241 VP.n26 B 0.029345f
C242 VP.t4 B 0.117657f
C243 VP.n27 B 0.05841f
C244 VP.n28 B 0.029345f
C245 VP.n29 B 0.054418f
C246 VP.t5 B 0.398224f
C247 VP.n30 B 0.275628f
C248 VP.t0 B 0.117657f
C249 VP.n31 B 0.192682f
C250 VP.n32 B 0.029165f
C251 VP.n33 B 0.372641f
C252 VP.n34 B 0.029345f
C253 VP.n35 B 0.029345f
C254 VP.n36 B 0.054418f
C255 VP.n37 B 0.057539f
C256 VP.n38 B 0.023785f
C257 VP.n39 B 0.029345f
C258 VP.n40 B 0.029345f
C259 VP.n41 B 0.029345f
C260 VP.n42 B 0.054418f
C261 VP.n43 B 0.054418f
C262 VP.n44 B 0.127447f
C263 VP.n45 B 0.029345f
C264 VP.n46 B 0.029345f
C265 VP.n47 B 0.029345f
C266 VP.n48 B 0.054418f
C267 VP.n49 B 0.05841f
C268 VP.n50 B 0.023785f
C269 VP.n51 B 0.029345f
C270 VP.n52 B 0.029345f
C271 VP.n53 B 0.029345f
C272 VP.n54 B 0.054418f
C273 VP.n55 B 0.054418f
C274 VP.t9 B 0.117657f
C275 VP.n56 B 0.099894f
C276 VP.n57 B 0.029165f
C277 VP.n58 B 0.029345f
C278 VP.n59 B 0.029345f
C279 VP.n60 B 0.029345f
C280 VP.n61 B 0.054418f
C281 VP.n62 B 0.058902f
C282 VP.n63 B 0.024468f
C283 VP.n64 B 0.029345f
C284 VP.n65 B 0.029345f
C285 VP.n66 B 0.029345f
C286 VP.n67 B 0.054418f
C287 VP.n68 B 0.054418f
C288 VP.n69 B 0.030777f
C289 VP.n70 B 0.047355f
C290 VP.n71 B 1.71376f
C291 VP.n72 B 1.73468f
C292 VP.t3 B 0.117657f
C293 VP.n73 B 0.20662f
C294 VP.n74 B 0.030777f
C295 VP.n75 B 0.047355f
C296 VP.n76 B 0.029345f
C297 VP.n77 B 0.029345f
C298 VP.n78 B 0.054418f
C299 VP.n79 B 0.056364f
C300 VP.n80 B 0.024468f
C301 VP.n81 B 0.029345f
C302 VP.n82 B 0.029345f
C303 VP.n83 B 0.029345f
C304 VP.n84 B 0.054418f
C305 VP.n85 B 0.052806f
C306 VP.n86 B 0.099894f
C307 VP.n87 B 0.029165f
C308 VP.n88 B 0.029345f
C309 VP.n89 B 0.029345f
C310 VP.n90 B 0.029345f
C311 VP.n91 B 0.054418f
C312 VP.n92 B 0.057539f
C313 VP.n93 B 0.023785f
C314 VP.n94 B 0.029345f
C315 VP.n95 B 0.029345f
C316 VP.n96 B 0.029345f
C317 VP.n97 B 0.054418f
C318 VP.n98 B 0.054418f
C319 VP.n99 B 0.127447f
C320 VP.n100 B 0.029345f
C321 VP.n101 B 0.029345f
C322 VP.n102 B 0.029345f
C323 VP.n103 B 0.054418f
C324 VP.n104 B 0.05841f
C325 VP.n105 B 0.023785f
C326 VP.n106 B 0.029345f
C327 VP.n107 B 0.029345f
C328 VP.n108 B 0.029345f
C329 VP.n109 B 0.054418f
C330 VP.n110 B 0.054418f
C331 VP.t8 B 0.117657f
C332 VP.n111 B 0.099894f
C333 VP.n112 B 0.029165f
C334 VP.n113 B 0.029345f
C335 VP.n114 B 0.029345f
C336 VP.n115 B 0.029345f
C337 VP.n116 B 0.054418f
C338 VP.n117 B 0.058902f
C339 VP.n118 B 0.024468f
C340 VP.n119 B 0.029345f
C341 VP.n120 B 0.029345f
C342 VP.n121 B 0.029345f
C343 VP.n122 B 0.054418f
C344 VP.n123 B 0.054418f
C345 VP.n124 B 0.030777f
C346 VP.n125 B 0.047355f
C347 VP.n126 B 0.088349f
.ends

