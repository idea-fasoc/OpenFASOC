* NGSPICE file created from diff_pair_sample_0501.ext - technology: sky130A

.subckt diff_pair_sample_0501 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0 ps=0 w=1.12 l=2.87
X1 VDD1.t5 VP.t0 VTAIL.t7 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0.1848 ps=1.45 w=1.12 l=2.87
X2 VTAIL.t9 VP.t1 VDD1.t4 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.1848 ps=1.45 w=1.12 l=2.87
X3 VDD2.t5 VN.t0 VTAIL.t11 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0.1848 ps=1.45 w=1.12 l=2.87
X4 VTAIL.t2 VN.t1 VDD2.t4 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.1848 ps=1.45 w=1.12 l=2.87
X5 VDD1.t3 VP.t2 VTAIL.t5 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.4368 ps=3.02 w=1.12 l=2.87
X6 VDD1.t2 VP.t3 VTAIL.t10 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.4368 ps=3.02 w=1.12 l=2.87
X7 B.t8 B.t6 B.t7 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0 ps=0 w=1.12 l=2.87
X8 VDD2.t3 VN.t2 VTAIL.t0 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.4368 ps=3.02 w=1.12 l=2.87
X9 VDD2.t2 VN.t3 VTAIL.t1 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.4368 ps=3.02 w=1.12 l=2.87
X10 VTAIL.t8 VP.t4 VDD1.t1 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.1848 ps=1.45 w=1.12 l=2.87
X11 VDD1.t0 VP.t5 VTAIL.t6 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0.1848 ps=1.45 w=1.12 l=2.87
X12 VTAIL.t4 VN.t4 VDD2.t1 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.1848 ps=1.45 w=1.12 l=2.87
X13 B.t5 B.t3 B.t4 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0 ps=0 w=1.12 l=2.87
X14 B.t2 B.t0 B.t1 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0 ps=0 w=1.12 l=2.87
X15 VDD2.t0 VN.t5 VTAIL.t3 w_n3530_n1192# sky130_fd_pr__pfet_01v8 ad=0.4368 pd=3.02 as=0.1848 ps=1.45 w=1.12 l=2.87
R0 B.n241 B.n240 585
R1 B.n239 B.n90 585
R2 B.n238 B.n237 585
R3 B.n236 B.n91 585
R4 B.n235 B.n234 585
R5 B.n233 B.n92 585
R6 B.n232 B.n231 585
R7 B.n230 B.n93 585
R8 B.n229 B.n228 585
R9 B.n227 B.n94 585
R10 B.n226 B.n225 585
R11 B.n221 B.n95 585
R12 B.n220 B.n219 585
R13 B.n218 B.n96 585
R14 B.n217 B.n216 585
R15 B.n215 B.n97 585
R16 B.n214 B.n213 585
R17 B.n212 B.n98 585
R18 B.n211 B.n210 585
R19 B.n208 B.n99 585
R20 B.n207 B.n206 585
R21 B.n205 B.n102 585
R22 B.n204 B.n203 585
R23 B.n202 B.n103 585
R24 B.n201 B.n200 585
R25 B.n199 B.n104 585
R26 B.n198 B.n197 585
R27 B.n196 B.n105 585
R28 B.n195 B.n194 585
R29 B.n242 B.n89 585
R30 B.n244 B.n243 585
R31 B.n245 B.n88 585
R32 B.n247 B.n246 585
R33 B.n248 B.n87 585
R34 B.n250 B.n249 585
R35 B.n251 B.n86 585
R36 B.n253 B.n252 585
R37 B.n254 B.n85 585
R38 B.n256 B.n255 585
R39 B.n257 B.n84 585
R40 B.n259 B.n258 585
R41 B.n260 B.n83 585
R42 B.n262 B.n261 585
R43 B.n263 B.n82 585
R44 B.n265 B.n264 585
R45 B.n266 B.n81 585
R46 B.n268 B.n267 585
R47 B.n269 B.n80 585
R48 B.n271 B.n270 585
R49 B.n272 B.n79 585
R50 B.n274 B.n273 585
R51 B.n275 B.n78 585
R52 B.n277 B.n276 585
R53 B.n278 B.n77 585
R54 B.n280 B.n279 585
R55 B.n281 B.n76 585
R56 B.n283 B.n282 585
R57 B.n284 B.n75 585
R58 B.n286 B.n285 585
R59 B.n287 B.n74 585
R60 B.n289 B.n288 585
R61 B.n290 B.n73 585
R62 B.n292 B.n291 585
R63 B.n293 B.n72 585
R64 B.n295 B.n294 585
R65 B.n296 B.n71 585
R66 B.n298 B.n297 585
R67 B.n299 B.n70 585
R68 B.n301 B.n300 585
R69 B.n302 B.n69 585
R70 B.n304 B.n303 585
R71 B.n305 B.n68 585
R72 B.n307 B.n306 585
R73 B.n308 B.n67 585
R74 B.n310 B.n309 585
R75 B.n311 B.n66 585
R76 B.n313 B.n312 585
R77 B.n314 B.n65 585
R78 B.n316 B.n315 585
R79 B.n317 B.n64 585
R80 B.n319 B.n318 585
R81 B.n320 B.n63 585
R82 B.n322 B.n321 585
R83 B.n323 B.n62 585
R84 B.n325 B.n324 585
R85 B.n326 B.n61 585
R86 B.n328 B.n327 585
R87 B.n329 B.n60 585
R88 B.n331 B.n330 585
R89 B.n332 B.n59 585
R90 B.n334 B.n333 585
R91 B.n335 B.n58 585
R92 B.n337 B.n336 585
R93 B.n338 B.n57 585
R94 B.n340 B.n339 585
R95 B.n341 B.n56 585
R96 B.n343 B.n342 585
R97 B.n344 B.n55 585
R98 B.n346 B.n345 585
R99 B.n347 B.n54 585
R100 B.n349 B.n348 585
R101 B.n350 B.n53 585
R102 B.n352 B.n351 585
R103 B.n353 B.n52 585
R104 B.n355 B.n354 585
R105 B.n356 B.n51 585
R106 B.n358 B.n357 585
R107 B.n359 B.n50 585
R108 B.n361 B.n360 585
R109 B.n362 B.n49 585
R110 B.n364 B.n363 585
R111 B.n365 B.n48 585
R112 B.n367 B.n366 585
R113 B.n368 B.n47 585
R114 B.n370 B.n369 585
R115 B.n371 B.n46 585
R116 B.n373 B.n372 585
R117 B.n374 B.n45 585
R118 B.n376 B.n375 585
R119 B.n377 B.n44 585
R120 B.n379 B.n378 585
R121 B.n424 B.n423 585
R122 B.n422 B.n25 585
R123 B.n421 B.n420 585
R124 B.n419 B.n26 585
R125 B.n418 B.n417 585
R126 B.n416 B.n27 585
R127 B.n415 B.n414 585
R128 B.n413 B.n28 585
R129 B.n412 B.n411 585
R130 B.n410 B.n29 585
R131 B.n408 B.n407 585
R132 B.n406 B.n32 585
R133 B.n405 B.n404 585
R134 B.n403 B.n33 585
R135 B.n402 B.n401 585
R136 B.n400 B.n34 585
R137 B.n399 B.n398 585
R138 B.n397 B.n35 585
R139 B.n396 B.n395 585
R140 B.n394 B.n393 585
R141 B.n392 B.n39 585
R142 B.n391 B.n390 585
R143 B.n389 B.n40 585
R144 B.n388 B.n387 585
R145 B.n386 B.n41 585
R146 B.n385 B.n384 585
R147 B.n383 B.n42 585
R148 B.n382 B.n381 585
R149 B.n380 B.n43 585
R150 B.n425 B.n24 585
R151 B.n427 B.n426 585
R152 B.n428 B.n23 585
R153 B.n430 B.n429 585
R154 B.n431 B.n22 585
R155 B.n433 B.n432 585
R156 B.n434 B.n21 585
R157 B.n436 B.n435 585
R158 B.n437 B.n20 585
R159 B.n439 B.n438 585
R160 B.n440 B.n19 585
R161 B.n442 B.n441 585
R162 B.n443 B.n18 585
R163 B.n445 B.n444 585
R164 B.n446 B.n17 585
R165 B.n448 B.n447 585
R166 B.n449 B.n16 585
R167 B.n451 B.n450 585
R168 B.n452 B.n15 585
R169 B.n454 B.n453 585
R170 B.n455 B.n14 585
R171 B.n457 B.n456 585
R172 B.n458 B.n13 585
R173 B.n460 B.n459 585
R174 B.n461 B.n12 585
R175 B.n463 B.n462 585
R176 B.n464 B.n11 585
R177 B.n466 B.n465 585
R178 B.n467 B.n10 585
R179 B.n469 B.n468 585
R180 B.n470 B.n9 585
R181 B.n472 B.n471 585
R182 B.n473 B.n8 585
R183 B.n475 B.n474 585
R184 B.n476 B.n7 585
R185 B.n478 B.n477 585
R186 B.n479 B.n6 585
R187 B.n481 B.n480 585
R188 B.n482 B.n5 585
R189 B.n484 B.n483 585
R190 B.n485 B.n4 585
R191 B.n487 B.n486 585
R192 B.n488 B.n3 585
R193 B.n490 B.n489 585
R194 B.n491 B.n0 585
R195 B.n2 B.n1 585
R196 B.n129 B.n128 585
R197 B.n130 B.n127 585
R198 B.n132 B.n131 585
R199 B.n133 B.n126 585
R200 B.n135 B.n134 585
R201 B.n136 B.n125 585
R202 B.n138 B.n137 585
R203 B.n139 B.n124 585
R204 B.n141 B.n140 585
R205 B.n142 B.n123 585
R206 B.n144 B.n143 585
R207 B.n145 B.n122 585
R208 B.n147 B.n146 585
R209 B.n148 B.n121 585
R210 B.n150 B.n149 585
R211 B.n151 B.n120 585
R212 B.n153 B.n152 585
R213 B.n154 B.n119 585
R214 B.n156 B.n155 585
R215 B.n157 B.n118 585
R216 B.n159 B.n158 585
R217 B.n160 B.n117 585
R218 B.n162 B.n161 585
R219 B.n163 B.n116 585
R220 B.n165 B.n164 585
R221 B.n166 B.n115 585
R222 B.n168 B.n167 585
R223 B.n169 B.n114 585
R224 B.n171 B.n170 585
R225 B.n172 B.n113 585
R226 B.n174 B.n173 585
R227 B.n175 B.n112 585
R228 B.n177 B.n176 585
R229 B.n178 B.n111 585
R230 B.n180 B.n179 585
R231 B.n181 B.n110 585
R232 B.n183 B.n182 585
R233 B.n184 B.n109 585
R234 B.n186 B.n185 585
R235 B.n187 B.n108 585
R236 B.n189 B.n188 585
R237 B.n190 B.n107 585
R238 B.n192 B.n191 585
R239 B.n193 B.n106 585
R240 B.n194 B.n193 526.135
R241 B.n240 B.n89 526.135
R242 B.n378 B.n43 526.135
R243 B.n425 B.n424 526.135
R244 B.n100 B.t10 425.587
R245 B.n222 B.t7 425.587
R246 B.n36 B.t2 425.587
R247 B.n30 B.t5 425.587
R248 B.n101 B.t11 363.526
R249 B.n223 B.t8 363.526
R250 B.n37 B.t1 363.526
R251 B.n31 B.t4 363.526
R252 B.n493 B.n492 256.663
R253 B.n492 B.n491 235.042
R254 B.n492 B.n2 235.042
R255 B.n100 B.t9 209.167
R256 B.n222 B.t6 209.167
R257 B.n36 B.t0 209.167
R258 B.n30 B.t3 209.167
R259 B.n194 B.n105 163.367
R260 B.n198 B.n105 163.367
R261 B.n199 B.n198 163.367
R262 B.n200 B.n199 163.367
R263 B.n200 B.n103 163.367
R264 B.n204 B.n103 163.367
R265 B.n205 B.n204 163.367
R266 B.n206 B.n205 163.367
R267 B.n206 B.n99 163.367
R268 B.n211 B.n99 163.367
R269 B.n212 B.n211 163.367
R270 B.n213 B.n212 163.367
R271 B.n213 B.n97 163.367
R272 B.n217 B.n97 163.367
R273 B.n218 B.n217 163.367
R274 B.n219 B.n218 163.367
R275 B.n219 B.n95 163.367
R276 B.n226 B.n95 163.367
R277 B.n227 B.n226 163.367
R278 B.n228 B.n227 163.367
R279 B.n228 B.n93 163.367
R280 B.n232 B.n93 163.367
R281 B.n233 B.n232 163.367
R282 B.n234 B.n233 163.367
R283 B.n234 B.n91 163.367
R284 B.n238 B.n91 163.367
R285 B.n239 B.n238 163.367
R286 B.n240 B.n239 163.367
R287 B.n378 B.n377 163.367
R288 B.n377 B.n376 163.367
R289 B.n376 B.n45 163.367
R290 B.n372 B.n45 163.367
R291 B.n372 B.n371 163.367
R292 B.n371 B.n370 163.367
R293 B.n370 B.n47 163.367
R294 B.n366 B.n47 163.367
R295 B.n366 B.n365 163.367
R296 B.n365 B.n364 163.367
R297 B.n364 B.n49 163.367
R298 B.n360 B.n49 163.367
R299 B.n360 B.n359 163.367
R300 B.n359 B.n358 163.367
R301 B.n358 B.n51 163.367
R302 B.n354 B.n51 163.367
R303 B.n354 B.n353 163.367
R304 B.n353 B.n352 163.367
R305 B.n352 B.n53 163.367
R306 B.n348 B.n53 163.367
R307 B.n348 B.n347 163.367
R308 B.n347 B.n346 163.367
R309 B.n346 B.n55 163.367
R310 B.n342 B.n55 163.367
R311 B.n342 B.n341 163.367
R312 B.n341 B.n340 163.367
R313 B.n340 B.n57 163.367
R314 B.n336 B.n57 163.367
R315 B.n336 B.n335 163.367
R316 B.n335 B.n334 163.367
R317 B.n334 B.n59 163.367
R318 B.n330 B.n59 163.367
R319 B.n330 B.n329 163.367
R320 B.n329 B.n328 163.367
R321 B.n328 B.n61 163.367
R322 B.n324 B.n61 163.367
R323 B.n324 B.n323 163.367
R324 B.n323 B.n322 163.367
R325 B.n322 B.n63 163.367
R326 B.n318 B.n63 163.367
R327 B.n318 B.n317 163.367
R328 B.n317 B.n316 163.367
R329 B.n316 B.n65 163.367
R330 B.n312 B.n65 163.367
R331 B.n312 B.n311 163.367
R332 B.n311 B.n310 163.367
R333 B.n310 B.n67 163.367
R334 B.n306 B.n67 163.367
R335 B.n306 B.n305 163.367
R336 B.n305 B.n304 163.367
R337 B.n304 B.n69 163.367
R338 B.n300 B.n69 163.367
R339 B.n300 B.n299 163.367
R340 B.n299 B.n298 163.367
R341 B.n298 B.n71 163.367
R342 B.n294 B.n71 163.367
R343 B.n294 B.n293 163.367
R344 B.n293 B.n292 163.367
R345 B.n292 B.n73 163.367
R346 B.n288 B.n73 163.367
R347 B.n288 B.n287 163.367
R348 B.n287 B.n286 163.367
R349 B.n286 B.n75 163.367
R350 B.n282 B.n75 163.367
R351 B.n282 B.n281 163.367
R352 B.n281 B.n280 163.367
R353 B.n280 B.n77 163.367
R354 B.n276 B.n77 163.367
R355 B.n276 B.n275 163.367
R356 B.n275 B.n274 163.367
R357 B.n274 B.n79 163.367
R358 B.n270 B.n79 163.367
R359 B.n270 B.n269 163.367
R360 B.n269 B.n268 163.367
R361 B.n268 B.n81 163.367
R362 B.n264 B.n81 163.367
R363 B.n264 B.n263 163.367
R364 B.n263 B.n262 163.367
R365 B.n262 B.n83 163.367
R366 B.n258 B.n83 163.367
R367 B.n258 B.n257 163.367
R368 B.n257 B.n256 163.367
R369 B.n256 B.n85 163.367
R370 B.n252 B.n85 163.367
R371 B.n252 B.n251 163.367
R372 B.n251 B.n250 163.367
R373 B.n250 B.n87 163.367
R374 B.n246 B.n87 163.367
R375 B.n246 B.n245 163.367
R376 B.n245 B.n244 163.367
R377 B.n244 B.n89 163.367
R378 B.n424 B.n25 163.367
R379 B.n420 B.n25 163.367
R380 B.n420 B.n419 163.367
R381 B.n419 B.n418 163.367
R382 B.n418 B.n27 163.367
R383 B.n414 B.n27 163.367
R384 B.n414 B.n413 163.367
R385 B.n413 B.n412 163.367
R386 B.n412 B.n29 163.367
R387 B.n407 B.n29 163.367
R388 B.n407 B.n406 163.367
R389 B.n406 B.n405 163.367
R390 B.n405 B.n33 163.367
R391 B.n401 B.n33 163.367
R392 B.n401 B.n400 163.367
R393 B.n400 B.n399 163.367
R394 B.n399 B.n35 163.367
R395 B.n395 B.n35 163.367
R396 B.n395 B.n394 163.367
R397 B.n394 B.n39 163.367
R398 B.n390 B.n39 163.367
R399 B.n390 B.n389 163.367
R400 B.n389 B.n388 163.367
R401 B.n388 B.n41 163.367
R402 B.n384 B.n41 163.367
R403 B.n384 B.n383 163.367
R404 B.n383 B.n382 163.367
R405 B.n382 B.n43 163.367
R406 B.n426 B.n425 163.367
R407 B.n426 B.n23 163.367
R408 B.n430 B.n23 163.367
R409 B.n431 B.n430 163.367
R410 B.n432 B.n431 163.367
R411 B.n432 B.n21 163.367
R412 B.n436 B.n21 163.367
R413 B.n437 B.n436 163.367
R414 B.n438 B.n437 163.367
R415 B.n438 B.n19 163.367
R416 B.n442 B.n19 163.367
R417 B.n443 B.n442 163.367
R418 B.n444 B.n443 163.367
R419 B.n444 B.n17 163.367
R420 B.n448 B.n17 163.367
R421 B.n449 B.n448 163.367
R422 B.n450 B.n449 163.367
R423 B.n450 B.n15 163.367
R424 B.n454 B.n15 163.367
R425 B.n455 B.n454 163.367
R426 B.n456 B.n455 163.367
R427 B.n456 B.n13 163.367
R428 B.n460 B.n13 163.367
R429 B.n461 B.n460 163.367
R430 B.n462 B.n461 163.367
R431 B.n462 B.n11 163.367
R432 B.n466 B.n11 163.367
R433 B.n467 B.n466 163.367
R434 B.n468 B.n467 163.367
R435 B.n468 B.n9 163.367
R436 B.n472 B.n9 163.367
R437 B.n473 B.n472 163.367
R438 B.n474 B.n473 163.367
R439 B.n474 B.n7 163.367
R440 B.n478 B.n7 163.367
R441 B.n479 B.n478 163.367
R442 B.n480 B.n479 163.367
R443 B.n480 B.n5 163.367
R444 B.n484 B.n5 163.367
R445 B.n485 B.n484 163.367
R446 B.n486 B.n485 163.367
R447 B.n486 B.n3 163.367
R448 B.n490 B.n3 163.367
R449 B.n491 B.n490 163.367
R450 B.n128 B.n2 163.367
R451 B.n128 B.n127 163.367
R452 B.n132 B.n127 163.367
R453 B.n133 B.n132 163.367
R454 B.n134 B.n133 163.367
R455 B.n134 B.n125 163.367
R456 B.n138 B.n125 163.367
R457 B.n139 B.n138 163.367
R458 B.n140 B.n139 163.367
R459 B.n140 B.n123 163.367
R460 B.n144 B.n123 163.367
R461 B.n145 B.n144 163.367
R462 B.n146 B.n145 163.367
R463 B.n146 B.n121 163.367
R464 B.n150 B.n121 163.367
R465 B.n151 B.n150 163.367
R466 B.n152 B.n151 163.367
R467 B.n152 B.n119 163.367
R468 B.n156 B.n119 163.367
R469 B.n157 B.n156 163.367
R470 B.n158 B.n157 163.367
R471 B.n158 B.n117 163.367
R472 B.n162 B.n117 163.367
R473 B.n163 B.n162 163.367
R474 B.n164 B.n163 163.367
R475 B.n164 B.n115 163.367
R476 B.n168 B.n115 163.367
R477 B.n169 B.n168 163.367
R478 B.n170 B.n169 163.367
R479 B.n170 B.n113 163.367
R480 B.n174 B.n113 163.367
R481 B.n175 B.n174 163.367
R482 B.n176 B.n175 163.367
R483 B.n176 B.n111 163.367
R484 B.n180 B.n111 163.367
R485 B.n181 B.n180 163.367
R486 B.n182 B.n181 163.367
R487 B.n182 B.n109 163.367
R488 B.n186 B.n109 163.367
R489 B.n187 B.n186 163.367
R490 B.n188 B.n187 163.367
R491 B.n188 B.n107 163.367
R492 B.n192 B.n107 163.367
R493 B.n193 B.n192 163.367
R494 B.n101 B.n100 62.0611
R495 B.n223 B.n222 62.0611
R496 B.n37 B.n36 62.0611
R497 B.n31 B.n30 62.0611
R498 B.n209 B.n101 59.5399
R499 B.n224 B.n223 59.5399
R500 B.n38 B.n37 59.5399
R501 B.n409 B.n31 59.5399
R502 B.n423 B.n24 34.1859
R503 B.n380 B.n379 34.1859
R504 B.n242 B.n241 34.1859
R505 B.n195 B.n106 34.1859
R506 B B.n493 18.0485
R507 B.n427 B.n24 10.6151
R508 B.n428 B.n427 10.6151
R509 B.n429 B.n428 10.6151
R510 B.n429 B.n22 10.6151
R511 B.n433 B.n22 10.6151
R512 B.n434 B.n433 10.6151
R513 B.n435 B.n434 10.6151
R514 B.n435 B.n20 10.6151
R515 B.n439 B.n20 10.6151
R516 B.n440 B.n439 10.6151
R517 B.n441 B.n440 10.6151
R518 B.n441 B.n18 10.6151
R519 B.n445 B.n18 10.6151
R520 B.n446 B.n445 10.6151
R521 B.n447 B.n446 10.6151
R522 B.n447 B.n16 10.6151
R523 B.n451 B.n16 10.6151
R524 B.n452 B.n451 10.6151
R525 B.n453 B.n452 10.6151
R526 B.n453 B.n14 10.6151
R527 B.n457 B.n14 10.6151
R528 B.n458 B.n457 10.6151
R529 B.n459 B.n458 10.6151
R530 B.n459 B.n12 10.6151
R531 B.n463 B.n12 10.6151
R532 B.n464 B.n463 10.6151
R533 B.n465 B.n464 10.6151
R534 B.n465 B.n10 10.6151
R535 B.n469 B.n10 10.6151
R536 B.n470 B.n469 10.6151
R537 B.n471 B.n470 10.6151
R538 B.n471 B.n8 10.6151
R539 B.n475 B.n8 10.6151
R540 B.n476 B.n475 10.6151
R541 B.n477 B.n476 10.6151
R542 B.n477 B.n6 10.6151
R543 B.n481 B.n6 10.6151
R544 B.n482 B.n481 10.6151
R545 B.n483 B.n482 10.6151
R546 B.n483 B.n4 10.6151
R547 B.n487 B.n4 10.6151
R548 B.n488 B.n487 10.6151
R549 B.n489 B.n488 10.6151
R550 B.n489 B.n0 10.6151
R551 B.n423 B.n422 10.6151
R552 B.n422 B.n421 10.6151
R553 B.n421 B.n26 10.6151
R554 B.n417 B.n26 10.6151
R555 B.n417 B.n416 10.6151
R556 B.n416 B.n415 10.6151
R557 B.n415 B.n28 10.6151
R558 B.n411 B.n28 10.6151
R559 B.n411 B.n410 10.6151
R560 B.n408 B.n32 10.6151
R561 B.n404 B.n32 10.6151
R562 B.n404 B.n403 10.6151
R563 B.n403 B.n402 10.6151
R564 B.n402 B.n34 10.6151
R565 B.n398 B.n34 10.6151
R566 B.n398 B.n397 10.6151
R567 B.n397 B.n396 10.6151
R568 B.n393 B.n392 10.6151
R569 B.n392 B.n391 10.6151
R570 B.n391 B.n40 10.6151
R571 B.n387 B.n40 10.6151
R572 B.n387 B.n386 10.6151
R573 B.n386 B.n385 10.6151
R574 B.n385 B.n42 10.6151
R575 B.n381 B.n42 10.6151
R576 B.n381 B.n380 10.6151
R577 B.n379 B.n44 10.6151
R578 B.n375 B.n44 10.6151
R579 B.n375 B.n374 10.6151
R580 B.n374 B.n373 10.6151
R581 B.n373 B.n46 10.6151
R582 B.n369 B.n46 10.6151
R583 B.n369 B.n368 10.6151
R584 B.n368 B.n367 10.6151
R585 B.n367 B.n48 10.6151
R586 B.n363 B.n48 10.6151
R587 B.n363 B.n362 10.6151
R588 B.n362 B.n361 10.6151
R589 B.n361 B.n50 10.6151
R590 B.n357 B.n50 10.6151
R591 B.n357 B.n356 10.6151
R592 B.n356 B.n355 10.6151
R593 B.n355 B.n52 10.6151
R594 B.n351 B.n52 10.6151
R595 B.n351 B.n350 10.6151
R596 B.n350 B.n349 10.6151
R597 B.n349 B.n54 10.6151
R598 B.n345 B.n54 10.6151
R599 B.n345 B.n344 10.6151
R600 B.n344 B.n343 10.6151
R601 B.n343 B.n56 10.6151
R602 B.n339 B.n56 10.6151
R603 B.n339 B.n338 10.6151
R604 B.n338 B.n337 10.6151
R605 B.n337 B.n58 10.6151
R606 B.n333 B.n58 10.6151
R607 B.n333 B.n332 10.6151
R608 B.n332 B.n331 10.6151
R609 B.n331 B.n60 10.6151
R610 B.n327 B.n60 10.6151
R611 B.n327 B.n326 10.6151
R612 B.n326 B.n325 10.6151
R613 B.n325 B.n62 10.6151
R614 B.n321 B.n62 10.6151
R615 B.n321 B.n320 10.6151
R616 B.n320 B.n319 10.6151
R617 B.n319 B.n64 10.6151
R618 B.n315 B.n64 10.6151
R619 B.n315 B.n314 10.6151
R620 B.n314 B.n313 10.6151
R621 B.n313 B.n66 10.6151
R622 B.n309 B.n66 10.6151
R623 B.n309 B.n308 10.6151
R624 B.n308 B.n307 10.6151
R625 B.n307 B.n68 10.6151
R626 B.n303 B.n68 10.6151
R627 B.n303 B.n302 10.6151
R628 B.n302 B.n301 10.6151
R629 B.n301 B.n70 10.6151
R630 B.n297 B.n70 10.6151
R631 B.n297 B.n296 10.6151
R632 B.n296 B.n295 10.6151
R633 B.n295 B.n72 10.6151
R634 B.n291 B.n72 10.6151
R635 B.n291 B.n290 10.6151
R636 B.n290 B.n289 10.6151
R637 B.n289 B.n74 10.6151
R638 B.n285 B.n74 10.6151
R639 B.n285 B.n284 10.6151
R640 B.n284 B.n283 10.6151
R641 B.n283 B.n76 10.6151
R642 B.n279 B.n76 10.6151
R643 B.n279 B.n278 10.6151
R644 B.n278 B.n277 10.6151
R645 B.n277 B.n78 10.6151
R646 B.n273 B.n78 10.6151
R647 B.n273 B.n272 10.6151
R648 B.n272 B.n271 10.6151
R649 B.n271 B.n80 10.6151
R650 B.n267 B.n80 10.6151
R651 B.n267 B.n266 10.6151
R652 B.n266 B.n265 10.6151
R653 B.n265 B.n82 10.6151
R654 B.n261 B.n82 10.6151
R655 B.n261 B.n260 10.6151
R656 B.n260 B.n259 10.6151
R657 B.n259 B.n84 10.6151
R658 B.n255 B.n84 10.6151
R659 B.n255 B.n254 10.6151
R660 B.n254 B.n253 10.6151
R661 B.n253 B.n86 10.6151
R662 B.n249 B.n86 10.6151
R663 B.n249 B.n248 10.6151
R664 B.n248 B.n247 10.6151
R665 B.n247 B.n88 10.6151
R666 B.n243 B.n88 10.6151
R667 B.n243 B.n242 10.6151
R668 B.n129 B.n1 10.6151
R669 B.n130 B.n129 10.6151
R670 B.n131 B.n130 10.6151
R671 B.n131 B.n126 10.6151
R672 B.n135 B.n126 10.6151
R673 B.n136 B.n135 10.6151
R674 B.n137 B.n136 10.6151
R675 B.n137 B.n124 10.6151
R676 B.n141 B.n124 10.6151
R677 B.n142 B.n141 10.6151
R678 B.n143 B.n142 10.6151
R679 B.n143 B.n122 10.6151
R680 B.n147 B.n122 10.6151
R681 B.n148 B.n147 10.6151
R682 B.n149 B.n148 10.6151
R683 B.n149 B.n120 10.6151
R684 B.n153 B.n120 10.6151
R685 B.n154 B.n153 10.6151
R686 B.n155 B.n154 10.6151
R687 B.n155 B.n118 10.6151
R688 B.n159 B.n118 10.6151
R689 B.n160 B.n159 10.6151
R690 B.n161 B.n160 10.6151
R691 B.n161 B.n116 10.6151
R692 B.n165 B.n116 10.6151
R693 B.n166 B.n165 10.6151
R694 B.n167 B.n166 10.6151
R695 B.n167 B.n114 10.6151
R696 B.n171 B.n114 10.6151
R697 B.n172 B.n171 10.6151
R698 B.n173 B.n172 10.6151
R699 B.n173 B.n112 10.6151
R700 B.n177 B.n112 10.6151
R701 B.n178 B.n177 10.6151
R702 B.n179 B.n178 10.6151
R703 B.n179 B.n110 10.6151
R704 B.n183 B.n110 10.6151
R705 B.n184 B.n183 10.6151
R706 B.n185 B.n184 10.6151
R707 B.n185 B.n108 10.6151
R708 B.n189 B.n108 10.6151
R709 B.n190 B.n189 10.6151
R710 B.n191 B.n190 10.6151
R711 B.n191 B.n106 10.6151
R712 B.n196 B.n195 10.6151
R713 B.n197 B.n196 10.6151
R714 B.n197 B.n104 10.6151
R715 B.n201 B.n104 10.6151
R716 B.n202 B.n201 10.6151
R717 B.n203 B.n202 10.6151
R718 B.n203 B.n102 10.6151
R719 B.n207 B.n102 10.6151
R720 B.n208 B.n207 10.6151
R721 B.n210 B.n98 10.6151
R722 B.n214 B.n98 10.6151
R723 B.n215 B.n214 10.6151
R724 B.n216 B.n215 10.6151
R725 B.n216 B.n96 10.6151
R726 B.n220 B.n96 10.6151
R727 B.n221 B.n220 10.6151
R728 B.n225 B.n221 10.6151
R729 B.n229 B.n94 10.6151
R730 B.n230 B.n229 10.6151
R731 B.n231 B.n230 10.6151
R732 B.n231 B.n92 10.6151
R733 B.n235 B.n92 10.6151
R734 B.n236 B.n235 10.6151
R735 B.n237 B.n236 10.6151
R736 B.n237 B.n90 10.6151
R737 B.n241 B.n90 10.6151
R738 B.n493 B.n0 8.11757
R739 B.n493 B.n1 8.11757
R740 B.n409 B.n408 6.5566
R741 B.n396 B.n38 6.5566
R742 B.n210 B.n209 6.5566
R743 B.n225 B.n224 6.5566
R744 B.n410 B.n409 4.05904
R745 B.n393 B.n38 4.05904
R746 B.n209 B.n208 4.05904
R747 B.n224 B.n94 4.05904
R748 VP.n13 VP.n10 161.3
R749 VP.n15 VP.n14 161.3
R750 VP.n16 VP.n9 161.3
R751 VP.n18 VP.n17 161.3
R752 VP.n19 VP.n8 161.3
R753 VP.n21 VP.n20 161.3
R754 VP.n43 VP.n42 161.3
R755 VP.n41 VP.n1 161.3
R756 VP.n40 VP.n39 161.3
R757 VP.n38 VP.n2 161.3
R758 VP.n37 VP.n36 161.3
R759 VP.n35 VP.n3 161.3
R760 VP.n33 VP.n32 161.3
R761 VP.n31 VP.n4 161.3
R762 VP.n30 VP.n29 161.3
R763 VP.n28 VP.n5 161.3
R764 VP.n27 VP.n26 161.3
R765 VP.n25 VP.n6 161.3
R766 VP.n24 VP.n23 68.1129
R767 VP.n44 VP.n0 68.1129
R768 VP.n22 VP.n7 68.1129
R769 VP.n12 VP.n11 61.6887
R770 VP.n29 VP.n28 55.1086
R771 VP.n40 VP.n2 55.1086
R772 VP.n18 VP.n9 55.1086
R773 VP.n24 VP.n22 41.6132
R774 VP.n11 VP.t0 41.2847
R775 VP.n28 VP.n27 26.0455
R776 VP.n41 VP.n40 26.0455
R777 VP.n19 VP.n18 26.0455
R778 VP.n27 VP.n6 24.5923
R779 VP.n29 VP.n4 24.5923
R780 VP.n33 VP.n4 24.5923
R781 VP.n36 VP.n35 24.5923
R782 VP.n36 VP.n2 24.5923
R783 VP.n42 VP.n41 24.5923
R784 VP.n20 VP.n19 24.5923
R785 VP.n14 VP.n13 24.5923
R786 VP.n14 VP.n9 24.5923
R787 VP.n23 VP.n6 22.1332
R788 VP.n42 VP.n0 22.1332
R789 VP.n20 VP.n7 22.1332
R790 VP.n34 VP.n33 12.2964
R791 VP.n35 VP.n34 12.2964
R792 VP.n13 VP.n12 12.2964
R793 VP.n23 VP.t5 9.40538
R794 VP.n34 VP.t4 9.40538
R795 VP.n0 VP.t2 9.40538
R796 VP.n7 VP.t3 9.40538
R797 VP.n12 VP.t1 9.40538
R798 VP.n11 VP.n10 5.38463
R799 VP.n22 VP.n21 0.354861
R800 VP.n25 VP.n24 0.354861
R801 VP.n44 VP.n43 0.354861
R802 VP VP.n44 0.267071
R803 VP.n15 VP.n10 0.189894
R804 VP.n16 VP.n15 0.189894
R805 VP.n17 VP.n16 0.189894
R806 VP.n17 VP.n8 0.189894
R807 VP.n21 VP.n8 0.189894
R808 VP.n26 VP.n25 0.189894
R809 VP.n26 VP.n5 0.189894
R810 VP.n30 VP.n5 0.189894
R811 VP.n31 VP.n30 0.189894
R812 VP.n32 VP.n31 0.189894
R813 VP.n32 VP.n3 0.189894
R814 VP.n37 VP.n3 0.189894
R815 VP.n38 VP.n37 0.189894
R816 VP.n39 VP.n38 0.189894
R817 VP.n39 VP.n1 0.189894
R818 VP.n43 VP.n1 0.189894
R819 VTAIL.n11 VTAIL.t1 372.911
R820 VTAIL.n2 VTAIL.t5 372.911
R821 VTAIL.n10 VTAIL.t10 372.911
R822 VTAIL.n7 VTAIL.t0 372.911
R823 VTAIL.n1 VTAIL.n0 329.974
R824 VTAIL.n4 VTAIL.n3 329.974
R825 VTAIL.n9 VTAIL.n8 329.973
R826 VTAIL.n6 VTAIL.n5 329.973
R827 VTAIL.n0 VTAIL.t3 29.0228
R828 VTAIL.n0 VTAIL.t2 29.0228
R829 VTAIL.n3 VTAIL.t6 29.0228
R830 VTAIL.n3 VTAIL.t8 29.0228
R831 VTAIL.n8 VTAIL.t7 29.0228
R832 VTAIL.n8 VTAIL.t9 29.0228
R833 VTAIL.n5 VTAIL.t11 29.0228
R834 VTAIL.n5 VTAIL.t4 29.0228
R835 VTAIL.n6 VTAIL.n4 18.8496
R836 VTAIL.n11 VTAIL.n10 16.091
R837 VTAIL.n7 VTAIL.n6 2.75912
R838 VTAIL.n10 VTAIL.n9 2.75912
R839 VTAIL.n4 VTAIL.n2 2.75912
R840 VTAIL VTAIL.n11 2.01128
R841 VTAIL.n9 VTAIL.n7 1.84964
R842 VTAIL.n2 VTAIL.n1 1.84964
R843 VTAIL VTAIL.n1 0.748345
R844 VDD1 VDD1.t5 391.716
R845 VDD1.n1 VDD1.t0 391.603
R846 VDD1.n1 VDD1.n0 347.286
R847 VDD1.n3 VDD1.n2 346.651
R848 VDD1.n3 VDD1.n1 35.6087
R849 VDD1.n2 VDD1.t4 29.0228
R850 VDD1.n2 VDD1.t2 29.0228
R851 VDD1.n0 VDD1.t1 29.0228
R852 VDD1.n0 VDD1.t3 29.0228
R853 VDD1 VDD1.n3 0.631965
R854 VN.n30 VN.n29 161.3
R855 VN.n28 VN.n17 161.3
R856 VN.n27 VN.n26 161.3
R857 VN.n25 VN.n18 161.3
R858 VN.n24 VN.n23 161.3
R859 VN.n22 VN.n19 161.3
R860 VN.n14 VN.n13 161.3
R861 VN.n12 VN.n1 161.3
R862 VN.n11 VN.n10 161.3
R863 VN.n9 VN.n2 161.3
R864 VN.n8 VN.n7 161.3
R865 VN.n6 VN.n3 161.3
R866 VN.n15 VN.n0 68.1129
R867 VN.n31 VN.n16 68.1129
R868 VN.n5 VN.n4 61.6886
R869 VN.n21 VN.n20 61.6886
R870 VN.n11 VN.n2 55.1086
R871 VN.n27 VN.n18 55.1086
R872 VN VN.n31 41.7784
R873 VN.n4 VN.t5 41.2849
R874 VN.n20 VN.t2 41.2849
R875 VN.n12 VN.n11 26.0455
R876 VN.n28 VN.n27 26.0455
R877 VN.n7 VN.n6 24.5923
R878 VN.n7 VN.n2 24.5923
R879 VN.n13 VN.n12 24.5923
R880 VN.n23 VN.n18 24.5923
R881 VN.n23 VN.n22 24.5923
R882 VN.n29 VN.n28 24.5923
R883 VN.n13 VN.n0 22.1332
R884 VN.n29 VN.n16 22.1332
R885 VN.n6 VN.n5 12.2964
R886 VN.n22 VN.n21 12.2964
R887 VN.n5 VN.t1 9.40538
R888 VN.n0 VN.t3 9.40538
R889 VN.n21 VN.t4 9.40538
R890 VN.n16 VN.t0 9.40538
R891 VN.n4 VN.n3 5.38467
R892 VN.n20 VN.n19 5.38467
R893 VN.n31 VN.n30 0.354861
R894 VN.n15 VN.n14 0.354861
R895 VN VN.n15 0.267071
R896 VN.n30 VN.n17 0.189894
R897 VN.n26 VN.n17 0.189894
R898 VN.n26 VN.n25 0.189894
R899 VN.n25 VN.n24 0.189894
R900 VN.n24 VN.n19 0.189894
R901 VN.n8 VN.n3 0.189894
R902 VN.n9 VN.n8 0.189894
R903 VN.n10 VN.n9 0.189894
R904 VN.n10 VN.n1 0.189894
R905 VN.n14 VN.n1 0.189894
R906 VDD2.n1 VDD2.t0 391.603
R907 VDD2.n2 VDD2.t5 389.589
R908 VDD2.n1 VDD2.n0 347.286
R909 VDD2 VDD2.n3 347.284
R910 VDD2.n2 VDD2.n1 33.6463
R911 VDD2.n3 VDD2.t1 29.0228
R912 VDD2.n3 VDD2.t3 29.0228
R913 VDD2.n0 VDD2.t4 29.0228
R914 VDD2.n0 VDD2.t2 29.0228
R915 VDD2 VDD2.n2 2.12766
C0 B VN 1.05897f
C1 VTAIL VN 2.06838f
C2 B VDD1 1.29781f
C3 VTAIL VDD1 3.98287f
C4 B w_n3530_n1192# 7.07453f
C5 w_n3530_n1192# VTAIL 1.41988f
C6 B VDD2 1.379f
C7 VDD2 VTAIL 4.03808f
C8 B VP 1.82238f
C9 VTAIL VP 2.0825f
C10 VN VDD1 0.159162f
C11 w_n3530_n1192# VN 6.55562f
C12 VDD2 VN 0.997558f
C13 w_n3530_n1192# VDD1 1.59606f
C14 VN VP 5.18077f
C15 VDD2 VDD1 1.51151f
C16 w_n3530_n1192# VDD2 1.68871f
C17 VP VDD1 1.32509f
C18 w_n3530_n1192# VP 7.00541f
C19 B VTAIL 1.15525f
C20 VDD2 VP 0.490111f
C21 VDD2 VSUBS 1.076125f
C22 VDD1 VSUBS 1.54596f
C23 VTAIL VSUBS 0.563283f
C24 VN VSUBS 6.33185f
C25 VP VSUBS 2.56535f
C26 B VSUBS 3.743083f
C27 w_n3530_n1192# VSUBS 54.1784f
C28 VDD2.t0 VSUBS 0.089974f
C29 VDD2.t4 VSUBS 0.016206f
C30 VDD2.t2 VSUBS 0.016206f
C31 VDD2.n0 VSUBS 0.054492f
C32 VDD2.n1 VSUBS 1.70426f
C33 VDD2.t5 VSUBS 0.088519f
C34 VDD2.n2 VSUBS 1.42696f
C35 VDD2.t1 VSUBS 0.016206f
C36 VDD2.t3 VSUBS 0.016206f
C37 VDD2.n3 VSUBS 0.054487f
C38 VN.t3 VSUBS 0.369537f
C39 VN.n0 VSUBS 0.457392f
C40 VN.n1 VSUBS 0.058404f
C41 VN.n2 VSUBS 0.100607f
C42 VN.n3 VSUBS 0.620567f
C43 VN.t1 VSUBS 0.369537f
C44 VN.t5 VSUBS 0.841674f
C45 VN.n4 VSUBS 0.426264f
C46 VN.n5 VSUBS 0.409085f
C47 VN.n6 VSUBS 0.081572f
C48 VN.n7 VSUBS 0.108305f
C49 VN.n8 VSUBS 0.058404f
C50 VN.n9 VSUBS 0.058404f
C51 VN.n10 VSUBS 0.058404f
C52 VN.n11 VSUBS 0.066388f
C53 VN.n12 VSUBS 0.111109f
C54 VN.n13 VSUBS 0.102959f
C55 VN.n14 VSUBS 0.094248f
C56 VN.n15 VSUBS 0.113654f
C57 VN.t0 VSUBS 0.369537f
C58 VN.n16 VSUBS 0.457392f
C59 VN.n17 VSUBS 0.058404f
C60 VN.n18 VSUBS 0.100607f
C61 VN.n19 VSUBS 0.620567f
C62 VN.t4 VSUBS 0.369537f
C63 VN.t2 VSUBS 0.841674f
C64 VN.n20 VSUBS 0.426264f
C65 VN.n21 VSUBS 0.409085f
C66 VN.n22 VSUBS 0.081572f
C67 VN.n23 VSUBS 0.108305f
C68 VN.n24 VSUBS 0.058404f
C69 VN.n25 VSUBS 0.058404f
C70 VN.n26 VSUBS 0.058404f
C71 VN.n27 VSUBS 0.066388f
C72 VN.n28 VSUBS 0.111109f
C73 VN.n29 VSUBS 0.102959f
C74 VN.n30 VSUBS 0.094248f
C75 VN.n31 VSUBS 2.51635f
C76 VDD1.t5 VSUBS 0.088593f
C77 VDD1.t0 VSUBS 0.088478f
C78 VDD1.t1 VSUBS 0.015937f
C79 VDD1.t3 VSUBS 0.015937f
C80 VDD1.n0 VSUBS 0.053585f
C81 VDD1.n1 VSUBS 1.76138f
C82 VDD1.t4 VSUBS 0.015937f
C83 VDD1.t2 VSUBS 0.015937f
C84 VDD1.n2 VSUBS 0.052948f
C85 VDD1.n3 VSUBS 1.4482f
C86 VTAIL.t3 VSUBS 0.034984f
C87 VTAIL.t2 VSUBS 0.034984f
C88 VTAIL.n0 VSUBS 0.100572f
C89 VTAIL.n1 VSUBS 0.609925f
C90 VTAIL.t5 VSUBS 0.176309f
C91 VTAIL.n2 VSUBS 0.885703f
C92 VTAIL.t6 VSUBS 0.034984f
C93 VTAIL.t8 VSUBS 0.034984f
C94 VTAIL.n3 VSUBS 0.100572f
C95 VTAIL.n4 VSUBS 1.99312f
C96 VTAIL.t11 VSUBS 0.034984f
C97 VTAIL.t4 VSUBS 0.034984f
C98 VTAIL.n5 VSUBS 0.100572f
C99 VTAIL.n6 VSUBS 1.99312f
C100 VTAIL.t0 VSUBS 0.176309f
C101 VTAIL.n7 VSUBS 0.885703f
C102 VTAIL.t7 VSUBS 0.034984f
C103 VTAIL.t9 VSUBS 0.034984f
C104 VTAIL.n8 VSUBS 0.100572f
C105 VTAIL.n9 VSUBS 0.866029f
C106 VTAIL.t10 VSUBS 0.176309f
C107 VTAIL.n10 VSUBS 1.66144f
C108 VTAIL.t1 VSUBS 0.176309f
C109 VTAIL.n11 VSUBS 1.5662f
C110 VP.t2 VSUBS 0.38243f
C111 VP.n0 VSUBS 0.473351f
C112 VP.n1 VSUBS 0.060442f
C113 VP.n2 VSUBS 0.104117f
C114 VP.n3 VSUBS 0.060442f
C115 VP.t4 VSUBS 0.38243f
C116 VP.n4 VSUBS 0.112084f
C117 VP.n5 VSUBS 0.060442f
C118 VP.n6 VSUBS 0.106551f
C119 VP.t3 VSUBS 0.38243f
C120 VP.n7 VSUBS 0.473351f
C121 VP.n8 VSUBS 0.060442f
C122 VP.n9 VSUBS 0.104117f
C123 VP.n10 VSUBS 0.642219f
C124 VP.t1 VSUBS 0.38243f
C125 VP.t0 VSUBS 0.871038f
C126 VP.n11 VSUBS 0.441137f
C127 VP.n12 VSUBS 0.423358f
C128 VP.n13 VSUBS 0.084417f
C129 VP.n14 VSUBS 0.112084f
C130 VP.n15 VSUBS 0.060442f
C131 VP.n16 VSUBS 0.060442f
C132 VP.n17 VSUBS 0.060442f
C133 VP.n18 VSUBS 0.068704f
C134 VP.n19 VSUBS 0.114986f
C135 VP.n20 VSUBS 0.106551f
C136 VP.n21 VSUBS 0.097537f
C137 VP.n22 VSUBS 2.57769f
C138 VP.t5 VSUBS 0.38243f
C139 VP.n23 VSUBS 0.473351f
C140 VP.n24 VSUBS 2.63005f
C141 VP.n25 VSUBS 0.097537f
C142 VP.n26 VSUBS 0.060442f
C143 VP.n27 VSUBS 0.114986f
C144 VP.n28 VSUBS 0.068704f
C145 VP.n29 VSUBS 0.104117f
C146 VP.n30 VSUBS 0.060442f
C147 VP.n31 VSUBS 0.060442f
C148 VP.n32 VSUBS 0.060442f
C149 VP.n33 VSUBS 0.084417f
C150 VP.n34 VSUBS 0.236825f
C151 VP.n35 VSUBS 0.084417f
C152 VP.n36 VSUBS 0.112084f
C153 VP.n37 VSUBS 0.060442f
C154 VP.n38 VSUBS 0.060442f
C155 VP.n39 VSUBS 0.060442f
C156 VP.n40 VSUBS 0.068704f
C157 VP.n41 VSUBS 0.114986f
C158 VP.n42 VSUBS 0.106551f
C159 VP.n43 VSUBS 0.097537f
C160 VP.n44 VSUBS 0.117619f
C161 B.n0 VSUBS 0.008935f
C162 B.n1 VSUBS 0.008935f
C163 B.n2 VSUBS 0.013214f
C164 B.n3 VSUBS 0.010126f
C165 B.n4 VSUBS 0.010126f
C166 B.n5 VSUBS 0.010126f
C167 B.n6 VSUBS 0.010126f
C168 B.n7 VSUBS 0.010126f
C169 B.n8 VSUBS 0.010126f
C170 B.n9 VSUBS 0.010126f
C171 B.n10 VSUBS 0.010126f
C172 B.n11 VSUBS 0.010126f
C173 B.n12 VSUBS 0.010126f
C174 B.n13 VSUBS 0.010126f
C175 B.n14 VSUBS 0.010126f
C176 B.n15 VSUBS 0.010126f
C177 B.n16 VSUBS 0.010126f
C178 B.n17 VSUBS 0.010126f
C179 B.n18 VSUBS 0.010126f
C180 B.n19 VSUBS 0.010126f
C181 B.n20 VSUBS 0.010126f
C182 B.n21 VSUBS 0.010126f
C183 B.n22 VSUBS 0.010126f
C184 B.n23 VSUBS 0.010126f
C185 B.n24 VSUBS 0.023544f
C186 B.n25 VSUBS 0.010126f
C187 B.n26 VSUBS 0.010126f
C188 B.n27 VSUBS 0.010126f
C189 B.n28 VSUBS 0.010126f
C190 B.n29 VSUBS 0.010126f
C191 B.t4 VSUBS 0.030511f
C192 B.t5 VSUBS 0.038851f
C193 B.t3 VSUBS 0.235054f
C194 B.n30 VSUBS 0.093562f
C195 B.n31 VSUBS 0.071635f
C196 B.n32 VSUBS 0.010126f
C197 B.n33 VSUBS 0.010126f
C198 B.n34 VSUBS 0.010126f
C199 B.n35 VSUBS 0.010126f
C200 B.t1 VSUBS 0.030511f
C201 B.t2 VSUBS 0.038851f
C202 B.t0 VSUBS 0.235054f
C203 B.n36 VSUBS 0.093562f
C204 B.n37 VSUBS 0.071635f
C205 B.n38 VSUBS 0.023461f
C206 B.n39 VSUBS 0.010126f
C207 B.n40 VSUBS 0.010126f
C208 B.n41 VSUBS 0.010126f
C209 B.n42 VSUBS 0.010126f
C210 B.n43 VSUBS 0.0253f
C211 B.n44 VSUBS 0.010126f
C212 B.n45 VSUBS 0.010126f
C213 B.n46 VSUBS 0.010126f
C214 B.n47 VSUBS 0.010126f
C215 B.n48 VSUBS 0.010126f
C216 B.n49 VSUBS 0.010126f
C217 B.n50 VSUBS 0.010126f
C218 B.n51 VSUBS 0.010126f
C219 B.n52 VSUBS 0.010126f
C220 B.n53 VSUBS 0.010126f
C221 B.n54 VSUBS 0.010126f
C222 B.n55 VSUBS 0.010126f
C223 B.n56 VSUBS 0.010126f
C224 B.n57 VSUBS 0.010126f
C225 B.n58 VSUBS 0.010126f
C226 B.n59 VSUBS 0.010126f
C227 B.n60 VSUBS 0.010126f
C228 B.n61 VSUBS 0.010126f
C229 B.n62 VSUBS 0.010126f
C230 B.n63 VSUBS 0.010126f
C231 B.n64 VSUBS 0.010126f
C232 B.n65 VSUBS 0.010126f
C233 B.n66 VSUBS 0.010126f
C234 B.n67 VSUBS 0.010126f
C235 B.n68 VSUBS 0.010126f
C236 B.n69 VSUBS 0.010126f
C237 B.n70 VSUBS 0.010126f
C238 B.n71 VSUBS 0.010126f
C239 B.n72 VSUBS 0.010126f
C240 B.n73 VSUBS 0.010126f
C241 B.n74 VSUBS 0.010126f
C242 B.n75 VSUBS 0.010126f
C243 B.n76 VSUBS 0.010126f
C244 B.n77 VSUBS 0.010126f
C245 B.n78 VSUBS 0.010126f
C246 B.n79 VSUBS 0.010126f
C247 B.n80 VSUBS 0.010126f
C248 B.n81 VSUBS 0.010126f
C249 B.n82 VSUBS 0.010126f
C250 B.n83 VSUBS 0.010126f
C251 B.n84 VSUBS 0.010126f
C252 B.n85 VSUBS 0.010126f
C253 B.n86 VSUBS 0.010126f
C254 B.n87 VSUBS 0.010126f
C255 B.n88 VSUBS 0.010126f
C256 B.n89 VSUBS 0.023544f
C257 B.n90 VSUBS 0.010126f
C258 B.n91 VSUBS 0.010126f
C259 B.n92 VSUBS 0.010126f
C260 B.n93 VSUBS 0.010126f
C261 B.n94 VSUBS 0.006999f
C262 B.n95 VSUBS 0.010126f
C263 B.n96 VSUBS 0.010126f
C264 B.n97 VSUBS 0.010126f
C265 B.n98 VSUBS 0.010126f
C266 B.n99 VSUBS 0.010126f
C267 B.t11 VSUBS 0.030511f
C268 B.t10 VSUBS 0.038851f
C269 B.t9 VSUBS 0.235054f
C270 B.n100 VSUBS 0.093562f
C271 B.n101 VSUBS 0.071635f
C272 B.n102 VSUBS 0.010126f
C273 B.n103 VSUBS 0.010126f
C274 B.n104 VSUBS 0.010126f
C275 B.n105 VSUBS 0.010126f
C276 B.n106 VSUBS 0.023544f
C277 B.n107 VSUBS 0.010126f
C278 B.n108 VSUBS 0.010126f
C279 B.n109 VSUBS 0.010126f
C280 B.n110 VSUBS 0.010126f
C281 B.n111 VSUBS 0.010126f
C282 B.n112 VSUBS 0.010126f
C283 B.n113 VSUBS 0.010126f
C284 B.n114 VSUBS 0.010126f
C285 B.n115 VSUBS 0.010126f
C286 B.n116 VSUBS 0.010126f
C287 B.n117 VSUBS 0.010126f
C288 B.n118 VSUBS 0.010126f
C289 B.n119 VSUBS 0.010126f
C290 B.n120 VSUBS 0.010126f
C291 B.n121 VSUBS 0.010126f
C292 B.n122 VSUBS 0.010126f
C293 B.n123 VSUBS 0.010126f
C294 B.n124 VSUBS 0.010126f
C295 B.n125 VSUBS 0.010126f
C296 B.n126 VSUBS 0.010126f
C297 B.n127 VSUBS 0.010126f
C298 B.n128 VSUBS 0.010126f
C299 B.n129 VSUBS 0.010126f
C300 B.n130 VSUBS 0.010126f
C301 B.n131 VSUBS 0.010126f
C302 B.n132 VSUBS 0.010126f
C303 B.n133 VSUBS 0.010126f
C304 B.n134 VSUBS 0.010126f
C305 B.n135 VSUBS 0.010126f
C306 B.n136 VSUBS 0.010126f
C307 B.n137 VSUBS 0.010126f
C308 B.n138 VSUBS 0.010126f
C309 B.n139 VSUBS 0.010126f
C310 B.n140 VSUBS 0.010126f
C311 B.n141 VSUBS 0.010126f
C312 B.n142 VSUBS 0.010126f
C313 B.n143 VSUBS 0.010126f
C314 B.n144 VSUBS 0.010126f
C315 B.n145 VSUBS 0.010126f
C316 B.n146 VSUBS 0.010126f
C317 B.n147 VSUBS 0.010126f
C318 B.n148 VSUBS 0.010126f
C319 B.n149 VSUBS 0.010126f
C320 B.n150 VSUBS 0.010126f
C321 B.n151 VSUBS 0.010126f
C322 B.n152 VSUBS 0.010126f
C323 B.n153 VSUBS 0.010126f
C324 B.n154 VSUBS 0.010126f
C325 B.n155 VSUBS 0.010126f
C326 B.n156 VSUBS 0.010126f
C327 B.n157 VSUBS 0.010126f
C328 B.n158 VSUBS 0.010126f
C329 B.n159 VSUBS 0.010126f
C330 B.n160 VSUBS 0.010126f
C331 B.n161 VSUBS 0.010126f
C332 B.n162 VSUBS 0.010126f
C333 B.n163 VSUBS 0.010126f
C334 B.n164 VSUBS 0.010126f
C335 B.n165 VSUBS 0.010126f
C336 B.n166 VSUBS 0.010126f
C337 B.n167 VSUBS 0.010126f
C338 B.n168 VSUBS 0.010126f
C339 B.n169 VSUBS 0.010126f
C340 B.n170 VSUBS 0.010126f
C341 B.n171 VSUBS 0.010126f
C342 B.n172 VSUBS 0.010126f
C343 B.n173 VSUBS 0.010126f
C344 B.n174 VSUBS 0.010126f
C345 B.n175 VSUBS 0.010126f
C346 B.n176 VSUBS 0.010126f
C347 B.n177 VSUBS 0.010126f
C348 B.n178 VSUBS 0.010126f
C349 B.n179 VSUBS 0.010126f
C350 B.n180 VSUBS 0.010126f
C351 B.n181 VSUBS 0.010126f
C352 B.n182 VSUBS 0.010126f
C353 B.n183 VSUBS 0.010126f
C354 B.n184 VSUBS 0.010126f
C355 B.n185 VSUBS 0.010126f
C356 B.n186 VSUBS 0.010126f
C357 B.n187 VSUBS 0.010126f
C358 B.n188 VSUBS 0.010126f
C359 B.n189 VSUBS 0.010126f
C360 B.n190 VSUBS 0.010126f
C361 B.n191 VSUBS 0.010126f
C362 B.n192 VSUBS 0.010126f
C363 B.n193 VSUBS 0.023544f
C364 B.n194 VSUBS 0.0253f
C365 B.n195 VSUBS 0.0253f
C366 B.n196 VSUBS 0.010126f
C367 B.n197 VSUBS 0.010126f
C368 B.n198 VSUBS 0.010126f
C369 B.n199 VSUBS 0.010126f
C370 B.n200 VSUBS 0.010126f
C371 B.n201 VSUBS 0.010126f
C372 B.n202 VSUBS 0.010126f
C373 B.n203 VSUBS 0.010126f
C374 B.n204 VSUBS 0.010126f
C375 B.n205 VSUBS 0.010126f
C376 B.n206 VSUBS 0.010126f
C377 B.n207 VSUBS 0.010126f
C378 B.n208 VSUBS 0.006999f
C379 B.n209 VSUBS 0.023461f
C380 B.n210 VSUBS 0.00819f
C381 B.n211 VSUBS 0.010126f
C382 B.n212 VSUBS 0.010126f
C383 B.n213 VSUBS 0.010126f
C384 B.n214 VSUBS 0.010126f
C385 B.n215 VSUBS 0.010126f
C386 B.n216 VSUBS 0.010126f
C387 B.n217 VSUBS 0.010126f
C388 B.n218 VSUBS 0.010126f
C389 B.n219 VSUBS 0.010126f
C390 B.n220 VSUBS 0.010126f
C391 B.n221 VSUBS 0.010126f
C392 B.t8 VSUBS 0.030511f
C393 B.t7 VSUBS 0.038851f
C394 B.t6 VSUBS 0.235054f
C395 B.n222 VSUBS 0.093562f
C396 B.n223 VSUBS 0.071635f
C397 B.n224 VSUBS 0.023461f
C398 B.n225 VSUBS 0.00819f
C399 B.n226 VSUBS 0.010126f
C400 B.n227 VSUBS 0.010126f
C401 B.n228 VSUBS 0.010126f
C402 B.n229 VSUBS 0.010126f
C403 B.n230 VSUBS 0.010126f
C404 B.n231 VSUBS 0.010126f
C405 B.n232 VSUBS 0.010126f
C406 B.n233 VSUBS 0.010126f
C407 B.n234 VSUBS 0.010126f
C408 B.n235 VSUBS 0.010126f
C409 B.n236 VSUBS 0.010126f
C410 B.n237 VSUBS 0.010126f
C411 B.n238 VSUBS 0.010126f
C412 B.n239 VSUBS 0.010126f
C413 B.n240 VSUBS 0.0253f
C414 B.n241 VSUBS 0.024157f
C415 B.n242 VSUBS 0.024687f
C416 B.n243 VSUBS 0.010126f
C417 B.n244 VSUBS 0.010126f
C418 B.n245 VSUBS 0.010126f
C419 B.n246 VSUBS 0.010126f
C420 B.n247 VSUBS 0.010126f
C421 B.n248 VSUBS 0.010126f
C422 B.n249 VSUBS 0.010126f
C423 B.n250 VSUBS 0.010126f
C424 B.n251 VSUBS 0.010126f
C425 B.n252 VSUBS 0.010126f
C426 B.n253 VSUBS 0.010126f
C427 B.n254 VSUBS 0.010126f
C428 B.n255 VSUBS 0.010126f
C429 B.n256 VSUBS 0.010126f
C430 B.n257 VSUBS 0.010126f
C431 B.n258 VSUBS 0.010126f
C432 B.n259 VSUBS 0.010126f
C433 B.n260 VSUBS 0.010126f
C434 B.n261 VSUBS 0.010126f
C435 B.n262 VSUBS 0.010126f
C436 B.n263 VSUBS 0.010126f
C437 B.n264 VSUBS 0.010126f
C438 B.n265 VSUBS 0.010126f
C439 B.n266 VSUBS 0.010126f
C440 B.n267 VSUBS 0.010126f
C441 B.n268 VSUBS 0.010126f
C442 B.n269 VSUBS 0.010126f
C443 B.n270 VSUBS 0.010126f
C444 B.n271 VSUBS 0.010126f
C445 B.n272 VSUBS 0.010126f
C446 B.n273 VSUBS 0.010126f
C447 B.n274 VSUBS 0.010126f
C448 B.n275 VSUBS 0.010126f
C449 B.n276 VSUBS 0.010126f
C450 B.n277 VSUBS 0.010126f
C451 B.n278 VSUBS 0.010126f
C452 B.n279 VSUBS 0.010126f
C453 B.n280 VSUBS 0.010126f
C454 B.n281 VSUBS 0.010126f
C455 B.n282 VSUBS 0.010126f
C456 B.n283 VSUBS 0.010126f
C457 B.n284 VSUBS 0.010126f
C458 B.n285 VSUBS 0.010126f
C459 B.n286 VSUBS 0.010126f
C460 B.n287 VSUBS 0.010126f
C461 B.n288 VSUBS 0.010126f
C462 B.n289 VSUBS 0.010126f
C463 B.n290 VSUBS 0.010126f
C464 B.n291 VSUBS 0.010126f
C465 B.n292 VSUBS 0.010126f
C466 B.n293 VSUBS 0.010126f
C467 B.n294 VSUBS 0.010126f
C468 B.n295 VSUBS 0.010126f
C469 B.n296 VSUBS 0.010126f
C470 B.n297 VSUBS 0.010126f
C471 B.n298 VSUBS 0.010126f
C472 B.n299 VSUBS 0.010126f
C473 B.n300 VSUBS 0.010126f
C474 B.n301 VSUBS 0.010126f
C475 B.n302 VSUBS 0.010126f
C476 B.n303 VSUBS 0.010126f
C477 B.n304 VSUBS 0.010126f
C478 B.n305 VSUBS 0.010126f
C479 B.n306 VSUBS 0.010126f
C480 B.n307 VSUBS 0.010126f
C481 B.n308 VSUBS 0.010126f
C482 B.n309 VSUBS 0.010126f
C483 B.n310 VSUBS 0.010126f
C484 B.n311 VSUBS 0.010126f
C485 B.n312 VSUBS 0.010126f
C486 B.n313 VSUBS 0.010126f
C487 B.n314 VSUBS 0.010126f
C488 B.n315 VSUBS 0.010126f
C489 B.n316 VSUBS 0.010126f
C490 B.n317 VSUBS 0.010126f
C491 B.n318 VSUBS 0.010126f
C492 B.n319 VSUBS 0.010126f
C493 B.n320 VSUBS 0.010126f
C494 B.n321 VSUBS 0.010126f
C495 B.n322 VSUBS 0.010126f
C496 B.n323 VSUBS 0.010126f
C497 B.n324 VSUBS 0.010126f
C498 B.n325 VSUBS 0.010126f
C499 B.n326 VSUBS 0.010126f
C500 B.n327 VSUBS 0.010126f
C501 B.n328 VSUBS 0.010126f
C502 B.n329 VSUBS 0.010126f
C503 B.n330 VSUBS 0.010126f
C504 B.n331 VSUBS 0.010126f
C505 B.n332 VSUBS 0.010126f
C506 B.n333 VSUBS 0.010126f
C507 B.n334 VSUBS 0.010126f
C508 B.n335 VSUBS 0.010126f
C509 B.n336 VSUBS 0.010126f
C510 B.n337 VSUBS 0.010126f
C511 B.n338 VSUBS 0.010126f
C512 B.n339 VSUBS 0.010126f
C513 B.n340 VSUBS 0.010126f
C514 B.n341 VSUBS 0.010126f
C515 B.n342 VSUBS 0.010126f
C516 B.n343 VSUBS 0.010126f
C517 B.n344 VSUBS 0.010126f
C518 B.n345 VSUBS 0.010126f
C519 B.n346 VSUBS 0.010126f
C520 B.n347 VSUBS 0.010126f
C521 B.n348 VSUBS 0.010126f
C522 B.n349 VSUBS 0.010126f
C523 B.n350 VSUBS 0.010126f
C524 B.n351 VSUBS 0.010126f
C525 B.n352 VSUBS 0.010126f
C526 B.n353 VSUBS 0.010126f
C527 B.n354 VSUBS 0.010126f
C528 B.n355 VSUBS 0.010126f
C529 B.n356 VSUBS 0.010126f
C530 B.n357 VSUBS 0.010126f
C531 B.n358 VSUBS 0.010126f
C532 B.n359 VSUBS 0.010126f
C533 B.n360 VSUBS 0.010126f
C534 B.n361 VSUBS 0.010126f
C535 B.n362 VSUBS 0.010126f
C536 B.n363 VSUBS 0.010126f
C537 B.n364 VSUBS 0.010126f
C538 B.n365 VSUBS 0.010126f
C539 B.n366 VSUBS 0.010126f
C540 B.n367 VSUBS 0.010126f
C541 B.n368 VSUBS 0.010126f
C542 B.n369 VSUBS 0.010126f
C543 B.n370 VSUBS 0.010126f
C544 B.n371 VSUBS 0.010126f
C545 B.n372 VSUBS 0.010126f
C546 B.n373 VSUBS 0.010126f
C547 B.n374 VSUBS 0.010126f
C548 B.n375 VSUBS 0.010126f
C549 B.n376 VSUBS 0.010126f
C550 B.n377 VSUBS 0.010126f
C551 B.n378 VSUBS 0.023544f
C552 B.n379 VSUBS 0.023544f
C553 B.n380 VSUBS 0.0253f
C554 B.n381 VSUBS 0.010126f
C555 B.n382 VSUBS 0.010126f
C556 B.n383 VSUBS 0.010126f
C557 B.n384 VSUBS 0.010126f
C558 B.n385 VSUBS 0.010126f
C559 B.n386 VSUBS 0.010126f
C560 B.n387 VSUBS 0.010126f
C561 B.n388 VSUBS 0.010126f
C562 B.n389 VSUBS 0.010126f
C563 B.n390 VSUBS 0.010126f
C564 B.n391 VSUBS 0.010126f
C565 B.n392 VSUBS 0.010126f
C566 B.n393 VSUBS 0.006999f
C567 B.n394 VSUBS 0.010126f
C568 B.n395 VSUBS 0.010126f
C569 B.n396 VSUBS 0.00819f
C570 B.n397 VSUBS 0.010126f
C571 B.n398 VSUBS 0.010126f
C572 B.n399 VSUBS 0.010126f
C573 B.n400 VSUBS 0.010126f
C574 B.n401 VSUBS 0.010126f
C575 B.n402 VSUBS 0.010126f
C576 B.n403 VSUBS 0.010126f
C577 B.n404 VSUBS 0.010126f
C578 B.n405 VSUBS 0.010126f
C579 B.n406 VSUBS 0.010126f
C580 B.n407 VSUBS 0.010126f
C581 B.n408 VSUBS 0.00819f
C582 B.n409 VSUBS 0.023461f
C583 B.n410 VSUBS 0.006999f
C584 B.n411 VSUBS 0.010126f
C585 B.n412 VSUBS 0.010126f
C586 B.n413 VSUBS 0.010126f
C587 B.n414 VSUBS 0.010126f
C588 B.n415 VSUBS 0.010126f
C589 B.n416 VSUBS 0.010126f
C590 B.n417 VSUBS 0.010126f
C591 B.n418 VSUBS 0.010126f
C592 B.n419 VSUBS 0.010126f
C593 B.n420 VSUBS 0.010126f
C594 B.n421 VSUBS 0.010126f
C595 B.n422 VSUBS 0.010126f
C596 B.n423 VSUBS 0.0253f
C597 B.n424 VSUBS 0.0253f
C598 B.n425 VSUBS 0.023544f
C599 B.n426 VSUBS 0.010126f
C600 B.n427 VSUBS 0.010126f
C601 B.n428 VSUBS 0.010126f
C602 B.n429 VSUBS 0.010126f
C603 B.n430 VSUBS 0.010126f
C604 B.n431 VSUBS 0.010126f
C605 B.n432 VSUBS 0.010126f
C606 B.n433 VSUBS 0.010126f
C607 B.n434 VSUBS 0.010126f
C608 B.n435 VSUBS 0.010126f
C609 B.n436 VSUBS 0.010126f
C610 B.n437 VSUBS 0.010126f
C611 B.n438 VSUBS 0.010126f
C612 B.n439 VSUBS 0.010126f
C613 B.n440 VSUBS 0.010126f
C614 B.n441 VSUBS 0.010126f
C615 B.n442 VSUBS 0.010126f
C616 B.n443 VSUBS 0.010126f
C617 B.n444 VSUBS 0.010126f
C618 B.n445 VSUBS 0.010126f
C619 B.n446 VSUBS 0.010126f
C620 B.n447 VSUBS 0.010126f
C621 B.n448 VSUBS 0.010126f
C622 B.n449 VSUBS 0.010126f
C623 B.n450 VSUBS 0.010126f
C624 B.n451 VSUBS 0.010126f
C625 B.n452 VSUBS 0.010126f
C626 B.n453 VSUBS 0.010126f
C627 B.n454 VSUBS 0.010126f
C628 B.n455 VSUBS 0.010126f
C629 B.n456 VSUBS 0.010126f
C630 B.n457 VSUBS 0.010126f
C631 B.n458 VSUBS 0.010126f
C632 B.n459 VSUBS 0.010126f
C633 B.n460 VSUBS 0.010126f
C634 B.n461 VSUBS 0.010126f
C635 B.n462 VSUBS 0.010126f
C636 B.n463 VSUBS 0.010126f
C637 B.n464 VSUBS 0.010126f
C638 B.n465 VSUBS 0.010126f
C639 B.n466 VSUBS 0.010126f
C640 B.n467 VSUBS 0.010126f
C641 B.n468 VSUBS 0.010126f
C642 B.n469 VSUBS 0.010126f
C643 B.n470 VSUBS 0.010126f
C644 B.n471 VSUBS 0.010126f
C645 B.n472 VSUBS 0.010126f
C646 B.n473 VSUBS 0.010126f
C647 B.n474 VSUBS 0.010126f
C648 B.n475 VSUBS 0.010126f
C649 B.n476 VSUBS 0.010126f
C650 B.n477 VSUBS 0.010126f
C651 B.n478 VSUBS 0.010126f
C652 B.n479 VSUBS 0.010126f
C653 B.n480 VSUBS 0.010126f
C654 B.n481 VSUBS 0.010126f
C655 B.n482 VSUBS 0.010126f
C656 B.n483 VSUBS 0.010126f
C657 B.n484 VSUBS 0.010126f
C658 B.n485 VSUBS 0.010126f
C659 B.n486 VSUBS 0.010126f
C660 B.n487 VSUBS 0.010126f
C661 B.n488 VSUBS 0.010126f
C662 B.n489 VSUBS 0.010126f
C663 B.n490 VSUBS 0.010126f
C664 B.n491 VSUBS 0.013214f
C665 B.n492 VSUBS 0.014076f
C666 B.n493 VSUBS 0.027992f
.ends

