* NGSPICE file created from diff_pair_sample_0220.ext - technology: sky130A

.subckt diff_pair_sample_0220 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=1.4079 ps=8 w=3.61 l=1.84
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0.59565 ps=3.94 w=3.61 l=1.84
X2 VTAIL.t0 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=0.59565 ps=3.94 w=3.61 l=1.84
X3 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0 ps=0 w=3.61 l=1.84
X4 VDD2.t4 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0.59565 ps=3.94 w=3.61 l=1.84
X5 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0.59565 ps=3.94 w=3.61 l=1.84
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0 ps=0 w=3.61 l=1.84
X7 VTAIL.t11 VP.t2 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=0.59565 ps=3.94 w=3.61 l=1.84
X8 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=1.4079 ps=8 w=3.61 l=1.84
X9 VTAIL.t7 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=0.59565 ps=3.94 w=3.61 l=1.84
X10 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=1.4079 ps=8 w=3.61 l=1.84
X11 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0 ps=0 w=3.61 l=1.84
X12 VDD1.t1 VP.t4 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0.59565 ps=3.94 w=3.61 l=1.84
X13 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=0.59565 ps=3.94 w=3.61 l=1.84
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4079 pd=8 as=0 ps=0 w=3.61 l=1.84
X15 VDD1.t0 VP.t5 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.59565 pd=3.94 as=1.4079 ps=8 w=3.61 l=1.84
R0 VP.n9 VP.n8 161.3
R1 VP.n10 VP.n5 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n13 VP.n4 161.3
R4 VP.n30 VP.n0 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n27 VP.n1 161.3
R7 VP.n26 VP.n25 161.3
R8 VP.n23 VP.n2 161.3
R9 VP.n22 VP.n21 161.3
R10 VP.n20 VP.n3 161.3
R11 VP.n19 VP.n18 161.3
R12 VP.n17 VP.n16 90.2042
R13 VP.n32 VP.n31 90.2042
R14 VP.n15 VP.n14 90.2042
R15 VP.n6 VP.t4 77.7446
R16 VP.n7 VP.n6 57.6509
R17 VP.n22 VP.n3 56.5193
R18 VP.n29 VP.n1 56.5193
R19 VP.n12 VP.n5 56.5193
R20 VP.n17 VP.t1 47.2837
R21 VP.n24 VP.t3 47.2837
R22 VP.n31 VP.t5 47.2837
R23 VP.n14 VP.t0 47.2837
R24 VP.n7 VP.t2 47.2837
R25 VP.n16 VP.n15 39.3367
R26 VP.n18 VP.n3 24.4675
R27 VP.n23 VP.n22 24.4675
R28 VP.n25 VP.n1 24.4675
R29 VP.n30 VP.n29 24.4675
R30 VP.n13 VP.n12 24.4675
R31 VP.n8 VP.n5 24.4675
R32 VP.n18 VP.n17 20.5528
R33 VP.n31 VP.n30 20.5528
R34 VP.n14 VP.n13 20.5528
R35 VP.n9 VP.n6 13.2264
R36 VP.n24 VP.n23 12.234
R37 VP.n25 VP.n24 12.234
R38 VP.n8 VP.n7 12.234
R39 VP.n15 VP.n4 0.278367
R40 VP.n19 VP.n16 0.278367
R41 VP.n32 VP.n0 0.278367
R42 VP.n10 VP.n9 0.189894
R43 VP.n11 VP.n10 0.189894
R44 VP.n11 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n21 VP.n20 0.189894
R47 VP.n21 VP.n2 0.189894
R48 VP.n26 VP.n2 0.189894
R49 VP.n27 VP.n26 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n28 VP.n0 0.189894
R52 VP VP.n32 0.153454
R53 VTAIL.n7 VTAIL.t5 66.6877
R54 VTAIL.n11 VTAIL.t4 66.6877
R55 VTAIL.n2 VTAIL.t8 66.6877
R56 VTAIL.n10 VTAIL.t9 66.6877
R57 VTAIL.n9 VTAIL.n8 61.2031
R58 VTAIL.n6 VTAIL.n5 61.2031
R59 VTAIL.n1 VTAIL.n0 61.2028
R60 VTAIL.n4 VTAIL.n3 61.2028
R61 VTAIL.n6 VTAIL.n4 19.2203
R62 VTAIL.n11 VTAIL.n10 17.3496
R63 VTAIL.n0 VTAIL.t1 5.48526
R64 VTAIL.n0 VTAIL.t2 5.48526
R65 VTAIL.n3 VTAIL.t10 5.48526
R66 VTAIL.n3 VTAIL.t7 5.48526
R67 VTAIL.n8 VTAIL.t6 5.48526
R68 VTAIL.n8 VTAIL.t11 5.48526
R69 VTAIL.n5 VTAIL.t3 5.48526
R70 VTAIL.n5 VTAIL.t0 5.48526
R71 VTAIL.n7 VTAIL.n6 1.87119
R72 VTAIL.n10 VTAIL.n9 1.87119
R73 VTAIL.n4 VTAIL.n2 1.87119
R74 VTAIL.n9 VTAIL.n7 1.40567
R75 VTAIL.n2 VTAIL.n1 1.40567
R76 VTAIL VTAIL.n11 1.34533
R77 VTAIL VTAIL.n1 0.526362
R78 VDD1 VDD1.t1 84.8277
R79 VDD1.n1 VDD1.t4 84.7142
R80 VDD1.n1 VDD1.n0 78.2939
R81 VDD1.n3 VDD1.n2 77.8817
R82 VDD1.n3 VDD1.n1 34.4255
R83 VDD1.n2 VDD1.t3 5.48526
R84 VDD1.n2 VDD1.t5 5.48526
R85 VDD1.n0 VDD1.t2 5.48526
R86 VDD1.n0 VDD1.t0 5.48526
R87 VDD1 VDD1.n3 0.409983
R88 B.n496 B.n495 585
R89 B.n497 B.n496 585
R90 B.n174 B.n85 585
R91 B.n173 B.n172 585
R92 B.n171 B.n170 585
R93 B.n169 B.n168 585
R94 B.n167 B.n166 585
R95 B.n165 B.n164 585
R96 B.n163 B.n162 585
R97 B.n161 B.n160 585
R98 B.n159 B.n158 585
R99 B.n157 B.n156 585
R100 B.n155 B.n154 585
R101 B.n153 B.n152 585
R102 B.n151 B.n150 585
R103 B.n149 B.n148 585
R104 B.n147 B.n146 585
R105 B.n145 B.n144 585
R106 B.n143 B.n142 585
R107 B.n141 B.n140 585
R108 B.n139 B.n138 585
R109 B.n137 B.n136 585
R110 B.n135 B.n134 585
R111 B.n133 B.n132 585
R112 B.n131 B.n130 585
R113 B.n129 B.n128 585
R114 B.n127 B.n126 585
R115 B.n124 B.n123 585
R116 B.n122 B.n121 585
R117 B.n120 B.n119 585
R118 B.n118 B.n117 585
R119 B.n116 B.n115 585
R120 B.n114 B.n113 585
R121 B.n112 B.n111 585
R122 B.n110 B.n109 585
R123 B.n108 B.n107 585
R124 B.n106 B.n105 585
R125 B.n104 B.n103 585
R126 B.n102 B.n101 585
R127 B.n100 B.n99 585
R128 B.n98 B.n97 585
R129 B.n96 B.n95 585
R130 B.n94 B.n93 585
R131 B.n92 B.n91 585
R132 B.n494 B.n63 585
R133 B.n498 B.n63 585
R134 B.n493 B.n62 585
R135 B.n499 B.n62 585
R136 B.n492 B.n491 585
R137 B.n491 B.n58 585
R138 B.n490 B.n57 585
R139 B.n505 B.n57 585
R140 B.n489 B.n56 585
R141 B.n506 B.n56 585
R142 B.n488 B.n55 585
R143 B.n507 B.n55 585
R144 B.n487 B.n486 585
R145 B.n486 B.n54 585
R146 B.n485 B.n50 585
R147 B.n513 B.n50 585
R148 B.n484 B.n49 585
R149 B.n514 B.n49 585
R150 B.n483 B.n48 585
R151 B.n515 B.n48 585
R152 B.n482 B.n481 585
R153 B.n481 B.n44 585
R154 B.n480 B.n43 585
R155 B.n521 B.n43 585
R156 B.n479 B.n42 585
R157 B.n522 B.n42 585
R158 B.n478 B.n41 585
R159 B.n523 B.n41 585
R160 B.n477 B.n476 585
R161 B.n476 B.n37 585
R162 B.n475 B.n36 585
R163 B.n529 B.n36 585
R164 B.n474 B.n35 585
R165 B.n530 B.n35 585
R166 B.n473 B.n34 585
R167 B.n531 B.n34 585
R168 B.n472 B.n471 585
R169 B.n471 B.n30 585
R170 B.n470 B.n29 585
R171 B.n537 B.n29 585
R172 B.n469 B.n28 585
R173 B.n538 B.n28 585
R174 B.n468 B.n27 585
R175 B.n539 B.n27 585
R176 B.n467 B.n466 585
R177 B.n466 B.n26 585
R178 B.n465 B.n22 585
R179 B.n545 B.n22 585
R180 B.n464 B.n21 585
R181 B.n546 B.n21 585
R182 B.n463 B.n20 585
R183 B.n547 B.n20 585
R184 B.n462 B.n461 585
R185 B.n461 B.n16 585
R186 B.n460 B.n15 585
R187 B.n553 B.n15 585
R188 B.n459 B.n14 585
R189 B.n554 B.n14 585
R190 B.n458 B.n13 585
R191 B.n555 B.n13 585
R192 B.n457 B.n456 585
R193 B.n456 B.n12 585
R194 B.n455 B.n454 585
R195 B.n455 B.n8 585
R196 B.n453 B.n7 585
R197 B.n562 B.n7 585
R198 B.n452 B.n6 585
R199 B.n563 B.n6 585
R200 B.n451 B.n5 585
R201 B.n564 B.n5 585
R202 B.n450 B.n449 585
R203 B.n449 B.n4 585
R204 B.n448 B.n175 585
R205 B.n448 B.n447 585
R206 B.n438 B.n176 585
R207 B.n177 B.n176 585
R208 B.n440 B.n439 585
R209 B.n441 B.n440 585
R210 B.n437 B.n181 585
R211 B.n185 B.n181 585
R212 B.n436 B.n435 585
R213 B.n435 B.n434 585
R214 B.n183 B.n182 585
R215 B.n184 B.n183 585
R216 B.n427 B.n426 585
R217 B.n428 B.n427 585
R218 B.n425 B.n190 585
R219 B.n190 B.n189 585
R220 B.n424 B.n423 585
R221 B.n423 B.n422 585
R222 B.n192 B.n191 585
R223 B.n415 B.n192 585
R224 B.n414 B.n413 585
R225 B.n416 B.n414 585
R226 B.n412 B.n197 585
R227 B.n197 B.n196 585
R228 B.n411 B.n410 585
R229 B.n410 B.n409 585
R230 B.n199 B.n198 585
R231 B.n200 B.n199 585
R232 B.n402 B.n401 585
R233 B.n403 B.n402 585
R234 B.n400 B.n205 585
R235 B.n205 B.n204 585
R236 B.n399 B.n398 585
R237 B.n398 B.n397 585
R238 B.n207 B.n206 585
R239 B.n208 B.n207 585
R240 B.n390 B.n389 585
R241 B.n391 B.n390 585
R242 B.n388 B.n213 585
R243 B.n213 B.n212 585
R244 B.n387 B.n386 585
R245 B.n386 B.n385 585
R246 B.n215 B.n214 585
R247 B.n216 B.n215 585
R248 B.n378 B.n377 585
R249 B.n379 B.n378 585
R250 B.n376 B.n221 585
R251 B.n221 B.n220 585
R252 B.n375 B.n374 585
R253 B.n374 B.n373 585
R254 B.n223 B.n222 585
R255 B.n366 B.n223 585
R256 B.n365 B.n364 585
R257 B.n367 B.n365 585
R258 B.n363 B.n228 585
R259 B.n228 B.n227 585
R260 B.n362 B.n361 585
R261 B.n361 B.n360 585
R262 B.n230 B.n229 585
R263 B.n231 B.n230 585
R264 B.n353 B.n352 585
R265 B.n354 B.n353 585
R266 B.n351 B.n236 585
R267 B.n236 B.n235 585
R268 B.n345 B.n344 585
R269 B.n343 B.n259 585
R270 B.n342 B.n258 585
R271 B.n347 B.n258 585
R272 B.n341 B.n340 585
R273 B.n339 B.n338 585
R274 B.n337 B.n336 585
R275 B.n335 B.n334 585
R276 B.n333 B.n332 585
R277 B.n331 B.n330 585
R278 B.n329 B.n328 585
R279 B.n327 B.n326 585
R280 B.n325 B.n324 585
R281 B.n323 B.n322 585
R282 B.n321 B.n320 585
R283 B.n319 B.n318 585
R284 B.n317 B.n316 585
R285 B.n315 B.n314 585
R286 B.n313 B.n312 585
R287 B.n311 B.n310 585
R288 B.n309 B.n308 585
R289 B.n307 B.n306 585
R290 B.n305 B.n304 585
R291 B.n303 B.n302 585
R292 B.n301 B.n300 585
R293 B.n299 B.n298 585
R294 B.n297 B.n296 585
R295 B.n294 B.n293 585
R296 B.n292 B.n291 585
R297 B.n290 B.n289 585
R298 B.n288 B.n287 585
R299 B.n286 B.n285 585
R300 B.n284 B.n283 585
R301 B.n282 B.n281 585
R302 B.n280 B.n279 585
R303 B.n278 B.n277 585
R304 B.n276 B.n275 585
R305 B.n274 B.n273 585
R306 B.n272 B.n271 585
R307 B.n270 B.n269 585
R308 B.n268 B.n267 585
R309 B.n266 B.n265 585
R310 B.n238 B.n237 585
R311 B.n350 B.n349 585
R312 B.n234 B.n233 585
R313 B.n235 B.n234 585
R314 B.n356 B.n355 585
R315 B.n355 B.n354 585
R316 B.n357 B.n232 585
R317 B.n232 B.n231 585
R318 B.n359 B.n358 585
R319 B.n360 B.n359 585
R320 B.n226 B.n225 585
R321 B.n227 B.n226 585
R322 B.n369 B.n368 585
R323 B.n368 B.n367 585
R324 B.n370 B.n224 585
R325 B.n366 B.n224 585
R326 B.n372 B.n371 585
R327 B.n373 B.n372 585
R328 B.n219 B.n218 585
R329 B.n220 B.n219 585
R330 B.n381 B.n380 585
R331 B.n380 B.n379 585
R332 B.n382 B.n217 585
R333 B.n217 B.n216 585
R334 B.n384 B.n383 585
R335 B.n385 B.n384 585
R336 B.n211 B.n210 585
R337 B.n212 B.n211 585
R338 B.n393 B.n392 585
R339 B.n392 B.n391 585
R340 B.n394 B.n209 585
R341 B.n209 B.n208 585
R342 B.n396 B.n395 585
R343 B.n397 B.n396 585
R344 B.n203 B.n202 585
R345 B.n204 B.n203 585
R346 B.n405 B.n404 585
R347 B.n404 B.n403 585
R348 B.n406 B.n201 585
R349 B.n201 B.n200 585
R350 B.n408 B.n407 585
R351 B.n409 B.n408 585
R352 B.n195 B.n194 585
R353 B.n196 B.n195 585
R354 B.n418 B.n417 585
R355 B.n417 B.n416 585
R356 B.n419 B.n193 585
R357 B.n415 B.n193 585
R358 B.n421 B.n420 585
R359 B.n422 B.n421 585
R360 B.n188 B.n187 585
R361 B.n189 B.n188 585
R362 B.n430 B.n429 585
R363 B.n429 B.n428 585
R364 B.n431 B.n186 585
R365 B.n186 B.n184 585
R366 B.n433 B.n432 585
R367 B.n434 B.n433 585
R368 B.n180 B.n179 585
R369 B.n185 B.n180 585
R370 B.n443 B.n442 585
R371 B.n442 B.n441 585
R372 B.n444 B.n178 585
R373 B.n178 B.n177 585
R374 B.n446 B.n445 585
R375 B.n447 B.n446 585
R376 B.n3 B.n0 585
R377 B.n4 B.n3 585
R378 B.n561 B.n1 585
R379 B.n562 B.n561 585
R380 B.n560 B.n559 585
R381 B.n560 B.n8 585
R382 B.n558 B.n9 585
R383 B.n12 B.n9 585
R384 B.n557 B.n556 585
R385 B.n556 B.n555 585
R386 B.n11 B.n10 585
R387 B.n554 B.n11 585
R388 B.n552 B.n551 585
R389 B.n553 B.n552 585
R390 B.n550 B.n17 585
R391 B.n17 B.n16 585
R392 B.n549 B.n548 585
R393 B.n548 B.n547 585
R394 B.n19 B.n18 585
R395 B.n546 B.n19 585
R396 B.n544 B.n543 585
R397 B.n545 B.n544 585
R398 B.n542 B.n23 585
R399 B.n26 B.n23 585
R400 B.n541 B.n540 585
R401 B.n540 B.n539 585
R402 B.n25 B.n24 585
R403 B.n538 B.n25 585
R404 B.n536 B.n535 585
R405 B.n537 B.n536 585
R406 B.n534 B.n31 585
R407 B.n31 B.n30 585
R408 B.n533 B.n532 585
R409 B.n532 B.n531 585
R410 B.n33 B.n32 585
R411 B.n530 B.n33 585
R412 B.n528 B.n527 585
R413 B.n529 B.n528 585
R414 B.n526 B.n38 585
R415 B.n38 B.n37 585
R416 B.n525 B.n524 585
R417 B.n524 B.n523 585
R418 B.n40 B.n39 585
R419 B.n522 B.n40 585
R420 B.n520 B.n519 585
R421 B.n521 B.n520 585
R422 B.n518 B.n45 585
R423 B.n45 B.n44 585
R424 B.n517 B.n516 585
R425 B.n516 B.n515 585
R426 B.n47 B.n46 585
R427 B.n514 B.n47 585
R428 B.n512 B.n511 585
R429 B.n513 B.n512 585
R430 B.n510 B.n51 585
R431 B.n54 B.n51 585
R432 B.n509 B.n508 585
R433 B.n508 B.n507 585
R434 B.n53 B.n52 585
R435 B.n506 B.n53 585
R436 B.n504 B.n503 585
R437 B.n505 B.n504 585
R438 B.n502 B.n59 585
R439 B.n59 B.n58 585
R440 B.n501 B.n500 585
R441 B.n500 B.n499 585
R442 B.n61 B.n60 585
R443 B.n498 B.n61 585
R444 B.n565 B.n564 585
R445 B.n563 B.n2 585
R446 B.n91 B.n61 559.769
R447 B.n496 B.n63 559.769
R448 B.n349 B.n236 559.769
R449 B.n345 B.n234 559.769
R450 B.n497 B.n84 256.663
R451 B.n497 B.n83 256.663
R452 B.n497 B.n82 256.663
R453 B.n497 B.n81 256.663
R454 B.n497 B.n80 256.663
R455 B.n497 B.n79 256.663
R456 B.n497 B.n78 256.663
R457 B.n497 B.n77 256.663
R458 B.n497 B.n76 256.663
R459 B.n497 B.n75 256.663
R460 B.n497 B.n74 256.663
R461 B.n497 B.n73 256.663
R462 B.n497 B.n72 256.663
R463 B.n497 B.n71 256.663
R464 B.n497 B.n70 256.663
R465 B.n497 B.n69 256.663
R466 B.n497 B.n68 256.663
R467 B.n497 B.n67 256.663
R468 B.n497 B.n66 256.663
R469 B.n497 B.n65 256.663
R470 B.n497 B.n64 256.663
R471 B.n347 B.n346 256.663
R472 B.n347 B.n239 256.663
R473 B.n347 B.n240 256.663
R474 B.n347 B.n241 256.663
R475 B.n347 B.n242 256.663
R476 B.n347 B.n243 256.663
R477 B.n347 B.n244 256.663
R478 B.n347 B.n245 256.663
R479 B.n347 B.n246 256.663
R480 B.n347 B.n247 256.663
R481 B.n347 B.n248 256.663
R482 B.n347 B.n249 256.663
R483 B.n347 B.n250 256.663
R484 B.n347 B.n251 256.663
R485 B.n347 B.n252 256.663
R486 B.n347 B.n253 256.663
R487 B.n347 B.n254 256.663
R488 B.n347 B.n255 256.663
R489 B.n347 B.n256 256.663
R490 B.n347 B.n257 256.663
R491 B.n348 B.n347 256.663
R492 B.n567 B.n566 256.663
R493 B.n89 B.t13 253.798
R494 B.n86 B.t17 253.798
R495 B.n263 B.t6 253.798
R496 B.n260 B.t10 253.798
R497 B.n347 B.n235 164.661
R498 B.n498 B.n497 164.661
R499 B.n95 B.n94 163.367
R500 B.n99 B.n98 163.367
R501 B.n103 B.n102 163.367
R502 B.n107 B.n106 163.367
R503 B.n111 B.n110 163.367
R504 B.n115 B.n114 163.367
R505 B.n119 B.n118 163.367
R506 B.n123 B.n122 163.367
R507 B.n128 B.n127 163.367
R508 B.n132 B.n131 163.367
R509 B.n136 B.n135 163.367
R510 B.n140 B.n139 163.367
R511 B.n144 B.n143 163.367
R512 B.n148 B.n147 163.367
R513 B.n152 B.n151 163.367
R514 B.n156 B.n155 163.367
R515 B.n160 B.n159 163.367
R516 B.n164 B.n163 163.367
R517 B.n168 B.n167 163.367
R518 B.n172 B.n171 163.367
R519 B.n496 B.n85 163.367
R520 B.n353 B.n236 163.367
R521 B.n353 B.n230 163.367
R522 B.n361 B.n230 163.367
R523 B.n361 B.n228 163.367
R524 B.n365 B.n228 163.367
R525 B.n365 B.n223 163.367
R526 B.n374 B.n223 163.367
R527 B.n374 B.n221 163.367
R528 B.n378 B.n221 163.367
R529 B.n378 B.n215 163.367
R530 B.n386 B.n215 163.367
R531 B.n386 B.n213 163.367
R532 B.n390 B.n213 163.367
R533 B.n390 B.n207 163.367
R534 B.n398 B.n207 163.367
R535 B.n398 B.n205 163.367
R536 B.n402 B.n205 163.367
R537 B.n402 B.n199 163.367
R538 B.n410 B.n199 163.367
R539 B.n410 B.n197 163.367
R540 B.n414 B.n197 163.367
R541 B.n414 B.n192 163.367
R542 B.n423 B.n192 163.367
R543 B.n423 B.n190 163.367
R544 B.n427 B.n190 163.367
R545 B.n427 B.n183 163.367
R546 B.n435 B.n183 163.367
R547 B.n435 B.n181 163.367
R548 B.n440 B.n181 163.367
R549 B.n440 B.n176 163.367
R550 B.n448 B.n176 163.367
R551 B.n449 B.n448 163.367
R552 B.n449 B.n5 163.367
R553 B.n6 B.n5 163.367
R554 B.n7 B.n6 163.367
R555 B.n455 B.n7 163.367
R556 B.n456 B.n455 163.367
R557 B.n456 B.n13 163.367
R558 B.n14 B.n13 163.367
R559 B.n15 B.n14 163.367
R560 B.n461 B.n15 163.367
R561 B.n461 B.n20 163.367
R562 B.n21 B.n20 163.367
R563 B.n22 B.n21 163.367
R564 B.n466 B.n22 163.367
R565 B.n466 B.n27 163.367
R566 B.n28 B.n27 163.367
R567 B.n29 B.n28 163.367
R568 B.n471 B.n29 163.367
R569 B.n471 B.n34 163.367
R570 B.n35 B.n34 163.367
R571 B.n36 B.n35 163.367
R572 B.n476 B.n36 163.367
R573 B.n476 B.n41 163.367
R574 B.n42 B.n41 163.367
R575 B.n43 B.n42 163.367
R576 B.n481 B.n43 163.367
R577 B.n481 B.n48 163.367
R578 B.n49 B.n48 163.367
R579 B.n50 B.n49 163.367
R580 B.n486 B.n50 163.367
R581 B.n486 B.n55 163.367
R582 B.n56 B.n55 163.367
R583 B.n57 B.n56 163.367
R584 B.n491 B.n57 163.367
R585 B.n491 B.n62 163.367
R586 B.n63 B.n62 163.367
R587 B.n259 B.n258 163.367
R588 B.n340 B.n258 163.367
R589 B.n338 B.n337 163.367
R590 B.n334 B.n333 163.367
R591 B.n330 B.n329 163.367
R592 B.n326 B.n325 163.367
R593 B.n322 B.n321 163.367
R594 B.n318 B.n317 163.367
R595 B.n314 B.n313 163.367
R596 B.n310 B.n309 163.367
R597 B.n306 B.n305 163.367
R598 B.n302 B.n301 163.367
R599 B.n298 B.n297 163.367
R600 B.n293 B.n292 163.367
R601 B.n289 B.n288 163.367
R602 B.n285 B.n284 163.367
R603 B.n281 B.n280 163.367
R604 B.n277 B.n276 163.367
R605 B.n273 B.n272 163.367
R606 B.n269 B.n268 163.367
R607 B.n265 B.n238 163.367
R608 B.n355 B.n234 163.367
R609 B.n355 B.n232 163.367
R610 B.n359 B.n232 163.367
R611 B.n359 B.n226 163.367
R612 B.n368 B.n226 163.367
R613 B.n368 B.n224 163.367
R614 B.n372 B.n224 163.367
R615 B.n372 B.n219 163.367
R616 B.n380 B.n219 163.367
R617 B.n380 B.n217 163.367
R618 B.n384 B.n217 163.367
R619 B.n384 B.n211 163.367
R620 B.n392 B.n211 163.367
R621 B.n392 B.n209 163.367
R622 B.n396 B.n209 163.367
R623 B.n396 B.n203 163.367
R624 B.n404 B.n203 163.367
R625 B.n404 B.n201 163.367
R626 B.n408 B.n201 163.367
R627 B.n408 B.n195 163.367
R628 B.n417 B.n195 163.367
R629 B.n417 B.n193 163.367
R630 B.n421 B.n193 163.367
R631 B.n421 B.n188 163.367
R632 B.n429 B.n188 163.367
R633 B.n429 B.n186 163.367
R634 B.n433 B.n186 163.367
R635 B.n433 B.n180 163.367
R636 B.n442 B.n180 163.367
R637 B.n442 B.n178 163.367
R638 B.n446 B.n178 163.367
R639 B.n446 B.n3 163.367
R640 B.n565 B.n3 163.367
R641 B.n561 B.n2 163.367
R642 B.n561 B.n560 163.367
R643 B.n560 B.n9 163.367
R644 B.n556 B.n9 163.367
R645 B.n556 B.n11 163.367
R646 B.n552 B.n11 163.367
R647 B.n552 B.n17 163.367
R648 B.n548 B.n17 163.367
R649 B.n548 B.n19 163.367
R650 B.n544 B.n19 163.367
R651 B.n544 B.n23 163.367
R652 B.n540 B.n23 163.367
R653 B.n540 B.n25 163.367
R654 B.n536 B.n25 163.367
R655 B.n536 B.n31 163.367
R656 B.n532 B.n31 163.367
R657 B.n532 B.n33 163.367
R658 B.n528 B.n33 163.367
R659 B.n528 B.n38 163.367
R660 B.n524 B.n38 163.367
R661 B.n524 B.n40 163.367
R662 B.n520 B.n40 163.367
R663 B.n520 B.n45 163.367
R664 B.n516 B.n45 163.367
R665 B.n516 B.n47 163.367
R666 B.n512 B.n47 163.367
R667 B.n512 B.n51 163.367
R668 B.n508 B.n51 163.367
R669 B.n508 B.n53 163.367
R670 B.n504 B.n53 163.367
R671 B.n504 B.n59 163.367
R672 B.n500 B.n59 163.367
R673 B.n500 B.n61 163.367
R674 B.n86 B.t18 118.603
R675 B.n263 B.t9 118.603
R676 B.n89 B.t15 118.602
R677 B.n260 B.t12 118.602
R678 B.n354 B.n235 84.1873
R679 B.n354 B.n231 84.1873
R680 B.n360 B.n231 84.1873
R681 B.n360 B.n227 84.1873
R682 B.n367 B.n227 84.1873
R683 B.n367 B.n366 84.1873
R684 B.n373 B.n220 84.1873
R685 B.n379 B.n220 84.1873
R686 B.n379 B.n216 84.1873
R687 B.n385 B.n216 84.1873
R688 B.n385 B.n212 84.1873
R689 B.n391 B.n212 84.1873
R690 B.n391 B.n208 84.1873
R691 B.n397 B.n208 84.1873
R692 B.n403 B.n204 84.1873
R693 B.n403 B.n200 84.1873
R694 B.n409 B.n200 84.1873
R695 B.n409 B.n196 84.1873
R696 B.n416 B.n196 84.1873
R697 B.n416 B.n415 84.1873
R698 B.n422 B.n189 84.1873
R699 B.n428 B.n189 84.1873
R700 B.n428 B.n184 84.1873
R701 B.n434 B.n184 84.1873
R702 B.n434 B.n185 84.1873
R703 B.n441 B.n177 84.1873
R704 B.n447 B.n177 84.1873
R705 B.n447 B.n4 84.1873
R706 B.n564 B.n4 84.1873
R707 B.n564 B.n563 84.1873
R708 B.n563 B.n562 84.1873
R709 B.n562 B.n8 84.1873
R710 B.n12 B.n8 84.1873
R711 B.n555 B.n12 84.1873
R712 B.n554 B.n553 84.1873
R713 B.n553 B.n16 84.1873
R714 B.n547 B.n16 84.1873
R715 B.n547 B.n546 84.1873
R716 B.n546 B.n545 84.1873
R717 B.n539 B.n26 84.1873
R718 B.n539 B.n538 84.1873
R719 B.n538 B.n537 84.1873
R720 B.n537 B.n30 84.1873
R721 B.n531 B.n30 84.1873
R722 B.n531 B.n530 84.1873
R723 B.n529 B.n37 84.1873
R724 B.n523 B.n37 84.1873
R725 B.n523 B.n522 84.1873
R726 B.n522 B.n521 84.1873
R727 B.n521 B.n44 84.1873
R728 B.n515 B.n44 84.1873
R729 B.n515 B.n514 84.1873
R730 B.n514 B.n513 84.1873
R731 B.n507 B.n54 84.1873
R732 B.n507 B.n506 84.1873
R733 B.n506 B.n505 84.1873
R734 B.n505 B.n58 84.1873
R735 B.n499 B.n58 84.1873
R736 B.n499 B.n498 84.1873
R737 B.n397 B.t3 79.2352
R738 B.t4 B.n529 79.2352
R739 B.n87 B.t19 76.5191
R740 B.n264 B.t8 76.5191
R741 B.n90 B.t16 76.5161
R742 B.n261 B.t11 76.5161
R743 B.n91 B.n64 71.676
R744 B.n95 B.n65 71.676
R745 B.n99 B.n66 71.676
R746 B.n103 B.n67 71.676
R747 B.n107 B.n68 71.676
R748 B.n111 B.n69 71.676
R749 B.n115 B.n70 71.676
R750 B.n119 B.n71 71.676
R751 B.n123 B.n72 71.676
R752 B.n128 B.n73 71.676
R753 B.n132 B.n74 71.676
R754 B.n136 B.n75 71.676
R755 B.n140 B.n76 71.676
R756 B.n144 B.n77 71.676
R757 B.n148 B.n78 71.676
R758 B.n152 B.n79 71.676
R759 B.n156 B.n80 71.676
R760 B.n160 B.n81 71.676
R761 B.n164 B.n82 71.676
R762 B.n168 B.n83 71.676
R763 B.n172 B.n84 71.676
R764 B.n85 B.n84 71.676
R765 B.n171 B.n83 71.676
R766 B.n167 B.n82 71.676
R767 B.n163 B.n81 71.676
R768 B.n159 B.n80 71.676
R769 B.n155 B.n79 71.676
R770 B.n151 B.n78 71.676
R771 B.n147 B.n77 71.676
R772 B.n143 B.n76 71.676
R773 B.n139 B.n75 71.676
R774 B.n135 B.n74 71.676
R775 B.n131 B.n73 71.676
R776 B.n127 B.n72 71.676
R777 B.n122 B.n71 71.676
R778 B.n118 B.n70 71.676
R779 B.n114 B.n69 71.676
R780 B.n110 B.n68 71.676
R781 B.n106 B.n67 71.676
R782 B.n102 B.n66 71.676
R783 B.n98 B.n65 71.676
R784 B.n94 B.n64 71.676
R785 B.n346 B.n345 71.676
R786 B.n340 B.n239 71.676
R787 B.n337 B.n240 71.676
R788 B.n333 B.n241 71.676
R789 B.n329 B.n242 71.676
R790 B.n325 B.n243 71.676
R791 B.n321 B.n244 71.676
R792 B.n317 B.n245 71.676
R793 B.n313 B.n246 71.676
R794 B.n309 B.n247 71.676
R795 B.n305 B.n248 71.676
R796 B.n301 B.n249 71.676
R797 B.n297 B.n250 71.676
R798 B.n292 B.n251 71.676
R799 B.n288 B.n252 71.676
R800 B.n284 B.n253 71.676
R801 B.n280 B.n254 71.676
R802 B.n276 B.n255 71.676
R803 B.n272 B.n256 71.676
R804 B.n268 B.n257 71.676
R805 B.n348 B.n238 71.676
R806 B.n346 B.n259 71.676
R807 B.n338 B.n239 71.676
R808 B.n334 B.n240 71.676
R809 B.n330 B.n241 71.676
R810 B.n326 B.n242 71.676
R811 B.n322 B.n243 71.676
R812 B.n318 B.n244 71.676
R813 B.n314 B.n245 71.676
R814 B.n310 B.n246 71.676
R815 B.n306 B.n247 71.676
R816 B.n302 B.n248 71.676
R817 B.n298 B.n249 71.676
R818 B.n293 B.n250 71.676
R819 B.n289 B.n251 71.676
R820 B.n285 B.n252 71.676
R821 B.n281 B.n253 71.676
R822 B.n277 B.n254 71.676
R823 B.n273 B.n255 71.676
R824 B.n269 B.n256 71.676
R825 B.n265 B.n257 71.676
R826 B.n349 B.n348 71.676
R827 B.n566 B.n565 71.676
R828 B.n566 B.n2 71.676
R829 B.n125 B.n90 59.5399
R830 B.n88 B.n87 59.5399
R831 B.n295 B.n264 59.5399
R832 B.n262 B.n261 59.5399
R833 B.n185 B.t5 59.4265
R834 B.t1 B.n554 59.4265
R835 B.n422 B.t0 56.9504
R836 B.n545 B.t2 56.9504
R837 B.n373 B.t7 54.4743
R838 B.n513 B.t14 54.4743
R839 B.n90 B.n89 42.0853
R840 B.n87 B.n86 42.0853
R841 B.n264 B.n263 42.0853
R842 B.n261 B.n260 42.0853
R843 B.n344 B.n233 36.3712
R844 B.n351 B.n350 36.3712
R845 B.n92 B.n60 36.3712
R846 B.n495 B.n494 36.3712
R847 B.n366 B.t7 29.7135
R848 B.n54 B.t14 29.7135
R849 B.n415 B.t0 27.2374
R850 B.n26 B.t2 27.2374
R851 B.n441 B.t5 24.7613
R852 B.n555 B.t1 24.7613
R853 B B.n567 18.0485
R854 B.n356 B.n233 10.6151
R855 B.n357 B.n356 10.6151
R856 B.n358 B.n357 10.6151
R857 B.n358 B.n225 10.6151
R858 B.n369 B.n225 10.6151
R859 B.n370 B.n369 10.6151
R860 B.n371 B.n370 10.6151
R861 B.n371 B.n218 10.6151
R862 B.n381 B.n218 10.6151
R863 B.n382 B.n381 10.6151
R864 B.n383 B.n382 10.6151
R865 B.n383 B.n210 10.6151
R866 B.n393 B.n210 10.6151
R867 B.n394 B.n393 10.6151
R868 B.n395 B.n394 10.6151
R869 B.n395 B.n202 10.6151
R870 B.n405 B.n202 10.6151
R871 B.n406 B.n405 10.6151
R872 B.n407 B.n406 10.6151
R873 B.n407 B.n194 10.6151
R874 B.n418 B.n194 10.6151
R875 B.n419 B.n418 10.6151
R876 B.n420 B.n419 10.6151
R877 B.n420 B.n187 10.6151
R878 B.n430 B.n187 10.6151
R879 B.n431 B.n430 10.6151
R880 B.n432 B.n431 10.6151
R881 B.n432 B.n179 10.6151
R882 B.n443 B.n179 10.6151
R883 B.n444 B.n443 10.6151
R884 B.n445 B.n444 10.6151
R885 B.n445 B.n0 10.6151
R886 B.n344 B.n343 10.6151
R887 B.n343 B.n342 10.6151
R888 B.n342 B.n341 10.6151
R889 B.n341 B.n339 10.6151
R890 B.n339 B.n336 10.6151
R891 B.n336 B.n335 10.6151
R892 B.n335 B.n332 10.6151
R893 B.n332 B.n331 10.6151
R894 B.n331 B.n328 10.6151
R895 B.n328 B.n327 10.6151
R896 B.n327 B.n324 10.6151
R897 B.n324 B.n323 10.6151
R898 B.n323 B.n320 10.6151
R899 B.n320 B.n319 10.6151
R900 B.n319 B.n316 10.6151
R901 B.n316 B.n315 10.6151
R902 B.n312 B.n311 10.6151
R903 B.n311 B.n308 10.6151
R904 B.n308 B.n307 10.6151
R905 B.n307 B.n304 10.6151
R906 B.n304 B.n303 10.6151
R907 B.n303 B.n300 10.6151
R908 B.n300 B.n299 10.6151
R909 B.n299 B.n296 10.6151
R910 B.n294 B.n291 10.6151
R911 B.n291 B.n290 10.6151
R912 B.n290 B.n287 10.6151
R913 B.n287 B.n286 10.6151
R914 B.n286 B.n283 10.6151
R915 B.n283 B.n282 10.6151
R916 B.n282 B.n279 10.6151
R917 B.n279 B.n278 10.6151
R918 B.n278 B.n275 10.6151
R919 B.n275 B.n274 10.6151
R920 B.n274 B.n271 10.6151
R921 B.n271 B.n270 10.6151
R922 B.n270 B.n267 10.6151
R923 B.n267 B.n266 10.6151
R924 B.n266 B.n237 10.6151
R925 B.n350 B.n237 10.6151
R926 B.n352 B.n351 10.6151
R927 B.n352 B.n229 10.6151
R928 B.n362 B.n229 10.6151
R929 B.n363 B.n362 10.6151
R930 B.n364 B.n363 10.6151
R931 B.n364 B.n222 10.6151
R932 B.n375 B.n222 10.6151
R933 B.n376 B.n375 10.6151
R934 B.n377 B.n376 10.6151
R935 B.n377 B.n214 10.6151
R936 B.n387 B.n214 10.6151
R937 B.n388 B.n387 10.6151
R938 B.n389 B.n388 10.6151
R939 B.n389 B.n206 10.6151
R940 B.n399 B.n206 10.6151
R941 B.n400 B.n399 10.6151
R942 B.n401 B.n400 10.6151
R943 B.n401 B.n198 10.6151
R944 B.n411 B.n198 10.6151
R945 B.n412 B.n411 10.6151
R946 B.n413 B.n412 10.6151
R947 B.n413 B.n191 10.6151
R948 B.n424 B.n191 10.6151
R949 B.n425 B.n424 10.6151
R950 B.n426 B.n425 10.6151
R951 B.n426 B.n182 10.6151
R952 B.n436 B.n182 10.6151
R953 B.n437 B.n436 10.6151
R954 B.n439 B.n437 10.6151
R955 B.n439 B.n438 10.6151
R956 B.n438 B.n175 10.6151
R957 B.n450 B.n175 10.6151
R958 B.n451 B.n450 10.6151
R959 B.n452 B.n451 10.6151
R960 B.n453 B.n452 10.6151
R961 B.n454 B.n453 10.6151
R962 B.n457 B.n454 10.6151
R963 B.n458 B.n457 10.6151
R964 B.n459 B.n458 10.6151
R965 B.n460 B.n459 10.6151
R966 B.n462 B.n460 10.6151
R967 B.n463 B.n462 10.6151
R968 B.n464 B.n463 10.6151
R969 B.n465 B.n464 10.6151
R970 B.n467 B.n465 10.6151
R971 B.n468 B.n467 10.6151
R972 B.n469 B.n468 10.6151
R973 B.n470 B.n469 10.6151
R974 B.n472 B.n470 10.6151
R975 B.n473 B.n472 10.6151
R976 B.n474 B.n473 10.6151
R977 B.n475 B.n474 10.6151
R978 B.n477 B.n475 10.6151
R979 B.n478 B.n477 10.6151
R980 B.n479 B.n478 10.6151
R981 B.n480 B.n479 10.6151
R982 B.n482 B.n480 10.6151
R983 B.n483 B.n482 10.6151
R984 B.n484 B.n483 10.6151
R985 B.n485 B.n484 10.6151
R986 B.n487 B.n485 10.6151
R987 B.n488 B.n487 10.6151
R988 B.n489 B.n488 10.6151
R989 B.n490 B.n489 10.6151
R990 B.n492 B.n490 10.6151
R991 B.n493 B.n492 10.6151
R992 B.n494 B.n493 10.6151
R993 B.n559 B.n1 10.6151
R994 B.n559 B.n558 10.6151
R995 B.n558 B.n557 10.6151
R996 B.n557 B.n10 10.6151
R997 B.n551 B.n10 10.6151
R998 B.n551 B.n550 10.6151
R999 B.n550 B.n549 10.6151
R1000 B.n549 B.n18 10.6151
R1001 B.n543 B.n18 10.6151
R1002 B.n543 B.n542 10.6151
R1003 B.n542 B.n541 10.6151
R1004 B.n541 B.n24 10.6151
R1005 B.n535 B.n24 10.6151
R1006 B.n535 B.n534 10.6151
R1007 B.n534 B.n533 10.6151
R1008 B.n533 B.n32 10.6151
R1009 B.n527 B.n32 10.6151
R1010 B.n527 B.n526 10.6151
R1011 B.n526 B.n525 10.6151
R1012 B.n525 B.n39 10.6151
R1013 B.n519 B.n39 10.6151
R1014 B.n519 B.n518 10.6151
R1015 B.n518 B.n517 10.6151
R1016 B.n517 B.n46 10.6151
R1017 B.n511 B.n46 10.6151
R1018 B.n511 B.n510 10.6151
R1019 B.n510 B.n509 10.6151
R1020 B.n509 B.n52 10.6151
R1021 B.n503 B.n52 10.6151
R1022 B.n503 B.n502 10.6151
R1023 B.n502 B.n501 10.6151
R1024 B.n501 B.n60 10.6151
R1025 B.n93 B.n92 10.6151
R1026 B.n96 B.n93 10.6151
R1027 B.n97 B.n96 10.6151
R1028 B.n100 B.n97 10.6151
R1029 B.n101 B.n100 10.6151
R1030 B.n104 B.n101 10.6151
R1031 B.n105 B.n104 10.6151
R1032 B.n108 B.n105 10.6151
R1033 B.n109 B.n108 10.6151
R1034 B.n112 B.n109 10.6151
R1035 B.n113 B.n112 10.6151
R1036 B.n116 B.n113 10.6151
R1037 B.n117 B.n116 10.6151
R1038 B.n120 B.n117 10.6151
R1039 B.n121 B.n120 10.6151
R1040 B.n124 B.n121 10.6151
R1041 B.n129 B.n126 10.6151
R1042 B.n130 B.n129 10.6151
R1043 B.n133 B.n130 10.6151
R1044 B.n134 B.n133 10.6151
R1045 B.n137 B.n134 10.6151
R1046 B.n138 B.n137 10.6151
R1047 B.n141 B.n138 10.6151
R1048 B.n142 B.n141 10.6151
R1049 B.n146 B.n145 10.6151
R1050 B.n149 B.n146 10.6151
R1051 B.n150 B.n149 10.6151
R1052 B.n153 B.n150 10.6151
R1053 B.n154 B.n153 10.6151
R1054 B.n157 B.n154 10.6151
R1055 B.n158 B.n157 10.6151
R1056 B.n161 B.n158 10.6151
R1057 B.n162 B.n161 10.6151
R1058 B.n165 B.n162 10.6151
R1059 B.n166 B.n165 10.6151
R1060 B.n169 B.n166 10.6151
R1061 B.n170 B.n169 10.6151
R1062 B.n173 B.n170 10.6151
R1063 B.n174 B.n173 10.6151
R1064 B.n495 B.n174 10.6151
R1065 B.n567 B.n0 8.11757
R1066 B.n567 B.n1 8.11757
R1067 B.n312 B.n262 6.5566
R1068 B.n296 B.n295 6.5566
R1069 B.n126 B.n125 6.5566
R1070 B.n142 B.n88 6.5566
R1071 B.t3 B.n204 4.95267
R1072 B.n530 B.t4 4.95267
R1073 B.n315 B.n262 4.05904
R1074 B.n295 B.n294 4.05904
R1075 B.n125 B.n124 4.05904
R1076 B.n145 B.n88 4.05904
R1077 VN.n21 VN.n12 161.3
R1078 VN.n20 VN.n19 161.3
R1079 VN.n18 VN.n13 161.3
R1080 VN.n17 VN.n16 161.3
R1081 VN.n9 VN.n0 161.3
R1082 VN.n8 VN.n7 161.3
R1083 VN.n6 VN.n1 161.3
R1084 VN.n5 VN.n4 161.3
R1085 VN.n11 VN.n10 90.2042
R1086 VN.n23 VN.n22 90.2042
R1087 VN.n2 VN.t1 77.7446
R1088 VN.n14 VN.t4 77.7446
R1089 VN.n3 VN.n2 57.6509
R1090 VN.n15 VN.n14 57.6509
R1091 VN.n8 VN.n1 56.5193
R1092 VN.n20 VN.n13 56.5193
R1093 VN.n3 VN.t5 47.2837
R1094 VN.n10 VN.t3 47.2837
R1095 VN.n15 VN.t0 47.2837
R1096 VN.n22 VN.t2 47.2837
R1097 VN VN.n23 39.6156
R1098 VN.n4 VN.n1 24.4675
R1099 VN.n9 VN.n8 24.4675
R1100 VN.n16 VN.n13 24.4675
R1101 VN.n21 VN.n20 24.4675
R1102 VN.n10 VN.n9 20.5528
R1103 VN.n22 VN.n21 20.5528
R1104 VN.n17 VN.n14 13.2264
R1105 VN.n5 VN.n2 13.2264
R1106 VN.n4 VN.n3 12.234
R1107 VN.n16 VN.n15 12.234
R1108 VN.n23 VN.n12 0.278367
R1109 VN.n11 VN.n0 0.278367
R1110 VN.n19 VN.n12 0.189894
R1111 VN.n19 VN.n18 0.189894
R1112 VN.n18 VN.n17 0.189894
R1113 VN.n6 VN.n5 0.189894
R1114 VN.n7 VN.n6 0.189894
R1115 VN.n7 VN.n0 0.189894
R1116 VN VN.n11 0.153454
R1117 VDD2.n1 VDD2.t4 84.7142
R1118 VDD2.n2 VDD2.t3 83.3665
R1119 VDD2.n1 VDD2.n0 78.2939
R1120 VDD2 VDD2.n3 78.2912
R1121 VDD2.n2 VDD2.n1 32.9071
R1122 VDD2.n3 VDD2.t5 5.48526
R1123 VDD2.n3 VDD2.t1 5.48526
R1124 VDD2.n0 VDD2.t0 5.48526
R1125 VDD2.n0 VDD2.t2 5.48526
R1126 VDD2 VDD2.n2 1.46171
C0 VP VDD1 2.3725f
C1 VN VDD1 0.154326f
C2 VDD2 VTAIL 4.32238f
C3 VDD2 VP 0.398255f
C4 VP VTAIL 2.61974f
C5 VDD2 VN 2.1308f
C6 VN VTAIL 2.60555f
C7 VN VP 4.6441f
C8 VDD2 VDD1 1.13501f
C9 VTAIL VDD1 4.27502f
C10 VDD2 B 3.865075f
C11 VDD1 B 4.145934f
C12 VTAIL B 3.745247f
C13 VN B 9.88097f
C14 VP B 8.489309f
C15 VDD2.t4 B 0.62272f
C16 VDD2.t0 B 0.062955f
C17 VDD2.t2 B 0.062955f
C18 VDD2.n0 B 0.486899f
C19 VDD2.n1 B 1.79576f
C20 VDD2.t3 B 0.617723f
C21 VDD2.n2 B 1.66585f
C22 VDD2.t5 B 0.062955f
C23 VDD2.t1 B 0.062955f
C24 VDD2.n3 B 0.486878f
C25 VN.n0 B 0.043925f
C26 VN.t3 B 0.562933f
C27 VN.n1 B 0.056531f
C28 VN.t1 B 0.715946f
C29 VN.n2 B 0.312197f
C30 VN.t5 B 0.562933f
C31 VN.n3 B 0.312539f
C32 VN.n4 B 0.046766f
C33 VN.n5 B 0.244657f
C34 VN.n6 B 0.033317f
C35 VN.n7 B 0.033317f
C36 VN.n8 B 0.040749f
C37 VN.n9 B 0.05719f
C38 VN.n10 B 0.332899f
C39 VN.n11 B 0.038894f
C40 VN.n12 B 0.043925f
C41 VN.t2 B 0.562933f
C42 VN.n13 B 0.056531f
C43 VN.t4 B 0.715946f
C44 VN.n14 B 0.312197f
C45 VN.t0 B 0.562933f
C46 VN.n15 B 0.312539f
C47 VN.n16 B 0.046766f
C48 VN.n17 B 0.244657f
C49 VN.n18 B 0.033317f
C50 VN.n19 B 0.033317f
C51 VN.n20 B 0.040749f
C52 VN.n21 B 0.05719f
C53 VN.n22 B 0.332899f
C54 VN.n23 B 1.27414f
C55 VDD1.t1 B 0.644279f
C56 VDD1.t4 B 0.643711f
C57 VDD1.t2 B 0.065077f
C58 VDD1.t0 B 0.065077f
C59 VDD1.n0 B 0.503312f
C60 VDD1.n1 B 1.9454f
C61 VDD1.t3 B 0.065077f
C62 VDD1.t5 B 0.065077f
C63 VDD1.n2 B 0.501446f
C64 VDD1.n3 B 1.73697f
C65 VTAIL.t1 B 0.082441f
C66 VTAIL.t2 B 0.082441f
C67 VTAIL.n0 B 0.576044f
C68 VTAIL.n1 B 0.422467f
C69 VTAIL.t8 B 0.741793f
C70 VTAIL.n2 B 0.606786f
C71 VTAIL.t10 B 0.082441f
C72 VTAIL.t7 B 0.082441f
C73 VTAIL.n3 B 0.576044f
C74 VTAIL.n4 B 1.44759f
C75 VTAIL.t3 B 0.082441f
C76 VTAIL.t0 B 0.082441f
C77 VTAIL.n5 B 0.576047f
C78 VTAIL.n6 B 1.44759f
C79 VTAIL.t5 B 0.741798f
C80 VTAIL.n7 B 0.606782f
C81 VTAIL.t6 B 0.082441f
C82 VTAIL.t11 B 0.082441f
C83 VTAIL.n8 B 0.576047f
C84 VTAIL.n9 B 0.547693f
C85 VTAIL.t9 B 0.741793f
C86 VTAIL.n10 B 1.33249f
C87 VTAIL.t4 B 0.741793f
C88 VTAIL.n11 B 1.28352f
C89 VP.n0 B 0.045572f
C90 VP.t5 B 0.584034f
C91 VP.n1 B 0.05865f
C92 VP.n2 B 0.034566f
C93 VP.t3 B 0.584034f
C94 VP.n3 B 0.042276f
C95 VP.n4 B 0.045572f
C96 VP.t0 B 0.584034f
C97 VP.n5 B 0.05865f
C98 VP.t4 B 0.742782f
C99 VP.n6 B 0.323899f
C100 VP.t2 B 0.584034f
C101 VP.n7 B 0.324254f
C102 VP.n8 B 0.048519f
C103 VP.n9 B 0.253827f
C104 VP.n10 B 0.034566f
C105 VP.n11 B 0.034566f
C106 VP.n12 B 0.042276f
C107 VP.n13 B 0.059333f
C108 VP.n14 B 0.345377f
C109 VP.n15 B 1.30252f
C110 VP.n16 B 1.33411f
C111 VP.t1 B 0.584034f
C112 VP.n17 B 0.345377f
C113 VP.n18 B 0.059333f
C114 VP.n19 B 0.045572f
C115 VP.n20 B 0.034566f
C116 VP.n21 B 0.034566f
C117 VP.n22 B 0.05865f
C118 VP.n23 B 0.048519f
C119 VP.n24 B 0.246288f
C120 VP.n25 B 0.048519f
C121 VP.n26 B 0.034566f
C122 VP.n27 B 0.034566f
C123 VP.n28 B 0.034566f
C124 VP.n29 B 0.042276f
C125 VP.n30 B 0.059333f
C126 VP.n31 B 0.345377f
C127 VP.n32 B 0.040352f
.ends

