* NGSPICE file created from diff_pair_sample_0030.ext - technology: sky130A

.subckt diff_pair_sample_0030 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=3.11355 ps=19.2 w=18.87 l=0.82
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=0 ps=0 w=18.87 l=0.82
X2 VDD2.t1 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.11355 pd=19.2 as=7.3593 ps=38.52 w=18.87 l=0.82
X3 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.11355 pd=19.2 as=7.3593 ps=38.52 w=18.87 l=0.82
X4 VTAIL.t5 VN.t2 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=3.11355 ps=19.2 w=18.87 l=0.82
X5 VDD1.t2 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.11355 pd=19.2 as=7.3593 ps=38.52 w=18.87 l=0.82
X6 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=3.11355 ps=19.2 w=18.87 l=0.82
X7 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=0 ps=0 w=18.87 l=0.82
X8 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=3.11355 ps=19.2 w=18.87 l=0.82
X9 VDD2.t3 VN.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.11355 pd=19.2 as=7.3593 ps=38.52 w=18.87 l=0.82
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=0 ps=0 w=18.87 l=0.82
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3593 pd=38.52 as=0 ps=0 w=18.87 l=0.82
R0 VN.n0 VN.t0 623.79
R1 VN.n1 VN.t3 623.79
R2 VN.n0 VN.t1 623.74
R3 VN.n1 VN.t2 623.74
R4 VN VN.n1 91.111
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 101.832
R7 VDD2.n2 VDD2.n1 58.8764
R8 VDD2.n1 VDD2.t0 1.04978
R9 VDD2.n1 VDD2.t3 1.04978
R10 VDD2.n0 VDD2.t2 1.04978
R11 VDD2.n0 VDD2.t1 1.04978
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n842 VTAIL.n742 289.615
R14 VTAIL.n100 VTAIL.n0 289.615
R15 VTAIL.n206 VTAIL.n106 289.615
R16 VTAIL.n312 VTAIL.n212 289.615
R17 VTAIL.n736 VTAIL.n636 289.615
R18 VTAIL.n630 VTAIL.n530 289.615
R19 VTAIL.n524 VTAIL.n424 289.615
R20 VTAIL.n418 VTAIL.n318 289.615
R21 VTAIL.n777 VTAIL.n776 185
R22 VTAIL.n774 VTAIL.n773 185
R23 VTAIL.n783 VTAIL.n782 185
R24 VTAIL.n785 VTAIL.n784 185
R25 VTAIL.n770 VTAIL.n769 185
R26 VTAIL.n791 VTAIL.n790 185
R27 VTAIL.n793 VTAIL.n792 185
R28 VTAIL.n766 VTAIL.n765 185
R29 VTAIL.n799 VTAIL.n798 185
R30 VTAIL.n801 VTAIL.n800 185
R31 VTAIL.n762 VTAIL.n761 185
R32 VTAIL.n807 VTAIL.n806 185
R33 VTAIL.n809 VTAIL.n808 185
R34 VTAIL.n758 VTAIL.n757 185
R35 VTAIL.n815 VTAIL.n814 185
R36 VTAIL.n818 VTAIL.n817 185
R37 VTAIL.n816 VTAIL.n754 185
R38 VTAIL.n823 VTAIL.n753 185
R39 VTAIL.n825 VTAIL.n824 185
R40 VTAIL.n827 VTAIL.n826 185
R41 VTAIL.n750 VTAIL.n749 185
R42 VTAIL.n833 VTAIL.n832 185
R43 VTAIL.n835 VTAIL.n834 185
R44 VTAIL.n746 VTAIL.n745 185
R45 VTAIL.n841 VTAIL.n840 185
R46 VTAIL.n843 VTAIL.n842 185
R47 VTAIL.n35 VTAIL.n34 185
R48 VTAIL.n32 VTAIL.n31 185
R49 VTAIL.n41 VTAIL.n40 185
R50 VTAIL.n43 VTAIL.n42 185
R51 VTAIL.n28 VTAIL.n27 185
R52 VTAIL.n49 VTAIL.n48 185
R53 VTAIL.n51 VTAIL.n50 185
R54 VTAIL.n24 VTAIL.n23 185
R55 VTAIL.n57 VTAIL.n56 185
R56 VTAIL.n59 VTAIL.n58 185
R57 VTAIL.n20 VTAIL.n19 185
R58 VTAIL.n65 VTAIL.n64 185
R59 VTAIL.n67 VTAIL.n66 185
R60 VTAIL.n16 VTAIL.n15 185
R61 VTAIL.n73 VTAIL.n72 185
R62 VTAIL.n76 VTAIL.n75 185
R63 VTAIL.n74 VTAIL.n12 185
R64 VTAIL.n81 VTAIL.n11 185
R65 VTAIL.n83 VTAIL.n82 185
R66 VTAIL.n85 VTAIL.n84 185
R67 VTAIL.n8 VTAIL.n7 185
R68 VTAIL.n91 VTAIL.n90 185
R69 VTAIL.n93 VTAIL.n92 185
R70 VTAIL.n4 VTAIL.n3 185
R71 VTAIL.n99 VTAIL.n98 185
R72 VTAIL.n101 VTAIL.n100 185
R73 VTAIL.n141 VTAIL.n140 185
R74 VTAIL.n138 VTAIL.n137 185
R75 VTAIL.n147 VTAIL.n146 185
R76 VTAIL.n149 VTAIL.n148 185
R77 VTAIL.n134 VTAIL.n133 185
R78 VTAIL.n155 VTAIL.n154 185
R79 VTAIL.n157 VTAIL.n156 185
R80 VTAIL.n130 VTAIL.n129 185
R81 VTAIL.n163 VTAIL.n162 185
R82 VTAIL.n165 VTAIL.n164 185
R83 VTAIL.n126 VTAIL.n125 185
R84 VTAIL.n171 VTAIL.n170 185
R85 VTAIL.n173 VTAIL.n172 185
R86 VTAIL.n122 VTAIL.n121 185
R87 VTAIL.n179 VTAIL.n178 185
R88 VTAIL.n182 VTAIL.n181 185
R89 VTAIL.n180 VTAIL.n118 185
R90 VTAIL.n187 VTAIL.n117 185
R91 VTAIL.n189 VTAIL.n188 185
R92 VTAIL.n191 VTAIL.n190 185
R93 VTAIL.n114 VTAIL.n113 185
R94 VTAIL.n197 VTAIL.n196 185
R95 VTAIL.n199 VTAIL.n198 185
R96 VTAIL.n110 VTAIL.n109 185
R97 VTAIL.n205 VTAIL.n204 185
R98 VTAIL.n207 VTAIL.n206 185
R99 VTAIL.n247 VTAIL.n246 185
R100 VTAIL.n244 VTAIL.n243 185
R101 VTAIL.n253 VTAIL.n252 185
R102 VTAIL.n255 VTAIL.n254 185
R103 VTAIL.n240 VTAIL.n239 185
R104 VTAIL.n261 VTAIL.n260 185
R105 VTAIL.n263 VTAIL.n262 185
R106 VTAIL.n236 VTAIL.n235 185
R107 VTAIL.n269 VTAIL.n268 185
R108 VTAIL.n271 VTAIL.n270 185
R109 VTAIL.n232 VTAIL.n231 185
R110 VTAIL.n277 VTAIL.n276 185
R111 VTAIL.n279 VTAIL.n278 185
R112 VTAIL.n228 VTAIL.n227 185
R113 VTAIL.n285 VTAIL.n284 185
R114 VTAIL.n288 VTAIL.n287 185
R115 VTAIL.n286 VTAIL.n224 185
R116 VTAIL.n293 VTAIL.n223 185
R117 VTAIL.n295 VTAIL.n294 185
R118 VTAIL.n297 VTAIL.n296 185
R119 VTAIL.n220 VTAIL.n219 185
R120 VTAIL.n303 VTAIL.n302 185
R121 VTAIL.n305 VTAIL.n304 185
R122 VTAIL.n216 VTAIL.n215 185
R123 VTAIL.n311 VTAIL.n310 185
R124 VTAIL.n313 VTAIL.n312 185
R125 VTAIL.n737 VTAIL.n736 185
R126 VTAIL.n735 VTAIL.n734 185
R127 VTAIL.n640 VTAIL.n639 185
R128 VTAIL.n729 VTAIL.n728 185
R129 VTAIL.n727 VTAIL.n726 185
R130 VTAIL.n644 VTAIL.n643 185
R131 VTAIL.n721 VTAIL.n720 185
R132 VTAIL.n719 VTAIL.n718 185
R133 VTAIL.n717 VTAIL.n647 185
R134 VTAIL.n651 VTAIL.n648 185
R135 VTAIL.n712 VTAIL.n711 185
R136 VTAIL.n710 VTAIL.n709 185
R137 VTAIL.n653 VTAIL.n652 185
R138 VTAIL.n704 VTAIL.n703 185
R139 VTAIL.n702 VTAIL.n701 185
R140 VTAIL.n657 VTAIL.n656 185
R141 VTAIL.n696 VTAIL.n695 185
R142 VTAIL.n694 VTAIL.n693 185
R143 VTAIL.n661 VTAIL.n660 185
R144 VTAIL.n688 VTAIL.n687 185
R145 VTAIL.n686 VTAIL.n685 185
R146 VTAIL.n665 VTAIL.n664 185
R147 VTAIL.n680 VTAIL.n679 185
R148 VTAIL.n678 VTAIL.n677 185
R149 VTAIL.n669 VTAIL.n668 185
R150 VTAIL.n672 VTAIL.n671 185
R151 VTAIL.n631 VTAIL.n630 185
R152 VTAIL.n629 VTAIL.n628 185
R153 VTAIL.n534 VTAIL.n533 185
R154 VTAIL.n623 VTAIL.n622 185
R155 VTAIL.n621 VTAIL.n620 185
R156 VTAIL.n538 VTAIL.n537 185
R157 VTAIL.n615 VTAIL.n614 185
R158 VTAIL.n613 VTAIL.n612 185
R159 VTAIL.n611 VTAIL.n541 185
R160 VTAIL.n545 VTAIL.n542 185
R161 VTAIL.n606 VTAIL.n605 185
R162 VTAIL.n604 VTAIL.n603 185
R163 VTAIL.n547 VTAIL.n546 185
R164 VTAIL.n598 VTAIL.n597 185
R165 VTAIL.n596 VTAIL.n595 185
R166 VTAIL.n551 VTAIL.n550 185
R167 VTAIL.n590 VTAIL.n589 185
R168 VTAIL.n588 VTAIL.n587 185
R169 VTAIL.n555 VTAIL.n554 185
R170 VTAIL.n582 VTAIL.n581 185
R171 VTAIL.n580 VTAIL.n579 185
R172 VTAIL.n559 VTAIL.n558 185
R173 VTAIL.n574 VTAIL.n573 185
R174 VTAIL.n572 VTAIL.n571 185
R175 VTAIL.n563 VTAIL.n562 185
R176 VTAIL.n566 VTAIL.n565 185
R177 VTAIL.n525 VTAIL.n524 185
R178 VTAIL.n523 VTAIL.n522 185
R179 VTAIL.n428 VTAIL.n427 185
R180 VTAIL.n517 VTAIL.n516 185
R181 VTAIL.n515 VTAIL.n514 185
R182 VTAIL.n432 VTAIL.n431 185
R183 VTAIL.n509 VTAIL.n508 185
R184 VTAIL.n507 VTAIL.n506 185
R185 VTAIL.n505 VTAIL.n435 185
R186 VTAIL.n439 VTAIL.n436 185
R187 VTAIL.n500 VTAIL.n499 185
R188 VTAIL.n498 VTAIL.n497 185
R189 VTAIL.n441 VTAIL.n440 185
R190 VTAIL.n492 VTAIL.n491 185
R191 VTAIL.n490 VTAIL.n489 185
R192 VTAIL.n445 VTAIL.n444 185
R193 VTAIL.n484 VTAIL.n483 185
R194 VTAIL.n482 VTAIL.n481 185
R195 VTAIL.n449 VTAIL.n448 185
R196 VTAIL.n476 VTAIL.n475 185
R197 VTAIL.n474 VTAIL.n473 185
R198 VTAIL.n453 VTAIL.n452 185
R199 VTAIL.n468 VTAIL.n467 185
R200 VTAIL.n466 VTAIL.n465 185
R201 VTAIL.n457 VTAIL.n456 185
R202 VTAIL.n460 VTAIL.n459 185
R203 VTAIL.n419 VTAIL.n418 185
R204 VTAIL.n417 VTAIL.n416 185
R205 VTAIL.n322 VTAIL.n321 185
R206 VTAIL.n411 VTAIL.n410 185
R207 VTAIL.n409 VTAIL.n408 185
R208 VTAIL.n326 VTAIL.n325 185
R209 VTAIL.n403 VTAIL.n402 185
R210 VTAIL.n401 VTAIL.n400 185
R211 VTAIL.n399 VTAIL.n329 185
R212 VTAIL.n333 VTAIL.n330 185
R213 VTAIL.n394 VTAIL.n393 185
R214 VTAIL.n392 VTAIL.n391 185
R215 VTAIL.n335 VTAIL.n334 185
R216 VTAIL.n386 VTAIL.n385 185
R217 VTAIL.n384 VTAIL.n383 185
R218 VTAIL.n339 VTAIL.n338 185
R219 VTAIL.n378 VTAIL.n377 185
R220 VTAIL.n376 VTAIL.n375 185
R221 VTAIL.n343 VTAIL.n342 185
R222 VTAIL.n370 VTAIL.n369 185
R223 VTAIL.n368 VTAIL.n367 185
R224 VTAIL.n347 VTAIL.n346 185
R225 VTAIL.n362 VTAIL.n361 185
R226 VTAIL.n360 VTAIL.n359 185
R227 VTAIL.n351 VTAIL.n350 185
R228 VTAIL.n354 VTAIL.n353 185
R229 VTAIL.t1 VTAIL.n670 147.659
R230 VTAIL.t2 VTAIL.n564 147.659
R231 VTAIL.t4 VTAIL.n458 147.659
R232 VTAIL.t5 VTAIL.n352 147.659
R233 VTAIL.t6 VTAIL.n775 147.659
R234 VTAIL.t7 VTAIL.n33 147.659
R235 VTAIL.t3 VTAIL.n139 147.659
R236 VTAIL.t0 VTAIL.n245 147.659
R237 VTAIL.n776 VTAIL.n773 104.615
R238 VTAIL.n783 VTAIL.n773 104.615
R239 VTAIL.n784 VTAIL.n783 104.615
R240 VTAIL.n784 VTAIL.n769 104.615
R241 VTAIL.n791 VTAIL.n769 104.615
R242 VTAIL.n792 VTAIL.n791 104.615
R243 VTAIL.n792 VTAIL.n765 104.615
R244 VTAIL.n799 VTAIL.n765 104.615
R245 VTAIL.n800 VTAIL.n799 104.615
R246 VTAIL.n800 VTAIL.n761 104.615
R247 VTAIL.n807 VTAIL.n761 104.615
R248 VTAIL.n808 VTAIL.n807 104.615
R249 VTAIL.n808 VTAIL.n757 104.615
R250 VTAIL.n815 VTAIL.n757 104.615
R251 VTAIL.n817 VTAIL.n815 104.615
R252 VTAIL.n817 VTAIL.n816 104.615
R253 VTAIL.n816 VTAIL.n753 104.615
R254 VTAIL.n825 VTAIL.n753 104.615
R255 VTAIL.n826 VTAIL.n825 104.615
R256 VTAIL.n826 VTAIL.n749 104.615
R257 VTAIL.n833 VTAIL.n749 104.615
R258 VTAIL.n834 VTAIL.n833 104.615
R259 VTAIL.n834 VTAIL.n745 104.615
R260 VTAIL.n841 VTAIL.n745 104.615
R261 VTAIL.n842 VTAIL.n841 104.615
R262 VTAIL.n34 VTAIL.n31 104.615
R263 VTAIL.n41 VTAIL.n31 104.615
R264 VTAIL.n42 VTAIL.n41 104.615
R265 VTAIL.n42 VTAIL.n27 104.615
R266 VTAIL.n49 VTAIL.n27 104.615
R267 VTAIL.n50 VTAIL.n49 104.615
R268 VTAIL.n50 VTAIL.n23 104.615
R269 VTAIL.n57 VTAIL.n23 104.615
R270 VTAIL.n58 VTAIL.n57 104.615
R271 VTAIL.n58 VTAIL.n19 104.615
R272 VTAIL.n65 VTAIL.n19 104.615
R273 VTAIL.n66 VTAIL.n65 104.615
R274 VTAIL.n66 VTAIL.n15 104.615
R275 VTAIL.n73 VTAIL.n15 104.615
R276 VTAIL.n75 VTAIL.n73 104.615
R277 VTAIL.n75 VTAIL.n74 104.615
R278 VTAIL.n74 VTAIL.n11 104.615
R279 VTAIL.n83 VTAIL.n11 104.615
R280 VTAIL.n84 VTAIL.n83 104.615
R281 VTAIL.n84 VTAIL.n7 104.615
R282 VTAIL.n91 VTAIL.n7 104.615
R283 VTAIL.n92 VTAIL.n91 104.615
R284 VTAIL.n92 VTAIL.n3 104.615
R285 VTAIL.n99 VTAIL.n3 104.615
R286 VTAIL.n100 VTAIL.n99 104.615
R287 VTAIL.n140 VTAIL.n137 104.615
R288 VTAIL.n147 VTAIL.n137 104.615
R289 VTAIL.n148 VTAIL.n147 104.615
R290 VTAIL.n148 VTAIL.n133 104.615
R291 VTAIL.n155 VTAIL.n133 104.615
R292 VTAIL.n156 VTAIL.n155 104.615
R293 VTAIL.n156 VTAIL.n129 104.615
R294 VTAIL.n163 VTAIL.n129 104.615
R295 VTAIL.n164 VTAIL.n163 104.615
R296 VTAIL.n164 VTAIL.n125 104.615
R297 VTAIL.n171 VTAIL.n125 104.615
R298 VTAIL.n172 VTAIL.n171 104.615
R299 VTAIL.n172 VTAIL.n121 104.615
R300 VTAIL.n179 VTAIL.n121 104.615
R301 VTAIL.n181 VTAIL.n179 104.615
R302 VTAIL.n181 VTAIL.n180 104.615
R303 VTAIL.n180 VTAIL.n117 104.615
R304 VTAIL.n189 VTAIL.n117 104.615
R305 VTAIL.n190 VTAIL.n189 104.615
R306 VTAIL.n190 VTAIL.n113 104.615
R307 VTAIL.n197 VTAIL.n113 104.615
R308 VTAIL.n198 VTAIL.n197 104.615
R309 VTAIL.n198 VTAIL.n109 104.615
R310 VTAIL.n205 VTAIL.n109 104.615
R311 VTAIL.n206 VTAIL.n205 104.615
R312 VTAIL.n246 VTAIL.n243 104.615
R313 VTAIL.n253 VTAIL.n243 104.615
R314 VTAIL.n254 VTAIL.n253 104.615
R315 VTAIL.n254 VTAIL.n239 104.615
R316 VTAIL.n261 VTAIL.n239 104.615
R317 VTAIL.n262 VTAIL.n261 104.615
R318 VTAIL.n262 VTAIL.n235 104.615
R319 VTAIL.n269 VTAIL.n235 104.615
R320 VTAIL.n270 VTAIL.n269 104.615
R321 VTAIL.n270 VTAIL.n231 104.615
R322 VTAIL.n277 VTAIL.n231 104.615
R323 VTAIL.n278 VTAIL.n277 104.615
R324 VTAIL.n278 VTAIL.n227 104.615
R325 VTAIL.n285 VTAIL.n227 104.615
R326 VTAIL.n287 VTAIL.n285 104.615
R327 VTAIL.n287 VTAIL.n286 104.615
R328 VTAIL.n286 VTAIL.n223 104.615
R329 VTAIL.n295 VTAIL.n223 104.615
R330 VTAIL.n296 VTAIL.n295 104.615
R331 VTAIL.n296 VTAIL.n219 104.615
R332 VTAIL.n303 VTAIL.n219 104.615
R333 VTAIL.n304 VTAIL.n303 104.615
R334 VTAIL.n304 VTAIL.n215 104.615
R335 VTAIL.n311 VTAIL.n215 104.615
R336 VTAIL.n312 VTAIL.n311 104.615
R337 VTAIL.n736 VTAIL.n735 104.615
R338 VTAIL.n735 VTAIL.n639 104.615
R339 VTAIL.n728 VTAIL.n639 104.615
R340 VTAIL.n728 VTAIL.n727 104.615
R341 VTAIL.n727 VTAIL.n643 104.615
R342 VTAIL.n720 VTAIL.n643 104.615
R343 VTAIL.n720 VTAIL.n719 104.615
R344 VTAIL.n719 VTAIL.n647 104.615
R345 VTAIL.n651 VTAIL.n647 104.615
R346 VTAIL.n711 VTAIL.n651 104.615
R347 VTAIL.n711 VTAIL.n710 104.615
R348 VTAIL.n710 VTAIL.n652 104.615
R349 VTAIL.n703 VTAIL.n652 104.615
R350 VTAIL.n703 VTAIL.n702 104.615
R351 VTAIL.n702 VTAIL.n656 104.615
R352 VTAIL.n695 VTAIL.n656 104.615
R353 VTAIL.n695 VTAIL.n694 104.615
R354 VTAIL.n694 VTAIL.n660 104.615
R355 VTAIL.n687 VTAIL.n660 104.615
R356 VTAIL.n687 VTAIL.n686 104.615
R357 VTAIL.n686 VTAIL.n664 104.615
R358 VTAIL.n679 VTAIL.n664 104.615
R359 VTAIL.n679 VTAIL.n678 104.615
R360 VTAIL.n678 VTAIL.n668 104.615
R361 VTAIL.n671 VTAIL.n668 104.615
R362 VTAIL.n630 VTAIL.n629 104.615
R363 VTAIL.n629 VTAIL.n533 104.615
R364 VTAIL.n622 VTAIL.n533 104.615
R365 VTAIL.n622 VTAIL.n621 104.615
R366 VTAIL.n621 VTAIL.n537 104.615
R367 VTAIL.n614 VTAIL.n537 104.615
R368 VTAIL.n614 VTAIL.n613 104.615
R369 VTAIL.n613 VTAIL.n541 104.615
R370 VTAIL.n545 VTAIL.n541 104.615
R371 VTAIL.n605 VTAIL.n545 104.615
R372 VTAIL.n605 VTAIL.n604 104.615
R373 VTAIL.n604 VTAIL.n546 104.615
R374 VTAIL.n597 VTAIL.n546 104.615
R375 VTAIL.n597 VTAIL.n596 104.615
R376 VTAIL.n596 VTAIL.n550 104.615
R377 VTAIL.n589 VTAIL.n550 104.615
R378 VTAIL.n589 VTAIL.n588 104.615
R379 VTAIL.n588 VTAIL.n554 104.615
R380 VTAIL.n581 VTAIL.n554 104.615
R381 VTAIL.n581 VTAIL.n580 104.615
R382 VTAIL.n580 VTAIL.n558 104.615
R383 VTAIL.n573 VTAIL.n558 104.615
R384 VTAIL.n573 VTAIL.n572 104.615
R385 VTAIL.n572 VTAIL.n562 104.615
R386 VTAIL.n565 VTAIL.n562 104.615
R387 VTAIL.n524 VTAIL.n523 104.615
R388 VTAIL.n523 VTAIL.n427 104.615
R389 VTAIL.n516 VTAIL.n427 104.615
R390 VTAIL.n516 VTAIL.n515 104.615
R391 VTAIL.n515 VTAIL.n431 104.615
R392 VTAIL.n508 VTAIL.n431 104.615
R393 VTAIL.n508 VTAIL.n507 104.615
R394 VTAIL.n507 VTAIL.n435 104.615
R395 VTAIL.n439 VTAIL.n435 104.615
R396 VTAIL.n499 VTAIL.n439 104.615
R397 VTAIL.n499 VTAIL.n498 104.615
R398 VTAIL.n498 VTAIL.n440 104.615
R399 VTAIL.n491 VTAIL.n440 104.615
R400 VTAIL.n491 VTAIL.n490 104.615
R401 VTAIL.n490 VTAIL.n444 104.615
R402 VTAIL.n483 VTAIL.n444 104.615
R403 VTAIL.n483 VTAIL.n482 104.615
R404 VTAIL.n482 VTAIL.n448 104.615
R405 VTAIL.n475 VTAIL.n448 104.615
R406 VTAIL.n475 VTAIL.n474 104.615
R407 VTAIL.n474 VTAIL.n452 104.615
R408 VTAIL.n467 VTAIL.n452 104.615
R409 VTAIL.n467 VTAIL.n466 104.615
R410 VTAIL.n466 VTAIL.n456 104.615
R411 VTAIL.n459 VTAIL.n456 104.615
R412 VTAIL.n418 VTAIL.n417 104.615
R413 VTAIL.n417 VTAIL.n321 104.615
R414 VTAIL.n410 VTAIL.n321 104.615
R415 VTAIL.n410 VTAIL.n409 104.615
R416 VTAIL.n409 VTAIL.n325 104.615
R417 VTAIL.n402 VTAIL.n325 104.615
R418 VTAIL.n402 VTAIL.n401 104.615
R419 VTAIL.n401 VTAIL.n329 104.615
R420 VTAIL.n333 VTAIL.n329 104.615
R421 VTAIL.n393 VTAIL.n333 104.615
R422 VTAIL.n393 VTAIL.n392 104.615
R423 VTAIL.n392 VTAIL.n334 104.615
R424 VTAIL.n385 VTAIL.n334 104.615
R425 VTAIL.n385 VTAIL.n384 104.615
R426 VTAIL.n384 VTAIL.n338 104.615
R427 VTAIL.n377 VTAIL.n338 104.615
R428 VTAIL.n377 VTAIL.n376 104.615
R429 VTAIL.n376 VTAIL.n342 104.615
R430 VTAIL.n369 VTAIL.n342 104.615
R431 VTAIL.n369 VTAIL.n368 104.615
R432 VTAIL.n368 VTAIL.n346 104.615
R433 VTAIL.n361 VTAIL.n346 104.615
R434 VTAIL.n361 VTAIL.n360 104.615
R435 VTAIL.n360 VTAIL.n350 104.615
R436 VTAIL.n353 VTAIL.n350 104.615
R437 VTAIL.n776 VTAIL.t6 52.3082
R438 VTAIL.n34 VTAIL.t7 52.3082
R439 VTAIL.n140 VTAIL.t3 52.3082
R440 VTAIL.n246 VTAIL.t0 52.3082
R441 VTAIL.n671 VTAIL.t1 52.3082
R442 VTAIL.n565 VTAIL.t2 52.3082
R443 VTAIL.n459 VTAIL.t4 52.3082
R444 VTAIL.n353 VTAIL.t5 52.3082
R445 VTAIL.n847 VTAIL.n846 30.4399
R446 VTAIL.n105 VTAIL.n104 30.4399
R447 VTAIL.n211 VTAIL.n210 30.4399
R448 VTAIL.n317 VTAIL.n316 30.4399
R449 VTAIL.n741 VTAIL.n740 30.4399
R450 VTAIL.n635 VTAIL.n634 30.4399
R451 VTAIL.n529 VTAIL.n528 30.4399
R452 VTAIL.n423 VTAIL.n422 30.4399
R453 VTAIL.n847 VTAIL.n741 29.6255
R454 VTAIL.n423 VTAIL.n317 29.6255
R455 VTAIL.n777 VTAIL.n775 15.6677
R456 VTAIL.n35 VTAIL.n33 15.6677
R457 VTAIL.n141 VTAIL.n139 15.6677
R458 VTAIL.n247 VTAIL.n245 15.6677
R459 VTAIL.n672 VTAIL.n670 15.6677
R460 VTAIL.n566 VTAIL.n564 15.6677
R461 VTAIL.n460 VTAIL.n458 15.6677
R462 VTAIL.n354 VTAIL.n352 15.6677
R463 VTAIL.n824 VTAIL.n823 13.1884
R464 VTAIL.n82 VTAIL.n81 13.1884
R465 VTAIL.n188 VTAIL.n187 13.1884
R466 VTAIL.n294 VTAIL.n293 13.1884
R467 VTAIL.n718 VTAIL.n717 13.1884
R468 VTAIL.n612 VTAIL.n611 13.1884
R469 VTAIL.n506 VTAIL.n505 13.1884
R470 VTAIL.n400 VTAIL.n399 13.1884
R471 VTAIL.n778 VTAIL.n774 12.8005
R472 VTAIL.n822 VTAIL.n754 12.8005
R473 VTAIL.n827 VTAIL.n752 12.8005
R474 VTAIL.n36 VTAIL.n32 12.8005
R475 VTAIL.n80 VTAIL.n12 12.8005
R476 VTAIL.n85 VTAIL.n10 12.8005
R477 VTAIL.n142 VTAIL.n138 12.8005
R478 VTAIL.n186 VTAIL.n118 12.8005
R479 VTAIL.n191 VTAIL.n116 12.8005
R480 VTAIL.n248 VTAIL.n244 12.8005
R481 VTAIL.n292 VTAIL.n224 12.8005
R482 VTAIL.n297 VTAIL.n222 12.8005
R483 VTAIL.n721 VTAIL.n646 12.8005
R484 VTAIL.n716 VTAIL.n648 12.8005
R485 VTAIL.n673 VTAIL.n669 12.8005
R486 VTAIL.n615 VTAIL.n540 12.8005
R487 VTAIL.n610 VTAIL.n542 12.8005
R488 VTAIL.n567 VTAIL.n563 12.8005
R489 VTAIL.n509 VTAIL.n434 12.8005
R490 VTAIL.n504 VTAIL.n436 12.8005
R491 VTAIL.n461 VTAIL.n457 12.8005
R492 VTAIL.n403 VTAIL.n328 12.8005
R493 VTAIL.n398 VTAIL.n330 12.8005
R494 VTAIL.n355 VTAIL.n351 12.8005
R495 VTAIL.n782 VTAIL.n781 12.0247
R496 VTAIL.n819 VTAIL.n818 12.0247
R497 VTAIL.n828 VTAIL.n750 12.0247
R498 VTAIL.n40 VTAIL.n39 12.0247
R499 VTAIL.n77 VTAIL.n76 12.0247
R500 VTAIL.n86 VTAIL.n8 12.0247
R501 VTAIL.n146 VTAIL.n145 12.0247
R502 VTAIL.n183 VTAIL.n182 12.0247
R503 VTAIL.n192 VTAIL.n114 12.0247
R504 VTAIL.n252 VTAIL.n251 12.0247
R505 VTAIL.n289 VTAIL.n288 12.0247
R506 VTAIL.n298 VTAIL.n220 12.0247
R507 VTAIL.n722 VTAIL.n644 12.0247
R508 VTAIL.n713 VTAIL.n712 12.0247
R509 VTAIL.n677 VTAIL.n676 12.0247
R510 VTAIL.n616 VTAIL.n538 12.0247
R511 VTAIL.n607 VTAIL.n606 12.0247
R512 VTAIL.n571 VTAIL.n570 12.0247
R513 VTAIL.n510 VTAIL.n432 12.0247
R514 VTAIL.n501 VTAIL.n500 12.0247
R515 VTAIL.n465 VTAIL.n464 12.0247
R516 VTAIL.n404 VTAIL.n326 12.0247
R517 VTAIL.n395 VTAIL.n394 12.0247
R518 VTAIL.n359 VTAIL.n358 12.0247
R519 VTAIL.n785 VTAIL.n772 11.249
R520 VTAIL.n814 VTAIL.n756 11.249
R521 VTAIL.n832 VTAIL.n831 11.249
R522 VTAIL.n43 VTAIL.n30 11.249
R523 VTAIL.n72 VTAIL.n14 11.249
R524 VTAIL.n90 VTAIL.n89 11.249
R525 VTAIL.n149 VTAIL.n136 11.249
R526 VTAIL.n178 VTAIL.n120 11.249
R527 VTAIL.n196 VTAIL.n195 11.249
R528 VTAIL.n255 VTAIL.n242 11.249
R529 VTAIL.n284 VTAIL.n226 11.249
R530 VTAIL.n302 VTAIL.n301 11.249
R531 VTAIL.n726 VTAIL.n725 11.249
R532 VTAIL.n709 VTAIL.n650 11.249
R533 VTAIL.n680 VTAIL.n667 11.249
R534 VTAIL.n620 VTAIL.n619 11.249
R535 VTAIL.n603 VTAIL.n544 11.249
R536 VTAIL.n574 VTAIL.n561 11.249
R537 VTAIL.n514 VTAIL.n513 11.249
R538 VTAIL.n497 VTAIL.n438 11.249
R539 VTAIL.n468 VTAIL.n455 11.249
R540 VTAIL.n408 VTAIL.n407 11.249
R541 VTAIL.n391 VTAIL.n332 11.249
R542 VTAIL.n362 VTAIL.n349 11.249
R543 VTAIL.n786 VTAIL.n770 10.4732
R544 VTAIL.n813 VTAIL.n758 10.4732
R545 VTAIL.n835 VTAIL.n748 10.4732
R546 VTAIL.n44 VTAIL.n28 10.4732
R547 VTAIL.n71 VTAIL.n16 10.4732
R548 VTAIL.n93 VTAIL.n6 10.4732
R549 VTAIL.n150 VTAIL.n134 10.4732
R550 VTAIL.n177 VTAIL.n122 10.4732
R551 VTAIL.n199 VTAIL.n112 10.4732
R552 VTAIL.n256 VTAIL.n240 10.4732
R553 VTAIL.n283 VTAIL.n228 10.4732
R554 VTAIL.n305 VTAIL.n218 10.4732
R555 VTAIL.n729 VTAIL.n642 10.4732
R556 VTAIL.n708 VTAIL.n653 10.4732
R557 VTAIL.n681 VTAIL.n665 10.4732
R558 VTAIL.n623 VTAIL.n536 10.4732
R559 VTAIL.n602 VTAIL.n547 10.4732
R560 VTAIL.n575 VTAIL.n559 10.4732
R561 VTAIL.n517 VTAIL.n430 10.4732
R562 VTAIL.n496 VTAIL.n441 10.4732
R563 VTAIL.n469 VTAIL.n453 10.4732
R564 VTAIL.n411 VTAIL.n324 10.4732
R565 VTAIL.n390 VTAIL.n335 10.4732
R566 VTAIL.n363 VTAIL.n347 10.4732
R567 VTAIL.n790 VTAIL.n789 9.69747
R568 VTAIL.n810 VTAIL.n809 9.69747
R569 VTAIL.n836 VTAIL.n746 9.69747
R570 VTAIL.n48 VTAIL.n47 9.69747
R571 VTAIL.n68 VTAIL.n67 9.69747
R572 VTAIL.n94 VTAIL.n4 9.69747
R573 VTAIL.n154 VTAIL.n153 9.69747
R574 VTAIL.n174 VTAIL.n173 9.69747
R575 VTAIL.n200 VTAIL.n110 9.69747
R576 VTAIL.n260 VTAIL.n259 9.69747
R577 VTAIL.n280 VTAIL.n279 9.69747
R578 VTAIL.n306 VTAIL.n216 9.69747
R579 VTAIL.n730 VTAIL.n640 9.69747
R580 VTAIL.n705 VTAIL.n704 9.69747
R581 VTAIL.n685 VTAIL.n684 9.69747
R582 VTAIL.n624 VTAIL.n534 9.69747
R583 VTAIL.n599 VTAIL.n598 9.69747
R584 VTAIL.n579 VTAIL.n578 9.69747
R585 VTAIL.n518 VTAIL.n428 9.69747
R586 VTAIL.n493 VTAIL.n492 9.69747
R587 VTAIL.n473 VTAIL.n472 9.69747
R588 VTAIL.n412 VTAIL.n322 9.69747
R589 VTAIL.n387 VTAIL.n386 9.69747
R590 VTAIL.n367 VTAIL.n366 9.69747
R591 VTAIL.n846 VTAIL.n845 9.45567
R592 VTAIL.n104 VTAIL.n103 9.45567
R593 VTAIL.n210 VTAIL.n209 9.45567
R594 VTAIL.n316 VTAIL.n315 9.45567
R595 VTAIL.n740 VTAIL.n739 9.45567
R596 VTAIL.n634 VTAIL.n633 9.45567
R597 VTAIL.n528 VTAIL.n527 9.45567
R598 VTAIL.n422 VTAIL.n421 9.45567
R599 VTAIL.n744 VTAIL.n743 9.3005
R600 VTAIL.n839 VTAIL.n838 9.3005
R601 VTAIL.n837 VTAIL.n836 9.3005
R602 VTAIL.n748 VTAIL.n747 9.3005
R603 VTAIL.n831 VTAIL.n830 9.3005
R604 VTAIL.n829 VTAIL.n828 9.3005
R605 VTAIL.n752 VTAIL.n751 9.3005
R606 VTAIL.n797 VTAIL.n796 9.3005
R607 VTAIL.n795 VTAIL.n794 9.3005
R608 VTAIL.n768 VTAIL.n767 9.3005
R609 VTAIL.n789 VTAIL.n788 9.3005
R610 VTAIL.n787 VTAIL.n786 9.3005
R611 VTAIL.n772 VTAIL.n771 9.3005
R612 VTAIL.n781 VTAIL.n780 9.3005
R613 VTAIL.n779 VTAIL.n778 9.3005
R614 VTAIL.n764 VTAIL.n763 9.3005
R615 VTAIL.n803 VTAIL.n802 9.3005
R616 VTAIL.n805 VTAIL.n804 9.3005
R617 VTAIL.n760 VTAIL.n759 9.3005
R618 VTAIL.n811 VTAIL.n810 9.3005
R619 VTAIL.n813 VTAIL.n812 9.3005
R620 VTAIL.n756 VTAIL.n755 9.3005
R621 VTAIL.n820 VTAIL.n819 9.3005
R622 VTAIL.n822 VTAIL.n821 9.3005
R623 VTAIL.n845 VTAIL.n844 9.3005
R624 VTAIL.n2 VTAIL.n1 9.3005
R625 VTAIL.n97 VTAIL.n96 9.3005
R626 VTAIL.n95 VTAIL.n94 9.3005
R627 VTAIL.n6 VTAIL.n5 9.3005
R628 VTAIL.n89 VTAIL.n88 9.3005
R629 VTAIL.n87 VTAIL.n86 9.3005
R630 VTAIL.n10 VTAIL.n9 9.3005
R631 VTAIL.n55 VTAIL.n54 9.3005
R632 VTAIL.n53 VTAIL.n52 9.3005
R633 VTAIL.n26 VTAIL.n25 9.3005
R634 VTAIL.n47 VTAIL.n46 9.3005
R635 VTAIL.n45 VTAIL.n44 9.3005
R636 VTAIL.n30 VTAIL.n29 9.3005
R637 VTAIL.n39 VTAIL.n38 9.3005
R638 VTAIL.n37 VTAIL.n36 9.3005
R639 VTAIL.n22 VTAIL.n21 9.3005
R640 VTAIL.n61 VTAIL.n60 9.3005
R641 VTAIL.n63 VTAIL.n62 9.3005
R642 VTAIL.n18 VTAIL.n17 9.3005
R643 VTAIL.n69 VTAIL.n68 9.3005
R644 VTAIL.n71 VTAIL.n70 9.3005
R645 VTAIL.n14 VTAIL.n13 9.3005
R646 VTAIL.n78 VTAIL.n77 9.3005
R647 VTAIL.n80 VTAIL.n79 9.3005
R648 VTAIL.n103 VTAIL.n102 9.3005
R649 VTAIL.n108 VTAIL.n107 9.3005
R650 VTAIL.n203 VTAIL.n202 9.3005
R651 VTAIL.n201 VTAIL.n200 9.3005
R652 VTAIL.n112 VTAIL.n111 9.3005
R653 VTAIL.n195 VTAIL.n194 9.3005
R654 VTAIL.n193 VTAIL.n192 9.3005
R655 VTAIL.n116 VTAIL.n115 9.3005
R656 VTAIL.n161 VTAIL.n160 9.3005
R657 VTAIL.n159 VTAIL.n158 9.3005
R658 VTAIL.n132 VTAIL.n131 9.3005
R659 VTAIL.n153 VTAIL.n152 9.3005
R660 VTAIL.n151 VTAIL.n150 9.3005
R661 VTAIL.n136 VTAIL.n135 9.3005
R662 VTAIL.n145 VTAIL.n144 9.3005
R663 VTAIL.n143 VTAIL.n142 9.3005
R664 VTAIL.n128 VTAIL.n127 9.3005
R665 VTAIL.n167 VTAIL.n166 9.3005
R666 VTAIL.n169 VTAIL.n168 9.3005
R667 VTAIL.n124 VTAIL.n123 9.3005
R668 VTAIL.n175 VTAIL.n174 9.3005
R669 VTAIL.n177 VTAIL.n176 9.3005
R670 VTAIL.n120 VTAIL.n119 9.3005
R671 VTAIL.n184 VTAIL.n183 9.3005
R672 VTAIL.n186 VTAIL.n185 9.3005
R673 VTAIL.n209 VTAIL.n208 9.3005
R674 VTAIL.n214 VTAIL.n213 9.3005
R675 VTAIL.n309 VTAIL.n308 9.3005
R676 VTAIL.n307 VTAIL.n306 9.3005
R677 VTAIL.n218 VTAIL.n217 9.3005
R678 VTAIL.n301 VTAIL.n300 9.3005
R679 VTAIL.n299 VTAIL.n298 9.3005
R680 VTAIL.n222 VTAIL.n221 9.3005
R681 VTAIL.n267 VTAIL.n266 9.3005
R682 VTAIL.n265 VTAIL.n264 9.3005
R683 VTAIL.n238 VTAIL.n237 9.3005
R684 VTAIL.n259 VTAIL.n258 9.3005
R685 VTAIL.n257 VTAIL.n256 9.3005
R686 VTAIL.n242 VTAIL.n241 9.3005
R687 VTAIL.n251 VTAIL.n250 9.3005
R688 VTAIL.n249 VTAIL.n248 9.3005
R689 VTAIL.n234 VTAIL.n233 9.3005
R690 VTAIL.n273 VTAIL.n272 9.3005
R691 VTAIL.n275 VTAIL.n274 9.3005
R692 VTAIL.n230 VTAIL.n229 9.3005
R693 VTAIL.n281 VTAIL.n280 9.3005
R694 VTAIL.n283 VTAIL.n282 9.3005
R695 VTAIL.n226 VTAIL.n225 9.3005
R696 VTAIL.n290 VTAIL.n289 9.3005
R697 VTAIL.n292 VTAIL.n291 9.3005
R698 VTAIL.n315 VTAIL.n314 9.3005
R699 VTAIL.n698 VTAIL.n697 9.3005
R700 VTAIL.n700 VTAIL.n699 9.3005
R701 VTAIL.n655 VTAIL.n654 9.3005
R702 VTAIL.n706 VTAIL.n705 9.3005
R703 VTAIL.n708 VTAIL.n707 9.3005
R704 VTAIL.n650 VTAIL.n649 9.3005
R705 VTAIL.n714 VTAIL.n713 9.3005
R706 VTAIL.n716 VTAIL.n715 9.3005
R707 VTAIL.n739 VTAIL.n738 9.3005
R708 VTAIL.n638 VTAIL.n637 9.3005
R709 VTAIL.n733 VTAIL.n732 9.3005
R710 VTAIL.n731 VTAIL.n730 9.3005
R711 VTAIL.n642 VTAIL.n641 9.3005
R712 VTAIL.n725 VTAIL.n724 9.3005
R713 VTAIL.n723 VTAIL.n722 9.3005
R714 VTAIL.n646 VTAIL.n645 9.3005
R715 VTAIL.n659 VTAIL.n658 9.3005
R716 VTAIL.n692 VTAIL.n691 9.3005
R717 VTAIL.n690 VTAIL.n689 9.3005
R718 VTAIL.n663 VTAIL.n662 9.3005
R719 VTAIL.n684 VTAIL.n683 9.3005
R720 VTAIL.n682 VTAIL.n681 9.3005
R721 VTAIL.n667 VTAIL.n666 9.3005
R722 VTAIL.n676 VTAIL.n675 9.3005
R723 VTAIL.n674 VTAIL.n673 9.3005
R724 VTAIL.n592 VTAIL.n591 9.3005
R725 VTAIL.n594 VTAIL.n593 9.3005
R726 VTAIL.n549 VTAIL.n548 9.3005
R727 VTAIL.n600 VTAIL.n599 9.3005
R728 VTAIL.n602 VTAIL.n601 9.3005
R729 VTAIL.n544 VTAIL.n543 9.3005
R730 VTAIL.n608 VTAIL.n607 9.3005
R731 VTAIL.n610 VTAIL.n609 9.3005
R732 VTAIL.n633 VTAIL.n632 9.3005
R733 VTAIL.n532 VTAIL.n531 9.3005
R734 VTAIL.n627 VTAIL.n626 9.3005
R735 VTAIL.n625 VTAIL.n624 9.3005
R736 VTAIL.n536 VTAIL.n535 9.3005
R737 VTAIL.n619 VTAIL.n618 9.3005
R738 VTAIL.n617 VTAIL.n616 9.3005
R739 VTAIL.n540 VTAIL.n539 9.3005
R740 VTAIL.n553 VTAIL.n552 9.3005
R741 VTAIL.n586 VTAIL.n585 9.3005
R742 VTAIL.n584 VTAIL.n583 9.3005
R743 VTAIL.n557 VTAIL.n556 9.3005
R744 VTAIL.n578 VTAIL.n577 9.3005
R745 VTAIL.n576 VTAIL.n575 9.3005
R746 VTAIL.n561 VTAIL.n560 9.3005
R747 VTAIL.n570 VTAIL.n569 9.3005
R748 VTAIL.n568 VTAIL.n567 9.3005
R749 VTAIL.n486 VTAIL.n485 9.3005
R750 VTAIL.n488 VTAIL.n487 9.3005
R751 VTAIL.n443 VTAIL.n442 9.3005
R752 VTAIL.n494 VTAIL.n493 9.3005
R753 VTAIL.n496 VTAIL.n495 9.3005
R754 VTAIL.n438 VTAIL.n437 9.3005
R755 VTAIL.n502 VTAIL.n501 9.3005
R756 VTAIL.n504 VTAIL.n503 9.3005
R757 VTAIL.n527 VTAIL.n526 9.3005
R758 VTAIL.n426 VTAIL.n425 9.3005
R759 VTAIL.n521 VTAIL.n520 9.3005
R760 VTAIL.n519 VTAIL.n518 9.3005
R761 VTAIL.n430 VTAIL.n429 9.3005
R762 VTAIL.n513 VTAIL.n512 9.3005
R763 VTAIL.n511 VTAIL.n510 9.3005
R764 VTAIL.n434 VTAIL.n433 9.3005
R765 VTAIL.n447 VTAIL.n446 9.3005
R766 VTAIL.n480 VTAIL.n479 9.3005
R767 VTAIL.n478 VTAIL.n477 9.3005
R768 VTAIL.n451 VTAIL.n450 9.3005
R769 VTAIL.n472 VTAIL.n471 9.3005
R770 VTAIL.n470 VTAIL.n469 9.3005
R771 VTAIL.n455 VTAIL.n454 9.3005
R772 VTAIL.n464 VTAIL.n463 9.3005
R773 VTAIL.n462 VTAIL.n461 9.3005
R774 VTAIL.n380 VTAIL.n379 9.3005
R775 VTAIL.n382 VTAIL.n381 9.3005
R776 VTAIL.n337 VTAIL.n336 9.3005
R777 VTAIL.n388 VTAIL.n387 9.3005
R778 VTAIL.n390 VTAIL.n389 9.3005
R779 VTAIL.n332 VTAIL.n331 9.3005
R780 VTAIL.n396 VTAIL.n395 9.3005
R781 VTAIL.n398 VTAIL.n397 9.3005
R782 VTAIL.n421 VTAIL.n420 9.3005
R783 VTAIL.n320 VTAIL.n319 9.3005
R784 VTAIL.n415 VTAIL.n414 9.3005
R785 VTAIL.n413 VTAIL.n412 9.3005
R786 VTAIL.n324 VTAIL.n323 9.3005
R787 VTAIL.n407 VTAIL.n406 9.3005
R788 VTAIL.n405 VTAIL.n404 9.3005
R789 VTAIL.n328 VTAIL.n327 9.3005
R790 VTAIL.n341 VTAIL.n340 9.3005
R791 VTAIL.n374 VTAIL.n373 9.3005
R792 VTAIL.n372 VTAIL.n371 9.3005
R793 VTAIL.n345 VTAIL.n344 9.3005
R794 VTAIL.n366 VTAIL.n365 9.3005
R795 VTAIL.n364 VTAIL.n363 9.3005
R796 VTAIL.n349 VTAIL.n348 9.3005
R797 VTAIL.n358 VTAIL.n357 9.3005
R798 VTAIL.n356 VTAIL.n355 9.3005
R799 VTAIL.n793 VTAIL.n768 8.92171
R800 VTAIL.n806 VTAIL.n760 8.92171
R801 VTAIL.n840 VTAIL.n839 8.92171
R802 VTAIL.n51 VTAIL.n26 8.92171
R803 VTAIL.n64 VTAIL.n18 8.92171
R804 VTAIL.n98 VTAIL.n97 8.92171
R805 VTAIL.n157 VTAIL.n132 8.92171
R806 VTAIL.n170 VTAIL.n124 8.92171
R807 VTAIL.n204 VTAIL.n203 8.92171
R808 VTAIL.n263 VTAIL.n238 8.92171
R809 VTAIL.n276 VTAIL.n230 8.92171
R810 VTAIL.n310 VTAIL.n309 8.92171
R811 VTAIL.n734 VTAIL.n733 8.92171
R812 VTAIL.n701 VTAIL.n655 8.92171
R813 VTAIL.n688 VTAIL.n663 8.92171
R814 VTAIL.n628 VTAIL.n627 8.92171
R815 VTAIL.n595 VTAIL.n549 8.92171
R816 VTAIL.n582 VTAIL.n557 8.92171
R817 VTAIL.n522 VTAIL.n521 8.92171
R818 VTAIL.n489 VTAIL.n443 8.92171
R819 VTAIL.n476 VTAIL.n451 8.92171
R820 VTAIL.n416 VTAIL.n415 8.92171
R821 VTAIL.n383 VTAIL.n337 8.92171
R822 VTAIL.n370 VTAIL.n345 8.92171
R823 VTAIL.n794 VTAIL.n766 8.14595
R824 VTAIL.n805 VTAIL.n762 8.14595
R825 VTAIL.n843 VTAIL.n744 8.14595
R826 VTAIL.n52 VTAIL.n24 8.14595
R827 VTAIL.n63 VTAIL.n20 8.14595
R828 VTAIL.n101 VTAIL.n2 8.14595
R829 VTAIL.n158 VTAIL.n130 8.14595
R830 VTAIL.n169 VTAIL.n126 8.14595
R831 VTAIL.n207 VTAIL.n108 8.14595
R832 VTAIL.n264 VTAIL.n236 8.14595
R833 VTAIL.n275 VTAIL.n232 8.14595
R834 VTAIL.n313 VTAIL.n214 8.14595
R835 VTAIL.n737 VTAIL.n638 8.14595
R836 VTAIL.n700 VTAIL.n657 8.14595
R837 VTAIL.n689 VTAIL.n661 8.14595
R838 VTAIL.n631 VTAIL.n532 8.14595
R839 VTAIL.n594 VTAIL.n551 8.14595
R840 VTAIL.n583 VTAIL.n555 8.14595
R841 VTAIL.n525 VTAIL.n426 8.14595
R842 VTAIL.n488 VTAIL.n445 8.14595
R843 VTAIL.n477 VTAIL.n449 8.14595
R844 VTAIL.n419 VTAIL.n320 8.14595
R845 VTAIL.n382 VTAIL.n339 8.14595
R846 VTAIL.n371 VTAIL.n343 8.14595
R847 VTAIL.n798 VTAIL.n797 7.3702
R848 VTAIL.n802 VTAIL.n801 7.3702
R849 VTAIL.n844 VTAIL.n742 7.3702
R850 VTAIL.n56 VTAIL.n55 7.3702
R851 VTAIL.n60 VTAIL.n59 7.3702
R852 VTAIL.n102 VTAIL.n0 7.3702
R853 VTAIL.n162 VTAIL.n161 7.3702
R854 VTAIL.n166 VTAIL.n165 7.3702
R855 VTAIL.n208 VTAIL.n106 7.3702
R856 VTAIL.n268 VTAIL.n267 7.3702
R857 VTAIL.n272 VTAIL.n271 7.3702
R858 VTAIL.n314 VTAIL.n212 7.3702
R859 VTAIL.n738 VTAIL.n636 7.3702
R860 VTAIL.n697 VTAIL.n696 7.3702
R861 VTAIL.n693 VTAIL.n692 7.3702
R862 VTAIL.n632 VTAIL.n530 7.3702
R863 VTAIL.n591 VTAIL.n590 7.3702
R864 VTAIL.n587 VTAIL.n586 7.3702
R865 VTAIL.n526 VTAIL.n424 7.3702
R866 VTAIL.n485 VTAIL.n484 7.3702
R867 VTAIL.n481 VTAIL.n480 7.3702
R868 VTAIL.n420 VTAIL.n318 7.3702
R869 VTAIL.n379 VTAIL.n378 7.3702
R870 VTAIL.n375 VTAIL.n374 7.3702
R871 VTAIL.n798 VTAIL.n764 6.59444
R872 VTAIL.n801 VTAIL.n764 6.59444
R873 VTAIL.n846 VTAIL.n742 6.59444
R874 VTAIL.n56 VTAIL.n22 6.59444
R875 VTAIL.n59 VTAIL.n22 6.59444
R876 VTAIL.n104 VTAIL.n0 6.59444
R877 VTAIL.n162 VTAIL.n128 6.59444
R878 VTAIL.n165 VTAIL.n128 6.59444
R879 VTAIL.n210 VTAIL.n106 6.59444
R880 VTAIL.n268 VTAIL.n234 6.59444
R881 VTAIL.n271 VTAIL.n234 6.59444
R882 VTAIL.n316 VTAIL.n212 6.59444
R883 VTAIL.n740 VTAIL.n636 6.59444
R884 VTAIL.n696 VTAIL.n659 6.59444
R885 VTAIL.n693 VTAIL.n659 6.59444
R886 VTAIL.n634 VTAIL.n530 6.59444
R887 VTAIL.n590 VTAIL.n553 6.59444
R888 VTAIL.n587 VTAIL.n553 6.59444
R889 VTAIL.n528 VTAIL.n424 6.59444
R890 VTAIL.n484 VTAIL.n447 6.59444
R891 VTAIL.n481 VTAIL.n447 6.59444
R892 VTAIL.n422 VTAIL.n318 6.59444
R893 VTAIL.n378 VTAIL.n341 6.59444
R894 VTAIL.n375 VTAIL.n341 6.59444
R895 VTAIL.n797 VTAIL.n766 5.81868
R896 VTAIL.n802 VTAIL.n762 5.81868
R897 VTAIL.n844 VTAIL.n843 5.81868
R898 VTAIL.n55 VTAIL.n24 5.81868
R899 VTAIL.n60 VTAIL.n20 5.81868
R900 VTAIL.n102 VTAIL.n101 5.81868
R901 VTAIL.n161 VTAIL.n130 5.81868
R902 VTAIL.n166 VTAIL.n126 5.81868
R903 VTAIL.n208 VTAIL.n207 5.81868
R904 VTAIL.n267 VTAIL.n236 5.81868
R905 VTAIL.n272 VTAIL.n232 5.81868
R906 VTAIL.n314 VTAIL.n313 5.81868
R907 VTAIL.n738 VTAIL.n737 5.81868
R908 VTAIL.n697 VTAIL.n657 5.81868
R909 VTAIL.n692 VTAIL.n661 5.81868
R910 VTAIL.n632 VTAIL.n631 5.81868
R911 VTAIL.n591 VTAIL.n551 5.81868
R912 VTAIL.n586 VTAIL.n555 5.81868
R913 VTAIL.n526 VTAIL.n525 5.81868
R914 VTAIL.n485 VTAIL.n445 5.81868
R915 VTAIL.n480 VTAIL.n449 5.81868
R916 VTAIL.n420 VTAIL.n419 5.81868
R917 VTAIL.n379 VTAIL.n339 5.81868
R918 VTAIL.n374 VTAIL.n343 5.81868
R919 VTAIL.n794 VTAIL.n793 5.04292
R920 VTAIL.n806 VTAIL.n805 5.04292
R921 VTAIL.n840 VTAIL.n744 5.04292
R922 VTAIL.n52 VTAIL.n51 5.04292
R923 VTAIL.n64 VTAIL.n63 5.04292
R924 VTAIL.n98 VTAIL.n2 5.04292
R925 VTAIL.n158 VTAIL.n157 5.04292
R926 VTAIL.n170 VTAIL.n169 5.04292
R927 VTAIL.n204 VTAIL.n108 5.04292
R928 VTAIL.n264 VTAIL.n263 5.04292
R929 VTAIL.n276 VTAIL.n275 5.04292
R930 VTAIL.n310 VTAIL.n214 5.04292
R931 VTAIL.n734 VTAIL.n638 5.04292
R932 VTAIL.n701 VTAIL.n700 5.04292
R933 VTAIL.n689 VTAIL.n688 5.04292
R934 VTAIL.n628 VTAIL.n532 5.04292
R935 VTAIL.n595 VTAIL.n594 5.04292
R936 VTAIL.n583 VTAIL.n582 5.04292
R937 VTAIL.n522 VTAIL.n426 5.04292
R938 VTAIL.n489 VTAIL.n488 5.04292
R939 VTAIL.n477 VTAIL.n476 5.04292
R940 VTAIL.n416 VTAIL.n320 5.04292
R941 VTAIL.n383 VTAIL.n382 5.04292
R942 VTAIL.n371 VTAIL.n370 5.04292
R943 VTAIL.n674 VTAIL.n670 4.38563
R944 VTAIL.n568 VTAIL.n564 4.38563
R945 VTAIL.n462 VTAIL.n458 4.38563
R946 VTAIL.n356 VTAIL.n352 4.38563
R947 VTAIL.n779 VTAIL.n775 4.38563
R948 VTAIL.n37 VTAIL.n33 4.38563
R949 VTAIL.n143 VTAIL.n139 4.38563
R950 VTAIL.n249 VTAIL.n245 4.38563
R951 VTAIL.n790 VTAIL.n768 4.26717
R952 VTAIL.n809 VTAIL.n760 4.26717
R953 VTAIL.n839 VTAIL.n746 4.26717
R954 VTAIL.n48 VTAIL.n26 4.26717
R955 VTAIL.n67 VTAIL.n18 4.26717
R956 VTAIL.n97 VTAIL.n4 4.26717
R957 VTAIL.n154 VTAIL.n132 4.26717
R958 VTAIL.n173 VTAIL.n124 4.26717
R959 VTAIL.n203 VTAIL.n110 4.26717
R960 VTAIL.n260 VTAIL.n238 4.26717
R961 VTAIL.n279 VTAIL.n230 4.26717
R962 VTAIL.n309 VTAIL.n216 4.26717
R963 VTAIL.n733 VTAIL.n640 4.26717
R964 VTAIL.n704 VTAIL.n655 4.26717
R965 VTAIL.n685 VTAIL.n663 4.26717
R966 VTAIL.n627 VTAIL.n534 4.26717
R967 VTAIL.n598 VTAIL.n549 4.26717
R968 VTAIL.n579 VTAIL.n557 4.26717
R969 VTAIL.n521 VTAIL.n428 4.26717
R970 VTAIL.n492 VTAIL.n443 4.26717
R971 VTAIL.n473 VTAIL.n451 4.26717
R972 VTAIL.n415 VTAIL.n322 4.26717
R973 VTAIL.n386 VTAIL.n337 4.26717
R974 VTAIL.n367 VTAIL.n345 4.26717
R975 VTAIL.n789 VTAIL.n770 3.49141
R976 VTAIL.n810 VTAIL.n758 3.49141
R977 VTAIL.n836 VTAIL.n835 3.49141
R978 VTAIL.n47 VTAIL.n28 3.49141
R979 VTAIL.n68 VTAIL.n16 3.49141
R980 VTAIL.n94 VTAIL.n93 3.49141
R981 VTAIL.n153 VTAIL.n134 3.49141
R982 VTAIL.n174 VTAIL.n122 3.49141
R983 VTAIL.n200 VTAIL.n199 3.49141
R984 VTAIL.n259 VTAIL.n240 3.49141
R985 VTAIL.n280 VTAIL.n228 3.49141
R986 VTAIL.n306 VTAIL.n305 3.49141
R987 VTAIL.n730 VTAIL.n729 3.49141
R988 VTAIL.n705 VTAIL.n653 3.49141
R989 VTAIL.n684 VTAIL.n665 3.49141
R990 VTAIL.n624 VTAIL.n623 3.49141
R991 VTAIL.n599 VTAIL.n547 3.49141
R992 VTAIL.n578 VTAIL.n559 3.49141
R993 VTAIL.n518 VTAIL.n517 3.49141
R994 VTAIL.n493 VTAIL.n441 3.49141
R995 VTAIL.n472 VTAIL.n453 3.49141
R996 VTAIL.n412 VTAIL.n411 3.49141
R997 VTAIL.n387 VTAIL.n335 3.49141
R998 VTAIL.n366 VTAIL.n347 3.49141
R999 VTAIL.n786 VTAIL.n785 2.71565
R1000 VTAIL.n814 VTAIL.n813 2.71565
R1001 VTAIL.n832 VTAIL.n748 2.71565
R1002 VTAIL.n44 VTAIL.n43 2.71565
R1003 VTAIL.n72 VTAIL.n71 2.71565
R1004 VTAIL.n90 VTAIL.n6 2.71565
R1005 VTAIL.n150 VTAIL.n149 2.71565
R1006 VTAIL.n178 VTAIL.n177 2.71565
R1007 VTAIL.n196 VTAIL.n112 2.71565
R1008 VTAIL.n256 VTAIL.n255 2.71565
R1009 VTAIL.n284 VTAIL.n283 2.71565
R1010 VTAIL.n302 VTAIL.n218 2.71565
R1011 VTAIL.n726 VTAIL.n642 2.71565
R1012 VTAIL.n709 VTAIL.n708 2.71565
R1013 VTAIL.n681 VTAIL.n680 2.71565
R1014 VTAIL.n620 VTAIL.n536 2.71565
R1015 VTAIL.n603 VTAIL.n602 2.71565
R1016 VTAIL.n575 VTAIL.n574 2.71565
R1017 VTAIL.n514 VTAIL.n430 2.71565
R1018 VTAIL.n497 VTAIL.n496 2.71565
R1019 VTAIL.n469 VTAIL.n468 2.71565
R1020 VTAIL.n408 VTAIL.n324 2.71565
R1021 VTAIL.n391 VTAIL.n390 2.71565
R1022 VTAIL.n363 VTAIL.n362 2.71565
R1023 VTAIL.n782 VTAIL.n772 1.93989
R1024 VTAIL.n818 VTAIL.n756 1.93989
R1025 VTAIL.n831 VTAIL.n750 1.93989
R1026 VTAIL.n40 VTAIL.n30 1.93989
R1027 VTAIL.n76 VTAIL.n14 1.93989
R1028 VTAIL.n89 VTAIL.n8 1.93989
R1029 VTAIL.n146 VTAIL.n136 1.93989
R1030 VTAIL.n182 VTAIL.n120 1.93989
R1031 VTAIL.n195 VTAIL.n114 1.93989
R1032 VTAIL.n252 VTAIL.n242 1.93989
R1033 VTAIL.n288 VTAIL.n226 1.93989
R1034 VTAIL.n301 VTAIL.n220 1.93989
R1035 VTAIL.n725 VTAIL.n644 1.93989
R1036 VTAIL.n712 VTAIL.n650 1.93989
R1037 VTAIL.n677 VTAIL.n667 1.93989
R1038 VTAIL.n619 VTAIL.n538 1.93989
R1039 VTAIL.n606 VTAIL.n544 1.93989
R1040 VTAIL.n571 VTAIL.n561 1.93989
R1041 VTAIL.n513 VTAIL.n432 1.93989
R1042 VTAIL.n500 VTAIL.n438 1.93989
R1043 VTAIL.n465 VTAIL.n455 1.93989
R1044 VTAIL.n407 VTAIL.n326 1.93989
R1045 VTAIL.n394 VTAIL.n332 1.93989
R1046 VTAIL.n359 VTAIL.n349 1.93989
R1047 VTAIL.n781 VTAIL.n774 1.16414
R1048 VTAIL.n819 VTAIL.n754 1.16414
R1049 VTAIL.n828 VTAIL.n827 1.16414
R1050 VTAIL.n39 VTAIL.n32 1.16414
R1051 VTAIL.n77 VTAIL.n12 1.16414
R1052 VTAIL.n86 VTAIL.n85 1.16414
R1053 VTAIL.n145 VTAIL.n138 1.16414
R1054 VTAIL.n183 VTAIL.n118 1.16414
R1055 VTAIL.n192 VTAIL.n191 1.16414
R1056 VTAIL.n251 VTAIL.n244 1.16414
R1057 VTAIL.n289 VTAIL.n224 1.16414
R1058 VTAIL.n298 VTAIL.n297 1.16414
R1059 VTAIL.n722 VTAIL.n721 1.16414
R1060 VTAIL.n713 VTAIL.n648 1.16414
R1061 VTAIL.n676 VTAIL.n669 1.16414
R1062 VTAIL.n616 VTAIL.n615 1.16414
R1063 VTAIL.n607 VTAIL.n542 1.16414
R1064 VTAIL.n570 VTAIL.n563 1.16414
R1065 VTAIL.n510 VTAIL.n509 1.16414
R1066 VTAIL.n501 VTAIL.n436 1.16414
R1067 VTAIL.n464 VTAIL.n457 1.16414
R1068 VTAIL.n404 VTAIL.n403 1.16414
R1069 VTAIL.n395 VTAIL.n330 1.16414
R1070 VTAIL.n358 VTAIL.n351 1.16414
R1071 VTAIL.n529 VTAIL.n423 0.991879
R1072 VTAIL.n741 VTAIL.n635 0.991879
R1073 VTAIL.n317 VTAIL.n211 0.991879
R1074 VTAIL VTAIL.n105 0.554379
R1075 VTAIL.n635 VTAIL.n529 0.470328
R1076 VTAIL.n211 VTAIL.n105 0.470328
R1077 VTAIL VTAIL.n847 0.438
R1078 VTAIL.n778 VTAIL.n777 0.388379
R1079 VTAIL.n823 VTAIL.n822 0.388379
R1080 VTAIL.n824 VTAIL.n752 0.388379
R1081 VTAIL.n36 VTAIL.n35 0.388379
R1082 VTAIL.n81 VTAIL.n80 0.388379
R1083 VTAIL.n82 VTAIL.n10 0.388379
R1084 VTAIL.n142 VTAIL.n141 0.388379
R1085 VTAIL.n187 VTAIL.n186 0.388379
R1086 VTAIL.n188 VTAIL.n116 0.388379
R1087 VTAIL.n248 VTAIL.n247 0.388379
R1088 VTAIL.n293 VTAIL.n292 0.388379
R1089 VTAIL.n294 VTAIL.n222 0.388379
R1090 VTAIL.n718 VTAIL.n646 0.388379
R1091 VTAIL.n717 VTAIL.n716 0.388379
R1092 VTAIL.n673 VTAIL.n672 0.388379
R1093 VTAIL.n612 VTAIL.n540 0.388379
R1094 VTAIL.n611 VTAIL.n610 0.388379
R1095 VTAIL.n567 VTAIL.n566 0.388379
R1096 VTAIL.n506 VTAIL.n434 0.388379
R1097 VTAIL.n505 VTAIL.n504 0.388379
R1098 VTAIL.n461 VTAIL.n460 0.388379
R1099 VTAIL.n400 VTAIL.n328 0.388379
R1100 VTAIL.n399 VTAIL.n398 0.388379
R1101 VTAIL.n355 VTAIL.n354 0.388379
R1102 VTAIL.n780 VTAIL.n779 0.155672
R1103 VTAIL.n780 VTAIL.n771 0.155672
R1104 VTAIL.n787 VTAIL.n771 0.155672
R1105 VTAIL.n788 VTAIL.n787 0.155672
R1106 VTAIL.n788 VTAIL.n767 0.155672
R1107 VTAIL.n795 VTAIL.n767 0.155672
R1108 VTAIL.n796 VTAIL.n795 0.155672
R1109 VTAIL.n796 VTAIL.n763 0.155672
R1110 VTAIL.n803 VTAIL.n763 0.155672
R1111 VTAIL.n804 VTAIL.n803 0.155672
R1112 VTAIL.n804 VTAIL.n759 0.155672
R1113 VTAIL.n811 VTAIL.n759 0.155672
R1114 VTAIL.n812 VTAIL.n811 0.155672
R1115 VTAIL.n812 VTAIL.n755 0.155672
R1116 VTAIL.n820 VTAIL.n755 0.155672
R1117 VTAIL.n821 VTAIL.n820 0.155672
R1118 VTAIL.n821 VTAIL.n751 0.155672
R1119 VTAIL.n829 VTAIL.n751 0.155672
R1120 VTAIL.n830 VTAIL.n829 0.155672
R1121 VTAIL.n830 VTAIL.n747 0.155672
R1122 VTAIL.n837 VTAIL.n747 0.155672
R1123 VTAIL.n838 VTAIL.n837 0.155672
R1124 VTAIL.n838 VTAIL.n743 0.155672
R1125 VTAIL.n845 VTAIL.n743 0.155672
R1126 VTAIL.n38 VTAIL.n37 0.155672
R1127 VTAIL.n38 VTAIL.n29 0.155672
R1128 VTAIL.n45 VTAIL.n29 0.155672
R1129 VTAIL.n46 VTAIL.n45 0.155672
R1130 VTAIL.n46 VTAIL.n25 0.155672
R1131 VTAIL.n53 VTAIL.n25 0.155672
R1132 VTAIL.n54 VTAIL.n53 0.155672
R1133 VTAIL.n54 VTAIL.n21 0.155672
R1134 VTAIL.n61 VTAIL.n21 0.155672
R1135 VTAIL.n62 VTAIL.n61 0.155672
R1136 VTAIL.n62 VTAIL.n17 0.155672
R1137 VTAIL.n69 VTAIL.n17 0.155672
R1138 VTAIL.n70 VTAIL.n69 0.155672
R1139 VTAIL.n70 VTAIL.n13 0.155672
R1140 VTAIL.n78 VTAIL.n13 0.155672
R1141 VTAIL.n79 VTAIL.n78 0.155672
R1142 VTAIL.n79 VTAIL.n9 0.155672
R1143 VTAIL.n87 VTAIL.n9 0.155672
R1144 VTAIL.n88 VTAIL.n87 0.155672
R1145 VTAIL.n88 VTAIL.n5 0.155672
R1146 VTAIL.n95 VTAIL.n5 0.155672
R1147 VTAIL.n96 VTAIL.n95 0.155672
R1148 VTAIL.n96 VTAIL.n1 0.155672
R1149 VTAIL.n103 VTAIL.n1 0.155672
R1150 VTAIL.n144 VTAIL.n143 0.155672
R1151 VTAIL.n144 VTAIL.n135 0.155672
R1152 VTAIL.n151 VTAIL.n135 0.155672
R1153 VTAIL.n152 VTAIL.n151 0.155672
R1154 VTAIL.n152 VTAIL.n131 0.155672
R1155 VTAIL.n159 VTAIL.n131 0.155672
R1156 VTAIL.n160 VTAIL.n159 0.155672
R1157 VTAIL.n160 VTAIL.n127 0.155672
R1158 VTAIL.n167 VTAIL.n127 0.155672
R1159 VTAIL.n168 VTAIL.n167 0.155672
R1160 VTAIL.n168 VTAIL.n123 0.155672
R1161 VTAIL.n175 VTAIL.n123 0.155672
R1162 VTAIL.n176 VTAIL.n175 0.155672
R1163 VTAIL.n176 VTAIL.n119 0.155672
R1164 VTAIL.n184 VTAIL.n119 0.155672
R1165 VTAIL.n185 VTAIL.n184 0.155672
R1166 VTAIL.n185 VTAIL.n115 0.155672
R1167 VTAIL.n193 VTAIL.n115 0.155672
R1168 VTAIL.n194 VTAIL.n193 0.155672
R1169 VTAIL.n194 VTAIL.n111 0.155672
R1170 VTAIL.n201 VTAIL.n111 0.155672
R1171 VTAIL.n202 VTAIL.n201 0.155672
R1172 VTAIL.n202 VTAIL.n107 0.155672
R1173 VTAIL.n209 VTAIL.n107 0.155672
R1174 VTAIL.n250 VTAIL.n249 0.155672
R1175 VTAIL.n250 VTAIL.n241 0.155672
R1176 VTAIL.n257 VTAIL.n241 0.155672
R1177 VTAIL.n258 VTAIL.n257 0.155672
R1178 VTAIL.n258 VTAIL.n237 0.155672
R1179 VTAIL.n265 VTAIL.n237 0.155672
R1180 VTAIL.n266 VTAIL.n265 0.155672
R1181 VTAIL.n266 VTAIL.n233 0.155672
R1182 VTAIL.n273 VTAIL.n233 0.155672
R1183 VTAIL.n274 VTAIL.n273 0.155672
R1184 VTAIL.n274 VTAIL.n229 0.155672
R1185 VTAIL.n281 VTAIL.n229 0.155672
R1186 VTAIL.n282 VTAIL.n281 0.155672
R1187 VTAIL.n282 VTAIL.n225 0.155672
R1188 VTAIL.n290 VTAIL.n225 0.155672
R1189 VTAIL.n291 VTAIL.n290 0.155672
R1190 VTAIL.n291 VTAIL.n221 0.155672
R1191 VTAIL.n299 VTAIL.n221 0.155672
R1192 VTAIL.n300 VTAIL.n299 0.155672
R1193 VTAIL.n300 VTAIL.n217 0.155672
R1194 VTAIL.n307 VTAIL.n217 0.155672
R1195 VTAIL.n308 VTAIL.n307 0.155672
R1196 VTAIL.n308 VTAIL.n213 0.155672
R1197 VTAIL.n315 VTAIL.n213 0.155672
R1198 VTAIL.n739 VTAIL.n637 0.155672
R1199 VTAIL.n732 VTAIL.n637 0.155672
R1200 VTAIL.n732 VTAIL.n731 0.155672
R1201 VTAIL.n731 VTAIL.n641 0.155672
R1202 VTAIL.n724 VTAIL.n641 0.155672
R1203 VTAIL.n724 VTAIL.n723 0.155672
R1204 VTAIL.n723 VTAIL.n645 0.155672
R1205 VTAIL.n715 VTAIL.n645 0.155672
R1206 VTAIL.n715 VTAIL.n714 0.155672
R1207 VTAIL.n714 VTAIL.n649 0.155672
R1208 VTAIL.n707 VTAIL.n649 0.155672
R1209 VTAIL.n707 VTAIL.n706 0.155672
R1210 VTAIL.n706 VTAIL.n654 0.155672
R1211 VTAIL.n699 VTAIL.n654 0.155672
R1212 VTAIL.n699 VTAIL.n698 0.155672
R1213 VTAIL.n698 VTAIL.n658 0.155672
R1214 VTAIL.n691 VTAIL.n658 0.155672
R1215 VTAIL.n691 VTAIL.n690 0.155672
R1216 VTAIL.n690 VTAIL.n662 0.155672
R1217 VTAIL.n683 VTAIL.n662 0.155672
R1218 VTAIL.n683 VTAIL.n682 0.155672
R1219 VTAIL.n682 VTAIL.n666 0.155672
R1220 VTAIL.n675 VTAIL.n666 0.155672
R1221 VTAIL.n675 VTAIL.n674 0.155672
R1222 VTAIL.n633 VTAIL.n531 0.155672
R1223 VTAIL.n626 VTAIL.n531 0.155672
R1224 VTAIL.n626 VTAIL.n625 0.155672
R1225 VTAIL.n625 VTAIL.n535 0.155672
R1226 VTAIL.n618 VTAIL.n535 0.155672
R1227 VTAIL.n618 VTAIL.n617 0.155672
R1228 VTAIL.n617 VTAIL.n539 0.155672
R1229 VTAIL.n609 VTAIL.n539 0.155672
R1230 VTAIL.n609 VTAIL.n608 0.155672
R1231 VTAIL.n608 VTAIL.n543 0.155672
R1232 VTAIL.n601 VTAIL.n543 0.155672
R1233 VTAIL.n601 VTAIL.n600 0.155672
R1234 VTAIL.n600 VTAIL.n548 0.155672
R1235 VTAIL.n593 VTAIL.n548 0.155672
R1236 VTAIL.n593 VTAIL.n592 0.155672
R1237 VTAIL.n592 VTAIL.n552 0.155672
R1238 VTAIL.n585 VTAIL.n552 0.155672
R1239 VTAIL.n585 VTAIL.n584 0.155672
R1240 VTAIL.n584 VTAIL.n556 0.155672
R1241 VTAIL.n577 VTAIL.n556 0.155672
R1242 VTAIL.n577 VTAIL.n576 0.155672
R1243 VTAIL.n576 VTAIL.n560 0.155672
R1244 VTAIL.n569 VTAIL.n560 0.155672
R1245 VTAIL.n569 VTAIL.n568 0.155672
R1246 VTAIL.n527 VTAIL.n425 0.155672
R1247 VTAIL.n520 VTAIL.n425 0.155672
R1248 VTAIL.n520 VTAIL.n519 0.155672
R1249 VTAIL.n519 VTAIL.n429 0.155672
R1250 VTAIL.n512 VTAIL.n429 0.155672
R1251 VTAIL.n512 VTAIL.n511 0.155672
R1252 VTAIL.n511 VTAIL.n433 0.155672
R1253 VTAIL.n503 VTAIL.n433 0.155672
R1254 VTAIL.n503 VTAIL.n502 0.155672
R1255 VTAIL.n502 VTAIL.n437 0.155672
R1256 VTAIL.n495 VTAIL.n437 0.155672
R1257 VTAIL.n495 VTAIL.n494 0.155672
R1258 VTAIL.n494 VTAIL.n442 0.155672
R1259 VTAIL.n487 VTAIL.n442 0.155672
R1260 VTAIL.n487 VTAIL.n486 0.155672
R1261 VTAIL.n486 VTAIL.n446 0.155672
R1262 VTAIL.n479 VTAIL.n446 0.155672
R1263 VTAIL.n479 VTAIL.n478 0.155672
R1264 VTAIL.n478 VTAIL.n450 0.155672
R1265 VTAIL.n471 VTAIL.n450 0.155672
R1266 VTAIL.n471 VTAIL.n470 0.155672
R1267 VTAIL.n470 VTAIL.n454 0.155672
R1268 VTAIL.n463 VTAIL.n454 0.155672
R1269 VTAIL.n463 VTAIL.n462 0.155672
R1270 VTAIL.n421 VTAIL.n319 0.155672
R1271 VTAIL.n414 VTAIL.n319 0.155672
R1272 VTAIL.n414 VTAIL.n413 0.155672
R1273 VTAIL.n413 VTAIL.n323 0.155672
R1274 VTAIL.n406 VTAIL.n323 0.155672
R1275 VTAIL.n406 VTAIL.n405 0.155672
R1276 VTAIL.n405 VTAIL.n327 0.155672
R1277 VTAIL.n397 VTAIL.n327 0.155672
R1278 VTAIL.n397 VTAIL.n396 0.155672
R1279 VTAIL.n396 VTAIL.n331 0.155672
R1280 VTAIL.n389 VTAIL.n331 0.155672
R1281 VTAIL.n389 VTAIL.n388 0.155672
R1282 VTAIL.n388 VTAIL.n336 0.155672
R1283 VTAIL.n381 VTAIL.n336 0.155672
R1284 VTAIL.n381 VTAIL.n380 0.155672
R1285 VTAIL.n380 VTAIL.n340 0.155672
R1286 VTAIL.n373 VTAIL.n340 0.155672
R1287 VTAIL.n373 VTAIL.n372 0.155672
R1288 VTAIL.n372 VTAIL.n344 0.155672
R1289 VTAIL.n365 VTAIL.n344 0.155672
R1290 VTAIL.n365 VTAIL.n364 0.155672
R1291 VTAIL.n364 VTAIL.n348 0.155672
R1292 VTAIL.n357 VTAIL.n348 0.155672
R1293 VTAIL.n357 VTAIL.n356 0.155672
R1294 B.n182 B.t8 756.255
R1295 B.n175 B.t4 756.255
R1296 B.n68 B.t11 756.255
R1297 B.n76 B.t15 756.255
R1298 B.n558 B.n557 585
R1299 B.n558 B.n36 585
R1300 B.n561 B.n560 585
R1301 B.n562 B.n107 585
R1302 B.n564 B.n563 585
R1303 B.n566 B.n106 585
R1304 B.n569 B.n568 585
R1305 B.n570 B.n105 585
R1306 B.n572 B.n571 585
R1307 B.n574 B.n104 585
R1308 B.n577 B.n576 585
R1309 B.n578 B.n103 585
R1310 B.n580 B.n579 585
R1311 B.n582 B.n102 585
R1312 B.n585 B.n584 585
R1313 B.n586 B.n101 585
R1314 B.n588 B.n587 585
R1315 B.n590 B.n100 585
R1316 B.n593 B.n592 585
R1317 B.n594 B.n99 585
R1318 B.n596 B.n595 585
R1319 B.n598 B.n98 585
R1320 B.n601 B.n600 585
R1321 B.n602 B.n97 585
R1322 B.n604 B.n603 585
R1323 B.n606 B.n96 585
R1324 B.n609 B.n608 585
R1325 B.n610 B.n95 585
R1326 B.n612 B.n611 585
R1327 B.n614 B.n94 585
R1328 B.n617 B.n616 585
R1329 B.n618 B.n93 585
R1330 B.n620 B.n619 585
R1331 B.n622 B.n92 585
R1332 B.n625 B.n624 585
R1333 B.n626 B.n91 585
R1334 B.n628 B.n627 585
R1335 B.n630 B.n90 585
R1336 B.n633 B.n632 585
R1337 B.n634 B.n89 585
R1338 B.n636 B.n635 585
R1339 B.n638 B.n88 585
R1340 B.n641 B.n640 585
R1341 B.n642 B.n87 585
R1342 B.n644 B.n643 585
R1343 B.n646 B.n86 585
R1344 B.n649 B.n648 585
R1345 B.n650 B.n85 585
R1346 B.n652 B.n651 585
R1347 B.n654 B.n84 585
R1348 B.n657 B.n656 585
R1349 B.n658 B.n83 585
R1350 B.n660 B.n659 585
R1351 B.n662 B.n82 585
R1352 B.n665 B.n664 585
R1353 B.n666 B.n81 585
R1354 B.n668 B.n667 585
R1355 B.n670 B.n80 585
R1356 B.n673 B.n672 585
R1357 B.n674 B.n79 585
R1358 B.n676 B.n675 585
R1359 B.n678 B.n78 585
R1360 B.n681 B.n680 585
R1361 B.n683 B.n75 585
R1362 B.n685 B.n684 585
R1363 B.n687 B.n74 585
R1364 B.n690 B.n689 585
R1365 B.n691 B.n73 585
R1366 B.n693 B.n692 585
R1367 B.n695 B.n72 585
R1368 B.n697 B.n696 585
R1369 B.n699 B.n698 585
R1370 B.n702 B.n701 585
R1371 B.n703 B.n67 585
R1372 B.n705 B.n704 585
R1373 B.n707 B.n66 585
R1374 B.n710 B.n709 585
R1375 B.n711 B.n65 585
R1376 B.n713 B.n712 585
R1377 B.n715 B.n64 585
R1378 B.n718 B.n717 585
R1379 B.n719 B.n63 585
R1380 B.n721 B.n720 585
R1381 B.n723 B.n62 585
R1382 B.n726 B.n725 585
R1383 B.n727 B.n61 585
R1384 B.n729 B.n728 585
R1385 B.n731 B.n60 585
R1386 B.n734 B.n733 585
R1387 B.n735 B.n59 585
R1388 B.n737 B.n736 585
R1389 B.n739 B.n58 585
R1390 B.n742 B.n741 585
R1391 B.n743 B.n57 585
R1392 B.n745 B.n744 585
R1393 B.n747 B.n56 585
R1394 B.n750 B.n749 585
R1395 B.n751 B.n55 585
R1396 B.n753 B.n752 585
R1397 B.n755 B.n54 585
R1398 B.n758 B.n757 585
R1399 B.n759 B.n53 585
R1400 B.n761 B.n760 585
R1401 B.n763 B.n52 585
R1402 B.n766 B.n765 585
R1403 B.n767 B.n51 585
R1404 B.n769 B.n768 585
R1405 B.n771 B.n50 585
R1406 B.n774 B.n773 585
R1407 B.n775 B.n49 585
R1408 B.n777 B.n776 585
R1409 B.n779 B.n48 585
R1410 B.n782 B.n781 585
R1411 B.n783 B.n47 585
R1412 B.n785 B.n784 585
R1413 B.n787 B.n46 585
R1414 B.n790 B.n789 585
R1415 B.n791 B.n45 585
R1416 B.n793 B.n792 585
R1417 B.n795 B.n44 585
R1418 B.n798 B.n797 585
R1419 B.n799 B.n43 585
R1420 B.n801 B.n800 585
R1421 B.n803 B.n42 585
R1422 B.n806 B.n805 585
R1423 B.n807 B.n41 585
R1424 B.n809 B.n808 585
R1425 B.n811 B.n40 585
R1426 B.n814 B.n813 585
R1427 B.n815 B.n39 585
R1428 B.n817 B.n816 585
R1429 B.n819 B.n38 585
R1430 B.n822 B.n821 585
R1431 B.n823 B.n37 585
R1432 B.n556 B.n35 585
R1433 B.n826 B.n35 585
R1434 B.n555 B.n34 585
R1435 B.n827 B.n34 585
R1436 B.n554 B.n33 585
R1437 B.n828 B.n33 585
R1438 B.n553 B.n552 585
R1439 B.n552 B.n29 585
R1440 B.n551 B.n28 585
R1441 B.n834 B.n28 585
R1442 B.n550 B.n27 585
R1443 B.n835 B.n27 585
R1444 B.n549 B.n26 585
R1445 B.n836 B.n26 585
R1446 B.n548 B.n547 585
R1447 B.n547 B.n22 585
R1448 B.n546 B.n21 585
R1449 B.n842 B.n21 585
R1450 B.n545 B.n20 585
R1451 B.n843 B.n20 585
R1452 B.n544 B.n19 585
R1453 B.n844 B.n19 585
R1454 B.n543 B.n542 585
R1455 B.n542 B.n18 585
R1456 B.n541 B.n14 585
R1457 B.n850 B.n14 585
R1458 B.n540 B.n13 585
R1459 B.n851 B.n13 585
R1460 B.n539 B.n12 585
R1461 B.n852 B.n12 585
R1462 B.n538 B.n537 585
R1463 B.n537 B.n8 585
R1464 B.n536 B.n7 585
R1465 B.n858 B.n7 585
R1466 B.n535 B.n6 585
R1467 B.n859 B.n6 585
R1468 B.n534 B.n5 585
R1469 B.n860 B.n5 585
R1470 B.n533 B.n532 585
R1471 B.n532 B.n4 585
R1472 B.n531 B.n108 585
R1473 B.n531 B.n530 585
R1474 B.n521 B.n109 585
R1475 B.n110 B.n109 585
R1476 B.n523 B.n522 585
R1477 B.n524 B.n523 585
R1478 B.n520 B.n115 585
R1479 B.n115 B.n114 585
R1480 B.n519 B.n518 585
R1481 B.n518 B.n517 585
R1482 B.n117 B.n116 585
R1483 B.n510 B.n117 585
R1484 B.n509 B.n508 585
R1485 B.n511 B.n509 585
R1486 B.n507 B.n122 585
R1487 B.n122 B.n121 585
R1488 B.n506 B.n505 585
R1489 B.n505 B.n504 585
R1490 B.n124 B.n123 585
R1491 B.n125 B.n124 585
R1492 B.n497 B.n496 585
R1493 B.n498 B.n497 585
R1494 B.n495 B.n130 585
R1495 B.n130 B.n129 585
R1496 B.n494 B.n493 585
R1497 B.n493 B.n492 585
R1498 B.n132 B.n131 585
R1499 B.n133 B.n132 585
R1500 B.n485 B.n484 585
R1501 B.n486 B.n485 585
R1502 B.n483 B.n138 585
R1503 B.n138 B.n137 585
R1504 B.n482 B.n481 585
R1505 B.n481 B.n480 585
R1506 B.n477 B.n142 585
R1507 B.n476 B.n475 585
R1508 B.n473 B.n143 585
R1509 B.n473 B.n141 585
R1510 B.n472 B.n471 585
R1511 B.n470 B.n469 585
R1512 B.n468 B.n145 585
R1513 B.n466 B.n465 585
R1514 B.n464 B.n146 585
R1515 B.n463 B.n462 585
R1516 B.n460 B.n147 585
R1517 B.n458 B.n457 585
R1518 B.n456 B.n148 585
R1519 B.n455 B.n454 585
R1520 B.n452 B.n149 585
R1521 B.n450 B.n449 585
R1522 B.n448 B.n150 585
R1523 B.n447 B.n446 585
R1524 B.n444 B.n151 585
R1525 B.n442 B.n441 585
R1526 B.n440 B.n152 585
R1527 B.n439 B.n438 585
R1528 B.n436 B.n153 585
R1529 B.n434 B.n433 585
R1530 B.n432 B.n154 585
R1531 B.n431 B.n430 585
R1532 B.n428 B.n155 585
R1533 B.n426 B.n425 585
R1534 B.n424 B.n156 585
R1535 B.n423 B.n422 585
R1536 B.n420 B.n157 585
R1537 B.n418 B.n417 585
R1538 B.n416 B.n158 585
R1539 B.n415 B.n414 585
R1540 B.n412 B.n159 585
R1541 B.n410 B.n409 585
R1542 B.n408 B.n160 585
R1543 B.n407 B.n406 585
R1544 B.n404 B.n161 585
R1545 B.n402 B.n401 585
R1546 B.n400 B.n162 585
R1547 B.n399 B.n398 585
R1548 B.n396 B.n163 585
R1549 B.n394 B.n393 585
R1550 B.n392 B.n164 585
R1551 B.n391 B.n390 585
R1552 B.n388 B.n165 585
R1553 B.n386 B.n385 585
R1554 B.n384 B.n166 585
R1555 B.n383 B.n382 585
R1556 B.n380 B.n167 585
R1557 B.n378 B.n377 585
R1558 B.n376 B.n168 585
R1559 B.n375 B.n374 585
R1560 B.n372 B.n169 585
R1561 B.n370 B.n369 585
R1562 B.n368 B.n170 585
R1563 B.n367 B.n366 585
R1564 B.n364 B.n171 585
R1565 B.n362 B.n361 585
R1566 B.n360 B.n172 585
R1567 B.n359 B.n358 585
R1568 B.n356 B.n173 585
R1569 B.n354 B.n353 585
R1570 B.n352 B.n174 585
R1571 B.n351 B.n350 585
R1572 B.n348 B.n178 585
R1573 B.n346 B.n345 585
R1574 B.n344 B.n179 585
R1575 B.n343 B.n342 585
R1576 B.n340 B.n180 585
R1577 B.n338 B.n337 585
R1578 B.n335 B.n181 585
R1579 B.n334 B.n333 585
R1580 B.n331 B.n184 585
R1581 B.n329 B.n328 585
R1582 B.n327 B.n185 585
R1583 B.n326 B.n325 585
R1584 B.n323 B.n186 585
R1585 B.n321 B.n320 585
R1586 B.n319 B.n187 585
R1587 B.n318 B.n317 585
R1588 B.n315 B.n188 585
R1589 B.n313 B.n312 585
R1590 B.n311 B.n189 585
R1591 B.n310 B.n309 585
R1592 B.n307 B.n190 585
R1593 B.n305 B.n304 585
R1594 B.n303 B.n191 585
R1595 B.n302 B.n301 585
R1596 B.n299 B.n192 585
R1597 B.n297 B.n296 585
R1598 B.n295 B.n193 585
R1599 B.n294 B.n293 585
R1600 B.n291 B.n194 585
R1601 B.n289 B.n288 585
R1602 B.n287 B.n195 585
R1603 B.n286 B.n285 585
R1604 B.n283 B.n196 585
R1605 B.n281 B.n280 585
R1606 B.n279 B.n197 585
R1607 B.n278 B.n277 585
R1608 B.n275 B.n198 585
R1609 B.n273 B.n272 585
R1610 B.n271 B.n199 585
R1611 B.n270 B.n269 585
R1612 B.n267 B.n200 585
R1613 B.n265 B.n264 585
R1614 B.n263 B.n201 585
R1615 B.n262 B.n261 585
R1616 B.n259 B.n202 585
R1617 B.n257 B.n256 585
R1618 B.n255 B.n203 585
R1619 B.n254 B.n253 585
R1620 B.n251 B.n204 585
R1621 B.n249 B.n248 585
R1622 B.n247 B.n205 585
R1623 B.n246 B.n245 585
R1624 B.n243 B.n206 585
R1625 B.n241 B.n240 585
R1626 B.n239 B.n207 585
R1627 B.n238 B.n237 585
R1628 B.n235 B.n208 585
R1629 B.n233 B.n232 585
R1630 B.n231 B.n209 585
R1631 B.n230 B.n229 585
R1632 B.n227 B.n210 585
R1633 B.n225 B.n224 585
R1634 B.n223 B.n211 585
R1635 B.n222 B.n221 585
R1636 B.n219 B.n212 585
R1637 B.n217 B.n216 585
R1638 B.n215 B.n214 585
R1639 B.n140 B.n139 585
R1640 B.n479 B.n478 585
R1641 B.n480 B.n479 585
R1642 B.n136 B.n135 585
R1643 B.n137 B.n136 585
R1644 B.n488 B.n487 585
R1645 B.n487 B.n486 585
R1646 B.n489 B.n134 585
R1647 B.n134 B.n133 585
R1648 B.n491 B.n490 585
R1649 B.n492 B.n491 585
R1650 B.n128 B.n127 585
R1651 B.n129 B.n128 585
R1652 B.n500 B.n499 585
R1653 B.n499 B.n498 585
R1654 B.n501 B.n126 585
R1655 B.n126 B.n125 585
R1656 B.n503 B.n502 585
R1657 B.n504 B.n503 585
R1658 B.n120 B.n119 585
R1659 B.n121 B.n120 585
R1660 B.n513 B.n512 585
R1661 B.n512 B.n511 585
R1662 B.n514 B.n118 585
R1663 B.n510 B.n118 585
R1664 B.n516 B.n515 585
R1665 B.n517 B.n516 585
R1666 B.n113 B.n112 585
R1667 B.n114 B.n113 585
R1668 B.n526 B.n525 585
R1669 B.n525 B.n524 585
R1670 B.n527 B.n111 585
R1671 B.n111 B.n110 585
R1672 B.n529 B.n528 585
R1673 B.n530 B.n529 585
R1674 B.n2 B.n0 585
R1675 B.n4 B.n2 585
R1676 B.n3 B.n1 585
R1677 B.n859 B.n3 585
R1678 B.n857 B.n856 585
R1679 B.n858 B.n857 585
R1680 B.n855 B.n9 585
R1681 B.n9 B.n8 585
R1682 B.n854 B.n853 585
R1683 B.n853 B.n852 585
R1684 B.n11 B.n10 585
R1685 B.n851 B.n11 585
R1686 B.n849 B.n848 585
R1687 B.n850 B.n849 585
R1688 B.n847 B.n15 585
R1689 B.n18 B.n15 585
R1690 B.n846 B.n845 585
R1691 B.n845 B.n844 585
R1692 B.n17 B.n16 585
R1693 B.n843 B.n17 585
R1694 B.n841 B.n840 585
R1695 B.n842 B.n841 585
R1696 B.n839 B.n23 585
R1697 B.n23 B.n22 585
R1698 B.n838 B.n837 585
R1699 B.n837 B.n836 585
R1700 B.n25 B.n24 585
R1701 B.n835 B.n25 585
R1702 B.n833 B.n832 585
R1703 B.n834 B.n833 585
R1704 B.n831 B.n30 585
R1705 B.n30 B.n29 585
R1706 B.n830 B.n829 585
R1707 B.n829 B.n828 585
R1708 B.n32 B.n31 585
R1709 B.n827 B.n32 585
R1710 B.n825 B.n824 585
R1711 B.n826 B.n825 585
R1712 B.n862 B.n861 585
R1713 B.n861 B.n860 585
R1714 B.n479 B.n142 559.769
R1715 B.n825 B.n37 559.769
R1716 B.n481 B.n140 559.769
R1717 B.n558 B.n35 559.769
R1718 B.n182 B.t10 422.793
R1719 B.n76 B.t16 422.793
R1720 B.n175 B.t7 422.793
R1721 B.n68 B.t13 422.793
R1722 B.n183 B.t9 400.49
R1723 B.n77 B.t17 400.49
R1724 B.n176 B.t6 400.49
R1725 B.n69 B.t14 400.49
R1726 B.n559 B.n36 256.663
R1727 B.n565 B.n36 256.663
R1728 B.n567 B.n36 256.663
R1729 B.n573 B.n36 256.663
R1730 B.n575 B.n36 256.663
R1731 B.n581 B.n36 256.663
R1732 B.n583 B.n36 256.663
R1733 B.n589 B.n36 256.663
R1734 B.n591 B.n36 256.663
R1735 B.n597 B.n36 256.663
R1736 B.n599 B.n36 256.663
R1737 B.n605 B.n36 256.663
R1738 B.n607 B.n36 256.663
R1739 B.n613 B.n36 256.663
R1740 B.n615 B.n36 256.663
R1741 B.n621 B.n36 256.663
R1742 B.n623 B.n36 256.663
R1743 B.n629 B.n36 256.663
R1744 B.n631 B.n36 256.663
R1745 B.n637 B.n36 256.663
R1746 B.n639 B.n36 256.663
R1747 B.n645 B.n36 256.663
R1748 B.n647 B.n36 256.663
R1749 B.n653 B.n36 256.663
R1750 B.n655 B.n36 256.663
R1751 B.n661 B.n36 256.663
R1752 B.n663 B.n36 256.663
R1753 B.n669 B.n36 256.663
R1754 B.n671 B.n36 256.663
R1755 B.n677 B.n36 256.663
R1756 B.n679 B.n36 256.663
R1757 B.n686 B.n36 256.663
R1758 B.n688 B.n36 256.663
R1759 B.n694 B.n36 256.663
R1760 B.n71 B.n36 256.663
R1761 B.n700 B.n36 256.663
R1762 B.n706 B.n36 256.663
R1763 B.n708 B.n36 256.663
R1764 B.n714 B.n36 256.663
R1765 B.n716 B.n36 256.663
R1766 B.n722 B.n36 256.663
R1767 B.n724 B.n36 256.663
R1768 B.n730 B.n36 256.663
R1769 B.n732 B.n36 256.663
R1770 B.n738 B.n36 256.663
R1771 B.n740 B.n36 256.663
R1772 B.n746 B.n36 256.663
R1773 B.n748 B.n36 256.663
R1774 B.n754 B.n36 256.663
R1775 B.n756 B.n36 256.663
R1776 B.n762 B.n36 256.663
R1777 B.n764 B.n36 256.663
R1778 B.n770 B.n36 256.663
R1779 B.n772 B.n36 256.663
R1780 B.n778 B.n36 256.663
R1781 B.n780 B.n36 256.663
R1782 B.n786 B.n36 256.663
R1783 B.n788 B.n36 256.663
R1784 B.n794 B.n36 256.663
R1785 B.n796 B.n36 256.663
R1786 B.n802 B.n36 256.663
R1787 B.n804 B.n36 256.663
R1788 B.n810 B.n36 256.663
R1789 B.n812 B.n36 256.663
R1790 B.n818 B.n36 256.663
R1791 B.n820 B.n36 256.663
R1792 B.n474 B.n141 256.663
R1793 B.n144 B.n141 256.663
R1794 B.n467 B.n141 256.663
R1795 B.n461 B.n141 256.663
R1796 B.n459 B.n141 256.663
R1797 B.n453 B.n141 256.663
R1798 B.n451 B.n141 256.663
R1799 B.n445 B.n141 256.663
R1800 B.n443 B.n141 256.663
R1801 B.n437 B.n141 256.663
R1802 B.n435 B.n141 256.663
R1803 B.n429 B.n141 256.663
R1804 B.n427 B.n141 256.663
R1805 B.n421 B.n141 256.663
R1806 B.n419 B.n141 256.663
R1807 B.n413 B.n141 256.663
R1808 B.n411 B.n141 256.663
R1809 B.n405 B.n141 256.663
R1810 B.n403 B.n141 256.663
R1811 B.n397 B.n141 256.663
R1812 B.n395 B.n141 256.663
R1813 B.n389 B.n141 256.663
R1814 B.n387 B.n141 256.663
R1815 B.n381 B.n141 256.663
R1816 B.n379 B.n141 256.663
R1817 B.n373 B.n141 256.663
R1818 B.n371 B.n141 256.663
R1819 B.n365 B.n141 256.663
R1820 B.n363 B.n141 256.663
R1821 B.n357 B.n141 256.663
R1822 B.n355 B.n141 256.663
R1823 B.n349 B.n141 256.663
R1824 B.n347 B.n141 256.663
R1825 B.n341 B.n141 256.663
R1826 B.n339 B.n141 256.663
R1827 B.n332 B.n141 256.663
R1828 B.n330 B.n141 256.663
R1829 B.n324 B.n141 256.663
R1830 B.n322 B.n141 256.663
R1831 B.n316 B.n141 256.663
R1832 B.n314 B.n141 256.663
R1833 B.n308 B.n141 256.663
R1834 B.n306 B.n141 256.663
R1835 B.n300 B.n141 256.663
R1836 B.n298 B.n141 256.663
R1837 B.n292 B.n141 256.663
R1838 B.n290 B.n141 256.663
R1839 B.n284 B.n141 256.663
R1840 B.n282 B.n141 256.663
R1841 B.n276 B.n141 256.663
R1842 B.n274 B.n141 256.663
R1843 B.n268 B.n141 256.663
R1844 B.n266 B.n141 256.663
R1845 B.n260 B.n141 256.663
R1846 B.n258 B.n141 256.663
R1847 B.n252 B.n141 256.663
R1848 B.n250 B.n141 256.663
R1849 B.n244 B.n141 256.663
R1850 B.n242 B.n141 256.663
R1851 B.n236 B.n141 256.663
R1852 B.n234 B.n141 256.663
R1853 B.n228 B.n141 256.663
R1854 B.n226 B.n141 256.663
R1855 B.n220 B.n141 256.663
R1856 B.n218 B.n141 256.663
R1857 B.n213 B.n141 256.663
R1858 B.n479 B.n136 163.367
R1859 B.n487 B.n136 163.367
R1860 B.n487 B.n134 163.367
R1861 B.n491 B.n134 163.367
R1862 B.n491 B.n128 163.367
R1863 B.n499 B.n128 163.367
R1864 B.n499 B.n126 163.367
R1865 B.n503 B.n126 163.367
R1866 B.n503 B.n120 163.367
R1867 B.n512 B.n120 163.367
R1868 B.n512 B.n118 163.367
R1869 B.n516 B.n118 163.367
R1870 B.n516 B.n113 163.367
R1871 B.n525 B.n113 163.367
R1872 B.n525 B.n111 163.367
R1873 B.n529 B.n111 163.367
R1874 B.n529 B.n2 163.367
R1875 B.n861 B.n2 163.367
R1876 B.n861 B.n3 163.367
R1877 B.n857 B.n3 163.367
R1878 B.n857 B.n9 163.367
R1879 B.n853 B.n9 163.367
R1880 B.n853 B.n11 163.367
R1881 B.n849 B.n11 163.367
R1882 B.n849 B.n15 163.367
R1883 B.n845 B.n15 163.367
R1884 B.n845 B.n17 163.367
R1885 B.n841 B.n17 163.367
R1886 B.n841 B.n23 163.367
R1887 B.n837 B.n23 163.367
R1888 B.n837 B.n25 163.367
R1889 B.n833 B.n25 163.367
R1890 B.n833 B.n30 163.367
R1891 B.n829 B.n30 163.367
R1892 B.n829 B.n32 163.367
R1893 B.n825 B.n32 163.367
R1894 B.n475 B.n473 163.367
R1895 B.n473 B.n472 163.367
R1896 B.n469 B.n468 163.367
R1897 B.n466 B.n146 163.367
R1898 B.n462 B.n460 163.367
R1899 B.n458 B.n148 163.367
R1900 B.n454 B.n452 163.367
R1901 B.n450 B.n150 163.367
R1902 B.n446 B.n444 163.367
R1903 B.n442 B.n152 163.367
R1904 B.n438 B.n436 163.367
R1905 B.n434 B.n154 163.367
R1906 B.n430 B.n428 163.367
R1907 B.n426 B.n156 163.367
R1908 B.n422 B.n420 163.367
R1909 B.n418 B.n158 163.367
R1910 B.n414 B.n412 163.367
R1911 B.n410 B.n160 163.367
R1912 B.n406 B.n404 163.367
R1913 B.n402 B.n162 163.367
R1914 B.n398 B.n396 163.367
R1915 B.n394 B.n164 163.367
R1916 B.n390 B.n388 163.367
R1917 B.n386 B.n166 163.367
R1918 B.n382 B.n380 163.367
R1919 B.n378 B.n168 163.367
R1920 B.n374 B.n372 163.367
R1921 B.n370 B.n170 163.367
R1922 B.n366 B.n364 163.367
R1923 B.n362 B.n172 163.367
R1924 B.n358 B.n356 163.367
R1925 B.n354 B.n174 163.367
R1926 B.n350 B.n348 163.367
R1927 B.n346 B.n179 163.367
R1928 B.n342 B.n340 163.367
R1929 B.n338 B.n181 163.367
R1930 B.n333 B.n331 163.367
R1931 B.n329 B.n185 163.367
R1932 B.n325 B.n323 163.367
R1933 B.n321 B.n187 163.367
R1934 B.n317 B.n315 163.367
R1935 B.n313 B.n189 163.367
R1936 B.n309 B.n307 163.367
R1937 B.n305 B.n191 163.367
R1938 B.n301 B.n299 163.367
R1939 B.n297 B.n193 163.367
R1940 B.n293 B.n291 163.367
R1941 B.n289 B.n195 163.367
R1942 B.n285 B.n283 163.367
R1943 B.n281 B.n197 163.367
R1944 B.n277 B.n275 163.367
R1945 B.n273 B.n199 163.367
R1946 B.n269 B.n267 163.367
R1947 B.n265 B.n201 163.367
R1948 B.n261 B.n259 163.367
R1949 B.n257 B.n203 163.367
R1950 B.n253 B.n251 163.367
R1951 B.n249 B.n205 163.367
R1952 B.n245 B.n243 163.367
R1953 B.n241 B.n207 163.367
R1954 B.n237 B.n235 163.367
R1955 B.n233 B.n209 163.367
R1956 B.n229 B.n227 163.367
R1957 B.n225 B.n211 163.367
R1958 B.n221 B.n219 163.367
R1959 B.n217 B.n214 163.367
R1960 B.n481 B.n138 163.367
R1961 B.n485 B.n138 163.367
R1962 B.n485 B.n132 163.367
R1963 B.n493 B.n132 163.367
R1964 B.n493 B.n130 163.367
R1965 B.n497 B.n130 163.367
R1966 B.n497 B.n124 163.367
R1967 B.n505 B.n124 163.367
R1968 B.n505 B.n122 163.367
R1969 B.n509 B.n122 163.367
R1970 B.n509 B.n117 163.367
R1971 B.n518 B.n117 163.367
R1972 B.n518 B.n115 163.367
R1973 B.n523 B.n115 163.367
R1974 B.n523 B.n109 163.367
R1975 B.n531 B.n109 163.367
R1976 B.n532 B.n531 163.367
R1977 B.n532 B.n5 163.367
R1978 B.n6 B.n5 163.367
R1979 B.n7 B.n6 163.367
R1980 B.n537 B.n7 163.367
R1981 B.n537 B.n12 163.367
R1982 B.n13 B.n12 163.367
R1983 B.n14 B.n13 163.367
R1984 B.n542 B.n14 163.367
R1985 B.n542 B.n19 163.367
R1986 B.n20 B.n19 163.367
R1987 B.n21 B.n20 163.367
R1988 B.n547 B.n21 163.367
R1989 B.n547 B.n26 163.367
R1990 B.n27 B.n26 163.367
R1991 B.n28 B.n27 163.367
R1992 B.n552 B.n28 163.367
R1993 B.n552 B.n33 163.367
R1994 B.n34 B.n33 163.367
R1995 B.n35 B.n34 163.367
R1996 B.n821 B.n819 163.367
R1997 B.n817 B.n39 163.367
R1998 B.n813 B.n811 163.367
R1999 B.n809 B.n41 163.367
R2000 B.n805 B.n803 163.367
R2001 B.n801 B.n43 163.367
R2002 B.n797 B.n795 163.367
R2003 B.n793 B.n45 163.367
R2004 B.n789 B.n787 163.367
R2005 B.n785 B.n47 163.367
R2006 B.n781 B.n779 163.367
R2007 B.n777 B.n49 163.367
R2008 B.n773 B.n771 163.367
R2009 B.n769 B.n51 163.367
R2010 B.n765 B.n763 163.367
R2011 B.n761 B.n53 163.367
R2012 B.n757 B.n755 163.367
R2013 B.n753 B.n55 163.367
R2014 B.n749 B.n747 163.367
R2015 B.n745 B.n57 163.367
R2016 B.n741 B.n739 163.367
R2017 B.n737 B.n59 163.367
R2018 B.n733 B.n731 163.367
R2019 B.n729 B.n61 163.367
R2020 B.n725 B.n723 163.367
R2021 B.n721 B.n63 163.367
R2022 B.n717 B.n715 163.367
R2023 B.n713 B.n65 163.367
R2024 B.n709 B.n707 163.367
R2025 B.n705 B.n67 163.367
R2026 B.n701 B.n699 163.367
R2027 B.n696 B.n695 163.367
R2028 B.n693 B.n73 163.367
R2029 B.n689 B.n687 163.367
R2030 B.n685 B.n75 163.367
R2031 B.n680 B.n678 163.367
R2032 B.n676 B.n79 163.367
R2033 B.n672 B.n670 163.367
R2034 B.n668 B.n81 163.367
R2035 B.n664 B.n662 163.367
R2036 B.n660 B.n83 163.367
R2037 B.n656 B.n654 163.367
R2038 B.n652 B.n85 163.367
R2039 B.n648 B.n646 163.367
R2040 B.n644 B.n87 163.367
R2041 B.n640 B.n638 163.367
R2042 B.n636 B.n89 163.367
R2043 B.n632 B.n630 163.367
R2044 B.n628 B.n91 163.367
R2045 B.n624 B.n622 163.367
R2046 B.n620 B.n93 163.367
R2047 B.n616 B.n614 163.367
R2048 B.n612 B.n95 163.367
R2049 B.n608 B.n606 163.367
R2050 B.n604 B.n97 163.367
R2051 B.n600 B.n598 163.367
R2052 B.n596 B.n99 163.367
R2053 B.n592 B.n590 163.367
R2054 B.n588 B.n101 163.367
R2055 B.n584 B.n582 163.367
R2056 B.n580 B.n103 163.367
R2057 B.n576 B.n574 163.367
R2058 B.n572 B.n105 163.367
R2059 B.n568 B.n566 163.367
R2060 B.n564 B.n107 163.367
R2061 B.n560 B.n558 163.367
R2062 B.n474 B.n142 71.676
R2063 B.n472 B.n144 71.676
R2064 B.n468 B.n467 71.676
R2065 B.n461 B.n146 71.676
R2066 B.n460 B.n459 71.676
R2067 B.n453 B.n148 71.676
R2068 B.n452 B.n451 71.676
R2069 B.n445 B.n150 71.676
R2070 B.n444 B.n443 71.676
R2071 B.n437 B.n152 71.676
R2072 B.n436 B.n435 71.676
R2073 B.n429 B.n154 71.676
R2074 B.n428 B.n427 71.676
R2075 B.n421 B.n156 71.676
R2076 B.n420 B.n419 71.676
R2077 B.n413 B.n158 71.676
R2078 B.n412 B.n411 71.676
R2079 B.n405 B.n160 71.676
R2080 B.n404 B.n403 71.676
R2081 B.n397 B.n162 71.676
R2082 B.n396 B.n395 71.676
R2083 B.n389 B.n164 71.676
R2084 B.n388 B.n387 71.676
R2085 B.n381 B.n166 71.676
R2086 B.n380 B.n379 71.676
R2087 B.n373 B.n168 71.676
R2088 B.n372 B.n371 71.676
R2089 B.n365 B.n170 71.676
R2090 B.n364 B.n363 71.676
R2091 B.n357 B.n172 71.676
R2092 B.n356 B.n355 71.676
R2093 B.n349 B.n174 71.676
R2094 B.n348 B.n347 71.676
R2095 B.n341 B.n179 71.676
R2096 B.n340 B.n339 71.676
R2097 B.n332 B.n181 71.676
R2098 B.n331 B.n330 71.676
R2099 B.n324 B.n185 71.676
R2100 B.n323 B.n322 71.676
R2101 B.n316 B.n187 71.676
R2102 B.n315 B.n314 71.676
R2103 B.n308 B.n189 71.676
R2104 B.n307 B.n306 71.676
R2105 B.n300 B.n191 71.676
R2106 B.n299 B.n298 71.676
R2107 B.n292 B.n193 71.676
R2108 B.n291 B.n290 71.676
R2109 B.n284 B.n195 71.676
R2110 B.n283 B.n282 71.676
R2111 B.n276 B.n197 71.676
R2112 B.n275 B.n274 71.676
R2113 B.n268 B.n199 71.676
R2114 B.n267 B.n266 71.676
R2115 B.n260 B.n201 71.676
R2116 B.n259 B.n258 71.676
R2117 B.n252 B.n203 71.676
R2118 B.n251 B.n250 71.676
R2119 B.n244 B.n205 71.676
R2120 B.n243 B.n242 71.676
R2121 B.n236 B.n207 71.676
R2122 B.n235 B.n234 71.676
R2123 B.n228 B.n209 71.676
R2124 B.n227 B.n226 71.676
R2125 B.n220 B.n211 71.676
R2126 B.n219 B.n218 71.676
R2127 B.n214 B.n213 71.676
R2128 B.n820 B.n37 71.676
R2129 B.n819 B.n818 71.676
R2130 B.n812 B.n39 71.676
R2131 B.n811 B.n810 71.676
R2132 B.n804 B.n41 71.676
R2133 B.n803 B.n802 71.676
R2134 B.n796 B.n43 71.676
R2135 B.n795 B.n794 71.676
R2136 B.n788 B.n45 71.676
R2137 B.n787 B.n786 71.676
R2138 B.n780 B.n47 71.676
R2139 B.n779 B.n778 71.676
R2140 B.n772 B.n49 71.676
R2141 B.n771 B.n770 71.676
R2142 B.n764 B.n51 71.676
R2143 B.n763 B.n762 71.676
R2144 B.n756 B.n53 71.676
R2145 B.n755 B.n754 71.676
R2146 B.n748 B.n55 71.676
R2147 B.n747 B.n746 71.676
R2148 B.n740 B.n57 71.676
R2149 B.n739 B.n738 71.676
R2150 B.n732 B.n59 71.676
R2151 B.n731 B.n730 71.676
R2152 B.n724 B.n61 71.676
R2153 B.n723 B.n722 71.676
R2154 B.n716 B.n63 71.676
R2155 B.n715 B.n714 71.676
R2156 B.n708 B.n65 71.676
R2157 B.n707 B.n706 71.676
R2158 B.n700 B.n67 71.676
R2159 B.n699 B.n71 71.676
R2160 B.n695 B.n694 71.676
R2161 B.n688 B.n73 71.676
R2162 B.n687 B.n686 71.676
R2163 B.n679 B.n75 71.676
R2164 B.n678 B.n677 71.676
R2165 B.n671 B.n79 71.676
R2166 B.n670 B.n669 71.676
R2167 B.n663 B.n81 71.676
R2168 B.n662 B.n661 71.676
R2169 B.n655 B.n83 71.676
R2170 B.n654 B.n653 71.676
R2171 B.n647 B.n85 71.676
R2172 B.n646 B.n645 71.676
R2173 B.n639 B.n87 71.676
R2174 B.n638 B.n637 71.676
R2175 B.n631 B.n89 71.676
R2176 B.n630 B.n629 71.676
R2177 B.n623 B.n91 71.676
R2178 B.n622 B.n621 71.676
R2179 B.n615 B.n93 71.676
R2180 B.n614 B.n613 71.676
R2181 B.n607 B.n95 71.676
R2182 B.n606 B.n605 71.676
R2183 B.n599 B.n97 71.676
R2184 B.n598 B.n597 71.676
R2185 B.n591 B.n99 71.676
R2186 B.n590 B.n589 71.676
R2187 B.n583 B.n101 71.676
R2188 B.n582 B.n581 71.676
R2189 B.n575 B.n103 71.676
R2190 B.n574 B.n573 71.676
R2191 B.n567 B.n105 71.676
R2192 B.n566 B.n565 71.676
R2193 B.n559 B.n107 71.676
R2194 B.n560 B.n559 71.676
R2195 B.n565 B.n564 71.676
R2196 B.n568 B.n567 71.676
R2197 B.n573 B.n572 71.676
R2198 B.n576 B.n575 71.676
R2199 B.n581 B.n580 71.676
R2200 B.n584 B.n583 71.676
R2201 B.n589 B.n588 71.676
R2202 B.n592 B.n591 71.676
R2203 B.n597 B.n596 71.676
R2204 B.n600 B.n599 71.676
R2205 B.n605 B.n604 71.676
R2206 B.n608 B.n607 71.676
R2207 B.n613 B.n612 71.676
R2208 B.n616 B.n615 71.676
R2209 B.n621 B.n620 71.676
R2210 B.n624 B.n623 71.676
R2211 B.n629 B.n628 71.676
R2212 B.n632 B.n631 71.676
R2213 B.n637 B.n636 71.676
R2214 B.n640 B.n639 71.676
R2215 B.n645 B.n644 71.676
R2216 B.n648 B.n647 71.676
R2217 B.n653 B.n652 71.676
R2218 B.n656 B.n655 71.676
R2219 B.n661 B.n660 71.676
R2220 B.n664 B.n663 71.676
R2221 B.n669 B.n668 71.676
R2222 B.n672 B.n671 71.676
R2223 B.n677 B.n676 71.676
R2224 B.n680 B.n679 71.676
R2225 B.n686 B.n685 71.676
R2226 B.n689 B.n688 71.676
R2227 B.n694 B.n693 71.676
R2228 B.n696 B.n71 71.676
R2229 B.n701 B.n700 71.676
R2230 B.n706 B.n705 71.676
R2231 B.n709 B.n708 71.676
R2232 B.n714 B.n713 71.676
R2233 B.n717 B.n716 71.676
R2234 B.n722 B.n721 71.676
R2235 B.n725 B.n724 71.676
R2236 B.n730 B.n729 71.676
R2237 B.n733 B.n732 71.676
R2238 B.n738 B.n737 71.676
R2239 B.n741 B.n740 71.676
R2240 B.n746 B.n745 71.676
R2241 B.n749 B.n748 71.676
R2242 B.n754 B.n753 71.676
R2243 B.n757 B.n756 71.676
R2244 B.n762 B.n761 71.676
R2245 B.n765 B.n764 71.676
R2246 B.n770 B.n769 71.676
R2247 B.n773 B.n772 71.676
R2248 B.n778 B.n777 71.676
R2249 B.n781 B.n780 71.676
R2250 B.n786 B.n785 71.676
R2251 B.n789 B.n788 71.676
R2252 B.n794 B.n793 71.676
R2253 B.n797 B.n796 71.676
R2254 B.n802 B.n801 71.676
R2255 B.n805 B.n804 71.676
R2256 B.n810 B.n809 71.676
R2257 B.n813 B.n812 71.676
R2258 B.n818 B.n817 71.676
R2259 B.n821 B.n820 71.676
R2260 B.n475 B.n474 71.676
R2261 B.n469 B.n144 71.676
R2262 B.n467 B.n466 71.676
R2263 B.n462 B.n461 71.676
R2264 B.n459 B.n458 71.676
R2265 B.n454 B.n453 71.676
R2266 B.n451 B.n450 71.676
R2267 B.n446 B.n445 71.676
R2268 B.n443 B.n442 71.676
R2269 B.n438 B.n437 71.676
R2270 B.n435 B.n434 71.676
R2271 B.n430 B.n429 71.676
R2272 B.n427 B.n426 71.676
R2273 B.n422 B.n421 71.676
R2274 B.n419 B.n418 71.676
R2275 B.n414 B.n413 71.676
R2276 B.n411 B.n410 71.676
R2277 B.n406 B.n405 71.676
R2278 B.n403 B.n402 71.676
R2279 B.n398 B.n397 71.676
R2280 B.n395 B.n394 71.676
R2281 B.n390 B.n389 71.676
R2282 B.n387 B.n386 71.676
R2283 B.n382 B.n381 71.676
R2284 B.n379 B.n378 71.676
R2285 B.n374 B.n373 71.676
R2286 B.n371 B.n370 71.676
R2287 B.n366 B.n365 71.676
R2288 B.n363 B.n362 71.676
R2289 B.n358 B.n357 71.676
R2290 B.n355 B.n354 71.676
R2291 B.n350 B.n349 71.676
R2292 B.n347 B.n346 71.676
R2293 B.n342 B.n341 71.676
R2294 B.n339 B.n338 71.676
R2295 B.n333 B.n332 71.676
R2296 B.n330 B.n329 71.676
R2297 B.n325 B.n324 71.676
R2298 B.n322 B.n321 71.676
R2299 B.n317 B.n316 71.676
R2300 B.n314 B.n313 71.676
R2301 B.n309 B.n308 71.676
R2302 B.n306 B.n305 71.676
R2303 B.n301 B.n300 71.676
R2304 B.n298 B.n297 71.676
R2305 B.n293 B.n292 71.676
R2306 B.n290 B.n289 71.676
R2307 B.n285 B.n284 71.676
R2308 B.n282 B.n281 71.676
R2309 B.n277 B.n276 71.676
R2310 B.n274 B.n273 71.676
R2311 B.n269 B.n268 71.676
R2312 B.n266 B.n265 71.676
R2313 B.n261 B.n260 71.676
R2314 B.n258 B.n257 71.676
R2315 B.n253 B.n252 71.676
R2316 B.n250 B.n249 71.676
R2317 B.n245 B.n244 71.676
R2318 B.n242 B.n241 71.676
R2319 B.n237 B.n236 71.676
R2320 B.n234 B.n233 71.676
R2321 B.n229 B.n228 71.676
R2322 B.n226 B.n225 71.676
R2323 B.n221 B.n220 71.676
R2324 B.n218 B.n217 71.676
R2325 B.n213 B.n140 71.676
R2326 B.n480 B.n141 64.2374
R2327 B.n826 B.n36 64.2374
R2328 B.n336 B.n183 59.5399
R2329 B.n177 B.n176 59.5399
R2330 B.n70 B.n69 59.5399
R2331 B.n682 B.n77 59.5399
R2332 B.n557 B.n556 36.3712
R2333 B.n824 B.n823 36.3712
R2334 B.n482 B.n139 36.3712
R2335 B.n478 B.n477 36.3712
R2336 B.n480 B.n137 30.98
R2337 B.n486 B.n137 30.98
R2338 B.n486 B.n133 30.98
R2339 B.n492 B.n133 30.98
R2340 B.n498 B.n129 30.98
R2341 B.n498 B.n125 30.98
R2342 B.n504 B.n125 30.98
R2343 B.n504 B.n121 30.98
R2344 B.n511 B.n121 30.98
R2345 B.n511 B.n510 30.98
R2346 B.n517 B.n114 30.98
R2347 B.n524 B.n114 30.98
R2348 B.n530 B.n110 30.98
R2349 B.n530 B.n4 30.98
R2350 B.n860 B.n4 30.98
R2351 B.n860 B.n859 30.98
R2352 B.n859 B.n858 30.98
R2353 B.n858 B.n8 30.98
R2354 B.n852 B.n851 30.98
R2355 B.n851 B.n850 30.98
R2356 B.n844 B.n18 30.98
R2357 B.n844 B.n843 30.98
R2358 B.n843 B.n842 30.98
R2359 B.n842 B.n22 30.98
R2360 B.n836 B.n22 30.98
R2361 B.n836 B.n835 30.98
R2362 B.n834 B.n29 30.98
R2363 B.n828 B.n29 30.98
R2364 B.n828 B.n827 30.98
R2365 B.n827 B.n826 30.98
R2366 B.n492 B.t5 22.7795
R2367 B.t12 B.n834 22.7795
R2368 B.n183 B.n182 22.3035
R2369 B.n176 B.n175 22.3035
R2370 B.n69 B.n68 22.3035
R2371 B.n77 B.n76 22.3035
R2372 B.n524 B.t3 21.8684
R2373 B.n852 B.t2 21.8684
R2374 B.n517 B.t0 20.9572
R2375 B.n850 B.t1 20.9572
R2376 B B.n862 18.0485
R2377 B.n823 B.n822 10.6151
R2378 B.n822 B.n38 10.6151
R2379 B.n816 B.n38 10.6151
R2380 B.n816 B.n815 10.6151
R2381 B.n815 B.n814 10.6151
R2382 B.n814 B.n40 10.6151
R2383 B.n808 B.n40 10.6151
R2384 B.n808 B.n807 10.6151
R2385 B.n807 B.n806 10.6151
R2386 B.n806 B.n42 10.6151
R2387 B.n800 B.n42 10.6151
R2388 B.n800 B.n799 10.6151
R2389 B.n799 B.n798 10.6151
R2390 B.n798 B.n44 10.6151
R2391 B.n792 B.n44 10.6151
R2392 B.n792 B.n791 10.6151
R2393 B.n791 B.n790 10.6151
R2394 B.n790 B.n46 10.6151
R2395 B.n784 B.n46 10.6151
R2396 B.n784 B.n783 10.6151
R2397 B.n783 B.n782 10.6151
R2398 B.n782 B.n48 10.6151
R2399 B.n776 B.n48 10.6151
R2400 B.n776 B.n775 10.6151
R2401 B.n775 B.n774 10.6151
R2402 B.n774 B.n50 10.6151
R2403 B.n768 B.n50 10.6151
R2404 B.n768 B.n767 10.6151
R2405 B.n767 B.n766 10.6151
R2406 B.n766 B.n52 10.6151
R2407 B.n760 B.n52 10.6151
R2408 B.n760 B.n759 10.6151
R2409 B.n759 B.n758 10.6151
R2410 B.n758 B.n54 10.6151
R2411 B.n752 B.n54 10.6151
R2412 B.n752 B.n751 10.6151
R2413 B.n751 B.n750 10.6151
R2414 B.n750 B.n56 10.6151
R2415 B.n744 B.n56 10.6151
R2416 B.n744 B.n743 10.6151
R2417 B.n743 B.n742 10.6151
R2418 B.n742 B.n58 10.6151
R2419 B.n736 B.n58 10.6151
R2420 B.n736 B.n735 10.6151
R2421 B.n735 B.n734 10.6151
R2422 B.n734 B.n60 10.6151
R2423 B.n728 B.n60 10.6151
R2424 B.n728 B.n727 10.6151
R2425 B.n727 B.n726 10.6151
R2426 B.n726 B.n62 10.6151
R2427 B.n720 B.n62 10.6151
R2428 B.n720 B.n719 10.6151
R2429 B.n719 B.n718 10.6151
R2430 B.n718 B.n64 10.6151
R2431 B.n712 B.n64 10.6151
R2432 B.n712 B.n711 10.6151
R2433 B.n711 B.n710 10.6151
R2434 B.n710 B.n66 10.6151
R2435 B.n704 B.n66 10.6151
R2436 B.n704 B.n703 10.6151
R2437 B.n703 B.n702 10.6151
R2438 B.n698 B.n697 10.6151
R2439 B.n697 B.n72 10.6151
R2440 B.n692 B.n72 10.6151
R2441 B.n692 B.n691 10.6151
R2442 B.n691 B.n690 10.6151
R2443 B.n690 B.n74 10.6151
R2444 B.n684 B.n74 10.6151
R2445 B.n684 B.n683 10.6151
R2446 B.n681 B.n78 10.6151
R2447 B.n675 B.n78 10.6151
R2448 B.n675 B.n674 10.6151
R2449 B.n674 B.n673 10.6151
R2450 B.n673 B.n80 10.6151
R2451 B.n667 B.n80 10.6151
R2452 B.n667 B.n666 10.6151
R2453 B.n666 B.n665 10.6151
R2454 B.n665 B.n82 10.6151
R2455 B.n659 B.n82 10.6151
R2456 B.n659 B.n658 10.6151
R2457 B.n658 B.n657 10.6151
R2458 B.n657 B.n84 10.6151
R2459 B.n651 B.n84 10.6151
R2460 B.n651 B.n650 10.6151
R2461 B.n650 B.n649 10.6151
R2462 B.n649 B.n86 10.6151
R2463 B.n643 B.n86 10.6151
R2464 B.n643 B.n642 10.6151
R2465 B.n642 B.n641 10.6151
R2466 B.n641 B.n88 10.6151
R2467 B.n635 B.n88 10.6151
R2468 B.n635 B.n634 10.6151
R2469 B.n634 B.n633 10.6151
R2470 B.n633 B.n90 10.6151
R2471 B.n627 B.n90 10.6151
R2472 B.n627 B.n626 10.6151
R2473 B.n626 B.n625 10.6151
R2474 B.n625 B.n92 10.6151
R2475 B.n619 B.n92 10.6151
R2476 B.n619 B.n618 10.6151
R2477 B.n618 B.n617 10.6151
R2478 B.n617 B.n94 10.6151
R2479 B.n611 B.n94 10.6151
R2480 B.n611 B.n610 10.6151
R2481 B.n610 B.n609 10.6151
R2482 B.n609 B.n96 10.6151
R2483 B.n603 B.n96 10.6151
R2484 B.n603 B.n602 10.6151
R2485 B.n602 B.n601 10.6151
R2486 B.n601 B.n98 10.6151
R2487 B.n595 B.n98 10.6151
R2488 B.n595 B.n594 10.6151
R2489 B.n594 B.n593 10.6151
R2490 B.n593 B.n100 10.6151
R2491 B.n587 B.n100 10.6151
R2492 B.n587 B.n586 10.6151
R2493 B.n586 B.n585 10.6151
R2494 B.n585 B.n102 10.6151
R2495 B.n579 B.n102 10.6151
R2496 B.n579 B.n578 10.6151
R2497 B.n578 B.n577 10.6151
R2498 B.n577 B.n104 10.6151
R2499 B.n571 B.n104 10.6151
R2500 B.n571 B.n570 10.6151
R2501 B.n570 B.n569 10.6151
R2502 B.n569 B.n106 10.6151
R2503 B.n563 B.n106 10.6151
R2504 B.n563 B.n562 10.6151
R2505 B.n562 B.n561 10.6151
R2506 B.n561 B.n557 10.6151
R2507 B.n483 B.n482 10.6151
R2508 B.n484 B.n483 10.6151
R2509 B.n484 B.n131 10.6151
R2510 B.n494 B.n131 10.6151
R2511 B.n495 B.n494 10.6151
R2512 B.n496 B.n495 10.6151
R2513 B.n496 B.n123 10.6151
R2514 B.n506 B.n123 10.6151
R2515 B.n507 B.n506 10.6151
R2516 B.n508 B.n507 10.6151
R2517 B.n508 B.n116 10.6151
R2518 B.n519 B.n116 10.6151
R2519 B.n520 B.n519 10.6151
R2520 B.n522 B.n520 10.6151
R2521 B.n522 B.n521 10.6151
R2522 B.n521 B.n108 10.6151
R2523 B.n533 B.n108 10.6151
R2524 B.n534 B.n533 10.6151
R2525 B.n535 B.n534 10.6151
R2526 B.n536 B.n535 10.6151
R2527 B.n538 B.n536 10.6151
R2528 B.n539 B.n538 10.6151
R2529 B.n540 B.n539 10.6151
R2530 B.n541 B.n540 10.6151
R2531 B.n543 B.n541 10.6151
R2532 B.n544 B.n543 10.6151
R2533 B.n545 B.n544 10.6151
R2534 B.n546 B.n545 10.6151
R2535 B.n548 B.n546 10.6151
R2536 B.n549 B.n548 10.6151
R2537 B.n550 B.n549 10.6151
R2538 B.n551 B.n550 10.6151
R2539 B.n553 B.n551 10.6151
R2540 B.n554 B.n553 10.6151
R2541 B.n555 B.n554 10.6151
R2542 B.n556 B.n555 10.6151
R2543 B.n477 B.n476 10.6151
R2544 B.n476 B.n143 10.6151
R2545 B.n471 B.n143 10.6151
R2546 B.n471 B.n470 10.6151
R2547 B.n470 B.n145 10.6151
R2548 B.n465 B.n145 10.6151
R2549 B.n465 B.n464 10.6151
R2550 B.n464 B.n463 10.6151
R2551 B.n463 B.n147 10.6151
R2552 B.n457 B.n147 10.6151
R2553 B.n457 B.n456 10.6151
R2554 B.n456 B.n455 10.6151
R2555 B.n455 B.n149 10.6151
R2556 B.n449 B.n149 10.6151
R2557 B.n449 B.n448 10.6151
R2558 B.n448 B.n447 10.6151
R2559 B.n447 B.n151 10.6151
R2560 B.n441 B.n151 10.6151
R2561 B.n441 B.n440 10.6151
R2562 B.n440 B.n439 10.6151
R2563 B.n439 B.n153 10.6151
R2564 B.n433 B.n153 10.6151
R2565 B.n433 B.n432 10.6151
R2566 B.n432 B.n431 10.6151
R2567 B.n431 B.n155 10.6151
R2568 B.n425 B.n155 10.6151
R2569 B.n425 B.n424 10.6151
R2570 B.n424 B.n423 10.6151
R2571 B.n423 B.n157 10.6151
R2572 B.n417 B.n157 10.6151
R2573 B.n417 B.n416 10.6151
R2574 B.n416 B.n415 10.6151
R2575 B.n415 B.n159 10.6151
R2576 B.n409 B.n159 10.6151
R2577 B.n409 B.n408 10.6151
R2578 B.n408 B.n407 10.6151
R2579 B.n407 B.n161 10.6151
R2580 B.n401 B.n161 10.6151
R2581 B.n401 B.n400 10.6151
R2582 B.n400 B.n399 10.6151
R2583 B.n399 B.n163 10.6151
R2584 B.n393 B.n163 10.6151
R2585 B.n393 B.n392 10.6151
R2586 B.n392 B.n391 10.6151
R2587 B.n391 B.n165 10.6151
R2588 B.n385 B.n165 10.6151
R2589 B.n385 B.n384 10.6151
R2590 B.n384 B.n383 10.6151
R2591 B.n383 B.n167 10.6151
R2592 B.n377 B.n167 10.6151
R2593 B.n377 B.n376 10.6151
R2594 B.n376 B.n375 10.6151
R2595 B.n375 B.n169 10.6151
R2596 B.n369 B.n169 10.6151
R2597 B.n369 B.n368 10.6151
R2598 B.n368 B.n367 10.6151
R2599 B.n367 B.n171 10.6151
R2600 B.n361 B.n171 10.6151
R2601 B.n361 B.n360 10.6151
R2602 B.n360 B.n359 10.6151
R2603 B.n359 B.n173 10.6151
R2604 B.n353 B.n352 10.6151
R2605 B.n352 B.n351 10.6151
R2606 B.n351 B.n178 10.6151
R2607 B.n345 B.n178 10.6151
R2608 B.n345 B.n344 10.6151
R2609 B.n344 B.n343 10.6151
R2610 B.n343 B.n180 10.6151
R2611 B.n337 B.n180 10.6151
R2612 B.n335 B.n334 10.6151
R2613 B.n334 B.n184 10.6151
R2614 B.n328 B.n184 10.6151
R2615 B.n328 B.n327 10.6151
R2616 B.n327 B.n326 10.6151
R2617 B.n326 B.n186 10.6151
R2618 B.n320 B.n186 10.6151
R2619 B.n320 B.n319 10.6151
R2620 B.n319 B.n318 10.6151
R2621 B.n318 B.n188 10.6151
R2622 B.n312 B.n188 10.6151
R2623 B.n312 B.n311 10.6151
R2624 B.n311 B.n310 10.6151
R2625 B.n310 B.n190 10.6151
R2626 B.n304 B.n190 10.6151
R2627 B.n304 B.n303 10.6151
R2628 B.n303 B.n302 10.6151
R2629 B.n302 B.n192 10.6151
R2630 B.n296 B.n192 10.6151
R2631 B.n296 B.n295 10.6151
R2632 B.n295 B.n294 10.6151
R2633 B.n294 B.n194 10.6151
R2634 B.n288 B.n194 10.6151
R2635 B.n288 B.n287 10.6151
R2636 B.n287 B.n286 10.6151
R2637 B.n286 B.n196 10.6151
R2638 B.n280 B.n196 10.6151
R2639 B.n280 B.n279 10.6151
R2640 B.n279 B.n278 10.6151
R2641 B.n278 B.n198 10.6151
R2642 B.n272 B.n198 10.6151
R2643 B.n272 B.n271 10.6151
R2644 B.n271 B.n270 10.6151
R2645 B.n270 B.n200 10.6151
R2646 B.n264 B.n200 10.6151
R2647 B.n264 B.n263 10.6151
R2648 B.n263 B.n262 10.6151
R2649 B.n262 B.n202 10.6151
R2650 B.n256 B.n202 10.6151
R2651 B.n256 B.n255 10.6151
R2652 B.n255 B.n254 10.6151
R2653 B.n254 B.n204 10.6151
R2654 B.n248 B.n204 10.6151
R2655 B.n248 B.n247 10.6151
R2656 B.n247 B.n246 10.6151
R2657 B.n246 B.n206 10.6151
R2658 B.n240 B.n206 10.6151
R2659 B.n240 B.n239 10.6151
R2660 B.n239 B.n238 10.6151
R2661 B.n238 B.n208 10.6151
R2662 B.n232 B.n208 10.6151
R2663 B.n232 B.n231 10.6151
R2664 B.n231 B.n230 10.6151
R2665 B.n230 B.n210 10.6151
R2666 B.n224 B.n210 10.6151
R2667 B.n224 B.n223 10.6151
R2668 B.n223 B.n222 10.6151
R2669 B.n222 B.n212 10.6151
R2670 B.n216 B.n212 10.6151
R2671 B.n216 B.n215 10.6151
R2672 B.n215 B.n139 10.6151
R2673 B.n478 B.n135 10.6151
R2674 B.n488 B.n135 10.6151
R2675 B.n489 B.n488 10.6151
R2676 B.n490 B.n489 10.6151
R2677 B.n490 B.n127 10.6151
R2678 B.n500 B.n127 10.6151
R2679 B.n501 B.n500 10.6151
R2680 B.n502 B.n501 10.6151
R2681 B.n502 B.n119 10.6151
R2682 B.n513 B.n119 10.6151
R2683 B.n514 B.n513 10.6151
R2684 B.n515 B.n514 10.6151
R2685 B.n515 B.n112 10.6151
R2686 B.n526 B.n112 10.6151
R2687 B.n527 B.n526 10.6151
R2688 B.n528 B.n527 10.6151
R2689 B.n528 B.n0 10.6151
R2690 B.n856 B.n1 10.6151
R2691 B.n856 B.n855 10.6151
R2692 B.n855 B.n854 10.6151
R2693 B.n854 B.n10 10.6151
R2694 B.n848 B.n10 10.6151
R2695 B.n848 B.n847 10.6151
R2696 B.n847 B.n846 10.6151
R2697 B.n846 B.n16 10.6151
R2698 B.n840 B.n16 10.6151
R2699 B.n840 B.n839 10.6151
R2700 B.n839 B.n838 10.6151
R2701 B.n838 B.n24 10.6151
R2702 B.n832 B.n24 10.6151
R2703 B.n832 B.n831 10.6151
R2704 B.n831 B.n830 10.6151
R2705 B.n830 B.n31 10.6151
R2706 B.n824 B.n31 10.6151
R2707 B.n510 B.t0 10.0233
R2708 B.n18 B.t1 10.0233
R2709 B.t3 B.n110 9.11212
R2710 B.t2 B.n8 9.11212
R2711 B.t5 B.n129 8.20096
R2712 B.n835 B.t12 8.20096
R2713 B.n698 B.n70 6.5566
R2714 B.n683 B.n682 6.5566
R2715 B.n353 B.n177 6.5566
R2716 B.n337 B.n336 6.5566
R2717 B.n702 B.n70 4.05904
R2718 B.n682 B.n681 4.05904
R2719 B.n177 B.n173 4.05904
R2720 B.n336 B.n335 4.05904
R2721 B.n862 B.n0 2.81026
R2722 B.n862 B.n1 2.81026
R2723 VP.n1 VP.t3 623.79
R2724 VP.n1 VP.t1 623.74
R2725 VP.n3 VP.t2 602.794
R2726 VP.n5 VP.t0 602.794
R2727 VP.n6 VP.n5 161.3
R2728 VP.n4 VP.n0 161.3
R2729 VP.n3 VP.n2 161.3
R2730 VP.n2 VP.n1 90.7303
R2731 VP.n4 VP.n3 24.1005
R2732 VP.n5 VP.n4 24.1005
R2733 VP.n2 VP.n0 0.189894
R2734 VP.n6 VP.n0 0.189894
R2735 VP VP.n6 0.0516364
R2736 VDD1 VDD1.n1 102.358
R2737 VDD1 VDD1.n0 58.9345
R2738 VDD1.n0 VDD1.t0 1.04978
R2739 VDD1.n0 VDD1.t2 1.04978
R2740 VDD1.n1 VDD1.t1 1.04978
R2741 VDD1.n1 VDD1.t3 1.04978
C0 VDD1 VDD2 0.594122f
C1 VP VDD1 5.29417f
C2 VN VTAIL 4.51273f
C3 VN VDD2 5.16081f
C4 VN VP 6.17879f
C5 VTAIL VDD2 9.27675f
C6 VTAIL VP 4.52683f
C7 VN VDD1 0.147199f
C8 VTAIL VDD1 9.23448f
C9 VP VDD2 0.280849f
C10 VDD2 B 3.304307f
C11 VDD1 B 7.76201f
C12 VTAIL B 12.8129f
C13 VN B 9.24083f
C14 VP B 5.613331f
C15 VDD1.t0 B 0.413685f
C16 VDD1.t2 B 0.413685f
C17 VDD1.n0 B 3.77272f
C18 VDD1.t1 B 0.413685f
C19 VDD1.t3 B 0.413685f
C20 VDD1.n1 B 4.68387f
C21 VP.n0 B 0.046719f
C22 VP.t1 B 2.07458f
C23 VP.t3 B 2.07465f
C24 VP.n1 B 2.67761f
C25 VP.n2 B 3.43098f
C26 VP.t2 B 2.04883f
C27 VP.n3 B 0.763469f
C28 VP.n4 B 0.010602f
C29 VP.t0 B 2.04883f
C30 VP.n5 B 0.763469f
C31 VP.n6 B 0.036206f
C32 VTAIL.n0 B 0.021215f
C33 VTAIL.n1 B 0.015464f
C34 VTAIL.n2 B 0.00831f
C35 VTAIL.n3 B 0.019641f
C36 VTAIL.n4 B 0.008799f
C37 VTAIL.n5 B 0.015464f
C38 VTAIL.n6 B 0.00831f
C39 VTAIL.n7 B 0.019641f
C40 VTAIL.n8 B 0.008799f
C41 VTAIL.n9 B 0.015464f
C42 VTAIL.n10 B 0.00831f
C43 VTAIL.n11 B 0.019641f
C44 VTAIL.n12 B 0.008799f
C45 VTAIL.n13 B 0.015464f
C46 VTAIL.n14 B 0.00831f
C47 VTAIL.n15 B 0.019641f
C48 VTAIL.n16 B 0.008799f
C49 VTAIL.n17 B 0.015464f
C50 VTAIL.n18 B 0.00831f
C51 VTAIL.n19 B 0.019641f
C52 VTAIL.n20 B 0.008799f
C53 VTAIL.n21 B 0.015464f
C54 VTAIL.n22 B 0.00831f
C55 VTAIL.n23 B 0.019641f
C56 VTAIL.n24 B 0.008799f
C57 VTAIL.n25 B 0.015464f
C58 VTAIL.n26 B 0.00831f
C59 VTAIL.n27 B 0.019641f
C60 VTAIL.n28 B 0.008799f
C61 VTAIL.n29 B 0.015464f
C62 VTAIL.n30 B 0.00831f
C63 VTAIL.n31 B 0.019641f
C64 VTAIL.n32 B 0.008799f
C65 VTAIL.n33 B 0.115865f
C66 VTAIL.t7 B 0.032591f
C67 VTAIL.n34 B 0.014731f
C68 VTAIL.n35 B 0.011603f
C69 VTAIL.n36 B 0.00831f
C70 VTAIL.n37 B 1.28039f
C71 VTAIL.n38 B 0.015464f
C72 VTAIL.n39 B 0.00831f
C73 VTAIL.n40 B 0.008799f
C74 VTAIL.n41 B 0.019641f
C75 VTAIL.n42 B 0.019641f
C76 VTAIL.n43 B 0.008799f
C77 VTAIL.n44 B 0.00831f
C78 VTAIL.n45 B 0.015464f
C79 VTAIL.n46 B 0.015464f
C80 VTAIL.n47 B 0.00831f
C81 VTAIL.n48 B 0.008799f
C82 VTAIL.n49 B 0.019641f
C83 VTAIL.n50 B 0.019641f
C84 VTAIL.n51 B 0.008799f
C85 VTAIL.n52 B 0.00831f
C86 VTAIL.n53 B 0.015464f
C87 VTAIL.n54 B 0.015464f
C88 VTAIL.n55 B 0.00831f
C89 VTAIL.n56 B 0.008799f
C90 VTAIL.n57 B 0.019641f
C91 VTAIL.n58 B 0.019641f
C92 VTAIL.n59 B 0.008799f
C93 VTAIL.n60 B 0.00831f
C94 VTAIL.n61 B 0.015464f
C95 VTAIL.n62 B 0.015464f
C96 VTAIL.n63 B 0.00831f
C97 VTAIL.n64 B 0.008799f
C98 VTAIL.n65 B 0.019641f
C99 VTAIL.n66 B 0.019641f
C100 VTAIL.n67 B 0.008799f
C101 VTAIL.n68 B 0.00831f
C102 VTAIL.n69 B 0.015464f
C103 VTAIL.n70 B 0.015464f
C104 VTAIL.n71 B 0.00831f
C105 VTAIL.n72 B 0.008799f
C106 VTAIL.n73 B 0.019641f
C107 VTAIL.n74 B 0.019641f
C108 VTAIL.n75 B 0.019641f
C109 VTAIL.n76 B 0.008799f
C110 VTAIL.n77 B 0.00831f
C111 VTAIL.n78 B 0.015464f
C112 VTAIL.n79 B 0.015464f
C113 VTAIL.n80 B 0.00831f
C114 VTAIL.n81 B 0.008554f
C115 VTAIL.n82 B 0.008554f
C116 VTAIL.n83 B 0.019641f
C117 VTAIL.n84 B 0.019641f
C118 VTAIL.n85 B 0.008799f
C119 VTAIL.n86 B 0.00831f
C120 VTAIL.n87 B 0.015464f
C121 VTAIL.n88 B 0.015464f
C122 VTAIL.n89 B 0.00831f
C123 VTAIL.n90 B 0.008799f
C124 VTAIL.n91 B 0.019641f
C125 VTAIL.n92 B 0.019641f
C126 VTAIL.n93 B 0.008799f
C127 VTAIL.n94 B 0.00831f
C128 VTAIL.n95 B 0.015464f
C129 VTAIL.n96 B 0.015464f
C130 VTAIL.n97 B 0.00831f
C131 VTAIL.n98 B 0.008799f
C132 VTAIL.n99 B 0.019641f
C133 VTAIL.n100 B 0.041597f
C134 VTAIL.n101 B 0.008799f
C135 VTAIL.n102 B 0.00831f
C136 VTAIL.n103 B 0.033843f
C137 VTAIL.n104 B 0.023121f
C138 VTAIL.n105 B 0.063146f
C139 VTAIL.n106 B 0.021215f
C140 VTAIL.n107 B 0.015464f
C141 VTAIL.n108 B 0.00831f
C142 VTAIL.n109 B 0.019641f
C143 VTAIL.n110 B 0.008799f
C144 VTAIL.n111 B 0.015464f
C145 VTAIL.n112 B 0.00831f
C146 VTAIL.n113 B 0.019641f
C147 VTAIL.n114 B 0.008799f
C148 VTAIL.n115 B 0.015464f
C149 VTAIL.n116 B 0.00831f
C150 VTAIL.n117 B 0.019641f
C151 VTAIL.n118 B 0.008799f
C152 VTAIL.n119 B 0.015464f
C153 VTAIL.n120 B 0.00831f
C154 VTAIL.n121 B 0.019641f
C155 VTAIL.n122 B 0.008799f
C156 VTAIL.n123 B 0.015464f
C157 VTAIL.n124 B 0.00831f
C158 VTAIL.n125 B 0.019641f
C159 VTAIL.n126 B 0.008799f
C160 VTAIL.n127 B 0.015464f
C161 VTAIL.n128 B 0.00831f
C162 VTAIL.n129 B 0.019641f
C163 VTAIL.n130 B 0.008799f
C164 VTAIL.n131 B 0.015464f
C165 VTAIL.n132 B 0.00831f
C166 VTAIL.n133 B 0.019641f
C167 VTAIL.n134 B 0.008799f
C168 VTAIL.n135 B 0.015464f
C169 VTAIL.n136 B 0.00831f
C170 VTAIL.n137 B 0.019641f
C171 VTAIL.n138 B 0.008799f
C172 VTAIL.n139 B 0.115865f
C173 VTAIL.t3 B 0.032591f
C174 VTAIL.n140 B 0.014731f
C175 VTAIL.n141 B 0.011603f
C176 VTAIL.n142 B 0.00831f
C177 VTAIL.n143 B 1.28039f
C178 VTAIL.n144 B 0.015464f
C179 VTAIL.n145 B 0.00831f
C180 VTAIL.n146 B 0.008799f
C181 VTAIL.n147 B 0.019641f
C182 VTAIL.n148 B 0.019641f
C183 VTAIL.n149 B 0.008799f
C184 VTAIL.n150 B 0.00831f
C185 VTAIL.n151 B 0.015464f
C186 VTAIL.n152 B 0.015464f
C187 VTAIL.n153 B 0.00831f
C188 VTAIL.n154 B 0.008799f
C189 VTAIL.n155 B 0.019641f
C190 VTAIL.n156 B 0.019641f
C191 VTAIL.n157 B 0.008799f
C192 VTAIL.n158 B 0.00831f
C193 VTAIL.n159 B 0.015464f
C194 VTAIL.n160 B 0.015464f
C195 VTAIL.n161 B 0.00831f
C196 VTAIL.n162 B 0.008799f
C197 VTAIL.n163 B 0.019641f
C198 VTAIL.n164 B 0.019641f
C199 VTAIL.n165 B 0.008799f
C200 VTAIL.n166 B 0.00831f
C201 VTAIL.n167 B 0.015464f
C202 VTAIL.n168 B 0.015464f
C203 VTAIL.n169 B 0.00831f
C204 VTAIL.n170 B 0.008799f
C205 VTAIL.n171 B 0.019641f
C206 VTAIL.n172 B 0.019641f
C207 VTAIL.n173 B 0.008799f
C208 VTAIL.n174 B 0.00831f
C209 VTAIL.n175 B 0.015464f
C210 VTAIL.n176 B 0.015464f
C211 VTAIL.n177 B 0.00831f
C212 VTAIL.n178 B 0.008799f
C213 VTAIL.n179 B 0.019641f
C214 VTAIL.n180 B 0.019641f
C215 VTAIL.n181 B 0.019641f
C216 VTAIL.n182 B 0.008799f
C217 VTAIL.n183 B 0.00831f
C218 VTAIL.n184 B 0.015464f
C219 VTAIL.n185 B 0.015464f
C220 VTAIL.n186 B 0.00831f
C221 VTAIL.n187 B 0.008554f
C222 VTAIL.n188 B 0.008554f
C223 VTAIL.n189 B 0.019641f
C224 VTAIL.n190 B 0.019641f
C225 VTAIL.n191 B 0.008799f
C226 VTAIL.n192 B 0.00831f
C227 VTAIL.n193 B 0.015464f
C228 VTAIL.n194 B 0.015464f
C229 VTAIL.n195 B 0.00831f
C230 VTAIL.n196 B 0.008799f
C231 VTAIL.n197 B 0.019641f
C232 VTAIL.n198 B 0.019641f
C233 VTAIL.n199 B 0.008799f
C234 VTAIL.n200 B 0.00831f
C235 VTAIL.n201 B 0.015464f
C236 VTAIL.n202 B 0.015464f
C237 VTAIL.n203 B 0.00831f
C238 VTAIL.n204 B 0.008799f
C239 VTAIL.n205 B 0.019641f
C240 VTAIL.n206 B 0.041597f
C241 VTAIL.n207 B 0.008799f
C242 VTAIL.n208 B 0.00831f
C243 VTAIL.n209 B 0.033843f
C244 VTAIL.n210 B 0.023121f
C245 VTAIL.n211 B 0.084946f
C246 VTAIL.n212 B 0.021215f
C247 VTAIL.n213 B 0.015464f
C248 VTAIL.n214 B 0.00831f
C249 VTAIL.n215 B 0.019641f
C250 VTAIL.n216 B 0.008799f
C251 VTAIL.n217 B 0.015464f
C252 VTAIL.n218 B 0.00831f
C253 VTAIL.n219 B 0.019641f
C254 VTAIL.n220 B 0.008799f
C255 VTAIL.n221 B 0.015464f
C256 VTAIL.n222 B 0.00831f
C257 VTAIL.n223 B 0.019641f
C258 VTAIL.n224 B 0.008799f
C259 VTAIL.n225 B 0.015464f
C260 VTAIL.n226 B 0.00831f
C261 VTAIL.n227 B 0.019641f
C262 VTAIL.n228 B 0.008799f
C263 VTAIL.n229 B 0.015464f
C264 VTAIL.n230 B 0.00831f
C265 VTAIL.n231 B 0.019641f
C266 VTAIL.n232 B 0.008799f
C267 VTAIL.n233 B 0.015464f
C268 VTAIL.n234 B 0.00831f
C269 VTAIL.n235 B 0.019641f
C270 VTAIL.n236 B 0.008799f
C271 VTAIL.n237 B 0.015464f
C272 VTAIL.n238 B 0.00831f
C273 VTAIL.n239 B 0.019641f
C274 VTAIL.n240 B 0.008799f
C275 VTAIL.n241 B 0.015464f
C276 VTAIL.n242 B 0.00831f
C277 VTAIL.n243 B 0.019641f
C278 VTAIL.n244 B 0.008799f
C279 VTAIL.n245 B 0.115865f
C280 VTAIL.t0 B 0.032591f
C281 VTAIL.n246 B 0.014731f
C282 VTAIL.n247 B 0.011603f
C283 VTAIL.n248 B 0.00831f
C284 VTAIL.n249 B 1.28039f
C285 VTAIL.n250 B 0.015464f
C286 VTAIL.n251 B 0.00831f
C287 VTAIL.n252 B 0.008799f
C288 VTAIL.n253 B 0.019641f
C289 VTAIL.n254 B 0.019641f
C290 VTAIL.n255 B 0.008799f
C291 VTAIL.n256 B 0.00831f
C292 VTAIL.n257 B 0.015464f
C293 VTAIL.n258 B 0.015464f
C294 VTAIL.n259 B 0.00831f
C295 VTAIL.n260 B 0.008799f
C296 VTAIL.n261 B 0.019641f
C297 VTAIL.n262 B 0.019641f
C298 VTAIL.n263 B 0.008799f
C299 VTAIL.n264 B 0.00831f
C300 VTAIL.n265 B 0.015464f
C301 VTAIL.n266 B 0.015464f
C302 VTAIL.n267 B 0.00831f
C303 VTAIL.n268 B 0.008799f
C304 VTAIL.n269 B 0.019641f
C305 VTAIL.n270 B 0.019641f
C306 VTAIL.n271 B 0.008799f
C307 VTAIL.n272 B 0.00831f
C308 VTAIL.n273 B 0.015464f
C309 VTAIL.n274 B 0.015464f
C310 VTAIL.n275 B 0.00831f
C311 VTAIL.n276 B 0.008799f
C312 VTAIL.n277 B 0.019641f
C313 VTAIL.n278 B 0.019641f
C314 VTAIL.n279 B 0.008799f
C315 VTAIL.n280 B 0.00831f
C316 VTAIL.n281 B 0.015464f
C317 VTAIL.n282 B 0.015464f
C318 VTAIL.n283 B 0.00831f
C319 VTAIL.n284 B 0.008799f
C320 VTAIL.n285 B 0.019641f
C321 VTAIL.n286 B 0.019641f
C322 VTAIL.n287 B 0.019641f
C323 VTAIL.n288 B 0.008799f
C324 VTAIL.n289 B 0.00831f
C325 VTAIL.n290 B 0.015464f
C326 VTAIL.n291 B 0.015464f
C327 VTAIL.n292 B 0.00831f
C328 VTAIL.n293 B 0.008554f
C329 VTAIL.n294 B 0.008554f
C330 VTAIL.n295 B 0.019641f
C331 VTAIL.n296 B 0.019641f
C332 VTAIL.n297 B 0.008799f
C333 VTAIL.n298 B 0.00831f
C334 VTAIL.n299 B 0.015464f
C335 VTAIL.n300 B 0.015464f
C336 VTAIL.n301 B 0.00831f
C337 VTAIL.n302 B 0.008799f
C338 VTAIL.n303 B 0.019641f
C339 VTAIL.n304 B 0.019641f
C340 VTAIL.n305 B 0.008799f
C341 VTAIL.n306 B 0.00831f
C342 VTAIL.n307 B 0.015464f
C343 VTAIL.n308 B 0.015464f
C344 VTAIL.n309 B 0.00831f
C345 VTAIL.n310 B 0.008799f
C346 VTAIL.n311 B 0.019641f
C347 VTAIL.n312 B 0.041597f
C348 VTAIL.n313 B 0.008799f
C349 VTAIL.n314 B 0.00831f
C350 VTAIL.n315 B 0.033843f
C351 VTAIL.n316 B 0.023121f
C352 VTAIL.n317 B 1.13157f
C353 VTAIL.n318 B 0.021215f
C354 VTAIL.n319 B 0.015464f
C355 VTAIL.n320 B 0.00831f
C356 VTAIL.n321 B 0.019641f
C357 VTAIL.n322 B 0.008799f
C358 VTAIL.n323 B 0.015464f
C359 VTAIL.n324 B 0.00831f
C360 VTAIL.n325 B 0.019641f
C361 VTAIL.n326 B 0.008799f
C362 VTAIL.n327 B 0.015464f
C363 VTAIL.n328 B 0.00831f
C364 VTAIL.n329 B 0.019641f
C365 VTAIL.n330 B 0.008799f
C366 VTAIL.n331 B 0.015464f
C367 VTAIL.n332 B 0.00831f
C368 VTAIL.n333 B 0.019641f
C369 VTAIL.n334 B 0.019641f
C370 VTAIL.n335 B 0.008799f
C371 VTAIL.n336 B 0.015464f
C372 VTAIL.n337 B 0.00831f
C373 VTAIL.n338 B 0.019641f
C374 VTAIL.n339 B 0.008799f
C375 VTAIL.n340 B 0.015464f
C376 VTAIL.n341 B 0.00831f
C377 VTAIL.n342 B 0.019641f
C378 VTAIL.n343 B 0.008799f
C379 VTAIL.n344 B 0.015464f
C380 VTAIL.n345 B 0.00831f
C381 VTAIL.n346 B 0.019641f
C382 VTAIL.n347 B 0.008799f
C383 VTAIL.n348 B 0.015464f
C384 VTAIL.n349 B 0.00831f
C385 VTAIL.n350 B 0.019641f
C386 VTAIL.n351 B 0.008799f
C387 VTAIL.n352 B 0.115865f
C388 VTAIL.t5 B 0.032591f
C389 VTAIL.n353 B 0.014731f
C390 VTAIL.n354 B 0.011603f
C391 VTAIL.n355 B 0.00831f
C392 VTAIL.n356 B 1.28039f
C393 VTAIL.n357 B 0.015464f
C394 VTAIL.n358 B 0.00831f
C395 VTAIL.n359 B 0.008799f
C396 VTAIL.n360 B 0.019641f
C397 VTAIL.n361 B 0.019641f
C398 VTAIL.n362 B 0.008799f
C399 VTAIL.n363 B 0.00831f
C400 VTAIL.n364 B 0.015464f
C401 VTAIL.n365 B 0.015464f
C402 VTAIL.n366 B 0.00831f
C403 VTAIL.n367 B 0.008799f
C404 VTAIL.n368 B 0.019641f
C405 VTAIL.n369 B 0.019641f
C406 VTAIL.n370 B 0.008799f
C407 VTAIL.n371 B 0.00831f
C408 VTAIL.n372 B 0.015464f
C409 VTAIL.n373 B 0.015464f
C410 VTAIL.n374 B 0.00831f
C411 VTAIL.n375 B 0.008799f
C412 VTAIL.n376 B 0.019641f
C413 VTAIL.n377 B 0.019641f
C414 VTAIL.n378 B 0.008799f
C415 VTAIL.n379 B 0.00831f
C416 VTAIL.n380 B 0.015464f
C417 VTAIL.n381 B 0.015464f
C418 VTAIL.n382 B 0.00831f
C419 VTAIL.n383 B 0.008799f
C420 VTAIL.n384 B 0.019641f
C421 VTAIL.n385 B 0.019641f
C422 VTAIL.n386 B 0.008799f
C423 VTAIL.n387 B 0.00831f
C424 VTAIL.n388 B 0.015464f
C425 VTAIL.n389 B 0.015464f
C426 VTAIL.n390 B 0.00831f
C427 VTAIL.n391 B 0.008799f
C428 VTAIL.n392 B 0.019641f
C429 VTAIL.n393 B 0.019641f
C430 VTAIL.n394 B 0.008799f
C431 VTAIL.n395 B 0.00831f
C432 VTAIL.n396 B 0.015464f
C433 VTAIL.n397 B 0.015464f
C434 VTAIL.n398 B 0.00831f
C435 VTAIL.n399 B 0.008554f
C436 VTAIL.n400 B 0.008554f
C437 VTAIL.n401 B 0.019641f
C438 VTAIL.n402 B 0.019641f
C439 VTAIL.n403 B 0.008799f
C440 VTAIL.n404 B 0.00831f
C441 VTAIL.n405 B 0.015464f
C442 VTAIL.n406 B 0.015464f
C443 VTAIL.n407 B 0.00831f
C444 VTAIL.n408 B 0.008799f
C445 VTAIL.n409 B 0.019641f
C446 VTAIL.n410 B 0.019641f
C447 VTAIL.n411 B 0.008799f
C448 VTAIL.n412 B 0.00831f
C449 VTAIL.n413 B 0.015464f
C450 VTAIL.n414 B 0.015464f
C451 VTAIL.n415 B 0.00831f
C452 VTAIL.n416 B 0.008799f
C453 VTAIL.n417 B 0.019641f
C454 VTAIL.n418 B 0.041597f
C455 VTAIL.n419 B 0.008799f
C456 VTAIL.n420 B 0.00831f
C457 VTAIL.n421 B 0.033843f
C458 VTAIL.n422 B 0.023121f
C459 VTAIL.n423 B 1.13157f
C460 VTAIL.n424 B 0.021215f
C461 VTAIL.n425 B 0.015464f
C462 VTAIL.n426 B 0.00831f
C463 VTAIL.n427 B 0.019641f
C464 VTAIL.n428 B 0.008799f
C465 VTAIL.n429 B 0.015464f
C466 VTAIL.n430 B 0.00831f
C467 VTAIL.n431 B 0.019641f
C468 VTAIL.n432 B 0.008799f
C469 VTAIL.n433 B 0.015464f
C470 VTAIL.n434 B 0.00831f
C471 VTAIL.n435 B 0.019641f
C472 VTAIL.n436 B 0.008799f
C473 VTAIL.n437 B 0.015464f
C474 VTAIL.n438 B 0.00831f
C475 VTAIL.n439 B 0.019641f
C476 VTAIL.n440 B 0.019641f
C477 VTAIL.n441 B 0.008799f
C478 VTAIL.n442 B 0.015464f
C479 VTAIL.n443 B 0.00831f
C480 VTAIL.n444 B 0.019641f
C481 VTAIL.n445 B 0.008799f
C482 VTAIL.n446 B 0.015464f
C483 VTAIL.n447 B 0.00831f
C484 VTAIL.n448 B 0.019641f
C485 VTAIL.n449 B 0.008799f
C486 VTAIL.n450 B 0.015464f
C487 VTAIL.n451 B 0.00831f
C488 VTAIL.n452 B 0.019641f
C489 VTAIL.n453 B 0.008799f
C490 VTAIL.n454 B 0.015464f
C491 VTAIL.n455 B 0.00831f
C492 VTAIL.n456 B 0.019641f
C493 VTAIL.n457 B 0.008799f
C494 VTAIL.n458 B 0.115865f
C495 VTAIL.t4 B 0.032591f
C496 VTAIL.n459 B 0.014731f
C497 VTAIL.n460 B 0.011603f
C498 VTAIL.n461 B 0.00831f
C499 VTAIL.n462 B 1.28039f
C500 VTAIL.n463 B 0.015464f
C501 VTAIL.n464 B 0.00831f
C502 VTAIL.n465 B 0.008799f
C503 VTAIL.n466 B 0.019641f
C504 VTAIL.n467 B 0.019641f
C505 VTAIL.n468 B 0.008799f
C506 VTAIL.n469 B 0.00831f
C507 VTAIL.n470 B 0.015464f
C508 VTAIL.n471 B 0.015464f
C509 VTAIL.n472 B 0.00831f
C510 VTAIL.n473 B 0.008799f
C511 VTAIL.n474 B 0.019641f
C512 VTAIL.n475 B 0.019641f
C513 VTAIL.n476 B 0.008799f
C514 VTAIL.n477 B 0.00831f
C515 VTAIL.n478 B 0.015464f
C516 VTAIL.n479 B 0.015464f
C517 VTAIL.n480 B 0.00831f
C518 VTAIL.n481 B 0.008799f
C519 VTAIL.n482 B 0.019641f
C520 VTAIL.n483 B 0.019641f
C521 VTAIL.n484 B 0.008799f
C522 VTAIL.n485 B 0.00831f
C523 VTAIL.n486 B 0.015464f
C524 VTAIL.n487 B 0.015464f
C525 VTAIL.n488 B 0.00831f
C526 VTAIL.n489 B 0.008799f
C527 VTAIL.n490 B 0.019641f
C528 VTAIL.n491 B 0.019641f
C529 VTAIL.n492 B 0.008799f
C530 VTAIL.n493 B 0.00831f
C531 VTAIL.n494 B 0.015464f
C532 VTAIL.n495 B 0.015464f
C533 VTAIL.n496 B 0.00831f
C534 VTAIL.n497 B 0.008799f
C535 VTAIL.n498 B 0.019641f
C536 VTAIL.n499 B 0.019641f
C537 VTAIL.n500 B 0.008799f
C538 VTAIL.n501 B 0.00831f
C539 VTAIL.n502 B 0.015464f
C540 VTAIL.n503 B 0.015464f
C541 VTAIL.n504 B 0.00831f
C542 VTAIL.n505 B 0.008554f
C543 VTAIL.n506 B 0.008554f
C544 VTAIL.n507 B 0.019641f
C545 VTAIL.n508 B 0.019641f
C546 VTAIL.n509 B 0.008799f
C547 VTAIL.n510 B 0.00831f
C548 VTAIL.n511 B 0.015464f
C549 VTAIL.n512 B 0.015464f
C550 VTAIL.n513 B 0.00831f
C551 VTAIL.n514 B 0.008799f
C552 VTAIL.n515 B 0.019641f
C553 VTAIL.n516 B 0.019641f
C554 VTAIL.n517 B 0.008799f
C555 VTAIL.n518 B 0.00831f
C556 VTAIL.n519 B 0.015464f
C557 VTAIL.n520 B 0.015464f
C558 VTAIL.n521 B 0.00831f
C559 VTAIL.n522 B 0.008799f
C560 VTAIL.n523 B 0.019641f
C561 VTAIL.n524 B 0.041597f
C562 VTAIL.n525 B 0.008799f
C563 VTAIL.n526 B 0.00831f
C564 VTAIL.n527 B 0.033843f
C565 VTAIL.n528 B 0.023121f
C566 VTAIL.n529 B 0.084946f
C567 VTAIL.n530 B 0.021215f
C568 VTAIL.n531 B 0.015464f
C569 VTAIL.n532 B 0.00831f
C570 VTAIL.n533 B 0.019641f
C571 VTAIL.n534 B 0.008799f
C572 VTAIL.n535 B 0.015464f
C573 VTAIL.n536 B 0.00831f
C574 VTAIL.n537 B 0.019641f
C575 VTAIL.n538 B 0.008799f
C576 VTAIL.n539 B 0.015464f
C577 VTAIL.n540 B 0.00831f
C578 VTAIL.n541 B 0.019641f
C579 VTAIL.n542 B 0.008799f
C580 VTAIL.n543 B 0.015464f
C581 VTAIL.n544 B 0.00831f
C582 VTAIL.n545 B 0.019641f
C583 VTAIL.n546 B 0.019641f
C584 VTAIL.n547 B 0.008799f
C585 VTAIL.n548 B 0.015464f
C586 VTAIL.n549 B 0.00831f
C587 VTAIL.n550 B 0.019641f
C588 VTAIL.n551 B 0.008799f
C589 VTAIL.n552 B 0.015464f
C590 VTAIL.n553 B 0.00831f
C591 VTAIL.n554 B 0.019641f
C592 VTAIL.n555 B 0.008799f
C593 VTAIL.n556 B 0.015464f
C594 VTAIL.n557 B 0.00831f
C595 VTAIL.n558 B 0.019641f
C596 VTAIL.n559 B 0.008799f
C597 VTAIL.n560 B 0.015464f
C598 VTAIL.n561 B 0.00831f
C599 VTAIL.n562 B 0.019641f
C600 VTAIL.n563 B 0.008799f
C601 VTAIL.n564 B 0.115865f
C602 VTAIL.t2 B 0.032591f
C603 VTAIL.n565 B 0.014731f
C604 VTAIL.n566 B 0.011603f
C605 VTAIL.n567 B 0.00831f
C606 VTAIL.n568 B 1.28039f
C607 VTAIL.n569 B 0.015464f
C608 VTAIL.n570 B 0.00831f
C609 VTAIL.n571 B 0.008799f
C610 VTAIL.n572 B 0.019641f
C611 VTAIL.n573 B 0.019641f
C612 VTAIL.n574 B 0.008799f
C613 VTAIL.n575 B 0.00831f
C614 VTAIL.n576 B 0.015464f
C615 VTAIL.n577 B 0.015464f
C616 VTAIL.n578 B 0.00831f
C617 VTAIL.n579 B 0.008799f
C618 VTAIL.n580 B 0.019641f
C619 VTAIL.n581 B 0.019641f
C620 VTAIL.n582 B 0.008799f
C621 VTAIL.n583 B 0.00831f
C622 VTAIL.n584 B 0.015464f
C623 VTAIL.n585 B 0.015464f
C624 VTAIL.n586 B 0.00831f
C625 VTAIL.n587 B 0.008799f
C626 VTAIL.n588 B 0.019641f
C627 VTAIL.n589 B 0.019641f
C628 VTAIL.n590 B 0.008799f
C629 VTAIL.n591 B 0.00831f
C630 VTAIL.n592 B 0.015464f
C631 VTAIL.n593 B 0.015464f
C632 VTAIL.n594 B 0.00831f
C633 VTAIL.n595 B 0.008799f
C634 VTAIL.n596 B 0.019641f
C635 VTAIL.n597 B 0.019641f
C636 VTAIL.n598 B 0.008799f
C637 VTAIL.n599 B 0.00831f
C638 VTAIL.n600 B 0.015464f
C639 VTAIL.n601 B 0.015464f
C640 VTAIL.n602 B 0.00831f
C641 VTAIL.n603 B 0.008799f
C642 VTAIL.n604 B 0.019641f
C643 VTAIL.n605 B 0.019641f
C644 VTAIL.n606 B 0.008799f
C645 VTAIL.n607 B 0.00831f
C646 VTAIL.n608 B 0.015464f
C647 VTAIL.n609 B 0.015464f
C648 VTAIL.n610 B 0.00831f
C649 VTAIL.n611 B 0.008554f
C650 VTAIL.n612 B 0.008554f
C651 VTAIL.n613 B 0.019641f
C652 VTAIL.n614 B 0.019641f
C653 VTAIL.n615 B 0.008799f
C654 VTAIL.n616 B 0.00831f
C655 VTAIL.n617 B 0.015464f
C656 VTAIL.n618 B 0.015464f
C657 VTAIL.n619 B 0.00831f
C658 VTAIL.n620 B 0.008799f
C659 VTAIL.n621 B 0.019641f
C660 VTAIL.n622 B 0.019641f
C661 VTAIL.n623 B 0.008799f
C662 VTAIL.n624 B 0.00831f
C663 VTAIL.n625 B 0.015464f
C664 VTAIL.n626 B 0.015464f
C665 VTAIL.n627 B 0.00831f
C666 VTAIL.n628 B 0.008799f
C667 VTAIL.n629 B 0.019641f
C668 VTAIL.n630 B 0.041597f
C669 VTAIL.n631 B 0.008799f
C670 VTAIL.n632 B 0.00831f
C671 VTAIL.n633 B 0.033843f
C672 VTAIL.n634 B 0.023121f
C673 VTAIL.n635 B 0.084946f
C674 VTAIL.n636 B 0.021215f
C675 VTAIL.n637 B 0.015464f
C676 VTAIL.n638 B 0.00831f
C677 VTAIL.n639 B 0.019641f
C678 VTAIL.n640 B 0.008799f
C679 VTAIL.n641 B 0.015464f
C680 VTAIL.n642 B 0.00831f
C681 VTAIL.n643 B 0.019641f
C682 VTAIL.n644 B 0.008799f
C683 VTAIL.n645 B 0.015464f
C684 VTAIL.n646 B 0.00831f
C685 VTAIL.n647 B 0.019641f
C686 VTAIL.n648 B 0.008799f
C687 VTAIL.n649 B 0.015464f
C688 VTAIL.n650 B 0.00831f
C689 VTAIL.n651 B 0.019641f
C690 VTAIL.n652 B 0.019641f
C691 VTAIL.n653 B 0.008799f
C692 VTAIL.n654 B 0.015464f
C693 VTAIL.n655 B 0.00831f
C694 VTAIL.n656 B 0.019641f
C695 VTAIL.n657 B 0.008799f
C696 VTAIL.n658 B 0.015464f
C697 VTAIL.n659 B 0.00831f
C698 VTAIL.n660 B 0.019641f
C699 VTAIL.n661 B 0.008799f
C700 VTAIL.n662 B 0.015464f
C701 VTAIL.n663 B 0.00831f
C702 VTAIL.n664 B 0.019641f
C703 VTAIL.n665 B 0.008799f
C704 VTAIL.n666 B 0.015464f
C705 VTAIL.n667 B 0.00831f
C706 VTAIL.n668 B 0.019641f
C707 VTAIL.n669 B 0.008799f
C708 VTAIL.n670 B 0.115865f
C709 VTAIL.t1 B 0.032591f
C710 VTAIL.n671 B 0.014731f
C711 VTAIL.n672 B 0.011603f
C712 VTAIL.n673 B 0.00831f
C713 VTAIL.n674 B 1.28039f
C714 VTAIL.n675 B 0.015464f
C715 VTAIL.n676 B 0.00831f
C716 VTAIL.n677 B 0.008799f
C717 VTAIL.n678 B 0.019641f
C718 VTAIL.n679 B 0.019641f
C719 VTAIL.n680 B 0.008799f
C720 VTAIL.n681 B 0.00831f
C721 VTAIL.n682 B 0.015464f
C722 VTAIL.n683 B 0.015464f
C723 VTAIL.n684 B 0.00831f
C724 VTAIL.n685 B 0.008799f
C725 VTAIL.n686 B 0.019641f
C726 VTAIL.n687 B 0.019641f
C727 VTAIL.n688 B 0.008799f
C728 VTAIL.n689 B 0.00831f
C729 VTAIL.n690 B 0.015464f
C730 VTAIL.n691 B 0.015464f
C731 VTAIL.n692 B 0.00831f
C732 VTAIL.n693 B 0.008799f
C733 VTAIL.n694 B 0.019641f
C734 VTAIL.n695 B 0.019641f
C735 VTAIL.n696 B 0.008799f
C736 VTAIL.n697 B 0.00831f
C737 VTAIL.n698 B 0.015464f
C738 VTAIL.n699 B 0.015464f
C739 VTAIL.n700 B 0.00831f
C740 VTAIL.n701 B 0.008799f
C741 VTAIL.n702 B 0.019641f
C742 VTAIL.n703 B 0.019641f
C743 VTAIL.n704 B 0.008799f
C744 VTAIL.n705 B 0.00831f
C745 VTAIL.n706 B 0.015464f
C746 VTAIL.n707 B 0.015464f
C747 VTAIL.n708 B 0.00831f
C748 VTAIL.n709 B 0.008799f
C749 VTAIL.n710 B 0.019641f
C750 VTAIL.n711 B 0.019641f
C751 VTAIL.n712 B 0.008799f
C752 VTAIL.n713 B 0.00831f
C753 VTAIL.n714 B 0.015464f
C754 VTAIL.n715 B 0.015464f
C755 VTAIL.n716 B 0.00831f
C756 VTAIL.n717 B 0.008554f
C757 VTAIL.n718 B 0.008554f
C758 VTAIL.n719 B 0.019641f
C759 VTAIL.n720 B 0.019641f
C760 VTAIL.n721 B 0.008799f
C761 VTAIL.n722 B 0.00831f
C762 VTAIL.n723 B 0.015464f
C763 VTAIL.n724 B 0.015464f
C764 VTAIL.n725 B 0.00831f
C765 VTAIL.n726 B 0.008799f
C766 VTAIL.n727 B 0.019641f
C767 VTAIL.n728 B 0.019641f
C768 VTAIL.n729 B 0.008799f
C769 VTAIL.n730 B 0.00831f
C770 VTAIL.n731 B 0.015464f
C771 VTAIL.n732 B 0.015464f
C772 VTAIL.n733 B 0.00831f
C773 VTAIL.n734 B 0.008799f
C774 VTAIL.n735 B 0.019641f
C775 VTAIL.n736 B 0.041597f
C776 VTAIL.n737 B 0.008799f
C777 VTAIL.n738 B 0.00831f
C778 VTAIL.n739 B 0.033843f
C779 VTAIL.n740 B 0.023121f
C780 VTAIL.n741 B 1.13157f
C781 VTAIL.n742 B 0.021215f
C782 VTAIL.n743 B 0.015464f
C783 VTAIL.n744 B 0.00831f
C784 VTAIL.n745 B 0.019641f
C785 VTAIL.n746 B 0.008799f
C786 VTAIL.n747 B 0.015464f
C787 VTAIL.n748 B 0.00831f
C788 VTAIL.n749 B 0.019641f
C789 VTAIL.n750 B 0.008799f
C790 VTAIL.n751 B 0.015464f
C791 VTAIL.n752 B 0.00831f
C792 VTAIL.n753 B 0.019641f
C793 VTAIL.n754 B 0.008799f
C794 VTAIL.n755 B 0.015464f
C795 VTAIL.n756 B 0.00831f
C796 VTAIL.n757 B 0.019641f
C797 VTAIL.n758 B 0.008799f
C798 VTAIL.n759 B 0.015464f
C799 VTAIL.n760 B 0.00831f
C800 VTAIL.n761 B 0.019641f
C801 VTAIL.n762 B 0.008799f
C802 VTAIL.n763 B 0.015464f
C803 VTAIL.n764 B 0.00831f
C804 VTAIL.n765 B 0.019641f
C805 VTAIL.n766 B 0.008799f
C806 VTAIL.n767 B 0.015464f
C807 VTAIL.n768 B 0.00831f
C808 VTAIL.n769 B 0.019641f
C809 VTAIL.n770 B 0.008799f
C810 VTAIL.n771 B 0.015464f
C811 VTAIL.n772 B 0.00831f
C812 VTAIL.n773 B 0.019641f
C813 VTAIL.n774 B 0.008799f
C814 VTAIL.n775 B 0.115865f
C815 VTAIL.t6 B 0.032591f
C816 VTAIL.n776 B 0.014731f
C817 VTAIL.n777 B 0.011603f
C818 VTAIL.n778 B 0.00831f
C819 VTAIL.n779 B 1.28039f
C820 VTAIL.n780 B 0.015464f
C821 VTAIL.n781 B 0.00831f
C822 VTAIL.n782 B 0.008799f
C823 VTAIL.n783 B 0.019641f
C824 VTAIL.n784 B 0.019641f
C825 VTAIL.n785 B 0.008799f
C826 VTAIL.n786 B 0.00831f
C827 VTAIL.n787 B 0.015464f
C828 VTAIL.n788 B 0.015464f
C829 VTAIL.n789 B 0.00831f
C830 VTAIL.n790 B 0.008799f
C831 VTAIL.n791 B 0.019641f
C832 VTAIL.n792 B 0.019641f
C833 VTAIL.n793 B 0.008799f
C834 VTAIL.n794 B 0.00831f
C835 VTAIL.n795 B 0.015464f
C836 VTAIL.n796 B 0.015464f
C837 VTAIL.n797 B 0.00831f
C838 VTAIL.n798 B 0.008799f
C839 VTAIL.n799 B 0.019641f
C840 VTAIL.n800 B 0.019641f
C841 VTAIL.n801 B 0.008799f
C842 VTAIL.n802 B 0.00831f
C843 VTAIL.n803 B 0.015464f
C844 VTAIL.n804 B 0.015464f
C845 VTAIL.n805 B 0.00831f
C846 VTAIL.n806 B 0.008799f
C847 VTAIL.n807 B 0.019641f
C848 VTAIL.n808 B 0.019641f
C849 VTAIL.n809 B 0.008799f
C850 VTAIL.n810 B 0.00831f
C851 VTAIL.n811 B 0.015464f
C852 VTAIL.n812 B 0.015464f
C853 VTAIL.n813 B 0.00831f
C854 VTAIL.n814 B 0.008799f
C855 VTAIL.n815 B 0.019641f
C856 VTAIL.n816 B 0.019641f
C857 VTAIL.n817 B 0.019641f
C858 VTAIL.n818 B 0.008799f
C859 VTAIL.n819 B 0.00831f
C860 VTAIL.n820 B 0.015464f
C861 VTAIL.n821 B 0.015464f
C862 VTAIL.n822 B 0.00831f
C863 VTAIL.n823 B 0.008554f
C864 VTAIL.n824 B 0.008554f
C865 VTAIL.n825 B 0.019641f
C866 VTAIL.n826 B 0.019641f
C867 VTAIL.n827 B 0.008799f
C868 VTAIL.n828 B 0.00831f
C869 VTAIL.n829 B 0.015464f
C870 VTAIL.n830 B 0.015464f
C871 VTAIL.n831 B 0.00831f
C872 VTAIL.n832 B 0.008799f
C873 VTAIL.n833 B 0.019641f
C874 VTAIL.n834 B 0.019641f
C875 VTAIL.n835 B 0.008799f
C876 VTAIL.n836 B 0.00831f
C877 VTAIL.n837 B 0.015464f
C878 VTAIL.n838 B 0.015464f
C879 VTAIL.n839 B 0.00831f
C880 VTAIL.n840 B 0.008799f
C881 VTAIL.n841 B 0.019641f
C882 VTAIL.n842 B 0.041597f
C883 VTAIL.n843 B 0.008799f
C884 VTAIL.n844 B 0.00831f
C885 VTAIL.n845 B 0.033843f
C886 VTAIL.n846 B 0.023121f
C887 VTAIL.n847 B 1.10397f
C888 VDD2.t2 B 0.416629f
C889 VDD2.t1 B 0.416629f
C890 VDD2.n0 B 4.68729f
C891 VDD2.t0 B 0.416629f
C892 VDD2.t3 B 0.416629f
C893 VDD2.n1 B 3.79924f
C894 VDD2.n2 B 4.25169f
C895 VN.t0 B 2.05325f
C896 VN.t1 B 2.05319f
C897 VN.n0 B 1.47114f
C898 VN.t3 B 2.05325f
C899 VN.t2 B 2.05319f
C900 VN.n1 B 2.67017f
.ends

