* NGSPICE file created from diff_pair_sample_0084.ext - technology: sky130A

.subckt diff_pair_sample_0084 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=4.0794 ps=21.7 w=10.46 l=2.54
X1 VTAIL.t9 VN.t1 VDD2.t6 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=1.7259 ps=10.79 w=10.46 l=2.54
X2 VTAIL.t8 VN.t2 VDD2.t5 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X3 B.t11 B.t9 B.t10 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=0 ps=0 w=10.46 l=2.54
X4 VTAIL.t6 VP.t0 VDD1.t7 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X5 VTAIL.t3 VP.t1 VDD1.t6 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=1.7259 ps=10.79 w=10.46 l=2.54
X6 VTAIL.t11 VN.t3 VDD2.t4 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=1.7259 ps=10.79 w=10.46 l=2.54
X7 VTAIL.t15 VN.t4 VDD2.t3 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X8 VDD2.t2 VN.t5 VTAIL.t10 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=4.0794 ps=21.7 w=10.46 l=2.54
X9 VDD1.t5 VP.t2 VTAIL.t1 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=4.0794 ps=21.7 w=10.46 l=2.54
X10 VTAIL.t2 VP.t3 VDD1.t4 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X11 B.t8 B.t6 B.t7 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=0 ps=0 w=10.46 l=2.54
X12 B.t5 B.t3 B.t4 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=0 ps=0 w=10.46 l=2.54
X13 VDD2.t1 VN.t6 VTAIL.t14 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X14 VDD1.t3 VP.t4 VTAIL.t5 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=4.0794 ps=21.7 w=10.46 l=2.54
X15 VDD2.t0 VN.t7 VTAIL.t13 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X16 VDD1.t2 VP.t5 VTAIL.t0 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X17 VTAIL.t7 VP.t6 VDD1.t1 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=1.7259 ps=10.79 w=10.46 l=2.54
X18 VDD1.t0 VP.t7 VTAIL.t4 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=1.7259 pd=10.79 as=1.7259 ps=10.79 w=10.46 l=2.54
X19 B.t2 B.t0 B.t1 w_n3840_n3060# sky130_fd_pr__pfet_01v8 ad=4.0794 pd=21.7 as=0 ps=0 w=10.46 l=2.54
R0 VN.n55 VN.n29 161.3
R1 VN.n54 VN.n53 161.3
R2 VN.n52 VN.n30 161.3
R3 VN.n51 VN.n50 161.3
R4 VN.n49 VN.n31 161.3
R5 VN.n48 VN.n47 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n26 VN.n0 161.3
R13 VN.n25 VN.n24 161.3
R14 VN.n23 VN.n1 161.3
R15 VN.n22 VN.n21 161.3
R16 VN.n20 VN.n2 161.3
R17 VN.n19 VN.n18 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n7 VN.t1 130.329
R25 VN.n36 VN.t5 130.329
R26 VN.n28 VN.n27 107.928
R27 VN.n57 VN.n56 107.928
R28 VN.n8 VN.t7 99.247
R29 VN.n3 VN.t4 99.247
R30 VN.n27 VN.t0 99.247
R31 VN.n37 VN.t2 99.247
R32 VN.n32 VN.t6 99.247
R33 VN.n56 VN.t3 99.247
R34 VN.n8 VN.n7 63.2583
R35 VN.n37 VN.n36 63.2583
R36 VN.n14 VN.n5 56.4773
R37 VN.n43 VN.n34 56.4773
R38 VN.n21 VN.n1 52.0954
R39 VN.n50 VN.n30 52.0954
R40 VN VN.n57 49.6193
R41 VN.n21 VN.n20 28.7258
R42 VN.n50 VN.n49 28.7258
R43 VN.n10 VN.n9 24.3439
R44 VN.n10 VN.n5 24.3439
R45 VN.n15 VN.n14 24.3439
R46 VN.n16 VN.n15 24.3439
R47 VN.n20 VN.n19 24.3439
R48 VN.n25 VN.n1 24.3439
R49 VN.n26 VN.n25 24.3439
R50 VN.n39 VN.n34 24.3439
R51 VN.n39 VN.n38 24.3439
R52 VN.n49 VN.n48 24.3439
R53 VN.n45 VN.n44 24.3439
R54 VN.n44 VN.n43 24.3439
R55 VN.n55 VN.n54 24.3439
R56 VN.n54 VN.n30 24.3439
R57 VN.n19 VN.n3 15.3369
R58 VN.n48 VN.n32 15.3369
R59 VN.n9 VN.n8 9.00757
R60 VN.n16 VN.n3 9.00757
R61 VN.n38 VN.n37 9.00757
R62 VN.n45 VN.n32 9.00757
R63 VN.n36 VN.n35 7.32939
R64 VN.n7 VN.n6 7.32939
R65 VN.n27 VN.n26 2.67828
R66 VN.n56 VN.n55 2.67828
R67 VN.n57 VN.n29 0.278398
R68 VN.n28 VN.n0 0.278398
R69 VN.n53 VN.n29 0.189894
R70 VN.n53 VN.n52 0.189894
R71 VN.n52 VN.n51 0.189894
R72 VN.n51 VN.n31 0.189894
R73 VN.n47 VN.n31 0.189894
R74 VN.n47 VN.n46 0.189894
R75 VN.n46 VN.n33 0.189894
R76 VN.n42 VN.n33 0.189894
R77 VN.n42 VN.n41 0.189894
R78 VN.n41 VN.n40 0.189894
R79 VN.n40 VN.n35 0.189894
R80 VN.n11 VN.n6 0.189894
R81 VN.n12 VN.n11 0.189894
R82 VN.n13 VN.n12 0.189894
R83 VN.n13 VN.n4 0.189894
R84 VN.n17 VN.n4 0.189894
R85 VN.n18 VN.n17 0.189894
R86 VN.n18 VN.n2 0.189894
R87 VN.n22 VN.n2 0.189894
R88 VN.n23 VN.n22 0.189894
R89 VN.n24 VN.n23 0.189894
R90 VN.n24 VN.n0 0.189894
R91 VN VN.n28 0.153422
R92 VTAIL.n11 VTAIL.t3 65.6126
R93 VTAIL.n10 VTAIL.t10 65.6126
R94 VTAIL.n7 VTAIL.t11 65.6126
R95 VTAIL.n14 VTAIL.t5 65.6124
R96 VTAIL.n15 VTAIL.t12 65.6124
R97 VTAIL.n2 VTAIL.t9 65.6124
R98 VTAIL.n3 VTAIL.t1 65.6124
R99 VTAIL.n6 VTAIL.t7 65.6124
R100 VTAIL.n13 VTAIL.n12 62.5051
R101 VTAIL.n9 VTAIL.n8 62.5051
R102 VTAIL.n1 VTAIL.n0 62.5048
R103 VTAIL.n5 VTAIL.n4 62.5048
R104 VTAIL.n15 VTAIL.n14 23.8583
R105 VTAIL.n7 VTAIL.n6 23.8583
R106 VTAIL.n0 VTAIL.t13 3.10805
R107 VTAIL.n0 VTAIL.t15 3.10805
R108 VTAIL.n4 VTAIL.t0 3.10805
R109 VTAIL.n4 VTAIL.t2 3.10805
R110 VTAIL.n12 VTAIL.t4 3.10805
R111 VTAIL.n12 VTAIL.t6 3.10805
R112 VTAIL.n8 VTAIL.t14 3.10805
R113 VTAIL.n8 VTAIL.t8 3.10805
R114 VTAIL.n9 VTAIL.n7 2.47464
R115 VTAIL.n10 VTAIL.n9 2.47464
R116 VTAIL.n13 VTAIL.n11 2.47464
R117 VTAIL.n14 VTAIL.n13 2.47464
R118 VTAIL.n6 VTAIL.n5 2.47464
R119 VTAIL.n5 VTAIL.n3 2.47464
R120 VTAIL.n2 VTAIL.n1 2.47464
R121 VTAIL VTAIL.n15 2.41645
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 80.3653
R126 VDD2.n2 VDD2.n0 80.3653
R127 VDD2 VDD2.n5 80.3625
R128 VDD2.n4 VDD2.n3 79.1839
R129 VDD2.n4 VDD2.n2 43.8662
R130 VDD2.n5 VDD2.t5 3.10805
R131 VDD2.n5 VDD2.t2 3.10805
R132 VDD2.n3 VDD2.t4 3.10805
R133 VDD2.n3 VDD2.t1 3.10805
R134 VDD2.n1 VDD2.t3 3.10805
R135 VDD2.n1 VDD2.t7 3.10805
R136 VDD2.n0 VDD2.t6 3.10805
R137 VDD2.n0 VDD2.t0 3.10805
R138 VDD2 VDD2.n4 1.29576
R139 B.n396 B.n125 585
R140 B.n395 B.n394 585
R141 B.n393 B.n126 585
R142 B.n392 B.n391 585
R143 B.n390 B.n127 585
R144 B.n389 B.n388 585
R145 B.n387 B.n128 585
R146 B.n386 B.n385 585
R147 B.n384 B.n129 585
R148 B.n383 B.n382 585
R149 B.n381 B.n130 585
R150 B.n380 B.n379 585
R151 B.n378 B.n131 585
R152 B.n377 B.n376 585
R153 B.n375 B.n132 585
R154 B.n374 B.n373 585
R155 B.n372 B.n133 585
R156 B.n371 B.n370 585
R157 B.n369 B.n134 585
R158 B.n368 B.n367 585
R159 B.n366 B.n135 585
R160 B.n365 B.n364 585
R161 B.n363 B.n136 585
R162 B.n362 B.n361 585
R163 B.n360 B.n137 585
R164 B.n359 B.n358 585
R165 B.n357 B.n138 585
R166 B.n356 B.n355 585
R167 B.n354 B.n139 585
R168 B.n353 B.n352 585
R169 B.n351 B.n140 585
R170 B.n350 B.n349 585
R171 B.n348 B.n141 585
R172 B.n347 B.n346 585
R173 B.n345 B.n142 585
R174 B.n344 B.n343 585
R175 B.n342 B.n143 585
R176 B.n341 B.n340 585
R177 B.n336 B.n144 585
R178 B.n335 B.n334 585
R179 B.n333 B.n145 585
R180 B.n332 B.n331 585
R181 B.n330 B.n146 585
R182 B.n329 B.n328 585
R183 B.n327 B.n147 585
R184 B.n326 B.n325 585
R185 B.n324 B.n148 585
R186 B.n322 B.n321 585
R187 B.n320 B.n151 585
R188 B.n319 B.n318 585
R189 B.n317 B.n152 585
R190 B.n316 B.n315 585
R191 B.n314 B.n153 585
R192 B.n313 B.n312 585
R193 B.n311 B.n154 585
R194 B.n310 B.n309 585
R195 B.n308 B.n155 585
R196 B.n307 B.n306 585
R197 B.n305 B.n156 585
R198 B.n304 B.n303 585
R199 B.n302 B.n157 585
R200 B.n301 B.n300 585
R201 B.n299 B.n158 585
R202 B.n298 B.n297 585
R203 B.n296 B.n159 585
R204 B.n295 B.n294 585
R205 B.n293 B.n160 585
R206 B.n292 B.n291 585
R207 B.n290 B.n161 585
R208 B.n289 B.n288 585
R209 B.n287 B.n162 585
R210 B.n286 B.n285 585
R211 B.n284 B.n163 585
R212 B.n283 B.n282 585
R213 B.n281 B.n164 585
R214 B.n280 B.n279 585
R215 B.n278 B.n165 585
R216 B.n277 B.n276 585
R217 B.n275 B.n166 585
R218 B.n274 B.n273 585
R219 B.n272 B.n167 585
R220 B.n271 B.n270 585
R221 B.n269 B.n168 585
R222 B.n268 B.n267 585
R223 B.n398 B.n397 585
R224 B.n399 B.n124 585
R225 B.n401 B.n400 585
R226 B.n402 B.n123 585
R227 B.n404 B.n403 585
R228 B.n405 B.n122 585
R229 B.n407 B.n406 585
R230 B.n408 B.n121 585
R231 B.n410 B.n409 585
R232 B.n411 B.n120 585
R233 B.n413 B.n412 585
R234 B.n414 B.n119 585
R235 B.n416 B.n415 585
R236 B.n417 B.n118 585
R237 B.n419 B.n418 585
R238 B.n420 B.n117 585
R239 B.n422 B.n421 585
R240 B.n423 B.n116 585
R241 B.n425 B.n424 585
R242 B.n426 B.n115 585
R243 B.n428 B.n427 585
R244 B.n429 B.n114 585
R245 B.n431 B.n430 585
R246 B.n432 B.n113 585
R247 B.n434 B.n433 585
R248 B.n435 B.n112 585
R249 B.n437 B.n436 585
R250 B.n438 B.n111 585
R251 B.n440 B.n439 585
R252 B.n441 B.n110 585
R253 B.n443 B.n442 585
R254 B.n444 B.n109 585
R255 B.n446 B.n445 585
R256 B.n447 B.n108 585
R257 B.n449 B.n448 585
R258 B.n450 B.n107 585
R259 B.n452 B.n451 585
R260 B.n453 B.n106 585
R261 B.n455 B.n454 585
R262 B.n456 B.n105 585
R263 B.n458 B.n457 585
R264 B.n459 B.n104 585
R265 B.n461 B.n460 585
R266 B.n462 B.n103 585
R267 B.n464 B.n463 585
R268 B.n465 B.n102 585
R269 B.n467 B.n466 585
R270 B.n468 B.n101 585
R271 B.n470 B.n469 585
R272 B.n471 B.n100 585
R273 B.n473 B.n472 585
R274 B.n474 B.n99 585
R275 B.n476 B.n475 585
R276 B.n477 B.n98 585
R277 B.n479 B.n478 585
R278 B.n480 B.n97 585
R279 B.n482 B.n481 585
R280 B.n483 B.n96 585
R281 B.n485 B.n484 585
R282 B.n486 B.n95 585
R283 B.n488 B.n487 585
R284 B.n489 B.n94 585
R285 B.n491 B.n490 585
R286 B.n492 B.n93 585
R287 B.n494 B.n493 585
R288 B.n495 B.n92 585
R289 B.n497 B.n496 585
R290 B.n498 B.n91 585
R291 B.n500 B.n499 585
R292 B.n501 B.n90 585
R293 B.n503 B.n502 585
R294 B.n504 B.n89 585
R295 B.n506 B.n505 585
R296 B.n507 B.n88 585
R297 B.n509 B.n508 585
R298 B.n510 B.n87 585
R299 B.n512 B.n511 585
R300 B.n513 B.n86 585
R301 B.n515 B.n514 585
R302 B.n516 B.n85 585
R303 B.n518 B.n517 585
R304 B.n519 B.n84 585
R305 B.n521 B.n520 585
R306 B.n522 B.n83 585
R307 B.n524 B.n523 585
R308 B.n525 B.n82 585
R309 B.n527 B.n526 585
R310 B.n528 B.n81 585
R311 B.n530 B.n529 585
R312 B.n531 B.n80 585
R313 B.n533 B.n532 585
R314 B.n534 B.n79 585
R315 B.n536 B.n535 585
R316 B.n537 B.n78 585
R317 B.n539 B.n538 585
R318 B.n540 B.n77 585
R319 B.n542 B.n541 585
R320 B.n543 B.n76 585
R321 B.n545 B.n544 585
R322 B.n546 B.n75 585
R323 B.n548 B.n547 585
R324 B.n549 B.n74 585
R325 B.n676 B.n27 585
R326 B.n675 B.n674 585
R327 B.n673 B.n28 585
R328 B.n672 B.n671 585
R329 B.n670 B.n29 585
R330 B.n669 B.n668 585
R331 B.n667 B.n30 585
R332 B.n666 B.n665 585
R333 B.n664 B.n31 585
R334 B.n663 B.n662 585
R335 B.n661 B.n32 585
R336 B.n660 B.n659 585
R337 B.n658 B.n33 585
R338 B.n657 B.n656 585
R339 B.n655 B.n34 585
R340 B.n654 B.n653 585
R341 B.n652 B.n35 585
R342 B.n651 B.n650 585
R343 B.n649 B.n36 585
R344 B.n648 B.n647 585
R345 B.n646 B.n37 585
R346 B.n645 B.n644 585
R347 B.n643 B.n38 585
R348 B.n642 B.n641 585
R349 B.n640 B.n39 585
R350 B.n639 B.n638 585
R351 B.n637 B.n40 585
R352 B.n636 B.n635 585
R353 B.n634 B.n41 585
R354 B.n633 B.n632 585
R355 B.n631 B.n42 585
R356 B.n630 B.n629 585
R357 B.n628 B.n43 585
R358 B.n627 B.n626 585
R359 B.n625 B.n44 585
R360 B.n624 B.n623 585
R361 B.n622 B.n45 585
R362 B.n620 B.n619 585
R363 B.n618 B.n48 585
R364 B.n617 B.n616 585
R365 B.n615 B.n49 585
R366 B.n614 B.n613 585
R367 B.n612 B.n50 585
R368 B.n611 B.n610 585
R369 B.n609 B.n51 585
R370 B.n608 B.n607 585
R371 B.n606 B.n52 585
R372 B.n605 B.n604 585
R373 B.n603 B.n53 585
R374 B.n602 B.n601 585
R375 B.n600 B.n57 585
R376 B.n599 B.n598 585
R377 B.n597 B.n58 585
R378 B.n596 B.n595 585
R379 B.n594 B.n59 585
R380 B.n593 B.n592 585
R381 B.n591 B.n60 585
R382 B.n590 B.n589 585
R383 B.n588 B.n61 585
R384 B.n587 B.n586 585
R385 B.n585 B.n62 585
R386 B.n584 B.n583 585
R387 B.n582 B.n63 585
R388 B.n581 B.n580 585
R389 B.n579 B.n64 585
R390 B.n578 B.n577 585
R391 B.n576 B.n65 585
R392 B.n575 B.n574 585
R393 B.n573 B.n66 585
R394 B.n572 B.n571 585
R395 B.n570 B.n67 585
R396 B.n569 B.n568 585
R397 B.n567 B.n68 585
R398 B.n566 B.n565 585
R399 B.n564 B.n69 585
R400 B.n563 B.n562 585
R401 B.n561 B.n70 585
R402 B.n560 B.n559 585
R403 B.n558 B.n71 585
R404 B.n557 B.n556 585
R405 B.n555 B.n72 585
R406 B.n554 B.n553 585
R407 B.n552 B.n73 585
R408 B.n551 B.n550 585
R409 B.n678 B.n677 585
R410 B.n679 B.n26 585
R411 B.n681 B.n680 585
R412 B.n682 B.n25 585
R413 B.n684 B.n683 585
R414 B.n685 B.n24 585
R415 B.n687 B.n686 585
R416 B.n688 B.n23 585
R417 B.n690 B.n689 585
R418 B.n691 B.n22 585
R419 B.n693 B.n692 585
R420 B.n694 B.n21 585
R421 B.n696 B.n695 585
R422 B.n697 B.n20 585
R423 B.n699 B.n698 585
R424 B.n700 B.n19 585
R425 B.n702 B.n701 585
R426 B.n703 B.n18 585
R427 B.n705 B.n704 585
R428 B.n706 B.n17 585
R429 B.n708 B.n707 585
R430 B.n709 B.n16 585
R431 B.n711 B.n710 585
R432 B.n712 B.n15 585
R433 B.n714 B.n713 585
R434 B.n715 B.n14 585
R435 B.n717 B.n716 585
R436 B.n718 B.n13 585
R437 B.n720 B.n719 585
R438 B.n721 B.n12 585
R439 B.n723 B.n722 585
R440 B.n724 B.n11 585
R441 B.n726 B.n725 585
R442 B.n727 B.n10 585
R443 B.n729 B.n728 585
R444 B.n730 B.n9 585
R445 B.n732 B.n731 585
R446 B.n733 B.n8 585
R447 B.n735 B.n734 585
R448 B.n736 B.n7 585
R449 B.n738 B.n737 585
R450 B.n739 B.n6 585
R451 B.n741 B.n740 585
R452 B.n742 B.n5 585
R453 B.n744 B.n743 585
R454 B.n745 B.n4 585
R455 B.n747 B.n746 585
R456 B.n748 B.n3 585
R457 B.n750 B.n749 585
R458 B.n751 B.n0 585
R459 B.n2 B.n1 585
R460 B.n194 B.n193 585
R461 B.n196 B.n195 585
R462 B.n197 B.n192 585
R463 B.n199 B.n198 585
R464 B.n200 B.n191 585
R465 B.n202 B.n201 585
R466 B.n203 B.n190 585
R467 B.n205 B.n204 585
R468 B.n206 B.n189 585
R469 B.n208 B.n207 585
R470 B.n209 B.n188 585
R471 B.n211 B.n210 585
R472 B.n212 B.n187 585
R473 B.n214 B.n213 585
R474 B.n215 B.n186 585
R475 B.n217 B.n216 585
R476 B.n218 B.n185 585
R477 B.n220 B.n219 585
R478 B.n221 B.n184 585
R479 B.n223 B.n222 585
R480 B.n224 B.n183 585
R481 B.n226 B.n225 585
R482 B.n227 B.n182 585
R483 B.n229 B.n228 585
R484 B.n230 B.n181 585
R485 B.n232 B.n231 585
R486 B.n233 B.n180 585
R487 B.n235 B.n234 585
R488 B.n236 B.n179 585
R489 B.n238 B.n237 585
R490 B.n239 B.n178 585
R491 B.n241 B.n240 585
R492 B.n242 B.n177 585
R493 B.n244 B.n243 585
R494 B.n245 B.n176 585
R495 B.n247 B.n246 585
R496 B.n248 B.n175 585
R497 B.n250 B.n249 585
R498 B.n251 B.n174 585
R499 B.n253 B.n252 585
R500 B.n254 B.n173 585
R501 B.n256 B.n255 585
R502 B.n257 B.n172 585
R503 B.n259 B.n258 585
R504 B.n260 B.n171 585
R505 B.n262 B.n261 585
R506 B.n263 B.n170 585
R507 B.n265 B.n264 585
R508 B.n266 B.n169 585
R509 B.n267 B.n266 449.257
R510 B.n397 B.n396 449.257
R511 B.n551 B.n74 449.257
R512 B.n678 B.n27 449.257
R513 B.n149 B.t3 307.202
R514 B.n337 B.t0 307.202
R515 B.n54 B.t6 307.202
R516 B.n46 B.t9 307.202
R517 B.n753 B.n752 256.663
R518 B.n752 B.n751 235.042
R519 B.n752 B.n2 235.042
R520 B.n337 B.t1 168.226
R521 B.n54 B.t8 168.226
R522 B.n149 B.t4 168.214
R523 B.n46 B.t11 168.214
R524 B.n267 B.n168 163.367
R525 B.n271 B.n168 163.367
R526 B.n272 B.n271 163.367
R527 B.n273 B.n272 163.367
R528 B.n273 B.n166 163.367
R529 B.n277 B.n166 163.367
R530 B.n278 B.n277 163.367
R531 B.n279 B.n278 163.367
R532 B.n279 B.n164 163.367
R533 B.n283 B.n164 163.367
R534 B.n284 B.n283 163.367
R535 B.n285 B.n284 163.367
R536 B.n285 B.n162 163.367
R537 B.n289 B.n162 163.367
R538 B.n290 B.n289 163.367
R539 B.n291 B.n290 163.367
R540 B.n291 B.n160 163.367
R541 B.n295 B.n160 163.367
R542 B.n296 B.n295 163.367
R543 B.n297 B.n296 163.367
R544 B.n297 B.n158 163.367
R545 B.n301 B.n158 163.367
R546 B.n302 B.n301 163.367
R547 B.n303 B.n302 163.367
R548 B.n303 B.n156 163.367
R549 B.n307 B.n156 163.367
R550 B.n308 B.n307 163.367
R551 B.n309 B.n308 163.367
R552 B.n309 B.n154 163.367
R553 B.n313 B.n154 163.367
R554 B.n314 B.n313 163.367
R555 B.n315 B.n314 163.367
R556 B.n315 B.n152 163.367
R557 B.n319 B.n152 163.367
R558 B.n320 B.n319 163.367
R559 B.n321 B.n320 163.367
R560 B.n321 B.n148 163.367
R561 B.n326 B.n148 163.367
R562 B.n327 B.n326 163.367
R563 B.n328 B.n327 163.367
R564 B.n328 B.n146 163.367
R565 B.n332 B.n146 163.367
R566 B.n333 B.n332 163.367
R567 B.n334 B.n333 163.367
R568 B.n334 B.n144 163.367
R569 B.n341 B.n144 163.367
R570 B.n342 B.n341 163.367
R571 B.n343 B.n342 163.367
R572 B.n343 B.n142 163.367
R573 B.n347 B.n142 163.367
R574 B.n348 B.n347 163.367
R575 B.n349 B.n348 163.367
R576 B.n349 B.n140 163.367
R577 B.n353 B.n140 163.367
R578 B.n354 B.n353 163.367
R579 B.n355 B.n354 163.367
R580 B.n355 B.n138 163.367
R581 B.n359 B.n138 163.367
R582 B.n360 B.n359 163.367
R583 B.n361 B.n360 163.367
R584 B.n361 B.n136 163.367
R585 B.n365 B.n136 163.367
R586 B.n366 B.n365 163.367
R587 B.n367 B.n366 163.367
R588 B.n367 B.n134 163.367
R589 B.n371 B.n134 163.367
R590 B.n372 B.n371 163.367
R591 B.n373 B.n372 163.367
R592 B.n373 B.n132 163.367
R593 B.n377 B.n132 163.367
R594 B.n378 B.n377 163.367
R595 B.n379 B.n378 163.367
R596 B.n379 B.n130 163.367
R597 B.n383 B.n130 163.367
R598 B.n384 B.n383 163.367
R599 B.n385 B.n384 163.367
R600 B.n385 B.n128 163.367
R601 B.n389 B.n128 163.367
R602 B.n390 B.n389 163.367
R603 B.n391 B.n390 163.367
R604 B.n391 B.n126 163.367
R605 B.n395 B.n126 163.367
R606 B.n396 B.n395 163.367
R607 B.n547 B.n74 163.367
R608 B.n547 B.n546 163.367
R609 B.n546 B.n545 163.367
R610 B.n545 B.n76 163.367
R611 B.n541 B.n76 163.367
R612 B.n541 B.n540 163.367
R613 B.n540 B.n539 163.367
R614 B.n539 B.n78 163.367
R615 B.n535 B.n78 163.367
R616 B.n535 B.n534 163.367
R617 B.n534 B.n533 163.367
R618 B.n533 B.n80 163.367
R619 B.n529 B.n80 163.367
R620 B.n529 B.n528 163.367
R621 B.n528 B.n527 163.367
R622 B.n527 B.n82 163.367
R623 B.n523 B.n82 163.367
R624 B.n523 B.n522 163.367
R625 B.n522 B.n521 163.367
R626 B.n521 B.n84 163.367
R627 B.n517 B.n84 163.367
R628 B.n517 B.n516 163.367
R629 B.n516 B.n515 163.367
R630 B.n515 B.n86 163.367
R631 B.n511 B.n86 163.367
R632 B.n511 B.n510 163.367
R633 B.n510 B.n509 163.367
R634 B.n509 B.n88 163.367
R635 B.n505 B.n88 163.367
R636 B.n505 B.n504 163.367
R637 B.n504 B.n503 163.367
R638 B.n503 B.n90 163.367
R639 B.n499 B.n90 163.367
R640 B.n499 B.n498 163.367
R641 B.n498 B.n497 163.367
R642 B.n497 B.n92 163.367
R643 B.n493 B.n92 163.367
R644 B.n493 B.n492 163.367
R645 B.n492 B.n491 163.367
R646 B.n491 B.n94 163.367
R647 B.n487 B.n94 163.367
R648 B.n487 B.n486 163.367
R649 B.n486 B.n485 163.367
R650 B.n485 B.n96 163.367
R651 B.n481 B.n96 163.367
R652 B.n481 B.n480 163.367
R653 B.n480 B.n479 163.367
R654 B.n479 B.n98 163.367
R655 B.n475 B.n98 163.367
R656 B.n475 B.n474 163.367
R657 B.n474 B.n473 163.367
R658 B.n473 B.n100 163.367
R659 B.n469 B.n100 163.367
R660 B.n469 B.n468 163.367
R661 B.n468 B.n467 163.367
R662 B.n467 B.n102 163.367
R663 B.n463 B.n102 163.367
R664 B.n463 B.n462 163.367
R665 B.n462 B.n461 163.367
R666 B.n461 B.n104 163.367
R667 B.n457 B.n104 163.367
R668 B.n457 B.n456 163.367
R669 B.n456 B.n455 163.367
R670 B.n455 B.n106 163.367
R671 B.n451 B.n106 163.367
R672 B.n451 B.n450 163.367
R673 B.n450 B.n449 163.367
R674 B.n449 B.n108 163.367
R675 B.n445 B.n108 163.367
R676 B.n445 B.n444 163.367
R677 B.n444 B.n443 163.367
R678 B.n443 B.n110 163.367
R679 B.n439 B.n110 163.367
R680 B.n439 B.n438 163.367
R681 B.n438 B.n437 163.367
R682 B.n437 B.n112 163.367
R683 B.n433 B.n112 163.367
R684 B.n433 B.n432 163.367
R685 B.n432 B.n431 163.367
R686 B.n431 B.n114 163.367
R687 B.n427 B.n114 163.367
R688 B.n427 B.n426 163.367
R689 B.n426 B.n425 163.367
R690 B.n425 B.n116 163.367
R691 B.n421 B.n116 163.367
R692 B.n421 B.n420 163.367
R693 B.n420 B.n419 163.367
R694 B.n419 B.n118 163.367
R695 B.n415 B.n118 163.367
R696 B.n415 B.n414 163.367
R697 B.n414 B.n413 163.367
R698 B.n413 B.n120 163.367
R699 B.n409 B.n120 163.367
R700 B.n409 B.n408 163.367
R701 B.n408 B.n407 163.367
R702 B.n407 B.n122 163.367
R703 B.n403 B.n122 163.367
R704 B.n403 B.n402 163.367
R705 B.n402 B.n401 163.367
R706 B.n401 B.n124 163.367
R707 B.n397 B.n124 163.367
R708 B.n674 B.n27 163.367
R709 B.n674 B.n673 163.367
R710 B.n673 B.n672 163.367
R711 B.n672 B.n29 163.367
R712 B.n668 B.n29 163.367
R713 B.n668 B.n667 163.367
R714 B.n667 B.n666 163.367
R715 B.n666 B.n31 163.367
R716 B.n662 B.n31 163.367
R717 B.n662 B.n661 163.367
R718 B.n661 B.n660 163.367
R719 B.n660 B.n33 163.367
R720 B.n656 B.n33 163.367
R721 B.n656 B.n655 163.367
R722 B.n655 B.n654 163.367
R723 B.n654 B.n35 163.367
R724 B.n650 B.n35 163.367
R725 B.n650 B.n649 163.367
R726 B.n649 B.n648 163.367
R727 B.n648 B.n37 163.367
R728 B.n644 B.n37 163.367
R729 B.n644 B.n643 163.367
R730 B.n643 B.n642 163.367
R731 B.n642 B.n39 163.367
R732 B.n638 B.n39 163.367
R733 B.n638 B.n637 163.367
R734 B.n637 B.n636 163.367
R735 B.n636 B.n41 163.367
R736 B.n632 B.n41 163.367
R737 B.n632 B.n631 163.367
R738 B.n631 B.n630 163.367
R739 B.n630 B.n43 163.367
R740 B.n626 B.n43 163.367
R741 B.n626 B.n625 163.367
R742 B.n625 B.n624 163.367
R743 B.n624 B.n45 163.367
R744 B.n619 B.n45 163.367
R745 B.n619 B.n618 163.367
R746 B.n618 B.n617 163.367
R747 B.n617 B.n49 163.367
R748 B.n613 B.n49 163.367
R749 B.n613 B.n612 163.367
R750 B.n612 B.n611 163.367
R751 B.n611 B.n51 163.367
R752 B.n607 B.n51 163.367
R753 B.n607 B.n606 163.367
R754 B.n606 B.n605 163.367
R755 B.n605 B.n53 163.367
R756 B.n601 B.n53 163.367
R757 B.n601 B.n600 163.367
R758 B.n600 B.n599 163.367
R759 B.n599 B.n58 163.367
R760 B.n595 B.n58 163.367
R761 B.n595 B.n594 163.367
R762 B.n594 B.n593 163.367
R763 B.n593 B.n60 163.367
R764 B.n589 B.n60 163.367
R765 B.n589 B.n588 163.367
R766 B.n588 B.n587 163.367
R767 B.n587 B.n62 163.367
R768 B.n583 B.n62 163.367
R769 B.n583 B.n582 163.367
R770 B.n582 B.n581 163.367
R771 B.n581 B.n64 163.367
R772 B.n577 B.n64 163.367
R773 B.n577 B.n576 163.367
R774 B.n576 B.n575 163.367
R775 B.n575 B.n66 163.367
R776 B.n571 B.n66 163.367
R777 B.n571 B.n570 163.367
R778 B.n570 B.n569 163.367
R779 B.n569 B.n68 163.367
R780 B.n565 B.n68 163.367
R781 B.n565 B.n564 163.367
R782 B.n564 B.n563 163.367
R783 B.n563 B.n70 163.367
R784 B.n559 B.n70 163.367
R785 B.n559 B.n558 163.367
R786 B.n558 B.n557 163.367
R787 B.n557 B.n72 163.367
R788 B.n553 B.n72 163.367
R789 B.n553 B.n552 163.367
R790 B.n552 B.n551 163.367
R791 B.n679 B.n678 163.367
R792 B.n680 B.n679 163.367
R793 B.n680 B.n25 163.367
R794 B.n684 B.n25 163.367
R795 B.n685 B.n684 163.367
R796 B.n686 B.n685 163.367
R797 B.n686 B.n23 163.367
R798 B.n690 B.n23 163.367
R799 B.n691 B.n690 163.367
R800 B.n692 B.n691 163.367
R801 B.n692 B.n21 163.367
R802 B.n696 B.n21 163.367
R803 B.n697 B.n696 163.367
R804 B.n698 B.n697 163.367
R805 B.n698 B.n19 163.367
R806 B.n702 B.n19 163.367
R807 B.n703 B.n702 163.367
R808 B.n704 B.n703 163.367
R809 B.n704 B.n17 163.367
R810 B.n708 B.n17 163.367
R811 B.n709 B.n708 163.367
R812 B.n710 B.n709 163.367
R813 B.n710 B.n15 163.367
R814 B.n714 B.n15 163.367
R815 B.n715 B.n714 163.367
R816 B.n716 B.n715 163.367
R817 B.n716 B.n13 163.367
R818 B.n720 B.n13 163.367
R819 B.n721 B.n720 163.367
R820 B.n722 B.n721 163.367
R821 B.n722 B.n11 163.367
R822 B.n726 B.n11 163.367
R823 B.n727 B.n726 163.367
R824 B.n728 B.n727 163.367
R825 B.n728 B.n9 163.367
R826 B.n732 B.n9 163.367
R827 B.n733 B.n732 163.367
R828 B.n734 B.n733 163.367
R829 B.n734 B.n7 163.367
R830 B.n738 B.n7 163.367
R831 B.n739 B.n738 163.367
R832 B.n740 B.n739 163.367
R833 B.n740 B.n5 163.367
R834 B.n744 B.n5 163.367
R835 B.n745 B.n744 163.367
R836 B.n746 B.n745 163.367
R837 B.n746 B.n3 163.367
R838 B.n750 B.n3 163.367
R839 B.n751 B.n750 163.367
R840 B.n194 B.n2 163.367
R841 B.n195 B.n194 163.367
R842 B.n195 B.n192 163.367
R843 B.n199 B.n192 163.367
R844 B.n200 B.n199 163.367
R845 B.n201 B.n200 163.367
R846 B.n201 B.n190 163.367
R847 B.n205 B.n190 163.367
R848 B.n206 B.n205 163.367
R849 B.n207 B.n206 163.367
R850 B.n207 B.n188 163.367
R851 B.n211 B.n188 163.367
R852 B.n212 B.n211 163.367
R853 B.n213 B.n212 163.367
R854 B.n213 B.n186 163.367
R855 B.n217 B.n186 163.367
R856 B.n218 B.n217 163.367
R857 B.n219 B.n218 163.367
R858 B.n219 B.n184 163.367
R859 B.n223 B.n184 163.367
R860 B.n224 B.n223 163.367
R861 B.n225 B.n224 163.367
R862 B.n225 B.n182 163.367
R863 B.n229 B.n182 163.367
R864 B.n230 B.n229 163.367
R865 B.n231 B.n230 163.367
R866 B.n231 B.n180 163.367
R867 B.n235 B.n180 163.367
R868 B.n236 B.n235 163.367
R869 B.n237 B.n236 163.367
R870 B.n237 B.n178 163.367
R871 B.n241 B.n178 163.367
R872 B.n242 B.n241 163.367
R873 B.n243 B.n242 163.367
R874 B.n243 B.n176 163.367
R875 B.n247 B.n176 163.367
R876 B.n248 B.n247 163.367
R877 B.n249 B.n248 163.367
R878 B.n249 B.n174 163.367
R879 B.n253 B.n174 163.367
R880 B.n254 B.n253 163.367
R881 B.n255 B.n254 163.367
R882 B.n255 B.n172 163.367
R883 B.n259 B.n172 163.367
R884 B.n260 B.n259 163.367
R885 B.n261 B.n260 163.367
R886 B.n261 B.n170 163.367
R887 B.n265 B.n170 163.367
R888 B.n266 B.n265 163.367
R889 B.n338 B.t2 112.567
R890 B.n55 B.t7 112.567
R891 B.n150 B.t5 112.555
R892 B.n47 B.t10 112.555
R893 B.n323 B.n150 59.5399
R894 B.n339 B.n338 59.5399
R895 B.n56 B.n55 59.5399
R896 B.n621 B.n47 59.5399
R897 B.n150 B.n149 55.6611
R898 B.n338 B.n337 55.6611
R899 B.n55 B.n54 55.6611
R900 B.n47 B.n46 55.6611
R901 B.n677 B.n676 29.1907
R902 B.n550 B.n549 29.1907
R903 B.n268 B.n169 29.1907
R904 B.n398 B.n125 29.1907
R905 B B.n753 18.0485
R906 B.n677 B.n26 10.6151
R907 B.n681 B.n26 10.6151
R908 B.n682 B.n681 10.6151
R909 B.n683 B.n682 10.6151
R910 B.n683 B.n24 10.6151
R911 B.n687 B.n24 10.6151
R912 B.n688 B.n687 10.6151
R913 B.n689 B.n688 10.6151
R914 B.n689 B.n22 10.6151
R915 B.n693 B.n22 10.6151
R916 B.n694 B.n693 10.6151
R917 B.n695 B.n694 10.6151
R918 B.n695 B.n20 10.6151
R919 B.n699 B.n20 10.6151
R920 B.n700 B.n699 10.6151
R921 B.n701 B.n700 10.6151
R922 B.n701 B.n18 10.6151
R923 B.n705 B.n18 10.6151
R924 B.n706 B.n705 10.6151
R925 B.n707 B.n706 10.6151
R926 B.n707 B.n16 10.6151
R927 B.n711 B.n16 10.6151
R928 B.n712 B.n711 10.6151
R929 B.n713 B.n712 10.6151
R930 B.n713 B.n14 10.6151
R931 B.n717 B.n14 10.6151
R932 B.n718 B.n717 10.6151
R933 B.n719 B.n718 10.6151
R934 B.n719 B.n12 10.6151
R935 B.n723 B.n12 10.6151
R936 B.n724 B.n723 10.6151
R937 B.n725 B.n724 10.6151
R938 B.n725 B.n10 10.6151
R939 B.n729 B.n10 10.6151
R940 B.n730 B.n729 10.6151
R941 B.n731 B.n730 10.6151
R942 B.n731 B.n8 10.6151
R943 B.n735 B.n8 10.6151
R944 B.n736 B.n735 10.6151
R945 B.n737 B.n736 10.6151
R946 B.n737 B.n6 10.6151
R947 B.n741 B.n6 10.6151
R948 B.n742 B.n741 10.6151
R949 B.n743 B.n742 10.6151
R950 B.n743 B.n4 10.6151
R951 B.n747 B.n4 10.6151
R952 B.n748 B.n747 10.6151
R953 B.n749 B.n748 10.6151
R954 B.n749 B.n0 10.6151
R955 B.n676 B.n675 10.6151
R956 B.n675 B.n28 10.6151
R957 B.n671 B.n28 10.6151
R958 B.n671 B.n670 10.6151
R959 B.n670 B.n669 10.6151
R960 B.n669 B.n30 10.6151
R961 B.n665 B.n30 10.6151
R962 B.n665 B.n664 10.6151
R963 B.n664 B.n663 10.6151
R964 B.n663 B.n32 10.6151
R965 B.n659 B.n32 10.6151
R966 B.n659 B.n658 10.6151
R967 B.n658 B.n657 10.6151
R968 B.n657 B.n34 10.6151
R969 B.n653 B.n34 10.6151
R970 B.n653 B.n652 10.6151
R971 B.n652 B.n651 10.6151
R972 B.n651 B.n36 10.6151
R973 B.n647 B.n36 10.6151
R974 B.n647 B.n646 10.6151
R975 B.n646 B.n645 10.6151
R976 B.n645 B.n38 10.6151
R977 B.n641 B.n38 10.6151
R978 B.n641 B.n640 10.6151
R979 B.n640 B.n639 10.6151
R980 B.n639 B.n40 10.6151
R981 B.n635 B.n40 10.6151
R982 B.n635 B.n634 10.6151
R983 B.n634 B.n633 10.6151
R984 B.n633 B.n42 10.6151
R985 B.n629 B.n42 10.6151
R986 B.n629 B.n628 10.6151
R987 B.n628 B.n627 10.6151
R988 B.n627 B.n44 10.6151
R989 B.n623 B.n44 10.6151
R990 B.n623 B.n622 10.6151
R991 B.n620 B.n48 10.6151
R992 B.n616 B.n48 10.6151
R993 B.n616 B.n615 10.6151
R994 B.n615 B.n614 10.6151
R995 B.n614 B.n50 10.6151
R996 B.n610 B.n50 10.6151
R997 B.n610 B.n609 10.6151
R998 B.n609 B.n608 10.6151
R999 B.n608 B.n52 10.6151
R1000 B.n604 B.n603 10.6151
R1001 B.n603 B.n602 10.6151
R1002 B.n602 B.n57 10.6151
R1003 B.n598 B.n57 10.6151
R1004 B.n598 B.n597 10.6151
R1005 B.n597 B.n596 10.6151
R1006 B.n596 B.n59 10.6151
R1007 B.n592 B.n59 10.6151
R1008 B.n592 B.n591 10.6151
R1009 B.n591 B.n590 10.6151
R1010 B.n590 B.n61 10.6151
R1011 B.n586 B.n61 10.6151
R1012 B.n586 B.n585 10.6151
R1013 B.n585 B.n584 10.6151
R1014 B.n584 B.n63 10.6151
R1015 B.n580 B.n63 10.6151
R1016 B.n580 B.n579 10.6151
R1017 B.n579 B.n578 10.6151
R1018 B.n578 B.n65 10.6151
R1019 B.n574 B.n65 10.6151
R1020 B.n574 B.n573 10.6151
R1021 B.n573 B.n572 10.6151
R1022 B.n572 B.n67 10.6151
R1023 B.n568 B.n67 10.6151
R1024 B.n568 B.n567 10.6151
R1025 B.n567 B.n566 10.6151
R1026 B.n566 B.n69 10.6151
R1027 B.n562 B.n69 10.6151
R1028 B.n562 B.n561 10.6151
R1029 B.n561 B.n560 10.6151
R1030 B.n560 B.n71 10.6151
R1031 B.n556 B.n71 10.6151
R1032 B.n556 B.n555 10.6151
R1033 B.n555 B.n554 10.6151
R1034 B.n554 B.n73 10.6151
R1035 B.n550 B.n73 10.6151
R1036 B.n549 B.n548 10.6151
R1037 B.n548 B.n75 10.6151
R1038 B.n544 B.n75 10.6151
R1039 B.n544 B.n543 10.6151
R1040 B.n543 B.n542 10.6151
R1041 B.n542 B.n77 10.6151
R1042 B.n538 B.n77 10.6151
R1043 B.n538 B.n537 10.6151
R1044 B.n537 B.n536 10.6151
R1045 B.n536 B.n79 10.6151
R1046 B.n532 B.n79 10.6151
R1047 B.n532 B.n531 10.6151
R1048 B.n531 B.n530 10.6151
R1049 B.n530 B.n81 10.6151
R1050 B.n526 B.n81 10.6151
R1051 B.n526 B.n525 10.6151
R1052 B.n525 B.n524 10.6151
R1053 B.n524 B.n83 10.6151
R1054 B.n520 B.n83 10.6151
R1055 B.n520 B.n519 10.6151
R1056 B.n519 B.n518 10.6151
R1057 B.n518 B.n85 10.6151
R1058 B.n514 B.n85 10.6151
R1059 B.n514 B.n513 10.6151
R1060 B.n513 B.n512 10.6151
R1061 B.n512 B.n87 10.6151
R1062 B.n508 B.n87 10.6151
R1063 B.n508 B.n507 10.6151
R1064 B.n507 B.n506 10.6151
R1065 B.n506 B.n89 10.6151
R1066 B.n502 B.n89 10.6151
R1067 B.n502 B.n501 10.6151
R1068 B.n501 B.n500 10.6151
R1069 B.n500 B.n91 10.6151
R1070 B.n496 B.n91 10.6151
R1071 B.n496 B.n495 10.6151
R1072 B.n495 B.n494 10.6151
R1073 B.n494 B.n93 10.6151
R1074 B.n490 B.n93 10.6151
R1075 B.n490 B.n489 10.6151
R1076 B.n489 B.n488 10.6151
R1077 B.n488 B.n95 10.6151
R1078 B.n484 B.n95 10.6151
R1079 B.n484 B.n483 10.6151
R1080 B.n483 B.n482 10.6151
R1081 B.n482 B.n97 10.6151
R1082 B.n478 B.n97 10.6151
R1083 B.n478 B.n477 10.6151
R1084 B.n477 B.n476 10.6151
R1085 B.n476 B.n99 10.6151
R1086 B.n472 B.n99 10.6151
R1087 B.n472 B.n471 10.6151
R1088 B.n471 B.n470 10.6151
R1089 B.n470 B.n101 10.6151
R1090 B.n466 B.n101 10.6151
R1091 B.n466 B.n465 10.6151
R1092 B.n465 B.n464 10.6151
R1093 B.n464 B.n103 10.6151
R1094 B.n460 B.n103 10.6151
R1095 B.n460 B.n459 10.6151
R1096 B.n459 B.n458 10.6151
R1097 B.n458 B.n105 10.6151
R1098 B.n454 B.n105 10.6151
R1099 B.n454 B.n453 10.6151
R1100 B.n453 B.n452 10.6151
R1101 B.n452 B.n107 10.6151
R1102 B.n448 B.n107 10.6151
R1103 B.n448 B.n447 10.6151
R1104 B.n447 B.n446 10.6151
R1105 B.n446 B.n109 10.6151
R1106 B.n442 B.n109 10.6151
R1107 B.n442 B.n441 10.6151
R1108 B.n441 B.n440 10.6151
R1109 B.n440 B.n111 10.6151
R1110 B.n436 B.n111 10.6151
R1111 B.n436 B.n435 10.6151
R1112 B.n435 B.n434 10.6151
R1113 B.n434 B.n113 10.6151
R1114 B.n430 B.n113 10.6151
R1115 B.n430 B.n429 10.6151
R1116 B.n429 B.n428 10.6151
R1117 B.n428 B.n115 10.6151
R1118 B.n424 B.n115 10.6151
R1119 B.n424 B.n423 10.6151
R1120 B.n423 B.n422 10.6151
R1121 B.n422 B.n117 10.6151
R1122 B.n418 B.n117 10.6151
R1123 B.n418 B.n417 10.6151
R1124 B.n417 B.n416 10.6151
R1125 B.n416 B.n119 10.6151
R1126 B.n412 B.n119 10.6151
R1127 B.n412 B.n411 10.6151
R1128 B.n411 B.n410 10.6151
R1129 B.n410 B.n121 10.6151
R1130 B.n406 B.n121 10.6151
R1131 B.n406 B.n405 10.6151
R1132 B.n405 B.n404 10.6151
R1133 B.n404 B.n123 10.6151
R1134 B.n400 B.n123 10.6151
R1135 B.n400 B.n399 10.6151
R1136 B.n399 B.n398 10.6151
R1137 B.n193 B.n1 10.6151
R1138 B.n196 B.n193 10.6151
R1139 B.n197 B.n196 10.6151
R1140 B.n198 B.n197 10.6151
R1141 B.n198 B.n191 10.6151
R1142 B.n202 B.n191 10.6151
R1143 B.n203 B.n202 10.6151
R1144 B.n204 B.n203 10.6151
R1145 B.n204 B.n189 10.6151
R1146 B.n208 B.n189 10.6151
R1147 B.n209 B.n208 10.6151
R1148 B.n210 B.n209 10.6151
R1149 B.n210 B.n187 10.6151
R1150 B.n214 B.n187 10.6151
R1151 B.n215 B.n214 10.6151
R1152 B.n216 B.n215 10.6151
R1153 B.n216 B.n185 10.6151
R1154 B.n220 B.n185 10.6151
R1155 B.n221 B.n220 10.6151
R1156 B.n222 B.n221 10.6151
R1157 B.n222 B.n183 10.6151
R1158 B.n226 B.n183 10.6151
R1159 B.n227 B.n226 10.6151
R1160 B.n228 B.n227 10.6151
R1161 B.n228 B.n181 10.6151
R1162 B.n232 B.n181 10.6151
R1163 B.n233 B.n232 10.6151
R1164 B.n234 B.n233 10.6151
R1165 B.n234 B.n179 10.6151
R1166 B.n238 B.n179 10.6151
R1167 B.n239 B.n238 10.6151
R1168 B.n240 B.n239 10.6151
R1169 B.n240 B.n177 10.6151
R1170 B.n244 B.n177 10.6151
R1171 B.n245 B.n244 10.6151
R1172 B.n246 B.n245 10.6151
R1173 B.n246 B.n175 10.6151
R1174 B.n250 B.n175 10.6151
R1175 B.n251 B.n250 10.6151
R1176 B.n252 B.n251 10.6151
R1177 B.n252 B.n173 10.6151
R1178 B.n256 B.n173 10.6151
R1179 B.n257 B.n256 10.6151
R1180 B.n258 B.n257 10.6151
R1181 B.n258 B.n171 10.6151
R1182 B.n262 B.n171 10.6151
R1183 B.n263 B.n262 10.6151
R1184 B.n264 B.n263 10.6151
R1185 B.n264 B.n169 10.6151
R1186 B.n269 B.n268 10.6151
R1187 B.n270 B.n269 10.6151
R1188 B.n270 B.n167 10.6151
R1189 B.n274 B.n167 10.6151
R1190 B.n275 B.n274 10.6151
R1191 B.n276 B.n275 10.6151
R1192 B.n276 B.n165 10.6151
R1193 B.n280 B.n165 10.6151
R1194 B.n281 B.n280 10.6151
R1195 B.n282 B.n281 10.6151
R1196 B.n282 B.n163 10.6151
R1197 B.n286 B.n163 10.6151
R1198 B.n287 B.n286 10.6151
R1199 B.n288 B.n287 10.6151
R1200 B.n288 B.n161 10.6151
R1201 B.n292 B.n161 10.6151
R1202 B.n293 B.n292 10.6151
R1203 B.n294 B.n293 10.6151
R1204 B.n294 B.n159 10.6151
R1205 B.n298 B.n159 10.6151
R1206 B.n299 B.n298 10.6151
R1207 B.n300 B.n299 10.6151
R1208 B.n300 B.n157 10.6151
R1209 B.n304 B.n157 10.6151
R1210 B.n305 B.n304 10.6151
R1211 B.n306 B.n305 10.6151
R1212 B.n306 B.n155 10.6151
R1213 B.n310 B.n155 10.6151
R1214 B.n311 B.n310 10.6151
R1215 B.n312 B.n311 10.6151
R1216 B.n312 B.n153 10.6151
R1217 B.n316 B.n153 10.6151
R1218 B.n317 B.n316 10.6151
R1219 B.n318 B.n317 10.6151
R1220 B.n318 B.n151 10.6151
R1221 B.n322 B.n151 10.6151
R1222 B.n325 B.n324 10.6151
R1223 B.n325 B.n147 10.6151
R1224 B.n329 B.n147 10.6151
R1225 B.n330 B.n329 10.6151
R1226 B.n331 B.n330 10.6151
R1227 B.n331 B.n145 10.6151
R1228 B.n335 B.n145 10.6151
R1229 B.n336 B.n335 10.6151
R1230 B.n340 B.n336 10.6151
R1231 B.n344 B.n143 10.6151
R1232 B.n345 B.n344 10.6151
R1233 B.n346 B.n345 10.6151
R1234 B.n346 B.n141 10.6151
R1235 B.n350 B.n141 10.6151
R1236 B.n351 B.n350 10.6151
R1237 B.n352 B.n351 10.6151
R1238 B.n352 B.n139 10.6151
R1239 B.n356 B.n139 10.6151
R1240 B.n357 B.n356 10.6151
R1241 B.n358 B.n357 10.6151
R1242 B.n358 B.n137 10.6151
R1243 B.n362 B.n137 10.6151
R1244 B.n363 B.n362 10.6151
R1245 B.n364 B.n363 10.6151
R1246 B.n364 B.n135 10.6151
R1247 B.n368 B.n135 10.6151
R1248 B.n369 B.n368 10.6151
R1249 B.n370 B.n369 10.6151
R1250 B.n370 B.n133 10.6151
R1251 B.n374 B.n133 10.6151
R1252 B.n375 B.n374 10.6151
R1253 B.n376 B.n375 10.6151
R1254 B.n376 B.n131 10.6151
R1255 B.n380 B.n131 10.6151
R1256 B.n381 B.n380 10.6151
R1257 B.n382 B.n381 10.6151
R1258 B.n382 B.n129 10.6151
R1259 B.n386 B.n129 10.6151
R1260 B.n387 B.n386 10.6151
R1261 B.n388 B.n387 10.6151
R1262 B.n388 B.n127 10.6151
R1263 B.n392 B.n127 10.6151
R1264 B.n393 B.n392 10.6151
R1265 B.n394 B.n393 10.6151
R1266 B.n394 B.n125 10.6151
R1267 B.n622 B.n621 9.36635
R1268 B.n604 B.n56 9.36635
R1269 B.n323 B.n322 9.36635
R1270 B.n339 B.n143 9.36635
R1271 B.n753 B.n0 8.11757
R1272 B.n753 B.n1 8.11757
R1273 B.n621 B.n620 1.24928
R1274 B.n56 B.n52 1.24928
R1275 B.n324 B.n323 1.24928
R1276 B.n340 B.n339 1.24928
R1277 VP.n19 VP.n16 161.3
R1278 VP.n21 VP.n20 161.3
R1279 VP.n22 VP.n15 161.3
R1280 VP.n24 VP.n23 161.3
R1281 VP.n25 VP.n14 161.3
R1282 VP.n27 VP.n26 161.3
R1283 VP.n29 VP.n28 161.3
R1284 VP.n30 VP.n12 161.3
R1285 VP.n32 VP.n31 161.3
R1286 VP.n33 VP.n11 161.3
R1287 VP.n35 VP.n34 161.3
R1288 VP.n36 VP.n10 161.3
R1289 VP.n68 VP.n0 161.3
R1290 VP.n67 VP.n66 161.3
R1291 VP.n65 VP.n1 161.3
R1292 VP.n64 VP.n63 161.3
R1293 VP.n62 VP.n2 161.3
R1294 VP.n61 VP.n60 161.3
R1295 VP.n59 VP.n58 161.3
R1296 VP.n57 VP.n4 161.3
R1297 VP.n56 VP.n55 161.3
R1298 VP.n54 VP.n5 161.3
R1299 VP.n53 VP.n52 161.3
R1300 VP.n51 VP.n6 161.3
R1301 VP.n49 VP.n48 161.3
R1302 VP.n47 VP.n7 161.3
R1303 VP.n46 VP.n45 161.3
R1304 VP.n44 VP.n8 161.3
R1305 VP.n43 VP.n42 161.3
R1306 VP.n41 VP.n9 161.3
R1307 VP.n17 VP.t1 130.329
R1308 VP.n40 VP.n39 107.928
R1309 VP.n70 VP.n69 107.928
R1310 VP.n38 VP.n37 107.928
R1311 VP.n39 VP.t6 99.247
R1312 VP.n50 VP.t5 99.247
R1313 VP.n3 VP.t3 99.247
R1314 VP.n69 VP.t2 99.247
R1315 VP.n37 VP.t4 99.247
R1316 VP.n13 VP.t0 99.247
R1317 VP.n18 VP.t7 99.247
R1318 VP.n18 VP.n17 63.2583
R1319 VP.n56 VP.n5 56.4773
R1320 VP.n24 VP.n15 56.4773
R1321 VP.n45 VP.n44 52.0954
R1322 VP.n63 VP.n1 52.0954
R1323 VP.n31 VP.n11 52.0954
R1324 VP.n40 VP.n38 49.3404
R1325 VP.n45 VP.n7 28.7258
R1326 VP.n63 VP.n62 28.7258
R1327 VP.n31 VP.n30 28.7258
R1328 VP.n43 VP.n9 24.3439
R1329 VP.n44 VP.n43 24.3439
R1330 VP.n49 VP.n7 24.3439
R1331 VP.n52 VP.n51 24.3439
R1332 VP.n52 VP.n5 24.3439
R1333 VP.n57 VP.n56 24.3439
R1334 VP.n58 VP.n57 24.3439
R1335 VP.n62 VP.n61 24.3439
R1336 VP.n67 VP.n1 24.3439
R1337 VP.n68 VP.n67 24.3439
R1338 VP.n35 VP.n11 24.3439
R1339 VP.n36 VP.n35 24.3439
R1340 VP.n25 VP.n24 24.3439
R1341 VP.n26 VP.n25 24.3439
R1342 VP.n30 VP.n29 24.3439
R1343 VP.n20 VP.n19 24.3439
R1344 VP.n20 VP.n15 24.3439
R1345 VP.n50 VP.n49 15.3369
R1346 VP.n61 VP.n3 15.3369
R1347 VP.n29 VP.n13 15.3369
R1348 VP.n51 VP.n50 9.00757
R1349 VP.n58 VP.n3 9.00757
R1350 VP.n26 VP.n13 9.00757
R1351 VP.n19 VP.n18 9.00757
R1352 VP.n17 VP.n16 7.32939
R1353 VP.n39 VP.n9 2.67828
R1354 VP.n69 VP.n68 2.67828
R1355 VP.n37 VP.n36 2.67828
R1356 VP.n38 VP.n10 0.278398
R1357 VP.n41 VP.n40 0.278398
R1358 VP.n70 VP.n0 0.278398
R1359 VP.n21 VP.n16 0.189894
R1360 VP.n22 VP.n21 0.189894
R1361 VP.n23 VP.n22 0.189894
R1362 VP.n23 VP.n14 0.189894
R1363 VP.n27 VP.n14 0.189894
R1364 VP.n28 VP.n27 0.189894
R1365 VP.n28 VP.n12 0.189894
R1366 VP.n32 VP.n12 0.189894
R1367 VP.n33 VP.n32 0.189894
R1368 VP.n34 VP.n33 0.189894
R1369 VP.n34 VP.n10 0.189894
R1370 VP.n42 VP.n41 0.189894
R1371 VP.n42 VP.n8 0.189894
R1372 VP.n46 VP.n8 0.189894
R1373 VP.n47 VP.n46 0.189894
R1374 VP.n48 VP.n47 0.189894
R1375 VP.n48 VP.n6 0.189894
R1376 VP.n53 VP.n6 0.189894
R1377 VP.n54 VP.n53 0.189894
R1378 VP.n55 VP.n54 0.189894
R1379 VP.n55 VP.n4 0.189894
R1380 VP.n59 VP.n4 0.189894
R1381 VP.n60 VP.n59 0.189894
R1382 VP.n60 VP.n2 0.189894
R1383 VP.n64 VP.n2 0.189894
R1384 VP.n65 VP.n64 0.189894
R1385 VP.n66 VP.n65 0.189894
R1386 VP.n66 VP.n0 0.189894
R1387 VP VP.n70 0.153422
R1388 VDD1 VDD1.n0 80.4791
R1389 VDD1.n3 VDD1.n2 80.3653
R1390 VDD1.n3 VDD1.n1 80.3653
R1391 VDD1.n5 VDD1.n4 79.1837
R1392 VDD1.n5 VDD1.n3 44.4492
R1393 VDD1.n4 VDD1.t7 3.10805
R1394 VDD1.n4 VDD1.t3 3.10805
R1395 VDD1.n0 VDD1.t6 3.10805
R1396 VDD1.n0 VDD1.t0 3.10805
R1397 VDD1.n2 VDD1.t4 3.10805
R1398 VDD1.n2 VDD1.t5 3.10805
R1399 VDD1.n1 VDD1.t1 3.10805
R1400 VDD1.n1 VDD1.t2 3.10805
R1401 VDD1 VDD1.n5 1.17938
C0 w_n3840_n3060# VTAIL 3.86347f
C1 VP VDD2 0.51288f
C2 B VN 1.18945f
C3 VDD1 VN 0.151213f
C4 VP w_n3840_n3060# 8.28706f
C5 B VDD1 1.58836f
C6 VP VTAIL 8.053619f
C7 VN VDD2 7.59865f
C8 B VDD2 1.6825f
C9 VDD1 VDD2 1.74561f
C10 w_n3840_n3060# VN 7.78873f
C11 B w_n3840_n3060# 9.59226f
C12 VTAIL VN 8.03951f
C13 B VTAIL 4.45223f
C14 VDD1 w_n3840_n3060# 1.89383f
C15 VDD1 VTAIL 7.5435f
C16 VP VN 7.31458f
C17 B VP 2.02451f
C18 w_n3840_n3060# VDD2 2.00602f
C19 VDD1 VP 7.95895f
C20 VTAIL VDD2 7.597519f
C21 VDD2 VSUBS 1.835193f
C22 VDD1 VSUBS 2.355709f
C23 VTAIL VSUBS 1.257576f
C24 VN VSUBS 6.60199f
C25 VP VSUBS 3.462167f
C26 B VSUBS 4.809645f
C27 w_n3840_n3060# VSUBS 0.145014p
C28 VDD1.t6 VSUBS 0.203641f
C29 VDD1.t0 VSUBS 0.203641f
C30 VDD1.n0 VSUBS 1.57052f
C31 VDD1.t1 VSUBS 0.203641f
C32 VDD1.t2 VSUBS 0.203641f
C33 VDD1.n1 VSUBS 1.56935f
C34 VDD1.t4 VSUBS 0.203641f
C35 VDD1.t5 VSUBS 0.203641f
C36 VDD1.n2 VSUBS 1.56935f
C37 VDD1.n3 VSUBS 3.62798f
C38 VDD1.t7 VSUBS 0.203641f
C39 VDD1.t3 VSUBS 0.203641f
C40 VDD1.n4 VSUBS 1.55842f
C41 VDD1.n5 VSUBS 3.03984f
C42 VP.n0 VSUBS 0.044313f
C43 VP.t2 VSUBS 2.42271f
C44 VP.n1 VSUBS 0.060635f
C45 VP.n2 VSUBS 0.033609f
C46 VP.t3 VSUBS 2.42271f
C47 VP.n3 VSUBS 0.865234f
C48 VP.n4 VSUBS 0.033609f
C49 VP.n5 VSUBS 0.049277f
C50 VP.n6 VSUBS 0.033609f
C51 VP.t5 VSUBS 2.42271f
C52 VP.n7 VSUBS 0.066841f
C53 VP.n8 VSUBS 0.033609f
C54 VP.n9 VSUBS 0.03529f
C55 VP.n10 VSUBS 0.044313f
C56 VP.t4 VSUBS 2.42271f
C57 VP.n11 VSUBS 0.060635f
C58 VP.n12 VSUBS 0.033609f
C59 VP.t0 VSUBS 2.42271f
C60 VP.n13 VSUBS 0.865234f
C61 VP.n14 VSUBS 0.033609f
C62 VP.n15 VSUBS 0.049277f
C63 VP.n16 VSUBS 0.321833f
C64 VP.t7 VSUBS 2.42271f
C65 VP.t1 VSUBS 2.67732f
C66 VP.n17 VSUBS 0.944644f
C67 VP.n18 VSUBS 0.957983f
C68 VP.n19 VSUBS 0.043371f
C69 VP.n20 VSUBS 0.062953f
C70 VP.n21 VSUBS 0.033609f
C71 VP.n22 VSUBS 0.033609f
C72 VP.n23 VSUBS 0.033609f
C73 VP.n24 VSUBS 0.049277f
C74 VP.n25 VSUBS 0.062953f
C75 VP.n26 VSUBS 0.043371f
C76 VP.n27 VSUBS 0.033609f
C77 VP.n28 VSUBS 0.033609f
C78 VP.n29 VSUBS 0.051453f
C79 VP.n30 VSUBS 0.066841f
C80 VP.n31 VSUBS 0.034031f
C81 VP.n32 VSUBS 0.033609f
C82 VP.n33 VSUBS 0.033609f
C83 VP.n34 VSUBS 0.033609f
C84 VP.n35 VSUBS 0.062953f
C85 VP.n36 VSUBS 0.03529f
C86 VP.n37 VSUBS 0.963011f
C87 VP.n38 VSUBS 1.83683f
C88 VP.t6 VSUBS 2.42271f
C89 VP.n39 VSUBS 0.963011f
C90 VP.n40 VSUBS 1.86124f
C91 VP.n41 VSUBS 0.044313f
C92 VP.n42 VSUBS 0.033609f
C93 VP.n43 VSUBS 0.062953f
C94 VP.n44 VSUBS 0.060635f
C95 VP.n45 VSUBS 0.034031f
C96 VP.n46 VSUBS 0.033609f
C97 VP.n47 VSUBS 0.033609f
C98 VP.n48 VSUBS 0.033609f
C99 VP.n49 VSUBS 0.051453f
C100 VP.n50 VSUBS 0.865234f
C101 VP.n51 VSUBS 0.043371f
C102 VP.n52 VSUBS 0.062953f
C103 VP.n53 VSUBS 0.033609f
C104 VP.n54 VSUBS 0.033609f
C105 VP.n55 VSUBS 0.033609f
C106 VP.n56 VSUBS 0.049277f
C107 VP.n57 VSUBS 0.062953f
C108 VP.n58 VSUBS 0.043371f
C109 VP.n59 VSUBS 0.033609f
C110 VP.n60 VSUBS 0.033609f
C111 VP.n61 VSUBS 0.051453f
C112 VP.n62 VSUBS 0.066841f
C113 VP.n63 VSUBS 0.034031f
C114 VP.n64 VSUBS 0.033609f
C115 VP.n65 VSUBS 0.033609f
C116 VP.n66 VSUBS 0.033609f
C117 VP.n67 VSUBS 0.062953f
C118 VP.n68 VSUBS 0.03529f
C119 VP.n69 VSUBS 0.963011f
C120 VP.n70 VSUBS 0.059342f
C121 B.n0 VSUBS 0.007066f
C122 B.n1 VSUBS 0.007066f
C123 B.n2 VSUBS 0.010451f
C124 B.n3 VSUBS 0.008009f
C125 B.n4 VSUBS 0.008009f
C126 B.n5 VSUBS 0.008009f
C127 B.n6 VSUBS 0.008009f
C128 B.n7 VSUBS 0.008009f
C129 B.n8 VSUBS 0.008009f
C130 B.n9 VSUBS 0.008009f
C131 B.n10 VSUBS 0.008009f
C132 B.n11 VSUBS 0.008009f
C133 B.n12 VSUBS 0.008009f
C134 B.n13 VSUBS 0.008009f
C135 B.n14 VSUBS 0.008009f
C136 B.n15 VSUBS 0.008009f
C137 B.n16 VSUBS 0.008009f
C138 B.n17 VSUBS 0.008009f
C139 B.n18 VSUBS 0.008009f
C140 B.n19 VSUBS 0.008009f
C141 B.n20 VSUBS 0.008009f
C142 B.n21 VSUBS 0.008009f
C143 B.n22 VSUBS 0.008009f
C144 B.n23 VSUBS 0.008009f
C145 B.n24 VSUBS 0.008009f
C146 B.n25 VSUBS 0.008009f
C147 B.n26 VSUBS 0.008009f
C148 B.n27 VSUBS 0.017882f
C149 B.n28 VSUBS 0.008009f
C150 B.n29 VSUBS 0.008009f
C151 B.n30 VSUBS 0.008009f
C152 B.n31 VSUBS 0.008009f
C153 B.n32 VSUBS 0.008009f
C154 B.n33 VSUBS 0.008009f
C155 B.n34 VSUBS 0.008009f
C156 B.n35 VSUBS 0.008009f
C157 B.n36 VSUBS 0.008009f
C158 B.n37 VSUBS 0.008009f
C159 B.n38 VSUBS 0.008009f
C160 B.n39 VSUBS 0.008009f
C161 B.n40 VSUBS 0.008009f
C162 B.n41 VSUBS 0.008009f
C163 B.n42 VSUBS 0.008009f
C164 B.n43 VSUBS 0.008009f
C165 B.n44 VSUBS 0.008009f
C166 B.n45 VSUBS 0.008009f
C167 B.t10 VSUBS 0.383843f
C168 B.t11 VSUBS 0.407105f
C169 B.t9 VSUBS 1.39395f
C170 B.n46 VSUBS 0.21293f
C171 B.n47 VSUBS 0.081726f
C172 B.n48 VSUBS 0.008009f
C173 B.n49 VSUBS 0.008009f
C174 B.n50 VSUBS 0.008009f
C175 B.n51 VSUBS 0.008009f
C176 B.n52 VSUBS 0.004475f
C177 B.n53 VSUBS 0.008009f
C178 B.t7 VSUBS 0.383837f
C179 B.t8 VSUBS 0.4071f
C180 B.t6 VSUBS 1.39395f
C181 B.n54 VSUBS 0.212936f
C182 B.n55 VSUBS 0.081731f
C183 B.n56 VSUBS 0.018555f
C184 B.n57 VSUBS 0.008009f
C185 B.n58 VSUBS 0.008009f
C186 B.n59 VSUBS 0.008009f
C187 B.n60 VSUBS 0.008009f
C188 B.n61 VSUBS 0.008009f
C189 B.n62 VSUBS 0.008009f
C190 B.n63 VSUBS 0.008009f
C191 B.n64 VSUBS 0.008009f
C192 B.n65 VSUBS 0.008009f
C193 B.n66 VSUBS 0.008009f
C194 B.n67 VSUBS 0.008009f
C195 B.n68 VSUBS 0.008009f
C196 B.n69 VSUBS 0.008009f
C197 B.n70 VSUBS 0.008009f
C198 B.n71 VSUBS 0.008009f
C199 B.n72 VSUBS 0.008009f
C200 B.n73 VSUBS 0.008009f
C201 B.n74 VSUBS 0.016979f
C202 B.n75 VSUBS 0.008009f
C203 B.n76 VSUBS 0.008009f
C204 B.n77 VSUBS 0.008009f
C205 B.n78 VSUBS 0.008009f
C206 B.n79 VSUBS 0.008009f
C207 B.n80 VSUBS 0.008009f
C208 B.n81 VSUBS 0.008009f
C209 B.n82 VSUBS 0.008009f
C210 B.n83 VSUBS 0.008009f
C211 B.n84 VSUBS 0.008009f
C212 B.n85 VSUBS 0.008009f
C213 B.n86 VSUBS 0.008009f
C214 B.n87 VSUBS 0.008009f
C215 B.n88 VSUBS 0.008009f
C216 B.n89 VSUBS 0.008009f
C217 B.n90 VSUBS 0.008009f
C218 B.n91 VSUBS 0.008009f
C219 B.n92 VSUBS 0.008009f
C220 B.n93 VSUBS 0.008009f
C221 B.n94 VSUBS 0.008009f
C222 B.n95 VSUBS 0.008009f
C223 B.n96 VSUBS 0.008009f
C224 B.n97 VSUBS 0.008009f
C225 B.n98 VSUBS 0.008009f
C226 B.n99 VSUBS 0.008009f
C227 B.n100 VSUBS 0.008009f
C228 B.n101 VSUBS 0.008009f
C229 B.n102 VSUBS 0.008009f
C230 B.n103 VSUBS 0.008009f
C231 B.n104 VSUBS 0.008009f
C232 B.n105 VSUBS 0.008009f
C233 B.n106 VSUBS 0.008009f
C234 B.n107 VSUBS 0.008009f
C235 B.n108 VSUBS 0.008009f
C236 B.n109 VSUBS 0.008009f
C237 B.n110 VSUBS 0.008009f
C238 B.n111 VSUBS 0.008009f
C239 B.n112 VSUBS 0.008009f
C240 B.n113 VSUBS 0.008009f
C241 B.n114 VSUBS 0.008009f
C242 B.n115 VSUBS 0.008009f
C243 B.n116 VSUBS 0.008009f
C244 B.n117 VSUBS 0.008009f
C245 B.n118 VSUBS 0.008009f
C246 B.n119 VSUBS 0.008009f
C247 B.n120 VSUBS 0.008009f
C248 B.n121 VSUBS 0.008009f
C249 B.n122 VSUBS 0.008009f
C250 B.n123 VSUBS 0.008009f
C251 B.n124 VSUBS 0.008009f
C252 B.n125 VSUBS 0.016824f
C253 B.n126 VSUBS 0.008009f
C254 B.n127 VSUBS 0.008009f
C255 B.n128 VSUBS 0.008009f
C256 B.n129 VSUBS 0.008009f
C257 B.n130 VSUBS 0.008009f
C258 B.n131 VSUBS 0.008009f
C259 B.n132 VSUBS 0.008009f
C260 B.n133 VSUBS 0.008009f
C261 B.n134 VSUBS 0.008009f
C262 B.n135 VSUBS 0.008009f
C263 B.n136 VSUBS 0.008009f
C264 B.n137 VSUBS 0.008009f
C265 B.n138 VSUBS 0.008009f
C266 B.n139 VSUBS 0.008009f
C267 B.n140 VSUBS 0.008009f
C268 B.n141 VSUBS 0.008009f
C269 B.n142 VSUBS 0.008009f
C270 B.n143 VSUBS 0.007538f
C271 B.n144 VSUBS 0.008009f
C272 B.n145 VSUBS 0.008009f
C273 B.n146 VSUBS 0.008009f
C274 B.n147 VSUBS 0.008009f
C275 B.n148 VSUBS 0.008009f
C276 B.t5 VSUBS 0.383843f
C277 B.t4 VSUBS 0.407105f
C278 B.t3 VSUBS 1.39395f
C279 B.n149 VSUBS 0.21293f
C280 B.n150 VSUBS 0.081726f
C281 B.n151 VSUBS 0.008009f
C282 B.n152 VSUBS 0.008009f
C283 B.n153 VSUBS 0.008009f
C284 B.n154 VSUBS 0.008009f
C285 B.n155 VSUBS 0.008009f
C286 B.n156 VSUBS 0.008009f
C287 B.n157 VSUBS 0.008009f
C288 B.n158 VSUBS 0.008009f
C289 B.n159 VSUBS 0.008009f
C290 B.n160 VSUBS 0.008009f
C291 B.n161 VSUBS 0.008009f
C292 B.n162 VSUBS 0.008009f
C293 B.n163 VSUBS 0.008009f
C294 B.n164 VSUBS 0.008009f
C295 B.n165 VSUBS 0.008009f
C296 B.n166 VSUBS 0.008009f
C297 B.n167 VSUBS 0.008009f
C298 B.n168 VSUBS 0.008009f
C299 B.n169 VSUBS 0.016979f
C300 B.n170 VSUBS 0.008009f
C301 B.n171 VSUBS 0.008009f
C302 B.n172 VSUBS 0.008009f
C303 B.n173 VSUBS 0.008009f
C304 B.n174 VSUBS 0.008009f
C305 B.n175 VSUBS 0.008009f
C306 B.n176 VSUBS 0.008009f
C307 B.n177 VSUBS 0.008009f
C308 B.n178 VSUBS 0.008009f
C309 B.n179 VSUBS 0.008009f
C310 B.n180 VSUBS 0.008009f
C311 B.n181 VSUBS 0.008009f
C312 B.n182 VSUBS 0.008009f
C313 B.n183 VSUBS 0.008009f
C314 B.n184 VSUBS 0.008009f
C315 B.n185 VSUBS 0.008009f
C316 B.n186 VSUBS 0.008009f
C317 B.n187 VSUBS 0.008009f
C318 B.n188 VSUBS 0.008009f
C319 B.n189 VSUBS 0.008009f
C320 B.n190 VSUBS 0.008009f
C321 B.n191 VSUBS 0.008009f
C322 B.n192 VSUBS 0.008009f
C323 B.n193 VSUBS 0.008009f
C324 B.n194 VSUBS 0.008009f
C325 B.n195 VSUBS 0.008009f
C326 B.n196 VSUBS 0.008009f
C327 B.n197 VSUBS 0.008009f
C328 B.n198 VSUBS 0.008009f
C329 B.n199 VSUBS 0.008009f
C330 B.n200 VSUBS 0.008009f
C331 B.n201 VSUBS 0.008009f
C332 B.n202 VSUBS 0.008009f
C333 B.n203 VSUBS 0.008009f
C334 B.n204 VSUBS 0.008009f
C335 B.n205 VSUBS 0.008009f
C336 B.n206 VSUBS 0.008009f
C337 B.n207 VSUBS 0.008009f
C338 B.n208 VSUBS 0.008009f
C339 B.n209 VSUBS 0.008009f
C340 B.n210 VSUBS 0.008009f
C341 B.n211 VSUBS 0.008009f
C342 B.n212 VSUBS 0.008009f
C343 B.n213 VSUBS 0.008009f
C344 B.n214 VSUBS 0.008009f
C345 B.n215 VSUBS 0.008009f
C346 B.n216 VSUBS 0.008009f
C347 B.n217 VSUBS 0.008009f
C348 B.n218 VSUBS 0.008009f
C349 B.n219 VSUBS 0.008009f
C350 B.n220 VSUBS 0.008009f
C351 B.n221 VSUBS 0.008009f
C352 B.n222 VSUBS 0.008009f
C353 B.n223 VSUBS 0.008009f
C354 B.n224 VSUBS 0.008009f
C355 B.n225 VSUBS 0.008009f
C356 B.n226 VSUBS 0.008009f
C357 B.n227 VSUBS 0.008009f
C358 B.n228 VSUBS 0.008009f
C359 B.n229 VSUBS 0.008009f
C360 B.n230 VSUBS 0.008009f
C361 B.n231 VSUBS 0.008009f
C362 B.n232 VSUBS 0.008009f
C363 B.n233 VSUBS 0.008009f
C364 B.n234 VSUBS 0.008009f
C365 B.n235 VSUBS 0.008009f
C366 B.n236 VSUBS 0.008009f
C367 B.n237 VSUBS 0.008009f
C368 B.n238 VSUBS 0.008009f
C369 B.n239 VSUBS 0.008009f
C370 B.n240 VSUBS 0.008009f
C371 B.n241 VSUBS 0.008009f
C372 B.n242 VSUBS 0.008009f
C373 B.n243 VSUBS 0.008009f
C374 B.n244 VSUBS 0.008009f
C375 B.n245 VSUBS 0.008009f
C376 B.n246 VSUBS 0.008009f
C377 B.n247 VSUBS 0.008009f
C378 B.n248 VSUBS 0.008009f
C379 B.n249 VSUBS 0.008009f
C380 B.n250 VSUBS 0.008009f
C381 B.n251 VSUBS 0.008009f
C382 B.n252 VSUBS 0.008009f
C383 B.n253 VSUBS 0.008009f
C384 B.n254 VSUBS 0.008009f
C385 B.n255 VSUBS 0.008009f
C386 B.n256 VSUBS 0.008009f
C387 B.n257 VSUBS 0.008009f
C388 B.n258 VSUBS 0.008009f
C389 B.n259 VSUBS 0.008009f
C390 B.n260 VSUBS 0.008009f
C391 B.n261 VSUBS 0.008009f
C392 B.n262 VSUBS 0.008009f
C393 B.n263 VSUBS 0.008009f
C394 B.n264 VSUBS 0.008009f
C395 B.n265 VSUBS 0.008009f
C396 B.n266 VSUBS 0.016979f
C397 B.n267 VSUBS 0.017882f
C398 B.n268 VSUBS 0.017882f
C399 B.n269 VSUBS 0.008009f
C400 B.n270 VSUBS 0.008009f
C401 B.n271 VSUBS 0.008009f
C402 B.n272 VSUBS 0.008009f
C403 B.n273 VSUBS 0.008009f
C404 B.n274 VSUBS 0.008009f
C405 B.n275 VSUBS 0.008009f
C406 B.n276 VSUBS 0.008009f
C407 B.n277 VSUBS 0.008009f
C408 B.n278 VSUBS 0.008009f
C409 B.n279 VSUBS 0.008009f
C410 B.n280 VSUBS 0.008009f
C411 B.n281 VSUBS 0.008009f
C412 B.n282 VSUBS 0.008009f
C413 B.n283 VSUBS 0.008009f
C414 B.n284 VSUBS 0.008009f
C415 B.n285 VSUBS 0.008009f
C416 B.n286 VSUBS 0.008009f
C417 B.n287 VSUBS 0.008009f
C418 B.n288 VSUBS 0.008009f
C419 B.n289 VSUBS 0.008009f
C420 B.n290 VSUBS 0.008009f
C421 B.n291 VSUBS 0.008009f
C422 B.n292 VSUBS 0.008009f
C423 B.n293 VSUBS 0.008009f
C424 B.n294 VSUBS 0.008009f
C425 B.n295 VSUBS 0.008009f
C426 B.n296 VSUBS 0.008009f
C427 B.n297 VSUBS 0.008009f
C428 B.n298 VSUBS 0.008009f
C429 B.n299 VSUBS 0.008009f
C430 B.n300 VSUBS 0.008009f
C431 B.n301 VSUBS 0.008009f
C432 B.n302 VSUBS 0.008009f
C433 B.n303 VSUBS 0.008009f
C434 B.n304 VSUBS 0.008009f
C435 B.n305 VSUBS 0.008009f
C436 B.n306 VSUBS 0.008009f
C437 B.n307 VSUBS 0.008009f
C438 B.n308 VSUBS 0.008009f
C439 B.n309 VSUBS 0.008009f
C440 B.n310 VSUBS 0.008009f
C441 B.n311 VSUBS 0.008009f
C442 B.n312 VSUBS 0.008009f
C443 B.n313 VSUBS 0.008009f
C444 B.n314 VSUBS 0.008009f
C445 B.n315 VSUBS 0.008009f
C446 B.n316 VSUBS 0.008009f
C447 B.n317 VSUBS 0.008009f
C448 B.n318 VSUBS 0.008009f
C449 B.n319 VSUBS 0.008009f
C450 B.n320 VSUBS 0.008009f
C451 B.n321 VSUBS 0.008009f
C452 B.n322 VSUBS 0.007538f
C453 B.n323 VSUBS 0.018555f
C454 B.n324 VSUBS 0.004475f
C455 B.n325 VSUBS 0.008009f
C456 B.n326 VSUBS 0.008009f
C457 B.n327 VSUBS 0.008009f
C458 B.n328 VSUBS 0.008009f
C459 B.n329 VSUBS 0.008009f
C460 B.n330 VSUBS 0.008009f
C461 B.n331 VSUBS 0.008009f
C462 B.n332 VSUBS 0.008009f
C463 B.n333 VSUBS 0.008009f
C464 B.n334 VSUBS 0.008009f
C465 B.n335 VSUBS 0.008009f
C466 B.n336 VSUBS 0.008009f
C467 B.t2 VSUBS 0.383837f
C468 B.t1 VSUBS 0.4071f
C469 B.t0 VSUBS 1.39395f
C470 B.n337 VSUBS 0.212936f
C471 B.n338 VSUBS 0.081731f
C472 B.n339 VSUBS 0.018555f
C473 B.n340 VSUBS 0.004475f
C474 B.n341 VSUBS 0.008009f
C475 B.n342 VSUBS 0.008009f
C476 B.n343 VSUBS 0.008009f
C477 B.n344 VSUBS 0.008009f
C478 B.n345 VSUBS 0.008009f
C479 B.n346 VSUBS 0.008009f
C480 B.n347 VSUBS 0.008009f
C481 B.n348 VSUBS 0.008009f
C482 B.n349 VSUBS 0.008009f
C483 B.n350 VSUBS 0.008009f
C484 B.n351 VSUBS 0.008009f
C485 B.n352 VSUBS 0.008009f
C486 B.n353 VSUBS 0.008009f
C487 B.n354 VSUBS 0.008009f
C488 B.n355 VSUBS 0.008009f
C489 B.n356 VSUBS 0.008009f
C490 B.n357 VSUBS 0.008009f
C491 B.n358 VSUBS 0.008009f
C492 B.n359 VSUBS 0.008009f
C493 B.n360 VSUBS 0.008009f
C494 B.n361 VSUBS 0.008009f
C495 B.n362 VSUBS 0.008009f
C496 B.n363 VSUBS 0.008009f
C497 B.n364 VSUBS 0.008009f
C498 B.n365 VSUBS 0.008009f
C499 B.n366 VSUBS 0.008009f
C500 B.n367 VSUBS 0.008009f
C501 B.n368 VSUBS 0.008009f
C502 B.n369 VSUBS 0.008009f
C503 B.n370 VSUBS 0.008009f
C504 B.n371 VSUBS 0.008009f
C505 B.n372 VSUBS 0.008009f
C506 B.n373 VSUBS 0.008009f
C507 B.n374 VSUBS 0.008009f
C508 B.n375 VSUBS 0.008009f
C509 B.n376 VSUBS 0.008009f
C510 B.n377 VSUBS 0.008009f
C511 B.n378 VSUBS 0.008009f
C512 B.n379 VSUBS 0.008009f
C513 B.n380 VSUBS 0.008009f
C514 B.n381 VSUBS 0.008009f
C515 B.n382 VSUBS 0.008009f
C516 B.n383 VSUBS 0.008009f
C517 B.n384 VSUBS 0.008009f
C518 B.n385 VSUBS 0.008009f
C519 B.n386 VSUBS 0.008009f
C520 B.n387 VSUBS 0.008009f
C521 B.n388 VSUBS 0.008009f
C522 B.n389 VSUBS 0.008009f
C523 B.n390 VSUBS 0.008009f
C524 B.n391 VSUBS 0.008009f
C525 B.n392 VSUBS 0.008009f
C526 B.n393 VSUBS 0.008009f
C527 B.n394 VSUBS 0.008009f
C528 B.n395 VSUBS 0.008009f
C529 B.n396 VSUBS 0.017882f
C530 B.n397 VSUBS 0.016979f
C531 B.n398 VSUBS 0.018037f
C532 B.n399 VSUBS 0.008009f
C533 B.n400 VSUBS 0.008009f
C534 B.n401 VSUBS 0.008009f
C535 B.n402 VSUBS 0.008009f
C536 B.n403 VSUBS 0.008009f
C537 B.n404 VSUBS 0.008009f
C538 B.n405 VSUBS 0.008009f
C539 B.n406 VSUBS 0.008009f
C540 B.n407 VSUBS 0.008009f
C541 B.n408 VSUBS 0.008009f
C542 B.n409 VSUBS 0.008009f
C543 B.n410 VSUBS 0.008009f
C544 B.n411 VSUBS 0.008009f
C545 B.n412 VSUBS 0.008009f
C546 B.n413 VSUBS 0.008009f
C547 B.n414 VSUBS 0.008009f
C548 B.n415 VSUBS 0.008009f
C549 B.n416 VSUBS 0.008009f
C550 B.n417 VSUBS 0.008009f
C551 B.n418 VSUBS 0.008009f
C552 B.n419 VSUBS 0.008009f
C553 B.n420 VSUBS 0.008009f
C554 B.n421 VSUBS 0.008009f
C555 B.n422 VSUBS 0.008009f
C556 B.n423 VSUBS 0.008009f
C557 B.n424 VSUBS 0.008009f
C558 B.n425 VSUBS 0.008009f
C559 B.n426 VSUBS 0.008009f
C560 B.n427 VSUBS 0.008009f
C561 B.n428 VSUBS 0.008009f
C562 B.n429 VSUBS 0.008009f
C563 B.n430 VSUBS 0.008009f
C564 B.n431 VSUBS 0.008009f
C565 B.n432 VSUBS 0.008009f
C566 B.n433 VSUBS 0.008009f
C567 B.n434 VSUBS 0.008009f
C568 B.n435 VSUBS 0.008009f
C569 B.n436 VSUBS 0.008009f
C570 B.n437 VSUBS 0.008009f
C571 B.n438 VSUBS 0.008009f
C572 B.n439 VSUBS 0.008009f
C573 B.n440 VSUBS 0.008009f
C574 B.n441 VSUBS 0.008009f
C575 B.n442 VSUBS 0.008009f
C576 B.n443 VSUBS 0.008009f
C577 B.n444 VSUBS 0.008009f
C578 B.n445 VSUBS 0.008009f
C579 B.n446 VSUBS 0.008009f
C580 B.n447 VSUBS 0.008009f
C581 B.n448 VSUBS 0.008009f
C582 B.n449 VSUBS 0.008009f
C583 B.n450 VSUBS 0.008009f
C584 B.n451 VSUBS 0.008009f
C585 B.n452 VSUBS 0.008009f
C586 B.n453 VSUBS 0.008009f
C587 B.n454 VSUBS 0.008009f
C588 B.n455 VSUBS 0.008009f
C589 B.n456 VSUBS 0.008009f
C590 B.n457 VSUBS 0.008009f
C591 B.n458 VSUBS 0.008009f
C592 B.n459 VSUBS 0.008009f
C593 B.n460 VSUBS 0.008009f
C594 B.n461 VSUBS 0.008009f
C595 B.n462 VSUBS 0.008009f
C596 B.n463 VSUBS 0.008009f
C597 B.n464 VSUBS 0.008009f
C598 B.n465 VSUBS 0.008009f
C599 B.n466 VSUBS 0.008009f
C600 B.n467 VSUBS 0.008009f
C601 B.n468 VSUBS 0.008009f
C602 B.n469 VSUBS 0.008009f
C603 B.n470 VSUBS 0.008009f
C604 B.n471 VSUBS 0.008009f
C605 B.n472 VSUBS 0.008009f
C606 B.n473 VSUBS 0.008009f
C607 B.n474 VSUBS 0.008009f
C608 B.n475 VSUBS 0.008009f
C609 B.n476 VSUBS 0.008009f
C610 B.n477 VSUBS 0.008009f
C611 B.n478 VSUBS 0.008009f
C612 B.n479 VSUBS 0.008009f
C613 B.n480 VSUBS 0.008009f
C614 B.n481 VSUBS 0.008009f
C615 B.n482 VSUBS 0.008009f
C616 B.n483 VSUBS 0.008009f
C617 B.n484 VSUBS 0.008009f
C618 B.n485 VSUBS 0.008009f
C619 B.n486 VSUBS 0.008009f
C620 B.n487 VSUBS 0.008009f
C621 B.n488 VSUBS 0.008009f
C622 B.n489 VSUBS 0.008009f
C623 B.n490 VSUBS 0.008009f
C624 B.n491 VSUBS 0.008009f
C625 B.n492 VSUBS 0.008009f
C626 B.n493 VSUBS 0.008009f
C627 B.n494 VSUBS 0.008009f
C628 B.n495 VSUBS 0.008009f
C629 B.n496 VSUBS 0.008009f
C630 B.n497 VSUBS 0.008009f
C631 B.n498 VSUBS 0.008009f
C632 B.n499 VSUBS 0.008009f
C633 B.n500 VSUBS 0.008009f
C634 B.n501 VSUBS 0.008009f
C635 B.n502 VSUBS 0.008009f
C636 B.n503 VSUBS 0.008009f
C637 B.n504 VSUBS 0.008009f
C638 B.n505 VSUBS 0.008009f
C639 B.n506 VSUBS 0.008009f
C640 B.n507 VSUBS 0.008009f
C641 B.n508 VSUBS 0.008009f
C642 B.n509 VSUBS 0.008009f
C643 B.n510 VSUBS 0.008009f
C644 B.n511 VSUBS 0.008009f
C645 B.n512 VSUBS 0.008009f
C646 B.n513 VSUBS 0.008009f
C647 B.n514 VSUBS 0.008009f
C648 B.n515 VSUBS 0.008009f
C649 B.n516 VSUBS 0.008009f
C650 B.n517 VSUBS 0.008009f
C651 B.n518 VSUBS 0.008009f
C652 B.n519 VSUBS 0.008009f
C653 B.n520 VSUBS 0.008009f
C654 B.n521 VSUBS 0.008009f
C655 B.n522 VSUBS 0.008009f
C656 B.n523 VSUBS 0.008009f
C657 B.n524 VSUBS 0.008009f
C658 B.n525 VSUBS 0.008009f
C659 B.n526 VSUBS 0.008009f
C660 B.n527 VSUBS 0.008009f
C661 B.n528 VSUBS 0.008009f
C662 B.n529 VSUBS 0.008009f
C663 B.n530 VSUBS 0.008009f
C664 B.n531 VSUBS 0.008009f
C665 B.n532 VSUBS 0.008009f
C666 B.n533 VSUBS 0.008009f
C667 B.n534 VSUBS 0.008009f
C668 B.n535 VSUBS 0.008009f
C669 B.n536 VSUBS 0.008009f
C670 B.n537 VSUBS 0.008009f
C671 B.n538 VSUBS 0.008009f
C672 B.n539 VSUBS 0.008009f
C673 B.n540 VSUBS 0.008009f
C674 B.n541 VSUBS 0.008009f
C675 B.n542 VSUBS 0.008009f
C676 B.n543 VSUBS 0.008009f
C677 B.n544 VSUBS 0.008009f
C678 B.n545 VSUBS 0.008009f
C679 B.n546 VSUBS 0.008009f
C680 B.n547 VSUBS 0.008009f
C681 B.n548 VSUBS 0.008009f
C682 B.n549 VSUBS 0.016979f
C683 B.n550 VSUBS 0.017882f
C684 B.n551 VSUBS 0.017882f
C685 B.n552 VSUBS 0.008009f
C686 B.n553 VSUBS 0.008009f
C687 B.n554 VSUBS 0.008009f
C688 B.n555 VSUBS 0.008009f
C689 B.n556 VSUBS 0.008009f
C690 B.n557 VSUBS 0.008009f
C691 B.n558 VSUBS 0.008009f
C692 B.n559 VSUBS 0.008009f
C693 B.n560 VSUBS 0.008009f
C694 B.n561 VSUBS 0.008009f
C695 B.n562 VSUBS 0.008009f
C696 B.n563 VSUBS 0.008009f
C697 B.n564 VSUBS 0.008009f
C698 B.n565 VSUBS 0.008009f
C699 B.n566 VSUBS 0.008009f
C700 B.n567 VSUBS 0.008009f
C701 B.n568 VSUBS 0.008009f
C702 B.n569 VSUBS 0.008009f
C703 B.n570 VSUBS 0.008009f
C704 B.n571 VSUBS 0.008009f
C705 B.n572 VSUBS 0.008009f
C706 B.n573 VSUBS 0.008009f
C707 B.n574 VSUBS 0.008009f
C708 B.n575 VSUBS 0.008009f
C709 B.n576 VSUBS 0.008009f
C710 B.n577 VSUBS 0.008009f
C711 B.n578 VSUBS 0.008009f
C712 B.n579 VSUBS 0.008009f
C713 B.n580 VSUBS 0.008009f
C714 B.n581 VSUBS 0.008009f
C715 B.n582 VSUBS 0.008009f
C716 B.n583 VSUBS 0.008009f
C717 B.n584 VSUBS 0.008009f
C718 B.n585 VSUBS 0.008009f
C719 B.n586 VSUBS 0.008009f
C720 B.n587 VSUBS 0.008009f
C721 B.n588 VSUBS 0.008009f
C722 B.n589 VSUBS 0.008009f
C723 B.n590 VSUBS 0.008009f
C724 B.n591 VSUBS 0.008009f
C725 B.n592 VSUBS 0.008009f
C726 B.n593 VSUBS 0.008009f
C727 B.n594 VSUBS 0.008009f
C728 B.n595 VSUBS 0.008009f
C729 B.n596 VSUBS 0.008009f
C730 B.n597 VSUBS 0.008009f
C731 B.n598 VSUBS 0.008009f
C732 B.n599 VSUBS 0.008009f
C733 B.n600 VSUBS 0.008009f
C734 B.n601 VSUBS 0.008009f
C735 B.n602 VSUBS 0.008009f
C736 B.n603 VSUBS 0.008009f
C737 B.n604 VSUBS 0.007538f
C738 B.n605 VSUBS 0.008009f
C739 B.n606 VSUBS 0.008009f
C740 B.n607 VSUBS 0.008009f
C741 B.n608 VSUBS 0.008009f
C742 B.n609 VSUBS 0.008009f
C743 B.n610 VSUBS 0.008009f
C744 B.n611 VSUBS 0.008009f
C745 B.n612 VSUBS 0.008009f
C746 B.n613 VSUBS 0.008009f
C747 B.n614 VSUBS 0.008009f
C748 B.n615 VSUBS 0.008009f
C749 B.n616 VSUBS 0.008009f
C750 B.n617 VSUBS 0.008009f
C751 B.n618 VSUBS 0.008009f
C752 B.n619 VSUBS 0.008009f
C753 B.n620 VSUBS 0.004475f
C754 B.n621 VSUBS 0.018555f
C755 B.n622 VSUBS 0.007538f
C756 B.n623 VSUBS 0.008009f
C757 B.n624 VSUBS 0.008009f
C758 B.n625 VSUBS 0.008009f
C759 B.n626 VSUBS 0.008009f
C760 B.n627 VSUBS 0.008009f
C761 B.n628 VSUBS 0.008009f
C762 B.n629 VSUBS 0.008009f
C763 B.n630 VSUBS 0.008009f
C764 B.n631 VSUBS 0.008009f
C765 B.n632 VSUBS 0.008009f
C766 B.n633 VSUBS 0.008009f
C767 B.n634 VSUBS 0.008009f
C768 B.n635 VSUBS 0.008009f
C769 B.n636 VSUBS 0.008009f
C770 B.n637 VSUBS 0.008009f
C771 B.n638 VSUBS 0.008009f
C772 B.n639 VSUBS 0.008009f
C773 B.n640 VSUBS 0.008009f
C774 B.n641 VSUBS 0.008009f
C775 B.n642 VSUBS 0.008009f
C776 B.n643 VSUBS 0.008009f
C777 B.n644 VSUBS 0.008009f
C778 B.n645 VSUBS 0.008009f
C779 B.n646 VSUBS 0.008009f
C780 B.n647 VSUBS 0.008009f
C781 B.n648 VSUBS 0.008009f
C782 B.n649 VSUBS 0.008009f
C783 B.n650 VSUBS 0.008009f
C784 B.n651 VSUBS 0.008009f
C785 B.n652 VSUBS 0.008009f
C786 B.n653 VSUBS 0.008009f
C787 B.n654 VSUBS 0.008009f
C788 B.n655 VSUBS 0.008009f
C789 B.n656 VSUBS 0.008009f
C790 B.n657 VSUBS 0.008009f
C791 B.n658 VSUBS 0.008009f
C792 B.n659 VSUBS 0.008009f
C793 B.n660 VSUBS 0.008009f
C794 B.n661 VSUBS 0.008009f
C795 B.n662 VSUBS 0.008009f
C796 B.n663 VSUBS 0.008009f
C797 B.n664 VSUBS 0.008009f
C798 B.n665 VSUBS 0.008009f
C799 B.n666 VSUBS 0.008009f
C800 B.n667 VSUBS 0.008009f
C801 B.n668 VSUBS 0.008009f
C802 B.n669 VSUBS 0.008009f
C803 B.n670 VSUBS 0.008009f
C804 B.n671 VSUBS 0.008009f
C805 B.n672 VSUBS 0.008009f
C806 B.n673 VSUBS 0.008009f
C807 B.n674 VSUBS 0.008009f
C808 B.n675 VSUBS 0.008009f
C809 B.n676 VSUBS 0.017882f
C810 B.n677 VSUBS 0.016979f
C811 B.n678 VSUBS 0.016979f
C812 B.n679 VSUBS 0.008009f
C813 B.n680 VSUBS 0.008009f
C814 B.n681 VSUBS 0.008009f
C815 B.n682 VSUBS 0.008009f
C816 B.n683 VSUBS 0.008009f
C817 B.n684 VSUBS 0.008009f
C818 B.n685 VSUBS 0.008009f
C819 B.n686 VSUBS 0.008009f
C820 B.n687 VSUBS 0.008009f
C821 B.n688 VSUBS 0.008009f
C822 B.n689 VSUBS 0.008009f
C823 B.n690 VSUBS 0.008009f
C824 B.n691 VSUBS 0.008009f
C825 B.n692 VSUBS 0.008009f
C826 B.n693 VSUBS 0.008009f
C827 B.n694 VSUBS 0.008009f
C828 B.n695 VSUBS 0.008009f
C829 B.n696 VSUBS 0.008009f
C830 B.n697 VSUBS 0.008009f
C831 B.n698 VSUBS 0.008009f
C832 B.n699 VSUBS 0.008009f
C833 B.n700 VSUBS 0.008009f
C834 B.n701 VSUBS 0.008009f
C835 B.n702 VSUBS 0.008009f
C836 B.n703 VSUBS 0.008009f
C837 B.n704 VSUBS 0.008009f
C838 B.n705 VSUBS 0.008009f
C839 B.n706 VSUBS 0.008009f
C840 B.n707 VSUBS 0.008009f
C841 B.n708 VSUBS 0.008009f
C842 B.n709 VSUBS 0.008009f
C843 B.n710 VSUBS 0.008009f
C844 B.n711 VSUBS 0.008009f
C845 B.n712 VSUBS 0.008009f
C846 B.n713 VSUBS 0.008009f
C847 B.n714 VSUBS 0.008009f
C848 B.n715 VSUBS 0.008009f
C849 B.n716 VSUBS 0.008009f
C850 B.n717 VSUBS 0.008009f
C851 B.n718 VSUBS 0.008009f
C852 B.n719 VSUBS 0.008009f
C853 B.n720 VSUBS 0.008009f
C854 B.n721 VSUBS 0.008009f
C855 B.n722 VSUBS 0.008009f
C856 B.n723 VSUBS 0.008009f
C857 B.n724 VSUBS 0.008009f
C858 B.n725 VSUBS 0.008009f
C859 B.n726 VSUBS 0.008009f
C860 B.n727 VSUBS 0.008009f
C861 B.n728 VSUBS 0.008009f
C862 B.n729 VSUBS 0.008009f
C863 B.n730 VSUBS 0.008009f
C864 B.n731 VSUBS 0.008009f
C865 B.n732 VSUBS 0.008009f
C866 B.n733 VSUBS 0.008009f
C867 B.n734 VSUBS 0.008009f
C868 B.n735 VSUBS 0.008009f
C869 B.n736 VSUBS 0.008009f
C870 B.n737 VSUBS 0.008009f
C871 B.n738 VSUBS 0.008009f
C872 B.n739 VSUBS 0.008009f
C873 B.n740 VSUBS 0.008009f
C874 B.n741 VSUBS 0.008009f
C875 B.n742 VSUBS 0.008009f
C876 B.n743 VSUBS 0.008009f
C877 B.n744 VSUBS 0.008009f
C878 B.n745 VSUBS 0.008009f
C879 B.n746 VSUBS 0.008009f
C880 B.n747 VSUBS 0.008009f
C881 B.n748 VSUBS 0.008009f
C882 B.n749 VSUBS 0.008009f
C883 B.n750 VSUBS 0.008009f
C884 B.n751 VSUBS 0.010451f
C885 B.n752 VSUBS 0.011133f
C886 B.n753 VSUBS 0.022139f
C887 VDD2.t6 VSUBS 0.227311f
C888 VDD2.t0 VSUBS 0.227311f
C889 VDD2.n0 VSUBS 1.75175f
C890 VDD2.t3 VSUBS 0.227311f
C891 VDD2.t7 VSUBS 0.227311f
C892 VDD2.n1 VSUBS 1.75175f
C893 VDD2.n2 VSUBS 3.99228f
C894 VDD2.t4 VSUBS 0.227311f
C895 VDD2.t1 VSUBS 0.227311f
C896 VDD2.n3 VSUBS 1.73957f
C897 VDD2.n4 VSUBS 3.35928f
C898 VDD2.t5 VSUBS 0.227311f
C899 VDD2.t2 VSUBS 0.227311f
C900 VDD2.n5 VSUBS 1.75171f
C901 VTAIL.t13 VSUBS 0.212472f
C902 VTAIL.t15 VSUBS 0.212472f
C903 VTAIL.n0 VSUBS 1.50427f
C904 VTAIL.n1 VSUBS 0.757647f
C905 VTAIL.t9 VSUBS 1.99512f
C906 VTAIL.n2 VSUBS 0.88037f
C907 VTAIL.t1 VSUBS 1.99512f
C908 VTAIL.n3 VSUBS 0.88037f
C909 VTAIL.t0 VSUBS 0.212472f
C910 VTAIL.t2 VSUBS 0.212472f
C911 VTAIL.n4 VSUBS 1.50427f
C912 VTAIL.n5 VSUBS 0.957753f
C913 VTAIL.t7 VSUBS 1.99512f
C914 VTAIL.n6 VSUBS 2.14243f
C915 VTAIL.t11 VSUBS 1.99512f
C916 VTAIL.n7 VSUBS 2.14242f
C917 VTAIL.t14 VSUBS 0.212472f
C918 VTAIL.t8 VSUBS 0.212472f
C919 VTAIL.n8 VSUBS 1.50428f
C920 VTAIL.n9 VSUBS 0.957747f
C921 VTAIL.t10 VSUBS 1.99512f
C922 VTAIL.n10 VSUBS 0.880364f
C923 VTAIL.t3 VSUBS 1.99512f
C924 VTAIL.n11 VSUBS 0.880364f
C925 VTAIL.t4 VSUBS 0.212472f
C926 VTAIL.t6 VSUBS 0.212472f
C927 VTAIL.n12 VSUBS 1.50428f
C928 VTAIL.n13 VSUBS 0.957747f
C929 VTAIL.t5 VSUBS 1.99512f
C930 VTAIL.n14 VSUBS 2.14243f
C931 VTAIL.t12 VSUBS 1.99512f
C932 VTAIL.n15 VSUBS 2.13761f
C933 VN.n0 VSUBS 0.040312f
C934 VN.t0 VSUBS 2.20395f
C935 VN.n1 VSUBS 0.05516f
C936 VN.n2 VSUBS 0.030574f
C937 VN.t4 VSUBS 2.20395f
C938 VN.n3 VSUBS 0.787107f
C939 VN.n4 VSUBS 0.030574f
C940 VN.n5 VSUBS 0.044828f
C941 VN.n6 VSUBS 0.292772f
C942 VN.t7 VSUBS 2.20395f
C943 VN.t1 VSUBS 2.43557f
C944 VN.n7 VSUBS 0.859346f
C945 VN.n8 VSUBS 0.871481f
C946 VN.n9 VSUBS 0.039455f
C947 VN.n10 VSUBS 0.057269f
C948 VN.n11 VSUBS 0.030574f
C949 VN.n12 VSUBS 0.030574f
C950 VN.n13 VSUBS 0.030574f
C951 VN.n14 VSUBS 0.044827f
C952 VN.n15 VSUBS 0.057269f
C953 VN.n16 VSUBS 0.039455f
C954 VN.n17 VSUBS 0.030574f
C955 VN.n18 VSUBS 0.030574f
C956 VN.n19 VSUBS 0.046807f
C957 VN.n20 VSUBS 0.060806f
C958 VN.n21 VSUBS 0.030958f
C959 VN.n22 VSUBS 0.030574f
C960 VN.n23 VSUBS 0.030574f
C961 VN.n24 VSUBS 0.030574f
C962 VN.n25 VSUBS 0.057269f
C963 VN.n26 VSUBS 0.032104f
C964 VN.n27 VSUBS 0.876054f
C965 VN.n28 VSUBS 0.053984f
C966 VN.n29 VSUBS 0.040312f
C967 VN.t3 VSUBS 2.20395f
C968 VN.n30 VSUBS 0.05516f
C969 VN.n31 VSUBS 0.030574f
C970 VN.t6 VSUBS 2.20395f
C971 VN.n32 VSUBS 0.787107f
C972 VN.n33 VSUBS 0.030574f
C973 VN.n34 VSUBS 0.044828f
C974 VN.n35 VSUBS 0.292772f
C975 VN.t2 VSUBS 2.20395f
C976 VN.t5 VSUBS 2.43557f
C977 VN.n36 VSUBS 0.859346f
C978 VN.n37 VSUBS 0.871481f
C979 VN.n38 VSUBS 0.039455f
C980 VN.n39 VSUBS 0.057269f
C981 VN.n40 VSUBS 0.030574f
C982 VN.n41 VSUBS 0.030574f
C983 VN.n42 VSUBS 0.030574f
C984 VN.n43 VSUBS 0.044827f
C985 VN.n44 VSUBS 0.057269f
C986 VN.n45 VSUBS 0.039455f
C987 VN.n46 VSUBS 0.030574f
C988 VN.n47 VSUBS 0.030574f
C989 VN.n48 VSUBS 0.046807f
C990 VN.n49 VSUBS 0.060806f
C991 VN.n50 VSUBS 0.030958f
C992 VN.n51 VSUBS 0.030574f
C993 VN.n52 VSUBS 0.030574f
C994 VN.n53 VSUBS 0.030574f
C995 VN.n54 VSUBS 0.057269f
C996 VN.n55 VSUBS 0.032104f
C997 VN.n56 VSUBS 0.876054f
C998 VN.n57 VSUBS 1.68744f
.ends

