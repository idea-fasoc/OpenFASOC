* NGSPICE file created from diff_pair_sample_1181.ext - technology: sky130A

.subckt diff_pair_sample_1181 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X1 B.t11 B.t9 B.t10 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0 ps=0 w=3.65 l=2.56
X2 VTAIL.t10 VN.t1 VDD2.t6 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X3 VTAIL.t6 VP.t0 VDD1.t7 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0.60225 ps=3.98 w=3.65 l=2.56
X4 VDD2.t5 VN.t2 VTAIL.t9 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=1.4235 ps=8.08 w=3.65 l=2.56
X5 B.t8 B.t6 B.t7 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0 ps=0 w=3.65 l=2.56
X6 VDD1.t6 VP.t1 VTAIL.t3 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X7 VDD2.t4 VN.t3 VTAIL.t15 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X8 VTAIL.t2 VP.t2 VDD1.t5 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X9 VTAIL.t12 VN.t4 VDD2.t3 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0.60225 ps=3.98 w=3.65 l=2.56
X10 B.t5 B.t3 B.t4 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0 ps=0 w=3.65 l=2.56
X11 VDD2.t2 VN.t5 VTAIL.t13 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=1.4235 ps=8.08 w=3.65 l=2.56
X12 VDD1.t4 VP.t3 VTAIL.t1 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=1.4235 ps=8.08 w=3.65 l=2.56
X13 B.t2 B.t0 B.t1 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0 ps=0 w=3.65 l=2.56
X14 VDD1.t3 VP.t4 VTAIL.t7 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X15 VTAIL.t5 VP.t5 VDD1.t2 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X16 VTAIL.t14 VN.t6 VDD2.t1 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0.60225 ps=3.98 w=3.65 l=2.56
X17 VDD1.t1 VP.t6 VTAIL.t4 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=1.4235 ps=8.08 w=3.65 l=2.56
X18 VTAIL.t11 VN.t7 VDD2.t0 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=0.60225 pd=3.98 as=0.60225 ps=3.98 w=3.65 l=2.56
X19 VTAIL.t0 VP.t7 VDD1.t0 w_n3860_n1698# sky130_fd_pr__pfet_01v8 ad=1.4235 pd=8.08 as=0.60225 ps=3.98 w=3.65 l=2.56
R0 VN.n55 VN.n29 161.3
R1 VN.n54 VN.n53 161.3
R2 VN.n52 VN.n30 161.3
R3 VN.n51 VN.n50 161.3
R4 VN.n49 VN.n31 161.3
R5 VN.n48 VN.n47 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n26 VN.n0 161.3
R13 VN.n25 VN.n24 161.3
R14 VN.n23 VN.n1 161.3
R15 VN.n22 VN.n21 161.3
R16 VN.n20 VN.n2 161.3
R17 VN.n19 VN.n18 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n28 VN.n27 106.597
R25 VN.n57 VN.n56 106.597
R26 VN.n7 VN.t6 66.0837
R27 VN.n36 VN.t5 66.0837
R28 VN.n8 VN.n7 62.8231
R29 VN.n37 VN.n36 62.8231
R30 VN.n14 VN.n5 56.5193
R31 VN.n43 VN.n34 56.5193
R32 VN.n21 VN.n1 54.0911
R33 VN.n50 VN.n30 54.0911
R34 VN VN.n57 44.5815
R35 VN.n8 VN.t3 34.3618
R36 VN.n3 VN.t1 34.3618
R37 VN.n27 VN.t2 34.3618
R38 VN.n37 VN.t7 34.3618
R39 VN.n32 VN.t0 34.3618
R40 VN.n56 VN.t4 34.3618
R41 VN.n21 VN.n20 26.8957
R42 VN.n50 VN.n49 26.8957
R43 VN.n10 VN.n9 24.4675
R44 VN.n10 VN.n5 24.4675
R45 VN.n15 VN.n14 24.4675
R46 VN.n16 VN.n15 24.4675
R47 VN.n20 VN.n19 24.4675
R48 VN.n25 VN.n1 24.4675
R49 VN.n26 VN.n25 24.4675
R50 VN.n39 VN.n34 24.4675
R51 VN.n39 VN.n38 24.4675
R52 VN.n49 VN.n48 24.4675
R53 VN.n45 VN.n44 24.4675
R54 VN.n44 VN.n43 24.4675
R55 VN.n55 VN.n54 24.4675
R56 VN.n54 VN.n30 24.4675
R57 VN.n19 VN.n3 14.9254
R58 VN.n48 VN.n32 14.9254
R59 VN.n9 VN.n8 9.54263
R60 VN.n16 VN.n3 9.54263
R61 VN.n38 VN.n37 9.54263
R62 VN.n45 VN.n32 9.54263
R63 VN.n36 VN.n35 7.21701
R64 VN.n7 VN.n6 7.21701
R65 VN.n27 VN.n26 4.15989
R66 VN.n56 VN.n55 4.15989
R67 VN.n57 VN.n29 0.278367
R68 VN.n28 VN.n0 0.278367
R69 VN.n53 VN.n29 0.189894
R70 VN.n53 VN.n52 0.189894
R71 VN.n52 VN.n51 0.189894
R72 VN.n51 VN.n31 0.189894
R73 VN.n47 VN.n31 0.189894
R74 VN.n47 VN.n46 0.189894
R75 VN.n46 VN.n33 0.189894
R76 VN.n42 VN.n33 0.189894
R77 VN.n42 VN.n41 0.189894
R78 VN.n41 VN.n40 0.189894
R79 VN.n40 VN.n35 0.189894
R80 VN.n11 VN.n6 0.189894
R81 VN.n12 VN.n11 0.189894
R82 VN.n13 VN.n12 0.189894
R83 VN.n13 VN.n4 0.189894
R84 VN.n17 VN.n4 0.189894
R85 VN.n18 VN.n17 0.189894
R86 VN.n18 VN.n2 0.189894
R87 VN.n22 VN.n2 0.189894
R88 VN.n23 VN.n22 0.189894
R89 VN.n24 VN.n23 0.189894
R90 VN.n24 VN.n0 0.189894
R91 VN VN.n28 0.153454
R92 VTAIL.n11 VTAIL.t0 115.431
R93 VTAIL.n10 VTAIL.t13 115.431
R94 VTAIL.n7 VTAIL.t12 115.431
R95 VTAIL.n15 VTAIL.t9 115.431
R96 VTAIL.n2 VTAIL.t14 115.431
R97 VTAIL.n3 VTAIL.t4 115.431
R98 VTAIL.n6 VTAIL.t6 115.431
R99 VTAIL.n14 VTAIL.t1 115.431
R100 VTAIL.n13 VTAIL.n12 106.526
R101 VTAIL.n9 VTAIL.n8 106.526
R102 VTAIL.n1 VTAIL.n0 106.526
R103 VTAIL.n5 VTAIL.n4 106.526
R104 VTAIL.n15 VTAIL.n14 18.0048
R105 VTAIL.n7 VTAIL.n6 18.0048
R106 VTAIL.n0 VTAIL.t15 8.90598
R107 VTAIL.n0 VTAIL.t10 8.90598
R108 VTAIL.n4 VTAIL.t7 8.90598
R109 VTAIL.n4 VTAIL.t2 8.90598
R110 VTAIL.n12 VTAIL.t3 8.90598
R111 VTAIL.n12 VTAIL.t5 8.90598
R112 VTAIL.n8 VTAIL.t8 8.90598
R113 VTAIL.n8 VTAIL.t11 8.90598
R114 VTAIL.n9 VTAIL.n7 2.49188
R115 VTAIL.n10 VTAIL.n9 2.49188
R116 VTAIL.n13 VTAIL.n11 2.49188
R117 VTAIL.n14 VTAIL.n13 2.49188
R118 VTAIL.n6 VTAIL.n5 2.49188
R119 VTAIL.n5 VTAIL.n3 2.49188
R120 VTAIL.n2 VTAIL.n1 2.49188
R121 VTAIL VTAIL.n15 2.43369
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 124.395
R126 VDD2.n2 VDD2.n0 124.395
R127 VDD2 VDD2.n5 124.392
R128 VDD2.n4 VDD2.n3 123.206
R129 VDD2.n4 VDD2.n2 38.0731
R130 VDD2.n5 VDD2.t0 8.90598
R131 VDD2.n5 VDD2.t2 8.90598
R132 VDD2.n3 VDD2.t3 8.90598
R133 VDD2.n3 VDD2.t7 8.90598
R134 VDD2.n1 VDD2.t6 8.90598
R135 VDD2.n1 VDD2.t5 8.90598
R136 VDD2.n0 VDD2.t1 8.90598
R137 VDD2.n0 VDD2.t4 8.90598
R138 VDD2 VDD2.n4 1.30438
R139 B.n296 B.n105 585
R140 B.n295 B.n294 585
R141 B.n293 B.n106 585
R142 B.n292 B.n291 585
R143 B.n290 B.n107 585
R144 B.n289 B.n288 585
R145 B.n287 B.n108 585
R146 B.n286 B.n285 585
R147 B.n284 B.n109 585
R148 B.n283 B.n282 585
R149 B.n281 B.n110 585
R150 B.n280 B.n279 585
R151 B.n278 B.n111 585
R152 B.n277 B.n276 585
R153 B.n275 B.n112 585
R154 B.n274 B.n273 585
R155 B.n272 B.n113 585
R156 B.n271 B.n270 585
R157 B.n266 B.n114 585
R158 B.n265 B.n264 585
R159 B.n263 B.n115 585
R160 B.n262 B.n261 585
R161 B.n260 B.n116 585
R162 B.n259 B.n258 585
R163 B.n257 B.n117 585
R164 B.n256 B.n255 585
R165 B.n254 B.n118 585
R166 B.n252 B.n251 585
R167 B.n250 B.n121 585
R168 B.n249 B.n248 585
R169 B.n247 B.n122 585
R170 B.n246 B.n245 585
R171 B.n244 B.n123 585
R172 B.n243 B.n242 585
R173 B.n241 B.n124 585
R174 B.n240 B.n239 585
R175 B.n238 B.n125 585
R176 B.n237 B.n236 585
R177 B.n235 B.n126 585
R178 B.n234 B.n233 585
R179 B.n232 B.n127 585
R180 B.n231 B.n230 585
R181 B.n229 B.n128 585
R182 B.n228 B.n227 585
R183 B.n298 B.n297 585
R184 B.n299 B.n104 585
R185 B.n301 B.n300 585
R186 B.n302 B.n103 585
R187 B.n304 B.n303 585
R188 B.n305 B.n102 585
R189 B.n307 B.n306 585
R190 B.n308 B.n101 585
R191 B.n310 B.n309 585
R192 B.n311 B.n100 585
R193 B.n313 B.n312 585
R194 B.n314 B.n99 585
R195 B.n316 B.n315 585
R196 B.n317 B.n98 585
R197 B.n319 B.n318 585
R198 B.n320 B.n97 585
R199 B.n322 B.n321 585
R200 B.n323 B.n96 585
R201 B.n325 B.n324 585
R202 B.n326 B.n95 585
R203 B.n328 B.n327 585
R204 B.n329 B.n94 585
R205 B.n331 B.n330 585
R206 B.n332 B.n93 585
R207 B.n334 B.n333 585
R208 B.n335 B.n92 585
R209 B.n337 B.n336 585
R210 B.n338 B.n91 585
R211 B.n340 B.n339 585
R212 B.n341 B.n90 585
R213 B.n343 B.n342 585
R214 B.n344 B.n89 585
R215 B.n346 B.n345 585
R216 B.n347 B.n88 585
R217 B.n349 B.n348 585
R218 B.n350 B.n87 585
R219 B.n352 B.n351 585
R220 B.n353 B.n86 585
R221 B.n355 B.n354 585
R222 B.n356 B.n85 585
R223 B.n358 B.n357 585
R224 B.n359 B.n84 585
R225 B.n361 B.n360 585
R226 B.n362 B.n83 585
R227 B.n364 B.n363 585
R228 B.n365 B.n82 585
R229 B.n367 B.n366 585
R230 B.n368 B.n81 585
R231 B.n370 B.n369 585
R232 B.n371 B.n80 585
R233 B.n373 B.n372 585
R234 B.n374 B.n79 585
R235 B.n376 B.n375 585
R236 B.n377 B.n78 585
R237 B.n379 B.n378 585
R238 B.n380 B.n77 585
R239 B.n382 B.n381 585
R240 B.n383 B.n76 585
R241 B.n385 B.n384 585
R242 B.n386 B.n75 585
R243 B.n388 B.n387 585
R244 B.n389 B.n74 585
R245 B.n391 B.n390 585
R246 B.n392 B.n73 585
R247 B.n394 B.n393 585
R248 B.n395 B.n72 585
R249 B.n397 B.n396 585
R250 B.n398 B.n71 585
R251 B.n400 B.n399 585
R252 B.n401 B.n70 585
R253 B.n403 B.n402 585
R254 B.n404 B.n69 585
R255 B.n406 B.n405 585
R256 B.n407 B.n68 585
R257 B.n409 B.n408 585
R258 B.n410 B.n67 585
R259 B.n412 B.n411 585
R260 B.n413 B.n66 585
R261 B.n415 B.n414 585
R262 B.n416 B.n65 585
R263 B.n418 B.n417 585
R264 B.n419 B.n64 585
R265 B.n421 B.n420 585
R266 B.n422 B.n63 585
R267 B.n424 B.n423 585
R268 B.n425 B.n62 585
R269 B.n427 B.n426 585
R270 B.n428 B.n61 585
R271 B.n430 B.n429 585
R272 B.n431 B.n60 585
R273 B.n433 B.n432 585
R274 B.n434 B.n59 585
R275 B.n436 B.n435 585
R276 B.n437 B.n58 585
R277 B.n439 B.n438 585
R278 B.n440 B.n57 585
R279 B.n442 B.n441 585
R280 B.n443 B.n56 585
R281 B.n445 B.n444 585
R282 B.n446 B.n55 585
R283 B.n448 B.n447 585
R284 B.n449 B.n54 585
R285 B.n516 B.n27 585
R286 B.n515 B.n514 585
R287 B.n513 B.n28 585
R288 B.n512 B.n511 585
R289 B.n510 B.n29 585
R290 B.n509 B.n508 585
R291 B.n507 B.n30 585
R292 B.n506 B.n505 585
R293 B.n504 B.n31 585
R294 B.n503 B.n502 585
R295 B.n501 B.n32 585
R296 B.n500 B.n499 585
R297 B.n498 B.n33 585
R298 B.n497 B.n496 585
R299 B.n495 B.n34 585
R300 B.n494 B.n493 585
R301 B.n492 B.n35 585
R302 B.n490 B.n489 585
R303 B.n488 B.n38 585
R304 B.n487 B.n486 585
R305 B.n485 B.n39 585
R306 B.n484 B.n483 585
R307 B.n482 B.n40 585
R308 B.n481 B.n480 585
R309 B.n479 B.n41 585
R310 B.n478 B.n477 585
R311 B.n476 B.n42 585
R312 B.n475 B.n474 585
R313 B.n473 B.n43 585
R314 B.n472 B.n471 585
R315 B.n470 B.n47 585
R316 B.n469 B.n468 585
R317 B.n467 B.n48 585
R318 B.n466 B.n465 585
R319 B.n464 B.n49 585
R320 B.n463 B.n462 585
R321 B.n461 B.n50 585
R322 B.n460 B.n459 585
R323 B.n458 B.n51 585
R324 B.n457 B.n456 585
R325 B.n455 B.n52 585
R326 B.n454 B.n453 585
R327 B.n452 B.n53 585
R328 B.n451 B.n450 585
R329 B.n518 B.n517 585
R330 B.n519 B.n26 585
R331 B.n521 B.n520 585
R332 B.n522 B.n25 585
R333 B.n524 B.n523 585
R334 B.n525 B.n24 585
R335 B.n527 B.n526 585
R336 B.n528 B.n23 585
R337 B.n530 B.n529 585
R338 B.n531 B.n22 585
R339 B.n533 B.n532 585
R340 B.n534 B.n21 585
R341 B.n536 B.n535 585
R342 B.n537 B.n20 585
R343 B.n539 B.n538 585
R344 B.n540 B.n19 585
R345 B.n542 B.n541 585
R346 B.n543 B.n18 585
R347 B.n545 B.n544 585
R348 B.n546 B.n17 585
R349 B.n548 B.n547 585
R350 B.n549 B.n16 585
R351 B.n551 B.n550 585
R352 B.n552 B.n15 585
R353 B.n554 B.n553 585
R354 B.n555 B.n14 585
R355 B.n557 B.n556 585
R356 B.n558 B.n13 585
R357 B.n560 B.n559 585
R358 B.n561 B.n12 585
R359 B.n563 B.n562 585
R360 B.n564 B.n11 585
R361 B.n566 B.n565 585
R362 B.n567 B.n10 585
R363 B.n569 B.n568 585
R364 B.n570 B.n9 585
R365 B.n572 B.n571 585
R366 B.n573 B.n8 585
R367 B.n575 B.n574 585
R368 B.n576 B.n7 585
R369 B.n578 B.n577 585
R370 B.n579 B.n6 585
R371 B.n581 B.n580 585
R372 B.n582 B.n5 585
R373 B.n584 B.n583 585
R374 B.n585 B.n4 585
R375 B.n587 B.n586 585
R376 B.n588 B.n3 585
R377 B.n590 B.n589 585
R378 B.n591 B.n0 585
R379 B.n2 B.n1 585
R380 B.n154 B.n153 585
R381 B.n156 B.n155 585
R382 B.n157 B.n152 585
R383 B.n159 B.n158 585
R384 B.n160 B.n151 585
R385 B.n162 B.n161 585
R386 B.n163 B.n150 585
R387 B.n165 B.n164 585
R388 B.n166 B.n149 585
R389 B.n168 B.n167 585
R390 B.n169 B.n148 585
R391 B.n171 B.n170 585
R392 B.n172 B.n147 585
R393 B.n174 B.n173 585
R394 B.n175 B.n146 585
R395 B.n177 B.n176 585
R396 B.n178 B.n145 585
R397 B.n180 B.n179 585
R398 B.n181 B.n144 585
R399 B.n183 B.n182 585
R400 B.n184 B.n143 585
R401 B.n186 B.n185 585
R402 B.n187 B.n142 585
R403 B.n189 B.n188 585
R404 B.n190 B.n141 585
R405 B.n192 B.n191 585
R406 B.n193 B.n140 585
R407 B.n195 B.n194 585
R408 B.n196 B.n139 585
R409 B.n198 B.n197 585
R410 B.n199 B.n138 585
R411 B.n201 B.n200 585
R412 B.n202 B.n137 585
R413 B.n204 B.n203 585
R414 B.n205 B.n136 585
R415 B.n207 B.n206 585
R416 B.n208 B.n135 585
R417 B.n210 B.n209 585
R418 B.n211 B.n134 585
R419 B.n213 B.n212 585
R420 B.n214 B.n133 585
R421 B.n216 B.n215 585
R422 B.n217 B.n132 585
R423 B.n219 B.n218 585
R424 B.n220 B.n131 585
R425 B.n222 B.n221 585
R426 B.n223 B.n130 585
R427 B.n225 B.n224 585
R428 B.n226 B.n129 585
R429 B.n227 B.n226 492.5
R430 B.n297 B.n296 492.5
R431 B.n451 B.n54 492.5
R432 B.n518 B.n27 492.5
R433 B.n593 B.n592 256.663
R434 B.n119 B.t6 242.347
R435 B.n267 B.t0 242.347
R436 B.n44 B.t3 242.347
R437 B.n36 B.t9 242.347
R438 B.n592 B.n591 235.042
R439 B.n592 B.n2 235.042
R440 B.n267 B.t1 186.871
R441 B.n44 B.t5 186.871
R442 B.n119 B.t7 186.869
R443 B.n36 B.t11 186.869
R444 B.n227 B.n128 163.367
R445 B.n231 B.n128 163.367
R446 B.n232 B.n231 163.367
R447 B.n233 B.n232 163.367
R448 B.n233 B.n126 163.367
R449 B.n237 B.n126 163.367
R450 B.n238 B.n237 163.367
R451 B.n239 B.n238 163.367
R452 B.n239 B.n124 163.367
R453 B.n243 B.n124 163.367
R454 B.n244 B.n243 163.367
R455 B.n245 B.n244 163.367
R456 B.n245 B.n122 163.367
R457 B.n249 B.n122 163.367
R458 B.n250 B.n249 163.367
R459 B.n251 B.n250 163.367
R460 B.n251 B.n118 163.367
R461 B.n256 B.n118 163.367
R462 B.n257 B.n256 163.367
R463 B.n258 B.n257 163.367
R464 B.n258 B.n116 163.367
R465 B.n262 B.n116 163.367
R466 B.n263 B.n262 163.367
R467 B.n264 B.n263 163.367
R468 B.n264 B.n114 163.367
R469 B.n271 B.n114 163.367
R470 B.n272 B.n271 163.367
R471 B.n273 B.n272 163.367
R472 B.n273 B.n112 163.367
R473 B.n277 B.n112 163.367
R474 B.n278 B.n277 163.367
R475 B.n279 B.n278 163.367
R476 B.n279 B.n110 163.367
R477 B.n283 B.n110 163.367
R478 B.n284 B.n283 163.367
R479 B.n285 B.n284 163.367
R480 B.n285 B.n108 163.367
R481 B.n289 B.n108 163.367
R482 B.n290 B.n289 163.367
R483 B.n291 B.n290 163.367
R484 B.n291 B.n106 163.367
R485 B.n295 B.n106 163.367
R486 B.n296 B.n295 163.367
R487 B.n447 B.n54 163.367
R488 B.n447 B.n446 163.367
R489 B.n446 B.n445 163.367
R490 B.n445 B.n56 163.367
R491 B.n441 B.n56 163.367
R492 B.n441 B.n440 163.367
R493 B.n440 B.n439 163.367
R494 B.n439 B.n58 163.367
R495 B.n435 B.n58 163.367
R496 B.n435 B.n434 163.367
R497 B.n434 B.n433 163.367
R498 B.n433 B.n60 163.367
R499 B.n429 B.n60 163.367
R500 B.n429 B.n428 163.367
R501 B.n428 B.n427 163.367
R502 B.n427 B.n62 163.367
R503 B.n423 B.n62 163.367
R504 B.n423 B.n422 163.367
R505 B.n422 B.n421 163.367
R506 B.n421 B.n64 163.367
R507 B.n417 B.n64 163.367
R508 B.n417 B.n416 163.367
R509 B.n416 B.n415 163.367
R510 B.n415 B.n66 163.367
R511 B.n411 B.n66 163.367
R512 B.n411 B.n410 163.367
R513 B.n410 B.n409 163.367
R514 B.n409 B.n68 163.367
R515 B.n405 B.n68 163.367
R516 B.n405 B.n404 163.367
R517 B.n404 B.n403 163.367
R518 B.n403 B.n70 163.367
R519 B.n399 B.n70 163.367
R520 B.n399 B.n398 163.367
R521 B.n398 B.n397 163.367
R522 B.n397 B.n72 163.367
R523 B.n393 B.n72 163.367
R524 B.n393 B.n392 163.367
R525 B.n392 B.n391 163.367
R526 B.n391 B.n74 163.367
R527 B.n387 B.n74 163.367
R528 B.n387 B.n386 163.367
R529 B.n386 B.n385 163.367
R530 B.n385 B.n76 163.367
R531 B.n381 B.n76 163.367
R532 B.n381 B.n380 163.367
R533 B.n380 B.n379 163.367
R534 B.n379 B.n78 163.367
R535 B.n375 B.n78 163.367
R536 B.n375 B.n374 163.367
R537 B.n374 B.n373 163.367
R538 B.n373 B.n80 163.367
R539 B.n369 B.n80 163.367
R540 B.n369 B.n368 163.367
R541 B.n368 B.n367 163.367
R542 B.n367 B.n82 163.367
R543 B.n363 B.n82 163.367
R544 B.n363 B.n362 163.367
R545 B.n362 B.n361 163.367
R546 B.n361 B.n84 163.367
R547 B.n357 B.n84 163.367
R548 B.n357 B.n356 163.367
R549 B.n356 B.n355 163.367
R550 B.n355 B.n86 163.367
R551 B.n351 B.n86 163.367
R552 B.n351 B.n350 163.367
R553 B.n350 B.n349 163.367
R554 B.n349 B.n88 163.367
R555 B.n345 B.n88 163.367
R556 B.n345 B.n344 163.367
R557 B.n344 B.n343 163.367
R558 B.n343 B.n90 163.367
R559 B.n339 B.n90 163.367
R560 B.n339 B.n338 163.367
R561 B.n338 B.n337 163.367
R562 B.n337 B.n92 163.367
R563 B.n333 B.n92 163.367
R564 B.n333 B.n332 163.367
R565 B.n332 B.n331 163.367
R566 B.n331 B.n94 163.367
R567 B.n327 B.n94 163.367
R568 B.n327 B.n326 163.367
R569 B.n326 B.n325 163.367
R570 B.n325 B.n96 163.367
R571 B.n321 B.n96 163.367
R572 B.n321 B.n320 163.367
R573 B.n320 B.n319 163.367
R574 B.n319 B.n98 163.367
R575 B.n315 B.n98 163.367
R576 B.n315 B.n314 163.367
R577 B.n314 B.n313 163.367
R578 B.n313 B.n100 163.367
R579 B.n309 B.n100 163.367
R580 B.n309 B.n308 163.367
R581 B.n308 B.n307 163.367
R582 B.n307 B.n102 163.367
R583 B.n303 B.n102 163.367
R584 B.n303 B.n302 163.367
R585 B.n302 B.n301 163.367
R586 B.n301 B.n104 163.367
R587 B.n297 B.n104 163.367
R588 B.n514 B.n27 163.367
R589 B.n514 B.n513 163.367
R590 B.n513 B.n512 163.367
R591 B.n512 B.n29 163.367
R592 B.n508 B.n29 163.367
R593 B.n508 B.n507 163.367
R594 B.n507 B.n506 163.367
R595 B.n506 B.n31 163.367
R596 B.n502 B.n31 163.367
R597 B.n502 B.n501 163.367
R598 B.n501 B.n500 163.367
R599 B.n500 B.n33 163.367
R600 B.n496 B.n33 163.367
R601 B.n496 B.n495 163.367
R602 B.n495 B.n494 163.367
R603 B.n494 B.n35 163.367
R604 B.n489 B.n35 163.367
R605 B.n489 B.n488 163.367
R606 B.n488 B.n487 163.367
R607 B.n487 B.n39 163.367
R608 B.n483 B.n39 163.367
R609 B.n483 B.n482 163.367
R610 B.n482 B.n481 163.367
R611 B.n481 B.n41 163.367
R612 B.n477 B.n41 163.367
R613 B.n477 B.n476 163.367
R614 B.n476 B.n475 163.367
R615 B.n475 B.n43 163.367
R616 B.n471 B.n43 163.367
R617 B.n471 B.n470 163.367
R618 B.n470 B.n469 163.367
R619 B.n469 B.n48 163.367
R620 B.n465 B.n48 163.367
R621 B.n465 B.n464 163.367
R622 B.n464 B.n463 163.367
R623 B.n463 B.n50 163.367
R624 B.n459 B.n50 163.367
R625 B.n459 B.n458 163.367
R626 B.n458 B.n457 163.367
R627 B.n457 B.n52 163.367
R628 B.n453 B.n52 163.367
R629 B.n453 B.n452 163.367
R630 B.n452 B.n451 163.367
R631 B.n519 B.n518 163.367
R632 B.n520 B.n519 163.367
R633 B.n520 B.n25 163.367
R634 B.n524 B.n25 163.367
R635 B.n525 B.n524 163.367
R636 B.n526 B.n525 163.367
R637 B.n526 B.n23 163.367
R638 B.n530 B.n23 163.367
R639 B.n531 B.n530 163.367
R640 B.n532 B.n531 163.367
R641 B.n532 B.n21 163.367
R642 B.n536 B.n21 163.367
R643 B.n537 B.n536 163.367
R644 B.n538 B.n537 163.367
R645 B.n538 B.n19 163.367
R646 B.n542 B.n19 163.367
R647 B.n543 B.n542 163.367
R648 B.n544 B.n543 163.367
R649 B.n544 B.n17 163.367
R650 B.n548 B.n17 163.367
R651 B.n549 B.n548 163.367
R652 B.n550 B.n549 163.367
R653 B.n550 B.n15 163.367
R654 B.n554 B.n15 163.367
R655 B.n555 B.n554 163.367
R656 B.n556 B.n555 163.367
R657 B.n556 B.n13 163.367
R658 B.n560 B.n13 163.367
R659 B.n561 B.n560 163.367
R660 B.n562 B.n561 163.367
R661 B.n562 B.n11 163.367
R662 B.n566 B.n11 163.367
R663 B.n567 B.n566 163.367
R664 B.n568 B.n567 163.367
R665 B.n568 B.n9 163.367
R666 B.n572 B.n9 163.367
R667 B.n573 B.n572 163.367
R668 B.n574 B.n573 163.367
R669 B.n574 B.n7 163.367
R670 B.n578 B.n7 163.367
R671 B.n579 B.n578 163.367
R672 B.n580 B.n579 163.367
R673 B.n580 B.n5 163.367
R674 B.n584 B.n5 163.367
R675 B.n585 B.n584 163.367
R676 B.n586 B.n585 163.367
R677 B.n586 B.n3 163.367
R678 B.n590 B.n3 163.367
R679 B.n591 B.n590 163.367
R680 B.n154 B.n2 163.367
R681 B.n155 B.n154 163.367
R682 B.n155 B.n152 163.367
R683 B.n159 B.n152 163.367
R684 B.n160 B.n159 163.367
R685 B.n161 B.n160 163.367
R686 B.n161 B.n150 163.367
R687 B.n165 B.n150 163.367
R688 B.n166 B.n165 163.367
R689 B.n167 B.n166 163.367
R690 B.n167 B.n148 163.367
R691 B.n171 B.n148 163.367
R692 B.n172 B.n171 163.367
R693 B.n173 B.n172 163.367
R694 B.n173 B.n146 163.367
R695 B.n177 B.n146 163.367
R696 B.n178 B.n177 163.367
R697 B.n179 B.n178 163.367
R698 B.n179 B.n144 163.367
R699 B.n183 B.n144 163.367
R700 B.n184 B.n183 163.367
R701 B.n185 B.n184 163.367
R702 B.n185 B.n142 163.367
R703 B.n189 B.n142 163.367
R704 B.n190 B.n189 163.367
R705 B.n191 B.n190 163.367
R706 B.n191 B.n140 163.367
R707 B.n195 B.n140 163.367
R708 B.n196 B.n195 163.367
R709 B.n197 B.n196 163.367
R710 B.n197 B.n138 163.367
R711 B.n201 B.n138 163.367
R712 B.n202 B.n201 163.367
R713 B.n203 B.n202 163.367
R714 B.n203 B.n136 163.367
R715 B.n207 B.n136 163.367
R716 B.n208 B.n207 163.367
R717 B.n209 B.n208 163.367
R718 B.n209 B.n134 163.367
R719 B.n213 B.n134 163.367
R720 B.n214 B.n213 163.367
R721 B.n215 B.n214 163.367
R722 B.n215 B.n132 163.367
R723 B.n219 B.n132 163.367
R724 B.n220 B.n219 163.367
R725 B.n221 B.n220 163.367
R726 B.n221 B.n130 163.367
R727 B.n225 B.n130 163.367
R728 B.n226 B.n225 163.367
R729 B.n268 B.t2 130.822
R730 B.n45 B.t4 130.822
R731 B.n120 B.t8 130.82
R732 B.n37 B.t10 130.82
R733 B.n253 B.n120 59.5399
R734 B.n269 B.n268 59.5399
R735 B.n46 B.n45 59.5399
R736 B.n491 B.n37 59.5399
R737 B.n120 B.n119 56.049
R738 B.n268 B.n267 56.049
R739 B.n45 B.n44 56.049
R740 B.n37 B.n36 56.049
R741 B.n517 B.n516 32.0005
R742 B.n450 B.n449 32.0005
R743 B.n298 B.n105 32.0005
R744 B.n228 B.n129 32.0005
R745 B B.n593 18.0485
R746 B.n517 B.n26 10.6151
R747 B.n521 B.n26 10.6151
R748 B.n522 B.n521 10.6151
R749 B.n523 B.n522 10.6151
R750 B.n523 B.n24 10.6151
R751 B.n527 B.n24 10.6151
R752 B.n528 B.n527 10.6151
R753 B.n529 B.n528 10.6151
R754 B.n529 B.n22 10.6151
R755 B.n533 B.n22 10.6151
R756 B.n534 B.n533 10.6151
R757 B.n535 B.n534 10.6151
R758 B.n535 B.n20 10.6151
R759 B.n539 B.n20 10.6151
R760 B.n540 B.n539 10.6151
R761 B.n541 B.n540 10.6151
R762 B.n541 B.n18 10.6151
R763 B.n545 B.n18 10.6151
R764 B.n546 B.n545 10.6151
R765 B.n547 B.n546 10.6151
R766 B.n547 B.n16 10.6151
R767 B.n551 B.n16 10.6151
R768 B.n552 B.n551 10.6151
R769 B.n553 B.n552 10.6151
R770 B.n553 B.n14 10.6151
R771 B.n557 B.n14 10.6151
R772 B.n558 B.n557 10.6151
R773 B.n559 B.n558 10.6151
R774 B.n559 B.n12 10.6151
R775 B.n563 B.n12 10.6151
R776 B.n564 B.n563 10.6151
R777 B.n565 B.n564 10.6151
R778 B.n565 B.n10 10.6151
R779 B.n569 B.n10 10.6151
R780 B.n570 B.n569 10.6151
R781 B.n571 B.n570 10.6151
R782 B.n571 B.n8 10.6151
R783 B.n575 B.n8 10.6151
R784 B.n576 B.n575 10.6151
R785 B.n577 B.n576 10.6151
R786 B.n577 B.n6 10.6151
R787 B.n581 B.n6 10.6151
R788 B.n582 B.n581 10.6151
R789 B.n583 B.n582 10.6151
R790 B.n583 B.n4 10.6151
R791 B.n587 B.n4 10.6151
R792 B.n588 B.n587 10.6151
R793 B.n589 B.n588 10.6151
R794 B.n589 B.n0 10.6151
R795 B.n516 B.n515 10.6151
R796 B.n515 B.n28 10.6151
R797 B.n511 B.n28 10.6151
R798 B.n511 B.n510 10.6151
R799 B.n510 B.n509 10.6151
R800 B.n509 B.n30 10.6151
R801 B.n505 B.n30 10.6151
R802 B.n505 B.n504 10.6151
R803 B.n504 B.n503 10.6151
R804 B.n503 B.n32 10.6151
R805 B.n499 B.n32 10.6151
R806 B.n499 B.n498 10.6151
R807 B.n498 B.n497 10.6151
R808 B.n497 B.n34 10.6151
R809 B.n493 B.n34 10.6151
R810 B.n493 B.n492 10.6151
R811 B.n490 B.n38 10.6151
R812 B.n486 B.n38 10.6151
R813 B.n486 B.n485 10.6151
R814 B.n485 B.n484 10.6151
R815 B.n484 B.n40 10.6151
R816 B.n480 B.n40 10.6151
R817 B.n480 B.n479 10.6151
R818 B.n479 B.n478 10.6151
R819 B.n478 B.n42 10.6151
R820 B.n474 B.n473 10.6151
R821 B.n473 B.n472 10.6151
R822 B.n472 B.n47 10.6151
R823 B.n468 B.n47 10.6151
R824 B.n468 B.n467 10.6151
R825 B.n467 B.n466 10.6151
R826 B.n466 B.n49 10.6151
R827 B.n462 B.n49 10.6151
R828 B.n462 B.n461 10.6151
R829 B.n461 B.n460 10.6151
R830 B.n460 B.n51 10.6151
R831 B.n456 B.n51 10.6151
R832 B.n456 B.n455 10.6151
R833 B.n455 B.n454 10.6151
R834 B.n454 B.n53 10.6151
R835 B.n450 B.n53 10.6151
R836 B.n449 B.n448 10.6151
R837 B.n448 B.n55 10.6151
R838 B.n444 B.n55 10.6151
R839 B.n444 B.n443 10.6151
R840 B.n443 B.n442 10.6151
R841 B.n442 B.n57 10.6151
R842 B.n438 B.n57 10.6151
R843 B.n438 B.n437 10.6151
R844 B.n437 B.n436 10.6151
R845 B.n436 B.n59 10.6151
R846 B.n432 B.n59 10.6151
R847 B.n432 B.n431 10.6151
R848 B.n431 B.n430 10.6151
R849 B.n430 B.n61 10.6151
R850 B.n426 B.n61 10.6151
R851 B.n426 B.n425 10.6151
R852 B.n425 B.n424 10.6151
R853 B.n424 B.n63 10.6151
R854 B.n420 B.n63 10.6151
R855 B.n420 B.n419 10.6151
R856 B.n419 B.n418 10.6151
R857 B.n418 B.n65 10.6151
R858 B.n414 B.n65 10.6151
R859 B.n414 B.n413 10.6151
R860 B.n413 B.n412 10.6151
R861 B.n412 B.n67 10.6151
R862 B.n408 B.n67 10.6151
R863 B.n408 B.n407 10.6151
R864 B.n407 B.n406 10.6151
R865 B.n406 B.n69 10.6151
R866 B.n402 B.n69 10.6151
R867 B.n402 B.n401 10.6151
R868 B.n401 B.n400 10.6151
R869 B.n400 B.n71 10.6151
R870 B.n396 B.n71 10.6151
R871 B.n396 B.n395 10.6151
R872 B.n395 B.n394 10.6151
R873 B.n394 B.n73 10.6151
R874 B.n390 B.n73 10.6151
R875 B.n390 B.n389 10.6151
R876 B.n389 B.n388 10.6151
R877 B.n388 B.n75 10.6151
R878 B.n384 B.n75 10.6151
R879 B.n384 B.n383 10.6151
R880 B.n383 B.n382 10.6151
R881 B.n382 B.n77 10.6151
R882 B.n378 B.n77 10.6151
R883 B.n378 B.n377 10.6151
R884 B.n377 B.n376 10.6151
R885 B.n376 B.n79 10.6151
R886 B.n372 B.n79 10.6151
R887 B.n372 B.n371 10.6151
R888 B.n371 B.n370 10.6151
R889 B.n370 B.n81 10.6151
R890 B.n366 B.n81 10.6151
R891 B.n366 B.n365 10.6151
R892 B.n365 B.n364 10.6151
R893 B.n364 B.n83 10.6151
R894 B.n360 B.n83 10.6151
R895 B.n360 B.n359 10.6151
R896 B.n359 B.n358 10.6151
R897 B.n358 B.n85 10.6151
R898 B.n354 B.n85 10.6151
R899 B.n354 B.n353 10.6151
R900 B.n353 B.n352 10.6151
R901 B.n352 B.n87 10.6151
R902 B.n348 B.n87 10.6151
R903 B.n348 B.n347 10.6151
R904 B.n347 B.n346 10.6151
R905 B.n346 B.n89 10.6151
R906 B.n342 B.n89 10.6151
R907 B.n342 B.n341 10.6151
R908 B.n341 B.n340 10.6151
R909 B.n340 B.n91 10.6151
R910 B.n336 B.n91 10.6151
R911 B.n336 B.n335 10.6151
R912 B.n335 B.n334 10.6151
R913 B.n334 B.n93 10.6151
R914 B.n330 B.n93 10.6151
R915 B.n330 B.n329 10.6151
R916 B.n329 B.n328 10.6151
R917 B.n328 B.n95 10.6151
R918 B.n324 B.n95 10.6151
R919 B.n324 B.n323 10.6151
R920 B.n323 B.n322 10.6151
R921 B.n322 B.n97 10.6151
R922 B.n318 B.n97 10.6151
R923 B.n318 B.n317 10.6151
R924 B.n317 B.n316 10.6151
R925 B.n316 B.n99 10.6151
R926 B.n312 B.n99 10.6151
R927 B.n312 B.n311 10.6151
R928 B.n311 B.n310 10.6151
R929 B.n310 B.n101 10.6151
R930 B.n306 B.n101 10.6151
R931 B.n306 B.n305 10.6151
R932 B.n305 B.n304 10.6151
R933 B.n304 B.n103 10.6151
R934 B.n300 B.n103 10.6151
R935 B.n300 B.n299 10.6151
R936 B.n299 B.n298 10.6151
R937 B.n153 B.n1 10.6151
R938 B.n156 B.n153 10.6151
R939 B.n157 B.n156 10.6151
R940 B.n158 B.n157 10.6151
R941 B.n158 B.n151 10.6151
R942 B.n162 B.n151 10.6151
R943 B.n163 B.n162 10.6151
R944 B.n164 B.n163 10.6151
R945 B.n164 B.n149 10.6151
R946 B.n168 B.n149 10.6151
R947 B.n169 B.n168 10.6151
R948 B.n170 B.n169 10.6151
R949 B.n170 B.n147 10.6151
R950 B.n174 B.n147 10.6151
R951 B.n175 B.n174 10.6151
R952 B.n176 B.n175 10.6151
R953 B.n176 B.n145 10.6151
R954 B.n180 B.n145 10.6151
R955 B.n181 B.n180 10.6151
R956 B.n182 B.n181 10.6151
R957 B.n182 B.n143 10.6151
R958 B.n186 B.n143 10.6151
R959 B.n187 B.n186 10.6151
R960 B.n188 B.n187 10.6151
R961 B.n188 B.n141 10.6151
R962 B.n192 B.n141 10.6151
R963 B.n193 B.n192 10.6151
R964 B.n194 B.n193 10.6151
R965 B.n194 B.n139 10.6151
R966 B.n198 B.n139 10.6151
R967 B.n199 B.n198 10.6151
R968 B.n200 B.n199 10.6151
R969 B.n200 B.n137 10.6151
R970 B.n204 B.n137 10.6151
R971 B.n205 B.n204 10.6151
R972 B.n206 B.n205 10.6151
R973 B.n206 B.n135 10.6151
R974 B.n210 B.n135 10.6151
R975 B.n211 B.n210 10.6151
R976 B.n212 B.n211 10.6151
R977 B.n212 B.n133 10.6151
R978 B.n216 B.n133 10.6151
R979 B.n217 B.n216 10.6151
R980 B.n218 B.n217 10.6151
R981 B.n218 B.n131 10.6151
R982 B.n222 B.n131 10.6151
R983 B.n223 B.n222 10.6151
R984 B.n224 B.n223 10.6151
R985 B.n224 B.n129 10.6151
R986 B.n229 B.n228 10.6151
R987 B.n230 B.n229 10.6151
R988 B.n230 B.n127 10.6151
R989 B.n234 B.n127 10.6151
R990 B.n235 B.n234 10.6151
R991 B.n236 B.n235 10.6151
R992 B.n236 B.n125 10.6151
R993 B.n240 B.n125 10.6151
R994 B.n241 B.n240 10.6151
R995 B.n242 B.n241 10.6151
R996 B.n242 B.n123 10.6151
R997 B.n246 B.n123 10.6151
R998 B.n247 B.n246 10.6151
R999 B.n248 B.n247 10.6151
R1000 B.n248 B.n121 10.6151
R1001 B.n252 B.n121 10.6151
R1002 B.n255 B.n254 10.6151
R1003 B.n255 B.n117 10.6151
R1004 B.n259 B.n117 10.6151
R1005 B.n260 B.n259 10.6151
R1006 B.n261 B.n260 10.6151
R1007 B.n261 B.n115 10.6151
R1008 B.n265 B.n115 10.6151
R1009 B.n266 B.n265 10.6151
R1010 B.n270 B.n266 10.6151
R1011 B.n274 B.n113 10.6151
R1012 B.n275 B.n274 10.6151
R1013 B.n276 B.n275 10.6151
R1014 B.n276 B.n111 10.6151
R1015 B.n280 B.n111 10.6151
R1016 B.n281 B.n280 10.6151
R1017 B.n282 B.n281 10.6151
R1018 B.n282 B.n109 10.6151
R1019 B.n286 B.n109 10.6151
R1020 B.n287 B.n286 10.6151
R1021 B.n288 B.n287 10.6151
R1022 B.n288 B.n107 10.6151
R1023 B.n292 B.n107 10.6151
R1024 B.n293 B.n292 10.6151
R1025 B.n294 B.n293 10.6151
R1026 B.n294 B.n105 10.6151
R1027 B.n492 B.n491 9.36635
R1028 B.n474 B.n46 9.36635
R1029 B.n253 B.n252 9.36635
R1030 B.n269 B.n113 9.36635
R1031 B.n593 B.n0 8.11757
R1032 B.n593 B.n1 8.11757
R1033 B.n491 B.n490 1.24928
R1034 B.n46 B.n42 1.24928
R1035 B.n254 B.n253 1.24928
R1036 B.n270 B.n269 1.24928
R1037 VP.n19 VP.n16 161.3
R1038 VP.n21 VP.n20 161.3
R1039 VP.n22 VP.n15 161.3
R1040 VP.n24 VP.n23 161.3
R1041 VP.n25 VP.n14 161.3
R1042 VP.n27 VP.n26 161.3
R1043 VP.n29 VP.n28 161.3
R1044 VP.n30 VP.n12 161.3
R1045 VP.n32 VP.n31 161.3
R1046 VP.n33 VP.n11 161.3
R1047 VP.n35 VP.n34 161.3
R1048 VP.n36 VP.n10 161.3
R1049 VP.n68 VP.n0 161.3
R1050 VP.n67 VP.n66 161.3
R1051 VP.n65 VP.n1 161.3
R1052 VP.n64 VP.n63 161.3
R1053 VP.n62 VP.n2 161.3
R1054 VP.n61 VP.n60 161.3
R1055 VP.n59 VP.n58 161.3
R1056 VP.n57 VP.n4 161.3
R1057 VP.n56 VP.n55 161.3
R1058 VP.n54 VP.n5 161.3
R1059 VP.n53 VP.n52 161.3
R1060 VP.n51 VP.n6 161.3
R1061 VP.n49 VP.n48 161.3
R1062 VP.n47 VP.n7 161.3
R1063 VP.n46 VP.n45 161.3
R1064 VP.n44 VP.n8 161.3
R1065 VP.n43 VP.n42 161.3
R1066 VP.n41 VP.n9 161.3
R1067 VP.n40 VP.n39 106.597
R1068 VP.n70 VP.n69 106.597
R1069 VP.n38 VP.n37 106.597
R1070 VP.n17 VP.t7 66.0837
R1071 VP.n18 VP.n17 62.8231
R1072 VP.n56 VP.n5 56.5193
R1073 VP.n24 VP.n15 56.5193
R1074 VP.n45 VP.n44 54.0911
R1075 VP.n63 VP.n1 54.0911
R1076 VP.n31 VP.n11 54.0911
R1077 VP.n40 VP.n38 44.3026
R1078 VP.n39 VP.t0 34.3618
R1079 VP.n50 VP.t4 34.3618
R1080 VP.n3 VP.t2 34.3618
R1081 VP.n69 VP.t6 34.3618
R1082 VP.n37 VP.t3 34.3618
R1083 VP.n13 VP.t5 34.3618
R1084 VP.n18 VP.t1 34.3618
R1085 VP.n45 VP.n7 26.8957
R1086 VP.n63 VP.n62 26.8957
R1087 VP.n31 VP.n30 26.8957
R1088 VP.n43 VP.n9 24.4675
R1089 VP.n44 VP.n43 24.4675
R1090 VP.n49 VP.n7 24.4675
R1091 VP.n52 VP.n51 24.4675
R1092 VP.n52 VP.n5 24.4675
R1093 VP.n57 VP.n56 24.4675
R1094 VP.n58 VP.n57 24.4675
R1095 VP.n62 VP.n61 24.4675
R1096 VP.n67 VP.n1 24.4675
R1097 VP.n68 VP.n67 24.4675
R1098 VP.n35 VP.n11 24.4675
R1099 VP.n36 VP.n35 24.4675
R1100 VP.n25 VP.n24 24.4675
R1101 VP.n26 VP.n25 24.4675
R1102 VP.n30 VP.n29 24.4675
R1103 VP.n20 VP.n19 24.4675
R1104 VP.n20 VP.n15 24.4675
R1105 VP.n50 VP.n49 14.9254
R1106 VP.n61 VP.n3 14.9254
R1107 VP.n29 VP.n13 14.9254
R1108 VP.n51 VP.n50 9.54263
R1109 VP.n58 VP.n3 9.54263
R1110 VP.n26 VP.n13 9.54263
R1111 VP.n19 VP.n18 9.54263
R1112 VP.n17 VP.n16 7.21701
R1113 VP.n39 VP.n9 4.15989
R1114 VP.n69 VP.n68 4.15989
R1115 VP.n37 VP.n36 4.15989
R1116 VP.n38 VP.n10 0.278367
R1117 VP.n41 VP.n40 0.278367
R1118 VP.n70 VP.n0 0.278367
R1119 VP.n21 VP.n16 0.189894
R1120 VP.n22 VP.n21 0.189894
R1121 VP.n23 VP.n22 0.189894
R1122 VP.n23 VP.n14 0.189894
R1123 VP.n27 VP.n14 0.189894
R1124 VP.n28 VP.n27 0.189894
R1125 VP.n28 VP.n12 0.189894
R1126 VP.n32 VP.n12 0.189894
R1127 VP.n33 VP.n32 0.189894
R1128 VP.n34 VP.n33 0.189894
R1129 VP.n34 VP.n10 0.189894
R1130 VP.n42 VP.n41 0.189894
R1131 VP.n42 VP.n8 0.189894
R1132 VP.n46 VP.n8 0.189894
R1133 VP.n47 VP.n46 0.189894
R1134 VP.n48 VP.n47 0.189894
R1135 VP.n48 VP.n6 0.189894
R1136 VP.n53 VP.n6 0.189894
R1137 VP.n54 VP.n53 0.189894
R1138 VP.n55 VP.n54 0.189894
R1139 VP.n55 VP.n4 0.189894
R1140 VP.n59 VP.n4 0.189894
R1141 VP.n60 VP.n59 0.189894
R1142 VP.n60 VP.n2 0.189894
R1143 VP.n64 VP.n2 0.189894
R1144 VP.n65 VP.n64 0.189894
R1145 VP.n66 VP.n65 0.189894
R1146 VP.n66 VP.n0 0.189894
R1147 VP VP.n70 0.153454
R1148 VDD1 VDD1.n0 124.51
R1149 VDD1.n3 VDD1.n2 124.395
R1150 VDD1.n3 VDD1.n1 124.395
R1151 VDD1.n5 VDD1.n4 123.206
R1152 VDD1.n5 VDD1.n3 38.6561
R1153 VDD1.n4 VDD1.t2 8.90598
R1154 VDD1.n4 VDD1.t4 8.90598
R1155 VDD1.n0 VDD1.t0 8.90598
R1156 VDD1.n0 VDD1.t6 8.90598
R1157 VDD1.n2 VDD1.t5 8.90598
R1158 VDD1.n2 VDD1.t1 8.90598
R1159 VDD1.n1 VDD1.t7 8.90598
R1160 VDD1.n1 VDD1.t3 8.90598
R1161 VDD1 VDD1.n5 1.188
C0 B VP 1.98021f
C1 VDD1 B 1.41065f
C2 VDD1 VP 3.31182f
C3 w_n3860_n1698# VN 7.704f
C4 VTAIL VN 3.91302f
C5 VTAIL w_n3860_n1698# 2.3105f
C6 VN VDD2 2.94959f
C7 w_n3860_n1698# VDD2 1.82931f
C8 VTAIL VDD2 5.29226f
C9 B VN 1.14086f
C10 VP VN 6.0767f
C11 B w_n3860_n1698# 7.73635f
C12 VP w_n3860_n1698# 8.203639f
C13 VDD1 VN 0.156172f
C14 VTAIL B 2.18719f
C15 VTAIL VP 3.92713f
C16 VDD1 w_n3860_n1698# 1.71669f
C17 VDD1 VTAIL 5.23812f
C18 B VDD2 1.50559f
C19 VP VDD2 0.520593f
C20 VDD1 VDD2 1.75652f
C21 VDD2 VSUBS 1.446048f
C22 VDD1 VSUBS 2.099092f
C23 VTAIL VSUBS 0.625343f
C24 VN VSUBS 6.46845f
C25 VP VSUBS 2.971938f
C26 B VSUBS 4.004032f
C27 w_n3860_n1698# VSUBS 82.681206f
C28 VDD1.t0 VSUBS 0.071202f
C29 VDD1.t6 VSUBS 0.071202f
C30 VDD1.n0 VSUBS 0.409463f
C31 VDD1.t7 VSUBS 0.071202f
C32 VDD1.t3 VSUBS 0.071202f
C33 VDD1.n1 VSUBS 0.408793f
C34 VDD1.t5 VSUBS 0.071202f
C35 VDD1.t1 VSUBS 0.071202f
C36 VDD1.n2 VSUBS 0.408793f
C37 VDD1.n3 VSUBS 3.03655f
C38 VDD1.t2 VSUBS 0.071202f
C39 VDD1.t4 VSUBS 0.071202f
C40 VDD1.n4 VSUBS 0.40266f
C41 VDD1.n5 VSUBS 2.42327f
C42 VP.n0 VSUBS 0.06011f
C43 VP.t6 VSUBS 1.08488f
C44 VP.n1 VSUBS 0.079915f
C45 VP.n2 VSUBS 0.045593f
C46 VP.t2 VSUBS 1.08488f
C47 VP.n3 VSUBS 0.439917f
C48 VP.n4 VSUBS 0.045593f
C49 VP.n5 VSUBS 0.066557f
C50 VP.n6 VSUBS 0.045593f
C51 VP.t4 VSUBS 1.08488f
C52 VP.n7 VSUBS 0.08838f
C53 VP.n8 VSUBS 0.045593f
C54 VP.n9 VSUBS 0.050152f
C55 VP.n10 VSUBS 0.06011f
C56 VP.t3 VSUBS 1.08488f
C57 VP.n11 VSUBS 0.079915f
C58 VP.n12 VSUBS 0.045593f
C59 VP.t5 VSUBS 1.08488f
C60 VP.n13 VSUBS 0.439917f
C61 VP.n14 VSUBS 0.045593f
C62 VP.n15 VSUBS 0.066557f
C63 VP.n16 VSUBS 0.437945f
C64 VP.t1 VSUBS 1.08488f
C65 VP.t7 VSUBS 1.42812f
C66 VP.n17 VSUBS 0.553376f
C67 VP.n18 VSUBS 0.566011f
C68 VP.n19 VSUBS 0.059381f
C69 VP.n20 VSUBS 0.084974f
C70 VP.n21 VSUBS 0.045593f
C71 VP.n22 VSUBS 0.045593f
C72 VP.n23 VSUBS 0.045593f
C73 VP.n24 VSUBS 0.066557f
C74 VP.n25 VSUBS 0.084974f
C75 VP.n26 VSUBS 0.059381f
C76 VP.n27 VSUBS 0.045593f
C77 VP.n28 VSUBS 0.045593f
C78 VP.n29 VSUBS 0.06861f
C79 VP.n30 VSUBS 0.08838f
C80 VP.n31 VSUBS 0.049793f
C81 VP.n32 VSUBS 0.045593f
C82 VP.n33 VSUBS 0.045593f
C83 VP.n34 VSUBS 0.045593f
C84 VP.n35 VSUBS 0.084974f
C85 VP.n36 VSUBS 0.050152f
C86 VP.n37 VSUBS 0.576218f
C87 VP.n38 VSUBS 2.1156f
C88 VP.t0 VSUBS 1.08488f
C89 VP.n39 VSUBS 0.576218f
C90 VP.n40 VSUBS 2.1526f
C91 VP.n41 VSUBS 0.06011f
C92 VP.n42 VSUBS 0.045593f
C93 VP.n43 VSUBS 0.084974f
C94 VP.n44 VSUBS 0.079915f
C95 VP.n45 VSUBS 0.049793f
C96 VP.n46 VSUBS 0.045593f
C97 VP.n47 VSUBS 0.045593f
C98 VP.n48 VSUBS 0.045593f
C99 VP.n49 VSUBS 0.06861f
C100 VP.n50 VSUBS 0.439917f
C101 VP.n51 VSUBS 0.059381f
C102 VP.n52 VSUBS 0.084974f
C103 VP.n53 VSUBS 0.045593f
C104 VP.n54 VSUBS 0.045593f
C105 VP.n55 VSUBS 0.045593f
C106 VP.n56 VSUBS 0.066557f
C107 VP.n57 VSUBS 0.084974f
C108 VP.n58 VSUBS 0.059381f
C109 VP.n59 VSUBS 0.045593f
C110 VP.n60 VSUBS 0.045593f
C111 VP.n61 VSUBS 0.06861f
C112 VP.n62 VSUBS 0.08838f
C113 VP.n63 VSUBS 0.049793f
C114 VP.n64 VSUBS 0.045593f
C115 VP.n65 VSUBS 0.045593f
C116 VP.n66 VSUBS 0.045593f
C117 VP.n67 VSUBS 0.084974f
C118 VP.n68 VSUBS 0.050152f
C119 VP.n69 VSUBS 0.576218f
C120 VP.n70 VSUBS 0.079558f
C121 B.n0 VSUBS 0.008111f
C122 B.n1 VSUBS 0.008111f
C123 B.n2 VSUBS 0.011995f
C124 B.n3 VSUBS 0.009192f
C125 B.n4 VSUBS 0.009192f
C126 B.n5 VSUBS 0.009192f
C127 B.n6 VSUBS 0.009192f
C128 B.n7 VSUBS 0.009192f
C129 B.n8 VSUBS 0.009192f
C130 B.n9 VSUBS 0.009192f
C131 B.n10 VSUBS 0.009192f
C132 B.n11 VSUBS 0.009192f
C133 B.n12 VSUBS 0.009192f
C134 B.n13 VSUBS 0.009192f
C135 B.n14 VSUBS 0.009192f
C136 B.n15 VSUBS 0.009192f
C137 B.n16 VSUBS 0.009192f
C138 B.n17 VSUBS 0.009192f
C139 B.n18 VSUBS 0.009192f
C140 B.n19 VSUBS 0.009192f
C141 B.n20 VSUBS 0.009192f
C142 B.n21 VSUBS 0.009192f
C143 B.n22 VSUBS 0.009192f
C144 B.n23 VSUBS 0.009192f
C145 B.n24 VSUBS 0.009192f
C146 B.n25 VSUBS 0.009192f
C147 B.n26 VSUBS 0.009192f
C148 B.n27 VSUBS 0.021994f
C149 B.n28 VSUBS 0.009192f
C150 B.n29 VSUBS 0.009192f
C151 B.n30 VSUBS 0.009192f
C152 B.n31 VSUBS 0.009192f
C153 B.n32 VSUBS 0.009192f
C154 B.n33 VSUBS 0.009192f
C155 B.n34 VSUBS 0.009192f
C156 B.n35 VSUBS 0.009192f
C157 B.t10 VSUBS 0.122244f
C158 B.t11 VSUBS 0.14498f
C159 B.t9 VSUBS 0.592166f
C160 B.n36 VSUBS 0.115683f
C161 B.n37 VSUBS 0.088914f
C162 B.n38 VSUBS 0.009192f
C163 B.n39 VSUBS 0.009192f
C164 B.n40 VSUBS 0.009192f
C165 B.n41 VSUBS 0.009192f
C166 B.n42 VSUBS 0.005137f
C167 B.n43 VSUBS 0.009192f
C168 B.t4 VSUBS 0.122244f
C169 B.t5 VSUBS 0.14498f
C170 B.t3 VSUBS 0.592166f
C171 B.n44 VSUBS 0.115683f
C172 B.n45 VSUBS 0.088914f
C173 B.n46 VSUBS 0.021297f
C174 B.n47 VSUBS 0.009192f
C175 B.n48 VSUBS 0.009192f
C176 B.n49 VSUBS 0.009192f
C177 B.n50 VSUBS 0.009192f
C178 B.n51 VSUBS 0.009192f
C179 B.n52 VSUBS 0.009192f
C180 B.n53 VSUBS 0.009192f
C181 B.n54 VSUBS 0.020453f
C182 B.n55 VSUBS 0.009192f
C183 B.n56 VSUBS 0.009192f
C184 B.n57 VSUBS 0.009192f
C185 B.n58 VSUBS 0.009192f
C186 B.n59 VSUBS 0.009192f
C187 B.n60 VSUBS 0.009192f
C188 B.n61 VSUBS 0.009192f
C189 B.n62 VSUBS 0.009192f
C190 B.n63 VSUBS 0.009192f
C191 B.n64 VSUBS 0.009192f
C192 B.n65 VSUBS 0.009192f
C193 B.n66 VSUBS 0.009192f
C194 B.n67 VSUBS 0.009192f
C195 B.n68 VSUBS 0.009192f
C196 B.n69 VSUBS 0.009192f
C197 B.n70 VSUBS 0.009192f
C198 B.n71 VSUBS 0.009192f
C199 B.n72 VSUBS 0.009192f
C200 B.n73 VSUBS 0.009192f
C201 B.n74 VSUBS 0.009192f
C202 B.n75 VSUBS 0.009192f
C203 B.n76 VSUBS 0.009192f
C204 B.n77 VSUBS 0.009192f
C205 B.n78 VSUBS 0.009192f
C206 B.n79 VSUBS 0.009192f
C207 B.n80 VSUBS 0.009192f
C208 B.n81 VSUBS 0.009192f
C209 B.n82 VSUBS 0.009192f
C210 B.n83 VSUBS 0.009192f
C211 B.n84 VSUBS 0.009192f
C212 B.n85 VSUBS 0.009192f
C213 B.n86 VSUBS 0.009192f
C214 B.n87 VSUBS 0.009192f
C215 B.n88 VSUBS 0.009192f
C216 B.n89 VSUBS 0.009192f
C217 B.n90 VSUBS 0.009192f
C218 B.n91 VSUBS 0.009192f
C219 B.n92 VSUBS 0.009192f
C220 B.n93 VSUBS 0.009192f
C221 B.n94 VSUBS 0.009192f
C222 B.n95 VSUBS 0.009192f
C223 B.n96 VSUBS 0.009192f
C224 B.n97 VSUBS 0.009192f
C225 B.n98 VSUBS 0.009192f
C226 B.n99 VSUBS 0.009192f
C227 B.n100 VSUBS 0.009192f
C228 B.n101 VSUBS 0.009192f
C229 B.n102 VSUBS 0.009192f
C230 B.n103 VSUBS 0.009192f
C231 B.n104 VSUBS 0.009192f
C232 B.n105 VSUBS 0.020885f
C233 B.n106 VSUBS 0.009192f
C234 B.n107 VSUBS 0.009192f
C235 B.n108 VSUBS 0.009192f
C236 B.n109 VSUBS 0.009192f
C237 B.n110 VSUBS 0.009192f
C238 B.n111 VSUBS 0.009192f
C239 B.n112 VSUBS 0.009192f
C240 B.n113 VSUBS 0.008652f
C241 B.n114 VSUBS 0.009192f
C242 B.n115 VSUBS 0.009192f
C243 B.n116 VSUBS 0.009192f
C244 B.n117 VSUBS 0.009192f
C245 B.n118 VSUBS 0.009192f
C246 B.t8 VSUBS 0.122244f
C247 B.t7 VSUBS 0.14498f
C248 B.t6 VSUBS 0.592166f
C249 B.n119 VSUBS 0.115683f
C250 B.n120 VSUBS 0.088914f
C251 B.n121 VSUBS 0.009192f
C252 B.n122 VSUBS 0.009192f
C253 B.n123 VSUBS 0.009192f
C254 B.n124 VSUBS 0.009192f
C255 B.n125 VSUBS 0.009192f
C256 B.n126 VSUBS 0.009192f
C257 B.n127 VSUBS 0.009192f
C258 B.n128 VSUBS 0.009192f
C259 B.n129 VSUBS 0.020453f
C260 B.n130 VSUBS 0.009192f
C261 B.n131 VSUBS 0.009192f
C262 B.n132 VSUBS 0.009192f
C263 B.n133 VSUBS 0.009192f
C264 B.n134 VSUBS 0.009192f
C265 B.n135 VSUBS 0.009192f
C266 B.n136 VSUBS 0.009192f
C267 B.n137 VSUBS 0.009192f
C268 B.n138 VSUBS 0.009192f
C269 B.n139 VSUBS 0.009192f
C270 B.n140 VSUBS 0.009192f
C271 B.n141 VSUBS 0.009192f
C272 B.n142 VSUBS 0.009192f
C273 B.n143 VSUBS 0.009192f
C274 B.n144 VSUBS 0.009192f
C275 B.n145 VSUBS 0.009192f
C276 B.n146 VSUBS 0.009192f
C277 B.n147 VSUBS 0.009192f
C278 B.n148 VSUBS 0.009192f
C279 B.n149 VSUBS 0.009192f
C280 B.n150 VSUBS 0.009192f
C281 B.n151 VSUBS 0.009192f
C282 B.n152 VSUBS 0.009192f
C283 B.n153 VSUBS 0.009192f
C284 B.n154 VSUBS 0.009192f
C285 B.n155 VSUBS 0.009192f
C286 B.n156 VSUBS 0.009192f
C287 B.n157 VSUBS 0.009192f
C288 B.n158 VSUBS 0.009192f
C289 B.n159 VSUBS 0.009192f
C290 B.n160 VSUBS 0.009192f
C291 B.n161 VSUBS 0.009192f
C292 B.n162 VSUBS 0.009192f
C293 B.n163 VSUBS 0.009192f
C294 B.n164 VSUBS 0.009192f
C295 B.n165 VSUBS 0.009192f
C296 B.n166 VSUBS 0.009192f
C297 B.n167 VSUBS 0.009192f
C298 B.n168 VSUBS 0.009192f
C299 B.n169 VSUBS 0.009192f
C300 B.n170 VSUBS 0.009192f
C301 B.n171 VSUBS 0.009192f
C302 B.n172 VSUBS 0.009192f
C303 B.n173 VSUBS 0.009192f
C304 B.n174 VSUBS 0.009192f
C305 B.n175 VSUBS 0.009192f
C306 B.n176 VSUBS 0.009192f
C307 B.n177 VSUBS 0.009192f
C308 B.n178 VSUBS 0.009192f
C309 B.n179 VSUBS 0.009192f
C310 B.n180 VSUBS 0.009192f
C311 B.n181 VSUBS 0.009192f
C312 B.n182 VSUBS 0.009192f
C313 B.n183 VSUBS 0.009192f
C314 B.n184 VSUBS 0.009192f
C315 B.n185 VSUBS 0.009192f
C316 B.n186 VSUBS 0.009192f
C317 B.n187 VSUBS 0.009192f
C318 B.n188 VSUBS 0.009192f
C319 B.n189 VSUBS 0.009192f
C320 B.n190 VSUBS 0.009192f
C321 B.n191 VSUBS 0.009192f
C322 B.n192 VSUBS 0.009192f
C323 B.n193 VSUBS 0.009192f
C324 B.n194 VSUBS 0.009192f
C325 B.n195 VSUBS 0.009192f
C326 B.n196 VSUBS 0.009192f
C327 B.n197 VSUBS 0.009192f
C328 B.n198 VSUBS 0.009192f
C329 B.n199 VSUBS 0.009192f
C330 B.n200 VSUBS 0.009192f
C331 B.n201 VSUBS 0.009192f
C332 B.n202 VSUBS 0.009192f
C333 B.n203 VSUBS 0.009192f
C334 B.n204 VSUBS 0.009192f
C335 B.n205 VSUBS 0.009192f
C336 B.n206 VSUBS 0.009192f
C337 B.n207 VSUBS 0.009192f
C338 B.n208 VSUBS 0.009192f
C339 B.n209 VSUBS 0.009192f
C340 B.n210 VSUBS 0.009192f
C341 B.n211 VSUBS 0.009192f
C342 B.n212 VSUBS 0.009192f
C343 B.n213 VSUBS 0.009192f
C344 B.n214 VSUBS 0.009192f
C345 B.n215 VSUBS 0.009192f
C346 B.n216 VSUBS 0.009192f
C347 B.n217 VSUBS 0.009192f
C348 B.n218 VSUBS 0.009192f
C349 B.n219 VSUBS 0.009192f
C350 B.n220 VSUBS 0.009192f
C351 B.n221 VSUBS 0.009192f
C352 B.n222 VSUBS 0.009192f
C353 B.n223 VSUBS 0.009192f
C354 B.n224 VSUBS 0.009192f
C355 B.n225 VSUBS 0.009192f
C356 B.n226 VSUBS 0.020453f
C357 B.n227 VSUBS 0.021994f
C358 B.n228 VSUBS 0.021994f
C359 B.n229 VSUBS 0.009192f
C360 B.n230 VSUBS 0.009192f
C361 B.n231 VSUBS 0.009192f
C362 B.n232 VSUBS 0.009192f
C363 B.n233 VSUBS 0.009192f
C364 B.n234 VSUBS 0.009192f
C365 B.n235 VSUBS 0.009192f
C366 B.n236 VSUBS 0.009192f
C367 B.n237 VSUBS 0.009192f
C368 B.n238 VSUBS 0.009192f
C369 B.n239 VSUBS 0.009192f
C370 B.n240 VSUBS 0.009192f
C371 B.n241 VSUBS 0.009192f
C372 B.n242 VSUBS 0.009192f
C373 B.n243 VSUBS 0.009192f
C374 B.n244 VSUBS 0.009192f
C375 B.n245 VSUBS 0.009192f
C376 B.n246 VSUBS 0.009192f
C377 B.n247 VSUBS 0.009192f
C378 B.n248 VSUBS 0.009192f
C379 B.n249 VSUBS 0.009192f
C380 B.n250 VSUBS 0.009192f
C381 B.n251 VSUBS 0.009192f
C382 B.n252 VSUBS 0.008652f
C383 B.n253 VSUBS 0.021297f
C384 B.n254 VSUBS 0.005137f
C385 B.n255 VSUBS 0.009192f
C386 B.n256 VSUBS 0.009192f
C387 B.n257 VSUBS 0.009192f
C388 B.n258 VSUBS 0.009192f
C389 B.n259 VSUBS 0.009192f
C390 B.n260 VSUBS 0.009192f
C391 B.n261 VSUBS 0.009192f
C392 B.n262 VSUBS 0.009192f
C393 B.n263 VSUBS 0.009192f
C394 B.n264 VSUBS 0.009192f
C395 B.n265 VSUBS 0.009192f
C396 B.n266 VSUBS 0.009192f
C397 B.t2 VSUBS 0.122244f
C398 B.t1 VSUBS 0.14498f
C399 B.t0 VSUBS 0.592166f
C400 B.n267 VSUBS 0.115683f
C401 B.n268 VSUBS 0.088914f
C402 B.n269 VSUBS 0.021297f
C403 B.n270 VSUBS 0.005137f
C404 B.n271 VSUBS 0.009192f
C405 B.n272 VSUBS 0.009192f
C406 B.n273 VSUBS 0.009192f
C407 B.n274 VSUBS 0.009192f
C408 B.n275 VSUBS 0.009192f
C409 B.n276 VSUBS 0.009192f
C410 B.n277 VSUBS 0.009192f
C411 B.n278 VSUBS 0.009192f
C412 B.n279 VSUBS 0.009192f
C413 B.n280 VSUBS 0.009192f
C414 B.n281 VSUBS 0.009192f
C415 B.n282 VSUBS 0.009192f
C416 B.n283 VSUBS 0.009192f
C417 B.n284 VSUBS 0.009192f
C418 B.n285 VSUBS 0.009192f
C419 B.n286 VSUBS 0.009192f
C420 B.n287 VSUBS 0.009192f
C421 B.n288 VSUBS 0.009192f
C422 B.n289 VSUBS 0.009192f
C423 B.n290 VSUBS 0.009192f
C424 B.n291 VSUBS 0.009192f
C425 B.n292 VSUBS 0.009192f
C426 B.n293 VSUBS 0.009192f
C427 B.n294 VSUBS 0.009192f
C428 B.n295 VSUBS 0.009192f
C429 B.n296 VSUBS 0.021994f
C430 B.n297 VSUBS 0.020453f
C431 B.n298 VSUBS 0.021561f
C432 B.n299 VSUBS 0.009192f
C433 B.n300 VSUBS 0.009192f
C434 B.n301 VSUBS 0.009192f
C435 B.n302 VSUBS 0.009192f
C436 B.n303 VSUBS 0.009192f
C437 B.n304 VSUBS 0.009192f
C438 B.n305 VSUBS 0.009192f
C439 B.n306 VSUBS 0.009192f
C440 B.n307 VSUBS 0.009192f
C441 B.n308 VSUBS 0.009192f
C442 B.n309 VSUBS 0.009192f
C443 B.n310 VSUBS 0.009192f
C444 B.n311 VSUBS 0.009192f
C445 B.n312 VSUBS 0.009192f
C446 B.n313 VSUBS 0.009192f
C447 B.n314 VSUBS 0.009192f
C448 B.n315 VSUBS 0.009192f
C449 B.n316 VSUBS 0.009192f
C450 B.n317 VSUBS 0.009192f
C451 B.n318 VSUBS 0.009192f
C452 B.n319 VSUBS 0.009192f
C453 B.n320 VSUBS 0.009192f
C454 B.n321 VSUBS 0.009192f
C455 B.n322 VSUBS 0.009192f
C456 B.n323 VSUBS 0.009192f
C457 B.n324 VSUBS 0.009192f
C458 B.n325 VSUBS 0.009192f
C459 B.n326 VSUBS 0.009192f
C460 B.n327 VSUBS 0.009192f
C461 B.n328 VSUBS 0.009192f
C462 B.n329 VSUBS 0.009192f
C463 B.n330 VSUBS 0.009192f
C464 B.n331 VSUBS 0.009192f
C465 B.n332 VSUBS 0.009192f
C466 B.n333 VSUBS 0.009192f
C467 B.n334 VSUBS 0.009192f
C468 B.n335 VSUBS 0.009192f
C469 B.n336 VSUBS 0.009192f
C470 B.n337 VSUBS 0.009192f
C471 B.n338 VSUBS 0.009192f
C472 B.n339 VSUBS 0.009192f
C473 B.n340 VSUBS 0.009192f
C474 B.n341 VSUBS 0.009192f
C475 B.n342 VSUBS 0.009192f
C476 B.n343 VSUBS 0.009192f
C477 B.n344 VSUBS 0.009192f
C478 B.n345 VSUBS 0.009192f
C479 B.n346 VSUBS 0.009192f
C480 B.n347 VSUBS 0.009192f
C481 B.n348 VSUBS 0.009192f
C482 B.n349 VSUBS 0.009192f
C483 B.n350 VSUBS 0.009192f
C484 B.n351 VSUBS 0.009192f
C485 B.n352 VSUBS 0.009192f
C486 B.n353 VSUBS 0.009192f
C487 B.n354 VSUBS 0.009192f
C488 B.n355 VSUBS 0.009192f
C489 B.n356 VSUBS 0.009192f
C490 B.n357 VSUBS 0.009192f
C491 B.n358 VSUBS 0.009192f
C492 B.n359 VSUBS 0.009192f
C493 B.n360 VSUBS 0.009192f
C494 B.n361 VSUBS 0.009192f
C495 B.n362 VSUBS 0.009192f
C496 B.n363 VSUBS 0.009192f
C497 B.n364 VSUBS 0.009192f
C498 B.n365 VSUBS 0.009192f
C499 B.n366 VSUBS 0.009192f
C500 B.n367 VSUBS 0.009192f
C501 B.n368 VSUBS 0.009192f
C502 B.n369 VSUBS 0.009192f
C503 B.n370 VSUBS 0.009192f
C504 B.n371 VSUBS 0.009192f
C505 B.n372 VSUBS 0.009192f
C506 B.n373 VSUBS 0.009192f
C507 B.n374 VSUBS 0.009192f
C508 B.n375 VSUBS 0.009192f
C509 B.n376 VSUBS 0.009192f
C510 B.n377 VSUBS 0.009192f
C511 B.n378 VSUBS 0.009192f
C512 B.n379 VSUBS 0.009192f
C513 B.n380 VSUBS 0.009192f
C514 B.n381 VSUBS 0.009192f
C515 B.n382 VSUBS 0.009192f
C516 B.n383 VSUBS 0.009192f
C517 B.n384 VSUBS 0.009192f
C518 B.n385 VSUBS 0.009192f
C519 B.n386 VSUBS 0.009192f
C520 B.n387 VSUBS 0.009192f
C521 B.n388 VSUBS 0.009192f
C522 B.n389 VSUBS 0.009192f
C523 B.n390 VSUBS 0.009192f
C524 B.n391 VSUBS 0.009192f
C525 B.n392 VSUBS 0.009192f
C526 B.n393 VSUBS 0.009192f
C527 B.n394 VSUBS 0.009192f
C528 B.n395 VSUBS 0.009192f
C529 B.n396 VSUBS 0.009192f
C530 B.n397 VSUBS 0.009192f
C531 B.n398 VSUBS 0.009192f
C532 B.n399 VSUBS 0.009192f
C533 B.n400 VSUBS 0.009192f
C534 B.n401 VSUBS 0.009192f
C535 B.n402 VSUBS 0.009192f
C536 B.n403 VSUBS 0.009192f
C537 B.n404 VSUBS 0.009192f
C538 B.n405 VSUBS 0.009192f
C539 B.n406 VSUBS 0.009192f
C540 B.n407 VSUBS 0.009192f
C541 B.n408 VSUBS 0.009192f
C542 B.n409 VSUBS 0.009192f
C543 B.n410 VSUBS 0.009192f
C544 B.n411 VSUBS 0.009192f
C545 B.n412 VSUBS 0.009192f
C546 B.n413 VSUBS 0.009192f
C547 B.n414 VSUBS 0.009192f
C548 B.n415 VSUBS 0.009192f
C549 B.n416 VSUBS 0.009192f
C550 B.n417 VSUBS 0.009192f
C551 B.n418 VSUBS 0.009192f
C552 B.n419 VSUBS 0.009192f
C553 B.n420 VSUBS 0.009192f
C554 B.n421 VSUBS 0.009192f
C555 B.n422 VSUBS 0.009192f
C556 B.n423 VSUBS 0.009192f
C557 B.n424 VSUBS 0.009192f
C558 B.n425 VSUBS 0.009192f
C559 B.n426 VSUBS 0.009192f
C560 B.n427 VSUBS 0.009192f
C561 B.n428 VSUBS 0.009192f
C562 B.n429 VSUBS 0.009192f
C563 B.n430 VSUBS 0.009192f
C564 B.n431 VSUBS 0.009192f
C565 B.n432 VSUBS 0.009192f
C566 B.n433 VSUBS 0.009192f
C567 B.n434 VSUBS 0.009192f
C568 B.n435 VSUBS 0.009192f
C569 B.n436 VSUBS 0.009192f
C570 B.n437 VSUBS 0.009192f
C571 B.n438 VSUBS 0.009192f
C572 B.n439 VSUBS 0.009192f
C573 B.n440 VSUBS 0.009192f
C574 B.n441 VSUBS 0.009192f
C575 B.n442 VSUBS 0.009192f
C576 B.n443 VSUBS 0.009192f
C577 B.n444 VSUBS 0.009192f
C578 B.n445 VSUBS 0.009192f
C579 B.n446 VSUBS 0.009192f
C580 B.n447 VSUBS 0.009192f
C581 B.n448 VSUBS 0.009192f
C582 B.n449 VSUBS 0.020453f
C583 B.n450 VSUBS 0.021994f
C584 B.n451 VSUBS 0.021994f
C585 B.n452 VSUBS 0.009192f
C586 B.n453 VSUBS 0.009192f
C587 B.n454 VSUBS 0.009192f
C588 B.n455 VSUBS 0.009192f
C589 B.n456 VSUBS 0.009192f
C590 B.n457 VSUBS 0.009192f
C591 B.n458 VSUBS 0.009192f
C592 B.n459 VSUBS 0.009192f
C593 B.n460 VSUBS 0.009192f
C594 B.n461 VSUBS 0.009192f
C595 B.n462 VSUBS 0.009192f
C596 B.n463 VSUBS 0.009192f
C597 B.n464 VSUBS 0.009192f
C598 B.n465 VSUBS 0.009192f
C599 B.n466 VSUBS 0.009192f
C600 B.n467 VSUBS 0.009192f
C601 B.n468 VSUBS 0.009192f
C602 B.n469 VSUBS 0.009192f
C603 B.n470 VSUBS 0.009192f
C604 B.n471 VSUBS 0.009192f
C605 B.n472 VSUBS 0.009192f
C606 B.n473 VSUBS 0.009192f
C607 B.n474 VSUBS 0.008652f
C608 B.n475 VSUBS 0.009192f
C609 B.n476 VSUBS 0.009192f
C610 B.n477 VSUBS 0.009192f
C611 B.n478 VSUBS 0.009192f
C612 B.n479 VSUBS 0.009192f
C613 B.n480 VSUBS 0.009192f
C614 B.n481 VSUBS 0.009192f
C615 B.n482 VSUBS 0.009192f
C616 B.n483 VSUBS 0.009192f
C617 B.n484 VSUBS 0.009192f
C618 B.n485 VSUBS 0.009192f
C619 B.n486 VSUBS 0.009192f
C620 B.n487 VSUBS 0.009192f
C621 B.n488 VSUBS 0.009192f
C622 B.n489 VSUBS 0.009192f
C623 B.n490 VSUBS 0.005137f
C624 B.n491 VSUBS 0.021297f
C625 B.n492 VSUBS 0.008652f
C626 B.n493 VSUBS 0.009192f
C627 B.n494 VSUBS 0.009192f
C628 B.n495 VSUBS 0.009192f
C629 B.n496 VSUBS 0.009192f
C630 B.n497 VSUBS 0.009192f
C631 B.n498 VSUBS 0.009192f
C632 B.n499 VSUBS 0.009192f
C633 B.n500 VSUBS 0.009192f
C634 B.n501 VSUBS 0.009192f
C635 B.n502 VSUBS 0.009192f
C636 B.n503 VSUBS 0.009192f
C637 B.n504 VSUBS 0.009192f
C638 B.n505 VSUBS 0.009192f
C639 B.n506 VSUBS 0.009192f
C640 B.n507 VSUBS 0.009192f
C641 B.n508 VSUBS 0.009192f
C642 B.n509 VSUBS 0.009192f
C643 B.n510 VSUBS 0.009192f
C644 B.n511 VSUBS 0.009192f
C645 B.n512 VSUBS 0.009192f
C646 B.n513 VSUBS 0.009192f
C647 B.n514 VSUBS 0.009192f
C648 B.n515 VSUBS 0.009192f
C649 B.n516 VSUBS 0.021994f
C650 B.n517 VSUBS 0.020453f
C651 B.n518 VSUBS 0.020453f
C652 B.n519 VSUBS 0.009192f
C653 B.n520 VSUBS 0.009192f
C654 B.n521 VSUBS 0.009192f
C655 B.n522 VSUBS 0.009192f
C656 B.n523 VSUBS 0.009192f
C657 B.n524 VSUBS 0.009192f
C658 B.n525 VSUBS 0.009192f
C659 B.n526 VSUBS 0.009192f
C660 B.n527 VSUBS 0.009192f
C661 B.n528 VSUBS 0.009192f
C662 B.n529 VSUBS 0.009192f
C663 B.n530 VSUBS 0.009192f
C664 B.n531 VSUBS 0.009192f
C665 B.n532 VSUBS 0.009192f
C666 B.n533 VSUBS 0.009192f
C667 B.n534 VSUBS 0.009192f
C668 B.n535 VSUBS 0.009192f
C669 B.n536 VSUBS 0.009192f
C670 B.n537 VSUBS 0.009192f
C671 B.n538 VSUBS 0.009192f
C672 B.n539 VSUBS 0.009192f
C673 B.n540 VSUBS 0.009192f
C674 B.n541 VSUBS 0.009192f
C675 B.n542 VSUBS 0.009192f
C676 B.n543 VSUBS 0.009192f
C677 B.n544 VSUBS 0.009192f
C678 B.n545 VSUBS 0.009192f
C679 B.n546 VSUBS 0.009192f
C680 B.n547 VSUBS 0.009192f
C681 B.n548 VSUBS 0.009192f
C682 B.n549 VSUBS 0.009192f
C683 B.n550 VSUBS 0.009192f
C684 B.n551 VSUBS 0.009192f
C685 B.n552 VSUBS 0.009192f
C686 B.n553 VSUBS 0.009192f
C687 B.n554 VSUBS 0.009192f
C688 B.n555 VSUBS 0.009192f
C689 B.n556 VSUBS 0.009192f
C690 B.n557 VSUBS 0.009192f
C691 B.n558 VSUBS 0.009192f
C692 B.n559 VSUBS 0.009192f
C693 B.n560 VSUBS 0.009192f
C694 B.n561 VSUBS 0.009192f
C695 B.n562 VSUBS 0.009192f
C696 B.n563 VSUBS 0.009192f
C697 B.n564 VSUBS 0.009192f
C698 B.n565 VSUBS 0.009192f
C699 B.n566 VSUBS 0.009192f
C700 B.n567 VSUBS 0.009192f
C701 B.n568 VSUBS 0.009192f
C702 B.n569 VSUBS 0.009192f
C703 B.n570 VSUBS 0.009192f
C704 B.n571 VSUBS 0.009192f
C705 B.n572 VSUBS 0.009192f
C706 B.n573 VSUBS 0.009192f
C707 B.n574 VSUBS 0.009192f
C708 B.n575 VSUBS 0.009192f
C709 B.n576 VSUBS 0.009192f
C710 B.n577 VSUBS 0.009192f
C711 B.n578 VSUBS 0.009192f
C712 B.n579 VSUBS 0.009192f
C713 B.n580 VSUBS 0.009192f
C714 B.n581 VSUBS 0.009192f
C715 B.n582 VSUBS 0.009192f
C716 B.n583 VSUBS 0.009192f
C717 B.n584 VSUBS 0.009192f
C718 B.n585 VSUBS 0.009192f
C719 B.n586 VSUBS 0.009192f
C720 B.n587 VSUBS 0.009192f
C721 B.n588 VSUBS 0.009192f
C722 B.n589 VSUBS 0.009192f
C723 B.n590 VSUBS 0.009192f
C724 B.n591 VSUBS 0.011995f
C725 B.n592 VSUBS 0.012778f
C726 B.n593 VSUBS 0.025411f
C727 VDD2.t1 VSUBS 0.069434f
C728 VDD2.t4 VSUBS 0.069434f
C729 VDD2.n0 VSUBS 0.398642f
C730 VDD2.t6 VSUBS 0.069434f
C731 VDD2.t5 VSUBS 0.069434f
C732 VDD2.n1 VSUBS 0.398642f
C733 VDD2.n2 VSUBS 2.91078f
C734 VDD2.t3 VSUBS 0.069434f
C735 VDD2.t7 VSUBS 0.069434f
C736 VDD2.n3 VSUBS 0.392662f
C737 VDD2.n4 VSUBS 2.33357f
C738 VDD2.t0 VSUBS 0.069434f
C739 VDD2.t2 VSUBS 0.069434f
C740 VDD2.n5 VSUBS 0.398621f
C741 VTAIL.t15 VSUBS 0.095161f
C742 VTAIL.t10 VSUBS 0.095161f
C743 VTAIL.n0 VSUBS 0.468479f
C744 VTAIL.n1 VSUBS 0.747139f
C745 VTAIL.t14 VSUBS 0.679184f
C746 VTAIL.n2 VSUBS 0.839725f
C747 VTAIL.t4 VSUBS 0.679184f
C748 VTAIL.n3 VSUBS 0.839725f
C749 VTAIL.t7 VSUBS 0.095161f
C750 VTAIL.t2 VSUBS 0.095161f
C751 VTAIL.n4 VSUBS 0.468479f
C752 VTAIL.n5 VSUBS 1.00581f
C753 VTAIL.t6 VSUBS 0.679184f
C754 VTAIL.n6 VSUBS 1.8373f
C755 VTAIL.t12 VSUBS 0.679187f
C756 VTAIL.n7 VSUBS 1.8373f
C757 VTAIL.t8 VSUBS 0.095161f
C758 VTAIL.t11 VSUBS 0.095161f
C759 VTAIL.n8 VSUBS 0.468481f
C760 VTAIL.n9 VSUBS 1.00581f
C761 VTAIL.t13 VSUBS 0.679187f
C762 VTAIL.n10 VSUBS 0.839721f
C763 VTAIL.t0 VSUBS 0.679187f
C764 VTAIL.n11 VSUBS 0.839721f
C765 VTAIL.t3 VSUBS 0.095161f
C766 VTAIL.t5 VSUBS 0.095161f
C767 VTAIL.n12 VSUBS 0.468481f
C768 VTAIL.n13 VSUBS 1.00581f
C769 VTAIL.t1 VSUBS 0.679184f
C770 VTAIL.n14 VSUBS 1.8373f
C771 VTAIL.t9 VSUBS 0.679184f
C772 VTAIL.n15 VSUBS 1.83111f
C773 VN.n0 VSUBS 0.057422f
C774 VN.t2 VSUBS 1.03637f
C775 VN.n1 VSUBS 0.076342f
C776 VN.n2 VSUBS 0.043555f
C777 VN.t1 VSUBS 1.03637f
C778 VN.n3 VSUBS 0.420249f
C779 VN.n4 VSUBS 0.043555f
C780 VN.n5 VSUBS 0.063582f
C781 VN.n6 VSUBS 0.418365f
C782 VN.t3 VSUBS 1.03637f
C783 VN.t6 VSUBS 1.36427f
C784 VN.n7 VSUBS 0.528636f
C785 VN.n8 VSUBS 0.540706f
C786 VN.n9 VSUBS 0.056726f
C787 VN.n10 VSUBS 0.081175f
C788 VN.n11 VSUBS 0.043555f
C789 VN.n12 VSUBS 0.043555f
C790 VN.n13 VSUBS 0.043555f
C791 VN.n14 VSUBS 0.063582f
C792 VN.n15 VSUBS 0.081175f
C793 VN.n16 VSUBS 0.056726f
C794 VN.n17 VSUBS 0.043555f
C795 VN.n18 VSUBS 0.043555f
C796 VN.n19 VSUBS 0.065543f
C797 VN.n20 VSUBS 0.084429f
C798 VN.n21 VSUBS 0.047567f
C799 VN.n22 VSUBS 0.043555f
C800 VN.n23 VSUBS 0.043555f
C801 VN.n24 VSUBS 0.043555f
C802 VN.n25 VSUBS 0.081175f
C803 VN.n26 VSUBS 0.047909f
C804 VN.n27 VSUBS 0.550456f
C805 VN.n28 VSUBS 0.076001f
C806 VN.n29 VSUBS 0.057422f
C807 VN.t4 VSUBS 1.03637f
C808 VN.n30 VSUBS 0.076342f
C809 VN.n31 VSUBS 0.043555f
C810 VN.t0 VSUBS 1.03637f
C811 VN.n32 VSUBS 0.420249f
C812 VN.n33 VSUBS 0.043555f
C813 VN.n34 VSUBS 0.063582f
C814 VN.n35 VSUBS 0.418365f
C815 VN.t7 VSUBS 1.03637f
C816 VN.t5 VSUBS 1.36427f
C817 VN.n36 VSUBS 0.528636f
C818 VN.n37 VSUBS 0.540706f
C819 VN.n38 VSUBS 0.056726f
C820 VN.n39 VSUBS 0.081175f
C821 VN.n40 VSUBS 0.043555f
C822 VN.n41 VSUBS 0.043555f
C823 VN.n42 VSUBS 0.043555f
C824 VN.n43 VSUBS 0.063582f
C825 VN.n44 VSUBS 0.081175f
C826 VN.n45 VSUBS 0.056726f
C827 VN.n46 VSUBS 0.043555f
C828 VN.n47 VSUBS 0.043555f
C829 VN.n48 VSUBS 0.065543f
C830 VN.n49 VSUBS 0.084429f
C831 VN.n50 VSUBS 0.047567f
C832 VN.n51 VSUBS 0.043555f
C833 VN.n52 VSUBS 0.043555f
C834 VN.n53 VSUBS 0.043555f
C835 VN.n54 VSUBS 0.081175f
C836 VN.n55 VSUBS 0.047909f
C837 VN.n56 VSUBS 0.550456f
C838 VN.n57 VSUBS 2.0449f
.ends

