* NGSPICE file created from diff_pair_sample_1767.ext - technology: sky130A

.subckt diff_pair_sample_1767 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=0 ps=0 w=11.96 l=1.87
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=0 ps=0 w=11.96 l=1.87
X2 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=4.6644 ps=24.7 w=11.96 l=1.87
X3 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=4.6644 ps=24.7 w=11.96 l=1.87
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=4.6644 ps=24.7 w=11.96 l=1.87
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=0 ps=0 w=11.96 l=1.87
X6 VDD1.t0 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=4.6644 ps=24.7 w=11.96 l=1.87
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.6644 pd=24.7 as=0 ps=0 w=11.96 l=1.87
R0 B.n647 B.n646 585
R1 B.n648 B.n647 585
R2 B.n277 B.n88 585
R3 B.n276 B.n275 585
R4 B.n274 B.n273 585
R5 B.n272 B.n271 585
R6 B.n270 B.n269 585
R7 B.n268 B.n267 585
R8 B.n266 B.n265 585
R9 B.n264 B.n263 585
R10 B.n262 B.n261 585
R11 B.n260 B.n259 585
R12 B.n258 B.n257 585
R13 B.n256 B.n255 585
R14 B.n254 B.n253 585
R15 B.n252 B.n251 585
R16 B.n250 B.n249 585
R17 B.n248 B.n247 585
R18 B.n246 B.n245 585
R19 B.n244 B.n243 585
R20 B.n242 B.n241 585
R21 B.n240 B.n239 585
R22 B.n238 B.n237 585
R23 B.n236 B.n235 585
R24 B.n234 B.n233 585
R25 B.n232 B.n231 585
R26 B.n230 B.n229 585
R27 B.n228 B.n227 585
R28 B.n226 B.n225 585
R29 B.n224 B.n223 585
R30 B.n222 B.n221 585
R31 B.n220 B.n219 585
R32 B.n218 B.n217 585
R33 B.n216 B.n215 585
R34 B.n214 B.n213 585
R35 B.n212 B.n211 585
R36 B.n210 B.n209 585
R37 B.n208 B.n207 585
R38 B.n206 B.n205 585
R39 B.n204 B.n203 585
R40 B.n202 B.n201 585
R41 B.n200 B.n199 585
R42 B.n198 B.n197 585
R43 B.n195 B.n194 585
R44 B.n193 B.n192 585
R45 B.n191 B.n190 585
R46 B.n189 B.n188 585
R47 B.n187 B.n186 585
R48 B.n185 B.n184 585
R49 B.n183 B.n182 585
R50 B.n181 B.n180 585
R51 B.n179 B.n178 585
R52 B.n177 B.n176 585
R53 B.n175 B.n174 585
R54 B.n173 B.n172 585
R55 B.n171 B.n170 585
R56 B.n169 B.n168 585
R57 B.n167 B.n166 585
R58 B.n165 B.n164 585
R59 B.n163 B.n162 585
R60 B.n161 B.n160 585
R61 B.n159 B.n158 585
R62 B.n157 B.n156 585
R63 B.n155 B.n154 585
R64 B.n153 B.n152 585
R65 B.n151 B.n150 585
R66 B.n149 B.n148 585
R67 B.n147 B.n146 585
R68 B.n145 B.n144 585
R69 B.n143 B.n142 585
R70 B.n141 B.n140 585
R71 B.n139 B.n138 585
R72 B.n137 B.n136 585
R73 B.n135 B.n134 585
R74 B.n133 B.n132 585
R75 B.n131 B.n130 585
R76 B.n129 B.n128 585
R77 B.n127 B.n126 585
R78 B.n125 B.n124 585
R79 B.n123 B.n122 585
R80 B.n121 B.n120 585
R81 B.n119 B.n118 585
R82 B.n117 B.n116 585
R83 B.n115 B.n114 585
R84 B.n113 B.n112 585
R85 B.n111 B.n110 585
R86 B.n109 B.n108 585
R87 B.n107 B.n106 585
R88 B.n105 B.n104 585
R89 B.n103 B.n102 585
R90 B.n101 B.n100 585
R91 B.n99 B.n98 585
R92 B.n97 B.n96 585
R93 B.n95 B.n94 585
R94 B.n645 B.n41 585
R95 B.n649 B.n41 585
R96 B.n644 B.n40 585
R97 B.n650 B.n40 585
R98 B.n643 B.n642 585
R99 B.n642 B.n36 585
R100 B.n641 B.n35 585
R101 B.n656 B.n35 585
R102 B.n640 B.n34 585
R103 B.n657 B.n34 585
R104 B.n639 B.n33 585
R105 B.n658 B.n33 585
R106 B.n638 B.n637 585
R107 B.n637 B.n32 585
R108 B.n636 B.n28 585
R109 B.n664 B.n28 585
R110 B.n635 B.n27 585
R111 B.n665 B.n27 585
R112 B.n634 B.n26 585
R113 B.n666 B.n26 585
R114 B.n633 B.n632 585
R115 B.n632 B.n22 585
R116 B.n631 B.n21 585
R117 B.n672 B.n21 585
R118 B.n630 B.n20 585
R119 B.n673 B.n20 585
R120 B.n629 B.n19 585
R121 B.n674 B.n19 585
R122 B.n628 B.n627 585
R123 B.n627 B.n15 585
R124 B.n626 B.n14 585
R125 B.n680 B.n14 585
R126 B.n625 B.n13 585
R127 B.n681 B.n13 585
R128 B.n624 B.n12 585
R129 B.n682 B.n12 585
R130 B.n623 B.n622 585
R131 B.n622 B.n8 585
R132 B.n621 B.n7 585
R133 B.n688 B.n7 585
R134 B.n620 B.n6 585
R135 B.n689 B.n6 585
R136 B.n619 B.n5 585
R137 B.n690 B.n5 585
R138 B.n618 B.n617 585
R139 B.n617 B.n4 585
R140 B.n616 B.n278 585
R141 B.n616 B.n615 585
R142 B.n606 B.n279 585
R143 B.n280 B.n279 585
R144 B.n608 B.n607 585
R145 B.n609 B.n608 585
R146 B.n605 B.n284 585
R147 B.n288 B.n284 585
R148 B.n604 B.n603 585
R149 B.n603 B.n602 585
R150 B.n286 B.n285 585
R151 B.n287 B.n286 585
R152 B.n595 B.n594 585
R153 B.n596 B.n595 585
R154 B.n593 B.n293 585
R155 B.n293 B.n292 585
R156 B.n592 B.n591 585
R157 B.n591 B.n590 585
R158 B.n295 B.n294 585
R159 B.n296 B.n295 585
R160 B.n583 B.n582 585
R161 B.n584 B.n583 585
R162 B.n581 B.n301 585
R163 B.n301 B.n300 585
R164 B.n580 B.n579 585
R165 B.n579 B.n578 585
R166 B.n303 B.n302 585
R167 B.n571 B.n303 585
R168 B.n570 B.n569 585
R169 B.n572 B.n570 585
R170 B.n568 B.n308 585
R171 B.n308 B.n307 585
R172 B.n567 B.n566 585
R173 B.n566 B.n565 585
R174 B.n310 B.n309 585
R175 B.n311 B.n310 585
R176 B.n558 B.n557 585
R177 B.n559 B.n558 585
R178 B.n556 B.n316 585
R179 B.n316 B.n315 585
R180 B.n550 B.n549 585
R181 B.n548 B.n364 585
R182 B.n547 B.n363 585
R183 B.n552 B.n363 585
R184 B.n546 B.n545 585
R185 B.n544 B.n543 585
R186 B.n542 B.n541 585
R187 B.n540 B.n539 585
R188 B.n538 B.n537 585
R189 B.n536 B.n535 585
R190 B.n534 B.n533 585
R191 B.n532 B.n531 585
R192 B.n530 B.n529 585
R193 B.n528 B.n527 585
R194 B.n526 B.n525 585
R195 B.n524 B.n523 585
R196 B.n522 B.n521 585
R197 B.n520 B.n519 585
R198 B.n518 B.n517 585
R199 B.n516 B.n515 585
R200 B.n514 B.n513 585
R201 B.n512 B.n511 585
R202 B.n510 B.n509 585
R203 B.n508 B.n507 585
R204 B.n506 B.n505 585
R205 B.n504 B.n503 585
R206 B.n502 B.n501 585
R207 B.n500 B.n499 585
R208 B.n498 B.n497 585
R209 B.n496 B.n495 585
R210 B.n494 B.n493 585
R211 B.n492 B.n491 585
R212 B.n490 B.n489 585
R213 B.n488 B.n487 585
R214 B.n486 B.n485 585
R215 B.n484 B.n483 585
R216 B.n482 B.n481 585
R217 B.n480 B.n479 585
R218 B.n478 B.n477 585
R219 B.n476 B.n475 585
R220 B.n474 B.n473 585
R221 B.n472 B.n471 585
R222 B.n470 B.n469 585
R223 B.n467 B.n466 585
R224 B.n465 B.n464 585
R225 B.n463 B.n462 585
R226 B.n461 B.n460 585
R227 B.n459 B.n458 585
R228 B.n457 B.n456 585
R229 B.n455 B.n454 585
R230 B.n453 B.n452 585
R231 B.n451 B.n450 585
R232 B.n449 B.n448 585
R233 B.n447 B.n446 585
R234 B.n445 B.n444 585
R235 B.n443 B.n442 585
R236 B.n441 B.n440 585
R237 B.n439 B.n438 585
R238 B.n437 B.n436 585
R239 B.n435 B.n434 585
R240 B.n433 B.n432 585
R241 B.n431 B.n430 585
R242 B.n429 B.n428 585
R243 B.n427 B.n426 585
R244 B.n425 B.n424 585
R245 B.n423 B.n422 585
R246 B.n421 B.n420 585
R247 B.n419 B.n418 585
R248 B.n417 B.n416 585
R249 B.n415 B.n414 585
R250 B.n413 B.n412 585
R251 B.n411 B.n410 585
R252 B.n409 B.n408 585
R253 B.n407 B.n406 585
R254 B.n405 B.n404 585
R255 B.n403 B.n402 585
R256 B.n401 B.n400 585
R257 B.n399 B.n398 585
R258 B.n397 B.n396 585
R259 B.n395 B.n394 585
R260 B.n393 B.n392 585
R261 B.n391 B.n390 585
R262 B.n389 B.n388 585
R263 B.n387 B.n386 585
R264 B.n385 B.n384 585
R265 B.n383 B.n382 585
R266 B.n381 B.n380 585
R267 B.n379 B.n378 585
R268 B.n377 B.n376 585
R269 B.n375 B.n374 585
R270 B.n373 B.n372 585
R271 B.n371 B.n370 585
R272 B.n318 B.n317 585
R273 B.n555 B.n554 585
R274 B.n314 B.n313 585
R275 B.n315 B.n314 585
R276 B.n561 B.n560 585
R277 B.n560 B.n559 585
R278 B.n562 B.n312 585
R279 B.n312 B.n311 585
R280 B.n564 B.n563 585
R281 B.n565 B.n564 585
R282 B.n306 B.n305 585
R283 B.n307 B.n306 585
R284 B.n574 B.n573 585
R285 B.n573 B.n572 585
R286 B.n575 B.n304 585
R287 B.n571 B.n304 585
R288 B.n577 B.n576 585
R289 B.n578 B.n577 585
R290 B.n299 B.n298 585
R291 B.n300 B.n299 585
R292 B.n586 B.n585 585
R293 B.n585 B.n584 585
R294 B.n587 B.n297 585
R295 B.n297 B.n296 585
R296 B.n589 B.n588 585
R297 B.n590 B.n589 585
R298 B.n291 B.n290 585
R299 B.n292 B.n291 585
R300 B.n598 B.n597 585
R301 B.n597 B.n596 585
R302 B.n599 B.n289 585
R303 B.n289 B.n287 585
R304 B.n601 B.n600 585
R305 B.n602 B.n601 585
R306 B.n283 B.n282 585
R307 B.n288 B.n283 585
R308 B.n611 B.n610 585
R309 B.n610 B.n609 585
R310 B.n612 B.n281 585
R311 B.n281 B.n280 585
R312 B.n614 B.n613 585
R313 B.n615 B.n614 585
R314 B.n2 B.n0 585
R315 B.n4 B.n2 585
R316 B.n3 B.n1 585
R317 B.n689 B.n3 585
R318 B.n687 B.n686 585
R319 B.n688 B.n687 585
R320 B.n685 B.n9 585
R321 B.n9 B.n8 585
R322 B.n684 B.n683 585
R323 B.n683 B.n682 585
R324 B.n11 B.n10 585
R325 B.n681 B.n11 585
R326 B.n679 B.n678 585
R327 B.n680 B.n679 585
R328 B.n677 B.n16 585
R329 B.n16 B.n15 585
R330 B.n676 B.n675 585
R331 B.n675 B.n674 585
R332 B.n18 B.n17 585
R333 B.n673 B.n18 585
R334 B.n671 B.n670 585
R335 B.n672 B.n671 585
R336 B.n669 B.n23 585
R337 B.n23 B.n22 585
R338 B.n668 B.n667 585
R339 B.n667 B.n666 585
R340 B.n25 B.n24 585
R341 B.n665 B.n25 585
R342 B.n663 B.n662 585
R343 B.n664 B.n663 585
R344 B.n661 B.n29 585
R345 B.n32 B.n29 585
R346 B.n660 B.n659 585
R347 B.n659 B.n658 585
R348 B.n31 B.n30 585
R349 B.n657 B.n31 585
R350 B.n655 B.n654 585
R351 B.n656 B.n655 585
R352 B.n653 B.n37 585
R353 B.n37 B.n36 585
R354 B.n652 B.n651 585
R355 B.n651 B.n650 585
R356 B.n39 B.n38 585
R357 B.n649 B.n39 585
R358 B.n692 B.n691 585
R359 B.n691 B.n690 585
R360 B.n550 B.n314 473.281
R361 B.n94 B.n39 473.281
R362 B.n554 B.n316 473.281
R363 B.n647 B.n41 473.281
R364 B.n367 B.t6 360.733
R365 B.n365 B.t10 360.733
R366 B.n91 B.t13 360.733
R367 B.n89 B.t2 360.733
R368 B.n367 B.t9 323.899
R369 B.n89 B.t4 323.899
R370 B.n365 B.t12 323.899
R371 B.n91 B.t14 323.899
R372 B.n368 B.t8 281.233
R373 B.n90 B.t5 281.233
R374 B.n366 B.t11 281.233
R375 B.n92 B.t15 281.233
R376 B.n648 B.n87 256.663
R377 B.n648 B.n86 256.663
R378 B.n648 B.n85 256.663
R379 B.n648 B.n84 256.663
R380 B.n648 B.n83 256.663
R381 B.n648 B.n82 256.663
R382 B.n648 B.n81 256.663
R383 B.n648 B.n80 256.663
R384 B.n648 B.n79 256.663
R385 B.n648 B.n78 256.663
R386 B.n648 B.n77 256.663
R387 B.n648 B.n76 256.663
R388 B.n648 B.n75 256.663
R389 B.n648 B.n74 256.663
R390 B.n648 B.n73 256.663
R391 B.n648 B.n72 256.663
R392 B.n648 B.n71 256.663
R393 B.n648 B.n70 256.663
R394 B.n648 B.n69 256.663
R395 B.n648 B.n68 256.663
R396 B.n648 B.n67 256.663
R397 B.n648 B.n66 256.663
R398 B.n648 B.n65 256.663
R399 B.n648 B.n64 256.663
R400 B.n648 B.n63 256.663
R401 B.n648 B.n62 256.663
R402 B.n648 B.n61 256.663
R403 B.n648 B.n60 256.663
R404 B.n648 B.n59 256.663
R405 B.n648 B.n58 256.663
R406 B.n648 B.n57 256.663
R407 B.n648 B.n56 256.663
R408 B.n648 B.n55 256.663
R409 B.n648 B.n54 256.663
R410 B.n648 B.n53 256.663
R411 B.n648 B.n52 256.663
R412 B.n648 B.n51 256.663
R413 B.n648 B.n50 256.663
R414 B.n648 B.n49 256.663
R415 B.n648 B.n48 256.663
R416 B.n648 B.n47 256.663
R417 B.n648 B.n46 256.663
R418 B.n648 B.n45 256.663
R419 B.n648 B.n44 256.663
R420 B.n648 B.n43 256.663
R421 B.n648 B.n42 256.663
R422 B.n552 B.n551 256.663
R423 B.n552 B.n319 256.663
R424 B.n552 B.n320 256.663
R425 B.n552 B.n321 256.663
R426 B.n552 B.n322 256.663
R427 B.n552 B.n323 256.663
R428 B.n552 B.n324 256.663
R429 B.n552 B.n325 256.663
R430 B.n552 B.n326 256.663
R431 B.n552 B.n327 256.663
R432 B.n552 B.n328 256.663
R433 B.n552 B.n329 256.663
R434 B.n552 B.n330 256.663
R435 B.n552 B.n331 256.663
R436 B.n552 B.n332 256.663
R437 B.n552 B.n333 256.663
R438 B.n552 B.n334 256.663
R439 B.n552 B.n335 256.663
R440 B.n552 B.n336 256.663
R441 B.n552 B.n337 256.663
R442 B.n552 B.n338 256.663
R443 B.n552 B.n339 256.663
R444 B.n552 B.n340 256.663
R445 B.n552 B.n341 256.663
R446 B.n552 B.n342 256.663
R447 B.n552 B.n343 256.663
R448 B.n552 B.n344 256.663
R449 B.n552 B.n345 256.663
R450 B.n552 B.n346 256.663
R451 B.n552 B.n347 256.663
R452 B.n552 B.n348 256.663
R453 B.n552 B.n349 256.663
R454 B.n552 B.n350 256.663
R455 B.n552 B.n351 256.663
R456 B.n552 B.n352 256.663
R457 B.n552 B.n353 256.663
R458 B.n552 B.n354 256.663
R459 B.n552 B.n355 256.663
R460 B.n552 B.n356 256.663
R461 B.n552 B.n357 256.663
R462 B.n552 B.n358 256.663
R463 B.n552 B.n359 256.663
R464 B.n552 B.n360 256.663
R465 B.n552 B.n361 256.663
R466 B.n552 B.n362 256.663
R467 B.n553 B.n552 256.663
R468 B.n560 B.n314 163.367
R469 B.n560 B.n312 163.367
R470 B.n564 B.n312 163.367
R471 B.n564 B.n306 163.367
R472 B.n573 B.n306 163.367
R473 B.n573 B.n304 163.367
R474 B.n577 B.n304 163.367
R475 B.n577 B.n299 163.367
R476 B.n585 B.n299 163.367
R477 B.n585 B.n297 163.367
R478 B.n589 B.n297 163.367
R479 B.n589 B.n291 163.367
R480 B.n597 B.n291 163.367
R481 B.n597 B.n289 163.367
R482 B.n601 B.n289 163.367
R483 B.n601 B.n283 163.367
R484 B.n610 B.n283 163.367
R485 B.n610 B.n281 163.367
R486 B.n614 B.n281 163.367
R487 B.n614 B.n2 163.367
R488 B.n691 B.n2 163.367
R489 B.n691 B.n3 163.367
R490 B.n687 B.n3 163.367
R491 B.n687 B.n9 163.367
R492 B.n683 B.n9 163.367
R493 B.n683 B.n11 163.367
R494 B.n679 B.n11 163.367
R495 B.n679 B.n16 163.367
R496 B.n675 B.n16 163.367
R497 B.n675 B.n18 163.367
R498 B.n671 B.n18 163.367
R499 B.n671 B.n23 163.367
R500 B.n667 B.n23 163.367
R501 B.n667 B.n25 163.367
R502 B.n663 B.n25 163.367
R503 B.n663 B.n29 163.367
R504 B.n659 B.n29 163.367
R505 B.n659 B.n31 163.367
R506 B.n655 B.n31 163.367
R507 B.n655 B.n37 163.367
R508 B.n651 B.n37 163.367
R509 B.n651 B.n39 163.367
R510 B.n364 B.n363 163.367
R511 B.n545 B.n363 163.367
R512 B.n543 B.n542 163.367
R513 B.n539 B.n538 163.367
R514 B.n535 B.n534 163.367
R515 B.n531 B.n530 163.367
R516 B.n527 B.n526 163.367
R517 B.n523 B.n522 163.367
R518 B.n519 B.n518 163.367
R519 B.n515 B.n514 163.367
R520 B.n511 B.n510 163.367
R521 B.n507 B.n506 163.367
R522 B.n503 B.n502 163.367
R523 B.n499 B.n498 163.367
R524 B.n495 B.n494 163.367
R525 B.n491 B.n490 163.367
R526 B.n487 B.n486 163.367
R527 B.n483 B.n482 163.367
R528 B.n479 B.n478 163.367
R529 B.n475 B.n474 163.367
R530 B.n471 B.n470 163.367
R531 B.n466 B.n465 163.367
R532 B.n462 B.n461 163.367
R533 B.n458 B.n457 163.367
R534 B.n454 B.n453 163.367
R535 B.n450 B.n449 163.367
R536 B.n446 B.n445 163.367
R537 B.n442 B.n441 163.367
R538 B.n438 B.n437 163.367
R539 B.n434 B.n433 163.367
R540 B.n430 B.n429 163.367
R541 B.n426 B.n425 163.367
R542 B.n422 B.n421 163.367
R543 B.n418 B.n417 163.367
R544 B.n414 B.n413 163.367
R545 B.n410 B.n409 163.367
R546 B.n406 B.n405 163.367
R547 B.n402 B.n401 163.367
R548 B.n398 B.n397 163.367
R549 B.n394 B.n393 163.367
R550 B.n390 B.n389 163.367
R551 B.n386 B.n385 163.367
R552 B.n382 B.n381 163.367
R553 B.n378 B.n377 163.367
R554 B.n374 B.n373 163.367
R555 B.n370 B.n318 163.367
R556 B.n558 B.n316 163.367
R557 B.n558 B.n310 163.367
R558 B.n566 B.n310 163.367
R559 B.n566 B.n308 163.367
R560 B.n570 B.n308 163.367
R561 B.n570 B.n303 163.367
R562 B.n579 B.n303 163.367
R563 B.n579 B.n301 163.367
R564 B.n583 B.n301 163.367
R565 B.n583 B.n295 163.367
R566 B.n591 B.n295 163.367
R567 B.n591 B.n293 163.367
R568 B.n595 B.n293 163.367
R569 B.n595 B.n286 163.367
R570 B.n603 B.n286 163.367
R571 B.n603 B.n284 163.367
R572 B.n608 B.n284 163.367
R573 B.n608 B.n279 163.367
R574 B.n616 B.n279 163.367
R575 B.n617 B.n616 163.367
R576 B.n617 B.n5 163.367
R577 B.n6 B.n5 163.367
R578 B.n7 B.n6 163.367
R579 B.n622 B.n7 163.367
R580 B.n622 B.n12 163.367
R581 B.n13 B.n12 163.367
R582 B.n14 B.n13 163.367
R583 B.n627 B.n14 163.367
R584 B.n627 B.n19 163.367
R585 B.n20 B.n19 163.367
R586 B.n21 B.n20 163.367
R587 B.n632 B.n21 163.367
R588 B.n632 B.n26 163.367
R589 B.n27 B.n26 163.367
R590 B.n28 B.n27 163.367
R591 B.n637 B.n28 163.367
R592 B.n637 B.n33 163.367
R593 B.n34 B.n33 163.367
R594 B.n35 B.n34 163.367
R595 B.n642 B.n35 163.367
R596 B.n642 B.n40 163.367
R597 B.n41 B.n40 163.367
R598 B.n98 B.n97 163.367
R599 B.n102 B.n101 163.367
R600 B.n106 B.n105 163.367
R601 B.n110 B.n109 163.367
R602 B.n114 B.n113 163.367
R603 B.n118 B.n117 163.367
R604 B.n122 B.n121 163.367
R605 B.n126 B.n125 163.367
R606 B.n130 B.n129 163.367
R607 B.n134 B.n133 163.367
R608 B.n138 B.n137 163.367
R609 B.n142 B.n141 163.367
R610 B.n146 B.n145 163.367
R611 B.n150 B.n149 163.367
R612 B.n154 B.n153 163.367
R613 B.n158 B.n157 163.367
R614 B.n162 B.n161 163.367
R615 B.n166 B.n165 163.367
R616 B.n170 B.n169 163.367
R617 B.n174 B.n173 163.367
R618 B.n178 B.n177 163.367
R619 B.n182 B.n181 163.367
R620 B.n186 B.n185 163.367
R621 B.n190 B.n189 163.367
R622 B.n194 B.n193 163.367
R623 B.n199 B.n198 163.367
R624 B.n203 B.n202 163.367
R625 B.n207 B.n206 163.367
R626 B.n211 B.n210 163.367
R627 B.n215 B.n214 163.367
R628 B.n219 B.n218 163.367
R629 B.n223 B.n222 163.367
R630 B.n227 B.n226 163.367
R631 B.n231 B.n230 163.367
R632 B.n235 B.n234 163.367
R633 B.n239 B.n238 163.367
R634 B.n243 B.n242 163.367
R635 B.n247 B.n246 163.367
R636 B.n251 B.n250 163.367
R637 B.n255 B.n254 163.367
R638 B.n259 B.n258 163.367
R639 B.n263 B.n262 163.367
R640 B.n267 B.n266 163.367
R641 B.n271 B.n270 163.367
R642 B.n275 B.n274 163.367
R643 B.n647 B.n88 163.367
R644 B.n552 B.n315 81.0565
R645 B.n649 B.n648 81.0565
R646 B.n551 B.n550 71.676
R647 B.n545 B.n319 71.676
R648 B.n542 B.n320 71.676
R649 B.n538 B.n321 71.676
R650 B.n534 B.n322 71.676
R651 B.n530 B.n323 71.676
R652 B.n526 B.n324 71.676
R653 B.n522 B.n325 71.676
R654 B.n518 B.n326 71.676
R655 B.n514 B.n327 71.676
R656 B.n510 B.n328 71.676
R657 B.n506 B.n329 71.676
R658 B.n502 B.n330 71.676
R659 B.n498 B.n331 71.676
R660 B.n494 B.n332 71.676
R661 B.n490 B.n333 71.676
R662 B.n486 B.n334 71.676
R663 B.n482 B.n335 71.676
R664 B.n478 B.n336 71.676
R665 B.n474 B.n337 71.676
R666 B.n470 B.n338 71.676
R667 B.n465 B.n339 71.676
R668 B.n461 B.n340 71.676
R669 B.n457 B.n341 71.676
R670 B.n453 B.n342 71.676
R671 B.n449 B.n343 71.676
R672 B.n445 B.n344 71.676
R673 B.n441 B.n345 71.676
R674 B.n437 B.n346 71.676
R675 B.n433 B.n347 71.676
R676 B.n429 B.n348 71.676
R677 B.n425 B.n349 71.676
R678 B.n421 B.n350 71.676
R679 B.n417 B.n351 71.676
R680 B.n413 B.n352 71.676
R681 B.n409 B.n353 71.676
R682 B.n405 B.n354 71.676
R683 B.n401 B.n355 71.676
R684 B.n397 B.n356 71.676
R685 B.n393 B.n357 71.676
R686 B.n389 B.n358 71.676
R687 B.n385 B.n359 71.676
R688 B.n381 B.n360 71.676
R689 B.n377 B.n361 71.676
R690 B.n373 B.n362 71.676
R691 B.n553 B.n318 71.676
R692 B.n94 B.n42 71.676
R693 B.n98 B.n43 71.676
R694 B.n102 B.n44 71.676
R695 B.n106 B.n45 71.676
R696 B.n110 B.n46 71.676
R697 B.n114 B.n47 71.676
R698 B.n118 B.n48 71.676
R699 B.n122 B.n49 71.676
R700 B.n126 B.n50 71.676
R701 B.n130 B.n51 71.676
R702 B.n134 B.n52 71.676
R703 B.n138 B.n53 71.676
R704 B.n142 B.n54 71.676
R705 B.n146 B.n55 71.676
R706 B.n150 B.n56 71.676
R707 B.n154 B.n57 71.676
R708 B.n158 B.n58 71.676
R709 B.n162 B.n59 71.676
R710 B.n166 B.n60 71.676
R711 B.n170 B.n61 71.676
R712 B.n174 B.n62 71.676
R713 B.n178 B.n63 71.676
R714 B.n182 B.n64 71.676
R715 B.n186 B.n65 71.676
R716 B.n190 B.n66 71.676
R717 B.n194 B.n67 71.676
R718 B.n199 B.n68 71.676
R719 B.n203 B.n69 71.676
R720 B.n207 B.n70 71.676
R721 B.n211 B.n71 71.676
R722 B.n215 B.n72 71.676
R723 B.n219 B.n73 71.676
R724 B.n223 B.n74 71.676
R725 B.n227 B.n75 71.676
R726 B.n231 B.n76 71.676
R727 B.n235 B.n77 71.676
R728 B.n239 B.n78 71.676
R729 B.n243 B.n79 71.676
R730 B.n247 B.n80 71.676
R731 B.n251 B.n81 71.676
R732 B.n255 B.n82 71.676
R733 B.n259 B.n83 71.676
R734 B.n263 B.n84 71.676
R735 B.n267 B.n85 71.676
R736 B.n271 B.n86 71.676
R737 B.n275 B.n87 71.676
R738 B.n88 B.n87 71.676
R739 B.n274 B.n86 71.676
R740 B.n270 B.n85 71.676
R741 B.n266 B.n84 71.676
R742 B.n262 B.n83 71.676
R743 B.n258 B.n82 71.676
R744 B.n254 B.n81 71.676
R745 B.n250 B.n80 71.676
R746 B.n246 B.n79 71.676
R747 B.n242 B.n78 71.676
R748 B.n238 B.n77 71.676
R749 B.n234 B.n76 71.676
R750 B.n230 B.n75 71.676
R751 B.n226 B.n74 71.676
R752 B.n222 B.n73 71.676
R753 B.n218 B.n72 71.676
R754 B.n214 B.n71 71.676
R755 B.n210 B.n70 71.676
R756 B.n206 B.n69 71.676
R757 B.n202 B.n68 71.676
R758 B.n198 B.n67 71.676
R759 B.n193 B.n66 71.676
R760 B.n189 B.n65 71.676
R761 B.n185 B.n64 71.676
R762 B.n181 B.n63 71.676
R763 B.n177 B.n62 71.676
R764 B.n173 B.n61 71.676
R765 B.n169 B.n60 71.676
R766 B.n165 B.n59 71.676
R767 B.n161 B.n58 71.676
R768 B.n157 B.n57 71.676
R769 B.n153 B.n56 71.676
R770 B.n149 B.n55 71.676
R771 B.n145 B.n54 71.676
R772 B.n141 B.n53 71.676
R773 B.n137 B.n52 71.676
R774 B.n133 B.n51 71.676
R775 B.n129 B.n50 71.676
R776 B.n125 B.n49 71.676
R777 B.n121 B.n48 71.676
R778 B.n117 B.n47 71.676
R779 B.n113 B.n46 71.676
R780 B.n109 B.n45 71.676
R781 B.n105 B.n44 71.676
R782 B.n101 B.n43 71.676
R783 B.n97 B.n42 71.676
R784 B.n551 B.n364 71.676
R785 B.n543 B.n319 71.676
R786 B.n539 B.n320 71.676
R787 B.n535 B.n321 71.676
R788 B.n531 B.n322 71.676
R789 B.n527 B.n323 71.676
R790 B.n523 B.n324 71.676
R791 B.n519 B.n325 71.676
R792 B.n515 B.n326 71.676
R793 B.n511 B.n327 71.676
R794 B.n507 B.n328 71.676
R795 B.n503 B.n329 71.676
R796 B.n499 B.n330 71.676
R797 B.n495 B.n331 71.676
R798 B.n491 B.n332 71.676
R799 B.n487 B.n333 71.676
R800 B.n483 B.n334 71.676
R801 B.n479 B.n335 71.676
R802 B.n475 B.n336 71.676
R803 B.n471 B.n337 71.676
R804 B.n466 B.n338 71.676
R805 B.n462 B.n339 71.676
R806 B.n458 B.n340 71.676
R807 B.n454 B.n341 71.676
R808 B.n450 B.n342 71.676
R809 B.n446 B.n343 71.676
R810 B.n442 B.n344 71.676
R811 B.n438 B.n345 71.676
R812 B.n434 B.n346 71.676
R813 B.n430 B.n347 71.676
R814 B.n426 B.n348 71.676
R815 B.n422 B.n349 71.676
R816 B.n418 B.n350 71.676
R817 B.n414 B.n351 71.676
R818 B.n410 B.n352 71.676
R819 B.n406 B.n353 71.676
R820 B.n402 B.n354 71.676
R821 B.n398 B.n355 71.676
R822 B.n394 B.n356 71.676
R823 B.n390 B.n357 71.676
R824 B.n386 B.n358 71.676
R825 B.n382 B.n359 71.676
R826 B.n378 B.n360 71.676
R827 B.n374 B.n361 71.676
R828 B.n370 B.n362 71.676
R829 B.n554 B.n553 71.676
R830 B.n369 B.n368 59.5399
R831 B.n468 B.n366 59.5399
R832 B.n93 B.n92 59.5399
R833 B.n196 B.n90 59.5399
R834 B.n559 B.n315 43.4006
R835 B.n559 B.n311 43.4006
R836 B.n565 B.n311 43.4006
R837 B.n565 B.n307 43.4006
R838 B.n572 B.n307 43.4006
R839 B.n572 B.n571 43.4006
R840 B.n578 B.n300 43.4006
R841 B.n584 B.n300 43.4006
R842 B.n584 B.n296 43.4006
R843 B.n590 B.n296 43.4006
R844 B.n590 B.n292 43.4006
R845 B.n596 B.n292 43.4006
R846 B.n596 B.n287 43.4006
R847 B.n602 B.n287 43.4006
R848 B.n602 B.n288 43.4006
R849 B.n609 B.n280 43.4006
R850 B.n615 B.n280 43.4006
R851 B.n615 B.n4 43.4006
R852 B.n690 B.n4 43.4006
R853 B.n690 B.n689 43.4006
R854 B.n689 B.n688 43.4006
R855 B.n688 B.n8 43.4006
R856 B.n682 B.n8 43.4006
R857 B.n681 B.n680 43.4006
R858 B.n680 B.n15 43.4006
R859 B.n674 B.n15 43.4006
R860 B.n674 B.n673 43.4006
R861 B.n673 B.n672 43.4006
R862 B.n672 B.n22 43.4006
R863 B.n666 B.n22 43.4006
R864 B.n666 B.n665 43.4006
R865 B.n665 B.n664 43.4006
R866 B.n658 B.n32 43.4006
R867 B.n658 B.n657 43.4006
R868 B.n657 B.n656 43.4006
R869 B.n656 B.n36 43.4006
R870 B.n650 B.n36 43.4006
R871 B.n650 B.n649 43.4006
R872 B.n368 B.n367 42.6672
R873 B.n366 B.n365 42.6672
R874 B.n92 B.n91 42.6672
R875 B.n90 B.n89 42.6672
R876 B.n609 B.t0 36.38
R877 B.n682 B.t1 36.38
R878 B.n646 B.n645 30.7517
R879 B.n95 B.n38 30.7517
R880 B.n556 B.n555 30.7517
R881 B.n549 B.n313 30.7517
R882 B.n578 B.t7 22.3388
R883 B.n664 B.t3 22.3388
R884 B.n571 B.t7 21.0623
R885 B.n32 B.t3 21.0623
R886 B B.n692 18.0485
R887 B.n96 B.n95 10.6151
R888 B.n99 B.n96 10.6151
R889 B.n100 B.n99 10.6151
R890 B.n103 B.n100 10.6151
R891 B.n104 B.n103 10.6151
R892 B.n107 B.n104 10.6151
R893 B.n108 B.n107 10.6151
R894 B.n111 B.n108 10.6151
R895 B.n112 B.n111 10.6151
R896 B.n115 B.n112 10.6151
R897 B.n116 B.n115 10.6151
R898 B.n119 B.n116 10.6151
R899 B.n120 B.n119 10.6151
R900 B.n123 B.n120 10.6151
R901 B.n124 B.n123 10.6151
R902 B.n127 B.n124 10.6151
R903 B.n128 B.n127 10.6151
R904 B.n131 B.n128 10.6151
R905 B.n132 B.n131 10.6151
R906 B.n135 B.n132 10.6151
R907 B.n136 B.n135 10.6151
R908 B.n139 B.n136 10.6151
R909 B.n140 B.n139 10.6151
R910 B.n143 B.n140 10.6151
R911 B.n144 B.n143 10.6151
R912 B.n147 B.n144 10.6151
R913 B.n148 B.n147 10.6151
R914 B.n151 B.n148 10.6151
R915 B.n152 B.n151 10.6151
R916 B.n155 B.n152 10.6151
R917 B.n156 B.n155 10.6151
R918 B.n159 B.n156 10.6151
R919 B.n160 B.n159 10.6151
R920 B.n163 B.n160 10.6151
R921 B.n164 B.n163 10.6151
R922 B.n167 B.n164 10.6151
R923 B.n168 B.n167 10.6151
R924 B.n171 B.n168 10.6151
R925 B.n172 B.n171 10.6151
R926 B.n175 B.n172 10.6151
R927 B.n176 B.n175 10.6151
R928 B.n180 B.n179 10.6151
R929 B.n183 B.n180 10.6151
R930 B.n184 B.n183 10.6151
R931 B.n187 B.n184 10.6151
R932 B.n188 B.n187 10.6151
R933 B.n191 B.n188 10.6151
R934 B.n192 B.n191 10.6151
R935 B.n195 B.n192 10.6151
R936 B.n200 B.n197 10.6151
R937 B.n201 B.n200 10.6151
R938 B.n204 B.n201 10.6151
R939 B.n205 B.n204 10.6151
R940 B.n208 B.n205 10.6151
R941 B.n209 B.n208 10.6151
R942 B.n212 B.n209 10.6151
R943 B.n213 B.n212 10.6151
R944 B.n216 B.n213 10.6151
R945 B.n217 B.n216 10.6151
R946 B.n220 B.n217 10.6151
R947 B.n221 B.n220 10.6151
R948 B.n224 B.n221 10.6151
R949 B.n225 B.n224 10.6151
R950 B.n228 B.n225 10.6151
R951 B.n229 B.n228 10.6151
R952 B.n232 B.n229 10.6151
R953 B.n233 B.n232 10.6151
R954 B.n236 B.n233 10.6151
R955 B.n237 B.n236 10.6151
R956 B.n240 B.n237 10.6151
R957 B.n241 B.n240 10.6151
R958 B.n244 B.n241 10.6151
R959 B.n245 B.n244 10.6151
R960 B.n248 B.n245 10.6151
R961 B.n249 B.n248 10.6151
R962 B.n252 B.n249 10.6151
R963 B.n253 B.n252 10.6151
R964 B.n256 B.n253 10.6151
R965 B.n257 B.n256 10.6151
R966 B.n260 B.n257 10.6151
R967 B.n261 B.n260 10.6151
R968 B.n264 B.n261 10.6151
R969 B.n265 B.n264 10.6151
R970 B.n268 B.n265 10.6151
R971 B.n269 B.n268 10.6151
R972 B.n272 B.n269 10.6151
R973 B.n273 B.n272 10.6151
R974 B.n276 B.n273 10.6151
R975 B.n277 B.n276 10.6151
R976 B.n646 B.n277 10.6151
R977 B.n557 B.n556 10.6151
R978 B.n557 B.n309 10.6151
R979 B.n567 B.n309 10.6151
R980 B.n568 B.n567 10.6151
R981 B.n569 B.n568 10.6151
R982 B.n569 B.n302 10.6151
R983 B.n580 B.n302 10.6151
R984 B.n581 B.n580 10.6151
R985 B.n582 B.n581 10.6151
R986 B.n582 B.n294 10.6151
R987 B.n592 B.n294 10.6151
R988 B.n593 B.n592 10.6151
R989 B.n594 B.n593 10.6151
R990 B.n594 B.n285 10.6151
R991 B.n604 B.n285 10.6151
R992 B.n605 B.n604 10.6151
R993 B.n607 B.n605 10.6151
R994 B.n607 B.n606 10.6151
R995 B.n606 B.n278 10.6151
R996 B.n618 B.n278 10.6151
R997 B.n619 B.n618 10.6151
R998 B.n620 B.n619 10.6151
R999 B.n621 B.n620 10.6151
R1000 B.n623 B.n621 10.6151
R1001 B.n624 B.n623 10.6151
R1002 B.n625 B.n624 10.6151
R1003 B.n626 B.n625 10.6151
R1004 B.n628 B.n626 10.6151
R1005 B.n629 B.n628 10.6151
R1006 B.n630 B.n629 10.6151
R1007 B.n631 B.n630 10.6151
R1008 B.n633 B.n631 10.6151
R1009 B.n634 B.n633 10.6151
R1010 B.n635 B.n634 10.6151
R1011 B.n636 B.n635 10.6151
R1012 B.n638 B.n636 10.6151
R1013 B.n639 B.n638 10.6151
R1014 B.n640 B.n639 10.6151
R1015 B.n641 B.n640 10.6151
R1016 B.n643 B.n641 10.6151
R1017 B.n644 B.n643 10.6151
R1018 B.n645 B.n644 10.6151
R1019 B.n549 B.n548 10.6151
R1020 B.n548 B.n547 10.6151
R1021 B.n547 B.n546 10.6151
R1022 B.n546 B.n544 10.6151
R1023 B.n544 B.n541 10.6151
R1024 B.n541 B.n540 10.6151
R1025 B.n540 B.n537 10.6151
R1026 B.n537 B.n536 10.6151
R1027 B.n536 B.n533 10.6151
R1028 B.n533 B.n532 10.6151
R1029 B.n532 B.n529 10.6151
R1030 B.n529 B.n528 10.6151
R1031 B.n528 B.n525 10.6151
R1032 B.n525 B.n524 10.6151
R1033 B.n524 B.n521 10.6151
R1034 B.n521 B.n520 10.6151
R1035 B.n520 B.n517 10.6151
R1036 B.n517 B.n516 10.6151
R1037 B.n516 B.n513 10.6151
R1038 B.n513 B.n512 10.6151
R1039 B.n512 B.n509 10.6151
R1040 B.n509 B.n508 10.6151
R1041 B.n508 B.n505 10.6151
R1042 B.n505 B.n504 10.6151
R1043 B.n504 B.n501 10.6151
R1044 B.n501 B.n500 10.6151
R1045 B.n500 B.n497 10.6151
R1046 B.n497 B.n496 10.6151
R1047 B.n496 B.n493 10.6151
R1048 B.n493 B.n492 10.6151
R1049 B.n492 B.n489 10.6151
R1050 B.n489 B.n488 10.6151
R1051 B.n488 B.n485 10.6151
R1052 B.n485 B.n484 10.6151
R1053 B.n484 B.n481 10.6151
R1054 B.n481 B.n480 10.6151
R1055 B.n480 B.n477 10.6151
R1056 B.n477 B.n476 10.6151
R1057 B.n476 B.n473 10.6151
R1058 B.n473 B.n472 10.6151
R1059 B.n472 B.n469 10.6151
R1060 B.n467 B.n464 10.6151
R1061 B.n464 B.n463 10.6151
R1062 B.n463 B.n460 10.6151
R1063 B.n460 B.n459 10.6151
R1064 B.n459 B.n456 10.6151
R1065 B.n456 B.n455 10.6151
R1066 B.n455 B.n452 10.6151
R1067 B.n452 B.n451 10.6151
R1068 B.n448 B.n447 10.6151
R1069 B.n447 B.n444 10.6151
R1070 B.n444 B.n443 10.6151
R1071 B.n443 B.n440 10.6151
R1072 B.n440 B.n439 10.6151
R1073 B.n439 B.n436 10.6151
R1074 B.n436 B.n435 10.6151
R1075 B.n435 B.n432 10.6151
R1076 B.n432 B.n431 10.6151
R1077 B.n431 B.n428 10.6151
R1078 B.n428 B.n427 10.6151
R1079 B.n427 B.n424 10.6151
R1080 B.n424 B.n423 10.6151
R1081 B.n423 B.n420 10.6151
R1082 B.n420 B.n419 10.6151
R1083 B.n419 B.n416 10.6151
R1084 B.n416 B.n415 10.6151
R1085 B.n415 B.n412 10.6151
R1086 B.n412 B.n411 10.6151
R1087 B.n411 B.n408 10.6151
R1088 B.n408 B.n407 10.6151
R1089 B.n407 B.n404 10.6151
R1090 B.n404 B.n403 10.6151
R1091 B.n403 B.n400 10.6151
R1092 B.n400 B.n399 10.6151
R1093 B.n399 B.n396 10.6151
R1094 B.n396 B.n395 10.6151
R1095 B.n395 B.n392 10.6151
R1096 B.n392 B.n391 10.6151
R1097 B.n391 B.n388 10.6151
R1098 B.n388 B.n387 10.6151
R1099 B.n387 B.n384 10.6151
R1100 B.n384 B.n383 10.6151
R1101 B.n383 B.n380 10.6151
R1102 B.n380 B.n379 10.6151
R1103 B.n379 B.n376 10.6151
R1104 B.n376 B.n375 10.6151
R1105 B.n375 B.n372 10.6151
R1106 B.n372 B.n371 10.6151
R1107 B.n371 B.n317 10.6151
R1108 B.n555 B.n317 10.6151
R1109 B.n561 B.n313 10.6151
R1110 B.n562 B.n561 10.6151
R1111 B.n563 B.n562 10.6151
R1112 B.n563 B.n305 10.6151
R1113 B.n574 B.n305 10.6151
R1114 B.n575 B.n574 10.6151
R1115 B.n576 B.n575 10.6151
R1116 B.n576 B.n298 10.6151
R1117 B.n586 B.n298 10.6151
R1118 B.n587 B.n586 10.6151
R1119 B.n588 B.n587 10.6151
R1120 B.n588 B.n290 10.6151
R1121 B.n598 B.n290 10.6151
R1122 B.n599 B.n598 10.6151
R1123 B.n600 B.n599 10.6151
R1124 B.n600 B.n282 10.6151
R1125 B.n611 B.n282 10.6151
R1126 B.n612 B.n611 10.6151
R1127 B.n613 B.n612 10.6151
R1128 B.n613 B.n0 10.6151
R1129 B.n686 B.n1 10.6151
R1130 B.n686 B.n685 10.6151
R1131 B.n685 B.n684 10.6151
R1132 B.n684 B.n10 10.6151
R1133 B.n678 B.n10 10.6151
R1134 B.n678 B.n677 10.6151
R1135 B.n677 B.n676 10.6151
R1136 B.n676 B.n17 10.6151
R1137 B.n670 B.n17 10.6151
R1138 B.n670 B.n669 10.6151
R1139 B.n669 B.n668 10.6151
R1140 B.n668 B.n24 10.6151
R1141 B.n662 B.n24 10.6151
R1142 B.n662 B.n661 10.6151
R1143 B.n661 B.n660 10.6151
R1144 B.n660 B.n30 10.6151
R1145 B.n654 B.n30 10.6151
R1146 B.n654 B.n653 10.6151
R1147 B.n653 B.n652 10.6151
R1148 B.n652 B.n38 10.6151
R1149 B.n288 B.t0 7.0211
R1150 B.t1 B.n681 7.0211
R1151 B.n179 B.n93 6.5566
R1152 B.n196 B.n195 6.5566
R1153 B.n468 B.n467 6.5566
R1154 B.n451 B.n369 6.5566
R1155 B.n176 B.n93 4.05904
R1156 B.n197 B.n196 4.05904
R1157 B.n469 B.n468 4.05904
R1158 B.n448 B.n369 4.05904
R1159 B.n692 B.n0 2.81026
R1160 B.n692 B.n1 2.81026
R1161 VN VN.t1 255.855
R1162 VN VN.t0 213.214
R1163 VTAIL.n262 VTAIL.n261 289.615
R1164 VTAIL.n64 VTAIL.n63 289.615
R1165 VTAIL.n196 VTAIL.n195 289.615
R1166 VTAIL.n130 VTAIL.n129 289.615
R1167 VTAIL.n221 VTAIL.n220 185
R1168 VTAIL.n223 VTAIL.n222 185
R1169 VTAIL.n216 VTAIL.n215 185
R1170 VTAIL.n229 VTAIL.n228 185
R1171 VTAIL.n231 VTAIL.n230 185
R1172 VTAIL.n212 VTAIL.n211 185
R1173 VTAIL.n237 VTAIL.n236 185
R1174 VTAIL.n239 VTAIL.n238 185
R1175 VTAIL.n208 VTAIL.n207 185
R1176 VTAIL.n245 VTAIL.n244 185
R1177 VTAIL.n247 VTAIL.n246 185
R1178 VTAIL.n204 VTAIL.n203 185
R1179 VTAIL.n253 VTAIL.n252 185
R1180 VTAIL.n255 VTAIL.n254 185
R1181 VTAIL.n200 VTAIL.n199 185
R1182 VTAIL.n261 VTAIL.n260 185
R1183 VTAIL.n23 VTAIL.n22 185
R1184 VTAIL.n25 VTAIL.n24 185
R1185 VTAIL.n18 VTAIL.n17 185
R1186 VTAIL.n31 VTAIL.n30 185
R1187 VTAIL.n33 VTAIL.n32 185
R1188 VTAIL.n14 VTAIL.n13 185
R1189 VTAIL.n39 VTAIL.n38 185
R1190 VTAIL.n41 VTAIL.n40 185
R1191 VTAIL.n10 VTAIL.n9 185
R1192 VTAIL.n47 VTAIL.n46 185
R1193 VTAIL.n49 VTAIL.n48 185
R1194 VTAIL.n6 VTAIL.n5 185
R1195 VTAIL.n55 VTAIL.n54 185
R1196 VTAIL.n57 VTAIL.n56 185
R1197 VTAIL.n2 VTAIL.n1 185
R1198 VTAIL.n63 VTAIL.n62 185
R1199 VTAIL.n195 VTAIL.n194 185
R1200 VTAIL.n134 VTAIL.n133 185
R1201 VTAIL.n189 VTAIL.n188 185
R1202 VTAIL.n187 VTAIL.n186 185
R1203 VTAIL.n138 VTAIL.n137 185
R1204 VTAIL.n181 VTAIL.n180 185
R1205 VTAIL.n179 VTAIL.n178 185
R1206 VTAIL.n142 VTAIL.n141 185
R1207 VTAIL.n173 VTAIL.n172 185
R1208 VTAIL.n171 VTAIL.n170 185
R1209 VTAIL.n146 VTAIL.n145 185
R1210 VTAIL.n165 VTAIL.n164 185
R1211 VTAIL.n163 VTAIL.n162 185
R1212 VTAIL.n150 VTAIL.n149 185
R1213 VTAIL.n157 VTAIL.n156 185
R1214 VTAIL.n155 VTAIL.n154 185
R1215 VTAIL.n129 VTAIL.n128 185
R1216 VTAIL.n68 VTAIL.n67 185
R1217 VTAIL.n123 VTAIL.n122 185
R1218 VTAIL.n121 VTAIL.n120 185
R1219 VTAIL.n72 VTAIL.n71 185
R1220 VTAIL.n115 VTAIL.n114 185
R1221 VTAIL.n113 VTAIL.n112 185
R1222 VTAIL.n76 VTAIL.n75 185
R1223 VTAIL.n107 VTAIL.n106 185
R1224 VTAIL.n105 VTAIL.n104 185
R1225 VTAIL.n80 VTAIL.n79 185
R1226 VTAIL.n99 VTAIL.n98 185
R1227 VTAIL.n97 VTAIL.n96 185
R1228 VTAIL.n84 VTAIL.n83 185
R1229 VTAIL.n91 VTAIL.n90 185
R1230 VTAIL.n89 VTAIL.n88 185
R1231 VTAIL.n87 VTAIL.t2 147.659
R1232 VTAIL.n219 VTAIL.t3 147.659
R1233 VTAIL.n21 VTAIL.t1 147.659
R1234 VTAIL.n153 VTAIL.t0 147.659
R1235 VTAIL.n222 VTAIL.n221 104.615
R1236 VTAIL.n222 VTAIL.n215 104.615
R1237 VTAIL.n229 VTAIL.n215 104.615
R1238 VTAIL.n230 VTAIL.n229 104.615
R1239 VTAIL.n230 VTAIL.n211 104.615
R1240 VTAIL.n237 VTAIL.n211 104.615
R1241 VTAIL.n238 VTAIL.n237 104.615
R1242 VTAIL.n238 VTAIL.n207 104.615
R1243 VTAIL.n245 VTAIL.n207 104.615
R1244 VTAIL.n246 VTAIL.n245 104.615
R1245 VTAIL.n246 VTAIL.n203 104.615
R1246 VTAIL.n253 VTAIL.n203 104.615
R1247 VTAIL.n254 VTAIL.n253 104.615
R1248 VTAIL.n254 VTAIL.n199 104.615
R1249 VTAIL.n261 VTAIL.n199 104.615
R1250 VTAIL.n24 VTAIL.n23 104.615
R1251 VTAIL.n24 VTAIL.n17 104.615
R1252 VTAIL.n31 VTAIL.n17 104.615
R1253 VTAIL.n32 VTAIL.n31 104.615
R1254 VTAIL.n32 VTAIL.n13 104.615
R1255 VTAIL.n39 VTAIL.n13 104.615
R1256 VTAIL.n40 VTAIL.n39 104.615
R1257 VTAIL.n40 VTAIL.n9 104.615
R1258 VTAIL.n47 VTAIL.n9 104.615
R1259 VTAIL.n48 VTAIL.n47 104.615
R1260 VTAIL.n48 VTAIL.n5 104.615
R1261 VTAIL.n55 VTAIL.n5 104.615
R1262 VTAIL.n56 VTAIL.n55 104.615
R1263 VTAIL.n56 VTAIL.n1 104.615
R1264 VTAIL.n63 VTAIL.n1 104.615
R1265 VTAIL.n195 VTAIL.n133 104.615
R1266 VTAIL.n188 VTAIL.n133 104.615
R1267 VTAIL.n188 VTAIL.n187 104.615
R1268 VTAIL.n187 VTAIL.n137 104.615
R1269 VTAIL.n180 VTAIL.n137 104.615
R1270 VTAIL.n180 VTAIL.n179 104.615
R1271 VTAIL.n179 VTAIL.n141 104.615
R1272 VTAIL.n172 VTAIL.n141 104.615
R1273 VTAIL.n172 VTAIL.n171 104.615
R1274 VTAIL.n171 VTAIL.n145 104.615
R1275 VTAIL.n164 VTAIL.n145 104.615
R1276 VTAIL.n164 VTAIL.n163 104.615
R1277 VTAIL.n163 VTAIL.n149 104.615
R1278 VTAIL.n156 VTAIL.n149 104.615
R1279 VTAIL.n156 VTAIL.n155 104.615
R1280 VTAIL.n129 VTAIL.n67 104.615
R1281 VTAIL.n122 VTAIL.n67 104.615
R1282 VTAIL.n122 VTAIL.n121 104.615
R1283 VTAIL.n121 VTAIL.n71 104.615
R1284 VTAIL.n114 VTAIL.n71 104.615
R1285 VTAIL.n114 VTAIL.n113 104.615
R1286 VTAIL.n113 VTAIL.n75 104.615
R1287 VTAIL.n106 VTAIL.n75 104.615
R1288 VTAIL.n106 VTAIL.n105 104.615
R1289 VTAIL.n105 VTAIL.n79 104.615
R1290 VTAIL.n98 VTAIL.n79 104.615
R1291 VTAIL.n98 VTAIL.n97 104.615
R1292 VTAIL.n97 VTAIL.n83 104.615
R1293 VTAIL.n90 VTAIL.n83 104.615
R1294 VTAIL.n90 VTAIL.n89 104.615
R1295 VTAIL.n221 VTAIL.t3 52.3082
R1296 VTAIL.n23 VTAIL.t1 52.3082
R1297 VTAIL.n155 VTAIL.t0 52.3082
R1298 VTAIL.n89 VTAIL.t2 52.3082
R1299 VTAIL.n263 VTAIL.n262 34.9005
R1300 VTAIL.n65 VTAIL.n64 34.9005
R1301 VTAIL.n197 VTAIL.n196 34.9005
R1302 VTAIL.n131 VTAIL.n130 34.9005
R1303 VTAIL.n131 VTAIL.n65 26.4703
R1304 VTAIL.n263 VTAIL.n197 24.5738
R1305 VTAIL.n220 VTAIL.n219 15.6677
R1306 VTAIL.n22 VTAIL.n21 15.6677
R1307 VTAIL.n154 VTAIL.n153 15.6677
R1308 VTAIL.n88 VTAIL.n87 15.6677
R1309 VTAIL.n223 VTAIL.n218 12.8005
R1310 VTAIL.n25 VTAIL.n20 12.8005
R1311 VTAIL.n157 VTAIL.n152 12.8005
R1312 VTAIL.n91 VTAIL.n86 12.8005
R1313 VTAIL.n224 VTAIL.n216 12.0247
R1314 VTAIL.n260 VTAIL.n198 12.0247
R1315 VTAIL.n26 VTAIL.n18 12.0247
R1316 VTAIL.n62 VTAIL.n0 12.0247
R1317 VTAIL.n194 VTAIL.n132 12.0247
R1318 VTAIL.n158 VTAIL.n150 12.0247
R1319 VTAIL.n128 VTAIL.n66 12.0247
R1320 VTAIL.n92 VTAIL.n84 12.0247
R1321 VTAIL.n228 VTAIL.n227 11.249
R1322 VTAIL.n259 VTAIL.n200 11.249
R1323 VTAIL.n30 VTAIL.n29 11.249
R1324 VTAIL.n61 VTAIL.n2 11.249
R1325 VTAIL.n193 VTAIL.n134 11.249
R1326 VTAIL.n162 VTAIL.n161 11.249
R1327 VTAIL.n127 VTAIL.n68 11.249
R1328 VTAIL.n96 VTAIL.n95 11.249
R1329 VTAIL.n231 VTAIL.n214 10.4732
R1330 VTAIL.n256 VTAIL.n255 10.4732
R1331 VTAIL.n33 VTAIL.n16 10.4732
R1332 VTAIL.n58 VTAIL.n57 10.4732
R1333 VTAIL.n190 VTAIL.n189 10.4732
R1334 VTAIL.n165 VTAIL.n148 10.4732
R1335 VTAIL.n124 VTAIL.n123 10.4732
R1336 VTAIL.n99 VTAIL.n82 10.4732
R1337 VTAIL.n232 VTAIL.n212 9.69747
R1338 VTAIL.n252 VTAIL.n202 9.69747
R1339 VTAIL.n34 VTAIL.n14 9.69747
R1340 VTAIL.n54 VTAIL.n4 9.69747
R1341 VTAIL.n186 VTAIL.n136 9.69747
R1342 VTAIL.n166 VTAIL.n146 9.69747
R1343 VTAIL.n120 VTAIL.n70 9.69747
R1344 VTAIL.n100 VTAIL.n80 9.69747
R1345 VTAIL.n258 VTAIL.n198 9.45567
R1346 VTAIL.n60 VTAIL.n0 9.45567
R1347 VTAIL.n192 VTAIL.n132 9.45567
R1348 VTAIL.n126 VTAIL.n66 9.45567
R1349 VTAIL.n243 VTAIL.n242 9.3005
R1350 VTAIL.n206 VTAIL.n205 9.3005
R1351 VTAIL.n249 VTAIL.n248 9.3005
R1352 VTAIL.n251 VTAIL.n250 9.3005
R1353 VTAIL.n202 VTAIL.n201 9.3005
R1354 VTAIL.n257 VTAIL.n256 9.3005
R1355 VTAIL.n259 VTAIL.n258 9.3005
R1356 VTAIL.n210 VTAIL.n209 9.3005
R1357 VTAIL.n235 VTAIL.n234 9.3005
R1358 VTAIL.n233 VTAIL.n232 9.3005
R1359 VTAIL.n214 VTAIL.n213 9.3005
R1360 VTAIL.n227 VTAIL.n226 9.3005
R1361 VTAIL.n225 VTAIL.n224 9.3005
R1362 VTAIL.n218 VTAIL.n217 9.3005
R1363 VTAIL.n241 VTAIL.n240 9.3005
R1364 VTAIL.n45 VTAIL.n44 9.3005
R1365 VTAIL.n8 VTAIL.n7 9.3005
R1366 VTAIL.n51 VTAIL.n50 9.3005
R1367 VTAIL.n53 VTAIL.n52 9.3005
R1368 VTAIL.n4 VTAIL.n3 9.3005
R1369 VTAIL.n59 VTAIL.n58 9.3005
R1370 VTAIL.n61 VTAIL.n60 9.3005
R1371 VTAIL.n12 VTAIL.n11 9.3005
R1372 VTAIL.n37 VTAIL.n36 9.3005
R1373 VTAIL.n35 VTAIL.n34 9.3005
R1374 VTAIL.n16 VTAIL.n15 9.3005
R1375 VTAIL.n29 VTAIL.n28 9.3005
R1376 VTAIL.n27 VTAIL.n26 9.3005
R1377 VTAIL.n20 VTAIL.n19 9.3005
R1378 VTAIL.n43 VTAIL.n42 9.3005
R1379 VTAIL.n193 VTAIL.n192 9.3005
R1380 VTAIL.n191 VTAIL.n190 9.3005
R1381 VTAIL.n136 VTAIL.n135 9.3005
R1382 VTAIL.n185 VTAIL.n184 9.3005
R1383 VTAIL.n183 VTAIL.n182 9.3005
R1384 VTAIL.n140 VTAIL.n139 9.3005
R1385 VTAIL.n177 VTAIL.n176 9.3005
R1386 VTAIL.n175 VTAIL.n174 9.3005
R1387 VTAIL.n144 VTAIL.n143 9.3005
R1388 VTAIL.n169 VTAIL.n168 9.3005
R1389 VTAIL.n167 VTAIL.n166 9.3005
R1390 VTAIL.n148 VTAIL.n147 9.3005
R1391 VTAIL.n161 VTAIL.n160 9.3005
R1392 VTAIL.n159 VTAIL.n158 9.3005
R1393 VTAIL.n152 VTAIL.n151 9.3005
R1394 VTAIL.n74 VTAIL.n73 9.3005
R1395 VTAIL.n117 VTAIL.n116 9.3005
R1396 VTAIL.n119 VTAIL.n118 9.3005
R1397 VTAIL.n70 VTAIL.n69 9.3005
R1398 VTAIL.n125 VTAIL.n124 9.3005
R1399 VTAIL.n127 VTAIL.n126 9.3005
R1400 VTAIL.n111 VTAIL.n110 9.3005
R1401 VTAIL.n109 VTAIL.n108 9.3005
R1402 VTAIL.n78 VTAIL.n77 9.3005
R1403 VTAIL.n103 VTAIL.n102 9.3005
R1404 VTAIL.n101 VTAIL.n100 9.3005
R1405 VTAIL.n82 VTAIL.n81 9.3005
R1406 VTAIL.n95 VTAIL.n94 9.3005
R1407 VTAIL.n93 VTAIL.n92 9.3005
R1408 VTAIL.n86 VTAIL.n85 9.3005
R1409 VTAIL.n236 VTAIL.n235 8.92171
R1410 VTAIL.n251 VTAIL.n204 8.92171
R1411 VTAIL.n38 VTAIL.n37 8.92171
R1412 VTAIL.n53 VTAIL.n6 8.92171
R1413 VTAIL.n185 VTAIL.n138 8.92171
R1414 VTAIL.n170 VTAIL.n169 8.92171
R1415 VTAIL.n119 VTAIL.n72 8.92171
R1416 VTAIL.n104 VTAIL.n103 8.92171
R1417 VTAIL.n239 VTAIL.n210 8.14595
R1418 VTAIL.n248 VTAIL.n247 8.14595
R1419 VTAIL.n41 VTAIL.n12 8.14595
R1420 VTAIL.n50 VTAIL.n49 8.14595
R1421 VTAIL.n182 VTAIL.n181 8.14595
R1422 VTAIL.n173 VTAIL.n144 8.14595
R1423 VTAIL.n116 VTAIL.n115 8.14595
R1424 VTAIL.n107 VTAIL.n78 8.14595
R1425 VTAIL.n240 VTAIL.n208 7.3702
R1426 VTAIL.n244 VTAIL.n206 7.3702
R1427 VTAIL.n42 VTAIL.n10 7.3702
R1428 VTAIL.n46 VTAIL.n8 7.3702
R1429 VTAIL.n178 VTAIL.n140 7.3702
R1430 VTAIL.n174 VTAIL.n142 7.3702
R1431 VTAIL.n112 VTAIL.n74 7.3702
R1432 VTAIL.n108 VTAIL.n76 7.3702
R1433 VTAIL.n243 VTAIL.n208 6.59444
R1434 VTAIL.n244 VTAIL.n243 6.59444
R1435 VTAIL.n45 VTAIL.n10 6.59444
R1436 VTAIL.n46 VTAIL.n45 6.59444
R1437 VTAIL.n178 VTAIL.n177 6.59444
R1438 VTAIL.n177 VTAIL.n142 6.59444
R1439 VTAIL.n112 VTAIL.n111 6.59444
R1440 VTAIL.n111 VTAIL.n76 6.59444
R1441 VTAIL.n240 VTAIL.n239 5.81868
R1442 VTAIL.n247 VTAIL.n206 5.81868
R1443 VTAIL.n42 VTAIL.n41 5.81868
R1444 VTAIL.n49 VTAIL.n8 5.81868
R1445 VTAIL.n181 VTAIL.n140 5.81868
R1446 VTAIL.n174 VTAIL.n173 5.81868
R1447 VTAIL.n115 VTAIL.n74 5.81868
R1448 VTAIL.n108 VTAIL.n107 5.81868
R1449 VTAIL.n236 VTAIL.n210 5.04292
R1450 VTAIL.n248 VTAIL.n204 5.04292
R1451 VTAIL.n38 VTAIL.n12 5.04292
R1452 VTAIL.n50 VTAIL.n6 5.04292
R1453 VTAIL.n182 VTAIL.n138 5.04292
R1454 VTAIL.n170 VTAIL.n144 5.04292
R1455 VTAIL.n116 VTAIL.n72 5.04292
R1456 VTAIL.n104 VTAIL.n78 5.04292
R1457 VTAIL.n87 VTAIL.n85 4.38563
R1458 VTAIL.n219 VTAIL.n217 4.38563
R1459 VTAIL.n21 VTAIL.n19 4.38563
R1460 VTAIL.n153 VTAIL.n151 4.38563
R1461 VTAIL.n235 VTAIL.n212 4.26717
R1462 VTAIL.n252 VTAIL.n251 4.26717
R1463 VTAIL.n37 VTAIL.n14 4.26717
R1464 VTAIL.n54 VTAIL.n53 4.26717
R1465 VTAIL.n186 VTAIL.n185 4.26717
R1466 VTAIL.n169 VTAIL.n146 4.26717
R1467 VTAIL.n120 VTAIL.n119 4.26717
R1468 VTAIL.n103 VTAIL.n80 4.26717
R1469 VTAIL.n232 VTAIL.n231 3.49141
R1470 VTAIL.n255 VTAIL.n202 3.49141
R1471 VTAIL.n34 VTAIL.n33 3.49141
R1472 VTAIL.n57 VTAIL.n4 3.49141
R1473 VTAIL.n189 VTAIL.n136 3.49141
R1474 VTAIL.n166 VTAIL.n165 3.49141
R1475 VTAIL.n123 VTAIL.n70 3.49141
R1476 VTAIL.n100 VTAIL.n99 3.49141
R1477 VTAIL.n228 VTAIL.n214 2.71565
R1478 VTAIL.n256 VTAIL.n200 2.71565
R1479 VTAIL.n30 VTAIL.n16 2.71565
R1480 VTAIL.n58 VTAIL.n2 2.71565
R1481 VTAIL.n190 VTAIL.n134 2.71565
R1482 VTAIL.n162 VTAIL.n148 2.71565
R1483 VTAIL.n124 VTAIL.n68 2.71565
R1484 VTAIL.n96 VTAIL.n82 2.71565
R1485 VTAIL.n227 VTAIL.n216 1.93989
R1486 VTAIL.n260 VTAIL.n259 1.93989
R1487 VTAIL.n29 VTAIL.n18 1.93989
R1488 VTAIL.n62 VTAIL.n61 1.93989
R1489 VTAIL.n194 VTAIL.n193 1.93989
R1490 VTAIL.n161 VTAIL.n150 1.93989
R1491 VTAIL.n128 VTAIL.n127 1.93989
R1492 VTAIL.n95 VTAIL.n84 1.93989
R1493 VTAIL.n197 VTAIL.n131 1.4186
R1494 VTAIL.n224 VTAIL.n223 1.16414
R1495 VTAIL.n262 VTAIL.n198 1.16414
R1496 VTAIL.n26 VTAIL.n25 1.16414
R1497 VTAIL.n64 VTAIL.n0 1.16414
R1498 VTAIL.n196 VTAIL.n132 1.16414
R1499 VTAIL.n158 VTAIL.n157 1.16414
R1500 VTAIL.n130 VTAIL.n66 1.16414
R1501 VTAIL.n92 VTAIL.n91 1.16414
R1502 VTAIL VTAIL.n65 1.00266
R1503 VTAIL VTAIL.n263 0.416448
R1504 VTAIL.n220 VTAIL.n218 0.388379
R1505 VTAIL.n22 VTAIL.n20 0.388379
R1506 VTAIL.n154 VTAIL.n152 0.388379
R1507 VTAIL.n88 VTAIL.n86 0.388379
R1508 VTAIL.n225 VTAIL.n217 0.155672
R1509 VTAIL.n226 VTAIL.n225 0.155672
R1510 VTAIL.n226 VTAIL.n213 0.155672
R1511 VTAIL.n233 VTAIL.n213 0.155672
R1512 VTAIL.n234 VTAIL.n233 0.155672
R1513 VTAIL.n234 VTAIL.n209 0.155672
R1514 VTAIL.n241 VTAIL.n209 0.155672
R1515 VTAIL.n242 VTAIL.n241 0.155672
R1516 VTAIL.n242 VTAIL.n205 0.155672
R1517 VTAIL.n249 VTAIL.n205 0.155672
R1518 VTAIL.n250 VTAIL.n249 0.155672
R1519 VTAIL.n250 VTAIL.n201 0.155672
R1520 VTAIL.n257 VTAIL.n201 0.155672
R1521 VTAIL.n258 VTAIL.n257 0.155672
R1522 VTAIL.n27 VTAIL.n19 0.155672
R1523 VTAIL.n28 VTAIL.n27 0.155672
R1524 VTAIL.n28 VTAIL.n15 0.155672
R1525 VTAIL.n35 VTAIL.n15 0.155672
R1526 VTAIL.n36 VTAIL.n35 0.155672
R1527 VTAIL.n36 VTAIL.n11 0.155672
R1528 VTAIL.n43 VTAIL.n11 0.155672
R1529 VTAIL.n44 VTAIL.n43 0.155672
R1530 VTAIL.n44 VTAIL.n7 0.155672
R1531 VTAIL.n51 VTAIL.n7 0.155672
R1532 VTAIL.n52 VTAIL.n51 0.155672
R1533 VTAIL.n52 VTAIL.n3 0.155672
R1534 VTAIL.n59 VTAIL.n3 0.155672
R1535 VTAIL.n60 VTAIL.n59 0.155672
R1536 VTAIL.n192 VTAIL.n191 0.155672
R1537 VTAIL.n191 VTAIL.n135 0.155672
R1538 VTAIL.n184 VTAIL.n135 0.155672
R1539 VTAIL.n184 VTAIL.n183 0.155672
R1540 VTAIL.n183 VTAIL.n139 0.155672
R1541 VTAIL.n176 VTAIL.n139 0.155672
R1542 VTAIL.n176 VTAIL.n175 0.155672
R1543 VTAIL.n175 VTAIL.n143 0.155672
R1544 VTAIL.n168 VTAIL.n143 0.155672
R1545 VTAIL.n168 VTAIL.n167 0.155672
R1546 VTAIL.n167 VTAIL.n147 0.155672
R1547 VTAIL.n160 VTAIL.n147 0.155672
R1548 VTAIL.n160 VTAIL.n159 0.155672
R1549 VTAIL.n159 VTAIL.n151 0.155672
R1550 VTAIL.n126 VTAIL.n125 0.155672
R1551 VTAIL.n125 VTAIL.n69 0.155672
R1552 VTAIL.n118 VTAIL.n69 0.155672
R1553 VTAIL.n118 VTAIL.n117 0.155672
R1554 VTAIL.n117 VTAIL.n73 0.155672
R1555 VTAIL.n110 VTAIL.n73 0.155672
R1556 VTAIL.n110 VTAIL.n109 0.155672
R1557 VTAIL.n109 VTAIL.n77 0.155672
R1558 VTAIL.n102 VTAIL.n77 0.155672
R1559 VTAIL.n102 VTAIL.n101 0.155672
R1560 VTAIL.n101 VTAIL.n81 0.155672
R1561 VTAIL.n94 VTAIL.n81 0.155672
R1562 VTAIL.n94 VTAIL.n93 0.155672
R1563 VTAIL.n93 VTAIL.n85 0.155672
R1564 VDD2.n129 VDD2.n128 289.615
R1565 VDD2.n64 VDD2.n63 289.615
R1566 VDD2.n128 VDD2.n127 185
R1567 VDD2.n67 VDD2.n66 185
R1568 VDD2.n122 VDD2.n121 185
R1569 VDD2.n120 VDD2.n119 185
R1570 VDD2.n71 VDD2.n70 185
R1571 VDD2.n114 VDD2.n113 185
R1572 VDD2.n112 VDD2.n111 185
R1573 VDD2.n75 VDD2.n74 185
R1574 VDD2.n106 VDD2.n105 185
R1575 VDD2.n104 VDD2.n103 185
R1576 VDD2.n79 VDD2.n78 185
R1577 VDD2.n98 VDD2.n97 185
R1578 VDD2.n96 VDD2.n95 185
R1579 VDD2.n83 VDD2.n82 185
R1580 VDD2.n90 VDD2.n89 185
R1581 VDD2.n88 VDD2.n87 185
R1582 VDD2.n23 VDD2.n22 185
R1583 VDD2.n25 VDD2.n24 185
R1584 VDD2.n18 VDD2.n17 185
R1585 VDD2.n31 VDD2.n30 185
R1586 VDD2.n33 VDD2.n32 185
R1587 VDD2.n14 VDD2.n13 185
R1588 VDD2.n39 VDD2.n38 185
R1589 VDD2.n41 VDD2.n40 185
R1590 VDD2.n10 VDD2.n9 185
R1591 VDD2.n47 VDD2.n46 185
R1592 VDD2.n49 VDD2.n48 185
R1593 VDD2.n6 VDD2.n5 185
R1594 VDD2.n55 VDD2.n54 185
R1595 VDD2.n57 VDD2.n56 185
R1596 VDD2.n2 VDD2.n1 185
R1597 VDD2.n63 VDD2.n62 185
R1598 VDD2.n86 VDD2.t0 147.659
R1599 VDD2.n21 VDD2.t1 147.659
R1600 VDD2.n128 VDD2.n66 104.615
R1601 VDD2.n121 VDD2.n66 104.615
R1602 VDD2.n121 VDD2.n120 104.615
R1603 VDD2.n120 VDD2.n70 104.615
R1604 VDD2.n113 VDD2.n70 104.615
R1605 VDD2.n113 VDD2.n112 104.615
R1606 VDD2.n112 VDD2.n74 104.615
R1607 VDD2.n105 VDD2.n74 104.615
R1608 VDD2.n105 VDD2.n104 104.615
R1609 VDD2.n104 VDD2.n78 104.615
R1610 VDD2.n97 VDD2.n78 104.615
R1611 VDD2.n97 VDD2.n96 104.615
R1612 VDD2.n96 VDD2.n82 104.615
R1613 VDD2.n89 VDD2.n82 104.615
R1614 VDD2.n89 VDD2.n88 104.615
R1615 VDD2.n24 VDD2.n23 104.615
R1616 VDD2.n24 VDD2.n17 104.615
R1617 VDD2.n31 VDD2.n17 104.615
R1618 VDD2.n32 VDD2.n31 104.615
R1619 VDD2.n32 VDD2.n13 104.615
R1620 VDD2.n39 VDD2.n13 104.615
R1621 VDD2.n40 VDD2.n39 104.615
R1622 VDD2.n40 VDD2.n9 104.615
R1623 VDD2.n47 VDD2.n9 104.615
R1624 VDD2.n48 VDD2.n47 104.615
R1625 VDD2.n48 VDD2.n5 104.615
R1626 VDD2.n55 VDD2.n5 104.615
R1627 VDD2.n56 VDD2.n55 104.615
R1628 VDD2.n56 VDD2.n1 104.615
R1629 VDD2.n63 VDD2.n1 104.615
R1630 VDD2.n130 VDD2.n64 89.3422
R1631 VDD2.n88 VDD2.t0 52.3082
R1632 VDD2.n23 VDD2.t1 52.3082
R1633 VDD2.n130 VDD2.n129 51.5793
R1634 VDD2.n87 VDD2.n86 15.6677
R1635 VDD2.n22 VDD2.n21 15.6677
R1636 VDD2.n90 VDD2.n85 12.8005
R1637 VDD2.n25 VDD2.n20 12.8005
R1638 VDD2.n127 VDD2.n65 12.0247
R1639 VDD2.n91 VDD2.n83 12.0247
R1640 VDD2.n26 VDD2.n18 12.0247
R1641 VDD2.n62 VDD2.n0 12.0247
R1642 VDD2.n126 VDD2.n67 11.249
R1643 VDD2.n95 VDD2.n94 11.249
R1644 VDD2.n30 VDD2.n29 11.249
R1645 VDD2.n61 VDD2.n2 11.249
R1646 VDD2.n123 VDD2.n122 10.4732
R1647 VDD2.n98 VDD2.n81 10.4732
R1648 VDD2.n33 VDD2.n16 10.4732
R1649 VDD2.n58 VDD2.n57 10.4732
R1650 VDD2.n119 VDD2.n69 9.69747
R1651 VDD2.n99 VDD2.n79 9.69747
R1652 VDD2.n34 VDD2.n14 9.69747
R1653 VDD2.n54 VDD2.n4 9.69747
R1654 VDD2.n125 VDD2.n65 9.45567
R1655 VDD2.n60 VDD2.n0 9.45567
R1656 VDD2.n126 VDD2.n125 9.3005
R1657 VDD2.n124 VDD2.n123 9.3005
R1658 VDD2.n69 VDD2.n68 9.3005
R1659 VDD2.n118 VDD2.n117 9.3005
R1660 VDD2.n116 VDD2.n115 9.3005
R1661 VDD2.n73 VDD2.n72 9.3005
R1662 VDD2.n110 VDD2.n109 9.3005
R1663 VDD2.n108 VDD2.n107 9.3005
R1664 VDD2.n77 VDD2.n76 9.3005
R1665 VDD2.n102 VDD2.n101 9.3005
R1666 VDD2.n100 VDD2.n99 9.3005
R1667 VDD2.n81 VDD2.n80 9.3005
R1668 VDD2.n94 VDD2.n93 9.3005
R1669 VDD2.n92 VDD2.n91 9.3005
R1670 VDD2.n85 VDD2.n84 9.3005
R1671 VDD2.n45 VDD2.n44 9.3005
R1672 VDD2.n8 VDD2.n7 9.3005
R1673 VDD2.n51 VDD2.n50 9.3005
R1674 VDD2.n53 VDD2.n52 9.3005
R1675 VDD2.n4 VDD2.n3 9.3005
R1676 VDD2.n59 VDD2.n58 9.3005
R1677 VDD2.n61 VDD2.n60 9.3005
R1678 VDD2.n12 VDD2.n11 9.3005
R1679 VDD2.n37 VDD2.n36 9.3005
R1680 VDD2.n35 VDD2.n34 9.3005
R1681 VDD2.n16 VDD2.n15 9.3005
R1682 VDD2.n29 VDD2.n28 9.3005
R1683 VDD2.n27 VDD2.n26 9.3005
R1684 VDD2.n20 VDD2.n19 9.3005
R1685 VDD2.n43 VDD2.n42 9.3005
R1686 VDD2.n118 VDD2.n71 8.92171
R1687 VDD2.n103 VDD2.n102 8.92171
R1688 VDD2.n38 VDD2.n37 8.92171
R1689 VDD2.n53 VDD2.n6 8.92171
R1690 VDD2.n115 VDD2.n114 8.14595
R1691 VDD2.n106 VDD2.n77 8.14595
R1692 VDD2.n41 VDD2.n12 8.14595
R1693 VDD2.n50 VDD2.n49 8.14595
R1694 VDD2.n111 VDD2.n73 7.3702
R1695 VDD2.n107 VDD2.n75 7.3702
R1696 VDD2.n42 VDD2.n10 7.3702
R1697 VDD2.n46 VDD2.n8 7.3702
R1698 VDD2.n111 VDD2.n110 6.59444
R1699 VDD2.n110 VDD2.n75 6.59444
R1700 VDD2.n45 VDD2.n10 6.59444
R1701 VDD2.n46 VDD2.n45 6.59444
R1702 VDD2.n114 VDD2.n73 5.81868
R1703 VDD2.n107 VDD2.n106 5.81868
R1704 VDD2.n42 VDD2.n41 5.81868
R1705 VDD2.n49 VDD2.n8 5.81868
R1706 VDD2.n115 VDD2.n71 5.04292
R1707 VDD2.n103 VDD2.n77 5.04292
R1708 VDD2.n38 VDD2.n12 5.04292
R1709 VDD2.n50 VDD2.n6 5.04292
R1710 VDD2.n86 VDD2.n84 4.38563
R1711 VDD2.n21 VDD2.n19 4.38563
R1712 VDD2.n119 VDD2.n118 4.26717
R1713 VDD2.n102 VDD2.n79 4.26717
R1714 VDD2.n37 VDD2.n14 4.26717
R1715 VDD2.n54 VDD2.n53 4.26717
R1716 VDD2.n122 VDD2.n69 3.49141
R1717 VDD2.n99 VDD2.n98 3.49141
R1718 VDD2.n34 VDD2.n33 3.49141
R1719 VDD2.n57 VDD2.n4 3.49141
R1720 VDD2.n123 VDD2.n67 2.71565
R1721 VDD2.n95 VDD2.n81 2.71565
R1722 VDD2.n30 VDD2.n16 2.71565
R1723 VDD2.n58 VDD2.n2 2.71565
R1724 VDD2.n127 VDD2.n126 1.93989
R1725 VDD2.n94 VDD2.n83 1.93989
R1726 VDD2.n29 VDD2.n18 1.93989
R1727 VDD2.n62 VDD2.n61 1.93989
R1728 VDD2.n129 VDD2.n65 1.16414
R1729 VDD2.n91 VDD2.n90 1.16414
R1730 VDD2.n26 VDD2.n25 1.16414
R1731 VDD2.n64 VDD2.n0 1.16414
R1732 VDD2 VDD2.n130 0.532828
R1733 VDD2.n87 VDD2.n85 0.388379
R1734 VDD2.n22 VDD2.n20 0.388379
R1735 VDD2.n125 VDD2.n124 0.155672
R1736 VDD2.n124 VDD2.n68 0.155672
R1737 VDD2.n117 VDD2.n68 0.155672
R1738 VDD2.n117 VDD2.n116 0.155672
R1739 VDD2.n116 VDD2.n72 0.155672
R1740 VDD2.n109 VDD2.n72 0.155672
R1741 VDD2.n109 VDD2.n108 0.155672
R1742 VDD2.n108 VDD2.n76 0.155672
R1743 VDD2.n101 VDD2.n76 0.155672
R1744 VDD2.n101 VDD2.n100 0.155672
R1745 VDD2.n100 VDD2.n80 0.155672
R1746 VDD2.n93 VDD2.n80 0.155672
R1747 VDD2.n93 VDD2.n92 0.155672
R1748 VDD2.n92 VDD2.n84 0.155672
R1749 VDD2.n27 VDD2.n19 0.155672
R1750 VDD2.n28 VDD2.n27 0.155672
R1751 VDD2.n28 VDD2.n15 0.155672
R1752 VDD2.n35 VDD2.n15 0.155672
R1753 VDD2.n36 VDD2.n35 0.155672
R1754 VDD2.n36 VDD2.n11 0.155672
R1755 VDD2.n43 VDD2.n11 0.155672
R1756 VDD2.n44 VDD2.n43 0.155672
R1757 VDD2.n44 VDD2.n7 0.155672
R1758 VDD2.n51 VDD2.n7 0.155672
R1759 VDD2.n52 VDD2.n51 0.155672
R1760 VDD2.n52 VDD2.n3 0.155672
R1761 VDD2.n59 VDD2.n3 0.155672
R1762 VDD2.n60 VDD2.n59 0.155672
R1763 VP.n0 VP.t0 255.663
R1764 VP.n0 VP.t1 212.974
R1765 VP VP.n0 0.241678
R1766 VDD1.n64 VDD1.n63 289.615
R1767 VDD1.n129 VDD1.n128 289.615
R1768 VDD1.n63 VDD1.n62 185
R1769 VDD1.n2 VDD1.n1 185
R1770 VDD1.n57 VDD1.n56 185
R1771 VDD1.n55 VDD1.n54 185
R1772 VDD1.n6 VDD1.n5 185
R1773 VDD1.n49 VDD1.n48 185
R1774 VDD1.n47 VDD1.n46 185
R1775 VDD1.n10 VDD1.n9 185
R1776 VDD1.n41 VDD1.n40 185
R1777 VDD1.n39 VDD1.n38 185
R1778 VDD1.n14 VDD1.n13 185
R1779 VDD1.n33 VDD1.n32 185
R1780 VDD1.n31 VDD1.n30 185
R1781 VDD1.n18 VDD1.n17 185
R1782 VDD1.n25 VDD1.n24 185
R1783 VDD1.n23 VDD1.n22 185
R1784 VDD1.n88 VDD1.n87 185
R1785 VDD1.n90 VDD1.n89 185
R1786 VDD1.n83 VDD1.n82 185
R1787 VDD1.n96 VDD1.n95 185
R1788 VDD1.n98 VDD1.n97 185
R1789 VDD1.n79 VDD1.n78 185
R1790 VDD1.n104 VDD1.n103 185
R1791 VDD1.n106 VDD1.n105 185
R1792 VDD1.n75 VDD1.n74 185
R1793 VDD1.n112 VDD1.n111 185
R1794 VDD1.n114 VDD1.n113 185
R1795 VDD1.n71 VDD1.n70 185
R1796 VDD1.n120 VDD1.n119 185
R1797 VDD1.n122 VDD1.n121 185
R1798 VDD1.n67 VDD1.n66 185
R1799 VDD1.n128 VDD1.n127 185
R1800 VDD1.n21 VDD1.t1 147.659
R1801 VDD1.n86 VDD1.t0 147.659
R1802 VDD1.n63 VDD1.n1 104.615
R1803 VDD1.n56 VDD1.n1 104.615
R1804 VDD1.n56 VDD1.n55 104.615
R1805 VDD1.n55 VDD1.n5 104.615
R1806 VDD1.n48 VDD1.n5 104.615
R1807 VDD1.n48 VDD1.n47 104.615
R1808 VDD1.n47 VDD1.n9 104.615
R1809 VDD1.n40 VDD1.n9 104.615
R1810 VDD1.n40 VDD1.n39 104.615
R1811 VDD1.n39 VDD1.n13 104.615
R1812 VDD1.n32 VDD1.n13 104.615
R1813 VDD1.n32 VDD1.n31 104.615
R1814 VDD1.n31 VDD1.n17 104.615
R1815 VDD1.n24 VDD1.n17 104.615
R1816 VDD1.n24 VDD1.n23 104.615
R1817 VDD1.n89 VDD1.n88 104.615
R1818 VDD1.n89 VDD1.n82 104.615
R1819 VDD1.n96 VDD1.n82 104.615
R1820 VDD1.n97 VDD1.n96 104.615
R1821 VDD1.n97 VDD1.n78 104.615
R1822 VDD1.n104 VDD1.n78 104.615
R1823 VDD1.n105 VDD1.n104 104.615
R1824 VDD1.n105 VDD1.n74 104.615
R1825 VDD1.n112 VDD1.n74 104.615
R1826 VDD1.n113 VDD1.n112 104.615
R1827 VDD1.n113 VDD1.n70 104.615
R1828 VDD1.n120 VDD1.n70 104.615
R1829 VDD1.n121 VDD1.n120 104.615
R1830 VDD1.n121 VDD1.n66 104.615
R1831 VDD1.n128 VDD1.n66 104.615
R1832 VDD1 VDD1.n129 90.3411
R1833 VDD1.n23 VDD1.t1 52.3082
R1834 VDD1.n88 VDD1.t0 52.3082
R1835 VDD1 VDD1.n64 52.1116
R1836 VDD1.n22 VDD1.n21 15.6677
R1837 VDD1.n87 VDD1.n86 15.6677
R1838 VDD1.n25 VDD1.n20 12.8005
R1839 VDD1.n90 VDD1.n85 12.8005
R1840 VDD1.n62 VDD1.n0 12.0247
R1841 VDD1.n26 VDD1.n18 12.0247
R1842 VDD1.n91 VDD1.n83 12.0247
R1843 VDD1.n127 VDD1.n65 12.0247
R1844 VDD1.n61 VDD1.n2 11.249
R1845 VDD1.n30 VDD1.n29 11.249
R1846 VDD1.n95 VDD1.n94 11.249
R1847 VDD1.n126 VDD1.n67 11.249
R1848 VDD1.n58 VDD1.n57 10.4732
R1849 VDD1.n33 VDD1.n16 10.4732
R1850 VDD1.n98 VDD1.n81 10.4732
R1851 VDD1.n123 VDD1.n122 10.4732
R1852 VDD1.n54 VDD1.n4 9.69747
R1853 VDD1.n34 VDD1.n14 9.69747
R1854 VDD1.n99 VDD1.n79 9.69747
R1855 VDD1.n119 VDD1.n69 9.69747
R1856 VDD1.n60 VDD1.n0 9.45567
R1857 VDD1.n125 VDD1.n65 9.45567
R1858 VDD1.n61 VDD1.n60 9.3005
R1859 VDD1.n59 VDD1.n58 9.3005
R1860 VDD1.n4 VDD1.n3 9.3005
R1861 VDD1.n53 VDD1.n52 9.3005
R1862 VDD1.n51 VDD1.n50 9.3005
R1863 VDD1.n8 VDD1.n7 9.3005
R1864 VDD1.n45 VDD1.n44 9.3005
R1865 VDD1.n43 VDD1.n42 9.3005
R1866 VDD1.n12 VDD1.n11 9.3005
R1867 VDD1.n37 VDD1.n36 9.3005
R1868 VDD1.n35 VDD1.n34 9.3005
R1869 VDD1.n16 VDD1.n15 9.3005
R1870 VDD1.n29 VDD1.n28 9.3005
R1871 VDD1.n27 VDD1.n26 9.3005
R1872 VDD1.n20 VDD1.n19 9.3005
R1873 VDD1.n110 VDD1.n109 9.3005
R1874 VDD1.n73 VDD1.n72 9.3005
R1875 VDD1.n116 VDD1.n115 9.3005
R1876 VDD1.n118 VDD1.n117 9.3005
R1877 VDD1.n69 VDD1.n68 9.3005
R1878 VDD1.n124 VDD1.n123 9.3005
R1879 VDD1.n126 VDD1.n125 9.3005
R1880 VDD1.n77 VDD1.n76 9.3005
R1881 VDD1.n102 VDD1.n101 9.3005
R1882 VDD1.n100 VDD1.n99 9.3005
R1883 VDD1.n81 VDD1.n80 9.3005
R1884 VDD1.n94 VDD1.n93 9.3005
R1885 VDD1.n92 VDD1.n91 9.3005
R1886 VDD1.n85 VDD1.n84 9.3005
R1887 VDD1.n108 VDD1.n107 9.3005
R1888 VDD1.n53 VDD1.n6 8.92171
R1889 VDD1.n38 VDD1.n37 8.92171
R1890 VDD1.n103 VDD1.n102 8.92171
R1891 VDD1.n118 VDD1.n71 8.92171
R1892 VDD1.n50 VDD1.n49 8.14595
R1893 VDD1.n41 VDD1.n12 8.14595
R1894 VDD1.n106 VDD1.n77 8.14595
R1895 VDD1.n115 VDD1.n114 8.14595
R1896 VDD1.n46 VDD1.n8 7.3702
R1897 VDD1.n42 VDD1.n10 7.3702
R1898 VDD1.n107 VDD1.n75 7.3702
R1899 VDD1.n111 VDD1.n73 7.3702
R1900 VDD1.n46 VDD1.n45 6.59444
R1901 VDD1.n45 VDD1.n10 6.59444
R1902 VDD1.n110 VDD1.n75 6.59444
R1903 VDD1.n111 VDD1.n110 6.59444
R1904 VDD1.n49 VDD1.n8 5.81868
R1905 VDD1.n42 VDD1.n41 5.81868
R1906 VDD1.n107 VDD1.n106 5.81868
R1907 VDD1.n114 VDD1.n73 5.81868
R1908 VDD1.n50 VDD1.n6 5.04292
R1909 VDD1.n38 VDD1.n12 5.04292
R1910 VDD1.n103 VDD1.n77 5.04292
R1911 VDD1.n115 VDD1.n71 5.04292
R1912 VDD1.n21 VDD1.n19 4.38563
R1913 VDD1.n86 VDD1.n84 4.38563
R1914 VDD1.n54 VDD1.n53 4.26717
R1915 VDD1.n37 VDD1.n14 4.26717
R1916 VDD1.n102 VDD1.n79 4.26717
R1917 VDD1.n119 VDD1.n118 4.26717
R1918 VDD1.n57 VDD1.n4 3.49141
R1919 VDD1.n34 VDD1.n33 3.49141
R1920 VDD1.n99 VDD1.n98 3.49141
R1921 VDD1.n122 VDD1.n69 3.49141
R1922 VDD1.n58 VDD1.n2 2.71565
R1923 VDD1.n30 VDD1.n16 2.71565
R1924 VDD1.n95 VDD1.n81 2.71565
R1925 VDD1.n123 VDD1.n67 2.71565
R1926 VDD1.n62 VDD1.n61 1.93989
R1927 VDD1.n29 VDD1.n18 1.93989
R1928 VDD1.n94 VDD1.n83 1.93989
R1929 VDD1.n127 VDD1.n126 1.93989
R1930 VDD1.n64 VDD1.n0 1.16414
R1931 VDD1.n26 VDD1.n25 1.16414
R1932 VDD1.n91 VDD1.n90 1.16414
R1933 VDD1.n129 VDD1.n65 1.16414
R1934 VDD1.n22 VDD1.n20 0.388379
R1935 VDD1.n87 VDD1.n85 0.388379
R1936 VDD1.n60 VDD1.n59 0.155672
R1937 VDD1.n59 VDD1.n3 0.155672
R1938 VDD1.n52 VDD1.n3 0.155672
R1939 VDD1.n52 VDD1.n51 0.155672
R1940 VDD1.n51 VDD1.n7 0.155672
R1941 VDD1.n44 VDD1.n7 0.155672
R1942 VDD1.n44 VDD1.n43 0.155672
R1943 VDD1.n43 VDD1.n11 0.155672
R1944 VDD1.n36 VDD1.n11 0.155672
R1945 VDD1.n36 VDD1.n35 0.155672
R1946 VDD1.n35 VDD1.n15 0.155672
R1947 VDD1.n28 VDD1.n15 0.155672
R1948 VDD1.n28 VDD1.n27 0.155672
R1949 VDD1.n27 VDD1.n19 0.155672
R1950 VDD1.n92 VDD1.n84 0.155672
R1951 VDD1.n93 VDD1.n92 0.155672
R1952 VDD1.n93 VDD1.n80 0.155672
R1953 VDD1.n100 VDD1.n80 0.155672
R1954 VDD1.n101 VDD1.n100 0.155672
R1955 VDD1.n101 VDD1.n76 0.155672
R1956 VDD1.n108 VDD1.n76 0.155672
R1957 VDD1.n109 VDD1.n108 0.155672
R1958 VDD1.n109 VDD1.n72 0.155672
R1959 VDD1.n116 VDD1.n72 0.155672
R1960 VDD1.n117 VDD1.n116 0.155672
R1961 VDD1.n117 VDD1.n68 0.155672
R1962 VDD1.n124 VDD1.n68 0.155672
R1963 VDD1.n125 VDD1.n124 0.155672
C0 VN VP 5.10828f
C1 VP VTAIL 2.24307f
C2 VDD2 VDD1 0.588267f
C3 VN VDD1 0.147453f
C4 VTAIL VDD1 5.00944f
C5 VN VDD2 2.61472f
C6 VTAIL VDD2 5.05419f
C7 VP VDD1 2.7664f
C8 VN VTAIL 2.22871f
C9 VP VDD2 0.302127f
C10 VDD2 B 4.168139f
C11 VDD1 B 6.775219f
C12 VTAIL B 6.982545f
C13 VN B 9.97795f
C14 VP B 5.487463f
C15 VDD1.n0 B 0.01147f
C16 VDD1.n1 B 0.025839f
C17 VDD1.n2 B 0.011575f
C18 VDD1.n3 B 0.020344f
C19 VDD1.n4 B 0.010932f
C20 VDD1.n5 B 0.025839f
C21 VDD1.n6 B 0.011575f
C22 VDD1.n7 B 0.020344f
C23 VDD1.n8 B 0.010932f
C24 VDD1.n9 B 0.025839f
C25 VDD1.n10 B 0.011575f
C26 VDD1.n11 B 0.020344f
C27 VDD1.n12 B 0.010932f
C28 VDD1.n13 B 0.025839f
C29 VDD1.n14 B 0.011575f
C30 VDD1.n15 B 0.020344f
C31 VDD1.n16 B 0.010932f
C32 VDD1.n17 B 0.025839f
C33 VDD1.n18 B 0.011575f
C34 VDD1.n19 B 1.04017f
C35 VDD1.n20 B 0.010932f
C36 VDD1.t1 B 0.042394f
C37 VDD1.n21 B 0.117182f
C38 VDD1.n22 B 0.015264f
C39 VDD1.n23 B 0.019379f
C40 VDD1.n24 B 0.025839f
C41 VDD1.n25 B 0.011575f
C42 VDD1.n26 B 0.010932f
C43 VDD1.n27 B 0.020344f
C44 VDD1.n28 B 0.020344f
C45 VDD1.n29 B 0.010932f
C46 VDD1.n30 B 0.011575f
C47 VDD1.n31 B 0.025839f
C48 VDD1.n32 B 0.025839f
C49 VDD1.n33 B 0.011575f
C50 VDD1.n34 B 0.010932f
C51 VDD1.n35 B 0.020344f
C52 VDD1.n36 B 0.020344f
C53 VDD1.n37 B 0.010932f
C54 VDD1.n38 B 0.011575f
C55 VDD1.n39 B 0.025839f
C56 VDD1.n40 B 0.025839f
C57 VDD1.n41 B 0.011575f
C58 VDD1.n42 B 0.010932f
C59 VDD1.n43 B 0.020344f
C60 VDD1.n44 B 0.020344f
C61 VDD1.n45 B 0.010932f
C62 VDD1.n46 B 0.011575f
C63 VDD1.n47 B 0.025839f
C64 VDD1.n48 B 0.025839f
C65 VDD1.n49 B 0.011575f
C66 VDD1.n50 B 0.010932f
C67 VDD1.n51 B 0.020344f
C68 VDD1.n52 B 0.020344f
C69 VDD1.n53 B 0.010932f
C70 VDD1.n54 B 0.011575f
C71 VDD1.n55 B 0.025839f
C72 VDD1.n56 B 0.025839f
C73 VDD1.n57 B 0.011575f
C74 VDD1.n58 B 0.010932f
C75 VDD1.n59 B 0.020344f
C76 VDD1.n60 B 0.052583f
C77 VDD1.n61 B 0.010932f
C78 VDD1.n62 B 0.011575f
C79 VDD1.n63 B 0.052054f
C80 VDD1.n64 B 0.058919f
C81 VDD1.n65 B 0.01147f
C82 VDD1.n66 B 0.025839f
C83 VDD1.n67 B 0.011575f
C84 VDD1.n68 B 0.020344f
C85 VDD1.n69 B 0.010932f
C86 VDD1.n70 B 0.025839f
C87 VDD1.n71 B 0.011575f
C88 VDD1.n72 B 0.020344f
C89 VDD1.n73 B 0.010932f
C90 VDD1.n74 B 0.025839f
C91 VDD1.n75 B 0.011575f
C92 VDD1.n76 B 0.020344f
C93 VDD1.n77 B 0.010932f
C94 VDD1.n78 B 0.025839f
C95 VDD1.n79 B 0.011575f
C96 VDD1.n80 B 0.020344f
C97 VDD1.n81 B 0.010932f
C98 VDD1.n82 B 0.025839f
C99 VDD1.n83 B 0.011575f
C100 VDD1.n84 B 1.04017f
C101 VDD1.n85 B 0.010932f
C102 VDD1.t0 B 0.042394f
C103 VDD1.n86 B 0.117182f
C104 VDD1.n87 B 0.015264f
C105 VDD1.n88 B 0.019379f
C106 VDD1.n89 B 0.025839f
C107 VDD1.n90 B 0.011575f
C108 VDD1.n91 B 0.010932f
C109 VDD1.n92 B 0.020344f
C110 VDD1.n93 B 0.020344f
C111 VDD1.n94 B 0.010932f
C112 VDD1.n95 B 0.011575f
C113 VDD1.n96 B 0.025839f
C114 VDD1.n97 B 0.025839f
C115 VDD1.n98 B 0.011575f
C116 VDD1.n99 B 0.010932f
C117 VDD1.n100 B 0.020344f
C118 VDD1.n101 B 0.020344f
C119 VDD1.n102 B 0.010932f
C120 VDD1.n103 B 0.011575f
C121 VDD1.n104 B 0.025839f
C122 VDD1.n105 B 0.025839f
C123 VDD1.n106 B 0.011575f
C124 VDD1.n107 B 0.010932f
C125 VDD1.n108 B 0.020344f
C126 VDD1.n109 B 0.020344f
C127 VDD1.n110 B 0.010932f
C128 VDD1.n111 B 0.011575f
C129 VDD1.n112 B 0.025839f
C130 VDD1.n113 B 0.025839f
C131 VDD1.n114 B 0.011575f
C132 VDD1.n115 B 0.010932f
C133 VDD1.n116 B 0.020344f
C134 VDD1.n117 B 0.020344f
C135 VDD1.n118 B 0.010932f
C136 VDD1.n119 B 0.011575f
C137 VDD1.n120 B 0.025839f
C138 VDD1.n121 B 0.025839f
C139 VDD1.n122 B 0.011575f
C140 VDD1.n123 B 0.010932f
C141 VDD1.n124 B 0.020344f
C142 VDD1.n125 B 0.052583f
C143 VDD1.n126 B 0.010932f
C144 VDD1.n127 B 0.011575f
C145 VDD1.n128 B 0.052054f
C146 VDD1.n129 B 0.590517f
C147 VP.t0 B 3.00151f
C148 VP.t1 B 2.59407f
C149 VP.n0 B 4.44458f
C150 VDD2.n0 B 0.011433f
C151 VDD2.n1 B 0.025756f
C152 VDD2.n2 B 0.011538f
C153 VDD2.n3 B 0.020279f
C154 VDD2.n4 B 0.010897f
C155 VDD2.n5 B 0.025756f
C156 VDD2.n6 B 0.011538f
C157 VDD2.n7 B 0.020279f
C158 VDD2.n8 B 0.010897f
C159 VDD2.n9 B 0.025756f
C160 VDD2.n10 B 0.011538f
C161 VDD2.n11 B 0.020279f
C162 VDD2.n12 B 0.010897f
C163 VDD2.n13 B 0.025756f
C164 VDD2.n14 B 0.011538f
C165 VDD2.n15 B 0.020279f
C166 VDD2.n16 B 0.010897f
C167 VDD2.n17 B 0.025756f
C168 VDD2.n18 B 0.011538f
C169 VDD2.n19 B 1.03682f
C170 VDD2.n20 B 0.010897f
C171 VDD2.t1 B 0.042257f
C172 VDD2.n21 B 0.116805f
C173 VDD2.n22 B 0.015215f
C174 VDD2.n23 B 0.019317f
C175 VDD2.n24 B 0.025756f
C176 VDD2.n25 B 0.011538f
C177 VDD2.n26 B 0.010897f
C178 VDD2.n27 B 0.020279f
C179 VDD2.n28 B 0.020279f
C180 VDD2.n29 B 0.010897f
C181 VDD2.n30 B 0.011538f
C182 VDD2.n31 B 0.025756f
C183 VDD2.n32 B 0.025756f
C184 VDD2.n33 B 0.011538f
C185 VDD2.n34 B 0.010897f
C186 VDD2.n35 B 0.020279f
C187 VDD2.n36 B 0.020279f
C188 VDD2.n37 B 0.010897f
C189 VDD2.n38 B 0.011538f
C190 VDD2.n39 B 0.025756f
C191 VDD2.n40 B 0.025756f
C192 VDD2.n41 B 0.011538f
C193 VDD2.n42 B 0.010897f
C194 VDD2.n43 B 0.020279f
C195 VDD2.n44 B 0.020279f
C196 VDD2.n45 B 0.010897f
C197 VDD2.n46 B 0.011538f
C198 VDD2.n47 B 0.025756f
C199 VDD2.n48 B 0.025756f
C200 VDD2.n49 B 0.011538f
C201 VDD2.n50 B 0.010897f
C202 VDD2.n51 B 0.020279f
C203 VDD2.n52 B 0.020279f
C204 VDD2.n53 B 0.010897f
C205 VDD2.n54 B 0.011538f
C206 VDD2.n55 B 0.025756f
C207 VDD2.n56 B 0.025756f
C208 VDD2.n57 B 0.011538f
C209 VDD2.n58 B 0.010897f
C210 VDD2.n59 B 0.020279f
C211 VDD2.n60 B 0.052413f
C212 VDD2.n61 B 0.010897f
C213 VDD2.n62 B 0.011538f
C214 VDD2.n63 B 0.051886f
C215 VDD2.n64 B 0.554804f
C216 VDD2.n65 B 0.011433f
C217 VDD2.n66 B 0.025756f
C218 VDD2.n67 B 0.011538f
C219 VDD2.n68 B 0.020279f
C220 VDD2.n69 B 0.010897f
C221 VDD2.n70 B 0.025756f
C222 VDD2.n71 B 0.011538f
C223 VDD2.n72 B 0.020279f
C224 VDD2.n73 B 0.010897f
C225 VDD2.n74 B 0.025756f
C226 VDD2.n75 B 0.011538f
C227 VDD2.n76 B 0.020279f
C228 VDD2.n77 B 0.010897f
C229 VDD2.n78 B 0.025756f
C230 VDD2.n79 B 0.011538f
C231 VDD2.n80 B 0.020279f
C232 VDD2.n81 B 0.010897f
C233 VDD2.n82 B 0.025756f
C234 VDD2.n83 B 0.011538f
C235 VDD2.n84 B 1.03682f
C236 VDD2.n85 B 0.010897f
C237 VDD2.t0 B 0.042257f
C238 VDD2.n86 B 0.116805f
C239 VDD2.n87 B 0.015215f
C240 VDD2.n88 B 0.019317f
C241 VDD2.n89 B 0.025756f
C242 VDD2.n90 B 0.011538f
C243 VDD2.n91 B 0.010897f
C244 VDD2.n92 B 0.020279f
C245 VDD2.n93 B 0.020279f
C246 VDD2.n94 B 0.010897f
C247 VDD2.n95 B 0.011538f
C248 VDD2.n96 B 0.025756f
C249 VDD2.n97 B 0.025756f
C250 VDD2.n98 B 0.011538f
C251 VDD2.n99 B 0.010897f
C252 VDD2.n100 B 0.020279f
C253 VDD2.n101 B 0.020279f
C254 VDD2.n102 B 0.010897f
C255 VDD2.n103 B 0.011538f
C256 VDD2.n104 B 0.025756f
C257 VDD2.n105 B 0.025756f
C258 VDD2.n106 B 0.011538f
C259 VDD2.n107 B 0.010897f
C260 VDD2.n108 B 0.020279f
C261 VDD2.n109 B 0.020279f
C262 VDD2.n110 B 0.010897f
C263 VDD2.n111 B 0.011538f
C264 VDD2.n112 B 0.025756f
C265 VDD2.n113 B 0.025756f
C266 VDD2.n114 B 0.011538f
C267 VDD2.n115 B 0.010897f
C268 VDD2.n116 B 0.020279f
C269 VDD2.n117 B 0.020279f
C270 VDD2.n118 B 0.010897f
C271 VDD2.n119 B 0.011538f
C272 VDD2.n120 B 0.025756f
C273 VDD2.n121 B 0.025756f
C274 VDD2.n122 B 0.011538f
C275 VDD2.n123 B 0.010897f
C276 VDD2.n124 B 0.020279f
C277 VDD2.n125 B 0.052413f
C278 VDD2.n126 B 0.010897f
C279 VDD2.n127 B 0.011538f
C280 VDD2.n128 B 0.051886f
C281 VDD2.n129 B 0.057953f
C282 VDD2.n130 B 2.37619f
C283 VTAIL.n0 B 0.011518f
C284 VTAIL.n1 B 0.025949f
C285 VTAIL.n2 B 0.011624f
C286 VTAIL.n3 B 0.02043f
C287 VTAIL.n4 B 0.010978f
C288 VTAIL.n5 B 0.025949f
C289 VTAIL.n6 B 0.011624f
C290 VTAIL.n7 B 0.02043f
C291 VTAIL.n8 B 0.010978f
C292 VTAIL.n9 B 0.025949f
C293 VTAIL.n10 B 0.011624f
C294 VTAIL.n11 B 0.02043f
C295 VTAIL.n12 B 0.010978f
C296 VTAIL.n13 B 0.025949f
C297 VTAIL.n14 B 0.011624f
C298 VTAIL.n15 B 0.02043f
C299 VTAIL.n16 B 0.010978f
C300 VTAIL.n17 B 0.025949f
C301 VTAIL.n18 B 0.011624f
C302 VTAIL.n19 B 1.04458f
C303 VTAIL.n20 B 0.010978f
C304 VTAIL.t1 B 0.042574f
C305 VTAIL.n21 B 0.117679f
C306 VTAIL.n22 B 0.015329f
C307 VTAIL.n23 B 0.019462f
C308 VTAIL.n24 B 0.025949f
C309 VTAIL.n25 B 0.011624f
C310 VTAIL.n26 B 0.010978f
C311 VTAIL.n27 B 0.02043f
C312 VTAIL.n28 B 0.02043f
C313 VTAIL.n29 B 0.010978f
C314 VTAIL.n30 B 0.011624f
C315 VTAIL.n31 B 0.025949f
C316 VTAIL.n32 B 0.025949f
C317 VTAIL.n33 B 0.011624f
C318 VTAIL.n34 B 0.010978f
C319 VTAIL.n35 B 0.02043f
C320 VTAIL.n36 B 0.02043f
C321 VTAIL.n37 B 0.010978f
C322 VTAIL.n38 B 0.011624f
C323 VTAIL.n39 B 0.025949f
C324 VTAIL.n40 B 0.025949f
C325 VTAIL.n41 B 0.011624f
C326 VTAIL.n42 B 0.010978f
C327 VTAIL.n43 B 0.02043f
C328 VTAIL.n44 B 0.02043f
C329 VTAIL.n45 B 0.010978f
C330 VTAIL.n46 B 0.011624f
C331 VTAIL.n47 B 0.025949f
C332 VTAIL.n48 B 0.025949f
C333 VTAIL.n49 B 0.011624f
C334 VTAIL.n50 B 0.010978f
C335 VTAIL.n51 B 0.02043f
C336 VTAIL.n52 B 0.02043f
C337 VTAIL.n53 B 0.010978f
C338 VTAIL.n54 B 0.011624f
C339 VTAIL.n55 B 0.025949f
C340 VTAIL.n56 B 0.025949f
C341 VTAIL.n57 B 0.011624f
C342 VTAIL.n58 B 0.010978f
C343 VTAIL.n59 B 0.02043f
C344 VTAIL.n60 B 0.052806f
C345 VTAIL.n61 B 0.010978f
C346 VTAIL.n62 B 0.011624f
C347 VTAIL.n63 B 0.052275f
C348 VTAIL.n64 B 0.044308f
C349 VTAIL.n65 B 1.2916f
C350 VTAIL.n66 B 0.011518f
C351 VTAIL.n67 B 0.025949f
C352 VTAIL.n68 B 0.011624f
C353 VTAIL.n69 B 0.02043f
C354 VTAIL.n70 B 0.010978f
C355 VTAIL.n71 B 0.025949f
C356 VTAIL.n72 B 0.011624f
C357 VTAIL.n73 B 0.02043f
C358 VTAIL.n74 B 0.010978f
C359 VTAIL.n75 B 0.025949f
C360 VTAIL.n76 B 0.011624f
C361 VTAIL.n77 B 0.02043f
C362 VTAIL.n78 B 0.010978f
C363 VTAIL.n79 B 0.025949f
C364 VTAIL.n80 B 0.011624f
C365 VTAIL.n81 B 0.02043f
C366 VTAIL.n82 B 0.010978f
C367 VTAIL.n83 B 0.025949f
C368 VTAIL.n84 B 0.011624f
C369 VTAIL.n85 B 1.04458f
C370 VTAIL.n86 B 0.010978f
C371 VTAIL.t2 B 0.042574f
C372 VTAIL.n87 B 0.117679f
C373 VTAIL.n88 B 0.015329f
C374 VTAIL.n89 B 0.019462f
C375 VTAIL.n90 B 0.025949f
C376 VTAIL.n91 B 0.011624f
C377 VTAIL.n92 B 0.010978f
C378 VTAIL.n93 B 0.02043f
C379 VTAIL.n94 B 0.02043f
C380 VTAIL.n95 B 0.010978f
C381 VTAIL.n96 B 0.011624f
C382 VTAIL.n97 B 0.025949f
C383 VTAIL.n98 B 0.025949f
C384 VTAIL.n99 B 0.011624f
C385 VTAIL.n100 B 0.010978f
C386 VTAIL.n101 B 0.02043f
C387 VTAIL.n102 B 0.02043f
C388 VTAIL.n103 B 0.010978f
C389 VTAIL.n104 B 0.011624f
C390 VTAIL.n105 B 0.025949f
C391 VTAIL.n106 B 0.025949f
C392 VTAIL.n107 B 0.011624f
C393 VTAIL.n108 B 0.010978f
C394 VTAIL.n109 B 0.02043f
C395 VTAIL.n110 B 0.02043f
C396 VTAIL.n111 B 0.010978f
C397 VTAIL.n112 B 0.011624f
C398 VTAIL.n113 B 0.025949f
C399 VTAIL.n114 B 0.025949f
C400 VTAIL.n115 B 0.011624f
C401 VTAIL.n116 B 0.010978f
C402 VTAIL.n117 B 0.02043f
C403 VTAIL.n118 B 0.02043f
C404 VTAIL.n119 B 0.010978f
C405 VTAIL.n120 B 0.011624f
C406 VTAIL.n121 B 0.025949f
C407 VTAIL.n122 B 0.025949f
C408 VTAIL.n123 B 0.011624f
C409 VTAIL.n124 B 0.010978f
C410 VTAIL.n125 B 0.02043f
C411 VTAIL.n126 B 0.052806f
C412 VTAIL.n127 B 0.010978f
C413 VTAIL.n128 B 0.011624f
C414 VTAIL.n129 B 0.052275f
C415 VTAIL.n130 B 0.044308f
C416 VTAIL.n131 B 1.31898f
C417 VTAIL.n132 B 0.011518f
C418 VTAIL.n133 B 0.025949f
C419 VTAIL.n134 B 0.011624f
C420 VTAIL.n135 B 0.02043f
C421 VTAIL.n136 B 0.010978f
C422 VTAIL.n137 B 0.025949f
C423 VTAIL.n138 B 0.011624f
C424 VTAIL.n139 B 0.02043f
C425 VTAIL.n140 B 0.010978f
C426 VTAIL.n141 B 0.025949f
C427 VTAIL.n142 B 0.011624f
C428 VTAIL.n143 B 0.02043f
C429 VTAIL.n144 B 0.010978f
C430 VTAIL.n145 B 0.025949f
C431 VTAIL.n146 B 0.011624f
C432 VTAIL.n147 B 0.02043f
C433 VTAIL.n148 B 0.010978f
C434 VTAIL.n149 B 0.025949f
C435 VTAIL.n150 B 0.011624f
C436 VTAIL.n151 B 1.04458f
C437 VTAIL.n152 B 0.010978f
C438 VTAIL.t0 B 0.042574f
C439 VTAIL.n153 B 0.117679f
C440 VTAIL.n154 B 0.015329f
C441 VTAIL.n155 B 0.019462f
C442 VTAIL.n156 B 0.025949f
C443 VTAIL.n157 B 0.011624f
C444 VTAIL.n158 B 0.010978f
C445 VTAIL.n159 B 0.02043f
C446 VTAIL.n160 B 0.02043f
C447 VTAIL.n161 B 0.010978f
C448 VTAIL.n162 B 0.011624f
C449 VTAIL.n163 B 0.025949f
C450 VTAIL.n164 B 0.025949f
C451 VTAIL.n165 B 0.011624f
C452 VTAIL.n166 B 0.010978f
C453 VTAIL.n167 B 0.02043f
C454 VTAIL.n168 B 0.02043f
C455 VTAIL.n169 B 0.010978f
C456 VTAIL.n170 B 0.011624f
C457 VTAIL.n171 B 0.025949f
C458 VTAIL.n172 B 0.025949f
C459 VTAIL.n173 B 0.011624f
C460 VTAIL.n174 B 0.010978f
C461 VTAIL.n175 B 0.02043f
C462 VTAIL.n176 B 0.02043f
C463 VTAIL.n177 B 0.010978f
C464 VTAIL.n178 B 0.011624f
C465 VTAIL.n179 B 0.025949f
C466 VTAIL.n180 B 0.025949f
C467 VTAIL.n181 B 0.011624f
C468 VTAIL.n182 B 0.010978f
C469 VTAIL.n183 B 0.02043f
C470 VTAIL.n184 B 0.02043f
C471 VTAIL.n185 B 0.010978f
C472 VTAIL.n186 B 0.011624f
C473 VTAIL.n187 B 0.025949f
C474 VTAIL.n188 B 0.025949f
C475 VTAIL.n189 B 0.011624f
C476 VTAIL.n190 B 0.010978f
C477 VTAIL.n191 B 0.02043f
C478 VTAIL.n192 B 0.052806f
C479 VTAIL.n193 B 0.010978f
C480 VTAIL.n194 B 0.011624f
C481 VTAIL.n195 B 0.052275f
C482 VTAIL.n196 B 0.044308f
C483 VTAIL.n197 B 1.19413f
C484 VTAIL.n198 B 0.011518f
C485 VTAIL.n199 B 0.025949f
C486 VTAIL.n200 B 0.011624f
C487 VTAIL.n201 B 0.02043f
C488 VTAIL.n202 B 0.010978f
C489 VTAIL.n203 B 0.025949f
C490 VTAIL.n204 B 0.011624f
C491 VTAIL.n205 B 0.02043f
C492 VTAIL.n206 B 0.010978f
C493 VTAIL.n207 B 0.025949f
C494 VTAIL.n208 B 0.011624f
C495 VTAIL.n209 B 0.02043f
C496 VTAIL.n210 B 0.010978f
C497 VTAIL.n211 B 0.025949f
C498 VTAIL.n212 B 0.011624f
C499 VTAIL.n213 B 0.02043f
C500 VTAIL.n214 B 0.010978f
C501 VTAIL.n215 B 0.025949f
C502 VTAIL.n216 B 0.011624f
C503 VTAIL.n217 B 1.04458f
C504 VTAIL.n218 B 0.010978f
C505 VTAIL.t3 B 0.042574f
C506 VTAIL.n219 B 0.117679f
C507 VTAIL.n220 B 0.015329f
C508 VTAIL.n221 B 0.019462f
C509 VTAIL.n222 B 0.025949f
C510 VTAIL.n223 B 0.011624f
C511 VTAIL.n224 B 0.010978f
C512 VTAIL.n225 B 0.02043f
C513 VTAIL.n226 B 0.02043f
C514 VTAIL.n227 B 0.010978f
C515 VTAIL.n228 B 0.011624f
C516 VTAIL.n229 B 0.025949f
C517 VTAIL.n230 B 0.025949f
C518 VTAIL.n231 B 0.011624f
C519 VTAIL.n232 B 0.010978f
C520 VTAIL.n233 B 0.02043f
C521 VTAIL.n234 B 0.02043f
C522 VTAIL.n235 B 0.010978f
C523 VTAIL.n236 B 0.011624f
C524 VTAIL.n237 B 0.025949f
C525 VTAIL.n238 B 0.025949f
C526 VTAIL.n239 B 0.011624f
C527 VTAIL.n240 B 0.010978f
C528 VTAIL.n241 B 0.02043f
C529 VTAIL.n242 B 0.02043f
C530 VTAIL.n243 B 0.010978f
C531 VTAIL.n244 B 0.011624f
C532 VTAIL.n245 B 0.025949f
C533 VTAIL.n246 B 0.025949f
C534 VTAIL.n247 B 0.011624f
C535 VTAIL.n248 B 0.010978f
C536 VTAIL.n249 B 0.02043f
C537 VTAIL.n250 B 0.02043f
C538 VTAIL.n251 B 0.010978f
C539 VTAIL.n252 B 0.011624f
C540 VTAIL.n253 B 0.025949f
C541 VTAIL.n254 B 0.025949f
C542 VTAIL.n255 B 0.011624f
C543 VTAIL.n256 B 0.010978f
C544 VTAIL.n257 B 0.02043f
C545 VTAIL.n258 B 0.052806f
C546 VTAIL.n259 B 0.010978f
C547 VTAIL.n260 B 0.011624f
C548 VTAIL.n261 B 0.052275f
C549 VTAIL.n262 B 0.044308f
C550 VTAIL.n263 B 1.12815f
C551 VN.t0 B 2.53029f
C552 VN.t1 B 2.93097f
.ends

