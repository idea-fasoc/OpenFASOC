* NGSPICE file created from diff_pair_sample_1227.ext - technology: sky130A

.subckt diff_pair_sample_1227 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=1.72425 ps=10.78 w=10.45 l=3.29
X1 VDD1.t7 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X2 VDD1.t6 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=4.0755 ps=21.68 w=10.45 l=3.29
X3 VDD1.t5 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X4 VDD1.t4 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=4.0755 ps=21.68 w=10.45 l=3.29
X5 VTAIL.t14 VN.t1 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=1.72425 ps=10.78 w=10.45 l=3.29
X6 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=0 ps=0 w=10.45 l=3.29
X7 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=0 ps=0 w=10.45 l=3.29
X8 VTAIL.t13 VN.t2 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X9 VDD2.t2 VN.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=4.0755 ps=21.68 w=10.45 l=3.29
X10 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=0 ps=0 w=10.45 l=3.29
X11 VTAIL.t11 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X12 VTAIL.t4 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=0 ps=0 w=10.45 l=3.29
X14 VTAIL.t7 VP.t5 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=1.72425 ps=10.78 w=10.45 l=3.29
X15 VDD2.t4 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X16 VTAIL.t2 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.0755 pd=21.68 as=1.72425 ps=10.78 w=10.45 l=3.29
X17 VTAIL.t6 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
X18 VDD2.t5 VN.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=4.0755 ps=21.68 w=10.45 l=3.29
X19 VDD2.t0 VN.t7 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.72425 pd=10.78 as=1.72425 ps=10.78 w=10.45 l=3.29
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n56 161.3
R8 VN.n55 VN.n40 161.3
R9 VN.n54 VN.n53 161.3
R10 VN.n52 VN.n41 161.3
R11 VN.n51 VN.n50 161.3
R12 VN.n49 VN.n42 161.3
R13 VN.n48 VN.n47 161.3
R14 VN.n46 VN.n43 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n21 161.3
R23 VN.n20 VN.n5 161.3
R24 VN.n19 VN.n18 161.3
R25 VN.n17 VN.n6 161.3
R26 VN.n16 VN.n15 161.3
R27 VN.n14 VN.n7 161.3
R28 VN.n13 VN.n12 161.3
R29 VN.n11 VN.n8 161.3
R30 VN.n45 VN.t3 108.425
R31 VN.n10 VN.t1 108.425
R32 VN.n34 VN.n0 81.2593
R33 VN.n69 VN.n35 81.2593
R34 VN.n9 VN.t7 76.5491
R35 VN.n4 VN.t2 76.5491
R36 VN.n0 VN.t6 76.5491
R37 VN.n44 VN.t4 76.5491
R38 VN.n39 VN.t5 76.5491
R39 VN.n35 VN.t0 76.5491
R40 VN.n45 VN.n44 71.6409
R41 VN.n10 VN.n9 71.6408
R42 VN.n15 VN.n6 56.5193
R43 VN.n50 VN.n41 56.5193
R44 VN VN.n69 53.1344
R45 VN.n26 VN.n2 53.1199
R46 VN.n61 VN.n37 53.1199
R47 VN.n30 VN.n2 27.8669
R48 VN.n65 VN.n37 27.8669
R49 VN.n13 VN.n8 24.4675
R50 VN.n14 VN.n13 24.4675
R51 VN.n15 VN.n14 24.4675
R52 VN.n19 VN.n6 24.4675
R53 VN.n20 VN.n19 24.4675
R54 VN.n21 VN.n20 24.4675
R55 VN.n25 VN.n24 24.4675
R56 VN.n26 VN.n25 24.4675
R57 VN.n31 VN.n30 24.4675
R58 VN.n32 VN.n31 24.4675
R59 VN.n50 VN.n49 24.4675
R60 VN.n49 VN.n48 24.4675
R61 VN.n48 VN.n43 24.4675
R62 VN.n61 VN.n60 24.4675
R63 VN.n60 VN.n59 24.4675
R64 VN.n56 VN.n55 24.4675
R65 VN.n55 VN.n54 24.4675
R66 VN.n54 VN.n41 24.4675
R67 VN.n67 VN.n66 24.4675
R68 VN.n66 VN.n65 24.4675
R69 VN.n24 VN.n4 21.5315
R70 VN.n59 VN.n39 21.5315
R71 VN.n32 VN.n0 8.80862
R72 VN.n67 VN.n35 8.80862
R73 VN.n46 VN.n45 4.46857
R74 VN.n11 VN.n10 4.46857
R75 VN.n9 VN.n8 2.93654
R76 VN.n21 VN.n4 2.93654
R77 VN.n44 VN.n43 2.93654
R78 VN.n56 VN.n39 2.93654
R79 VN.n69 VN.n68 0.354971
R80 VN.n34 VN.n33 0.354971
R81 VN VN.n34 0.26696
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n40 0.189894
R90 VN.n53 VN.n40 0.189894
R91 VN.n53 VN.n52 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n42 0.189894
R94 VN.n47 VN.n42 0.189894
R95 VN.n47 VN.n46 0.189894
R96 VN.n12 VN.n11 0.189894
R97 VN.n12 VN.n7 0.189894
R98 VN.n16 VN.n7 0.189894
R99 VN.n17 VN.n16 0.189894
R100 VN.n18 VN.n17 0.189894
R101 VN.n18 VN.n5 0.189894
R102 VN.n22 VN.n5 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VDD2.n2 VDD2.n1 66.509
R111 VDD2.n2 VDD2.n0 66.509
R112 VDD2 VDD2.n5 66.5062
R113 VDD2.n4 VDD2.n3 65.0042
R114 VDD2.n4 VDD2.n2 46.767
R115 VDD2.n5 VDD2.t3 1.89524
R116 VDD2.n5 VDD2.t2 1.89524
R117 VDD2.n3 VDD2.t6 1.89524
R118 VDD2.n3 VDD2.t4 1.89524
R119 VDD2.n1 VDD2.t1 1.89524
R120 VDD2.n1 VDD2.t5 1.89524
R121 VDD2.n0 VDD2.t7 1.89524
R122 VDD2.n0 VDD2.t0 1.89524
R123 VDD2 VDD2.n4 1.61903
R124 VTAIL.n11 VTAIL.t7 50.2202
R125 VTAIL.n10 VTAIL.t12 50.2202
R126 VTAIL.n7 VTAIL.t15 50.2202
R127 VTAIL.n15 VTAIL.t9 50.2199
R128 VTAIL.n2 VTAIL.t14 50.2199
R129 VTAIL.n3 VTAIL.t1 50.2199
R130 VTAIL.n6 VTAIL.t2 50.2199
R131 VTAIL.n14 VTAIL.t3 50.2199
R132 VTAIL.n13 VTAIL.n12 48.3254
R133 VTAIL.n9 VTAIL.n8 48.3254
R134 VTAIL.n1 VTAIL.n0 48.3252
R135 VTAIL.n5 VTAIL.n4 48.3252
R136 VTAIL.n15 VTAIL.n14 24.4962
R137 VTAIL.n7 VTAIL.n6 24.4962
R138 VTAIL.n9 VTAIL.n7 3.12119
R139 VTAIL.n10 VTAIL.n9 3.12119
R140 VTAIL.n13 VTAIL.n11 3.12119
R141 VTAIL.n14 VTAIL.n13 3.12119
R142 VTAIL.n6 VTAIL.n5 3.12119
R143 VTAIL.n5 VTAIL.n3 3.12119
R144 VTAIL.n2 VTAIL.n1 3.12119
R145 VTAIL VTAIL.n15 3.063
R146 VTAIL.n0 VTAIL.t8 1.89524
R147 VTAIL.n0 VTAIL.t13 1.89524
R148 VTAIL.n4 VTAIL.t0 1.89524
R149 VTAIL.n4 VTAIL.t4 1.89524
R150 VTAIL.n12 VTAIL.t5 1.89524
R151 VTAIL.n12 VTAIL.t6 1.89524
R152 VTAIL.n8 VTAIL.t10 1.89524
R153 VTAIL.n8 VTAIL.t11 1.89524
R154 VTAIL.n11 VTAIL.n10 0.470328
R155 VTAIL.n3 VTAIL.n2 0.470328
R156 VTAIL VTAIL.n1 0.0586897
R157 B.n924 B.n923 585
R158 B.n325 B.n154 585
R159 B.n324 B.n323 585
R160 B.n322 B.n321 585
R161 B.n320 B.n319 585
R162 B.n318 B.n317 585
R163 B.n316 B.n315 585
R164 B.n314 B.n313 585
R165 B.n312 B.n311 585
R166 B.n310 B.n309 585
R167 B.n308 B.n307 585
R168 B.n306 B.n305 585
R169 B.n304 B.n303 585
R170 B.n302 B.n301 585
R171 B.n300 B.n299 585
R172 B.n298 B.n297 585
R173 B.n296 B.n295 585
R174 B.n294 B.n293 585
R175 B.n292 B.n291 585
R176 B.n290 B.n289 585
R177 B.n288 B.n287 585
R178 B.n286 B.n285 585
R179 B.n284 B.n283 585
R180 B.n282 B.n281 585
R181 B.n280 B.n279 585
R182 B.n278 B.n277 585
R183 B.n276 B.n275 585
R184 B.n274 B.n273 585
R185 B.n272 B.n271 585
R186 B.n270 B.n269 585
R187 B.n268 B.n267 585
R188 B.n266 B.n265 585
R189 B.n264 B.n263 585
R190 B.n262 B.n261 585
R191 B.n260 B.n259 585
R192 B.n258 B.n257 585
R193 B.n256 B.n255 585
R194 B.n253 B.n252 585
R195 B.n251 B.n250 585
R196 B.n249 B.n248 585
R197 B.n247 B.n246 585
R198 B.n245 B.n244 585
R199 B.n243 B.n242 585
R200 B.n241 B.n240 585
R201 B.n239 B.n238 585
R202 B.n237 B.n236 585
R203 B.n235 B.n234 585
R204 B.n232 B.n231 585
R205 B.n230 B.n229 585
R206 B.n228 B.n227 585
R207 B.n226 B.n225 585
R208 B.n224 B.n223 585
R209 B.n222 B.n221 585
R210 B.n220 B.n219 585
R211 B.n218 B.n217 585
R212 B.n216 B.n215 585
R213 B.n214 B.n213 585
R214 B.n212 B.n211 585
R215 B.n210 B.n209 585
R216 B.n208 B.n207 585
R217 B.n206 B.n205 585
R218 B.n204 B.n203 585
R219 B.n202 B.n201 585
R220 B.n200 B.n199 585
R221 B.n198 B.n197 585
R222 B.n196 B.n195 585
R223 B.n194 B.n193 585
R224 B.n192 B.n191 585
R225 B.n190 B.n189 585
R226 B.n188 B.n187 585
R227 B.n186 B.n185 585
R228 B.n184 B.n183 585
R229 B.n182 B.n181 585
R230 B.n180 B.n179 585
R231 B.n178 B.n177 585
R232 B.n176 B.n175 585
R233 B.n174 B.n173 585
R234 B.n172 B.n171 585
R235 B.n170 B.n169 585
R236 B.n168 B.n167 585
R237 B.n166 B.n165 585
R238 B.n164 B.n163 585
R239 B.n162 B.n161 585
R240 B.n160 B.n159 585
R241 B.n922 B.n112 585
R242 B.n927 B.n112 585
R243 B.n921 B.n111 585
R244 B.n928 B.n111 585
R245 B.n920 B.n919 585
R246 B.n919 B.n107 585
R247 B.n918 B.n106 585
R248 B.n934 B.n106 585
R249 B.n917 B.n105 585
R250 B.n935 B.n105 585
R251 B.n916 B.n104 585
R252 B.n936 B.n104 585
R253 B.n915 B.n914 585
R254 B.n914 B.n100 585
R255 B.n913 B.n99 585
R256 B.n942 B.n99 585
R257 B.n912 B.n98 585
R258 B.n943 B.n98 585
R259 B.n911 B.n97 585
R260 B.n944 B.n97 585
R261 B.n910 B.n909 585
R262 B.n909 B.n93 585
R263 B.n908 B.n92 585
R264 B.n950 B.n92 585
R265 B.n907 B.n91 585
R266 B.n951 B.n91 585
R267 B.n906 B.n90 585
R268 B.n952 B.n90 585
R269 B.n905 B.n904 585
R270 B.n904 B.n86 585
R271 B.n903 B.n85 585
R272 B.n958 B.n85 585
R273 B.n902 B.n84 585
R274 B.n959 B.n84 585
R275 B.n901 B.n83 585
R276 B.n960 B.n83 585
R277 B.n900 B.n899 585
R278 B.n899 B.n79 585
R279 B.n898 B.n78 585
R280 B.n966 B.n78 585
R281 B.n897 B.n77 585
R282 B.n967 B.n77 585
R283 B.n896 B.n76 585
R284 B.n968 B.n76 585
R285 B.n895 B.n894 585
R286 B.n894 B.n75 585
R287 B.n893 B.n71 585
R288 B.n974 B.n71 585
R289 B.n892 B.n70 585
R290 B.n975 B.n70 585
R291 B.n891 B.n69 585
R292 B.n976 B.n69 585
R293 B.n890 B.n889 585
R294 B.n889 B.n65 585
R295 B.n888 B.n64 585
R296 B.n982 B.n64 585
R297 B.n887 B.n63 585
R298 B.n983 B.n63 585
R299 B.n886 B.n62 585
R300 B.n984 B.n62 585
R301 B.n885 B.n884 585
R302 B.n884 B.n58 585
R303 B.n883 B.n57 585
R304 B.n990 B.n57 585
R305 B.n882 B.n56 585
R306 B.n991 B.n56 585
R307 B.n881 B.n55 585
R308 B.n992 B.n55 585
R309 B.n880 B.n879 585
R310 B.n879 B.n51 585
R311 B.n878 B.n50 585
R312 B.n998 B.n50 585
R313 B.n877 B.n49 585
R314 B.n999 B.n49 585
R315 B.n876 B.n48 585
R316 B.n1000 B.n48 585
R317 B.n875 B.n874 585
R318 B.n874 B.n44 585
R319 B.n873 B.n43 585
R320 B.n1006 B.n43 585
R321 B.n872 B.n42 585
R322 B.n1007 B.n42 585
R323 B.n871 B.n41 585
R324 B.n1008 B.n41 585
R325 B.n870 B.n869 585
R326 B.n869 B.n37 585
R327 B.n868 B.n36 585
R328 B.n1014 B.n36 585
R329 B.n867 B.n35 585
R330 B.n1015 B.n35 585
R331 B.n866 B.n34 585
R332 B.n1016 B.n34 585
R333 B.n865 B.n864 585
R334 B.n864 B.n30 585
R335 B.n863 B.n29 585
R336 B.n1022 B.n29 585
R337 B.n862 B.n28 585
R338 B.n1023 B.n28 585
R339 B.n861 B.n27 585
R340 B.n1024 B.n27 585
R341 B.n860 B.n859 585
R342 B.n859 B.n23 585
R343 B.n858 B.n22 585
R344 B.n1030 B.n22 585
R345 B.n857 B.n21 585
R346 B.n1031 B.n21 585
R347 B.n856 B.n20 585
R348 B.n1032 B.n20 585
R349 B.n855 B.n854 585
R350 B.n854 B.n19 585
R351 B.n853 B.n15 585
R352 B.n1038 B.n15 585
R353 B.n852 B.n14 585
R354 B.n1039 B.n14 585
R355 B.n851 B.n13 585
R356 B.n1040 B.n13 585
R357 B.n850 B.n849 585
R358 B.n849 B.n12 585
R359 B.n848 B.n847 585
R360 B.n848 B.n8 585
R361 B.n846 B.n7 585
R362 B.n1047 B.n7 585
R363 B.n845 B.n6 585
R364 B.n1048 B.n6 585
R365 B.n844 B.n5 585
R366 B.n1049 B.n5 585
R367 B.n843 B.n842 585
R368 B.n842 B.n4 585
R369 B.n841 B.n326 585
R370 B.n841 B.n840 585
R371 B.n831 B.n327 585
R372 B.n328 B.n327 585
R373 B.n833 B.n832 585
R374 B.n834 B.n833 585
R375 B.n830 B.n333 585
R376 B.n333 B.n332 585
R377 B.n829 B.n828 585
R378 B.n828 B.n827 585
R379 B.n335 B.n334 585
R380 B.n820 B.n335 585
R381 B.n819 B.n818 585
R382 B.n821 B.n819 585
R383 B.n817 B.n340 585
R384 B.n340 B.n339 585
R385 B.n816 B.n815 585
R386 B.n815 B.n814 585
R387 B.n342 B.n341 585
R388 B.n343 B.n342 585
R389 B.n807 B.n806 585
R390 B.n808 B.n807 585
R391 B.n805 B.n348 585
R392 B.n348 B.n347 585
R393 B.n804 B.n803 585
R394 B.n803 B.n802 585
R395 B.n350 B.n349 585
R396 B.n351 B.n350 585
R397 B.n795 B.n794 585
R398 B.n796 B.n795 585
R399 B.n793 B.n356 585
R400 B.n356 B.n355 585
R401 B.n792 B.n791 585
R402 B.n791 B.n790 585
R403 B.n358 B.n357 585
R404 B.n359 B.n358 585
R405 B.n783 B.n782 585
R406 B.n784 B.n783 585
R407 B.n781 B.n364 585
R408 B.n364 B.n363 585
R409 B.n780 B.n779 585
R410 B.n779 B.n778 585
R411 B.n366 B.n365 585
R412 B.n367 B.n366 585
R413 B.n771 B.n770 585
R414 B.n772 B.n771 585
R415 B.n769 B.n372 585
R416 B.n372 B.n371 585
R417 B.n768 B.n767 585
R418 B.n767 B.n766 585
R419 B.n374 B.n373 585
R420 B.n375 B.n374 585
R421 B.n759 B.n758 585
R422 B.n760 B.n759 585
R423 B.n757 B.n380 585
R424 B.n380 B.n379 585
R425 B.n756 B.n755 585
R426 B.n755 B.n754 585
R427 B.n382 B.n381 585
R428 B.n383 B.n382 585
R429 B.n747 B.n746 585
R430 B.n748 B.n747 585
R431 B.n745 B.n388 585
R432 B.n388 B.n387 585
R433 B.n744 B.n743 585
R434 B.n743 B.n742 585
R435 B.n390 B.n389 585
R436 B.n391 B.n390 585
R437 B.n735 B.n734 585
R438 B.n736 B.n735 585
R439 B.n733 B.n396 585
R440 B.n396 B.n395 585
R441 B.n732 B.n731 585
R442 B.n731 B.n730 585
R443 B.n398 B.n397 585
R444 B.n723 B.n398 585
R445 B.n722 B.n721 585
R446 B.n724 B.n722 585
R447 B.n720 B.n403 585
R448 B.n403 B.n402 585
R449 B.n719 B.n718 585
R450 B.n718 B.n717 585
R451 B.n405 B.n404 585
R452 B.n406 B.n405 585
R453 B.n710 B.n709 585
R454 B.n711 B.n710 585
R455 B.n708 B.n411 585
R456 B.n411 B.n410 585
R457 B.n707 B.n706 585
R458 B.n706 B.n705 585
R459 B.n413 B.n412 585
R460 B.n414 B.n413 585
R461 B.n698 B.n697 585
R462 B.n699 B.n698 585
R463 B.n696 B.n419 585
R464 B.n419 B.n418 585
R465 B.n695 B.n694 585
R466 B.n694 B.n693 585
R467 B.n421 B.n420 585
R468 B.n422 B.n421 585
R469 B.n686 B.n685 585
R470 B.n687 B.n686 585
R471 B.n684 B.n426 585
R472 B.n430 B.n426 585
R473 B.n683 B.n682 585
R474 B.n682 B.n681 585
R475 B.n428 B.n427 585
R476 B.n429 B.n428 585
R477 B.n674 B.n673 585
R478 B.n675 B.n674 585
R479 B.n672 B.n435 585
R480 B.n435 B.n434 585
R481 B.n671 B.n670 585
R482 B.n670 B.n669 585
R483 B.n437 B.n436 585
R484 B.n438 B.n437 585
R485 B.n662 B.n661 585
R486 B.n663 B.n662 585
R487 B.n660 B.n443 585
R488 B.n443 B.n442 585
R489 B.n655 B.n654 585
R490 B.n653 B.n487 585
R491 B.n652 B.n486 585
R492 B.n657 B.n486 585
R493 B.n651 B.n650 585
R494 B.n649 B.n648 585
R495 B.n647 B.n646 585
R496 B.n645 B.n644 585
R497 B.n643 B.n642 585
R498 B.n641 B.n640 585
R499 B.n639 B.n638 585
R500 B.n637 B.n636 585
R501 B.n635 B.n634 585
R502 B.n633 B.n632 585
R503 B.n631 B.n630 585
R504 B.n629 B.n628 585
R505 B.n627 B.n626 585
R506 B.n625 B.n624 585
R507 B.n623 B.n622 585
R508 B.n621 B.n620 585
R509 B.n619 B.n618 585
R510 B.n617 B.n616 585
R511 B.n615 B.n614 585
R512 B.n613 B.n612 585
R513 B.n611 B.n610 585
R514 B.n609 B.n608 585
R515 B.n607 B.n606 585
R516 B.n605 B.n604 585
R517 B.n603 B.n602 585
R518 B.n601 B.n600 585
R519 B.n599 B.n598 585
R520 B.n597 B.n596 585
R521 B.n595 B.n594 585
R522 B.n593 B.n592 585
R523 B.n591 B.n590 585
R524 B.n589 B.n588 585
R525 B.n587 B.n586 585
R526 B.n585 B.n584 585
R527 B.n583 B.n582 585
R528 B.n581 B.n580 585
R529 B.n579 B.n578 585
R530 B.n577 B.n576 585
R531 B.n575 B.n574 585
R532 B.n573 B.n572 585
R533 B.n571 B.n570 585
R534 B.n569 B.n568 585
R535 B.n567 B.n566 585
R536 B.n565 B.n564 585
R537 B.n563 B.n562 585
R538 B.n561 B.n560 585
R539 B.n559 B.n558 585
R540 B.n557 B.n556 585
R541 B.n555 B.n554 585
R542 B.n553 B.n552 585
R543 B.n551 B.n550 585
R544 B.n549 B.n548 585
R545 B.n547 B.n546 585
R546 B.n545 B.n544 585
R547 B.n543 B.n542 585
R548 B.n541 B.n540 585
R549 B.n539 B.n538 585
R550 B.n537 B.n536 585
R551 B.n535 B.n534 585
R552 B.n533 B.n532 585
R553 B.n531 B.n530 585
R554 B.n529 B.n528 585
R555 B.n527 B.n526 585
R556 B.n525 B.n524 585
R557 B.n523 B.n522 585
R558 B.n521 B.n520 585
R559 B.n519 B.n518 585
R560 B.n517 B.n516 585
R561 B.n515 B.n514 585
R562 B.n513 B.n512 585
R563 B.n511 B.n510 585
R564 B.n509 B.n508 585
R565 B.n507 B.n506 585
R566 B.n505 B.n504 585
R567 B.n503 B.n502 585
R568 B.n501 B.n500 585
R569 B.n499 B.n498 585
R570 B.n497 B.n496 585
R571 B.n495 B.n494 585
R572 B.n445 B.n444 585
R573 B.n659 B.n658 585
R574 B.n658 B.n657 585
R575 B.n441 B.n440 585
R576 B.n442 B.n441 585
R577 B.n665 B.n664 585
R578 B.n664 B.n663 585
R579 B.n666 B.n439 585
R580 B.n439 B.n438 585
R581 B.n668 B.n667 585
R582 B.n669 B.n668 585
R583 B.n433 B.n432 585
R584 B.n434 B.n433 585
R585 B.n677 B.n676 585
R586 B.n676 B.n675 585
R587 B.n678 B.n431 585
R588 B.n431 B.n429 585
R589 B.n680 B.n679 585
R590 B.n681 B.n680 585
R591 B.n425 B.n424 585
R592 B.n430 B.n425 585
R593 B.n689 B.n688 585
R594 B.n688 B.n687 585
R595 B.n690 B.n423 585
R596 B.n423 B.n422 585
R597 B.n692 B.n691 585
R598 B.n693 B.n692 585
R599 B.n417 B.n416 585
R600 B.n418 B.n417 585
R601 B.n701 B.n700 585
R602 B.n700 B.n699 585
R603 B.n702 B.n415 585
R604 B.n415 B.n414 585
R605 B.n704 B.n703 585
R606 B.n705 B.n704 585
R607 B.n409 B.n408 585
R608 B.n410 B.n409 585
R609 B.n713 B.n712 585
R610 B.n712 B.n711 585
R611 B.n714 B.n407 585
R612 B.n407 B.n406 585
R613 B.n716 B.n715 585
R614 B.n717 B.n716 585
R615 B.n401 B.n400 585
R616 B.n402 B.n401 585
R617 B.n726 B.n725 585
R618 B.n725 B.n724 585
R619 B.n727 B.n399 585
R620 B.n723 B.n399 585
R621 B.n729 B.n728 585
R622 B.n730 B.n729 585
R623 B.n394 B.n393 585
R624 B.n395 B.n394 585
R625 B.n738 B.n737 585
R626 B.n737 B.n736 585
R627 B.n739 B.n392 585
R628 B.n392 B.n391 585
R629 B.n741 B.n740 585
R630 B.n742 B.n741 585
R631 B.n386 B.n385 585
R632 B.n387 B.n386 585
R633 B.n750 B.n749 585
R634 B.n749 B.n748 585
R635 B.n751 B.n384 585
R636 B.n384 B.n383 585
R637 B.n753 B.n752 585
R638 B.n754 B.n753 585
R639 B.n378 B.n377 585
R640 B.n379 B.n378 585
R641 B.n762 B.n761 585
R642 B.n761 B.n760 585
R643 B.n763 B.n376 585
R644 B.n376 B.n375 585
R645 B.n765 B.n764 585
R646 B.n766 B.n765 585
R647 B.n370 B.n369 585
R648 B.n371 B.n370 585
R649 B.n774 B.n773 585
R650 B.n773 B.n772 585
R651 B.n775 B.n368 585
R652 B.n368 B.n367 585
R653 B.n777 B.n776 585
R654 B.n778 B.n777 585
R655 B.n362 B.n361 585
R656 B.n363 B.n362 585
R657 B.n786 B.n785 585
R658 B.n785 B.n784 585
R659 B.n787 B.n360 585
R660 B.n360 B.n359 585
R661 B.n789 B.n788 585
R662 B.n790 B.n789 585
R663 B.n354 B.n353 585
R664 B.n355 B.n354 585
R665 B.n798 B.n797 585
R666 B.n797 B.n796 585
R667 B.n799 B.n352 585
R668 B.n352 B.n351 585
R669 B.n801 B.n800 585
R670 B.n802 B.n801 585
R671 B.n346 B.n345 585
R672 B.n347 B.n346 585
R673 B.n810 B.n809 585
R674 B.n809 B.n808 585
R675 B.n811 B.n344 585
R676 B.n344 B.n343 585
R677 B.n813 B.n812 585
R678 B.n814 B.n813 585
R679 B.n338 B.n337 585
R680 B.n339 B.n338 585
R681 B.n823 B.n822 585
R682 B.n822 B.n821 585
R683 B.n824 B.n336 585
R684 B.n820 B.n336 585
R685 B.n826 B.n825 585
R686 B.n827 B.n826 585
R687 B.n331 B.n330 585
R688 B.n332 B.n331 585
R689 B.n836 B.n835 585
R690 B.n835 B.n834 585
R691 B.n837 B.n329 585
R692 B.n329 B.n328 585
R693 B.n839 B.n838 585
R694 B.n840 B.n839 585
R695 B.n3 B.n0 585
R696 B.n4 B.n3 585
R697 B.n1046 B.n1 585
R698 B.n1047 B.n1046 585
R699 B.n1045 B.n1044 585
R700 B.n1045 B.n8 585
R701 B.n1043 B.n9 585
R702 B.n12 B.n9 585
R703 B.n1042 B.n1041 585
R704 B.n1041 B.n1040 585
R705 B.n11 B.n10 585
R706 B.n1039 B.n11 585
R707 B.n1037 B.n1036 585
R708 B.n1038 B.n1037 585
R709 B.n1035 B.n16 585
R710 B.n19 B.n16 585
R711 B.n1034 B.n1033 585
R712 B.n1033 B.n1032 585
R713 B.n18 B.n17 585
R714 B.n1031 B.n18 585
R715 B.n1029 B.n1028 585
R716 B.n1030 B.n1029 585
R717 B.n1027 B.n24 585
R718 B.n24 B.n23 585
R719 B.n1026 B.n1025 585
R720 B.n1025 B.n1024 585
R721 B.n26 B.n25 585
R722 B.n1023 B.n26 585
R723 B.n1021 B.n1020 585
R724 B.n1022 B.n1021 585
R725 B.n1019 B.n31 585
R726 B.n31 B.n30 585
R727 B.n1018 B.n1017 585
R728 B.n1017 B.n1016 585
R729 B.n33 B.n32 585
R730 B.n1015 B.n33 585
R731 B.n1013 B.n1012 585
R732 B.n1014 B.n1013 585
R733 B.n1011 B.n38 585
R734 B.n38 B.n37 585
R735 B.n1010 B.n1009 585
R736 B.n1009 B.n1008 585
R737 B.n40 B.n39 585
R738 B.n1007 B.n40 585
R739 B.n1005 B.n1004 585
R740 B.n1006 B.n1005 585
R741 B.n1003 B.n45 585
R742 B.n45 B.n44 585
R743 B.n1002 B.n1001 585
R744 B.n1001 B.n1000 585
R745 B.n47 B.n46 585
R746 B.n999 B.n47 585
R747 B.n997 B.n996 585
R748 B.n998 B.n997 585
R749 B.n995 B.n52 585
R750 B.n52 B.n51 585
R751 B.n994 B.n993 585
R752 B.n993 B.n992 585
R753 B.n54 B.n53 585
R754 B.n991 B.n54 585
R755 B.n989 B.n988 585
R756 B.n990 B.n989 585
R757 B.n987 B.n59 585
R758 B.n59 B.n58 585
R759 B.n986 B.n985 585
R760 B.n985 B.n984 585
R761 B.n61 B.n60 585
R762 B.n983 B.n61 585
R763 B.n981 B.n980 585
R764 B.n982 B.n981 585
R765 B.n979 B.n66 585
R766 B.n66 B.n65 585
R767 B.n978 B.n977 585
R768 B.n977 B.n976 585
R769 B.n68 B.n67 585
R770 B.n975 B.n68 585
R771 B.n973 B.n972 585
R772 B.n974 B.n973 585
R773 B.n971 B.n72 585
R774 B.n75 B.n72 585
R775 B.n970 B.n969 585
R776 B.n969 B.n968 585
R777 B.n74 B.n73 585
R778 B.n967 B.n74 585
R779 B.n965 B.n964 585
R780 B.n966 B.n965 585
R781 B.n963 B.n80 585
R782 B.n80 B.n79 585
R783 B.n962 B.n961 585
R784 B.n961 B.n960 585
R785 B.n82 B.n81 585
R786 B.n959 B.n82 585
R787 B.n957 B.n956 585
R788 B.n958 B.n957 585
R789 B.n955 B.n87 585
R790 B.n87 B.n86 585
R791 B.n954 B.n953 585
R792 B.n953 B.n952 585
R793 B.n89 B.n88 585
R794 B.n951 B.n89 585
R795 B.n949 B.n948 585
R796 B.n950 B.n949 585
R797 B.n947 B.n94 585
R798 B.n94 B.n93 585
R799 B.n946 B.n945 585
R800 B.n945 B.n944 585
R801 B.n96 B.n95 585
R802 B.n943 B.n96 585
R803 B.n941 B.n940 585
R804 B.n942 B.n941 585
R805 B.n939 B.n101 585
R806 B.n101 B.n100 585
R807 B.n938 B.n937 585
R808 B.n937 B.n936 585
R809 B.n103 B.n102 585
R810 B.n935 B.n103 585
R811 B.n933 B.n932 585
R812 B.n934 B.n933 585
R813 B.n931 B.n108 585
R814 B.n108 B.n107 585
R815 B.n930 B.n929 585
R816 B.n929 B.n928 585
R817 B.n110 B.n109 585
R818 B.n927 B.n110 585
R819 B.n1050 B.n1049 585
R820 B.n1048 B.n2 585
R821 B.n159 B.n110 449.257
R822 B.n924 B.n112 449.257
R823 B.n658 B.n443 449.257
R824 B.n655 B.n441 449.257
R825 B.n157 B.t12 285.443
R826 B.n155 B.t8 285.443
R827 B.n491 B.t15 285.443
R828 B.n488 B.t19 285.443
R829 B.n926 B.n925 256.663
R830 B.n926 B.n153 256.663
R831 B.n926 B.n152 256.663
R832 B.n926 B.n151 256.663
R833 B.n926 B.n150 256.663
R834 B.n926 B.n149 256.663
R835 B.n926 B.n148 256.663
R836 B.n926 B.n147 256.663
R837 B.n926 B.n146 256.663
R838 B.n926 B.n145 256.663
R839 B.n926 B.n144 256.663
R840 B.n926 B.n143 256.663
R841 B.n926 B.n142 256.663
R842 B.n926 B.n141 256.663
R843 B.n926 B.n140 256.663
R844 B.n926 B.n139 256.663
R845 B.n926 B.n138 256.663
R846 B.n926 B.n137 256.663
R847 B.n926 B.n136 256.663
R848 B.n926 B.n135 256.663
R849 B.n926 B.n134 256.663
R850 B.n926 B.n133 256.663
R851 B.n926 B.n132 256.663
R852 B.n926 B.n131 256.663
R853 B.n926 B.n130 256.663
R854 B.n926 B.n129 256.663
R855 B.n926 B.n128 256.663
R856 B.n926 B.n127 256.663
R857 B.n926 B.n126 256.663
R858 B.n926 B.n125 256.663
R859 B.n926 B.n124 256.663
R860 B.n926 B.n123 256.663
R861 B.n926 B.n122 256.663
R862 B.n926 B.n121 256.663
R863 B.n926 B.n120 256.663
R864 B.n926 B.n119 256.663
R865 B.n926 B.n118 256.663
R866 B.n926 B.n117 256.663
R867 B.n926 B.n116 256.663
R868 B.n926 B.n115 256.663
R869 B.n926 B.n114 256.663
R870 B.n926 B.n113 256.663
R871 B.n657 B.n656 256.663
R872 B.n657 B.n446 256.663
R873 B.n657 B.n447 256.663
R874 B.n657 B.n448 256.663
R875 B.n657 B.n449 256.663
R876 B.n657 B.n450 256.663
R877 B.n657 B.n451 256.663
R878 B.n657 B.n452 256.663
R879 B.n657 B.n453 256.663
R880 B.n657 B.n454 256.663
R881 B.n657 B.n455 256.663
R882 B.n657 B.n456 256.663
R883 B.n657 B.n457 256.663
R884 B.n657 B.n458 256.663
R885 B.n657 B.n459 256.663
R886 B.n657 B.n460 256.663
R887 B.n657 B.n461 256.663
R888 B.n657 B.n462 256.663
R889 B.n657 B.n463 256.663
R890 B.n657 B.n464 256.663
R891 B.n657 B.n465 256.663
R892 B.n657 B.n466 256.663
R893 B.n657 B.n467 256.663
R894 B.n657 B.n468 256.663
R895 B.n657 B.n469 256.663
R896 B.n657 B.n470 256.663
R897 B.n657 B.n471 256.663
R898 B.n657 B.n472 256.663
R899 B.n657 B.n473 256.663
R900 B.n657 B.n474 256.663
R901 B.n657 B.n475 256.663
R902 B.n657 B.n476 256.663
R903 B.n657 B.n477 256.663
R904 B.n657 B.n478 256.663
R905 B.n657 B.n479 256.663
R906 B.n657 B.n480 256.663
R907 B.n657 B.n481 256.663
R908 B.n657 B.n482 256.663
R909 B.n657 B.n483 256.663
R910 B.n657 B.n484 256.663
R911 B.n657 B.n485 256.663
R912 B.n1052 B.n1051 256.663
R913 B.n163 B.n162 163.367
R914 B.n167 B.n166 163.367
R915 B.n171 B.n170 163.367
R916 B.n175 B.n174 163.367
R917 B.n179 B.n178 163.367
R918 B.n183 B.n182 163.367
R919 B.n187 B.n186 163.367
R920 B.n191 B.n190 163.367
R921 B.n195 B.n194 163.367
R922 B.n199 B.n198 163.367
R923 B.n203 B.n202 163.367
R924 B.n207 B.n206 163.367
R925 B.n211 B.n210 163.367
R926 B.n215 B.n214 163.367
R927 B.n219 B.n218 163.367
R928 B.n223 B.n222 163.367
R929 B.n227 B.n226 163.367
R930 B.n231 B.n230 163.367
R931 B.n236 B.n235 163.367
R932 B.n240 B.n239 163.367
R933 B.n244 B.n243 163.367
R934 B.n248 B.n247 163.367
R935 B.n252 B.n251 163.367
R936 B.n257 B.n256 163.367
R937 B.n261 B.n260 163.367
R938 B.n265 B.n264 163.367
R939 B.n269 B.n268 163.367
R940 B.n273 B.n272 163.367
R941 B.n277 B.n276 163.367
R942 B.n281 B.n280 163.367
R943 B.n285 B.n284 163.367
R944 B.n289 B.n288 163.367
R945 B.n293 B.n292 163.367
R946 B.n297 B.n296 163.367
R947 B.n301 B.n300 163.367
R948 B.n305 B.n304 163.367
R949 B.n309 B.n308 163.367
R950 B.n313 B.n312 163.367
R951 B.n317 B.n316 163.367
R952 B.n321 B.n320 163.367
R953 B.n323 B.n154 163.367
R954 B.n662 B.n443 163.367
R955 B.n662 B.n437 163.367
R956 B.n670 B.n437 163.367
R957 B.n670 B.n435 163.367
R958 B.n674 B.n435 163.367
R959 B.n674 B.n428 163.367
R960 B.n682 B.n428 163.367
R961 B.n682 B.n426 163.367
R962 B.n686 B.n426 163.367
R963 B.n686 B.n421 163.367
R964 B.n694 B.n421 163.367
R965 B.n694 B.n419 163.367
R966 B.n698 B.n419 163.367
R967 B.n698 B.n413 163.367
R968 B.n706 B.n413 163.367
R969 B.n706 B.n411 163.367
R970 B.n710 B.n411 163.367
R971 B.n710 B.n405 163.367
R972 B.n718 B.n405 163.367
R973 B.n718 B.n403 163.367
R974 B.n722 B.n403 163.367
R975 B.n722 B.n398 163.367
R976 B.n731 B.n398 163.367
R977 B.n731 B.n396 163.367
R978 B.n735 B.n396 163.367
R979 B.n735 B.n390 163.367
R980 B.n743 B.n390 163.367
R981 B.n743 B.n388 163.367
R982 B.n747 B.n388 163.367
R983 B.n747 B.n382 163.367
R984 B.n755 B.n382 163.367
R985 B.n755 B.n380 163.367
R986 B.n759 B.n380 163.367
R987 B.n759 B.n374 163.367
R988 B.n767 B.n374 163.367
R989 B.n767 B.n372 163.367
R990 B.n771 B.n372 163.367
R991 B.n771 B.n366 163.367
R992 B.n779 B.n366 163.367
R993 B.n779 B.n364 163.367
R994 B.n783 B.n364 163.367
R995 B.n783 B.n358 163.367
R996 B.n791 B.n358 163.367
R997 B.n791 B.n356 163.367
R998 B.n795 B.n356 163.367
R999 B.n795 B.n350 163.367
R1000 B.n803 B.n350 163.367
R1001 B.n803 B.n348 163.367
R1002 B.n807 B.n348 163.367
R1003 B.n807 B.n342 163.367
R1004 B.n815 B.n342 163.367
R1005 B.n815 B.n340 163.367
R1006 B.n819 B.n340 163.367
R1007 B.n819 B.n335 163.367
R1008 B.n828 B.n335 163.367
R1009 B.n828 B.n333 163.367
R1010 B.n833 B.n333 163.367
R1011 B.n833 B.n327 163.367
R1012 B.n841 B.n327 163.367
R1013 B.n842 B.n841 163.367
R1014 B.n842 B.n5 163.367
R1015 B.n6 B.n5 163.367
R1016 B.n7 B.n6 163.367
R1017 B.n848 B.n7 163.367
R1018 B.n849 B.n848 163.367
R1019 B.n849 B.n13 163.367
R1020 B.n14 B.n13 163.367
R1021 B.n15 B.n14 163.367
R1022 B.n854 B.n15 163.367
R1023 B.n854 B.n20 163.367
R1024 B.n21 B.n20 163.367
R1025 B.n22 B.n21 163.367
R1026 B.n859 B.n22 163.367
R1027 B.n859 B.n27 163.367
R1028 B.n28 B.n27 163.367
R1029 B.n29 B.n28 163.367
R1030 B.n864 B.n29 163.367
R1031 B.n864 B.n34 163.367
R1032 B.n35 B.n34 163.367
R1033 B.n36 B.n35 163.367
R1034 B.n869 B.n36 163.367
R1035 B.n869 B.n41 163.367
R1036 B.n42 B.n41 163.367
R1037 B.n43 B.n42 163.367
R1038 B.n874 B.n43 163.367
R1039 B.n874 B.n48 163.367
R1040 B.n49 B.n48 163.367
R1041 B.n50 B.n49 163.367
R1042 B.n879 B.n50 163.367
R1043 B.n879 B.n55 163.367
R1044 B.n56 B.n55 163.367
R1045 B.n57 B.n56 163.367
R1046 B.n884 B.n57 163.367
R1047 B.n884 B.n62 163.367
R1048 B.n63 B.n62 163.367
R1049 B.n64 B.n63 163.367
R1050 B.n889 B.n64 163.367
R1051 B.n889 B.n69 163.367
R1052 B.n70 B.n69 163.367
R1053 B.n71 B.n70 163.367
R1054 B.n894 B.n71 163.367
R1055 B.n894 B.n76 163.367
R1056 B.n77 B.n76 163.367
R1057 B.n78 B.n77 163.367
R1058 B.n899 B.n78 163.367
R1059 B.n899 B.n83 163.367
R1060 B.n84 B.n83 163.367
R1061 B.n85 B.n84 163.367
R1062 B.n904 B.n85 163.367
R1063 B.n904 B.n90 163.367
R1064 B.n91 B.n90 163.367
R1065 B.n92 B.n91 163.367
R1066 B.n909 B.n92 163.367
R1067 B.n909 B.n97 163.367
R1068 B.n98 B.n97 163.367
R1069 B.n99 B.n98 163.367
R1070 B.n914 B.n99 163.367
R1071 B.n914 B.n104 163.367
R1072 B.n105 B.n104 163.367
R1073 B.n106 B.n105 163.367
R1074 B.n919 B.n106 163.367
R1075 B.n919 B.n111 163.367
R1076 B.n112 B.n111 163.367
R1077 B.n487 B.n486 163.367
R1078 B.n650 B.n486 163.367
R1079 B.n648 B.n647 163.367
R1080 B.n644 B.n643 163.367
R1081 B.n640 B.n639 163.367
R1082 B.n636 B.n635 163.367
R1083 B.n632 B.n631 163.367
R1084 B.n628 B.n627 163.367
R1085 B.n624 B.n623 163.367
R1086 B.n620 B.n619 163.367
R1087 B.n616 B.n615 163.367
R1088 B.n612 B.n611 163.367
R1089 B.n608 B.n607 163.367
R1090 B.n604 B.n603 163.367
R1091 B.n600 B.n599 163.367
R1092 B.n596 B.n595 163.367
R1093 B.n592 B.n591 163.367
R1094 B.n588 B.n587 163.367
R1095 B.n584 B.n583 163.367
R1096 B.n580 B.n579 163.367
R1097 B.n576 B.n575 163.367
R1098 B.n572 B.n571 163.367
R1099 B.n568 B.n567 163.367
R1100 B.n564 B.n563 163.367
R1101 B.n560 B.n559 163.367
R1102 B.n556 B.n555 163.367
R1103 B.n552 B.n551 163.367
R1104 B.n548 B.n547 163.367
R1105 B.n544 B.n543 163.367
R1106 B.n540 B.n539 163.367
R1107 B.n536 B.n535 163.367
R1108 B.n532 B.n531 163.367
R1109 B.n528 B.n527 163.367
R1110 B.n524 B.n523 163.367
R1111 B.n520 B.n519 163.367
R1112 B.n516 B.n515 163.367
R1113 B.n512 B.n511 163.367
R1114 B.n508 B.n507 163.367
R1115 B.n504 B.n503 163.367
R1116 B.n500 B.n499 163.367
R1117 B.n496 B.n495 163.367
R1118 B.n658 B.n445 163.367
R1119 B.n664 B.n441 163.367
R1120 B.n664 B.n439 163.367
R1121 B.n668 B.n439 163.367
R1122 B.n668 B.n433 163.367
R1123 B.n676 B.n433 163.367
R1124 B.n676 B.n431 163.367
R1125 B.n680 B.n431 163.367
R1126 B.n680 B.n425 163.367
R1127 B.n688 B.n425 163.367
R1128 B.n688 B.n423 163.367
R1129 B.n692 B.n423 163.367
R1130 B.n692 B.n417 163.367
R1131 B.n700 B.n417 163.367
R1132 B.n700 B.n415 163.367
R1133 B.n704 B.n415 163.367
R1134 B.n704 B.n409 163.367
R1135 B.n712 B.n409 163.367
R1136 B.n712 B.n407 163.367
R1137 B.n716 B.n407 163.367
R1138 B.n716 B.n401 163.367
R1139 B.n725 B.n401 163.367
R1140 B.n725 B.n399 163.367
R1141 B.n729 B.n399 163.367
R1142 B.n729 B.n394 163.367
R1143 B.n737 B.n394 163.367
R1144 B.n737 B.n392 163.367
R1145 B.n741 B.n392 163.367
R1146 B.n741 B.n386 163.367
R1147 B.n749 B.n386 163.367
R1148 B.n749 B.n384 163.367
R1149 B.n753 B.n384 163.367
R1150 B.n753 B.n378 163.367
R1151 B.n761 B.n378 163.367
R1152 B.n761 B.n376 163.367
R1153 B.n765 B.n376 163.367
R1154 B.n765 B.n370 163.367
R1155 B.n773 B.n370 163.367
R1156 B.n773 B.n368 163.367
R1157 B.n777 B.n368 163.367
R1158 B.n777 B.n362 163.367
R1159 B.n785 B.n362 163.367
R1160 B.n785 B.n360 163.367
R1161 B.n789 B.n360 163.367
R1162 B.n789 B.n354 163.367
R1163 B.n797 B.n354 163.367
R1164 B.n797 B.n352 163.367
R1165 B.n801 B.n352 163.367
R1166 B.n801 B.n346 163.367
R1167 B.n809 B.n346 163.367
R1168 B.n809 B.n344 163.367
R1169 B.n813 B.n344 163.367
R1170 B.n813 B.n338 163.367
R1171 B.n822 B.n338 163.367
R1172 B.n822 B.n336 163.367
R1173 B.n826 B.n336 163.367
R1174 B.n826 B.n331 163.367
R1175 B.n835 B.n331 163.367
R1176 B.n835 B.n329 163.367
R1177 B.n839 B.n329 163.367
R1178 B.n839 B.n3 163.367
R1179 B.n1050 B.n3 163.367
R1180 B.n1046 B.n2 163.367
R1181 B.n1046 B.n1045 163.367
R1182 B.n1045 B.n9 163.367
R1183 B.n1041 B.n9 163.367
R1184 B.n1041 B.n11 163.367
R1185 B.n1037 B.n11 163.367
R1186 B.n1037 B.n16 163.367
R1187 B.n1033 B.n16 163.367
R1188 B.n1033 B.n18 163.367
R1189 B.n1029 B.n18 163.367
R1190 B.n1029 B.n24 163.367
R1191 B.n1025 B.n24 163.367
R1192 B.n1025 B.n26 163.367
R1193 B.n1021 B.n26 163.367
R1194 B.n1021 B.n31 163.367
R1195 B.n1017 B.n31 163.367
R1196 B.n1017 B.n33 163.367
R1197 B.n1013 B.n33 163.367
R1198 B.n1013 B.n38 163.367
R1199 B.n1009 B.n38 163.367
R1200 B.n1009 B.n40 163.367
R1201 B.n1005 B.n40 163.367
R1202 B.n1005 B.n45 163.367
R1203 B.n1001 B.n45 163.367
R1204 B.n1001 B.n47 163.367
R1205 B.n997 B.n47 163.367
R1206 B.n997 B.n52 163.367
R1207 B.n993 B.n52 163.367
R1208 B.n993 B.n54 163.367
R1209 B.n989 B.n54 163.367
R1210 B.n989 B.n59 163.367
R1211 B.n985 B.n59 163.367
R1212 B.n985 B.n61 163.367
R1213 B.n981 B.n61 163.367
R1214 B.n981 B.n66 163.367
R1215 B.n977 B.n66 163.367
R1216 B.n977 B.n68 163.367
R1217 B.n973 B.n68 163.367
R1218 B.n973 B.n72 163.367
R1219 B.n969 B.n72 163.367
R1220 B.n969 B.n74 163.367
R1221 B.n965 B.n74 163.367
R1222 B.n965 B.n80 163.367
R1223 B.n961 B.n80 163.367
R1224 B.n961 B.n82 163.367
R1225 B.n957 B.n82 163.367
R1226 B.n957 B.n87 163.367
R1227 B.n953 B.n87 163.367
R1228 B.n953 B.n89 163.367
R1229 B.n949 B.n89 163.367
R1230 B.n949 B.n94 163.367
R1231 B.n945 B.n94 163.367
R1232 B.n945 B.n96 163.367
R1233 B.n941 B.n96 163.367
R1234 B.n941 B.n101 163.367
R1235 B.n937 B.n101 163.367
R1236 B.n937 B.n103 163.367
R1237 B.n933 B.n103 163.367
R1238 B.n933 B.n108 163.367
R1239 B.n929 B.n108 163.367
R1240 B.n929 B.n110 163.367
R1241 B.n155 B.t10 143.087
R1242 B.n491 B.t18 143.087
R1243 B.n157 B.t13 143.073
R1244 B.n488 B.t21 143.073
R1245 B.n657 B.n442 79.0466
R1246 B.n927 B.n926 79.0466
R1247 B.n156 B.t11 72.8806
R1248 B.n492 B.t17 72.8806
R1249 B.n158 B.t14 72.8679
R1250 B.n489 B.t20 72.8679
R1251 B.n159 B.n113 71.676
R1252 B.n163 B.n114 71.676
R1253 B.n167 B.n115 71.676
R1254 B.n171 B.n116 71.676
R1255 B.n175 B.n117 71.676
R1256 B.n179 B.n118 71.676
R1257 B.n183 B.n119 71.676
R1258 B.n187 B.n120 71.676
R1259 B.n191 B.n121 71.676
R1260 B.n195 B.n122 71.676
R1261 B.n199 B.n123 71.676
R1262 B.n203 B.n124 71.676
R1263 B.n207 B.n125 71.676
R1264 B.n211 B.n126 71.676
R1265 B.n215 B.n127 71.676
R1266 B.n219 B.n128 71.676
R1267 B.n223 B.n129 71.676
R1268 B.n227 B.n130 71.676
R1269 B.n231 B.n131 71.676
R1270 B.n236 B.n132 71.676
R1271 B.n240 B.n133 71.676
R1272 B.n244 B.n134 71.676
R1273 B.n248 B.n135 71.676
R1274 B.n252 B.n136 71.676
R1275 B.n257 B.n137 71.676
R1276 B.n261 B.n138 71.676
R1277 B.n265 B.n139 71.676
R1278 B.n269 B.n140 71.676
R1279 B.n273 B.n141 71.676
R1280 B.n277 B.n142 71.676
R1281 B.n281 B.n143 71.676
R1282 B.n285 B.n144 71.676
R1283 B.n289 B.n145 71.676
R1284 B.n293 B.n146 71.676
R1285 B.n297 B.n147 71.676
R1286 B.n301 B.n148 71.676
R1287 B.n305 B.n149 71.676
R1288 B.n309 B.n150 71.676
R1289 B.n313 B.n151 71.676
R1290 B.n317 B.n152 71.676
R1291 B.n321 B.n153 71.676
R1292 B.n925 B.n154 71.676
R1293 B.n925 B.n924 71.676
R1294 B.n323 B.n153 71.676
R1295 B.n320 B.n152 71.676
R1296 B.n316 B.n151 71.676
R1297 B.n312 B.n150 71.676
R1298 B.n308 B.n149 71.676
R1299 B.n304 B.n148 71.676
R1300 B.n300 B.n147 71.676
R1301 B.n296 B.n146 71.676
R1302 B.n292 B.n145 71.676
R1303 B.n288 B.n144 71.676
R1304 B.n284 B.n143 71.676
R1305 B.n280 B.n142 71.676
R1306 B.n276 B.n141 71.676
R1307 B.n272 B.n140 71.676
R1308 B.n268 B.n139 71.676
R1309 B.n264 B.n138 71.676
R1310 B.n260 B.n137 71.676
R1311 B.n256 B.n136 71.676
R1312 B.n251 B.n135 71.676
R1313 B.n247 B.n134 71.676
R1314 B.n243 B.n133 71.676
R1315 B.n239 B.n132 71.676
R1316 B.n235 B.n131 71.676
R1317 B.n230 B.n130 71.676
R1318 B.n226 B.n129 71.676
R1319 B.n222 B.n128 71.676
R1320 B.n218 B.n127 71.676
R1321 B.n214 B.n126 71.676
R1322 B.n210 B.n125 71.676
R1323 B.n206 B.n124 71.676
R1324 B.n202 B.n123 71.676
R1325 B.n198 B.n122 71.676
R1326 B.n194 B.n121 71.676
R1327 B.n190 B.n120 71.676
R1328 B.n186 B.n119 71.676
R1329 B.n182 B.n118 71.676
R1330 B.n178 B.n117 71.676
R1331 B.n174 B.n116 71.676
R1332 B.n170 B.n115 71.676
R1333 B.n166 B.n114 71.676
R1334 B.n162 B.n113 71.676
R1335 B.n656 B.n655 71.676
R1336 B.n650 B.n446 71.676
R1337 B.n647 B.n447 71.676
R1338 B.n643 B.n448 71.676
R1339 B.n639 B.n449 71.676
R1340 B.n635 B.n450 71.676
R1341 B.n631 B.n451 71.676
R1342 B.n627 B.n452 71.676
R1343 B.n623 B.n453 71.676
R1344 B.n619 B.n454 71.676
R1345 B.n615 B.n455 71.676
R1346 B.n611 B.n456 71.676
R1347 B.n607 B.n457 71.676
R1348 B.n603 B.n458 71.676
R1349 B.n599 B.n459 71.676
R1350 B.n595 B.n460 71.676
R1351 B.n591 B.n461 71.676
R1352 B.n587 B.n462 71.676
R1353 B.n583 B.n463 71.676
R1354 B.n579 B.n464 71.676
R1355 B.n575 B.n465 71.676
R1356 B.n571 B.n466 71.676
R1357 B.n567 B.n467 71.676
R1358 B.n563 B.n468 71.676
R1359 B.n559 B.n469 71.676
R1360 B.n555 B.n470 71.676
R1361 B.n551 B.n471 71.676
R1362 B.n547 B.n472 71.676
R1363 B.n543 B.n473 71.676
R1364 B.n539 B.n474 71.676
R1365 B.n535 B.n475 71.676
R1366 B.n531 B.n476 71.676
R1367 B.n527 B.n477 71.676
R1368 B.n523 B.n478 71.676
R1369 B.n519 B.n479 71.676
R1370 B.n515 B.n480 71.676
R1371 B.n511 B.n481 71.676
R1372 B.n507 B.n482 71.676
R1373 B.n503 B.n483 71.676
R1374 B.n499 B.n484 71.676
R1375 B.n495 B.n485 71.676
R1376 B.n656 B.n487 71.676
R1377 B.n648 B.n446 71.676
R1378 B.n644 B.n447 71.676
R1379 B.n640 B.n448 71.676
R1380 B.n636 B.n449 71.676
R1381 B.n632 B.n450 71.676
R1382 B.n628 B.n451 71.676
R1383 B.n624 B.n452 71.676
R1384 B.n620 B.n453 71.676
R1385 B.n616 B.n454 71.676
R1386 B.n612 B.n455 71.676
R1387 B.n608 B.n456 71.676
R1388 B.n604 B.n457 71.676
R1389 B.n600 B.n458 71.676
R1390 B.n596 B.n459 71.676
R1391 B.n592 B.n460 71.676
R1392 B.n588 B.n461 71.676
R1393 B.n584 B.n462 71.676
R1394 B.n580 B.n463 71.676
R1395 B.n576 B.n464 71.676
R1396 B.n572 B.n465 71.676
R1397 B.n568 B.n466 71.676
R1398 B.n564 B.n467 71.676
R1399 B.n560 B.n468 71.676
R1400 B.n556 B.n469 71.676
R1401 B.n552 B.n470 71.676
R1402 B.n548 B.n471 71.676
R1403 B.n544 B.n472 71.676
R1404 B.n540 B.n473 71.676
R1405 B.n536 B.n474 71.676
R1406 B.n532 B.n475 71.676
R1407 B.n528 B.n476 71.676
R1408 B.n524 B.n477 71.676
R1409 B.n520 B.n478 71.676
R1410 B.n516 B.n479 71.676
R1411 B.n512 B.n480 71.676
R1412 B.n508 B.n481 71.676
R1413 B.n504 B.n482 71.676
R1414 B.n500 B.n483 71.676
R1415 B.n496 B.n484 71.676
R1416 B.n485 B.n445 71.676
R1417 B.n1051 B.n1050 71.676
R1418 B.n1051 B.n2 71.676
R1419 B.n158 B.n157 70.2066
R1420 B.n156 B.n155 70.2066
R1421 B.n492 B.n491 70.2066
R1422 B.n489 B.n488 70.2066
R1423 B.n233 B.n158 59.5399
R1424 B.n254 B.n156 59.5399
R1425 B.n493 B.n492 59.5399
R1426 B.n490 B.n489 59.5399
R1427 B.n663 B.n442 47.5681
R1428 B.n663 B.n438 47.5681
R1429 B.n669 B.n438 47.5681
R1430 B.n669 B.n434 47.5681
R1431 B.n675 B.n434 47.5681
R1432 B.n675 B.n429 47.5681
R1433 B.n681 B.n429 47.5681
R1434 B.n681 B.n430 47.5681
R1435 B.n687 B.n422 47.5681
R1436 B.n693 B.n422 47.5681
R1437 B.n693 B.n418 47.5681
R1438 B.n699 B.n418 47.5681
R1439 B.n699 B.n414 47.5681
R1440 B.n705 B.n414 47.5681
R1441 B.n705 B.n410 47.5681
R1442 B.n711 B.n410 47.5681
R1443 B.n711 B.n406 47.5681
R1444 B.n717 B.n406 47.5681
R1445 B.n717 B.n402 47.5681
R1446 B.n724 B.n402 47.5681
R1447 B.n724 B.n723 47.5681
R1448 B.n730 B.n395 47.5681
R1449 B.n736 B.n395 47.5681
R1450 B.n736 B.n391 47.5681
R1451 B.n742 B.n391 47.5681
R1452 B.n742 B.n387 47.5681
R1453 B.n748 B.n387 47.5681
R1454 B.n748 B.n383 47.5681
R1455 B.n754 B.n383 47.5681
R1456 B.n754 B.n379 47.5681
R1457 B.n760 B.n379 47.5681
R1458 B.n766 B.n375 47.5681
R1459 B.n766 B.n371 47.5681
R1460 B.n772 B.n371 47.5681
R1461 B.n772 B.n367 47.5681
R1462 B.n778 B.n367 47.5681
R1463 B.n778 B.n363 47.5681
R1464 B.n784 B.n363 47.5681
R1465 B.n784 B.n359 47.5681
R1466 B.n790 B.n359 47.5681
R1467 B.n796 B.n355 47.5681
R1468 B.n796 B.n351 47.5681
R1469 B.n802 B.n351 47.5681
R1470 B.n802 B.n347 47.5681
R1471 B.n808 B.n347 47.5681
R1472 B.n808 B.n343 47.5681
R1473 B.n814 B.n343 47.5681
R1474 B.n814 B.n339 47.5681
R1475 B.n821 B.n339 47.5681
R1476 B.n821 B.n820 47.5681
R1477 B.n827 B.n332 47.5681
R1478 B.n834 B.n332 47.5681
R1479 B.n834 B.n328 47.5681
R1480 B.n840 B.n328 47.5681
R1481 B.n840 B.n4 47.5681
R1482 B.n1049 B.n4 47.5681
R1483 B.n1049 B.n1048 47.5681
R1484 B.n1048 B.n1047 47.5681
R1485 B.n1047 B.n8 47.5681
R1486 B.n12 B.n8 47.5681
R1487 B.n1040 B.n12 47.5681
R1488 B.n1040 B.n1039 47.5681
R1489 B.n1039 B.n1038 47.5681
R1490 B.n1032 B.n19 47.5681
R1491 B.n1032 B.n1031 47.5681
R1492 B.n1031 B.n1030 47.5681
R1493 B.n1030 B.n23 47.5681
R1494 B.n1024 B.n23 47.5681
R1495 B.n1024 B.n1023 47.5681
R1496 B.n1023 B.n1022 47.5681
R1497 B.n1022 B.n30 47.5681
R1498 B.n1016 B.n30 47.5681
R1499 B.n1016 B.n1015 47.5681
R1500 B.n1014 B.n37 47.5681
R1501 B.n1008 B.n37 47.5681
R1502 B.n1008 B.n1007 47.5681
R1503 B.n1007 B.n1006 47.5681
R1504 B.n1006 B.n44 47.5681
R1505 B.n1000 B.n44 47.5681
R1506 B.n1000 B.n999 47.5681
R1507 B.n999 B.n998 47.5681
R1508 B.n998 B.n51 47.5681
R1509 B.n992 B.n991 47.5681
R1510 B.n991 B.n990 47.5681
R1511 B.n990 B.n58 47.5681
R1512 B.n984 B.n58 47.5681
R1513 B.n984 B.n983 47.5681
R1514 B.n983 B.n982 47.5681
R1515 B.n982 B.n65 47.5681
R1516 B.n976 B.n65 47.5681
R1517 B.n976 B.n975 47.5681
R1518 B.n975 B.n974 47.5681
R1519 B.n968 B.n75 47.5681
R1520 B.n968 B.n967 47.5681
R1521 B.n967 B.n966 47.5681
R1522 B.n966 B.n79 47.5681
R1523 B.n960 B.n79 47.5681
R1524 B.n960 B.n959 47.5681
R1525 B.n959 B.n958 47.5681
R1526 B.n958 B.n86 47.5681
R1527 B.n952 B.n86 47.5681
R1528 B.n952 B.n951 47.5681
R1529 B.n951 B.n950 47.5681
R1530 B.n950 B.n93 47.5681
R1531 B.n944 B.n93 47.5681
R1532 B.n943 B.n942 47.5681
R1533 B.n942 B.n100 47.5681
R1534 B.n936 B.n100 47.5681
R1535 B.n936 B.n935 47.5681
R1536 B.n935 B.n934 47.5681
R1537 B.n934 B.n107 47.5681
R1538 B.n928 B.n107 47.5681
R1539 B.n928 B.n927 47.5681
R1540 B.n790 B.t4 44.0705
R1541 B.t5 B.n1014 44.0705
R1542 B.n430 B.t16 37.0752
R1543 B.t9 B.n943 37.0752
R1544 B.t0 B.n375 34.2771
R1545 B.t6 B.n51 34.2771
R1546 B.n723 B.t2 30.08
R1547 B.n75 B.t3 30.08
R1548 B.n654 B.n440 29.1907
R1549 B.n660 B.n659 29.1907
R1550 B.n923 B.n922 29.1907
R1551 B.n160 B.n109 29.1907
R1552 B.n820 B.t1 27.2819
R1553 B.n19 B.t7 27.2819
R1554 B.n827 B.t1 20.2867
R1555 B.n1038 B.t7 20.2867
R1556 B B.n1052 18.0485
R1557 B.n730 B.t2 17.4886
R1558 B.n974 B.t3 17.4886
R1559 B.n760 B.t0 13.2914
R1560 B.n992 B.t6 13.2914
R1561 B.n665 B.n440 10.6151
R1562 B.n666 B.n665 10.6151
R1563 B.n667 B.n666 10.6151
R1564 B.n667 B.n432 10.6151
R1565 B.n677 B.n432 10.6151
R1566 B.n678 B.n677 10.6151
R1567 B.n679 B.n678 10.6151
R1568 B.n679 B.n424 10.6151
R1569 B.n689 B.n424 10.6151
R1570 B.n690 B.n689 10.6151
R1571 B.n691 B.n690 10.6151
R1572 B.n691 B.n416 10.6151
R1573 B.n701 B.n416 10.6151
R1574 B.n702 B.n701 10.6151
R1575 B.n703 B.n702 10.6151
R1576 B.n703 B.n408 10.6151
R1577 B.n713 B.n408 10.6151
R1578 B.n714 B.n713 10.6151
R1579 B.n715 B.n714 10.6151
R1580 B.n715 B.n400 10.6151
R1581 B.n726 B.n400 10.6151
R1582 B.n727 B.n726 10.6151
R1583 B.n728 B.n727 10.6151
R1584 B.n728 B.n393 10.6151
R1585 B.n738 B.n393 10.6151
R1586 B.n739 B.n738 10.6151
R1587 B.n740 B.n739 10.6151
R1588 B.n740 B.n385 10.6151
R1589 B.n750 B.n385 10.6151
R1590 B.n751 B.n750 10.6151
R1591 B.n752 B.n751 10.6151
R1592 B.n752 B.n377 10.6151
R1593 B.n762 B.n377 10.6151
R1594 B.n763 B.n762 10.6151
R1595 B.n764 B.n763 10.6151
R1596 B.n764 B.n369 10.6151
R1597 B.n774 B.n369 10.6151
R1598 B.n775 B.n774 10.6151
R1599 B.n776 B.n775 10.6151
R1600 B.n776 B.n361 10.6151
R1601 B.n786 B.n361 10.6151
R1602 B.n787 B.n786 10.6151
R1603 B.n788 B.n787 10.6151
R1604 B.n788 B.n353 10.6151
R1605 B.n798 B.n353 10.6151
R1606 B.n799 B.n798 10.6151
R1607 B.n800 B.n799 10.6151
R1608 B.n800 B.n345 10.6151
R1609 B.n810 B.n345 10.6151
R1610 B.n811 B.n810 10.6151
R1611 B.n812 B.n811 10.6151
R1612 B.n812 B.n337 10.6151
R1613 B.n823 B.n337 10.6151
R1614 B.n824 B.n823 10.6151
R1615 B.n825 B.n824 10.6151
R1616 B.n825 B.n330 10.6151
R1617 B.n836 B.n330 10.6151
R1618 B.n837 B.n836 10.6151
R1619 B.n838 B.n837 10.6151
R1620 B.n838 B.n0 10.6151
R1621 B.n654 B.n653 10.6151
R1622 B.n653 B.n652 10.6151
R1623 B.n652 B.n651 10.6151
R1624 B.n651 B.n649 10.6151
R1625 B.n649 B.n646 10.6151
R1626 B.n646 B.n645 10.6151
R1627 B.n645 B.n642 10.6151
R1628 B.n642 B.n641 10.6151
R1629 B.n641 B.n638 10.6151
R1630 B.n638 B.n637 10.6151
R1631 B.n637 B.n634 10.6151
R1632 B.n634 B.n633 10.6151
R1633 B.n633 B.n630 10.6151
R1634 B.n630 B.n629 10.6151
R1635 B.n629 B.n626 10.6151
R1636 B.n626 B.n625 10.6151
R1637 B.n625 B.n622 10.6151
R1638 B.n622 B.n621 10.6151
R1639 B.n621 B.n618 10.6151
R1640 B.n618 B.n617 10.6151
R1641 B.n617 B.n614 10.6151
R1642 B.n614 B.n613 10.6151
R1643 B.n613 B.n610 10.6151
R1644 B.n610 B.n609 10.6151
R1645 B.n609 B.n606 10.6151
R1646 B.n606 B.n605 10.6151
R1647 B.n605 B.n602 10.6151
R1648 B.n602 B.n601 10.6151
R1649 B.n601 B.n598 10.6151
R1650 B.n598 B.n597 10.6151
R1651 B.n597 B.n594 10.6151
R1652 B.n594 B.n593 10.6151
R1653 B.n593 B.n590 10.6151
R1654 B.n590 B.n589 10.6151
R1655 B.n589 B.n586 10.6151
R1656 B.n586 B.n585 10.6151
R1657 B.n582 B.n581 10.6151
R1658 B.n581 B.n578 10.6151
R1659 B.n578 B.n577 10.6151
R1660 B.n577 B.n574 10.6151
R1661 B.n574 B.n573 10.6151
R1662 B.n573 B.n570 10.6151
R1663 B.n570 B.n569 10.6151
R1664 B.n569 B.n566 10.6151
R1665 B.n566 B.n565 10.6151
R1666 B.n562 B.n561 10.6151
R1667 B.n561 B.n558 10.6151
R1668 B.n558 B.n557 10.6151
R1669 B.n557 B.n554 10.6151
R1670 B.n554 B.n553 10.6151
R1671 B.n553 B.n550 10.6151
R1672 B.n550 B.n549 10.6151
R1673 B.n549 B.n546 10.6151
R1674 B.n546 B.n545 10.6151
R1675 B.n545 B.n542 10.6151
R1676 B.n542 B.n541 10.6151
R1677 B.n541 B.n538 10.6151
R1678 B.n538 B.n537 10.6151
R1679 B.n537 B.n534 10.6151
R1680 B.n534 B.n533 10.6151
R1681 B.n533 B.n530 10.6151
R1682 B.n530 B.n529 10.6151
R1683 B.n529 B.n526 10.6151
R1684 B.n526 B.n525 10.6151
R1685 B.n525 B.n522 10.6151
R1686 B.n522 B.n521 10.6151
R1687 B.n521 B.n518 10.6151
R1688 B.n518 B.n517 10.6151
R1689 B.n517 B.n514 10.6151
R1690 B.n514 B.n513 10.6151
R1691 B.n513 B.n510 10.6151
R1692 B.n510 B.n509 10.6151
R1693 B.n509 B.n506 10.6151
R1694 B.n506 B.n505 10.6151
R1695 B.n505 B.n502 10.6151
R1696 B.n502 B.n501 10.6151
R1697 B.n501 B.n498 10.6151
R1698 B.n498 B.n497 10.6151
R1699 B.n497 B.n494 10.6151
R1700 B.n494 B.n444 10.6151
R1701 B.n659 B.n444 10.6151
R1702 B.n661 B.n660 10.6151
R1703 B.n661 B.n436 10.6151
R1704 B.n671 B.n436 10.6151
R1705 B.n672 B.n671 10.6151
R1706 B.n673 B.n672 10.6151
R1707 B.n673 B.n427 10.6151
R1708 B.n683 B.n427 10.6151
R1709 B.n684 B.n683 10.6151
R1710 B.n685 B.n684 10.6151
R1711 B.n685 B.n420 10.6151
R1712 B.n695 B.n420 10.6151
R1713 B.n696 B.n695 10.6151
R1714 B.n697 B.n696 10.6151
R1715 B.n697 B.n412 10.6151
R1716 B.n707 B.n412 10.6151
R1717 B.n708 B.n707 10.6151
R1718 B.n709 B.n708 10.6151
R1719 B.n709 B.n404 10.6151
R1720 B.n719 B.n404 10.6151
R1721 B.n720 B.n719 10.6151
R1722 B.n721 B.n720 10.6151
R1723 B.n721 B.n397 10.6151
R1724 B.n732 B.n397 10.6151
R1725 B.n733 B.n732 10.6151
R1726 B.n734 B.n733 10.6151
R1727 B.n734 B.n389 10.6151
R1728 B.n744 B.n389 10.6151
R1729 B.n745 B.n744 10.6151
R1730 B.n746 B.n745 10.6151
R1731 B.n746 B.n381 10.6151
R1732 B.n756 B.n381 10.6151
R1733 B.n757 B.n756 10.6151
R1734 B.n758 B.n757 10.6151
R1735 B.n758 B.n373 10.6151
R1736 B.n768 B.n373 10.6151
R1737 B.n769 B.n768 10.6151
R1738 B.n770 B.n769 10.6151
R1739 B.n770 B.n365 10.6151
R1740 B.n780 B.n365 10.6151
R1741 B.n781 B.n780 10.6151
R1742 B.n782 B.n781 10.6151
R1743 B.n782 B.n357 10.6151
R1744 B.n792 B.n357 10.6151
R1745 B.n793 B.n792 10.6151
R1746 B.n794 B.n793 10.6151
R1747 B.n794 B.n349 10.6151
R1748 B.n804 B.n349 10.6151
R1749 B.n805 B.n804 10.6151
R1750 B.n806 B.n805 10.6151
R1751 B.n806 B.n341 10.6151
R1752 B.n816 B.n341 10.6151
R1753 B.n817 B.n816 10.6151
R1754 B.n818 B.n817 10.6151
R1755 B.n818 B.n334 10.6151
R1756 B.n829 B.n334 10.6151
R1757 B.n830 B.n829 10.6151
R1758 B.n832 B.n830 10.6151
R1759 B.n832 B.n831 10.6151
R1760 B.n831 B.n326 10.6151
R1761 B.n843 B.n326 10.6151
R1762 B.n844 B.n843 10.6151
R1763 B.n845 B.n844 10.6151
R1764 B.n846 B.n845 10.6151
R1765 B.n847 B.n846 10.6151
R1766 B.n850 B.n847 10.6151
R1767 B.n851 B.n850 10.6151
R1768 B.n852 B.n851 10.6151
R1769 B.n853 B.n852 10.6151
R1770 B.n855 B.n853 10.6151
R1771 B.n856 B.n855 10.6151
R1772 B.n857 B.n856 10.6151
R1773 B.n858 B.n857 10.6151
R1774 B.n860 B.n858 10.6151
R1775 B.n861 B.n860 10.6151
R1776 B.n862 B.n861 10.6151
R1777 B.n863 B.n862 10.6151
R1778 B.n865 B.n863 10.6151
R1779 B.n866 B.n865 10.6151
R1780 B.n867 B.n866 10.6151
R1781 B.n868 B.n867 10.6151
R1782 B.n870 B.n868 10.6151
R1783 B.n871 B.n870 10.6151
R1784 B.n872 B.n871 10.6151
R1785 B.n873 B.n872 10.6151
R1786 B.n875 B.n873 10.6151
R1787 B.n876 B.n875 10.6151
R1788 B.n877 B.n876 10.6151
R1789 B.n878 B.n877 10.6151
R1790 B.n880 B.n878 10.6151
R1791 B.n881 B.n880 10.6151
R1792 B.n882 B.n881 10.6151
R1793 B.n883 B.n882 10.6151
R1794 B.n885 B.n883 10.6151
R1795 B.n886 B.n885 10.6151
R1796 B.n887 B.n886 10.6151
R1797 B.n888 B.n887 10.6151
R1798 B.n890 B.n888 10.6151
R1799 B.n891 B.n890 10.6151
R1800 B.n892 B.n891 10.6151
R1801 B.n893 B.n892 10.6151
R1802 B.n895 B.n893 10.6151
R1803 B.n896 B.n895 10.6151
R1804 B.n897 B.n896 10.6151
R1805 B.n898 B.n897 10.6151
R1806 B.n900 B.n898 10.6151
R1807 B.n901 B.n900 10.6151
R1808 B.n902 B.n901 10.6151
R1809 B.n903 B.n902 10.6151
R1810 B.n905 B.n903 10.6151
R1811 B.n906 B.n905 10.6151
R1812 B.n907 B.n906 10.6151
R1813 B.n908 B.n907 10.6151
R1814 B.n910 B.n908 10.6151
R1815 B.n911 B.n910 10.6151
R1816 B.n912 B.n911 10.6151
R1817 B.n913 B.n912 10.6151
R1818 B.n915 B.n913 10.6151
R1819 B.n916 B.n915 10.6151
R1820 B.n917 B.n916 10.6151
R1821 B.n918 B.n917 10.6151
R1822 B.n920 B.n918 10.6151
R1823 B.n921 B.n920 10.6151
R1824 B.n922 B.n921 10.6151
R1825 B.n1044 B.n1 10.6151
R1826 B.n1044 B.n1043 10.6151
R1827 B.n1043 B.n1042 10.6151
R1828 B.n1042 B.n10 10.6151
R1829 B.n1036 B.n10 10.6151
R1830 B.n1036 B.n1035 10.6151
R1831 B.n1035 B.n1034 10.6151
R1832 B.n1034 B.n17 10.6151
R1833 B.n1028 B.n17 10.6151
R1834 B.n1028 B.n1027 10.6151
R1835 B.n1027 B.n1026 10.6151
R1836 B.n1026 B.n25 10.6151
R1837 B.n1020 B.n25 10.6151
R1838 B.n1020 B.n1019 10.6151
R1839 B.n1019 B.n1018 10.6151
R1840 B.n1018 B.n32 10.6151
R1841 B.n1012 B.n32 10.6151
R1842 B.n1012 B.n1011 10.6151
R1843 B.n1011 B.n1010 10.6151
R1844 B.n1010 B.n39 10.6151
R1845 B.n1004 B.n39 10.6151
R1846 B.n1004 B.n1003 10.6151
R1847 B.n1003 B.n1002 10.6151
R1848 B.n1002 B.n46 10.6151
R1849 B.n996 B.n46 10.6151
R1850 B.n996 B.n995 10.6151
R1851 B.n995 B.n994 10.6151
R1852 B.n994 B.n53 10.6151
R1853 B.n988 B.n53 10.6151
R1854 B.n988 B.n987 10.6151
R1855 B.n987 B.n986 10.6151
R1856 B.n986 B.n60 10.6151
R1857 B.n980 B.n60 10.6151
R1858 B.n980 B.n979 10.6151
R1859 B.n979 B.n978 10.6151
R1860 B.n978 B.n67 10.6151
R1861 B.n972 B.n67 10.6151
R1862 B.n972 B.n971 10.6151
R1863 B.n971 B.n970 10.6151
R1864 B.n970 B.n73 10.6151
R1865 B.n964 B.n73 10.6151
R1866 B.n964 B.n963 10.6151
R1867 B.n963 B.n962 10.6151
R1868 B.n962 B.n81 10.6151
R1869 B.n956 B.n81 10.6151
R1870 B.n956 B.n955 10.6151
R1871 B.n955 B.n954 10.6151
R1872 B.n954 B.n88 10.6151
R1873 B.n948 B.n88 10.6151
R1874 B.n948 B.n947 10.6151
R1875 B.n947 B.n946 10.6151
R1876 B.n946 B.n95 10.6151
R1877 B.n940 B.n95 10.6151
R1878 B.n940 B.n939 10.6151
R1879 B.n939 B.n938 10.6151
R1880 B.n938 B.n102 10.6151
R1881 B.n932 B.n102 10.6151
R1882 B.n932 B.n931 10.6151
R1883 B.n931 B.n930 10.6151
R1884 B.n930 B.n109 10.6151
R1885 B.n161 B.n160 10.6151
R1886 B.n164 B.n161 10.6151
R1887 B.n165 B.n164 10.6151
R1888 B.n168 B.n165 10.6151
R1889 B.n169 B.n168 10.6151
R1890 B.n172 B.n169 10.6151
R1891 B.n173 B.n172 10.6151
R1892 B.n176 B.n173 10.6151
R1893 B.n177 B.n176 10.6151
R1894 B.n180 B.n177 10.6151
R1895 B.n181 B.n180 10.6151
R1896 B.n184 B.n181 10.6151
R1897 B.n185 B.n184 10.6151
R1898 B.n188 B.n185 10.6151
R1899 B.n189 B.n188 10.6151
R1900 B.n192 B.n189 10.6151
R1901 B.n193 B.n192 10.6151
R1902 B.n196 B.n193 10.6151
R1903 B.n197 B.n196 10.6151
R1904 B.n200 B.n197 10.6151
R1905 B.n201 B.n200 10.6151
R1906 B.n204 B.n201 10.6151
R1907 B.n205 B.n204 10.6151
R1908 B.n208 B.n205 10.6151
R1909 B.n209 B.n208 10.6151
R1910 B.n212 B.n209 10.6151
R1911 B.n213 B.n212 10.6151
R1912 B.n216 B.n213 10.6151
R1913 B.n217 B.n216 10.6151
R1914 B.n220 B.n217 10.6151
R1915 B.n221 B.n220 10.6151
R1916 B.n224 B.n221 10.6151
R1917 B.n225 B.n224 10.6151
R1918 B.n228 B.n225 10.6151
R1919 B.n229 B.n228 10.6151
R1920 B.n232 B.n229 10.6151
R1921 B.n237 B.n234 10.6151
R1922 B.n238 B.n237 10.6151
R1923 B.n241 B.n238 10.6151
R1924 B.n242 B.n241 10.6151
R1925 B.n245 B.n242 10.6151
R1926 B.n246 B.n245 10.6151
R1927 B.n249 B.n246 10.6151
R1928 B.n250 B.n249 10.6151
R1929 B.n253 B.n250 10.6151
R1930 B.n258 B.n255 10.6151
R1931 B.n259 B.n258 10.6151
R1932 B.n262 B.n259 10.6151
R1933 B.n263 B.n262 10.6151
R1934 B.n266 B.n263 10.6151
R1935 B.n267 B.n266 10.6151
R1936 B.n270 B.n267 10.6151
R1937 B.n271 B.n270 10.6151
R1938 B.n274 B.n271 10.6151
R1939 B.n275 B.n274 10.6151
R1940 B.n278 B.n275 10.6151
R1941 B.n279 B.n278 10.6151
R1942 B.n282 B.n279 10.6151
R1943 B.n283 B.n282 10.6151
R1944 B.n286 B.n283 10.6151
R1945 B.n287 B.n286 10.6151
R1946 B.n290 B.n287 10.6151
R1947 B.n291 B.n290 10.6151
R1948 B.n294 B.n291 10.6151
R1949 B.n295 B.n294 10.6151
R1950 B.n298 B.n295 10.6151
R1951 B.n299 B.n298 10.6151
R1952 B.n302 B.n299 10.6151
R1953 B.n303 B.n302 10.6151
R1954 B.n306 B.n303 10.6151
R1955 B.n307 B.n306 10.6151
R1956 B.n310 B.n307 10.6151
R1957 B.n311 B.n310 10.6151
R1958 B.n314 B.n311 10.6151
R1959 B.n315 B.n314 10.6151
R1960 B.n318 B.n315 10.6151
R1961 B.n319 B.n318 10.6151
R1962 B.n322 B.n319 10.6151
R1963 B.n324 B.n322 10.6151
R1964 B.n325 B.n324 10.6151
R1965 B.n923 B.n325 10.6151
R1966 B.n687 B.t16 10.4933
R1967 B.n944 B.t9 10.4933
R1968 B.n585 B.n490 9.36635
R1969 B.n562 B.n493 9.36635
R1970 B.n233 B.n232 9.36635
R1971 B.n255 B.n254 9.36635
R1972 B.n1052 B.n0 8.11757
R1973 B.n1052 B.n1 8.11757
R1974 B.t4 B.n355 3.49812
R1975 B.n1015 B.t5 3.49812
R1976 B.n582 B.n490 1.24928
R1977 B.n565 B.n493 1.24928
R1978 B.n234 B.n233 1.24928
R1979 B.n254 B.n253 1.24928
R1980 VP.n24 VP.n21 161.3
R1981 VP.n26 VP.n25 161.3
R1982 VP.n27 VP.n20 161.3
R1983 VP.n29 VP.n28 161.3
R1984 VP.n30 VP.n19 161.3
R1985 VP.n32 VP.n31 161.3
R1986 VP.n33 VP.n18 161.3
R1987 VP.n35 VP.n34 161.3
R1988 VP.n37 VP.n36 161.3
R1989 VP.n38 VP.n16 161.3
R1990 VP.n40 VP.n39 161.3
R1991 VP.n41 VP.n15 161.3
R1992 VP.n43 VP.n42 161.3
R1993 VP.n44 VP.n14 161.3
R1994 VP.n46 VP.n45 161.3
R1995 VP.n83 VP.n82 161.3
R1996 VP.n81 VP.n1 161.3
R1997 VP.n80 VP.n79 161.3
R1998 VP.n78 VP.n2 161.3
R1999 VP.n77 VP.n76 161.3
R2000 VP.n75 VP.n3 161.3
R2001 VP.n74 VP.n73 161.3
R2002 VP.n72 VP.n71 161.3
R2003 VP.n70 VP.n5 161.3
R2004 VP.n69 VP.n68 161.3
R2005 VP.n67 VP.n6 161.3
R2006 VP.n66 VP.n65 161.3
R2007 VP.n64 VP.n7 161.3
R2008 VP.n63 VP.n62 161.3
R2009 VP.n61 VP.n8 161.3
R2010 VP.n60 VP.n59 161.3
R2011 VP.n57 VP.n9 161.3
R2012 VP.n56 VP.n55 161.3
R2013 VP.n54 VP.n10 161.3
R2014 VP.n53 VP.n52 161.3
R2015 VP.n51 VP.n11 161.3
R2016 VP.n50 VP.n49 161.3
R2017 VP.n23 VP.t5 108.425
R2018 VP.n48 VP.n12 81.2593
R2019 VP.n84 VP.n0 81.2593
R2020 VP.n47 VP.n13 81.2593
R2021 VP.n12 VP.t6 76.5491
R2022 VP.n58 VP.t0 76.5491
R2023 VP.n4 VP.t4 76.5491
R2024 VP.n0 VP.t3 76.5491
R2025 VP.n13 VP.t1 76.5491
R2026 VP.n17 VP.t7 76.5491
R2027 VP.n22 VP.t2 76.5491
R2028 VP.n23 VP.n22 71.6409
R2029 VP.n65 VP.n6 56.5193
R2030 VP.n28 VP.n19 56.5193
R2031 VP.n56 VP.n10 53.1199
R2032 VP.n76 VP.n2 53.1199
R2033 VP.n39 VP.n15 53.1199
R2034 VP.n48 VP.n47 52.969
R2035 VP.n52 VP.n10 27.8669
R2036 VP.n80 VP.n2 27.8669
R2037 VP.n43 VP.n15 27.8669
R2038 VP.n51 VP.n50 24.4675
R2039 VP.n52 VP.n51 24.4675
R2040 VP.n57 VP.n56 24.4675
R2041 VP.n59 VP.n57 24.4675
R2042 VP.n63 VP.n8 24.4675
R2043 VP.n64 VP.n63 24.4675
R2044 VP.n65 VP.n64 24.4675
R2045 VP.n69 VP.n6 24.4675
R2046 VP.n70 VP.n69 24.4675
R2047 VP.n71 VP.n70 24.4675
R2048 VP.n75 VP.n74 24.4675
R2049 VP.n76 VP.n75 24.4675
R2050 VP.n81 VP.n80 24.4675
R2051 VP.n82 VP.n81 24.4675
R2052 VP.n44 VP.n43 24.4675
R2053 VP.n45 VP.n44 24.4675
R2054 VP.n32 VP.n19 24.4675
R2055 VP.n33 VP.n32 24.4675
R2056 VP.n34 VP.n33 24.4675
R2057 VP.n38 VP.n37 24.4675
R2058 VP.n39 VP.n38 24.4675
R2059 VP.n26 VP.n21 24.4675
R2060 VP.n27 VP.n26 24.4675
R2061 VP.n28 VP.n27 24.4675
R2062 VP.n59 VP.n58 21.5315
R2063 VP.n74 VP.n4 21.5315
R2064 VP.n37 VP.n17 21.5315
R2065 VP.n50 VP.n12 8.80862
R2066 VP.n82 VP.n0 8.80862
R2067 VP.n45 VP.n13 8.80862
R2068 VP.n24 VP.n23 4.46855
R2069 VP.n58 VP.n8 2.93654
R2070 VP.n71 VP.n4 2.93654
R2071 VP.n34 VP.n17 2.93654
R2072 VP.n22 VP.n21 2.93654
R2073 VP.n47 VP.n46 0.354971
R2074 VP.n49 VP.n48 0.354971
R2075 VP.n84 VP.n83 0.354971
R2076 VP VP.n84 0.26696
R2077 VP.n25 VP.n24 0.189894
R2078 VP.n25 VP.n20 0.189894
R2079 VP.n29 VP.n20 0.189894
R2080 VP.n30 VP.n29 0.189894
R2081 VP.n31 VP.n30 0.189894
R2082 VP.n31 VP.n18 0.189894
R2083 VP.n35 VP.n18 0.189894
R2084 VP.n36 VP.n35 0.189894
R2085 VP.n36 VP.n16 0.189894
R2086 VP.n40 VP.n16 0.189894
R2087 VP.n41 VP.n40 0.189894
R2088 VP.n42 VP.n41 0.189894
R2089 VP.n42 VP.n14 0.189894
R2090 VP.n46 VP.n14 0.189894
R2091 VP.n49 VP.n11 0.189894
R2092 VP.n53 VP.n11 0.189894
R2093 VP.n54 VP.n53 0.189894
R2094 VP.n55 VP.n54 0.189894
R2095 VP.n55 VP.n9 0.189894
R2096 VP.n60 VP.n9 0.189894
R2097 VP.n61 VP.n60 0.189894
R2098 VP.n62 VP.n61 0.189894
R2099 VP.n62 VP.n7 0.189894
R2100 VP.n66 VP.n7 0.189894
R2101 VP.n67 VP.n66 0.189894
R2102 VP.n68 VP.n67 0.189894
R2103 VP.n68 VP.n5 0.189894
R2104 VP.n72 VP.n5 0.189894
R2105 VP.n73 VP.n72 0.189894
R2106 VP.n73 VP.n3 0.189894
R2107 VP.n77 VP.n3 0.189894
R2108 VP.n78 VP.n77 0.189894
R2109 VP.n79 VP.n78 0.189894
R2110 VP.n79 VP.n1 0.189894
R2111 VP.n83 VP.n1 0.189894
R2112 VDD1 VDD1.n0 66.6227
R2113 VDD1.n3 VDD1.n2 66.509
R2114 VDD1.n3 VDD1.n1 66.509
R2115 VDD1.n5 VDD1.n4 65.004
R2116 VDD1.n5 VDD1.n3 47.35
R2117 VDD1.n4 VDD1.t0 1.89524
R2118 VDD1.n4 VDD1.t6 1.89524
R2119 VDD1.n0 VDD1.t2 1.89524
R2120 VDD1.n0 VDD1.t5 1.89524
R2121 VDD1.n2 VDD1.t3 1.89524
R2122 VDD1.n2 VDD1.t4 1.89524
R2123 VDD1.n1 VDD1.t1 1.89524
R2124 VDD1.n1 VDD1.t7 1.89524
R2125 VDD1 VDD1.n5 1.50266
C0 VDD2 VN 7.9499f
C1 VP VN 8.22459f
C2 VTAIL VN 8.64771f
C3 VP VDD2 0.593083f
C4 VN VDD1 0.152964f
C5 VTAIL VDD2 7.9184f
C6 VTAIL VP 8.661819f
C7 VDD2 VDD1 2.13412f
C8 VP VDD1 8.388269f
C9 VTAIL VDD1 7.85935f
C10 VDD2 B 5.984487f
C11 VDD1 B 6.504629f
C12 VTAIL B 10.024788f
C13 VN B 18.050268f
C14 VP B 16.709137f
C15 VDD1.t2 B 0.229504f
C16 VDD1.t5 B 0.229504f
C17 VDD1.n0 B 2.04542f
C18 VDD1.t1 B 0.229504f
C19 VDD1.t7 B 0.229504f
C20 VDD1.n1 B 2.0441f
C21 VDD1.t3 B 0.229504f
C22 VDD1.t4 B 0.229504f
C23 VDD1.n2 B 2.0441f
C24 VDD1.n3 B 4.03121f
C25 VDD1.t0 B 0.229504f
C26 VDD1.t6 B 0.229504f
C27 VDD1.n4 B 2.02936f
C28 VDD1.n5 B 3.44565f
C29 VP.t3 B 1.84992f
C30 VP.n0 B 0.726168f
C31 VP.n1 B 0.019833f
C32 VP.n2 B 0.020801f
C33 VP.n3 B 0.019833f
C34 VP.t4 B 1.84992f
C35 VP.n4 B 0.655208f
C36 VP.n5 B 0.019833f
C37 VP.n6 B 0.028952f
C38 VP.n7 B 0.019833f
C39 VP.n8 B 0.020904f
C40 VP.n9 B 0.019833f
C41 VP.n10 B 0.020801f
C42 VP.n11 B 0.019833f
C43 VP.t6 B 1.84992f
C44 VP.n12 B 0.726168f
C45 VP.t1 B 1.84992f
C46 VP.n13 B 0.726168f
C47 VP.n14 B 0.019833f
C48 VP.n15 B 0.020801f
C49 VP.n16 B 0.019833f
C50 VP.t7 B 1.84992f
C51 VP.n17 B 0.655208f
C52 VP.n18 B 0.019833f
C53 VP.n19 B 0.028952f
C54 VP.n20 B 0.019833f
C55 VP.n21 B 0.020904f
C56 VP.t5 B 2.08301f
C57 VP.t2 B 1.84992f
C58 VP.n22 B 0.715465f
C59 VP.n23 B 0.686079f
C60 VP.n24 B 0.234423f
C61 VP.n25 B 0.019833f
C62 VP.n26 B 0.036963f
C63 VP.n27 B 0.036963f
C64 VP.n28 B 0.028952f
C65 VP.n29 B 0.019833f
C66 VP.n30 B 0.019833f
C67 VP.n31 B 0.019833f
C68 VP.n32 B 0.036963f
C69 VP.n33 B 0.036963f
C70 VP.n34 B 0.020904f
C71 VP.n35 B 0.019833f
C72 VP.n36 B 0.019833f
C73 VP.n37 B 0.034773f
C74 VP.n38 B 0.036963f
C75 VP.n39 B 0.035189f
C76 VP.n40 B 0.019833f
C77 VP.n41 B 0.019833f
C78 VP.n42 B 0.019833f
C79 VP.n43 B 0.038876f
C80 VP.n44 B 0.036963f
C81 VP.n45 B 0.025284f
C82 VP.n46 B 0.032009f
C83 VP.n47 B 1.2269f
C84 VP.n48 B 1.24036f
C85 VP.n49 B 0.032009f
C86 VP.n50 B 0.025284f
C87 VP.n51 B 0.036963f
C88 VP.n52 B 0.038876f
C89 VP.n53 B 0.019833f
C90 VP.n54 B 0.019833f
C91 VP.n55 B 0.019833f
C92 VP.n56 B 0.035189f
C93 VP.n57 B 0.036963f
C94 VP.t0 B 1.84992f
C95 VP.n58 B 0.655208f
C96 VP.n59 B 0.034773f
C97 VP.n60 B 0.019833f
C98 VP.n61 B 0.019833f
C99 VP.n62 B 0.019833f
C100 VP.n63 B 0.036963f
C101 VP.n64 B 0.036963f
C102 VP.n65 B 0.028952f
C103 VP.n66 B 0.019833f
C104 VP.n67 B 0.019833f
C105 VP.n68 B 0.019833f
C106 VP.n69 B 0.036963f
C107 VP.n70 B 0.036963f
C108 VP.n71 B 0.020904f
C109 VP.n72 B 0.019833f
C110 VP.n73 B 0.019833f
C111 VP.n74 B 0.034773f
C112 VP.n75 B 0.036963f
C113 VP.n76 B 0.035189f
C114 VP.n77 B 0.019833f
C115 VP.n78 B 0.019833f
C116 VP.n79 B 0.019833f
C117 VP.n80 B 0.038876f
C118 VP.n81 B 0.036963f
C119 VP.n82 B 0.025284f
C120 VP.n83 B 0.032009f
C121 VP.n84 B 0.05205f
C122 VTAIL.t8 B 0.172891f
C123 VTAIL.t13 B 0.172891f
C124 VTAIL.n0 B 1.47162f
C125 VTAIL.n1 B 0.412739f
C126 VTAIL.t14 B 1.87635f
C127 VTAIL.n2 B 0.507299f
C128 VTAIL.t1 B 1.87635f
C129 VTAIL.n3 B 0.507299f
C130 VTAIL.t0 B 0.172891f
C131 VTAIL.t4 B 0.172891f
C132 VTAIL.n4 B 1.47162f
C133 VTAIL.n5 B 0.619341f
C134 VTAIL.t2 B 1.87635f
C135 VTAIL.n6 B 1.57827f
C136 VTAIL.t15 B 1.87635f
C137 VTAIL.n7 B 1.57826f
C138 VTAIL.t10 B 0.172891f
C139 VTAIL.t11 B 0.172891f
C140 VTAIL.n8 B 1.47162f
C141 VTAIL.n9 B 0.619337f
C142 VTAIL.t12 B 1.87635f
C143 VTAIL.n10 B 0.507294f
C144 VTAIL.t7 B 1.87635f
C145 VTAIL.n11 B 0.507294f
C146 VTAIL.t5 B 0.172891f
C147 VTAIL.t6 B 0.172891f
C148 VTAIL.n12 B 1.47162f
C149 VTAIL.n13 B 0.619337f
C150 VTAIL.t3 B 1.87635f
C151 VTAIL.n14 B 1.57827f
C152 VTAIL.t9 B 1.87635f
C153 VTAIL.n15 B 1.57434f
C154 VDD2.t7 B 0.22452f
C155 VDD2.t0 B 0.22452f
C156 VDD2.n0 B 1.99971f
C157 VDD2.t1 B 0.22452f
C158 VDD2.t5 B 0.22452f
C159 VDD2.n1 B 1.99971f
C160 VDD2.n2 B 3.88738f
C161 VDD2.t6 B 0.22452f
C162 VDD2.t4 B 0.22452f
C163 VDD2.n3 B 1.9853f
C164 VDD2.n4 B 3.33687f
C165 VDD2.t3 B 0.22452f
C166 VDD2.t2 B 0.22452f
C167 VDD2.n5 B 1.99966f
C168 VN.t6 B 1.80406f
C169 VN.n0 B 0.708167f
C170 VN.n1 B 0.019341f
C171 VN.n2 B 0.020286f
C172 VN.n3 B 0.019341f
C173 VN.t2 B 1.80406f
C174 VN.n4 B 0.638965f
C175 VN.n5 B 0.019341f
C176 VN.n6 B 0.028234f
C177 VN.n7 B 0.019341f
C178 VN.n8 B 0.020386f
C179 VN.t7 B 1.80406f
C180 VN.n9 B 0.697729f
C181 VN.t1 B 2.03137f
C182 VN.n10 B 0.66907f
C183 VN.n11 B 0.228612f
C184 VN.n12 B 0.019341f
C185 VN.n13 B 0.036047f
C186 VN.n14 B 0.036047f
C187 VN.n15 B 0.028234f
C188 VN.n16 B 0.019341f
C189 VN.n17 B 0.019341f
C190 VN.n18 B 0.019341f
C191 VN.n19 B 0.036047f
C192 VN.n20 B 0.036047f
C193 VN.n21 B 0.020386f
C194 VN.n22 B 0.019341f
C195 VN.n23 B 0.019341f
C196 VN.n24 B 0.033911f
C197 VN.n25 B 0.036047f
C198 VN.n26 B 0.034317f
C199 VN.n27 B 0.019341f
C200 VN.n28 B 0.019341f
C201 VN.n29 B 0.019341f
C202 VN.n30 B 0.037913f
C203 VN.n31 B 0.036047f
C204 VN.n32 B 0.024657f
C205 VN.n33 B 0.031216f
C206 VN.n34 B 0.05076f
C207 VN.t0 B 1.80406f
C208 VN.n35 B 0.708167f
C209 VN.n36 B 0.019341f
C210 VN.n37 B 0.020286f
C211 VN.n38 B 0.019341f
C212 VN.t5 B 1.80406f
C213 VN.n39 B 0.638965f
C214 VN.n40 B 0.019341f
C215 VN.n41 B 0.028234f
C216 VN.n42 B 0.019341f
C217 VN.n43 B 0.020386f
C218 VN.t3 B 2.03137f
C219 VN.t4 B 1.80406f
C220 VN.n44 B 0.697729f
C221 VN.n45 B 0.66907f
C222 VN.n46 B 0.228612f
C223 VN.n47 B 0.019341f
C224 VN.n48 B 0.036047f
C225 VN.n49 B 0.036047f
C226 VN.n50 B 0.028234f
C227 VN.n51 B 0.019341f
C228 VN.n52 B 0.019341f
C229 VN.n53 B 0.019341f
C230 VN.n54 B 0.036047f
C231 VN.n55 B 0.036047f
C232 VN.n56 B 0.020386f
C233 VN.n57 B 0.019341f
C234 VN.n58 B 0.019341f
C235 VN.n59 B 0.033911f
C236 VN.n60 B 0.036047f
C237 VN.n61 B 0.034317f
C238 VN.n62 B 0.019341f
C239 VN.n63 B 0.019341f
C240 VN.n64 B 0.019341f
C241 VN.n65 B 0.037913f
C242 VN.n66 B 0.036047f
C243 VN.n67 B 0.024657f
C244 VN.n68 B 0.031216f
C245 VN.n69 B 1.20425f
.ends

