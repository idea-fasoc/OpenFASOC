* NGSPICE file created from diff_pair_sample_0638.ext - technology: sky130A

.subckt diff_pair_sample_0638 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=0.9372 ps=6.01 w=5.68 l=3.26
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=2.2152 ps=12.14 w=5.68 l=3.26
X2 VDD1.t3 VP.t2 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0.9372 ps=6.01 w=5.68 l=3.26
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=3.26
X4 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=2.2152 ps=12.14 w=5.68 l=3.26
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=3.26
X6 VTAIL.t8 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=0.9372 ps=6.01 w=5.68 l=3.26
X7 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=2.2152 ps=12.14 w=5.68 l=3.26
X8 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=3.26
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=3.26
X10 VTAIL.t2 VN.t2 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=0.9372 ps=6.01 w=5.68 l=3.26
X11 VTAIL.t1 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=0.9372 ps=6.01 w=5.68 l=3.26
X12 VDD1.t5 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0.9372 ps=6.01 w=5.68 l=3.26
X13 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0.9372 ps=6.01 w=5.68 l=3.26
X14 VDD1.t1 VP.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9372 pd=6.01 as=2.2152 ps=12.14 w=5.68 l=3.26
X15 VDD2.t0 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2152 pd=12.14 as=0.9372 ps=6.01 w=5.68 l=3.26
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t4 75.2139
R22 VP.n27 VP.n8 73.5231
R23 VP.n50 VP.n0 73.5231
R24 VP.n26 VP.n9 73.5231
R25 VP.n14 VP.n13 62.2205
R26 VP.n27 VP.n26 46.6094
R27 VP.n31 VP.n6 44.9365
R28 VP.n46 VP.n2 44.9365
R29 VP.n22 VP.n11 44.9365
R30 VP.n8 VP.t2 41.9907
R31 VP.n4 VP.t3 41.9907
R32 VP.n0 VP.t1 41.9907
R33 VP.n9 VP.t5 41.9907
R34 VP.n13 VP.t0 41.9907
R35 VP.n35 VP.n6 36.2176
R36 VP.n42 VP.n2 36.2176
R37 VP.n18 VP.n11 36.2176
R38 VP.n30 VP.n29 24.5923
R39 VP.n31 VP.n30 24.5923
R40 VP.n36 VP.n35 24.5923
R41 VP.n37 VP.n36 24.5923
R42 VP.n41 VP.n40 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n47 VP.n46 24.5923
R45 VP.n48 VP.n47 24.5923
R46 VP.n23 VP.n22 24.5923
R47 VP.n24 VP.n23 24.5923
R48 VP.n17 VP.n16 24.5923
R49 VP.n18 VP.n17 24.5923
R50 VP.n29 VP.n8 16.7229
R51 VP.n48 VP.n0 16.7229
R52 VP.n24 VP.n9 16.7229
R53 VP.n37 VP.n4 12.2964
R54 VP.n40 VP.n4 12.2964
R55 VP.n16 VP.n13 12.2964
R56 VP.n15 VP.n14 4.04952
R57 VP.n26 VP.n25 0.354861
R58 VP.n28 VP.n27 0.354861
R59 VP.n50 VP.n49 0.354861
R60 VP VP.n50 0.267071
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VDD1 VDD1.t5 74.511
R81 VDD1.n1 VDD1.t3 74.3973
R82 VDD1.n1 VDD1.n0 69.3639
R83 VDD1.n3 VDD1.n2 68.6456
R84 VDD1.n3 VDD1.n1 40.8005
R85 VDD1.n2 VDD1.t2 3.48642
R86 VDD1.n2 VDD1.t1 3.48642
R87 VDD1.n0 VDD1.t0 3.48642
R88 VDD1.n0 VDD1.t4 3.48642
R89 VDD1 VDD1.n3 0.716017
R90 VTAIL.n7 VTAIL.t3 55.4529
R91 VTAIL.n11 VTAIL.t4 55.4527
R92 VTAIL.n2 VTAIL.t10 55.4527
R93 VTAIL.n10 VTAIL.t6 55.4527
R94 VTAIL.n9 VTAIL.n8 51.967
R95 VTAIL.n6 VTAIL.n5 51.967
R96 VTAIL.n1 VTAIL.n0 51.9668
R97 VTAIL.n4 VTAIL.n3 51.9668
R98 VTAIL.n6 VTAIL.n4 23.4531
R99 VTAIL.n11 VTAIL.n10 20.3583
R100 VTAIL.n0 VTAIL.t5 3.48642
R101 VTAIL.n0 VTAIL.t1 3.48642
R102 VTAIL.n3 VTAIL.t9 3.48642
R103 VTAIL.n3 VTAIL.t8 3.48642
R104 VTAIL.n8 VTAIL.t7 3.48642
R105 VTAIL.n8 VTAIL.t11 3.48642
R106 VTAIL.n5 VTAIL.t0 3.48642
R107 VTAIL.n5 VTAIL.t2 3.48642
R108 VTAIL.n7 VTAIL.n6 3.09533
R109 VTAIL.n10 VTAIL.n9 3.09533
R110 VTAIL.n4 VTAIL.n2 3.09533
R111 VTAIL VTAIL.n11 2.26343
R112 VTAIL.n9 VTAIL.n7 2.01774
R113 VTAIL.n2 VTAIL.n1 2.01774
R114 VTAIL VTAIL.n1 0.832397
R115 B.n586 B.n585 585
R116 B.n588 B.n126 585
R117 B.n591 B.n590 585
R118 B.n592 B.n125 585
R119 B.n594 B.n593 585
R120 B.n596 B.n124 585
R121 B.n599 B.n598 585
R122 B.n600 B.n123 585
R123 B.n602 B.n601 585
R124 B.n604 B.n122 585
R125 B.n607 B.n606 585
R126 B.n608 B.n121 585
R127 B.n610 B.n609 585
R128 B.n612 B.n120 585
R129 B.n615 B.n614 585
R130 B.n616 B.n119 585
R131 B.n618 B.n617 585
R132 B.n620 B.n118 585
R133 B.n623 B.n622 585
R134 B.n624 B.n117 585
R135 B.n626 B.n625 585
R136 B.n628 B.n116 585
R137 B.n631 B.n630 585
R138 B.n633 B.n113 585
R139 B.n635 B.n634 585
R140 B.n637 B.n112 585
R141 B.n640 B.n639 585
R142 B.n641 B.n111 585
R143 B.n643 B.n642 585
R144 B.n645 B.n110 585
R145 B.n648 B.n647 585
R146 B.n649 B.n106 585
R147 B.n651 B.n650 585
R148 B.n653 B.n105 585
R149 B.n656 B.n655 585
R150 B.n657 B.n104 585
R151 B.n659 B.n658 585
R152 B.n661 B.n103 585
R153 B.n664 B.n663 585
R154 B.n665 B.n102 585
R155 B.n667 B.n666 585
R156 B.n669 B.n101 585
R157 B.n672 B.n671 585
R158 B.n673 B.n100 585
R159 B.n675 B.n674 585
R160 B.n677 B.n99 585
R161 B.n680 B.n679 585
R162 B.n681 B.n98 585
R163 B.n683 B.n682 585
R164 B.n685 B.n97 585
R165 B.n688 B.n687 585
R166 B.n689 B.n96 585
R167 B.n691 B.n690 585
R168 B.n693 B.n95 585
R169 B.n696 B.n695 585
R170 B.n697 B.n94 585
R171 B.n584 B.n92 585
R172 B.n700 B.n92 585
R173 B.n583 B.n91 585
R174 B.n701 B.n91 585
R175 B.n582 B.n90 585
R176 B.n702 B.n90 585
R177 B.n581 B.n580 585
R178 B.n580 B.n86 585
R179 B.n579 B.n85 585
R180 B.n708 B.n85 585
R181 B.n578 B.n84 585
R182 B.n709 B.n84 585
R183 B.n577 B.n83 585
R184 B.n710 B.n83 585
R185 B.n576 B.n575 585
R186 B.n575 B.n79 585
R187 B.n574 B.n78 585
R188 B.n716 B.n78 585
R189 B.n573 B.n77 585
R190 B.n717 B.n77 585
R191 B.n572 B.n76 585
R192 B.n718 B.n76 585
R193 B.n571 B.n570 585
R194 B.n570 B.n72 585
R195 B.n569 B.n71 585
R196 B.n724 B.n71 585
R197 B.n568 B.n70 585
R198 B.n725 B.n70 585
R199 B.n567 B.n69 585
R200 B.n726 B.n69 585
R201 B.n566 B.n565 585
R202 B.n565 B.n65 585
R203 B.n564 B.n64 585
R204 B.n732 B.n64 585
R205 B.n563 B.n63 585
R206 B.n733 B.n63 585
R207 B.n562 B.n62 585
R208 B.n734 B.n62 585
R209 B.n561 B.n560 585
R210 B.n560 B.n58 585
R211 B.n559 B.n57 585
R212 B.n740 B.n57 585
R213 B.n558 B.n56 585
R214 B.n741 B.n56 585
R215 B.n557 B.n55 585
R216 B.n742 B.n55 585
R217 B.n556 B.n555 585
R218 B.n555 B.n51 585
R219 B.n554 B.n50 585
R220 B.n748 B.n50 585
R221 B.n553 B.n49 585
R222 B.n749 B.n49 585
R223 B.n552 B.n48 585
R224 B.n750 B.n48 585
R225 B.n551 B.n550 585
R226 B.n550 B.n44 585
R227 B.n549 B.n43 585
R228 B.n756 B.n43 585
R229 B.n548 B.n42 585
R230 B.n757 B.n42 585
R231 B.n547 B.n41 585
R232 B.n758 B.n41 585
R233 B.n546 B.n545 585
R234 B.n545 B.n37 585
R235 B.n544 B.n36 585
R236 B.n764 B.n36 585
R237 B.n543 B.n35 585
R238 B.n765 B.n35 585
R239 B.n542 B.n34 585
R240 B.n766 B.n34 585
R241 B.n541 B.n540 585
R242 B.n540 B.n30 585
R243 B.n539 B.n29 585
R244 B.n772 B.n29 585
R245 B.n538 B.n28 585
R246 B.n773 B.n28 585
R247 B.n537 B.n27 585
R248 B.n774 B.n27 585
R249 B.n536 B.n535 585
R250 B.n535 B.n23 585
R251 B.n534 B.n22 585
R252 B.n780 B.n22 585
R253 B.n533 B.n21 585
R254 B.n781 B.n21 585
R255 B.n532 B.n20 585
R256 B.n782 B.n20 585
R257 B.n531 B.n530 585
R258 B.n530 B.n19 585
R259 B.n529 B.n15 585
R260 B.n788 B.n15 585
R261 B.n528 B.n14 585
R262 B.n789 B.n14 585
R263 B.n527 B.n13 585
R264 B.n790 B.n13 585
R265 B.n526 B.n525 585
R266 B.n525 B.n12 585
R267 B.n524 B.n523 585
R268 B.n524 B.n8 585
R269 B.n522 B.n7 585
R270 B.n797 B.n7 585
R271 B.n521 B.n6 585
R272 B.n798 B.n6 585
R273 B.n520 B.n5 585
R274 B.n799 B.n5 585
R275 B.n519 B.n518 585
R276 B.n518 B.n4 585
R277 B.n517 B.n127 585
R278 B.n517 B.n516 585
R279 B.n507 B.n128 585
R280 B.n129 B.n128 585
R281 B.n509 B.n508 585
R282 B.n510 B.n509 585
R283 B.n506 B.n134 585
R284 B.n134 B.n133 585
R285 B.n505 B.n504 585
R286 B.n504 B.n503 585
R287 B.n136 B.n135 585
R288 B.n496 B.n136 585
R289 B.n495 B.n494 585
R290 B.n497 B.n495 585
R291 B.n493 B.n141 585
R292 B.n141 B.n140 585
R293 B.n492 B.n491 585
R294 B.n491 B.n490 585
R295 B.n143 B.n142 585
R296 B.n144 B.n143 585
R297 B.n483 B.n482 585
R298 B.n484 B.n483 585
R299 B.n481 B.n149 585
R300 B.n149 B.n148 585
R301 B.n480 B.n479 585
R302 B.n479 B.n478 585
R303 B.n151 B.n150 585
R304 B.n152 B.n151 585
R305 B.n471 B.n470 585
R306 B.n472 B.n471 585
R307 B.n469 B.n156 585
R308 B.n160 B.n156 585
R309 B.n468 B.n467 585
R310 B.n467 B.n466 585
R311 B.n158 B.n157 585
R312 B.n159 B.n158 585
R313 B.n459 B.n458 585
R314 B.n460 B.n459 585
R315 B.n457 B.n165 585
R316 B.n165 B.n164 585
R317 B.n456 B.n455 585
R318 B.n455 B.n454 585
R319 B.n167 B.n166 585
R320 B.n168 B.n167 585
R321 B.n447 B.n446 585
R322 B.n448 B.n447 585
R323 B.n445 B.n173 585
R324 B.n173 B.n172 585
R325 B.n444 B.n443 585
R326 B.n443 B.n442 585
R327 B.n175 B.n174 585
R328 B.n176 B.n175 585
R329 B.n435 B.n434 585
R330 B.n436 B.n435 585
R331 B.n433 B.n181 585
R332 B.n181 B.n180 585
R333 B.n432 B.n431 585
R334 B.n431 B.n430 585
R335 B.n183 B.n182 585
R336 B.n184 B.n183 585
R337 B.n423 B.n422 585
R338 B.n424 B.n423 585
R339 B.n421 B.n189 585
R340 B.n189 B.n188 585
R341 B.n420 B.n419 585
R342 B.n419 B.n418 585
R343 B.n191 B.n190 585
R344 B.n192 B.n191 585
R345 B.n411 B.n410 585
R346 B.n412 B.n411 585
R347 B.n409 B.n197 585
R348 B.n197 B.n196 585
R349 B.n408 B.n407 585
R350 B.n407 B.n406 585
R351 B.n199 B.n198 585
R352 B.n200 B.n199 585
R353 B.n399 B.n398 585
R354 B.n400 B.n399 585
R355 B.n397 B.n205 585
R356 B.n205 B.n204 585
R357 B.n396 B.n395 585
R358 B.n395 B.n394 585
R359 B.n207 B.n206 585
R360 B.n208 B.n207 585
R361 B.n387 B.n386 585
R362 B.n388 B.n387 585
R363 B.n385 B.n213 585
R364 B.n213 B.n212 585
R365 B.n384 B.n383 585
R366 B.n383 B.n382 585
R367 B.n215 B.n214 585
R368 B.n216 B.n215 585
R369 B.n375 B.n374 585
R370 B.n376 B.n375 585
R371 B.n373 B.n221 585
R372 B.n221 B.n220 585
R373 B.n372 B.n371 585
R374 B.n371 B.n370 585
R375 B.n367 B.n225 585
R376 B.n366 B.n365 585
R377 B.n363 B.n226 585
R378 B.n363 B.n224 585
R379 B.n362 B.n361 585
R380 B.n360 B.n359 585
R381 B.n358 B.n228 585
R382 B.n356 B.n355 585
R383 B.n354 B.n229 585
R384 B.n353 B.n352 585
R385 B.n350 B.n230 585
R386 B.n348 B.n347 585
R387 B.n346 B.n231 585
R388 B.n345 B.n344 585
R389 B.n342 B.n232 585
R390 B.n340 B.n339 585
R391 B.n338 B.n233 585
R392 B.n337 B.n336 585
R393 B.n334 B.n234 585
R394 B.n332 B.n331 585
R395 B.n330 B.n235 585
R396 B.n329 B.n328 585
R397 B.n326 B.n236 585
R398 B.n324 B.n323 585
R399 B.n321 B.n237 585
R400 B.n320 B.n319 585
R401 B.n317 B.n240 585
R402 B.n315 B.n314 585
R403 B.n313 B.n241 585
R404 B.n312 B.n311 585
R405 B.n309 B.n242 585
R406 B.n307 B.n306 585
R407 B.n305 B.n243 585
R408 B.n304 B.n303 585
R409 B.n301 B.n300 585
R410 B.n299 B.n298 585
R411 B.n297 B.n248 585
R412 B.n295 B.n294 585
R413 B.n293 B.n249 585
R414 B.n292 B.n291 585
R415 B.n289 B.n250 585
R416 B.n287 B.n286 585
R417 B.n285 B.n251 585
R418 B.n284 B.n283 585
R419 B.n281 B.n252 585
R420 B.n279 B.n278 585
R421 B.n277 B.n253 585
R422 B.n276 B.n275 585
R423 B.n273 B.n254 585
R424 B.n271 B.n270 585
R425 B.n269 B.n255 585
R426 B.n268 B.n267 585
R427 B.n265 B.n256 585
R428 B.n263 B.n262 585
R429 B.n261 B.n257 585
R430 B.n260 B.n259 585
R431 B.n223 B.n222 585
R432 B.n224 B.n223 585
R433 B.n369 B.n368 585
R434 B.n370 B.n369 585
R435 B.n219 B.n218 585
R436 B.n220 B.n219 585
R437 B.n378 B.n377 585
R438 B.n377 B.n376 585
R439 B.n379 B.n217 585
R440 B.n217 B.n216 585
R441 B.n381 B.n380 585
R442 B.n382 B.n381 585
R443 B.n211 B.n210 585
R444 B.n212 B.n211 585
R445 B.n390 B.n389 585
R446 B.n389 B.n388 585
R447 B.n391 B.n209 585
R448 B.n209 B.n208 585
R449 B.n393 B.n392 585
R450 B.n394 B.n393 585
R451 B.n203 B.n202 585
R452 B.n204 B.n203 585
R453 B.n402 B.n401 585
R454 B.n401 B.n400 585
R455 B.n403 B.n201 585
R456 B.n201 B.n200 585
R457 B.n405 B.n404 585
R458 B.n406 B.n405 585
R459 B.n195 B.n194 585
R460 B.n196 B.n195 585
R461 B.n414 B.n413 585
R462 B.n413 B.n412 585
R463 B.n415 B.n193 585
R464 B.n193 B.n192 585
R465 B.n417 B.n416 585
R466 B.n418 B.n417 585
R467 B.n187 B.n186 585
R468 B.n188 B.n187 585
R469 B.n426 B.n425 585
R470 B.n425 B.n424 585
R471 B.n427 B.n185 585
R472 B.n185 B.n184 585
R473 B.n429 B.n428 585
R474 B.n430 B.n429 585
R475 B.n179 B.n178 585
R476 B.n180 B.n179 585
R477 B.n438 B.n437 585
R478 B.n437 B.n436 585
R479 B.n439 B.n177 585
R480 B.n177 B.n176 585
R481 B.n441 B.n440 585
R482 B.n442 B.n441 585
R483 B.n171 B.n170 585
R484 B.n172 B.n171 585
R485 B.n450 B.n449 585
R486 B.n449 B.n448 585
R487 B.n451 B.n169 585
R488 B.n169 B.n168 585
R489 B.n453 B.n452 585
R490 B.n454 B.n453 585
R491 B.n163 B.n162 585
R492 B.n164 B.n163 585
R493 B.n462 B.n461 585
R494 B.n461 B.n460 585
R495 B.n463 B.n161 585
R496 B.n161 B.n159 585
R497 B.n465 B.n464 585
R498 B.n466 B.n465 585
R499 B.n155 B.n154 585
R500 B.n160 B.n155 585
R501 B.n474 B.n473 585
R502 B.n473 B.n472 585
R503 B.n475 B.n153 585
R504 B.n153 B.n152 585
R505 B.n477 B.n476 585
R506 B.n478 B.n477 585
R507 B.n147 B.n146 585
R508 B.n148 B.n147 585
R509 B.n486 B.n485 585
R510 B.n485 B.n484 585
R511 B.n487 B.n145 585
R512 B.n145 B.n144 585
R513 B.n489 B.n488 585
R514 B.n490 B.n489 585
R515 B.n139 B.n138 585
R516 B.n140 B.n139 585
R517 B.n499 B.n498 585
R518 B.n498 B.n497 585
R519 B.n500 B.n137 585
R520 B.n496 B.n137 585
R521 B.n502 B.n501 585
R522 B.n503 B.n502 585
R523 B.n132 B.n131 585
R524 B.n133 B.n132 585
R525 B.n512 B.n511 585
R526 B.n511 B.n510 585
R527 B.n513 B.n130 585
R528 B.n130 B.n129 585
R529 B.n515 B.n514 585
R530 B.n516 B.n515 585
R531 B.n3 B.n0 585
R532 B.n4 B.n3 585
R533 B.n796 B.n1 585
R534 B.n797 B.n796 585
R535 B.n795 B.n794 585
R536 B.n795 B.n8 585
R537 B.n793 B.n9 585
R538 B.n12 B.n9 585
R539 B.n792 B.n791 585
R540 B.n791 B.n790 585
R541 B.n11 B.n10 585
R542 B.n789 B.n11 585
R543 B.n787 B.n786 585
R544 B.n788 B.n787 585
R545 B.n785 B.n16 585
R546 B.n19 B.n16 585
R547 B.n784 B.n783 585
R548 B.n783 B.n782 585
R549 B.n18 B.n17 585
R550 B.n781 B.n18 585
R551 B.n779 B.n778 585
R552 B.n780 B.n779 585
R553 B.n777 B.n24 585
R554 B.n24 B.n23 585
R555 B.n776 B.n775 585
R556 B.n775 B.n774 585
R557 B.n26 B.n25 585
R558 B.n773 B.n26 585
R559 B.n771 B.n770 585
R560 B.n772 B.n771 585
R561 B.n769 B.n31 585
R562 B.n31 B.n30 585
R563 B.n768 B.n767 585
R564 B.n767 B.n766 585
R565 B.n33 B.n32 585
R566 B.n765 B.n33 585
R567 B.n763 B.n762 585
R568 B.n764 B.n763 585
R569 B.n761 B.n38 585
R570 B.n38 B.n37 585
R571 B.n760 B.n759 585
R572 B.n759 B.n758 585
R573 B.n40 B.n39 585
R574 B.n757 B.n40 585
R575 B.n755 B.n754 585
R576 B.n756 B.n755 585
R577 B.n753 B.n45 585
R578 B.n45 B.n44 585
R579 B.n752 B.n751 585
R580 B.n751 B.n750 585
R581 B.n47 B.n46 585
R582 B.n749 B.n47 585
R583 B.n747 B.n746 585
R584 B.n748 B.n747 585
R585 B.n745 B.n52 585
R586 B.n52 B.n51 585
R587 B.n744 B.n743 585
R588 B.n743 B.n742 585
R589 B.n54 B.n53 585
R590 B.n741 B.n54 585
R591 B.n739 B.n738 585
R592 B.n740 B.n739 585
R593 B.n737 B.n59 585
R594 B.n59 B.n58 585
R595 B.n736 B.n735 585
R596 B.n735 B.n734 585
R597 B.n61 B.n60 585
R598 B.n733 B.n61 585
R599 B.n731 B.n730 585
R600 B.n732 B.n731 585
R601 B.n729 B.n66 585
R602 B.n66 B.n65 585
R603 B.n728 B.n727 585
R604 B.n727 B.n726 585
R605 B.n68 B.n67 585
R606 B.n725 B.n68 585
R607 B.n723 B.n722 585
R608 B.n724 B.n723 585
R609 B.n721 B.n73 585
R610 B.n73 B.n72 585
R611 B.n720 B.n719 585
R612 B.n719 B.n718 585
R613 B.n75 B.n74 585
R614 B.n717 B.n75 585
R615 B.n715 B.n714 585
R616 B.n716 B.n715 585
R617 B.n713 B.n80 585
R618 B.n80 B.n79 585
R619 B.n712 B.n711 585
R620 B.n711 B.n710 585
R621 B.n82 B.n81 585
R622 B.n709 B.n82 585
R623 B.n707 B.n706 585
R624 B.n708 B.n707 585
R625 B.n705 B.n87 585
R626 B.n87 B.n86 585
R627 B.n704 B.n703 585
R628 B.n703 B.n702 585
R629 B.n89 B.n88 585
R630 B.n701 B.n89 585
R631 B.n699 B.n698 585
R632 B.n700 B.n699 585
R633 B.n800 B.n799 585
R634 B.n798 B.n2 585
R635 B.n699 B.n94 444.452
R636 B.n586 B.n92 444.452
R637 B.n371 B.n223 444.452
R638 B.n369 B.n225 444.452
R639 B.n587 B.n93 256.663
R640 B.n589 B.n93 256.663
R641 B.n595 B.n93 256.663
R642 B.n597 B.n93 256.663
R643 B.n603 B.n93 256.663
R644 B.n605 B.n93 256.663
R645 B.n611 B.n93 256.663
R646 B.n613 B.n93 256.663
R647 B.n619 B.n93 256.663
R648 B.n621 B.n93 256.663
R649 B.n627 B.n93 256.663
R650 B.n629 B.n93 256.663
R651 B.n636 B.n93 256.663
R652 B.n638 B.n93 256.663
R653 B.n644 B.n93 256.663
R654 B.n646 B.n93 256.663
R655 B.n652 B.n93 256.663
R656 B.n654 B.n93 256.663
R657 B.n660 B.n93 256.663
R658 B.n662 B.n93 256.663
R659 B.n668 B.n93 256.663
R660 B.n670 B.n93 256.663
R661 B.n676 B.n93 256.663
R662 B.n678 B.n93 256.663
R663 B.n684 B.n93 256.663
R664 B.n686 B.n93 256.663
R665 B.n692 B.n93 256.663
R666 B.n694 B.n93 256.663
R667 B.n364 B.n224 256.663
R668 B.n227 B.n224 256.663
R669 B.n357 B.n224 256.663
R670 B.n351 B.n224 256.663
R671 B.n349 B.n224 256.663
R672 B.n343 B.n224 256.663
R673 B.n341 B.n224 256.663
R674 B.n335 B.n224 256.663
R675 B.n333 B.n224 256.663
R676 B.n327 B.n224 256.663
R677 B.n325 B.n224 256.663
R678 B.n318 B.n224 256.663
R679 B.n316 B.n224 256.663
R680 B.n310 B.n224 256.663
R681 B.n308 B.n224 256.663
R682 B.n302 B.n224 256.663
R683 B.n247 B.n224 256.663
R684 B.n296 B.n224 256.663
R685 B.n290 B.n224 256.663
R686 B.n288 B.n224 256.663
R687 B.n282 B.n224 256.663
R688 B.n280 B.n224 256.663
R689 B.n274 B.n224 256.663
R690 B.n272 B.n224 256.663
R691 B.n266 B.n224 256.663
R692 B.n264 B.n224 256.663
R693 B.n258 B.n224 256.663
R694 B.n802 B.n801 256.663
R695 B.n107 B.t17 250.855
R696 B.n114 B.t10 250.855
R697 B.n244 B.t6 250.855
R698 B.n238 B.t14 250.855
R699 B.n695 B.n693 163.367
R700 B.n691 B.n96 163.367
R701 B.n687 B.n685 163.367
R702 B.n683 B.n98 163.367
R703 B.n679 B.n677 163.367
R704 B.n675 B.n100 163.367
R705 B.n671 B.n669 163.367
R706 B.n667 B.n102 163.367
R707 B.n663 B.n661 163.367
R708 B.n659 B.n104 163.367
R709 B.n655 B.n653 163.367
R710 B.n651 B.n106 163.367
R711 B.n647 B.n645 163.367
R712 B.n643 B.n111 163.367
R713 B.n639 B.n637 163.367
R714 B.n635 B.n113 163.367
R715 B.n630 B.n628 163.367
R716 B.n626 B.n117 163.367
R717 B.n622 B.n620 163.367
R718 B.n618 B.n119 163.367
R719 B.n614 B.n612 163.367
R720 B.n610 B.n121 163.367
R721 B.n606 B.n604 163.367
R722 B.n602 B.n123 163.367
R723 B.n598 B.n596 163.367
R724 B.n594 B.n125 163.367
R725 B.n590 B.n588 163.367
R726 B.n371 B.n221 163.367
R727 B.n375 B.n221 163.367
R728 B.n375 B.n215 163.367
R729 B.n383 B.n215 163.367
R730 B.n383 B.n213 163.367
R731 B.n387 B.n213 163.367
R732 B.n387 B.n207 163.367
R733 B.n395 B.n207 163.367
R734 B.n395 B.n205 163.367
R735 B.n399 B.n205 163.367
R736 B.n399 B.n199 163.367
R737 B.n407 B.n199 163.367
R738 B.n407 B.n197 163.367
R739 B.n411 B.n197 163.367
R740 B.n411 B.n191 163.367
R741 B.n419 B.n191 163.367
R742 B.n419 B.n189 163.367
R743 B.n423 B.n189 163.367
R744 B.n423 B.n183 163.367
R745 B.n431 B.n183 163.367
R746 B.n431 B.n181 163.367
R747 B.n435 B.n181 163.367
R748 B.n435 B.n175 163.367
R749 B.n443 B.n175 163.367
R750 B.n443 B.n173 163.367
R751 B.n447 B.n173 163.367
R752 B.n447 B.n167 163.367
R753 B.n455 B.n167 163.367
R754 B.n455 B.n165 163.367
R755 B.n459 B.n165 163.367
R756 B.n459 B.n158 163.367
R757 B.n467 B.n158 163.367
R758 B.n467 B.n156 163.367
R759 B.n471 B.n156 163.367
R760 B.n471 B.n151 163.367
R761 B.n479 B.n151 163.367
R762 B.n479 B.n149 163.367
R763 B.n483 B.n149 163.367
R764 B.n483 B.n143 163.367
R765 B.n491 B.n143 163.367
R766 B.n491 B.n141 163.367
R767 B.n495 B.n141 163.367
R768 B.n495 B.n136 163.367
R769 B.n504 B.n136 163.367
R770 B.n504 B.n134 163.367
R771 B.n509 B.n134 163.367
R772 B.n509 B.n128 163.367
R773 B.n517 B.n128 163.367
R774 B.n518 B.n517 163.367
R775 B.n518 B.n5 163.367
R776 B.n6 B.n5 163.367
R777 B.n7 B.n6 163.367
R778 B.n524 B.n7 163.367
R779 B.n525 B.n524 163.367
R780 B.n525 B.n13 163.367
R781 B.n14 B.n13 163.367
R782 B.n15 B.n14 163.367
R783 B.n530 B.n15 163.367
R784 B.n530 B.n20 163.367
R785 B.n21 B.n20 163.367
R786 B.n22 B.n21 163.367
R787 B.n535 B.n22 163.367
R788 B.n535 B.n27 163.367
R789 B.n28 B.n27 163.367
R790 B.n29 B.n28 163.367
R791 B.n540 B.n29 163.367
R792 B.n540 B.n34 163.367
R793 B.n35 B.n34 163.367
R794 B.n36 B.n35 163.367
R795 B.n545 B.n36 163.367
R796 B.n545 B.n41 163.367
R797 B.n42 B.n41 163.367
R798 B.n43 B.n42 163.367
R799 B.n550 B.n43 163.367
R800 B.n550 B.n48 163.367
R801 B.n49 B.n48 163.367
R802 B.n50 B.n49 163.367
R803 B.n555 B.n50 163.367
R804 B.n555 B.n55 163.367
R805 B.n56 B.n55 163.367
R806 B.n57 B.n56 163.367
R807 B.n560 B.n57 163.367
R808 B.n560 B.n62 163.367
R809 B.n63 B.n62 163.367
R810 B.n64 B.n63 163.367
R811 B.n565 B.n64 163.367
R812 B.n565 B.n69 163.367
R813 B.n70 B.n69 163.367
R814 B.n71 B.n70 163.367
R815 B.n570 B.n71 163.367
R816 B.n570 B.n76 163.367
R817 B.n77 B.n76 163.367
R818 B.n78 B.n77 163.367
R819 B.n575 B.n78 163.367
R820 B.n575 B.n83 163.367
R821 B.n84 B.n83 163.367
R822 B.n85 B.n84 163.367
R823 B.n580 B.n85 163.367
R824 B.n580 B.n90 163.367
R825 B.n91 B.n90 163.367
R826 B.n92 B.n91 163.367
R827 B.n365 B.n363 163.367
R828 B.n363 B.n362 163.367
R829 B.n359 B.n358 163.367
R830 B.n356 B.n229 163.367
R831 B.n352 B.n350 163.367
R832 B.n348 B.n231 163.367
R833 B.n344 B.n342 163.367
R834 B.n340 B.n233 163.367
R835 B.n336 B.n334 163.367
R836 B.n332 B.n235 163.367
R837 B.n328 B.n326 163.367
R838 B.n324 B.n237 163.367
R839 B.n319 B.n317 163.367
R840 B.n315 B.n241 163.367
R841 B.n311 B.n309 163.367
R842 B.n307 B.n243 163.367
R843 B.n303 B.n301 163.367
R844 B.n298 B.n297 163.367
R845 B.n295 B.n249 163.367
R846 B.n291 B.n289 163.367
R847 B.n287 B.n251 163.367
R848 B.n283 B.n281 163.367
R849 B.n279 B.n253 163.367
R850 B.n275 B.n273 163.367
R851 B.n271 B.n255 163.367
R852 B.n267 B.n265 163.367
R853 B.n263 B.n257 163.367
R854 B.n259 B.n223 163.367
R855 B.n369 B.n219 163.367
R856 B.n377 B.n219 163.367
R857 B.n377 B.n217 163.367
R858 B.n381 B.n217 163.367
R859 B.n381 B.n211 163.367
R860 B.n389 B.n211 163.367
R861 B.n389 B.n209 163.367
R862 B.n393 B.n209 163.367
R863 B.n393 B.n203 163.367
R864 B.n401 B.n203 163.367
R865 B.n401 B.n201 163.367
R866 B.n405 B.n201 163.367
R867 B.n405 B.n195 163.367
R868 B.n413 B.n195 163.367
R869 B.n413 B.n193 163.367
R870 B.n417 B.n193 163.367
R871 B.n417 B.n187 163.367
R872 B.n425 B.n187 163.367
R873 B.n425 B.n185 163.367
R874 B.n429 B.n185 163.367
R875 B.n429 B.n179 163.367
R876 B.n437 B.n179 163.367
R877 B.n437 B.n177 163.367
R878 B.n441 B.n177 163.367
R879 B.n441 B.n171 163.367
R880 B.n449 B.n171 163.367
R881 B.n449 B.n169 163.367
R882 B.n453 B.n169 163.367
R883 B.n453 B.n163 163.367
R884 B.n461 B.n163 163.367
R885 B.n461 B.n161 163.367
R886 B.n465 B.n161 163.367
R887 B.n465 B.n155 163.367
R888 B.n473 B.n155 163.367
R889 B.n473 B.n153 163.367
R890 B.n477 B.n153 163.367
R891 B.n477 B.n147 163.367
R892 B.n485 B.n147 163.367
R893 B.n485 B.n145 163.367
R894 B.n489 B.n145 163.367
R895 B.n489 B.n139 163.367
R896 B.n498 B.n139 163.367
R897 B.n498 B.n137 163.367
R898 B.n502 B.n137 163.367
R899 B.n502 B.n132 163.367
R900 B.n511 B.n132 163.367
R901 B.n511 B.n130 163.367
R902 B.n515 B.n130 163.367
R903 B.n515 B.n3 163.367
R904 B.n800 B.n3 163.367
R905 B.n796 B.n2 163.367
R906 B.n796 B.n795 163.367
R907 B.n795 B.n9 163.367
R908 B.n791 B.n9 163.367
R909 B.n791 B.n11 163.367
R910 B.n787 B.n11 163.367
R911 B.n787 B.n16 163.367
R912 B.n783 B.n16 163.367
R913 B.n783 B.n18 163.367
R914 B.n779 B.n18 163.367
R915 B.n779 B.n24 163.367
R916 B.n775 B.n24 163.367
R917 B.n775 B.n26 163.367
R918 B.n771 B.n26 163.367
R919 B.n771 B.n31 163.367
R920 B.n767 B.n31 163.367
R921 B.n767 B.n33 163.367
R922 B.n763 B.n33 163.367
R923 B.n763 B.n38 163.367
R924 B.n759 B.n38 163.367
R925 B.n759 B.n40 163.367
R926 B.n755 B.n40 163.367
R927 B.n755 B.n45 163.367
R928 B.n751 B.n45 163.367
R929 B.n751 B.n47 163.367
R930 B.n747 B.n47 163.367
R931 B.n747 B.n52 163.367
R932 B.n743 B.n52 163.367
R933 B.n743 B.n54 163.367
R934 B.n739 B.n54 163.367
R935 B.n739 B.n59 163.367
R936 B.n735 B.n59 163.367
R937 B.n735 B.n61 163.367
R938 B.n731 B.n61 163.367
R939 B.n731 B.n66 163.367
R940 B.n727 B.n66 163.367
R941 B.n727 B.n68 163.367
R942 B.n723 B.n68 163.367
R943 B.n723 B.n73 163.367
R944 B.n719 B.n73 163.367
R945 B.n719 B.n75 163.367
R946 B.n715 B.n75 163.367
R947 B.n715 B.n80 163.367
R948 B.n711 B.n80 163.367
R949 B.n711 B.n82 163.367
R950 B.n707 B.n82 163.367
R951 B.n707 B.n87 163.367
R952 B.n703 B.n87 163.367
R953 B.n703 B.n89 163.367
R954 B.n699 B.n89 163.367
R955 B.n114 B.t12 143.929
R956 B.n244 B.t9 143.929
R957 B.n107 B.t18 143.923
R958 B.n238 B.t16 143.923
R959 B.n370 B.n224 113.465
R960 B.n700 B.n93 113.465
R961 B.n115 B.t13 74.3048
R962 B.n245 B.t8 74.3048
R963 B.n108 B.t19 74.299
R964 B.n239 B.t15 74.299
R965 B.n694 B.n94 71.676
R966 B.n693 B.n692 71.676
R967 B.n686 B.n96 71.676
R968 B.n685 B.n684 71.676
R969 B.n678 B.n98 71.676
R970 B.n677 B.n676 71.676
R971 B.n670 B.n100 71.676
R972 B.n669 B.n668 71.676
R973 B.n662 B.n102 71.676
R974 B.n661 B.n660 71.676
R975 B.n654 B.n104 71.676
R976 B.n653 B.n652 71.676
R977 B.n646 B.n106 71.676
R978 B.n645 B.n644 71.676
R979 B.n638 B.n111 71.676
R980 B.n637 B.n636 71.676
R981 B.n629 B.n113 71.676
R982 B.n628 B.n627 71.676
R983 B.n621 B.n117 71.676
R984 B.n620 B.n619 71.676
R985 B.n613 B.n119 71.676
R986 B.n612 B.n611 71.676
R987 B.n605 B.n121 71.676
R988 B.n604 B.n603 71.676
R989 B.n597 B.n123 71.676
R990 B.n596 B.n595 71.676
R991 B.n589 B.n125 71.676
R992 B.n588 B.n587 71.676
R993 B.n587 B.n586 71.676
R994 B.n590 B.n589 71.676
R995 B.n595 B.n594 71.676
R996 B.n598 B.n597 71.676
R997 B.n603 B.n602 71.676
R998 B.n606 B.n605 71.676
R999 B.n611 B.n610 71.676
R1000 B.n614 B.n613 71.676
R1001 B.n619 B.n618 71.676
R1002 B.n622 B.n621 71.676
R1003 B.n627 B.n626 71.676
R1004 B.n630 B.n629 71.676
R1005 B.n636 B.n635 71.676
R1006 B.n639 B.n638 71.676
R1007 B.n644 B.n643 71.676
R1008 B.n647 B.n646 71.676
R1009 B.n652 B.n651 71.676
R1010 B.n655 B.n654 71.676
R1011 B.n660 B.n659 71.676
R1012 B.n663 B.n662 71.676
R1013 B.n668 B.n667 71.676
R1014 B.n671 B.n670 71.676
R1015 B.n676 B.n675 71.676
R1016 B.n679 B.n678 71.676
R1017 B.n684 B.n683 71.676
R1018 B.n687 B.n686 71.676
R1019 B.n692 B.n691 71.676
R1020 B.n695 B.n694 71.676
R1021 B.n364 B.n225 71.676
R1022 B.n362 B.n227 71.676
R1023 B.n358 B.n357 71.676
R1024 B.n351 B.n229 71.676
R1025 B.n350 B.n349 71.676
R1026 B.n343 B.n231 71.676
R1027 B.n342 B.n341 71.676
R1028 B.n335 B.n233 71.676
R1029 B.n334 B.n333 71.676
R1030 B.n327 B.n235 71.676
R1031 B.n326 B.n325 71.676
R1032 B.n318 B.n237 71.676
R1033 B.n317 B.n316 71.676
R1034 B.n310 B.n241 71.676
R1035 B.n309 B.n308 71.676
R1036 B.n302 B.n243 71.676
R1037 B.n301 B.n247 71.676
R1038 B.n297 B.n296 71.676
R1039 B.n290 B.n249 71.676
R1040 B.n289 B.n288 71.676
R1041 B.n282 B.n251 71.676
R1042 B.n281 B.n280 71.676
R1043 B.n274 B.n253 71.676
R1044 B.n273 B.n272 71.676
R1045 B.n266 B.n255 71.676
R1046 B.n265 B.n264 71.676
R1047 B.n258 B.n257 71.676
R1048 B.n365 B.n364 71.676
R1049 B.n359 B.n227 71.676
R1050 B.n357 B.n356 71.676
R1051 B.n352 B.n351 71.676
R1052 B.n349 B.n348 71.676
R1053 B.n344 B.n343 71.676
R1054 B.n341 B.n340 71.676
R1055 B.n336 B.n335 71.676
R1056 B.n333 B.n332 71.676
R1057 B.n328 B.n327 71.676
R1058 B.n325 B.n324 71.676
R1059 B.n319 B.n318 71.676
R1060 B.n316 B.n315 71.676
R1061 B.n311 B.n310 71.676
R1062 B.n308 B.n307 71.676
R1063 B.n303 B.n302 71.676
R1064 B.n298 B.n247 71.676
R1065 B.n296 B.n295 71.676
R1066 B.n291 B.n290 71.676
R1067 B.n288 B.n287 71.676
R1068 B.n283 B.n282 71.676
R1069 B.n280 B.n279 71.676
R1070 B.n275 B.n274 71.676
R1071 B.n272 B.n271 71.676
R1072 B.n267 B.n266 71.676
R1073 B.n264 B.n263 71.676
R1074 B.n259 B.n258 71.676
R1075 B.n801 B.n800 71.676
R1076 B.n801 B.n2 71.676
R1077 B.n108 B.n107 69.6247
R1078 B.n115 B.n114 69.6247
R1079 B.n245 B.n244 69.6247
R1080 B.n239 B.n238 69.6247
R1081 B.n370 B.n220 68.2798
R1082 B.n376 B.n220 68.2798
R1083 B.n376 B.n216 68.2798
R1084 B.n382 B.n216 68.2798
R1085 B.n382 B.n212 68.2798
R1086 B.n388 B.n212 68.2798
R1087 B.n388 B.n208 68.2798
R1088 B.n394 B.n208 68.2798
R1089 B.n400 B.n204 68.2798
R1090 B.n400 B.n200 68.2798
R1091 B.n406 B.n200 68.2798
R1092 B.n406 B.n196 68.2798
R1093 B.n412 B.n196 68.2798
R1094 B.n412 B.n192 68.2798
R1095 B.n418 B.n192 68.2798
R1096 B.n418 B.n188 68.2798
R1097 B.n424 B.n188 68.2798
R1098 B.n424 B.n184 68.2798
R1099 B.n430 B.n184 68.2798
R1100 B.n430 B.n180 68.2798
R1101 B.n436 B.n180 68.2798
R1102 B.n442 B.n176 68.2798
R1103 B.n442 B.n172 68.2798
R1104 B.n448 B.n172 68.2798
R1105 B.n448 B.n168 68.2798
R1106 B.n454 B.n168 68.2798
R1107 B.n454 B.n164 68.2798
R1108 B.n460 B.n164 68.2798
R1109 B.n460 B.n159 68.2798
R1110 B.n466 B.n159 68.2798
R1111 B.n466 B.n160 68.2798
R1112 B.n472 B.n152 68.2798
R1113 B.n478 B.n152 68.2798
R1114 B.n478 B.n148 68.2798
R1115 B.n484 B.n148 68.2798
R1116 B.n484 B.n144 68.2798
R1117 B.n490 B.n144 68.2798
R1118 B.n490 B.n140 68.2798
R1119 B.n497 B.n140 68.2798
R1120 B.n497 B.n496 68.2798
R1121 B.n503 B.n133 68.2798
R1122 B.n510 B.n133 68.2798
R1123 B.n510 B.n129 68.2798
R1124 B.n516 B.n129 68.2798
R1125 B.n516 B.n4 68.2798
R1126 B.n799 B.n4 68.2798
R1127 B.n799 B.n798 68.2798
R1128 B.n798 B.n797 68.2798
R1129 B.n797 B.n8 68.2798
R1130 B.n12 B.n8 68.2798
R1131 B.n790 B.n12 68.2798
R1132 B.n790 B.n789 68.2798
R1133 B.n789 B.n788 68.2798
R1134 B.n782 B.n19 68.2798
R1135 B.n782 B.n781 68.2798
R1136 B.n781 B.n780 68.2798
R1137 B.n780 B.n23 68.2798
R1138 B.n774 B.n23 68.2798
R1139 B.n774 B.n773 68.2798
R1140 B.n773 B.n772 68.2798
R1141 B.n772 B.n30 68.2798
R1142 B.n766 B.n30 68.2798
R1143 B.n765 B.n764 68.2798
R1144 B.n764 B.n37 68.2798
R1145 B.n758 B.n37 68.2798
R1146 B.n758 B.n757 68.2798
R1147 B.n757 B.n756 68.2798
R1148 B.n756 B.n44 68.2798
R1149 B.n750 B.n44 68.2798
R1150 B.n750 B.n749 68.2798
R1151 B.n749 B.n748 68.2798
R1152 B.n748 B.n51 68.2798
R1153 B.n742 B.n741 68.2798
R1154 B.n741 B.n740 68.2798
R1155 B.n740 B.n58 68.2798
R1156 B.n734 B.n58 68.2798
R1157 B.n734 B.n733 68.2798
R1158 B.n733 B.n732 68.2798
R1159 B.n732 B.n65 68.2798
R1160 B.n726 B.n65 68.2798
R1161 B.n726 B.n725 68.2798
R1162 B.n725 B.n724 68.2798
R1163 B.n724 B.n72 68.2798
R1164 B.n718 B.n72 68.2798
R1165 B.n718 B.n717 68.2798
R1166 B.n716 B.n79 68.2798
R1167 B.n710 B.n79 68.2798
R1168 B.n710 B.n709 68.2798
R1169 B.n709 B.n708 68.2798
R1170 B.n708 B.n86 68.2798
R1171 B.n702 B.n86 68.2798
R1172 B.n702 B.n701 68.2798
R1173 B.n701 B.n700 68.2798
R1174 B.n472 B.t2 64.2634
R1175 B.n766 B.t1 64.2634
R1176 B.n109 B.n108 59.5399
R1177 B.n632 B.n115 59.5399
R1178 B.n246 B.n245 59.5399
R1179 B.n322 B.n239 59.5399
R1180 B.n394 B.t7 50.2059
R1181 B.t11 B.n716 50.2059
R1182 B.n496 B.t3 42.173
R1183 B.n19 B.t5 42.173
R1184 B.n436 B.t0 34.1402
R1185 B.t0 B.n176 34.1402
R1186 B.t4 B.n51 34.1402
R1187 B.n742 B.t4 34.1402
R1188 B.n368 B.n367 28.8785
R1189 B.n372 B.n222 28.8785
R1190 B.n585 B.n584 28.8785
R1191 B.n698 B.n697 28.8785
R1192 B.n503 B.t3 26.1073
R1193 B.n788 B.t5 26.1073
R1194 B.t7 B.n204 18.0744
R1195 B.n717 B.t11 18.0744
R1196 B B.n802 18.0485
R1197 B.n368 B.n218 10.6151
R1198 B.n378 B.n218 10.6151
R1199 B.n379 B.n378 10.6151
R1200 B.n380 B.n379 10.6151
R1201 B.n380 B.n210 10.6151
R1202 B.n390 B.n210 10.6151
R1203 B.n391 B.n390 10.6151
R1204 B.n392 B.n391 10.6151
R1205 B.n392 B.n202 10.6151
R1206 B.n402 B.n202 10.6151
R1207 B.n403 B.n402 10.6151
R1208 B.n404 B.n403 10.6151
R1209 B.n404 B.n194 10.6151
R1210 B.n414 B.n194 10.6151
R1211 B.n415 B.n414 10.6151
R1212 B.n416 B.n415 10.6151
R1213 B.n416 B.n186 10.6151
R1214 B.n426 B.n186 10.6151
R1215 B.n427 B.n426 10.6151
R1216 B.n428 B.n427 10.6151
R1217 B.n428 B.n178 10.6151
R1218 B.n438 B.n178 10.6151
R1219 B.n439 B.n438 10.6151
R1220 B.n440 B.n439 10.6151
R1221 B.n440 B.n170 10.6151
R1222 B.n450 B.n170 10.6151
R1223 B.n451 B.n450 10.6151
R1224 B.n452 B.n451 10.6151
R1225 B.n452 B.n162 10.6151
R1226 B.n462 B.n162 10.6151
R1227 B.n463 B.n462 10.6151
R1228 B.n464 B.n463 10.6151
R1229 B.n464 B.n154 10.6151
R1230 B.n474 B.n154 10.6151
R1231 B.n475 B.n474 10.6151
R1232 B.n476 B.n475 10.6151
R1233 B.n476 B.n146 10.6151
R1234 B.n486 B.n146 10.6151
R1235 B.n487 B.n486 10.6151
R1236 B.n488 B.n487 10.6151
R1237 B.n488 B.n138 10.6151
R1238 B.n499 B.n138 10.6151
R1239 B.n500 B.n499 10.6151
R1240 B.n501 B.n500 10.6151
R1241 B.n501 B.n131 10.6151
R1242 B.n512 B.n131 10.6151
R1243 B.n513 B.n512 10.6151
R1244 B.n514 B.n513 10.6151
R1245 B.n514 B.n0 10.6151
R1246 B.n367 B.n366 10.6151
R1247 B.n366 B.n226 10.6151
R1248 B.n361 B.n226 10.6151
R1249 B.n361 B.n360 10.6151
R1250 B.n360 B.n228 10.6151
R1251 B.n355 B.n228 10.6151
R1252 B.n355 B.n354 10.6151
R1253 B.n354 B.n353 10.6151
R1254 B.n353 B.n230 10.6151
R1255 B.n347 B.n230 10.6151
R1256 B.n347 B.n346 10.6151
R1257 B.n346 B.n345 10.6151
R1258 B.n345 B.n232 10.6151
R1259 B.n339 B.n232 10.6151
R1260 B.n339 B.n338 10.6151
R1261 B.n338 B.n337 10.6151
R1262 B.n337 B.n234 10.6151
R1263 B.n331 B.n234 10.6151
R1264 B.n331 B.n330 10.6151
R1265 B.n330 B.n329 10.6151
R1266 B.n329 B.n236 10.6151
R1267 B.n323 B.n236 10.6151
R1268 B.n321 B.n320 10.6151
R1269 B.n320 B.n240 10.6151
R1270 B.n314 B.n240 10.6151
R1271 B.n314 B.n313 10.6151
R1272 B.n313 B.n312 10.6151
R1273 B.n312 B.n242 10.6151
R1274 B.n306 B.n242 10.6151
R1275 B.n306 B.n305 10.6151
R1276 B.n305 B.n304 10.6151
R1277 B.n300 B.n299 10.6151
R1278 B.n299 B.n248 10.6151
R1279 B.n294 B.n248 10.6151
R1280 B.n294 B.n293 10.6151
R1281 B.n293 B.n292 10.6151
R1282 B.n292 B.n250 10.6151
R1283 B.n286 B.n250 10.6151
R1284 B.n286 B.n285 10.6151
R1285 B.n285 B.n284 10.6151
R1286 B.n284 B.n252 10.6151
R1287 B.n278 B.n252 10.6151
R1288 B.n278 B.n277 10.6151
R1289 B.n277 B.n276 10.6151
R1290 B.n276 B.n254 10.6151
R1291 B.n270 B.n254 10.6151
R1292 B.n270 B.n269 10.6151
R1293 B.n269 B.n268 10.6151
R1294 B.n268 B.n256 10.6151
R1295 B.n262 B.n256 10.6151
R1296 B.n262 B.n261 10.6151
R1297 B.n261 B.n260 10.6151
R1298 B.n260 B.n222 10.6151
R1299 B.n373 B.n372 10.6151
R1300 B.n374 B.n373 10.6151
R1301 B.n374 B.n214 10.6151
R1302 B.n384 B.n214 10.6151
R1303 B.n385 B.n384 10.6151
R1304 B.n386 B.n385 10.6151
R1305 B.n386 B.n206 10.6151
R1306 B.n396 B.n206 10.6151
R1307 B.n397 B.n396 10.6151
R1308 B.n398 B.n397 10.6151
R1309 B.n398 B.n198 10.6151
R1310 B.n408 B.n198 10.6151
R1311 B.n409 B.n408 10.6151
R1312 B.n410 B.n409 10.6151
R1313 B.n410 B.n190 10.6151
R1314 B.n420 B.n190 10.6151
R1315 B.n421 B.n420 10.6151
R1316 B.n422 B.n421 10.6151
R1317 B.n422 B.n182 10.6151
R1318 B.n432 B.n182 10.6151
R1319 B.n433 B.n432 10.6151
R1320 B.n434 B.n433 10.6151
R1321 B.n434 B.n174 10.6151
R1322 B.n444 B.n174 10.6151
R1323 B.n445 B.n444 10.6151
R1324 B.n446 B.n445 10.6151
R1325 B.n446 B.n166 10.6151
R1326 B.n456 B.n166 10.6151
R1327 B.n457 B.n456 10.6151
R1328 B.n458 B.n457 10.6151
R1329 B.n458 B.n157 10.6151
R1330 B.n468 B.n157 10.6151
R1331 B.n469 B.n468 10.6151
R1332 B.n470 B.n469 10.6151
R1333 B.n470 B.n150 10.6151
R1334 B.n480 B.n150 10.6151
R1335 B.n481 B.n480 10.6151
R1336 B.n482 B.n481 10.6151
R1337 B.n482 B.n142 10.6151
R1338 B.n492 B.n142 10.6151
R1339 B.n493 B.n492 10.6151
R1340 B.n494 B.n493 10.6151
R1341 B.n494 B.n135 10.6151
R1342 B.n505 B.n135 10.6151
R1343 B.n506 B.n505 10.6151
R1344 B.n508 B.n506 10.6151
R1345 B.n508 B.n507 10.6151
R1346 B.n507 B.n127 10.6151
R1347 B.n519 B.n127 10.6151
R1348 B.n520 B.n519 10.6151
R1349 B.n521 B.n520 10.6151
R1350 B.n522 B.n521 10.6151
R1351 B.n523 B.n522 10.6151
R1352 B.n526 B.n523 10.6151
R1353 B.n527 B.n526 10.6151
R1354 B.n528 B.n527 10.6151
R1355 B.n529 B.n528 10.6151
R1356 B.n531 B.n529 10.6151
R1357 B.n532 B.n531 10.6151
R1358 B.n533 B.n532 10.6151
R1359 B.n534 B.n533 10.6151
R1360 B.n536 B.n534 10.6151
R1361 B.n537 B.n536 10.6151
R1362 B.n538 B.n537 10.6151
R1363 B.n539 B.n538 10.6151
R1364 B.n541 B.n539 10.6151
R1365 B.n542 B.n541 10.6151
R1366 B.n543 B.n542 10.6151
R1367 B.n544 B.n543 10.6151
R1368 B.n546 B.n544 10.6151
R1369 B.n547 B.n546 10.6151
R1370 B.n548 B.n547 10.6151
R1371 B.n549 B.n548 10.6151
R1372 B.n551 B.n549 10.6151
R1373 B.n552 B.n551 10.6151
R1374 B.n553 B.n552 10.6151
R1375 B.n554 B.n553 10.6151
R1376 B.n556 B.n554 10.6151
R1377 B.n557 B.n556 10.6151
R1378 B.n558 B.n557 10.6151
R1379 B.n559 B.n558 10.6151
R1380 B.n561 B.n559 10.6151
R1381 B.n562 B.n561 10.6151
R1382 B.n563 B.n562 10.6151
R1383 B.n564 B.n563 10.6151
R1384 B.n566 B.n564 10.6151
R1385 B.n567 B.n566 10.6151
R1386 B.n568 B.n567 10.6151
R1387 B.n569 B.n568 10.6151
R1388 B.n571 B.n569 10.6151
R1389 B.n572 B.n571 10.6151
R1390 B.n573 B.n572 10.6151
R1391 B.n574 B.n573 10.6151
R1392 B.n576 B.n574 10.6151
R1393 B.n577 B.n576 10.6151
R1394 B.n578 B.n577 10.6151
R1395 B.n579 B.n578 10.6151
R1396 B.n581 B.n579 10.6151
R1397 B.n582 B.n581 10.6151
R1398 B.n583 B.n582 10.6151
R1399 B.n584 B.n583 10.6151
R1400 B.n794 B.n1 10.6151
R1401 B.n794 B.n793 10.6151
R1402 B.n793 B.n792 10.6151
R1403 B.n792 B.n10 10.6151
R1404 B.n786 B.n10 10.6151
R1405 B.n786 B.n785 10.6151
R1406 B.n785 B.n784 10.6151
R1407 B.n784 B.n17 10.6151
R1408 B.n778 B.n17 10.6151
R1409 B.n778 B.n777 10.6151
R1410 B.n777 B.n776 10.6151
R1411 B.n776 B.n25 10.6151
R1412 B.n770 B.n25 10.6151
R1413 B.n770 B.n769 10.6151
R1414 B.n769 B.n768 10.6151
R1415 B.n768 B.n32 10.6151
R1416 B.n762 B.n32 10.6151
R1417 B.n762 B.n761 10.6151
R1418 B.n761 B.n760 10.6151
R1419 B.n760 B.n39 10.6151
R1420 B.n754 B.n39 10.6151
R1421 B.n754 B.n753 10.6151
R1422 B.n753 B.n752 10.6151
R1423 B.n752 B.n46 10.6151
R1424 B.n746 B.n46 10.6151
R1425 B.n746 B.n745 10.6151
R1426 B.n745 B.n744 10.6151
R1427 B.n744 B.n53 10.6151
R1428 B.n738 B.n53 10.6151
R1429 B.n738 B.n737 10.6151
R1430 B.n737 B.n736 10.6151
R1431 B.n736 B.n60 10.6151
R1432 B.n730 B.n60 10.6151
R1433 B.n730 B.n729 10.6151
R1434 B.n729 B.n728 10.6151
R1435 B.n728 B.n67 10.6151
R1436 B.n722 B.n67 10.6151
R1437 B.n722 B.n721 10.6151
R1438 B.n721 B.n720 10.6151
R1439 B.n720 B.n74 10.6151
R1440 B.n714 B.n74 10.6151
R1441 B.n714 B.n713 10.6151
R1442 B.n713 B.n712 10.6151
R1443 B.n712 B.n81 10.6151
R1444 B.n706 B.n81 10.6151
R1445 B.n706 B.n705 10.6151
R1446 B.n705 B.n704 10.6151
R1447 B.n704 B.n88 10.6151
R1448 B.n698 B.n88 10.6151
R1449 B.n697 B.n696 10.6151
R1450 B.n696 B.n95 10.6151
R1451 B.n690 B.n95 10.6151
R1452 B.n690 B.n689 10.6151
R1453 B.n689 B.n688 10.6151
R1454 B.n688 B.n97 10.6151
R1455 B.n682 B.n97 10.6151
R1456 B.n682 B.n681 10.6151
R1457 B.n681 B.n680 10.6151
R1458 B.n680 B.n99 10.6151
R1459 B.n674 B.n99 10.6151
R1460 B.n674 B.n673 10.6151
R1461 B.n673 B.n672 10.6151
R1462 B.n672 B.n101 10.6151
R1463 B.n666 B.n101 10.6151
R1464 B.n666 B.n665 10.6151
R1465 B.n665 B.n664 10.6151
R1466 B.n664 B.n103 10.6151
R1467 B.n658 B.n103 10.6151
R1468 B.n658 B.n657 10.6151
R1469 B.n657 B.n656 10.6151
R1470 B.n656 B.n105 10.6151
R1471 B.n650 B.n649 10.6151
R1472 B.n649 B.n648 10.6151
R1473 B.n648 B.n110 10.6151
R1474 B.n642 B.n110 10.6151
R1475 B.n642 B.n641 10.6151
R1476 B.n641 B.n640 10.6151
R1477 B.n640 B.n112 10.6151
R1478 B.n634 B.n112 10.6151
R1479 B.n634 B.n633 10.6151
R1480 B.n631 B.n116 10.6151
R1481 B.n625 B.n116 10.6151
R1482 B.n625 B.n624 10.6151
R1483 B.n624 B.n623 10.6151
R1484 B.n623 B.n118 10.6151
R1485 B.n617 B.n118 10.6151
R1486 B.n617 B.n616 10.6151
R1487 B.n616 B.n615 10.6151
R1488 B.n615 B.n120 10.6151
R1489 B.n609 B.n120 10.6151
R1490 B.n609 B.n608 10.6151
R1491 B.n608 B.n607 10.6151
R1492 B.n607 B.n122 10.6151
R1493 B.n601 B.n122 10.6151
R1494 B.n601 B.n600 10.6151
R1495 B.n600 B.n599 10.6151
R1496 B.n599 B.n124 10.6151
R1497 B.n593 B.n124 10.6151
R1498 B.n593 B.n592 10.6151
R1499 B.n592 B.n591 10.6151
R1500 B.n591 B.n126 10.6151
R1501 B.n585 B.n126 10.6151
R1502 B.n323 B.n322 9.36635
R1503 B.n300 B.n246 9.36635
R1504 B.n109 B.n105 9.36635
R1505 B.n632 B.n631 9.36635
R1506 B.n802 B.n0 8.11757
R1507 B.n802 B.n1 8.11757
R1508 B.n160 B.t2 4.01693
R1509 B.t1 B.n765 4.01693
R1510 B.n322 B.n321 1.24928
R1511 B.n304 B.n246 1.24928
R1512 B.n650 B.n109 1.24928
R1513 B.n633 B.n632 1.24928
R1514 VN.n34 VN.n33 161.3
R1515 VN.n32 VN.n19 161.3
R1516 VN.n31 VN.n30 161.3
R1517 VN.n29 VN.n20 161.3
R1518 VN.n28 VN.n27 161.3
R1519 VN.n26 VN.n21 161.3
R1520 VN.n25 VN.n24 161.3
R1521 VN.n16 VN.n15 161.3
R1522 VN.n14 VN.n1 161.3
R1523 VN.n13 VN.n12 161.3
R1524 VN.n11 VN.n2 161.3
R1525 VN.n10 VN.n9 161.3
R1526 VN.n8 VN.n3 161.3
R1527 VN.n7 VN.n6 161.3
R1528 VN.n23 VN.t1 75.2141
R1529 VN.n5 VN.t5 75.2141
R1530 VN.n17 VN.n0 73.5231
R1531 VN.n35 VN.n18 73.5231
R1532 VN.n5 VN.n4 62.2204
R1533 VN.n23 VN.n22 62.2204
R1534 VN VN.n35 46.7746
R1535 VN.n13 VN.n2 44.9365
R1536 VN.n31 VN.n20 44.9365
R1537 VN.n4 VN.t3 41.9907
R1538 VN.n0 VN.t0 41.9907
R1539 VN.n22 VN.t2 41.9907
R1540 VN.n18 VN.t4 41.9907
R1541 VN.n9 VN.n2 36.2176
R1542 VN.n27 VN.n20 36.2176
R1543 VN.n8 VN.n7 24.5923
R1544 VN.n9 VN.n8 24.5923
R1545 VN.n14 VN.n13 24.5923
R1546 VN.n15 VN.n14 24.5923
R1547 VN.n27 VN.n26 24.5923
R1548 VN.n26 VN.n25 24.5923
R1549 VN.n33 VN.n32 24.5923
R1550 VN.n32 VN.n31 24.5923
R1551 VN.n15 VN.n0 16.7229
R1552 VN.n33 VN.n18 16.7229
R1553 VN.n7 VN.n4 12.2964
R1554 VN.n25 VN.n22 12.2964
R1555 VN.n24 VN.n23 4.04954
R1556 VN.n6 VN.n5 4.04954
R1557 VN.n35 VN.n34 0.354861
R1558 VN.n17 VN.n16 0.354861
R1559 VN VN.n17 0.267071
R1560 VN.n34 VN.n19 0.189894
R1561 VN.n30 VN.n19 0.189894
R1562 VN.n30 VN.n29 0.189894
R1563 VN.n29 VN.n28 0.189894
R1564 VN.n28 VN.n21 0.189894
R1565 VN.n24 VN.n21 0.189894
R1566 VN.n6 VN.n3 0.189894
R1567 VN.n10 VN.n3 0.189894
R1568 VN.n11 VN.n10 0.189894
R1569 VN.n12 VN.n11 0.189894
R1570 VN.n12 VN.n1 0.189894
R1571 VN.n16 VN.n1 0.189894
R1572 VDD2.n1 VDD2.t0 74.3973
R1573 VDD2.n2 VDD2.t1 72.1317
R1574 VDD2.n1 VDD2.n0 69.3639
R1575 VDD2 VDD2.n3 69.3611
R1576 VDD2.n2 VDD2.n1 38.67
R1577 VDD2.n3 VDD2.t3 3.48642
R1578 VDD2.n3 VDD2.t4 3.48642
R1579 VDD2.n0 VDD2.t2 3.48642
R1580 VDD2.n0 VDD2.t5 3.48642
R1581 VDD2 VDD2.n2 2.37981
C0 VDD2 VN 3.52321f
C1 VN VTAIL 4.31303f
C2 VDD2 VP 0.514066f
C3 VP VTAIL 4.32721f
C4 VDD2 VTAIL 5.86494f
C5 VN VDD1 0.151845f
C6 VDD1 VP 3.88327f
C7 VDD2 VDD1 1.66292f
C8 VDD1 VTAIL 5.80791f
C9 VN VP 6.39236f
C10 VDD2 B 5.368536f
C11 VDD1 B 5.720341f
C12 VTAIL B 5.297209f
C13 VN B 14.20774f
C14 VP B 12.899021f
C15 VDD2.t0 B 1.0486f
C16 VDD2.t2 B 0.098456f
C17 VDD2.t5 B 0.098456f
C18 VDD2.n0 B 0.820457f
C19 VDD2.n1 B 2.447f
C20 VDD2.t1 B 1.03661f
C21 VDD2.n2 B 2.16399f
C22 VDD2.t3 B 0.098456f
C23 VDD2.t4 B 0.098456f
C24 VDD2.n3 B 0.820428f
C25 VN.t0 B 1.1408f
C26 VN.n0 B 0.518605f
C27 VN.n1 B 0.023354f
C28 VN.n2 B 0.019473f
C29 VN.n3 B 0.023354f
C30 VN.t3 B 1.1408f
C31 VN.n4 B 0.50233f
C32 VN.t5 B 1.40231f
C33 VN.n5 B 0.47891f
C34 VN.n6 B 0.272305f
C35 VN.n7 B 0.032618f
C36 VN.n8 B 0.043308f
C37 VN.n9 B 0.046877f
C38 VN.n10 B 0.023354f
C39 VN.n11 B 0.023354f
C40 VN.n12 B 0.023354f
C41 VN.n13 B 0.044857f
C42 VN.n14 B 0.043308f
C43 VN.n15 B 0.036467f
C44 VN.n16 B 0.037687f
C45 VN.n17 B 0.054188f
C46 VN.t4 B 1.1408f
C47 VN.n18 B 0.518605f
C48 VN.n19 B 0.023354f
C49 VN.n20 B 0.019473f
C50 VN.n21 B 0.023354f
C51 VN.t2 B 1.1408f
C52 VN.n22 B 0.50233f
C53 VN.t1 B 1.40231f
C54 VN.n23 B 0.47891f
C55 VN.n24 B 0.272305f
C56 VN.n25 B 0.032618f
C57 VN.n26 B 0.043308f
C58 VN.n27 B 0.046877f
C59 VN.n28 B 0.023354f
C60 VN.n29 B 0.023354f
C61 VN.n30 B 0.023354f
C62 VN.n31 B 0.044857f
C63 VN.n32 B 0.043308f
C64 VN.n33 B 0.036467f
C65 VN.n34 B 0.037687f
C66 VN.n35 B 1.20691f
C67 VTAIL.t5 B 0.126712f
C68 VTAIL.t1 B 0.126712f
C69 VTAIL.n0 B 0.978502f
C70 VTAIL.n1 B 0.519815f
C71 VTAIL.t10 B 1.24881f
C72 VTAIL.n2 B 0.800932f
C73 VTAIL.t9 B 0.126712f
C74 VTAIL.t8 B 0.126712f
C75 VTAIL.n3 B 0.978502f
C76 VTAIL.n4 B 1.93409f
C77 VTAIL.t0 B 0.126712f
C78 VTAIL.t2 B 0.126712f
C79 VTAIL.n5 B 0.978508f
C80 VTAIL.n6 B 1.93409f
C81 VTAIL.t3 B 1.24882f
C82 VTAIL.n7 B 0.800927f
C83 VTAIL.t7 B 0.126712f
C84 VTAIL.t11 B 0.126712f
C85 VTAIL.n8 B 0.978508f
C86 VTAIL.n9 B 0.725656f
C87 VTAIL.t6 B 1.24881f
C88 VTAIL.n10 B 1.72784f
C89 VTAIL.t4 B 1.24881f
C90 VTAIL.n11 B 1.65217f
C91 VDD1.t5 B 1.07367f
C92 VDD1.t3 B 1.07282f
C93 VDD1.t0 B 0.10073f
C94 VDD1.t4 B 0.10073f
C95 VDD1.n0 B 0.839407f
C96 VDD1.n1 B 2.62464f
C97 VDD1.t2 B 0.10073f
C98 VDD1.t1 B 0.10073f
C99 VDD1.n2 B 0.834575f
C100 VDD1.n3 B 2.23048f
C101 VP.t1 B 1.17565f
C102 VP.n0 B 0.534449f
C103 VP.n1 B 0.024068f
C104 VP.n2 B 0.020067f
C105 VP.n3 B 0.024068f
C106 VP.t3 B 1.17565f
C107 VP.n4 B 0.43835f
C108 VP.n5 B 0.024068f
C109 VP.n6 B 0.020067f
C110 VP.n7 B 0.024068f
C111 VP.t2 B 1.17565f
C112 VP.n8 B 0.534449f
C113 VP.t5 B 1.17565f
C114 VP.n9 B 0.534449f
C115 VP.n10 B 0.024068f
C116 VP.n11 B 0.020067f
C117 VP.n12 B 0.024068f
C118 VP.t0 B 1.17565f
C119 VP.n13 B 0.517677f
C120 VP.t4 B 1.44515f
C121 VP.n14 B 0.493543f
C122 VP.n15 B 0.280624f
C123 VP.n16 B 0.033615f
C124 VP.n17 B 0.044632f
C125 VP.n18 B 0.048309f
C126 VP.n19 B 0.024068f
C127 VP.n20 B 0.024068f
C128 VP.n21 B 0.024068f
C129 VP.n22 B 0.046228f
C130 VP.n23 B 0.044632f
C131 VP.n24 B 0.037581f
C132 VP.n25 B 0.038839f
C133 VP.n26 B 1.2337f
C134 VP.n27 B 1.25231f
C135 VP.n28 B 0.038839f
C136 VP.n29 B 0.037581f
C137 VP.n30 B 0.044632f
C138 VP.n31 B 0.046228f
C139 VP.n32 B 0.024068f
C140 VP.n33 B 0.024068f
C141 VP.n34 B 0.024068f
C142 VP.n35 B 0.048309f
C143 VP.n36 B 0.044632f
C144 VP.n37 B 0.033615f
C145 VP.n38 B 0.024068f
C146 VP.n39 B 0.024068f
C147 VP.n40 B 0.033615f
C148 VP.n41 B 0.044632f
C149 VP.n42 B 0.048309f
C150 VP.n43 B 0.024068f
C151 VP.n44 B 0.024068f
C152 VP.n45 B 0.024068f
C153 VP.n46 B 0.046228f
C154 VP.n47 B 0.044632f
C155 VP.n48 B 0.037581f
C156 VP.n49 B 0.038839f
C157 VP.n50 B 0.055844f
.ends

