* NGSPICE file created from diff_pair_sample_0112.ext - technology: sky130A

.subckt diff_pair_sample_0112 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X1 B.t11 B.t9 B.t10 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=0 ps=0 w=14.34 l=2.61
X2 VTAIL.t8 VN.t0 VDD2.t9 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X3 VDD2.t8 VN.t1 VTAIL.t7 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=2.3661 ps=14.67 w=14.34 l=2.61
X4 B.t8 B.t6 B.t7 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=0 ps=0 w=14.34 l=2.61
X5 VDD1.t8 VP.t1 VTAIL.t17 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=2.3661 ps=14.67 w=14.34 l=2.61
X6 VDD2.t7 VN.t2 VTAIL.t6 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=5.5926 ps=29.46 w=14.34 l=2.61
X7 VTAIL.t13 VP.t2 VDD1.t7 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X8 VDD2.t6 VN.t3 VTAIL.t0 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=5.5926 ps=29.46 w=14.34 l=2.61
X9 VDD1.t6 VP.t3 VTAIL.t12 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=5.5926 ps=29.46 w=14.34 l=2.61
X10 VDD2.t5 VN.t4 VTAIL.t5 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=2.3661 ps=14.67 w=14.34 l=2.61
X11 VTAIL.t4 VN.t5 VDD2.t4 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X12 VDD1.t5 VP.t4 VTAIL.t10 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=5.5926 ps=29.46 w=14.34 l=2.61
X13 VTAIL.t3 VN.t6 VDD2.t3 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X14 B.t5 B.t3 B.t4 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=0 ps=0 w=14.34 l=2.61
X15 VDD1.t4 VP.t5 VTAIL.t18 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=2.3661 ps=14.67 w=14.34 l=2.61
X16 B.t2 B.t0 B.t1 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=5.5926 pd=29.46 as=0 ps=0 w=14.34 l=2.61
X17 VTAIL.t15 VP.t6 VDD1.t3 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X18 VTAIL.t16 VP.t7 VDD1.t2 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X19 VTAIL.t9 VP.t8 VDD1.t1 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X20 VDD2.t2 VN.t7 VTAIL.t2 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X21 VDD1.t0 VP.t9 VTAIL.t14 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X22 VTAIL.t19 VN.t8 VDD2.t1 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
X23 VDD2.t0 VN.t9 VTAIL.t1 w_n4498_n3836# sky130_fd_pr__pfet_01v8 ad=2.3661 pd=14.67 as=2.3661 ps=14.67 w=14.34 l=2.61
R0 VP.n24 VP.t5 164.99
R1 VP.n25 VP.n22 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n21 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n20 161.3
R6 VP.n33 VP.n32 161.3
R7 VP.n35 VP.n19 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n18 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n17 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n15 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n14 161.3
R17 VP.n51 VP.n50 161.3
R18 VP.n52 VP.n13 161.3
R19 VP.n94 VP.n0 161.3
R20 VP.n93 VP.n92 161.3
R21 VP.n91 VP.n1 161.3
R22 VP.n90 VP.n89 161.3
R23 VP.n88 VP.n2 161.3
R24 VP.n87 VP.n86 161.3
R25 VP.n85 VP.n84 161.3
R26 VP.n83 VP.n4 161.3
R27 VP.n82 VP.n81 161.3
R28 VP.n80 VP.n5 161.3
R29 VP.n79 VP.n78 161.3
R30 VP.n77 VP.n6 161.3
R31 VP.n75 VP.n74 161.3
R32 VP.n73 VP.n7 161.3
R33 VP.n72 VP.n71 161.3
R34 VP.n70 VP.n8 161.3
R35 VP.n69 VP.n68 161.3
R36 VP.n67 VP.n9 161.3
R37 VP.n66 VP.n65 161.3
R38 VP.n63 VP.n10 161.3
R39 VP.n62 VP.n61 161.3
R40 VP.n60 VP.n11 161.3
R41 VP.n59 VP.n58 161.3
R42 VP.n57 VP.n12 161.3
R43 VP.n56 VP.t1 132.411
R44 VP.n64 VP.t2 132.411
R45 VP.n76 VP.t0 132.411
R46 VP.n3 VP.t8 132.411
R47 VP.n95 VP.t3 132.411
R48 VP.n53 VP.t4 132.411
R49 VP.n16 VP.t6 132.411
R50 VP.n34 VP.t9 132.411
R51 VP.n23 VP.t7 132.411
R52 VP.n56 VP.n55 104.514
R53 VP.n96 VP.n95 104.514
R54 VP.n54 VP.n53 104.514
R55 VP.n24 VP.n23 63.1649
R56 VP.n71 VP.n70 56.5617
R57 VP.n82 VP.n5 56.5617
R58 VP.n40 VP.n18 56.5617
R59 VP.n29 VP.n28 56.5617
R60 VP.n62 VP.n11 56.0773
R61 VP.n89 VP.n1 56.0773
R62 VP.n47 VP.n14 56.0773
R63 VP.n55 VP.n54 54.9087
R64 VP.n63 VP.n62 25.0767
R65 VP.n89 VP.n88 25.0767
R66 VP.n47 VP.n46 25.0767
R67 VP.n58 VP.n57 24.5923
R68 VP.n58 VP.n11 24.5923
R69 VP.n65 VP.n63 24.5923
R70 VP.n69 VP.n9 24.5923
R71 VP.n70 VP.n69 24.5923
R72 VP.n71 VP.n7 24.5923
R73 VP.n75 VP.n7 24.5923
R74 VP.n78 VP.n77 24.5923
R75 VP.n78 VP.n5 24.5923
R76 VP.n83 VP.n82 24.5923
R77 VP.n84 VP.n83 24.5923
R78 VP.n88 VP.n87 24.5923
R79 VP.n93 VP.n1 24.5923
R80 VP.n94 VP.n93 24.5923
R81 VP.n51 VP.n14 24.5923
R82 VP.n52 VP.n51 24.5923
R83 VP.n41 VP.n40 24.5923
R84 VP.n42 VP.n41 24.5923
R85 VP.n46 VP.n45 24.5923
R86 VP.n29 VP.n20 24.5923
R87 VP.n33 VP.n20 24.5923
R88 VP.n36 VP.n35 24.5923
R89 VP.n36 VP.n18 24.5923
R90 VP.n27 VP.n22 24.5923
R91 VP.n28 VP.n27 24.5923
R92 VP.n65 VP.n64 15.2474
R93 VP.n87 VP.n3 15.2474
R94 VP.n45 VP.n16 15.2474
R95 VP.n76 VP.n75 12.2964
R96 VP.n77 VP.n76 12.2964
R97 VP.n34 VP.n33 12.2964
R98 VP.n35 VP.n34 12.2964
R99 VP.n64 VP.n9 9.3454
R100 VP.n84 VP.n3 9.3454
R101 VP.n42 VP.n16 9.3454
R102 VP.n23 VP.n22 9.3454
R103 VP.n25 VP.n24 7.05922
R104 VP.n57 VP.n56 6.39438
R105 VP.n95 VP.n94 6.39438
R106 VP.n53 VP.n52 6.39438
R107 VP.n54 VP.n13 0.278335
R108 VP.n55 VP.n12 0.278335
R109 VP.n96 VP.n0 0.278335
R110 VP.n26 VP.n25 0.189894
R111 VP.n26 VP.n21 0.189894
R112 VP.n30 VP.n21 0.189894
R113 VP.n31 VP.n30 0.189894
R114 VP.n32 VP.n31 0.189894
R115 VP.n32 VP.n19 0.189894
R116 VP.n37 VP.n19 0.189894
R117 VP.n38 VP.n37 0.189894
R118 VP.n39 VP.n38 0.189894
R119 VP.n39 VP.n17 0.189894
R120 VP.n43 VP.n17 0.189894
R121 VP.n44 VP.n43 0.189894
R122 VP.n44 VP.n15 0.189894
R123 VP.n48 VP.n15 0.189894
R124 VP.n49 VP.n48 0.189894
R125 VP.n50 VP.n49 0.189894
R126 VP.n50 VP.n13 0.189894
R127 VP.n59 VP.n12 0.189894
R128 VP.n60 VP.n59 0.189894
R129 VP.n61 VP.n60 0.189894
R130 VP.n61 VP.n10 0.189894
R131 VP.n66 VP.n10 0.189894
R132 VP.n67 VP.n66 0.189894
R133 VP.n68 VP.n67 0.189894
R134 VP.n68 VP.n8 0.189894
R135 VP.n72 VP.n8 0.189894
R136 VP.n73 VP.n72 0.189894
R137 VP.n74 VP.n73 0.189894
R138 VP.n74 VP.n6 0.189894
R139 VP.n79 VP.n6 0.189894
R140 VP.n80 VP.n79 0.189894
R141 VP.n81 VP.n80 0.189894
R142 VP.n81 VP.n4 0.189894
R143 VP.n85 VP.n4 0.189894
R144 VP.n86 VP.n85 0.189894
R145 VP.n86 VP.n2 0.189894
R146 VP.n90 VP.n2 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n92 VP.n91 0.189894
R149 VP.n92 VP.n0 0.189894
R150 VP VP.n96 0.153485
R151 VTAIL.n11 VTAIL.t0 57.7941
R152 VTAIL.n17 VTAIL.t6 57.794
R153 VTAIL.n2 VTAIL.t12 57.794
R154 VTAIL.n16 VTAIL.t10 57.794
R155 VTAIL.n15 VTAIL.n14 55.5274
R156 VTAIL.n13 VTAIL.n12 55.5274
R157 VTAIL.n10 VTAIL.n9 55.5274
R158 VTAIL.n8 VTAIL.n7 55.5274
R159 VTAIL.n19 VTAIL.n18 55.5272
R160 VTAIL.n1 VTAIL.n0 55.5272
R161 VTAIL.n4 VTAIL.n3 55.5272
R162 VTAIL.n6 VTAIL.n5 55.5272
R163 VTAIL.n8 VTAIL.n6 29.7979
R164 VTAIL.n17 VTAIL.n16 27.2634
R165 VTAIL.n10 VTAIL.n8 2.53498
R166 VTAIL.n11 VTAIL.n10 2.53498
R167 VTAIL.n15 VTAIL.n13 2.53498
R168 VTAIL.n16 VTAIL.n15 2.53498
R169 VTAIL.n6 VTAIL.n4 2.53498
R170 VTAIL.n4 VTAIL.n2 2.53498
R171 VTAIL.n19 VTAIL.n17 2.53498
R172 VTAIL.n18 VTAIL.t1 2.26724
R173 VTAIL.n18 VTAIL.t8 2.26724
R174 VTAIL.n0 VTAIL.t7 2.26724
R175 VTAIL.n0 VTAIL.t4 2.26724
R176 VTAIL.n3 VTAIL.t11 2.26724
R177 VTAIL.n3 VTAIL.t9 2.26724
R178 VTAIL.n5 VTAIL.t17 2.26724
R179 VTAIL.n5 VTAIL.t13 2.26724
R180 VTAIL.n14 VTAIL.t14 2.26724
R181 VTAIL.n14 VTAIL.t15 2.26724
R182 VTAIL.n12 VTAIL.t18 2.26724
R183 VTAIL.n12 VTAIL.t16 2.26724
R184 VTAIL.n9 VTAIL.t2 2.26724
R185 VTAIL.n9 VTAIL.t3 2.26724
R186 VTAIL.n7 VTAIL.t5 2.26724
R187 VTAIL.n7 VTAIL.t19 2.26724
R188 VTAIL VTAIL.n1 1.95955
R189 VTAIL.n13 VTAIL.n11 1.73757
R190 VTAIL.n2 VTAIL.n1 1.73757
R191 VTAIL VTAIL.n19 0.575931
R192 VDD1.n1 VDD1.t4 77.0074
R193 VDD1.n3 VDD1.t8 77.0073
R194 VDD1.n5 VDD1.n4 74.0515
R195 VDD1.n1 VDD1.n0 72.2062
R196 VDD1.n7 VDD1.n6 72.206
R197 VDD1.n3 VDD1.n2 72.206
R198 VDD1.n7 VDD1.n5 49.9664
R199 VDD1.n6 VDD1.t3 2.26724
R200 VDD1.n6 VDD1.t5 2.26724
R201 VDD1.n0 VDD1.t2 2.26724
R202 VDD1.n0 VDD1.t0 2.26724
R203 VDD1.n4 VDD1.t1 2.26724
R204 VDD1.n4 VDD1.t6 2.26724
R205 VDD1.n2 VDD1.t7 2.26724
R206 VDD1.n2 VDD1.t9 2.26724
R207 VDD1 VDD1.n7 1.84317
R208 VDD1 VDD1.n1 0.69231
R209 VDD1.n5 VDD1.n3 0.578775
R210 B.n671 B.n90 585
R211 B.n673 B.n672 585
R212 B.n674 B.n89 585
R213 B.n676 B.n675 585
R214 B.n677 B.n88 585
R215 B.n679 B.n678 585
R216 B.n680 B.n87 585
R217 B.n682 B.n681 585
R218 B.n683 B.n86 585
R219 B.n685 B.n684 585
R220 B.n686 B.n85 585
R221 B.n688 B.n687 585
R222 B.n689 B.n84 585
R223 B.n691 B.n690 585
R224 B.n692 B.n83 585
R225 B.n694 B.n693 585
R226 B.n695 B.n82 585
R227 B.n697 B.n696 585
R228 B.n698 B.n81 585
R229 B.n700 B.n699 585
R230 B.n701 B.n80 585
R231 B.n703 B.n702 585
R232 B.n704 B.n79 585
R233 B.n706 B.n705 585
R234 B.n707 B.n78 585
R235 B.n709 B.n708 585
R236 B.n710 B.n77 585
R237 B.n712 B.n711 585
R238 B.n713 B.n76 585
R239 B.n715 B.n714 585
R240 B.n716 B.n75 585
R241 B.n718 B.n717 585
R242 B.n719 B.n74 585
R243 B.n721 B.n720 585
R244 B.n722 B.n73 585
R245 B.n724 B.n723 585
R246 B.n725 B.n72 585
R247 B.n727 B.n726 585
R248 B.n728 B.n71 585
R249 B.n730 B.n729 585
R250 B.n731 B.n70 585
R251 B.n733 B.n732 585
R252 B.n734 B.n69 585
R253 B.n736 B.n735 585
R254 B.n737 B.n68 585
R255 B.n739 B.n738 585
R256 B.n740 B.n67 585
R257 B.n742 B.n741 585
R258 B.n743 B.n64 585
R259 B.n746 B.n745 585
R260 B.n747 B.n63 585
R261 B.n749 B.n748 585
R262 B.n750 B.n62 585
R263 B.n752 B.n751 585
R264 B.n753 B.n61 585
R265 B.n755 B.n754 585
R266 B.n756 B.n57 585
R267 B.n758 B.n757 585
R268 B.n759 B.n56 585
R269 B.n761 B.n760 585
R270 B.n762 B.n55 585
R271 B.n764 B.n763 585
R272 B.n765 B.n54 585
R273 B.n767 B.n766 585
R274 B.n768 B.n53 585
R275 B.n770 B.n769 585
R276 B.n771 B.n52 585
R277 B.n773 B.n772 585
R278 B.n774 B.n51 585
R279 B.n776 B.n775 585
R280 B.n777 B.n50 585
R281 B.n779 B.n778 585
R282 B.n780 B.n49 585
R283 B.n782 B.n781 585
R284 B.n783 B.n48 585
R285 B.n785 B.n784 585
R286 B.n786 B.n47 585
R287 B.n788 B.n787 585
R288 B.n789 B.n46 585
R289 B.n791 B.n790 585
R290 B.n792 B.n45 585
R291 B.n794 B.n793 585
R292 B.n795 B.n44 585
R293 B.n797 B.n796 585
R294 B.n798 B.n43 585
R295 B.n800 B.n799 585
R296 B.n801 B.n42 585
R297 B.n803 B.n802 585
R298 B.n804 B.n41 585
R299 B.n806 B.n805 585
R300 B.n807 B.n40 585
R301 B.n809 B.n808 585
R302 B.n810 B.n39 585
R303 B.n812 B.n811 585
R304 B.n813 B.n38 585
R305 B.n815 B.n814 585
R306 B.n816 B.n37 585
R307 B.n818 B.n817 585
R308 B.n819 B.n36 585
R309 B.n821 B.n820 585
R310 B.n822 B.n35 585
R311 B.n824 B.n823 585
R312 B.n825 B.n34 585
R313 B.n827 B.n826 585
R314 B.n828 B.n33 585
R315 B.n830 B.n829 585
R316 B.n831 B.n32 585
R317 B.n670 B.n669 585
R318 B.n668 B.n91 585
R319 B.n667 B.n666 585
R320 B.n665 B.n92 585
R321 B.n664 B.n663 585
R322 B.n662 B.n93 585
R323 B.n661 B.n660 585
R324 B.n659 B.n94 585
R325 B.n658 B.n657 585
R326 B.n656 B.n95 585
R327 B.n655 B.n654 585
R328 B.n653 B.n96 585
R329 B.n652 B.n651 585
R330 B.n650 B.n97 585
R331 B.n649 B.n648 585
R332 B.n647 B.n98 585
R333 B.n646 B.n645 585
R334 B.n644 B.n99 585
R335 B.n643 B.n642 585
R336 B.n641 B.n100 585
R337 B.n640 B.n639 585
R338 B.n638 B.n101 585
R339 B.n637 B.n636 585
R340 B.n635 B.n102 585
R341 B.n634 B.n633 585
R342 B.n632 B.n103 585
R343 B.n631 B.n630 585
R344 B.n629 B.n104 585
R345 B.n628 B.n627 585
R346 B.n626 B.n105 585
R347 B.n625 B.n624 585
R348 B.n623 B.n106 585
R349 B.n622 B.n621 585
R350 B.n620 B.n107 585
R351 B.n619 B.n618 585
R352 B.n617 B.n108 585
R353 B.n616 B.n615 585
R354 B.n614 B.n109 585
R355 B.n613 B.n612 585
R356 B.n611 B.n110 585
R357 B.n610 B.n609 585
R358 B.n608 B.n111 585
R359 B.n607 B.n606 585
R360 B.n605 B.n112 585
R361 B.n604 B.n603 585
R362 B.n602 B.n113 585
R363 B.n601 B.n600 585
R364 B.n599 B.n114 585
R365 B.n598 B.n597 585
R366 B.n596 B.n115 585
R367 B.n595 B.n594 585
R368 B.n593 B.n116 585
R369 B.n592 B.n591 585
R370 B.n590 B.n117 585
R371 B.n589 B.n588 585
R372 B.n587 B.n118 585
R373 B.n586 B.n585 585
R374 B.n584 B.n119 585
R375 B.n583 B.n582 585
R376 B.n581 B.n120 585
R377 B.n580 B.n579 585
R378 B.n578 B.n121 585
R379 B.n577 B.n576 585
R380 B.n575 B.n122 585
R381 B.n574 B.n573 585
R382 B.n572 B.n123 585
R383 B.n571 B.n570 585
R384 B.n569 B.n124 585
R385 B.n568 B.n567 585
R386 B.n566 B.n125 585
R387 B.n565 B.n564 585
R388 B.n563 B.n126 585
R389 B.n562 B.n561 585
R390 B.n560 B.n127 585
R391 B.n559 B.n558 585
R392 B.n557 B.n128 585
R393 B.n556 B.n555 585
R394 B.n554 B.n129 585
R395 B.n553 B.n552 585
R396 B.n551 B.n130 585
R397 B.n550 B.n549 585
R398 B.n548 B.n131 585
R399 B.n547 B.n546 585
R400 B.n545 B.n132 585
R401 B.n544 B.n543 585
R402 B.n542 B.n133 585
R403 B.n541 B.n540 585
R404 B.n539 B.n134 585
R405 B.n538 B.n537 585
R406 B.n536 B.n135 585
R407 B.n535 B.n534 585
R408 B.n533 B.n136 585
R409 B.n532 B.n531 585
R410 B.n530 B.n137 585
R411 B.n529 B.n528 585
R412 B.n527 B.n138 585
R413 B.n526 B.n525 585
R414 B.n524 B.n139 585
R415 B.n523 B.n522 585
R416 B.n521 B.n140 585
R417 B.n520 B.n519 585
R418 B.n518 B.n141 585
R419 B.n517 B.n516 585
R420 B.n515 B.n142 585
R421 B.n514 B.n513 585
R422 B.n512 B.n143 585
R423 B.n511 B.n510 585
R424 B.n509 B.n144 585
R425 B.n508 B.n507 585
R426 B.n506 B.n145 585
R427 B.n505 B.n504 585
R428 B.n503 B.n146 585
R429 B.n502 B.n501 585
R430 B.n500 B.n147 585
R431 B.n499 B.n498 585
R432 B.n497 B.n148 585
R433 B.n496 B.n495 585
R434 B.n494 B.n149 585
R435 B.n493 B.n492 585
R436 B.n491 B.n150 585
R437 B.n490 B.n489 585
R438 B.n325 B.n206 585
R439 B.n327 B.n326 585
R440 B.n328 B.n205 585
R441 B.n330 B.n329 585
R442 B.n331 B.n204 585
R443 B.n333 B.n332 585
R444 B.n334 B.n203 585
R445 B.n336 B.n335 585
R446 B.n337 B.n202 585
R447 B.n339 B.n338 585
R448 B.n340 B.n201 585
R449 B.n342 B.n341 585
R450 B.n343 B.n200 585
R451 B.n345 B.n344 585
R452 B.n346 B.n199 585
R453 B.n348 B.n347 585
R454 B.n349 B.n198 585
R455 B.n351 B.n350 585
R456 B.n352 B.n197 585
R457 B.n354 B.n353 585
R458 B.n355 B.n196 585
R459 B.n357 B.n356 585
R460 B.n358 B.n195 585
R461 B.n360 B.n359 585
R462 B.n361 B.n194 585
R463 B.n363 B.n362 585
R464 B.n364 B.n193 585
R465 B.n366 B.n365 585
R466 B.n367 B.n192 585
R467 B.n369 B.n368 585
R468 B.n370 B.n191 585
R469 B.n372 B.n371 585
R470 B.n373 B.n190 585
R471 B.n375 B.n374 585
R472 B.n376 B.n189 585
R473 B.n378 B.n377 585
R474 B.n379 B.n188 585
R475 B.n381 B.n380 585
R476 B.n382 B.n187 585
R477 B.n384 B.n383 585
R478 B.n385 B.n186 585
R479 B.n387 B.n386 585
R480 B.n388 B.n185 585
R481 B.n390 B.n389 585
R482 B.n391 B.n184 585
R483 B.n393 B.n392 585
R484 B.n394 B.n183 585
R485 B.n396 B.n395 585
R486 B.n397 B.n180 585
R487 B.n400 B.n399 585
R488 B.n401 B.n179 585
R489 B.n403 B.n402 585
R490 B.n404 B.n178 585
R491 B.n406 B.n405 585
R492 B.n407 B.n177 585
R493 B.n409 B.n408 585
R494 B.n410 B.n176 585
R495 B.n415 B.n414 585
R496 B.n416 B.n175 585
R497 B.n418 B.n417 585
R498 B.n419 B.n174 585
R499 B.n421 B.n420 585
R500 B.n422 B.n173 585
R501 B.n424 B.n423 585
R502 B.n425 B.n172 585
R503 B.n427 B.n426 585
R504 B.n428 B.n171 585
R505 B.n430 B.n429 585
R506 B.n431 B.n170 585
R507 B.n433 B.n432 585
R508 B.n434 B.n169 585
R509 B.n436 B.n435 585
R510 B.n437 B.n168 585
R511 B.n439 B.n438 585
R512 B.n440 B.n167 585
R513 B.n442 B.n441 585
R514 B.n443 B.n166 585
R515 B.n445 B.n444 585
R516 B.n446 B.n165 585
R517 B.n448 B.n447 585
R518 B.n449 B.n164 585
R519 B.n451 B.n450 585
R520 B.n452 B.n163 585
R521 B.n454 B.n453 585
R522 B.n455 B.n162 585
R523 B.n457 B.n456 585
R524 B.n458 B.n161 585
R525 B.n460 B.n459 585
R526 B.n461 B.n160 585
R527 B.n463 B.n462 585
R528 B.n464 B.n159 585
R529 B.n466 B.n465 585
R530 B.n467 B.n158 585
R531 B.n469 B.n468 585
R532 B.n470 B.n157 585
R533 B.n472 B.n471 585
R534 B.n473 B.n156 585
R535 B.n475 B.n474 585
R536 B.n476 B.n155 585
R537 B.n478 B.n477 585
R538 B.n479 B.n154 585
R539 B.n481 B.n480 585
R540 B.n482 B.n153 585
R541 B.n484 B.n483 585
R542 B.n485 B.n152 585
R543 B.n487 B.n486 585
R544 B.n488 B.n151 585
R545 B.n324 B.n323 585
R546 B.n322 B.n207 585
R547 B.n321 B.n320 585
R548 B.n319 B.n208 585
R549 B.n318 B.n317 585
R550 B.n316 B.n209 585
R551 B.n315 B.n314 585
R552 B.n313 B.n210 585
R553 B.n312 B.n311 585
R554 B.n310 B.n211 585
R555 B.n309 B.n308 585
R556 B.n307 B.n212 585
R557 B.n306 B.n305 585
R558 B.n304 B.n213 585
R559 B.n303 B.n302 585
R560 B.n301 B.n214 585
R561 B.n300 B.n299 585
R562 B.n298 B.n215 585
R563 B.n297 B.n296 585
R564 B.n295 B.n216 585
R565 B.n294 B.n293 585
R566 B.n292 B.n217 585
R567 B.n291 B.n290 585
R568 B.n289 B.n218 585
R569 B.n288 B.n287 585
R570 B.n286 B.n219 585
R571 B.n285 B.n284 585
R572 B.n283 B.n220 585
R573 B.n282 B.n281 585
R574 B.n280 B.n221 585
R575 B.n279 B.n278 585
R576 B.n277 B.n222 585
R577 B.n276 B.n275 585
R578 B.n274 B.n223 585
R579 B.n273 B.n272 585
R580 B.n271 B.n224 585
R581 B.n270 B.n269 585
R582 B.n268 B.n225 585
R583 B.n267 B.n266 585
R584 B.n265 B.n226 585
R585 B.n264 B.n263 585
R586 B.n262 B.n227 585
R587 B.n261 B.n260 585
R588 B.n259 B.n228 585
R589 B.n258 B.n257 585
R590 B.n256 B.n229 585
R591 B.n255 B.n254 585
R592 B.n253 B.n230 585
R593 B.n252 B.n251 585
R594 B.n250 B.n231 585
R595 B.n249 B.n248 585
R596 B.n247 B.n232 585
R597 B.n246 B.n245 585
R598 B.n244 B.n233 585
R599 B.n243 B.n242 585
R600 B.n241 B.n234 585
R601 B.n240 B.n239 585
R602 B.n238 B.n235 585
R603 B.n237 B.n236 585
R604 B.n2 B.n0 585
R605 B.n921 B.n1 585
R606 B.n920 B.n919 585
R607 B.n918 B.n3 585
R608 B.n917 B.n916 585
R609 B.n915 B.n4 585
R610 B.n914 B.n913 585
R611 B.n912 B.n5 585
R612 B.n911 B.n910 585
R613 B.n909 B.n6 585
R614 B.n908 B.n907 585
R615 B.n906 B.n7 585
R616 B.n905 B.n904 585
R617 B.n903 B.n8 585
R618 B.n902 B.n901 585
R619 B.n900 B.n9 585
R620 B.n899 B.n898 585
R621 B.n897 B.n10 585
R622 B.n896 B.n895 585
R623 B.n894 B.n11 585
R624 B.n893 B.n892 585
R625 B.n891 B.n12 585
R626 B.n890 B.n889 585
R627 B.n888 B.n13 585
R628 B.n887 B.n886 585
R629 B.n885 B.n14 585
R630 B.n884 B.n883 585
R631 B.n882 B.n15 585
R632 B.n881 B.n880 585
R633 B.n879 B.n16 585
R634 B.n878 B.n877 585
R635 B.n876 B.n17 585
R636 B.n875 B.n874 585
R637 B.n873 B.n18 585
R638 B.n872 B.n871 585
R639 B.n870 B.n19 585
R640 B.n869 B.n868 585
R641 B.n867 B.n20 585
R642 B.n866 B.n865 585
R643 B.n864 B.n21 585
R644 B.n863 B.n862 585
R645 B.n861 B.n22 585
R646 B.n860 B.n859 585
R647 B.n858 B.n23 585
R648 B.n857 B.n856 585
R649 B.n855 B.n24 585
R650 B.n854 B.n853 585
R651 B.n852 B.n25 585
R652 B.n851 B.n850 585
R653 B.n849 B.n26 585
R654 B.n848 B.n847 585
R655 B.n846 B.n27 585
R656 B.n845 B.n844 585
R657 B.n843 B.n28 585
R658 B.n842 B.n841 585
R659 B.n840 B.n29 585
R660 B.n839 B.n838 585
R661 B.n837 B.n30 585
R662 B.n836 B.n835 585
R663 B.n834 B.n31 585
R664 B.n833 B.n832 585
R665 B.n923 B.n922 585
R666 B.n323 B.n206 463.671
R667 B.n832 B.n831 463.671
R668 B.n489 B.n488 463.671
R669 B.n669 B.n90 463.671
R670 B.n411 B.t0 340.474
R671 B.n181 B.t9 340.474
R672 B.n58 B.t6 340.474
R673 B.n65 B.t3 340.474
R674 B.n411 B.t2 164.843
R675 B.n65 B.t4 164.843
R676 B.n181 B.t11 164.825
R677 B.n58 B.t7 164.825
R678 B.n323 B.n322 163.367
R679 B.n322 B.n321 163.367
R680 B.n321 B.n208 163.367
R681 B.n317 B.n208 163.367
R682 B.n317 B.n316 163.367
R683 B.n316 B.n315 163.367
R684 B.n315 B.n210 163.367
R685 B.n311 B.n210 163.367
R686 B.n311 B.n310 163.367
R687 B.n310 B.n309 163.367
R688 B.n309 B.n212 163.367
R689 B.n305 B.n212 163.367
R690 B.n305 B.n304 163.367
R691 B.n304 B.n303 163.367
R692 B.n303 B.n214 163.367
R693 B.n299 B.n214 163.367
R694 B.n299 B.n298 163.367
R695 B.n298 B.n297 163.367
R696 B.n297 B.n216 163.367
R697 B.n293 B.n216 163.367
R698 B.n293 B.n292 163.367
R699 B.n292 B.n291 163.367
R700 B.n291 B.n218 163.367
R701 B.n287 B.n218 163.367
R702 B.n287 B.n286 163.367
R703 B.n286 B.n285 163.367
R704 B.n285 B.n220 163.367
R705 B.n281 B.n220 163.367
R706 B.n281 B.n280 163.367
R707 B.n280 B.n279 163.367
R708 B.n279 B.n222 163.367
R709 B.n275 B.n222 163.367
R710 B.n275 B.n274 163.367
R711 B.n274 B.n273 163.367
R712 B.n273 B.n224 163.367
R713 B.n269 B.n224 163.367
R714 B.n269 B.n268 163.367
R715 B.n268 B.n267 163.367
R716 B.n267 B.n226 163.367
R717 B.n263 B.n226 163.367
R718 B.n263 B.n262 163.367
R719 B.n262 B.n261 163.367
R720 B.n261 B.n228 163.367
R721 B.n257 B.n228 163.367
R722 B.n257 B.n256 163.367
R723 B.n256 B.n255 163.367
R724 B.n255 B.n230 163.367
R725 B.n251 B.n230 163.367
R726 B.n251 B.n250 163.367
R727 B.n250 B.n249 163.367
R728 B.n249 B.n232 163.367
R729 B.n245 B.n232 163.367
R730 B.n245 B.n244 163.367
R731 B.n244 B.n243 163.367
R732 B.n243 B.n234 163.367
R733 B.n239 B.n234 163.367
R734 B.n239 B.n238 163.367
R735 B.n238 B.n237 163.367
R736 B.n237 B.n2 163.367
R737 B.n922 B.n2 163.367
R738 B.n922 B.n921 163.367
R739 B.n921 B.n920 163.367
R740 B.n920 B.n3 163.367
R741 B.n916 B.n3 163.367
R742 B.n916 B.n915 163.367
R743 B.n915 B.n914 163.367
R744 B.n914 B.n5 163.367
R745 B.n910 B.n5 163.367
R746 B.n910 B.n909 163.367
R747 B.n909 B.n908 163.367
R748 B.n908 B.n7 163.367
R749 B.n904 B.n7 163.367
R750 B.n904 B.n903 163.367
R751 B.n903 B.n902 163.367
R752 B.n902 B.n9 163.367
R753 B.n898 B.n9 163.367
R754 B.n898 B.n897 163.367
R755 B.n897 B.n896 163.367
R756 B.n896 B.n11 163.367
R757 B.n892 B.n11 163.367
R758 B.n892 B.n891 163.367
R759 B.n891 B.n890 163.367
R760 B.n890 B.n13 163.367
R761 B.n886 B.n13 163.367
R762 B.n886 B.n885 163.367
R763 B.n885 B.n884 163.367
R764 B.n884 B.n15 163.367
R765 B.n880 B.n15 163.367
R766 B.n880 B.n879 163.367
R767 B.n879 B.n878 163.367
R768 B.n878 B.n17 163.367
R769 B.n874 B.n17 163.367
R770 B.n874 B.n873 163.367
R771 B.n873 B.n872 163.367
R772 B.n872 B.n19 163.367
R773 B.n868 B.n19 163.367
R774 B.n868 B.n867 163.367
R775 B.n867 B.n866 163.367
R776 B.n866 B.n21 163.367
R777 B.n862 B.n21 163.367
R778 B.n862 B.n861 163.367
R779 B.n861 B.n860 163.367
R780 B.n860 B.n23 163.367
R781 B.n856 B.n23 163.367
R782 B.n856 B.n855 163.367
R783 B.n855 B.n854 163.367
R784 B.n854 B.n25 163.367
R785 B.n850 B.n25 163.367
R786 B.n850 B.n849 163.367
R787 B.n849 B.n848 163.367
R788 B.n848 B.n27 163.367
R789 B.n844 B.n27 163.367
R790 B.n844 B.n843 163.367
R791 B.n843 B.n842 163.367
R792 B.n842 B.n29 163.367
R793 B.n838 B.n29 163.367
R794 B.n838 B.n837 163.367
R795 B.n837 B.n836 163.367
R796 B.n836 B.n31 163.367
R797 B.n832 B.n31 163.367
R798 B.n327 B.n206 163.367
R799 B.n328 B.n327 163.367
R800 B.n329 B.n328 163.367
R801 B.n329 B.n204 163.367
R802 B.n333 B.n204 163.367
R803 B.n334 B.n333 163.367
R804 B.n335 B.n334 163.367
R805 B.n335 B.n202 163.367
R806 B.n339 B.n202 163.367
R807 B.n340 B.n339 163.367
R808 B.n341 B.n340 163.367
R809 B.n341 B.n200 163.367
R810 B.n345 B.n200 163.367
R811 B.n346 B.n345 163.367
R812 B.n347 B.n346 163.367
R813 B.n347 B.n198 163.367
R814 B.n351 B.n198 163.367
R815 B.n352 B.n351 163.367
R816 B.n353 B.n352 163.367
R817 B.n353 B.n196 163.367
R818 B.n357 B.n196 163.367
R819 B.n358 B.n357 163.367
R820 B.n359 B.n358 163.367
R821 B.n359 B.n194 163.367
R822 B.n363 B.n194 163.367
R823 B.n364 B.n363 163.367
R824 B.n365 B.n364 163.367
R825 B.n365 B.n192 163.367
R826 B.n369 B.n192 163.367
R827 B.n370 B.n369 163.367
R828 B.n371 B.n370 163.367
R829 B.n371 B.n190 163.367
R830 B.n375 B.n190 163.367
R831 B.n376 B.n375 163.367
R832 B.n377 B.n376 163.367
R833 B.n377 B.n188 163.367
R834 B.n381 B.n188 163.367
R835 B.n382 B.n381 163.367
R836 B.n383 B.n382 163.367
R837 B.n383 B.n186 163.367
R838 B.n387 B.n186 163.367
R839 B.n388 B.n387 163.367
R840 B.n389 B.n388 163.367
R841 B.n389 B.n184 163.367
R842 B.n393 B.n184 163.367
R843 B.n394 B.n393 163.367
R844 B.n395 B.n394 163.367
R845 B.n395 B.n180 163.367
R846 B.n400 B.n180 163.367
R847 B.n401 B.n400 163.367
R848 B.n402 B.n401 163.367
R849 B.n402 B.n178 163.367
R850 B.n406 B.n178 163.367
R851 B.n407 B.n406 163.367
R852 B.n408 B.n407 163.367
R853 B.n408 B.n176 163.367
R854 B.n415 B.n176 163.367
R855 B.n416 B.n415 163.367
R856 B.n417 B.n416 163.367
R857 B.n417 B.n174 163.367
R858 B.n421 B.n174 163.367
R859 B.n422 B.n421 163.367
R860 B.n423 B.n422 163.367
R861 B.n423 B.n172 163.367
R862 B.n427 B.n172 163.367
R863 B.n428 B.n427 163.367
R864 B.n429 B.n428 163.367
R865 B.n429 B.n170 163.367
R866 B.n433 B.n170 163.367
R867 B.n434 B.n433 163.367
R868 B.n435 B.n434 163.367
R869 B.n435 B.n168 163.367
R870 B.n439 B.n168 163.367
R871 B.n440 B.n439 163.367
R872 B.n441 B.n440 163.367
R873 B.n441 B.n166 163.367
R874 B.n445 B.n166 163.367
R875 B.n446 B.n445 163.367
R876 B.n447 B.n446 163.367
R877 B.n447 B.n164 163.367
R878 B.n451 B.n164 163.367
R879 B.n452 B.n451 163.367
R880 B.n453 B.n452 163.367
R881 B.n453 B.n162 163.367
R882 B.n457 B.n162 163.367
R883 B.n458 B.n457 163.367
R884 B.n459 B.n458 163.367
R885 B.n459 B.n160 163.367
R886 B.n463 B.n160 163.367
R887 B.n464 B.n463 163.367
R888 B.n465 B.n464 163.367
R889 B.n465 B.n158 163.367
R890 B.n469 B.n158 163.367
R891 B.n470 B.n469 163.367
R892 B.n471 B.n470 163.367
R893 B.n471 B.n156 163.367
R894 B.n475 B.n156 163.367
R895 B.n476 B.n475 163.367
R896 B.n477 B.n476 163.367
R897 B.n477 B.n154 163.367
R898 B.n481 B.n154 163.367
R899 B.n482 B.n481 163.367
R900 B.n483 B.n482 163.367
R901 B.n483 B.n152 163.367
R902 B.n487 B.n152 163.367
R903 B.n488 B.n487 163.367
R904 B.n489 B.n150 163.367
R905 B.n493 B.n150 163.367
R906 B.n494 B.n493 163.367
R907 B.n495 B.n494 163.367
R908 B.n495 B.n148 163.367
R909 B.n499 B.n148 163.367
R910 B.n500 B.n499 163.367
R911 B.n501 B.n500 163.367
R912 B.n501 B.n146 163.367
R913 B.n505 B.n146 163.367
R914 B.n506 B.n505 163.367
R915 B.n507 B.n506 163.367
R916 B.n507 B.n144 163.367
R917 B.n511 B.n144 163.367
R918 B.n512 B.n511 163.367
R919 B.n513 B.n512 163.367
R920 B.n513 B.n142 163.367
R921 B.n517 B.n142 163.367
R922 B.n518 B.n517 163.367
R923 B.n519 B.n518 163.367
R924 B.n519 B.n140 163.367
R925 B.n523 B.n140 163.367
R926 B.n524 B.n523 163.367
R927 B.n525 B.n524 163.367
R928 B.n525 B.n138 163.367
R929 B.n529 B.n138 163.367
R930 B.n530 B.n529 163.367
R931 B.n531 B.n530 163.367
R932 B.n531 B.n136 163.367
R933 B.n535 B.n136 163.367
R934 B.n536 B.n535 163.367
R935 B.n537 B.n536 163.367
R936 B.n537 B.n134 163.367
R937 B.n541 B.n134 163.367
R938 B.n542 B.n541 163.367
R939 B.n543 B.n542 163.367
R940 B.n543 B.n132 163.367
R941 B.n547 B.n132 163.367
R942 B.n548 B.n547 163.367
R943 B.n549 B.n548 163.367
R944 B.n549 B.n130 163.367
R945 B.n553 B.n130 163.367
R946 B.n554 B.n553 163.367
R947 B.n555 B.n554 163.367
R948 B.n555 B.n128 163.367
R949 B.n559 B.n128 163.367
R950 B.n560 B.n559 163.367
R951 B.n561 B.n560 163.367
R952 B.n561 B.n126 163.367
R953 B.n565 B.n126 163.367
R954 B.n566 B.n565 163.367
R955 B.n567 B.n566 163.367
R956 B.n567 B.n124 163.367
R957 B.n571 B.n124 163.367
R958 B.n572 B.n571 163.367
R959 B.n573 B.n572 163.367
R960 B.n573 B.n122 163.367
R961 B.n577 B.n122 163.367
R962 B.n578 B.n577 163.367
R963 B.n579 B.n578 163.367
R964 B.n579 B.n120 163.367
R965 B.n583 B.n120 163.367
R966 B.n584 B.n583 163.367
R967 B.n585 B.n584 163.367
R968 B.n585 B.n118 163.367
R969 B.n589 B.n118 163.367
R970 B.n590 B.n589 163.367
R971 B.n591 B.n590 163.367
R972 B.n591 B.n116 163.367
R973 B.n595 B.n116 163.367
R974 B.n596 B.n595 163.367
R975 B.n597 B.n596 163.367
R976 B.n597 B.n114 163.367
R977 B.n601 B.n114 163.367
R978 B.n602 B.n601 163.367
R979 B.n603 B.n602 163.367
R980 B.n603 B.n112 163.367
R981 B.n607 B.n112 163.367
R982 B.n608 B.n607 163.367
R983 B.n609 B.n608 163.367
R984 B.n609 B.n110 163.367
R985 B.n613 B.n110 163.367
R986 B.n614 B.n613 163.367
R987 B.n615 B.n614 163.367
R988 B.n615 B.n108 163.367
R989 B.n619 B.n108 163.367
R990 B.n620 B.n619 163.367
R991 B.n621 B.n620 163.367
R992 B.n621 B.n106 163.367
R993 B.n625 B.n106 163.367
R994 B.n626 B.n625 163.367
R995 B.n627 B.n626 163.367
R996 B.n627 B.n104 163.367
R997 B.n631 B.n104 163.367
R998 B.n632 B.n631 163.367
R999 B.n633 B.n632 163.367
R1000 B.n633 B.n102 163.367
R1001 B.n637 B.n102 163.367
R1002 B.n638 B.n637 163.367
R1003 B.n639 B.n638 163.367
R1004 B.n639 B.n100 163.367
R1005 B.n643 B.n100 163.367
R1006 B.n644 B.n643 163.367
R1007 B.n645 B.n644 163.367
R1008 B.n645 B.n98 163.367
R1009 B.n649 B.n98 163.367
R1010 B.n650 B.n649 163.367
R1011 B.n651 B.n650 163.367
R1012 B.n651 B.n96 163.367
R1013 B.n655 B.n96 163.367
R1014 B.n656 B.n655 163.367
R1015 B.n657 B.n656 163.367
R1016 B.n657 B.n94 163.367
R1017 B.n661 B.n94 163.367
R1018 B.n662 B.n661 163.367
R1019 B.n663 B.n662 163.367
R1020 B.n663 B.n92 163.367
R1021 B.n667 B.n92 163.367
R1022 B.n668 B.n667 163.367
R1023 B.n669 B.n668 163.367
R1024 B.n831 B.n830 163.367
R1025 B.n830 B.n33 163.367
R1026 B.n826 B.n33 163.367
R1027 B.n826 B.n825 163.367
R1028 B.n825 B.n824 163.367
R1029 B.n824 B.n35 163.367
R1030 B.n820 B.n35 163.367
R1031 B.n820 B.n819 163.367
R1032 B.n819 B.n818 163.367
R1033 B.n818 B.n37 163.367
R1034 B.n814 B.n37 163.367
R1035 B.n814 B.n813 163.367
R1036 B.n813 B.n812 163.367
R1037 B.n812 B.n39 163.367
R1038 B.n808 B.n39 163.367
R1039 B.n808 B.n807 163.367
R1040 B.n807 B.n806 163.367
R1041 B.n806 B.n41 163.367
R1042 B.n802 B.n41 163.367
R1043 B.n802 B.n801 163.367
R1044 B.n801 B.n800 163.367
R1045 B.n800 B.n43 163.367
R1046 B.n796 B.n43 163.367
R1047 B.n796 B.n795 163.367
R1048 B.n795 B.n794 163.367
R1049 B.n794 B.n45 163.367
R1050 B.n790 B.n45 163.367
R1051 B.n790 B.n789 163.367
R1052 B.n789 B.n788 163.367
R1053 B.n788 B.n47 163.367
R1054 B.n784 B.n47 163.367
R1055 B.n784 B.n783 163.367
R1056 B.n783 B.n782 163.367
R1057 B.n782 B.n49 163.367
R1058 B.n778 B.n49 163.367
R1059 B.n778 B.n777 163.367
R1060 B.n777 B.n776 163.367
R1061 B.n776 B.n51 163.367
R1062 B.n772 B.n51 163.367
R1063 B.n772 B.n771 163.367
R1064 B.n771 B.n770 163.367
R1065 B.n770 B.n53 163.367
R1066 B.n766 B.n53 163.367
R1067 B.n766 B.n765 163.367
R1068 B.n765 B.n764 163.367
R1069 B.n764 B.n55 163.367
R1070 B.n760 B.n55 163.367
R1071 B.n760 B.n759 163.367
R1072 B.n759 B.n758 163.367
R1073 B.n758 B.n57 163.367
R1074 B.n754 B.n57 163.367
R1075 B.n754 B.n753 163.367
R1076 B.n753 B.n752 163.367
R1077 B.n752 B.n62 163.367
R1078 B.n748 B.n62 163.367
R1079 B.n748 B.n747 163.367
R1080 B.n747 B.n746 163.367
R1081 B.n746 B.n64 163.367
R1082 B.n741 B.n64 163.367
R1083 B.n741 B.n740 163.367
R1084 B.n740 B.n739 163.367
R1085 B.n739 B.n68 163.367
R1086 B.n735 B.n68 163.367
R1087 B.n735 B.n734 163.367
R1088 B.n734 B.n733 163.367
R1089 B.n733 B.n70 163.367
R1090 B.n729 B.n70 163.367
R1091 B.n729 B.n728 163.367
R1092 B.n728 B.n727 163.367
R1093 B.n727 B.n72 163.367
R1094 B.n723 B.n72 163.367
R1095 B.n723 B.n722 163.367
R1096 B.n722 B.n721 163.367
R1097 B.n721 B.n74 163.367
R1098 B.n717 B.n74 163.367
R1099 B.n717 B.n716 163.367
R1100 B.n716 B.n715 163.367
R1101 B.n715 B.n76 163.367
R1102 B.n711 B.n76 163.367
R1103 B.n711 B.n710 163.367
R1104 B.n710 B.n709 163.367
R1105 B.n709 B.n78 163.367
R1106 B.n705 B.n78 163.367
R1107 B.n705 B.n704 163.367
R1108 B.n704 B.n703 163.367
R1109 B.n703 B.n80 163.367
R1110 B.n699 B.n80 163.367
R1111 B.n699 B.n698 163.367
R1112 B.n698 B.n697 163.367
R1113 B.n697 B.n82 163.367
R1114 B.n693 B.n82 163.367
R1115 B.n693 B.n692 163.367
R1116 B.n692 B.n691 163.367
R1117 B.n691 B.n84 163.367
R1118 B.n687 B.n84 163.367
R1119 B.n687 B.n686 163.367
R1120 B.n686 B.n685 163.367
R1121 B.n685 B.n86 163.367
R1122 B.n681 B.n86 163.367
R1123 B.n681 B.n680 163.367
R1124 B.n680 B.n679 163.367
R1125 B.n679 B.n88 163.367
R1126 B.n675 B.n88 163.367
R1127 B.n675 B.n674 163.367
R1128 B.n674 B.n673 163.367
R1129 B.n673 B.n90 163.367
R1130 B.n412 B.t1 107.825
R1131 B.n66 B.t5 107.825
R1132 B.n182 B.t10 107.806
R1133 B.n59 B.t8 107.806
R1134 B.n413 B.n412 59.5399
R1135 B.n398 B.n182 59.5399
R1136 B.n60 B.n59 59.5399
R1137 B.n744 B.n66 59.5399
R1138 B.n412 B.n411 57.0187
R1139 B.n182 B.n181 57.0187
R1140 B.n59 B.n58 57.0187
R1141 B.n66 B.n65 57.0187
R1142 B.n671 B.n670 30.1273
R1143 B.n833 B.n32 30.1273
R1144 B.n490 B.n151 30.1273
R1145 B.n325 B.n324 30.1273
R1146 B B.n923 18.0485
R1147 B.n829 B.n32 10.6151
R1148 B.n829 B.n828 10.6151
R1149 B.n828 B.n827 10.6151
R1150 B.n827 B.n34 10.6151
R1151 B.n823 B.n34 10.6151
R1152 B.n823 B.n822 10.6151
R1153 B.n822 B.n821 10.6151
R1154 B.n821 B.n36 10.6151
R1155 B.n817 B.n36 10.6151
R1156 B.n817 B.n816 10.6151
R1157 B.n816 B.n815 10.6151
R1158 B.n815 B.n38 10.6151
R1159 B.n811 B.n38 10.6151
R1160 B.n811 B.n810 10.6151
R1161 B.n810 B.n809 10.6151
R1162 B.n809 B.n40 10.6151
R1163 B.n805 B.n40 10.6151
R1164 B.n805 B.n804 10.6151
R1165 B.n804 B.n803 10.6151
R1166 B.n803 B.n42 10.6151
R1167 B.n799 B.n42 10.6151
R1168 B.n799 B.n798 10.6151
R1169 B.n798 B.n797 10.6151
R1170 B.n797 B.n44 10.6151
R1171 B.n793 B.n44 10.6151
R1172 B.n793 B.n792 10.6151
R1173 B.n792 B.n791 10.6151
R1174 B.n791 B.n46 10.6151
R1175 B.n787 B.n46 10.6151
R1176 B.n787 B.n786 10.6151
R1177 B.n786 B.n785 10.6151
R1178 B.n785 B.n48 10.6151
R1179 B.n781 B.n48 10.6151
R1180 B.n781 B.n780 10.6151
R1181 B.n780 B.n779 10.6151
R1182 B.n779 B.n50 10.6151
R1183 B.n775 B.n50 10.6151
R1184 B.n775 B.n774 10.6151
R1185 B.n774 B.n773 10.6151
R1186 B.n773 B.n52 10.6151
R1187 B.n769 B.n52 10.6151
R1188 B.n769 B.n768 10.6151
R1189 B.n768 B.n767 10.6151
R1190 B.n767 B.n54 10.6151
R1191 B.n763 B.n54 10.6151
R1192 B.n763 B.n762 10.6151
R1193 B.n762 B.n761 10.6151
R1194 B.n761 B.n56 10.6151
R1195 B.n757 B.n756 10.6151
R1196 B.n756 B.n755 10.6151
R1197 B.n755 B.n61 10.6151
R1198 B.n751 B.n61 10.6151
R1199 B.n751 B.n750 10.6151
R1200 B.n750 B.n749 10.6151
R1201 B.n749 B.n63 10.6151
R1202 B.n745 B.n63 10.6151
R1203 B.n743 B.n742 10.6151
R1204 B.n742 B.n67 10.6151
R1205 B.n738 B.n67 10.6151
R1206 B.n738 B.n737 10.6151
R1207 B.n737 B.n736 10.6151
R1208 B.n736 B.n69 10.6151
R1209 B.n732 B.n69 10.6151
R1210 B.n732 B.n731 10.6151
R1211 B.n731 B.n730 10.6151
R1212 B.n730 B.n71 10.6151
R1213 B.n726 B.n71 10.6151
R1214 B.n726 B.n725 10.6151
R1215 B.n725 B.n724 10.6151
R1216 B.n724 B.n73 10.6151
R1217 B.n720 B.n73 10.6151
R1218 B.n720 B.n719 10.6151
R1219 B.n719 B.n718 10.6151
R1220 B.n718 B.n75 10.6151
R1221 B.n714 B.n75 10.6151
R1222 B.n714 B.n713 10.6151
R1223 B.n713 B.n712 10.6151
R1224 B.n712 B.n77 10.6151
R1225 B.n708 B.n77 10.6151
R1226 B.n708 B.n707 10.6151
R1227 B.n707 B.n706 10.6151
R1228 B.n706 B.n79 10.6151
R1229 B.n702 B.n79 10.6151
R1230 B.n702 B.n701 10.6151
R1231 B.n701 B.n700 10.6151
R1232 B.n700 B.n81 10.6151
R1233 B.n696 B.n81 10.6151
R1234 B.n696 B.n695 10.6151
R1235 B.n695 B.n694 10.6151
R1236 B.n694 B.n83 10.6151
R1237 B.n690 B.n83 10.6151
R1238 B.n690 B.n689 10.6151
R1239 B.n689 B.n688 10.6151
R1240 B.n688 B.n85 10.6151
R1241 B.n684 B.n85 10.6151
R1242 B.n684 B.n683 10.6151
R1243 B.n683 B.n682 10.6151
R1244 B.n682 B.n87 10.6151
R1245 B.n678 B.n87 10.6151
R1246 B.n678 B.n677 10.6151
R1247 B.n677 B.n676 10.6151
R1248 B.n676 B.n89 10.6151
R1249 B.n672 B.n89 10.6151
R1250 B.n672 B.n671 10.6151
R1251 B.n491 B.n490 10.6151
R1252 B.n492 B.n491 10.6151
R1253 B.n492 B.n149 10.6151
R1254 B.n496 B.n149 10.6151
R1255 B.n497 B.n496 10.6151
R1256 B.n498 B.n497 10.6151
R1257 B.n498 B.n147 10.6151
R1258 B.n502 B.n147 10.6151
R1259 B.n503 B.n502 10.6151
R1260 B.n504 B.n503 10.6151
R1261 B.n504 B.n145 10.6151
R1262 B.n508 B.n145 10.6151
R1263 B.n509 B.n508 10.6151
R1264 B.n510 B.n509 10.6151
R1265 B.n510 B.n143 10.6151
R1266 B.n514 B.n143 10.6151
R1267 B.n515 B.n514 10.6151
R1268 B.n516 B.n515 10.6151
R1269 B.n516 B.n141 10.6151
R1270 B.n520 B.n141 10.6151
R1271 B.n521 B.n520 10.6151
R1272 B.n522 B.n521 10.6151
R1273 B.n522 B.n139 10.6151
R1274 B.n526 B.n139 10.6151
R1275 B.n527 B.n526 10.6151
R1276 B.n528 B.n527 10.6151
R1277 B.n528 B.n137 10.6151
R1278 B.n532 B.n137 10.6151
R1279 B.n533 B.n532 10.6151
R1280 B.n534 B.n533 10.6151
R1281 B.n534 B.n135 10.6151
R1282 B.n538 B.n135 10.6151
R1283 B.n539 B.n538 10.6151
R1284 B.n540 B.n539 10.6151
R1285 B.n540 B.n133 10.6151
R1286 B.n544 B.n133 10.6151
R1287 B.n545 B.n544 10.6151
R1288 B.n546 B.n545 10.6151
R1289 B.n546 B.n131 10.6151
R1290 B.n550 B.n131 10.6151
R1291 B.n551 B.n550 10.6151
R1292 B.n552 B.n551 10.6151
R1293 B.n552 B.n129 10.6151
R1294 B.n556 B.n129 10.6151
R1295 B.n557 B.n556 10.6151
R1296 B.n558 B.n557 10.6151
R1297 B.n558 B.n127 10.6151
R1298 B.n562 B.n127 10.6151
R1299 B.n563 B.n562 10.6151
R1300 B.n564 B.n563 10.6151
R1301 B.n564 B.n125 10.6151
R1302 B.n568 B.n125 10.6151
R1303 B.n569 B.n568 10.6151
R1304 B.n570 B.n569 10.6151
R1305 B.n570 B.n123 10.6151
R1306 B.n574 B.n123 10.6151
R1307 B.n575 B.n574 10.6151
R1308 B.n576 B.n575 10.6151
R1309 B.n576 B.n121 10.6151
R1310 B.n580 B.n121 10.6151
R1311 B.n581 B.n580 10.6151
R1312 B.n582 B.n581 10.6151
R1313 B.n582 B.n119 10.6151
R1314 B.n586 B.n119 10.6151
R1315 B.n587 B.n586 10.6151
R1316 B.n588 B.n587 10.6151
R1317 B.n588 B.n117 10.6151
R1318 B.n592 B.n117 10.6151
R1319 B.n593 B.n592 10.6151
R1320 B.n594 B.n593 10.6151
R1321 B.n594 B.n115 10.6151
R1322 B.n598 B.n115 10.6151
R1323 B.n599 B.n598 10.6151
R1324 B.n600 B.n599 10.6151
R1325 B.n600 B.n113 10.6151
R1326 B.n604 B.n113 10.6151
R1327 B.n605 B.n604 10.6151
R1328 B.n606 B.n605 10.6151
R1329 B.n606 B.n111 10.6151
R1330 B.n610 B.n111 10.6151
R1331 B.n611 B.n610 10.6151
R1332 B.n612 B.n611 10.6151
R1333 B.n612 B.n109 10.6151
R1334 B.n616 B.n109 10.6151
R1335 B.n617 B.n616 10.6151
R1336 B.n618 B.n617 10.6151
R1337 B.n618 B.n107 10.6151
R1338 B.n622 B.n107 10.6151
R1339 B.n623 B.n622 10.6151
R1340 B.n624 B.n623 10.6151
R1341 B.n624 B.n105 10.6151
R1342 B.n628 B.n105 10.6151
R1343 B.n629 B.n628 10.6151
R1344 B.n630 B.n629 10.6151
R1345 B.n630 B.n103 10.6151
R1346 B.n634 B.n103 10.6151
R1347 B.n635 B.n634 10.6151
R1348 B.n636 B.n635 10.6151
R1349 B.n636 B.n101 10.6151
R1350 B.n640 B.n101 10.6151
R1351 B.n641 B.n640 10.6151
R1352 B.n642 B.n641 10.6151
R1353 B.n642 B.n99 10.6151
R1354 B.n646 B.n99 10.6151
R1355 B.n647 B.n646 10.6151
R1356 B.n648 B.n647 10.6151
R1357 B.n648 B.n97 10.6151
R1358 B.n652 B.n97 10.6151
R1359 B.n653 B.n652 10.6151
R1360 B.n654 B.n653 10.6151
R1361 B.n654 B.n95 10.6151
R1362 B.n658 B.n95 10.6151
R1363 B.n659 B.n658 10.6151
R1364 B.n660 B.n659 10.6151
R1365 B.n660 B.n93 10.6151
R1366 B.n664 B.n93 10.6151
R1367 B.n665 B.n664 10.6151
R1368 B.n666 B.n665 10.6151
R1369 B.n666 B.n91 10.6151
R1370 B.n670 B.n91 10.6151
R1371 B.n326 B.n325 10.6151
R1372 B.n326 B.n205 10.6151
R1373 B.n330 B.n205 10.6151
R1374 B.n331 B.n330 10.6151
R1375 B.n332 B.n331 10.6151
R1376 B.n332 B.n203 10.6151
R1377 B.n336 B.n203 10.6151
R1378 B.n337 B.n336 10.6151
R1379 B.n338 B.n337 10.6151
R1380 B.n338 B.n201 10.6151
R1381 B.n342 B.n201 10.6151
R1382 B.n343 B.n342 10.6151
R1383 B.n344 B.n343 10.6151
R1384 B.n344 B.n199 10.6151
R1385 B.n348 B.n199 10.6151
R1386 B.n349 B.n348 10.6151
R1387 B.n350 B.n349 10.6151
R1388 B.n350 B.n197 10.6151
R1389 B.n354 B.n197 10.6151
R1390 B.n355 B.n354 10.6151
R1391 B.n356 B.n355 10.6151
R1392 B.n356 B.n195 10.6151
R1393 B.n360 B.n195 10.6151
R1394 B.n361 B.n360 10.6151
R1395 B.n362 B.n361 10.6151
R1396 B.n362 B.n193 10.6151
R1397 B.n366 B.n193 10.6151
R1398 B.n367 B.n366 10.6151
R1399 B.n368 B.n367 10.6151
R1400 B.n368 B.n191 10.6151
R1401 B.n372 B.n191 10.6151
R1402 B.n373 B.n372 10.6151
R1403 B.n374 B.n373 10.6151
R1404 B.n374 B.n189 10.6151
R1405 B.n378 B.n189 10.6151
R1406 B.n379 B.n378 10.6151
R1407 B.n380 B.n379 10.6151
R1408 B.n380 B.n187 10.6151
R1409 B.n384 B.n187 10.6151
R1410 B.n385 B.n384 10.6151
R1411 B.n386 B.n385 10.6151
R1412 B.n386 B.n185 10.6151
R1413 B.n390 B.n185 10.6151
R1414 B.n391 B.n390 10.6151
R1415 B.n392 B.n391 10.6151
R1416 B.n392 B.n183 10.6151
R1417 B.n396 B.n183 10.6151
R1418 B.n397 B.n396 10.6151
R1419 B.n399 B.n179 10.6151
R1420 B.n403 B.n179 10.6151
R1421 B.n404 B.n403 10.6151
R1422 B.n405 B.n404 10.6151
R1423 B.n405 B.n177 10.6151
R1424 B.n409 B.n177 10.6151
R1425 B.n410 B.n409 10.6151
R1426 B.n414 B.n410 10.6151
R1427 B.n418 B.n175 10.6151
R1428 B.n419 B.n418 10.6151
R1429 B.n420 B.n419 10.6151
R1430 B.n420 B.n173 10.6151
R1431 B.n424 B.n173 10.6151
R1432 B.n425 B.n424 10.6151
R1433 B.n426 B.n425 10.6151
R1434 B.n426 B.n171 10.6151
R1435 B.n430 B.n171 10.6151
R1436 B.n431 B.n430 10.6151
R1437 B.n432 B.n431 10.6151
R1438 B.n432 B.n169 10.6151
R1439 B.n436 B.n169 10.6151
R1440 B.n437 B.n436 10.6151
R1441 B.n438 B.n437 10.6151
R1442 B.n438 B.n167 10.6151
R1443 B.n442 B.n167 10.6151
R1444 B.n443 B.n442 10.6151
R1445 B.n444 B.n443 10.6151
R1446 B.n444 B.n165 10.6151
R1447 B.n448 B.n165 10.6151
R1448 B.n449 B.n448 10.6151
R1449 B.n450 B.n449 10.6151
R1450 B.n450 B.n163 10.6151
R1451 B.n454 B.n163 10.6151
R1452 B.n455 B.n454 10.6151
R1453 B.n456 B.n455 10.6151
R1454 B.n456 B.n161 10.6151
R1455 B.n460 B.n161 10.6151
R1456 B.n461 B.n460 10.6151
R1457 B.n462 B.n461 10.6151
R1458 B.n462 B.n159 10.6151
R1459 B.n466 B.n159 10.6151
R1460 B.n467 B.n466 10.6151
R1461 B.n468 B.n467 10.6151
R1462 B.n468 B.n157 10.6151
R1463 B.n472 B.n157 10.6151
R1464 B.n473 B.n472 10.6151
R1465 B.n474 B.n473 10.6151
R1466 B.n474 B.n155 10.6151
R1467 B.n478 B.n155 10.6151
R1468 B.n479 B.n478 10.6151
R1469 B.n480 B.n479 10.6151
R1470 B.n480 B.n153 10.6151
R1471 B.n484 B.n153 10.6151
R1472 B.n485 B.n484 10.6151
R1473 B.n486 B.n485 10.6151
R1474 B.n486 B.n151 10.6151
R1475 B.n324 B.n207 10.6151
R1476 B.n320 B.n207 10.6151
R1477 B.n320 B.n319 10.6151
R1478 B.n319 B.n318 10.6151
R1479 B.n318 B.n209 10.6151
R1480 B.n314 B.n209 10.6151
R1481 B.n314 B.n313 10.6151
R1482 B.n313 B.n312 10.6151
R1483 B.n312 B.n211 10.6151
R1484 B.n308 B.n211 10.6151
R1485 B.n308 B.n307 10.6151
R1486 B.n307 B.n306 10.6151
R1487 B.n306 B.n213 10.6151
R1488 B.n302 B.n213 10.6151
R1489 B.n302 B.n301 10.6151
R1490 B.n301 B.n300 10.6151
R1491 B.n300 B.n215 10.6151
R1492 B.n296 B.n215 10.6151
R1493 B.n296 B.n295 10.6151
R1494 B.n295 B.n294 10.6151
R1495 B.n294 B.n217 10.6151
R1496 B.n290 B.n217 10.6151
R1497 B.n290 B.n289 10.6151
R1498 B.n289 B.n288 10.6151
R1499 B.n288 B.n219 10.6151
R1500 B.n284 B.n219 10.6151
R1501 B.n284 B.n283 10.6151
R1502 B.n283 B.n282 10.6151
R1503 B.n282 B.n221 10.6151
R1504 B.n278 B.n221 10.6151
R1505 B.n278 B.n277 10.6151
R1506 B.n277 B.n276 10.6151
R1507 B.n276 B.n223 10.6151
R1508 B.n272 B.n223 10.6151
R1509 B.n272 B.n271 10.6151
R1510 B.n271 B.n270 10.6151
R1511 B.n270 B.n225 10.6151
R1512 B.n266 B.n225 10.6151
R1513 B.n266 B.n265 10.6151
R1514 B.n265 B.n264 10.6151
R1515 B.n264 B.n227 10.6151
R1516 B.n260 B.n227 10.6151
R1517 B.n260 B.n259 10.6151
R1518 B.n259 B.n258 10.6151
R1519 B.n258 B.n229 10.6151
R1520 B.n254 B.n229 10.6151
R1521 B.n254 B.n253 10.6151
R1522 B.n253 B.n252 10.6151
R1523 B.n252 B.n231 10.6151
R1524 B.n248 B.n231 10.6151
R1525 B.n248 B.n247 10.6151
R1526 B.n247 B.n246 10.6151
R1527 B.n246 B.n233 10.6151
R1528 B.n242 B.n233 10.6151
R1529 B.n242 B.n241 10.6151
R1530 B.n241 B.n240 10.6151
R1531 B.n240 B.n235 10.6151
R1532 B.n236 B.n235 10.6151
R1533 B.n236 B.n0 10.6151
R1534 B.n919 B.n1 10.6151
R1535 B.n919 B.n918 10.6151
R1536 B.n918 B.n917 10.6151
R1537 B.n917 B.n4 10.6151
R1538 B.n913 B.n4 10.6151
R1539 B.n913 B.n912 10.6151
R1540 B.n912 B.n911 10.6151
R1541 B.n911 B.n6 10.6151
R1542 B.n907 B.n6 10.6151
R1543 B.n907 B.n906 10.6151
R1544 B.n906 B.n905 10.6151
R1545 B.n905 B.n8 10.6151
R1546 B.n901 B.n8 10.6151
R1547 B.n901 B.n900 10.6151
R1548 B.n900 B.n899 10.6151
R1549 B.n899 B.n10 10.6151
R1550 B.n895 B.n10 10.6151
R1551 B.n895 B.n894 10.6151
R1552 B.n894 B.n893 10.6151
R1553 B.n893 B.n12 10.6151
R1554 B.n889 B.n12 10.6151
R1555 B.n889 B.n888 10.6151
R1556 B.n888 B.n887 10.6151
R1557 B.n887 B.n14 10.6151
R1558 B.n883 B.n14 10.6151
R1559 B.n883 B.n882 10.6151
R1560 B.n882 B.n881 10.6151
R1561 B.n881 B.n16 10.6151
R1562 B.n877 B.n16 10.6151
R1563 B.n877 B.n876 10.6151
R1564 B.n876 B.n875 10.6151
R1565 B.n875 B.n18 10.6151
R1566 B.n871 B.n18 10.6151
R1567 B.n871 B.n870 10.6151
R1568 B.n870 B.n869 10.6151
R1569 B.n869 B.n20 10.6151
R1570 B.n865 B.n20 10.6151
R1571 B.n865 B.n864 10.6151
R1572 B.n864 B.n863 10.6151
R1573 B.n863 B.n22 10.6151
R1574 B.n859 B.n22 10.6151
R1575 B.n859 B.n858 10.6151
R1576 B.n858 B.n857 10.6151
R1577 B.n857 B.n24 10.6151
R1578 B.n853 B.n24 10.6151
R1579 B.n853 B.n852 10.6151
R1580 B.n852 B.n851 10.6151
R1581 B.n851 B.n26 10.6151
R1582 B.n847 B.n26 10.6151
R1583 B.n847 B.n846 10.6151
R1584 B.n846 B.n845 10.6151
R1585 B.n845 B.n28 10.6151
R1586 B.n841 B.n28 10.6151
R1587 B.n841 B.n840 10.6151
R1588 B.n840 B.n839 10.6151
R1589 B.n839 B.n30 10.6151
R1590 B.n835 B.n30 10.6151
R1591 B.n835 B.n834 10.6151
R1592 B.n834 B.n833 10.6151
R1593 B.n757 B.n60 6.5566
R1594 B.n745 B.n744 6.5566
R1595 B.n399 B.n398 6.5566
R1596 B.n414 B.n413 6.5566
R1597 B.n60 B.n56 4.05904
R1598 B.n744 B.n743 4.05904
R1599 B.n398 B.n397 4.05904
R1600 B.n413 B.n175 4.05904
R1601 B.n923 B.n0 2.81026
R1602 B.n923 B.n1 2.81026
R1603 VN.n11 VN.t1 164.99
R1604 VN.n53 VN.t3 164.99
R1605 VN.n81 VN.n42 161.3
R1606 VN.n80 VN.n79 161.3
R1607 VN.n78 VN.n43 161.3
R1608 VN.n77 VN.n76 161.3
R1609 VN.n75 VN.n44 161.3
R1610 VN.n74 VN.n73 161.3
R1611 VN.n72 VN.n71 161.3
R1612 VN.n70 VN.n46 161.3
R1613 VN.n69 VN.n68 161.3
R1614 VN.n67 VN.n47 161.3
R1615 VN.n66 VN.n65 161.3
R1616 VN.n64 VN.n48 161.3
R1617 VN.n62 VN.n61 161.3
R1618 VN.n60 VN.n49 161.3
R1619 VN.n59 VN.n58 161.3
R1620 VN.n57 VN.n50 161.3
R1621 VN.n56 VN.n55 161.3
R1622 VN.n54 VN.n51 161.3
R1623 VN.n39 VN.n0 161.3
R1624 VN.n38 VN.n37 161.3
R1625 VN.n36 VN.n1 161.3
R1626 VN.n35 VN.n34 161.3
R1627 VN.n33 VN.n2 161.3
R1628 VN.n32 VN.n31 161.3
R1629 VN.n30 VN.n29 161.3
R1630 VN.n28 VN.n4 161.3
R1631 VN.n27 VN.n26 161.3
R1632 VN.n25 VN.n5 161.3
R1633 VN.n24 VN.n23 161.3
R1634 VN.n22 VN.n6 161.3
R1635 VN.n20 VN.n19 161.3
R1636 VN.n18 VN.n7 161.3
R1637 VN.n17 VN.n16 161.3
R1638 VN.n15 VN.n8 161.3
R1639 VN.n14 VN.n13 161.3
R1640 VN.n12 VN.n9 161.3
R1641 VN.n10 VN.t5 132.411
R1642 VN.n21 VN.t9 132.411
R1643 VN.n3 VN.t0 132.411
R1644 VN.n40 VN.t2 132.411
R1645 VN.n52 VN.t6 132.411
R1646 VN.n63 VN.t7 132.411
R1647 VN.n45 VN.t8 132.411
R1648 VN.n82 VN.t4 132.411
R1649 VN.n41 VN.n40 104.514
R1650 VN.n83 VN.n82 104.514
R1651 VN.n11 VN.n10 63.1649
R1652 VN.n53 VN.n52 63.1649
R1653 VN.n16 VN.n15 56.5617
R1654 VN.n27 VN.n5 56.5617
R1655 VN.n58 VN.n57 56.5617
R1656 VN.n69 VN.n47 56.5617
R1657 VN.n34 VN.n1 56.0773
R1658 VN.n76 VN.n43 56.0773
R1659 VN VN.n83 55.1876
R1660 VN.n34 VN.n33 25.0767
R1661 VN.n76 VN.n75 25.0767
R1662 VN.n14 VN.n9 24.5923
R1663 VN.n15 VN.n14 24.5923
R1664 VN.n16 VN.n7 24.5923
R1665 VN.n20 VN.n7 24.5923
R1666 VN.n23 VN.n22 24.5923
R1667 VN.n23 VN.n5 24.5923
R1668 VN.n28 VN.n27 24.5923
R1669 VN.n29 VN.n28 24.5923
R1670 VN.n33 VN.n32 24.5923
R1671 VN.n38 VN.n1 24.5923
R1672 VN.n39 VN.n38 24.5923
R1673 VN.n57 VN.n56 24.5923
R1674 VN.n56 VN.n51 24.5923
R1675 VN.n65 VN.n47 24.5923
R1676 VN.n65 VN.n64 24.5923
R1677 VN.n62 VN.n49 24.5923
R1678 VN.n58 VN.n49 24.5923
R1679 VN.n75 VN.n74 24.5923
R1680 VN.n71 VN.n70 24.5923
R1681 VN.n70 VN.n69 24.5923
R1682 VN.n81 VN.n80 24.5923
R1683 VN.n80 VN.n43 24.5923
R1684 VN.n32 VN.n3 15.2474
R1685 VN.n74 VN.n45 15.2474
R1686 VN.n21 VN.n20 12.2964
R1687 VN.n22 VN.n21 12.2964
R1688 VN.n64 VN.n63 12.2964
R1689 VN.n63 VN.n62 12.2964
R1690 VN.n10 VN.n9 9.3454
R1691 VN.n29 VN.n3 9.3454
R1692 VN.n52 VN.n51 9.3454
R1693 VN.n71 VN.n45 9.3454
R1694 VN.n54 VN.n53 7.05922
R1695 VN.n12 VN.n11 7.05922
R1696 VN.n40 VN.n39 6.39438
R1697 VN.n82 VN.n81 6.39438
R1698 VN.n83 VN.n42 0.278335
R1699 VN.n41 VN.n0 0.278335
R1700 VN.n79 VN.n42 0.189894
R1701 VN.n79 VN.n78 0.189894
R1702 VN.n78 VN.n77 0.189894
R1703 VN.n77 VN.n44 0.189894
R1704 VN.n73 VN.n44 0.189894
R1705 VN.n73 VN.n72 0.189894
R1706 VN.n72 VN.n46 0.189894
R1707 VN.n68 VN.n46 0.189894
R1708 VN.n68 VN.n67 0.189894
R1709 VN.n67 VN.n66 0.189894
R1710 VN.n66 VN.n48 0.189894
R1711 VN.n61 VN.n48 0.189894
R1712 VN.n61 VN.n60 0.189894
R1713 VN.n60 VN.n59 0.189894
R1714 VN.n59 VN.n50 0.189894
R1715 VN.n55 VN.n50 0.189894
R1716 VN.n55 VN.n54 0.189894
R1717 VN.n13 VN.n12 0.189894
R1718 VN.n13 VN.n8 0.189894
R1719 VN.n17 VN.n8 0.189894
R1720 VN.n18 VN.n17 0.189894
R1721 VN.n19 VN.n18 0.189894
R1722 VN.n19 VN.n6 0.189894
R1723 VN.n24 VN.n6 0.189894
R1724 VN.n25 VN.n24 0.189894
R1725 VN.n26 VN.n25 0.189894
R1726 VN.n26 VN.n4 0.189894
R1727 VN.n30 VN.n4 0.189894
R1728 VN.n31 VN.n30 0.189894
R1729 VN.n31 VN.n2 0.189894
R1730 VN.n35 VN.n2 0.189894
R1731 VN.n36 VN.n35 0.189894
R1732 VN.n37 VN.n36 0.189894
R1733 VN.n37 VN.n0 0.189894
R1734 VN VN.n41 0.153485
R1735 VDD2.n1 VDD2.t8 77.0073
R1736 VDD2.n4 VDD2.t5 74.4729
R1737 VDD2.n3 VDD2.n2 74.0515
R1738 VDD2 VDD2.n7 74.0487
R1739 VDD2.n6 VDD2.n5 72.2062
R1740 VDD2.n1 VDD2.n0 72.206
R1741 VDD2.n4 VDD2.n3 48.1162
R1742 VDD2.n6 VDD2.n4 2.53498
R1743 VDD2.n7 VDD2.t3 2.26724
R1744 VDD2.n7 VDD2.t6 2.26724
R1745 VDD2.n5 VDD2.t1 2.26724
R1746 VDD2.n5 VDD2.t2 2.26724
R1747 VDD2.n2 VDD2.t9 2.26724
R1748 VDD2.n2 VDD2.t7 2.26724
R1749 VDD2.n0 VDD2.t4 2.26724
R1750 VDD2.n0 VDD2.t0 2.26724
R1751 VDD2 VDD2.n6 0.69231
R1752 VDD2.n3 VDD2.n1 0.578775
C0 w_n4498_n3836# VN 9.65243f
C1 VTAIL B 4.25988f
C2 VDD2 VP 0.585515f
C3 VDD1 VDD2 2.18217f
C4 VDD2 w_n4498_n3836# 3.10184f
C5 VDD1 VP 13.0811f
C6 w_n4498_n3836# VP 10.2381f
C7 VDD1 w_n4498_n3836# 2.95778f
C8 VTAIL VN 13.1946f
C9 B VN 1.31715f
C10 VDD2 VTAIL 11.5226f
C11 VDD2 B 2.78743f
C12 VTAIL VP 13.2089f
C13 B VP 2.30201f
C14 VDD1 VTAIL 11.4721f
C15 VDD1 B 2.66912f
C16 VTAIL w_n4498_n3836# 3.54358f
C17 B w_n4498_n3836# 11.22f
C18 VDD2 VN 12.6537f
C19 VP VN 8.84078f
C20 VDD1 VN 0.153857f
C21 VDD2 VSUBS 2.22168f
C22 VDD1 VSUBS 2.026722f
C23 VTAIL VSUBS 1.377824f
C24 VN VSUBS 7.770279f
C25 VP VSUBS 4.332897f
C26 B VSUBS 5.57828f
C27 w_n4498_n3836# VSUBS 0.211748p
C28 VDD2.t8 VSUBS 3.51753f
C29 VDD2.t4 VSUBS 0.331998f
C30 VDD2.t0 VSUBS 0.331998f
C31 VDD2.n0 VSUBS 2.68147f
C32 VDD2.n1 VSUBS 1.71966f
C33 VDD2.t9 VSUBS 0.331998f
C34 VDD2.t7 VSUBS 0.331998f
C35 VDD2.n2 VSUBS 2.70584f
C36 VDD2.n3 VSUBS 3.88717f
C37 VDD2.t5 VSUBS 3.48786f
C38 VDD2.n4 VSUBS 4.20851f
C39 VDD2.t1 VSUBS 0.331998f
C40 VDD2.t2 VSUBS 0.331998f
C41 VDD2.n5 VSUBS 2.68147f
C42 VDD2.n6 VSUBS 0.856662f
C43 VDD2.t3 VSUBS 0.331998f
C44 VDD2.t6 VSUBS 0.331998f
C45 VDD2.n7 VSUBS 2.70578f
C46 VN.n0 VSUBS 0.035369f
C47 VN.t2 VSUBS 2.74867f
C48 VN.n1 VSUBS 0.045615f
C49 VN.n2 VSUBS 0.026829f
C50 VN.t0 VSUBS 2.74867f
C51 VN.n3 VSUBS 0.96259f
C52 VN.n4 VSUBS 0.026829f
C53 VN.n5 VSUBS 0.036773f
C54 VN.n6 VSUBS 0.026829f
C55 VN.t9 VSUBS 2.74867f
C56 VN.n7 VSUBS 0.049752f
C57 VN.n8 VSUBS 0.026829f
C58 VN.n9 VSUBS 0.034524f
C59 VN.t1 VSUBS 2.97113f
C60 VN.t5 VSUBS 2.74867f
C61 VN.n10 VSUBS 1.03677f
C62 VN.n11 VSUBS 1.01496f
C63 VN.n12 VSUBS 0.259375f
C64 VN.n13 VSUBS 0.026829f
C65 VN.n14 VSUBS 0.049752f
C66 VN.n15 VSUBS 0.041227f
C67 VN.n16 VSUBS 0.036773f
C68 VN.n17 VSUBS 0.026829f
C69 VN.n18 VSUBS 0.026829f
C70 VN.n19 VSUBS 0.026829f
C71 VN.n20 VSUBS 0.037471f
C72 VN.n21 VSUBS 0.96259f
C73 VN.n22 VSUBS 0.037471f
C74 VN.n23 VSUBS 0.049752f
C75 VN.n24 VSUBS 0.026829f
C76 VN.n25 VSUBS 0.026829f
C77 VN.n26 VSUBS 0.026829f
C78 VN.n27 VSUBS 0.041227f
C79 VN.n28 VSUBS 0.049752f
C80 VN.n29 VSUBS 0.034524f
C81 VN.n30 VSUBS 0.026829f
C82 VN.n31 VSUBS 0.026829f
C83 VN.n32 VSUBS 0.040419f
C84 VN.n33 VSUBS 0.050217f
C85 VN.n34 VSUBS 0.031921f
C86 VN.n35 VSUBS 0.026829f
C87 VN.n36 VSUBS 0.026829f
C88 VN.n37 VSUBS 0.026829f
C89 VN.n38 VSUBS 0.049752f
C90 VN.n39 VSUBS 0.031577f
C91 VN.n40 VSUBS 1.04708f
C92 VN.n41 VSUBS 0.046056f
C93 VN.n42 VSUBS 0.035369f
C94 VN.t4 VSUBS 2.74867f
C95 VN.n43 VSUBS 0.045615f
C96 VN.n44 VSUBS 0.026829f
C97 VN.t8 VSUBS 2.74867f
C98 VN.n45 VSUBS 0.96259f
C99 VN.n46 VSUBS 0.026829f
C100 VN.n47 VSUBS 0.036773f
C101 VN.n48 VSUBS 0.026829f
C102 VN.t7 VSUBS 2.74867f
C103 VN.n49 VSUBS 0.049752f
C104 VN.n50 VSUBS 0.026829f
C105 VN.n51 VSUBS 0.034524f
C106 VN.t3 VSUBS 2.97113f
C107 VN.t6 VSUBS 2.74867f
C108 VN.n52 VSUBS 1.03677f
C109 VN.n53 VSUBS 1.01496f
C110 VN.n54 VSUBS 0.259375f
C111 VN.n55 VSUBS 0.026829f
C112 VN.n56 VSUBS 0.049752f
C113 VN.n57 VSUBS 0.041227f
C114 VN.n58 VSUBS 0.036773f
C115 VN.n59 VSUBS 0.026829f
C116 VN.n60 VSUBS 0.026829f
C117 VN.n61 VSUBS 0.026829f
C118 VN.n62 VSUBS 0.037471f
C119 VN.n63 VSUBS 0.96259f
C120 VN.n64 VSUBS 0.037471f
C121 VN.n65 VSUBS 0.049752f
C122 VN.n66 VSUBS 0.026829f
C123 VN.n67 VSUBS 0.026829f
C124 VN.n68 VSUBS 0.026829f
C125 VN.n69 VSUBS 0.041227f
C126 VN.n70 VSUBS 0.049752f
C127 VN.n71 VSUBS 0.034524f
C128 VN.n72 VSUBS 0.026829f
C129 VN.n73 VSUBS 0.026829f
C130 VN.n74 VSUBS 0.040419f
C131 VN.n75 VSUBS 0.050217f
C132 VN.n76 VSUBS 0.031921f
C133 VN.n77 VSUBS 0.026829f
C134 VN.n78 VSUBS 0.026829f
C135 VN.n79 VSUBS 0.026829f
C136 VN.n80 VSUBS 0.049752f
C137 VN.n81 VSUBS 0.031577f
C138 VN.n82 VSUBS 1.04708f
C139 VN.n83 VSUBS 1.72422f
C140 B.n0 VSUBS 0.005557f
C141 B.n1 VSUBS 0.005557f
C142 B.n2 VSUBS 0.008787f
C143 B.n3 VSUBS 0.008787f
C144 B.n4 VSUBS 0.008787f
C145 B.n5 VSUBS 0.008787f
C146 B.n6 VSUBS 0.008787f
C147 B.n7 VSUBS 0.008787f
C148 B.n8 VSUBS 0.008787f
C149 B.n9 VSUBS 0.008787f
C150 B.n10 VSUBS 0.008787f
C151 B.n11 VSUBS 0.008787f
C152 B.n12 VSUBS 0.008787f
C153 B.n13 VSUBS 0.008787f
C154 B.n14 VSUBS 0.008787f
C155 B.n15 VSUBS 0.008787f
C156 B.n16 VSUBS 0.008787f
C157 B.n17 VSUBS 0.008787f
C158 B.n18 VSUBS 0.008787f
C159 B.n19 VSUBS 0.008787f
C160 B.n20 VSUBS 0.008787f
C161 B.n21 VSUBS 0.008787f
C162 B.n22 VSUBS 0.008787f
C163 B.n23 VSUBS 0.008787f
C164 B.n24 VSUBS 0.008787f
C165 B.n25 VSUBS 0.008787f
C166 B.n26 VSUBS 0.008787f
C167 B.n27 VSUBS 0.008787f
C168 B.n28 VSUBS 0.008787f
C169 B.n29 VSUBS 0.008787f
C170 B.n30 VSUBS 0.008787f
C171 B.n31 VSUBS 0.008787f
C172 B.n32 VSUBS 0.02024f
C173 B.n33 VSUBS 0.008787f
C174 B.n34 VSUBS 0.008787f
C175 B.n35 VSUBS 0.008787f
C176 B.n36 VSUBS 0.008787f
C177 B.n37 VSUBS 0.008787f
C178 B.n38 VSUBS 0.008787f
C179 B.n39 VSUBS 0.008787f
C180 B.n40 VSUBS 0.008787f
C181 B.n41 VSUBS 0.008787f
C182 B.n42 VSUBS 0.008787f
C183 B.n43 VSUBS 0.008787f
C184 B.n44 VSUBS 0.008787f
C185 B.n45 VSUBS 0.008787f
C186 B.n46 VSUBS 0.008787f
C187 B.n47 VSUBS 0.008787f
C188 B.n48 VSUBS 0.008787f
C189 B.n49 VSUBS 0.008787f
C190 B.n50 VSUBS 0.008787f
C191 B.n51 VSUBS 0.008787f
C192 B.n52 VSUBS 0.008787f
C193 B.n53 VSUBS 0.008787f
C194 B.n54 VSUBS 0.008787f
C195 B.n55 VSUBS 0.008787f
C196 B.n56 VSUBS 0.006073f
C197 B.n57 VSUBS 0.008787f
C198 B.t8 VSUBS 0.596895f
C199 B.t7 VSUBS 0.623828f
C200 B.t6 VSUBS 2.11647f
C201 B.n58 VSUBS 0.331144f
C202 B.n59 VSUBS 0.090388f
C203 B.n60 VSUBS 0.020359f
C204 B.n61 VSUBS 0.008787f
C205 B.n62 VSUBS 0.008787f
C206 B.n63 VSUBS 0.008787f
C207 B.n64 VSUBS 0.008787f
C208 B.t5 VSUBS 0.596879f
C209 B.t4 VSUBS 0.623814f
C210 B.t3 VSUBS 2.11647f
C211 B.n65 VSUBS 0.331157f
C212 B.n66 VSUBS 0.090404f
C213 B.n67 VSUBS 0.008787f
C214 B.n68 VSUBS 0.008787f
C215 B.n69 VSUBS 0.008787f
C216 B.n70 VSUBS 0.008787f
C217 B.n71 VSUBS 0.008787f
C218 B.n72 VSUBS 0.008787f
C219 B.n73 VSUBS 0.008787f
C220 B.n74 VSUBS 0.008787f
C221 B.n75 VSUBS 0.008787f
C222 B.n76 VSUBS 0.008787f
C223 B.n77 VSUBS 0.008787f
C224 B.n78 VSUBS 0.008787f
C225 B.n79 VSUBS 0.008787f
C226 B.n80 VSUBS 0.008787f
C227 B.n81 VSUBS 0.008787f
C228 B.n82 VSUBS 0.008787f
C229 B.n83 VSUBS 0.008787f
C230 B.n84 VSUBS 0.008787f
C231 B.n85 VSUBS 0.008787f
C232 B.n86 VSUBS 0.008787f
C233 B.n87 VSUBS 0.008787f
C234 B.n88 VSUBS 0.008787f
C235 B.n89 VSUBS 0.008787f
C236 B.n90 VSUBS 0.02024f
C237 B.n91 VSUBS 0.008787f
C238 B.n92 VSUBS 0.008787f
C239 B.n93 VSUBS 0.008787f
C240 B.n94 VSUBS 0.008787f
C241 B.n95 VSUBS 0.008787f
C242 B.n96 VSUBS 0.008787f
C243 B.n97 VSUBS 0.008787f
C244 B.n98 VSUBS 0.008787f
C245 B.n99 VSUBS 0.008787f
C246 B.n100 VSUBS 0.008787f
C247 B.n101 VSUBS 0.008787f
C248 B.n102 VSUBS 0.008787f
C249 B.n103 VSUBS 0.008787f
C250 B.n104 VSUBS 0.008787f
C251 B.n105 VSUBS 0.008787f
C252 B.n106 VSUBS 0.008787f
C253 B.n107 VSUBS 0.008787f
C254 B.n108 VSUBS 0.008787f
C255 B.n109 VSUBS 0.008787f
C256 B.n110 VSUBS 0.008787f
C257 B.n111 VSUBS 0.008787f
C258 B.n112 VSUBS 0.008787f
C259 B.n113 VSUBS 0.008787f
C260 B.n114 VSUBS 0.008787f
C261 B.n115 VSUBS 0.008787f
C262 B.n116 VSUBS 0.008787f
C263 B.n117 VSUBS 0.008787f
C264 B.n118 VSUBS 0.008787f
C265 B.n119 VSUBS 0.008787f
C266 B.n120 VSUBS 0.008787f
C267 B.n121 VSUBS 0.008787f
C268 B.n122 VSUBS 0.008787f
C269 B.n123 VSUBS 0.008787f
C270 B.n124 VSUBS 0.008787f
C271 B.n125 VSUBS 0.008787f
C272 B.n126 VSUBS 0.008787f
C273 B.n127 VSUBS 0.008787f
C274 B.n128 VSUBS 0.008787f
C275 B.n129 VSUBS 0.008787f
C276 B.n130 VSUBS 0.008787f
C277 B.n131 VSUBS 0.008787f
C278 B.n132 VSUBS 0.008787f
C279 B.n133 VSUBS 0.008787f
C280 B.n134 VSUBS 0.008787f
C281 B.n135 VSUBS 0.008787f
C282 B.n136 VSUBS 0.008787f
C283 B.n137 VSUBS 0.008787f
C284 B.n138 VSUBS 0.008787f
C285 B.n139 VSUBS 0.008787f
C286 B.n140 VSUBS 0.008787f
C287 B.n141 VSUBS 0.008787f
C288 B.n142 VSUBS 0.008787f
C289 B.n143 VSUBS 0.008787f
C290 B.n144 VSUBS 0.008787f
C291 B.n145 VSUBS 0.008787f
C292 B.n146 VSUBS 0.008787f
C293 B.n147 VSUBS 0.008787f
C294 B.n148 VSUBS 0.008787f
C295 B.n149 VSUBS 0.008787f
C296 B.n150 VSUBS 0.008787f
C297 B.n151 VSUBS 0.02024f
C298 B.n152 VSUBS 0.008787f
C299 B.n153 VSUBS 0.008787f
C300 B.n154 VSUBS 0.008787f
C301 B.n155 VSUBS 0.008787f
C302 B.n156 VSUBS 0.008787f
C303 B.n157 VSUBS 0.008787f
C304 B.n158 VSUBS 0.008787f
C305 B.n159 VSUBS 0.008787f
C306 B.n160 VSUBS 0.008787f
C307 B.n161 VSUBS 0.008787f
C308 B.n162 VSUBS 0.008787f
C309 B.n163 VSUBS 0.008787f
C310 B.n164 VSUBS 0.008787f
C311 B.n165 VSUBS 0.008787f
C312 B.n166 VSUBS 0.008787f
C313 B.n167 VSUBS 0.008787f
C314 B.n168 VSUBS 0.008787f
C315 B.n169 VSUBS 0.008787f
C316 B.n170 VSUBS 0.008787f
C317 B.n171 VSUBS 0.008787f
C318 B.n172 VSUBS 0.008787f
C319 B.n173 VSUBS 0.008787f
C320 B.n174 VSUBS 0.008787f
C321 B.n175 VSUBS 0.006073f
C322 B.n176 VSUBS 0.008787f
C323 B.n177 VSUBS 0.008787f
C324 B.n178 VSUBS 0.008787f
C325 B.n179 VSUBS 0.008787f
C326 B.n180 VSUBS 0.008787f
C327 B.t10 VSUBS 0.596895f
C328 B.t11 VSUBS 0.623828f
C329 B.t9 VSUBS 2.11647f
C330 B.n181 VSUBS 0.331144f
C331 B.n182 VSUBS 0.090388f
C332 B.n183 VSUBS 0.008787f
C333 B.n184 VSUBS 0.008787f
C334 B.n185 VSUBS 0.008787f
C335 B.n186 VSUBS 0.008787f
C336 B.n187 VSUBS 0.008787f
C337 B.n188 VSUBS 0.008787f
C338 B.n189 VSUBS 0.008787f
C339 B.n190 VSUBS 0.008787f
C340 B.n191 VSUBS 0.008787f
C341 B.n192 VSUBS 0.008787f
C342 B.n193 VSUBS 0.008787f
C343 B.n194 VSUBS 0.008787f
C344 B.n195 VSUBS 0.008787f
C345 B.n196 VSUBS 0.008787f
C346 B.n197 VSUBS 0.008787f
C347 B.n198 VSUBS 0.008787f
C348 B.n199 VSUBS 0.008787f
C349 B.n200 VSUBS 0.008787f
C350 B.n201 VSUBS 0.008787f
C351 B.n202 VSUBS 0.008787f
C352 B.n203 VSUBS 0.008787f
C353 B.n204 VSUBS 0.008787f
C354 B.n205 VSUBS 0.008787f
C355 B.n206 VSUBS 0.02024f
C356 B.n207 VSUBS 0.008787f
C357 B.n208 VSUBS 0.008787f
C358 B.n209 VSUBS 0.008787f
C359 B.n210 VSUBS 0.008787f
C360 B.n211 VSUBS 0.008787f
C361 B.n212 VSUBS 0.008787f
C362 B.n213 VSUBS 0.008787f
C363 B.n214 VSUBS 0.008787f
C364 B.n215 VSUBS 0.008787f
C365 B.n216 VSUBS 0.008787f
C366 B.n217 VSUBS 0.008787f
C367 B.n218 VSUBS 0.008787f
C368 B.n219 VSUBS 0.008787f
C369 B.n220 VSUBS 0.008787f
C370 B.n221 VSUBS 0.008787f
C371 B.n222 VSUBS 0.008787f
C372 B.n223 VSUBS 0.008787f
C373 B.n224 VSUBS 0.008787f
C374 B.n225 VSUBS 0.008787f
C375 B.n226 VSUBS 0.008787f
C376 B.n227 VSUBS 0.008787f
C377 B.n228 VSUBS 0.008787f
C378 B.n229 VSUBS 0.008787f
C379 B.n230 VSUBS 0.008787f
C380 B.n231 VSUBS 0.008787f
C381 B.n232 VSUBS 0.008787f
C382 B.n233 VSUBS 0.008787f
C383 B.n234 VSUBS 0.008787f
C384 B.n235 VSUBS 0.008787f
C385 B.n236 VSUBS 0.008787f
C386 B.n237 VSUBS 0.008787f
C387 B.n238 VSUBS 0.008787f
C388 B.n239 VSUBS 0.008787f
C389 B.n240 VSUBS 0.008787f
C390 B.n241 VSUBS 0.008787f
C391 B.n242 VSUBS 0.008787f
C392 B.n243 VSUBS 0.008787f
C393 B.n244 VSUBS 0.008787f
C394 B.n245 VSUBS 0.008787f
C395 B.n246 VSUBS 0.008787f
C396 B.n247 VSUBS 0.008787f
C397 B.n248 VSUBS 0.008787f
C398 B.n249 VSUBS 0.008787f
C399 B.n250 VSUBS 0.008787f
C400 B.n251 VSUBS 0.008787f
C401 B.n252 VSUBS 0.008787f
C402 B.n253 VSUBS 0.008787f
C403 B.n254 VSUBS 0.008787f
C404 B.n255 VSUBS 0.008787f
C405 B.n256 VSUBS 0.008787f
C406 B.n257 VSUBS 0.008787f
C407 B.n258 VSUBS 0.008787f
C408 B.n259 VSUBS 0.008787f
C409 B.n260 VSUBS 0.008787f
C410 B.n261 VSUBS 0.008787f
C411 B.n262 VSUBS 0.008787f
C412 B.n263 VSUBS 0.008787f
C413 B.n264 VSUBS 0.008787f
C414 B.n265 VSUBS 0.008787f
C415 B.n266 VSUBS 0.008787f
C416 B.n267 VSUBS 0.008787f
C417 B.n268 VSUBS 0.008787f
C418 B.n269 VSUBS 0.008787f
C419 B.n270 VSUBS 0.008787f
C420 B.n271 VSUBS 0.008787f
C421 B.n272 VSUBS 0.008787f
C422 B.n273 VSUBS 0.008787f
C423 B.n274 VSUBS 0.008787f
C424 B.n275 VSUBS 0.008787f
C425 B.n276 VSUBS 0.008787f
C426 B.n277 VSUBS 0.008787f
C427 B.n278 VSUBS 0.008787f
C428 B.n279 VSUBS 0.008787f
C429 B.n280 VSUBS 0.008787f
C430 B.n281 VSUBS 0.008787f
C431 B.n282 VSUBS 0.008787f
C432 B.n283 VSUBS 0.008787f
C433 B.n284 VSUBS 0.008787f
C434 B.n285 VSUBS 0.008787f
C435 B.n286 VSUBS 0.008787f
C436 B.n287 VSUBS 0.008787f
C437 B.n288 VSUBS 0.008787f
C438 B.n289 VSUBS 0.008787f
C439 B.n290 VSUBS 0.008787f
C440 B.n291 VSUBS 0.008787f
C441 B.n292 VSUBS 0.008787f
C442 B.n293 VSUBS 0.008787f
C443 B.n294 VSUBS 0.008787f
C444 B.n295 VSUBS 0.008787f
C445 B.n296 VSUBS 0.008787f
C446 B.n297 VSUBS 0.008787f
C447 B.n298 VSUBS 0.008787f
C448 B.n299 VSUBS 0.008787f
C449 B.n300 VSUBS 0.008787f
C450 B.n301 VSUBS 0.008787f
C451 B.n302 VSUBS 0.008787f
C452 B.n303 VSUBS 0.008787f
C453 B.n304 VSUBS 0.008787f
C454 B.n305 VSUBS 0.008787f
C455 B.n306 VSUBS 0.008787f
C456 B.n307 VSUBS 0.008787f
C457 B.n308 VSUBS 0.008787f
C458 B.n309 VSUBS 0.008787f
C459 B.n310 VSUBS 0.008787f
C460 B.n311 VSUBS 0.008787f
C461 B.n312 VSUBS 0.008787f
C462 B.n313 VSUBS 0.008787f
C463 B.n314 VSUBS 0.008787f
C464 B.n315 VSUBS 0.008787f
C465 B.n316 VSUBS 0.008787f
C466 B.n317 VSUBS 0.008787f
C467 B.n318 VSUBS 0.008787f
C468 B.n319 VSUBS 0.008787f
C469 B.n320 VSUBS 0.008787f
C470 B.n321 VSUBS 0.008787f
C471 B.n322 VSUBS 0.008787f
C472 B.n323 VSUBS 0.018785f
C473 B.n324 VSUBS 0.018785f
C474 B.n325 VSUBS 0.02024f
C475 B.n326 VSUBS 0.008787f
C476 B.n327 VSUBS 0.008787f
C477 B.n328 VSUBS 0.008787f
C478 B.n329 VSUBS 0.008787f
C479 B.n330 VSUBS 0.008787f
C480 B.n331 VSUBS 0.008787f
C481 B.n332 VSUBS 0.008787f
C482 B.n333 VSUBS 0.008787f
C483 B.n334 VSUBS 0.008787f
C484 B.n335 VSUBS 0.008787f
C485 B.n336 VSUBS 0.008787f
C486 B.n337 VSUBS 0.008787f
C487 B.n338 VSUBS 0.008787f
C488 B.n339 VSUBS 0.008787f
C489 B.n340 VSUBS 0.008787f
C490 B.n341 VSUBS 0.008787f
C491 B.n342 VSUBS 0.008787f
C492 B.n343 VSUBS 0.008787f
C493 B.n344 VSUBS 0.008787f
C494 B.n345 VSUBS 0.008787f
C495 B.n346 VSUBS 0.008787f
C496 B.n347 VSUBS 0.008787f
C497 B.n348 VSUBS 0.008787f
C498 B.n349 VSUBS 0.008787f
C499 B.n350 VSUBS 0.008787f
C500 B.n351 VSUBS 0.008787f
C501 B.n352 VSUBS 0.008787f
C502 B.n353 VSUBS 0.008787f
C503 B.n354 VSUBS 0.008787f
C504 B.n355 VSUBS 0.008787f
C505 B.n356 VSUBS 0.008787f
C506 B.n357 VSUBS 0.008787f
C507 B.n358 VSUBS 0.008787f
C508 B.n359 VSUBS 0.008787f
C509 B.n360 VSUBS 0.008787f
C510 B.n361 VSUBS 0.008787f
C511 B.n362 VSUBS 0.008787f
C512 B.n363 VSUBS 0.008787f
C513 B.n364 VSUBS 0.008787f
C514 B.n365 VSUBS 0.008787f
C515 B.n366 VSUBS 0.008787f
C516 B.n367 VSUBS 0.008787f
C517 B.n368 VSUBS 0.008787f
C518 B.n369 VSUBS 0.008787f
C519 B.n370 VSUBS 0.008787f
C520 B.n371 VSUBS 0.008787f
C521 B.n372 VSUBS 0.008787f
C522 B.n373 VSUBS 0.008787f
C523 B.n374 VSUBS 0.008787f
C524 B.n375 VSUBS 0.008787f
C525 B.n376 VSUBS 0.008787f
C526 B.n377 VSUBS 0.008787f
C527 B.n378 VSUBS 0.008787f
C528 B.n379 VSUBS 0.008787f
C529 B.n380 VSUBS 0.008787f
C530 B.n381 VSUBS 0.008787f
C531 B.n382 VSUBS 0.008787f
C532 B.n383 VSUBS 0.008787f
C533 B.n384 VSUBS 0.008787f
C534 B.n385 VSUBS 0.008787f
C535 B.n386 VSUBS 0.008787f
C536 B.n387 VSUBS 0.008787f
C537 B.n388 VSUBS 0.008787f
C538 B.n389 VSUBS 0.008787f
C539 B.n390 VSUBS 0.008787f
C540 B.n391 VSUBS 0.008787f
C541 B.n392 VSUBS 0.008787f
C542 B.n393 VSUBS 0.008787f
C543 B.n394 VSUBS 0.008787f
C544 B.n395 VSUBS 0.008787f
C545 B.n396 VSUBS 0.008787f
C546 B.n397 VSUBS 0.006073f
C547 B.n398 VSUBS 0.020359f
C548 B.n399 VSUBS 0.007107f
C549 B.n400 VSUBS 0.008787f
C550 B.n401 VSUBS 0.008787f
C551 B.n402 VSUBS 0.008787f
C552 B.n403 VSUBS 0.008787f
C553 B.n404 VSUBS 0.008787f
C554 B.n405 VSUBS 0.008787f
C555 B.n406 VSUBS 0.008787f
C556 B.n407 VSUBS 0.008787f
C557 B.n408 VSUBS 0.008787f
C558 B.n409 VSUBS 0.008787f
C559 B.n410 VSUBS 0.008787f
C560 B.t1 VSUBS 0.596879f
C561 B.t2 VSUBS 0.623814f
C562 B.t0 VSUBS 2.11647f
C563 B.n411 VSUBS 0.331157f
C564 B.n412 VSUBS 0.090404f
C565 B.n413 VSUBS 0.020359f
C566 B.n414 VSUBS 0.007107f
C567 B.n415 VSUBS 0.008787f
C568 B.n416 VSUBS 0.008787f
C569 B.n417 VSUBS 0.008787f
C570 B.n418 VSUBS 0.008787f
C571 B.n419 VSUBS 0.008787f
C572 B.n420 VSUBS 0.008787f
C573 B.n421 VSUBS 0.008787f
C574 B.n422 VSUBS 0.008787f
C575 B.n423 VSUBS 0.008787f
C576 B.n424 VSUBS 0.008787f
C577 B.n425 VSUBS 0.008787f
C578 B.n426 VSUBS 0.008787f
C579 B.n427 VSUBS 0.008787f
C580 B.n428 VSUBS 0.008787f
C581 B.n429 VSUBS 0.008787f
C582 B.n430 VSUBS 0.008787f
C583 B.n431 VSUBS 0.008787f
C584 B.n432 VSUBS 0.008787f
C585 B.n433 VSUBS 0.008787f
C586 B.n434 VSUBS 0.008787f
C587 B.n435 VSUBS 0.008787f
C588 B.n436 VSUBS 0.008787f
C589 B.n437 VSUBS 0.008787f
C590 B.n438 VSUBS 0.008787f
C591 B.n439 VSUBS 0.008787f
C592 B.n440 VSUBS 0.008787f
C593 B.n441 VSUBS 0.008787f
C594 B.n442 VSUBS 0.008787f
C595 B.n443 VSUBS 0.008787f
C596 B.n444 VSUBS 0.008787f
C597 B.n445 VSUBS 0.008787f
C598 B.n446 VSUBS 0.008787f
C599 B.n447 VSUBS 0.008787f
C600 B.n448 VSUBS 0.008787f
C601 B.n449 VSUBS 0.008787f
C602 B.n450 VSUBS 0.008787f
C603 B.n451 VSUBS 0.008787f
C604 B.n452 VSUBS 0.008787f
C605 B.n453 VSUBS 0.008787f
C606 B.n454 VSUBS 0.008787f
C607 B.n455 VSUBS 0.008787f
C608 B.n456 VSUBS 0.008787f
C609 B.n457 VSUBS 0.008787f
C610 B.n458 VSUBS 0.008787f
C611 B.n459 VSUBS 0.008787f
C612 B.n460 VSUBS 0.008787f
C613 B.n461 VSUBS 0.008787f
C614 B.n462 VSUBS 0.008787f
C615 B.n463 VSUBS 0.008787f
C616 B.n464 VSUBS 0.008787f
C617 B.n465 VSUBS 0.008787f
C618 B.n466 VSUBS 0.008787f
C619 B.n467 VSUBS 0.008787f
C620 B.n468 VSUBS 0.008787f
C621 B.n469 VSUBS 0.008787f
C622 B.n470 VSUBS 0.008787f
C623 B.n471 VSUBS 0.008787f
C624 B.n472 VSUBS 0.008787f
C625 B.n473 VSUBS 0.008787f
C626 B.n474 VSUBS 0.008787f
C627 B.n475 VSUBS 0.008787f
C628 B.n476 VSUBS 0.008787f
C629 B.n477 VSUBS 0.008787f
C630 B.n478 VSUBS 0.008787f
C631 B.n479 VSUBS 0.008787f
C632 B.n480 VSUBS 0.008787f
C633 B.n481 VSUBS 0.008787f
C634 B.n482 VSUBS 0.008787f
C635 B.n483 VSUBS 0.008787f
C636 B.n484 VSUBS 0.008787f
C637 B.n485 VSUBS 0.008787f
C638 B.n486 VSUBS 0.008787f
C639 B.n487 VSUBS 0.008787f
C640 B.n488 VSUBS 0.02024f
C641 B.n489 VSUBS 0.018785f
C642 B.n490 VSUBS 0.018785f
C643 B.n491 VSUBS 0.008787f
C644 B.n492 VSUBS 0.008787f
C645 B.n493 VSUBS 0.008787f
C646 B.n494 VSUBS 0.008787f
C647 B.n495 VSUBS 0.008787f
C648 B.n496 VSUBS 0.008787f
C649 B.n497 VSUBS 0.008787f
C650 B.n498 VSUBS 0.008787f
C651 B.n499 VSUBS 0.008787f
C652 B.n500 VSUBS 0.008787f
C653 B.n501 VSUBS 0.008787f
C654 B.n502 VSUBS 0.008787f
C655 B.n503 VSUBS 0.008787f
C656 B.n504 VSUBS 0.008787f
C657 B.n505 VSUBS 0.008787f
C658 B.n506 VSUBS 0.008787f
C659 B.n507 VSUBS 0.008787f
C660 B.n508 VSUBS 0.008787f
C661 B.n509 VSUBS 0.008787f
C662 B.n510 VSUBS 0.008787f
C663 B.n511 VSUBS 0.008787f
C664 B.n512 VSUBS 0.008787f
C665 B.n513 VSUBS 0.008787f
C666 B.n514 VSUBS 0.008787f
C667 B.n515 VSUBS 0.008787f
C668 B.n516 VSUBS 0.008787f
C669 B.n517 VSUBS 0.008787f
C670 B.n518 VSUBS 0.008787f
C671 B.n519 VSUBS 0.008787f
C672 B.n520 VSUBS 0.008787f
C673 B.n521 VSUBS 0.008787f
C674 B.n522 VSUBS 0.008787f
C675 B.n523 VSUBS 0.008787f
C676 B.n524 VSUBS 0.008787f
C677 B.n525 VSUBS 0.008787f
C678 B.n526 VSUBS 0.008787f
C679 B.n527 VSUBS 0.008787f
C680 B.n528 VSUBS 0.008787f
C681 B.n529 VSUBS 0.008787f
C682 B.n530 VSUBS 0.008787f
C683 B.n531 VSUBS 0.008787f
C684 B.n532 VSUBS 0.008787f
C685 B.n533 VSUBS 0.008787f
C686 B.n534 VSUBS 0.008787f
C687 B.n535 VSUBS 0.008787f
C688 B.n536 VSUBS 0.008787f
C689 B.n537 VSUBS 0.008787f
C690 B.n538 VSUBS 0.008787f
C691 B.n539 VSUBS 0.008787f
C692 B.n540 VSUBS 0.008787f
C693 B.n541 VSUBS 0.008787f
C694 B.n542 VSUBS 0.008787f
C695 B.n543 VSUBS 0.008787f
C696 B.n544 VSUBS 0.008787f
C697 B.n545 VSUBS 0.008787f
C698 B.n546 VSUBS 0.008787f
C699 B.n547 VSUBS 0.008787f
C700 B.n548 VSUBS 0.008787f
C701 B.n549 VSUBS 0.008787f
C702 B.n550 VSUBS 0.008787f
C703 B.n551 VSUBS 0.008787f
C704 B.n552 VSUBS 0.008787f
C705 B.n553 VSUBS 0.008787f
C706 B.n554 VSUBS 0.008787f
C707 B.n555 VSUBS 0.008787f
C708 B.n556 VSUBS 0.008787f
C709 B.n557 VSUBS 0.008787f
C710 B.n558 VSUBS 0.008787f
C711 B.n559 VSUBS 0.008787f
C712 B.n560 VSUBS 0.008787f
C713 B.n561 VSUBS 0.008787f
C714 B.n562 VSUBS 0.008787f
C715 B.n563 VSUBS 0.008787f
C716 B.n564 VSUBS 0.008787f
C717 B.n565 VSUBS 0.008787f
C718 B.n566 VSUBS 0.008787f
C719 B.n567 VSUBS 0.008787f
C720 B.n568 VSUBS 0.008787f
C721 B.n569 VSUBS 0.008787f
C722 B.n570 VSUBS 0.008787f
C723 B.n571 VSUBS 0.008787f
C724 B.n572 VSUBS 0.008787f
C725 B.n573 VSUBS 0.008787f
C726 B.n574 VSUBS 0.008787f
C727 B.n575 VSUBS 0.008787f
C728 B.n576 VSUBS 0.008787f
C729 B.n577 VSUBS 0.008787f
C730 B.n578 VSUBS 0.008787f
C731 B.n579 VSUBS 0.008787f
C732 B.n580 VSUBS 0.008787f
C733 B.n581 VSUBS 0.008787f
C734 B.n582 VSUBS 0.008787f
C735 B.n583 VSUBS 0.008787f
C736 B.n584 VSUBS 0.008787f
C737 B.n585 VSUBS 0.008787f
C738 B.n586 VSUBS 0.008787f
C739 B.n587 VSUBS 0.008787f
C740 B.n588 VSUBS 0.008787f
C741 B.n589 VSUBS 0.008787f
C742 B.n590 VSUBS 0.008787f
C743 B.n591 VSUBS 0.008787f
C744 B.n592 VSUBS 0.008787f
C745 B.n593 VSUBS 0.008787f
C746 B.n594 VSUBS 0.008787f
C747 B.n595 VSUBS 0.008787f
C748 B.n596 VSUBS 0.008787f
C749 B.n597 VSUBS 0.008787f
C750 B.n598 VSUBS 0.008787f
C751 B.n599 VSUBS 0.008787f
C752 B.n600 VSUBS 0.008787f
C753 B.n601 VSUBS 0.008787f
C754 B.n602 VSUBS 0.008787f
C755 B.n603 VSUBS 0.008787f
C756 B.n604 VSUBS 0.008787f
C757 B.n605 VSUBS 0.008787f
C758 B.n606 VSUBS 0.008787f
C759 B.n607 VSUBS 0.008787f
C760 B.n608 VSUBS 0.008787f
C761 B.n609 VSUBS 0.008787f
C762 B.n610 VSUBS 0.008787f
C763 B.n611 VSUBS 0.008787f
C764 B.n612 VSUBS 0.008787f
C765 B.n613 VSUBS 0.008787f
C766 B.n614 VSUBS 0.008787f
C767 B.n615 VSUBS 0.008787f
C768 B.n616 VSUBS 0.008787f
C769 B.n617 VSUBS 0.008787f
C770 B.n618 VSUBS 0.008787f
C771 B.n619 VSUBS 0.008787f
C772 B.n620 VSUBS 0.008787f
C773 B.n621 VSUBS 0.008787f
C774 B.n622 VSUBS 0.008787f
C775 B.n623 VSUBS 0.008787f
C776 B.n624 VSUBS 0.008787f
C777 B.n625 VSUBS 0.008787f
C778 B.n626 VSUBS 0.008787f
C779 B.n627 VSUBS 0.008787f
C780 B.n628 VSUBS 0.008787f
C781 B.n629 VSUBS 0.008787f
C782 B.n630 VSUBS 0.008787f
C783 B.n631 VSUBS 0.008787f
C784 B.n632 VSUBS 0.008787f
C785 B.n633 VSUBS 0.008787f
C786 B.n634 VSUBS 0.008787f
C787 B.n635 VSUBS 0.008787f
C788 B.n636 VSUBS 0.008787f
C789 B.n637 VSUBS 0.008787f
C790 B.n638 VSUBS 0.008787f
C791 B.n639 VSUBS 0.008787f
C792 B.n640 VSUBS 0.008787f
C793 B.n641 VSUBS 0.008787f
C794 B.n642 VSUBS 0.008787f
C795 B.n643 VSUBS 0.008787f
C796 B.n644 VSUBS 0.008787f
C797 B.n645 VSUBS 0.008787f
C798 B.n646 VSUBS 0.008787f
C799 B.n647 VSUBS 0.008787f
C800 B.n648 VSUBS 0.008787f
C801 B.n649 VSUBS 0.008787f
C802 B.n650 VSUBS 0.008787f
C803 B.n651 VSUBS 0.008787f
C804 B.n652 VSUBS 0.008787f
C805 B.n653 VSUBS 0.008787f
C806 B.n654 VSUBS 0.008787f
C807 B.n655 VSUBS 0.008787f
C808 B.n656 VSUBS 0.008787f
C809 B.n657 VSUBS 0.008787f
C810 B.n658 VSUBS 0.008787f
C811 B.n659 VSUBS 0.008787f
C812 B.n660 VSUBS 0.008787f
C813 B.n661 VSUBS 0.008787f
C814 B.n662 VSUBS 0.008787f
C815 B.n663 VSUBS 0.008787f
C816 B.n664 VSUBS 0.008787f
C817 B.n665 VSUBS 0.008787f
C818 B.n666 VSUBS 0.008787f
C819 B.n667 VSUBS 0.008787f
C820 B.n668 VSUBS 0.008787f
C821 B.n669 VSUBS 0.018785f
C822 B.n670 VSUBS 0.019911f
C823 B.n671 VSUBS 0.019115f
C824 B.n672 VSUBS 0.008787f
C825 B.n673 VSUBS 0.008787f
C826 B.n674 VSUBS 0.008787f
C827 B.n675 VSUBS 0.008787f
C828 B.n676 VSUBS 0.008787f
C829 B.n677 VSUBS 0.008787f
C830 B.n678 VSUBS 0.008787f
C831 B.n679 VSUBS 0.008787f
C832 B.n680 VSUBS 0.008787f
C833 B.n681 VSUBS 0.008787f
C834 B.n682 VSUBS 0.008787f
C835 B.n683 VSUBS 0.008787f
C836 B.n684 VSUBS 0.008787f
C837 B.n685 VSUBS 0.008787f
C838 B.n686 VSUBS 0.008787f
C839 B.n687 VSUBS 0.008787f
C840 B.n688 VSUBS 0.008787f
C841 B.n689 VSUBS 0.008787f
C842 B.n690 VSUBS 0.008787f
C843 B.n691 VSUBS 0.008787f
C844 B.n692 VSUBS 0.008787f
C845 B.n693 VSUBS 0.008787f
C846 B.n694 VSUBS 0.008787f
C847 B.n695 VSUBS 0.008787f
C848 B.n696 VSUBS 0.008787f
C849 B.n697 VSUBS 0.008787f
C850 B.n698 VSUBS 0.008787f
C851 B.n699 VSUBS 0.008787f
C852 B.n700 VSUBS 0.008787f
C853 B.n701 VSUBS 0.008787f
C854 B.n702 VSUBS 0.008787f
C855 B.n703 VSUBS 0.008787f
C856 B.n704 VSUBS 0.008787f
C857 B.n705 VSUBS 0.008787f
C858 B.n706 VSUBS 0.008787f
C859 B.n707 VSUBS 0.008787f
C860 B.n708 VSUBS 0.008787f
C861 B.n709 VSUBS 0.008787f
C862 B.n710 VSUBS 0.008787f
C863 B.n711 VSUBS 0.008787f
C864 B.n712 VSUBS 0.008787f
C865 B.n713 VSUBS 0.008787f
C866 B.n714 VSUBS 0.008787f
C867 B.n715 VSUBS 0.008787f
C868 B.n716 VSUBS 0.008787f
C869 B.n717 VSUBS 0.008787f
C870 B.n718 VSUBS 0.008787f
C871 B.n719 VSUBS 0.008787f
C872 B.n720 VSUBS 0.008787f
C873 B.n721 VSUBS 0.008787f
C874 B.n722 VSUBS 0.008787f
C875 B.n723 VSUBS 0.008787f
C876 B.n724 VSUBS 0.008787f
C877 B.n725 VSUBS 0.008787f
C878 B.n726 VSUBS 0.008787f
C879 B.n727 VSUBS 0.008787f
C880 B.n728 VSUBS 0.008787f
C881 B.n729 VSUBS 0.008787f
C882 B.n730 VSUBS 0.008787f
C883 B.n731 VSUBS 0.008787f
C884 B.n732 VSUBS 0.008787f
C885 B.n733 VSUBS 0.008787f
C886 B.n734 VSUBS 0.008787f
C887 B.n735 VSUBS 0.008787f
C888 B.n736 VSUBS 0.008787f
C889 B.n737 VSUBS 0.008787f
C890 B.n738 VSUBS 0.008787f
C891 B.n739 VSUBS 0.008787f
C892 B.n740 VSUBS 0.008787f
C893 B.n741 VSUBS 0.008787f
C894 B.n742 VSUBS 0.008787f
C895 B.n743 VSUBS 0.006073f
C896 B.n744 VSUBS 0.020359f
C897 B.n745 VSUBS 0.007107f
C898 B.n746 VSUBS 0.008787f
C899 B.n747 VSUBS 0.008787f
C900 B.n748 VSUBS 0.008787f
C901 B.n749 VSUBS 0.008787f
C902 B.n750 VSUBS 0.008787f
C903 B.n751 VSUBS 0.008787f
C904 B.n752 VSUBS 0.008787f
C905 B.n753 VSUBS 0.008787f
C906 B.n754 VSUBS 0.008787f
C907 B.n755 VSUBS 0.008787f
C908 B.n756 VSUBS 0.008787f
C909 B.n757 VSUBS 0.007107f
C910 B.n758 VSUBS 0.008787f
C911 B.n759 VSUBS 0.008787f
C912 B.n760 VSUBS 0.008787f
C913 B.n761 VSUBS 0.008787f
C914 B.n762 VSUBS 0.008787f
C915 B.n763 VSUBS 0.008787f
C916 B.n764 VSUBS 0.008787f
C917 B.n765 VSUBS 0.008787f
C918 B.n766 VSUBS 0.008787f
C919 B.n767 VSUBS 0.008787f
C920 B.n768 VSUBS 0.008787f
C921 B.n769 VSUBS 0.008787f
C922 B.n770 VSUBS 0.008787f
C923 B.n771 VSUBS 0.008787f
C924 B.n772 VSUBS 0.008787f
C925 B.n773 VSUBS 0.008787f
C926 B.n774 VSUBS 0.008787f
C927 B.n775 VSUBS 0.008787f
C928 B.n776 VSUBS 0.008787f
C929 B.n777 VSUBS 0.008787f
C930 B.n778 VSUBS 0.008787f
C931 B.n779 VSUBS 0.008787f
C932 B.n780 VSUBS 0.008787f
C933 B.n781 VSUBS 0.008787f
C934 B.n782 VSUBS 0.008787f
C935 B.n783 VSUBS 0.008787f
C936 B.n784 VSUBS 0.008787f
C937 B.n785 VSUBS 0.008787f
C938 B.n786 VSUBS 0.008787f
C939 B.n787 VSUBS 0.008787f
C940 B.n788 VSUBS 0.008787f
C941 B.n789 VSUBS 0.008787f
C942 B.n790 VSUBS 0.008787f
C943 B.n791 VSUBS 0.008787f
C944 B.n792 VSUBS 0.008787f
C945 B.n793 VSUBS 0.008787f
C946 B.n794 VSUBS 0.008787f
C947 B.n795 VSUBS 0.008787f
C948 B.n796 VSUBS 0.008787f
C949 B.n797 VSUBS 0.008787f
C950 B.n798 VSUBS 0.008787f
C951 B.n799 VSUBS 0.008787f
C952 B.n800 VSUBS 0.008787f
C953 B.n801 VSUBS 0.008787f
C954 B.n802 VSUBS 0.008787f
C955 B.n803 VSUBS 0.008787f
C956 B.n804 VSUBS 0.008787f
C957 B.n805 VSUBS 0.008787f
C958 B.n806 VSUBS 0.008787f
C959 B.n807 VSUBS 0.008787f
C960 B.n808 VSUBS 0.008787f
C961 B.n809 VSUBS 0.008787f
C962 B.n810 VSUBS 0.008787f
C963 B.n811 VSUBS 0.008787f
C964 B.n812 VSUBS 0.008787f
C965 B.n813 VSUBS 0.008787f
C966 B.n814 VSUBS 0.008787f
C967 B.n815 VSUBS 0.008787f
C968 B.n816 VSUBS 0.008787f
C969 B.n817 VSUBS 0.008787f
C970 B.n818 VSUBS 0.008787f
C971 B.n819 VSUBS 0.008787f
C972 B.n820 VSUBS 0.008787f
C973 B.n821 VSUBS 0.008787f
C974 B.n822 VSUBS 0.008787f
C975 B.n823 VSUBS 0.008787f
C976 B.n824 VSUBS 0.008787f
C977 B.n825 VSUBS 0.008787f
C978 B.n826 VSUBS 0.008787f
C979 B.n827 VSUBS 0.008787f
C980 B.n828 VSUBS 0.008787f
C981 B.n829 VSUBS 0.008787f
C982 B.n830 VSUBS 0.008787f
C983 B.n831 VSUBS 0.02024f
C984 B.n832 VSUBS 0.018785f
C985 B.n833 VSUBS 0.018785f
C986 B.n834 VSUBS 0.008787f
C987 B.n835 VSUBS 0.008787f
C988 B.n836 VSUBS 0.008787f
C989 B.n837 VSUBS 0.008787f
C990 B.n838 VSUBS 0.008787f
C991 B.n839 VSUBS 0.008787f
C992 B.n840 VSUBS 0.008787f
C993 B.n841 VSUBS 0.008787f
C994 B.n842 VSUBS 0.008787f
C995 B.n843 VSUBS 0.008787f
C996 B.n844 VSUBS 0.008787f
C997 B.n845 VSUBS 0.008787f
C998 B.n846 VSUBS 0.008787f
C999 B.n847 VSUBS 0.008787f
C1000 B.n848 VSUBS 0.008787f
C1001 B.n849 VSUBS 0.008787f
C1002 B.n850 VSUBS 0.008787f
C1003 B.n851 VSUBS 0.008787f
C1004 B.n852 VSUBS 0.008787f
C1005 B.n853 VSUBS 0.008787f
C1006 B.n854 VSUBS 0.008787f
C1007 B.n855 VSUBS 0.008787f
C1008 B.n856 VSUBS 0.008787f
C1009 B.n857 VSUBS 0.008787f
C1010 B.n858 VSUBS 0.008787f
C1011 B.n859 VSUBS 0.008787f
C1012 B.n860 VSUBS 0.008787f
C1013 B.n861 VSUBS 0.008787f
C1014 B.n862 VSUBS 0.008787f
C1015 B.n863 VSUBS 0.008787f
C1016 B.n864 VSUBS 0.008787f
C1017 B.n865 VSUBS 0.008787f
C1018 B.n866 VSUBS 0.008787f
C1019 B.n867 VSUBS 0.008787f
C1020 B.n868 VSUBS 0.008787f
C1021 B.n869 VSUBS 0.008787f
C1022 B.n870 VSUBS 0.008787f
C1023 B.n871 VSUBS 0.008787f
C1024 B.n872 VSUBS 0.008787f
C1025 B.n873 VSUBS 0.008787f
C1026 B.n874 VSUBS 0.008787f
C1027 B.n875 VSUBS 0.008787f
C1028 B.n876 VSUBS 0.008787f
C1029 B.n877 VSUBS 0.008787f
C1030 B.n878 VSUBS 0.008787f
C1031 B.n879 VSUBS 0.008787f
C1032 B.n880 VSUBS 0.008787f
C1033 B.n881 VSUBS 0.008787f
C1034 B.n882 VSUBS 0.008787f
C1035 B.n883 VSUBS 0.008787f
C1036 B.n884 VSUBS 0.008787f
C1037 B.n885 VSUBS 0.008787f
C1038 B.n886 VSUBS 0.008787f
C1039 B.n887 VSUBS 0.008787f
C1040 B.n888 VSUBS 0.008787f
C1041 B.n889 VSUBS 0.008787f
C1042 B.n890 VSUBS 0.008787f
C1043 B.n891 VSUBS 0.008787f
C1044 B.n892 VSUBS 0.008787f
C1045 B.n893 VSUBS 0.008787f
C1046 B.n894 VSUBS 0.008787f
C1047 B.n895 VSUBS 0.008787f
C1048 B.n896 VSUBS 0.008787f
C1049 B.n897 VSUBS 0.008787f
C1050 B.n898 VSUBS 0.008787f
C1051 B.n899 VSUBS 0.008787f
C1052 B.n900 VSUBS 0.008787f
C1053 B.n901 VSUBS 0.008787f
C1054 B.n902 VSUBS 0.008787f
C1055 B.n903 VSUBS 0.008787f
C1056 B.n904 VSUBS 0.008787f
C1057 B.n905 VSUBS 0.008787f
C1058 B.n906 VSUBS 0.008787f
C1059 B.n907 VSUBS 0.008787f
C1060 B.n908 VSUBS 0.008787f
C1061 B.n909 VSUBS 0.008787f
C1062 B.n910 VSUBS 0.008787f
C1063 B.n911 VSUBS 0.008787f
C1064 B.n912 VSUBS 0.008787f
C1065 B.n913 VSUBS 0.008787f
C1066 B.n914 VSUBS 0.008787f
C1067 B.n915 VSUBS 0.008787f
C1068 B.n916 VSUBS 0.008787f
C1069 B.n917 VSUBS 0.008787f
C1070 B.n918 VSUBS 0.008787f
C1071 B.n919 VSUBS 0.008787f
C1072 B.n920 VSUBS 0.008787f
C1073 B.n921 VSUBS 0.008787f
C1074 B.n922 VSUBS 0.008787f
C1075 B.n923 VSUBS 0.019897f
C1076 VDD1.t4 VSUBS 3.52752f
C1077 VDD1.t2 VSUBS 0.332938f
C1078 VDD1.t0 VSUBS 0.332938f
C1079 VDD1.n0 VSUBS 2.68907f
C1080 VDD1.n1 VSUBS 1.73408f
C1081 VDD1.t8 VSUBS 3.5275f
C1082 VDD1.t7 VSUBS 0.332938f
C1083 VDD1.t9 VSUBS 0.332938f
C1084 VDD1.n2 VSUBS 2.68906f
C1085 VDD1.n3 VSUBS 1.72453f
C1086 VDD1.t1 VSUBS 0.332938f
C1087 VDD1.t6 VSUBS 0.332938f
C1088 VDD1.n4 VSUBS 2.7135f
C1089 VDD1.n5 VSUBS 4.04726f
C1090 VDD1.t3 VSUBS 0.332938f
C1091 VDD1.t5 VSUBS 0.332938f
C1092 VDD1.n6 VSUBS 2.68906f
C1093 VDD1.n7 VSUBS 4.25497f
C1094 VTAIL.t7 VSUBS 0.319495f
C1095 VTAIL.t4 VSUBS 0.319495f
C1096 VTAIL.n0 VSUBS 2.42251f
C1097 VTAIL.n1 VSUBS 0.986743f
C1098 VTAIL.t12 VSUBS 3.17719f
C1099 VTAIL.n2 VSUBS 1.15569f
C1100 VTAIL.t11 VSUBS 0.319495f
C1101 VTAIL.t9 VSUBS 0.319495f
C1102 VTAIL.n3 VSUBS 2.42251f
C1103 VTAIL.n4 VSUBS 1.11146f
C1104 VTAIL.t17 VSUBS 0.319495f
C1105 VTAIL.t13 VSUBS 0.319495f
C1106 VTAIL.n5 VSUBS 2.42251f
C1107 VTAIL.n6 VSUBS 2.84778f
C1108 VTAIL.t5 VSUBS 0.319495f
C1109 VTAIL.t19 VSUBS 0.319495f
C1110 VTAIL.n7 VSUBS 2.42252f
C1111 VTAIL.n8 VSUBS 2.84777f
C1112 VTAIL.t2 VSUBS 0.319495f
C1113 VTAIL.t3 VSUBS 0.319495f
C1114 VTAIL.n9 VSUBS 2.42252f
C1115 VTAIL.n10 VSUBS 1.11146f
C1116 VTAIL.t0 VSUBS 3.17722f
C1117 VTAIL.n11 VSUBS 1.15566f
C1118 VTAIL.t18 VSUBS 0.319495f
C1119 VTAIL.t16 VSUBS 0.319495f
C1120 VTAIL.n12 VSUBS 2.42252f
C1121 VTAIL.n13 VSUBS 1.03901f
C1122 VTAIL.t14 VSUBS 0.319495f
C1123 VTAIL.t15 VSUBS 0.319495f
C1124 VTAIL.n14 VSUBS 2.42252f
C1125 VTAIL.n15 VSUBS 1.11146f
C1126 VTAIL.t10 VSUBS 3.17719f
C1127 VTAIL.n16 VSUBS 2.73419f
C1128 VTAIL.t6 VSUBS 3.17719f
C1129 VTAIL.n17 VSUBS 2.73419f
C1130 VTAIL.t1 VSUBS 0.319495f
C1131 VTAIL.t8 VSUBS 0.319495f
C1132 VTAIL.n18 VSUBS 2.42251f
C1133 VTAIL.n19 VSUBS 0.933487f
C1134 VP.n0 VSUBS 0.037951f
C1135 VP.t3 VSUBS 2.94928f
C1136 VP.n1 VSUBS 0.048944f
C1137 VP.n2 VSUBS 0.028787f
C1138 VP.t8 VSUBS 2.94928f
C1139 VP.n3 VSUBS 1.03284f
C1140 VP.n4 VSUBS 0.028787f
C1141 VP.n5 VSUBS 0.039457f
C1142 VP.n6 VSUBS 0.028787f
C1143 VP.t0 VSUBS 2.94928f
C1144 VP.n7 VSUBS 0.053383f
C1145 VP.n8 VSUBS 0.028787f
C1146 VP.n9 VSUBS 0.037044f
C1147 VP.n10 VSUBS 0.028787f
C1148 VP.n11 VSUBS 0.048944f
C1149 VP.n12 VSUBS 0.037951f
C1150 VP.t1 VSUBS 2.94928f
C1151 VP.n13 VSUBS 0.037951f
C1152 VP.t4 VSUBS 2.94928f
C1153 VP.n14 VSUBS 0.048944f
C1154 VP.n15 VSUBS 0.028787f
C1155 VP.t6 VSUBS 2.94928f
C1156 VP.n16 VSUBS 1.03284f
C1157 VP.n17 VSUBS 0.028787f
C1158 VP.n18 VSUBS 0.039457f
C1159 VP.n19 VSUBS 0.028787f
C1160 VP.t9 VSUBS 2.94928f
C1161 VP.n20 VSUBS 0.053383f
C1162 VP.n21 VSUBS 0.028787f
C1163 VP.n22 VSUBS 0.037044f
C1164 VP.t5 VSUBS 3.18797f
C1165 VP.t7 VSUBS 2.94928f
C1166 VP.n23 VSUBS 1.11243f
C1167 VP.n24 VSUBS 1.08904f
C1168 VP.n25 VSUBS 0.278306f
C1169 VP.n26 VSUBS 0.028787f
C1170 VP.n27 VSUBS 0.053383f
C1171 VP.n28 VSUBS 0.044236f
C1172 VP.n29 VSUBS 0.039457f
C1173 VP.n30 VSUBS 0.028787f
C1174 VP.n31 VSUBS 0.028787f
C1175 VP.n32 VSUBS 0.028787f
C1176 VP.n33 VSUBS 0.040206f
C1177 VP.n34 VSUBS 1.03284f
C1178 VP.n35 VSUBS 0.040206f
C1179 VP.n36 VSUBS 0.053383f
C1180 VP.n37 VSUBS 0.028787f
C1181 VP.n38 VSUBS 0.028787f
C1182 VP.n39 VSUBS 0.028787f
C1183 VP.n40 VSUBS 0.044236f
C1184 VP.n41 VSUBS 0.053383f
C1185 VP.n42 VSUBS 0.037044f
C1186 VP.n43 VSUBS 0.028787f
C1187 VP.n44 VSUBS 0.028787f
C1188 VP.n45 VSUBS 0.043369f
C1189 VP.n46 VSUBS 0.053882f
C1190 VP.n47 VSUBS 0.03425f
C1191 VP.n48 VSUBS 0.028787f
C1192 VP.n49 VSUBS 0.028787f
C1193 VP.n50 VSUBS 0.028787f
C1194 VP.n51 VSUBS 0.053383f
C1195 VP.n52 VSUBS 0.033881f
C1196 VP.n53 VSUBS 1.1235f
C1197 VP.n54 VSUBS 1.83481f
C1198 VP.n55 VSUBS 1.85371f
C1199 VP.n56 VSUBS 1.1235f
C1200 VP.n57 VSUBS 0.033881f
C1201 VP.n58 VSUBS 0.053383f
C1202 VP.n59 VSUBS 0.028787f
C1203 VP.n60 VSUBS 0.028787f
C1204 VP.n61 VSUBS 0.028787f
C1205 VP.n62 VSUBS 0.03425f
C1206 VP.n63 VSUBS 0.053882f
C1207 VP.t2 VSUBS 2.94928f
C1208 VP.n64 VSUBS 1.03284f
C1209 VP.n65 VSUBS 0.043369f
C1210 VP.n66 VSUBS 0.028787f
C1211 VP.n67 VSUBS 0.028787f
C1212 VP.n68 VSUBS 0.028787f
C1213 VP.n69 VSUBS 0.053383f
C1214 VP.n70 VSUBS 0.044236f
C1215 VP.n71 VSUBS 0.039457f
C1216 VP.n72 VSUBS 0.028787f
C1217 VP.n73 VSUBS 0.028787f
C1218 VP.n74 VSUBS 0.028787f
C1219 VP.n75 VSUBS 0.040206f
C1220 VP.n76 VSUBS 1.03284f
C1221 VP.n77 VSUBS 0.040206f
C1222 VP.n78 VSUBS 0.053383f
C1223 VP.n79 VSUBS 0.028787f
C1224 VP.n80 VSUBS 0.028787f
C1225 VP.n81 VSUBS 0.028787f
C1226 VP.n82 VSUBS 0.044236f
C1227 VP.n83 VSUBS 0.053383f
C1228 VP.n84 VSUBS 0.037044f
C1229 VP.n85 VSUBS 0.028787f
C1230 VP.n86 VSUBS 0.028787f
C1231 VP.n87 VSUBS 0.043369f
C1232 VP.n88 VSUBS 0.053882f
C1233 VP.n89 VSUBS 0.03425f
C1234 VP.n90 VSUBS 0.028787f
C1235 VP.n91 VSUBS 0.028787f
C1236 VP.n92 VSUBS 0.028787f
C1237 VP.n93 VSUBS 0.053383f
C1238 VP.n94 VSUBS 0.033881f
C1239 VP.n95 VSUBS 1.1235f
C1240 VP.n96 VSUBS 0.049417f
.ends

