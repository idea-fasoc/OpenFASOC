* NGSPICE file created from diff_pair_sample_0103.ext - technology: sky130A

.subckt diff_pair_sample_0103 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t2 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X1 VDD2.t9 VN.t0 VTAIL.t6 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X2 VDD2.t8 VN.t1 VTAIL.t5 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X3 VDD2.t7 VN.t2 VTAIL.t4 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=2.2308 ps=13.85 w=13.52 l=3.08
X4 VDD2.t6 VN.t3 VTAIL.t19 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=5.2728 ps=27.82 w=13.52 l=3.08
X5 B.t11 B.t9 B.t10 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=3.08
X6 B.t8 B.t6 B.t7 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=3.08
X7 VTAIL.t2 VN.t4 VDD2.t5 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X8 VTAIL.t8 VN.t5 VDD2.t4 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X9 VDD1.t7 VP.t1 VTAIL.t17 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=5.2728 ps=27.82 w=13.52 l=3.08
X10 VTAIL.t16 VP.t2 VDD1.t6 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X11 VTAIL.t0 VN.t6 VDD2.t3 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X12 VDD1.t4 VP.t3 VTAIL.t15 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=2.2308 ps=13.85 w=13.52 l=3.08
X13 VTAIL.t7 VN.t7 VDD2.t2 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X14 VTAIL.t14 VP.t4 VDD1.t3 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X15 VDD1.t9 VP.t5 VTAIL.t13 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=2.2308 ps=13.85 w=13.52 l=3.08
X16 B.t5 B.t3 B.t4 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=3.08
X17 VDD2.t1 VN.t8 VTAIL.t1 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=5.2728 ps=27.82 w=13.52 l=3.08
X18 VTAIL.t12 VP.t6 VDD1.t8 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X19 VDD1.t1 VP.t7 VTAIL.t11 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X20 VDD1.t0 VP.t8 VTAIL.t10 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=2.2308 ps=13.85 w=13.52 l=3.08
X21 VDD1.t5 VP.t9 VTAIL.t9 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=2.2308 pd=13.85 as=5.2728 ps=27.82 w=13.52 l=3.08
X22 B.t2 B.t0 B.t1 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=3.08
X23 VDD2.t0 VN.t9 VTAIL.t3 w_n5062_n3672# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=2.2308 ps=13.85 w=13.52 l=3.08
R0 VP.n29 VP.n28 161.3
R1 VP.n30 VP.n25 161.3
R2 VP.n32 VP.n31 161.3
R3 VP.n33 VP.n24 161.3
R4 VP.n35 VP.n34 161.3
R5 VP.n36 VP.n23 161.3
R6 VP.n38 VP.n37 161.3
R7 VP.n39 VP.n22 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n42 VP.n21 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n45 VP.n20 161.3
R12 VP.n47 VP.n46 161.3
R13 VP.n49 VP.n48 161.3
R14 VP.n50 VP.n18 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n17 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n16 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n94 VP.n93 161.3
R27 VP.n92 VP.n91 161.3
R28 VP.n90 VP.n5 161.3
R29 VP.n89 VP.n88 161.3
R30 VP.n87 VP.n6 161.3
R31 VP.n86 VP.n85 161.3
R32 VP.n84 VP.n7 161.3
R33 VP.n83 VP.n82 161.3
R34 VP.n81 VP.n8 161.3
R35 VP.n80 VP.n79 161.3
R36 VP.n78 VP.n9 161.3
R37 VP.n77 VP.n76 161.3
R38 VP.n75 VP.n10 161.3
R39 VP.n74 VP.n73 161.3
R40 VP.n71 VP.n11 161.3
R41 VP.n70 VP.n69 161.3
R42 VP.n68 VP.n12 161.3
R43 VP.n67 VP.n66 161.3
R44 VP.n65 VP.n13 161.3
R45 VP.n64 VP.n63 161.3
R46 VP.n62 VP.n14 161.3
R47 VP.n26 VP.t3 139.006
R48 VP.n83 VP.t8 105.79
R49 VP.n60 VP.t5 105.79
R50 VP.n72 VP.t4 105.79
R51 VP.n4 VP.t6 105.79
R52 VP.n0 VP.t1 105.79
R53 VP.n38 VP.t7 105.79
R54 VP.n15 VP.t9 105.79
R55 VP.n19 VP.t2 105.79
R56 VP.n27 VP.t0 105.79
R57 VP.n61 VP.n60 74.5068
R58 VP.n104 VP.n0 74.5068
R59 VP.n59 VP.n15 74.5068
R60 VP.n61 VP.n59 56.9503
R61 VP.n78 VP.n77 56.5617
R62 VP.n89 VP.n6 56.5617
R63 VP.n44 VP.n21 56.5617
R64 VP.n33 VP.n32 56.5617
R65 VP.n27 VP.n26 53.9797
R66 VP.n66 VP.n65 51.7179
R67 VP.n100 VP.n2 51.7179
R68 VP.n55 VP.n17 51.7179
R69 VP.n66 VP.n12 29.4362
R70 VP.n96 VP.n2 29.4362
R71 VP.n51 VP.n17 29.4362
R72 VP.n64 VP.n14 24.5923
R73 VP.n65 VP.n64 24.5923
R74 VP.n70 VP.n12 24.5923
R75 VP.n71 VP.n70 24.5923
R76 VP.n73 VP.n10 24.5923
R77 VP.n77 VP.n10 24.5923
R78 VP.n79 VP.n78 24.5923
R79 VP.n79 VP.n8 24.5923
R80 VP.n83 VP.n8 24.5923
R81 VP.n84 VP.n83 24.5923
R82 VP.n85 VP.n84 24.5923
R83 VP.n85 VP.n6 24.5923
R84 VP.n90 VP.n89 24.5923
R85 VP.n91 VP.n90 24.5923
R86 VP.n95 VP.n94 24.5923
R87 VP.n96 VP.n95 24.5923
R88 VP.n101 VP.n100 24.5923
R89 VP.n102 VP.n101 24.5923
R90 VP.n56 VP.n55 24.5923
R91 VP.n57 VP.n56 24.5923
R92 VP.n45 VP.n44 24.5923
R93 VP.n46 VP.n45 24.5923
R94 VP.n50 VP.n49 24.5923
R95 VP.n51 VP.n50 24.5923
R96 VP.n34 VP.n33 24.5923
R97 VP.n34 VP.n23 24.5923
R98 VP.n38 VP.n23 24.5923
R99 VP.n39 VP.n38 24.5923
R100 VP.n40 VP.n39 24.5923
R101 VP.n40 VP.n21 24.5923
R102 VP.n28 VP.n25 24.5923
R103 VP.n32 VP.n25 24.5923
R104 VP.n73 VP.n72 20.1658
R105 VP.n91 VP.n4 20.1658
R106 VP.n46 VP.n19 20.1658
R107 VP.n28 VP.n27 20.1658
R108 VP.n60 VP.n14 15.7393
R109 VP.n102 VP.n0 15.7393
R110 VP.n57 VP.n15 15.7393
R111 VP.n72 VP.n71 4.42703
R112 VP.n94 VP.n4 4.42703
R113 VP.n49 VP.n19 4.42703
R114 VP.n29 VP.n26 4.1008
R115 VP.n59 VP.n58 0.354861
R116 VP.n62 VP.n61 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n30 VP.n29 0.189894
R120 VP.n31 VP.n30 0.189894
R121 VP.n31 VP.n24 0.189894
R122 VP.n35 VP.n24 0.189894
R123 VP.n36 VP.n35 0.189894
R124 VP.n37 VP.n36 0.189894
R125 VP.n37 VP.n22 0.189894
R126 VP.n41 VP.n22 0.189894
R127 VP.n42 VP.n41 0.189894
R128 VP.n43 VP.n42 0.189894
R129 VP.n43 VP.n20 0.189894
R130 VP.n47 VP.n20 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n18 0.189894
R133 VP.n52 VP.n18 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n16 0.189894
R137 VP.n58 VP.n16 0.189894
R138 VP.n63 VP.n62 0.189894
R139 VP.n63 VP.n13 0.189894
R140 VP.n67 VP.n13 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n69 VP.n68 0.189894
R143 VP.n69 VP.n11 0.189894
R144 VP.n74 VP.n11 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n76 VP.n75 0.189894
R147 VP.n76 VP.n9 0.189894
R148 VP.n80 VP.n9 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n82 VP.n81 0.189894
R151 VP.n82 VP.n7 0.189894
R152 VP.n86 VP.n7 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n88 VP.n87 0.189894
R155 VP.n88 VP.n5 0.189894
R156 VP.n92 VP.n5 0.189894
R157 VP.n93 VP.n92 0.189894
R158 VP.n93 VP.n3 0.189894
R159 VP.n97 VP.n3 0.189894
R160 VP.n98 VP.n97 0.189894
R161 VP.n99 VP.n98 0.189894
R162 VP.n99 VP.n1 0.189894
R163 VP.n103 VP.n1 0.189894
R164 VDD1.n68 VDD1.n0 756.745
R165 VDD1.n143 VDD1.n75 756.745
R166 VDD1.n69 VDD1.n68 585
R167 VDD1.n67 VDD1.n66 585
R168 VDD1.n4 VDD1.n3 585
R169 VDD1.n61 VDD1.n60 585
R170 VDD1.n59 VDD1.n58 585
R171 VDD1.n8 VDD1.n7 585
R172 VDD1.n53 VDD1.n52 585
R173 VDD1.n51 VDD1.n50 585
R174 VDD1.n12 VDD1.n11 585
R175 VDD1.n16 VDD1.n14 585
R176 VDD1.n45 VDD1.n44 585
R177 VDD1.n43 VDD1.n42 585
R178 VDD1.n18 VDD1.n17 585
R179 VDD1.n37 VDD1.n36 585
R180 VDD1.n35 VDD1.n34 585
R181 VDD1.n22 VDD1.n21 585
R182 VDD1.n29 VDD1.n28 585
R183 VDD1.n27 VDD1.n26 585
R184 VDD1.n100 VDD1.n99 585
R185 VDD1.n102 VDD1.n101 585
R186 VDD1.n95 VDD1.n94 585
R187 VDD1.n108 VDD1.n107 585
R188 VDD1.n110 VDD1.n109 585
R189 VDD1.n91 VDD1.n90 585
R190 VDD1.n117 VDD1.n116 585
R191 VDD1.n118 VDD1.n89 585
R192 VDD1.n120 VDD1.n119 585
R193 VDD1.n87 VDD1.n86 585
R194 VDD1.n126 VDD1.n125 585
R195 VDD1.n128 VDD1.n127 585
R196 VDD1.n83 VDD1.n82 585
R197 VDD1.n134 VDD1.n133 585
R198 VDD1.n136 VDD1.n135 585
R199 VDD1.n79 VDD1.n78 585
R200 VDD1.n142 VDD1.n141 585
R201 VDD1.n144 VDD1.n143 585
R202 VDD1.n25 VDD1.t4 329.036
R203 VDD1.n98 VDD1.t9 329.036
R204 VDD1.n68 VDD1.n67 171.744
R205 VDD1.n67 VDD1.n3 171.744
R206 VDD1.n60 VDD1.n3 171.744
R207 VDD1.n60 VDD1.n59 171.744
R208 VDD1.n59 VDD1.n7 171.744
R209 VDD1.n52 VDD1.n7 171.744
R210 VDD1.n52 VDD1.n51 171.744
R211 VDD1.n51 VDD1.n11 171.744
R212 VDD1.n16 VDD1.n11 171.744
R213 VDD1.n44 VDD1.n16 171.744
R214 VDD1.n44 VDD1.n43 171.744
R215 VDD1.n43 VDD1.n17 171.744
R216 VDD1.n36 VDD1.n17 171.744
R217 VDD1.n36 VDD1.n35 171.744
R218 VDD1.n35 VDD1.n21 171.744
R219 VDD1.n28 VDD1.n21 171.744
R220 VDD1.n28 VDD1.n27 171.744
R221 VDD1.n101 VDD1.n100 171.744
R222 VDD1.n101 VDD1.n94 171.744
R223 VDD1.n108 VDD1.n94 171.744
R224 VDD1.n109 VDD1.n108 171.744
R225 VDD1.n109 VDD1.n90 171.744
R226 VDD1.n117 VDD1.n90 171.744
R227 VDD1.n118 VDD1.n117 171.744
R228 VDD1.n119 VDD1.n118 171.744
R229 VDD1.n119 VDD1.n86 171.744
R230 VDD1.n126 VDD1.n86 171.744
R231 VDD1.n127 VDD1.n126 171.744
R232 VDD1.n127 VDD1.n82 171.744
R233 VDD1.n134 VDD1.n82 171.744
R234 VDD1.n135 VDD1.n134 171.744
R235 VDD1.n135 VDD1.n78 171.744
R236 VDD1.n142 VDD1.n78 171.744
R237 VDD1.n143 VDD1.n142 171.744
R238 VDD1.n27 VDD1.t4 85.8723
R239 VDD1.n100 VDD1.t9 85.8723
R240 VDD1.n151 VDD1.n150 73.6543
R241 VDD1.n74 VDD1.n73 71.5051
R242 VDD1.n153 VDD1.n152 71.5049
R243 VDD1.n149 VDD1.n148 71.5049
R244 VDD1.n153 VDD1.n151 51.3867
R245 VDD1.n74 VDD1.n72 51.028
R246 VDD1.n149 VDD1.n147 51.028
R247 VDD1.n14 VDD1.n12 13.1884
R248 VDD1.n120 VDD1.n87 13.1884
R249 VDD1.n50 VDD1.n49 12.8005
R250 VDD1.n46 VDD1.n45 12.8005
R251 VDD1.n121 VDD1.n89 12.8005
R252 VDD1.n125 VDD1.n124 12.8005
R253 VDD1.n53 VDD1.n10 12.0247
R254 VDD1.n42 VDD1.n15 12.0247
R255 VDD1.n116 VDD1.n115 12.0247
R256 VDD1.n128 VDD1.n85 12.0247
R257 VDD1.n54 VDD1.n8 11.249
R258 VDD1.n41 VDD1.n18 11.249
R259 VDD1.n114 VDD1.n91 11.249
R260 VDD1.n129 VDD1.n83 11.249
R261 VDD1.n26 VDD1.n25 10.7239
R262 VDD1.n99 VDD1.n98 10.7239
R263 VDD1.n58 VDD1.n57 10.4732
R264 VDD1.n38 VDD1.n37 10.4732
R265 VDD1.n111 VDD1.n110 10.4732
R266 VDD1.n133 VDD1.n132 10.4732
R267 VDD1.n61 VDD1.n6 9.69747
R268 VDD1.n34 VDD1.n20 9.69747
R269 VDD1.n107 VDD1.n93 9.69747
R270 VDD1.n136 VDD1.n81 9.69747
R271 VDD1.n72 VDD1.n71 9.45567
R272 VDD1.n147 VDD1.n146 9.45567
R273 VDD1.n24 VDD1.n23 9.3005
R274 VDD1.n31 VDD1.n30 9.3005
R275 VDD1.n33 VDD1.n32 9.3005
R276 VDD1.n20 VDD1.n19 9.3005
R277 VDD1.n39 VDD1.n38 9.3005
R278 VDD1.n41 VDD1.n40 9.3005
R279 VDD1.n15 VDD1.n13 9.3005
R280 VDD1.n47 VDD1.n46 9.3005
R281 VDD1.n71 VDD1.n70 9.3005
R282 VDD1.n2 VDD1.n1 9.3005
R283 VDD1.n65 VDD1.n64 9.3005
R284 VDD1.n63 VDD1.n62 9.3005
R285 VDD1.n6 VDD1.n5 9.3005
R286 VDD1.n57 VDD1.n56 9.3005
R287 VDD1.n55 VDD1.n54 9.3005
R288 VDD1.n10 VDD1.n9 9.3005
R289 VDD1.n49 VDD1.n48 9.3005
R290 VDD1.n146 VDD1.n145 9.3005
R291 VDD1.n140 VDD1.n139 9.3005
R292 VDD1.n138 VDD1.n137 9.3005
R293 VDD1.n81 VDD1.n80 9.3005
R294 VDD1.n132 VDD1.n131 9.3005
R295 VDD1.n130 VDD1.n129 9.3005
R296 VDD1.n85 VDD1.n84 9.3005
R297 VDD1.n124 VDD1.n123 9.3005
R298 VDD1.n97 VDD1.n96 9.3005
R299 VDD1.n104 VDD1.n103 9.3005
R300 VDD1.n106 VDD1.n105 9.3005
R301 VDD1.n93 VDD1.n92 9.3005
R302 VDD1.n112 VDD1.n111 9.3005
R303 VDD1.n114 VDD1.n113 9.3005
R304 VDD1.n115 VDD1.n88 9.3005
R305 VDD1.n122 VDD1.n121 9.3005
R306 VDD1.n77 VDD1.n76 9.3005
R307 VDD1.n62 VDD1.n4 8.92171
R308 VDD1.n33 VDD1.n22 8.92171
R309 VDD1.n106 VDD1.n95 8.92171
R310 VDD1.n137 VDD1.n79 8.92171
R311 VDD1.n66 VDD1.n65 8.14595
R312 VDD1.n30 VDD1.n29 8.14595
R313 VDD1.n103 VDD1.n102 8.14595
R314 VDD1.n141 VDD1.n140 8.14595
R315 VDD1.n72 VDD1.n0 7.3702
R316 VDD1.n69 VDD1.n2 7.3702
R317 VDD1.n26 VDD1.n24 7.3702
R318 VDD1.n99 VDD1.n97 7.3702
R319 VDD1.n144 VDD1.n77 7.3702
R320 VDD1.n147 VDD1.n75 7.3702
R321 VDD1.n70 VDD1.n0 6.59444
R322 VDD1.n70 VDD1.n69 6.59444
R323 VDD1.n145 VDD1.n144 6.59444
R324 VDD1.n145 VDD1.n75 6.59444
R325 VDD1.n66 VDD1.n2 5.81868
R326 VDD1.n29 VDD1.n24 5.81868
R327 VDD1.n102 VDD1.n97 5.81868
R328 VDD1.n141 VDD1.n77 5.81868
R329 VDD1.n65 VDD1.n4 5.04292
R330 VDD1.n30 VDD1.n22 5.04292
R331 VDD1.n103 VDD1.n95 5.04292
R332 VDD1.n140 VDD1.n79 5.04292
R333 VDD1.n62 VDD1.n61 4.26717
R334 VDD1.n34 VDD1.n33 4.26717
R335 VDD1.n107 VDD1.n106 4.26717
R336 VDD1.n137 VDD1.n136 4.26717
R337 VDD1.n58 VDD1.n6 3.49141
R338 VDD1.n37 VDD1.n20 3.49141
R339 VDD1.n110 VDD1.n93 3.49141
R340 VDD1.n133 VDD1.n81 3.49141
R341 VDD1.n57 VDD1.n8 2.71565
R342 VDD1.n38 VDD1.n18 2.71565
R343 VDD1.n111 VDD1.n91 2.71565
R344 VDD1.n132 VDD1.n83 2.71565
R345 VDD1.n25 VDD1.n23 2.41282
R346 VDD1.n98 VDD1.n96 2.41282
R347 VDD1.n152 VDD1.t6 2.40472
R348 VDD1.n152 VDD1.t5 2.40472
R349 VDD1.n73 VDD1.t2 2.40472
R350 VDD1.n73 VDD1.t1 2.40472
R351 VDD1.n150 VDD1.t8 2.40472
R352 VDD1.n150 VDD1.t7 2.40472
R353 VDD1.n148 VDD1.t3 2.40472
R354 VDD1.n148 VDD1.t0 2.40472
R355 VDD1 VDD1.n153 2.14705
R356 VDD1.n54 VDD1.n53 1.93989
R357 VDD1.n42 VDD1.n41 1.93989
R358 VDD1.n116 VDD1.n114 1.93989
R359 VDD1.n129 VDD1.n128 1.93989
R360 VDD1.n50 VDD1.n10 1.16414
R361 VDD1.n45 VDD1.n15 1.16414
R362 VDD1.n115 VDD1.n89 1.16414
R363 VDD1.n125 VDD1.n85 1.16414
R364 VDD1 VDD1.n74 0.793603
R365 VDD1.n151 VDD1.n149 0.680068
R366 VDD1.n49 VDD1.n12 0.388379
R367 VDD1.n46 VDD1.n14 0.388379
R368 VDD1.n121 VDD1.n120 0.388379
R369 VDD1.n124 VDD1.n87 0.388379
R370 VDD1.n71 VDD1.n1 0.155672
R371 VDD1.n64 VDD1.n1 0.155672
R372 VDD1.n64 VDD1.n63 0.155672
R373 VDD1.n63 VDD1.n5 0.155672
R374 VDD1.n56 VDD1.n5 0.155672
R375 VDD1.n56 VDD1.n55 0.155672
R376 VDD1.n55 VDD1.n9 0.155672
R377 VDD1.n48 VDD1.n9 0.155672
R378 VDD1.n48 VDD1.n47 0.155672
R379 VDD1.n47 VDD1.n13 0.155672
R380 VDD1.n40 VDD1.n13 0.155672
R381 VDD1.n40 VDD1.n39 0.155672
R382 VDD1.n39 VDD1.n19 0.155672
R383 VDD1.n32 VDD1.n19 0.155672
R384 VDD1.n32 VDD1.n31 0.155672
R385 VDD1.n31 VDD1.n23 0.155672
R386 VDD1.n104 VDD1.n96 0.155672
R387 VDD1.n105 VDD1.n104 0.155672
R388 VDD1.n105 VDD1.n92 0.155672
R389 VDD1.n112 VDD1.n92 0.155672
R390 VDD1.n113 VDD1.n112 0.155672
R391 VDD1.n113 VDD1.n88 0.155672
R392 VDD1.n122 VDD1.n88 0.155672
R393 VDD1.n123 VDD1.n122 0.155672
R394 VDD1.n123 VDD1.n84 0.155672
R395 VDD1.n130 VDD1.n84 0.155672
R396 VDD1.n131 VDD1.n130 0.155672
R397 VDD1.n131 VDD1.n80 0.155672
R398 VDD1.n138 VDD1.n80 0.155672
R399 VDD1.n139 VDD1.n138 0.155672
R400 VDD1.n139 VDD1.n76 0.155672
R401 VDD1.n146 VDD1.n76 0.155672
R402 VTAIL.n304 VTAIL.n236 756.745
R403 VTAIL.n70 VTAIL.n2 756.745
R404 VTAIL.n230 VTAIL.n162 756.745
R405 VTAIL.n152 VTAIL.n84 756.745
R406 VTAIL.n261 VTAIL.n260 585
R407 VTAIL.n263 VTAIL.n262 585
R408 VTAIL.n256 VTAIL.n255 585
R409 VTAIL.n269 VTAIL.n268 585
R410 VTAIL.n271 VTAIL.n270 585
R411 VTAIL.n252 VTAIL.n251 585
R412 VTAIL.n278 VTAIL.n277 585
R413 VTAIL.n279 VTAIL.n250 585
R414 VTAIL.n281 VTAIL.n280 585
R415 VTAIL.n248 VTAIL.n247 585
R416 VTAIL.n287 VTAIL.n286 585
R417 VTAIL.n289 VTAIL.n288 585
R418 VTAIL.n244 VTAIL.n243 585
R419 VTAIL.n295 VTAIL.n294 585
R420 VTAIL.n297 VTAIL.n296 585
R421 VTAIL.n240 VTAIL.n239 585
R422 VTAIL.n303 VTAIL.n302 585
R423 VTAIL.n305 VTAIL.n304 585
R424 VTAIL.n27 VTAIL.n26 585
R425 VTAIL.n29 VTAIL.n28 585
R426 VTAIL.n22 VTAIL.n21 585
R427 VTAIL.n35 VTAIL.n34 585
R428 VTAIL.n37 VTAIL.n36 585
R429 VTAIL.n18 VTAIL.n17 585
R430 VTAIL.n44 VTAIL.n43 585
R431 VTAIL.n45 VTAIL.n16 585
R432 VTAIL.n47 VTAIL.n46 585
R433 VTAIL.n14 VTAIL.n13 585
R434 VTAIL.n53 VTAIL.n52 585
R435 VTAIL.n55 VTAIL.n54 585
R436 VTAIL.n10 VTAIL.n9 585
R437 VTAIL.n61 VTAIL.n60 585
R438 VTAIL.n63 VTAIL.n62 585
R439 VTAIL.n6 VTAIL.n5 585
R440 VTAIL.n69 VTAIL.n68 585
R441 VTAIL.n71 VTAIL.n70 585
R442 VTAIL.n231 VTAIL.n230 585
R443 VTAIL.n229 VTAIL.n228 585
R444 VTAIL.n166 VTAIL.n165 585
R445 VTAIL.n223 VTAIL.n222 585
R446 VTAIL.n221 VTAIL.n220 585
R447 VTAIL.n170 VTAIL.n169 585
R448 VTAIL.n215 VTAIL.n214 585
R449 VTAIL.n213 VTAIL.n212 585
R450 VTAIL.n174 VTAIL.n173 585
R451 VTAIL.n178 VTAIL.n176 585
R452 VTAIL.n207 VTAIL.n206 585
R453 VTAIL.n205 VTAIL.n204 585
R454 VTAIL.n180 VTAIL.n179 585
R455 VTAIL.n199 VTAIL.n198 585
R456 VTAIL.n197 VTAIL.n196 585
R457 VTAIL.n184 VTAIL.n183 585
R458 VTAIL.n191 VTAIL.n190 585
R459 VTAIL.n189 VTAIL.n188 585
R460 VTAIL.n153 VTAIL.n152 585
R461 VTAIL.n151 VTAIL.n150 585
R462 VTAIL.n88 VTAIL.n87 585
R463 VTAIL.n145 VTAIL.n144 585
R464 VTAIL.n143 VTAIL.n142 585
R465 VTAIL.n92 VTAIL.n91 585
R466 VTAIL.n137 VTAIL.n136 585
R467 VTAIL.n135 VTAIL.n134 585
R468 VTAIL.n96 VTAIL.n95 585
R469 VTAIL.n100 VTAIL.n98 585
R470 VTAIL.n129 VTAIL.n128 585
R471 VTAIL.n127 VTAIL.n126 585
R472 VTAIL.n102 VTAIL.n101 585
R473 VTAIL.n121 VTAIL.n120 585
R474 VTAIL.n119 VTAIL.n118 585
R475 VTAIL.n106 VTAIL.n105 585
R476 VTAIL.n113 VTAIL.n112 585
R477 VTAIL.n111 VTAIL.n110 585
R478 VTAIL.n259 VTAIL.t19 329.036
R479 VTAIL.n25 VTAIL.t17 329.036
R480 VTAIL.n187 VTAIL.t9 329.036
R481 VTAIL.n109 VTAIL.t1 329.036
R482 VTAIL.n262 VTAIL.n261 171.744
R483 VTAIL.n262 VTAIL.n255 171.744
R484 VTAIL.n269 VTAIL.n255 171.744
R485 VTAIL.n270 VTAIL.n269 171.744
R486 VTAIL.n270 VTAIL.n251 171.744
R487 VTAIL.n278 VTAIL.n251 171.744
R488 VTAIL.n279 VTAIL.n278 171.744
R489 VTAIL.n280 VTAIL.n279 171.744
R490 VTAIL.n280 VTAIL.n247 171.744
R491 VTAIL.n287 VTAIL.n247 171.744
R492 VTAIL.n288 VTAIL.n287 171.744
R493 VTAIL.n288 VTAIL.n243 171.744
R494 VTAIL.n295 VTAIL.n243 171.744
R495 VTAIL.n296 VTAIL.n295 171.744
R496 VTAIL.n296 VTAIL.n239 171.744
R497 VTAIL.n303 VTAIL.n239 171.744
R498 VTAIL.n304 VTAIL.n303 171.744
R499 VTAIL.n28 VTAIL.n27 171.744
R500 VTAIL.n28 VTAIL.n21 171.744
R501 VTAIL.n35 VTAIL.n21 171.744
R502 VTAIL.n36 VTAIL.n35 171.744
R503 VTAIL.n36 VTAIL.n17 171.744
R504 VTAIL.n44 VTAIL.n17 171.744
R505 VTAIL.n45 VTAIL.n44 171.744
R506 VTAIL.n46 VTAIL.n45 171.744
R507 VTAIL.n46 VTAIL.n13 171.744
R508 VTAIL.n53 VTAIL.n13 171.744
R509 VTAIL.n54 VTAIL.n53 171.744
R510 VTAIL.n54 VTAIL.n9 171.744
R511 VTAIL.n61 VTAIL.n9 171.744
R512 VTAIL.n62 VTAIL.n61 171.744
R513 VTAIL.n62 VTAIL.n5 171.744
R514 VTAIL.n69 VTAIL.n5 171.744
R515 VTAIL.n70 VTAIL.n69 171.744
R516 VTAIL.n230 VTAIL.n229 171.744
R517 VTAIL.n229 VTAIL.n165 171.744
R518 VTAIL.n222 VTAIL.n165 171.744
R519 VTAIL.n222 VTAIL.n221 171.744
R520 VTAIL.n221 VTAIL.n169 171.744
R521 VTAIL.n214 VTAIL.n169 171.744
R522 VTAIL.n214 VTAIL.n213 171.744
R523 VTAIL.n213 VTAIL.n173 171.744
R524 VTAIL.n178 VTAIL.n173 171.744
R525 VTAIL.n206 VTAIL.n178 171.744
R526 VTAIL.n206 VTAIL.n205 171.744
R527 VTAIL.n205 VTAIL.n179 171.744
R528 VTAIL.n198 VTAIL.n179 171.744
R529 VTAIL.n198 VTAIL.n197 171.744
R530 VTAIL.n197 VTAIL.n183 171.744
R531 VTAIL.n190 VTAIL.n183 171.744
R532 VTAIL.n190 VTAIL.n189 171.744
R533 VTAIL.n152 VTAIL.n151 171.744
R534 VTAIL.n151 VTAIL.n87 171.744
R535 VTAIL.n144 VTAIL.n87 171.744
R536 VTAIL.n144 VTAIL.n143 171.744
R537 VTAIL.n143 VTAIL.n91 171.744
R538 VTAIL.n136 VTAIL.n91 171.744
R539 VTAIL.n136 VTAIL.n135 171.744
R540 VTAIL.n135 VTAIL.n95 171.744
R541 VTAIL.n100 VTAIL.n95 171.744
R542 VTAIL.n128 VTAIL.n100 171.744
R543 VTAIL.n128 VTAIL.n127 171.744
R544 VTAIL.n127 VTAIL.n101 171.744
R545 VTAIL.n120 VTAIL.n101 171.744
R546 VTAIL.n120 VTAIL.n119 171.744
R547 VTAIL.n119 VTAIL.n105 171.744
R548 VTAIL.n112 VTAIL.n105 171.744
R549 VTAIL.n112 VTAIL.n111 171.744
R550 VTAIL.n261 VTAIL.t19 85.8723
R551 VTAIL.n27 VTAIL.t17 85.8723
R552 VTAIL.n189 VTAIL.t9 85.8723
R553 VTAIL.n111 VTAIL.t1 85.8723
R554 VTAIL.n161 VTAIL.n160 54.8263
R555 VTAIL.n159 VTAIL.n158 54.8263
R556 VTAIL.n83 VTAIL.n82 54.8263
R557 VTAIL.n81 VTAIL.n80 54.8263
R558 VTAIL.n311 VTAIL.n310 54.8261
R559 VTAIL.n1 VTAIL.n0 54.8261
R560 VTAIL.n77 VTAIL.n76 54.8261
R561 VTAIL.n79 VTAIL.n78 54.8261
R562 VTAIL.n309 VTAIL.n308 31.4096
R563 VTAIL.n75 VTAIL.n74 31.4096
R564 VTAIL.n235 VTAIL.n234 31.4096
R565 VTAIL.n157 VTAIL.n156 31.4096
R566 VTAIL.n81 VTAIL.n79 29.9014
R567 VTAIL.n309 VTAIL.n235 26.9617
R568 VTAIL.n281 VTAIL.n248 13.1884
R569 VTAIL.n47 VTAIL.n14 13.1884
R570 VTAIL.n176 VTAIL.n174 13.1884
R571 VTAIL.n98 VTAIL.n96 13.1884
R572 VTAIL.n282 VTAIL.n250 12.8005
R573 VTAIL.n286 VTAIL.n285 12.8005
R574 VTAIL.n48 VTAIL.n16 12.8005
R575 VTAIL.n52 VTAIL.n51 12.8005
R576 VTAIL.n212 VTAIL.n211 12.8005
R577 VTAIL.n208 VTAIL.n207 12.8005
R578 VTAIL.n134 VTAIL.n133 12.8005
R579 VTAIL.n130 VTAIL.n129 12.8005
R580 VTAIL.n277 VTAIL.n276 12.0247
R581 VTAIL.n289 VTAIL.n246 12.0247
R582 VTAIL.n43 VTAIL.n42 12.0247
R583 VTAIL.n55 VTAIL.n12 12.0247
R584 VTAIL.n215 VTAIL.n172 12.0247
R585 VTAIL.n204 VTAIL.n177 12.0247
R586 VTAIL.n137 VTAIL.n94 12.0247
R587 VTAIL.n126 VTAIL.n99 12.0247
R588 VTAIL.n275 VTAIL.n252 11.249
R589 VTAIL.n290 VTAIL.n244 11.249
R590 VTAIL.n41 VTAIL.n18 11.249
R591 VTAIL.n56 VTAIL.n10 11.249
R592 VTAIL.n216 VTAIL.n170 11.249
R593 VTAIL.n203 VTAIL.n180 11.249
R594 VTAIL.n138 VTAIL.n92 11.249
R595 VTAIL.n125 VTAIL.n102 11.249
R596 VTAIL.n260 VTAIL.n259 10.7239
R597 VTAIL.n26 VTAIL.n25 10.7239
R598 VTAIL.n188 VTAIL.n187 10.7239
R599 VTAIL.n110 VTAIL.n109 10.7239
R600 VTAIL.n272 VTAIL.n271 10.4732
R601 VTAIL.n294 VTAIL.n293 10.4732
R602 VTAIL.n38 VTAIL.n37 10.4732
R603 VTAIL.n60 VTAIL.n59 10.4732
R604 VTAIL.n220 VTAIL.n219 10.4732
R605 VTAIL.n200 VTAIL.n199 10.4732
R606 VTAIL.n142 VTAIL.n141 10.4732
R607 VTAIL.n122 VTAIL.n121 10.4732
R608 VTAIL.n268 VTAIL.n254 9.69747
R609 VTAIL.n297 VTAIL.n242 9.69747
R610 VTAIL.n34 VTAIL.n20 9.69747
R611 VTAIL.n63 VTAIL.n8 9.69747
R612 VTAIL.n223 VTAIL.n168 9.69747
R613 VTAIL.n196 VTAIL.n182 9.69747
R614 VTAIL.n145 VTAIL.n90 9.69747
R615 VTAIL.n118 VTAIL.n104 9.69747
R616 VTAIL.n308 VTAIL.n307 9.45567
R617 VTAIL.n74 VTAIL.n73 9.45567
R618 VTAIL.n234 VTAIL.n233 9.45567
R619 VTAIL.n156 VTAIL.n155 9.45567
R620 VTAIL.n307 VTAIL.n306 9.3005
R621 VTAIL.n301 VTAIL.n300 9.3005
R622 VTAIL.n299 VTAIL.n298 9.3005
R623 VTAIL.n242 VTAIL.n241 9.3005
R624 VTAIL.n293 VTAIL.n292 9.3005
R625 VTAIL.n291 VTAIL.n290 9.3005
R626 VTAIL.n246 VTAIL.n245 9.3005
R627 VTAIL.n285 VTAIL.n284 9.3005
R628 VTAIL.n258 VTAIL.n257 9.3005
R629 VTAIL.n265 VTAIL.n264 9.3005
R630 VTAIL.n267 VTAIL.n266 9.3005
R631 VTAIL.n254 VTAIL.n253 9.3005
R632 VTAIL.n273 VTAIL.n272 9.3005
R633 VTAIL.n275 VTAIL.n274 9.3005
R634 VTAIL.n276 VTAIL.n249 9.3005
R635 VTAIL.n283 VTAIL.n282 9.3005
R636 VTAIL.n238 VTAIL.n237 9.3005
R637 VTAIL.n73 VTAIL.n72 9.3005
R638 VTAIL.n67 VTAIL.n66 9.3005
R639 VTAIL.n65 VTAIL.n64 9.3005
R640 VTAIL.n8 VTAIL.n7 9.3005
R641 VTAIL.n59 VTAIL.n58 9.3005
R642 VTAIL.n57 VTAIL.n56 9.3005
R643 VTAIL.n12 VTAIL.n11 9.3005
R644 VTAIL.n51 VTAIL.n50 9.3005
R645 VTAIL.n24 VTAIL.n23 9.3005
R646 VTAIL.n31 VTAIL.n30 9.3005
R647 VTAIL.n33 VTAIL.n32 9.3005
R648 VTAIL.n20 VTAIL.n19 9.3005
R649 VTAIL.n39 VTAIL.n38 9.3005
R650 VTAIL.n41 VTAIL.n40 9.3005
R651 VTAIL.n42 VTAIL.n15 9.3005
R652 VTAIL.n49 VTAIL.n48 9.3005
R653 VTAIL.n4 VTAIL.n3 9.3005
R654 VTAIL.n186 VTAIL.n185 9.3005
R655 VTAIL.n193 VTAIL.n192 9.3005
R656 VTAIL.n195 VTAIL.n194 9.3005
R657 VTAIL.n182 VTAIL.n181 9.3005
R658 VTAIL.n201 VTAIL.n200 9.3005
R659 VTAIL.n203 VTAIL.n202 9.3005
R660 VTAIL.n177 VTAIL.n175 9.3005
R661 VTAIL.n209 VTAIL.n208 9.3005
R662 VTAIL.n233 VTAIL.n232 9.3005
R663 VTAIL.n164 VTAIL.n163 9.3005
R664 VTAIL.n227 VTAIL.n226 9.3005
R665 VTAIL.n225 VTAIL.n224 9.3005
R666 VTAIL.n168 VTAIL.n167 9.3005
R667 VTAIL.n219 VTAIL.n218 9.3005
R668 VTAIL.n217 VTAIL.n216 9.3005
R669 VTAIL.n172 VTAIL.n171 9.3005
R670 VTAIL.n211 VTAIL.n210 9.3005
R671 VTAIL.n108 VTAIL.n107 9.3005
R672 VTAIL.n115 VTAIL.n114 9.3005
R673 VTAIL.n117 VTAIL.n116 9.3005
R674 VTAIL.n104 VTAIL.n103 9.3005
R675 VTAIL.n123 VTAIL.n122 9.3005
R676 VTAIL.n125 VTAIL.n124 9.3005
R677 VTAIL.n99 VTAIL.n97 9.3005
R678 VTAIL.n131 VTAIL.n130 9.3005
R679 VTAIL.n155 VTAIL.n154 9.3005
R680 VTAIL.n86 VTAIL.n85 9.3005
R681 VTAIL.n149 VTAIL.n148 9.3005
R682 VTAIL.n147 VTAIL.n146 9.3005
R683 VTAIL.n90 VTAIL.n89 9.3005
R684 VTAIL.n141 VTAIL.n140 9.3005
R685 VTAIL.n139 VTAIL.n138 9.3005
R686 VTAIL.n94 VTAIL.n93 9.3005
R687 VTAIL.n133 VTAIL.n132 9.3005
R688 VTAIL.n267 VTAIL.n256 8.92171
R689 VTAIL.n298 VTAIL.n240 8.92171
R690 VTAIL.n33 VTAIL.n22 8.92171
R691 VTAIL.n64 VTAIL.n6 8.92171
R692 VTAIL.n224 VTAIL.n166 8.92171
R693 VTAIL.n195 VTAIL.n184 8.92171
R694 VTAIL.n146 VTAIL.n88 8.92171
R695 VTAIL.n117 VTAIL.n106 8.92171
R696 VTAIL.n264 VTAIL.n263 8.14595
R697 VTAIL.n302 VTAIL.n301 8.14595
R698 VTAIL.n30 VTAIL.n29 8.14595
R699 VTAIL.n68 VTAIL.n67 8.14595
R700 VTAIL.n228 VTAIL.n227 8.14595
R701 VTAIL.n192 VTAIL.n191 8.14595
R702 VTAIL.n150 VTAIL.n149 8.14595
R703 VTAIL.n114 VTAIL.n113 8.14595
R704 VTAIL.n260 VTAIL.n258 7.3702
R705 VTAIL.n305 VTAIL.n238 7.3702
R706 VTAIL.n308 VTAIL.n236 7.3702
R707 VTAIL.n26 VTAIL.n24 7.3702
R708 VTAIL.n71 VTAIL.n4 7.3702
R709 VTAIL.n74 VTAIL.n2 7.3702
R710 VTAIL.n234 VTAIL.n162 7.3702
R711 VTAIL.n231 VTAIL.n164 7.3702
R712 VTAIL.n188 VTAIL.n186 7.3702
R713 VTAIL.n156 VTAIL.n84 7.3702
R714 VTAIL.n153 VTAIL.n86 7.3702
R715 VTAIL.n110 VTAIL.n108 7.3702
R716 VTAIL.n306 VTAIL.n305 6.59444
R717 VTAIL.n306 VTAIL.n236 6.59444
R718 VTAIL.n72 VTAIL.n71 6.59444
R719 VTAIL.n72 VTAIL.n2 6.59444
R720 VTAIL.n232 VTAIL.n162 6.59444
R721 VTAIL.n232 VTAIL.n231 6.59444
R722 VTAIL.n154 VTAIL.n84 6.59444
R723 VTAIL.n154 VTAIL.n153 6.59444
R724 VTAIL.n263 VTAIL.n258 5.81868
R725 VTAIL.n302 VTAIL.n238 5.81868
R726 VTAIL.n29 VTAIL.n24 5.81868
R727 VTAIL.n68 VTAIL.n4 5.81868
R728 VTAIL.n228 VTAIL.n164 5.81868
R729 VTAIL.n191 VTAIL.n186 5.81868
R730 VTAIL.n150 VTAIL.n86 5.81868
R731 VTAIL.n113 VTAIL.n108 5.81868
R732 VTAIL.n264 VTAIL.n256 5.04292
R733 VTAIL.n301 VTAIL.n240 5.04292
R734 VTAIL.n30 VTAIL.n22 5.04292
R735 VTAIL.n67 VTAIL.n6 5.04292
R736 VTAIL.n227 VTAIL.n166 5.04292
R737 VTAIL.n192 VTAIL.n184 5.04292
R738 VTAIL.n149 VTAIL.n88 5.04292
R739 VTAIL.n114 VTAIL.n106 5.04292
R740 VTAIL.n268 VTAIL.n267 4.26717
R741 VTAIL.n298 VTAIL.n297 4.26717
R742 VTAIL.n34 VTAIL.n33 4.26717
R743 VTAIL.n64 VTAIL.n63 4.26717
R744 VTAIL.n224 VTAIL.n223 4.26717
R745 VTAIL.n196 VTAIL.n195 4.26717
R746 VTAIL.n146 VTAIL.n145 4.26717
R747 VTAIL.n118 VTAIL.n117 4.26717
R748 VTAIL.n271 VTAIL.n254 3.49141
R749 VTAIL.n294 VTAIL.n242 3.49141
R750 VTAIL.n37 VTAIL.n20 3.49141
R751 VTAIL.n60 VTAIL.n8 3.49141
R752 VTAIL.n220 VTAIL.n168 3.49141
R753 VTAIL.n199 VTAIL.n182 3.49141
R754 VTAIL.n142 VTAIL.n90 3.49141
R755 VTAIL.n121 VTAIL.n104 3.49141
R756 VTAIL.n83 VTAIL.n81 2.94016
R757 VTAIL.n157 VTAIL.n83 2.94016
R758 VTAIL.n161 VTAIL.n159 2.94016
R759 VTAIL.n235 VTAIL.n161 2.94016
R760 VTAIL.n79 VTAIL.n77 2.94016
R761 VTAIL.n77 VTAIL.n75 2.94016
R762 VTAIL.n311 VTAIL.n309 2.94016
R763 VTAIL.n272 VTAIL.n252 2.71565
R764 VTAIL.n293 VTAIL.n244 2.71565
R765 VTAIL.n38 VTAIL.n18 2.71565
R766 VTAIL.n59 VTAIL.n10 2.71565
R767 VTAIL.n219 VTAIL.n170 2.71565
R768 VTAIL.n200 VTAIL.n180 2.71565
R769 VTAIL.n141 VTAIL.n92 2.71565
R770 VTAIL.n122 VTAIL.n102 2.71565
R771 VTAIL.n259 VTAIL.n257 2.41282
R772 VTAIL.n25 VTAIL.n23 2.41282
R773 VTAIL.n187 VTAIL.n185 2.41282
R774 VTAIL.n109 VTAIL.n107 2.41282
R775 VTAIL.n310 VTAIL.t6 2.40472
R776 VTAIL.n310 VTAIL.t0 2.40472
R777 VTAIL.n0 VTAIL.t3 2.40472
R778 VTAIL.n0 VTAIL.t2 2.40472
R779 VTAIL.n76 VTAIL.t10 2.40472
R780 VTAIL.n76 VTAIL.t12 2.40472
R781 VTAIL.n78 VTAIL.t13 2.40472
R782 VTAIL.n78 VTAIL.t14 2.40472
R783 VTAIL.n160 VTAIL.t11 2.40472
R784 VTAIL.n160 VTAIL.t16 2.40472
R785 VTAIL.n158 VTAIL.t15 2.40472
R786 VTAIL.n158 VTAIL.t18 2.40472
R787 VTAIL.n82 VTAIL.t5 2.40472
R788 VTAIL.n82 VTAIL.t8 2.40472
R789 VTAIL.n80 VTAIL.t4 2.40472
R790 VTAIL.n80 VTAIL.t7 2.40472
R791 VTAIL VTAIL.n1 2.26343
R792 VTAIL.n159 VTAIL.n157 1.94016
R793 VTAIL.n75 VTAIL.n1 1.94016
R794 VTAIL.n277 VTAIL.n275 1.93989
R795 VTAIL.n290 VTAIL.n289 1.93989
R796 VTAIL.n43 VTAIL.n41 1.93989
R797 VTAIL.n56 VTAIL.n55 1.93989
R798 VTAIL.n216 VTAIL.n215 1.93989
R799 VTAIL.n204 VTAIL.n203 1.93989
R800 VTAIL.n138 VTAIL.n137 1.93989
R801 VTAIL.n126 VTAIL.n125 1.93989
R802 VTAIL.n276 VTAIL.n250 1.16414
R803 VTAIL.n286 VTAIL.n246 1.16414
R804 VTAIL.n42 VTAIL.n16 1.16414
R805 VTAIL.n52 VTAIL.n12 1.16414
R806 VTAIL.n212 VTAIL.n172 1.16414
R807 VTAIL.n207 VTAIL.n177 1.16414
R808 VTAIL.n134 VTAIL.n94 1.16414
R809 VTAIL.n129 VTAIL.n99 1.16414
R810 VTAIL VTAIL.n311 0.677224
R811 VTAIL.n282 VTAIL.n281 0.388379
R812 VTAIL.n285 VTAIL.n248 0.388379
R813 VTAIL.n48 VTAIL.n47 0.388379
R814 VTAIL.n51 VTAIL.n14 0.388379
R815 VTAIL.n211 VTAIL.n174 0.388379
R816 VTAIL.n208 VTAIL.n176 0.388379
R817 VTAIL.n133 VTAIL.n96 0.388379
R818 VTAIL.n130 VTAIL.n98 0.388379
R819 VTAIL.n265 VTAIL.n257 0.155672
R820 VTAIL.n266 VTAIL.n265 0.155672
R821 VTAIL.n266 VTAIL.n253 0.155672
R822 VTAIL.n273 VTAIL.n253 0.155672
R823 VTAIL.n274 VTAIL.n273 0.155672
R824 VTAIL.n274 VTAIL.n249 0.155672
R825 VTAIL.n283 VTAIL.n249 0.155672
R826 VTAIL.n284 VTAIL.n283 0.155672
R827 VTAIL.n284 VTAIL.n245 0.155672
R828 VTAIL.n291 VTAIL.n245 0.155672
R829 VTAIL.n292 VTAIL.n291 0.155672
R830 VTAIL.n292 VTAIL.n241 0.155672
R831 VTAIL.n299 VTAIL.n241 0.155672
R832 VTAIL.n300 VTAIL.n299 0.155672
R833 VTAIL.n300 VTAIL.n237 0.155672
R834 VTAIL.n307 VTAIL.n237 0.155672
R835 VTAIL.n31 VTAIL.n23 0.155672
R836 VTAIL.n32 VTAIL.n31 0.155672
R837 VTAIL.n32 VTAIL.n19 0.155672
R838 VTAIL.n39 VTAIL.n19 0.155672
R839 VTAIL.n40 VTAIL.n39 0.155672
R840 VTAIL.n40 VTAIL.n15 0.155672
R841 VTAIL.n49 VTAIL.n15 0.155672
R842 VTAIL.n50 VTAIL.n49 0.155672
R843 VTAIL.n50 VTAIL.n11 0.155672
R844 VTAIL.n57 VTAIL.n11 0.155672
R845 VTAIL.n58 VTAIL.n57 0.155672
R846 VTAIL.n58 VTAIL.n7 0.155672
R847 VTAIL.n65 VTAIL.n7 0.155672
R848 VTAIL.n66 VTAIL.n65 0.155672
R849 VTAIL.n66 VTAIL.n3 0.155672
R850 VTAIL.n73 VTAIL.n3 0.155672
R851 VTAIL.n233 VTAIL.n163 0.155672
R852 VTAIL.n226 VTAIL.n163 0.155672
R853 VTAIL.n226 VTAIL.n225 0.155672
R854 VTAIL.n225 VTAIL.n167 0.155672
R855 VTAIL.n218 VTAIL.n167 0.155672
R856 VTAIL.n218 VTAIL.n217 0.155672
R857 VTAIL.n217 VTAIL.n171 0.155672
R858 VTAIL.n210 VTAIL.n171 0.155672
R859 VTAIL.n210 VTAIL.n209 0.155672
R860 VTAIL.n209 VTAIL.n175 0.155672
R861 VTAIL.n202 VTAIL.n175 0.155672
R862 VTAIL.n202 VTAIL.n201 0.155672
R863 VTAIL.n201 VTAIL.n181 0.155672
R864 VTAIL.n194 VTAIL.n181 0.155672
R865 VTAIL.n194 VTAIL.n193 0.155672
R866 VTAIL.n193 VTAIL.n185 0.155672
R867 VTAIL.n155 VTAIL.n85 0.155672
R868 VTAIL.n148 VTAIL.n85 0.155672
R869 VTAIL.n148 VTAIL.n147 0.155672
R870 VTAIL.n147 VTAIL.n89 0.155672
R871 VTAIL.n140 VTAIL.n89 0.155672
R872 VTAIL.n140 VTAIL.n139 0.155672
R873 VTAIL.n139 VTAIL.n93 0.155672
R874 VTAIL.n132 VTAIL.n93 0.155672
R875 VTAIL.n132 VTAIL.n131 0.155672
R876 VTAIL.n131 VTAIL.n97 0.155672
R877 VTAIL.n124 VTAIL.n97 0.155672
R878 VTAIL.n124 VTAIL.n123 0.155672
R879 VTAIL.n123 VTAIL.n103 0.155672
R880 VTAIL.n116 VTAIL.n103 0.155672
R881 VTAIL.n116 VTAIL.n115 0.155672
R882 VTAIL.n115 VTAIL.n107 0.155672
R883 VN.n88 VN.n87 161.3
R884 VN.n86 VN.n46 161.3
R885 VN.n85 VN.n84 161.3
R886 VN.n83 VN.n47 161.3
R887 VN.n82 VN.n81 161.3
R888 VN.n80 VN.n48 161.3
R889 VN.n79 VN.n78 161.3
R890 VN.n77 VN.n76 161.3
R891 VN.n75 VN.n50 161.3
R892 VN.n74 VN.n73 161.3
R893 VN.n72 VN.n51 161.3
R894 VN.n71 VN.n70 161.3
R895 VN.n69 VN.n52 161.3
R896 VN.n68 VN.n67 161.3
R897 VN.n66 VN.n53 161.3
R898 VN.n65 VN.n64 161.3
R899 VN.n63 VN.n54 161.3
R900 VN.n62 VN.n61 161.3
R901 VN.n60 VN.n55 161.3
R902 VN.n59 VN.n58 161.3
R903 VN.n43 VN.n42 161.3
R904 VN.n41 VN.n1 161.3
R905 VN.n40 VN.n39 161.3
R906 VN.n38 VN.n2 161.3
R907 VN.n37 VN.n36 161.3
R908 VN.n35 VN.n3 161.3
R909 VN.n34 VN.n33 161.3
R910 VN.n32 VN.n31 161.3
R911 VN.n30 VN.n5 161.3
R912 VN.n29 VN.n28 161.3
R913 VN.n27 VN.n6 161.3
R914 VN.n26 VN.n25 161.3
R915 VN.n24 VN.n7 161.3
R916 VN.n23 VN.n22 161.3
R917 VN.n21 VN.n8 161.3
R918 VN.n20 VN.n19 161.3
R919 VN.n18 VN.n9 161.3
R920 VN.n17 VN.n16 161.3
R921 VN.n15 VN.n10 161.3
R922 VN.n14 VN.n13 161.3
R923 VN.n56 VN.t8 139.006
R924 VN.n11 VN.t9 139.006
R925 VN.n23 VN.t0 105.79
R926 VN.n12 VN.t4 105.79
R927 VN.n4 VN.t6 105.79
R928 VN.n0 VN.t3 105.79
R929 VN.n68 VN.t1 105.79
R930 VN.n57 VN.t5 105.79
R931 VN.n49 VN.t7 105.79
R932 VN.n45 VN.t2 105.79
R933 VN.n44 VN.n0 74.5068
R934 VN.n89 VN.n45 74.5068
R935 VN VN.n89 57.1156
R936 VN.n18 VN.n17 56.5617
R937 VN.n29 VN.n6 56.5617
R938 VN.n63 VN.n62 56.5617
R939 VN.n74 VN.n51 56.5617
R940 VN.n12 VN.n11 53.9797
R941 VN.n57 VN.n56 53.9797
R942 VN.n40 VN.n2 51.7179
R943 VN.n85 VN.n47 51.7179
R944 VN.n36 VN.n2 29.4362
R945 VN.n81 VN.n47 29.4362
R946 VN.n13 VN.n10 24.5923
R947 VN.n17 VN.n10 24.5923
R948 VN.n19 VN.n18 24.5923
R949 VN.n19 VN.n8 24.5923
R950 VN.n23 VN.n8 24.5923
R951 VN.n24 VN.n23 24.5923
R952 VN.n25 VN.n24 24.5923
R953 VN.n25 VN.n6 24.5923
R954 VN.n30 VN.n29 24.5923
R955 VN.n31 VN.n30 24.5923
R956 VN.n35 VN.n34 24.5923
R957 VN.n36 VN.n35 24.5923
R958 VN.n41 VN.n40 24.5923
R959 VN.n42 VN.n41 24.5923
R960 VN.n62 VN.n55 24.5923
R961 VN.n58 VN.n55 24.5923
R962 VN.n70 VN.n51 24.5923
R963 VN.n70 VN.n69 24.5923
R964 VN.n69 VN.n68 24.5923
R965 VN.n68 VN.n53 24.5923
R966 VN.n64 VN.n53 24.5923
R967 VN.n64 VN.n63 24.5923
R968 VN.n81 VN.n80 24.5923
R969 VN.n80 VN.n79 24.5923
R970 VN.n76 VN.n75 24.5923
R971 VN.n75 VN.n74 24.5923
R972 VN.n87 VN.n86 24.5923
R973 VN.n86 VN.n85 24.5923
R974 VN.n13 VN.n12 20.1658
R975 VN.n31 VN.n4 20.1658
R976 VN.n58 VN.n57 20.1658
R977 VN.n76 VN.n49 20.1658
R978 VN.n42 VN.n0 15.7393
R979 VN.n87 VN.n45 15.7393
R980 VN.n34 VN.n4 4.42703
R981 VN.n79 VN.n49 4.42703
R982 VN.n59 VN.n56 4.10082
R983 VN.n14 VN.n11 4.10082
R984 VN.n89 VN.n88 0.354861
R985 VN.n44 VN.n43 0.354861
R986 VN VN.n44 0.267071
R987 VN.n88 VN.n46 0.189894
R988 VN.n84 VN.n46 0.189894
R989 VN.n84 VN.n83 0.189894
R990 VN.n83 VN.n82 0.189894
R991 VN.n82 VN.n48 0.189894
R992 VN.n78 VN.n48 0.189894
R993 VN.n78 VN.n77 0.189894
R994 VN.n77 VN.n50 0.189894
R995 VN.n73 VN.n50 0.189894
R996 VN.n73 VN.n72 0.189894
R997 VN.n72 VN.n71 0.189894
R998 VN.n71 VN.n52 0.189894
R999 VN.n67 VN.n52 0.189894
R1000 VN.n67 VN.n66 0.189894
R1001 VN.n66 VN.n65 0.189894
R1002 VN.n65 VN.n54 0.189894
R1003 VN.n61 VN.n54 0.189894
R1004 VN.n61 VN.n60 0.189894
R1005 VN.n60 VN.n59 0.189894
R1006 VN.n15 VN.n14 0.189894
R1007 VN.n16 VN.n15 0.189894
R1008 VN.n16 VN.n9 0.189894
R1009 VN.n20 VN.n9 0.189894
R1010 VN.n21 VN.n20 0.189894
R1011 VN.n22 VN.n21 0.189894
R1012 VN.n22 VN.n7 0.189894
R1013 VN.n26 VN.n7 0.189894
R1014 VN.n27 VN.n26 0.189894
R1015 VN.n28 VN.n27 0.189894
R1016 VN.n28 VN.n5 0.189894
R1017 VN.n32 VN.n5 0.189894
R1018 VN.n33 VN.n32 0.189894
R1019 VN.n33 VN.n3 0.189894
R1020 VN.n37 VN.n3 0.189894
R1021 VN.n38 VN.n37 0.189894
R1022 VN.n39 VN.n38 0.189894
R1023 VN.n39 VN.n1 0.189894
R1024 VN.n43 VN.n1 0.189894
R1025 VDD2.n145 VDD2.n77 756.745
R1026 VDD2.n68 VDD2.n0 756.745
R1027 VDD2.n146 VDD2.n145 585
R1028 VDD2.n144 VDD2.n143 585
R1029 VDD2.n81 VDD2.n80 585
R1030 VDD2.n138 VDD2.n137 585
R1031 VDD2.n136 VDD2.n135 585
R1032 VDD2.n85 VDD2.n84 585
R1033 VDD2.n130 VDD2.n129 585
R1034 VDD2.n128 VDD2.n127 585
R1035 VDD2.n89 VDD2.n88 585
R1036 VDD2.n93 VDD2.n91 585
R1037 VDD2.n122 VDD2.n121 585
R1038 VDD2.n120 VDD2.n119 585
R1039 VDD2.n95 VDD2.n94 585
R1040 VDD2.n114 VDD2.n113 585
R1041 VDD2.n112 VDD2.n111 585
R1042 VDD2.n99 VDD2.n98 585
R1043 VDD2.n106 VDD2.n105 585
R1044 VDD2.n104 VDD2.n103 585
R1045 VDD2.n25 VDD2.n24 585
R1046 VDD2.n27 VDD2.n26 585
R1047 VDD2.n20 VDD2.n19 585
R1048 VDD2.n33 VDD2.n32 585
R1049 VDD2.n35 VDD2.n34 585
R1050 VDD2.n16 VDD2.n15 585
R1051 VDD2.n42 VDD2.n41 585
R1052 VDD2.n43 VDD2.n14 585
R1053 VDD2.n45 VDD2.n44 585
R1054 VDD2.n12 VDD2.n11 585
R1055 VDD2.n51 VDD2.n50 585
R1056 VDD2.n53 VDD2.n52 585
R1057 VDD2.n8 VDD2.n7 585
R1058 VDD2.n59 VDD2.n58 585
R1059 VDD2.n61 VDD2.n60 585
R1060 VDD2.n4 VDD2.n3 585
R1061 VDD2.n67 VDD2.n66 585
R1062 VDD2.n69 VDD2.n68 585
R1063 VDD2.n102 VDD2.t7 329.036
R1064 VDD2.n23 VDD2.t0 329.036
R1065 VDD2.n145 VDD2.n144 171.744
R1066 VDD2.n144 VDD2.n80 171.744
R1067 VDD2.n137 VDD2.n80 171.744
R1068 VDD2.n137 VDD2.n136 171.744
R1069 VDD2.n136 VDD2.n84 171.744
R1070 VDD2.n129 VDD2.n84 171.744
R1071 VDD2.n129 VDD2.n128 171.744
R1072 VDD2.n128 VDD2.n88 171.744
R1073 VDD2.n93 VDD2.n88 171.744
R1074 VDD2.n121 VDD2.n93 171.744
R1075 VDD2.n121 VDD2.n120 171.744
R1076 VDD2.n120 VDD2.n94 171.744
R1077 VDD2.n113 VDD2.n94 171.744
R1078 VDD2.n113 VDD2.n112 171.744
R1079 VDD2.n112 VDD2.n98 171.744
R1080 VDD2.n105 VDD2.n98 171.744
R1081 VDD2.n105 VDD2.n104 171.744
R1082 VDD2.n26 VDD2.n25 171.744
R1083 VDD2.n26 VDD2.n19 171.744
R1084 VDD2.n33 VDD2.n19 171.744
R1085 VDD2.n34 VDD2.n33 171.744
R1086 VDD2.n34 VDD2.n15 171.744
R1087 VDD2.n42 VDD2.n15 171.744
R1088 VDD2.n43 VDD2.n42 171.744
R1089 VDD2.n44 VDD2.n43 171.744
R1090 VDD2.n44 VDD2.n11 171.744
R1091 VDD2.n51 VDD2.n11 171.744
R1092 VDD2.n52 VDD2.n51 171.744
R1093 VDD2.n52 VDD2.n7 171.744
R1094 VDD2.n59 VDD2.n7 171.744
R1095 VDD2.n60 VDD2.n59 171.744
R1096 VDD2.n60 VDD2.n3 171.744
R1097 VDD2.n67 VDD2.n3 171.744
R1098 VDD2.n68 VDD2.n67 171.744
R1099 VDD2.n104 VDD2.t7 85.8723
R1100 VDD2.n25 VDD2.t0 85.8723
R1101 VDD2.n76 VDD2.n75 73.6543
R1102 VDD2 VDD2.n153 73.6515
R1103 VDD2.n152 VDD2.n151 71.5051
R1104 VDD2.n74 VDD2.n73 71.5049
R1105 VDD2.n74 VDD2.n72 51.028
R1106 VDD2.n150 VDD2.n76 49.3338
R1107 VDD2.n150 VDD2.n149 48.0884
R1108 VDD2.n91 VDD2.n89 13.1884
R1109 VDD2.n45 VDD2.n12 13.1884
R1110 VDD2.n127 VDD2.n126 12.8005
R1111 VDD2.n123 VDD2.n122 12.8005
R1112 VDD2.n46 VDD2.n14 12.8005
R1113 VDD2.n50 VDD2.n49 12.8005
R1114 VDD2.n130 VDD2.n87 12.0247
R1115 VDD2.n119 VDD2.n92 12.0247
R1116 VDD2.n41 VDD2.n40 12.0247
R1117 VDD2.n53 VDD2.n10 12.0247
R1118 VDD2.n131 VDD2.n85 11.249
R1119 VDD2.n118 VDD2.n95 11.249
R1120 VDD2.n39 VDD2.n16 11.249
R1121 VDD2.n54 VDD2.n8 11.249
R1122 VDD2.n103 VDD2.n102 10.7239
R1123 VDD2.n24 VDD2.n23 10.7239
R1124 VDD2.n135 VDD2.n134 10.4732
R1125 VDD2.n115 VDD2.n114 10.4732
R1126 VDD2.n36 VDD2.n35 10.4732
R1127 VDD2.n58 VDD2.n57 10.4732
R1128 VDD2.n138 VDD2.n83 9.69747
R1129 VDD2.n111 VDD2.n97 9.69747
R1130 VDD2.n32 VDD2.n18 9.69747
R1131 VDD2.n61 VDD2.n6 9.69747
R1132 VDD2.n149 VDD2.n148 9.45567
R1133 VDD2.n72 VDD2.n71 9.45567
R1134 VDD2.n101 VDD2.n100 9.3005
R1135 VDD2.n108 VDD2.n107 9.3005
R1136 VDD2.n110 VDD2.n109 9.3005
R1137 VDD2.n97 VDD2.n96 9.3005
R1138 VDD2.n116 VDD2.n115 9.3005
R1139 VDD2.n118 VDD2.n117 9.3005
R1140 VDD2.n92 VDD2.n90 9.3005
R1141 VDD2.n124 VDD2.n123 9.3005
R1142 VDD2.n148 VDD2.n147 9.3005
R1143 VDD2.n79 VDD2.n78 9.3005
R1144 VDD2.n142 VDD2.n141 9.3005
R1145 VDD2.n140 VDD2.n139 9.3005
R1146 VDD2.n83 VDD2.n82 9.3005
R1147 VDD2.n134 VDD2.n133 9.3005
R1148 VDD2.n132 VDD2.n131 9.3005
R1149 VDD2.n87 VDD2.n86 9.3005
R1150 VDD2.n126 VDD2.n125 9.3005
R1151 VDD2.n71 VDD2.n70 9.3005
R1152 VDD2.n65 VDD2.n64 9.3005
R1153 VDD2.n63 VDD2.n62 9.3005
R1154 VDD2.n6 VDD2.n5 9.3005
R1155 VDD2.n57 VDD2.n56 9.3005
R1156 VDD2.n55 VDD2.n54 9.3005
R1157 VDD2.n10 VDD2.n9 9.3005
R1158 VDD2.n49 VDD2.n48 9.3005
R1159 VDD2.n22 VDD2.n21 9.3005
R1160 VDD2.n29 VDD2.n28 9.3005
R1161 VDD2.n31 VDD2.n30 9.3005
R1162 VDD2.n18 VDD2.n17 9.3005
R1163 VDD2.n37 VDD2.n36 9.3005
R1164 VDD2.n39 VDD2.n38 9.3005
R1165 VDD2.n40 VDD2.n13 9.3005
R1166 VDD2.n47 VDD2.n46 9.3005
R1167 VDD2.n2 VDD2.n1 9.3005
R1168 VDD2.n139 VDD2.n81 8.92171
R1169 VDD2.n110 VDD2.n99 8.92171
R1170 VDD2.n31 VDD2.n20 8.92171
R1171 VDD2.n62 VDD2.n4 8.92171
R1172 VDD2.n143 VDD2.n142 8.14595
R1173 VDD2.n107 VDD2.n106 8.14595
R1174 VDD2.n28 VDD2.n27 8.14595
R1175 VDD2.n66 VDD2.n65 8.14595
R1176 VDD2.n149 VDD2.n77 7.3702
R1177 VDD2.n146 VDD2.n79 7.3702
R1178 VDD2.n103 VDD2.n101 7.3702
R1179 VDD2.n24 VDD2.n22 7.3702
R1180 VDD2.n69 VDD2.n2 7.3702
R1181 VDD2.n72 VDD2.n0 7.3702
R1182 VDD2.n147 VDD2.n77 6.59444
R1183 VDD2.n147 VDD2.n146 6.59444
R1184 VDD2.n70 VDD2.n69 6.59444
R1185 VDD2.n70 VDD2.n0 6.59444
R1186 VDD2.n143 VDD2.n79 5.81868
R1187 VDD2.n106 VDD2.n101 5.81868
R1188 VDD2.n27 VDD2.n22 5.81868
R1189 VDD2.n66 VDD2.n2 5.81868
R1190 VDD2.n142 VDD2.n81 5.04292
R1191 VDD2.n107 VDD2.n99 5.04292
R1192 VDD2.n28 VDD2.n20 5.04292
R1193 VDD2.n65 VDD2.n4 5.04292
R1194 VDD2.n139 VDD2.n138 4.26717
R1195 VDD2.n111 VDD2.n110 4.26717
R1196 VDD2.n32 VDD2.n31 4.26717
R1197 VDD2.n62 VDD2.n61 4.26717
R1198 VDD2.n135 VDD2.n83 3.49141
R1199 VDD2.n114 VDD2.n97 3.49141
R1200 VDD2.n35 VDD2.n18 3.49141
R1201 VDD2.n58 VDD2.n6 3.49141
R1202 VDD2.n152 VDD2.n150 2.94016
R1203 VDD2.n134 VDD2.n85 2.71565
R1204 VDD2.n115 VDD2.n95 2.71565
R1205 VDD2.n36 VDD2.n16 2.71565
R1206 VDD2.n57 VDD2.n8 2.71565
R1207 VDD2.n102 VDD2.n100 2.41282
R1208 VDD2.n23 VDD2.n21 2.41282
R1209 VDD2.n153 VDD2.t4 2.40472
R1210 VDD2.n153 VDD2.t1 2.40472
R1211 VDD2.n151 VDD2.t2 2.40472
R1212 VDD2.n151 VDD2.t8 2.40472
R1213 VDD2.n75 VDD2.t3 2.40472
R1214 VDD2.n75 VDD2.t6 2.40472
R1215 VDD2.n73 VDD2.t5 2.40472
R1216 VDD2.n73 VDD2.t9 2.40472
R1217 VDD2.n131 VDD2.n130 1.93989
R1218 VDD2.n119 VDD2.n118 1.93989
R1219 VDD2.n41 VDD2.n39 1.93989
R1220 VDD2.n54 VDD2.n53 1.93989
R1221 VDD2.n127 VDD2.n87 1.16414
R1222 VDD2.n122 VDD2.n92 1.16414
R1223 VDD2.n40 VDD2.n14 1.16414
R1224 VDD2.n50 VDD2.n10 1.16414
R1225 VDD2 VDD2.n152 0.793603
R1226 VDD2.n76 VDD2.n74 0.680068
R1227 VDD2.n126 VDD2.n89 0.388379
R1228 VDD2.n123 VDD2.n91 0.388379
R1229 VDD2.n46 VDD2.n45 0.388379
R1230 VDD2.n49 VDD2.n12 0.388379
R1231 VDD2.n148 VDD2.n78 0.155672
R1232 VDD2.n141 VDD2.n78 0.155672
R1233 VDD2.n141 VDD2.n140 0.155672
R1234 VDD2.n140 VDD2.n82 0.155672
R1235 VDD2.n133 VDD2.n82 0.155672
R1236 VDD2.n133 VDD2.n132 0.155672
R1237 VDD2.n132 VDD2.n86 0.155672
R1238 VDD2.n125 VDD2.n86 0.155672
R1239 VDD2.n125 VDD2.n124 0.155672
R1240 VDD2.n124 VDD2.n90 0.155672
R1241 VDD2.n117 VDD2.n90 0.155672
R1242 VDD2.n117 VDD2.n116 0.155672
R1243 VDD2.n116 VDD2.n96 0.155672
R1244 VDD2.n109 VDD2.n96 0.155672
R1245 VDD2.n109 VDD2.n108 0.155672
R1246 VDD2.n108 VDD2.n100 0.155672
R1247 VDD2.n29 VDD2.n21 0.155672
R1248 VDD2.n30 VDD2.n29 0.155672
R1249 VDD2.n30 VDD2.n17 0.155672
R1250 VDD2.n37 VDD2.n17 0.155672
R1251 VDD2.n38 VDD2.n37 0.155672
R1252 VDD2.n38 VDD2.n13 0.155672
R1253 VDD2.n47 VDD2.n13 0.155672
R1254 VDD2.n48 VDD2.n47 0.155672
R1255 VDD2.n48 VDD2.n9 0.155672
R1256 VDD2.n55 VDD2.n9 0.155672
R1257 VDD2.n56 VDD2.n55 0.155672
R1258 VDD2.n56 VDD2.n5 0.155672
R1259 VDD2.n63 VDD2.n5 0.155672
R1260 VDD2.n64 VDD2.n63 0.155672
R1261 VDD2.n64 VDD2.n1 0.155672
R1262 VDD2.n71 VDD2.n1 0.155672
R1263 B.n710 B.n91 585
R1264 B.n712 B.n711 585
R1265 B.n713 B.n90 585
R1266 B.n715 B.n714 585
R1267 B.n716 B.n89 585
R1268 B.n718 B.n717 585
R1269 B.n719 B.n88 585
R1270 B.n721 B.n720 585
R1271 B.n722 B.n87 585
R1272 B.n724 B.n723 585
R1273 B.n725 B.n86 585
R1274 B.n727 B.n726 585
R1275 B.n728 B.n85 585
R1276 B.n730 B.n729 585
R1277 B.n731 B.n84 585
R1278 B.n733 B.n732 585
R1279 B.n734 B.n83 585
R1280 B.n736 B.n735 585
R1281 B.n737 B.n82 585
R1282 B.n739 B.n738 585
R1283 B.n740 B.n81 585
R1284 B.n742 B.n741 585
R1285 B.n743 B.n80 585
R1286 B.n745 B.n744 585
R1287 B.n746 B.n79 585
R1288 B.n748 B.n747 585
R1289 B.n749 B.n78 585
R1290 B.n751 B.n750 585
R1291 B.n752 B.n77 585
R1292 B.n754 B.n753 585
R1293 B.n755 B.n76 585
R1294 B.n757 B.n756 585
R1295 B.n758 B.n75 585
R1296 B.n760 B.n759 585
R1297 B.n761 B.n74 585
R1298 B.n763 B.n762 585
R1299 B.n764 B.n73 585
R1300 B.n766 B.n765 585
R1301 B.n767 B.n72 585
R1302 B.n769 B.n768 585
R1303 B.n770 B.n71 585
R1304 B.n772 B.n771 585
R1305 B.n773 B.n70 585
R1306 B.n775 B.n774 585
R1307 B.n776 B.n69 585
R1308 B.n778 B.n777 585
R1309 B.n780 B.n779 585
R1310 B.n781 B.n65 585
R1311 B.n783 B.n782 585
R1312 B.n784 B.n64 585
R1313 B.n786 B.n785 585
R1314 B.n787 B.n63 585
R1315 B.n789 B.n788 585
R1316 B.n790 B.n62 585
R1317 B.n792 B.n791 585
R1318 B.n793 B.n59 585
R1319 B.n796 B.n795 585
R1320 B.n797 B.n58 585
R1321 B.n799 B.n798 585
R1322 B.n800 B.n57 585
R1323 B.n802 B.n801 585
R1324 B.n803 B.n56 585
R1325 B.n805 B.n804 585
R1326 B.n806 B.n55 585
R1327 B.n808 B.n807 585
R1328 B.n809 B.n54 585
R1329 B.n811 B.n810 585
R1330 B.n812 B.n53 585
R1331 B.n814 B.n813 585
R1332 B.n815 B.n52 585
R1333 B.n817 B.n816 585
R1334 B.n818 B.n51 585
R1335 B.n820 B.n819 585
R1336 B.n821 B.n50 585
R1337 B.n823 B.n822 585
R1338 B.n824 B.n49 585
R1339 B.n826 B.n825 585
R1340 B.n827 B.n48 585
R1341 B.n829 B.n828 585
R1342 B.n830 B.n47 585
R1343 B.n832 B.n831 585
R1344 B.n833 B.n46 585
R1345 B.n835 B.n834 585
R1346 B.n836 B.n45 585
R1347 B.n838 B.n837 585
R1348 B.n839 B.n44 585
R1349 B.n841 B.n840 585
R1350 B.n842 B.n43 585
R1351 B.n844 B.n843 585
R1352 B.n845 B.n42 585
R1353 B.n847 B.n846 585
R1354 B.n848 B.n41 585
R1355 B.n850 B.n849 585
R1356 B.n851 B.n40 585
R1357 B.n853 B.n852 585
R1358 B.n854 B.n39 585
R1359 B.n856 B.n855 585
R1360 B.n857 B.n38 585
R1361 B.n859 B.n858 585
R1362 B.n860 B.n37 585
R1363 B.n862 B.n861 585
R1364 B.n863 B.n36 585
R1365 B.n709 B.n708 585
R1366 B.n707 B.n92 585
R1367 B.n706 B.n705 585
R1368 B.n704 B.n93 585
R1369 B.n703 B.n702 585
R1370 B.n701 B.n94 585
R1371 B.n700 B.n699 585
R1372 B.n698 B.n95 585
R1373 B.n697 B.n696 585
R1374 B.n695 B.n96 585
R1375 B.n694 B.n693 585
R1376 B.n692 B.n97 585
R1377 B.n691 B.n690 585
R1378 B.n689 B.n98 585
R1379 B.n688 B.n687 585
R1380 B.n686 B.n99 585
R1381 B.n685 B.n684 585
R1382 B.n683 B.n100 585
R1383 B.n682 B.n681 585
R1384 B.n680 B.n101 585
R1385 B.n679 B.n678 585
R1386 B.n677 B.n102 585
R1387 B.n676 B.n675 585
R1388 B.n674 B.n103 585
R1389 B.n673 B.n672 585
R1390 B.n671 B.n104 585
R1391 B.n670 B.n669 585
R1392 B.n668 B.n105 585
R1393 B.n667 B.n666 585
R1394 B.n665 B.n106 585
R1395 B.n664 B.n663 585
R1396 B.n662 B.n107 585
R1397 B.n661 B.n660 585
R1398 B.n659 B.n108 585
R1399 B.n658 B.n657 585
R1400 B.n656 B.n109 585
R1401 B.n655 B.n654 585
R1402 B.n653 B.n110 585
R1403 B.n652 B.n651 585
R1404 B.n650 B.n111 585
R1405 B.n649 B.n648 585
R1406 B.n647 B.n112 585
R1407 B.n646 B.n645 585
R1408 B.n644 B.n113 585
R1409 B.n643 B.n642 585
R1410 B.n641 B.n114 585
R1411 B.n640 B.n639 585
R1412 B.n638 B.n115 585
R1413 B.n637 B.n636 585
R1414 B.n635 B.n116 585
R1415 B.n634 B.n633 585
R1416 B.n632 B.n117 585
R1417 B.n631 B.n630 585
R1418 B.n629 B.n118 585
R1419 B.n628 B.n627 585
R1420 B.n626 B.n119 585
R1421 B.n625 B.n624 585
R1422 B.n623 B.n120 585
R1423 B.n622 B.n621 585
R1424 B.n620 B.n121 585
R1425 B.n619 B.n618 585
R1426 B.n617 B.n122 585
R1427 B.n616 B.n615 585
R1428 B.n614 B.n123 585
R1429 B.n613 B.n612 585
R1430 B.n611 B.n124 585
R1431 B.n610 B.n609 585
R1432 B.n608 B.n125 585
R1433 B.n607 B.n606 585
R1434 B.n605 B.n126 585
R1435 B.n604 B.n603 585
R1436 B.n602 B.n127 585
R1437 B.n601 B.n600 585
R1438 B.n599 B.n128 585
R1439 B.n598 B.n597 585
R1440 B.n596 B.n129 585
R1441 B.n595 B.n594 585
R1442 B.n593 B.n130 585
R1443 B.n592 B.n591 585
R1444 B.n590 B.n131 585
R1445 B.n589 B.n588 585
R1446 B.n587 B.n132 585
R1447 B.n586 B.n585 585
R1448 B.n584 B.n133 585
R1449 B.n583 B.n582 585
R1450 B.n581 B.n134 585
R1451 B.n580 B.n579 585
R1452 B.n578 B.n135 585
R1453 B.n577 B.n576 585
R1454 B.n575 B.n136 585
R1455 B.n574 B.n573 585
R1456 B.n572 B.n137 585
R1457 B.n571 B.n570 585
R1458 B.n569 B.n138 585
R1459 B.n568 B.n567 585
R1460 B.n566 B.n139 585
R1461 B.n565 B.n564 585
R1462 B.n563 B.n140 585
R1463 B.n562 B.n561 585
R1464 B.n560 B.n141 585
R1465 B.n559 B.n558 585
R1466 B.n557 B.n142 585
R1467 B.n556 B.n555 585
R1468 B.n554 B.n143 585
R1469 B.n553 B.n552 585
R1470 B.n551 B.n144 585
R1471 B.n550 B.n549 585
R1472 B.n548 B.n145 585
R1473 B.n547 B.n546 585
R1474 B.n545 B.n146 585
R1475 B.n544 B.n543 585
R1476 B.n542 B.n147 585
R1477 B.n541 B.n540 585
R1478 B.n539 B.n148 585
R1479 B.n538 B.n537 585
R1480 B.n536 B.n149 585
R1481 B.n535 B.n534 585
R1482 B.n533 B.n150 585
R1483 B.n532 B.n531 585
R1484 B.n530 B.n151 585
R1485 B.n529 B.n528 585
R1486 B.n527 B.n152 585
R1487 B.n526 B.n525 585
R1488 B.n524 B.n153 585
R1489 B.n523 B.n522 585
R1490 B.n521 B.n154 585
R1491 B.n520 B.n519 585
R1492 B.n518 B.n155 585
R1493 B.n517 B.n516 585
R1494 B.n515 B.n156 585
R1495 B.n514 B.n513 585
R1496 B.n512 B.n157 585
R1497 B.n511 B.n510 585
R1498 B.n509 B.n158 585
R1499 B.n508 B.n507 585
R1500 B.n506 B.n159 585
R1501 B.n505 B.n504 585
R1502 B.n350 B.n215 585
R1503 B.n352 B.n351 585
R1504 B.n353 B.n214 585
R1505 B.n355 B.n354 585
R1506 B.n356 B.n213 585
R1507 B.n358 B.n357 585
R1508 B.n359 B.n212 585
R1509 B.n361 B.n360 585
R1510 B.n362 B.n211 585
R1511 B.n364 B.n363 585
R1512 B.n365 B.n210 585
R1513 B.n367 B.n366 585
R1514 B.n368 B.n209 585
R1515 B.n370 B.n369 585
R1516 B.n371 B.n208 585
R1517 B.n373 B.n372 585
R1518 B.n374 B.n207 585
R1519 B.n376 B.n375 585
R1520 B.n377 B.n206 585
R1521 B.n379 B.n378 585
R1522 B.n380 B.n205 585
R1523 B.n382 B.n381 585
R1524 B.n383 B.n204 585
R1525 B.n385 B.n384 585
R1526 B.n386 B.n203 585
R1527 B.n388 B.n387 585
R1528 B.n389 B.n202 585
R1529 B.n391 B.n390 585
R1530 B.n392 B.n201 585
R1531 B.n394 B.n393 585
R1532 B.n395 B.n200 585
R1533 B.n397 B.n396 585
R1534 B.n398 B.n199 585
R1535 B.n400 B.n399 585
R1536 B.n401 B.n198 585
R1537 B.n403 B.n402 585
R1538 B.n404 B.n197 585
R1539 B.n406 B.n405 585
R1540 B.n407 B.n196 585
R1541 B.n409 B.n408 585
R1542 B.n410 B.n195 585
R1543 B.n412 B.n411 585
R1544 B.n413 B.n194 585
R1545 B.n415 B.n414 585
R1546 B.n416 B.n193 585
R1547 B.n418 B.n417 585
R1548 B.n420 B.n419 585
R1549 B.n421 B.n189 585
R1550 B.n423 B.n422 585
R1551 B.n424 B.n188 585
R1552 B.n426 B.n425 585
R1553 B.n427 B.n187 585
R1554 B.n429 B.n428 585
R1555 B.n430 B.n186 585
R1556 B.n432 B.n431 585
R1557 B.n433 B.n183 585
R1558 B.n436 B.n435 585
R1559 B.n437 B.n182 585
R1560 B.n439 B.n438 585
R1561 B.n440 B.n181 585
R1562 B.n442 B.n441 585
R1563 B.n443 B.n180 585
R1564 B.n445 B.n444 585
R1565 B.n446 B.n179 585
R1566 B.n448 B.n447 585
R1567 B.n449 B.n178 585
R1568 B.n451 B.n450 585
R1569 B.n452 B.n177 585
R1570 B.n454 B.n453 585
R1571 B.n455 B.n176 585
R1572 B.n457 B.n456 585
R1573 B.n458 B.n175 585
R1574 B.n460 B.n459 585
R1575 B.n461 B.n174 585
R1576 B.n463 B.n462 585
R1577 B.n464 B.n173 585
R1578 B.n466 B.n465 585
R1579 B.n467 B.n172 585
R1580 B.n469 B.n468 585
R1581 B.n470 B.n171 585
R1582 B.n472 B.n471 585
R1583 B.n473 B.n170 585
R1584 B.n475 B.n474 585
R1585 B.n476 B.n169 585
R1586 B.n478 B.n477 585
R1587 B.n479 B.n168 585
R1588 B.n481 B.n480 585
R1589 B.n482 B.n167 585
R1590 B.n484 B.n483 585
R1591 B.n485 B.n166 585
R1592 B.n487 B.n486 585
R1593 B.n488 B.n165 585
R1594 B.n490 B.n489 585
R1595 B.n491 B.n164 585
R1596 B.n493 B.n492 585
R1597 B.n494 B.n163 585
R1598 B.n496 B.n495 585
R1599 B.n497 B.n162 585
R1600 B.n499 B.n498 585
R1601 B.n500 B.n161 585
R1602 B.n502 B.n501 585
R1603 B.n503 B.n160 585
R1604 B.n349 B.n348 585
R1605 B.n347 B.n216 585
R1606 B.n346 B.n345 585
R1607 B.n344 B.n217 585
R1608 B.n343 B.n342 585
R1609 B.n341 B.n218 585
R1610 B.n340 B.n339 585
R1611 B.n338 B.n219 585
R1612 B.n337 B.n336 585
R1613 B.n335 B.n220 585
R1614 B.n334 B.n333 585
R1615 B.n332 B.n221 585
R1616 B.n331 B.n330 585
R1617 B.n329 B.n222 585
R1618 B.n328 B.n327 585
R1619 B.n326 B.n223 585
R1620 B.n325 B.n324 585
R1621 B.n323 B.n224 585
R1622 B.n322 B.n321 585
R1623 B.n320 B.n225 585
R1624 B.n319 B.n318 585
R1625 B.n317 B.n226 585
R1626 B.n316 B.n315 585
R1627 B.n314 B.n227 585
R1628 B.n313 B.n312 585
R1629 B.n311 B.n228 585
R1630 B.n310 B.n309 585
R1631 B.n308 B.n229 585
R1632 B.n307 B.n306 585
R1633 B.n305 B.n230 585
R1634 B.n304 B.n303 585
R1635 B.n302 B.n231 585
R1636 B.n301 B.n300 585
R1637 B.n299 B.n232 585
R1638 B.n298 B.n297 585
R1639 B.n296 B.n233 585
R1640 B.n295 B.n294 585
R1641 B.n293 B.n234 585
R1642 B.n292 B.n291 585
R1643 B.n290 B.n235 585
R1644 B.n289 B.n288 585
R1645 B.n287 B.n236 585
R1646 B.n286 B.n285 585
R1647 B.n284 B.n237 585
R1648 B.n283 B.n282 585
R1649 B.n281 B.n238 585
R1650 B.n280 B.n279 585
R1651 B.n278 B.n239 585
R1652 B.n277 B.n276 585
R1653 B.n275 B.n240 585
R1654 B.n274 B.n273 585
R1655 B.n272 B.n241 585
R1656 B.n271 B.n270 585
R1657 B.n269 B.n242 585
R1658 B.n268 B.n267 585
R1659 B.n266 B.n243 585
R1660 B.n265 B.n264 585
R1661 B.n263 B.n244 585
R1662 B.n262 B.n261 585
R1663 B.n260 B.n245 585
R1664 B.n259 B.n258 585
R1665 B.n257 B.n246 585
R1666 B.n256 B.n255 585
R1667 B.n254 B.n247 585
R1668 B.n253 B.n252 585
R1669 B.n251 B.n248 585
R1670 B.n250 B.n249 585
R1671 B.n2 B.n0 585
R1672 B.n965 B.n1 585
R1673 B.n964 B.n963 585
R1674 B.n962 B.n3 585
R1675 B.n961 B.n960 585
R1676 B.n959 B.n4 585
R1677 B.n958 B.n957 585
R1678 B.n956 B.n5 585
R1679 B.n955 B.n954 585
R1680 B.n953 B.n6 585
R1681 B.n952 B.n951 585
R1682 B.n950 B.n7 585
R1683 B.n949 B.n948 585
R1684 B.n947 B.n8 585
R1685 B.n946 B.n945 585
R1686 B.n944 B.n9 585
R1687 B.n943 B.n942 585
R1688 B.n941 B.n10 585
R1689 B.n940 B.n939 585
R1690 B.n938 B.n11 585
R1691 B.n937 B.n936 585
R1692 B.n935 B.n12 585
R1693 B.n934 B.n933 585
R1694 B.n932 B.n13 585
R1695 B.n931 B.n930 585
R1696 B.n929 B.n14 585
R1697 B.n928 B.n927 585
R1698 B.n926 B.n15 585
R1699 B.n925 B.n924 585
R1700 B.n923 B.n16 585
R1701 B.n922 B.n921 585
R1702 B.n920 B.n17 585
R1703 B.n919 B.n918 585
R1704 B.n917 B.n18 585
R1705 B.n916 B.n915 585
R1706 B.n914 B.n19 585
R1707 B.n913 B.n912 585
R1708 B.n911 B.n20 585
R1709 B.n910 B.n909 585
R1710 B.n908 B.n21 585
R1711 B.n907 B.n906 585
R1712 B.n905 B.n22 585
R1713 B.n904 B.n903 585
R1714 B.n902 B.n23 585
R1715 B.n901 B.n900 585
R1716 B.n899 B.n24 585
R1717 B.n898 B.n897 585
R1718 B.n896 B.n25 585
R1719 B.n895 B.n894 585
R1720 B.n893 B.n26 585
R1721 B.n892 B.n891 585
R1722 B.n890 B.n27 585
R1723 B.n889 B.n888 585
R1724 B.n887 B.n28 585
R1725 B.n886 B.n885 585
R1726 B.n884 B.n29 585
R1727 B.n883 B.n882 585
R1728 B.n881 B.n30 585
R1729 B.n880 B.n879 585
R1730 B.n878 B.n31 585
R1731 B.n877 B.n876 585
R1732 B.n875 B.n32 585
R1733 B.n874 B.n873 585
R1734 B.n872 B.n33 585
R1735 B.n871 B.n870 585
R1736 B.n869 B.n34 585
R1737 B.n868 B.n867 585
R1738 B.n866 B.n35 585
R1739 B.n865 B.n864 585
R1740 B.n967 B.n966 585
R1741 B.n348 B.n215 526.135
R1742 B.n864 B.n863 526.135
R1743 B.n504 B.n503 526.135
R1744 B.n708 B.n91 526.135
R1745 B.n184 B.t5 469.26
R1746 B.n66 B.t7 469.26
R1747 B.n190 B.t11 469.26
R1748 B.n60 B.t1 469.26
R1749 B.n185 B.t4 403.127
R1750 B.n67 B.t8 403.127
R1751 B.n191 B.t10 403.127
R1752 B.n61 B.t2 403.127
R1753 B.n184 B.t3 314.462
R1754 B.n190 B.t9 314.462
R1755 B.n60 B.t0 314.462
R1756 B.n66 B.t6 314.462
R1757 B.n348 B.n347 163.367
R1758 B.n347 B.n346 163.367
R1759 B.n346 B.n217 163.367
R1760 B.n342 B.n217 163.367
R1761 B.n342 B.n341 163.367
R1762 B.n341 B.n340 163.367
R1763 B.n340 B.n219 163.367
R1764 B.n336 B.n219 163.367
R1765 B.n336 B.n335 163.367
R1766 B.n335 B.n334 163.367
R1767 B.n334 B.n221 163.367
R1768 B.n330 B.n221 163.367
R1769 B.n330 B.n329 163.367
R1770 B.n329 B.n328 163.367
R1771 B.n328 B.n223 163.367
R1772 B.n324 B.n223 163.367
R1773 B.n324 B.n323 163.367
R1774 B.n323 B.n322 163.367
R1775 B.n322 B.n225 163.367
R1776 B.n318 B.n225 163.367
R1777 B.n318 B.n317 163.367
R1778 B.n317 B.n316 163.367
R1779 B.n316 B.n227 163.367
R1780 B.n312 B.n227 163.367
R1781 B.n312 B.n311 163.367
R1782 B.n311 B.n310 163.367
R1783 B.n310 B.n229 163.367
R1784 B.n306 B.n229 163.367
R1785 B.n306 B.n305 163.367
R1786 B.n305 B.n304 163.367
R1787 B.n304 B.n231 163.367
R1788 B.n300 B.n231 163.367
R1789 B.n300 B.n299 163.367
R1790 B.n299 B.n298 163.367
R1791 B.n298 B.n233 163.367
R1792 B.n294 B.n233 163.367
R1793 B.n294 B.n293 163.367
R1794 B.n293 B.n292 163.367
R1795 B.n292 B.n235 163.367
R1796 B.n288 B.n235 163.367
R1797 B.n288 B.n287 163.367
R1798 B.n287 B.n286 163.367
R1799 B.n286 B.n237 163.367
R1800 B.n282 B.n237 163.367
R1801 B.n282 B.n281 163.367
R1802 B.n281 B.n280 163.367
R1803 B.n280 B.n239 163.367
R1804 B.n276 B.n239 163.367
R1805 B.n276 B.n275 163.367
R1806 B.n275 B.n274 163.367
R1807 B.n274 B.n241 163.367
R1808 B.n270 B.n241 163.367
R1809 B.n270 B.n269 163.367
R1810 B.n269 B.n268 163.367
R1811 B.n268 B.n243 163.367
R1812 B.n264 B.n243 163.367
R1813 B.n264 B.n263 163.367
R1814 B.n263 B.n262 163.367
R1815 B.n262 B.n245 163.367
R1816 B.n258 B.n245 163.367
R1817 B.n258 B.n257 163.367
R1818 B.n257 B.n256 163.367
R1819 B.n256 B.n247 163.367
R1820 B.n252 B.n247 163.367
R1821 B.n252 B.n251 163.367
R1822 B.n251 B.n250 163.367
R1823 B.n250 B.n2 163.367
R1824 B.n966 B.n2 163.367
R1825 B.n966 B.n965 163.367
R1826 B.n965 B.n964 163.367
R1827 B.n964 B.n3 163.367
R1828 B.n960 B.n3 163.367
R1829 B.n960 B.n959 163.367
R1830 B.n959 B.n958 163.367
R1831 B.n958 B.n5 163.367
R1832 B.n954 B.n5 163.367
R1833 B.n954 B.n953 163.367
R1834 B.n953 B.n952 163.367
R1835 B.n952 B.n7 163.367
R1836 B.n948 B.n7 163.367
R1837 B.n948 B.n947 163.367
R1838 B.n947 B.n946 163.367
R1839 B.n946 B.n9 163.367
R1840 B.n942 B.n9 163.367
R1841 B.n942 B.n941 163.367
R1842 B.n941 B.n940 163.367
R1843 B.n940 B.n11 163.367
R1844 B.n936 B.n11 163.367
R1845 B.n936 B.n935 163.367
R1846 B.n935 B.n934 163.367
R1847 B.n934 B.n13 163.367
R1848 B.n930 B.n13 163.367
R1849 B.n930 B.n929 163.367
R1850 B.n929 B.n928 163.367
R1851 B.n928 B.n15 163.367
R1852 B.n924 B.n15 163.367
R1853 B.n924 B.n923 163.367
R1854 B.n923 B.n922 163.367
R1855 B.n922 B.n17 163.367
R1856 B.n918 B.n17 163.367
R1857 B.n918 B.n917 163.367
R1858 B.n917 B.n916 163.367
R1859 B.n916 B.n19 163.367
R1860 B.n912 B.n19 163.367
R1861 B.n912 B.n911 163.367
R1862 B.n911 B.n910 163.367
R1863 B.n910 B.n21 163.367
R1864 B.n906 B.n21 163.367
R1865 B.n906 B.n905 163.367
R1866 B.n905 B.n904 163.367
R1867 B.n904 B.n23 163.367
R1868 B.n900 B.n23 163.367
R1869 B.n900 B.n899 163.367
R1870 B.n899 B.n898 163.367
R1871 B.n898 B.n25 163.367
R1872 B.n894 B.n25 163.367
R1873 B.n894 B.n893 163.367
R1874 B.n893 B.n892 163.367
R1875 B.n892 B.n27 163.367
R1876 B.n888 B.n27 163.367
R1877 B.n888 B.n887 163.367
R1878 B.n887 B.n886 163.367
R1879 B.n886 B.n29 163.367
R1880 B.n882 B.n29 163.367
R1881 B.n882 B.n881 163.367
R1882 B.n881 B.n880 163.367
R1883 B.n880 B.n31 163.367
R1884 B.n876 B.n31 163.367
R1885 B.n876 B.n875 163.367
R1886 B.n875 B.n874 163.367
R1887 B.n874 B.n33 163.367
R1888 B.n870 B.n33 163.367
R1889 B.n870 B.n869 163.367
R1890 B.n869 B.n868 163.367
R1891 B.n868 B.n35 163.367
R1892 B.n864 B.n35 163.367
R1893 B.n352 B.n215 163.367
R1894 B.n353 B.n352 163.367
R1895 B.n354 B.n353 163.367
R1896 B.n354 B.n213 163.367
R1897 B.n358 B.n213 163.367
R1898 B.n359 B.n358 163.367
R1899 B.n360 B.n359 163.367
R1900 B.n360 B.n211 163.367
R1901 B.n364 B.n211 163.367
R1902 B.n365 B.n364 163.367
R1903 B.n366 B.n365 163.367
R1904 B.n366 B.n209 163.367
R1905 B.n370 B.n209 163.367
R1906 B.n371 B.n370 163.367
R1907 B.n372 B.n371 163.367
R1908 B.n372 B.n207 163.367
R1909 B.n376 B.n207 163.367
R1910 B.n377 B.n376 163.367
R1911 B.n378 B.n377 163.367
R1912 B.n378 B.n205 163.367
R1913 B.n382 B.n205 163.367
R1914 B.n383 B.n382 163.367
R1915 B.n384 B.n383 163.367
R1916 B.n384 B.n203 163.367
R1917 B.n388 B.n203 163.367
R1918 B.n389 B.n388 163.367
R1919 B.n390 B.n389 163.367
R1920 B.n390 B.n201 163.367
R1921 B.n394 B.n201 163.367
R1922 B.n395 B.n394 163.367
R1923 B.n396 B.n395 163.367
R1924 B.n396 B.n199 163.367
R1925 B.n400 B.n199 163.367
R1926 B.n401 B.n400 163.367
R1927 B.n402 B.n401 163.367
R1928 B.n402 B.n197 163.367
R1929 B.n406 B.n197 163.367
R1930 B.n407 B.n406 163.367
R1931 B.n408 B.n407 163.367
R1932 B.n408 B.n195 163.367
R1933 B.n412 B.n195 163.367
R1934 B.n413 B.n412 163.367
R1935 B.n414 B.n413 163.367
R1936 B.n414 B.n193 163.367
R1937 B.n418 B.n193 163.367
R1938 B.n419 B.n418 163.367
R1939 B.n419 B.n189 163.367
R1940 B.n423 B.n189 163.367
R1941 B.n424 B.n423 163.367
R1942 B.n425 B.n424 163.367
R1943 B.n425 B.n187 163.367
R1944 B.n429 B.n187 163.367
R1945 B.n430 B.n429 163.367
R1946 B.n431 B.n430 163.367
R1947 B.n431 B.n183 163.367
R1948 B.n436 B.n183 163.367
R1949 B.n437 B.n436 163.367
R1950 B.n438 B.n437 163.367
R1951 B.n438 B.n181 163.367
R1952 B.n442 B.n181 163.367
R1953 B.n443 B.n442 163.367
R1954 B.n444 B.n443 163.367
R1955 B.n444 B.n179 163.367
R1956 B.n448 B.n179 163.367
R1957 B.n449 B.n448 163.367
R1958 B.n450 B.n449 163.367
R1959 B.n450 B.n177 163.367
R1960 B.n454 B.n177 163.367
R1961 B.n455 B.n454 163.367
R1962 B.n456 B.n455 163.367
R1963 B.n456 B.n175 163.367
R1964 B.n460 B.n175 163.367
R1965 B.n461 B.n460 163.367
R1966 B.n462 B.n461 163.367
R1967 B.n462 B.n173 163.367
R1968 B.n466 B.n173 163.367
R1969 B.n467 B.n466 163.367
R1970 B.n468 B.n467 163.367
R1971 B.n468 B.n171 163.367
R1972 B.n472 B.n171 163.367
R1973 B.n473 B.n472 163.367
R1974 B.n474 B.n473 163.367
R1975 B.n474 B.n169 163.367
R1976 B.n478 B.n169 163.367
R1977 B.n479 B.n478 163.367
R1978 B.n480 B.n479 163.367
R1979 B.n480 B.n167 163.367
R1980 B.n484 B.n167 163.367
R1981 B.n485 B.n484 163.367
R1982 B.n486 B.n485 163.367
R1983 B.n486 B.n165 163.367
R1984 B.n490 B.n165 163.367
R1985 B.n491 B.n490 163.367
R1986 B.n492 B.n491 163.367
R1987 B.n492 B.n163 163.367
R1988 B.n496 B.n163 163.367
R1989 B.n497 B.n496 163.367
R1990 B.n498 B.n497 163.367
R1991 B.n498 B.n161 163.367
R1992 B.n502 B.n161 163.367
R1993 B.n503 B.n502 163.367
R1994 B.n504 B.n159 163.367
R1995 B.n508 B.n159 163.367
R1996 B.n509 B.n508 163.367
R1997 B.n510 B.n509 163.367
R1998 B.n510 B.n157 163.367
R1999 B.n514 B.n157 163.367
R2000 B.n515 B.n514 163.367
R2001 B.n516 B.n515 163.367
R2002 B.n516 B.n155 163.367
R2003 B.n520 B.n155 163.367
R2004 B.n521 B.n520 163.367
R2005 B.n522 B.n521 163.367
R2006 B.n522 B.n153 163.367
R2007 B.n526 B.n153 163.367
R2008 B.n527 B.n526 163.367
R2009 B.n528 B.n527 163.367
R2010 B.n528 B.n151 163.367
R2011 B.n532 B.n151 163.367
R2012 B.n533 B.n532 163.367
R2013 B.n534 B.n533 163.367
R2014 B.n534 B.n149 163.367
R2015 B.n538 B.n149 163.367
R2016 B.n539 B.n538 163.367
R2017 B.n540 B.n539 163.367
R2018 B.n540 B.n147 163.367
R2019 B.n544 B.n147 163.367
R2020 B.n545 B.n544 163.367
R2021 B.n546 B.n545 163.367
R2022 B.n546 B.n145 163.367
R2023 B.n550 B.n145 163.367
R2024 B.n551 B.n550 163.367
R2025 B.n552 B.n551 163.367
R2026 B.n552 B.n143 163.367
R2027 B.n556 B.n143 163.367
R2028 B.n557 B.n556 163.367
R2029 B.n558 B.n557 163.367
R2030 B.n558 B.n141 163.367
R2031 B.n562 B.n141 163.367
R2032 B.n563 B.n562 163.367
R2033 B.n564 B.n563 163.367
R2034 B.n564 B.n139 163.367
R2035 B.n568 B.n139 163.367
R2036 B.n569 B.n568 163.367
R2037 B.n570 B.n569 163.367
R2038 B.n570 B.n137 163.367
R2039 B.n574 B.n137 163.367
R2040 B.n575 B.n574 163.367
R2041 B.n576 B.n575 163.367
R2042 B.n576 B.n135 163.367
R2043 B.n580 B.n135 163.367
R2044 B.n581 B.n580 163.367
R2045 B.n582 B.n581 163.367
R2046 B.n582 B.n133 163.367
R2047 B.n586 B.n133 163.367
R2048 B.n587 B.n586 163.367
R2049 B.n588 B.n587 163.367
R2050 B.n588 B.n131 163.367
R2051 B.n592 B.n131 163.367
R2052 B.n593 B.n592 163.367
R2053 B.n594 B.n593 163.367
R2054 B.n594 B.n129 163.367
R2055 B.n598 B.n129 163.367
R2056 B.n599 B.n598 163.367
R2057 B.n600 B.n599 163.367
R2058 B.n600 B.n127 163.367
R2059 B.n604 B.n127 163.367
R2060 B.n605 B.n604 163.367
R2061 B.n606 B.n605 163.367
R2062 B.n606 B.n125 163.367
R2063 B.n610 B.n125 163.367
R2064 B.n611 B.n610 163.367
R2065 B.n612 B.n611 163.367
R2066 B.n612 B.n123 163.367
R2067 B.n616 B.n123 163.367
R2068 B.n617 B.n616 163.367
R2069 B.n618 B.n617 163.367
R2070 B.n618 B.n121 163.367
R2071 B.n622 B.n121 163.367
R2072 B.n623 B.n622 163.367
R2073 B.n624 B.n623 163.367
R2074 B.n624 B.n119 163.367
R2075 B.n628 B.n119 163.367
R2076 B.n629 B.n628 163.367
R2077 B.n630 B.n629 163.367
R2078 B.n630 B.n117 163.367
R2079 B.n634 B.n117 163.367
R2080 B.n635 B.n634 163.367
R2081 B.n636 B.n635 163.367
R2082 B.n636 B.n115 163.367
R2083 B.n640 B.n115 163.367
R2084 B.n641 B.n640 163.367
R2085 B.n642 B.n641 163.367
R2086 B.n642 B.n113 163.367
R2087 B.n646 B.n113 163.367
R2088 B.n647 B.n646 163.367
R2089 B.n648 B.n647 163.367
R2090 B.n648 B.n111 163.367
R2091 B.n652 B.n111 163.367
R2092 B.n653 B.n652 163.367
R2093 B.n654 B.n653 163.367
R2094 B.n654 B.n109 163.367
R2095 B.n658 B.n109 163.367
R2096 B.n659 B.n658 163.367
R2097 B.n660 B.n659 163.367
R2098 B.n660 B.n107 163.367
R2099 B.n664 B.n107 163.367
R2100 B.n665 B.n664 163.367
R2101 B.n666 B.n665 163.367
R2102 B.n666 B.n105 163.367
R2103 B.n670 B.n105 163.367
R2104 B.n671 B.n670 163.367
R2105 B.n672 B.n671 163.367
R2106 B.n672 B.n103 163.367
R2107 B.n676 B.n103 163.367
R2108 B.n677 B.n676 163.367
R2109 B.n678 B.n677 163.367
R2110 B.n678 B.n101 163.367
R2111 B.n682 B.n101 163.367
R2112 B.n683 B.n682 163.367
R2113 B.n684 B.n683 163.367
R2114 B.n684 B.n99 163.367
R2115 B.n688 B.n99 163.367
R2116 B.n689 B.n688 163.367
R2117 B.n690 B.n689 163.367
R2118 B.n690 B.n97 163.367
R2119 B.n694 B.n97 163.367
R2120 B.n695 B.n694 163.367
R2121 B.n696 B.n695 163.367
R2122 B.n696 B.n95 163.367
R2123 B.n700 B.n95 163.367
R2124 B.n701 B.n700 163.367
R2125 B.n702 B.n701 163.367
R2126 B.n702 B.n93 163.367
R2127 B.n706 B.n93 163.367
R2128 B.n707 B.n706 163.367
R2129 B.n708 B.n707 163.367
R2130 B.n863 B.n862 163.367
R2131 B.n862 B.n37 163.367
R2132 B.n858 B.n37 163.367
R2133 B.n858 B.n857 163.367
R2134 B.n857 B.n856 163.367
R2135 B.n856 B.n39 163.367
R2136 B.n852 B.n39 163.367
R2137 B.n852 B.n851 163.367
R2138 B.n851 B.n850 163.367
R2139 B.n850 B.n41 163.367
R2140 B.n846 B.n41 163.367
R2141 B.n846 B.n845 163.367
R2142 B.n845 B.n844 163.367
R2143 B.n844 B.n43 163.367
R2144 B.n840 B.n43 163.367
R2145 B.n840 B.n839 163.367
R2146 B.n839 B.n838 163.367
R2147 B.n838 B.n45 163.367
R2148 B.n834 B.n45 163.367
R2149 B.n834 B.n833 163.367
R2150 B.n833 B.n832 163.367
R2151 B.n832 B.n47 163.367
R2152 B.n828 B.n47 163.367
R2153 B.n828 B.n827 163.367
R2154 B.n827 B.n826 163.367
R2155 B.n826 B.n49 163.367
R2156 B.n822 B.n49 163.367
R2157 B.n822 B.n821 163.367
R2158 B.n821 B.n820 163.367
R2159 B.n820 B.n51 163.367
R2160 B.n816 B.n51 163.367
R2161 B.n816 B.n815 163.367
R2162 B.n815 B.n814 163.367
R2163 B.n814 B.n53 163.367
R2164 B.n810 B.n53 163.367
R2165 B.n810 B.n809 163.367
R2166 B.n809 B.n808 163.367
R2167 B.n808 B.n55 163.367
R2168 B.n804 B.n55 163.367
R2169 B.n804 B.n803 163.367
R2170 B.n803 B.n802 163.367
R2171 B.n802 B.n57 163.367
R2172 B.n798 B.n57 163.367
R2173 B.n798 B.n797 163.367
R2174 B.n797 B.n796 163.367
R2175 B.n796 B.n59 163.367
R2176 B.n791 B.n59 163.367
R2177 B.n791 B.n790 163.367
R2178 B.n790 B.n789 163.367
R2179 B.n789 B.n63 163.367
R2180 B.n785 B.n63 163.367
R2181 B.n785 B.n784 163.367
R2182 B.n784 B.n783 163.367
R2183 B.n783 B.n65 163.367
R2184 B.n779 B.n65 163.367
R2185 B.n779 B.n778 163.367
R2186 B.n778 B.n69 163.367
R2187 B.n774 B.n69 163.367
R2188 B.n774 B.n773 163.367
R2189 B.n773 B.n772 163.367
R2190 B.n772 B.n71 163.367
R2191 B.n768 B.n71 163.367
R2192 B.n768 B.n767 163.367
R2193 B.n767 B.n766 163.367
R2194 B.n766 B.n73 163.367
R2195 B.n762 B.n73 163.367
R2196 B.n762 B.n761 163.367
R2197 B.n761 B.n760 163.367
R2198 B.n760 B.n75 163.367
R2199 B.n756 B.n75 163.367
R2200 B.n756 B.n755 163.367
R2201 B.n755 B.n754 163.367
R2202 B.n754 B.n77 163.367
R2203 B.n750 B.n77 163.367
R2204 B.n750 B.n749 163.367
R2205 B.n749 B.n748 163.367
R2206 B.n748 B.n79 163.367
R2207 B.n744 B.n79 163.367
R2208 B.n744 B.n743 163.367
R2209 B.n743 B.n742 163.367
R2210 B.n742 B.n81 163.367
R2211 B.n738 B.n81 163.367
R2212 B.n738 B.n737 163.367
R2213 B.n737 B.n736 163.367
R2214 B.n736 B.n83 163.367
R2215 B.n732 B.n83 163.367
R2216 B.n732 B.n731 163.367
R2217 B.n731 B.n730 163.367
R2218 B.n730 B.n85 163.367
R2219 B.n726 B.n85 163.367
R2220 B.n726 B.n725 163.367
R2221 B.n725 B.n724 163.367
R2222 B.n724 B.n87 163.367
R2223 B.n720 B.n87 163.367
R2224 B.n720 B.n719 163.367
R2225 B.n719 B.n718 163.367
R2226 B.n718 B.n89 163.367
R2227 B.n714 B.n89 163.367
R2228 B.n714 B.n713 163.367
R2229 B.n713 B.n712 163.367
R2230 B.n712 B.n91 163.367
R2231 B.n185 B.n184 66.1338
R2232 B.n191 B.n190 66.1338
R2233 B.n61 B.n60 66.1338
R2234 B.n67 B.n66 66.1338
R2235 B.n434 B.n185 59.5399
R2236 B.n192 B.n191 59.5399
R2237 B.n794 B.n61 59.5399
R2238 B.n68 B.n67 59.5399
R2239 B.n865 B.n36 34.1859
R2240 B.n710 B.n709 34.1859
R2241 B.n505 B.n160 34.1859
R2242 B.n350 B.n349 34.1859
R2243 B B.n967 18.0485
R2244 B.n861 B.n36 10.6151
R2245 B.n861 B.n860 10.6151
R2246 B.n860 B.n859 10.6151
R2247 B.n859 B.n38 10.6151
R2248 B.n855 B.n38 10.6151
R2249 B.n855 B.n854 10.6151
R2250 B.n854 B.n853 10.6151
R2251 B.n853 B.n40 10.6151
R2252 B.n849 B.n40 10.6151
R2253 B.n849 B.n848 10.6151
R2254 B.n848 B.n847 10.6151
R2255 B.n847 B.n42 10.6151
R2256 B.n843 B.n42 10.6151
R2257 B.n843 B.n842 10.6151
R2258 B.n842 B.n841 10.6151
R2259 B.n841 B.n44 10.6151
R2260 B.n837 B.n44 10.6151
R2261 B.n837 B.n836 10.6151
R2262 B.n836 B.n835 10.6151
R2263 B.n835 B.n46 10.6151
R2264 B.n831 B.n46 10.6151
R2265 B.n831 B.n830 10.6151
R2266 B.n830 B.n829 10.6151
R2267 B.n829 B.n48 10.6151
R2268 B.n825 B.n48 10.6151
R2269 B.n825 B.n824 10.6151
R2270 B.n824 B.n823 10.6151
R2271 B.n823 B.n50 10.6151
R2272 B.n819 B.n50 10.6151
R2273 B.n819 B.n818 10.6151
R2274 B.n818 B.n817 10.6151
R2275 B.n817 B.n52 10.6151
R2276 B.n813 B.n52 10.6151
R2277 B.n813 B.n812 10.6151
R2278 B.n812 B.n811 10.6151
R2279 B.n811 B.n54 10.6151
R2280 B.n807 B.n54 10.6151
R2281 B.n807 B.n806 10.6151
R2282 B.n806 B.n805 10.6151
R2283 B.n805 B.n56 10.6151
R2284 B.n801 B.n56 10.6151
R2285 B.n801 B.n800 10.6151
R2286 B.n800 B.n799 10.6151
R2287 B.n799 B.n58 10.6151
R2288 B.n795 B.n58 10.6151
R2289 B.n793 B.n792 10.6151
R2290 B.n792 B.n62 10.6151
R2291 B.n788 B.n62 10.6151
R2292 B.n788 B.n787 10.6151
R2293 B.n787 B.n786 10.6151
R2294 B.n786 B.n64 10.6151
R2295 B.n782 B.n64 10.6151
R2296 B.n782 B.n781 10.6151
R2297 B.n781 B.n780 10.6151
R2298 B.n777 B.n776 10.6151
R2299 B.n776 B.n775 10.6151
R2300 B.n775 B.n70 10.6151
R2301 B.n771 B.n70 10.6151
R2302 B.n771 B.n770 10.6151
R2303 B.n770 B.n769 10.6151
R2304 B.n769 B.n72 10.6151
R2305 B.n765 B.n72 10.6151
R2306 B.n765 B.n764 10.6151
R2307 B.n764 B.n763 10.6151
R2308 B.n763 B.n74 10.6151
R2309 B.n759 B.n74 10.6151
R2310 B.n759 B.n758 10.6151
R2311 B.n758 B.n757 10.6151
R2312 B.n757 B.n76 10.6151
R2313 B.n753 B.n76 10.6151
R2314 B.n753 B.n752 10.6151
R2315 B.n752 B.n751 10.6151
R2316 B.n751 B.n78 10.6151
R2317 B.n747 B.n78 10.6151
R2318 B.n747 B.n746 10.6151
R2319 B.n746 B.n745 10.6151
R2320 B.n745 B.n80 10.6151
R2321 B.n741 B.n80 10.6151
R2322 B.n741 B.n740 10.6151
R2323 B.n740 B.n739 10.6151
R2324 B.n739 B.n82 10.6151
R2325 B.n735 B.n82 10.6151
R2326 B.n735 B.n734 10.6151
R2327 B.n734 B.n733 10.6151
R2328 B.n733 B.n84 10.6151
R2329 B.n729 B.n84 10.6151
R2330 B.n729 B.n728 10.6151
R2331 B.n728 B.n727 10.6151
R2332 B.n727 B.n86 10.6151
R2333 B.n723 B.n86 10.6151
R2334 B.n723 B.n722 10.6151
R2335 B.n722 B.n721 10.6151
R2336 B.n721 B.n88 10.6151
R2337 B.n717 B.n88 10.6151
R2338 B.n717 B.n716 10.6151
R2339 B.n716 B.n715 10.6151
R2340 B.n715 B.n90 10.6151
R2341 B.n711 B.n90 10.6151
R2342 B.n711 B.n710 10.6151
R2343 B.n506 B.n505 10.6151
R2344 B.n507 B.n506 10.6151
R2345 B.n507 B.n158 10.6151
R2346 B.n511 B.n158 10.6151
R2347 B.n512 B.n511 10.6151
R2348 B.n513 B.n512 10.6151
R2349 B.n513 B.n156 10.6151
R2350 B.n517 B.n156 10.6151
R2351 B.n518 B.n517 10.6151
R2352 B.n519 B.n518 10.6151
R2353 B.n519 B.n154 10.6151
R2354 B.n523 B.n154 10.6151
R2355 B.n524 B.n523 10.6151
R2356 B.n525 B.n524 10.6151
R2357 B.n525 B.n152 10.6151
R2358 B.n529 B.n152 10.6151
R2359 B.n530 B.n529 10.6151
R2360 B.n531 B.n530 10.6151
R2361 B.n531 B.n150 10.6151
R2362 B.n535 B.n150 10.6151
R2363 B.n536 B.n535 10.6151
R2364 B.n537 B.n536 10.6151
R2365 B.n537 B.n148 10.6151
R2366 B.n541 B.n148 10.6151
R2367 B.n542 B.n541 10.6151
R2368 B.n543 B.n542 10.6151
R2369 B.n543 B.n146 10.6151
R2370 B.n547 B.n146 10.6151
R2371 B.n548 B.n547 10.6151
R2372 B.n549 B.n548 10.6151
R2373 B.n549 B.n144 10.6151
R2374 B.n553 B.n144 10.6151
R2375 B.n554 B.n553 10.6151
R2376 B.n555 B.n554 10.6151
R2377 B.n555 B.n142 10.6151
R2378 B.n559 B.n142 10.6151
R2379 B.n560 B.n559 10.6151
R2380 B.n561 B.n560 10.6151
R2381 B.n561 B.n140 10.6151
R2382 B.n565 B.n140 10.6151
R2383 B.n566 B.n565 10.6151
R2384 B.n567 B.n566 10.6151
R2385 B.n567 B.n138 10.6151
R2386 B.n571 B.n138 10.6151
R2387 B.n572 B.n571 10.6151
R2388 B.n573 B.n572 10.6151
R2389 B.n573 B.n136 10.6151
R2390 B.n577 B.n136 10.6151
R2391 B.n578 B.n577 10.6151
R2392 B.n579 B.n578 10.6151
R2393 B.n579 B.n134 10.6151
R2394 B.n583 B.n134 10.6151
R2395 B.n584 B.n583 10.6151
R2396 B.n585 B.n584 10.6151
R2397 B.n585 B.n132 10.6151
R2398 B.n589 B.n132 10.6151
R2399 B.n590 B.n589 10.6151
R2400 B.n591 B.n590 10.6151
R2401 B.n591 B.n130 10.6151
R2402 B.n595 B.n130 10.6151
R2403 B.n596 B.n595 10.6151
R2404 B.n597 B.n596 10.6151
R2405 B.n597 B.n128 10.6151
R2406 B.n601 B.n128 10.6151
R2407 B.n602 B.n601 10.6151
R2408 B.n603 B.n602 10.6151
R2409 B.n603 B.n126 10.6151
R2410 B.n607 B.n126 10.6151
R2411 B.n608 B.n607 10.6151
R2412 B.n609 B.n608 10.6151
R2413 B.n609 B.n124 10.6151
R2414 B.n613 B.n124 10.6151
R2415 B.n614 B.n613 10.6151
R2416 B.n615 B.n614 10.6151
R2417 B.n615 B.n122 10.6151
R2418 B.n619 B.n122 10.6151
R2419 B.n620 B.n619 10.6151
R2420 B.n621 B.n620 10.6151
R2421 B.n621 B.n120 10.6151
R2422 B.n625 B.n120 10.6151
R2423 B.n626 B.n625 10.6151
R2424 B.n627 B.n626 10.6151
R2425 B.n627 B.n118 10.6151
R2426 B.n631 B.n118 10.6151
R2427 B.n632 B.n631 10.6151
R2428 B.n633 B.n632 10.6151
R2429 B.n633 B.n116 10.6151
R2430 B.n637 B.n116 10.6151
R2431 B.n638 B.n637 10.6151
R2432 B.n639 B.n638 10.6151
R2433 B.n639 B.n114 10.6151
R2434 B.n643 B.n114 10.6151
R2435 B.n644 B.n643 10.6151
R2436 B.n645 B.n644 10.6151
R2437 B.n645 B.n112 10.6151
R2438 B.n649 B.n112 10.6151
R2439 B.n650 B.n649 10.6151
R2440 B.n651 B.n650 10.6151
R2441 B.n651 B.n110 10.6151
R2442 B.n655 B.n110 10.6151
R2443 B.n656 B.n655 10.6151
R2444 B.n657 B.n656 10.6151
R2445 B.n657 B.n108 10.6151
R2446 B.n661 B.n108 10.6151
R2447 B.n662 B.n661 10.6151
R2448 B.n663 B.n662 10.6151
R2449 B.n663 B.n106 10.6151
R2450 B.n667 B.n106 10.6151
R2451 B.n668 B.n667 10.6151
R2452 B.n669 B.n668 10.6151
R2453 B.n669 B.n104 10.6151
R2454 B.n673 B.n104 10.6151
R2455 B.n674 B.n673 10.6151
R2456 B.n675 B.n674 10.6151
R2457 B.n675 B.n102 10.6151
R2458 B.n679 B.n102 10.6151
R2459 B.n680 B.n679 10.6151
R2460 B.n681 B.n680 10.6151
R2461 B.n681 B.n100 10.6151
R2462 B.n685 B.n100 10.6151
R2463 B.n686 B.n685 10.6151
R2464 B.n687 B.n686 10.6151
R2465 B.n687 B.n98 10.6151
R2466 B.n691 B.n98 10.6151
R2467 B.n692 B.n691 10.6151
R2468 B.n693 B.n692 10.6151
R2469 B.n693 B.n96 10.6151
R2470 B.n697 B.n96 10.6151
R2471 B.n698 B.n697 10.6151
R2472 B.n699 B.n698 10.6151
R2473 B.n699 B.n94 10.6151
R2474 B.n703 B.n94 10.6151
R2475 B.n704 B.n703 10.6151
R2476 B.n705 B.n704 10.6151
R2477 B.n705 B.n92 10.6151
R2478 B.n709 B.n92 10.6151
R2479 B.n351 B.n350 10.6151
R2480 B.n351 B.n214 10.6151
R2481 B.n355 B.n214 10.6151
R2482 B.n356 B.n355 10.6151
R2483 B.n357 B.n356 10.6151
R2484 B.n357 B.n212 10.6151
R2485 B.n361 B.n212 10.6151
R2486 B.n362 B.n361 10.6151
R2487 B.n363 B.n362 10.6151
R2488 B.n363 B.n210 10.6151
R2489 B.n367 B.n210 10.6151
R2490 B.n368 B.n367 10.6151
R2491 B.n369 B.n368 10.6151
R2492 B.n369 B.n208 10.6151
R2493 B.n373 B.n208 10.6151
R2494 B.n374 B.n373 10.6151
R2495 B.n375 B.n374 10.6151
R2496 B.n375 B.n206 10.6151
R2497 B.n379 B.n206 10.6151
R2498 B.n380 B.n379 10.6151
R2499 B.n381 B.n380 10.6151
R2500 B.n381 B.n204 10.6151
R2501 B.n385 B.n204 10.6151
R2502 B.n386 B.n385 10.6151
R2503 B.n387 B.n386 10.6151
R2504 B.n387 B.n202 10.6151
R2505 B.n391 B.n202 10.6151
R2506 B.n392 B.n391 10.6151
R2507 B.n393 B.n392 10.6151
R2508 B.n393 B.n200 10.6151
R2509 B.n397 B.n200 10.6151
R2510 B.n398 B.n397 10.6151
R2511 B.n399 B.n398 10.6151
R2512 B.n399 B.n198 10.6151
R2513 B.n403 B.n198 10.6151
R2514 B.n404 B.n403 10.6151
R2515 B.n405 B.n404 10.6151
R2516 B.n405 B.n196 10.6151
R2517 B.n409 B.n196 10.6151
R2518 B.n410 B.n409 10.6151
R2519 B.n411 B.n410 10.6151
R2520 B.n411 B.n194 10.6151
R2521 B.n415 B.n194 10.6151
R2522 B.n416 B.n415 10.6151
R2523 B.n417 B.n416 10.6151
R2524 B.n421 B.n420 10.6151
R2525 B.n422 B.n421 10.6151
R2526 B.n422 B.n188 10.6151
R2527 B.n426 B.n188 10.6151
R2528 B.n427 B.n426 10.6151
R2529 B.n428 B.n427 10.6151
R2530 B.n428 B.n186 10.6151
R2531 B.n432 B.n186 10.6151
R2532 B.n433 B.n432 10.6151
R2533 B.n435 B.n182 10.6151
R2534 B.n439 B.n182 10.6151
R2535 B.n440 B.n439 10.6151
R2536 B.n441 B.n440 10.6151
R2537 B.n441 B.n180 10.6151
R2538 B.n445 B.n180 10.6151
R2539 B.n446 B.n445 10.6151
R2540 B.n447 B.n446 10.6151
R2541 B.n447 B.n178 10.6151
R2542 B.n451 B.n178 10.6151
R2543 B.n452 B.n451 10.6151
R2544 B.n453 B.n452 10.6151
R2545 B.n453 B.n176 10.6151
R2546 B.n457 B.n176 10.6151
R2547 B.n458 B.n457 10.6151
R2548 B.n459 B.n458 10.6151
R2549 B.n459 B.n174 10.6151
R2550 B.n463 B.n174 10.6151
R2551 B.n464 B.n463 10.6151
R2552 B.n465 B.n464 10.6151
R2553 B.n465 B.n172 10.6151
R2554 B.n469 B.n172 10.6151
R2555 B.n470 B.n469 10.6151
R2556 B.n471 B.n470 10.6151
R2557 B.n471 B.n170 10.6151
R2558 B.n475 B.n170 10.6151
R2559 B.n476 B.n475 10.6151
R2560 B.n477 B.n476 10.6151
R2561 B.n477 B.n168 10.6151
R2562 B.n481 B.n168 10.6151
R2563 B.n482 B.n481 10.6151
R2564 B.n483 B.n482 10.6151
R2565 B.n483 B.n166 10.6151
R2566 B.n487 B.n166 10.6151
R2567 B.n488 B.n487 10.6151
R2568 B.n489 B.n488 10.6151
R2569 B.n489 B.n164 10.6151
R2570 B.n493 B.n164 10.6151
R2571 B.n494 B.n493 10.6151
R2572 B.n495 B.n494 10.6151
R2573 B.n495 B.n162 10.6151
R2574 B.n499 B.n162 10.6151
R2575 B.n500 B.n499 10.6151
R2576 B.n501 B.n500 10.6151
R2577 B.n501 B.n160 10.6151
R2578 B.n349 B.n216 10.6151
R2579 B.n345 B.n216 10.6151
R2580 B.n345 B.n344 10.6151
R2581 B.n344 B.n343 10.6151
R2582 B.n343 B.n218 10.6151
R2583 B.n339 B.n218 10.6151
R2584 B.n339 B.n338 10.6151
R2585 B.n338 B.n337 10.6151
R2586 B.n337 B.n220 10.6151
R2587 B.n333 B.n220 10.6151
R2588 B.n333 B.n332 10.6151
R2589 B.n332 B.n331 10.6151
R2590 B.n331 B.n222 10.6151
R2591 B.n327 B.n222 10.6151
R2592 B.n327 B.n326 10.6151
R2593 B.n326 B.n325 10.6151
R2594 B.n325 B.n224 10.6151
R2595 B.n321 B.n224 10.6151
R2596 B.n321 B.n320 10.6151
R2597 B.n320 B.n319 10.6151
R2598 B.n319 B.n226 10.6151
R2599 B.n315 B.n226 10.6151
R2600 B.n315 B.n314 10.6151
R2601 B.n314 B.n313 10.6151
R2602 B.n313 B.n228 10.6151
R2603 B.n309 B.n228 10.6151
R2604 B.n309 B.n308 10.6151
R2605 B.n308 B.n307 10.6151
R2606 B.n307 B.n230 10.6151
R2607 B.n303 B.n230 10.6151
R2608 B.n303 B.n302 10.6151
R2609 B.n302 B.n301 10.6151
R2610 B.n301 B.n232 10.6151
R2611 B.n297 B.n232 10.6151
R2612 B.n297 B.n296 10.6151
R2613 B.n296 B.n295 10.6151
R2614 B.n295 B.n234 10.6151
R2615 B.n291 B.n234 10.6151
R2616 B.n291 B.n290 10.6151
R2617 B.n290 B.n289 10.6151
R2618 B.n289 B.n236 10.6151
R2619 B.n285 B.n236 10.6151
R2620 B.n285 B.n284 10.6151
R2621 B.n284 B.n283 10.6151
R2622 B.n283 B.n238 10.6151
R2623 B.n279 B.n238 10.6151
R2624 B.n279 B.n278 10.6151
R2625 B.n278 B.n277 10.6151
R2626 B.n277 B.n240 10.6151
R2627 B.n273 B.n240 10.6151
R2628 B.n273 B.n272 10.6151
R2629 B.n272 B.n271 10.6151
R2630 B.n271 B.n242 10.6151
R2631 B.n267 B.n242 10.6151
R2632 B.n267 B.n266 10.6151
R2633 B.n266 B.n265 10.6151
R2634 B.n265 B.n244 10.6151
R2635 B.n261 B.n244 10.6151
R2636 B.n261 B.n260 10.6151
R2637 B.n260 B.n259 10.6151
R2638 B.n259 B.n246 10.6151
R2639 B.n255 B.n246 10.6151
R2640 B.n255 B.n254 10.6151
R2641 B.n254 B.n253 10.6151
R2642 B.n253 B.n248 10.6151
R2643 B.n249 B.n248 10.6151
R2644 B.n249 B.n0 10.6151
R2645 B.n963 B.n1 10.6151
R2646 B.n963 B.n962 10.6151
R2647 B.n962 B.n961 10.6151
R2648 B.n961 B.n4 10.6151
R2649 B.n957 B.n4 10.6151
R2650 B.n957 B.n956 10.6151
R2651 B.n956 B.n955 10.6151
R2652 B.n955 B.n6 10.6151
R2653 B.n951 B.n6 10.6151
R2654 B.n951 B.n950 10.6151
R2655 B.n950 B.n949 10.6151
R2656 B.n949 B.n8 10.6151
R2657 B.n945 B.n8 10.6151
R2658 B.n945 B.n944 10.6151
R2659 B.n944 B.n943 10.6151
R2660 B.n943 B.n10 10.6151
R2661 B.n939 B.n10 10.6151
R2662 B.n939 B.n938 10.6151
R2663 B.n938 B.n937 10.6151
R2664 B.n937 B.n12 10.6151
R2665 B.n933 B.n12 10.6151
R2666 B.n933 B.n932 10.6151
R2667 B.n932 B.n931 10.6151
R2668 B.n931 B.n14 10.6151
R2669 B.n927 B.n14 10.6151
R2670 B.n927 B.n926 10.6151
R2671 B.n926 B.n925 10.6151
R2672 B.n925 B.n16 10.6151
R2673 B.n921 B.n16 10.6151
R2674 B.n921 B.n920 10.6151
R2675 B.n920 B.n919 10.6151
R2676 B.n919 B.n18 10.6151
R2677 B.n915 B.n18 10.6151
R2678 B.n915 B.n914 10.6151
R2679 B.n914 B.n913 10.6151
R2680 B.n913 B.n20 10.6151
R2681 B.n909 B.n20 10.6151
R2682 B.n909 B.n908 10.6151
R2683 B.n908 B.n907 10.6151
R2684 B.n907 B.n22 10.6151
R2685 B.n903 B.n22 10.6151
R2686 B.n903 B.n902 10.6151
R2687 B.n902 B.n901 10.6151
R2688 B.n901 B.n24 10.6151
R2689 B.n897 B.n24 10.6151
R2690 B.n897 B.n896 10.6151
R2691 B.n896 B.n895 10.6151
R2692 B.n895 B.n26 10.6151
R2693 B.n891 B.n26 10.6151
R2694 B.n891 B.n890 10.6151
R2695 B.n890 B.n889 10.6151
R2696 B.n889 B.n28 10.6151
R2697 B.n885 B.n28 10.6151
R2698 B.n885 B.n884 10.6151
R2699 B.n884 B.n883 10.6151
R2700 B.n883 B.n30 10.6151
R2701 B.n879 B.n30 10.6151
R2702 B.n879 B.n878 10.6151
R2703 B.n878 B.n877 10.6151
R2704 B.n877 B.n32 10.6151
R2705 B.n873 B.n32 10.6151
R2706 B.n873 B.n872 10.6151
R2707 B.n872 B.n871 10.6151
R2708 B.n871 B.n34 10.6151
R2709 B.n867 B.n34 10.6151
R2710 B.n867 B.n866 10.6151
R2711 B.n866 B.n865 10.6151
R2712 B.n795 B.n794 9.36635
R2713 B.n777 B.n68 9.36635
R2714 B.n417 B.n192 9.36635
R2715 B.n435 B.n434 9.36635
R2716 B.n967 B.n0 2.81026
R2717 B.n967 B.n1 2.81026
R2718 B.n794 B.n793 1.24928
R2719 B.n780 B.n68 1.24928
R2720 B.n420 B.n192 1.24928
R2721 B.n434 B.n433 1.24928
C0 VDD1 VDD2 2.48765f
C1 VP VTAIL 13.1274f
C2 B VP 2.5408f
C3 w_n5062_n3672# VP 11.6539f
C4 VN VTAIL 13.1132f
C5 B VN 1.42744f
C6 w_n5062_n3672# VN 10.9934f
C7 B VTAIL 4.27265f
C8 w_n5062_n3672# VTAIL 3.48926f
C9 w_n5062_n3672# B 11.780299f
C10 VDD1 VP 12.8195f
C11 VDD1 VN 0.15486f
C12 VDD2 VP 0.645324f
C13 VDD2 VN 12.3332f
C14 VDD1 VTAIL 11.2078f
C15 VDD1 B 2.78919f
C16 VDD1 w_n5062_n3672# 3.07708f
C17 VDD2 VTAIL 11.262099f
C18 VDD2 B 2.9258f
C19 VDD2 w_n5062_n3672# 3.24558f
C20 VP VN 9.38375f
C21 VDD2 VSUBS 2.3833f
C22 VDD1 VSUBS 2.195699f
C23 VTAIL VSUBS 1.472211f
C24 VN VSUBS 8.52637f
C25 VP VSUBS 4.912086f
C26 B VSUBS 6.090661f
C27 w_n5062_n3672# VSUBS 0.228337p
C28 B.n0 VSUBS 0.005507f
C29 B.n1 VSUBS 0.005507f
C30 B.n2 VSUBS 0.008709f
C31 B.n3 VSUBS 0.008709f
C32 B.n4 VSUBS 0.008709f
C33 B.n5 VSUBS 0.008709f
C34 B.n6 VSUBS 0.008709f
C35 B.n7 VSUBS 0.008709f
C36 B.n8 VSUBS 0.008709f
C37 B.n9 VSUBS 0.008709f
C38 B.n10 VSUBS 0.008709f
C39 B.n11 VSUBS 0.008709f
C40 B.n12 VSUBS 0.008709f
C41 B.n13 VSUBS 0.008709f
C42 B.n14 VSUBS 0.008709f
C43 B.n15 VSUBS 0.008709f
C44 B.n16 VSUBS 0.008709f
C45 B.n17 VSUBS 0.008709f
C46 B.n18 VSUBS 0.008709f
C47 B.n19 VSUBS 0.008709f
C48 B.n20 VSUBS 0.008709f
C49 B.n21 VSUBS 0.008709f
C50 B.n22 VSUBS 0.008709f
C51 B.n23 VSUBS 0.008709f
C52 B.n24 VSUBS 0.008709f
C53 B.n25 VSUBS 0.008709f
C54 B.n26 VSUBS 0.008709f
C55 B.n27 VSUBS 0.008709f
C56 B.n28 VSUBS 0.008709f
C57 B.n29 VSUBS 0.008709f
C58 B.n30 VSUBS 0.008709f
C59 B.n31 VSUBS 0.008709f
C60 B.n32 VSUBS 0.008709f
C61 B.n33 VSUBS 0.008709f
C62 B.n34 VSUBS 0.008709f
C63 B.n35 VSUBS 0.008709f
C64 B.n36 VSUBS 0.021808f
C65 B.n37 VSUBS 0.008709f
C66 B.n38 VSUBS 0.008709f
C67 B.n39 VSUBS 0.008709f
C68 B.n40 VSUBS 0.008709f
C69 B.n41 VSUBS 0.008709f
C70 B.n42 VSUBS 0.008709f
C71 B.n43 VSUBS 0.008709f
C72 B.n44 VSUBS 0.008709f
C73 B.n45 VSUBS 0.008709f
C74 B.n46 VSUBS 0.008709f
C75 B.n47 VSUBS 0.008709f
C76 B.n48 VSUBS 0.008709f
C77 B.n49 VSUBS 0.008709f
C78 B.n50 VSUBS 0.008709f
C79 B.n51 VSUBS 0.008709f
C80 B.n52 VSUBS 0.008709f
C81 B.n53 VSUBS 0.008709f
C82 B.n54 VSUBS 0.008709f
C83 B.n55 VSUBS 0.008709f
C84 B.n56 VSUBS 0.008709f
C85 B.n57 VSUBS 0.008709f
C86 B.n58 VSUBS 0.008709f
C87 B.n59 VSUBS 0.008709f
C88 B.t2 VSUBS 0.30543f
C89 B.t1 VSUBS 0.351778f
C90 B.t0 VSUBS 2.3693f
C91 B.n60 VSUBS 0.556789f
C92 B.n61 VSUBS 0.341293f
C93 B.n62 VSUBS 0.008709f
C94 B.n63 VSUBS 0.008709f
C95 B.n64 VSUBS 0.008709f
C96 B.n65 VSUBS 0.008709f
C97 B.t8 VSUBS 0.305434f
C98 B.t7 VSUBS 0.351782f
C99 B.t6 VSUBS 2.3693f
C100 B.n66 VSUBS 0.556786f
C101 B.n67 VSUBS 0.341289f
C102 B.n68 VSUBS 0.020178f
C103 B.n69 VSUBS 0.008709f
C104 B.n70 VSUBS 0.008709f
C105 B.n71 VSUBS 0.008709f
C106 B.n72 VSUBS 0.008709f
C107 B.n73 VSUBS 0.008709f
C108 B.n74 VSUBS 0.008709f
C109 B.n75 VSUBS 0.008709f
C110 B.n76 VSUBS 0.008709f
C111 B.n77 VSUBS 0.008709f
C112 B.n78 VSUBS 0.008709f
C113 B.n79 VSUBS 0.008709f
C114 B.n80 VSUBS 0.008709f
C115 B.n81 VSUBS 0.008709f
C116 B.n82 VSUBS 0.008709f
C117 B.n83 VSUBS 0.008709f
C118 B.n84 VSUBS 0.008709f
C119 B.n85 VSUBS 0.008709f
C120 B.n86 VSUBS 0.008709f
C121 B.n87 VSUBS 0.008709f
C122 B.n88 VSUBS 0.008709f
C123 B.n89 VSUBS 0.008709f
C124 B.n90 VSUBS 0.008709f
C125 B.n91 VSUBS 0.021808f
C126 B.n92 VSUBS 0.008709f
C127 B.n93 VSUBS 0.008709f
C128 B.n94 VSUBS 0.008709f
C129 B.n95 VSUBS 0.008709f
C130 B.n96 VSUBS 0.008709f
C131 B.n97 VSUBS 0.008709f
C132 B.n98 VSUBS 0.008709f
C133 B.n99 VSUBS 0.008709f
C134 B.n100 VSUBS 0.008709f
C135 B.n101 VSUBS 0.008709f
C136 B.n102 VSUBS 0.008709f
C137 B.n103 VSUBS 0.008709f
C138 B.n104 VSUBS 0.008709f
C139 B.n105 VSUBS 0.008709f
C140 B.n106 VSUBS 0.008709f
C141 B.n107 VSUBS 0.008709f
C142 B.n108 VSUBS 0.008709f
C143 B.n109 VSUBS 0.008709f
C144 B.n110 VSUBS 0.008709f
C145 B.n111 VSUBS 0.008709f
C146 B.n112 VSUBS 0.008709f
C147 B.n113 VSUBS 0.008709f
C148 B.n114 VSUBS 0.008709f
C149 B.n115 VSUBS 0.008709f
C150 B.n116 VSUBS 0.008709f
C151 B.n117 VSUBS 0.008709f
C152 B.n118 VSUBS 0.008709f
C153 B.n119 VSUBS 0.008709f
C154 B.n120 VSUBS 0.008709f
C155 B.n121 VSUBS 0.008709f
C156 B.n122 VSUBS 0.008709f
C157 B.n123 VSUBS 0.008709f
C158 B.n124 VSUBS 0.008709f
C159 B.n125 VSUBS 0.008709f
C160 B.n126 VSUBS 0.008709f
C161 B.n127 VSUBS 0.008709f
C162 B.n128 VSUBS 0.008709f
C163 B.n129 VSUBS 0.008709f
C164 B.n130 VSUBS 0.008709f
C165 B.n131 VSUBS 0.008709f
C166 B.n132 VSUBS 0.008709f
C167 B.n133 VSUBS 0.008709f
C168 B.n134 VSUBS 0.008709f
C169 B.n135 VSUBS 0.008709f
C170 B.n136 VSUBS 0.008709f
C171 B.n137 VSUBS 0.008709f
C172 B.n138 VSUBS 0.008709f
C173 B.n139 VSUBS 0.008709f
C174 B.n140 VSUBS 0.008709f
C175 B.n141 VSUBS 0.008709f
C176 B.n142 VSUBS 0.008709f
C177 B.n143 VSUBS 0.008709f
C178 B.n144 VSUBS 0.008709f
C179 B.n145 VSUBS 0.008709f
C180 B.n146 VSUBS 0.008709f
C181 B.n147 VSUBS 0.008709f
C182 B.n148 VSUBS 0.008709f
C183 B.n149 VSUBS 0.008709f
C184 B.n150 VSUBS 0.008709f
C185 B.n151 VSUBS 0.008709f
C186 B.n152 VSUBS 0.008709f
C187 B.n153 VSUBS 0.008709f
C188 B.n154 VSUBS 0.008709f
C189 B.n155 VSUBS 0.008709f
C190 B.n156 VSUBS 0.008709f
C191 B.n157 VSUBS 0.008709f
C192 B.n158 VSUBS 0.008709f
C193 B.n159 VSUBS 0.008709f
C194 B.n160 VSUBS 0.021808f
C195 B.n161 VSUBS 0.008709f
C196 B.n162 VSUBS 0.008709f
C197 B.n163 VSUBS 0.008709f
C198 B.n164 VSUBS 0.008709f
C199 B.n165 VSUBS 0.008709f
C200 B.n166 VSUBS 0.008709f
C201 B.n167 VSUBS 0.008709f
C202 B.n168 VSUBS 0.008709f
C203 B.n169 VSUBS 0.008709f
C204 B.n170 VSUBS 0.008709f
C205 B.n171 VSUBS 0.008709f
C206 B.n172 VSUBS 0.008709f
C207 B.n173 VSUBS 0.008709f
C208 B.n174 VSUBS 0.008709f
C209 B.n175 VSUBS 0.008709f
C210 B.n176 VSUBS 0.008709f
C211 B.n177 VSUBS 0.008709f
C212 B.n178 VSUBS 0.008709f
C213 B.n179 VSUBS 0.008709f
C214 B.n180 VSUBS 0.008709f
C215 B.n181 VSUBS 0.008709f
C216 B.n182 VSUBS 0.008709f
C217 B.n183 VSUBS 0.008709f
C218 B.t4 VSUBS 0.305434f
C219 B.t5 VSUBS 0.351782f
C220 B.t3 VSUBS 2.3693f
C221 B.n184 VSUBS 0.556786f
C222 B.n185 VSUBS 0.341289f
C223 B.n186 VSUBS 0.008709f
C224 B.n187 VSUBS 0.008709f
C225 B.n188 VSUBS 0.008709f
C226 B.n189 VSUBS 0.008709f
C227 B.t10 VSUBS 0.30543f
C228 B.t11 VSUBS 0.351778f
C229 B.t9 VSUBS 2.3693f
C230 B.n190 VSUBS 0.556789f
C231 B.n191 VSUBS 0.341293f
C232 B.n192 VSUBS 0.020178f
C233 B.n193 VSUBS 0.008709f
C234 B.n194 VSUBS 0.008709f
C235 B.n195 VSUBS 0.008709f
C236 B.n196 VSUBS 0.008709f
C237 B.n197 VSUBS 0.008709f
C238 B.n198 VSUBS 0.008709f
C239 B.n199 VSUBS 0.008709f
C240 B.n200 VSUBS 0.008709f
C241 B.n201 VSUBS 0.008709f
C242 B.n202 VSUBS 0.008709f
C243 B.n203 VSUBS 0.008709f
C244 B.n204 VSUBS 0.008709f
C245 B.n205 VSUBS 0.008709f
C246 B.n206 VSUBS 0.008709f
C247 B.n207 VSUBS 0.008709f
C248 B.n208 VSUBS 0.008709f
C249 B.n209 VSUBS 0.008709f
C250 B.n210 VSUBS 0.008709f
C251 B.n211 VSUBS 0.008709f
C252 B.n212 VSUBS 0.008709f
C253 B.n213 VSUBS 0.008709f
C254 B.n214 VSUBS 0.008709f
C255 B.n215 VSUBS 0.021808f
C256 B.n216 VSUBS 0.008709f
C257 B.n217 VSUBS 0.008709f
C258 B.n218 VSUBS 0.008709f
C259 B.n219 VSUBS 0.008709f
C260 B.n220 VSUBS 0.008709f
C261 B.n221 VSUBS 0.008709f
C262 B.n222 VSUBS 0.008709f
C263 B.n223 VSUBS 0.008709f
C264 B.n224 VSUBS 0.008709f
C265 B.n225 VSUBS 0.008709f
C266 B.n226 VSUBS 0.008709f
C267 B.n227 VSUBS 0.008709f
C268 B.n228 VSUBS 0.008709f
C269 B.n229 VSUBS 0.008709f
C270 B.n230 VSUBS 0.008709f
C271 B.n231 VSUBS 0.008709f
C272 B.n232 VSUBS 0.008709f
C273 B.n233 VSUBS 0.008709f
C274 B.n234 VSUBS 0.008709f
C275 B.n235 VSUBS 0.008709f
C276 B.n236 VSUBS 0.008709f
C277 B.n237 VSUBS 0.008709f
C278 B.n238 VSUBS 0.008709f
C279 B.n239 VSUBS 0.008709f
C280 B.n240 VSUBS 0.008709f
C281 B.n241 VSUBS 0.008709f
C282 B.n242 VSUBS 0.008709f
C283 B.n243 VSUBS 0.008709f
C284 B.n244 VSUBS 0.008709f
C285 B.n245 VSUBS 0.008709f
C286 B.n246 VSUBS 0.008709f
C287 B.n247 VSUBS 0.008709f
C288 B.n248 VSUBS 0.008709f
C289 B.n249 VSUBS 0.008709f
C290 B.n250 VSUBS 0.008709f
C291 B.n251 VSUBS 0.008709f
C292 B.n252 VSUBS 0.008709f
C293 B.n253 VSUBS 0.008709f
C294 B.n254 VSUBS 0.008709f
C295 B.n255 VSUBS 0.008709f
C296 B.n256 VSUBS 0.008709f
C297 B.n257 VSUBS 0.008709f
C298 B.n258 VSUBS 0.008709f
C299 B.n259 VSUBS 0.008709f
C300 B.n260 VSUBS 0.008709f
C301 B.n261 VSUBS 0.008709f
C302 B.n262 VSUBS 0.008709f
C303 B.n263 VSUBS 0.008709f
C304 B.n264 VSUBS 0.008709f
C305 B.n265 VSUBS 0.008709f
C306 B.n266 VSUBS 0.008709f
C307 B.n267 VSUBS 0.008709f
C308 B.n268 VSUBS 0.008709f
C309 B.n269 VSUBS 0.008709f
C310 B.n270 VSUBS 0.008709f
C311 B.n271 VSUBS 0.008709f
C312 B.n272 VSUBS 0.008709f
C313 B.n273 VSUBS 0.008709f
C314 B.n274 VSUBS 0.008709f
C315 B.n275 VSUBS 0.008709f
C316 B.n276 VSUBS 0.008709f
C317 B.n277 VSUBS 0.008709f
C318 B.n278 VSUBS 0.008709f
C319 B.n279 VSUBS 0.008709f
C320 B.n280 VSUBS 0.008709f
C321 B.n281 VSUBS 0.008709f
C322 B.n282 VSUBS 0.008709f
C323 B.n283 VSUBS 0.008709f
C324 B.n284 VSUBS 0.008709f
C325 B.n285 VSUBS 0.008709f
C326 B.n286 VSUBS 0.008709f
C327 B.n287 VSUBS 0.008709f
C328 B.n288 VSUBS 0.008709f
C329 B.n289 VSUBS 0.008709f
C330 B.n290 VSUBS 0.008709f
C331 B.n291 VSUBS 0.008709f
C332 B.n292 VSUBS 0.008709f
C333 B.n293 VSUBS 0.008709f
C334 B.n294 VSUBS 0.008709f
C335 B.n295 VSUBS 0.008709f
C336 B.n296 VSUBS 0.008709f
C337 B.n297 VSUBS 0.008709f
C338 B.n298 VSUBS 0.008709f
C339 B.n299 VSUBS 0.008709f
C340 B.n300 VSUBS 0.008709f
C341 B.n301 VSUBS 0.008709f
C342 B.n302 VSUBS 0.008709f
C343 B.n303 VSUBS 0.008709f
C344 B.n304 VSUBS 0.008709f
C345 B.n305 VSUBS 0.008709f
C346 B.n306 VSUBS 0.008709f
C347 B.n307 VSUBS 0.008709f
C348 B.n308 VSUBS 0.008709f
C349 B.n309 VSUBS 0.008709f
C350 B.n310 VSUBS 0.008709f
C351 B.n311 VSUBS 0.008709f
C352 B.n312 VSUBS 0.008709f
C353 B.n313 VSUBS 0.008709f
C354 B.n314 VSUBS 0.008709f
C355 B.n315 VSUBS 0.008709f
C356 B.n316 VSUBS 0.008709f
C357 B.n317 VSUBS 0.008709f
C358 B.n318 VSUBS 0.008709f
C359 B.n319 VSUBS 0.008709f
C360 B.n320 VSUBS 0.008709f
C361 B.n321 VSUBS 0.008709f
C362 B.n322 VSUBS 0.008709f
C363 B.n323 VSUBS 0.008709f
C364 B.n324 VSUBS 0.008709f
C365 B.n325 VSUBS 0.008709f
C366 B.n326 VSUBS 0.008709f
C367 B.n327 VSUBS 0.008709f
C368 B.n328 VSUBS 0.008709f
C369 B.n329 VSUBS 0.008709f
C370 B.n330 VSUBS 0.008709f
C371 B.n331 VSUBS 0.008709f
C372 B.n332 VSUBS 0.008709f
C373 B.n333 VSUBS 0.008709f
C374 B.n334 VSUBS 0.008709f
C375 B.n335 VSUBS 0.008709f
C376 B.n336 VSUBS 0.008709f
C377 B.n337 VSUBS 0.008709f
C378 B.n338 VSUBS 0.008709f
C379 B.n339 VSUBS 0.008709f
C380 B.n340 VSUBS 0.008709f
C381 B.n341 VSUBS 0.008709f
C382 B.n342 VSUBS 0.008709f
C383 B.n343 VSUBS 0.008709f
C384 B.n344 VSUBS 0.008709f
C385 B.n345 VSUBS 0.008709f
C386 B.n346 VSUBS 0.008709f
C387 B.n347 VSUBS 0.008709f
C388 B.n348 VSUBS 0.020201f
C389 B.n349 VSUBS 0.020201f
C390 B.n350 VSUBS 0.021808f
C391 B.n351 VSUBS 0.008709f
C392 B.n352 VSUBS 0.008709f
C393 B.n353 VSUBS 0.008709f
C394 B.n354 VSUBS 0.008709f
C395 B.n355 VSUBS 0.008709f
C396 B.n356 VSUBS 0.008709f
C397 B.n357 VSUBS 0.008709f
C398 B.n358 VSUBS 0.008709f
C399 B.n359 VSUBS 0.008709f
C400 B.n360 VSUBS 0.008709f
C401 B.n361 VSUBS 0.008709f
C402 B.n362 VSUBS 0.008709f
C403 B.n363 VSUBS 0.008709f
C404 B.n364 VSUBS 0.008709f
C405 B.n365 VSUBS 0.008709f
C406 B.n366 VSUBS 0.008709f
C407 B.n367 VSUBS 0.008709f
C408 B.n368 VSUBS 0.008709f
C409 B.n369 VSUBS 0.008709f
C410 B.n370 VSUBS 0.008709f
C411 B.n371 VSUBS 0.008709f
C412 B.n372 VSUBS 0.008709f
C413 B.n373 VSUBS 0.008709f
C414 B.n374 VSUBS 0.008709f
C415 B.n375 VSUBS 0.008709f
C416 B.n376 VSUBS 0.008709f
C417 B.n377 VSUBS 0.008709f
C418 B.n378 VSUBS 0.008709f
C419 B.n379 VSUBS 0.008709f
C420 B.n380 VSUBS 0.008709f
C421 B.n381 VSUBS 0.008709f
C422 B.n382 VSUBS 0.008709f
C423 B.n383 VSUBS 0.008709f
C424 B.n384 VSUBS 0.008709f
C425 B.n385 VSUBS 0.008709f
C426 B.n386 VSUBS 0.008709f
C427 B.n387 VSUBS 0.008709f
C428 B.n388 VSUBS 0.008709f
C429 B.n389 VSUBS 0.008709f
C430 B.n390 VSUBS 0.008709f
C431 B.n391 VSUBS 0.008709f
C432 B.n392 VSUBS 0.008709f
C433 B.n393 VSUBS 0.008709f
C434 B.n394 VSUBS 0.008709f
C435 B.n395 VSUBS 0.008709f
C436 B.n396 VSUBS 0.008709f
C437 B.n397 VSUBS 0.008709f
C438 B.n398 VSUBS 0.008709f
C439 B.n399 VSUBS 0.008709f
C440 B.n400 VSUBS 0.008709f
C441 B.n401 VSUBS 0.008709f
C442 B.n402 VSUBS 0.008709f
C443 B.n403 VSUBS 0.008709f
C444 B.n404 VSUBS 0.008709f
C445 B.n405 VSUBS 0.008709f
C446 B.n406 VSUBS 0.008709f
C447 B.n407 VSUBS 0.008709f
C448 B.n408 VSUBS 0.008709f
C449 B.n409 VSUBS 0.008709f
C450 B.n410 VSUBS 0.008709f
C451 B.n411 VSUBS 0.008709f
C452 B.n412 VSUBS 0.008709f
C453 B.n413 VSUBS 0.008709f
C454 B.n414 VSUBS 0.008709f
C455 B.n415 VSUBS 0.008709f
C456 B.n416 VSUBS 0.008709f
C457 B.n417 VSUBS 0.008197f
C458 B.n418 VSUBS 0.008709f
C459 B.n419 VSUBS 0.008709f
C460 B.n420 VSUBS 0.004867f
C461 B.n421 VSUBS 0.008709f
C462 B.n422 VSUBS 0.008709f
C463 B.n423 VSUBS 0.008709f
C464 B.n424 VSUBS 0.008709f
C465 B.n425 VSUBS 0.008709f
C466 B.n426 VSUBS 0.008709f
C467 B.n427 VSUBS 0.008709f
C468 B.n428 VSUBS 0.008709f
C469 B.n429 VSUBS 0.008709f
C470 B.n430 VSUBS 0.008709f
C471 B.n431 VSUBS 0.008709f
C472 B.n432 VSUBS 0.008709f
C473 B.n433 VSUBS 0.004867f
C474 B.n434 VSUBS 0.020178f
C475 B.n435 VSUBS 0.008197f
C476 B.n436 VSUBS 0.008709f
C477 B.n437 VSUBS 0.008709f
C478 B.n438 VSUBS 0.008709f
C479 B.n439 VSUBS 0.008709f
C480 B.n440 VSUBS 0.008709f
C481 B.n441 VSUBS 0.008709f
C482 B.n442 VSUBS 0.008709f
C483 B.n443 VSUBS 0.008709f
C484 B.n444 VSUBS 0.008709f
C485 B.n445 VSUBS 0.008709f
C486 B.n446 VSUBS 0.008709f
C487 B.n447 VSUBS 0.008709f
C488 B.n448 VSUBS 0.008709f
C489 B.n449 VSUBS 0.008709f
C490 B.n450 VSUBS 0.008709f
C491 B.n451 VSUBS 0.008709f
C492 B.n452 VSUBS 0.008709f
C493 B.n453 VSUBS 0.008709f
C494 B.n454 VSUBS 0.008709f
C495 B.n455 VSUBS 0.008709f
C496 B.n456 VSUBS 0.008709f
C497 B.n457 VSUBS 0.008709f
C498 B.n458 VSUBS 0.008709f
C499 B.n459 VSUBS 0.008709f
C500 B.n460 VSUBS 0.008709f
C501 B.n461 VSUBS 0.008709f
C502 B.n462 VSUBS 0.008709f
C503 B.n463 VSUBS 0.008709f
C504 B.n464 VSUBS 0.008709f
C505 B.n465 VSUBS 0.008709f
C506 B.n466 VSUBS 0.008709f
C507 B.n467 VSUBS 0.008709f
C508 B.n468 VSUBS 0.008709f
C509 B.n469 VSUBS 0.008709f
C510 B.n470 VSUBS 0.008709f
C511 B.n471 VSUBS 0.008709f
C512 B.n472 VSUBS 0.008709f
C513 B.n473 VSUBS 0.008709f
C514 B.n474 VSUBS 0.008709f
C515 B.n475 VSUBS 0.008709f
C516 B.n476 VSUBS 0.008709f
C517 B.n477 VSUBS 0.008709f
C518 B.n478 VSUBS 0.008709f
C519 B.n479 VSUBS 0.008709f
C520 B.n480 VSUBS 0.008709f
C521 B.n481 VSUBS 0.008709f
C522 B.n482 VSUBS 0.008709f
C523 B.n483 VSUBS 0.008709f
C524 B.n484 VSUBS 0.008709f
C525 B.n485 VSUBS 0.008709f
C526 B.n486 VSUBS 0.008709f
C527 B.n487 VSUBS 0.008709f
C528 B.n488 VSUBS 0.008709f
C529 B.n489 VSUBS 0.008709f
C530 B.n490 VSUBS 0.008709f
C531 B.n491 VSUBS 0.008709f
C532 B.n492 VSUBS 0.008709f
C533 B.n493 VSUBS 0.008709f
C534 B.n494 VSUBS 0.008709f
C535 B.n495 VSUBS 0.008709f
C536 B.n496 VSUBS 0.008709f
C537 B.n497 VSUBS 0.008709f
C538 B.n498 VSUBS 0.008709f
C539 B.n499 VSUBS 0.008709f
C540 B.n500 VSUBS 0.008709f
C541 B.n501 VSUBS 0.008709f
C542 B.n502 VSUBS 0.008709f
C543 B.n503 VSUBS 0.021808f
C544 B.n504 VSUBS 0.020201f
C545 B.n505 VSUBS 0.020201f
C546 B.n506 VSUBS 0.008709f
C547 B.n507 VSUBS 0.008709f
C548 B.n508 VSUBS 0.008709f
C549 B.n509 VSUBS 0.008709f
C550 B.n510 VSUBS 0.008709f
C551 B.n511 VSUBS 0.008709f
C552 B.n512 VSUBS 0.008709f
C553 B.n513 VSUBS 0.008709f
C554 B.n514 VSUBS 0.008709f
C555 B.n515 VSUBS 0.008709f
C556 B.n516 VSUBS 0.008709f
C557 B.n517 VSUBS 0.008709f
C558 B.n518 VSUBS 0.008709f
C559 B.n519 VSUBS 0.008709f
C560 B.n520 VSUBS 0.008709f
C561 B.n521 VSUBS 0.008709f
C562 B.n522 VSUBS 0.008709f
C563 B.n523 VSUBS 0.008709f
C564 B.n524 VSUBS 0.008709f
C565 B.n525 VSUBS 0.008709f
C566 B.n526 VSUBS 0.008709f
C567 B.n527 VSUBS 0.008709f
C568 B.n528 VSUBS 0.008709f
C569 B.n529 VSUBS 0.008709f
C570 B.n530 VSUBS 0.008709f
C571 B.n531 VSUBS 0.008709f
C572 B.n532 VSUBS 0.008709f
C573 B.n533 VSUBS 0.008709f
C574 B.n534 VSUBS 0.008709f
C575 B.n535 VSUBS 0.008709f
C576 B.n536 VSUBS 0.008709f
C577 B.n537 VSUBS 0.008709f
C578 B.n538 VSUBS 0.008709f
C579 B.n539 VSUBS 0.008709f
C580 B.n540 VSUBS 0.008709f
C581 B.n541 VSUBS 0.008709f
C582 B.n542 VSUBS 0.008709f
C583 B.n543 VSUBS 0.008709f
C584 B.n544 VSUBS 0.008709f
C585 B.n545 VSUBS 0.008709f
C586 B.n546 VSUBS 0.008709f
C587 B.n547 VSUBS 0.008709f
C588 B.n548 VSUBS 0.008709f
C589 B.n549 VSUBS 0.008709f
C590 B.n550 VSUBS 0.008709f
C591 B.n551 VSUBS 0.008709f
C592 B.n552 VSUBS 0.008709f
C593 B.n553 VSUBS 0.008709f
C594 B.n554 VSUBS 0.008709f
C595 B.n555 VSUBS 0.008709f
C596 B.n556 VSUBS 0.008709f
C597 B.n557 VSUBS 0.008709f
C598 B.n558 VSUBS 0.008709f
C599 B.n559 VSUBS 0.008709f
C600 B.n560 VSUBS 0.008709f
C601 B.n561 VSUBS 0.008709f
C602 B.n562 VSUBS 0.008709f
C603 B.n563 VSUBS 0.008709f
C604 B.n564 VSUBS 0.008709f
C605 B.n565 VSUBS 0.008709f
C606 B.n566 VSUBS 0.008709f
C607 B.n567 VSUBS 0.008709f
C608 B.n568 VSUBS 0.008709f
C609 B.n569 VSUBS 0.008709f
C610 B.n570 VSUBS 0.008709f
C611 B.n571 VSUBS 0.008709f
C612 B.n572 VSUBS 0.008709f
C613 B.n573 VSUBS 0.008709f
C614 B.n574 VSUBS 0.008709f
C615 B.n575 VSUBS 0.008709f
C616 B.n576 VSUBS 0.008709f
C617 B.n577 VSUBS 0.008709f
C618 B.n578 VSUBS 0.008709f
C619 B.n579 VSUBS 0.008709f
C620 B.n580 VSUBS 0.008709f
C621 B.n581 VSUBS 0.008709f
C622 B.n582 VSUBS 0.008709f
C623 B.n583 VSUBS 0.008709f
C624 B.n584 VSUBS 0.008709f
C625 B.n585 VSUBS 0.008709f
C626 B.n586 VSUBS 0.008709f
C627 B.n587 VSUBS 0.008709f
C628 B.n588 VSUBS 0.008709f
C629 B.n589 VSUBS 0.008709f
C630 B.n590 VSUBS 0.008709f
C631 B.n591 VSUBS 0.008709f
C632 B.n592 VSUBS 0.008709f
C633 B.n593 VSUBS 0.008709f
C634 B.n594 VSUBS 0.008709f
C635 B.n595 VSUBS 0.008709f
C636 B.n596 VSUBS 0.008709f
C637 B.n597 VSUBS 0.008709f
C638 B.n598 VSUBS 0.008709f
C639 B.n599 VSUBS 0.008709f
C640 B.n600 VSUBS 0.008709f
C641 B.n601 VSUBS 0.008709f
C642 B.n602 VSUBS 0.008709f
C643 B.n603 VSUBS 0.008709f
C644 B.n604 VSUBS 0.008709f
C645 B.n605 VSUBS 0.008709f
C646 B.n606 VSUBS 0.008709f
C647 B.n607 VSUBS 0.008709f
C648 B.n608 VSUBS 0.008709f
C649 B.n609 VSUBS 0.008709f
C650 B.n610 VSUBS 0.008709f
C651 B.n611 VSUBS 0.008709f
C652 B.n612 VSUBS 0.008709f
C653 B.n613 VSUBS 0.008709f
C654 B.n614 VSUBS 0.008709f
C655 B.n615 VSUBS 0.008709f
C656 B.n616 VSUBS 0.008709f
C657 B.n617 VSUBS 0.008709f
C658 B.n618 VSUBS 0.008709f
C659 B.n619 VSUBS 0.008709f
C660 B.n620 VSUBS 0.008709f
C661 B.n621 VSUBS 0.008709f
C662 B.n622 VSUBS 0.008709f
C663 B.n623 VSUBS 0.008709f
C664 B.n624 VSUBS 0.008709f
C665 B.n625 VSUBS 0.008709f
C666 B.n626 VSUBS 0.008709f
C667 B.n627 VSUBS 0.008709f
C668 B.n628 VSUBS 0.008709f
C669 B.n629 VSUBS 0.008709f
C670 B.n630 VSUBS 0.008709f
C671 B.n631 VSUBS 0.008709f
C672 B.n632 VSUBS 0.008709f
C673 B.n633 VSUBS 0.008709f
C674 B.n634 VSUBS 0.008709f
C675 B.n635 VSUBS 0.008709f
C676 B.n636 VSUBS 0.008709f
C677 B.n637 VSUBS 0.008709f
C678 B.n638 VSUBS 0.008709f
C679 B.n639 VSUBS 0.008709f
C680 B.n640 VSUBS 0.008709f
C681 B.n641 VSUBS 0.008709f
C682 B.n642 VSUBS 0.008709f
C683 B.n643 VSUBS 0.008709f
C684 B.n644 VSUBS 0.008709f
C685 B.n645 VSUBS 0.008709f
C686 B.n646 VSUBS 0.008709f
C687 B.n647 VSUBS 0.008709f
C688 B.n648 VSUBS 0.008709f
C689 B.n649 VSUBS 0.008709f
C690 B.n650 VSUBS 0.008709f
C691 B.n651 VSUBS 0.008709f
C692 B.n652 VSUBS 0.008709f
C693 B.n653 VSUBS 0.008709f
C694 B.n654 VSUBS 0.008709f
C695 B.n655 VSUBS 0.008709f
C696 B.n656 VSUBS 0.008709f
C697 B.n657 VSUBS 0.008709f
C698 B.n658 VSUBS 0.008709f
C699 B.n659 VSUBS 0.008709f
C700 B.n660 VSUBS 0.008709f
C701 B.n661 VSUBS 0.008709f
C702 B.n662 VSUBS 0.008709f
C703 B.n663 VSUBS 0.008709f
C704 B.n664 VSUBS 0.008709f
C705 B.n665 VSUBS 0.008709f
C706 B.n666 VSUBS 0.008709f
C707 B.n667 VSUBS 0.008709f
C708 B.n668 VSUBS 0.008709f
C709 B.n669 VSUBS 0.008709f
C710 B.n670 VSUBS 0.008709f
C711 B.n671 VSUBS 0.008709f
C712 B.n672 VSUBS 0.008709f
C713 B.n673 VSUBS 0.008709f
C714 B.n674 VSUBS 0.008709f
C715 B.n675 VSUBS 0.008709f
C716 B.n676 VSUBS 0.008709f
C717 B.n677 VSUBS 0.008709f
C718 B.n678 VSUBS 0.008709f
C719 B.n679 VSUBS 0.008709f
C720 B.n680 VSUBS 0.008709f
C721 B.n681 VSUBS 0.008709f
C722 B.n682 VSUBS 0.008709f
C723 B.n683 VSUBS 0.008709f
C724 B.n684 VSUBS 0.008709f
C725 B.n685 VSUBS 0.008709f
C726 B.n686 VSUBS 0.008709f
C727 B.n687 VSUBS 0.008709f
C728 B.n688 VSUBS 0.008709f
C729 B.n689 VSUBS 0.008709f
C730 B.n690 VSUBS 0.008709f
C731 B.n691 VSUBS 0.008709f
C732 B.n692 VSUBS 0.008709f
C733 B.n693 VSUBS 0.008709f
C734 B.n694 VSUBS 0.008709f
C735 B.n695 VSUBS 0.008709f
C736 B.n696 VSUBS 0.008709f
C737 B.n697 VSUBS 0.008709f
C738 B.n698 VSUBS 0.008709f
C739 B.n699 VSUBS 0.008709f
C740 B.n700 VSUBS 0.008709f
C741 B.n701 VSUBS 0.008709f
C742 B.n702 VSUBS 0.008709f
C743 B.n703 VSUBS 0.008709f
C744 B.n704 VSUBS 0.008709f
C745 B.n705 VSUBS 0.008709f
C746 B.n706 VSUBS 0.008709f
C747 B.n707 VSUBS 0.008709f
C748 B.n708 VSUBS 0.020201f
C749 B.n709 VSUBS 0.021184f
C750 B.n710 VSUBS 0.020825f
C751 B.n711 VSUBS 0.008709f
C752 B.n712 VSUBS 0.008709f
C753 B.n713 VSUBS 0.008709f
C754 B.n714 VSUBS 0.008709f
C755 B.n715 VSUBS 0.008709f
C756 B.n716 VSUBS 0.008709f
C757 B.n717 VSUBS 0.008709f
C758 B.n718 VSUBS 0.008709f
C759 B.n719 VSUBS 0.008709f
C760 B.n720 VSUBS 0.008709f
C761 B.n721 VSUBS 0.008709f
C762 B.n722 VSUBS 0.008709f
C763 B.n723 VSUBS 0.008709f
C764 B.n724 VSUBS 0.008709f
C765 B.n725 VSUBS 0.008709f
C766 B.n726 VSUBS 0.008709f
C767 B.n727 VSUBS 0.008709f
C768 B.n728 VSUBS 0.008709f
C769 B.n729 VSUBS 0.008709f
C770 B.n730 VSUBS 0.008709f
C771 B.n731 VSUBS 0.008709f
C772 B.n732 VSUBS 0.008709f
C773 B.n733 VSUBS 0.008709f
C774 B.n734 VSUBS 0.008709f
C775 B.n735 VSUBS 0.008709f
C776 B.n736 VSUBS 0.008709f
C777 B.n737 VSUBS 0.008709f
C778 B.n738 VSUBS 0.008709f
C779 B.n739 VSUBS 0.008709f
C780 B.n740 VSUBS 0.008709f
C781 B.n741 VSUBS 0.008709f
C782 B.n742 VSUBS 0.008709f
C783 B.n743 VSUBS 0.008709f
C784 B.n744 VSUBS 0.008709f
C785 B.n745 VSUBS 0.008709f
C786 B.n746 VSUBS 0.008709f
C787 B.n747 VSUBS 0.008709f
C788 B.n748 VSUBS 0.008709f
C789 B.n749 VSUBS 0.008709f
C790 B.n750 VSUBS 0.008709f
C791 B.n751 VSUBS 0.008709f
C792 B.n752 VSUBS 0.008709f
C793 B.n753 VSUBS 0.008709f
C794 B.n754 VSUBS 0.008709f
C795 B.n755 VSUBS 0.008709f
C796 B.n756 VSUBS 0.008709f
C797 B.n757 VSUBS 0.008709f
C798 B.n758 VSUBS 0.008709f
C799 B.n759 VSUBS 0.008709f
C800 B.n760 VSUBS 0.008709f
C801 B.n761 VSUBS 0.008709f
C802 B.n762 VSUBS 0.008709f
C803 B.n763 VSUBS 0.008709f
C804 B.n764 VSUBS 0.008709f
C805 B.n765 VSUBS 0.008709f
C806 B.n766 VSUBS 0.008709f
C807 B.n767 VSUBS 0.008709f
C808 B.n768 VSUBS 0.008709f
C809 B.n769 VSUBS 0.008709f
C810 B.n770 VSUBS 0.008709f
C811 B.n771 VSUBS 0.008709f
C812 B.n772 VSUBS 0.008709f
C813 B.n773 VSUBS 0.008709f
C814 B.n774 VSUBS 0.008709f
C815 B.n775 VSUBS 0.008709f
C816 B.n776 VSUBS 0.008709f
C817 B.n777 VSUBS 0.008197f
C818 B.n778 VSUBS 0.008709f
C819 B.n779 VSUBS 0.008709f
C820 B.n780 VSUBS 0.004867f
C821 B.n781 VSUBS 0.008709f
C822 B.n782 VSUBS 0.008709f
C823 B.n783 VSUBS 0.008709f
C824 B.n784 VSUBS 0.008709f
C825 B.n785 VSUBS 0.008709f
C826 B.n786 VSUBS 0.008709f
C827 B.n787 VSUBS 0.008709f
C828 B.n788 VSUBS 0.008709f
C829 B.n789 VSUBS 0.008709f
C830 B.n790 VSUBS 0.008709f
C831 B.n791 VSUBS 0.008709f
C832 B.n792 VSUBS 0.008709f
C833 B.n793 VSUBS 0.004867f
C834 B.n794 VSUBS 0.020178f
C835 B.n795 VSUBS 0.008197f
C836 B.n796 VSUBS 0.008709f
C837 B.n797 VSUBS 0.008709f
C838 B.n798 VSUBS 0.008709f
C839 B.n799 VSUBS 0.008709f
C840 B.n800 VSUBS 0.008709f
C841 B.n801 VSUBS 0.008709f
C842 B.n802 VSUBS 0.008709f
C843 B.n803 VSUBS 0.008709f
C844 B.n804 VSUBS 0.008709f
C845 B.n805 VSUBS 0.008709f
C846 B.n806 VSUBS 0.008709f
C847 B.n807 VSUBS 0.008709f
C848 B.n808 VSUBS 0.008709f
C849 B.n809 VSUBS 0.008709f
C850 B.n810 VSUBS 0.008709f
C851 B.n811 VSUBS 0.008709f
C852 B.n812 VSUBS 0.008709f
C853 B.n813 VSUBS 0.008709f
C854 B.n814 VSUBS 0.008709f
C855 B.n815 VSUBS 0.008709f
C856 B.n816 VSUBS 0.008709f
C857 B.n817 VSUBS 0.008709f
C858 B.n818 VSUBS 0.008709f
C859 B.n819 VSUBS 0.008709f
C860 B.n820 VSUBS 0.008709f
C861 B.n821 VSUBS 0.008709f
C862 B.n822 VSUBS 0.008709f
C863 B.n823 VSUBS 0.008709f
C864 B.n824 VSUBS 0.008709f
C865 B.n825 VSUBS 0.008709f
C866 B.n826 VSUBS 0.008709f
C867 B.n827 VSUBS 0.008709f
C868 B.n828 VSUBS 0.008709f
C869 B.n829 VSUBS 0.008709f
C870 B.n830 VSUBS 0.008709f
C871 B.n831 VSUBS 0.008709f
C872 B.n832 VSUBS 0.008709f
C873 B.n833 VSUBS 0.008709f
C874 B.n834 VSUBS 0.008709f
C875 B.n835 VSUBS 0.008709f
C876 B.n836 VSUBS 0.008709f
C877 B.n837 VSUBS 0.008709f
C878 B.n838 VSUBS 0.008709f
C879 B.n839 VSUBS 0.008709f
C880 B.n840 VSUBS 0.008709f
C881 B.n841 VSUBS 0.008709f
C882 B.n842 VSUBS 0.008709f
C883 B.n843 VSUBS 0.008709f
C884 B.n844 VSUBS 0.008709f
C885 B.n845 VSUBS 0.008709f
C886 B.n846 VSUBS 0.008709f
C887 B.n847 VSUBS 0.008709f
C888 B.n848 VSUBS 0.008709f
C889 B.n849 VSUBS 0.008709f
C890 B.n850 VSUBS 0.008709f
C891 B.n851 VSUBS 0.008709f
C892 B.n852 VSUBS 0.008709f
C893 B.n853 VSUBS 0.008709f
C894 B.n854 VSUBS 0.008709f
C895 B.n855 VSUBS 0.008709f
C896 B.n856 VSUBS 0.008709f
C897 B.n857 VSUBS 0.008709f
C898 B.n858 VSUBS 0.008709f
C899 B.n859 VSUBS 0.008709f
C900 B.n860 VSUBS 0.008709f
C901 B.n861 VSUBS 0.008709f
C902 B.n862 VSUBS 0.008709f
C903 B.n863 VSUBS 0.021808f
C904 B.n864 VSUBS 0.020201f
C905 B.n865 VSUBS 0.020201f
C906 B.n866 VSUBS 0.008709f
C907 B.n867 VSUBS 0.008709f
C908 B.n868 VSUBS 0.008709f
C909 B.n869 VSUBS 0.008709f
C910 B.n870 VSUBS 0.008709f
C911 B.n871 VSUBS 0.008709f
C912 B.n872 VSUBS 0.008709f
C913 B.n873 VSUBS 0.008709f
C914 B.n874 VSUBS 0.008709f
C915 B.n875 VSUBS 0.008709f
C916 B.n876 VSUBS 0.008709f
C917 B.n877 VSUBS 0.008709f
C918 B.n878 VSUBS 0.008709f
C919 B.n879 VSUBS 0.008709f
C920 B.n880 VSUBS 0.008709f
C921 B.n881 VSUBS 0.008709f
C922 B.n882 VSUBS 0.008709f
C923 B.n883 VSUBS 0.008709f
C924 B.n884 VSUBS 0.008709f
C925 B.n885 VSUBS 0.008709f
C926 B.n886 VSUBS 0.008709f
C927 B.n887 VSUBS 0.008709f
C928 B.n888 VSUBS 0.008709f
C929 B.n889 VSUBS 0.008709f
C930 B.n890 VSUBS 0.008709f
C931 B.n891 VSUBS 0.008709f
C932 B.n892 VSUBS 0.008709f
C933 B.n893 VSUBS 0.008709f
C934 B.n894 VSUBS 0.008709f
C935 B.n895 VSUBS 0.008709f
C936 B.n896 VSUBS 0.008709f
C937 B.n897 VSUBS 0.008709f
C938 B.n898 VSUBS 0.008709f
C939 B.n899 VSUBS 0.008709f
C940 B.n900 VSUBS 0.008709f
C941 B.n901 VSUBS 0.008709f
C942 B.n902 VSUBS 0.008709f
C943 B.n903 VSUBS 0.008709f
C944 B.n904 VSUBS 0.008709f
C945 B.n905 VSUBS 0.008709f
C946 B.n906 VSUBS 0.008709f
C947 B.n907 VSUBS 0.008709f
C948 B.n908 VSUBS 0.008709f
C949 B.n909 VSUBS 0.008709f
C950 B.n910 VSUBS 0.008709f
C951 B.n911 VSUBS 0.008709f
C952 B.n912 VSUBS 0.008709f
C953 B.n913 VSUBS 0.008709f
C954 B.n914 VSUBS 0.008709f
C955 B.n915 VSUBS 0.008709f
C956 B.n916 VSUBS 0.008709f
C957 B.n917 VSUBS 0.008709f
C958 B.n918 VSUBS 0.008709f
C959 B.n919 VSUBS 0.008709f
C960 B.n920 VSUBS 0.008709f
C961 B.n921 VSUBS 0.008709f
C962 B.n922 VSUBS 0.008709f
C963 B.n923 VSUBS 0.008709f
C964 B.n924 VSUBS 0.008709f
C965 B.n925 VSUBS 0.008709f
C966 B.n926 VSUBS 0.008709f
C967 B.n927 VSUBS 0.008709f
C968 B.n928 VSUBS 0.008709f
C969 B.n929 VSUBS 0.008709f
C970 B.n930 VSUBS 0.008709f
C971 B.n931 VSUBS 0.008709f
C972 B.n932 VSUBS 0.008709f
C973 B.n933 VSUBS 0.008709f
C974 B.n934 VSUBS 0.008709f
C975 B.n935 VSUBS 0.008709f
C976 B.n936 VSUBS 0.008709f
C977 B.n937 VSUBS 0.008709f
C978 B.n938 VSUBS 0.008709f
C979 B.n939 VSUBS 0.008709f
C980 B.n940 VSUBS 0.008709f
C981 B.n941 VSUBS 0.008709f
C982 B.n942 VSUBS 0.008709f
C983 B.n943 VSUBS 0.008709f
C984 B.n944 VSUBS 0.008709f
C985 B.n945 VSUBS 0.008709f
C986 B.n946 VSUBS 0.008709f
C987 B.n947 VSUBS 0.008709f
C988 B.n948 VSUBS 0.008709f
C989 B.n949 VSUBS 0.008709f
C990 B.n950 VSUBS 0.008709f
C991 B.n951 VSUBS 0.008709f
C992 B.n952 VSUBS 0.008709f
C993 B.n953 VSUBS 0.008709f
C994 B.n954 VSUBS 0.008709f
C995 B.n955 VSUBS 0.008709f
C996 B.n956 VSUBS 0.008709f
C997 B.n957 VSUBS 0.008709f
C998 B.n958 VSUBS 0.008709f
C999 B.n959 VSUBS 0.008709f
C1000 B.n960 VSUBS 0.008709f
C1001 B.n961 VSUBS 0.008709f
C1002 B.n962 VSUBS 0.008709f
C1003 B.n963 VSUBS 0.008709f
C1004 B.n964 VSUBS 0.008709f
C1005 B.n965 VSUBS 0.008709f
C1006 B.n966 VSUBS 0.008709f
C1007 B.n967 VSUBS 0.019721f
C1008 VDD2.n0 VSUBS 0.033213f
C1009 VDD2.n1 VSUBS 0.029879f
C1010 VDD2.n2 VSUBS 0.016056f
C1011 VDD2.n3 VSUBS 0.03795f
C1012 VDD2.n4 VSUBS 0.017f
C1013 VDD2.n5 VSUBS 0.029879f
C1014 VDD2.n6 VSUBS 0.016056f
C1015 VDD2.n7 VSUBS 0.03795f
C1016 VDD2.n8 VSUBS 0.017f
C1017 VDD2.n9 VSUBS 0.029879f
C1018 VDD2.n10 VSUBS 0.016056f
C1019 VDD2.n11 VSUBS 0.03795f
C1020 VDD2.n12 VSUBS 0.016528f
C1021 VDD2.n13 VSUBS 0.029879f
C1022 VDD2.n14 VSUBS 0.017f
C1023 VDD2.n15 VSUBS 0.03795f
C1024 VDD2.n16 VSUBS 0.017f
C1025 VDD2.n17 VSUBS 0.029879f
C1026 VDD2.n18 VSUBS 0.016056f
C1027 VDD2.n19 VSUBS 0.03795f
C1028 VDD2.n20 VSUBS 0.017f
C1029 VDD2.n21 VSUBS 1.66707f
C1030 VDD2.n22 VSUBS 0.016056f
C1031 VDD2.t0 VSUBS 0.081929f
C1032 VDD2.n23 VSUBS 0.25585f
C1033 VDD2.n24 VSUBS 0.028548f
C1034 VDD2.n25 VSUBS 0.028463f
C1035 VDD2.n26 VSUBS 0.03795f
C1036 VDD2.n27 VSUBS 0.017f
C1037 VDD2.n28 VSUBS 0.016056f
C1038 VDD2.n29 VSUBS 0.029879f
C1039 VDD2.n30 VSUBS 0.029879f
C1040 VDD2.n31 VSUBS 0.016056f
C1041 VDD2.n32 VSUBS 0.017f
C1042 VDD2.n33 VSUBS 0.03795f
C1043 VDD2.n34 VSUBS 0.03795f
C1044 VDD2.n35 VSUBS 0.017f
C1045 VDD2.n36 VSUBS 0.016056f
C1046 VDD2.n37 VSUBS 0.029879f
C1047 VDD2.n38 VSUBS 0.029879f
C1048 VDD2.n39 VSUBS 0.016056f
C1049 VDD2.n40 VSUBS 0.016056f
C1050 VDD2.n41 VSUBS 0.017f
C1051 VDD2.n42 VSUBS 0.03795f
C1052 VDD2.n43 VSUBS 0.03795f
C1053 VDD2.n44 VSUBS 0.03795f
C1054 VDD2.n45 VSUBS 0.016528f
C1055 VDD2.n46 VSUBS 0.016056f
C1056 VDD2.n47 VSUBS 0.029879f
C1057 VDD2.n48 VSUBS 0.029879f
C1058 VDD2.n49 VSUBS 0.016056f
C1059 VDD2.n50 VSUBS 0.017f
C1060 VDD2.n51 VSUBS 0.03795f
C1061 VDD2.n52 VSUBS 0.03795f
C1062 VDD2.n53 VSUBS 0.017f
C1063 VDD2.n54 VSUBS 0.016056f
C1064 VDD2.n55 VSUBS 0.029879f
C1065 VDD2.n56 VSUBS 0.029879f
C1066 VDD2.n57 VSUBS 0.016056f
C1067 VDD2.n58 VSUBS 0.017f
C1068 VDD2.n59 VSUBS 0.03795f
C1069 VDD2.n60 VSUBS 0.03795f
C1070 VDD2.n61 VSUBS 0.017f
C1071 VDD2.n62 VSUBS 0.016056f
C1072 VDD2.n63 VSUBS 0.029879f
C1073 VDD2.n64 VSUBS 0.029879f
C1074 VDD2.n65 VSUBS 0.016056f
C1075 VDD2.n66 VSUBS 0.017f
C1076 VDD2.n67 VSUBS 0.03795f
C1077 VDD2.n68 VSUBS 0.093173f
C1078 VDD2.n69 VSUBS 0.017f
C1079 VDD2.n70 VSUBS 0.016056f
C1080 VDD2.n71 VSUBS 0.067432f
C1081 VDD2.n72 VSUBS 0.087073f
C1082 VDD2.t5 VSUBS 0.319228f
C1083 VDD2.t9 VSUBS 0.319228f
C1084 VDD2.n73 VSUBS 2.53544f
C1085 VDD2.n74 VSUBS 1.24762f
C1086 VDD2.t3 VSUBS 0.319228f
C1087 VDD2.t6 VSUBS 0.319228f
C1088 VDD2.n75 VSUBS 2.56697f
C1089 VDD2.n76 VSUBS 4.21011f
C1090 VDD2.n77 VSUBS 0.033213f
C1091 VDD2.n78 VSUBS 0.029879f
C1092 VDD2.n79 VSUBS 0.016056f
C1093 VDD2.n80 VSUBS 0.03795f
C1094 VDD2.n81 VSUBS 0.017f
C1095 VDD2.n82 VSUBS 0.029879f
C1096 VDD2.n83 VSUBS 0.016056f
C1097 VDD2.n84 VSUBS 0.03795f
C1098 VDD2.n85 VSUBS 0.017f
C1099 VDD2.n86 VSUBS 0.029879f
C1100 VDD2.n87 VSUBS 0.016056f
C1101 VDD2.n88 VSUBS 0.03795f
C1102 VDD2.n89 VSUBS 0.016528f
C1103 VDD2.n90 VSUBS 0.029879f
C1104 VDD2.n91 VSUBS 0.016528f
C1105 VDD2.n92 VSUBS 0.016056f
C1106 VDD2.n93 VSUBS 0.03795f
C1107 VDD2.n94 VSUBS 0.03795f
C1108 VDD2.n95 VSUBS 0.017f
C1109 VDD2.n96 VSUBS 0.029879f
C1110 VDD2.n97 VSUBS 0.016056f
C1111 VDD2.n98 VSUBS 0.03795f
C1112 VDD2.n99 VSUBS 0.017f
C1113 VDD2.n100 VSUBS 1.66707f
C1114 VDD2.n101 VSUBS 0.016056f
C1115 VDD2.t7 VSUBS 0.081929f
C1116 VDD2.n102 VSUBS 0.25585f
C1117 VDD2.n103 VSUBS 0.028548f
C1118 VDD2.n104 VSUBS 0.028463f
C1119 VDD2.n105 VSUBS 0.03795f
C1120 VDD2.n106 VSUBS 0.017f
C1121 VDD2.n107 VSUBS 0.016056f
C1122 VDD2.n108 VSUBS 0.029879f
C1123 VDD2.n109 VSUBS 0.029879f
C1124 VDD2.n110 VSUBS 0.016056f
C1125 VDD2.n111 VSUBS 0.017f
C1126 VDD2.n112 VSUBS 0.03795f
C1127 VDD2.n113 VSUBS 0.03795f
C1128 VDD2.n114 VSUBS 0.017f
C1129 VDD2.n115 VSUBS 0.016056f
C1130 VDD2.n116 VSUBS 0.029879f
C1131 VDD2.n117 VSUBS 0.029879f
C1132 VDD2.n118 VSUBS 0.016056f
C1133 VDD2.n119 VSUBS 0.017f
C1134 VDD2.n120 VSUBS 0.03795f
C1135 VDD2.n121 VSUBS 0.03795f
C1136 VDD2.n122 VSUBS 0.017f
C1137 VDD2.n123 VSUBS 0.016056f
C1138 VDD2.n124 VSUBS 0.029879f
C1139 VDD2.n125 VSUBS 0.029879f
C1140 VDD2.n126 VSUBS 0.016056f
C1141 VDD2.n127 VSUBS 0.017f
C1142 VDD2.n128 VSUBS 0.03795f
C1143 VDD2.n129 VSUBS 0.03795f
C1144 VDD2.n130 VSUBS 0.017f
C1145 VDD2.n131 VSUBS 0.016056f
C1146 VDD2.n132 VSUBS 0.029879f
C1147 VDD2.n133 VSUBS 0.029879f
C1148 VDD2.n134 VSUBS 0.016056f
C1149 VDD2.n135 VSUBS 0.017f
C1150 VDD2.n136 VSUBS 0.03795f
C1151 VDD2.n137 VSUBS 0.03795f
C1152 VDD2.n138 VSUBS 0.017f
C1153 VDD2.n139 VSUBS 0.016056f
C1154 VDD2.n140 VSUBS 0.029879f
C1155 VDD2.n141 VSUBS 0.029879f
C1156 VDD2.n142 VSUBS 0.016056f
C1157 VDD2.n143 VSUBS 0.017f
C1158 VDD2.n144 VSUBS 0.03795f
C1159 VDD2.n145 VSUBS 0.093173f
C1160 VDD2.n146 VSUBS 0.017f
C1161 VDD2.n147 VSUBS 0.016056f
C1162 VDD2.n148 VSUBS 0.067432f
C1163 VDD2.n149 VSUBS 0.067507f
C1164 VDD2.n150 VSUBS 3.81607f
C1165 VDD2.t2 VSUBS 0.319228f
C1166 VDD2.t8 VSUBS 0.319228f
C1167 VDD2.n151 VSUBS 2.53546f
C1168 VDD2.n152 VSUBS 0.93746f
C1169 VDD2.t4 VSUBS 0.319228f
C1170 VDD2.t1 VSUBS 0.319228f
C1171 VDD2.n153 VSUBS 2.56692f
C1172 VN.t3 VSUBS 2.83139f
C1173 VN.n0 VSUBS 1.08328f
C1174 VN.n1 VSUBS 0.024876f
C1175 VN.n2 VSUBS 0.024627f
C1176 VN.n3 VSUBS 0.024876f
C1177 VN.t6 VSUBS 2.83139f
C1178 VN.n4 VSUBS 0.990428f
C1179 VN.n5 VSUBS 0.024876f
C1180 VN.n6 VSUBS 0.033064f
C1181 VN.n7 VSUBS 0.024876f
C1182 VN.t0 VSUBS 2.83139f
C1183 VN.n8 VSUBS 0.046129f
C1184 VN.n9 VSUBS 0.024876f
C1185 VN.n10 VSUBS 0.046129f
C1186 VN.t9 VSUBS 3.10887f
C1187 VN.n11 VSUBS 1.02739f
C1188 VN.t4 VSUBS 2.83139f
C1189 VN.n12 VSUBS 1.07784f
C1190 VN.n13 VSUBS 0.04203f
C1191 VN.n14 VSUBS 0.28509f
C1192 VN.n15 VSUBS 0.024876f
C1193 VN.n16 VSUBS 0.024876f
C1194 VN.n17 VSUBS 0.039258f
C1195 VN.n18 VSUBS 0.033064f
C1196 VN.n19 VSUBS 0.046129f
C1197 VN.n20 VSUBS 0.024876f
C1198 VN.n21 VSUBS 0.024876f
C1199 VN.n22 VSUBS 0.024876f
C1200 VN.n23 VSUBS 1.01378f
C1201 VN.n24 VSUBS 0.046129f
C1202 VN.n25 VSUBS 0.046129f
C1203 VN.n26 VSUBS 0.024876f
C1204 VN.n27 VSUBS 0.024876f
C1205 VN.n28 VSUBS 0.024876f
C1206 VN.n29 VSUBS 0.039258f
C1207 VN.n30 VSUBS 0.046129f
C1208 VN.n31 VSUBS 0.04203f
C1209 VN.n32 VSUBS 0.024876f
C1210 VN.n33 VSUBS 0.024876f
C1211 VN.n34 VSUBS 0.027456f
C1212 VN.n35 VSUBS 0.046129f
C1213 VN.n36 VSUBS 0.049127f
C1214 VN.n37 VSUBS 0.024876f
C1215 VN.n38 VSUBS 0.024876f
C1216 VN.n39 VSUBS 0.024876f
C1217 VN.n40 VSUBS 0.044696f
C1218 VN.n41 VSUBS 0.046129f
C1219 VN.n42 VSUBS 0.037931f
C1220 VN.n43 VSUBS 0.040142f
C1221 VN.n44 VSUBS 0.056973f
C1222 VN.t2 VSUBS 2.83139f
C1223 VN.n45 VSUBS 1.08328f
C1224 VN.n46 VSUBS 0.024876f
C1225 VN.n47 VSUBS 0.024627f
C1226 VN.n48 VSUBS 0.024876f
C1227 VN.t7 VSUBS 2.83139f
C1228 VN.n49 VSUBS 0.990428f
C1229 VN.n50 VSUBS 0.024876f
C1230 VN.n51 VSUBS 0.033064f
C1231 VN.n52 VSUBS 0.024876f
C1232 VN.t1 VSUBS 2.83139f
C1233 VN.n53 VSUBS 0.046129f
C1234 VN.n54 VSUBS 0.024876f
C1235 VN.n55 VSUBS 0.046129f
C1236 VN.t8 VSUBS 3.10887f
C1237 VN.n56 VSUBS 1.02739f
C1238 VN.t5 VSUBS 2.83139f
C1239 VN.n57 VSUBS 1.07784f
C1240 VN.n58 VSUBS 0.04203f
C1241 VN.n59 VSUBS 0.28509f
C1242 VN.n60 VSUBS 0.024876f
C1243 VN.n61 VSUBS 0.024876f
C1244 VN.n62 VSUBS 0.039258f
C1245 VN.n63 VSUBS 0.033064f
C1246 VN.n64 VSUBS 0.046129f
C1247 VN.n65 VSUBS 0.024876f
C1248 VN.n66 VSUBS 0.024876f
C1249 VN.n67 VSUBS 0.024876f
C1250 VN.n68 VSUBS 1.01378f
C1251 VN.n69 VSUBS 0.046129f
C1252 VN.n70 VSUBS 0.046129f
C1253 VN.n71 VSUBS 0.024876f
C1254 VN.n72 VSUBS 0.024876f
C1255 VN.n73 VSUBS 0.024876f
C1256 VN.n74 VSUBS 0.039258f
C1257 VN.n75 VSUBS 0.046129f
C1258 VN.n76 VSUBS 0.04203f
C1259 VN.n77 VSUBS 0.024876f
C1260 VN.n78 VSUBS 0.024876f
C1261 VN.n79 VSUBS 0.027456f
C1262 VN.n80 VSUBS 0.046129f
C1263 VN.n81 VSUBS 0.049127f
C1264 VN.n82 VSUBS 0.024876f
C1265 VN.n83 VSUBS 0.024876f
C1266 VN.n84 VSUBS 0.024876f
C1267 VN.n85 VSUBS 0.044696f
C1268 VN.n86 VSUBS 0.046129f
C1269 VN.n87 VSUBS 0.037931f
C1270 VN.n88 VSUBS 0.040142f
C1271 VN.n89 VSUBS 1.70266f
C1272 VTAIL.t3 VSUBS 0.308047f
C1273 VTAIL.t2 VSUBS 0.308047f
C1274 VTAIL.n0 VSUBS 2.27861f
C1275 VTAIL.n1 VSUBS 1.07713f
C1276 VTAIL.n2 VSUBS 0.032049f
C1277 VTAIL.n3 VSUBS 0.028833f
C1278 VTAIL.n4 VSUBS 0.015494f
C1279 VTAIL.n5 VSUBS 0.036621f
C1280 VTAIL.n6 VSUBS 0.016405f
C1281 VTAIL.n7 VSUBS 0.028833f
C1282 VTAIL.n8 VSUBS 0.015494f
C1283 VTAIL.n9 VSUBS 0.036621f
C1284 VTAIL.n10 VSUBS 0.016405f
C1285 VTAIL.n11 VSUBS 0.028833f
C1286 VTAIL.n12 VSUBS 0.015494f
C1287 VTAIL.n13 VSUBS 0.036621f
C1288 VTAIL.n14 VSUBS 0.015949f
C1289 VTAIL.n15 VSUBS 0.028833f
C1290 VTAIL.n16 VSUBS 0.016405f
C1291 VTAIL.n17 VSUBS 0.036621f
C1292 VTAIL.n18 VSUBS 0.016405f
C1293 VTAIL.n19 VSUBS 0.028833f
C1294 VTAIL.n20 VSUBS 0.015494f
C1295 VTAIL.n21 VSUBS 0.036621f
C1296 VTAIL.n22 VSUBS 0.016405f
C1297 VTAIL.n23 VSUBS 1.60868f
C1298 VTAIL.n24 VSUBS 0.015494f
C1299 VTAIL.t17 VSUBS 0.079059f
C1300 VTAIL.n25 VSUBS 0.246889f
C1301 VTAIL.n26 VSUBS 0.027548f
C1302 VTAIL.n27 VSUBS 0.027466f
C1303 VTAIL.n28 VSUBS 0.036621f
C1304 VTAIL.n29 VSUBS 0.016405f
C1305 VTAIL.n30 VSUBS 0.015494f
C1306 VTAIL.n31 VSUBS 0.028833f
C1307 VTAIL.n32 VSUBS 0.028833f
C1308 VTAIL.n33 VSUBS 0.015494f
C1309 VTAIL.n34 VSUBS 0.016405f
C1310 VTAIL.n35 VSUBS 0.036621f
C1311 VTAIL.n36 VSUBS 0.036621f
C1312 VTAIL.n37 VSUBS 0.016405f
C1313 VTAIL.n38 VSUBS 0.015494f
C1314 VTAIL.n39 VSUBS 0.028833f
C1315 VTAIL.n40 VSUBS 0.028833f
C1316 VTAIL.n41 VSUBS 0.015494f
C1317 VTAIL.n42 VSUBS 0.015494f
C1318 VTAIL.n43 VSUBS 0.016405f
C1319 VTAIL.n44 VSUBS 0.036621f
C1320 VTAIL.n45 VSUBS 0.036621f
C1321 VTAIL.n46 VSUBS 0.036621f
C1322 VTAIL.n47 VSUBS 0.015949f
C1323 VTAIL.n48 VSUBS 0.015494f
C1324 VTAIL.n49 VSUBS 0.028833f
C1325 VTAIL.n50 VSUBS 0.028833f
C1326 VTAIL.n51 VSUBS 0.015494f
C1327 VTAIL.n52 VSUBS 0.016405f
C1328 VTAIL.n53 VSUBS 0.036621f
C1329 VTAIL.n54 VSUBS 0.036621f
C1330 VTAIL.n55 VSUBS 0.016405f
C1331 VTAIL.n56 VSUBS 0.015494f
C1332 VTAIL.n57 VSUBS 0.028833f
C1333 VTAIL.n58 VSUBS 0.028833f
C1334 VTAIL.n59 VSUBS 0.015494f
C1335 VTAIL.n60 VSUBS 0.016405f
C1336 VTAIL.n61 VSUBS 0.036621f
C1337 VTAIL.n62 VSUBS 0.036621f
C1338 VTAIL.n63 VSUBS 0.016405f
C1339 VTAIL.n64 VSUBS 0.015494f
C1340 VTAIL.n65 VSUBS 0.028833f
C1341 VTAIL.n66 VSUBS 0.028833f
C1342 VTAIL.n67 VSUBS 0.015494f
C1343 VTAIL.n68 VSUBS 0.016405f
C1344 VTAIL.n69 VSUBS 0.036621f
C1345 VTAIL.n70 VSUBS 0.08991f
C1346 VTAIL.n71 VSUBS 0.016405f
C1347 VTAIL.n72 VSUBS 0.015494f
C1348 VTAIL.n73 VSUBS 0.06507f
C1349 VTAIL.n74 VSUBS 0.045222f
C1350 VTAIL.n75 VSUBS 0.477052f
C1351 VTAIL.t10 VSUBS 0.308047f
C1352 VTAIL.t12 VSUBS 0.308047f
C1353 VTAIL.n76 VSUBS 2.27861f
C1354 VTAIL.n77 VSUBS 1.23291f
C1355 VTAIL.t13 VSUBS 0.308047f
C1356 VTAIL.t14 VSUBS 0.308047f
C1357 VTAIL.n78 VSUBS 2.27861f
C1358 VTAIL.n79 VSUBS 2.98051f
C1359 VTAIL.t4 VSUBS 0.308047f
C1360 VTAIL.t7 VSUBS 0.308047f
C1361 VTAIL.n80 VSUBS 2.27862f
C1362 VTAIL.n81 VSUBS 2.9805f
C1363 VTAIL.t5 VSUBS 0.308047f
C1364 VTAIL.t8 VSUBS 0.308047f
C1365 VTAIL.n82 VSUBS 2.27862f
C1366 VTAIL.n83 VSUBS 1.23289f
C1367 VTAIL.n84 VSUBS 0.032049f
C1368 VTAIL.n85 VSUBS 0.028833f
C1369 VTAIL.n86 VSUBS 0.015494f
C1370 VTAIL.n87 VSUBS 0.036621f
C1371 VTAIL.n88 VSUBS 0.016405f
C1372 VTAIL.n89 VSUBS 0.028833f
C1373 VTAIL.n90 VSUBS 0.015494f
C1374 VTAIL.n91 VSUBS 0.036621f
C1375 VTAIL.n92 VSUBS 0.016405f
C1376 VTAIL.n93 VSUBS 0.028833f
C1377 VTAIL.n94 VSUBS 0.015494f
C1378 VTAIL.n95 VSUBS 0.036621f
C1379 VTAIL.n96 VSUBS 0.015949f
C1380 VTAIL.n97 VSUBS 0.028833f
C1381 VTAIL.n98 VSUBS 0.015949f
C1382 VTAIL.n99 VSUBS 0.015494f
C1383 VTAIL.n100 VSUBS 0.036621f
C1384 VTAIL.n101 VSUBS 0.036621f
C1385 VTAIL.n102 VSUBS 0.016405f
C1386 VTAIL.n103 VSUBS 0.028833f
C1387 VTAIL.n104 VSUBS 0.015494f
C1388 VTAIL.n105 VSUBS 0.036621f
C1389 VTAIL.n106 VSUBS 0.016405f
C1390 VTAIL.n107 VSUBS 1.60868f
C1391 VTAIL.n108 VSUBS 0.015494f
C1392 VTAIL.t1 VSUBS 0.079059f
C1393 VTAIL.n109 VSUBS 0.246889f
C1394 VTAIL.n110 VSUBS 0.027548f
C1395 VTAIL.n111 VSUBS 0.027466f
C1396 VTAIL.n112 VSUBS 0.036621f
C1397 VTAIL.n113 VSUBS 0.016405f
C1398 VTAIL.n114 VSUBS 0.015494f
C1399 VTAIL.n115 VSUBS 0.028833f
C1400 VTAIL.n116 VSUBS 0.028833f
C1401 VTAIL.n117 VSUBS 0.015494f
C1402 VTAIL.n118 VSUBS 0.016405f
C1403 VTAIL.n119 VSUBS 0.036621f
C1404 VTAIL.n120 VSUBS 0.036621f
C1405 VTAIL.n121 VSUBS 0.016405f
C1406 VTAIL.n122 VSUBS 0.015494f
C1407 VTAIL.n123 VSUBS 0.028833f
C1408 VTAIL.n124 VSUBS 0.028833f
C1409 VTAIL.n125 VSUBS 0.015494f
C1410 VTAIL.n126 VSUBS 0.016405f
C1411 VTAIL.n127 VSUBS 0.036621f
C1412 VTAIL.n128 VSUBS 0.036621f
C1413 VTAIL.n129 VSUBS 0.016405f
C1414 VTAIL.n130 VSUBS 0.015494f
C1415 VTAIL.n131 VSUBS 0.028833f
C1416 VTAIL.n132 VSUBS 0.028833f
C1417 VTAIL.n133 VSUBS 0.015494f
C1418 VTAIL.n134 VSUBS 0.016405f
C1419 VTAIL.n135 VSUBS 0.036621f
C1420 VTAIL.n136 VSUBS 0.036621f
C1421 VTAIL.n137 VSUBS 0.016405f
C1422 VTAIL.n138 VSUBS 0.015494f
C1423 VTAIL.n139 VSUBS 0.028833f
C1424 VTAIL.n140 VSUBS 0.028833f
C1425 VTAIL.n141 VSUBS 0.015494f
C1426 VTAIL.n142 VSUBS 0.016405f
C1427 VTAIL.n143 VSUBS 0.036621f
C1428 VTAIL.n144 VSUBS 0.036621f
C1429 VTAIL.n145 VSUBS 0.016405f
C1430 VTAIL.n146 VSUBS 0.015494f
C1431 VTAIL.n147 VSUBS 0.028833f
C1432 VTAIL.n148 VSUBS 0.028833f
C1433 VTAIL.n149 VSUBS 0.015494f
C1434 VTAIL.n150 VSUBS 0.016405f
C1435 VTAIL.n151 VSUBS 0.036621f
C1436 VTAIL.n152 VSUBS 0.08991f
C1437 VTAIL.n153 VSUBS 0.016405f
C1438 VTAIL.n154 VSUBS 0.015494f
C1439 VTAIL.n155 VSUBS 0.06507f
C1440 VTAIL.n156 VSUBS 0.045222f
C1441 VTAIL.n157 VSUBS 0.477052f
C1442 VTAIL.t15 VSUBS 0.308047f
C1443 VTAIL.t18 VSUBS 0.308047f
C1444 VTAIL.n158 VSUBS 2.27862f
C1445 VTAIL.n159 VSUBS 1.13999f
C1446 VTAIL.t11 VSUBS 0.308047f
C1447 VTAIL.t16 VSUBS 0.308047f
C1448 VTAIL.n160 VSUBS 2.27862f
C1449 VTAIL.n161 VSUBS 1.23289f
C1450 VTAIL.n162 VSUBS 0.032049f
C1451 VTAIL.n163 VSUBS 0.028833f
C1452 VTAIL.n164 VSUBS 0.015494f
C1453 VTAIL.n165 VSUBS 0.036621f
C1454 VTAIL.n166 VSUBS 0.016405f
C1455 VTAIL.n167 VSUBS 0.028833f
C1456 VTAIL.n168 VSUBS 0.015494f
C1457 VTAIL.n169 VSUBS 0.036621f
C1458 VTAIL.n170 VSUBS 0.016405f
C1459 VTAIL.n171 VSUBS 0.028833f
C1460 VTAIL.n172 VSUBS 0.015494f
C1461 VTAIL.n173 VSUBS 0.036621f
C1462 VTAIL.n174 VSUBS 0.015949f
C1463 VTAIL.n175 VSUBS 0.028833f
C1464 VTAIL.n176 VSUBS 0.015949f
C1465 VTAIL.n177 VSUBS 0.015494f
C1466 VTAIL.n178 VSUBS 0.036621f
C1467 VTAIL.n179 VSUBS 0.036621f
C1468 VTAIL.n180 VSUBS 0.016405f
C1469 VTAIL.n181 VSUBS 0.028833f
C1470 VTAIL.n182 VSUBS 0.015494f
C1471 VTAIL.n183 VSUBS 0.036621f
C1472 VTAIL.n184 VSUBS 0.016405f
C1473 VTAIL.n185 VSUBS 1.60868f
C1474 VTAIL.n186 VSUBS 0.015494f
C1475 VTAIL.t9 VSUBS 0.079059f
C1476 VTAIL.n187 VSUBS 0.246889f
C1477 VTAIL.n188 VSUBS 0.027548f
C1478 VTAIL.n189 VSUBS 0.027466f
C1479 VTAIL.n190 VSUBS 0.036621f
C1480 VTAIL.n191 VSUBS 0.016405f
C1481 VTAIL.n192 VSUBS 0.015494f
C1482 VTAIL.n193 VSUBS 0.028833f
C1483 VTAIL.n194 VSUBS 0.028833f
C1484 VTAIL.n195 VSUBS 0.015494f
C1485 VTAIL.n196 VSUBS 0.016405f
C1486 VTAIL.n197 VSUBS 0.036621f
C1487 VTAIL.n198 VSUBS 0.036621f
C1488 VTAIL.n199 VSUBS 0.016405f
C1489 VTAIL.n200 VSUBS 0.015494f
C1490 VTAIL.n201 VSUBS 0.028833f
C1491 VTAIL.n202 VSUBS 0.028833f
C1492 VTAIL.n203 VSUBS 0.015494f
C1493 VTAIL.n204 VSUBS 0.016405f
C1494 VTAIL.n205 VSUBS 0.036621f
C1495 VTAIL.n206 VSUBS 0.036621f
C1496 VTAIL.n207 VSUBS 0.016405f
C1497 VTAIL.n208 VSUBS 0.015494f
C1498 VTAIL.n209 VSUBS 0.028833f
C1499 VTAIL.n210 VSUBS 0.028833f
C1500 VTAIL.n211 VSUBS 0.015494f
C1501 VTAIL.n212 VSUBS 0.016405f
C1502 VTAIL.n213 VSUBS 0.036621f
C1503 VTAIL.n214 VSUBS 0.036621f
C1504 VTAIL.n215 VSUBS 0.016405f
C1505 VTAIL.n216 VSUBS 0.015494f
C1506 VTAIL.n217 VSUBS 0.028833f
C1507 VTAIL.n218 VSUBS 0.028833f
C1508 VTAIL.n219 VSUBS 0.015494f
C1509 VTAIL.n220 VSUBS 0.016405f
C1510 VTAIL.n221 VSUBS 0.036621f
C1511 VTAIL.n222 VSUBS 0.036621f
C1512 VTAIL.n223 VSUBS 0.016405f
C1513 VTAIL.n224 VSUBS 0.015494f
C1514 VTAIL.n225 VSUBS 0.028833f
C1515 VTAIL.n226 VSUBS 0.028833f
C1516 VTAIL.n227 VSUBS 0.015494f
C1517 VTAIL.n228 VSUBS 0.016405f
C1518 VTAIL.n229 VSUBS 0.036621f
C1519 VTAIL.n230 VSUBS 0.08991f
C1520 VTAIL.n231 VSUBS 0.016405f
C1521 VTAIL.n232 VSUBS 0.015494f
C1522 VTAIL.n233 VSUBS 0.06507f
C1523 VTAIL.n234 VSUBS 0.045222f
C1524 VTAIL.n235 VSUBS 2.04445f
C1525 VTAIL.n236 VSUBS 0.032049f
C1526 VTAIL.n237 VSUBS 0.028833f
C1527 VTAIL.n238 VSUBS 0.015494f
C1528 VTAIL.n239 VSUBS 0.036621f
C1529 VTAIL.n240 VSUBS 0.016405f
C1530 VTAIL.n241 VSUBS 0.028833f
C1531 VTAIL.n242 VSUBS 0.015494f
C1532 VTAIL.n243 VSUBS 0.036621f
C1533 VTAIL.n244 VSUBS 0.016405f
C1534 VTAIL.n245 VSUBS 0.028833f
C1535 VTAIL.n246 VSUBS 0.015494f
C1536 VTAIL.n247 VSUBS 0.036621f
C1537 VTAIL.n248 VSUBS 0.015949f
C1538 VTAIL.n249 VSUBS 0.028833f
C1539 VTAIL.n250 VSUBS 0.016405f
C1540 VTAIL.n251 VSUBS 0.036621f
C1541 VTAIL.n252 VSUBS 0.016405f
C1542 VTAIL.n253 VSUBS 0.028833f
C1543 VTAIL.n254 VSUBS 0.015494f
C1544 VTAIL.n255 VSUBS 0.036621f
C1545 VTAIL.n256 VSUBS 0.016405f
C1546 VTAIL.n257 VSUBS 1.60868f
C1547 VTAIL.n258 VSUBS 0.015494f
C1548 VTAIL.t19 VSUBS 0.079059f
C1549 VTAIL.n259 VSUBS 0.246889f
C1550 VTAIL.n260 VSUBS 0.027548f
C1551 VTAIL.n261 VSUBS 0.027466f
C1552 VTAIL.n262 VSUBS 0.036621f
C1553 VTAIL.n263 VSUBS 0.016405f
C1554 VTAIL.n264 VSUBS 0.015494f
C1555 VTAIL.n265 VSUBS 0.028833f
C1556 VTAIL.n266 VSUBS 0.028833f
C1557 VTAIL.n267 VSUBS 0.015494f
C1558 VTAIL.n268 VSUBS 0.016405f
C1559 VTAIL.n269 VSUBS 0.036621f
C1560 VTAIL.n270 VSUBS 0.036621f
C1561 VTAIL.n271 VSUBS 0.016405f
C1562 VTAIL.n272 VSUBS 0.015494f
C1563 VTAIL.n273 VSUBS 0.028833f
C1564 VTAIL.n274 VSUBS 0.028833f
C1565 VTAIL.n275 VSUBS 0.015494f
C1566 VTAIL.n276 VSUBS 0.015494f
C1567 VTAIL.n277 VSUBS 0.016405f
C1568 VTAIL.n278 VSUBS 0.036621f
C1569 VTAIL.n279 VSUBS 0.036621f
C1570 VTAIL.n280 VSUBS 0.036621f
C1571 VTAIL.n281 VSUBS 0.015949f
C1572 VTAIL.n282 VSUBS 0.015494f
C1573 VTAIL.n283 VSUBS 0.028833f
C1574 VTAIL.n284 VSUBS 0.028833f
C1575 VTAIL.n285 VSUBS 0.015494f
C1576 VTAIL.n286 VSUBS 0.016405f
C1577 VTAIL.n287 VSUBS 0.036621f
C1578 VTAIL.n288 VSUBS 0.036621f
C1579 VTAIL.n289 VSUBS 0.016405f
C1580 VTAIL.n290 VSUBS 0.015494f
C1581 VTAIL.n291 VSUBS 0.028833f
C1582 VTAIL.n292 VSUBS 0.028833f
C1583 VTAIL.n293 VSUBS 0.015494f
C1584 VTAIL.n294 VSUBS 0.016405f
C1585 VTAIL.n295 VSUBS 0.036621f
C1586 VTAIL.n296 VSUBS 0.036621f
C1587 VTAIL.n297 VSUBS 0.016405f
C1588 VTAIL.n298 VSUBS 0.015494f
C1589 VTAIL.n299 VSUBS 0.028833f
C1590 VTAIL.n300 VSUBS 0.028833f
C1591 VTAIL.n301 VSUBS 0.015494f
C1592 VTAIL.n302 VSUBS 0.016405f
C1593 VTAIL.n303 VSUBS 0.036621f
C1594 VTAIL.n304 VSUBS 0.08991f
C1595 VTAIL.n305 VSUBS 0.016405f
C1596 VTAIL.n306 VSUBS 0.015494f
C1597 VTAIL.n307 VSUBS 0.06507f
C1598 VTAIL.n308 VSUBS 0.045222f
C1599 VTAIL.n309 VSUBS 2.04445f
C1600 VTAIL.t6 VSUBS 0.308047f
C1601 VTAIL.t0 VSUBS 0.308047f
C1602 VTAIL.n310 VSUBS 2.27861f
C1603 VTAIL.n311 VSUBS 1.02267f
C1604 VDD1.n0 VSUBS 0.033305f
C1605 VDD1.n1 VSUBS 0.029962f
C1606 VDD1.n2 VSUBS 0.0161f
C1607 VDD1.n3 VSUBS 0.038055f
C1608 VDD1.n4 VSUBS 0.017048f
C1609 VDD1.n5 VSUBS 0.029962f
C1610 VDD1.n6 VSUBS 0.0161f
C1611 VDD1.n7 VSUBS 0.038055f
C1612 VDD1.n8 VSUBS 0.017048f
C1613 VDD1.n9 VSUBS 0.029962f
C1614 VDD1.n10 VSUBS 0.0161f
C1615 VDD1.n11 VSUBS 0.038055f
C1616 VDD1.n12 VSUBS 0.016574f
C1617 VDD1.n13 VSUBS 0.029962f
C1618 VDD1.n14 VSUBS 0.016574f
C1619 VDD1.n15 VSUBS 0.0161f
C1620 VDD1.n16 VSUBS 0.038055f
C1621 VDD1.n17 VSUBS 0.038055f
C1622 VDD1.n18 VSUBS 0.017048f
C1623 VDD1.n19 VSUBS 0.029962f
C1624 VDD1.n20 VSUBS 0.0161f
C1625 VDD1.n21 VSUBS 0.038055f
C1626 VDD1.n22 VSUBS 0.017048f
C1627 VDD1.n23 VSUBS 1.6717f
C1628 VDD1.n24 VSUBS 0.0161f
C1629 VDD1.t4 VSUBS 0.082156f
C1630 VDD1.n25 VSUBS 0.25656f
C1631 VDD1.n26 VSUBS 0.028627f
C1632 VDD1.n27 VSUBS 0.028542f
C1633 VDD1.n28 VSUBS 0.038055f
C1634 VDD1.n29 VSUBS 0.017048f
C1635 VDD1.n30 VSUBS 0.0161f
C1636 VDD1.n31 VSUBS 0.029962f
C1637 VDD1.n32 VSUBS 0.029962f
C1638 VDD1.n33 VSUBS 0.0161f
C1639 VDD1.n34 VSUBS 0.017048f
C1640 VDD1.n35 VSUBS 0.038055f
C1641 VDD1.n36 VSUBS 0.038055f
C1642 VDD1.n37 VSUBS 0.017048f
C1643 VDD1.n38 VSUBS 0.0161f
C1644 VDD1.n39 VSUBS 0.029962f
C1645 VDD1.n40 VSUBS 0.029962f
C1646 VDD1.n41 VSUBS 0.0161f
C1647 VDD1.n42 VSUBS 0.017048f
C1648 VDD1.n43 VSUBS 0.038055f
C1649 VDD1.n44 VSUBS 0.038055f
C1650 VDD1.n45 VSUBS 0.017048f
C1651 VDD1.n46 VSUBS 0.0161f
C1652 VDD1.n47 VSUBS 0.029962f
C1653 VDD1.n48 VSUBS 0.029962f
C1654 VDD1.n49 VSUBS 0.0161f
C1655 VDD1.n50 VSUBS 0.017048f
C1656 VDD1.n51 VSUBS 0.038055f
C1657 VDD1.n52 VSUBS 0.038055f
C1658 VDD1.n53 VSUBS 0.017048f
C1659 VDD1.n54 VSUBS 0.0161f
C1660 VDD1.n55 VSUBS 0.029962f
C1661 VDD1.n56 VSUBS 0.029962f
C1662 VDD1.n57 VSUBS 0.0161f
C1663 VDD1.n58 VSUBS 0.017048f
C1664 VDD1.n59 VSUBS 0.038055f
C1665 VDD1.n60 VSUBS 0.038055f
C1666 VDD1.n61 VSUBS 0.017048f
C1667 VDD1.n62 VSUBS 0.0161f
C1668 VDD1.n63 VSUBS 0.029962f
C1669 VDD1.n64 VSUBS 0.029962f
C1670 VDD1.n65 VSUBS 0.0161f
C1671 VDD1.n66 VSUBS 0.017048f
C1672 VDD1.n67 VSUBS 0.038055f
C1673 VDD1.n68 VSUBS 0.093432f
C1674 VDD1.n69 VSUBS 0.017048f
C1675 VDD1.n70 VSUBS 0.0161f
C1676 VDD1.n71 VSUBS 0.067619f
C1677 VDD1.n72 VSUBS 0.087315f
C1678 VDD1.t2 VSUBS 0.320114f
C1679 VDD1.t1 VSUBS 0.320114f
C1680 VDD1.n73 VSUBS 2.54249f
C1681 VDD1.n74 VSUBS 1.26101f
C1682 VDD1.n75 VSUBS 0.033305f
C1683 VDD1.n76 VSUBS 0.029962f
C1684 VDD1.n77 VSUBS 0.0161f
C1685 VDD1.n78 VSUBS 0.038055f
C1686 VDD1.n79 VSUBS 0.017048f
C1687 VDD1.n80 VSUBS 0.029962f
C1688 VDD1.n81 VSUBS 0.0161f
C1689 VDD1.n82 VSUBS 0.038055f
C1690 VDD1.n83 VSUBS 0.017048f
C1691 VDD1.n84 VSUBS 0.029962f
C1692 VDD1.n85 VSUBS 0.0161f
C1693 VDD1.n86 VSUBS 0.038055f
C1694 VDD1.n87 VSUBS 0.016574f
C1695 VDD1.n88 VSUBS 0.029962f
C1696 VDD1.n89 VSUBS 0.017048f
C1697 VDD1.n90 VSUBS 0.038055f
C1698 VDD1.n91 VSUBS 0.017048f
C1699 VDD1.n92 VSUBS 0.029962f
C1700 VDD1.n93 VSUBS 0.0161f
C1701 VDD1.n94 VSUBS 0.038055f
C1702 VDD1.n95 VSUBS 0.017048f
C1703 VDD1.n96 VSUBS 1.6717f
C1704 VDD1.n97 VSUBS 0.0161f
C1705 VDD1.t9 VSUBS 0.082156f
C1706 VDD1.n98 VSUBS 0.25656f
C1707 VDD1.n99 VSUBS 0.028627f
C1708 VDD1.n100 VSUBS 0.028542f
C1709 VDD1.n101 VSUBS 0.038055f
C1710 VDD1.n102 VSUBS 0.017048f
C1711 VDD1.n103 VSUBS 0.0161f
C1712 VDD1.n104 VSUBS 0.029962f
C1713 VDD1.n105 VSUBS 0.029962f
C1714 VDD1.n106 VSUBS 0.0161f
C1715 VDD1.n107 VSUBS 0.017048f
C1716 VDD1.n108 VSUBS 0.038055f
C1717 VDD1.n109 VSUBS 0.038055f
C1718 VDD1.n110 VSUBS 0.017048f
C1719 VDD1.n111 VSUBS 0.0161f
C1720 VDD1.n112 VSUBS 0.029962f
C1721 VDD1.n113 VSUBS 0.029962f
C1722 VDD1.n114 VSUBS 0.0161f
C1723 VDD1.n115 VSUBS 0.0161f
C1724 VDD1.n116 VSUBS 0.017048f
C1725 VDD1.n117 VSUBS 0.038055f
C1726 VDD1.n118 VSUBS 0.038055f
C1727 VDD1.n119 VSUBS 0.038055f
C1728 VDD1.n120 VSUBS 0.016574f
C1729 VDD1.n121 VSUBS 0.0161f
C1730 VDD1.n122 VSUBS 0.029962f
C1731 VDD1.n123 VSUBS 0.029962f
C1732 VDD1.n124 VSUBS 0.0161f
C1733 VDD1.n125 VSUBS 0.017048f
C1734 VDD1.n126 VSUBS 0.038055f
C1735 VDD1.n127 VSUBS 0.038055f
C1736 VDD1.n128 VSUBS 0.017048f
C1737 VDD1.n129 VSUBS 0.0161f
C1738 VDD1.n130 VSUBS 0.029962f
C1739 VDD1.n131 VSUBS 0.029962f
C1740 VDD1.n132 VSUBS 0.0161f
C1741 VDD1.n133 VSUBS 0.017048f
C1742 VDD1.n134 VSUBS 0.038055f
C1743 VDD1.n135 VSUBS 0.038055f
C1744 VDD1.n136 VSUBS 0.017048f
C1745 VDD1.n137 VSUBS 0.0161f
C1746 VDD1.n138 VSUBS 0.029962f
C1747 VDD1.n139 VSUBS 0.029962f
C1748 VDD1.n140 VSUBS 0.0161f
C1749 VDD1.n141 VSUBS 0.017048f
C1750 VDD1.n142 VSUBS 0.038055f
C1751 VDD1.n143 VSUBS 0.093432f
C1752 VDD1.n144 VSUBS 0.017048f
C1753 VDD1.n145 VSUBS 0.0161f
C1754 VDD1.n146 VSUBS 0.067619f
C1755 VDD1.n147 VSUBS 0.087315f
C1756 VDD1.t3 VSUBS 0.320114f
C1757 VDD1.t0 VSUBS 0.320114f
C1758 VDD1.n148 VSUBS 2.54248f
C1759 VDD1.n149 VSUBS 1.25108f
C1760 VDD1.t8 VSUBS 0.320114f
C1761 VDD1.t7 VSUBS 0.320114f
C1762 VDD1.n150 VSUBS 2.5741f
C1763 VDD1.n151 VSUBS 4.38863f
C1764 VDD1.t6 VSUBS 0.320114f
C1765 VDD1.t5 VSUBS 0.320114f
C1766 VDD1.n152 VSUBS 2.54248f
C1767 VDD1.n153 VSUBS 4.51273f
C1768 VP.t1 VSUBS 3.06247f
C1769 VP.n0 VSUBS 1.17169f
C1770 VP.n1 VSUBS 0.026906f
C1771 VP.n2 VSUBS 0.026637f
C1772 VP.n3 VSUBS 0.026906f
C1773 VP.t6 VSUBS 3.06247f
C1774 VP.n4 VSUBS 1.07126f
C1775 VP.n5 VSUBS 0.026906f
C1776 VP.n6 VSUBS 0.035762f
C1777 VP.n7 VSUBS 0.026906f
C1778 VP.t8 VSUBS 3.06247f
C1779 VP.n8 VSUBS 0.049894f
C1780 VP.n9 VSUBS 0.026906f
C1781 VP.n10 VSUBS 0.049894f
C1782 VP.n11 VSUBS 0.026906f
C1783 VP.t4 VSUBS 3.06247f
C1784 VP.n12 VSUBS 0.053137f
C1785 VP.n13 VSUBS 0.026906f
C1786 VP.n14 VSUBS 0.041027f
C1787 VP.t9 VSUBS 3.06247f
C1788 VP.n15 VSUBS 1.17169f
C1789 VP.n16 VSUBS 0.026906f
C1790 VP.n17 VSUBS 0.026637f
C1791 VP.n18 VSUBS 0.026906f
C1792 VP.t2 VSUBS 3.06247f
C1793 VP.n19 VSUBS 1.07126f
C1794 VP.n20 VSUBS 0.026906f
C1795 VP.n21 VSUBS 0.035762f
C1796 VP.n22 VSUBS 0.026906f
C1797 VP.t7 VSUBS 3.06247f
C1798 VP.n23 VSUBS 0.049894f
C1799 VP.n24 VSUBS 0.026906f
C1800 VP.n25 VSUBS 0.049894f
C1801 VP.t3 VSUBS 3.36258f
C1802 VP.n26 VSUBS 1.11124f
C1803 VP.t0 VSUBS 3.06247f
C1804 VP.n27 VSUBS 1.1658f
C1805 VP.n28 VSUBS 0.045461f
C1806 VP.n29 VSUBS 0.308357f
C1807 VP.n30 VSUBS 0.026906f
C1808 VP.n31 VSUBS 0.026906f
C1809 VP.n32 VSUBS 0.042461f
C1810 VP.n33 VSUBS 0.035762f
C1811 VP.n34 VSUBS 0.049894f
C1812 VP.n35 VSUBS 0.026906f
C1813 VP.n36 VSUBS 0.026906f
C1814 VP.n37 VSUBS 0.026906f
C1815 VP.n38 VSUBS 1.09652f
C1816 VP.n39 VSUBS 0.049894f
C1817 VP.n40 VSUBS 0.049894f
C1818 VP.n41 VSUBS 0.026906f
C1819 VP.n42 VSUBS 0.026906f
C1820 VP.n43 VSUBS 0.026906f
C1821 VP.n44 VSUBS 0.042461f
C1822 VP.n45 VSUBS 0.049894f
C1823 VP.n46 VSUBS 0.045461f
C1824 VP.n47 VSUBS 0.026906f
C1825 VP.n48 VSUBS 0.026906f
C1826 VP.n49 VSUBS 0.029696f
C1827 VP.n50 VSUBS 0.049894f
C1828 VP.n51 VSUBS 0.053137f
C1829 VP.n52 VSUBS 0.026906f
C1830 VP.n53 VSUBS 0.026906f
C1831 VP.n54 VSUBS 0.026906f
C1832 VP.n55 VSUBS 0.048344f
C1833 VP.n56 VSUBS 0.049894f
C1834 VP.n57 VSUBS 0.041027f
C1835 VP.n58 VSUBS 0.043418f
C1836 VP.n59 VSUBS 1.83107f
C1837 VP.t5 VSUBS 3.06247f
C1838 VP.n60 VSUBS 1.17169f
C1839 VP.n61 VSUBS 1.8481f
C1840 VP.n62 VSUBS 0.043418f
C1841 VP.n63 VSUBS 0.026906f
C1842 VP.n64 VSUBS 0.049894f
C1843 VP.n65 VSUBS 0.048344f
C1844 VP.n66 VSUBS 0.026637f
C1845 VP.n67 VSUBS 0.026906f
C1846 VP.n68 VSUBS 0.026906f
C1847 VP.n69 VSUBS 0.026906f
C1848 VP.n70 VSUBS 0.049894f
C1849 VP.n71 VSUBS 0.029696f
C1850 VP.n72 VSUBS 1.07126f
C1851 VP.n73 VSUBS 0.045461f
C1852 VP.n74 VSUBS 0.026906f
C1853 VP.n75 VSUBS 0.026906f
C1854 VP.n76 VSUBS 0.026906f
C1855 VP.n77 VSUBS 0.042461f
C1856 VP.n78 VSUBS 0.035762f
C1857 VP.n79 VSUBS 0.049894f
C1858 VP.n80 VSUBS 0.026906f
C1859 VP.n81 VSUBS 0.026906f
C1860 VP.n82 VSUBS 0.026906f
C1861 VP.n83 VSUBS 1.09652f
C1862 VP.n84 VSUBS 0.049894f
C1863 VP.n85 VSUBS 0.049894f
C1864 VP.n86 VSUBS 0.026906f
C1865 VP.n87 VSUBS 0.026906f
C1866 VP.n88 VSUBS 0.026906f
C1867 VP.n89 VSUBS 0.042461f
C1868 VP.n90 VSUBS 0.049894f
C1869 VP.n91 VSUBS 0.045461f
C1870 VP.n92 VSUBS 0.026906f
C1871 VP.n93 VSUBS 0.026906f
C1872 VP.n94 VSUBS 0.029696f
C1873 VP.n95 VSUBS 0.049894f
C1874 VP.n96 VSUBS 0.053137f
C1875 VP.n97 VSUBS 0.026906f
C1876 VP.n98 VSUBS 0.026906f
C1877 VP.n99 VSUBS 0.026906f
C1878 VP.n100 VSUBS 0.048344f
C1879 VP.n101 VSUBS 0.049894f
C1880 VP.n102 VSUBS 0.041027f
C1881 VP.n103 VSUBS 0.043418f
C1882 VP.n104 VSUBS 0.061623f
.ends

