* NGSPICE file created from diff_pair_sample_1399.ext - technology: sky130A

.subckt diff_pair_sample_1399 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.35
X1 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.35
X2 VDD1.t6 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.35
X3 VDD2.t2 VN.t1 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X4 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.35
X5 VTAIL.t7 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X6 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.35
X7 VDD2.t3 VN.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.35
X8 VTAIL.t12 VN.t3 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.35
X10 VTAIL.t11 VN.t4 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.35
X11 VDD2.t0 VN.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X12 VDD1.t3 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X13 VTAIL.t9 VN.t6 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.35
X15 VTAIL.t6 VP.t5 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X16 VDD1.t1 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.35
X17 VTAIL.t5 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.35
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.35
X19 VDD2.t5 VN.t7 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.35
R0 VN.n1 VN.t0 305.515
R1 VN.n7 VN.t2 305.515
R2 VN.n4 VN.t7 289.993
R3 VN.n10 VN.t4 289.993
R4 VN.n2 VN.t1 276.118
R5 VN.n3 VN.t6 276.118
R6 VN.n8 VN.t3 276.118
R7 VN.n9 VN.t5 276.118
R8 VN.n5 VN.n4 161.3
R9 VN.n11 VN.n10 161.3
R10 VN.n9 VN.n6 161.3
R11 VN.n3 VN.n0 161.3
R12 VN.n7 VN.n6 73.1314
R13 VN.n1 VN.n0 73.1314
R14 VN.n3 VN.n2 48.2005
R15 VN.n9 VN.n8 48.2005
R16 VN.n4 VN.n3 34.3247
R17 VN.n10 VN.n9 34.3247
R18 VN VN.n11 33.5251
R19 VN.n8 VN.n7 15.5045
R20 VN.n2 VN.n1 15.5045
R21 VN.n11 VN.n6 0.189894
R22 VN.n5 VN.n0 0.189894
R23 VN VN.n5 0.0516364
R24 VDD2.n2 VDD2.n1 92.1306
R25 VDD2.n2 VDD2.n0 92.1306
R26 VDD2 VDD2.n5 92.1278
R27 VDD2.n4 VDD2.n3 91.8929
R28 VDD2.n4 VDD2.n2 28.3963
R29 VDD2.n5 VDD2.t1 8.35493
R30 VDD2.n5 VDD2.t3 8.35493
R31 VDD2.n3 VDD2.t6 8.35493
R32 VDD2.n3 VDD2.t0 8.35493
R33 VDD2.n1 VDD2.t7 8.35493
R34 VDD2.n1 VDD2.t5 8.35493
R35 VDD2.n0 VDD2.t4 8.35493
R36 VDD2.n0 VDD2.t2 8.35493
R37 VDD2 VDD2.n4 0.351793
R38 VTAIL.n14 VTAIL.t1 83.5685
R39 VTAIL.n11 VTAIL.t5 83.5685
R40 VTAIL.n10 VTAIL.t13 83.5685
R41 VTAIL.n7 VTAIL.t11 83.5685
R42 VTAIL.n15 VTAIL.t8 83.5684
R43 VTAIL.n2 VTAIL.t15 83.5684
R44 VTAIL.n3 VTAIL.t0 83.5684
R45 VTAIL.n6 VTAIL.t4 83.5684
R46 VTAIL.n13 VTAIL.n12 75.2141
R47 VTAIL.n9 VTAIL.n8 75.2141
R48 VTAIL.n1 VTAIL.n0 75.214
R49 VTAIL.n5 VTAIL.n4 75.214
R50 VTAIL.n15 VTAIL.n14 14.9962
R51 VTAIL.n7 VTAIL.n6 14.9962
R52 VTAIL.n0 VTAIL.t14 8.35493
R53 VTAIL.n0 VTAIL.t9 8.35493
R54 VTAIL.n4 VTAIL.t2 8.35493
R55 VTAIL.n4 VTAIL.t7 8.35493
R56 VTAIL.n12 VTAIL.t3 8.35493
R57 VTAIL.n12 VTAIL.t6 8.35493
R58 VTAIL.n8 VTAIL.t10 8.35493
R59 VTAIL.n8 VTAIL.t12 8.35493
R60 VTAIL.n9 VTAIL.n7 0.586707
R61 VTAIL.n10 VTAIL.n9 0.586707
R62 VTAIL.n13 VTAIL.n11 0.586707
R63 VTAIL.n14 VTAIL.n13 0.586707
R64 VTAIL.n6 VTAIL.n5 0.586707
R65 VTAIL.n5 VTAIL.n3 0.586707
R66 VTAIL.n2 VTAIL.n1 0.586707
R67 VTAIL VTAIL.n15 0.528517
R68 VTAIL.n11 VTAIL.n10 0.470328
R69 VTAIL.n3 VTAIL.n2 0.470328
R70 VTAIL VTAIL.n1 0.0586897
R71 B.n267 B.n266 585
R72 B.n269 B.n59 585
R73 B.n272 B.n271 585
R74 B.n273 B.n58 585
R75 B.n275 B.n274 585
R76 B.n277 B.n57 585
R77 B.n280 B.n279 585
R78 B.n281 B.n56 585
R79 B.n283 B.n282 585
R80 B.n285 B.n55 585
R81 B.n288 B.n287 585
R82 B.n289 B.n51 585
R83 B.n291 B.n290 585
R84 B.n293 B.n50 585
R85 B.n296 B.n295 585
R86 B.n297 B.n49 585
R87 B.n299 B.n298 585
R88 B.n301 B.n48 585
R89 B.n304 B.n303 585
R90 B.n305 B.n47 585
R91 B.n307 B.n306 585
R92 B.n309 B.n46 585
R93 B.n312 B.n311 585
R94 B.n314 B.n43 585
R95 B.n316 B.n315 585
R96 B.n318 B.n42 585
R97 B.n321 B.n320 585
R98 B.n322 B.n41 585
R99 B.n324 B.n323 585
R100 B.n326 B.n40 585
R101 B.n329 B.n328 585
R102 B.n330 B.n39 585
R103 B.n332 B.n331 585
R104 B.n334 B.n38 585
R105 B.n337 B.n336 585
R106 B.n338 B.n37 585
R107 B.n265 B.n35 585
R108 B.n341 B.n35 585
R109 B.n264 B.n34 585
R110 B.n342 B.n34 585
R111 B.n263 B.n33 585
R112 B.n343 B.n33 585
R113 B.n262 B.n261 585
R114 B.n261 B.n29 585
R115 B.n260 B.n28 585
R116 B.n349 B.n28 585
R117 B.n259 B.n27 585
R118 B.n350 B.n27 585
R119 B.n258 B.n26 585
R120 B.n351 B.n26 585
R121 B.n257 B.n256 585
R122 B.n256 B.n22 585
R123 B.n255 B.n21 585
R124 B.n357 B.n21 585
R125 B.n254 B.n20 585
R126 B.n358 B.n20 585
R127 B.n253 B.n19 585
R128 B.n359 B.n19 585
R129 B.n252 B.n251 585
R130 B.n251 B.n18 585
R131 B.n250 B.n14 585
R132 B.n365 B.n14 585
R133 B.n249 B.n13 585
R134 B.n366 B.n13 585
R135 B.n248 B.n12 585
R136 B.n367 B.n12 585
R137 B.n247 B.n246 585
R138 B.n246 B.n11 585
R139 B.n245 B.n7 585
R140 B.n373 B.n7 585
R141 B.n244 B.n6 585
R142 B.n374 B.n6 585
R143 B.n243 B.n5 585
R144 B.n375 B.n5 585
R145 B.n242 B.n241 585
R146 B.n241 B.n4 585
R147 B.n240 B.n60 585
R148 B.n240 B.n239 585
R149 B.n229 B.n61 585
R150 B.n232 B.n61 585
R151 B.n231 B.n230 585
R152 B.n233 B.n231 585
R153 B.n228 B.n65 585
R154 B.n68 B.n65 585
R155 B.n227 B.n226 585
R156 B.n226 B.n225 585
R157 B.n67 B.n66 585
R158 B.n218 B.n67 585
R159 B.n217 B.n216 585
R160 B.n219 B.n217 585
R161 B.n215 B.n72 585
R162 B.n76 B.n72 585
R163 B.n214 B.n213 585
R164 B.n213 B.n212 585
R165 B.n74 B.n73 585
R166 B.n75 B.n74 585
R167 B.n205 B.n204 585
R168 B.n206 B.n205 585
R169 B.n203 B.n81 585
R170 B.n81 B.n80 585
R171 B.n202 B.n201 585
R172 B.n201 B.n200 585
R173 B.n83 B.n82 585
R174 B.n84 B.n83 585
R175 B.n193 B.n192 585
R176 B.n194 B.n193 585
R177 B.n191 B.n89 585
R178 B.n89 B.n88 585
R179 B.n190 B.n189 585
R180 B.n189 B.n188 585
R181 B.n185 B.n93 585
R182 B.n184 B.n183 585
R183 B.n181 B.n94 585
R184 B.n181 B.n92 585
R185 B.n180 B.n179 585
R186 B.n178 B.n177 585
R187 B.n176 B.n96 585
R188 B.n174 B.n173 585
R189 B.n172 B.n97 585
R190 B.n171 B.n170 585
R191 B.n168 B.n98 585
R192 B.n166 B.n165 585
R193 B.n164 B.n99 585
R194 B.n163 B.n162 585
R195 B.n160 B.n159 585
R196 B.n158 B.n157 585
R197 B.n156 B.n104 585
R198 B.n154 B.n153 585
R199 B.n152 B.n105 585
R200 B.n151 B.n150 585
R201 B.n148 B.n106 585
R202 B.n146 B.n145 585
R203 B.n144 B.n107 585
R204 B.n143 B.n142 585
R205 B.n140 B.n139 585
R206 B.n138 B.n137 585
R207 B.n136 B.n112 585
R208 B.n134 B.n133 585
R209 B.n132 B.n113 585
R210 B.n131 B.n130 585
R211 B.n128 B.n114 585
R212 B.n126 B.n125 585
R213 B.n124 B.n115 585
R214 B.n123 B.n122 585
R215 B.n120 B.n116 585
R216 B.n118 B.n117 585
R217 B.n91 B.n90 585
R218 B.n92 B.n91 585
R219 B.n187 B.n186 585
R220 B.n188 B.n187 585
R221 B.n87 B.n86 585
R222 B.n88 B.n87 585
R223 B.n196 B.n195 585
R224 B.n195 B.n194 585
R225 B.n197 B.n85 585
R226 B.n85 B.n84 585
R227 B.n199 B.n198 585
R228 B.n200 B.n199 585
R229 B.n79 B.n78 585
R230 B.n80 B.n79 585
R231 B.n208 B.n207 585
R232 B.n207 B.n206 585
R233 B.n209 B.n77 585
R234 B.n77 B.n75 585
R235 B.n211 B.n210 585
R236 B.n212 B.n211 585
R237 B.n71 B.n70 585
R238 B.n76 B.n71 585
R239 B.n221 B.n220 585
R240 B.n220 B.n219 585
R241 B.n222 B.n69 585
R242 B.n218 B.n69 585
R243 B.n224 B.n223 585
R244 B.n225 B.n224 585
R245 B.n64 B.n63 585
R246 B.n68 B.n64 585
R247 B.n235 B.n234 585
R248 B.n234 B.n233 585
R249 B.n236 B.n62 585
R250 B.n232 B.n62 585
R251 B.n238 B.n237 585
R252 B.n239 B.n238 585
R253 B.n2 B.n0 585
R254 B.n4 B.n2 585
R255 B.n3 B.n1 585
R256 B.n374 B.n3 585
R257 B.n372 B.n371 585
R258 B.n373 B.n372 585
R259 B.n370 B.n8 585
R260 B.n11 B.n8 585
R261 B.n369 B.n368 585
R262 B.n368 B.n367 585
R263 B.n10 B.n9 585
R264 B.n366 B.n10 585
R265 B.n364 B.n363 585
R266 B.n365 B.n364 585
R267 B.n362 B.n15 585
R268 B.n18 B.n15 585
R269 B.n361 B.n360 585
R270 B.n360 B.n359 585
R271 B.n17 B.n16 585
R272 B.n358 B.n17 585
R273 B.n356 B.n355 585
R274 B.n357 B.n356 585
R275 B.n354 B.n23 585
R276 B.n23 B.n22 585
R277 B.n353 B.n352 585
R278 B.n352 B.n351 585
R279 B.n25 B.n24 585
R280 B.n350 B.n25 585
R281 B.n348 B.n347 585
R282 B.n349 B.n348 585
R283 B.n346 B.n30 585
R284 B.n30 B.n29 585
R285 B.n345 B.n344 585
R286 B.n344 B.n343 585
R287 B.n32 B.n31 585
R288 B.n342 B.n32 585
R289 B.n340 B.n339 585
R290 B.n341 B.n340 585
R291 B.n377 B.n376 585
R292 B.n376 B.n375 585
R293 B.n187 B.n93 530.939
R294 B.n340 B.n37 530.939
R295 B.n189 B.n91 530.939
R296 B.n267 B.n35 530.939
R297 B.n108 B.t12 374.764
R298 B.n100 B.t19 374.764
R299 B.n44 B.t16 374.764
R300 B.n52 B.t8 374.764
R301 B.n268 B.n36 256.663
R302 B.n270 B.n36 256.663
R303 B.n276 B.n36 256.663
R304 B.n278 B.n36 256.663
R305 B.n284 B.n36 256.663
R306 B.n286 B.n36 256.663
R307 B.n292 B.n36 256.663
R308 B.n294 B.n36 256.663
R309 B.n300 B.n36 256.663
R310 B.n302 B.n36 256.663
R311 B.n308 B.n36 256.663
R312 B.n310 B.n36 256.663
R313 B.n317 B.n36 256.663
R314 B.n319 B.n36 256.663
R315 B.n325 B.n36 256.663
R316 B.n327 B.n36 256.663
R317 B.n333 B.n36 256.663
R318 B.n335 B.n36 256.663
R319 B.n182 B.n92 256.663
R320 B.n95 B.n92 256.663
R321 B.n175 B.n92 256.663
R322 B.n169 B.n92 256.663
R323 B.n167 B.n92 256.663
R324 B.n161 B.n92 256.663
R325 B.n103 B.n92 256.663
R326 B.n155 B.n92 256.663
R327 B.n149 B.n92 256.663
R328 B.n147 B.n92 256.663
R329 B.n141 B.n92 256.663
R330 B.n111 B.n92 256.663
R331 B.n135 B.n92 256.663
R332 B.n129 B.n92 256.663
R333 B.n127 B.n92 256.663
R334 B.n121 B.n92 256.663
R335 B.n119 B.n92 256.663
R336 B.n188 B.n92 188.489
R337 B.n341 B.n36 188.489
R338 B.n187 B.n87 163.367
R339 B.n195 B.n87 163.367
R340 B.n195 B.n85 163.367
R341 B.n199 B.n85 163.367
R342 B.n199 B.n79 163.367
R343 B.n207 B.n79 163.367
R344 B.n207 B.n77 163.367
R345 B.n211 B.n77 163.367
R346 B.n211 B.n71 163.367
R347 B.n220 B.n71 163.367
R348 B.n220 B.n69 163.367
R349 B.n224 B.n69 163.367
R350 B.n224 B.n64 163.367
R351 B.n234 B.n64 163.367
R352 B.n234 B.n62 163.367
R353 B.n238 B.n62 163.367
R354 B.n238 B.n2 163.367
R355 B.n376 B.n2 163.367
R356 B.n376 B.n3 163.367
R357 B.n372 B.n3 163.367
R358 B.n372 B.n8 163.367
R359 B.n368 B.n8 163.367
R360 B.n368 B.n10 163.367
R361 B.n364 B.n10 163.367
R362 B.n364 B.n15 163.367
R363 B.n360 B.n15 163.367
R364 B.n360 B.n17 163.367
R365 B.n356 B.n17 163.367
R366 B.n356 B.n23 163.367
R367 B.n352 B.n23 163.367
R368 B.n352 B.n25 163.367
R369 B.n348 B.n25 163.367
R370 B.n348 B.n30 163.367
R371 B.n344 B.n30 163.367
R372 B.n344 B.n32 163.367
R373 B.n340 B.n32 163.367
R374 B.n183 B.n181 163.367
R375 B.n181 B.n180 163.367
R376 B.n177 B.n176 163.367
R377 B.n174 B.n97 163.367
R378 B.n170 B.n168 163.367
R379 B.n166 B.n99 163.367
R380 B.n162 B.n160 163.367
R381 B.n157 B.n156 163.367
R382 B.n154 B.n105 163.367
R383 B.n150 B.n148 163.367
R384 B.n146 B.n107 163.367
R385 B.n142 B.n140 163.367
R386 B.n137 B.n136 163.367
R387 B.n134 B.n113 163.367
R388 B.n130 B.n128 163.367
R389 B.n126 B.n115 163.367
R390 B.n122 B.n120 163.367
R391 B.n118 B.n91 163.367
R392 B.n189 B.n89 163.367
R393 B.n193 B.n89 163.367
R394 B.n193 B.n83 163.367
R395 B.n201 B.n83 163.367
R396 B.n201 B.n81 163.367
R397 B.n205 B.n81 163.367
R398 B.n205 B.n74 163.367
R399 B.n213 B.n74 163.367
R400 B.n213 B.n72 163.367
R401 B.n217 B.n72 163.367
R402 B.n217 B.n67 163.367
R403 B.n226 B.n67 163.367
R404 B.n226 B.n65 163.367
R405 B.n231 B.n65 163.367
R406 B.n231 B.n61 163.367
R407 B.n240 B.n61 163.367
R408 B.n241 B.n240 163.367
R409 B.n241 B.n5 163.367
R410 B.n6 B.n5 163.367
R411 B.n7 B.n6 163.367
R412 B.n246 B.n7 163.367
R413 B.n246 B.n12 163.367
R414 B.n13 B.n12 163.367
R415 B.n14 B.n13 163.367
R416 B.n251 B.n14 163.367
R417 B.n251 B.n19 163.367
R418 B.n20 B.n19 163.367
R419 B.n21 B.n20 163.367
R420 B.n256 B.n21 163.367
R421 B.n256 B.n26 163.367
R422 B.n27 B.n26 163.367
R423 B.n28 B.n27 163.367
R424 B.n261 B.n28 163.367
R425 B.n261 B.n33 163.367
R426 B.n34 B.n33 163.367
R427 B.n35 B.n34 163.367
R428 B.n336 B.n334 163.367
R429 B.n332 B.n39 163.367
R430 B.n328 B.n326 163.367
R431 B.n324 B.n41 163.367
R432 B.n320 B.n318 163.367
R433 B.n316 B.n43 163.367
R434 B.n311 B.n309 163.367
R435 B.n307 B.n47 163.367
R436 B.n303 B.n301 163.367
R437 B.n299 B.n49 163.367
R438 B.n295 B.n293 163.367
R439 B.n291 B.n51 163.367
R440 B.n287 B.n285 163.367
R441 B.n283 B.n56 163.367
R442 B.n279 B.n277 163.367
R443 B.n275 B.n58 163.367
R444 B.n271 B.n269 163.367
R445 B.n108 B.t15 101.547
R446 B.n52 B.t10 101.547
R447 B.n100 B.t21 101.546
R448 B.n44 B.t17 101.546
R449 B.n188 B.n88 97.8422
R450 B.n194 B.n88 97.8422
R451 B.n194 B.n84 97.8422
R452 B.n200 B.n84 97.8422
R453 B.n206 B.n80 97.8422
R454 B.n206 B.n75 97.8422
R455 B.n212 B.n75 97.8422
R456 B.n212 B.n76 97.8422
R457 B.n219 B.n218 97.8422
R458 B.n225 B.n68 97.8422
R459 B.n233 B.n232 97.8422
R460 B.n239 B.n4 97.8422
R461 B.n375 B.n4 97.8422
R462 B.n375 B.n374 97.8422
R463 B.n374 B.n373 97.8422
R464 B.n367 B.n11 97.8422
R465 B.n366 B.n365 97.8422
R466 B.n359 B.n18 97.8422
R467 B.n358 B.n357 97.8422
R468 B.n357 B.n22 97.8422
R469 B.n351 B.n22 97.8422
R470 B.n351 B.n350 97.8422
R471 B.n349 B.n29 97.8422
R472 B.n343 B.n29 97.8422
R473 B.n343 B.n342 97.8422
R474 B.n342 B.n341 97.8422
R475 B.n109 B.t14 88.3592
R476 B.n53 B.t11 88.3592
R477 B.n101 B.t20 88.3589
R478 B.n45 B.t18 88.3589
R479 B.t13 B.n80 79.1372
R480 B.n350 B.t9 79.1372
R481 B.n182 B.n93 71.676
R482 B.n180 B.n95 71.676
R483 B.n176 B.n175 71.676
R484 B.n169 B.n97 71.676
R485 B.n168 B.n167 71.676
R486 B.n161 B.n99 71.676
R487 B.n160 B.n103 71.676
R488 B.n156 B.n155 71.676
R489 B.n149 B.n105 71.676
R490 B.n148 B.n147 71.676
R491 B.n141 B.n107 71.676
R492 B.n140 B.n111 71.676
R493 B.n136 B.n135 71.676
R494 B.n129 B.n113 71.676
R495 B.n128 B.n127 71.676
R496 B.n121 B.n115 71.676
R497 B.n120 B.n119 71.676
R498 B.n335 B.n37 71.676
R499 B.n334 B.n333 71.676
R500 B.n327 B.n39 71.676
R501 B.n326 B.n325 71.676
R502 B.n319 B.n41 71.676
R503 B.n318 B.n317 71.676
R504 B.n310 B.n43 71.676
R505 B.n309 B.n308 71.676
R506 B.n302 B.n47 71.676
R507 B.n301 B.n300 71.676
R508 B.n294 B.n49 71.676
R509 B.n293 B.n292 71.676
R510 B.n286 B.n51 71.676
R511 B.n285 B.n284 71.676
R512 B.n278 B.n56 71.676
R513 B.n277 B.n276 71.676
R514 B.n270 B.n58 71.676
R515 B.n269 B.n268 71.676
R516 B.n268 B.n267 71.676
R517 B.n271 B.n270 71.676
R518 B.n276 B.n275 71.676
R519 B.n279 B.n278 71.676
R520 B.n284 B.n283 71.676
R521 B.n287 B.n286 71.676
R522 B.n292 B.n291 71.676
R523 B.n295 B.n294 71.676
R524 B.n300 B.n299 71.676
R525 B.n303 B.n302 71.676
R526 B.n308 B.n307 71.676
R527 B.n311 B.n310 71.676
R528 B.n317 B.n316 71.676
R529 B.n320 B.n319 71.676
R530 B.n325 B.n324 71.676
R531 B.n328 B.n327 71.676
R532 B.n333 B.n332 71.676
R533 B.n336 B.n335 71.676
R534 B.n183 B.n182 71.676
R535 B.n177 B.n95 71.676
R536 B.n175 B.n174 71.676
R537 B.n170 B.n169 71.676
R538 B.n167 B.n166 71.676
R539 B.n162 B.n161 71.676
R540 B.n157 B.n103 71.676
R541 B.n155 B.n154 71.676
R542 B.n150 B.n149 71.676
R543 B.n147 B.n146 71.676
R544 B.n142 B.n141 71.676
R545 B.n137 B.n111 71.676
R546 B.n135 B.n134 71.676
R547 B.n130 B.n129 71.676
R548 B.n127 B.n126 71.676
R549 B.n122 B.n121 71.676
R550 B.n119 B.n118 71.676
R551 B.n110 B.n109 59.5399
R552 B.n102 B.n101 59.5399
R553 B.n313 B.n45 59.5399
R554 B.n54 B.n53 59.5399
R555 B.n219 B.t4 58.9933
R556 B.n225 B.t2 58.9933
R557 B.n233 B.t7 58.9933
R558 B.n239 B.t0 58.9933
R559 B.n373 B.t5 58.9933
R560 B.n367 B.t3 58.9933
R561 B.n365 B.t6 58.9933
R562 B.n359 B.t1 58.9933
R563 B.n76 B.t4 38.8494
R564 B.n218 B.t2 38.8494
R565 B.n68 B.t7 38.8494
R566 B.n232 B.t0 38.8494
R567 B.n11 B.t5 38.8494
R568 B.t3 B.n366 38.8494
R569 B.n18 B.t6 38.8494
R570 B.t1 B.n358 38.8494
R571 B.n339 B.n338 34.4981
R572 B.n266 B.n265 34.4981
R573 B.n190 B.n90 34.4981
R574 B.n186 B.n185 34.4981
R575 B.n200 B.t13 18.7055
R576 B.t9 B.n349 18.7055
R577 B B.n377 18.0485
R578 B.n109 B.n108 13.1884
R579 B.n101 B.n100 13.1884
R580 B.n45 B.n44 13.1884
R581 B.n53 B.n52 13.1884
R582 B.n338 B.n337 10.6151
R583 B.n337 B.n38 10.6151
R584 B.n331 B.n38 10.6151
R585 B.n331 B.n330 10.6151
R586 B.n330 B.n329 10.6151
R587 B.n329 B.n40 10.6151
R588 B.n323 B.n40 10.6151
R589 B.n323 B.n322 10.6151
R590 B.n322 B.n321 10.6151
R591 B.n321 B.n42 10.6151
R592 B.n315 B.n42 10.6151
R593 B.n315 B.n314 10.6151
R594 B.n312 B.n46 10.6151
R595 B.n306 B.n46 10.6151
R596 B.n306 B.n305 10.6151
R597 B.n305 B.n304 10.6151
R598 B.n304 B.n48 10.6151
R599 B.n298 B.n48 10.6151
R600 B.n298 B.n297 10.6151
R601 B.n297 B.n296 10.6151
R602 B.n296 B.n50 10.6151
R603 B.n290 B.n289 10.6151
R604 B.n289 B.n288 10.6151
R605 B.n288 B.n55 10.6151
R606 B.n282 B.n55 10.6151
R607 B.n282 B.n281 10.6151
R608 B.n281 B.n280 10.6151
R609 B.n280 B.n57 10.6151
R610 B.n274 B.n57 10.6151
R611 B.n274 B.n273 10.6151
R612 B.n273 B.n272 10.6151
R613 B.n272 B.n59 10.6151
R614 B.n266 B.n59 10.6151
R615 B.n191 B.n190 10.6151
R616 B.n192 B.n191 10.6151
R617 B.n192 B.n82 10.6151
R618 B.n202 B.n82 10.6151
R619 B.n203 B.n202 10.6151
R620 B.n204 B.n203 10.6151
R621 B.n204 B.n73 10.6151
R622 B.n214 B.n73 10.6151
R623 B.n215 B.n214 10.6151
R624 B.n216 B.n215 10.6151
R625 B.n216 B.n66 10.6151
R626 B.n227 B.n66 10.6151
R627 B.n228 B.n227 10.6151
R628 B.n230 B.n228 10.6151
R629 B.n230 B.n229 10.6151
R630 B.n229 B.n60 10.6151
R631 B.n242 B.n60 10.6151
R632 B.n243 B.n242 10.6151
R633 B.n244 B.n243 10.6151
R634 B.n245 B.n244 10.6151
R635 B.n247 B.n245 10.6151
R636 B.n248 B.n247 10.6151
R637 B.n249 B.n248 10.6151
R638 B.n250 B.n249 10.6151
R639 B.n252 B.n250 10.6151
R640 B.n253 B.n252 10.6151
R641 B.n254 B.n253 10.6151
R642 B.n255 B.n254 10.6151
R643 B.n257 B.n255 10.6151
R644 B.n258 B.n257 10.6151
R645 B.n259 B.n258 10.6151
R646 B.n260 B.n259 10.6151
R647 B.n262 B.n260 10.6151
R648 B.n263 B.n262 10.6151
R649 B.n264 B.n263 10.6151
R650 B.n265 B.n264 10.6151
R651 B.n185 B.n184 10.6151
R652 B.n184 B.n94 10.6151
R653 B.n179 B.n94 10.6151
R654 B.n179 B.n178 10.6151
R655 B.n178 B.n96 10.6151
R656 B.n173 B.n96 10.6151
R657 B.n173 B.n172 10.6151
R658 B.n172 B.n171 10.6151
R659 B.n171 B.n98 10.6151
R660 B.n165 B.n98 10.6151
R661 B.n165 B.n164 10.6151
R662 B.n164 B.n163 10.6151
R663 B.n159 B.n158 10.6151
R664 B.n158 B.n104 10.6151
R665 B.n153 B.n104 10.6151
R666 B.n153 B.n152 10.6151
R667 B.n152 B.n151 10.6151
R668 B.n151 B.n106 10.6151
R669 B.n145 B.n106 10.6151
R670 B.n145 B.n144 10.6151
R671 B.n144 B.n143 10.6151
R672 B.n139 B.n138 10.6151
R673 B.n138 B.n112 10.6151
R674 B.n133 B.n112 10.6151
R675 B.n133 B.n132 10.6151
R676 B.n132 B.n131 10.6151
R677 B.n131 B.n114 10.6151
R678 B.n125 B.n114 10.6151
R679 B.n125 B.n124 10.6151
R680 B.n124 B.n123 10.6151
R681 B.n123 B.n116 10.6151
R682 B.n117 B.n116 10.6151
R683 B.n117 B.n90 10.6151
R684 B.n186 B.n86 10.6151
R685 B.n196 B.n86 10.6151
R686 B.n197 B.n196 10.6151
R687 B.n198 B.n197 10.6151
R688 B.n198 B.n78 10.6151
R689 B.n208 B.n78 10.6151
R690 B.n209 B.n208 10.6151
R691 B.n210 B.n209 10.6151
R692 B.n210 B.n70 10.6151
R693 B.n221 B.n70 10.6151
R694 B.n222 B.n221 10.6151
R695 B.n223 B.n222 10.6151
R696 B.n223 B.n63 10.6151
R697 B.n235 B.n63 10.6151
R698 B.n236 B.n235 10.6151
R699 B.n237 B.n236 10.6151
R700 B.n237 B.n0 10.6151
R701 B.n371 B.n1 10.6151
R702 B.n371 B.n370 10.6151
R703 B.n370 B.n369 10.6151
R704 B.n369 B.n9 10.6151
R705 B.n363 B.n9 10.6151
R706 B.n363 B.n362 10.6151
R707 B.n362 B.n361 10.6151
R708 B.n361 B.n16 10.6151
R709 B.n355 B.n16 10.6151
R710 B.n355 B.n354 10.6151
R711 B.n354 B.n353 10.6151
R712 B.n353 B.n24 10.6151
R713 B.n347 B.n24 10.6151
R714 B.n347 B.n346 10.6151
R715 B.n346 B.n345 10.6151
R716 B.n345 B.n31 10.6151
R717 B.n339 B.n31 10.6151
R718 B.n314 B.n313 9.36635
R719 B.n290 B.n54 9.36635
R720 B.n163 B.n102 9.36635
R721 B.n139 B.n110 9.36635
R722 B.n377 B.n0 2.81026
R723 B.n377 B.n1 2.81026
R724 B.n313 B.n312 1.24928
R725 B.n54 B.n50 1.24928
R726 B.n159 B.n102 1.24928
R727 B.n143 B.n110 1.24928
R728 VP.n3 VP.t7 305.515
R729 VP.n12 VP.t1 289.993
R730 VP.n1 VP.t2 289.993
R731 VP.n6 VP.t0 289.993
R732 VP.n10 VP.t4 276.118
R733 VP.n11 VP.t3 276.118
R734 VP.n5 VP.t5 276.118
R735 VP.n4 VP.t6 276.118
R736 VP.n13 VP.n12 161.3
R737 VP.n5 VP.n2 161.3
R738 VP.n7 VP.n6 161.3
R739 VP.n11 VP.n0 161.3
R740 VP.n10 VP.n9 161.3
R741 VP.n8 VP.n1 161.3
R742 VP.n3 VP.n2 73.1314
R743 VP.n11 VP.n10 48.2005
R744 VP.n5 VP.n4 48.2005
R745 VP.n10 VP.n1 34.3247
R746 VP.n12 VP.n11 34.3247
R747 VP.n6 VP.n5 34.3247
R748 VP.n8 VP.n7 33.1444
R749 VP.n4 VP.n3 15.5045
R750 VP.n7 VP.n2 0.189894
R751 VP.n9 VP.n8 0.189894
R752 VP.n9 VP.n0 0.189894
R753 VP.n13 VP.n0 0.189894
R754 VP VP.n13 0.0516364
R755 VDD1 VDD1.n0 92.2442
R756 VDD1.n3 VDD1.n2 92.1306
R757 VDD1.n3 VDD1.n1 92.1306
R758 VDD1.n5 VDD1.n4 91.8929
R759 VDD1.n5 VDD1.n3 28.9793
R760 VDD1.n4 VDD1.t2 8.35493
R761 VDD1.n4 VDD1.t7 8.35493
R762 VDD1.n0 VDD1.t0 8.35493
R763 VDD1.n0 VDD1.t1 8.35493
R764 VDD1.n2 VDD1.t4 8.35493
R765 VDD1.n2 VDD1.t6 8.35493
R766 VDD1.n1 VDD1.t5 8.35493
R767 VDD1.n1 VDD1.t3 8.35493
R768 VDD1 VDD1.n5 0.235414
C0 VTAIL VDD2 4.51169f
C1 VN VDD1 0.152804f
C2 VDD1 VP 1.14985f
C3 VDD2 VDD1 0.653877f
C4 VN VP 3.13392f
C5 VTAIL VDD1 4.47236f
C6 VDD2 VN 1.01754f
C7 VDD2 VP 0.285974f
C8 VTAIL VN 1.08685f
C9 VTAIL VP 1.10096f
C10 VDD2 B 2.305961f
C11 VDD1 B 2.495898f
C12 VTAIL B 3.110554f
C13 VN B 5.466835f
C14 VP B 4.477253f
C15 VDD1.t0 B 0.043803f
C16 VDD1.t1 B 0.043803f
C17 VDD1.n0 B 0.293773f
C18 VDD1.t5 B 0.043803f
C19 VDD1.t3 B 0.043803f
C20 VDD1.n1 B 0.293432f
C21 VDD1.t4 B 0.043803f
C22 VDD1.t6 B 0.043803f
C23 VDD1.n2 B 0.293432f
C24 VDD1.n3 B 1.34768f
C25 VDD1.t2 B 0.043803f
C26 VDD1.t7 B 0.043803f
C27 VDD1.n4 B 0.292769f
C28 VDD1.n5 B 1.32172f
C29 VP.n0 B 0.032232f
C30 VP.t2 B 0.084118f
C31 VP.n1 B 0.055971f
C32 VP.n2 B 0.104212f
C33 VP.t5 B 0.081672f
C34 VP.t6 B 0.081672f
C35 VP.t7 B 0.086964f
C36 VP.n3 B 0.053359f
C37 VP.n4 B 0.061198f
C38 VP.n5 B 0.061198f
C39 VP.t0 B 0.084118f
C40 VP.n6 B 0.055971f
C41 VP.n7 B 0.862158f
C42 VP.n8 B 0.897115f
C43 VP.n9 B 0.032232f
C44 VP.t4 B 0.081672f
C45 VP.n10 B 0.061198f
C46 VP.t3 B 0.081672f
C47 VP.n11 B 0.061198f
C48 VP.t1 B 0.084118f
C49 VP.n12 B 0.055971f
C50 VP.n13 B 0.024978f
C51 VTAIL.t14 B 0.041271f
C52 VTAIL.t9 B 0.041271f
C53 VTAIL.n0 B 0.238429f
C54 VTAIL.n1 B 0.226145f
C55 VTAIL.t15 B 0.320023f
C56 VTAIL.n2 B 0.286336f
C57 VTAIL.t0 B 0.320023f
C58 VTAIL.n3 B 0.286336f
C59 VTAIL.t2 B 0.041271f
C60 VTAIL.t7 B 0.041271f
C61 VTAIL.n4 B 0.238429f
C62 VTAIL.n5 B 0.263637f
C63 VTAIL.t4 B 0.320023f
C64 VTAIL.n6 B 0.73901f
C65 VTAIL.t11 B 0.320024f
C66 VTAIL.n7 B 0.739009f
C67 VTAIL.t10 B 0.041271f
C68 VTAIL.t12 B 0.041271f
C69 VTAIL.n8 B 0.238431f
C70 VTAIL.n9 B 0.263635f
C71 VTAIL.t13 B 0.320024f
C72 VTAIL.n10 B 0.286335f
C73 VTAIL.t5 B 0.320024f
C74 VTAIL.n11 B 0.286335f
C75 VTAIL.t3 B 0.041271f
C76 VTAIL.t6 B 0.041271f
C77 VTAIL.n12 B 0.238431f
C78 VTAIL.n13 B 0.263635f
C79 VTAIL.t1 B 0.320024f
C80 VTAIL.n14 B 0.739009f
C81 VTAIL.t8 B 0.320023f
C82 VTAIL.n15 B 0.734879f
C83 VDD2.t4 B 0.04466f
C84 VDD2.t2 B 0.04466f
C85 VDD2.n0 B 0.299175f
C86 VDD2.t7 B 0.04466f
C87 VDD2.t5 B 0.04466f
C88 VDD2.n1 B 0.299175f
C89 VDD2.n2 B 1.32268f
C90 VDD2.t6 B 0.04466f
C91 VDD2.t0 B 0.04466f
C92 VDD2.n3 B 0.298499f
C93 VDD2.n4 B 1.31983f
C94 VDD2.t1 B 0.04466f
C95 VDD2.t3 B 0.04466f
C96 VDD2.n5 B 0.299162f
C97 VN.n0 B 0.102711f
C98 VN.t0 B 0.085711f
C99 VN.n1 B 0.05259f
C100 VN.t1 B 0.080496f
C101 VN.n2 B 0.060317f
C102 VN.t6 B 0.080496f
C103 VN.n3 B 0.060317f
C104 VN.t7 B 0.082906f
C105 VN.n4 B 0.055165f
C106 VN.n5 B 0.024619f
C107 VN.n6 B 0.102711f
C108 VN.t4 B 0.082906f
C109 VN.t3 B 0.080496f
C110 VN.t2 B 0.085711f
C111 VN.n7 B 0.05259f
C112 VN.n8 B 0.060317f
C113 VN.t5 B 0.080496f
C114 VN.n9 B 0.060317f
C115 VN.n10 B 0.055165f
C116 VN.n11 B 0.870943f
.ends

