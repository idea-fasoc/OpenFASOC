* NGSPICE file created from diff_pair_sample_0211.ext - technology: sky130A

.subckt diff_pair_sample_0211 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0 ps=0 w=2.43 l=1.59
X2 VDD2.t7 VN.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.9477 ps=5.64 w=2.43 l=1.59
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0 ps=0 w=2.43 l=1.59
X4 VTAIL.t1 VN.t1 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X5 VTAIL.t15 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X6 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0 ps=0 w=2.43 l=1.59
X7 VTAIL.t3 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0.40095 ps=2.76 w=2.43 l=1.59
X8 VDD2.t4 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X9 VDD1.t5 VP.t2 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.9477 ps=5.64 w=2.43 l=1.59
X10 VDD2.t3 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.9477 ps=5.64 w=2.43 l=1.59
X11 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X12 VTAIL.t5 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0.40095 ps=2.76 w=2.43 l=1.59
X13 VTAIL.t6 VN.t7 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X14 VDD1.t4 VP.t3 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.9477 ps=5.64 w=2.43 l=1.59
X15 VTAIL.t12 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X16 VDD1.t2 VP.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.40095 pd=2.76 as=0.40095 ps=2.76 w=2.43 l=1.59
X17 VTAIL.t9 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0.40095 ps=2.76 w=2.43 l=1.59
X18 VTAIL.t8 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0.40095 ps=2.76 w=2.43 l=1.59
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9477 pd=5.64 as=0 ps=0 w=2.43 l=1.59
R0 VP.n28 VP.n27 179.406
R1 VP.n50 VP.n49 179.406
R2 VP.n26 VP.n25 179.406
R3 VP.n13 VP.n12 161.3
R4 VP.n14 VP.n9 161.3
R5 VP.n16 VP.n15 161.3
R6 VP.n17 VP.n8 161.3
R7 VP.n20 VP.n19 161.3
R8 VP.n21 VP.n7 161.3
R9 VP.n23 VP.n22 161.3
R10 VP.n24 VP.n6 161.3
R11 VP.n48 VP.n0 161.3
R12 VP.n47 VP.n46 161.3
R13 VP.n45 VP.n1 161.3
R14 VP.n44 VP.n43 161.3
R15 VP.n41 VP.n2 161.3
R16 VP.n40 VP.n39 161.3
R17 VP.n38 VP.n3 161.3
R18 VP.n37 VP.n36 161.3
R19 VP.n34 VP.n4 161.3
R20 VP.n33 VP.n32 161.3
R21 VP.n31 VP.n5 161.3
R22 VP.n30 VP.n29 161.3
R23 VP.n10 VP.t6 68.617
R24 VP.n33 VP.n5 56.5193
R25 VP.n47 VP.n1 56.5193
R26 VP.n23 VP.n7 56.5193
R27 VP.n40 VP.n3 56.5193
R28 VP.n16 VP.n9 56.5193
R29 VP.n11 VP.n10 55.7366
R30 VP.n27 VP.n26 38.8111
R31 VP.n28 VP.t7 36.8326
R32 VP.n35 VP.t0 36.8326
R33 VP.n42 VP.t1 36.8326
R34 VP.n49 VP.t2 36.8326
R35 VP.n25 VP.t3 36.8326
R36 VP.n18 VP.t4 36.8326
R37 VP.n11 VP.t5 36.8326
R38 VP.n29 VP.n5 24.4675
R39 VP.n34 VP.n33 24.4675
R40 VP.n36 VP.n3 24.4675
R41 VP.n41 VP.n40 24.4675
R42 VP.n43 VP.n1 24.4675
R43 VP.n48 VP.n47 24.4675
R44 VP.n24 VP.n23 24.4675
R45 VP.n17 VP.n16 24.4675
R46 VP.n19 VP.n7 24.4675
R47 VP.n12 VP.n9 24.4675
R48 VP.n13 VP.n10 18.144
R49 VP.n35 VP.n34 14.1914
R50 VP.n43 VP.n42 14.1914
R51 VP.n19 VP.n18 14.1914
R52 VP.n36 VP.n35 10.2766
R53 VP.n42 VP.n41 10.2766
R54 VP.n18 VP.n17 10.2766
R55 VP.n12 VP.n11 10.2766
R56 VP.n29 VP.n28 6.36192
R57 VP.n49 VP.n48 6.36192
R58 VP.n25 VP.n24 6.36192
R59 VP.n14 VP.n13 0.189894
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n8 0.189894
R62 VP.n20 VP.n8 0.189894
R63 VP.n21 VP.n20 0.189894
R64 VP.n22 VP.n21 0.189894
R65 VP.n22 VP.n6 0.189894
R66 VP.n26 VP.n6 0.189894
R67 VP.n30 VP.n27 0.189894
R68 VP.n31 VP.n30 0.189894
R69 VP.n32 VP.n31 0.189894
R70 VP.n32 VP.n4 0.189894
R71 VP.n37 VP.n4 0.189894
R72 VP.n38 VP.n37 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP.n50 VP.n0 0.189894
R80 VP VP.n50 0.0516364
R81 VTAIL.n98 VTAIL.n92 289.615
R82 VTAIL.n8 VTAIL.n2 289.615
R83 VTAIL.n20 VTAIL.n14 289.615
R84 VTAIL.n34 VTAIL.n28 289.615
R85 VTAIL.n86 VTAIL.n80 289.615
R86 VTAIL.n72 VTAIL.n66 289.615
R87 VTAIL.n60 VTAIL.n54 289.615
R88 VTAIL.n46 VTAIL.n40 289.615
R89 VTAIL.n97 VTAIL.n96 185
R90 VTAIL.n99 VTAIL.n98 185
R91 VTAIL.n7 VTAIL.n6 185
R92 VTAIL.n9 VTAIL.n8 185
R93 VTAIL.n19 VTAIL.n18 185
R94 VTAIL.n21 VTAIL.n20 185
R95 VTAIL.n33 VTAIL.n32 185
R96 VTAIL.n35 VTAIL.n34 185
R97 VTAIL.n87 VTAIL.n86 185
R98 VTAIL.n85 VTAIL.n84 185
R99 VTAIL.n73 VTAIL.n72 185
R100 VTAIL.n71 VTAIL.n70 185
R101 VTAIL.n61 VTAIL.n60 185
R102 VTAIL.n59 VTAIL.n58 185
R103 VTAIL.n47 VTAIL.n46 185
R104 VTAIL.n45 VTAIL.n44 185
R105 VTAIL.n95 VTAIL.t7 151.613
R106 VTAIL.n5 VTAIL.t5 151.613
R107 VTAIL.n17 VTAIL.t11 151.613
R108 VTAIL.n31 VTAIL.t8 151.613
R109 VTAIL.n83 VTAIL.t13 151.613
R110 VTAIL.n69 VTAIL.t9 151.613
R111 VTAIL.n57 VTAIL.t2 151.613
R112 VTAIL.n43 VTAIL.t3 151.613
R113 VTAIL.n98 VTAIL.n97 104.615
R114 VTAIL.n8 VTAIL.n7 104.615
R115 VTAIL.n20 VTAIL.n19 104.615
R116 VTAIL.n34 VTAIL.n33 104.615
R117 VTAIL.n86 VTAIL.n85 104.615
R118 VTAIL.n72 VTAIL.n71 104.615
R119 VTAIL.n60 VTAIL.n59 104.615
R120 VTAIL.n46 VTAIL.n45 104.615
R121 VTAIL.n79 VTAIL.n78 68.8623
R122 VTAIL.n53 VTAIL.n52 68.8623
R123 VTAIL.n1 VTAIL.n0 68.8622
R124 VTAIL.n27 VTAIL.n26 68.8622
R125 VTAIL.n97 VTAIL.t7 52.3082
R126 VTAIL.n7 VTAIL.t5 52.3082
R127 VTAIL.n19 VTAIL.t11 52.3082
R128 VTAIL.n33 VTAIL.t8 52.3082
R129 VTAIL.n85 VTAIL.t13 52.3082
R130 VTAIL.n71 VTAIL.t9 52.3082
R131 VTAIL.n59 VTAIL.t2 52.3082
R132 VTAIL.n45 VTAIL.t3 52.3082
R133 VTAIL.n103 VTAIL.n102 32.7672
R134 VTAIL.n13 VTAIL.n12 32.7672
R135 VTAIL.n25 VTAIL.n24 32.7672
R136 VTAIL.n39 VTAIL.n38 32.7672
R137 VTAIL.n91 VTAIL.n90 32.7672
R138 VTAIL.n77 VTAIL.n76 32.7672
R139 VTAIL.n65 VTAIL.n64 32.7672
R140 VTAIL.n51 VTAIL.n50 32.7672
R141 VTAIL.n103 VTAIL.n91 16.1169
R142 VTAIL.n51 VTAIL.n39 16.1169
R143 VTAIL.n96 VTAIL.n95 15.3979
R144 VTAIL.n6 VTAIL.n5 15.3979
R145 VTAIL.n18 VTAIL.n17 15.3979
R146 VTAIL.n32 VTAIL.n31 15.3979
R147 VTAIL.n84 VTAIL.n83 15.3979
R148 VTAIL.n70 VTAIL.n69 15.3979
R149 VTAIL.n58 VTAIL.n57 15.3979
R150 VTAIL.n44 VTAIL.n43 15.3979
R151 VTAIL.n99 VTAIL.n94 12.8005
R152 VTAIL.n9 VTAIL.n4 12.8005
R153 VTAIL.n21 VTAIL.n16 12.8005
R154 VTAIL.n35 VTAIL.n30 12.8005
R155 VTAIL.n87 VTAIL.n82 12.8005
R156 VTAIL.n73 VTAIL.n68 12.8005
R157 VTAIL.n61 VTAIL.n56 12.8005
R158 VTAIL.n47 VTAIL.n42 12.8005
R159 VTAIL.n100 VTAIL.n92 12.0247
R160 VTAIL.n10 VTAIL.n2 12.0247
R161 VTAIL.n22 VTAIL.n14 12.0247
R162 VTAIL.n36 VTAIL.n28 12.0247
R163 VTAIL.n88 VTAIL.n80 12.0247
R164 VTAIL.n74 VTAIL.n66 12.0247
R165 VTAIL.n62 VTAIL.n54 12.0247
R166 VTAIL.n48 VTAIL.n40 12.0247
R167 VTAIL.n102 VTAIL.n101 9.45567
R168 VTAIL.n12 VTAIL.n11 9.45567
R169 VTAIL.n24 VTAIL.n23 9.45567
R170 VTAIL.n38 VTAIL.n37 9.45567
R171 VTAIL.n90 VTAIL.n89 9.45567
R172 VTAIL.n76 VTAIL.n75 9.45567
R173 VTAIL.n64 VTAIL.n63 9.45567
R174 VTAIL.n50 VTAIL.n49 9.45567
R175 VTAIL.n101 VTAIL.n100 9.3005
R176 VTAIL.n94 VTAIL.n93 9.3005
R177 VTAIL.n11 VTAIL.n10 9.3005
R178 VTAIL.n4 VTAIL.n3 9.3005
R179 VTAIL.n23 VTAIL.n22 9.3005
R180 VTAIL.n16 VTAIL.n15 9.3005
R181 VTAIL.n37 VTAIL.n36 9.3005
R182 VTAIL.n30 VTAIL.n29 9.3005
R183 VTAIL.n89 VTAIL.n88 9.3005
R184 VTAIL.n82 VTAIL.n81 9.3005
R185 VTAIL.n75 VTAIL.n74 9.3005
R186 VTAIL.n68 VTAIL.n67 9.3005
R187 VTAIL.n63 VTAIL.n62 9.3005
R188 VTAIL.n56 VTAIL.n55 9.3005
R189 VTAIL.n49 VTAIL.n48 9.3005
R190 VTAIL.n42 VTAIL.n41 9.3005
R191 VTAIL.n0 VTAIL.t0 8.14865
R192 VTAIL.n0 VTAIL.t1 8.14865
R193 VTAIL.n26 VTAIL.t14 8.14865
R194 VTAIL.n26 VTAIL.t15 8.14865
R195 VTAIL.n78 VTAIL.t10 8.14865
R196 VTAIL.n78 VTAIL.t12 8.14865
R197 VTAIL.n52 VTAIL.t4 8.14865
R198 VTAIL.n52 VTAIL.t6 8.14865
R199 VTAIL.n95 VTAIL.n93 4.69785
R200 VTAIL.n5 VTAIL.n3 4.69785
R201 VTAIL.n17 VTAIL.n15 4.69785
R202 VTAIL.n31 VTAIL.n29 4.69785
R203 VTAIL.n83 VTAIL.n81 4.69785
R204 VTAIL.n69 VTAIL.n67 4.69785
R205 VTAIL.n57 VTAIL.n55 4.69785
R206 VTAIL.n43 VTAIL.n41 4.69785
R207 VTAIL.n102 VTAIL.n92 1.93989
R208 VTAIL.n12 VTAIL.n2 1.93989
R209 VTAIL.n24 VTAIL.n14 1.93989
R210 VTAIL.n38 VTAIL.n28 1.93989
R211 VTAIL.n90 VTAIL.n80 1.93989
R212 VTAIL.n76 VTAIL.n66 1.93989
R213 VTAIL.n64 VTAIL.n54 1.93989
R214 VTAIL.n50 VTAIL.n40 1.93989
R215 VTAIL.n53 VTAIL.n51 1.65567
R216 VTAIL.n65 VTAIL.n53 1.65567
R217 VTAIL.n79 VTAIL.n77 1.65567
R218 VTAIL.n91 VTAIL.n79 1.65567
R219 VTAIL.n39 VTAIL.n27 1.65567
R220 VTAIL.n27 VTAIL.n25 1.65567
R221 VTAIL.n13 VTAIL.n1 1.65567
R222 VTAIL VTAIL.n103 1.59748
R223 VTAIL.n100 VTAIL.n99 1.16414
R224 VTAIL.n10 VTAIL.n9 1.16414
R225 VTAIL.n22 VTAIL.n21 1.16414
R226 VTAIL.n36 VTAIL.n35 1.16414
R227 VTAIL.n88 VTAIL.n87 1.16414
R228 VTAIL.n74 VTAIL.n73 1.16414
R229 VTAIL.n62 VTAIL.n61 1.16414
R230 VTAIL.n48 VTAIL.n47 1.16414
R231 VTAIL.n77 VTAIL.n65 0.470328
R232 VTAIL.n25 VTAIL.n13 0.470328
R233 VTAIL.n96 VTAIL.n94 0.388379
R234 VTAIL.n6 VTAIL.n4 0.388379
R235 VTAIL.n18 VTAIL.n16 0.388379
R236 VTAIL.n32 VTAIL.n30 0.388379
R237 VTAIL.n84 VTAIL.n82 0.388379
R238 VTAIL.n70 VTAIL.n68 0.388379
R239 VTAIL.n58 VTAIL.n56 0.388379
R240 VTAIL.n44 VTAIL.n42 0.388379
R241 VTAIL.n101 VTAIL.n93 0.155672
R242 VTAIL.n11 VTAIL.n3 0.155672
R243 VTAIL.n23 VTAIL.n15 0.155672
R244 VTAIL.n37 VTAIL.n29 0.155672
R245 VTAIL.n89 VTAIL.n81 0.155672
R246 VTAIL.n75 VTAIL.n67 0.155672
R247 VTAIL.n63 VTAIL.n55 0.155672
R248 VTAIL.n49 VTAIL.n41 0.155672
R249 VTAIL VTAIL.n1 0.0586897
R250 VDD1 VDD1.n0 86.4269
R251 VDD1.n3 VDD1.n2 86.3132
R252 VDD1.n3 VDD1.n1 86.3132
R253 VDD1.n5 VDD1.n4 85.541
R254 VDD1.n5 VDD1.n3 33.8414
R255 VDD1.n4 VDD1.t3 8.14865
R256 VDD1.n4 VDD1.t4 8.14865
R257 VDD1.n0 VDD1.t1 8.14865
R258 VDD1.n0 VDD1.t2 8.14865
R259 VDD1.n2 VDD1.t6 8.14865
R260 VDD1.n2 VDD1.t5 8.14865
R261 VDD1.n1 VDD1.t0 8.14865
R262 VDD1.n1 VDD1.t7 8.14865
R263 VDD1 VDD1.n5 0.769897
R264 B.n489 B.n488 585
R265 B.n490 B.n489 585
R266 B.n162 B.n87 585
R267 B.n161 B.n160 585
R268 B.n159 B.n158 585
R269 B.n157 B.n156 585
R270 B.n155 B.n154 585
R271 B.n153 B.n152 585
R272 B.n151 B.n150 585
R273 B.n149 B.n148 585
R274 B.n147 B.n146 585
R275 B.n145 B.n144 585
R276 B.n143 B.n142 585
R277 B.n141 B.n140 585
R278 B.n139 B.n138 585
R279 B.n136 B.n135 585
R280 B.n134 B.n133 585
R281 B.n132 B.n131 585
R282 B.n130 B.n129 585
R283 B.n128 B.n127 585
R284 B.n126 B.n125 585
R285 B.n124 B.n123 585
R286 B.n122 B.n121 585
R287 B.n120 B.n119 585
R288 B.n118 B.n117 585
R289 B.n116 B.n115 585
R290 B.n114 B.n113 585
R291 B.n112 B.n111 585
R292 B.n110 B.n109 585
R293 B.n108 B.n107 585
R294 B.n106 B.n105 585
R295 B.n104 B.n103 585
R296 B.n102 B.n101 585
R297 B.n100 B.n99 585
R298 B.n98 B.n97 585
R299 B.n96 B.n95 585
R300 B.n94 B.n93 585
R301 B.n67 B.n66 585
R302 B.n487 B.n68 585
R303 B.n491 B.n68 585
R304 B.n486 B.n485 585
R305 B.n485 B.n64 585
R306 B.n484 B.n63 585
R307 B.n497 B.n63 585
R308 B.n483 B.n62 585
R309 B.n498 B.n62 585
R310 B.n482 B.n61 585
R311 B.n499 B.n61 585
R312 B.n481 B.n480 585
R313 B.n480 B.n57 585
R314 B.n479 B.n56 585
R315 B.n505 B.n56 585
R316 B.n478 B.n55 585
R317 B.n506 B.n55 585
R318 B.n477 B.n54 585
R319 B.n507 B.n54 585
R320 B.n476 B.n475 585
R321 B.n475 B.n50 585
R322 B.n474 B.n49 585
R323 B.n513 B.n49 585
R324 B.n473 B.n48 585
R325 B.n514 B.n48 585
R326 B.n472 B.n47 585
R327 B.n515 B.n47 585
R328 B.n471 B.n470 585
R329 B.n470 B.n43 585
R330 B.n469 B.n42 585
R331 B.n521 B.n42 585
R332 B.n468 B.n41 585
R333 B.n522 B.n41 585
R334 B.n467 B.n40 585
R335 B.n523 B.n40 585
R336 B.n466 B.n465 585
R337 B.n465 B.n36 585
R338 B.n464 B.n35 585
R339 B.n529 B.n35 585
R340 B.n463 B.n34 585
R341 B.n530 B.n34 585
R342 B.n462 B.n33 585
R343 B.n531 B.n33 585
R344 B.n461 B.n460 585
R345 B.n460 B.n29 585
R346 B.n459 B.n28 585
R347 B.n537 B.n28 585
R348 B.n458 B.n27 585
R349 B.n538 B.n27 585
R350 B.n457 B.n26 585
R351 B.n539 B.n26 585
R352 B.n456 B.n455 585
R353 B.n455 B.n22 585
R354 B.n454 B.n21 585
R355 B.n545 B.n21 585
R356 B.n453 B.n20 585
R357 B.n546 B.n20 585
R358 B.n452 B.n19 585
R359 B.n547 B.n19 585
R360 B.n451 B.n450 585
R361 B.n450 B.n15 585
R362 B.n449 B.n14 585
R363 B.n553 B.n14 585
R364 B.n448 B.n13 585
R365 B.n554 B.n13 585
R366 B.n447 B.n12 585
R367 B.n555 B.n12 585
R368 B.n446 B.n445 585
R369 B.n445 B.n444 585
R370 B.n443 B.n442 585
R371 B.n443 B.n8 585
R372 B.n441 B.n7 585
R373 B.n562 B.n7 585
R374 B.n440 B.n6 585
R375 B.n563 B.n6 585
R376 B.n439 B.n5 585
R377 B.n564 B.n5 585
R378 B.n438 B.n437 585
R379 B.n437 B.n4 585
R380 B.n436 B.n163 585
R381 B.n436 B.n435 585
R382 B.n426 B.n164 585
R383 B.n165 B.n164 585
R384 B.n428 B.n427 585
R385 B.n429 B.n428 585
R386 B.n425 B.n170 585
R387 B.n170 B.n169 585
R388 B.n424 B.n423 585
R389 B.n423 B.n422 585
R390 B.n172 B.n171 585
R391 B.n173 B.n172 585
R392 B.n415 B.n414 585
R393 B.n416 B.n415 585
R394 B.n413 B.n178 585
R395 B.n178 B.n177 585
R396 B.n412 B.n411 585
R397 B.n411 B.n410 585
R398 B.n180 B.n179 585
R399 B.n181 B.n180 585
R400 B.n403 B.n402 585
R401 B.n404 B.n403 585
R402 B.n401 B.n186 585
R403 B.n186 B.n185 585
R404 B.n400 B.n399 585
R405 B.n399 B.n398 585
R406 B.n188 B.n187 585
R407 B.n189 B.n188 585
R408 B.n391 B.n390 585
R409 B.n392 B.n391 585
R410 B.n389 B.n194 585
R411 B.n194 B.n193 585
R412 B.n388 B.n387 585
R413 B.n387 B.n386 585
R414 B.n196 B.n195 585
R415 B.n197 B.n196 585
R416 B.n379 B.n378 585
R417 B.n380 B.n379 585
R418 B.n377 B.n201 585
R419 B.n205 B.n201 585
R420 B.n376 B.n375 585
R421 B.n375 B.n374 585
R422 B.n203 B.n202 585
R423 B.n204 B.n203 585
R424 B.n367 B.n366 585
R425 B.n368 B.n367 585
R426 B.n365 B.n210 585
R427 B.n210 B.n209 585
R428 B.n364 B.n363 585
R429 B.n363 B.n362 585
R430 B.n212 B.n211 585
R431 B.n213 B.n212 585
R432 B.n355 B.n354 585
R433 B.n356 B.n355 585
R434 B.n353 B.n218 585
R435 B.n218 B.n217 585
R436 B.n352 B.n351 585
R437 B.n351 B.n350 585
R438 B.n220 B.n219 585
R439 B.n221 B.n220 585
R440 B.n343 B.n342 585
R441 B.n344 B.n343 585
R442 B.n341 B.n226 585
R443 B.n226 B.n225 585
R444 B.n340 B.n339 585
R445 B.n339 B.n338 585
R446 B.n228 B.n227 585
R447 B.n229 B.n228 585
R448 B.n331 B.n330 585
R449 B.n332 B.n331 585
R450 B.n232 B.n231 585
R451 B.n257 B.n255 585
R452 B.n258 B.n254 585
R453 B.n258 B.n233 585
R454 B.n261 B.n260 585
R455 B.n262 B.n253 585
R456 B.n264 B.n263 585
R457 B.n266 B.n252 585
R458 B.n269 B.n268 585
R459 B.n270 B.n251 585
R460 B.n272 B.n271 585
R461 B.n274 B.n250 585
R462 B.n277 B.n276 585
R463 B.n278 B.n249 585
R464 B.n283 B.n282 585
R465 B.n285 B.n248 585
R466 B.n288 B.n287 585
R467 B.n289 B.n247 585
R468 B.n291 B.n290 585
R469 B.n293 B.n246 585
R470 B.n296 B.n295 585
R471 B.n297 B.n245 585
R472 B.n299 B.n298 585
R473 B.n301 B.n244 585
R474 B.n304 B.n303 585
R475 B.n305 B.n240 585
R476 B.n307 B.n306 585
R477 B.n309 B.n239 585
R478 B.n312 B.n311 585
R479 B.n313 B.n238 585
R480 B.n315 B.n314 585
R481 B.n317 B.n237 585
R482 B.n320 B.n319 585
R483 B.n321 B.n236 585
R484 B.n323 B.n322 585
R485 B.n325 B.n235 585
R486 B.n328 B.n327 585
R487 B.n329 B.n234 585
R488 B.n334 B.n333 585
R489 B.n333 B.n332 585
R490 B.n335 B.n230 585
R491 B.n230 B.n229 585
R492 B.n337 B.n336 585
R493 B.n338 B.n337 585
R494 B.n224 B.n223 585
R495 B.n225 B.n224 585
R496 B.n346 B.n345 585
R497 B.n345 B.n344 585
R498 B.n347 B.n222 585
R499 B.n222 B.n221 585
R500 B.n349 B.n348 585
R501 B.n350 B.n349 585
R502 B.n216 B.n215 585
R503 B.n217 B.n216 585
R504 B.n358 B.n357 585
R505 B.n357 B.n356 585
R506 B.n359 B.n214 585
R507 B.n214 B.n213 585
R508 B.n361 B.n360 585
R509 B.n362 B.n361 585
R510 B.n208 B.n207 585
R511 B.n209 B.n208 585
R512 B.n370 B.n369 585
R513 B.n369 B.n368 585
R514 B.n371 B.n206 585
R515 B.n206 B.n204 585
R516 B.n373 B.n372 585
R517 B.n374 B.n373 585
R518 B.n200 B.n199 585
R519 B.n205 B.n200 585
R520 B.n382 B.n381 585
R521 B.n381 B.n380 585
R522 B.n383 B.n198 585
R523 B.n198 B.n197 585
R524 B.n385 B.n384 585
R525 B.n386 B.n385 585
R526 B.n192 B.n191 585
R527 B.n193 B.n192 585
R528 B.n394 B.n393 585
R529 B.n393 B.n392 585
R530 B.n395 B.n190 585
R531 B.n190 B.n189 585
R532 B.n397 B.n396 585
R533 B.n398 B.n397 585
R534 B.n184 B.n183 585
R535 B.n185 B.n184 585
R536 B.n406 B.n405 585
R537 B.n405 B.n404 585
R538 B.n407 B.n182 585
R539 B.n182 B.n181 585
R540 B.n409 B.n408 585
R541 B.n410 B.n409 585
R542 B.n176 B.n175 585
R543 B.n177 B.n176 585
R544 B.n418 B.n417 585
R545 B.n417 B.n416 585
R546 B.n419 B.n174 585
R547 B.n174 B.n173 585
R548 B.n421 B.n420 585
R549 B.n422 B.n421 585
R550 B.n168 B.n167 585
R551 B.n169 B.n168 585
R552 B.n431 B.n430 585
R553 B.n430 B.n429 585
R554 B.n432 B.n166 585
R555 B.n166 B.n165 585
R556 B.n434 B.n433 585
R557 B.n435 B.n434 585
R558 B.n3 B.n0 585
R559 B.n4 B.n3 585
R560 B.n561 B.n1 585
R561 B.n562 B.n561 585
R562 B.n560 B.n559 585
R563 B.n560 B.n8 585
R564 B.n558 B.n9 585
R565 B.n444 B.n9 585
R566 B.n557 B.n556 585
R567 B.n556 B.n555 585
R568 B.n11 B.n10 585
R569 B.n554 B.n11 585
R570 B.n552 B.n551 585
R571 B.n553 B.n552 585
R572 B.n550 B.n16 585
R573 B.n16 B.n15 585
R574 B.n549 B.n548 585
R575 B.n548 B.n547 585
R576 B.n18 B.n17 585
R577 B.n546 B.n18 585
R578 B.n544 B.n543 585
R579 B.n545 B.n544 585
R580 B.n542 B.n23 585
R581 B.n23 B.n22 585
R582 B.n541 B.n540 585
R583 B.n540 B.n539 585
R584 B.n25 B.n24 585
R585 B.n538 B.n25 585
R586 B.n536 B.n535 585
R587 B.n537 B.n536 585
R588 B.n534 B.n30 585
R589 B.n30 B.n29 585
R590 B.n533 B.n532 585
R591 B.n532 B.n531 585
R592 B.n32 B.n31 585
R593 B.n530 B.n32 585
R594 B.n528 B.n527 585
R595 B.n529 B.n528 585
R596 B.n526 B.n37 585
R597 B.n37 B.n36 585
R598 B.n525 B.n524 585
R599 B.n524 B.n523 585
R600 B.n39 B.n38 585
R601 B.n522 B.n39 585
R602 B.n520 B.n519 585
R603 B.n521 B.n520 585
R604 B.n518 B.n44 585
R605 B.n44 B.n43 585
R606 B.n517 B.n516 585
R607 B.n516 B.n515 585
R608 B.n46 B.n45 585
R609 B.n514 B.n46 585
R610 B.n512 B.n511 585
R611 B.n513 B.n512 585
R612 B.n510 B.n51 585
R613 B.n51 B.n50 585
R614 B.n509 B.n508 585
R615 B.n508 B.n507 585
R616 B.n53 B.n52 585
R617 B.n506 B.n53 585
R618 B.n504 B.n503 585
R619 B.n505 B.n504 585
R620 B.n502 B.n58 585
R621 B.n58 B.n57 585
R622 B.n501 B.n500 585
R623 B.n500 B.n499 585
R624 B.n60 B.n59 585
R625 B.n498 B.n60 585
R626 B.n496 B.n495 585
R627 B.n497 B.n496 585
R628 B.n494 B.n65 585
R629 B.n65 B.n64 585
R630 B.n493 B.n492 585
R631 B.n492 B.n491 585
R632 B.n565 B.n564 585
R633 B.n563 B.n2 585
R634 B.n492 B.n67 434.841
R635 B.n489 B.n68 434.841
R636 B.n331 B.n234 434.841
R637 B.n333 B.n232 434.841
R638 B.n490 B.n86 256.663
R639 B.n490 B.n85 256.663
R640 B.n490 B.n84 256.663
R641 B.n490 B.n83 256.663
R642 B.n490 B.n82 256.663
R643 B.n490 B.n81 256.663
R644 B.n490 B.n80 256.663
R645 B.n490 B.n79 256.663
R646 B.n490 B.n78 256.663
R647 B.n490 B.n77 256.663
R648 B.n490 B.n76 256.663
R649 B.n490 B.n75 256.663
R650 B.n490 B.n74 256.663
R651 B.n490 B.n73 256.663
R652 B.n490 B.n72 256.663
R653 B.n490 B.n71 256.663
R654 B.n490 B.n70 256.663
R655 B.n490 B.n69 256.663
R656 B.n256 B.n233 256.663
R657 B.n259 B.n233 256.663
R658 B.n265 B.n233 256.663
R659 B.n267 B.n233 256.663
R660 B.n273 B.n233 256.663
R661 B.n275 B.n233 256.663
R662 B.n284 B.n233 256.663
R663 B.n286 B.n233 256.663
R664 B.n292 B.n233 256.663
R665 B.n294 B.n233 256.663
R666 B.n300 B.n233 256.663
R667 B.n302 B.n233 256.663
R668 B.n308 B.n233 256.663
R669 B.n310 B.n233 256.663
R670 B.n316 B.n233 256.663
R671 B.n318 B.n233 256.663
R672 B.n324 B.n233 256.663
R673 B.n326 B.n233 256.663
R674 B.n567 B.n566 256.663
R675 B.n90 B.t19 242.593
R676 B.n88 B.t12 242.593
R677 B.n241 B.t8 242.593
R678 B.n279 B.t16 242.593
R679 B.n95 B.n94 163.367
R680 B.n99 B.n98 163.367
R681 B.n103 B.n102 163.367
R682 B.n107 B.n106 163.367
R683 B.n111 B.n110 163.367
R684 B.n115 B.n114 163.367
R685 B.n119 B.n118 163.367
R686 B.n123 B.n122 163.367
R687 B.n127 B.n126 163.367
R688 B.n131 B.n130 163.367
R689 B.n135 B.n134 163.367
R690 B.n140 B.n139 163.367
R691 B.n144 B.n143 163.367
R692 B.n148 B.n147 163.367
R693 B.n152 B.n151 163.367
R694 B.n156 B.n155 163.367
R695 B.n160 B.n159 163.367
R696 B.n489 B.n87 163.367
R697 B.n331 B.n228 163.367
R698 B.n339 B.n228 163.367
R699 B.n339 B.n226 163.367
R700 B.n343 B.n226 163.367
R701 B.n343 B.n220 163.367
R702 B.n351 B.n220 163.367
R703 B.n351 B.n218 163.367
R704 B.n355 B.n218 163.367
R705 B.n355 B.n212 163.367
R706 B.n363 B.n212 163.367
R707 B.n363 B.n210 163.367
R708 B.n367 B.n210 163.367
R709 B.n367 B.n203 163.367
R710 B.n375 B.n203 163.367
R711 B.n375 B.n201 163.367
R712 B.n379 B.n201 163.367
R713 B.n379 B.n196 163.367
R714 B.n387 B.n196 163.367
R715 B.n387 B.n194 163.367
R716 B.n391 B.n194 163.367
R717 B.n391 B.n188 163.367
R718 B.n399 B.n188 163.367
R719 B.n399 B.n186 163.367
R720 B.n403 B.n186 163.367
R721 B.n403 B.n180 163.367
R722 B.n411 B.n180 163.367
R723 B.n411 B.n178 163.367
R724 B.n415 B.n178 163.367
R725 B.n415 B.n172 163.367
R726 B.n423 B.n172 163.367
R727 B.n423 B.n170 163.367
R728 B.n428 B.n170 163.367
R729 B.n428 B.n164 163.367
R730 B.n436 B.n164 163.367
R731 B.n437 B.n436 163.367
R732 B.n437 B.n5 163.367
R733 B.n6 B.n5 163.367
R734 B.n7 B.n6 163.367
R735 B.n443 B.n7 163.367
R736 B.n445 B.n443 163.367
R737 B.n445 B.n12 163.367
R738 B.n13 B.n12 163.367
R739 B.n14 B.n13 163.367
R740 B.n450 B.n14 163.367
R741 B.n450 B.n19 163.367
R742 B.n20 B.n19 163.367
R743 B.n21 B.n20 163.367
R744 B.n455 B.n21 163.367
R745 B.n455 B.n26 163.367
R746 B.n27 B.n26 163.367
R747 B.n28 B.n27 163.367
R748 B.n460 B.n28 163.367
R749 B.n460 B.n33 163.367
R750 B.n34 B.n33 163.367
R751 B.n35 B.n34 163.367
R752 B.n465 B.n35 163.367
R753 B.n465 B.n40 163.367
R754 B.n41 B.n40 163.367
R755 B.n42 B.n41 163.367
R756 B.n470 B.n42 163.367
R757 B.n470 B.n47 163.367
R758 B.n48 B.n47 163.367
R759 B.n49 B.n48 163.367
R760 B.n475 B.n49 163.367
R761 B.n475 B.n54 163.367
R762 B.n55 B.n54 163.367
R763 B.n56 B.n55 163.367
R764 B.n480 B.n56 163.367
R765 B.n480 B.n61 163.367
R766 B.n62 B.n61 163.367
R767 B.n63 B.n62 163.367
R768 B.n485 B.n63 163.367
R769 B.n485 B.n68 163.367
R770 B.n258 B.n257 163.367
R771 B.n260 B.n258 163.367
R772 B.n264 B.n253 163.367
R773 B.n268 B.n266 163.367
R774 B.n272 B.n251 163.367
R775 B.n276 B.n274 163.367
R776 B.n283 B.n249 163.367
R777 B.n287 B.n285 163.367
R778 B.n291 B.n247 163.367
R779 B.n295 B.n293 163.367
R780 B.n299 B.n245 163.367
R781 B.n303 B.n301 163.367
R782 B.n307 B.n240 163.367
R783 B.n311 B.n309 163.367
R784 B.n315 B.n238 163.367
R785 B.n319 B.n317 163.367
R786 B.n323 B.n236 163.367
R787 B.n327 B.n325 163.367
R788 B.n333 B.n230 163.367
R789 B.n337 B.n230 163.367
R790 B.n337 B.n224 163.367
R791 B.n345 B.n224 163.367
R792 B.n345 B.n222 163.367
R793 B.n349 B.n222 163.367
R794 B.n349 B.n216 163.367
R795 B.n357 B.n216 163.367
R796 B.n357 B.n214 163.367
R797 B.n361 B.n214 163.367
R798 B.n361 B.n208 163.367
R799 B.n369 B.n208 163.367
R800 B.n369 B.n206 163.367
R801 B.n373 B.n206 163.367
R802 B.n373 B.n200 163.367
R803 B.n381 B.n200 163.367
R804 B.n381 B.n198 163.367
R805 B.n385 B.n198 163.367
R806 B.n385 B.n192 163.367
R807 B.n393 B.n192 163.367
R808 B.n393 B.n190 163.367
R809 B.n397 B.n190 163.367
R810 B.n397 B.n184 163.367
R811 B.n405 B.n184 163.367
R812 B.n405 B.n182 163.367
R813 B.n409 B.n182 163.367
R814 B.n409 B.n176 163.367
R815 B.n417 B.n176 163.367
R816 B.n417 B.n174 163.367
R817 B.n421 B.n174 163.367
R818 B.n421 B.n168 163.367
R819 B.n430 B.n168 163.367
R820 B.n430 B.n166 163.367
R821 B.n434 B.n166 163.367
R822 B.n434 B.n3 163.367
R823 B.n565 B.n3 163.367
R824 B.n561 B.n2 163.367
R825 B.n561 B.n560 163.367
R826 B.n560 B.n9 163.367
R827 B.n556 B.n9 163.367
R828 B.n556 B.n11 163.367
R829 B.n552 B.n11 163.367
R830 B.n552 B.n16 163.367
R831 B.n548 B.n16 163.367
R832 B.n548 B.n18 163.367
R833 B.n544 B.n18 163.367
R834 B.n544 B.n23 163.367
R835 B.n540 B.n23 163.367
R836 B.n540 B.n25 163.367
R837 B.n536 B.n25 163.367
R838 B.n536 B.n30 163.367
R839 B.n532 B.n30 163.367
R840 B.n532 B.n32 163.367
R841 B.n528 B.n32 163.367
R842 B.n528 B.n37 163.367
R843 B.n524 B.n37 163.367
R844 B.n524 B.n39 163.367
R845 B.n520 B.n39 163.367
R846 B.n520 B.n44 163.367
R847 B.n516 B.n44 163.367
R848 B.n516 B.n46 163.367
R849 B.n512 B.n46 163.367
R850 B.n512 B.n51 163.367
R851 B.n508 B.n51 163.367
R852 B.n508 B.n53 163.367
R853 B.n504 B.n53 163.367
R854 B.n504 B.n58 163.367
R855 B.n500 B.n58 163.367
R856 B.n500 B.n60 163.367
R857 B.n496 B.n60 163.367
R858 B.n496 B.n65 163.367
R859 B.n492 B.n65 163.367
R860 B.n332 B.n233 161.325
R861 B.n491 B.n490 161.325
R862 B.n88 B.t14 158.577
R863 B.n241 B.t11 158.577
R864 B.n90 B.t20 158.577
R865 B.n279 B.t18 158.577
R866 B.n89 B.t15 121.341
R867 B.n242 B.t10 121.341
R868 B.n91 B.t21 121.341
R869 B.n280 B.t17 121.341
R870 B.n332 B.n229 97.0803
R871 B.n338 B.n229 97.0803
R872 B.n338 B.n225 97.0803
R873 B.n344 B.n225 97.0803
R874 B.n344 B.n221 97.0803
R875 B.n350 B.n221 97.0803
R876 B.n356 B.n217 97.0803
R877 B.n356 B.n213 97.0803
R878 B.n362 B.n213 97.0803
R879 B.n362 B.n209 97.0803
R880 B.n368 B.n209 97.0803
R881 B.n368 B.n204 97.0803
R882 B.n374 B.n204 97.0803
R883 B.n374 B.n205 97.0803
R884 B.n380 B.n197 97.0803
R885 B.n386 B.n197 97.0803
R886 B.n386 B.n193 97.0803
R887 B.n392 B.n193 97.0803
R888 B.n398 B.n189 97.0803
R889 B.n398 B.n185 97.0803
R890 B.n404 B.n185 97.0803
R891 B.n404 B.n181 97.0803
R892 B.n410 B.n181 97.0803
R893 B.n416 B.n177 97.0803
R894 B.n416 B.n173 97.0803
R895 B.n422 B.n173 97.0803
R896 B.n422 B.n169 97.0803
R897 B.n429 B.n169 97.0803
R898 B.n435 B.n165 97.0803
R899 B.n435 B.n4 97.0803
R900 B.n564 B.n4 97.0803
R901 B.n564 B.n563 97.0803
R902 B.n563 B.n562 97.0803
R903 B.n562 B.n8 97.0803
R904 B.n444 B.n8 97.0803
R905 B.n555 B.n554 97.0803
R906 B.n554 B.n553 97.0803
R907 B.n553 B.n15 97.0803
R908 B.n547 B.n15 97.0803
R909 B.n547 B.n546 97.0803
R910 B.n545 B.n22 97.0803
R911 B.n539 B.n22 97.0803
R912 B.n539 B.n538 97.0803
R913 B.n538 B.n537 97.0803
R914 B.n537 B.n29 97.0803
R915 B.n531 B.n530 97.0803
R916 B.n530 B.n529 97.0803
R917 B.n529 B.n36 97.0803
R918 B.n523 B.n36 97.0803
R919 B.n522 B.n521 97.0803
R920 B.n521 B.n43 97.0803
R921 B.n515 B.n43 97.0803
R922 B.n515 B.n514 97.0803
R923 B.n514 B.n513 97.0803
R924 B.n513 B.n50 97.0803
R925 B.n507 B.n50 97.0803
R926 B.n507 B.n506 97.0803
R927 B.n505 B.n57 97.0803
R928 B.n499 B.n57 97.0803
R929 B.n499 B.n498 97.0803
R930 B.n498 B.n497 97.0803
R931 B.n497 B.n64 97.0803
R932 B.n491 B.n64 97.0803
R933 B.t2 B.n165 89.9421
R934 B.n444 B.t5 89.9421
R935 B.n380 B.t3 84.2315
R936 B.n523 B.t7 84.2315
R937 B.n392 B.t4 75.6657
R938 B.n531 B.t1 75.6657
R939 B.n69 B.n67 71.676
R940 B.n95 B.n70 71.676
R941 B.n99 B.n71 71.676
R942 B.n103 B.n72 71.676
R943 B.n107 B.n73 71.676
R944 B.n111 B.n74 71.676
R945 B.n115 B.n75 71.676
R946 B.n119 B.n76 71.676
R947 B.n123 B.n77 71.676
R948 B.n127 B.n78 71.676
R949 B.n131 B.n79 71.676
R950 B.n135 B.n80 71.676
R951 B.n140 B.n81 71.676
R952 B.n144 B.n82 71.676
R953 B.n148 B.n83 71.676
R954 B.n152 B.n84 71.676
R955 B.n156 B.n85 71.676
R956 B.n160 B.n86 71.676
R957 B.n87 B.n86 71.676
R958 B.n159 B.n85 71.676
R959 B.n155 B.n84 71.676
R960 B.n151 B.n83 71.676
R961 B.n147 B.n82 71.676
R962 B.n143 B.n81 71.676
R963 B.n139 B.n80 71.676
R964 B.n134 B.n79 71.676
R965 B.n130 B.n78 71.676
R966 B.n126 B.n77 71.676
R967 B.n122 B.n76 71.676
R968 B.n118 B.n75 71.676
R969 B.n114 B.n74 71.676
R970 B.n110 B.n73 71.676
R971 B.n106 B.n72 71.676
R972 B.n102 B.n71 71.676
R973 B.n98 B.n70 71.676
R974 B.n94 B.n69 71.676
R975 B.n256 B.n232 71.676
R976 B.n260 B.n259 71.676
R977 B.n265 B.n264 71.676
R978 B.n268 B.n267 71.676
R979 B.n273 B.n272 71.676
R980 B.n276 B.n275 71.676
R981 B.n284 B.n283 71.676
R982 B.n287 B.n286 71.676
R983 B.n292 B.n291 71.676
R984 B.n295 B.n294 71.676
R985 B.n300 B.n299 71.676
R986 B.n303 B.n302 71.676
R987 B.n308 B.n307 71.676
R988 B.n311 B.n310 71.676
R989 B.n316 B.n315 71.676
R990 B.n319 B.n318 71.676
R991 B.n324 B.n323 71.676
R992 B.n327 B.n326 71.676
R993 B.n257 B.n256 71.676
R994 B.n259 B.n253 71.676
R995 B.n266 B.n265 71.676
R996 B.n267 B.n251 71.676
R997 B.n274 B.n273 71.676
R998 B.n275 B.n249 71.676
R999 B.n285 B.n284 71.676
R1000 B.n286 B.n247 71.676
R1001 B.n293 B.n292 71.676
R1002 B.n294 B.n245 71.676
R1003 B.n301 B.n300 71.676
R1004 B.n302 B.n240 71.676
R1005 B.n309 B.n308 71.676
R1006 B.n310 B.n238 71.676
R1007 B.n317 B.n316 71.676
R1008 B.n318 B.n236 71.676
R1009 B.n325 B.n324 71.676
R1010 B.n326 B.n234 71.676
R1011 B.n566 B.n565 71.676
R1012 B.n566 B.n2 71.676
R1013 B.t9 B.n217 69.9551
R1014 B.n506 B.t13 69.9551
R1015 B.n92 B.n91 59.5399
R1016 B.n137 B.n89 59.5399
R1017 B.n243 B.n242 59.5399
R1018 B.n281 B.n280 59.5399
R1019 B.t6 B.n177 55.6786
R1020 B.n546 B.t0 55.6786
R1021 B.n410 B.t6 41.4022
R1022 B.t0 B.n545 41.4022
R1023 B.n91 B.n90 37.2369
R1024 B.n89 B.n88 37.2369
R1025 B.n242 B.n241 37.2369
R1026 B.n280 B.n279 37.2369
R1027 B.n488 B.n487 28.2542
R1028 B.n334 B.n231 28.2542
R1029 B.n330 B.n329 28.2542
R1030 B.n493 B.n66 28.2542
R1031 B.n350 B.t9 27.1257
R1032 B.t13 B.n505 27.1257
R1033 B.t4 B.n189 21.4152
R1034 B.t1 B.n29 21.4152
R1035 B B.n567 18.0485
R1036 B.n205 B.t3 12.8493
R1037 B.t7 B.n522 12.8493
R1038 B.n335 B.n334 10.6151
R1039 B.n336 B.n335 10.6151
R1040 B.n336 B.n223 10.6151
R1041 B.n346 B.n223 10.6151
R1042 B.n347 B.n346 10.6151
R1043 B.n348 B.n347 10.6151
R1044 B.n348 B.n215 10.6151
R1045 B.n358 B.n215 10.6151
R1046 B.n359 B.n358 10.6151
R1047 B.n360 B.n359 10.6151
R1048 B.n360 B.n207 10.6151
R1049 B.n370 B.n207 10.6151
R1050 B.n371 B.n370 10.6151
R1051 B.n372 B.n371 10.6151
R1052 B.n372 B.n199 10.6151
R1053 B.n382 B.n199 10.6151
R1054 B.n383 B.n382 10.6151
R1055 B.n384 B.n383 10.6151
R1056 B.n384 B.n191 10.6151
R1057 B.n394 B.n191 10.6151
R1058 B.n395 B.n394 10.6151
R1059 B.n396 B.n395 10.6151
R1060 B.n396 B.n183 10.6151
R1061 B.n406 B.n183 10.6151
R1062 B.n407 B.n406 10.6151
R1063 B.n408 B.n407 10.6151
R1064 B.n408 B.n175 10.6151
R1065 B.n418 B.n175 10.6151
R1066 B.n419 B.n418 10.6151
R1067 B.n420 B.n419 10.6151
R1068 B.n420 B.n167 10.6151
R1069 B.n431 B.n167 10.6151
R1070 B.n432 B.n431 10.6151
R1071 B.n433 B.n432 10.6151
R1072 B.n433 B.n0 10.6151
R1073 B.n255 B.n231 10.6151
R1074 B.n255 B.n254 10.6151
R1075 B.n261 B.n254 10.6151
R1076 B.n262 B.n261 10.6151
R1077 B.n263 B.n262 10.6151
R1078 B.n263 B.n252 10.6151
R1079 B.n269 B.n252 10.6151
R1080 B.n270 B.n269 10.6151
R1081 B.n271 B.n270 10.6151
R1082 B.n271 B.n250 10.6151
R1083 B.n277 B.n250 10.6151
R1084 B.n278 B.n277 10.6151
R1085 B.n282 B.n278 10.6151
R1086 B.n288 B.n248 10.6151
R1087 B.n289 B.n288 10.6151
R1088 B.n290 B.n289 10.6151
R1089 B.n290 B.n246 10.6151
R1090 B.n296 B.n246 10.6151
R1091 B.n297 B.n296 10.6151
R1092 B.n298 B.n297 10.6151
R1093 B.n298 B.n244 10.6151
R1094 B.n305 B.n304 10.6151
R1095 B.n306 B.n305 10.6151
R1096 B.n306 B.n239 10.6151
R1097 B.n312 B.n239 10.6151
R1098 B.n313 B.n312 10.6151
R1099 B.n314 B.n313 10.6151
R1100 B.n314 B.n237 10.6151
R1101 B.n320 B.n237 10.6151
R1102 B.n321 B.n320 10.6151
R1103 B.n322 B.n321 10.6151
R1104 B.n322 B.n235 10.6151
R1105 B.n328 B.n235 10.6151
R1106 B.n329 B.n328 10.6151
R1107 B.n330 B.n227 10.6151
R1108 B.n340 B.n227 10.6151
R1109 B.n341 B.n340 10.6151
R1110 B.n342 B.n341 10.6151
R1111 B.n342 B.n219 10.6151
R1112 B.n352 B.n219 10.6151
R1113 B.n353 B.n352 10.6151
R1114 B.n354 B.n353 10.6151
R1115 B.n354 B.n211 10.6151
R1116 B.n364 B.n211 10.6151
R1117 B.n365 B.n364 10.6151
R1118 B.n366 B.n365 10.6151
R1119 B.n366 B.n202 10.6151
R1120 B.n376 B.n202 10.6151
R1121 B.n377 B.n376 10.6151
R1122 B.n378 B.n377 10.6151
R1123 B.n378 B.n195 10.6151
R1124 B.n388 B.n195 10.6151
R1125 B.n389 B.n388 10.6151
R1126 B.n390 B.n389 10.6151
R1127 B.n390 B.n187 10.6151
R1128 B.n400 B.n187 10.6151
R1129 B.n401 B.n400 10.6151
R1130 B.n402 B.n401 10.6151
R1131 B.n402 B.n179 10.6151
R1132 B.n412 B.n179 10.6151
R1133 B.n413 B.n412 10.6151
R1134 B.n414 B.n413 10.6151
R1135 B.n414 B.n171 10.6151
R1136 B.n424 B.n171 10.6151
R1137 B.n425 B.n424 10.6151
R1138 B.n427 B.n425 10.6151
R1139 B.n427 B.n426 10.6151
R1140 B.n426 B.n163 10.6151
R1141 B.n438 B.n163 10.6151
R1142 B.n439 B.n438 10.6151
R1143 B.n440 B.n439 10.6151
R1144 B.n441 B.n440 10.6151
R1145 B.n442 B.n441 10.6151
R1146 B.n446 B.n442 10.6151
R1147 B.n447 B.n446 10.6151
R1148 B.n448 B.n447 10.6151
R1149 B.n449 B.n448 10.6151
R1150 B.n451 B.n449 10.6151
R1151 B.n452 B.n451 10.6151
R1152 B.n453 B.n452 10.6151
R1153 B.n454 B.n453 10.6151
R1154 B.n456 B.n454 10.6151
R1155 B.n457 B.n456 10.6151
R1156 B.n458 B.n457 10.6151
R1157 B.n459 B.n458 10.6151
R1158 B.n461 B.n459 10.6151
R1159 B.n462 B.n461 10.6151
R1160 B.n463 B.n462 10.6151
R1161 B.n464 B.n463 10.6151
R1162 B.n466 B.n464 10.6151
R1163 B.n467 B.n466 10.6151
R1164 B.n468 B.n467 10.6151
R1165 B.n469 B.n468 10.6151
R1166 B.n471 B.n469 10.6151
R1167 B.n472 B.n471 10.6151
R1168 B.n473 B.n472 10.6151
R1169 B.n474 B.n473 10.6151
R1170 B.n476 B.n474 10.6151
R1171 B.n477 B.n476 10.6151
R1172 B.n478 B.n477 10.6151
R1173 B.n479 B.n478 10.6151
R1174 B.n481 B.n479 10.6151
R1175 B.n482 B.n481 10.6151
R1176 B.n483 B.n482 10.6151
R1177 B.n484 B.n483 10.6151
R1178 B.n486 B.n484 10.6151
R1179 B.n487 B.n486 10.6151
R1180 B.n559 B.n1 10.6151
R1181 B.n559 B.n558 10.6151
R1182 B.n558 B.n557 10.6151
R1183 B.n557 B.n10 10.6151
R1184 B.n551 B.n10 10.6151
R1185 B.n551 B.n550 10.6151
R1186 B.n550 B.n549 10.6151
R1187 B.n549 B.n17 10.6151
R1188 B.n543 B.n17 10.6151
R1189 B.n543 B.n542 10.6151
R1190 B.n542 B.n541 10.6151
R1191 B.n541 B.n24 10.6151
R1192 B.n535 B.n24 10.6151
R1193 B.n535 B.n534 10.6151
R1194 B.n534 B.n533 10.6151
R1195 B.n533 B.n31 10.6151
R1196 B.n527 B.n31 10.6151
R1197 B.n527 B.n526 10.6151
R1198 B.n526 B.n525 10.6151
R1199 B.n525 B.n38 10.6151
R1200 B.n519 B.n38 10.6151
R1201 B.n519 B.n518 10.6151
R1202 B.n518 B.n517 10.6151
R1203 B.n517 B.n45 10.6151
R1204 B.n511 B.n45 10.6151
R1205 B.n511 B.n510 10.6151
R1206 B.n510 B.n509 10.6151
R1207 B.n509 B.n52 10.6151
R1208 B.n503 B.n52 10.6151
R1209 B.n503 B.n502 10.6151
R1210 B.n502 B.n501 10.6151
R1211 B.n501 B.n59 10.6151
R1212 B.n495 B.n59 10.6151
R1213 B.n495 B.n494 10.6151
R1214 B.n494 B.n493 10.6151
R1215 B.n93 B.n66 10.6151
R1216 B.n96 B.n93 10.6151
R1217 B.n97 B.n96 10.6151
R1218 B.n100 B.n97 10.6151
R1219 B.n101 B.n100 10.6151
R1220 B.n104 B.n101 10.6151
R1221 B.n105 B.n104 10.6151
R1222 B.n108 B.n105 10.6151
R1223 B.n109 B.n108 10.6151
R1224 B.n112 B.n109 10.6151
R1225 B.n113 B.n112 10.6151
R1226 B.n116 B.n113 10.6151
R1227 B.n117 B.n116 10.6151
R1228 B.n121 B.n120 10.6151
R1229 B.n124 B.n121 10.6151
R1230 B.n125 B.n124 10.6151
R1231 B.n128 B.n125 10.6151
R1232 B.n129 B.n128 10.6151
R1233 B.n132 B.n129 10.6151
R1234 B.n133 B.n132 10.6151
R1235 B.n136 B.n133 10.6151
R1236 B.n141 B.n138 10.6151
R1237 B.n142 B.n141 10.6151
R1238 B.n145 B.n142 10.6151
R1239 B.n146 B.n145 10.6151
R1240 B.n149 B.n146 10.6151
R1241 B.n150 B.n149 10.6151
R1242 B.n153 B.n150 10.6151
R1243 B.n154 B.n153 10.6151
R1244 B.n157 B.n154 10.6151
R1245 B.n158 B.n157 10.6151
R1246 B.n161 B.n158 10.6151
R1247 B.n162 B.n161 10.6151
R1248 B.n488 B.n162 10.6151
R1249 B.n567 B.n0 8.11757
R1250 B.n567 B.n1 8.11757
R1251 B.n429 B.t2 7.13872
R1252 B.n555 B.t5 7.13872
R1253 B.n281 B.n248 6.5566
R1254 B.n244 B.n243 6.5566
R1255 B.n120 B.n92 6.5566
R1256 B.n137 B.n136 6.5566
R1257 B.n282 B.n281 4.05904
R1258 B.n304 B.n243 4.05904
R1259 B.n117 B.n92 4.05904
R1260 B.n138 B.n137 4.05904
R1261 VN.n20 VN.n19 179.406
R1262 VN.n41 VN.n40 179.406
R1263 VN.n39 VN.n21 161.3
R1264 VN.n38 VN.n37 161.3
R1265 VN.n36 VN.n22 161.3
R1266 VN.n35 VN.n34 161.3
R1267 VN.n32 VN.n23 161.3
R1268 VN.n31 VN.n30 161.3
R1269 VN.n29 VN.n24 161.3
R1270 VN.n28 VN.n27 161.3
R1271 VN.n18 VN.n0 161.3
R1272 VN.n17 VN.n16 161.3
R1273 VN.n15 VN.n1 161.3
R1274 VN.n14 VN.n13 161.3
R1275 VN.n11 VN.n2 161.3
R1276 VN.n10 VN.n9 161.3
R1277 VN.n8 VN.n3 161.3
R1278 VN.n7 VN.n6 161.3
R1279 VN.n4 VN.t6 68.617
R1280 VN.n25 VN.t4 68.617
R1281 VN.n17 VN.n1 56.5193
R1282 VN.n38 VN.n22 56.5193
R1283 VN.n10 VN.n3 56.5193
R1284 VN.n31 VN.n24 56.5193
R1285 VN.n5 VN.n4 55.7366
R1286 VN.n26 VN.n25 55.7366
R1287 VN VN.n41 39.1918
R1288 VN.n5 VN.t3 36.8326
R1289 VN.n12 VN.t1 36.8326
R1290 VN.n19 VN.t0 36.8326
R1291 VN.n26 VN.t7 36.8326
R1292 VN.n33 VN.t5 36.8326
R1293 VN.n40 VN.t2 36.8326
R1294 VN.n6 VN.n3 24.4675
R1295 VN.n11 VN.n10 24.4675
R1296 VN.n13 VN.n1 24.4675
R1297 VN.n18 VN.n17 24.4675
R1298 VN.n27 VN.n24 24.4675
R1299 VN.n34 VN.n22 24.4675
R1300 VN.n32 VN.n31 24.4675
R1301 VN.n39 VN.n38 24.4675
R1302 VN.n28 VN.n25 18.144
R1303 VN.n7 VN.n4 18.144
R1304 VN.n13 VN.n12 14.1914
R1305 VN.n34 VN.n33 14.1914
R1306 VN.n6 VN.n5 10.2766
R1307 VN.n12 VN.n11 10.2766
R1308 VN.n27 VN.n26 10.2766
R1309 VN.n33 VN.n32 10.2766
R1310 VN.n19 VN.n18 6.36192
R1311 VN.n40 VN.n39 6.36192
R1312 VN.n41 VN.n21 0.189894
R1313 VN.n37 VN.n21 0.189894
R1314 VN.n37 VN.n36 0.189894
R1315 VN.n36 VN.n35 0.189894
R1316 VN.n35 VN.n23 0.189894
R1317 VN.n30 VN.n23 0.189894
R1318 VN.n30 VN.n29 0.189894
R1319 VN.n29 VN.n28 0.189894
R1320 VN.n8 VN.n7 0.189894
R1321 VN.n9 VN.n8 0.189894
R1322 VN.n9 VN.n2 0.189894
R1323 VN.n14 VN.n2 0.189894
R1324 VN.n15 VN.n14 0.189894
R1325 VN.n16 VN.n15 0.189894
R1326 VN.n16 VN.n0 0.189894
R1327 VN.n20 VN.n0 0.189894
R1328 VN VN.n20 0.0516364
R1329 VDD2.n2 VDD2.n1 86.3132
R1330 VDD2.n2 VDD2.n0 86.3132
R1331 VDD2 VDD2.n5 86.3104
R1332 VDD2.n4 VDD2.n3 85.5411
R1333 VDD2.n4 VDD2.n2 33.2584
R1334 VDD2.n5 VDD2.t0 8.14865
R1335 VDD2.n5 VDD2.t3 8.14865
R1336 VDD2.n3 VDD2.t5 8.14865
R1337 VDD2.n3 VDD2.t2 8.14865
R1338 VDD2.n1 VDD2.t6 8.14865
R1339 VDD2.n1 VDD2.t7 8.14865
R1340 VDD2.n0 VDD2.t1 8.14865
R1341 VDD2.n0 VDD2.t4 8.14865
R1342 VDD2 VDD2.n4 0.886276
C0 VN VP 4.66297f
C1 VDD2 VP 0.418501f
C2 VTAIL VP 2.54699f
C3 VDD2 VN 1.89511f
C4 VDD1 VP 2.15637f
C5 VTAIL VN 2.53289f
C6 VDD2 VTAIL 4.14009f
C7 VDD1 VN 0.155385f
C8 VDD2 VDD1 1.2552f
C9 VDD1 VTAIL 4.09245f
C10 VDD2 B 3.434032f
C11 VDD1 B 3.935894f
C12 VTAIL B 3.821585f
C13 VN B 10.46622f
C14 VP B 9.276098f
C15 VDD2.t1 B 0.03196f
C16 VDD2.t4 B 0.03196f
C17 VDD2.n0 B 0.228409f
C18 VDD2.t6 B 0.03196f
C19 VDD2.t7 B 0.03196f
C20 VDD2.n1 B 0.228409f
C21 VDD2.n2 B 1.3783f
C22 VDD2.t5 B 0.03196f
C23 VDD2.t2 B 0.03196f
C24 VDD2.n3 B 0.226104f
C25 VDD2.n4 B 1.21114f
C26 VDD2.t0 B 0.03196f
C27 VDD2.t3 B 0.03196f
C28 VDD2.n5 B 0.228395f
C29 VN.n0 B 0.028302f
C30 VN.t0 B 0.264418f
C31 VN.n1 B 0.035007f
C32 VN.n2 B 0.028302f
C33 VN.t1 B 0.264418f
C34 VN.n3 B 0.041316f
C35 VN.t6 B 0.376712f
C36 VN.n4 B 0.181629f
C37 VN.t3 B 0.264418f
C38 VN.n5 B 0.181111f
C39 VN.n6 B 0.037644f
C40 VN.n7 B 0.179403f
C41 VN.n8 B 0.028302f
C42 VN.n9 B 0.028302f
C43 VN.n10 B 0.041316f
C44 VN.n11 B 0.037644f
C45 VN.n12 B 0.128194f
C46 VN.n13 B 0.041811f
C47 VN.n14 B 0.028302f
C48 VN.n15 B 0.028302f
C49 VN.n16 B 0.028302f
C50 VN.n17 B 0.047626f
C51 VN.n18 B 0.033477f
C52 VN.n19 B 0.185922f
C53 VN.n20 B 0.028413f
C54 VN.n21 B 0.028302f
C55 VN.t2 B 0.264418f
C56 VN.n22 B 0.035007f
C57 VN.n23 B 0.028302f
C58 VN.t5 B 0.264418f
C59 VN.n24 B 0.041316f
C60 VN.t4 B 0.376712f
C61 VN.n25 B 0.181629f
C62 VN.t7 B 0.264418f
C63 VN.n26 B 0.181111f
C64 VN.n27 B 0.037644f
C65 VN.n28 B 0.179403f
C66 VN.n29 B 0.028302f
C67 VN.n30 B 0.028302f
C68 VN.n31 B 0.041316f
C69 VN.n32 B 0.037644f
C70 VN.n33 B 0.128194f
C71 VN.n34 B 0.041811f
C72 VN.n35 B 0.028302f
C73 VN.n36 B 0.028302f
C74 VN.n37 B 0.028302f
C75 VN.n38 B 0.047626f
C76 VN.n39 B 0.033477f
C77 VN.n40 B 0.185922f
C78 VN.n41 B 1.04549f
C79 VDD1.t1 B 0.048384f
C80 VDD1.t2 B 0.048384f
C81 VDD1.n0 B 0.346382f
C82 VDD1.t0 B 0.048384f
C83 VDD1.t7 B 0.048384f
C84 VDD1.n1 B 0.345786f
C85 VDD1.t6 B 0.048384f
C86 VDD1.t5 B 0.048384f
C87 VDD1.n2 B 0.345786f
C88 VDD1.n3 B 2.13993f
C89 VDD1.t3 B 0.048384f
C90 VDD1.t4 B 0.048384f
C91 VDD1.n4 B 0.342295f
C92 VDD1.n5 B 1.86381f
C93 VTAIL.t0 B 0.052284f
C94 VTAIL.t1 B 0.052284f
C95 VTAIL.n0 B 0.323454f
C96 VTAIL.n1 B 0.356634f
C97 VTAIL.n2 B 0.035148f
C98 VTAIL.n3 B 0.198373f
C99 VTAIL.n4 B 0.014631f
C100 VTAIL.t5 B 0.05893f
C101 VTAIL.n5 B 0.094099f
C102 VTAIL.n6 B 0.019576f
C103 VTAIL.n7 B 0.025937f
C104 VTAIL.n8 B 0.069343f
C105 VTAIL.n9 B 0.015492f
C106 VTAIL.n10 B 0.014631f
C107 VTAIL.n11 B 0.064052f
C108 VTAIL.n12 B 0.038266f
C109 VTAIL.n13 B 0.210319f
C110 VTAIL.n14 B 0.035148f
C111 VTAIL.n15 B 0.198373f
C112 VTAIL.n16 B 0.014631f
C113 VTAIL.t11 B 0.05893f
C114 VTAIL.n17 B 0.094099f
C115 VTAIL.n18 B 0.019576f
C116 VTAIL.n19 B 0.025937f
C117 VTAIL.n20 B 0.069343f
C118 VTAIL.n21 B 0.015492f
C119 VTAIL.n22 B 0.014631f
C120 VTAIL.n23 B 0.064052f
C121 VTAIL.n24 B 0.038266f
C122 VTAIL.n25 B 0.210319f
C123 VTAIL.t14 B 0.052284f
C124 VTAIL.t15 B 0.052284f
C125 VTAIL.n26 B 0.323454f
C126 VTAIL.n27 B 0.496743f
C127 VTAIL.n28 B 0.035148f
C128 VTAIL.n29 B 0.198373f
C129 VTAIL.n30 B 0.014631f
C130 VTAIL.t8 B 0.05893f
C131 VTAIL.n31 B 0.094099f
C132 VTAIL.n32 B 0.019576f
C133 VTAIL.n33 B 0.025937f
C134 VTAIL.n34 B 0.069343f
C135 VTAIL.n35 B 0.015492f
C136 VTAIL.n36 B 0.014631f
C137 VTAIL.n37 B 0.064052f
C138 VTAIL.n38 B 0.038266f
C139 VTAIL.n39 B 0.867959f
C140 VTAIL.n40 B 0.035148f
C141 VTAIL.n41 B 0.198373f
C142 VTAIL.n42 B 0.014631f
C143 VTAIL.t3 B 0.05893f
C144 VTAIL.n43 B 0.094099f
C145 VTAIL.n44 B 0.019576f
C146 VTAIL.n45 B 0.025937f
C147 VTAIL.n46 B 0.069343f
C148 VTAIL.n47 B 0.015492f
C149 VTAIL.n48 B 0.014631f
C150 VTAIL.n49 B 0.064052f
C151 VTAIL.n50 B 0.038266f
C152 VTAIL.n51 B 0.867959f
C153 VTAIL.t4 B 0.052284f
C154 VTAIL.t6 B 0.052284f
C155 VTAIL.n52 B 0.323457f
C156 VTAIL.n53 B 0.496741f
C157 VTAIL.n54 B 0.035148f
C158 VTAIL.n55 B 0.198373f
C159 VTAIL.n56 B 0.014631f
C160 VTAIL.t2 B 0.05893f
C161 VTAIL.n57 B 0.094099f
C162 VTAIL.n58 B 0.019576f
C163 VTAIL.n59 B 0.025937f
C164 VTAIL.n60 B 0.069343f
C165 VTAIL.n61 B 0.015492f
C166 VTAIL.n62 B 0.014631f
C167 VTAIL.n63 B 0.064052f
C168 VTAIL.n64 B 0.038266f
C169 VTAIL.n65 B 0.210319f
C170 VTAIL.n66 B 0.035148f
C171 VTAIL.n67 B 0.198373f
C172 VTAIL.n68 B 0.014631f
C173 VTAIL.t9 B 0.05893f
C174 VTAIL.n69 B 0.094099f
C175 VTAIL.n70 B 0.019576f
C176 VTAIL.n71 B 0.025937f
C177 VTAIL.n72 B 0.069343f
C178 VTAIL.n73 B 0.015492f
C179 VTAIL.n74 B 0.014631f
C180 VTAIL.n75 B 0.064052f
C181 VTAIL.n76 B 0.038266f
C182 VTAIL.n77 B 0.210319f
C183 VTAIL.t10 B 0.052284f
C184 VTAIL.t12 B 0.052284f
C185 VTAIL.n78 B 0.323457f
C186 VTAIL.n79 B 0.496741f
C187 VTAIL.n80 B 0.035148f
C188 VTAIL.n81 B 0.198373f
C189 VTAIL.n82 B 0.014631f
C190 VTAIL.t13 B 0.05893f
C191 VTAIL.n83 B 0.094099f
C192 VTAIL.n84 B 0.019576f
C193 VTAIL.n85 B 0.025937f
C194 VTAIL.n86 B 0.069343f
C195 VTAIL.n87 B 0.015492f
C196 VTAIL.n88 B 0.014631f
C197 VTAIL.n89 B 0.064052f
C198 VTAIL.n90 B 0.038266f
C199 VTAIL.n91 B 0.867959f
C200 VTAIL.n92 B 0.035148f
C201 VTAIL.n93 B 0.198373f
C202 VTAIL.n94 B 0.014631f
C203 VTAIL.t7 B 0.05893f
C204 VTAIL.n95 B 0.094099f
C205 VTAIL.n96 B 0.019576f
C206 VTAIL.n97 B 0.025937f
C207 VTAIL.n98 B 0.069343f
C208 VTAIL.n99 B 0.015492f
C209 VTAIL.n100 B 0.014631f
C210 VTAIL.n101 B 0.064052f
C211 VTAIL.n102 B 0.038266f
C212 VTAIL.n103 B 0.862854f
C213 VP.n0 B 0.037156f
C214 VP.t2 B 0.34713f
C215 VP.n1 B 0.045957f
C216 VP.n2 B 0.037156f
C217 VP.t1 B 0.34713f
C218 VP.n3 B 0.054241f
C219 VP.n4 B 0.037156f
C220 VP.t0 B 0.34713f
C221 VP.n5 B 0.062524f
C222 VP.n6 B 0.037156f
C223 VP.t3 B 0.34713f
C224 VP.n7 B 0.045957f
C225 VP.n8 B 0.037156f
C226 VP.t4 B 0.34713f
C227 VP.n9 B 0.054241f
C228 VP.t6 B 0.494552f
C229 VP.n10 B 0.238444f
C230 VP.t5 B 0.34713f
C231 VP.n11 B 0.237764f
C232 VP.n12 B 0.049419f
C233 VP.n13 B 0.235523f
C234 VP.n14 B 0.037156f
C235 VP.n15 B 0.037156f
C236 VP.n16 B 0.054241f
C237 VP.n17 B 0.049419f
C238 VP.n18 B 0.168294f
C239 VP.n19 B 0.05489f
C240 VP.n20 B 0.037156f
C241 VP.n21 B 0.037156f
C242 VP.n22 B 0.037156f
C243 VP.n23 B 0.062524f
C244 VP.n24 B 0.043949f
C245 VP.n25 B 0.24408f
C246 VP.n26 B 1.34802f
C247 VP.n27 B 1.38243f
C248 VP.t7 B 0.34713f
C249 VP.n28 B 0.24408f
C250 VP.n29 B 0.043949f
C251 VP.n30 B 0.037156f
C252 VP.n31 B 0.037156f
C253 VP.n32 B 0.037156f
C254 VP.n33 B 0.045957f
C255 VP.n34 B 0.05489f
C256 VP.n35 B 0.168294f
C257 VP.n36 B 0.049419f
C258 VP.n37 B 0.037156f
C259 VP.n38 B 0.037156f
C260 VP.n39 B 0.037156f
C261 VP.n40 B 0.054241f
C262 VP.n41 B 0.049419f
C263 VP.n42 B 0.168294f
C264 VP.n43 B 0.05489f
C265 VP.n44 B 0.037156f
C266 VP.n45 B 0.037156f
C267 VP.n46 B 0.037156f
C268 VP.n47 B 0.062524f
C269 VP.n48 B 0.043949f
C270 VP.n49 B 0.24408f
C271 VP.n50 B 0.037301f
.ends

