* NGSPICE file created from diff_pair_sample_0702.ext - technology: sky130A

.subckt diff_pair_sample_0702 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=2.21595 ps=13.76 w=13.43 l=1.01
X1 VDD2.t9 VN.t0 VTAIL.t3 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X2 VDD2.t8 VN.t1 VTAIL.t5 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X3 VDD2.t7 VN.t2 VTAIL.t4 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=2.21595 ps=13.76 w=13.43 l=1.01
X4 VTAIL.t9 VN.t3 VDD2.t6 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X5 VTAIL.t2 VN.t4 VDD2.t5 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X6 VTAIL.t17 VP.t1 VDD1.t8 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X7 VDD2.t4 VN.t5 VTAIL.t1 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=2.21595 ps=13.76 w=13.43 l=1.01
X8 B.t11 B.t9 B.t10 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=0 ps=0 w=13.43 l=1.01
X9 VDD2.t3 VN.t6 VTAIL.t0 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=5.2377 ps=27.64 w=13.43 l=1.01
X10 B.t8 B.t6 B.t7 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=0 ps=0 w=13.43 l=1.01
X11 VDD2.t2 VN.t7 VTAIL.t8 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=5.2377 ps=27.64 w=13.43 l=1.01
X12 VTAIL.t15 VP.t2 VDD1.t7 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X13 VDD1.t6 VP.t3 VTAIL.t16 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=2.21595 ps=13.76 w=13.43 l=1.01
X14 B.t5 B.t3 B.t4 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=0 ps=0 w=13.43 l=1.01
X15 VDD1.t5 VP.t4 VTAIL.t13 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=5.2377 ps=27.64 w=13.43 l=1.01
X16 VTAIL.t7 VN.t8 VDD2.t1 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X17 VDD1.t4 VP.t5 VTAIL.t11 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X18 VTAIL.t10 VP.t6 VDD1.t3 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X19 VDD1.t2 VP.t7 VTAIL.t12 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=5.2377 ps=27.64 w=13.43 l=1.01
X20 VTAIL.t19 VP.t8 VDD1.t1 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X21 B.t2 B.t0 B.t1 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=5.2377 pd=27.64 as=0 ps=0 w=13.43 l=1.01
X22 VDD1.t0 VP.t9 VTAIL.t14 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
X23 VTAIL.t6 VN.t9 VDD2.t0 w_n2578_n3654# sky130_fd_pr__pfet_01v8 ad=2.21595 pd=13.76 as=2.21595 ps=13.76 w=13.43 l=1.01
R0 VP.n9 VP.t0 374.082
R1 VP.n25 VP.t3 359.591
R2 VP.n41 VP.t4 359.591
R3 VP.n22 VP.t7 359.591
R4 VP.n26 VP.t8 320.459
R5 VP.n33 VP.t5 320.459
R6 VP.n39 VP.t6 320.459
R7 VP.n20 VP.t1 320.459
R8 VP.n14 VP.t9 320.459
R9 VP.n8 VP.t2 320.459
R10 VP.n10 VP.n7 161.3
R11 VP.n12 VP.n11 161.3
R12 VP.n13 VP.n6 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n5 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n21 VP.n4 161.3
R17 VP.n40 VP.n0 161.3
R18 VP.n38 VP.n37 161.3
R19 VP.n36 VP.n1 161.3
R20 VP.n35 VP.n34 161.3
R21 VP.n32 VP.n2 161.3
R22 VP.n31 VP.n30 161.3
R23 VP.n29 VP.n3 161.3
R24 VP.n28 VP.n27 161.3
R25 VP.n23 VP.n22 80.6037
R26 VP.n42 VP.n41 80.6037
R27 VP.n25 VP.n24 80.6037
R28 VP.n27 VP.n25 52.8492
R29 VP.n41 VP.n40 52.8492
R30 VP.n22 VP.n21 52.8492
R31 VP.n9 VP.n8 48.957
R32 VP.n32 VP.n31 48.2635
R33 VP.n34 VP.n1 48.2635
R34 VP.n15 VP.n5 48.2635
R35 VP.n13 VP.n12 48.2635
R36 VP.n24 VP.n23 45.7211
R37 VP.n10 VP.n9 44.4127
R38 VP.n31 VP.n3 32.7233
R39 VP.n38 VP.n1 32.7233
R40 VP.n19 VP.n5 32.7233
R41 VP.n12 VP.n7 32.7233
R42 VP.n27 VP.n26 20.0634
R43 VP.n40 VP.n39 20.0634
R44 VP.n21 VP.n20 20.0634
R45 VP.n33 VP.n32 12.234
R46 VP.n34 VP.n33 12.234
R47 VP.n14 VP.n13 12.234
R48 VP.n15 VP.n14 12.234
R49 VP.n26 VP.n3 4.40456
R50 VP.n39 VP.n38 4.40456
R51 VP.n20 VP.n19 4.40456
R52 VP.n8 VP.n7 4.40456
R53 VP.n23 VP.n4 0.285035
R54 VP.n28 VP.n24 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n11 VP.n10 0.189894
R57 VP.n11 VP.n6 0.189894
R58 VP.n16 VP.n6 0.189894
R59 VP.n17 VP.n16 0.189894
R60 VP.n18 VP.n17 0.189894
R61 VP.n18 VP.n4 0.189894
R62 VP.n29 VP.n28 0.189894
R63 VP.n30 VP.n29 0.189894
R64 VP.n30 VP.n2 0.189894
R65 VP.n35 VP.n2 0.189894
R66 VP.n36 VP.n35 0.189894
R67 VP.n37 VP.n36 0.189894
R68 VP.n37 VP.n0 0.189894
R69 VP VP.n42 0.146778
R70 VTAIL.n255 VTAIL.n254 585
R71 VTAIL.n257 VTAIL.n256 585
R72 VTAIL.n250 VTAIL.n249 585
R73 VTAIL.n263 VTAIL.n262 585
R74 VTAIL.n265 VTAIL.n264 585
R75 VTAIL.n246 VTAIL.n245 585
R76 VTAIL.n271 VTAIL.n270 585
R77 VTAIL.n273 VTAIL.n272 585
R78 VTAIL.n242 VTAIL.n241 585
R79 VTAIL.n279 VTAIL.n278 585
R80 VTAIL.n281 VTAIL.n280 585
R81 VTAIL.n238 VTAIL.n237 585
R82 VTAIL.n287 VTAIL.n286 585
R83 VTAIL.n289 VTAIL.n288 585
R84 VTAIL.n234 VTAIL.n233 585
R85 VTAIL.n295 VTAIL.n294 585
R86 VTAIL.n297 VTAIL.n296 585
R87 VTAIL.n27 VTAIL.n26 585
R88 VTAIL.n29 VTAIL.n28 585
R89 VTAIL.n22 VTAIL.n21 585
R90 VTAIL.n35 VTAIL.n34 585
R91 VTAIL.n37 VTAIL.n36 585
R92 VTAIL.n18 VTAIL.n17 585
R93 VTAIL.n43 VTAIL.n42 585
R94 VTAIL.n45 VTAIL.n44 585
R95 VTAIL.n14 VTAIL.n13 585
R96 VTAIL.n51 VTAIL.n50 585
R97 VTAIL.n53 VTAIL.n52 585
R98 VTAIL.n10 VTAIL.n9 585
R99 VTAIL.n59 VTAIL.n58 585
R100 VTAIL.n61 VTAIL.n60 585
R101 VTAIL.n6 VTAIL.n5 585
R102 VTAIL.n67 VTAIL.n66 585
R103 VTAIL.n69 VTAIL.n68 585
R104 VTAIL.n225 VTAIL.n224 585
R105 VTAIL.n223 VTAIL.n222 585
R106 VTAIL.n162 VTAIL.n161 585
R107 VTAIL.n217 VTAIL.n216 585
R108 VTAIL.n215 VTAIL.n214 585
R109 VTAIL.n166 VTAIL.n165 585
R110 VTAIL.n209 VTAIL.n208 585
R111 VTAIL.n207 VTAIL.n206 585
R112 VTAIL.n170 VTAIL.n169 585
R113 VTAIL.n201 VTAIL.n200 585
R114 VTAIL.n199 VTAIL.n198 585
R115 VTAIL.n174 VTAIL.n173 585
R116 VTAIL.n193 VTAIL.n192 585
R117 VTAIL.n191 VTAIL.n190 585
R118 VTAIL.n178 VTAIL.n177 585
R119 VTAIL.n185 VTAIL.n184 585
R120 VTAIL.n183 VTAIL.n182 585
R121 VTAIL.n149 VTAIL.n148 585
R122 VTAIL.n147 VTAIL.n146 585
R123 VTAIL.n86 VTAIL.n85 585
R124 VTAIL.n141 VTAIL.n140 585
R125 VTAIL.n139 VTAIL.n138 585
R126 VTAIL.n90 VTAIL.n89 585
R127 VTAIL.n133 VTAIL.n132 585
R128 VTAIL.n131 VTAIL.n130 585
R129 VTAIL.n94 VTAIL.n93 585
R130 VTAIL.n125 VTAIL.n124 585
R131 VTAIL.n123 VTAIL.n122 585
R132 VTAIL.n98 VTAIL.n97 585
R133 VTAIL.n117 VTAIL.n116 585
R134 VTAIL.n115 VTAIL.n114 585
R135 VTAIL.n102 VTAIL.n101 585
R136 VTAIL.n109 VTAIL.n108 585
R137 VTAIL.n107 VTAIL.n106 585
R138 VTAIL.n296 VTAIL.n230 498.474
R139 VTAIL.n68 VTAIL.n2 498.474
R140 VTAIL.n224 VTAIL.n158 498.474
R141 VTAIL.n148 VTAIL.n82 498.474
R142 VTAIL.n253 VTAIL.t0 327.466
R143 VTAIL.n25 VTAIL.t13 327.466
R144 VTAIL.n181 VTAIL.t12 327.466
R145 VTAIL.n105 VTAIL.t8 327.466
R146 VTAIL.n256 VTAIL.n255 171.744
R147 VTAIL.n256 VTAIL.n249 171.744
R148 VTAIL.n263 VTAIL.n249 171.744
R149 VTAIL.n264 VTAIL.n263 171.744
R150 VTAIL.n264 VTAIL.n245 171.744
R151 VTAIL.n271 VTAIL.n245 171.744
R152 VTAIL.n272 VTAIL.n271 171.744
R153 VTAIL.n272 VTAIL.n241 171.744
R154 VTAIL.n279 VTAIL.n241 171.744
R155 VTAIL.n280 VTAIL.n279 171.744
R156 VTAIL.n280 VTAIL.n237 171.744
R157 VTAIL.n287 VTAIL.n237 171.744
R158 VTAIL.n288 VTAIL.n287 171.744
R159 VTAIL.n288 VTAIL.n233 171.744
R160 VTAIL.n295 VTAIL.n233 171.744
R161 VTAIL.n296 VTAIL.n295 171.744
R162 VTAIL.n28 VTAIL.n27 171.744
R163 VTAIL.n28 VTAIL.n21 171.744
R164 VTAIL.n35 VTAIL.n21 171.744
R165 VTAIL.n36 VTAIL.n35 171.744
R166 VTAIL.n36 VTAIL.n17 171.744
R167 VTAIL.n43 VTAIL.n17 171.744
R168 VTAIL.n44 VTAIL.n43 171.744
R169 VTAIL.n44 VTAIL.n13 171.744
R170 VTAIL.n51 VTAIL.n13 171.744
R171 VTAIL.n52 VTAIL.n51 171.744
R172 VTAIL.n52 VTAIL.n9 171.744
R173 VTAIL.n59 VTAIL.n9 171.744
R174 VTAIL.n60 VTAIL.n59 171.744
R175 VTAIL.n60 VTAIL.n5 171.744
R176 VTAIL.n67 VTAIL.n5 171.744
R177 VTAIL.n68 VTAIL.n67 171.744
R178 VTAIL.n224 VTAIL.n223 171.744
R179 VTAIL.n223 VTAIL.n161 171.744
R180 VTAIL.n216 VTAIL.n161 171.744
R181 VTAIL.n216 VTAIL.n215 171.744
R182 VTAIL.n215 VTAIL.n165 171.744
R183 VTAIL.n208 VTAIL.n165 171.744
R184 VTAIL.n208 VTAIL.n207 171.744
R185 VTAIL.n207 VTAIL.n169 171.744
R186 VTAIL.n200 VTAIL.n169 171.744
R187 VTAIL.n200 VTAIL.n199 171.744
R188 VTAIL.n199 VTAIL.n173 171.744
R189 VTAIL.n192 VTAIL.n173 171.744
R190 VTAIL.n192 VTAIL.n191 171.744
R191 VTAIL.n191 VTAIL.n177 171.744
R192 VTAIL.n184 VTAIL.n177 171.744
R193 VTAIL.n184 VTAIL.n183 171.744
R194 VTAIL.n148 VTAIL.n147 171.744
R195 VTAIL.n147 VTAIL.n85 171.744
R196 VTAIL.n140 VTAIL.n85 171.744
R197 VTAIL.n140 VTAIL.n139 171.744
R198 VTAIL.n139 VTAIL.n89 171.744
R199 VTAIL.n132 VTAIL.n89 171.744
R200 VTAIL.n132 VTAIL.n131 171.744
R201 VTAIL.n131 VTAIL.n93 171.744
R202 VTAIL.n124 VTAIL.n93 171.744
R203 VTAIL.n124 VTAIL.n123 171.744
R204 VTAIL.n123 VTAIL.n97 171.744
R205 VTAIL.n116 VTAIL.n97 171.744
R206 VTAIL.n116 VTAIL.n115 171.744
R207 VTAIL.n115 VTAIL.n101 171.744
R208 VTAIL.n108 VTAIL.n101 171.744
R209 VTAIL.n108 VTAIL.n107 171.744
R210 VTAIL.n255 VTAIL.t0 85.8723
R211 VTAIL.n27 VTAIL.t13 85.8723
R212 VTAIL.n183 VTAIL.t12 85.8723
R213 VTAIL.n107 VTAIL.t8 85.8723
R214 VTAIL.n157 VTAIL.n156 59.7484
R215 VTAIL.n155 VTAIL.n154 59.7484
R216 VTAIL.n81 VTAIL.n80 59.7484
R217 VTAIL.n79 VTAIL.n78 59.7484
R218 VTAIL.n303 VTAIL.n302 59.7482
R219 VTAIL.n1 VTAIL.n0 59.7482
R220 VTAIL.n75 VTAIL.n74 59.7482
R221 VTAIL.n77 VTAIL.n76 59.7482
R222 VTAIL.n301 VTAIL.n300 36.646
R223 VTAIL.n73 VTAIL.n72 36.646
R224 VTAIL.n229 VTAIL.n228 36.646
R225 VTAIL.n153 VTAIL.n152 36.646
R226 VTAIL.n79 VTAIL.n77 26.2548
R227 VTAIL.n301 VTAIL.n229 25.0996
R228 VTAIL.n254 VTAIL.n253 16.3895
R229 VTAIL.n26 VTAIL.n25 16.3895
R230 VTAIL.n182 VTAIL.n181 16.3895
R231 VTAIL.n106 VTAIL.n105 16.3895
R232 VTAIL.n257 VTAIL.n252 12.8005
R233 VTAIL.n298 VTAIL.n297 12.8005
R234 VTAIL.n29 VTAIL.n24 12.8005
R235 VTAIL.n70 VTAIL.n69 12.8005
R236 VTAIL.n226 VTAIL.n225 12.8005
R237 VTAIL.n185 VTAIL.n180 12.8005
R238 VTAIL.n150 VTAIL.n149 12.8005
R239 VTAIL.n109 VTAIL.n104 12.8005
R240 VTAIL.n258 VTAIL.n250 12.0247
R241 VTAIL.n294 VTAIL.n232 12.0247
R242 VTAIL.n30 VTAIL.n22 12.0247
R243 VTAIL.n66 VTAIL.n4 12.0247
R244 VTAIL.n222 VTAIL.n160 12.0247
R245 VTAIL.n186 VTAIL.n178 12.0247
R246 VTAIL.n146 VTAIL.n84 12.0247
R247 VTAIL.n110 VTAIL.n102 12.0247
R248 VTAIL.n262 VTAIL.n261 11.249
R249 VTAIL.n293 VTAIL.n234 11.249
R250 VTAIL.n34 VTAIL.n33 11.249
R251 VTAIL.n65 VTAIL.n6 11.249
R252 VTAIL.n221 VTAIL.n162 11.249
R253 VTAIL.n190 VTAIL.n189 11.249
R254 VTAIL.n145 VTAIL.n86 11.249
R255 VTAIL.n114 VTAIL.n113 11.249
R256 VTAIL.n265 VTAIL.n248 10.4732
R257 VTAIL.n290 VTAIL.n289 10.4732
R258 VTAIL.n37 VTAIL.n20 10.4732
R259 VTAIL.n62 VTAIL.n61 10.4732
R260 VTAIL.n218 VTAIL.n217 10.4732
R261 VTAIL.n193 VTAIL.n176 10.4732
R262 VTAIL.n142 VTAIL.n141 10.4732
R263 VTAIL.n117 VTAIL.n100 10.4732
R264 VTAIL.n266 VTAIL.n246 9.69747
R265 VTAIL.n286 VTAIL.n236 9.69747
R266 VTAIL.n38 VTAIL.n18 9.69747
R267 VTAIL.n58 VTAIL.n8 9.69747
R268 VTAIL.n214 VTAIL.n164 9.69747
R269 VTAIL.n194 VTAIL.n174 9.69747
R270 VTAIL.n138 VTAIL.n88 9.69747
R271 VTAIL.n118 VTAIL.n98 9.69747
R272 VTAIL.n300 VTAIL.n299 9.45567
R273 VTAIL.n72 VTAIL.n71 9.45567
R274 VTAIL.n228 VTAIL.n227 9.45567
R275 VTAIL.n152 VTAIL.n151 9.45567
R276 VTAIL.n275 VTAIL.n274 9.3005
R277 VTAIL.n244 VTAIL.n243 9.3005
R278 VTAIL.n269 VTAIL.n268 9.3005
R279 VTAIL.n267 VTAIL.n266 9.3005
R280 VTAIL.n248 VTAIL.n247 9.3005
R281 VTAIL.n261 VTAIL.n260 9.3005
R282 VTAIL.n259 VTAIL.n258 9.3005
R283 VTAIL.n252 VTAIL.n251 9.3005
R284 VTAIL.n277 VTAIL.n276 9.3005
R285 VTAIL.n240 VTAIL.n239 9.3005
R286 VTAIL.n283 VTAIL.n282 9.3005
R287 VTAIL.n285 VTAIL.n284 9.3005
R288 VTAIL.n236 VTAIL.n235 9.3005
R289 VTAIL.n291 VTAIL.n290 9.3005
R290 VTAIL.n293 VTAIL.n292 9.3005
R291 VTAIL.n232 VTAIL.n231 9.3005
R292 VTAIL.n299 VTAIL.n298 9.3005
R293 VTAIL.n47 VTAIL.n46 9.3005
R294 VTAIL.n16 VTAIL.n15 9.3005
R295 VTAIL.n41 VTAIL.n40 9.3005
R296 VTAIL.n39 VTAIL.n38 9.3005
R297 VTAIL.n20 VTAIL.n19 9.3005
R298 VTAIL.n33 VTAIL.n32 9.3005
R299 VTAIL.n31 VTAIL.n30 9.3005
R300 VTAIL.n24 VTAIL.n23 9.3005
R301 VTAIL.n49 VTAIL.n48 9.3005
R302 VTAIL.n12 VTAIL.n11 9.3005
R303 VTAIL.n55 VTAIL.n54 9.3005
R304 VTAIL.n57 VTAIL.n56 9.3005
R305 VTAIL.n8 VTAIL.n7 9.3005
R306 VTAIL.n63 VTAIL.n62 9.3005
R307 VTAIL.n65 VTAIL.n64 9.3005
R308 VTAIL.n4 VTAIL.n3 9.3005
R309 VTAIL.n71 VTAIL.n70 9.3005
R310 VTAIL.n168 VTAIL.n167 9.3005
R311 VTAIL.n211 VTAIL.n210 9.3005
R312 VTAIL.n213 VTAIL.n212 9.3005
R313 VTAIL.n164 VTAIL.n163 9.3005
R314 VTAIL.n219 VTAIL.n218 9.3005
R315 VTAIL.n221 VTAIL.n220 9.3005
R316 VTAIL.n160 VTAIL.n159 9.3005
R317 VTAIL.n227 VTAIL.n226 9.3005
R318 VTAIL.n205 VTAIL.n204 9.3005
R319 VTAIL.n203 VTAIL.n202 9.3005
R320 VTAIL.n172 VTAIL.n171 9.3005
R321 VTAIL.n197 VTAIL.n196 9.3005
R322 VTAIL.n195 VTAIL.n194 9.3005
R323 VTAIL.n176 VTAIL.n175 9.3005
R324 VTAIL.n189 VTAIL.n188 9.3005
R325 VTAIL.n187 VTAIL.n186 9.3005
R326 VTAIL.n180 VTAIL.n179 9.3005
R327 VTAIL.n92 VTAIL.n91 9.3005
R328 VTAIL.n135 VTAIL.n134 9.3005
R329 VTAIL.n137 VTAIL.n136 9.3005
R330 VTAIL.n88 VTAIL.n87 9.3005
R331 VTAIL.n143 VTAIL.n142 9.3005
R332 VTAIL.n145 VTAIL.n144 9.3005
R333 VTAIL.n84 VTAIL.n83 9.3005
R334 VTAIL.n151 VTAIL.n150 9.3005
R335 VTAIL.n129 VTAIL.n128 9.3005
R336 VTAIL.n127 VTAIL.n126 9.3005
R337 VTAIL.n96 VTAIL.n95 9.3005
R338 VTAIL.n121 VTAIL.n120 9.3005
R339 VTAIL.n119 VTAIL.n118 9.3005
R340 VTAIL.n100 VTAIL.n99 9.3005
R341 VTAIL.n113 VTAIL.n112 9.3005
R342 VTAIL.n111 VTAIL.n110 9.3005
R343 VTAIL.n104 VTAIL.n103 9.3005
R344 VTAIL.n270 VTAIL.n269 8.92171
R345 VTAIL.n285 VTAIL.n238 8.92171
R346 VTAIL.n42 VTAIL.n41 8.92171
R347 VTAIL.n57 VTAIL.n10 8.92171
R348 VTAIL.n213 VTAIL.n166 8.92171
R349 VTAIL.n198 VTAIL.n197 8.92171
R350 VTAIL.n137 VTAIL.n90 8.92171
R351 VTAIL.n122 VTAIL.n121 8.92171
R352 VTAIL.n273 VTAIL.n244 8.14595
R353 VTAIL.n282 VTAIL.n281 8.14595
R354 VTAIL.n45 VTAIL.n16 8.14595
R355 VTAIL.n54 VTAIL.n53 8.14595
R356 VTAIL.n210 VTAIL.n209 8.14595
R357 VTAIL.n201 VTAIL.n172 8.14595
R358 VTAIL.n134 VTAIL.n133 8.14595
R359 VTAIL.n125 VTAIL.n96 8.14595
R360 VTAIL.n300 VTAIL.n230 7.75445
R361 VTAIL.n72 VTAIL.n2 7.75445
R362 VTAIL.n228 VTAIL.n158 7.75445
R363 VTAIL.n152 VTAIL.n82 7.75445
R364 VTAIL.n274 VTAIL.n242 7.3702
R365 VTAIL.n278 VTAIL.n240 7.3702
R366 VTAIL.n46 VTAIL.n14 7.3702
R367 VTAIL.n50 VTAIL.n12 7.3702
R368 VTAIL.n206 VTAIL.n168 7.3702
R369 VTAIL.n202 VTAIL.n170 7.3702
R370 VTAIL.n130 VTAIL.n92 7.3702
R371 VTAIL.n126 VTAIL.n94 7.3702
R372 VTAIL.n277 VTAIL.n242 6.59444
R373 VTAIL.n278 VTAIL.n277 6.59444
R374 VTAIL.n49 VTAIL.n14 6.59444
R375 VTAIL.n50 VTAIL.n49 6.59444
R376 VTAIL.n206 VTAIL.n205 6.59444
R377 VTAIL.n205 VTAIL.n170 6.59444
R378 VTAIL.n130 VTAIL.n129 6.59444
R379 VTAIL.n129 VTAIL.n94 6.59444
R380 VTAIL.n298 VTAIL.n230 6.08283
R381 VTAIL.n70 VTAIL.n2 6.08283
R382 VTAIL.n226 VTAIL.n158 6.08283
R383 VTAIL.n150 VTAIL.n82 6.08283
R384 VTAIL.n274 VTAIL.n273 5.81868
R385 VTAIL.n281 VTAIL.n240 5.81868
R386 VTAIL.n46 VTAIL.n45 5.81868
R387 VTAIL.n53 VTAIL.n12 5.81868
R388 VTAIL.n209 VTAIL.n168 5.81868
R389 VTAIL.n202 VTAIL.n201 5.81868
R390 VTAIL.n133 VTAIL.n92 5.81868
R391 VTAIL.n126 VTAIL.n125 5.81868
R392 VTAIL.n270 VTAIL.n244 5.04292
R393 VTAIL.n282 VTAIL.n238 5.04292
R394 VTAIL.n42 VTAIL.n16 5.04292
R395 VTAIL.n54 VTAIL.n10 5.04292
R396 VTAIL.n210 VTAIL.n166 5.04292
R397 VTAIL.n198 VTAIL.n172 5.04292
R398 VTAIL.n134 VTAIL.n90 5.04292
R399 VTAIL.n122 VTAIL.n96 5.04292
R400 VTAIL.n269 VTAIL.n246 4.26717
R401 VTAIL.n286 VTAIL.n285 4.26717
R402 VTAIL.n41 VTAIL.n18 4.26717
R403 VTAIL.n58 VTAIL.n57 4.26717
R404 VTAIL.n214 VTAIL.n213 4.26717
R405 VTAIL.n197 VTAIL.n174 4.26717
R406 VTAIL.n138 VTAIL.n137 4.26717
R407 VTAIL.n121 VTAIL.n98 4.26717
R408 VTAIL.n253 VTAIL.n251 3.70982
R409 VTAIL.n25 VTAIL.n23 3.70982
R410 VTAIL.n181 VTAIL.n179 3.70982
R411 VTAIL.n105 VTAIL.n103 3.70982
R412 VTAIL.n266 VTAIL.n265 3.49141
R413 VTAIL.n289 VTAIL.n236 3.49141
R414 VTAIL.n38 VTAIL.n37 3.49141
R415 VTAIL.n61 VTAIL.n8 3.49141
R416 VTAIL.n217 VTAIL.n164 3.49141
R417 VTAIL.n194 VTAIL.n193 3.49141
R418 VTAIL.n141 VTAIL.n88 3.49141
R419 VTAIL.n118 VTAIL.n117 3.49141
R420 VTAIL.n262 VTAIL.n248 2.71565
R421 VTAIL.n290 VTAIL.n234 2.71565
R422 VTAIL.n34 VTAIL.n20 2.71565
R423 VTAIL.n62 VTAIL.n6 2.71565
R424 VTAIL.n218 VTAIL.n162 2.71565
R425 VTAIL.n190 VTAIL.n176 2.71565
R426 VTAIL.n142 VTAIL.n86 2.71565
R427 VTAIL.n114 VTAIL.n100 2.71565
R428 VTAIL.n302 VTAIL.t5 2.42083
R429 VTAIL.n302 VTAIL.t9 2.42083
R430 VTAIL.n0 VTAIL.t4 2.42083
R431 VTAIL.n0 VTAIL.t2 2.42083
R432 VTAIL.n74 VTAIL.t11 2.42083
R433 VTAIL.n74 VTAIL.t10 2.42083
R434 VTAIL.n76 VTAIL.t16 2.42083
R435 VTAIL.n76 VTAIL.t19 2.42083
R436 VTAIL.n156 VTAIL.t14 2.42083
R437 VTAIL.n156 VTAIL.t17 2.42083
R438 VTAIL.n154 VTAIL.t18 2.42083
R439 VTAIL.n154 VTAIL.t15 2.42083
R440 VTAIL.n80 VTAIL.t3 2.42083
R441 VTAIL.n80 VTAIL.t6 2.42083
R442 VTAIL.n78 VTAIL.t1 2.42083
R443 VTAIL.n78 VTAIL.t7 2.42083
R444 VTAIL.n261 VTAIL.n250 1.93989
R445 VTAIL.n294 VTAIL.n293 1.93989
R446 VTAIL.n33 VTAIL.n22 1.93989
R447 VTAIL.n66 VTAIL.n65 1.93989
R448 VTAIL.n222 VTAIL.n221 1.93989
R449 VTAIL.n189 VTAIL.n178 1.93989
R450 VTAIL.n146 VTAIL.n145 1.93989
R451 VTAIL.n113 VTAIL.n102 1.93989
R452 VTAIL.n258 VTAIL.n257 1.16414
R453 VTAIL.n297 VTAIL.n232 1.16414
R454 VTAIL.n30 VTAIL.n29 1.16414
R455 VTAIL.n69 VTAIL.n4 1.16414
R456 VTAIL.n225 VTAIL.n160 1.16414
R457 VTAIL.n186 VTAIL.n185 1.16414
R458 VTAIL.n149 VTAIL.n84 1.16414
R459 VTAIL.n110 VTAIL.n109 1.16414
R460 VTAIL.n81 VTAIL.n79 1.15567
R461 VTAIL.n153 VTAIL.n81 1.15567
R462 VTAIL.n157 VTAIL.n155 1.15567
R463 VTAIL.n229 VTAIL.n157 1.15567
R464 VTAIL.n77 VTAIL.n75 1.15567
R465 VTAIL.n75 VTAIL.n73 1.15567
R466 VTAIL.n303 VTAIL.n301 1.15567
R467 VTAIL.n155 VTAIL.n153 1.04791
R468 VTAIL.n73 VTAIL.n1 1.04791
R469 VTAIL VTAIL.n1 0.925069
R470 VTAIL.n254 VTAIL.n252 0.388379
R471 VTAIL.n26 VTAIL.n24 0.388379
R472 VTAIL.n182 VTAIL.n180 0.388379
R473 VTAIL.n106 VTAIL.n104 0.388379
R474 VTAIL VTAIL.n303 0.231103
R475 VTAIL.n259 VTAIL.n251 0.155672
R476 VTAIL.n260 VTAIL.n259 0.155672
R477 VTAIL.n260 VTAIL.n247 0.155672
R478 VTAIL.n267 VTAIL.n247 0.155672
R479 VTAIL.n268 VTAIL.n267 0.155672
R480 VTAIL.n268 VTAIL.n243 0.155672
R481 VTAIL.n275 VTAIL.n243 0.155672
R482 VTAIL.n276 VTAIL.n275 0.155672
R483 VTAIL.n276 VTAIL.n239 0.155672
R484 VTAIL.n283 VTAIL.n239 0.155672
R485 VTAIL.n284 VTAIL.n283 0.155672
R486 VTAIL.n284 VTAIL.n235 0.155672
R487 VTAIL.n291 VTAIL.n235 0.155672
R488 VTAIL.n292 VTAIL.n291 0.155672
R489 VTAIL.n292 VTAIL.n231 0.155672
R490 VTAIL.n299 VTAIL.n231 0.155672
R491 VTAIL.n31 VTAIL.n23 0.155672
R492 VTAIL.n32 VTAIL.n31 0.155672
R493 VTAIL.n32 VTAIL.n19 0.155672
R494 VTAIL.n39 VTAIL.n19 0.155672
R495 VTAIL.n40 VTAIL.n39 0.155672
R496 VTAIL.n40 VTAIL.n15 0.155672
R497 VTAIL.n47 VTAIL.n15 0.155672
R498 VTAIL.n48 VTAIL.n47 0.155672
R499 VTAIL.n48 VTAIL.n11 0.155672
R500 VTAIL.n55 VTAIL.n11 0.155672
R501 VTAIL.n56 VTAIL.n55 0.155672
R502 VTAIL.n56 VTAIL.n7 0.155672
R503 VTAIL.n63 VTAIL.n7 0.155672
R504 VTAIL.n64 VTAIL.n63 0.155672
R505 VTAIL.n64 VTAIL.n3 0.155672
R506 VTAIL.n71 VTAIL.n3 0.155672
R507 VTAIL.n227 VTAIL.n159 0.155672
R508 VTAIL.n220 VTAIL.n159 0.155672
R509 VTAIL.n220 VTAIL.n219 0.155672
R510 VTAIL.n219 VTAIL.n163 0.155672
R511 VTAIL.n212 VTAIL.n163 0.155672
R512 VTAIL.n212 VTAIL.n211 0.155672
R513 VTAIL.n211 VTAIL.n167 0.155672
R514 VTAIL.n204 VTAIL.n167 0.155672
R515 VTAIL.n204 VTAIL.n203 0.155672
R516 VTAIL.n203 VTAIL.n171 0.155672
R517 VTAIL.n196 VTAIL.n171 0.155672
R518 VTAIL.n196 VTAIL.n195 0.155672
R519 VTAIL.n195 VTAIL.n175 0.155672
R520 VTAIL.n188 VTAIL.n175 0.155672
R521 VTAIL.n188 VTAIL.n187 0.155672
R522 VTAIL.n187 VTAIL.n179 0.155672
R523 VTAIL.n151 VTAIL.n83 0.155672
R524 VTAIL.n144 VTAIL.n83 0.155672
R525 VTAIL.n144 VTAIL.n143 0.155672
R526 VTAIL.n143 VTAIL.n87 0.155672
R527 VTAIL.n136 VTAIL.n87 0.155672
R528 VTAIL.n136 VTAIL.n135 0.155672
R529 VTAIL.n135 VTAIL.n91 0.155672
R530 VTAIL.n128 VTAIL.n91 0.155672
R531 VTAIL.n128 VTAIL.n127 0.155672
R532 VTAIL.n127 VTAIL.n95 0.155672
R533 VTAIL.n120 VTAIL.n95 0.155672
R534 VTAIL.n120 VTAIL.n119 0.155672
R535 VTAIL.n119 VTAIL.n99 0.155672
R536 VTAIL.n112 VTAIL.n99 0.155672
R537 VTAIL.n112 VTAIL.n111 0.155672
R538 VTAIL.n111 VTAIL.n103 0.155672
R539 VDD1.n67 VDD1.n66 585
R540 VDD1.n65 VDD1.n64 585
R541 VDD1.n4 VDD1.n3 585
R542 VDD1.n59 VDD1.n58 585
R543 VDD1.n57 VDD1.n56 585
R544 VDD1.n8 VDD1.n7 585
R545 VDD1.n51 VDD1.n50 585
R546 VDD1.n49 VDD1.n48 585
R547 VDD1.n12 VDD1.n11 585
R548 VDD1.n43 VDD1.n42 585
R549 VDD1.n41 VDD1.n40 585
R550 VDD1.n16 VDD1.n15 585
R551 VDD1.n35 VDD1.n34 585
R552 VDD1.n33 VDD1.n32 585
R553 VDD1.n20 VDD1.n19 585
R554 VDD1.n27 VDD1.n26 585
R555 VDD1.n25 VDD1.n24 585
R556 VDD1.n98 VDD1.n97 585
R557 VDD1.n100 VDD1.n99 585
R558 VDD1.n93 VDD1.n92 585
R559 VDD1.n106 VDD1.n105 585
R560 VDD1.n108 VDD1.n107 585
R561 VDD1.n89 VDD1.n88 585
R562 VDD1.n114 VDD1.n113 585
R563 VDD1.n116 VDD1.n115 585
R564 VDD1.n85 VDD1.n84 585
R565 VDD1.n122 VDD1.n121 585
R566 VDD1.n124 VDD1.n123 585
R567 VDD1.n81 VDD1.n80 585
R568 VDD1.n130 VDD1.n129 585
R569 VDD1.n132 VDD1.n131 585
R570 VDD1.n77 VDD1.n76 585
R571 VDD1.n138 VDD1.n137 585
R572 VDD1.n140 VDD1.n139 585
R573 VDD1.n66 VDD1.n0 498.474
R574 VDD1.n139 VDD1.n73 498.474
R575 VDD1.n23 VDD1.t9 327.466
R576 VDD1.n96 VDD1.t6 327.466
R577 VDD1.n66 VDD1.n65 171.744
R578 VDD1.n65 VDD1.n3 171.744
R579 VDD1.n58 VDD1.n3 171.744
R580 VDD1.n58 VDD1.n57 171.744
R581 VDD1.n57 VDD1.n7 171.744
R582 VDD1.n50 VDD1.n7 171.744
R583 VDD1.n50 VDD1.n49 171.744
R584 VDD1.n49 VDD1.n11 171.744
R585 VDD1.n42 VDD1.n11 171.744
R586 VDD1.n42 VDD1.n41 171.744
R587 VDD1.n41 VDD1.n15 171.744
R588 VDD1.n34 VDD1.n15 171.744
R589 VDD1.n34 VDD1.n33 171.744
R590 VDD1.n33 VDD1.n19 171.744
R591 VDD1.n26 VDD1.n19 171.744
R592 VDD1.n26 VDD1.n25 171.744
R593 VDD1.n99 VDD1.n98 171.744
R594 VDD1.n99 VDD1.n92 171.744
R595 VDD1.n106 VDD1.n92 171.744
R596 VDD1.n107 VDD1.n106 171.744
R597 VDD1.n107 VDD1.n88 171.744
R598 VDD1.n114 VDD1.n88 171.744
R599 VDD1.n115 VDD1.n114 171.744
R600 VDD1.n115 VDD1.n84 171.744
R601 VDD1.n122 VDD1.n84 171.744
R602 VDD1.n123 VDD1.n122 171.744
R603 VDD1.n123 VDD1.n80 171.744
R604 VDD1.n130 VDD1.n80 171.744
R605 VDD1.n131 VDD1.n130 171.744
R606 VDD1.n131 VDD1.n76 171.744
R607 VDD1.n138 VDD1.n76 171.744
R608 VDD1.n139 VDD1.n138 171.744
R609 VDD1.n25 VDD1.t9 85.8723
R610 VDD1.n98 VDD1.t6 85.8723
R611 VDD1.n147 VDD1.n146 77.238
R612 VDD1.n72 VDD1.n71 76.4272
R613 VDD1.n149 VDD1.n148 76.427
R614 VDD1.n145 VDD1.n144 76.427
R615 VDD1.n72 VDD1.n70 54.4799
R616 VDD1.n145 VDD1.n143 54.4799
R617 VDD1.n149 VDD1.n147 41.9405
R618 VDD1.n24 VDD1.n23 16.3895
R619 VDD1.n97 VDD1.n96 16.3895
R620 VDD1.n68 VDD1.n67 12.8005
R621 VDD1.n27 VDD1.n22 12.8005
R622 VDD1.n100 VDD1.n95 12.8005
R623 VDD1.n141 VDD1.n140 12.8005
R624 VDD1.n64 VDD1.n2 12.0247
R625 VDD1.n28 VDD1.n20 12.0247
R626 VDD1.n101 VDD1.n93 12.0247
R627 VDD1.n137 VDD1.n75 12.0247
R628 VDD1.n63 VDD1.n4 11.249
R629 VDD1.n32 VDD1.n31 11.249
R630 VDD1.n105 VDD1.n104 11.249
R631 VDD1.n136 VDD1.n77 11.249
R632 VDD1.n60 VDD1.n59 10.4732
R633 VDD1.n35 VDD1.n18 10.4732
R634 VDD1.n108 VDD1.n91 10.4732
R635 VDD1.n133 VDD1.n132 10.4732
R636 VDD1.n56 VDD1.n6 9.69747
R637 VDD1.n36 VDD1.n16 9.69747
R638 VDD1.n109 VDD1.n89 9.69747
R639 VDD1.n129 VDD1.n79 9.69747
R640 VDD1.n70 VDD1.n69 9.45567
R641 VDD1.n143 VDD1.n142 9.45567
R642 VDD1.n10 VDD1.n9 9.3005
R643 VDD1.n53 VDD1.n52 9.3005
R644 VDD1.n55 VDD1.n54 9.3005
R645 VDD1.n6 VDD1.n5 9.3005
R646 VDD1.n61 VDD1.n60 9.3005
R647 VDD1.n63 VDD1.n62 9.3005
R648 VDD1.n2 VDD1.n1 9.3005
R649 VDD1.n69 VDD1.n68 9.3005
R650 VDD1.n47 VDD1.n46 9.3005
R651 VDD1.n45 VDD1.n44 9.3005
R652 VDD1.n14 VDD1.n13 9.3005
R653 VDD1.n39 VDD1.n38 9.3005
R654 VDD1.n37 VDD1.n36 9.3005
R655 VDD1.n18 VDD1.n17 9.3005
R656 VDD1.n31 VDD1.n30 9.3005
R657 VDD1.n29 VDD1.n28 9.3005
R658 VDD1.n22 VDD1.n21 9.3005
R659 VDD1.n118 VDD1.n117 9.3005
R660 VDD1.n87 VDD1.n86 9.3005
R661 VDD1.n112 VDD1.n111 9.3005
R662 VDD1.n110 VDD1.n109 9.3005
R663 VDD1.n91 VDD1.n90 9.3005
R664 VDD1.n104 VDD1.n103 9.3005
R665 VDD1.n102 VDD1.n101 9.3005
R666 VDD1.n95 VDD1.n94 9.3005
R667 VDD1.n120 VDD1.n119 9.3005
R668 VDD1.n83 VDD1.n82 9.3005
R669 VDD1.n126 VDD1.n125 9.3005
R670 VDD1.n128 VDD1.n127 9.3005
R671 VDD1.n79 VDD1.n78 9.3005
R672 VDD1.n134 VDD1.n133 9.3005
R673 VDD1.n136 VDD1.n135 9.3005
R674 VDD1.n75 VDD1.n74 9.3005
R675 VDD1.n142 VDD1.n141 9.3005
R676 VDD1.n55 VDD1.n8 8.92171
R677 VDD1.n40 VDD1.n39 8.92171
R678 VDD1.n113 VDD1.n112 8.92171
R679 VDD1.n128 VDD1.n81 8.92171
R680 VDD1.n52 VDD1.n51 8.14595
R681 VDD1.n43 VDD1.n14 8.14595
R682 VDD1.n116 VDD1.n87 8.14595
R683 VDD1.n125 VDD1.n124 8.14595
R684 VDD1.n70 VDD1.n0 7.75445
R685 VDD1.n143 VDD1.n73 7.75445
R686 VDD1.n48 VDD1.n10 7.3702
R687 VDD1.n44 VDD1.n12 7.3702
R688 VDD1.n117 VDD1.n85 7.3702
R689 VDD1.n121 VDD1.n83 7.3702
R690 VDD1.n48 VDD1.n47 6.59444
R691 VDD1.n47 VDD1.n12 6.59444
R692 VDD1.n120 VDD1.n85 6.59444
R693 VDD1.n121 VDD1.n120 6.59444
R694 VDD1.n68 VDD1.n0 6.08283
R695 VDD1.n141 VDD1.n73 6.08283
R696 VDD1.n51 VDD1.n10 5.81868
R697 VDD1.n44 VDD1.n43 5.81868
R698 VDD1.n117 VDD1.n116 5.81868
R699 VDD1.n124 VDD1.n83 5.81868
R700 VDD1.n52 VDD1.n8 5.04292
R701 VDD1.n40 VDD1.n14 5.04292
R702 VDD1.n113 VDD1.n87 5.04292
R703 VDD1.n125 VDD1.n81 5.04292
R704 VDD1.n56 VDD1.n55 4.26717
R705 VDD1.n39 VDD1.n16 4.26717
R706 VDD1.n112 VDD1.n89 4.26717
R707 VDD1.n129 VDD1.n128 4.26717
R708 VDD1.n23 VDD1.n21 3.70982
R709 VDD1.n96 VDD1.n94 3.70982
R710 VDD1.n59 VDD1.n6 3.49141
R711 VDD1.n36 VDD1.n35 3.49141
R712 VDD1.n109 VDD1.n108 3.49141
R713 VDD1.n132 VDD1.n79 3.49141
R714 VDD1.n60 VDD1.n4 2.71565
R715 VDD1.n32 VDD1.n18 2.71565
R716 VDD1.n105 VDD1.n91 2.71565
R717 VDD1.n133 VDD1.n77 2.71565
R718 VDD1.n148 VDD1.t8 2.42083
R719 VDD1.n148 VDD1.t2 2.42083
R720 VDD1.n71 VDD1.t7 2.42083
R721 VDD1.n71 VDD1.t0 2.42083
R722 VDD1.n146 VDD1.t3 2.42083
R723 VDD1.n146 VDD1.t5 2.42083
R724 VDD1.n144 VDD1.t1 2.42083
R725 VDD1.n144 VDD1.t4 2.42083
R726 VDD1.n64 VDD1.n63 1.93989
R727 VDD1.n31 VDD1.n20 1.93989
R728 VDD1.n104 VDD1.n93 1.93989
R729 VDD1.n137 VDD1.n136 1.93989
R730 VDD1.n67 VDD1.n2 1.16414
R731 VDD1.n28 VDD1.n27 1.16414
R732 VDD1.n101 VDD1.n100 1.16414
R733 VDD1.n140 VDD1.n75 1.16414
R734 VDD1 VDD1.n149 0.80869
R735 VDD1.n24 VDD1.n22 0.388379
R736 VDD1.n97 VDD1.n95 0.388379
R737 VDD1 VDD1.n72 0.347483
R738 VDD1.n147 VDD1.n145 0.233947
R739 VDD1.n69 VDD1.n1 0.155672
R740 VDD1.n62 VDD1.n1 0.155672
R741 VDD1.n62 VDD1.n61 0.155672
R742 VDD1.n61 VDD1.n5 0.155672
R743 VDD1.n54 VDD1.n5 0.155672
R744 VDD1.n54 VDD1.n53 0.155672
R745 VDD1.n53 VDD1.n9 0.155672
R746 VDD1.n46 VDD1.n9 0.155672
R747 VDD1.n46 VDD1.n45 0.155672
R748 VDD1.n45 VDD1.n13 0.155672
R749 VDD1.n38 VDD1.n13 0.155672
R750 VDD1.n38 VDD1.n37 0.155672
R751 VDD1.n37 VDD1.n17 0.155672
R752 VDD1.n30 VDD1.n17 0.155672
R753 VDD1.n30 VDD1.n29 0.155672
R754 VDD1.n29 VDD1.n21 0.155672
R755 VDD1.n102 VDD1.n94 0.155672
R756 VDD1.n103 VDD1.n102 0.155672
R757 VDD1.n103 VDD1.n90 0.155672
R758 VDD1.n110 VDD1.n90 0.155672
R759 VDD1.n111 VDD1.n110 0.155672
R760 VDD1.n111 VDD1.n86 0.155672
R761 VDD1.n118 VDD1.n86 0.155672
R762 VDD1.n119 VDD1.n118 0.155672
R763 VDD1.n119 VDD1.n82 0.155672
R764 VDD1.n126 VDD1.n82 0.155672
R765 VDD1.n127 VDD1.n126 0.155672
R766 VDD1.n127 VDD1.n78 0.155672
R767 VDD1.n134 VDD1.n78 0.155672
R768 VDD1.n135 VDD1.n134 0.155672
R769 VDD1.n135 VDD1.n74 0.155672
R770 VDD1.n142 VDD1.n74 0.155672
R771 VN.n5 VN.t2 374.082
R772 VN.n25 VN.t7 374.082
R773 VN.n18 VN.t6 359.591
R774 VN.n38 VN.t5 359.591
R775 VN.n4 VN.t4 320.459
R776 VN.n10 VN.t1 320.459
R777 VN.n16 VN.t3 320.459
R778 VN.n24 VN.t9 320.459
R779 VN.n30 VN.t0 320.459
R780 VN.n36 VN.t8 320.459
R781 VN.n37 VN.n20 161.3
R782 VN.n35 VN.n34 161.3
R783 VN.n33 VN.n21 161.3
R784 VN.n32 VN.n31 161.3
R785 VN.n29 VN.n22 161.3
R786 VN.n28 VN.n27 161.3
R787 VN.n26 VN.n23 161.3
R788 VN.n17 VN.n0 161.3
R789 VN.n15 VN.n14 161.3
R790 VN.n13 VN.n1 161.3
R791 VN.n12 VN.n11 161.3
R792 VN.n9 VN.n2 161.3
R793 VN.n8 VN.n7 161.3
R794 VN.n6 VN.n3 161.3
R795 VN.n39 VN.n38 80.6037
R796 VN.n19 VN.n18 80.6037
R797 VN.n18 VN.n17 52.8492
R798 VN.n38 VN.n37 52.8492
R799 VN.n5 VN.n4 48.957
R800 VN.n25 VN.n24 48.957
R801 VN.n9 VN.n8 48.2635
R802 VN.n11 VN.n1 48.2635
R803 VN.n29 VN.n28 48.2635
R804 VN.n31 VN.n21 48.2635
R805 VN VN.n39 46.0066
R806 VN.n26 VN.n25 44.4127
R807 VN.n6 VN.n5 44.4127
R808 VN.n8 VN.n3 32.7233
R809 VN.n15 VN.n1 32.7233
R810 VN.n28 VN.n23 32.7233
R811 VN.n35 VN.n21 32.7233
R812 VN.n17 VN.n16 20.0634
R813 VN.n37 VN.n36 20.0634
R814 VN.n10 VN.n9 12.234
R815 VN.n11 VN.n10 12.234
R816 VN.n31 VN.n30 12.234
R817 VN.n30 VN.n29 12.234
R818 VN.n4 VN.n3 4.40456
R819 VN.n16 VN.n15 4.40456
R820 VN.n24 VN.n23 4.40456
R821 VN.n36 VN.n35 4.40456
R822 VN.n39 VN.n20 0.285035
R823 VN.n19 VN.n0 0.285035
R824 VN.n34 VN.n20 0.189894
R825 VN.n34 VN.n33 0.189894
R826 VN.n33 VN.n32 0.189894
R827 VN.n32 VN.n22 0.189894
R828 VN.n27 VN.n22 0.189894
R829 VN.n27 VN.n26 0.189894
R830 VN.n7 VN.n6 0.189894
R831 VN.n7 VN.n2 0.189894
R832 VN.n12 VN.n2 0.189894
R833 VN.n13 VN.n12 0.189894
R834 VN.n14 VN.n13 0.189894
R835 VN.n14 VN.n0 0.189894
R836 VN VN.n19 0.146778
R837 VDD2.n142 VDD2.n141 585
R838 VDD2.n140 VDD2.n139 585
R839 VDD2.n79 VDD2.n78 585
R840 VDD2.n134 VDD2.n133 585
R841 VDD2.n132 VDD2.n131 585
R842 VDD2.n83 VDD2.n82 585
R843 VDD2.n126 VDD2.n125 585
R844 VDD2.n124 VDD2.n123 585
R845 VDD2.n87 VDD2.n86 585
R846 VDD2.n118 VDD2.n117 585
R847 VDD2.n116 VDD2.n115 585
R848 VDD2.n91 VDD2.n90 585
R849 VDD2.n110 VDD2.n109 585
R850 VDD2.n108 VDD2.n107 585
R851 VDD2.n95 VDD2.n94 585
R852 VDD2.n102 VDD2.n101 585
R853 VDD2.n100 VDD2.n99 585
R854 VDD2.n25 VDD2.n24 585
R855 VDD2.n27 VDD2.n26 585
R856 VDD2.n20 VDD2.n19 585
R857 VDD2.n33 VDD2.n32 585
R858 VDD2.n35 VDD2.n34 585
R859 VDD2.n16 VDD2.n15 585
R860 VDD2.n41 VDD2.n40 585
R861 VDD2.n43 VDD2.n42 585
R862 VDD2.n12 VDD2.n11 585
R863 VDD2.n49 VDD2.n48 585
R864 VDD2.n51 VDD2.n50 585
R865 VDD2.n8 VDD2.n7 585
R866 VDD2.n57 VDD2.n56 585
R867 VDD2.n59 VDD2.n58 585
R868 VDD2.n4 VDD2.n3 585
R869 VDD2.n65 VDD2.n64 585
R870 VDD2.n67 VDD2.n66 585
R871 VDD2.n141 VDD2.n75 498.474
R872 VDD2.n66 VDD2.n0 498.474
R873 VDD2.n98 VDD2.t4 327.466
R874 VDD2.n23 VDD2.t7 327.466
R875 VDD2.n141 VDD2.n140 171.744
R876 VDD2.n140 VDD2.n78 171.744
R877 VDD2.n133 VDD2.n78 171.744
R878 VDD2.n133 VDD2.n132 171.744
R879 VDD2.n132 VDD2.n82 171.744
R880 VDD2.n125 VDD2.n82 171.744
R881 VDD2.n125 VDD2.n124 171.744
R882 VDD2.n124 VDD2.n86 171.744
R883 VDD2.n117 VDD2.n86 171.744
R884 VDD2.n117 VDD2.n116 171.744
R885 VDD2.n116 VDD2.n90 171.744
R886 VDD2.n109 VDD2.n90 171.744
R887 VDD2.n109 VDD2.n108 171.744
R888 VDD2.n108 VDD2.n94 171.744
R889 VDD2.n101 VDD2.n94 171.744
R890 VDD2.n101 VDD2.n100 171.744
R891 VDD2.n26 VDD2.n25 171.744
R892 VDD2.n26 VDD2.n19 171.744
R893 VDD2.n33 VDD2.n19 171.744
R894 VDD2.n34 VDD2.n33 171.744
R895 VDD2.n34 VDD2.n15 171.744
R896 VDD2.n41 VDD2.n15 171.744
R897 VDD2.n42 VDD2.n41 171.744
R898 VDD2.n42 VDD2.n11 171.744
R899 VDD2.n49 VDD2.n11 171.744
R900 VDD2.n50 VDD2.n49 171.744
R901 VDD2.n50 VDD2.n7 171.744
R902 VDD2.n57 VDD2.n7 171.744
R903 VDD2.n58 VDD2.n57 171.744
R904 VDD2.n58 VDD2.n3 171.744
R905 VDD2.n65 VDD2.n3 171.744
R906 VDD2.n66 VDD2.n65 171.744
R907 VDD2.n100 VDD2.t4 85.8723
R908 VDD2.n25 VDD2.t7 85.8723
R909 VDD2.n74 VDD2.n73 77.238
R910 VDD2 VDD2.n149 77.2352
R911 VDD2.n148 VDD2.n147 76.4272
R912 VDD2.n72 VDD2.n71 76.427
R913 VDD2.n72 VDD2.n70 54.4799
R914 VDD2.n146 VDD2.n145 53.3247
R915 VDD2.n146 VDD2.n74 40.7799
R916 VDD2.n99 VDD2.n98 16.3895
R917 VDD2.n24 VDD2.n23 16.3895
R918 VDD2.n143 VDD2.n142 12.8005
R919 VDD2.n102 VDD2.n97 12.8005
R920 VDD2.n27 VDD2.n22 12.8005
R921 VDD2.n68 VDD2.n67 12.8005
R922 VDD2.n139 VDD2.n77 12.0247
R923 VDD2.n103 VDD2.n95 12.0247
R924 VDD2.n28 VDD2.n20 12.0247
R925 VDD2.n64 VDD2.n2 12.0247
R926 VDD2.n138 VDD2.n79 11.249
R927 VDD2.n107 VDD2.n106 11.249
R928 VDD2.n32 VDD2.n31 11.249
R929 VDD2.n63 VDD2.n4 11.249
R930 VDD2.n135 VDD2.n134 10.4732
R931 VDD2.n110 VDD2.n93 10.4732
R932 VDD2.n35 VDD2.n18 10.4732
R933 VDD2.n60 VDD2.n59 10.4732
R934 VDD2.n131 VDD2.n81 9.69747
R935 VDD2.n111 VDD2.n91 9.69747
R936 VDD2.n36 VDD2.n16 9.69747
R937 VDD2.n56 VDD2.n6 9.69747
R938 VDD2.n145 VDD2.n144 9.45567
R939 VDD2.n70 VDD2.n69 9.45567
R940 VDD2.n85 VDD2.n84 9.3005
R941 VDD2.n128 VDD2.n127 9.3005
R942 VDD2.n130 VDD2.n129 9.3005
R943 VDD2.n81 VDD2.n80 9.3005
R944 VDD2.n136 VDD2.n135 9.3005
R945 VDD2.n138 VDD2.n137 9.3005
R946 VDD2.n77 VDD2.n76 9.3005
R947 VDD2.n144 VDD2.n143 9.3005
R948 VDD2.n122 VDD2.n121 9.3005
R949 VDD2.n120 VDD2.n119 9.3005
R950 VDD2.n89 VDD2.n88 9.3005
R951 VDD2.n114 VDD2.n113 9.3005
R952 VDD2.n112 VDD2.n111 9.3005
R953 VDD2.n93 VDD2.n92 9.3005
R954 VDD2.n106 VDD2.n105 9.3005
R955 VDD2.n104 VDD2.n103 9.3005
R956 VDD2.n97 VDD2.n96 9.3005
R957 VDD2.n45 VDD2.n44 9.3005
R958 VDD2.n14 VDD2.n13 9.3005
R959 VDD2.n39 VDD2.n38 9.3005
R960 VDD2.n37 VDD2.n36 9.3005
R961 VDD2.n18 VDD2.n17 9.3005
R962 VDD2.n31 VDD2.n30 9.3005
R963 VDD2.n29 VDD2.n28 9.3005
R964 VDD2.n22 VDD2.n21 9.3005
R965 VDD2.n47 VDD2.n46 9.3005
R966 VDD2.n10 VDD2.n9 9.3005
R967 VDD2.n53 VDD2.n52 9.3005
R968 VDD2.n55 VDD2.n54 9.3005
R969 VDD2.n6 VDD2.n5 9.3005
R970 VDD2.n61 VDD2.n60 9.3005
R971 VDD2.n63 VDD2.n62 9.3005
R972 VDD2.n2 VDD2.n1 9.3005
R973 VDD2.n69 VDD2.n68 9.3005
R974 VDD2.n130 VDD2.n83 8.92171
R975 VDD2.n115 VDD2.n114 8.92171
R976 VDD2.n40 VDD2.n39 8.92171
R977 VDD2.n55 VDD2.n8 8.92171
R978 VDD2.n127 VDD2.n126 8.14595
R979 VDD2.n118 VDD2.n89 8.14595
R980 VDD2.n43 VDD2.n14 8.14595
R981 VDD2.n52 VDD2.n51 8.14595
R982 VDD2.n145 VDD2.n75 7.75445
R983 VDD2.n70 VDD2.n0 7.75445
R984 VDD2.n123 VDD2.n85 7.3702
R985 VDD2.n119 VDD2.n87 7.3702
R986 VDD2.n44 VDD2.n12 7.3702
R987 VDD2.n48 VDD2.n10 7.3702
R988 VDD2.n123 VDD2.n122 6.59444
R989 VDD2.n122 VDD2.n87 6.59444
R990 VDD2.n47 VDD2.n12 6.59444
R991 VDD2.n48 VDD2.n47 6.59444
R992 VDD2.n143 VDD2.n75 6.08283
R993 VDD2.n68 VDD2.n0 6.08283
R994 VDD2.n126 VDD2.n85 5.81868
R995 VDD2.n119 VDD2.n118 5.81868
R996 VDD2.n44 VDD2.n43 5.81868
R997 VDD2.n51 VDD2.n10 5.81868
R998 VDD2.n127 VDD2.n83 5.04292
R999 VDD2.n115 VDD2.n89 5.04292
R1000 VDD2.n40 VDD2.n14 5.04292
R1001 VDD2.n52 VDD2.n8 5.04292
R1002 VDD2.n131 VDD2.n130 4.26717
R1003 VDD2.n114 VDD2.n91 4.26717
R1004 VDD2.n39 VDD2.n16 4.26717
R1005 VDD2.n56 VDD2.n55 4.26717
R1006 VDD2.n98 VDD2.n96 3.70982
R1007 VDD2.n23 VDD2.n21 3.70982
R1008 VDD2.n134 VDD2.n81 3.49141
R1009 VDD2.n111 VDD2.n110 3.49141
R1010 VDD2.n36 VDD2.n35 3.49141
R1011 VDD2.n59 VDD2.n6 3.49141
R1012 VDD2.n135 VDD2.n79 2.71565
R1013 VDD2.n107 VDD2.n93 2.71565
R1014 VDD2.n32 VDD2.n18 2.71565
R1015 VDD2.n60 VDD2.n4 2.71565
R1016 VDD2.n149 VDD2.t0 2.42083
R1017 VDD2.n149 VDD2.t2 2.42083
R1018 VDD2.n147 VDD2.t1 2.42083
R1019 VDD2.n147 VDD2.t9 2.42083
R1020 VDD2.n73 VDD2.t6 2.42083
R1021 VDD2.n73 VDD2.t3 2.42083
R1022 VDD2.n71 VDD2.t5 2.42083
R1023 VDD2.n71 VDD2.t8 2.42083
R1024 VDD2.n139 VDD2.n138 1.93989
R1025 VDD2.n106 VDD2.n95 1.93989
R1026 VDD2.n31 VDD2.n20 1.93989
R1027 VDD2.n64 VDD2.n63 1.93989
R1028 VDD2.n142 VDD2.n77 1.16414
R1029 VDD2.n103 VDD2.n102 1.16414
R1030 VDD2.n28 VDD2.n27 1.16414
R1031 VDD2.n67 VDD2.n2 1.16414
R1032 VDD2.n148 VDD2.n146 1.15567
R1033 VDD2.n99 VDD2.n97 0.388379
R1034 VDD2.n24 VDD2.n22 0.388379
R1035 VDD2 VDD2.n148 0.347483
R1036 VDD2.n74 VDD2.n72 0.233947
R1037 VDD2.n144 VDD2.n76 0.155672
R1038 VDD2.n137 VDD2.n76 0.155672
R1039 VDD2.n137 VDD2.n136 0.155672
R1040 VDD2.n136 VDD2.n80 0.155672
R1041 VDD2.n129 VDD2.n80 0.155672
R1042 VDD2.n129 VDD2.n128 0.155672
R1043 VDD2.n128 VDD2.n84 0.155672
R1044 VDD2.n121 VDD2.n84 0.155672
R1045 VDD2.n121 VDD2.n120 0.155672
R1046 VDD2.n120 VDD2.n88 0.155672
R1047 VDD2.n113 VDD2.n88 0.155672
R1048 VDD2.n113 VDD2.n112 0.155672
R1049 VDD2.n112 VDD2.n92 0.155672
R1050 VDD2.n105 VDD2.n92 0.155672
R1051 VDD2.n105 VDD2.n104 0.155672
R1052 VDD2.n104 VDD2.n96 0.155672
R1053 VDD2.n29 VDD2.n21 0.155672
R1054 VDD2.n30 VDD2.n29 0.155672
R1055 VDD2.n30 VDD2.n17 0.155672
R1056 VDD2.n37 VDD2.n17 0.155672
R1057 VDD2.n38 VDD2.n37 0.155672
R1058 VDD2.n38 VDD2.n13 0.155672
R1059 VDD2.n45 VDD2.n13 0.155672
R1060 VDD2.n46 VDD2.n45 0.155672
R1061 VDD2.n46 VDD2.n9 0.155672
R1062 VDD2.n53 VDD2.n9 0.155672
R1063 VDD2.n54 VDD2.n53 0.155672
R1064 VDD2.n54 VDD2.n5 0.155672
R1065 VDD2.n61 VDD2.n5 0.155672
R1066 VDD2.n62 VDD2.n61 0.155672
R1067 VDD2.n62 VDD2.n1 0.155672
R1068 VDD2.n69 VDD2.n1 0.155672
R1069 B.n372 B.n105 585
R1070 B.n371 B.n370 585
R1071 B.n369 B.n106 585
R1072 B.n368 B.n367 585
R1073 B.n366 B.n107 585
R1074 B.n365 B.n364 585
R1075 B.n363 B.n108 585
R1076 B.n362 B.n361 585
R1077 B.n360 B.n109 585
R1078 B.n359 B.n358 585
R1079 B.n357 B.n110 585
R1080 B.n356 B.n355 585
R1081 B.n354 B.n111 585
R1082 B.n353 B.n352 585
R1083 B.n351 B.n112 585
R1084 B.n350 B.n349 585
R1085 B.n348 B.n113 585
R1086 B.n347 B.n346 585
R1087 B.n345 B.n114 585
R1088 B.n344 B.n343 585
R1089 B.n342 B.n115 585
R1090 B.n341 B.n340 585
R1091 B.n339 B.n116 585
R1092 B.n338 B.n337 585
R1093 B.n336 B.n117 585
R1094 B.n335 B.n334 585
R1095 B.n333 B.n118 585
R1096 B.n332 B.n331 585
R1097 B.n330 B.n119 585
R1098 B.n329 B.n328 585
R1099 B.n327 B.n120 585
R1100 B.n326 B.n325 585
R1101 B.n324 B.n121 585
R1102 B.n323 B.n322 585
R1103 B.n321 B.n122 585
R1104 B.n320 B.n319 585
R1105 B.n318 B.n123 585
R1106 B.n317 B.n316 585
R1107 B.n315 B.n124 585
R1108 B.n314 B.n313 585
R1109 B.n312 B.n125 585
R1110 B.n311 B.n310 585
R1111 B.n309 B.n126 585
R1112 B.n308 B.n307 585
R1113 B.n306 B.n127 585
R1114 B.n305 B.n304 585
R1115 B.n302 B.n128 585
R1116 B.n301 B.n300 585
R1117 B.n299 B.n131 585
R1118 B.n298 B.n297 585
R1119 B.n296 B.n132 585
R1120 B.n295 B.n294 585
R1121 B.n293 B.n133 585
R1122 B.n292 B.n291 585
R1123 B.n290 B.n134 585
R1124 B.n288 B.n287 585
R1125 B.n286 B.n137 585
R1126 B.n285 B.n284 585
R1127 B.n283 B.n138 585
R1128 B.n282 B.n281 585
R1129 B.n280 B.n139 585
R1130 B.n279 B.n278 585
R1131 B.n277 B.n140 585
R1132 B.n276 B.n275 585
R1133 B.n274 B.n141 585
R1134 B.n273 B.n272 585
R1135 B.n271 B.n142 585
R1136 B.n270 B.n269 585
R1137 B.n268 B.n143 585
R1138 B.n267 B.n266 585
R1139 B.n265 B.n144 585
R1140 B.n264 B.n263 585
R1141 B.n262 B.n145 585
R1142 B.n261 B.n260 585
R1143 B.n259 B.n146 585
R1144 B.n258 B.n257 585
R1145 B.n256 B.n147 585
R1146 B.n255 B.n254 585
R1147 B.n253 B.n148 585
R1148 B.n252 B.n251 585
R1149 B.n250 B.n149 585
R1150 B.n249 B.n248 585
R1151 B.n247 B.n150 585
R1152 B.n246 B.n245 585
R1153 B.n244 B.n151 585
R1154 B.n243 B.n242 585
R1155 B.n241 B.n152 585
R1156 B.n240 B.n239 585
R1157 B.n238 B.n153 585
R1158 B.n237 B.n236 585
R1159 B.n235 B.n154 585
R1160 B.n234 B.n233 585
R1161 B.n232 B.n155 585
R1162 B.n231 B.n230 585
R1163 B.n229 B.n156 585
R1164 B.n228 B.n227 585
R1165 B.n226 B.n157 585
R1166 B.n225 B.n224 585
R1167 B.n223 B.n158 585
R1168 B.n222 B.n221 585
R1169 B.n220 B.n159 585
R1170 B.n374 B.n373 585
R1171 B.n375 B.n104 585
R1172 B.n377 B.n376 585
R1173 B.n378 B.n103 585
R1174 B.n380 B.n379 585
R1175 B.n381 B.n102 585
R1176 B.n383 B.n382 585
R1177 B.n384 B.n101 585
R1178 B.n386 B.n385 585
R1179 B.n387 B.n100 585
R1180 B.n389 B.n388 585
R1181 B.n390 B.n99 585
R1182 B.n392 B.n391 585
R1183 B.n393 B.n98 585
R1184 B.n395 B.n394 585
R1185 B.n396 B.n97 585
R1186 B.n398 B.n397 585
R1187 B.n399 B.n96 585
R1188 B.n401 B.n400 585
R1189 B.n402 B.n95 585
R1190 B.n404 B.n403 585
R1191 B.n405 B.n94 585
R1192 B.n407 B.n406 585
R1193 B.n408 B.n93 585
R1194 B.n410 B.n409 585
R1195 B.n411 B.n92 585
R1196 B.n413 B.n412 585
R1197 B.n414 B.n91 585
R1198 B.n416 B.n415 585
R1199 B.n417 B.n90 585
R1200 B.n419 B.n418 585
R1201 B.n420 B.n89 585
R1202 B.n422 B.n421 585
R1203 B.n423 B.n88 585
R1204 B.n425 B.n424 585
R1205 B.n426 B.n87 585
R1206 B.n428 B.n427 585
R1207 B.n429 B.n86 585
R1208 B.n431 B.n430 585
R1209 B.n432 B.n85 585
R1210 B.n434 B.n433 585
R1211 B.n435 B.n84 585
R1212 B.n437 B.n436 585
R1213 B.n438 B.n83 585
R1214 B.n440 B.n439 585
R1215 B.n441 B.n82 585
R1216 B.n443 B.n442 585
R1217 B.n444 B.n81 585
R1218 B.n446 B.n445 585
R1219 B.n447 B.n80 585
R1220 B.n449 B.n448 585
R1221 B.n450 B.n79 585
R1222 B.n452 B.n451 585
R1223 B.n453 B.n78 585
R1224 B.n455 B.n454 585
R1225 B.n456 B.n77 585
R1226 B.n458 B.n457 585
R1227 B.n459 B.n76 585
R1228 B.n461 B.n460 585
R1229 B.n462 B.n75 585
R1230 B.n464 B.n463 585
R1231 B.n465 B.n74 585
R1232 B.n467 B.n466 585
R1233 B.n468 B.n73 585
R1234 B.n621 B.n620 585
R1235 B.n619 B.n18 585
R1236 B.n618 B.n617 585
R1237 B.n616 B.n19 585
R1238 B.n615 B.n614 585
R1239 B.n613 B.n20 585
R1240 B.n612 B.n611 585
R1241 B.n610 B.n21 585
R1242 B.n609 B.n608 585
R1243 B.n607 B.n22 585
R1244 B.n606 B.n605 585
R1245 B.n604 B.n23 585
R1246 B.n603 B.n602 585
R1247 B.n601 B.n24 585
R1248 B.n600 B.n599 585
R1249 B.n598 B.n25 585
R1250 B.n597 B.n596 585
R1251 B.n595 B.n26 585
R1252 B.n594 B.n593 585
R1253 B.n592 B.n27 585
R1254 B.n591 B.n590 585
R1255 B.n589 B.n28 585
R1256 B.n588 B.n587 585
R1257 B.n586 B.n29 585
R1258 B.n585 B.n584 585
R1259 B.n583 B.n30 585
R1260 B.n582 B.n581 585
R1261 B.n580 B.n31 585
R1262 B.n579 B.n578 585
R1263 B.n577 B.n32 585
R1264 B.n576 B.n575 585
R1265 B.n574 B.n33 585
R1266 B.n573 B.n572 585
R1267 B.n571 B.n34 585
R1268 B.n570 B.n569 585
R1269 B.n568 B.n35 585
R1270 B.n567 B.n566 585
R1271 B.n565 B.n36 585
R1272 B.n564 B.n563 585
R1273 B.n562 B.n37 585
R1274 B.n561 B.n560 585
R1275 B.n559 B.n38 585
R1276 B.n558 B.n557 585
R1277 B.n556 B.n39 585
R1278 B.n555 B.n554 585
R1279 B.n553 B.n40 585
R1280 B.n552 B.n551 585
R1281 B.n550 B.n41 585
R1282 B.n549 B.n548 585
R1283 B.n547 B.n45 585
R1284 B.n546 B.n545 585
R1285 B.n544 B.n46 585
R1286 B.n543 B.n542 585
R1287 B.n541 B.n47 585
R1288 B.n540 B.n539 585
R1289 B.n537 B.n48 585
R1290 B.n536 B.n535 585
R1291 B.n534 B.n51 585
R1292 B.n533 B.n532 585
R1293 B.n531 B.n52 585
R1294 B.n530 B.n529 585
R1295 B.n528 B.n53 585
R1296 B.n527 B.n526 585
R1297 B.n525 B.n54 585
R1298 B.n524 B.n523 585
R1299 B.n522 B.n55 585
R1300 B.n521 B.n520 585
R1301 B.n519 B.n56 585
R1302 B.n518 B.n517 585
R1303 B.n516 B.n57 585
R1304 B.n515 B.n514 585
R1305 B.n513 B.n58 585
R1306 B.n512 B.n511 585
R1307 B.n510 B.n59 585
R1308 B.n509 B.n508 585
R1309 B.n507 B.n60 585
R1310 B.n506 B.n505 585
R1311 B.n504 B.n61 585
R1312 B.n503 B.n502 585
R1313 B.n501 B.n62 585
R1314 B.n500 B.n499 585
R1315 B.n498 B.n63 585
R1316 B.n497 B.n496 585
R1317 B.n495 B.n64 585
R1318 B.n494 B.n493 585
R1319 B.n492 B.n65 585
R1320 B.n491 B.n490 585
R1321 B.n489 B.n66 585
R1322 B.n488 B.n487 585
R1323 B.n486 B.n67 585
R1324 B.n485 B.n484 585
R1325 B.n483 B.n68 585
R1326 B.n482 B.n481 585
R1327 B.n480 B.n69 585
R1328 B.n479 B.n478 585
R1329 B.n477 B.n70 585
R1330 B.n476 B.n475 585
R1331 B.n474 B.n71 585
R1332 B.n473 B.n472 585
R1333 B.n471 B.n72 585
R1334 B.n470 B.n469 585
R1335 B.n622 B.n17 585
R1336 B.n624 B.n623 585
R1337 B.n625 B.n16 585
R1338 B.n627 B.n626 585
R1339 B.n628 B.n15 585
R1340 B.n630 B.n629 585
R1341 B.n631 B.n14 585
R1342 B.n633 B.n632 585
R1343 B.n634 B.n13 585
R1344 B.n636 B.n635 585
R1345 B.n637 B.n12 585
R1346 B.n639 B.n638 585
R1347 B.n640 B.n11 585
R1348 B.n642 B.n641 585
R1349 B.n643 B.n10 585
R1350 B.n645 B.n644 585
R1351 B.n646 B.n9 585
R1352 B.n648 B.n647 585
R1353 B.n649 B.n8 585
R1354 B.n651 B.n650 585
R1355 B.n652 B.n7 585
R1356 B.n654 B.n653 585
R1357 B.n655 B.n6 585
R1358 B.n657 B.n656 585
R1359 B.n658 B.n5 585
R1360 B.n660 B.n659 585
R1361 B.n661 B.n4 585
R1362 B.n663 B.n662 585
R1363 B.n664 B.n3 585
R1364 B.n666 B.n665 585
R1365 B.n667 B.n0 585
R1366 B.n2 B.n1 585
R1367 B.n175 B.n174 585
R1368 B.n177 B.n176 585
R1369 B.n178 B.n173 585
R1370 B.n180 B.n179 585
R1371 B.n181 B.n172 585
R1372 B.n183 B.n182 585
R1373 B.n184 B.n171 585
R1374 B.n186 B.n185 585
R1375 B.n187 B.n170 585
R1376 B.n189 B.n188 585
R1377 B.n190 B.n169 585
R1378 B.n192 B.n191 585
R1379 B.n193 B.n168 585
R1380 B.n195 B.n194 585
R1381 B.n196 B.n167 585
R1382 B.n198 B.n197 585
R1383 B.n199 B.n166 585
R1384 B.n201 B.n200 585
R1385 B.n202 B.n165 585
R1386 B.n204 B.n203 585
R1387 B.n205 B.n164 585
R1388 B.n207 B.n206 585
R1389 B.n208 B.n163 585
R1390 B.n210 B.n209 585
R1391 B.n211 B.n162 585
R1392 B.n213 B.n212 585
R1393 B.n214 B.n161 585
R1394 B.n216 B.n215 585
R1395 B.n217 B.n160 585
R1396 B.n219 B.n218 585
R1397 B.n220 B.n219 559.769
R1398 B.n373 B.n372 559.769
R1399 B.n469 B.n468 559.769
R1400 B.n620 B.n17 559.769
R1401 B.n135 B.t0 523.452
R1402 B.n129 B.t9 523.452
R1403 B.n49 B.t3 523.452
R1404 B.n42 B.t6 523.452
R1405 B.n129 B.t10 427.37
R1406 B.n49 B.t5 427.37
R1407 B.n135 B.t1 427.37
R1408 B.n42 B.t8 427.37
R1409 B.n130 B.t11 401.382
R1410 B.n50 B.t4 401.382
R1411 B.n136 B.t2 401.382
R1412 B.n43 B.t7 401.382
R1413 B.n669 B.n668 256.663
R1414 B.n668 B.n667 235.042
R1415 B.n668 B.n2 235.042
R1416 B.n221 B.n220 163.367
R1417 B.n221 B.n158 163.367
R1418 B.n225 B.n158 163.367
R1419 B.n226 B.n225 163.367
R1420 B.n227 B.n226 163.367
R1421 B.n227 B.n156 163.367
R1422 B.n231 B.n156 163.367
R1423 B.n232 B.n231 163.367
R1424 B.n233 B.n232 163.367
R1425 B.n233 B.n154 163.367
R1426 B.n237 B.n154 163.367
R1427 B.n238 B.n237 163.367
R1428 B.n239 B.n238 163.367
R1429 B.n239 B.n152 163.367
R1430 B.n243 B.n152 163.367
R1431 B.n244 B.n243 163.367
R1432 B.n245 B.n244 163.367
R1433 B.n245 B.n150 163.367
R1434 B.n249 B.n150 163.367
R1435 B.n250 B.n249 163.367
R1436 B.n251 B.n250 163.367
R1437 B.n251 B.n148 163.367
R1438 B.n255 B.n148 163.367
R1439 B.n256 B.n255 163.367
R1440 B.n257 B.n256 163.367
R1441 B.n257 B.n146 163.367
R1442 B.n261 B.n146 163.367
R1443 B.n262 B.n261 163.367
R1444 B.n263 B.n262 163.367
R1445 B.n263 B.n144 163.367
R1446 B.n267 B.n144 163.367
R1447 B.n268 B.n267 163.367
R1448 B.n269 B.n268 163.367
R1449 B.n269 B.n142 163.367
R1450 B.n273 B.n142 163.367
R1451 B.n274 B.n273 163.367
R1452 B.n275 B.n274 163.367
R1453 B.n275 B.n140 163.367
R1454 B.n279 B.n140 163.367
R1455 B.n280 B.n279 163.367
R1456 B.n281 B.n280 163.367
R1457 B.n281 B.n138 163.367
R1458 B.n285 B.n138 163.367
R1459 B.n286 B.n285 163.367
R1460 B.n287 B.n286 163.367
R1461 B.n287 B.n134 163.367
R1462 B.n292 B.n134 163.367
R1463 B.n293 B.n292 163.367
R1464 B.n294 B.n293 163.367
R1465 B.n294 B.n132 163.367
R1466 B.n298 B.n132 163.367
R1467 B.n299 B.n298 163.367
R1468 B.n300 B.n299 163.367
R1469 B.n300 B.n128 163.367
R1470 B.n305 B.n128 163.367
R1471 B.n306 B.n305 163.367
R1472 B.n307 B.n306 163.367
R1473 B.n307 B.n126 163.367
R1474 B.n311 B.n126 163.367
R1475 B.n312 B.n311 163.367
R1476 B.n313 B.n312 163.367
R1477 B.n313 B.n124 163.367
R1478 B.n317 B.n124 163.367
R1479 B.n318 B.n317 163.367
R1480 B.n319 B.n318 163.367
R1481 B.n319 B.n122 163.367
R1482 B.n323 B.n122 163.367
R1483 B.n324 B.n323 163.367
R1484 B.n325 B.n324 163.367
R1485 B.n325 B.n120 163.367
R1486 B.n329 B.n120 163.367
R1487 B.n330 B.n329 163.367
R1488 B.n331 B.n330 163.367
R1489 B.n331 B.n118 163.367
R1490 B.n335 B.n118 163.367
R1491 B.n336 B.n335 163.367
R1492 B.n337 B.n336 163.367
R1493 B.n337 B.n116 163.367
R1494 B.n341 B.n116 163.367
R1495 B.n342 B.n341 163.367
R1496 B.n343 B.n342 163.367
R1497 B.n343 B.n114 163.367
R1498 B.n347 B.n114 163.367
R1499 B.n348 B.n347 163.367
R1500 B.n349 B.n348 163.367
R1501 B.n349 B.n112 163.367
R1502 B.n353 B.n112 163.367
R1503 B.n354 B.n353 163.367
R1504 B.n355 B.n354 163.367
R1505 B.n355 B.n110 163.367
R1506 B.n359 B.n110 163.367
R1507 B.n360 B.n359 163.367
R1508 B.n361 B.n360 163.367
R1509 B.n361 B.n108 163.367
R1510 B.n365 B.n108 163.367
R1511 B.n366 B.n365 163.367
R1512 B.n367 B.n366 163.367
R1513 B.n367 B.n106 163.367
R1514 B.n371 B.n106 163.367
R1515 B.n372 B.n371 163.367
R1516 B.n468 B.n467 163.367
R1517 B.n467 B.n74 163.367
R1518 B.n463 B.n74 163.367
R1519 B.n463 B.n462 163.367
R1520 B.n462 B.n461 163.367
R1521 B.n461 B.n76 163.367
R1522 B.n457 B.n76 163.367
R1523 B.n457 B.n456 163.367
R1524 B.n456 B.n455 163.367
R1525 B.n455 B.n78 163.367
R1526 B.n451 B.n78 163.367
R1527 B.n451 B.n450 163.367
R1528 B.n450 B.n449 163.367
R1529 B.n449 B.n80 163.367
R1530 B.n445 B.n80 163.367
R1531 B.n445 B.n444 163.367
R1532 B.n444 B.n443 163.367
R1533 B.n443 B.n82 163.367
R1534 B.n439 B.n82 163.367
R1535 B.n439 B.n438 163.367
R1536 B.n438 B.n437 163.367
R1537 B.n437 B.n84 163.367
R1538 B.n433 B.n84 163.367
R1539 B.n433 B.n432 163.367
R1540 B.n432 B.n431 163.367
R1541 B.n431 B.n86 163.367
R1542 B.n427 B.n86 163.367
R1543 B.n427 B.n426 163.367
R1544 B.n426 B.n425 163.367
R1545 B.n425 B.n88 163.367
R1546 B.n421 B.n88 163.367
R1547 B.n421 B.n420 163.367
R1548 B.n420 B.n419 163.367
R1549 B.n419 B.n90 163.367
R1550 B.n415 B.n90 163.367
R1551 B.n415 B.n414 163.367
R1552 B.n414 B.n413 163.367
R1553 B.n413 B.n92 163.367
R1554 B.n409 B.n92 163.367
R1555 B.n409 B.n408 163.367
R1556 B.n408 B.n407 163.367
R1557 B.n407 B.n94 163.367
R1558 B.n403 B.n94 163.367
R1559 B.n403 B.n402 163.367
R1560 B.n402 B.n401 163.367
R1561 B.n401 B.n96 163.367
R1562 B.n397 B.n96 163.367
R1563 B.n397 B.n396 163.367
R1564 B.n396 B.n395 163.367
R1565 B.n395 B.n98 163.367
R1566 B.n391 B.n98 163.367
R1567 B.n391 B.n390 163.367
R1568 B.n390 B.n389 163.367
R1569 B.n389 B.n100 163.367
R1570 B.n385 B.n100 163.367
R1571 B.n385 B.n384 163.367
R1572 B.n384 B.n383 163.367
R1573 B.n383 B.n102 163.367
R1574 B.n379 B.n102 163.367
R1575 B.n379 B.n378 163.367
R1576 B.n378 B.n377 163.367
R1577 B.n377 B.n104 163.367
R1578 B.n373 B.n104 163.367
R1579 B.n620 B.n619 163.367
R1580 B.n619 B.n618 163.367
R1581 B.n618 B.n19 163.367
R1582 B.n614 B.n19 163.367
R1583 B.n614 B.n613 163.367
R1584 B.n613 B.n612 163.367
R1585 B.n612 B.n21 163.367
R1586 B.n608 B.n21 163.367
R1587 B.n608 B.n607 163.367
R1588 B.n607 B.n606 163.367
R1589 B.n606 B.n23 163.367
R1590 B.n602 B.n23 163.367
R1591 B.n602 B.n601 163.367
R1592 B.n601 B.n600 163.367
R1593 B.n600 B.n25 163.367
R1594 B.n596 B.n25 163.367
R1595 B.n596 B.n595 163.367
R1596 B.n595 B.n594 163.367
R1597 B.n594 B.n27 163.367
R1598 B.n590 B.n27 163.367
R1599 B.n590 B.n589 163.367
R1600 B.n589 B.n588 163.367
R1601 B.n588 B.n29 163.367
R1602 B.n584 B.n29 163.367
R1603 B.n584 B.n583 163.367
R1604 B.n583 B.n582 163.367
R1605 B.n582 B.n31 163.367
R1606 B.n578 B.n31 163.367
R1607 B.n578 B.n577 163.367
R1608 B.n577 B.n576 163.367
R1609 B.n576 B.n33 163.367
R1610 B.n572 B.n33 163.367
R1611 B.n572 B.n571 163.367
R1612 B.n571 B.n570 163.367
R1613 B.n570 B.n35 163.367
R1614 B.n566 B.n35 163.367
R1615 B.n566 B.n565 163.367
R1616 B.n565 B.n564 163.367
R1617 B.n564 B.n37 163.367
R1618 B.n560 B.n37 163.367
R1619 B.n560 B.n559 163.367
R1620 B.n559 B.n558 163.367
R1621 B.n558 B.n39 163.367
R1622 B.n554 B.n39 163.367
R1623 B.n554 B.n553 163.367
R1624 B.n553 B.n552 163.367
R1625 B.n552 B.n41 163.367
R1626 B.n548 B.n41 163.367
R1627 B.n548 B.n547 163.367
R1628 B.n547 B.n546 163.367
R1629 B.n546 B.n46 163.367
R1630 B.n542 B.n46 163.367
R1631 B.n542 B.n541 163.367
R1632 B.n541 B.n540 163.367
R1633 B.n540 B.n48 163.367
R1634 B.n535 B.n48 163.367
R1635 B.n535 B.n534 163.367
R1636 B.n534 B.n533 163.367
R1637 B.n533 B.n52 163.367
R1638 B.n529 B.n52 163.367
R1639 B.n529 B.n528 163.367
R1640 B.n528 B.n527 163.367
R1641 B.n527 B.n54 163.367
R1642 B.n523 B.n54 163.367
R1643 B.n523 B.n522 163.367
R1644 B.n522 B.n521 163.367
R1645 B.n521 B.n56 163.367
R1646 B.n517 B.n56 163.367
R1647 B.n517 B.n516 163.367
R1648 B.n516 B.n515 163.367
R1649 B.n515 B.n58 163.367
R1650 B.n511 B.n58 163.367
R1651 B.n511 B.n510 163.367
R1652 B.n510 B.n509 163.367
R1653 B.n509 B.n60 163.367
R1654 B.n505 B.n60 163.367
R1655 B.n505 B.n504 163.367
R1656 B.n504 B.n503 163.367
R1657 B.n503 B.n62 163.367
R1658 B.n499 B.n62 163.367
R1659 B.n499 B.n498 163.367
R1660 B.n498 B.n497 163.367
R1661 B.n497 B.n64 163.367
R1662 B.n493 B.n64 163.367
R1663 B.n493 B.n492 163.367
R1664 B.n492 B.n491 163.367
R1665 B.n491 B.n66 163.367
R1666 B.n487 B.n66 163.367
R1667 B.n487 B.n486 163.367
R1668 B.n486 B.n485 163.367
R1669 B.n485 B.n68 163.367
R1670 B.n481 B.n68 163.367
R1671 B.n481 B.n480 163.367
R1672 B.n480 B.n479 163.367
R1673 B.n479 B.n70 163.367
R1674 B.n475 B.n70 163.367
R1675 B.n475 B.n474 163.367
R1676 B.n474 B.n473 163.367
R1677 B.n473 B.n72 163.367
R1678 B.n469 B.n72 163.367
R1679 B.n624 B.n17 163.367
R1680 B.n625 B.n624 163.367
R1681 B.n626 B.n625 163.367
R1682 B.n626 B.n15 163.367
R1683 B.n630 B.n15 163.367
R1684 B.n631 B.n630 163.367
R1685 B.n632 B.n631 163.367
R1686 B.n632 B.n13 163.367
R1687 B.n636 B.n13 163.367
R1688 B.n637 B.n636 163.367
R1689 B.n638 B.n637 163.367
R1690 B.n638 B.n11 163.367
R1691 B.n642 B.n11 163.367
R1692 B.n643 B.n642 163.367
R1693 B.n644 B.n643 163.367
R1694 B.n644 B.n9 163.367
R1695 B.n648 B.n9 163.367
R1696 B.n649 B.n648 163.367
R1697 B.n650 B.n649 163.367
R1698 B.n650 B.n7 163.367
R1699 B.n654 B.n7 163.367
R1700 B.n655 B.n654 163.367
R1701 B.n656 B.n655 163.367
R1702 B.n656 B.n5 163.367
R1703 B.n660 B.n5 163.367
R1704 B.n661 B.n660 163.367
R1705 B.n662 B.n661 163.367
R1706 B.n662 B.n3 163.367
R1707 B.n666 B.n3 163.367
R1708 B.n667 B.n666 163.367
R1709 B.n174 B.n2 163.367
R1710 B.n177 B.n174 163.367
R1711 B.n178 B.n177 163.367
R1712 B.n179 B.n178 163.367
R1713 B.n179 B.n172 163.367
R1714 B.n183 B.n172 163.367
R1715 B.n184 B.n183 163.367
R1716 B.n185 B.n184 163.367
R1717 B.n185 B.n170 163.367
R1718 B.n189 B.n170 163.367
R1719 B.n190 B.n189 163.367
R1720 B.n191 B.n190 163.367
R1721 B.n191 B.n168 163.367
R1722 B.n195 B.n168 163.367
R1723 B.n196 B.n195 163.367
R1724 B.n197 B.n196 163.367
R1725 B.n197 B.n166 163.367
R1726 B.n201 B.n166 163.367
R1727 B.n202 B.n201 163.367
R1728 B.n203 B.n202 163.367
R1729 B.n203 B.n164 163.367
R1730 B.n207 B.n164 163.367
R1731 B.n208 B.n207 163.367
R1732 B.n209 B.n208 163.367
R1733 B.n209 B.n162 163.367
R1734 B.n213 B.n162 163.367
R1735 B.n214 B.n213 163.367
R1736 B.n215 B.n214 163.367
R1737 B.n215 B.n160 163.367
R1738 B.n219 B.n160 163.367
R1739 B.n289 B.n136 59.5399
R1740 B.n303 B.n130 59.5399
R1741 B.n538 B.n50 59.5399
R1742 B.n44 B.n43 59.5399
R1743 B.n374 B.n105 36.3712
R1744 B.n622 B.n621 36.3712
R1745 B.n470 B.n73 36.3712
R1746 B.n218 B.n159 36.3712
R1747 B.n136 B.n135 25.9884
R1748 B.n130 B.n129 25.9884
R1749 B.n50 B.n49 25.9884
R1750 B.n43 B.n42 25.9884
R1751 B B.n669 18.0485
R1752 B.n623 B.n622 10.6151
R1753 B.n623 B.n16 10.6151
R1754 B.n627 B.n16 10.6151
R1755 B.n628 B.n627 10.6151
R1756 B.n629 B.n628 10.6151
R1757 B.n629 B.n14 10.6151
R1758 B.n633 B.n14 10.6151
R1759 B.n634 B.n633 10.6151
R1760 B.n635 B.n634 10.6151
R1761 B.n635 B.n12 10.6151
R1762 B.n639 B.n12 10.6151
R1763 B.n640 B.n639 10.6151
R1764 B.n641 B.n640 10.6151
R1765 B.n641 B.n10 10.6151
R1766 B.n645 B.n10 10.6151
R1767 B.n646 B.n645 10.6151
R1768 B.n647 B.n646 10.6151
R1769 B.n647 B.n8 10.6151
R1770 B.n651 B.n8 10.6151
R1771 B.n652 B.n651 10.6151
R1772 B.n653 B.n652 10.6151
R1773 B.n653 B.n6 10.6151
R1774 B.n657 B.n6 10.6151
R1775 B.n658 B.n657 10.6151
R1776 B.n659 B.n658 10.6151
R1777 B.n659 B.n4 10.6151
R1778 B.n663 B.n4 10.6151
R1779 B.n664 B.n663 10.6151
R1780 B.n665 B.n664 10.6151
R1781 B.n665 B.n0 10.6151
R1782 B.n621 B.n18 10.6151
R1783 B.n617 B.n18 10.6151
R1784 B.n617 B.n616 10.6151
R1785 B.n616 B.n615 10.6151
R1786 B.n615 B.n20 10.6151
R1787 B.n611 B.n20 10.6151
R1788 B.n611 B.n610 10.6151
R1789 B.n610 B.n609 10.6151
R1790 B.n609 B.n22 10.6151
R1791 B.n605 B.n22 10.6151
R1792 B.n605 B.n604 10.6151
R1793 B.n604 B.n603 10.6151
R1794 B.n603 B.n24 10.6151
R1795 B.n599 B.n24 10.6151
R1796 B.n599 B.n598 10.6151
R1797 B.n598 B.n597 10.6151
R1798 B.n597 B.n26 10.6151
R1799 B.n593 B.n26 10.6151
R1800 B.n593 B.n592 10.6151
R1801 B.n592 B.n591 10.6151
R1802 B.n591 B.n28 10.6151
R1803 B.n587 B.n28 10.6151
R1804 B.n587 B.n586 10.6151
R1805 B.n586 B.n585 10.6151
R1806 B.n585 B.n30 10.6151
R1807 B.n581 B.n30 10.6151
R1808 B.n581 B.n580 10.6151
R1809 B.n580 B.n579 10.6151
R1810 B.n579 B.n32 10.6151
R1811 B.n575 B.n32 10.6151
R1812 B.n575 B.n574 10.6151
R1813 B.n574 B.n573 10.6151
R1814 B.n573 B.n34 10.6151
R1815 B.n569 B.n34 10.6151
R1816 B.n569 B.n568 10.6151
R1817 B.n568 B.n567 10.6151
R1818 B.n567 B.n36 10.6151
R1819 B.n563 B.n36 10.6151
R1820 B.n563 B.n562 10.6151
R1821 B.n562 B.n561 10.6151
R1822 B.n561 B.n38 10.6151
R1823 B.n557 B.n38 10.6151
R1824 B.n557 B.n556 10.6151
R1825 B.n556 B.n555 10.6151
R1826 B.n555 B.n40 10.6151
R1827 B.n551 B.n550 10.6151
R1828 B.n550 B.n549 10.6151
R1829 B.n549 B.n45 10.6151
R1830 B.n545 B.n45 10.6151
R1831 B.n545 B.n544 10.6151
R1832 B.n544 B.n543 10.6151
R1833 B.n543 B.n47 10.6151
R1834 B.n539 B.n47 10.6151
R1835 B.n537 B.n536 10.6151
R1836 B.n536 B.n51 10.6151
R1837 B.n532 B.n51 10.6151
R1838 B.n532 B.n531 10.6151
R1839 B.n531 B.n530 10.6151
R1840 B.n530 B.n53 10.6151
R1841 B.n526 B.n53 10.6151
R1842 B.n526 B.n525 10.6151
R1843 B.n525 B.n524 10.6151
R1844 B.n524 B.n55 10.6151
R1845 B.n520 B.n55 10.6151
R1846 B.n520 B.n519 10.6151
R1847 B.n519 B.n518 10.6151
R1848 B.n518 B.n57 10.6151
R1849 B.n514 B.n57 10.6151
R1850 B.n514 B.n513 10.6151
R1851 B.n513 B.n512 10.6151
R1852 B.n512 B.n59 10.6151
R1853 B.n508 B.n59 10.6151
R1854 B.n508 B.n507 10.6151
R1855 B.n507 B.n506 10.6151
R1856 B.n506 B.n61 10.6151
R1857 B.n502 B.n61 10.6151
R1858 B.n502 B.n501 10.6151
R1859 B.n501 B.n500 10.6151
R1860 B.n500 B.n63 10.6151
R1861 B.n496 B.n63 10.6151
R1862 B.n496 B.n495 10.6151
R1863 B.n495 B.n494 10.6151
R1864 B.n494 B.n65 10.6151
R1865 B.n490 B.n65 10.6151
R1866 B.n490 B.n489 10.6151
R1867 B.n489 B.n488 10.6151
R1868 B.n488 B.n67 10.6151
R1869 B.n484 B.n67 10.6151
R1870 B.n484 B.n483 10.6151
R1871 B.n483 B.n482 10.6151
R1872 B.n482 B.n69 10.6151
R1873 B.n478 B.n69 10.6151
R1874 B.n478 B.n477 10.6151
R1875 B.n477 B.n476 10.6151
R1876 B.n476 B.n71 10.6151
R1877 B.n472 B.n71 10.6151
R1878 B.n472 B.n471 10.6151
R1879 B.n471 B.n470 10.6151
R1880 B.n466 B.n73 10.6151
R1881 B.n466 B.n465 10.6151
R1882 B.n465 B.n464 10.6151
R1883 B.n464 B.n75 10.6151
R1884 B.n460 B.n75 10.6151
R1885 B.n460 B.n459 10.6151
R1886 B.n459 B.n458 10.6151
R1887 B.n458 B.n77 10.6151
R1888 B.n454 B.n77 10.6151
R1889 B.n454 B.n453 10.6151
R1890 B.n453 B.n452 10.6151
R1891 B.n452 B.n79 10.6151
R1892 B.n448 B.n79 10.6151
R1893 B.n448 B.n447 10.6151
R1894 B.n447 B.n446 10.6151
R1895 B.n446 B.n81 10.6151
R1896 B.n442 B.n81 10.6151
R1897 B.n442 B.n441 10.6151
R1898 B.n441 B.n440 10.6151
R1899 B.n440 B.n83 10.6151
R1900 B.n436 B.n83 10.6151
R1901 B.n436 B.n435 10.6151
R1902 B.n435 B.n434 10.6151
R1903 B.n434 B.n85 10.6151
R1904 B.n430 B.n85 10.6151
R1905 B.n430 B.n429 10.6151
R1906 B.n429 B.n428 10.6151
R1907 B.n428 B.n87 10.6151
R1908 B.n424 B.n87 10.6151
R1909 B.n424 B.n423 10.6151
R1910 B.n423 B.n422 10.6151
R1911 B.n422 B.n89 10.6151
R1912 B.n418 B.n89 10.6151
R1913 B.n418 B.n417 10.6151
R1914 B.n417 B.n416 10.6151
R1915 B.n416 B.n91 10.6151
R1916 B.n412 B.n91 10.6151
R1917 B.n412 B.n411 10.6151
R1918 B.n411 B.n410 10.6151
R1919 B.n410 B.n93 10.6151
R1920 B.n406 B.n93 10.6151
R1921 B.n406 B.n405 10.6151
R1922 B.n405 B.n404 10.6151
R1923 B.n404 B.n95 10.6151
R1924 B.n400 B.n95 10.6151
R1925 B.n400 B.n399 10.6151
R1926 B.n399 B.n398 10.6151
R1927 B.n398 B.n97 10.6151
R1928 B.n394 B.n97 10.6151
R1929 B.n394 B.n393 10.6151
R1930 B.n393 B.n392 10.6151
R1931 B.n392 B.n99 10.6151
R1932 B.n388 B.n99 10.6151
R1933 B.n388 B.n387 10.6151
R1934 B.n387 B.n386 10.6151
R1935 B.n386 B.n101 10.6151
R1936 B.n382 B.n101 10.6151
R1937 B.n382 B.n381 10.6151
R1938 B.n381 B.n380 10.6151
R1939 B.n380 B.n103 10.6151
R1940 B.n376 B.n103 10.6151
R1941 B.n376 B.n375 10.6151
R1942 B.n375 B.n374 10.6151
R1943 B.n175 B.n1 10.6151
R1944 B.n176 B.n175 10.6151
R1945 B.n176 B.n173 10.6151
R1946 B.n180 B.n173 10.6151
R1947 B.n181 B.n180 10.6151
R1948 B.n182 B.n181 10.6151
R1949 B.n182 B.n171 10.6151
R1950 B.n186 B.n171 10.6151
R1951 B.n187 B.n186 10.6151
R1952 B.n188 B.n187 10.6151
R1953 B.n188 B.n169 10.6151
R1954 B.n192 B.n169 10.6151
R1955 B.n193 B.n192 10.6151
R1956 B.n194 B.n193 10.6151
R1957 B.n194 B.n167 10.6151
R1958 B.n198 B.n167 10.6151
R1959 B.n199 B.n198 10.6151
R1960 B.n200 B.n199 10.6151
R1961 B.n200 B.n165 10.6151
R1962 B.n204 B.n165 10.6151
R1963 B.n205 B.n204 10.6151
R1964 B.n206 B.n205 10.6151
R1965 B.n206 B.n163 10.6151
R1966 B.n210 B.n163 10.6151
R1967 B.n211 B.n210 10.6151
R1968 B.n212 B.n211 10.6151
R1969 B.n212 B.n161 10.6151
R1970 B.n216 B.n161 10.6151
R1971 B.n217 B.n216 10.6151
R1972 B.n218 B.n217 10.6151
R1973 B.n222 B.n159 10.6151
R1974 B.n223 B.n222 10.6151
R1975 B.n224 B.n223 10.6151
R1976 B.n224 B.n157 10.6151
R1977 B.n228 B.n157 10.6151
R1978 B.n229 B.n228 10.6151
R1979 B.n230 B.n229 10.6151
R1980 B.n230 B.n155 10.6151
R1981 B.n234 B.n155 10.6151
R1982 B.n235 B.n234 10.6151
R1983 B.n236 B.n235 10.6151
R1984 B.n236 B.n153 10.6151
R1985 B.n240 B.n153 10.6151
R1986 B.n241 B.n240 10.6151
R1987 B.n242 B.n241 10.6151
R1988 B.n242 B.n151 10.6151
R1989 B.n246 B.n151 10.6151
R1990 B.n247 B.n246 10.6151
R1991 B.n248 B.n247 10.6151
R1992 B.n248 B.n149 10.6151
R1993 B.n252 B.n149 10.6151
R1994 B.n253 B.n252 10.6151
R1995 B.n254 B.n253 10.6151
R1996 B.n254 B.n147 10.6151
R1997 B.n258 B.n147 10.6151
R1998 B.n259 B.n258 10.6151
R1999 B.n260 B.n259 10.6151
R2000 B.n260 B.n145 10.6151
R2001 B.n264 B.n145 10.6151
R2002 B.n265 B.n264 10.6151
R2003 B.n266 B.n265 10.6151
R2004 B.n266 B.n143 10.6151
R2005 B.n270 B.n143 10.6151
R2006 B.n271 B.n270 10.6151
R2007 B.n272 B.n271 10.6151
R2008 B.n272 B.n141 10.6151
R2009 B.n276 B.n141 10.6151
R2010 B.n277 B.n276 10.6151
R2011 B.n278 B.n277 10.6151
R2012 B.n278 B.n139 10.6151
R2013 B.n282 B.n139 10.6151
R2014 B.n283 B.n282 10.6151
R2015 B.n284 B.n283 10.6151
R2016 B.n284 B.n137 10.6151
R2017 B.n288 B.n137 10.6151
R2018 B.n291 B.n290 10.6151
R2019 B.n291 B.n133 10.6151
R2020 B.n295 B.n133 10.6151
R2021 B.n296 B.n295 10.6151
R2022 B.n297 B.n296 10.6151
R2023 B.n297 B.n131 10.6151
R2024 B.n301 B.n131 10.6151
R2025 B.n302 B.n301 10.6151
R2026 B.n304 B.n127 10.6151
R2027 B.n308 B.n127 10.6151
R2028 B.n309 B.n308 10.6151
R2029 B.n310 B.n309 10.6151
R2030 B.n310 B.n125 10.6151
R2031 B.n314 B.n125 10.6151
R2032 B.n315 B.n314 10.6151
R2033 B.n316 B.n315 10.6151
R2034 B.n316 B.n123 10.6151
R2035 B.n320 B.n123 10.6151
R2036 B.n321 B.n320 10.6151
R2037 B.n322 B.n321 10.6151
R2038 B.n322 B.n121 10.6151
R2039 B.n326 B.n121 10.6151
R2040 B.n327 B.n326 10.6151
R2041 B.n328 B.n327 10.6151
R2042 B.n328 B.n119 10.6151
R2043 B.n332 B.n119 10.6151
R2044 B.n333 B.n332 10.6151
R2045 B.n334 B.n333 10.6151
R2046 B.n334 B.n117 10.6151
R2047 B.n338 B.n117 10.6151
R2048 B.n339 B.n338 10.6151
R2049 B.n340 B.n339 10.6151
R2050 B.n340 B.n115 10.6151
R2051 B.n344 B.n115 10.6151
R2052 B.n345 B.n344 10.6151
R2053 B.n346 B.n345 10.6151
R2054 B.n346 B.n113 10.6151
R2055 B.n350 B.n113 10.6151
R2056 B.n351 B.n350 10.6151
R2057 B.n352 B.n351 10.6151
R2058 B.n352 B.n111 10.6151
R2059 B.n356 B.n111 10.6151
R2060 B.n357 B.n356 10.6151
R2061 B.n358 B.n357 10.6151
R2062 B.n358 B.n109 10.6151
R2063 B.n362 B.n109 10.6151
R2064 B.n363 B.n362 10.6151
R2065 B.n364 B.n363 10.6151
R2066 B.n364 B.n107 10.6151
R2067 B.n368 B.n107 10.6151
R2068 B.n369 B.n368 10.6151
R2069 B.n370 B.n369 10.6151
R2070 B.n370 B.n105 10.6151
R2071 B.n669 B.n0 8.11757
R2072 B.n669 B.n1 8.11757
R2073 B.n551 B.n44 6.5566
R2074 B.n539 B.n538 6.5566
R2075 B.n290 B.n289 6.5566
R2076 B.n303 B.n302 6.5566
R2077 B.n44 B.n40 4.05904
R2078 B.n538 B.n537 4.05904
R2079 B.n289 B.n288 4.05904
R2080 B.n304 B.n303 4.05904
C0 VN VDD1 0.149699f
C1 VP w_n2578_n3654# 5.38684f
C2 B VDD1 1.94322f
C3 VDD2 w_n2578_n3654# 2.33751f
C4 VDD2 VP 0.381163f
C5 VTAIL VN 8.79786f
C6 VTAIL B 3.20202f
C7 w_n2578_n3654# VDD1 2.27659f
C8 VP VDD1 9.100691f
C9 B VN 0.895045f
C10 VDD2 VDD1 1.16782f
C11 VTAIL w_n2578_n3654# 3.24884f
C12 VTAIL VP 8.81243f
C13 VDD2 VTAIL 13.425f
C14 w_n2578_n3654# VN 5.05611f
C15 VP VN 6.31928f
C16 B w_n2578_n3654# 8.2743f
C17 VP B 1.44243f
C18 VTAIL VDD1 13.3884f
C19 VDD2 VN 8.87405f
C20 VDD2 B 1.9994f
C21 VDD2 VSUBS 1.545862f
C22 VDD1 VSUBS 1.322206f
C23 VTAIL VSUBS 0.932902f
C24 VN VSUBS 5.40042f
C25 VP VSUBS 2.286016f
C26 B VSUBS 3.514493f
C27 w_n2578_n3654# VSUBS 0.115732p
C28 B.n0 VSUBS 0.006088f
C29 B.n1 VSUBS 0.006088f
C30 B.n2 VSUBS 0.009003f
C31 B.n3 VSUBS 0.006899f
C32 B.n4 VSUBS 0.006899f
C33 B.n5 VSUBS 0.006899f
C34 B.n6 VSUBS 0.006899f
C35 B.n7 VSUBS 0.006899f
C36 B.n8 VSUBS 0.006899f
C37 B.n9 VSUBS 0.006899f
C38 B.n10 VSUBS 0.006899f
C39 B.n11 VSUBS 0.006899f
C40 B.n12 VSUBS 0.006899f
C41 B.n13 VSUBS 0.006899f
C42 B.n14 VSUBS 0.006899f
C43 B.n15 VSUBS 0.006899f
C44 B.n16 VSUBS 0.006899f
C45 B.n17 VSUBS 0.016912f
C46 B.n18 VSUBS 0.006899f
C47 B.n19 VSUBS 0.006899f
C48 B.n20 VSUBS 0.006899f
C49 B.n21 VSUBS 0.006899f
C50 B.n22 VSUBS 0.006899f
C51 B.n23 VSUBS 0.006899f
C52 B.n24 VSUBS 0.006899f
C53 B.n25 VSUBS 0.006899f
C54 B.n26 VSUBS 0.006899f
C55 B.n27 VSUBS 0.006899f
C56 B.n28 VSUBS 0.006899f
C57 B.n29 VSUBS 0.006899f
C58 B.n30 VSUBS 0.006899f
C59 B.n31 VSUBS 0.006899f
C60 B.n32 VSUBS 0.006899f
C61 B.n33 VSUBS 0.006899f
C62 B.n34 VSUBS 0.006899f
C63 B.n35 VSUBS 0.006899f
C64 B.n36 VSUBS 0.006899f
C65 B.n37 VSUBS 0.006899f
C66 B.n38 VSUBS 0.006899f
C67 B.n39 VSUBS 0.006899f
C68 B.n40 VSUBS 0.004769f
C69 B.n41 VSUBS 0.006899f
C70 B.t7 VSUBS 0.23979f
C71 B.t8 VSUBS 0.255056f
C72 B.t6 VSUBS 0.562448f
C73 B.n42 VSUBS 0.361f
C74 B.n43 VSUBS 0.26088f
C75 B.n44 VSUBS 0.015985f
C76 B.n45 VSUBS 0.006899f
C77 B.n46 VSUBS 0.006899f
C78 B.n47 VSUBS 0.006899f
C79 B.n48 VSUBS 0.006899f
C80 B.t4 VSUBS 0.239794f
C81 B.t5 VSUBS 0.255059f
C82 B.t3 VSUBS 0.562448f
C83 B.n49 VSUBS 0.360997f
C84 B.n50 VSUBS 0.260877f
C85 B.n51 VSUBS 0.006899f
C86 B.n52 VSUBS 0.006899f
C87 B.n53 VSUBS 0.006899f
C88 B.n54 VSUBS 0.006899f
C89 B.n55 VSUBS 0.006899f
C90 B.n56 VSUBS 0.006899f
C91 B.n57 VSUBS 0.006899f
C92 B.n58 VSUBS 0.006899f
C93 B.n59 VSUBS 0.006899f
C94 B.n60 VSUBS 0.006899f
C95 B.n61 VSUBS 0.006899f
C96 B.n62 VSUBS 0.006899f
C97 B.n63 VSUBS 0.006899f
C98 B.n64 VSUBS 0.006899f
C99 B.n65 VSUBS 0.006899f
C100 B.n66 VSUBS 0.006899f
C101 B.n67 VSUBS 0.006899f
C102 B.n68 VSUBS 0.006899f
C103 B.n69 VSUBS 0.006899f
C104 B.n70 VSUBS 0.006899f
C105 B.n71 VSUBS 0.006899f
C106 B.n72 VSUBS 0.006899f
C107 B.n73 VSUBS 0.016912f
C108 B.n74 VSUBS 0.006899f
C109 B.n75 VSUBS 0.006899f
C110 B.n76 VSUBS 0.006899f
C111 B.n77 VSUBS 0.006899f
C112 B.n78 VSUBS 0.006899f
C113 B.n79 VSUBS 0.006899f
C114 B.n80 VSUBS 0.006899f
C115 B.n81 VSUBS 0.006899f
C116 B.n82 VSUBS 0.006899f
C117 B.n83 VSUBS 0.006899f
C118 B.n84 VSUBS 0.006899f
C119 B.n85 VSUBS 0.006899f
C120 B.n86 VSUBS 0.006899f
C121 B.n87 VSUBS 0.006899f
C122 B.n88 VSUBS 0.006899f
C123 B.n89 VSUBS 0.006899f
C124 B.n90 VSUBS 0.006899f
C125 B.n91 VSUBS 0.006899f
C126 B.n92 VSUBS 0.006899f
C127 B.n93 VSUBS 0.006899f
C128 B.n94 VSUBS 0.006899f
C129 B.n95 VSUBS 0.006899f
C130 B.n96 VSUBS 0.006899f
C131 B.n97 VSUBS 0.006899f
C132 B.n98 VSUBS 0.006899f
C133 B.n99 VSUBS 0.006899f
C134 B.n100 VSUBS 0.006899f
C135 B.n101 VSUBS 0.006899f
C136 B.n102 VSUBS 0.006899f
C137 B.n103 VSUBS 0.006899f
C138 B.n104 VSUBS 0.006899f
C139 B.n105 VSUBS 0.017055f
C140 B.n106 VSUBS 0.006899f
C141 B.n107 VSUBS 0.006899f
C142 B.n108 VSUBS 0.006899f
C143 B.n109 VSUBS 0.006899f
C144 B.n110 VSUBS 0.006899f
C145 B.n111 VSUBS 0.006899f
C146 B.n112 VSUBS 0.006899f
C147 B.n113 VSUBS 0.006899f
C148 B.n114 VSUBS 0.006899f
C149 B.n115 VSUBS 0.006899f
C150 B.n116 VSUBS 0.006899f
C151 B.n117 VSUBS 0.006899f
C152 B.n118 VSUBS 0.006899f
C153 B.n119 VSUBS 0.006899f
C154 B.n120 VSUBS 0.006899f
C155 B.n121 VSUBS 0.006899f
C156 B.n122 VSUBS 0.006899f
C157 B.n123 VSUBS 0.006899f
C158 B.n124 VSUBS 0.006899f
C159 B.n125 VSUBS 0.006899f
C160 B.n126 VSUBS 0.006899f
C161 B.n127 VSUBS 0.006899f
C162 B.n128 VSUBS 0.006899f
C163 B.t11 VSUBS 0.239794f
C164 B.t10 VSUBS 0.255059f
C165 B.t9 VSUBS 0.562448f
C166 B.n129 VSUBS 0.360997f
C167 B.n130 VSUBS 0.260877f
C168 B.n131 VSUBS 0.006899f
C169 B.n132 VSUBS 0.006899f
C170 B.n133 VSUBS 0.006899f
C171 B.n134 VSUBS 0.006899f
C172 B.t2 VSUBS 0.23979f
C173 B.t1 VSUBS 0.255056f
C174 B.t0 VSUBS 0.562448f
C175 B.n135 VSUBS 0.361f
C176 B.n136 VSUBS 0.26088f
C177 B.n137 VSUBS 0.006899f
C178 B.n138 VSUBS 0.006899f
C179 B.n139 VSUBS 0.006899f
C180 B.n140 VSUBS 0.006899f
C181 B.n141 VSUBS 0.006899f
C182 B.n142 VSUBS 0.006899f
C183 B.n143 VSUBS 0.006899f
C184 B.n144 VSUBS 0.006899f
C185 B.n145 VSUBS 0.006899f
C186 B.n146 VSUBS 0.006899f
C187 B.n147 VSUBS 0.006899f
C188 B.n148 VSUBS 0.006899f
C189 B.n149 VSUBS 0.006899f
C190 B.n150 VSUBS 0.006899f
C191 B.n151 VSUBS 0.006899f
C192 B.n152 VSUBS 0.006899f
C193 B.n153 VSUBS 0.006899f
C194 B.n154 VSUBS 0.006899f
C195 B.n155 VSUBS 0.006899f
C196 B.n156 VSUBS 0.006899f
C197 B.n157 VSUBS 0.006899f
C198 B.n158 VSUBS 0.006899f
C199 B.n159 VSUBS 0.017787f
C200 B.n160 VSUBS 0.006899f
C201 B.n161 VSUBS 0.006899f
C202 B.n162 VSUBS 0.006899f
C203 B.n163 VSUBS 0.006899f
C204 B.n164 VSUBS 0.006899f
C205 B.n165 VSUBS 0.006899f
C206 B.n166 VSUBS 0.006899f
C207 B.n167 VSUBS 0.006899f
C208 B.n168 VSUBS 0.006899f
C209 B.n169 VSUBS 0.006899f
C210 B.n170 VSUBS 0.006899f
C211 B.n171 VSUBS 0.006899f
C212 B.n172 VSUBS 0.006899f
C213 B.n173 VSUBS 0.006899f
C214 B.n174 VSUBS 0.006899f
C215 B.n175 VSUBS 0.006899f
C216 B.n176 VSUBS 0.006899f
C217 B.n177 VSUBS 0.006899f
C218 B.n178 VSUBS 0.006899f
C219 B.n179 VSUBS 0.006899f
C220 B.n180 VSUBS 0.006899f
C221 B.n181 VSUBS 0.006899f
C222 B.n182 VSUBS 0.006899f
C223 B.n183 VSUBS 0.006899f
C224 B.n184 VSUBS 0.006899f
C225 B.n185 VSUBS 0.006899f
C226 B.n186 VSUBS 0.006899f
C227 B.n187 VSUBS 0.006899f
C228 B.n188 VSUBS 0.006899f
C229 B.n189 VSUBS 0.006899f
C230 B.n190 VSUBS 0.006899f
C231 B.n191 VSUBS 0.006899f
C232 B.n192 VSUBS 0.006899f
C233 B.n193 VSUBS 0.006899f
C234 B.n194 VSUBS 0.006899f
C235 B.n195 VSUBS 0.006899f
C236 B.n196 VSUBS 0.006899f
C237 B.n197 VSUBS 0.006899f
C238 B.n198 VSUBS 0.006899f
C239 B.n199 VSUBS 0.006899f
C240 B.n200 VSUBS 0.006899f
C241 B.n201 VSUBS 0.006899f
C242 B.n202 VSUBS 0.006899f
C243 B.n203 VSUBS 0.006899f
C244 B.n204 VSUBS 0.006899f
C245 B.n205 VSUBS 0.006899f
C246 B.n206 VSUBS 0.006899f
C247 B.n207 VSUBS 0.006899f
C248 B.n208 VSUBS 0.006899f
C249 B.n209 VSUBS 0.006899f
C250 B.n210 VSUBS 0.006899f
C251 B.n211 VSUBS 0.006899f
C252 B.n212 VSUBS 0.006899f
C253 B.n213 VSUBS 0.006899f
C254 B.n214 VSUBS 0.006899f
C255 B.n215 VSUBS 0.006899f
C256 B.n216 VSUBS 0.006899f
C257 B.n217 VSUBS 0.006899f
C258 B.n218 VSUBS 0.016912f
C259 B.n219 VSUBS 0.016912f
C260 B.n220 VSUBS 0.017787f
C261 B.n221 VSUBS 0.006899f
C262 B.n222 VSUBS 0.006899f
C263 B.n223 VSUBS 0.006899f
C264 B.n224 VSUBS 0.006899f
C265 B.n225 VSUBS 0.006899f
C266 B.n226 VSUBS 0.006899f
C267 B.n227 VSUBS 0.006899f
C268 B.n228 VSUBS 0.006899f
C269 B.n229 VSUBS 0.006899f
C270 B.n230 VSUBS 0.006899f
C271 B.n231 VSUBS 0.006899f
C272 B.n232 VSUBS 0.006899f
C273 B.n233 VSUBS 0.006899f
C274 B.n234 VSUBS 0.006899f
C275 B.n235 VSUBS 0.006899f
C276 B.n236 VSUBS 0.006899f
C277 B.n237 VSUBS 0.006899f
C278 B.n238 VSUBS 0.006899f
C279 B.n239 VSUBS 0.006899f
C280 B.n240 VSUBS 0.006899f
C281 B.n241 VSUBS 0.006899f
C282 B.n242 VSUBS 0.006899f
C283 B.n243 VSUBS 0.006899f
C284 B.n244 VSUBS 0.006899f
C285 B.n245 VSUBS 0.006899f
C286 B.n246 VSUBS 0.006899f
C287 B.n247 VSUBS 0.006899f
C288 B.n248 VSUBS 0.006899f
C289 B.n249 VSUBS 0.006899f
C290 B.n250 VSUBS 0.006899f
C291 B.n251 VSUBS 0.006899f
C292 B.n252 VSUBS 0.006899f
C293 B.n253 VSUBS 0.006899f
C294 B.n254 VSUBS 0.006899f
C295 B.n255 VSUBS 0.006899f
C296 B.n256 VSUBS 0.006899f
C297 B.n257 VSUBS 0.006899f
C298 B.n258 VSUBS 0.006899f
C299 B.n259 VSUBS 0.006899f
C300 B.n260 VSUBS 0.006899f
C301 B.n261 VSUBS 0.006899f
C302 B.n262 VSUBS 0.006899f
C303 B.n263 VSUBS 0.006899f
C304 B.n264 VSUBS 0.006899f
C305 B.n265 VSUBS 0.006899f
C306 B.n266 VSUBS 0.006899f
C307 B.n267 VSUBS 0.006899f
C308 B.n268 VSUBS 0.006899f
C309 B.n269 VSUBS 0.006899f
C310 B.n270 VSUBS 0.006899f
C311 B.n271 VSUBS 0.006899f
C312 B.n272 VSUBS 0.006899f
C313 B.n273 VSUBS 0.006899f
C314 B.n274 VSUBS 0.006899f
C315 B.n275 VSUBS 0.006899f
C316 B.n276 VSUBS 0.006899f
C317 B.n277 VSUBS 0.006899f
C318 B.n278 VSUBS 0.006899f
C319 B.n279 VSUBS 0.006899f
C320 B.n280 VSUBS 0.006899f
C321 B.n281 VSUBS 0.006899f
C322 B.n282 VSUBS 0.006899f
C323 B.n283 VSUBS 0.006899f
C324 B.n284 VSUBS 0.006899f
C325 B.n285 VSUBS 0.006899f
C326 B.n286 VSUBS 0.006899f
C327 B.n287 VSUBS 0.006899f
C328 B.n288 VSUBS 0.004769f
C329 B.n289 VSUBS 0.015985f
C330 B.n290 VSUBS 0.00558f
C331 B.n291 VSUBS 0.006899f
C332 B.n292 VSUBS 0.006899f
C333 B.n293 VSUBS 0.006899f
C334 B.n294 VSUBS 0.006899f
C335 B.n295 VSUBS 0.006899f
C336 B.n296 VSUBS 0.006899f
C337 B.n297 VSUBS 0.006899f
C338 B.n298 VSUBS 0.006899f
C339 B.n299 VSUBS 0.006899f
C340 B.n300 VSUBS 0.006899f
C341 B.n301 VSUBS 0.006899f
C342 B.n302 VSUBS 0.00558f
C343 B.n303 VSUBS 0.015985f
C344 B.n304 VSUBS 0.004769f
C345 B.n305 VSUBS 0.006899f
C346 B.n306 VSUBS 0.006899f
C347 B.n307 VSUBS 0.006899f
C348 B.n308 VSUBS 0.006899f
C349 B.n309 VSUBS 0.006899f
C350 B.n310 VSUBS 0.006899f
C351 B.n311 VSUBS 0.006899f
C352 B.n312 VSUBS 0.006899f
C353 B.n313 VSUBS 0.006899f
C354 B.n314 VSUBS 0.006899f
C355 B.n315 VSUBS 0.006899f
C356 B.n316 VSUBS 0.006899f
C357 B.n317 VSUBS 0.006899f
C358 B.n318 VSUBS 0.006899f
C359 B.n319 VSUBS 0.006899f
C360 B.n320 VSUBS 0.006899f
C361 B.n321 VSUBS 0.006899f
C362 B.n322 VSUBS 0.006899f
C363 B.n323 VSUBS 0.006899f
C364 B.n324 VSUBS 0.006899f
C365 B.n325 VSUBS 0.006899f
C366 B.n326 VSUBS 0.006899f
C367 B.n327 VSUBS 0.006899f
C368 B.n328 VSUBS 0.006899f
C369 B.n329 VSUBS 0.006899f
C370 B.n330 VSUBS 0.006899f
C371 B.n331 VSUBS 0.006899f
C372 B.n332 VSUBS 0.006899f
C373 B.n333 VSUBS 0.006899f
C374 B.n334 VSUBS 0.006899f
C375 B.n335 VSUBS 0.006899f
C376 B.n336 VSUBS 0.006899f
C377 B.n337 VSUBS 0.006899f
C378 B.n338 VSUBS 0.006899f
C379 B.n339 VSUBS 0.006899f
C380 B.n340 VSUBS 0.006899f
C381 B.n341 VSUBS 0.006899f
C382 B.n342 VSUBS 0.006899f
C383 B.n343 VSUBS 0.006899f
C384 B.n344 VSUBS 0.006899f
C385 B.n345 VSUBS 0.006899f
C386 B.n346 VSUBS 0.006899f
C387 B.n347 VSUBS 0.006899f
C388 B.n348 VSUBS 0.006899f
C389 B.n349 VSUBS 0.006899f
C390 B.n350 VSUBS 0.006899f
C391 B.n351 VSUBS 0.006899f
C392 B.n352 VSUBS 0.006899f
C393 B.n353 VSUBS 0.006899f
C394 B.n354 VSUBS 0.006899f
C395 B.n355 VSUBS 0.006899f
C396 B.n356 VSUBS 0.006899f
C397 B.n357 VSUBS 0.006899f
C398 B.n358 VSUBS 0.006899f
C399 B.n359 VSUBS 0.006899f
C400 B.n360 VSUBS 0.006899f
C401 B.n361 VSUBS 0.006899f
C402 B.n362 VSUBS 0.006899f
C403 B.n363 VSUBS 0.006899f
C404 B.n364 VSUBS 0.006899f
C405 B.n365 VSUBS 0.006899f
C406 B.n366 VSUBS 0.006899f
C407 B.n367 VSUBS 0.006899f
C408 B.n368 VSUBS 0.006899f
C409 B.n369 VSUBS 0.006899f
C410 B.n370 VSUBS 0.006899f
C411 B.n371 VSUBS 0.006899f
C412 B.n372 VSUBS 0.017787f
C413 B.n373 VSUBS 0.016912f
C414 B.n374 VSUBS 0.017645f
C415 B.n375 VSUBS 0.006899f
C416 B.n376 VSUBS 0.006899f
C417 B.n377 VSUBS 0.006899f
C418 B.n378 VSUBS 0.006899f
C419 B.n379 VSUBS 0.006899f
C420 B.n380 VSUBS 0.006899f
C421 B.n381 VSUBS 0.006899f
C422 B.n382 VSUBS 0.006899f
C423 B.n383 VSUBS 0.006899f
C424 B.n384 VSUBS 0.006899f
C425 B.n385 VSUBS 0.006899f
C426 B.n386 VSUBS 0.006899f
C427 B.n387 VSUBS 0.006899f
C428 B.n388 VSUBS 0.006899f
C429 B.n389 VSUBS 0.006899f
C430 B.n390 VSUBS 0.006899f
C431 B.n391 VSUBS 0.006899f
C432 B.n392 VSUBS 0.006899f
C433 B.n393 VSUBS 0.006899f
C434 B.n394 VSUBS 0.006899f
C435 B.n395 VSUBS 0.006899f
C436 B.n396 VSUBS 0.006899f
C437 B.n397 VSUBS 0.006899f
C438 B.n398 VSUBS 0.006899f
C439 B.n399 VSUBS 0.006899f
C440 B.n400 VSUBS 0.006899f
C441 B.n401 VSUBS 0.006899f
C442 B.n402 VSUBS 0.006899f
C443 B.n403 VSUBS 0.006899f
C444 B.n404 VSUBS 0.006899f
C445 B.n405 VSUBS 0.006899f
C446 B.n406 VSUBS 0.006899f
C447 B.n407 VSUBS 0.006899f
C448 B.n408 VSUBS 0.006899f
C449 B.n409 VSUBS 0.006899f
C450 B.n410 VSUBS 0.006899f
C451 B.n411 VSUBS 0.006899f
C452 B.n412 VSUBS 0.006899f
C453 B.n413 VSUBS 0.006899f
C454 B.n414 VSUBS 0.006899f
C455 B.n415 VSUBS 0.006899f
C456 B.n416 VSUBS 0.006899f
C457 B.n417 VSUBS 0.006899f
C458 B.n418 VSUBS 0.006899f
C459 B.n419 VSUBS 0.006899f
C460 B.n420 VSUBS 0.006899f
C461 B.n421 VSUBS 0.006899f
C462 B.n422 VSUBS 0.006899f
C463 B.n423 VSUBS 0.006899f
C464 B.n424 VSUBS 0.006899f
C465 B.n425 VSUBS 0.006899f
C466 B.n426 VSUBS 0.006899f
C467 B.n427 VSUBS 0.006899f
C468 B.n428 VSUBS 0.006899f
C469 B.n429 VSUBS 0.006899f
C470 B.n430 VSUBS 0.006899f
C471 B.n431 VSUBS 0.006899f
C472 B.n432 VSUBS 0.006899f
C473 B.n433 VSUBS 0.006899f
C474 B.n434 VSUBS 0.006899f
C475 B.n435 VSUBS 0.006899f
C476 B.n436 VSUBS 0.006899f
C477 B.n437 VSUBS 0.006899f
C478 B.n438 VSUBS 0.006899f
C479 B.n439 VSUBS 0.006899f
C480 B.n440 VSUBS 0.006899f
C481 B.n441 VSUBS 0.006899f
C482 B.n442 VSUBS 0.006899f
C483 B.n443 VSUBS 0.006899f
C484 B.n444 VSUBS 0.006899f
C485 B.n445 VSUBS 0.006899f
C486 B.n446 VSUBS 0.006899f
C487 B.n447 VSUBS 0.006899f
C488 B.n448 VSUBS 0.006899f
C489 B.n449 VSUBS 0.006899f
C490 B.n450 VSUBS 0.006899f
C491 B.n451 VSUBS 0.006899f
C492 B.n452 VSUBS 0.006899f
C493 B.n453 VSUBS 0.006899f
C494 B.n454 VSUBS 0.006899f
C495 B.n455 VSUBS 0.006899f
C496 B.n456 VSUBS 0.006899f
C497 B.n457 VSUBS 0.006899f
C498 B.n458 VSUBS 0.006899f
C499 B.n459 VSUBS 0.006899f
C500 B.n460 VSUBS 0.006899f
C501 B.n461 VSUBS 0.006899f
C502 B.n462 VSUBS 0.006899f
C503 B.n463 VSUBS 0.006899f
C504 B.n464 VSUBS 0.006899f
C505 B.n465 VSUBS 0.006899f
C506 B.n466 VSUBS 0.006899f
C507 B.n467 VSUBS 0.006899f
C508 B.n468 VSUBS 0.016912f
C509 B.n469 VSUBS 0.017787f
C510 B.n470 VSUBS 0.017787f
C511 B.n471 VSUBS 0.006899f
C512 B.n472 VSUBS 0.006899f
C513 B.n473 VSUBS 0.006899f
C514 B.n474 VSUBS 0.006899f
C515 B.n475 VSUBS 0.006899f
C516 B.n476 VSUBS 0.006899f
C517 B.n477 VSUBS 0.006899f
C518 B.n478 VSUBS 0.006899f
C519 B.n479 VSUBS 0.006899f
C520 B.n480 VSUBS 0.006899f
C521 B.n481 VSUBS 0.006899f
C522 B.n482 VSUBS 0.006899f
C523 B.n483 VSUBS 0.006899f
C524 B.n484 VSUBS 0.006899f
C525 B.n485 VSUBS 0.006899f
C526 B.n486 VSUBS 0.006899f
C527 B.n487 VSUBS 0.006899f
C528 B.n488 VSUBS 0.006899f
C529 B.n489 VSUBS 0.006899f
C530 B.n490 VSUBS 0.006899f
C531 B.n491 VSUBS 0.006899f
C532 B.n492 VSUBS 0.006899f
C533 B.n493 VSUBS 0.006899f
C534 B.n494 VSUBS 0.006899f
C535 B.n495 VSUBS 0.006899f
C536 B.n496 VSUBS 0.006899f
C537 B.n497 VSUBS 0.006899f
C538 B.n498 VSUBS 0.006899f
C539 B.n499 VSUBS 0.006899f
C540 B.n500 VSUBS 0.006899f
C541 B.n501 VSUBS 0.006899f
C542 B.n502 VSUBS 0.006899f
C543 B.n503 VSUBS 0.006899f
C544 B.n504 VSUBS 0.006899f
C545 B.n505 VSUBS 0.006899f
C546 B.n506 VSUBS 0.006899f
C547 B.n507 VSUBS 0.006899f
C548 B.n508 VSUBS 0.006899f
C549 B.n509 VSUBS 0.006899f
C550 B.n510 VSUBS 0.006899f
C551 B.n511 VSUBS 0.006899f
C552 B.n512 VSUBS 0.006899f
C553 B.n513 VSUBS 0.006899f
C554 B.n514 VSUBS 0.006899f
C555 B.n515 VSUBS 0.006899f
C556 B.n516 VSUBS 0.006899f
C557 B.n517 VSUBS 0.006899f
C558 B.n518 VSUBS 0.006899f
C559 B.n519 VSUBS 0.006899f
C560 B.n520 VSUBS 0.006899f
C561 B.n521 VSUBS 0.006899f
C562 B.n522 VSUBS 0.006899f
C563 B.n523 VSUBS 0.006899f
C564 B.n524 VSUBS 0.006899f
C565 B.n525 VSUBS 0.006899f
C566 B.n526 VSUBS 0.006899f
C567 B.n527 VSUBS 0.006899f
C568 B.n528 VSUBS 0.006899f
C569 B.n529 VSUBS 0.006899f
C570 B.n530 VSUBS 0.006899f
C571 B.n531 VSUBS 0.006899f
C572 B.n532 VSUBS 0.006899f
C573 B.n533 VSUBS 0.006899f
C574 B.n534 VSUBS 0.006899f
C575 B.n535 VSUBS 0.006899f
C576 B.n536 VSUBS 0.006899f
C577 B.n537 VSUBS 0.004769f
C578 B.n538 VSUBS 0.015985f
C579 B.n539 VSUBS 0.00558f
C580 B.n540 VSUBS 0.006899f
C581 B.n541 VSUBS 0.006899f
C582 B.n542 VSUBS 0.006899f
C583 B.n543 VSUBS 0.006899f
C584 B.n544 VSUBS 0.006899f
C585 B.n545 VSUBS 0.006899f
C586 B.n546 VSUBS 0.006899f
C587 B.n547 VSUBS 0.006899f
C588 B.n548 VSUBS 0.006899f
C589 B.n549 VSUBS 0.006899f
C590 B.n550 VSUBS 0.006899f
C591 B.n551 VSUBS 0.00558f
C592 B.n552 VSUBS 0.006899f
C593 B.n553 VSUBS 0.006899f
C594 B.n554 VSUBS 0.006899f
C595 B.n555 VSUBS 0.006899f
C596 B.n556 VSUBS 0.006899f
C597 B.n557 VSUBS 0.006899f
C598 B.n558 VSUBS 0.006899f
C599 B.n559 VSUBS 0.006899f
C600 B.n560 VSUBS 0.006899f
C601 B.n561 VSUBS 0.006899f
C602 B.n562 VSUBS 0.006899f
C603 B.n563 VSUBS 0.006899f
C604 B.n564 VSUBS 0.006899f
C605 B.n565 VSUBS 0.006899f
C606 B.n566 VSUBS 0.006899f
C607 B.n567 VSUBS 0.006899f
C608 B.n568 VSUBS 0.006899f
C609 B.n569 VSUBS 0.006899f
C610 B.n570 VSUBS 0.006899f
C611 B.n571 VSUBS 0.006899f
C612 B.n572 VSUBS 0.006899f
C613 B.n573 VSUBS 0.006899f
C614 B.n574 VSUBS 0.006899f
C615 B.n575 VSUBS 0.006899f
C616 B.n576 VSUBS 0.006899f
C617 B.n577 VSUBS 0.006899f
C618 B.n578 VSUBS 0.006899f
C619 B.n579 VSUBS 0.006899f
C620 B.n580 VSUBS 0.006899f
C621 B.n581 VSUBS 0.006899f
C622 B.n582 VSUBS 0.006899f
C623 B.n583 VSUBS 0.006899f
C624 B.n584 VSUBS 0.006899f
C625 B.n585 VSUBS 0.006899f
C626 B.n586 VSUBS 0.006899f
C627 B.n587 VSUBS 0.006899f
C628 B.n588 VSUBS 0.006899f
C629 B.n589 VSUBS 0.006899f
C630 B.n590 VSUBS 0.006899f
C631 B.n591 VSUBS 0.006899f
C632 B.n592 VSUBS 0.006899f
C633 B.n593 VSUBS 0.006899f
C634 B.n594 VSUBS 0.006899f
C635 B.n595 VSUBS 0.006899f
C636 B.n596 VSUBS 0.006899f
C637 B.n597 VSUBS 0.006899f
C638 B.n598 VSUBS 0.006899f
C639 B.n599 VSUBS 0.006899f
C640 B.n600 VSUBS 0.006899f
C641 B.n601 VSUBS 0.006899f
C642 B.n602 VSUBS 0.006899f
C643 B.n603 VSUBS 0.006899f
C644 B.n604 VSUBS 0.006899f
C645 B.n605 VSUBS 0.006899f
C646 B.n606 VSUBS 0.006899f
C647 B.n607 VSUBS 0.006899f
C648 B.n608 VSUBS 0.006899f
C649 B.n609 VSUBS 0.006899f
C650 B.n610 VSUBS 0.006899f
C651 B.n611 VSUBS 0.006899f
C652 B.n612 VSUBS 0.006899f
C653 B.n613 VSUBS 0.006899f
C654 B.n614 VSUBS 0.006899f
C655 B.n615 VSUBS 0.006899f
C656 B.n616 VSUBS 0.006899f
C657 B.n617 VSUBS 0.006899f
C658 B.n618 VSUBS 0.006899f
C659 B.n619 VSUBS 0.006899f
C660 B.n620 VSUBS 0.017787f
C661 B.n621 VSUBS 0.017787f
C662 B.n622 VSUBS 0.016912f
C663 B.n623 VSUBS 0.006899f
C664 B.n624 VSUBS 0.006899f
C665 B.n625 VSUBS 0.006899f
C666 B.n626 VSUBS 0.006899f
C667 B.n627 VSUBS 0.006899f
C668 B.n628 VSUBS 0.006899f
C669 B.n629 VSUBS 0.006899f
C670 B.n630 VSUBS 0.006899f
C671 B.n631 VSUBS 0.006899f
C672 B.n632 VSUBS 0.006899f
C673 B.n633 VSUBS 0.006899f
C674 B.n634 VSUBS 0.006899f
C675 B.n635 VSUBS 0.006899f
C676 B.n636 VSUBS 0.006899f
C677 B.n637 VSUBS 0.006899f
C678 B.n638 VSUBS 0.006899f
C679 B.n639 VSUBS 0.006899f
C680 B.n640 VSUBS 0.006899f
C681 B.n641 VSUBS 0.006899f
C682 B.n642 VSUBS 0.006899f
C683 B.n643 VSUBS 0.006899f
C684 B.n644 VSUBS 0.006899f
C685 B.n645 VSUBS 0.006899f
C686 B.n646 VSUBS 0.006899f
C687 B.n647 VSUBS 0.006899f
C688 B.n648 VSUBS 0.006899f
C689 B.n649 VSUBS 0.006899f
C690 B.n650 VSUBS 0.006899f
C691 B.n651 VSUBS 0.006899f
C692 B.n652 VSUBS 0.006899f
C693 B.n653 VSUBS 0.006899f
C694 B.n654 VSUBS 0.006899f
C695 B.n655 VSUBS 0.006899f
C696 B.n656 VSUBS 0.006899f
C697 B.n657 VSUBS 0.006899f
C698 B.n658 VSUBS 0.006899f
C699 B.n659 VSUBS 0.006899f
C700 B.n660 VSUBS 0.006899f
C701 B.n661 VSUBS 0.006899f
C702 B.n662 VSUBS 0.006899f
C703 B.n663 VSUBS 0.006899f
C704 B.n664 VSUBS 0.006899f
C705 B.n665 VSUBS 0.006899f
C706 B.n666 VSUBS 0.006899f
C707 B.n667 VSUBS 0.009003f
C708 B.n668 VSUBS 0.009591f
C709 B.n669 VSUBS 0.019072f
C710 VDD2.n0 VSUBS 0.028643f
C711 VDD2.n1 VSUBS 0.025624f
C712 VDD2.n2 VSUBS 0.013769f
C713 VDD2.n3 VSUBS 0.032546f
C714 VDD2.n4 VSUBS 0.014579f
C715 VDD2.n5 VSUBS 0.025624f
C716 VDD2.n6 VSUBS 0.013769f
C717 VDD2.n7 VSUBS 0.032546f
C718 VDD2.n8 VSUBS 0.014579f
C719 VDD2.n9 VSUBS 0.025624f
C720 VDD2.n10 VSUBS 0.013769f
C721 VDD2.n11 VSUBS 0.032546f
C722 VDD2.n12 VSUBS 0.014579f
C723 VDD2.n13 VSUBS 0.025624f
C724 VDD2.n14 VSUBS 0.013769f
C725 VDD2.n15 VSUBS 0.032546f
C726 VDD2.n16 VSUBS 0.014579f
C727 VDD2.n17 VSUBS 0.025624f
C728 VDD2.n18 VSUBS 0.013769f
C729 VDD2.n19 VSUBS 0.032546f
C730 VDD2.n20 VSUBS 0.014579f
C731 VDD2.n21 VSUBS 1.45353f
C732 VDD2.n22 VSUBS 0.013769f
C733 VDD2.t7 VSUBS 0.069576f
C734 VDD2.n23 VSUBS 0.168765f
C735 VDD2.n24 VSUBS 0.020704f
C736 VDD2.n25 VSUBS 0.024409f
C737 VDD2.n26 VSUBS 0.032546f
C738 VDD2.n27 VSUBS 0.014579f
C739 VDD2.n28 VSUBS 0.013769f
C740 VDD2.n29 VSUBS 0.025624f
C741 VDD2.n30 VSUBS 0.025624f
C742 VDD2.n31 VSUBS 0.013769f
C743 VDD2.n32 VSUBS 0.014579f
C744 VDD2.n33 VSUBS 0.032546f
C745 VDD2.n34 VSUBS 0.032546f
C746 VDD2.n35 VSUBS 0.014579f
C747 VDD2.n36 VSUBS 0.013769f
C748 VDD2.n37 VSUBS 0.025624f
C749 VDD2.n38 VSUBS 0.025624f
C750 VDD2.n39 VSUBS 0.013769f
C751 VDD2.n40 VSUBS 0.014579f
C752 VDD2.n41 VSUBS 0.032546f
C753 VDD2.n42 VSUBS 0.032546f
C754 VDD2.n43 VSUBS 0.014579f
C755 VDD2.n44 VSUBS 0.013769f
C756 VDD2.n45 VSUBS 0.025624f
C757 VDD2.n46 VSUBS 0.025624f
C758 VDD2.n47 VSUBS 0.013769f
C759 VDD2.n48 VSUBS 0.014579f
C760 VDD2.n49 VSUBS 0.032546f
C761 VDD2.n50 VSUBS 0.032546f
C762 VDD2.n51 VSUBS 0.014579f
C763 VDD2.n52 VSUBS 0.013769f
C764 VDD2.n53 VSUBS 0.025624f
C765 VDD2.n54 VSUBS 0.025624f
C766 VDD2.n55 VSUBS 0.013769f
C767 VDD2.n56 VSUBS 0.014579f
C768 VDD2.n57 VSUBS 0.032546f
C769 VDD2.n58 VSUBS 0.032546f
C770 VDD2.n59 VSUBS 0.014579f
C771 VDD2.n60 VSUBS 0.013769f
C772 VDD2.n61 VSUBS 0.025624f
C773 VDD2.n62 VSUBS 0.025624f
C774 VDD2.n63 VSUBS 0.013769f
C775 VDD2.n64 VSUBS 0.014579f
C776 VDD2.n65 VSUBS 0.032546f
C777 VDD2.n66 VSUBS 0.082738f
C778 VDD2.n67 VSUBS 0.014579f
C779 VDD2.n68 VSUBS 0.02704f
C780 VDD2.n69 VSUBS 0.067281f
C781 VDD2.n70 VSUBS 0.085194f
C782 VDD2.t5 VSUBS 0.271946f
C783 VDD2.t8 VSUBS 0.271946f
C784 VDD2.n71 VSUBS 2.18736f
C785 VDD2.n72 VSUBS 0.728809f
C786 VDD2.t6 VSUBS 0.271946f
C787 VDD2.t3 VSUBS 0.271946f
C788 VDD2.n73 VSUBS 2.19407f
C789 VDD2.n74 VSUBS 2.46273f
C790 VDD2.n75 VSUBS 0.028643f
C791 VDD2.n76 VSUBS 0.025624f
C792 VDD2.n77 VSUBS 0.013769f
C793 VDD2.n78 VSUBS 0.032546f
C794 VDD2.n79 VSUBS 0.014579f
C795 VDD2.n80 VSUBS 0.025624f
C796 VDD2.n81 VSUBS 0.013769f
C797 VDD2.n82 VSUBS 0.032546f
C798 VDD2.n83 VSUBS 0.014579f
C799 VDD2.n84 VSUBS 0.025624f
C800 VDD2.n85 VSUBS 0.013769f
C801 VDD2.n86 VSUBS 0.032546f
C802 VDD2.n87 VSUBS 0.014579f
C803 VDD2.n88 VSUBS 0.025624f
C804 VDD2.n89 VSUBS 0.013769f
C805 VDD2.n90 VSUBS 0.032546f
C806 VDD2.n91 VSUBS 0.014579f
C807 VDD2.n92 VSUBS 0.025624f
C808 VDD2.n93 VSUBS 0.013769f
C809 VDD2.n94 VSUBS 0.032546f
C810 VDD2.n95 VSUBS 0.014579f
C811 VDD2.n96 VSUBS 1.45353f
C812 VDD2.n97 VSUBS 0.013769f
C813 VDD2.t4 VSUBS 0.069576f
C814 VDD2.n98 VSUBS 0.168765f
C815 VDD2.n99 VSUBS 0.020704f
C816 VDD2.n100 VSUBS 0.024409f
C817 VDD2.n101 VSUBS 0.032546f
C818 VDD2.n102 VSUBS 0.014579f
C819 VDD2.n103 VSUBS 0.013769f
C820 VDD2.n104 VSUBS 0.025624f
C821 VDD2.n105 VSUBS 0.025624f
C822 VDD2.n106 VSUBS 0.013769f
C823 VDD2.n107 VSUBS 0.014579f
C824 VDD2.n108 VSUBS 0.032546f
C825 VDD2.n109 VSUBS 0.032546f
C826 VDD2.n110 VSUBS 0.014579f
C827 VDD2.n111 VSUBS 0.013769f
C828 VDD2.n112 VSUBS 0.025624f
C829 VDD2.n113 VSUBS 0.025624f
C830 VDD2.n114 VSUBS 0.013769f
C831 VDD2.n115 VSUBS 0.014579f
C832 VDD2.n116 VSUBS 0.032546f
C833 VDD2.n117 VSUBS 0.032546f
C834 VDD2.n118 VSUBS 0.014579f
C835 VDD2.n119 VSUBS 0.013769f
C836 VDD2.n120 VSUBS 0.025624f
C837 VDD2.n121 VSUBS 0.025624f
C838 VDD2.n122 VSUBS 0.013769f
C839 VDD2.n123 VSUBS 0.014579f
C840 VDD2.n124 VSUBS 0.032546f
C841 VDD2.n125 VSUBS 0.032546f
C842 VDD2.n126 VSUBS 0.014579f
C843 VDD2.n127 VSUBS 0.013769f
C844 VDD2.n128 VSUBS 0.025624f
C845 VDD2.n129 VSUBS 0.025624f
C846 VDD2.n130 VSUBS 0.013769f
C847 VDD2.n131 VSUBS 0.014579f
C848 VDD2.n132 VSUBS 0.032546f
C849 VDD2.n133 VSUBS 0.032546f
C850 VDD2.n134 VSUBS 0.014579f
C851 VDD2.n135 VSUBS 0.013769f
C852 VDD2.n136 VSUBS 0.025624f
C853 VDD2.n137 VSUBS 0.025624f
C854 VDD2.n138 VSUBS 0.013769f
C855 VDD2.n139 VSUBS 0.014579f
C856 VDD2.n140 VSUBS 0.032546f
C857 VDD2.n141 VSUBS 0.082738f
C858 VDD2.n142 VSUBS 0.014579f
C859 VDD2.n143 VSUBS 0.02704f
C860 VDD2.n144 VSUBS 0.067281f
C861 VDD2.n145 VSUBS 0.082028f
C862 VDD2.n146 VSUBS 2.44916f
C863 VDD2.t1 VSUBS 0.271946f
C864 VDD2.t9 VSUBS 0.271946f
C865 VDD2.n147 VSUBS 2.18737f
C866 VDD2.n148 VSUBS 0.589462f
C867 VDD2.t0 VSUBS 0.271946f
C868 VDD2.t2 VSUBS 0.271946f
C869 VDD2.n149 VSUBS 2.19404f
C870 VN.n0 VSUBS 0.059087f
C871 VN.t3 VSUBS 1.64149f
C872 VN.n1 VSUBS 0.039576f
C873 VN.n2 VSUBS 0.044281f
C874 VN.t1 VSUBS 1.64149f
C875 VN.n3 VSUBS 0.055899f
C876 VN.t2 VSUBS 1.73596f
C877 VN.t4 VSUBS 1.64149f
C878 VN.n4 VSUBS 0.63575f
C879 VN.n5 VSUBS 0.668242f
C880 VN.n6 VSUBS 0.186322f
C881 VN.n7 VSUBS 0.044281f
C882 VN.n8 VSUBS 0.039576f
C883 VN.n9 VSUBS 0.062554f
C884 VN.n10 VSUBS 0.601835f
C885 VN.n11 VSUBS 0.062554f
C886 VN.n12 VSUBS 0.044281f
C887 VN.n13 VSUBS 0.044281f
C888 VN.n14 VSUBS 0.044281f
C889 VN.n15 VSUBS 0.055899f
C890 VN.n16 VSUBS 0.601835f
C891 VN.n17 VSUBS 0.057465f
C892 VN.t6 VSUBS 1.71001f
C893 VN.n18 VSUBS 0.669742f
C894 VN.n19 VSUBS 0.041471f
C895 VN.n20 VSUBS 0.059087f
C896 VN.t8 VSUBS 1.64149f
C897 VN.n21 VSUBS 0.039576f
C898 VN.n22 VSUBS 0.044281f
C899 VN.t0 VSUBS 1.64149f
C900 VN.n23 VSUBS 0.055899f
C901 VN.t7 VSUBS 1.73596f
C902 VN.t9 VSUBS 1.64149f
C903 VN.n24 VSUBS 0.63575f
C904 VN.n25 VSUBS 0.668242f
C905 VN.n26 VSUBS 0.186322f
C906 VN.n27 VSUBS 0.044281f
C907 VN.n28 VSUBS 0.039576f
C908 VN.n29 VSUBS 0.062554f
C909 VN.n30 VSUBS 0.601835f
C910 VN.n31 VSUBS 0.062554f
C911 VN.n32 VSUBS 0.044281f
C912 VN.n33 VSUBS 0.044281f
C913 VN.n34 VSUBS 0.044281f
C914 VN.n35 VSUBS 0.055899f
C915 VN.n36 VSUBS 0.601835f
C916 VN.n37 VSUBS 0.057465f
C917 VN.t5 VSUBS 1.71001f
C918 VN.n38 VSUBS 0.669742f
C919 VN.n39 VSUBS 2.13777f
C920 VDD1.n0 VSUBS 0.028765f
C921 VDD1.n1 VSUBS 0.025734f
C922 VDD1.n2 VSUBS 0.013828f
C923 VDD1.n3 VSUBS 0.032685f
C924 VDD1.n4 VSUBS 0.014642f
C925 VDD1.n5 VSUBS 0.025734f
C926 VDD1.n6 VSUBS 0.013828f
C927 VDD1.n7 VSUBS 0.032685f
C928 VDD1.n8 VSUBS 0.014642f
C929 VDD1.n9 VSUBS 0.025734f
C930 VDD1.n10 VSUBS 0.013828f
C931 VDD1.n11 VSUBS 0.032685f
C932 VDD1.n12 VSUBS 0.014642f
C933 VDD1.n13 VSUBS 0.025734f
C934 VDD1.n14 VSUBS 0.013828f
C935 VDD1.n15 VSUBS 0.032685f
C936 VDD1.n16 VSUBS 0.014642f
C937 VDD1.n17 VSUBS 0.025734f
C938 VDD1.n18 VSUBS 0.013828f
C939 VDD1.n19 VSUBS 0.032685f
C940 VDD1.n20 VSUBS 0.014642f
C941 VDD1.n21 VSUBS 1.45973f
C942 VDD1.n22 VSUBS 0.013828f
C943 VDD1.t9 VSUBS 0.069872f
C944 VDD1.n23 VSUBS 0.169485f
C945 VDD1.n24 VSUBS 0.020792f
C946 VDD1.n25 VSUBS 0.024514f
C947 VDD1.n26 VSUBS 0.032685f
C948 VDD1.n27 VSUBS 0.014642f
C949 VDD1.n28 VSUBS 0.013828f
C950 VDD1.n29 VSUBS 0.025734f
C951 VDD1.n30 VSUBS 0.025734f
C952 VDD1.n31 VSUBS 0.013828f
C953 VDD1.n32 VSUBS 0.014642f
C954 VDD1.n33 VSUBS 0.032685f
C955 VDD1.n34 VSUBS 0.032685f
C956 VDD1.n35 VSUBS 0.014642f
C957 VDD1.n36 VSUBS 0.013828f
C958 VDD1.n37 VSUBS 0.025734f
C959 VDD1.n38 VSUBS 0.025734f
C960 VDD1.n39 VSUBS 0.013828f
C961 VDD1.n40 VSUBS 0.014642f
C962 VDD1.n41 VSUBS 0.032685f
C963 VDD1.n42 VSUBS 0.032685f
C964 VDD1.n43 VSUBS 0.014642f
C965 VDD1.n44 VSUBS 0.013828f
C966 VDD1.n45 VSUBS 0.025734f
C967 VDD1.n46 VSUBS 0.025734f
C968 VDD1.n47 VSUBS 0.013828f
C969 VDD1.n48 VSUBS 0.014642f
C970 VDD1.n49 VSUBS 0.032685f
C971 VDD1.n50 VSUBS 0.032685f
C972 VDD1.n51 VSUBS 0.014642f
C973 VDD1.n52 VSUBS 0.013828f
C974 VDD1.n53 VSUBS 0.025734f
C975 VDD1.n54 VSUBS 0.025734f
C976 VDD1.n55 VSUBS 0.013828f
C977 VDD1.n56 VSUBS 0.014642f
C978 VDD1.n57 VSUBS 0.032685f
C979 VDD1.n58 VSUBS 0.032685f
C980 VDD1.n59 VSUBS 0.014642f
C981 VDD1.n60 VSUBS 0.013828f
C982 VDD1.n61 VSUBS 0.025734f
C983 VDD1.n62 VSUBS 0.025734f
C984 VDD1.n63 VSUBS 0.013828f
C985 VDD1.n64 VSUBS 0.014642f
C986 VDD1.n65 VSUBS 0.032685f
C987 VDD1.n66 VSUBS 0.083091f
C988 VDD1.n67 VSUBS 0.014642f
C989 VDD1.n68 VSUBS 0.027155f
C990 VDD1.n69 VSUBS 0.067568f
C991 VDD1.n70 VSUBS 0.085557f
C992 VDD1.t7 VSUBS 0.273106f
C993 VDD1.t0 VSUBS 0.273106f
C994 VDD1.n71 VSUBS 2.19671f
C995 VDD1.n72 VSUBS 0.738767f
C996 VDD1.n73 VSUBS 0.028765f
C997 VDD1.n74 VSUBS 0.025734f
C998 VDD1.n75 VSUBS 0.013828f
C999 VDD1.n76 VSUBS 0.032685f
C1000 VDD1.n77 VSUBS 0.014642f
C1001 VDD1.n78 VSUBS 0.025734f
C1002 VDD1.n79 VSUBS 0.013828f
C1003 VDD1.n80 VSUBS 0.032685f
C1004 VDD1.n81 VSUBS 0.014642f
C1005 VDD1.n82 VSUBS 0.025734f
C1006 VDD1.n83 VSUBS 0.013828f
C1007 VDD1.n84 VSUBS 0.032685f
C1008 VDD1.n85 VSUBS 0.014642f
C1009 VDD1.n86 VSUBS 0.025734f
C1010 VDD1.n87 VSUBS 0.013828f
C1011 VDD1.n88 VSUBS 0.032685f
C1012 VDD1.n89 VSUBS 0.014642f
C1013 VDD1.n90 VSUBS 0.025734f
C1014 VDD1.n91 VSUBS 0.013828f
C1015 VDD1.n92 VSUBS 0.032685f
C1016 VDD1.n93 VSUBS 0.014642f
C1017 VDD1.n94 VSUBS 1.45973f
C1018 VDD1.n95 VSUBS 0.013828f
C1019 VDD1.t6 VSUBS 0.069872f
C1020 VDD1.n96 VSUBS 0.169485f
C1021 VDD1.n97 VSUBS 0.020792f
C1022 VDD1.n98 VSUBS 0.024514f
C1023 VDD1.n99 VSUBS 0.032685f
C1024 VDD1.n100 VSUBS 0.014642f
C1025 VDD1.n101 VSUBS 0.013828f
C1026 VDD1.n102 VSUBS 0.025734f
C1027 VDD1.n103 VSUBS 0.025734f
C1028 VDD1.n104 VSUBS 0.013828f
C1029 VDD1.n105 VSUBS 0.014642f
C1030 VDD1.n106 VSUBS 0.032685f
C1031 VDD1.n107 VSUBS 0.032685f
C1032 VDD1.n108 VSUBS 0.014642f
C1033 VDD1.n109 VSUBS 0.013828f
C1034 VDD1.n110 VSUBS 0.025734f
C1035 VDD1.n111 VSUBS 0.025734f
C1036 VDD1.n112 VSUBS 0.013828f
C1037 VDD1.n113 VSUBS 0.014642f
C1038 VDD1.n114 VSUBS 0.032685f
C1039 VDD1.n115 VSUBS 0.032685f
C1040 VDD1.n116 VSUBS 0.014642f
C1041 VDD1.n117 VSUBS 0.013828f
C1042 VDD1.n118 VSUBS 0.025734f
C1043 VDD1.n119 VSUBS 0.025734f
C1044 VDD1.n120 VSUBS 0.013828f
C1045 VDD1.n121 VSUBS 0.014642f
C1046 VDD1.n122 VSUBS 0.032685f
C1047 VDD1.n123 VSUBS 0.032685f
C1048 VDD1.n124 VSUBS 0.014642f
C1049 VDD1.n125 VSUBS 0.013828f
C1050 VDD1.n126 VSUBS 0.025734f
C1051 VDD1.n127 VSUBS 0.025734f
C1052 VDD1.n128 VSUBS 0.013828f
C1053 VDD1.n129 VSUBS 0.014642f
C1054 VDD1.n130 VSUBS 0.032685f
C1055 VDD1.n131 VSUBS 0.032685f
C1056 VDD1.n132 VSUBS 0.014642f
C1057 VDD1.n133 VSUBS 0.013828f
C1058 VDD1.n134 VSUBS 0.025734f
C1059 VDD1.n135 VSUBS 0.025734f
C1060 VDD1.n136 VSUBS 0.013828f
C1061 VDD1.n137 VSUBS 0.014642f
C1062 VDD1.n138 VSUBS 0.032685f
C1063 VDD1.n139 VSUBS 0.083091f
C1064 VDD1.n140 VSUBS 0.014642f
C1065 VDD1.n141 VSUBS 0.027155f
C1066 VDD1.n142 VSUBS 0.067568f
C1067 VDD1.n143 VSUBS 0.085557f
C1068 VDD1.t1 VSUBS 0.273106f
C1069 VDD1.t4 VSUBS 0.273106f
C1070 VDD1.n144 VSUBS 2.1967f
C1071 VDD1.n145 VSUBS 0.731918f
C1072 VDD1.t3 VSUBS 0.273106f
C1073 VDD1.t5 VSUBS 0.273106f
C1074 VDD1.n146 VSUBS 2.20343f
C1075 VDD1.n147 VSUBS 2.56064f
C1076 VDD1.t8 VSUBS 0.273106f
C1077 VDD1.t2 VSUBS 0.273106f
C1078 VDD1.n148 VSUBS 2.1967f
C1079 VDD1.n149 VSUBS 2.95788f
C1080 VTAIL.t4 VSUBS 0.297773f
C1081 VTAIL.t2 VSUBS 0.297773f
C1082 VTAIL.n0 VSUBS 2.25432f
C1083 VTAIL.n1 VSUBS 0.790575f
C1084 VTAIL.n2 VSUBS 0.031363f
C1085 VTAIL.n3 VSUBS 0.028058f
C1086 VTAIL.n4 VSUBS 0.015077f
C1087 VTAIL.n5 VSUBS 0.035637f
C1088 VTAIL.n6 VSUBS 0.015964f
C1089 VTAIL.n7 VSUBS 0.028058f
C1090 VTAIL.n8 VSUBS 0.015077f
C1091 VTAIL.n9 VSUBS 0.035637f
C1092 VTAIL.n10 VSUBS 0.015964f
C1093 VTAIL.n11 VSUBS 0.028058f
C1094 VTAIL.n12 VSUBS 0.015077f
C1095 VTAIL.n13 VSUBS 0.035637f
C1096 VTAIL.n14 VSUBS 0.015964f
C1097 VTAIL.n15 VSUBS 0.028058f
C1098 VTAIL.n16 VSUBS 0.015077f
C1099 VTAIL.n17 VSUBS 0.035637f
C1100 VTAIL.n18 VSUBS 0.015964f
C1101 VTAIL.n19 VSUBS 0.028058f
C1102 VTAIL.n20 VSUBS 0.015077f
C1103 VTAIL.n21 VSUBS 0.035637f
C1104 VTAIL.n22 VSUBS 0.015964f
C1105 VTAIL.n23 VSUBS 1.59157f
C1106 VTAIL.n24 VSUBS 0.015077f
C1107 VTAIL.t13 VSUBS 0.076183f
C1108 VTAIL.n25 VSUBS 0.184793f
C1109 VTAIL.n26 VSUBS 0.02267f
C1110 VTAIL.n27 VSUBS 0.026728f
C1111 VTAIL.n28 VSUBS 0.035637f
C1112 VTAIL.n29 VSUBS 0.015964f
C1113 VTAIL.n30 VSUBS 0.015077f
C1114 VTAIL.n31 VSUBS 0.028058f
C1115 VTAIL.n32 VSUBS 0.028058f
C1116 VTAIL.n33 VSUBS 0.015077f
C1117 VTAIL.n34 VSUBS 0.015964f
C1118 VTAIL.n35 VSUBS 0.035637f
C1119 VTAIL.n36 VSUBS 0.035637f
C1120 VTAIL.n37 VSUBS 0.015964f
C1121 VTAIL.n38 VSUBS 0.015077f
C1122 VTAIL.n39 VSUBS 0.028058f
C1123 VTAIL.n40 VSUBS 0.028058f
C1124 VTAIL.n41 VSUBS 0.015077f
C1125 VTAIL.n42 VSUBS 0.015964f
C1126 VTAIL.n43 VSUBS 0.035637f
C1127 VTAIL.n44 VSUBS 0.035637f
C1128 VTAIL.n45 VSUBS 0.015964f
C1129 VTAIL.n46 VSUBS 0.015077f
C1130 VTAIL.n47 VSUBS 0.028058f
C1131 VTAIL.n48 VSUBS 0.028058f
C1132 VTAIL.n49 VSUBS 0.015077f
C1133 VTAIL.n50 VSUBS 0.015964f
C1134 VTAIL.n51 VSUBS 0.035637f
C1135 VTAIL.n52 VSUBS 0.035637f
C1136 VTAIL.n53 VSUBS 0.015964f
C1137 VTAIL.n54 VSUBS 0.015077f
C1138 VTAIL.n55 VSUBS 0.028058f
C1139 VTAIL.n56 VSUBS 0.028058f
C1140 VTAIL.n57 VSUBS 0.015077f
C1141 VTAIL.n58 VSUBS 0.015964f
C1142 VTAIL.n59 VSUBS 0.035637f
C1143 VTAIL.n60 VSUBS 0.035637f
C1144 VTAIL.n61 VSUBS 0.015964f
C1145 VTAIL.n62 VSUBS 0.015077f
C1146 VTAIL.n63 VSUBS 0.028058f
C1147 VTAIL.n64 VSUBS 0.028058f
C1148 VTAIL.n65 VSUBS 0.015077f
C1149 VTAIL.n66 VSUBS 0.015964f
C1150 VTAIL.n67 VSUBS 0.035637f
C1151 VTAIL.n68 VSUBS 0.090596f
C1152 VTAIL.n69 VSUBS 0.015964f
C1153 VTAIL.n70 VSUBS 0.029608f
C1154 VTAIL.n71 VSUBS 0.07367f
C1155 VTAIL.n72 VSUBS 0.070504f
C1156 VTAIL.n73 VSUBS 0.228088f
C1157 VTAIL.t11 VSUBS 0.297773f
C1158 VTAIL.t10 VSUBS 0.297773f
C1159 VTAIL.n74 VSUBS 2.25432f
C1160 VTAIL.n75 VSUBS 0.821166f
C1161 VTAIL.t16 VSUBS 0.297773f
C1162 VTAIL.t19 VSUBS 0.297773f
C1163 VTAIL.n76 VSUBS 2.25432f
C1164 VTAIL.n77 VSUBS 2.35345f
C1165 VTAIL.t1 VSUBS 0.297773f
C1166 VTAIL.t7 VSUBS 0.297773f
C1167 VTAIL.n78 VSUBS 2.25434f
C1168 VTAIL.n79 VSUBS 2.35344f
C1169 VTAIL.t3 VSUBS 0.297773f
C1170 VTAIL.t6 VSUBS 0.297773f
C1171 VTAIL.n80 VSUBS 2.25434f
C1172 VTAIL.n81 VSUBS 0.821151f
C1173 VTAIL.n82 VSUBS 0.031363f
C1174 VTAIL.n83 VSUBS 0.028058f
C1175 VTAIL.n84 VSUBS 0.015077f
C1176 VTAIL.n85 VSUBS 0.035637f
C1177 VTAIL.n86 VSUBS 0.015964f
C1178 VTAIL.n87 VSUBS 0.028058f
C1179 VTAIL.n88 VSUBS 0.015077f
C1180 VTAIL.n89 VSUBS 0.035637f
C1181 VTAIL.n90 VSUBS 0.015964f
C1182 VTAIL.n91 VSUBS 0.028058f
C1183 VTAIL.n92 VSUBS 0.015077f
C1184 VTAIL.n93 VSUBS 0.035637f
C1185 VTAIL.n94 VSUBS 0.015964f
C1186 VTAIL.n95 VSUBS 0.028058f
C1187 VTAIL.n96 VSUBS 0.015077f
C1188 VTAIL.n97 VSUBS 0.035637f
C1189 VTAIL.n98 VSUBS 0.015964f
C1190 VTAIL.n99 VSUBS 0.028058f
C1191 VTAIL.n100 VSUBS 0.015077f
C1192 VTAIL.n101 VSUBS 0.035637f
C1193 VTAIL.n102 VSUBS 0.015964f
C1194 VTAIL.n103 VSUBS 1.59157f
C1195 VTAIL.n104 VSUBS 0.015077f
C1196 VTAIL.t8 VSUBS 0.076183f
C1197 VTAIL.n105 VSUBS 0.184793f
C1198 VTAIL.n106 VSUBS 0.02267f
C1199 VTAIL.n107 VSUBS 0.026728f
C1200 VTAIL.n108 VSUBS 0.035637f
C1201 VTAIL.n109 VSUBS 0.015964f
C1202 VTAIL.n110 VSUBS 0.015077f
C1203 VTAIL.n111 VSUBS 0.028058f
C1204 VTAIL.n112 VSUBS 0.028058f
C1205 VTAIL.n113 VSUBS 0.015077f
C1206 VTAIL.n114 VSUBS 0.015964f
C1207 VTAIL.n115 VSUBS 0.035637f
C1208 VTAIL.n116 VSUBS 0.035637f
C1209 VTAIL.n117 VSUBS 0.015964f
C1210 VTAIL.n118 VSUBS 0.015077f
C1211 VTAIL.n119 VSUBS 0.028058f
C1212 VTAIL.n120 VSUBS 0.028058f
C1213 VTAIL.n121 VSUBS 0.015077f
C1214 VTAIL.n122 VSUBS 0.015964f
C1215 VTAIL.n123 VSUBS 0.035637f
C1216 VTAIL.n124 VSUBS 0.035637f
C1217 VTAIL.n125 VSUBS 0.015964f
C1218 VTAIL.n126 VSUBS 0.015077f
C1219 VTAIL.n127 VSUBS 0.028058f
C1220 VTAIL.n128 VSUBS 0.028058f
C1221 VTAIL.n129 VSUBS 0.015077f
C1222 VTAIL.n130 VSUBS 0.015964f
C1223 VTAIL.n131 VSUBS 0.035637f
C1224 VTAIL.n132 VSUBS 0.035637f
C1225 VTAIL.n133 VSUBS 0.015964f
C1226 VTAIL.n134 VSUBS 0.015077f
C1227 VTAIL.n135 VSUBS 0.028058f
C1228 VTAIL.n136 VSUBS 0.028058f
C1229 VTAIL.n137 VSUBS 0.015077f
C1230 VTAIL.n138 VSUBS 0.015964f
C1231 VTAIL.n139 VSUBS 0.035637f
C1232 VTAIL.n140 VSUBS 0.035637f
C1233 VTAIL.n141 VSUBS 0.015964f
C1234 VTAIL.n142 VSUBS 0.015077f
C1235 VTAIL.n143 VSUBS 0.028058f
C1236 VTAIL.n144 VSUBS 0.028058f
C1237 VTAIL.n145 VSUBS 0.015077f
C1238 VTAIL.n146 VSUBS 0.015964f
C1239 VTAIL.n147 VSUBS 0.035637f
C1240 VTAIL.n148 VSUBS 0.090596f
C1241 VTAIL.n149 VSUBS 0.015964f
C1242 VTAIL.n150 VSUBS 0.029608f
C1243 VTAIL.n151 VSUBS 0.07367f
C1244 VTAIL.n152 VSUBS 0.070504f
C1245 VTAIL.n153 VSUBS 0.228088f
C1246 VTAIL.t18 VSUBS 0.297773f
C1247 VTAIL.t15 VSUBS 0.297773f
C1248 VTAIL.n154 VSUBS 2.25434f
C1249 VTAIL.n155 VSUBS 0.811408f
C1250 VTAIL.t14 VSUBS 0.297773f
C1251 VTAIL.t17 VSUBS 0.297773f
C1252 VTAIL.n156 VSUBS 2.25434f
C1253 VTAIL.n157 VSUBS 0.821151f
C1254 VTAIL.n158 VSUBS 0.031363f
C1255 VTAIL.n159 VSUBS 0.028058f
C1256 VTAIL.n160 VSUBS 0.015077f
C1257 VTAIL.n161 VSUBS 0.035637f
C1258 VTAIL.n162 VSUBS 0.015964f
C1259 VTAIL.n163 VSUBS 0.028058f
C1260 VTAIL.n164 VSUBS 0.015077f
C1261 VTAIL.n165 VSUBS 0.035637f
C1262 VTAIL.n166 VSUBS 0.015964f
C1263 VTAIL.n167 VSUBS 0.028058f
C1264 VTAIL.n168 VSUBS 0.015077f
C1265 VTAIL.n169 VSUBS 0.035637f
C1266 VTAIL.n170 VSUBS 0.015964f
C1267 VTAIL.n171 VSUBS 0.028058f
C1268 VTAIL.n172 VSUBS 0.015077f
C1269 VTAIL.n173 VSUBS 0.035637f
C1270 VTAIL.n174 VSUBS 0.015964f
C1271 VTAIL.n175 VSUBS 0.028058f
C1272 VTAIL.n176 VSUBS 0.015077f
C1273 VTAIL.n177 VSUBS 0.035637f
C1274 VTAIL.n178 VSUBS 0.015964f
C1275 VTAIL.n179 VSUBS 1.59157f
C1276 VTAIL.n180 VSUBS 0.015077f
C1277 VTAIL.t12 VSUBS 0.076183f
C1278 VTAIL.n181 VSUBS 0.184793f
C1279 VTAIL.n182 VSUBS 0.02267f
C1280 VTAIL.n183 VSUBS 0.026728f
C1281 VTAIL.n184 VSUBS 0.035637f
C1282 VTAIL.n185 VSUBS 0.015964f
C1283 VTAIL.n186 VSUBS 0.015077f
C1284 VTAIL.n187 VSUBS 0.028058f
C1285 VTAIL.n188 VSUBS 0.028058f
C1286 VTAIL.n189 VSUBS 0.015077f
C1287 VTAIL.n190 VSUBS 0.015964f
C1288 VTAIL.n191 VSUBS 0.035637f
C1289 VTAIL.n192 VSUBS 0.035637f
C1290 VTAIL.n193 VSUBS 0.015964f
C1291 VTAIL.n194 VSUBS 0.015077f
C1292 VTAIL.n195 VSUBS 0.028058f
C1293 VTAIL.n196 VSUBS 0.028058f
C1294 VTAIL.n197 VSUBS 0.015077f
C1295 VTAIL.n198 VSUBS 0.015964f
C1296 VTAIL.n199 VSUBS 0.035637f
C1297 VTAIL.n200 VSUBS 0.035637f
C1298 VTAIL.n201 VSUBS 0.015964f
C1299 VTAIL.n202 VSUBS 0.015077f
C1300 VTAIL.n203 VSUBS 0.028058f
C1301 VTAIL.n204 VSUBS 0.028058f
C1302 VTAIL.n205 VSUBS 0.015077f
C1303 VTAIL.n206 VSUBS 0.015964f
C1304 VTAIL.n207 VSUBS 0.035637f
C1305 VTAIL.n208 VSUBS 0.035637f
C1306 VTAIL.n209 VSUBS 0.015964f
C1307 VTAIL.n210 VSUBS 0.015077f
C1308 VTAIL.n211 VSUBS 0.028058f
C1309 VTAIL.n212 VSUBS 0.028058f
C1310 VTAIL.n213 VSUBS 0.015077f
C1311 VTAIL.n214 VSUBS 0.015964f
C1312 VTAIL.n215 VSUBS 0.035637f
C1313 VTAIL.n216 VSUBS 0.035637f
C1314 VTAIL.n217 VSUBS 0.015964f
C1315 VTAIL.n218 VSUBS 0.015077f
C1316 VTAIL.n219 VSUBS 0.028058f
C1317 VTAIL.n220 VSUBS 0.028058f
C1318 VTAIL.n221 VSUBS 0.015077f
C1319 VTAIL.n222 VSUBS 0.015964f
C1320 VTAIL.n223 VSUBS 0.035637f
C1321 VTAIL.n224 VSUBS 0.090596f
C1322 VTAIL.n225 VSUBS 0.015964f
C1323 VTAIL.n226 VSUBS 0.029608f
C1324 VTAIL.n227 VSUBS 0.07367f
C1325 VTAIL.n228 VSUBS 0.070504f
C1326 VTAIL.n229 VSUBS 1.66568f
C1327 VTAIL.n230 VSUBS 0.031363f
C1328 VTAIL.n231 VSUBS 0.028058f
C1329 VTAIL.n232 VSUBS 0.015077f
C1330 VTAIL.n233 VSUBS 0.035637f
C1331 VTAIL.n234 VSUBS 0.015964f
C1332 VTAIL.n235 VSUBS 0.028058f
C1333 VTAIL.n236 VSUBS 0.015077f
C1334 VTAIL.n237 VSUBS 0.035637f
C1335 VTAIL.n238 VSUBS 0.015964f
C1336 VTAIL.n239 VSUBS 0.028058f
C1337 VTAIL.n240 VSUBS 0.015077f
C1338 VTAIL.n241 VSUBS 0.035637f
C1339 VTAIL.n242 VSUBS 0.015964f
C1340 VTAIL.n243 VSUBS 0.028058f
C1341 VTAIL.n244 VSUBS 0.015077f
C1342 VTAIL.n245 VSUBS 0.035637f
C1343 VTAIL.n246 VSUBS 0.015964f
C1344 VTAIL.n247 VSUBS 0.028058f
C1345 VTAIL.n248 VSUBS 0.015077f
C1346 VTAIL.n249 VSUBS 0.035637f
C1347 VTAIL.n250 VSUBS 0.015964f
C1348 VTAIL.n251 VSUBS 1.59157f
C1349 VTAIL.n252 VSUBS 0.015077f
C1350 VTAIL.t0 VSUBS 0.076183f
C1351 VTAIL.n253 VSUBS 0.184793f
C1352 VTAIL.n254 VSUBS 0.02267f
C1353 VTAIL.n255 VSUBS 0.026728f
C1354 VTAIL.n256 VSUBS 0.035637f
C1355 VTAIL.n257 VSUBS 0.015964f
C1356 VTAIL.n258 VSUBS 0.015077f
C1357 VTAIL.n259 VSUBS 0.028058f
C1358 VTAIL.n260 VSUBS 0.028058f
C1359 VTAIL.n261 VSUBS 0.015077f
C1360 VTAIL.n262 VSUBS 0.015964f
C1361 VTAIL.n263 VSUBS 0.035637f
C1362 VTAIL.n264 VSUBS 0.035637f
C1363 VTAIL.n265 VSUBS 0.015964f
C1364 VTAIL.n266 VSUBS 0.015077f
C1365 VTAIL.n267 VSUBS 0.028058f
C1366 VTAIL.n268 VSUBS 0.028058f
C1367 VTAIL.n269 VSUBS 0.015077f
C1368 VTAIL.n270 VSUBS 0.015964f
C1369 VTAIL.n271 VSUBS 0.035637f
C1370 VTAIL.n272 VSUBS 0.035637f
C1371 VTAIL.n273 VSUBS 0.015964f
C1372 VTAIL.n274 VSUBS 0.015077f
C1373 VTAIL.n275 VSUBS 0.028058f
C1374 VTAIL.n276 VSUBS 0.028058f
C1375 VTAIL.n277 VSUBS 0.015077f
C1376 VTAIL.n278 VSUBS 0.015964f
C1377 VTAIL.n279 VSUBS 0.035637f
C1378 VTAIL.n280 VSUBS 0.035637f
C1379 VTAIL.n281 VSUBS 0.015964f
C1380 VTAIL.n282 VSUBS 0.015077f
C1381 VTAIL.n283 VSUBS 0.028058f
C1382 VTAIL.n284 VSUBS 0.028058f
C1383 VTAIL.n285 VSUBS 0.015077f
C1384 VTAIL.n286 VSUBS 0.015964f
C1385 VTAIL.n287 VSUBS 0.035637f
C1386 VTAIL.n288 VSUBS 0.035637f
C1387 VTAIL.n289 VSUBS 0.015964f
C1388 VTAIL.n290 VSUBS 0.015077f
C1389 VTAIL.n291 VSUBS 0.028058f
C1390 VTAIL.n292 VSUBS 0.028058f
C1391 VTAIL.n293 VSUBS 0.015077f
C1392 VTAIL.n294 VSUBS 0.015964f
C1393 VTAIL.n295 VSUBS 0.035637f
C1394 VTAIL.n296 VSUBS 0.090596f
C1395 VTAIL.n297 VSUBS 0.015964f
C1396 VTAIL.n298 VSUBS 0.029608f
C1397 VTAIL.n299 VSUBS 0.07367f
C1398 VTAIL.n300 VSUBS 0.070504f
C1399 VTAIL.n301 VSUBS 1.66568f
C1400 VTAIL.t5 VSUBS 0.297773f
C1401 VTAIL.t9 VSUBS 0.297773f
C1402 VTAIL.n302 VSUBS 2.25432f
C1403 VTAIL.n303 VSUBS 0.737576f
C1404 VP.n0 VSUBS 0.060231f
C1405 VP.t6 VSUBS 1.67328f
C1406 VP.n1 VSUBS 0.040342f
C1407 VP.n2 VSUBS 0.045138f
C1408 VP.t5 VSUBS 1.67328f
C1409 VP.n3 VSUBS 0.056982f
C1410 VP.n4 VSUBS 0.060231f
C1411 VP.t7 VSUBS 1.74312f
C1412 VP.t1 VSUBS 1.67328f
C1413 VP.n5 VSUBS 0.040342f
C1414 VP.n6 VSUBS 0.045138f
C1415 VP.t9 VSUBS 1.67328f
C1416 VP.n7 VSUBS 0.056982f
C1417 VP.t2 VSUBS 1.67328f
C1418 VP.n8 VSUBS 0.64806f
C1419 VP.t0 VSUBS 1.76958f
C1420 VP.n9 VSUBS 0.681181f
C1421 VP.n10 VSUBS 0.189929f
C1422 VP.n11 VSUBS 0.045138f
C1423 VP.n12 VSUBS 0.040342f
C1424 VP.n13 VSUBS 0.063765f
C1425 VP.n14 VSUBS 0.613488f
C1426 VP.n15 VSUBS 0.063765f
C1427 VP.n16 VSUBS 0.045138f
C1428 VP.n17 VSUBS 0.045138f
C1429 VP.n18 VSUBS 0.045138f
C1430 VP.n19 VSUBS 0.056982f
C1431 VP.n20 VSUBS 0.613488f
C1432 VP.n21 VSUBS 0.058577f
C1433 VP.n22 VSUBS 0.68271f
C1434 VP.n23 VSUBS 2.1542f
C1435 VP.n24 VSUBS 2.18968f
C1436 VP.t3 VSUBS 1.74312f
C1437 VP.n25 VSUBS 0.68271f
C1438 VP.t8 VSUBS 1.67328f
C1439 VP.n26 VSUBS 0.613488f
C1440 VP.n27 VSUBS 0.058577f
C1441 VP.n28 VSUBS 0.060231f
C1442 VP.n29 VSUBS 0.045138f
C1443 VP.n30 VSUBS 0.045138f
C1444 VP.n31 VSUBS 0.040342f
C1445 VP.n32 VSUBS 0.063765f
C1446 VP.n33 VSUBS 0.613488f
C1447 VP.n34 VSUBS 0.063765f
C1448 VP.n35 VSUBS 0.045138f
C1449 VP.n36 VSUBS 0.045138f
C1450 VP.n37 VSUBS 0.045138f
C1451 VP.n38 VSUBS 0.056982f
C1452 VP.n39 VSUBS 0.613488f
C1453 VP.n40 VSUBS 0.058577f
C1454 VP.t4 VSUBS 1.74312f
C1455 VP.n41 VSUBS 0.68271f
C1456 VP.n42 VSUBS 0.042274f
.ends

