* NGSPICE file created from diff_pair_sample_0959.ext - technology: sky130A

.subckt diff_pair_sample_0959 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X1 VDD1.t7 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=1.716 ps=9.58 w=4.4 l=1.86
X2 VTAIL.t14 VN.t1 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0.726 ps=4.73 w=4.4 l=1.86
X3 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0 ps=0 w=4.4 l=1.86
X4 VTAIL.t2 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0.726 ps=4.73 w=4.4 l=1.86
X5 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X6 VTAIL.t13 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0.726 ps=4.73 w=4.4 l=1.86
X7 VTAIL.t7 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X8 VDD2.t7 VN.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X9 VTAIL.t5 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0.726 ps=4.73 w=4.4 l=1.86
X10 VDD2.t6 VN.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=1.716 ps=9.58 w=4.4 l=1.86
X11 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0 ps=0 w=4.4 l=1.86
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0 ps=0 w=4.4 l=1.86
X13 VDD2.t5 VN.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=1.716 ps=9.58 w=4.4 l=1.86
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.716 pd=9.58 as=0 ps=0 w=4.4 l=1.86
X15 VDD1.t2 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X16 VDD2.t2 VN.t6 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X17 VTAIL.t8 VN.t7 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
X18 VDD1.t1 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=1.716 ps=9.58 w=4.4 l=1.86
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.726 pd=4.73 as=0.726 ps=4.73 w=4.4 l=1.86
R0 VN.n22 VN.n21 184.171
R1 VN.n45 VN.n44 184.171
R2 VN.n43 VN.n23 161.3
R3 VN.n42 VN.n41 161.3
R4 VN.n40 VN.n24 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n25 161.3
R7 VN.n35 VN.n34 161.3
R8 VN.n33 VN.n26 161.3
R9 VN.n32 VN.n31 161.3
R10 VN.n30 VN.n27 161.3
R11 VN.n20 VN.n0 161.3
R12 VN.n19 VN.n18 161.3
R13 VN.n17 VN.n1 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n14 VN.n2 161.3
R16 VN.n12 VN.n11 161.3
R17 VN.n10 VN.n3 161.3
R18 VN.n9 VN.n8 161.3
R19 VN.n7 VN.n4 161.3
R20 VN.n5 VN.t1 89.9794
R21 VN.n28 VN.t5 89.9794
R22 VN.n6 VN.t3 57.0113
R23 VN.n13 VN.t7 57.0113
R24 VN.n21 VN.t4 57.0113
R25 VN.n29 VN.t0 57.0113
R26 VN.n36 VN.t6 57.0113
R27 VN.n44 VN.t2 57.0113
R28 VN.n8 VN.n3 56.5617
R29 VN.n31 VN.n26 56.5617
R30 VN.n6 VN.n5 53.0172
R31 VN.n29 VN.n28 53.0172
R32 VN.n15 VN.n1 46.3896
R33 VN.n38 VN.n24 46.3896
R34 VN VN.n45 41.9418
R35 VN.n19 VN.n1 34.7644
R36 VN.n42 VN.n24 34.7644
R37 VN.n8 VN.n7 24.5923
R38 VN.n12 VN.n3 24.5923
R39 VN.n15 VN.n14 24.5923
R40 VN.n20 VN.n19 24.5923
R41 VN.n31 VN.n30 24.5923
R42 VN.n38 VN.n37 24.5923
R43 VN.n35 VN.n26 24.5923
R44 VN.n43 VN.n42 24.5923
R45 VN.n7 VN.n6 16.9689
R46 VN.n13 VN.n12 16.9689
R47 VN.n30 VN.n29 16.9689
R48 VN.n36 VN.n35 16.9689
R49 VN.n28 VN.n27 12.4356
R50 VN.n5 VN.n4 12.4356
R51 VN.n14 VN.n13 7.62397
R52 VN.n37 VN.n36 7.62397
R53 VN.n21 VN.n20 1.72193
R54 VN.n44 VN.n43 1.72193
R55 VN.n45 VN.n23 0.189894
R56 VN.n41 VN.n23 0.189894
R57 VN.n41 VN.n40 0.189894
R58 VN.n40 VN.n39 0.189894
R59 VN.n39 VN.n25 0.189894
R60 VN.n34 VN.n25 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n32 0.189894
R63 VN.n32 VN.n27 0.189894
R64 VN.n9 VN.n4 0.189894
R65 VN.n10 VN.n9 0.189894
R66 VN.n11 VN.n10 0.189894
R67 VN.n11 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n18 VN.n17 0.189894
R71 VN.n18 VN.n0 0.189894
R72 VN.n22 VN.n0 0.189894
R73 VN VN.n22 0.0516364
R74 VDD2.n2 VDD2.n1 76.6856
R75 VDD2.n2 VDD2.n0 76.6856
R76 VDD2 VDD2.n5 76.6829
R77 VDD2.n4 VDD2.n3 75.7972
R78 VDD2.n4 VDD2.n2 36.0041
R79 VDD2.n5 VDD2.t4 4.5005
R80 VDD2.n5 VDD2.t5 4.5005
R81 VDD2.n3 VDD2.t1 4.5005
R82 VDD2.n3 VDD2.t2 4.5005
R83 VDD2.n1 VDD2.t3 4.5005
R84 VDD2.n1 VDD2.t6 4.5005
R85 VDD2.n0 VDD2.t0 4.5005
R86 VDD2.n0 VDD2.t7 4.5005
R87 VDD2 VDD2.n4 1.00266
R88 VTAIL.n11 VTAIL.t5 63.6184
R89 VTAIL.n10 VTAIL.t10 63.6184
R90 VTAIL.n7 VTAIL.t13 63.6184
R91 VTAIL.n15 VTAIL.t11 63.6182
R92 VTAIL.n2 VTAIL.t14 63.6182
R93 VTAIL.n3 VTAIL.t3 63.6182
R94 VTAIL.n6 VTAIL.t2 63.6182
R95 VTAIL.n14 VTAIL.t6 63.6182
R96 VTAIL.n13 VTAIL.n12 59.1184
R97 VTAIL.n9 VTAIL.n8 59.1184
R98 VTAIL.n1 VTAIL.n0 59.1182
R99 VTAIL.n5 VTAIL.n4 59.1182
R100 VTAIL.n15 VTAIL.n14 18.0479
R101 VTAIL.n7 VTAIL.n6 18.0479
R102 VTAIL.n0 VTAIL.t12 4.5005
R103 VTAIL.n0 VTAIL.t8 4.5005
R104 VTAIL.n4 VTAIL.t0 4.5005
R105 VTAIL.n4 VTAIL.t7 4.5005
R106 VTAIL.n12 VTAIL.t4 4.5005
R107 VTAIL.n12 VTAIL.t1 4.5005
R108 VTAIL.n8 VTAIL.t9 4.5005
R109 VTAIL.n8 VTAIL.t15 4.5005
R110 VTAIL.n9 VTAIL.n7 1.88843
R111 VTAIL.n10 VTAIL.n9 1.88843
R112 VTAIL.n13 VTAIL.n11 1.88843
R113 VTAIL.n14 VTAIL.n13 1.88843
R114 VTAIL.n6 VTAIL.n5 1.88843
R115 VTAIL.n5 VTAIL.n3 1.88843
R116 VTAIL.n2 VTAIL.n1 1.88843
R117 VTAIL VTAIL.n15 1.83024
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 B.n575 B.n574 585
R122 B.n197 B.n100 585
R123 B.n196 B.n195 585
R124 B.n194 B.n193 585
R125 B.n192 B.n191 585
R126 B.n190 B.n189 585
R127 B.n188 B.n187 585
R128 B.n186 B.n185 585
R129 B.n184 B.n183 585
R130 B.n182 B.n181 585
R131 B.n180 B.n179 585
R132 B.n178 B.n177 585
R133 B.n176 B.n175 585
R134 B.n174 B.n173 585
R135 B.n172 B.n171 585
R136 B.n170 B.n169 585
R137 B.n168 B.n167 585
R138 B.n166 B.n165 585
R139 B.n164 B.n163 585
R140 B.n161 B.n160 585
R141 B.n159 B.n158 585
R142 B.n157 B.n156 585
R143 B.n155 B.n154 585
R144 B.n153 B.n152 585
R145 B.n151 B.n150 585
R146 B.n149 B.n148 585
R147 B.n147 B.n146 585
R148 B.n145 B.n144 585
R149 B.n143 B.n142 585
R150 B.n140 B.n139 585
R151 B.n138 B.n137 585
R152 B.n136 B.n135 585
R153 B.n134 B.n133 585
R154 B.n132 B.n131 585
R155 B.n130 B.n129 585
R156 B.n128 B.n127 585
R157 B.n126 B.n125 585
R158 B.n124 B.n123 585
R159 B.n122 B.n121 585
R160 B.n120 B.n119 585
R161 B.n118 B.n117 585
R162 B.n116 B.n115 585
R163 B.n114 B.n113 585
R164 B.n112 B.n111 585
R165 B.n110 B.n109 585
R166 B.n108 B.n107 585
R167 B.n106 B.n105 585
R168 B.n75 B.n74 585
R169 B.n573 B.n76 585
R170 B.n578 B.n76 585
R171 B.n572 B.n571 585
R172 B.n571 B.n72 585
R173 B.n570 B.n71 585
R174 B.n584 B.n71 585
R175 B.n569 B.n70 585
R176 B.n585 B.n70 585
R177 B.n568 B.n69 585
R178 B.n586 B.n69 585
R179 B.n567 B.n566 585
R180 B.n566 B.n65 585
R181 B.n565 B.n64 585
R182 B.n592 B.n64 585
R183 B.n564 B.n63 585
R184 B.n593 B.n63 585
R185 B.n563 B.n62 585
R186 B.n594 B.n62 585
R187 B.n562 B.n561 585
R188 B.n561 B.n58 585
R189 B.n560 B.n57 585
R190 B.n600 B.n57 585
R191 B.n559 B.n56 585
R192 B.n601 B.n56 585
R193 B.n558 B.n55 585
R194 B.n602 B.n55 585
R195 B.n557 B.n556 585
R196 B.n556 B.n51 585
R197 B.n555 B.n50 585
R198 B.n608 B.n50 585
R199 B.n554 B.n49 585
R200 B.n609 B.n49 585
R201 B.n553 B.n48 585
R202 B.n610 B.n48 585
R203 B.n552 B.n551 585
R204 B.n551 B.n44 585
R205 B.n550 B.n43 585
R206 B.n616 B.n43 585
R207 B.n549 B.n42 585
R208 B.n617 B.n42 585
R209 B.n548 B.n41 585
R210 B.n618 B.n41 585
R211 B.n547 B.n546 585
R212 B.n546 B.n37 585
R213 B.n545 B.n36 585
R214 B.n624 B.n36 585
R215 B.n544 B.n35 585
R216 B.n625 B.n35 585
R217 B.n543 B.n34 585
R218 B.n626 B.n34 585
R219 B.n542 B.n541 585
R220 B.n541 B.n30 585
R221 B.n540 B.n29 585
R222 B.n632 B.n29 585
R223 B.n539 B.n28 585
R224 B.n633 B.n28 585
R225 B.n538 B.n27 585
R226 B.n634 B.n27 585
R227 B.n537 B.n536 585
R228 B.n536 B.n26 585
R229 B.n535 B.n22 585
R230 B.n640 B.n22 585
R231 B.n534 B.n21 585
R232 B.n641 B.n21 585
R233 B.n533 B.n20 585
R234 B.n642 B.n20 585
R235 B.n532 B.n531 585
R236 B.n531 B.n16 585
R237 B.n530 B.n15 585
R238 B.n648 B.n15 585
R239 B.n529 B.n14 585
R240 B.n649 B.n14 585
R241 B.n528 B.n13 585
R242 B.n650 B.n13 585
R243 B.n527 B.n526 585
R244 B.n526 B.n12 585
R245 B.n525 B.n524 585
R246 B.n525 B.n8 585
R247 B.n523 B.n7 585
R248 B.n657 B.n7 585
R249 B.n522 B.n6 585
R250 B.n658 B.n6 585
R251 B.n521 B.n5 585
R252 B.n659 B.n5 585
R253 B.n520 B.n519 585
R254 B.n519 B.n4 585
R255 B.n518 B.n198 585
R256 B.n518 B.n517 585
R257 B.n508 B.n199 585
R258 B.n200 B.n199 585
R259 B.n510 B.n509 585
R260 B.n511 B.n510 585
R261 B.n507 B.n204 585
R262 B.n208 B.n204 585
R263 B.n506 B.n505 585
R264 B.n505 B.n504 585
R265 B.n206 B.n205 585
R266 B.n207 B.n206 585
R267 B.n497 B.n496 585
R268 B.n498 B.n497 585
R269 B.n495 B.n213 585
R270 B.n213 B.n212 585
R271 B.n494 B.n493 585
R272 B.n493 B.n492 585
R273 B.n215 B.n214 585
R274 B.n485 B.n215 585
R275 B.n484 B.n483 585
R276 B.n486 B.n484 585
R277 B.n482 B.n220 585
R278 B.n220 B.n219 585
R279 B.n481 B.n480 585
R280 B.n480 B.n479 585
R281 B.n222 B.n221 585
R282 B.n223 B.n222 585
R283 B.n472 B.n471 585
R284 B.n473 B.n472 585
R285 B.n470 B.n228 585
R286 B.n228 B.n227 585
R287 B.n469 B.n468 585
R288 B.n468 B.n467 585
R289 B.n230 B.n229 585
R290 B.n231 B.n230 585
R291 B.n460 B.n459 585
R292 B.n461 B.n460 585
R293 B.n458 B.n236 585
R294 B.n236 B.n235 585
R295 B.n457 B.n456 585
R296 B.n456 B.n455 585
R297 B.n238 B.n237 585
R298 B.n239 B.n238 585
R299 B.n448 B.n447 585
R300 B.n449 B.n448 585
R301 B.n446 B.n244 585
R302 B.n244 B.n243 585
R303 B.n445 B.n444 585
R304 B.n444 B.n443 585
R305 B.n246 B.n245 585
R306 B.n247 B.n246 585
R307 B.n436 B.n435 585
R308 B.n437 B.n436 585
R309 B.n434 B.n252 585
R310 B.n252 B.n251 585
R311 B.n433 B.n432 585
R312 B.n432 B.n431 585
R313 B.n254 B.n253 585
R314 B.n255 B.n254 585
R315 B.n424 B.n423 585
R316 B.n425 B.n424 585
R317 B.n422 B.n260 585
R318 B.n260 B.n259 585
R319 B.n421 B.n420 585
R320 B.n420 B.n419 585
R321 B.n262 B.n261 585
R322 B.n263 B.n262 585
R323 B.n412 B.n411 585
R324 B.n413 B.n412 585
R325 B.n410 B.n268 585
R326 B.n268 B.n267 585
R327 B.n409 B.n408 585
R328 B.n408 B.n407 585
R329 B.n270 B.n269 585
R330 B.n271 B.n270 585
R331 B.n400 B.n399 585
R332 B.n401 B.n400 585
R333 B.n274 B.n273 585
R334 B.n307 B.n306 585
R335 B.n308 B.n304 585
R336 B.n304 B.n275 585
R337 B.n310 B.n309 585
R338 B.n312 B.n303 585
R339 B.n315 B.n314 585
R340 B.n316 B.n302 585
R341 B.n318 B.n317 585
R342 B.n320 B.n301 585
R343 B.n323 B.n322 585
R344 B.n324 B.n300 585
R345 B.n326 B.n325 585
R346 B.n328 B.n299 585
R347 B.n331 B.n330 585
R348 B.n332 B.n298 585
R349 B.n334 B.n333 585
R350 B.n336 B.n297 585
R351 B.n339 B.n338 585
R352 B.n340 B.n294 585
R353 B.n343 B.n342 585
R354 B.n345 B.n293 585
R355 B.n348 B.n347 585
R356 B.n349 B.n292 585
R357 B.n351 B.n350 585
R358 B.n353 B.n291 585
R359 B.n356 B.n355 585
R360 B.n357 B.n290 585
R361 B.n359 B.n358 585
R362 B.n361 B.n289 585
R363 B.n364 B.n363 585
R364 B.n365 B.n285 585
R365 B.n367 B.n366 585
R366 B.n369 B.n284 585
R367 B.n372 B.n371 585
R368 B.n373 B.n283 585
R369 B.n375 B.n374 585
R370 B.n377 B.n282 585
R371 B.n380 B.n379 585
R372 B.n381 B.n281 585
R373 B.n383 B.n382 585
R374 B.n385 B.n280 585
R375 B.n388 B.n387 585
R376 B.n389 B.n279 585
R377 B.n391 B.n390 585
R378 B.n393 B.n278 585
R379 B.n394 B.n277 585
R380 B.n397 B.n396 585
R381 B.n398 B.n276 585
R382 B.n276 B.n275 585
R383 B.n403 B.n402 585
R384 B.n402 B.n401 585
R385 B.n404 B.n272 585
R386 B.n272 B.n271 585
R387 B.n406 B.n405 585
R388 B.n407 B.n406 585
R389 B.n266 B.n265 585
R390 B.n267 B.n266 585
R391 B.n415 B.n414 585
R392 B.n414 B.n413 585
R393 B.n416 B.n264 585
R394 B.n264 B.n263 585
R395 B.n418 B.n417 585
R396 B.n419 B.n418 585
R397 B.n258 B.n257 585
R398 B.n259 B.n258 585
R399 B.n427 B.n426 585
R400 B.n426 B.n425 585
R401 B.n428 B.n256 585
R402 B.n256 B.n255 585
R403 B.n430 B.n429 585
R404 B.n431 B.n430 585
R405 B.n250 B.n249 585
R406 B.n251 B.n250 585
R407 B.n439 B.n438 585
R408 B.n438 B.n437 585
R409 B.n440 B.n248 585
R410 B.n248 B.n247 585
R411 B.n442 B.n441 585
R412 B.n443 B.n442 585
R413 B.n242 B.n241 585
R414 B.n243 B.n242 585
R415 B.n451 B.n450 585
R416 B.n450 B.n449 585
R417 B.n452 B.n240 585
R418 B.n240 B.n239 585
R419 B.n454 B.n453 585
R420 B.n455 B.n454 585
R421 B.n234 B.n233 585
R422 B.n235 B.n234 585
R423 B.n463 B.n462 585
R424 B.n462 B.n461 585
R425 B.n464 B.n232 585
R426 B.n232 B.n231 585
R427 B.n466 B.n465 585
R428 B.n467 B.n466 585
R429 B.n226 B.n225 585
R430 B.n227 B.n226 585
R431 B.n475 B.n474 585
R432 B.n474 B.n473 585
R433 B.n476 B.n224 585
R434 B.n224 B.n223 585
R435 B.n478 B.n477 585
R436 B.n479 B.n478 585
R437 B.n218 B.n217 585
R438 B.n219 B.n218 585
R439 B.n488 B.n487 585
R440 B.n487 B.n486 585
R441 B.n489 B.n216 585
R442 B.n485 B.n216 585
R443 B.n491 B.n490 585
R444 B.n492 B.n491 585
R445 B.n211 B.n210 585
R446 B.n212 B.n211 585
R447 B.n500 B.n499 585
R448 B.n499 B.n498 585
R449 B.n501 B.n209 585
R450 B.n209 B.n207 585
R451 B.n503 B.n502 585
R452 B.n504 B.n503 585
R453 B.n203 B.n202 585
R454 B.n208 B.n203 585
R455 B.n513 B.n512 585
R456 B.n512 B.n511 585
R457 B.n514 B.n201 585
R458 B.n201 B.n200 585
R459 B.n516 B.n515 585
R460 B.n517 B.n516 585
R461 B.n3 B.n0 585
R462 B.n4 B.n3 585
R463 B.n656 B.n1 585
R464 B.n657 B.n656 585
R465 B.n655 B.n654 585
R466 B.n655 B.n8 585
R467 B.n653 B.n9 585
R468 B.n12 B.n9 585
R469 B.n652 B.n651 585
R470 B.n651 B.n650 585
R471 B.n11 B.n10 585
R472 B.n649 B.n11 585
R473 B.n647 B.n646 585
R474 B.n648 B.n647 585
R475 B.n645 B.n17 585
R476 B.n17 B.n16 585
R477 B.n644 B.n643 585
R478 B.n643 B.n642 585
R479 B.n19 B.n18 585
R480 B.n641 B.n19 585
R481 B.n639 B.n638 585
R482 B.n640 B.n639 585
R483 B.n637 B.n23 585
R484 B.n26 B.n23 585
R485 B.n636 B.n635 585
R486 B.n635 B.n634 585
R487 B.n25 B.n24 585
R488 B.n633 B.n25 585
R489 B.n631 B.n630 585
R490 B.n632 B.n631 585
R491 B.n629 B.n31 585
R492 B.n31 B.n30 585
R493 B.n628 B.n627 585
R494 B.n627 B.n626 585
R495 B.n33 B.n32 585
R496 B.n625 B.n33 585
R497 B.n623 B.n622 585
R498 B.n624 B.n623 585
R499 B.n621 B.n38 585
R500 B.n38 B.n37 585
R501 B.n620 B.n619 585
R502 B.n619 B.n618 585
R503 B.n40 B.n39 585
R504 B.n617 B.n40 585
R505 B.n615 B.n614 585
R506 B.n616 B.n615 585
R507 B.n613 B.n45 585
R508 B.n45 B.n44 585
R509 B.n612 B.n611 585
R510 B.n611 B.n610 585
R511 B.n47 B.n46 585
R512 B.n609 B.n47 585
R513 B.n607 B.n606 585
R514 B.n608 B.n607 585
R515 B.n605 B.n52 585
R516 B.n52 B.n51 585
R517 B.n604 B.n603 585
R518 B.n603 B.n602 585
R519 B.n54 B.n53 585
R520 B.n601 B.n54 585
R521 B.n599 B.n598 585
R522 B.n600 B.n599 585
R523 B.n597 B.n59 585
R524 B.n59 B.n58 585
R525 B.n596 B.n595 585
R526 B.n595 B.n594 585
R527 B.n61 B.n60 585
R528 B.n593 B.n61 585
R529 B.n591 B.n590 585
R530 B.n592 B.n591 585
R531 B.n589 B.n66 585
R532 B.n66 B.n65 585
R533 B.n588 B.n587 585
R534 B.n587 B.n586 585
R535 B.n68 B.n67 585
R536 B.n585 B.n68 585
R537 B.n583 B.n582 585
R538 B.n584 B.n583 585
R539 B.n581 B.n73 585
R540 B.n73 B.n72 585
R541 B.n580 B.n579 585
R542 B.n579 B.n578 585
R543 B.n660 B.n659 585
R544 B.n658 B.n2 585
R545 B.n579 B.n75 478.086
R546 B.n575 B.n76 478.086
R547 B.n400 B.n276 478.086
R548 B.n402 B.n274 478.086
R549 B.n103 B.t12 263.579
R550 B.n101 B.t16 263.579
R551 B.n286 B.t8 263.579
R552 B.n295 B.t19 263.579
R553 B.n577 B.n576 256.663
R554 B.n577 B.n99 256.663
R555 B.n577 B.n98 256.663
R556 B.n577 B.n97 256.663
R557 B.n577 B.n96 256.663
R558 B.n577 B.n95 256.663
R559 B.n577 B.n94 256.663
R560 B.n577 B.n93 256.663
R561 B.n577 B.n92 256.663
R562 B.n577 B.n91 256.663
R563 B.n577 B.n90 256.663
R564 B.n577 B.n89 256.663
R565 B.n577 B.n88 256.663
R566 B.n577 B.n87 256.663
R567 B.n577 B.n86 256.663
R568 B.n577 B.n85 256.663
R569 B.n577 B.n84 256.663
R570 B.n577 B.n83 256.663
R571 B.n577 B.n82 256.663
R572 B.n577 B.n81 256.663
R573 B.n577 B.n80 256.663
R574 B.n577 B.n79 256.663
R575 B.n577 B.n78 256.663
R576 B.n577 B.n77 256.663
R577 B.n305 B.n275 256.663
R578 B.n311 B.n275 256.663
R579 B.n313 B.n275 256.663
R580 B.n319 B.n275 256.663
R581 B.n321 B.n275 256.663
R582 B.n327 B.n275 256.663
R583 B.n329 B.n275 256.663
R584 B.n335 B.n275 256.663
R585 B.n337 B.n275 256.663
R586 B.n344 B.n275 256.663
R587 B.n346 B.n275 256.663
R588 B.n352 B.n275 256.663
R589 B.n354 B.n275 256.663
R590 B.n360 B.n275 256.663
R591 B.n362 B.n275 256.663
R592 B.n368 B.n275 256.663
R593 B.n370 B.n275 256.663
R594 B.n376 B.n275 256.663
R595 B.n378 B.n275 256.663
R596 B.n384 B.n275 256.663
R597 B.n386 B.n275 256.663
R598 B.n392 B.n275 256.663
R599 B.n395 B.n275 256.663
R600 B.n662 B.n661 256.663
R601 B.n107 B.n106 163.367
R602 B.n111 B.n110 163.367
R603 B.n115 B.n114 163.367
R604 B.n119 B.n118 163.367
R605 B.n123 B.n122 163.367
R606 B.n127 B.n126 163.367
R607 B.n131 B.n130 163.367
R608 B.n135 B.n134 163.367
R609 B.n139 B.n138 163.367
R610 B.n144 B.n143 163.367
R611 B.n148 B.n147 163.367
R612 B.n152 B.n151 163.367
R613 B.n156 B.n155 163.367
R614 B.n160 B.n159 163.367
R615 B.n165 B.n164 163.367
R616 B.n169 B.n168 163.367
R617 B.n173 B.n172 163.367
R618 B.n177 B.n176 163.367
R619 B.n181 B.n180 163.367
R620 B.n185 B.n184 163.367
R621 B.n189 B.n188 163.367
R622 B.n193 B.n192 163.367
R623 B.n195 B.n100 163.367
R624 B.n400 B.n270 163.367
R625 B.n408 B.n270 163.367
R626 B.n408 B.n268 163.367
R627 B.n412 B.n268 163.367
R628 B.n412 B.n262 163.367
R629 B.n420 B.n262 163.367
R630 B.n420 B.n260 163.367
R631 B.n424 B.n260 163.367
R632 B.n424 B.n254 163.367
R633 B.n432 B.n254 163.367
R634 B.n432 B.n252 163.367
R635 B.n436 B.n252 163.367
R636 B.n436 B.n246 163.367
R637 B.n444 B.n246 163.367
R638 B.n444 B.n244 163.367
R639 B.n448 B.n244 163.367
R640 B.n448 B.n238 163.367
R641 B.n456 B.n238 163.367
R642 B.n456 B.n236 163.367
R643 B.n460 B.n236 163.367
R644 B.n460 B.n230 163.367
R645 B.n468 B.n230 163.367
R646 B.n468 B.n228 163.367
R647 B.n472 B.n228 163.367
R648 B.n472 B.n222 163.367
R649 B.n480 B.n222 163.367
R650 B.n480 B.n220 163.367
R651 B.n484 B.n220 163.367
R652 B.n484 B.n215 163.367
R653 B.n493 B.n215 163.367
R654 B.n493 B.n213 163.367
R655 B.n497 B.n213 163.367
R656 B.n497 B.n206 163.367
R657 B.n505 B.n206 163.367
R658 B.n505 B.n204 163.367
R659 B.n510 B.n204 163.367
R660 B.n510 B.n199 163.367
R661 B.n518 B.n199 163.367
R662 B.n519 B.n518 163.367
R663 B.n519 B.n5 163.367
R664 B.n6 B.n5 163.367
R665 B.n7 B.n6 163.367
R666 B.n525 B.n7 163.367
R667 B.n526 B.n525 163.367
R668 B.n526 B.n13 163.367
R669 B.n14 B.n13 163.367
R670 B.n15 B.n14 163.367
R671 B.n531 B.n15 163.367
R672 B.n531 B.n20 163.367
R673 B.n21 B.n20 163.367
R674 B.n22 B.n21 163.367
R675 B.n536 B.n22 163.367
R676 B.n536 B.n27 163.367
R677 B.n28 B.n27 163.367
R678 B.n29 B.n28 163.367
R679 B.n541 B.n29 163.367
R680 B.n541 B.n34 163.367
R681 B.n35 B.n34 163.367
R682 B.n36 B.n35 163.367
R683 B.n546 B.n36 163.367
R684 B.n546 B.n41 163.367
R685 B.n42 B.n41 163.367
R686 B.n43 B.n42 163.367
R687 B.n551 B.n43 163.367
R688 B.n551 B.n48 163.367
R689 B.n49 B.n48 163.367
R690 B.n50 B.n49 163.367
R691 B.n556 B.n50 163.367
R692 B.n556 B.n55 163.367
R693 B.n56 B.n55 163.367
R694 B.n57 B.n56 163.367
R695 B.n561 B.n57 163.367
R696 B.n561 B.n62 163.367
R697 B.n63 B.n62 163.367
R698 B.n64 B.n63 163.367
R699 B.n566 B.n64 163.367
R700 B.n566 B.n69 163.367
R701 B.n70 B.n69 163.367
R702 B.n71 B.n70 163.367
R703 B.n571 B.n71 163.367
R704 B.n571 B.n76 163.367
R705 B.n306 B.n304 163.367
R706 B.n310 B.n304 163.367
R707 B.n314 B.n312 163.367
R708 B.n318 B.n302 163.367
R709 B.n322 B.n320 163.367
R710 B.n326 B.n300 163.367
R711 B.n330 B.n328 163.367
R712 B.n334 B.n298 163.367
R713 B.n338 B.n336 163.367
R714 B.n343 B.n294 163.367
R715 B.n347 B.n345 163.367
R716 B.n351 B.n292 163.367
R717 B.n355 B.n353 163.367
R718 B.n359 B.n290 163.367
R719 B.n363 B.n361 163.367
R720 B.n367 B.n285 163.367
R721 B.n371 B.n369 163.367
R722 B.n375 B.n283 163.367
R723 B.n379 B.n377 163.367
R724 B.n383 B.n281 163.367
R725 B.n387 B.n385 163.367
R726 B.n391 B.n279 163.367
R727 B.n394 B.n393 163.367
R728 B.n396 B.n276 163.367
R729 B.n402 B.n272 163.367
R730 B.n406 B.n272 163.367
R731 B.n406 B.n266 163.367
R732 B.n414 B.n266 163.367
R733 B.n414 B.n264 163.367
R734 B.n418 B.n264 163.367
R735 B.n418 B.n258 163.367
R736 B.n426 B.n258 163.367
R737 B.n426 B.n256 163.367
R738 B.n430 B.n256 163.367
R739 B.n430 B.n250 163.367
R740 B.n438 B.n250 163.367
R741 B.n438 B.n248 163.367
R742 B.n442 B.n248 163.367
R743 B.n442 B.n242 163.367
R744 B.n450 B.n242 163.367
R745 B.n450 B.n240 163.367
R746 B.n454 B.n240 163.367
R747 B.n454 B.n234 163.367
R748 B.n462 B.n234 163.367
R749 B.n462 B.n232 163.367
R750 B.n466 B.n232 163.367
R751 B.n466 B.n226 163.367
R752 B.n474 B.n226 163.367
R753 B.n474 B.n224 163.367
R754 B.n478 B.n224 163.367
R755 B.n478 B.n218 163.367
R756 B.n487 B.n218 163.367
R757 B.n487 B.n216 163.367
R758 B.n491 B.n216 163.367
R759 B.n491 B.n211 163.367
R760 B.n499 B.n211 163.367
R761 B.n499 B.n209 163.367
R762 B.n503 B.n209 163.367
R763 B.n503 B.n203 163.367
R764 B.n512 B.n203 163.367
R765 B.n512 B.n201 163.367
R766 B.n516 B.n201 163.367
R767 B.n516 B.n3 163.367
R768 B.n660 B.n3 163.367
R769 B.n656 B.n2 163.367
R770 B.n656 B.n655 163.367
R771 B.n655 B.n9 163.367
R772 B.n651 B.n9 163.367
R773 B.n651 B.n11 163.367
R774 B.n647 B.n11 163.367
R775 B.n647 B.n17 163.367
R776 B.n643 B.n17 163.367
R777 B.n643 B.n19 163.367
R778 B.n639 B.n19 163.367
R779 B.n639 B.n23 163.367
R780 B.n635 B.n23 163.367
R781 B.n635 B.n25 163.367
R782 B.n631 B.n25 163.367
R783 B.n631 B.n31 163.367
R784 B.n627 B.n31 163.367
R785 B.n627 B.n33 163.367
R786 B.n623 B.n33 163.367
R787 B.n623 B.n38 163.367
R788 B.n619 B.n38 163.367
R789 B.n619 B.n40 163.367
R790 B.n615 B.n40 163.367
R791 B.n615 B.n45 163.367
R792 B.n611 B.n45 163.367
R793 B.n611 B.n47 163.367
R794 B.n607 B.n47 163.367
R795 B.n607 B.n52 163.367
R796 B.n603 B.n52 163.367
R797 B.n603 B.n54 163.367
R798 B.n599 B.n54 163.367
R799 B.n599 B.n59 163.367
R800 B.n595 B.n59 163.367
R801 B.n595 B.n61 163.367
R802 B.n591 B.n61 163.367
R803 B.n591 B.n66 163.367
R804 B.n587 B.n66 163.367
R805 B.n587 B.n68 163.367
R806 B.n583 B.n68 163.367
R807 B.n583 B.n73 163.367
R808 B.n579 B.n73 163.367
R809 B.n401 B.n275 126.203
R810 B.n578 B.n577 126.203
R811 B.n101 B.t17 119.594
R812 B.n286 B.t11 119.594
R813 B.n103 B.t14 119.59
R814 B.n295 B.t21 119.59
R815 B.n401 B.n271 77.3132
R816 B.n407 B.n271 77.3132
R817 B.n407 B.n267 77.3132
R818 B.n413 B.n267 77.3132
R819 B.n413 B.n263 77.3132
R820 B.n419 B.n263 77.3132
R821 B.n425 B.n259 77.3132
R822 B.n425 B.n255 77.3132
R823 B.n431 B.n255 77.3132
R824 B.n431 B.n251 77.3132
R825 B.n437 B.n251 77.3132
R826 B.n437 B.n247 77.3132
R827 B.n443 B.n247 77.3132
R828 B.n443 B.n243 77.3132
R829 B.n449 B.n243 77.3132
R830 B.n455 B.n239 77.3132
R831 B.n455 B.n235 77.3132
R832 B.n461 B.n235 77.3132
R833 B.n461 B.n231 77.3132
R834 B.n467 B.n231 77.3132
R835 B.n473 B.n227 77.3132
R836 B.n473 B.n223 77.3132
R837 B.n479 B.n223 77.3132
R838 B.n479 B.n219 77.3132
R839 B.n486 B.n219 77.3132
R840 B.n486 B.n485 77.3132
R841 B.n492 B.n212 77.3132
R842 B.n498 B.n212 77.3132
R843 B.n498 B.n207 77.3132
R844 B.n504 B.n207 77.3132
R845 B.n504 B.n208 77.3132
R846 B.n511 B.n200 77.3132
R847 B.n517 B.n200 77.3132
R848 B.n517 B.n4 77.3132
R849 B.n659 B.n4 77.3132
R850 B.n659 B.n658 77.3132
R851 B.n658 B.n657 77.3132
R852 B.n657 B.n8 77.3132
R853 B.n12 B.n8 77.3132
R854 B.n650 B.n12 77.3132
R855 B.n649 B.n648 77.3132
R856 B.n648 B.n16 77.3132
R857 B.n642 B.n16 77.3132
R858 B.n642 B.n641 77.3132
R859 B.n641 B.n640 77.3132
R860 B.n634 B.n26 77.3132
R861 B.n634 B.n633 77.3132
R862 B.n633 B.n632 77.3132
R863 B.n632 B.n30 77.3132
R864 B.n626 B.n30 77.3132
R865 B.n626 B.n625 77.3132
R866 B.n624 B.n37 77.3132
R867 B.n618 B.n37 77.3132
R868 B.n618 B.n617 77.3132
R869 B.n617 B.n616 77.3132
R870 B.n616 B.n44 77.3132
R871 B.n610 B.n609 77.3132
R872 B.n609 B.n608 77.3132
R873 B.n608 B.n51 77.3132
R874 B.n602 B.n51 77.3132
R875 B.n602 B.n601 77.3132
R876 B.n601 B.n600 77.3132
R877 B.n600 B.n58 77.3132
R878 B.n594 B.n58 77.3132
R879 B.n594 B.n593 77.3132
R880 B.n592 B.n65 77.3132
R881 B.n586 B.n65 77.3132
R882 B.n586 B.n585 77.3132
R883 B.n585 B.n584 77.3132
R884 B.n584 B.n72 77.3132
R885 B.n578 B.n72 77.3132
R886 B.n102 B.t18 77.1206
R887 B.n287 B.t10 77.1206
R888 B.n104 B.t15 77.1167
R889 B.n296 B.t20 77.1167
R890 B.n77 B.n75 71.676
R891 B.n107 B.n78 71.676
R892 B.n111 B.n79 71.676
R893 B.n115 B.n80 71.676
R894 B.n119 B.n81 71.676
R895 B.n123 B.n82 71.676
R896 B.n127 B.n83 71.676
R897 B.n131 B.n84 71.676
R898 B.n135 B.n85 71.676
R899 B.n139 B.n86 71.676
R900 B.n144 B.n87 71.676
R901 B.n148 B.n88 71.676
R902 B.n152 B.n89 71.676
R903 B.n156 B.n90 71.676
R904 B.n160 B.n91 71.676
R905 B.n165 B.n92 71.676
R906 B.n169 B.n93 71.676
R907 B.n173 B.n94 71.676
R908 B.n177 B.n95 71.676
R909 B.n181 B.n96 71.676
R910 B.n185 B.n97 71.676
R911 B.n189 B.n98 71.676
R912 B.n193 B.n99 71.676
R913 B.n576 B.n100 71.676
R914 B.n576 B.n575 71.676
R915 B.n195 B.n99 71.676
R916 B.n192 B.n98 71.676
R917 B.n188 B.n97 71.676
R918 B.n184 B.n96 71.676
R919 B.n180 B.n95 71.676
R920 B.n176 B.n94 71.676
R921 B.n172 B.n93 71.676
R922 B.n168 B.n92 71.676
R923 B.n164 B.n91 71.676
R924 B.n159 B.n90 71.676
R925 B.n155 B.n89 71.676
R926 B.n151 B.n88 71.676
R927 B.n147 B.n87 71.676
R928 B.n143 B.n86 71.676
R929 B.n138 B.n85 71.676
R930 B.n134 B.n84 71.676
R931 B.n130 B.n83 71.676
R932 B.n126 B.n82 71.676
R933 B.n122 B.n81 71.676
R934 B.n118 B.n80 71.676
R935 B.n114 B.n79 71.676
R936 B.n110 B.n78 71.676
R937 B.n106 B.n77 71.676
R938 B.n305 B.n274 71.676
R939 B.n311 B.n310 71.676
R940 B.n314 B.n313 71.676
R941 B.n319 B.n318 71.676
R942 B.n322 B.n321 71.676
R943 B.n327 B.n326 71.676
R944 B.n330 B.n329 71.676
R945 B.n335 B.n334 71.676
R946 B.n338 B.n337 71.676
R947 B.n344 B.n343 71.676
R948 B.n347 B.n346 71.676
R949 B.n352 B.n351 71.676
R950 B.n355 B.n354 71.676
R951 B.n360 B.n359 71.676
R952 B.n363 B.n362 71.676
R953 B.n368 B.n367 71.676
R954 B.n371 B.n370 71.676
R955 B.n376 B.n375 71.676
R956 B.n379 B.n378 71.676
R957 B.n384 B.n383 71.676
R958 B.n387 B.n386 71.676
R959 B.n392 B.n391 71.676
R960 B.n395 B.n394 71.676
R961 B.n306 B.n305 71.676
R962 B.n312 B.n311 71.676
R963 B.n313 B.n302 71.676
R964 B.n320 B.n319 71.676
R965 B.n321 B.n300 71.676
R966 B.n328 B.n327 71.676
R967 B.n329 B.n298 71.676
R968 B.n336 B.n335 71.676
R969 B.n337 B.n294 71.676
R970 B.n345 B.n344 71.676
R971 B.n346 B.n292 71.676
R972 B.n353 B.n352 71.676
R973 B.n354 B.n290 71.676
R974 B.n361 B.n360 71.676
R975 B.n362 B.n285 71.676
R976 B.n369 B.n368 71.676
R977 B.n370 B.n283 71.676
R978 B.n377 B.n376 71.676
R979 B.n378 B.n281 71.676
R980 B.n385 B.n384 71.676
R981 B.n386 B.n279 71.676
R982 B.n393 B.n392 71.676
R983 B.n396 B.n395 71.676
R984 B.n661 B.n660 71.676
R985 B.n661 B.n2 71.676
R986 B.n467 B.t0 61.3958
R987 B.t1 B.n624 61.3958
R988 B.n141 B.n104 59.5399
R989 B.n162 B.n102 59.5399
R990 B.n288 B.n287 59.5399
R991 B.n341 B.n296 59.5399
R992 B.n492 B.t7 59.1219
R993 B.n640 B.t4 59.1219
R994 B.n419 B.t9 54.5741
R995 B.t13 B.n592 54.5741
R996 B.n208 B.t3 52.3002
R997 B.t5 B.n649 52.3002
R998 B.t2 B.n239 50.0263
R999 B.t6 B.n44 50.0263
R1000 B.n104 B.n103 42.4732
R1001 B.n102 B.n101 42.4732
R1002 B.n287 B.n286 42.4732
R1003 B.n296 B.n295 42.4732
R1004 B.n403 B.n273 31.0639
R1005 B.n399 B.n398 31.0639
R1006 B.n574 B.n573 31.0639
R1007 B.n580 B.n74 31.0639
R1008 B.n449 B.t2 27.2873
R1009 B.n610 B.t6 27.2873
R1010 B.n511 B.t3 25.0134
R1011 B.n650 B.t5 25.0134
R1012 B.t9 B.n259 22.7395
R1013 B.n593 B.t13 22.7395
R1014 B.n485 B.t7 18.1917
R1015 B.n26 B.t4 18.1917
R1016 B B.n662 18.0485
R1017 B.t0 B.n227 15.9178
R1018 B.n625 B.t1 15.9178
R1019 B.n404 B.n403 10.6151
R1020 B.n405 B.n404 10.6151
R1021 B.n405 B.n265 10.6151
R1022 B.n415 B.n265 10.6151
R1023 B.n416 B.n415 10.6151
R1024 B.n417 B.n416 10.6151
R1025 B.n417 B.n257 10.6151
R1026 B.n427 B.n257 10.6151
R1027 B.n428 B.n427 10.6151
R1028 B.n429 B.n428 10.6151
R1029 B.n429 B.n249 10.6151
R1030 B.n439 B.n249 10.6151
R1031 B.n440 B.n439 10.6151
R1032 B.n441 B.n440 10.6151
R1033 B.n441 B.n241 10.6151
R1034 B.n451 B.n241 10.6151
R1035 B.n452 B.n451 10.6151
R1036 B.n453 B.n452 10.6151
R1037 B.n453 B.n233 10.6151
R1038 B.n463 B.n233 10.6151
R1039 B.n464 B.n463 10.6151
R1040 B.n465 B.n464 10.6151
R1041 B.n465 B.n225 10.6151
R1042 B.n475 B.n225 10.6151
R1043 B.n476 B.n475 10.6151
R1044 B.n477 B.n476 10.6151
R1045 B.n477 B.n217 10.6151
R1046 B.n488 B.n217 10.6151
R1047 B.n489 B.n488 10.6151
R1048 B.n490 B.n489 10.6151
R1049 B.n490 B.n210 10.6151
R1050 B.n500 B.n210 10.6151
R1051 B.n501 B.n500 10.6151
R1052 B.n502 B.n501 10.6151
R1053 B.n502 B.n202 10.6151
R1054 B.n513 B.n202 10.6151
R1055 B.n514 B.n513 10.6151
R1056 B.n515 B.n514 10.6151
R1057 B.n515 B.n0 10.6151
R1058 B.n307 B.n273 10.6151
R1059 B.n308 B.n307 10.6151
R1060 B.n309 B.n308 10.6151
R1061 B.n309 B.n303 10.6151
R1062 B.n315 B.n303 10.6151
R1063 B.n316 B.n315 10.6151
R1064 B.n317 B.n316 10.6151
R1065 B.n317 B.n301 10.6151
R1066 B.n323 B.n301 10.6151
R1067 B.n324 B.n323 10.6151
R1068 B.n325 B.n324 10.6151
R1069 B.n325 B.n299 10.6151
R1070 B.n331 B.n299 10.6151
R1071 B.n332 B.n331 10.6151
R1072 B.n333 B.n332 10.6151
R1073 B.n333 B.n297 10.6151
R1074 B.n339 B.n297 10.6151
R1075 B.n340 B.n339 10.6151
R1076 B.n342 B.n293 10.6151
R1077 B.n348 B.n293 10.6151
R1078 B.n349 B.n348 10.6151
R1079 B.n350 B.n349 10.6151
R1080 B.n350 B.n291 10.6151
R1081 B.n356 B.n291 10.6151
R1082 B.n357 B.n356 10.6151
R1083 B.n358 B.n357 10.6151
R1084 B.n358 B.n289 10.6151
R1085 B.n365 B.n364 10.6151
R1086 B.n366 B.n365 10.6151
R1087 B.n366 B.n284 10.6151
R1088 B.n372 B.n284 10.6151
R1089 B.n373 B.n372 10.6151
R1090 B.n374 B.n373 10.6151
R1091 B.n374 B.n282 10.6151
R1092 B.n380 B.n282 10.6151
R1093 B.n381 B.n380 10.6151
R1094 B.n382 B.n381 10.6151
R1095 B.n382 B.n280 10.6151
R1096 B.n388 B.n280 10.6151
R1097 B.n389 B.n388 10.6151
R1098 B.n390 B.n389 10.6151
R1099 B.n390 B.n278 10.6151
R1100 B.n278 B.n277 10.6151
R1101 B.n397 B.n277 10.6151
R1102 B.n398 B.n397 10.6151
R1103 B.n399 B.n269 10.6151
R1104 B.n409 B.n269 10.6151
R1105 B.n410 B.n409 10.6151
R1106 B.n411 B.n410 10.6151
R1107 B.n411 B.n261 10.6151
R1108 B.n421 B.n261 10.6151
R1109 B.n422 B.n421 10.6151
R1110 B.n423 B.n422 10.6151
R1111 B.n423 B.n253 10.6151
R1112 B.n433 B.n253 10.6151
R1113 B.n434 B.n433 10.6151
R1114 B.n435 B.n434 10.6151
R1115 B.n435 B.n245 10.6151
R1116 B.n445 B.n245 10.6151
R1117 B.n446 B.n445 10.6151
R1118 B.n447 B.n446 10.6151
R1119 B.n447 B.n237 10.6151
R1120 B.n457 B.n237 10.6151
R1121 B.n458 B.n457 10.6151
R1122 B.n459 B.n458 10.6151
R1123 B.n459 B.n229 10.6151
R1124 B.n469 B.n229 10.6151
R1125 B.n470 B.n469 10.6151
R1126 B.n471 B.n470 10.6151
R1127 B.n471 B.n221 10.6151
R1128 B.n481 B.n221 10.6151
R1129 B.n482 B.n481 10.6151
R1130 B.n483 B.n482 10.6151
R1131 B.n483 B.n214 10.6151
R1132 B.n494 B.n214 10.6151
R1133 B.n495 B.n494 10.6151
R1134 B.n496 B.n495 10.6151
R1135 B.n496 B.n205 10.6151
R1136 B.n506 B.n205 10.6151
R1137 B.n507 B.n506 10.6151
R1138 B.n509 B.n507 10.6151
R1139 B.n509 B.n508 10.6151
R1140 B.n508 B.n198 10.6151
R1141 B.n520 B.n198 10.6151
R1142 B.n521 B.n520 10.6151
R1143 B.n522 B.n521 10.6151
R1144 B.n523 B.n522 10.6151
R1145 B.n524 B.n523 10.6151
R1146 B.n527 B.n524 10.6151
R1147 B.n528 B.n527 10.6151
R1148 B.n529 B.n528 10.6151
R1149 B.n530 B.n529 10.6151
R1150 B.n532 B.n530 10.6151
R1151 B.n533 B.n532 10.6151
R1152 B.n534 B.n533 10.6151
R1153 B.n535 B.n534 10.6151
R1154 B.n537 B.n535 10.6151
R1155 B.n538 B.n537 10.6151
R1156 B.n539 B.n538 10.6151
R1157 B.n540 B.n539 10.6151
R1158 B.n542 B.n540 10.6151
R1159 B.n543 B.n542 10.6151
R1160 B.n544 B.n543 10.6151
R1161 B.n545 B.n544 10.6151
R1162 B.n547 B.n545 10.6151
R1163 B.n548 B.n547 10.6151
R1164 B.n549 B.n548 10.6151
R1165 B.n550 B.n549 10.6151
R1166 B.n552 B.n550 10.6151
R1167 B.n553 B.n552 10.6151
R1168 B.n554 B.n553 10.6151
R1169 B.n555 B.n554 10.6151
R1170 B.n557 B.n555 10.6151
R1171 B.n558 B.n557 10.6151
R1172 B.n559 B.n558 10.6151
R1173 B.n560 B.n559 10.6151
R1174 B.n562 B.n560 10.6151
R1175 B.n563 B.n562 10.6151
R1176 B.n564 B.n563 10.6151
R1177 B.n565 B.n564 10.6151
R1178 B.n567 B.n565 10.6151
R1179 B.n568 B.n567 10.6151
R1180 B.n569 B.n568 10.6151
R1181 B.n570 B.n569 10.6151
R1182 B.n572 B.n570 10.6151
R1183 B.n573 B.n572 10.6151
R1184 B.n654 B.n1 10.6151
R1185 B.n654 B.n653 10.6151
R1186 B.n653 B.n652 10.6151
R1187 B.n652 B.n10 10.6151
R1188 B.n646 B.n10 10.6151
R1189 B.n646 B.n645 10.6151
R1190 B.n645 B.n644 10.6151
R1191 B.n644 B.n18 10.6151
R1192 B.n638 B.n18 10.6151
R1193 B.n638 B.n637 10.6151
R1194 B.n637 B.n636 10.6151
R1195 B.n636 B.n24 10.6151
R1196 B.n630 B.n24 10.6151
R1197 B.n630 B.n629 10.6151
R1198 B.n629 B.n628 10.6151
R1199 B.n628 B.n32 10.6151
R1200 B.n622 B.n32 10.6151
R1201 B.n622 B.n621 10.6151
R1202 B.n621 B.n620 10.6151
R1203 B.n620 B.n39 10.6151
R1204 B.n614 B.n39 10.6151
R1205 B.n614 B.n613 10.6151
R1206 B.n613 B.n612 10.6151
R1207 B.n612 B.n46 10.6151
R1208 B.n606 B.n46 10.6151
R1209 B.n606 B.n605 10.6151
R1210 B.n605 B.n604 10.6151
R1211 B.n604 B.n53 10.6151
R1212 B.n598 B.n53 10.6151
R1213 B.n598 B.n597 10.6151
R1214 B.n597 B.n596 10.6151
R1215 B.n596 B.n60 10.6151
R1216 B.n590 B.n60 10.6151
R1217 B.n590 B.n589 10.6151
R1218 B.n589 B.n588 10.6151
R1219 B.n588 B.n67 10.6151
R1220 B.n582 B.n67 10.6151
R1221 B.n582 B.n581 10.6151
R1222 B.n581 B.n580 10.6151
R1223 B.n105 B.n74 10.6151
R1224 B.n108 B.n105 10.6151
R1225 B.n109 B.n108 10.6151
R1226 B.n112 B.n109 10.6151
R1227 B.n113 B.n112 10.6151
R1228 B.n116 B.n113 10.6151
R1229 B.n117 B.n116 10.6151
R1230 B.n120 B.n117 10.6151
R1231 B.n121 B.n120 10.6151
R1232 B.n124 B.n121 10.6151
R1233 B.n125 B.n124 10.6151
R1234 B.n128 B.n125 10.6151
R1235 B.n129 B.n128 10.6151
R1236 B.n132 B.n129 10.6151
R1237 B.n133 B.n132 10.6151
R1238 B.n136 B.n133 10.6151
R1239 B.n137 B.n136 10.6151
R1240 B.n140 B.n137 10.6151
R1241 B.n145 B.n142 10.6151
R1242 B.n146 B.n145 10.6151
R1243 B.n149 B.n146 10.6151
R1244 B.n150 B.n149 10.6151
R1245 B.n153 B.n150 10.6151
R1246 B.n154 B.n153 10.6151
R1247 B.n157 B.n154 10.6151
R1248 B.n158 B.n157 10.6151
R1249 B.n161 B.n158 10.6151
R1250 B.n166 B.n163 10.6151
R1251 B.n167 B.n166 10.6151
R1252 B.n170 B.n167 10.6151
R1253 B.n171 B.n170 10.6151
R1254 B.n174 B.n171 10.6151
R1255 B.n175 B.n174 10.6151
R1256 B.n178 B.n175 10.6151
R1257 B.n179 B.n178 10.6151
R1258 B.n182 B.n179 10.6151
R1259 B.n183 B.n182 10.6151
R1260 B.n186 B.n183 10.6151
R1261 B.n187 B.n186 10.6151
R1262 B.n190 B.n187 10.6151
R1263 B.n191 B.n190 10.6151
R1264 B.n194 B.n191 10.6151
R1265 B.n196 B.n194 10.6151
R1266 B.n197 B.n196 10.6151
R1267 B.n574 B.n197 10.6151
R1268 B.n341 B.n340 9.36635
R1269 B.n364 B.n288 9.36635
R1270 B.n141 B.n140 9.36635
R1271 B.n163 B.n162 9.36635
R1272 B.n662 B.n0 8.11757
R1273 B.n662 B.n1 8.11757
R1274 B.n342 B.n341 1.24928
R1275 B.n289 B.n288 1.24928
R1276 B.n142 B.n141 1.24928
R1277 B.n162 B.n161 1.24928
R1278 VP.n31 VP.n7 184.171
R1279 VP.n56 VP.n55 184.171
R1280 VP.n30 VP.n29 184.171
R1281 VP.n15 VP.n12 161.3
R1282 VP.n17 VP.n16 161.3
R1283 VP.n18 VP.n11 161.3
R1284 VP.n20 VP.n19 161.3
R1285 VP.n22 VP.n10 161.3
R1286 VP.n24 VP.n23 161.3
R1287 VP.n25 VP.n9 161.3
R1288 VP.n27 VP.n26 161.3
R1289 VP.n28 VP.n8 161.3
R1290 VP.n54 VP.n0 161.3
R1291 VP.n53 VP.n52 161.3
R1292 VP.n51 VP.n1 161.3
R1293 VP.n50 VP.n49 161.3
R1294 VP.n48 VP.n2 161.3
R1295 VP.n46 VP.n45 161.3
R1296 VP.n44 VP.n3 161.3
R1297 VP.n43 VP.n42 161.3
R1298 VP.n41 VP.n4 161.3
R1299 VP.n39 VP.n38 161.3
R1300 VP.n37 VP.n5 161.3
R1301 VP.n36 VP.n35 161.3
R1302 VP.n34 VP.n6 161.3
R1303 VP.n33 VP.n32 161.3
R1304 VP.n13 VP.t4 89.9794
R1305 VP.n7 VP.t1 57.0113
R1306 VP.n40 VP.t7 57.0113
R1307 VP.n47 VP.t3 57.0113
R1308 VP.n55 VP.t0 57.0113
R1309 VP.n29 VP.t6 57.0113
R1310 VP.n21 VP.t2 57.0113
R1311 VP.n14 VP.t5 57.0113
R1312 VP.n42 VP.n3 56.5617
R1313 VP.n16 VP.n11 56.5617
R1314 VP.n14 VP.n13 53.0172
R1315 VP.n35 VP.n5 46.3896
R1316 VP.n49 VP.n1 46.3896
R1317 VP.n23 VP.n9 46.3896
R1318 VP.n31 VP.n30 41.5611
R1319 VP.n35 VP.n34 34.7644
R1320 VP.n53 VP.n1 34.7644
R1321 VP.n27 VP.n9 34.7644
R1322 VP.n34 VP.n33 24.5923
R1323 VP.n39 VP.n5 24.5923
R1324 VP.n42 VP.n41 24.5923
R1325 VP.n46 VP.n3 24.5923
R1326 VP.n49 VP.n48 24.5923
R1327 VP.n54 VP.n53 24.5923
R1328 VP.n28 VP.n27 24.5923
R1329 VP.n20 VP.n11 24.5923
R1330 VP.n23 VP.n22 24.5923
R1331 VP.n16 VP.n15 24.5923
R1332 VP.n41 VP.n40 16.9689
R1333 VP.n47 VP.n46 16.9689
R1334 VP.n21 VP.n20 16.9689
R1335 VP.n15 VP.n14 16.9689
R1336 VP.n13 VP.n12 12.4356
R1337 VP.n40 VP.n39 7.62397
R1338 VP.n48 VP.n47 7.62397
R1339 VP.n22 VP.n21 7.62397
R1340 VP.n33 VP.n7 1.72193
R1341 VP.n55 VP.n54 1.72193
R1342 VP.n29 VP.n28 1.72193
R1343 VP.n17 VP.n12 0.189894
R1344 VP.n18 VP.n17 0.189894
R1345 VP.n19 VP.n18 0.189894
R1346 VP.n19 VP.n10 0.189894
R1347 VP.n24 VP.n10 0.189894
R1348 VP.n25 VP.n24 0.189894
R1349 VP.n26 VP.n25 0.189894
R1350 VP.n26 VP.n8 0.189894
R1351 VP.n30 VP.n8 0.189894
R1352 VP.n32 VP.n31 0.189894
R1353 VP.n32 VP.n6 0.189894
R1354 VP.n36 VP.n6 0.189894
R1355 VP.n37 VP.n36 0.189894
R1356 VP.n38 VP.n37 0.189894
R1357 VP.n38 VP.n4 0.189894
R1358 VP.n43 VP.n4 0.189894
R1359 VP.n44 VP.n43 0.189894
R1360 VP.n45 VP.n44 0.189894
R1361 VP.n45 VP.n2 0.189894
R1362 VP.n50 VP.n2 0.189894
R1363 VP.n51 VP.n50 0.189894
R1364 VP.n52 VP.n51 0.189894
R1365 VP.n52 VP.n0 0.189894
R1366 VP.n56 VP.n0 0.189894
R1367 VP VP.n56 0.0516364
R1368 VDD1 VDD1.n0 76.7994
R1369 VDD1.n3 VDD1.n2 76.6856
R1370 VDD1.n3 VDD1.n1 76.6856
R1371 VDD1.n5 VDD1.n4 75.7971
R1372 VDD1.n5 VDD1.n3 36.5871
R1373 VDD1.n4 VDD1.t5 4.5005
R1374 VDD1.n4 VDD1.t1 4.5005
R1375 VDD1.n0 VDD1.t3 4.5005
R1376 VDD1.n0 VDD1.t2 4.5005
R1377 VDD1.n2 VDD1.t4 4.5005
R1378 VDD1.n2 VDD1.t7 4.5005
R1379 VDD1.n1 VDD1.t6 4.5005
R1380 VDD1.n1 VDD1.t0 4.5005
R1381 VDD1 VDD1.n5 0.886276
C0 VP VN 5.3503f
C1 VDD1 VTAIL 5.07247f
C2 VDD2 VDD1 1.39021f
C3 VDD2 VTAIL 5.12193f
C4 VDD1 VN 0.154495f
C5 VP VDD1 3.52161f
C6 VN VTAIL 3.84862f
C7 VDD2 VN 3.23217f
C8 VP VTAIL 3.86273f
C9 VDD2 VP 0.445484f
C10 VDD2 B 4.023432f
C11 VDD1 B 4.390216f
C12 VTAIL B 5.166425f
C13 VN B 11.89497f
C14 VP B 10.467248f
C15 VDD1.t3 B 0.086753f
C16 VDD1.t2 B 0.086753f
C17 VDD1.n0 B 0.697967f
C18 VDD1.t6 B 0.086753f
C19 VDD1.t0 B 0.086753f
C20 VDD1.n1 B 0.697225f
C21 VDD1.t4 B 0.086753f
C22 VDD1.t7 B 0.086753f
C23 VDD1.n2 B 0.697225f
C24 VDD1.n3 B 2.4199f
C25 VDD1.t5 B 0.086753f
C26 VDD1.t1 B 0.086753f
C27 VDD1.n4 B 0.692233f
C28 VDD1.n5 B 2.11625f
C29 VP.n0 B 0.031925f
C30 VP.t0 B 0.676747f
C31 VP.n1 B 0.027281f
C32 VP.n2 B 0.031925f
C33 VP.t3 B 0.676747f
C34 VP.n3 B 0.046408f
C35 VP.n4 B 0.031925f
C36 VP.t7 B 0.676747f
C37 VP.n5 B 0.060576f
C38 VP.n6 B 0.031925f
C39 VP.t1 B 0.676747f
C40 VP.n7 B 0.345372f
C41 VP.n8 B 0.031925f
C42 VP.t6 B 0.676747f
C43 VP.n9 B 0.027281f
C44 VP.n10 B 0.031925f
C45 VP.t2 B 0.676747f
C46 VP.n11 B 0.046408f
C47 VP.n12 B 0.235718f
C48 VP.t5 B 0.676747f
C49 VP.t4 B 0.833107f
C50 VP.n13 B 0.340875f
C51 VP.n14 B 0.350955f
C52 VP.n15 B 0.050142f
C53 VP.n16 B 0.046408f
C54 VP.n17 B 0.031925f
C55 VP.n18 B 0.031925f
C56 VP.n19 B 0.031925f
C57 VP.n20 B 0.050142f
C58 VP.n21 B 0.2733f
C59 VP.n22 B 0.039036f
C60 VP.n23 B 0.060576f
C61 VP.n24 B 0.031925f
C62 VP.n25 B 0.031925f
C63 VP.n26 B 0.031925f
C64 VP.n27 B 0.064163f
C65 VP.n28 B 0.032022f
C66 VP.n29 B 0.345372f
C67 VP.n30 B 1.305f
C68 VP.n31 B 1.3327f
C69 VP.n32 B 0.031925f
C70 VP.n33 B 0.032022f
C71 VP.n34 B 0.064163f
C72 VP.n35 B 0.027281f
C73 VP.n36 B 0.031925f
C74 VP.n37 B 0.031925f
C75 VP.n38 B 0.031925f
C76 VP.n39 B 0.039036f
C77 VP.n40 B 0.2733f
C78 VP.n41 B 0.050142f
C79 VP.n42 B 0.046408f
C80 VP.n43 B 0.031925f
C81 VP.n44 B 0.031925f
C82 VP.n45 B 0.031925f
C83 VP.n46 B 0.050142f
C84 VP.n47 B 0.2733f
C85 VP.n48 B 0.039036f
C86 VP.n49 B 0.060576f
C87 VP.n50 B 0.031925f
C88 VP.n51 B 0.031925f
C89 VP.n52 B 0.031925f
C90 VP.n53 B 0.064163f
C91 VP.n54 B 0.032022f
C92 VP.n55 B 0.345372f
C93 VP.n56 B 0.03496f
C94 VTAIL.t12 B 0.083445f
C95 VTAIL.t8 B 0.083445f
C96 VTAIL.n0 B 0.613742f
C97 VTAIL.n1 B 0.359194f
C98 VTAIL.t14 B 0.787712f
C99 VTAIL.n2 B 0.444634f
C100 VTAIL.t3 B 0.787712f
C101 VTAIL.n3 B 0.444634f
C102 VTAIL.t0 B 0.083445f
C103 VTAIL.t7 B 0.083445f
C104 VTAIL.n4 B 0.613742f
C105 VTAIL.n5 B 0.500689f
C106 VTAIL.t2 B 0.787712f
C107 VTAIL.n6 B 1.17362f
C108 VTAIL.t13 B 0.787715f
C109 VTAIL.n7 B 1.17362f
C110 VTAIL.t9 B 0.083445f
C111 VTAIL.t15 B 0.083445f
C112 VTAIL.n8 B 0.613745f
C113 VTAIL.n9 B 0.500686f
C114 VTAIL.t10 B 0.787715f
C115 VTAIL.n10 B 0.444632f
C116 VTAIL.t5 B 0.787715f
C117 VTAIL.n11 B 0.444632f
C118 VTAIL.t4 B 0.083445f
C119 VTAIL.t1 B 0.083445f
C120 VTAIL.n12 B 0.613745f
C121 VTAIL.n13 B 0.500686f
C122 VTAIL.t6 B 0.787712f
C123 VTAIL.n14 B 1.17362f
C124 VTAIL.t11 B 0.787712f
C125 VTAIL.n15 B 1.16912f
C126 VDD2.t0 B 0.084634f
C127 VDD2.t7 B 0.084634f
C128 VDD2.n0 B 0.680191f
C129 VDD2.t3 B 0.084634f
C130 VDD2.t6 B 0.084634f
C131 VDD2.n1 B 0.680191f
C132 VDD2.n2 B 2.30943f
C133 VDD2.t1 B 0.084634f
C134 VDD2.t2 B 0.084634f
C135 VDD2.n3 B 0.675325f
C136 VDD2.n4 B 2.03512f
C137 VDD2.t4 B 0.084634f
C138 VDD2.t5 B 0.084634f
C139 VDD2.n5 B 0.680165f
C140 VN.n0 B 0.030819f
C141 VN.t4 B 0.653309f
C142 VN.n1 B 0.026336f
C143 VN.n2 B 0.030819f
C144 VN.t7 B 0.653309f
C145 VN.n3 B 0.044801f
C146 VN.n4 B 0.227554f
C147 VN.t3 B 0.653309f
C148 VN.t1 B 0.804253f
C149 VN.n5 B 0.329069f
C150 VN.n6 B 0.3388f
C151 VN.n7 B 0.048405f
C152 VN.n8 B 0.044801f
C153 VN.n9 B 0.030819f
C154 VN.n10 B 0.030819f
C155 VN.n11 B 0.030819f
C156 VN.n12 B 0.048405f
C157 VN.n13 B 0.263834f
C158 VN.n14 B 0.037684f
C159 VN.n15 B 0.058478f
C160 VN.n16 B 0.030819f
C161 VN.n17 B 0.030819f
C162 VN.n18 B 0.030819f
C163 VN.n19 B 0.06194f
C164 VN.n20 B 0.030912f
C165 VN.n21 B 0.33341f
C166 VN.n22 B 0.033749f
C167 VN.n23 B 0.030819f
C168 VN.t2 B 0.653309f
C169 VN.n24 B 0.026336f
C170 VN.n25 B 0.030819f
C171 VN.t6 B 0.653309f
C172 VN.n26 B 0.044801f
C173 VN.n27 B 0.227554f
C174 VN.t0 B 0.653309f
C175 VN.t5 B 0.804253f
C176 VN.n28 B 0.329069f
C177 VN.n29 B 0.3388f
C178 VN.n30 B 0.048405f
C179 VN.n31 B 0.044801f
C180 VN.n32 B 0.030819f
C181 VN.n33 B 0.030819f
C182 VN.n34 B 0.030819f
C183 VN.n35 B 0.048405f
C184 VN.n36 B 0.263834f
C185 VN.n37 B 0.037684f
C186 VN.n38 B 0.058478f
C187 VN.n39 B 0.030819f
C188 VN.n40 B 0.030819f
C189 VN.n41 B 0.030819f
C190 VN.n42 B 0.06194f
C191 VN.n43 B 0.030912f
C192 VN.n44 B 0.33341f
C193 VN.n45 B 1.28005f
.ends

