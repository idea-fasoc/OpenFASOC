* NGSPICE file created from diff_pair_sample_0671.ext - technology: sky130A

.subckt diff_pair_sample_0671 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=5.3079 ps=28 w=13.61 l=0.84
X1 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=5.3079 ps=28 w=13.61 l=0.84
X2 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=0 ps=0 w=13.61 l=0.84
X3 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=5.3079 ps=28 w=13.61 l=0.84
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=0 ps=0 w=13.61 l=0.84
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=0 ps=0 w=13.61 l=0.84
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=5.3079 ps=28 w=13.61 l=0.84
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3079 pd=28 as=0 ps=0 w=13.61 l=0.84
R0 VN VN.t0 640.434
R1 VN VN.t1 598.881
R2 VTAIL.n1 VTAIL.t0 46.8128
R3 VTAIL.n3 VTAIL.t1 46.8127
R4 VTAIL.n0 VTAIL.t3 46.8127
R5 VTAIL.n2 VTAIL.t2 46.8127
R6 VTAIL.n1 VTAIL.n0 26.1341
R7 VTAIL.n3 VTAIL.n2 25.1255
R8 VTAIL.n2 VTAIL.n1 0.974638
R9 VTAIL VTAIL.n0 0.780672
R10 VTAIL VTAIL.n3 0.194466
R11 VDD2.n0 VDD2.t0 100.918
R12 VDD2.n0 VDD2.t1 63.4914
R13 VDD2 VDD2.n0 0.310845
R14 B.n370 B.t13 592.179
R15 B.n368 B.t2 592.179
R16 B.n87 B.t10 592.179
R17 B.n84 B.t6 592.179
R18 B.n640 B.n639 585
R19 B.n286 B.n82 585
R20 B.n285 B.n284 585
R21 B.n283 B.n282 585
R22 B.n281 B.n280 585
R23 B.n279 B.n278 585
R24 B.n277 B.n276 585
R25 B.n275 B.n274 585
R26 B.n273 B.n272 585
R27 B.n271 B.n270 585
R28 B.n269 B.n268 585
R29 B.n267 B.n266 585
R30 B.n265 B.n264 585
R31 B.n263 B.n262 585
R32 B.n261 B.n260 585
R33 B.n259 B.n258 585
R34 B.n257 B.n256 585
R35 B.n255 B.n254 585
R36 B.n253 B.n252 585
R37 B.n251 B.n250 585
R38 B.n249 B.n248 585
R39 B.n247 B.n246 585
R40 B.n245 B.n244 585
R41 B.n243 B.n242 585
R42 B.n241 B.n240 585
R43 B.n239 B.n238 585
R44 B.n237 B.n236 585
R45 B.n235 B.n234 585
R46 B.n233 B.n232 585
R47 B.n231 B.n230 585
R48 B.n229 B.n228 585
R49 B.n227 B.n226 585
R50 B.n225 B.n224 585
R51 B.n223 B.n222 585
R52 B.n221 B.n220 585
R53 B.n219 B.n218 585
R54 B.n217 B.n216 585
R55 B.n215 B.n214 585
R56 B.n213 B.n212 585
R57 B.n211 B.n210 585
R58 B.n209 B.n208 585
R59 B.n207 B.n206 585
R60 B.n205 B.n204 585
R61 B.n203 B.n202 585
R62 B.n201 B.n200 585
R63 B.n199 B.n198 585
R64 B.n197 B.n196 585
R65 B.n195 B.n194 585
R66 B.n193 B.n192 585
R67 B.n191 B.n190 585
R68 B.n189 B.n188 585
R69 B.n187 B.n186 585
R70 B.n185 B.n184 585
R71 B.n183 B.n182 585
R72 B.n181 B.n180 585
R73 B.n179 B.n178 585
R74 B.n177 B.n176 585
R75 B.n175 B.n174 585
R76 B.n173 B.n172 585
R77 B.n171 B.n170 585
R78 B.n169 B.n168 585
R79 B.n167 B.n166 585
R80 B.n165 B.n164 585
R81 B.n163 B.n162 585
R82 B.n161 B.n160 585
R83 B.n159 B.n158 585
R84 B.n157 B.n156 585
R85 B.n155 B.n154 585
R86 B.n153 B.n152 585
R87 B.n151 B.n150 585
R88 B.n149 B.n148 585
R89 B.n147 B.n146 585
R90 B.n145 B.n144 585
R91 B.n143 B.n142 585
R92 B.n141 B.n140 585
R93 B.n139 B.n138 585
R94 B.n137 B.n136 585
R95 B.n135 B.n134 585
R96 B.n133 B.n132 585
R97 B.n131 B.n130 585
R98 B.n129 B.n128 585
R99 B.n127 B.n126 585
R100 B.n125 B.n124 585
R101 B.n123 B.n122 585
R102 B.n121 B.n120 585
R103 B.n119 B.n118 585
R104 B.n117 B.n116 585
R105 B.n115 B.n114 585
R106 B.n113 B.n112 585
R107 B.n111 B.n110 585
R108 B.n109 B.n108 585
R109 B.n107 B.n106 585
R110 B.n105 B.n104 585
R111 B.n103 B.n102 585
R112 B.n101 B.n100 585
R113 B.n99 B.n98 585
R114 B.n97 B.n96 585
R115 B.n95 B.n94 585
R116 B.n93 B.n92 585
R117 B.n91 B.n90 585
R118 B.n32 B.n31 585
R119 B.n645 B.n644 585
R120 B.n638 B.n83 585
R121 B.n83 B.n29 585
R122 B.n637 B.n28 585
R123 B.n649 B.n28 585
R124 B.n636 B.n27 585
R125 B.n650 B.n27 585
R126 B.n635 B.n26 585
R127 B.n651 B.n26 585
R128 B.n634 B.n633 585
R129 B.n633 B.n22 585
R130 B.n632 B.n21 585
R131 B.n657 B.n21 585
R132 B.n631 B.n20 585
R133 B.n658 B.n20 585
R134 B.n630 B.n19 585
R135 B.n659 B.n19 585
R136 B.n629 B.n628 585
R137 B.n628 B.n15 585
R138 B.n627 B.n14 585
R139 B.n665 B.n14 585
R140 B.n626 B.n13 585
R141 B.n666 B.n13 585
R142 B.n625 B.n12 585
R143 B.n667 B.n12 585
R144 B.n624 B.n623 585
R145 B.n623 B.n8 585
R146 B.n622 B.n7 585
R147 B.n673 B.n7 585
R148 B.n621 B.n6 585
R149 B.n674 B.n6 585
R150 B.n620 B.n5 585
R151 B.n675 B.n5 585
R152 B.n619 B.n618 585
R153 B.n618 B.n4 585
R154 B.n617 B.n287 585
R155 B.n617 B.n616 585
R156 B.n607 B.n288 585
R157 B.n289 B.n288 585
R158 B.n609 B.n608 585
R159 B.n610 B.n609 585
R160 B.n606 B.n294 585
R161 B.n294 B.n293 585
R162 B.n605 B.n604 585
R163 B.n604 B.n603 585
R164 B.n296 B.n295 585
R165 B.n297 B.n296 585
R166 B.n596 B.n595 585
R167 B.n597 B.n596 585
R168 B.n594 B.n302 585
R169 B.n302 B.n301 585
R170 B.n593 B.n592 585
R171 B.n592 B.n591 585
R172 B.n304 B.n303 585
R173 B.n305 B.n304 585
R174 B.n584 B.n583 585
R175 B.n585 B.n584 585
R176 B.n582 B.n310 585
R177 B.n310 B.n309 585
R178 B.n581 B.n580 585
R179 B.n580 B.n579 585
R180 B.n312 B.n311 585
R181 B.n313 B.n312 585
R182 B.n575 B.n574 585
R183 B.n316 B.n315 585
R184 B.n571 B.n570 585
R185 B.n572 B.n571 585
R186 B.n569 B.n367 585
R187 B.n568 B.n567 585
R188 B.n566 B.n565 585
R189 B.n564 B.n563 585
R190 B.n562 B.n561 585
R191 B.n560 B.n559 585
R192 B.n558 B.n557 585
R193 B.n556 B.n555 585
R194 B.n554 B.n553 585
R195 B.n552 B.n551 585
R196 B.n550 B.n549 585
R197 B.n548 B.n547 585
R198 B.n546 B.n545 585
R199 B.n544 B.n543 585
R200 B.n542 B.n541 585
R201 B.n540 B.n539 585
R202 B.n538 B.n537 585
R203 B.n536 B.n535 585
R204 B.n534 B.n533 585
R205 B.n532 B.n531 585
R206 B.n530 B.n529 585
R207 B.n528 B.n527 585
R208 B.n526 B.n525 585
R209 B.n524 B.n523 585
R210 B.n522 B.n521 585
R211 B.n520 B.n519 585
R212 B.n518 B.n517 585
R213 B.n516 B.n515 585
R214 B.n514 B.n513 585
R215 B.n512 B.n511 585
R216 B.n510 B.n509 585
R217 B.n508 B.n507 585
R218 B.n506 B.n505 585
R219 B.n504 B.n503 585
R220 B.n502 B.n501 585
R221 B.n500 B.n499 585
R222 B.n498 B.n497 585
R223 B.n496 B.n495 585
R224 B.n494 B.n493 585
R225 B.n492 B.n491 585
R226 B.n490 B.n489 585
R227 B.n488 B.n487 585
R228 B.n486 B.n485 585
R229 B.n483 B.n482 585
R230 B.n481 B.n480 585
R231 B.n479 B.n478 585
R232 B.n477 B.n476 585
R233 B.n475 B.n474 585
R234 B.n473 B.n472 585
R235 B.n471 B.n470 585
R236 B.n469 B.n468 585
R237 B.n467 B.n466 585
R238 B.n465 B.n464 585
R239 B.n462 B.n461 585
R240 B.n460 B.n459 585
R241 B.n458 B.n457 585
R242 B.n456 B.n455 585
R243 B.n454 B.n453 585
R244 B.n452 B.n451 585
R245 B.n450 B.n449 585
R246 B.n448 B.n447 585
R247 B.n446 B.n445 585
R248 B.n444 B.n443 585
R249 B.n442 B.n441 585
R250 B.n440 B.n439 585
R251 B.n438 B.n437 585
R252 B.n436 B.n435 585
R253 B.n434 B.n433 585
R254 B.n432 B.n431 585
R255 B.n430 B.n429 585
R256 B.n428 B.n427 585
R257 B.n426 B.n425 585
R258 B.n424 B.n423 585
R259 B.n422 B.n421 585
R260 B.n420 B.n419 585
R261 B.n418 B.n417 585
R262 B.n416 B.n415 585
R263 B.n414 B.n413 585
R264 B.n412 B.n411 585
R265 B.n410 B.n409 585
R266 B.n408 B.n407 585
R267 B.n406 B.n405 585
R268 B.n404 B.n403 585
R269 B.n402 B.n401 585
R270 B.n400 B.n399 585
R271 B.n398 B.n397 585
R272 B.n396 B.n395 585
R273 B.n394 B.n393 585
R274 B.n392 B.n391 585
R275 B.n390 B.n389 585
R276 B.n388 B.n387 585
R277 B.n386 B.n385 585
R278 B.n384 B.n383 585
R279 B.n382 B.n381 585
R280 B.n380 B.n379 585
R281 B.n378 B.n377 585
R282 B.n376 B.n375 585
R283 B.n374 B.n373 585
R284 B.n372 B.n366 585
R285 B.n572 B.n366 585
R286 B.n576 B.n314 585
R287 B.n314 B.n313 585
R288 B.n578 B.n577 585
R289 B.n579 B.n578 585
R290 B.n308 B.n307 585
R291 B.n309 B.n308 585
R292 B.n587 B.n586 585
R293 B.n586 B.n585 585
R294 B.n588 B.n306 585
R295 B.n306 B.n305 585
R296 B.n590 B.n589 585
R297 B.n591 B.n590 585
R298 B.n300 B.n299 585
R299 B.n301 B.n300 585
R300 B.n599 B.n598 585
R301 B.n598 B.n597 585
R302 B.n600 B.n298 585
R303 B.n298 B.n297 585
R304 B.n602 B.n601 585
R305 B.n603 B.n602 585
R306 B.n292 B.n291 585
R307 B.n293 B.n292 585
R308 B.n612 B.n611 585
R309 B.n611 B.n610 585
R310 B.n613 B.n290 585
R311 B.n290 B.n289 585
R312 B.n615 B.n614 585
R313 B.n616 B.n615 585
R314 B.n2 B.n0 585
R315 B.n4 B.n2 585
R316 B.n3 B.n1 585
R317 B.n674 B.n3 585
R318 B.n672 B.n671 585
R319 B.n673 B.n672 585
R320 B.n670 B.n9 585
R321 B.n9 B.n8 585
R322 B.n669 B.n668 585
R323 B.n668 B.n667 585
R324 B.n11 B.n10 585
R325 B.n666 B.n11 585
R326 B.n664 B.n663 585
R327 B.n665 B.n664 585
R328 B.n662 B.n16 585
R329 B.n16 B.n15 585
R330 B.n661 B.n660 585
R331 B.n660 B.n659 585
R332 B.n18 B.n17 585
R333 B.n658 B.n18 585
R334 B.n656 B.n655 585
R335 B.n657 B.n656 585
R336 B.n654 B.n23 585
R337 B.n23 B.n22 585
R338 B.n653 B.n652 585
R339 B.n652 B.n651 585
R340 B.n25 B.n24 585
R341 B.n650 B.n25 585
R342 B.n648 B.n647 585
R343 B.n649 B.n648 585
R344 B.n646 B.n30 585
R345 B.n30 B.n29 585
R346 B.n677 B.n676 585
R347 B.n676 B.n675 585
R348 B.n574 B.n314 530.939
R349 B.n644 B.n30 530.939
R350 B.n366 B.n312 530.939
R351 B.n640 B.n83 530.939
R352 B.n642 B.n641 256.663
R353 B.n642 B.n81 256.663
R354 B.n642 B.n80 256.663
R355 B.n642 B.n79 256.663
R356 B.n642 B.n78 256.663
R357 B.n642 B.n77 256.663
R358 B.n642 B.n76 256.663
R359 B.n642 B.n75 256.663
R360 B.n642 B.n74 256.663
R361 B.n642 B.n73 256.663
R362 B.n642 B.n72 256.663
R363 B.n642 B.n71 256.663
R364 B.n642 B.n70 256.663
R365 B.n642 B.n69 256.663
R366 B.n642 B.n68 256.663
R367 B.n642 B.n67 256.663
R368 B.n642 B.n66 256.663
R369 B.n642 B.n65 256.663
R370 B.n642 B.n64 256.663
R371 B.n642 B.n63 256.663
R372 B.n642 B.n62 256.663
R373 B.n642 B.n61 256.663
R374 B.n642 B.n60 256.663
R375 B.n642 B.n59 256.663
R376 B.n642 B.n58 256.663
R377 B.n642 B.n57 256.663
R378 B.n642 B.n56 256.663
R379 B.n642 B.n55 256.663
R380 B.n642 B.n54 256.663
R381 B.n642 B.n53 256.663
R382 B.n642 B.n52 256.663
R383 B.n642 B.n51 256.663
R384 B.n642 B.n50 256.663
R385 B.n642 B.n49 256.663
R386 B.n642 B.n48 256.663
R387 B.n642 B.n47 256.663
R388 B.n642 B.n46 256.663
R389 B.n642 B.n45 256.663
R390 B.n642 B.n44 256.663
R391 B.n642 B.n43 256.663
R392 B.n642 B.n42 256.663
R393 B.n642 B.n41 256.663
R394 B.n642 B.n40 256.663
R395 B.n642 B.n39 256.663
R396 B.n642 B.n38 256.663
R397 B.n642 B.n37 256.663
R398 B.n642 B.n36 256.663
R399 B.n642 B.n35 256.663
R400 B.n642 B.n34 256.663
R401 B.n642 B.n33 256.663
R402 B.n643 B.n642 256.663
R403 B.n573 B.n572 256.663
R404 B.n572 B.n317 256.663
R405 B.n572 B.n318 256.663
R406 B.n572 B.n319 256.663
R407 B.n572 B.n320 256.663
R408 B.n572 B.n321 256.663
R409 B.n572 B.n322 256.663
R410 B.n572 B.n323 256.663
R411 B.n572 B.n324 256.663
R412 B.n572 B.n325 256.663
R413 B.n572 B.n326 256.663
R414 B.n572 B.n327 256.663
R415 B.n572 B.n328 256.663
R416 B.n572 B.n329 256.663
R417 B.n572 B.n330 256.663
R418 B.n572 B.n331 256.663
R419 B.n572 B.n332 256.663
R420 B.n572 B.n333 256.663
R421 B.n572 B.n334 256.663
R422 B.n572 B.n335 256.663
R423 B.n572 B.n336 256.663
R424 B.n572 B.n337 256.663
R425 B.n572 B.n338 256.663
R426 B.n572 B.n339 256.663
R427 B.n572 B.n340 256.663
R428 B.n572 B.n341 256.663
R429 B.n572 B.n342 256.663
R430 B.n572 B.n343 256.663
R431 B.n572 B.n344 256.663
R432 B.n572 B.n345 256.663
R433 B.n572 B.n346 256.663
R434 B.n572 B.n347 256.663
R435 B.n572 B.n348 256.663
R436 B.n572 B.n349 256.663
R437 B.n572 B.n350 256.663
R438 B.n572 B.n351 256.663
R439 B.n572 B.n352 256.663
R440 B.n572 B.n353 256.663
R441 B.n572 B.n354 256.663
R442 B.n572 B.n355 256.663
R443 B.n572 B.n356 256.663
R444 B.n572 B.n357 256.663
R445 B.n572 B.n358 256.663
R446 B.n572 B.n359 256.663
R447 B.n572 B.n360 256.663
R448 B.n572 B.n361 256.663
R449 B.n572 B.n362 256.663
R450 B.n572 B.n363 256.663
R451 B.n572 B.n364 256.663
R452 B.n572 B.n365 256.663
R453 B.n578 B.n314 163.367
R454 B.n578 B.n308 163.367
R455 B.n586 B.n308 163.367
R456 B.n586 B.n306 163.367
R457 B.n590 B.n306 163.367
R458 B.n590 B.n300 163.367
R459 B.n598 B.n300 163.367
R460 B.n598 B.n298 163.367
R461 B.n602 B.n298 163.367
R462 B.n602 B.n292 163.367
R463 B.n611 B.n292 163.367
R464 B.n611 B.n290 163.367
R465 B.n615 B.n290 163.367
R466 B.n615 B.n2 163.367
R467 B.n676 B.n2 163.367
R468 B.n676 B.n3 163.367
R469 B.n672 B.n3 163.367
R470 B.n672 B.n9 163.367
R471 B.n668 B.n9 163.367
R472 B.n668 B.n11 163.367
R473 B.n664 B.n11 163.367
R474 B.n664 B.n16 163.367
R475 B.n660 B.n16 163.367
R476 B.n660 B.n18 163.367
R477 B.n656 B.n18 163.367
R478 B.n656 B.n23 163.367
R479 B.n652 B.n23 163.367
R480 B.n652 B.n25 163.367
R481 B.n648 B.n25 163.367
R482 B.n648 B.n30 163.367
R483 B.n571 B.n316 163.367
R484 B.n571 B.n367 163.367
R485 B.n567 B.n566 163.367
R486 B.n563 B.n562 163.367
R487 B.n559 B.n558 163.367
R488 B.n555 B.n554 163.367
R489 B.n551 B.n550 163.367
R490 B.n547 B.n546 163.367
R491 B.n543 B.n542 163.367
R492 B.n539 B.n538 163.367
R493 B.n535 B.n534 163.367
R494 B.n531 B.n530 163.367
R495 B.n527 B.n526 163.367
R496 B.n523 B.n522 163.367
R497 B.n519 B.n518 163.367
R498 B.n515 B.n514 163.367
R499 B.n511 B.n510 163.367
R500 B.n507 B.n506 163.367
R501 B.n503 B.n502 163.367
R502 B.n499 B.n498 163.367
R503 B.n495 B.n494 163.367
R504 B.n491 B.n490 163.367
R505 B.n487 B.n486 163.367
R506 B.n482 B.n481 163.367
R507 B.n478 B.n477 163.367
R508 B.n474 B.n473 163.367
R509 B.n470 B.n469 163.367
R510 B.n466 B.n465 163.367
R511 B.n461 B.n460 163.367
R512 B.n457 B.n456 163.367
R513 B.n453 B.n452 163.367
R514 B.n449 B.n448 163.367
R515 B.n445 B.n444 163.367
R516 B.n441 B.n440 163.367
R517 B.n437 B.n436 163.367
R518 B.n433 B.n432 163.367
R519 B.n429 B.n428 163.367
R520 B.n425 B.n424 163.367
R521 B.n421 B.n420 163.367
R522 B.n417 B.n416 163.367
R523 B.n413 B.n412 163.367
R524 B.n409 B.n408 163.367
R525 B.n405 B.n404 163.367
R526 B.n401 B.n400 163.367
R527 B.n397 B.n396 163.367
R528 B.n393 B.n392 163.367
R529 B.n389 B.n388 163.367
R530 B.n385 B.n384 163.367
R531 B.n381 B.n380 163.367
R532 B.n377 B.n376 163.367
R533 B.n373 B.n366 163.367
R534 B.n580 B.n312 163.367
R535 B.n580 B.n310 163.367
R536 B.n584 B.n310 163.367
R537 B.n584 B.n304 163.367
R538 B.n592 B.n304 163.367
R539 B.n592 B.n302 163.367
R540 B.n596 B.n302 163.367
R541 B.n596 B.n296 163.367
R542 B.n604 B.n296 163.367
R543 B.n604 B.n294 163.367
R544 B.n609 B.n294 163.367
R545 B.n609 B.n288 163.367
R546 B.n617 B.n288 163.367
R547 B.n618 B.n617 163.367
R548 B.n618 B.n5 163.367
R549 B.n6 B.n5 163.367
R550 B.n7 B.n6 163.367
R551 B.n623 B.n7 163.367
R552 B.n623 B.n12 163.367
R553 B.n13 B.n12 163.367
R554 B.n14 B.n13 163.367
R555 B.n628 B.n14 163.367
R556 B.n628 B.n19 163.367
R557 B.n20 B.n19 163.367
R558 B.n21 B.n20 163.367
R559 B.n633 B.n21 163.367
R560 B.n633 B.n26 163.367
R561 B.n27 B.n26 163.367
R562 B.n28 B.n27 163.367
R563 B.n83 B.n28 163.367
R564 B.n90 B.n32 163.367
R565 B.n94 B.n93 163.367
R566 B.n98 B.n97 163.367
R567 B.n102 B.n101 163.367
R568 B.n106 B.n105 163.367
R569 B.n110 B.n109 163.367
R570 B.n114 B.n113 163.367
R571 B.n118 B.n117 163.367
R572 B.n122 B.n121 163.367
R573 B.n126 B.n125 163.367
R574 B.n130 B.n129 163.367
R575 B.n134 B.n133 163.367
R576 B.n138 B.n137 163.367
R577 B.n142 B.n141 163.367
R578 B.n146 B.n145 163.367
R579 B.n150 B.n149 163.367
R580 B.n154 B.n153 163.367
R581 B.n158 B.n157 163.367
R582 B.n162 B.n161 163.367
R583 B.n166 B.n165 163.367
R584 B.n170 B.n169 163.367
R585 B.n174 B.n173 163.367
R586 B.n178 B.n177 163.367
R587 B.n182 B.n181 163.367
R588 B.n186 B.n185 163.367
R589 B.n190 B.n189 163.367
R590 B.n194 B.n193 163.367
R591 B.n198 B.n197 163.367
R592 B.n202 B.n201 163.367
R593 B.n206 B.n205 163.367
R594 B.n210 B.n209 163.367
R595 B.n214 B.n213 163.367
R596 B.n218 B.n217 163.367
R597 B.n222 B.n221 163.367
R598 B.n226 B.n225 163.367
R599 B.n230 B.n229 163.367
R600 B.n234 B.n233 163.367
R601 B.n238 B.n237 163.367
R602 B.n242 B.n241 163.367
R603 B.n246 B.n245 163.367
R604 B.n250 B.n249 163.367
R605 B.n254 B.n253 163.367
R606 B.n258 B.n257 163.367
R607 B.n262 B.n261 163.367
R608 B.n266 B.n265 163.367
R609 B.n270 B.n269 163.367
R610 B.n274 B.n273 163.367
R611 B.n278 B.n277 163.367
R612 B.n282 B.n281 163.367
R613 B.n284 B.n82 163.367
R614 B.n370 B.t15 90.4821
R615 B.n84 B.t8 90.4821
R616 B.n368 B.t5 90.4643
R617 B.n87 B.t11 90.4643
R618 B.n574 B.n573 71.676
R619 B.n367 B.n317 71.676
R620 B.n566 B.n318 71.676
R621 B.n562 B.n319 71.676
R622 B.n558 B.n320 71.676
R623 B.n554 B.n321 71.676
R624 B.n550 B.n322 71.676
R625 B.n546 B.n323 71.676
R626 B.n542 B.n324 71.676
R627 B.n538 B.n325 71.676
R628 B.n534 B.n326 71.676
R629 B.n530 B.n327 71.676
R630 B.n526 B.n328 71.676
R631 B.n522 B.n329 71.676
R632 B.n518 B.n330 71.676
R633 B.n514 B.n331 71.676
R634 B.n510 B.n332 71.676
R635 B.n506 B.n333 71.676
R636 B.n502 B.n334 71.676
R637 B.n498 B.n335 71.676
R638 B.n494 B.n336 71.676
R639 B.n490 B.n337 71.676
R640 B.n486 B.n338 71.676
R641 B.n481 B.n339 71.676
R642 B.n477 B.n340 71.676
R643 B.n473 B.n341 71.676
R644 B.n469 B.n342 71.676
R645 B.n465 B.n343 71.676
R646 B.n460 B.n344 71.676
R647 B.n456 B.n345 71.676
R648 B.n452 B.n346 71.676
R649 B.n448 B.n347 71.676
R650 B.n444 B.n348 71.676
R651 B.n440 B.n349 71.676
R652 B.n436 B.n350 71.676
R653 B.n432 B.n351 71.676
R654 B.n428 B.n352 71.676
R655 B.n424 B.n353 71.676
R656 B.n420 B.n354 71.676
R657 B.n416 B.n355 71.676
R658 B.n412 B.n356 71.676
R659 B.n408 B.n357 71.676
R660 B.n404 B.n358 71.676
R661 B.n400 B.n359 71.676
R662 B.n396 B.n360 71.676
R663 B.n392 B.n361 71.676
R664 B.n388 B.n362 71.676
R665 B.n384 B.n363 71.676
R666 B.n380 B.n364 71.676
R667 B.n376 B.n365 71.676
R668 B.n644 B.n643 71.676
R669 B.n90 B.n33 71.676
R670 B.n94 B.n34 71.676
R671 B.n98 B.n35 71.676
R672 B.n102 B.n36 71.676
R673 B.n106 B.n37 71.676
R674 B.n110 B.n38 71.676
R675 B.n114 B.n39 71.676
R676 B.n118 B.n40 71.676
R677 B.n122 B.n41 71.676
R678 B.n126 B.n42 71.676
R679 B.n130 B.n43 71.676
R680 B.n134 B.n44 71.676
R681 B.n138 B.n45 71.676
R682 B.n142 B.n46 71.676
R683 B.n146 B.n47 71.676
R684 B.n150 B.n48 71.676
R685 B.n154 B.n49 71.676
R686 B.n158 B.n50 71.676
R687 B.n162 B.n51 71.676
R688 B.n166 B.n52 71.676
R689 B.n170 B.n53 71.676
R690 B.n174 B.n54 71.676
R691 B.n178 B.n55 71.676
R692 B.n182 B.n56 71.676
R693 B.n186 B.n57 71.676
R694 B.n190 B.n58 71.676
R695 B.n194 B.n59 71.676
R696 B.n198 B.n60 71.676
R697 B.n202 B.n61 71.676
R698 B.n206 B.n62 71.676
R699 B.n210 B.n63 71.676
R700 B.n214 B.n64 71.676
R701 B.n218 B.n65 71.676
R702 B.n222 B.n66 71.676
R703 B.n226 B.n67 71.676
R704 B.n230 B.n68 71.676
R705 B.n234 B.n69 71.676
R706 B.n238 B.n70 71.676
R707 B.n242 B.n71 71.676
R708 B.n246 B.n72 71.676
R709 B.n250 B.n73 71.676
R710 B.n254 B.n74 71.676
R711 B.n258 B.n75 71.676
R712 B.n262 B.n76 71.676
R713 B.n266 B.n77 71.676
R714 B.n270 B.n78 71.676
R715 B.n274 B.n79 71.676
R716 B.n278 B.n80 71.676
R717 B.n282 B.n81 71.676
R718 B.n641 B.n82 71.676
R719 B.n641 B.n640 71.676
R720 B.n284 B.n81 71.676
R721 B.n281 B.n80 71.676
R722 B.n277 B.n79 71.676
R723 B.n273 B.n78 71.676
R724 B.n269 B.n77 71.676
R725 B.n265 B.n76 71.676
R726 B.n261 B.n75 71.676
R727 B.n257 B.n74 71.676
R728 B.n253 B.n73 71.676
R729 B.n249 B.n72 71.676
R730 B.n245 B.n71 71.676
R731 B.n241 B.n70 71.676
R732 B.n237 B.n69 71.676
R733 B.n233 B.n68 71.676
R734 B.n229 B.n67 71.676
R735 B.n225 B.n66 71.676
R736 B.n221 B.n65 71.676
R737 B.n217 B.n64 71.676
R738 B.n213 B.n63 71.676
R739 B.n209 B.n62 71.676
R740 B.n205 B.n61 71.676
R741 B.n201 B.n60 71.676
R742 B.n197 B.n59 71.676
R743 B.n193 B.n58 71.676
R744 B.n189 B.n57 71.676
R745 B.n185 B.n56 71.676
R746 B.n181 B.n55 71.676
R747 B.n177 B.n54 71.676
R748 B.n173 B.n53 71.676
R749 B.n169 B.n52 71.676
R750 B.n165 B.n51 71.676
R751 B.n161 B.n50 71.676
R752 B.n157 B.n49 71.676
R753 B.n153 B.n48 71.676
R754 B.n149 B.n47 71.676
R755 B.n145 B.n46 71.676
R756 B.n141 B.n45 71.676
R757 B.n137 B.n44 71.676
R758 B.n133 B.n43 71.676
R759 B.n129 B.n42 71.676
R760 B.n125 B.n41 71.676
R761 B.n121 B.n40 71.676
R762 B.n117 B.n39 71.676
R763 B.n113 B.n38 71.676
R764 B.n109 B.n37 71.676
R765 B.n105 B.n36 71.676
R766 B.n101 B.n35 71.676
R767 B.n97 B.n34 71.676
R768 B.n93 B.n33 71.676
R769 B.n643 B.n32 71.676
R770 B.n573 B.n316 71.676
R771 B.n567 B.n317 71.676
R772 B.n563 B.n318 71.676
R773 B.n559 B.n319 71.676
R774 B.n555 B.n320 71.676
R775 B.n551 B.n321 71.676
R776 B.n547 B.n322 71.676
R777 B.n543 B.n323 71.676
R778 B.n539 B.n324 71.676
R779 B.n535 B.n325 71.676
R780 B.n531 B.n326 71.676
R781 B.n527 B.n327 71.676
R782 B.n523 B.n328 71.676
R783 B.n519 B.n329 71.676
R784 B.n515 B.n330 71.676
R785 B.n511 B.n331 71.676
R786 B.n507 B.n332 71.676
R787 B.n503 B.n333 71.676
R788 B.n499 B.n334 71.676
R789 B.n495 B.n335 71.676
R790 B.n491 B.n336 71.676
R791 B.n487 B.n337 71.676
R792 B.n482 B.n338 71.676
R793 B.n478 B.n339 71.676
R794 B.n474 B.n340 71.676
R795 B.n470 B.n341 71.676
R796 B.n466 B.n342 71.676
R797 B.n461 B.n343 71.676
R798 B.n457 B.n344 71.676
R799 B.n453 B.n345 71.676
R800 B.n449 B.n346 71.676
R801 B.n445 B.n347 71.676
R802 B.n441 B.n348 71.676
R803 B.n437 B.n349 71.676
R804 B.n433 B.n350 71.676
R805 B.n429 B.n351 71.676
R806 B.n425 B.n352 71.676
R807 B.n421 B.n353 71.676
R808 B.n417 B.n354 71.676
R809 B.n413 B.n355 71.676
R810 B.n409 B.n356 71.676
R811 B.n405 B.n357 71.676
R812 B.n401 B.n358 71.676
R813 B.n397 B.n359 71.676
R814 B.n393 B.n360 71.676
R815 B.n389 B.n361 71.676
R816 B.n385 B.n362 71.676
R817 B.n381 B.n363 71.676
R818 B.n377 B.n364 71.676
R819 B.n373 B.n365 71.676
R820 B.n572 B.n313 71.5689
R821 B.n642 B.n29 71.5689
R822 B.n371 B.t14 67.7911
R823 B.n85 B.t9 67.7911
R824 B.n369 B.t4 67.7734
R825 B.n88 B.t12 67.7734
R826 B.n463 B.n371 59.5399
R827 B.n484 B.n369 59.5399
R828 B.n89 B.n88 59.5399
R829 B.n86 B.n85 59.5399
R830 B.n579 B.n313 39.5668
R831 B.n579 B.n309 39.5668
R832 B.n585 B.n309 39.5668
R833 B.n585 B.n305 39.5668
R834 B.n591 B.n305 39.5668
R835 B.n597 B.n301 39.5668
R836 B.n597 B.n297 39.5668
R837 B.n603 B.n297 39.5668
R838 B.n603 B.n293 39.5668
R839 B.n610 B.n293 39.5668
R840 B.n616 B.n289 39.5668
R841 B.n616 B.n4 39.5668
R842 B.n675 B.n4 39.5668
R843 B.n675 B.n674 39.5668
R844 B.n674 B.n673 39.5668
R845 B.n673 B.n8 39.5668
R846 B.n667 B.n666 39.5668
R847 B.n666 B.n665 39.5668
R848 B.n665 B.n15 39.5668
R849 B.n659 B.n15 39.5668
R850 B.n659 B.n658 39.5668
R851 B.n657 B.n22 39.5668
R852 B.n651 B.n22 39.5668
R853 B.n651 B.n650 39.5668
R854 B.n650 B.n649 39.5668
R855 B.n649 B.n29 39.5668
R856 B.t3 B.n301 38.403
R857 B.n658 B.t7 38.403
R858 B.n646 B.n645 34.4981
R859 B.n639 B.n638 34.4981
R860 B.n372 B.n311 34.4981
R861 B.n576 B.n575 34.4981
R862 B.n610 B.t1 26.7659
R863 B.n667 B.t0 26.7659
R864 B.n371 B.n370 22.6914
R865 B.n369 B.n368 22.6914
R866 B.n88 B.n87 22.6914
R867 B.n85 B.n84 22.6914
R868 B B.n677 18.0485
R869 B.t1 B.n289 12.8013
R870 B.t0 B.n8 12.8013
R871 B.n645 B.n31 10.6151
R872 B.n91 B.n31 10.6151
R873 B.n92 B.n91 10.6151
R874 B.n95 B.n92 10.6151
R875 B.n96 B.n95 10.6151
R876 B.n99 B.n96 10.6151
R877 B.n100 B.n99 10.6151
R878 B.n103 B.n100 10.6151
R879 B.n104 B.n103 10.6151
R880 B.n107 B.n104 10.6151
R881 B.n108 B.n107 10.6151
R882 B.n111 B.n108 10.6151
R883 B.n112 B.n111 10.6151
R884 B.n115 B.n112 10.6151
R885 B.n116 B.n115 10.6151
R886 B.n119 B.n116 10.6151
R887 B.n120 B.n119 10.6151
R888 B.n123 B.n120 10.6151
R889 B.n124 B.n123 10.6151
R890 B.n127 B.n124 10.6151
R891 B.n128 B.n127 10.6151
R892 B.n131 B.n128 10.6151
R893 B.n132 B.n131 10.6151
R894 B.n135 B.n132 10.6151
R895 B.n136 B.n135 10.6151
R896 B.n139 B.n136 10.6151
R897 B.n140 B.n139 10.6151
R898 B.n143 B.n140 10.6151
R899 B.n144 B.n143 10.6151
R900 B.n147 B.n144 10.6151
R901 B.n148 B.n147 10.6151
R902 B.n151 B.n148 10.6151
R903 B.n152 B.n151 10.6151
R904 B.n155 B.n152 10.6151
R905 B.n156 B.n155 10.6151
R906 B.n159 B.n156 10.6151
R907 B.n160 B.n159 10.6151
R908 B.n163 B.n160 10.6151
R909 B.n164 B.n163 10.6151
R910 B.n167 B.n164 10.6151
R911 B.n168 B.n167 10.6151
R912 B.n171 B.n168 10.6151
R913 B.n172 B.n171 10.6151
R914 B.n175 B.n172 10.6151
R915 B.n176 B.n175 10.6151
R916 B.n180 B.n179 10.6151
R917 B.n183 B.n180 10.6151
R918 B.n184 B.n183 10.6151
R919 B.n187 B.n184 10.6151
R920 B.n188 B.n187 10.6151
R921 B.n191 B.n188 10.6151
R922 B.n192 B.n191 10.6151
R923 B.n195 B.n192 10.6151
R924 B.n196 B.n195 10.6151
R925 B.n200 B.n199 10.6151
R926 B.n203 B.n200 10.6151
R927 B.n204 B.n203 10.6151
R928 B.n207 B.n204 10.6151
R929 B.n208 B.n207 10.6151
R930 B.n211 B.n208 10.6151
R931 B.n212 B.n211 10.6151
R932 B.n215 B.n212 10.6151
R933 B.n216 B.n215 10.6151
R934 B.n219 B.n216 10.6151
R935 B.n220 B.n219 10.6151
R936 B.n223 B.n220 10.6151
R937 B.n224 B.n223 10.6151
R938 B.n227 B.n224 10.6151
R939 B.n228 B.n227 10.6151
R940 B.n231 B.n228 10.6151
R941 B.n232 B.n231 10.6151
R942 B.n235 B.n232 10.6151
R943 B.n236 B.n235 10.6151
R944 B.n239 B.n236 10.6151
R945 B.n240 B.n239 10.6151
R946 B.n243 B.n240 10.6151
R947 B.n244 B.n243 10.6151
R948 B.n247 B.n244 10.6151
R949 B.n248 B.n247 10.6151
R950 B.n251 B.n248 10.6151
R951 B.n252 B.n251 10.6151
R952 B.n255 B.n252 10.6151
R953 B.n256 B.n255 10.6151
R954 B.n259 B.n256 10.6151
R955 B.n260 B.n259 10.6151
R956 B.n263 B.n260 10.6151
R957 B.n264 B.n263 10.6151
R958 B.n267 B.n264 10.6151
R959 B.n268 B.n267 10.6151
R960 B.n271 B.n268 10.6151
R961 B.n272 B.n271 10.6151
R962 B.n275 B.n272 10.6151
R963 B.n276 B.n275 10.6151
R964 B.n279 B.n276 10.6151
R965 B.n280 B.n279 10.6151
R966 B.n283 B.n280 10.6151
R967 B.n285 B.n283 10.6151
R968 B.n286 B.n285 10.6151
R969 B.n639 B.n286 10.6151
R970 B.n581 B.n311 10.6151
R971 B.n582 B.n581 10.6151
R972 B.n583 B.n582 10.6151
R973 B.n583 B.n303 10.6151
R974 B.n593 B.n303 10.6151
R975 B.n594 B.n593 10.6151
R976 B.n595 B.n594 10.6151
R977 B.n595 B.n295 10.6151
R978 B.n605 B.n295 10.6151
R979 B.n606 B.n605 10.6151
R980 B.n608 B.n606 10.6151
R981 B.n608 B.n607 10.6151
R982 B.n607 B.n287 10.6151
R983 B.n619 B.n287 10.6151
R984 B.n620 B.n619 10.6151
R985 B.n621 B.n620 10.6151
R986 B.n622 B.n621 10.6151
R987 B.n624 B.n622 10.6151
R988 B.n625 B.n624 10.6151
R989 B.n626 B.n625 10.6151
R990 B.n627 B.n626 10.6151
R991 B.n629 B.n627 10.6151
R992 B.n630 B.n629 10.6151
R993 B.n631 B.n630 10.6151
R994 B.n632 B.n631 10.6151
R995 B.n634 B.n632 10.6151
R996 B.n635 B.n634 10.6151
R997 B.n636 B.n635 10.6151
R998 B.n637 B.n636 10.6151
R999 B.n638 B.n637 10.6151
R1000 B.n575 B.n315 10.6151
R1001 B.n570 B.n315 10.6151
R1002 B.n570 B.n569 10.6151
R1003 B.n569 B.n568 10.6151
R1004 B.n568 B.n565 10.6151
R1005 B.n565 B.n564 10.6151
R1006 B.n564 B.n561 10.6151
R1007 B.n561 B.n560 10.6151
R1008 B.n560 B.n557 10.6151
R1009 B.n557 B.n556 10.6151
R1010 B.n556 B.n553 10.6151
R1011 B.n553 B.n552 10.6151
R1012 B.n552 B.n549 10.6151
R1013 B.n549 B.n548 10.6151
R1014 B.n548 B.n545 10.6151
R1015 B.n545 B.n544 10.6151
R1016 B.n544 B.n541 10.6151
R1017 B.n541 B.n540 10.6151
R1018 B.n540 B.n537 10.6151
R1019 B.n537 B.n536 10.6151
R1020 B.n536 B.n533 10.6151
R1021 B.n533 B.n532 10.6151
R1022 B.n532 B.n529 10.6151
R1023 B.n529 B.n528 10.6151
R1024 B.n528 B.n525 10.6151
R1025 B.n525 B.n524 10.6151
R1026 B.n524 B.n521 10.6151
R1027 B.n521 B.n520 10.6151
R1028 B.n520 B.n517 10.6151
R1029 B.n517 B.n516 10.6151
R1030 B.n516 B.n513 10.6151
R1031 B.n513 B.n512 10.6151
R1032 B.n512 B.n509 10.6151
R1033 B.n509 B.n508 10.6151
R1034 B.n508 B.n505 10.6151
R1035 B.n505 B.n504 10.6151
R1036 B.n504 B.n501 10.6151
R1037 B.n501 B.n500 10.6151
R1038 B.n500 B.n497 10.6151
R1039 B.n497 B.n496 10.6151
R1040 B.n496 B.n493 10.6151
R1041 B.n493 B.n492 10.6151
R1042 B.n492 B.n489 10.6151
R1043 B.n489 B.n488 10.6151
R1044 B.n488 B.n485 10.6151
R1045 B.n483 B.n480 10.6151
R1046 B.n480 B.n479 10.6151
R1047 B.n479 B.n476 10.6151
R1048 B.n476 B.n475 10.6151
R1049 B.n475 B.n472 10.6151
R1050 B.n472 B.n471 10.6151
R1051 B.n471 B.n468 10.6151
R1052 B.n468 B.n467 10.6151
R1053 B.n467 B.n464 10.6151
R1054 B.n462 B.n459 10.6151
R1055 B.n459 B.n458 10.6151
R1056 B.n458 B.n455 10.6151
R1057 B.n455 B.n454 10.6151
R1058 B.n454 B.n451 10.6151
R1059 B.n451 B.n450 10.6151
R1060 B.n450 B.n447 10.6151
R1061 B.n447 B.n446 10.6151
R1062 B.n446 B.n443 10.6151
R1063 B.n443 B.n442 10.6151
R1064 B.n442 B.n439 10.6151
R1065 B.n439 B.n438 10.6151
R1066 B.n438 B.n435 10.6151
R1067 B.n435 B.n434 10.6151
R1068 B.n434 B.n431 10.6151
R1069 B.n431 B.n430 10.6151
R1070 B.n430 B.n427 10.6151
R1071 B.n427 B.n426 10.6151
R1072 B.n426 B.n423 10.6151
R1073 B.n423 B.n422 10.6151
R1074 B.n422 B.n419 10.6151
R1075 B.n419 B.n418 10.6151
R1076 B.n418 B.n415 10.6151
R1077 B.n415 B.n414 10.6151
R1078 B.n414 B.n411 10.6151
R1079 B.n411 B.n410 10.6151
R1080 B.n410 B.n407 10.6151
R1081 B.n407 B.n406 10.6151
R1082 B.n406 B.n403 10.6151
R1083 B.n403 B.n402 10.6151
R1084 B.n402 B.n399 10.6151
R1085 B.n399 B.n398 10.6151
R1086 B.n398 B.n395 10.6151
R1087 B.n395 B.n394 10.6151
R1088 B.n394 B.n391 10.6151
R1089 B.n391 B.n390 10.6151
R1090 B.n390 B.n387 10.6151
R1091 B.n387 B.n386 10.6151
R1092 B.n386 B.n383 10.6151
R1093 B.n383 B.n382 10.6151
R1094 B.n382 B.n379 10.6151
R1095 B.n379 B.n378 10.6151
R1096 B.n378 B.n375 10.6151
R1097 B.n375 B.n374 10.6151
R1098 B.n374 B.n372 10.6151
R1099 B.n577 B.n576 10.6151
R1100 B.n577 B.n307 10.6151
R1101 B.n587 B.n307 10.6151
R1102 B.n588 B.n587 10.6151
R1103 B.n589 B.n588 10.6151
R1104 B.n589 B.n299 10.6151
R1105 B.n599 B.n299 10.6151
R1106 B.n600 B.n599 10.6151
R1107 B.n601 B.n600 10.6151
R1108 B.n601 B.n291 10.6151
R1109 B.n612 B.n291 10.6151
R1110 B.n613 B.n612 10.6151
R1111 B.n614 B.n613 10.6151
R1112 B.n614 B.n0 10.6151
R1113 B.n671 B.n1 10.6151
R1114 B.n671 B.n670 10.6151
R1115 B.n670 B.n669 10.6151
R1116 B.n669 B.n10 10.6151
R1117 B.n663 B.n10 10.6151
R1118 B.n663 B.n662 10.6151
R1119 B.n662 B.n661 10.6151
R1120 B.n661 B.n17 10.6151
R1121 B.n655 B.n17 10.6151
R1122 B.n655 B.n654 10.6151
R1123 B.n654 B.n653 10.6151
R1124 B.n653 B.n24 10.6151
R1125 B.n647 B.n24 10.6151
R1126 B.n647 B.n646 10.6151
R1127 B.n176 B.n89 8.74196
R1128 B.n199 B.n86 8.74196
R1129 B.n485 B.n484 8.74196
R1130 B.n463 B.n462 8.74196
R1131 B.n677 B.n0 2.81026
R1132 B.n677 B.n1 2.81026
R1133 B.n179 B.n89 1.87367
R1134 B.n196 B.n86 1.87367
R1135 B.n484 B.n483 1.87367
R1136 B.n464 B.n463 1.87367
R1137 B.n591 B.t3 1.16421
R1138 B.t7 B.n657 1.16421
R1139 VP.n0 VP.t1 640.053
R1140 VP.n0 VP.t0 598.831
R1141 VP VP.n0 0.0516364
R1142 VDD1 VDD1.t1 101.695
R1143 VDD1 VDD1.t0 63.8018
C0 VTAIL VDD2 6.05322f
C1 VN VTAIL 1.81092f
C2 VP VDD1 2.47428f
C3 VP VDD2 0.261046f
C4 VDD1 VDD2 0.476243f
C5 VP VN 4.92315f
C6 VN VDD1 0.148652f
C7 VN VDD2 2.36653f
C8 VP VTAIL 1.82554f
C9 VDD1 VTAIL 6.01874f
C10 VDD2 B 4.097591f
C11 VDD1 B 7.04177f
C12 VTAIL B 7.064014f
C13 VN B 8.51563f
C14 VP B 4.306966f
C15 VDD1.t0 B 2.5506f
C16 VDD1.t1 B 3.08566f
C17 VP.t1 B 1.6876f
C18 VP.t0 B 1.55038f
C19 VP.n0 B 4.14326f
C20 VDD2.t0 B 3.08687f
C21 VDD2.t1 B 2.57246f
C22 VDD2.n0 B 2.78541f
C23 VTAIL.t3 B 1.88344f
C24 VTAIL.n0 B 1.15729f
C25 VTAIL.t0 B 1.88344f
C26 VTAIL.n1 B 1.16712f
C27 VTAIL.t2 B 1.88344f
C28 VTAIL.n2 B 1.116f
C29 VTAIL.t1 B 1.88344f
C30 VTAIL.n3 B 1.07646f
C31 VN.t1 B 1.51702f
C32 VN.t0 B 1.65422f
.ends

