* NGSPICE file created from diff_pair_sample_1309.ext - technology: sky130A

.subckt diff_pair_sample_1309 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=3.32
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=3.32
X2 B.t8 B.t6 B.t7 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=3.32
X3 VDD1.t1 VP.t0 VTAIL.t3 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=3.32
X4 B.t5 B.t3 B.t4 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=3.32
X5 B.t2 B.t0 B.t1 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=3.32
X6 VDD2.t0 VN.t1 VTAIL.t1 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=3.32
X7 VDD1.t0 VP.t1 VTAIL.t2 w_n2430_n4308# sky130_fd_pr__pfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=3.32
R0 B.n412 B.n111 585
R1 B.n411 B.n410 585
R2 B.n409 B.n112 585
R3 B.n408 B.n407 585
R4 B.n406 B.n113 585
R5 B.n405 B.n404 585
R6 B.n403 B.n114 585
R7 B.n402 B.n401 585
R8 B.n400 B.n115 585
R9 B.n399 B.n398 585
R10 B.n397 B.n116 585
R11 B.n396 B.n395 585
R12 B.n394 B.n117 585
R13 B.n393 B.n392 585
R14 B.n391 B.n118 585
R15 B.n390 B.n389 585
R16 B.n388 B.n119 585
R17 B.n387 B.n386 585
R18 B.n385 B.n120 585
R19 B.n384 B.n383 585
R20 B.n382 B.n121 585
R21 B.n381 B.n380 585
R22 B.n379 B.n122 585
R23 B.n378 B.n377 585
R24 B.n376 B.n123 585
R25 B.n375 B.n374 585
R26 B.n373 B.n124 585
R27 B.n372 B.n371 585
R28 B.n370 B.n125 585
R29 B.n369 B.n368 585
R30 B.n367 B.n126 585
R31 B.n366 B.n365 585
R32 B.n364 B.n127 585
R33 B.n363 B.n362 585
R34 B.n361 B.n128 585
R35 B.n360 B.n359 585
R36 B.n358 B.n129 585
R37 B.n357 B.n356 585
R38 B.n355 B.n130 585
R39 B.n354 B.n353 585
R40 B.n352 B.n131 585
R41 B.n351 B.n350 585
R42 B.n349 B.n132 585
R43 B.n348 B.n347 585
R44 B.n346 B.n133 585
R45 B.n345 B.n344 585
R46 B.n343 B.n134 585
R47 B.n342 B.n341 585
R48 B.n340 B.n135 585
R49 B.n339 B.n338 585
R50 B.n337 B.n136 585
R51 B.n336 B.n335 585
R52 B.n334 B.n137 585
R53 B.n333 B.n332 585
R54 B.n331 B.n138 585
R55 B.n330 B.n329 585
R56 B.n325 B.n139 585
R57 B.n324 B.n323 585
R58 B.n322 B.n140 585
R59 B.n321 B.n320 585
R60 B.n319 B.n141 585
R61 B.n318 B.n317 585
R62 B.n316 B.n142 585
R63 B.n315 B.n314 585
R64 B.n313 B.n143 585
R65 B.n311 B.n310 585
R66 B.n309 B.n146 585
R67 B.n308 B.n307 585
R68 B.n306 B.n147 585
R69 B.n305 B.n304 585
R70 B.n303 B.n148 585
R71 B.n302 B.n301 585
R72 B.n300 B.n149 585
R73 B.n299 B.n298 585
R74 B.n297 B.n150 585
R75 B.n296 B.n295 585
R76 B.n294 B.n151 585
R77 B.n293 B.n292 585
R78 B.n291 B.n152 585
R79 B.n290 B.n289 585
R80 B.n288 B.n153 585
R81 B.n287 B.n286 585
R82 B.n285 B.n154 585
R83 B.n284 B.n283 585
R84 B.n282 B.n155 585
R85 B.n281 B.n280 585
R86 B.n279 B.n156 585
R87 B.n278 B.n277 585
R88 B.n276 B.n157 585
R89 B.n275 B.n274 585
R90 B.n273 B.n158 585
R91 B.n272 B.n271 585
R92 B.n270 B.n159 585
R93 B.n269 B.n268 585
R94 B.n267 B.n160 585
R95 B.n266 B.n265 585
R96 B.n264 B.n161 585
R97 B.n263 B.n262 585
R98 B.n261 B.n162 585
R99 B.n260 B.n259 585
R100 B.n258 B.n163 585
R101 B.n257 B.n256 585
R102 B.n255 B.n164 585
R103 B.n254 B.n253 585
R104 B.n252 B.n165 585
R105 B.n251 B.n250 585
R106 B.n249 B.n166 585
R107 B.n248 B.n247 585
R108 B.n246 B.n167 585
R109 B.n245 B.n244 585
R110 B.n243 B.n168 585
R111 B.n242 B.n241 585
R112 B.n240 B.n169 585
R113 B.n239 B.n238 585
R114 B.n237 B.n170 585
R115 B.n236 B.n235 585
R116 B.n234 B.n171 585
R117 B.n233 B.n232 585
R118 B.n231 B.n172 585
R119 B.n230 B.n229 585
R120 B.n414 B.n413 585
R121 B.n415 B.n110 585
R122 B.n417 B.n416 585
R123 B.n418 B.n109 585
R124 B.n420 B.n419 585
R125 B.n421 B.n108 585
R126 B.n423 B.n422 585
R127 B.n424 B.n107 585
R128 B.n426 B.n425 585
R129 B.n427 B.n106 585
R130 B.n429 B.n428 585
R131 B.n430 B.n105 585
R132 B.n432 B.n431 585
R133 B.n433 B.n104 585
R134 B.n435 B.n434 585
R135 B.n436 B.n103 585
R136 B.n438 B.n437 585
R137 B.n439 B.n102 585
R138 B.n441 B.n440 585
R139 B.n442 B.n101 585
R140 B.n444 B.n443 585
R141 B.n445 B.n100 585
R142 B.n447 B.n446 585
R143 B.n448 B.n99 585
R144 B.n450 B.n449 585
R145 B.n451 B.n98 585
R146 B.n453 B.n452 585
R147 B.n454 B.n97 585
R148 B.n456 B.n455 585
R149 B.n457 B.n96 585
R150 B.n459 B.n458 585
R151 B.n460 B.n95 585
R152 B.n462 B.n461 585
R153 B.n463 B.n94 585
R154 B.n465 B.n464 585
R155 B.n466 B.n93 585
R156 B.n468 B.n467 585
R157 B.n469 B.n92 585
R158 B.n471 B.n470 585
R159 B.n472 B.n91 585
R160 B.n474 B.n473 585
R161 B.n475 B.n90 585
R162 B.n477 B.n476 585
R163 B.n478 B.n89 585
R164 B.n480 B.n479 585
R165 B.n481 B.n88 585
R166 B.n483 B.n482 585
R167 B.n484 B.n87 585
R168 B.n486 B.n485 585
R169 B.n487 B.n86 585
R170 B.n489 B.n488 585
R171 B.n490 B.n85 585
R172 B.n492 B.n491 585
R173 B.n493 B.n84 585
R174 B.n495 B.n494 585
R175 B.n496 B.n83 585
R176 B.n498 B.n497 585
R177 B.n499 B.n82 585
R178 B.n501 B.n500 585
R179 B.n502 B.n81 585
R180 B.n684 B.n683 585
R181 B.n682 B.n17 585
R182 B.n681 B.n680 585
R183 B.n679 B.n18 585
R184 B.n678 B.n677 585
R185 B.n676 B.n19 585
R186 B.n675 B.n674 585
R187 B.n673 B.n20 585
R188 B.n672 B.n671 585
R189 B.n670 B.n21 585
R190 B.n669 B.n668 585
R191 B.n667 B.n22 585
R192 B.n666 B.n665 585
R193 B.n664 B.n23 585
R194 B.n663 B.n662 585
R195 B.n661 B.n24 585
R196 B.n660 B.n659 585
R197 B.n658 B.n25 585
R198 B.n657 B.n656 585
R199 B.n655 B.n26 585
R200 B.n654 B.n653 585
R201 B.n652 B.n27 585
R202 B.n651 B.n650 585
R203 B.n649 B.n28 585
R204 B.n648 B.n647 585
R205 B.n646 B.n29 585
R206 B.n645 B.n644 585
R207 B.n643 B.n30 585
R208 B.n642 B.n641 585
R209 B.n640 B.n31 585
R210 B.n639 B.n638 585
R211 B.n637 B.n32 585
R212 B.n636 B.n635 585
R213 B.n634 B.n33 585
R214 B.n633 B.n632 585
R215 B.n631 B.n34 585
R216 B.n630 B.n629 585
R217 B.n628 B.n35 585
R218 B.n627 B.n626 585
R219 B.n625 B.n36 585
R220 B.n624 B.n623 585
R221 B.n622 B.n37 585
R222 B.n621 B.n620 585
R223 B.n619 B.n38 585
R224 B.n618 B.n617 585
R225 B.n616 B.n39 585
R226 B.n615 B.n614 585
R227 B.n613 B.n40 585
R228 B.n612 B.n611 585
R229 B.n610 B.n41 585
R230 B.n609 B.n608 585
R231 B.n607 B.n42 585
R232 B.n606 B.n605 585
R233 B.n604 B.n43 585
R234 B.n603 B.n602 585
R235 B.n601 B.n600 585
R236 B.n599 B.n47 585
R237 B.n598 B.n597 585
R238 B.n596 B.n48 585
R239 B.n595 B.n594 585
R240 B.n593 B.n49 585
R241 B.n592 B.n591 585
R242 B.n590 B.n50 585
R243 B.n589 B.n588 585
R244 B.n587 B.n51 585
R245 B.n585 B.n584 585
R246 B.n583 B.n54 585
R247 B.n582 B.n581 585
R248 B.n580 B.n55 585
R249 B.n579 B.n578 585
R250 B.n577 B.n56 585
R251 B.n576 B.n575 585
R252 B.n574 B.n57 585
R253 B.n573 B.n572 585
R254 B.n571 B.n58 585
R255 B.n570 B.n569 585
R256 B.n568 B.n59 585
R257 B.n567 B.n566 585
R258 B.n565 B.n60 585
R259 B.n564 B.n563 585
R260 B.n562 B.n61 585
R261 B.n561 B.n560 585
R262 B.n559 B.n62 585
R263 B.n558 B.n557 585
R264 B.n556 B.n63 585
R265 B.n555 B.n554 585
R266 B.n553 B.n64 585
R267 B.n552 B.n551 585
R268 B.n550 B.n65 585
R269 B.n549 B.n548 585
R270 B.n547 B.n66 585
R271 B.n546 B.n545 585
R272 B.n544 B.n67 585
R273 B.n543 B.n542 585
R274 B.n541 B.n68 585
R275 B.n540 B.n539 585
R276 B.n538 B.n69 585
R277 B.n537 B.n536 585
R278 B.n535 B.n70 585
R279 B.n534 B.n533 585
R280 B.n532 B.n71 585
R281 B.n531 B.n530 585
R282 B.n529 B.n72 585
R283 B.n528 B.n527 585
R284 B.n526 B.n73 585
R285 B.n525 B.n524 585
R286 B.n523 B.n74 585
R287 B.n522 B.n521 585
R288 B.n520 B.n75 585
R289 B.n519 B.n518 585
R290 B.n517 B.n76 585
R291 B.n516 B.n515 585
R292 B.n514 B.n77 585
R293 B.n513 B.n512 585
R294 B.n511 B.n78 585
R295 B.n510 B.n509 585
R296 B.n508 B.n79 585
R297 B.n507 B.n506 585
R298 B.n505 B.n80 585
R299 B.n504 B.n503 585
R300 B.n685 B.n16 585
R301 B.n687 B.n686 585
R302 B.n688 B.n15 585
R303 B.n690 B.n689 585
R304 B.n691 B.n14 585
R305 B.n693 B.n692 585
R306 B.n694 B.n13 585
R307 B.n696 B.n695 585
R308 B.n697 B.n12 585
R309 B.n699 B.n698 585
R310 B.n700 B.n11 585
R311 B.n702 B.n701 585
R312 B.n703 B.n10 585
R313 B.n705 B.n704 585
R314 B.n706 B.n9 585
R315 B.n708 B.n707 585
R316 B.n709 B.n8 585
R317 B.n711 B.n710 585
R318 B.n712 B.n7 585
R319 B.n714 B.n713 585
R320 B.n715 B.n6 585
R321 B.n717 B.n716 585
R322 B.n718 B.n5 585
R323 B.n720 B.n719 585
R324 B.n721 B.n4 585
R325 B.n723 B.n722 585
R326 B.n724 B.n3 585
R327 B.n726 B.n725 585
R328 B.n727 B.n0 585
R329 B.n2 B.n1 585
R330 B.n188 B.n187 585
R331 B.n189 B.n186 585
R332 B.n191 B.n190 585
R333 B.n192 B.n185 585
R334 B.n194 B.n193 585
R335 B.n195 B.n184 585
R336 B.n197 B.n196 585
R337 B.n198 B.n183 585
R338 B.n200 B.n199 585
R339 B.n201 B.n182 585
R340 B.n203 B.n202 585
R341 B.n204 B.n181 585
R342 B.n206 B.n205 585
R343 B.n207 B.n180 585
R344 B.n209 B.n208 585
R345 B.n210 B.n179 585
R346 B.n212 B.n211 585
R347 B.n213 B.n178 585
R348 B.n215 B.n214 585
R349 B.n216 B.n177 585
R350 B.n218 B.n217 585
R351 B.n219 B.n176 585
R352 B.n221 B.n220 585
R353 B.n222 B.n175 585
R354 B.n224 B.n223 585
R355 B.n225 B.n174 585
R356 B.n227 B.n226 585
R357 B.n228 B.n173 585
R358 B.n230 B.n173 550.159
R359 B.n414 B.n111 550.159
R360 B.n504 B.n81 550.159
R361 B.n685 B.n684 550.159
R362 B.n326 B.t7 530.889
R363 B.n52 B.t2 530.889
R364 B.n144 B.t4 530.889
R365 B.n44 B.t11 530.889
R366 B.n327 B.t8 460.101
R367 B.n53 B.t1 460.101
R368 B.n145 B.t5 460.101
R369 B.n45 B.t10 460.101
R370 B.n144 B.t3 330.151
R371 B.n326 B.t6 330.151
R372 B.n52 B.t0 330.151
R373 B.n44 B.t9 330.151
R374 B.n729 B.n728 256.663
R375 B.n728 B.n727 235.042
R376 B.n728 B.n2 235.042
R377 B.n231 B.n230 163.367
R378 B.n232 B.n231 163.367
R379 B.n232 B.n171 163.367
R380 B.n236 B.n171 163.367
R381 B.n237 B.n236 163.367
R382 B.n238 B.n237 163.367
R383 B.n238 B.n169 163.367
R384 B.n242 B.n169 163.367
R385 B.n243 B.n242 163.367
R386 B.n244 B.n243 163.367
R387 B.n244 B.n167 163.367
R388 B.n248 B.n167 163.367
R389 B.n249 B.n248 163.367
R390 B.n250 B.n249 163.367
R391 B.n250 B.n165 163.367
R392 B.n254 B.n165 163.367
R393 B.n255 B.n254 163.367
R394 B.n256 B.n255 163.367
R395 B.n256 B.n163 163.367
R396 B.n260 B.n163 163.367
R397 B.n261 B.n260 163.367
R398 B.n262 B.n261 163.367
R399 B.n262 B.n161 163.367
R400 B.n266 B.n161 163.367
R401 B.n267 B.n266 163.367
R402 B.n268 B.n267 163.367
R403 B.n268 B.n159 163.367
R404 B.n272 B.n159 163.367
R405 B.n273 B.n272 163.367
R406 B.n274 B.n273 163.367
R407 B.n274 B.n157 163.367
R408 B.n278 B.n157 163.367
R409 B.n279 B.n278 163.367
R410 B.n280 B.n279 163.367
R411 B.n280 B.n155 163.367
R412 B.n284 B.n155 163.367
R413 B.n285 B.n284 163.367
R414 B.n286 B.n285 163.367
R415 B.n286 B.n153 163.367
R416 B.n290 B.n153 163.367
R417 B.n291 B.n290 163.367
R418 B.n292 B.n291 163.367
R419 B.n292 B.n151 163.367
R420 B.n296 B.n151 163.367
R421 B.n297 B.n296 163.367
R422 B.n298 B.n297 163.367
R423 B.n298 B.n149 163.367
R424 B.n302 B.n149 163.367
R425 B.n303 B.n302 163.367
R426 B.n304 B.n303 163.367
R427 B.n304 B.n147 163.367
R428 B.n308 B.n147 163.367
R429 B.n309 B.n308 163.367
R430 B.n310 B.n309 163.367
R431 B.n310 B.n143 163.367
R432 B.n315 B.n143 163.367
R433 B.n316 B.n315 163.367
R434 B.n317 B.n316 163.367
R435 B.n317 B.n141 163.367
R436 B.n321 B.n141 163.367
R437 B.n322 B.n321 163.367
R438 B.n323 B.n322 163.367
R439 B.n323 B.n139 163.367
R440 B.n330 B.n139 163.367
R441 B.n331 B.n330 163.367
R442 B.n332 B.n331 163.367
R443 B.n332 B.n137 163.367
R444 B.n336 B.n137 163.367
R445 B.n337 B.n336 163.367
R446 B.n338 B.n337 163.367
R447 B.n338 B.n135 163.367
R448 B.n342 B.n135 163.367
R449 B.n343 B.n342 163.367
R450 B.n344 B.n343 163.367
R451 B.n344 B.n133 163.367
R452 B.n348 B.n133 163.367
R453 B.n349 B.n348 163.367
R454 B.n350 B.n349 163.367
R455 B.n350 B.n131 163.367
R456 B.n354 B.n131 163.367
R457 B.n355 B.n354 163.367
R458 B.n356 B.n355 163.367
R459 B.n356 B.n129 163.367
R460 B.n360 B.n129 163.367
R461 B.n361 B.n360 163.367
R462 B.n362 B.n361 163.367
R463 B.n362 B.n127 163.367
R464 B.n366 B.n127 163.367
R465 B.n367 B.n366 163.367
R466 B.n368 B.n367 163.367
R467 B.n368 B.n125 163.367
R468 B.n372 B.n125 163.367
R469 B.n373 B.n372 163.367
R470 B.n374 B.n373 163.367
R471 B.n374 B.n123 163.367
R472 B.n378 B.n123 163.367
R473 B.n379 B.n378 163.367
R474 B.n380 B.n379 163.367
R475 B.n380 B.n121 163.367
R476 B.n384 B.n121 163.367
R477 B.n385 B.n384 163.367
R478 B.n386 B.n385 163.367
R479 B.n386 B.n119 163.367
R480 B.n390 B.n119 163.367
R481 B.n391 B.n390 163.367
R482 B.n392 B.n391 163.367
R483 B.n392 B.n117 163.367
R484 B.n396 B.n117 163.367
R485 B.n397 B.n396 163.367
R486 B.n398 B.n397 163.367
R487 B.n398 B.n115 163.367
R488 B.n402 B.n115 163.367
R489 B.n403 B.n402 163.367
R490 B.n404 B.n403 163.367
R491 B.n404 B.n113 163.367
R492 B.n408 B.n113 163.367
R493 B.n409 B.n408 163.367
R494 B.n410 B.n409 163.367
R495 B.n410 B.n111 163.367
R496 B.n500 B.n81 163.367
R497 B.n500 B.n499 163.367
R498 B.n499 B.n498 163.367
R499 B.n498 B.n83 163.367
R500 B.n494 B.n83 163.367
R501 B.n494 B.n493 163.367
R502 B.n493 B.n492 163.367
R503 B.n492 B.n85 163.367
R504 B.n488 B.n85 163.367
R505 B.n488 B.n487 163.367
R506 B.n487 B.n486 163.367
R507 B.n486 B.n87 163.367
R508 B.n482 B.n87 163.367
R509 B.n482 B.n481 163.367
R510 B.n481 B.n480 163.367
R511 B.n480 B.n89 163.367
R512 B.n476 B.n89 163.367
R513 B.n476 B.n475 163.367
R514 B.n475 B.n474 163.367
R515 B.n474 B.n91 163.367
R516 B.n470 B.n91 163.367
R517 B.n470 B.n469 163.367
R518 B.n469 B.n468 163.367
R519 B.n468 B.n93 163.367
R520 B.n464 B.n93 163.367
R521 B.n464 B.n463 163.367
R522 B.n463 B.n462 163.367
R523 B.n462 B.n95 163.367
R524 B.n458 B.n95 163.367
R525 B.n458 B.n457 163.367
R526 B.n457 B.n456 163.367
R527 B.n456 B.n97 163.367
R528 B.n452 B.n97 163.367
R529 B.n452 B.n451 163.367
R530 B.n451 B.n450 163.367
R531 B.n450 B.n99 163.367
R532 B.n446 B.n99 163.367
R533 B.n446 B.n445 163.367
R534 B.n445 B.n444 163.367
R535 B.n444 B.n101 163.367
R536 B.n440 B.n101 163.367
R537 B.n440 B.n439 163.367
R538 B.n439 B.n438 163.367
R539 B.n438 B.n103 163.367
R540 B.n434 B.n103 163.367
R541 B.n434 B.n433 163.367
R542 B.n433 B.n432 163.367
R543 B.n432 B.n105 163.367
R544 B.n428 B.n105 163.367
R545 B.n428 B.n427 163.367
R546 B.n427 B.n426 163.367
R547 B.n426 B.n107 163.367
R548 B.n422 B.n107 163.367
R549 B.n422 B.n421 163.367
R550 B.n421 B.n420 163.367
R551 B.n420 B.n109 163.367
R552 B.n416 B.n109 163.367
R553 B.n416 B.n415 163.367
R554 B.n415 B.n414 163.367
R555 B.n684 B.n17 163.367
R556 B.n680 B.n17 163.367
R557 B.n680 B.n679 163.367
R558 B.n679 B.n678 163.367
R559 B.n678 B.n19 163.367
R560 B.n674 B.n19 163.367
R561 B.n674 B.n673 163.367
R562 B.n673 B.n672 163.367
R563 B.n672 B.n21 163.367
R564 B.n668 B.n21 163.367
R565 B.n668 B.n667 163.367
R566 B.n667 B.n666 163.367
R567 B.n666 B.n23 163.367
R568 B.n662 B.n23 163.367
R569 B.n662 B.n661 163.367
R570 B.n661 B.n660 163.367
R571 B.n660 B.n25 163.367
R572 B.n656 B.n25 163.367
R573 B.n656 B.n655 163.367
R574 B.n655 B.n654 163.367
R575 B.n654 B.n27 163.367
R576 B.n650 B.n27 163.367
R577 B.n650 B.n649 163.367
R578 B.n649 B.n648 163.367
R579 B.n648 B.n29 163.367
R580 B.n644 B.n29 163.367
R581 B.n644 B.n643 163.367
R582 B.n643 B.n642 163.367
R583 B.n642 B.n31 163.367
R584 B.n638 B.n31 163.367
R585 B.n638 B.n637 163.367
R586 B.n637 B.n636 163.367
R587 B.n636 B.n33 163.367
R588 B.n632 B.n33 163.367
R589 B.n632 B.n631 163.367
R590 B.n631 B.n630 163.367
R591 B.n630 B.n35 163.367
R592 B.n626 B.n35 163.367
R593 B.n626 B.n625 163.367
R594 B.n625 B.n624 163.367
R595 B.n624 B.n37 163.367
R596 B.n620 B.n37 163.367
R597 B.n620 B.n619 163.367
R598 B.n619 B.n618 163.367
R599 B.n618 B.n39 163.367
R600 B.n614 B.n39 163.367
R601 B.n614 B.n613 163.367
R602 B.n613 B.n612 163.367
R603 B.n612 B.n41 163.367
R604 B.n608 B.n41 163.367
R605 B.n608 B.n607 163.367
R606 B.n607 B.n606 163.367
R607 B.n606 B.n43 163.367
R608 B.n602 B.n43 163.367
R609 B.n602 B.n601 163.367
R610 B.n601 B.n47 163.367
R611 B.n597 B.n47 163.367
R612 B.n597 B.n596 163.367
R613 B.n596 B.n595 163.367
R614 B.n595 B.n49 163.367
R615 B.n591 B.n49 163.367
R616 B.n591 B.n590 163.367
R617 B.n590 B.n589 163.367
R618 B.n589 B.n51 163.367
R619 B.n584 B.n51 163.367
R620 B.n584 B.n583 163.367
R621 B.n583 B.n582 163.367
R622 B.n582 B.n55 163.367
R623 B.n578 B.n55 163.367
R624 B.n578 B.n577 163.367
R625 B.n577 B.n576 163.367
R626 B.n576 B.n57 163.367
R627 B.n572 B.n57 163.367
R628 B.n572 B.n571 163.367
R629 B.n571 B.n570 163.367
R630 B.n570 B.n59 163.367
R631 B.n566 B.n59 163.367
R632 B.n566 B.n565 163.367
R633 B.n565 B.n564 163.367
R634 B.n564 B.n61 163.367
R635 B.n560 B.n61 163.367
R636 B.n560 B.n559 163.367
R637 B.n559 B.n558 163.367
R638 B.n558 B.n63 163.367
R639 B.n554 B.n63 163.367
R640 B.n554 B.n553 163.367
R641 B.n553 B.n552 163.367
R642 B.n552 B.n65 163.367
R643 B.n548 B.n65 163.367
R644 B.n548 B.n547 163.367
R645 B.n547 B.n546 163.367
R646 B.n546 B.n67 163.367
R647 B.n542 B.n67 163.367
R648 B.n542 B.n541 163.367
R649 B.n541 B.n540 163.367
R650 B.n540 B.n69 163.367
R651 B.n536 B.n69 163.367
R652 B.n536 B.n535 163.367
R653 B.n535 B.n534 163.367
R654 B.n534 B.n71 163.367
R655 B.n530 B.n71 163.367
R656 B.n530 B.n529 163.367
R657 B.n529 B.n528 163.367
R658 B.n528 B.n73 163.367
R659 B.n524 B.n73 163.367
R660 B.n524 B.n523 163.367
R661 B.n523 B.n522 163.367
R662 B.n522 B.n75 163.367
R663 B.n518 B.n75 163.367
R664 B.n518 B.n517 163.367
R665 B.n517 B.n516 163.367
R666 B.n516 B.n77 163.367
R667 B.n512 B.n77 163.367
R668 B.n512 B.n511 163.367
R669 B.n511 B.n510 163.367
R670 B.n510 B.n79 163.367
R671 B.n506 B.n79 163.367
R672 B.n506 B.n505 163.367
R673 B.n505 B.n504 163.367
R674 B.n686 B.n685 163.367
R675 B.n686 B.n15 163.367
R676 B.n690 B.n15 163.367
R677 B.n691 B.n690 163.367
R678 B.n692 B.n691 163.367
R679 B.n692 B.n13 163.367
R680 B.n696 B.n13 163.367
R681 B.n697 B.n696 163.367
R682 B.n698 B.n697 163.367
R683 B.n698 B.n11 163.367
R684 B.n702 B.n11 163.367
R685 B.n703 B.n702 163.367
R686 B.n704 B.n703 163.367
R687 B.n704 B.n9 163.367
R688 B.n708 B.n9 163.367
R689 B.n709 B.n708 163.367
R690 B.n710 B.n709 163.367
R691 B.n710 B.n7 163.367
R692 B.n714 B.n7 163.367
R693 B.n715 B.n714 163.367
R694 B.n716 B.n715 163.367
R695 B.n716 B.n5 163.367
R696 B.n720 B.n5 163.367
R697 B.n721 B.n720 163.367
R698 B.n722 B.n721 163.367
R699 B.n722 B.n3 163.367
R700 B.n726 B.n3 163.367
R701 B.n727 B.n726 163.367
R702 B.n188 B.n2 163.367
R703 B.n189 B.n188 163.367
R704 B.n190 B.n189 163.367
R705 B.n190 B.n185 163.367
R706 B.n194 B.n185 163.367
R707 B.n195 B.n194 163.367
R708 B.n196 B.n195 163.367
R709 B.n196 B.n183 163.367
R710 B.n200 B.n183 163.367
R711 B.n201 B.n200 163.367
R712 B.n202 B.n201 163.367
R713 B.n202 B.n181 163.367
R714 B.n206 B.n181 163.367
R715 B.n207 B.n206 163.367
R716 B.n208 B.n207 163.367
R717 B.n208 B.n179 163.367
R718 B.n212 B.n179 163.367
R719 B.n213 B.n212 163.367
R720 B.n214 B.n213 163.367
R721 B.n214 B.n177 163.367
R722 B.n218 B.n177 163.367
R723 B.n219 B.n218 163.367
R724 B.n220 B.n219 163.367
R725 B.n220 B.n175 163.367
R726 B.n224 B.n175 163.367
R727 B.n225 B.n224 163.367
R728 B.n226 B.n225 163.367
R729 B.n226 B.n173 163.367
R730 B.n145 B.n144 70.7884
R731 B.n327 B.n326 70.7884
R732 B.n53 B.n52 70.7884
R733 B.n45 B.n44 70.7884
R734 B.n312 B.n145 59.5399
R735 B.n328 B.n327 59.5399
R736 B.n586 B.n53 59.5399
R737 B.n46 B.n45 59.5399
R738 B.n683 B.n16 35.7468
R739 B.n503 B.n502 35.7468
R740 B.n229 B.n228 35.7468
R741 B.n413 B.n412 35.7468
R742 B B.n729 18.0485
R743 B.n687 B.n16 10.6151
R744 B.n688 B.n687 10.6151
R745 B.n689 B.n688 10.6151
R746 B.n689 B.n14 10.6151
R747 B.n693 B.n14 10.6151
R748 B.n694 B.n693 10.6151
R749 B.n695 B.n694 10.6151
R750 B.n695 B.n12 10.6151
R751 B.n699 B.n12 10.6151
R752 B.n700 B.n699 10.6151
R753 B.n701 B.n700 10.6151
R754 B.n701 B.n10 10.6151
R755 B.n705 B.n10 10.6151
R756 B.n706 B.n705 10.6151
R757 B.n707 B.n706 10.6151
R758 B.n707 B.n8 10.6151
R759 B.n711 B.n8 10.6151
R760 B.n712 B.n711 10.6151
R761 B.n713 B.n712 10.6151
R762 B.n713 B.n6 10.6151
R763 B.n717 B.n6 10.6151
R764 B.n718 B.n717 10.6151
R765 B.n719 B.n718 10.6151
R766 B.n719 B.n4 10.6151
R767 B.n723 B.n4 10.6151
R768 B.n724 B.n723 10.6151
R769 B.n725 B.n724 10.6151
R770 B.n725 B.n0 10.6151
R771 B.n683 B.n682 10.6151
R772 B.n682 B.n681 10.6151
R773 B.n681 B.n18 10.6151
R774 B.n677 B.n18 10.6151
R775 B.n677 B.n676 10.6151
R776 B.n676 B.n675 10.6151
R777 B.n675 B.n20 10.6151
R778 B.n671 B.n20 10.6151
R779 B.n671 B.n670 10.6151
R780 B.n670 B.n669 10.6151
R781 B.n669 B.n22 10.6151
R782 B.n665 B.n22 10.6151
R783 B.n665 B.n664 10.6151
R784 B.n664 B.n663 10.6151
R785 B.n663 B.n24 10.6151
R786 B.n659 B.n24 10.6151
R787 B.n659 B.n658 10.6151
R788 B.n658 B.n657 10.6151
R789 B.n657 B.n26 10.6151
R790 B.n653 B.n26 10.6151
R791 B.n653 B.n652 10.6151
R792 B.n652 B.n651 10.6151
R793 B.n651 B.n28 10.6151
R794 B.n647 B.n28 10.6151
R795 B.n647 B.n646 10.6151
R796 B.n646 B.n645 10.6151
R797 B.n645 B.n30 10.6151
R798 B.n641 B.n30 10.6151
R799 B.n641 B.n640 10.6151
R800 B.n640 B.n639 10.6151
R801 B.n639 B.n32 10.6151
R802 B.n635 B.n32 10.6151
R803 B.n635 B.n634 10.6151
R804 B.n634 B.n633 10.6151
R805 B.n633 B.n34 10.6151
R806 B.n629 B.n34 10.6151
R807 B.n629 B.n628 10.6151
R808 B.n628 B.n627 10.6151
R809 B.n627 B.n36 10.6151
R810 B.n623 B.n36 10.6151
R811 B.n623 B.n622 10.6151
R812 B.n622 B.n621 10.6151
R813 B.n621 B.n38 10.6151
R814 B.n617 B.n38 10.6151
R815 B.n617 B.n616 10.6151
R816 B.n616 B.n615 10.6151
R817 B.n615 B.n40 10.6151
R818 B.n611 B.n40 10.6151
R819 B.n611 B.n610 10.6151
R820 B.n610 B.n609 10.6151
R821 B.n609 B.n42 10.6151
R822 B.n605 B.n42 10.6151
R823 B.n605 B.n604 10.6151
R824 B.n604 B.n603 10.6151
R825 B.n600 B.n599 10.6151
R826 B.n599 B.n598 10.6151
R827 B.n598 B.n48 10.6151
R828 B.n594 B.n48 10.6151
R829 B.n594 B.n593 10.6151
R830 B.n593 B.n592 10.6151
R831 B.n592 B.n50 10.6151
R832 B.n588 B.n50 10.6151
R833 B.n588 B.n587 10.6151
R834 B.n585 B.n54 10.6151
R835 B.n581 B.n54 10.6151
R836 B.n581 B.n580 10.6151
R837 B.n580 B.n579 10.6151
R838 B.n579 B.n56 10.6151
R839 B.n575 B.n56 10.6151
R840 B.n575 B.n574 10.6151
R841 B.n574 B.n573 10.6151
R842 B.n573 B.n58 10.6151
R843 B.n569 B.n58 10.6151
R844 B.n569 B.n568 10.6151
R845 B.n568 B.n567 10.6151
R846 B.n567 B.n60 10.6151
R847 B.n563 B.n60 10.6151
R848 B.n563 B.n562 10.6151
R849 B.n562 B.n561 10.6151
R850 B.n561 B.n62 10.6151
R851 B.n557 B.n62 10.6151
R852 B.n557 B.n556 10.6151
R853 B.n556 B.n555 10.6151
R854 B.n555 B.n64 10.6151
R855 B.n551 B.n64 10.6151
R856 B.n551 B.n550 10.6151
R857 B.n550 B.n549 10.6151
R858 B.n549 B.n66 10.6151
R859 B.n545 B.n66 10.6151
R860 B.n545 B.n544 10.6151
R861 B.n544 B.n543 10.6151
R862 B.n543 B.n68 10.6151
R863 B.n539 B.n68 10.6151
R864 B.n539 B.n538 10.6151
R865 B.n538 B.n537 10.6151
R866 B.n537 B.n70 10.6151
R867 B.n533 B.n70 10.6151
R868 B.n533 B.n532 10.6151
R869 B.n532 B.n531 10.6151
R870 B.n531 B.n72 10.6151
R871 B.n527 B.n72 10.6151
R872 B.n527 B.n526 10.6151
R873 B.n526 B.n525 10.6151
R874 B.n525 B.n74 10.6151
R875 B.n521 B.n74 10.6151
R876 B.n521 B.n520 10.6151
R877 B.n520 B.n519 10.6151
R878 B.n519 B.n76 10.6151
R879 B.n515 B.n76 10.6151
R880 B.n515 B.n514 10.6151
R881 B.n514 B.n513 10.6151
R882 B.n513 B.n78 10.6151
R883 B.n509 B.n78 10.6151
R884 B.n509 B.n508 10.6151
R885 B.n508 B.n507 10.6151
R886 B.n507 B.n80 10.6151
R887 B.n503 B.n80 10.6151
R888 B.n502 B.n501 10.6151
R889 B.n501 B.n82 10.6151
R890 B.n497 B.n82 10.6151
R891 B.n497 B.n496 10.6151
R892 B.n496 B.n495 10.6151
R893 B.n495 B.n84 10.6151
R894 B.n491 B.n84 10.6151
R895 B.n491 B.n490 10.6151
R896 B.n490 B.n489 10.6151
R897 B.n489 B.n86 10.6151
R898 B.n485 B.n86 10.6151
R899 B.n485 B.n484 10.6151
R900 B.n484 B.n483 10.6151
R901 B.n483 B.n88 10.6151
R902 B.n479 B.n88 10.6151
R903 B.n479 B.n478 10.6151
R904 B.n478 B.n477 10.6151
R905 B.n477 B.n90 10.6151
R906 B.n473 B.n90 10.6151
R907 B.n473 B.n472 10.6151
R908 B.n472 B.n471 10.6151
R909 B.n471 B.n92 10.6151
R910 B.n467 B.n92 10.6151
R911 B.n467 B.n466 10.6151
R912 B.n466 B.n465 10.6151
R913 B.n465 B.n94 10.6151
R914 B.n461 B.n94 10.6151
R915 B.n461 B.n460 10.6151
R916 B.n460 B.n459 10.6151
R917 B.n459 B.n96 10.6151
R918 B.n455 B.n96 10.6151
R919 B.n455 B.n454 10.6151
R920 B.n454 B.n453 10.6151
R921 B.n453 B.n98 10.6151
R922 B.n449 B.n98 10.6151
R923 B.n449 B.n448 10.6151
R924 B.n448 B.n447 10.6151
R925 B.n447 B.n100 10.6151
R926 B.n443 B.n100 10.6151
R927 B.n443 B.n442 10.6151
R928 B.n442 B.n441 10.6151
R929 B.n441 B.n102 10.6151
R930 B.n437 B.n102 10.6151
R931 B.n437 B.n436 10.6151
R932 B.n436 B.n435 10.6151
R933 B.n435 B.n104 10.6151
R934 B.n431 B.n104 10.6151
R935 B.n431 B.n430 10.6151
R936 B.n430 B.n429 10.6151
R937 B.n429 B.n106 10.6151
R938 B.n425 B.n106 10.6151
R939 B.n425 B.n424 10.6151
R940 B.n424 B.n423 10.6151
R941 B.n423 B.n108 10.6151
R942 B.n419 B.n108 10.6151
R943 B.n419 B.n418 10.6151
R944 B.n418 B.n417 10.6151
R945 B.n417 B.n110 10.6151
R946 B.n413 B.n110 10.6151
R947 B.n187 B.n1 10.6151
R948 B.n187 B.n186 10.6151
R949 B.n191 B.n186 10.6151
R950 B.n192 B.n191 10.6151
R951 B.n193 B.n192 10.6151
R952 B.n193 B.n184 10.6151
R953 B.n197 B.n184 10.6151
R954 B.n198 B.n197 10.6151
R955 B.n199 B.n198 10.6151
R956 B.n199 B.n182 10.6151
R957 B.n203 B.n182 10.6151
R958 B.n204 B.n203 10.6151
R959 B.n205 B.n204 10.6151
R960 B.n205 B.n180 10.6151
R961 B.n209 B.n180 10.6151
R962 B.n210 B.n209 10.6151
R963 B.n211 B.n210 10.6151
R964 B.n211 B.n178 10.6151
R965 B.n215 B.n178 10.6151
R966 B.n216 B.n215 10.6151
R967 B.n217 B.n216 10.6151
R968 B.n217 B.n176 10.6151
R969 B.n221 B.n176 10.6151
R970 B.n222 B.n221 10.6151
R971 B.n223 B.n222 10.6151
R972 B.n223 B.n174 10.6151
R973 B.n227 B.n174 10.6151
R974 B.n228 B.n227 10.6151
R975 B.n229 B.n172 10.6151
R976 B.n233 B.n172 10.6151
R977 B.n234 B.n233 10.6151
R978 B.n235 B.n234 10.6151
R979 B.n235 B.n170 10.6151
R980 B.n239 B.n170 10.6151
R981 B.n240 B.n239 10.6151
R982 B.n241 B.n240 10.6151
R983 B.n241 B.n168 10.6151
R984 B.n245 B.n168 10.6151
R985 B.n246 B.n245 10.6151
R986 B.n247 B.n246 10.6151
R987 B.n247 B.n166 10.6151
R988 B.n251 B.n166 10.6151
R989 B.n252 B.n251 10.6151
R990 B.n253 B.n252 10.6151
R991 B.n253 B.n164 10.6151
R992 B.n257 B.n164 10.6151
R993 B.n258 B.n257 10.6151
R994 B.n259 B.n258 10.6151
R995 B.n259 B.n162 10.6151
R996 B.n263 B.n162 10.6151
R997 B.n264 B.n263 10.6151
R998 B.n265 B.n264 10.6151
R999 B.n265 B.n160 10.6151
R1000 B.n269 B.n160 10.6151
R1001 B.n270 B.n269 10.6151
R1002 B.n271 B.n270 10.6151
R1003 B.n271 B.n158 10.6151
R1004 B.n275 B.n158 10.6151
R1005 B.n276 B.n275 10.6151
R1006 B.n277 B.n276 10.6151
R1007 B.n277 B.n156 10.6151
R1008 B.n281 B.n156 10.6151
R1009 B.n282 B.n281 10.6151
R1010 B.n283 B.n282 10.6151
R1011 B.n283 B.n154 10.6151
R1012 B.n287 B.n154 10.6151
R1013 B.n288 B.n287 10.6151
R1014 B.n289 B.n288 10.6151
R1015 B.n289 B.n152 10.6151
R1016 B.n293 B.n152 10.6151
R1017 B.n294 B.n293 10.6151
R1018 B.n295 B.n294 10.6151
R1019 B.n295 B.n150 10.6151
R1020 B.n299 B.n150 10.6151
R1021 B.n300 B.n299 10.6151
R1022 B.n301 B.n300 10.6151
R1023 B.n301 B.n148 10.6151
R1024 B.n305 B.n148 10.6151
R1025 B.n306 B.n305 10.6151
R1026 B.n307 B.n306 10.6151
R1027 B.n307 B.n146 10.6151
R1028 B.n311 B.n146 10.6151
R1029 B.n314 B.n313 10.6151
R1030 B.n314 B.n142 10.6151
R1031 B.n318 B.n142 10.6151
R1032 B.n319 B.n318 10.6151
R1033 B.n320 B.n319 10.6151
R1034 B.n320 B.n140 10.6151
R1035 B.n324 B.n140 10.6151
R1036 B.n325 B.n324 10.6151
R1037 B.n329 B.n325 10.6151
R1038 B.n333 B.n138 10.6151
R1039 B.n334 B.n333 10.6151
R1040 B.n335 B.n334 10.6151
R1041 B.n335 B.n136 10.6151
R1042 B.n339 B.n136 10.6151
R1043 B.n340 B.n339 10.6151
R1044 B.n341 B.n340 10.6151
R1045 B.n341 B.n134 10.6151
R1046 B.n345 B.n134 10.6151
R1047 B.n346 B.n345 10.6151
R1048 B.n347 B.n346 10.6151
R1049 B.n347 B.n132 10.6151
R1050 B.n351 B.n132 10.6151
R1051 B.n352 B.n351 10.6151
R1052 B.n353 B.n352 10.6151
R1053 B.n353 B.n130 10.6151
R1054 B.n357 B.n130 10.6151
R1055 B.n358 B.n357 10.6151
R1056 B.n359 B.n358 10.6151
R1057 B.n359 B.n128 10.6151
R1058 B.n363 B.n128 10.6151
R1059 B.n364 B.n363 10.6151
R1060 B.n365 B.n364 10.6151
R1061 B.n365 B.n126 10.6151
R1062 B.n369 B.n126 10.6151
R1063 B.n370 B.n369 10.6151
R1064 B.n371 B.n370 10.6151
R1065 B.n371 B.n124 10.6151
R1066 B.n375 B.n124 10.6151
R1067 B.n376 B.n375 10.6151
R1068 B.n377 B.n376 10.6151
R1069 B.n377 B.n122 10.6151
R1070 B.n381 B.n122 10.6151
R1071 B.n382 B.n381 10.6151
R1072 B.n383 B.n382 10.6151
R1073 B.n383 B.n120 10.6151
R1074 B.n387 B.n120 10.6151
R1075 B.n388 B.n387 10.6151
R1076 B.n389 B.n388 10.6151
R1077 B.n389 B.n118 10.6151
R1078 B.n393 B.n118 10.6151
R1079 B.n394 B.n393 10.6151
R1080 B.n395 B.n394 10.6151
R1081 B.n395 B.n116 10.6151
R1082 B.n399 B.n116 10.6151
R1083 B.n400 B.n399 10.6151
R1084 B.n401 B.n400 10.6151
R1085 B.n401 B.n114 10.6151
R1086 B.n405 B.n114 10.6151
R1087 B.n406 B.n405 10.6151
R1088 B.n407 B.n406 10.6151
R1089 B.n407 B.n112 10.6151
R1090 B.n411 B.n112 10.6151
R1091 B.n412 B.n411 10.6151
R1092 B.n603 B.n46 9.36635
R1093 B.n586 B.n585 9.36635
R1094 B.n312 B.n311 9.36635
R1095 B.n328 B.n138 9.36635
R1096 B.n729 B.n0 8.11757
R1097 B.n729 B.n1 8.11757
R1098 B.n600 B.n46 1.24928
R1099 B.n587 B.n586 1.24928
R1100 B.n313 B.n312 1.24928
R1101 B.n329 B.n328 1.24928
R1102 VN VN.t0 210.106
R1103 VN VN.t1 160.597
R1104 VTAIL.n370 VTAIL.n282 756.745
R1105 VTAIL.n88 VTAIL.n0 756.745
R1106 VTAIL.n276 VTAIL.n188 756.745
R1107 VTAIL.n182 VTAIL.n94 756.745
R1108 VTAIL.n313 VTAIL.n312 585
R1109 VTAIL.n310 VTAIL.n309 585
R1110 VTAIL.n319 VTAIL.n318 585
R1111 VTAIL.n321 VTAIL.n320 585
R1112 VTAIL.n306 VTAIL.n305 585
R1113 VTAIL.n327 VTAIL.n326 585
R1114 VTAIL.n329 VTAIL.n328 585
R1115 VTAIL.n302 VTAIL.n301 585
R1116 VTAIL.n335 VTAIL.n334 585
R1117 VTAIL.n337 VTAIL.n336 585
R1118 VTAIL.n298 VTAIL.n297 585
R1119 VTAIL.n343 VTAIL.n342 585
R1120 VTAIL.n345 VTAIL.n344 585
R1121 VTAIL.n294 VTAIL.n293 585
R1122 VTAIL.n351 VTAIL.n350 585
R1123 VTAIL.n354 VTAIL.n353 585
R1124 VTAIL.n352 VTAIL.n290 585
R1125 VTAIL.n359 VTAIL.n289 585
R1126 VTAIL.n361 VTAIL.n360 585
R1127 VTAIL.n363 VTAIL.n362 585
R1128 VTAIL.n286 VTAIL.n285 585
R1129 VTAIL.n369 VTAIL.n368 585
R1130 VTAIL.n371 VTAIL.n370 585
R1131 VTAIL.n31 VTAIL.n30 585
R1132 VTAIL.n28 VTAIL.n27 585
R1133 VTAIL.n37 VTAIL.n36 585
R1134 VTAIL.n39 VTAIL.n38 585
R1135 VTAIL.n24 VTAIL.n23 585
R1136 VTAIL.n45 VTAIL.n44 585
R1137 VTAIL.n47 VTAIL.n46 585
R1138 VTAIL.n20 VTAIL.n19 585
R1139 VTAIL.n53 VTAIL.n52 585
R1140 VTAIL.n55 VTAIL.n54 585
R1141 VTAIL.n16 VTAIL.n15 585
R1142 VTAIL.n61 VTAIL.n60 585
R1143 VTAIL.n63 VTAIL.n62 585
R1144 VTAIL.n12 VTAIL.n11 585
R1145 VTAIL.n69 VTAIL.n68 585
R1146 VTAIL.n72 VTAIL.n71 585
R1147 VTAIL.n70 VTAIL.n8 585
R1148 VTAIL.n77 VTAIL.n7 585
R1149 VTAIL.n79 VTAIL.n78 585
R1150 VTAIL.n81 VTAIL.n80 585
R1151 VTAIL.n4 VTAIL.n3 585
R1152 VTAIL.n87 VTAIL.n86 585
R1153 VTAIL.n89 VTAIL.n88 585
R1154 VTAIL.n277 VTAIL.n276 585
R1155 VTAIL.n275 VTAIL.n274 585
R1156 VTAIL.n192 VTAIL.n191 585
R1157 VTAIL.n269 VTAIL.n268 585
R1158 VTAIL.n267 VTAIL.n266 585
R1159 VTAIL.n265 VTAIL.n195 585
R1160 VTAIL.n199 VTAIL.n196 585
R1161 VTAIL.n260 VTAIL.n259 585
R1162 VTAIL.n258 VTAIL.n257 585
R1163 VTAIL.n201 VTAIL.n200 585
R1164 VTAIL.n252 VTAIL.n251 585
R1165 VTAIL.n250 VTAIL.n249 585
R1166 VTAIL.n205 VTAIL.n204 585
R1167 VTAIL.n244 VTAIL.n243 585
R1168 VTAIL.n242 VTAIL.n241 585
R1169 VTAIL.n209 VTAIL.n208 585
R1170 VTAIL.n236 VTAIL.n235 585
R1171 VTAIL.n234 VTAIL.n233 585
R1172 VTAIL.n213 VTAIL.n212 585
R1173 VTAIL.n228 VTAIL.n227 585
R1174 VTAIL.n226 VTAIL.n225 585
R1175 VTAIL.n217 VTAIL.n216 585
R1176 VTAIL.n220 VTAIL.n219 585
R1177 VTAIL.n183 VTAIL.n182 585
R1178 VTAIL.n181 VTAIL.n180 585
R1179 VTAIL.n98 VTAIL.n97 585
R1180 VTAIL.n175 VTAIL.n174 585
R1181 VTAIL.n173 VTAIL.n172 585
R1182 VTAIL.n171 VTAIL.n101 585
R1183 VTAIL.n105 VTAIL.n102 585
R1184 VTAIL.n166 VTAIL.n165 585
R1185 VTAIL.n164 VTAIL.n163 585
R1186 VTAIL.n107 VTAIL.n106 585
R1187 VTAIL.n158 VTAIL.n157 585
R1188 VTAIL.n156 VTAIL.n155 585
R1189 VTAIL.n111 VTAIL.n110 585
R1190 VTAIL.n150 VTAIL.n149 585
R1191 VTAIL.n148 VTAIL.n147 585
R1192 VTAIL.n115 VTAIL.n114 585
R1193 VTAIL.n142 VTAIL.n141 585
R1194 VTAIL.n140 VTAIL.n139 585
R1195 VTAIL.n119 VTAIL.n118 585
R1196 VTAIL.n134 VTAIL.n133 585
R1197 VTAIL.n132 VTAIL.n131 585
R1198 VTAIL.n123 VTAIL.n122 585
R1199 VTAIL.n126 VTAIL.n125 585
R1200 VTAIL.t2 VTAIL.n218 327.466
R1201 VTAIL.t0 VTAIL.n124 327.466
R1202 VTAIL.t1 VTAIL.n311 327.466
R1203 VTAIL.t3 VTAIL.n29 327.466
R1204 VTAIL.n312 VTAIL.n309 171.744
R1205 VTAIL.n319 VTAIL.n309 171.744
R1206 VTAIL.n320 VTAIL.n319 171.744
R1207 VTAIL.n320 VTAIL.n305 171.744
R1208 VTAIL.n327 VTAIL.n305 171.744
R1209 VTAIL.n328 VTAIL.n327 171.744
R1210 VTAIL.n328 VTAIL.n301 171.744
R1211 VTAIL.n335 VTAIL.n301 171.744
R1212 VTAIL.n336 VTAIL.n335 171.744
R1213 VTAIL.n336 VTAIL.n297 171.744
R1214 VTAIL.n343 VTAIL.n297 171.744
R1215 VTAIL.n344 VTAIL.n343 171.744
R1216 VTAIL.n344 VTAIL.n293 171.744
R1217 VTAIL.n351 VTAIL.n293 171.744
R1218 VTAIL.n353 VTAIL.n351 171.744
R1219 VTAIL.n353 VTAIL.n352 171.744
R1220 VTAIL.n352 VTAIL.n289 171.744
R1221 VTAIL.n361 VTAIL.n289 171.744
R1222 VTAIL.n362 VTAIL.n361 171.744
R1223 VTAIL.n362 VTAIL.n285 171.744
R1224 VTAIL.n369 VTAIL.n285 171.744
R1225 VTAIL.n370 VTAIL.n369 171.744
R1226 VTAIL.n30 VTAIL.n27 171.744
R1227 VTAIL.n37 VTAIL.n27 171.744
R1228 VTAIL.n38 VTAIL.n37 171.744
R1229 VTAIL.n38 VTAIL.n23 171.744
R1230 VTAIL.n45 VTAIL.n23 171.744
R1231 VTAIL.n46 VTAIL.n45 171.744
R1232 VTAIL.n46 VTAIL.n19 171.744
R1233 VTAIL.n53 VTAIL.n19 171.744
R1234 VTAIL.n54 VTAIL.n53 171.744
R1235 VTAIL.n54 VTAIL.n15 171.744
R1236 VTAIL.n61 VTAIL.n15 171.744
R1237 VTAIL.n62 VTAIL.n61 171.744
R1238 VTAIL.n62 VTAIL.n11 171.744
R1239 VTAIL.n69 VTAIL.n11 171.744
R1240 VTAIL.n71 VTAIL.n69 171.744
R1241 VTAIL.n71 VTAIL.n70 171.744
R1242 VTAIL.n70 VTAIL.n7 171.744
R1243 VTAIL.n79 VTAIL.n7 171.744
R1244 VTAIL.n80 VTAIL.n79 171.744
R1245 VTAIL.n80 VTAIL.n3 171.744
R1246 VTAIL.n87 VTAIL.n3 171.744
R1247 VTAIL.n88 VTAIL.n87 171.744
R1248 VTAIL.n276 VTAIL.n275 171.744
R1249 VTAIL.n275 VTAIL.n191 171.744
R1250 VTAIL.n268 VTAIL.n191 171.744
R1251 VTAIL.n268 VTAIL.n267 171.744
R1252 VTAIL.n267 VTAIL.n195 171.744
R1253 VTAIL.n199 VTAIL.n195 171.744
R1254 VTAIL.n259 VTAIL.n199 171.744
R1255 VTAIL.n259 VTAIL.n258 171.744
R1256 VTAIL.n258 VTAIL.n200 171.744
R1257 VTAIL.n251 VTAIL.n200 171.744
R1258 VTAIL.n251 VTAIL.n250 171.744
R1259 VTAIL.n250 VTAIL.n204 171.744
R1260 VTAIL.n243 VTAIL.n204 171.744
R1261 VTAIL.n243 VTAIL.n242 171.744
R1262 VTAIL.n242 VTAIL.n208 171.744
R1263 VTAIL.n235 VTAIL.n208 171.744
R1264 VTAIL.n235 VTAIL.n234 171.744
R1265 VTAIL.n234 VTAIL.n212 171.744
R1266 VTAIL.n227 VTAIL.n212 171.744
R1267 VTAIL.n227 VTAIL.n226 171.744
R1268 VTAIL.n226 VTAIL.n216 171.744
R1269 VTAIL.n219 VTAIL.n216 171.744
R1270 VTAIL.n182 VTAIL.n181 171.744
R1271 VTAIL.n181 VTAIL.n97 171.744
R1272 VTAIL.n174 VTAIL.n97 171.744
R1273 VTAIL.n174 VTAIL.n173 171.744
R1274 VTAIL.n173 VTAIL.n101 171.744
R1275 VTAIL.n105 VTAIL.n101 171.744
R1276 VTAIL.n165 VTAIL.n105 171.744
R1277 VTAIL.n165 VTAIL.n164 171.744
R1278 VTAIL.n164 VTAIL.n106 171.744
R1279 VTAIL.n157 VTAIL.n106 171.744
R1280 VTAIL.n157 VTAIL.n156 171.744
R1281 VTAIL.n156 VTAIL.n110 171.744
R1282 VTAIL.n149 VTAIL.n110 171.744
R1283 VTAIL.n149 VTAIL.n148 171.744
R1284 VTAIL.n148 VTAIL.n114 171.744
R1285 VTAIL.n141 VTAIL.n114 171.744
R1286 VTAIL.n141 VTAIL.n140 171.744
R1287 VTAIL.n140 VTAIL.n118 171.744
R1288 VTAIL.n133 VTAIL.n118 171.744
R1289 VTAIL.n133 VTAIL.n132 171.744
R1290 VTAIL.n132 VTAIL.n122 171.744
R1291 VTAIL.n125 VTAIL.n122 171.744
R1292 VTAIL.n312 VTAIL.t1 85.8723
R1293 VTAIL.n30 VTAIL.t3 85.8723
R1294 VTAIL.n219 VTAIL.t2 85.8723
R1295 VTAIL.n125 VTAIL.t0 85.8723
R1296 VTAIL.n187 VTAIL.n93 33.0565
R1297 VTAIL.n375 VTAIL.n374 30.246
R1298 VTAIL.n93 VTAIL.n92 30.246
R1299 VTAIL.n281 VTAIL.n280 30.246
R1300 VTAIL.n187 VTAIL.n186 30.246
R1301 VTAIL.n375 VTAIL.n281 29.91
R1302 VTAIL.n313 VTAIL.n311 16.3895
R1303 VTAIL.n31 VTAIL.n29 16.3895
R1304 VTAIL.n220 VTAIL.n218 16.3895
R1305 VTAIL.n126 VTAIL.n124 16.3895
R1306 VTAIL.n360 VTAIL.n359 13.1884
R1307 VTAIL.n78 VTAIL.n77 13.1884
R1308 VTAIL.n266 VTAIL.n265 13.1884
R1309 VTAIL.n172 VTAIL.n171 13.1884
R1310 VTAIL.n314 VTAIL.n310 12.8005
R1311 VTAIL.n358 VTAIL.n290 12.8005
R1312 VTAIL.n363 VTAIL.n288 12.8005
R1313 VTAIL.n32 VTAIL.n28 12.8005
R1314 VTAIL.n76 VTAIL.n8 12.8005
R1315 VTAIL.n81 VTAIL.n6 12.8005
R1316 VTAIL.n269 VTAIL.n194 12.8005
R1317 VTAIL.n264 VTAIL.n196 12.8005
R1318 VTAIL.n221 VTAIL.n217 12.8005
R1319 VTAIL.n175 VTAIL.n100 12.8005
R1320 VTAIL.n170 VTAIL.n102 12.8005
R1321 VTAIL.n127 VTAIL.n123 12.8005
R1322 VTAIL.n318 VTAIL.n317 12.0247
R1323 VTAIL.n355 VTAIL.n354 12.0247
R1324 VTAIL.n364 VTAIL.n286 12.0247
R1325 VTAIL.n36 VTAIL.n35 12.0247
R1326 VTAIL.n73 VTAIL.n72 12.0247
R1327 VTAIL.n82 VTAIL.n4 12.0247
R1328 VTAIL.n270 VTAIL.n192 12.0247
R1329 VTAIL.n261 VTAIL.n260 12.0247
R1330 VTAIL.n225 VTAIL.n224 12.0247
R1331 VTAIL.n176 VTAIL.n98 12.0247
R1332 VTAIL.n167 VTAIL.n166 12.0247
R1333 VTAIL.n131 VTAIL.n130 12.0247
R1334 VTAIL.n321 VTAIL.n308 11.249
R1335 VTAIL.n350 VTAIL.n292 11.249
R1336 VTAIL.n368 VTAIL.n367 11.249
R1337 VTAIL.n39 VTAIL.n26 11.249
R1338 VTAIL.n68 VTAIL.n10 11.249
R1339 VTAIL.n86 VTAIL.n85 11.249
R1340 VTAIL.n274 VTAIL.n273 11.249
R1341 VTAIL.n257 VTAIL.n198 11.249
R1342 VTAIL.n228 VTAIL.n215 11.249
R1343 VTAIL.n180 VTAIL.n179 11.249
R1344 VTAIL.n163 VTAIL.n104 11.249
R1345 VTAIL.n134 VTAIL.n121 11.249
R1346 VTAIL.n322 VTAIL.n306 10.4732
R1347 VTAIL.n349 VTAIL.n294 10.4732
R1348 VTAIL.n371 VTAIL.n284 10.4732
R1349 VTAIL.n40 VTAIL.n24 10.4732
R1350 VTAIL.n67 VTAIL.n12 10.4732
R1351 VTAIL.n89 VTAIL.n2 10.4732
R1352 VTAIL.n277 VTAIL.n190 10.4732
R1353 VTAIL.n256 VTAIL.n201 10.4732
R1354 VTAIL.n229 VTAIL.n213 10.4732
R1355 VTAIL.n183 VTAIL.n96 10.4732
R1356 VTAIL.n162 VTAIL.n107 10.4732
R1357 VTAIL.n135 VTAIL.n119 10.4732
R1358 VTAIL.n326 VTAIL.n325 9.69747
R1359 VTAIL.n346 VTAIL.n345 9.69747
R1360 VTAIL.n372 VTAIL.n282 9.69747
R1361 VTAIL.n44 VTAIL.n43 9.69747
R1362 VTAIL.n64 VTAIL.n63 9.69747
R1363 VTAIL.n90 VTAIL.n0 9.69747
R1364 VTAIL.n278 VTAIL.n188 9.69747
R1365 VTAIL.n253 VTAIL.n252 9.69747
R1366 VTAIL.n233 VTAIL.n232 9.69747
R1367 VTAIL.n184 VTAIL.n94 9.69747
R1368 VTAIL.n159 VTAIL.n158 9.69747
R1369 VTAIL.n139 VTAIL.n138 9.69747
R1370 VTAIL.n374 VTAIL.n373 9.45567
R1371 VTAIL.n92 VTAIL.n91 9.45567
R1372 VTAIL.n280 VTAIL.n279 9.45567
R1373 VTAIL.n186 VTAIL.n185 9.45567
R1374 VTAIL.n373 VTAIL.n372 9.3005
R1375 VTAIL.n284 VTAIL.n283 9.3005
R1376 VTAIL.n367 VTAIL.n366 9.3005
R1377 VTAIL.n365 VTAIL.n364 9.3005
R1378 VTAIL.n288 VTAIL.n287 9.3005
R1379 VTAIL.n333 VTAIL.n332 9.3005
R1380 VTAIL.n331 VTAIL.n330 9.3005
R1381 VTAIL.n304 VTAIL.n303 9.3005
R1382 VTAIL.n325 VTAIL.n324 9.3005
R1383 VTAIL.n323 VTAIL.n322 9.3005
R1384 VTAIL.n308 VTAIL.n307 9.3005
R1385 VTAIL.n317 VTAIL.n316 9.3005
R1386 VTAIL.n315 VTAIL.n314 9.3005
R1387 VTAIL.n300 VTAIL.n299 9.3005
R1388 VTAIL.n339 VTAIL.n338 9.3005
R1389 VTAIL.n341 VTAIL.n340 9.3005
R1390 VTAIL.n296 VTAIL.n295 9.3005
R1391 VTAIL.n347 VTAIL.n346 9.3005
R1392 VTAIL.n349 VTAIL.n348 9.3005
R1393 VTAIL.n292 VTAIL.n291 9.3005
R1394 VTAIL.n356 VTAIL.n355 9.3005
R1395 VTAIL.n358 VTAIL.n357 9.3005
R1396 VTAIL.n91 VTAIL.n90 9.3005
R1397 VTAIL.n2 VTAIL.n1 9.3005
R1398 VTAIL.n85 VTAIL.n84 9.3005
R1399 VTAIL.n83 VTAIL.n82 9.3005
R1400 VTAIL.n6 VTAIL.n5 9.3005
R1401 VTAIL.n51 VTAIL.n50 9.3005
R1402 VTAIL.n49 VTAIL.n48 9.3005
R1403 VTAIL.n22 VTAIL.n21 9.3005
R1404 VTAIL.n43 VTAIL.n42 9.3005
R1405 VTAIL.n41 VTAIL.n40 9.3005
R1406 VTAIL.n26 VTAIL.n25 9.3005
R1407 VTAIL.n35 VTAIL.n34 9.3005
R1408 VTAIL.n33 VTAIL.n32 9.3005
R1409 VTAIL.n18 VTAIL.n17 9.3005
R1410 VTAIL.n57 VTAIL.n56 9.3005
R1411 VTAIL.n59 VTAIL.n58 9.3005
R1412 VTAIL.n14 VTAIL.n13 9.3005
R1413 VTAIL.n65 VTAIL.n64 9.3005
R1414 VTAIL.n67 VTAIL.n66 9.3005
R1415 VTAIL.n10 VTAIL.n9 9.3005
R1416 VTAIL.n74 VTAIL.n73 9.3005
R1417 VTAIL.n76 VTAIL.n75 9.3005
R1418 VTAIL.n246 VTAIL.n245 9.3005
R1419 VTAIL.n248 VTAIL.n247 9.3005
R1420 VTAIL.n203 VTAIL.n202 9.3005
R1421 VTAIL.n254 VTAIL.n253 9.3005
R1422 VTAIL.n256 VTAIL.n255 9.3005
R1423 VTAIL.n198 VTAIL.n197 9.3005
R1424 VTAIL.n262 VTAIL.n261 9.3005
R1425 VTAIL.n264 VTAIL.n263 9.3005
R1426 VTAIL.n279 VTAIL.n278 9.3005
R1427 VTAIL.n190 VTAIL.n189 9.3005
R1428 VTAIL.n273 VTAIL.n272 9.3005
R1429 VTAIL.n271 VTAIL.n270 9.3005
R1430 VTAIL.n194 VTAIL.n193 9.3005
R1431 VTAIL.n207 VTAIL.n206 9.3005
R1432 VTAIL.n240 VTAIL.n239 9.3005
R1433 VTAIL.n238 VTAIL.n237 9.3005
R1434 VTAIL.n211 VTAIL.n210 9.3005
R1435 VTAIL.n232 VTAIL.n231 9.3005
R1436 VTAIL.n230 VTAIL.n229 9.3005
R1437 VTAIL.n215 VTAIL.n214 9.3005
R1438 VTAIL.n224 VTAIL.n223 9.3005
R1439 VTAIL.n222 VTAIL.n221 9.3005
R1440 VTAIL.n152 VTAIL.n151 9.3005
R1441 VTAIL.n154 VTAIL.n153 9.3005
R1442 VTAIL.n109 VTAIL.n108 9.3005
R1443 VTAIL.n160 VTAIL.n159 9.3005
R1444 VTAIL.n162 VTAIL.n161 9.3005
R1445 VTAIL.n104 VTAIL.n103 9.3005
R1446 VTAIL.n168 VTAIL.n167 9.3005
R1447 VTAIL.n170 VTAIL.n169 9.3005
R1448 VTAIL.n185 VTAIL.n184 9.3005
R1449 VTAIL.n96 VTAIL.n95 9.3005
R1450 VTAIL.n179 VTAIL.n178 9.3005
R1451 VTAIL.n177 VTAIL.n176 9.3005
R1452 VTAIL.n100 VTAIL.n99 9.3005
R1453 VTAIL.n113 VTAIL.n112 9.3005
R1454 VTAIL.n146 VTAIL.n145 9.3005
R1455 VTAIL.n144 VTAIL.n143 9.3005
R1456 VTAIL.n117 VTAIL.n116 9.3005
R1457 VTAIL.n138 VTAIL.n137 9.3005
R1458 VTAIL.n136 VTAIL.n135 9.3005
R1459 VTAIL.n121 VTAIL.n120 9.3005
R1460 VTAIL.n130 VTAIL.n129 9.3005
R1461 VTAIL.n128 VTAIL.n127 9.3005
R1462 VTAIL.n329 VTAIL.n304 8.92171
R1463 VTAIL.n342 VTAIL.n296 8.92171
R1464 VTAIL.n47 VTAIL.n22 8.92171
R1465 VTAIL.n60 VTAIL.n14 8.92171
R1466 VTAIL.n249 VTAIL.n203 8.92171
R1467 VTAIL.n236 VTAIL.n211 8.92171
R1468 VTAIL.n155 VTAIL.n109 8.92171
R1469 VTAIL.n142 VTAIL.n117 8.92171
R1470 VTAIL.n330 VTAIL.n302 8.14595
R1471 VTAIL.n341 VTAIL.n298 8.14595
R1472 VTAIL.n48 VTAIL.n20 8.14595
R1473 VTAIL.n59 VTAIL.n16 8.14595
R1474 VTAIL.n248 VTAIL.n205 8.14595
R1475 VTAIL.n237 VTAIL.n209 8.14595
R1476 VTAIL.n154 VTAIL.n111 8.14595
R1477 VTAIL.n143 VTAIL.n115 8.14595
R1478 VTAIL.n334 VTAIL.n333 7.3702
R1479 VTAIL.n338 VTAIL.n337 7.3702
R1480 VTAIL.n52 VTAIL.n51 7.3702
R1481 VTAIL.n56 VTAIL.n55 7.3702
R1482 VTAIL.n245 VTAIL.n244 7.3702
R1483 VTAIL.n241 VTAIL.n240 7.3702
R1484 VTAIL.n151 VTAIL.n150 7.3702
R1485 VTAIL.n147 VTAIL.n146 7.3702
R1486 VTAIL.n334 VTAIL.n300 6.59444
R1487 VTAIL.n337 VTAIL.n300 6.59444
R1488 VTAIL.n52 VTAIL.n18 6.59444
R1489 VTAIL.n55 VTAIL.n18 6.59444
R1490 VTAIL.n244 VTAIL.n207 6.59444
R1491 VTAIL.n241 VTAIL.n207 6.59444
R1492 VTAIL.n150 VTAIL.n113 6.59444
R1493 VTAIL.n147 VTAIL.n113 6.59444
R1494 VTAIL.n333 VTAIL.n302 5.81868
R1495 VTAIL.n338 VTAIL.n298 5.81868
R1496 VTAIL.n51 VTAIL.n20 5.81868
R1497 VTAIL.n56 VTAIL.n16 5.81868
R1498 VTAIL.n245 VTAIL.n205 5.81868
R1499 VTAIL.n240 VTAIL.n209 5.81868
R1500 VTAIL.n151 VTAIL.n111 5.81868
R1501 VTAIL.n146 VTAIL.n115 5.81868
R1502 VTAIL.n330 VTAIL.n329 5.04292
R1503 VTAIL.n342 VTAIL.n341 5.04292
R1504 VTAIL.n48 VTAIL.n47 5.04292
R1505 VTAIL.n60 VTAIL.n59 5.04292
R1506 VTAIL.n249 VTAIL.n248 5.04292
R1507 VTAIL.n237 VTAIL.n236 5.04292
R1508 VTAIL.n155 VTAIL.n154 5.04292
R1509 VTAIL.n143 VTAIL.n142 5.04292
R1510 VTAIL.n326 VTAIL.n304 4.26717
R1511 VTAIL.n345 VTAIL.n296 4.26717
R1512 VTAIL.n374 VTAIL.n282 4.26717
R1513 VTAIL.n44 VTAIL.n22 4.26717
R1514 VTAIL.n63 VTAIL.n14 4.26717
R1515 VTAIL.n92 VTAIL.n0 4.26717
R1516 VTAIL.n280 VTAIL.n188 4.26717
R1517 VTAIL.n252 VTAIL.n203 4.26717
R1518 VTAIL.n233 VTAIL.n211 4.26717
R1519 VTAIL.n186 VTAIL.n94 4.26717
R1520 VTAIL.n158 VTAIL.n109 4.26717
R1521 VTAIL.n139 VTAIL.n117 4.26717
R1522 VTAIL.n315 VTAIL.n311 3.70982
R1523 VTAIL.n33 VTAIL.n29 3.70982
R1524 VTAIL.n222 VTAIL.n218 3.70982
R1525 VTAIL.n128 VTAIL.n124 3.70982
R1526 VTAIL.n325 VTAIL.n306 3.49141
R1527 VTAIL.n346 VTAIL.n294 3.49141
R1528 VTAIL.n372 VTAIL.n371 3.49141
R1529 VTAIL.n43 VTAIL.n24 3.49141
R1530 VTAIL.n64 VTAIL.n12 3.49141
R1531 VTAIL.n90 VTAIL.n89 3.49141
R1532 VTAIL.n278 VTAIL.n277 3.49141
R1533 VTAIL.n253 VTAIL.n201 3.49141
R1534 VTAIL.n232 VTAIL.n213 3.49141
R1535 VTAIL.n184 VTAIL.n183 3.49141
R1536 VTAIL.n159 VTAIL.n107 3.49141
R1537 VTAIL.n138 VTAIL.n119 3.49141
R1538 VTAIL.n322 VTAIL.n321 2.71565
R1539 VTAIL.n350 VTAIL.n349 2.71565
R1540 VTAIL.n368 VTAIL.n284 2.71565
R1541 VTAIL.n40 VTAIL.n39 2.71565
R1542 VTAIL.n68 VTAIL.n67 2.71565
R1543 VTAIL.n86 VTAIL.n2 2.71565
R1544 VTAIL.n274 VTAIL.n190 2.71565
R1545 VTAIL.n257 VTAIL.n256 2.71565
R1546 VTAIL.n229 VTAIL.n228 2.71565
R1547 VTAIL.n180 VTAIL.n96 2.71565
R1548 VTAIL.n163 VTAIL.n162 2.71565
R1549 VTAIL.n135 VTAIL.n134 2.71565
R1550 VTAIL.n281 VTAIL.n187 2.0436
R1551 VTAIL.n318 VTAIL.n308 1.93989
R1552 VTAIL.n354 VTAIL.n292 1.93989
R1553 VTAIL.n367 VTAIL.n286 1.93989
R1554 VTAIL.n36 VTAIL.n26 1.93989
R1555 VTAIL.n72 VTAIL.n10 1.93989
R1556 VTAIL.n85 VTAIL.n4 1.93989
R1557 VTAIL.n273 VTAIL.n192 1.93989
R1558 VTAIL.n260 VTAIL.n198 1.93989
R1559 VTAIL.n225 VTAIL.n215 1.93989
R1560 VTAIL.n179 VTAIL.n98 1.93989
R1561 VTAIL.n166 VTAIL.n104 1.93989
R1562 VTAIL.n131 VTAIL.n121 1.93989
R1563 VTAIL VTAIL.n93 1.31516
R1564 VTAIL.n317 VTAIL.n310 1.16414
R1565 VTAIL.n355 VTAIL.n290 1.16414
R1566 VTAIL.n364 VTAIL.n363 1.16414
R1567 VTAIL.n35 VTAIL.n28 1.16414
R1568 VTAIL.n73 VTAIL.n8 1.16414
R1569 VTAIL.n82 VTAIL.n81 1.16414
R1570 VTAIL.n270 VTAIL.n269 1.16414
R1571 VTAIL.n261 VTAIL.n196 1.16414
R1572 VTAIL.n224 VTAIL.n217 1.16414
R1573 VTAIL.n176 VTAIL.n175 1.16414
R1574 VTAIL.n167 VTAIL.n102 1.16414
R1575 VTAIL.n130 VTAIL.n123 1.16414
R1576 VTAIL VTAIL.n375 0.728948
R1577 VTAIL.n314 VTAIL.n313 0.388379
R1578 VTAIL.n359 VTAIL.n358 0.388379
R1579 VTAIL.n360 VTAIL.n288 0.388379
R1580 VTAIL.n32 VTAIL.n31 0.388379
R1581 VTAIL.n77 VTAIL.n76 0.388379
R1582 VTAIL.n78 VTAIL.n6 0.388379
R1583 VTAIL.n266 VTAIL.n194 0.388379
R1584 VTAIL.n265 VTAIL.n264 0.388379
R1585 VTAIL.n221 VTAIL.n220 0.388379
R1586 VTAIL.n172 VTAIL.n100 0.388379
R1587 VTAIL.n171 VTAIL.n170 0.388379
R1588 VTAIL.n127 VTAIL.n126 0.388379
R1589 VTAIL.n316 VTAIL.n315 0.155672
R1590 VTAIL.n316 VTAIL.n307 0.155672
R1591 VTAIL.n323 VTAIL.n307 0.155672
R1592 VTAIL.n324 VTAIL.n323 0.155672
R1593 VTAIL.n324 VTAIL.n303 0.155672
R1594 VTAIL.n331 VTAIL.n303 0.155672
R1595 VTAIL.n332 VTAIL.n331 0.155672
R1596 VTAIL.n332 VTAIL.n299 0.155672
R1597 VTAIL.n339 VTAIL.n299 0.155672
R1598 VTAIL.n340 VTAIL.n339 0.155672
R1599 VTAIL.n340 VTAIL.n295 0.155672
R1600 VTAIL.n347 VTAIL.n295 0.155672
R1601 VTAIL.n348 VTAIL.n347 0.155672
R1602 VTAIL.n348 VTAIL.n291 0.155672
R1603 VTAIL.n356 VTAIL.n291 0.155672
R1604 VTAIL.n357 VTAIL.n356 0.155672
R1605 VTAIL.n357 VTAIL.n287 0.155672
R1606 VTAIL.n365 VTAIL.n287 0.155672
R1607 VTAIL.n366 VTAIL.n365 0.155672
R1608 VTAIL.n366 VTAIL.n283 0.155672
R1609 VTAIL.n373 VTAIL.n283 0.155672
R1610 VTAIL.n34 VTAIL.n33 0.155672
R1611 VTAIL.n34 VTAIL.n25 0.155672
R1612 VTAIL.n41 VTAIL.n25 0.155672
R1613 VTAIL.n42 VTAIL.n41 0.155672
R1614 VTAIL.n42 VTAIL.n21 0.155672
R1615 VTAIL.n49 VTAIL.n21 0.155672
R1616 VTAIL.n50 VTAIL.n49 0.155672
R1617 VTAIL.n50 VTAIL.n17 0.155672
R1618 VTAIL.n57 VTAIL.n17 0.155672
R1619 VTAIL.n58 VTAIL.n57 0.155672
R1620 VTAIL.n58 VTAIL.n13 0.155672
R1621 VTAIL.n65 VTAIL.n13 0.155672
R1622 VTAIL.n66 VTAIL.n65 0.155672
R1623 VTAIL.n66 VTAIL.n9 0.155672
R1624 VTAIL.n74 VTAIL.n9 0.155672
R1625 VTAIL.n75 VTAIL.n74 0.155672
R1626 VTAIL.n75 VTAIL.n5 0.155672
R1627 VTAIL.n83 VTAIL.n5 0.155672
R1628 VTAIL.n84 VTAIL.n83 0.155672
R1629 VTAIL.n84 VTAIL.n1 0.155672
R1630 VTAIL.n91 VTAIL.n1 0.155672
R1631 VTAIL.n279 VTAIL.n189 0.155672
R1632 VTAIL.n272 VTAIL.n189 0.155672
R1633 VTAIL.n272 VTAIL.n271 0.155672
R1634 VTAIL.n271 VTAIL.n193 0.155672
R1635 VTAIL.n263 VTAIL.n193 0.155672
R1636 VTAIL.n263 VTAIL.n262 0.155672
R1637 VTAIL.n262 VTAIL.n197 0.155672
R1638 VTAIL.n255 VTAIL.n197 0.155672
R1639 VTAIL.n255 VTAIL.n254 0.155672
R1640 VTAIL.n254 VTAIL.n202 0.155672
R1641 VTAIL.n247 VTAIL.n202 0.155672
R1642 VTAIL.n247 VTAIL.n246 0.155672
R1643 VTAIL.n246 VTAIL.n206 0.155672
R1644 VTAIL.n239 VTAIL.n206 0.155672
R1645 VTAIL.n239 VTAIL.n238 0.155672
R1646 VTAIL.n238 VTAIL.n210 0.155672
R1647 VTAIL.n231 VTAIL.n210 0.155672
R1648 VTAIL.n231 VTAIL.n230 0.155672
R1649 VTAIL.n230 VTAIL.n214 0.155672
R1650 VTAIL.n223 VTAIL.n214 0.155672
R1651 VTAIL.n223 VTAIL.n222 0.155672
R1652 VTAIL.n185 VTAIL.n95 0.155672
R1653 VTAIL.n178 VTAIL.n95 0.155672
R1654 VTAIL.n178 VTAIL.n177 0.155672
R1655 VTAIL.n177 VTAIL.n99 0.155672
R1656 VTAIL.n169 VTAIL.n99 0.155672
R1657 VTAIL.n169 VTAIL.n168 0.155672
R1658 VTAIL.n168 VTAIL.n103 0.155672
R1659 VTAIL.n161 VTAIL.n103 0.155672
R1660 VTAIL.n161 VTAIL.n160 0.155672
R1661 VTAIL.n160 VTAIL.n108 0.155672
R1662 VTAIL.n153 VTAIL.n108 0.155672
R1663 VTAIL.n153 VTAIL.n152 0.155672
R1664 VTAIL.n152 VTAIL.n112 0.155672
R1665 VTAIL.n145 VTAIL.n112 0.155672
R1666 VTAIL.n145 VTAIL.n144 0.155672
R1667 VTAIL.n144 VTAIL.n116 0.155672
R1668 VTAIL.n137 VTAIL.n116 0.155672
R1669 VTAIL.n137 VTAIL.n136 0.155672
R1670 VTAIL.n136 VTAIL.n120 0.155672
R1671 VTAIL.n129 VTAIL.n120 0.155672
R1672 VTAIL.n129 VTAIL.n128 0.155672
R1673 VDD2.n181 VDD2.n93 756.745
R1674 VDD2.n88 VDD2.n0 756.745
R1675 VDD2.n182 VDD2.n181 585
R1676 VDD2.n180 VDD2.n179 585
R1677 VDD2.n97 VDD2.n96 585
R1678 VDD2.n174 VDD2.n173 585
R1679 VDD2.n172 VDD2.n171 585
R1680 VDD2.n170 VDD2.n100 585
R1681 VDD2.n104 VDD2.n101 585
R1682 VDD2.n165 VDD2.n164 585
R1683 VDD2.n163 VDD2.n162 585
R1684 VDD2.n106 VDD2.n105 585
R1685 VDD2.n157 VDD2.n156 585
R1686 VDD2.n155 VDD2.n154 585
R1687 VDD2.n110 VDD2.n109 585
R1688 VDD2.n149 VDD2.n148 585
R1689 VDD2.n147 VDD2.n146 585
R1690 VDD2.n114 VDD2.n113 585
R1691 VDD2.n141 VDD2.n140 585
R1692 VDD2.n139 VDD2.n138 585
R1693 VDD2.n118 VDD2.n117 585
R1694 VDD2.n133 VDD2.n132 585
R1695 VDD2.n131 VDD2.n130 585
R1696 VDD2.n122 VDD2.n121 585
R1697 VDD2.n125 VDD2.n124 585
R1698 VDD2.n31 VDD2.n30 585
R1699 VDD2.n28 VDD2.n27 585
R1700 VDD2.n37 VDD2.n36 585
R1701 VDD2.n39 VDD2.n38 585
R1702 VDD2.n24 VDD2.n23 585
R1703 VDD2.n45 VDD2.n44 585
R1704 VDD2.n47 VDD2.n46 585
R1705 VDD2.n20 VDD2.n19 585
R1706 VDD2.n53 VDD2.n52 585
R1707 VDD2.n55 VDD2.n54 585
R1708 VDD2.n16 VDD2.n15 585
R1709 VDD2.n61 VDD2.n60 585
R1710 VDD2.n63 VDD2.n62 585
R1711 VDD2.n12 VDD2.n11 585
R1712 VDD2.n69 VDD2.n68 585
R1713 VDD2.n72 VDD2.n71 585
R1714 VDD2.n70 VDD2.n8 585
R1715 VDD2.n77 VDD2.n7 585
R1716 VDD2.n79 VDD2.n78 585
R1717 VDD2.n81 VDD2.n80 585
R1718 VDD2.n4 VDD2.n3 585
R1719 VDD2.n87 VDD2.n86 585
R1720 VDD2.n89 VDD2.n88 585
R1721 VDD2.t1 VDD2.n123 327.466
R1722 VDD2.t0 VDD2.n29 327.466
R1723 VDD2.n181 VDD2.n180 171.744
R1724 VDD2.n180 VDD2.n96 171.744
R1725 VDD2.n173 VDD2.n96 171.744
R1726 VDD2.n173 VDD2.n172 171.744
R1727 VDD2.n172 VDD2.n100 171.744
R1728 VDD2.n104 VDD2.n100 171.744
R1729 VDD2.n164 VDD2.n104 171.744
R1730 VDD2.n164 VDD2.n163 171.744
R1731 VDD2.n163 VDD2.n105 171.744
R1732 VDD2.n156 VDD2.n105 171.744
R1733 VDD2.n156 VDD2.n155 171.744
R1734 VDD2.n155 VDD2.n109 171.744
R1735 VDD2.n148 VDD2.n109 171.744
R1736 VDD2.n148 VDD2.n147 171.744
R1737 VDD2.n147 VDD2.n113 171.744
R1738 VDD2.n140 VDD2.n113 171.744
R1739 VDD2.n140 VDD2.n139 171.744
R1740 VDD2.n139 VDD2.n117 171.744
R1741 VDD2.n132 VDD2.n117 171.744
R1742 VDD2.n132 VDD2.n131 171.744
R1743 VDD2.n131 VDD2.n121 171.744
R1744 VDD2.n124 VDD2.n121 171.744
R1745 VDD2.n30 VDD2.n27 171.744
R1746 VDD2.n37 VDD2.n27 171.744
R1747 VDD2.n38 VDD2.n37 171.744
R1748 VDD2.n38 VDD2.n23 171.744
R1749 VDD2.n45 VDD2.n23 171.744
R1750 VDD2.n46 VDD2.n45 171.744
R1751 VDD2.n46 VDD2.n19 171.744
R1752 VDD2.n53 VDD2.n19 171.744
R1753 VDD2.n54 VDD2.n53 171.744
R1754 VDD2.n54 VDD2.n15 171.744
R1755 VDD2.n61 VDD2.n15 171.744
R1756 VDD2.n62 VDD2.n61 171.744
R1757 VDD2.n62 VDD2.n11 171.744
R1758 VDD2.n69 VDD2.n11 171.744
R1759 VDD2.n71 VDD2.n69 171.744
R1760 VDD2.n71 VDD2.n70 171.744
R1761 VDD2.n70 VDD2.n7 171.744
R1762 VDD2.n79 VDD2.n7 171.744
R1763 VDD2.n80 VDD2.n79 171.744
R1764 VDD2.n80 VDD2.n3 171.744
R1765 VDD2.n87 VDD2.n3 171.744
R1766 VDD2.n88 VDD2.n87 171.744
R1767 VDD2.n186 VDD2.n92 91.2739
R1768 VDD2.n124 VDD2.t1 85.8723
R1769 VDD2.n30 VDD2.t0 85.8723
R1770 VDD2.n186 VDD2.n185 46.9247
R1771 VDD2.n125 VDD2.n123 16.3895
R1772 VDD2.n31 VDD2.n29 16.3895
R1773 VDD2.n171 VDD2.n170 13.1884
R1774 VDD2.n78 VDD2.n77 13.1884
R1775 VDD2.n174 VDD2.n99 12.8005
R1776 VDD2.n169 VDD2.n101 12.8005
R1777 VDD2.n126 VDD2.n122 12.8005
R1778 VDD2.n32 VDD2.n28 12.8005
R1779 VDD2.n76 VDD2.n8 12.8005
R1780 VDD2.n81 VDD2.n6 12.8005
R1781 VDD2.n175 VDD2.n97 12.0247
R1782 VDD2.n166 VDD2.n165 12.0247
R1783 VDD2.n130 VDD2.n129 12.0247
R1784 VDD2.n36 VDD2.n35 12.0247
R1785 VDD2.n73 VDD2.n72 12.0247
R1786 VDD2.n82 VDD2.n4 12.0247
R1787 VDD2.n179 VDD2.n178 11.249
R1788 VDD2.n162 VDD2.n103 11.249
R1789 VDD2.n133 VDD2.n120 11.249
R1790 VDD2.n39 VDD2.n26 11.249
R1791 VDD2.n68 VDD2.n10 11.249
R1792 VDD2.n86 VDD2.n85 11.249
R1793 VDD2.n182 VDD2.n95 10.4732
R1794 VDD2.n161 VDD2.n106 10.4732
R1795 VDD2.n134 VDD2.n118 10.4732
R1796 VDD2.n40 VDD2.n24 10.4732
R1797 VDD2.n67 VDD2.n12 10.4732
R1798 VDD2.n89 VDD2.n2 10.4732
R1799 VDD2.n183 VDD2.n93 9.69747
R1800 VDD2.n158 VDD2.n157 9.69747
R1801 VDD2.n138 VDD2.n137 9.69747
R1802 VDD2.n44 VDD2.n43 9.69747
R1803 VDD2.n64 VDD2.n63 9.69747
R1804 VDD2.n90 VDD2.n0 9.69747
R1805 VDD2.n185 VDD2.n184 9.45567
R1806 VDD2.n92 VDD2.n91 9.45567
R1807 VDD2.n151 VDD2.n150 9.3005
R1808 VDD2.n153 VDD2.n152 9.3005
R1809 VDD2.n108 VDD2.n107 9.3005
R1810 VDD2.n159 VDD2.n158 9.3005
R1811 VDD2.n161 VDD2.n160 9.3005
R1812 VDD2.n103 VDD2.n102 9.3005
R1813 VDD2.n167 VDD2.n166 9.3005
R1814 VDD2.n169 VDD2.n168 9.3005
R1815 VDD2.n184 VDD2.n183 9.3005
R1816 VDD2.n95 VDD2.n94 9.3005
R1817 VDD2.n178 VDD2.n177 9.3005
R1818 VDD2.n176 VDD2.n175 9.3005
R1819 VDD2.n99 VDD2.n98 9.3005
R1820 VDD2.n112 VDD2.n111 9.3005
R1821 VDD2.n145 VDD2.n144 9.3005
R1822 VDD2.n143 VDD2.n142 9.3005
R1823 VDD2.n116 VDD2.n115 9.3005
R1824 VDD2.n137 VDD2.n136 9.3005
R1825 VDD2.n135 VDD2.n134 9.3005
R1826 VDD2.n120 VDD2.n119 9.3005
R1827 VDD2.n129 VDD2.n128 9.3005
R1828 VDD2.n127 VDD2.n126 9.3005
R1829 VDD2.n91 VDD2.n90 9.3005
R1830 VDD2.n2 VDD2.n1 9.3005
R1831 VDD2.n85 VDD2.n84 9.3005
R1832 VDD2.n83 VDD2.n82 9.3005
R1833 VDD2.n6 VDD2.n5 9.3005
R1834 VDD2.n51 VDD2.n50 9.3005
R1835 VDD2.n49 VDD2.n48 9.3005
R1836 VDD2.n22 VDD2.n21 9.3005
R1837 VDD2.n43 VDD2.n42 9.3005
R1838 VDD2.n41 VDD2.n40 9.3005
R1839 VDD2.n26 VDD2.n25 9.3005
R1840 VDD2.n35 VDD2.n34 9.3005
R1841 VDD2.n33 VDD2.n32 9.3005
R1842 VDD2.n18 VDD2.n17 9.3005
R1843 VDD2.n57 VDD2.n56 9.3005
R1844 VDD2.n59 VDD2.n58 9.3005
R1845 VDD2.n14 VDD2.n13 9.3005
R1846 VDD2.n65 VDD2.n64 9.3005
R1847 VDD2.n67 VDD2.n66 9.3005
R1848 VDD2.n10 VDD2.n9 9.3005
R1849 VDD2.n74 VDD2.n73 9.3005
R1850 VDD2.n76 VDD2.n75 9.3005
R1851 VDD2.n154 VDD2.n108 8.92171
R1852 VDD2.n141 VDD2.n116 8.92171
R1853 VDD2.n47 VDD2.n22 8.92171
R1854 VDD2.n60 VDD2.n14 8.92171
R1855 VDD2.n153 VDD2.n110 8.14595
R1856 VDD2.n142 VDD2.n114 8.14595
R1857 VDD2.n48 VDD2.n20 8.14595
R1858 VDD2.n59 VDD2.n16 8.14595
R1859 VDD2.n150 VDD2.n149 7.3702
R1860 VDD2.n146 VDD2.n145 7.3702
R1861 VDD2.n52 VDD2.n51 7.3702
R1862 VDD2.n56 VDD2.n55 7.3702
R1863 VDD2.n149 VDD2.n112 6.59444
R1864 VDD2.n146 VDD2.n112 6.59444
R1865 VDD2.n52 VDD2.n18 6.59444
R1866 VDD2.n55 VDD2.n18 6.59444
R1867 VDD2.n150 VDD2.n110 5.81868
R1868 VDD2.n145 VDD2.n114 5.81868
R1869 VDD2.n51 VDD2.n20 5.81868
R1870 VDD2.n56 VDD2.n16 5.81868
R1871 VDD2.n154 VDD2.n153 5.04292
R1872 VDD2.n142 VDD2.n141 5.04292
R1873 VDD2.n48 VDD2.n47 5.04292
R1874 VDD2.n60 VDD2.n59 5.04292
R1875 VDD2.n185 VDD2.n93 4.26717
R1876 VDD2.n157 VDD2.n108 4.26717
R1877 VDD2.n138 VDD2.n116 4.26717
R1878 VDD2.n44 VDD2.n22 4.26717
R1879 VDD2.n63 VDD2.n14 4.26717
R1880 VDD2.n92 VDD2.n0 4.26717
R1881 VDD2.n127 VDD2.n123 3.70982
R1882 VDD2.n33 VDD2.n29 3.70982
R1883 VDD2.n183 VDD2.n182 3.49141
R1884 VDD2.n158 VDD2.n106 3.49141
R1885 VDD2.n137 VDD2.n118 3.49141
R1886 VDD2.n43 VDD2.n24 3.49141
R1887 VDD2.n64 VDD2.n12 3.49141
R1888 VDD2.n90 VDD2.n89 3.49141
R1889 VDD2.n179 VDD2.n95 2.71565
R1890 VDD2.n162 VDD2.n161 2.71565
R1891 VDD2.n134 VDD2.n133 2.71565
R1892 VDD2.n40 VDD2.n39 2.71565
R1893 VDD2.n68 VDD2.n67 2.71565
R1894 VDD2.n86 VDD2.n2 2.71565
R1895 VDD2.n178 VDD2.n97 1.93989
R1896 VDD2.n165 VDD2.n103 1.93989
R1897 VDD2.n130 VDD2.n120 1.93989
R1898 VDD2.n36 VDD2.n26 1.93989
R1899 VDD2.n72 VDD2.n10 1.93989
R1900 VDD2.n85 VDD2.n4 1.93989
R1901 VDD2.n175 VDD2.n174 1.16414
R1902 VDD2.n166 VDD2.n101 1.16414
R1903 VDD2.n129 VDD2.n122 1.16414
R1904 VDD2.n35 VDD2.n28 1.16414
R1905 VDD2.n73 VDD2.n8 1.16414
R1906 VDD2.n82 VDD2.n81 1.16414
R1907 VDD2 VDD2.n186 0.845328
R1908 VDD2.n171 VDD2.n99 0.388379
R1909 VDD2.n170 VDD2.n169 0.388379
R1910 VDD2.n126 VDD2.n125 0.388379
R1911 VDD2.n32 VDD2.n31 0.388379
R1912 VDD2.n77 VDD2.n76 0.388379
R1913 VDD2.n78 VDD2.n6 0.388379
R1914 VDD2.n184 VDD2.n94 0.155672
R1915 VDD2.n177 VDD2.n94 0.155672
R1916 VDD2.n177 VDD2.n176 0.155672
R1917 VDD2.n176 VDD2.n98 0.155672
R1918 VDD2.n168 VDD2.n98 0.155672
R1919 VDD2.n168 VDD2.n167 0.155672
R1920 VDD2.n167 VDD2.n102 0.155672
R1921 VDD2.n160 VDD2.n102 0.155672
R1922 VDD2.n160 VDD2.n159 0.155672
R1923 VDD2.n159 VDD2.n107 0.155672
R1924 VDD2.n152 VDD2.n107 0.155672
R1925 VDD2.n152 VDD2.n151 0.155672
R1926 VDD2.n151 VDD2.n111 0.155672
R1927 VDD2.n144 VDD2.n111 0.155672
R1928 VDD2.n144 VDD2.n143 0.155672
R1929 VDD2.n143 VDD2.n115 0.155672
R1930 VDD2.n136 VDD2.n115 0.155672
R1931 VDD2.n136 VDD2.n135 0.155672
R1932 VDD2.n135 VDD2.n119 0.155672
R1933 VDD2.n128 VDD2.n119 0.155672
R1934 VDD2.n128 VDD2.n127 0.155672
R1935 VDD2.n34 VDD2.n33 0.155672
R1936 VDD2.n34 VDD2.n25 0.155672
R1937 VDD2.n41 VDD2.n25 0.155672
R1938 VDD2.n42 VDD2.n41 0.155672
R1939 VDD2.n42 VDD2.n21 0.155672
R1940 VDD2.n49 VDD2.n21 0.155672
R1941 VDD2.n50 VDD2.n49 0.155672
R1942 VDD2.n50 VDD2.n17 0.155672
R1943 VDD2.n57 VDD2.n17 0.155672
R1944 VDD2.n58 VDD2.n57 0.155672
R1945 VDD2.n58 VDD2.n13 0.155672
R1946 VDD2.n65 VDD2.n13 0.155672
R1947 VDD2.n66 VDD2.n65 0.155672
R1948 VDD2.n66 VDD2.n9 0.155672
R1949 VDD2.n74 VDD2.n9 0.155672
R1950 VDD2.n75 VDD2.n74 0.155672
R1951 VDD2.n75 VDD2.n5 0.155672
R1952 VDD2.n83 VDD2.n5 0.155672
R1953 VDD2.n84 VDD2.n83 0.155672
R1954 VDD2.n84 VDD2.n1 0.155672
R1955 VDD2.n91 VDD2.n1 0.155672
R1956 VP.n0 VP.t1 210.198
R1957 VP.n0 VP.t0 160.072
R1958 VP VP.n0 0.526373
R1959 VDD1.n88 VDD1.n0 756.745
R1960 VDD1.n181 VDD1.n93 756.745
R1961 VDD1.n89 VDD1.n88 585
R1962 VDD1.n87 VDD1.n86 585
R1963 VDD1.n4 VDD1.n3 585
R1964 VDD1.n81 VDD1.n80 585
R1965 VDD1.n79 VDD1.n78 585
R1966 VDD1.n77 VDD1.n7 585
R1967 VDD1.n11 VDD1.n8 585
R1968 VDD1.n72 VDD1.n71 585
R1969 VDD1.n70 VDD1.n69 585
R1970 VDD1.n13 VDD1.n12 585
R1971 VDD1.n64 VDD1.n63 585
R1972 VDD1.n62 VDD1.n61 585
R1973 VDD1.n17 VDD1.n16 585
R1974 VDD1.n56 VDD1.n55 585
R1975 VDD1.n54 VDD1.n53 585
R1976 VDD1.n21 VDD1.n20 585
R1977 VDD1.n48 VDD1.n47 585
R1978 VDD1.n46 VDD1.n45 585
R1979 VDD1.n25 VDD1.n24 585
R1980 VDD1.n40 VDD1.n39 585
R1981 VDD1.n38 VDD1.n37 585
R1982 VDD1.n29 VDD1.n28 585
R1983 VDD1.n32 VDD1.n31 585
R1984 VDD1.n124 VDD1.n123 585
R1985 VDD1.n121 VDD1.n120 585
R1986 VDD1.n130 VDD1.n129 585
R1987 VDD1.n132 VDD1.n131 585
R1988 VDD1.n117 VDD1.n116 585
R1989 VDD1.n138 VDD1.n137 585
R1990 VDD1.n140 VDD1.n139 585
R1991 VDD1.n113 VDD1.n112 585
R1992 VDD1.n146 VDD1.n145 585
R1993 VDD1.n148 VDD1.n147 585
R1994 VDD1.n109 VDD1.n108 585
R1995 VDD1.n154 VDD1.n153 585
R1996 VDD1.n156 VDD1.n155 585
R1997 VDD1.n105 VDD1.n104 585
R1998 VDD1.n162 VDD1.n161 585
R1999 VDD1.n165 VDD1.n164 585
R2000 VDD1.n163 VDD1.n101 585
R2001 VDD1.n170 VDD1.n100 585
R2002 VDD1.n172 VDD1.n171 585
R2003 VDD1.n174 VDD1.n173 585
R2004 VDD1.n97 VDD1.n96 585
R2005 VDD1.n180 VDD1.n179 585
R2006 VDD1.n182 VDD1.n181 585
R2007 VDD1.t0 VDD1.n30 327.466
R2008 VDD1.t1 VDD1.n122 327.466
R2009 VDD1.n88 VDD1.n87 171.744
R2010 VDD1.n87 VDD1.n3 171.744
R2011 VDD1.n80 VDD1.n3 171.744
R2012 VDD1.n80 VDD1.n79 171.744
R2013 VDD1.n79 VDD1.n7 171.744
R2014 VDD1.n11 VDD1.n7 171.744
R2015 VDD1.n71 VDD1.n11 171.744
R2016 VDD1.n71 VDD1.n70 171.744
R2017 VDD1.n70 VDD1.n12 171.744
R2018 VDD1.n63 VDD1.n12 171.744
R2019 VDD1.n63 VDD1.n62 171.744
R2020 VDD1.n62 VDD1.n16 171.744
R2021 VDD1.n55 VDD1.n16 171.744
R2022 VDD1.n55 VDD1.n54 171.744
R2023 VDD1.n54 VDD1.n20 171.744
R2024 VDD1.n47 VDD1.n20 171.744
R2025 VDD1.n47 VDD1.n46 171.744
R2026 VDD1.n46 VDD1.n24 171.744
R2027 VDD1.n39 VDD1.n24 171.744
R2028 VDD1.n39 VDD1.n38 171.744
R2029 VDD1.n38 VDD1.n28 171.744
R2030 VDD1.n31 VDD1.n28 171.744
R2031 VDD1.n123 VDD1.n120 171.744
R2032 VDD1.n130 VDD1.n120 171.744
R2033 VDD1.n131 VDD1.n130 171.744
R2034 VDD1.n131 VDD1.n116 171.744
R2035 VDD1.n138 VDD1.n116 171.744
R2036 VDD1.n139 VDD1.n138 171.744
R2037 VDD1.n139 VDD1.n112 171.744
R2038 VDD1.n146 VDD1.n112 171.744
R2039 VDD1.n147 VDD1.n146 171.744
R2040 VDD1.n147 VDD1.n108 171.744
R2041 VDD1.n154 VDD1.n108 171.744
R2042 VDD1.n155 VDD1.n154 171.744
R2043 VDD1.n155 VDD1.n104 171.744
R2044 VDD1.n162 VDD1.n104 171.744
R2045 VDD1.n164 VDD1.n162 171.744
R2046 VDD1.n164 VDD1.n163 171.744
R2047 VDD1.n163 VDD1.n100 171.744
R2048 VDD1.n172 VDD1.n100 171.744
R2049 VDD1.n173 VDD1.n172 171.744
R2050 VDD1.n173 VDD1.n96 171.744
R2051 VDD1.n180 VDD1.n96 171.744
R2052 VDD1.n181 VDD1.n180 171.744
R2053 VDD1 VDD1.n185 92.5853
R2054 VDD1.n31 VDD1.t0 85.8723
R2055 VDD1.n123 VDD1.t1 85.8723
R2056 VDD1 VDD1.n92 47.7696
R2057 VDD1.n32 VDD1.n30 16.3895
R2058 VDD1.n124 VDD1.n122 16.3895
R2059 VDD1.n78 VDD1.n77 13.1884
R2060 VDD1.n171 VDD1.n170 13.1884
R2061 VDD1.n81 VDD1.n6 12.8005
R2062 VDD1.n76 VDD1.n8 12.8005
R2063 VDD1.n33 VDD1.n29 12.8005
R2064 VDD1.n125 VDD1.n121 12.8005
R2065 VDD1.n169 VDD1.n101 12.8005
R2066 VDD1.n174 VDD1.n99 12.8005
R2067 VDD1.n82 VDD1.n4 12.0247
R2068 VDD1.n73 VDD1.n72 12.0247
R2069 VDD1.n37 VDD1.n36 12.0247
R2070 VDD1.n129 VDD1.n128 12.0247
R2071 VDD1.n166 VDD1.n165 12.0247
R2072 VDD1.n175 VDD1.n97 12.0247
R2073 VDD1.n86 VDD1.n85 11.249
R2074 VDD1.n69 VDD1.n10 11.249
R2075 VDD1.n40 VDD1.n27 11.249
R2076 VDD1.n132 VDD1.n119 11.249
R2077 VDD1.n161 VDD1.n103 11.249
R2078 VDD1.n179 VDD1.n178 11.249
R2079 VDD1.n89 VDD1.n2 10.4732
R2080 VDD1.n68 VDD1.n13 10.4732
R2081 VDD1.n41 VDD1.n25 10.4732
R2082 VDD1.n133 VDD1.n117 10.4732
R2083 VDD1.n160 VDD1.n105 10.4732
R2084 VDD1.n182 VDD1.n95 10.4732
R2085 VDD1.n90 VDD1.n0 9.69747
R2086 VDD1.n65 VDD1.n64 9.69747
R2087 VDD1.n45 VDD1.n44 9.69747
R2088 VDD1.n137 VDD1.n136 9.69747
R2089 VDD1.n157 VDD1.n156 9.69747
R2090 VDD1.n183 VDD1.n93 9.69747
R2091 VDD1.n92 VDD1.n91 9.45567
R2092 VDD1.n185 VDD1.n184 9.45567
R2093 VDD1.n58 VDD1.n57 9.3005
R2094 VDD1.n60 VDD1.n59 9.3005
R2095 VDD1.n15 VDD1.n14 9.3005
R2096 VDD1.n66 VDD1.n65 9.3005
R2097 VDD1.n68 VDD1.n67 9.3005
R2098 VDD1.n10 VDD1.n9 9.3005
R2099 VDD1.n74 VDD1.n73 9.3005
R2100 VDD1.n76 VDD1.n75 9.3005
R2101 VDD1.n91 VDD1.n90 9.3005
R2102 VDD1.n2 VDD1.n1 9.3005
R2103 VDD1.n85 VDD1.n84 9.3005
R2104 VDD1.n83 VDD1.n82 9.3005
R2105 VDD1.n6 VDD1.n5 9.3005
R2106 VDD1.n19 VDD1.n18 9.3005
R2107 VDD1.n52 VDD1.n51 9.3005
R2108 VDD1.n50 VDD1.n49 9.3005
R2109 VDD1.n23 VDD1.n22 9.3005
R2110 VDD1.n44 VDD1.n43 9.3005
R2111 VDD1.n42 VDD1.n41 9.3005
R2112 VDD1.n27 VDD1.n26 9.3005
R2113 VDD1.n36 VDD1.n35 9.3005
R2114 VDD1.n34 VDD1.n33 9.3005
R2115 VDD1.n184 VDD1.n183 9.3005
R2116 VDD1.n95 VDD1.n94 9.3005
R2117 VDD1.n178 VDD1.n177 9.3005
R2118 VDD1.n176 VDD1.n175 9.3005
R2119 VDD1.n99 VDD1.n98 9.3005
R2120 VDD1.n144 VDD1.n143 9.3005
R2121 VDD1.n142 VDD1.n141 9.3005
R2122 VDD1.n115 VDD1.n114 9.3005
R2123 VDD1.n136 VDD1.n135 9.3005
R2124 VDD1.n134 VDD1.n133 9.3005
R2125 VDD1.n119 VDD1.n118 9.3005
R2126 VDD1.n128 VDD1.n127 9.3005
R2127 VDD1.n126 VDD1.n125 9.3005
R2128 VDD1.n111 VDD1.n110 9.3005
R2129 VDD1.n150 VDD1.n149 9.3005
R2130 VDD1.n152 VDD1.n151 9.3005
R2131 VDD1.n107 VDD1.n106 9.3005
R2132 VDD1.n158 VDD1.n157 9.3005
R2133 VDD1.n160 VDD1.n159 9.3005
R2134 VDD1.n103 VDD1.n102 9.3005
R2135 VDD1.n167 VDD1.n166 9.3005
R2136 VDD1.n169 VDD1.n168 9.3005
R2137 VDD1.n61 VDD1.n15 8.92171
R2138 VDD1.n48 VDD1.n23 8.92171
R2139 VDD1.n140 VDD1.n115 8.92171
R2140 VDD1.n153 VDD1.n107 8.92171
R2141 VDD1.n60 VDD1.n17 8.14595
R2142 VDD1.n49 VDD1.n21 8.14595
R2143 VDD1.n141 VDD1.n113 8.14595
R2144 VDD1.n152 VDD1.n109 8.14595
R2145 VDD1.n57 VDD1.n56 7.3702
R2146 VDD1.n53 VDD1.n52 7.3702
R2147 VDD1.n145 VDD1.n144 7.3702
R2148 VDD1.n149 VDD1.n148 7.3702
R2149 VDD1.n56 VDD1.n19 6.59444
R2150 VDD1.n53 VDD1.n19 6.59444
R2151 VDD1.n145 VDD1.n111 6.59444
R2152 VDD1.n148 VDD1.n111 6.59444
R2153 VDD1.n57 VDD1.n17 5.81868
R2154 VDD1.n52 VDD1.n21 5.81868
R2155 VDD1.n144 VDD1.n113 5.81868
R2156 VDD1.n149 VDD1.n109 5.81868
R2157 VDD1.n61 VDD1.n60 5.04292
R2158 VDD1.n49 VDD1.n48 5.04292
R2159 VDD1.n141 VDD1.n140 5.04292
R2160 VDD1.n153 VDD1.n152 5.04292
R2161 VDD1.n92 VDD1.n0 4.26717
R2162 VDD1.n64 VDD1.n15 4.26717
R2163 VDD1.n45 VDD1.n23 4.26717
R2164 VDD1.n137 VDD1.n115 4.26717
R2165 VDD1.n156 VDD1.n107 4.26717
R2166 VDD1.n185 VDD1.n93 4.26717
R2167 VDD1.n34 VDD1.n30 3.70982
R2168 VDD1.n126 VDD1.n122 3.70982
R2169 VDD1.n90 VDD1.n89 3.49141
R2170 VDD1.n65 VDD1.n13 3.49141
R2171 VDD1.n44 VDD1.n25 3.49141
R2172 VDD1.n136 VDD1.n117 3.49141
R2173 VDD1.n157 VDD1.n105 3.49141
R2174 VDD1.n183 VDD1.n182 3.49141
R2175 VDD1.n86 VDD1.n2 2.71565
R2176 VDD1.n69 VDD1.n68 2.71565
R2177 VDD1.n41 VDD1.n40 2.71565
R2178 VDD1.n133 VDD1.n132 2.71565
R2179 VDD1.n161 VDD1.n160 2.71565
R2180 VDD1.n179 VDD1.n95 2.71565
R2181 VDD1.n85 VDD1.n4 1.93989
R2182 VDD1.n72 VDD1.n10 1.93989
R2183 VDD1.n37 VDD1.n27 1.93989
R2184 VDD1.n129 VDD1.n119 1.93989
R2185 VDD1.n165 VDD1.n103 1.93989
R2186 VDD1.n178 VDD1.n97 1.93989
R2187 VDD1.n82 VDD1.n81 1.16414
R2188 VDD1.n73 VDD1.n8 1.16414
R2189 VDD1.n36 VDD1.n29 1.16414
R2190 VDD1.n128 VDD1.n121 1.16414
R2191 VDD1.n166 VDD1.n101 1.16414
R2192 VDD1.n175 VDD1.n174 1.16414
R2193 VDD1.n78 VDD1.n6 0.388379
R2194 VDD1.n77 VDD1.n76 0.388379
R2195 VDD1.n33 VDD1.n32 0.388379
R2196 VDD1.n125 VDD1.n124 0.388379
R2197 VDD1.n170 VDD1.n169 0.388379
R2198 VDD1.n171 VDD1.n99 0.388379
R2199 VDD1.n91 VDD1.n1 0.155672
R2200 VDD1.n84 VDD1.n1 0.155672
R2201 VDD1.n84 VDD1.n83 0.155672
R2202 VDD1.n83 VDD1.n5 0.155672
R2203 VDD1.n75 VDD1.n5 0.155672
R2204 VDD1.n75 VDD1.n74 0.155672
R2205 VDD1.n74 VDD1.n9 0.155672
R2206 VDD1.n67 VDD1.n9 0.155672
R2207 VDD1.n67 VDD1.n66 0.155672
R2208 VDD1.n66 VDD1.n14 0.155672
R2209 VDD1.n59 VDD1.n14 0.155672
R2210 VDD1.n59 VDD1.n58 0.155672
R2211 VDD1.n58 VDD1.n18 0.155672
R2212 VDD1.n51 VDD1.n18 0.155672
R2213 VDD1.n51 VDD1.n50 0.155672
R2214 VDD1.n50 VDD1.n22 0.155672
R2215 VDD1.n43 VDD1.n22 0.155672
R2216 VDD1.n43 VDD1.n42 0.155672
R2217 VDD1.n42 VDD1.n26 0.155672
R2218 VDD1.n35 VDD1.n26 0.155672
R2219 VDD1.n35 VDD1.n34 0.155672
R2220 VDD1.n127 VDD1.n126 0.155672
R2221 VDD1.n127 VDD1.n118 0.155672
R2222 VDD1.n134 VDD1.n118 0.155672
R2223 VDD1.n135 VDD1.n134 0.155672
R2224 VDD1.n135 VDD1.n114 0.155672
R2225 VDD1.n142 VDD1.n114 0.155672
R2226 VDD1.n143 VDD1.n142 0.155672
R2227 VDD1.n143 VDD1.n110 0.155672
R2228 VDD1.n150 VDD1.n110 0.155672
R2229 VDD1.n151 VDD1.n150 0.155672
R2230 VDD1.n151 VDD1.n106 0.155672
R2231 VDD1.n158 VDD1.n106 0.155672
R2232 VDD1.n159 VDD1.n158 0.155672
R2233 VDD1.n159 VDD1.n102 0.155672
R2234 VDD1.n167 VDD1.n102 0.155672
R2235 VDD1.n168 VDD1.n167 0.155672
R2236 VDD1.n168 VDD1.n98 0.155672
R2237 VDD1.n176 VDD1.n98 0.155672
R2238 VDD1.n177 VDD1.n176 0.155672
R2239 VDD1.n177 VDD1.n94 0.155672
R2240 VDD1.n184 VDD1.n94 0.155672
C0 VDD1 VDD2 0.76283f
C1 VN VDD1 0.148787f
C2 B VTAIL 5.02664f
C3 B w_n2430_n4308# 10.904401f
C4 VN VDD2 3.90234f
C5 VTAIL VDD1 6.39223f
C6 B VP 1.74485f
C7 VDD1 w_n2430_n4308# 2.18508f
C8 VTAIL VDD2 6.44747f
C9 VN VTAIL 3.3974f
C10 VDD2 w_n2430_n4308# 2.21989f
C11 VN w_n2430_n4308# 3.5143f
C12 VP VDD1 4.11461f
C13 VP VDD2 0.363955f
C14 VP VN 6.66215f
C15 VTAIL w_n2430_n4308# 3.40127f
C16 B VDD1 2.17826f
C17 B VDD2 2.21474f
C18 VP VTAIL 3.41169f
C19 B VN 1.23052f
C20 VP w_n2430_n4308# 3.82539f
C21 VDD2 VSUBS 1.153672f
C22 VDD1 VSUBS 5.666619f
C23 VTAIL VSUBS 1.263411f
C24 VN VSUBS 8.99157f
C25 VP VSUBS 2.067739f
C26 B VSUBS 4.835219f
C27 w_n2430_n4308# VSUBS 0.128158p
C28 VDD1.n0 VSUBS 0.029202f
C29 VDD1.n1 VSUBS 0.028677f
C30 VDD1.n2 VSUBS 0.01541f
C31 VDD1.n3 VSUBS 0.036423f
C32 VDD1.n4 VSUBS 0.016316f
C33 VDD1.n5 VSUBS 0.028677f
C34 VDD1.n6 VSUBS 0.01541f
C35 VDD1.n7 VSUBS 0.036423f
C36 VDD1.n8 VSUBS 0.016316f
C37 VDD1.n9 VSUBS 0.028677f
C38 VDD1.n10 VSUBS 0.01541f
C39 VDD1.n11 VSUBS 0.036423f
C40 VDD1.n12 VSUBS 0.036423f
C41 VDD1.n13 VSUBS 0.016316f
C42 VDD1.n14 VSUBS 0.028677f
C43 VDD1.n15 VSUBS 0.01541f
C44 VDD1.n16 VSUBS 0.036423f
C45 VDD1.n17 VSUBS 0.016316f
C46 VDD1.n18 VSUBS 0.028677f
C47 VDD1.n19 VSUBS 0.01541f
C48 VDD1.n20 VSUBS 0.036423f
C49 VDD1.n21 VSUBS 0.016316f
C50 VDD1.n22 VSUBS 0.028677f
C51 VDD1.n23 VSUBS 0.01541f
C52 VDD1.n24 VSUBS 0.036423f
C53 VDD1.n25 VSUBS 0.016316f
C54 VDD1.n26 VSUBS 0.028677f
C55 VDD1.n27 VSUBS 0.01541f
C56 VDD1.n28 VSUBS 0.036423f
C57 VDD1.n29 VSUBS 0.016316f
C58 VDD1.n30 VSUBS 0.216529f
C59 VDD1.t0 VSUBS 0.078096f
C60 VDD1.n31 VSUBS 0.027317f
C61 VDD1.n32 VSUBS 0.023171f
C62 VDD1.n33 VSUBS 0.01541f
C63 VDD1.n34 VSUBS 2.05241f
C64 VDD1.n35 VSUBS 0.028677f
C65 VDD1.n36 VSUBS 0.01541f
C66 VDD1.n37 VSUBS 0.016316f
C67 VDD1.n38 VSUBS 0.036423f
C68 VDD1.n39 VSUBS 0.036423f
C69 VDD1.n40 VSUBS 0.016316f
C70 VDD1.n41 VSUBS 0.01541f
C71 VDD1.n42 VSUBS 0.028677f
C72 VDD1.n43 VSUBS 0.028677f
C73 VDD1.n44 VSUBS 0.01541f
C74 VDD1.n45 VSUBS 0.016316f
C75 VDD1.n46 VSUBS 0.036423f
C76 VDD1.n47 VSUBS 0.036423f
C77 VDD1.n48 VSUBS 0.016316f
C78 VDD1.n49 VSUBS 0.01541f
C79 VDD1.n50 VSUBS 0.028677f
C80 VDD1.n51 VSUBS 0.028677f
C81 VDD1.n52 VSUBS 0.01541f
C82 VDD1.n53 VSUBS 0.016316f
C83 VDD1.n54 VSUBS 0.036423f
C84 VDD1.n55 VSUBS 0.036423f
C85 VDD1.n56 VSUBS 0.016316f
C86 VDD1.n57 VSUBS 0.01541f
C87 VDD1.n58 VSUBS 0.028677f
C88 VDD1.n59 VSUBS 0.028677f
C89 VDD1.n60 VSUBS 0.01541f
C90 VDD1.n61 VSUBS 0.016316f
C91 VDD1.n62 VSUBS 0.036423f
C92 VDD1.n63 VSUBS 0.036423f
C93 VDD1.n64 VSUBS 0.016316f
C94 VDD1.n65 VSUBS 0.01541f
C95 VDD1.n66 VSUBS 0.028677f
C96 VDD1.n67 VSUBS 0.028677f
C97 VDD1.n68 VSUBS 0.01541f
C98 VDD1.n69 VSUBS 0.016316f
C99 VDD1.n70 VSUBS 0.036423f
C100 VDD1.n71 VSUBS 0.036423f
C101 VDD1.n72 VSUBS 0.016316f
C102 VDD1.n73 VSUBS 0.01541f
C103 VDD1.n74 VSUBS 0.028677f
C104 VDD1.n75 VSUBS 0.028677f
C105 VDD1.n76 VSUBS 0.01541f
C106 VDD1.n77 VSUBS 0.015863f
C107 VDD1.n78 VSUBS 0.015863f
C108 VDD1.n79 VSUBS 0.036423f
C109 VDD1.n80 VSUBS 0.036423f
C110 VDD1.n81 VSUBS 0.016316f
C111 VDD1.n82 VSUBS 0.01541f
C112 VDD1.n83 VSUBS 0.028677f
C113 VDD1.n84 VSUBS 0.028677f
C114 VDD1.n85 VSUBS 0.01541f
C115 VDD1.n86 VSUBS 0.016316f
C116 VDD1.n87 VSUBS 0.036423f
C117 VDD1.n88 VSUBS 0.080315f
C118 VDD1.n89 VSUBS 0.016316f
C119 VDD1.n90 VSUBS 0.01541f
C120 VDD1.n91 VSUBS 0.062368f
C121 VDD1.n92 VSUBS 0.062069f
C122 VDD1.n93 VSUBS 0.029202f
C123 VDD1.n94 VSUBS 0.028677f
C124 VDD1.n95 VSUBS 0.01541f
C125 VDD1.n96 VSUBS 0.036423f
C126 VDD1.n97 VSUBS 0.016316f
C127 VDD1.n98 VSUBS 0.028677f
C128 VDD1.n99 VSUBS 0.01541f
C129 VDD1.n100 VSUBS 0.036423f
C130 VDD1.n101 VSUBS 0.016316f
C131 VDD1.n102 VSUBS 0.028677f
C132 VDD1.n103 VSUBS 0.01541f
C133 VDD1.n104 VSUBS 0.036423f
C134 VDD1.n105 VSUBS 0.016316f
C135 VDD1.n106 VSUBS 0.028677f
C136 VDD1.n107 VSUBS 0.01541f
C137 VDD1.n108 VSUBS 0.036423f
C138 VDD1.n109 VSUBS 0.016316f
C139 VDD1.n110 VSUBS 0.028677f
C140 VDD1.n111 VSUBS 0.01541f
C141 VDD1.n112 VSUBS 0.036423f
C142 VDD1.n113 VSUBS 0.016316f
C143 VDD1.n114 VSUBS 0.028677f
C144 VDD1.n115 VSUBS 0.01541f
C145 VDD1.n116 VSUBS 0.036423f
C146 VDD1.n117 VSUBS 0.016316f
C147 VDD1.n118 VSUBS 0.028677f
C148 VDD1.n119 VSUBS 0.01541f
C149 VDD1.n120 VSUBS 0.036423f
C150 VDD1.n121 VSUBS 0.016316f
C151 VDD1.n122 VSUBS 0.216529f
C152 VDD1.t1 VSUBS 0.078096f
C153 VDD1.n123 VSUBS 0.027317f
C154 VDD1.n124 VSUBS 0.023171f
C155 VDD1.n125 VSUBS 0.01541f
C156 VDD1.n126 VSUBS 2.05242f
C157 VDD1.n127 VSUBS 0.028677f
C158 VDD1.n128 VSUBS 0.01541f
C159 VDD1.n129 VSUBS 0.016316f
C160 VDD1.n130 VSUBS 0.036423f
C161 VDD1.n131 VSUBS 0.036423f
C162 VDD1.n132 VSUBS 0.016316f
C163 VDD1.n133 VSUBS 0.01541f
C164 VDD1.n134 VSUBS 0.028677f
C165 VDD1.n135 VSUBS 0.028677f
C166 VDD1.n136 VSUBS 0.01541f
C167 VDD1.n137 VSUBS 0.016316f
C168 VDD1.n138 VSUBS 0.036423f
C169 VDD1.n139 VSUBS 0.036423f
C170 VDD1.n140 VSUBS 0.016316f
C171 VDD1.n141 VSUBS 0.01541f
C172 VDD1.n142 VSUBS 0.028677f
C173 VDD1.n143 VSUBS 0.028677f
C174 VDD1.n144 VSUBS 0.01541f
C175 VDD1.n145 VSUBS 0.016316f
C176 VDD1.n146 VSUBS 0.036423f
C177 VDD1.n147 VSUBS 0.036423f
C178 VDD1.n148 VSUBS 0.016316f
C179 VDD1.n149 VSUBS 0.01541f
C180 VDD1.n150 VSUBS 0.028677f
C181 VDD1.n151 VSUBS 0.028677f
C182 VDD1.n152 VSUBS 0.01541f
C183 VDD1.n153 VSUBS 0.016316f
C184 VDD1.n154 VSUBS 0.036423f
C185 VDD1.n155 VSUBS 0.036423f
C186 VDD1.n156 VSUBS 0.016316f
C187 VDD1.n157 VSUBS 0.01541f
C188 VDD1.n158 VSUBS 0.028677f
C189 VDD1.n159 VSUBS 0.028677f
C190 VDD1.n160 VSUBS 0.01541f
C191 VDD1.n161 VSUBS 0.016316f
C192 VDD1.n162 VSUBS 0.036423f
C193 VDD1.n163 VSUBS 0.036423f
C194 VDD1.n164 VSUBS 0.036423f
C195 VDD1.n165 VSUBS 0.016316f
C196 VDD1.n166 VSUBS 0.01541f
C197 VDD1.n167 VSUBS 0.028677f
C198 VDD1.n168 VSUBS 0.028677f
C199 VDD1.n169 VSUBS 0.01541f
C200 VDD1.n170 VSUBS 0.015863f
C201 VDD1.n171 VSUBS 0.015863f
C202 VDD1.n172 VSUBS 0.036423f
C203 VDD1.n173 VSUBS 0.036423f
C204 VDD1.n174 VSUBS 0.016316f
C205 VDD1.n175 VSUBS 0.01541f
C206 VDD1.n176 VSUBS 0.028677f
C207 VDD1.n177 VSUBS 0.028677f
C208 VDD1.n178 VSUBS 0.01541f
C209 VDD1.n179 VSUBS 0.016316f
C210 VDD1.n180 VSUBS 0.036423f
C211 VDD1.n181 VSUBS 0.080315f
C212 VDD1.n182 VSUBS 0.016316f
C213 VDD1.n183 VSUBS 0.01541f
C214 VDD1.n184 VSUBS 0.062368f
C215 VDD1.n185 VSUBS 1.18706f
C216 VP.t1 VSUBS 6.30382f
C217 VP.t0 VSUBS 5.46319f
C218 VP.n0 VSUBS 6.11776f
C219 VDD2.n0 VSUBS 0.029016f
C220 VDD2.n1 VSUBS 0.028495f
C221 VDD2.n2 VSUBS 0.015312f
C222 VDD2.n3 VSUBS 0.036192f
C223 VDD2.n4 VSUBS 0.016213f
C224 VDD2.n5 VSUBS 0.028495f
C225 VDD2.n6 VSUBS 0.015312f
C226 VDD2.n7 VSUBS 0.036192f
C227 VDD2.n8 VSUBS 0.016213f
C228 VDD2.n9 VSUBS 0.028495f
C229 VDD2.n10 VSUBS 0.015312f
C230 VDD2.n11 VSUBS 0.036192f
C231 VDD2.n12 VSUBS 0.016213f
C232 VDD2.n13 VSUBS 0.028495f
C233 VDD2.n14 VSUBS 0.015312f
C234 VDD2.n15 VSUBS 0.036192f
C235 VDD2.n16 VSUBS 0.016213f
C236 VDD2.n17 VSUBS 0.028495f
C237 VDD2.n18 VSUBS 0.015312f
C238 VDD2.n19 VSUBS 0.036192f
C239 VDD2.n20 VSUBS 0.016213f
C240 VDD2.n21 VSUBS 0.028495f
C241 VDD2.n22 VSUBS 0.015312f
C242 VDD2.n23 VSUBS 0.036192f
C243 VDD2.n24 VSUBS 0.016213f
C244 VDD2.n25 VSUBS 0.028495f
C245 VDD2.n26 VSUBS 0.015312f
C246 VDD2.n27 VSUBS 0.036192f
C247 VDD2.n28 VSUBS 0.016213f
C248 VDD2.n29 VSUBS 0.215152f
C249 VDD2.t0 VSUBS 0.0776f
C250 VDD2.n30 VSUBS 0.027144f
C251 VDD2.n31 VSUBS 0.023024f
C252 VDD2.n32 VSUBS 0.015312f
C253 VDD2.n33 VSUBS 2.03936f
C254 VDD2.n34 VSUBS 0.028495f
C255 VDD2.n35 VSUBS 0.015312f
C256 VDD2.n36 VSUBS 0.016213f
C257 VDD2.n37 VSUBS 0.036192f
C258 VDD2.n38 VSUBS 0.036192f
C259 VDD2.n39 VSUBS 0.016213f
C260 VDD2.n40 VSUBS 0.015312f
C261 VDD2.n41 VSUBS 0.028495f
C262 VDD2.n42 VSUBS 0.028495f
C263 VDD2.n43 VSUBS 0.015312f
C264 VDD2.n44 VSUBS 0.016213f
C265 VDD2.n45 VSUBS 0.036192f
C266 VDD2.n46 VSUBS 0.036192f
C267 VDD2.n47 VSUBS 0.016213f
C268 VDD2.n48 VSUBS 0.015312f
C269 VDD2.n49 VSUBS 0.028495f
C270 VDD2.n50 VSUBS 0.028495f
C271 VDD2.n51 VSUBS 0.015312f
C272 VDD2.n52 VSUBS 0.016213f
C273 VDD2.n53 VSUBS 0.036192f
C274 VDD2.n54 VSUBS 0.036192f
C275 VDD2.n55 VSUBS 0.016213f
C276 VDD2.n56 VSUBS 0.015312f
C277 VDD2.n57 VSUBS 0.028495f
C278 VDD2.n58 VSUBS 0.028495f
C279 VDD2.n59 VSUBS 0.015312f
C280 VDD2.n60 VSUBS 0.016213f
C281 VDD2.n61 VSUBS 0.036192f
C282 VDD2.n62 VSUBS 0.036192f
C283 VDD2.n63 VSUBS 0.016213f
C284 VDD2.n64 VSUBS 0.015312f
C285 VDD2.n65 VSUBS 0.028495f
C286 VDD2.n66 VSUBS 0.028495f
C287 VDD2.n67 VSUBS 0.015312f
C288 VDD2.n68 VSUBS 0.016213f
C289 VDD2.n69 VSUBS 0.036192f
C290 VDD2.n70 VSUBS 0.036192f
C291 VDD2.n71 VSUBS 0.036192f
C292 VDD2.n72 VSUBS 0.016213f
C293 VDD2.n73 VSUBS 0.015312f
C294 VDD2.n74 VSUBS 0.028495f
C295 VDD2.n75 VSUBS 0.028495f
C296 VDD2.n76 VSUBS 0.015312f
C297 VDD2.n77 VSUBS 0.015762f
C298 VDD2.n78 VSUBS 0.015762f
C299 VDD2.n79 VSUBS 0.036192f
C300 VDD2.n80 VSUBS 0.036192f
C301 VDD2.n81 VSUBS 0.016213f
C302 VDD2.n82 VSUBS 0.015312f
C303 VDD2.n83 VSUBS 0.028495f
C304 VDD2.n84 VSUBS 0.028495f
C305 VDD2.n85 VSUBS 0.015312f
C306 VDD2.n86 VSUBS 0.016213f
C307 VDD2.n87 VSUBS 0.036192f
C308 VDD2.n88 VSUBS 0.079805f
C309 VDD2.n89 VSUBS 0.016213f
C310 VDD2.n90 VSUBS 0.015312f
C311 VDD2.n91 VSUBS 0.061972f
C312 VDD2.n92 VSUBS 1.11037f
C313 VDD2.n93 VSUBS 0.029016f
C314 VDD2.n94 VSUBS 0.028495f
C315 VDD2.n95 VSUBS 0.015312f
C316 VDD2.n96 VSUBS 0.036192f
C317 VDD2.n97 VSUBS 0.016213f
C318 VDD2.n98 VSUBS 0.028495f
C319 VDD2.n99 VSUBS 0.015312f
C320 VDD2.n100 VSUBS 0.036192f
C321 VDD2.n101 VSUBS 0.016213f
C322 VDD2.n102 VSUBS 0.028495f
C323 VDD2.n103 VSUBS 0.015312f
C324 VDD2.n104 VSUBS 0.036192f
C325 VDD2.n105 VSUBS 0.036192f
C326 VDD2.n106 VSUBS 0.016213f
C327 VDD2.n107 VSUBS 0.028495f
C328 VDD2.n108 VSUBS 0.015312f
C329 VDD2.n109 VSUBS 0.036192f
C330 VDD2.n110 VSUBS 0.016213f
C331 VDD2.n111 VSUBS 0.028495f
C332 VDD2.n112 VSUBS 0.015312f
C333 VDD2.n113 VSUBS 0.036192f
C334 VDD2.n114 VSUBS 0.016213f
C335 VDD2.n115 VSUBS 0.028495f
C336 VDD2.n116 VSUBS 0.015312f
C337 VDD2.n117 VSUBS 0.036192f
C338 VDD2.n118 VSUBS 0.016213f
C339 VDD2.n119 VSUBS 0.028495f
C340 VDD2.n120 VSUBS 0.015312f
C341 VDD2.n121 VSUBS 0.036192f
C342 VDD2.n122 VSUBS 0.016213f
C343 VDD2.n123 VSUBS 0.215152f
C344 VDD2.t1 VSUBS 0.0776f
C345 VDD2.n124 VSUBS 0.027144f
C346 VDD2.n125 VSUBS 0.023024f
C347 VDD2.n126 VSUBS 0.015312f
C348 VDD2.n127 VSUBS 2.03936f
C349 VDD2.n128 VSUBS 0.028495f
C350 VDD2.n129 VSUBS 0.015312f
C351 VDD2.n130 VSUBS 0.016213f
C352 VDD2.n131 VSUBS 0.036192f
C353 VDD2.n132 VSUBS 0.036192f
C354 VDD2.n133 VSUBS 0.016213f
C355 VDD2.n134 VSUBS 0.015312f
C356 VDD2.n135 VSUBS 0.028495f
C357 VDD2.n136 VSUBS 0.028495f
C358 VDD2.n137 VSUBS 0.015312f
C359 VDD2.n138 VSUBS 0.016213f
C360 VDD2.n139 VSUBS 0.036192f
C361 VDD2.n140 VSUBS 0.036192f
C362 VDD2.n141 VSUBS 0.016213f
C363 VDD2.n142 VSUBS 0.015312f
C364 VDD2.n143 VSUBS 0.028495f
C365 VDD2.n144 VSUBS 0.028495f
C366 VDD2.n145 VSUBS 0.015312f
C367 VDD2.n146 VSUBS 0.016213f
C368 VDD2.n147 VSUBS 0.036192f
C369 VDD2.n148 VSUBS 0.036192f
C370 VDD2.n149 VSUBS 0.016213f
C371 VDD2.n150 VSUBS 0.015312f
C372 VDD2.n151 VSUBS 0.028495f
C373 VDD2.n152 VSUBS 0.028495f
C374 VDD2.n153 VSUBS 0.015312f
C375 VDD2.n154 VSUBS 0.016213f
C376 VDD2.n155 VSUBS 0.036192f
C377 VDD2.n156 VSUBS 0.036192f
C378 VDD2.n157 VSUBS 0.016213f
C379 VDD2.n158 VSUBS 0.015312f
C380 VDD2.n159 VSUBS 0.028495f
C381 VDD2.n160 VSUBS 0.028495f
C382 VDD2.n161 VSUBS 0.015312f
C383 VDD2.n162 VSUBS 0.016213f
C384 VDD2.n163 VSUBS 0.036192f
C385 VDD2.n164 VSUBS 0.036192f
C386 VDD2.n165 VSUBS 0.016213f
C387 VDD2.n166 VSUBS 0.015312f
C388 VDD2.n167 VSUBS 0.028495f
C389 VDD2.n168 VSUBS 0.028495f
C390 VDD2.n169 VSUBS 0.015312f
C391 VDD2.n170 VSUBS 0.015762f
C392 VDD2.n171 VSUBS 0.015762f
C393 VDD2.n172 VSUBS 0.036192f
C394 VDD2.n173 VSUBS 0.036192f
C395 VDD2.n174 VSUBS 0.016213f
C396 VDD2.n175 VSUBS 0.015312f
C397 VDD2.n176 VSUBS 0.028495f
C398 VDD2.n177 VSUBS 0.028495f
C399 VDD2.n178 VSUBS 0.015312f
C400 VDD2.n179 VSUBS 0.016213f
C401 VDD2.n180 VSUBS 0.036192f
C402 VDD2.n181 VSUBS 0.079805f
C403 VDD2.n182 VSUBS 0.016213f
C404 VDD2.n183 VSUBS 0.015312f
C405 VDD2.n184 VSUBS 0.061972f
C406 VDD2.n185 VSUBS 0.059371f
C407 VDD2.n186 VSUBS 4.15617f
C408 VTAIL.n0 VSUBS 0.029153f
C409 VTAIL.n1 VSUBS 0.028629f
C410 VTAIL.n2 VSUBS 0.015384f
C411 VTAIL.n3 VSUBS 0.036362f
C412 VTAIL.n4 VSUBS 0.016289f
C413 VTAIL.n5 VSUBS 0.028629f
C414 VTAIL.n6 VSUBS 0.015384f
C415 VTAIL.n7 VSUBS 0.036362f
C416 VTAIL.n8 VSUBS 0.016289f
C417 VTAIL.n9 VSUBS 0.028629f
C418 VTAIL.n10 VSUBS 0.015384f
C419 VTAIL.n11 VSUBS 0.036362f
C420 VTAIL.n12 VSUBS 0.016289f
C421 VTAIL.n13 VSUBS 0.028629f
C422 VTAIL.n14 VSUBS 0.015384f
C423 VTAIL.n15 VSUBS 0.036362f
C424 VTAIL.n16 VSUBS 0.016289f
C425 VTAIL.n17 VSUBS 0.028629f
C426 VTAIL.n18 VSUBS 0.015384f
C427 VTAIL.n19 VSUBS 0.036362f
C428 VTAIL.n20 VSUBS 0.016289f
C429 VTAIL.n21 VSUBS 0.028629f
C430 VTAIL.n22 VSUBS 0.015384f
C431 VTAIL.n23 VSUBS 0.036362f
C432 VTAIL.n24 VSUBS 0.016289f
C433 VTAIL.n25 VSUBS 0.028629f
C434 VTAIL.n26 VSUBS 0.015384f
C435 VTAIL.n27 VSUBS 0.036362f
C436 VTAIL.n28 VSUBS 0.016289f
C437 VTAIL.n29 VSUBS 0.216161f
C438 VTAIL.t3 VSUBS 0.077964f
C439 VTAIL.n30 VSUBS 0.027271f
C440 VTAIL.n31 VSUBS 0.023132f
C441 VTAIL.n32 VSUBS 0.015384f
C442 VTAIL.n33 VSUBS 2.04893f
C443 VTAIL.n34 VSUBS 0.028629f
C444 VTAIL.n35 VSUBS 0.015384f
C445 VTAIL.n36 VSUBS 0.016289f
C446 VTAIL.n37 VSUBS 0.036362f
C447 VTAIL.n38 VSUBS 0.036362f
C448 VTAIL.n39 VSUBS 0.016289f
C449 VTAIL.n40 VSUBS 0.015384f
C450 VTAIL.n41 VSUBS 0.028629f
C451 VTAIL.n42 VSUBS 0.028629f
C452 VTAIL.n43 VSUBS 0.015384f
C453 VTAIL.n44 VSUBS 0.016289f
C454 VTAIL.n45 VSUBS 0.036362f
C455 VTAIL.n46 VSUBS 0.036362f
C456 VTAIL.n47 VSUBS 0.016289f
C457 VTAIL.n48 VSUBS 0.015384f
C458 VTAIL.n49 VSUBS 0.028629f
C459 VTAIL.n50 VSUBS 0.028629f
C460 VTAIL.n51 VSUBS 0.015384f
C461 VTAIL.n52 VSUBS 0.016289f
C462 VTAIL.n53 VSUBS 0.036362f
C463 VTAIL.n54 VSUBS 0.036362f
C464 VTAIL.n55 VSUBS 0.016289f
C465 VTAIL.n56 VSUBS 0.015384f
C466 VTAIL.n57 VSUBS 0.028629f
C467 VTAIL.n58 VSUBS 0.028629f
C468 VTAIL.n59 VSUBS 0.015384f
C469 VTAIL.n60 VSUBS 0.016289f
C470 VTAIL.n61 VSUBS 0.036362f
C471 VTAIL.n62 VSUBS 0.036362f
C472 VTAIL.n63 VSUBS 0.016289f
C473 VTAIL.n64 VSUBS 0.015384f
C474 VTAIL.n65 VSUBS 0.028629f
C475 VTAIL.n66 VSUBS 0.028629f
C476 VTAIL.n67 VSUBS 0.015384f
C477 VTAIL.n68 VSUBS 0.016289f
C478 VTAIL.n69 VSUBS 0.036362f
C479 VTAIL.n70 VSUBS 0.036362f
C480 VTAIL.n71 VSUBS 0.036362f
C481 VTAIL.n72 VSUBS 0.016289f
C482 VTAIL.n73 VSUBS 0.015384f
C483 VTAIL.n74 VSUBS 0.028629f
C484 VTAIL.n75 VSUBS 0.028629f
C485 VTAIL.n76 VSUBS 0.015384f
C486 VTAIL.n77 VSUBS 0.015836f
C487 VTAIL.n78 VSUBS 0.015836f
C488 VTAIL.n79 VSUBS 0.036362f
C489 VTAIL.n80 VSUBS 0.036362f
C490 VTAIL.n81 VSUBS 0.016289f
C491 VTAIL.n82 VSUBS 0.015384f
C492 VTAIL.n83 VSUBS 0.028629f
C493 VTAIL.n84 VSUBS 0.028629f
C494 VTAIL.n85 VSUBS 0.015384f
C495 VTAIL.n86 VSUBS 0.016289f
C496 VTAIL.n87 VSUBS 0.036362f
C497 VTAIL.n88 VSUBS 0.080179f
C498 VTAIL.n89 VSUBS 0.016289f
C499 VTAIL.n90 VSUBS 0.015384f
C500 VTAIL.n91 VSUBS 0.062263f
C501 VTAIL.n92 VSUBS 0.039849f
C502 VTAIL.n93 VSUBS 2.44098f
C503 VTAIL.n94 VSUBS 0.029153f
C504 VTAIL.n95 VSUBS 0.028629f
C505 VTAIL.n96 VSUBS 0.015384f
C506 VTAIL.n97 VSUBS 0.036362f
C507 VTAIL.n98 VSUBS 0.016289f
C508 VTAIL.n99 VSUBS 0.028629f
C509 VTAIL.n100 VSUBS 0.015384f
C510 VTAIL.n101 VSUBS 0.036362f
C511 VTAIL.n102 VSUBS 0.016289f
C512 VTAIL.n103 VSUBS 0.028629f
C513 VTAIL.n104 VSUBS 0.015384f
C514 VTAIL.n105 VSUBS 0.036362f
C515 VTAIL.n106 VSUBS 0.036362f
C516 VTAIL.n107 VSUBS 0.016289f
C517 VTAIL.n108 VSUBS 0.028629f
C518 VTAIL.n109 VSUBS 0.015384f
C519 VTAIL.n110 VSUBS 0.036362f
C520 VTAIL.n111 VSUBS 0.016289f
C521 VTAIL.n112 VSUBS 0.028629f
C522 VTAIL.n113 VSUBS 0.015384f
C523 VTAIL.n114 VSUBS 0.036362f
C524 VTAIL.n115 VSUBS 0.016289f
C525 VTAIL.n116 VSUBS 0.028629f
C526 VTAIL.n117 VSUBS 0.015384f
C527 VTAIL.n118 VSUBS 0.036362f
C528 VTAIL.n119 VSUBS 0.016289f
C529 VTAIL.n120 VSUBS 0.028629f
C530 VTAIL.n121 VSUBS 0.015384f
C531 VTAIL.n122 VSUBS 0.036362f
C532 VTAIL.n123 VSUBS 0.016289f
C533 VTAIL.n124 VSUBS 0.216161f
C534 VTAIL.t0 VSUBS 0.077964f
C535 VTAIL.n125 VSUBS 0.027271f
C536 VTAIL.n126 VSUBS 0.023132f
C537 VTAIL.n127 VSUBS 0.015384f
C538 VTAIL.n128 VSUBS 2.04893f
C539 VTAIL.n129 VSUBS 0.028629f
C540 VTAIL.n130 VSUBS 0.015384f
C541 VTAIL.n131 VSUBS 0.016289f
C542 VTAIL.n132 VSUBS 0.036362f
C543 VTAIL.n133 VSUBS 0.036362f
C544 VTAIL.n134 VSUBS 0.016289f
C545 VTAIL.n135 VSUBS 0.015384f
C546 VTAIL.n136 VSUBS 0.028629f
C547 VTAIL.n137 VSUBS 0.028629f
C548 VTAIL.n138 VSUBS 0.015384f
C549 VTAIL.n139 VSUBS 0.016289f
C550 VTAIL.n140 VSUBS 0.036362f
C551 VTAIL.n141 VSUBS 0.036362f
C552 VTAIL.n142 VSUBS 0.016289f
C553 VTAIL.n143 VSUBS 0.015384f
C554 VTAIL.n144 VSUBS 0.028629f
C555 VTAIL.n145 VSUBS 0.028629f
C556 VTAIL.n146 VSUBS 0.015384f
C557 VTAIL.n147 VSUBS 0.016289f
C558 VTAIL.n148 VSUBS 0.036362f
C559 VTAIL.n149 VSUBS 0.036362f
C560 VTAIL.n150 VSUBS 0.016289f
C561 VTAIL.n151 VSUBS 0.015384f
C562 VTAIL.n152 VSUBS 0.028629f
C563 VTAIL.n153 VSUBS 0.028629f
C564 VTAIL.n154 VSUBS 0.015384f
C565 VTAIL.n155 VSUBS 0.016289f
C566 VTAIL.n156 VSUBS 0.036362f
C567 VTAIL.n157 VSUBS 0.036362f
C568 VTAIL.n158 VSUBS 0.016289f
C569 VTAIL.n159 VSUBS 0.015384f
C570 VTAIL.n160 VSUBS 0.028629f
C571 VTAIL.n161 VSUBS 0.028629f
C572 VTAIL.n162 VSUBS 0.015384f
C573 VTAIL.n163 VSUBS 0.016289f
C574 VTAIL.n164 VSUBS 0.036362f
C575 VTAIL.n165 VSUBS 0.036362f
C576 VTAIL.n166 VSUBS 0.016289f
C577 VTAIL.n167 VSUBS 0.015384f
C578 VTAIL.n168 VSUBS 0.028629f
C579 VTAIL.n169 VSUBS 0.028629f
C580 VTAIL.n170 VSUBS 0.015384f
C581 VTAIL.n171 VSUBS 0.015836f
C582 VTAIL.n172 VSUBS 0.015836f
C583 VTAIL.n173 VSUBS 0.036362f
C584 VTAIL.n174 VSUBS 0.036362f
C585 VTAIL.n175 VSUBS 0.016289f
C586 VTAIL.n176 VSUBS 0.015384f
C587 VTAIL.n177 VSUBS 0.028629f
C588 VTAIL.n178 VSUBS 0.028629f
C589 VTAIL.n179 VSUBS 0.015384f
C590 VTAIL.n180 VSUBS 0.016289f
C591 VTAIL.n181 VSUBS 0.036362f
C592 VTAIL.n182 VSUBS 0.080179f
C593 VTAIL.n183 VSUBS 0.016289f
C594 VTAIL.n184 VSUBS 0.015384f
C595 VTAIL.n185 VSUBS 0.062263f
C596 VTAIL.n186 VSUBS 0.039849f
C597 VTAIL.n187 VSUBS 2.50817f
C598 VTAIL.n188 VSUBS 0.029153f
C599 VTAIL.n189 VSUBS 0.028629f
C600 VTAIL.n190 VSUBS 0.015384f
C601 VTAIL.n191 VSUBS 0.036362f
C602 VTAIL.n192 VSUBS 0.016289f
C603 VTAIL.n193 VSUBS 0.028629f
C604 VTAIL.n194 VSUBS 0.015384f
C605 VTAIL.n195 VSUBS 0.036362f
C606 VTAIL.n196 VSUBS 0.016289f
C607 VTAIL.n197 VSUBS 0.028629f
C608 VTAIL.n198 VSUBS 0.015384f
C609 VTAIL.n199 VSUBS 0.036362f
C610 VTAIL.n200 VSUBS 0.036362f
C611 VTAIL.n201 VSUBS 0.016289f
C612 VTAIL.n202 VSUBS 0.028629f
C613 VTAIL.n203 VSUBS 0.015384f
C614 VTAIL.n204 VSUBS 0.036362f
C615 VTAIL.n205 VSUBS 0.016289f
C616 VTAIL.n206 VSUBS 0.028629f
C617 VTAIL.n207 VSUBS 0.015384f
C618 VTAIL.n208 VSUBS 0.036362f
C619 VTAIL.n209 VSUBS 0.016289f
C620 VTAIL.n210 VSUBS 0.028629f
C621 VTAIL.n211 VSUBS 0.015384f
C622 VTAIL.n212 VSUBS 0.036362f
C623 VTAIL.n213 VSUBS 0.016289f
C624 VTAIL.n214 VSUBS 0.028629f
C625 VTAIL.n215 VSUBS 0.015384f
C626 VTAIL.n216 VSUBS 0.036362f
C627 VTAIL.n217 VSUBS 0.016289f
C628 VTAIL.n218 VSUBS 0.216161f
C629 VTAIL.t2 VSUBS 0.077964f
C630 VTAIL.n219 VSUBS 0.027271f
C631 VTAIL.n220 VSUBS 0.023132f
C632 VTAIL.n221 VSUBS 0.015384f
C633 VTAIL.n222 VSUBS 2.04893f
C634 VTAIL.n223 VSUBS 0.028629f
C635 VTAIL.n224 VSUBS 0.015384f
C636 VTAIL.n225 VSUBS 0.016289f
C637 VTAIL.n226 VSUBS 0.036362f
C638 VTAIL.n227 VSUBS 0.036362f
C639 VTAIL.n228 VSUBS 0.016289f
C640 VTAIL.n229 VSUBS 0.015384f
C641 VTAIL.n230 VSUBS 0.028629f
C642 VTAIL.n231 VSUBS 0.028629f
C643 VTAIL.n232 VSUBS 0.015384f
C644 VTAIL.n233 VSUBS 0.016289f
C645 VTAIL.n234 VSUBS 0.036362f
C646 VTAIL.n235 VSUBS 0.036362f
C647 VTAIL.n236 VSUBS 0.016289f
C648 VTAIL.n237 VSUBS 0.015384f
C649 VTAIL.n238 VSUBS 0.028629f
C650 VTAIL.n239 VSUBS 0.028629f
C651 VTAIL.n240 VSUBS 0.015384f
C652 VTAIL.n241 VSUBS 0.016289f
C653 VTAIL.n242 VSUBS 0.036362f
C654 VTAIL.n243 VSUBS 0.036362f
C655 VTAIL.n244 VSUBS 0.016289f
C656 VTAIL.n245 VSUBS 0.015384f
C657 VTAIL.n246 VSUBS 0.028629f
C658 VTAIL.n247 VSUBS 0.028629f
C659 VTAIL.n248 VSUBS 0.015384f
C660 VTAIL.n249 VSUBS 0.016289f
C661 VTAIL.n250 VSUBS 0.036362f
C662 VTAIL.n251 VSUBS 0.036362f
C663 VTAIL.n252 VSUBS 0.016289f
C664 VTAIL.n253 VSUBS 0.015384f
C665 VTAIL.n254 VSUBS 0.028629f
C666 VTAIL.n255 VSUBS 0.028629f
C667 VTAIL.n256 VSUBS 0.015384f
C668 VTAIL.n257 VSUBS 0.016289f
C669 VTAIL.n258 VSUBS 0.036362f
C670 VTAIL.n259 VSUBS 0.036362f
C671 VTAIL.n260 VSUBS 0.016289f
C672 VTAIL.n261 VSUBS 0.015384f
C673 VTAIL.n262 VSUBS 0.028629f
C674 VTAIL.n263 VSUBS 0.028629f
C675 VTAIL.n264 VSUBS 0.015384f
C676 VTAIL.n265 VSUBS 0.015836f
C677 VTAIL.n266 VSUBS 0.015836f
C678 VTAIL.n267 VSUBS 0.036362f
C679 VTAIL.n268 VSUBS 0.036362f
C680 VTAIL.n269 VSUBS 0.016289f
C681 VTAIL.n270 VSUBS 0.015384f
C682 VTAIL.n271 VSUBS 0.028629f
C683 VTAIL.n272 VSUBS 0.028629f
C684 VTAIL.n273 VSUBS 0.015384f
C685 VTAIL.n274 VSUBS 0.016289f
C686 VTAIL.n275 VSUBS 0.036362f
C687 VTAIL.n276 VSUBS 0.080179f
C688 VTAIL.n277 VSUBS 0.016289f
C689 VTAIL.n278 VSUBS 0.015384f
C690 VTAIL.n279 VSUBS 0.062263f
C691 VTAIL.n280 VSUBS 0.039849f
C692 VTAIL.n281 VSUBS 2.21791f
C693 VTAIL.n282 VSUBS 0.029153f
C694 VTAIL.n283 VSUBS 0.028629f
C695 VTAIL.n284 VSUBS 0.015384f
C696 VTAIL.n285 VSUBS 0.036362f
C697 VTAIL.n286 VSUBS 0.016289f
C698 VTAIL.n287 VSUBS 0.028629f
C699 VTAIL.n288 VSUBS 0.015384f
C700 VTAIL.n289 VSUBS 0.036362f
C701 VTAIL.n290 VSUBS 0.016289f
C702 VTAIL.n291 VSUBS 0.028629f
C703 VTAIL.n292 VSUBS 0.015384f
C704 VTAIL.n293 VSUBS 0.036362f
C705 VTAIL.n294 VSUBS 0.016289f
C706 VTAIL.n295 VSUBS 0.028629f
C707 VTAIL.n296 VSUBS 0.015384f
C708 VTAIL.n297 VSUBS 0.036362f
C709 VTAIL.n298 VSUBS 0.016289f
C710 VTAIL.n299 VSUBS 0.028629f
C711 VTAIL.n300 VSUBS 0.015384f
C712 VTAIL.n301 VSUBS 0.036362f
C713 VTAIL.n302 VSUBS 0.016289f
C714 VTAIL.n303 VSUBS 0.028629f
C715 VTAIL.n304 VSUBS 0.015384f
C716 VTAIL.n305 VSUBS 0.036362f
C717 VTAIL.n306 VSUBS 0.016289f
C718 VTAIL.n307 VSUBS 0.028629f
C719 VTAIL.n308 VSUBS 0.015384f
C720 VTAIL.n309 VSUBS 0.036362f
C721 VTAIL.n310 VSUBS 0.016289f
C722 VTAIL.n311 VSUBS 0.216161f
C723 VTAIL.t1 VSUBS 0.077964f
C724 VTAIL.n312 VSUBS 0.027271f
C725 VTAIL.n313 VSUBS 0.023132f
C726 VTAIL.n314 VSUBS 0.015384f
C727 VTAIL.n315 VSUBS 2.04893f
C728 VTAIL.n316 VSUBS 0.028629f
C729 VTAIL.n317 VSUBS 0.015384f
C730 VTAIL.n318 VSUBS 0.016289f
C731 VTAIL.n319 VSUBS 0.036362f
C732 VTAIL.n320 VSUBS 0.036362f
C733 VTAIL.n321 VSUBS 0.016289f
C734 VTAIL.n322 VSUBS 0.015384f
C735 VTAIL.n323 VSUBS 0.028629f
C736 VTAIL.n324 VSUBS 0.028629f
C737 VTAIL.n325 VSUBS 0.015384f
C738 VTAIL.n326 VSUBS 0.016289f
C739 VTAIL.n327 VSUBS 0.036362f
C740 VTAIL.n328 VSUBS 0.036362f
C741 VTAIL.n329 VSUBS 0.016289f
C742 VTAIL.n330 VSUBS 0.015384f
C743 VTAIL.n331 VSUBS 0.028629f
C744 VTAIL.n332 VSUBS 0.028629f
C745 VTAIL.n333 VSUBS 0.015384f
C746 VTAIL.n334 VSUBS 0.016289f
C747 VTAIL.n335 VSUBS 0.036362f
C748 VTAIL.n336 VSUBS 0.036362f
C749 VTAIL.n337 VSUBS 0.016289f
C750 VTAIL.n338 VSUBS 0.015384f
C751 VTAIL.n339 VSUBS 0.028629f
C752 VTAIL.n340 VSUBS 0.028629f
C753 VTAIL.n341 VSUBS 0.015384f
C754 VTAIL.n342 VSUBS 0.016289f
C755 VTAIL.n343 VSUBS 0.036362f
C756 VTAIL.n344 VSUBS 0.036362f
C757 VTAIL.n345 VSUBS 0.016289f
C758 VTAIL.n346 VSUBS 0.015384f
C759 VTAIL.n347 VSUBS 0.028629f
C760 VTAIL.n348 VSUBS 0.028629f
C761 VTAIL.n349 VSUBS 0.015384f
C762 VTAIL.n350 VSUBS 0.016289f
C763 VTAIL.n351 VSUBS 0.036362f
C764 VTAIL.n352 VSUBS 0.036362f
C765 VTAIL.n353 VSUBS 0.036362f
C766 VTAIL.n354 VSUBS 0.016289f
C767 VTAIL.n355 VSUBS 0.015384f
C768 VTAIL.n356 VSUBS 0.028629f
C769 VTAIL.n357 VSUBS 0.028629f
C770 VTAIL.n358 VSUBS 0.015384f
C771 VTAIL.n359 VSUBS 0.015836f
C772 VTAIL.n360 VSUBS 0.015836f
C773 VTAIL.n361 VSUBS 0.036362f
C774 VTAIL.n362 VSUBS 0.036362f
C775 VTAIL.n363 VSUBS 0.016289f
C776 VTAIL.n364 VSUBS 0.015384f
C777 VTAIL.n365 VSUBS 0.028629f
C778 VTAIL.n366 VSUBS 0.028629f
C779 VTAIL.n367 VSUBS 0.015384f
C780 VTAIL.n368 VSUBS 0.016289f
C781 VTAIL.n369 VSUBS 0.036362f
C782 VTAIL.n370 VSUBS 0.080179f
C783 VTAIL.n371 VSUBS 0.016289f
C784 VTAIL.n372 VSUBS 0.015384f
C785 VTAIL.n373 VSUBS 0.062263f
C786 VTAIL.n374 VSUBS 0.039849f
C787 VTAIL.n375 VSUBS 2.09664f
C788 VN.t1 VSUBS 5.30333f
C789 VN.t0 VSUBS 6.11275f
C790 B.n0 VSUBS 0.005806f
C791 B.n1 VSUBS 0.005806f
C792 B.n2 VSUBS 0.008587f
C793 B.n3 VSUBS 0.00658f
C794 B.n4 VSUBS 0.00658f
C795 B.n5 VSUBS 0.00658f
C796 B.n6 VSUBS 0.00658f
C797 B.n7 VSUBS 0.00658f
C798 B.n8 VSUBS 0.00658f
C799 B.n9 VSUBS 0.00658f
C800 B.n10 VSUBS 0.00658f
C801 B.n11 VSUBS 0.00658f
C802 B.n12 VSUBS 0.00658f
C803 B.n13 VSUBS 0.00658f
C804 B.n14 VSUBS 0.00658f
C805 B.n15 VSUBS 0.00658f
C806 B.n16 VSUBS 0.016102f
C807 B.n17 VSUBS 0.00658f
C808 B.n18 VSUBS 0.00658f
C809 B.n19 VSUBS 0.00658f
C810 B.n20 VSUBS 0.00658f
C811 B.n21 VSUBS 0.00658f
C812 B.n22 VSUBS 0.00658f
C813 B.n23 VSUBS 0.00658f
C814 B.n24 VSUBS 0.00658f
C815 B.n25 VSUBS 0.00658f
C816 B.n26 VSUBS 0.00658f
C817 B.n27 VSUBS 0.00658f
C818 B.n28 VSUBS 0.00658f
C819 B.n29 VSUBS 0.00658f
C820 B.n30 VSUBS 0.00658f
C821 B.n31 VSUBS 0.00658f
C822 B.n32 VSUBS 0.00658f
C823 B.n33 VSUBS 0.00658f
C824 B.n34 VSUBS 0.00658f
C825 B.n35 VSUBS 0.00658f
C826 B.n36 VSUBS 0.00658f
C827 B.n37 VSUBS 0.00658f
C828 B.n38 VSUBS 0.00658f
C829 B.n39 VSUBS 0.00658f
C830 B.n40 VSUBS 0.00658f
C831 B.n41 VSUBS 0.00658f
C832 B.n42 VSUBS 0.00658f
C833 B.n43 VSUBS 0.00658f
C834 B.t10 VSUBS 0.300459f
C835 B.t11 VSUBS 0.338833f
C836 B.t9 VSUBS 2.36439f
C837 B.n44 VSUBS 0.535724f
C838 B.n45 VSUBS 0.297174f
C839 B.n46 VSUBS 0.015245f
C840 B.n47 VSUBS 0.00658f
C841 B.n48 VSUBS 0.00658f
C842 B.n49 VSUBS 0.00658f
C843 B.n50 VSUBS 0.00658f
C844 B.n51 VSUBS 0.00658f
C845 B.t1 VSUBS 0.300463f
C846 B.t2 VSUBS 0.338836f
C847 B.t0 VSUBS 2.36439f
C848 B.n52 VSUBS 0.535721f
C849 B.n53 VSUBS 0.297171f
C850 B.n54 VSUBS 0.00658f
C851 B.n55 VSUBS 0.00658f
C852 B.n56 VSUBS 0.00658f
C853 B.n57 VSUBS 0.00658f
C854 B.n58 VSUBS 0.00658f
C855 B.n59 VSUBS 0.00658f
C856 B.n60 VSUBS 0.00658f
C857 B.n61 VSUBS 0.00658f
C858 B.n62 VSUBS 0.00658f
C859 B.n63 VSUBS 0.00658f
C860 B.n64 VSUBS 0.00658f
C861 B.n65 VSUBS 0.00658f
C862 B.n66 VSUBS 0.00658f
C863 B.n67 VSUBS 0.00658f
C864 B.n68 VSUBS 0.00658f
C865 B.n69 VSUBS 0.00658f
C866 B.n70 VSUBS 0.00658f
C867 B.n71 VSUBS 0.00658f
C868 B.n72 VSUBS 0.00658f
C869 B.n73 VSUBS 0.00658f
C870 B.n74 VSUBS 0.00658f
C871 B.n75 VSUBS 0.00658f
C872 B.n76 VSUBS 0.00658f
C873 B.n77 VSUBS 0.00658f
C874 B.n78 VSUBS 0.00658f
C875 B.n79 VSUBS 0.00658f
C876 B.n80 VSUBS 0.00658f
C877 B.n81 VSUBS 0.016102f
C878 B.n82 VSUBS 0.00658f
C879 B.n83 VSUBS 0.00658f
C880 B.n84 VSUBS 0.00658f
C881 B.n85 VSUBS 0.00658f
C882 B.n86 VSUBS 0.00658f
C883 B.n87 VSUBS 0.00658f
C884 B.n88 VSUBS 0.00658f
C885 B.n89 VSUBS 0.00658f
C886 B.n90 VSUBS 0.00658f
C887 B.n91 VSUBS 0.00658f
C888 B.n92 VSUBS 0.00658f
C889 B.n93 VSUBS 0.00658f
C890 B.n94 VSUBS 0.00658f
C891 B.n95 VSUBS 0.00658f
C892 B.n96 VSUBS 0.00658f
C893 B.n97 VSUBS 0.00658f
C894 B.n98 VSUBS 0.00658f
C895 B.n99 VSUBS 0.00658f
C896 B.n100 VSUBS 0.00658f
C897 B.n101 VSUBS 0.00658f
C898 B.n102 VSUBS 0.00658f
C899 B.n103 VSUBS 0.00658f
C900 B.n104 VSUBS 0.00658f
C901 B.n105 VSUBS 0.00658f
C902 B.n106 VSUBS 0.00658f
C903 B.n107 VSUBS 0.00658f
C904 B.n108 VSUBS 0.00658f
C905 B.n109 VSUBS 0.00658f
C906 B.n110 VSUBS 0.00658f
C907 B.n111 VSUBS 0.016605f
C908 B.n112 VSUBS 0.00658f
C909 B.n113 VSUBS 0.00658f
C910 B.n114 VSUBS 0.00658f
C911 B.n115 VSUBS 0.00658f
C912 B.n116 VSUBS 0.00658f
C913 B.n117 VSUBS 0.00658f
C914 B.n118 VSUBS 0.00658f
C915 B.n119 VSUBS 0.00658f
C916 B.n120 VSUBS 0.00658f
C917 B.n121 VSUBS 0.00658f
C918 B.n122 VSUBS 0.00658f
C919 B.n123 VSUBS 0.00658f
C920 B.n124 VSUBS 0.00658f
C921 B.n125 VSUBS 0.00658f
C922 B.n126 VSUBS 0.00658f
C923 B.n127 VSUBS 0.00658f
C924 B.n128 VSUBS 0.00658f
C925 B.n129 VSUBS 0.00658f
C926 B.n130 VSUBS 0.00658f
C927 B.n131 VSUBS 0.00658f
C928 B.n132 VSUBS 0.00658f
C929 B.n133 VSUBS 0.00658f
C930 B.n134 VSUBS 0.00658f
C931 B.n135 VSUBS 0.00658f
C932 B.n136 VSUBS 0.00658f
C933 B.n137 VSUBS 0.00658f
C934 B.n138 VSUBS 0.006193f
C935 B.n139 VSUBS 0.00658f
C936 B.n140 VSUBS 0.00658f
C937 B.n141 VSUBS 0.00658f
C938 B.n142 VSUBS 0.00658f
C939 B.n143 VSUBS 0.00658f
C940 B.t5 VSUBS 0.300459f
C941 B.t4 VSUBS 0.338833f
C942 B.t3 VSUBS 2.36439f
C943 B.n144 VSUBS 0.535724f
C944 B.n145 VSUBS 0.297174f
C945 B.n146 VSUBS 0.00658f
C946 B.n147 VSUBS 0.00658f
C947 B.n148 VSUBS 0.00658f
C948 B.n149 VSUBS 0.00658f
C949 B.n150 VSUBS 0.00658f
C950 B.n151 VSUBS 0.00658f
C951 B.n152 VSUBS 0.00658f
C952 B.n153 VSUBS 0.00658f
C953 B.n154 VSUBS 0.00658f
C954 B.n155 VSUBS 0.00658f
C955 B.n156 VSUBS 0.00658f
C956 B.n157 VSUBS 0.00658f
C957 B.n158 VSUBS 0.00658f
C958 B.n159 VSUBS 0.00658f
C959 B.n160 VSUBS 0.00658f
C960 B.n161 VSUBS 0.00658f
C961 B.n162 VSUBS 0.00658f
C962 B.n163 VSUBS 0.00658f
C963 B.n164 VSUBS 0.00658f
C964 B.n165 VSUBS 0.00658f
C965 B.n166 VSUBS 0.00658f
C966 B.n167 VSUBS 0.00658f
C967 B.n168 VSUBS 0.00658f
C968 B.n169 VSUBS 0.00658f
C969 B.n170 VSUBS 0.00658f
C970 B.n171 VSUBS 0.00658f
C971 B.n172 VSUBS 0.00658f
C972 B.n173 VSUBS 0.016102f
C973 B.n174 VSUBS 0.00658f
C974 B.n175 VSUBS 0.00658f
C975 B.n176 VSUBS 0.00658f
C976 B.n177 VSUBS 0.00658f
C977 B.n178 VSUBS 0.00658f
C978 B.n179 VSUBS 0.00658f
C979 B.n180 VSUBS 0.00658f
C980 B.n181 VSUBS 0.00658f
C981 B.n182 VSUBS 0.00658f
C982 B.n183 VSUBS 0.00658f
C983 B.n184 VSUBS 0.00658f
C984 B.n185 VSUBS 0.00658f
C985 B.n186 VSUBS 0.00658f
C986 B.n187 VSUBS 0.00658f
C987 B.n188 VSUBS 0.00658f
C988 B.n189 VSUBS 0.00658f
C989 B.n190 VSUBS 0.00658f
C990 B.n191 VSUBS 0.00658f
C991 B.n192 VSUBS 0.00658f
C992 B.n193 VSUBS 0.00658f
C993 B.n194 VSUBS 0.00658f
C994 B.n195 VSUBS 0.00658f
C995 B.n196 VSUBS 0.00658f
C996 B.n197 VSUBS 0.00658f
C997 B.n198 VSUBS 0.00658f
C998 B.n199 VSUBS 0.00658f
C999 B.n200 VSUBS 0.00658f
C1000 B.n201 VSUBS 0.00658f
C1001 B.n202 VSUBS 0.00658f
C1002 B.n203 VSUBS 0.00658f
C1003 B.n204 VSUBS 0.00658f
C1004 B.n205 VSUBS 0.00658f
C1005 B.n206 VSUBS 0.00658f
C1006 B.n207 VSUBS 0.00658f
C1007 B.n208 VSUBS 0.00658f
C1008 B.n209 VSUBS 0.00658f
C1009 B.n210 VSUBS 0.00658f
C1010 B.n211 VSUBS 0.00658f
C1011 B.n212 VSUBS 0.00658f
C1012 B.n213 VSUBS 0.00658f
C1013 B.n214 VSUBS 0.00658f
C1014 B.n215 VSUBS 0.00658f
C1015 B.n216 VSUBS 0.00658f
C1016 B.n217 VSUBS 0.00658f
C1017 B.n218 VSUBS 0.00658f
C1018 B.n219 VSUBS 0.00658f
C1019 B.n220 VSUBS 0.00658f
C1020 B.n221 VSUBS 0.00658f
C1021 B.n222 VSUBS 0.00658f
C1022 B.n223 VSUBS 0.00658f
C1023 B.n224 VSUBS 0.00658f
C1024 B.n225 VSUBS 0.00658f
C1025 B.n226 VSUBS 0.00658f
C1026 B.n227 VSUBS 0.00658f
C1027 B.n228 VSUBS 0.016102f
C1028 B.n229 VSUBS 0.016605f
C1029 B.n230 VSUBS 0.016605f
C1030 B.n231 VSUBS 0.00658f
C1031 B.n232 VSUBS 0.00658f
C1032 B.n233 VSUBS 0.00658f
C1033 B.n234 VSUBS 0.00658f
C1034 B.n235 VSUBS 0.00658f
C1035 B.n236 VSUBS 0.00658f
C1036 B.n237 VSUBS 0.00658f
C1037 B.n238 VSUBS 0.00658f
C1038 B.n239 VSUBS 0.00658f
C1039 B.n240 VSUBS 0.00658f
C1040 B.n241 VSUBS 0.00658f
C1041 B.n242 VSUBS 0.00658f
C1042 B.n243 VSUBS 0.00658f
C1043 B.n244 VSUBS 0.00658f
C1044 B.n245 VSUBS 0.00658f
C1045 B.n246 VSUBS 0.00658f
C1046 B.n247 VSUBS 0.00658f
C1047 B.n248 VSUBS 0.00658f
C1048 B.n249 VSUBS 0.00658f
C1049 B.n250 VSUBS 0.00658f
C1050 B.n251 VSUBS 0.00658f
C1051 B.n252 VSUBS 0.00658f
C1052 B.n253 VSUBS 0.00658f
C1053 B.n254 VSUBS 0.00658f
C1054 B.n255 VSUBS 0.00658f
C1055 B.n256 VSUBS 0.00658f
C1056 B.n257 VSUBS 0.00658f
C1057 B.n258 VSUBS 0.00658f
C1058 B.n259 VSUBS 0.00658f
C1059 B.n260 VSUBS 0.00658f
C1060 B.n261 VSUBS 0.00658f
C1061 B.n262 VSUBS 0.00658f
C1062 B.n263 VSUBS 0.00658f
C1063 B.n264 VSUBS 0.00658f
C1064 B.n265 VSUBS 0.00658f
C1065 B.n266 VSUBS 0.00658f
C1066 B.n267 VSUBS 0.00658f
C1067 B.n268 VSUBS 0.00658f
C1068 B.n269 VSUBS 0.00658f
C1069 B.n270 VSUBS 0.00658f
C1070 B.n271 VSUBS 0.00658f
C1071 B.n272 VSUBS 0.00658f
C1072 B.n273 VSUBS 0.00658f
C1073 B.n274 VSUBS 0.00658f
C1074 B.n275 VSUBS 0.00658f
C1075 B.n276 VSUBS 0.00658f
C1076 B.n277 VSUBS 0.00658f
C1077 B.n278 VSUBS 0.00658f
C1078 B.n279 VSUBS 0.00658f
C1079 B.n280 VSUBS 0.00658f
C1080 B.n281 VSUBS 0.00658f
C1081 B.n282 VSUBS 0.00658f
C1082 B.n283 VSUBS 0.00658f
C1083 B.n284 VSUBS 0.00658f
C1084 B.n285 VSUBS 0.00658f
C1085 B.n286 VSUBS 0.00658f
C1086 B.n287 VSUBS 0.00658f
C1087 B.n288 VSUBS 0.00658f
C1088 B.n289 VSUBS 0.00658f
C1089 B.n290 VSUBS 0.00658f
C1090 B.n291 VSUBS 0.00658f
C1091 B.n292 VSUBS 0.00658f
C1092 B.n293 VSUBS 0.00658f
C1093 B.n294 VSUBS 0.00658f
C1094 B.n295 VSUBS 0.00658f
C1095 B.n296 VSUBS 0.00658f
C1096 B.n297 VSUBS 0.00658f
C1097 B.n298 VSUBS 0.00658f
C1098 B.n299 VSUBS 0.00658f
C1099 B.n300 VSUBS 0.00658f
C1100 B.n301 VSUBS 0.00658f
C1101 B.n302 VSUBS 0.00658f
C1102 B.n303 VSUBS 0.00658f
C1103 B.n304 VSUBS 0.00658f
C1104 B.n305 VSUBS 0.00658f
C1105 B.n306 VSUBS 0.00658f
C1106 B.n307 VSUBS 0.00658f
C1107 B.n308 VSUBS 0.00658f
C1108 B.n309 VSUBS 0.00658f
C1109 B.n310 VSUBS 0.00658f
C1110 B.n311 VSUBS 0.006193f
C1111 B.n312 VSUBS 0.015245f
C1112 B.n313 VSUBS 0.003677f
C1113 B.n314 VSUBS 0.00658f
C1114 B.n315 VSUBS 0.00658f
C1115 B.n316 VSUBS 0.00658f
C1116 B.n317 VSUBS 0.00658f
C1117 B.n318 VSUBS 0.00658f
C1118 B.n319 VSUBS 0.00658f
C1119 B.n320 VSUBS 0.00658f
C1120 B.n321 VSUBS 0.00658f
C1121 B.n322 VSUBS 0.00658f
C1122 B.n323 VSUBS 0.00658f
C1123 B.n324 VSUBS 0.00658f
C1124 B.n325 VSUBS 0.00658f
C1125 B.t8 VSUBS 0.300463f
C1126 B.t7 VSUBS 0.338836f
C1127 B.t6 VSUBS 2.36439f
C1128 B.n326 VSUBS 0.535721f
C1129 B.n327 VSUBS 0.297171f
C1130 B.n328 VSUBS 0.015245f
C1131 B.n329 VSUBS 0.003677f
C1132 B.n330 VSUBS 0.00658f
C1133 B.n331 VSUBS 0.00658f
C1134 B.n332 VSUBS 0.00658f
C1135 B.n333 VSUBS 0.00658f
C1136 B.n334 VSUBS 0.00658f
C1137 B.n335 VSUBS 0.00658f
C1138 B.n336 VSUBS 0.00658f
C1139 B.n337 VSUBS 0.00658f
C1140 B.n338 VSUBS 0.00658f
C1141 B.n339 VSUBS 0.00658f
C1142 B.n340 VSUBS 0.00658f
C1143 B.n341 VSUBS 0.00658f
C1144 B.n342 VSUBS 0.00658f
C1145 B.n343 VSUBS 0.00658f
C1146 B.n344 VSUBS 0.00658f
C1147 B.n345 VSUBS 0.00658f
C1148 B.n346 VSUBS 0.00658f
C1149 B.n347 VSUBS 0.00658f
C1150 B.n348 VSUBS 0.00658f
C1151 B.n349 VSUBS 0.00658f
C1152 B.n350 VSUBS 0.00658f
C1153 B.n351 VSUBS 0.00658f
C1154 B.n352 VSUBS 0.00658f
C1155 B.n353 VSUBS 0.00658f
C1156 B.n354 VSUBS 0.00658f
C1157 B.n355 VSUBS 0.00658f
C1158 B.n356 VSUBS 0.00658f
C1159 B.n357 VSUBS 0.00658f
C1160 B.n358 VSUBS 0.00658f
C1161 B.n359 VSUBS 0.00658f
C1162 B.n360 VSUBS 0.00658f
C1163 B.n361 VSUBS 0.00658f
C1164 B.n362 VSUBS 0.00658f
C1165 B.n363 VSUBS 0.00658f
C1166 B.n364 VSUBS 0.00658f
C1167 B.n365 VSUBS 0.00658f
C1168 B.n366 VSUBS 0.00658f
C1169 B.n367 VSUBS 0.00658f
C1170 B.n368 VSUBS 0.00658f
C1171 B.n369 VSUBS 0.00658f
C1172 B.n370 VSUBS 0.00658f
C1173 B.n371 VSUBS 0.00658f
C1174 B.n372 VSUBS 0.00658f
C1175 B.n373 VSUBS 0.00658f
C1176 B.n374 VSUBS 0.00658f
C1177 B.n375 VSUBS 0.00658f
C1178 B.n376 VSUBS 0.00658f
C1179 B.n377 VSUBS 0.00658f
C1180 B.n378 VSUBS 0.00658f
C1181 B.n379 VSUBS 0.00658f
C1182 B.n380 VSUBS 0.00658f
C1183 B.n381 VSUBS 0.00658f
C1184 B.n382 VSUBS 0.00658f
C1185 B.n383 VSUBS 0.00658f
C1186 B.n384 VSUBS 0.00658f
C1187 B.n385 VSUBS 0.00658f
C1188 B.n386 VSUBS 0.00658f
C1189 B.n387 VSUBS 0.00658f
C1190 B.n388 VSUBS 0.00658f
C1191 B.n389 VSUBS 0.00658f
C1192 B.n390 VSUBS 0.00658f
C1193 B.n391 VSUBS 0.00658f
C1194 B.n392 VSUBS 0.00658f
C1195 B.n393 VSUBS 0.00658f
C1196 B.n394 VSUBS 0.00658f
C1197 B.n395 VSUBS 0.00658f
C1198 B.n396 VSUBS 0.00658f
C1199 B.n397 VSUBS 0.00658f
C1200 B.n398 VSUBS 0.00658f
C1201 B.n399 VSUBS 0.00658f
C1202 B.n400 VSUBS 0.00658f
C1203 B.n401 VSUBS 0.00658f
C1204 B.n402 VSUBS 0.00658f
C1205 B.n403 VSUBS 0.00658f
C1206 B.n404 VSUBS 0.00658f
C1207 B.n405 VSUBS 0.00658f
C1208 B.n406 VSUBS 0.00658f
C1209 B.n407 VSUBS 0.00658f
C1210 B.n408 VSUBS 0.00658f
C1211 B.n409 VSUBS 0.00658f
C1212 B.n410 VSUBS 0.00658f
C1213 B.n411 VSUBS 0.00658f
C1214 B.n412 VSUBS 0.015894f
C1215 B.n413 VSUBS 0.016813f
C1216 B.n414 VSUBS 0.016102f
C1217 B.n415 VSUBS 0.00658f
C1218 B.n416 VSUBS 0.00658f
C1219 B.n417 VSUBS 0.00658f
C1220 B.n418 VSUBS 0.00658f
C1221 B.n419 VSUBS 0.00658f
C1222 B.n420 VSUBS 0.00658f
C1223 B.n421 VSUBS 0.00658f
C1224 B.n422 VSUBS 0.00658f
C1225 B.n423 VSUBS 0.00658f
C1226 B.n424 VSUBS 0.00658f
C1227 B.n425 VSUBS 0.00658f
C1228 B.n426 VSUBS 0.00658f
C1229 B.n427 VSUBS 0.00658f
C1230 B.n428 VSUBS 0.00658f
C1231 B.n429 VSUBS 0.00658f
C1232 B.n430 VSUBS 0.00658f
C1233 B.n431 VSUBS 0.00658f
C1234 B.n432 VSUBS 0.00658f
C1235 B.n433 VSUBS 0.00658f
C1236 B.n434 VSUBS 0.00658f
C1237 B.n435 VSUBS 0.00658f
C1238 B.n436 VSUBS 0.00658f
C1239 B.n437 VSUBS 0.00658f
C1240 B.n438 VSUBS 0.00658f
C1241 B.n439 VSUBS 0.00658f
C1242 B.n440 VSUBS 0.00658f
C1243 B.n441 VSUBS 0.00658f
C1244 B.n442 VSUBS 0.00658f
C1245 B.n443 VSUBS 0.00658f
C1246 B.n444 VSUBS 0.00658f
C1247 B.n445 VSUBS 0.00658f
C1248 B.n446 VSUBS 0.00658f
C1249 B.n447 VSUBS 0.00658f
C1250 B.n448 VSUBS 0.00658f
C1251 B.n449 VSUBS 0.00658f
C1252 B.n450 VSUBS 0.00658f
C1253 B.n451 VSUBS 0.00658f
C1254 B.n452 VSUBS 0.00658f
C1255 B.n453 VSUBS 0.00658f
C1256 B.n454 VSUBS 0.00658f
C1257 B.n455 VSUBS 0.00658f
C1258 B.n456 VSUBS 0.00658f
C1259 B.n457 VSUBS 0.00658f
C1260 B.n458 VSUBS 0.00658f
C1261 B.n459 VSUBS 0.00658f
C1262 B.n460 VSUBS 0.00658f
C1263 B.n461 VSUBS 0.00658f
C1264 B.n462 VSUBS 0.00658f
C1265 B.n463 VSUBS 0.00658f
C1266 B.n464 VSUBS 0.00658f
C1267 B.n465 VSUBS 0.00658f
C1268 B.n466 VSUBS 0.00658f
C1269 B.n467 VSUBS 0.00658f
C1270 B.n468 VSUBS 0.00658f
C1271 B.n469 VSUBS 0.00658f
C1272 B.n470 VSUBS 0.00658f
C1273 B.n471 VSUBS 0.00658f
C1274 B.n472 VSUBS 0.00658f
C1275 B.n473 VSUBS 0.00658f
C1276 B.n474 VSUBS 0.00658f
C1277 B.n475 VSUBS 0.00658f
C1278 B.n476 VSUBS 0.00658f
C1279 B.n477 VSUBS 0.00658f
C1280 B.n478 VSUBS 0.00658f
C1281 B.n479 VSUBS 0.00658f
C1282 B.n480 VSUBS 0.00658f
C1283 B.n481 VSUBS 0.00658f
C1284 B.n482 VSUBS 0.00658f
C1285 B.n483 VSUBS 0.00658f
C1286 B.n484 VSUBS 0.00658f
C1287 B.n485 VSUBS 0.00658f
C1288 B.n486 VSUBS 0.00658f
C1289 B.n487 VSUBS 0.00658f
C1290 B.n488 VSUBS 0.00658f
C1291 B.n489 VSUBS 0.00658f
C1292 B.n490 VSUBS 0.00658f
C1293 B.n491 VSUBS 0.00658f
C1294 B.n492 VSUBS 0.00658f
C1295 B.n493 VSUBS 0.00658f
C1296 B.n494 VSUBS 0.00658f
C1297 B.n495 VSUBS 0.00658f
C1298 B.n496 VSUBS 0.00658f
C1299 B.n497 VSUBS 0.00658f
C1300 B.n498 VSUBS 0.00658f
C1301 B.n499 VSUBS 0.00658f
C1302 B.n500 VSUBS 0.00658f
C1303 B.n501 VSUBS 0.00658f
C1304 B.n502 VSUBS 0.016102f
C1305 B.n503 VSUBS 0.016605f
C1306 B.n504 VSUBS 0.016605f
C1307 B.n505 VSUBS 0.00658f
C1308 B.n506 VSUBS 0.00658f
C1309 B.n507 VSUBS 0.00658f
C1310 B.n508 VSUBS 0.00658f
C1311 B.n509 VSUBS 0.00658f
C1312 B.n510 VSUBS 0.00658f
C1313 B.n511 VSUBS 0.00658f
C1314 B.n512 VSUBS 0.00658f
C1315 B.n513 VSUBS 0.00658f
C1316 B.n514 VSUBS 0.00658f
C1317 B.n515 VSUBS 0.00658f
C1318 B.n516 VSUBS 0.00658f
C1319 B.n517 VSUBS 0.00658f
C1320 B.n518 VSUBS 0.00658f
C1321 B.n519 VSUBS 0.00658f
C1322 B.n520 VSUBS 0.00658f
C1323 B.n521 VSUBS 0.00658f
C1324 B.n522 VSUBS 0.00658f
C1325 B.n523 VSUBS 0.00658f
C1326 B.n524 VSUBS 0.00658f
C1327 B.n525 VSUBS 0.00658f
C1328 B.n526 VSUBS 0.00658f
C1329 B.n527 VSUBS 0.00658f
C1330 B.n528 VSUBS 0.00658f
C1331 B.n529 VSUBS 0.00658f
C1332 B.n530 VSUBS 0.00658f
C1333 B.n531 VSUBS 0.00658f
C1334 B.n532 VSUBS 0.00658f
C1335 B.n533 VSUBS 0.00658f
C1336 B.n534 VSUBS 0.00658f
C1337 B.n535 VSUBS 0.00658f
C1338 B.n536 VSUBS 0.00658f
C1339 B.n537 VSUBS 0.00658f
C1340 B.n538 VSUBS 0.00658f
C1341 B.n539 VSUBS 0.00658f
C1342 B.n540 VSUBS 0.00658f
C1343 B.n541 VSUBS 0.00658f
C1344 B.n542 VSUBS 0.00658f
C1345 B.n543 VSUBS 0.00658f
C1346 B.n544 VSUBS 0.00658f
C1347 B.n545 VSUBS 0.00658f
C1348 B.n546 VSUBS 0.00658f
C1349 B.n547 VSUBS 0.00658f
C1350 B.n548 VSUBS 0.00658f
C1351 B.n549 VSUBS 0.00658f
C1352 B.n550 VSUBS 0.00658f
C1353 B.n551 VSUBS 0.00658f
C1354 B.n552 VSUBS 0.00658f
C1355 B.n553 VSUBS 0.00658f
C1356 B.n554 VSUBS 0.00658f
C1357 B.n555 VSUBS 0.00658f
C1358 B.n556 VSUBS 0.00658f
C1359 B.n557 VSUBS 0.00658f
C1360 B.n558 VSUBS 0.00658f
C1361 B.n559 VSUBS 0.00658f
C1362 B.n560 VSUBS 0.00658f
C1363 B.n561 VSUBS 0.00658f
C1364 B.n562 VSUBS 0.00658f
C1365 B.n563 VSUBS 0.00658f
C1366 B.n564 VSUBS 0.00658f
C1367 B.n565 VSUBS 0.00658f
C1368 B.n566 VSUBS 0.00658f
C1369 B.n567 VSUBS 0.00658f
C1370 B.n568 VSUBS 0.00658f
C1371 B.n569 VSUBS 0.00658f
C1372 B.n570 VSUBS 0.00658f
C1373 B.n571 VSUBS 0.00658f
C1374 B.n572 VSUBS 0.00658f
C1375 B.n573 VSUBS 0.00658f
C1376 B.n574 VSUBS 0.00658f
C1377 B.n575 VSUBS 0.00658f
C1378 B.n576 VSUBS 0.00658f
C1379 B.n577 VSUBS 0.00658f
C1380 B.n578 VSUBS 0.00658f
C1381 B.n579 VSUBS 0.00658f
C1382 B.n580 VSUBS 0.00658f
C1383 B.n581 VSUBS 0.00658f
C1384 B.n582 VSUBS 0.00658f
C1385 B.n583 VSUBS 0.00658f
C1386 B.n584 VSUBS 0.00658f
C1387 B.n585 VSUBS 0.006193f
C1388 B.n586 VSUBS 0.015245f
C1389 B.n587 VSUBS 0.003677f
C1390 B.n588 VSUBS 0.00658f
C1391 B.n589 VSUBS 0.00658f
C1392 B.n590 VSUBS 0.00658f
C1393 B.n591 VSUBS 0.00658f
C1394 B.n592 VSUBS 0.00658f
C1395 B.n593 VSUBS 0.00658f
C1396 B.n594 VSUBS 0.00658f
C1397 B.n595 VSUBS 0.00658f
C1398 B.n596 VSUBS 0.00658f
C1399 B.n597 VSUBS 0.00658f
C1400 B.n598 VSUBS 0.00658f
C1401 B.n599 VSUBS 0.00658f
C1402 B.n600 VSUBS 0.003677f
C1403 B.n601 VSUBS 0.00658f
C1404 B.n602 VSUBS 0.00658f
C1405 B.n603 VSUBS 0.006193f
C1406 B.n604 VSUBS 0.00658f
C1407 B.n605 VSUBS 0.00658f
C1408 B.n606 VSUBS 0.00658f
C1409 B.n607 VSUBS 0.00658f
C1410 B.n608 VSUBS 0.00658f
C1411 B.n609 VSUBS 0.00658f
C1412 B.n610 VSUBS 0.00658f
C1413 B.n611 VSUBS 0.00658f
C1414 B.n612 VSUBS 0.00658f
C1415 B.n613 VSUBS 0.00658f
C1416 B.n614 VSUBS 0.00658f
C1417 B.n615 VSUBS 0.00658f
C1418 B.n616 VSUBS 0.00658f
C1419 B.n617 VSUBS 0.00658f
C1420 B.n618 VSUBS 0.00658f
C1421 B.n619 VSUBS 0.00658f
C1422 B.n620 VSUBS 0.00658f
C1423 B.n621 VSUBS 0.00658f
C1424 B.n622 VSUBS 0.00658f
C1425 B.n623 VSUBS 0.00658f
C1426 B.n624 VSUBS 0.00658f
C1427 B.n625 VSUBS 0.00658f
C1428 B.n626 VSUBS 0.00658f
C1429 B.n627 VSUBS 0.00658f
C1430 B.n628 VSUBS 0.00658f
C1431 B.n629 VSUBS 0.00658f
C1432 B.n630 VSUBS 0.00658f
C1433 B.n631 VSUBS 0.00658f
C1434 B.n632 VSUBS 0.00658f
C1435 B.n633 VSUBS 0.00658f
C1436 B.n634 VSUBS 0.00658f
C1437 B.n635 VSUBS 0.00658f
C1438 B.n636 VSUBS 0.00658f
C1439 B.n637 VSUBS 0.00658f
C1440 B.n638 VSUBS 0.00658f
C1441 B.n639 VSUBS 0.00658f
C1442 B.n640 VSUBS 0.00658f
C1443 B.n641 VSUBS 0.00658f
C1444 B.n642 VSUBS 0.00658f
C1445 B.n643 VSUBS 0.00658f
C1446 B.n644 VSUBS 0.00658f
C1447 B.n645 VSUBS 0.00658f
C1448 B.n646 VSUBS 0.00658f
C1449 B.n647 VSUBS 0.00658f
C1450 B.n648 VSUBS 0.00658f
C1451 B.n649 VSUBS 0.00658f
C1452 B.n650 VSUBS 0.00658f
C1453 B.n651 VSUBS 0.00658f
C1454 B.n652 VSUBS 0.00658f
C1455 B.n653 VSUBS 0.00658f
C1456 B.n654 VSUBS 0.00658f
C1457 B.n655 VSUBS 0.00658f
C1458 B.n656 VSUBS 0.00658f
C1459 B.n657 VSUBS 0.00658f
C1460 B.n658 VSUBS 0.00658f
C1461 B.n659 VSUBS 0.00658f
C1462 B.n660 VSUBS 0.00658f
C1463 B.n661 VSUBS 0.00658f
C1464 B.n662 VSUBS 0.00658f
C1465 B.n663 VSUBS 0.00658f
C1466 B.n664 VSUBS 0.00658f
C1467 B.n665 VSUBS 0.00658f
C1468 B.n666 VSUBS 0.00658f
C1469 B.n667 VSUBS 0.00658f
C1470 B.n668 VSUBS 0.00658f
C1471 B.n669 VSUBS 0.00658f
C1472 B.n670 VSUBS 0.00658f
C1473 B.n671 VSUBS 0.00658f
C1474 B.n672 VSUBS 0.00658f
C1475 B.n673 VSUBS 0.00658f
C1476 B.n674 VSUBS 0.00658f
C1477 B.n675 VSUBS 0.00658f
C1478 B.n676 VSUBS 0.00658f
C1479 B.n677 VSUBS 0.00658f
C1480 B.n678 VSUBS 0.00658f
C1481 B.n679 VSUBS 0.00658f
C1482 B.n680 VSUBS 0.00658f
C1483 B.n681 VSUBS 0.00658f
C1484 B.n682 VSUBS 0.00658f
C1485 B.n683 VSUBS 0.016605f
C1486 B.n684 VSUBS 0.016605f
C1487 B.n685 VSUBS 0.016102f
C1488 B.n686 VSUBS 0.00658f
C1489 B.n687 VSUBS 0.00658f
C1490 B.n688 VSUBS 0.00658f
C1491 B.n689 VSUBS 0.00658f
C1492 B.n690 VSUBS 0.00658f
C1493 B.n691 VSUBS 0.00658f
C1494 B.n692 VSUBS 0.00658f
C1495 B.n693 VSUBS 0.00658f
C1496 B.n694 VSUBS 0.00658f
C1497 B.n695 VSUBS 0.00658f
C1498 B.n696 VSUBS 0.00658f
C1499 B.n697 VSUBS 0.00658f
C1500 B.n698 VSUBS 0.00658f
C1501 B.n699 VSUBS 0.00658f
C1502 B.n700 VSUBS 0.00658f
C1503 B.n701 VSUBS 0.00658f
C1504 B.n702 VSUBS 0.00658f
C1505 B.n703 VSUBS 0.00658f
C1506 B.n704 VSUBS 0.00658f
C1507 B.n705 VSUBS 0.00658f
C1508 B.n706 VSUBS 0.00658f
C1509 B.n707 VSUBS 0.00658f
C1510 B.n708 VSUBS 0.00658f
C1511 B.n709 VSUBS 0.00658f
C1512 B.n710 VSUBS 0.00658f
C1513 B.n711 VSUBS 0.00658f
C1514 B.n712 VSUBS 0.00658f
C1515 B.n713 VSUBS 0.00658f
C1516 B.n714 VSUBS 0.00658f
C1517 B.n715 VSUBS 0.00658f
C1518 B.n716 VSUBS 0.00658f
C1519 B.n717 VSUBS 0.00658f
C1520 B.n718 VSUBS 0.00658f
C1521 B.n719 VSUBS 0.00658f
C1522 B.n720 VSUBS 0.00658f
C1523 B.n721 VSUBS 0.00658f
C1524 B.n722 VSUBS 0.00658f
C1525 B.n723 VSUBS 0.00658f
C1526 B.n724 VSUBS 0.00658f
C1527 B.n725 VSUBS 0.00658f
C1528 B.n726 VSUBS 0.00658f
C1529 B.n727 VSUBS 0.008587f
C1530 B.n728 VSUBS 0.009147f
C1531 B.n729 VSUBS 0.01819f
.ends

