* NGSPICE file created from diff_pair_sample_0807.ext - technology: sky130A

.subckt diff_pair_sample_0807 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.11
X1 VTAIL.t13 VP.t1 VDD1.t8 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X2 VDD2.t9 VN.t0 VTAIL.t17 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.11
X3 B.t11 B.t9 B.t10 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.11
X4 VDD2.t8 VN.t1 VTAIL.t14 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X5 VTAIL.t3 VN.t2 VDD2.t7 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X6 B.t8 B.t6 B.t7 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.11
X7 VDD2.t6 VN.t3 VTAIL.t16 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.11
X8 VTAIL.t19 VN.t4 VDD2.t5 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X9 VDD1.t7 VP.t2 VTAIL.t8 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.11
X10 VDD2.t4 VN.t5 VTAIL.t18 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.11
X11 VDD1.t6 VP.t3 VTAIL.t7 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.11
X12 VTAIL.t4 VP.t4 VDD1.t5 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X13 B.t5 B.t3 B.t4 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.11
X14 VDD2.t3 VN.t6 VTAIL.t15 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X15 VTAIL.t5 VP.t5 VDD1.t4 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X16 VDD1.t3 VP.t6 VTAIL.t6 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X17 VTAIL.t2 VN.t7 VDD2.t2 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X18 VTAIL.t0 VN.t8 VDD2.t1 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X19 VDD1.t2 VP.t7 VTAIL.t12 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.11
X20 VDD2.t0 VN.t9 VTAIL.t1 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.11
X21 VDD1.t1 VP.t8 VTAIL.t11 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
X22 B.t2 B.t0 B.t1 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.11
X23 VTAIL.t9 VP.t9 VDD1.t0 w_n5098_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.11
R0 VP.n26 VP.t2 183.764
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n25 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n24 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n23 161.3
R7 VP.n38 VP.n37 161.3
R8 VP.n39 VP.n22 161.3
R9 VP.n41 VP.n40 161.3
R10 VP.n42 VP.n21 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n45 VP.n20 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n49 VP.n48 161.3
R15 VP.n50 VP.n18 161.3
R16 VP.n52 VP.n51 161.3
R17 VP.n53 VP.n17 161.3
R18 VP.n55 VP.n54 161.3
R19 VP.n56 VP.n16 161.3
R20 VP.n58 VP.n57 161.3
R21 VP.n103 VP.n102 161.3
R22 VP.n101 VP.n1 161.3
R23 VP.n100 VP.n99 161.3
R24 VP.n98 VP.n2 161.3
R25 VP.n97 VP.n96 161.3
R26 VP.n95 VP.n3 161.3
R27 VP.n94 VP.n93 161.3
R28 VP.n92 VP.n91 161.3
R29 VP.n90 VP.n5 161.3
R30 VP.n89 VP.n88 161.3
R31 VP.n87 VP.n6 161.3
R32 VP.n86 VP.n85 161.3
R33 VP.n84 VP.n7 161.3
R34 VP.n83 VP.n82 161.3
R35 VP.n81 VP.n8 161.3
R36 VP.n80 VP.n79 161.3
R37 VP.n78 VP.n9 161.3
R38 VP.n77 VP.n76 161.3
R39 VP.n75 VP.n10 161.3
R40 VP.n74 VP.n73 161.3
R41 VP.n71 VP.n11 161.3
R42 VP.n70 VP.n69 161.3
R43 VP.n68 VP.n12 161.3
R44 VP.n67 VP.n66 161.3
R45 VP.n65 VP.n13 161.3
R46 VP.n64 VP.n63 161.3
R47 VP.n62 VP.n14 161.3
R48 VP.n83 VP.t8 150.412
R49 VP.n60 VP.t7 150.412
R50 VP.n72 VP.t9 150.412
R51 VP.n4 VP.t5 150.412
R52 VP.n0 VP.t3 150.412
R53 VP.n38 VP.t6 150.412
R54 VP.n15 VP.t0 150.412
R55 VP.n19 VP.t4 150.412
R56 VP.n27 VP.t1 150.412
R57 VP.n61 VP.n60 71.4725
R58 VP.n104 VP.n0 71.4725
R59 VP.n59 VP.n15 71.4725
R60 VP.n61 VP.n59 61.6281
R61 VP.n78 VP.n77 56.5193
R62 VP.n89 VP.n6 56.5193
R63 VP.n44 VP.n21 56.5193
R64 VP.n33 VP.n32 56.5193
R65 VP.n66 VP.n65 56.0336
R66 VP.n100 VP.n2 56.0336
R67 VP.n55 VP.n17 56.0336
R68 VP.n27 VP.n26 52.2938
R69 VP.n66 VP.n12 24.9531
R70 VP.n96 VP.n2 24.9531
R71 VP.n51 VP.n17 24.9531
R72 VP.n64 VP.n14 24.4675
R73 VP.n65 VP.n64 24.4675
R74 VP.n70 VP.n12 24.4675
R75 VP.n71 VP.n70 24.4675
R76 VP.n73 VP.n10 24.4675
R77 VP.n77 VP.n10 24.4675
R78 VP.n79 VP.n78 24.4675
R79 VP.n79 VP.n8 24.4675
R80 VP.n83 VP.n8 24.4675
R81 VP.n84 VP.n83 24.4675
R82 VP.n85 VP.n84 24.4675
R83 VP.n85 VP.n6 24.4675
R84 VP.n90 VP.n89 24.4675
R85 VP.n91 VP.n90 24.4675
R86 VP.n95 VP.n94 24.4675
R87 VP.n96 VP.n95 24.4675
R88 VP.n101 VP.n100 24.4675
R89 VP.n102 VP.n101 24.4675
R90 VP.n56 VP.n55 24.4675
R91 VP.n57 VP.n56 24.4675
R92 VP.n45 VP.n44 24.4675
R93 VP.n46 VP.n45 24.4675
R94 VP.n50 VP.n49 24.4675
R95 VP.n51 VP.n50 24.4675
R96 VP.n34 VP.n33 24.4675
R97 VP.n34 VP.n23 24.4675
R98 VP.n38 VP.n23 24.4675
R99 VP.n39 VP.n38 24.4675
R100 VP.n40 VP.n39 24.4675
R101 VP.n40 VP.n21 24.4675
R102 VP.n28 VP.n25 24.4675
R103 VP.n32 VP.n25 24.4675
R104 VP.n73 VP.n72 21.5315
R105 VP.n91 VP.n4 21.5315
R106 VP.n46 VP.n19 21.5315
R107 VP.n28 VP.n27 21.5315
R108 VP.n60 VP.n14 18.5954
R109 VP.n102 VP.n0 18.5954
R110 VP.n57 VP.n15 18.5954
R111 VP.n29 VP.n26 3.98136
R112 VP.n72 VP.n71 2.93654
R113 VP.n94 VP.n4 2.93654
R114 VP.n49 VP.n19 2.93654
R115 VP.n59 VP.n58 0.354971
R116 VP.n62 VP.n61 0.354971
R117 VP.n104 VP.n103 0.354971
R118 VP VP.n104 0.26696
R119 VP.n30 VP.n29 0.189894
R120 VP.n31 VP.n30 0.189894
R121 VP.n31 VP.n24 0.189894
R122 VP.n35 VP.n24 0.189894
R123 VP.n36 VP.n35 0.189894
R124 VP.n37 VP.n36 0.189894
R125 VP.n37 VP.n22 0.189894
R126 VP.n41 VP.n22 0.189894
R127 VP.n42 VP.n41 0.189894
R128 VP.n43 VP.n42 0.189894
R129 VP.n43 VP.n20 0.189894
R130 VP.n47 VP.n20 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n18 0.189894
R133 VP.n52 VP.n18 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n16 0.189894
R137 VP.n58 VP.n16 0.189894
R138 VP.n63 VP.n62 0.189894
R139 VP.n63 VP.n13 0.189894
R140 VP.n67 VP.n13 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n69 VP.n68 0.189894
R143 VP.n69 VP.n11 0.189894
R144 VP.n74 VP.n11 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n76 VP.n75 0.189894
R147 VP.n76 VP.n9 0.189894
R148 VP.n80 VP.n9 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n82 VP.n81 0.189894
R151 VP.n82 VP.n7 0.189894
R152 VP.n86 VP.n7 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n88 VP.n87 0.189894
R155 VP.n88 VP.n5 0.189894
R156 VP.n92 VP.n5 0.189894
R157 VP.n93 VP.n92 0.189894
R158 VP.n93 VP.n3 0.189894
R159 VP.n97 VP.n3 0.189894
R160 VP.n98 VP.n97 0.189894
R161 VP.n99 VP.n98 0.189894
R162 VP.n99 VP.n1 0.189894
R163 VP.n103 VP.n1 0.189894
R164 VTAIL.n367 VTAIL.n366 585
R165 VTAIL.n364 VTAIL.n363 585
R166 VTAIL.n373 VTAIL.n372 585
R167 VTAIL.n375 VTAIL.n374 585
R168 VTAIL.n360 VTAIL.n359 585
R169 VTAIL.n381 VTAIL.n380 585
R170 VTAIL.n384 VTAIL.n383 585
R171 VTAIL.n382 VTAIL.n356 585
R172 VTAIL.n389 VTAIL.n355 585
R173 VTAIL.n391 VTAIL.n390 585
R174 VTAIL.n393 VTAIL.n392 585
R175 VTAIL.n352 VTAIL.n351 585
R176 VTAIL.n399 VTAIL.n398 585
R177 VTAIL.n401 VTAIL.n400 585
R178 VTAIL.n348 VTAIL.n347 585
R179 VTAIL.n407 VTAIL.n406 585
R180 VTAIL.n409 VTAIL.n408 585
R181 VTAIL.n344 VTAIL.n343 585
R182 VTAIL.n415 VTAIL.n414 585
R183 VTAIL.n417 VTAIL.n416 585
R184 VTAIL.n340 VTAIL.n339 585
R185 VTAIL.n423 VTAIL.n422 585
R186 VTAIL.n425 VTAIL.n424 585
R187 VTAIL.n336 VTAIL.n335 585
R188 VTAIL.n431 VTAIL.n430 585
R189 VTAIL.n433 VTAIL.n432 585
R190 VTAIL.n37 VTAIL.n36 585
R191 VTAIL.n34 VTAIL.n33 585
R192 VTAIL.n43 VTAIL.n42 585
R193 VTAIL.n45 VTAIL.n44 585
R194 VTAIL.n30 VTAIL.n29 585
R195 VTAIL.n51 VTAIL.n50 585
R196 VTAIL.n54 VTAIL.n53 585
R197 VTAIL.n52 VTAIL.n26 585
R198 VTAIL.n59 VTAIL.n25 585
R199 VTAIL.n61 VTAIL.n60 585
R200 VTAIL.n63 VTAIL.n62 585
R201 VTAIL.n22 VTAIL.n21 585
R202 VTAIL.n69 VTAIL.n68 585
R203 VTAIL.n71 VTAIL.n70 585
R204 VTAIL.n18 VTAIL.n17 585
R205 VTAIL.n77 VTAIL.n76 585
R206 VTAIL.n79 VTAIL.n78 585
R207 VTAIL.n14 VTAIL.n13 585
R208 VTAIL.n85 VTAIL.n84 585
R209 VTAIL.n87 VTAIL.n86 585
R210 VTAIL.n10 VTAIL.n9 585
R211 VTAIL.n93 VTAIL.n92 585
R212 VTAIL.n95 VTAIL.n94 585
R213 VTAIL.n6 VTAIL.n5 585
R214 VTAIL.n101 VTAIL.n100 585
R215 VTAIL.n103 VTAIL.n102 585
R216 VTAIL.n327 VTAIL.n326 585
R217 VTAIL.n325 VTAIL.n324 585
R218 VTAIL.n230 VTAIL.n229 585
R219 VTAIL.n319 VTAIL.n318 585
R220 VTAIL.n317 VTAIL.n316 585
R221 VTAIL.n234 VTAIL.n233 585
R222 VTAIL.n311 VTAIL.n310 585
R223 VTAIL.n309 VTAIL.n308 585
R224 VTAIL.n238 VTAIL.n237 585
R225 VTAIL.n303 VTAIL.n302 585
R226 VTAIL.n301 VTAIL.n300 585
R227 VTAIL.n242 VTAIL.n241 585
R228 VTAIL.n295 VTAIL.n294 585
R229 VTAIL.n293 VTAIL.n292 585
R230 VTAIL.n246 VTAIL.n245 585
R231 VTAIL.n287 VTAIL.n286 585
R232 VTAIL.n285 VTAIL.n284 585
R233 VTAIL.n283 VTAIL.n249 585
R234 VTAIL.n253 VTAIL.n250 585
R235 VTAIL.n278 VTAIL.n277 585
R236 VTAIL.n276 VTAIL.n275 585
R237 VTAIL.n255 VTAIL.n254 585
R238 VTAIL.n270 VTAIL.n269 585
R239 VTAIL.n268 VTAIL.n267 585
R240 VTAIL.n259 VTAIL.n258 585
R241 VTAIL.n262 VTAIL.n261 585
R242 VTAIL.n217 VTAIL.n216 585
R243 VTAIL.n215 VTAIL.n214 585
R244 VTAIL.n120 VTAIL.n119 585
R245 VTAIL.n209 VTAIL.n208 585
R246 VTAIL.n207 VTAIL.n206 585
R247 VTAIL.n124 VTAIL.n123 585
R248 VTAIL.n201 VTAIL.n200 585
R249 VTAIL.n199 VTAIL.n198 585
R250 VTAIL.n128 VTAIL.n127 585
R251 VTAIL.n193 VTAIL.n192 585
R252 VTAIL.n191 VTAIL.n190 585
R253 VTAIL.n132 VTAIL.n131 585
R254 VTAIL.n185 VTAIL.n184 585
R255 VTAIL.n183 VTAIL.n182 585
R256 VTAIL.n136 VTAIL.n135 585
R257 VTAIL.n177 VTAIL.n176 585
R258 VTAIL.n175 VTAIL.n174 585
R259 VTAIL.n173 VTAIL.n139 585
R260 VTAIL.n143 VTAIL.n140 585
R261 VTAIL.n168 VTAIL.n167 585
R262 VTAIL.n166 VTAIL.n165 585
R263 VTAIL.n145 VTAIL.n144 585
R264 VTAIL.n160 VTAIL.n159 585
R265 VTAIL.n158 VTAIL.n157 585
R266 VTAIL.n149 VTAIL.n148 585
R267 VTAIL.n152 VTAIL.n151 585
R268 VTAIL.n432 VTAIL.n332 498.474
R269 VTAIL.n102 VTAIL.n2 498.474
R270 VTAIL.n326 VTAIL.n226 498.474
R271 VTAIL.n216 VTAIL.n116 498.474
R272 VTAIL.t1 VTAIL.n365 329.036
R273 VTAIL.t7 VTAIL.n35 329.036
R274 VTAIL.t10 VTAIL.n260 329.036
R275 VTAIL.t18 VTAIL.n150 329.036
R276 VTAIL.n366 VTAIL.n363 171.744
R277 VTAIL.n373 VTAIL.n363 171.744
R278 VTAIL.n374 VTAIL.n373 171.744
R279 VTAIL.n374 VTAIL.n359 171.744
R280 VTAIL.n381 VTAIL.n359 171.744
R281 VTAIL.n383 VTAIL.n381 171.744
R282 VTAIL.n383 VTAIL.n382 171.744
R283 VTAIL.n382 VTAIL.n355 171.744
R284 VTAIL.n391 VTAIL.n355 171.744
R285 VTAIL.n392 VTAIL.n391 171.744
R286 VTAIL.n392 VTAIL.n351 171.744
R287 VTAIL.n399 VTAIL.n351 171.744
R288 VTAIL.n400 VTAIL.n399 171.744
R289 VTAIL.n400 VTAIL.n347 171.744
R290 VTAIL.n407 VTAIL.n347 171.744
R291 VTAIL.n408 VTAIL.n407 171.744
R292 VTAIL.n408 VTAIL.n343 171.744
R293 VTAIL.n415 VTAIL.n343 171.744
R294 VTAIL.n416 VTAIL.n415 171.744
R295 VTAIL.n416 VTAIL.n339 171.744
R296 VTAIL.n423 VTAIL.n339 171.744
R297 VTAIL.n424 VTAIL.n423 171.744
R298 VTAIL.n424 VTAIL.n335 171.744
R299 VTAIL.n431 VTAIL.n335 171.744
R300 VTAIL.n432 VTAIL.n431 171.744
R301 VTAIL.n36 VTAIL.n33 171.744
R302 VTAIL.n43 VTAIL.n33 171.744
R303 VTAIL.n44 VTAIL.n43 171.744
R304 VTAIL.n44 VTAIL.n29 171.744
R305 VTAIL.n51 VTAIL.n29 171.744
R306 VTAIL.n53 VTAIL.n51 171.744
R307 VTAIL.n53 VTAIL.n52 171.744
R308 VTAIL.n52 VTAIL.n25 171.744
R309 VTAIL.n61 VTAIL.n25 171.744
R310 VTAIL.n62 VTAIL.n61 171.744
R311 VTAIL.n62 VTAIL.n21 171.744
R312 VTAIL.n69 VTAIL.n21 171.744
R313 VTAIL.n70 VTAIL.n69 171.744
R314 VTAIL.n70 VTAIL.n17 171.744
R315 VTAIL.n77 VTAIL.n17 171.744
R316 VTAIL.n78 VTAIL.n77 171.744
R317 VTAIL.n78 VTAIL.n13 171.744
R318 VTAIL.n85 VTAIL.n13 171.744
R319 VTAIL.n86 VTAIL.n85 171.744
R320 VTAIL.n86 VTAIL.n9 171.744
R321 VTAIL.n93 VTAIL.n9 171.744
R322 VTAIL.n94 VTAIL.n93 171.744
R323 VTAIL.n94 VTAIL.n5 171.744
R324 VTAIL.n101 VTAIL.n5 171.744
R325 VTAIL.n102 VTAIL.n101 171.744
R326 VTAIL.n326 VTAIL.n325 171.744
R327 VTAIL.n325 VTAIL.n229 171.744
R328 VTAIL.n318 VTAIL.n229 171.744
R329 VTAIL.n318 VTAIL.n317 171.744
R330 VTAIL.n317 VTAIL.n233 171.744
R331 VTAIL.n310 VTAIL.n233 171.744
R332 VTAIL.n310 VTAIL.n309 171.744
R333 VTAIL.n309 VTAIL.n237 171.744
R334 VTAIL.n302 VTAIL.n237 171.744
R335 VTAIL.n302 VTAIL.n301 171.744
R336 VTAIL.n301 VTAIL.n241 171.744
R337 VTAIL.n294 VTAIL.n241 171.744
R338 VTAIL.n294 VTAIL.n293 171.744
R339 VTAIL.n293 VTAIL.n245 171.744
R340 VTAIL.n286 VTAIL.n245 171.744
R341 VTAIL.n286 VTAIL.n285 171.744
R342 VTAIL.n285 VTAIL.n249 171.744
R343 VTAIL.n253 VTAIL.n249 171.744
R344 VTAIL.n277 VTAIL.n253 171.744
R345 VTAIL.n277 VTAIL.n276 171.744
R346 VTAIL.n276 VTAIL.n254 171.744
R347 VTAIL.n269 VTAIL.n254 171.744
R348 VTAIL.n269 VTAIL.n268 171.744
R349 VTAIL.n268 VTAIL.n258 171.744
R350 VTAIL.n261 VTAIL.n258 171.744
R351 VTAIL.n216 VTAIL.n215 171.744
R352 VTAIL.n215 VTAIL.n119 171.744
R353 VTAIL.n208 VTAIL.n119 171.744
R354 VTAIL.n208 VTAIL.n207 171.744
R355 VTAIL.n207 VTAIL.n123 171.744
R356 VTAIL.n200 VTAIL.n123 171.744
R357 VTAIL.n200 VTAIL.n199 171.744
R358 VTAIL.n199 VTAIL.n127 171.744
R359 VTAIL.n192 VTAIL.n127 171.744
R360 VTAIL.n192 VTAIL.n191 171.744
R361 VTAIL.n191 VTAIL.n131 171.744
R362 VTAIL.n184 VTAIL.n131 171.744
R363 VTAIL.n184 VTAIL.n183 171.744
R364 VTAIL.n183 VTAIL.n135 171.744
R365 VTAIL.n176 VTAIL.n135 171.744
R366 VTAIL.n176 VTAIL.n175 171.744
R367 VTAIL.n175 VTAIL.n139 171.744
R368 VTAIL.n143 VTAIL.n139 171.744
R369 VTAIL.n167 VTAIL.n143 171.744
R370 VTAIL.n167 VTAIL.n166 171.744
R371 VTAIL.n166 VTAIL.n144 171.744
R372 VTAIL.n159 VTAIL.n144 171.744
R373 VTAIL.n159 VTAIL.n158 171.744
R374 VTAIL.n158 VTAIL.n148 171.744
R375 VTAIL.n151 VTAIL.n148 171.744
R376 VTAIL.n366 VTAIL.t1 85.8723
R377 VTAIL.n36 VTAIL.t7 85.8723
R378 VTAIL.n261 VTAIL.t10 85.8723
R379 VTAIL.n151 VTAIL.t18 85.8723
R380 VTAIL.n225 VTAIL.n224 52.9099
R381 VTAIL.n223 VTAIL.n222 52.9099
R382 VTAIL.n115 VTAIL.n114 52.9099
R383 VTAIL.n113 VTAIL.n112 52.9099
R384 VTAIL.n439 VTAIL.n438 52.9097
R385 VTAIL.n1 VTAIL.n0 52.9097
R386 VTAIL.n109 VTAIL.n108 52.9097
R387 VTAIL.n111 VTAIL.n110 52.9097
R388 VTAIL.n113 VTAIL.n111 35.0307
R389 VTAIL.n437 VTAIL.n436 33.9308
R390 VTAIL.n107 VTAIL.n106 33.9308
R391 VTAIL.n331 VTAIL.n330 33.9308
R392 VTAIL.n221 VTAIL.n220 33.9308
R393 VTAIL.n437 VTAIL.n331 32.0652
R394 VTAIL.n390 VTAIL.n389 13.1884
R395 VTAIL.n60 VTAIL.n59 13.1884
R396 VTAIL.n284 VTAIL.n283 13.1884
R397 VTAIL.n174 VTAIL.n173 13.1884
R398 VTAIL.n388 VTAIL.n356 12.8005
R399 VTAIL.n393 VTAIL.n354 12.8005
R400 VTAIL.n434 VTAIL.n433 12.8005
R401 VTAIL.n58 VTAIL.n26 12.8005
R402 VTAIL.n63 VTAIL.n24 12.8005
R403 VTAIL.n104 VTAIL.n103 12.8005
R404 VTAIL.n328 VTAIL.n327 12.8005
R405 VTAIL.n287 VTAIL.n248 12.8005
R406 VTAIL.n282 VTAIL.n250 12.8005
R407 VTAIL.n218 VTAIL.n217 12.8005
R408 VTAIL.n177 VTAIL.n138 12.8005
R409 VTAIL.n172 VTAIL.n140 12.8005
R410 VTAIL.n385 VTAIL.n384 12.0247
R411 VTAIL.n394 VTAIL.n352 12.0247
R412 VTAIL.n430 VTAIL.n334 12.0247
R413 VTAIL.n55 VTAIL.n54 12.0247
R414 VTAIL.n64 VTAIL.n22 12.0247
R415 VTAIL.n100 VTAIL.n4 12.0247
R416 VTAIL.n324 VTAIL.n228 12.0247
R417 VTAIL.n288 VTAIL.n246 12.0247
R418 VTAIL.n279 VTAIL.n278 12.0247
R419 VTAIL.n214 VTAIL.n118 12.0247
R420 VTAIL.n178 VTAIL.n136 12.0247
R421 VTAIL.n169 VTAIL.n168 12.0247
R422 VTAIL.n380 VTAIL.n358 11.249
R423 VTAIL.n398 VTAIL.n397 11.249
R424 VTAIL.n429 VTAIL.n336 11.249
R425 VTAIL.n50 VTAIL.n28 11.249
R426 VTAIL.n68 VTAIL.n67 11.249
R427 VTAIL.n99 VTAIL.n6 11.249
R428 VTAIL.n323 VTAIL.n230 11.249
R429 VTAIL.n292 VTAIL.n291 11.249
R430 VTAIL.n275 VTAIL.n252 11.249
R431 VTAIL.n213 VTAIL.n120 11.249
R432 VTAIL.n182 VTAIL.n181 11.249
R433 VTAIL.n165 VTAIL.n142 11.249
R434 VTAIL.n367 VTAIL.n365 10.7239
R435 VTAIL.n37 VTAIL.n35 10.7239
R436 VTAIL.n262 VTAIL.n260 10.7239
R437 VTAIL.n152 VTAIL.n150 10.7239
R438 VTAIL.n379 VTAIL.n360 10.4732
R439 VTAIL.n401 VTAIL.n350 10.4732
R440 VTAIL.n426 VTAIL.n425 10.4732
R441 VTAIL.n49 VTAIL.n30 10.4732
R442 VTAIL.n71 VTAIL.n20 10.4732
R443 VTAIL.n96 VTAIL.n95 10.4732
R444 VTAIL.n320 VTAIL.n319 10.4732
R445 VTAIL.n295 VTAIL.n244 10.4732
R446 VTAIL.n274 VTAIL.n255 10.4732
R447 VTAIL.n210 VTAIL.n209 10.4732
R448 VTAIL.n185 VTAIL.n134 10.4732
R449 VTAIL.n164 VTAIL.n145 10.4732
R450 VTAIL.n376 VTAIL.n375 9.69747
R451 VTAIL.n402 VTAIL.n348 9.69747
R452 VTAIL.n422 VTAIL.n338 9.69747
R453 VTAIL.n46 VTAIL.n45 9.69747
R454 VTAIL.n72 VTAIL.n18 9.69747
R455 VTAIL.n92 VTAIL.n8 9.69747
R456 VTAIL.n316 VTAIL.n232 9.69747
R457 VTAIL.n296 VTAIL.n242 9.69747
R458 VTAIL.n271 VTAIL.n270 9.69747
R459 VTAIL.n206 VTAIL.n122 9.69747
R460 VTAIL.n186 VTAIL.n132 9.69747
R461 VTAIL.n161 VTAIL.n160 9.69747
R462 VTAIL.n436 VTAIL.n435 9.45567
R463 VTAIL.n106 VTAIL.n105 9.45567
R464 VTAIL.n330 VTAIL.n329 9.45567
R465 VTAIL.n220 VTAIL.n219 9.45567
R466 VTAIL.n411 VTAIL.n410 9.3005
R467 VTAIL.n346 VTAIL.n345 9.3005
R468 VTAIL.n405 VTAIL.n404 9.3005
R469 VTAIL.n403 VTAIL.n402 9.3005
R470 VTAIL.n350 VTAIL.n349 9.3005
R471 VTAIL.n397 VTAIL.n396 9.3005
R472 VTAIL.n395 VTAIL.n394 9.3005
R473 VTAIL.n354 VTAIL.n353 9.3005
R474 VTAIL.n369 VTAIL.n368 9.3005
R475 VTAIL.n371 VTAIL.n370 9.3005
R476 VTAIL.n362 VTAIL.n361 9.3005
R477 VTAIL.n377 VTAIL.n376 9.3005
R478 VTAIL.n379 VTAIL.n378 9.3005
R479 VTAIL.n358 VTAIL.n357 9.3005
R480 VTAIL.n386 VTAIL.n385 9.3005
R481 VTAIL.n388 VTAIL.n387 9.3005
R482 VTAIL.n413 VTAIL.n412 9.3005
R483 VTAIL.n342 VTAIL.n341 9.3005
R484 VTAIL.n419 VTAIL.n418 9.3005
R485 VTAIL.n421 VTAIL.n420 9.3005
R486 VTAIL.n338 VTAIL.n337 9.3005
R487 VTAIL.n427 VTAIL.n426 9.3005
R488 VTAIL.n429 VTAIL.n428 9.3005
R489 VTAIL.n334 VTAIL.n333 9.3005
R490 VTAIL.n435 VTAIL.n434 9.3005
R491 VTAIL.n81 VTAIL.n80 9.3005
R492 VTAIL.n16 VTAIL.n15 9.3005
R493 VTAIL.n75 VTAIL.n74 9.3005
R494 VTAIL.n73 VTAIL.n72 9.3005
R495 VTAIL.n20 VTAIL.n19 9.3005
R496 VTAIL.n67 VTAIL.n66 9.3005
R497 VTAIL.n65 VTAIL.n64 9.3005
R498 VTAIL.n24 VTAIL.n23 9.3005
R499 VTAIL.n39 VTAIL.n38 9.3005
R500 VTAIL.n41 VTAIL.n40 9.3005
R501 VTAIL.n32 VTAIL.n31 9.3005
R502 VTAIL.n47 VTAIL.n46 9.3005
R503 VTAIL.n49 VTAIL.n48 9.3005
R504 VTAIL.n28 VTAIL.n27 9.3005
R505 VTAIL.n56 VTAIL.n55 9.3005
R506 VTAIL.n58 VTAIL.n57 9.3005
R507 VTAIL.n83 VTAIL.n82 9.3005
R508 VTAIL.n12 VTAIL.n11 9.3005
R509 VTAIL.n89 VTAIL.n88 9.3005
R510 VTAIL.n91 VTAIL.n90 9.3005
R511 VTAIL.n8 VTAIL.n7 9.3005
R512 VTAIL.n97 VTAIL.n96 9.3005
R513 VTAIL.n99 VTAIL.n98 9.3005
R514 VTAIL.n4 VTAIL.n3 9.3005
R515 VTAIL.n105 VTAIL.n104 9.3005
R516 VTAIL.n264 VTAIL.n263 9.3005
R517 VTAIL.n266 VTAIL.n265 9.3005
R518 VTAIL.n257 VTAIL.n256 9.3005
R519 VTAIL.n272 VTAIL.n271 9.3005
R520 VTAIL.n274 VTAIL.n273 9.3005
R521 VTAIL.n252 VTAIL.n251 9.3005
R522 VTAIL.n280 VTAIL.n279 9.3005
R523 VTAIL.n282 VTAIL.n281 9.3005
R524 VTAIL.n236 VTAIL.n235 9.3005
R525 VTAIL.n313 VTAIL.n312 9.3005
R526 VTAIL.n315 VTAIL.n314 9.3005
R527 VTAIL.n232 VTAIL.n231 9.3005
R528 VTAIL.n321 VTAIL.n320 9.3005
R529 VTAIL.n323 VTAIL.n322 9.3005
R530 VTAIL.n228 VTAIL.n227 9.3005
R531 VTAIL.n329 VTAIL.n328 9.3005
R532 VTAIL.n307 VTAIL.n306 9.3005
R533 VTAIL.n305 VTAIL.n304 9.3005
R534 VTAIL.n240 VTAIL.n239 9.3005
R535 VTAIL.n299 VTAIL.n298 9.3005
R536 VTAIL.n297 VTAIL.n296 9.3005
R537 VTAIL.n244 VTAIL.n243 9.3005
R538 VTAIL.n291 VTAIL.n290 9.3005
R539 VTAIL.n289 VTAIL.n288 9.3005
R540 VTAIL.n248 VTAIL.n247 9.3005
R541 VTAIL.n154 VTAIL.n153 9.3005
R542 VTAIL.n156 VTAIL.n155 9.3005
R543 VTAIL.n147 VTAIL.n146 9.3005
R544 VTAIL.n162 VTAIL.n161 9.3005
R545 VTAIL.n164 VTAIL.n163 9.3005
R546 VTAIL.n142 VTAIL.n141 9.3005
R547 VTAIL.n170 VTAIL.n169 9.3005
R548 VTAIL.n172 VTAIL.n171 9.3005
R549 VTAIL.n126 VTAIL.n125 9.3005
R550 VTAIL.n203 VTAIL.n202 9.3005
R551 VTAIL.n205 VTAIL.n204 9.3005
R552 VTAIL.n122 VTAIL.n121 9.3005
R553 VTAIL.n211 VTAIL.n210 9.3005
R554 VTAIL.n213 VTAIL.n212 9.3005
R555 VTAIL.n118 VTAIL.n117 9.3005
R556 VTAIL.n219 VTAIL.n218 9.3005
R557 VTAIL.n197 VTAIL.n196 9.3005
R558 VTAIL.n195 VTAIL.n194 9.3005
R559 VTAIL.n130 VTAIL.n129 9.3005
R560 VTAIL.n189 VTAIL.n188 9.3005
R561 VTAIL.n187 VTAIL.n186 9.3005
R562 VTAIL.n134 VTAIL.n133 9.3005
R563 VTAIL.n181 VTAIL.n180 9.3005
R564 VTAIL.n179 VTAIL.n178 9.3005
R565 VTAIL.n138 VTAIL.n137 9.3005
R566 VTAIL.n372 VTAIL.n362 8.92171
R567 VTAIL.n406 VTAIL.n405 8.92171
R568 VTAIL.n421 VTAIL.n340 8.92171
R569 VTAIL.n42 VTAIL.n32 8.92171
R570 VTAIL.n76 VTAIL.n75 8.92171
R571 VTAIL.n91 VTAIL.n10 8.92171
R572 VTAIL.n315 VTAIL.n234 8.92171
R573 VTAIL.n300 VTAIL.n299 8.92171
R574 VTAIL.n267 VTAIL.n257 8.92171
R575 VTAIL.n205 VTAIL.n124 8.92171
R576 VTAIL.n190 VTAIL.n189 8.92171
R577 VTAIL.n157 VTAIL.n147 8.92171
R578 VTAIL.n371 VTAIL.n364 8.14595
R579 VTAIL.n409 VTAIL.n346 8.14595
R580 VTAIL.n418 VTAIL.n417 8.14595
R581 VTAIL.n41 VTAIL.n34 8.14595
R582 VTAIL.n79 VTAIL.n16 8.14595
R583 VTAIL.n88 VTAIL.n87 8.14595
R584 VTAIL.n312 VTAIL.n311 8.14595
R585 VTAIL.n303 VTAIL.n240 8.14595
R586 VTAIL.n266 VTAIL.n259 8.14595
R587 VTAIL.n202 VTAIL.n201 8.14595
R588 VTAIL.n193 VTAIL.n130 8.14595
R589 VTAIL.n156 VTAIL.n149 8.14595
R590 VTAIL.n436 VTAIL.n332 7.75445
R591 VTAIL.n106 VTAIL.n2 7.75445
R592 VTAIL.n330 VTAIL.n226 7.75445
R593 VTAIL.n220 VTAIL.n116 7.75445
R594 VTAIL.n368 VTAIL.n367 7.3702
R595 VTAIL.n410 VTAIL.n344 7.3702
R596 VTAIL.n414 VTAIL.n342 7.3702
R597 VTAIL.n38 VTAIL.n37 7.3702
R598 VTAIL.n80 VTAIL.n14 7.3702
R599 VTAIL.n84 VTAIL.n12 7.3702
R600 VTAIL.n308 VTAIL.n236 7.3702
R601 VTAIL.n304 VTAIL.n238 7.3702
R602 VTAIL.n263 VTAIL.n262 7.3702
R603 VTAIL.n198 VTAIL.n126 7.3702
R604 VTAIL.n194 VTAIL.n128 7.3702
R605 VTAIL.n153 VTAIL.n152 7.3702
R606 VTAIL.n413 VTAIL.n344 6.59444
R607 VTAIL.n414 VTAIL.n413 6.59444
R608 VTAIL.n83 VTAIL.n14 6.59444
R609 VTAIL.n84 VTAIL.n83 6.59444
R610 VTAIL.n308 VTAIL.n307 6.59444
R611 VTAIL.n307 VTAIL.n238 6.59444
R612 VTAIL.n198 VTAIL.n197 6.59444
R613 VTAIL.n197 VTAIL.n128 6.59444
R614 VTAIL.n434 VTAIL.n332 6.08283
R615 VTAIL.n104 VTAIL.n2 6.08283
R616 VTAIL.n328 VTAIL.n226 6.08283
R617 VTAIL.n218 VTAIL.n116 6.08283
R618 VTAIL.n368 VTAIL.n364 5.81868
R619 VTAIL.n410 VTAIL.n409 5.81868
R620 VTAIL.n417 VTAIL.n342 5.81868
R621 VTAIL.n38 VTAIL.n34 5.81868
R622 VTAIL.n80 VTAIL.n79 5.81868
R623 VTAIL.n87 VTAIL.n12 5.81868
R624 VTAIL.n311 VTAIL.n236 5.81868
R625 VTAIL.n304 VTAIL.n303 5.81868
R626 VTAIL.n263 VTAIL.n259 5.81868
R627 VTAIL.n201 VTAIL.n126 5.81868
R628 VTAIL.n194 VTAIL.n193 5.81868
R629 VTAIL.n153 VTAIL.n149 5.81868
R630 VTAIL.n372 VTAIL.n371 5.04292
R631 VTAIL.n406 VTAIL.n346 5.04292
R632 VTAIL.n418 VTAIL.n340 5.04292
R633 VTAIL.n42 VTAIL.n41 5.04292
R634 VTAIL.n76 VTAIL.n16 5.04292
R635 VTAIL.n88 VTAIL.n10 5.04292
R636 VTAIL.n312 VTAIL.n234 5.04292
R637 VTAIL.n300 VTAIL.n240 5.04292
R638 VTAIL.n267 VTAIL.n266 5.04292
R639 VTAIL.n202 VTAIL.n124 5.04292
R640 VTAIL.n190 VTAIL.n130 5.04292
R641 VTAIL.n157 VTAIL.n156 5.04292
R642 VTAIL.n375 VTAIL.n362 4.26717
R643 VTAIL.n405 VTAIL.n348 4.26717
R644 VTAIL.n422 VTAIL.n421 4.26717
R645 VTAIL.n45 VTAIL.n32 4.26717
R646 VTAIL.n75 VTAIL.n18 4.26717
R647 VTAIL.n92 VTAIL.n91 4.26717
R648 VTAIL.n316 VTAIL.n315 4.26717
R649 VTAIL.n299 VTAIL.n242 4.26717
R650 VTAIL.n270 VTAIL.n257 4.26717
R651 VTAIL.n206 VTAIL.n205 4.26717
R652 VTAIL.n189 VTAIL.n132 4.26717
R653 VTAIL.n160 VTAIL.n147 4.26717
R654 VTAIL.n376 VTAIL.n360 3.49141
R655 VTAIL.n402 VTAIL.n401 3.49141
R656 VTAIL.n425 VTAIL.n338 3.49141
R657 VTAIL.n46 VTAIL.n30 3.49141
R658 VTAIL.n72 VTAIL.n71 3.49141
R659 VTAIL.n95 VTAIL.n8 3.49141
R660 VTAIL.n319 VTAIL.n232 3.49141
R661 VTAIL.n296 VTAIL.n295 3.49141
R662 VTAIL.n271 VTAIL.n255 3.49141
R663 VTAIL.n209 VTAIL.n122 3.49141
R664 VTAIL.n186 VTAIL.n185 3.49141
R665 VTAIL.n161 VTAIL.n145 3.49141
R666 VTAIL.n115 VTAIL.n113 2.96602
R667 VTAIL.n221 VTAIL.n115 2.96602
R668 VTAIL.n225 VTAIL.n223 2.96602
R669 VTAIL.n331 VTAIL.n225 2.96602
R670 VTAIL.n111 VTAIL.n109 2.96602
R671 VTAIL.n109 VTAIL.n107 2.96602
R672 VTAIL.n439 VTAIL.n437 2.96602
R673 VTAIL.n380 VTAIL.n379 2.71565
R674 VTAIL.n398 VTAIL.n350 2.71565
R675 VTAIL.n426 VTAIL.n336 2.71565
R676 VTAIL.n50 VTAIL.n49 2.71565
R677 VTAIL.n68 VTAIL.n20 2.71565
R678 VTAIL.n96 VTAIL.n6 2.71565
R679 VTAIL.n320 VTAIL.n230 2.71565
R680 VTAIL.n292 VTAIL.n244 2.71565
R681 VTAIL.n275 VTAIL.n274 2.71565
R682 VTAIL.n210 VTAIL.n120 2.71565
R683 VTAIL.n182 VTAIL.n134 2.71565
R684 VTAIL.n165 VTAIL.n164 2.71565
R685 VTAIL.n264 VTAIL.n260 2.41282
R686 VTAIL.n154 VTAIL.n150 2.41282
R687 VTAIL.n369 VTAIL.n365 2.41282
R688 VTAIL.n39 VTAIL.n35 2.41282
R689 VTAIL VTAIL.n1 2.28283
R690 VTAIL.n223 VTAIL.n221 1.95309
R691 VTAIL.n107 VTAIL.n1 1.95309
R692 VTAIL.n384 VTAIL.n358 1.93989
R693 VTAIL.n397 VTAIL.n352 1.93989
R694 VTAIL.n430 VTAIL.n429 1.93989
R695 VTAIL.n54 VTAIL.n28 1.93989
R696 VTAIL.n67 VTAIL.n22 1.93989
R697 VTAIL.n100 VTAIL.n99 1.93989
R698 VTAIL.n324 VTAIL.n323 1.93989
R699 VTAIL.n291 VTAIL.n246 1.93989
R700 VTAIL.n278 VTAIL.n252 1.93989
R701 VTAIL.n214 VTAIL.n213 1.93989
R702 VTAIL.n181 VTAIL.n136 1.93989
R703 VTAIL.n168 VTAIL.n142 1.93989
R704 VTAIL.n438 VTAIL.t15 1.67515
R705 VTAIL.n438 VTAIL.t0 1.67515
R706 VTAIL.n0 VTAIL.t17 1.67515
R707 VTAIL.n0 VTAIL.t19 1.67515
R708 VTAIL.n108 VTAIL.t11 1.67515
R709 VTAIL.n108 VTAIL.t5 1.67515
R710 VTAIL.n110 VTAIL.t12 1.67515
R711 VTAIL.n110 VTAIL.t9 1.67515
R712 VTAIL.n224 VTAIL.t6 1.67515
R713 VTAIL.n224 VTAIL.t4 1.67515
R714 VTAIL.n222 VTAIL.t8 1.67515
R715 VTAIL.n222 VTAIL.t13 1.67515
R716 VTAIL.n114 VTAIL.t14 1.67515
R717 VTAIL.n114 VTAIL.t3 1.67515
R718 VTAIL.n112 VTAIL.t16 1.67515
R719 VTAIL.n112 VTAIL.t2 1.67515
R720 VTAIL.n385 VTAIL.n356 1.16414
R721 VTAIL.n394 VTAIL.n393 1.16414
R722 VTAIL.n433 VTAIL.n334 1.16414
R723 VTAIL.n55 VTAIL.n26 1.16414
R724 VTAIL.n64 VTAIL.n63 1.16414
R725 VTAIL.n103 VTAIL.n4 1.16414
R726 VTAIL.n327 VTAIL.n228 1.16414
R727 VTAIL.n288 VTAIL.n287 1.16414
R728 VTAIL.n279 VTAIL.n250 1.16414
R729 VTAIL.n217 VTAIL.n118 1.16414
R730 VTAIL.n178 VTAIL.n177 1.16414
R731 VTAIL.n169 VTAIL.n140 1.16414
R732 VTAIL VTAIL.n439 0.68369
R733 VTAIL.n389 VTAIL.n388 0.388379
R734 VTAIL.n390 VTAIL.n354 0.388379
R735 VTAIL.n59 VTAIL.n58 0.388379
R736 VTAIL.n60 VTAIL.n24 0.388379
R737 VTAIL.n284 VTAIL.n248 0.388379
R738 VTAIL.n283 VTAIL.n282 0.388379
R739 VTAIL.n174 VTAIL.n138 0.388379
R740 VTAIL.n173 VTAIL.n172 0.388379
R741 VTAIL.n370 VTAIL.n369 0.155672
R742 VTAIL.n370 VTAIL.n361 0.155672
R743 VTAIL.n377 VTAIL.n361 0.155672
R744 VTAIL.n378 VTAIL.n377 0.155672
R745 VTAIL.n378 VTAIL.n357 0.155672
R746 VTAIL.n386 VTAIL.n357 0.155672
R747 VTAIL.n387 VTAIL.n386 0.155672
R748 VTAIL.n387 VTAIL.n353 0.155672
R749 VTAIL.n395 VTAIL.n353 0.155672
R750 VTAIL.n396 VTAIL.n395 0.155672
R751 VTAIL.n396 VTAIL.n349 0.155672
R752 VTAIL.n403 VTAIL.n349 0.155672
R753 VTAIL.n404 VTAIL.n403 0.155672
R754 VTAIL.n404 VTAIL.n345 0.155672
R755 VTAIL.n411 VTAIL.n345 0.155672
R756 VTAIL.n412 VTAIL.n411 0.155672
R757 VTAIL.n412 VTAIL.n341 0.155672
R758 VTAIL.n419 VTAIL.n341 0.155672
R759 VTAIL.n420 VTAIL.n419 0.155672
R760 VTAIL.n420 VTAIL.n337 0.155672
R761 VTAIL.n427 VTAIL.n337 0.155672
R762 VTAIL.n428 VTAIL.n427 0.155672
R763 VTAIL.n428 VTAIL.n333 0.155672
R764 VTAIL.n435 VTAIL.n333 0.155672
R765 VTAIL.n40 VTAIL.n39 0.155672
R766 VTAIL.n40 VTAIL.n31 0.155672
R767 VTAIL.n47 VTAIL.n31 0.155672
R768 VTAIL.n48 VTAIL.n47 0.155672
R769 VTAIL.n48 VTAIL.n27 0.155672
R770 VTAIL.n56 VTAIL.n27 0.155672
R771 VTAIL.n57 VTAIL.n56 0.155672
R772 VTAIL.n57 VTAIL.n23 0.155672
R773 VTAIL.n65 VTAIL.n23 0.155672
R774 VTAIL.n66 VTAIL.n65 0.155672
R775 VTAIL.n66 VTAIL.n19 0.155672
R776 VTAIL.n73 VTAIL.n19 0.155672
R777 VTAIL.n74 VTAIL.n73 0.155672
R778 VTAIL.n74 VTAIL.n15 0.155672
R779 VTAIL.n81 VTAIL.n15 0.155672
R780 VTAIL.n82 VTAIL.n81 0.155672
R781 VTAIL.n82 VTAIL.n11 0.155672
R782 VTAIL.n89 VTAIL.n11 0.155672
R783 VTAIL.n90 VTAIL.n89 0.155672
R784 VTAIL.n90 VTAIL.n7 0.155672
R785 VTAIL.n97 VTAIL.n7 0.155672
R786 VTAIL.n98 VTAIL.n97 0.155672
R787 VTAIL.n98 VTAIL.n3 0.155672
R788 VTAIL.n105 VTAIL.n3 0.155672
R789 VTAIL.n329 VTAIL.n227 0.155672
R790 VTAIL.n322 VTAIL.n227 0.155672
R791 VTAIL.n322 VTAIL.n321 0.155672
R792 VTAIL.n321 VTAIL.n231 0.155672
R793 VTAIL.n314 VTAIL.n231 0.155672
R794 VTAIL.n314 VTAIL.n313 0.155672
R795 VTAIL.n313 VTAIL.n235 0.155672
R796 VTAIL.n306 VTAIL.n235 0.155672
R797 VTAIL.n306 VTAIL.n305 0.155672
R798 VTAIL.n305 VTAIL.n239 0.155672
R799 VTAIL.n298 VTAIL.n239 0.155672
R800 VTAIL.n298 VTAIL.n297 0.155672
R801 VTAIL.n297 VTAIL.n243 0.155672
R802 VTAIL.n290 VTAIL.n243 0.155672
R803 VTAIL.n290 VTAIL.n289 0.155672
R804 VTAIL.n289 VTAIL.n247 0.155672
R805 VTAIL.n281 VTAIL.n247 0.155672
R806 VTAIL.n281 VTAIL.n280 0.155672
R807 VTAIL.n280 VTAIL.n251 0.155672
R808 VTAIL.n273 VTAIL.n251 0.155672
R809 VTAIL.n273 VTAIL.n272 0.155672
R810 VTAIL.n272 VTAIL.n256 0.155672
R811 VTAIL.n265 VTAIL.n256 0.155672
R812 VTAIL.n265 VTAIL.n264 0.155672
R813 VTAIL.n219 VTAIL.n117 0.155672
R814 VTAIL.n212 VTAIL.n117 0.155672
R815 VTAIL.n212 VTAIL.n211 0.155672
R816 VTAIL.n211 VTAIL.n121 0.155672
R817 VTAIL.n204 VTAIL.n121 0.155672
R818 VTAIL.n204 VTAIL.n203 0.155672
R819 VTAIL.n203 VTAIL.n125 0.155672
R820 VTAIL.n196 VTAIL.n125 0.155672
R821 VTAIL.n196 VTAIL.n195 0.155672
R822 VTAIL.n195 VTAIL.n129 0.155672
R823 VTAIL.n188 VTAIL.n129 0.155672
R824 VTAIL.n188 VTAIL.n187 0.155672
R825 VTAIL.n187 VTAIL.n133 0.155672
R826 VTAIL.n180 VTAIL.n133 0.155672
R827 VTAIL.n180 VTAIL.n179 0.155672
R828 VTAIL.n179 VTAIL.n137 0.155672
R829 VTAIL.n171 VTAIL.n137 0.155672
R830 VTAIL.n171 VTAIL.n170 0.155672
R831 VTAIL.n170 VTAIL.n141 0.155672
R832 VTAIL.n163 VTAIL.n141 0.155672
R833 VTAIL.n163 VTAIL.n162 0.155672
R834 VTAIL.n162 VTAIL.n146 0.155672
R835 VTAIL.n155 VTAIL.n146 0.155672
R836 VTAIL.n155 VTAIL.n154 0.155672
R837 VDD1.n101 VDD1.n100 585
R838 VDD1.n99 VDD1.n98 585
R839 VDD1.n4 VDD1.n3 585
R840 VDD1.n93 VDD1.n92 585
R841 VDD1.n91 VDD1.n90 585
R842 VDD1.n8 VDD1.n7 585
R843 VDD1.n85 VDD1.n84 585
R844 VDD1.n83 VDD1.n82 585
R845 VDD1.n12 VDD1.n11 585
R846 VDD1.n77 VDD1.n76 585
R847 VDD1.n75 VDD1.n74 585
R848 VDD1.n16 VDD1.n15 585
R849 VDD1.n69 VDD1.n68 585
R850 VDD1.n67 VDD1.n66 585
R851 VDD1.n20 VDD1.n19 585
R852 VDD1.n61 VDD1.n60 585
R853 VDD1.n59 VDD1.n58 585
R854 VDD1.n57 VDD1.n23 585
R855 VDD1.n27 VDD1.n24 585
R856 VDD1.n52 VDD1.n51 585
R857 VDD1.n50 VDD1.n49 585
R858 VDD1.n29 VDD1.n28 585
R859 VDD1.n44 VDD1.n43 585
R860 VDD1.n42 VDD1.n41 585
R861 VDD1.n33 VDD1.n32 585
R862 VDD1.n36 VDD1.n35 585
R863 VDD1.n142 VDD1.n141 585
R864 VDD1.n139 VDD1.n138 585
R865 VDD1.n148 VDD1.n147 585
R866 VDD1.n150 VDD1.n149 585
R867 VDD1.n135 VDD1.n134 585
R868 VDD1.n156 VDD1.n155 585
R869 VDD1.n159 VDD1.n158 585
R870 VDD1.n157 VDD1.n131 585
R871 VDD1.n164 VDD1.n130 585
R872 VDD1.n166 VDD1.n165 585
R873 VDD1.n168 VDD1.n167 585
R874 VDD1.n127 VDD1.n126 585
R875 VDD1.n174 VDD1.n173 585
R876 VDD1.n176 VDD1.n175 585
R877 VDD1.n123 VDD1.n122 585
R878 VDD1.n182 VDD1.n181 585
R879 VDD1.n184 VDD1.n183 585
R880 VDD1.n119 VDD1.n118 585
R881 VDD1.n190 VDD1.n189 585
R882 VDD1.n192 VDD1.n191 585
R883 VDD1.n115 VDD1.n114 585
R884 VDD1.n198 VDD1.n197 585
R885 VDD1.n200 VDD1.n199 585
R886 VDD1.n111 VDD1.n110 585
R887 VDD1.n206 VDD1.n205 585
R888 VDD1.n208 VDD1.n207 585
R889 VDD1.n100 VDD1.n0 498.474
R890 VDD1.n207 VDD1.n107 498.474
R891 VDD1.t7 VDD1.n34 329.036
R892 VDD1.t2 VDD1.n140 329.036
R893 VDD1.n100 VDD1.n99 171.744
R894 VDD1.n99 VDD1.n3 171.744
R895 VDD1.n92 VDD1.n3 171.744
R896 VDD1.n92 VDD1.n91 171.744
R897 VDD1.n91 VDD1.n7 171.744
R898 VDD1.n84 VDD1.n7 171.744
R899 VDD1.n84 VDD1.n83 171.744
R900 VDD1.n83 VDD1.n11 171.744
R901 VDD1.n76 VDD1.n11 171.744
R902 VDD1.n76 VDD1.n75 171.744
R903 VDD1.n75 VDD1.n15 171.744
R904 VDD1.n68 VDD1.n15 171.744
R905 VDD1.n68 VDD1.n67 171.744
R906 VDD1.n67 VDD1.n19 171.744
R907 VDD1.n60 VDD1.n19 171.744
R908 VDD1.n60 VDD1.n59 171.744
R909 VDD1.n59 VDD1.n23 171.744
R910 VDD1.n27 VDD1.n23 171.744
R911 VDD1.n51 VDD1.n27 171.744
R912 VDD1.n51 VDD1.n50 171.744
R913 VDD1.n50 VDD1.n28 171.744
R914 VDD1.n43 VDD1.n28 171.744
R915 VDD1.n43 VDD1.n42 171.744
R916 VDD1.n42 VDD1.n32 171.744
R917 VDD1.n35 VDD1.n32 171.744
R918 VDD1.n141 VDD1.n138 171.744
R919 VDD1.n148 VDD1.n138 171.744
R920 VDD1.n149 VDD1.n148 171.744
R921 VDD1.n149 VDD1.n134 171.744
R922 VDD1.n156 VDD1.n134 171.744
R923 VDD1.n158 VDD1.n156 171.744
R924 VDD1.n158 VDD1.n157 171.744
R925 VDD1.n157 VDD1.n130 171.744
R926 VDD1.n166 VDD1.n130 171.744
R927 VDD1.n167 VDD1.n166 171.744
R928 VDD1.n167 VDD1.n126 171.744
R929 VDD1.n174 VDD1.n126 171.744
R930 VDD1.n175 VDD1.n174 171.744
R931 VDD1.n175 VDD1.n122 171.744
R932 VDD1.n182 VDD1.n122 171.744
R933 VDD1.n183 VDD1.n182 171.744
R934 VDD1.n183 VDD1.n118 171.744
R935 VDD1.n190 VDD1.n118 171.744
R936 VDD1.n191 VDD1.n190 171.744
R937 VDD1.n191 VDD1.n114 171.744
R938 VDD1.n198 VDD1.n114 171.744
R939 VDD1.n199 VDD1.n198 171.744
R940 VDD1.n199 VDD1.n110 171.744
R941 VDD1.n206 VDD1.n110 171.744
R942 VDD1.n207 VDD1.n206 171.744
R943 VDD1.n35 VDD1.t7 85.8723
R944 VDD1.n141 VDD1.t2 85.8723
R945 VDD1.n215 VDD1.n214 71.7573
R946 VDD1.n106 VDD1.n105 69.5887
R947 VDD1.n217 VDD1.n216 69.5885
R948 VDD1.n213 VDD1.n212 69.5885
R949 VDD1.n217 VDD1.n215 56.6
R950 VDD1.n106 VDD1.n104 53.5751
R951 VDD1.n213 VDD1.n211 53.5751
R952 VDD1.n58 VDD1.n57 13.1884
R953 VDD1.n165 VDD1.n164 13.1884
R954 VDD1.n102 VDD1.n101 12.8005
R955 VDD1.n61 VDD1.n22 12.8005
R956 VDD1.n56 VDD1.n24 12.8005
R957 VDD1.n163 VDD1.n131 12.8005
R958 VDD1.n168 VDD1.n129 12.8005
R959 VDD1.n209 VDD1.n208 12.8005
R960 VDD1.n98 VDD1.n2 12.0247
R961 VDD1.n62 VDD1.n20 12.0247
R962 VDD1.n53 VDD1.n52 12.0247
R963 VDD1.n160 VDD1.n159 12.0247
R964 VDD1.n169 VDD1.n127 12.0247
R965 VDD1.n205 VDD1.n109 12.0247
R966 VDD1.n97 VDD1.n4 11.249
R967 VDD1.n66 VDD1.n65 11.249
R968 VDD1.n49 VDD1.n26 11.249
R969 VDD1.n155 VDD1.n133 11.249
R970 VDD1.n173 VDD1.n172 11.249
R971 VDD1.n204 VDD1.n111 11.249
R972 VDD1.n36 VDD1.n34 10.7239
R973 VDD1.n142 VDD1.n140 10.7239
R974 VDD1.n94 VDD1.n93 10.4732
R975 VDD1.n69 VDD1.n18 10.4732
R976 VDD1.n48 VDD1.n29 10.4732
R977 VDD1.n154 VDD1.n135 10.4732
R978 VDD1.n176 VDD1.n125 10.4732
R979 VDD1.n201 VDD1.n200 10.4732
R980 VDD1.n90 VDD1.n6 9.69747
R981 VDD1.n70 VDD1.n16 9.69747
R982 VDD1.n45 VDD1.n44 9.69747
R983 VDD1.n151 VDD1.n150 9.69747
R984 VDD1.n177 VDD1.n123 9.69747
R985 VDD1.n197 VDD1.n113 9.69747
R986 VDD1.n104 VDD1.n103 9.45567
R987 VDD1.n211 VDD1.n210 9.45567
R988 VDD1.n38 VDD1.n37 9.3005
R989 VDD1.n40 VDD1.n39 9.3005
R990 VDD1.n31 VDD1.n30 9.3005
R991 VDD1.n46 VDD1.n45 9.3005
R992 VDD1.n48 VDD1.n47 9.3005
R993 VDD1.n26 VDD1.n25 9.3005
R994 VDD1.n54 VDD1.n53 9.3005
R995 VDD1.n56 VDD1.n55 9.3005
R996 VDD1.n10 VDD1.n9 9.3005
R997 VDD1.n87 VDD1.n86 9.3005
R998 VDD1.n89 VDD1.n88 9.3005
R999 VDD1.n6 VDD1.n5 9.3005
R1000 VDD1.n95 VDD1.n94 9.3005
R1001 VDD1.n97 VDD1.n96 9.3005
R1002 VDD1.n2 VDD1.n1 9.3005
R1003 VDD1.n103 VDD1.n102 9.3005
R1004 VDD1.n81 VDD1.n80 9.3005
R1005 VDD1.n79 VDD1.n78 9.3005
R1006 VDD1.n14 VDD1.n13 9.3005
R1007 VDD1.n73 VDD1.n72 9.3005
R1008 VDD1.n71 VDD1.n70 9.3005
R1009 VDD1.n18 VDD1.n17 9.3005
R1010 VDD1.n65 VDD1.n64 9.3005
R1011 VDD1.n63 VDD1.n62 9.3005
R1012 VDD1.n22 VDD1.n21 9.3005
R1013 VDD1.n186 VDD1.n185 9.3005
R1014 VDD1.n121 VDD1.n120 9.3005
R1015 VDD1.n180 VDD1.n179 9.3005
R1016 VDD1.n178 VDD1.n177 9.3005
R1017 VDD1.n125 VDD1.n124 9.3005
R1018 VDD1.n172 VDD1.n171 9.3005
R1019 VDD1.n170 VDD1.n169 9.3005
R1020 VDD1.n129 VDD1.n128 9.3005
R1021 VDD1.n144 VDD1.n143 9.3005
R1022 VDD1.n146 VDD1.n145 9.3005
R1023 VDD1.n137 VDD1.n136 9.3005
R1024 VDD1.n152 VDD1.n151 9.3005
R1025 VDD1.n154 VDD1.n153 9.3005
R1026 VDD1.n133 VDD1.n132 9.3005
R1027 VDD1.n161 VDD1.n160 9.3005
R1028 VDD1.n163 VDD1.n162 9.3005
R1029 VDD1.n188 VDD1.n187 9.3005
R1030 VDD1.n117 VDD1.n116 9.3005
R1031 VDD1.n194 VDD1.n193 9.3005
R1032 VDD1.n196 VDD1.n195 9.3005
R1033 VDD1.n113 VDD1.n112 9.3005
R1034 VDD1.n202 VDD1.n201 9.3005
R1035 VDD1.n204 VDD1.n203 9.3005
R1036 VDD1.n109 VDD1.n108 9.3005
R1037 VDD1.n210 VDD1.n209 9.3005
R1038 VDD1.n89 VDD1.n8 8.92171
R1039 VDD1.n74 VDD1.n73 8.92171
R1040 VDD1.n41 VDD1.n31 8.92171
R1041 VDD1.n147 VDD1.n137 8.92171
R1042 VDD1.n181 VDD1.n180 8.92171
R1043 VDD1.n196 VDD1.n115 8.92171
R1044 VDD1.n86 VDD1.n85 8.14595
R1045 VDD1.n77 VDD1.n14 8.14595
R1046 VDD1.n40 VDD1.n33 8.14595
R1047 VDD1.n146 VDD1.n139 8.14595
R1048 VDD1.n184 VDD1.n121 8.14595
R1049 VDD1.n193 VDD1.n192 8.14595
R1050 VDD1.n104 VDD1.n0 7.75445
R1051 VDD1.n211 VDD1.n107 7.75445
R1052 VDD1.n82 VDD1.n10 7.3702
R1053 VDD1.n78 VDD1.n12 7.3702
R1054 VDD1.n37 VDD1.n36 7.3702
R1055 VDD1.n143 VDD1.n142 7.3702
R1056 VDD1.n185 VDD1.n119 7.3702
R1057 VDD1.n189 VDD1.n117 7.3702
R1058 VDD1.n82 VDD1.n81 6.59444
R1059 VDD1.n81 VDD1.n12 6.59444
R1060 VDD1.n188 VDD1.n119 6.59444
R1061 VDD1.n189 VDD1.n188 6.59444
R1062 VDD1.n102 VDD1.n0 6.08283
R1063 VDD1.n209 VDD1.n107 6.08283
R1064 VDD1.n85 VDD1.n10 5.81868
R1065 VDD1.n78 VDD1.n77 5.81868
R1066 VDD1.n37 VDD1.n33 5.81868
R1067 VDD1.n143 VDD1.n139 5.81868
R1068 VDD1.n185 VDD1.n184 5.81868
R1069 VDD1.n192 VDD1.n117 5.81868
R1070 VDD1.n86 VDD1.n8 5.04292
R1071 VDD1.n74 VDD1.n14 5.04292
R1072 VDD1.n41 VDD1.n40 5.04292
R1073 VDD1.n147 VDD1.n146 5.04292
R1074 VDD1.n181 VDD1.n121 5.04292
R1075 VDD1.n193 VDD1.n115 5.04292
R1076 VDD1.n90 VDD1.n89 4.26717
R1077 VDD1.n73 VDD1.n16 4.26717
R1078 VDD1.n44 VDD1.n31 4.26717
R1079 VDD1.n150 VDD1.n137 4.26717
R1080 VDD1.n180 VDD1.n123 4.26717
R1081 VDD1.n197 VDD1.n196 4.26717
R1082 VDD1.n93 VDD1.n6 3.49141
R1083 VDD1.n70 VDD1.n69 3.49141
R1084 VDD1.n45 VDD1.n29 3.49141
R1085 VDD1.n151 VDD1.n135 3.49141
R1086 VDD1.n177 VDD1.n176 3.49141
R1087 VDD1.n200 VDD1.n113 3.49141
R1088 VDD1.n94 VDD1.n4 2.71565
R1089 VDD1.n66 VDD1.n18 2.71565
R1090 VDD1.n49 VDD1.n48 2.71565
R1091 VDD1.n155 VDD1.n154 2.71565
R1092 VDD1.n173 VDD1.n125 2.71565
R1093 VDD1.n201 VDD1.n111 2.71565
R1094 VDD1.n38 VDD1.n34 2.41282
R1095 VDD1.n144 VDD1.n140 2.41282
R1096 VDD1 VDD1.n217 2.16645
R1097 VDD1.n98 VDD1.n97 1.93989
R1098 VDD1.n65 VDD1.n20 1.93989
R1099 VDD1.n52 VDD1.n26 1.93989
R1100 VDD1.n159 VDD1.n133 1.93989
R1101 VDD1.n172 VDD1.n127 1.93989
R1102 VDD1.n205 VDD1.n204 1.93989
R1103 VDD1.n216 VDD1.t5 1.67515
R1104 VDD1.n216 VDD1.t9 1.67515
R1105 VDD1.n105 VDD1.t8 1.67515
R1106 VDD1.n105 VDD1.t3 1.67515
R1107 VDD1.n214 VDD1.t4 1.67515
R1108 VDD1.n214 VDD1.t6 1.67515
R1109 VDD1.n212 VDD1.t0 1.67515
R1110 VDD1.n212 VDD1.t1 1.67515
R1111 VDD1.n101 VDD1.n2 1.16414
R1112 VDD1.n62 VDD1.n61 1.16414
R1113 VDD1.n53 VDD1.n24 1.16414
R1114 VDD1.n160 VDD1.n131 1.16414
R1115 VDD1.n169 VDD1.n168 1.16414
R1116 VDD1.n208 VDD1.n109 1.16414
R1117 VDD1 VDD1.n106 0.800069
R1118 VDD1.n215 VDD1.n213 0.686533
R1119 VDD1.n58 VDD1.n22 0.388379
R1120 VDD1.n57 VDD1.n56 0.388379
R1121 VDD1.n164 VDD1.n163 0.388379
R1122 VDD1.n165 VDD1.n129 0.388379
R1123 VDD1.n103 VDD1.n1 0.155672
R1124 VDD1.n96 VDD1.n1 0.155672
R1125 VDD1.n96 VDD1.n95 0.155672
R1126 VDD1.n95 VDD1.n5 0.155672
R1127 VDD1.n88 VDD1.n5 0.155672
R1128 VDD1.n88 VDD1.n87 0.155672
R1129 VDD1.n87 VDD1.n9 0.155672
R1130 VDD1.n80 VDD1.n9 0.155672
R1131 VDD1.n80 VDD1.n79 0.155672
R1132 VDD1.n79 VDD1.n13 0.155672
R1133 VDD1.n72 VDD1.n13 0.155672
R1134 VDD1.n72 VDD1.n71 0.155672
R1135 VDD1.n71 VDD1.n17 0.155672
R1136 VDD1.n64 VDD1.n17 0.155672
R1137 VDD1.n64 VDD1.n63 0.155672
R1138 VDD1.n63 VDD1.n21 0.155672
R1139 VDD1.n55 VDD1.n21 0.155672
R1140 VDD1.n55 VDD1.n54 0.155672
R1141 VDD1.n54 VDD1.n25 0.155672
R1142 VDD1.n47 VDD1.n25 0.155672
R1143 VDD1.n47 VDD1.n46 0.155672
R1144 VDD1.n46 VDD1.n30 0.155672
R1145 VDD1.n39 VDD1.n30 0.155672
R1146 VDD1.n39 VDD1.n38 0.155672
R1147 VDD1.n145 VDD1.n144 0.155672
R1148 VDD1.n145 VDD1.n136 0.155672
R1149 VDD1.n152 VDD1.n136 0.155672
R1150 VDD1.n153 VDD1.n152 0.155672
R1151 VDD1.n153 VDD1.n132 0.155672
R1152 VDD1.n161 VDD1.n132 0.155672
R1153 VDD1.n162 VDD1.n161 0.155672
R1154 VDD1.n162 VDD1.n128 0.155672
R1155 VDD1.n170 VDD1.n128 0.155672
R1156 VDD1.n171 VDD1.n170 0.155672
R1157 VDD1.n171 VDD1.n124 0.155672
R1158 VDD1.n178 VDD1.n124 0.155672
R1159 VDD1.n179 VDD1.n178 0.155672
R1160 VDD1.n179 VDD1.n120 0.155672
R1161 VDD1.n186 VDD1.n120 0.155672
R1162 VDD1.n187 VDD1.n186 0.155672
R1163 VDD1.n187 VDD1.n116 0.155672
R1164 VDD1.n194 VDD1.n116 0.155672
R1165 VDD1.n195 VDD1.n194 0.155672
R1166 VDD1.n195 VDD1.n112 0.155672
R1167 VDD1.n202 VDD1.n112 0.155672
R1168 VDD1.n203 VDD1.n202 0.155672
R1169 VDD1.n203 VDD1.n108 0.155672
R1170 VDD1.n210 VDD1.n108 0.155672
R1171 VN.n56 VN.t5 183.764
R1172 VN.n11 VN.t0 183.764
R1173 VN.n88 VN.n87 161.3
R1174 VN.n86 VN.n46 161.3
R1175 VN.n85 VN.n84 161.3
R1176 VN.n83 VN.n47 161.3
R1177 VN.n82 VN.n81 161.3
R1178 VN.n80 VN.n48 161.3
R1179 VN.n79 VN.n78 161.3
R1180 VN.n77 VN.n76 161.3
R1181 VN.n75 VN.n50 161.3
R1182 VN.n74 VN.n73 161.3
R1183 VN.n72 VN.n51 161.3
R1184 VN.n71 VN.n70 161.3
R1185 VN.n69 VN.n52 161.3
R1186 VN.n68 VN.n67 161.3
R1187 VN.n66 VN.n53 161.3
R1188 VN.n65 VN.n64 161.3
R1189 VN.n63 VN.n54 161.3
R1190 VN.n62 VN.n61 161.3
R1191 VN.n60 VN.n55 161.3
R1192 VN.n59 VN.n58 161.3
R1193 VN.n43 VN.n42 161.3
R1194 VN.n41 VN.n1 161.3
R1195 VN.n40 VN.n39 161.3
R1196 VN.n38 VN.n2 161.3
R1197 VN.n37 VN.n36 161.3
R1198 VN.n35 VN.n3 161.3
R1199 VN.n34 VN.n33 161.3
R1200 VN.n32 VN.n31 161.3
R1201 VN.n30 VN.n5 161.3
R1202 VN.n29 VN.n28 161.3
R1203 VN.n27 VN.n6 161.3
R1204 VN.n26 VN.n25 161.3
R1205 VN.n24 VN.n7 161.3
R1206 VN.n23 VN.n22 161.3
R1207 VN.n21 VN.n8 161.3
R1208 VN.n20 VN.n19 161.3
R1209 VN.n18 VN.n9 161.3
R1210 VN.n17 VN.n16 161.3
R1211 VN.n15 VN.n10 161.3
R1212 VN.n14 VN.n13 161.3
R1213 VN.n23 VN.t6 150.412
R1214 VN.n12 VN.t4 150.412
R1215 VN.n4 VN.t8 150.412
R1216 VN.n0 VN.t9 150.412
R1217 VN.n68 VN.t1 150.412
R1218 VN.n57 VN.t2 150.412
R1219 VN.n49 VN.t7 150.412
R1220 VN.n45 VN.t3 150.412
R1221 VN.n44 VN.n0 71.4725
R1222 VN.n89 VN.n45 71.4725
R1223 VN VN.n89 61.7935
R1224 VN.n18 VN.n17 56.5193
R1225 VN.n29 VN.n6 56.5193
R1226 VN.n63 VN.n62 56.5193
R1227 VN.n74 VN.n51 56.5193
R1228 VN.n40 VN.n2 56.0336
R1229 VN.n85 VN.n47 56.0336
R1230 VN.n12 VN.n11 52.2938
R1231 VN.n57 VN.n56 52.2938
R1232 VN.n36 VN.n2 24.9531
R1233 VN.n81 VN.n47 24.9531
R1234 VN.n13 VN.n10 24.4675
R1235 VN.n17 VN.n10 24.4675
R1236 VN.n19 VN.n18 24.4675
R1237 VN.n19 VN.n8 24.4675
R1238 VN.n23 VN.n8 24.4675
R1239 VN.n24 VN.n23 24.4675
R1240 VN.n25 VN.n24 24.4675
R1241 VN.n25 VN.n6 24.4675
R1242 VN.n30 VN.n29 24.4675
R1243 VN.n31 VN.n30 24.4675
R1244 VN.n35 VN.n34 24.4675
R1245 VN.n36 VN.n35 24.4675
R1246 VN.n41 VN.n40 24.4675
R1247 VN.n42 VN.n41 24.4675
R1248 VN.n62 VN.n55 24.4675
R1249 VN.n58 VN.n55 24.4675
R1250 VN.n70 VN.n51 24.4675
R1251 VN.n70 VN.n69 24.4675
R1252 VN.n69 VN.n68 24.4675
R1253 VN.n68 VN.n53 24.4675
R1254 VN.n64 VN.n53 24.4675
R1255 VN.n64 VN.n63 24.4675
R1256 VN.n81 VN.n80 24.4675
R1257 VN.n80 VN.n79 24.4675
R1258 VN.n76 VN.n75 24.4675
R1259 VN.n75 VN.n74 24.4675
R1260 VN.n87 VN.n86 24.4675
R1261 VN.n86 VN.n85 24.4675
R1262 VN.n13 VN.n12 21.5315
R1263 VN.n31 VN.n4 21.5315
R1264 VN.n58 VN.n57 21.5315
R1265 VN.n76 VN.n49 21.5315
R1266 VN.n42 VN.n0 18.5954
R1267 VN.n87 VN.n45 18.5954
R1268 VN.n59 VN.n56 3.98138
R1269 VN.n14 VN.n11 3.98138
R1270 VN.n34 VN.n4 2.93654
R1271 VN.n79 VN.n49 2.93654
R1272 VN.n89 VN.n88 0.354971
R1273 VN.n44 VN.n43 0.354971
R1274 VN VN.n44 0.26696
R1275 VN.n88 VN.n46 0.189894
R1276 VN.n84 VN.n46 0.189894
R1277 VN.n84 VN.n83 0.189894
R1278 VN.n83 VN.n82 0.189894
R1279 VN.n82 VN.n48 0.189894
R1280 VN.n78 VN.n48 0.189894
R1281 VN.n78 VN.n77 0.189894
R1282 VN.n77 VN.n50 0.189894
R1283 VN.n73 VN.n50 0.189894
R1284 VN.n73 VN.n72 0.189894
R1285 VN.n72 VN.n71 0.189894
R1286 VN.n71 VN.n52 0.189894
R1287 VN.n67 VN.n52 0.189894
R1288 VN.n67 VN.n66 0.189894
R1289 VN.n66 VN.n65 0.189894
R1290 VN.n65 VN.n54 0.189894
R1291 VN.n61 VN.n54 0.189894
R1292 VN.n61 VN.n60 0.189894
R1293 VN.n60 VN.n59 0.189894
R1294 VN.n15 VN.n14 0.189894
R1295 VN.n16 VN.n15 0.189894
R1296 VN.n16 VN.n9 0.189894
R1297 VN.n20 VN.n9 0.189894
R1298 VN.n21 VN.n20 0.189894
R1299 VN.n22 VN.n21 0.189894
R1300 VN.n22 VN.n7 0.189894
R1301 VN.n26 VN.n7 0.189894
R1302 VN.n27 VN.n26 0.189894
R1303 VN.n28 VN.n27 0.189894
R1304 VN.n28 VN.n5 0.189894
R1305 VN.n32 VN.n5 0.189894
R1306 VN.n33 VN.n32 0.189894
R1307 VN.n33 VN.n3 0.189894
R1308 VN.n37 VN.n3 0.189894
R1309 VN.n38 VN.n37 0.189894
R1310 VN.n39 VN.n38 0.189894
R1311 VN.n39 VN.n1 0.189894
R1312 VN.n43 VN.n1 0.189894
R1313 VDD2.n210 VDD2.n209 585
R1314 VDD2.n208 VDD2.n207 585
R1315 VDD2.n113 VDD2.n112 585
R1316 VDD2.n202 VDD2.n201 585
R1317 VDD2.n200 VDD2.n199 585
R1318 VDD2.n117 VDD2.n116 585
R1319 VDD2.n194 VDD2.n193 585
R1320 VDD2.n192 VDD2.n191 585
R1321 VDD2.n121 VDD2.n120 585
R1322 VDD2.n186 VDD2.n185 585
R1323 VDD2.n184 VDD2.n183 585
R1324 VDD2.n125 VDD2.n124 585
R1325 VDD2.n178 VDD2.n177 585
R1326 VDD2.n176 VDD2.n175 585
R1327 VDD2.n129 VDD2.n128 585
R1328 VDD2.n170 VDD2.n169 585
R1329 VDD2.n168 VDD2.n167 585
R1330 VDD2.n166 VDD2.n132 585
R1331 VDD2.n136 VDD2.n133 585
R1332 VDD2.n161 VDD2.n160 585
R1333 VDD2.n159 VDD2.n158 585
R1334 VDD2.n138 VDD2.n137 585
R1335 VDD2.n153 VDD2.n152 585
R1336 VDD2.n151 VDD2.n150 585
R1337 VDD2.n142 VDD2.n141 585
R1338 VDD2.n145 VDD2.n144 585
R1339 VDD2.n35 VDD2.n34 585
R1340 VDD2.n32 VDD2.n31 585
R1341 VDD2.n41 VDD2.n40 585
R1342 VDD2.n43 VDD2.n42 585
R1343 VDD2.n28 VDD2.n27 585
R1344 VDD2.n49 VDD2.n48 585
R1345 VDD2.n52 VDD2.n51 585
R1346 VDD2.n50 VDD2.n24 585
R1347 VDD2.n57 VDD2.n23 585
R1348 VDD2.n59 VDD2.n58 585
R1349 VDD2.n61 VDD2.n60 585
R1350 VDD2.n20 VDD2.n19 585
R1351 VDD2.n67 VDD2.n66 585
R1352 VDD2.n69 VDD2.n68 585
R1353 VDD2.n16 VDD2.n15 585
R1354 VDD2.n75 VDD2.n74 585
R1355 VDD2.n77 VDD2.n76 585
R1356 VDD2.n12 VDD2.n11 585
R1357 VDD2.n83 VDD2.n82 585
R1358 VDD2.n85 VDD2.n84 585
R1359 VDD2.n8 VDD2.n7 585
R1360 VDD2.n91 VDD2.n90 585
R1361 VDD2.n93 VDD2.n92 585
R1362 VDD2.n4 VDD2.n3 585
R1363 VDD2.n99 VDD2.n98 585
R1364 VDD2.n101 VDD2.n100 585
R1365 VDD2.n209 VDD2.n109 498.474
R1366 VDD2.n100 VDD2.n0 498.474
R1367 VDD2.t6 VDD2.n143 329.036
R1368 VDD2.t9 VDD2.n33 329.036
R1369 VDD2.n209 VDD2.n208 171.744
R1370 VDD2.n208 VDD2.n112 171.744
R1371 VDD2.n201 VDD2.n112 171.744
R1372 VDD2.n201 VDD2.n200 171.744
R1373 VDD2.n200 VDD2.n116 171.744
R1374 VDD2.n193 VDD2.n116 171.744
R1375 VDD2.n193 VDD2.n192 171.744
R1376 VDD2.n192 VDD2.n120 171.744
R1377 VDD2.n185 VDD2.n120 171.744
R1378 VDD2.n185 VDD2.n184 171.744
R1379 VDD2.n184 VDD2.n124 171.744
R1380 VDD2.n177 VDD2.n124 171.744
R1381 VDD2.n177 VDD2.n176 171.744
R1382 VDD2.n176 VDD2.n128 171.744
R1383 VDD2.n169 VDD2.n128 171.744
R1384 VDD2.n169 VDD2.n168 171.744
R1385 VDD2.n168 VDD2.n132 171.744
R1386 VDD2.n136 VDD2.n132 171.744
R1387 VDD2.n160 VDD2.n136 171.744
R1388 VDD2.n160 VDD2.n159 171.744
R1389 VDD2.n159 VDD2.n137 171.744
R1390 VDD2.n152 VDD2.n137 171.744
R1391 VDD2.n152 VDD2.n151 171.744
R1392 VDD2.n151 VDD2.n141 171.744
R1393 VDD2.n144 VDD2.n141 171.744
R1394 VDD2.n34 VDD2.n31 171.744
R1395 VDD2.n41 VDD2.n31 171.744
R1396 VDD2.n42 VDD2.n41 171.744
R1397 VDD2.n42 VDD2.n27 171.744
R1398 VDD2.n49 VDD2.n27 171.744
R1399 VDD2.n51 VDD2.n49 171.744
R1400 VDD2.n51 VDD2.n50 171.744
R1401 VDD2.n50 VDD2.n23 171.744
R1402 VDD2.n59 VDD2.n23 171.744
R1403 VDD2.n60 VDD2.n59 171.744
R1404 VDD2.n60 VDD2.n19 171.744
R1405 VDD2.n67 VDD2.n19 171.744
R1406 VDD2.n68 VDD2.n67 171.744
R1407 VDD2.n68 VDD2.n15 171.744
R1408 VDD2.n75 VDD2.n15 171.744
R1409 VDD2.n76 VDD2.n75 171.744
R1410 VDD2.n76 VDD2.n11 171.744
R1411 VDD2.n83 VDD2.n11 171.744
R1412 VDD2.n84 VDD2.n83 171.744
R1413 VDD2.n84 VDD2.n7 171.744
R1414 VDD2.n91 VDD2.n7 171.744
R1415 VDD2.n92 VDD2.n91 171.744
R1416 VDD2.n92 VDD2.n3 171.744
R1417 VDD2.n99 VDD2.n3 171.744
R1418 VDD2.n100 VDD2.n99 171.744
R1419 VDD2.n144 VDD2.t6 85.8723
R1420 VDD2.n34 VDD2.t9 85.8723
R1421 VDD2.n108 VDD2.n107 71.7573
R1422 VDD2 VDD2.n217 71.7545
R1423 VDD2.n216 VDD2.n215 69.5887
R1424 VDD2.n106 VDD2.n105 69.5885
R1425 VDD2.n214 VDD2.n108 54.5343
R1426 VDD2.n106 VDD2.n104 53.5751
R1427 VDD2.n214 VDD2.n213 50.6096
R1428 VDD2.n167 VDD2.n166 13.1884
R1429 VDD2.n58 VDD2.n57 13.1884
R1430 VDD2.n211 VDD2.n210 12.8005
R1431 VDD2.n170 VDD2.n131 12.8005
R1432 VDD2.n165 VDD2.n133 12.8005
R1433 VDD2.n56 VDD2.n24 12.8005
R1434 VDD2.n61 VDD2.n22 12.8005
R1435 VDD2.n102 VDD2.n101 12.8005
R1436 VDD2.n207 VDD2.n111 12.0247
R1437 VDD2.n171 VDD2.n129 12.0247
R1438 VDD2.n162 VDD2.n161 12.0247
R1439 VDD2.n53 VDD2.n52 12.0247
R1440 VDD2.n62 VDD2.n20 12.0247
R1441 VDD2.n98 VDD2.n2 12.0247
R1442 VDD2.n206 VDD2.n113 11.249
R1443 VDD2.n175 VDD2.n174 11.249
R1444 VDD2.n158 VDD2.n135 11.249
R1445 VDD2.n48 VDD2.n26 11.249
R1446 VDD2.n66 VDD2.n65 11.249
R1447 VDD2.n97 VDD2.n4 11.249
R1448 VDD2.n145 VDD2.n143 10.7239
R1449 VDD2.n35 VDD2.n33 10.7239
R1450 VDD2.n203 VDD2.n202 10.4732
R1451 VDD2.n178 VDD2.n127 10.4732
R1452 VDD2.n157 VDD2.n138 10.4732
R1453 VDD2.n47 VDD2.n28 10.4732
R1454 VDD2.n69 VDD2.n18 10.4732
R1455 VDD2.n94 VDD2.n93 10.4732
R1456 VDD2.n199 VDD2.n115 9.69747
R1457 VDD2.n179 VDD2.n125 9.69747
R1458 VDD2.n154 VDD2.n153 9.69747
R1459 VDD2.n44 VDD2.n43 9.69747
R1460 VDD2.n70 VDD2.n16 9.69747
R1461 VDD2.n90 VDD2.n6 9.69747
R1462 VDD2.n213 VDD2.n212 9.45567
R1463 VDD2.n104 VDD2.n103 9.45567
R1464 VDD2.n147 VDD2.n146 9.3005
R1465 VDD2.n149 VDD2.n148 9.3005
R1466 VDD2.n140 VDD2.n139 9.3005
R1467 VDD2.n155 VDD2.n154 9.3005
R1468 VDD2.n157 VDD2.n156 9.3005
R1469 VDD2.n135 VDD2.n134 9.3005
R1470 VDD2.n163 VDD2.n162 9.3005
R1471 VDD2.n165 VDD2.n164 9.3005
R1472 VDD2.n119 VDD2.n118 9.3005
R1473 VDD2.n196 VDD2.n195 9.3005
R1474 VDD2.n198 VDD2.n197 9.3005
R1475 VDD2.n115 VDD2.n114 9.3005
R1476 VDD2.n204 VDD2.n203 9.3005
R1477 VDD2.n206 VDD2.n205 9.3005
R1478 VDD2.n111 VDD2.n110 9.3005
R1479 VDD2.n212 VDD2.n211 9.3005
R1480 VDD2.n190 VDD2.n189 9.3005
R1481 VDD2.n188 VDD2.n187 9.3005
R1482 VDD2.n123 VDD2.n122 9.3005
R1483 VDD2.n182 VDD2.n181 9.3005
R1484 VDD2.n180 VDD2.n179 9.3005
R1485 VDD2.n127 VDD2.n126 9.3005
R1486 VDD2.n174 VDD2.n173 9.3005
R1487 VDD2.n172 VDD2.n171 9.3005
R1488 VDD2.n131 VDD2.n130 9.3005
R1489 VDD2.n79 VDD2.n78 9.3005
R1490 VDD2.n14 VDD2.n13 9.3005
R1491 VDD2.n73 VDD2.n72 9.3005
R1492 VDD2.n71 VDD2.n70 9.3005
R1493 VDD2.n18 VDD2.n17 9.3005
R1494 VDD2.n65 VDD2.n64 9.3005
R1495 VDD2.n63 VDD2.n62 9.3005
R1496 VDD2.n22 VDD2.n21 9.3005
R1497 VDD2.n37 VDD2.n36 9.3005
R1498 VDD2.n39 VDD2.n38 9.3005
R1499 VDD2.n30 VDD2.n29 9.3005
R1500 VDD2.n45 VDD2.n44 9.3005
R1501 VDD2.n47 VDD2.n46 9.3005
R1502 VDD2.n26 VDD2.n25 9.3005
R1503 VDD2.n54 VDD2.n53 9.3005
R1504 VDD2.n56 VDD2.n55 9.3005
R1505 VDD2.n81 VDD2.n80 9.3005
R1506 VDD2.n10 VDD2.n9 9.3005
R1507 VDD2.n87 VDD2.n86 9.3005
R1508 VDD2.n89 VDD2.n88 9.3005
R1509 VDD2.n6 VDD2.n5 9.3005
R1510 VDD2.n95 VDD2.n94 9.3005
R1511 VDD2.n97 VDD2.n96 9.3005
R1512 VDD2.n2 VDD2.n1 9.3005
R1513 VDD2.n103 VDD2.n102 9.3005
R1514 VDD2.n198 VDD2.n117 8.92171
R1515 VDD2.n183 VDD2.n182 8.92171
R1516 VDD2.n150 VDD2.n140 8.92171
R1517 VDD2.n40 VDD2.n30 8.92171
R1518 VDD2.n74 VDD2.n73 8.92171
R1519 VDD2.n89 VDD2.n8 8.92171
R1520 VDD2.n195 VDD2.n194 8.14595
R1521 VDD2.n186 VDD2.n123 8.14595
R1522 VDD2.n149 VDD2.n142 8.14595
R1523 VDD2.n39 VDD2.n32 8.14595
R1524 VDD2.n77 VDD2.n14 8.14595
R1525 VDD2.n86 VDD2.n85 8.14595
R1526 VDD2.n213 VDD2.n109 7.75445
R1527 VDD2.n104 VDD2.n0 7.75445
R1528 VDD2.n191 VDD2.n119 7.3702
R1529 VDD2.n187 VDD2.n121 7.3702
R1530 VDD2.n146 VDD2.n145 7.3702
R1531 VDD2.n36 VDD2.n35 7.3702
R1532 VDD2.n78 VDD2.n12 7.3702
R1533 VDD2.n82 VDD2.n10 7.3702
R1534 VDD2.n191 VDD2.n190 6.59444
R1535 VDD2.n190 VDD2.n121 6.59444
R1536 VDD2.n81 VDD2.n12 6.59444
R1537 VDD2.n82 VDD2.n81 6.59444
R1538 VDD2.n211 VDD2.n109 6.08283
R1539 VDD2.n102 VDD2.n0 6.08283
R1540 VDD2.n194 VDD2.n119 5.81868
R1541 VDD2.n187 VDD2.n186 5.81868
R1542 VDD2.n146 VDD2.n142 5.81868
R1543 VDD2.n36 VDD2.n32 5.81868
R1544 VDD2.n78 VDD2.n77 5.81868
R1545 VDD2.n85 VDD2.n10 5.81868
R1546 VDD2.n195 VDD2.n117 5.04292
R1547 VDD2.n183 VDD2.n123 5.04292
R1548 VDD2.n150 VDD2.n149 5.04292
R1549 VDD2.n40 VDD2.n39 5.04292
R1550 VDD2.n74 VDD2.n14 5.04292
R1551 VDD2.n86 VDD2.n8 5.04292
R1552 VDD2.n199 VDD2.n198 4.26717
R1553 VDD2.n182 VDD2.n125 4.26717
R1554 VDD2.n153 VDD2.n140 4.26717
R1555 VDD2.n43 VDD2.n30 4.26717
R1556 VDD2.n73 VDD2.n16 4.26717
R1557 VDD2.n90 VDD2.n89 4.26717
R1558 VDD2.n202 VDD2.n115 3.49141
R1559 VDD2.n179 VDD2.n178 3.49141
R1560 VDD2.n154 VDD2.n138 3.49141
R1561 VDD2.n44 VDD2.n28 3.49141
R1562 VDD2.n70 VDD2.n69 3.49141
R1563 VDD2.n93 VDD2.n6 3.49141
R1564 VDD2.n216 VDD2.n214 2.96602
R1565 VDD2.n203 VDD2.n113 2.71565
R1566 VDD2.n175 VDD2.n127 2.71565
R1567 VDD2.n158 VDD2.n157 2.71565
R1568 VDD2.n48 VDD2.n47 2.71565
R1569 VDD2.n66 VDD2.n18 2.71565
R1570 VDD2.n94 VDD2.n4 2.71565
R1571 VDD2.n147 VDD2.n143 2.41282
R1572 VDD2.n37 VDD2.n33 2.41282
R1573 VDD2.n207 VDD2.n206 1.93989
R1574 VDD2.n174 VDD2.n129 1.93989
R1575 VDD2.n161 VDD2.n135 1.93989
R1576 VDD2.n52 VDD2.n26 1.93989
R1577 VDD2.n65 VDD2.n20 1.93989
R1578 VDD2.n98 VDD2.n97 1.93989
R1579 VDD2.n217 VDD2.t7 1.67515
R1580 VDD2.n217 VDD2.t4 1.67515
R1581 VDD2.n215 VDD2.t2 1.67515
R1582 VDD2.n215 VDD2.t8 1.67515
R1583 VDD2.n107 VDD2.t1 1.67515
R1584 VDD2.n107 VDD2.t0 1.67515
R1585 VDD2.n105 VDD2.t5 1.67515
R1586 VDD2.n105 VDD2.t3 1.67515
R1587 VDD2.n210 VDD2.n111 1.16414
R1588 VDD2.n171 VDD2.n170 1.16414
R1589 VDD2.n162 VDD2.n133 1.16414
R1590 VDD2.n53 VDD2.n24 1.16414
R1591 VDD2.n62 VDD2.n61 1.16414
R1592 VDD2.n101 VDD2.n2 1.16414
R1593 VDD2 VDD2.n216 0.800069
R1594 VDD2.n108 VDD2.n106 0.686533
R1595 VDD2.n167 VDD2.n131 0.388379
R1596 VDD2.n166 VDD2.n165 0.388379
R1597 VDD2.n57 VDD2.n56 0.388379
R1598 VDD2.n58 VDD2.n22 0.388379
R1599 VDD2.n212 VDD2.n110 0.155672
R1600 VDD2.n205 VDD2.n110 0.155672
R1601 VDD2.n205 VDD2.n204 0.155672
R1602 VDD2.n204 VDD2.n114 0.155672
R1603 VDD2.n197 VDD2.n114 0.155672
R1604 VDD2.n197 VDD2.n196 0.155672
R1605 VDD2.n196 VDD2.n118 0.155672
R1606 VDD2.n189 VDD2.n118 0.155672
R1607 VDD2.n189 VDD2.n188 0.155672
R1608 VDD2.n188 VDD2.n122 0.155672
R1609 VDD2.n181 VDD2.n122 0.155672
R1610 VDD2.n181 VDD2.n180 0.155672
R1611 VDD2.n180 VDD2.n126 0.155672
R1612 VDD2.n173 VDD2.n126 0.155672
R1613 VDD2.n173 VDD2.n172 0.155672
R1614 VDD2.n172 VDD2.n130 0.155672
R1615 VDD2.n164 VDD2.n130 0.155672
R1616 VDD2.n164 VDD2.n163 0.155672
R1617 VDD2.n163 VDD2.n134 0.155672
R1618 VDD2.n156 VDD2.n134 0.155672
R1619 VDD2.n156 VDD2.n155 0.155672
R1620 VDD2.n155 VDD2.n139 0.155672
R1621 VDD2.n148 VDD2.n139 0.155672
R1622 VDD2.n148 VDD2.n147 0.155672
R1623 VDD2.n38 VDD2.n37 0.155672
R1624 VDD2.n38 VDD2.n29 0.155672
R1625 VDD2.n45 VDD2.n29 0.155672
R1626 VDD2.n46 VDD2.n45 0.155672
R1627 VDD2.n46 VDD2.n25 0.155672
R1628 VDD2.n54 VDD2.n25 0.155672
R1629 VDD2.n55 VDD2.n54 0.155672
R1630 VDD2.n55 VDD2.n21 0.155672
R1631 VDD2.n63 VDD2.n21 0.155672
R1632 VDD2.n64 VDD2.n63 0.155672
R1633 VDD2.n64 VDD2.n17 0.155672
R1634 VDD2.n71 VDD2.n17 0.155672
R1635 VDD2.n72 VDD2.n71 0.155672
R1636 VDD2.n72 VDD2.n13 0.155672
R1637 VDD2.n79 VDD2.n13 0.155672
R1638 VDD2.n80 VDD2.n79 0.155672
R1639 VDD2.n80 VDD2.n9 0.155672
R1640 VDD2.n87 VDD2.n9 0.155672
R1641 VDD2.n88 VDD2.n87 0.155672
R1642 VDD2.n88 VDD2.n5 0.155672
R1643 VDD2.n95 VDD2.n5 0.155672
R1644 VDD2.n96 VDD2.n95 0.155672
R1645 VDD2.n96 VDD2.n1 0.155672
R1646 VDD2.n103 VDD2.n1 0.155672
R1647 B.n802 B.n801 585
R1648 B.n803 B.n108 585
R1649 B.n805 B.n804 585
R1650 B.n806 B.n107 585
R1651 B.n808 B.n807 585
R1652 B.n809 B.n106 585
R1653 B.n811 B.n810 585
R1654 B.n812 B.n105 585
R1655 B.n814 B.n813 585
R1656 B.n815 B.n104 585
R1657 B.n817 B.n816 585
R1658 B.n818 B.n103 585
R1659 B.n820 B.n819 585
R1660 B.n821 B.n102 585
R1661 B.n823 B.n822 585
R1662 B.n824 B.n101 585
R1663 B.n826 B.n825 585
R1664 B.n827 B.n100 585
R1665 B.n829 B.n828 585
R1666 B.n830 B.n99 585
R1667 B.n832 B.n831 585
R1668 B.n833 B.n98 585
R1669 B.n835 B.n834 585
R1670 B.n836 B.n97 585
R1671 B.n838 B.n837 585
R1672 B.n839 B.n96 585
R1673 B.n841 B.n840 585
R1674 B.n842 B.n95 585
R1675 B.n844 B.n843 585
R1676 B.n845 B.n94 585
R1677 B.n847 B.n846 585
R1678 B.n848 B.n93 585
R1679 B.n850 B.n849 585
R1680 B.n851 B.n92 585
R1681 B.n853 B.n852 585
R1682 B.n854 B.n91 585
R1683 B.n856 B.n855 585
R1684 B.n857 B.n90 585
R1685 B.n859 B.n858 585
R1686 B.n860 B.n89 585
R1687 B.n862 B.n861 585
R1688 B.n863 B.n88 585
R1689 B.n865 B.n864 585
R1690 B.n866 B.n87 585
R1691 B.n868 B.n867 585
R1692 B.n869 B.n86 585
R1693 B.n871 B.n870 585
R1694 B.n872 B.n85 585
R1695 B.n874 B.n873 585
R1696 B.n875 B.n84 585
R1697 B.n877 B.n876 585
R1698 B.n878 B.n83 585
R1699 B.n880 B.n879 585
R1700 B.n881 B.n82 585
R1701 B.n883 B.n882 585
R1702 B.n884 B.n81 585
R1703 B.n886 B.n885 585
R1704 B.n887 B.n80 585
R1705 B.n889 B.n888 585
R1706 B.n890 B.n79 585
R1707 B.n892 B.n891 585
R1708 B.n893 B.n78 585
R1709 B.n895 B.n894 585
R1710 B.n897 B.n75 585
R1711 B.n899 B.n898 585
R1712 B.n900 B.n74 585
R1713 B.n902 B.n901 585
R1714 B.n903 B.n73 585
R1715 B.n905 B.n904 585
R1716 B.n906 B.n72 585
R1717 B.n908 B.n907 585
R1718 B.n909 B.n71 585
R1719 B.n911 B.n910 585
R1720 B.n913 B.n912 585
R1721 B.n914 B.n67 585
R1722 B.n916 B.n915 585
R1723 B.n917 B.n66 585
R1724 B.n919 B.n918 585
R1725 B.n920 B.n65 585
R1726 B.n922 B.n921 585
R1727 B.n923 B.n64 585
R1728 B.n925 B.n924 585
R1729 B.n926 B.n63 585
R1730 B.n928 B.n927 585
R1731 B.n929 B.n62 585
R1732 B.n931 B.n930 585
R1733 B.n932 B.n61 585
R1734 B.n934 B.n933 585
R1735 B.n935 B.n60 585
R1736 B.n937 B.n936 585
R1737 B.n938 B.n59 585
R1738 B.n940 B.n939 585
R1739 B.n941 B.n58 585
R1740 B.n943 B.n942 585
R1741 B.n944 B.n57 585
R1742 B.n946 B.n945 585
R1743 B.n947 B.n56 585
R1744 B.n949 B.n948 585
R1745 B.n950 B.n55 585
R1746 B.n952 B.n951 585
R1747 B.n953 B.n54 585
R1748 B.n955 B.n954 585
R1749 B.n956 B.n53 585
R1750 B.n958 B.n957 585
R1751 B.n959 B.n52 585
R1752 B.n961 B.n960 585
R1753 B.n962 B.n51 585
R1754 B.n964 B.n963 585
R1755 B.n965 B.n50 585
R1756 B.n967 B.n966 585
R1757 B.n968 B.n49 585
R1758 B.n970 B.n969 585
R1759 B.n971 B.n48 585
R1760 B.n973 B.n972 585
R1761 B.n974 B.n47 585
R1762 B.n976 B.n975 585
R1763 B.n977 B.n46 585
R1764 B.n979 B.n978 585
R1765 B.n980 B.n45 585
R1766 B.n982 B.n981 585
R1767 B.n983 B.n44 585
R1768 B.n985 B.n984 585
R1769 B.n986 B.n43 585
R1770 B.n988 B.n987 585
R1771 B.n989 B.n42 585
R1772 B.n991 B.n990 585
R1773 B.n992 B.n41 585
R1774 B.n994 B.n993 585
R1775 B.n995 B.n40 585
R1776 B.n997 B.n996 585
R1777 B.n998 B.n39 585
R1778 B.n1000 B.n999 585
R1779 B.n1001 B.n38 585
R1780 B.n1003 B.n1002 585
R1781 B.n1004 B.n37 585
R1782 B.n1006 B.n1005 585
R1783 B.n800 B.n109 585
R1784 B.n799 B.n798 585
R1785 B.n797 B.n110 585
R1786 B.n796 B.n795 585
R1787 B.n794 B.n111 585
R1788 B.n793 B.n792 585
R1789 B.n791 B.n112 585
R1790 B.n790 B.n789 585
R1791 B.n788 B.n113 585
R1792 B.n787 B.n786 585
R1793 B.n785 B.n114 585
R1794 B.n784 B.n783 585
R1795 B.n782 B.n115 585
R1796 B.n781 B.n780 585
R1797 B.n779 B.n116 585
R1798 B.n778 B.n777 585
R1799 B.n776 B.n117 585
R1800 B.n775 B.n774 585
R1801 B.n773 B.n118 585
R1802 B.n772 B.n771 585
R1803 B.n770 B.n119 585
R1804 B.n769 B.n768 585
R1805 B.n767 B.n120 585
R1806 B.n766 B.n765 585
R1807 B.n764 B.n121 585
R1808 B.n763 B.n762 585
R1809 B.n761 B.n122 585
R1810 B.n760 B.n759 585
R1811 B.n758 B.n123 585
R1812 B.n757 B.n756 585
R1813 B.n755 B.n124 585
R1814 B.n754 B.n753 585
R1815 B.n752 B.n125 585
R1816 B.n751 B.n750 585
R1817 B.n749 B.n126 585
R1818 B.n748 B.n747 585
R1819 B.n746 B.n127 585
R1820 B.n745 B.n744 585
R1821 B.n743 B.n128 585
R1822 B.n742 B.n741 585
R1823 B.n740 B.n129 585
R1824 B.n739 B.n738 585
R1825 B.n737 B.n130 585
R1826 B.n736 B.n735 585
R1827 B.n734 B.n131 585
R1828 B.n733 B.n732 585
R1829 B.n731 B.n132 585
R1830 B.n730 B.n729 585
R1831 B.n728 B.n133 585
R1832 B.n727 B.n726 585
R1833 B.n725 B.n134 585
R1834 B.n724 B.n723 585
R1835 B.n722 B.n135 585
R1836 B.n721 B.n720 585
R1837 B.n719 B.n136 585
R1838 B.n718 B.n717 585
R1839 B.n716 B.n137 585
R1840 B.n715 B.n714 585
R1841 B.n713 B.n138 585
R1842 B.n712 B.n711 585
R1843 B.n710 B.n139 585
R1844 B.n709 B.n708 585
R1845 B.n707 B.n140 585
R1846 B.n706 B.n705 585
R1847 B.n704 B.n141 585
R1848 B.n703 B.n702 585
R1849 B.n701 B.n142 585
R1850 B.n700 B.n699 585
R1851 B.n698 B.n143 585
R1852 B.n697 B.n696 585
R1853 B.n695 B.n144 585
R1854 B.n694 B.n693 585
R1855 B.n692 B.n145 585
R1856 B.n691 B.n690 585
R1857 B.n689 B.n146 585
R1858 B.n688 B.n687 585
R1859 B.n686 B.n147 585
R1860 B.n685 B.n684 585
R1861 B.n683 B.n148 585
R1862 B.n682 B.n681 585
R1863 B.n680 B.n149 585
R1864 B.n679 B.n678 585
R1865 B.n677 B.n150 585
R1866 B.n676 B.n675 585
R1867 B.n674 B.n151 585
R1868 B.n673 B.n672 585
R1869 B.n671 B.n152 585
R1870 B.n670 B.n669 585
R1871 B.n668 B.n153 585
R1872 B.n667 B.n666 585
R1873 B.n665 B.n154 585
R1874 B.n664 B.n663 585
R1875 B.n662 B.n155 585
R1876 B.n661 B.n660 585
R1877 B.n659 B.n156 585
R1878 B.n658 B.n657 585
R1879 B.n656 B.n157 585
R1880 B.n655 B.n654 585
R1881 B.n653 B.n158 585
R1882 B.n652 B.n651 585
R1883 B.n650 B.n159 585
R1884 B.n649 B.n648 585
R1885 B.n647 B.n160 585
R1886 B.n646 B.n645 585
R1887 B.n644 B.n161 585
R1888 B.n643 B.n642 585
R1889 B.n641 B.n162 585
R1890 B.n640 B.n639 585
R1891 B.n638 B.n163 585
R1892 B.n637 B.n636 585
R1893 B.n635 B.n164 585
R1894 B.n634 B.n633 585
R1895 B.n632 B.n165 585
R1896 B.n631 B.n630 585
R1897 B.n629 B.n166 585
R1898 B.n628 B.n627 585
R1899 B.n626 B.n167 585
R1900 B.n625 B.n624 585
R1901 B.n623 B.n168 585
R1902 B.n622 B.n621 585
R1903 B.n620 B.n169 585
R1904 B.n619 B.n618 585
R1905 B.n617 B.n170 585
R1906 B.n616 B.n615 585
R1907 B.n614 B.n171 585
R1908 B.n613 B.n612 585
R1909 B.n611 B.n172 585
R1910 B.n610 B.n609 585
R1911 B.n608 B.n173 585
R1912 B.n607 B.n606 585
R1913 B.n605 B.n174 585
R1914 B.n604 B.n603 585
R1915 B.n602 B.n175 585
R1916 B.n601 B.n600 585
R1917 B.n599 B.n176 585
R1918 B.n598 B.n597 585
R1919 B.n596 B.n177 585
R1920 B.n595 B.n594 585
R1921 B.n593 B.n178 585
R1922 B.n388 B.n387 585
R1923 B.n389 B.n250 585
R1924 B.n391 B.n390 585
R1925 B.n392 B.n249 585
R1926 B.n394 B.n393 585
R1927 B.n395 B.n248 585
R1928 B.n397 B.n396 585
R1929 B.n398 B.n247 585
R1930 B.n400 B.n399 585
R1931 B.n401 B.n246 585
R1932 B.n403 B.n402 585
R1933 B.n404 B.n245 585
R1934 B.n406 B.n405 585
R1935 B.n407 B.n244 585
R1936 B.n409 B.n408 585
R1937 B.n410 B.n243 585
R1938 B.n412 B.n411 585
R1939 B.n413 B.n242 585
R1940 B.n415 B.n414 585
R1941 B.n416 B.n241 585
R1942 B.n418 B.n417 585
R1943 B.n419 B.n240 585
R1944 B.n421 B.n420 585
R1945 B.n422 B.n239 585
R1946 B.n424 B.n423 585
R1947 B.n425 B.n238 585
R1948 B.n427 B.n426 585
R1949 B.n428 B.n237 585
R1950 B.n430 B.n429 585
R1951 B.n431 B.n236 585
R1952 B.n433 B.n432 585
R1953 B.n434 B.n235 585
R1954 B.n436 B.n435 585
R1955 B.n437 B.n234 585
R1956 B.n439 B.n438 585
R1957 B.n440 B.n233 585
R1958 B.n442 B.n441 585
R1959 B.n443 B.n232 585
R1960 B.n445 B.n444 585
R1961 B.n446 B.n231 585
R1962 B.n448 B.n447 585
R1963 B.n449 B.n230 585
R1964 B.n451 B.n450 585
R1965 B.n452 B.n229 585
R1966 B.n454 B.n453 585
R1967 B.n455 B.n228 585
R1968 B.n457 B.n456 585
R1969 B.n458 B.n227 585
R1970 B.n460 B.n459 585
R1971 B.n461 B.n226 585
R1972 B.n463 B.n462 585
R1973 B.n464 B.n225 585
R1974 B.n466 B.n465 585
R1975 B.n467 B.n224 585
R1976 B.n469 B.n468 585
R1977 B.n470 B.n223 585
R1978 B.n472 B.n471 585
R1979 B.n473 B.n222 585
R1980 B.n475 B.n474 585
R1981 B.n476 B.n221 585
R1982 B.n478 B.n477 585
R1983 B.n479 B.n220 585
R1984 B.n481 B.n480 585
R1985 B.n483 B.n217 585
R1986 B.n485 B.n484 585
R1987 B.n486 B.n216 585
R1988 B.n488 B.n487 585
R1989 B.n489 B.n215 585
R1990 B.n491 B.n490 585
R1991 B.n492 B.n214 585
R1992 B.n494 B.n493 585
R1993 B.n495 B.n213 585
R1994 B.n497 B.n496 585
R1995 B.n499 B.n498 585
R1996 B.n500 B.n209 585
R1997 B.n502 B.n501 585
R1998 B.n503 B.n208 585
R1999 B.n505 B.n504 585
R2000 B.n506 B.n207 585
R2001 B.n508 B.n507 585
R2002 B.n509 B.n206 585
R2003 B.n511 B.n510 585
R2004 B.n512 B.n205 585
R2005 B.n514 B.n513 585
R2006 B.n515 B.n204 585
R2007 B.n517 B.n516 585
R2008 B.n518 B.n203 585
R2009 B.n520 B.n519 585
R2010 B.n521 B.n202 585
R2011 B.n523 B.n522 585
R2012 B.n524 B.n201 585
R2013 B.n526 B.n525 585
R2014 B.n527 B.n200 585
R2015 B.n529 B.n528 585
R2016 B.n530 B.n199 585
R2017 B.n532 B.n531 585
R2018 B.n533 B.n198 585
R2019 B.n535 B.n534 585
R2020 B.n536 B.n197 585
R2021 B.n538 B.n537 585
R2022 B.n539 B.n196 585
R2023 B.n541 B.n540 585
R2024 B.n542 B.n195 585
R2025 B.n544 B.n543 585
R2026 B.n545 B.n194 585
R2027 B.n547 B.n546 585
R2028 B.n548 B.n193 585
R2029 B.n550 B.n549 585
R2030 B.n551 B.n192 585
R2031 B.n553 B.n552 585
R2032 B.n554 B.n191 585
R2033 B.n556 B.n555 585
R2034 B.n557 B.n190 585
R2035 B.n559 B.n558 585
R2036 B.n560 B.n189 585
R2037 B.n562 B.n561 585
R2038 B.n563 B.n188 585
R2039 B.n565 B.n564 585
R2040 B.n566 B.n187 585
R2041 B.n568 B.n567 585
R2042 B.n569 B.n186 585
R2043 B.n571 B.n570 585
R2044 B.n572 B.n185 585
R2045 B.n574 B.n573 585
R2046 B.n575 B.n184 585
R2047 B.n577 B.n576 585
R2048 B.n578 B.n183 585
R2049 B.n580 B.n579 585
R2050 B.n581 B.n182 585
R2051 B.n583 B.n582 585
R2052 B.n584 B.n181 585
R2053 B.n586 B.n585 585
R2054 B.n587 B.n180 585
R2055 B.n589 B.n588 585
R2056 B.n590 B.n179 585
R2057 B.n592 B.n591 585
R2058 B.n386 B.n251 585
R2059 B.n385 B.n384 585
R2060 B.n383 B.n252 585
R2061 B.n382 B.n381 585
R2062 B.n380 B.n253 585
R2063 B.n379 B.n378 585
R2064 B.n377 B.n254 585
R2065 B.n376 B.n375 585
R2066 B.n374 B.n255 585
R2067 B.n373 B.n372 585
R2068 B.n371 B.n256 585
R2069 B.n370 B.n369 585
R2070 B.n368 B.n257 585
R2071 B.n367 B.n366 585
R2072 B.n365 B.n258 585
R2073 B.n364 B.n363 585
R2074 B.n362 B.n259 585
R2075 B.n361 B.n360 585
R2076 B.n359 B.n260 585
R2077 B.n358 B.n357 585
R2078 B.n356 B.n261 585
R2079 B.n355 B.n354 585
R2080 B.n353 B.n262 585
R2081 B.n352 B.n351 585
R2082 B.n350 B.n263 585
R2083 B.n349 B.n348 585
R2084 B.n347 B.n264 585
R2085 B.n346 B.n345 585
R2086 B.n344 B.n265 585
R2087 B.n343 B.n342 585
R2088 B.n341 B.n266 585
R2089 B.n340 B.n339 585
R2090 B.n338 B.n267 585
R2091 B.n337 B.n336 585
R2092 B.n335 B.n268 585
R2093 B.n334 B.n333 585
R2094 B.n332 B.n269 585
R2095 B.n331 B.n330 585
R2096 B.n329 B.n270 585
R2097 B.n328 B.n327 585
R2098 B.n326 B.n271 585
R2099 B.n325 B.n324 585
R2100 B.n323 B.n272 585
R2101 B.n322 B.n321 585
R2102 B.n320 B.n273 585
R2103 B.n319 B.n318 585
R2104 B.n317 B.n274 585
R2105 B.n316 B.n315 585
R2106 B.n314 B.n275 585
R2107 B.n313 B.n312 585
R2108 B.n311 B.n276 585
R2109 B.n310 B.n309 585
R2110 B.n308 B.n277 585
R2111 B.n307 B.n306 585
R2112 B.n305 B.n278 585
R2113 B.n304 B.n303 585
R2114 B.n302 B.n279 585
R2115 B.n301 B.n300 585
R2116 B.n299 B.n280 585
R2117 B.n298 B.n297 585
R2118 B.n296 B.n281 585
R2119 B.n295 B.n294 585
R2120 B.n293 B.n282 585
R2121 B.n292 B.n291 585
R2122 B.n290 B.n283 585
R2123 B.n289 B.n288 585
R2124 B.n287 B.n284 585
R2125 B.n286 B.n285 585
R2126 B.n2 B.n0 585
R2127 B.n1109 B.n1 585
R2128 B.n1108 B.n1107 585
R2129 B.n1106 B.n3 585
R2130 B.n1105 B.n1104 585
R2131 B.n1103 B.n4 585
R2132 B.n1102 B.n1101 585
R2133 B.n1100 B.n5 585
R2134 B.n1099 B.n1098 585
R2135 B.n1097 B.n6 585
R2136 B.n1096 B.n1095 585
R2137 B.n1094 B.n7 585
R2138 B.n1093 B.n1092 585
R2139 B.n1091 B.n8 585
R2140 B.n1090 B.n1089 585
R2141 B.n1088 B.n9 585
R2142 B.n1087 B.n1086 585
R2143 B.n1085 B.n10 585
R2144 B.n1084 B.n1083 585
R2145 B.n1082 B.n11 585
R2146 B.n1081 B.n1080 585
R2147 B.n1079 B.n12 585
R2148 B.n1078 B.n1077 585
R2149 B.n1076 B.n13 585
R2150 B.n1075 B.n1074 585
R2151 B.n1073 B.n14 585
R2152 B.n1072 B.n1071 585
R2153 B.n1070 B.n15 585
R2154 B.n1069 B.n1068 585
R2155 B.n1067 B.n16 585
R2156 B.n1066 B.n1065 585
R2157 B.n1064 B.n17 585
R2158 B.n1063 B.n1062 585
R2159 B.n1061 B.n18 585
R2160 B.n1060 B.n1059 585
R2161 B.n1058 B.n19 585
R2162 B.n1057 B.n1056 585
R2163 B.n1055 B.n20 585
R2164 B.n1054 B.n1053 585
R2165 B.n1052 B.n21 585
R2166 B.n1051 B.n1050 585
R2167 B.n1049 B.n22 585
R2168 B.n1048 B.n1047 585
R2169 B.n1046 B.n23 585
R2170 B.n1045 B.n1044 585
R2171 B.n1043 B.n24 585
R2172 B.n1042 B.n1041 585
R2173 B.n1040 B.n25 585
R2174 B.n1039 B.n1038 585
R2175 B.n1037 B.n26 585
R2176 B.n1036 B.n1035 585
R2177 B.n1034 B.n27 585
R2178 B.n1033 B.n1032 585
R2179 B.n1031 B.n28 585
R2180 B.n1030 B.n1029 585
R2181 B.n1028 B.n29 585
R2182 B.n1027 B.n1026 585
R2183 B.n1025 B.n30 585
R2184 B.n1024 B.n1023 585
R2185 B.n1022 B.n31 585
R2186 B.n1021 B.n1020 585
R2187 B.n1019 B.n32 585
R2188 B.n1018 B.n1017 585
R2189 B.n1016 B.n33 585
R2190 B.n1015 B.n1014 585
R2191 B.n1013 B.n34 585
R2192 B.n1012 B.n1011 585
R2193 B.n1010 B.n35 585
R2194 B.n1009 B.n1008 585
R2195 B.n1007 B.n36 585
R2196 B.n1111 B.n1110 585
R2197 B.n210 B.t8 575.615
R2198 B.n76 B.t1 575.615
R2199 B.n218 B.t5 575.615
R2200 B.n68 B.t10 575.615
R2201 B.n211 B.t7 508.901
R2202 B.n77 B.t2 508.901
R2203 B.n219 B.t4 508.901
R2204 B.n69 B.t11 508.901
R2205 B.n388 B.n251 502.111
R2206 B.n1007 B.n1006 502.111
R2207 B.n593 B.n592 502.111
R2208 B.n802 B.n109 502.111
R2209 B.n210 B.t6 359.118
R2210 B.n218 B.t3 359.118
R2211 B.n68 B.t9 359.118
R2212 B.n76 B.t0 359.118
R2213 B.n384 B.n251 163.367
R2214 B.n384 B.n383 163.367
R2215 B.n383 B.n382 163.367
R2216 B.n382 B.n253 163.367
R2217 B.n378 B.n253 163.367
R2218 B.n378 B.n377 163.367
R2219 B.n377 B.n376 163.367
R2220 B.n376 B.n255 163.367
R2221 B.n372 B.n255 163.367
R2222 B.n372 B.n371 163.367
R2223 B.n371 B.n370 163.367
R2224 B.n370 B.n257 163.367
R2225 B.n366 B.n257 163.367
R2226 B.n366 B.n365 163.367
R2227 B.n365 B.n364 163.367
R2228 B.n364 B.n259 163.367
R2229 B.n360 B.n259 163.367
R2230 B.n360 B.n359 163.367
R2231 B.n359 B.n358 163.367
R2232 B.n358 B.n261 163.367
R2233 B.n354 B.n261 163.367
R2234 B.n354 B.n353 163.367
R2235 B.n353 B.n352 163.367
R2236 B.n352 B.n263 163.367
R2237 B.n348 B.n263 163.367
R2238 B.n348 B.n347 163.367
R2239 B.n347 B.n346 163.367
R2240 B.n346 B.n265 163.367
R2241 B.n342 B.n265 163.367
R2242 B.n342 B.n341 163.367
R2243 B.n341 B.n340 163.367
R2244 B.n340 B.n267 163.367
R2245 B.n336 B.n267 163.367
R2246 B.n336 B.n335 163.367
R2247 B.n335 B.n334 163.367
R2248 B.n334 B.n269 163.367
R2249 B.n330 B.n269 163.367
R2250 B.n330 B.n329 163.367
R2251 B.n329 B.n328 163.367
R2252 B.n328 B.n271 163.367
R2253 B.n324 B.n271 163.367
R2254 B.n324 B.n323 163.367
R2255 B.n323 B.n322 163.367
R2256 B.n322 B.n273 163.367
R2257 B.n318 B.n273 163.367
R2258 B.n318 B.n317 163.367
R2259 B.n317 B.n316 163.367
R2260 B.n316 B.n275 163.367
R2261 B.n312 B.n275 163.367
R2262 B.n312 B.n311 163.367
R2263 B.n311 B.n310 163.367
R2264 B.n310 B.n277 163.367
R2265 B.n306 B.n277 163.367
R2266 B.n306 B.n305 163.367
R2267 B.n305 B.n304 163.367
R2268 B.n304 B.n279 163.367
R2269 B.n300 B.n279 163.367
R2270 B.n300 B.n299 163.367
R2271 B.n299 B.n298 163.367
R2272 B.n298 B.n281 163.367
R2273 B.n294 B.n281 163.367
R2274 B.n294 B.n293 163.367
R2275 B.n293 B.n292 163.367
R2276 B.n292 B.n283 163.367
R2277 B.n288 B.n283 163.367
R2278 B.n288 B.n287 163.367
R2279 B.n287 B.n286 163.367
R2280 B.n286 B.n2 163.367
R2281 B.n1110 B.n2 163.367
R2282 B.n1110 B.n1109 163.367
R2283 B.n1109 B.n1108 163.367
R2284 B.n1108 B.n3 163.367
R2285 B.n1104 B.n3 163.367
R2286 B.n1104 B.n1103 163.367
R2287 B.n1103 B.n1102 163.367
R2288 B.n1102 B.n5 163.367
R2289 B.n1098 B.n5 163.367
R2290 B.n1098 B.n1097 163.367
R2291 B.n1097 B.n1096 163.367
R2292 B.n1096 B.n7 163.367
R2293 B.n1092 B.n7 163.367
R2294 B.n1092 B.n1091 163.367
R2295 B.n1091 B.n1090 163.367
R2296 B.n1090 B.n9 163.367
R2297 B.n1086 B.n9 163.367
R2298 B.n1086 B.n1085 163.367
R2299 B.n1085 B.n1084 163.367
R2300 B.n1084 B.n11 163.367
R2301 B.n1080 B.n11 163.367
R2302 B.n1080 B.n1079 163.367
R2303 B.n1079 B.n1078 163.367
R2304 B.n1078 B.n13 163.367
R2305 B.n1074 B.n13 163.367
R2306 B.n1074 B.n1073 163.367
R2307 B.n1073 B.n1072 163.367
R2308 B.n1072 B.n15 163.367
R2309 B.n1068 B.n15 163.367
R2310 B.n1068 B.n1067 163.367
R2311 B.n1067 B.n1066 163.367
R2312 B.n1066 B.n17 163.367
R2313 B.n1062 B.n17 163.367
R2314 B.n1062 B.n1061 163.367
R2315 B.n1061 B.n1060 163.367
R2316 B.n1060 B.n19 163.367
R2317 B.n1056 B.n19 163.367
R2318 B.n1056 B.n1055 163.367
R2319 B.n1055 B.n1054 163.367
R2320 B.n1054 B.n21 163.367
R2321 B.n1050 B.n21 163.367
R2322 B.n1050 B.n1049 163.367
R2323 B.n1049 B.n1048 163.367
R2324 B.n1048 B.n23 163.367
R2325 B.n1044 B.n23 163.367
R2326 B.n1044 B.n1043 163.367
R2327 B.n1043 B.n1042 163.367
R2328 B.n1042 B.n25 163.367
R2329 B.n1038 B.n25 163.367
R2330 B.n1038 B.n1037 163.367
R2331 B.n1037 B.n1036 163.367
R2332 B.n1036 B.n27 163.367
R2333 B.n1032 B.n27 163.367
R2334 B.n1032 B.n1031 163.367
R2335 B.n1031 B.n1030 163.367
R2336 B.n1030 B.n29 163.367
R2337 B.n1026 B.n29 163.367
R2338 B.n1026 B.n1025 163.367
R2339 B.n1025 B.n1024 163.367
R2340 B.n1024 B.n31 163.367
R2341 B.n1020 B.n31 163.367
R2342 B.n1020 B.n1019 163.367
R2343 B.n1019 B.n1018 163.367
R2344 B.n1018 B.n33 163.367
R2345 B.n1014 B.n33 163.367
R2346 B.n1014 B.n1013 163.367
R2347 B.n1013 B.n1012 163.367
R2348 B.n1012 B.n35 163.367
R2349 B.n1008 B.n35 163.367
R2350 B.n1008 B.n1007 163.367
R2351 B.n389 B.n388 163.367
R2352 B.n390 B.n389 163.367
R2353 B.n390 B.n249 163.367
R2354 B.n394 B.n249 163.367
R2355 B.n395 B.n394 163.367
R2356 B.n396 B.n395 163.367
R2357 B.n396 B.n247 163.367
R2358 B.n400 B.n247 163.367
R2359 B.n401 B.n400 163.367
R2360 B.n402 B.n401 163.367
R2361 B.n402 B.n245 163.367
R2362 B.n406 B.n245 163.367
R2363 B.n407 B.n406 163.367
R2364 B.n408 B.n407 163.367
R2365 B.n408 B.n243 163.367
R2366 B.n412 B.n243 163.367
R2367 B.n413 B.n412 163.367
R2368 B.n414 B.n413 163.367
R2369 B.n414 B.n241 163.367
R2370 B.n418 B.n241 163.367
R2371 B.n419 B.n418 163.367
R2372 B.n420 B.n419 163.367
R2373 B.n420 B.n239 163.367
R2374 B.n424 B.n239 163.367
R2375 B.n425 B.n424 163.367
R2376 B.n426 B.n425 163.367
R2377 B.n426 B.n237 163.367
R2378 B.n430 B.n237 163.367
R2379 B.n431 B.n430 163.367
R2380 B.n432 B.n431 163.367
R2381 B.n432 B.n235 163.367
R2382 B.n436 B.n235 163.367
R2383 B.n437 B.n436 163.367
R2384 B.n438 B.n437 163.367
R2385 B.n438 B.n233 163.367
R2386 B.n442 B.n233 163.367
R2387 B.n443 B.n442 163.367
R2388 B.n444 B.n443 163.367
R2389 B.n444 B.n231 163.367
R2390 B.n448 B.n231 163.367
R2391 B.n449 B.n448 163.367
R2392 B.n450 B.n449 163.367
R2393 B.n450 B.n229 163.367
R2394 B.n454 B.n229 163.367
R2395 B.n455 B.n454 163.367
R2396 B.n456 B.n455 163.367
R2397 B.n456 B.n227 163.367
R2398 B.n460 B.n227 163.367
R2399 B.n461 B.n460 163.367
R2400 B.n462 B.n461 163.367
R2401 B.n462 B.n225 163.367
R2402 B.n466 B.n225 163.367
R2403 B.n467 B.n466 163.367
R2404 B.n468 B.n467 163.367
R2405 B.n468 B.n223 163.367
R2406 B.n472 B.n223 163.367
R2407 B.n473 B.n472 163.367
R2408 B.n474 B.n473 163.367
R2409 B.n474 B.n221 163.367
R2410 B.n478 B.n221 163.367
R2411 B.n479 B.n478 163.367
R2412 B.n480 B.n479 163.367
R2413 B.n480 B.n217 163.367
R2414 B.n485 B.n217 163.367
R2415 B.n486 B.n485 163.367
R2416 B.n487 B.n486 163.367
R2417 B.n487 B.n215 163.367
R2418 B.n491 B.n215 163.367
R2419 B.n492 B.n491 163.367
R2420 B.n493 B.n492 163.367
R2421 B.n493 B.n213 163.367
R2422 B.n497 B.n213 163.367
R2423 B.n498 B.n497 163.367
R2424 B.n498 B.n209 163.367
R2425 B.n502 B.n209 163.367
R2426 B.n503 B.n502 163.367
R2427 B.n504 B.n503 163.367
R2428 B.n504 B.n207 163.367
R2429 B.n508 B.n207 163.367
R2430 B.n509 B.n508 163.367
R2431 B.n510 B.n509 163.367
R2432 B.n510 B.n205 163.367
R2433 B.n514 B.n205 163.367
R2434 B.n515 B.n514 163.367
R2435 B.n516 B.n515 163.367
R2436 B.n516 B.n203 163.367
R2437 B.n520 B.n203 163.367
R2438 B.n521 B.n520 163.367
R2439 B.n522 B.n521 163.367
R2440 B.n522 B.n201 163.367
R2441 B.n526 B.n201 163.367
R2442 B.n527 B.n526 163.367
R2443 B.n528 B.n527 163.367
R2444 B.n528 B.n199 163.367
R2445 B.n532 B.n199 163.367
R2446 B.n533 B.n532 163.367
R2447 B.n534 B.n533 163.367
R2448 B.n534 B.n197 163.367
R2449 B.n538 B.n197 163.367
R2450 B.n539 B.n538 163.367
R2451 B.n540 B.n539 163.367
R2452 B.n540 B.n195 163.367
R2453 B.n544 B.n195 163.367
R2454 B.n545 B.n544 163.367
R2455 B.n546 B.n545 163.367
R2456 B.n546 B.n193 163.367
R2457 B.n550 B.n193 163.367
R2458 B.n551 B.n550 163.367
R2459 B.n552 B.n551 163.367
R2460 B.n552 B.n191 163.367
R2461 B.n556 B.n191 163.367
R2462 B.n557 B.n556 163.367
R2463 B.n558 B.n557 163.367
R2464 B.n558 B.n189 163.367
R2465 B.n562 B.n189 163.367
R2466 B.n563 B.n562 163.367
R2467 B.n564 B.n563 163.367
R2468 B.n564 B.n187 163.367
R2469 B.n568 B.n187 163.367
R2470 B.n569 B.n568 163.367
R2471 B.n570 B.n569 163.367
R2472 B.n570 B.n185 163.367
R2473 B.n574 B.n185 163.367
R2474 B.n575 B.n574 163.367
R2475 B.n576 B.n575 163.367
R2476 B.n576 B.n183 163.367
R2477 B.n580 B.n183 163.367
R2478 B.n581 B.n580 163.367
R2479 B.n582 B.n581 163.367
R2480 B.n582 B.n181 163.367
R2481 B.n586 B.n181 163.367
R2482 B.n587 B.n586 163.367
R2483 B.n588 B.n587 163.367
R2484 B.n588 B.n179 163.367
R2485 B.n592 B.n179 163.367
R2486 B.n594 B.n593 163.367
R2487 B.n594 B.n177 163.367
R2488 B.n598 B.n177 163.367
R2489 B.n599 B.n598 163.367
R2490 B.n600 B.n599 163.367
R2491 B.n600 B.n175 163.367
R2492 B.n604 B.n175 163.367
R2493 B.n605 B.n604 163.367
R2494 B.n606 B.n605 163.367
R2495 B.n606 B.n173 163.367
R2496 B.n610 B.n173 163.367
R2497 B.n611 B.n610 163.367
R2498 B.n612 B.n611 163.367
R2499 B.n612 B.n171 163.367
R2500 B.n616 B.n171 163.367
R2501 B.n617 B.n616 163.367
R2502 B.n618 B.n617 163.367
R2503 B.n618 B.n169 163.367
R2504 B.n622 B.n169 163.367
R2505 B.n623 B.n622 163.367
R2506 B.n624 B.n623 163.367
R2507 B.n624 B.n167 163.367
R2508 B.n628 B.n167 163.367
R2509 B.n629 B.n628 163.367
R2510 B.n630 B.n629 163.367
R2511 B.n630 B.n165 163.367
R2512 B.n634 B.n165 163.367
R2513 B.n635 B.n634 163.367
R2514 B.n636 B.n635 163.367
R2515 B.n636 B.n163 163.367
R2516 B.n640 B.n163 163.367
R2517 B.n641 B.n640 163.367
R2518 B.n642 B.n641 163.367
R2519 B.n642 B.n161 163.367
R2520 B.n646 B.n161 163.367
R2521 B.n647 B.n646 163.367
R2522 B.n648 B.n647 163.367
R2523 B.n648 B.n159 163.367
R2524 B.n652 B.n159 163.367
R2525 B.n653 B.n652 163.367
R2526 B.n654 B.n653 163.367
R2527 B.n654 B.n157 163.367
R2528 B.n658 B.n157 163.367
R2529 B.n659 B.n658 163.367
R2530 B.n660 B.n659 163.367
R2531 B.n660 B.n155 163.367
R2532 B.n664 B.n155 163.367
R2533 B.n665 B.n664 163.367
R2534 B.n666 B.n665 163.367
R2535 B.n666 B.n153 163.367
R2536 B.n670 B.n153 163.367
R2537 B.n671 B.n670 163.367
R2538 B.n672 B.n671 163.367
R2539 B.n672 B.n151 163.367
R2540 B.n676 B.n151 163.367
R2541 B.n677 B.n676 163.367
R2542 B.n678 B.n677 163.367
R2543 B.n678 B.n149 163.367
R2544 B.n682 B.n149 163.367
R2545 B.n683 B.n682 163.367
R2546 B.n684 B.n683 163.367
R2547 B.n684 B.n147 163.367
R2548 B.n688 B.n147 163.367
R2549 B.n689 B.n688 163.367
R2550 B.n690 B.n689 163.367
R2551 B.n690 B.n145 163.367
R2552 B.n694 B.n145 163.367
R2553 B.n695 B.n694 163.367
R2554 B.n696 B.n695 163.367
R2555 B.n696 B.n143 163.367
R2556 B.n700 B.n143 163.367
R2557 B.n701 B.n700 163.367
R2558 B.n702 B.n701 163.367
R2559 B.n702 B.n141 163.367
R2560 B.n706 B.n141 163.367
R2561 B.n707 B.n706 163.367
R2562 B.n708 B.n707 163.367
R2563 B.n708 B.n139 163.367
R2564 B.n712 B.n139 163.367
R2565 B.n713 B.n712 163.367
R2566 B.n714 B.n713 163.367
R2567 B.n714 B.n137 163.367
R2568 B.n718 B.n137 163.367
R2569 B.n719 B.n718 163.367
R2570 B.n720 B.n719 163.367
R2571 B.n720 B.n135 163.367
R2572 B.n724 B.n135 163.367
R2573 B.n725 B.n724 163.367
R2574 B.n726 B.n725 163.367
R2575 B.n726 B.n133 163.367
R2576 B.n730 B.n133 163.367
R2577 B.n731 B.n730 163.367
R2578 B.n732 B.n731 163.367
R2579 B.n732 B.n131 163.367
R2580 B.n736 B.n131 163.367
R2581 B.n737 B.n736 163.367
R2582 B.n738 B.n737 163.367
R2583 B.n738 B.n129 163.367
R2584 B.n742 B.n129 163.367
R2585 B.n743 B.n742 163.367
R2586 B.n744 B.n743 163.367
R2587 B.n744 B.n127 163.367
R2588 B.n748 B.n127 163.367
R2589 B.n749 B.n748 163.367
R2590 B.n750 B.n749 163.367
R2591 B.n750 B.n125 163.367
R2592 B.n754 B.n125 163.367
R2593 B.n755 B.n754 163.367
R2594 B.n756 B.n755 163.367
R2595 B.n756 B.n123 163.367
R2596 B.n760 B.n123 163.367
R2597 B.n761 B.n760 163.367
R2598 B.n762 B.n761 163.367
R2599 B.n762 B.n121 163.367
R2600 B.n766 B.n121 163.367
R2601 B.n767 B.n766 163.367
R2602 B.n768 B.n767 163.367
R2603 B.n768 B.n119 163.367
R2604 B.n772 B.n119 163.367
R2605 B.n773 B.n772 163.367
R2606 B.n774 B.n773 163.367
R2607 B.n774 B.n117 163.367
R2608 B.n778 B.n117 163.367
R2609 B.n779 B.n778 163.367
R2610 B.n780 B.n779 163.367
R2611 B.n780 B.n115 163.367
R2612 B.n784 B.n115 163.367
R2613 B.n785 B.n784 163.367
R2614 B.n786 B.n785 163.367
R2615 B.n786 B.n113 163.367
R2616 B.n790 B.n113 163.367
R2617 B.n791 B.n790 163.367
R2618 B.n792 B.n791 163.367
R2619 B.n792 B.n111 163.367
R2620 B.n796 B.n111 163.367
R2621 B.n797 B.n796 163.367
R2622 B.n798 B.n797 163.367
R2623 B.n798 B.n109 163.367
R2624 B.n1006 B.n37 163.367
R2625 B.n1002 B.n37 163.367
R2626 B.n1002 B.n1001 163.367
R2627 B.n1001 B.n1000 163.367
R2628 B.n1000 B.n39 163.367
R2629 B.n996 B.n39 163.367
R2630 B.n996 B.n995 163.367
R2631 B.n995 B.n994 163.367
R2632 B.n994 B.n41 163.367
R2633 B.n990 B.n41 163.367
R2634 B.n990 B.n989 163.367
R2635 B.n989 B.n988 163.367
R2636 B.n988 B.n43 163.367
R2637 B.n984 B.n43 163.367
R2638 B.n984 B.n983 163.367
R2639 B.n983 B.n982 163.367
R2640 B.n982 B.n45 163.367
R2641 B.n978 B.n45 163.367
R2642 B.n978 B.n977 163.367
R2643 B.n977 B.n976 163.367
R2644 B.n976 B.n47 163.367
R2645 B.n972 B.n47 163.367
R2646 B.n972 B.n971 163.367
R2647 B.n971 B.n970 163.367
R2648 B.n970 B.n49 163.367
R2649 B.n966 B.n49 163.367
R2650 B.n966 B.n965 163.367
R2651 B.n965 B.n964 163.367
R2652 B.n964 B.n51 163.367
R2653 B.n960 B.n51 163.367
R2654 B.n960 B.n959 163.367
R2655 B.n959 B.n958 163.367
R2656 B.n958 B.n53 163.367
R2657 B.n954 B.n53 163.367
R2658 B.n954 B.n953 163.367
R2659 B.n953 B.n952 163.367
R2660 B.n952 B.n55 163.367
R2661 B.n948 B.n55 163.367
R2662 B.n948 B.n947 163.367
R2663 B.n947 B.n946 163.367
R2664 B.n946 B.n57 163.367
R2665 B.n942 B.n57 163.367
R2666 B.n942 B.n941 163.367
R2667 B.n941 B.n940 163.367
R2668 B.n940 B.n59 163.367
R2669 B.n936 B.n59 163.367
R2670 B.n936 B.n935 163.367
R2671 B.n935 B.n934 163.367
R2672 B.n934 B.n61 163.367
R2673 B.n930 B.n61 163.367
R2674 B.n930 B.n929 163.367
R2675 B.n929 B.n928 163.367
R2676 B.n928 B.n63 163.367
R2677 B.n924 B.n63 163.367
R2678 B.n924 B.n923 163.367
R2679 B.n923 B.n922 163.367
R2680 B.n922 B.n65 163.367
R2681 B.n918 B.n65 163.367
R2682 B.n918 B.n917 163.367
R2683 B.n917 B.n916 163.367
R2684 B.n916 B.n67 163.367
R2685 B.n912 B.n67 163.367
R2686 B.n912 B.n911 163.367
R2687 B.n911 B.n71 163.367
R2688 B.n907 B.n71 163.367
R2689 B.n907 B.n906 163.367
R2690 B.n906 B.n905 163.367
R2691 B.n905 B.n73 163.367
R2692 B.n901 B.n73 163.367
R2693 B.n901 B.n900 163.367
R2694 B.n900 B.n899 163.367
R2695 B.n899 B.n75 163.367
R2696 B.n894 B.n75 163.367
R2697 B.n894 B.n893 163.367
R2698 B.n893 B.n892 163.367
R2699 B.n892 B.n79 163.367
R2700 B.n888 B.n79 163.367
R2701 B.n888 B.n887 163.367
R2702 B.n887 B.n886 163.367
R2703 B.n886 B.n81 163.367
R2704 B.n882 B.n81 163.367
R2705 B.n882 B.n881 163.367
R2706 B.n881 B.n880 163.367
R2707 B.n880 B.n83 163.367
R2708 B.n876 B.n83 163.367
R2709 B.n876 B.n875 163.367
R2710 B.n875 B.n874 163.367
R2711 B.n874 B.n85 163.367
R2712 B.n870 B.n85 163.367
R2713 B.n870 B.n869 163.367
R2714 B.n869 B.n868 163.367
R2715 B.n868 B.n87 163.367
R2716 B.n864 B.n87 163.367
R2717 B.n864 B.n863 163.367
R2718 B.n863 B.n862 163.367
R2719 B.n862 B.n89 163.367
R2720 B.n858 B.n89 163.367
R2721 B.n858 B.n857 163.367
R2722 B.n857 B.n856 163.367
R2723 B.n856 B.n91 163.367
R2724 B.n852 B.n91 163.367
R2725 B.n852 B.n851 163.367
R2726 B.n851 B.n850 163.367
R2727 B.n850 B.n93 163.367
R2728 B.n846 B.n93 163.367
R2729 B.n846 B.n845 163.367
R2730 B.n845 B.n844 163.367
R2731 B.n844 B.n95 163.367
R2732 B.n840 B.n95 163.367
R2733 B.n840 B.n839 163.367
R2734 B.n839 B.n838 163.367
R2735 B.n838 B.n97 163.367
R2736 B.n834 B.n97 163.367
R2737 B.n834 B.n833 163.367
R2738 B.n833 B.n832 163.367
R2739 B.n832 B.n99 163.367
R2740 B.n828 B.n99 163.367
R2741 B.n828 B.n827 163.367
R2742 B.n827 B.n826 163.367
R2743 B.n826 B.n101 163.367
R2744 B.n822 B.n101 163.367
R2745 B.n822 B.n821 163.367
R2746 B.n821 B.n820 163.367
R2747 B.n820 B.n103 163.367
R2748 B.n816 B.n103 163.367
R2749 B.n816 B.n815 163.367
R2750 B.n815 B.n814 163.367
R2751 B.n814 B.n105 163.367
R2752 B.n810 B.n105 163.367
R2753 B.n810 B.n809 163.367
R2754 B.n809 B.n808 163.367
R2755 B.n808 B.n107 163.367
R2756 B.n804 B.n107 163.367
R2757 B.n804 B.n803 163.367
R2758 B.n803 B.n802 163.367
R2759 B.n211 B.n210 66.7156
R2760 B.n219 B.n218 66.7156
R2761 B.n69 B.n68 66.7156
R2762 B.n77 B.n76 66.7156
R2763 B.n212 B.n211 59.5399
R2764 B.n482 B.n219 59.5399
R2765 B.n70 B.n69 59.5399
R2766 B.n896 B.n77 59.5399
R2767 B.n1005 B.n36 32.6249
R2768 B.n801 B.n800 32.6249
R2769 B.n591 B.n178 32.6249
R2770 B.n387 B.n386 32.6249
R2771 B B.n1111 18.0485
R2772 B.n1005 B.n1004 10.6151
R2773 B.n1004 B.n1003 10.6151
R2774 B.n1003 B.n38 10.6151
R2775 B.n999 B.n38 10.6151
R2776 B.n999 B.n998 10.6151
R2777 B.n998 B.n997 10.6151
R2778 B.n997 B.n40 10.6151
R2779 B.n993 B.n40 10.6151
R2780 B.n993 B.n992 10.6151
R2781 B.n992 B.n991 10.6151
R2782 B.n991 B.n42 10.6151
R2783 B.n987 B.n42 10.6151
R2784 B.n987 B.n986 10.6151
R2785 B.n986 B.n985 10.6151
R2786 B.n985 B.n44 10.6151
R2787 B.n981 B.n44 10.6151
R2788 B.n981 B.n980 10.6151
R2789 B.n980 B.n979 10.6151
R2790 B.n979 B.n46 10.6151
R2791 B.n975 B.n46 10.6151
R2792 B.n975 B.n974 10.6151
R2793 B.n974 B.n973 10.6151
R2794 B.n973 B.n48 10.6151
R2795 B.n969 B.n48 10.6151
R2796 B.n969 B.n968 10.6151
R2797 B.n968 B.n967 10.6151
R2798 B.n967 B.n50 10.6151
R2799 B.n963 B.n50 10.6151
R2800 B.n963 B.n962 10.6151
R2801 B.n962 B.n961 10.6151
R2802 B.n961 B.n52 10.6151
R2803 B.n957 B.n52 10.6151
R2804 B.n957 B.n956 10.6151
R2805 B.n956 B.n955 10.6151
R2806 B.n955 B.n54 10.6151
R2807 B.n951 B.n54 10.6151
R2808 B.n951 B.n950 10.6151
R2809 B.n950 B.n949 10.6151
R2810 B.n949 B.n56 10.6151
R2811 B.n945 B.n56 10.6151
R2812 B.n945 B.n944 10.6151
R2813 B.n944 B.n943 10.6151
R2814 B.n943 B.n58 10.6151
R2815 B.n939 B.n58 10.6151
R2816 B.n939 B.n938 10.6151
R2817 B.n938 B.n937 10.6151
R2818 B.n937 B.n60 10.6151
R2819 B.n933 B.n60 10.6151
R2820 B.n933 B.n932 10.6151
R2821 B.n932 B.n931 10.6151
R2822 B.n931 B.n62 10.6151
R2823 B.n927 B.n62 10.6151
R2824 B.n927 B.n926 10.6151
R2825 B.n926 B.n925 10.6151
R2826 B.n925 B.n64 10.6151
R2827 B.n921 B.n64 10.6151
R2828 B.n921 B.n920 10.6151
R2829 B.n920 B.n919 10.6151
R2830 B.n919 B.n66 10.6151
R2831 B.n915 B.n66 10.6151
R2832 B.n915 B.n914 10.6151
R2833 B.n914 B.n913 10.6151
R2834 B.n910 B.n909 10.6151
R2835 B.n909 B.n908 10.6151
R2836 B.n908 B.n72 10.6151
R2837 B.n904 B.n72 10.6151
R2838 B.n904 B.n903 10.6151
R2839 B.n903 B.n902 10.6151
R2840 B.n902 B.n74 10.6151
R2841 B.n898 B.n74 10.6151
R2842 B.n898 B.n897 10.6151
R2843 B.n895 B.n78 10.6151
R2844 B.n891 B.n78 10.6151
R2845 B.n891 B.n890 10.6151
R2846 B.n890 B.n889 10.6151
R2847 B.n889 B.n80 10.6151
R2848 B.n885 B.n80 10.6151
R2849 B.n885 B.n884 10.6151
R2850 B.n884 B.n883 10.6151
R2851 B.n883 B.n82 10.6151
R2852 B.n879 B.n82 10.6151
R2853 B.n879 B.n878 10.6151
R2854 B.n878 B.n877 10.6151
R2855 B.n877 B.n84 10.6151
R2856 B.n873 B.n84 10.6151
R2857 B.n873 B.n872 10.6151
R2858 B.n872 B.n871 10.6151
R2859 B.n871 B.n86 10.6151
R2860 B.n867 B.n86 10.6151
R2861 B.n867 B.n866 10.6151
R2862 B.n866 B.n865 10.6151
R2863 B.n865 B.n88 10.6151
R2864 B.n861 B.n88 10.6151
R2865 B.n861 B.n860 10.6151
R2866 B.n860 B.n859 10.6151
R2867 B.n859 B.n90 10.6151
R2868 B.n855 B.n90 10.6151
R2869 B.n855 B.n854 10.6151
R2870 B.n854 B.n853 10.6151
R2871 B.n853 B.n92 10.6151
R2872 B.n849 B.n92 10.6151
R2873 B.n849 B.n848 10.6151
R2874 B.n848 B.n847 10.6151
R2875 B.n847 B.n94 10.6151
R2876 B.n843 B.n94 10.6151
R2877 B.n843 B.n842 10.6151
R2878 B.n842 B.n841 10.6151
R2879 B.n841 B.n96 10.6151
R2880 B.n837 B.n96 10.6151
R2881 B.n837 B.n836 10.6151
R2882 B.n836 B.n835 10.6151
R2883 B.n835 B.n98 10.6151
R2884 B.n831 B.n98 10.6151
R2885 B.n831 B.n830 10.6151
R2886 B.n830 B.n829 10.6151
R2887 B.n829 B.n100 10.6151
R2888 B.n825 B.n100 10.6151
R2889 B.n825 B.n824 10.6151
R2890 B.n824 B.n823 10.6151
R2891 B.n823 B.n102 10.6151
R2892 B.n819 B.n102 10.6151
R2893 B.n819 B.n818 10.6151
R2894 B.n818 B.n817 10.6151
R2895 B.n817 B.n104 10.6151
R2896 B.n813 B.n104 10.6151
R2897 B.n813 B.n812 10.6151
R2898 B.n812 B.n811 10.6151
R2899 B.n811 B.n106 10.6151
R2900 B.n807 B.n106 10.6151
R2901 B.n807 B.n806 10.6151
R2902 B.n806 B.n805 10.6151
R2903 B.n805 B.n108 10.6151
R2904 B.n801 B.n108 10.6151
R2905 B.n595 B.n178 10.6151
R2906 B.n596 B.n595 10.6151
R2907 B.n597 B.n596 10.6151
R2908 B.n597 B.n176 10.6151
R2909 B.n601 B.n176 10.6151
R2910 B.n602 B.n601 10.6151
R2911 B.n603 B.n602 10.6151
R2912 B.n603 B.n174 10.6151
R2913 B.n607 B.n174 10.6151
R2914 B.n608 B.n607 10.6151
R2915 B.n609 B.n608 10.6151
R2916 B.n609 B.n172 10.6151
R2917 B.n613 B.n172 10.6151
R2918 B.n614 B.n613 10.6151
R2919 B.n615 B.n614 10.6151
R2920 B.n615 B.n170 10.6151
R2921 B.n619 B.n170 10.6151
R2922 B.n620 B.n619 10.6151
R2923 B.n621 B.n620 10.6151
R2924 B.n621 B.n168 10.6151
R2925 B.n625 B.n168 10.6151
R2926 B.n626 B.n625 10.6151
R2927 B.n627 B.n626 10.6151
R2928 B.n627 B.n166 10.6151
R2929 B.n631 B.n166 10.6151
R2930 B.n632 B.n631 10.6151
R2931 B.n633 B.n632 10.6151
R2932 B.n633 B.n164 10.6151
R2933 B.n637 B.n164 10.6151
R2934 B.n638 B.n637 10.6151
R2935 B.n639 B.n638 10.6151
R2936 B.n639 B.n162 10.6151
R2937 B.n643 B.n162 10.6151
R2938 B.n644 B.n643 10.6151
R2939 B.n645 B.n644 10.6151
R2940 B.n645 B.n160 10.6151
R2941 B.n649 B.n160 10.6151
R2942 B.n650 B.n649 10.6151
R2943 B.n651 B.n650 10.6151
R2944 B.n651 B.n158 10.6151
R2945 B.n655 B.n158 10.6151
R2946 B.n656 B.n655 10.6151
R2947 B.n657 B.n656 10.6151
R2948 B.n657 B.n156 10.6151
R2949 B.n661 B.n156 10.6151
R2950 B.n662 B.n661 10.6151
R2951 B.n663 B.n662 10.6151
R2952 B.n663 B.n154 10.6151
R2953 B.n667 B.n154 10.6151
R2954 B.n668 B.n667 10.6151
R2955 B.n669 B.n668 10.6151
R2956 B.n669 B.n152 10.6151
R2957 B.n673 B.n152 10.6151
R2958 B.n674 B.n673 10.6151
R2959 B.n675 B.n674 10.6151
R2960 B.n675 B.n150 10.6151
R2961 B.n679 B.n150 10.6151
R2962 B.n680 B.n679 10.6151
R2963 B.n681 B.n680 10.6151
R2964 B.n681 B.n148 10.6151
R2965 B.n685 B.n148 10.6151
R2966 B.n686 B.n685 10.6151
R2967 B.n687 B.n686 10.6151
R2968 B.n687 B.n146 10.6151
R2969 B.n691 B.n146 10.6151
R2970 B.n692 B.n691 10.6151
R2971 B.n693 B.n692 10.6151
R2972 B.n693 B.n144 10.6151
R2973 B.n697 B.n144 10.6151
R2974 B.n698 B.n697 10.6151
R2975 B.n699 B.n698 10.6151
R2976 B.n699 B.n142 10.6151
R2977 B.n703 B.n142 10.6151
R2978 B.n704 B.n703 10.6151
R2979 B.n705 B.n704 10.6151
R2980 B.n705 B.n140 10.6151
R2981 B.n709 B.n140 10.6151
R2982 B.n710 B.n709 10.6151
R2983 B.n711 B.n710 10.6151
R2984 B.n711 B.n138 10.6151
R2985 B.n715 B.n138 10.6151
R2986 B.n716 B.n715 10.6151
R2987 B.n717 B.n716 10.6151
R2988 B.n717 B.n136 10.6151
R2989 B.n721 B.n136 10.6151
R2990 B.n722 B.n721 10.6151
R2991 B.n723 B.n722 10.6151
R2992 B.n723 B.n134 10.6151
R2993 B.n727 B.n134 10.6151
R2994 B.n728 B.n727 10.6151
R2995 B.n729 B.n728 10.6151
R2996 B.n729 B.n132 10.6151
R2997 B.n733 B.n132 10.6151
R2998 B.n734 B.n733 10.6151
R2999 B.n735 B.n734 10.6151
R3000 B.n735 B.n130 10.6151
R3001 B.n739 B.n130 10.6151
R3002 B.n740 B.n739 10.6151
R3003 B.n741 B.n740 10.6151
R3004 B.n741 B.n128 10.6151
R3005 B.n745 B.n128 10.6151
R3006 B.n746 B.n745 10.6151
R3007 B.n747 B.n746 10.6151
R3008 B.n747 B.n126 10.6151
R3009 B.n751 B.n126 10.6151
R3010 B.n752 B.n751 10.6151
R3011 B.n753 B.n752 10.6151
R3012 B.n753 B.n124 10.6151
R3013 B.n757 B.n124 10.6151
R3014 B.n758 B.n757 10.6151
R3015 B.n759 B.n758 10.6151
R3016 B.n759 B.n122 10.6151
R3017 B.n763 B.n122 10.6151
R3018 B.n764 B.n763 10.6151
R3019 B.n765 B.n764 10.6151
R3020 B.n765 B.n120 10.6151
R3021 B.n769 B.n120 10.6151
R3022 B.n770 B.n769 10.6151
R3023 B.n771 B.n770 10.6151
R3024 B.n771 B.n118 10.6151
R3025 B.n775 B.n118 10.6151
R3026 B.n776 B.n775 10.6151
R3027 B.n777 B.n776 10.6151
R3028 B.n777 B.n116 10.6151
R3029 B.n781 B.n116 10.6151
R3030 B.n782 B.n781 10.6151
R3031 B.n783 B.n782 10.6151
R3032 B.n783 B.n114 10.6151
R3033 B.n787 B.n114 10.6151
R3034 B.n788 B.n787 10.6151
R3035 B.n789 B.n788 10.6151
R3036 B.n789 B.n112 10.6151
R3037 B.n793 B.n112 10.6151
R3038 B.n794 B.n793 10.6151
R3039 B.n795 B.n794 10.6151
R3040 B.n795 B.n110 10.6151
R3041 B.n799 B.n110 10.6151
R3042 B.n800 B.n799 10.6151
R3043 B.n387 B.n250 10.6151
R3044 B.n391 B.n250 10.6151
R3045 B.n392 B.n391 10.6151
R3046 B.n393 B.n392 10.6151
R3047 B.n393 B.n248 10.6151
R3048 B.n397 B.n248 10.6151
R3049 B.n398 B.n397 10.6151
R3050 B.n399 B.n398 10.6151
R3051 B.n399 B.n246 10.6151
R3052 B.n403 B.n246 10.6151
R3053 B.n404 B.n403 10.6151
R3054 B.n405 B.n404 10.6151
R3055 B.n405 B.n244 10.6151
R3056 B.n409 B.n244 10.6151
R3057 B.n410 B.n409 10.6151
R3058 B.n411 B.n410 10.6151
R3059 B.n411 B.n242 10.6151
R3060 B.n415 B.n242 10.6151
R3061 B.n416 B.n415 10.6151
R3062 B.n417 B.n416 10.6151
R3063 B.n417 B.n240 10.6151
R3064 B.n421 B.n240 10.6151
R3065 B.n422 B.n421 10.6151
R3066 B.n423 B.n422 10.6151
R3067 B.n423 B.n238 10.6151
R3068 B.n427 B.n238 10.6151
R3069 B.n428 B.n427 10.6151
R3070 B.n429 B.n428 10.6151
R3071 B.n429 B.n236 10.6151
R3072 B.n433 B.n236 10.6151
R3073 B.n434 B.n433 10.6151
R3074 B.n435 B.n434 10.6151
R3075 B.n435 B.n234 10.6151
R3076 B.n439 B.n234 10.6151
R3077 B.n440 B.n439 10.6151
R3078 B.n441 B.n440 10.6151
R3079 B.n441 B.n232 10.6151
R3080 B.n445 B.n232 10.6151
R3081 B.n446 B.n445 10.6151
R3082 B.n447 B.n446 10.6151
R3083 B.n447 B.n230 10.6151
R3084 B.n451 B.n230 10.6151
R3085 B.n452 B.n451 10.6151
R3086 B.n453 B.n452 10.6151
R3087 B.n453 B.n228 10.6151
R3088 B.n457 B.n228 10.6151
R3089 B.n458 B.n457 10.6151
R3090 B.n459 B.n458 10.6151
R3091 B.n459 B.n226 10.6151
R3092 B.n463 B.n226 10.6151
R3093 B.n464 B.n463 10.6151
R3094 B.n465 B.n464 10.6151
R3095 B.n465 B.n224 10.6151
R3096 B.n469 B.n224 10.6151
R3097 B.n470 B.n469 10.6151
R3098 B.n471 B.n470 10.6151
R3099 B.n471 B.n222 10.6151
R3100 B.n475 B.n222 10.6151
R3101 B.n476 B.n475 10.6151
R3102 B.n477 B.n476 10.6151
R3103 B.n477 B.n220 10.6151
R3104 B.n481 B.n220 10.6151
R3105 B.n484 B.n483 10.6151
R3106 B.n484 B.n216 10.6151
R3107 B.n488 B.n216 10.6151
R3108 B.n489 B.n488 10.6151
R3109 B.n490 B.n489 10.6151
R3110 B.n490 B.n214 10.6151
R3111 B.n494 B.n214 10.6151
R3112 B.n495 B.n494 10.6151
R3113 B.n496 B.n495 10.6151
R3114 B.n500 B.n499 10.6151
R3115 B.n501 B.n500 10.6151
R3116 B.n501 B.n208 10.6151
R3117 B.n505 B.n208 10.6151
R3118 B.n506 B.n505 10.6151
R3119 B.n507 B.n506 10.6151
R3120 B.n507 B.n206 10.6151
R3121 B.n511 B.n206 10.6151
R3122 B.n512 B.n511 10.6151
R3123 B.n513 B.n512 10.6151
R3124 B.n513 B.n204 10.6151
R3125 B.n517 B.n204 10.6151
R3126 B.n518 B.n517 10.6151
R3127 B.n519 B.n518 10.6151
R3128 B.n519 B.n202 10.6151
R3129 B.n523 B.n202 10.6151
R3130 B.n524 B.n523 10.6151
R3131 B.n525 B.n524 10.6151
R3132 B.n525 B.n200 10.6151
R3133 B.n529 B.n200 10.6151
R3134 B.n530 B.n529 10.6151
R3135 B.n531 B.n530 10.6151
R3136 B.n531 B.n198 10.6151
R3137 B.n535 B.n198 10.6151
R3138 B.n536 B.n535 10.6151
R3139 B.n537 B.n536 10.6151
R3140 B.n537 B.n196 10.6151
R3141 B.n541 B.n196 10.6151
R3142 B.n542 B.n541 10.6151
R3143 B.n543 B.n542 10.6151
R3144 B.n543 B.n194 10.6151
R3145 B.n547 B.n194 10.6151
R3146 B.n548 B.n547 10.6151
R3147 B.n549 B.n548 10.6151
R3148 B.n549 B.n192 10.6151
R3149 B.n553 B.n192 10.6151
R3150 B.n554 B.n553 10.6151
R3151 B.n555 B.n554 10.6151
R3152 B.n555 B.n190 10.6151
R3153 B.n559 B.n190 10.6151
R3154 B.n560 B.n559 10.6151
R3155 B.n561 B.n560 10.6151
R3156 B.n561 B.n188 10.6151
R3157 B.n565 B.n188 10.6151
R3158 B.n566 B.n565 10.6151
R3159 B.n567 B.n566 10.6151
R3160 B.n567 B.n186 10.6151
R3161 B.n571 B.n186 10.6151
R3162 B.n572 B.n571 10.6151
R3163 B.n573 B.n572 10.6151
R3164 B.n573 B.n184 10.6151
R3165 B.n577 B.n184 10.6151
R3166 B.n578 B.n577 10.6151
R3167 B.n579 B.n578 10.6151
R3168 B.n579 B.n182 10.6151
R3169 B.n583 B.n182 10.6151
R3170 B.n584 B.n583 10.6151
R3171 B.n585 B.n584 10.6151
R3172 B.n585 B.n180 10.6151
R3173 B.n589 B.n180 10.6151
R3174 B.n590 B.n589 10.6151
R3175 B.n591 B.n590 10.6151
R3176 B.n386 B.n385 10.6151
R3177 B.n385 B.n252 10.6151
R3178 B.n381 B.n252 10.6151
R3179 B.n381 B.n380 10.6151
R3180 B.n380 B.n379 10.6151
R3181 B.n379 B.n254 10.6151
R3182 B.n375 B.n254 10.6151
R3183 B.n375 B.n374 10.6151
R3184 B.n374 B.n373 10.6151
R3185 B.n373 B.n256 10.6151
R3186 B.n369 B.n256 10.6151
R3187 B.n369 B.n368 10.6151
R3188 B.n368 B.n367 10.6151
R3189 B.n367 B.n258 10.6151
R3190 B.n363 B.n258 10.6151
R3191 B.n363 B.n362 10.6151
R3192 B.n362 B.n361 10.6151
R3193 B.n361 B.n260 10.6151
R3194 B.n357 B.n260 10.6151
R3195 B.n357 B.n356 10.6151
R3196 B.n356 B.n355 10.6151
R3197 B.n355 B.n262 10.6151
R3198 B.n351 B.n262 10.6151
R3199 B.n351 B.n350 10.6151
R3200 B.n350 B.n349 10.6151
R3201 B.n349 B.n264 10.6151
R3202 B.n345 B.n264 10.6151
R3203 B.n345 B.n344 10.6151
R3204 B.n344 B.n343 10.6151
R3205 B.n343 B.n266 10.6151
R3206 B.n339 B.n266 10.6151
R3207 B.n339 B.n338 10.6151
R3208 B.n338 B.n337 10.6151
R3209 B.n337 B.n268 10.6151
R3210 B.n333 B.n268 10.6151
R3211 B.n333 B.n332 10.6151
R3212 B.n332 B.n331 10.6151
R3213 B.n331 B.n270 10.6151
R3214 B.n327 B.n270 10.6151
R3215 B.n327 B.n326 10.6151
R3216 B.n326 B.n325 10.6151
R3217 B.n325 B.n272 10.6151
R3218 B.n321 B.n272 10.6151
R3219 B.n321 B.n320 10.6151
R3220 B.n320 B.n319 10.6151
R3221 B.n319 B.n274 10.6151
R3222 B.n315 B.n274 10.6151
R3223 B.n315 B.n314 10.6151
R3224 B.n314 B.n313 10.6151
R3225 B.n313 B.n276 10.6151
R3226 B.n309 B.n276 10.6151
R3227 B.n309 B.n308 10.6151
R3228 B.n308 B.n307 10.6151
R3229 B.n307 B.n278 10.6151
R3230 B.n303 B.n278 10.6151
R3231 B.n303 B.n302 10.6151
R3232 B.n302 B.n301 10.6151
R3233 B.n301 B.n280 10.6151
R3234 B.n297 B.n280 10.6151
R3235 B.n297 B.n296 10.6151
R3236 B.n296 B.n295 10.6151
R3237 B.n295 B.n282 10.6151
R3238 B.n291 B.n282 10.6151
R3239 B.n291 B.n290 10.6151
R3240 B.n290 B.n289 10.6151
R3241 B.n289 B.n284 10.6151
R3242 B.n285 B.n284 10.6151
R3243 B.n285 B.n0 10.6151
R3244 B.n1107 B.n1 10.6151
R3245 B.n1107 B.n1106 10.6151
R3246 B.n1106 B.n1105 10.6151
R3247 B.n1105 B.n4 10.6151
R3248 B.n1101 B.n4 10.6151
R3249 B.n1101 B.n1100 10.6151
R3250 B.n1100 B.n1099 10.6151
R3251 B.n1099 B.n6 10.6151
R3252 B.n1095 B.n6 10.6151
R3253 B.n1095 B.n1094 10.6151
R3254 B.n1094 B.n1093 10.6151
R3255 B.n1093 B.n8 10.6151
R3256 B.n1089 B.n8 10.6151
R3257 B.n1089 B.n1088 10.6151
R3258 B.n1088 B.n1087 10.6151
R3259 B.n1087 B.n10 10.6151
R3260 B.n1083 B.n10 10.6151
R3261 B.n1083 B.n1082 10.6151
R3262 B.n1082 B.n1081 10.6151
R3263 B.n1081 B.n12 10.6151
R3264 B.n1077 B.n12 10.6151
R3265 B.n1077 B.n1076 10.6151
R3266 B.n1076 B.n1075 10.6151
R3267 B.n1075 B.n14 10.6151
R3268 B.n1071 B.n14 10.6151
R3269 B.n1071 B.n1070 10.6151
R3270 B.n1070 B.n1069 10.6151
R3271 B.n1069 B.n16 10.6151
R3272 B.n1065 B.n16 10.6151
R3273 B.n1065 B.n1064 10.6151
R3274 B.n1064 B.n1063 10.6151
R3275 B.n1063 B.n18 10.6151
R3276 B.n1059 B.n18 10.6151
R3277 B.n1059 B.n1058 10.6151
R3278 B.n1058 B.n1057 10.6151
R3279 B.n1057 B.n20 10.6151
R3280 B.n1053 B.n20 10.6151
R3281 B.n1053 B.n1052 10.6151
R3282 B.n1052 B.n1051 10.6151
R3283 B.n1051 B.n22 10.6151
R3284 B.n1047 B.n22 10.6151
R3285 B.n1047 B.n1046 10.6151
R3286 B.n1046 B.n1045 10.6151
R3287 B.n1045 B.n24 10.6151
R3288 B.n1041 B.n24 10.6151
R3289 B.n1041 B.n1040 10.6151
R3290 B.n1040 B.n1039 10.6151
R3291 B.n1039 B.n26 10.6151
R3292 B.n1035 B.n26 10.6151
R3293 B.n1035 B.n1034 10.6151
R3294 B.n1034 B.n1033 10.6151
R3295 B.n1033 B.n28 10.6151
R3296 B.n1029 B.n28 10.6151
R3297 B.n1029 B.n1028 10.6151
R3298 B.n1028 B.n1027 10.6151
R3299 B.n1027 B.n30 10.6151
R3300 B.n1023 B.n30 10.6151
R3301 B.n1023 B.n1022 10.6151
R3302 B.n1022 B.n1021 10.6151
R3303 B.n1021 B.n32 10.6151
R3304 B.n1017 B.n32 10.6151
R3305 B.n1017 B.n1016 10.6151
R3306 B.n1016 B.n1015 10.6151
R3307 B.n1015 B.n34 10.6151
R3308 B.n1011 B.n34 10.6151
R3309 B.n1011 B.n1010 10.6151
R3310 B.n1010 B.n1009 10.6151
R3311 B.n1009 B.n36 10.6151
R3312 B.n913 B.n70 9.36635
R3313 B.n896 B.n895 9.36635
R3314 B.n482 B.n481 9.36635
R3315 B.n499 B.n212 9.36635
R3316 B.n1111 B.n0 2.81026
R3317 B.n1111 B.n1 2.81026
R3318 B.n910 B.n70 1.24928
R3319 B.n897 B.n896 1.24928
R3320 B.n483 B.n482 1.24928
R3321 B.n496 B.n212 1.24928
C0 VP VTAIL 18.0401f
C1 w_n5098_n4850# VDD1 3.49538f
C2 VN VTAIL 18.0258f
C3 w_n5098_n4850# VDD2 3.66544f
C4 B VDD1 3.27143f
C5 VP VDD1 17.9935f
C6 B VDD2 3.4092f
C7 VN VDD1 0.154676f
C8 VP VDD2 0.649307f
C9 w_n5098_n4850# B 13.4821f
C10 VTAIL VDD1 13.7122f
C11 VN VDD2 17.5038f
C12 w_n5098_n4850# VP 11.8606f
C13 VTAIL VDD2 13.7656f
C14 w_n5098_n4850# VN 11.1953f
C15 w_n5098_n4850# VTAIL 4.30409f
C16 B VP 2.62161f
C17 B VN 1.50005f
C18 VDD1 VDD2 2.50833f
C19 B VTAIL 5.6464f
C20 VP VN 10.524f
C21 VDD2 VSUBS 2.49365f
C22 VDD1 VSUBS 2.361803f
C23 VTAIL VSUBS 1.682656f
C24 VN VSUBS 8.79991f
C25 VP VSUBS 5.167387f
C26 B VSUBS 6.624949f
C27 w_n5098_n4850# VSUBS 0.302026p
C28 B.n0 VSUBS 0.004836f
C29 B.n1 VSUBS 0.004836f
C30 B.n2 VSUBS 0.007647f
C31 B.n3 VSUBS 0.007647f
C32 B.n4 VSUBS 0.007647f
C33 B.n5 VSUBS 0.007647f
C34 B.n6 VSUBS 0.007647f
C35 B.n7 VSUBS 0.007647f
C36 B.n8 VSUBS 0.007647f
C37 B.n9 VSUBS 0.007647f
C38 B.n10 VSUBS 0.007647f
C39 B.n11 VSUBS 0.007647f
C40 B.n12 VSUBS 0.007647f
C41 B.n13 VSUBS 0.007647f
C42 B.n14 VSUBS 0.007647f
C43 B.n15 VSUBS 0.007647f
C44 B.n16 VSUBS 0.007647f
C45 B.n17 VSUBS 0.007647f
C46 B.n18 VSUBS 0.007647f
C47 B.n19 VSUBS 0.007647f
C48 B.n20 VSUBS 0.007647f
C49 B.n21 VSUBS 0.007647f
C50 B.n22 VSUBS 0.007647f
C51 B.n23 VSUBS 0.007647f
C52 B.n24 VSUBS 0.007647f
C53 B.n25 VSUBS 0.007647f
C54 B.n26 VSUBS 0.007647f
C55 B.n27 VSUBS 0.007647f
C56 B.n28 VSUBS 0.007647f
C57 B.n29 VSUBS 0.007647f
C58 B.n30 VSUBS 0.007647f
C59 B.n31 VSUBS 0.007647f
C60 B.n32 VSUBS 0.007647f
C61 B.n33 VSUBS 0.007647f
C62 B.n34 VSUBS 0.007647f
C63 B.n35 VSUBS 0.007647f
C64 B.n36 VSUBS 0.017737f
C65 B.n37 VSUBS 0.007647f
C66 B.n38 VSUBS 0.007647f
C67 B.n39 VSUBS 0.007647f
C68 B.n40 VSUBS 0.007647f
C69 B.n41 VSUBS 0.007647f
C70 B.n42 VSUBS 0.007647f
C71 B.n43 VSUBS 0.007647f
C72 B.n44 VSUBS 0.007647f
C73 B.n45 VSUBS 0.007647f
C74 B.n46 VSUBS 0.007647f
C75 B.n47 VSUBS 0.007647f
C76 B.n48 VSUBS 0.007647f
C77 B.n49 VSUBS 0.007647f
C78 B.n50 VSUBS 0.007647f
C79 B.n51 VSUBS 0.007647f
C80 B.n52 VSUBS 0.007647f
C81 B.n53 VSUBS 0.007647f
C82 B.n54 VSUBS 0.007647f
C83 B.n55 VSUBS 0.007647f
C84 B.n56 VSUBS 0.007647f
C85 B.n57 VSUBS 0.007647f
C86 B.n58 VSUBS 0.007647f
C87 B.n59 VSUBS 0.007647f
C88 B.n60 VSUBS 0.007647f
C89 B.n61 VSUBS 0.007647f
C90 B.n62 VSUBS 0.007647f
C91 B.n63 VSUBS 0.007647f
C92 B.n64 VSUBS 0.007647f
C93 B.n65 VSUBS 0.007647f
C94 B.n66 VSUBS 0.007647f
C95 B.n67 VSUBS 0.007647f
C96 B.t11 VSUBS 0.42078f
C97 B.t10 VSUBS 0.463539f
C98 B.t9 VSUBS 2.94886f
C99 B.n68 VSUBS 0.725822f
C100 B.n69 VSUBS 0.379834f
C101 B.n70 VSUBS 0.017717f
C102 B.n71 VSUBS 0.007647f
C103 B.n72 VSUBS 0.007647f
C104 B.n73 VSUBS 0.007647f
C105 B.n74 VSUBS 0.007647f
C106 B.n75 VSUBS 0.007647f
C107 B.t2 VSUBS 0.420784f
C108 B.t1 VSUBS 0.463543f
C109 B.t0 VSUBS 2.94886f
C110 B.n76 VSUBS 0.725819f
C111 B.n77 VSUBS 0.37983f
C112 B.n78 VSUBS 0.007647f
C113 B.n79 VSUBS 0.007647f
C114 B.n80 VSUBS 0.007647f
C115 B.n81 VSUBS 0.007647f
C116 B.n82 VSUBS 0.007647f
C117 B.n83 VSUBS 0.007647f
C118 B.n84 VSUBS 0.007647f
C119 B.n85 VSUBS 0.007647f
C120 B.n86 VSUBS 0.007647f
C121 B.n87 VSUBS 0.007647f
C122 B.n88 VSUBS 0.007647f
C123 B.n89 VSUBS 0.007647f
C124 B.n90 VSUBS 0.007647f
C125 B.n91 VSUBS 0.007647f
C126 B.n92 VSUBS 0.007647f
C127 B.n93 VSUBS 0.007647f
C128 B.n94 VSUBS 0.007647f
C129 B.n95 VSUBS 0.007647f
C130 B.n96 VSUBS 0.007647f
C131 B.n97 VSUBS 0.007647f
C132 B.n98 VSUBS 0.007647f
C133 B.n99 VSUBS 0.007647f
C134 B.n100 VSUBS 0.007647f
C135 B.n101 VSUBS 0.007647f
C136 B.n102 VSUBS 0.007647f
C137 B.n103 VSUBS 0.007647f
C138 B.n104 VSUBS 0.007647f
C139 B.n105 VSUBS 0.007647f
C140 B.n106 VSUBS 0.007647f
C141 B.n107 VSUBS 0.007647f
C142 B.n108 VSUBS 0.007647f
C143 B.n109 VSUBS 0.017737f
C144 B.n110 VSUBS 0.007647f
C145 B.n111 VSUBS 0.007647f
C146 B.n112 VSUBS 0.007647f
C147 B.n113 VSUBS 0.007647f
C148 B.n114 VSUBS 0.007647f
C149 B.n115 VSUBS 0.007647f
C150 B.n116 VSUBS 0.007647f
C151 B.n117 VSUBS 0.007647f
C152 B.n118 VSUBS 0.007647f
C153 B.n119 VSUBS 0.007647f
C154 B.n120 VSUBS 0.007647f
C155 B.n121 VSUBS 0.007647f
C156 B.n122 VSUBS 0.007647f
C157 B.n123 VSUBS 0.007647f
C158 B.n124 VSUBS 0.007647f
C159 B.n125 VSUBS 0.007647f
C160 B.n126 VSUBS 0.007647f
C161 B.n127 VSUBS 0.007647f
C162 B.n128 VSUBS 0.007647f
C163 B.n129 VSUBS 0.007647f
C164 B.n130 VSUBS 0.007647f
C165 B.n131 VSUBS 0.007647f
C166 B.n132 VSUBS 0.007647f
C167 B.n133 VSUBS 0.007647f
C168 B.n134 VSUBS 0.007647f
C169 B.n135 VSUBS 0.007647f
C170 B.n136 VSUBS 0.007647f
C171 B.n137 VSUBS 0.007647f
C172 B.n138 VSUBS 0.007647f
C173 B.n139 VSUBS 0.007647f
C174 B.n140 VSUBS 0.007647f
C175 B.n141 VSUBS 0.007647f
C176 B.n142 VSUBS 0.007647f
C177 B.n143 VSUBS 0.007647f
C178 B.n144 VSUBS 0.007647f
C179 B.n145 VSUBS 0.007647f
C180 B.n146 VSUBS 0.007647f
C181 B.n147 VSUBS 0.007647f
C182 B.n148 VSUBS 0.007647f
C183 B.n149 VSUBS 0.007647f
C184 B.n150 VSUBS 0.007647f
C185 B.n151 VSUBS 0.007647f
C186 B.n152 VSUBS 0.007647f
C187 B.n153 VSUBS 0.007647f
C188 B.n154 VSUBS 0.007647f
C189 B.n155 VSUBS 0.007647f
C190 B.n156 VSUBS 0.007647f
C191 B.n157 VSUBS 0.007647f
C192 B.n158 VSUBS 0.007647f
C193 B.n159 VSUBS 0.007647f
C194 B.n160 VSUBS 0.007647f
C195 B.n161 VSUBS 0.007647f
C196 B.n162 VSUBS 0.007647f
C197 B.n163 VSUBS 0.007647f
C198 B.n164 VSUBS 0.007647f
C199 B.n165 VSUBS 0.007647f
C200 B.n166 VSUBS 0.007647f
C201 B.n167 VSUBS 0.007647f
C202 B.n168 VSUBS 0.007647f
C203 B.n169 VSUBS 0.007647f
C204 B.n170 VSUBS 0.007647f
C205 B.n171 VSUBS 0.007647f
C206 B.n172 VSUBS 0.007647f
C207 B.n173 VSUBS 0.007647f
C208 B.n174 VSUBS 0.007647f
C209 B.n175 VSUBS 0.007647f
C210 B.n176 VSUBS 0.007647f
C211 B.n177 VSUBS 0.007647f
C212 B.n178 VSUBS 0.017737f
C213 B.n179 VSUBS 0.007647f
C214 B.n180 VSUBS 0.007647f
C215 B.n181 VSUBS 0.007647f
C216 B.n182 VSUBS 0.007647f
C217 B.n183 VSUBS 0.007647f
C218 B.n184 VSUBS 0.007647f
C219 B.n185 VSUBS 0.007647f
C220 B.n186 VSUBS 0.007647f
C221 B.n187 VSUBS 0.007647f
C222 B.n188 VSUBS 0.007647f
C223 B.n189 VSUBS 0.007647f
C224 B.n190 VSUBS 0.007647f
C225 B.n191 VSUBS 0.007647f
C226 B.n192 VSUBS 0.007647f
C227 B.n193 VSUBS 0.007647f
C228 B.n194 VSUBS 0.007647f
C229 B.n195 VSUBS 0.007647f
C230 B.n196 VSUBS 0.007647f
C231 B.n197 VSUBS 0.007647f
C232 B.n198 VSUBS 0.007647f
C233 B.n199 VSUBS 0.007647f
C234 B.n200 VSUBS 0.007647f
C235 B.n201 VSUBS 0.007647f
C236 B.n202 VSUBS 0.007647f
C237 B.n203 VSUBS 0.007647f
C238 B.n204 VSUBS 0.007647f
C239 B.n205 VSUBS 0.007647f
C240 B.n206 VSUBS 0.007647f
C241 B.n207 VSUBS 0.007647f
C242 B.n208 VSUBS 0.007647f
C243 B.n209 VSUBS 0.007647f
C244 B.t7 VSUBS 0.420784f
C245 B.t8 VSUBS 0.463543f
C246 B.t6 VSUBS 2.94886f
C247 B.n210 VSUBS 0.725819f
C248 B.n211 VSUBS 0.37983f
C249 B.n212 VSUBS 0.017717f
C250 B.n213 VSUBS 0.007647f
C251 B.n214 VSUBS 0.007647f
C252 B.n215 VSUBS 0.007647f
C253 B.n216 VSUBS 0.007647f
C254 B.n217 VSUBS 0.007647f
C255 B.t4 VSUBS 0.42078f
C256 B.t5 VSUBS 0.463539f
C257 B.t3 VSUBS 2.94886f
C258 B.n218 VSUBS 0.725822f
C259 B.n219 VSUBS 0.379834f
C260 B.n220 VSUBS 0.007647f
C261 B.n221 VSUBS 0.007647f
C262 B.n222 VSUBS 0.007647f
C263 B.n223 VSUBS 0.007647f
C264 B.n224 VSUBS 0.007647f
C265 B.n225 VSUBS 0.007647f
C266 B.n226 VSUBS 0.007647f
C267 B.n227 VSUBS 0.007647f
C268 B.n228 VSUBS 0.007647f
C269 B.n229 VSUBS 0.007647f
C270 B.n230 VSUBS 0.007647f
C271 B.n231 VSUBS 0.007647f
C272 B.n232 VSUBS 0.007647f
C273 B.n233 VSUBS 0.007647f
C274 B.n234 VSUBS 0.007647f
C275 B.n235 VSUBS 0.007647f
C276 B.n236 VSUBS 0.007647f
C277 B.n237 VSUBS 0.007647f
C278 B.n238 VSUBS 0.007647f
C279 B.n239 VSUBS 0.007647f
C280 B.n240 VSUBS 0.007647f
C281 B.n241 VSUBS 0.007647f
C282 B.n242 VSUBS 0.007647f
C283 B.n243 VSUBS 0.007647f
C284 B.n244 VSUBS 0.007647f
C285 B.n245 VSUBS 0.007647f
C286 B.n246 VSUBS 0.007647f
C287 B.n247 VSUBS 0.007647f
C288 B.n248 VSUBS 0.007647f
C289 B.n249 VSUBS 0.007647f
C290 B.n250 VSUBS 0.007647f
C291 B.n251 VSUBS 0.017737f
C292 B.n252 VSUBS 0.007647f
C293 B.n253 VSUBS 0.007647f
C294 B.n254 VSUBS 0.007647f
C295 B.n255 VSUBS 0.007647f
C296 B.n256 VSUBS 0.007647f
C297 B.n257 VSUBS 0.007647f
C298 B.n258 VSUBS 0.007647f
C299 B.n259 VSUBS 0.007647f
C300 B.n260 VSUBS 0.007647f
C301 B.n261 VSUBS 0.007647f
C302 B.n262 VSUBS 0.007647f
C303 B.n263 VSUBS 0.007647f
C304 B.n264 VSUBS 0.007647f
C305 B.n265 VSUBS 0.007647f
C306 B.n266 VSUBS 0.007647f
C307 B.n267 VSUBS 0.007647f
C308 B.n268 VSUBS 0.007647f
C309 B.n269 VSUBS 0.007647f
C310 B.n270 VSUBS 0.007647f
C311 B.n271 VSUBS 0.007647f
C312 B.n272 VSUBS 0.007647f
C313 B.n273 VSUBS 0.007647f
C314 B.n274 VSUBS 0.007647f
C315 B.n275 VSUBS 0.007647f
C316 B.n276 VSUBS 0.007647f
C317 B.n277 VSUBS 0.007647f
C318 B.n278 VSUBS 0.007647f
C319 B.n279 VSUBS 0.007647f
C320 B.n280 VSUBS 0.007647f
C321 B.n281 VSUBS 0.007647f
C322 B.n282 VSUBS 0.007647f
C323 B.n283 VSUBS 0.007647f
C324 B.n284 VSUBS 0.007647f
C325 B.n285 VSUBS 0.007647f
C326 B.n286 VSUBS 0.007647f
C327 B.n287 VSUBS 0.007647f
C328 B.n288 VSUBS 0.007647f
C329 B.n289 VSUBS 0.007647f
C330 B.n290 VSUBS 0.007647f
C331 B.n291 VSUBS 0.007647f
C332 B.n292 VSUBS 0.007647f
C333 B.n293 VSUBS 0.007647f
C334 B.n294 VSUBS 0.007647f
C335 B.n295 VSUBS 0.007647f
C336 B.n296 VSUBS 0.007647f
C337 B.n297 VSUBS 0.007647f
C338 B.n298 VSUBS 0.007647f
C339 B.n299 VSUBS 0.007647f
C340 B.n300 VSUBS 0.007647f
C341 B.n301 VSUBS 0.007647f
C342 B.n302 VSUBS 0.007647f
C343 B.n303 VSUBS 0.007647f
C344 B.n304 VSUBS 0.007647f
C345 B.n305 VSUBS 0.007647f
C346 B.n306 VSUBS 0.007647f
C347 B.n307 VSUBS 0.007647f
C348 B.n308 VSUBS 0.007647f
C349 B.n309 VSUBS 0.007647f
C350 B.n310 VSUBS 0.007647f
C351 B.n311 VSUBS 0.007647f
C352 B.n312 VSUBS 0.007647f
C353 B.n313 VSUBS 0.007647f
C354 B.n314 VSUBS 0.007647f
C355 B.n315 VSUBS 0.007647f
C356 B.n316 VSUBS 0.007647f
C357 B.n317 VSUBS 0.007647f
C358 B.n318 VSUBS 0.007647f
C359 B.n319 VSUBS 0.007647f
C360 B.n320 VSUBS 0.007647f
C361 B.n321 VSUBS 0.007647f
C362 B.n322 VSUBS 0.007647f
C363 B.n323 VSUBS 0.007647f
C364 B.n324 VSUBS 0.007647f
C365 B.n325 VSUBS 0.007647f
C366 B.n326 VSUBS 0.007647f
C367 B.n327 VSUBS 0.007647f
C368 B.n328 VSUBS 0.007647f
C369 B.n329 VSUBS 0.007647f
C370 B.n330 VSUBS 0.007647f
C371 B.n331 VSUBS 0.007647f
C372 B.n332 VSUBS 0.007647f
C373 B.n333 VSUBS 0.007647f
C374 B.n334 VSUBS 0.007647f
C375 B.n335 VSUBS 0.007647f
C376 B.n336 VSUBS 0.007647f
C377 B.n337 VSUBS 0.007647f
C378 B.n338 VSUBS 0.007647f
C379 B.n339 VSUBS 0.007647f
C380 B.n340 VSUBS 0.007647f
C381 B.n341 VSUBS 0.007647f
C382 B.n342 VSUBS 0.007647f
C383 B.n343 VSUBS 0.007647f
C384 B.n344 VSUBS 0.007647f
C385 B.n345 VSUBS 0.007647f
C386 B.n346 VSUBS 0.007647f
C387 B.n347 VSUBS 0.007647f
C388 B.n348 VSUBS 0.007647f
C389 B.n349 VSUBS 0.007647f
C390 B.n350 VSUBS 0.007647f
C391 B.n351 VSUBS 0.007647f
C392 B.n352 VSUBS 0.007647f
C393 B.n353 VSUBS 0.007647f
C394 B.n354 VSUBS 0.007647f
C395 B.n355 VSUBS 0.007647f
C396 B.n356 VSUBS 0.007647f
C397 B.n357 VSUBS 0.007647f
C398 B.n358 VSUBS 0.007647f
C399 B.n359 VSUBS 0.007647f
C400 B.n360 VSUBS 0.007647f
C401 B.n361 VSUBS 0.007647f
C402 B.n362 VSUBS 0.007647f
C403 B.n363 VSUBS 0.007647f
C404 B.n364 VSUBS 0.007647f
C405 B.n365 VSUBS 0.007647f
C406 B.n366 VSUBS 0.007647f
C407 B.n367 VSUBS 0.007647f
C408 B.n368 VSUBS 0.007647f
C409 B.n369 VSUBS 0.007647f
C410 B.n370 VSUBS 0.007647f
C411 B.n371 VSUBS 0.007647f
C412 B.n372 VSUBS 0.007647f
C413 B.n373 VSUBS 0.007647f
C414 B.n374 VSUBS 0.007647f
C415 B.n375 VSUBS 0.007647f
C416 B.n376 VSUBS 0.007647f
C417 B.n377 VSUBS 0.007647f
C418 B.n378 VSUBS 0.007647f
C419 B.n379 VSUBS 0.007647f
C420 B.n380 VSUBS 0.007647f
C421 B.n381 VSUBS 0.007647f
C422 B.n382 VSUBS 0.007647f
C423 B.n383 VSUBS 0.007647f
C424 B.n384 VSUBS 0.007647f
C425 B.n385 VSUBS 0.007647f
C426 B.n386 VSUBS 0.017737f
C427 B.n387 VSUBS 0.018024f
C428 B.n388 VSUBS 0.018024f
C429 B.n389 VSUBS 0.007647f
C430 B.n390 VSUBS 0.007647f
C431 B.n391 VSUBS 0.007647f
C432 B.n392 VSUBS 0.007647f
C433 B.n393 VSUBS 0.007647f
C434 B.n394 VSUBS 0.007647f
C435 B.n395 VSUBS 0.007647f
C436 B.n396 VSUBS 0.007647f
C437 B.n397 VSUBS 0.007647f
C438 B.n398 VSUBS 0.007647f
C439 B.n399 VSUBS 0.007647f
C440 B.n400 VSUBS 0.007647f
C441 B.n401 VSUBS 0.007647f
C442 B.n402 VSUBS 0.007647f
C443 B.n403 VSUBS 0.007647f
C444 B.n404 VSUBS 0.007647f
C445 B.n405 VSUBS 0.007647f
C446 B.n406 VSUBS 0.007647f
C447 B.n407 VSUBS 0.007647f
C448 B.n408 VSUBS 0.007647f
C449 B.n409 VSUBS 0.007647f
C450 B.n410 VSUBS 0.007647f
C451 B.n411 VSUBS 0.007647f
C452 B.n412 VSUBS 0.007647f
C453 B.n413 VSUBS 0.007647f
C454 B.n414 VSUBS 0.007647f
C455 B.n415 VSUBS 0.007647f
C456 B.n416 VSUBS 0.007647f
C457 B.n417 VSUBS 0.007647f
C458 B.n418 VSUBS 0.007647f
C459 B.n419 VSUBS 0.007647f
C460 B.n420 VSUBS 0.007647f
C461 B.n421 VSUBS 0.007647f
C462 B.n422 VSUBS 0.007647f
C463 B.n423 VSUBS 0.007647f
C464 B.n424 VSUBS 0.007647f
C465 B.n425 VSUBS 0.007647f
C466 B.n426 VSUBS 0.007647f
C467 B.n427 VSUBS 0.007647f
C468 B.n428 VSUBS 0.007647f
C469 B.n429 VSUBS 0.007647f
C470 B.n430 VSUBS 0.007647f
C471 B.n431 VSUBS 0.007647f
C472 B.n432 VSUBS 0.007647f
C473 B.n433 VSUBS 0.007647f
C474 B.n434 VSUBS 0.007647f
C475 B.n435 VSUBS 0.007647f
C476 B.n436 VSUBS 0.007647f
C477 B.n437 VSUBS 0.007647f
C478 B.n438 VSUBS 0.007647f
C479 B.n439 VSUBS 0.007647f
C480 B.n440 VSUBS 0.007647f
C481 B.n441 VSUBS 0.007647f
C482 B.n442 VSUBS 0.007647f
C483 B.n443 VSUBS 0.007647f
C484 B.n444 VSUBS 0.007647f
C485 B.n445 VSUBS 0.007647f
C486 B.n446 VSUBS 0.007647f
C487 B.n447 VSUBS 0.007647f
C488 B.n448 VSUBS 0.007647f
C489 B.n449 VSUBS 0.007647f
C490 B.n450 VSUBS 0.007647f
C491 B.n451 VSUBS 0.007647f
C492 B.n452 VSUBS 0.007647f
C493 B.n453 VSUBS 0.007647f
C494 B.n454 VSUBS 0.007647f
C495 B.n455 VSUBS 0.007647f
C496 B.n456 VSUBS 0.007647f
C497 B.n457 VSUBS 0.007647f
C498 B.n458 VSUBS 0.007647f
C499 B.n459 VSUBS 0.007647f
C500 B.n460 VSUBS 0.007647f
C501 B.n461 VSUBS 0.007647f
C502 B.n462 VSUBS 0.007647f
C503 B.n463 VSUBS 0.007647f
C504 B.n464 VSUBS 0.007647f
C505 B.n465 VSUBS 0.007647f
C506 B.n466 VSUBS 0.007647f
C507 B.n467 VSUBS 0.007647f
C508 B.n468 VSUBS 0.007647f
C509 B.n469 VSUBS 0.007647f
C510 B.n470 VSUBS 0.007647f
C511 B.n471 VSUBS 0.007647f
C512 B.n472 VSUBS 0.007647f
C513 B.n473 VSUBS 0.007647f
C514 B.n474 VSUBS 0.007647f
C515 B.n475 VSUBS 0.007647f
C516 B.n476 VSUBS 0.007647f
C517 B.n477 VSUBS 0.007647f
C518 B.n478 VSUBS 0.007647f
C519 B.n479 VSUBS 0.007647f
C520 B.n480 VSUBS 0.007647f
C521 B.n481 VSUBS 0.007197f
C522 B.n482 VSUBS 0.017717f
C523 B.n483 VSUBS 0.004273f
C524 B.n484 VSUBS 0.007647f
C525 B.n485 VSUBS 0.007647f
C526 B.n486 VSUBS 0.007647f
C527 B.n487 VSUBS 0.007647f
C528 B.n488 VSUBS 0.007647f
C529 B.n489 VSUBS 0.007647f
C530 B.n490 VSUBS 0.007647f
C531 B.n491 VSUBS 0.007647f
C532 B.n492 VSUBS 0.007647f
C533 B.n493 VSUBS 0.007647f
C534 B.n494 VSUBS 0.007647f
C535 B.n495 VSUBS 0.007647f
C536 B.n496 VSUBS 0.004273f
C537 B.n497 VSUBS 0.007647f
C538 B.n498 VSUBS 0.007647f
C539 B.n499 VSUBS 0.007197f
C540 B.n500 VSUBS 0.007647f
C541 B.n501 VSUBS 0.007647f
C542 B.n502 VSUBS 0.007647f
C543 B.n503 VSUBS 0.007647f
C544 B.n504 VSUBS 0.007647f
C545 B.n505 VSUBS 0.007647f
C546 B.n506 VSUBS 0.007647f
C547 B.n507 VSUBS 0.007647f
C548 B.n508 VSUBS 0.007647f
C549 B.n509 VSUBS 0.007647f
C550 B.n510 VSUBS 0.007647f
C551 B.n511 VSUBS 0.007647f
C552 B.n512 VSUBS 0.007647f
C553 B.n513 VSUBS 0.007647f
C554 B.n514 VSUBS 0.007647f
C555 B.n515 VSUBS 0.007647f
C556 B.n516 VSUBS 0.007647f
C557 B.n517 VSUBS 0.007647f
C558 B.n518 VSUBS 0.007647f
C559 B.n519 VSUBS 0.007647f
C560 B.n520 VSUBS 0.007647f
C561 B.n521 VSUBS 0.007647f
C562 B.n522 VSUBS 0.007647f
C563 B.n523 VSUBS 0.007647f
C564 B.n524 VSUBS 0.007647f
C565 B.n525 VSUBS 0.007647f
C566 B.n526 VSUBS 0.007647f
C567 B.n527 VSUBS 0.007647f
C568 B.n528 VSUBS 0.007647f
C569 B.n529 VSUBS 0.007647f
C570 B.n530 VSUBS 0.007647f
C571 B.n531 VSUBS 0.007647f
C572 B.n532 VSUBS 0.007647f
C573 B.n533 VSUBS 0.007647f
C574 B.n534 VSUBS 0.007647f
C575 B.n535 VSUBS 0.007647f
C576 B.n536 VSUBS 0.007647f
C577 B.n537 VSUBS 0.007647f
C578 B.n538 VSUBS 0.007647f
C579 B.n539 VSUBS 0.007647f
C580 B.n540 VSUBS 0.007647f
C581 B.n541 VSUBS 0.007647f
C582 B.n542 VSUBS 0.007647f
C583 B.n543 VSUBS 0.007647f
C584 B.n544 VSUBS 0.007647f
C585 B.n545 VSUBS 0.007647f
C586 B.n546 VSUBS 0.007647f
C587 B.n547 VSUBS 0.007647f
C588 B.n548 VSUBS 0.007647f
C589 B.n549 VSUBS 0.007647f
C590 B.n550 VSUBS 0.007647f
C591 B.n551 VSUBS 0.007647f
C592 B.n552 VSUBS 0.007647f
C593 B.n553 VSUBS 0.007647f
C594 B.n554 VSUBS 0.007647f
C595 B.n555 VSUBS 0.007647f
C596 B.n556 VSUBS 0.007647f
C597 B.n557 VSUBS 0.007647f
C598 B.n558 VSUBS 0.007647f
C599 B.n559 VSUBS 0.007647f
C600 B.n560 VSUBS 0.007647f
C601 B.n561 VSUBS 0.007647f
C602 B.n562 VSUBS 0.007647f
C603 B.n563 VSUBS 0.007647f
C604 B.n564 VSUBS 0.007647f
C605 B.n565 VSUBS 0.007647f
C606 B.n566 VSUBS 0.007647f
C607 B.n567 VSUBS 0.007647f
C608 B.n568 VSUBS 0.007647f
C609 B.n569 VSUBS 0.007647f
C610 B.n570 VSUBS 0.007647f
C611 B.n571 VSUBS 0.007647f
C612 B.n572 VSUBS 0.007647f
C613 B.n573 VSUBS 0.007647f
C614 B.n574 VSUBS 0.007647f
C615 B.n575 VSUBS 0.007647f
C616 B.n576 VSUBS 0.007647f
C617 B.n577 VSUBS 0.007647f
C618 B.n578 VSUBS 0.007647f
C619 B.n579 VSUBS 0.007647f
C620 B.n580 VSUBS 0.007647f
C621 B.n581 VSUBS 0.007647f
C622 B.n582 VSUBS 0.007647f
C623 B.n583 VSUBS 0.007647f
C624 B.n584 VSUBS 0.007647f
C625 B.n585 VSUBS 0.007647f
C626 B.n586 VSUBS 0.007647f
C627 B.n587 VSUBS 0.007647f
C628 B.n588 VSUBS 0.007647f
C629 B.n589 VSUBS 0.007647f
C630 B.n590 VSUBS 0.007647f
C631 B.n591 VSUBS 0.018024f
C632 B.n592 VSUBS 0.018024f
C633 B.n593 VSUBS 0.017737f
C634 B.n594 VSUBS 0.007647f
C635 B.n595 VSUBS 0.007647f
C636 B.n596 VSUBS 0.007647f
C637 B.n597 VSUBS 0.007647f
C638 B.n598 VSUBS 0.007647f
C639 B.n599 VSUBS 0.007647f
C640 B.n600 VSUBS 0.007647f
C641 B.n601 VSUBS 0.007647f
C642 B.n602 VSUBS 0.007647f
C643 B.n603 VSUBS 0.007647f
C644 B.n604 VSUBS 0.007647f
C645 B.n605 VSUBS 0.007647f
C646 B.n606 VSUBS 0.007647f
C647 B.n607 VSUBS 0.007647f
C648 B.n608 VSUBS 0.007647f
C649 B.n609 VSUBS 0.007647f
C650 B.n610 VSUBS 0.007647f
C651 B.n611 VSUBS 0.007647f
C652 B.n612 VSUBS 0.007647f
C653 B.n613 VSUBS 0.007647f
C654 B.n614 VSUBS 0.007647f
C655 B.n615 VSUBS 0.007647f
C656 B.n616 VSUBS 0.007647f
C657 B.n617 VSUBS 0.007647f
C658 B.n618 VSUBS 0.007647f
C659 B.n619 VSUBS 0.007647f
C660 B.n620 VSUBS 0.007647f
C661 B.n621 VSUBS 0.007647f
C662 B.n622 VSUBS 0.007647f
C663 B.n623 VSUBS 0.007647f
C664 B.n624 VSUBS 0.007647f
C665 B.n625 VSUBS 0.007647f
C666 B.n626 VSUBS 0.007647f
C667 B.n627 VSUBS 0.007647f
C668 B.n628 VSUBS 0.007647f
C669 B.n629 VSUBS 0.007647f
C670 B.n630 VSUBS 0.007647f
C671 B.n631 VSUBS 0.007647f
C672 B.n632 VSUBS 0.007647f
C673 B.n633 VSUBS 0.007647f
C674 B.n634 VSUBS 0.007647f
C675 B.n635 VSUBS 0.007647f
C676 B.n636 VSUBS 0.007647f
C677 B.n637 VSUBS 0.007647f
C678 B.n638 VSUBS 0.007647f
C679 B.n639 VSUBS 0.007647f
C680 B.n640 VSUBS 0.007647f
C681 B.n641 VSUBS 0.007647f
C682 B.n642 VSUBS 0.007647f
C683 B.n643 VSUBS 0.007647f
C684 B.n644 VSUBS 0.007647f
C685 B.n645 VSUBS 0.007647f
C686 B.n646 VSUBS 0.007647f
C687 B.n647 VSUBS 0.007647f
C688 B.n648 VSUBS 0.007647f
C689 B.n649 VSUBS 0.007647f
C690 B.n650 VSUBS 0.007647f
C691 B.n651 VSUBS 0.007647f
C692 B.n652 VSUBS 0.007647f
C693 B.n653 VSUBS 0.007647f
C694 B.n654 VSUBS 0.007647f
C695 B.n655 VSUBS 0.007647f
C696 B.n656 VSUBS 0.007647f
C697 B.n657 VSUBS 0.007647f
C698 B.n658 VSUBS 0.007647f
C699 B.n659 VSUBS 0.007647f
C700 B.n660 VSUBS 0.007647f
C701 B.n661 VSUBS 0.007647f
C702 B.n662 VSUBS 0.007647f
C703 B.n663 VSUBS 0.007647f
C704 B.n664 VSUBS 0.007647f
C705 B.n665 VSUBS 0.007647f
C706 B.n666 VSUBS 0.007647f
C707 B.n667 VSUBS 0.007647f
C708 B.n668 VSUBS 0.007647f
C709 B.n669 VSUBS 0.007647f
C710 B.n670 VSUBS 0.007647f
C711 B.n671 VSUBS 0.007647f
C712 B.n672 VSUBS 0.007647f
C713 B.n673 VSUBS 0.007647f
C714 B.n674 VSUBS 0.007647f
C715 B.n675 VSUBS 0.007647f
C716 B.n676 VSUBS 0.007647f
C717 B.n677 VSUBS 0.007647f
C718 B.n678 VSUBS 0.007647f
C719 B.n679 VSUBS 0.007647f
C720 B.n680 VSUBS 0.007647f
C721 B.n681 VSUBS 0.007647f
C722 B.n682 VSUBS 0.007647f
C723 B.n683 VSUBS 0.007647f
C724 B.n684 VSUBS 0.007647f
C725 B.n685 VSUBS 0.007647f
C726 B.n686 VSUBS 0.007647f
C727 B.n687 VSUBS 0.007647f
C728 B.n688 VSUBS 0.007647f
C729 B.n689 VSUBS 0.007647f
C730 B.n690 VSUBS 0.007647f
C731 B.n691 VSUBS 0.007647f
C732 B.n692 VSUBS 0.007647f
C733 B.n693 VSUBS 0.007647f
C734 B.n694 VSUBS 0.007647f
C735 B.n695 VSUBS 0.007647f
C736 B.n696 VSUBS 0.007647f
C737 B.n697 VSUBS 0.007647f
C738 B.n698 VSUBS 0.007647f
C739 B.n699 VSUBS 0.007647f
C740 B.n700 VSUBS 0.007647f
C741 B.n701 VSUBS 0.007647f
C742 B.n702 VSUBS 0.007647f
C743 B.n703 VSUBS 0.007647f
C744 B.n704 VSUBS 0.007647f
C745 B.n705 VSUBS 0.007647f
C746 B.n706 VSUBS 0.007647f
C747 B.n707 VSUBS 0.007647f
C748 B.n708 VSUBS 0.007647f
C749 B.n709 VSUBS 0.007647f
C750 B.n710 VSUBS 0.007647f
C751 B.n711 VSUBS 0.007647f
C752 B.n712 VSUBS 0.007647f
C753 B.n713 VSUBS 0.007647f
C754 B.n714 VSUBS 0.007647f
C755 B.n715 VSUBS 0.007647f
C756 B.n716 VSUBS 0.007647f
C757 B.n717 VSUBS 0.007647f
C758 B.n718 VSUBS 0.007647f
C759 B.n719 VSUBS 0.007647f
C760 B.n720 VSUBS 0.007647f
C761 B.n721 VSUBS 0.007647f
C762 B.n722 VSUBS 0.007647f
C763 B.n723 VSUBS 0.007647f
C764 B.n724 VSUBS 0.007647f
C765 B.n725 VSUBS 0.007647f
C766 B.n726 VSUBS 0.007647f
C767 B.n727 VSUBS 0.007647f
C768 B.n728 VSUBS 0.007647f
C769 B.n729 VSUBS 0.007647f
C770 B.n730 VSUBS 0.007647f
C771 B.n731 VSUBS 0.007647f
C772 B.n732 VSUBS 0.007647f
C773 B.n733 VSUBS 0.007647f
C774 B.n734 VSUBS 0.007647f
C775 B.n735 VSUBS 0.007647f
C776 B.n736 VSUBS 0.007647f
C777 B.n737 VSUBS 0.007647f
C778 B.n738 VSUBS 0.007647f
C779 B.n739 VSUBS 0.007647f
C780 B.n740 VSUBS 0.007647f
C781 B.n741 VSUBS 0.007647f
C782 B.n742 VSUBS 0.007647f
C783 B.n743 VSUBS 0.007647f
C784 B.n744 VSUBS 0.007647f
C785 B.n745 VSUBS 0.007647f
C786 B.n746 VSUBS 0.007647f
C787 B.n747 VSUBS 0.007647f
C788 B.n748 VSUBS 0.007647f
C789 B.n749 VSUBS 0.007647f
C790 B.n750 VSUBS 0.007647f
C791 B.n751 VSUBS 0.007647f
C792 B.n752 VSUBS 0.007647f
C793 B.n753 VSUBS 0.007647f
C794 B.n754 VSUBS 0.007647f
C795 B.n755 VSUBS 0.007647f
C796 B.n756 VSUBS 0.007647f
C797 B.n757 VSUBS 0.007647f
C798 B.n758 VSUBS 0.007647f
C799 B.n759 VSUBS 0.007647f
C800 B.n760 VSUBS 0.007647f
C801 B.n761 VSUBS 0.007647f
C802 B.n762 VSUBS 0.007647f
C803 B.n763 VSUBS 0.007647f
C804 B.n764 VSUBS 0.007647f
C805 B.n765 VSUBS 0.007647f
C806 B.n766 VSUBS 0.007647f
C807 B.n767 VSUBS 0.007647f
C808 B.n768 VSUBS 0.007647f
C809 B.n769 VSUBS 0.007647f
C810 B.n770 VSUBS 0.007647f
C811 B.n771 VSUBS 0.007647f
C812 B.n772 VSUBS 0.007647f
C813 B.n773 VSUBS 0.007647f
C814 B.n774 VSUBS 0.007647f
C815 B.n775 VSUBS 0.007647f
C816 B.n776 VSUBS 0.007647f
C817 B.n777 VSUBS 0.007647f
C818 B.n778 VSUBS 0.007647f
C819 B.n779 VSUBS 0.007647f
C820 B.n780 VSUBS 0.007647f
C821 B.n781 VSUBS 0.007647f
C822 B.n782 VSUBS 0.007647f
C823 B.n783 VSUBS 0.007647f
C824 B.n784 VSUBS 0.007647f
C825 B.n785 VSUBS 0.007647f
C826 B.n786 VSUBS 0.007647f
C827 B.n787 VSUBS 0.007647f
C828 B.n788 VSUBS 0.007647f
C829 B.n789 VSUBS 0.007647f
C830 B.n790 VSUBS 0.007647f
C831 B.n791 VSUBS 0.007647f
C832 B.n792 VSUBS 0.007647f
C833 B.n793 VSUBS 0.007647f
C834 B.n794 VSUBS 0.007647f
C835 B.n795 VSUBS 0.007647f
C836 B.n796 VSUBS 0.007647f
C837 B.n797 VSUBS 0.007647f
C838 B.n798 VSUBS 0.007647f
C839 B.n799 VSUBS 0.007647f
C840 B.n800 VSUBS 0.018642f
C841 B.n801 VSUBS 0.017119f
C842 B.n802 VSUBS 0.018024f
C843 B.n803 VSUBS 0.007647f
C844 B.n804 VSUBS 0.007647f
C845 B.n805 VSUBS 0.007647f
C846 B.n806 VSUBS 0.007647f
C847 B.n807 VSUBS 0.007647f
C848 B.n808 VSUBS 0.007647f
C849 B.n809 VSUBS 0.007647f
C850 B.n810 VSUBS 0.007647f
C851 B.n811 VSUBS 0.007647f
C852 B.n812 VSUBS 0.007647f
C853 B.n813 VSUBS 0.007647f
C854 B.n814 VSUBS 0.007647f
C855 B.n815 VSUBS 0.007647f
C856 B.n816 VSUBS 0.007647f
C857 B.n817 VSUBS 0.007647f
C858 B.n818 VSUBS 0.007647f
C859 B.n819 VSUBS 0.007647f
C860 B.n820 VSUBS 0.007647f
C861 B.n821 VSUBS 0.007647f
C862 B.n822 VSUBS 0.007647f
C863 B.n823 VSUBS 0.007647f
C864 B.n824 VSUBS 0.007647f
C865 B.n825 VSUBS 0.007647f
C866 B.n826 VSUBS 0.007647f
C867 B.n827 VSUBS 0.007647f
C868 B.n828 VSUBS 0.007647f
C869 B.n829 VSUBS 0.007647f
C870 B.n830 VSUBS 0.007647f
C871 B.n831 VSUBS 0.007647f
C872 B.n832 VSUBS 0.007647f
C873 B.n833 VSUBS 0.007647f
C874 B.n834 VSUBS 0.007647f
C875 B.n835 VSUBS 0.007647f
C876 B.n836 VSUBS 0.007647f
C877 B.n837 VSUBS 0.007647f
C878 B.n838 VSUBS 0.007647f
C879 B.n839 VSUBS 0.007647f
C880 B.n840 VSUBS 0.007647f
C881 B.n841 VSUBS 0.007647f
C882 B.n842 VSUBS 0.007647f
C883 B.n843 VSUBS 0.007647f
C884 B.n844 VSUBS 0.007647f
C885 B.n845 VSUBS 0.007647f
C886 B.n846 VSUBS 0.007647f
C887 B.n847 VSUBS 0.007647f
C888 B.n848 VSUBS 0.007647f
C889 B.n849 VSUBS 0.007647f
C890 B.n850 VSUBS 0.007647f
C891 B.n851 VSUBS 0.007647f
C892 B.n852 VSUBS 0.007647f
C893 B.n853 VSUBS 0.007647f
C894 B.n854 VSUBS 0.007647f
C895 B.n855 VSUBS 0.007647f
C896 B.n856 VSUBS 0.007647f
C897 B.n857 VSUBS 0.007647f
C898 B.n858 VSUBS 0.007647f
C899 B.n859 VSUBS 0.007647f
C900 B.n860 VSUBS 0.007647f
C901 B.n861 VSUBS 0.007647f
C902 B.n862 VSUBS 0.007647f
C903 B.n863 VSUBS 0.007647f
C904 B.n864 VSUBS 0.007647f
C905 B.n865 VSUBS 0.007647f
C906 B.n866 VSUBS 0.007647f
C907 B.n867 VSUBS 0.007647f
C908 B.n868 VSUBS 0.007647f
C909 B.n869 VSUBS 0.007647f
C910 B.n870 VSUBS 0.007647f
C911 B.n871 VSUBS 0.007647f
C912 B.n872 VSUBS 0.007647f
C913 B.n873 VSUBS 0.007647f
C914 B.n874 VSUBS 0.007647f
C915 B.n875 VSUBS 0.007647f
C916 B.n876 VSUBS 0.007647f
C917 B.n877 VSUBS 0.007647f
C918 B.n878 VSUBS 0.007647f
C919 B.n879 VSUBS 0.007647f
C920 B.n880 VSUBS 0.007647f
C921 B.n881 VSUBS 0.007647f
C922 B.n882 VSUBS 0.007647f
C923 B.n883 VSUBS 0.007647f
C924 B.n884 VSUBS 0.007647f
C925 B.n885 VSUBS 0.007647f
C926 B.n886 VSUBS 0.007647f
C927 B.n887 VSUBS 0.007647f
C928 B.n888 VSUBS 0.007647f
C929 B.n889 VSUBS 0.007647f
C930 B.n890 VSUBS 0.007647f
C931 B.n891 VSUBS 0.007647f
C932 B.n892 VSUBS 0.007647f
C933 B.n893 VSUBS 0.007647f
C934 B.n894 VSUBS 0.007647f
C935 B.n895 VSUBS 0.007197f
C936 B.n896 VSUBS 0.017717f
C937 B.n897 VSUBS 0.004273f
C938 B.n898 VSUBS 0.007647f
C939 B.n899 VSUBS 0.007647f
C940 B.n900 VSUBS 0.007647f
C941 B.n901 VSUBS 0.007647f
C942 B.n902 VSUBS 0.007647f
C943 B.n903 VSUBS 0.007647f
C944 B.n904 VSUBS 0.007647f
C945 B.n905 VSUBS 0.007647f
C946 B.n906 VSUBS 0.007647f
C947 B.n907 VSUBS 0.007647f
C948 B.n908 VSUBS 0.007647f
C949 B.n909 VSUBS 0.007647f
C950 B.n910 VSUBS 0.004273f
C951 B.n911 VSUBS 0.007647f
C952 B.n912 VSUBS 0.007647f
C953 B.n913 VSUBS 0.007197f
C954 B.n914 VSUBS 0.007647f
C955 B.n915 VSUBS 0.007647f
C956 B.n916 VSUBS 0.007647f
C957 B.n917 VSUBS 0.007647f
C958 B.n918 VSUBS 0.007647f
C959 B.n919 VSUBS 0.007647f
C960 B.n920 VSUBS 0.007647f
C961 B.n921 VSUBS 0.007647f
C962 B.n922 VSUBS 0.007647f
C963 B.n923 VSUBS 0.007647f
C964 B.n924 VSUBS 0.007647f
C965 B.n925 VSUBS 0.007647f
C966 B.n926 VSUBS 0.007647f
C967 B.n927 VSUBS 0.007647f
C968 B.n928 VSUBS 0.007647f
C969 B.n929 VSUBS 0.007647f
C970 B.n930 VSUBS 0.007647f
C971 B.n931 VSUBS 0.007647f
C972 B.n932 VSUBS 0.007647f
C973 B.n933 VSUBS 0.007647f
C974 B.n934 VSUBS 0.007647f
C975 B.n935 VSUBS 0.007647f
C976 B.n936 VSUBS 0.007647f
C977 B.n937 VSUBS 0.007647f
C978 B.n938 VSUBS 0.007647f
C979 B.n939 VSUBS 0.007647f
C980 B.n940 VSUBS 0.007647f
C981 B.n941 VSUBS 0.007647f
C982 B.n942 VSUBS 0.007647f
C983 B.n943 VSUBS 0.007647f
C984 B.n944 VSUBS 0.007647f
C985 B.n945 VSUBS 0.007647f
C986 B.n946 VSUBS 0.007647f
C987 B.n947 VSUBS 0.007647f
C988 B.n948 VSUBS 0.007647f
C989 B.n949 VSUBS 0.007647f
C990 B.n950 VSUBS 0.007647f
C991 B.n951 VSUBS 0.007647f
C992 B.n952 VSUBS 0.007647f
C993 B.n953 VSUBS 0.007647f
C994 B.n954 VSUBS 0.007647f
C995 B.n955 VSUBS 0.007647f
C996 B.n956 VSUBS 0.007647f
C997 B.n957 VSUBS 0.007647f
C998 B.n958 VSUBS 0.007647f
C999 B.n959 VSUBS 0.007647f
C1000 B.n960 VSUBS 0.007647f
C1001 B.n961 VSUBS 0.007647f
C1002 B.n962 VSUBS 0.007647f
C1003 B.n963 VSUBS 0.007647f
C1004 B.n964 VSUBS 0.007647f
C1005 B.n965 VSUBS 0.007647f
C1006 B.n966 VSUBS 0.007647f
C1007 B.n967 VSUBS 0.007647f
C1008 B.n968 VSUBS 0.007647f
C1009 B.n969 VSUBS 0.007647f
C1010 B.n970 VSUBS 0.007647f
C1011 B.n971 VSUBS 0.007647f
C1012 B.n972 VSUBS 0.007647f
C1013 B.n973 VSUBS 0.007647f
C1014 B.n974 VSUBS 0.007647f
C1015 B.n975 VSUBS 0.007647f
C1016 B.n976 VSUBS 0.007647f
C1017 B.n977 VSUBS 0.007647f
C1018 B.n978 VSUBS 0.007647f
C1019 B.n979 VSUBS 0.007647f
C1020 B.n980 VSUBS 0.007647f
C1021 B.n981 VSUBS 0.007647f
C1022 B.n982 VSUBS 0.007647f
C1023 B.n983 VSUBS 0.007647f
C1024 B.n984 VSUBS 0.007647f
C1025 B.n985 VSUBS 0.007647f
C1026 B.n986 VSUBS 0.007647f
C1027 B.n987 VSUBS 0.007647f
C1028 B.n988 VSUBS 0.007647f
C1029 B.n989 VSUBS 0.007647f
C1030 B.n990 VSUBS 0.007647f
C1031 B.n991 VSUBS 0.007647f
C1032 B.n992 VSUBS 0.007647f
C1033 B.n993 VSUBS 0.007647f
C1034 B.n994 VSUBS 0.007647f
C1035 B.n995 VSUBS 0.007647f
C1036 B.n996 VSUBS 0.007647f
C1037 B.n997 VSUBS 0.007647f
C1038 B.n998 VSUBS 0.007647f
C1039 B.n999 VSUBS 0.007647f
C1040 B.n1000 VSUBS 0.007647f
C1041 B.n1001 VSUBS 0.007647f
C1042 B.n1002 VSUBS 0.007647f
C1043 B.n1003 VSUBS 0.007647f
C1044 B.n1004 VSUBS 0.007647f
C1045 B.n1005 VSUBS 0.018024f
C1046 B.n1006 VSUBS 0.018024f
C1047 B.n1007 VSUBS 0.017737f
C1048 B.n1008 VSUBS 0.007647f
C1049 B.n1009 VSUBS 0.007647f
C1050 B.n1010 VSUBS 0.007647f
C1051 B.n1011 VSUBS 0.007647f
C1052 B.n1012 VSUBS 0.007647f
C1053 B.n1013 VSUBS 0.007647f
C1054 B.n1014 VSUBS 0.007647f
C1055 B.n1015 VSUBS 0.007647f
C1056 B.n1016 VSUBS 0.007647f
C1057 B.n1017 VSUBS 0.007647f
C1058 B.n1018 VSUBS 0.007647f
C1059 B.n1019 VSUBS 0.007647f
C1060 B.n1020 VSUBS 0.007647f
C1061 B.n1021 VSUBS 0.007647f
C1062 B.n1022 VSUBS 0.007647f
C1063 B.n1023 VSUBS 0.007647f
C1064 B.n1024 VSUBS 0.007647f
C1065 B.n1025 VSUBS 0.007647f
C1066 B.n1026 VSUBS 0.007647f
C1067 B.n1027 VSUBS 0.007647f
C1068 B.n1028 VSUBS 0.007647f
C1069 B.n1029 VSUBS 0.007647f
C1070 B.n1030 VSUBS 0.007647f
C1071 B.n1031 VSUBS 0.007647f
C1072 B.n1032 VSUBS 0.007647f
C1073 B.n1033 VSUBS 0.007647f
C1074 B.n1034 VSUBS 0.007647f
C1075 B.n1035 VSUBS 0.007647f
C1076 B.n1036 VSUBS 0.007647f
C1077 B.n1037 VSUBS 0.007647f
C1078 B.n1038 VSUBS 0.007647f
C1079 B.n1039 VSUBS 0.007647f
C1080 B.n1040 VSUBS 0.007647f
C1081 B.n1041 VSUBS 0.007647f
C1082 B.n1042 VSUBS 0.007647f
C1083 B.n1043 VSUBS 0.007647f
C1084 B.n1044 VSUBS 0.007647f
C1085 B.n1045 VSUBS 0.007647f
C1086 B.n1046 VSUBS 0.007647f
C1087 B.n1047 VSUBS 0.007647f
C1088 B.n1048 VSUBS 0.007647f
C1089 B.n1049 VSUBS 0.007647f
C1090 B.n1050 VSUBS 0.007647f
C1091 B.n1051 VSUBS 0.007647f
C1092 B.n1052 VSUBS 0.007647f
C1093 B.n1053 VSUBS 0.007647f
C1094 B.n1054 VSUBS 0.007647f
C1095 B.n1055 VSUBS 0.007647f
C1096 B.n1056 VSUBS 0.007647f
C1097 B.n1057 VSUBS 0.007647f
C1098 B.n1058 VSUBS 0.007647f
C1099 B.n1059 VSUBS 0.007647f
C1100 B.n1060 VSUBS 0.007647f
C1101 B.n1061 VSUBS 0.007647f
C1102 B.n1062 VSUBS 0.007647f
C1103 B.n1063 VSUBS 0.007647f
C1104 B.n1064 VSUBS 0.007647f
C1105 B.n1065 VSUBS 0.007647f
C1106 B.n1066 VSUBS 0.007647f
C1107 B.n1067 VSUBS 0.007647f
C1108 B.n1068 VSUBS 0.007647f
C1109 B.n1069 VSUBS 0.007647f
C1110 B.n1070 VSUBS 0.007647f
C1111 B.n1071 VSUBS 0.007647f
C1112 B.n1072 VSUBS 0.007647f
C1113 B.n1073 VSUBS 0.007647f
C1114 B.n1074 VSUBS 0.007647f
C1115 B.n1075 VSUBS 0.007647f
C1116 B.n1076 VSUBS 0.007647f
C1117 B.n1077 VSUBS 0.007647f
C1118 B.n1078 VSUBS 0.007647f
C1119 B.n1079 VSUBS 0.007647f
C1120 B.n1080 VSUBS 0.007647f
C1121 B.n1081 VSUBS 0.007647f
C1122 B.n1082 VSUBS 0.007647f
C1123 B.n1083 VSUBS 0.007647f
C1124 B.n1084 VSUBS 0.007647f
C1125 B.n1085 VSUBS 0.007647f
C1126 B.n1086 VSUBS 0.007647f
C1127 B.n1087 VSUBS 0.007647f
C1128 B.n1088 VSUBS 0.007647f
C1129 B.n1089 VSUBS 0.007647f
C1130 B.n1090 VSUBS 0.007647f
C1131 B.n1091 VSUBS 0.007647f
C1132 B.n1092 VSUBS 0.007647f
C1133 B.n1093 VSUBS 0.007647f
C1134 B.n1094 VSUBS 0.007647f
C1135 B.n1095 VSUBS 0.007647f
C1136 B.n1096 VSUBS 0.007647f
C1137 B.n1097 VSUBS 0.007647f
C1138 B.n1098 VSUBS 0.007647f
C1139 B.n1099 VSUBS 0.007647f
C1140 B.n1100 VSUBS 0.007647f
C1141 B.n1101 VSUBS 0.007647f
C1142 B.n1102 VSUBS 0.007647f
C1143 B.n1103 VSUBS 0.007647f
C1144 B.n1104 VSUBS 0.007647f
C1145 B.n1105 VSUBS 0.007647f
C1146 B.n1106 VSUBS 0.007647f
C1147 B.n1107 VSUBS 0.007647f
C1148 B.n1108 VSUBS 0.007647f
C1149 B.n1109 VSUBS 0.007647f
C1150 B.n1110 VSUBS 0.007647f
C1151 B.n1111 VSUBS 0.017315f
C1152 VDD2.n0 VSUBS 0.029678f
C1153 VDD2.n1 VSUBS 0.028396f
C1154 VDD2.n2 VSUBS 0.015258f
C1155 VDD2.n3 VSUBS 0.036066f
C1156 VDD2.n4 VSUBS 0.016156f
C1157 VDD2.n5 VSUBS 0.028396f
C1158 VDD2.n6 VSUBS 0.015258f
C1159 VDD2.n7 VSUBS 0.036066f
C1160 VDD2.n8 VSUBS 0.016156f
C1161 VDD2.n9 VSUBS 0.028396f
C1162 VDD2.n10 VSUBS 0.015258f
C1163 VDD2.n11 VSUBS 0.036066f
C1164 VDD2.n12 VSUBS 0.016156f
C1165 VDD2.n13 VSUBS 0.028396f
C1166 VDD2.n14 VSUBS 0.015258f
C1167 VDD2.n15 VSUBS 0.036066f
C1168 VDD2.n16 VSUBS 0.016156f
C1169 VDD2.n17 VSUBS 0.028396f
C1170 VDD2.n18 VSUBS 0.015258f
C1171 VDD2.n19 VSUBS 0.036066f
C1172 VDD2.n20 VSUBS 0.016156f
C1173 VDD2.n21 VSUBS 0.028396f
C1174 VDD2.n22 VSUBS 0.015258f
C1175 VDD2.n23 VSUBS 0.036066f
C1176 VDD2.n24 VSUBS 0.016156f
C1177 VDD2.n25 VSUBS 0.028396f
C1178 VDD2.n26 VSUBS 0.015258f
C1179 VDD2.n27 VSUBS 0.036066f
C1180 VDD2.n28 VSUBS 0.016156f
C1181 VDD2.n29 VSUBS 0.028396f
C1182 VDD2.n30 VSUBS 0.015258f
C1183 VDD2.n31 VSUBS 0.036066f
C1184 VDD2.n32 VSUBS 0.016156f
C1185 VDD2.n33 VSUBS 0.318771f
C1186 VDD2.t9 VSUBS 0.078428f
C1187 VDD2.n34 VSUBS 0.027049f
C1188 VDD2.n35 VSUBS 0.02713f
C1189 VDD2.n36 VSUBS 0.015258f
C1190 VDD2.n37 VSUBS 2.31711f
C1191 VDD2.n38 VSUBS 0.028396f
C1192 VDD2.n39 VSUBS 0.015258f
C1193 VDD2.n40 VSUBS 0.016156f
C1194 VDD2.n41 VSUBS 0.036066f
C1195 VDD2.n42 VSUBS 0.036066f
C1196 VDD2.n43 VSUBS 0.016156f
C1197 VDD2.n44 VSUBS 0.015258f
C1198 VDD2.n45 VSUBS 0.028396f
C1199 VDD2.n46 VSUBS 0.028396f
C1200 VDD2.n47 VSUBS 0.015258f
C1201 VDD2.n48 VSUBS 0.016156f
C1202 VDD2.n49 VSUBS 0.036066f
C1203 VDD2.n50 VSUBS 0.036066f
C1204 VDD2.n51 VSUBS 0.036066f
C1205 VDD2.n52 VSUBS 0.016156f
C1206 VDD2.n53 VSUBS 0.015258f
C1207 VDD2.n54 VSUBS 0.028396f
C1208 VDD2.n55 VSUBS 0.028396f
C1209 VDD2.n56 VSUBS 0.015258f
C1210 VDD2.n57 VSUBS 0.015707f
C1211 VDD2.n58 VSUBS 0.015707f
C1212 VDD2.n59 VSUBS 0.036066f
C1213 VDD2.n60 VSUBS 0.036066f
C1214 VDD2.n61 VSUBS 0.016156f
C1215 VDD2.n62 VSUBS 0.015258f
C1216 VDD2.n63 VSUBS 0.028396f
C1217 VDD2.n64 VSUBS 0.028396f
C1218 VDD2.n65 VSUBS 0.015258f
C1219 VDD2.n66 VSUBS 0.016156f
C1220 VDD2.n67 VSUBS 0.036066f
C1221 VDD2.n68 VSUBS 0.036066f
C1222 VDD2.n69 VSUBS 0.016156f
C1223 VDD2.n70 VSUBS 0.015258f
C1224 VDD2.n71 VSUBS 0.028396f
C1225 VDD2.n72 VSUBS 0.028396f
C1226 VDD2.n73 VSUBS 0.015258f
C1227 VDD2.n74 VSUBS 0.016156f
C1228 VDD2.n75 VSUBS 0.036066f
C1229 VDD2.n76 VSUBS 0.036066f
C1230 VDD2.n77 VSUBS 0.016156f
C1231 VDD2.n78 VSUBS 0.015258f
C1232 VDD2.n79 VSUBS 0.028396f
C1233 VDD2.n80 VSUBS 0.028396f
C1234 VDD2.n81 VSUBS 0.015258f
C1235 VDD2.n82 VSUBS 0.016156f
C1236 VDD2.n83 VSUBS 0.036066f
C1237 VDD2.n84 VSUBS 0.036066f
C1238 VDD2.n85 VSUBS 0.016156f
C1239 VDD2.n86 VSUBS 0.015258f
C1240 VDD2.n87 VSUBS 0.028396f
C1241 VDD2.n88 VSUBS 0.028396f
C1242 VDD2.n89 VSUBS 0.015258f
C1243 VDD2.n90 VSUBS 0.016156f
C1244 VDD2.n91 VSUBS 0.036066f
C1245 VDD2.n92 VSUBS 0.036066f
C1246 VDD2.n93 VSUBS 0.016156f
C1247 VDD2.n94 VSUBS 0.015258f
C1248 VDD2.n95 VSUBS 0.028396f
C1249 VDD2.n96 VSUBS 0.028396f
C1250 VDD2.n97 VSUBS 0.015258f
C1251 VDD2.n98 VSUBS 0.016156f
C1252 VDD2.n99 VSUBS 0.036066f
C1253 VDD2.n100 VSUBS 0.087923f
C1254 VDD2.n101 VSUBS 0.016156f
C1255 VDD2.n102 VSUBS 0.029964f
C1256 VDD2.n103 VSUBS 0.069126f
C1257 VDD2.n104 VSUBS 0.104193f
C1258 VDD2.t5 VSUBS 0.435542f
C1259 VDD2.t3 VSUBS 0.435542f
C1260 VDD2.n105 VSUBS 3.66804f
C1261 VDD2.n106 VSUBS 1.19338f
C1262 VDD2.t1 VSUBS 0.435542f
C1263 VDD2.t0 VSUBS 0.435542f
C1264 VDD2.n107 VSUBS 3.69917f
C1265 VDD2.n108 VSUBS 4.43943f
C1266 VDD2.n109 VSUBS 0.029678f
C1267 VDD2.n110 VSUBS 0.028396f
C1268 VDD2.n111 VSUBS 0.015258f
C1269 VDD2.n112 VSUBS 0.036066f
C1270 VDD2.n113 VSUBS 0.016156f
C1271 VDD2.n114 VSUBS 0.028396f
C1272 VDD2.n115 VSUBS 0.015258f
C1273 VDD2.n116 VSUBS 0.036066f
C1274 VDD2.n117 VSUBS 0.016156f
C1275 VDD2.n118 VSUBS 0.028396f
C1276 VDD2.n119 VSUBS 0.015258f
C1277 VDD2.n120 VSUBS 0.036066f
C1278 VDD2.n121 VSUBS 0.016156f
C1279 VDD2.n122 VSUBS 0.028396f
C1280 VDD2.n123 VSUBS 0.015258f
C1281 VDD2.n124 VSUBS 0.036066f
C1282 VDD2.n125 VSUBS 0.016156f
C1283 VDD2.n126 VSUBS 0.028396f
C1284 VDD2.n127 VSUBS 0.015258f
C1285 VDD2.n128 VSUBS 0.036066f
C1286 VDD2.n129 VSUBS 0.016156f
C1287 VDD2.n130 VSUBS 0.028396f
C1288 VDD2.n131 VSUBS 0.015258f
C1289 VDD2.n132 VSUBS 0.036066f
C1290 VDD2.n133 VSUBS 0.016156f
C1291 VDD2.n134 VSUBS 0.028396f
C1292 VDD2.n135 VSUBS 0.015258f
C1293 VDD2.n136 VSUBS 0.036066f
C1294 VDD2.n137 VSUBS 0.036066f
C1295 VDD2.n138 VSUBS 0.016156f
C1296 VDD2.n139 VSUBS 0.028396f
C1297 VDD2.n140 VSUBS 0.015258f
C1298 VDD2.n141 VSUBS 0.036066f
C1299 VDD2.n142 VSUBS 0.016156f
C1300 VDD2.n143 VSUBS 0.318771f
C1301 VDD2.t6 VSUBS 0.078428f
C1302 VDD2.n144 VSUBS 0.027049f
C1303 VDD2.n145 VSUBS 0.02713f
C1304 VDD2.n146 VSUBS 0.015258f
C1305 VDD2.n147 VSUBS 2.31711f
C1306 VDD2.n148 VSUBS 0.028396f
C1307 VDD2.n149 VSUBS 0.015258f
C1308 VDD2.n150 VSUBS 0.016156f
C1309 VDD2.n151 VSUBS 0.036066f
C1310 VDD2.n152 VSUBS 0.036066f
C1311 VDD2.n153 VSUBS 0.016156f
C1312 VDD2.n154 VSUBS 0.015258f
C1313 VDD2.n155 VSUBS 0.028396f
C1314 VDD2.n156 VSUBS 0.028396f
C1315 VDD2.n157 VSUBS 0.015258f
C1316 VDD2.n158 VSUBS 0.016156f
C1317 VDD2.n159 VSUBS 0.036066f
C1318 VDD2.n160 VSUBS 0.036066f
C1319 VDD2.n161 VSUBS 0.016156f
C1320 VDD2.n162 VSUBS 0.015258f
C1321 VDD2.n163 VSUBS 0.028396f
C1322 VDD2.n164 VSUBS 0.028396f
C1323 VDD2.n165 VSUBS 0.015258f
C1324 VDD2.n166 VSUBS 0.015707f
C1325 VDD2.n167 VSUBS 0.015707f
C1326 VDD2.n168 VSUBS 0.036066f
C1327 VDD2.n169 VSUBS 0.036066f
C1328 VDD2.n170 VSUBS 0.016156f
C1329 VDD2.n171 VSUBS 0.015258f
C1330 VDD2.n172 VSUBS 0.028396f
C1331 VDD2.n173 VSUBS 0.028396f
C1332 VDD2.n174 VSUBS 0.015258f
C1333 VDD2.n175 VSUBS 0.016156f
C1334 VDD2.n176 VSUBS 0.036066f
C1335 VDD2.n177 VSUBS 0.036066f
C1336 VDD2.n178 VSUBS 0.016156f
C1337 VDD2.n179 VSUBS 0.015258f
C1338 VDD2.n180 VSUBS 0.028396f
C1339 VDD2.n181 VSUBS 0.028396f
C1340 VDD2.n182 VSUBS 0.015258f
C1341 VDD2.n183 VSUBS 0.016156f
C1342 VDD2.n184 VSUBS 0.036066f
C1343 VDD2.n185 VSUBS 0.036066f
C1344 VDD2.n186 VSUBS 0.016156f
C1345 VDD2.n187 VSUBS 0.015258f
C1346 VDD2.n188 VSUBS 0.028396f
C1347 VDD2.n189 VSUBS 0.028396f
C1348 VDD2.n190 VSUBS 0.015258f
C1349 VDD2.n191 VSUBS 0.016156f
C1350 VDD2.n192 VSUBS 0.036066f
C1351 VDD2.n193 VSUBS 0.036066f
C1352 VDD2.n194 VSUBS 0.016156f
C1353 VDD2.n195 VSUBS 0.015258f
C1354 VDD2.n196 VSUBS 0.028396f
C1355 VDD2.n197 VSUBS 0.028396f
C1356 VDD2.n198 VSUBS 0.015258f
C1357 VDD2.n199 VSUBS 0.016156f
C1358 VDD2.n200 VSUBS 0.036066f
C1359 VDD2.n201 VSUBS 0.036066f
C1360 VDD2.n202 VSUBS 0.016156f
C1361 VDD2.n203 VSUBS 0.015258f
C1362 VDD2.n204 VSUBS 0.028396f
C1363 VDD2.n205 VSUBS 0.028396f
C1364 VDD2.n206 VSUBS 0.015258f
C1365 VDD2.n207 VSUBS 0.016156f
C1366 VDD2.n208 VSUBS 0.036066f
C1367 VDD2.n209 VSUBS 0.087923f
C1368 VDD2.n210 VSUBS 0.016156f
C1369 VDD2.n211 VSUBS 0.029964f
C1370 VDD2.n212 VSUBS 0.069126f
C1371 VDD2.n213 VSUBS 0.086037f
C1372 VDD2.n214 VSUBS 4.1495f
C1373 VDD2.t2 VSUBS 0.435542f
C1374 VDD2.t8 VSUBS 0.435542f
C1375 VDD2.n215 VSUBS 3.66806f
C1376 VDD2.n216 VSUBS 0.892933f
C1377 VDD2.t7 VSUBS 0.435542f
C1378 VDD2.t4 VSUBS 0.435542f
C1379 VDD2.n217 VSUBS 3.69912f
C1380 VN.t9 VSUBS 3.71849f
C1381 VN.n0 VSUBS 1.37078f
C1382 VN.n1 VSUBS 0.022365f
C1383 VN.n2 VSUBS 0.026703f
C1384 VN.n3 VSUBS 0.022365f
C1385 VN.t8 VSUBS 3.71849f
C1386 VN.n4 VSUBS 1.28174f
C1387 VN.n5 VSUBS 0.022365f
C1388 VN.n6 VSUBS 0.030779f
C1389 VN.n7 VSUBS 0.022365f
C1390 VN.t6 VSUBS 3.71849f
C1391 VN.n8 VSUBS 0.041682f
C1392 VN.n9 VSUBS 0.022365f
C1393 VN.n10 VSUBS 0.041682f
C1394 VN.t0 VSUBS 3.97982f
C1395 VN.n11 VSUBS 1.31003f
C1396 VN.t4 VSUBS 3.71849f
C1397 VN.n12 VSUBS 1.36253f
C1398 VN.n13 VSUBS 0.039213f
C1399 VN.n14 VSUBS 0.256001f
C1400 VN.n15 VSUBS 0.022365f
C1401 VN.n16 VSUBS 0.022365f
C1402 VN.n17 VSUBS 0.034518f
C1403 VN.n18 VSUBS 0.030779f
C1404 VN.n19 VSUBS 0.041682f
C1405 VN.n20 VSUBS 0.022365f
C1406 VN.n21 VSUBS 0.022365f
C1407 VN.n22 VSUBS 0.022365f
C1408 VN.n23 VSUBS 1.30284f
C1409 VN.n24 VSUBS 0.041682f
C1410 VN.n25 VSUBS 0.041682f
C1411 VN.n26 VSUBS 0.022365f
C1412 VN.n27 VSUBS 0.022365f
C1413 VN.n28 VSUBS 0.022365f
C1414 VN.n29 VSUBS 0.034518f
C1415 VN.n30 VSUBS 0.041682f
C1416 VN.n31 VSUBS 0.039213f
C1417 VN.n32 VSUBS 0.022365f
C1418 VN.n33 VSUBS 0.022365f
C1419 VN.n34 VSUBS 0.023573f
C1420 VN.n35 VSUBS 0.041682f
C1421 VN.n36 VSUBS 0.042074f
C1422 VN.n37 VSUBS 0.022365f
C1423 VN.n38 VSUBS 0.022365f
C1424 VN.n39 VSUBS 0.022365f
C1425 VN.n40 VSUBS 0.038202f
C1426 VN.n41 VSUBS 0.041682f
C1427 VN.n42 VSUBS 0.036743f
C1428 VN.n43 VSUBS 0.036096f
C1429 VN.n44 VSUBS 0.048792f
C1430 VN.t3 VSUBS 3.71849f
C1431 VN.n45 VSUBS 1.37078f
C1432 VN.n46 VSUBS 0.022365f
C1433 VN.n47 VSUBS 0.026703f
C1434 VN.n48 VSUBS 0.022365f
C1435 VN.t7 VSUBS 3.71849f
C1436 VN.n49 VSUBS 1.28174f
C1437 VN.n50 VSUBS 0.022365f
C1438 VN.n51 VSUBS 0.030779f
C1439 VN.n52 VSUBS 0.022365f
C1440 VN.t1 VSUBS 3.71849f
C1441 VN.n53 VSUBS 0.041682f
C1442 VN.n54 VSUBS 0.022365f
C1443 VN.n55 VSUBS 0.041682f
C1444 VN.t5 VSUBS 3.97982f
C1445 VN.n56 VSUBS 1.31003f
C1446 VN.t2 VSUBS 3.71849f
C1447 VN.n57 VSUBS 1.36253f
C1448 VN.n58 VSUBS 0.039213f
C1449 VN.n59 VSUBS 0.256001f
C1450 VN.n60 VSUBS 0.022365f
C1451 VN.n61 VSUBS 0.022365f
C1452 VN.n62 VSUBS 0.034518f
C1453 VN.n63 VSUBS 0.030779f
C1454 VN.n64 VSUBS 0.041682f
C1455 VN.n65 VSUBS 0.022365f
C1456 VN.n66 VSUBS 0.022365f
C1457 VN.n67 VSUBS 0.022365f
C1458 VN.n68 VSUBS 1.30284f
C1459 VN.n69 VSUBS 0.041682f
C1460 VN.n70 VSUBS 0.041682f
C1461 VN.n71 VSUBS 0.022365f
C1462 VN.n72 VSUBS 0.022365f
C1463 VN.n73 VSUBS 0.022365f
C1464 VN.n74 VSUBS 0.034518f
C1465 VN.n75 VSUBS 0.041682f
C1466 VN.n76 VSUBS 0.039213f
C1467 VN.n77 VSUBS 0.022365f
C1468 VN.n78 VSUBS 0.022365f
C1469 VN.n79 VSUBS 0.023573f
C1470 VN.n80 VSUBS 0.041682f
C1471 VN.n81 VSUBS 0.042074f
C1472 VN.n82 VSUBS 0.022365f
C1473 VN.n83 VSUBS 0.022365f
C1474 VN.n84 VSUBS 0.022365f
C1475 VN.n85 VSUBS 0.038202f
C1476 VN.n86 VSUBS 0.041682f
C1477 VN.n87 VSUBS 0.036743f
C1478 VN.n88 VSUBS 0.036096f
C1479 VN.n89 VSUBS 1.70018f
C1480 VDD1.n0 VSUBS 0.029675f
C1481 VDD1.n1 VSUBS 0.028392f
C1482 VDD1.n2 VSUBS 0.015257f
C1483 VDD1.n3 VSUBS 0.036061f
C1484 VDD1.n4 VSUBS 0.016154f
C1485 VDD1.n5 VSUBS 0.028392f
C1486 VDD1.n6 VSUBS 0.015257f
C1487 VDD1.n7 VSUBS 0.036061f
C1488 VDD1.n8 VSUBS 0.016154f
C1489 VDD1.n9 VSUBS 0.028392f
C1490 VDD1.n10 VSUBS 0.015257f
C1491 VDD1.n11 VSUBS 0.036061f
C1492 VDD1.n12 VSUBS 0.016154f
C1493 VDD1.n13 VSUBS 0.028392f
C1494 VDD1.n14 VSUBS 0.015257f
C1495 VDD1.n15 VSUBS 0.036061f
C1496 VDD1.n16 VSUBS 0.016154f
C1497 VDD1.n17 VSUBS 0.028392f
C1498 VDD1.n18 VSUBS 0.015257f
C1499 VDD1.n19 VSUBS 0.036061f
C1500 VDD1.n20 VSUBS 0.016154f
C1501 VDD1.n21 VSUBS 0.028392f
C1502 VDD1.n22 VSUBS 0.015257f
C1503 VDD1.n23 VSUBS 0.036061f
C1504 VDD1.n24 VSUBS 0.016154f
C1505 VDD1.n25 VSUBS 0.028392f
C1506 VDD1.n26 VSUBS 0.015257f
C1507 VDD1.n27 VSUBS 0.036061f
C1508 VDD1.n28 VSUBS 0.036061f
C1509 VDD1.n29 VSUBS 0.016154f
C1510 VDD1.n30 VSUBS 0.028392f
C1511 VDD1.n31 VSUBS 0.015257f
C1512 VDD1.n32 VSUBS 0.036061f
C1513 VDD1.n33 VSUBS 0.016154f
C1514 VDD1.n34 VSUBS 0.318733f
C1515 VDD1.t7 VSUBS 0.078419f
C1516 VDD1.n35 VSUBS 0.027046f
C1517 VDD1.n36 VSUBS 0.027127f
C1518 VDD1.n37 VSUBS 0.015257f
C1519 VDD1.n38 VSUBS 2.31683f
C1520 VDD1.n39 VSUBS 0.028392f
C1521 VDD1.n40 VSUBS 0.015257f
C1522 VDD1.n41 VSUBS 0.016154f
C1523 VDD1.n42 VSUBS 0.036061f
C1524 VDD1.n43 VSUBS 0.036061f
C1525 VDD1.n44 VSUBS 0.016154f
C1526 VDD1.n45 VSUBS 0.015257f
C1527 VDD1.n46 VSUBS 0.028392f
C1528 VDD1.n47 VSUBS 0.028392f
C1529 VDD1.n48 VSUBS 0.015257f
C1530 VDD1.n49 VSUBS 0.016154f
C1531 VDD1.n50 VSUBS 0.036061f
C1532 VDD1.n51 VSUBS 0.036061f
C1533 VDD1.n52 VSUBS 0.016154f
C1534 VDD1.n53 VSUBS 0.015257f
C1535 VDD1.n54 VSUBS 0.028392f
C1536 VDD1.n55 VSUBS 0.028392f
C1537 VDD1.n56 VSUBS 0.015257f
C1538 VDD1.n57 VSUBS 0.015705f
C1539 VDD1.n58 VSUBS 0.015705f
C1540 VDD1.n59 VSUBS 0.036061f
C1541 VDD1.n60 VSUBS 0.036061f
C1542 VDD1.n61 VSUBS 0.016154f
C1543 VDD1.n62 VSUBS 0.015257f
C1544 VDD1.n63 VSUBS 0.028392f
C1545 VDD1.n64 VSUBS 0.028392f
C1546 VDD1.n65 VSUBS 0.015257f
C1547 VDD1.n66 VSUBS 0.016154f
C1548 VDD1.n67 VSUBS 0.036061f
C1549 VDD1.n68 VSUBS 0.036061f
C1550 VDD1.n69 VSUBS 0.016154f
C1551 VDD1.n70 VSUBS 0.015257f
C1552 VDD1.n71 VSUBS 0.028392f
C1553 VDD1.n72 VSUBS 0.028392f
C1554 VDD1.n73 VSUBS 0.015257f
C1555 VDD1.n74 VSUBS 0.016154f
C1556 VDD1.n75 VSUBS 0.036061f
C1557 VDD1.n76 VSUBS 0.036061f
C1558 VDD1.n77 VSUBS 0.016154f
C1559 VDD1.n78 VSUBS 0.015257f
C1560 VDD1.n79 VSUBS 0.028392f
C1561 VDD1.n80 VSUBS 0.028392f
C1562 VDD1.n81 VSUBS 0.015257f
C1563 VDD1.n82 VSUBS 0.016154f
C1564 VDD1.n83 VSUBS 0.036061f
C1565 VDD1.n84 VSUBS 0.036061f
C1566 VDD1.n85 VSUBS 0.016154f
C1567 VDD1.n86 VSUBS 0.015257f
C1568 VDD1.n87 VSUBS 0.028392f
C1569 VDD1.n88 VSUBS 0.028392f
C1570 VDD1.n89 VSUBS 0.015257f
C1571 VDD1.n90 VSUBS 0.016154f
C1572 VDD1.n91 VSUBS 0.036061f
C1573 VDD1.n92 VSUBS 0.036061f
C1574 VDD1.n93 VSUBS 0.016154f
C1575 VDD1.n94 VSUBS 0.015257f
C1576 VDD1.n95 VSUBS 0.028392f
C1577 VDD1.n96 VSUBS 0.028392f
C1578 VDD1.n97 VSUBS 0.015257f
C1579 VDD1.n98 VSUBS 0.016154f
C1580 VDD1.n99 VSUBS 0.036061f
C1581 VDD1.n100 VSUBS 0.087913f
C1582 VDD1.n101 VSUBS 0.016154f
C1583 VDD1.n102 VSUBS 0.029961f
C1584 VDD1.n103 VSUBS 0.069118f
C1585 VDD1.n104 VSUBS 0.104181f
C1586 VDD1.t8 VSUBS 0.43549f
C1587 VDD1.t3 VSUBS 0.43549f
C1588 VDD1.n105 VSUBS 3.66762f
C1589 VDD1.n106 VSUBS 1.20265f
C1590 VDD1.n107 VSUBS 0.029675f
C1591 VDD1.n108 VSUBS 0.028392f
C1592 VDD1.n109 VSUBS 0.015257f
C1593 VDD1.n110 VSUBS 0.036061f
C1594 VDD1.n111 VSUBS 0.016154f
C1595 VDD1.n112 VSUBS 0.028392f
C1596 VDD1.n113 VSUBS 0.015257f
C1597 VDD1.n114 VSUBS 0.036061f
C1598 VDD1.n115 VSUBS 0.016154f
C1599 VDD1.n116 VSUBS 0.028392f
C1600 VDD1.n117 VSUBS 0.015257f
C1601 VDD1.n118 VSUBS 0.036061f
C1602 VDD1.n119 VSUBS 0.016154f
C1603 VDD1.n120 VSUBS 0.028392f
C1604 VDD1.n121 VSUBS 0.015257f
C1605 VDD1.n122 VSUBS 0.036061f
C1606 VDD1.n123 VSUBS 0.016154f
C1607 VDD1.n124 VSUBS 0.028392f
C1608 VDD1.n125 VSUBS 0.015257f
C1609 VDD1.n126 VSUBS 0.036061f
C1610 VDD1.n127 VSUBS 0.016154f
C1611 VDD1.n128 VSUBS 0.028392f
C1612 VDD1.n129 VSUBS 0.015257f
C1613 VDD1.n130 VSUBS 0.036061f
C1614 VDD1.n131 VSUBS 0.016154f
C1615 VDD1.n132 VSUBS 0.028392f
C1616 VDD1.n133 VSUBS 0.015257f
C1617 VDD1.n134 VSUBS 0.036061f
C1618 VDD1.n135 VSUBS 0.016154f
C1619 VDD1.n136 VSUBS 0.028392f
C1620 VDD1.n137 VSUBS 0.015257f
C1621 VDD1.n138 VSUBS 0.036061f
C1622 VDD1.n139 VSUBS 0.016154f
C1623 VDD1.n140 VSUBS 0.318733f
C1624 VDD1.t2 VSUBS 0.078419f
C1625 VDD1.n141 VSUBS 0.027046f
C1626 VDD1.n142 VSUBS 0.027127f
C1627 VDD1.n143 VSUBS 0.015257f
C1628 VDD1.n144 VSUBS 2.31683f
C1629 VDD1.n145 VSUBS 0.028392f
C1630 VDD1.n146 VSUBS 0.015257f
C1631 VDD1.n147 VSUBS 0.016154f
C1632 VDD1.n148 VSUBS 0.036061f
C1633 VDD1.n149 VSUBS 0.036061f
C1634 VDD1.n150 VSUBS 0.016154f
C1635 VDD1.n151 VSUBS 0.015257f
C1636 VDD1.n152 VSUBS 0.028392f
C1637 VDD1.n153 VSUBS 0.028392f
C1638 VDD1.n154 VSUBS 0.015257f
C1639 VDD1.n155 VSUBS 0.016154f
C1640 VDD1.n156 VSUBS 0.036061f
C1641 VDD1.n157 VSUBS 0.036061f
C1642 VDD1.n158 VSUBS 0.036061f
C1643 VDD1.n159 VSUBS 0.016154f
C1644 VDD1.n160 VSUBS 0.015257f
C1645 VDD1.n161 VSUBS 0.028392f
C1646 VDD1.n162 VSUBS 0.028392f
C1647 VDD1.n163 VSUBS 0.015257f
C1648 VDD1.n164 VSUBS 0.015705f
C1649 VDD1.n165 VSUBS 0.015705f
C1650 VDD1.n166 VSUBS 0.036061f
C1651 VDD1.n167 VSUBS 0.036061f
C1652 VDD1.n168 VSUBS 0.016154f
C1653 VDD1.n169 VSUBS 0.015257f
C1654 VDD1.n170 VSUBS 0.028392f
C1655 VDD1.n171 VSUBS 0.028392f
C1656 VDD1.n172 VSUBS 0.015257f
C1657 VDD1.n173 VSUBS 0.016154f
C1658 VDD1.n174 VSUBS 0.036061f
C1659 VDD1.n175 VSUBS 0.036061f
C1660 VDD1.n176 VSUBS 0.016154f
C1661 VDD1.n177 VSUBS 0.015257f
C1662 VDD1.n178 VSUBS 0.028392f
C1663 VDD1.n179 VSUBS 0.028392f
C1664 VDD1.n180 VSUBS 0.015257f
C1665 VDD1.n181 VSUBS 0.016154f
C1666 VDD1.n182 VSUBS 0.036061f
C1667 VDD1.n183 VSUBS 0.036061f
C1668 VDD1.n184 VSUBS 0.016154f
C1669 VDD1.n185 VSUBS 0.015257f
C1670 VDD1.n186 VSUBS 0.028392f
C1671 VDD1.n187 VSUBS 0.028392f
C1672 VDD1.n188 VSUBS 0.015257f
C1673 VDD1.n189 VSUBS 0.016154f
C1674 VDD1.n190 VSUBS 0.036061f
C1675 VDD1.n191 VSUBS 0.036061f
C1676 VDD1.n192 VSUBS 0.016154f
C1677 VDD1.n193 VSUBS 0.015257f
C1678 VDD1.n194 VSUBS 0.028392f
C1679 VDD1.n195 VSUBS 0.028392f
C1680 VDD1.n196 VSUBS 0.015257f
C1681 VDD1.n197 VSUBS 0.016154f
C1682 VDD1.n198 VSUBS 0.036061f
C1683 VDD1.n199 VSUBS 0.036061f
C1684 VDD1.n200 VSUBS 0.016154f
C1685 VDD1.n201 VSUBS 0.015257f
C1686 VDD1.n202 VSUBS 0.028392f
C1687 VDD1.n203 VSUBS 0.028392f
C1688 VDD1.n204 VSUBS 0.015257f
C1689 VDD1.n205 VSUBS 0.016154f
C1690 VDD1.n206 VSUBS 0.036061f
C1691 VDD1.n207 VSUBS 0.087913f
C1692 VDD1.n208 VSUBS 0.016154f
C1693 VDD1.n209 VSUBS 0.029961f
C1694 VDD1.n210 VSUBS 0.069118f
C1695 VDD1.n211 VSUBS 0.104181f
C1696 VDD1.t0 VSUBS 0.43549f
C1697 VDD1.t1 VSUBS 0.43549f
C1698 VDD1.n212 VSUBS 3.66761f
C1699 VDD1.n213 VSUBS 1.19323f
C1700 VDD1.t4 VSUBS 0.43549f
C1701 VDD1.t6 VSUBS 0.43549f
C1702 VDD1.n214 VSUBS 3.69873f
C1703 VDD1.n215 VSUBS 4.60201f
C1704 VDD1.t5 VSUBS 0.43549f
C1705 VDD1.t9 VSUBS 0.43549f
C1706 VDD1.n216 VSUBS 3.66761f
C1707 VDD1.n217 VSUBS 4.79209f
C1708 VTAIL.t17 VSUBS 0.419506f
C1709 VTAIL.t19 VSUBS 0.419506f
C1710 VTAIL.n0 VSUBS 3.36811f
C1711 VTAIL.n1 VSUBS 1.02919f
C1712 VTAIL.n2 VSUBS 0.028586f
C1713 VTAIL.n3 VSUBS 0.02735f
C1714 VTAIL.n4 VSUBS 0.014697f
C1715 VTAIL.n5 VSUBS 0.034738f
C1716 VTAIL.n6 VSUBS 0.015561f
C1717 VTAIL.n7 VSUBS 0.02735f
C1718 VTAIL.n8 VSUBS 0.014697f
C1719 VTAIL.n9 VSUBS 0.034738f
C1720 VTAIL.n10 VSUBS 0.015561f
C1721 VTAIL.n11 VSUBS 0.02735f
C1722 VTAIL.n12 VSUBS 0.014697f
C1723 VTAIL.n13 VSUBS 0.034738f
C1724 VTAIL.n14 VSUBS 0.015561f
C1725 VTAIL.n15 VSUBS 0.02735f
C1726 VTAIL.n16 VSUBS 0.014697f
C1727 VTAIL.n17 VSUBS 0.034738f
C1728 VTAIL.n18 VSUBS 0.015561f
C1729 VTAIL.n19 VSUBS 0.02735f
C1730 VTAIL.n20 VSUBS 0.014697f
C1731 VTAIL.n21 VSUBS 0.034738f
C1732 VTAIL.n22 VSUBS 0.015561f
C1733 VTAIL.n23 VSUBS 0.02735f
C1734 VTAIL.n24 VSUBS 0.014697f
C1735 VTAIL.n25 VSUBS 0.034738f
C1736 VTAIL.n26 VSUBS 0.015561f
C1737 VTAIL.n27 VSUBS 0.02735f
C1738 VTAIL.n28 VSUBS 0.014697f
C1739 VTAIL.n29 VSUBS 0.034738f
C1740 VTAIL.n30 VSUBS 0.015561f
C1741 VTAIL.n31 VSUBS 0.02735f
C1742 VTAIL.n32 VSUBS 0.014697f
C1743 VTAIL.n33 VSUBS 0.034738f
C1744 VTAIL.n34 VSUBS 0.015561f
C1745 VTAIL.n35 VSUBS 0.307034f
C1746 VTAIL.t7 VSUBS 0.075541f
C1747 VTAIL.n36 VSUBS 0.026053f
C1748 VTAIL.n37 VSUBS 0.026132f
C1749 VTAIL.n38 VSUBS 0.014697f
C1750 VTAIL.n39 VSUBS 2.2318f
C1751 VTAIL.n40 VSUBS 0.02735f
C1752 VTAIL.n41 VSUBS 0.014697f
C1753 VTAIL.n42 VSUBS 0.015561f
C1754 VTAIL.n43 VSUBS 0.034738f
C1755 VTAIL.n44 VSUBS 0.034738f
C1756 VTAIL.n45 VSUBS 0.015561f
C1757 VTAIL.n46 VSUBS 0.014697f
C1758 VTAIL.n47 VSUBS 0.02735f
C1759 VTAIL.n48 VSUBS 0.02735f
C1760 VTAIL.n49 VSUBS 0.014697f
C1761 VTAIL.n50 VSUBS 0.015561f
C1762 VTAIL.n51 VSUBS 0.034738f
C1763 VTAIL.n52 VSUBS 0.034738f
C1764 VTAIL.n53 VSUBS 0.034738f
C1765 VTAIL.n54 VSUBS 0.015561f
C1766 VTAIL.n55 VSUBS 0.014697f
C1767 VTAIL.n56 VSUBS 0.02735f
C1768 VTAIL.n57 VSUBS 0.02735f
C1769 VTAIL.n58 VSUBS 0.014697f
C1770 VTAIL.n59 VSUBS 0.015129f
C1771 VTAIL.n60 VSUBS 0.015129f
C1772 VTAIL.n61 VSUBS 0.034738f
C1773 VTAIL.n62 VSUBS 0.034738f
C1774 VTAIL.n63 VSUBS 0.015561f
C1775 VTAIL.n64 VSUBS 0.014697f
C1776 VTAIL.n65 VSUBS 0.02735f
C1777 VTAIL.n66 VSUBS 0.02735f
C1778 VTAIL.n67 VSUBS 0.014697f
C1779 VTAIL.n68 VSUBS 0.015561f
C1780 VTAIL.n69 VSUBS 0.034738f
C1781 VTAIL.n70 VSUBS 0.034738f
C1782 VTAIL.n71 VSUBS 0.015561f
C1783 VTAIL.n72 VSUBS 0.014697f
C1784 VTAIL.n73 VSUBS 0.02735f
C1785 VTAIL.n74 VSUBS 0.02735f
C1786 VTAIL.n75 VSUBS 0.014697f
C1787 VTAIL.n76 VSUBS 0.015561f
C1788 VTAIL.n77 VSUBS 0.034738f
C1789 VTAIL.n78 VSUBS 0.034738f
C1790 VTAIL.n79 VSUBS 0.015561f
C1791 VTAIL.n80 VSUBS 0.014697f
C1792 VTAIL.n81 VSUBS 0.02735f
C1793 VTAIL.n82 VSUBS 0.02735f
C1794 VTAIL.n83 VSUBS 0.014697f
C1795 VTAIL.n84 VSUBS 0.015561f
C1796 VTAIL.n85 VSUBS 0.034738f
C1797 VTAIL.n86 VSUBS 0.034738f
C1798 VTAIL.n87 VSUBS 0.015561f
C1799 VTAIL.n88 VSUBS 0.014697f
C1800 VTAIL.n89 VSUBS 0.02735f
C1801 VTAIL.n90 VSUBS 0.02735f
C1802 VTAIL.n91 VSUBS 0.014697f
C1803 VTAIL.n92 VSUBS 0.015561f
C1804 VTAIL.n93 VSUBS 0.034738f
C1805 VTAIL.n94 VSUBS 0.034738f
C1806 VTAIL.n95 VSUBS 0.015561f
C1807 VTAIL.n96 VSUBS 0.014697f
C1808 VTAIL.n97 VSUBS 0.02735f
C1809 VTAIL.n98 VSUBS 0.02735f
C1810 VTAIL.n99 VSUBS 0.014697f
C1811 VTAIL.n100 VSUBS 0.015561f
C1812 VTAIL.n101 VSUBS 0.034738f
C1813 VTAIL.n102 VSUBS 0.084686f
C1814 VTAIL.n103 VSUBS 0.015561f
C1815 VTAIL.n104 VSUBS 0.028861f
C1816 VTAIL.n105 VSUBS 0.066581f
C1817 VTAIL.n106 VSUBS 0.064009f
C1818 VTAIL.n107 VSUBS 0.458683f
C1819 VTAIL.t11 VSUBS 0.419506f
C1820 VTAIL.t5 VSUBS 0.419506f
C1821 VTAIL.n108 VSUBS 3.36811f
C1822 VTAIL.n109 VSUBS 1.17866f
C1823 VTAIL.t12 VSUBS 0.419506f
C1824 VTAIL.t9 VSUBS 0.419506f
C1825 VTAIL.n110 VSUBS 3.36811f
C1826 VTAIL.n111 VSUBS 3.28615f
C1827 VTAIL.t16 VSUBS 0.419506f
C1828 VTAIL.t2 VSUBS 0.419506f
C1829 VTAIL.n112 VSUBS 3.36813f
C1830 VTAIL.n113 VSUBS 3.28613f
C1831 VTAIL.t14 VSUBS 0.419506f
C1832 VTAIL.t3 VSUBS 0.419506f
C1833 VTAIL.n114 VSUBS 3.36813f
C1834 VTAIL.n115 VSUBS 1.17864f
C1835 VTAIL.n116 VSUBS 0.028586f
C1836 VTAIL.n117 VSUBS 0.02735f
C1837 VTAIL.n118 VSUBS 0.014697f
C1838 VTAIL.n119 VSUBS 0.034738f
C1839 VTAIL.n120 VSUBS 0.015561f
C1840 VTAIL.n121 VSUBS 0.02735f
C1841 VTAIL.n122 VSUBS 0.014697f
C1842 VTAIL.n123 VSUBS 0.034738f
C1843 VTAIL.n124 VSUBS 0.015561f
C1844 VTAIL.n125 VSUBS 0.02735f
C1845 VTAIL.n126 VSUBS 0.014697f
C1846 VTAIL.n127 VSUBS 0.034738f
C1847 VTAIL.n128 VSUBS 0.015561f
C1848 VTAIL.n129 VSUBS 0.02735f
C1849 VTAIL.n130 VSUBS 0.014697f
C1850 VTAIL.n131 VSUBS 0.034738f
C1851 VTAIL.n132 VSUBS 0.015561f
C1852 VTAIL.n133 VSUBS 0.02735f
C1853 VTAIL.n134 VSUBS 0.014697f
C1854 VTAIL.n135 VSUBS 0.034738f
C1855 VTAIL.n136 VSUBS 0.015561f
C1856 VTAIL.n137 VSUBS 0.02735f
C1857 VTAIL.n138 VSUBS 0.014697f
C1858 VTAIL.n139 VSUBS 0.034738f
C1859 VTAIL.n140 VSUBS 0.015561f
C1860 VTAIL.n141 VSUBS 0.02735f
C1861 VTAIL.n142 VSUBS 0.014697f
C1862 VTAIL.n143 VSUBS 0.034738f
C1863 VTAIL.n144 VSUBS 0.034738f
C1864 VTAIL.n145 VSUBS 0.015561f
C1865 VTAIL.n146 VSUBS 0.02735f
C1866 VTAIL.n147 VSUBS 0.014697f
C1867 VTAIL.n148 VSUBS 0.034738f
C1868 VTAIL.n149 VSUBS 0.015561f
C1869 VTAIL.n150 VSUBS 0.307034f
C1870 VTAIL.t18 VSUBS 0.075541f
C1871 VTAIL.n151 VSUBS 0.026053f
C1872 VTAIL.n152 VSUBS 0.026132f
C1873 VTAIL.n153 VSUBS 0.014697f
C1874 VTAIL.n154 VSUBS 2.2318f
C1875 VTAIL.n155 VSUBS 0.02735f
C1876 VTAIL.n156 VSUBS 0.014697f
C1877 VTAIL.n157 VSUBS 0.015561f
C1878 VTAIL.n158 VSUBS 0.034738f
C1879 VTAIL.n159 VSUBS 0.034738f
C1880 VTAIL.n160 VSUBS 0.015561f
C1881 VTAIL.n161 VSUBS 0.014697f
C1882 VTAIL.n162 VSUBS 0.02735f
C1883 VTAIL.n163 VSUBS 0.02735f
C1884 VTAIL.n164 VSUBS 0.014697f
C1885 VTAIL.n165 VSUBS 0.015561f
C1886 VTAIL.n166 VSUBS 0.034738f
C1887 VTAIL.n167 VSUBS 0.034738f
C1888 VTAIL.n168 VSUBS 0.015561f
C1889 VTAIL.n169 VSUBS 0.014697f
C1890 VTAIL.n170 VSUBS 0.02735f
C1891 VTAIL.n171 VSUBS 0.02735f
C1892 VTAIL.n172 VSUBS 0.014697f
C1893 VTAIL.n173 VSUBS 0.015129f
C1894 VTAIL.n174 VSUBS 0.015129f
C1895 VTAIL.n175 VSUBS 0.034738f
C1896 VTAIL.n176 VSUBS 0.034738f
C1897 VTAIL.n177 VSUBS 0.015561f
C1898 VTAIL.n178 VSUBS 0.014697f
C1899 VTAIL.n179 VSUBS 0.02735f
C1900 VTAIL.n180 VSUBS 0.02735f
C1901 VTAIL.n181 VSUBS 0.014697f
C1902 VTAIL.n182 VSUBS 0.015561f
C1903 VTAIL.n183 VSUBS 0.034738f
C1904 VTAIL.n184 VSUBS 0.034738f
C1905 VTAIL.n185 VSUBS 0.015561f
C1906 VTAIL.n186 VSUBS 0.014697f
C1907 VTAIL.n187 VSUBS 0.02735f
C1908 VTAIL.n188 VSUBS 0.02735f
C1909 VTAIL.n189 VSUBS 0.014697f
C1910 VTAIL.n190 VSUBS 0.015561f
C1911 VTAIL.n191 VSUBS 0.034738f
C1912 VTAIL.n192 VSUBS 0.034738f
C1913 VTAIL.n193 VSUBS 0.015561f
C1914 VTAIL.n194 VSUBS 0.014697f
C1915 VTAIL.n195 VSUBS 0.02735f
C1916 VTAIL.n196 VSUBS 0.02735f
C1917 VTAIL.n197 VSUBS 0.014697f
C1918 VTAIL.n198 VSUBS 0.015561f
C1919 VTAIL.n199 VSUBS 0.034738f
C1920 VTAIL.n200 VSUBS 0.034738f
C1921 VTAIL.n201 VSUBS 0.015561f
C1922 VTAIL.n202 VSUBS 0.014697f
C1923 VTAIL.n203 VSUBS 0.02735f
C1924 VTAIL.n204 VSUBS 0.02735f
C1925 VTAIL.n205 VSUBS 0.014697f
C1926 VTAIL.n206 VSUBS 0.015561f
C1927 VTAIL.n207 VSUBS 0.034738f
C1928 VTAIL.n208 VSUBS 0.034738f
C1929 VTAIL.n209 VSUBS 0.015561f
C1930 VTAIL.n210 VSUBS 0.014697f
C1931 VTAIL.n211 VSUBS 0.02735f
C1932 VTAIL.n212 VSUBS 0.02735f
C1933 VTAIL.n213 VSUBS 0.014697f
C1934 VTAIL.n214 VSUBS 0.015561f
C1935 VTAIL.n215 VSUBS 0.034738f
C1936 VTAIL.n216 VSUBS 0.084686f
C1937 VTAIL.n217 VSUBS 0.015561f
C1938 VTAIL.n218 VSUBS 0.028861f
C1939 VTAIL.n219 VSUBS 0.066581f
C1940 VTAIL.n220 VSUBS 0.064009f
C1941 VTAIL.n221 VSUBS 0.458683f
C1942 VTAIL.t8 VSUBS 0.419506f
C1943 VTAIL.t13 VSUBS 0.419506f
C1944 VTAIL.n222 VSUBS 3.36813f
C1945 VTAIL.n223 VSUBS 1.08938f
C1946 VTAIL.t6 VSUBS 0.419506f
C1947 VTAIL.t4 VSUBS 0.419506f
C1948 VTAIL.n224 VSUBS 3.36813f
C1949 VTAIL.n225 VSUBS 1.17864f
C1950 VTAIL.n226 VSUBS 0.028586f
C1951 VTAIL.n227 VSUBS 0.02735f
C1952 VTAIL.n228 VSUBS 0.014697f
C1953 VTAIL.n229 VSUBS 0.034738f
C1954 VTAIL.n230 VSUBS 0.015561f
C1955 VTAIL.n231 VSUBS 0.02735f
C1956 VTAIL.n232 VSUBS 0.014697f
C1957 VTAIL.n233 VSUBS 0.034738f
C1958 VTAIL.n234 VSUBS 0.015561f
C1959 VTAIL.n235 VSUBS 0.02735f
C1960 VTAIL.n236 VSUBS 0.014697f
C1961 VTAIL.n237 VSUBS 0.034738f
C1962 VTAIL.n238 VSUBS 0.015561f
C1963 VTAIL.n239 VSUBS 0.02735f
C1964 VTAIL.n240 VSUBS 0.014697f
C1965 VTAIL.n241 VSUBS 0.034738f
C1966 VTAIL.n242 VSUBS 0.015561f
C1967 VTAIL.n243 VSUBS 0.02735f
C1968 VTAIL.n244 VSUBS 0.014697f
C1969 VTAIL.n245 VSUBS 0.034738f
C1970 VTAIL.n246 VSUBS 0.015561f
C1971 VTAIL.n247 VSUBS 0.02735f
C1972 VTAIL.n248 VSUBS 0.014697f
C1973 VTAIL.n249 VSUBS 0.034738f
C1974 VTAIL.n250 VSUBS 0.015561f
C1975 VTAIL.n251 VSUBS 0.02735f
C1976 VTAIL.n252 VSUBS 0.014697f
C1977 VTAIL.n253 VSUBS 0.034738f
C1978 VTAIL.n254 VSUBS 0.034738f
C1979 VTAIL.n255 VSUBS 0.015561f
C1980 VTAIL.n256 VSUBS 0.02735f
C1981 VTAIL.n257 VSUBS 0.014697f
C1982 VTAIL.n258 VSUBS 0.034738f
C1983 VTAIL.n259 VSUBS 0.015561f
C1984 VTAIL.n260 VSUBS 0.307034f
C1985 VTAIL.t10 VSUBS 0.075541f
C1986 VTAIL.n261 VSUBS 0.026053f
C1987 VTAIL.n262 VSUBS 0.026132f
C1988 VTAIL.n263 VSUBS 0.014697f
C1989 VTAIL.n264 VSUBS 2.2318f
C1990 VTAIL.n265 VSUBS 0.02735f
C1991 VTAIL.n266 VSUBS 0.014697f
C1992 VTAIL.n267 VSUBS 0.015561f
C1993 VTAIL.n268 VSUBS 0.034738f
C1994 VTAIL.n269 VSUBS 0.034738f
C1995 VTAIL.n270 VSUBS 0.015561f
C1996 VTAIL.n271 VSUBS 0.014697f
C1997 VTAIL.n272 VSUBS 0.02735f
C1998 VTAIL.n273 VSUBS 0.02735f
C1999 VTAIL.n274 VSUBS 0.014697f
C2000 VTAIL.n275 VSUBS 0.015561f
C2001 VTAIL.n276 VSUBS 0.034738f
C2002 VTAIL.n277 VSUBS 0.034738f
C2003 VTAIL.n278 VSUBS 0.015561f
C2004 VTAIL.n279 VSUBS 0.014697f
C2005 VTAIL.n280 VSUBS 0.02735f
C2006 VTAIL.n281 VSUBS 0.02735f
C2007 VTAIL.n282 VSUBS 0.014697f
C2008 VTAIL.n283 VSUBS 0.015129f
C2009 VTAIL.n284 VSUBS 0.015129f
C2010 VTAIL.n285 VSUBS 0.034738f
C2011 VTAIL.n286 VSUBS 0.034738f
C2012 VTAIL.n287 VSUBS 0.015561f
C2013 VTAIL.n288 VSUBS 0.014697f
C2014 VTAIL.n289 VSUBS 0.02735f
C2015 VTAIL.n290 VSUBS 0.02735f
C2016 VTAIL.n291 VSUBS 0.014697f
C2017 VTAIL.n292 VSUBS 0.015561f
C2018 VTAIL.n293 VSUBS 0.034738f
C2019 VTAIL.n294 VSUBS 0.034738f
C2020 VTAIL.n295 VSUBS 0.015561f
C2021 VTAIL.n296 VSUBS 0.014697f
C2022 VTAIL.n297 VSUBS 0.02735f
C2023 VTAIL.n298 VSUBS 0.02735f
C2024 VTAIL.n299 VSUBS 0.014697f
C2025 VTAIL.n300 VSUBS 0.015561f
C2026 VTAIL.n301 VSUBS 0.034738f
C2027 VTAIL.n302 VSUBS 0.034738f
C2028 VTAIL.n303 VSUBS 0.015561f
C2029 VTAIL.n304 VSUBS 0.014697f
C2030 VTAIL.n305 VSUBS 0.02735f
C2031 VTAIL.n306 VSUBS 0.02735f
C2032 VTAIL.n307 VSUBS 0.014697f
C2033 VTAIL.n308 VSUBS 0.015561f
C2034 VTAIL.n309 VSUBS 0.034738f
C2035 VTAIL.n310 VSUBS 0.034738f
C2036 VTAIL.n311 VSUBS 0.015561f
C2037 VTAIL.n312 VSUBS 0.014697f
C2038 VTAIL.n313 VSUBS 0.02735f
C2039 VTAIL.n314 VSUBS 0.02735f
C2040 VTAIL.n315 VSUBS 0.014697f
C2041 VTAIL.n316 VSUBS 0.015561f
C2042 VTAIL.n317 VSUBS 0.034738f
C2043 VTAIL.n318 VSUBS 0.034738f
C2044 VTAIL.n319 VSUBS 0.015561f
C2045 VTAIL.n320 VSUBS 0.014697f
C2046 VTAIL.n321 VSUBS 0.02735f
C2047 VTAIL.n322 VSUBS 0.02735f
C2048 VTAIL.n323 VSUBS 0.014697f
C2049 VTAIL.n324 VSUBS 0.015561f
C2050 VTAIL.n325 VSUBS 0.034738f
C2051 VTAIL.n326 VSUBS 0.084686f
C2052 VTAIL.n327 VSUBS 0.015561f
C2053 VTAIL.n328 VSUBS 0.028861f
C2054 VTAIL.n329 VSUBS 0.066581f
C2055 VTAIL.n330 VSUBS 0.064009f
C2056 VTAIL.n331 VSUBS 2.3941f
C2057 VTAIL.n332 VSUBS 0.028586f
C2058 VTAIL.n333 VSUBS 0.02735f
C2059 VTAIL.n334 VSUBS 0.014697f
C2060 VTAIL.n335 VSUBS 0.034738f
C2061 VTAIL.n336 VSUBS 0.015561f
C2062 VTAIL.n337 VSUBS 0.02735f
C2063 VTAIL.n338 VSUBS 0.014697f
C2064 VTAIL.n339 VSUBS 0.034738f
C2065 VTAIL.n340 VSUBS 0.015561f
C2066 VTAIL.n341 VSUBS 0.02735f
C2067 VTAIL.n342 VSUBS 0.014697f
C2068 VTAIL.n343 VSUBS 0.034738f
C2069 VTAIL.n344 VSUBS 0.015561f
C2070 VTAIL.n345 VSUBS 0.02735f
C2071 VTAIL.n346 VSUBS 0.014697f
C2072 VTAIL.n347 VSUBS 0.034738f
C2073 VTAIL.n348 VSUBS 0.015561f
C2074 VTAIL.n349 VSUBS 0.02735f
C2075 VTAIL.n350 VSUBS 0.014697f
C2076 VTAIL.n351 VSUBS 0.034738f
C2077 VTAIL.n352 VSUBS 0.015561f
C2078 VTAIL.n353 VSUBS 0.02735f
C2079 VTAIL.n354 VSUBS 0.014697f
C2080 VTAIL.n355 VSUBS 0.034738f
C2081 VTAIL.n356 VSUBS 0.015561f
C2082 VTAIL.n357 VSUBS 0.02735f
C2083 VTAIL.n358 VSUBS 0.014697f
C2084 VTAIL.n359 VSUBS 0.034738f
C2085 VTAIL.n360 VSUBS 0.015561f
C2086 VTAIL.n361 VSUBS 0.02735f
C2087 VTAIL.n362 VSUBS 0.014697f
C2088 VTAIL.n363 VSUBS 0.034738f
C2089 VTAIL.n364 VSUBS 0.015561f
C2090 VTAIL.n365 VSUBS 0.307034f
C2091 VTAIL.t1 VSUBS 0.075541f
C2092 VTAIL.n366 VSUBS 0.026053f
C2093 VTAIL.n367 VSUBS 0.026132f
C2094 VTAIL.n368 VSUBS 0.014697f
C2095 VTAIL.n369 VSUBS 2.2318f
C2096 VTAIL.n370 VSUBS 0.02735f
C2097 VTAIL.n371 VSUBS 0.014697f
C2098 VTAIL.n372 VSUBS 0.015561f
C2099 VTAIL.n373 VSUBS 0.034738f
C2100 VTAIL.n374 VSUBS 0.034738f
C2101 VTAIL.n375 VSUBS 0.015561f
C2102 VTAIL.n376 VSUBS 0.014697f
C2103 VTAIL.n377 VSUBS 0.02735f
C2104 VTAIL.n378 VSUBS 0.02735f
C2105 VTAIL.n379 VSUBS 0.014697f
C2106 VTAIL.n380 VSUBS 0.015561f
C2107 VTAIL.n381 VSUBS 0.034738f
C2108 VTAIL.n382 VSUBS 0.034738f
C2109 VTAIL.n383 VSUBS 0.034738f
C2110 VTAIL.n384 VSUBS 0.015561f
C2111 VTAIL.n385 VSUBS 0.014697f
C2112 VTAIL.n386 VSUBS 0.02735f
C2113 VTAIL.n387 VSUBS 0.02735f
C2114 VTAIL.n388 VSUBS 0.014697f
C2115 VTAIL.n389 VSUBS 0.015129f
C2116 VTAIL.n390 VSUBS 0.015129f
C2117 VTAIL.n391 VSUBS 0.034738f
C2118 VTAIL.n392 VSUBS 0.034738f
C2119 VTAIL.n393 VSUBS 0.015561f
C2120 VTAIL.n394 VSUBS 0.014697f
C2121 VTAIL.n395 VSUBS 0.02735f
C2122 VTAIL.n396 VSUBS 0.02735f
C2123 VTAIL.n397 VSUBS 0.014697f
C2124 VTAIL.n398 VSUBS 0.015561f
C2125 VTAIL.n399 VSUBS 0.034738f
C2126 VTAIL.n400 VSUBS 0.034738f
C2127 VTAIL.n401 VSUBS 0.015561f
C2128 VTAIL.n402 VSUBS 0.014697f
C2129 VTAIL.n403 VSUBS 0.02735f
C2130 VTAIL.n404 VSUBS 0.02735f
C2131 VTAIL.n405 VSUBS 0.014697f
C2132 VTAIL.n406 VSUBS 0.015561f
C2133 VTAIL.n407 VSUBS 0.034738f
C2134 VTAIL.n408 VSUBS 0.034738f
C2135 VTAIL.n409 VSUBS 0.015561f
C2136 VTAIL.n410 VSUBS 0.014697f
C2137 VTAIL.n411 VSUBS 0.02735f
C2138 VTAIL.n412 VSUBS 0.02735f
C2139 VTAIL.n413 VSUBS 0.014697f
C2140 VTAIL.n414 VSUBS 0.015561f
C2141 VTAIL.n415 VSUBS 0.034738f
C2142 VTAIL.n416 VSUBS 0.034738f
C2143 VTAIL.n417 VSUBS 0.015561f
C2144 VTAIL.n418 VSUBS 0.014697f
C2145 VTAIL.n419 VSUBS 0.02735f
C2146 VTAIL.n420 VSUBS 0.02735f
C2147 VTAIL.n421 VSUBS 0.014697f
C2148 VTAIL.n422 VSUBS 0.015561f
C2149 VTAIL.n423 VSUBS 0.034738f
C2150 VTAIL.n424 VSUBS 0.034738f
C2151 VTAIL.n425 VSUBS 0.015561f
C2152 VTAIL.n426 VSUBS 0.014697f
C2153 VTAIL.n427 VSUBS 0.02735f
C2154 VTAIL.n428 VSUBS 0.02735f
C2155 VTAIL.n429 VSUBS 0.014697f
C2156 VTAIL.n430 VSUBS 0.015561f
C2157 VTAIL.n431 VSUBS 0.034738f
C2158 VTAIL.n432 VSUBS 0.084686f
C2159 VTAIL.n433 VSUBS 0.015561f
C2160 VTAIL.n434 VSUBS 0.028861f
C2161 VTAIL.n435 VSUBS 0.066581f
C2162 VTAIL.n436 VSUBS 0.064009f
C2163 VTAIL.n437 VSUBS 2.3941f
C2164 VTAIL.t15 VSUBS 0.419506f
C2165 VTAIL.t0 VSUBS 0.419506f
C2166 VTAIL.n438 VSUBS 3.36811f
C2167 VTAIL.n439 VSUBS 0.977526f
C2168 VP.t3 VSUBS 3.96771f
C2169 VP.n0 VSUBS 1.46265f
C2170 VP.n1 VSUBS 0.023864f
C2171 VP.n2 VSUBS 0.028493f
C2172 VP.n3 VSUBS 0.023864f
C2173 VP.t5 VSUBS 3.96771f
C2174 VP.n4 VSUBS 1.36764f
C2175 VP.n5 VSUBS 0.023864f
C2176 VP.n6 VSUBS 0.032842f
C2177 VP.n7 VSUBS 0.023864f
C2178 VP.t8 VSUBS 3.96771f
C2179 VP.n8 VSUBS 0.044476f
C2180 VP.n9 VSUBS 0.023864f
C2181 VP.n10 VSUBS 0.044476f
C2182 VP.n11 VSUBS 0.023864f
C2183 VP.t9 VSUBS 3.96771f
C2184 VP.n12 VSUBS 0.044893f
C2185 VP.n13 VSUBS 0.023864f
C2186 VP.n14 VSUBS 0.039206f
C2187 VP.t0 VSUBS 3.96771f
C2188 VP.n15 VSUBS 1.46265f
C2189 VP.n16 VSUBS 0.023864f
C2190 VP.n17 VSUBS 0.028493f
C2191 VP.n18 VSUBS 0.023864f
C2192 VP.t4 VSUBS 3.96771f
C2193 VP.n19 VSUBS 1.36764f
C2194 VP.n20 VSUBS 0.023864f
C2195 VP.n21 VSUBS 0.032842f
C2196 VP.n22 VSUBS 0.023864f
C2197 VP.t6 VSUBS 3.96771f
C2198 VP.n23 VSUBS 0.044476f
C2199 VP.n24 VSUBS 0.023864f
C2200 VP.n25 VSUBS 0.044476f
C2201 VP.t2 VSUBS 4.24654f
C2202 VP.n26 VSUBS 1.39783f
C2203 VP.t1 VSUBS 3.96771f
C2204 VP.n27 VSUBS 1.45385f
C2205 VP.n28 VSUBS 0.041841f
C2206 VP.n29 VSUBS 0.273159f
C2207 VP.n30 VSUBS 0.023864f
C2208 VP.n31 VSUBS 0.023864f
C2209 VP.n32 VSUBS 0.036832f
C2210 VP.n33 VSUBS 0.032842f
C2211 VP.n34 VSUBS 0.044476f
C2212 VP.n35 VSUBS 0.023864f
C2213 VP.n36 VSUBS 0.023864f
C2214 VP.n37 VSUBS 0.023864f
C2215 VP.n38 VSUBS 1.39015f
C2216 VP.n39 VSUBS 0.044476f
C2217 VP.n40 VSUBS 0.044476f
C2218 VP.n41 VSUBS 0.023864f
C2219 VP.n42 VSUBS 0.023864f
C2220 VP.n43 VSUBS 0.023864f
C2221 VP.n44 VSUBS 0.036832f
C2222 VP.n45 VSUBS 0.044476f
C2223 VP.n46 VSUBS 0.041841f
C2224 VP.n47 VSUBS 0.023864f
C2225 VP.n48 VSUBS 0.023864f
C2226 VP.n49 VSUBS 0.025153f
C2227 VP.n50 VSUBS 0.044476f
C2228 VP.n51 VSUBS 0.044893f
C2229 VP.n52 VSUBS 0.023864f
C2230 VP.n53 VSUBS 0.023864f
C2231 VP.n54 VSUBS 0.023864f
C2232 VP.n55 VSUBS 0.040763f
C2233 VP.n56 VSUBS 0.044476f
C2234 VP.n57 VSUBS 0.039206f
C2235 VP.n58 VSUBS 0.038515f
C2236 VP.n59 VSUBS 1.80499f
C2237 VP.t7 VSUBS 3.96771f
C2238 VP.n60 VSUBS 1.46265f
C2239 VP.n61 VSUBS 1.81891f
C2240 VP.n62 VSUBS 0.038515f
C2241 VP.n63 VSUBS 0.023864f
C2242 VP.n64 VSUBS 0.044476f
C2243 VP.n65 VSUBS 0.040763f
C2244 VP.n66 VSUBS 0.028493f
C2245 VP.n67 VSUBS 0.023864f
C2246 VP.n68 VSUBS 0.023864f
C2247 VP.n69 VSUBS 0.023864f
C2248 VP.n70 VSUBS 0.044476f
C2249 VP.n71 VSUBS 0.025153f
C2250 VP.n72 VSUBS 1.36764f
C2251 VP.n73 VSUBS 0.041841f
C2252 VP.n74 VSUBS 0.023864f
C2253 VP.n75 VSUBS 0.023864f
C2254 VP.n76 VSUBS 0.023864f
C2255 VP.n77 VSUBS 0.036832f
C2256 VP.n78 VSUBS 0.032842f
C2257 VP.n79 VSUBS 0.044476f
C2258 VP.n80 VSUBS 0.023864f
C2259 VP.n81 VSUBS 0.023864f
C2260 VP.n82 VSUBS 0.023864f
C2261 VP.n83 VSUBS 1.39015f
C2262 VP.n84 VSUBS 0.044476f
C2263 VP.n85 VSUBS 0.044476f
C2264 VP.n86 VSUBS 0.023864f
C2265 VP.n87 VSUBS 0.023864f
C2266 VP.n88 VSUBS 0.023864f
C2267 VP.n89 VSUBS 0.036832f
C2268 VP.n90 VSUBS 0.044476f
C2269 VP.n91 VSUBS 0.041841f
C2270 VP.n92 VSUBS 0.023864f
C2271 VP.n93 VSUBS 0.023864f
C2272 VP.n94 VSUBS 0.025153f
C2273 VP.n95 VSUBS 0.044476f
C2274 VP.n96 VSUBS 0.044893f
C2275 VP.n97 VSUBS 0.023864f
C2276 VP.n98 VSUBS 0.023864f
C2277 VP.n99 VSUBS 0.023864f
C2278 VP.n100 VSUBS 0.040763f
C2279 VP.n101 VSUBS 0.044476f
C2280 VP.n102 VSUBS 0.039206f
C2281 VP.n103 VSUBS 0.038515f
C2282 VP.n104 VSUBS 0.052062f
.ends

