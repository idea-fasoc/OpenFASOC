* NGSPICE file created from diff_pair_sample_0553.ext - technology: sky130A

.subckt diff_pair_sample_0553 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0.4455 ps=3.03 w=2.7 l=1.6
X1 VDD2.t2 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4455 pd=3.03 as=1.053 ps=6.18 w=2.7 l=1.6
X2 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0.4455 ps=3.03 w=2.7 l=1.6
X3 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4455 pd=3.03 as=1.053 ps=6.18 w=2.7 l=1.6
X4 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0.4455 ps=3.03 w=2.7 l=1.6
X5 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0 ps=0 w=2.7 l=1.6
X6 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4455 pd=3.03 as=1.053 ps=6.18 w=2.7 l=1.6
X7 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4455 pd=3.03 as=1.053 ps=6.18 w=2.7 l=1.6
X8 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0 ps=0 w=2.7 l=1.6
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0 ps=0 w=2.7 l=1.6
X10 VTAIL.t4 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0.4455 ps=3.03 w=2.7 l=1.6
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.053 pd=6.18 as=0 ps=0 w=2.7 l=1.6
R0 VN.n0 VN.t3 78.549
R1 VN.n1 VN.t2 78.549
R2 VN.n0 VN.t1 78.2235
R3 VN.n1 VN.t0 78.2235
R4 VN VN.n1 49.2243
R5 VN VN.n0 12.6902
R6 VDD2.n2 VDD2.n0 116.288
R7 VDD2.n2 VDD2.n1 85.2545
R8 VDD2.n1 VDD2.t1 7.33383
R9 VDD2.n1 VDD2.t3 7.33383
R10 VDD2.n0 VDD2.t0 7.33383
R11 VDD2.n0 VDD2.t2 7.33383
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n90 VTAIL.n84 289.615
R14 VTAIL.n6 VTAIL.n0 289.615
R15 VTAIL.n18 VTAIL.n12 289.615
R16 VTAIL.n30 VTAIL.n24 289.615
R17 VTAIL.n78 VTAIL.n72 289.615
R18 VTAIL.n66 VTAIL.n60 289.615
R19 VTAIL.n54 VTAIL.n48 289.615
R20 VTAIL.n42 VTAIL.n36 289.615
R21 VTAIL.n89 VTAIL.n88 185
R22 VTAIL.n91 VTAIL.n90 185
R23 VTAIL.n5 VTAIL.n4 185
R24 VTAIL.n7 VTAIL.n6 185
R25 VTAIL.n17 VTAIL.n16 185
R26 VTAIL.n19 VTAIL.n18 185
R27 VTAIL.n29 VTAIL.n28 185
R28 VTAIL.n31 VTAIL.n30 185
R29 VTAIL.n79 VTAIL.n78 185
R30 VTAIL.n77 VTAIL.n76 185
R31 VTAIL.n67 VTAIL.n66 185
R32 VTAIL.n65 VTAIL.n64 185
R33 VTAIL.n55 VTAIL.n54 185
R34 VTAIL.n53 VTAIL.n52 185
R35 VTAIL.n43 VTAIL.n42 185
R36 VTAIL.n41 VTAIL.n40 185
R37 VTAIL.n87 VTAIL.t6 153.582
R38 VTAIL.n3 VTAIL.t4 153.582
R39 VTAIL.n15 VTAIL.t3 153.582
R40 VTAIL.n27 VTAIL.t2 153.582
R41 VTAIL.n75 VTAIL.t0 153.582
R42 VTAIL.n63 VTAIL.t1 153.582
R43 VTAIL.n51 VTAIL.t5 153.582
R44 VTAIL.n39 VTAIL.t7 153.582
R45 VTAIL.n90 VTAIL.n89 104.615
R46 VTAIL.n6 VTAIL.n5 104.615
R47 VTAIL.n18 VTAIL.n17 104.615
R48 VTAIL.n30 VTAIL.n29 104.615
R49 VTAIL.n78 VTAIL.n77 104.615
R50 VTAIL.n66 VTAIL.n65 104.615
R51 VTAIL.n54 VTAIL.n53 104.615
R52 VTAIL.n42 VTAIL.n41 104.615
R53 VTAIL.n89 VTAIL.t6 52.3082
R54 VTAIL.n5 VTAIL.t4 52.3082
R55 VTAIL.n17 VTAIL.t3 52.3082
R56 VTAIL.n29 VTAIL.t2 52.3082
R57 VTAIL.n77 VTAIL.t0 52.3082
R58 VTAIL.n65 VTAIL.t1 52.3082
R59 VTAIL.n53 VTAIL.t5 52.3082
R60 VTAIL.n41 VTAIL.t7 52.3082
R61 VTAIL.n95 VTAIL.n94 31.0217
R62 VTAIL.n11 VTAIL.n10 31.0217
R63 VTAIL.n23 VTAIL.n22 31.0217
R64 VTAIL.n35 VTAIL.n34 31.0217
R65 VTAIL.n83 VTAIL.n82 31.0217
R66 VTAIL.n71 VTAIL.n70 31.0217
R67 VTAIL.n59 VTAIL.n58 31.0217
R68 VTAIL.n47 VTAIL.n46 31.0217
R69 VTAIL.n95 VTAIL.n83 16.3583
R70 VTAIL.n47 VTAIL.n35 16.3583
R71 VTAIL.n88 VTAIL.n87 10.1164
R72 VTAIL.n4 VTAIL.n3 10.1164
R73 VTAIL.n16 VTAIL.n15 10.1164
R74 VTAIL.n28 VTAIL.n27 10.1164
R75 VTAIL.n76 VTAIL.n75 10.1164
R76 VTAIL.n64 VTAIL.n63 10.1164
R77 VTAIL.n52 VTAIL.n51 10.1164
R78 VTAIL.n40 VTAIL.n39 10.1164
R79 VTAIL.n94 VTAIL.n93 9.45567
R80 VTAIL.n10 VTAIL.n9 9.45567
R81 VTAIL.n22 VTAIL.n21 9.45567
R82 VTAIL.n34 VTAIL.n33 9.45567
R83 VTAIL.n82 VTAIL.n81 9.45567
R84 VTAIL.n70 VTAIL.n69 9.45567
R85 VTAIL.n58 VTAIL.n57 9.45567
R86 VTAIL.n46 VTAIL.n45 9.45567
R87 VTAIL.n86 VTAIL.n85 9.3005
R88 VTAIL.n93 VTAIL.n92 9.3005
R89 VTAIL.n2 VTAIL.n1 9.3005
R90 VTAIL.n9 VTAIL.n8 9.3005
R91 VTAIL.n14 VTAIL.n13 9.3005
R92 VTAIL.n21 VTAIL.n20 9.3005
R93 VTAIL.n26 VTAIL.n25 9.3005
R94 VTAIL.n33 VTAIL.n32 9.3005
R95 VTAIL.n74 VTAIL.n73 9.3005
R96 VTAIL.n81 VTAIL.n80 9.3005
R97 VTAIL.n69 VTAIL.n68 9.3005
R98 VTAIL.n62 VTAIL.n61 9.3005
R99 VTAIL.n57 VTAIL.n56 9.3005
R100 VTAIL.n50 VTAIL.n49 9.3005
R101 VTAIL.n45 VTAIL.n44 9.3005
R102 VTAIL.n38 VTAIL.n37 9.3005
R103 VTAIL.n94 VTAIL.n84 8.92171
R104 VTAIL.n10 VTAIL.n0 8.92171
R105 VTAIL.n22 VTAIL.n12 8.92171
R106 VTAIL.n34 VTAIL.n24 8.92171
R107 VTAIL.n82 VTAIL.n72 8.92171
R108 VTAIL.n70 VTAIL.n60 8.92171
R109 VTAIL.n58 VTAIL.n48 8.92171
R110 VTAIL.n46 VTAIL.n36 8.92171
R111 VTAIL.n92 VTAIL.n91 8.14595
R112 VTAIL.n8 VTAIL.n7 8.14595
R113 VTAIL.n20 VTAIL.n19 8.14595
R114 VTAIL.n32 VTAIL.n31 8.14595
R115 VTAIL.n80 VTAIL.n79 8.14595
R116 VTAIL.n68 VTAIL.n67 8.14595
R117 VTAIL.n56 VTAIL.n55 8.14595
R118 VTAIL.n44 VTAIL.n43 8.14595
R119 VTAIL.n88 VTAIL.n86 7.3702
R120 VTAIL.n4 VTAIL.n2 7.3702
R121 VTAIL.n16 VTAIL.n14 7.3702
R122 VTAIL.n28 VTAIL.n26 7.3702
R123 VTAIL.n76 VTAIL.n74 7.3702
R124 VTAIL.n64 VTAIL.n62 7.3702
R125 VTAIL.n52 VTAIL.n50 7.3702
R126 VTAIL.n40 VTAIL.n38 7.3702
R127 VTAIL.n91 VTAIL.n86 5.81868
R128 VTAIL.n7 VTAIL.n2 5.81868
R129 VTAIL.n19 VTAIL.n14 5.81868
R130 VTAIL.n31 VTAIL.n26 5.81868
R131 VTAIL.n79 VTAIL.n74 5.81868
R132 VTAIL.n67 VTAIL.n62 5.81868
R133 VTAIL.n55 VTAIL.n50 5.81868
R134 VTAIL.n43 VTAIL.n38 5.81868
R135 VTAIL.n92 VTAIL.n84 5.04292
R136 VTAIL.n8 VTAIL.n0 5.04292
R137 VTAIL.n20 VTAIL.n12 5.04292
R138 VTAIL.n32 VTAIL.n24 5.04292
R139 VTAIL.n80 VTAIL.n72 5.04292
R140 VTAIL.n68 VTAIL.n60 5.04292
R141 VTAIL.n56 VTAIL.n48 5.04292
R142 VTAIL.n44 VTAIL.n36 5.04292
R143 VTAIL.n63 VTAIL.n61 3.00987
R144 VTAIL.n51 VTAIL.n49 3.00987
R145 VTAIL.n39 VTAIL.n37 3.00987
R146 VTAIL.n87 VTAIL.n85 3.00987
R147 VTAIL.n3 VTAIL.n1 3.00987
R148 VTAIL.n15 VTAIL.n13 3.00987
R149 VTAIL.n27 VTAIL.n25 3.00987
R150 VTAIL.n75 VTAIL.n73 3.00987
R151 VTAIL.n59 VTAIL.n47 1.66429
R152 VTAIL.n83 VTAIL.n71 1.66429
R153 VTAIL.n35 VTAIL.n23 1.66429
R154 VTAIL VTAIL.n11 0.890586
R155 VTAIL VTAIL.n95 0.774207
R156 VTAIL.n71 VTAIL.n59 0.470328
R157 VTAIL.n23 VTAIL.n11 0.470328
R158 VTAIL.n93 VTAIL.n85 0.155672
R159 VTAIL.n9 VTAIL.n1 0.155672
R160 VTAIL.n21 VTAIL.n13 0.155672
R161 VTAIL.n33 VTAIL.n25 0.155672
R162 VTAIL.n81 VTAIL.n73 0.155672
R163 VTAIL.n69 VTAIL.n61 0.155672
R164 VTAIL.n57 VTAIL.n49 0.155672
R165 VTAIL.n45 VTAIL.n37 0.155672
R166 B.n401 B.n400 585
R167 B.n145 B.n66 585
R168 B.n144 B.n143 585
R169 B.n142 B.n141 585
R170 B.n140 B.n139 585
R171 B.n138 B.n137 585
R172 B.n136 B.n135 585
R173 B.n134 B.n133 585
R174 B.n132 B.n131 585
R175 B.n130 B.n129 585
R176 B.n128 B.n127 585
R177 B.n126 B.n125 585
R178 B.n124 B.n123 585
R179 B.n122 B.n121 585
R180 B.n120 B.n119 585
R181 B.n118 B.n117 585
R182 B.n116 B.n115 585
R183 B.n114 B.n113 585
R184 B.n112 B.n111 585
R185 B.n110 B.n109 585
R186 B.n108 B.n107 585
R187 B.n106 B.n105 585
R188 B.n104 B.n103 585
R189 B.n102 B.n101 585
R190 B.n100 B.n99 585
R191 B.n98 B.n97 585
R192 B.n96 B.n95 585
R193 B.n94 B.n93 585
R194 B.n92 B.n91 585
R195 B.n90 B.n89 585
R196 B.n88 B.n87 585
R197 B.n86 B.n85 585
R198 B.n84 B.n83 585
R199 B.n82 B.n81 585
R200 B.n80 B.n79 585
R201 B.n78 B.n77 585
R202 B.n76 B.n75 585
R203 B.n74 B.n73 585
R204 B.n399 B.n47 585
R205 B.n404 B.n47 585
R206 B.n398 B.n46 585
R207 B.n405 B.n46 585
R208 B.n397 B.n396 585
R209 B.n396 B.n42 585
R210 B.n395 B.n41 585
R211 B.n411 B.n41 585
R212 B.n394 B.n40 585
R213 B.n412 B.n40 585
R214 B.n393 B.n39 585
R215 B.n413 B.n39 585
R216 B.n392 B.n391 585
R217 B.n391 B.t12 585
R218 B.n390 B.n35 585
R219 B.n419 B.n35 585
R220 B.n389 B.n34 585
R221 B.n420 B.n34 585
R222 B.n388 B.n33 585
R223 B.n421 B.n33 585
R224 B.n387 B.n386 585
R225 B.n386 B.n29 585
R226 B.n385 B.n28 585
R227 B.n427 B.n28 585
R228 B.n384 B.n27 585
R229 B.n428 B.n27 585
R230 B.n383 B.n26 585
R231 B.n429 B.n26 585
R232 B.n382 B.n381 585
R233 B.n381 B.n25 585
R234 B.n380 B.n21 585
R235 B.n435 B.n21 585
R236 B.n379 B.n20 585
R237 B.n436 B.n20 585
R238 B.n378 B.n19 585
R239 B.n437 B.n19 585
R240 B.n377 B.n376 585
R241 B.n376 B.n15 585
R242 B.n375 B.n14 585
R243 B.n443 B.n14 585
R244 B.n374 B.n13 585
R245 B.n444 B.n13 585
R246 B.n373 B.n12 585
R247 B.n445 B.n12 585
R248 B.n372 B.n371 585
R249 B.n371 B.n8 585
R250 B.n370 B.n7 585
R251 B.n451 B.n7 585
R252 B.n369 B.n6 585
R253 B.n452 B.n6 585
R254 B.n368 B.n5 585
R255 B.n453 B.n5 585
R256 B.n367 B.n366 585
R257 B.n366 B.n4 585
R258 B.n365 B.n146 585
R259 B.n365 B.n364 585
R260 B.n355 B.n147 585
R261 B.n148 B.n147 585
R262 B.n357 B.n356 585
R263 B.n358 B.n357 585
R264 B.n354 B.n152 585
R265 B.n156 B.n152 585
R266 B.n353 B.n352 585
R267 B.n352 B.n351 585
R268 B.n154 B.n153 585
R269 B.n155 B.n154 585
R270 B.n344 B.n343 585
R271 B.n345 B.n344 585
R272 B.n342 B.n161 585
R273 B.n161 B.n160 585
R274 B.n341 B.n340 585
R275 B.n340 B.n339 585
R276 B.n163 B.n162 585
R277 B.n332 B.n163 585
R278 B.n331 B.n330 585
R279 B.n333 B.n331 585
R280 B.n329 B.n168 585
R281 B.n168 B.n167 585
R282 B.n328 B.n327 585
R283 B.n327 B.n326 585
R284 B.n170 B.n169 585
R285 B.n171 B.n170 585
R286 B.n319 B.n318 585
R287 B.n320 B.n319 585
R288 B.n317 B.n176 585
R289 B.n176 B.n175 585
R290 B.n316 B.n315 585
R291 B.n315 B.n314 585
R292 B.n178 B.n177 585
R293 B.t5 B.n178 585
R294 B.n307 B.n306 585
R295 B.n308 B.n307 585
R296 B.n305 B.n183 585
R297 B.n183 B.n182 585
R298 B.n304 B.n303 585
R299 B.n303 B.n302 585
R300 B.n185 B.n184 585
R301 B.n186 B.n185 585
R302 B.n295 B.n294 585
R303 B.n296 B.n295 585
R304 B.n293 B.n191 585
R305 B.n191 B.n190 585
R306 B.n288 B.n287 585
R307 B.n286 B.n212 585
R308 B.n285 B.n211 585
R309 B.n290 B.n211 585
R310 B.n284 B.n283 585
R311 B.n282 B.n281 585
R312 B.n280 B.n279 585
R313 B.n278 B.n277 585
R314 B.n276 B.n275 585
R315 B.n274 B.n273 585
R316 B.n272 B.n271 585
R317 B.n270 B.n269 585
R318 B.n268 B.n267 585
R319 B.n266 B.n265 585
R320 B.n264 B.n263 585
R321 B.n261 B.n260 585
R322 B.n259 B.n258 585
R323 B.n257 B.n256 585
R324 B.n255 B.n254 585
R325 B.n253 B.n252 585
R326 B.n251 B.n250 585
R327 B.n249 B.n248 585
R328 B.n247 B.n246 585
R329 B.n245 B.n244 585
R330 B.n243 B.n242 585
R331 B.n240 B.n239 585
R332 B.n238 B.n237 585
R333 B.n236 B.n235 585
R334 B.n234 B.n233 585
R335 B.n232 B.n231 585
R336 B.n230 B.n229 585
R337 B.n228 B.n227 585
R338 B.n226 B.n225 585
R339 B.n224 B.n223 585
R340 B.n222 B.n221 585
R341 B.n220 B.n219 585
R342 B.n218 B.n217 585
R343 B.n193 B.n192 585
R344 B.n292 B.n291 585
R345 B.n291 B.n290 585
R346 B.n189 B.n188 585
R347 B.n190 B.n189 585
R348 B.n298 B.n297 585
R349 B.n297 B.n296 585
R350 B.n299 B.n187 585
R351 B.n187 B.n186 585
R352 B.n301 B.n300 585
R353 B.n302 B.n301 585
R354 B.n181 B.n180 585
R355 B.n182 B.n181 585
R356 B.n310 B.n309 585
R357 B.n309 B.n308 585
R358 B.n311 B.n179 585
R359 B.n179 B.t5 585
R360 B.n313 B.n312 585
R361 B.n314 B.n313 585
R362 B.n174 B.n173 585
R363 B.n175 B.n174 585
R364 B.n322 B.n321 585
R365 B.n321 B.n320 585
R366 B.n323 B.n172 585
R367 B.n172 B.n171 585
R368 B.n325 B.n324 585
R369 B.n326 B.n325 585
R370 B.n166 B.n165 585
R371 B.n167 B.n166 585
R372 B.n335 B.n334 585
R373 B.n334 B.n333 585
R374 B.n336 B.n164 585
R375 B.n332 B.n164 585
R376 B.n338 B.n337 585
R377 B.n339 B.n338 585
R378 B.n159 B.n158 585
R379 B.n160 B.n159 585
R380 B.n347 B.n346 585
R381 B.n346 B.n345 585
R382 B.n348 B.n157 585
R383 B.n157 B.n155 585
R384 B.n350 B.n349 585
R385 B.n351 B.n350 585
R386 B.n151 B.n150 585
R387 B.n156 B.n151 585
R388 B.n360 B.n359 585
R389 B.n359 B.n358 585
R390 B.n361 B.n149 585
R391 B.n149 B.n148 585
R392 B.n363 B.n362 585
R393 B.n364 B.n363 585
R394 B.n2 B.n0 585
R395 B.n4 B.n2 585
R396 B.n3 B.n1 585
R397 B.n452 B.n3 585
R398 B.n450 B.n449 585
R399 B.n451 B.n450 585
R400 B.n448 B.n9 585
R401 B.n9 B.n8 585
R402 B.n447 B.n446 585
R403 B.n446 B.n445 585
R404 B.n11 B.n10 585
R405 B.n444 B.n11 585
R406 B.n442 B.n441 585
R407 B.n443 B.n442 585
R408 B.n440 B.n16 585
R409 B.n16 B.n15 585
R410 B.n439 B.n438 585
R411 B.n438 B.n437 585
R412 B.n18 B.n17 585
R413 B.n436 B.n18 585
R414 B.n434 B.n433 585
R415 B.n435 B.n434 585
R416 B.n432 B.n22 585
R417 B.n25 B.n22 585
R418 B.n431 B.n430 585
R419 B.n430 B.n429 585
R420 B.n24 B.n23 585
R421 B.n428 B.n24 585
R422 B.n426 B.n425 585
R423 B.n427 B.n426 585
R424 B.n424 B.n30 585
R425 B.n30 B.n29 585
R426 B.n423 B.n422 585
R427 B.n422 B.n421 585
R428 B.n32 B.n31 585
R429 B.n420 B.n32 585
R430 B.n418 B.n417 585
R431 B.n419 B.n418 585
R432 B.n416 B.n36 585
R433 B.n36 B.t12 585
R434 B.n415 B.n414 585
R435 B.n414 B.n413 585
R436 B.n38 B.n37 585
R437 B.n412 B.n38 585
R438 B.n410 B.n409 585
R439 B.n411 B.n410 585
R440 B.n408 B.n43 585
R441 B.n43 B.n42 585
R442 B.n407 B.n406 585
R443 B.n406 B.n405 585
R444 B.n45 B.n44 585
R445 B.n404 B.n45 585
R446 B.n455 B.n454 585
R447 B.n454 B.n453 585
R448 B.n288 B.n189 530.939
R449 B.n73 B.n45 530.939
R450 B.n291 B.n191 530.939
R451 B.n401 B.n47 530.939
R452 B.n403 B.n402 256.663
R453 B.n403 B.n65 256.663
R454 B.n403 B.n64 256.663
R455 B.n403 B.n63 256.663
R456 B.n403 B.n62 256.663
R457 B.n403 B.n61 256.663
R458 B.n403 B.n60 256.663
R459 B.n403 B.n59 256.663
R460 B.n403 B.n58 256.663
R461 B.n403 B.n57 256.663
R462 B.n403 B.n56 256.663
R463 B.n403 B.n55 256.663
R464 B.n403 B.n54 256.663
R465 B.n403 B.n53 256.663
R466 B.n403 B.n52 256.663
R467 B.n403 B.n51 256.663
R468 B.n403 B.n50 256.663
R469 B.n403 B.n49 256.663
R470 B.n403 B.n48 256.663
R471 B.n290 B.n289 256.663
R472 B.n290 B.n194 256.663
R473 B.n290 B.n195 256.663
R474 B.n290 B.n196 256.663
R475 B.n290 B.n197 256.663
R476 B.n290 B.n198 256.663
R477 B.n290 B.n199 256.663
R478 B.n290 B.n200 256.663
R479 B.n290 B.n201 256.663
R480 B.n290 B.n202 256.663
R481 B.n290 B.n203 256.663
R482 B.n290 B.n204 256.663
R483 B.n290 B.n205 256.663
R484 B.n290 B.n206 256.663
R485 B.n290 B.n207 256.663
R486 B.n290 B.n208 256.663
R487 B.n290 B.n209 256.663
R488 B.n290 B.n210 256.663
R489 B.n215 B.t4 246.463
R490 B.n213 B.t8 246.463
R491 B.n70 B.t15 246.463
R492 B.n67 B.t11 246.463
R493 B.n290 B.n190 183.448
R494 B.n404 B.n403 183.448
R495 B.n215 B.t7 164.008
R496 B.n67 B.t13 164.008
R497 B.n213 B.t10 164.008
R498 B.n70 B.t16 164.008
R499 B.n297 B.n189 163.367
R500 B.n297 B.n187 163.367
R501 B.n301 B.n187 163.367
R502 B.n301 B.n181 163.367
R503 B.n309 B.n181 163.367
R504 B.n309 B.n179 163.367
R505 B.n313 B.n179 163.367
R506 B.n313 B.n174 163.367
R507 B.n321 B.n174 163.367
R508 B.n321 B.n172 163.367
R509 B.n325 B.n172 163.367
R510 B.n325 B.n166 163.367
R511 B.n334 B.n166 163.367
R512 B.n334 B.n164 163.367
R513 B.n338 B.n164 163.367
R514 B.n338 B.n159 163.367
R515 B.n346 B.n159 163.367
R516 B.n346 B.n157 163.367
R517 B.n350 B.n157 163.367
R518 B.n350 B.n151 163.367
R519 B.n359 B.n151 163.367
R520 B.n359 B.n149 163.367
R521 B.n363 B.n149 163.367
R522 B.n363 B.n2 163.367
R523 B.n454 B.n2 163.367
R524 B.n454 B.n3 163.367
R525 B.n450 B.n3 163.367
R526 B.n450 B.n9 163.367
R527 B.n446 B.n9 163.367
R528 B.n446 B.n11 163.367
R529 B.n442 B.n11 163.367
R530 B.n442 B.n16 163.367
R531 B.n438 B.n16 163.367
R532 B.n438 B.n18 163.367
R533 B.n434 B.n18 163.367
R534 B.n434 B.n22 163.367
R535 B.n430 B.n22 163.367
R536 B.n430 B.n24 163.367
R537 B.n426 B.n24 163.367
R538 B.n426 B.n30 163.367
R539 B.n422 B.n30 163.367
R540 B.n422 B.n32 163.367
R541 B.n418 B.n32 163.367
R542 B.n418 B.n36 163.367
R543 B.n414 B.n36 163.367
R544 B.n414 B.n38 163.367
R545 B.n410 B.n38 163.367
R546 B.n410 B.n43 163.367
R547 B.n406 B.n43 163.367
R548 B.n406 B.n45 163.367
R549 B.n212 B.n211 163.367
R550 B.n283 B.n211 163.367
R551 B.n281 B.n280 163.367
R552 B.n277 B.n276 163.367
R553 B.n273 B.n272 163.367
R554 B.n269 B.n268 163.367
R555 B.n265 B.n264 163.367
R556 B.n260 B.n259 163.367
R557 B.n256 B.n255 163.367
R558 B.n252 B.n251 163.367
R559 B.n248 B.n247 163.367
R560 B.n244 B.n243 163.367
R561 B.n239 B.n238 163.367
R562 B.n235 B.n234 163.367
R563 B.n231 B.n230 163.367
R564 B.n227 B.n226 163.367
R565 B.n223 B.n222 163.367
R566 B.n219 B.n218 163.367
R567 B.n291 B.n193 163.367
R568 B.n295 B.n191 163.367
R569 B.n295 B.n185 163.367
R570 B.n303 B.n185 163.367
R571 B.n303 B.n183 163.367
R572 B.n307 B.n183 163.367
R573 B.n307 B.n178 163.367
R574 B.n315 B.n178 163.367
R575 B.n315 B.n176 163.367
R576 B.n319 B.n176 163.367
R577 B.n319 B.n170 163.367
R578 B.n327 B.n170 163.367
R579 B.n327 B.n168 163.367
R580 B.n331 B.n168 163.367
R581 B.n331 B.n163 163.367
R582 B.n340 B.n163 163.367
R583 B.n340 B.n161 163.367
R584 B.n344 B.n161 163.367
R585 B.n344 B.n154 163.367
R586 B.n352 B.n154 163.367
R587 B.n352 B.n152 163.367
R588 B.n357 B.n152 163.367
R589 B.n357 B.n147 163.367
R590 B.n365 B.n147 163.367
R591 B.n366 B.n365 163.367
R592 B.n366 B.n5 163.367
R593 B.n6 B.n5 163.367
R594 B.n7 B.n6 163.367
R595 B.n371 B.n7 163.367
R596 B.n371 B.n12 163.367
R597 B.n13 B.n12 163.367
R598 B.n14 B.n13 163.367
R599 B.n376 B.n14 163.367
R600 B.n376 B.n19 163.367
R601 B.n20 B.n19 163.367
R602 B.n21 B.n20 163.367
R603 B.n381 B.n21 163.367
R604 B.n381 B.n26 163.367
R605 B.n27 B.n26 163.367
R606 B.n28 B.n27 163.367
R607 B.n386 B.n28 163.367
R608 B.n386 B.n33 163.367
R609 B.n34 B.n33 163.367
R610 B.n35 B.n34 163.367
R611 B.n391 B.n35 163.367
R612 B.n391 B.n39 163.367
R613 B.n40 B.n39 163.367
R614 B.n41 B.n40 163.367
R615 B.n396 B.n41 163.367
R616 B.n396 B.n46 163.367
R617 B.n47 B.n46 163.367
R618 B.n77 B.n76 163.367
R619 B.n81 B.n80 163.367
R620 B.n85 B.n84 163.367
R621 B.n89 B.n88 163.367
R622 B.n93 B.n92 163.367
R623 B.n97 B.n96 163.367
R624 B.n101 B.n100 163.367
R625 B.n105 B.n104 163.367
R626 B.n109 B.n108 163.367
R627 B.n113 B.n112 163.367
R628 B.n117 B.n116 163.367
R629 B.n121 B.n120 163.367
R630 B.n125 B.n124 163.367
R631 B.n129 B.n128 163.367
R632 B.n133 B.n132 163.367
R633 B.n137 B.n136 163.367
R634 B.n141 B.n140 163.367
R635 B.n143 B.n66 163.367
R636 B.n216 B.t6 126.578
R637 B.n68 B.t14 126.578
R638 B.n214 B.t9 126.578
R639 B.n71 B.t17 126.578
R640 B.n296 B.n190 93.7936
R641 B.n296 B.n186 93.7936
R642 B.n302 B.n186 93.7936
R643 B.n302 B.n182 93.7936
R644 B.n308 B.n182 93.7936
R645 B.n308 B.t5 93.7936
R646 B.n314 B.t5 93.7936
R647 B.n314 B.n175 93.7936
R648 B.n320 B.n175 93.7936
R649 B.n320 B.n171 93.7936
R650 B.n326 B.n171 93.7936
R651 B.n326 B.n167 93.7936
R652 B.n333 B.n167 93.7936
R653 B.n333 B.n332 93.7936
R654 B.n339 B.n160 93.7936
R655 B.n345 B.n160 93.7936
R656 B.n345 B.n155 93.7936
R657 B.n351 B.n155 93.7936
R658 B.n351 B.n156 93.7936
R659 B.n358 B.n148 93.7936
R660 B.n364 B.n148 93.7936
R661 B.n364 B.n4 93.7936
R662 B.n453 B.n4 93.7936
R663 B.n453 B.n452 93.7936
R664 B.n452 B.n451 93.7936
R665 B.n451 B.n8 93.7936
R666 B.n445 B.n8 93.7936
R667 B.n444 B.n443 93.7936
R668 B.n443 B.n15 93.7936
R669 B.n437 B.n15 93.7936
R670 B.n437 B.n436 93.7936
R671 B.n436 B.n435 93.7936
R672 B.n429 B.n25 93.7936
R673 B.n429 B.n428 93.7936
R674 B.n428 B.n427 93.7936
R675 B.n427 B.n29 93.7936
R676 B.n421 B.n29 93.7936
R677 B.n421 B.n420 93.7936
R678 B.n420 B.n419 93.7936
R679 B.n419 B.t12 93.7936
R680 B.n413 B.t12 93.7936
R681 B.n413 B.n412 93.7936
R682 B.n412 B.n411 93.7936
R683 B.n411 B.n42 93.7936
R684 B.n405 B.n42 93.7936
R685 B.n405 B.n404 93.7936
R686 B.n332 B.t2 82.7591
R687 B.n25 B.t0 82.7591
R688 B.n289 B.n288 71.676
R689 B.n283 B.n194 71.676
R690 B.n280 B.n195 71.676
R691 B.n276 B.n196 71.676
R692 B.n272 B.n197 71.676
R693 B.n268 B.n198 71.676
R694 B.n264 B.n199 71.676
R695 B.n259 B.n200 71.676
R696 B.n255 B.n201 71.676
R697 B.n251 B.n202 71.676
R698 B.n247 B.n203 71.676
R699 B.n243 B.n204 71.676
R700 B.n238 B.n205 71.676
R701 B.n234 B.n206 71.676
R702 B.n230 B.n207 71.676
R703 B.n226 B.n208 71.676
R704 B.n222 B.n209 71.676
R705 B.n218 B.n210 71.676
R706 B.n73 B.n48 71.676
R707 B.n77 B.n49 71.676
R708 B.n81 B.n50 71.676
R709 B.n85 B.n51 71.676
R710 B.n89 B.n52 71.676
R711 B.n93 B.n53 71.676
R712 B.n97 B.n54 71.676
R713 B.n101 B.n55 71.676
R714 B.n105 B.n56 71.676
R715 B.n109 B.n57 71.676
R716 B.n113 B.n58 71.676
R717 B.n117 B.n59 71.676
R718 B.n121 B.n60 71.676
R719 B.n125 B.n61 71.676
R720 B.n129 B.n62 71.676
R721 B.n133 B.n63 71.676
R722 B.n137 B.n64 71.676
R723 B.n141 B.n65 71.676
R724 B.n402 B.n66 71.676
R725 B.n402 B.n401 71.676
R726 B.n143 B.n65 71.676
R727 B.n140 B.n64 71.676
R728 B.n136 B.n63 71.676
R729 B.n132 B.n62 71.676
R730 B.n128 B.n61 71.676
R731 B.n124 B.n60 71.676
R732 B.n120 B.n59 71.676
R733 B.n116 B.n58 71.676
R734 B.n112 B.n57 71.676
R735 B.n108 B.n56 71.676
R736 B.n104 B.n55 71.676
R737 B.n100 B.n54 71.676
R738 B.n96 B.n53 71.676
R739 B.n92 B.n52 71.676
R740 B.n88 B.n51 71.676
R741 B.n84 B.n50 71.676
R742 B.n80 B.n49 71.676
R743 B.n76 B.n48 71.676
R744 B.n289 B.n212 71.676
R745 B.n281 B.n194 71.676
R746 B.n277 B.n195 71.676
R747 B.n273 B.n196 71.676
R748 B.n269 B.n197 71.676
R749 B.n265 B.n198 71.676
R750 B.n260 B.n199 71.676
R751 B.n256 B.n200 71.676
R752 B.n252 B.n201 71.676
R753 B.n248 B.n202 71.676
R754 B.n244 B.n203 71.676
R755 B.n239 B.n204 71.676
R756 B.n235 B.n205 71.676
R757 B.n231 B.n206 71.676
R758 B.n227 B.n207 71.676
R759 B.n223 B.n208 71.676
R760 B.n219 B.n209 71.676
R761 B.n210 B.n193 71.676
R762 B.n241 B.n216 59.5399
R763 B.n262 B.n214 59.5399
R764 B.n72 B.n71 59.5399
R765 B.n69 B.n68 59.5399
R766 B.n156 B.t3 52.4143
R767 B.t1 B.n444 52.4143
R768 B.n358 B.t3 41.3798
R769 B.n445 B.t1 41.3798
R770 B.n216 B.n215 37.4308
R771 B.n214 B.n213 37.4308
R772 B.n71 B.n70 37.4308
R773 B.n68 B.n67 37.4308
R774 B.n74 B.n44 34.4981
R775 B.n400 B.n399 34.4981
R776 B.n293 B.n292 34.4981
R777 B.n287 B.n188 34.4981
R778 B B.n455 18.0485
R779 B.n339 B.t2 11.035
R780 B.n435 B.t0 11.035
R781 B.n75 B.n74 10.6151
R782 B.n78 B.n75 10.6151
R783 B.n79 B.n78 10.6151
R784 B.n82 B.n79 10.6151
R785 B.n83 B.n82 10.6151
R786 B.n86 B.n83 10.6151
R787 B.n87 B.n86 10.6151
R788 B.n90 B.n87 10.6151
R789 B.n91 B.n90 10.6151
R790 B.n94 B.n91 10.6151
R791 B.n95 B.n94 10.6151
R792 B.n98 B.n95 10.6151
R793 B.n99 B.n98 10.6151
R794 B.n103 B.n102 10.6151
R795 B.n106 B.n103 10.6151
R796 B.n107 B.n106 10.6151
R797 B.n110 B.n107 10.6151
R798 B.n111 B.n110 10.6151
R799 B.n114 B.n111 10.6151
R800 B.n115 B.n114 10.6151
R801 B.n118 B.n115 10.6151
R802 B.n119 B.n118 10.6151
R803 B.n123 B.n122 10.6151
R804 B.n126 B.n123 10.6151
R805 B.n127 B.n126 10.6151
R806 B.n130 B.n127 10.6151
R807 B.n131 B.n130 10.6151
R808 B.n134 B.n131 10.6151
R809 B.n135 B.n134 10.6151
R810 B.n138 B.n135 10.6151
R811 B.n139 B.n138 10.6151
R812 B.n142 B.n139 10.6151
R813 B.n144 B.n142 10.6151
R814 B.n145 B.n144 10.6151
R815 B.n400 B.n145 10.6151
R816 B.n294 B.n293 10.6151
R817 B.n294 B.n184 10.6151
R818 B.n304 B.n184 10.6151
R819 B.n305 B.n304 10.6151
R820 B.n306 B.n305 10.6151
R821 B.n306 B.n177 10.6151
R822 B.n316 B.n177 10.6151
R823 B.n317 B.n316 10.6151
R824 B.n318 B.n317 10.6151
R825 B.n318 B.n169 10.6151
R826 B.n328 B.n169 10.6151
R827 B.n329 B.n328 10.6151
R828 B.n330 B.n329 10.6151
R829 B.n330 B.n162 10.6151
R830 B.n341 B.n162 10.6151
R831 B.n342 B.n341 10.6151
R832 B.n343 B.n342 10.6151
R833 B.n343 B.n153 10.6151
R834 B.n353 B.n153 10.6151
R835 B.n354 B.n353 10.6151
R836 B.n356 B.n354 10.6151
R837 B.n356 B.n355 10.6151
R838 B.n355 B.n146 10.6151
R839 B.n367 B.n146 10.6151
R840 B.n368 B.n367 10.6151
R841 B.n369 B.n368 10.6151
R842 B.n370 B.n369 10.6151
R843 B.n372 B.n370 10.6151
R844 B.n373 B.n372 10.6151
R845 B.n374 B.n373 10.6151
R846 B.n375 B.n374 10.6151
R847 B.n377 B.n375 10.6151
R848 B.n378 B.n377 10.6151
R849 B.n379 B.n378 10.6151
R850 B.n380 B.n379 10.6151
R851 B.n382 B.n380 10.6151
R852 B.n383 B.n382 10.6151
R853 B.n384 B.n383 10.6151
R854 B.n385 B.n384 10.6151
R855 B.n387 B.n385 10.6151
R856 B.n388 B.n387 10.6151
R857 B.n389 B.n388 10.6151
R858 B.n390 B.n389 10.6151
R859 B.n392 B.n390 10.6151
R860 B.n393 B.n392 10.6151
R861 B.n394 B.n393 10.6151
R862 B.n395 B.n394 10.6151
R863 B.n397 B.n395 10.6151
R864 B.n398 B.n397 10.6151
R865 B.n399 B.n398 10.6151
R866 B.n287 B.n286 10.6151
R867 B.n286 B.n285 10.6151
R868 B.n285 B.n284 10.6151
R869 B.n284 B.n282 10.6151
R870 B.n282 B.n279 10.6151
R871 B.n279 B.n278 10.6151
R872 B.n278 B.n275 10.6151
R873 B.n275 B.n274 10.6151
R874 B.n274 B.n271 10.6151
R875 B.n271 B.n270 10.6151
R876 B.n270 B.n267 10.6151
R877 B.n267 B.n266 10.6151
R878 B.n266 B.n263 10.6151
R879 B.n261 B.n258 10.6151
R880 B.n258 B.n257 10.6151
R881 B.n257 B.n254 10.6151
R882 B.n254 B.n253 10.6151
R883 B.n253 B.n250 10.6151
R884 B.n250 B.n249 10.6151
R885 B.n249 B.n246 10.6151
R886 B.n246 B.n245 10.6151
R887 B.n245 B.n242 10.6151
R888 B.n240 B.n237 10.6151
R889 B.n237 B.n236 10.6151
R890 B.n236 B.n233 10.6151
R891 B.n233 B.n232 10.6151
R892 B.n232 B.n229 10.6151
R893 B.n229 B.n228 10.6151
R894 B.n228 B.n225 10.6151
R895 B.n225 B.n224 10.6151
R896 B.n224 B.n221 10.6151
R897 B.n221 B.n220 10.6151
R898 B.n220 B.n217 10.6151
R899 B.n217 B.n192 10.6151
R900 B.n292 B.n192 10.6151
R901 B.n298 B.n188 10.6151
R902 B.n299 B.n298 10.6151
R903 B.n300 B.n299 10.6151
R904 B.n300 B.n180 10.6151
R905 B.n310 B.n180 10.6151
R906 B.n311 B.n310 10.6151
R907 B.n312 B.n311 10.6151
R908 B.n312 B.n173 10.6151
R909 B.n322 B.n173 10.6151
R910 B.n323 B.n322 10.6151
R911 B.n324 B.n323 10.6151
R912 B.n324 B.n165 10.6151
R913 B.n335 B.n165 10.6151
R914 B.n336 B.n335 10.6151
R915 B.n337 B.n336 10.6151
R916 B.n337 B.n158 10.6151
R917 B.n347 B.n158 10.6151
R918 B.n348 B.n347 10.6151
R919 B.n349 B.n348 10.6151
R920 B.n349 B.n150 10.6151
R921 B.n360 B.n150 10.6151
R922 B.n361 B.n360 10.6151
R923 B.n362 B.n361 10.6151
R924 B.n362 B.n0 10.6151
R925 B.n449 B.n1 10.6151
R926 B.n449 B.n448 10.6151
R927 B.n448 B.n447 10.6151
R928 B.n447 B.n10 10.6151
R929 B.n441 B.n10 10.6151
R930 B.n441 B.n440 10.6151
R931 B.n440 B.n439 10.6151
R932 B.n439 B.n17 10.6151
R933 B.n433 B.n17 10.6151
R934 B.n433 B.n432 10.6151
R935 B.n432 B.n431 10.6151
R936 B.n431 B.n23 10.6151
R937 B.n425 B.n23 10.6151
R938 B.n425 B.n424 10.6151
R939 B.n424 B.n423 10.6151
R940 B.n423 B.n31 10.6151
R941 B.n417 B.n31 10.6151
R942 B.n417 B.n416 10.6151
R943 B.n416 B.n415 10.6151
R944 B.n415 B.n37 10.6151
R945 B.n409 B.n37 10.6151
R946 B.n409 B.n408 10.6151
R947 B.n408 B.n407 10.6151
R948 B.n407 B.n44 10.6151
R949 B.n99 B.n72 9.36635
R950 B.n122 B.n69 9.36635
R951 B.n263 B.n262 9.36635
R952 B.n241 B.n240 9.36635
R953 B.n455 B.n0 2.81026
R954 B.n455 B.n1 2.81026
R955 B.n102 B.n72 1.24928
R956 B.n119 B.n69 1.24928
R957 B.n262 B.n261 1.24928
R958 B.n242 B.n241 1.24928
R959 VP.n4 VP.n3 175.317
R960 VP.n12 VP.n11 175.317
R961 VP.n10 VP.n0 161.3
R962 VP.n9 VP.n8 161.3
R963 VP.n7 VP.n1 161.3
R964 VP.n6 VP.n5 161.3
R965 VP.n2 VP.t0 78.5491
R966 VP.n2 VP.t3 78.2235
R967 VP.n9 VP.n1 56.5617
R968 VP.n3 VP.n2 48.8436
R969 VP.n4 VP.t2 40.6693
R970 VP.n11 VP.t1 40.6693
R971 VP.n5 VP.n1 24.5923
R972 VP.n10 VP.n9 24.5923
R973 VP.n5 VP.n4 10.575
R974 VP.n11 VP.n10 10.575
R975 VP.n6 VP.n3 0.189894
R976 VP.n7 VP.n6 0.189894
R977 VP.n8 VP.n7 0.189894
R978 VP.n8 VP.n0 0.189894
R979 VP.n12 VP.n0 0.189894
R980 VP VP.n12 0.0516364
R981 VDD1 VDD1.n1 116.814
R982 VDD1 VDD1.n0 85.3127
R983 VDD1.n0 VDD1.t3 7.33383
R984 VDD1.n0 VDD1.t0 7.33383
R985 VDD1.n1 VDD1.t1 7.33383
R986 VDD1.n1 VDD1.t2 7.33383
C0 VP VTAIL 1.4865f
C1 VTAIL VN 1.4724f
C2 VDD2 VTAIL 2.81198f
C3 VP VDD1 1.37717f
C4 VN VDD1 0.153679f
C5 VDD2 VDD1 0.784429f
C6 VP VN 3.74935f
C7 VDD2 VN 1.19514f
C8 VDD2 VP 0.336856f
C9 VTAIL VDD1 2.76448f
C10 VDD2 B 2.429552f
C11 VDD1 B 4.42615f
C12 VTAIL B 3.721051f
C13 VN B 7.25193f
C14 VP B 5.997206f
C15 VDD1.t3 B 0.039992f
C16 VDD1.t0 B 0.039992f
C17 VDD1.n0 B 0.279475f
C18 VDD1.t1 B 0.039992f
C19 VDD1.t2 B 0.039992f
C20 VDD1.n1 B 0.478742f
C21 VP.n0 B 0.02337f
C22 VP.t1 B 0.248006f
C23 VP.n1 B 0.033972f
C24 VP.t0 B 0.351936f
C25 VP.t3 B 0.35106f
C26 VP.n2 B 0.909322f
C27 VP.n3 B 0.996445f
C28 VP.t2 B 0.248006f
C29 VP.n4 B 0.167981f
C30 VP.n5 B 0.031143f
C31 VP.n6 B 0.02337f
C32 VP.n7 B 0.02337f
C33 VP.n8 B 0.02337f
C34 VP.n9 B 0.033972f
C35 VP.n10 B 0.031143f
C36 VP.n11 B 0.167981f
C37 VP.n12 B 0.022654f
C38 VTAIL.n0 B 0.022105f
C39 VTAIL.n1 B 0.13134f
C40 VTAIL.n2 B 0.008064f
C41 VTAIL.t4 B 0.034835f
C42 VTAIL.n3 B 0.056609f
C43 VTAIL.n4 B 0.01305f
C44 VTAIL.n5 B 0.014295f
C45 VTAIL.n6 B 0.043052f
C46 VTAIL.n7 B 0.008538f
C47 VTAIL.n8 B 0.008064f
C48 VTAIL.n9 B 0.033457f
C49 VTAIL.n10 B 0.024235f
C50 VTAIL.n11 B 0.077881f
C51 VTAIL.n12 B 0.022105f
C52 VTAIL.n13 B 0.13134f
C53 VTAIL.n14 B 0.008064f
C54 VTAIL.t3 B 0.034835f
C55 VTAIL.n15 B 0.056609f
C56 VTAIL.n16 B 0.01305f
C57 VTAIL.n17 B 0.014295f
C58 VTAIL.n18 B 0.043052f
C59 VTAIL.n19 B 0.008538f
C60 VTAIL.n20 B 0.008064f
C61 VTAIL.n21 B 0.033457f
C62 VTAIL.n22 B 0.024235f
C63 VTAIL.n23 B 0.115292f
C64 VTAIL.n24 B 0.022105f
C65 VTAIL.n25 B 0.13134f
C66 VTAIL.n26 B 0.008064f
C67 VTAIL.t2 B 0.034835f
C68 VTAIL.n27 B 0.056609f
C69 VTAIL.n28 B 0.01305f
C70 VTAIL.n29 B 0.014295f
C71 VTAIL.n30 B 0.043052f
C72 VTAIL.n31 B 0.008538f
C73 VTAIL.n32 B 0.008064f
C74 VTAIL.n33 B 0.033457f
C75 VTAIL.n34 B 0.024235f
C76 VTAIL.n35 B 0.489419f
C77 VTAIL.n36 B 0.022105f
C78 VTAIL.n37 B 0.13134f
C79 VTAIL.n38 B 0.008064f
C80 VTAIL.t7 B 0.034835f
C81 VTAIL.n39 B 0.056609f
C82 VTAIL.n40 B 0.01305f
C83 VTAIL.n41 B 0.014295f
C84 VTAIL.n42 B 0.043052f
C85 VTAIL.n43 B 0.008538f
C86 VTAIL.n44 B 0.008064f
C87 VTAIL.n45 B 0.033457f
C88 VTAIL.n46 B 0.024235f
C89 VTAIL.n47 B 0.489419f
C90 VTAIL.n48 B 0.022105f
C91 VTAIL.n49 B 0.13134f
C92 VTAIL.n50 B 0.008064f
C93 VTAIL.t5 B 0.034835f
C94 VTAIL.n51 B 0.056609f
C95 VTAIL.n52 B 0.01305f
C96 VTAIL.n53 B 0.014295f
C97 VTAIL.n54 B 0.043052f
C98 VTAIL.n55 B 0.008538f
C99 VTAIL.n56 B 0.008064f
C100 VTAIL.n57 B 0.033457f
C101 VTAIL.n58 B 0.024235f
C102 VTAIL.n59 B 0.115292f
C103 VTAIL.n60 B 0.022105f
C104 VTAIL.n61 B 0.13134f
C105 VTAIL.n62 B 0.008064f
C106 VTAIL.t1 B 0.034835f
C107 VTAIL.n63 B 0.056609f
C108 VTAIL.n64 B 0.01305f
C109 VTAIL.n65 B 0.014295f
C110 VTAIL.n66 B 0.043052f
C111 VTAIL.n67 B 0.008538f
C112 VTAIL.n68 B 0.008064f
C113 VTAIL.n69 B 0.033457f
C114 VTAIL.n70 B 0.024235f
C115 VTAIL.n71 B 0.115292f
C116 VTAIL.n72 B 0.022105f
C117 VTAIL.n73 B 0.13134f
C118 VTAIL.n74 B 0.008064f
C119 VTAIL.t0 B 0.034835f
C120 VTAIL.n75 B 0.056609f
C121 VTAIL.n76 B 0.01305f
C122 VTAIL.n77 B 0.014295f
C123 VTAIL.n78 B 0.043052f
C124 VTAIL.n79 B 0.008538f
C125 VTAIL.n80 B 0.008064f
C126 VTAIL.n81 B 0.033457f
C127 VTAIL.n82 B 0.024235f
C128 VTAIL.n83 B 0.489419f
C129 VTAIL.n84 B 0.022105f
C130 VTAIL.n85 B 0.13134f
C131 VTAIL.n86 B 0.008064f
C132 VTAIL.t6 B 0.034835f
C133 VTAIL.n87 B 0.056609f
C134 VTAIL.n88 B 0.01305f
C135 VTAIL.n89 B 0.014295f
C136 VTAIL.n90 B 0.043052f
C137 VTAIL.n91 B 0.008538f
C138 VTAIL.n92 B 0.008064f
C139 VTAIL.n93 B 0.033457f
C140 VTAIL.n94 B 0.024235f
C141 VTAIL.n95 B 0.44638f
C142 VDD2.t0 B 0.041006f
C143 VDD2.t2 B 0.041006f
C144 VDD2.n0 B 0.477891f
C145 VDD2.t1 B 0.041006f
C146 VDD2.t3 B 0.041006f
C147 VDD2.n1 B 0.286378f
C148 VDD2.n2 B 1.76454f
C149 VN.t3 B 0.348839f
C150 VN.t1 B 0.34797f
C151 VN.n0 B 0.260081f
C152 VN.t2 B 0.348839f
C153 VN.t0 B 0.34797f
C154 VN.n1 B 0.914468f
.ends

