* NGSPICE file created from opamp_sample_0010.ext - technology: sky130A

.subckt opamp_sample_0010 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t166 GND.t163 GND.t165 GND.t164 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=0 ps=0 w=4.7 l=5.88
X1 VOUT.t15 CS_BIAS.t8 GND.t25 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X2 GND.t8 CS_BIAS.t9 VOUT.t14 GND.t6 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X3 VN.t6 GND.t160 GND.t162 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 VDD.t133 a_n11634_10845.t22 a_n11778_11043.t16 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X5 VOUT.t26 a_n8732_9422.t0 sky130_fd_pr__cap_mim_m3_1 l=18.34 w=7.84
X6 a_n3337_n4072.t3 DIFFPAIR_BIAS.t8 GND.t27 GND.t26 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X7 VOUT.t13 CS_BIAS.t10 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X8 a_n11634_10845.t21 VP.t7 a_n3337_n4072.t7 GND.t169 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=5.1336 ps=15.7 w=7.13 l=2.31
X9 VOUT.t25 a_n17232_8522.t12 VDD.t146 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X10 GND.t159 GND.t157 GND.t158 GND.t84 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X11 a_n11778_11043.t12 a_n11634_10845.t3 a_n11634_10845.t4 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X12 GND.t156 GND.t153 GND.t155 GND.t154 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=0 ps=0 w=4.7 l=5.88
X13 GND.t116 GND.t114 VP.t6 GND.t115 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X14 VDD.t127 a_n11634_10845.t23 a_n8732_9422.t8 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X15 VDD.t91 VDD.t89 VDD.t90 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X16 a_n11778_11043.t17 a_n11634_10845.t24 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X17 VDD.t88 VDD.t86 VDD.t87 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X18 a_n11778_11043.t11 a_n11634_10845.t5 a_n11634_10845.t6 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X19 VN.t5 GND.t150 GND.t152 GND.t151 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X20 VN.t4 GND.t147 GND.t149 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X21 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X22 VDD.t85 VDD.t83 VDD.t84 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X23 a_n11634_10845.t14 a_n11634_10845.t13 a_n11778_11043.t10 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X24 a_n11778_11043.t13 a_n11634_10845.t25 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X25 GND.t146 GND.t144 GND.t145 GND.t63 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X26 VOUT.t24 a_n17232_8522.t13 VDD.t145 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X27 VDD.t82 VDD.t80 VDD.t81 VDD.t22 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X28 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t168 GND.t167 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X29 GND.t143 GND.t141 GND.t142 GND.t77 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=0 ps=0 w=7.13 l=2.31
X30 VDD.t79 VDD.t77 VDD.t78 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X31 VDD.t76 VDD.t74 VDD.t75 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X32 CS_BIAS.t7 CS_BIAS.t6 GND.t9 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X33 a_n11634_10845.t8 a_n11634_10845.t7 a_n11778_11043.t9 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X34 VDD.t125 a_n11634_10845.t26 a_n8732_9422.t7 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X35 VDD.t73 VDD.t71 VDD.t72 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X36 a_n3337_n4072.t2 DIFFPAIR_BIAS.t9 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X37 GND.t140 GND.t138 GND.t139 GND.t67 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X38 a_n3337_n4072.t1 DIFFPAIR_BIAS.t10 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X39 GND.t137 GND.t135 GND.t136 GND.t84 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X40 GND.t29 CS_BIAS.t11 VOUT.t12 GND.t6 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X41 GND.t134 GND.t132 VP.t5 GND.t133 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X42 GND.t131 GND.t129 GND.t130 GND.t63 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X43 GND.t7 CS_BIAS.t12 VOUT.t11 GND.t6 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X44 VDD.t70 VDD.t68 VDD.t69 VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X45 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X46 GND.t128 GND.t126 GND.t127 GND.t63 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X47 GND.t119 GND.t117 VN.t3 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X48 GND.t125 GND.t123 GND.t124 GND.t53 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X49 GND.t122 GND.t120 GND.t121 GND.t53 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X50 GND.t28 CS_BIAS.t4 CS_BIAS.t5 GND.t18 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X51 VDD.t123 a_n11634_10845.t27 a_n11778_11043.t15 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X52 VDD.t67 VDD.t65 VDD.t66 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X53 a_n11778_11043.t8 a_n11634_10845.t11 a_n11634_10845.t12 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X54 a_n17232_8522.t9 a_n11634_10845.t28 a_n8732_9422.t10 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X55 a_n17232_8522.t8 a_n11634_10845.t29 a_n8732_9422.t11 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X56 VDD.t64 VDD.t62 VDD.t63 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X57 a_11906_11043# a_11906_11043# a_11906_11043# VDD.t147 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=3.6864 ps=13.12 w=2.56 l=5.82
X58 a_n11778_11043.t7 a_n11634_10845.t19 a_n11634_10845.t20 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X59 GND.t110 GND.t108 VP.t4 GND.t109 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X60 GND.t113 GND.t111 GND.t112 GND.t43 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=0 ps=0 w=7.13 l=2.31
X61 VOUT.t10 CS_BIAS.t13 GND.t35 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X62 VDD.t61 VDD.t59 VDD.t60 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X63 VOUT.t23 a_n17232_8522.t14 VDD.t144 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X64 a_n11634_10845.t0 VP.t8 a_n3337_n4072.t4 GND.t23 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=5.1336 ps=15.7 w=7.13 l=2.31
X65 a_n17232_8522.t7 a_n11634_10845.t30 a_n8732_9422.t12 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X66 GND.t107 GND.t105 VN.t2 GND.t106 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X67 VDD.t58 VDD.t56 VDD.t57 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X68 GND.t104 GND.t102 GND.t103 GND.t67 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X69 a_n3337_n4072.t0 DIFFPAIR_BIAS.t11 GND.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X70 GND.t33 CS_BIAS.t14 VOUT.t9 GND.t18 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X71 a_n17232_8522.t6 a_n11634_10845.t31 a_n8732_9422.t13 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X72 VDD.t55 VDD.t53 VDD.t54 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X73 GND.t30 CS_BIAS.t15 VOUT.t8 GND.t18 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X74 a_n8732_9422.t18 a_n11634_10845.t32 a_n17232_8522.t5 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X75 VOUT.t22 a_n17232_8522.t15 VDD.t143 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X76 VDD.t118 a_n11634_10845.t33 a_n8732_9422.t6 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X77 VOUT.t21 a_n17232_8522.t16 VDD.t142 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X78 GND.t101 GND.t99 GND.t100 GND.t63 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X79 a_n8732_9422.t14 a_n11634_10845.t34 a_n17232_8522.t4 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X80 a_n8732_9422.t15 a_n11634_10845.t35 a_n17232_8522.t3 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X81 VOUT.t7 CS_BIAS.t16 GND.t36 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X82 GND.t98 GND.t96 GND.t97 GND.t84 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X83 VOUT.t20 a_n17232_8522.t17 VDD.t141 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X84 VOUT.t6 CS_BIAS.t17 GND.t24 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X85 VDD.t100 a_n11634_10845.t36 a_n8732_9422.t5 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X86 GND.t95 GND.t93 GND.t94 GND.t84 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X87 a_n17232_8522.t11 VN.t7 a_n3337_n4072.t5 GND.t169 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=5.1336 ps=15.7 w=7.13 l=2.31
X88 VP.t3 GND.t90 GND.t92 GND.t91 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X89 a_n11778_11043.t0 a_n11634_10845.t37 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X90 VP.t2 GND.t87 GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X91 a_n17232_8522.t2 a_n11634_10845.t38 a_n8732_9422.t16 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X92 a_n8732_9422.t4 a_n11634_10845.t39 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X93 GND.t86 GND.t83 GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X94 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X95 CS_BIAS.t3 CS_BIAS.t2 GND.t17 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X96 VDD.t48 VDD.t46 VDD.t47 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X97 VDD.t45 VDD.t42 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X98 a_n13358_11043# a_n13358_11043# a_n13358_11043# VDD.t134 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=3.6864 ps=13.12 w=2.56 l=5.82
X99 VDD.t41 VDD.t39 VDD.t40 VDD.t29 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X100 VOUT.t19 a_n17232_8522.t18 VDD.t140 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X101 GND.t82 GND.t80 GND.t81 GND.t53 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X102 VDD.t38 VDD.t36 VDD.t37 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X103 GND.t34 CS_BIAS.t18 VOUT.t5 GND.t18 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X104 GND.t31 CS_BIAS.t0 CS_BIAS.t1 GND.t6 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X105 a_n11634_10845.t10 a_n11634_10845.t9 a_n11778_11043.t6 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X106 a_n8732_9422.t3 a_n11634_10845.t40 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X107 GND.t79 GND.t76 GND.t78 GND.t77 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=0 ps=0 w=7.13 l=2.31
X108 VP.t1 GND.t46 GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X109 GND.t75 GND.t73 GND.t74 GND.t67 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X110 VDD.t35 VDD.t32 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X111 VDD.t31 VDD.t28 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X112 VDD.t27 VDD.t25 VDD.t26 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X113 GND.t72 GND.t70 GND.t71 GND.t67 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X114 a_n11778_11043.t5 a_n11634_10845.t1 a_n11634_10845.t2 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X115 VDD.t24 VDD.t21 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X116 GND.t69 GND.t66 GND.t68 GND.t67 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X117 a_n8732_9422.t17 a_n11634_10845.t41 a_n17232_8522.t1 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X118 GND.t22 CS_BIAS.t19 VOUT.t4 GND.t6 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X119 GND.t65 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X120 GND.t61 GND.t59 GND.t60 GND.t53 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X121 GND.t55 GND.t52 GND.t54 GND.t53 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=0 ps=0 w=5.91 l=4.37
X122 VDD.t106 a_n11634_10845.t42 a_n11778_11043.t14 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=1.8432 ps=6.56 w=2.56 l=5.82
X123 GND.t58 GND.t56 VN.t1 GND.t57 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X124 VDD.t20 VDD.t17 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0 ps=0 w=2.56 l=5.82
X125 VOUT.t27 a_n8732_9422.t0 sky130_fd_pr__cap_mim_m3_1 l=18.34 w=7.84
X126 VDD.t16 VDD.t14 VDD.t15 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X127 VDD.t13 VDD.t10 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X128 GND.t51 GND.t49 VP.t0 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X129 a_n11778_11043.t4 a_n11634_10845.t15 a_n11634_10845.t16 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X130 VOUT.t3 CS_BIAS.t20 GND.t32 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X131 GND.t45 GND.t42 GND.t44 GND.t43 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=0 ps=0 w=7.13 l=2.31
X132 VOUT.t2 CS_BIAS.t21 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X133 a_n11634_10845.t18 a_n11634_10845.t17 a_n11778_11043.t3 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X134 VDD.t9 VDD.t7 VDD.t8 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X135 a_n11778_11043.t2 a_n11634_10845.t43 VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X136 a_n17232_8522.t10 VN.t8 a_n3337_n4072.t6 GND.t23 sky130_fd_pr__nfet_01v8 ad=5.1336 pd=15.7 as=5.1336 ps=15.7 w=7.13 l=2.31
X137 a_n8732_9422.t2 a_n11634_10845.t44 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X138 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=3.384 pd=10.84 as=3.384 ps=10.84 w=4.7 l=5.88
X139 VOUT.t18 a_n17232_8522.t19 VDD.t139 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X140 VOUT.t1 CS_BIAS.t22 GND.t12 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.9503 pd=6.57 as=4.2552 ps=13.26 w=5.91 l=4.37
X141 VDD.t6 VDD.t4 VDD.t5 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X142 VDD.t96 a_n11634_10845.t45 a_n11778_11043.t1 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X143 VDD.t3 VDD.t0 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=0 ps=0 w=2.43 l=5.92
X144 GND.t19 CS_BIAS.t23 VOUT.t0 GND.t18 sky130_fd_pr__nfet_01v8 ad=4.2552 pd=13.26 as=1.9503 ps=6.57 w=5.91 l=4.37
X145 a_n17232_8522.t0 a_n11634_10845.t46 a_n8732_9422.t9 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.8448 pd=3.22 as=0.8448 ps=3.22 w=2.56 l=5.82
X146 VOUT.t17 a_n17232_8522.t20 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X147 a_n8732_9422.t1 a_n11634_10845.t47 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=1.8432 pd=6.56 as=0.8448 ps=3.22 w=2.56 l=5.82
X148 VOUT.t16 a_n17232_8522.t21 VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.7496 pd=6.3 as=1.7496 ps=6.3 w=2.43 l=5.92
X149 GND.t41 GND.t39 VN.t0 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
R0 GND.n7594 GND.n7593 2254.37
R1 GND.n6503 GND.n1209 1000.86
R2 GND.n8010 GND.n149 857.672
R3 GND.n7876 GND.n289 857.672
R4 GND.n5440 GND.n2304 857.672
R5 GND.n5586 GND.n2316 857.672
R6 GND.n6272 GND.n1513 857.672
R7 GND.n4155 GND.n3288 857.672
R8 GND.n3777 GND.n3533 857.672
R9 GND.n3780 GND.n3524 857.672
R10 GND.n5642 GND.n2233 838.452
R11 GND.n5023 GND.n5022 838.452
R12 GND.n3114 GND.n3038 838.452
R13 GND.n4196 GND.n3036 838.452
R14 GND.n5250 GND.n144 833.646
R15 GND.n5292 GND.n290 833.646
R16 GND.n5041 GND.n2405 833.646
R17 GND.n5438 GND.n2433 833.646
R18 GND.n6380 GND.n1374 833.646
R19 GND.n1400 GND.n1372 833.646
R20 GND.n4153 GND.n1495 833.646
R21 GND.n6274 GND.n1464 833.646
R22 GND.n6626 GND.n1085 747.159
R23 GND.n7592 GND.n507 747.159
R24 GND.n7753 GND.n413 747.159
R25 GND.n6502 GND.n1210 747.159
R26 GND.n6625 GND.n1084 609.133
R27 GND.n6627 GND.n6626 585
R28 GND.n6626 GND.n6625 585
R29 GND.n1089 GND.n1088 585
R30 GND.n6624 GND.n1089 585
R31 GND.n6622 GND.n6621 585
R32 GND.n6623 GND.n6622 585
R33 GND.n6620 GND.n1091 585
R34 GND.n1091 GND.n1090 585
R35 GND.n6619 GND.n6618 585
R36 GND.n6618 GND.n6617 585
R37 GND.n1096 GND.n1095 585
R38 GND.n6616 GND.n1096 585
R39 GND.n6614 GND.n6613 585
R40 GND.n6615 GND.n6614 585
R41 GND.n6612 GND.n1098 585
R42 GND.n1098 GND.n1097 585
R43 GND.n6611 GND.n6610 585
R44 GND.n6610 GND.n6609 585
R45 GND.n1104 GND.n1103 585
R46 GND.n6608 GND.n1104 585
R47 GND.n6606 GND.n6605 585
R48 GND.n6607 GND.n6606 585
R49 GND.n6604 GND.n1106 585
R50 GND.n1106 GND.n1105 585
R51 GND.n6603 GND.n6602 585
R52 GND.n6602 GND.n6601 585
R53 GND.n1112 GND.n1111 585
R54 GND.n6600 GND.n1112 585
R55 GND.n6598 GND.n6597 585
R56 GND.n6599 GND.n6598 585
R57 GND.n6596 GND.n1114 585
R58 GND.n1114 GND.n1113 585
R59 GND.n6595 GND.n6594 585
R60 GND.n6594 GND.n6593 585
R61 GND.n1120 GND.n1119 585
R62 GND.n6592 GND.n1120 585
R63 GND.n6590 GND.n6589 585
R64 GND.n6591 GND.n6590 585
R65 GND.n6588 GND.n1122 585
R66 GND.n1122 GND.n1121 585
R67 GND.n6587 GND.n6586 585
R68 GND.n6586 GND.n6585 585
R69 GND.n1128 GND.n1127 585
R70 GND.n6584 GND.n1128 585
R71 GND.n6582 GND.n6581 585
R72 GND.n6583 GND.n6582 585
R73 GND.n6580 GND.n1130 585
R74 GND.n1130 GND.n1129 585
R75 GND.n6579 GND.n6578 585
R76 GND.n6578 GND.n6577 585
R77 GND.n1136 GND.n1135 585
R78 GND.n6576 GND.n1136 585
R79 GND.n6574 GND.n6573 585
R80 GND.n6575 GND.n6574 585
R81 GND.n6572 GND.n1138 585
R82 GND.n1138 GND.n1137 585
R83 GND.n6571 GND.n6570 585
R84 GND.n6570 GND.n6569 585
R85 GND.n1144 GND.n1143 585
R86 GND.n6568 GND.n1144 585
R87 GND.n6566 GND.n6565 585
R88 GND.n6567 GND.n6566 585
R89 GND.n6564 GND.n1146 585
R90 GND.n1146 GND.n1145 585
R91 GND.n6563 GND.n6562 585
R92 GND.n6562 GND.n6561 585
R93 GND.n1152 GND.n1151 585
R94 GND.n6560 GND.n1152 585
R95 GND.n6558 GND.n6557 585
R96 GND.n6559 GND.n6558 585
R97 GND.n6556 GND.n1154 585
R98 GND.n1154 GND.n1153 585
R99 GND.n6555 GND.n6554 585
R100 GND.n6554 GND.n6553 585
R101 GND.n1160 GND.n1159 585
R102 GND.n6552 GND.n1160 585
R103 GND.n6550 GND.n6549 585
R104 GND.n6551 GND.n6550 585
R105 GND.n6548 GND.n1162 585
R106 GND.n1162 GND.n1161 585
R107 GND.n6547 GND.n6546 585
R108 GND.n6546 GND.n6545 585
R109 GND.n1168 GND.n1167 585
R110 GND.n6544 GND.n1168 585
R111 GND.n6542 GND.n6541 585
R112 GND.n6543 GND.n6542 585
R113 GND.n6540 GND.n1170 585
R114 GND.n1170 GND.n1169 585
R115 GND.n6539 GND.n6538 585
R116 GND.n6538 GND.n6537 585
R117 GND.n1176 GND.n1175 585
R118 GND.n6536 GND.n1176 585
R119 GND.n6534 GND.n6533 585
R120 GND.n6535 GND.n6534 585
R121 GND.n6532 GND.n1178 585
R122 GND.n1178 GND.n1177 585
R123 GND.n6531 GND.n6530 585
R124 GND.n6530 GND.n6529 585
R125 GND.n1184 GND.n1183 585
R126 GND.n6528 GND.n1184 585
R127 GND.n6526 GND.n6525 585
R128 GND.n6527 GND.n6526 585
R129 GND.n6524 GND.n1186 585
R130 GND.n1186 GND.n1185 585
R131 GND.n6523 GND.n6522 585
R132 GND.n6522 GND.n6521 585
R133 GND.n1192 GND.n1191 585
R134 GND.n6520 GND.n1192 585
R135 GND.n6518 GND.n6517 585
R136 GND.n6519 GND.n6518 585
R137 GND.n6516 GND.n1194 585
R138 GND.n1194 GND.n1193 585
R139 GND.n6515 GND.n6514 585
R140 GND.n6514 GND.n6513 585
R141 GND.n1200 GND.n1199 585
R142 GND.n6512 GND.n1200 585
R143 GND.n6510 GND.n6509 585
R144 GND.n6511 GND.n6510 585
R145 GND.n6508 GND.n1202 585
R146 GND.n1202 GND.n1201 585
R147 GND.n6507 GND.n6506 585
R148 GND.n6506 GND.n6505 585
R149 GND.n1208 GND.n1207 585
R150 GND.n6504 GND.n1208 585
R151 GND.n6502 GND.n6501 585
R152 GND.n6503 GND.n6502 585
R153 GND.n1086 GND.n1085 585
R154 GND.n1085 GND.n1084 585
R155 GND.n6632 GND.n6631 585
R156 GND.n6633 GND.n6632 585
R157 GND.n1083 GND.n1082 585
R158 GND.n6634 GND.n1083 585
R159 GND.n6637 GND.n6636 585
R160 GND.n6636 GND.n6635 585
R161 GND.n1080 GND.n1079 585
R162 GND.n1079 GND.n1078 585
R163 GND.n6642 GND.n6641 585
R164 GND.n6643 GND.n6642 585
R165 GND.n1077 GND.n1076 585
R166 GND.n6644 GND.n1077 585
R167 GND.n6647 GND.n6646 585
R168 GND.n6646 GND.n6645 585
R169 GND.n1074 GND.n1073 585
R170 GND.n1073 GND.n1072 585
R171 GND.n6652 GND.n6651 585
R172 GND.n6653 GND.n6652 585
R173 GND.n1071 GND.n1070 585
R174 GND.n6654 GND.n1071 585
R175 GND.n6657 GND.n6656 585
R176 GND.n6656 GND.n6655 585
R177 GND.n1068 GND.n1067 585
R178 GND.n1067 GND.n1066 585
R179 GND.n6662 GND.n6661 585
R180 GND.n6663 GND.n6662 585
R181 GND.n1065 GND.n1064 585
R182 GND.n6664 GND.n1065 585
R183 GND.n6667 GND.n6666 585
R184 GND.n6666 GND.n6665 585
R185 GND.n1062 GND.n1061 585
R186 GND.n1061 GND.n1060 585
R187 GND.n6672 GND.n6671 585
R188 GND.n6673 GND.n6672 585
R189 GND.n1059 GND.n1058 585
R190 GND.n6674 GND.n1059 585
R191 GND.n6677 GND.n6676 585
R192 GND.n6676 GND.n6675 585
R193 GND.n1056 GND.n1055 585
R194 GND.n1055 GND.n1054 585
R195 GND.n6682 GND.n6681 585
R196 GND.n6683 GND.n6682 585
R197 GND.n1053 GND.n1052 585
R198 GND.n6684 GND.n1053 585
R199 GND.n6687 GND.n6686 585
R200 GND.n6686 GND.n6685 585
R201 GND.n1050 GND.n1049 585
R202 GND.n1049 GND.n1048 585
R203 GND.n6692 GND.n6691 585
R204 GND.n6693 GND.n6692 585
R205 GND.n1047 GND.n1046 585
R206 GND.n6694 GND.n1047 585
R207 GND.n6697 GND.n6696 585
R208 GND.n6696 GND.n6695 585
R209 GND.n1044 GND.n1043 585
R210 GND.n1043 GND.n1042 585
R211 GND.n6702 GND.n6701 585
R212 GND.n6703 GND.n6702 585
R213 GND.n1041 GND.n1040 585
R214 GND.n6704 GND.n1041 585
R215 GND.n6707 GND.n6706 585
R216 GND.n6706 GND.n6705 585
R217 GND.n1038 GND.n1037 585
R218 GND.n1037 GND.n1036 585
R219 GND.n6712 GND.n6711 585
R220 GND.n6713 GND.n6712 585
R221 GND.n1035 GND.n1034 585
R222 GND.n6714 GND.n1035 585
R223 GND.n6717 GND.n6716 585
R224 GND.n6716 GND.n6715 585
R225 GND.n1032 GND.n1031 585
R226 GND.n1031 GND.n1030 585
R227 GND.n6722 GND.n6721 585
R228 GND.n6723 GND.n6722 585
R229 GND.n1029 GND.n1028 585
R230 GND.n6724 GND.n1029 585
R231 GND.n6727 GND.n6726 585
R232 GND.n6726 GND.n6725 585
R233 GND.n1026 GND.n1025 585
R234 GND.n1025 GND.n1024 585
R235 GND.n6732 GND.n6731 585
R236 GND.n6733 GND.n6732 585
R237 GND.n1023 GND.n1022 585
R238 GND.n6734 GND.n1023 585
R239 GND.n6737 GND.n6736 585
R240 GND.n6736 GND.n6735 585
R241 GND.n1020 GND.n1019 585
R242 GND.n1019 GND.n1018 585
R243 GND.n6742 GND.n6741 585
R244 GND.n6743 GND.n6742 585
R245 GND.n1017 GND.n1016 585
R246 GND.n6744 GND.n1017 585
R247 GND.n6747 GND.n6746 585
R248 GND.n6746 GND.n6745 585
R249 GND.n1014 GND.n1013 585
R250 GND.n1013 GND.n1012 585
R251 GND.n6752 GND.n6751 585
R252 GND.n6753 GND.n6752 585
R253 GND.n1011 GND.n1010 585
R254 GND.n6754 GND.n1011 585
R255 GND.n6757 GND.n6756 585
R256 GND.n6756 GND.n6755 585
R257 GND.n1008 GND.n1007 585
R258 GND.n1007 GND.n1006 585
R259 GND.n6762 GND.n6761 585
R260 GND.n6763 GND.n6762 585
R261 GND.n1005 GND.n1004 585
R262 GND.n6764 GND.n1005 585
R263 GND.n6767 GND.n6766 585
R264 GND.n6766 GND.n6765 585
R265 GND.n1002 GND.n1001 585
R266 GND.n1001 GND.n1000 585
R267 GND.n6772 GND.n6771 585
R268 GND.n6773 GND.n6772 585
R269 GND.n999 GND.n998 585
R270 GND.n6774 GND.n999 585
R271 GND.n6777 GND.n6776 585
R272 GND.n6776 GND.n6775 585
R273 GND.n996 GND.n995 585
R274 GND.n995 GND.n994 585
R275 GND.n6782 GND.n6781 585
R276 GND.n6783 GND.n6782 585
R277 GND.n993 GND.n992 585
R278 GND.n6784 GND.n993 585
R279 GND.n6787 GND.n6786 585
R280 GND.n6786 GND.n6785 585
R281 GND.n990 GND.n989 585
R282 GND.n989 GND.n988 585
R283 GND.n6792 GND.n6791 585
R284 GND.n6793 GND.n6792 585
R285 GND.n987 GND.n986 585
R286 GND.n6794 GND.n987 585
R287 GND.n6797 GND.n6796 585
R288 GND.n6796 GND.n6795 585
R289 GND.n984 GND.n983 585
R290 GND.n983 GND.n982 585
R291 GND.n6802 GND.n6801 585
R292 GND.n6803 GND.n6802 585
R293 GND.n981 GND.n980 585
R294 GND.n6804 GND.n981 585
R295 GND.n6807 GND.n6806 585
R296 GND.n6806 GND.n6805 585
R297 GND.n978 GND.n977 585
R298 GND.n977 GND.n976 585
R299 GND.n6812 GND.n6811 585
R300 GND.n6813 GND.n6812 585
R301 GND.n975 GND.n974 585
R302 GND.n6814 GND.n975 585
R303 GND.n6817 GND.n6816 585
R304 GND.n6816 GND.n6815 585
R305 GND.n972 GND.n971 585
R306 GND.n971 GND.n970 585
R307 GND.n6822 GND.n6821 585
R308 GND.n6823 GND.n6822 585
R309 GND.n969 GND.n968 585
R310 GND.n6824 GND.n969 585
R311 GND.n6827 GND.n6826 585
R312 GND.n6826 GND.n6825 585
R313 GND.n966 GND.n965 585
R314 GND.n965 GND.n964 585
R315 GND.n6832 GND.n6831 585
R316 GND.n6833 GND.n6832 585
R317 GND.n963 GND.n962 585
R318 GND.n6834 GND.n963 585
R319 GND.n6837 GND.n6836 585
R320 GND.n6836 GND.n6835 585
R321 GND.n960 GND.n959 585
R322 GND.n959 GND.n958 585
R323 GND.n6842 GND.n6841 585
R324 GND.n6843 GND.n6842 585
R325 GND.n957 GND.n956 585
R326 GND.n6844 GND.n957 585
R327 GND.n6847 GND.n6846 585
R328 GND.n6846 GND.n6845 585
R329 GND.n954 GND.n953 585
R330 GND.n953 GND.n952 585
R331 GND.n6852 GND.n6851 585
R332 GND.n6853 GND.n6852 585
R333 GND.n951 GND.n950 585
R334 GND.n6854 GND.n951 585
R335 GND.n6857 GND.n6856 585
R336 GND.n6856 GND.n6855 585
R337 GND.n948 GND.n947 585
R338 GND.n947 GND.n946 585
R339 GND.n6862 GND.n6861 585
R340 GND.n6863 GND.n6862 585
R341 GND.n945 GND.n944 585
R342 GND.n6864 GND.n945 585
R343 GND.n6867 GND.n6866 585
R344 GND.n6866 GND.n6865 585
R345 GND.n942 GND.n941 585
R346 GND.n941 GND.n940 585
R347 GND.n6872 GND.n6871 585
R348 GND.n6873 GND.n6872 585
R349 GND.n939 GND.n938 585
R350 GND.n6874 GND.n939 585
R351 GND.n6877 GND.n6876 585
R352 GND.n6876 GND.n6875 585
R353 GND.n936 GND.n935 585
R354 GND.n935 GND.n934 585
R355 GND.n6882 GND.n6881 585
R356 GND.n6883 GND.n6882 585
R357 GND.n933 GND.n932 585
R358 GND.n6884 GND.n933 585
R359 GND.n6887 GND.n6886 585
R360 GND.n6886 GND.n6885 585
R361 GND.n930 GND.n929 585
R362 GND.n929 GND.n928 585
R363 GND.n6892 GND.n6891 585
R364 GND.n6893 GND.n6892 585
R365 GND.n927 GND.n926 585
R366 GND.n6894 GND.n927 585
R367 GND.n6897 GND.n6896 585
R368 GND.n6896 GND.n6895 585
R369 GND.n924 GND.n923 585
R370 GND.n923 GND.n922 585
R371 GND.n6902 GND.n6901 585
R372 GND.n6903 GND.n6902 585
R373 GND.n921 GND.n920 585
R374 GND.n6904 GND.n921 585
R375 GND.n6907 GND.n6906 585
R376 GND.n6906 GND.n6905 585
R377 GND.n918 GND.n917 585
R378 GND.n917 GND.n916 585
R379 GND.n6912 GND.n6911 585
R380 GND.n6913 GND.n6912 585
R381 GND.n915 GND.n914 585
R382 GND.n6914 GND.n915 585
R383 GND.n6917 GND.n6916 585
R384 GND.n6916 GND.n6915 585
R385 GND.n912 GND.n911 585
R386 GND.n911 GND.n910 585
R387 GND.n6922 GND.n6921 585
R388 GND.n6923 GND.n6922 585
R389 GND.n909 GND.n908 585
R390 GND.n6924 GND.n909 585
R391 GND.n6927 GND.n6926 585
R392 GND.n6926 GND.n6925 585
R393 GND.n906 GND.n905 585
R394 GND.n905 GND.n904 585
R395 GND.n6932 GND.n6931 585
R396 GND.n6933 GND.n6932 585
R397 GND.n903 GND.n902 585
R398 GND.n6934 GND.n903 585
R399 GND.n6937 GND.n6936 585
R400 GND.n6936 GND.n6935 585
R401 GND.n900 GND.n899 585
R402 GND.n899 GND.n898 585
R403 GND.n6942 GND.n6941 585
R404 GND.n6943 GND.n6942 585
R405 GND.n897 GND.n896 585
R406 GND.n6944 GND.n897 585
R407 GND.n6947 GND.n6946 585
R408 GND.n6946 GND.n6945 585
R409 GND.n894 GND.n893 585
R410 GND.n893 GND.n892 585
R411 GND.n6952 GND.n6951 585
R412 GND.n6953 GND.n6952 585
R413 GND.n891 GND.n890 585
R414 GND.n6954 GND.n891 585
R415 GND.n6957 GND.n6956 585
R416 GND.n6956 GND.n6955 585
R417 GND.n888 GND.n887 585
R418 GND.n887 GND.n886 585
R419 GND.n6962 GND.n6961 585
R420 GND.n6963 GND.n6962 585
R421 GND.n885 GND.n884 585
R422 GND.n6964 GND.n885 585
R423 GND.n6967 GND.n6966 585
R424 GND.n6966 GND.n6965 585
R425 GND.n882 GND.n881 585
R426 GND.n881 GND.n880 585
R427 GND.n6972 GND.n6971 585
R428 GND.n6973 GND.n6972 585
R429 GND.n879 GND.n878 585
R430 GND.n6974 GND.n879 585
R431 GND.n6977 GND.n6976 585
R432 GND.n6976 GND.n6975 585
R433 GND.n876 GND.n875 585
R434 GND.n875 GND.n874 585
R435 GND.n6982 GND.n6981 585
R436 GND.n6983 GND.n6982 585
R437 GND.n873 GND.n872 585
R438 GND.n6984 GND.n873 585
R439 GND.n6987 GND.n6986 585
R440 GND.n6986 GND.n6985 585
R441 GND.n870 GND.n869 585
R442 GND.n869 GND.n868 585
R443 GND.n6992 GND.n6991 585
R444 GND.n6993 GND.n6992 585
R445 GND.n867 GND.n866 585
R446 GND.n6994 GND.n867 585
R447 GND.n6997 GND.n6996 585
R448 GND.n6996 GND.n6995 585
R449 GND.n864 GND.n863 585
R450 GND.n863 GND.n862 585
R451 GND.n7002 GND.n7001 585
R452 GND.n7003 GND.n7002 585
R453 GND.n861 GND.n860 585
R454 GND.n7004 GND.n861 585
R455 GND.n7007 GND.n7006 585
R456 GND.n7006 GND.n7005 585
R457 GND.n858 GND.n857 585
R458 GND.n857 GND.n856 585
R459 GND.n7012 GND.n7011 585
R460 GND.n7013 GND.n7012 585
R461 GND.n855 GND.n854 585
R462 GND.n7014 GND.n855 585
R463 GND.n7017 GND.n7016 585
R464 GND.n7016 GND.n7015 585
R465 GND.n852 GND.n851 585
R466 GND.n851 GND.n850 585
R467 GND.n7022 GND.n7021 585
R468 GND.n7023 GND.n7022 585
R469 GND.n849 GND.n848 585
R470 GND.n7024 GND.n849 585
R471 GND.n7027 GND.n7026 585
R472 GND.n7026 GND.n7025 585
R473 GND.n846 GND.n845 585
R474 GND.n845 GND.n844 585
R475 GND.n7032 GND.n7031 585
R476 GND.n7033 GND.n7032 585
R477 GND.n843 GND.n842 585
R478 GND.n7034 GND.n843 585
R479 GND.n7037 GND.n7036 585
R480 GND.n7036 GND.n7035 585
R481 GND.n840 GND.n839 585
R482 GND.n839 GND.n838 585
R483 GND.n7042 GND.n7041 585
R484 GND.n7043 GND.n7042 585
R485 GND.n837 GND.n836 585
R486 GND.n7044 GND.n837 585
R487 GND.n7047 GND.n7046 585
R488 GND.n7046 GND.n7045 585
R489 GND.n834 GND.n833 585
R490 GND.n833 GND.n832 585
R491 GND.n7052 GND.n7051 585
R492 GND.n7053 GND.n7052 585
R493 GND.n831 GND.n830 585
R494 GND.n7054 GND.n831 585
R495 GND.n7057 GND.n7056 585
R496 GND.n7056 GND.n7055 585
R497 GND.n828 GND.n827 585
R498 GND.n827 GND.n826 585
R499 GND.n7062 GND.n7061 585
R500 GND.n7063 GND.n7062 585
R501 GND.n825 GND.n824 585
R502 GND.n7064 GND.n825 585
R503 GND.n7067 GND.n7066 585
R504 GND.n7066 GND.n7065 585
R505 GND.n822 GND.n821 585
R506 GND.n821 GND.n820 585
R507 GND.n7072 GND.n7071 585
R508 GND.n7073 GND.n7072 585
R509 GND.n819 GND.n818 585
R510 GND.n7074 GND.n819 585
R511 GND.n7077 GND.n7076 585
R512 GND.n7076 GND.n7075 585
R513 GND.n816 GND.n815 585
R514 GND.n815 GND.n814 585
R515 GND.n7082 GND.n7081 585
R516 GND.n7083 GND.n7082 585
R517 GND.n813 GND.n812 585
R518 GND.n7084 GND.n813 585
R519 GND.n7087 GND.n7086 585
R520 GND.n7086 GND.n7085 585
R521 GND.n810 GND.n809 585
R522 GND.n809 GND.n808 585
R523 GND.n7092 GND.n7091 585
R524 GND.n7093 GND.n7092 585
R525 GND.n807 GND.n806 585
R526 GND.n7094 GND.n807 585
R527 GND.n7097 GND.n7096 585
R528 GND.n7096 GND.n7095 585
R529 GND.n804 GND.n803 585
R530 GND.n803 GND.n802 585
R531 GND.n7102 GND.n7101 585
R532 GND.n7103 GND.n7102 585
R533 GND.n801 GND.n800 585
R534 GND.n7104 GND.n801 585
R535 GND.n7107 GND.n7106 585
R536 GND.n7106 GND.n7105 585
R537 GND.n798 GND.n797 585
R538 GND.n797 GND.n796 585
R539 GND.n7112 GND.n7111 585
R540 GND.n7113 GND.n7112 585
R541 GND.n795 GND.n794 585
R542 GND.n7114 GND.n795 585
R543 GND.n7117 GND.n7116 585
R544 GND.n7116 GND.n7115 585
R545 GND.n792 GND.n791 585
R546 GND.n791 GND.n790 585
R547 GND.n7122 GND.n7121 585
R548 GND.n7123 GND.n7122 585
R549 GND.n789 GND.n788 585
R550 GND.n7124 GND.n789 585
R551 GND.n7127 GND.n7126 585
R552 GND.n7126 GND.n7125 585
R553 GND.n786 GND.n785 585
R554 GND.n785 GND.n784 585
R555 GND.n7132 GND.n7131 585
R556 GND.n7133 GND.n7132 585
R557 GND.n783 GND.n782 585
R558 GND.n7134 GND.n783 585
R559 GND.n7137 GND.n7136 585
R560 GND.n7136 GND.n7135 585
R561 GND.n780 GND.n779 585
R562 GND.n779 GND.n778 585
R563 GND.n7142 GND.n7141 585
R564 GND.n7143 GND.n7142 585
R565 GND.n777 GND.n776 585
R566 GND.n7144 GND.n777 585
R567 GND.n7147 GND.n7146 585
R568 GND.n7146 GND.n7145 585
R569 GND.n774 GND.n773 585
R570 GND.n773 GND.n772 585
R571 GND.n7152 GND.n7151 585
R572 GND.n7153 GND.n7152 585
R573 GND.n771 GND.n770 585
R574 GND.n7154 GND.n771 585
R575 GND.n7157 GND.n7156 585
R576 GND.n7156 GND.n7155 585
R577 GND.n768 GND.n767 585
R578 GND.n767 GND.n766 585
R579 GND.n7162 GND.n7161 585
R580 GND.n7163 GND.n7162 585
R581 GND.n765 GND.n764 585
R582 GND.n7164 GND.n765 585
R583 GND.n7167 GND.n7166 585
R584 GND.n7166 GND.n7165 585
R585 GND.n762 GND.n761 585
R586 GND.n761 GND.n760 585
R587 GND.n7172 GND.n7171 585
R588 GND.n7173 GND.n7172 585
R589 GND.n759 GND.n758 585
R590 GND.n7174 GND.n759 585
R591 GND.n7177 GND.n7176 585
R592 GND.n7176 GND.n7175 585
R593 GND.n756 GND.n755 585
R594 GND.n755 GND.n754 585
R595 GND.n7182 GND.n7181 585
R596 GND.n7183 GND.n7182 585
R597 GND.n753 GND.n752 585
R598 GND.n7184 GND.n753 585
R599 GND.n7187 GND.n7186 585
R600 GND.n7186 GND.n7185 585
R601 GND.n750 GND.n749 585
R602 GND.n749 GND.n748 585
R603 GND.n7192 GND.n7191 585
R604 GND.n7193 GND.n7192 585
R605 GND.n747 GND.n746 585
R606 GND.n7194 GND.n747 585
R607 GND.n7197 GND.n7196 585
R608 GND.n7196 GND.n7195 585
R609 GND.n744 GND.n743 585
R610 GND.n743 GND.n742 585
R611 GND.n7202 GND.n7201 585
R612 GND.n7203 GND.n7202 585
R613 GND.n741 GND.n740 585
R614 GND.n7204 GND.n741 585
R615 GND.n7207 GND.n7206 585
R616 GND.n7206 GND.n7205 585
R617 GND.n738 GND.n737 585
R618 GND.n737 GND.n736 585
R619 GND.n7212 GND.n7211 585
R620 GND.n7213 GND.n7212 585
R621 GND.n735 GND.n734 585
R622 GND.n7214 GND.n735 585
R623 GND.n7217 GND.n7216 585
R624 GND.n7216 GND.n7215 585
R625 GND.n732 GND.n731 585
R626 GND.n731 GND.n730 585
R627 GND.n7222 GND.n7221 585
R628 GND.n7223 GND.n7222 585
R629 GND.n729 GND.n728 585
R630 GND.n7224 GND.n729 585
R631 GND.n7227 GND.n7226 585
R632 GND.n7226 GND.n7225 585
R633 GND.n726 GND.n725 585
R634 GND.n725 GND.n724 585
R635 GND.n7232 GND.n7231 585
R636 GND.n7233 GND.n7232 585
R637 GND.n723 GND.n722 585
R638 GND.n7234 GND.n723 585
R639 GND.n7237 GND.n7236 585
R640 GND.n7236 GND.n7235 585
R641 GND.n720 GND.n719 585
R642 GND.n719 GND.n718 585
R643 GND.n7242 GND.n7241 585
R644 GND.n7243 GND.n7242 585
R645 GND.n717 GND.n716 585
R646 GND.n7244 GND.n717 585
R647 GND.n7247 GND.n7246 585
R648 GND.n7246 GND.n7245 585
R649 GND.n714 GND.n713 585
R650 GND.n713 GND.n712 585
R651 GND.n7252 GND.n7251 585
R652 GND.n7253 GND.n7252 585
R653 GND.n711 GND.n710 585
R654 GND.n7254 GND.n711 585
R655 GND.n7257 GND.n7256 585
R656 GND.n7256 GND.n7255 585
R657 GND.n708 GND.n707 585
R658 GND.n707 GND.n706 585
R659 GND.n7262 GND.n7261 585
R660 GND.n7263 GND.n7262 585
R661 GND.n705 GND.n704 585
R662 GND.n7264 GND.n705 585
R663 GND.n7267 GND.n7266 585
R664 GND.n7266 GND.n7265 585
R665 GND.n702 GND.n701 585
R666 GND.n701 GND.n700 585
R667 GND.n7272 GND.n7271 585
R668 GND.n7273 GND.n7272 585
R669 GND.n699 GND.n698 585
R670 GND.n7274 GND.n699 585
R671 GND.n7277 GND.n7276 585
R672 GND.n7276 GND.n7275 585
R673 GND.n696 GND.n695 585
R674 GND.n695 GND.n694 585
R675 GND.n7282 GND.n7281 585
R676 GND.n7283 GND.n7282 585
R677 GND.n693 GND.n692 585
R678 GND.n7284 GND.n693 585
R679 GND.n7287 GND.n7286 585
R680 GND.n7286 GND.n7285 585
R681 GND.n690 GND.n689 585
R682 GND.n689 GND.n688 585
R683 GND.n7292 GND.n7291 585
R684 GND.n7293 GND.n7292 585
R685 GND.n687 GND.n686 585
R686 GND.n7294 GND.n687 585
R687 GND.n7297 GND.n7296 585
R688 GND.n7296 GND.n7295 585
R689 GND.n684 GND.n683 585
R690 GND.n683 GND.n682 585
R691 GND.n7302 GND.n7301 585
R692 GND.n7303 GND.n7302 585
R693 GND.n681 GND.n680 585
R694 GND.n7304 GND.n681 585
R695 GND.n7307 GND.n7306 585
R696 GND.n7306 GND.n7305 585
R697 GND.n678 GND.n677 585
R698 GND.n677 GND.n676 585
R699 GND.n7312 GND.n7311 585
R700 GND.n7313 GND.n7312 585
R701 GND.n675 GND.n674 585
R702 GND.n7314 GND.n675 585
R703 GND.n7317 GND.n7316 585
R704 GND.n7316 GND.n7315 585
R705 GND.n672 GND.n671 585
R706 GND.n671 GND.n670 585
R707 GND.n7322 GND.n7321 585
R708 GND.n7323 GND.n7322 585
R709 GND.n669 GND.n668 585
R710 GND.n7324 GND.n669 585
R711 GND.n7327 GND.n7326 585
R712 GND.n7326 GND.n7325 585
R713 GND.n666 GND.n665 585
R714 GND.n665 GND.n664 585
R715 GND.n7332 GND.n7331 585
R716 GND.n7333 GND.n7332 585
R717 GND.n663 GND.n662 585
R718 GND.n7334 GND.n663 585
R719 GND.n7337 GND.n7336 585
R720 GND.n7336 GND.n7335 585
R721 GND.n660 GND.n659 585
R722 GND.n659 GND.n658 585
R723 GND.n7342 GND.n7341 585
R724 GND.n7343 GND.n7342 585
R725 GND.n657 GND.n656 585
R726 GND.n7344 GND.n657 585
R727 GND.n7347 GND.n7346 585
R728 GND.n7346 GND.n7345 585
R729 GND.n654 GND.n653 585
R730 GND.n653 GND.n652 585
R731 GND.n7352 GND.n7351 585
R732 GND.n7353 GND.n7352 585
R733 GND.n651 GND.n650 585
R734 GND.n7354 GND.n651 585
R735 GND.n7357 GND.n7356 585
R736 GND.n7356 GND.n7355 585
R737 GND.n648 GND.n647 585
R738 GND.n647 GND.n646 585
R739 GND.n7362 GND.n7361 585
R740 GND.n7363 GND.n7362 585
R741 GND.n645 GND.n644 585
R742 GND.n7364 GND.n645 585
R743 GND.n7367 GND.n7366 585
R744 GND.n7366 GND.n7365 585
R745 GND.n642 GND.n641 585
R746 GND.n641 GND.n640 585
R747 GND.n7372 GND.n7371 585
R748 GND.n7373 GND.n7372 585
R749 GND.n639 GND.n638 585
R750 GND.n7374 GND.n639 585
R751 GND.n7377 GND.n7376 585
R752 GND.n7376 GND.n7375 585
R753 GND.n636 GND.n635 585
R754 GND.n635 GND.n634 585
R755 GND.n7382 GND.n7381 585
R756 GND.n7383 GND.n7382 585
R757 GND.n633 GND.n632 585
R758 GND.n7384 GND.n633 585
R759 GND.n7387 GND.n7386 585
R760 GND.n7386 GND.n7385 585
R761 GND.n630 GND.n629 585
R762 GND.n629 GND.n628 585
R763 GND.n7392 GND.n7391 585
R764 GND.n7393 GND.n7392 585
R765 GND.n627 GND.n626 585
R766 GND.n7394 GND.n627 585
R767 GND.n7397 GND.n7396 585
R768 GND.n7396 GND.n7395 585
R769 GND.n624 GND.n623 585
R770 GND.n623 GND.n622 585
R771 GND.n7402 GND.n7401 585
R772 GND.n7403 GND.n7402 585
R773 GND.n621 GND.n620 585
R774 GND.n7404 GND.n621 585
R775 GND.n7407 GND.n7406 585
R776 GND.n7406 GND.n7405 585
R777 GND.n618 GND.n617 585
R778 GND.n617 GND.n616 585
R779 GND.n7412 GND.n7411 585
R780 GND.n7413 GND.n7412 585
R781 GND.n615 GND.n614 585
R782 GND.n7414 GND.n615 585
R783 GND.n7417 GND.n7416 585
R784 GND.n7416 GND.n7415 585
R785 GND.n612 GND.n611 585
R786 GND.n611 GND.n610 585
R787 GND.n7422 GND.n7421 585
R788 GND.n7423 GND.n7422 585
R789 GND.n609 GND.n608 585
R790 GND.n7424 GND.n609 585
R791 GND.n7427 GND.n7426 585
R792 GND.n7426 GND.n7425 585
R793 GND.n606 GND.n605 585
R794 GND.n605 GND.n604 585
R795 GND.n7432 GND.n7431 585
R796 GND.n7433 GND.n7432 585
R797 GND.n603 GND.n602 585
R798 GND.n7434 GND.n603 585
R799 GND.n7437 GND.n7436 585
R800 GND.n7436 GND.n7435 585
R801 GND.n600 GND.n599 585
R802 GND.n599 GND.n598 585
R803 GND.n7442 GND.n7441 585
R804 GND.n7443 GND.n7442 585
R805 GND.n597 GND.n596 585
R806 GND.n7444 GND.n597 585
R807 GND.n7447 GND.n7446 585
R808 GND.n7446 GND.n7445 585
R809 GND.n594 GND.n593 585
R810 GND.n593 GND.n592 585
R811 GND.n7452 GND.n7451 585
R812 GND.n7453 GND.n7452 585
R813 GND.n591 GND.n590 585
R814 GND.n7454 GND.n591 585
R815 GND.n7457 GND.n7456 585
R816 GND.n7456 GND.n7455 585
R817 GND.n588 GND.n587 585
R818 GND.n587 GND.n586 585
R819 GND.n7462 GND.n7461 585
R820 GND.n7463 GND.n7462 585
R821 GND.n585 GND.n584 585
R822 GND.n7464 GND.n585 585
R823 GND.n7467 GND.n7466 585
R824 GND.n7466 GND.n7465 585
R825 GND.n582 GND.n581 585
R826 GND.n581 GND.n580 585
R827 GND.n7472 GND.n7471 585
R828 GND.n7473 GND.n7472 585
R829 GND.n579 GND.n578 585
R830 GND.n7474 GND.n579 585
R831 GND.n7477 GND.n7476 585
R832 GND.n7476 GND.n7475 585
R833 GND.n576 GND.n575 585
R834 GND.n575 GND.n574 585
R835 GND.n7482 GND.n7481 585
R836 GND.n7483 GND.n7482 585
R837 GND.n573 GND.n572 585
R838 GND.n7484 GND.n573 585
R839 GND.n7487 GND.n7486 585
R840 GND.n7486 GND.n7485 585
R841 GND.n570 GND.n569 585
R842 GND.n569 GND.n568 585
R843 GND.n7492 GND.n7491 585
R844 GND.n7493 GND.n7492 585
R845 GND.n567 GND.n566 585
R846 GND.n7494 GND.n567 585
R847 GND.n7497 GND.n7496 585
R848 GND.n7496 GND.n7495 585
R849 GND.n564 GND.n563 585
R850 GND.n563 GND.n562 585
R851 GND.n7502 GND.n7501 585
R852 GND.n7503 GND.n7502 585
R853 GND.n561 GND.n560 585
R854 GND.n7504 GND.n561 585
R855 GND.n7507 GND.n7506 585
R856 GND.n7506 GND.n7505 585
R857 GND.n558 GND.n557 585
R858 GND.n557 GND.n556 585
R859 GND.n7512 GND.n7511 585
R860 GND.n7513 GND.n7512 585
R861 GND.n555 GND.n554 585
R862 GND.n7514 GND.n555 585
R863 GND.n7517 GND.n7516 585
R864 GND.n7516 GND.n7515 585
R865 GND.n552 GND.n551 585
R866 GND.n551 GND.n550 585
R867 GND.n7522 GND.n7521 585
R868 GND.n7523 GND.n7522 585
R869 GND.n549 GND.n548 585
R870 GND.n7524 GND.n549 585
R871 GND.n7527 GND.n7526 585
R872 GND.n7526 GND.n7525 585
R873 GND.n546 GND.n545 585
R874 GND.n545 GND.n544 585
R875 GND.n7532 GND.n7531 585
R876 GND.n7533 GND.n7532 585
R877 GND.n543 GND.n542 585
R878 GND.n7534 GND.n543 585
R879 GND.n7537 GND.n7536 585
R880 GND.n7536 GND.n7535 585
R881 GND.n540 GND.n539 585
R882 GND.n539 GND.n538 585
R883 GND.n7542 GND.n7541 585
R884 GND.n7543 GND.n7542 585
R885 GND.n537 GND.n536 585
R886 GND.n7544 GND.n537 585
R887 GND.n7547 GND.n7546 585
R888 GND.n7546 GND.n7545 585
R889 GND.n534 GND.n533 585
R890 GND.n533 GND.n532 585
R891 GND.n7552 GND.n7551 585
R892 GND.n7553 GND.n7552 585
R893 GND.n531 GND.n530 585
R894 GND.n7554 GND.n531 585
R895 GND.n7557 GND.n7556 585
R896 GND.n7556 GND.n7555 585
R897 GND.n528 GND.n527 585
R898 GND.n527 GND.n526 585
R899 GND.n7562 GND.n7561 585
R900 GND.n7563 GND.n7562 585
R901 GND.n525 GND.n524 585
R902 GND.n7564 GND.n525 585
R903 GND.n7567 GND.n7566 585
R904 GND.n7566 GND.n7565 585
R905 GND.n522 GND.n521 585
R906 GND.n521 GND.n520 585
R907 GND.n7572 GND.n7571 585
R908 GND.n7573 GND.n7572 585
R909 GND.n519 GND.n518 585
R910 GND.n7574 GND.n519 585
R911 GND.n7577 GND.n7576 585
R912 GND.n7576 GND.n7575 585
R913 GND.n516 GND.n515 585
R914 GND.n515 GND.n514 585
R915 GND.n7582 GND.n7581 585
R916 GND.n7583 GND.n7582 585
R917 GND.n513 GND.n512 585
R918 GND.n7584 GND.n513 585
R919 GND.n7587 GND.n7586 585
R920 GND.n7586 GND.n7585 585
R921 GND.n510 GND.n509 585
R922 GND.n509 GND.n508 585
R923 GND.n7592 GND.n7591 585
R924 GND.n7593 GND.n7592 585
R925 GND.n7749 GND.n413 585
R926 GND.n413 GND.n412 585
R927 GND.n7748 GND.n7747 585
R928 GND.n7747 GND.n7746 585
R929 GND.n417 GND.n416 585
R930 GND.n7745 GND.n417 585
R931 GND.n7743 GND.n7742 585
R932 GND.n7744 GND.n7743 585
R933 GND.n420 GND.n419 585
R934 GND.n419 GND.n418 585
R935 GND.n7737 GND.n7736 585
R936 GND.n7736 GND.n7735 585
R937 GND.n423 GND.n422 585
R938 GND.n7734 GND.n423 585
R939 GND.n7732 GND.n7731 585
R940 GND.n7733 GND.n7732 585
R941 GND.n426 GND.n425 585
R942 GND.n425 GND.n424 585
R943 GND.n7727 GND.n7726 585
R944 GND.n7726 GND.n7725 585
R945 GND.n429 GND.n428 585
R946 GND.n7724 GND.n429 585
R947 GND.n7722 GND.n7721 585
R948 GND.n7723 GND.n7722 585
R949 GND.n432 GND.n431 585
R950 GND.n431 GND.n430 585
R951 GND.n7717 GND.n7716 585
R952 GND.n7716 GND.n7715 585
R953 GND.n435 GND.n434 585
R954 GND.n7714 GND.n435 585
R955 GND.n7712 GND.n7711 585
R956 GND.n7713 GND.n7712 585
R957 GND.n438 GND.n437 585
R958 GND.n437 GND.n436 585
R959 GND.n7707 GND.n7706 585
R960 GND.n7706 GND.n7705 585
R961 GND.n441 GND.n440 585
R962 GND.n7704 GND.n441 585
R963 GND.n7702 GND.n7701 585
R964 GND.n7703 GND.n7702 585
R965 GND.n444 GND.n443 585
R966 GND.n443 GND.n442 585
R967 GND.n7697 GND.n7696 585
R968 GND.n7696 GND.n7695 585
R969 GND.n447 GND.n446 585
R970 GND.n7694 GND.n447 585
R971 GND.n7692 GND.n7691 585
R972 GND.n7693 GND.n7692 585
R973 GND.n450 GND.n449 585
R974 GND.n449 GND.n448 585
R975 GND.n7687 GND.n7686 585
R976 GND.n7686 GND.n7685 585
R977 GND.n453 GND.n452 585
R978 GND.n7684 GND.n453 585
R979 GND.n7682 GND.n7681 585
R980 GND.n7683 GND.n7682 585
R981 GND.n456 GND.n455 585
R982 GND.n455 GND.n454 585
R983 GND.n7677 GND.n7676 585
R984 GND.n7676 GND.n7675 585
R985 GND.n459 GND.n458 585
R986 GND.n7674 GND.n459 585
R987 GND.n7672 GND.n7671 585
R988 GND.n7673 GND.n7672 585
R989 GND.n462 GND.n461 585
R990 GND.n461 GND.n460 585
R991 GND.n7667 GND.n7666 585
R992 GND.n7666 GND.n7665 585
R993 GND.n465 GND.n464 585
R994 GND.n7664 GND.n465 585
R995 GND.n7662 GND.n7661 585
R996 GND.n7663 GND.n7662 585
R997 GND.n468 GND.n467 585
R998 GND.n467 GND.n466 585
R999 GND.n7657 GND.n7656 585
R1000 GND.n7656 GND.n7655 585
R1001 GND.n471 GND.n470 585
R1002 GND.n7654 GND.n471 585
R1003 GND.n7652 GND.n7651 585
R1004 GND.n7653 GND.n7652 585
R1005 GND.n474 GND.n473 585
R1006 GND.n473 GND.n472 585
R1007 GND.n7647 GND.n7646 585
R1008 GND.n7646 GND.n7645 585
R1009 GND.n477 GND.n476 585
R1010 GND.n7644 GND.n477 585
R1011 GND.n7642 GND.n7641 585
R1012 GND.n7643 GND.n7642 585
R1013 GND.n480 GND.n479 585
R1014 GND.n479 GND.n478 585
R1015 GND.n7637 GND.n7636 585
R1016 GND.n7636 GND.n7635 585
R1017 GND.n483 GND.n482 585
R1018 GND.n7634 GND.n483 585
R1019 GND.n7632 GND.n7631 585
R1020 GND.n7633 GND.n7632 585
R1021 GND.n486 GND.n485 585
R1022 GND.n485 GND.n484 585
R1023 GND.n7627 GND.n7626 585
R1024 GND.n7626 GND.n7625 585
R1025 GND.n489 GND.n488 585
R1026 GND.n7624 GND.n489 585
R1027 GND.n7622 GND.n7621 585
R1028 GND.n7623 GND.n7622 585
R1029 GND.n492 GND.n491 585
R1030 GND.n491 GND.n490 585
R1031 GND.n7617 GND.n7616 585
R1032 GND.n7616 GND.n7615 585
R1033 GND.n495 GND.n494 585
R1034 GND.n7614 GND.n495 585
R1035 GND.n7612 GND.n7611 585
R1036 GND.n7613 GND.n7612 585
R1037 GND.n498 GND.n497 585
R1038 GND.n497 GND.n496 585
R1039 GND.n7607 GND.n7606 585
R1040 GND.n7606 GND.n7605 585
R1041 GND.n501 GND.n500 585
R1042 GND.n7604 GND.n501 585
R1043 GND.n7602 GND.n7601 585
R1044 GND.n7603 GND.n7602 585
R1045 GND.n504 GND.n503 585
R1046 GND.n503 GND.n502 585
R1047 GND.n7597 GND.n7596 585
R1048 GND.n7596 GND.n7595 585
R1049 GND.n507 GND.n506 585
R1050 GND.n7594 GND.n507 585
R1051 GND.n144 GND.n143 585
R1052 GND.n7875 GND.n144 585
R1053 GND.n8019 GND.n8018 585
R1054 GND.n8018 GND.n8017 585
R1055 GND.n8020 GND.n139 585
R1056 GND.n5300 GND.n139 585
R1057 GND.n8022 GND.n8021 585
R1058 GND.n8023 GND.n8022 585
R1059 GND.n123 GND.n122 585
R1060 GND.n5306 GND.n123 585
R1061 GND.n8031 GND.n8030 585
R1062 GND.n8030 GND.n8029 585
R1063 GND.n8032 GND.n118 585
R1064 GND.n5312 GND.n118 585
R1065 GND.n8034 GND.n8033 585
R1066 GND.n8035 GND.n8034 585
R1067 GND.n102 GND.n101 585
R1068 GND.n5318 GND.n102 585
R1069 GND.n8043 GND.n8042 585
R1070 GND.n8042 GND.n8041 585
R1071 GND.n8044 GND.n97 585
R1072 GND.n5324 GND.n97 585
R1073 GND.n8046 GND.n8045 585
R1074 GND.n8047 GND.n8046 585
R1075 GND.n81 GND.n80 585
R1076 GND.n5330 GND.n81 585
R1077 GND.n8055 GND.n8054 585
R1078 GND.n8054 GND.n8053 585
R1079 GND.n8056 GND.n76 585
R1080 GND.n5336 GND.n76 585
R1081 GND.n8058 GND.n8057 585
R1082 GND.n8059 GND.n8058 585
R1083 GND.n61 GND.n60 585
R1084 GND.n5342 GND.n61 585
R1085 GND.n8067 GND.n8066 585
R1086 GND.n8066 GND.n8065 585
R1087 GND.n8068 GND.n55 585
R1088 GND.n5348 GND.n55 585
R1089 GND.n8070 GND.n8069 585
R1090 GND.n8071 GND.n8070 585
R1091 GND.n56 GND.n54 585
R1092 GND.n5354 GND.n54 585
R1093 GND.n5360 GND.n5359 585
R1094 GND.n5363 GND.n5360 585
R1095 GND.n2557 GND.n2556 585
R1096 GND.n2556 GND.n2552 585
R1097 GND.n5131 GND.n35 585
R1098 GND.n8078 GND.n35 585
R1099 GND.n5130 GND.n5129 585
R1100 GND.n5129 GND.n2545 585
R1101 GND.n2537 GND.n2536 585
R1102 GND.n5373 GND.n2537 585
R1103 GND.n5378 GND.n5377 585
R1104 GND.n5377 GND.n5376 585
R1105 GND.n5379 GND.n2532 585
R1106 GND.n5122 GND.n2532 585
R1107 GND.n5381 GND.n5380 585
R1108 GND.n5382 GND.n5381 585
R1109 GND.n2518 GND.n2517 585
R1110 GND.n5110 GND.n2518 585
R1111 GND.n5390 GND.n5389 585
R1112 GND.n5389 GND.n5388 585
R1113 GND.n5391 GND.n2513 585
R1114 GND.n5103 GND.n2513 585
R1115 GND.n5393 GND.n5392 585
R1116 GND.n5394 GND.n5393 585
R1117 GND.n2497 GND.n2496 585
R1118 GND.n5095 GND.n2497 585
R1119 GND.n5402 GND.n5401 585
R1120 GND.n5401 GND.n5400 585
R1121 GND.n5403 GND.n2492 585
R1122 GND.n5088 GND.n2492 585
R1123 GND.n5405 GND.n5404 585
R1124 GND.n5406 GND.n5405 585
R1125 GND.n2476 GND.n2475 585
R1126 GND.n5080 GND.n2476 585
R1127 GND.n5414 GND.n5413 585
R1128 GND.n5413 GND.n5412 585
R1129 GND.n5415 GND.n2471 585
R1130 GND.n5073 GND.n2471 585
R1131 GND.n5417 GND.n5416 585
R1132 GND.n5418 GND.n5417 585
R1133 GND.n2456 GND.n2455 585
R1134 GND.n5065 GND.n2456 585
R1135 GND.n5426 GND.n5425 585
R1136 GND.n5425 GND.n5424 585
R1137 GND.n5427 GND.n2450 585
R1138 GND.n5058 GND.n2450 585
R1139 GND.n5429 GND.n5428 585
R1140 GND.n5430 GND.n5429 585
R1141 GND.n2451 GND.n2434 585
R1142 GND.n5050 GND.n2434 585
R1143 GND.n5437 GND.n2435 585
R1144 GND.n5437 GND.n5436 585
R1145 GND.n5438 GND.n2400 585
R1146 GND.n5439 GND.n5438 585
R1147 GND.n2433 GND.n2432 585
R1148 GND.n2431 GND.n2430 585
R1149 GND.n2429 GND.n2428 585
R1150 GND.n2427 GND.n2426 585
R1151 GND.n2425 GND.n2424 585
R1152 GND.n2423 GND.n2422 585
R1153 GND.n2421 GND.n2420 585
R1154 GND.n2419 GND.n2418 585
R1155 GND.n2417 GND.n2416 585
R1156 GND.n2266 GND.n2264 585
R1157 GND.n5591 GND.n5590 585
R1158 GND.n2267 GND.n2265 585
R1159 GND.n5031 GND.n5030 585
R1160 GND.n5034 GND.n5033 585
R1161 GND.n5032 GND.n2665 585
R1162 GND.n5039 GND.n2666 585
R1163 GND.n5040 GND.n2662 585
R1164 GND.n5042 GND.n5041 585
R1165 GND.n5293 GND.n5292 585
R1166 GND.n5290 GND.n5234 585
R1167 GND.n5289 GND.n5288 585
R1168 GND.n5282 GND.n5236 585
R1169 GND.n5284 GND.n5283 585
R1170 GND.n5280 GND.n5238 585
R1171 GND.n5279 GND.n5278 585
R1172 GND.n5272 GND.n5240 585
R1173 GND.n5274 GND.n5273 585
R1174 GND.n5270 GND.n5242 585
R1175 GND.n5269 GND.n5268 585
R1176 GND.n5262 GND.n5244 585
R1177 GND.n5264 GND.n5263 585
R1178 GND.n5260 GND.n5246 585
R1179 GND.n5259 GND.n5258 585
R1180 GND.n5252 GND.n5248 585
R1181 GND.n5254 GND.n5253 585
R1182 GND.n5250 GND.n5249 585
R1183 GND.n5296 GND.n290 585
R1184 GND.n7875 GND.n290 585
R1185 GND.n5297 GND.n147 585
R1186 GND.n8017 GND.n147 585
R1187 GND.n5302 GND.n5301 585
R1188 GND.n5301 GND.n5300 585
R1189 GND.n5303 GND.n137 585
R1190 GND.n8023 GND.n137 585
R1191 GND.n5305 GND.n5304 585
R1192 GND.n5306 GND.n5305 585
R1193 GND.n5223 GND.n126 585
R1194 GND.n8029 GND.n126 585
R1195 GND.n5314 GND.n5313 585
R1196 GND.n5313 GND.n5312 585
R1197 GND.n5315 GND.n116 585
R1198 GND.n8035 GND.n116 585
R1199 GND.n5317 GND.n5316 585
R1200 GND.n5318 GND.n5317 585
R1201 GND.n5216 GND.n105 585
R1202 GND.n8041 GND.n105 585
R1203 GND.n5326 GND.n5325 585
R1204 GND.n5325 GND.n5324 585
R1205 GND.n5327 GND.n95 585
R1206 GND.n8047 GND.n95 585
R1207 GND.n5329 GND.n5328 585
R1208 GND.n5330 GND.n5329 585
R1209 GND.n5209 GND.n84 585
R1210 GND.n8053 GND.n84 585
R1211 GND.n5338 GND.n5337 585
R1212 GND.n5337 GND.n5336 585
R1213 GND.n5339 GND.n74 585
R1214 GND.n8059 GND.n74 585
R1215 GND.n5341 GND.n5340 585
R1216 GND.n5342 GND.n5341 585
R1217 GND.n5142 GND.n64 585
R1218 GND.n8065 GND.n64 585
R1219 GND.n5350 GND.n5349 585
R1220 GND.n5349 GND.n5348 585
R1221 GND.n5351 GND.n53 585
R1222 GND.n8071 GND.n53 585
R1223 GND.n5353 GND.n5352 585
R1224 GND.n5354 GND.n5353 585
R1225 GND.n5137 GND.n2554 585
R1226 GND.n5363 GND.n2554 585
R1227 GND.n31 GND.n29 585
R1228 GND.n2552 GND.n31 585
R1229 GND.n8080 GND.n8079 585
R1230 GND.n8079 GND.n8078 585
R1231 GND.n30 GND.n28 585
R1232 GND.n2545 GND.n30 585
R1233 GND.n5118 GND.n2544 585
R1234 GND.n5373 GND.n2544 585
R1235 GND.n5119 GND.n2540 585
R1236 GND.n5376 GND.n2540 585
R1237 GND.n5121 GND.n5120 585
R1238 GND.n5122 GND.n5121 585
R1239 GND.n2563 GND.n2530 585
R1240 GND.n5382 GND.n2530 585
R1241 GND.n5112 GND.n5111 585
R1242 GND.n5111 GND.n5110 585
R1243 GND.n2565 GND.n2521 585
R1244 GND.n5388 GND.n2521 585
R1245 GND.n5102 GND.n5101 585
R1246 GND.n5103 GND.n5102 585
R1247 GND.n2567 GND.n2511 585
R1248 GND.n5394 GND.n2511 585
R1249 GND.n5097 GND.n5096 585
R1250 GND.n5096 GND.n5095 585
R1251 GND.n2569 GND.n2500 585
R1252 GND.n5400 GND.n2500 585
R1253 GND.n5087 GND.n5086 585
R1254 GND.n5088 GND.n5087 585
R1255 GND.n2571 GND.n2490 585
R1256 GND.n5406 GND.n2490 585
R1257 GND.n5082 GND.n5081 585
R1258 GND.n5081 GND.n5080 585
R1259 GND.n2573 GND.n2479 585
R1260 GND.n5412 GND.n2479 585
R1261 GND.n5072 GND.n5071 585
R1262 GND.n5073 GND.n5072 585
R1263 GND.n2575 GND.n2469 585
R1264 GND.n5418 GND.n2469 585
R1265 GND.n5067 GND.n5066 585
R1266 GND.n5066 GND.n5065 585
R1267 GND.n2577 GND.n2459 585
R1268 GND.n5424 GND.n2459 585
R1269 GND.n5057 GND.n5056 585
R1270 GND.n5058 GND.n5057 585
R1271 GND.n2659 GND.n2448 585
R1272 GND.n5430 GND.n2448 585
R1273 GND.n5052 GND.n5051 585
R1274 GND.n5051 GND.n5050 585
R1275 GND.n5046 GND.n2436 585
R1276 GND.n5436 GND.n2436 585
R1277 GND.n5045 GND.n2405 585
R1278 GND.n5439 GND.n2405 585
R1279 GND.n2236 GND.n2233 585
R1280 GND.n2233 GND.n2218 585
R1281 GND.n2203 GND.n2202 585
R1282 GND.n2206 GND.n2203 585
R1283 GND.n5654 GND.n5653 585
R1284 GND.n5653 GND.n5652 585
R1285 GND.n5655 GND.n2195 585
R1286 GND.n5014 GND.n2195 585
R1287 GND.n5657 GND.n5656 585
R1288 GND.n5658 GND.n5657 585
R1289 GND.n2196 GND.n2194 585
R1290 GND.n2194 GND.n2191 585
R1291 GND.n2177 GND.n2176 585
R1292 GND.n2179 GND.n2177 585
R1293 GND.n5668 GND.n5667 585
R1294 GND.n5667 GND.n5666 585
R1295 GND.n5669 GND.n2169 585
R1296 GND.n5003 GND.n2169 585
R1297 GND.n5671 GND.n5670 585
R1298 GND.n5672 GND.n5671 585
R1299 GND.n2170 GND.n2168 585
R1300 GND.n2168 GND.n2165 585
R1301 GND.n2150 GND.n2149 585
R1302 GND.n2153 GND.n2150 585
R1303 GND.n5682 GND.n5681 585
R1304 GND.n5681 GND.n5680 585
R1305 GND.n5683 GND.n2142 585
R1306 GND.n4991 GND.n2142 585
R1307 GND.n5685 GND.n5684 585
R1308 GND.n5686 GND.n5685 585
R1309 GND.n2143 GND.n2141 585
R1310 GND.n2141 GND.n2138 585
R1311 GND.n2123 GND.n2122 585
R1312 GND.n2126 GND.n2123 585
R1313 GND.n5696 GND.n5695 585
R1314 GND.n5695 GND.n5694 585
R1315 GND.n5697 GND.n2115 585
R1316 GND.n2679 GND.n2115 585
R1317 GND.n5699 GND.n5698 585
R1318 GND.n5700 GND.n5699 585
R1319 GND.n2116 GND.n2114 585
R1320 GND.n2114 GND.n2111 585
R1321 GND.n2096 GND.n2095 585
R1322 GND.n2099 GND.n2096 585
R1323 GND.n5710 GND.n5709 585
R1324 GND.n5709 GND.n5708 585
R1325 GND.n5711 GND.n2088 585
R1326 GND.n4969 GND.n2088 585
R1327 GND.n5713 GND.n5712 585
R1328 GND.n5714 GND.n5713 585
R1329 GND.n2089 GND.n2087 585
R1330 GND.n2087 GND.n2084 585
R1331 GND.n2069 GND.n2068 585
R1332 GND.n2072 GND.n2069 585
R1333 GND.n5724 GND.n5723 585
R1334 GND.n5723 GND.n5722 585
R1335 GND.n5725 GND.n2061 585
R1336 GND.n4958 GND.n2061 585
R1337 GND.n5727 GND.n5726 585
R1338 GND.n5728 GND.n5727 585
R1339 GND.n2062 GND.n2060 585
R1340 GND.n2060 GND.n2057 585
R1341 GND.n2042 GND.n2041 585
R1342 GND.n2045 GND.n2042 585
R1343 GND.n5738 GND.n5737 585
R1344 GND.n5737 GND.n5736 585
R1345 GND.n5739 GND.n2034 585
R1346 GND.n4947 GND.n2034 585
R1347 GND.n5741 GND.n5740 585
R1348 GND.n5742 GND.n5741 585
R1349 GND.n2035 GND.n2033 585
R1350 GND.n2033 GND.n2030 585
R1351 GND.n2015 GND.n2014 585
R1352 GND.n2018 GND.n2015 585
R1353 GND.n5752 GND.n5751 585
R1354 GND.n5751 GND.n5750 585
R1355 GND.n5753 GND.n2007 585
R1356 GND.n2692 GND.n2007 585
R1357 GND.n5755 GND.n5754 585
R1358 GND.n5756 GND.n5755 585
R1359 GND.n2008 GND.n2006 585
R1360 GND.n2006 GND.n2004 585
R1361 GND.n1989 GND.n1988 585
R1362 GND.n1992 GND.n1989 585
R1363 GND.n5766 GND.n5765 585
R1364 GND.n5765 GND.n5764 585
R1365 GND.n5767 GND.n1981 585
R1366 GND.n4925 GND.n1981 585
R1367 GND.n5769 GND.n5768 585
R1368 GND.n5770 GND.n5769 585
R1369 GND.n1982 GND.n1980 585
R1370 GND.n1980 GND.n1977 585
R1371 GND.n1962 GND.n1961 585
R1372 GND.n1965 GND.n1962 585
R1373 GND.n5780 GND.n5779 585
R1374 GND.n5779 GND.n5778 585
R1375 GND.n5781 GND.n1954 585
R1376 GND.n4914 GND.n1954 585
R1377 GND.n5783 GND.n5782 585
R1378 GND.n5784 GND.n5783 585
R1379 GND.n1955 GND.n1953 585
R1380 GND.n1953 GND.n1950 585
R1381 GND.n1935 GND.n1934 585
R1382 GND.n1938 GND.n1935 585
R1383 GND.n5794 GND.n5793 585
R1384 GND.n5793 GND.n5792 585
R1385 GND.n5795 GND.n1927 585
R1386 GND.n4903 GND.n1927 585
R1387 GND.n5797 GND.n5796 585
R1388 GND.n5798 GND.n5797 585
R1389 GND.n1928 GND.n1926 585
R1390 GND.n1926 GND.n1923 585
R1391 GND.n1911 GND.n1910 585
R1392 GND.n1914 GND.n1911 585
R1393 GND.n5808 GND.n5807 585
R1394 GND.n5807 GND.n5806 585
R1395 GND.n5809 GND.n1905 585
R1396 GND.n1905 GND.n1871 585
R1397 GND.n5811 GND.n5810 585
R1398 GND.n5811 GND.n1852 585
R1399 GND.n5812 GND.n1904 585
R1400 GND.n5812 GND.n1844 585
R1401 GND.n5814 GND.n5813 585
R1402 GND.n5813 GND.n1842 585
R1403 GND.n5815 GND.n1899 585
R1404 GND.n1899 GND.n1836 585
R1405 GND.n5817 GND.n5816 585
R1406 GND.n5818 GND.n5817 585
R1407 GND.n1900 GND.n1898 585
R1408 GND.n4879 GND.n1898 585
R1409 GND.n4876 GND.n4875 585
R1410 GND.n4877 GND.n4876 585
R1411 GND.n2715 GND.n2714 585
R1412 GND.n2714 GND.n1819 585
R1413 GND.n4870 GND.n4869 585
R1414 GND.n4869 GND.n4868 585
R1415 GND.n2718 GND.n2717 585
R1416 GND.n2723 GND.n2718 585
R1417 GND.n4853 GND.n2731 585
R1418 GND.n2731 GND.n1807 585
R1419 GND.n4855 GND.n4854 585
R1420 GND.n4856 GND.n4855 585
R1421 GND.n2732 GND.n2730 585
R1422 GND.n4841 GND.n2730 585
R1423 GND.n4848 GND.n4847 585
R1424 GND.n4847 GND.n4846 585
R1425 GND.n2735 GND.n2734 585
R1426 GND.n2735 GND.n1790 585
R1427 GND.n4805 GND.n4790 585
R1428 GND.n4790 GND.n1784 585
R1429 GND.n4807 GND.n4806 585
R1430 GND.n4808 GND.n4807 585
R1431 GND.n4791 GND.n4789 585
R1432 GND.n4789 GND.n2741 585
R1433 GND.n4800 GND.n4799 585
R1434 GND.n4799 GND.n1772 585
R1435 GND.n4798 GND.n4793 585
R1436 GND.n4798 GND.n1766 585
R1437 GND.n4797 GND.n4796 585
R1438 GND.n4797 GND.n1764 585
R1439 GND.n1747 GND.n1746 585
R1440 GND.n2755 GND.n1747 585
R1441 GND.n6091 GND.n6090 585
R1442 GND.n6090 GND.n6089 585
R1443 GND.n6092 GND.n1733 585
R1444 GND.n4763 GND.n1733 585
R1445 GND.n6094 GND.n6093 585
R1446 GND.n6095 GND.n6094 585
R1447 GND.n1734 GND.n1732 585
R1448 GND.n1732 GND.n1722 585
R1449 GND.n1740 GND.n1739 585
R1450 GND.n1739 GND.n1720 585
R1451 GND.n1738 GND.n1737 585
R1452 GND.n1738 GND.n1705 585
R1453 GND.n1695 GND.n1694 585
R1454 GND.t40 GND.n1695 585
R1455 GND.n6118 GND.n6117 585
R1456 GND.n6117 GND.n6116 585
R1457 GND.n6119 GND.n1684 585
R1458 GND.n4714 GND.n1684 585
R1459 GND.n6121 GND.n6120 585
R1460 GND.n6122 GND.n6121 585
R1461 GND.n1685 GND.n1683 585
R1462 GND.n4691 GND.n1683 585
R1463 GND.n1688 GND.n1687 585
R1464 GND.n1687 GND.n1671 585
R1465 GND.n1660 GND.n1659 585
R1466 GND.n1669 GND.n1660 585
R1467 GND.n6139 GND.n6138 585
R1468 GND.n6138 GND.n6137 585
R1469 GND.n6140 GND.n1654 585
R1470 GND.n4666 GND.n1654 585
R1471 GND.n6142 GND.n6141 585
R1472 GND.n6143 GND.n6142 585
R1473 GND.n1655 GND.n1653 585
R1474 GND.n4653 GND.n1653 585
R1475 GND.n4574 GND.n2780 585
R1476 GND.n2780 GND.n1578 585
R1477 GND.n4576 GND.n4575 585
R1478 GND.n4577 GND.n4576 585
R1479 GND.n2781 GND.n2779 585
R1480 GND.n2787 GND.n2779 585
R1481 GND.n4568 GND.n4567 585
R1482 GND.n4567 GND.n4566 585
R1483 GND.n2784 GND.n2783 585
R1484 GND.n4538 GND.n2784 585
R1485 GND.n4522 GND.n2803 585
R1486 GND.n2803 GND.n2794 585
R1487 GND.n4524 GND.n4523 585
R1488 GND.n4525 GND.n4524 585
R1489 GND.n2804 GND.n2802 585
R1490 GND.n2810 GND.n2802 585
R1491 GND.n4517 GND.n4516 585
R1492 GND.n4516 GND.n4515 585
R1493 GND.n2807 GND.n2806 585
R1494 GND.n4503 GND.n2807 585
R1495 GND.n4490 GND.n2826 585
R1496 GND.n2826 GND.n2817 585
R1497 GND.n4492 GND.n4491 585
R1498 GND.n4493 GND.n4492 585
R1499 GND.n2827 GND.n2825 585
R1500 GND.n2833 GND.n2825 585
R1501 GND.n4485 GND.n4484 585
R1502 GND.n4484 GND.n4483 585
R1503 GND.n2830 GND.n2829 585
R1504 GND.n4471 GND.n2830 585
R1505 GND.n4458 GND.n2849 585
R1506 GND.n2849 GND.n2840 585
R1507 GND.n4460 GND.n4459 585
R1508 GND.n4461 GND.n4460 585
R1509 GND.n2850 GND.n2848 585
R1510 GND.n2856 GND.n2848 585
R1511 GND.n4453 GND.n4452 585
R1512 GND.n4452 GND.n4451 585
R1513 GND.n2853 GND.n2852 585
R1514 GND.n4439 GND.n2853 585
R1515 GND.n4426 GND.n2872 585
R1516 GND.n2872 GND.n2863 585
R1517 GND.n4428 GND.n4427 585
R1518 GND.n4429 GND.n4428 585
R1519 GND.n2873 GND.n2871 585
R1520 GND.n2879 GND.n2871 585
R1521 GND.n4421 GND.n4420 585
R1522 GND.n4420 GND.n4419 585
R1523 GND.n2876 GND.n2875 585
R1524 GND.n4407 GND.n2876 585
R1525 GND.n4394 GND.n2895 585
R1526 GND.n2895 GND.n2886 585
R1527 GND.n4396 GND.n4395 585
R1528 GND.n4397 GND.n4396 585
R1529 GND.n2896 GND.n2894 585
R1530 GND.n2902 GND.n2894 585
R1531 GND.n4389 GND.n4388 585
R1532 GND.n4388 GND.n4387 585
R1533 GND.n2899 GND.n2898 585
R1534 GND.n4375 GND.n2899 585
R1535 GND.n4362 GND.n2918 585
R1536 GND.n2918 GND.n2909 585
R1537 GND.n4364 GND.n4363 585
R1538 GND.n4365 GND.n4364 585
R1539 GND.n2919 GND.n2917 585
R1540 GND.n2925 GND.n2917 585
R1541 GND.n4357 GND.n4356 585
R1542 GND.n4356 GND.n4355 585
R1543 GND.n2922 GND.n2921 585
R1544 GND.n4343 GND.n2922 585
R1545 GND.n4330 GND.n2941 585
R1546 GND.n2941 GND.n2940 585
R1547 GND.n4332 GND.n4331 585
R1548 GND.n4333 GND.n4332 585
R1549 GND.n2942 GND.n2939 585
R1550 GND.n2948 GND.n2939 585
R1551 GND.n4325 GND.n4324 585
R1552 GND.n4324 GND.n4323 585
R1553 GND.n2945 GND.n2944 585
R1554 GND.n4311 GND.n2945 585
R1555 GND.n4298 GND.n2964 585
R1556 GND.n2964 GND.n2955 585
R1557 GND.n4300 GND.n4299 585
R1558 GND.n4301 GND.n4300 585
R1559 GND.n2965 GND.n2963 585
R1560 GND.n2971 GND.n2963 585
R1561 GND.n4293 GND.n4292 585
R1562 GND.n4292 GND.n4291 585
R1563 GND.n2968 GND.n2967 585
R1564 GND.n4279 GND.n2968 585
R1565 GND.n4266 GND.n2987 585
R1566 GND.n2987 GND.n2978 585
R1567 GND.n4268 GND.n4267 585
R1568 GND.n4269 GND.n4268 585
R1569 GND.n2988 GND.n2986 585
R1570 GND.n2994 GND.n2986 585
R1571 GND.n4261 GND.n4260 585
R1572 GND.n4260 GND.n4259 585
R1573 GND.n2991 GND.n2990 585
R1574 GND.n4247 GND.n2991 585
R1575 GND.n4234 GND.n3010 585
R1576 GND.n3010 GND.n3001 585
R1577 GND.n4236 GND.n4235 585
R1578 GND.n4237 GND.n4236 585
R1579 GND.n3011 GND.n3009 585
R1580 GND.n3017 GND.n3009 585
R1581 GND.n4229 GND.n4228 585
R1582 GND.n4228 GND.n4227 585
R1583 GND.n3014 GND.n3013 585
R1584 GND.n4215 GND.n3014 585
R1585 GND.n4202 GND.n3033 585
R1586 GND.n3033 GND.n3024 585
R1587 GND.n4204 GND.n4203 585
R1588 GND.n4205 GND.n4204 585
R1589 GND.n3034 GND.n3032 585
R1590 GND.n3039 GND.n3032 585
R1591 GND.n4197 GND.n4196 585
R1592 GND.n4196 GND.n4195 585
R1593 GND.n3060 GND.n3036 585
R1594 GND.n4181 GND.n4180 585
R1595 GND.n4179 GND.n3059 585
R1596 GND.n4183 GND.n3059 585
R1597 GND.n4178 GND.n4177 585
R1598 GND.n4176 GND.n4175 585
R1599 GND.n4174 GND.n4173 585
R1600 GND.n4172 GND.n4171 585
R1601 GND.n4170 GND.n4169 585
R1602 GND.n4168 GND.n4167 585
R1603 GND.n4166 GND.n4165 585
R1604 GND.n4164 GND.n4163 585
R1605 GND.n4162 GND.n4161 585
R1606 GND.n3073 GND.n3071 585
R1607 GND.n3165 GND.n3074 585
R1608 GND.n3164 GND.n3075 585
R1609 GND.n3077 GND.n3076 585
R1610 GND.n3157 GND.n3085 585
R1611 GND.n3156 GND.n3086 585
R1612 GND.n3093 GND.n3087 585
R1613 GND.n3149 GND.n3094 585
R1614 GND.n3148 GND.n3095 585
R1615 GND.n3097 GND.n3096 585
R1616 GND.n3141 GND.n3105 585
R1617 GND.n3140 GND.n3137 585
R1618 GND.n3112 GND.n3106 585
R1619 GND.n3130 GND.n3113 585
R1620 GND.n3129 GND.n3114 585
R1621 GND.n5024 GND.n5023 585
R1622 GND.n5027 GND.n5026 585
R1623 GND.n5025 GND.n2259 585
R1624 GND.n5595 GND.n5594 585
R1625 GND.n5597 GND.n5596 585
R1626 GND.n5599 GND.n5598 585
R1627 GND.n5601 GND.n5600 585
R1628 GND.n5603 GND.n5602 585
R1629 GND.n5605 GND.n5604 585
R1630 GND.n5607 GND.n5606 585
R1631 GND.n5609 GND.n5608 585
R1632 GND.n5611 GND.n5610 585
R1633 GND.n5613 GND.n5612 585
R1634 GND.n5615 GND.n5614 585
R1635 GND.n5617 GND.n5616 585
R1636 GND.n5619 GND.n5618 585
R1637 GND.n5621 GND.n5620 585
R1638 GND.n5623 GND.n5622 585
R1639 GND.n5625 GND.n5624 585
R1640 GND.n5627 GND.n5626 585
R1641 GND.n5629 GND.n5628 585
R1642 GND.n5631 GND.n5630 585
R1643 GND.n5633 GND.n5632 585
R1644 GND.n5636 GND.n5635 585
R1645 GND.n5634 GND.n2239 585
R1646 GND.n5640 GND.n2234 585
R1647 GND.n5642 GND.n5641 585
R1648 GND.n5643 GND.n5642 585
R1649 GND.n5022 GND.n5021 585
R1650 GND.n5022 GND.n2218 585
R1651 GND.n5020 GND.n2670 585
R1652 GND.n2670 GND.n2206 585
R1653 GND.n2671 GND.n2205 585
R1654 GND.n5652 GND.n2205 585
R1655 GND.n5016 GND.n5015 585
R1656 GND.n5015 GND.n5014 585
R1657 GND.n5013 GND.n2192 585
R1658 GND.n5658 GND.n2192 585
R1659 GND.n5012 GND.n5011 585
R1660 GND.n5011 GND.n2191 585
R1661 GND.n5010 GND.n2673 585
R1662 GND.n5010 GND.n2179 585
R1663 GND.n5006 GND.n2178 585
R1664 GND.n5666 GND.n2178 585
R1665 GND.n5005 GND.n5004 585
R1666 GND.n5004 GND.n5003 585
R1667 GND.n5001 GND.n2166 585
R1668 GND.n5672 GND.n2166 585
R1669 GND.n4995 GND.n2675 585
R1670 GND.n4995 GND.n2165 585
R1671 GND.n4997 GND.n4996 585
R1672 GND.n4996 GND.n2153 585
R1673 GND.n4994 GND.n2152 585
R1674 GND.n5680 GND.n2152 585
R1675 GND.n4993 GND.n4992 585
R1676 GND.n4992 GND.n4991 585
R1677 GND.n2677 GND.n2139 585
R1678 GND.n5686 GND.n2139 585
R1679 GND.n4987 GND.n4986 585
R1680 GND.n4986 GND.n2138 585
R1681 GND.n4985 GND.n4984 585
R1682 GND.n4985 GND.n2126 585
R1683 GND.n4983 GND.n2125 585
R1684 GND.n5694 GND.n2125 585
R1685 GND.n2681 GND.n2680 585
R1686 GND.n2680 GND.n2679 585
R1687 GND.n4979 GND.n2112 585
R1688 GND.n5700 GND.n2112 585
R1689 GND.n4978 GND.n4977 585
R1690 GND.n4977 GND.n2111 585
R1691 GND.n4976 GND.n4975 585
R1692 GND.n4976 GND.n2099 585
R1693 GND.n2683 GND.n2098 585
R1694 GND.n5708 GND.n2098 585
R1695 GND.n4971 GND.n4970 585
R1696 GND.n4970 GND.n4969 585
R1697 GND.n4968 GND.n2085 585
R1698 GND.n5714 GND.n2085 585
R1699 GND.n4967 GND.n4966 585
R1700 GND.n4966 GND.n2084 585
R1701 GND.n4965 GND.n2685 585
R1702 GND.n4965 GND.n2072 585
R1703 GND.n4961 GND.n2071 585
R1704 GND.n5722 GND.n2071 585
R1705 GND.n4960 GND.n4959 585
R1706 GND.n4959 GND.n4958 585
R1707 GND.n4957 GND.n2058 585
R1708 GND.n5728 GND.n2058 585
R1709 GND.n4951 GND.n2687 585
R1710 GND.n4951 GND.n2057 585
R1711 GND.n4953 GND.n4952 585
R1712 GND.n4952 GND.n2045 585
R1713 GND.n4950 GND.n2044 585
R1714 GND.n5736 GND.n2044 585
R1715 GND.n4949 GND.n4948 585
R1716 GND.n4948 GND.n4947 585
R1717 GND.n2689 GND.n2031 585
R1718 GND.n5742 GND.n2031 585
R1719 GND.n4943 GND.n4942 585
R1720 GND.n4942 GND.n2030 585
R1721 GND.n4941 GND.n4940 585
R1722 GND.n4941 GND.n2018 585
R1723 GND.n4939 GND.n2017 585
R1724 GND.n5750 GND.n2017 585
R1725 GND.n2694 GND.n2693 585
R1726 GND.n2693 GND.n2692 585
R1727 GND.n4935 GND.n2005 585
R1728 GND.n5756 GND.n2005 585
R1729 GND.n4934 GND.n4933 585
R1730 GND.n4933 GND.n2004 585
R1731 GND.n4932 GND.n4931 585
R1732 GND.n4932 GND.n1992 585
R1733 GND.n2696 GND.n1991 585
R1734 GND.n5764 GND.n1991 585
R1735 GND.n4927 GND.n4926 585
R1736 GND.n4926 GND.n4925 585
R1737 GND.n4924 GND.n1978 585
R1738 GND.n5770 GND.n1978 585
R1739 GND.n4923 GND.n4922 585
R1740 GND.n4922 GND.n1977 585
R1741 GND.n4921 GND.n2698 585
R1742 GND.n4921 GND.n1965 585
R1743 GND.n4917 GND.n1964 585
R1744 GND.n5778 GND.n1964 585
R1745 GND.n4916 GND.n4915 585
R1746 GND.n4915 GND.n4914 585
R1747 GND.n4913 GND.n1951 585
R1748 GND.n5784 GND.n1951 585
R1749 GND.n4907 GND.n2700 585
R1750 GND.n4907 GND.n1950 585
R1751 GND.n4909 GND.n4908 585
R1752 GND.n4908 GND.n1938 585
R1753 GND.n4906 GND.n1937 585
R1754 GND.n5792 GND.n1937 585
R1755 GND.n4905 GND.n4904 585
R1756 GND.n4904 GND.n4903 585
R1757 GND.n2702 GND.n1924 585
R1758 GND.n5798 GND.n1924 585
R1759 GND.n4899 GND.n4898 585
R1760 GND.n4898 GND.n1923 585
R1761 GND.n4897 GND.n4896 585
R1762 GND.n4897 GND.n1914 585
R1763 GND.n4895 GND.n1913 585
R1764 GND.n5806 GND.n1913 585
R1765 GND.n4889 GND.n2704 585
R1766 GND.n4889 GND.n1871 585
R1767 GND.n4891 GND.n4890 585
R1768 GND.n4890 GND.n1852 585
R1769 GND.n4888 GND.n2706 585
R1770 GND.n4888 GND.n1844 585
R1771 GND.n4887 GND.n4886 585
R1772 GND.n4887 GND.n1842 585
R1773 GND.n2708 GND.n2707 585
R1774 GND.n2707 GND.n1836 585
R1775 GND.n4882 GND.n1897 585
R1776 GND.n5818 GND.n1897 585
R1777 GND.n4881 GND.n4880 585
R1778 GND.n4880 GND.n4879 585
R1779 GND.n4878 GND.n2710 585
R1780 GND.n4878 GND.n4877 585
R1781 GND.n4865 GND.n2711 585
R1782 GND.n2711 GND.n1819 585
R1783 GND.n4867 GND.n4866 585
R1784 GND.n4868 GND.n4867 585
R1785 GND.n2725 GND.n2724 585
R1786 GND.n2724 GND.n2723 585
R1787 GND.n4859 GND.n4858 585
R1788 GND.n4858 GND.n1807 585
R1789 GND.n4857 GND.n2727 585
R1790 GND.n4857 GND.n4856 585
R1791 GND.n4782 GND.n2728 585
R1792 GND.n4841 GND.n2728 585
R1793 GND.n4783 GND.n2736 585
R1794 GND.n4846 GND.n2736 585
R1795 GND.n4785 GND.n4784 585
R1796 GND.n4784 GND.n1790 585
R1797 GND.n4786 GND.n2743 585
R1798 GND.n2743 GND.n1784 585
R1799 GND.n4788 GND.n4787 585
R1800 GND.n4808 GND.n4788 585
R1801 GND.n2744 GND.n2742 585
R1802 GND.n2742 GND.n2741 585
R1803 GND.n4774 GND.n4773 585
R1804 GND.n4773 GND.n1772 585
R1805 GND.n4772 GND.n2746 585
R1806 GND.n4772 GND.n1766 585
R1807 GND.n4771 GND.n4770 585
R1808 GND.n4771 GND.n1764 585
R1809 GND.n2748 GND.n2747 585
R1810 GND.n2755 GND.n2747 585
R1811 GND.n4766 GND.n1749 585
R1812 GND.n6089 GND.n1749 585
R1813 GND.n4765 GND.n4764 585
R1814 GND.n4764 GND.n4763 585
R1815 GND.n2750 GND.n1730 585
R1816 GND.n6095 GND.n1730 585
R1817 GND.n4705 GND.n4700 585
R1818 GND.n4700 GND.n1722 585
R1819 GND.n4707 GND.n4706 585
R1820 GND.n4707 GND.n1720 585
R1821 GND.n4708 GND.n4699 585
R1822 GND.n4708 GND.n1705 585
R1823 GND.n4710 GND.n4709 585
R1824 GND.n4709 GND.t40 585
R1825 GND.n4711 GND.n1697 585
R1826 GND.n6116 GND.n1697 585
R1827 GND.n4713 GND.n4712 585
R1828 GND.n4714 GND.n4713 585
R1829 GND.n2761 GND.n1681 585
R1830 GND.n6122 GND.n1681 585
R1831 GND.n4693 GND.n4692 585
R1832 GND.n4692 GND.n4691 585
R1833 GND.n2764 GND.n2763 585
R1834 GND.n2764 GND.n1671 585
R1835 GND.n4662 GND.n4661 585
R1836 GND.n4661 GND.n1669 585
R1837 GND.n4663 GND.n1662 585
R1838 GND.n6137 GND.n1662 585
R1839 GND.n4665 GND.n4664 585
R1840 GND.n4666 GND.n4665 585
R1841 GND.n2772 GND.n1651 585
R1842 GND.n6143 GND.n1651 585
R1843 GND.n4655 GND.n4654 585
R1844 GND.n4654 GND.n4653 585
R1845 GND.n4579 GND.n2774 585
R1846 GND.n4579 GND.n1578 585
R1847 GND.n4578 GND.n2776 585
R1848 GND.n4578 GND.n4577 585
R1849 GND.n4534 GND.n2775 585
R1850 GND.n2787 GND.n2775 585
R1851 GND.n4535 GND.n2786 585
R1852 GND.n4566 GND.n2786 585
R1853 GND.n4537 GND.n4536 585
R1854 GND.n4538 GND.n4537 585
R1855 GND.n2796 GND.n2795 585
R1856 GND.n2795 GND.n2794 585
R1857 GND.n4527 GND.n4526 585
R1858 GND.n4526 GND.n4525 585
R1859 GND.n2799 GND.n2798 585
R1860 GND.n2810 GND.n2799 585
R1861 GND.n4500 GND.n2809 585
R1862 GND.n4515 GND.n2809 585
R1863 GND.n4502 GND.n4501 585
R1864 GND.n4503 GND.n4502 585
R1865 GND.n2819 GND.n2818 585
R1866 GND.n2818 GND.n2817 585
R1867 GND.n4495 GND.n4494 585
R1868 GND.n4494 GND.n4493 585
R1869 GND.n2822 GND.n2821 585
R1870 GND.n2833 GND.n2822 585
R1871 GND.n4468 GND.n2832 585
R1872 GND.n4483 GND.n2832 585
R1873 GND.n4470 GND.n4469 585
R1874 GND.n4471 GND.n4470 585
R1875 GND.n2842 GND.n2841 585
R1876 GND.n2841 GND.n2840 585
R1877 GND.n4463 GND.n4462 585
R1878 GND.n4462 GND.n4461 585
R1879 GND.n2845 GND.n2844 585
R1880 GND.n2856 GND.n2845 585
R1881 GND.n4436 GND.n2855 585
R1882 GND.n4451 GND.n2855 585
R1883 GND.n4438 GND.n4437 585
R1884 GND.n4439 GND.n4438 585
R1885 GND.n2865 GND.n2864 585
R1886 GND.n2864 GND.n2863 585
R1887 GND.n4431 GND.n4430 585
R1888 GND.n4430 GND.n4429 585
R1889 GND.n2868 GND.n2867 585
R1890 GND.n2879 GND.n2868 585
R1891 GND.n4404 GND.n2878 585
R1892 GND.n4419 GND.n2878 585
R1893 GND.n4406 GND.n4405 585
R1894 GND.n4407 GND.n4406 585
R1895 GND.n2888 GND.n2887 585
R1896 GND.n2887 GND.n2886 585
R1897 GND.n4399 GND.n4398 585
R1898 GND.n4398 GND.n4397 585
R1899 GND.n2891 GND.n2890 585
R1900 GND.n2902 GND.n2891 585
R1901 GND.n4372 GND.n2901 585
R1902 GND.n4387 GND.n2901 585
R1903 GND.n4374 GND.n4373 585
R1904 GND.n4375 GND.n4374 585
R1905 GND.n2911 GND.n2910 585
R1906 GND.n2910 GND.n2909 585
R1907 GND.n4367 GND.n4366 585
R1908 GND.n4366 GND.n4365 585
R1909 GND.n2914 GND.n2913 585
R1910 GND.n2925 GND.n2914 585
R1911 GND.n4340 GND.n2924 585
R1912 GND.n4355 GND.n2924 585
R1913 GND.n4342 GND.n4341 585
R1914 GND.n4343 GND.n4342 585
R1915 GND.n2933 GND.n2932 585
R1916 GND.n2940 GND.n2932 585
R1917 GND.n4335 GND.n4334 585
R1918 GND.n4334 GND.n4333 585
R1919 GND.n2936 GND.n2935 585
R1920 GND.n2948 GND.n2936 585
R1921 GND.n4308 GND.n2947 585
R1922 GND.n4323 GND.n2947 585
R1923 GND.n4310 GND.n4309 585
R1924 GND.n4311 GND.n4310 585
R1925 GND.n2957 GND.n2956 585
R1926 GND.n2956 GND.n2955 585
R1927 GND.n4303 GND.n4302 585
R1928 GND.n4302 GND.n4301 585
R1929 GND.n2960 GND.n2959 585
R1930 GND.n2971 GND.n2960 585
R1931 GND.n4276 GND.n2970 585
R1932 GND.n4291 GND.n2970 585
R1933 GND.n4278 GND.n4277 585
R1934 GND.n4279 GND.n4278 585
R1935 GND.n2980 GND.n2979 585
R1936 GND.n2979 GND.n2978 585
R1937 GND.n4271 GND.n4270 585
R1938 GND.n4270 GND.n4269 585
R1939 GND.n2983 GND.n2982 585
R1940 GND.n2994 GND.n2983 585
R1941 GND.n4244 GND.n2993 585
R1942 GND.n4259 GND.n2993 585
R1943 GND.n4246 GND.n4245 585
R1944 GND.n4247 GND.n4246 585
R1945 GND.n3003 GND.n3002 585
R1946 GND.n3002 GND.n3001 585
R1947 GND.n4239 GND.n4238 585
R1948 GND.n4238 GND.n4237 585
R1949 GND.n3006 GND.n3005 585
R1950 GND.n3017 GND.n3006 585
R1951 GND.n4212 GND.n3016 585
R1952 GND.n4227 GND.n3016 585
R1953 GND.n4214 GND.n4213 585
R1954 GND.n4215 GND.n4214 585
R1955 GND.n3026 GND.n3025 585
R1956 GND.n3025 GND.n3024 585
R1957 GND.n4207 GND.n4206 585
R1958 GND.n4206 GND.n4205 585
R1959 GND.n3029 GND.n3028 585
R1960 GND.n3039 GND.n3029 585
R1961 GND.n3120 GND.n3038 585
R1962 GND.n4195 GND.n3038 585
R1963 GND.n5938 GND.n5937 585
R1964 GND.n5939 GND.n5938 585
R1965 GND.n1841 GND.n1840 585
R1966 GND.n5833 GND.n1841 585
R1967 GND.n6021 GND.n6020 585
R1968 GND.n6020 GND.n6019 585
R1969 GND.n6022 GND.n1838 585
R1970 GND.n5827 GND.n1838 585
R1971 GND.n6024 GND.n6023 585
R1972 GND.n6025 GND.n6024 585
R1973 GND.n1839 GND.n1837 585
R1974 GND.n1837 GND.n1834 585
R1975 GND.n5820 GND.n5819 585
R1976 GND.n5821 GND.n5820 585
R1977 GND.n1824 GND.n1823 585
R1978 GND.n1826 GND.n1824 585
R1979 GND.n6035 GND.n6034 585
R1980 GND.n6034 GND.n6033 585
R1981 GND.n6036 GND.n1821 585
R1982 GND.n2713 GND.n1821 585
R1983 GND.n6038 GND.n6037 585
R1984 GND.n6039 GND.n6038 585
R1985 GND.n1822 GND.n1820 585
R1986 GND.n1820 GND.n1817 585
R1987 GND.n2720 GND.n2719 585
R1988 GND.n2721 GND.n2720 585
R1989 GND.n1806 GND.n1805 585
R1990 GND.n1809 GND.n1806 585
R1991 GND.n6049 GND.n6048 585
R1992 GND.n6048 GND.n6047 585
R1993 GND.n6050 GND.n1803 585
R1994 GND.n2729 GND.n1803 585
R1995 GND.n6052 GND.n6051 585
R1996 GND.n6053 GND.n6052 585
R1997 GND.n1804 GND.n1802 585
R1998 GND.n1802 GND.n1800 585
R1999 GND.n4844 GND.n4843 585
R2000 GND.n4845 GND.n4844 585
R2001 GND.n1789 GND.n1788 585
R2002 GND.n1792 GND.n1789 585
R2003 GND.n6063 GND.n6062 585
R2004 GND.n6062 GND.n6061 585
R2005 GND.n6064 GND.n1786 585
R2006 GND.n4818 GND.n1786 585
R2007 GND.n6066 GND.n6065 585
R2008 GND.n6067 GND.n6066 585
R2009 GND.n1787 GND.n1785 585
R2010 GND.n1785 GND.n1782 585
R2011 GND.n4811 GND.n4810 585
R2012 GND.n4812 GND.n4811 585
R2013 GND.n1771 GND.n1770 585
R2014 GND.n1774 GND.n1771 585
R2015 GND.n6077 GND.n6076 585
R2016 GND.n6076 GND.n6075 585
R2017 GND.n6078 GND.n1768 585
R2018 GND.n4747 GND.n1768 585
R2019 GND.n6080 GND.n6079 585
R2020 GND.n6081 GND.n6080 585
R2021 GND.n1769 GND.n1767 585
R2022 GND.n4753 GND.n1767 585
R2023 GND.n4756 GND.n2754 585
R2024 GND.n4756 GND.n4755 585
R2025 GND.n4758 GND.n4757 585
R2026 GND.n4757 GND.n1750 585
R2027 GND.n4759 GND.n2753 585
R2028 GND.n2753 GND.n1748 585
R2029 GND.n4761 GND.n4760 585
R2030 GND.n4762 GND.n4761 585
R2031 GND.n1727 GND.n1726 585
R2032 GND.n4735 GND.n1727 585
R2033 GND.n6098 GND.n6097 585
R2034 GND.n6097 GND.n6096 585
R2035 GND.n6099 GND.n1724 585
R2036 GND.n4731 GND.n1724 585
R2037 GND.n6101 GND.n6100 585
R2038 GND.n6102 GND.n6101 585
R2039 GND.n1725 GND.n1723 585
R2040 GND.n4727 GND.n1723 585
R2041 GND.n1704 GND.n1703 585
R2042 GND.n4725 GND.n1704 585
R2043 GND.n6111 GND.n6110 585
R2044 GND.n6110 GND.n6109 585
R2045 GND.n6112 GND.n1701 585
R2046 GND.n4719 GND.n1701 585
R2047 GND.n6114 GND.n6113 585
R2048 GND.n6115 GND.n6114 585
R2049 GND.n1702 GND.n1700 585
R2050 GND.n4715 GND.n1700 585
R2051 GND.n4684 GND.n4683 585
R2052 GND.n4684 GND.n2760 585
R2053 GND.n4686 GND.n4685 585
R2054 GND.n4685 GND.n1682 585
R2055 GND.n4687 GND.n4682 585
R2056 GND.n4682 GND.n1680 585
R2057 GND.n4689 GND.n4688 585
R2058 GND.n4690 GND.n4689 585
R2059 GND.n1668 GND.n1667 585
R2060 GND.n2766 GND.n1668 585
R2061 GND.n6132 GND.n6131 585
R2062 GND.n6131 GND.n6130 585
R2063 GND.n6133 GND.n1665 585
R2064 GND.n4672 GND.n1665 585
R2065 GND.n6135 GND.n6134 585
R2066 GND.n6136 GND.n6135 585
R2067 GND.n1666 GND.n1664 585
R2068 GND.n4667 GND.n1664 585
R2069 GND.n1648 GND.n1647 585
R2070 GND.n2771 GND.n1648 585
R2071 GND.n6146 GND.n6145 585
R2072 GND.n6145 GND.n6144 585
R2073 GND.n6147 GND.n1616 585
R2074 GND.n4652 GND.n1616 585
R2075 GND.n6213 GND.n6212 585
R2076 GND.n6211 GND.n1615 585
R2077 GND.n6210 GND.n1614 585
R2078 GND.n6215 GND.n1614 585
R2079 GND.n6209 GND.n6208 585
R2080 GND.n6207 GND.n6206 585
R2081 GND.n6205 GND.n6204 585
R2082 GND.n6203 GND.n6202 585
R2083 GND.n6201 GND.n6200 585
R2084 GND.n6199 GND.n6198 585
R2085 GND.n6197 GND.n6196 585
R2086 GND.n6195 GND.n6194 585
R2087 GND.n6193 GND.n6192 585
R2088 GND.n6191 GND.n6190 585
R2089 GND.n6189 GND.n6188 585
R2090 GND.n6187 GND.n6186 585
R2091 GND.n6185 GND.n6184 585
R2092 GND.n6183 GND.n6182 585
R2093 GND.n6181 GND.n6180 585
R2094 GND.n6179 GND.n6178 585
R2095 GND.n6177 GND.n6176 585
R2096 GND.n6175 GND.n6174 585
R2097 GND.n6173 GND.n6172 585
R2098 GND.n6171 GND.n6170 585
R2099 GND.n6169 GND.n6168 585
R2100 GND.n6167 GND.n6166 585
R2101 GND.n6165 GND.n6164 585
R2102 GND.n6163 GND.n6162 585
R2103 GND.n6161 GND.n6160 585
R2104 GND.n6159 GND.n6158 585
R2105 GND.n6157 GND.n6156 585
R2106 GND.n6155 GND.n6154 585
R2107 GND.n6153 GND.n6152 585
R2108 GND.n1577 GND.n1576 585
R2109 GND.n6218 GND.n6217 585
R2110 GND.n6219 GND.n1574 585
R2111 GND.n1595 GND.n1573 585
R2112 GND.n4584 GND.n4583 585
R2113 GND.n4586 GND.n4585 585
R2114 GND.n4589 GND.n4588 585
R2115 GND.n4591 GND.n4590 585
R2116 GND.n4593 GND.n4592 585
R2117 GND.n4595 GND.n4594 585
R2118 GND.n4597 GND.n4596 585
R2119 GND.n4599 GND.n4598 585
R2120 GND.n4601 GND.n4600 585
R2121 GND.n4603 GND.n4602 585
R2122 GND.n4605 GND.n4604 585
R2123 GND.n4607 GND.n4606 585
R2124 GND.n4609 GND.n4608 585
R2125 GND.n4611 GND.n4610 585
R2126 GND.n4613 GND.n4612 585
R2127 GND.n4615 GND.n4614 585
R2128 GND.n4617 GND.n4616 585
R2129 GND.n4619 GND.n4618 585
R2130 GND.n4621 GND.n4620 585
R2131 GND.n4623 GND.n4622 585
R2132 GND.n4625 GND.n4624 585
R2133 GND.n4627 GND.n4626 585
R2134 GND.n4629 GND.n4628 585
R2135 GND.n4631 GND.n4630 585
R2136 GND.n4633 GND.n4632 585
R2137 GND.n4635 GND.n4634 585
R2138 GND.n4637 GND.n4636 585
R2139 GND.n4639 GND.n4638 585
R2140 GND.n4641 GND.n4640 585
R2141 GND.n4643 GND.n4642 585
R2142 GND.n4645 GND.n4644 585
R2143 GND.n4647 GND.n4646 585
R2144 GND.n4648 GND.n4580 585
R2145 GND.n5942 GND.n5941 585
R2146 GND.n5944 GND.n5943 585
R2147 GND.n5946 GND.n5945 585
R2148 GND.n5948 GND.n5947 585
R2149 GND.n5950 GND.n5949 585
R2150 GND.n5952 GND.n5951 585
R2151 GND.n5954 GND.n5953 585
R2152 GND.n5956 GND.n5955 585
R2153 GND.n5958 GND.n5957 585
R2154 GND.n5960 GND.n5959 585
R2155 GND.n5962 GND.n5961 585
R2156 GND.n5964 GND.n5963 585
R2157 GND.n5966 GND.n5965 585
R2158 GND.n5968 GND.n5967 585
R2159 GND.n5970 GND.n5969 585
R2160 GND.n5972 GND.n5971 585
R2161 GND.n5974 GND.n5973 585
R2162 GND.n5976 GND.n5975 585
R2163 GND.n5978 GND.n5977 585
R2164 GND.n5980 GND.n5979 585
R2165 GND.n5982 GND.n5981 585
R2166 GND.n5984 GND.n5983 585
R2167 GND.n5986 GND.n5985 585
R2168 GND.n5988 GND.n5987 585
R2169 GND.n5990 GND.n5989 585
R2170 GND.n5992 GND.n5991 585
R2171 GND.n5994 GND.n5993 585
R2172 GND.n5996 GND.n5995 585
R2173 GND.n5998 GND.n5997 585
R2174 GND.n6000 GND.n5999 585
R2175 GND.n6002 GND.n6001 585
R2176 GND.n6005 GND.n6004 585
R2177 GND.n6007 GND.n6006 585
R2178 GND.n6009 GND.n6008 585
R2179 GND.n6011 GND.n6010 585
R2180 GND.n5867 GND.n1890 585
R2181 GND.n5869 GND.n5868 585
R2182 GND.n5871 GND.n5870 585
R2183 GND.n5873 GND.n5872 585
R2184 GND.n5876 GND.n5875 585
R2185 GND.n5878 GND.n5877 585
R2186 GND.n5880 GND.n5879 585
R2187 GND.n5882 GND.n5881 585
R2188 GND.n5884 GND.n5883 585
R2189 GND.n5886 GND.n5885 585
R2190 GND.n5888 GND.n5887 585
R2191 GND.n5890 GND.n5889 585
R2192 GND.n5892 GND.n5891 585
R2193 GND.n5894 GND.n5893 585
R2194 GND.n5896 GND.n5895 585
R2195 GND.n5898 GND.n5897 585
R2196 GND.n5900 GND.n5899 585
R2197 GND.n5902 GND.n5901 585
R2198 GND.n5904 GND.n5903 585
R2199 GND.n5906 GND.n5905 585
R2200 GND.n5908 GND.n5907 585
R2201 GND.n5910 GND.n5909 585
R2202 GND.n5912 GND.n5911 585
R2203 GND.n5914 GND.n5913 585
R2204 GND.n5916 GND.n5915 585
R2205 GND.n5918 GND.n5917 585
R2206 GND.n5920 GND.n5919 585
R2207 GND.n5922 GND.n5921 585
R2208 GND.n5924 GND.n5923 585
R2209 GND.n5926 GND.n5925 585
R2210 GND.n5928 GND.n5927 585
R2211 GND.n5930 GND.n5929 585
R2212 GND.n5932 GND.n5931 585
R2213 GND.n5934 GND.n5933 585
R2214 GND.n5935 GND.n5835 585
R2215 GND.n5940 GND.n1893 585
R2216 GND.n5940 GND.n5939 585
R2217 GND.n5832 GND.n5831 585
R2218 GND.n5833 GND.n5832 585
R2219 GND.n5830 GND.n1843 585
R2220 GND.n6019 GND.n1843 585
R2221 GND.n5829 GND.n5828 585
R2222 GND.n5828 GND.n5827 585
R2223 GND.n5825 GND.n1835 585
R2224 GND.n6025 GND.n1835 585
R2225 GND.n5824 GND.n5823 585
R2226 GND.n5823 GND.n1834 585
R2227 GND.n5822 GND.n1894 585
R2228 GND.n5822 GND.n5821 585
R2229 GND.n4824 GND.n1895 585
R2230 GND.n1895 GND.n1826 585
R2231 GND.n4825 GND.n1825 585
R2232 GND.n6033 GND.n1825 585
R2233 GND.n4827 GND.n4826 585
R2234 GND.n4826 GND.n2713 585
R2235 GND.n4828 GND.n1818 585
R2236 GND.n6039 GND.n1818 585
R2237 GND.n4830 GND.n4829 585
R2238 GND.n4830 GND.n1817 585
R2239 GND.n4831 GND.n4823 585
R2240 GND.n4831 GND.n2721 585
R2241 GND.n4833 GND.n4832 585
R2242 GND.n4832 GND.n1809 585
R2243 GND.n4834 GND.n1808 585
R2244 GND.n6047 GND.n1808 585
R2245 GND.n4836 GND.n4835 585
R2246 GND.n4835 GND.n2729 585
R2247 GND.n4837 GND.n1801 585
R2248 GND.n6053 GND.n1801 585
R2249 GND.n4838 GND.n2738 585
R2250 GND.n2738 GND.n1800 585
R2251 GND.n4840 GND.n4839 585
R2252 GND.n4845 GND.n4840 585
R2253 GND.n4822 GND.n2737 585
R2254 GND.n2737 GND.n1792 585
R2255 GND.n4821 GND.n1791 585
R2256 GND.n6061 GND.n1791 585
R2257 GND.n4820 GND.n4819 585
R2258 GND.n4819 GND.n4818 585
R2259 GND.n4816 GND.n1783 585
R2260 GND.n6067 GND.n1783 585
R2261 GND.n4815 GND.n4814 585
R2262 GND.n4814 GND.n1782 585
R2263 GND.n4813 GND.n2739 585
R2264 GND.n4813 GND.n4812 585
R2265 GND.n4744 GND.n2740 585
R2266 GND.n2740 GND.n1774 585
R2267 GND.n4745 GND.n1773 585
R2268 GND.n6075 GND.n1773 585
R2269 GND.n4749 GND.n4748 585
R2270 GND.n4748 GND.n4747 585
R2271 GND.n4750 GND.n1765 585
R2272 GND.n6081 GND.n1765 585
R2273 GND.n4752 GND.n4751 585
R2274 GND.n4753 GND.n4752 585
R2275 GND.n4743 GND.n2756 585
R2276 GND.n4755 GND.n2756 585
R2277 GND.n4742 GND.n4741 585
R2278 GND.n4741 GND.n1750 585
R2279 GND.n4740 GND.n4739 585
R2280 GND.n4740 GND.n1748 585
R2281 GND.n4738 GND.n2751 585
R2282 GND.n4762 GND.n2751 585
R2283 GND.n4737 GND.n4736 585
R2284 GND.n4736 GND.n4735 585
R2285 GND.n4734 GND.n1729 585
R2286 GND.n6096 GND.n1729 585
R2287 GND.n4733 GND.n4732 585
R2288 GND.n4732 GND.n4731 585
R2289 GND.n4730 GND.n1721 585
R2290 GND.n6102 GND.n1721 585
R2291 GND.n4729 GND.n4728 585
R2292 GND.n4728 GND.n4727 585
R2293 GND.n4724 GND.n4723 585
R2294 GND.n4725 GND.n4724 585
R2295 GND.n4722 GND.n1706 585
R2296 GND.n6109 GND.n1706 585
R2297 GND.n4721 GND.n4720 585
R2298 GND.n4720 GND.n4719 585
R2299 GND.n4718 GND.n1698 585
R2300 GND.n6115 GND.n1698 585
R2301 GND.n4717 GND.n4716 585
R2302 GND.n4716 GND.n4715 585
R2303 GND.n2758 GND.n2757 585
R2304 GND.n2760 GND.n2758 585
R2305 GND.n4678 GND.n4677 585
R2306 GND.n4677 GND.n1682 585
R2307 GND.n4679 GND.n2768 585
R2308 GND.n2768 GND.n1680 585
R2309 GND.n4681 GND.n4680 585
R2310 GND.n4690 GND.n4681 585
R2311 GND.n4676 GND.n2767 585
R2312 GND.n2767 GND.n2766 585
R2313 GND.n4675 GND.n1670 585
R2314 GND.n6130 GND.n1670 585
R2315 GND.n4674 GND.n4673 585
R2316 GND.n4673 GND.n4672 585
R2317 GND.n4670 GND.n1663 585
R2318 GND.n6136 GND.n1663 585
R2319 GND.n4669 GND.n4668 585
R2320 GND.n4668 GND.n4667 585
R2321 GND.n2770 GND.n2769 585
R2322 GND.n2771 GND.n2770 585
R2323 GND.n4649 GND.n1650 585
R2324 GND.n6144 GND.n1650 585
R2325 GND.n4651 GND.n4650 585
R2326 GND.n4652 GND.n4651 585
R2327 GND.n4148 GND.n1513 585
R2328 GND.n4154 GND.n1513 585
R2329 GND.n4150 GND.n4149 585
R2330 GND.n4151 GND.n4150 585
R2331 GND.n3295 GND.n3294 585
R2332 GND.n4135 GND.n3294 585
R2333 GND.n4144 GND.n4143 585
R2334 GND.n4143 GND.n4142 585
R2335 GND.n3298 GND.n3297 585
R2336 GND.n4132 GND.n3298 585
R2337 GND.n4094 GND.n3321 585
R2338 GND.n3321 GND.n3309 585
R2339 GND.n4096 GND.n4095 585
R2340 GND.n4097 GND.n4096 585
R2341 GND.n3322 GND.n3320 585
R2342 GND.n3320 GND.n3316 585
R2343 GND.n4089 GND.n4088 585
R2344 GND.n4088 GND.n4087 585
R2345 GND.n3325 GND.n3324 585
R2346 GND.n4072 GND.n3325 585
R2347 GND.n4057 GND.n3351 585
R2348 GND.n3351 GND.n3338 585
R2349 GND.n4059 GND.n4058 585
R2350 GND.n4060 GND.n4059 585
R2351 GND.n3352 GND.n3350 585
R2352 GND.n3350 GND.n3346 585
R2353 GND.n4052 GND.n4051 585
R2354 GND.n4051 GND.n4050 585
R2355 GND.n3355 GND.n3354 585
R2356 GND.n4035 GND.n3355 585
R2357 GND.n4020 GND.n3380 585
R2358 GND.n3380 GND.n3367 585
R2359 GND.n4022 GND.n4021 585
R2360 GND.n4023 GND.n4022 585
R2361 GND.n3381 GND.n3379 585
R2362 GND.n3379 GND.n3374 585
R2363 GND.n4015 GND.n4014 585
R2364 GND.n4014 GND.n4013 585
R2365 GND.n3384 GND.n3383 585
R2366 GND.n3998 GND.n3384 585
R2367 GND.n3964 GND.n3930 585
R2368 GND.n3930 GND.n3929 585
R2369 GND.n3967 GND.n3966 585
R2370 GND.n3968 GND.n3967 585
R2371 GND.n3963 GND.n3923 585
R2372 GND.n3956 GND.n3923 585
R2373 GND.n3961 GND.n3960 585
R2374 GND.n3960 GND.n3959 585
R2375 GND.n3933 GND.n3932 585
R2376 GND.n3954 GND.n3933 585
R2377 GND.n3416 GND.n3415 585
R2378 GND.n3937 GND.n3416 585
R2379 GND.n3983 GND.n3982 585
R2380 GND.n3982 GND.n3981 585
R2381 GND.n3984 GND.n3413 585
R2382 GND.n3909 GND.n3413 585
R2383 GND.n3987 GND.n3986 585
R2384 GND.n3988 GND.n3987 585
R2385 GND.n3414 GND.n3412 585
R2386 GND.n3412 GND.n3407 585
R2387 GND.n3901 GND.n3900 585
R2388 GND.n3902 GND.n3901 585
R2389 GND.n3435 GND.n3434 585
R2390 GND.n3884 GND.n3434 585
R2391 GND.n3895 GND.n3894 585
R2392 GND.n3894 GND.n3893 585
R2393 GND.n3438 GND.n3437 585
R2394 GND.n3881 GND.n3438 585
R2395 GND.n3860 GND.n3463 585
R2396 GND.n3463 GND.n3450 585
R2397 GND.n3862 GND.n3861 585
R2398 GND.n3863 GND.n3862 585
R2399 GND.n3464 GND.n3462 585
R2400 GND.n3462 GND.n3458 585
R2401 GND.n3855 GND.n3854 585
R2402 GND.n3854 GND.n3853 585
R2403 GND.n3467 GND.n3466 585
R2404 GND.n3838 GND.n3467 585
R2405 GND.n3823 GND.n3492 585
R2406 GND.n3492 GND.n3479 585
R2407 GND.n3825 GND.n3824 585
R2408 GND.n3826 GND.n3825 585
R2409 GND.n3493 GND.n3491 585
R2410 GND.n3491 GND.n3486 585
R2411 GND.n3818 GND.n3817 585
R2412 GND.n3817 GND.n3816 585
R2413 GND.n3496 GND.n3495 585
R2414 GND.n3801 GND.n3496 585
R2415 GND.n3786 GND.n3521 585
R2416 GND.n3521 GND.n3509 585
R2417 GND.n3788 GND.n3787 585
R2418 GND.n3789 GND.n3788 585
R2419 GND.n3522 GND.n3520 585
R2420 GND.n3520 GND.n3516 585
R2421 GND.n3781 GND.n3780 585
R2422 GND.n3780 GND.n3779 585
R2423 GND.n3576 GND.n3524 585
R2424 GND.n3579 GND.n3578 585
R2425 GND.n3577 GND.n3575 585
R2426 GND.n3584 GND.n3583 585
R2427 GND.n3586 GND.n3585 585
R2428 GND.n3589 GND.n3588 585
R2429 GND.n3587 GND.n3573 585
R2430 GND.n3594 GND.n3593 585
R2431 GND.n3596 GND.n3595 585
R2432 GND.n3599 GND.n3598 585
R2433 GND.n3597 GND.n3571 585
R2434 GND.n3604 GND.n3603 585
R2435 GND.n3606 GND.n3605 585
R2436 GND.n3609 GND.n3608 585
R2437 GND.n3607 GND.n3569 585
R2438 GND.n3614 GND.n3613 585
R2439 GND.n3618 GND.n3615 585
R2440 GND.n3621 GND.n3620 585
R2441 GND.n3619 GND.n3567 585
R2442 GND.n3626 GND.n3625 585
R2443 GND.n3628 GND.n3627 585
R2444 GND.n3631 GND.n3630 585
R2445 GND.n3629 GND.n3565 585
R2446 GND.n3636 GND.n3635 585
R2447 GND.n3638 GND.n3637 585
R2448 GND.n3641 GND.n3640 585
R2449 GND.n3639 GND.n3563 585
R2450 GND.n3646 GND.n3645 585
R2451 GND.n3648 GND.n3647 585
R2452 GND.n3651 GND.n3650 585
R2453 GND.n3649 GND.n3561 585
R2454 GND.n3656 GND.n3655 585
R2455 GND.n3658 GND.n3657 585
R2456 GND.n3661 GND.n3660 585
R2457 GND.n3659 GND.n3559 585
R2458 GND.n3668 GND.n3667 585
R2459 GND.n3670 GND.n3669 585
R2460 GND.n3673 GND.n3672 585
R2461 GND.n3671 GND.n3557 585
R2462 GND.n3678 GND.n3677 585
R2463 GND.n3680 GND.n3679 585
R2464 GND.n3683 GND.n3682 585
R2465 GND.n3681 GND.n3555 585
R2466 GND.n3688 GND.n3687 585
R2467 GND.n3690 GND.n3689 585
R2468 GND.n3693 GND.n3692 585
R2469 GND.n3691 GND.n3553 585
R2470 GND.n3698 GND.n3697 585
R2471 GND.n3700 GND.n3699 585
R2472 GND.n3703 GND.n3702 585
R2473 GND.n3701 GND.n3551 585
R2474 GND.n3708 GND.n3707 585
R2475 GND.n3710 GND.n3709 585
R2476 GND.n3716 GND.n3715 585
R2477 GND.n3714 GND.n3549 585
R2478 GND.n3721 GND.n3720 585
R2479 GND.n3723 GND.n3722 585
R2480 GND.n3726 GND.n3725 585
R2481 GND.n3724 GND.n3547 585
R2482 GND.n3731 GND.n3730 585
R2483 GND.n3733 GND.n3732 585
R2484 GND.n3736 GND.n3735 585
R2485 GND.n3734 GND.n3545 585
R2486 GND.n3741 GND.n3740 585
R2487 GND.n3743 GND.n3742 585
R2488 GND.n3746 GND.n3745 585
R2489 GND.n3744 GND.n3543 585
R2490 GND.n3751 GND.n3750 585
R2491 GND.n3753 GND.n3752 585
R2492 GND.n3756 GND.n3755 585
R2493 GND.n3754 GND.n3540 585
R2494 GND.n3760 GND.n3541 585
R2495 GND.n3761 GND.n3537 585
R2496 GND.n3762 GND.n3533 585
R2497 GND.n3288 GND.n3287 585
R2498 GND.n3286 GND.n3285 585
R2499 GND.n3284 GND.n3173 585
R2500 GND.n3280 GND.n3279 585
R2501 GND.n3278 GND.n3277 585
R2502 GND.n3276 GND.n3179 585
R2503 GND.n3178 GND.n3177 585
R2504 GND.n3272 GND.n3271 585
R2505 GND.n3270 GND.n3269 585
R2506 GND.n3268 GND.n3183 585
R2507 GND.n3182 GND.n3181 585
R2508 GND.n3264 GND.n3263 585
R2509 GND.n3262 GND.n3261 585
R2510 GND.n3260 GND.n3187 585
R2511 GND.n3186 GND.n3185 585
R2512 GND.n3256 GND.n3255 585
R2513 GND.n3254 GND.n3253 585
R2514 GND.n3252 GND.n3191 585
R2515 GND.n3190 GND.n3189 585
R2516 GND.n3248 GND.n3247 585
R2517 GND.n3246 GND.n3245 585
R2518 GND.n3244 GND.n3198 585
R2519 GND.n3197 GND.n3196 585
R2520 GND.n3240 GND.n3239 585
R2521 GND.n3238 GND.n3237 585
R2522 GND.n3236 GND.n3202 585
R2523 GND.n3201 GND.n3200 585
R2524 GND.n3232 GND.n3231 585
R2525 GND.n3230 GND.n3229 585
R2526 GND.n3228 GND.n3206 585
R2527 GND.n3205 GND.n3204 585
R2528 GND.n3224 GND.n3223 585
R2529 GND.n3222 GND.n3221 585
R2530 GND.n3220 GND.n3210 585
R2531 GND.n3209 GND.n3208 585
R2532 GND.n3216 GND.n3215 585
R2533 GND.n3214 GND.n3213 585
R2534 GND.n1568 GND.n1567 585
R2535 GND.n6273 GND.n1466 585
R2536 GND.n6222 GND.n6221 585
R2537 GND.n6223 GND.n1565 585
R2538 GND.n6224 GND.n1564 585
R2539 GND.n1563 GND.n1561 585
R2540 GND.n6228 GND.n1560 585
R2541 GND.n6229 GND.n1559 585
R2542 GND.n6230 GND.n1558 585
R2543 GND.n1557 GND.n1555 585
R2544 GND.n6234 GND.n1554 585
R2545 GND.n6235 GND.n1553 585
R2546 GND.n6236 GND.n1552 585
R2547 GND.n1551 GND.n1549 585
R2548 GND.n6240 GND.n1548 585
R2549 GND.n6241 GND.n1547 585
R2550 GND.n6242 GND.n1546 585
R2551 GND.n1545 GND.n1543 585
R2552 GND.n6246 GND.n1542 585
R2553 GND.n6247 GND.n1541 585
R2554 GND.n6248 GND.n1537 585
R2555 GND.n6249 GND.n1536 585
R2556 GND.n1534 GND.n1533 585
R2557 GND.n6253 GND.n1532 585
R2558 GND.n6254 GND.n1531 585
R2559 GND.n6255 GND.n1530 585
R2560 GND.n1528 GND.n1527 585
R2561 GND.n6259 GND.n1526 585
R2562 GND.n6260 GND.n1525 585
R2563 GND.n6261 GND.n1524 585
R2564 GND.n1522 GND.n1521 585
R2565 GND.n6265 GND.n1520 585
R2566 GND.n6266 GND.n1519 585
R2567 GND.n6267 GND.n1518 585
R2568 GND.n1515 GND.n1514 585
R2569 GND.n6272 GND.n6271 585
R2570 GND.n6273 GND.n6272 585
R2571 GND.n4156 GND.n4155 585
R2572 GND.n4155 GND.n4154 585
R2573 GND.n3172 GND.n3171 585
R2574 GND.n4151 GND.n3172 585
R2575 GND.n4137 GND.n4136 585
R2576 GND.n4136 GND.n4135 585
R2577 GND.n4138 GND.n3300 585
R2578 GND.n4142 GND.n3300 585
R2579 GND.n4134 GND.n4133 585
R2580 GND.n4133 GND.n4132 585
R2581 GND.n3308 GND.n3307 585
R2582 GND.n3309 GND.n3308 585
R2583 GND.n4081 GND.n3317 585
R2584 GND.n4097 GND.n3317 585
R2585 GND.n4082 GND.n4075 585
R2586 GND.n4075 GND.n3316 585
R2587 GND.n4083 GND.n3327 585
R2588 GND.n4087 GND.n3327 585
R2589 GND.n4074 GND.n4073 585
R2590 GND.n4073 GND.n4072 585
R2591 GND.n3337 GND.n3336 585
R2592 GND.n3338 GND.n3337 585
R2593 GND.n4044 GND.n3347 585
R2594 GND.n4060 GND.n3347 585
R2595 GND.n4045 GND.n4038 585
R2596 GND.n4038 GND.n3346 585
R2597 GND.n4046 GND.n3357 585
R2598 GND.n4050 GND.n3357 585
R2599 GND.n4037 GND.n4036 585
R2600 GND.n4036 GND.n4035 585
R2601 GND.n3366 GND.n3365 585
R2602 GND.n3367 GND.n3366 585
R2603 GND.n4007 GND.n3375 585
R2604 GND.n4023 GND.n3375 585
R2605 GND.n4008 GND.n4001 585
R2606 GND.n4001 GND.n3374 585
R2607 GND.n4009 GND.n3385 585
R2608 GND.n4013 GND.n3385 585
R2609 GND.n4000 GND.n3999 585
R2610 GND.n3999 GND.n3998 585
R2611 GND.n3394 GND.n3393 585
R2612 GND.n3929 GND.n3394 585
R2613 GND.n3970 GND.n3969 585
R2614 GND.n3969 GND.n3968 585
R2615 GND.n3971 GND.n3919 585
R2616 GND.n3956 GND.n3919 585
R2617 GND.n3935 GND.n3914 585
R2618 GND.n3959 GND.n3935 585
R2619 GND.n3975 GND.n3913 585
R2620 GND.n3954 GND.n3913 585
R2621 GND.n3976 GND.n3912 585
R2622 GND.n3937 GND.n3912 585
R2623 GND.n3977 GND.n3418 585
R2624 GND.n3981 GND.n3418 585
R2625 GND.n3911 GND.n3910 585
R2626 GND.n3910 GND.n3909 585
R2627 GND.n3908 GND.n3408 585
R2628 GND.n3988 GND.n3408 585
R2629 GND.n3431 GND.n3426 585
R2630 GND.n3431 GND.n3407 585
R2631 GND.n3887 GND.n3432 585
R2632 GND.n3902 GND.n3432 585
R2633 GND.n3888 GND.n3885 585
R2634 GND.n3885 GND.n3884 585
R2635 GND.n3889 GND.n3440 585
R2636 GND.n3893 GND.n3440 585
R2637 GND.n3883 GND.n3882 585
R2638 GND.n3882 GND.n3881 585
R2639 GND.n3449 GND.n3448 585
R2640 GND.n3450 GND.n3449 585
R2641 GND.n3847 GND.n3459 585
R2642 GND.n3863 GND.n3459 585
R2643 GND.n3848 GND.n3841 585
R2644 GND.n3841 GND.n3458 585
R2645 GND.n3849 GND.n3469 585
R2646 GND.n3853 GND.n3469 585
R2647 GND.n3840 GND.n3839 585
R2648 GND.n3839 GND.n3838 585
R2649 GND.n3478 GND.n3477 585
R2650 GND.n3479 GND.n3478 585
R2651 GND.n3810 GND.n3487 585
R2652 GND.n3826 GND.n3487 585
R2653 GND.n3811 GND.n3804 585
R2654 GND.n3804 GND.n3486 585
R2655 GND.n3812 GND.n3498 585
R2656 GND.n3816 GND.n3498 585
R2657 GND.n3803 GND.n3802 585
R2658 GND.n3802 GND.n3801 585
R2659 GND.n3507 GND.n3506 585
R2660 GND.n3509 GND.n3507 585
R2661 GND.n3772 GND.n3517 585
R2662 GND.n3789 GND.n3517 585
R2663 GND.n3535 GND.n3534 585
R2664 GND.n3534 GND.n3516 585
R2665 GND.n3777 GND.n3776 585
R2666 GND.n3779 GND.n3777 585
R2667 GND.n8014 GND.n149 585
R2668 GND.n7875 GND.n149 585
R2669 GND.n8016 GND.n8015 585
R2670 GND.n8017 GND.n8016 585
R2671 GND.n134 GND.n133 585
R2672 GND.n5300 GND.n134 585
R2673 GND.n8025 GND.n8024 585
R2674 GND.n8024 GND.n8023 585
R2675 GND.n8026 GND.n128 585
R2676 GND.n5306 GND.n128 585
R2677 GND.n8028 GND.n8027 585
R2678 GND.n8029 GND.n8028 585
R2679 GND.n113 GND.n112 585
R2680 GND.n5312 GND.n113 585
R2681 GND.n8037 GND.n8036 585
R2682 GND.n8036 GND.n8035 585
R2683 GND.n8038 GND.n107 585
R2684 GND.n5318 GND.n107 585
R2685 GND.n8040 GND.n8039 585
R2686 GND.n8041 GND.n8040 585
R2687 GND.n92 GND.n91 585
R2688 GND.n5324 GND.n92 585
R2689 GND.n8049 GND.n8048 585
R2690 GND.n8048 GND.n8047 585
R2691 GND.n8050 GND.n86 585
R2692 GND.n5330 GND.n86 585
R2693 GND.n8052 GND.n8051 585
R2694 GND.n8053 GND.n8052 585
R2695 GND.n71 GND.n70 585
R2696 GND.n5336 GND.n71 585
R2697 GND.n8061 GND.n8060 585
R2698 GND.n8060 GND.n8059 585
R2699 GND.n8062 GND.n66 585
R2700 GND.n5342 GND.n66 585
R2701 GND.n8064 GND.n8063 585
R2702 GND.n8065 GND.n8064 585
R2703 GND.n50 GND.n48 585
R2704 GND.n5348 GND.n50 585
R2705 GND.n8073 GND.n8072 585
R2706 GND.n8072 GND.n8071 585
R2707 GND.n49 GND.n47 585
R2708 GND.n5354 GND.n49 585
R2709 GND.n5362 GND.n5361 585
R2710 GND.n5363 GND.n5362 585
R2711 GND.n39 GND.n37 585
R2712 GND.n2552 GND.n37 585
R2713 GND.n8077 GND.n8076 585
R2714 GND.n8078 GND.n8077 585
R2715 GND.n38 GND.n36 585
R2716 GND.n2545 GND.n36 585
R2717 GND.n5374 GND.n2542 585
R2718 GND.n5374 GND.n5373 585
R2719 GND.n5375 GND.n45 585
R2720 GND.n5376 GND.n5375 585
R2721 GND.n2527 GND.n2526 585
R2722 GND.n5122 GND.n2527 585
R2723 GND.n5384 GND.n5383 585
R2724 GND.n5383 GND.n5382 585
R2725 GND.n5385 GND.n2523 585
R2726 GND.n5110 GND.n2523 585
R2727 GND.n5387 GND.n5386 585
R2728 GND.n5388 GND.n5387 585
R2729 GND.n2508 GND.n2507 585
R2730 GND.n5103 GND.n2508 585
R2731 GND.n5396 GND.n5395 585
R2732 GND.n5395 GND.n5394 585
R2733 GND.n5397 GND.n2502 585
R2734 GND.n5095 GND.n2502 585
R2735 GND.n5399 GND.n5398 585
R2736 GND.n5400 GND.n5399 585
R2737 GND.n2487 GND.n2486 585
R2738 GND.n5088 GND.n2487 585
R2739 GND.n5408 GND.n5407 585
R2740 GND.n5407 GND.n5406 585
R2741 GND.n5409 GND.n2481 585
R2742 GND.n5080 GND.n2481 585
R2743 GND.n5411 GND.n5410 585
R2744 GND.n5412 GND.n5411 585
R2745 GND.n2466 GND.n2465 585
R2746 GND.n5073 GND.n2466 585
R2747 GND.n5420 GND.n5419 585
R2748 GND.n5419 GND.n5418 585
R2749 GND.n5421 GND.n2460 585
R2750 GND.n5065 GND.n2460 585
R2751 GND.n5423 GND.n5422 585
R2752 GND.n5424 GND.n5423 585
R2753 GND.n2445 GND.n2444 585
R2754 GND.n5058 GND.n2445 585
R2755 GND.n5432 GND.n5431 585
R2756 GND.n5431 GND.n5430 585
R2757 GND.n5433 GND.n2438 585
R2758 GND.n5050 GND.n2438 585
R2759 GND.n5435 GND.n5434 585
R2760 GND.n5436 GND.n5435 585
R2761 GND.n2439 GND.n2316 585
R2762 GND.n5439 GND.n2316 585
R2763 GND.n5586 GND.n5585 585
R2764 GND.n5584 GND.n2315 585
R2765 GND.n5583 GND.n2314 585
R2766 GND.n5588 GND.n2314 585
R2767 GND.n5582 GND.n5581 585
R2768 GND.n5580 GND.n5579 585
R2769 GND.n5578 GND.n5577 585
R2770 GND.n5576 GND.n5575 585
R2771 GND.n5574 GND.n5573 585
R2772 GND.n5572 GND.n5571 585
R2773 GND.n5570 GND.n5569 585
R2774 GND.n5568 GND.n5567 585
R2775 GND.n5566 GND.n5565 585
R2776 GND.n5564 GND.n5563 585
R2777 GND.n5562 GND.n5561 585
R2778 GND.n5560 GND.n5559 585
R2779 GND.n5558 GND.n5557 585
R2780 GND.n5556 GND.n2333 585
R2781 GND.n5555 GND.n5554 585
R2782 GND.n5553 GND.n5552 585
R2783 GND.n5551 GND.n5550 585
R2784 GND.n5549 GND.n5548 585
R2785 GND.n5547 GND.n5546 585
R2786 GND.n5545 GND.n5544 585
R2787 GND.n5543 GND.n5542 585
R2788 GND.n5541 GND.n5540 585
R2789 GND.n5539 GND.n5538 585
R2790 GND.n5537 GND.n5536 585
R2791 GND.n5535 GND.n5534 585
R2792 GND.n5533 GND.n5532 585
R2793 GND.n5531 GND.n5530 585
R2794 GND.n5529 GND.n5528 585
R2795 GND.n5527 GND.n5526 585
R2796 GND.n5525 GND.n5524 585
R2797 GND.n5523 GND.n5522 585
R2798 GND.n5520 GND.n5519 585
R2799 GND.n5518 GND.n5517 585
R2800 GND.n5516 GND.n5515 585
R2801 GND.n5514 GND.n5513 585
R2802 GND.n5512 GND.n5511 585
R2803 GND.n5510 GND.n5509 585
R2804 GND.n5508 GND.n5507 585
R2805 GND.n5506 GND.n5505 585
R2806 GND.n5504 GND.n5503 585
R2807 GND.n5502 GND.n5501 585
R2808 GND.n5500 GND.n5499 585
R2809 GND.n5498 GND.n5497 585
R2810 GND.n5496 GND.n5495 585
R2811 GND.n5494 GND.n5493 585
R2812 GND.n5492 GND.n5491 585
R2813 GND.n5490 GND.n5489 585
R2814 GND.n5488 GND.n5487 585
R2815 GND.n5486 GND.n5485 585
R2816 GND.n5483 GND.n5482 585
R2817 GND.n5481 GND.n5480 585
R2818 GND.n5479 GND.n5478 585
R2819 GND.n5477 GND.n5476 585
R2820 GND.n5475 GND.n5474 585
R2821 GND.n5473 GND.n5472 585
R2822 GND.n5471 GND.n5470 585
R2823 GND.n5469 GND.n5468 585
R2824 GND.n5467 GND.n5466 585
R2825 GND.n5465 GND.n5464 585
R2826 GND.n5463 GND.n5462 585
R2827 GND.n5461 GND.n5460 585
R2828 GND.n5459 GND.n5458 585
R2829 GND.n5457 GND.n5456 585
R2830 GND.n5455 GND.n5454 585
R2831 GND.n5453 GND.n5452 585
R2832 GND.n5451 GND.n5450 585
R2833 GND.n5449 GND.n5448 585
R2834 GND.n2398 GND.n2395 585
R2835 GND.n5444 GND.n2304 585
R2836 GND.n5588 GND.n2304 585
R2837 GND.n289 GND.n283 585
R2838 GND.n7882 GND.n280 585
R2839 GND.n7884 GND.n7883 585
R2840 GND.n7886 GND.n278 585
R2841 GND.n7888 GND.n7887 585
R2842 GND.n7889 GND.n273 585
R2843 GND.n7891 GND.n7890 585
R2844 GND.n7893 GND.n271 585
R2845 GND.n7895 GND.n7894 585
R2846 GND.n7896 GND.n266 585
R2847 GND.n7898 GND.n7897 585
R2848 GND.n7900 GND.n264 585
R2849 GND.n7902 GND.n7901 585
R2850 GND.n7903 GND.n259 585
R2851 GND.n7905 GND.n7904 585
R2852 GND.n7907 GND.n257 585
R2853 GND.n7909 GND.n7908 585
R2854 GND.n7910 GND.n252 585
R2855 GND.n7912 GND.n7911 585
R2856 GND.n7914 GND.n251 585
R2857 GND.n7916 GND.n7915 585
R2858 GND.n7917 GND.n242 585
R2859 GND.n7919 GND.n7918 585
R2860 GND.n7921 GND.n240 585
R2861 GND.n7923 GND.n7922 585
R2862 GND.n7924 GND.n235 585
R2863 GND.n7926 GND.n7925 585
R2864 GND.n7928 GND.n233 585
R2865 GND.n7930 GND.n7929 585
R2866 GND.n7931 GND.n228 585
R2867 GND.n7933 GND.n7932 585
R2868 GND.n7935 GND.n226 585
R2869 GND.n7937 GND.n7936 585
R2870 GND.n7938 GND.n222 585
R2871 GND.n7940 GND.n7939 585
R2872 GND.n7942 GND.n219 585
R2873 GND.n7944 GND.n7943 585
R2874 GND.n220 GND.n213 585
R2875 GND.n7948 GND.n217 585
R2876 GND.n7949 GND.n209 585
R2877 GND.n7951 GND.n7950 585
R2878 GND.n7953 GND.n207 585
R2879 GND.n7955 GND.n7954 585
R2880 GND.n7956 GND.n202 585
R2881 GND.n7958 GND.n7957 585
R2882 GND.n7960 GND.n200 585
R2883 GND.n7962 GND.n7961 585
R2884 GND.n7963 GND.n195 585
R2885 GND.n7965 GND.n7964 585
R2886 GND.n7967 GND.n193 585
R2887 GND.n7969 GND.n7968 585
R2888 GND.n7970 GND.n188 585
R2889 GND.n7972 GND.n7971 585
R2890 GND.n7974 GND.n187 585
R2891 GND.n7975 GND.n184 585
R2892 GND.n7978 GND.n7977 585
R2893 GND.n186 GND.n180 585
R2894 GND.n7982 GND.n177 585
R2895 GND.n7984 GND.n7983 585
R2896 GND.n7986 GND.n175 585
R2897 GND.n7988 GND.n7987 585
R2898 GND.n7989 GND.n170 585
R2899 GND.n7991 GND.n7990 585
R2900 GND.n7993 GND.n168 585
R2901 GND.n7995 GND.n7994 585
R2902 GND.n7996 GND.n163 585
R2903 GND.n7998 GND.n7997 585
R2904 GND.n8000 GND.n161 585
R2905 GND.n8002 GND.n8001 585
R2906 GND.n8003 GND.n156 585
R2907 GND.n8005 GND.n8004 585
R2908 GND.n8007 GND.n155 585
R2909 GND.n8008 GND.n153 585
R2910 GND.n8011 GND.n8010 585
R2911 GND.n7877 GND.n7876 585
R2912 GND.n7876 GND.n7875 585
R2913 GND.n287 GND.n146 585
R2914 GND.n8017 GND.n146 585
R2915 GND.n5299 GND.n5298 585
R2916 GND.n5300 GND.n5299 585
R2917 GND.n5225 GND.n136 585
R2918 GND.n8023 GND.n136 585
R2919 GND.n5308 GND.n5307 585
R2920 GND.n5307 GND.n5306 585
R2921 GND.n5309 GND.n125 585
R2922 GND.n8029 GND.n125 585
R2923 GND.n5311 GND.n5310 585
R2924 GND.n5312 GND.n5311 585
R2925 GND.n5218 GND.n115 585
R2926 GND.n8035 GND.n115 585
R2927 GND.n5320 GND.n5319 585
R2928 GND.n5319 GND.n5318 585
R2929 GND.n5321 GND.n104 585
R2930 GND.n8041 GND.n104 585
R2931 GND.n5323 GND.n5322 585
R2932 GND.n5324 GND.n5323 585
R2933 GND.n5211 GND.n94 585
R2934 GND.n8047 GND.n94 585
R2935 GND.n5332 GND.n5331 585
R2936 GND.n5331 GND.n5330 585
R2937 GND.n5333 GND.n83 585
R2938 GND.n8053 GND.n83 585
R2939 GND.n5335 GND.n5334 585
R2940 GND.n5336 GND.n5335 585
R2941 GND.n5204 GND.n73 585
R2942 GND.n8059 GND.n73 585
R2943 GND.n5344 GND.n5343 585
R2944 GND.n5343 GND.n5342 585
R2945 GND.n5345 GND.n63 585
R2946 GND.n8065 GND.n63 585
R2947 GND.n5347 GND.n5346 585
R2948 GND.n5348 GND.n5347 585
R2949 GND.n5136 GND.n52 585
R2950 GND.n8071 GND.n52 585
R2951 GND.n5356 GND.n5355 585
R2952 GND.n5355 GND.n5354 585
R2953 GND.n5357 GND.n2553 585
R2954 GND.n5363 GND.n2553 585
R2955 GND.n5135 GND.n5134 585
R2956 GND.n5134 GND.n2552 585
R2957 GND.n5133 GND.n33 585
R2958 GND.n8078 GND.n33 585
R2959 GND.n2561 GND.n2560 585
R2960 GND.n2560 GND.n2545 585
R2961 GND.n5126 GND.n2543 585
R2962 GND.n5373 GND.n2543 585
R2963 GND.n5125 GND.n2539 585
R2964 GND.n5376 GND.n2539 585
R2965 GND.n5124 GND.n5123 585
R2966 GND.n5123 GND.n5122 585
R2967 GND.n2562 GND.n2529 585
R2968 GND.n5382 GND.n2529 585
R2969 GND.n5109 GND.n5108 585
R2970 GND.n5110 GND.n5109 585
R2971 GND.n5106 GND.n2520 585
R2972 GND.n5388 GND.n2520 585
R2973 GND.n5105 GND.n5104 585
R2974 GND.n5104 GND.n5103 585
R2975 GND.n2566 GND.n2510 585
R2976 GND.n5394 GND.n2510 585
R2977 GND.n5094 GND.n5093 585
R2978 GND.n5095 GND.n5094 585
R2979 GND.n5091 GND.n2499 585
R2980 GND.n5400 GND.n2499 585
R2981 GND.n5090 GND.n5089 585
R2982 GND.n5089 GND.n5088 585
R2983 GND.n2570 GND.n2489 585
R2984 GND.n5406 GND.n2489 585
R2985 GND.n5079 GND.n5078 585
R2986 GND.n5080 GND.n5079 585
R2987 GND.n5076 GND.n2478 585
R2988 GND.n5412 GND.n2478 585
R2989 GND.n5075 GND.n5074 585
R2990 GND.n5074 GND.n5073 585
R2991 GND.n2574 GND.n2468 585
R2992 GND.n5418 GND.n2468 585
R2993 GND.n5064 GND.n5063 585
R2994 GND.n5065 GND.n5064 585
R2995 GND.n5061 GND.n2458 585
R2996 GND.n5424 GND.n2458 585
R2997 GND.n5060 GND.n5059 585
R2998 GND.n5059 GND.n5058 585
R2999 GND.n2658 GND.n2447 585
R3000 GND.n5430 GND.n2447 585
R3001 GND.n5049 GND.n5048 585
R3002 GND.n5050 GND.n5049 585
R3003 GND.n2403 GND.n2402 585
R3004 GND.n5436 GND.n2403 585
R3005 GND.n5441 GND.n5440 585
R3006 GND.n5440 GND.n5439 585
R3007 GND.n7753 GND.n7752 585
R3008 GND.n7754 GND.n7753 585
R3009 GND.n411 GND.n410 585
R3010 GND.n7755 GND.n411 585
R3011 GND.n7758 GND.n7757 585
R3012 GND.n7757 GND.n7756 585
R3013 GND.n7759 GND.n405 585
R3014 GND.n405 GND.n404 585
R3015 GND.n7761 GND.n7760 585
R3016 GND.n7762 GND.n7761 585
R3017 GND.n403 GND.n402 585
R3018 GND.n7763 GND.n403 585
R3019 GND.n7766 GND.n7765 585
R3020 GND.n7765 GND.n7764 585
R3021 GND.n7767 GND.n397 585
R3022 GND.n397 GND.n396 585
R3023 GND.n7769 GND.n7768 585
R3024 GND.n7770 GND.n7769 585
R3025 GND.n395 GND.n394 585
R3026 GND.n7771 GND.n395 585
R3027 GND.n7774 GND.n7773 585
R3028 GND.n7773 GND.n7772 585
R3029 GND.n7775 GND.n389 585
R3030 GND.n389 GND.n388 585
R3031 GND.n7777 GND.n7776 585
R3032 GND.n7778 GND.n7777 585
R3033 GND.n387 GND.n386 585
R3034 GND.n7779 GND.n387 585
R3035 GND.n7782 GND.n7781 585
R3036 GND.n7781 GND.n7780 585
R3037 GND.n7783 GND.n381 585
R3038 GND.n381 GND.n380 585
R3039 GND.n7785 GND.n7784 585
R3040 GND.n7786 GND.n7785 585
R3041 GND.n379 GND.n378 585
R3042 GND.n7787 GND.n379 585
R3043 GND.n7790 GND.n7789 585
R3044 GND.n7789 GND.n7788 585
R3045 GND.n7791 GND.n373 585
R3046 GND.n373 GND.n372 585
R3047 GND.n7793 GND.n7792 585
R3048 GND.n7794 GND.n7793 585
R3049 GND.n371 GND.n370 585
R3050 GND.n7795 GND.n371 585
R3051 GND.n7798 GND.n7797 585
R3052 GND.n7797 GND.n7796 585
R3053 GND.n7799 GND.n365 585
R3054 GND.n365 GND.n364 585
R3055 GND.n7801 GND.n7800 585
R3056 GND.n7802 GND.n7801 585
R3057 GND.n363 GND.n362 585
R3058 GND.n7803 GND.n363 585
R3059 GND.n7806 GND.n7805 585
R3060 GND.n7805 GND.n7804 585
R3061 GND.n7807 GND.n357 585
R3062 GND.n357 GND.n356 585
R3063 GND.n7809 GND.n7808 585
R3064 GND.n7810 GND.n7809 585
R3065 GND.n355 GND.n354 585
R3066 GND.n7811 GND.n355 585
R3067 GND.n7814 GND.n7813 585
R3068 GND.n7813 GND.n7812 585
R3069 GND.n7815 GND.n349 585
R3070 GND.n349 GND.n348 585
R3071 GND.n7817 GND.n7816 585
R3072 GND.n7818 GND.n7817 585
R3073 GND.n347 GND.n346 585
R3074 GND.n7819 GND.n347 585
R3075 GND.n7822 GND.n7821 585
R3076 GND.n7821 GND.n7820 585
R3077 GND.n7823 GND.n341 585
R3078 GND.n341 GND.n340 585
R3079 GND.n7825 GND.n7824 585
R3080 GND.n7826 GND.n7825 585
R3081 GND.n339 GND.n338 585
R3082 GND.n7827 GND.n339 585
R3083 GND.n7830 GND.n7829 585
R3084 GND.n7829 GND.n7828 585
R3085 GND.n7831 GND.n333 585
R3086 GND.n333 GND.n332 585
R3087 GND.n7833 GND.n7832 585
R3088 GND.n7834 GND.n7833 585
R3089 GND.n331 GND.n330 585
R3090 GND.n7835 GND.n331 585
R3091 GND.n7838 GND.n7837 585
R3092 GND.n7837 GND.n7836 585
R3093 GND.n7839 GND.n325 585
R3094 GND.n325 GND.n324 585
R3095 GND.n7841 GND.n7840 585
R3096 GND.n7842 GND.n7841 585
R3097 GND.n323 GND.n322 585
R3098 GND.n7843 GND.n323 585
R3099 GND.n7846 GND.n7845 585
R3100 GND.n7845 GND.n7844 585
R3101 GND.n7847 GND.n317 585
R3102 GND.n317 GND.n316 585
R3103 GND.n7849 GND.n7848 585
R3104 GND.n7850 GND.n7849 585
R3105 GND.n315 GND.n314 585
R3106 GND.n7851 GND.n315 585
R3107 GND.n7854 GND.n7853 585
R3108 GND.n7853 GND.n7852 585
R3109 GND.n7855 GND.n309 585
R3110 GND.n309 GND.n308 585
R3111 GND.n7857 GND.n7856 585
R3112 GND.n7858 GND.n7857 585
R3113 GND.n307 GND.n306 585
R3114 GND.n7859 GND.n307 585
R3115 GND.n7862 GND.n7861 585
R3116 GND.n7861 GND.n7860 585
R3117 GND.n7863 GND.n301 585
R3118 GND.n301 GND.n300 585
R3119 GND.n7865 GND.n7864 585
R3120 GND.n7866 GND.n7865 585
R3121 GND.n299 GND.n298 585
R3122 GND.n7867 GND.n299 585
R3123 GND.n7870 GND.n7869 585
R3124 GND.n7869 GND.n7868 585
R3125 GND.n7871 GND.n293 585
R3126 GND.n293 GND.n291 585
R3127 GND.n7873 GND.n7872 585
R3128 GND.n7874 GND.n7873 585
R3129 GND.n294 GND.n292 585
R3130 GND.n292 GND.n148 585
R3131 GND.n5175 GND.n5170 585
R3132 GND.n5170 GND.n145 585
R3133 GND.n5177 GND.n5176 585
R3134 GND.n5177 GND.n138 585
R3135 GND.n5178 GND.n5169 585
R3136 GND.n5178 GND.n135 585
R3137 GND.n5180 GND.n5179 585
R3138 GND.n5179 GND.n127 585
R3139 GND.n5181 GND.n5164 585
R3140 GND.n5164 GND.n124 585
R3141 GND.n5183 GND.n5182 585
R3142 GND.n5183 GND.n117 585
R3143 GND.n5184 GND.n5163 585
R3144 GND.n5184 GND.n114 585
R3145 GND.n5186 GND.n5185 585
R3146 GND.n5185 GND.n106 585
R3147 GND.n5187 GND.n5158 585
R3148 GND.n5158 GND.n103 585
R3149 GND.n5189 GND.n5188 585
R3150 GND.n5189 GND.n96 585
R3151 GND.n5190 GND.n5157 585
R3152 GND.n5190 GND.n93 585
R3153 GND.n5192 GND.n5191 585
R3154 GND.n5191 GND.n85 585
R3155 GND.n5193 GND.n5152 585
R3156 GND.n5152 GND.n82 585
R3157 GND.n5195 GND.n5194 585
R3158 GND.n5195 GND.n75 585
R3159 GND.n5196 GND.n5151 585
R3160 GND.n5196 GND.n72 585
R3161 GND.n5198 GND.n5197 585
R3162 GND.n5197 GND.n65 585
R3163 GND.n5199 GND.n5144 585
R3164 GND.n5144 GND.n62 585
R3165 GND.n5201 GND.n5200 585
R3166 GND.n5202 GND.n5201 585
R3167 GND.n5147 GND.n5143 585
R3168 GND.n5143 GND.n51 585
R3169 GND.n5145 GND.n2550 585
R3170 GND.n2555 GND.n2550 585
R3171 GND.n5365 GND.n2551 585
R3172 GND.n5365 GND.n5364 585
R3173 GND.n5367 GND.n5366 585
R3174 GND.n5366 GND.n34 585
R3175 GND.n5368 GND.n2547 585
R3176 GND.n2547 GND.n32 585
R3177 GND.n5371 GND.n5370 585
R3178 GND.n5372 GND.n5371 585
R3179 GND.n2548 GND.n2546 585
R3180 GND.n2546 GND.n2541 585
R3181 GND.n2632 GND.n2631 585
R3182 GND.n2632 GND.n2538 585
R3183 GND.n2634 GND.n2633 585
R3184 GND.n2633 GND.n2531 585
R3185 GND.n2636 GND.n2627 585
R3186 GND.n2627 GND.n2528 585
R3187 GND.n2638 GND.n2637 585
R3188 GND.n2638 GND.n2522 585
R3189 GND.n2639 GND.n2626 585
R3190 GND.n2639 GND.n2519 585
R3191 GND.n2641 GND.n2640 585
R3192 GND.n2640 GND.n2512 585
R3193 GND.n2642 GND.n2621 585
R3194 GND.n2621 GND.n2509 585
R3195 GND.n2644 GND.n2643 585
R3196 GND.n2644 GND.n2501 585
R3197 GND.n2645 GND.n2620 585
R3198 GND.n2645 GND.n2498 585
R3199 GND.n2647 GND.n2646 585
R3200 GND.n2646 GND.n2491 585
R3201 GND.n2648 GND.n2615 585
R3202 GND.n2615 GND.n2488 585
R3203 GND.n2650 GND.n2649 585
R3204 GND.n2650 GND.n2480 585
R3205 GND.n2651 GND.n2614 585
R3206 GND.n2651 GND.n2477 585
R3207 GND.n2653 GND.n2652 585
R3208 GND.n2652 GND.n2470 585
R3209 GND.n2654 GND.n2579 585
R3210 GND.n2579 GND.n2467 585
R3211 GND.n2656 GND.n2655 585
R3212 GND.n2657 GND.n2656 585
R3213 GND.n2580 GND.n2578 585
R3214 GND.n2578 GND.n2457 585
R3215 GND.n2608 GND.n2607 585
R3216 GND.n2607 GND.n2449 585
R3217 GND.n2606 GND.n2582 585
R3218 GND.n2606 GND.n2446 585
R3219 GND.n2605 GND.n2604 585
R3220 GND.n2605 GND.n2437 585
R3221 GND.n2584 GND.n2583 585
R3222 GND.n2583 GND.n2406 585
R3223 GND.n2600 GND.n2599 585
R3224 GND.n2599 GND.n2404 585
R3225 GND.n2598 GND.n2586 585
R3226 GND.n2598 GND.n2305 585
R3227 GND.n2597 GND.n2596 585
R3228 GND.n2597 GND.n2268 585
R3229 GND.n2589 GND.n2588 585
R3230 GND.n2588 GND.n2587 585
R3231 GND.n2592 GND.n2591 585
R3232 GND.n2591 GND.n2219 585
R3233 GND.n2216 GND.n2215 585
R3234 GND.n5644 GND.n2216 585
R3235 GND.n5647 GND.n5646 585
R3236 GND.n5646 GND.n5645 585
R3237 GND.n5648 GND.n2208 585
R3238 GND.n2217 GND.n2208 585
R3239 GND.n5650 GND.n5649 585
R3240 GND.n5651 GND.n5650 585
R3241 GND.n2209 GND.n2207 585
R3242 GND.n2207 GND.n2204 585
R3243 GND.n2189 GND.n2188 585
R3244 GND.n2193 GND.n2189 585
R3245 GND.n5661 GND.n5660 585
R3246 GND.n5660 GND.n5659 585
R3247 GND.n5662 GND.n2181 585
R3248 GND.n2190 GND.n2181 585
R3249 GND.n5664 GND.n5663 585
R3250 GND.n5665 GND.n5664 585
R3251 GND.n2182 GND.n2180 585
R3252 GND.n5002 GND.n2180 585
R3253 GND.n2163 GND.n2162 585
R3254 GND.n2167 GND.n2163 585
R3255 GND.n5675 GND.n5674 585
R3256 GND.n5674 GND.n5673 585
R3257 GND.n5676 GND.n2155 585
R3258 GND.n2164 GND.n2155 585
R3259 GND.n5678 GND.n5677 585
R3260 GND.n5679 GND.n5678 585
R3261 GND.n2156 GND.n2154 585
R3262 GND.n2154 GND.n2151 585
R3263 GND.n2136 GND.n2135 585
R3264 GND.n2140 GND.n2136 585
R3265 GND.n5689 GND.n5688 585
R3266 GND.n5688 GND.n5687 585
R3267 GND.n5690 GND.n2128 585
R3268 GND.n2137 GND.n2128 585
R3269 GND.n5692 GND.n5691 585
R3270 GND.n5693 GND.n5692 585
R3271 GND.n2129 GND.n2127 585
R3272 GND.n2127 GND.n2124 585
R3273 GND.n2109 GND.n2108 585
R3274 GND.n2113 GND.n2109 585
R3275 GND.n5703 GND.n5702 585
R3276 GND.n5702 GND.n5701 585
R3277 GND.n5704 GND.n2101 585
R3278 GND.n2110 GND.n2101 585
R3279 GND.n5706 GND.n5705 585
R3280 GND.n5707 GND.n5706 585
R3281 GND.n2102 GND.n2100 585
R3282 GND.n2100 GND.n2097 585
R3283 GND.n2082 GND.n2081 585
R3284 GND.n2086 GND.n2082 585
R3285 GND.n5717 GND.n5716 585
R3286 GND.n5716 GND.n5715 585
R3287 GND.n5718 GND.n2074 585
R3288 GND.n2083 GND.n2074 585
R3289 GND.n5720 GND.n5719 585
R3290 GND.n5721 GND.n5720 585
R3291 GND.n2075 GND.n2073 585
R3292 GND.n2073 GND.n2070 585
R3293 GND.n2055 GND.n2054 585
R3294 GND.n2059 GND.n2055 585
R3295 GND.n5731 GND.n5730 585
R3296 GND.n5730 GND.n5729 585
R3297 GND.n5732 GND.n2047 585
R3298 GND.n2056 GND.n2047 585
R3299 GND.n5734 GND.n5733 585
R3300 GND.n5735 GND.n5734 585
R3301 GND.n2048 GND.n2046 585
R3302 GND.n2046 GND.n2043 585
R3303 GND.n2028 GND.n2027 585
R3304 GND.n2032 GND.n2028 585
R3305 GND.n5745 GND.n5744 585
R3306 GND.n5744 GND.n5743 585
R3307 GND.n5746 GND.n2020 585
R3308 GND.n2029 GND.n2020 585
R3309 GND.n5748 GND.n5747 585
R3310 GND.n5749 GND.n5748 585
R3311 GND.n2021 GND.n2019 585
R3312 GND.n2019 GND.n2016 585
R3313 GND.n2002 GND.n2001 585
R3314 GND.n2691 GND.n2002 585
R3315 GND.n5759 GND.n5758 585
R3316 GND.n5758 GND.n5757 585
R3317 GND.n5760 GND.n1994 585
R3318 GND.n2003 GND.n1994 585
R3319 GND.n5762 GND.n5761 585
R3320 GND.n5763 GND.n5762 585
R3321 GND.n1995 GND.n1993 585
R3322 GND.n1993 GND.n1990 585
R3323 GND.n1975 GND.n1974 585
R3324 GND.n1979 GND.n1975 585
R3325 GND.n5773 GND.n5772 585
R3326 GND.n5772 GND.n5771 585
R3327 GND.n5774 GND.n1967 585
R3328 GND.n1976 GND.n1967 585
R3329 GND.n5776 GND.n5775 585
R3330 GND.n5777 GND.n5776 585
R3331 GND.n1968 GND.n1966 585
R3332 GND.n1966 GND.n1963 585
R3333 GND.n1948 GND.n1947 585
R3334 GND.n1952 GND.n1948 585
R3335 GND.n5787 GND.n5786 585
R3336 GND.n5786 GND.n5785 585
R3337 GND.n5788 GND.n1940 585
R3338 GND.n1949 GND.n1940 585
R3339 GND.n5790 GND.n5789 585
R3340 GND.n5791 GND.n5790 585
R3341 GND.n1941 GND.n1939 585
R3342 GND.n1939 GND.n1936 585
R3343 GND.n1921 GND.n1920 585
R3344 GND.n1925 GND.n1921 585
R3345 GND.n5801 GND.n5800 585
R3346 GND.n5800 GND.n5799 585
R3347 GND.n5802 GND.n1915 585
R3348 GND.n1922 GND.n1915 585
R3349 GND.n5804 GND.n5803 585
R3350 GND.n5805 GND.n5804 585
R3351 GND.n1851 GND.n1850 585
R3352 GND.n1912 GND.n1851 585
R3353 GND.n6014 GND.n6013 585
R3354 GND.n6013 GND.n6012 585
R3355 GND.n6015 GND.n1845 585
R3356 GND.n5834 GND.n1845 585
R3357 GND.n6017 GND.n6016 585
R3358 GND.n6018 GND.n6017 585
R3359 GND.n1833 GND.n1832 585
R3360 GND.n5826 GND.n1833 585
R3361 GND.n6028 GND.n6027 585
R3362 GND.n6027 GND.n6026 585
R3363 GND.n6029 GND.n1827 585
R3364 GND.n1896 GND.n1827 585
R3365 GND.n6031 GND.n6030 585
R3366 GND.n6032 GND.n6031 585
R3367 GND.n1816 GND.n1815 585
R3368 GND.n2712 GND.n1816 585
R3369 GND.n6042 GND.n6041 585
R3370 GND.n6041 GND.n6040 585
R3371 GND.n6043 GND.n1810 585
R3372 GND.n2722 GND.n1810 585
R3373 GND.n6045 GND.n6044 585
R3374 GND.n6046 GND.n6045 585
R3375 GND.n1799 GND.n1798 585
R3376 GND.n2729 GND.n1799 585
R3377 GND.n6056 GND.n6055 585
R3378 GND.n6055 GND.n6054 585
R3379 GND.n6057 GND.n1793 585
R3380 GND.n4842 GND.n1793 585
R3381 GND.n6059 GND.n6058 585
R3382 GND.n6060 GND.n6059 585
R3383 GND.n1781 GND.n1780 585
R3384 GND.n4817 GND.n1781 585
R3385 GND.n6070 GND.n6069 585
R3386 GND.n6069 GND.n6068 585
R3387 GND.n6071 GND.n1775 585
R3388 GND.n4809 GND.n1775 585
R3389 GND.n6073 GND.n6072 585
R3390 GND.n6074 GND.n6073 585
R3391 GND.n1763 GND.n1762 585
R3392 GND.n4746 GND.n1763 585
R3393 GND.n6084 GND.n6083 585
R3394 GND.n6083 GND.n6082 585
R3395 GND.n6085 GND.n1752 585
R3396 GND.n4754 GND.n1752 585
R3397 GND.n6087 GND.n6086 585
R3398 GND.n6088 GND.n6087 585
R3399 GND.n1753 GND.n1751 585
R3400 GND.n2752 GND.n1751 585
R3401 GND.n1756 GND.n1755 585
R3402 GND.n1755 GND.n1731 585
R3403 GND.n1719 GND.n1718 585
R3404 GND.n1728 GND.n1719 585
R3405 GND.n6105 GND.n6104 585
R3406 GND.n6104 GND.n6103 585
R3407 GND.n6106 GND.n1708 585
R3408 GND.n4726 GND.n1708 585
R3409 GND.n6108 GND.n6107 585
R3410 GND.n6109 GND.n6108 585
R3411 GND.n1709 GND.n1707 585
R3412 GND.n1707 GND.n1699 585
R3413 GND.n1712 GND.n1711 585
R3414 GND.n1711 GND.n1696 585
R3415 GND.n1679 GND.n1678 585
R3416 GND.n2759 GND.n1679 585
R3417 GND.n6125 GND.n6124 585
R3418 GND.n6124 GND.n6123 585
R3419 GND.n6126 GND.n1673 585
R3420 GND.n2765 GND.n1673 585
R3421 GND.n6128 GND.n6127 585
R3422 GND.n6129 GND.n6128 585
R3423 GND.n1674 GND.n1672 585
R3424 GND.n4671 GND.n1672 585
R3425 GND.n4555 GND.n4554 585
R3426 GND.n4554 GND.n1661 585
R3427 GND.n4556 GND.n4548 585
R3428 GND.n4548 GND.n1652 585
R3429 GND.n4558 GND.n4557 585
R3430 GND.n4558 GND.n1649 585
R3431 GND.n4559 GND.n4547 585
R3432 GND.n4559 GND.n1613 585
R3433 GND.n4561 GND.n4560 585
R3434 GND.n4560 GND.n2778 585
R3435 GND.n4562 GND.n2789 585
R3436 GND.n2789 GND.n2777 585
R3437 GND.n4564 GND.n4563 585
R3438 GND.n4565 GND.n4564 585
R3439 GND.n2790 GND.n2788 585
R3440 GND.n2788 GND.n2785 585
R3441 GND.n4541 GND.n4540 585
R3442 GND.n4540 GND.n4539 585
R3443 GND.n2793 GND.n2792 585
R3444 GND.n2801 GND.n2793 585
R3445 GND.n4511 GND.n2812 585
R3446 GND.n2812 GND.n2800 585
R3447 GND.n4513 GND.n4512 585
R3448 GND.n4514 GND.n4513 585
R3449 GND.n2813 GND.n2811 585
R3450 GND.n2811 GND.n2808 585
R3451 GND.n4506 GND.n4505 585
R3452 GND.n4505 GND.n4504 585
R3453 GND.n2816 GND.n2815 585
R3454 GND.n2824 GND.n2816 585
R3455 GND.n4479 GND.n2835 585
R3456 GND.n2835 GND.n2823 585
R3457 GND.n4481 GND.n4480 585
R3458 GND.n4482 GND.n4481 585
R3459 GND.n2836 GND.n2834 585
R3460 GND.n2834 GND.n2831 585
R3461 GND.n4474 GND.n4473 585
R3462 GND.n4473 GND.n4472 585
R3463 GND.n2839 GND.n2838 585
R3464 GND.n2847 GND.n2839 585
R3465 GND.n4447 GND.n2858 585
R3466 GND.n2858 GND.n2846 585
R3467 GND.n4449 GND.n4448 585
R3468 GND.n4450 GND.n4449 585
R3469 GND.n2859 GND.n2857 585
R3470 GND.n2857 GND.n2854 585
R3471 GND.n4442 GND.n4441 585
R3472 GND.n4441 GND.n4440 585
R3473 GND.n2862 GND.n2861 585
R3474 GND.n2870 GND.n2862 585
R3475 GND.n4415 GND.n2881 585
R3476 GND.n2881 GND.n2869 585
R3477 GND.n4417 GND.n4416 585
R3478 GND.n4418 GND.n4417 585
R3479 GND.n2882 GND.n2880 585
R3480 GND.n2880 GND.n2877 585
R3481 GND.n4410 GND.n4409 585
R3482 GND.n4409 GND.n4408 585
R3483 GND.n2885 GND.n2884 585
R3484 GND.n2893 GND.n2885 585
R3485 GND.n4383 GND.n2904 585
R3486 GND.n2904 GND.n2892 585
R3487 GND.n4385 GND.n4384 585
R3488 GND.n4386 GND.n4385 585
R3489 GND.n2905 GND.n2903 585
R3490 GND.n2903 GND.n2900 585
R3491 GND.n4378 GND.n4377 585
R3492 GND.n4377 GND.n4376 585
R3493 GND.n2908 GND.n2907 585
R3494 GND.n2916 GND.n2908 585
R3495 GND.n4351 GND.n2927 585
R3496 GND.n2927 GND.n2915 585
R3497 GND.n4353 GND.n4352 585
R3498 GND.n4354 GND.n4353 585
R3499 GND.n2928 GND.n2926 585
R3500 GND.n2926 GND.n2923 585
R3501 GND.n4346 GND.n4345 585
R3502 GND.n4345 GND.n4344 585
R3503 GND.n2931 GND.n2930 585
R3504 GND.n2938 GND.n2931 585
R3505 GND.n4319 GND.n2950 585
R3506 GND.n2950 GND.n2937 585
R3507 GND.n4321 GND.n4320 585
R3508 GND.n4322 GND.n4321 585
R3509 GND.n2951 GND.n2949 585
R3510 GND.n2949 GND.n2946 585
R3511 GND.n4314 GND.n4313 585
R3512 GND.n4313 GND.n4312 585
R3513 GND.n2954 GND.n2953 585
R3514 GND.n2962 GND.n2954 585
R3515 GND.n4287 GND.n2973 585
R3516 GND.n2973 GND.n2961 585
R3517 GND.n4289 GND.n4288 585
R3518 GND.n4290 GND.n4289 585
R3519 GND.n2974 GND.n2972 585
R3520 GND.n2972 GND.n2969 585
R3521 GND.n4282 GND.n4281 585
R3522 GND.n4281 GND.n4280 585
R3523 GND.n2977 GND.n2976 585
R3524 GND.n2985 GND.n2977 585
R3525 GND.n4255 GND.n2996 585
R3526 GND.n2996 GND.n2984 585
R3527 GND.n4257 GND.n4256 585
R3528 GND.n4258 GND.n4257 585
R3529 GND.n2997 GND.n2995 585
R3530 GND.n2995 GND.n2992 585
R3531 GND.n4250 GND.n4249 585
R3532 GND.n4249 GND.n4248 585
R3533 GND.n3000 GND.n2999 585
R3534 GND.n3008 GND.n3000 585
R3535 GND.n4223 GND.n3019 585
R3536 GND.n3019 GND.n3007 585
R3537 GND.n4225 GND.n4224 585
R3538 GND.n4226 GND.n4225 585
R3539 GND.n3020 GND.n3018 585
R3540 GND.n3018 GND.n3015 585
R3541 GND.n4218 GND.n4217 585
R3542 GND.n4217 GND.n4216 585
R3543 GND.n3023 GND.n3022 585
R3544 GND.n3031 GND.n3023 585
R3545 GND.n4191 GND.n3041 585
R3546 GND.n3041 GND.n3030 585
R3547 GND.n4193 GND.n4192 585
R3548 GND.n4194 GND.n4193 585
R3549 GND.n3042 GND.n3040 585
R3550 GND.n3040 GND.n3037 585
R3551 GND.n4186 GND.n4185 585
R3552 GND.n4185 GND.n4184 585
R3553 GND.n3045 GND.n3044 585
R3554 GND.n3046 GND.n3045 585
R3555 GND.n4117 GND.n4115 585
R3556 GND.n4117 GND.n4116 585
R3557 GND.n4118 GND.n4112 585
R3558 GND.n4118 GND.n1494 585
R3559 GND.n4120 GND.n4119 585
R3560 GND.n4119 GND.n1465 585
R3561 GND.n4121 GND.n4107 585
R3562 GND.n4107 GND.n3290 585
R3563 GND.n4123 GND.n4122 585
R3564 GND.n4123 GND.n3289 585
R3565 GND.n4124 GND.n4106 585
R3566 GND.n4124 GND.n3293 585
R3567 GND.n4126 GND.n4125 585
R3568 GND.n4125 GND.n3301 585
R3569 GND.n4127 GND.n3311 585
R3570 GND.n3311 GND.n3299 585
R3571 GND.n4129 GND.n4128 585
R3572 GND.n4130 GND.n4129 585
R3573 GND.n3312 GND.n3310 585
R3574 GND.n3318 GND.n3310 585
R3575 GND.n4100 GND.n4099 585
R3576 GND.n4099 GND.n4098 585
R3577 GND.n3315 GND.n3314 585
R3578 GND.n3329 GND.n3315 585
R3579 GND.n4068 GND.n3340 585
R3580 GND.n3340 GND.n3326 585
R3581 GND.n4070 GND.n4069 585
R3582 GND.n4071 GND.n4070 585
R3583 GND.n3341 GND.n3339 585
R3584 GND.n3348 GND.n3339 585
R3585 GND.n4063 GND.n4062 585
R3586 GND.n4062 GND.n4061 585
R3587 GND.n3344 GND.n3343 585
R3588 GND.n3358 GND.n3344 585
R3589 GND.n4031 GND.n3369 585
R3590 GND.n3369 GND.n3356 585
R3591 GND.n4033 GND.n4032 585
R3592 GND.n4034 GND.n4033 585
R3593 GND.n3370 GND.n3368 585
R3594 GND.n3377 GND.n3368 585
R3595 GND.n4026 GND.n4025 585
R3596 GND.n4025 GND.n4024 585
R3597 GND.n3373 GND.n3372 585
R3598 GND.n3386 GND.n3373 585
R3599 GND.n3996 GND.n3995 585
R3600 GND.n3997 GND.n3996 585
R3601 GND.n3397 GND.n3396 585
R3602 GND.n3396 GND.n3395 585
R3603 GND.n3943 GND.n3942 585
R3604 GND.n3943 GND.n3921 585
R3605 GND.n3945 GND.n3944 585
R3606 GND.n3944 GND.n3920 585
R3607 GND.n3947 GND.n3946 585
R3608 GND.n3947 GND.n3936 585
R3609 GND.n3949 GND.n3948 585
R3610 GND.n3948 GND.n3934 585
R3611 GND.n3951 GND.n3950 585
R3612 GND.n3952 GND.n3951 585
R3613 GND.n3941 GND.n3940 585
R3614 GND.n3941 GND.n3419 585
R3615 GND.n3939 GND.n3938 585
R3616 GND.n3938 GND.n3417 585
R3617 GND.n3406 GND.n3404 585
R3618 GND.n3410 GND.n3406 585
R3619 GND.n3991 GND.n3990 585
R3620 GND.n3990 GND.n3989 585
R3621 GND.n3405 GND.n3403 585
R3622 GND.n3433 GND.n3405 585
R3623 GND.n3874 GND.n3873 585
R3624 GND.n3874 GND.n3430 585
R3625 GND.n3876 GND.n3875 585
R3626 GND.n3875 GND.n3442 585
R3627 GND.n3877 GND.n3452 585
R3628 GND.n3452 GND.n3439 585
R3629 GND.n3879 GND.n3878 585
R3630 GND.n3880 GND.n3879 585
R3631 GND.n3453 GND.n3451 585
R3632 GND.n3460 GND.n3451 585
R3633 GND.n3866 GND.n3865 585
R3634 GND.n3865 GND.n3864 585
R3635 GND.n3456 GND.n3455 585
R3636 GND.n3470 GND.n3456 585
R3637 GND.n3834 GND.n3481 585
R3638 GND.n3481 GND.n3468 585
R3639 GND.n3836 GND.n3835 585
R3640 GND.n3837 GND.n3836 585
R3641 GND.n3482 GND.n3480 585
R3642 GND.n3489 GND.n3480 585
R3643 GND.n3829 GND.n3828 585
R3644 GND.n3828 GND.n3827 585
R3645 GND.n3485 GND.n3484 585
R3646 GND.n3499 GND.n3485 585
R3647 GND.n3797 GND.n3511 585
R3648 GND.n3511 GND.n3497 585
R3649 GND.n3799 GND.n3798 585
R3650 GND.n3800 GND.n3799 585
R3651 GND.n3512 GND.n3510 585
R3652 GND.n3518 GND.n3510 585
R3653 GND.n3792 GND.n3791 585
R3654 GND.n3791 GND.n3790 585
R3655 GND.n3515 GND.n3514 585
R3656 GND.n3778 GND.n3515 585
R3657 GND.n3531 GND.n3530 585
R3658 GND.n3532 GND.n3531 585
R3659 GND.n3526 GND.n3525 585
R3660 GND.n3525 GND.n1373 585
R3661 GND.n1326 GND.n1325 585
R3662 GND.n6382 GND.n1326 585
R3663 GND.n6385 GND.n6384 585
R3664 GND.n6384 GND.n6383 585
R3665 GND.n6386 GND.n1320 585
R3666 GND.n1320 GND.n1319 585
R3667 GND.n6388 GND.n6387 585
R3668 GND.n6389 GND.n6388 585
R3669 GND.n1318 GND.n1317 585
R3670 GND.n6390 GND.n1318 585
R3671 GND.n6393 GND.n6392 585
R3672 GND.n6392 GND.n6391 585
R3673 GND.n6394 GND.n1312 585
R3674 GND.n1312 GND.n1311 585
R3675 GND.n6396 GND.n6395 585
R3676 GND.n6397 GND.n6396 585
R3677 GND.n1310 GND.n1309 585
R3678 GND.n6398 GND.n1310 585
R3679 GND.n6401 GND.n6400 585
R3680 GND.n6400 GND.n6399 585
R3681 GND.n6402 GND.n1304 585
R3682 GND.n1304 GND.n1303 585
R3683 GND.n6404 GND.n6403 585
R3684 GND.n6405 GND.n6404 585
R3685 GND.n1302 GND.n1301 585
R3686 GND.n6406 GND.n1302 585
R3687 GND.n6409 GND.n6408 585
R3688 GND.n6408 GND.n6407 585
R3689 GND.n6410 GND.n1296 585
R3690 GND.n1296 GND.n1295 585
R3691 GND.n6412 GND.n6411 585
R3692 GND.n6413 GND.n6412 585
R3693 GND.n1294 GND.n1293 585
R3694 GND.n6414 GND.n1294 585
R3695 GND.n6417 GND.n6416 585
R3696 GND.n6416 GND.n6415 585
R3697 GND.n6418 GND.n1288 585
R3698 GND.n1288 GND.n1287 585
R3699 GND.n6420 GND.n6419 585
R3700 GND.n6421 GND.n6420 585
R3701 GND.n1286 GND.n1285 585
R3702 GND.n6422 GND.n1286 585
R3703 GND.n6425 GND.n6424 585
R3704 GND.n6424 GND.n6423 585
R3705 GND.n6426 GND.n1280 585
R3706 GND.n1280 GND.n1279 585
R3707 GND.n6428 GND.n6427 585
R3708 GND.n6429 GND.n6428 585
R3709 GND.n1278 GND.n1277 585
R3710 GND.n6430 GND.n1278 585
R3711 GND.n6433 GND.n6432 585
R3712 GND.n6432 GND.n6431 585
R3713 GND.n6434 GND.n1272 585
R3714 GND.n1272 GND.n1271 585
R3715 GND.n6436 GND.n6435 585
R3716 GND.n6437 GND.n6436 585
R3717 GND.n1270 GND.n1269 585
R3718 GND.n6438 GND.n1270 585
R3719 GND.n6441 GND.n6440 585
R3720 GND.n6440 GND.n6439 585
R3721 GND.n6442 GND.n1264 585
R3722 GND.n1264 GND.n1263 585
R3723 GND.n6444 GND.n6443 585
R3724 GND.n6445 GND.n6444 585
R3725 GND.n1262 GND.n1261 585
R3726 GND.n6446 GND.n1262 585
R3727 GND.n6449 GND.n6448 585
R3728 GND.n6448 GND.n6447 585
R3729 GND.n6450 GND.n1256 585
R3730 GND.n1256 GND.n1255 585
R3731 GND.n6452 GND.n6451 585
R3732 GND.n6453 GND.n6452 585
R3733 GND.n1254 GND.n1253 585
R3734 GND.n6454 GND.n1254 585
R3735 GND.n6457 GND.n6456 585
R3736 GND.n6456 GND.n6455 585
R3737 GND.n6458 GND.n1248 585
R3738 GND.n1248 GND.n1247 585
R3739 GND.n6460 GND.n6459 585
R3740 GND.n6461 GND.n6460 585
R3741 GND.n1246 GND.n1245 585
R3742 GND.n6462 GND.n1246 585
R3743 GND.n6465 GND.n6464 585
R3744 GND.n6464 GND.n6463 585
R3745 GND.n6466 GND.n1240 585
R3746 GND.n1240 GND.n1239 585
R3747 GND.n6468 GND.n6467 585
R3748 GND.n6469 GND.n6468 585
R3749 GND.n1238 GND.n1237 585
R3750 GND.n6470 GND.n1238 585
R3751 GND.n6473 GND.n6472 585
R3752 GND.n6472 GND.n6471 585
R3753 GND.n6474 GND.n1232 585
R3754 GND.n1232 GND.n1231 585
R3755 GND.n6476 GND.n6475 585
R3756 GND.n6477 GND.n6476 585
R3757 GND.n1230 GND.n1229 585
R3758 GND.n6478 GND.n1230 585
R3759 GND.n6481 GND.n6480 585
R3760 GND.n6480 GND.n6479 585
R3761 GND.n6482 GND.n1224 585
R3762 GND.n1224 GND.n1223 585
R3763 GND.n6484 GND.n6483 585
R3764 GND.n6485 GND.n6484 585
R3765 GND.n1222 GND.n1221 585
R3766 GND.n6486 GND.n1222 585
R3767 GND.n6489 GND.n6488 585
R3768 GND.n6488 GND.n6487 585
R3769 GND.n6490 GND.n1216 585
R3770 GND.n1216 GND.n1215 585
R3771 GND.n6492 GND.n6491 585
R3772 GND.n6493 GND.n6492 585
R3773 GND.n1214 GND.n1213 585
R3774 GND.n6494 GND.n1214 585
R3775 GND.n6497 GND.n6496 585
R3776 GND.n6496 GND.n6495 585
R3777 GND.n6498 GND.n1210 585
R3778 GND.n1210 GND.n1209 585
R3779 GND.n6380 GND.n6379 585
R3780 GND.n6381 GND.n6380 585
R3781 GND.n6378 GND.n1375 585
R3782 GND.n1379 GND.n1377 585
R3783 GND.n6374 GND.n1380 585
R3784 GND.n6373 GND.n1381 585
R3785 GND.n6372 GND.n1382 585
R3786 GND.n1385 GND.n1383 585
R3787 GND.n6368 GND.n1386 585
R3788 GND.n6367 GND.n1387 585
R3789 GND.n6366 GND.n1388 585
R3790 GND.n1391 GND.n1389 585
R3791 GND.n6362 GND.n1392 585
R3792 GND.n6361 GND.n1393 585
R3793 GND.n6360 GND.n1394 585
R3794 GND.n1397 GND.n1395 585
R3795 GND.n6356 GND.n1398 585
R3796 GND.n6355 GND.n6352 585
R3797 GND.n6351 GND.n1372 585
R3798 GND.n6381 GND.n1372 585
R3799 GND.n4153 GND.n3170 585
R3800 GND.n4154 GND.n4153 585
R3801 GND.n4152 GND.n3292 585
R3802 GND.n4152 GND.n4151 585
R3803 GND.n3304 GND.n3291 585
R3804 GND.n4135 GND.n3291 585
R3805 GND.n4141 GND.n4140 585
R3806 GND.n4142 GND.n4141 585
R3807 GND.n3303 GND.n3302 585
R3808 GND.n4132 GND.n3302 585
R3809 GND.n4078 GND.n4077 585
R3810 GND.n4077 GND.n3309 585
R3811 GND.n4076 GND.n3319 585
R3812 GND.n4097 GND.n3319 585
R3813 GND.n3333 GND.n3331 585
R3814 GND.n3331 GND.n3316 585
R3815 GND.n4086 GND.n4085 585
R3816 GND.n4087 GND.n4086 585
R3817 GND.n3332 GND.n3330 585
R3818 GND.n4072 GND.n3330 585
R3819 GND.n4041 GND.n4040 585
R3820 GND.n4040 GND.n3338 585
R3821 GND.n4039 GND.n3349 585
R3822 GND.n4060 GND.n3349 585
R3823 GND.n3362 GND.n3360 585
R3824 GND.n3360 GND.n3346 585
R3825 GND.n4049 GND.n4048 585
R3826 GND.n4050 GND.n4049 585
R3827 GND.n3361 GND.n3359 585
R3828 GND.n4035 GND.n3359 585
R3829 GND.n4004 GND.n4003 585
R3830 GND.n4003 GND.n3367 585
R3831 GND.n4002 GND.n3378 585
R3832 GND.n4023 GND.n3378 585
R3833 GND.n3390 GND.n3388 585
R3834 GND.n3388 GND.n3374 585
R3835 GND.n4012 GND.n4011 585
R3836 GND.n4013 GND.n4012 585
R3837 GND.n3389 GND.n3387 585
R3838 GND.n3998 GND.n3387 585
R3839 GND.n3928 GND.n3927 585
R3840 GND.n3929 GND.n3928 585
R3841 GND.n3925 GND.n3922 585
R3842 GND.n3968 GND.n3922 585
R3843 GND.n3957 GND.n3917 585
R3844 GND.n3957 GND.n3956 585
R3845 GND.n3958 GND.n3916 585
R3846 GND.n3959 GND.n3958 585
R3847 GND.n3955 GND.n3915 585
R3848 GND.n3955 GND.n3954 585
R3849 GND.n3423 GND.n3421 585
R3850 GND.n3937 GND.n3421 585
R3851 GND.n3980 GND.n3979 585
R3852 GND.n3981 GND.n3980 585
R3853 GND.n3422 GND.n3420 585
R3854 GND.n3909 GND.n3420 585
R3855 GND.n3906 GND.n3411 585
R3856 GND.n3988 GND.n3411 585
R3857 GND.n3905 GND.n3904 585
R3858 GND.n3904 GND.n3407 585
R3859 GND.n3903 GND.n3428 585
R3860 GND.n3903 GND.n3902 585
R3861 GND.n3445 GND.n3429 585
R3862 GND.n3884 GND.n3429 585
R3863 GND.n3892 GND.n3891 585
R3864 GND.n3893 GND.n3892 585
R3865 GND.n3444 GND.n3443 585
R3866 GND.n3881 GND.n3443 585
R3867 GND.n3844 GND.n3843 585
R3868 GND.n3843 GND.n3450 585
R3869 GND.n3842 GND.n3461 585
R3870 GND.n3863 GND.n3461 585
R3871 GND.n3474 GND.n3472 585
R3872 GND.n3472 GND.n3458 585
R3873 GND.n3852 GND.n3851 585
R3874 GND.n3853 GND.n3852 585
R3875 GND.n3473 GND.n3471 585
R3876 GND.n3838 GND.n3471 585
R3877 GND.n3807 GND.n3806 585
R3878 GND.n3806 GND.n3479 585
R3879 GND.n3805 GND.n3490 585
R3880 GND.n3826 GND.n3490 585
R3881 GND.n3503 GND.n3501 585
R3882 GND.n3501 GND.n3486 585
R3883 GND.n3815 GND.n3814 585
R3884 GND.n3816 GND.n3815 585
R3885 GND.n3502 GND.n3500 585
R3886 GND.n3801 GND.n3500 585
R3887 GND.n3770 GND.n3769 585
R3888 GND.n3769 GND.n3509 585
R3889 GND.n3768 GND.n3519 585
R3890 GND.n3789 GND.n3519 585
R3891 GND.n3767 GND.n3766 585
R3892 GND.n3766 GND.n3516 585
R3893 GND.n3765 GND.n1374 585
R3894 GND.n3779 GND.n1374 585
R3895 GND.n6275 GND.n6274 585
R3896 GND.n6274 GND.n6273 585
R3897 GND.n1463 GND.n1462 585
R3898 GND.n3124 GND.n3119 585
R3899 GND.n3125 GND.n3118 585
R3900 GND.n3126 GND.n3117 585
R3901 GND.n3116 GND.n3110 585
R3902 GND.n3133 GND.n3109 585
R3903 GND.n3134 GND.n3108 585
R3904 GND.n3103 GND.n3102 585
R3905 GND.n3144 GND.n3101 585
R3906 GND.n3145 GND.n3100 585
R3907 GND.n3099 GND.n3091 585
R3908 GND.n3152 GND.n3090 585
R3909 GND.n3153 GND.n3089 585
R3910 GND.n3083 GND.n3082 585
R3911 GND.n3160 GND.n3081 585
R3912 GND.n3161 GND.n3080 585
R3913 GND.n3079 GND.n1495 585
R3914 GND.n6273 GND.n1495 585
R3915 GND.n1464 GND.n1458 585
R3916 GND.n4154 GND.n1464 585
R3917 GND.n6279 GND.n1457 585
R3918 GND.n4151 GND.n1457 585
R3919 GND.n6280 GND.n1456 585
R3920 GND.n4135 GND.n1456 585
R3921 GND.n6281 GND.n1455 585
R3922 GND.n4142 GND.n1455 585
R3923 GND.n4131 GND.n1453 585
R3924 GND.n4132 GND.n4131 585
R3925 GND.n6285 GND.n1452 585
R3926 GND.n3309 GND.n1452 585
R3927 GND.n6286 GND.n1451 585
R3928 GND.n4097 GND.n1451 585
R3929 GND.n6287 GND.n1450 585
R3930 GND.n3316 GND.n1450 585
R3931 GND.n3328 GND.n1448 585
R3932 GND.n4087 GND.n3328 585
R3933 GND.n6291 GND.n1447 585
R3934 GND.n4072 GND.n1447 585
R3935 GND.n6292 GND.n1446 585
R3936 GND.n3338 GND.n1446 585
R3937 GND.n6293 GND.n1445 585
R3938 GND.n4060 GND.n1445 585
R3939 GND.n3345 GND.n1443 585
R3940 GND.n3346 GND.n3345 585
R3941 GND.n6297 GND.n1442 585
R3942 GND.n4050 GND.n1442 585
R3943 GND.n6298 GND.n1441 585
R3944 GND.n4035 GND.n1441 585
R3945 GND.n6299 GND.n1440 585
R3946 GND.n3367 GND.n1440 585
R3947 GND.n3376 GND.n1438 585
R3948 GND.n4023 GND.n3376 585
R3949 GND.n6303 GND.n1437 585
R3950 GND.n3374 GND.n1437 585
R3951 GND.n6304 GND.n1436 585
R3952 GND.n4013 GND.n1436 585
R3953 GND.n6305 GND.n1435 585
R3954 GND.n3998 GND.n1435 585
R3955 GND.n3924 GND.n1433 585
R3956 GND.n3929 GND.n3924 585
R3957 GND.n6309 GND.n1432 585
R3958 GND.n3968 GND.n1432 585
R3959 GND.n6310 GND.n1431 585
R3960 GND.n3956 GND.n1431 585
R3961 GND.n6311 GND.n1430 585
R3962 GND.n3959 GND.n1430 585
R3963 GND.n3953 GND.n1428 585
R3964 GND.n3954 GND.n3953 585
R3965 GND.n6316 GND.n1427 585
R3966 GND.n3937 GND.n1427 585
R3967 GND.n6317 GND.n1426 585
R3968 GND.n3981 GND.n1426 585
R3969 GND.n6318 GND.n1425 585
R3970 GND.n3909 GND.n1425 585
R3971 GND.n3409 GND.n1423 585
R3972 GND.n3988 GND.n3409 585
R3973 GND.n6322 GND.n1422 585
R3974 GND.n3407 GND.n1422 585
R3975 GND.n6323 GND.n1421 585
R3976 GND.n3902 GND.n1421 585
R3977 GND.n6324 GND.n1420 585
R3978 GND.n3884 GND.n1420 585
R3979 GND.n3441 GND.n1418 585
R3980 GND.n3893 GND.n3441 585
R3981 GND.n6328 GND.n1417 585
R3982 GND.n3881 GND.n1417 585
R3983 GND.n6329 GND.n1416 585
R3984 GND.n3450 GND.n1416 585
R3985 GND.n6330 GND.n1415 585
R3986 GND.n3863 GND.n1415 585
R3987 GND.n3457 GND.n1413 585
R3988 GND.n3458 GND.n3457 585
R3989 GND.n6334 GND.n1412 585
R3990 GND.n3853 GND.n1412 585
R3991 GND.n6335 GND.n1411 585
R3992 GND.n3838 GND.n1411 585
R3993 GND.n6336 GND.n1410 585
R3994 GND.n3479 GND.n1410 585
R3995 GND.n3488 GND.n1408 585
R3996 GND.n3826 GND.n3488 585
R3997 GND.n6340 GND.n1407 585
R3998 GND.n3486 GND.n1407 585
R3999 GND.n6341 GND.n1406 585
R4000 GND.n3816 GND.n1406 585
R4001 GND.n6342 GND.n1405 585
R4002 GND.n3801 GND.n1405 585
R4003 GND.n3508 GND.n1403 585
R4004 GND.n3509 GND.n3508 585
R4005 GND.n6346 GND.n1402 585
R4006 GND.n3789 GND.n1402 585
R4007 GND.n6347 GND.n1401 585
R4008 GND.n3516 GND.n1401 585
R4009 GND.n6348 GND.n1400 585
R4010 GND.n3779 GND.n1400 585
R4011 GND.n5938 GND.n5835 502.111
R4012 GND.n5941 GND.n5940 502.111
R4013 GND.n4651 GND.n4580 502.111
R4014 GND.n6213 GND.n1616 502.111
R4015 GND.n6220 GND.n6219 402.176
R4016 GND.n5521 GND.n1890 402.176
R4017 GND.n7754 GND.n412 395.481
R4018 GND.n7595 GND.n7594 301.784
R4019 GND.n7595 GND.n502 301.784
R4020 GND.n7603 GND.n502 301.784
R4021 GND.n7604 GND.n7603 301.784
R4022 GND.n7605 GND.n7604 301.784
R4023 GND.n7605 GND.n496 301.784
R4024 GND.n7613 GND.n496 301.784
R4025 GND.n7614 GND.n7613 301.784
R4026 GND.n7615 GND.n7614 301.784
R4027 GND.n7615 GND.n490 301.784
R4028 GND.n7623 GND.n490 301.784
R4029 GND.n7624 GND.n7623 301.784
R4030 GND.n7625 GND.n7624 301.784
R4031 GND.n7625 GND.n484 301.784
R4032 GND.n7633 GND.n484 301.784
R4033 GND.n7634 GND.n7633 301.784
R4034 GND.n7635 GND.n7634 301.784
R4035 GND.n7635 GND.n478 301.784
R4036 GND.n7643 GND.n478 301.784
R4037 GND.n7644 GND.n7643 301.784
R4038 GND.n7645 GND.n7644 301.784
R4039 GND.n7645 GND.n472 301.784
R4040 GND.n7653 GND.n472 301.784
R4041 GND.n7654 GND.n7653 301.784
R4042 GND.n7655 GND.n7654 301.784
R4043 GND.n7655 GND.n466 301.784
R4044 GND.n7663 GND.n466 301.784
R4045 GND.n7664 GND.n7663 301.784
R4046 GND.n7665 GND.n7664 301.784
R4047 GND.n7665 GND.n460 301.784
R4048 GND.n7673 GND.n460 301.784
R4049 GND.n7674 GND.n7673 301.784
R4050 GND.n7675 GND.n7674 301.784
R4051 GND.n7675 GND.n454 301.784
R4052 GND.n7683 GND.n454 301.784
R4053 GND.n7684 GND.n7683 301.784
R4054 GND.n7685 GND.n7684 301.784
R4055 GND.n7685 GND.n448 301.784
R4056 GND.n7693 GND.n448 301.784
R4057 GND.n7694 GND.n7693 301.784
R4058 GND.n7695 GND.n7694 301.784
R4059 GND.n7695 GND.n442 301.784
R4060 GND.n7703 GND.n442 301.784
R4061 GND.n7704 GND.n7703 301.784
R4062 GND.n7705 GND.n7704 301.784
R4063 GND.n7705 GND.n436 301.784
R4064 GND.n7713 GND.n436 301.784
R4065 GND.n7714 GND.n7713 301.784
R4066 GND.n7715 GND.n7714 301.784
R4067 GND.n7715 GND.n430 301.784
R4068 GND.n7723 GND.n430 301.784
R4069 GND.n7724 GND.n7723 301.784
R4070 GND.n7725 GND.n7724 301.784
R4071 GND.n7725 GND.n424 301.784
R4072 GND.n7733 GND.n424 301.784
R4073 GND.n7734 GND.n7733 301.784
R4074 GND.n7735 GND.n7734 301.784
R4075 GND.n7735 GND.n418 301.784
R4076 GND.n7744 GND.n418 301.784
R4077 GND.n7745 GND.n7744 301.784
R4078 GND.n7746 GND.n7745 301.784
R4079 GND.n7746 GND.n412 301.784
R4080 GND.n6149 GND.t141 281.95
R4081 GND.n4581 GND.t76 281.95
R4082 GND.n1891 GND.t111 281.95
R4083 GND.n5865 GND.t42 281.95
R4084 GND.n6633 GND.n1084 280.613
R4085 GND.n6634 GND.n6633 280.613
R4086 GND.n6635 GND.n6634 280.613
R4087 GND.n6635 GND.n1078 280.613
R4088 GND.n6643 GND.n1078 280.613
R4089 GND.n6644 GND.n6643 280.613
R4090 GND.n6645 GND.n6644 280.613
R4091 GND.n6645 GND.n1072 280.613
R4092 GND.n6653 GND.n1072 280.613
R4093 GND.n6654 GND.n6653 280.613
R4094 GND.n6655 GND.n6654 280.613
R4095 GND.n6655 GND.n1066 280.613
R4096 GND.n6663 GND.n1066 280.613
R4097 GND.n6664 GND.n6663 280.613
R4098 GND.n6665 GND.n6664 280.613
R4099 GND.n6665 GND.n1060 280.613
R4100 GND.n6673 GND.n1060 280.613
R4101 GND.n6674 GND.n6673 280.613
R4102 GND.n6675 GND.n6674 280.613
R4103 GND.n6675 GND.n1054 280.613
R4104 GND.n6683 GND.n1054 280.613
R4105 GND.n6684 GND.n6683 280.613
R4106 GND.n6685 GND.n6684 280.613
R4107 GND.n6685 GND.n1048 280.613
R4108 GND.n6693 GND.n1048 280.613
R4109 GND.n6694 GND.n6693 280.613
R4110 GND.n6695 GND.n6694 280.613
R4111 GND.n6695 GND.n1042 280.613
R4112 GND.n6703 GND.n1042 280.613
R4113 GND.n6704 GND.n6703 280.613
R4114 GND.n6705 GND.n6704 280.613
R4115 GND.n6705 GND.n1036 280.613
R4116 GND.n6713 GND.n1036 280.613
R4117 GND.n6714 GND.n6713 280.613
R4118 GND.n6715 GND.n6714 280.613
R4119 GND.n6715 GND.n1030 280.613
R4120 GND.n6723 GND.n1030 280.613
R4121 GND.n6724 GND.n6723 280.613
R4122 GND.n6725 GND.n6724 280.613
R4123 GND.n6725 GND.n1024 280.613
R4124 GND.n6733 GND.n1024 280.613
R4125 GND.n6734 GND.n6733 280.613
R4126 GND.n6735 GND.n6734 280.613
R4127 GND.n6735 GND.n1018 280.613
R4128 GND.n6743 GND.n1018 280.613
R4129 GND.n6744 GND.n6743 280.613
R4130 GND.n6745 GND.n6744 280.613
R4131 GND.n6745 GND.n1012 280.613
R4132 GND.n6753 GND.n1012 280.613
R4133 GND.n6754 GND.n6753 280.613
R4134 GND.n6755 GND.n6754 280.613
R4135 GND.n6755 GND.n1006 280.613
R4136 GND.n6763 GND.n1006 280.613
R4137 GND.n6764 GND.n6763 280.613
R4138 GND.n6765 GND.n6764 280.613
R4139 GND.n6765 GND.n1000 280.613
R4140 GND.n6773 GND.n1000 280.613
R4141 GND.n6774 GND.n6773 280.613
R4142 GND.n6775 GND.n6774 280.613
R4143 GND.n6775 GND.n994 280.613
R4144 GND.n6783 GND.n994 280.613
R4145 GND.n6784 GND.n6783 280.613
R4146 GND.n6785 GND.n6784 280.613
R4147 GND.n6785 GND.n988 280.613
R4148 GND.n6793 GND.n988 280.613
R4149 GND.n6794 GND.n6793 280.613
R4150 GND.n6795 GND.n6794 280.613
R4151 GND.n6795 GND.n982 280.613
R4152 GND.n6803 GND.n982 280.613
R4153 GND.n6804 GND.n6803 280.613
R4154 GND.n6805 GND.n6804 280.613
R4155 GND.n6805 GND.n976 280.613
R4156 GND.n6813 GND.n976 280.613
R4157 GND.n6814 GND.n6813 280.613
R4158 GND.n6815 GND.n6814 280.613
R4159 GND.n6815 GND.n970 280.613
R4160 GND.n6823 GND.n970 280.613
R4161 GND.n6824 GND.n6823 280.613
R4162 GND.n6825 GND.n6824 280.613
R4163 GND.n6825 GND.n964 280.613
R4164 GND.n6833 GND.n964 280.613
R4165 GND.n6834 GND.n6833 280.613
R4166 GND.n6835 GND.n6834 280.613
R4167 GND.n6835 GND.n958 280.613
R4168 GND.n6843 GND.n958 280.613
R4169 GND.n6844 GND.n6843 280.613
R4170 GND.n6845 GND.n6844 280.613
R4171 GND.n6845 GND.n952 280.613
R4172 GND.n6853 GND.n952 280.613
R4173 GND.n6854 GND.n6853 280.613
R4174 GND.n6855 GND.n6854 280.613
R4175 GND.n6855 GND.n946 280.613
R4176 GND.n6863 GND.n946 280.613
R4177 GND.n6864 GND.n6863 280.613
R4178 GND.n6865 GND.n6864 280.613
R4179 GND.n6865 GND.n940 280.613
R4180 GND.n6873 GND.n940 280.613
R4181 GND.n6874 GND.n6873 280.613
R4182 GND.n6875 GND.n6874 280.613
R4183 GND.n6875 GND.n934 280.613
R4184 GND.n6883 GND.n934 280.613
R4185 GND.n6884 GND.n6883 280.613
R4186 GND.n6885 GND.n6884 280.613
R4187 GND.n6885 GND.n928 280.613
R4188 GND.n6893 GND.n928 280.613
R4189 GND.n6894 GND.n6893 280.613
R4190 GND.n6895 GND.n6894 280.613
R4191 GND.n6895 GND.n922 280.613
R4192 GND.n6903 GND.n922 280.613
R4193 GND.n6904 GND.n6903 280.613
R4194 GND.n6905 GND.n6904 280.613
R4195 GND.n6905 GND.n916 280.613
R4196 GND.n6913 GND.n916 280.613
R4197 GND.n6914 GND.n6913 280.613
R4198 GND.n6915 GND.n6914 280.613
R4199 GND.n6915 GND.n910 280.613
R4200 GND.n6923 GND.n910 280.613
R4201 GND.n6924 GND.n6923 280.613
R4202 GND.n6925 GND.n6924 280.613
R4203 GND.n6925 GND.n904 280.613
R4204 GND.n6933 GND.n904 280.613
R4205 GND.n6934 GND.n6933 280.613
R4206 GND.n6935 GND.n6934 280.613
R4207 GND.n6935 GND.n898 280.613
R4208 GND.n6943 GND.n898 280.613
R4209 GND.n6944 GND.n6943 280.613
R4210 GND.n6945 GND.n6944 280.613
R4211 GND.n6945 GND.n892 280.613
R4212 GND.n6953 GND.n892 280.613
R4213 GND.n6954 GND.n6953 280.613
R4214 GND.n6955 GND.n6954 280.613
R4215 GND.n6955 GND.n886 280.613
R4216 GND.n6963 GND.n886 280.613
R4217 GND.n6964 GND.n6963 280.613
R4218 GND.n6965 GND.n6964 280.613
R4219 GND.n6965 GND.n880 280.613
R4220 GND.n6973 GND.n880 280.613
R4221 GND.n6974 GND.n6973 280.613
R4222 GND.n6975 GND.n6974 280.613
R4223 GND.n6975 GND.n874 280.613
R4224 GND.n6983 GND.n874 280.613
R4225 GND.n6984 GND.n6983 280.613
R4226 GND.n6985 GND.n6984 280.613
R4227 GND.n6985 GND.n868 280.613
R4228 GND.n6993 GND.n868 280.613
R4229 GND.n6994 GND.n6993 280.613
R4230 GND.n6995 GND.n6994 280.613
R4231 GND.n6995 GND.n862 280.613
R4232 GND.n7003 GND.n862 280.613
R4233 GND.n7004 GND.n7003 280.613
R4234 GND.n7005 GND.n7004 280.613
R4235 GND.n7005 GND.n856 280.613
R4236 GND.n7013 GND.n856 280.613
R4237 GND.n7014 GND.n7013 280.613
R4238 GND.n7015 GND.n7014 280.613
R4239 GND.n7015 GND.n850 280.613
R4240 GND.n7023 GND.n850 280.613
R4241 GND.n7024 GND.n7023 280.613
R4242 GND.n7025 GND.n7024 280.613
R4243 GND.n7025 GND.n844 280.613
R4244 GND.n7033 GND.n844 280.613
R4245 GND.n7034 GND.n7033 280.613
R4246 GND.n7035 GND.n7034 280.613
R4247 GND.n7035 GND.n838 280.613
R4248 GND.n7043 GND.n838 280.613
R4249 GND.n7044 GND.n7043 280.613
R4250 GND.n7045 GND.n7044 280.613
R4251 GND.n7045 GND.n832 280.613
R4252 GND.n7053 GND.n832 280.613
R4253 GND.n7054 GND.n7053 280.613
R4254 GND.n7055 GND.n7054 280.613
R4255 GND.n7055 GND.n826 280.613
R4256 GND.n7063 GND.n826 280.613
R4257 GND.n7064 GND.n7063 280.613
R4258 GND.n7065 GND.n7064 280.613
R4259 GND.n7065 GND.n820 280.613
R4260 GND.n7073 GND.n820 280.613
R4261 GND.n7074 GND.n7073 280.613
R4262 GND.n7075 GND.n7074 280.613
R4263 GND.n7075 GND.n814 280.613
R4264 GND.n7083 GND.n814 280.613
R4265 GND.n7084 GND.n7083 280.613
R4266 GND.n7085 GND.n7084 280.613
R4267 GND.n7085 GND.n808 280.613
R4268 GND.n7093 GND.n808 280.613
R4269 GND.n7094 GND.n7093 280.613
R4270 GND.n7095 GND.n7094 280.613
R4271 GND.n7095 GND.n802 280.613
R4272 GND.n7103 GND.n802 280.613
R4273 GND.n7104 GND.n7103 280.613
R4274 GND.n7105 GND.n7104 280.613
R4275 GND.n7105 GND.n796 280.613
R4276 GND.n7113 GND.n796 280.613
R4277 GND.n7114 GND.n7113 280.613
R4278 GND.n7115 GND.n7114 280.613
R4279 GND.n7115 GND.n790 280.613
R4280 GND.n7123 GND.n790 280.613
R4281 GND.n7124 GND.n7123 280.613
R4282 GND.n7125 GND.n7124 280.613
R4283 GND.n7125 GND.n784 280.613
R4284 GND.n7133 GND.n784 280.613
R4285 GND.n7134 GND.n7133 280.613
R4286 GND.n7135 GND.n7134 280.613
R4287 GND.n7135 GND.n778 280.613
R4288 GND.n7143 GND.n778 280.613
R4289 GND.n7144 GND.n7143 280.613
R4290 GND.n7145 GND.n7144 280.613
R4291 GND.n7145 GND.n772 280.613
R4292 GND.n7153 GND.n772 280.613
R4293 GND.n7154 GND.n7153 280.613
R4294 GND.n7155 GND.n7154 280.613
R4295 GND.n7155 GND.n766 280.613
R4296 GND.n7163 GND.n766 280.613
R4297 GND.n7164 GND.n7163 280.613
R4298 GND.n7165 GND.n7164 280.613
R4299 GND.n7165 GND.n760 280.613
R4300 GND.n7173 GND.n760 280.613
R4301 GND.n7174 GND.n7173 280.613
R4302 GND.n7175 GND.n7174 280.613
R4303 GND.n7175 GND.n754 280.613
R4304 GND.n7183 GND.n754 280.613
R4305 GND.n7184 GND.n7183 280.613
R4306 GND.n7185 GND.n7184 280.613
R4307 GND.n7185 GND.n748 280.613
R4308 GND.n7193 GND.n748 280.613
R4309 GND.n7194 GND.n7193 280.613
R4310 GND.n7195 GND.n7194 280.613
R4311 GND.n7195 GND.n742 280.613
R4312 GND.n7203 GND.n742 280.613
R4313 GND.n7204 GND.n7203 280.613
R4314 GND.n7205 GND.n7204 280.613
R4315 GND.n7205 GND.n736 280.613
R4316 GND.n7213 GND.n736 280.613
R4317 GND.n7214 GND.n7213 280.613
R4318 GND.n7215 GND.n7214 280.613
R4319 GND.n7215 GND.n730 280.613
R4320 GND.n7223 GND.n730 280.613
R4321 GND.n7224 GND.n7223 280.613
R4322 GND.n7225 GND.n7224 280.613
R4323 GND.n7225 GND.n724 280.613
R4324 GND.n7233 GND.n724 280.613
R4325 GND.n7234 GND.n7233 280.613
R4326 GND.n7235 GND.n7234 280.613
R4327 GND.n7235 GND.n718 280.613
R4328 GND.n7243 GND.n718 280.613
R4329 GND.n7244 GND.n7243 280.613
R4330 GND.n7245 GND.n7244 280.613
R4331 GND.n7245 GND.n712 280.613
R4332 GND.n7253 GND.n712 280.613
R4333 GND.n7254 GND.n7253 280.613
R4334 GND.n7255 GND.n7254 280.613
R4335 GND.n7255 GND.n706 280.613
R4336 GND.n7263 GND.n706 280.613
R4337 GND.n7264 GND.n7263 280.613
R4338 GND.n7265 GND.n7264 280.613
R4339 GND.n7265 GND.n700 280.613
R4340 GND.n7273 GND.n700 280.613
R4341 GND.n7274 GND.n7273 280.613
R4342 GND.n7275 GND.n7274 280.613
R4343 GND.n7275 GND.n694 280.613
R4344 GND.n7283 GND.n694 280.613
R4345 GND.n7284 GND.n7283 280.613
R4346 GND.n7285 GND.n7284 280.613
R4347 GND.n7285 GND.n688 280.613
R4348 GND.n7293 GND.n688 280.613
R4349 GND.n7294 GND.n7293 280.613
R4350 GND.n7295 GND.n7294 280.613
R4351 GND.n7295 GND.n682 280.613
R4352 GND.n7303 GND.n682 280.613
R4353 GND.n7304 GND.n7303 280.613
R4354 GND.n7305 GND.n7304 280.613
R4355 GND.n7305 GND.n676 280.613
R4356 GND.n7313 GND.n676 280.613
R4357 GND.n7314 GND.n7313 280.613
R4358 GND.n7315 GND.n7314 280.613
R4359 GND.n7315 GND.n670 280.613
R4360 GND.n7323 GND.n670 280.613
R4361 GND.n7324 GND.n7323 280.613
R4362 GND.n7325 GND.n7324 280.613
R4363 GND.n7325 GND.n664 280.613
R4364 GND.n7333 GND.n664 280.613
R4365 GND.n7334 GND.n7333 280.613
R4366 GND.n7335 GND.n7334 280.613
R4367 GND.n7335 GND.n658 280.613
R4368 GND.n7343 GND.n658 280.613
R4369 GND.n7344 GND.n7343 280.613
R4370 GND.n7345 GND.n7344 280.613
R4371 GND.n7345 GND.n652 280.613
R4372 GND.n7353 GND.n652 280.613
R4373 GND.n7354 GND.n7353 280.613
R4374 GND.n7355 GND.n7354 280.613
R4375 GND.n7355 GND.n646 280.613
R4376 GND.n7363 GND.n646 280.613
R4377 GND.n7364 GND.n7363 280.613
R4378 GND.n7365 GND.n7364 280.613
R4379 GND.n7365 GND.n640 280.613
R4380 GND.n7373 GND.n640 280.613
R4381 GND.n7374 GND.n7373 280.613
R4382 GND.n7375 GND.n7374 280.613
R4383 GND.n7375 GND.n634 280.613
R4384 GND.n7383 GND.n634 280.613
R4385 GND.n7384 GND.n7383 280.613
R4386 GND.n7385 GND.n7384 280.613
R4387 GND.n7385 GND.n628 280.613
R4388 GND.n7393 GND.n628 280.613
R4389 GND.n7394 GND.n7393 280.613
R4390 GND.n7395 GND.n7394 280.613
R4391 GND.n7395 GND.n622 280.613
R4392 GND.n7403 GND.n622 280.613
R4393 GND.n7404 GND.n7403 280.613
R4394 GND.n7405 GND.n7404 280.613
R4395 GND.n7405 GND.n616 280.613
R4396 GND.n7413 GND.n616 280.613
R4397 GND.n7414 GND.n7413 280.613
R4398 GND.n7415 GND.n7414 280.613
R4399 GND.n7415 GND.n610 280.613
R4400 GND.n7423 GND.n610 280.613
R4401 GND.n7424 GND.n7423 280.613
R4402 GND.n7425 GND.n7424 280.613
R4403 GND.n7425 GND.n604 280.613
R4404 GND.n7433 GND.n604 280.613
R4405 GND.n7434 GND.n7433 280.613
R4406 GND.n7435 GND.n7434 280.613
R4407 GND.n7435 GND.n598 280.613
R4408 GND.n7443 GND.n598 280.613
R4409 GND.n7444 GND.n7443 280.613
R4410 GND.n7445 GND.n7444 280.613
R4411 GND.n7445 GND.n592 280.613
R4412 GND.n7453 GND.n592 280.613
R4413 GND.n7454 GND.n7453 280.613
R4414 GND.n7455 GND.n7454 280.613
R4415 GND.n7455 GND.n586 280.613
R4416 GND.n7463 GND.n586 280.613
R4417 GND.n7464 GND.n7463 280.613
R4418 GND.n7465 GND.n7464 280.613
R4419 GND.n7465 GND.n580 280.613
R4420 GND.n7473 GND.n580 280.613
R4421 GND.n7474 GND.n7473 280.613
R4422 GND.n7475 GND.n7474 280.613
R4423 GND.n7475 GND.n574 280.613
R4424 GND.n7483 GND.n574 280.613
R4425 GND.n7484 GND.n7483 280.613
R4426 GND.n7485 GND.n7484 280.613
R4427 GND.n7485 GND.n568 280.613
R4428 GND.n7493 GND.n568 280.613
R4429 GND.n7494 GND.n7493 280.613
R4430 GND.n7495 GND.n7494 280.613
R4431 GND.n7495 GND.n562 280.613
R4432 GND.n7503 GND.n562 280.613
R4433 GND.n7504 GND.n7503 280.613
R4434 GND.n7505 GND.n7504 280.613
R4435 GND.n7505 GND.n556 280.613
R4436 GND.n7513 GND.n556 280.613
R4437 GND.n7514 GND.n7513 280.613
R4438 GND.n7515 GND.n7514 280.613
R4439 GND.n7515 GND.n550 280.613
R4440 GND.n7523 GND.n550 280.613
R4441 GND.n7524 GND.n7523 280.613
R4442 GND.n7525 GND.n7524 280.613
R4443 GND.n7525 GND.n544 280.613
R4444 GND.n7533 GND.n544 280.613
R4445 GND.n7534 GND.n7533 280.613
R4446 GND.n7535 GND.n7534 280.613
R4447 GND.n7535 GND.n538 280.613
R4448 GND.n7543 GND.n538 280.613
R4449 GND.n7544 GND.n7543 280.613
R4450 GND.n7545 GND.n7544 280.613
R4451 GND.n7545 GND.n532 280.613
R4452 GND.n7553 GND.n532 280.613
R4453 GND.n7554 GND.n7553 280.613
R4454 GND.n7555 GND.n7554 280.613
R4455 GND.n7555 GND.n526 280.613
R4456 GND.n7563 GND.n526 280.613
R4457 GND.n7564 GND.n7563 280.613
R4458 GND.n7565 GND.n7564 280.613
R4459 GND.n7565 GND.n520 280.613
R4460 GND.n7573 GND.n520 280.613
R4461 GND.n7574 GND.n7573 280.613
R4462 GND.n7575 GND.n7574 280.613
R4463 GND.n7575 GND.n514 280.613
R4464 GND.n7583 GND.n514 280.613
R4465 GND.n7584 GND.n7583 280.613
R4466 GND.n7585 GND.n7584 280.613
R4467 GND.n7585 GND.n508 280.613
R4468 GND.n7593 GND.n508 280.613
R4469 GND.n1625 GND.t119 260.649
R4470 GND.n5855 GND.t110 260.649
R4471 GND.n6215 GND.n6214 256.663
R4472 GND.n6215 GND.n1579 256.663
R4473 GND.n6215 GND.n1580 256.663
R4474 GND.n6215 GND.n1581 256.663
R4475 GND.n6215 GND.n1582 256.663
R4476 GND.n6215 GND.n1583 256.663
R4477 GND.n6215 GND.n1584 256.663
R4478 GND.n6215 GND.n1585 256.663
R4479 GND.n6215 GND.n1586 256.663
R4480 GND.n6215 GND.n1587 256.663
R4481 GND.n6215 GND.n1588 256.663
R4482 GND.n6215 GND.n1589 256.663
R4483 GND.n6215 GND.n1590 256.663
R4484 GND.n6215 GND.n1591 256.663
R4485 GND.n6215 GND.n1592 256.663
R4486 GND.n6215 GND.n1593 256.663
R4487 GND.n6216 GND.n6215 256.663
R4488 GND.n6219 GND.n1575 256.663
R4489 GND.n6215 GND.n1594 256.663
R4490 GND.n6215 GND.n1596 256.663
R4491 GND.n6215 GND.n1597 256.663
R4492 GND.n6215 GND.n1598 256.663
R4493 GND.n6215 GND.n1599 256.663
R4494 GND.n6215 GND.n1600 256.663
R4495 GND.n6215 GND.n1601 256.663
R4496 GND.n6215 GND.n1602 256.663
R4497 GND.n6215 GND.n1603 256.663
R4498 GND.n6215 GND.n1604 256.663
R4499 GND.n6215 GND.n1605 256.663
R4500 GND.n6215 GND.n1606 256.663
R4501 GND.n6215 GND.n1607 256.663
R4502 GND.n6215 GND.n1608 256.663
R4503 GND.n6215 GND.n1609 256.663
R4504 GND.n6215 GND.n1610 256.663
R4505 GND.n6215 GND.n1611 256.663
R4506 GND.n6215 GND.n1612 256.663
R4507 GND.n6011 GND.n1872 256.663
R4508 GND.n6011 GND.n1873 256.663
R4509 GND.n6011 GND.n1874 256.663
R4510 GND.n6011 GND.n1875 256.663
R4511 GND.n6011 GND.n1876 256.663
R4512 GND.n6011 GND.n1877 256.663
R4513 GND.n6011 GND.n1878 256.663
R4514 GND.n6011 GND.n1879 256.663
R4515 GND.n6011 GND.n1880 256.663
R4516 GND.n6011 GND.n1881 256.663
R4517 GND.n6011 GND.n1882 256.663
R4518 GND.n6011 GND.n1883 256.663
R4519 GND.n6011 GND.n1884 256.663
R4520 GND.n6011 GND.n1885 256.663
R4521 GND.n6011 GND.n1886 256.663
R4522 GND.n6011 GND.n1887 256.663
R4523 GND.n6011 GND.n1888 256.663
R4524 GND.n1890 GND.n1889 256.663
R4525 GND.n6011 GND.n1870 256.663
R4526 GND.n6011 GND.n1869 256.663
R4527 GND.n6011 GND.n1868 256.663
R4528 GND.n6011 GND.n1867 256.663
R4529 GND.n6011 GND.n1866 256.663
R4530 GND.n6011 GND.n1865 256.663
R4531 GND.n6011 GND.n1864 256.663
R4532 GND.n6011 GND.n1863 256.663
R4533 GND.n6011 GND.n1862 256.663
R4534 GND.n6011 GND.n1861 256.663
R4535 GND.n6011 GND.n1860 256.663
R4536 GND.n6011 GND.n1859 256.663
R4537 GND.n6011 GND.n1858 256.663
R4538 GND.n6011 GND.n1857 256.663
R4539 GND.n6011 GND.n1856 256.663
R4540 GND.n6011 GND.n1855 256.663
R4541 GND.n6011 GND.n1854 256.663
R4542 GND.n6011 GND.n1853 256.663
R4543 GND.n5588 GND.n2313 242.672
R4544 GND.n5588 GND.n2312 242.672
R4545 GND.n5588 GND.n2311 242.672
R4546 GND.n5588 GND.n2310 242.672
R4547 GND.n5588 GND.n2309 242.672
R4548 GND.n5589 GND.n5588 242.672
R4549 GND.n5588 GND.n2308 242.672
R4550 GND.n5588 GND.n2307 242.672
R4551 GND.n5588 GND.n2306 242.672
R4552 GND.n5291 GND.n154 242.672
R4553 GND.n5235 GND.n154 242.672
R4554 GND.n5281 GND.n154 242.672
R4555 GND.n5239 GND.n154 242.672
R4556 GND.n5271 GND.n154 242.672
R4557 GND.n5243 GND.n154 242.672
R4558 GND.n5261 GND.n154 242.672
R4559 GND.n5247 GND.n154 242.672
R4560 GND.n5251 GND.n154 242.672
R4561 GND.n4183 GND.n4182 242.672
R4562 GND.n4183 GND.n3047 242.672
R4563 GND.n4183 GND.n3048 242.672
R4564 GND.n4183 GND.n3049 242.672
R4565 GND.n4183 GND.n3050 242.672
R4566 GND.n4183 GND.n3051 242.672
R4567 GND.n4183 GND.n3052 242.672
R4568 GND.n4183 GND.n3053 242.672
R4569 GND.n4183 GND.n3054 242.672
R4570 GND.n4183 GND.n3055 242.672
R4571 GND.n4183 GND.n3056 242.672
R4572 GND.n4183 GND.n3057 242.672
R4573 GND.n4183 GND.n3058 242.672
R4574 GND.n5643 GND.n2220 242.672
R4575 GND.n5643 GND.n2221 242.672
R4576 GND.n5643 GND.n2222 242.672
R4577 GND.n5643 GND.n2223 242.672
R4578 GND.n5643 GND.n2224 242.672
R4579 GND.n5643 GND.n2225 242.672
R4580 GND.n5643 GND.n2226 242.672
R4581 GND.n5643 GND.n2227 242.672
R4582 GND.n5643 GND.n2228 242.672
R4583 GND.n5643 GND.n2229 242.672
R4584 GND.n5643 GND.n2230 242.672
R4585 GND.n5643 GND.n2231 242.672
R4586 GND.n5643 GND.n2232 242.672
R4587 GND.n6381 GND.n1327 242.672
R4588 GND.n6381 GND.n1328 242.672
R4589 GND.n6381 GND.n1329 242.672
R4590 GND.n6381 GND.n1330 242.672
R4591 GND.n6381 GND.n1331 242.672
R4592 GND.n6381 GND.n1332 242.672
R4593 GND.n6381 GND.n1333 242.672
R4594 GND.n6381 GND.n1334 242.672
R4595 GND.n6381 GND.n1335 242.672
R4596 GND.n6381 GND.n1336 242.672
R4597 GND.n6381 GND.n1337 242.672
R4598 GND.n6381 GND.n1338 242.672
R4599 GND.n6381 GND.n1339 242.672
R4600 GND.n6381 GND.n1340 242.672
R4601 GND.n6381 GND.n1341 242.672
R4602 GND.n6381 GND.n1342 242.672
R4603 GND.n6381 GND.n1343 242.672
R4604 GND.n6381 GND.n1344 242.672
R4605 GND.n6381 GND.n1345 242.672
R4606 GND.n6381 GND.n1346 242.672
R4607 GND.n6381 GND.n1347 242.672
R4608 GND.n6381 GND.n1348 242.672
R4609 GND.n6381 GND.n1349 242.672
R4610 GND.n6381 GND.n1350 242.672
R4611 GND.n6381 GND.n1351 242.672
R4612 GND.n6381 GND.n1352 242.672
R4613 GND.n6381 GND.n1353 242.672
R4614 GND.n6381 GND.n1354 242.672
R4615 GND.n6381 GND.n1355 242.672
R4616 GND.n6381 GND.n1356 242.672
R4617 GND.n6381 GND.n1357 242.672
R4618 GND.n6381 GND.n1358 242.672
R4619 GND.n6381 GND.n1359 242.672
R4620 GND.n6381 GND.n1360 242.672
R4621 GND.n6381 GND.n1361 242.672
R4622 GND.n6381 GND.n1362 242.672
R4623 GND.n6381 GND.n1363 242.672
R4624 GND.n6273 GND.n1485 242.672
R4625 GND.n6273 GND.n1484 242.672
R4626 GND.n6273 GND.n1483 242.672
R4627 GND.n6273 GND.n1482 242.672
R4628 GND.n6273 GND.n1481 242.672
R4629 GND.n6273 GND.n1480 242.672
R4630 GND.n6273 GND.n1479 242.672
R4631 GND.n6273 GND.n1478 242.672
R4632 GND.n6273 GND.n1477 242.672
R4633 GND.n6273 GND.n1476 242.672
R4634 GND.n6273 GND.n1475 242.672
R4635 GND.n6273 GND.n1474 242.672
R4636 GND.n6273 GND.n1473 242.672
R4637 GND.n6273 GND.n1472 242.672
R4638 GND.n6273 GND.n1471 242.672
R4639 GND.n6273 GND.n1470 242.672
R4640 GND.n6273 GND.n1469 242.672
R4641 GND.n6273 GND.n1468 242.672
R4642 GND.n6273 GND.n1467 242.672
R4643 GND.n6220 GND.n1572 242.672
R4644 GND.n6273 GND.n1496 242.672
R4645 GND.n6273 GND.n1497 242.672
R4646 GND.n6273 GND.n1498 242.672
R4647 GND.n6273 GND.n1499 242.672
R4648 GND.n6273 GND.n1500 242.672
R4649 GND.n6273 GND.n1501 242.672
R4650 GND.n6273 GND.n1502 242.672
R4651 GND.n6273 GND.n1503 242.672
R4652 GND.n6273 GND.n1504 242.672
R4653 GND.n6273 GND.n1505 242.672
R4654 GND.n6273 GND.n1506 242.672
R4655 GND.n6273 GND.n1507 242.672
R4656 GND.n6273 GND.n1508 242.672
R4657 GND.n6273 GND.n1509 242.672
R4658 GND.n6273 GND.n1510 242.672
R4659 GND.n6273 GND.n1511 242.672
R4660 GND.n6273 GND.n1512 242.672
R4661 GND.n5588 GND.n5587 242.672
R4662 GND.n5588 GND.n2269 242.672
R4663 GND.n5588 GND.n2270 242.672
R4664 GND.n5588 GND.n2271 242.672
R4665 GND.n5588 GND.n2272 242.672
R4666 GND.n5588 GND.n2273 242.672
R4667 GND.n5588 GND.n2274 242.672
R4668 GND.n5588 GND.n2275 242.672
R4669 GND.n5588 GND.n2276 242.672
R4670 GND.n5588 GND.n2277 242.672
R4671 GND.n5588 GND.n2278 242.672
R4672 GND.n5588 GND.n2279 242.672
R4673 GND.n5588 GND.n2280 242.672
R4674 GND.n5588 GND.n2281 242.672
R4675 GND.n5588 GND.n2282 242.672
R4676 GND.n5588 GND.n2283 242.672
R4677 GND.n5588 GND.n2284 242.672
R4678 GND.n5521 GND.n2354 242.672
R4679 GND.n5588 GND.n2285 242.672
R4680 GND.n5588 GND.n2286 242.672
R4681 GND.n5588 GND.n2287 242.672
R4682 GND.n5588 GND.n2288 242.672
R4683 GND.n5588 GND.n2289 242.672
R4684 GND.n5588 GND.n2290 242.672
R4685 GND.n5588 GND.n2291 242.672
R4686 GND.n5588 GND.n2292 242.672
R4687 GND.n5588 GND.n2293 242.672
R4688 GND.n5588 GND.n2294 242.672
R4689 GND.n5588 GND.n2295 242.672
R4690 GND.n5588 GND.n2296 242.672
R4691 GND.n5588 GND.n2297 242.672
R4692 GND.n5588 GND.n2298 242.672
R4693 GND.n5588 GND.n2299 242.672
R4694 GND.n5588 GND.n2300 242.672
R4695 GND.n5588 GND.n2301 242.672
R4696 GND.n5588 GND.n2302 242.672
R4697 GND.n5588 GND.n2303 242.672
R4698 GND.n288 GND.n154 242.672
R4699 GND.n7885 GND.n154 242.672
R4700 GND.n279 GND.n154 242.672
R4701 GND.n7892 GND.n154 242.672
R4702 GND.n272 GND.n154 242.672
R4703 GND.n7899 GND.n154 242.672
R4704 GND.n265 GND.n154 242.672
R4705 GND.n7906 GND.n154 242.672
R4706 GND.n258 GND.n154 242.672
R4707 GND.n7913 GND.n154 242.672
R4708 GND.n250 GND.n154 242.672
R4709 GND.n7920 GND.n154 242.672
R4710 GND.n241 GND.n154 242.672
R4711 GND.n7927 GND.n154 242.672
R4712 GND.n234 GND.n154 242.672
R4713 GND.n7934 GND.n154 242.672
R4714 GND.n227 GND.n154 242.672
R4715 GND.n7941 GND.n154 242.672
R4716 GND.n221 GND.n154 242.672
R4717 GND.n216 GND.n154 242.672
R4718 GND.n7952 GND.n154 242.672
R4719 GND.n208 GND.n154 242.672
R4720 GND.n7959 GND.n154 242.672
R4721 GND.n201 GND.n154 242.672
R4722 GND.n7966 GND.n154 242.672
R4723 GND.n194 GND.n154 242.672
R4724 GND.n7973 GND.n154 242.672
R4725 GND.n7976 GND.n154 242.672
R4726 GND.n185 GND.n154 242.672
R4727 GND.n7985 GND.n154 242.672
R4728 GND.n176 GND.n154 242.672
R4729 GND.n7992 GND.n154 242.672
R4730 GND.n169 GND.n154 242.672
R4731 GND.n7999 GND.n154 242.672
R4732 GND.n162 GND.n154 242.672
R4733 GND.n8006 GND.n154 242.672
R4734 GND.n8009 GND.n154 242.672
R4735 GND.n6381 GND.n1364 242.672
R4736 GND.n6381 GND.n1365 242.672
R4737 GND.n6381 GND.n1366 242.672
R4738 GND.n6381 GND.n1367 242.672
R4739 GND.n6381 GND.n1368 242.672
R4740 GND.n6381 GND.n1369 242.672
R4741 GND.n6381 GND.n1370 242.672
R4742 GND.n6381 GND.n1371 242.672
R4743 GND.n6273 GND.n1493 242.672
R4744 GND.n6273 GND.n1492 242.672
R4745 GND.n6273 GND.n1491 242.672
R4746 GND.n6273 GND.n1490 242.672
R4747 GND.n6273 GND.n1489 242.672
R4748 GND.n6273 GND.n1488 242.672
R4749 GND.n6273 GND.n1487 242.672
R4750 GND.n6273 GND.n1486 242.672
R4751 GND.n1460 GND.t135 242.326
R4752 GND.n1538 GND.t96 242.326
R4753 GND.n3193 GND.t93 242.326
R4754 GND.n3174 GND.t83 242.326
R4755 GND.n1569 GND.t157 242.326
R4756 GND.n2335 GND.t59 242.326
R4757 GND.n2356 GND.t120 242.326
R4758 GND.n2376 GND.t52 242.326
R4759 GND.n2396 GND.t80 242.326
R4760 GND.n284 GND.t66 242.326
R4761 GND.n247 GND.t70 242.326
R4762 GND.n214 GND.t138 242.326
R4763 GND.n181 GND.t73 242.326
R4764 GND.n5232 GND.t102 242.326
R4765 GND.n2663 GND.t123 242.326
R4766 GND.n3616 GND.t129 242.326
R4767 GND.n3665 GND.t62 242.326
R4768 GND.n3711 GND.t126 242.326
R4769 GND.n3538 GND.t99 242.326
R4770 GND.n6353 GND.t144 242.326
R4771 GND.n8008 GND.n8007 240.244
R4772 GND.n8005 GND.n156 240.244
R4773 GND.n8001 GND.n8000 240.244
R4774 GND.n7998 GND.n163 240.244
R4775 GND.n7994 GND.n7993 240.244
R4776 GND.n7991 GND.n170 240.244
R4777 GND.n7987 GND.n7986 240.244
R4778 GND.n7984 GND.n177 240.244
R4779 GND.n7977 GND.n186 240.244
R4780 GND.n7975 GND.n7974 240.244
R4781 GND.n7972 GND.n188 240.244
R4782 GND.n7968 GND.n7967 240.244
R4783 GND.n7965 GND.n195 240.244
R4784 GND.n7961 GND.n7960 240.244
R4785 GND.n7958 GND.n202 240.244
R4786 GND.n7954 GND.n7953 240.244
R4787 GND.n7951 GND.n209 240.244
R4788 GND.n220 GND.n217 240.244
R4789 GND.n7943 GND.n7942 240.244
R4790 GND.n7940 GND.n222 240.244
R4791 GND.n7936 GND.n7935 240.244
R4792 GND.n7933 GND.n228 240.244
R4793 GND.n7929 GND.n7928 240.244
R4794 GND.n7926 GND.n235 240.244
R4795 GND.n7922 GND.n7921 240.244
R4796 GND.n7919 GND.n242 240.244
R4797 GND.n7915 GND.n7914 240.244
R4798 GND.n7912 GND.n252 240.244
R4799 GND.n7908 GND.n7907 240.244
R4800 GND.n7905 GND.n259 240.244
R4801 GND.n7901 GND.n7900 240.244
R4802 GND.n7898 GND.n266 240.244
R4803 GND.n7894 GND.n7893 240.244
R4804 GND.n7891 GND.n273 240.244
R4805 GND.n7887 GND.n7886 240.244
R4806 GND.n7884 GND.n280 240.244
R4807 GND.n5440 GND.n2403 240.244
R4808 GND.n5049 GND.n2403 240.244
R4809 GND.n5049 GND.n2447 240.244
R4810 GND.n5059 GND.n2447 240.244
R4811 GND.n5059 GND.n2458 240.244
R4812 GND.n5064 GND.n2458 240.244
R4813 GND.n5064 GND.n2468 240.244
R4814 GND.n5074 GND.n2468 240.244
R4815 GND.n5074 GND.n2478 240.244
R4816 GND.n5079 GND.n2478 240.244
R4817 GND.n5079 GND.n2489 240.244
R4818 GND.n5089 GND.n2489 240.244
R4819 GND.n5089 GND.n2499 240.244
R4820 GND.n5094 GND.n2499 240.244
R4821 GND.n5094 GND.n2510 240.244
R4822 GND.n5104 GND.n2510 240.244
R4823 GND.n5104 GND.n2520 240.244
R4824 GND.n5109 GND.n2520 240.244
R4825 GND.n5109 GND.n2529 240.244
R4826 GND.n5123 GND.n2529 240.244
R4827 GND.n5123 GND.n2539 240.244
R4828 GND.n2543 GND.n2539 240.244
R4829 GND.n2560 GND.n2543 240.244
R4830 GND.n2560 GND.n33 240.244
R4831 GND.n5134 GND.n33 240.244
R4832 GND.n5134 GND.n2553 240.244
R4833 GND.n5355 GND.n2553 240.244
R4834 GND.n5355 GND.n52 240.244
R4835 GND.n5347 GND.n52 240.244
R4836 GND.n5347 GND.n63 240.244
R4837 GND.n5343 GND.n63 240.244
R4838 GND.n5343 GND.n73 240.244
R4839 GND.n5335 GND.n73 240.244
R4840 GND.n5335 GND.n83 240.244
R4841 GND.n5331 GND.n83 240.244
R4842 GND.n5331 GND.n94 240.244
R4843 GND.n5323 GND.n94 240.244
R4844 GND.n5323 GND.n104 240.244
R4845 GND.n5319 GND.n104 240.244
R4846 GND.n5319 GND.n115 240.244
R4847 GND.n5311 GND.n115 240.244
R4848 GND.n5311 GND.n125 240.244
R4849 GND.n5307 GND.n125 240.244
R4850 GND.n5307 GND.n136 240.244
R4851 GND.n5299 GND.n136 240.244
R4852 GND.n5299 GND.n146 240.244
R4853 GND.n7876 GND.n146 240.244
R4854 GND.n2315 GND.n2314 240.244
R4855 GND.n5581 GND.n2314 240.244
R4856 GND.n5579 GND.n5578 240.244
R4857 GND.n5575 GND.n5574 240.244
R4858 GND.n5571 GND.n5570 240.244
R4859 GND.n5567 GND.n5566 240.244
R4860 GND.n5563 GND.n5562 240.244
R4861 GND.n5559 GND.n5558 240.244
R4862 GND.n5554 GND.n2333 240.244
R4863 GND.n5552 GND.n5551 240.244
R4864 GND.n5548 GND.n5547 240.244
R4865 GND.n5544 GND.n5543 240.244
R4866 GND.n5540 GND.n5539 240.244
R4867 GND.n5536 GND.n5535 240.244
R4868 GND.n5532 GND.n5531 240.244
R4869 GND.n5528 GND.n5527 240.244
R4870 GND.n5524 GND.n5523 240.244
R4871 GND.n5519 GND.n5518 240.244
R4872 GND.n5515 GND.n5514 240.244
R4873 GND.n5511 GND.n5510 240.244
R4874 GND.n5507 GND.n5506 240.244
R4875 GND.n5503 GND.n5502 240.244
R4876 GND.n5499 GND.n5498 240.244
R4877 GND.n5495 GND.n5494 240.244
R4878 GND.n5491 GND.n5490 240.244
R4879 GND.n5487 GND.n5486 240.244
R4880 GND.n5482 GND.n5481 240.244
R4881 GND.n5478 GND.n5477 240.244
R4882 GND.n5474 GND.n5473 240.244
R4883 GND.n5470 GND.n5469 240.244
R4884 GND.n5466 GND.n5465 240.244
R4885 GND.n5462 GND.n5461 240.244
R4886 GND.n5458 GND.n5457 240.244
R4887 GND.n5454 GND.n5453 240.244
R4888 GND.n5450 GND.n5449 240.244
R4889 GND.n2395 GND.n2304 240.244
R4890 GND.n5435 GND.n2316 240.244
R4891 GND.n5435 GND.n2438 240.244
R4892 GND.n5431 GND.n2438 240.244
R4893 GND.n5431 GND.n2445 240.244
R4894 GND.n5423 GND.n2445 240.244
R4895 GND.n5423 GND.n2460 240.244
R4896 GND.n5419 GND.n2460 240.244
R4897 GND.n5419 GND.n2466 240.244
R4898 GND.n5411 GND.n2466 240.244
R4899 GND.n5411 GND.n2481 240.244
R4900 GND.n5407 GND.n2481 240.244
R4901 GND.n5407 GND.n2487 240.244
R4902 GND.n5399 GND.n2487 240.244
R4903 GND.n5399 GND.n2502 240.244
R4904 GND.n5395 GND.n2502 240.244
R4905 GND.n5395 GND.n2508 240.244
R4906 GND.n5387 GND.n2508 240.244
R4907 GND.n5387 GND.n2523 240.244
R4908 GND.n5383 GND.n2523 240.244
R4909 GND.n5383 GND.n2527 240.244
R4910 GND.n5375 GND.n2527 240.244
R4911 GND.n5375 GND.n5374 240.244
R4912 GND.n5374 GND.n36 240.244
R4913 GND.n8077 GND.n36 240.244
R4914 GND.n8077 GND.n37 240.244
R4915 GND.n5362 GND.n37 240.244
R4916 GND.n5362 GND.n49 240.244
R4917 GND.n8072 GND.n49 240.244
R4918 GND.n8072 GND.n50 240.244
R4919 GND.n8064 GND.n50 240.244
R4920 GND.n8064 GND.n66 240.244
R4921 GND.n8060 GND.n66 240.244
R4922 GND.n8060 GND.n71 240.244
R4923 GND.n8052 GND.n71 240.244
R4924 GND.n8052 GND.n86 240.244
R4925 GND.n8048 GND.n86 240.244
R4926 GND.n8048 GND.n92 240.244
R4927 GND.n8040 GND.n92 240.244
R4928 GND.n8040 GND.n107 240.244
R4929 GND.n8036 GND.n107 240.244
R4930 GND.n8036 GND.n113 240.244
R4931 GND.n8028 GND.n113 240.244
R4932 GND.n8028 GND.n128 240.244
R4933 GND.n8024 GND.n128 240.244
R4934 GND.n8024 GND.n134 240.244
R4935 GND.n8016 GND.n134 240.244
R4936 GND.n8016 GND.n149 240.244
R4937 GND.n6272 GND.n1514 240.244
R4938 GND.n1519 GND.n1518 240.244
R4939 GND.n1521 GND.n1520 240.244
R4940 GND.n1525 GND.n1524 240.244
R4941 GND.n1527 GND.n1526 240.244
R4942 GND.n1531 GND.n1530 240.244
R4943 GND.n1533 GND.n1532 240.244
R4944 GND.n1537 GND.n1536 240.244
R4945 GND.n1542 GND.n1541 240.244
R4946 GND.n1546 GND.n1545 240.244
R4947 GND.n1548 GND.n1547 240.244
R4948 GND.n1552 GND.n1551 240.244
R4949 GND.n1554 GND.n1553 240.244
R4950 GND.n1558 GND.n1557 240.244
R4951 GND.n1560 GND.n1559 240.244
R4952 GND.n1564 GND.n1563 240.244
R4953 GND.n6221 GND.n1565 240.244
R4954 GND.n1567 GND.n1466 240.244
R4955 GND.n3215 GND.n3214 240.244
R4956 GND.n3210 GND.n3209 240.244
R4957 GND.n3223 GND.n3222 240.244
R4958 GND.n3206 GND.n3205 240.244
R4959 GND.n3231 GND.n3230 240.244
R4960 GND.n3202 GND.n3201 240.244
R4961 GND.n3239 GND.n3238 240.244
R4962 GND.n3198 GND.n3197 240.244
R4963 GND.n3247 GND.n3246 240.244
R4964 GND.n3191 GND.n3190 240.244
R4965 GND.n3255 GND.n3254 240.244
R4966 GND.n3187 GND.n3186 240.244
R4967 GND.n3263 GND.n3262 240.244
R4968 GND.n3183 GND.n3182 240.244
R4969 GND.n3271 GND.n3270 240.244
R4970 GND.n3179 GND.n3178 240.244
R4971 GND.n3279 GND.n3278 240.244
R4972 GND.n3285 GND.n3284 240.244
R4973 GND.n3777 GND.n3534 240.244
R4974 GND.n3534 GND.n3517 240.244
R4975 GND.n3517 GND.n3507 240.244
R4976 GND.n3802 GND.n3507 240.244
R4977 GND.n3802 GND.n3498 240.244
R4978 GND.n3804 GND.n3498 240.244
R4979 GND.n3804 GND.n3487 240.244
R4980 GND.n3487 GND.n3478 240.244
R4981 GND.n3839 GND.n3478 240.244
R4982 GND.n3839 GND.n3469 240.244
R4983 GND.n3841 GND.n3469 240.244
R4984 GND.n3841 GND.n3459 240.244
R4985 GND.n3459 GND.n3449 240.244
R4986 GND.n3882 GND.n3449 240.244
R4987 GND.n3882 GND.n3440 240.244
R4988 GND.n3885 GND.n3440 240.244
R4989 GND.n3885 GND.n3432 240.244
R4990 GND.n3432 GND.n3431 240.244
R4991 GND.n3431 GND.n3408 240.244
R4992 GND.n3910 GND.n3408 240.244
R4993 GND.n3910 GND.n3418 240.244
R4994 GND.n3912 GND.n3418 240.244
R4995 GND.n3913 GND.n3912 240.244
R4996 GND.n3935 GND.n3913 240.244
R4997 GND.n3935 GND.n3919 240.244
R4998 GND.n3969 GND.n3919 240.244
R4999 GND.n3969 GND.n3394 240.244
R5000 GND.n3999 GND.n3394 240.244
R5001 GND.n3999 GND.n3385 240.244
R5002 GND.n4001 GND.n3385 240.244
R5003 GND.n4001 GND.n3375 240.244
R5004 GND.n3375 GND.n3366 240.244
R5005 GND.n4036 GND.n3366 240.244
R5006 GND.n4036 GND.n3357 240.244
R5007 GND.n4038 GND.n3357 240.244
R5008 GND.n4038 GND.n3347 240.244
R5009 GND.n3347 GND.n3337 240.244
R5010 GND.n4073 GND.n3337 240.244
R5011 GND.n4073 GND.n3327 240.244
R5012 GND.n4075 GND.n3327 240.244
R5013 GND.n4075 GND.n3317 240.244
R5014 GND.n3317 GND.n3308 240.244
R5015 GND.n4133 GND.n3308 240.244
R5016 GND.n4133 GND.n3300 240.244
R5017 GND.n4136 GND.n3300 240.244
R5018 GND.n4136 GND.n3172 240.244
R5019 GND.n4155 GND.n3172 240.244
R5020 GND.n3578 GND.n3577 240.244
R5021 GND.n3585 GND.n3584 240.244
R5022 GND.n3588 GND.n3587 240.244
R5023 GND.n3595 GND.n3594 240.244
R5024 GND.n3598 GND.n3597 240.244
R5025 GND.n3605 GND.n3604 240.244
R5026 GND.n3608 GND.n3607 240.244
R5027 GND.n3615 GND.n3614 240.244
R5028 GND.n3620 GND.n3619 240.244
R5029 GND.n3627 GND.n3626 240.244
R5030 GND.n3630 GND.n3629 240.244
R5031 GND.n3637 GND.n3636 240.244
R5032 GND.n3640 GND.n3639 240.244
R5033 GND.n3647 GND.n3646 240.244
R5034 GND.n3650 GND.n3649 240.244
R5035 GND.n3657 GND.n3656 240.244
R5036 GND.n3660 GND.n3659 240.244
R5037 GND.n3669 GND.n3668 240.244
R5038 GND.n3672 GND.n3671 240.244
R5039 GND.n3679 GND.n3678 240.244
R5040 GND.n3682 GND.n3681 240.244
R5041 GND.n3689 GND.n3688 240.244
R5042 GND.n3692 GND.n3691 240.244
R5043 GND.n3699 GND.n3698 240.244
R5044 GND.n3702 GND.n3701 240.244
R5045 GND.n3709 GND.n3708 240.244
R5046 GND.n3715 GND.n3714 240.244
R5047 GND.n3722 GND.n3721 240.244
R5048 GND.n3725 GND.n3724 240.244
R5049 GND.n3732 GND.n3731 240.244
R5050 GND.n3735 GND.n3734 240.244
R5051 GND.n3742 GND.n3741 240.244
R5052 GND.n3745 GND.n3744 240.244
R5053 GND.n3752 GND.n3751 240.244
R5054 GND.n3755 GND.n3754 240.244
R5055 GND.n3541 GND.n3537 240.244
R5056 GND.n3780 GND.n3520 240.244
R5057 GND.n3788 GND.n3520 240.244
R5058 GND.n3788 GND.n3521 240.244
R5059 GND.n3521 GND.n3496 240.244
R5060 GND.n3817 GND.n3496 240.244
R5061 GND.n3817 GND.n3491 240.244
R5062 GND.n3825 GND.n3491 240.244
R5063 GND.n3825 GND.n3492 240.244
R5064 GND.n3492 GND.n3467 240.244
R5065 GND.n3854 GND.n3467 240.244
R5066 GND.n3854 GND.n3462 240.244
R5067 GND.n3862 GND.n3462 240.244
R5068 GND.n3862 GND.n3463 240.244
R5069 GND.n3463 GND.n3438 240.244
R5070 GND.n3894 GND.n3438 240.244
R5071 GND.n3894 GND.n3434 240.244
R5072 GND.n3901 GND.n3434 240.244
R5073 GND.n3901 GND.n3412 240.244
R5074 GND.n3987 GND.n3412 240.244
R5075 GND.n3987 GND.n3413 240.244
R5076 GND.n3982 GND.n3413 240.244
R5077 GND.n3982 GND.n3416 240.244
R5078 GND.n3933 GND.n3416 240.244
R5079 GND.n3960 GND.n3933 240.244
R5080 GND.n3960 GND.n3923 240.244
R5081 GND.n3967 GND.n3923 240.244
R5082 GND.n3967 GND.n3930 240.244
R5083 GND.n3930 GND.n3384 240.244
R5084 GND.n4014 GND.n3384 240.244
R5085 GND.n4014 GND.n3379 240.244
R5086 GND.n4022 GND.n3379 240.244
R5087 GND.n4022 GND.n3380 240.244
R5088 GND.n3380 GND.n3355 240.244
R5089 GND.n4051 GND.n3355 240.244
R5090 GND.n4051 GND.n3350 240.244
R5091 GND.n4059 GND.n3350 240.244
R5092 GND.n4059 GND.n3351 240.244
R5093 GND.n3351 GND.n3325 240.244
R5094 GND.n4088 GND.n3325 240.244
R5095 GND.n4088 GND.n3320 240.244
R5096 GND.n4096 GND.n3320 240.244
R5097 GND.n4096 GND.n3321 240.244
R5098 GND.n3321 GND.n3298 240.244
R5099 GND.n4143 GND.n3298 240.244
R5100 GND.n4143 GND.n3294 240.244
R5101 GND.n4150 GND.n3294 240.244
R5102 GND.n4150 GND.n1513 240.244
R5103 GND.n5642 GND.n2234 240.244
R5104 GND.n5635 GND.n5634 240.244
R5105 GND.n5632 GND.n5631 240.244
R5106 GND.n5628 GND.n5627 240.244
R5107 GND.n5624 GND.n5623 240.244
R5108 GND.n5620 GND.n5619 240.244
R5109 GND.n5616 GND.n5615 240.244
R5110 GND.n5612 GND.n5611 240.244
R5111 GND.n5608 GND.n5607 240.244
R5112 GND.n5604 GND.n5603 240.244
R5113 GND.n5600 GND.n5599 240.244
R5114 GND.n5596 GND.n5595 240.244
R5115 GND.n5026 GND.n5025 240.244
R5116 GND.n3038 GND.n3029 240.244
R5117 GND.n4206 GND.n3029 240.244
R5118 GND.n4206 GND.n3025 240.244
R5119 GND.n4214 GND.n3025 240.244
R5120 GND.n4214 GND.n3016 240.244
R5121 GND.n3016 GND.n3006 240.244
R5122 GND.n4238 GND.n3006 240.244
R5123 GND.n4238 GND.n3002 240.244
R5124 GND.n4246 GND.n3002 240.244
R5125 GND.n4246 GND.n2993 240.244
R5126 GND.n2993 GND.n2983 240.244
R5127 GND.n4270 GND.n2983 240.244
R5128 GND.n4270 GND.n2979 240.244
R5129 GND.n4278 GND.n2979 240.244
R5130 GND.n4278 GND.n2970 240.244
R5131 GND.n2970 GND.n2960 240.244
R5132 GND.n4302 GND.n2960 240.244
R5133 GND.n4302 GND.n2956 240.244
R5134 GND.n4310 GND.n2956 240.244
R5135 GND.n4310 GND.n2947 240.244
R5136 GND.n2947 GND.n2936 240.244
R5137 GND.n4334 GND.n2936 240.244
R5138 GND.n4334 GND.n2932 240.244
R5139 GND.n4342 GND.n2932 240.244
R5140 GND.n4342 GND.n2924 240.244
R5141 GND.n2924 GND.n2914 240.244
R5142 GND.n4366 GND.n2914 240.244
R5143 GND.n4366 GND.n2910 240.244
R5144 GND.n4374 GND.n2910 240.244
R5145 GND.n4374 GND.n2901 240.244
R5146 GND.n2901 GND.n2891 240.244
R5147 GND.n4398 GND.n2891 240.244
R5148 GND.n4398 GND.n2887 240.244
R5149 GND.n4406 GND.n2887 240.244
R5150 GND.n4406 GND.n2878 240.244
R5151 GND.n2878 GND.n2868 240.244
R5152 GND.n4430 GND.n2868 240.244
R5153 GND.n4430 GND.n2864 240.244
R5154 GND.n4438 GND.n2864 240.244
R5155 GND.n4438 GND.n2855 240.244
R5156 GND.n2855 GND.n2845 240.244
R5157 GND.n4462 GND.n2845 240.244
R5158 GND.n4462 GND.n2841 240.244
R5159 GND.n4470 GND.n2841 240.244
R5160 GND.n4470 GND.n2832 240.244
R5161 GND.n2832 GND.n2822 240.244
R5162 GND.n4494 GND.n2822 240.244
R5163 GND.n4494 GND.n2818 240.244
R5164 GND.n4502 GND.n2818 240.244
R5165 GND.n4502 GND.n2809 240.244
R5166 GND.n2809 GND.n2799 240.244
R5167 GND.n4526 GND.n2799 240.244
R5168 GND.n4526 GND.n2795 240.244
R5169 GND.n4537 GND.n2795 240.244
R5170 GND.n4537 GND.n2786 240.244
R5171 GND.n2786 GND.n2775 240.244
R5172 GND.n4578 GND.n2775 240.244
R5173 GND.n4579 GND.n4578 240.244
R5174 GND.n4654 GND.n4579 240.244
R5175 GND.n4654 GND.n1651 240.244
R5176 GND.n4665 GND.n1651 240.244
R5177 GND.n4665 GND.n1662 240.244
R5178 GND.n4661 GND.n1662 240.244
R5179 GND.n4661 GND.n2764 240.244
R5180 GND.n4692 GND.n2764 240.244
R5181 GND.n4692 GND.n1681 240.244
R5182 GND.n4713 GND.n1681 240.244
R5183 GND.n4713 GND.n1697 240.244
R5184 GND.n4709 GND.n1697 240.244
R5185 GND.n4709 GND.n4708 240.244
R5186 GND.n4708 GND.n4707 240.244
R5187 GND.n4707 GND.n4700 240.244
R5188 GND.n4700 GND.n1730 240.244
R5189 GND.n4764 GND.n1730 240.244
R5190 GND.n4764 GND.n1749 240.244
R5191 GND.n2747 GND.n1749 240.244
R5192 GND.n4771 GND.n2747 240.244
R5193 GND.n4772 GND.n4771 240.244
R5194 GND.n4773 GND.n4772 240.244
R5195 GND.n4773 GND.n2742 240.244
R5196 GND.n4788 GND.n2742 240.244
R5197 GND.n4788 GND.n2743 240.244
R5198 GND.n4784 GND.n2743 240.244
R5199 GND.n4784 GND.n2736 240.244
R5200 GND.n2736 GND.n2728 240.244
R5201 GND.n4857 GND.n2728 240.244
R5202 GND.n4858 GND.n4857 240.244
R5203 GND.n4858 GND.n2724 240.244
R5204 GND.n4867 GND.n2724 240.244
R5205 GND.n4867 GND.n2711 240.244
R5206 GND.n4878 GND.n2711 240.244
R5207 GND.n4880 GND.n4878 240.244
R5208 GND.n4880 GND.n1897 240.244
R5209 GND.n2707 GND.n1897 240.244
R5210 GND.n4887 GND.n2707 240.244
R5211 GND.n4888 GND.n4887 240.244
R5212 GND.n4890 GND.n4888 240.244
R5213 GND.n4890 GND.n4889 240.244
R5214 GND.n4889 GND.n1913 240.244
R5215 GND.n4897 GND.n1913 240.244
R5216 GND.n4898 GND.n4897 240.244
R5217 GND.n4898 GND.n1924 240.244
R5218 GND.n4904 GND.n1924 240.244
R5219 GND.n4904 GND.n1937 240.244
R5220 GND.n4908 GND.n1937 240.244
R5221 GND.n4908 GND.n4907 240.244
R5222 GND.n4907 GND.n1951 240.244
R5223 GND.n4915 GND.n1951 240.244
R5224 GND.n4915 GND.n1964 240.244
R5225 GND.n4921 GND.n1964 240.244
R5226 GND.n4922 GND.n4921 240.244
R5227 GND.n4922 GND.n1978 240.244
R5228 GND.n4926 GND.n1978 240.244
R5229 GND.n4926 GND.n1991 240.244
R5230 GND.n4932 GND.n1991 240.244
R5231 GND.n4933 GND.n4932 240.244
R5232 GND.n4933 GND.n2005 240.244
R5233 GND.n2693 GND.n2005 240.244
R5234 GND.n2693 GND.n2017 240.244
R5235 GND.n4941 GND.n2017 240.244
R5236 GND.n4942 GND.n4941 240.244
R5237 GND.n4942 GND.n2031 240.244
R5238 GND.n4948 GND.n2031 240.244
R5239 GND.n4948 GND.n2044 240.244
R5240 GND.n4952 GND.n2044 240.244
R5241 GND.n4952 GND.n4951 240.244
R5242 GND.n4951 GND.n2058 240.244
R5243 GND.n4959 GND.n2058 240.244
R5244 GND.n4959 GND.n2071 240.244
R5245 GND.n4965 GND.n2071 240.244
R5246 GND.n4966 GND.n4965 240.244
R5247 GND.n4966 GND.n2085 240.244
R5248 GND.n4970 GND.n2085 240.244
R5249 GND.n4970 GND.n2098 240.244
R5250 GND.n4976 GND.n2098 240.244
R5251 GND.n4977 GND.n4976 240.244
R5252 GND.n4977 GND.n2112 240.244
R5253 GND.n2680 GND.n2112 240.244
R5254 GND.n2680 GND.n2125 240.244
R5255 GND.n4985 GND.n2125 240.244
R5256 GND.n4986 GND.n4985 240.244
R5257 GND.n4986 GND.n2139 240.244
R5258 GND.n4992 GND.n2139 240.244
R5259 GND.n4992 GND.n2152 240.244
R5260 GND.n4996 GND.n2152 240.244
R5261 GND.n4996 GND.n4995 240.244
R5262 GND.n4995 GND.n2166 240.244
R5263 GND.n5004 GND.n2166 240.244
R5264 GND.n5004 GND.n2178 240.244
R5265 GND.n5010 GND.n2178 240.244
R5266 GND.n5011 GND.n5010 240.244
R5267 GND.n5011 GND.n2192 240.244
R5268 GND.n5015 GND.n2192 240.244
R5269 GND.n5015 GND.n2205 240.244
R5270 GND.n2670 GND.n2205 240.244
R5271 GND.n5022 GND.n2670 240.244
R5272 GND.n4181 GND.n3059 240.244
R5273 GND.n4177 GND.n3059 240.244
R5274 GND.n4175 GND.n4174 240.244
R5275 GND.n4171 GND.n4170 240.244
R5276 GND.n4167 GND.n4166 240.244
R5277 GND.n4163 GND.n4162 240.244
R5278 GND.n3074 GND.n3073 240.244
R5279 GND.n3076 GND.n3075 240.244
R5280 GND.n3086 GND.n3085 240.244
R5281 GND.n3094 GND.n3093 240.244
R5282 GND.n3096 GND.n3095 240.244
R5283 GND.n3137 GND.n3105 240.244
R5284 GND.n3113 GND.n3112 240.244
R5285 GND.n4196 GND.n3032 240.244
R5286 GND.n4204 GND.n3032 240.244
R5287 GND.n4204 GND.n3033 240.244
R5288 GND.n3033 GND.n3014 240.244
R5289 GND.n4228 GND.n3014 240.244
R5290 GND.n4228 GND.n3009 240.244
R5291 GND.n4236 GND.n3009 240.244
R5292 GND.n4236 GND.n3010 240.244
R5293 GND.n3010 GND.n2991 240.244
R5294 GND.n4260 GND.n2991 240.244
R5295 GND.n4260 GND.n2986 240.244
R5296 GND.n4268 GND.n2986 240.244
R5297 GND.n4268 GND.n2987 240.244
R5298 GND.n2987 GND.n2968 240.244
R5299 GND.n4292 GND.n2968 240.244
R5300 GND.n4292 GND.n2963 240.244
R5301 GND.n4300 GND.n2963 240.244
R5302 GND.n4300 GND.n2964 240.244
R5303 GND.n2964 GND.n2945 240.244
R5304 GND.n4324 GND.n2945 240.244
R5305 GND.n4324 GND.n2939 240.244
R5306 GND.n4332 GND.n2939 240.244
R5307 GND.n4332 GND.n2941 240.244
R5308 GND.n2941 GND.n2922 240.244
R5309 GND.n4356 GND.n2922 240.244
R5310 GND.n4356 GND.n2917 240.244
R5311 GND.n4364 GND.n2917 240.244
R5312 GND.n4364 GND.n2918 240.244
R5313 GND.n2918 GND.n2899 240.244
R5314 GND.n4388 GND.n2899 240.244
R5315 GND.n4388 GND.n2894 240.244
R5316 GND.n4396 GND.n2894 240.244
R5317 GND.n4396 GND.n2895 240.244
R5318 GND.n2895 GND.n2876 240.244
R5319 GND.n4420 GND.n2876 240.244
R5320 GND.n4420 GND.n2871 240.244
R5321 GND.n4428 GND.n2871 240.244
R5322 GND.n4428 GND.n2872 240.244
R5323 GND.n2872 GND.n2853 240.244
R5324 GND.n4452 GND.n2853 240.244
R5325 GND.n4452 GND.n2848 240.244
R5326 GND.n4460 GND.n2848 240.244
R5327 GND.n4460 GND.n2849 240.244
R5328 GND.n2849 GND.n2830 240.244
R5329 GND.n4484 GND.n2830 240.244
R5330 GND.n4484 GND.n2825 240.244
R5331 GND.n4492 GND.n2825 240.244
R5332 GND.n4492 GND.n2826 240.244
R5333 GND.n2826 GND.n2807 240.244
R5334 GND.n4516 GND.n2807 240.244
R5335 GND.n4516 GND.n2802 240.244
R5336 GND.n4524 GND.n2802 240.244
R5337 GND.n4524 GND.n2803 240.244
R5338 GND.n2803 GND.n2784 240.244
R5339 GND.n4567 GND.n2784 240.244
R5340 GND.n4567 GND.n2779 240.244
R5341 GND.n4576 GND.n2779 240.244
R5342 GND.n4576 GND.n2780 240.244
R5343 GND.n2780 GND.n1653 240.244
R5344 GND.n6142 GND.n1653 240.244
R5345 GND.n6142 GND.n1654 240.244
R5346 GND.n6138 GND.n1654 240.244
R5347 GND.n6138 GND.n1660 240.244
R5348 GND.n1687 GND.n1660 240.244
R5349 GND.n1687 GND.n1683 240.244
R5350 GND.n6121 GND.n1683 240.244
R5351 GND.n6121 GND.n1684 240.244
R5352 GND.n6117 GND.n1684 240.244
R5353 GND.n6117 GND.n1695 240.244
R5354 GND.n1738 GND.n1695 240.244
R5355 GND.n1739 GND.n1738 240.244
R5356 GND.n1739 GND.n1732 240.244
R5357 GND.n6094 GND.n1732 240.244
R5358 GND.n6094 GND.n1733 240.244
R5359 GND.n6090 GND.n1733 240.244
R5360 GND.n6090 GND.n1747 240.244
R5361 GND.n4797 GND.n1747 240.244
R5362 GND.n4798 GND.n4797 240.244
R5363 GND.n4799 GND.n4798 240.244
R5364 GND.n4799 GND.n4789 240.244
R5365 GND.n4807 GND.n4789 240.244
R5366 GND.n4807 GND.n4790 240.244
R5367 GND.n4790 GND.n2735 240.244
R5368 GND.n4847 GND.n2735 240.244
R5369 GND.n4847 GND.n2730 240.244
R5370 GND.n4855 GND.n2730 240.244
R5371 GND.n4855 GND.n2731 240.244
R5372 GND.n2731 GND.n2718 240.244
R5373 GND.n4869 GND.n2718 240.244
R5374 GND.n4869 GND.n2714 240.244
R5375 GND.n4876 GND.n2714 240.244
R5376 GND.n4876 GND.n1898 240.244
R5377 GND.n5817 GND.n1898 240.244
R5378 GND.n5817 GND.n1899 240.244
R5379 GND.n5813 GND.n1899 240.244
R5380 GND.n5813 GND.n5812 240.244
R5381 GND.n5812 GND.n5811 240.244
R5382 GND.n5811 GND.n1905 240.244
R5383 GND.n5807 GND.n1905 240.244
R5384 GND.n5807 GND.n1911 240.244
R5385 GND.n1926 GND.n1911 240.244
R5386 GND.n5797 GND.n1926 240.244
R5387 GND.n5797 GND.n1927 240.244
R5388 GND.n5793 GND.n1927 240.244
R5389 GND.n5793 GND.n1935 240.244
R5390 GND.n1953 GND.n1935 240.244
R5391 GND.n5783 GND.n1953 240.244
R5392 GND.n5783 GND.n1954 240.244
R5393 GND.n5779 GND.n1954 240.244
R5394 GND.n5779 GND.n1962 240.244
R5395 GND.n1980 GND.n1962 240.244
R5396 GND.n5769 GND.n1980 240.244
R5397 GND.n5769 GND.n1981 240.244
R5398 GND.n5765 GND.n1981 240.244
R5399 GND.n5765 GND.n1989 240.244
R5400 GND.n2006 GND.n1989 240.244
R5401 GND.n5755 GND.n2006 240.244
R5402 GND.n5755 GND.n2007 240.244
R5403 GND.n5751 GND.n2007 240.244
R5404 GND.n5751 GND.n2015 240.244
R5405 GND.n2033 GND.n2015 240.244
R5406 GND.n5741 GND.n2033 240.244
R5407 GND.n5741 GND.n2034 240.244
R5408 GND.n5737 GND.n2034 240.244
R5409 GND.n5737 GND.n2042 240.244
R5410 GND.n2060 GND.n2042 240.244
R5411 GND.n5727 GND.n2060 240.244
R5412 GND.n5727 GND.n2061 240.244
R5413 GND.n5723 GND.n2061 240.244
R5414 GND.n5723 GND.n2069 240.244
R5415 GND.n2087 GND.n2069 240.244
R5416 GND.n5713 GND.n2087 240.244
R5417 GND.n5713 GND.n2088 240.244
R5418 GND.n5709 GND.n2088 240.244
R5419 GND.n5709 GND.n2096 240.244
R5420 GND.n2114 GND.n2096 240.244
R5421 GND.n5699 GND.n2114 240.244
R5422 GND.n5699 GND.n2115 240.244
R5423 GND.n5695 GND.n2115 240.244
R5424 GND.n5695 GND.n2123 240.244
R5425 GND.n2141 GND.n2123 240.244
R5426 GND.n5685 GND.n2141 240.244
R5427 GND.n5685 GND.n2142 240.244
R5428 GND.n5681 GND.n2142 240.244
R5429 GND.n5681 GND.n2150 240.244
R5430 GND.n2168 GND.n2150 240.244
R5431 GND.n5671 GND.n2168 240.244
R5432 GND.n5671 GND.n2169 240.244
R5433 GND.n5667 GND.n2169 240.244
R5434 GND.n5667 GND.n2177 240.244
R5435 GND.n2194 GND.n2177 240.244
R5436 GND.n5657 GND.n2194 240.244
R5437 GND.n5657 GND.n2195 240.244
R5438 GND.n5653 GND.n2195 240.244
R5439 GND.n5653 GND.n2203 240.244
R5440 GND.n2233 GND.n2203 240.244
R5441 GND.n5253 GND.n5252 240.244
R5442 GND.n5260 GND.n5259 240.244
R5443 GND.n5263 GND.n5262 240.244
R5444 GND.n5270 GND.n5269 240.244
R5445 GND.n5273 GND.n5272 240.244
R5446 GND.n5280 GND.n5279 240.244
R5447 GND.n5283 GND.n5282 240.244
R5448 GND.n5290 GND.n5289 240.244
R5449 GND.n2436 GND.n2405 240.244
R5450 GND.n5051 GND.n2436 240.244
R5451 GND.n5051 GND.n2448 240.244
R5452 GND.n5057 GND.n2448 240.244
R5453 GND.n5057 GND.n2459 240.244
R5454 GND.n5066 GND.n2459 240.244
R5455 GND.n5066 GND.n2469 240.244
R5456 GND.n5072 GND.n2469 240.244
R5457 GND.n5072 GND.n2479 240.244
R5458 GND.n5081 GND.n2479 240.244
R5459 GND.n5081 GND.n2490 240.244
R5460 GND.n5087 GND.n2490 240.244
R5461 GND.n5087 GND.n2500 240.244
R5462 GND.n5096 GND.n2500 240.244
R5463 GND.n5096 GND.n2511 240.244
R5464 GND.n5102 GND.n2511 240.244
R5465 GND.n5102 GND.n2521 240.244
R5466 GND.n5111 GND.n2521 240.244
R5467 GND.n5111 GND.n2530 240.244
R5468 GND.n5121 GND.n2530 240.244
R5469 GND.n5121 GND.n2540 240.244
R5470 GND.n2544 GND.n2540 240.244
R5471 GND.n2544 GND.n30 240.244
R5472 GND.n8079 GND.n30 240.244
R5473 GND.n8079 GND.n31 240.244
R5474 GND.n2554 GND.n31 240.244
R5475 GND.n5353 GND.n2554 240.244
R5476 GND.n5353 GND.n53 240.244
R5477 GND.n5349 GND.n53 240.244
R5478 GND.n5349 GND.n64 240.244
R5479 GND.n5341 GND.n64 240.244
R5480 GND.n5341 GND.n74 240.244
R5481 GND.n5337 GND.n74 240.244
R5482 GND.n5337 GND.n84 240.244
R5483 GND.n5329 GND.n84 240.244
R5484 GND.n5329 GND.n95 240.244
R5485 GND.n5325 GND.n95 240.244
R5486 GND.n5325 GND.n105 240.244
R5487 GND.n5317 GND.n105 240.244
R5488 GND.n5317 GND.n116 240.244
R5489 GND.n5313 GND.n116 240.244
R5490 GND.n5313 GND.n126 240.244
R5491 GND.n5305 GND.n126 240.244
R5492 GND.n5305 GND.n137 240.244
R5493 GND.n5301 GND.n137 240.244
R5494 GND.n5301 GND.n147 240.244
R5495 GND.n290 GND.n147 240.244
R5496 GND.n2430 GND.n2429 240.244
R5497 GND.n2426 GND.n2425 240.244
R5498 GND.n2422 GND.n2421 240.244
R5499 GND.n2418 GND.n2417 240.244
R5500 GND.n5590 GND.n2266 240.244
R5501 GND.n5030 GND.n2267 240.244
R5502 GND.n5033 GND.n5032 240.244
R5503 GND.n2666 GND.n2662 240.244
R5504 GND.n5438 GND.n5437 240.244
R5505 GND.n5437 GND.n2434 240.244
R5506 GND.n5429 GND.n2434 240.244
R5507 GND.n5429 GND.n2450 240.244
R5508 GND.n5425 GND.n2450 240.244
R5509 GND.n5425 GND.n2456 240.244
R5510 GND.n5417 GND.n2456 240.244
R5511 GND.n5417 GND.n2471 240.244
R5512 GND.n5413 GND.n2471 240.244
R5513 GND.n5413 GND.n2476 240.244
R5514 GND.n5405 GND.n2476 240.244
R5515 GND.n5405 GND.n2492 240.244
R5516 GND.n5401 GND.n2492 240.244
R5517 GND.n5401 GND.n2497 240.244
R5518 GND.n5393 GND.n2497 240.244
R5519 GND.n5393 GND.n2513 240.244
R5520 GND.n5389 GND.n2513 240.244
R5521 GND.n5389 GND.n2518 240.244
R5522 GND.n5381 GND.n2518 240.244
R5523 GND.n5381 GND.n2532 240.244
R5524 GND.n5377 GND.n2532 240.244
R5525 GND.n5377 GND.n2537 240.244
R5526 GND.n5129 GND.n2537 240.244
R5527 GND.n5129 GND.n35 240.244
R5528 GND.n2556 GND.n35 240.244
R5529 GND.n5360 GND.n2556 240.244
R5530 GND.n5360 GND.n54 240.244
R5531 GND.n8070 GND.n54 240.244
R5532 GND.n8070 GND.n55 240.244
R5533 GND.n8066 GND.n55 240.244
R5534 GND.n8066 GND.n61 240.244
R5535 GND.n8058 GND.n61 240.244
R5536 GND.n8058 GND.n76 240.244
R5537 GND.n8054 GND.n76 240.244
R5538 GND.n8054 GND.n81 240.244
R5539 GND.n8046 GND.n81 240.244
R5540 GND.n8046 GND.n97 240.244
R5541 GND.n8042 GND.n97 240.244
R5542 GND.n8042 GND.n102 240.244
R5543 GND.n8034 GND.n102 240.244
R5544 GND.n8034 GND.n118 240.244
R5545 GND.n8030 GND.n118 240.244
R5546 GND.n8030 GND.n123 240.244
R5547 GND.n8022 GND.n123 240.244
R5548 GND.n8022 GND.n139 240.244
R5549 GND.n8018 GND.n139 240.244
R5550 GND.n8018 GND.n144 240.244
R5551 GND.n6632 GND.n1085 240.244
R5552 GND.n6632 GND.n1083 240.244
R5553 GND.n6636 GND.n1083 240.244
R5554 GND.n6636 GND.n1079 240.244
R5555 GND.n6642 GND.n1079 240.244
R5556 GND.n6642 GND.n1077 240.244
R5557 GND.n6646 GND.n1077 240.244
R5558 GND.n6646 GND.n1073 240.244
R5559 GND.n6652 GND.n1073 240.244
R5560 GND.n6652 GND.n1071 240.244
R5561 GND.n6656 GND.n1071 240.244
R5562 GND.n6656 GND.n1067 240.244
R5563 GND.n6662 GND.n1067 240.244
R5564 GND.n6662 GND.n1065 240.244
R5565 GND.n6666 GND.n1065 240.244
R5566 GND.n6666 GND.n1061 240.244
R5567 GND.n6672 GND.n1061 240.244
R5568 GND.n6672 GND.n1059 240.244
R5569 GND.n6676 GND.n1059 240.244
R5570 GND.n6676 GND.n1055 240.244
R5571 GND.n6682 GND.n1055 240.244
R5572 GND.n6682 GND.n1053 240.244
R5573 GND.n6686 GND.n1053 240.244
R5574 GND.n6686 GND.n1049 240.244
R5575 GND.n6692 GND.n1049 240.244
R5576 GND.n6692 GND.n1047 240.244
R5577 GND.n6696 GND.n1047 240.244
R5578 GND.n6696 GND.n1043 240.244
R5579 GND.n6702 GND.n1043 240.244
R5580 GND.n6702 GND.n1041 240.244
R5581 GND.n6706 GND.n1041 240.244
R5582 GND.n6706 GND.n1037 240.244
R5583 GND.n6712 GND.n1037 240.244
R5584 GND.n6712 GND.n1035 240.244
R5585 GND.n6716 GND.n1035 240.244
R5586 GND.n6716 GND.n1031 240.244
R5587 GND.n6722 GND.n1031 240.244
R5588 GND.n6722 GND.n1029 240.244
R5589 GND.n6726 GND.n1029 240.244
R5590 GND.n6726 GND.n1025 240.244
R5591 GND.n6732 GND.n1025 240.244
R5592 GND.n6732 GND.n1023 240.244
R5593 GND.n6736 GND.n1023 240.244
R5594 GND.n6736 GND.n1019 240.244
R5595 GND.n6742 GND.n1019 240.244
R5596 GND.n6742 GND.n1017 240.244
R5597 GND.n6746 GND.n1017 240.244
R5598 GND.n6746 GND.n1013 240.244
R5599 GND.n6752 GND.n1013 240.244
R5600 GND.n6752 GND.n1011 240.244
R5601 GND.n6756 GND.n1011 240.244
R5602 GND.n6756 GND.n1007 240.244
R5603 GND.n6762 GND.n1007 240.244
R5604 GND.n6762 GND.n1005 240.244
R5605 GND.n6766 GND.n1005 240.244
R5606 GND.n6766 GND.n1001 240.244
R5607 GND.n6772 GND.n1001 240.244
R5608 GND.n6772 GND.n999 240.244
R5609 GND.n6776 GND.n999 240.244
R5610 GND.n6776 GND.n995 240.244
R5611 GND.n6782 GND.n995 240.244
R5612 GND.n6782 GND.n993 240.244
R5613 GND.n6786 GND.n993 240.244
R5614 GND.n6786 GND.n989 240.244
R5615 GND.n6792 GND.n989 240.244
R5616 GND.n6792 GND.n987 240.244
R5617 GND.n6796 GND.n987 240.244
R5618 GND.n6796 GND.n983 240.244
R5619 GND.n6802 GND.n983 240.244
R5620 GND.n6802 GND.n981 240.244
R5621 GND.n6806 GND.n981 240.244
R5622 GND.n6806 GND.n977 240.244
R5623 GND.n6812 GND.n977 240.244
R5624 GND.n6812 GND.n975 240.244
R5625 GND.n6816 GND.n975 240.244
R5626 GND.n6816 GND.n971 240.244
R5627 GND.n6822 GND.n971 240.244
R5628 GND.n6822 GND.n969 240.244
R5629 GND.n6826 GND.n969 240.244
R5630 GND.n6826 GND.n965 240.244
R5631 GND.n6832 GND.n965 240.244
R5632 GND.n6832 GND.n963 240.244
R5633 GND.n6836 GND.n963 240.244
R5634 GND.n6836 GND.n959 240.244
R5635 GND.n6842 GND.n959 240.244
R5636 GND.n6842 GND.n957 240.244
R5637 GND.n6846 GND.n957 240.244
R5638 GND.n6846 GND.n953 240.244
R5639 GND.n6852 GND.n953 240.244
R5640 GND.n6852 GND.n951 240.244
R5641 GND.n6856 GND.n951 240.244
R5642 GND.n6856 GND.n947 240.244
R5643 GND.n6862 GND.n947 240.244
R5644 GND.n6862 GND.n945 240.244
R5645 GND.n6866 GND.n945 240.244
R5646 GND.n6866 GND.n941 240.244
R5647 GND.n6872 GND.n941 240.244
R5648 GND.n6872 GND.n939 240.244
R5649 GND.n6876 GND.n939 240.244
R5650 GND.n6876 GND.n935 240.244
R5651 GND.n6882 GND.n935 240.244
R5652 GND.n6882 GND.n933 240.244
R5653 GND.n6886 GND.n933 240.244
R5654 GND.n6886 GND.n929 240.244
R5655 GND.n6892 GND.n929 240.244
R5656 GND.n6892 GND.n927 240.244
R5657 GND.n6896 GND.n927 240.244
R5658 GND.n6896 GND.n923 240.244
R5659 GND.n6902 GND.n923 240.244
R5660 GND.n6902 GND.n921 240.244
R5661 GND.n6906 GND.n921 240.244
R5662 GND.n6906 GND.n917 240.244
R5663 GND.n6912 GND.n917 240.244
R5664 GND.n6912 GND.n915 240.244
R5665 GND.n6916 GND.n915 240.244
R5666 GND.n6916 GND.n911 240.244
R5667 GND.n6922 GND.n911 240.244
R5668 GND.n6922 GND.n909 240.244
R5669 GND.n6926 GND.n909 240.244
R5670 GND.n6926 GND.n905 240.244
R5671 GND.n6932 GND.n905 240.244
R5672 GND.n6932 GND.n903 240.244
R5673 GND.n6936 GND.n903 240.244
R5674 GND.n6936 GND.n899 240.244
R5675 GND.n6942 GND.n899 240.244
R5676 GND.n6942 GND.n897 240.244
R5677 GND.n6946 GND.n897 240.244
R5678 GND.n6946 GND.n893 240.244
R5679 GND.n6952 GND.n893 240.244
R5680 GND.n6952 GND.n891 240.244
R5681 GND.n6956 GND.n891 240.244
R5682 GND.n6956 GND.n887 240.244
R5683 GND.n6962 GND.n887 240.244
R5684 GND.n6962 GND.n885 240.244
R5685 GND.n6966 GND.n885 240.244
R5686 GND.n6966 GND.n881 240.244
R5687 GND.n6972 GND.n881 240.244
R5688 GND.n6972 GND.n879 240.244
R5689 GND.n6976 GND.n879 240.244
R5690 GND.n6976 GND.n875 240.244
R5691 GND.n6982 GND.n875 240.244
R5692 GND.n6982 GND.n873 240.244
R5693 GND.n6986 GND.n873 240.244
R5694 GND.n6986 GND.n869 240.244
R5695 GND.n6992 GND.n869 240.244
R5696 GND.n6992 GND.n867 240.244
R5697 GND.n6996 GND.n867 240.244
R5698 GND.n6996 GND.n863 240.244
R5699 GND.n7002 GND.n863 240.244
R5700 GND.n7002 GND.n861 240.244
R5701 GND.n7006 GND.n861 240.244
R5702 GND.n7006 GND.n857 240.244
R5703 GND.n7012 GND.n857 240.244
R5704 GND.n7012 GND.n855 240.244
R5705 GND.n7016 GND.n855 240.244
R5706 GND.n7016 GND.n851 240.244
R5707 GND.n7022 GND.n851 240.244
R5708 GND.n7022 GND.n849 240.244
R5709 GND.n7026 GND.n849 240.244
R5710 GND.n7026 GND.n845 240.244
R5711 GND.n7032 GND.n845 240.244
R5712 GND.n7032 GND.n843 240.244
R5713 GND.n7036 GND.n843 240.244
R5714 GND.n7036 GND.n839 240.244
R5715 GND.n7042 GND.n839 240.244
R5716 GND.n7042 GND.n837 240.244
R5717 GND.n7046 GND.n837 240.244
R5718 GND.n7046 GND.n833 240.244
R5719 GND.n7052 GND.n833 240.244
R5720 GND.n7052 GND.n831 240.244
R5721 GND.n7056 GND.n831 240.244
R5722 GND.n7056 GND.n827 240.244
R5723 GND.n7062 GND.n827 240.244
R5724 GND.n7062 GND.n825 240.244
R5725 GND.n7066 GND.n825 240.244
R5726 GND.n7066 GND.n821 240.244
R5727 GND.n7072 GND.n821 240.244
R5728 GND.n7072 GND.n819 240.244
R5729 GND.n7076 GND.n819 240.244
R5730 GND.n7076 GND.n815 240.244
R5731 GND.n7082 GND.n815 240.244
R5732 GND.n7082 GND.n813 240.244
R5733 GND.n7086 GND.n813 240.244
R5734 GND.n7086 GND.n809 240.244
R5735 GND.n7092 GND.n809 240.244
R5736 GND.n7092 GND.n807 240.244
R5737 GND.n7096 GND.n807 240.244
R5738 GND.n7096 GND.n803 240.244
R5739 GND.n7102 GND.n803 240.244
R5740 GND.n7102 GND.n801 240.244
R5741 GND.n7106 GND.n801 240.244
R5742 GND.n7106 GND.n797 240.244
R5743 GND.n7112 GND.n797 240.244
R5744 GND.n7112 GND.n795 240.244
R5745 GND.n7116 GND.n795 240.244
R5746 GND.n7116 GND.n791 240.244
R5747 GND.n7122 GND.n791 240.244
R5748 GND.n7122 GND.n789 240.244
R5749 GND.n7126 GND.n789 240.244
R5750 GND.n7126 GND.n785 240.244
R5751 GND.n7132 GND.n785 240.244
R5752 GND.n7132 GND.n783 240.244
R5753 GND.n7136 GND.n783 240.244
R5754 GND.n7136 GND.n779 240.244
R5755 GND.n7142 GND.n779 240.244
R5756 GND.n7142 GND.n777 240.244
R5757 GND.n7146 GND.n777 240.244
R5758 GND.n7146 GND.n773 240.244
R5759 GND.n7152 GND.n773 240.244
R5760 GND.n7152 GND.n771 240.244
R5761 GND.n7156 GND.n771 240.244
R5762 GND.n7156 GND.n767 240.244
R5763 GND.n7162 GND.n767 240.244
R5764 GND.n7162 GND.n765 240.244
R5765 GND.n7166 GND.n765 240.244
R5766 GND.n7166 GND.n761 240.244
R5767 GND.n7172 GND.n761 240.244
R5768 GND.n7172 GND.n759 240.244
R5769 GND.n7176 GND.n759 240.244
R5770 GND.n7176 GND.n755 240.244
R5771 GND.n7182 GND.n755 240.244
R5772 GND.n7182 GND.n753 240.244
R5773 GND.n7186 GND.n753 240.244
R5774 GND.n7186 GND.n749 240.244
R5775 GND.n7192 GND.n749 240.244
R5776 GND.n7192 GND.n747 240.244
R5777 GND.n7196 GND.n747 240.244
R5778 GND.n7196 GND.n743 240.244
R5779 GND.n7202 GND.n743 240.244
R5780 GND.n7202 GND.n741 240.244
R5781 GND.n7206 GND.n741 240.244
R5782 GND.n7206 GND.n737 240.244
R5783 GND.n7212 GND.n737 240.244
R5784 GND.n7212 GND.n735 240.244
R5785 GND.n7216 GND.n735 240.244
R5786 GND.n7216 GND.n731 240.244
R5787 GND.n7222 GND.n731 240.244
R5788 GND.n7222 GND.n729 240.244
R5789 GND.n7226 GND.n729 240.244
R5790 GND.n7226 GND.n725 240.244
R5791 GND.n7232 GND.n725 240.244
R5792 GND.n7232 GND.n723 240.244
R5793 GND.n7236 GND.n723 240.244
R5794 GND.n7236 GND.n719 240.244
R5795 GND.n7242 GND.n719 240.244
R5796 GND.n7242 GND.n717 240.244
R5797 GND.n7246 GND.n717 240.244
R5798 GND.n7246 GND.n713 240.244
R5799 GND.n7252 GND.n713 240.244
R5800 GND.n7252 GND.n711 240.244
R5801 GND.n7256 GND.n711 240.244
R5802 GND.n7256 GND.n707 240.244
R5803 GND.n7262 GND.n707 240.244
R5804 GND.n7262 GND.n705 240.244
R5805 GND.n7266 GND.n705 240.244
R5806 GND.n7266 GND.n701 240.244
R5807 GND.n7272 GND.n701 240.244
R5808 GND.n7272 GND.n699 240.244
R5809 GND.n7276 GND.n699 240.244
R5810 GND.n7276 GND.n695 240.244
R5811 GND.n7282 GND.n695 240.244
R5812 GND.n7282 GND.n693 240.244
R5813 GND.n7286 GND.n693 240.244
R5814 GND.n7286 GND.n689 240.244
R5815 GND.n7292 GND.n689 240.244
R5816 GND.n7292 GND.n687 240.244
R5817 GND.n7296 GND.n687 240.244
R5818 GND.n7296 GND.n683 240.244
R5819 GND.n7302 GND.n683 240.244
R5820 GND.n7302 GND.n681 240.244
R5821 GND.n7306 GND.n681 240.244
R5822 GND.n7306 GND.n677 240.244
R5823 GND.n7312 GND.n677 240.244
R5824 GND.n7312 GND.n675 240.244
R5825 GND.n7316 GND.n675 240.244
R5826 GND.n7316 GND.n671 240.244
R5827 GND.n7322 GND.n671 240.244
R5828 GND.n7322 GND.n669 240.244
R5829 GND.n7326 GND.n669 240.244
R5830 GND.n7326 GND.n665 240.244
R5831 GND.n7332 GND.n665 240.244
R5832 GND.n7332 GND.n663 240.244
R5833 GND.n7336 GND.n663 240.244
R5834 GND.n7336 GND.n659 240.244
R5835 GND.n7342 GND.n659 240.244
R5836 GND.n7342 GND.n657 240.244
R5837 GND.n7346 GND.n657 240.244
R5838 GND.n7346 GND.n653 240.244
R5839 GND.n7352 GND.n653 240.244
R5840 GND.n7352 GND.n651 240.244
R5841 GND.n7356 GND.n651 240.244
R5842 GND.n7356 GND.n647 240.244
R5843 GND.n7362 GND.n647 240.244
R5844 GND.n7362 GND.n645 240.244
R5845 GND.n7366 GND.n645 240.244
R5846 GND.n7366 GND.n641 240.244
R5847 GND.n7372 GND.n641 240.244
R5848 GND.n7372 GND.n639 240.244
R5849 GND.n7376 GND.n639 240.244
R5850 GND.n7376 GND.n635 240.244
R5851 GND.n7382 GND.n635 240.244
R5852 GND.n7382 GND.n633 240.244
R5853 GND.n7386 GND.n633 240.244
R5854 GND.n7386 GND.n629 240.244
R5855 GND.n7392 GND.n629 240.244
R5856 GND.n7392 GND.n627 240.244
R5857 GND.n7396 GND.n627 240.244
R5858 GND.n7396 GND.n623 240.244
R5859 GND.n7402 GND.n623 240.244
R5860 GND.n7402 GND.n621 240.244
R5861 GND.n7406 GND.n621 240.244
R5862 GND.n7406 GND.n617 240.244
R5863 GND.n7412 GND.n617 240.244
R5864 GND.n7412 GND.n615 240.244
R5865 GND.n7416 GND.n615 240.244
R5866 GND.n7416 GND.n611 240.244
R5867 GND.n7422 GND.n611 240.244
R5868 GND.n7422 GND.n609 240.244
R5869 GND.n7426 GND.n609 240.244
R5870 GND.n7426 GND.n605 240.244
R5871 GND.n7432 GND.n605 240.244
R5872 GND.n7432 GND.n603 240.244
R5873 GND.n7436 GND.n603 240.244
R5874 GND.n7436 GND.n599 240.244
R5875 GND.n7442 GND.n599 240.244
R5876 GND.n7442 GND.n597 240.244
R5877 GND.n7446 GND.n597 240.244
R5878 GND.n7446 GND.n593 240.244
R5879 GND.n7452 GND.n593 240.244
R5880 GND.n7452 GND.n591 240.244
R5881 GND.n7456 GND.n591 240.244
R5882 GND.n7456 GND.n587 240.244
R5883 GND.n7462 GND.n587 240.244
R5884 GND.n7462 GND.n585 240.244
R5885 GND.n7466 GND.n585 240.244
R5886 GND.n7466 GND.n581 240.244
R5887 GND.n7472 GND.n581 240.244
R5888 GND.n7472 GND.n579 240.244
R5889 GND.n7476 GND.n579 240.244
R5890 GND.n7476 GND.n575 240.244
R5891 GND.n7482 GND.n575 240.244
R5892 GND.n7482 GND.n573 240.244
R5893 GND.n7486 GND.n573 240.244
R5894 GND.n7486 GND.n569 240.244
R5895 GND.n7492 GND.n569 240.244
R5896 GND.n7492 GND.n567 240.244
R5897 GND.n7496 GND.n567 240.244
R5898 GND.n7496 GND.n563 240.244
R5899 GND.n7502 GND.n563 240.244
R5900 GND.n7502 GND.n561 240.244
R5901 GND.n7506 GND.n561 240.244
R5902 GND.n7506 GND.n557 240.244
R5903 GND.n7512 GND.n557 240.244
R5904 GND.n7512 GND.n555 240.244
R5905 GND.n7516 GND.n555 240.244
R5906 GND.n7516 GND.n551 240.244
R5907 GND.n7522 GND.n551 240.244
R5908 GND.n7522 GND.n549 240.244
R5909 GND.n7526 GND.n549 240.244
R5910 GND.n7526 GND.n545 240.244
R5911 GND.n7532 GND.n545 240.244
R5912 GND.n7532 GND.n543 240.244
R5913 GND.n7536 GND.n543 240.244
R5914 GND.n7536 GND.n539 240.244
R5915 GND.n7542 GND.n539 240.244
R5916 GND.n7542 GND.n537 240.244
R5917 GND.n7546 GND.n537 240.244
R5918 GND.n7546 GND.n533 240.244
R5919 GND.n7552 GND.n533 240.244
R5920 GND.n7552 GND.n531 240.244
R5921 GND.n7556 GND.n531 240.244
R5922 GND.n7556 GND.n527 240.244
R5923 GND.n7562 GND.n527 240.244
R5924 GND.n7562 GND.n525 240.244
R5925 GND.n7566 GND.n525 240.244
R5926 GND.n7566 GND.n521 240.244
R5927 GND.n7572 GND.n521 240.244
R5928 GND.n7572 GND.n519 240.244
R5929 GND.n7576 GND.n519 240.244
R5930 GND.n7576 GND.n515 240.244
R5931 GND.n7582 GND.n515 240.244
R5932 GND.n7582 GND.n513 240.244
R5933 GND.n7586 GND.n513 240.244
R5934 GND.n7586 GND.n509 240.244
R5935 GND.n7592 GND.n509 240.244
R5936 GND.n7596 GND.n507 240.244
R5937 GND.n7596 GND.n503 240.244
R5938 GND.n7602 GND.n503 240.244
R5939 GND.n7602 GND.n501 240.244
R5940 GND.n7606 GND.n501 240.244
R5941 GND.n7606 GND.n497 240.244
R5942 GND.n7612 GND.n497 240.244
R5943 GND.n7612 GND.n495 240.244
R5944 GND.n7616 GND.n495 240.244
R5945 GND.n7616 GND.n491 240.244
R5946 GND.n7622 GND.n491 240.244
R5947 GND.n7622 GND.n489 240.244
R5948 GND.n7626 GND.n489 240.244
R5949 GND.n7626 GND.n485 240.244
R5950 GND.n7632 GND.n485 240.244
R5951 GND.n7632 GND.n483 240.244
R5952 GND.n7636 GND.n483 240.244
R5953 GND.n7636 GND.n479 240.244
R5954 GND.n7642 GND.n479 240.244
R5955 GND.n7642 GND.n477 240.244
R5956 GND.n7646 GND.n477 240.244
R5957 GND.n7646 GND.n473 240.244
R5958 GND.n7652 GND.n473 240.244
R5959 GND.n7652 GND.n471 240.244
R5960 GND.n7656 GND.n471 240.244
R5961 GND.n7656 GND.n467 240.244
R5962 GND.n7662 GND.n467 240.244
R5963 GND.n7662 GND.n465 240.244
R5964 GND.n7666 GND.n465 240.244
R5965 GND.n7666 GND.n461 240.244
R5966 GND.n7672 GND.n461 240.244
R5967 GND.n7672 GND.n459 240.244
R5968 GND.n7676 GND.n459 240.244
R5969 GND.n7676 GND.n455 240.244
R5970 GND.n7682 GND.n455 240.244
R5971 GND.n7682 GND.n453 240.244
R5972 GND.n7686 GND.n453 240.244
R5973 GND.n7686 GND.n449 240.244
R5974 GND.n7692 GND.n449 240.244
R5975 GND.n7692 GND.n447 240.244
R5976 GND.n7696 GND.n447 240.244
R5977 GND.n7696 GND.n443 240.244
R5978 GND.n7702 GND.n443 240.244
R5979 GND.n7702 GND.n441 240.244
R5980 GND.n7706 GND.n441 240.244
R5981 GND.n7706 GND.n437 240.244
R5982 GND.n7712 GND.n437 240.244
R5983 GND.n7712 GND.n435 240.244
R5984 GND.n7716 GND.n435 240.244
R5985 GND.n7716 GND.n431 240.244
R5986 GND.n7722 GND.n431 240.244
R5987 GND.n7722 GND.n429 240.244
R5988 GND.n7726 GND.n429 240.244
R5989 GND.n7726 GND.n425 240.244
R5990 GND.n7732 GND.n425 240.244
R5991 GND.n7732 GND.n423 240.244
R5992 GND.n7736 GND.n423 240.244
R5993 GND.n7736 GND.n419 240.244
R5994 GND.n7743 GND.n419 240.244
R5995 GND.n7743 GND.n417 240.244
R5996 GND.n7747 GND.n417 240.244
R5997 GND.n7747 GND.n413 240.244
R5998 GND.n6496 GND.n1210 240.244
R5999 GND.n6496 GND.n1214 240.244
R6000 GND.n6492 GND.n1214 240.244
R6001 GND.n6492 GND.n1216 240.244
R6002 GND.n6488 GND.n1216 240.244
R6003 GND.n6488 GND.n1222 240.244
R6004 GND.n6484 GND.n1222 240.244
R6005 GND.n6484 GND.n1224 240.244
R6006 GND.n6480 GND.n1224 240.244
R6007 GND.n6480 GND.n1230 240.244
R6008 GND.n6476 GND.n1230 240.244
R6009 GND.n6476 GND.n1232 240.244
R6010 GND.n6472 GND.n1232 240.244
R6011 GND.n6472 GND.n1238 240.244
R6012 GND.n6468 GND.n1238 240.244
R6013 GND.n6468 GND.n1240 240.244
R6014 GND.n6464 GND.n1240 240.244
R6015 GND.n6464 GND.n1246 240.244
R6016 GND.n6460 GND.n1246 240.244
R6017 GND.n6460 GND.n1248 240.244
R6018 GND.n6456 GND.n1248 240.244
R6019 GND.n6456 GND.n1254 240.244
R6020 GND.n6452 GND.n1254 240.244
R6021 GND.n6452 GND.n1256 240.244
R6022 GND.n6448 GND.n1256 240.244
R6023 GND.n6448 GND.n1262 240.244
R6024 GND.n6444 GND.n1262 240.244
R6025 GND.n6444 GND.n1264 240.244
R6026 GND.n6440 GND.n1264 240.244
R6027 GND.n6440 GND.n1270 240.244
R6028 GND.n6436 GND.n1270 240.244
R6029 GND.n6436 GND.n1272 240.244
R6030 GND.n6432 GND.n1272 240.244
R6031 GND.n6432 GND.n1278 240.244
R6032 GND.n6428 GND.n1278 240.244
R6033 GND.n6428 GND.n1280 240.244
R6034 GND.n6424 GND.n1280 240.244
R6035 GND.n6424 GND.n1286 240.244
R6036 GND.n6420 GND.n1286 240.244
R6037 GND.n6420 GND.n1288 240.244
R6038 GND.n6416 GND.n1288 240.244
R6039 GND.n6416 GND.n1294 240.244
R6040 GND.n6412 GND.n1294 240.244
R6041 GND.n6412 GND.n1296 240.244
R6042 GND.n6408 GND.n1296 240.244
R6043 GND.n6408 GND.n1302 240.244
R6044 GND.n6404 GND.n1302 240.244
R6045 GND.n6404 GND.n1304 240.244
R6046 GND.n6400 GND.n1304 240.244
R6047 GND.n6400 GND.n1310 240.244
R6048 GND.n6396 GND.n1310 240.244
R6049 GND.n6396 GND.n1312 240.244
R6050 GND.n6392 GND.n1312 240.244
R6051 GND.n6392 GND.n1318 240.244
R6052 GND.n6388 GND.n1318 240.244
R6053 GND.n6388 GND.n1320 240.244
R6054 GND.n6384 GND.n1320 240.244
R6055 GND.n6384 GND.n1326 240.244
R6056 GND.n3525 GND.n1326 240.244
R6057 GND.n3531 GND.n3525 240.244
R6058 GND.n3531 GND.n3515 240.244
R6059 GND.n3791 GND.n3515 240.244
R6060 GND.n3791 GND.n3510 240.244
R6061 GND.n3799 GND.n3510 240.244
R6062 GND.n3799 GND.n3511 240.244
R6063 GND.n3511 GND.n3485 240.244
R6064 GND.n3828 GND.n3485 240.244
R6065 GND.n3828 GND.n3480 240.244
R6066 GND.n3836 GND.n3480 240.244
R6067 GND.n3836 GND.n3481 240.244
R6068 GND.n3481 GND.n3456 240.244
R6069 GND.n3865 GND.n3456 240.244
R6070 GND.n3865 GND.n3451 240.244
R6071 GND.n3879 GND.n3451 240.244
R6072 GND.n3879 GND.n3452 240.244
R6073 GND.n3875 GND.n3452 240.244
R6074 GND.n3875 GND.n3874 240.244
R6075 GND.n3874 GND.n3405 240.244
R6076 GND.n3990 GND.n3405 240.244
R6077 GND.n3990 GND.n3406 240.244
R6078 GND.n3938 GND.n3406 240.244
R6079 GND.n3941 GND.n3938 240.244
R6080 GND.n3951 GND.n3941 240.244
R6081 GND.n3951 GND.n3948 240.244
R6082 GND.n3948 GND.n3947 240.244
R6083 GND.n3947 GND.n3944 240.244
R6084 GND.n3944 GND.n3943 240.244
R6085 GND.n3943 GND.n3396 240.244
R6086 GND.n3996 GND.n3396 240.244
R6087 GND.n3996 GND.n3373 240.244
R6088 GND.n4025 GND.n3373 240.244
R6089 GND.n4025 GND.n3368 240.244
R6090 GND.n4033 GND.n3368 240.244
R6091 GND.n4033 GND.n3369 240.244
R6092 GND.n3369 GND.n3344 240.244
R6093 GND.n4062 GND.n3344 240.244
R6094 GND.n4062 GND.n3339 240.244
R6095 GND.n4070 GND.n3339 240.244
R6096 GND.n4070 GND.n3340 240.244
R6097 GND.n3340 GND.n3315 240.244
R6098 GND.n4099 GND.n3315 240.244
R6099 GND.n4099 GND.n3310 240.244
R6100 GND.n4129 GND.n3310 240.244
R6101 GND.n4129 GND.n3311 240.244
R6102 GND.n4125 GND.n3311 240.244
R6103 GND.n4125 GND.n4124 240.244
R6104 GND.n4124 GND.n4123 240.244
R6105 GND.n4123 GND.n4107 240.244
R6106 GND.n4119 GND.n4107 240.244
R6107 GND.n4119 GND.n4118 240.244
R6108 GND.n4118 GND.n4117 240.244
R6109 GND.n4117 GND.n3045 240.244
R6110 GND.n4185 GND.n3045 240.244
R6111 GND.n4185 GND.n3040 240.244
R6112 GND.n4193 GND.n3040 240.244
R6113 GND.n4193 GND.n3041 240.244
R6114 GND.n3041 GND.n3023 240.244
R6115 GND.n4217 GND.n3023 240.244
R6116 GND.n4217 GND.n3018 240.244
R6117 GND.n4225 GND.n3018 240.244
R6118 GND.n4225 GND.n3019 240.244
R6119 GND.n3019 GND.n3000 240.244
R6120 GND.n4249 GND.n3000 240.244
R6121 GND.n4249 GND.n2995 240.244
R6122 GND.n4257 GND.n2995 240.244
R6123 GND.n4257 GND.n2996 240.244
R6124 GND.n2996 GND.n2977 240.244
R6125 GND.n4281 GND.n2977 240.244
R6126 GND.n4281 GND.n2972 240.244
R6127 GND.n4289 GND.n2972 240.244
R6128 GND.n4289 GND.n2973 240.244
R6129 GND.n2973 GND.n2954 240.244
R6130 GND.n4313 GND.n2954 240.244
R6131 GND.n4313 GND.n2949 240.244
R6132 GND.n4321 GND.n2949 240.244
R6133 GND.n4321 GND.n2950 240.244
R6134 GND.n2950 GND.n2931 240.244
R6135 GND.n4345 GND.n2931 240.244
R6136 GND.n4345 GND.n2926 240.244
R6137 GND.n4353 GND.n2926 240.244
R6138 GND.n4353 GND.n2927 240.244
R6139 GND.n2927 GND.n2908 240.244
R6140 GND.n4377 GND.n2908 240.244
R6141 GND.n4377 GND.n2903 240.244
R6142 GND.n4385 GND.n2903 240.244
R6143 GND.n4385 GND.n2904 240.244
R6144 GND.n2904 GND.n2885 240.244
R6145 GND.n4409 GND.n2885 240.244
R6146 GND.n4409 GND.n2880 240.244
R6147 GND.n4417 GND.n2880 240.244
R6148 GND.n4417 GND.n2881 240.244
R6149 GND.n2881 GND.n2862 240.244
R6150 GND.n4441 GND.n2862 240.244
R6151 GND.n4441 GND.n2857 240.244
R6152 GND.n4449 GND.n2857 240.244
R6153 GND.n4449 GND.n2858 240.244
R6154 GND.n2858 GND.n2839 240.244
R6155 GND.n4473 GND.n2839 240.244
R6156 GND.n4473 GND.n2834 240.244
R6157 GND.n4481 GND.n2834 240.244
R6158 GND.n4481 GND.n2835 240.244
R6159 GND.n2835 GND.n2816 240.244
R6160 GND.n4505 GND.n2816 240.244
R6161 GND.n4505 GND.n2811 240.244
R6162 GND.n4513 GND.n2811 240.244
R6163 GND.n4513 GND.n2812 240.244
R6164 GND.n2812 GND.n2793 240.244
R6165 GND.n4540 GND.n2793 240.244
R6166 GND.n4540 GND.n2788 240.244
R6167 GND.n4564 GND.n2788 240.244
R6168 GND.n4564 GND.n2789 240.244
R6169 GND.n4560 GND.n2789 240.244
R6170 GND.n4560 GND.n4559 240.244
R6171 GND.n4559 GND.n4558 240.244
R6172 GND.n4558 GND.n4548 240.244
R6173 GND.n4554 GND.n4548 240.244
R6174 GND.n4554 GND.n1672 240.244
R6175 GND.n6128 GND.n1672 240.244
R6176 GND.n6128 GND.n1673 240.244
R6177 GND.n6124 GND.n1673 240.244
R6178 GND.n6124 GND.n1679 240.244
R6179 GND.n1711 GND.n1679 240.244
R6180 GND.n1711 GND.n1707 240.244
R6181 GND.n6108 GND.n1707 240.244
R6182 GND.n6108 GND.n1708 240.244
R6183 GND.n6104 GND.n1708 240.244
R6184 GND.n6104 GND.n1719 240.244
R6185 GND.n1755 GND.n1719 240.244
R6186 GND.n1755 GND.n1751 240.244
R6187 GND.n6087 GND.n1751 240.244
R6188 GND.n6087 GND.n1752 240.244
R6189 GND.n6083 GND.n1752 240.244
R6190 GND.n6083 GND.n1763 240.244
R6191 GND.n6073 GND.n1763 240.244
R6192 GND.n6073 GND.n1775 240.244
R6193 GND.n6069 GND.n1775 240.244
R6194 GND.n6069 GND.n1781 240.244
R6195 GND.n6059 GND.n1781 240.244
R6196 GND.n6059 GND.n1793 240.244
R6197 GND.n6055 GND.n1793 240.244
R6198 GND.n6055 GND.n1799 240.244
R6199 GND.n6045 GND.n1799 240.244
R6200 GND.n6045 GND.n1810 240.244
R6201 GND.n6041 GND.n1810 240.244
R6202 GND.n6041 GND.n1816 240.244
R6203 GND.n6031 GND.n1816 240.244
R6204 GND.n6031 GND.n1827 240.244
R6205 GND.n6027 GND.n1827 240.244
R6206 GND.n6027 GND.n1833 240.244
R6207 GND.n6017 GND.n1833 240.244
R6208 GND.n6017 GND.n1845 240.244
R6209 GND.n6013 GND.n1845 240.244
R6210 GND.n6013 GND.n1851 240.244
R6211 GND.n5804 GND.n1851 240.244
R6212 GND.n5804 GND.n1915 240.244
R6213 GND.n5800 GND.n1915 240.244
R6214 GND.n5800 GND.n1921 240.244
R6215 GND.n1939 GND.n1921 240.244
R6216 GND.n5790 GND.n1939 240.244
R6217 GND.n5790 GND.n1940 240.244
R6218 GND.n5786 GND.n1940 240.244
R6219 GND.n5786 GND.n1948 240.244
R6220 GND.n1966 GND.n1948 240.244
R6221 GND.n5776 GND.n1966 240.244
R6222 GND.n5776 GND.n1967 240.244
R6223 GND.n5772 GND.n1967 240.244
R6224 GND.n5772 GND.n1975 240.244
R6225 GND.n1993 GND.n1975 240.244
R6226 GND.n5762 GND.n1993 240.244
R6227 GND.n5762 GND.n1994 240.244
R6228 GND.n5758 GND.n1994 240.244
R6229 GND.n5758 GND.n2002 240.244
R6230 GND.n2019 GND.n2002 240.244
R6231 GND.n5748 GND.n2019 240.244
R6232 GND.n5748 GND.n2020 240.244
R6233 GND.n5744 GND.n2020 240.244
R6234 GND.n5744 GND.n2028 240.244
R6235 GND.n2046 GND.n2028 240.244
R6236 GND.n5734 GND.n2046 240.244
R6237 GND.n5734 GND.n2047 240.244
R6238 GND.n5730 GND.n2047 240.244
R6239 GND.n5730 GND.n2055 240.244
R6240 GND.n2073 GND.n2055 240.244
R6241 GND.n5720 GND.n2073 240.244
R6242 GND.n5720 GND.n2074 240.244
R6243 GND.n5716 GND.n2074 240.244
R6244 GND.n5716 GND.n2082 240.244
R6245 GND.n2100 GND.n2082 240.244
R6246 GND.n5706 GND.n2100 240.244
R6247 GND.n5706 GND.n2101 240.244
R6248 GND.n5702 GND.n2101 240.244
R6249 GND.n5702 GND.n2109 240.244
R6250 GND.n2127 GND.n2109 240.244
R6251 GND.n5692 GND.n2127 240.244
R6252 GND.n5692 GND.n2128 240.244
R6253 GND.n5688 GND.n2128 240.244
R6254 GND.n5688 GND.n2136 240.244
R6255 GND.n2154 GND.n2136 240.244
R6256 GND.n5678 GND.n2154 240.244
R6257 GND.n5678 GND.n2155 240.244
R6258 GND.n5674 GND.n2155 240.244
R6259 GND.n5674 GND.n2163 240.244
R6260 GND.n2180 GND.n2163 240.244
R6261 GND.n5664 GND.n2180 240.244
R6262 GND.n5664 GND.n2181 240.244
R6263 GND.n5660 GND.n2181 240.244
R6264 GND.n5660 GND.n2189 240.244
R6265 GND.n2207 GND.n2189 240.244
R6266 GND.n5650 GND.n2207 240.244
R6267 GND.n5650 GND.n2208 240.244
R6268 GND.n5646 GND.n2208 240.244
R6269 GND.n5646 GND.n2216 240.244
R6270 GND.n2591 GND.n2216 240.244
R6271 GND.n2591 GND.n2588 240.244
R6272 GND.n2597 GND.n2588 240.244
R6273 GND.n2598 GND.n2597 240.244
R6274 GND.n2599 GND.n2598 240.244
R6275 GND.n2599 GND.n2583 240.244
R6276 GND.n2605 GND.n2583 240.244
R6277 GND.n2606 GND.n2605 240.244
R6278 GND.n2607 GND.n2606 240.244
R6279 GND.n2607 GND.n2578 240.244
R6280 GND.n2656 GND.n2578 240.244
R6281 GND.n2656 GND.n2579 240.244
R6282 GND.n2652 GND.n2579 240.244
R6283 GND.n2652 GND.n2651 240.244
R6284 GND.n2651 GND.n2650 240.244
R6285 GND.n2650 GND.n2615 240.244
R6286 GND.n2646 GND.n2615 240.244
R6287 GND.n2646 GND.n2645 240.244
R6288 GND.n2645 GND.n2644 240.244
R6289 GND.n2644 GND.n2621 240.244
R6290 GND.n2640 GND.n2621 240.244
R6291 GND.n2640 GND.n2639 240.244
R6292 GND.n2639 GND.n2638 240.244
R6293 GND.n2638 GND.n2627 240.244
R6294 GND.n2633 GND.n2627 240.244
R6295 GND.n2633 GND.n2632 240.244
R6296 GND.n2632 GND.n2546 240.244
R6297 GND.n5371 GND.n2546 240.244
R6298 GND.n5371 GND.n2547 240.244
R6299 GND.n5366 GND.n2547 240.244
R6300 GND.n5366 GND.n5365 240.244
R6301 GND.n5365 GND.n2550 240.244
R6302 GND.n5143 GND.n2550 240.244
R6303 GND.n5201 GND.n5143 240.244
R6304 GND.n5201 GND.n5144 240.244
R6305 GND.n5197 GND.n5144 240.244
R6306 GND.n5197 GND.n5196 240.244
R6307 GND.n5196 GND.n5195 240.244
R6308 GND.n5195 GND.n5152 240.244
R6309 GND.n5191 GND.n5152 240.244
R6310 GND.n5191 GND.n5190 240.244
R6311 GND.n5190 GND.n5189 240.244
R6312 GND.n5189 GND.n5158 240.244
R6313 GND.n5185 GND.n5158 240.244
R6314 GND.n5185 GND.n5184 240.244
R6315 GND.n5184 GND.n5183 240.244
R6316 GND.n5183 GND.n5164 240.244
R6317 GND.n5179 GND.n5164 240.244
R6318 GND.n5179 GND.n5178 240.244
R6319 GND.n5178 GND.n5177 240.244
R6320 GND.n5177 GND.n5170 240.244
R6321 GND.n5170 GND.n292 240.244
R6322 GND.n7873 GND.n292 240.244
R6323 GND.n7873 GND.n293 240.244
R6324 GND.n7869 GND.n293 240.244
R6325 GND.n7869 GND.n299 240.244
R6326 GND.n7865 GND.n299 240.244
R6327 GND.n7865 GND.n301 240.244
R6328 GND.n7861 GND.n301 240.244
R6329 GND.n7861 GND.n307 240.244
R6330 GND.n7857 GND.n307 240.244
R6331 GND.n7857 GND.n309 240.244
R6332 GND.n7853 GND.n309 240.244
R6333 GND.n7853 GND.n315 240.244
R6334 GND.n7849 GND.n315 240.244
R6335 GND.n7849 GND.n317 240.244
R6336 GND.n7845 GND.n317 240.244
R6337 GND.n7845 GND.n323 240.244
R6338 GND.n7841 GND.n323 240.244
R6339 GND.n7841 GND.n325 240.244
R6340 GND.n7837 GND.n325 240.244
R6341 GND.n7837 GND.n331 240.244
R6342 GND.n7833 GND.n331 240.244
R6343 GND.n7833 GND.n333 240.244
R6344 GND.n7829 GND.n333 240.244
R6345 GND.n7829 GND.n339 240.244
R6346 GND.n7825 GND.n339 240.244
R6347 GND.n7825 GND.n341 240.244
R6348 GND.n7821 GND.n341 240.244
R6349 GND.n7821 GND.n347 240.244
R6350 GND.n7817 GND.n347 240.244
R6351 GND.n7817 GND.n349 240.244
R6352 GND.n7813 GND.n349 240.244
R6353 GND.n7813 GND.n355 240.244
R6354 GND.n7809 GND.n355 240.244
R6355 GND.n7809 GND.n357 240.244
R6356 GND.n7805 GND.n357 240.244
R6357 GND.n7805 GND.n363 240.244
R6358 GND.n7801 GND.n363 240.244
R6359 GND.n7801 GND.n365 240.244
R6360 GND.n7797 GND.n365 240.244
R6361 GND.n7797 GND.n371 240.244
R6362 GND.n7793 GND.n371 240.244
R6363 GND.n7793 GND.n373 240.244
R6364 GND.n7789 GND.n373 240.244
R6365 GND.n7789 GND.n379 240.244
R6366 GND.n7785 GND.n379 240.244
R6367 GND.n7785 GND.n381 240.244
R6368 GND.n7781 GND.n381 240.244
R6369 GND.n7781 GND.n387 240.244
R6370 GND.n7777 GND.n387 240.244
R6371 GND.n7777 GND.n389 240.244
R6372 GND.n7773 GND.n389 240.244
R6373 GND.n7773 GND.n395 240.244
R6374 GND.n7769 GND.n395 240.244
R6375 GND.n7769 GND.n397 240.244
R6376 GND.n7765 GND.n397 240.244
R6377 GND.n7765 GND.n403 240.244
R6378 GND.n7761 GND.n403 240.244
R6379 GND.n7761 GND.n405 240.244
R6380 GND.n7757 GND.n405 240.244
R6381 GND.n7757 GND.n411 240.244
R6382 GND.n7753 GND.n411 240.244
R6383 GND.n6626 GND.n1089 240.244
R6384 GND.n6622 GND.n1089 240.244
R6385 GND.n6622 GND.n1091 240.244
R6386 GND.n6618 GND.n1091 240.244
R6387 GND.n6618 GND.n1096 240.244
R6388 GND.n6614 GND.n1096 240.244
R6389 GND.n6614 GND.n1098 240.244
R6390 GND.n6610 GND.n1098 240.244
R6391 GND.n6610 GND.n1104 240.244
R6392 GND.n6606 GND.n1104 240.244
R6393 GND.n6606 GND.n1106 240.244
R6394 GND.n6602 GND.n1106 240.244
R6395 GND.n6602 GND.n1112 240.244
R6396 GND.n6598 GND.n1112 240.244
R6397 GND.n6598 GND.n1114 240.244
R6398 GND.n6594 GND.n1114 240.244
R6399 GND.n6594 GND.n1120 240.244
R6400 GND.n6590 GND.n1120 240.244
R6401 GND.n6590 GND.n1122 240.244
R6402 GND.n6586 GND.n1122 240.244
R6403 GND.n6586 GND.n1128 240.244
R6404 GND.n6582 GND.n1128 240.244
R6405 GND.n6582 GND.n1130 240.244
R6406 GND.n6578 GND.n1130 240.244
R6407 GND.n6578 GND.n1136 240.244
R6408 GND.n6574 GND.n1136 240.244
R6409 GND.n6574 GND.n1138 240.244
R6410 GND.n6570 GND.n1138 240.244
R6411 GND.n6570 GND.n1144 240.244
R6412 GND.n6566 GND.n1144 240.244
R6413 GND.n6566 GND.n1146 240.244
R6414 GND.n6562 GND.n1146 240.244
R6415 GND.n6562 GND.n1152 240.244
R6416 GND.n6558 GND.n1152 240.244
R6417 GND.n6558 GND.n1154 240.244
R6418 GND.n6554 GND.n1154 240.244
R6419 GND.n6554 GND.n1160 240.244
R6420 GND.n6550 GND.n1160 240.244
R6421 GND.n6550 GND.n1162 240.244
R6422 GND.n6546 GND.n1162 240.244
R6423 GND.n6546 GND.n1168 240.244
R6424 GND.n6542 GND.n1168 240.244
R6425 GND.n6542 GND.n1170 240.244
R6426 GND.n6538 GND.n1170 240.244
R6427 GND.n6538 GND.n1176 240.244
R6428 GND.n6534 GND.n1176 240.244
R6429 GND.n6534 GND.n1178 240.244
R6430 GND.n6530 GND.n1178 240.244
R6431 GND.n6530 GND.n1184 240.244
R6432 GND.n6526 GND.n1184 240.244
R6433 GND.n6526 GND.n1186 240.244
R6434 GND.n6522 GND.n1186 240.244
R6435 GND.n6522 GND.n1192 240.244
R6436 GND.n6518 GND.n1192 240.244
R6437 GND.n6518 GND.n1194 240.244
R6438 GND.n6514 GND.n1194 240.244
R6439 GND.n6514 GND.n1200 240.244
R6440 GND.n6510 GND.n1200 240.244
R6441 GND.n6510 GND.n1202 240.244
R6442 GND.n6506 GND.n1202 240.244
R6443 GND.n6506 GND.n1208 240.244
R6444 GND.n6502 GND.n1208 240.244
R6445 GND.n6380 GND.n1375 240.244
R6446 GND.n1380 GND.n1379 240.244
R6447 GND.n1382 GND.n1381 240.244
R6448 GND.n1386 GND.n1385 240.244
R6449 GND.n1388 GND.n1387 240.244
R6450 GND.n1392 GND.n1391 240.244
R6451 GND.n1394 GND.n1393 240.244
R6452 GND.n1398 GND.n1397 240.244
R6453 GND.n6352 GND.n1372 240.244
R6454 GND.n3766 GND.n1374 240.244
R6455 GND.n3766 GND.n3519 240.244
R6456 GND.n3769 GND.n3519 240.244
R6457 GND.n3769 GND.n3500 240.244
R6458 GND.n3815 GND.n3500 240.244
R6459 GND.n3815 GND.n3501 240.244
R6460 GND.n3501 GND.n3490 240.244
R6461 GND.n3806 GND.n3490 240.244
R6462 GND.n3806 GND.n3471 240.244
R6463 GND.n3852 GND.n3471 240.244
R6464 GND.n3852 GND.n3472 240.244
R6465 GND.n3472 GND.n3461 240.244
R6466 GND.n3843 GND.n3461 240.244
R6467 GND.n3843 GND.n3443 240.244
R6468 GND.n3892 GND.n3443 240.244
R6469 GND.n3892 GND.n3429 240.244
R6470 GND.n3903 GND.n3429 240.244
R6471 GND.n3904 GND.n3903 240.244
R6472 GND.n3904 GND.n3411 240.244
R6473 GND.n3420 GND.n3411 240.244
R6474 GND.n3980 GND.n3420 240.244
R6475 GND.n3980 GND.n3421 240.244
R6476 GND.n3955 GND.n3421 240.244
R6477 GND.n3958 GND.n3955 240.244
R6478 GND.n3958 GND.n3957 240.244
R6479 GND.n3957 GND.n3922 240.244
R6480 GND.n3928 GND.n3922 240.244
R6481 GND.n3928 GND.n3387 240.244
R6482 GND.n4012 GND.n3387 240.244
R6483 GND.n4012 GND.n3388 240.244
R6484 GND.n3388 GND.n3378 240.244
R6485 GND.n4003 GND.n3378 240.244
R6486 GND.n4003 GND.n3359 240.244
R6487 GND.n4049 GND.n3359 240.244
R6488 GND.n4049 GND.n3360 240.244
R6489 GND.n3360 GND.n3349 240.244
R6490 GND.n4040 GND.n3349 240.244
R6491 GND.n4040 GND.n3330 240.244
R6492 GND.n4086 GND.n3330 240.244
R6493 GND.n4086 GND.n3331 240.244
R6494 GND.n3331 GND.n3319 240.244
R6495 GND.n4077 GND.n3319 240.244
R6496 GND.n4077 GND.n3302 240.244
R6497 GND.n4141 GND.n3302 240.244
R6498 GND.n4141 GND.n3291 240.244
R6499 GND.n4152 GND.n3291 240.244
R6500 GND.n4153 GND.n4152 240.244
R6501 GND.n3080 GND.n1495 240.244
R6502 GND.n3082 GND.n3081 240.244
R6503 GND.n3090 GND.n3089 240.244
R6504 GND.n3100 GND.n3099 240.244
R6505 GND.n3102 GND.n3101 240.244
R6506 GND.n3109 GND.n3108 240.244
R6507 GND.n3117 GND.n3116 240.244
R6508 GND.n3119 GND.n3118 240.244
R6509 GND.n6274 GND.n1463 240.244
R6510 GND.n1401 GND.n1400 240.244
R6511 GND.n1402 GND.n1401 240.244
R6512 GND.n3508 GND.n1402 240.244
R6513 GND.n3508 GND.n1405 240.244
R6514 GND.n1406 GND.n1405 240.244
R6515 GND.n1407 GND.n1406 240.244
R6516 GND.n3488 GND.n1407 240.244
R6517 GND.n3488 GND.n1410 240.244
R6518 GND.n1411 GND.n1410 240.244
R6519 GND.n1412 GND.n1411 240.244
R6520 GND.n3457 GND.n1412 240.244
R6521 GND.n3457 GND.n1415 240.244
R6522 GND.n1416 GND.n1415 240.244
R6523 GND.n1417 GND.n1416 240.244
R6524 GND.n3441 GND.n1417 240.244
R6525 GND.n3441 GND.n1420 240.244
R6526 GND.n1421 GND.n1420 240.244
R6527 GND.n1422 GND.n1421 240.244
R6528 GND.n3409 GND.n1422 240.244
R6529 GND.n3409 GND.n1425 240.244
R6530 GND.n1426 GND.n1425 240.244
R6531 GND.n1427 GND.n1426 240.244
R6532 GND.n3953 GND.n1427 240.244
R6533 GND.n3953 GND.n1430 240.244
R6534 GND.n1431 GND.n1430 240.244
R6535 GND.n1432 GND.n1431 240.244
R6536 GND.n3924 GND.n1432 240.244
R6537 GND.n3924 GND.n1435 240.244
R6538 GND.n1436 GND.n1435 240.244
R6539 GND.n1437 GND.n1436 240.244
R6540 GND.n3376 GND.n1437 240.244
R6541 GND.n3376 GND.n1440 240.244
R6542 GND.n1441 GND.n1440 240.244
R6543 GND.n1442 GND.n1441 240.244
R6544 GND.n3345 GND.n1442 240.244
R6545 GND.n3345 GND.n1445 240.244
R6546 GND.n1446 GND.n1445 240.244
R6547 GND.n1447 GND.n1446 240.244
R6548 GND.n3328 GND.n1447 240.244
R6549 GND.n3328 GND.n1450 240.244
R6550 GND.n1451 GND.n1450 240.244
R6551 GND.n1452 GND.n1451 240.244
R6552 GND.n4131 GND.n1452 240.244
R6553 GND.n4131 GND.n1455 240.244
R6554 GND.n1456 GND.n1455 240.244
R6555 GND.n1457 GND.n1456 240.244
R6556 GND.n1464 GND.n1457 240.244
R6557 GND.n1627 GND.n1626 240.132
R6558 GND.n1625 GND.n1624 240.132
R6559 GND.n5857 GND.n5856 240.132
R6560 GND.n5855 GND.n5854 240.132
R6561 GND.n2260 GND.t163 229.686
R6562 GND.n3138 GND.t153 229.686
R6563 GND.n2354 GND.n2284 199.319
R6564 GND.n2354 GND.n2285 199.319
R6565 GND.n1572 GND.n1496 199.319
R6566 GND.n1628 GND.n1623 186.49
R6567 GND.n5858 GND.n5853 186.49
R6568 GND.n2260 GND.t165 172.375
R6569 GND.n3138 GND.t156 172.375
R6570 GND.n5933 GND.n5932 163.367
R6571 GND.n5929 GND.n5928 163.367
R6572 GND.n5925 GND.n5924 163.367
R6573 GND.n5921 GND.n5920 163.367
R6574 GND.n5917 GND.n5916 163.367
R6575 GND.n5913 GND.n5912 163.367
R6576 GND.n5909 GND.n5908 163.367
R6577 GND.n5905 GND.n5904 163.367
R6578 GND.n5901 GND.n5900 163.367
R6579 GND.n5897 GND.n5896 163.367
R6580 GND.n5893 GND.n5892 163.367
R6581 GND.n5889 GND.n5888 163.367
R6582 GND.n5885 GND.n5884 163.367
R6583 GND.n5881 GND.n5880 163.367
R6584 GND.n5877 GND.n5876 163.367
R6585 GND.n5872 GND.n5871 163.367
R6586 GND.n5868 GND.n5867 163.367
R6587 GND.n6010 GND.n6009 163.367
R6588 GND.n6006 GND.n6005 163.367
R6589 GND.n6001 GND.n6000 163.367
R6590 GND.n5997 GND.n5996 163.367
R6591 GND.n5993 GND.n5992 163.367
R6592 GND.n5989 GND.n5988 163.367
R6593 GND.n5985 GND.n5984 163.367
R6594 GND.n5981 GND.n5980 163.367
R6595 GND.n5977 GND.n5976 163.367
R6596 GND.n5973 GND.n5972 163.367
R6597 GND.n5969 GND.n5968 163.367
R6598 GND.n5965 GND.n5964 163.367
R6599 GND.n5961 GND.n5960 163.367
R6600 GND.n5957 GND.n5956 163.367
R6601 GND.n5953 GND.n5952 163.367
R6602 GND.n5949 GND.n5948 163.367
R6603 GND.n5945 GND.n5944 163.367
R6604 GND.n4651 GND.n1650 163.367
R6605 GND.n2770 GND.n1650 163.367
R6606 GND.n4668 GND.n2770 163.367
R6607 GND.n4668 GND.n1663 163.367
R6608 GND.n4673 GND.n1663 163.367
R6609 GND.n4673 GND.n1670 163.367
R6610 GND.n2767 GND.n1670 163.367
R6611 GND.n4681 GND.n2767 163.367
R6612 GND.n4681 GND.n2768 163.367
R6613 GND.n4677 GND.n2768 163.367
R6614 GND.n4677 GND.n2758 163.367
R6615 GND.n4716 GND.n2758 163.367
R6616 GND.n4716 GND.n1698 163.367
R6617 GND.n4720 GND.n1698 163.367
R6618 GND.n4720 GND.n1706 163.367
R6619 GND.n4724 GND.n1706 163.367
R6620 GND.n4728 GND.n4724 163.367
R6621 GND.n4728 GND.n1721 163.367
R6622 GND.n4732 GND.n1721 163.367
R6623 GND.n4732 GND.n1729 163.367
R6624 GND.n4736 GND.n1729 163.367
R6625 GND.n4736 GND.n2751 163.367
R6626 GND.n4740 GND.n2751 163.367
R6627 GND.n4741 GND.n4740 163.367
R6628 GND.n4741 GND.n2756 163.367
R6629 GND.n4752 GND.n2756 163.367
R6630 GND.n4752 GND.n1765 163.367
R6631 GND.n4748 GND.n1765 163.367
R6632 GND.n4748 GND.n1773 163.367
R6633 GND.n2740 GND.n1773 163.367
R6634 GND.n4813 GND.n2740 163.367
R6635 GND.n4814 GND.n4813 163.367
R6636 GND.n4814 GND.n1783 163.367
R6637 GND.n4819 GND.n1783 163.367
R6638 GND.n4819 GND.n1791 163.367
R6639 GND.n2737 GND.n1791 163.367
R6640 GND.n4840 GND.n2737 163.367
R6641 GND.n4840 GND.n2738 163.367
R6642 GND.n2738 GND.n1801 163.367
R6643 GND.n4835 GND.n1801 163.367
R6644 GND.n4835 GND.n1808 163.367
R6645 GND.n4832 GND.n1808 163.367
R6646 GND.n4832 GND.n4831 163.367
R6647 GND.n4831 GND.n4830 163.367
R6648 GND.n4830 GND.n1818 163.367
R6649 GND.n4826 GND.n1818 163.367
R6650 GND.n4826 GND.n1825 163.367
R6651 GND.n1895 GND.n1825 163.367
R6652 GND.n5822 GND.n1895 163.367
R6653 GND.n5823 GND.n5822 163.367
R6654 GND.n5823 GND.n1835 163.367
R6655 GND.n5828 GND.n1835 163.367
R6656 GND.n5828 GND.n1843 163.367
R6657 GND.n5832 GND.n1843 163.367
R6658 GND.n5940 GND.n5832 163.367
R6659 GND.n1615 GND.n1614 163.367
R6660 GND.n6208 GND.n1614 163.367
R6661 GND.n6206 GND.n6205 163.367
R6662 GND.n6202 GND.n6201 163.367
R6663 GND.n6198 GND.n6197 163.367
R6664 GND.n6194 GND.n6193 163.367
R6665 GND.n6190 GND.n6189 163.367
R6666 GND.n6186 GND.n6185 163.367
R6667 GND.n6182 GND.n6181 163.367
R6668 GND.n6178 GND.n6177 163.367
R6669 GND.n6174 GND.n6173 163.367
R6670 GND.n6170 GND.n6169 163.367
R6671 GND.n6166 GND.n6165 163.367
R6672 GND.n6162 GND.n6161 163.367
R6673 GND.n6158 GND.n6157 163.367
R6674 GND.n6154 GND.n6153 163.367
R6675 GND.n6217 GND.n1577 163.367
R6676 GND.n1595 GND.n1574 163.367
R6677 GND.n4585 GND.n4584 163.367
R6678 GND.n4590 GND.n4589 163.367
R6679 GND.n4594 GND.n4593 163.367
R6680 GND.n4598 GND.n4597 163.367
R6681 GND.n4602 GND.n4601 163.367
R6682 GND.n4606 GND.n4605 163.367
R6683 GND.n4610 GND.n4609 163.367
R6684 GND.n4614 GND.n4613 163.367
R6685 GND.n4618 GND.n4617 163.367
R6686 GND.n4622 GND.n4621 163.367
R6687 GND.n4626 GND.n4625 163.367
R6688 GND.n4630 GND.n4629 163.367
R6689 GND.n4634 GND.n4633 163.367
R6690 GND.n4638 GND.n4637 163.367
R6691 GND.n4642 GND.n4641 163.367
R6692 GND.n4646 GND.n4645 163.367
R6693 GND.n6145 GND.n1616 163.367
R6694 GND.n6145 GND.n1648 163.367
R6695 GND.n1664 GND.n1648 163.367
R6696 GND.n6135 GND.n1664 163.367
R6697 GND.n6135 GND.n1665 163.367
R6698 GND.n6131 GND.n1665 163.367
R6699 GND.n6131 GND.n1668 163.367
R6700 GND.n4689 GND.n1668 163.367
R6701 GND.n4689 GND.n4682 163.367
R6702 GND.n4685 GND.n4682 163.367
R6703 GND.n4685 GND.n4684 163.367
R6704 GND.n4684 GND.n1700 163.367
R6705 GND.n6114 GND.n1700 163.367
R6706 GND.n6114 GND.n1701 163.367
R6707 GND.n6110 GND.n1701 163.367
R6708 GND.n6110 GND.n1704 163.367
R6709 GND.n1723 GND.n1704 163.367
R6710 GND.n6101 GND.n1723 163.367
R6711 GND.n6101 GND.n1724 163.367
R6712 GND.n6097 GND.n1724 163.367
R6713 GND.n6097 GND.n1727 163.367
R6714 GND.n4761 GND.n1727 163.367
R6715 GND.n4761 GND.n2753 163.367
R6716 GND.n4757 GND.n2753 163.367
R6717 GND.n4757 GND.n4756 163.367
R6718 GND.n4756 GND.n1767 163.367
R6719 GND.n6080 GND.n1767 163.367
R6720 GND.n6080 GND.n1768 163.367
R6721 GND.n6076 GND.n1768 163.367
R6722 GND.n6076 GND.n1771 163.367
R6723 GND.n4811 GND.n1771 163.367
R6724 GND.n4811 GND.n1785 163.367
R6725 GND.n6066 GND.n1785 163.367
R6726 GND.n6066 GND.n1786 163.367
R6727 GND.n6062 GND.n1786 163.367
R6728 GND.n6062 GND.n1789 163.367
R6729 GND.n4844 GND.n1789 163.367
R6730 GND.n4844 GND.n1802 163.367
R6731 GND.n6052 GND.n1802 163.367
R6732 GND.n6052 GND.n1803 163.367
R6733 GND.n6048 GND.n1803 163.367
R6734 GND.n6048 GND.n1806 163.367
R6735 GND.n2720 GND.n1806 163.367
R6736 GND.n2720 GND.n1820 163.367
R6737 GND.n6038 GND.n1820 163.367
R6738 GND.n6038 GND.n1821 163.367
R6739 GND.n6034 GND.n1821 163.367
R6740 GND.n6034 GND.n1824 163.367
R6741 GND.n5820 GND.n1824 163.367
R6742 GND.n5820 GND.n1837 163.367
R6743 GND.n6024 GND.n1837 163.367
R6744 GND.n6024 GND.n1838 163.367
R6745 GND.n6020 GND.n1838 163.367
R6746 GND.n6020 GND.n1841 163.367
R6747 GND.n5938 GND.n1841 163.367
R6748 GND.n5864 GND.n5863 157.237
R6749 GND.n1633 GND.n1632 152
R6750 GND.n1634 GND.n1621 152
R6751 GND.n1636 GND.n1635 152
R6752 GND.n1639 GND.n1638 152
R6753 GND.n1640 GND.n1619 152
R6754 GND.n1642 GND.n1641 152
R6755 GND.n1644 GND.n1617 152
R6756 GND.n1646 GND.n1645 152
R6757 GND.n5862 GND.n5836 152
R6758 GND.n5852 GND.n5837 152
R6759 GND.n5851 GND.n5850 152
R6760 GND.n5849 GND.n5838 152
R6761 GND.n5846 GND.n5839 152
R6762 GND.n5845 GND.n5844 152
R6763 GND.n5843 GND.n5840 152
R6764 GND.n5841 GND.t108 149.72
R6765 GND.n2376 GND.t55 148.911
R6766 GND.n284 GND.t68 148.911
R6767 GND.n1889 GND.n1870 143.351
R6768 GND.n6216 GND.n1575 143.351
R6769 GND.n1594 GND.n1575 143.351
R6770 GND.n1460 GND.t136 139.31
R6771 GND.n1538 GND.t97 139.31
R6772 GND.n3193 GND.t94 139.31
R6773 GND.n3174 GND.t85 139.31
R6774 GND.n1569 GND.t158 139.31
R6775 GND.n2335 GND.t61 139.31
R6776 GND.n2356 GND.t122 139.31
R6777 GND.n2396 GND.t82 139.31
R6778 GND.n247 GND.t71 139.31
R6779 GND.n214 GND.t139 139.31
R6780 GND.n181 GND.t74 139.31
R6781 GND.n5232 GND.t103 139.31
R6782 GND.n2663 GND.t125 139.31
R6783 GND.n3616 GND.t131 139.31
R6784 GND.n3665 GND.t65 139.31
R6785 GND.n3711 GND.t128 139.31
R6786 GND.n3538 GND.t101 139.31
R6787 GND.n6353 GND.t146 139.31
R6788 GND.n10 GND.t14 135.601
R6789 GND.n12 GND.t16 134.078
R6790 GND.n11 GND.t27 134.078
R6791 GND.n10 GND.t21 134.078
R6792 GND.n1630 GND.t39 129.018
R6793 GND.n1645 GND.t117 126.766
R6794 GND.n1643 GND.t150 126.766
R6795 GND.n1619 GND.t105 126.766
R6796 GND.n1637 GND.t160 126.766
R6797 GND.n1621 GND.t56 126.766
R6798 GND.n1631 GND.t147 126.766
R6799 GND.n5842 GND.t87 126.766
R6800 GND.n5844 GND.t132 126.766
R6801 GND.n5848 GND.t46 126.766
R6802 GND.n5850 GND.t49 126.766
R6803 GND.n5861 GND.t90 126.766
R6804 GND.n5863 GND.t114 126.766
R6805 GND.n2261 GND.n2260 114.037
R6806 GND.n3139 GND.n3138 114.037
R6807 GND.n4581 GND.t79 100.046
R6808 GND.n1891 GND.t112 100.046
R6809 GND.n6149 GND.t143 100.037
R6810 GND.n5865 GND.t44 100.037
R6811 GND.n8009 GND.n8008 99.6594
R6812 GND.n8006 GND.n8005 99.6594
R6813 GND.n8001 GND.n162 99.6594
R6814 GND.n7999 GND.n7998 99.6594
R6815 GND.n7994 GND.n169 99.6594
R6816 GND.n7992 GND.n7991 99.6594
R6817 GND.n7987 GND.n176 99.6594
R6818 GND.n7985 GND.n7984 99.6594
R6819 GND.n186 GND.n185 99.6594
R6820 GND.n7976 GND.n7975 99.6594
R6821 GND.n7973 GND.n7972 99.6594
R6822 GND.n7968 GND.n194 99.6594
R6823 GND.n7966 GND.n7965 99.6594
R6824 GND.n7961 GND.n201 99.6594
R6825 GND.n7959 GND.n7958 99.6594
R6826 GND.n7954 GND.n208 99.6594
R6827 GND.n7952 GND.n7951 99.6594
R6828 GND.n217 GND.n216 99.6594
R6829 GND.n7943 GND.n221 99.6594
R6830 GND.n7941 GND.n7940 99.6594
R6831 GND.n7936 GND.n227 99.6594
R6832 GND.n7934 GND.n7933 99.6594
R6833 GND.n7929 GND.n234 99.6594
R6834 GND.n7927 GND.n7926 99.6594
R6835 GND.n7922 GND.n241 99.6594
R6836 GND.n7920 GND.n7919 99.6594
R6837 GND.n7915 GND.n250 99.6594
R6838 GND.n7913 GND.n7912 99.6594
R6839 GND.n7908 GND.n258 99.6594
R6840 GND.n7906 GND.n7905 99.6594
R6841 GND.n7901 GND.n265 99.6594
R6842 GND.n7899 GND.n7898 99.6594
R6843 GND.n7894 GND.n272 99.6594
R6844 GND.n7892 GND.n7891 99.6594
R6845 GND.n7887 GND.n279 99.6594
R6846 GND.n7885 GND.n7884 99.6594
R6847 GND.n289 GND.n288 99.6594
R6848 GND.n5587 GND.n5586 99.6594
R6849 GND.n5581 GND.n2269 99.6594
R6850 GND.n5578 GND.n2270 99.6594
R6851 GND.n5574 GND.n2271 99.6594
R6852 GND.n5570 GND.n2272 99.6594
R6853 GND.n5566 GND.n2273 99.6594
R6854 GND.n5562 GND.n2274 99.6594
R6855 GND.n5558 GND.n2275 99.6594
R6856 GND.n5554 GND.n2276 99.6594
R6857 GND.n5551 GND.n2277 99.6594
R6858 GND.n5547 GND.n2278 99.6594
R6859 GND.n5543 GND.n2279 99.6594
R6860 GND.n5539 GND.n2280 99.6594
R6861 GND.n5535 GND.n2281 99.6594
R6862 GND.n5531 GND.n2282 99.6594
R6863 GND.n5527 GND.n2283 99.6594
R6864 GND.n5523 GND.n2284 99.6594
R6865 GND.n5518 GND.n2286 99.6594
R6866 GND.n5514 GND.n2287 99.6594
R6867 GND.n5510 GND.n2288 99.6594
R6868 GND.n5506 GND.n2289 99.6594
R6869 GND.n5502 GND.n2290 99.6594
R6870 GND.n5498 GND.n2291 99.6594
R6871 GND.n5494 GND.n2292 99.6594
R6872 GND.n5490 GND.n2293 99.6594
R6873 GND.n5486 GND.n2294 99.6594
R6874 GND.n5481 GND.n2295 99.6594
R6875 GND.n5477 GND.n2296 99.6594
R6876 GND.n5473 GND.n2297 99.6594
R6877 GND.n5469 GND.n2298 99.6594
R6878 GND.n5465 GND.n2299 99.6594
R6879 GND.n5461 GND.n2300 99.6594
R6880 GND.n5457 GND.n2301 99.6594
R6881 GND.n5453 GND.n2302 99.6594
R6882 GND.n5449 GND.n2303 99.6594
R6883 GND.n1518 GND.n1512 99.6594
R6884 GND.n1520 GND.n1511 99.6594
R6885 GND.n1524 GND.n1510 99.6594
R6886 GND.n1526 GND.n1509 99.6594
R6887 GND.n1530 GND.n1508 99.6594
R6888 GND.n1532 GND.n1507 99.6594
R6889 GND.n1536 GND.n1506 99.6594
R6890 GND.n1541 GND.n1505 99.6594
R6891 GND.n1545 GND.n1504 99.6594
R6892 GND.n1547 GND.n1503 99.6594
R6893 GND.n1551 GND.n1502 99.6594
R6894 GND.n1553 GND.n1501 99.6594
R6895 GND.n1557 GND.n1500 99.6594
R6896 GND.n1559 GND.n1499 99.6594
R6897 GND.n1563 GND.n1498 99.6594
R6898 GND.n1565 GND.n1497 99.6594
R6899 GND.n1572 GND.n1466 99.6594
R6900 GND.n3214 GND.n1467 99.6594
R6901 GND.n3209 GND.n1468 99.6594
R6902 GND.n3222 GND.n1469 99.6594
R6903 GND.n3205 GND.n1470 99.6594
R6904 GND.n3230 GND.n1471 99.6594
R6905 GND.n3201 GND.n1472 99.6594
R6906 GND.n3238 GND.n1473 99.6594
R6907 GND.n3197 GND.n1474 99.6594
R6908 GND.n3246 GND.n1475 99.6594
R6909 GND.n3190 GND.n1476 99.6594
R6910 GND.n3254 GND.n1477 99.6594
R6911 GND.n3186 GND.n1478 99.6594
R6912 GND.n3262 GND.n1479 99.6594
R6913 GND.n3182 GND.n1480 99.6594
R6914 GND.n3270 GND.n1481 99.6594
R6915 GND.n3178 GND.n1482 99.6594
R6916 GND.n3278 GND.n1483 99.6594
R6917 GND.n3284 GND.n1484 99.6594
R6918 GND.n3288 GND.n1485 99.6594
R6919 GND.n3524 GND.n1327 99.6594
R6920 GND.n3577 GND.n1328 99.6594
R6921 GND.n3585 GND.n1329 99.6594
R6922 GND.n3587 GND.n1330 99.6594
R6923 GND.n3595 GND.n1331 99.6594
R6924 GND.n3597 GND.n1332 99.6594
R6925 GND.n3605 GND.n1333 99.6594
R6926 GND.n3607 GND.n1334 99.6594
R6927 GND.n3615 GND.n1335 99.6594
R6928 GND.n3619 GND.n1336 99.6594
R6929 GND.n3627 GND.n1337 99.6594
R6930 GND.n3629 GND.n1338 99.6594
R6931 GND.n3637 GND.n1339 99.6594
R6932 GND.n3639 GND.n1340 99.6594
R6933 GND.n3647 GND.n1341 99.6594
R6934 GND.n3649 GND.n1342 99.6594
R6935 GND.n3657 GND.n1343 99.6594
R6936 GND.n3659 GND.n1344 99.6594
R6937 GND.n3669 GND.n1345 99.6594
R6938 GND.n3671 GND.n1346 99.6594
R6939 GND.n3679 GND.n1347 99.6594
R6940 GND.n3681 GND.n1348 99.6594
R6941 GND.n3689 GND.n1349 99.6594
R6942 GND.n3691 GND.n1350 99.6594
R6943 GND.n3699 GND.n1351 99.6594
R6944 GND.n3701 GND.n1352 99.6594
R6945 GND.n3709 GND.n1353 99.6594
R6946 GND.n3714 GND.n1354 99.6594
R6947 GND.n3722 GND.n1355 99.6594
R6948 GND.n3724 GND.n1356 99.6594
R6949 GND.n3732 GND.n1357 99.6594
R6950 GND.n3734 GND.n1358 99.6594
R6951 GND.n3742 GND.n1359 99.6594
R6952 GND.n3744 GND.n1360 99.6594
R6953 GND.n3752 GND.n1361 99.6594
R6954 GND.n3754 GND.n1362 99.6594
R6955 GND.n3537 GND.n1363 99.6594
R6956 GND.n5634 GND.n2232 99.6594
R6957 GND.n5632 GND.n2231 99.6594
R6958 GND.n5628 GND.n2230 99.6594
R6959 GND.n5624 GND.n2229 99.6594
R6960 GND.n5620 GND.n2228 99.6594
R6961 GND.n5616 GND.n2227 99.6594
R6962 GND.n5612 GND.n2226 99.6594
R6963 GND.n5608 GND.n2225 99.6594
R6964 GND.n5604 GND.n2224 99.6594
R6965 GND.n5600 GND.n2223 99.6594
R6966 GND.n5596 GND.n2222 99.6594
R6967 GND.n5025 GND.n2221 99.6594
R6968 GND.n5023 GND.n2220 99.6594
R6969 GND.n4182 GND.n3036 99.6594
R6970 GND.n4177 GND.n3047 99.6594
R6971 GND.n4174 GND.n3048 99.6594
R6972 GND.n4170 GND.n3049 99.6594
R6973 GND.n4166 GND.n3050 99.6594
R6974 GND.n4162 GND.n3051 99.6594
R6975 GND.n3074 GND.n3052 99.6594
R6976 GND.n3076 GND.n3053 99.6594
R6977 GND.n3086 GND.n3054 99.6594
R6978 GND.n3094 GND.n3055 99.6594
R6979 GND.n3096 GND.n3056 99.6594
R6980 GND.n3137 GND.n3057 99.6594
R6981 GND.n3113 GND.n3058 99.6594
R6982 GND.n5253 GND.n5251 99.6594
R6983 GND.n5259 GND.n5247 99.6594
R6984 GND.n5263 GND.n5261 99.6594
R6985 GND.n5269 GND.n5243 99.6594
R6986 GND.n5273 GND.n5271 99.6594
R6987 GND.n5279 GND.n5239 99.6594
R6988 GND.n5283 GND.n5281 99.6594
R6989 GND.n5289 GND.n5235 99.6594
R6990 GND.n5292 GND.n5291 99.6594
R6991 GND.n2433 GND.n2313 99.6594
R6992 GND.n2429 GND.n2312 99.6594
R6993 GND.n2425 GND.n2311 99.6594
R6994 GND.n2421 GND.n2310 99.6594
R6995 GND.n2417 GND.n2309 99.6594
R6996 GND.n5590 GND.n5589 99.6594
R6997 GND.n5030 GND.n2308 99.6594
R6998 GND.n5032 GND.n2307 99.6594
R6999 GND.n2662 GND.n2306 99.6594
R7000 GND.n2430 GND.n2313 99.6594
R7001 GND.n2426 GND.n2312 99.6594
R7002 GND.n2422 GND.n2311 99.6594
R7003 GND.n2418 GND.n2310 99.6594
R7004 GND.n2309 GND.n2266 99.6594
R7005 GND.n5589 GND.n2267 99.6594
R7006 GND.n5033 GND.n2308 99.6594
R7007 GND.n2666 GND.n2307 99.6594
R7008 GND.n5041 GND.n2306 99.6594
R7009 GND.n5291 GND.n5290 99.6594
R7010 GND.n5282 GND.n5235 99.6594
R7011 GND.n5281 GND.n5280 99.6594
R7012 GND.n5272 GND.n5239 99.6594
R7013 GND.n5271 GND.n5270 99.6594
R7014 GND.n5262 GND.n5243 99.6594
R7015 GND.n5261 GND.n5260 99.6594
R7016 GND.n5252 GND.n5247 99.6594
R7017 GND.n5251 GND.n5250 99.6594
R7018 GND.n4182 GND.n4181 99.6594
R7019 GND.n4175 GND.n3047 99.6594
R7020 GND.n4171 GND.n3048 99.6594
R7021 GND.n4167 GND.n3049 99.6594
R7022 GND.n4163 GND.n3050 99.6594
R7023 GND.n3073 GND.n3051 99.6594
R7024 GND.n3075 GND.n3052 99.6594
R7025 GND.n3085 GND.n3053 99.6594
R7026 GND.n3093 GND.n3054 99.6594
R7027 GND.n3095 GND.n3055 99.6594
R7028 GND.n3105 GND.n3056 99.6594
R7029 GND.n3112 GND.n3057 99.6594
R7030 GND.n3114 GND.n3058 99.6594
R7031 GND.n5026 GND.n2220 99.6594
R7032 GND.n5595 GND.n2221 99.6594
R7033 GND.n5599 GND.n2222 99.6594
R7034 GND.n5603 GND.n2223 99.6594
R7035 GND.n5607 GND.n2224 99.6594
R7036 GND.n5611 GND.n2225 99.6594
R7037 GND.n5615 GND.n2226 99.6594
R7038 GND.n5619 GND.n2227 99.6594
R7039 GND.n5623 GND.n2228 99.6594
R7040 GND.n5627 GND.n2229 99.6594
R7041 GND.n5631 GND.n2230 99.6594
R7042 GND.n5635 GND.n2231 99.6594
R7043 GND.n2234 GND.n2232 99.6594
R7044 GND.n3578 GND.n1327 99.6594
R7045 GND.n3584 GND.n1328 99.6594
R7046 GND.n3588 GND.n1329 99.6594
R7047 GND.n3594 GND.n1330 99.6594
R7048 GND.n3598 GND.n1331 99.6594
R7049 GND.n3604 GND.n1332 99.6594
R7050 GND.n3608 GND.n1333 99.6594
R7051 GND.n3614 GND.n1334 99.6594
R7052 GND.n3620 GND.n1335 99.6594
R7053 GND.n3626 GND.n1336 99.6594
R7054 GND.n3630 GND.n1337 99.6594
R7055 GND.n3636 GND.n1338 99.6594
R7056 GND.n3640 GND.n1339 99.6594
R7057 GND.n3646 GND.n1340 99.6594
R7058 GND.n3650 GND.n1341 99.6594
R7059 GND.n3656 GND.n1342 99.6594
R7060 GND.n3660 GND.n1343 99.6594
R7061 GND.n3668 GND.n1344 99.6594
R7062 GND.n3672 GND.n1345 99.6594
R7063 GND.n3678 GND.n1346 99.6594
R7064 GND.n3682 GND.n1347 99.6594
R7065 GND.n3688 GND.n1348 99.6594
R7066 GND.n3692 GND.n1349 99.6594
R7067 GND.n3698 GND.n1350 99.6594
R7068 GND.n3702 GND.n1351 99.6594
R7069 GND.n3708 GND.n1352 99.6594
R7070 GND.n3715 GND.n1353 99.6594
R7071 GND.n3721 GND.n1354 99.6594
R7072 GND.n3725 GND.n1355 99.6594
R7073 GND.n3731 GND.n1356 99.6594
R7074 GND.n3735 GND.n1357 99.6594
R7075 GND.n3741 GND.n1358 99.6594
R7076 GND.n3745 GND.n1359 99.6594
R7077 GND.n3751 GND.n1360 99.6594
R7078 GND.n3755 GND.n1361 99.6594
R7079 GND.n3541 GND.n1362 99.6594
R7080 GND.n3533 GND.n1363 99.6594
R7081 GND.n3285 GND.n1485 99.6594
R7082 GND.n3279 GND.n1484 99.6594
R7083 GND.n3179 GND.n1483 99.6594
R7084 GND.n3271 GND.n1482 99.6594
R7085 GND.n3183 GND.n1481 99.6594
R7086 GND.n3263 GND.n1480 99.6594
R7087 GND.n3187 GND.n1479 99.6594
R7088 GND.n3255 GND.n1478 99.6594
R7089 GND.n3191 GND.n1477 99.6594
R7090 GND.n3247 GND.n1476 99.6594
R7091 GND.n3198 GND.n1475 99.6594
R7092 GND.n3239 GND.n1474 99.6594
R7093 GND.n3202 GND.n1473 99.6594
R7094 GND.n3231 GND.n1472 99.6594
R7095 GND.n3206 GND.n1471 99.6594
R7096 GND.n3223 GND.n1470 99.6594
R7097 GND.n3210 GND.n1469 99.6594
R7098 GND.n3215 GND.n1468 99.6594
R7099 GND.n1567 GND.n1467 99.6594
R7100 GND.n6221 GND.n1496 99.6594
R7101 GND.n1564 GND.n1497 99.6594
R7102 GND.n1560 GND.n1498 99.6594
R7103 GND.n1558 GND.n1499 99.6594
R7104 GND.n1554 GND.n1500 99.6594
R7105 GND.n1552 GND.n1501 99.6594
R7106 GND.n1548 GND.n1502 99.6594
R7107 GND.n1546 GND.n1503 99.6594
R7108 GND.n1542 GND.n1504 99.6594
R7109 GND.n1537 GND.n1505 99.6594
R7110 GND.n1533 GND.n1506 99.6594
R7111 GND.n1531 GND.n1507 99.6594
R7112 GND.n1527 GND.n1508 99.6594
R7113 GND.n1525 GND.n1509 99.6594
R7114 GND.n1521 GND.n1510 99.6594
R7115 GND.n1519 GND.n1511 99.6594
R7116 GND.n1514 GND.n1512 99.6594
R7117 GND.n5587 GND.n2315 99.6594
R7118 GND.n5579 GND.n2269 99.6594
R7119 GND.n5575 GND.n2270 99.6594
R7120 GND.n5571 GND.n2271 99.6594
R7121 GND.n5567 GND.n2272 99.6594
R7122 GND.n5563 GND.n2273 99.6594
R7123 GND.n5559 GND.n2274 99.6594
R7124 GND.n2333 GND.n2275 99.6594
R7125 GND.n5552 GND.n2276 99.6594
R7126 GND.n5548 GND.n2277 99.6594
R7127 GND.n5544 GND.n2278 99.6594
R7128 GND.n5540 GND.n2279 99.6594
R7129 GND.n5536 GND.n2280 99.6594
R7130 GND.n5532 GND.n2281 99.6594
R7131 GND.n5528 GND.n2282 99.6594
R7132 GND.n5524 GND.n2283 99.6594
R7133 GND.n5519 GND.n2285 99.6594
R7134 GND.n5515 GND.n2286 99.6594
R7135 GND.n5511 GND.n2287 99.6594
R7136 GND.n5507 GND.n2288 99.6594
R7137 GND.n5503 GND.n2289 99.6594
R7138 GND.n5499 GND.n2290 99.6594
R7139 GND.n5495 GND.n2291 99.6594
R7140 GND.n5491 GND.n2292 99.6594
R7141 GND.n5487 GND.n2293 99.6594
R7142 GND.n5482 GND.n2294 99.6594
R7143 GND.n5478 GND.n2295 99.6594
R7144 GND.n5474 GND.n2296 99.6594
R7145 GND.n5470 GND.n2297 99.6594
R7146 GND.n5466 GND.n2298 99.6594
R7147 GND.n5462 GND.n2299 99.6594
R7148 GND.n5458 GND.n2300 99.6594
R7149 GND.n5454 GND.n2301 99.6594
R7150 GND.n5450 GND.n2302 99.6594
R7151 GND.n2395 GND.n2303 99.6594
R7152 GND.n288 GND.n280 99.6594
R7153 GND.n7886 GND.n7885 99.6594
R7154 GND.n279 GND.n273 99.6594
R7155 GND.n7893 GND.n7892 99.6594
R7156 GND.n272 GND.n266 99.6594
R7157 GND.n7900 GND.n7899 99.6594
R7158 GND.n265 GND.n259 99.6594
R7159 GND.n7907 GND.n7906 99.6594
R7160 GND.n258 GND.n252 99.6594
R7161 GND.n7914 GND.n7913 99.6594
R7162 GND.n250 GND.n242 99.6594
R7163 GND.n7921 GND.n7920 99.6594
R7164 GND.n241 GND.n235 99.6594
R7165 GND.n7928 GND.n7927 99.6594
R7166 GND.n234 GND.n228 99.6594
R7167 GND.n7935 GND.n7934 99.6594
R7168 GND.n227 GND.n222 99.6594
R7169 GND.n7942 GND.n7941 99.6594
R7170 GND.n221 GND.n220 99.6594
R7171 GND.n216 GND.n209 99.6594
R7172 GND.n7953 GND.n7952 99.6594
R7173 GND.n208 GND.n202 99.6594
R7174 GND.n7960 GND.n7959 99.6594
R7175 GND.n201 GND.n195 99.6594
R7176 GND.n7967 GND.n7966 99.6594
R7177 GND.n194 GND.n188 99.6594
R7178 GND.n7974 GND.n7973 99.6594
R7179 GND.n7977 GND.n7976 99.6594
R7180 GND.n185 GND.n177 99.6594
R7181 GND.n7986 GND.n7985 99.6594
R7182 GND.n176 GND.n170 99.6594
R7183 GND.n7993 GND.n7992 99.6594
R7184 GND.n169 GND.n163 99.6594
R7185 GND.n8000 GND.n7999 99.6594
R7186 GND.n162 GND.n156 99.6594
R7187 GND.n8007 GND.n8006 99.6594
R7188 GND.n8010 GND.n8009 99.6594
R7189 GND.n1375 GND.n1364 99.6594
R7190 GND.n1380 GND.n1365 99.6594
R7191 GND.n1382 GND.n1366 99.6594
R7192 GND.n1386 GND.n1367 99.6594
R7193 GND.n1388 GND.n1368 99.6594
R7194 GND.n1392 GND.n1369 99.6594
R7195 GND.n1394 GND.n1370 99.6594
R7196 GND.n1398 GND.n1371 99.6594
R7197 GND.n1379 GND.n1364 99.6594
R7198 GND.n1381 GND.n1365 99.6594
R7199 GND.n1385 GND.n1366 99.6594
R7200 GND.n1387 GND.n1367 99.6594
R7201 GND.n1391 GND.n1368 99.6594
R7202 GND.n1393 GND.n1369 99.6594
R7203 GND.n1397 GND.n1370 99.6594
R7204 GND.n6352 GND.n1371 99.6594
R7205 GND.n3080 GND.n1486 99.6594
R7206 GND.n3082 GND.n1487 99.6594
R7207 GND.n3090 GND.n1488 99.6594
R7208 GND.n3100 GND.n1489 99.6594
R7209 GND.n3102 GND.n1490 99.6594
R7210 GND.n3109 GND.n1491 99.6594
R7211 GND.n3117 GND.n1492 99.6594
R7212 GND.n3119 GND.n1493 99.6594
R7213 GND.n1493 GND.n1463 99.6594
R7214 GND.n3118 GND.n1492 99.6594
R7215 GND.n3116 GND.n1491 99.6594
R7216 GND.n3108 GND.n1490 99.6594
R7217 GND.n3101 GND.n1489 99.6594
R7218 GND.n3099 GND.n1488 99.6594
R7219 GND.n3089 GND.n1487 99.6594
R7220 GND.n3081 GND.n1486 99.6594
R7221 GND.n2377 GND.n2376 97.552
R7222 GND.n285 GND.n284 97.552
R7223 GND.n1461 GND.n1460 84.752
R7224 GND.n1539 GND.n1538 84.752
R7225 GND.n3194 GND.n3193 84.752
R7226 GND.n3175 GND.n3174 84.752
R7227 GND.n1570 GND.n1569 84.752
R7228 GND.n2336 GND.n2335 84.752
R7229 GND.n2357 GND.n2356 84.752
R7230 GND.n2397 GND.n2396 84.752
R7231 GND.n248 GND.n247 84.752
R7232 GND.n215 GND.n214 84.752
R7233 GND.n182 GND.n181 84.752
R7234 GND.n5233 GND.n5232 84.752
R7235 GND.n2664 GND.n2663 84.752
R7236 GND.n3617 GND.n3616 84.752
R7237 GND.n3666 GND.n3665 84.752
R7238 GND.n3712 GND.n3711 84.752
R7239 GND.n3539 GND.n3538 84.752
R7240 GND.n6354 GND.n6353 84.752
R7241 GND.n1630 GND.n1629 83.3186
R7242 GND.n1631 GND.n1622 72.8411
R7243 GND.n1637 GND.n1620 72.8411
R7244 GND.n1643 GND.n1618 72.8411
R7245 GND.n5861 GND.n5860 72.8411
R7246 GND.n5848 GND.n5847 72.8411
R7247 GND.n5933 GND.n1853 71.676
R7248 GND.n5929 GND.n1854 71.676
R7249 GND.n5925 GND.n1855 71.676
R7250 GND.n5921 GND.n1856 71.676
R7251 GND.n5917 GND.n1857 71.676
R7252 GND.n5913 GND.n1858 71.676
R7253 GND.n5909 GND.n1859 71.676
R7254 GND.n5905 GND.n1860 71.676
R7255 GND.n5901 GND.n1861 71.676
R7256 GND.n5897 GND.n1862 71.676
R7257 GND.n5893 GND.n1863 71.676
R7258 GND.n5889 GND.n1864 71.676
R7259 GND.n5885 GND.n1865 71.676
R7260 GND.n5881 GND.n1866 71.676
R7261 GND.n5877 GND.n1867 71.676
R7262 GND.n5872 GND.n1868 71.676
R7263 GND.n5868 GND.n1869 71.676
R7264 GND.n6010 GND.n1889 71.676
R7265 GND.n6006 GND.n1888 71.676
R7266 GND.n6001 GND.n1887 71.676
R7267 GND.n5997 GND.n1886 71.676
R7268 GND.n5993 GND.n1885 71.676
R7269 GND.n5989 GND.n1884 71.676
R7270 GND.n5985 GND.n1883 71.676
R7271 GND.n5981 GND.n1882 71.676
R7272 GND.n5977 GND.n1881 71.676
R7273 GND.n5973 GND.n1880 71.676
R7274 GND.n5969 GND.n1879 71.676
R7275 GND.n5965 GND.n1878 71.676
R7276 GND.n5961 GND.n1877 71.676
R7277 GND.n5957 GND.n1876 71.676
R7278 GND.n5953 GND.n1875 71.676
R7279 GND.n5949 GND.n1874 71.676
R7280 GND.n5945 GND.n1873 71.676
R7281 GND.n5941 GND.n1872 71.676
R7282 GND.n6214 GND.n6213 71.676
R7283 GND.n6208 GND.n1579 71.676
R7284 GND.n6205 GND.n1580 71.676
R7285 GND.n6201 GND.n1581 71.676
R7286 GND.n6197 GND.n1582 71.676
R7287 GND.n6193 GND.n1583 71.676
R7288 GND.n6189 GND.n1584 71.676
R7289 GND.n6185 GND.n1585 71.676
R7290 GND.n6181 GND.n1586 71.676
R7291 GND.n6177 GND.n1587 71.676
R7292 GND.n6173 GND.n1588 71.676
R7293 GND.n6169 GND.n1589 71.676
R7294 GND.n6165 GND.n1590 71.676
R7295 GND.n6161 GND.n1591 71.676
R7296 GND.n6157 GND.n1592 71.676
R7297 GND.n6153 GND.n1593 71.676
R7298 GND.n6217 GND.n6216 71.676
R7299 GND.n1596 GND.n1595 71.676
R7300 GND.n4585 GND.n1597 71.676
R7301 GND.n4590 GND.n1598 71.676
R7302 GND.n4594 GND.n1599 71.676
R7303 GND.n4598 GND.n1600 71.676
R7304 GND.n4602 GND.n1601 71.676
R7305 GND.n4606 GND.n1602 71.676
R7306 GND.n4610 GND.n1603 71.676
R7307 GND.n4614 GND.n1604 71.676
R7308 GND.n4618 GND.n1605 71.676
R7309 GND.n4622 GND.n1606 71.676
R7310 GND.n4626 GND.n1607 71.676
R7311 GND.n4630 GND.n1608 71.676
R7312 GND.n4634 GND.n1609 71.676
R7313 GND.n4638 GND.n1610 71.676
R7314 GND.n4642 GND.n1611 71.676
R7315 GND.n4646 GND.n1612 71.676
R7316 GND.n6214 GND.n1615 71.676
R7317 GND.n6206 GND.n1579 71.676
R7318 GND.n6202 GND.n1580 71.676
R7319 GND.n6198 GND.n1581 71.676
R7320 GND.n6194 GND.n1582 71.676
R7321 GND.n6190 GND.n1583 71.676
R7322 GND.n6186 GND.n1584 71.676
R7323 GND.n6182 GND.n1585 71.676
R7324 GND.n6178 GND.n1586 71.676
R7325 GND.n6174 GND.n1587 71.676
R7326 GND.n6170 GND.n1588 71.676
R7327 GND.n6166 GND.n1589 71.676
R7328 GND.n6162 GND.n1590 71.676
R7329 GND.n6158 GND.n1591 71.676
R7330 GND.n6154 GND.n1592 71.676
R7331 GND.n1593 GND.n1577 71.676
R7332 GND.n1594 GND.n1574 71.676
R7333 GND.n4584 GND.n1596 71.676
R7334 GND.n4589 GND.n1597 71.676
R7335 GND.n4593 GND.n1598 71.676
R7336 GND.n4597 GND.n1599 71.676
R7337 GND.n4601 GND.n1600 71.676
R7338 GND.n4605 GND.n1601 71.676
R7339 GND.n4609 GND.n1602 71.676
R7340 GND.n4613 GND.n1603 71.676
R7341 GND.n4617 GND.n1604 71.676
R7342 GND.n4621 GND.n1605 71.676
R7343 GND.n4625 GND.n1606 71.676
R7344 GND.n4629 GND.n1607 71.676
R7345 GND.n4633 GND.n1608 71.676
R7346 GND.n4637 GND.n1609 71.676
R7347 GND.n4641 GND.n1610 71.676
R7348 GND.n4645 GND.n1611 71.676
R7349 GND.n4580 GND.n1612 71.676
R7350 GND.n5944 GND.n1872 71.676
R7351 GND.n5948 GND.n1873 71.676
R7352 GND.n5952 GND.n1874 71.676
R7353 GND.n5956 GND.n1875 71.676
R7354 GND.n5960 GND.n1876 71.676
R7355 GND.n5964 GND.n1877 71.676
R7356 GND.n5968 GND.n1878 71.676
R7357 GND.n5972 GND.n1879 71.676
R7358 GND.n5976 GND.n1880 71.676
R7359 GND.n5980 GND.n1881 71.676
R7360 GND.n5984 GND.n1882 71.676
R7361 GND.n5988 GND.n1883 71.676
R7362 GND.n5992 GND.n1884 71.676
R7363 GND.n5996 GND.n1885 71.676
R7364 GND.n6000 GND.n1886 71.676
R7365 GND.n6005 GND.n1887 71.676
R7366 GND.n6009 GND.n1888 71.676
R7367 GND.n5867 GND.n1870 71.676
R7368 GND.n5871 GND.n1869 71.676
R7369 GND.n5876 GND.n1868 71.676
R7370 GND.n5880 GND.n1867 71.676
R7371 GND.n5884 GND.n1866 71.676
R7372 GND.n5888 GND.n1865 71.676
R7373 GND.n5892 GND.n1864 71.676
R7374 GND.n5896 GND.n1863 71.676
R7375 GND.n5900 GND.n1862 71.676
R7376 GND.n5904 GND.n1861 71.676
R7377 GND.n5908 GND.n1860 71.676
R7378 GND.n5912 GND.n1859 71.676
R7379 GND.n5916 GND.n1858 71.676
R7380 GND.n5920 GND.n1857 71.676
R7381 GND.n5924 GND.n1856 71.676
R7382 GND.n5928 GND.n1855 71.676
R7383 GND.n5932 GND.n1854 71.676
R7384 GND.n5835 GND.n1853 71.676
R7385 GND.n6625 GND.n6624 68.3447
R7386 GND.n6624 GND.n6623 68.3447
R7387 GND.n6623 GND.n1090 68.3447
R7388 GND.n6617 GND.n1090 68.3447
R7389 GND.n6617 GND.n6616 68.3447
R7390 GND.n6616 GND.n6615 68.3447
R7391 GND.n6615 GND.n1097 68.3447
R7392 GND.n6609 GND.n1097 68.3447
R7393 GND.n6609 GND.n6608 68.3447
R7394 GND.n6608 GND.n6607 68.3447
R7395 GND.n6607 GND.n1105 68.3447
R7396 GND.n6601 GND.n1105 68.3447
R7397 GND.n6601 GND.n6600 68.3447
R7398 GND.n6600 GND.n6599 68.3447
R7399 GND.n6599 GND.n1113 68.3447
R7400 GND.n6593 GND.n1113 68.3447
R7401 GND.n6593 GND.n6592 68.3447
R7402 GND.n6592 GND.n6591 68.3447
R7403 GND.n6591 GND.n1121 68.3447
R7404 GND.n6585 GND.n1121 68.3447
R7405 GND.n6585 GND.n6584 68.3447
R7406 GND.n6584 GND.n6583 68.3447
R7407 GND.n6583 GND.n1129 68.3447
R7408 GND.n6577 GND.n1129 68.3447
R7409 GND.n6577 GND.n6576 68.3447
R7410 GND.n6576 GND.n6575 68.3447
R7411 GND.n6575 GND.n1137 68.3447
R7412 GND.n6569 GND.n1137 68.3447
R7413 GND.n6569 GND.n6568 68.3447
R7414 GND.n6568 GND.n6567 68.3447
R7415 GND.n6567 GND.n1145 68.3447
R7416 GND.n6561 GND.n1145 68.3447
R7417 GND.n6561 GND.n6560 68.3447
R7418 GND.n6560 GND.n6559 68.3447
R7419 GND.n6559 GND.n1153 68.3447
R7420 GND.n6553 GND.n1153 68.3447
R7421 GND.n6553 GND.n6552 68.3447
R7422 GND.n6552 GND.n6551 68.3447
R7423 GND.n6551 GND.n1161 68.3447
R7424 GND.n6545 GND.n1161 68.3447
R7425 GND.n6545 GND.n6544 68.3447
R7426 GND.n6544 GND.n6543 68.3447
R7427 GND.n6543 GND.n1169 68.3447
R7428 GND.n6537 GND.n1169 68.3447
R7429 GND.n6537 GND.n6536 68.3447
R7430 GND.n6536 GND.n6535 68.3447
R7431 GND.n6535 GND.n1177 68.3447
R7432 GND.n6529 GND.n1177 68.3447
R7433 GND.n6529 GND.n6528 68.3447
R7434 GND.n6528 GND.n6527 68.3447
R7435 GND.n6527 GND.n1185 68.3447
R7436 GND.n6521 GND.n1185 68.3447
R7437 GND.n6521 GND.n6520 68.3447
R7438 GND.n6520 GND.n6519 68.3447
R7439 GND.n6519 GND.n1193 68.3447
R7440 GND.n6513 GND.n1193 68.3447
R7441 GND.n6513 GND.n6512 68.3447
R7442 GND.n6512 GND.n6511 68.3447
R7443 GND.n6511 GND.n1201 68.3447
R7444 GND.n6505 GND.n1201 68.3447
R7445 GND.n6505 GND.n6504 68.3447
R7446 GND.n6504 GND.n6503 68.3447
R7447 GND.n13 GND.t3 68.1093
R7448 GND.n15 GND.t5 66.588
R7449 GND.n14 GND.t168 66.588
R7450 GND.n13 GND.t38 66.588
R7451 GND.n6148 GND.n1646 58.4046
R7452 GND.n2261 GND.t166 58.3387
R7453 GND.n3139 GND.t155 58.3387
R7454 GND.n4582 GND.t78 55.2453
R7455 GND.n1892 GND.t113 55.2453
R7456 GND.n6150 GND.t142 55.2378
R7457 GND.n5866 GND.t45 55.2378
R7458 GND.n1461 GND.t137 54.5589
R7459 GND.n1539 GND.t98 54.5589
R7460 GND.n3194 GND.t95 54.5589
R7461 GND.n3175 GND.t86 54.5589
R7462 GND.n1570 GND.t159 54.5589
R7463 GND.n2336 GND.t60 54.5589
R7464 GND.n2357 GND.t121 54.5589
R7465 GND.n2397 GND.t81 54.5589
R7466 GND.n248 GND.t72 54.5589
R7467 GND.n215 GND.t140 54.5589
R7468 GND.n182 GND.t75 54.5589
R7469 GND.n5233 GND.t104 54.5589
R7470 GND.n2664 GND.t124 54.5589
R7471 GND.n3617 GND.t130 54.5589
R7472 GND.n3666 GND.t64 54.5589
R7473 GND.n3712 GND.t127 54.5589
R7474 GND.n3539 GND.t100 54.5589
R7475 GND.n6354 GND.t145 54.5589
R7476 GND.n1628 GND.n1627 54.358
R7477 GND.n5858 GND.n5857 54.358
R7478 GND.n6151 GND.n6150 53.1399
R7479 GND.n4587 GND.n4582 53.1399
R7480 GND.n6003 GND.n1892 53.1399
R7481 GND.n5874 GND.n5866 53.1399
R7482 GND.n5841 GND.n5840 52.3702
R7483 GND.n2377 GND.t54 51.3589
R7484 GND.n285 GND.t69 51.3589
R7485 GND.n1 GND.t25 50.6888
R7486 GND.n2 GND.t36 50.6888
R7487 GND.n4 GND.t1 50.6888
R7488 GND.n6 GND.t24 50.6888
R7489 GND.n0 GND.t9 50.6888
R7490 GND.n17 GND.t29 50.6888
R7491 GND.n18 GND.t22 50.6888
R7492 GND.n20 GND.t7 50.6888
R7493 GND.n22 GND.t8 50.6888
R7494 GND.n24 GND.t31 50.6888
R7495 GND.n1 GND.t33 49.2434
R7496 GND.n2 GND.t19 49.2434
R7497 GND.n4 GND.t30 49.2434
R7498 GND.n6 GND.t34 49.2434
R7499 GND.n0 GND.t28 49.2434
R7500 GND.n17 GND.t32 49.2434
R7501 GND.n18 GND.t35 49.2434
R7502 GND.n20 GND.t11 49.2434
R7503 GND.n22 GND.t12 49.2434
R7504 GND.n24 GND.t17 49.2434
R7505 GND.n5484 GND.n2377 48.6793
R7506 GND.n7882 GND.n285 48.6793
R7507 GND.n1631 GND.n1630 45.8904
R7508 GND.n6150 GND.n6149 44.8005
R7509 GND.n4582 GND.n4581 44.8005
R7510 GND.n1892 GND.n1891 44.8005
R7511 GND.n5866 GND.n5865 44.8005
R7512 GND.n5936 GND.n5864 44.3322
R7513 GND.n1644 GND.n1643 43.8187
R7514 GND.n5862 GND.n5861 43.8187
R7515 GND.n1629 GND.n1628 41.6274
R7516 GND.n5859 GND.n5858 41.6274
R7517 GND.n1638 GND.n1637 37.9763
R7518 GND.n1637 GND.n1636 37.9763
R7519 GND.n5848 GND.n5839 37.9763
R7520 GND.n5849 GND.n5848 37.9763
R7521 GND.n1462 GND.n1461 35.8793
R7522 GND.n6247 GND.n1539 35.8793
R7523 GND.n3195 GND.n3194 35.8793
R7524 GND.n3286 GND.n3175 35.8793
R7525 GND.n5556 GND.n2336 35.8793
R7526 GND.n2398 GND.n2397 35.8793
R7527 GND.n249 GND.n248 35.8793
R7528 GND.n7948 GND.n215 35.8793
R7529 GND.n7982 GND.n182 35.8793
R7530 GND.n5234 GND.n5233 35.8793
R7531 GND.n5040 GND.n2664 35.8793
R7532 GND.n5594 GND.n2261 35.8793
R7533 GND.n3140 GND.n3139 35.8793
R7534 GND.n3618 GND.n3617 35.8793
R7535 GND.n3667 GND.n3666 35.8793
R7536 GND.n3713 GND.n3712 35.8793
R7537 GND.n3761 GND.n3539 35.8793
R7538 GND.n6355 GND.n6354 35.8793
R7539 GND.n5942 GND.n1893 32.6249
R7540 GND.n4650 GND.n4648 32.6249
R7541 GND.n1643 GND.n1642 32.1338
R7542 GND.n1632 GND.n1631 32.1338
R7543 GND.n5843 GND.n5842 32.1338
R7544 GND.n5861 GND.n5837 32.1338
R7545 GND.n6220 GND.n1570 30.5518
R7546 GND.n5521 GND.n2357 30.5518
R7547 GND.n6495 GND.n1209 29.7503
R7548 GND.n6495 GND.n6494 29.7503
R7549 GND.n6494 GND.n6493 29.7503
R7550 GND.n6493 GND.n1215 29.7503
R7551 GND.n6487 GND.n1215 29.7503
R7552 GND.n6487 GND.n6486 29.7503
R7553 GND.n6486 GND.n6485 29.7503
R7554 GND.n6485 GND.n1223 29.7503
R7555 GND.n6479 GND.n1223 29.7503
R7556 GND.n6479 GND.n6478 29.7503
R7557 GND.n6478 GND.n6477 29.7503
R7558 GND.n6477 GND.n1231 29.7503
R7559 GND.n6471 GND.n1231 29.7503
R7560 GND.n6471 GND.n6470 29.7503
R7561 GND.n6470 GND.n6469 29.7503
R7562 GND.n6469 GND.n1239 29.7503
R7563 GND.n6463 GND.n1239 29.7503
R7564 GND.n6463 GND.n6462 29.7503
R7565 GND.n6462 GND.n6461 29.7503
R7566 GND.n6461 GND.n1247 29.7503
R7567 GND.n6455 GND.n1247 29.7503
R7568 GND.n6455 GND.n6454 29.7503
R7569 GND.n6454 GND.n6453 29.7503
R7570 GND.n6453 GND.n1255 29.7503
R7571 GND.n6447 GND.n1255 29.7503
R7572 GND.n6447 GND.n6446 29.7503
R7573 GND.n6446 GND.n6445 29.7503
R7574 GND.n6445 GND.n1263 29.7503
R7575 GND.n6439 GND.n1263 29.7503
R7576 GND.n6439 GND.n6438 29.7503
R7577 GND.n6438 GND.n6437 29.7503
R7578 GND.n6437 GND.n1271 29.7503
R7579 GND.n6431 GND.n1271 29.7503
R7580 GND.n6431 GND.n6430 29.7503
R7581 GND.n6430 GND.n6429 29.7503
R7582 GND.n6429 GND.n1279 29.7503
R7583 GND.n6423 GND.n1279 29.7503
R7584 GND.n6423 GND.n6422 29.7503
R7585 GND.n6422 GND.n6421 29.7503
R7586 GND.n6421 GND.n1287 29.7503
R7587 GND.n6415 GND.n1287 29.7503
R7588 GND.n6415 GND.n6414 29.7503
R7589 GND.n6414 GND.n6413 29.7503
R7590 GND.n6413 GND.n1295 29.7503
R7591 GND.n6407 GND.n1295 29.7503
R7592 GND.n6407 GND.n6406 29.7503
R7593 GND.n6406 GND.n6405 29.7503
R7594 GND.n6405 GND.n1303 29.7503
R7595 GND.n6399 GND.n1303 29.7503
R7596 GND.n6399 GND.n6398 29.7503
R7597 GND.n6398 GND.n6397 29.7503
R7598 GND.n6397 GND.n1311 29.7503
R7599 GND.n6391 GND.n1311 29.7503
R7600 GND.n6391 GND.n6390 29.7503
R7601 GND.n6390 GND.n6389 29.7503
R7602 GND.n6389 GND.n1319 29.7503
R7603 GND.n6383 GND.n1319 29.7503
R7604 GND.n6383 GND.n6382 29.7503
R7605 GND.n3532 GND.n1373 29.7503
R7606 GND.n3290 GND.n1465 29.7503
R7607 GND.n4116 GND.n1494 29.7503
R7608 GND.n4116 GND.n3046 29.7503
R7609 GND.n4184 GND.n3037 29.7503
R7610 GND.n5645 GND.n5644 29.7503
R7611 GND.n2587 GND.n2219 29.7503
R7612 GND.n2587 GND.n2268 29.7503
R7613 GND.n2404 GND.n2305 29.7503
R7614 GND.n7874 GND.n291 29.7503
R7615 GND.n7868 GND.n7867 29.7503
R7616 GND.n7867 GND.n7866 29.7503
R7617 GND.n7866 GND.n300 29.7503
R7618 GND.n7860 GND.n300 29.7503
R7619 GND.n7860 GND.n7859 29.7503
R7620 GND.n7859 GND.n7858 29.7503
R7621 GND.n7858 GND.n308 29.7503
R7622 GND.n7852 GND.n308 29.7503
R7623 GND.n7852 GND.n7851 29.7503
R7624 GND.n7851 GND.n7850 29.7503
R7625 GND.n7850 GND.n316 29.7503
R7626 GND.n7844 GND.n316 29.7503
R7627 GND.n7844 GND.n7843 29.7503
R7628 GND.n7843 GND.n7842 29.7503
R7629 GND.n7842 GND.n324 29.7503
R7630 GND.n7836 GND.n324 29.7503
R7631 GND.n7836 GND.n7835 29.7503
R7632 GND.n7835 GND.n7834 29.7503
R7633 GND.n7834 GND.n332 29.7503
R7634 GND.n7828 GND.n332 29.7503
R7635 GND.n7828 GND.n7827 29.7503
R7636 GND.n7827 GND.n7826 29.7503
R7637 GND.n7826 GND.n340 29.7503
R7638 GND.n7820 GND.n340 29.7503
R7639 GND.n7820 GND.n7819 29.7503
R7640 GND.n7819 GND.n7818 29.7503
R7641 GND.n7818 GND.n348 29.7503
R7642 GND.n7812 GND.n348 29.7503
R7643 GND.n7812 GND.n7811 29.7503
R7644 GND.n7811 GND.n7810 29.7503
R7645 GND.n7810 GND.n356 29.7503
R7646 GND.n7804 GND.n356 29.7503
R7647 GND.n7804 GND.n7803 29.7503
R7648 GND.n7803 GND.n7802 29.7503
R7649 GND.n7802 GND.n364 29.7503
R7650 GND.n7796 GND.n364 29.7503
R7651 GND.n7796 GND.n7795 29.7503
R7652 GND.n7795 GND.n7794 29.7503
R7653 GND.n7794 GND.n372 29.7503
R7654 GND.n7788 GND.n372 29.7503
R7655 GND.n7788 GND.n7787 29.7503
R7656 GND.n7787 GND.n7786 29.7503
R7657 GND.n7786 GND.n380 29.7503
R7658 GND.n7780 GND.n380 29.7503
R7659 GND.n7780 GND.n7779 29.7503
R7660 GND.n7779 GND.n7778 29.7503
R7661 GND.n7778 GND.n388 29.7503
R7662 GND.n7772 GND.n388 29.7503
R7663 GND.n7772 GND.n7771 29.7503
R7664 GND.n7771 GND.n7770 29.7503
R7665 GND.n7770 GND.n396 29.7503
R7666 GND.n7764 GND.n396 29.7503
R7667 GND.n7764 GND.n7763 29.7503
R7668 GND.n7763 GND.n7762 29.7503
R7669 GND.n7762 GND.n404 29.7503
R7670 GND.n7756 GND.n404 29.7503
R7671 GND.n7756 GND.n7755 29.7503
R7672 GND.n7755 GND.n7754 29.7503
R7673 GND.n6382 GND.n6381 22.9079
R7674 GND.n7868 GND.n154 22.9079
R7675 GND.n3779 GND.n3532 22.0154
R7676 GND.n3778 GND.n3516 22.0154
R7677 GND.n3790 GND.n3789 22.0154
R7678 GND.n3518 GND.n3509 22.0154
R7679 GND.n3801 GND.n3800 22.0154
R7680 GND.n3816 GND.n3497 22.0154
R7681 GND.n3827 GND.n3826 22.0154
R7682 GND.n3489 GND.n3479 22.0154
R7683 GND.n3838 GND.n3837 22.0154
R7684 GND.n3853 GND.n3468 22.0154
R7685 GND.n3470 GND.n3458 22.0154
R7686 GND.n3864 GND.n3863 22.0154
R7687 GND.n3460 GND.n3450 22.0154
R7688 GND.n3881 GND.n3880 22.0154
R7689 GND.n3893 GND.n3439 22.0154
R7690 GND.n3884 GND.n3442 22.0154
R7691 GND.n3902 GND.n3430 22.0154
R7692 GND.n3433 GND.n3407 22.0154
R7693 GND.n3909 GND.n3410 22.0154
R7694 GND.n3981 GND.n3417 22.0154
R7695 GND.n3937 GND.n3419 22.0154
R7696 GND.n3954 GND.n3952 22.0154
R7697 GND.n3959 GND.n3934 22.0154
R7698 GND.n3956 GND.n3936 22.0154
R7699 GND.n3968 GND.n3920 22.0154
R7700 GND.n3929 GND.n3921 22.0154
R7701 GND.n3998 GND.n3395 22.0154
R7702 GND.n3386 GND.n3374 22.0154
R7703 GND.n4024 GND.n4023 22.0154
R7704 GND.n3377 GND.n3367 22.0154
R7705 GND.n4035 GND.n4034 22.0154
R7706 GND.n4050 GND.n3356 22.0154
R7707 GND.n3358 GND.n3346 22.0154
R7708 GND.n4061 GND.n4060 22.0154
R7709 GND.n3348 GND.n3338 22.0154
R7710 GND.n4072 GND.n4071 22.0154
R7711 GND.n4087 GND.n3326 22.0154
R7712 GND.n3329 GND.n3316 22.0154
R7713 GND.n4098 GND.n4097 22.0154
R7714 GND.n4132 GND.n4130 22.0154
R7715 GND.n4142 GND.n3299 22.0154
R7716 GND.n4135 GND.n3301 22.0154
R7717 GND.n4151 GND.n3293 22.0154
R7718 GND.n4154 GND.n3289 22.0154
R7719 GND.n5439 GND.n2406 22.0154
R7720 GND.n5436 GND.n2437 22.0154
R7721 GND.n5050 GND.n2446 22.0154
R7722 GND.n5430 GND.n2449 22.0154
R7723 GND.n5058 GND.n2457 22.0154
R7724 GND.n5065 GND.n2467 22.0154
R7725 GND.n5418 GND.n2470 22.0154
R7726 GND.n5073 GND.n2477 22.0154
R7727 GND.n5412 GND.n2480 22.0154
R7728 GND.n5080 GND.n2488 22.0154
R7729 GND.n5406 GND.n2491 22.0154
R7730 GND.n5088 GND.n2498 22.0154
R7731 GND.n5400 GND.n2501 22.0154
R7732 GND.n5095 GND.n2509 22.0154
R7733 GND.n5394 GND.n2512 22.0154
R7734 GND.n5103 GND.n2519 22.0154
R7735 GND.n5388 GND.n2522 22.0154
R7736 GND.n5382 GND.n2531 22.0154
R7737 GND.n5122 GND.n2538 22.0154
R7738 GND.n5376 GND.n2541 22.0154
R7739 GND.n5373 GND.n5372 22.0154
R7740 GND.n2545 GND.n32 22.0154
R7741 GND.n8078 GND.n34 22.0154
R7742 GND.n5364 GND.n2552 22.0154
R7743 GND.n5363 GND.n2555 22.0154
R7744 GND.n5354 GND.n51 22.0154
R7745 GND.n5348 GND.n62 22.0154
R7746 GND.n8065 GND.n65 22.0154
R7747 GND.n5342 GND.n72 22.0154
R7748 GND.n8059 GND.n75 22.0154
R7749 GND.n5336 GND.n82 22.0154
R7750 GND.n8053 GND.n85 22.0154
R7751 GND.n5330 GND.n93 22.0154
R7752 GND.n8047 GND.n96 22.0154
R7753 GND.n5324 GND.n103 22.0154
R7754 GND.n8041 GND.n106 22.0154
R7755 GND.n5318 GND.n114 22.0154
R7756 GND.n8035 GND.n117 22.0154
R7757 GND.n8029 GND.n127 22.0154
R7758 GND.n5306 GND.n135 22.0154
R7759 GND.n8023 GND.n138 22.0154
R7760 GND.n5300 GND.n145 22.0154
R7761 GND.n8017 GND.n148 22.0154
R7762 GND.n7875 GND.n7874 22.0154
R7763 GND.n6273 GND.n1465 21.1229
R7764 GND.n5588 GND.n2305 21.1229
R7765 GND.n1626 GND.t162 19.8005
R7766 GND.n1626 GND.t58 19.8005
R7767 GND.n1624 GND.t152 19.8005
R7768 GND.n1624 GND.t107 19.8005
R7769 GND.n1623 GND.t149 19.8005
R7770 GND.n1623 GND.t41 19.8005
R7771 GND.n5856 GND.t48 19.8005
R7772 GND.n5856 GND.t51 19.8005
R7773 GND.n5854 GND.t89 19.8005
R7774 GND.n5854 GND.t134 19.8005
R7775 GND.n5853 GND.t92 19.8005
R7776 GND.n5853 GND.t116 19.8005
R7777 GND.n6148 GND.n6147 19.5127
R7778 GND.n5937 GND.n5936 19.5127
R7779 GND.n1618 GND.n1617 19.5087
R7780 GND.n1641 GND.n1618 19.5087
R7781 GND.n1639 GND.n1620 19.5087
R7782 GND.n1635 GND.n1620 19.5087
R7783 GND.n1633 GND.n1622 19.5087
R7784 GND.n5847 GND.n5846 19.5087
R7785 GND.n5847 GND.n5838 19.5087
R7786 GND.n5860 GND.n5852 19.5087
R7787 GND.n3161 GND.n3079 19.3944
R7788 GND.n3161 GND.n3160 19.3944
R7789 GND.n3160 GND.n3083 19.3944
R7790 GND.n3153 GND.n3083 19.3944
R7791 GND.n3153 GND.n3152 19.3944
R7792 GND.n3152 GND.n3091 19.3944
R7793 GND.n3145 GND.n3091 19.3944
R7794 GND.n3145 GND.n3144 19.3944
R7795 GND.n3144 GND.n3103 19.3944
R7796 GND.n3134 GND.n3103 19.3944
R7797 GND.n3134 GND.n3133 19.3944
R7798 GND.n3133 GND.n3110 19.3944
R7799 GND.n3126 GND.n3110 19.3944
R7800 GND.n3126 GND.n3125 19.3944
R7801 GND.n3125 GND.n3124 19.3944
R7802 GND.n3767 GND.n3765 19.3944
R7803 GND.n3768 GND.n3767 19.3944
R7804 GND.n3770 GND.n3768 19.3944
R7805 GND.n3770 GND.n3502 19.3944
R7806 GND.n3814 GND.n3502 19.3944
R7807 GND.n3814 GND.n3503 19.3944
R7808 GND.n3805 GND.n3503 19.3944
R7809 GND.n3807 GND.n3805 19.3944
R7810 GND.n3807 GND.n3473 19.3944
R7811 GND.n3851 GND.n3473 19.3944
R7812 GND.n3851 GND.n3474 19.3944
R7813 GND.n3842 GND.n3474 19.3944
R7814 GND.n3844 GND.n3842 19.3944
R7815 GND.n3844 GND.n3444 19.3944
R7816 GND.n3891 GND.n3444 19.3944
R7817 GND.n3891 GND.n3445 19.3944
R7818 GND.n3445 GND.n3428 19.3944
R7819 GND.n3905 GND.n3428 19.3944
R7820 GND.n3906 GND.n3905 19.3944
R7821 GND.n3906 GND.n3422 19.3944
R7822 GND.n3979 GND.n3422 19.3944
R7823 GND.n3979 GND.n3423 19.3944
R7824 GND.n3915 GND.n3423 19.3944
R7825 GND.n3916 GND.n3915 19.3944
R7826 GND.n3917 GND.n3916 19.3944
R7827 GND.n3925 GND.n3917 19.3944
R7828 GND.n3927 GND.n3925 19.3944
R7829 GND.n3927 GND.n3389 19.3944
R7830 GND.n4011 GND.n3389 19.3944
R7831 GND.n4011 GND.n3390 19.3944
R7832 GND.n4002 GND.n3390 19.3944
R7833 GND.n4004 GND.n4002 19.3944
R7834 GND.n4004 GND.n3361 19.3944
R7835 GND.n4048 GND.n3361 19.3944
R7836 GND.n4048 GND.n3362 19.3944
R7837 GND.n4039 GND.n3362 19.3944
R7838 GND.n4041 GND.n4039 19.3944
R7839 GND.n4041 GND.n3332 19.3944
R7840 GND.n4085 GND.n3332 19.3944
R7841 GND.n4085 GND.n3333 19.3944
R7842 GND.n4076 GND.n3333 19.3944
R7843 GND.n4078 GND.n4076 19.3944
R7844 GND.n4078 GND.n3303 19.3944
R7845 GND.n4140 GND.n3303 19.3944
R7846 GND.n4140 GND.n3304 19.3944
R7847 GND.n3304 GND.n3292 19.3944
R7848 GND.n3292 GND.n3170 19.3944
R7849 GND.n3776 GND.n3535 19.3944
R7850 GND.n3772 GND.n3535 19.3944
R7851 GND.n3772 GND.n3506 19.3944
R7852 GND.n3803 GND.n3506 19.3944
R7853 GND.n3812 GND.n3803 19.3944
R7854 GND.n3812 GND.n3811 19.3944
R7855 GND.n3811 GND.n3810 19.3944
R7856 GND.n3810 GND.n3477 19.3944
R7857 GND.n3840 GND.n3477 19.3944
R7858 GND.n3849 GND.n3840 19.3944
R7859 GND.n3849 GND.n3848 19.3944
R7860 GND.n3848 GND.n3847 19.3944
R7861 GND.n3847 GND.n3448 19.3944
R7862 GND.n3883 GND.n3448 19.3944
R7863 GND.n3889 GND.n3883 19.3944
R7864 GND.n3889 GND.n3888 19.3944
R7865 GND.n3888 GND.n3887 19.3944
R7866 GND.n3887 GND.n3426 19.3944
R7867 GND.n3908 GND.n3426 19.3944
R7868 GND.n3911 GND.n3908 19.3944
R7869 GND.n3977 GND.n3911 19.3944
R7870 GND.n3977 GND.n3976 19.3944
R7871 GND.n3976 GND.n3975 19.3944
R7872 GND.n3975 GND.n3914 19.3944
R7873 GND.n3971 GND.n3914 19.3944
R7874 GND.n3971 GND.n3970 19.3944
R7875 GND.n3970 GND.n3393 19.3944
R7876 GND.n4000 GND.n3393 19.3944
R7877 GND.n4009 GND.n4000 19.3944
R7878 GND.n4009 GND.n4008 19.3944
R7879 GND.n4008 GND.n4007 19.3944
R7880 GND.n4007 GND.n3365 19.3944
R7881 GND.n4037 GND.n3365 19.3944
R7882 GND.n4046 GND.n4037 19.3944
R7883 GND.n4046 GND.n4045 19.3944
R7884 GND.n4045 GND.n4044 19.3944
R7885 GND.n4044 GND.n3336 19.3944
R7886 GND.n4074 GND.n3336 19.3944
R7887 GND.n4083 GND.n4074 19.3944
R7888 GND.n4083 GND.n4082 19.3944
R7889 GND.n4082 GND.n4081 19.3944
R7890 GND.n4081 GND.n3307 19.3944
R7891 GND.n4134 GND.n3307 19.3944
R7892 GND.n4138 GND.n4134 19.3944
R7893 GND.n4138 GND.n4137 19.3944
R7894 GND.n4137 GND.n3171 19.3944
R7895 GND.n4156 GND.n3171 19.3944
R7896 GND.n6271 GND.n1515 19.3944
R7897 GND.n6267 GND.n1515 19.3944
R7898 GND.n6267 GND.n6266 19.3944
R7899 GND.n6266 GND.n6265 19.3944
R7900 GND.n6265 GND.n1522 19.3944
R7901 GND.n6261 GND.n1522 19.3944
R7902 GND.n6261 GND.n6260 19.3944
R7903 GND.n6260 GND.n6259 19.3944
R7904 GND.n6259 GND.n1528 19.3944
R7905 GND.n6255 GND.n1528 19.3944
R7906 GND.n6255 GND.n6254 19.3944
R7907 GND.n6254 GND.n6253 19.3944
R7908 GND.n6253 GND.n1534 19.3944
R7909 GND.n6249 GND.n1534 19.3944
R7910 GND.n6249 GND.n6248 19.3944
R7911 GND.n6246 GND.n1543 19.3944
R7912 GND.n6242 GND.n1543 19.3944
R7913 GND.n6242 GND.n6241 19.3944
R7914 GND.n6241 GND.n6240 19.3944
R7915 GND.n6240 GND.n1549 19.3944
R7916 GND.n6236 GND.n1549 19.3944
R7917 GND.n6236 GND.n6235 19.3944
R7918 GND.n6235 GND.n6234 19.3944
R7919 GND.n6234 GND.n1555 19.3944
R7920 GND.n6230 GND.n1555 19.3944
R7921 GND.n6230 GND.n6229 19.3944
R7922 GND.n6229 GND.n6228 19.3944
R7923 GND.n6228 GND.n1561 19.3944
R7924 GND.n6224 GND.n1561 19.3944
R7925 GND.n6224 GND.n6223 19.3944
R7926 GND.n6223 GND.n6222 19.3944
R7927 GND.n3213 GND.n1568 19.3944
R7928 GND.n3216 GND.n3213 19.3944
R7929 GND.n3216 GND.n3208 19.3944
R7930 GND.n3220 GND.n3208 19.3944
R7931 GND.n3221 GND.n3220 19.3944
R7932 GND.n3224 GND.n3221 19.3944
R7933 GND.n3224 GND.n3204 19.3944
R7934 GND.n3228 GND.n3204 19.3944
R7935 GND.n3229 GND.n3228 19.3944
R7936 GND.n3232 GND.n3229 19.3944
R7937 GND.n3232 GND.n3200 19.3944
R7938 GND.n3236 GND.n3200 19.3944
R7939 GND.n3237 GND.n3236 19.3944
R7940 GND.n3240 GND.n3237 19.3944
R7941 GND.n3240 GND.n3196 19.3944
R7942 GND.n3244 GND.n3196 19.3944
R7943 GND.n3245 GND.n3244 19.3944
R7944 GND.n3248 GND.n3189 19.3944
R7945 GND.n3252 GND.n3189 19.3944
R7946 GND.n3253 GND.n3252 19.3944
R7947 GND.n3256 GND.n3253 19.3944
R7948 GND.n3256 GND.n3185 19.3944
R7949 GND.n3260 GND.n3185 19.3944
R7950 GND.n3261 GND.n3260 19.3944
R7951 GND.n3264 GND.n3261 19.3944
R7952 GND.n3264 GND.n3181 19.3944
R7953 GND.n3268 GND.n3181 19.3944
R7954 GND.n3269 GND.n3268 19.3944
R7955 GND.n3272 GND.n3269 19.3944
R7956 GND.n3272 GND.n3177 19.3944
R7957 GND.n3276 GND.n3177 19.3944
R7958 GND.n3277 GND.n3276 19.3944
R7959 GND.n3280 GND.n3277 19.3944
R7960 GND.n3280 GND.n3173 19.3944
R7961 GND.n7597 GND.n506 19.3944
R7962 GND.n7597 GND.n504 19.3944
R7963 GND.n7601 GND.n504 19.3944
R7964 GND.n7601 GND.n500 19.3944
R7965 GND.n7607 GND.n500 19.3944
R7966 GND.n7607 GND.n498 19.3944
R7967 GND.n7611 GND.n498 19.3944
R7968 GND.n7611 GND.n494 19.3944
R7969 GND.n7617 GND.n494 19.3944
R7970 GND.n7617 GND.n492 19.3944
R7971 GND.n7621 GND.n492 19.3944
R7972 GND.n7621 GND.n488 19.3944
R7973 GND.n7627 GND.n488 19.3944
R7974 GND.n7627 GND.n486 19.3944
R7975 GND.n7631 GND.n486 19.3944
R7976 GND.n7631 GND.n482 19.3944
R7977 GND.n7637 GND.n482 19.3944
R7978 GND.n7637 GND.n480 19.3944
R7979 GND.n7641 GND.n480 19.3944
R7980 GND.n7641 GND.n476 19.3944
R7981 GND.n7647 GND.n476 19.3944
R7982 GND.n7647 GND.n474 19.3944
R7983 GND.n7651 GND.n474 19.3944
R7984 GND.n7651 GND.n470 19.3944
R7985 GND.n7657 GND.n470 19.3944
R7986 GND.n7657 GND.n468 19.3944
R7987 GND.n7661 GND.n468 19.3944
R7988 GND.n7661 GND.n464 19.3944
R7989 GND.n7667 GND.n464 19.3944
R7990 GND.n7667 GND.n462 19.3944
R7991 GND.n7671 GND.n462 19.3944
R7992 GND.n7671 GND.n458 19.3944
R7993 GND.n7677 GND.n458 19.3944
R7994 GND.n7677 GND.n456 19.3944
R7995 GND.n7681 GND.n456 19.3944
R7996 GND.n7681 GND.n452 19.3944
R7997 GND.n7687 GND.n452 19.3944
R7998 GND.n7687 GND.n450 19.3944
R7999 GND.n7691 GND.n450 19.3944
R8000 GND.n7691 GND.n446 19.3944
R8001 GND.n7697 GND.n446 19.3944
R8002 GND.n7697 GND.n444 19.3944
R8003 GND.n7701 GND.n444 19.3944
R8004 GND.n7701 GND.n440 19.3944
R8005 GND.n7707 GND.n440 19.3944
R8006 GND.n7707 GND.n438 19.3944
R8007 GND.n7711 GND.n438 19.3944
R8008 GND.n7711 GND.n434 19.3944
R8009 GND.n7717 GND.n434 19.3944
R8010 GND.n7717 GND.n432 19.3944
R8011 GND.n7721 GND.n432 19.3944
R8012 GND.n7721 GND.n428 19.3944
R8013 GND.n7727 GND.n428 19.3944
R8014 GND.n7727 GND.n426 19.3944
R8015 GND.n7731 GND.n426 19.3944
R8016 GND.n7731 GND.n422 19.3944
R8017 GND.n7737 GND.n422 19.3944
R8018 GND.n7737 GND.n420 19.3944
R8019 GND.n7742 GND.n420 19.3944
R8020 GND.n7742 GND.n416 19.3944
R8021 GND.n7748 GND.n416 19.3944
R8022 GND.n7749 GND.n7748 19.3944
R8023 GND.n6631 GND.n1086 19.3944
R8024 GND.n6631 GND.n1082 19.3944
R8025 GND.n6637 GND.n1082 19.3944
R8026 GND.n6637 GND.n1080 19.3944
R8027 GND.n6641 GND.n1080 19.3944
R8028 GND.n6641 GND.n1076 19.3944
R8029 GND.n6647 GND.n1076 19.3944
R8030 GND.n6647 GND.n1074 19.3944
R8031 GND.n6651 GND.n1074 19.3944
R8032 GND.n6651 GND.n1070 19.3944
R8033 GND.n6657 GND.n1070 19.3944
R8034 GND.n6657 GND.n1068 19.3944
R8035 GND.n6661 GND.n1068 19.3944
R8036 GND.n6661 GND.n1064 19.3944
R8037 GND.n6667 GND.n1064 19.3944
R8038 GND.n6667 GND.n1062 19.3944
R8039 GND.n6671 GND.n1062 19.3944
R8040 GND.n6671 GND.n1058 19.3944
R8041 GND.n6677 GND.n1058 19.3944
R8042 GND.n6677 GND.n1056 19.3944
R8043 GND.n6681 GND.n1056 19.3944
R8044 GND.n6681 GND.n1052 19.3944
R8045 GND.n6687 GND.n1052 19.3944
R8046 GND.n6687 GND.n1050 19.3944
R8047 GND.n6691 GND.n1050 19.3944
R8048 GND.n6691 GND.n1046 19.3944
R8049 GND.n6697 GND.n1046 19.3944
R8050 GND.n6697 GND.n1044 19.3944
R8051 GND.n6701 GND.n1044 19.3944
R8052 GND.n6701 GND.n1040 19.3944
R8053 GND.n6707 GND.n1040 19.3944
R8054 GND.n6707 GND.n1038 19.3944
R8055 GND.n6711 GND.n1038 19.3944
R8056 GND.n6711 GND.n1034 19.3944
R8057 GND.n6717 GND.n1034 19.3944
R8058 GND.n6717 GND.n1032 19.3944
R8059 GND.n6721 GND.n1032 19.3944
R8060 GND.n6721 GND.n1028 19.3944
R8061 GND.n6727 GND.n1028 19.3944
R8062 GND.n6727 GND.n1026 19.3944
R8063 GND.n6731 GND.n1026 19.3944
R8064 GND.n6731 GND.n1022 19.3944
R8065 GND.n6737 GND.n1022 19.3944
R8066 GND.n6737 GND.n1020 19.3944
R8067 GND.n6741 GND.n1020 19.3944
R8068 GND.n6741 GND.n1016 19.3944
R8069 GND.n6747 GND.n1016 19.3944
R8070 GND.n6747 GND.n1014 19.3944
R8071 GND.n6751 GND.n1014 19.3944
R8072 GND.n6751 GND.n1010 19.3944
R8073 GND.n6757 GND.n1010 19.3944
R8074 GND.n6757 GND.n1008 19.3944
R8075 GND.n6761 GND.n1008 19.3944
R8076 GND.n6761 GND.n1004 19.3944
R8077 GND.n6767 GND.n1004 19.3944
R8078 GND.n6767 GND.n1002 19.3944
R8079 GND.n6771 GND.n1002 19.3944
R8080 GND.n6771 GND.n998 19.3944
R8081 GND.n6777 GND.n998 19.3944
R8082 GND.n6777 GND.n996 19.3944
R8083 GND.n6781 GND.n996 19.3944
R8084 GND.n6781 GND.n992 19.3944
R8085 GND.n6787 GND.n992 19.3944
R8086 GND.n6787 GND.n990 19.3944
R8087 GND.n6791 GND.n990 19.3944
R8088 GND.n6791 GND.n986 19.3944
R8089 GND.n6797 GND.n986 19.3944
R8090 GND.n6797 GND.n984 19.3944
R8091 GND.n6801 GND.n984 19.3944
R8092 GND.n6801 GND.n980 19.3944
R8093 GND.n6807 GND.n980 19.3944
R8094 GND.n6807 GND.n978 19.3944
R8095 GND.n6811 GND.n978 19.3944
R8096 GND.n6811 GND.n974 19.3944
R8097 GND.n6817 GND.n974 19.3944
R8098 GND.n6817 GND.n972 19.3944
R8099 GND.n6821 GND.n972 19.3944
R8100 GND.n6821 GND.n968 19.3944
R8101 GND.n6827 GND.n968 19.3944
R8102 GND.n6827 GND.n966 19.3944
R8103 GND.n6831 GND.n966 19.3944
R8104 GND.n6831 GND.n962 19.3944
R8105 GND.n6837 GND.n962 19.3944
R8106 GND.n6837 GND.n960 19.3944
R8107 GND.n6841 GND.n960 19.3944
R8108 GND.n6841 GND.n956 19.3944
R8109 GND.n6847 GND.n956 19.3944
R8110 GND.n6847 GND.n954 19.3944
R8111 GND.n6851 GND.n954 19.3944
R8112 GND.n6851 GND.n950 19.3944
R8113 GND.n6857 GND.n950 19.3944
R8114 GND.n6857 GND.n948 19.3944
R8115 GND.n6861 GND.n948 19.3944
R8116 GND.n6861 GND.n944 19.3944
R8117 GND.n6867 GND.n944 19.3944
R8118 GND.n6867 GND.n942 19.3944
R8119 GND.n6871 GND.n942 19.3944
R8120 GND.n6871 GND.n938 19.3944
R8121 GND.n6877 GND.n938 19.3944
R8122 GND.n6877 GND.n936 19.3944
R8123 GND.n6881 GND.n936 19.3944
R8124 GND.n6881 GND.n932 19.3944
R8125 GND.n6887 GND.n932 19.3944
R8126 GND.n6887 GND.n930 19.3944
R8127 GND.n6891 GND.n930 19.3944
R8128 GND.n6891 GND.n926 19.3944
R8129 GND.n6897 GND.n926 19.3944
R8130 GND.n6897 GND.n924 19.3944
R8131 GND.n6901 GND.n924 19.3944
R8132 GND.n6901 GND.n920 19.3944
R8133 GND.n6907 GND.n920 19.3944
R8134 GND.n6907 GND.n918 19.3944
R8135 GND.n6911 GND.n918 19.3944
R8136 GND.n6911 GND.n914 19.3944
R8137 GND.n6917 GND.n914 19.3944
R8138 GND.n6917 GND.n912 19.3944
R8139 GND.n6921 GND.n912 19.3944
R8140 GND.n6921 GND.n908 19.3944
R8141 GND.n6927 GND.n908 19.3944
R8142 GND.n6927 GND.n906 19.3944
R8143 GND.n6931 GND.n906 19.3944
R8144 GND.n6931 GND.n902 19.3944
R8145 GND.n6937 GND.n902 19.3944
R8146 GND.n6937 GND.n900 19.3944
R8147 GND.n6941 GND.n900 19.3944
R8148 GND.n6941 GND.n896 19.3944
R8149 GND.n6947 GND.n896 19.3944
R8150 GND.n6947 GND.n894 19.3944
R8151 GND.n6951 GND.n894 19.3944
R8152 GND.n6951 GND.n890 19.3944
R8153 GND.n6957 GND.n890 19.3944
R8154 GND.n6957 GND.n888 19.3944
R8155 GND.n6961 GND.n888 19.3944
R8156 GND.n6961 GND.n884 19.3944
R8157 GND.n6967 GND.n884 19.3944
R8158 GND.n6967 GND.n882 19.3944
R8159 GND.n6971 GND.n882 19.3944
R8160 GND.n6971 GND.n878 19.3944
R8161 GND.n6977 GND.n878 19.3944
R8162 GND.n6977 GND.n876 19.3944
R8163 GND.n6981 GND.n876 19.3944
R8164 GND.n6981 GND.n872 19.3944
R8165 GND.n6987 GND.n872 19.3944
R8166 GND.n6987 GND.n870 19.3944
R8167 GND.n6991 GND.n870 19.3944
R8168 GND.n6991 GND.n866 19.3944
R8169 GND.n6997 GND.n866 19.3944
R8170 GND.n6997 GND.n864 19.3944
R8171 GND.n7001 GND.n864 19.3944
R8172 GND.n7001 GND.n860 19.3944
R8173 GND.n7007 GND.n860 19.3944
R8174 GND.n7007 GND.n858 19.3944
R8175 GND.n7011 GND.n858 19.3944
R8176 GND.n7011 GND.n854 19.3944
R8177 GND.n7017 GND.n854 19.3944
R8178 GND.n7017 GND.n852 19.3944
R8179 GND.n7021 GND.n852 19.3944
R8180 GND.n7021 GND.n848 19.3944
R8181 GND.n7027 GND.n848 19.3944
R8182 GND.n7027 GND.n846 19.3944
R8183 GND.n7031 GND.n846 19.3944
R8184 GND.n7031 GND.n842 19.3944
R8185 GND.n7037 GND.n842 19.3944
R8186 GND.n7037 GND.n840 19.3944
R8187 GND.n7041 GND.n840 19.3944
R8188 GND.n7041 GND.n836 19.3944
R8189 GND.n7047 GND.n836 19.3944
R8190 GND.n7047 GND.n834 19.3944
R8191 GND.n7051 GND.n834 19.3944
R8192 GND.n7051 GND.n830 19.3944
R8193 GND.n7057 GND.n830 19.3944
R8194 GND.n7057 GND.n828 19.3944
R8195 GND.n7061 GND.n828 19.3944
R8196 GND.n7061 GND.n824 19.3944
R8197 GND.n7067 GND.n824 19.3944
R8198 GND.n7067 GND.n822 19.3944
R8199 GND.n7071 GND.n822 19.3944
R8200 GND.n7071 GND.n818 19.3944
R8201 GND.n7077 GND.n818 19.3944
R8202 GND.n7077 GND.n816 19.3944
R8203 GND.n7081 GND.n816 19.3944
R8204 GND.n7081 GND.n812 19.3944
R8205 GND.n7087 GND.n812 19.3944
R8206 GND.n7087 GND.n810 19.3944
R8207 GND.n7091 GND.n810 19.3944
R8208 GND.n7091 GND.n806 19.3944
R8209 GND.n7097 GND.n806 19.3944
R8210 GND.n7097 GND.n804 19.3944
R8211 GND.n7101 GND.n804 19.3944
R8212 GND.n7101 GND.n800 19.3944
R8213 GND.n7107 GND.n800 19.3944
R8214 GND.n7107 GND.n798 19.3944
R8215 GND.n7111 GND.n798 19.3944
R8216 GND.n7111 GND.n794 19.3944
R8217 GND.n7117 GND.n794 19.3944
R8218 GND.n7117 GND.n792 19.3944
R8219 GND.n7121 GND.n792 19.3944
R8220 GND.n7121 GND.n788 19.3944
R8221 GND.n7127 GND.n788 19.3944
R8222 GND.n7127 GND.n786 19.3944
R8223 GND.n7131 GND.n786 19.3944
R8224 GND.n7131 GND.n782 19.3944
R8225 GND.n7137 GND.n782 19.3944
R8226 GND.n7137 GND.n780 19.3944
R8227 GND.n7141 GND.n780 19.3944
R8228 GND.n7141 GND.n776 19.3944
R8229 GND.n7147 GND.n776 19.3944
R8230 GND.n7147 GND.n774 19.3944
R8231 GND.n7151 GND.n774 19.3944
R8232 GND.n7151 GND.n770 19.3944
R8233 GND.n7157 GND.n770 19.3944
R8234 GND.n7157 GND.n768 19.3944
R8235 GND.n7161 GND.n768 19.3944
R8236 GND.n7161 GND.n764 19.3944
R8237 GND.n7167 GND.n764 19.3944
R8238 GND.n7167 GND.n762 19.3944
R8239 GND.n7171 GND.n762 19.3944
R8240 GND.n7171 GND.n758 19.3944
R8241 GND.n7177 GND.n758 19.3944
R8242 GND.n7177 GND.n756 19.3944
R8243 GND.n7181 GND.n756 19.3944
R8244 GND.n7181 GND.n752 19.3944
R8245 GND.n7187 GND.n752 19.3944
R8246 GND.n7187 GND.n750 19.3944
R8247 GND.n7191 GND.n750 19.3944
R8248 GND.n7191 GND.n746 19.3944
R8249 GND.n7197 GND.n746 19.3944
R8250 GND.n7197 GND.n744 19.3944
R8251 GND.n7201 GND.n744 19.3944
R8252 GND.n7201 GND.n740 19.3944
R8253 GND.n7207 GND.n740 19.3944
R8254 GND.n7207 GND.n738 19.3944
R8255 GND.n7211 GND.n738 19.3944
R8256 GND.n7211 GND.n734 19.3944
R8257 GND.n7217 GND.n734 19.3944
R8258 GND.n7217 GND.n732 19.3944
R8259 GND.n7221 GND.n732 19.3944
R8260 GND.n7221 GND.n728 19.3944
R8261 GND.n7227 GND.n728 19.3944
R8262 GND.n7227 GND.n726 19.3944
R8263 GND.n7231 GND.n726 19.3944
R8264 GND.n7231 GND.n722 19.3944
R8265 GND.n7237 GND.n722 19.3944
R8266 GND.n7237 GND.n720 19.3944
R8267 GND.n7241 GND.n720 19.3944
R8268 GND.n7241 GND.n716 19.3944
R8269 GND.n7247 GND.n716 19.3944
R8270 GND.n7247 GND.n714 19.3944
R8271 GND.n7251 GND.n714 19.3944
R8272 GND.n7251 GND.n710 19.3944
R8273 GND.n7257 GND.n710 19.3944
R8274 GND.n7257 GND.n708 19.3944
R8275 GND.n7261 GND.n708 19.3944
R8276 GND.n7261 GND.n704 19.3944
R8277 GND.n7267 GND.n704 19.3944
R8278 GND.n7267 GND.n702 19.3944
R8279 GND.n7271 GND.n702 19.3944
R8280 GND.n7271 GND.n698 19.3944
R8281 GND.n7277 GND.n698 19.3944
R8282 GND.n7277 GND.n696 19.3944
R8283 GND.n7281 GND.n696 19.3944
R8284 GND.n7281 GND.n692 19.3944
R8285 GND.n7287 GND.n692 19.3944
R8286 GND.n7287 GND.n690 19.3944
R8287 GND.n7291 GND.n690 19.3944
R8288 GND.n7291 GND.n686 19.3944
R8289 GND.n7297 GND.n686 19.3944
R8290 GND.n7297 GND.n684 19.3944
R8291 GND.n7301 GND.n684 19.3944
R8292 GND.n7301 GND.n680 19.3944
R8293 GND.n7307 GND.n680 19.3944
R8294 GND.n7307 GND.n678 19.3944
R8295 GND.n7311 GND.n678 19.3944
R8296 GND.n7311 GND.n674 19.3944
R8297 GND.n7317 GND.n674 19.3944
R8298 GND.n7317 GND.n672 19.3944
R8299 GND.n7321 GND.n672 19.3944
R8300 GND.n7321 GND.n668 19.3944
R8301 GND.n7327 GND.n668 19.3944
R8302 GND.n7327 GND.n666 19.3944
R8303 GND.n7331 GND.n666 19.3944
R8304 GND.n7331 GND.n662 19.3944
R8305 GND.n7337 GND.n662 19.3944
R8306 GND.n7337 GND.n660 19.3944
R8307 GND.n7341 GND.n660 19.3944
R8308 GND.n7341 GND.n656 19.3944
R8309 GND.n7347 GND.n656 19.3944
R8310 GND.n7347 GND.n654 19.3944
R8311 GND.n7351 GND.n654 19.3944
R8312 GND.n7351 GND.n650 19.3944
R8313 GND.n7357 GND.n650 19.3944
R8314 GND.n7357 GND.n648 19.3944
R8315 GND.n7361 GND.n648 19.3944
R8316 GND.n7361 GND.n644 19.3944
R8317 GND.n7367 GND.n644 19.3944
R8318 GND.n7367 GND.n642 19.3944
R8319 GND.n7371 GND.n642 19.3944
R8320 GND.n7371 GND.n638 19.3944
R8321 GND.n7377 GND.n638 19.3944
R8322 GND.n7377 GND.n636 19.3944
R8323 GND.n7381 GND.n636 19.3944
R8324 GND.n7381 GND.n632 19.3944
R8325 GND.n7387 GND.n632 19.3944
R8326 GND.n7387 GND.n630 19.3944
R8327 GND.n7391 GND.n630 19.3944
R8328 GND.n7391 GND.n626 19.3944
R8329 GND.n7397 GND.n626 19.3944
R8330 GND.n7397 GND.n624 19.3944
R8331 GND.n7401 GND.n624 19.3944
R8332 GND.n7401 GND.n620 19.3944
R8333 GND.n7407 GND.n620 19.3944
R8334 GND.n7407 GND.n618 19.3944
R8335 GND.n7411 GND.n618 19.3944
R8336 GND.n7411 GND.n614 19.3944
R8337 GND.n7417 GND.n614 19.3944
R8338 GND.n7417 GND.n612 19.3944
R8339 GND.n7421 GND.n612 19.3944
R8340 GND.n7421 GND.n608 19.3944
R8341 GND.n7427 GND.n608 19.3944
R8342 GND.n7427 GND.n606 19.3944
R8343 GND.n7431 GND.n606 19.3944
R8344 GND.n7431 GND.n602 19.3944
R8345 GND.n7437 GND.n602 19.3944
R8346 GND.n7437 GND.n600 19.3944
R8347 GND.n7441 GND.n600 19.3944
R8348 GND.n7441 GND.n596 19.3944
R8349 GND.n7447 GND.n596 19.3944
R8350 GND.n7447 GND.n594 19.3944
R8351 GND.n7451 GND.n594 19.3944
R8352 GND.n7451 GND.n590 19.3944
R8353 GND.n7457 GND.n590 19.3944
R8354 GND.n7457 GND.n588 19.3944
R8355 GND.n7461 GND.n588 19.3944
R8356 GND.n7461 GND.n584 19.3944
R8357 GND.n7467 GND.n584 19.3944
R8358 GND.n7467 GND.n582 19.3944
R8359 GND.n7471 GND.n582 19.3944
R8360 GND.n7471 GND.n578 19.3944
R8361 GND.n7477 GND.n578 19.3944
R8362 GND.n7477 GND.n576 19.3944
R8363 GND.n7481 GND.n576 19.3944
R8364 GND.n7481 GND.n572 19.3944
R8365 GND.n7487 GND.n572 19.3944
R8366 GND.n7487 GND.n570 19.3944
R8367 GND.n7491 GND.n570 19.3944
R8368 GND.n7491 GND.n566 19.3944
R8369 GND.n7497 GND.n566 19.3944
R8370 GND.n7497 GND.n564 19.3944
R8371 GND.n7501 GND.n564 19.3944
R8372 GND.n7501 GND.n560 19.3944
R8373 GND.n7507 GND.n560 19.3944
R8374 GND.n7507 GND.n558 19.3944
R8375 GND.n7511 GND.n558 19.3944
R8376 GND.n7511 GND.n554 19.3944
R8377 GND.n7517 GND.n554 19.3944
R8378 GND.n7517 GND.n552 19.3944
R8379 GND.n7521 GND.n552 19.3944
R8380 GND.n7521 GND.n548 19.3944
R8381 GND.n7527 GND.n548 19.3944
R8382 GND.n7527 GND.n546 19.3944
R8383 GND.n7531 GND.n546 19.3944
R8384 GND.n7531 GND.n542 19.3944
R8385 GND.n7537 GND.n542 19.3944
R8386 GND.n7537 GND.n540 19.3944
R8387 GND.n7541 GND.n540 19.3944
R8388 GND.n7541 GND.n536 19.3944
R8389 GND.n7547 GND.n536 19.3944
R8390 GND.n7547 GND.n534 19.3944
R8391 GND.n7551 GND.n534 19.3944
R8392 GND.n7551 GND.n530 19.3944
R8393 GND.n7557 GND.n530 19.3944
R8394 GND.n7557 GND.n528 19.3944
R8395 GND.n7561 GND.n528 19.3944
R8396 GND.n7561 GND.n524 19.3944
R8397 GND.n7567 GND.n524 19.3944
R8398 GND.n7567 GND.n522 19.3944
R8399 GND.n7571 GND.n522 19.3944
R8400 GND.n7571 GND.n518 19.3944
R8401 GND.n7577 GND.n518 19.3944
R8402 GND.n7577 GND.n516 19.3944
R8403 GND.n7581 GND.n516 19.3944
R8404 GND.n7581 GND.n512 19.3944
R8405 GND.n7587 GND.n512 19.3944
R8406 GND.n7587 GND.n510 19.3944
R8407 GND.n7591 GND.n510 19.3944
R8408 GND.n5585 GND.n5584 19.3944
R8409 GND.n5584 GND.n5583 19.3944
R8410 GND.n5583 GND.n5582 19.3944
R8411 GND.n5582 GND.n5580 19.3944
R8412 GND.n5580 GND.n5577 19.3944
R8413 GND.n5577 GND.n5576 19.3944
R8414 GND.n5576 GND.n5573 19.3944
R8415 GND.n5573 GND.n5572 19.3944
R8416 GND.n5572 GND.n5569 19.3944
R8417 GND.n5569 GND.n5568 19.3944
R8418 GND.n5568 GND.n5565 19.3944
R8419 GND.n5565 GND.n5564 19.3944
R8420 GND.n5564 GND.n5561 19.3944
R8421 GND.n5561 GND.n5560 19.3944
R8422 GND.n5560 GND.n5557 19.3944
R8423 GND.n5555 GND.n5553 19.3944
R8424 GND.n5553 GND.n5550 19.3944
R8425 GND.n5550 GND.n5549 19.3944
R8426 GND.n5549 GND.n5546 19.3944
R8427 GND.n5546 GND.n5545 19.3944
R8428 GND.n5545 GND.n5542 19.3944
R8429 GND.n5542 GND.n5541 19.3944
R8430 GND.n5541 GND.n5538 19.3944
R8431 GND.n5538 GND.n5537 19.3944
R8432 GND.n5537 GND.n5534 19.3944
R8433 GND.n5534 GND.n5533 19.3944
R8434 GND.n5533 GND.n5530 19.3944
R8435 GND.n5530 GND.n5529 19.3944
R8436 GND.n5529 GND.n5526 19.3944
R8437 GND.n5526 GND.n5525 19.3944
R8438 GND.n5525 GND.n5522 19.3944
R8439 GND.n5520 GND.n5517 19.3944
R8440 GND.n5517 GND.n5516 19.3944
R8441 GND.n5516 GND.n5513 19.3944
R8442 GND.n5513 GND.n5512 19.3944
R8443 GND.n5512 GND.n5509 19.3944
R8444 GND.n5509 GND.n5508 19.3944
R8445 GND.n5508 GND.n5505 19.3944
R8446 GND.n5505 GND.n5504 19.3944
R8447 GND.n5504 GND.n5501 19.3944
R8448 GND.n5501 GND.n5500 19.3944
R8449 GND.n5500 GND.n5497 19.3944
R8450 GND.n5497 GND.n5496 19.3944
R8451 GND.n5496 GND.n5493 19.3944
R8452 GND.n5493 GND.n5492 19.3944
R8453 GND.n5492 GND.n5489 19.3944
R8454 GND.n5489 GND.n5488 19.3944
R8455 GND.n5488 GND.n5485 19.3944
R8456 GND.n5483 GND.n5480 19.3944
R8457 GND.n5480 GND.n5479 19.3944
R8458 GND.n5479 GND.n5476 19.3944
R8459 GND.n5476 GND.n5475 19.3944
R8460 GND.n5475 GND.n5472 19.3944
R8461 GND.n5472 GND.n5471 19.3944
R8462 GND.n5471 GND.n5468 19.3944
R8463 GND.n5468 GND.n5467 19.3944
R8464 GND.n5467 GND.n5464 19.3944
R8465 GND.n5464 GND.n5463 19.3944
R8466 GND.n5463 GND.n5460 19.3944
R8467 GND.n5460 GND.n5459 19.3944
R8468 GND.n5459 GND.n5456 19.3944
R8469 GND.n5456 GND.n5455 19.3944
R8470 GND.n5455 GND.n5452 19.3944
R8471 GND.n5452 GND.n5451 19.3944
R8472 GND.n5451 GND.n5448 19.3944
R8473 GND.n5441 GND.n2402 19.3944
R8474 GND.n5048 GND.n2402 19.3944
R8475 GND.n5048 GND.n2658 19.3944
R8476 GND.n5060 GND.n2658 19.3944
R8477 GND.n5061 GND.n5060 19.3944
R8478 GND.n5063 GND.n5061 19.3944
R8479 GND.n5063 GND.n2574 19.3944
R8480 GND.n5075 GND.n2574 19.3944
R8481 GND.n5076 GND.n5075 19.3944
R8482 GND.n5078 GND.n5076 19.3944
R8483 GND.n5078 GND.n2570 19.3944
R8484 GND.n5090 GND.n2570 19.3944
R8485 GND.n5091 GND.n5090 19.3944
R8486 GND.n5093 GND.n5091 19.3944
R8487 GND.n5093 GND.n2566 19.3944
R8488 GND.n5105 GND.n2566 19.3944
R8489 GND.n5106 GND.n5105 19.3944
R8490 GND.n5108 GND.n5106 19.3944
R8491 GND.n5108 GND.n2562 19.3944
R8492 GND.n5124 GND.n2562 19.3944
R8493 GND.n5125 GND.n5124 19.3944
R8494 GND.n5126 GND.n5125 19.3944
R8495 GND.n5126 GND.n2561 19.3944
R8496 GND.n5133 GND.n2561 19.3944
R8497 GND.n5135 GND.n5133 19.3944
R8498 GND.n5357 GND.n5135 19.3944
R8499 GND.n5357 GND.n5356 19.3944
R8500 GND.n5356 GND.n5136 19.3944
R8501 GND.n5346 GND.n5136 19.3944
R8502 GND.n5346 GND.n5345 19.3944
R8503 GND.n5345 GND.n5344 19.3944
R8504 GND.n5344 GND.n5204 19.3944
R8505 GND.n5334 GND.n5204 19.3944
R8506 GND.n5334 GND.n5333 19.3944
R8507 GND.n5333 GND.n5332 19.3944
R8508 GND.n5332 GND.n5211 19.3944
R8509 GND.n5322 GND.n5211 19.3944
R8510 GND.n5322 GND.n5321 19.3944
R8511 GND.n5321 GND.n5320 19.3944
R8512 GND.n5320 GND.n5218 19.3944
R8513 GND.n5310 GND.n5218 19.3944
R8514 GND.n5310 GND.n5309 19.3944
R8515 GND.n5309 GND.n5308 19.3944
R8516 GND.n5308 GND.n5225 19.3944
R8517 GND.n5298 GND.n5225 19.3944
R8518 GND.n5298 GND.n287 19.3944
R8519 GND.n7877 GND.n287 19.3944
R8520 GND.n2435 GND.n2400 19.3944
R8521 GND.n2451 GND.n2435 19.3944
R8522 GND.n5428 GND.n2451 19.3944
R8523 GND.n5428 GND.n5427 19.3944
R8524 GND.n5427 GND.n5426 19.3944
R8525 GND.n5426 GND.n2455 19.3944
R8526 GND.n5416 GND.n2455 19.3944
R8527 GND.n5416 GND.n5415 19.3944
R8528 GND.n5415 GND.n5414 19.3944
R8529 GND.n5414 GND.n2475 19.3944
R8530 GND.n5404 GND.n2475 19.3944
R8531 GND.n5404 GND.n5403 19.3944
R8532 GND.n5403 GND.n5402 19.3944
R8533 GND.n5402 GND.n2496 19.3944
R8534 GND.n5392 GND.n2496 19.3944
R8535 GND.n5392 GND.n5391 19.3944
R8536 GND.n5391 GND.n5390 19.3944
R8537 GND.n5390 GND.n2517 19.3944
R8538 GND.n5380 GND.n2517 19.3944
R8539 GND.n5380 GND.n5379 19.3944
R8540 GND.n5379 GND.n5378 19.3944
R8541 GND.n5378 GND.n2536 19.3944
R8542 GND.n5130 GND.n2536 19.3944
R8543 GND.n5131 GND.n5130 19.3944
R8544 GND.n5131 GND.n2557 19.3944
R8545 GND.n5359 GND.n2557 19.3944
R8546 GND.n5359 GND.n56 19.3944
R8547 GND.n8069 GND.n56 19.3944
R8548 GND.n8069 GND.n8068 19.3944
R8549 GND.n8068 GND.n8067 19.3944
R8550 GND.n8067 GND.n60 19.3944
R8551 GND.n8057 GND.n60 19.3944
R8552 GND.n8057 GND.n8056 19.3944
R8553 GND.n8056 GND.n8055 19.3944
R8554 GND.n8055 GND.n80 19.3944
R8555 GND.n8045 GND.n80 19.3944
R8556 GND.n8045 GND.n8044 19.3944
R8557 GND.n8044 GND.n8043 19.3944
R8558 GND.n8043 GND.n101 19.3944
R8559 GND.n8033 GND.n101 19.3944
R8560 GND.n8033 GND.n8032 19.3944
R8561 GND.n8032 GND.n8031 19.3944
R8562 GND.n8031 GND.n122 19.3944
R8563 GND.n8021 GND.n122 19.3944
R8564 GND.n8021 GND.n8020 19.3944
R8565 GND.n8020 GND.n8019 19.3944
R8566 GND.n8019 GND.n143 19.3944
R8567 GND.n7911 GND.n251 19.3944
R8568 GND.n7911 GND.n7910 19.3944
R8569 GND.n7910 GND.n7909 19.3944
R8570 GND.n7909 GND.n257 19.3944
R8571 GND.n7904 GND.n257 19.3944
R8572 GND.n7904 GND.n7903 19.3944
R8573 GND.n7903 GND.n7902 19.3944
R8574 GND.n7902 GND.n264 19.3944
R8575 GND.n7897 GND.n264 19.3944
R8576 GND.n7897 GND.n7896 19.3944
R8577 GND.n7896 GND.n7895 19.3944
R8578 GND.n7895 GND.n271 19.3944
R8579 GND.n7890 GND.n271 19.3944
R8580 GND.n7890 GND.n7889 19.3944
R8581 GND.n7889 GND.n7888 19.3944
R8582 GND.n7888 GND.n278 19.3944
R8583 GND.n7883 GND.n278 19.3944
R8584 GND.n7944 GND.n213 19.3944
R8585 GND.n7944 GND.n219 19.3944
R8586 GND.n7939 GND.n219 19.3944
R8587 GND.n7939 GND.n7938 19.3944
R8588 GND.n7938 GND.n7937 19.3944
R8589 GND.n7937 GND.n226 19.3944
R8590 GND.n7932 GND.n226 19.3944
R8591 GND.n7932 GND.n7931 19.3944
R8592 GND.n7931 GND.n7930 19.3944
R8593 GND.n7930 GND.n233 19.3944
R8594 GND.n7925 GND.n233 19.3944
R8595 GND.n7925 GND.n7924 19.3944
R8596 GND.n7924 GND.n7923 19.3944
R8597 GND.n7923 GND.n240 19.3944
R8598 GND.n7918 GND.n240 19.3944
R8599 GND.n7918 GND.n7917 19.3944
R8600 GND.n7917 GND.n7916 19.3944
R8601 GND.n7978 GND.n180 19.3944
R8602 GND.n7978 GND.n184 19.3944
R8603 GND.n187 GND.n184 19.3944
R8604 GND.n7971 GND.n187 19.3944
R8605 GND.n7971 GND.n7970 19.3944
R8606 GND.n7970 GND.n7969 19.3944
R8607 GND.n7969 GND.n193 19.3944
R8608 GND.n7964 GND.n193 19.3944
R8609 GND.n7964 GND.n7963 19.3944
R8610 GND.n7963 GND.n7962 19.3944
R8611 GND.n7962 GND.n200 19.3944
R8612 GND.n7957 GND.n200 19.3944
R8613 GND.n7957 GND.n7956 19.3944
R8614 GND.n7956 GND.n7955 19.3944
R8615 GND.n7955 GND.n207 19.3944
R8616 GND.n7950 GND.n207 19.3944
R8617 GND.n7950 GND.n7949 19.3944
R8618 GND.n8011 GND.n153 19.3944
R8619 GND.n155 GND.n153 19.3944
R8620 GND.n8004 GND.n155 19.3944
R8621 GND.n8004 GND.n8003 19.3944
R8622 GND.n8003 GND.n8002 19.3944
R8623 GND.n8002 GND.n161 19.3944
R8624 GND.n7997 GND.n161 19.3944
R8625 GND.n7997 GND.n7996 19.3944
R8626 GND.n7996 GND.n7995 19.3944
R8627 GND.n7995 GND.n168 19.3944
R8628 GND.n7990 GND.n168 19.3944
R8629 GND.n7990 GND.n7989 19.3944
R8630 GND.n7989 GND.n7988 19.3944
R8631 GND.n7988 GND.n175 19.3944
R8632 GND.n7983 GND.n175 19.3944
R8633 GND.n5254 GND.n5249 19.3944
R8634 GND.n5254 GND.n5248 19.3944
R8635 GND.n5258 GND.n5248 19.3944
R8636 GND.n5258 GND.n5246 19.3944
R8637 GND.n5264 GND.n5246 19.3944
R8638 GND.n5264 GND.n5244 19.3944
R8639 GND.n5268 GND.n5244 19.3944
R8640 GND.n5268 GND.n5242 19.3944
R8641 GND.n5274 GND.n5242 19.3944
R8642 GND.n5274 GND.n5240 19.3944
R8643 GND.n5278 GND.n5240 19.3944
R8644 GND.n5278 GND.n5238 19.3944
R8645 GND.n5284 GND.n5238 19.3944
R8646 GND.n5284 GND.n5236 19.3944
R8647 GND.n5288 GND.n5236 19.3944
R8648 GND.n5046 GND.n5045 19.3944
R8649 GND.n5052 GND.n5046 19.3944
R8650 GND.n5052 GND.n2659 19.3944
R8651 GND.n5056 GND.n2659 19.3944
R8652 GND.n5056 GND.n2577 19.3944
R8653 GND.n5067 GND.n2577 19.3944
R8654 GND.n5067 GND.n2575 19.3944
R8655 GND.n5071 GND.n2575 19.3944
R8656 GND.n5071 GND.n2573 19.3944
R8657 GND.n5082 GND.n2573 19.3944
R8658 GND.n5082 GND.n2571 19.3944
R8659 GND.n5086 GND.n2571 19.3944
R8660 GND.n5086 GND.n2569 19.3944
R8661 GND.n5097 GND.n2569 19.3944
R8662 GND.n5097 GND.n2567 19.3944
R8663 GND.n5101 GND.n2567 19.3944
R8664 GND.n5101 GND.n2565 19.3944
R8665 GND.n5112 GND.n2565 19.3944
R8666 GND.n5112 GND.n2563 19.3944
R8667 GND.n5120 GND.n2563 19.3944
R8668 GND.n5120 GND.n5119 19.3944
R8669 GND.n5119 GND.n5118 19.3944
R8670 GND.n5118 GND.n28 19.3944
R8671 GND.n8080 GND.n28 19.3944
R8672 GND.n8080 GND.n29 19.3944
R8673 GND.n5137 GND.n29 19.3944
R8674 GND.n5352 GND.n5137 19.3944
R8675 GND.n5352 GND.n5351 19.3944
R8676 GND.n5351 GND.n5350 19.3944
R8677 GND.n5350 GND.n5142 19.3944
R8678 GND.n5340 GND.n5142 19.3944
R8679 GND.n5340 GND.n5339 19.3944
R8680 GND.n5339 GND.n5338 19.3944
R8681 GND.n5338 GND.n5209 19.3944
R8682 GND.n5328 GND.n5209 19.3944
R8683 GND.n5328 GND.n5327 19.3944
R8684 GND.n5327 GND.n5326 19.3944
R8685 GND.n5326 GND.n5216 19.3944
R8686 GND.n5316 GND.n5216 19.3944
R8687 GND.n5316 GND.n5315 19.3944
R8688 GND.n5315 GND.n5314 19.3944
R8689 GND.n5314 GND.n5223 19.3944
R8690 GND.n5304 GND.n5223 19.3944
R8691 GND.n5304 GND.n5303 19.3944
R8692 GND.n5303 GND.n5302 19.3944
R8693 GND.n5302 GND.n5297 19.3944
R8694 GND.n5297 GND.n5296 19.3944
R8695 GND.n2432 GND.n2431 19.3944
R8696 GND.n2431 GND.n2428 19.3944
R8697 GND.n2428 GND.n2427 19.3944
R8698 GND.n2427 GND.n2424 19.3944
R8699 GND.n2424 GND.n2423 19.3944
R8700 GND.n2423 GND.n2420 19.3944
R8701 GND.n2420 GND.n2419 19.3944
R8702 GND.n2419 GND.n2416 19.3944
R8703 GND.n2416 GND.n2264 19.3944
R8704 GND.n5591 GND.n2264 19.3944
R8705 GND.n5591 GND.n2265 19.3944
R8706 GND.n5031 GND.n2265 19.3944
R8707 GND.n5034 GND.n5031 19.3944
R8708 GND.n5034 GND.n2665 19.3944
R8709 GND.n5039 GND.n2665 19.3944
R8710 GND.n3120 GND.n3028 19.3944
R8711 GND.n4207 GND.n3028 19.3944
R8712 GND.n4207 GND.n3026 19.3944
R8713 GND.n4213 GND.n3026 19.3944
R8714 GND.n4213 GND.n4212 19.3944
R8715 GND.n4212 GND.n3005 19.3944
R8716 GND.n4239 GND.n3005 19.3944
R8717 GND.n4239 GND.n3003 19.3944
R8718 GND.n4245 GND.n3003 19.3944
R8719 GND.n4245 GND.n4244 19.3944
R8720 GND.n4244 GND.n2982 19.3944
R8721 GND.n4271 GND.n2982 19.3944
R8722 GND.n4271 GND.n2980 19.3944
R8723 GND.n4277 GND.n2980 19.3944
R8724 GND.n4277 GND.n4276 19.3944
R8725 GND.n4276 GND.n2959 19.3944
R8726 GND.n4303 GND.n2959 19.3944
R8727 GND.n4303 GND.n2957 19.3944
R8728 GND.n4309 GND.n2957 19.3944
R8729 GND.n4309 GND.n4308 19.3944
R8730 GND.n4308 GND.n2935 19.3944
R8731 GND.n4335 GND.n2935 19.3944
R8732 GND.n4335 GND.n2933 19.3944
R8733 GND.n4341 GND.n2933 19.3944
R8734 GND.n4341 GND.n4340 19.3944
R8735 GND.n4340 GND.n2913 19.3944
R8736 GND.n4367 GND.n2913 19.3944
R8737 GND.n4367 GND.n2911 19.3944
R8738 GND.n4373 GND.n2911 19.3944
R8739 GND.n4373 GND.n4372 19.3944
R8740 GND.n4372 GND.n2890 19.3944
R8741 GND.n4399 GND.n2890 19.3944
R8742 GND.n4399 GND.n2888 19.3944
R8743 GND.n4405 GND.n2888 19.3944
R8744 GND.n4405 GND.n4404 19.3944
R8745 GND.n4404 GND.n2867 19.3944
R8746 GND.n4431 GND.n2867 19.3944
R8747 GND.n4431 GND.n2865 19.3944
R8748 GND.n4437 GND.n2865 19.3944
R8749 GND.n4437 GND.n4436 19.3944
R8750 GND.n4436 GND.n2844 19.3944
R8751 GND.n4463 GND.n2844 19.3944
R8752 GND.n4463 GND.n2842 19.3944
R8753 GND.n4469 GND.n2842 19.3944
R8754 GND.n4469 GND.n4468 19.3944
R8755 GND.n4468 GND.n2821 19.3944
R8756 GND.n4495 GND.n2821 19.3944
R8757 GND.n4495 GND.n2819 19.3944
R8758 GND.n4501 GND.n2819 19.3944
R8759 GND.n4501 GND.n4500 19.3944
R8760 GND.n4500 GND.n2798 19.3944
R8761 GND.n4527 GND.n2798 19.3944
R8762 GND.n4527 GND.n2796 19.3944
R8763 GND.n4536 GND.n2796 19.3944
R8764 GND.n4536 GND.n4535 19.3944
R8765 GND.n4535 GND.n4534 19.3944
R8766 GND.n4534 GND.n2776 19.3944
R8767 GND.n2776 GND.n2774 19.3944
R8768 GND.n4655 GND.n2774 19.3944
R8769 GND.n4655 GND.n2772 19.3944
R8770 GND.n4664 GND.n2772 19.3944
R8771 GND.n4664 GND.n4663 19.3944
R8772 GND.n4663 GND.n4662 19.3944
R8773 GND.n4662 GND.n2763 19.3944
R8774 GND.n4693 GND.n2763 19.3944
R8775 GND.n4693 GND.n2761 19.3944
R8776 GND.n4712 GND.n2761 19.3944
R8777 GND.n4712 GND.n4711 19.3944
R8778 GND.n4711 GND.n4710 19.3944
R8779 GND.n4710 GND.n4699 19.3944
R8780 GND.n4706 GND.n4699 19.3944
R8781 GND.n4706 GND.n4705 19.3944
R8782 GND.n4705 GND.n2750 19.3944
R8783 GND.n4765 GND.n2750 19.3944
R8784 GND.n4766 GND.n4765 19.3944
R8785 GND.n4766 GND.n2748 19.3944
R8786 GND.n4770 GND.n2748 19.3944
R8787 GND.n4770 GND.n2746 19.3944
R8788 GND.n4774 GND.n2746 19.3944
R8789 GND.n4774 GND.n2744 19.3944
R8790 GND.n4787 GND.n2744 19.3944
R8791 GND.n4787 GND.n4786 19.3944
R8792 GND.n4786 GND.n4785 19.3944
R8793 GND.n4785 GND.n4783 19.3944
R8794 GND.n4783 GND.n4782 19.3944
R8795 GND.n4782 GND.n2727 19.3944
R8796 GND.n4859 GND.n2727 19.3944
R8797 GND.n4859 GND.n2725 19.3944
R8798 GND.n4866 GND.n2725 19.3944
R8799 GND.n4866 GND.n4865 19.3944
R8800 GND.n4865 GND.n2710 19.3944
R8801 GND.n4881 GND.n2710 19.3944
R8802 GND.n4882 GND.n4881 19.3944
R8803 GND.n4882 GND.n2708 19.3944
R8804 GND.n4886 GND.n2708 19.3944
R8805 GND.n4886 GND.n2706 19.3944
R8806 GND.n4891 GND.n2706 19.3944
R8807 GND.n4891 GND.n2704 19.3944
R8808 GND.n4895 GND.n2704 19.3944
R8809 GND.n4896 GND.n4895 19.3944
R8810 GND.n4899 GND.n4896 19.3944
R8811 GND.n4899 GND.n2702 19.3944
R8812 GND.n4905 GND.n2702 19.3944
R8813 GND.n4906 GND.n4905 19.3944
R8814 GND.n4909 GND.n4906 19.3944
R8815 GND.n4909 GND.n2700 19.3944
R8816 GND.n4913 GND.n2700 19.3944
R8817 GND.n4916 GND.n4913 19.3944
R8818 GND.n4917 GND.n4916 19.3944
R8819 GND.n4917 GND.n2698 19.3944
R8820 GND.n4923 GND.n2698 19.3944
R8821 GND.n4924 GND.n4923 19.3944
R8822 GND.n4927 GND.n4924 19.3944
R8823 GND.n4927 GND.n2696 19.3944
R8824 GND.n4931 GND.n2696 19.3944
R8825 GND.n4934 GND.n4931 19.3944
R8826 GND.n4935 GND.n4934 19.3944
R8827 GND.n4935 GND.n2694 19.3944
R8828 GND.n4939 GND.n2694 19.3944
R8829 GND.n4940 GND.n4939 19.3944
R8830 GND.n4943 GND.n4940 19.3944
R8831 GND.n4943 GND.n2689 19.3944
R8832 GND.n4949 GND.n2689 19.3944
R8833 GND.n4950 GND.n4949 19.3944
R8834 GND.n4953 GND.n4950 19.3944
R8835 GND.n4953 GND.n2687 19.3944
R8836 GND.n4957 GND.n2687 19.3944
R8837 GND.n4960 GND.n4957 19.3944
R8838 GND.n4961 GND.n4960 19.3944
R8839 GND.n4961 GND.n2685 19.3944
R8840 GND.n4967 GND.n2685 19.3944
R8841 GND.n4968 GND.n4967 19.3944
R8842 GND.n4971 GND.n4968 19.3944
R8843 GND.n4971 GND.n2683 19.3944
R8844 GND.n4975 GND.n2683 19.3944
R8845 GND.n4978 GND.n4975 19.3944
R8846 GND.n4979 GND.n4978 19.3944
R8847 GND.n4979 GND.n2681 19.3944
R8848 GND.n4983 GND.n2681 19.3944
R8849 GND.n4984 GND.n4983 19.3944
R8850 GND.n4987 GND.n4984 19.3944
R8851 GND.n4987 GND.n2677 19.3944
R8852 GND.n4993 GND.n2677 19.3944
R8853 GND.n4994 GND.n4993 19.3944
R8854 GND.n4997 GND.n4994 19.3944
R8855 GND.n4997 GND.n2675 19.3944
R8856 GND.n5001 GND.n2675 19.3944
R8857 GND.n5005 GND.n5001 19.3944
R8858 GND.n5006 GND.n5005 19.3944
R8859 GND.n5006 GND.n2673 19.3944
R8860 GND.n5012 GND.n2673 19.3944
R8861 GND.n5013 GND.n5012 19.3944
R8862 GND.n5016 GND.n5013 19.3944
R8863 GND.n5016 GND.n2671 19.3944
R8864 GND.n5020 GND.n2671 19.3944
R8865 GND.n5021 GND.n5020 19.3944
R8866 GND.n5027 GND.n2259 19.3944
R8867 GND.n5027 GND.n5024 19.3944
R8868 GND.n5641 GND.n5640 19.3944
R8869 GND.n5640 GND.n2239 19.3944
R8870 GND.n5636 GND.n2239 19.3944
R8871 GND.n5636 GND.n5633 19.3944
R8872 GND.n5633 GND.n5630 19.3944
R8873 GND.n5630 GND.n5629 19.3944
R8874 GND.n5629 GND.n5626 19.3944
R8875 GND.n5626 GND.n5625 19.3944
R8876 GND.n5625 GND.n5622 19.3944
R8877 GND.n5622 GND.n5621 19.3944
R8878 GND.n5621 GND.n5618 19.3944
R8879 GND.n5618 GND.n5617 19.3944
R8880 GND.n5617 GND.n5614 19.3944
R8881 GND.n5614 GND.n5613 19.3944
R8882 GND.n5613 GND.n5610 19.3944
R8883 GND.n5610 GND.n5609 19.3944
R8884 GND.n5609 GND.n5606 19.3944
R8885 GND.n5606 GND.n5605 19.3944
R8886 GND.n5605 GND.n5602 19.3944
R8887 GND.n5602 GND.n5601 19.3944
R8888 GND.n5601 GND.n5598 19.3944
R8889 GND.n5598 GND.n5597 19.3944
R8890 GND.n4197 GND.n3034 19.3944
R8891 GND.n4203 GND.n3034 19.3944
R8892 GND.n4203 GND.n4202 19.3944
R8893 GND.n4202 GND.n3013 19.3944
R8894 GND.n4229 GND.n3013 19.3944
R8895 GND.n4229 GND.n3011 19.3944
R8896 GND.n4235 GND.n3011 19.3944
R8897 GND.n4235 GND.n4234 19.3944
R8898 GND.n4234 GND.n2990 19.3944
R8899 GND.n4261 GND.n2990 19.3944
R8900 GND.n4261 GND.n2988 19.3944
R8901 GND.n4267 GND.n2988 19.3944
R8902 GND.n4267 GND.n4266 19.3944
R8903 GND.n4266 GND.n2967 19.3944
R8904 GND.n4293 GND.n2967 19.3944
R8905 GND.n4293 GND.n2965 19.3944
R8906 GND.n4299 GND.n2965 19.3944
R8907 GND.n4299 GND.n4298 19.3944
R8908 GND.n4298 GND.n2944 19.3944
R8909 GND.n4325 GND.n2944 19.3944
R8910 GND.n4325 GND.n2942 19.3944
R8911 GND.n4331 GND.n2942 19.3944
R8912 GND.n4331 GND.n4330 19.3944
R8913 GND.n4330 GND.n2921 19.3944
R8914 GND.n4357 GND.n2921 19.3944
R8915 GND.n4357 GND.n2919 19.3944
R8916 GND.n4363 GND.n2919 19.3944
R8917 GND.n4363 GND.n4362 19.3944
R8918 GND.n4362 GND.n2898 19.3944
R8919 GND.n4389 GND.n2898 19.3944
R8920 GND.n4389 GND.n2896 19.3944
R8921 GND.n4395 GND.n2896 19.3944
R8922 GND.n4395 GND.n4394 19.3944
R8923 GND.n4394 GND.n2875 19.3944
R8924 GND.n4421 GND.n2875 19.3944
R8925 GND.n4421 GND.n2873 19.3944
R8926 GND.n4427 GND.n2873 19.3944
R8927 GND.n4427 GND.n4426 19.3944
R8928 GND.n4426 GND.n2852 19.3944
R8929 GND.n4453 GND.n2852 19.3944
R8930 GND.n4453 GND.n2850 19.3944
R8931 GND.n4459 GND.n2850 19.3944
R8932 GND.n4459 GND.n4458 19.3944
R8933 GND.n4458 GND.n2829 19.3944
R8934 GND.n4485 GND.n2829 19.3944
R8935 GND.n4485 GND.n2827 19.3944
R8936 GND.n4491 GND.n2827 19.3944
R8937 GND.n4491 GND.n4490 19.3944
R8938 GND.n4490 GND.n2806 19.3944
R8939 GND.n4517 GND.n2806 19.3944
R8940 GND.n4517 GND.n2804 19.3944
R8941 GND.n4523 GND.n2804 19.3944
R8942 GND.n4523 GND.n4522 19.3944
R8943 GND.n4522 GND.n2783 19.3944
R8944 GND.n4568 GND.n2783 19.3944
R8945 GND.n4568 GND.n2781 19.3944
R8946 GND.n4575 GND.n2781 19.3944
R8947 GND.n4575 GND.n4574 19.3944
R8948 GND.n4574 GND.n1655 19.3944
R8949 GND.n6141 GND.n1655 19.3944
R8950 GND.n6141 GND.n6140 19.3944
R8951 GND.n6140 GND.n6139 19.3944
R8952 GND.n6139 GND.n1659 19.3944
R8953 GND.n1688 GND.n1659 19.3944
R8954 GND.n1688 GND.n1685 19.3944
R8955 GND.n6120 GND.n1685 19.3944
R8956 GND.n6120 GND.n6119 19.3944
R8957 GND.n6119 GND.n6118 19.3944
R8958 GND.n6118 GND.n1694 19.3944
R8959 GND.n1737 GND.n1694 19.3944
R8960 GND.n1740 GND.n1737 19.3944
R8961 GND.n1740 GND.n1734 19.3944
R8962 GND.n6093 GND.n1734 19.3944
R8963 GND.n6093 GND.n6092 19.3944
R8964 GND.n6092 GND.n6091 19.3944
R8965 GND.n6091 GND.n1746 19.3944
R8966 GND.n4796 GND.n1746 19.3944
R8967 GND.n4796 GND.n4793 19.3944
R8968 GND.n4800 GND.n4793 19.3944
R8969 GND.n4800 GND.n4791 19.3944
R8970 GND.n4806 GND.n4791 19.3944
R8971 GND.n4806 GND.n4805 19.3944
R8972 GND.n4805 GND.n2734 19.3944
R8973 GND.n4848 GND.n2734 19.3944
R8974 GND.n4848 GND.n2732 19.3944
R8975 GND.n4854 GND.n2732 19.3944
R8976 GND.n4854 GND.n4853 19.3944
R8977 GND.n4853 GND.n2717 19.3944
R8978 GND.n4870 GND.n2717 19.3944
R8979 GND.n4870 GND.n2715 19.3944
R8980 GND.n4875 GND.n2715 19.3944
R8981 GND.n4875 GND.n1900 19.3944
R8982 GND.n5816 GND.n1900 19.3944
R8983 GND.n5816 GND.n5815 19.3944
R8984 GND.n5815 GND.n5814 19.3944
R8985 GND.n5814 GND.n1904 19.3944
R8986 GND.n5810 GND.n1904 19.3944
R8987 GND.n5810 GND.n5809 19.3944
R8988 GND.n5809 GND.n5808 19.3944
R8989 GND.n5808 GND.n1910 19.3944
R8990 GND.n1928 GND.n1910 19.3944
R8991 GND.n5796 GND.n1928 19.3944
R8992 GND.n5796 GND.n5795 19.3944
R8993 GND.n5795 GND.n5794 19.3944
R8994 GND.n5794 GND.n1934 19.3944
R8995 GND.n1955 GND.n1934 19.3944
R8996 GND.n5782 GND.n1955 19.3944
R8997 GND.n5782 GND.n5781 19.3944
R8998 GND.n5781 GND.n5780 19.3944
R8999 GND.n5780 GND.n1961 19.3944
R9000 GND.n1982 GND.n1961 19.3944
R9001 GND.n5768 GND.n1982 19.3944
R9002 GND.n5768 GND.n5767 19.3944
R9003 GND.n5767 GND.n5766 19.3944
R9004 GND.n5766 GND.n1988 19.3944
R9005 GND.n2008 GND.n1988 19.3944
R9006 GND.n5754 GND.n2008 19.3944
R9007 GND.n5754 GND.n5753 19.3944
R9008 GND.n5753 GND.n5752 19.3944
R9009 GND.n5752 GND.n2014 19.3944
R9010 GND.n2035 GND.n2014 19.3944
R9011 GND.n5740 GND.n2035 19.3944
R9012 GND.n5740 GND.n5739 19.3944
R9013 GND.n5739 GND.n5738 19.3944
R9014 GND.n5738 GND.n2041 19.3944
R9015 GND.n2062 GND.n2041 19.3944
R9016 GND.n5726 GND.n2062 19.3944
R9017 GND.n5726 GND.n5725 19.3944
R9018 GND.n5725 GND.n5724 19.3944
R9019 GND.n5724 GND.n2068 19.3944
R9020 GND.n2089 GND.n2068 19.3944
R9021 GND.n5712 GND.n2089 19.3944
R9022 GND.n5712 GND.n5711 19.3944
R9023 GND.n5711 GND.n5710 19.3944
R9024 GND.n5710 GND.n2095 19.3944
R9025 GND.n2116 GND.n2095 19.3944
R9026 GND.n5698 GND.n2116 19.3944
R9027 GND.n5698 GND.n5697 19.3944
R9028 GND.n5697 GND.n5696 19.3944
R9029 GND.n5696 GND.n2122 19.3944
R9030 GND.n2143 GND.n2122 19.3944
R9031 GND.n5684 GND.n2143 19.3944
R9032 GND.n5684 GND.n5683 19.3944
R9033 GND.n5683 GND.n5682 19.3944
R9034 GND.n5682 GND.n2149 19.3944
R9035 GND.n2170 GND.n2149 19.3944
R9036 GND.n5670 GND.n2170 19.3944
R9037 GND.n5670 GND.n5669 19.3944
R9038 GND.n5669 GND.n5668 19.3944
R9039 GND.n5668 GND.n2176 19.3944
R9040 GND.n2196 GND.n2176 19.3944
R9041 GND.n5656 GND.n2196 19.3944
R9042 GND.n5656 GND.n5655 19.3944
R9043 GND.n5655 GND.n5654 19.3944
R9044 GND.n5654 GND.n2202 19.3944
R9045 GND.n2236 GND.n2202 19.3944
R9046 GND.n3130 GND.n3106 19.3944
R9047 GND.n3130 GND.n3129 19.3944
R9048 GND.n4180 GND.n3060 19.3944
R9049 GND.n4180 GND.n4179 19.3944
R9050 GND.n4179 GND.n4178 19.3944
R9051 GND.n4178 GND.n4176 19.3944
R9052 GND.n4176 GND.n4173 19.3944
R9053 GND.n4173 GND.n4172 19.3944
R9054 GND.n4172 GND.n4169 19.3944
R9055 GND.n4169 GND.n4168 19.3944
R9056 GND.n4168 GND.n4165 19.3944
R9057 GND.n4165 GND.n4164 19.3944
R9058 GND.n4164 GND.n4161 19.3944
R9059 GND.n4161 GND.n3071 19.3944
R9060 GND.n3165 GND.n3071 19.3944
R9061 GND.n3165 GND.n3164 19.3944
R9062 GND.n3164 GND.n3077 19.3944
R9063 GND.n3157 GND.n3077 19.3944
R9064 GND.n3157 GND.n3156 19.3944
R9065 GND.n3156 GND.n3087 19.3944
R9066 GND.n3149 GND.n3087 19.3944
R9067 GND.n3149 GND.n3148 19.3944
R9068 GND.n3148 GND.n3097 19.3944
R9069 GND.n3141 GND.n3097 19.3944
R9070 GND.n5434 GND.n2439 19.3944
R9071 GND.n5434 GND.n5433 19.3944
R9072 GND.n5433 GND.n5432 19.3944
R9073 GND.n5432 GND.n2444 19.3944
R9074 GND.n5422 GND.n2444 19.3944
R9075 GND.n5422 GND.n5421 19.3944
R9076 GND.n5421 GND.n5420 19.3944
R9077 GND.n5420 GND.n2465 19.3944
R9078 GND.n5410 GND.n2465 19.3944
R9079 GND.n5410 GND.n5409 19.3944
R9080 GND.n5409 GND.n5408 19.3944
R9081 GND.n5408 GND.n2486 19.3944
R9082 GND.n5398 GND.n2486 19.3944
R9083 GND.n5398 GND.n5397 19.3944
R9084 GND.n5397 GND.n5396 19.3944
R9085 GND.n5396 GND.n2507 19.3944
R9086 GND.n5386 GND.n2507 19.3944
R9087 GND.n5386 GND.n5385 19.3944
R9088 GND.n5385 GND.n5384 19.3944
R9089 GND.n2526 GND.n45 19.3944
R9090 GND.n2542 GND.n45 19.3944
R9091 GND.n8076 GND.n38 19.3944
R9092 GND.n5361 GND.n39 19.3944
R9093 GND.n8073 GND.n47 19.3944
R9094 GND.n8073 GND.n48 19.3944
R9095 GND.n8063 GND.n48 19.3944
R9096 GND.n8063 GND.n8062 19.3944
R9097 GND.n8062 GND.n8061 19.3944
R9098 GND.n8061 GND.n70 19.3944
R9099 GND.n8051 GND.n70 19.3944
R9100 GND.n8051 GND.n8050 19.3944
R9101 GND.n8050 GND.n8049 19.3944
R9102 GND.n8049 GND.n91 19.3944
R9103 GND.n8039 GND.n91 19.3944
R9104 GND.n8039 GND.n8038 19.3944
R9105 GND.n8038 GND.n8037 19.3944
R9106 GND.n8037 GND.n112 19.3944
R9107 GND.n8027 GND.n112 19.3944
R9108 GND.n8027 GND.n8026 19.3944
R9109 GND.n8026 GND.n8025 19.3944
R9110 GND.n8025 GND.n133 19.3944
R9111 GND.n8015 GND.n133 19.3944
R9112 GND.n8015 GND.n8014 19.3944
R9113 GND.n6498 GND.n6497 19.3944
R9114 GND.n6497 GND.n1213 19.3944
R9115 GND.n6491 GND.n1213 19.3944
R9116 GND.n6491 GND.n6490 19.3944
R9117 GND.n6490 GND.n6489 19.3944
R9118 GND.n6489 GND.n1221 19.3944
R9119 GND.n6483 GND.n1221 19.3944
R9120 GND.n6483 GND.n6482 19.3944
R9121 GND.n6482 GND.n6481 19.3944
R9122 GND.n6481 GND.n1229 19.3944
R9123 GND.n6475 GND.n1229 19.3944
R9124 GND.n6475 GND.n6474 19.3944
R9125 GND.n6474 GND.n6473 19.3944
R9126 GND.n6473 GND.n1237 19.3944
R9127 GND.n6467 GND.n1237 19.3944
R9128 GND.n6467 GND.n6466 19.3944
R9129 GND.n6466 GND.n6465 19.3944
R9130 GND.n6465 GND.n1245 19.3944
R9131 GND.n6459 GND.n1245 19.3944
R9132 GND.n6459 GND.n6458 19.3944
R9133 GND.n6458 GND.n6457 19.3944
R9134 GND.n6457 GND.n1253 19.3944
R9135 GND.n6451 GND.n1253 19.3944
R9136 GND.n6451 GND.n6450 19.3944
R9137 GND.n6450 GND.n6449 19.3944
R9138 GND.n6449 GND.n1261 19.3944
R9139 GND.n6443 GND.n1261 19.3944
R9140 GND.n6443 GND.n6442 19.3944
R9141 GND.n6442 GND.n6441 19.3944
R9142 GND.n6441 GND.n1269 19.3944
R9143 GND.n6435 GND.n1269 19.3944
R9144 GND.n6435 GND.n6434 19.3944
R9145 GND.n6434 GND.n6433 19.3944
R9146 GND.n6433 GND.n1277 19.3944
R9147 GND.n6427 GND.n1277 19.3944
R9148 GND.n6427 GND.n6426 19.3944
R9149 GND.n6426 GND.n6425 19.3944
R9150 GND.n6425 GND.n1285 19.3944
R9151 GND.n6419 GND.n1285 19.3944
R9152 GND.n6419 GND.n6418 19.3944
R9153 GND.n6418 GND.n6417 19.3944
R9154 GND.n6417 GND.n1293 19.3944
R9155 GND.n6411 GND.n1293 19.3944
R9156 GND.n6411 GND.n6410 19.3944
R9157 GND.n6410 GND.n6409 19.3944
R9158 GND.n6409 GND.n1301 19.3944
R9159 GND.n6403 GND.n1301 19.3944
R9160 GND.n6403 GND.n6402 19.3944
R9161 GND.n6402 GND.n6401 19.3944
R9162 GND.n6401 GND.n1309 19.3944
R9163 GND.n6395 GND.n1309 19.3944
R9164 GND.n6395 GND.n6394 19.3944
R9165 GND.n6394 GND.n6393 19.3944
R9166 GND.n6393 GND.n1317 19.3944
R9167 GND.n6387 GND.n1317 19.3944
R9168 GND.n6387 GND.n6386 19.3944
R9169 GND.n6386 GND.n6385 19.3944
R9170 GND.n6385 GND.n1325 19.3944
R9171 GND.n3526 GND.n1325 19.3944
R9172 GND.n3530 GND.n3526 19.3944
R9173 GND.n3530 GND.n3514 19.3944
R9174 GND.n3792 GND.n3514 19.3944
R9175 GND.n3792 GND.n3512 19.3944
R9176 GND.n3798 GND.n3512 19.3944
R9177 GND.n3798 GND.n3797 19.3944
R9178 GND.n3797 GND.n3484 19.3944
R9179 GND.n3829 GND.n3484 19.3944
R9180 GND.n3829 GND.n3482 19.3944
R9181 GND.n3835 GND.n3482 19.3944
R9182 GND.n3835 GND.n3834 19.3944
R9183 GND.n3834 GND.n3455 19.3944
R9184 GND.n3866 GND.n3455 19.3944
R9185 GND.n3866 GND.n3453 19.3944
R9186 GND.n3878 GND.n3453 19.3944
R9187 GND.n3878 GND.n3877 19.3944
R9188 GND.n3877 GND.n3876 19.3944
R9189 GND.n3876 GND.n3873 19.3944
R9190 GND.n3873 GND.n3403 19.3944
R9191 GND.n3991 GND.n3403 19.3944
R9192 GND.n3991 GND.n3404 19.3944
R9193 GND.n3940 GND.n3939 19.3944
R9194 GND.n3950 GND.n3949 19.3944
R9195 GND.n3946 GND.n3945 19.3944
R9196 GND.n3942 GND.n3397 19.3944
R9197 GND.n3995 GND.n3372 19.3944
R9198 GND.n4026 GND.n3372 19.3944
R9199 GND.n4026 GND.n3370 19.3944
R9200 GND.n4032 GND.n3370 19.3944
R9201 GND.n4032 GND.n4031 19.3944
R9202 GND.n4031 GND.n3343 19.3944
R9203 GND.n4063 GND.n3343 19.3944
R9204 GND.n4063 GND.n3341 19.3944
R9205 GND.n4069 GND.n3341 19.3944
R9206 GND.n4069 GND.n4068 19.3944
R9207 GND.n4068 GND.n3314 19.3944
R9208 GND.n4100 GND.n3314 19.3944
R9209 GND.n4100 GND.n3312 19.3944
R9210 GND.n4128 GND.n3312 19.3944
R9211 GND.n4128 GND.n4127 19.3944
R9212 GND.n4127 GND.n4126 19.3944
R9213 GND.n4126 GND.n4106 19.3944
R9214 GND.n4122 GND.n4106 19.3944
R9215 GND.n4122 GND.n4121 19.3944
R9216 GND.n4121 GND.n4120 19.3944
R9217 GND.n4120 GND.n4112 19.3944
R9218 GND.n4115 GND.n4112 19.3944
R9219 GND.n4115 GND.n3044 19.3944
R9220 GND.n4186 GND.n3044 19.3944
R9221 GND.n4186 GND.n3042 19.3944
R9222 GND.n4192 GND.n3042 19.3944
R9223 GND.n4192 GND.n4191 19.3944
R9224 GND.n4191 GND.n3022 19.3944
R9225 GND.n4218 GND.n3022 19.3944
R9226 GND.n4218 GND.n3020 19.3944
R9227 GND.n4224 GND.n3020 19.3944
R9228 GND.n4224 GND.n4223 19.3944
R9229 GND.n4223 GND.n2999 19.3944
R9230 GND.n4250 GND.n2999 19.3944
R9231 GND.n4250 GND.n2997 19.3944
R9232 GND.n4256 GND.n2997 19.3944
R9233 GND.n4256 GND.n4255 19.3944
R9234 GND.n4255 GND.n2976 19.3944
R9235 GND.n4282 GND.n2976 19.3944
R9236 GND.n4282 GND.n2974 19.3944
R9237 GND.n4288 GND.n2974 19.3944
R9238 GND.n4288 GND.n4287 19.3944
R9239 GND.n4287 GND.n2953 19.3944
R9240 GND.n4314 GND.n2953 19.3944
R9241 GND.n4314 GND.n2951 19.3944
R9242 GND.n4320 GND.n2951 19.3944
R9243 GND.n4320 GND.n4319 19.3944
R9244 GND.n4319 GND.n2930 19.3944
R9245 GND.n4346 GND.n2930 19.3944
R9246 GND.n4346 GND.n2928 19.3944
R9247 GND.n4352 GND.n2928 19.3944
R9248 GND.n4352 GND.n4351 19.3944
R9249 GND.n4351 GND.n2907 19.3944
R9250 GND.n4378 GND.n2907 19.3944
R9251 GND.n4378 GND.n2905 19.3944
R9252 GND.n4384 GND.n2905 19.3944
R9253 GND.n4384 GND.n4383 19.3944
R9254 GND.n4383 GND.n2884 19.3944
R9255 GND.n4410 GND.n2884 19.3944
R9256 GND.n4410 GND.n2882 19.3944
R9257 GND.n4416 GND.n2882 19.3944
R9258 GND.n4416 GND.n4415 19.3944
R9259 GND.n4415 GND.n2861 19.3944
R9260 GND.n4442 GND.n2861 19.3944
R9261 GND.n4442 GND.n2859 19.3944
R9262 GND.n4448 GND.n2859 19.3944
R9263 GND.n4448 GND.n4447 19.3944
R9264 GND.n4447 GND.n2838 19.3944
R9265 GND.n4474 GND.n2838 19.3944
R9266 GND.n4474 GND.n2836 19.3944
R9267 GND.n4480 GND.n2836 19.3944
R9268 GND.n4480 GND.n4479 19.3944
R9269 GND.n4479 GND.n2815 19.3944
R9270 GND.n4506 GND.n2815 19.3944
R9271 GND.n4506 GND.n2813 19.3944
R9272 GND.n4512 GND.n2813 19.3944
R9273 GND.n4512 GND.n4511 19.3944
R9274 GND.n4511 GND.n2792 19.3944
R9275 GND.n4541 GND.n2792 19.3944
R9276 GND.n4541 GND.n2790 19.3944
R9277 GND.n4563 GND.n2790 19.3944
R9278 GND.n4563 GND.n4562 19.3944
R9279 GND.n4562 GND.n4561 19.3944
R9280 GND.n4561 GND.n4547 19.3944
R9281 GND.n4557 GND.n4547 19.3944
R9282 GND.n4557 GND.n4556 19.3944
R9283 GND.n4556 GND.n4555 19.3944
R9284 GND.n4555 GND.n1674 19.3944
R9285 GND.n6127 GND.n1674 19.3944
R9286 GND.n6127 GND.n6126 19.3944
R9287 GND.n6126 GND.n6125 19.3944
R9288 GND.n6125 GND.n1678 19.3944
R9289 GND.n1712 GND.n1678 19.3944
R9290 GND.n1712 GND.n1709 19.3944
R9291 GND.n6107 GND.n1709 19.3944
R9292 GND.n6107 GND.n6106 19.3944
R9293 GND.n6106 GND.n6105 19.3944
R9294 GND.n6105 GND.n1718 19.3944
R9295 GND.n1756 GND.n1718 19.3944
R9296 GND.n1756 GND.n1753 19.3944
R9297 GND.n6086 GND.n1753 19.3944
R9298 GND.n6086 GND.n6085 19.3944
R9299 GND.n6085 GND.n6084 19.3944
R9300 GND.n6084 GND.n1762 19.3944
R9301 GND.n6072 GND.n1762 19.3944
R9302 GND.n6072 GND.n6071 19.3944
R9303 GND.n6071 GND.n6070 19.3944
R9304 GND.n6070 GND.n1780 19.3944
R9305 GND.n6058 GND.n1780 19.3944
R9306 GND.n6058 GND.n6057 19.3944
R9307 GND.n6057 GND.n6056 19.3944
R9308 GND.n6056 GND.n1798 19.3944
R9309 GND.n6044 GND.n1798 19.3944
R9310 GND.n6044 GND.n6043 19.3944
R9311 GND.n6043 GND.n6042 19.3944
R9312 GND.n6042 GND.n1815 19.3944
R9313 GND.n6030 GND.n1815 19.3944
R9314 GND.n6030 GND.n6029 19.3944
R9315 GND.n6029 GND.n6028 19.3944
R9316 GND.n6028 GND.n1832 19.3944
R9317 GND.n6016 GND.n1832 19.3944
R9318 GND.n6016 GND.n6015 19.3944
R9319 GND.n6015 GND.n6014 19.3944
R9320 GND.n6014 GND.n1850 19.3944
R9321 GND.n5803 GND.n1850 19.3944
R9322 GND.n5803 GND.n5802 19.3944
R9323 GND.n5802 GND.n5801 19.3944
R9324 GND.n5801 GND.n1920 19.3944
R9325 GND.n1941 GND.n1920 19.3944
R9326 GND.n5789 GND.n1941 19.3944
R9327 GND.n5789 GND.n5788 19.3944
R9328 GND.n5788 GND.n5787 19.3944
R9329 GND.n5787 GND.n1947 19.3944
R9330 GND.n1968 GND.n1947 19.3944
R9331 GND.n5775 GND.n1968 19.3944
R9332 GND.n5775 GND.n5774 19.3944
R9333 GND.n5774 GND.n5773 19.3944
R9334 GND.n5773 GND.n1974 19.3944
R9335 GND.n1995 GND.n1974 19.3944
R9336 GND.n5761 GND.n1995 19.3944
R9337 GND.n5761 GND.n5760 19.3944
R9338 GND.n5760 GND.n5759 19.3944
R9339 GND.n5759 GND.n2001 19.3944
R9340 GND.n2021 GND.n2001 19.3944
R9341 GND.n5747 GND.n2021 19.3944
R9342 GND.n5747 GND.n5746 19.3944
R9343 GND.n5746 GND.n5745 19.3944
R9344 GND.n5745 GND.n2027 19.3944
R9345 GND.n2048 GND.n2027 19.3944
R9346 GND.n5733 GND.n2048 19.3944
R9347 GND.n5733 GND.n5732 19.3944
R9348 GND.n5732 GND.n5731 19.3944
R9349 GND.n5731 GND.n2054 19.3944
R9350 GND.n2075 GND.n2054 19.3944
R9351 GND.n5719 GND.n2075 19.3944
R9352 GND.n5719 GND.n5718 19.3944
R9353 GND.n5718 GND.n5717 19.3944
R9354 GND.n5717 GND.n2081 19.3944
R9355 GND.n2102 GND.n2081 19.3944
R9356 GND.n5705 GND.n2102 19.3944
R9357 GND.n5705 GND.n5704 19.3944
R9358 GND.n5704 GND.n5703 19.3944
R9359 GND.n5703 GND.n2108 19.3944
R9360 GND.n2129 GND.n2108 19.3944
R9361 GND.n5691 GND.n2129 19.3944
R9362 GND.n5691 GND.n5690 19.3944
R9363 GND.n5690 GND.n5689 19.3944
R9364 GND.n5689 GND.n2135 19.3944
R9365 GND.n2156 GND.n2135 19.3944
R9366 GND.n5677 GND.n2156 19.3944
R9367 GND.n5677 GND.n5676 19.3944
R9368 GND.n5676 GND.n5675 19.3944
R9369 GND.n5675 GND.n2162 19.3944
R9370 GND.n2182 GND.n2162 19.3944
R9371 GND.n5663 GND.n2182 19.3944
R9372 GND.n5663 GND.n5662 19.3944
R9373 GND.n5662 GND.n5661 19.3944
R9374 GND.n5661 GND.n2188 19.3944
R9375 GND.n2209 GND.n2188 19.3944
R9376 GND.n5649 GND.n2209 19.3944
R9377 GND.n5649 GND.n5648 19.3944
R9378 GND.n5648 GND.n5647 19.3944
R9379 GND.n5647 GND.n2215 19.3944
R9380 GND.n2592 GND.n2215 19.3944
R9381 GND.n2592 GND.n2589 19.3944
R9382 GND.n2596 GND.n2589 19.3944
R9383 GND.n2596 GND.n2586 19.3944
R9384 GND.n2600 GND.n2586 19.3944
R9385 GND.n2600 GND.n2584 19.3944
R9386 GND.n2604 GND.n2584 19.3944
R9387 GND.n2604 GND.n2582 19.3944
R9388 GND.n2608 GND.n2582 19.3944
R9389 GND.n2608 GND.n2580 19.3944
R9390 GND.n2655 GND.n2580 19.3944
R9391 GND.n2655 GND.n2654 19.3944
R9392 GND.n2654 GND.n2653 19.3944
R9393 GND.n2653 GND.n2614 19.3944
R9394 GND.n2649 GND.n2614 19.3944
R9395 GND.n2649 GND.n2648 19.3944
R9396 GND.n2648 GND.n2647 19.3944
R9397 GND.n2647 GND.n2620 19.3944
R9398 GND.n2643 GND.n2620 19.3944
R9399 GND.n2643 GND.n2642 19.3944
R9400 GND.n2642 GND.n2641 19.3944
R9401 GND.n2641 GND.n2626 19.3944
R9402 GND.n2637 GND.n2626 19.3944
R9403 GND.n2637 GND.n2636 19.3944
R9404 GND.n2634 GND.n2631 19.3944
R9405 GND.n5370 GND.n2548 19.3944
R9406 GND.n5368 GND.n5367 19.3944
R9407 GND.n5145 GND.n2551 19.3944
R9408 GND.n5200 GND.n5147 19.3944
R9409 GND.n5200 GND.n5199 19.3944
R9410 GND.n5199 GND.n5198 19.3944
R9411 GND.n5198 GND.n5151 19.3944
R9412 GND.n5194 GND.n5151 19.3944
R9413 GND.n5194 GND.n5193 19.3944
R9414 GND.n5193 GND.n5192 19.3944
R9415 GND.n5192 GND.n5157 19.3944
R9416 GND.n5188 GND.n5157 19.3944
R9417 GND.n5188 GND.n5187 19.3944
R9418 GND.n5187 GND.n5186 19.3944
R9419 GND.n5186 GND.n5163 19.3944
R9420 GND.n5182 GND.n5163 19.3944
R9421 GND.n5182 GND.n5181 19.3944
R9422 GND.n5181 GND.n5180 19.3944
R9423 GND.n5180 GND.n5169 19.3944
R9424 GND.n5176 GND.n5169 19.3944
R9425 GND.n5176 GND.n5175 19.3944
R9426 GND.n5175 GND.n294 19.3944
R9427 GND.n7872 GND.n294 19.3944
R9428 GND.n7872 GND.n7871 19.3944
R9429 GND.n7871 GND.n7870 19.3944
R9430 GND.n7870 GND.n298 19.3944
R9431 GND.n7864 GND.n298 19.3944
R9432 GND.n7864 GND.n7863 19.3944
R9433 GND.n7863 GND.n7862 19.3944
R9434 GND.n7862 GND.n306 19.3944
R9435 GND.n7856 GND.n306 19.3944
R9436 GND.n7856 GND.n7855 19.3944
R9437 GND.n7855 GND.n7854 19.3944
R9438 GND.n7854 GND.n314 19.3944
R9439 GND.n7848 GND.n314 19.3944
R9440 GND.n7848 GND.n7847 19.3944
R9441 GND.n7847 GND.n7846 19.3944
R9442 GND.n7846 GND.n322 19.3944
R9443 GND.n7840 GND.n322 19.3944
R9444 GND.n7840 GND.n7839 19.3944
R9445 GND.n7839 GND.n7838 19.3944
R9446 GND.n7838 GND.n330 19.3944
R9447 GND.n7832 GND.n330 19.3944
R9448 GND.n7832 GND.n7831 19.3944
R9449 GND.n7831 GND.n7830 19.3944
R9450 GND.n7830 GND.n338 19.3944
R9451 GND.n7824 GND.n338 19.3944
R9452 GND.n7824 GND.n7823 19.3944
R9453 GND.n7823 GND.n7822 19.3944
R9454 GND.n7822 GND.n346 19.3944
R9455 GND.n7816 GND.n346 19.3944
R9456 GND.n7816 GND.n7815 19.3944
R9457 GND.n7815 GND.n7814 19.3944
R9458 GND.n7814 GND.n354 19.3944
R9459 GND.n7808 GND.n354 19.3944
R9460 GND.n7808 GND.n7807 19.3944
R9461 GND.n7807 GND.n7806 19.3944
R9462 GND.n7806 GND.n362 19.3944
R9463 GND.n7800 GND.n362 19.3944
R9464 GND.n7800 GND.n7799 19.3944
R9465 GND.n7799 GND.n7798 19.3944
R9466 GND.n7798 GND.n370 19.3944
R9467 GND.n7792 GND.n370 19.3944
R9468 GND.n7792 GND.n7791 19.3944
R9469 GND.n7791 GND.n7790 19.3944
R9470 GND.n7790 GND.n378 19.3944
R9471 GND.n7784 GND.n378 19.3944
R9472 GND.n7784 GND.n7783 19.3944
R9473 GND.n7783 GND.n7782 19.3944
R9474 GND.n7782 GND.n386 19.3944
R9475 GND.n7776 GND.n386 19.3944
R9476 GND.n7776 GND.n7775 19.3944
R9477 GND.n7775 GND.n7774 19.3944
R9478 GND.n7774 GND.n394 19.3944
R9479 GND.n7768 GND.n394 19.3944
R9480 GND.n7768 GND.n7767 19.3944
R9481 GND.n7767 GND.n7766 19.3944
R9482 GND.n7766 GND.n402 19.3944
R9483 GND.n7760 GND.n402 19.3944
R9484 GND.n7760 GND.n7759 19.3944
R9485 GND.n7759 GND.n7758 19.3944
R9486 GND.n7758 GND.n410 19.3944
R9487 GND.n7752 GND.n410 19.3944
R9488 GND.n3579 GND.n3576 19.3944
R9489 GND.n3579 GND.n3575 19.3944
R9490 GND.n3583 GND.n3575 19.3944
R9491 GND.n3586 GND.n3583 19.3944
R9492 GND.n3589 GND.n3586 19.3944
R9493 GND.n3589 GND.n3573 19.3944
R9494 GND.n3593 GND.n3573 19.3944
R9495 GND.n3596 GND.n3593 19.3944
R9496 GND.n3599 GND.n3596 19.3944
R9497 GND.n3599 GND.n3571 19.3944
R9498 GND.n3603 GND.n3571 19.3944
R9499 GND.n3606 GND.n3603 19.3944
R9500 GND.n3609 GND.n3606 19.3944
R9501 GND.n3609 GND.n3569 19.3944
R9502 GND.n3613 GND.n3569 19.3944
R9503 GND.n3621 GND.n3567 19.3944
R9504 GND.n3625 GND.n3567 19.3944
R9505 GND.n3628 GND.n3625 19.3944
R9506 GND.n3631 GND.n3628 19.3944
R9507 GND.n3631 GND.n3565 19.3944
R9508 GND.n3635 GND.n3565 19.3944
R9509 GND.n3638 GND.n3635 19.3944
R9510 GND.n3641 GND.n3638 19.3944
R9511 GND.n3641 GND.n3563 19.3944
R9512 GND.n3645 GND.n3563 19.3944
R9513 GND.n3648 GND.n3645 19.3944
R9514 GND.n3651 GND.n3648 19.3944
R9515 GND.n3651 GND.n3561 19.3944
R9516 GND.n3655 GND.n3561 19.3944
R9517 GND.n3658 GND.n3655 19.3944
R9518 GND.n3661 GND.n3658 19.3944
R9519 GND.n3661 GND.n3559 19.3944
R9520 GND.n3673 GND.n3670 19.3944
R9521 GND.n3673 GND.n3557 19.3944
R9522 GND.n3677 GND.n3557 19.3944
R9523 GND.n3680 GND.n3677 19.3944
R9524 GND.n3683 GND.n3680 19.3944
R9525 GND.n3683 GND.n3555 19.3944
R9526 GND.n3687 GND.n3555 19.3944
R9527 GND.n3690 GND.n3687 19.3944
R9528 GND.n3693 GND.n3690 19.3944
R9529 GND.n3693 GND.n3553 19.3944
R9530 GND.n3697 GND.n3553 19.3944
R9531 GND.n3700 GND.n3697 19.3944
R9532 GND.n3703 GND.n3700 19.3944
R9533 GND.n3703 GND.n3551 19.3944
R9534 GND.n3707 GND.n3551 19.3944
R9535 GND.n3710 GND.n3707 19.3944
R9536 GND.n3716 GND.n3710 19.3944
R9537 GND.n3720 GND.n3549 19.3944
R9538 GND.n3723 GND.n3720 19.3944
R9539 GND.n3726 GND.n3723 19.3944
R9540 GND.n3726 GND.n3547 19.3944
R9541 GND.n3730 GND.n3547 19.3944
R9542 GND.n3733 GND.n3730 19.3944
R9543 GND.n3736 GND.n3733 19.3944
R9544 GND.n3736 GND.n3545 19.3944
R9545 GND.n3740 GND.n3545 19.3944
R9546 GND.n3743 GND.n3740 19.3944
R9547 GND.n3746 GND.n3743 19.3944
R9548 GND.n3746 GND.n3543 19.3944
R9549 GND.n3750 GND.n3543 19.3944
R9550 GND.n3753 GND.n3750 19.3944
R9551 GND.n3756 GND.n3753 19.3944
R9552 GND.n3756 GND.n3540 19.3944
R9553 GND.n3760 GND.n3540 19.3944
R9554 GND.n3781 GND.n3522 19.3944
R9555 GND.n3787 GND.n3522 19.3944
R9556 GND.n3787 GND.n3786 19.3944
R9557 GND.n3786 GND.n3495 19.3944
R9558 GND.n3818 GND.n3495 19.3944
R9559 GND.n3818 GND.n3493 19.3944
R9560 GND.n3824 GND.n3493 19.3944
R9561 GND.n3824 GND.n3823 19.3944
R9562 GND.n3823 GND.n3466 19.3944
R9563 GND.n3855 GND.n3466 19.3944
R9564 GND.n3855 GND.n3464 19.3944
R9565 GND.n3861 GND.n3464 19.3944
R9566 GND.n3861 GND.n3860 19.3944
R9567 GND.n3860 GND.n3437 19.3944
R9568 GND.n3895 GND.n3437 19.3944
R9569 GND.n3895 GND.n3435 19.3944
R9570 GND.n3900 GND.n3435 19.3944
R9571 GND.n3900 GND.n3414 19.3944
R9572 GND.n3986 GND.n3414 19.3944
R9573 GND.n3984 GND.n3983 19.3944
R9574 GND.n3983 GND.n3415 19.3944
R9575 GND.n3961 GND.n3932 19.3944
R9576 GND.n3966 GND.n3963 19.3944
R9577 GND.n3964 GND.n3383 19.3944
R9578 GND.n4015 GND.n3383 19.3944
R9579 GND.n4015 GND.n3381 19.3944
R9580 GND.n4021 GND.n3381 19.3944
R9581 GND.n4021 GND.n4020 19.3944
R9582 GND.n4020 GND.n3354 19.3944
R9583 GND.n4052 GND.n3354 19.3944
R9584 GND.n4052 GND.n3352 19.3944
R9585 GND.n4058 GND.n3352 19.3944
R9586 GND.n4058 GND.n4057 19.3944
R9587 GND.n4057 GND.n3324 19.3944
R9588 GND.n4089 GND.n3324 19.3944
R9589 GND.n4089 GND.n3322 19.3944
R9590 GND.n4095 GND.n3322 19.3944
R9591 GND.n4095 GND.n4094 19.3944
R9592 GND.n4094 GND.n3297 19.3944
R9593 GND.n4144 GND.n3297 19.3944
R9594 GND.n4144 GND.n3295 19.3944
R9595 GND.n4149 GND.n3295 19.3944
R9596 GND.n4149 GND.n4148 19.3944
R9597 GND.n6627 GND.n1088 19.3944
R9598 GND.n6621 GND.n1088 19.3944
R9599 GND.n6621 GND.n6620 19.3944
R9600 GND.n6620 GND.n6619 19.3944
R9601 GND.n6619 GND.n1095 19.3944
R9602 GND.n6613 GND.n1095 19.3944
R9603 GND.n6613 GND.n6612 19.3944
R9604 GND.n6612 GND.n6611 19.3944
R9605 GND.n6611 GND.n1103 19.3944
R9606 GND.n6605 GND.n1103 19.3944
R9607 GND.n6605 GND.n6604 19.3944
R9608 GND.n6604 GND.n6603 19.3944
R9609 GND.n6603 GND.n1111 19.3944
R9610 GND.n6597 GND.n1111 19.3944
R9611 GND.n6597 GND.n6596 19.3944
R9612 GND.n6596 GND.n6595 19.3944
R9613 GND.n6595 GND.n1119 19.3944
R9614 GND.n6589 GND.n1119 19.3944
R9615 GND.n6589 GND.n6588 19.3944
R9616 GND.n6588 GND.n6587 19.3944
R9617 GND.n6587 GND.n1127 19.3944
R9618 GND.n6581 GND.n1127 19.3944
R9619 GND.n6581 GND.n6580 19.3944
R9620 GND.n6580 GND.n6579 19.3944
R9621 GND.n6579 GND.n1135 19.3944
R9622 GND.n6573 GND.n1135 19.3944
R9623 GND.n6573 GND.n6572 19.3944
R9624 GND.n6572 GND.n6571 19.3944
R9625 GND.n6571 GND.n1143 19.3944
R9626 GND.n6565 GND.n1143 19.3944
R9627 GND.n6565 GND.n6564 19.3944
R9628 GND.n6564 GND.n6563 19.3944
R9629 GND.n6563 GND.n1151 19.3944
R9630 GND.n6557 GND.n1151 19.3944
R9631 GND.n6557 GND.n6556 19.3944
R9632 GND.n6556 GND.n6555 19.3944
R9633 GND.n6555 GND.n1159 19.3944
R9634 GND.n6549 GND.n1159 19.3944
R9635 GND.n6549 GND.n6548 19.3944
R9636 GND.n6548 GND.n6547 19.3944
R9637 GND.n6547 GND.n1167 19.3944
R9638 GND.n6541 GND.n1167 19.3944
R9639 GND.n6541 GND.n6540 19.3944
R9640 GND.n6540 GND.n6539 19.3944
R9641 GND.n6539 GND.n1175 19.3944
R9642 GND.n6533 GND.n1175 19.3944
R9643 GND.n6533 GND.n6532 19.3944
R9644 GND.n6532 GND.n6531 19.3944
R9645 GND.n6531 GND.n1183 19.3944
R9646 GND.n6525 GND.n1183 19.3944
R9647 GND.n6525 GND.n6524 19.3944
R9648 GND.n6524 GND.n6523 19.3944
R9649 GND.n6523 GND.n1191 19.3944
R9650 GND.n6517 GND.n1191 19.3944
R9651 GND.n6517 GND.n6516 19.3944
R9652 GND.n6516 GND.n6515 19.3944
R9653 GND.n6515 GND.n1199 19.3944
R9654 GND.n6509 GND.n1199 19.3944
R9655 GND.n6509 GND.n6508 19.3944
R9656 GND.n6508 GND.n6507 19.3944
R9657 GND.n6507 GND.n1207 19.3944
R9658 GND.n6501 GND.n1207 19.3944
R9659 GND.n6379 GND.n6378 19.3944
R9660 GND.n6378 GND.n1377 19.3944
R9661 GND.n6374 GND.n1377 19.3944
R9662 GND.n6374 GND.n6373 19.3944
R9663 GND.n6373 GND.n6372 19.3944
R9664 GND.n6372 GND.n1383 19.3944
R9665 GND.n6368 GND.n1383 19.3944
R9666 GND.n6368 GND.n6367 19.3944
R9667 GND.n6367 GND.n6366 19.3944
R9668 GND.n6366 GND.n1389 19.3944
R9669 GND.n6362 GND.n1389 19.3944
R9670 GND.n6362 GND.n6361 19.3944
R9671 GND.n6361 GND.n6360 19.3944
R9672 GND.n6360 GND.n1395 19.3944
R9673 GND.n6356 GND.n1395 19.3944
R9674 GND.n6348 GND.n6347 19.3944
R9675 GND.n6347 GND.n6346 19.3944
R9676 GND.n6346 GND.n1403 19.3944
R9677 GND.n6342 GND.n1403 19.3944
R9678 GND.n6342 GND.n6341 19.3944
R9679 GND.n6341 GND.n6340 19.3944
R9680 GND.n6340 GND.n1408 19.3944
R9681 GND.n6336 GND.n1408 19.3944
R9682 GND.n6336 GND.n6335 19.3944
R9683 GND.n6335 GND.n6334 19.3944
R9684 GND.n6334 GND.n1413 19.3944
R9685 GND.n6330 GND.n1413 19.3944
R9686 GND.n6330 GND.n6329 19.3944
R9687 GND.n6329 GND.n6328 19.3944
R9688 GND.n6328 GND.n1418 19.3944
R9689 GND.n6324 GND.n1418 19.3944
R9690 GND.n6324 GND.n6323 19.3944
R9691 GND.n6323 GND.n6322 19.3944
R9692 GND.n6322 GND.n1423 19.3944
R9693 GND.n6318 GND.n1423 19.3944
R9694 GND.n6318 GND.n6317 19.3944
R9695 GND.n6317 GND.n6316 19.3944
R9696 GND.n6316 GND.n1428 19.3944
R9697 GND.n6311 GND.n1428 19.3944
R9698 GND.n6311 GND.n6310 19.3944
R9699 GND.n6310 GND.n6309 19.3944
R9700 GND.n6309 GND.n1433 19.3944
R9701 GND.n6305 GND.n1433 19.3944
R9702 GND.n6305 GND.n6304 19.3944
R9703 GND.n6304 GND.n6303 19.3944
R9704 GND.n6303 GND.n1438 19.3944
R9705 GND.n6299 GND.n1438 19.3944
R9706 GND.n6299 GND.n6298 19.3944
R9707 GND.n6298 GND.n6297 19.3944
R9708 GND.n6297 GND.n1443 19.3944
R9709 GND.n6293 GND.n1443 19.3944
R9710 GND.n6293 GND.n6292 19.3944
R9711 GND.n6292 GND.n6291 19.3944
R9712 GND.n6291 GND.n1448 19.3944
R9713 GND.n6287 GND.n1448 19.3944
R9714 GND.n6287 GND.n6286 19.3944
R9715 GND.n6286 GND.n6285 19.3944
R9716 GND.n6285 GND.n1453 19.3944
R9717 GND.n6281 GND.n1453 19.3944
R9718 GND.n6281 GND.n6280 19.3944
R9719 GND.n6280 GND.n6279 19.3944
R9720 GND.n6279 GND.n1458 19.3944
R9721 GND.n3124 GND.n1462 18.0369
R9722 GND.n5288 GND.n5234 18.0369
R9723 GND.n5040 GND.n5039 18.0369
R9724 GND.n6356 GND.n6355 18.0369
R9725 GND.n4183 GND.n3046 17.2554
R9726 GND.n5643 GND.n2219 17.2554
R9727 GND.t84 GND.n3309 16.9579
R9728 GND.n5424 GND.t53 16.9579
R9729 GND.n3286 GND.n3173 16.8732
R9730 GND.n5448 GND.n2398 16.8732
R9731 GND.n7883 GND.n7882 16.8732
R9732 GND.n3761 GND.n3760 16.8732
R9733 GND.n5594 GND.n2259 16.2914
R9734 GND.n3140 GND.n3106 16.2914
R9735 GND.n6248 GND.n6247 16.0975
R9736 GND.n5557 GND.n5556 16.0975
R9737 GND.n7948 GND.n213 16.0975
R9738 GND.n7983 GND.n7982 16.0975
R9739 GND.n3618 GND.n3613 16.0975
R9740 GND.n3670 GND.n3667 16.0975
R9741 GND.n1642 GND.n1619 16.0672
R9742 GND.n1632 GND.n1621 16.0672
R9743 GND.n5844 GND.n5843 16.0672
R9744 GND.n5850 GND.n5837 16.0672
R9745 GND.t18 GND.n3988 15.7679
R9746 GND.n8071 GND.t10 15.7679
R9747 GND.n5842 GND.n5841 15.4533
R9748 GND.n4195 GND.n3037 14.8754
R9749 GND.n4195 GND.n4194 14.8754
R9750 GND.n4194 GND.n3039 14.8754
R9751 GND.n3039 GND.n3030 14.8754
R9752 GND.n4205 GND.n3030 14.8754
R9753 GND.n4205 GND.n3031 14.8754
R9754 GND.n3031 GND.n3024 14.8754
R9755 GND.n4216 GND.n3024 14.8754
R9756 GND.n4216 GND.n4215 14.8754
R9757 GND.n4215 GND.n3015 14.8754
R9758 GND.n4227 GND.n3015 14.8754
R9759 GND.n4227 GND.n4226 14.8754
R9760 GND.n4226 GND.n3017 14.8754
R9761 GND.n3017 GND.n3007 14.8754
R9762 GND.n4237 GND.n3007 14.8754
R9763 GND.n3008 GND.n3001 14.8754
R9764 GND.n4248 GND.n3001 14.8754
R9765 GND.n4248 GND.n4247 14.8754
R9766 GND.n4247 GND.n2992 14.8754
R9767 GND.n4259 GND.n2992 14.8754
R9768 GND.n4259 GND.n4258 14.8754
R9769 GND.n4258 GND.n2994 14.8754
R9770 GND.n2994 GND.n2984 14.8754
R9771 GND.n4269 GND.n2984 14.8754
R9772 GND.n4269 GND.n2985 14.8754
R9773 GND.n2985 GND.n2978 14.8754
R9774 GND.n4280 GND.n2978 14.8754
R9775 GND.n4280 GND.n4279 14.8754
R9776 GND.n4279 GND.n2969 14.8754
R9777 GND.n4291 GND.n2969 14.8754
R9778 GND.n4291 GND.n4290 14.8754
R9779 GND.n4290 GND.n2971 14.8754
R9780 GND.n2971 GND.n2961 14.8754
R9781 GND.n4301 GND.n2961 14.8754
R9782 GND.n4301 GND.n2962 14.8754
R9783 GND.n2962 GND.n2955 14.8754
R9784 GND.n4312 GND.n2955 14.8754
R9785 GND.n4312 GND.n4311 14.8754
R9786 GND.n4311 GND.n2946 14.8754
R9787 GND.n4323 GND.n2946 14.8754
R9788 GND.n4323 GND.n4322 14.8754
R9789 GND.n4322 GND.n2948 14.8754
R9790 GND.n2948 GND.n2937 14.8754
R9791 GND.n4333 GND.n2937 14.8754
R9792 GND.n4333 GND.n2938 14.8754
R9793 GND.n2940 GND.n2938 14.8754
R9794 GND.n4344 GND.n4343 14.8754
R9795 GND.n4343 GND.n2923 14.8754
R9796 GND.n4355 GND.n2923 14.8754
R9797 GND.n4355 GND.n4354 14.8754
R9798 GND.n4354 GND.n2925 14.8754
R9799 GND.n2925 GND.n2915 14.8754
R9800 GND.n4365 GND.n2915 14.8754
R9801 GND.n4365 GND.n2916 14.8754
R9802 GND.n2916 GND.n2909 14.8754
R9803 GND.n4376 GND.n2909 14.8754
R9804 GND.n4376 GND.n4375 14.8754
R9805 GND.n4375 GND.n2900 14.8754
R9806 GND.n4387 GND.n2900 14.8754
R9807 GND.n4387 GND.n4386 14.8754
R9808 GND.n4386 GND.n2902 14.8754
R9809 GND.n2902 GND.n2892 14.8754
R9810 GND.n4397 GND.n2892 14.8754
R9811 GND.n4397 GND.n2893 14.8754
R9812 GND.n2893 GND.n2886 14.8754
R9813 GND.n4408 GND.n2886 14.8754
R9814 GND.n4408 GND.n4407 14.8754
R9815 GND.n4407 GND.n2877 14.8754
R9816 GND.n4419 GND.n2877 14.8754
R9817 GND.n4419 GND.n4418 14.8754
R9818 GND.n4418 GND.n2879 14.8754
R9819 GND.n2879 GND.n2869 14.8754
R9820 GND.n4429 GND.n2869 14.8754
R9821 GND.n4429 GND.n2870 14.8754
R9822 GND.n2870 GND.n2863 14.8754
R9823 GND.n4440 GND.n2863 14.8754
R9824 GND.n4439 GND.n2854 14.8754
R9825 GND.n4451 GND.n2854 14.8754
R9826 GND.n4451 GND.n4450 14.8754
R9827 GND.n4450 GND.n2856 14.8754
R9828 GND.n2856 GND.n2846 14.8754
R9829 GND.n4461 GND.n2846 14.8754
R9830 GND.n4461 GND.n2847 14.8754
R9831 GND.n2847 GND.n2840 14.8754
R9832 GND.n4472 GND.n2840 14.8754
R9833 GND.n4472 GND.n4471 14.8754
R9834 GND.n4471 GND.n2831 14.8754
R9835 GND.n4483 GND.n2831 14.8754
R9836 GND.n4483 GND.n4482 14.8754
R9837 GND.n4482 GND.n2833 14.8754
R9838 GND.n2833 GND.n2823 14.8754
R9839 GND.n4493 GND.n2823 14.8754
R9840 GND.n4493 GND.n2824 14.8754
R9841 GND.n2824 GND.n2817 14.8754
R9842 GND.n4504 GND.n2817 14.8754
R9843 GND.n4504 GND.n4503 14.8754
R9844 GND.n4503 GND.n2808 14.8754
R9845 GND.n4515 GND.n2808 14.8754
R9846 GND.n4515 GND.n4514 14.8754
R9847 GND.n4514 GND.n2810 14.8754
R9848 GND.n2810 GND.n2800 14.8754
R9849 GND.n4525 GND.n2800 14.8754
R9850 GND.n4525 GND.n2801 14.8754
R9851 GND.n2801 GND.n2794 14.8754
R9852 GND.n4539 GND.n2794 14.8754
R9853 GND.n4539 GND.n4538 14.8754
R9854 GND.n4566 GND.n2785 14.8754
R9855 GND.n4566 GND.n4565 14.8754
R9856 GND.n4565 GND.n2787 14.8754
R9857 GND.n2787 GND.n2777 14.8754
R9858 GND.n4577 GND.n2777 14.8754
R9859 GND.n4577 GND.n2778 14.8754
R9860 GND.n2778 GND.n1578 14.8754
R9861 GND.n4653 GND.n1613 14.8754
R9862 GND.n6143 GND.n1652 14.8754
R9863 GND.n6137 GND.n1661 14.8754
R9864 GND.n6129 GND.n1671 14.8754
R9865 GND.n6116 GND.n1696 14.8754
R9866 GND.n6109 GND.t40 14.8754
R9867 GND.n6109 GND.n1705 14.8754
R9868 GND.n6103 GND.n1720 14.8754
R9869 GND.n6095 GND.n1731 14.8754
R9870 GND.n6089 GND.n6088 14.8754
R9871 GND.n6082 GND.n1764 14.8754
R9872 GND.n4746 GND.n1772 14.8754
R9873 GND.n4809 GND.n4808 14.8754
R9874 GND.n4817 GND.n1790 14.8754
R9875 GND.n4842 GND.n4841 14.8754
R9876 GND.n4856 GND.n2729 14.8754
R9877 GND.n2729 GND.n1807 14.8754
R9878 GND.n2712 GND.n1819 14.8754
R9879 GND.n4879 GND.n1896 14.8754
R9880 GND.n5826 GND.n1836 14.8754
R9881 GND.n6018 GND.n1844 14.8754
R9882 GND.n6012 GND.n1852 14.8754
R9883 GND.n5806 GND.n1912 14.8754
R9884 GND.n5806 GND.n5805 14.8754
R9885 GND.n5805 GND.n1914 14.8754
R9886 GND.n1922 GND.n1914 14.8754
R9887 GND.n1923 GND.n1922 14.8754
R9888 GND.n5799 GND.n1923 14.8754
R9889 GND.n5798 GND.n1925 14.8754
R9890 GND.n4903 GND.n1925 14.8754
R9891 GND.n4903 GND.n1936 14.8754
R9892 GND.n5792 GND.n1936 14.8754
R9893 GND.n5792 GND.n5791 14.8754
R9894 GND.n5791 GND.n1938 14.8754
R9895 GND.n1949 GND.n1938 14.8754
R9896 GND.n1950 GND.n1949 14.8754
R9897 GND.n5785 GND.n1950 14.8754
R9898 GND.n5785 GND.n5784 14.8754
R9899 GND.n5784 GND.n1952 14.8754
R9900 GND.n4914 GND.n1952 14.8754
R9901 GND.n4914 GND.n1963 14.8754
R9902 GND.n5778 GND.n1963 14.8754
R9903 GND.n5778 GND.n5777 14.8754
R9904 GND.n5777 GND.n1965 14.8754
R9905 GND.n1976 GND.n1965 14.8754
R9906 GND.n1977 GND.n1976 14.8754
R9907 GND.n5771 GND.n1977 14.8754
R9908 GND.n5771 GND.n5770 14.8754
R9909 GND.n5770 GND.n1979 14.8754
R9910 GND.n4925 GND.n1979 14.8754
R9911 GND.n4925 GND.n1990 14.8754
R9912 GND.n5764 GND.n1990 14.8754
R9913 GND.n5764 GND.n5763 14.8754
R9914 GND.n5763 GND.n1992 14.8754
R9915 GND.n2003 GND.n1992 14.8754
R9916 GND.n2004 GND.n2003 14.8754
R9917 GND.n5757 GND.n2004 14.8754
R9918 GND.n5757 GND.n5756 14.8754
R9919 GND.n2692 GND.n2691 14.8754
R9920 GND.n2692 GND.n2016 14.8754
R9921 GND.n5750 GND.n2016 14.8754
R9922 GND.n5750 GND.n5749 14.8754
R9923 GND.n5749 GND.n2018 14.8754
R9924 GND.n2029 GND.n2018 14.8754
R9925 GND.n2030 GND.n2029 14.8754
R9926 GND.n5743 GND.n2030 14.8754
R9927 GND.n5743 GND.n5742 14.8754
R9928 GND.n5742 GND.n2032 14.8754
R9929 GND.n4947 GND.n2032 14.8754
R9930 GND.n4947 GND.n2043 14.8754
R9931 GND.n5736 GND.n2043 14.8754
R9932 GND.n5736 GND.n5735 14.8754
R9933 GND.n5735 GND.n2045 14.8754
R9934 GND.n2056 GND.n2045 14.8754
R9935 GND.n2057 GND.n2056 14.8754
R9936 GND.n5729 GND.n2057 14.8754
R9937 GND.n5729 GND.n5728 14.8754
R9938 GND.n5728 GND.n2059 14.8754
R9939 GND.n4958 GND.n2059 14.8754
R9940 GND.n4958 GND.n2070 14.8754
R9941 GND.n5722 GND.n2070 14.8754
R9942 GND.n5722 GND.n5721 14.8754
R9943 GND.n5721 GND.n2072 14.8754
R9944 GND.n2083 GND.n2072 14.8754
R9945 GND.n2084 GND.n2083 14.8754
R9946 GND.n5715 GND.n2084 14.8754
R9947 GND.n5715 GND.n5714 14.8754
R9948 GND.n5714 GND.n2086 14.8754
R9949 GND.n4969 GND.n2097 14.8754
R9950 GND.n5708 GND.n2097 14.8754
R9951 GND.n5708 GND.n5707 14.8754
R9952 GND.n5707 GND.n2099 14.8754
R9953 GND.n2110 GND.n2099 14.8754
R9954 GND.n2111 GND.n2110 14.8754
R9955 GND.n5701 GND.n2111 14.8754
R9956 GND.n5701 GND.n5700 14.8754
R9957 GND.n5700 GND.n2113 14.8754
R9958 GND.n2679 GND.n2113 14.8754
R9959 GND.n2679 GND.n2124 14.8754
R9960 GND.n5694 GND.n2124 14.8754
R9961 GND.n5694 GND.n5693 14.8754
R9962 GND.n5693 GND.n2126 14.8754
R9963 GND.n2137 GND.n2126 14.8754
R9964 GND.n2138 GND.n2137 14.8754
R9965 GND.n5687 GND.n2138 14.8754
R9966 GND.n5687 GND.n5686 14.8754
R9967 GND.n5686 GND.n2140 14.8754
R9968 GND.n4991 GND.n2140 14.8754
R9969 GND.n4991 GND.n2151 14.8754
R9970 GND.n5680 GND.n2151 14.8754
R9971 GND.n5680 GND.n5679 14.8754
R9972 GND.n5679 GND.n2153 14.8754
R9973 GND.n2164 GND.n2153 14.8754
R9974 GND.n2165 GND.n2164 14.8754
R9975 GND.n5673 GND.n2165 14.8754
R9976 GND.n5673 GND.n5672 14.8754
R9977 GND.n5672 GND.n2167 14.8754
R9978 GND.n5003 GND.n2167 14.8754
R9979 GND.n5003 GND.n5002 14.8754
R9980 GND.n5666 GND.n5665 14.8754
R9981 GND.n5665 GND.n2179 14.8754
R9982 GND.n2190 GND.n2179 14.8754
R9983 GND.n2191 GND.n2190 14.8754
R9984 GND.n5659 GND.n2191 14.8754
R9985 GND.n5659 GND.n5658 14.8754
R9986 GND.n5658 GND.n2193 14.8754
R9987 GND.n5014 GND.n2193 14.8754
R9988 GND.n5014 GND.n2204 14.8754
R9989 GND.n5652 GND.n2204 14.8754
R9990 GND.n5652 GND.n5651 14.8754
R9991 GND.n5651 GND.n2206 14.8754
R9992 GND.n2217 GND.n2206 14.8754
R9993 GND.n2218 GND.n2217 14.8754
R9994 GND.n5645 GND.n2218 14.8754
R9995 GND.n6144 GND.n1649 14.2804
R9996 GND.n4754 GND.n4753 14.2804
R9997 GND.n6075 GND.n6074 14.2804
R9998 GND.n6026 GND.n6025 14.2804
R9999 GND.n1629 GND.n1622 14.2723
R10000 GND.n5860 GND.n5859 14.2723
R10001 GND.n4013 GND.t0 13.9829
R10002 GND.n5110 GND.t6 13.9829
R10003 GND.n6102 GND.n1722 13.6854
R10004 GND.n4846 GND.n4845 13.6854
R10005 GND.n4868 GND.n2721 13.6854
R10006 GND.n4344 GND.t13 13.3879
R10007 GND.n4538 GND.t20 13.3879
R10008 GND.n6215 GND.n1613 13.3879
R10009 GND.n6012 GND.n6011 13.3879
R10010 GND.t167 GND.n5798 13.3879
R10011 GND.t4 GND.n2086 13.3879
R10012 GND.n1646 GND.n1617 13.1884
R10013 GND.n1641 GND.n1640 13.1884
R10014 GND.n1640 GND.n1639 13.1884
R10015 GND.n1635 GND.n1634 13.1884
R10016 GND.n1634 GND.n1633 13.1884
R10017 GND.n5845 GND.n5840 13.1884
R10018 GND.n5846 GND.n5845 13.1884
R10019 GND.n5851 GND.n5838 13.1884
R10020 GND.n5852 GND.n5851 13.1884
R10021 GND.n6212 GND.n6148 13.1127
R10022 GND.n5936 GND.n5935 13.1127
R10023 GND.n2766 GND.n2765 13.0904
R10024 GND.n2752 GND.n1748 13.0904
R10025 GND.n6068 GND.n1782 13.0904
R10026 GND.n6032 GND.n1826 13.0904
R10027 GND.t63 GND.n3486 12.7929
R10028 GND.n5312 GND.t67 12.7929
R10029 GND.n4184 GND.n4183 12.4954
R10030 GND.n4691 GND.n1680 12.4954
R10031 GND.n4877 GND.n2713 12.4954
R10032 GND.t91 GND.n5833 12.4954
R10033 GND.n5644 GND.n5643 12.4954
R10034 GND.n2759 GND.n1682 11.9004
R10035 GND.n6096 GND.n1728 11.9004
R10036 GND.n6061 GND.n6060 11.9004
R10037 GND.n1912 GND.t115 11.9004
R10038 GND.n4763 GND.t169 11.6029
R10039 GND.t23 GND.n1784 11.6029
R10040 GND.n6130 GND.n1669 11.3054
R10041 GND.n2755 GND.n1750 11.3054
R10042 GND.n4812 GND.n2741 11.3054
R10043 GND.n5821 GND.n5818 11.3054
R10044 GND.t154 GND.n3008 11.0079
R10045 GND.n5002 GND.t164 11.0079
R10046 GND.n6115 GND.n1699 10.7104
R10047 GND.n4727 GND.n4726 10.7104
R10048 GND.n6054 GND.n1800 10.7104
R10049 GND.n6046 GND.n1809 10.7104
R10050 GND.t109 GND.n2722 10.7104
R10051 GND.n6008 GND.n6007 10.6151
R10052 GND.n6007 GND.n6004 10.6151
R10053 GND.n6002 GND.n5999 10.6151
R10054 GND.n5999 GND.n5998 10.6151
R10055 GND.n5998 GND.n5995 10.6151
R10056 GND.n5995 GND.n5994 10.6151
R10057 GND.n5994 GND.n5991 10.6151
R10058 GND.n5991 GND.n5990 10.6151
R10059 GND.n5990 GND.n5987 10.6151
R10060 GND.n5987 GND.n5986 10.6151
R10061 GND.n5986 GND.n5983 10.6151
R10062 GND.n5983 GND.n5982 10.6151
R10063 GND.n5982 GND.n5979 10.6151
R10064 GND.n5979 GND.n5978 10.6151
R10065 GND.n5978 GND.n5975 10.6151
R10066 GND.n5975 GND.n5974 10.6151
R10067 GND.n5974 GND.n5971 10.6151
R10068 GND.n5971 GND.n5970 10.6151
R10069 GND.n5970 GND.n5967 10.6151
R10070 GND.n5967 GND.n5966 10.6151
R10071 GND.n5966 GND.n5963 10.6151
R10072 GND.n5963 GND.n5962 10.6151
R10073 GND.n5962 GND.n5959 10.6151
R10074 GND.n5959 GND.n5958 10.6151
R10075 GND.n5958 GND.n5955 10.6151
R10076 GND.n5955 GND.n5954 10.6151
R10077 GND.n5954 GND.n5951 10.6151
R10078 GND.n5951 GND.n5950 10.6151
R10079 GND.n5950 GND.n5947 10.6151
R10080 GND.n5947 GND.n5946 10.6151
R10081 GND.n5946 GND.n5943 10.6151
R10082 GND.n5943 GND.n5942 10.6151
R10083 GND.n4650 GND.n4649 10.6151
R10084 GND.n4649 GND.n2769 10.6151
R10085 GND.n4669 GND.n2769 10.6151
R10086 GND.n4670 GND.n4669 10.6151
R10087 GND.n4674 GND.n4670 10.6151
R10088 GND.n4675 GND.n4674 10.6151
R10089 GND.n4676 GND.n4675 10.6151
R10090 GND.n4680 GND.n4676 10.6151
R10091 GND.n4680 GND.n4679 10.6151
R10092 GND.n4679 GND.n4678 10.6151
R10093 GND.n4678 GND.n2757 10.6151
R10094 GND.n4717 GND.n2757 10.6151
R10095 GND.n4718 GND.n4717 10.6151
R10096 GND.n4721 GND.n4718 10.6151
R10097 GND.n4722 GND.n4721 10.6151
R10098 GND.n4723 GND.n4722 10.6151
R10099 GND.n4729 GND.n4723 10.6151
R10100 GND.n4730 GND.n4729 10.6151
R10101 GND.n4733 GND.n4730 10.6151
R10102 GND.n4734 GND.n4733 10.6151
R10103 GND.n4737 GND.n4734 10.6151
R10104 GND.n4738 GND.n4737 10.6151
R10105 GND.n4739 GND.n4738 10.6151
R10106 GND.n4742 GND.n4739 10.6151
R10107 GND.n4743 GND.n4742 10.6151
R10108 GND.n4751 GND.n4743 10.6151
R10109 GND.n4751 GND.n4750 10.6151
R10110 GND.n4750 GND.n4749 10.6151
R10111 GND.n4749 GND.n4745 10.6151
R10112 GND.n4745 GND.n4744 10.6151
R10113 GND.n4744 GND.n2739 10.6151
R10114 GND.n4815 GND.n2739 10.6151
R10115 GND.n4816 GND.n4815 10.6151
R10116 GND.n4820 GND.n4816 10.6151
R10117 GND.n4821 GND.n4820 10.6151
R10118 GND.n4822 GND.n4821 10.6151
R10119 GND.n4839 GND.n4822 10.6151
R10120 GND.n4839 GND.n4838 10.6151
R10121 GND.n4838 GND.n4837 10.6151
R10122 GND.n4837 GND.n4836 10.6151
R10123 GND.n4836 GND.n4834 10.6151
R10124 GND.n4834 GND.n4833 10.6151
R10125 GND.n4833 GND.n4823 10.6151
R10126 GND.n4829 GND.n4823 10.6151
R10127 GND.n4829 GND.n4828 10.6151
R10128 GND.n4828 GND.n4827 10.6151
R10129 GND.n4827 GND.n4825 10.6151
R10130 GND.n4825 GND.n4824 10.6151
R10131 GND.n4824 GND.n1894 10.6151
R10132 GND.n5824 GND.n1894 10.6151
R10133 GND.n5825 GND.n5824 10.6151
R10134 GND.n5829 GND.n5825 10.6151
R10135 GND.n5830 GND.n5829 10.6151
R10136 GND.n5831 GND.n5830 10.6151
R10137 GND.n5831 GND.n1893 10.6151
R10138 GND.n4583 GND.n1573 10.6151
R10139 GND.n4586 GND.n4583 10.6151
R10140 GND.n4591 GND.n4588 10.6151
R10141 GND.n4592 GND.n4591 10.6151
R10142 GND.n4595 GND.n4592 10.6151
R10143 GND.n4596 GND.n4595 10.6151
R10144 GND.n4599 GND.n4596 10.6151
R10145 GND.n4600 GND.n4599 10.6151
R10146 GND.n4603 GND.n4600 10.6151
R10147 GND.n4604 GND.n4603 10.6151
R10148 GND.n4607 GND.n4604 10.6151
R10149 GND.n4608 GND.n4607 10.6151
R10150 GND.n4611 GND.n4608 10.6151
R10151 GND.n4612 GND.n4611 10.6151
R10152 GND.n4615 GND.n4612 10.6151
R10153 GND.n4616 GND.n4615 10.6151
R10154 GND.n4619 GND.n4616 10.6151
R10155 GND.n4620 GND.n4619 10.6151
R10156 GND.n4623 GND.n4620 10.6151
R10157 GND.n4624 GND.n4623 10.6151
R10158 GND.n4627 GND.n4624 10.6151
R10159 GND.n4628 GND.n4627 10.6151
R10160 GND.n4631 GND.n4628 10.6151
R10161 GND.n4632 GND.n4631 10.6151
R10162 GND.n4635 GND.n4632 10.6151
R10163 GND.n4636 GND.n4635 10.6151
R10164 GND.n4639 GND.n4636 10.6151
R10165 GND.n4640 GND.n4639 10.6151
R10166 GND.n4643 GND.n4640 10.6151
R10167 GND.n4644 GND.n4643 10.6151
R10168 GND.n4647 GND.n4644 10.6151
R10169 GND.n4648 GND.n4647 10.6151
R10170 GND.n6212 GND.n6211 10.6151
R10171 GND.n6211 GND.n6210 10.6151
R10172 GND.n6210 GND.n6209 10.6151
R10173 GND.n6209 GND.n6207 10.6151
R10174 GND.n6207 GND.n6204 10.6151
R10175 GND.n6204 GND.n6203 10.6151
R10176 GND.n6203 GND.n6200 10.6151
R10177 GND.n6200 GND.n6199 10.6151
R10178 GND.n6199 GND.n6196 10.6151
R10179 GND.n6196 GND.n6195 10.6151
R10180 GND.n6195 GND.n6192 10.6151
R10181 GND.n6192 GND.n6191 10.6151
R10182 GND.n6191 GND.n6188 10.6151
R10183 GND.n6188 GND.n6187 10.6151
R10184 GND.n6187 GND.n6184 10.6151
R10185 GND.n6184 GND.n6183 10.6151
R10186 GND.n6183 GND.n6180 10.6151
R10187 GND.n6180 GND.n6179 10.6151
R10188 GND.n6179 GND.n6176 10.6151
R10189 GND.n6176 GND.n6175 10.6151
R10190 GND.n6175 GND.n6172 10.6151
R10191 GND.n6172 GND.n6171 10.6151
R10192 GND.n6171 GND.n6168 10.6151
R10193 GND.n6168 GND.n6167 10.6151
R10194 GND.n6167 GND.n6164 10.6151
R10195 GND.n6164 GND.n6163 10.6151
R10196 GND.n6163 GND.n6160 10.6151
R10197 GND.n6160 GND.n6159 10.6151
R10198 GND.n6159 GND.n6156 10.6151
R10199 GND.n6156 GND.n6155 10.6151
R10200 GND.n6152 GND.n1576 10.6151
R10201 GND.n6218 GND.n1576 10.6151
R10202 GND.n5935 GND.n5934 10.6151
R10203 GND.n5934 GND.n5931 10.6151
R10204 GND.n5931 GND.n5930 10.6151
R10205 GND.n5930 GND.n5927 10.6151
R10206 GND.n5927 GND.n5926 10.6151
R10207 GND.n5926 GND.n5923 10.6151
R10208 GND.n5923 GND.n5922 10.6151
R10209 GND.n5922 GND.n5919 10.6151
R10210 GND.n5919 GND.n5918 10.6151
R10211 GND.n5918 GND.n5915 10.6151
R10212 GND.n5915 GND.n5914 10.6151
R10213 GND.n5914 GND.n5911 10.6151
R10214 GND.n5911 GND.n5910 10.6151
R10215 GND.n5910 GND.n5907 10.6151
R10216 GND.n5907 GND.n5906 10.6151
R10217 GND.n5906 GND.n5903 10.6151
R10218 GND.n5903 GND.n5902 10.6151
R10219 GND.n5902 GND.n5899 10.6151
R10220 GND.n5899 GND.n5898 10.6151
R10221 GND.n5898 GND.n5895 10.6151
R10222 GND.n5895 GND.n5894 10.6151
R10223 GND.n5894 GND.n5891 10.6151
R10224 GND.n5891 GND.n5890 10.6151
R10225 GND.n5890 GND.n5887 10.6151
R10226 GND.n5887 GND.n5886 10.6151
R10227 GND.n5886 GND.n5883 10.6151
R10228 GND.n5883 GND.n5882 10.6151
R10229 GND.n5882 GND.n5879 10.6151
R10230 GND.n5879 GND.n5878 10.6151
R10231 GND.n5878 GND.n5875 10.6151
R10232 GND.n5873 GND.n5870 10.6151
R10233 GND.n5870 GND.n5869 10.6151
R10234 GND.n6147 GND.n6146 10.6151
R10235 GND.n6146 GND.n1647 10.6151
R10236 GND.n1666 GND.n1647 10.6151
R10237 GND.n6134 GND.n1666 10.6151
R10238 GND.n6134 GND.n6133 10.6151
R10239 GND.n6133 GND.n6132 10.6151
R10240 GND.n6132 GND.n1667 10.6151
R10241 GND.n4688 GND.n1667 10.6151
R10242 GND.n4688 GND.n4687 10.6151
R10243 GND.n4687 GND.n4686 10.6151
R10244 GND.n4686 GND.n4683 10.6151
R10245 GND.n4683 GND.n1702 10.6151
R10246 GND.n6113 GND.n1702 10.6151
R10247 GND.n6113 GND.n6112 10.6151
R10248 GND.n6112 GND.n6111 10.6151
R10249 GND.n6111 GND.n1703 10.6151
R10250 GND.n1725 GND.n1703 10.6151
R10251 GND.n6100 GND.n1725 10.6151
R10252 GND.n6100 GND.n6099 10.6151
R10253 GND.n6099 GND.n6098 10.6151
R10254 GND.n6098 GND.n1726 10.6151
R10255 GND.n4760 GND.n1726 10.6151
R10256 GND.n4760 GND.n4759 10.6151
R10257 GND.n4759 GND.n4758 10.6151
R10258 GND.n4758 GND.n2754 10.6151
R10259 GND.n2754 GND.n1769 10.6151
R10260 GND.n6079 GND.n1769 10.6151
R10261 GND.n6079 GND.n6078 10.6151
R10262 GND.n6078 GND.n6077 10.6151
R10263 GND.n6077 GND.n1770 10.6151
R10264 GND.n4810 GND.n1770 10.6151
R10265 GND.n4810 GND.n1787 10.6151
R10266 GND.n6065 GND.n1787 10.6151
R10267 GND.n6065 GND.n6064 10.6151
R10268 GND.n6064 GND.n6063 10.6151
R10269 GND.n6063 GND.n1788 10.6151
R10270 GND.n4843 GND.n1788 10.6151
R10271 GND.n4843 GND.n1804 10.6151
R10272 GND.n6051 GND.n1804 10.6151
R10273 GND.n6051 GND.n6050 10.6151
R10274 GND.n6050 GND.n6049 10.6151
R10275 GND.n6049 GND.n1805 10.6151
R10276 GND.n2719 GND.n1805 10.6151
R10277 GND.n2719 GND.n1822 10.6151
R10278 GND.n6037 GND.n1822 10.6151
R10279 GND.n6037 GND.n6036 10.6151
R10280 GND.n6036 GND.n6035 10.6151
R10281 GND.n6035 GND.n1823 10.6151
R10282 GND.n5819 GND.n1823 10.6151
R10283 GND.n5819 GND.n1839 10.6151
R10284 GND.n6023 GND.n1839 10.6151
R10285 GND.n6023 GND.n6022 10.6151
R10286 GND.n6022 GND.n6021 10.6151
R10287 GND.n6021 GND.n1840 10.6151
R10288 GND.n5937 GND.n1840 10.6151
R10289 GND.n6220 GND.n1568 10.4732
R10290 GND.n5521 GND.n5520 10.4732
R10291 GND.n1638 GND.n1619 10.2247
R10292 GND.n1636 GND.n1621 10.2247
R10293 GND.n5844 GND.n5839 10.2247
R10294 GND.n5850 GND.n5849 10.2247
R10295 GND.n4667 GND.n4666 10.1154
R10296 GND.n6136 GND.t106 10.1154
R10297 GND.t148 GND.n4714 10.1154
R10298 GND.n6081 GND.n1766 10.1154
R10299 GND.n4747 GND.n1766 10.1154
R10300 GND.n6019 GND.n1842 10.1154
R10301 GND.n6247 GND.n6246 9.89141
R10302 GND.n5556 GND.n5555 9.89141
R10303 GND.n7982 GND.n180 9.89141
R10304 GND.n7949 GND.n7948 9.89141
R10305 GND.n3621 GND.n3618 9.89141
R10306 GND.n3667 GND.n3559 9.89141
R10307 GND.n5597 GND.n5594 9.69747
R10308 GND.n3141 GND.n3140 9.69747
R10309 GND.t57 GND.n6122 9.52045
R10310 GND.n4719 GND.n1699 9.52045
R10311 GND.n4726 GND.n4725 9.52045
R10312 GND.n6054 GND.n6053 9.52045
R10313 GND.n6047 GND.n6046 9.52045
R10314 GND.n6629 GND.n1086 9.3005
R10315 GND.n6631 GND.n6630 9.3005
R10316 GND.n1082 GND.n1081 9.3005
R10317 GND.n6638 GND.n6637 9.3005
R10318 GND.n6639 GND.n1080 9.3005
R10319 GND.n6641 GND.n6640 9.3005
R10320 GND.n1076 GND.n1075 9.3005
R10321 GND.n6648 GND.n6647 9.3005
R10322 GND.n6649 GND.n1074 9.3005
R10323 GND.n6651 GND.n6650 9.3005
R10324 GND.n1070 GND.n1069 9.3005
R10325 GND.n6658 GND.n6657 9.3005
R10326 GND.n6659 GND.n1068 9.3005
R10327 GND.n6661 GND.n6660 9.3005
R10328 GND.n1064 GND.n1063 9.3005
R10329 GND.n6668 GND.n6667 9.3005
R10330 GND.n6669 GND.n1062 9.3005
R10331 GND.n6671 GND.n6670 9.3005
R10332 GND.n1058 GND.n1057 9.3005
R10333 GND.n6678 GND.n6677 9.3005
R10334 GND.n6679 GND.n1056 9.3005
R10335 GND.n6681 GND.n6680 9.3005
R10336 GND.n1052 GND.n1051 9.3005
R10337 GND.n6688 GND.n6687 9.3005
R10338 GND.n6689 GND.n1050 9.3005
R10339 GND.n6691 GND.n6690 9.3005
R10340 GND.n1046 GND.n1045 9.3005
R10341 GND.n6698 GND.n6697 9.3005
R10342 GND.n6699 GND.n1044 9.3005
R10343 GND.n6701 GND.n6700 9.3005
R10344 GND.n1040 GND.n1039 9.3005
R10345 GND.n6708 GND.n6707 9.3005
R10346 GND.n6709 GND.n1038 9.3005
R10347 GND.n6711 GND.n6710 9.3005
R10348 GND.n1034 GND.n1033 9.3005
R10349 GND.n6718 GND.n6717 9.3005
R10350 GND.n6719 GND.n1032 9.3005
R10351 GND.n6721 GND.n6720 9.3005
R10352 GND.n1028 GND.n1027 9.3005
R10353 GND.n6728 GND.n6727 9.3005
R10354 GND.n6729 GND.n1026 9.3005
R10355 GND.n6731 GND.n6730 9.3005
R10356 GND.n1022 GND.n1021 9.3005
R10357 GND.n6738 GND.n6737 9.3005
R10358 GND.n6739 GND.n1020 9.3005
R10359 GND.n6741 GND.n6740 9.3005
R10360 GND.n1016 GND.n1015 9.3005
R10361 GND.n6748 GND.n6747 9.3005
R10362 GND.n6749 GND.n1014 9.3005
R10363 GND.n6751 GND.n6750 9.3005
R10364 GND.n1010 GND.n1009 9.3005
R10365 GND.n6758 GND.n6757 9.3005
R10366 GND.n6759 GND.n1008 9.3005
R10367 GND.n6761 GND.n6760 9.3005
R10368 GND.n1004 GND.n1003 9.3005
R10369 GND.n6768 GND.n6767 9.3005
R10370 GND.n6769 GND.n1002 9.3005
R10371 GND.n6771 GND.n6770 9.3005
R10372 GND.n998 GND.n997 9.3005
R10373 GND.n6778 GND.n6777 9.3005
R10374 GND.n6779 GND.n996 9.3005
R10375 GND.n6781 GND.n6780 9.3005
R10376 GND.n992 GND.n991 9.3005
R10377 GND.n6788 GND.n6787 9.3005
R10378 GND.n6789 GND.n990 9.3005
R10379 GND.n6791 GND.n6790 9.3005
R10380 GND.n986 GND.n985 9.3005
R10381 GND.n6798 GND.n6797 9.3005
R10382 GND.n6799 GND.n984 9.3005
R10383 GND.n6801 GND.n6800 9.3005
R10384 GND.n980 GND.n979 9.3005
R10385 GND.n6808 GND.n6807 9.3005
R10386 GND.n6809 GND.n978 9.3005
R10387 GND.n6811 GND.n6810 9.3005
R10388 GND.n974 GND.n973 9.3005
R10389 GND.n6818 GND.n6817 9.3005
R10390 GND.n6819 GND.n972 9.3005
R10391 GND.n6821 GND.n6820 9.3005
R10392 GND.n968 GND.n967 9.3005
R10393 GND.n6828 GND.n6827 9.3005
R10394 GND.n6829 GND.n966 9.3005
R10395 GND.n6831 GND.n6830 9.3005
R10396 GND.n962 GND.n961 9.3005
R10397 GND.n6838 GND.n6837 9.3005
R10398 GND.n6839 GND.n960 9.3005
R10399 GND.n6841 GND.n6840 9.3005
R10400 GND.n956 GND.n955 9.3005
R10401 GND.n6848 GND.n6847 9.3005
R10402 GND.n6849 GND.n954 9.3005
R10403 GND.n6851 GND.n6850 9.3005
R10404 GND.n950 GND.n949 9.3005
R10405 GND.n6858 GND.n6857 9.3005
R10406 GND.n6859 GND.n948 9.3005
R10407 GND.n6861 GND.n6860 9.3005
R10408 GND.n944 GND.n943 9.3005
R10409 GND.n6868 GND.n6867 9.3005
R10410 GND.n6869 GND.n942 9.3005
R10411 GND.n6871 GND.n6870 9.3005
R10412 GND.n938 GND.n937 9.3005
R10413 GND.n6878 GND.n6877 9.3005
R10414 GND.n6879 GND.n936 9.3005
R10415 GND.n6881 GND.n6880 9.3005
R10416 GND.n932 GND.n931 9.3005
R10417 GND.n6888 GND.n6887 9.3005
R10418 GND.n6889 GND.n930 9.3005
R10419 GND.n6891 GND.n6890 9.3005
R10420 GND.n926 GND.n925 9.3005
R10421 GND.n6898 GND.n6897 9.3005
R10422 GND.n6899 GND.n924 9.3005
R10423 GND.n6901 GND.n6900 9.3005
R10424 GND.n920 GND.n919 9.3005
R10425 GND.n6908 GND.n6907 9.3005
R10426 GND.n6909 GND.n918 9.3005
R10427 GND.n6911 GND.n6910 9.3005
R10428 GND.n914 GND.n913 9.3005
R10429 GND.n6918 GND.n6917 9.3005
R10430 GND.n6919 GND.n912 9.3005
R10431 GND.n6921 GND.n6920 9.3005
R10432 GND.n908 GND.n907 9.3005
R10433 GND.n6928 GND.n6927 9.3005
R10434 GND.n6929 GND.n906 9.3005
R10435 GND.n6931 GND.n6930 9.3005
R10436 GND.n902 GND.n901 9.3005
R10437 GND.n6938 GND.n6937 9.3005
R10438 GND.n6939 GND.n900 9.3005
R10439 GND.n6941 GND.n6940 9.3005
R10440 GND.n896 GND.n895 9.3005
R10441 GND.n6948 GND.n6947 9.3005
R10442 GND.n6949 GND.n894 9.3005
R10443 GND.n6951 GND.n6950 9.3005
R10444 GND.n890 GND.n889 9.3005
R10445 GND.n6958 GND.n6957 9.3005
R10446 GND.n6959 GND.n888 9.3005
R10447 GND.n6961 GND.n6960 9.3005
R10448 GND.n884 GND.n883 9.3005
R10449 GND.n6968 GND.n6967 9.3005
R10450 GND.n6969 GND.n882 9.3005
R10451 GND.n6971 GND.n6970 9.3005
R10452 GND.n878 GND.n877 9.3005
R10453 GND.n6978 GND.n6977 9.3005
R10454 GND.n6979 GND.n876 9.3005
R10455 GND.n6981 GND.n6980 9.3005
R10456 GND.n872 GND.n871 9.3005
R10457 GND.n6988 GND.n6987 9.3005
R10458 GND.n6989 GND.n870 9.3005
R10459 GND.n6991 GND.n6990 9.3005
R10460 GND.n866 GND.n865 9.3005
R10461 GND.n6998 GND.n6997 9.3005
R10462 GND.n6999 GND.n864 9.3005
R10463 GND.n7001 GND.n7000 9.3005
R10464 GND.n860 GND.n859 9.3005
R10465 GND.n7008 GND.n7007 9.3005
R10466 GND.n7009 GND.n858 9.3005
R10467 GND.n7011 GND.n7010 9.3005
R10468 GND.n854 GND.n853 9.3005
R10469 GND.n7018 GND.n7017 9.3005
R10470 GND.n7019 GND.n852 9.3005
R10471 GND.n7021 GND.n7020 9.3005
R10472 GND.n848 GND.n847 9.3005
R10473 GND.n7028 GND.n7027 9.3005
R10474 GND.n7029 GND.n846 9.3005
R10475 GND.n7031 GND.n7030 9.3005
R10476 GND.n842 GND.n841 9.3005
R10477 GND.n7038 GND.n7037 9.3005
R10478 GND.n7039 GND.n840 9.3005
R10479 GND.n7041 GND.n7040 9.3005
R10480 GND.n836 GND.n835 9.3005
R10481 GND.n7048 GND.n7047 9.3005
R10482 GND.n7049 GND.n834 9.3005
R10483 GND.n7051 GND.n7050 9.3005
R10484 GND.n830 GND.n829 9.3005
R10485 GND.n7058 GND.n7057 9.3005
R10486 GND.n7059 GND.n828 9.3005
R10487 GND.n7061 GND.n7060 9.3005
R10488 GND.n824 GND.n823 9.3005
R10489 GND.n7068 GND.n7067 9.3005
R10490 GND.n7069 GND.n822 9.3005
R10491 GND.n7071 GND.n7070 9.3005
R10492 GND.n818 GND.n817 9.3005
R10493 GND.n7078 GND.n7077 9.3005
R10494 GND.n7079 GND.n816 9.3005
R10495 GND.n7081 GND.n7080 9.3005
R10496 GND.n812 GND.n811 9.3005
R10497 GND.n7088 GND.n7087 9.3005
R10498 GND.n7089 GND.n810 9.3005
R10499 GND.n7091 GND.n7090 9.3005
R10500 GND.n806 GND.n805 9.3005
R10501 GND.n7098 GND.n7097 9.3005
R10502 GND.n7099 GND.n804 9.3005
R10503 GND.n7101 GND.n7100 9.3005
R10504 GND.n800 GND.n799 9.3005
R10505 GND.n7108 GND.n7107 9.3005
R10506 GND.n7109 GND.n798 9.3005
R10507 GND.n7111 GND.n7110 9.3005
R10508 GND.n794 GND.n793 9.3005
R10509 GND.n7118 GND.n7117 9.3005
R10510 GND.n7119 GND.n792 9.3005
R10511 GND.n7121 GND.n7120 9.3005
R10512 GND.n788 GND.n787 9.3005
R10513 GND.n7128 GND.n7127 9.3005
R10514 GND.n7129 GND.n786 9.3005
R10515 GND.n7131 GND.n7130 9.3005
R10516 GND.n782 GND.n781 9.3005
R10517 GND.n7138 GND.n7137 9.3005
R10518 GND.n7139 GND.n780 9.3005
R10519 GND.n7141 GND.n7140 9.3005
R10520 GND.n776 GND.n775 9.3005
R10521 GND.n7148 GND.n7147 9.3005
R10522 GND.n7149 GND.n774 9.3005
R10523 GND.n7151 GND.n7150 9.3005
R10524 GND.n770 GND.n769 9.3005
R10525 GND.n7158 GND.n7157 9.3005
R10526 GND.n7159 GND.n768 9.3005
R10527 GND.n7161 GND.n7160 9.3005
R10528 GND.n764 GND.n763 9.3005
R10529 GND.n7168 GND.n7167 9.3005
R10530 GND.n7169 GND.n762 9.3005
R10531 GND.n7171 GND.n7170 9.3005
R10532 GND.n758 GND.n757 9.3005
R10533 GND.n7178 GND.n7177 9.3005
R10534 GND.n7179 GND.n756 9.3005
R10535 GND.n7181 GND.n7180 9.3005
R10536 GND.n752 GND.n751 9.3005
R10537 GND.n7188 GND.n7187 9.3005
R10538 GND.n7189 GND.n750 9.3005
R10539 GND.n7191 GND.n7190 9.3005
R10540 GND.n746 GND.n745 9.3005
R10541 GND.n7198 GND.n7197 9.3005
R10542 GND.n7199 GND.n744 9.3005
R10543 GND.n7201 GND.n7200 9.3005
R10544 GND.n740 GND.n739 9.3005
R10545 GND.n7208 GND.n7207 9.3005
R10546 GND.n7209 GND.n738 9.3005
R10547 GND.n7211 GND.n7210 9.3005
R10548 GND.n734 GND.n733 9.3005
R10549 GND.n7218 GND.n7217 9.3005
R10550 GND.n7219 GND.n732 9.3005
R10551 GND.n7221 GND.n7220 9.3005
R10552 GND.n728 GND.n727 9.3005
R10553 GND.n7228 GND.n7227 9.3005
R10554 GND.n7229 GND.n726 9.3005
R10555 GND.n7231 GND.n7230 9.3005
R10556 GND.n722 GND.n721 9.3005
R10557 GND.n7238 GND.n7237 9.3005
R10558 GND.n7239 GND.n720 9.3005
R10559 GND.n7241 GND.n7240 9.3005
R10560 GND.n716 GND.n715 9.3005
R10561 GND.n7248 GND.n7247 9.3005
R10562 GND.n7249 GND.n714 9.3005
R10563 GND.n7251 GND.n7250 9.3005
R10564 GND.n710 GND.n709 9.3005
R10565 GND.n7258 GND.n7257 9.3005
R10566 GND.n7259 GND.n708 9.3005
R10567 GND.n7261 GND.n7260 9.3005
R10568 GND.n704 GND.n703 9.3005
R10569 GND.n7268 GND.n7267 9.3005
R10570 GND.n7269 GND.n702 9.3005
R10571 GND.n7271 GND.n7270 9.3005
R10572 GND.n698 GND.n697 9.3005
R10573 GND.n7278 GND.n7277 9.3005
R10574 GND.n7279 GND.n696 9.3005
R10575 GND.n7281 GND.n7280 9.3005
R10576 GND.n692 GND.n691 9.3005
R10577 GND.n7288 GND.n7287 9.3005
R10578 GND.n7289 GND.n690 9.3005
R10579 GND.n7291 GND.n7290 9.3005
R10580 GND.n686 GND.n685 9.3005
R10581 GND.n7298 GND.n7297 9.3005
R10582 GND.n7299 GND.n684 9.3005
R10583 GND.n7301 GND.n7300 9.3005
R10584 GND.n680 GND.n679 9.3005
R10585 GND.n7308 GND.n7307 9.3005
R10586 GND.n7309 GND.n678 9.3005
R10587 GND.n7311 GND.n7310 9.3005
R10588 GND.n674 GND.n673 9.3005
R10589 GND.n7318 GND.n7317 9.3005
R10590 GND.n7319 GND.n672 9.3005
R10591 GND.n7321 GND.n7320 9.3005
R10592 GND.n668 GND.n667 9.3005
R10593 GND.n7328 GND.n7327 9.3005
R10594 GND.n7329 GND.n666 9.3005
R10595 GND.n7331 GND.n7330 9.3005
R10596 GND.n662 GND.n661 9.3005
R10597 GND.n7338 GND.n7337 9.3005
R10598 GND.n7339 GND.n660 9.3005
R10599 GND.n7341 GND.n7340 9.3005
R10600 GND.n656 GND.n655 9.3005
R10601 GND.n7348 GND.n7347 9.3005
R10602 GND.n7349 GND.n654 9.3005
R10603 GND.n7351 GND.n7350 9.3005
R10604 GND.n650 GND.n649 9.3005
R10605 GND.n7358 GND.n7357 9.3005
R10606 GND.n7359 GND.n648 9.3005
R10607 GND.n7361 GND.n7360 9.3005
R10608 GND.n644 GND.n643 9.3005
R10609 GND.n7368 GND.n7367 9.3005
R10610 GND.n7369 GND.n642 9.3005
R10611 GND.n7371 GND.n7370 9.3005
R10612 GND.n638 GND.n637 9.3005
R10613 GND.n7378 GND.n7377 9.3005
R10614 GND.n7379 GND.n636 9.3005
R10615 GND.n7381 GND.n7380 9.3005
R10616 GND.n632 GND.n631 9.3005
R10617 GND.n7388 GND.n7387 9.3005
R10618 GND.n7389 GND.n630 9.3005
R10619 GND.n7391 GND.n7390 9.3005
R10620 GND.n626 GND.n625 9.3005
R10621 GND.n7398 GND.n7397 9.3005
R10622 GND.n7399 GND.n624 9.3005
R10623 GND.n7401 GND.n7400 9.3005
R10624 GND.n620 GND.n619 9.3005
R10625 GND.n7408 GND.n7407 9.3005
R10626 GND.n7409 GND.n618 9.3005
R10627 GND.n7411 GND.n7410 9.3005
R10628 GND.n614 GND.n613 9.3005
R10629 GND.n7418 GND.n7417 9.3005
R10630 GND.n7419 GND.n612 9.3005
R10631 GND.n7421 GND.n7420 9.3005
R10632 GND.n608 GND.n607 9.3005
R10633 GND.n7428 GND.n7427 9.3005
R10634 GND.n7429 GND.n606 9.3005
R10635 GND.n7431 GND.n7430 9.3005
R10636 GND.n602 GND.n601 9.3005
R10637 GND.n7438 GND.n7437 9.3005
R10638 GND.n7439 GND.n600 9.3005
R10639 GND.n7441 GND.n7440 9.3005
R10640 GND.n596 GND.n595 9.3005
R10641 GND.n7448 GND.n7447 9.3005
R10642 GND.n7449 GND.n594 9.3005
R10643 GND.n7451 GND.n7450 9.3005
R10644 GND.n590 GND.n589 9.3005
R10645 GND.n7458 GND.n7457 9.3005
R10646 GND.n7459 GND.n588 9.3005
R10647 GND.n7461 GND.n7460 9.3005
R10648 GND.n584 GND.n583 9.3005
R10649 GND.n7468 GND.n7467 9.3005
R10650 GND.n7469 GND.n582 9.3005
R10651 GND.n7471 GND.n7470 9.3005
R10652 GND.n578 GND.n577 9.3005
R10653 GND.n7478 GND.n7477 9.3005
R10654 GND.n7479 GND.n576 9.3005
R10655 GND.n7481 GND.n7480 9.3005
R10656 GND.n572 GND.n571 9.3005
R10657 GND.n7488 GND.n7487 9.3005
R10658 GND.n7489 GND.n570 9.3005
R10659 GND.n7491 GND.n7490 9.3005
R10660 GND.n566 GND.n565 9.3005
R10661 GND.n7498 GND.n7497 9.3005
R10662 GND.n7499 GND.n564 9.3005
R10663 GND.n7501 GND.n7500 9.3005
R10664 GND.n560 GND.n559 9.3005
R10665 GND.n7508 GND.n7507 9.3005
R10666 GND.n7509 GND.n558 9.3005
R10667 GND.n7511 GND.n7510 9.3005
R10668 GND.n554 GND.n553 9.3005
R10669 GND.n7518 GND.n7517 9.3005
R10670 GND.n7519 GND.n552 9.3005
R10671 GND.n7521 GND.n7520 9.3005
R10672 GND.n548 GND.n547 9.3005
R10673 GND.n7528 GND.n7527 9.3005
R10674 GND.n7529 GND.n546 9.3005
R10675 GND.n7531 GND.n7530 9.3005
R10676 GND.n542 GND.n541 9.3005
R10677 GND.n7538 GND.n7537 9.3005
R10678 GND.n7539 GND.n540 9.3005
R10679 GND.n7541 GND.n7540 9.3005
R10680 GND.n536 GND.n535 9.3005
R10681 GND.n7548 GND.n7547 9.3005
R10682 GND.n7549 GND.n534 9.3005
R10683 GND.n7551 GND.n7550 9.3005
R10684 GND.n530 GND.n529 9.3005
R10685 GND.n7558 GND.n7557 9.3005
R10686 GND.n7559 GND.n528 9.3005
R10687 GND.n7561 GND.n7560 9.3005
R10688 GND.n524 GND.n523 9.3005
R10689 GND.n7568 GND.n7567 9.3005
R10690 GND.n7569 GND.n522 9.3005
R10691 GND.n7571 GND.n7570 9.3005
R10692 GND.n518 GND.n517 9.3005
R10693 GND.n7578 GND.n7577 9.3005
R10694 GND.n7579 GND.n516 9.3005
R10695 GND.n7581 GND.n7580 9.3005
R10696 GND.n512 GND.n511 9.3005
R10697 GND.n7588 GND.n7587 9.3005
R10698 GND.n7589 GND.n510 9.3005
R10699 GND.n7591 GND.n7590 9.3005
R10700 GND.n7598 GND.n7597 9.3005
R10701 GND.n7599 GND.n504 9.3005
R10702 GND.n7601 GND.n7600 9.3005
R10703 GND.n500 GND.n499 9.3005
R10704 GND.n7608 GND.n7607 9.3005
R10705 GND.n7609 GND.n498 9.3005
R10706 GND.n7611 GND.n7610 9.3005
R10707 GND.n494 GND.n493 9.3005
R10708 GND.n7618 GND.n7617 9.3005
R10709 GND.n7619 GND.n492 9.3005
R10710 GND.n7621 GND.n7620 9.3005
R10711 GND.n488 GND.n487 9.3005
R10712 GND.n7628 GND.n7627 9.3005
R10713 GND.n7629 GND.n486 9.3005
R10714 GND.n7631 GND.n7630 9.3005
R10715 GND.n482 GND.n481 9.3005
R10716 GND.n7638 GND.n7637 9.3005
R10717 GND.n7639 GND.n480 9.3005
R10718 GND.n7641 GND.n7640 9.3005
R10719 GND.n476 GND.n475 9.3005
R10720 GND.n7648 GND.n7647 9.3005
R10721 GND.n7649 GND.n474 9.3005
R10722 GND.n7651 GND.n7650 9.3005
R10723 GND.n470 GND.n469 9.3005
R10724 GND.n7658 GND.n7657 9.3005
R10725 GND.n7659 GND.n468 9.3005
R10726 GND.n7661 GND.n7660 9.3005
R10727 GND.n464 GND.n463 9.3005
R10728 GND.n7668 GND.n7667 9.3005
R10729 GND.n7669 GND.n462 9.3005
R10730 GND.n7671 GND.n7670 9.3005
R10731 GND.n458 GND.n457 9.3005
R10732 GND.n7678 GND.n7677 9.3005
R10733 GND.n7679 GND.n456 9.3005
R10734 GND.n7681 GND.n7680 9.3005
R10735 GND.n452 GND.n451 9.3005
R10736 GND.n7688 GND.n7687 9.3005
R10737 GND.n7689 GND.n450 9.3005
R10738 GND.n7691 GND.n7690 9.3005
R10739 GND.n446 GND.n445 9.3005
R10740 GND.n7698 GND.n7697 9.3005
R10741 GND.n7699 GND.n444 9.3005
R10742 GND.n7701 GND.n7700 9.3005
R10743 GND.n440 GND.n439 9.3005
R10744 GND.n7708 GND.n7707 9.3005
R10745 GND.n7709 GND.n438 9.3005
R10746 GND.n7711 GND.n7710 9.3005
R10747 GND.n434 GND.n433 9.3005
R10748 GND.n7718 GND.n7717 9.3005
R10749 GND.n7719 GND.n432 9.3005
R10750 GND.n7721 GND.n7720 9.3005
R10751 GND.n428 GND.n427 9.3005
R10752 GND.n7728 GND.n7727 9.3005
R10753 GND.n7729 GND.n426 9.3005
R10754 GND.n7731 GND.n7730 9.3005
R10755 GND.n422 GND.n421 9.3005
R10756 GND.n7738 GND.n7737 9.3005
R10757 GND.n7739 GND.n420 9.3005
R10758 GND.n7742 GND.n7741 9.3005
R10759 GND.n7740 GND.n416 9.3005
R10760 GND.n7748 GND.n415 9.3005
R10761 GND.n7750 GND.n7749 9.3005
R10762 GND.n506 GND.n505 9.3005
R10763 GND.n3028 GND.n3027 9.3005
R10764 GND.n4208 GND.n4207 9.3005
R10765 GND.n4209 GND.n3026 9.3005
R10766 GND.n4213 GND.n4210 9.3005
R10767 GND.n4212 GND.n4211 9.3005
R10768 GND.n3005 GND.n3004 9.3005
R10769 GND.n4240 GND.n4239 9.3005
R10770 GND.n4241 GND.n3003 9.3005
R10771 GND.n4245 GND.n4242 9.3005
R10772 GND.n4244 GND.n4243 9.3005
R10773 GND.n2982 GND.n2981 9.3005
R10774 GND.n4272 GND.n4271 9.3005
R10775 GND.n4273 GND.n2980 9.3005
R10776 GND.n4277 GND.n4274 9.3005
R10777 GND.n4276 GND.n4275 9.3005
R10778 GND.n2959 GND.n2958 9.3005
R10779 GND.n4304 GND.n4303 9.3005
R10780 GND.n4305 GND.n2957 9.3005
R10781 GND.n4309 GND.n4306 9.3005
R10782 GND.n4308 GND.n4307 9.3005
R10783 GND.n2935 GND.n2934 9.3005
R10784 GND.n4336 GND.n4335 9.3005
R10785 GND.n4337 GND.n2933 9.3005
R10786 GND.n4341 GND.n4338 9.3005
R10787 GND.n4340 GND.n4339 9.3005
R10788 GND.n2913 GND.n2912 9.3005
R10789 GND.n4368 GND.n4367 9.3005
R10790 GND.n4369 GND.n2911 9.3005
R10791 GND.n4373 GND.n4370 9.3005
R10792 GND.n4372 GND.n4371 9.3005
R10793 GND.n2890 GND.n2889 9.3005
R10794 GND.n4400 GND.n4399 9.3005
R10795 GND.n4401 GND.n2888 9.3005
R10796 GND.n4405 GND.n4402 9.3005
R10797 GND.n4404 GND.n4403 9.3005
R10798 GND.n2867 GND.n2866 9.3005
R10799 GND.n4432 GND.n4431 9.3005
R10800 GND.n4433 GND.n2865 9.3005
R10801 GND.n4437 GND.n4434 9.3005
R10802 GND.n4436 GND.n4435 9.3005
R10803 GND.n2844 GND.n2843 9.3005
R10804 GND.n4464 GND.n4463 9.3005
R10805 GND.n4465 GND.n2842 9.3005
R10806 GND.n4469 GND.n4466 9.3005
R10807 GND.n4468 GND.n4467 9.3005
R10808 GND.n2821 GND.n2820 9.3005
R10809 GND.n4496 GND.n4495 9.3005
R10810 GND.n4497 GND.n2819 9.3005
R10811 GND.n4501 GND.n4498 9.3005
R10812 GND.n4500 GND.n4499 9.3005
R10813 GND.n2798 GND.n2797 9.3005
R10814 GND.n4528 GND.n4527 9.3005
R10815 GND.n4529 GND.n2796 9.3005
R10816 GND.n4536 GND.n4530 9.3005
R10817 GND.n4535 GND.n4531 9.3005
R10818 GND.n4534 GND.n4533 9.3005
R10819 GND.n4532 GND.n2776 9.3005
R10820 GND.n2774 GND.n2773 9.3005
R10821 GND.n4656 GND.n4655 9.3005
R10822 GND.n4657 GND.n2772 9.3005
R10823 GND.n4664 GND.n4658 9.3005
R10824 GND.n4663 GND.n4659 9.3005
R10825 GND.n4662 GND.n4660 9.3005
R10826 GND.n2763 GND.n2762 9.3005
R10827 GND.n4694 GND.n4693 9.3005
R10828 GND.n4695 GND.n2761 9.3005
R10829 GND.n4712 GND.n4696 9.3005
R10830 GND.n4711 GND.n4697 9.3005
R10831 GND.n4710 GND.n4698 9.3005
R10832 GND.n4701 GND.n4699 9.3005
R10833 GND.n4706 GND.n4702 9.3005
R10834 GND.n4705 GND.n4704 9.3005
R10835 GND.n4703 GND.n2750 9.3005
R10836 GND.n4765 GND.n2749 9.3005
R10837 GND.n4767 GND.n4766 9.3005
R10838 GND.n4768 GND.n2748 9.3005
R10839 GND.n4770 GND.n4769 9.3005
R10840 GND.n2746 GND.n2745 9.3005
R10841 GND.n4775 GND.n4774 9.3005
R10842 GND.n4776 GND.n2744 9.3005
R10843 GND.n4787 GND.n4777 9.3005
R10844 GND.n4786 GND.n4778 9.3005
R10845 GND.n4785 GND.n4779 9.3005
R10846 GND.n4783 GND.n4780 9.3005
R10847 GND.n4782 GND.n4781 9.3005
R10848 GND.n2727 GND.n2726 9.3005
R10849 GND.n4860 GND.n4859 9.3005
R10850 GND.n4861 GND.n2725 9.3005
R10851 GND.n4866 GND.n4862 9.3005
R10852 GND.n4865 GND.n4864 9.3005
R10853 GND.n4863 GND.n2710 9.3005
R10854 GND.n4881 GND.n2709 9.3005
R10855 GND.n4883 GND.n4882 9.3005
R10856 GND.n4884 GND.n2708 9.3005
R10857 GND.n4886 GND.n4885 9.3005
R10858 GND.n2706 GND.n2705 9.3005
R10859 GND.n4892 GND.n4891 9.3005
R10860 GND.n4893 GND.n2704 9.3005
R10861 GND.n4895 GND.n4894 9.3005
R10862 GND.n4896 GND.n2703 9.3005
R10863 GND.n4900 GND.n4899 9.3005
R10864 GND.n4901 GND.n2702 9.3005
R10865 GND.n4905 GND.n4902 9.3005
R10866 GND.n4906 GND.n2701 9.3005
R10867 GND.n4910 GND.n4909 9.3005
R10868 GND.n4911 GND.n2700 9.3005
R10869 GND.n4913 GND.n4912 9.3005
R10870 GND.n4916 GND.n2699 9.3005
R10871 GND.n4918 GND.n4917 9.3005
R10872 GND.n4919 GND.n2698 9.3005
R10873 GND.n4923 GND.n4920 9.3005
R10874 GND.n4924 GND.n2697 9.3005
R10875 GND.n4928 GND.n4927 9.3005
R10876 GND.n4929 GND.n2696 9.3005
R10877 GND.n4931 GND.n4930 9.3005
R10878 GND.n4934 GND.n2695 9.3005
R10879 GND.n4936 GND.n4935 9.3005
R10880 GND.n4937 GND.n2694 9.3005
R10881 GND.n4939 GND.n4938 9.3005
R10882 GND.n4940 GND.n2690 9.3005
R10883 GND.n4944 GND.n4943 9.3005
R10884 GND.n4945 GND.n2689 9.3005
R10885 GND.n4949 GND.n4946 9.3005
R10886 GND.n4950 GND.n2688 9.3005
R10887 GND.n4954 GND.n4953 9.3005
R10888 GND.n4955 GND.n2687 9.3005
R10889 GND.n4957 GND.n4956 9.3005
R10890 GND.n4960 GND.n2686 9.3005
R10891 GND.n4962 GND.n4961 9.3005
R10892 GND.n4963 GND.n2685 9.3005
R10893 GND.n4967 GND.n4964 9.3005
R10894 GND.n4968 GND.n2684 9.3005
R10895 GND.n4972 GND.n4971 9.3005
R10896 GND.n4973 GND.n2683 9.3005
R10897 GND.n4975 GND.n4974 9.3005
R10898 GND.n4978 GND.n2682 9.3005
R10899 GND.n4980 GND.n4979 9.3005
R10900 GND.n4981 GND.n2681 9.3005
R10901 GND.n4983 GND.n4982 9.3005
R10902 GND.n4984 GND.n2678 9.3005
R10903 GND.n4988 GND.n4987 9.3005
R10904 GND.n4989 GND.n2677 9.3005
R10905 GND.n4993 GND.n4990 9.3005
R10906 GND.n4994 GND.n2676 9.3005
R10907 GND.n4998 GND.n4997 9.3005
R10908 GND.n4999 GND.n2675 9.3005
R10909 GND.n5001 GND.n5000 9.3005
R10910 GND.n5005 GND.n2674 9.3005
R10911 GND.n5007 GND.n5006 9.3005
R10912 GND.n5008 GND.n2673 9.3005
R10913 GND.n5012 GND.n5009 9.3005
R10914 GND.n5013 GND.n2672 9.3005
R10915 GND.n5017 GND.n5016 9.3005
R10916 GND.n5018 GND.n2671 9.3005
R10917 GND.n5020 GND.n5019 9.3005
R10918 GND.n5021 GND.n2667 9.3005
R10919 GND.n3121 GND.n3120 9.3005
R10920 GND.n4161 GND.n4160 9.3005
R10921 GND.n4164 GND.n3070 9.3005
R10922 GND.n4165 GND.n3069 9.3005
R10923 GND.n4168 GND.n3068 9.3005
R10924 GND.n4169 GND.n3067 9.3005
R10925 GND.n4172 GND.n3066 9.3005
R10926 GND.n4173 GND.n3065 9.3005
R10927 GND.n4176 GND.n3064 9.3005
R10928 GND.n4178 GND.n3063 9.3005
R10929 GND.n4179 GND.n3062 9.3005
R10930 GND.n4180 GND.n3061 9.3005
R10931 GND.n3060 GND.n3035 9.3005
R10932 GND.n4199 GND.n3034 9.3005
R10933 GND.n4203 GND.n4200 9.3005
R10934 GND.n4202 GND.n4201 9.3005
R10935 GND.n3013 GND.n3012 9.3005
R10936 GND.n4230 GND.n4229 9.3005
R10937 GND.n4231 GND.n3011 9.3005
R10938 GND.n4235 GND.n4232 9.3005
R10939 GND.n4234 GND.n4233 9.3005
R10940 GND.n2990 GND.n2989 9.3005
R10941 GND.n4262 GND.n4261 9.3005
R10942 GND.n4263 GND.n2988 9.3005
R10943 GND.n4267 GND.n4264 9.3005
R10944 GND.n4266 GND.n4265 9.3005
R10945 GND.n2967 GND.n2966 9.3005
R10946 GND.n4294 GND.n4293 9.3005
R10947 GND.n4295 GND.n2965 9.3005
R10948 GND.n4299 GND.n4296 9.3005
R10949 GND.n4298 GND.n4297 9.3005
R10950 GND.n2944 GND.n2943 9.3005
R10951 GND.n4326 GND.n4325 9.3005
R10952 GND.n4327 GND.n2942 9.3005
R10953 GND.n4331 GND.n4328 9.3005
R10954 GND.n4330 GND.n4329 9.3005
R10955 GND.n2921 GND.n2920 9.3005
R10956 GND.n4358 GND.n4357 9.3005
R10957 GND.n4359 GND.n2919 9.3005
R10958 GND.n4363 GND.n4360 9.3005
R10959 GND.n4362 GND.n4361 9.3005
R10960 GND.n2898 GND.n2897 9.3005
R10961 GND.n4390 GND.n4389 9.3005
R10962 GND.n4391 GND.n2896 9.3005
R10963 GND.n4395 GND.n4392 9.3005
R10964 GND.n4394 GND.n4393 9.3005
R10965 GND.n2875 GND.n2874 9.3005
R10966 GND.n4422 GND.n4421 9.3005
R10967 GND.n4423 GND.n2873 9.3005
R10968 GND.n4427 GND.n4424 9.3005
R10969 GND.n4426 GND.n4425 9.3005
R10970 GND.n2852 GND.n2851 9.3005
R10971 GND.n4454 GND.n4453 9.3005
R10972 GND.n4455 GND.n2850 9.3005
R10973 GND.n4459 GND.n4456 9.3005
R10974 GND.n4458 GND.n4457 9.3005
R10975 GND.n2829 GND.n2828 9.3005
R10976 GND.n4486 GND.n4485 9.3005
R10977 GND.n4487 GND.n2827 9.3005
R10978 GND.n4491 GND.n4488 9.3005
R10979 GND.n4490 GND.n4489 9.3005
R10980 GND.n2806 GND.n2805 9.3005
R10981 GND.n4518 GND.n4517 9.3005
R10982 GND.n4519 GND.n2804 9.3005
R10983 GND.n4523 GND.n4520 9.3005
R10984 GND.n4522 GND.n4521 9.3005
R10985 GND.n2783 GND.n2782 9.3005
R10986 GND.n4569 GND.n4568 9.3005
R10987 GND.n4570 GND.n2781 9.3005
R10988 GND.n4575 GND.n4571 9.3005
R10989 GND.n4574 GND.n4573 9.3005
R10990 GND.n4572 GND.n1655 9.3005
R10991 GND.n6141 GND.n1656 9.3005
R10992 GND.n6140 GND.n1657 9.3005
R10993 GND.n6139 GND.n1658 9.3005
R10994 GND.n1686 GND.n1659 9.3005
R10995 GND.n1689 GND.n1688 9.3005
R10996 GND.n1690 GND.n1685 9.3005
R10997 GND.n6120 GND.n1691 9.3005
R10998 GND.n6119 GND.n1692 9.3005
R10999 GND.n6118 GND.n1693 9.3005
R11000 GND.n1735 GND.n1694 9.3005
R11001 GND.n1737 GND.n1736 9.3005
R11002 GND.n1741 GND.n1740 9.3005
R11003 GND.n1742 GND.n1734 9.3005
R11004 GND.n6093 GND.n1743 9.3005
R11005 GND.n6092 GND.n1744 9.3005
R11006 GND.n6091 GND.n1745 9.3005
R11007 GND.n4794 GND.n1746 9.3005
R11008 GND.n4796 GND.n4795 9.3005
R11009 GND.n4793 GND.n4792 9.3005
R11010 GND.n4801 GND.n4800 9.3005
R11011 GND.n4802 GND.n4791 9.3005
R11012 GND.n4806 GND.n4803 9.3005
R11013 GND.n4805 GND.n4804 9.3005
R11014 GND.n2734 GND.n2733 9.3005
R11015 GND.n4849 GND.n4848 9.3005
R11016 GND.n4850 GND.n2732 9.3005
R11017 GND.n4854 GND.n4851 9.3005
R11018 GND.n4853 GND.n4852 9.3005
R11019 GND.n2717 GND.n2716 9.3005
R11020 GND.n4871 GND.n4870 9.3005
R11021 GND.n4872 GND.n2715 9.3005
R11022 GND.n4875 GND.n4874 9.3005
R11023 GND.n4873 GND.n1900 9.3005
R11024 GND.n5816 GND.n1901 9.3005
R11025 GND.n5815 GND.n1902 9.3005
R11026 GND.n5814 GND.n1903 9.3005
R11027 GND.n1906 GND.n1904 9.3005
R11028 GND.n5810 GND.n1907 9.3005
R11029 GND.n5809 GND.n1908 9.3005
R11030 GND.n5808 GND.n1909 9.3005
R11031 GND.n1929 GND.n1910 9.3005
R11032 GND.n1930 GND.n1928 9.3005
R11033 GND.n5796 GND.n1931 9.3005
R11034 GND.n5795 GND.n1932 9.3005
R11035 GND.n5794 GND.n1933 9.3005
R11036 GND.n1956 GND.n1934 9.3005
R11037 GND.n1957 GND.n1955 9.3005
R11038 GND.n5782 GND.n1958 9.3005
R11039 GND.n5781 GND.n1959 9.3005
R11040 GND.n5780 GND.n1960 9.3005
R11041 GND.n1983 GND.n1961 9.3005
R11042 GND.n1984 GND.n1982 9.3005
R11043 GND.n5768 GND.n1985 9.3005
R11044 GND.n5767 GND.n1986 9.3005
R11045 GND.n5766 GND.n1987 9.3005
R11046 GND.n2009 GND.n1988 9.3005
R11047 GND.n2010 GND.n2008 9.3005
R11048 GND.n5754 GND.n2011 9.3005
R11049 GND.n5753 GND.n2012 9.3005
R11050 GND.n5752 GND.n2013 9.3005
R11051 GND.n2036 GND.n2014 9.3005
R11052 GND.n2037 GND.n2035 9.3005
R11053 GND.n5740 GND.n2038 9.3005
R11054 GND.n5739 GND.n2039 9.3005
R11055 GND.n5738 GND.n2040 9.3005
R11056 GND.n2063 GND.n2041 9.3005
R11057 GND.n2064 GND.n2062 9.3005
R11058 GND.n5726 GND.n2065 9.3005
R11059 GND.n5725 GND.n2066 9.3005
R11060 GND.n5724 GND.n2067 9.3005
R11061 GND.n2090 GND.n2068 9.3005
R11062 GND.n2091 GND.n2089 9.3005
R11063 GND.n5712 GND.n2092 9.3005
R11064 GND.n5711 GND.n2093 9.3005
R11065 GND.n5710 GND.n2094 9.3005
R11066 GND.n2117 GND.n2095 9.3005
R11067 GND.n2118 GND.n2116 9.3005
R11068 GND.n5698 GND.n2119 9.3005
R11069 GND.n5697 GND.n2120 9.3005
R11070 GND.n5696 GND.n2121 9.3005
R11071 GND.n2144 GND.n2122 9.3005
R11072 GND.n2145 GND.n2143 9.3005
R11073 GND.n5684 GND.n2146 9.3005
R11074 GND.n5683 GND.n2147 9.3005
R11075 GND.n5682 GND.n2148 9.3005
R11076 GND.n2171 GND.n2149 9.3005
R11077 GND.n2172 GND.n2170 9.3005
R11078 GND.n5670 GND.n2173 9.3005
R11079 GND.n5669 GND.n2174 9.3005
R11080 GND.n5668 GND.n2175 9.3005
R11081 GND.n2197 GND.n2176 9.3005
R11082 GND.n2198 GND.n2196 9.3005
R11083 GND.n5656 GND.n2199 9.3005
R11084 GND.n5655 GND.n2200 9.3005
R11085 GND.n5654 GND.n2201 9.3005
R11086 GND.n2235 GND.n2202 9.3005
R11087 GND.n2237 GND.n2236 9.3005
R11088 GND.n4198 GND.n4197 9.3005
R11089 GND.n5640 GND.n5639 9.3005
R11090 GND.n5638 GND.n2239 9.3005
R11091 GND.n5637 GND.n5636 9.3005
R11092 GND.n5633 GND.n2240 9.3005
R11093 GND.n5630 GND.n2241 9.3005
R11094 GND.n5629 GND.n2242 9.3005
R11095 GND.n5626 GND.n2243 9.3005
R11096 GND.n5625 GND.n2244 9.3005
R11097 GND.n5622 GND.n2245 9.3005
R11098 GND.n5621 GND.n2246 9.3005
R11099 GND.n5618 GND.n2247 9.3005
R11100 GND.n5641 GND.n2238 9.3005
R11101 GND.n5039 GND.n5038 9.3005
R11102 GND.n5036 GND.n2665 9.3005
R11103 GND.n5035 GND.n5034 9.3005
R11104 GND.n5031 GND.n5029 9.3005
R11105 GND.n2669 GND.n2265 9.3005
R11106 GND.n5592 GND.n5591 9.3005
R11107 GND.n2264 GND.n2262 9.3005
R11108 GND.n2416 GND.n2415 9.3005
R11109 GND.n2419 GND.n2414 9.3005
R11110 GND.n2420 GND.n2413 9.3005
R11111 GND.n2423 GND.n2412 9.3005
R11112 GND.n2424 GND.n2411 9.3005
R11113 GND.n2427 GND.n2410 9.3005
R11114 GND.n2428 GND.n2409 9.3005
R11115 GND.n2431 GND.n2408 9.3005
R11116 GND.n2432 GND.n2407 9.3005
R11117 GND.n5617 GND.n2248 9.3005
R11118 GND.n5614 GND.n2249 9.3005
R11119 GND.n5613 GND.n2250 9.3005
R11120 GND.n5610 GND.n2251 9.3005
R11121 GND.n5609 GND.n2252 9.3005
R11122 GND.n5606 GND.n2253 9.3005
R11123 GND.n5605 GND.n2254 9.3005
R11124 GND.n5602 GND.n2255 9.3005
R11125 GND.n5601 GND.n2256 9.3005
R11126 GND.n5598 GND.n2257 9.3005
R11127 GND.n5597 GND.n2258 9.3005
R11128 GND.n5594 GND.n5593 9.3005
R11129 GND.n2263 GND.n2259 9.3005
R11130 GND.n5028 GND.n5027 9.3005
R11131 GND.n5024 GND.n2668 9.3005
R11132 GND.n5040 GND.n2661 9.3005
R11133 GND.n5043 GND.n5042 9.3005
R11134 GND.n5046 GND.n2660 9.3005
R11135 GND.n5053 GND.n5052 9.3005
R11136 GND.n5054 GND.n2659 9.3005
R11137 GND.n5056 GND.n5055 9.3005
R11138 GND.n2577 GND.n2576 9.3005
R11139 GND.n5068 GND.n5067 9.3005
R11140 GND.n5069 GND.n2575 9.3005
R11141 GND.n5071 GND.n5070 9.3005
R11142 GND.n2573 GND.n2572 9.3005
R11143 GND.n5083 GND.n5082 9.3005
R11144 GND.n5084 GND.n2571 9.3005
R11145 GND.n5086 GND.n5085 9.3005
R11146 GND.n2569 GND.n2568 9.3005
R11147 GND.n5098 GND.n5097 9.3005
R11148 GND.n5099 GND.n2567 9.3005
R11149 GND.n5101 GND.n5100 9.3005
R11150 GND.n2565 GND.n2564 9.3005
R11151 GND.n5113 GND.n5112 9.3005
R11152 GND.n5114 GND.n2563 9.3005
R11153 GND.n5120 GND.n5115 9.3005
R11154 GND.n5119 GND.n5116 9.3005
R11155 GND.n5118 GND.n5117 9.3005
R11156 GND.n28 GND.n26 9.3005
R11157 GND.n5045 GND.n5044 9.3005
R11158 GND.n8081 GND.n8080 9.3005
R11159 GND.n29 GND.n27 9.3005
R11160 GND.n5138 GND.n5137 9.3005
R11161 GND.n5352 GND.n5139 9.3005
R11162 GND.n5351 GND.n5140 9.3005
R11163 GND.n5350 GND.n5141 9.3005
R11164 GND.n5205 GND.n5142 9.3005
R11165 GND.n5340 GND.n5206 9.3005
R11166 GND.n5339 GND.n5207 9.3005
R11167 GND.n5338 GND.n5208 9.3005
R11168 GND.n5212 GND.n5209 9.3005
R11169 GND.n5328 GND.n5213 9.3005
R11170 GND.n5327 GND.n5214 9.3005
R11171 GND.n5326 GND.n5215 9.3005
R11172 GND.n5219 GND.n5216 9.3005
R11173 GND.n5316 GND.n5220 9.3005
R11174 GND.n5315 GND.n5221 9.3005
R11175 GND.n5314 GND.n5222 9.3005
R11176 GND.n5226 GND.n5223 9.3005
R11177 GND.n5304 GND.n5227 9.3005
R11178 GND.n5303 GND.n5228 9.3005
R11179 GND.n5302 GND.n5229 9.3005
R11180 GND.n5297 GND.n5230 9.3005
R11181 GND.n5296 GND.n5295 9.3005
R11182 GND.n5255 GND.n5254 9.3005
R11183 GND.n5256 GND.n5248 9.3005
R11184 GND.n5258 GND.n5257 9.3005
R11185 GND.n5246 GND.n5245 9.3005
R11186 GND.n5265 GND.n5264 9.3005
R11187 GND.n5266 GND.n5244 9.3005
R11188 GND.n5268 GND.n5267 9.3005
R11189 GND.n5242 GND.n5241 9.3005
R11190 GND.n5275 GND.n5274 9.3005
R11191 GND.n5276 GND.n5240 9.3005
R11192 GND.n5278 GND.n5277 9.3005
R11193 GND.n5238 GND.n5237 9.3005
R11194 GND.n5285 GND.n5284 9.3005
R11195 GND.n5286 GND.n5236 9.3005
R11196 GND.n5288 GND.n5287 9.3005
R11197 GND.n5234 GND.n5231 9.3005
R11198 GND.n5294 GND.n5293 9.3005
R11199 GND.n5249 GND.n286 9.3005
R11200 GND.n153 GND.n152 9.3005
R11201 GND.n157 GND.n155 9.3005
R11202 GND.n8004 GND.n158 9.3005
R11203 GND.n8003 GND.n159 9.3005
R11204 GND.n8002 GND.n160 9.3005
R11205 GND.n164 GND.n161 9.3005
R11206 GND.n7997 GND.n165 9.3005
R11207 GND.n7996 GND.n166 9.3005
R11208 GND.n7995 GND.n167 9.3005
R11209 GND.n171 GND.n168 9.3005
R11210 GND.n7990 GND.n172 9.3005
R11211 GND.n7989 GND.n173 9.3005
R11212 GND.n7988 GND.n174 9.3005
R11213 GND.n178 GND.n175 9.3005
R11214 GND.n7983 GND.n179 9.3005
R11215 GND.n7982 GND.n7981 9.3005
R11216 GND.n7980 GND.n180 9.3005
R11217 GND.n7979 GND.n7978 9.3005
R11218 GND.n184 GND.n183 9.3005
R11219 GND.n189 GND.n187 9.3005
R11220 GND.n7971 GND.n190 9.3005
R11221 GND.n7970 GND.n191 9.3005
R11222 GND.n7969 GND.n192 9.3005
R11223 GND.n196 GND.n193 9.3005
R11224 GND.n7964 GND.n197 9.3005
R11225 GND.n7963 GND.n198 9.3005
R11226 GND.n7962 GND.n199 9.3005
R11227 GND.n203 GND.n200 9.3005
R11228 GND.n7957 GND.n204 9.3005
R11229 GND.n7956 GND.n205 9.3005
R11230 GND.n7955 GND.n206 9.3005
R11231 GND.n210 GND.n207 9.3005
R11232 GND.n7950 GND.n211 9.3005
R11233 GND.n7949 GND.n212 9.3005
R11234 GND.n7948 GND.n7947 9.3005
R11235 GND.n7946 GND.n213 9.3005
R11236 GND.n7945 GND.n7944 9.3005
R11237 GND.n219 GND.n218 9.3005
R11238 GND.n7939 GND.n223 9.3005
R11239 GND.n7938 GND.n224 9.3005
R11240 GND.n7937 GND.n225 9.3005
R11241 GND.n229 GND.n226 9.3005
R11242 GND.n7932 GND.n230 9.3005
R11243 GND.n7931 GND.n231 9.3005
R11244 GND.n7930 GND.n232 9.3005
R11245 GND.n236 GND.n233 9.3005
R11246 GND.n7925 GND.n237 9.3005
R11247 GND.n7924 GND.n238 9.3005
R11248 GND.n7923 GND.n239 9.3005
R11249 GND.n243 GND.n240 9.3005
R11250 GND.n7918 GND.n244 9.3005
R11251 GND.n7917 GND.n245 9.3005
R11252 GND.n7916 GND.n246 9.3005
R11253 GND.n253 GND.n251 9.3005
R11254 GND.n7911 GND.n254 9.3005
R11255 GND.n7910 GND.n255 9.3005
R11256 GND.n7909 GND.n256 9.3005
R11257 GND.n260 GND.n257 9.3005
R11258 GND.n7904 GND.n261 9.3005
R11259 GND.n7903 GND.n262 9.3005
R11260 GND.n7902 GND.n263 9.3005
R11261 GND.n267 GND.n264 9.3005
R11262 GND.n7897 GND.n268 9.3005
R11263 GND.n7896 GND.n269 9.3005
R11264 GND.n7895 GND.n270 9.3005
R11265 GND.n274 GND.n271 9.3005
R11266 GND.n7890 GND.n275 9.3005
R11267 GND.n7889 GND.n276 9.3005
R11268 GND.n7888 GND.n277 9.3005
R11269 GND.n281 GND.n278 9.3005
R11270 GND.n7883 GND.n282 9.3005
R11271 GND.n7882 GND.n7881 9.3005
R11272 GND.n7880 GND.n283 9.3005
R11273 GND.n8012 GND.n8011 9.3005
R11274 GND.n2435 GND.n2401 9.3005
R11275 GND.n5047 GND.n2451 9.3005
R11276 GND.n5428 GND.n2452 9.3005
R11277 GND.n5427 GND.n2453 9.3005
R11278 GND.n5426 GND.n2454 9.3005
R11279 GND.n5062 GND.n2455 9.3005
R11280 GND.n5416 GND.n2472 9.3005
R11281 GND.n5415 GND.n2473 9.3005
R11282 GND.n5414 GND.n2474 9.3005
R11283 GND.n5077 GND.n2475 9.3005
R11284 GND.n5404 GND.n2493 9.3005
R11285 GND.n5403 GND.n2494 9.3005
R11286 GND.n5402 GND.n2495 9.3005
R11287 GND.n5092 GND.n2496 9.3005
R11288 GND.n5392 GND.n2514 9.3005
R11289 GND.n5391 GND.n2515 9.3005
R11290 GND.n5390 GND.n2516 9.3005
R11291 GND.n5107 GND.n2517 9.3005
R11292 GND.n5380 GND.n2533 9.3005
R11293 GND.n5379 GND.n2534 9.3005
R11294 GND.n5378 GND.n2535 9.3005
R11295 GND.n5127 GND.n2536 9.3005
R11296 GND.n5130 GND.n5128 9.3005
R11297 GND.n5132 GND.n5131 9.3005
R11298 GND.n2558 GND.n2557 9.3005
R11299 GND.n5359 GND.n5358 9.3005
R11300 GND.n2559 GND.n56 9.3005
R11301 GND.n8069 GND.n57 9.3005
R11302 GND.n8068 GND.n58 9.3005
R11303 GND.n8067 GND.n59 9.3005
R11304 GND.n5203 GND.n60 9.3005
R11305 GND.n8057 GND.n77 9.3005
R11306 GND.n8056 GND.n78 9.3005
R11307 GND.n8055 GND.n79 9.3005
R11308 GND.n5210 GND.n80 9.3005
R11309 GND.n8045 GND.n98 9.3005
R11310 GND.n8044 GND.n99 9.3005
R11311 GND.n8043 GND.n100 9.3005
R11312 GND.n5217 GND.n101 9.3005
R11313 GND.n8033 GND.n119 9.3005
R11314 GND.n8032 GND.n120 9.3005
R11315 GND.n8031 GND.n121 9.3005
R11316 GND.n5224 GND.n122 9.3005
R11317 GND.n8021 GND.n140 9.3005
R11318 GND.n8020 GND.n141 9.3005
R11319 GND.n8019 GND.n142 9.3005
R11320 GND.n7878 GND.n143 9.3005
R11321 GND.n5442 GND.n2400 9.3005
R11322 GND.n2402 GND.n2401 9.3005
R11323 GND.n5048 GND.n5047 9.3005
R11324 GND.n2658 GND.n2452 9.3005
R11325 GND.n5060 GND.n2453 9.3005
R11326 GND.n5061 GND.n2454 9.3005
R11327 GND.n5063 GND.n5062 9.3005
R11328 GND.n2574 GND.n2472 9.3005
R11329 GND.n5075 GND.n2473 9.3005
R11330 GND.n5076 GND.n2474 9.3005
R11331 GND.n5078 GND.n5077 9.3005
R11332 GND.n2570 GND.n2493 9.3005
R11333 GND.n5090 GND.n2494 9.3005
R11334 GND.n5091 GND.n2495 9.3005
R11335 GND.n5093 GND.n5092 9.3005
R11336 GND.n2566 GND.n2514 9.3005
R11337 GND.n5105 GND.n2515 9.3005
R11338 GND.n5106 GND.n2516 9.3005
R11339 GND.n5108 GND.n5107 9.3005
R11340 GND.n2562 GND.n2533 9.3005
R11341 GND.n5124 GND.n2534 9.3005
R11342 GND.n5125 GND.n2535 9.3005
R11343 GND.n5127 GND.n5126 9.3005
R11344 GND.n5128 GND.n2561 9.3005
R11345 GND.n5133 GND.n5132 9.3005
R11346 GND.n5135 GND.n2558 9.3005
R11347 GND.n5358 GND.n5357 9.3005
R11348 GND.n5356 GND.n2559 9.3005
R11349 GND.n5136 GND.n57 9.3005
R11350 GND.n5346 GND.n58 9.3005
R11351 GND.n5345 GND.n59 9.3005
R11352 GND.n5344 GND.n5203 9.3005
R11353 GND.n5204 GND.n77 9.3005
R11354 GND.n5334 GND.n78 9.3005
R11355 GND.n5333 GND.n79 9.3005
R11356 GND.n5332 GND.n5210 9.3005
R11357 GND.n5211 GND.n98 9.3005
R11358 GND.n5322 GND.n99 9.3005
R11359 GND.n5321 GND.n100 9.3005
R11360 GND.n5320 GND.n5217 9.3005
R11361 GND.n5218 GND.n119 9.3005
R11362 GND.n5310 GND.n120 9.3005
R11363 GND.n5309 GND.n121 9.3005
R11364 GND.n5308 GND.n5224 9.3005
R11365 GND.n5225 GND.n140 9.3005
R11366 GND.n5298 GND.n141 9.3005
R11367 GND.n287 GND.n142 9.3005
R11368 GND.n7878 GND.n7877 9.3005
R11369 GND.n5442 GND.n5441 9.3005
R11370 GND.n5448 GND.n5447 9.3005
R11371 GND.n5451 GND.n2394 9.3005
R11372 GND.n5452 GND.n2393 9.3005
R11373 GND.n5455 GND.n2392 9.3005
R11374 GND.n5456 GND.n2391 9.3005
R11375 GND.n5459 GND.n2390 9.3005
R11376 GND.n5460 GND.n2389 9.3005
R11377 GND.n5463 GND.n2388 9.3005
R11378 GND.n5464 GND.n2387 9.3005
R11379 GND.n5467 GND.n2386 9.3005
R11380 GND.n5468 GND.n2385 9.3005
R11381 GND.n5471 GND.n2384 9.3005
R11382 GND.n5472 GND.n2383 9.3005
R11383 GND.n5475 GND.n2382 9.3005
R11384 GND.n5476 GND.n2381 9.3005
R11385 GND.n5479 GND.n2380 9.3005
R11386 GND.n5480 GND.n2379 9.3005
R11387 GND.n5483 GND.n2378 9.3005
R11388 GND.n5485 GND.n2375 9.3005
R11389 GND.n5488 GND.n2374 9.3005
R11390 GND.n5489 GND.n2373 9.3005
R11391 GND.n5492 GND.n2372 9.3005
R11392 GND.n5493 GND.n2371 9.3005
R11393 GND.n5496 GND.n2370 9.3005
R11394 GND.n5497 GND.n2369 9.3005
R11395 GND.n5500 GND.n2368 9.3005
R11396 GND.n5501 GND.n2367 9.3005
R11397 GND.n5504 GND.n2366 9.3005
R11398 GND.n5505 GND.n2365 9.3005
R11399 GND.n5508 GND.n2364 9.3005
R11400 GND.n5509 GND.n2363 9.3005
R11401 GND.n5512 GND.n2362 9.3005
R11402 GND.n5513 GND.n2361 9.3005
R11403 GND.n5516 GND.n2360 9.3005
R11404 GND.n5517 GND.n2359 9.3005
R11405 GND.n5520 GND.n2358 9.3005
R11406 GND.n5522 GND.n2353 9.3005
R11407 GND.n5525 GND.n2352 9.3005
R11408 GND.n5526 GND.n2351 9.3005
R11409 GND.n5529 GND.n2350 9.3005
R11410 GND.n5530 GND.n2349 9.3005
R11411 GND.n5533 GND.n2348 9.3005
R11412 GND.n5534 GND.n2347 9.3005
R11413 GND.n5537 GND.n2346 9.3005
R11414 GND.n5538 GND.n2345 9.3005
R11415 GND.n5541 GND.n2344 9.3005
R11416 GND.n5542 GND.n2343 9.3005
R11417 GND.n5545 GND.n2342 9.3005
R11418 GND.n5546 GND.n2341 9.3005
R11419 GND.n5549 GND.n2340 9.3005
R11420 GND.n5550 GND.n2339 9.3005
R11421 GND.n5553 GND.n2338 9.3005
R11422 GND.n5555 GND.n2337 9.3005
R11423 GND.n5557 GND.n2332 9.3005
R11424 GND.n5560 GND.n2331 9.3005
R11425 GND.n5561 GND.n2330 9.3005
R11426 GND.n5564 GND.n2329 9.3005
R11427 GND.n5565 GND.n2328 9.3005
R11428 GND.n5568 GND.n2327 9.3005
R11429 GND.n5569 GND.n2326 9.3005
R11430 GND.n5572 GND.n2325 9.3005
R11431 GND.n5573 GND.n2324 9.3005
R11432 GND.n5576 GND.n2323 9.3005
R11433 GND.n5577 GND.n2322 9.3005
R11434 GND.n5580 GND.n2321 9.3005
R11435 GND.n5582 GND.n2320 9.3005
R11436 GND.n5583 GND.n2319 9.3005
R11437 GND.n5584 GND.n2318 9.3005
R11438 GND.n5585 GND.n2317 9.3005
R11439 GND.n5556 GND.n2334 9.3005
R11440 GND.n5446 GND.n2398 9.3005
R11441 GND.n5445 GND.n5444 9.3005
R11442 GND.n5434 GND.n2441 9.3005
R11443 GND.n5433 GND.n2442 9.3005
R11444 GND.n5432 GND.n2443 9.3005
R11445 GND.n2461 GND.n2444 9.3005
R11446 GND.n5422 GND.n2462 9.3005
R11447 GND.n5421 GND.n2463 9.3005
R11448 GND.n5420 GND.n2464 9.3005
R11449 GND.n2482 GND.n2465 9.3005
R11450 GND.n5410 GND.n2483 9.3005
R11451 GND.n5409 GND.n2484 9.3005
R11452 GND.n5408 GND.n2485 9.3005
R11453 GND.n2503 GND.n2486 9.3005
R11454 GND.n5398 GND.n2504 9.3005
R11455 GND.n5397 GND.n2505 9.3005
R11456 GND.n5396 GND.n2506 9.3005
R11457 GND.n2524 GND.n2507 9.3005
R11458 GND.n5386 GND.n2525 9.3005
R11459 GND.n5385 GND.n41 9.3005
R11460 GND.n48 GND.n40 9.3005
R11461 GND.n8063 GND.n67 9.3005
R11462 GND.n8062 GND.n68 9.3005
R11463 GND.n8061 GND.n69 9.3005
R11464 GND.n87 GND.n70 9.3005
R11465 GND.n8051 GND.n88 9.3005
R11466 GND.n8050 GND.n89 9.3005
R11467 GND.n8049 GND.n90 9.3005
R11468 GND.n108 GND.n91 9.3005
R11469 GND.n8039 GND.n109 9.3005
R11470 GND.n8038 GND.n110 9.3005
R11471 GND.n8037 GND.n111 9.3005
R11472 GND.n129 GND.n112 9.3005
R11473 GND.n8027 GND.n130 9.3005
R11474 GND.n8026 GND.n131 9.3005
R11475 GND.n8025 GND.n132 9.3005
R11476 GND.n150 GND.n133 9.3005
R11477 GND.n8015 GND.n151 9.3005
R11478 GND.n8014 GND.n8013 9.3005
R11479 GND.n2440 GND.n2439 9.3005
R11480 GND.n8074 GND.n45 9.3005
R11481 GND.n8074 GND.n8073 9.3005
R11482 GND.n3372 GND.n3371 9.3005
R11483 GND.n4027 GND.n4026 9.3005
R11484 GND.n4028 GND.n3370 9.3005
R11485 GND.n4032 GND.n4029 9.3005
R11486 GND.n4031 GND.n4030 9.3005
R11487 GND.n3343 GND.n3342 9.3005
R11488 GND.n4064 GND.n4063 9.3005
R11489 GND.n4065 GND.n3341 9.3005
R11490 GND.n4069 GND.n4066 9.3005
R11491 GND.n4068 GND.n4067 9.3005
R11492 GND.n3314 GND.n3313 9.3005
R11493 GND.n4101 GND.n4100 9.3005
R11494 GND.n4102 GND.n3312 9.3005
R11495 GND.n4128 GND.n4103 9.3005
R11496 GND.n4127 GND.n4104 9.3005
R11497 GND.n4126 GND.n4105 9.3005
R11498 GND.n4108 GND.n4106 9.3005
R11499 GND.n4122 GND.n4109 9.3005
R11500 GND.n4121 GND.n4110 9.3005
R11501 GND.n4120 GND.n4111 9.3005
R11502 GND.n4113 GND.n4112 9.3005
R11503 GND.n4115 GND.n4114 9.3005
R11504 GND.n3044 GND.n3043 9.3005
R11505 GND.n4187 GND.n4186 9.3005
R11506 GND.n4188 GND.n3042 9.3005
R11507 GND.n4192 GND.n4189 9.3005
R11508 GND.n4191 GND.n4190 9.3005
R11509 GND.n3022 GND.n3021 9.3005
R11510 GND.n4219 GND.n4218 9.3005
R11511 GND.n4220 GND.n3020 9.3005
R11512 GND.n4224 GND.n4221 9.3005
R11513 GND.n4223 GND.n4222 9.3005
R11514 GND.n2999 GND.n2998 9.3005
R11515 GND.n4251 GND.n4250 9.3005
R11516 GND.n4252 GND.n2997 9.3005
R11517 GND.n4256 GND.n4253 9.3005
R11518 GND.n4255 GND.n4254 9.3005
R11519 GND.n2976 GND.n2975 9.3005
R11520 GND.n4283 GND.n4282 9.3005
R11521 GND.n4284 GND.n2974 9.3005
R11522 GND.n4288 GND.n4285 9.3005
R11523 GND.n4287 GND.n4286 9.3005
R11524 GND.n2953 GND.n2952 9.3005
R11525 GND.n4315 GND.n4314 9.3005
R11526 GND.n4316 GND.n2951 9.3005
R11527 GND.n4320 GND.n4317 9.3005
R11528 GND.n4319 GND.n4318 9.3005
R11529 GND.n2930 GND.n2929 9.3005
R11530 GND.n4347 GND.n4346 9.3005
R11531 GND.n4348 GND.n2928 9.3005
R11532 GND.n4352 GND.n4349 9.3005
R11533 GND.n4351 GND.n4350 9.3005
R11534 GND.n2907 GND.n2906 9.3005
R11535 GND.n4379 GND.n4378 9.3005
R11536 GND.n4380 GND.n2905 9.3005
R11537 GND.n4384 GND.n4381 9.3005
R11538 GND.n4383 GND.n4382 9.3005
R11539 GND.n2884 GND.n2883 9.3005
R11540 GND.n4411 GND.n4410 9.3005
R11541 GND.n4412 GND.n2882 9.3005
R11542 GND.n4416 GND.n4413 9.3005
R11543 GND.n4415 GND.n4414 9.3005
R11544 GND.n2861 GND.n2860 9.3005
R11545 GND.n4443 GND.n4442 9.3005
R11546 GND.n4444 GND.n2859 9.3005
R11547 GND.n4448 GND.n4445 9.3005
R11548 GND.n4447 GND.n4446 9.3005
R11549 GND.n2838 GND.n2837 9.3005
R11550 GND.n4475 GND.n4474 9.3005
R11551 GND.n4476 GND.n2836 9.3005
R11552 GND.n4480 GND.n4477 9.3005
R11553 GND.n4479 GND.n4478 9.3005
R11554 GND.n2815 GND.n2814 9.3005
R11555 GND.n4507 GND.n4506 9.3005
R11556 GND.n4508 GND.n2813 9.3005
R11557 GND.n4512 GND.n4509 9.3005
R11558 GND.n4511 GND.n4510 9.3005
R11559 GND.n2792 GND.n2791 9.3005
R11560 GND.n4542 GND.n4541 9.3005
R11561 GND.n4543 GND.n2790 9.3005
R11562 GND.n4563 GND.n4544 9.3005
R11563 GND.n4562 GND.n4545 9.3005
R11564 GND.n4561 GND.n4546 9.3005
R11565 GND.n4549 GND.n4547 9.3005
R11566 GND.n4557 GND.n4550 9.3005
R11567 GND.n4556 GND.n4551 9.3005
R11568 GND.n4555 GND.n4553 9.3005
R11569 GND.n4552 GND.n1674 9.3005
R11570 GND.n6127 GND.n1675 9.3005
R11571 GND.n6126 GND.n1676 9.3005
R11572 GND.n6125 GND.n1677 9.3005
R11573 GND.n1710 GND.n1678 9.3005
R11574 GND.n1713 GND.n1712 9.3005
R11575 GND.n1714 GND.n1709 9.3005
R11576 GND.n6107 GND.n1715 9.3005
R11577 GND.n6106 GND.n1716 9.3005
R11578 GND.n6105 GND.n1717 9.3005
R11579 GND.n1754 GND.n1718 9.3005
R11580 GND.n1757 GND.n1756 9.3005
R11581 GND.n1758 GND.n1753 9.3005
R11582 GND.n6086 GND.n1759 9.3005
R11583 GND.n6085 GND.n1760 9.3005
R11584 GND.n6084 GND.n1761 9.3005
R11585 GND.n1776 GND.n1762 9.3005
R11586 GND.n6072 GND.n1777 9.3005
R11587 GND.n6071 GND.n1778 9.3005
R11588 GND.n6070 GND.n1779 9.3005
R11589 GND.n1794 GND.n1780 9.3005
R11590 GND.n6058 GND.n1795 9.3005
R11591 GND.n6057 GND.n1796 9.3005
R11592 GND.n6056 GND.n1797 9.3005
R11593 GND.n1811 GND.n1798 9.3005
R11594 GND.n6044 GND.n1812 9.3005
R11595 GND.n6043 GND.n1813 9.3005
R11596 GND.n6042 GND.n1814 9.3005
R11597 GND.n1828 GND.n1815 9.3005
R11598 GND.n6030 GND.n1829 9.3005
R11599 GND.n6029 GND.n1830 9.3005
R11600 GND.n6028 GND.n1831 9.3005
R11601 GND.n1846 GND.n1832 9.3005
R11602 GND.n6016 GND.n1847 9.3005
R11603 GND.n6015 GND.n1848 9.3005
R11604 GND.n6014 GND.n1849 9.3005
R11605 GND.n1916 GND.n1850 9.3005
R11606 GND.n5803 GND.n1917 9.3005
R11607 GND.n5802 GND.n1918 9.3005
R11608 GND.n5801 GND.n1919 9.3005
R11609 GND.n1942 GND.n1920 9.3005
R11610 GND.n1943 GND.n1941 9.3005
R11611 GND.n5789 GND.n1944 9.3005
R11612 GND.n5788 GND.n1945 9.3005
R11613 GND.n5787 GND.n1946 9.3005
R11614 GND.n1969 GND.n1947 9.3005
R11615 GND.n1970 GND.n1968 9.3005
R11616 GND.n5775 GND.n1971 9.3005
R11617 GND.n5774 GND.n1972 9.3005
R11618 GND.n5773 GND.n1973 9.3005
R11619 GND.n1996 GND.n1974 9.3005
R11620 GND.n1997 GND.n1995 9.3005
R11621 GND.n5761 GND.n1998 9.3005
R11622 GND.n5760 GND.n1999 9.3005
R11623 GND.n5759 GND.n2000 9.3005
R11624 GND.n2022 GND.n2001 9.3005
R11625 GND.n2023 GND.n2021 9.3005
R11626 GND.n5747 GND.n2024 9.3005
R11627 GND.n5746 GND.n2025 9.3005
R11628 GND.n5745 GND.n2026 9.3005
R11629 GND.n2049 GND.n2027 9.3005
R11630 GND.n2050 GND.n2048 9.3005
R11631 GND.n5733 GND.n2051 9.3005
R11632 GND.n5732 GND.n2052 9.3005
R11633 GND.n5731 GND.n2053 9.3005
R11634 GND.n2076 GND.n2054 9.3005
R11635 GND.n2077 GND.n2075 9.3005
R11636 GND.n5719 GND.n2078 9.3005
R11637 GND.n5718 GND.n2079 9.3005
R11638 GND.n5717 GND.n2080 9.3005
R11639 GND.n2103 GND.n2081 9.3005
R11640 GND.n2104 GND.n2102 9.3005
R11641 GND.n5705 GND.n2105 9.3005
R11642 GND.n5704 GND.n2106 9.3005
R11643 GND.n5703 GND.n2107 9.3005
R11644 GND.n2130 GND.n2108 9.3005
R11645 GND.n2131 GND.n2129 9.3005
R11646 GND.n5691 GND.n2132 9.3005
R11647 GND.n5690 GND.n2133 9.3005
R11648 GND.n5689 GND.n2134 9.3005
R11649 GND.n2157 GND.n2135 9.3005
R11650 GND.n2158 GND.n2156 9.3005
R11651 GND.n5677 GND.n2159 9.3005
R11652 GND.n5676 GND.n2160 9.3005
R11653 GND.n5675 GND.n2161 9.3005
R11654 GND.n2183 GND.n2162 9.3005
R11655 GND.n2184 GND.n2182 9.3005
R11656 GND.n5663 GND.n2185 9.3005
R11657 GND.n5662 GND.n2186 9.3005
R11658 GND.n5661 GND.n2187 9.3005
R11659 GND.n2210 GND.n2188 9.3005
R11660 GND.n2211 GND.n2209 9.3005
R11661 GND.n5649 GND.n2212 9.3005
R11662 GND.n5648 GND.n2213 9.3005
R11663 GND.n5647 GND.n2214 9.3005
R11664 GND.n2590 GND.n2215 9.3005
R11665 GND.n2593 GND.n2592 9.3005
R11666 GND.n2594 GND.n2589 9.3005
R11667 GND.n2596 GND.n2595 9.3005
R11668 GND.n2586 GND.n2585 9.3005
R11669 GND.n2601 GND.n2600 9.3005
R11670 GND.n2602 GND.n2584 9.3005
R11671 GND.n2604 GND.n2603 9.3005
R11672 GND.n2582 GND.n2581 9.3005
R11673 GND.n2609 GND.n2608 9.3005
R11674 GND.n2610 GND.n2580 9.3005
R11675 GND.n2655 GND.n2611 9.3005
R11676 GND.n2654 GND.n2612 9.3005
R11677 GND.n2653 GND.n2613 9.3005
R11678 GND.n2616 GND.n2614 9.3005
R11679 GND.n2649 GND.n2617 9.3005
R11680 GND.n2648 GND.n2618 9.3005
R11681 GND.n2647 GND.n2619 9.3005
R11682 GND.n2622 GND.n2620 9.3005
R11683 GND.n2643 GND.n2623 9.3005
R11684 GND.n2642 GND.n2624 9.3005
R11685 GND.n2641 GND.n2625 9.3005
R11686 GND.n2628 GND.n2626 9.3005
R11687 GND.n2637 GND.n2629 9.3005
R11688 GND.n5200 GND.n5148 9.3005
R11689 GND.n5199 GND.n5149 9.3005
R11690 GND.n5198 GND.n5150 9.3005
R11691 GND.n5153 GND.n5151 9.3005
R11692 GND.n5194 GND.n5154 9.3005
R11693 GND.n5193 GND.n5155 9.3005
R11694 GND.n5192 GND.n5156 9.3005
R11695 GND.n5159 GND.n5157 9.3005
R11696 GND.n5188 GND.n5160 9.3005
R11697 GND.n5187 GND.n5161 9.3005
R11698 GND.n5186 GND.n5162 9.3005
R11699 GND.n5165 GND.n5163 9.3005
R11700 GND.n5182 GND.n5166 9.3005
R11701 GND.n5181 GND.n5167 9.3005
R11702 GND.n5180 GND.n5168 9.3005
R11703 GND.n5171 GND.n5169 9.3005
R11704 GND.n5176 GND.n5172 9.3005
R11705 GND.n5175 GND.n5174 9.3005
R11706 GND.n5173 GND.n294 9.3005
R11707 GND.n7872 GND.n295 9.3005
R11708 GND.n7871 GND.n296 9.3005
R11709 GND.n7870 GND.n297 9.3005
R11710 GND.n302 GND.n298 9.3005
R11711 GND.n7864 GND.n303 9.3005
R11712 GND.n7863 GND.n304 9.3005
R11713 GND.n7862 GND.n305 9.3005
R11714 GND.n310 GND.n306 9.3005
R11715 GND.n7856 GND.n311 9.3005
R11716 GND.n7855 GND.n312 9.3005
R11717 GND.n7854 GND.n313 9.3005
R11718 GND.n318 GND.n314 9.3005
R11719 GND.n7848 GND.n319 9.3005
R11720 GND.n7847 GND.n320 9.3005
R11721 GND.n7846 GND.n321 9.3005
R11722 GND.n326 GND.n322 9.3005
R11723 GND.n7840 GND.n327 9.3005
R11724 GND.n7839 GND.n328 9.3005
R11725 GND.n7838 GND.n329 9.3005
R11726 GND.n334 GND.n330 9.3005
R11727 GND.n7832 GND.n335 9.3005
R11728 GND.n7831 GND.n336 9.3005
R11729 GND.n7830 GND.n337 9.3005
R11730 GND.n342 GND.n338 9.3005
R11731 GND.n7824 GND.n343 9.3005
R11732 GND.n7823 GND.n344 9.3005
R11733 GND.n7822 GND.n345 9.3005
R11734 GND.n350 GND.n346 9.3005
R11735 GND.n7816 GND.n351 9.3005
R11736 GND.n7815 GND.n352 9.3005
R11737 GND.n7814 GND.n353 9.3005
R11738 GND.n358 GND.n354 9.3005
R11739 GND.n7808 GND.n359 9.3005
R11740 GND.n7807 GND.n360 9.3005
R11741 GND.n7806 GND.n361 9.3005
R11742 GND.n366 GND.n362 9.3005
R11743 GND.n7800 GND.n367 9.3005
R11744 GND.n7799 GND.n368 9.3005
R11745 GND.n7798 GND.n369 9.3005
R11746 GND.n374 GND.n370 9.3005
R11747 GND.n7792 GND.n375 9.3005
R11748 GND.n7791 GND.n376 9.3005
R11749 GND.n7790 GND.n377 9.3005
R11750 GND.n382 GND.n378 9.3005
R11751 GND.n7784 GND.n383 9.3005
R11752 GND.n7783 GND.n384 9.3005
R11753 GND.n7782 GND.n385 9.3005
R11754 GND.n390 GND.n386 9.3005
R11755 GND.n7776 GND.n391 9.3005
R11756 GND.n7775 GND.n392 9.3005
R11757 GND.n7774 GND.n393 9.3005
R11758 GND.n398 GND.n394 9.3005
R11759 GND.n7768 GND.n399 9.3005
R11760 GND.n7767 GND.n400 9.3005
R11761 GND.n7766 GND.n401 9.3005
R11762 GND.n406 GND.n402 9.3005
R11763 GND.n7760 GND.n407 9.3005
R11764 GND.n7759 GND.n408 9.3005
R11765 GND.n7758 GND.n409 9.3005
R11766 GND.n414 GND.n410 9.3005
R11767 GND.n7752 GND.n7751 9.3005
R11768 GND.n3760 GND.n3759 9.3005
R11769 GND.n3758 GND.n3540 9.3005
R11770 GND.n3757 GND.n3756 9.3005
R11771 GND.n3753 GND.n3542 9.3005
R11772 GND.n3750 GND.n3749 9.3005
R11773 GND.n3748 GND.n3543 9.3005
R11774 GND.n3747 GND.n3746 9.3005
R11775 GND.n3743 GND.n3544 9.3005
R11776 GND.n3740 GND.n3739 9.3005
R11777 GND.n3738 GND.n3545 9.3005
R11778 GND.n3737 GND.n3736 9.3005
R11779 GND.n3733 GND.n3546 9.3005
R11780 GND.n3730 GND.n3729 9.3005
R11781 GND.n3728 GND.n3547 9.3005
R11782 GND.n3727 GND.n3726 9.3005
R11783 GND.n3723 GND.n3548 9.3005
R11784 GND.n3720 GND.n3719 9.3005
R11785 GND.n3718 GND.n3549 9.3005
R11786 GND.n3717 GND.n3716 9.3005
R11787 GND.n3710 GND.n3550 9.3005
R11788 GND.n3707 GND.n3706 9.3005
R11789 GND.n3705 GND.n3551 9.3005
R11790 GND.n3704 GND.n3703 9.3005
R11791 GND.n3700 GND.n3552 9.3005
R11792 GND.n3697 GND.n3696 9.3005
R11793 GND.n3695 GND.n3553 9.3005
R11794 GND.n3694 GND.n3693 9.3005
R11795 GND.n3690 GND.n3554 9.3005
R11796 GND.n3687 GND.n3686 9.3005
R11797 GND.n3685 GND.n3555 9.3005
R11798 GND.n3684 GND.n3683 9.3005
R11799 GND.n3680 GND.n3556 9.3005
R11800 GND.n3677 GND.n3676 9.3005
R11801 GND.n3675 GND.n3557 9.3005
R11802 GND.n3674 GND.n3673 9.3005
R11803 GND.n3670 GND.n3558 9.3005
R11804 GND.n3667 GND.n3664 9.3005
R11805 GND.n3663 GND.n3559 9.3005
R11806 GND.n3662 GND.n3661 9.3005
R11807 GND.n3658 GND.n3560 9.3005
R11808 GND.n3655 GND.n3654 9.3005
R11809 GND.n3653 GND.n3561 9.3005
R11810 GND.n3652 GND.n3651 9.3005
R11811 GND.n3648 GND.n3562 9.3005
R11812 GND.n3645 GND.n3644 9.3005
R11813 GND.n3643 GND.n3563 9.3005
R11814 GND.n3642 GND.n3641 9.3005
R11815 GND.n3638 GND.n3564 9.3005
R11816 GND.n3635 GND.n3634 9.3005
R11817 GND.n3633 GND.n3565 9.3005
R11818 GND.n3632 GND.n3631 9.3005
R11819 GND.n3628 GND.n3566 9.3005
R11820 GND.n3625 GND.n3624 9.3005
R11821 GND.n3623 GND.n3567 9.3005
R11822 GND.n3622 GND.n3621 9.3005
R11823 GND.n3613 GND.n3612 9.3005
R11824 GND.n3611 GND.n3569 9.3005
R11825 GND.n3610 GND.n3609 9.3005
R11826 GND.n3606 GND.n3570 9.3005
R11827 GND.n3603 GND.n3602 9.3005
R11828 GND.n3601 GND.n3571 9.3005
R11829 GND.n3600 GND.n3599 9.3005
R11830 GND.n3596 GND.n3572 9.3005
R11831 GND.n3593 GND.n3592 9.3005
R11832 GND.n3591 GND.n3573 9.3005
R11833 GND.n3590 GND.n3589 9.3005
R11834 GND.n3586 GND.n3574 9.3005
R11835 GND.n3583 GND.n3582 9.3005
R11836 GND.n3581 GND.n3575 9.3005
R11837 GND.n3580 GND.n3579 9.3005
R11838 GND.n3576 GND.n3523 9.3005
R11839 GND.n3618 GND.n3568 9.3005
R11840 GND.n3761 GND.n3536 9.3005
R11841 GND.n3763 GND.n3762 9.3005
R11842 GND.n3783 GND.n3522 9.3005
R11843 GND.n3787 GND.n3784 9.3005
R11844 GND.n3786 GND.n3785 9.3005
R11845 GND.n3495 GND.n3494 9.3005
R11846 GND.n3819 GND.n3818 9.3005
R11847 GND.n3820 GND.n3493 9.3005
R11848 GND.n3824 GND.n3821 9.3005
R11849 GND.n3823 GND.n3822 9.3005
R11850 GND.n3466 GND.n3465 9.3005
R11851 GND.n3856 GND.n3855 9.3005
R11852 GND.n3857 GND.n3464 9.3005
R11853 GND.n3861 GND.n3858 9.3005
R11854 GND.n3860 GND.n3859 9.3005
R11855 GND.n3437 GND.n3436 9.3005
R11856 GND.n3896 GND.n3895 9.3005
R11857 GND.n3897 GND.n3435 9.3005
R11858 GND.n3900 GND.n3899 9.3005
R11859 GND.n3898 GND.n3414 9.3005
R11860 GND.n4016 GND.n4015 9.3005
R11861 GND.n4017 GND.n3381 9.3005
R11862 GND.n4021 GND.n4018 9.3005
R11863 GND.n4020 GND.n4019 9.3005
R11864 GND.n3354 GND.n3353 9.3005
R11865 GND.n4053 GND.n4052 9.3005
R11866 GND.n4054 GND.n3352 9.3005
R11867 GND.n4058 GND.n4055 9.3005
R11868 GND.n4057 GND.n4056 9.3005
R11869 GND.n3324 GND.n3323 9.3005
R11870 GND.n4090 GND.n4089 9.3005
R11871 GND.n4091 GND.n3322 9.3005
R11872 GND.n4095 GND.n4092 9.3005
R11873 GND.n4094 GND.n4093 9.3005
R11874 GND.n3297 GND.n3296 9.3005
R11875 GND.n4145 GND.n4144 9.3005
R11876 GND.n4146 GND.n3295 9.3005
R11877 GND.n4149 GND.n4147 9.3005
R11878 GND.n4148 GND.n1516 9.3005
R11879 GND.n3782 GND.n3781 9.3005
R11880 GND.n3983 GND.n3382 9.3005
R11881 GND.n3383 GND.n3382 9.3005
R11882 GND.n6497 GND.n1212 9.3005
R11883 GND.n1217 GND.n1213 9.3005
R11884 GND.n6491 GND.n1218 9.3005
R11885 GND.n6490 GND.n1219 9.3005
R11886 GND.n6489 GND.n1220 9.3005
R11887 GND.n1225 GND.n1221 9.3005
R11888 GND.n6483 GND.n1226 9.3005
R11889 GND.n6482 GND.n1227 9.3005
R11890 GND.n6481 GND.n1228 9.3005
R11891 GND.n1233 GND.n1229 9.3005
R11892 GND.n6475 GND.n1234 9.3005
R11893 GND.n6474 GND.n1235 9.3005
R11894 GND.n6473 GND.n1236 9.3005
R11895 GND.n1241 GND.n1237 9.3005
R11896 GND.n6467 GND.n1242 9.3005
R11897 GND.n6466 GND.n1243 9.3005
R11898 GND.n6465 GND.n1244 9.3005
R11899 GND.n1249 GND.n1245 9.3005
R11900 GND.n6459 GND.n1250 9.3005
R11901 GND.n6458 GND.n1251 9.3005
R11902 GND.n6457 GND.n1252 9.3005
R11903 GND.n1257 GND.n1253 9.3005
R11904 GND.n6451 GND.n1258 9.3005
R11905 GND.n6450 GND.n1259 9.3005
R11906 GND.n6449 GND.n1260 9.3005
R11907 GND.n1265 GND.n1261 9.3005
R11908 GND.n6443 GND.n1266 9.3005
R11909 GND.n6442 GND.n1267 9.3005
R11910 GND.n6441 GND.n1268 9.3005
R11911 GND.n1273 GND.n1269 9.3005
R11912 GND.n6435 GND.n1274 9.3005
R11913 GND.n6434 GND.n1275 9.3005
R11914 GND.n6433 GND.n1276 9.3005
R11915 GND.n1281 GND.n1277 9.3005
R11916 GND.n6427 GND.n1282 9.3005
R11917 GND.n6426 GND.n1283 9.3005
R11918 GND.n6425 GND.n1284 9.3005
R11919 GND.n1289 GND.n1285 9.3005
R11920 GND.n6419 GND.n1290 9.3005
R11921 GND.n6418 GND.n1291 9.3005
R11922 GND.n6417 GND.n1292 9.3005
R11923 GND.n1297 GND.n1293 9.3005
R11924 GND.n6411 GND.n1298 9.3005
R11925 GND.n6410 GND.n1299 9.3005
R11926 GND.n6409 GND.n1300 9.3005
R11927 GND.n1305 GND.n1301 9.3005
R11928 GND.n6403 GND.n1306 9.3005
R11929 GND.n6402 GND.n1307 9.3005
R11930 GND.n6401 GND.n1308 9.3005
R11931 GND.n1313 GND.n1309 9.3005
R11932 GND.n6395 GND.n1314 9.3005
R11933 GND.n6394 GND.n1315 9.3005
R11934 GND.n6393 GND.n1316 9.3005
R11935 GND.n1321 GND.n1317 9.3005
R11936 GND.n6387 GND.n1322 9.3005
R11937 GND.n6386 GND.n1323 9.3005
R11938 GND.n6385 GND.n1324 9.3005
R11939 GND.n3527 GND.n1325 9.3005
R11940 GND.n3528 GND.n3526 9.3005
R11941 GND.n3530 GND.n3529 9.3005
R11942 GND.n3514 GND.n3513 9.3005
R11943 GND.n3793 GND.n3792 9.3005
R11944 GND.n3794 GND.n3512 9.3005
R11945 GND.n3798 GND.n3795 9.3005
R11946 GND.n3797 GND.n3796 9.3005
R11947 GND.n3484 GND.n3483 9.3005
R11948 GND.n3830 GND.n3829 9.3005
R11949 GND.n3831 GND.n3482 9.3005
R11950 GND.n3835 GND.n3832 9.3005
R11951 GND.n3834 GND.n3833 9.3005
R11952 GND.n3455 GND.n3454 9.3005
R11953 GND.n3867 GND.n3866 9.3005
R11954 GND.n3868 GND.n3453 9.3005
R11955 GND.n3878 GND.n3869 9.3005
R11956 GND.n3877 GND.n3870 9.3005
R11957 GND.n3876 GND.n3871 9.3005
R11958 GND.n3873 GND.n3872 9.3005
R11959 GND.n3403 GND.n3402 9.3005
R11960 GND.n3992 GND.n3991 9.3005
R11961 GND.n6499 GND.n6498 9.3005
R11962 GND.n1211 GND.n1207 9.3005
R11963 GND.n6507 GND.n1206 9.3005
R11964 GND.n6508 GND.n1205 9.3005
R11965 GND.n6509 GND.n1204 9.3005
R11966 GND.n1203 GND.n1199 9.3005
R11967 GND.n6515 GND.n1198 9.3005
R11968 GND.n6516 GND.n1197 9.3005
R11969 GND.n6517 GND.n1196 9.3005
R11970 GND.n1195 GND.n1191 9.3005
R11971 GND.n6523 GND.n1190 9.3005
R11972 GND.n6524 GND.n1189 9.3005
R11973 GND.n6525 GND.n1188 9.3005
R11974 GND.n1187 GND.n1183 9.3005
R11975 GND.n6531 GND.n1182 9.3005
R11976 GND.n6532 GND.n1181 9.3005
R11977 GND.n6533 GND.n1180 9.3005
R11978 GND.n1179 GND.n1175 9.3005
R11979 GND.n6539 GND.n1174 9.3005
R11980 GND.n6540 GND.n1173 9.3005
R11981 GND.n6541 GND.n1172 9.3005
R11982 GND.n1171 GND.n1167 9.3005
R11983 GND.n6547 GND.n1166 9.3005
R11984 GND.n6548 GND.n1165 9.3005
R11985 GND.n6549 GND.n1164 9.3005
R11986 GND.n1163 GND.n1159 9.3005
R11987 GND.n6555 GND.n1158 9.3005
R11988 GND.n6556 GND.n1157 9.3005
R11989 GND.n6557 GND.n1156 9.3005
R11990 GND.n1155 GND.n1151 9.3005
R11991 GND.n6563 GND.n1150 9.3005
R11992 GND.n6564 GND.n1149 9.3005
R11993 GND.n6565 GND.n1148 9.3005
R11994 GND.n1147 GND.n1143 9.3005
R11995 GND.n6571 GND.n1142 9.3005
R11996 GND.n6572 GND.n1141 9.3005
R11997 GND.n6573 GND.n1140 9.3005
R11998 GND.n1139 GND.n1135 9.3005
R11999 GND.n6579 GND.n1134 9.3005
R12000 GND.n6580 GND.n1133 9.3005
R12001 GND.n6581 GND.n1132 9.3005
R12002 GND.n1131 GND.n1127 9.3005
R12003 GND.n6587 GND.n1126 9.3005
R12004 GND.n6588 GND.n1125 9.3005
R12005 GND.n6589 GND.n1124 9.3005
R12006 GND.n1123 GND.n1119 9.3005
R12007 GND.n6595 GND.n1118 9.3005
R12008 GND.n6596 GND.n1117 9.3005
R12009 GND.n6597 GND.n1116 9.3005
R12010 GND.n1115 GND.n1111 9.3005
R12011 GND.n6603 GND.n1110 9.3005
R12012 GND.n6604 GND.n1109 9.3005
R12013 GND.n6605 GND.n1108 9.3005
R12014 GND.n1107 GND.n1103 9.3005
R12015 GND.n6611 GND.n1102 9.3005
R12016 GND.n6612 GND.n1101 9.3005
R12017 GND.n6613 GND.n1100 9.3005
R12018 GND.n1099 GND.n1095 9.3005
R12019 GND.n6619 GND.n1094 9.3005
R12020 GND.n6620 GND.n1093 9.3005
R12021 GND.n6621 GND.n1092 9.3005
R12022 GND.n1088 GND.n1087 9.3005
R12023 GND.n6628 GND.n6627 9.3005
R12024 GND.n6501 GND.n6500 9.3005
R12025 GND.n6312 GND.n6311 9.3005
R12026 GND.n6310 GND.n1429 9.3005
R12027 GND.n6309 GND.n6308 9.3005
R12028 GND.n6307 GND.n1433 9.3005
R12029 GND.n6306 GND.n6305 9.3005
R12030 GND.n6304 GND.n1434 9.3005
R12031 GND.n6303 GND.n6302 9.3005
R12032 GND.n6301 GND.n1438 9.3005
R12033 GND.n6300 GND.n6299 9.3005
R12034 GND.n6298 GND.n1439 9.3005
R12035 GND.n6297 GND.n6296 9.3005
R12036 GND.n6295 GND.n1443 9.3005
R12037 GND.n6294 GND.n6293 9.3005
R12038 GND.n6292 GND.n1444 9.3005
R12039 GND.n6291 GND.n6290 9.3005
R12040 GND.n6289 GND.n1448 9.3005
R12041 GND.n6288 GND.n6287 9.3005
R12042 GND.n6286 GND.n1449 9.3005
R12043 GND.n6285 GND.n6284 9.3005
R12044 GND.n6283 GND.n1453 9.3005
R12045 GND.n6282 GND.n6281 9.3005
R12046 GND.n6280 GND.n1454 9.3005
R12047 GND.n6279 GND.n6278 9.3005
R12048 GND.n6277 GND.n1458 9.3005
R12049 GND.n1462 GND.n1459 9.3005
R12050 GND.n6276 GND.n6275 9.3005
R12051 GND.n3162 GND.n3161 9.3005
R12052 GND.n3160 GND.n3159 9.3005
R12053 GND.n3084 GND.n3083 9.3005
R12054 GND.n3154 GND.n3153 9.3005
R12055 GND.n3152 GND.n3151 9.3005
R12056 GND.n3092 GND.n3091 9.3005
R12057 GND.n3146 GND.n3145 9.3005
R12058 GND.n3144 GND.n3143 9.3005
R12059 GND.n3104 GND.n3103 9.3005
R12060 GND.n3135 GND.n3134 9.3005
R12061 GND.n3133 GND.n3132 9.3005
R12062 GND.n3111 GND.n3110 9.3005
R12063 GND.n3127 GND.n3126 9.3005
R12064 GND.n3125 GND.n3115 9.3005
R12065 GND.n3124 GND.n3123 9.3005
R12066 GND.n3079 GND.n3072 9.3005
R12067 GND.n3131 GND.n3130 9.3005
R12068 GND.n3107 GND.n3106 9.3005
R12069 GND.n3140 GND.n3136 9.3005
R12070 GND.n3142 GND.n3141 9.3005
R12071 GND.n3098 GND.n3097 9.3005
R12072 GND.n3148 GND.n3147 9.3005
R12073 GND.n3150 GND.n3149 9.3005
R12074 GND.n3088 GND.n3087 9.3005
R12075 GND.n3156 GND.n3155 9.3005
R12076 GND.n3158 GND.n3157 9.3005
R12077 GND.n3078 GND.n3077 9.3005
R12078 GND.n3164 GND.n3163 9.3005
R12079 GND.n3166 GND.n3165 9.3005
R12080 GND.n3167 GND.n3071 9.3005
R12081 GND.n3129 GND.n3128 9.3005
R12082 GND.n6222 GND.n1566 9.3005
R12083 GND.n6223 GND.n1562 9.3005
R12084 GND.n6225 GND.n6224 9.3005
R12085 GND.n6226 GND.n1561 9.3005
R12086 GND.n6228 GND.n6227 9.3005
R12087 GND.n6229 GND.n1556 9.3005
R12088 GND.n6231 GND.n6230 9.3005
R12089 GND.n6232 GND.n1555 9.3005
R12090 GND.n6234 GND.n6233 9.3005
R12091 GND.n6235 GND.n1550 9.3005
R12092 GND.n6237 GND.n6236 9.3005
R12093 GND.n6238 GND.n1549 9.3005
R12094 GND.n6240 GND.n6239 9.3005
R12095 GND.n6241 GND.n1544 9.3005
R12096 GND.n6243 GND.n6242 9.3005
R12097 GND.n6244 GND.n1543 9.3005
R12098 GND.n6246 GND.n6245 9.3005
R12099 GND.n6247 GND.n1540 9.3005
R12100 GND.n6248 GND.n1535 9.3005
R12101 GND.n6250 GND.n6249 9.3005
R12102 GND.n6251 GND.n1534 9.3005
R12103 GND.n6253 GND.n6252 9.3005
R12104 GND.n6254 GND.n1529 9.3005
R12105 GND.n6256 GND.n6255 9.3005
R12106 GND.n6257 GND.n1528 9.3005
R12107 GND.n6259 GND.n6258 9.3005
R12108 GND.n6260 GND.n1523 9.3005
R12109 GND.n6262 GND.n6261 9.3005
R12110 GND.n6263 GND.n1522 9.3005
R12111 GND.n6265 GND.n6264 9.3005
R12112 GND.n6266 GND.n1517 9.3005
R12113 GND.n6268 GND.n6267 9.3005
R12114 GND.n6269 GND.n1515 9.3005
R12115 GND.n6271 GND.n6270 9.3005
R12116 GND.n3211 GND.n1568 9.3005
R12117 GND.n3213 GND.n3212 9.3005
R12118 GND.n3217 GND.n3216 9.3005
R12119 GND.n3218 GND.n3208 9.3005
R12120 GND.n3220 GND.n3219 9.3005
R12121 GND.n3221 GND.n3207 9.3005
R12122 GND.n3225 GND.n3224 9.3005
R12123 GND.n3226 GND.n3204 9.3005
R12124 GND.n3228 GND.n3227 9.3005
R12125 GND.n3229 GND.n3203 9.3005
R12126 GND.n3233 GND.n3232 9.3005
R12127 GND.n3234 GND.n3200 9.3005
R12128 GND.n3236 GND.n3235 9.3005
R12129 GND.n3237 GND.n3199 9.3005
R12130 GND.n3241 GND.n3240 9.3005
R12131 GND.n3242 GND.n3196 9.3005
R12132 GND.n3244 GND.n3243 9.3005
R12133 GND.n3245 GND.n3192 9.3005
R12134 GND.n3249 GND.n3248 9.3005
R12135 GND.n3250 GND.n3189 9.3005
R12136 GND.n3252 GND.n3251 9.3005
R12137 GND.n3253 GND.n3188 9.3005
R12138 GND.n3257 GND.n3256 9.3005
R12139 GND.n3258 GND.n3185 9.3005
R12140 GND.n3260 GND.n3259 9.3005
R12141 GND.n3261 GND.n3184 9.3005
R12142 GND.n3265 GND.n3264 9.3005
R12143 GND.n3266 GND.n3181 9.3005
R12144 GND.n3268 GND.n3267 9.3005
R12145 GND.n3269 GND.n3180 9.3005
R12146 GND.n3273 GND.n3272 9.3005
R12147 GND.n3274 GND.n3177 9.3005
R12148 GND.n3276 GND.n3275 9.3005
R12149 GND.n3277 GND.n3176 9.3005
R12150 GND.n3281 GND.n3280 9.3005
R12151 GND.n3282 GND.n3173 9.3005
R12152 GND.n3286 GND.n3283 9.3005
R12153 GND.n3287 GND.n3168 9.3005
R12154 GND.n3774 GND.n3767 9.3005
R12155 GND.n3773 GND.n3768 9.3005
R12156 GND.n3771 GND.n3770 9.3005
R12157 GND.n3504 GND.n3502 9.3005
R12158 GND.n3814 GND.n3813 9.3005
R12159 GND.n3505 GND.n3503 9.3005
R12160 GND.n3809 GND.n3805 9.3005
R12161 GND.n3808 GND.n3807 9.3005
R12162 GND.n3475 GND.n3473 9.3005
R12163 GND.n3851 GND.n3850 9.3005
R12164 GND.n3476 GND.n3474 9.3005
R12165 GND.n3846 GND.n3842 9.3005
R12166 GND.n3845 GND.n3844 9.3005
R12167 GND.n3446 GND.n3444 9.3005
R12168 GND.n3891 GND.n3890 9.3005
R12169 GND.n3447 GND.n3445 9.3005
R12170 GND.n3886 GND.n3428 9.3005
R12171 GND.n3905 GND.n3427 9.3005
R12172 GND.n3907 GND.n3906 9.3005
R12173 GND.n3424 GND.n3422 9.3005
R12174 GND.n3979 GND.n3978 9.3005
R12175 GND.n3425 GND.n3423 9.3005
R12176 GND.n3974 GND.n3915 9.3005
R12177 GND.n3973 GND.n3916 9.3005
R12178 GND.n3972 GND.n3917 9.3005
R12179 GND.n3925 GND.n3918 9.3005
R12180 GND.n3927 GND.n3926 9.3005
R12181 GND.n3391 GND.n3389 9.3005
R12182 GND.n4011 GND.n4010 9.3005
R12183 GND.n3392 GND.n3390 9.3005
R12184 GND.n4006 GND.n4002 9.3005
R12185 GND.n4005 GND.n4004 9.3005
R12186 GND.n3363 GND.n3361 9.3005
R12187 GND.n4048 GND.n4047 9.3005
R12188 GND.n3364 GND.n3362 9.3005
R12189 GND.n4043 GND.n4039 9.3005
R12190 GND.n4042 GND.n4041 9.3005
R12191 GND.n3334 GND.n3332 9.3005
R12192 GND.n4085 GND.n4084 9.3005
R12193 GND.n3335 GND.n3333 9.3005
R12194 GND.n4080 GND.n4076 9.3005
R12195 GND.n4079 GND.n4078 9.3005
R12196 GND.n3305 GND.n3303 9.3005
R12197 GND.n4140 GND.n4139 9.3005
R12198 GND.n3306 GND.n3304 9.3005
R12199 GND.n3292 GND.n3169 9.3005
R12200 GND.n4157 GND.n3170 9.3005
R12201 GND.n3775 GND.n3765 9.3005
R12202 GND.n3774 GND.n3535 9.3005
R12203 GND.n3773 GND.n3772 9.3005
R12204 GND.n3771 GND.n3506 9.3005
R12205 GND.n3803 GND.n3504 9.3005
R12206 GND.n3813 GND.n3812 9.3005
R12207 GND.n3811 GND.n3505 9.3005
R12208 GND.n3810 GND.n3809 9.3005
R12209 GND.n3808 GND.n3477 9.3005
R12210 GND.n3840 GND.n3475 9.3005
R12211 GND.n3850 GND.n3849 9.3005
R12212 GND.n3848 GND.n3476 9.3005
R12213 GND.n3847 GND.n3846 9.3005
R12214 GND.n3845 GND.n3448 9.3005
R12215 GND.n3883 GND.n3446 9.3005
R12216 GND.n3890 GND.n3889 9.3005
R12217 GND.n3888 GND.n3447 9.3005
R12218 GND.n3887 GND.n3886 9.3005
R12219 GND.n3427 GND.n3426 9.3005
R12220 GND.n3908 GND.n3907 9.3005
R12221 GND.n3911 GND.n3424 9.3005
R12222 GND.n3978 GND.n3977 9.3005
R12223 GND.n3976 GND.n3425 9.3005
R12224 GND.n3975 GND.n3974 9.3005
R12225 GND.n3973 GND.n3914 9.3005
R12226 GND.n3972 GND.n3971 9.3005
R12227 GND.n3970 GND.n3918 9.3005
R12228 GND.n3926 GND.n3393 9.3005
R12229 GND.n4000 GND.n3391 9.3005
R12230 GND.n4010 GND.n4009 9.3005
R12231 GND.n4008 GND.n3392 9.3005
R12232 GND.n4007 GND.n4006 9.3005
R12233 GND.n4005 GND.n3365 9.3005
R12234 GND.n4037 GND.n3363 9.3005
R12235 GND.n4047 GND.n4046 9.3005
R12236 GND.n4045 GND.n3364 9.3005
R12237 GND.n4044 GND.n4043 9.3005
R12238 GND.n4042 GND.n3336 9.3005
R12239 GND.n4074 GND.n3334 9.3005
R12240 GND.n4084 GND.n4083 9.3005
R12241 GND.n4082 GND.n3335 9.3005
R12242 GND.n4081 GND.n4080 9.3005
R12243 GND.n4079 GND.n3307 9.3005
R12244 GND.n4134 GND.n3305 9.3005
R12245 GND.n4139 GND.n4138 9.3005
R12246 GND.n4137 GND.n3306 9.3005
R12247 GND.n3171 GND.n3169 9.3005
R12248 GND.n4157 GND.n4156 9.3005
R12249 GND.n3776 GND.n3775 9.3005
R12250 GND.n6357 GND.n6356 9.3005
R12251 GND.n6358 GND.n1395 9.3005
R12252 GND.n6360 GND.n6359 9.3005
R12253 GND.n6361 GND.n1390 9.3005
R12254 GND.n6363 GND.n6362 9.3005
R12255 GND.n6364 GND.n1389 9.3005
R12256 GND.n6366 GND.n6365 9.3005
R12257 GND.n6367 GND.n1384 9.3005
R12258 GND.n6369 GND.n6368 9.3005
R12259 GND.n6370 GND.n1383 9.3005
R12260 GND.n6372 GND.n6371 9.3005
R12261 GND.n6373 GND.n1378 9.3005
R12262 GND.n6375 GND.n6374 9.3005
R12263 GND.n6376 GND.n1377 9.3005
R12264 GND.n6378 GND.n6377 9.3005
R12265 GND.n6379 GND.n1376 9.3005
R12266 GND.n6355 GND.n1396 9.3005
R12267 GND.n6351 GND.n6350 9.3005
R12268 GND.n6347 GND.n1399 9.3005
R12269 GND.n6346 GND.n6345 9.3005
R12270 GND.n6344 GND.n1403 9.3005
R12271 GND.n6343 GND.n6342 9.3005
R12272 GND.n6341 GND.n1404 9.3005
R12273 GND.n6340 GND.n6339 9.3005
R12274 GND.n6338 GND.n1408 9.3005
R12275 GND.n6337 GND.n6336 9.3005
R12276 GND.n6335 GND.n1409 9.3005
R12277 GND.n6334 GND.n6333 9.3005
R12278 GND.n6332 GND.n1413 9.3005
R12279 GND.n6331 GND.n6330 9.3005
R12280 GND.n6329 GND.n1414 9.3005
R12281 GND.n6328 GND.n6327 9.3005
R12282 GND.n6326 GND.n1418 9.3005
R12283 GND.n6325 GND.n6324 9.3005
R12284 GND.n6323 GND.n1419 9.3005
R12285 GND.n6322 GND.n6321 9.3005
R12286 GND.n6320 GND.n1423 9.3005
R12287 GND.n6319 GND.n6318 9.3005
R12288 GND.n6317 GND.n1424 9.3005
R12289 GND.n6316 GND.n6315 9.3005
R12290 GND.n6314 GND.n1428 9.3005
R12291 GND.n6349 GND.n6348 9.3005
R12292 GND.n3499 GND.t63 9.22295
R12293 GND.t67 GND.n124 9.22295
R12294 GND.n3287 GND.n3286 9.11565
R12295 GND.n5444 GND.n2398 9.11565
R12296 GND.n7882 GND.n283 9.11565
R12297 GND.n3762 GND.n3761 9.11565
R12298 GND.n4666 GND.t151 8.92545
R12299 GND.n4672 GND.n1669 8.92545
R12300 GND.n4755 GND.n2755 8.92545
R12301 GND.n2741 GND.n1774 8.92545
R12302 GND.n6040 GND.t88 8.92545
R12303 GND.n5939 GND.n1852 8.92545
R12304 GND.n6222 GND.n6220 8.92171
R12305 GND.n5522 GND.n5521 8.92171
R12306 GND.n6273 GND.n1494 8.62795
R12307 GND.n5588 GND.n2268 8.62795
R12308 GND.n2760 GND.n2759 8.33045
R12309 GND.n4731 GND.n1728 8.33045
R12310 GND.n6060 GND.n1792 8.33045
R12311 GND.n6040 GND.n1817 8.33045
R12312 GND.n8083 GND.n8082 8.09508
R12313 GND.n6313 GND.n9 8.09508
R12314 GND.n3997 GND.t0 8.03295
R12315 GND.t6 GND.n2528 8.03295
R12316 GND.n6275 GND.n1462 7.95202
R12317 GND.n5864 GND.n5836 7.95202
R12318 GND.n5293 GND.n5234 7.95202
R12319 GND.n5042 GND.n5040 7.95202
R12320 GND.n6355 GND.n6351 7.95202
R12321 GND.n3779 GND.n3778 7.73546
R12322 GND.n3790 GND.n3516 7.73546
R12323 GND.n3789 GND.n3518 7.73546
R12324 GND.n3800 GND.n3509 7.73546
R12325 GND.n3801 GND.n3497 7.73546
R12326 GND.n3816 GND.n3499 7.73546
R12327 GND.n3827 GND.n3486 7.73546
R12328 GND.n3826 GND.n3489 7.73546
R12329 GND.n3837 GND.n3479 7.73546
R12330 GND.n3838 GND.n3468 7.73546
R12331 GND.n3853 GND.n3470 7.73546
R12332 GND.n3864 GND.n3458 7.73546
R12333 GND.n3863 GND.n3460 7.73546
R12334 GND.n3880 GND.n3450 7.73546
R12335 GND.n3881 GND.n3439 7.73546
R12336 GND.n3893 GND.n3442 7.73546
R12337 GND.n3884 GND.n3430 7.73546
R12338 GND.n3902 GND.n3433 7.73546
R12339 GND.n3989 GND.n3407 7.73546
R12340 GND.n3988 GND.n3410 7.73546
R12341 GND.n3909 GND.n3417 7.73546
R12342 GND.n3981 GND.n3419 7.73546
R12343 GND.n3952 GND.n3937 7.73546
R12344 GND.n3954 GND.n3934 7.73546
R12345 GND.n3959 GND.n3936 7.73546
R12346 GND.n3956 GND.n3920 7.73546
R12347 GND.n3968 GND.n3921 7.73546
R12348 GND.n3929 GND.n3395 7.73546
R12349 GND.n3998 GND.n3997 7.73546
R12350 GND.n4013 GND.n3386 7.73546
R12351 GND.n4024 GND.n3374 7.73546
R12352 GND.n4023 GND.n3377 7.73546
R12353 GND.n4034 GND.n3367 7.73546
R12354 GND.n4035 GND.n3356 7.73546
R12355 GND.n4050 GND.n3358 7.73546
R12356 GND.n4061 GND.n3346 7.73546
R12357 GND.n4060 GND.n3348 7.73546
R12358 GND.n4071 GND.n3338 7.73546
R12359 GND.n4072 GND.n3326 7.73546
R12360 GND.n4087 GND.n3329 7.73546
R12361 GND.n4098 GND.n3316 7.73546
R12362 GND.n4097 GND.n3318 7.73546
R12363 GND.n4130 GND.n3309 7.73546
R12364 GND.n4132 GND.n3299 7.73546
R12365 GND.n4142 GND.n3301 7.73546
R12366 GND.n4135 GND.n3293 7.73546
R12367 GND.n4151 GND.n3289 7.73546
R12368 GND.n4154 GND.n3290 7.73546
R12369 GND.t118 GND.n4652 7.73546
R12370 GND.n4763 GND.n4762 7.73546
R12371 GND.n6067 GND.n1784 7.73546
R12372 GND.n5439 GND.n2404 7.73546
R12373 GND.n5436 GND.n2406 7.73546
R12374 GND.n5050 GND.n2437 7.73546
R12375 GND.n5430 GND.n2446 7.73546
R12376 GND.n5058 GND.n2449 7.73546
R12377 GND.n5424 GND.n2457 7.73546
R12378 GND.n5065 GND.n2657 7.73546
R12379 GND.n5418 GND.n2467 7.73546
R12380 GND.n5073 GND.n2470 7.73546
R12381 GND.n5412 GND.n2477 7.73546
R12382 GND.n5080 GND.n2480 7.73546
R12383 GND.n5406 GND.n2488 7.73546
R12384 GND.n5088 GND.n2491 7.73546
R12385 GND.n5400 GND.n2498 7.73546
R12386 GND.n5095 GND.n2501 7.73546
R12387 GND.n5394 GND.n2509 7.73546
R12388 GND.n5103 GND.n2512 7.73546
R12389 GND.n5388 GND.n2519 7.73546
R12390 GND.n5110 GND.n2522 7.73546
R12391 GND.n5382 GND.n2528 7.73546
R12392 GND.n5122 GND.n2531 7.73546
R12393 GND.n5376 GND.n2538 7.73546
R12394 GND.n5373 GND.n2541 7.73546
R12395 GND.n5372 GND.n2545 7.73546
R12396 GND.n8078 GND.n32 7.73546
R12397 GND.n2552 GND.n34 7.73546
R12398 GND.n5364 GND.n5363 7.73546
R12399 GND.n5354 GND.n2555 7.73546
R12400 GND.n8071 GND.n51 7.73546
R12401 GND.n5348 GND.n5202 7.73546
R12402 GND.n8065 GND.n62 7.73546
R12403 GND.n5342 GND.n65 7.73546
R12404 GND.n8059 GND.n72 7.73546
R12405 GND.n5336 GND.n75 7.73546
R12406 GND.n8053 GND.n82 7.73546
R12407 GND.n5330 GND.n85 7.73546
R12408 GND.n8047 GND.n93 7.73546
R12409 GND.n5324 GND.n96 7.73546
R12410 GND.n8041 GND.n103 7.73546
R12411 GND.n5318 GND.n106 7.73546
R12412 GND.n8035 GND.n114 7.73546
R12413 GND.n5312 GND.n117 7.73546
R12414 GND.n8029 GND.n124 7.73546
R12415 GND.n5306 GND.n127 7.73546
R12416 GND.n8023 GND.n135 7.73546
R12417 GND.n5300 GND.n138 7.73546
R12418 GND.n8017 GND.n145 7.73546
R12419 GND.n7875 GND.n148 7.73546
R12420 GND.n4440 GND.t2 7.43796
R12421 GND.t2 GND.n4439 7.43796
R12422 GND.n5756 GND.t15 7.43796
R12423 GND.n2691 GND.t15 7.43796
R12424 GND.n4690 GND.n2765 7.14046
R12425 GND.n4762 GND.n2752 7.14046
R12426 GND.n6068 GND.n6067 7.14046
R12427 GND.n6381 GND.n1373 6.84296
R12428 GND.n291 GND.n154 6.84296
R12429 GND.n6004 GND.n6003 6.5566
R12430 GND.n4587 GND.n4586 6.5566
R12431 GND.n6152 GND.n6151 6.5566
R12432 GND.n5874 GND.n5873 6.5566
R12433 GND.n4714 GND.n2760 6.54546
R12434 GND.n4731 GND.n1722 6.54546
R12435 GND.n4846 GND.n1792 6.54546
R12436 GND.n4868 GND.n1817 6.54546
R12437 GND.t50 GND.n1842 6.54546
R12438 GND.n3989 GND.t18 6.24796
R12439 GND.n5202 GND.t10 6.24796
R12440 GND.n3 GND.n1 5.98039
R12441 GND.n19 GND.n17 5.98039
R12442 GND.n4652 GND.n1649 5.95047
R12443 GND.n4672 GND.n4671 5.95047
R12444 GND.n4755 GND.n4754 5.95047
R12445 GND.n6074 GND.n1774 5.95047
R12446 GND.n6033 GND.t133 5.95047
R12447 GND.n6026 GND.n1834 5.95047
R12448 GND.n5939 GND.n5834 5.95047
R12449 GND.n6008 GND.n1890 5.62001
R12450 GND.n6219 GND.n1573 5.62001
R12451 GND.n6219 GND.n6218 5.62001
R12452 GND.n5869 GND.n1890 5.62001
R12453 GND.n6123 GND.t57 5.35547
R12454 GND.n4719 GND.t40 5.35547
R12455 GND.n6047 GND.n1807 5.35547
R12456 GND.t47 GND.n1834 5.35547
R12457 GND.n5859 GND.n5836 5.23686
R12458 GND.n3318 GND.t84 5.05797
R12459 GND.n4691 GND.t77 5.05797
R12460 GND.n4877 GND.t43 5.05797
R12461 GND.n2657 GND.t53 5.05797
R12462 GND.n9 GND.n8 4.95764
R12463 GND.n8083 GND.n25 4.95764
R12464 GND.n2771 GND.n1652 4.76047
R12465 GND.n4667 GND.n1661 4.76047
R12466 GND.n6082 GND.n6081 4.76047
R12467 GND.n4747 GND.n4746 4.76047
R12468 GND.n5827 GND.n5826 4.76047
R12469 GND.n6019 GND.n6018 4.76047
R12470 GND.n5384 GND.n46 4.74817
R12471 GND.n44 GND.n38 4.74817
R12472 GND.n8075 GND.n39 4.74817
R12473 GND.n47 GND.n43 4.74817
R12474 GND.n2526 GND.n46 4.74817
R12475 GND.n2542 GND.n44 4.74817
R12476 GND.n8076 GND.n8075 4.74817
R12477 GND.n5361 GND.n43 4.74817
R12478 GND.n3404 GND.n3401 4.74817
R12479 GND.n3950 GND.n3400 4.74817
R12480 GND.n3946 GND.n3399 4.74817
R12481 GND.n3942 GND.n3398 4.74817
R12482 GND.n3995 GND.n3994 4.74817
R12483 GND.n2635 GND.n2634 4.74817
R12484 GND.n2630 GND.n2548 4.74817
R12485 GND.n5369 GND.n5368 4.74817
R12486 GND.n2551 GND.n2549 4.74817
R12487 GND.n5147 GND.n5146 4.74817
R12488 GND.n2636 GND.n2635 4.74817
R12489 GND.n2631 GND.n2630 4.74817
R12490 GND.n5370 GND.n5369 4.74817
R12491 GND.n5367 GND.n2549 4.74817
R12492 GND.n5146 GND.n5145 4.74817
R12493 GND.n3986 GND.n3985 4.74817
R12494 GND.n3932 GND.n3931 4.74817
R12495 GND.n3963 GND.n3962 4.74817
R12496 GND.n3965 GND.n3964 4.74817
R12497 GND.n3985 GND.n3984 4.74817
R12498 GND.n3931 GND.n3415 4.74817
R12499 GND.n3962 GND.n3961 4.74817
R12500 GND.n3966 GND.n3965 4.74817
R12501 GND.n3939 GND.n3401 4.74817
R12502 GND.n3940 GND.n3400 4.74817
R12503 GND.n3949 GND.n3399 4.74817
R12504 GND.n3945 GND.n3398 4.74817
R12505 GND.n3994 GND.n3397 4.74817
R12506 GND.n8 GND.n0 4.70093
R12507 GND.n25 GND.n24 4.70093
R12508 GND.n3 GND.n2 4.63843
R12509 GND.n5 GND.n4 4.63843
R12510 GND.n7 GND.n6 4.63843
R12511 GND.n19 GND.n18 4.63843
R12512 GND.n21 GND.n20 4.63843
R12513 GND.n23 GND.n22 4.63843
R12514 GND.n5521 GND.n2355 4.6132
R12515 GND.n6220 GND.n1571 4.6132
R12516 GND.t37 GND.n1705 4.46297
R12517 GND.n4856 GND.t26 4.46297
R12518 GND.n16 GND.n12 4.40104
R12519 GND.n1645 GND.n1644 4.38232
R12520 GND.n5863 GND.n5862 4.38232
R12521 GND.n4671 GND.t106 4.16548
R12522 GND.n6116 GND.n6115 4.16548
R12523 GND.n4727 GND.n1720 4.16548
R12524 GND.n4841 GND.n1800 4.16548
R12525 GND.n2723 GND.n1809 4.16548
R12526 GND.n2723 GND.t109 4.16548
R12527 GND.n6003 GND.n6002 4.05904
R12528 GND.n4588 GND.n4587 4.05904
R12529 GND.n6155 GND.n6151 4.05904
R12530 GND.n5875 GND.n5874 4.05904
R12531 GND.n4237 GND.t154 3.86798
R12532 GND.n5666 GND.t164 3.86798
R12533 GND.n3245 GND.n3195 3.68535
R12534 GND.n5485 GND.n5484 3.68535
R12535 GND.n7916 GND.n249 3.68535
R12536 GND.n3716 GND.n3713 3.68535
R12537 GND.n6130 GND.n6129 3.57048
R12538 GND.n4715 GND.t148 3.57048
R12539 GND.n6088 GND.n1750 3.57048
R12540 GND.n4812 GND.n4809 3.57048
R12541 GND.n5821 GND.n1896 3.57048
R12542 GND.n5818 GND.t47 3.57048
R12543 GND.n5827 GND.t50 3.57048
R12544 GND.n16 GND.n15 3.53792
R12545 GND.n6122 GND.n1682 2.97548
R12546 GND.n6096 GND.n6095 2.97548
R12547 GND.n6061 GND.n1790 2.97548
R12548 GND.t88 GND.n6039 2.97548
R12549 GND.n6039 GND.n1819 2.97548
R12550 GND.t115 GND.n1871 2.97548
R12551 GND.n3248 GND.n3195 2.90959
R12552 GND.n5484 GND.n5483 2.90959
R12553 GND.n251 GND.n249 2.90959
R12554 GND.n3713 GND.n3549 2.90959
R12555 GND.t77 GND.n4690 2.67798
R12556 GND.n6033 GND.t43 2.67798
R12557 GND.n6123 GND.n1680 2.38049
R12558 GND.n4735 GND.n1731 2.38049
R12559 GND.n4818 GND.n4817 2.38049
R12560 GND.n2713 GND.n2712 2.38049
R12561 GND.n8074 GND.n46 2.27742
R12562 GND.n8074 GND.n44 2.27742
R12563 GND.n8075 GND.n8074 2.27742
R12564 GND.n8074 GND.n43 2.27742
R12565 GND.n2635 GND.n42 2.27742
R12566 GND.n2630 GND.n42 2.27742
R12567 GND.n5369 GND.n42 2.27742
R12568 GND.n2549 GND.n42 2.27742
R12569 GND.n5146 GND.n42 2.27742
R12570 GND.n3985 GND.n3382 2.27742
R12571 GND.n3931 GND.n3382 2.27742
R12572 GND.n3962 GND.n3382 2.27742
R12573 GND.n3965 GND.n3382 2.27742
R12574 GND.n3993 GND.n3401 2.27742
R12575 GND.n3993 GND.n3400 2.27742
R12576 GND.n3993 GND.n3399 2.27742
R12577 GND.n3993 GND.n3398 2.27742
R12578 GND.n3994 GND.n3993 2.27742
R12579 GND.n6089 GND.n1748 1.78549
R12580 GND.n4808 GND.n1782 1.78549
R12581 GND.n4879 GND.n1826 1.78549
R12582 GND.n5834 GND.t91 1.78549
R12583 GND.n8 GND.n7 1.68153
R12584 GND.n25 GND.n23 1.68153
R12585 GND GND.n9 1.67307
R12586 GND.n11 GND.n10 1.52182
R12587 GND.n12 GND.n11 1.52182
R12588 GND.n14 GND.n13 1.52182
R12589 GND.n15 GND.n14 1.52182
R12590 GND.n2940 GND.t13 1.48799
R12591 GND.t20 GND.n2785 1.48799
R12592 GND.n6215 GND.n1578 1.48799
R12593 GND.n6011 GND.n1871 1.48799
R12594 GND.n5799 GND.t167 1.48799
R12595 GND.n4969 GND.t4 1.48799
R12596 GND.n5 GND.n3 1.34245
R12597 GND.n7 GND.n5 1.34245
R12598 GND.n21 GND.n19 1.34245
R12599 GND.n23 GND.n21 1.34245
R12600 GND.n4653 GND.t118 1.19049
R12601 GND.t151 GND.n2771 1.19049
R12602 GND.n2766 GND.t161 1.19049
R12603 GND.n4715 GND.n1696 1.19049
R12604 GND.n6103 GND.n6102 1.19049
R12605 GND.n4845 GND.n4842 1.19049
R12606 GND.n2722 GND.n2721 1.19049
R12607 GND.t133 GND.n6032 1.19049
R12608 GND.n4725 GND.t37 0.892995
R12609 GND.n4735 GND.t169 0.892995
R12610 GND.n4818 GND.t23 0.892995
R12611 GND.n6053 GND.t26 0.892995
R12612 GND.n1627 GND.n1625 0.716017
R12613 GND.n5857 GND.n5855 0.716017
R12614 GND.n8084 GND.n8083 0.68811
R12615 GND.n6144 GND.n6143 0.595497
R12616 GND.n6137 GND.n6136 0.595497
R12617 GND.t161 GND.n1671 0.595497
R12618 GND.n4753 GND.n1764 0.595497
R12619 GND.n6075 GND.n1772 0.595497
R12620 GND.n6025 GND.n1836 0.595497
R12621 GND.n5833 GND.n1844 0.595497
R12622 GND.n8013 GND.n8012 0.544707
R12623 GND.n2440 GND.n2317 0.544707
R12624 GND.n6270 GND.n1516 0.544707
R12625 GND.n3782 GND.n3523 0.544707
R12626 GND.n4198 GND.n3035 0.532512
R12627 GND.n2238 GND.n2237 0.532512
R12628 GND.n5295 GND.n5294 0.529463
R12629 GND.n6350 GND.n6349 0.529463
R12630 GND GND.n8084 0.49494
R12631 GND.n6629 GND.n6628 0.474585
R12632 GND.n7590 GND.n505 0.474585
R12633 GND.n7751 GND.n7750 0.474585
R12634 GND.n6500 GND.n6499 0.474585
R12635 GND.n8074 GND.n42 0.389875
R12636 GND.n3993 GND.n3382 0.389875
R12637 GND.n5044 GND.n5043 0.366136
R12638 GND.n6277 GND.n6276 0.366136
R12639 GND.n8084 GND.n16 0.365377
R12640 GND.n7880 GND.n7879 0.306902
R12641 GND.n5445 GND.n5443 0.306902
R12642 GND.n3764 GND.n3763 0.306902
R12643 GND.n4158 GND.n3168 0.306902
R12644 GND.n7879 GND.n286 0.291659
R12645 GND.n3764 GND.n1376 0.291659
R12646 GND.n3122 GND.n3121 0.230683
R12647 GND.n5037 GND.n2667 0.230683
R12648 GND.n2355 GND.n2353 0.229039
R12649 GND.n2358 GND.n2355 0.229039
R12650 GND.n1571 GND.n1566 0.229039
R12651 GND.n3211 GND.n1571 0.229039
R12652 GND.n6630 GND.n6629 0.152939
R12653 GND.n6630 GND.n1081 0.152939
R12654 GND.n6638 GND.n1081 0.152939
R12655 GND.n6639 GND.n6638 0.152939
R12656 GND.n6640 GND.n6639 0.152939
R12657 GND.n6640 GND.n1075 0.152939
R12658 GND.n6648 GND.n1075 0.152939
R12659 GND.n6649 GND.n6648 0.152939
R12660 GND.n6650 GND.n6649 0.152939
R12661 GND.n6650 GND.n1069 0.152939
R12662 GND.n6658 GND.n1069 0.152939
R12663 GND.n6659 GND.n6658 0.152939
R12664 GND.n6660 GND.n6659 0.152939
R12665 GND.n6660 GND.n1063 0.152939
R12666 GND.n6668 GND.n1063 0.152939
R12667 GND.n6669 GND.n6668 0.152939
R12668 GND.n6670 GND.n6669 0.152939
R12669 GND.n6670 GND.n1057 0.152939
R12670 GND.n6678 GND.n1057 0.152939
R12671 GND.n6679 GND.n6678 0.152939
R12672 GND.n6680 GND.n6679 0.152939
R12673 GND.n6680 GND.n1051 0.152939
R12674 GND.n6688 GND.n1051 0.152939
R12675 GND.n6689 GND.n6688 0.152939
R12676 GND.n6690 GND.n6689 0.152939
R12677 GND.n6690 GND.n1045 0.152939
R12678 GND.n6698 GND.n1045 0.152939
R12679 GND.n6699 GND.n6698 0.152939
R12680 GND.n6700 GND.n6699 0.152939
R12681 GND.n6700 GND.n1039 0.152939
R12682 GND.n6708 GND.n1039 0.152939
R12683 GND.n6709 GND.n6708 0.152939
R12684 GND.n6710 GND.n6709 0.152939
R12685 GND.n6710 GND.n1033 0.152939
R12686 GND.n6718 GND.n1033 0.152939
R12687 GND.n6719 GND.n6718 0.152939
R12688 GND.n6720 GND.n6719 0.152939
R12689 GND.n6720 GND.n1027 0.152939
R12690 GND.n6728 GND.n1027 0.152939
R12691 GND.n6729 GND.n6728 0.152939
R12692 GND.n6730 GND.n6729 0.152939
R12693 GND.n6730 GND.n1021 0.152939
R12694 GND.n6738 GND.n1021 0.152939
R12695 GND.n6739 GND.n6738 0.152939
R12696 GND.n6740 GND.n6739 0.152939
R12697 GND.n6740 GND.n1015 0.152939
R12698 GND.n6748 GND.n1015 0.152939
R12699 GND.n6749 GND.n6748 0.152939
R12700 GND.n6750 GND.n6749 0.152939
R12701 GND.n6750 GND.n1009 0.152939
R12702 GND.n6758 GND.n1009 0.152939
R12703 GND.n6759 GND.n6758 0.152939
R12704 GND.n6760 GND.n6759 0.152939
R12705 GND.n6760 GND.n1003 0.152939
R12706 GND.n6768 GND.n1003 0.152939
R12707 GND.n6769 GND.n6768 0.152939
R12708 GND.n6770 GND.n6769 0.152939
R12709 GND.n6770 GND.n997 0.152939
R12710 GND.n6778 GND.n997 0.152939
R12711 GND.n6779 GND.n6778 0.152939
R12712 GND.n6780 GND.n6779 0.152939
R12713 GND.n6780 GND.n991 0.152939
R12714 GND.n6788 GND.n991 0.152939
R12715 GND.n6789 GND.n6788 0.152939
R12716 GND.n6790 GND.n6789 0.152939
R12717 GND.n6790 GND.n985 0.152939
R12718 GND.n6798 GND.n985 0.152939
R12719 GND.n6799 GND.n6798 0.152939
R12720 GND.n6800 GND.n6799 0.152939
R12721 GND.n6800 GND.n979 0.152939
R12722 GND.n6808 GND.n979 0.152939
R12723 GND.n6809 GND.n6808 0.152939
R12724 GND.n6810 GND.n6809 0.152939
R12725 GND.n6810 GND.n973 0.152939
R12726 GND.n6818 GND.n973 0.152939
R12727 GND.n6819 GND.n6818 0.152939
R12728 GND.n6820 GND.n6819 0.152939
R12729 GND.n6820 GND.n967 0.152939
R12730 GND.n6828 GND.n967 0.152939
R12731 GND.n6829 GND.n6828 0.152939
R12732 GND.n6830 GND.n6829 0.152939
R12733 GND.n6830 GND.n961 0.152939
R12734 GND.n6838 GND.n961 0.152939
R12735 GND.n6839 GND.n6838 0.152939
R12736 GND.n6840 GND.n6839 0.152939
R12737 GND.n6840 GND.n955 0.152939
R12738 GND.n6848 GND.n955 0.152939
R12739 GND.n6849 GND.n6848 0.152939
R12740 GND.n6850 GND.n6849 0.152939
R12741 GND.n6850 GND.n949 0.152939
R12742 GND.n6858 GND.n949 0.152939
R12743 GND.n6859 GND.n6858 0.152939
R12744 GND.n6860 GND.n6859 0.152939
R12745 GND.n6860 GND.n943 0.152939
R12746 GND.n6868 GND.n943 0.152939
R12747 GND.n6869 GND.n6868 0.152939
R12748 GND.n6870 GND.n6869 0.152939
R12749 GND.n6870 GND.n937 0.152939
R12750 GND.n6878 GND.n937 0.152939
R12751 GND.n6879 GND.n6878 0.152939
R12752 GND.n6880 GND.n6879 0.152939
R12753 GND.n6880 GND.n931 0.152939
R12754 GND.n6888 GND.n931 0.152939
R12755 GND.n6889 GND.n6888 0.152939
R12756 GND.n6890 GND.n6889 0.152939
R12757 GND.n6890 GND.n925 0.152939
R12758 GND.n6898 GND.n925 0.152939
R12759 GND.n6899 GND.n6898 0.152939
R12760 GND.n6900 GND.n6899 0.152939
R12761 GND.n6900 GND.n919 0.152939
R12762 GND.n6908 GND.n919 0.152939
R12763 GND.n6909 GND.n6908 0.152939
R12764 GND.n6910 GND.n6909 0.152939
R12765 GND.n6910 GND.n913 0.152939
R12766 GND.n6918 GND.n913 0.152939
R12767 GND.n6919 GND.n6918 0.152939
R12768 GND.n6920 GND.n6919 0.152939
R12769 GND.n6920 GND.n907 0.152939
R12770 GND.n6928 GND.n907 0.152939
R12771 GND.n6929 GND.n6928 0.152939
R12772 GND.n6930 GND.n6929 0.152939
R12773 GND.n6930 GND.n901 0.152939
R12774 GND.n6938 GND.n901 0.152939
R12775 GND.n6939 GND.n6938 0.152939
R12776 GND.n6940 GND.n6939 0.152939
R12777 GND.n6940 GND.n895 0.152939
R12778 GND.n6948 GND.n895 0.152939
R12779 GND.n6949 GND.n6948 0.152939
R12780 GND.n6950 GND.n6949 0.152939
R12781 GND.n6950 GND.n889 0.152939
R12782 GND.n6958 GND.n889 0.152939
R12783 GND.n6959 GND.n6958 0.152939
R12784 GND.n6960 GND.n6959 0.152939
R12785 GND.n6960 GND.n883 0.152939
R12786 GND.n6968 GND.n883 0.152939
R12787 GND.n6969 GND.n6968 0.152939
R12788 GND.n6970 GND.n6969 0.152939
R12789 GND.n6970 GND.n877 0.152939
R12790 GND.n6978 GND.n877 0.152939
R12791 GND.n6979 GND.n6978 0.152939
R12792 GND.n6980 GND.n6979 0.152939
R12793 GND.n6980 GND.n871 0.152939
R12794 GND.n6988 GND.n871 0.152939
R12795 GND.n6989 GND.n6988 0.152939
R12796 GND.n6990 GND.n6989 0.152939
R12797 GND.n6990 GND.n865 0.152939
R12798 GND.n6998 GND.n865 0.152939
R12799 GND.n6999 GND.n6998 0.152939
R12800 GND.n7000 GND.n6999 0.152939
R12801 GND.n7000 GND.n859 0.152939
R12802 GND.n7008 GND.n859 0.152939
R12803 GND.n7009 GND.n7008 0.152939
R12804 GND.n7010 GND.n7009 0.152939
R12805 GND.n7010 GND.n853 0.152939
R12806 GND.n7018 GND.n853 0.152939
R12807 GND.n7019 GND.n7018 0.152939
R12808 GND.n7020 GND.n7019 0.152939
R12809 GND.n7020 GND.n847 0.152939
R12810 GND.n7028 GND.n847 0.152939
R12811 GND.n7029 GND.n7028 0.152939
R12812 GND.n7030 GND.n7029 0.152939
R12813 GND.n7030 GND.n841 0.152939
R12814 GND.n7038 GND.n841 0.152939
R12815 GND.n7039 GND.n7038 0.152939
R12816 GND.n7040 GND.n7039 0.152939
R12817 GND.n7040 GND.n835 0.152939
R12818 GND.n7048 GND.n835 0.152939
R12819 GND.n7049 GND.n7048 0.152939
R12820 GND.n7050 GND.n7049 0.152939
R12821 GND.n7050 GND.n829 0.152939
R12822 GND.n7058 GND.n829 0.152939
R12823 GND.n7059 GND.n7058 0.152939
R12824 GND.n7060 GND.n7059 0.152939
R12825 GND.n7060 GND.n823 0.152939
R12826 GND.n7068 GND.n823 0.152939
R12827 GND.n7069 GND.n7068 0.152939
R12828 GND.n7070 GND.n7069 0.152939
R12829 GND.n7070 GND.n817 0.152939
R12830 GND.n7078 GND.n817 0.152939
R12831 GND.n7079 GND.n7078 0.152939
R12832 GND.n7080 GND.n7079 0.152939
R12833 GND.n7080 GND.n811 0.152939
R12834 GND.n7088 GND.n811 0.152939
R12835 GND.n7089 GND.n7088 0.152939
R12836 GND.n7090 GND.n7089 0.152939
R12837 GND.n7090 GND.n805 0.152939
R12838 GND.n7098 GND.n805 0.152939
R12839 GND.n7099 GND.n7098 0.152939
R12840 GND.n7100 GND.n7099 0.152939
R12841 GND.n7100 GND.n799 0.152939
R12842 GND.n7108 GND.n799 0.152939
R12843 GND.n7109 GND.n7108 0.152939
R12844 GND.n7110 GND.n7109 0.152939
R12845 GND.n7110 GND.n793 0.152939
R12846 GND.n7118 GND.n793 0.152939
R12847 GND.n7119 GND.n7118 0.152939
R12848 GND.n7120 GND.n7119 0.152939
R12849 GND.n7120 GND.n787 0.152939
R12850 GND.n7128 GND.n787 0.152939
R12851 GND.n7129 GND.n7128 0.152939
R12852 GND.n7130 GND.n7129 0.152939
R12853 GND.n7130 GND.n781 0.152939
R12854 GND.n7138 GND.n781 0.152939
R12855 GND.n7139 GND.n7138 0.152939
R12856 GND.n7140 GND.n7139 0.152939
R12857 GND.n7140 GND.n775 0.152939
R12858 GND.n7148 GND.n775 0.152939
R12859 GND.n7149 GND.n7148 0.152939
R12860 GND.n7150 GND.n7149 0.152939
R12861 GND.n7150 GND.n769 0.152939
R12862 GND.n7158 GND.n769 0.152939
R12863 GND.n7159 GND.n7158 0.152939
R12864 GND.n7160 GND.n7159 0.152939
R12865 GND.n7160 GND.n763 0.152939
R12866 GND.n7168 GND.n763 0.152939
R12867 GND.n7169 GND.n7168 0.152939
R12868 GND.n7170 GND.n7169 0.152939
R12869 GND.n7170 GND.n757 0.152939
R12870 GND.n7178 GND.n757 0.152939
R12871 GND.n7179 GND.n7178 0.152939
R12872 GND.n7180 GND.n7179 0.152939
R12873 GND.n7180 GND.n751 0.152939
R12874 GND.n7188 GND.n751 0.152939
R12875 GND.n7189 GND.n7188 0.152939
R12876 GND.n7190 GND.n7189 0.152939
R12877 GND.n7190 GND.n745 0.152939
R12878 GND.n7198 GND.n745 0.152939
R12879 GND.n7199 GND.n7198 0.152939
R12880 GND.n7200 GND.n7199 0.152939
R12881 GND.n7200 GND.n739 0.152939
R12882 GND.n7208 GND.n739 0.152939
R12883 GND.n7209 GND.n7208 0.152939
R12884 GND.n7210 GND.n7209 0.152939
R12885 GND.n7210 GND.n733 0.152939
R12886 GND.n7218 GND.n733 0.152939
R12887 GND.n7219 GND.n7218 0.152939
R12888 GND.n7220 GND.n7219 0.152939
R12889 GND.n7220 GND.n727 0.152939
R12890 GND.n7228 GND.n727 0.152939
R12891 GND.n7229 GND.n7228 0.152939
R12892 GND.n7230 GND.n7229 0.152939
R12893 GND.n7230 GND.n721 0.152939
R12894 GND.n7238 GND.n721 0.152939
R12895 GND.n7239 GND.n7238 0.152939
R12896 GND.n7240 GND.n7239 0.152939
R12897 GND.n7240 GND.n715 0.152939
R12898 GND.n7248 GND.n715 0.152939
R12899 GND.n7249 GND.n7248 0.152939
R12900 GND.n7250 GND.n7249 0.152939
R12901 GND.n7250 GND.n709 0.152939
R12902 GND.n7258 GND.n709 0.152939
R12903 GND.n7259 GND.n7258 0.152939
R12904 GND.n7260 GND.n7259 0.152939
R12905 GND.n7260 GND.n703 0.152939
R12906 GND.n7268 GND.n703 0.152939
R12907 GND.n7269 GND.n7268 0.152939
R12908 GND.n7270 GND.n7269 0.152939
R12909 GND.n7270 GND.n697 0.152939
R12910 GND.n7278 GND.n697 0.152939
R12911 GND.n7279 GND.n7278 0.152939
R12912 GND.n7280 GND.n7279 0.152939
R12913 GND.n7280 GND.n691 0.152939
R12914 GND.n7288 GND.n691 0.152939
R12915 GND.n7289 GND.n7288 0.152939
R12916 GND.n7290 GND.n7289 0.152939
R12917 GND.n7290 GND.n685 0.152939
R12918 GND.n7298 GND.n685 0.152939
R12919 GND.n7299 GND.n7298 0.152939
R12920 GND.n7300 GND.n7299 0.152939
R12921 GND.n7300 GND.n679 0.152939
R12922 GND.n7308 GND.n679 0.152939
R12923 GND.n7309 GND.n7308 0.152939
R12924 GND.n7310 GND.n7309 0.152939
R12925 GND.n7310 GND.n673 0.152939
R12926 GND.n7318 GND.n673 0.152939
R12927 GND.n7319 GND.n7318 0.152939
R12928 GND.n7320 GND.n7319 0.152939
R12929 GND.n7320 GND.n667 0.152939
R12930 GND.n7328 GND.n667 0.152939
R12931 GND.n7329 GND.n7328 0.152939
R12932 GND.n7330 GND.n7329 0.152939
R12933 GND.n7330 GND.n661 0.152939
R12934 GND.n7338 GND.n661 0.152939
R12935 GND.n7339 GND.n7338 0.152939
R12936 GND.n7340 GND.n7339 0.152939
R12937 GND.n7340 GND.n655 0.152939
R12938 GND.n7348 GND.n655 0.152939
R12939 GND.n7349 GND.n7348 0.152939
R12940 GND.n7350 GND.n7349 0.152939
R12941 GND.n7350 GND.n649 0.152939
R12942 GND.n7358 GND.n649 0.152939
R12943 GND.n7359 GND.n7358 0.152939
R12944 GND.n7360 GND.n7359 0.152939
R12945 GND.n7360 GND.n643 0.152939
R12946 GND.n7368 GND.n643 0.152939
R12947 GND.n7369 GND.n7368 0.152939
R12948 GND.n7370 GND.n7369 0.152939
R12949 GND.n7370 GND.n637 0.152939
R12950 GND.n7378 GND.n637 0.152939
R12951 GND.n7379 GND.n7378 0.152939
R12952 GND.n7380 GND.n7379 0.152939
R12953 GND.n7380 GND.n631 0.152939
R12954 GND.n7388 GND.n631 0.152939
R12955 GND.n7389 GND.n7388 0.152939
R12956 GND.n7390 GND.n7389 0.152939
R12957 GND.n7390 GND.n625 0.152939
R12958 GND.n7398 GND.n625 0.152939
R12959 GND.n7399 GND.n7398 0.152939
R12960 GND.n7400 GND.n7399 0.152939
R12961 GND.n7400 GND.n619 0.152939
R12962 GND.n7408 GND.n619 0.152939
R12963 GND.n7409 GND.n7408 0.152939
R12964 GND.n7410 GND.n7409 0.152939
R12965 GND.n7410 GND.n613 0.152939
R12966 GND.n7418 GND.n613 0.152939
R12967 GND.n7419 GND.n7418 0.152939
R12968 GND.n7420 GND.n7419 0.152939
R12969 GND.n7420 GND.n607 0.152939
R12970 GND.n7428 GND.n607 0.152939
R12971 GND.n7429 GND.n7428 0.152939
R12972 GND.n7430 GND.n7429 0.152939
R12973 GND.n7430 GND.n601 0.152939
R12974 GND.n7438 GND.n601 0.152939
R12975 GND.n7439 GND.n7438 0.152939
R12976 GND.n7440 GND.n7439 0.152939
R12977 GND.n7440 GND.n595 0.152939
R12978 GND.n7448 GND.n595 0.152939
R12979 GND.n7449 GND.n7448 0.152939
R12980 GND.n7450 GND.n7449 0.152939
R12981 GND.n7450 GND.n589 0.152939
R12982 GND.n7458 GND.n589 0.152939
R12983 GND.n7459 GND.n7458 0.152939
R12984 GND.n7460 GND.n7459 0.152939
R12985 GND.n7460 GND.n583 0.152939
R12986 GND.n7468 GND.n583 0.152939
R12987 GND.n7469 GND.n7468 0.152939
R12988 GND.n7470 GND.n7469 0.152939
R12989 GND.n7470 GND.n577 0.152939
R12990 GND.n7478 GND.n577 0.152939
R12991 GND.n7479 GND.n7478 0.152939
R12992 GND.n7480 GND.n7479 0.152939
R12993 GND.n7480 GND.n571 0.152939
R12994 GND.n7488 GND.n571 0.152939
R12995 GND.n7489 GND.n7488 0.152939
R12996 GND.n7490 GND.n7489 0.152939
R12997 GND.n7490 GND.n565 0.152939
R12998 GND.n7498 GND.n565 0.152939
R12999 GND.n7499 GND.n7498 0.152939
R13000 GND.n7500 GND.n7499 0.152939
R13001 GND.n7500 GND.n559 0.152939
R13002 GND.n7508 GND.n559 0.152939
R13003 GND.n7509 GND.n7508 0.152939
R13004 GND.n7510 GND.n7509 0.152939
R13005 GND.n7510 GND.n553 0.152939
R13006 GND.n7518 GND.n553 0.152939
R13007 GND.n7519 GND.n7518 0.152939
R13008 GND.n7520 GND.n7519 0.152939
R13009 GND.n7520 GND.n547 0.152939
R13010 GND.n7528 GND.n547 0.152939
R13011 GND.n7529 GND.n7528 0.152939
R13012 GND.n7530 GND.n7529 0.152939
R13013 GND.n7530 GND.n541 0.152939
R13014 GND.n7538 GND.n541 0.152939
R13015 GND.n7539 GND.n7538 0.152939
R13016 GND.n7540 GND.n7539 0.152939
R13017 GND.n7540 GND.n535 0.152939
R13018 GND.n7548 GND.n535 0.152939
R13019 GND.n7549 GND.n7548 0.152939
R13020 GND.n7550 GND.n7549 0.152939
R13021 GND.n7550 GND.n529 0.152939
R13022 GND.n7558 GND.n529 0.152939
R13023 GND.n7559 GND.n7558 0.152939
R13024 GND.n7560 GND.n7559 0.152939
R13025 GND.n7560 GND.n523 0.152939
R13026 GND.n7568 GND.n523 0.152939
R13027 GND.n7569 GND.n7568 0.152939
R13028 GND.n7570 GND.n7569 0.152939
R13029 GND.n7570 GND.n517 0.152939
R13030 GND.n7578 GND.n517 0.152939
R13031 GND.n7579 GND.n7578 0.152939
R13032 GND.n7580 GND.n7579 0.152939
R13033 GND.n7580 GND.n511 0.152939
R13034 GND.n7588 GND.n511 0.152939
R13035 GND.n7589 GND.n7588 0.152939
R13036 GND.n7590 GND.n7589 0.152939
R13037 GND.n7598 GND.n505 0.152939
R13038 GND.n7599 GND.n7598 0.152939
R13039 GND.n7600 GND.n7599 0.152939
R13040 GND.n7600 GND.n499 0.152939
R13041 GND.n7608 GND.n499 0.152939
R13042 GND.n7609 GND.n7608 0.152939
R13043 GND.n7610 GND.n7609 0.152939
R13044 GND.n7610 GND.n493 0.152939
R13045 GND.n7618 GND.n493 0.152939
R13046 GND.n7619 GND.n7618 0.152939
R13047 GND.n7620 GND.n7619 0.152939
R13048 GND.n7620 GND.n487 0.152939
R13049 GND.n7628 GND.n487 0.152939
R13050 GND.n7629 GND.n7628 0.152939
R13051 GND.n7630 GND.n7629 0.152939
R13052 GND.n7630 GND.n481 0.152939
R13053 GND.n7638 GND.n481 0.152939
R13054 GND.n7639 GND.n7638 0.152939
R13055 GND.n7640 GND.n7639 0.152939
R13056 GND.n7640 GND.n475 0.152939
R13057 GND.n7648 GND.n475 0.152939
R13058 GND.n7649 GND.n7648 0.152939
R13059 GND.n7650 GND.n7649 0.152939
R13060 GND.n7650 GND.n469 0.152939
R13061 GND.n7658 GND.n469 0.152939
R13062 GND.n7659 GND.n7658 0.152939
R13063 GND.n7660 GND.n7659 0.152939
R13064 GND.n7660 GND.n463 0.152939
R13065 GND.n7668 GND.n463 0.152939
R13066 GND.n7669 GND.n7668 0.152939
R13067 GND.n7670 GND.n7669 0.152939
R13068 GND.n7670 GND.n457 0.152939
R13069 GND.n7678 GND.n457 0.152939
R13070 GND.n7679 GND.n7678 0.152939
R13071 GND.n7680 GND.n7679 0.152939
R13072 GND.n7680 GND.n451 0.152939
R13073 GND.n7688 GND.n451 0.152939
R13074 GND.n7689 GND.n7688 0.152939
R13075 GND.n7690 GND.n7689 0.152939
R13076 GND.n7690 GND.n445 0.152939
R13077 GND.n7698 GND.n445 0.152939
R13078 GND.n7699 GND.n7698 0.152939
R13079 GND.n7700 GND.n7699 0.152939
R13080 GND.n7700 GND.n439 0.152939
R13081 GND.n7708 GND.n439 0.152939
R13082 GND.n7709 GND.n7708 0.152939
R13083 GND.n7710 GND.n7709 0.152939
R13084 GND.n7710 GND.n433 0.152939
R13085 GND.n7718 GND.n433 0.152939
R13086 GND.n7719 GND.n7718 0.152939
R13087 GND.n7720 GND.n7719 0.152939
R13088 GND.n7720 GND.n427 0.152939
R13089 GND.n7728 GND.n427 0.152939
R13090 GND.n7729 GND.n7728 0.152939
R13091 GND.n7730 GND.n7729 0.152939
R13092 GND.n7730 GND.n421 0.152939
R13093 GND.n7738 GND.n421 0.152939
R13094 GND.n7739 GND.n7738 0.152939
R13095 GND.n7741 GND.n7739 0.152939
R13096 GND.n7741 GND.n7740 0.152939
R13097 GND.n7740 GND.n415 0.152939
R13098 GND.n7750 GND.n415 0.152939
R13099 GND.n5149 GND.n5148 0.152939
R13100 GND.n5150 GND.n5149 0.152939
R13101 GND.n5153 GND.n5150 0.152939
R13102 GND.n5154 GND.n5153 0.152939
R13103 GND.n5155 GND.n5154 0.152939
R13104 GND.n5156 GND.n5155 0.152939
R13105 GND.n5159 GND.n5156 0.152939
R13106 GND.n5160 GND.n5159 0.152939
R13107 GND.n5161 GND.n5160 0.152939
R13108 GND.n5162 GND.n5161 0.152939
R13109 GND.n5165 GND.n5162 0.152939
R13110 GND.n5166 GND.n5165 0.152939
R13111 GND.n5167 GND.n5166 0.152939
R13112 GND.n5168 GND.n5167 0.152939
R13113 GND.n5171 GND.n5168 0.152939
R13114 GND.n5172 GND.n5171 0.152939
R13115 GND.n5174 GND.n5172 0.152939
R13116 GND.n5174 GND.n5173 0.152939
R13117 GND.n5173 GND.n295 0.152939
R13118 GND.n296 GND.n295 0.152939
R13119 GND.n297 GND.n296 0.152939
R13120 GND.n302 GND.n297 0.152939
R13121 GND.n303 GND.n302 0.152939
R13122 GND.n304 GND.n303 0.152939
R13123 GND.n305 GND.n304 0.152939
R13124 GND.n310 GND.n305 0.152939
R13125 GND.n311 GND.n310 0.152939
R13126 GND.n312 GND.n311 0.152939
R13127 GND.n313 GND.n312 0.152939
R13128 GND.n318 GND.n313 0.152939
R13129 GND.n319 GND.n318 0.152939
R13130 GND.n320 GND.n319 0.152939
R13131 GND.n321 GND.n320 0.152939
R13132 GND.n326 GND.n321 0.152939
R13133 GND.n327 GND.n326 0.152939
R13134 GND.n328 GND.n327 0.152939
R13135 GND.n329 GND.n328 0.152939
R13136 GND.n334 GND.n329 0.152939
R13137 GND.n335 GND.n334 0.152939
R13138 GND.n336 GND.n335 0.152939
R13139 GND.n337 GND.n336 0.152939
R13140 GND.n342 GND.n337 0.152939
R13141 GND.n343 GND.n342 0.152939
R13142 GND.n344 GND.n343 0.152939
R13143 GND.n345 GND.n344 0.152939
R13144 GND.n350 GND.n345 0.152939
R13145 GND.n351 GND.n350 0.152939
R13146 GND.n352 GND.n351 0.152939
R13147 GND.n353 GND.n352 0.152939
R13148 GND.n358 GND.n353 0.152939
R13149 GND.n359 GND.n358 0.152939
R13150 GND.n360 GND.n359 0.152939
R13151 GND.n361 GND.n360 0.152939
R13152 GND.n366 GND.n361 0.152939
R13153 GND.n367 GND.n366 0.152939
R13154 GND.n368 GND.n367 0.152939
R13155 GND.n369 GND.n368 0.152939
R13156 GND.n374 GND.n369 0.152939
R13157 GND.n375 GND.n374 0.152939
R13158 GND.n376 GND.n375 0.152939
R13159 GND.n377 GND.n376 0.152939
R13160 GND.n382 GND.n377 0.152939
R13161 GND.n383 GND.n382 0.152939
R13162 GND.n384 GND.n383 0.152939
R13163 GND.n385 GND.n384 0.152939
R13164 GND.n390 GND.n385 0.152939
R13165 GND.n391 GND.n390 0.152939
R13166 GND.n392 GND.n391 0.152939
R13167 GND.n393 GND.n392 0.152939
R13168 GND.n398 GND.n393 0.152939
R13169 GND.n399 GND.n398 0.152939
R13170 GND.n400 GND.n399 0.152939
R13171 GND.n401 GND.n400 0.152939
R13172 GND.n406 GND.n401 0.152939
R13173 GND.n407 GND.n406 0.152939
R13174 GND.n408 GND.n407 0.152939
R13175 GND.n409 GND.n408 0.152939
R13176 GND.n414 GND.n409 0.152939
R13177 GND.n7751 GND.n414 0.152939
R13178 GND.n67 GND.n40 0.152939
R13179 GND.n68 GND.n67 0.152939
R13180 GND.n69 GND.n68 0.152939
R13181 GND.n87 GND.n69 0.152939
R13182 GND.n88 GND.n87 0.152939
R13183 GND.n89 GND.n88 0.152939
R13184 GND.n90 GND.n89 0.152939
R13185 GND.n108 GND.n90 0.152939
R13186 GND.n109 GND.n108 0.152939
R13187 GND.n110 GND.n109 0.152939
R13188 GND.n111 GND.n110 0.152939
R13189 GND.n129 GND.n111 0.152939
R13190 GND.n130 GND.n129 0.152939
R13191 GND.n131 GND.n130 0.152939
R13192 GND.n132 GND.n131 0.152939
R13193 GND.n150 GND.n132 0.152939
R13194 GND.n151 GND.n150 0.152939
R13195 GND.n8013 GND.n151 0.152939
R13196 GND.n3121 GND.n3027 0.152939
R13197 GND.n4208 GND.n3027 0.152939
R13198 GND.n4209 GND.n4208 0.152939
R13199 GND.n4210 GND.n4209 0.152939
R13200 GND.n4211 GND.n4210 0.152939
R13201 GND.n4211 GND.n3004 0.152939
R13202 GND.n4240 GND.n3004 0.152939
R13203 GND.n4241 GND.n4240 0.152939
R13204 GND.n4242 GND.n4241 0.152939
R13205 GND.n4243 GND.n4242 0.152939
R13206 GND.n4243 GND.n2981 0.152939
R13207 GND.n4272 GND.n2981 0.152939
R13208 GND.n4273 GND.n4272 0.152939
R13209 GND.n4274 GND.n4273 0.152939
R13210 GND.n4275 GND.n4274 0.152939
R13211 GND.n4275 GND.n2958 0.152939
R13212 GND.n4304 GND.n2958 0.152939
R13213 GND.n4305 GND.n4304 0.152939
R13214 GND.n4306 GND.n4305 0.152939
R13215 GND.n4307 GND.n4306 0.152939
R13216 GND.n4307 GND.n2934 0.152939
R13217 GND.n4336 GND.n2934 0.152939
R13218 GND.n4337 GND.n4336 0.152939
R13219 GND.n4338 GND.n4337 0.152939
R13220 GND.n4339 GND.n4338 0.152939
R13221 GND.n4339 GND.n2912 0.152939
R13222 GND.n4368 GND.n2912 0.152939
R13223 GND.n4369 GND.n4368 0.152939
R13224 GND.n4370 GND.n4369 0.152939
R13225 GND.n4371 GND.n4370 0.152939
R13226 GND.n4371 GND.n2889 0.152939
R13227 GND.n4400 GND.n2889 0.152939
R13228 GND.n4401 GND.n4400 0.152939
R13229 GND.n4402 GND.n4401 0.152939
R13230 GND.n4403 GND.n4402 0.152939
R13231 GND.n4403 GND.n2866 0.152939
R13232 GND.n4432 GND.n2866 0.152939
R13233 GND.n4433 GND.n4432 0.152939
R13234 GND.n4434 GND.n4433 0.152939
R13235 GND.n4435 GND.n4434 0.152939
R13236 GND.n4435 GND.n2843 0.152939
R13237 GND.n4464 GND.n2843 0.152939
R13238 GND.n4465 GND.n4464 0.152939
R13239 GND.n4466 GND.n4465 0.152939
R13240 GND.n4467 GND.n4466 0.152939
R13241 GND.n4467 GND.n2820 0.152939
R13242 GND.n4496 GND.n2820 0.152939
R13243 GND.n4497 GND.n4496 0.152939
R13244 GND.n4498 GND.n4497 0.152939
R13245 GND.n4499 GND.n4498 0.152939
R13246 GND.n4499 GND.n2797 0.152939
R13247 GND.n4528 GND.n2797 0.152939
R13248 GND.n4529 GND.n4528 0.152939
R13249 GND.n4530 GND.n4529 0.152939
R13250 GND.n4531 GND.n4530 0.152939
R13251 GND.n4533 GND.n4531 0.152939
R13252 GND.n4533 GND.n4532 0.152939
R13253 GND.n4532 GND.n2773 0.152939
R13254 GND.n4656 GND.n2773 0.152939
R13255 GND.n4657 GND.n4656 0.152939
R13256 GND.n4658 GND.n4657 0.152939
R13257 GND.n4659 GND.n4658 0.152939
R13258 GND.n4660 GND.n4659 0.152939
R13259 GND.n4660 GND.n2762 0.152939
R13260 GND.n4694 GND.n2762 0.152939
R13261 GND.n4695 GND.n4694 0.152939
R13262 GND.n4696 GND.n4695 0.152939
R13263 GND.n4697 GND.n4696 0.152939
R13264 GND.n4698 GND.n4697 0.152939
R13265 GND.n4701 GND.n4698 0.152939
R13266 GND.n4702 GND.n4701 0.152939
R13267 GND.n4704 GND.n4702 0.152939
R13268 GND.n4704 GND.n4703 0.152939
R13269 GND.n4703 GND.n2749 0.152939
R13270 GND.n4767 GND.n2749 0.152939
R13271 GND.n4768 GND.n4767 0.152939
R13272 GND.n4769 GND.n4768 0.152939
R13273 GND.n4769 GND.n2745 0.152939
R13274 GND.n4775 GND.n2745 0.152939
R13275 GND.n4776 GND.n4775 0.152939
R13276 GND.n4777 GND.n4776 0.152939
R13277 GND.n4778 GND.n4777 0.152939
R13278 GND.n4779 GND.n4778 0.152939
R13279 GND.n4780 GND.n4779 0.152939
R13280 GND.n4781 GND.n4780 0.152939
R13281 GND.n4781 GND.n2726 0.152939
R13282 GND.n4860 GND.n2726 0.152939
R13283 GND.n4861 GND.n4860 0.152939
R13284 GND.n4862 GND.n4861 0.152939
R13285 GND.n4864 GND.n4862 0.152939
R13286 GND.n4864 GND.n4863 0.152939
R13287 GND.n4863 GND.n2709 0.152939
R13288 GND.n4883 GND.n2709 0.152939
R13289 GND.n4884 GND.n4883 0.152939
R13290 GND.n4885 GND.n4884 0.152939
R13291 GND.n4885 GND.n2705 0.152939
R13292 GND.n4892 GND.n2705 0.152939
R13293 GND.n4893 GND.n4892 0.152939
R13294 GND.n4894 GND.n4893 0.152939
R13295 GND.n4894 GND.n2703 0.152939
R13296 GND.n4900 GND.n2703 0.152939
R13297 GND.n4901 GND.n4900 0.152939
R13298 GND.n4902 GND.n4901 0.152939
R13299 GND.n4902 GND.n2701 0.152939
R13300 GND.n4910 GND.n2701 0.152939
R13301 GND.n4911 GND.n4910 0.152939
R13302 GND.n4912 GND.n4911 0.152939
R13303 GND.n4912 GND.n2699 0.152939
R13304 GND.n4918 GND.n2699 0.152939
R13305 GND.n4919 GND.n4918 0.152939
R13306 GND.n4920 GND.n4919 0.152939
R13307 GND.n4920 GND.n2697 0.152939
R13308 GND.n4928 GND.n2697 0.152939
R13309 GND.n4929 GND.n4928 0.152939
R13310 GND.n4930 GND.n4929 0.152939
R13311 GND.n4930 GND.n2695 0.152939
R13312 GND.n4936 GND.n2695 0.152939
R13313 GND.n4937 GND.n4936 0.152939
R13314 GND.n4938 GND.n4937 0.152939
R13315 GND.n4938 GND.n2690 0.152939
R13316 GND.n4944 GND.n2690 0.152939
R13317 GND.n4945 GND.n4944 0.152939
R13318 GND.n4946 GND.n4945 0.152939
R13319 GND.n4946 GND.n2688 0.152939
R13320 GND.n4954 GND.n2688 0.152939
R13321 GND.n4955 GND.n4954 0.152939
R13322 GND.n4956 GND.n4955 0.152939
R13323 GND.n4956 GND.n2686 0.152939
R13324 GND.n4962 GND.n2686 0.152939
R13325 GND.n4963 GND.n4962 0.152939
R13326 GND.n4964 GND.n4963 0.152939
R13327 GND.n4964 GND.n2684 0.152939
R13328 GND.n4972 GND.n2684 0.152939
R13329 GND.n4973 GND.n4972 0.152939
R13330 GND.n4974 GND.n4973 0.152939
R13331 GND.n4974 GND.n2682 0.152939
R13332 GND.n4980 GND.n2682 0.152939
R13333 GND.n4981 GND.n4980 0.152939
R13334 GND.n4982 GND.n4981 0.152939
R13335 GND.n4982 GND.n2678 0.152939
R13336 GND.n4988 GND.n2678 0.152939
R13337 GND.n4989 GND.n4988 0.152939
R13338 GND.n4990 GND.n4989 0.152939
R13339 GND.n4990 GND.n2676 0.152939
R13340 GND.n4998 GND.n2676 0.152939
R13341 GND.n4999 GND.n4998 0.152939
R13342 GND.n5000 GND.n4999 0.152939
R13343 GND.n5000 GND.n2674 0.152939
R13344 GND.n5007 GND.n2674 0.152939
R13345 GND.n5008 GND.n5007 0.152939
R13346 GND.n5009 GND.n5008 0.152939
R13347 GND.n5009 GND.n2672 0.152939
R13348 GND.n5017 GND.n2672 0.152939
R13349 GND.n5018 GND.n5017 0.152939
R13350 GND.n5019 GND.n5018 0.152939
R13351 GND.n5019 GND.n2667 0.152939
R13352 GND.n3061 GND.n3035 0.152939
R13353 GND.n3062 GND.n3061 0.152939
R13354 GND.n3063 GND.n3062 0.152939
R13355 GND.n3064 GND.n3063 0.152939
R13356 GND.n3065 GND.n3064 0.152939
R13357 GND.n3066 GND.n3065 0.152939
R13358 GND.n3067 GND.n3066 0.152939
R13359 GND.n3068 GND.n3067 0.152939
R13360 GND.n3069 GND.n3068 0.152939
R13361 GND.n3070 GND.n3069 0.152939
R13362 GND.n4160 GND.n3070 0.152939
R13363 GND.n4199 GND.n4198 0.152939
R13364 GND.n4200 GND.n4199 0.152939
R13365 GND.n4201 GND.n4200 0.152939
R13366 GND.n4201 GND.n3012 0.152939
R13367 GND.n4230 GND.n3012 0.152939
R13368 GND.n4231 GND.n4230 0.152939
R13369 GND.n4232 GND.n4231 0.152939
R13370 GND.n4233 GND.n4232 0.152939
R13371 GND.n4233 GND.n2989 0.152939
R13372 GND.n4262 GND.n2989 0.152939
R13373 GND.n4263 GND.n4262 0.152939
R13374 GND.n4264 GND.n4263 0.152939
R13375 GND.n4265 GND.n4264 0.152939
R13376 GND.n4265 GND.n2966 0.152939
R13377 GND.n4294 GND.n2966 0.152939
R13378 GND.n4295 GND.n4294 0.152939
R13379 GND.n4296 GND.n4295 0.152939
R13380 GND.n4297 GND.n4296 0.152939
R13381 GND.n4297 GND.n2943 0.152939
R13382 GND.n4326 GND.n2943 0.152939
R13383 GND.n4327 GND.n4326 0.152939
R13384 GND.n4328 GND.n4327 0.152939
R13385 GND.n4329 GND.n4328 0.152939
R13386 GND.n4329 GND.n2920 0.152939
R13387 GND.n4358 GND.n2920 0.152939
R13388 GND.n4359 GND.n4358 0.152939
R13389 GND.n4360 GND.n4359 0.152939
R13390 GND.n4361 GND.n4360 0.152939
R13391 GND.n4361 GND.n2897 0.152939
R13392 GND.n4390 GND.n2897 0.152939
R13393 GND.n4391 GND.n4390 0.152939
R13394 GND.n4392 GND.n4391 0.152939
R13395 GND.n4393 GND.n4392 0.152939
R13396 GND.n4393 GND.n2874 0.152939
R13397 GND.n4422 GND.n2874 0.152939
R13398 GND.n4423 GND.n4422 0.152939
R13399 GND.n4424 GND.n4423 0.152939
R13400 GND.n4425 GND.n4424 0.152939
R13401 GND.n4425 GND.n2851 0.152939
R13402 GND.n4454 GND.n2851 0.152939
R13403 GND.n4455 GND.n4454 0.152939
R13404 GND.n4456 GND.n4455 0.152939
R13405 GND.n4457 GND.n4456 0.152939
R13406 GND.n4457 GND.n2828 0.152939
R13407 GND.n4486 GND.n2828 0.152939
R13408 GND.n4487 GND.n4486 0.152939
R13409 GND.n4488 GND.n4487 0.152939
R13410 GND.n4489 GND.n4488 0.152939
R13411 GND.n4489 GND.n2805 0.152939
R13412 GND.n4518 GND.n2805 0.152939
R13413 GND.n4519 GND.n4518 0.152939
R13414 GND.n4520 GND.n4519 0.152939
R13415 GND.n4521 GND.n4520 0.152939
R13416 GND.n4521 GND.n2782 0.152939
R13417 GND.n4569 GND.n2782 0.152939
R13418 GND.n4570 GND.n4569 0.152939
R13419 GND.n4571 GND.n4570 0.152939
R13420 GND.n4573 GND.n4571 0.152939
R13421 GND.n4573 GND.n4572 0.152939
R13422 GND.n4572 GND.n1656 0.152939
R13423 GND.n1657 GND.n1656 0.152939
R13424 GND.n1658 GND.n1657 0.152939
R13425 GND.n1686 GND.n1658 0.152939
R13426 GND.n1689 GND.n1686 0.152939
R13427 GND.n1690 GND.n1689 0.152939
R13428 GND.n1691 GND.n1690 0.152939
R13429 GND.n1692 GND.n1691 0.152939
R13430 GND.n1693 GND.n1692 0.152939
R13431 GND.n1735 GND.n1693 0.152939
R13432 GND.n1736 GND.n1735 0.152939
R13433 GND.n1741 GND.n1736 0.152939
R13434 GND.n1742 GND.n1741 0.152939
R13435 GND.n1743 GND.n1742 0.152939
R13436 GND.n1744 GND.n1743 0.152939
R13437 GND.n1745 GND.n1744 0.152939
R13438 GND.n4794 GND.n1745 0.152939
R13439 GND.n4795 GND.n4794 0.152939
R13440 GND.n4795 GND.n4792 0.152939
R13441 GND.n4801 GND.n4792 0.152939
R13442 GND.n4802 GND.n4801 0.152939
R13443 GND.n4803 GND.n4802 0.152939
R13444 GND.n4804 GND.n4803 0.152939
R13445 GND.n4804 GND.n2733 0.152939
R13446 GND.n4849 GND.n2733 0.152939
R13447 GND.n4850 GND.n4849 0.152939
R13448 GND.n4851 GND.n4850 0.152939
R13449 GND.n4852 GND.n4851 0.152939
R13450 GND.n4852 GND.n2716 0.152939
R13451 GND.n4871 GND.n2716 0.152939
R13452 GND.n4872 GND.n4871 0.152939
R13453 GND.n4874 GND.n4872 0.152939
R13454 GND.n4874 GND.n4873 0.152939
R13455 GND.n4873 GND.n1901 0.152939
R13456 GND.n1902 GND.n1901 0.152939
R13457 GND.n1903 GND.n1902 0.152939
R13458 GND.n1906 GND.n1903 0.152939
R13459 GND.n1907 GND.n1906 0.152939
R13460 GND.n1908 GND.n1907 0.152939
R13461 GND.n1909 GND.n1908 0.152939
R13462 GND.n1929 GND.n1909 0.152939
R13463 GND.n1930 GND.n1929 0.152939
R13464 GND.n1931 GND.n1930 0.152939
R13465 GND.n1932 GND.n1931 0.152939
R13466 GND.n1933 GND.n1932 0.152939
R13467 GND.n1956 GND.n1933 0.152939
R13468 GND.n1957 GND.n1956 0.152939
R13469 GND.n1958 GND.n1957 0.152939
R13470 GND.n1959 GND.n1958 0.152939
R13471 GND.n1960 GND.n1959 0.152939
R13472 GND.n1983 GND.n1960 0.152939
R13473 GND.n1984 GND.n1983 0.152939
R13474 GND.n1985 GND.n1984 0.152939
R13475 GND.n1986 GND.n1985 0.152939
R13476 GND.n1987 GND.n1986 0.152939
R13477 GND.n2009 GND.n1987 0.152939
R13478 GND.n2010 GND.n2009 0.152939
R13479 GND.n2011 GND.n2010 0.152939
R13480 GND.n2012 GND.n2011 0.152939
R13481 GND.n2013 GND.n2012 0.152939
R13482 GND.n2036 GND.n2013 0.152939
R13483 GND.n2037 GND.n2036 0.152939
R13484 GND.n2038 GND.n2037 0.152939
R13485 GND.n2039 GND.n2038 0.152939
R13486 GND.n2040 GND.n2039 0.152939
R13487 GND.n2063 GND.n2040 0.152939
R13488 GND.n2064 GND.n2063 0.152939
R13489 GND.n2065 GND.n2064 0.152939
R13490 GND.n2066 GND.n2065 0.152939
R13491 GND.n2067 GND.n2066 0.152939
R13492 GND.n2090 GND.n2067 0.152939
R13493 GND.n2091 GND.n2090 0.152939
R13494 GND.n2092 GND.n2091 0.152939
R13495 GND.n2093 GND.n2092 0.152939
R13496 GND.n2094 GND.n2093 0.152939
R13497 GND.n2117 GND.n2094 0.152939
R13498 GND.n2118 GND.n2117 0.152939
R13499 GND.n2119 GND.n2118 0.152939
R13500 GND.n2120 GND.n2119 0.152939
R13501 GND.n2121 GND.n2120 0.152939
R13502 GND.n2144 GND.n2121 0.152939
R13503 GND.n2145 GND.n2144 0.152939
R13504 GND.n2146 GND.n2145 0.152939
R13505 GND.n2147 GND.n2146 0.152939
R13506 GND.n2148 GND.n2147 0.152939
R13507 GND.n2171 GND.n2148 0.152939
R13508 GND.n2172 GND.n2171 0.152939
R13509 GND.n2173 GND.n2172 0.152939
R13510 GND.n2174 GND.n2173 0.152939
R13511 GND.n2175 GND.n2174 0.152939
R13512 GND.n2197 GND.n2175 0.152939
R13513 GND.n2198 GND.n2197 0.152939
R13514 GND.n2199 GND.n2198 0.152939
R13515 GND.n2200 GND.n2199 0.152939
R13516 GND.n2201 GND.n2200 0.152939
R13517 GND.n2235 GND.n2201 0.152939
R13518 GND.n2237 GND.n2235 0.152939
R13519 GND.n5639 GND.n2238 0.152939
R13520 GND.n5639 GND.n5638 0.152939
R13521 GND.n5638 GND.n5637 0.152939
R13522 GND.n5637 GND.n2240 0.152939
R13523 GND.n2241 GND.n2240 0.152939
R13524 GND.n2242 GND.n2241 0.152939
R13525 GND.n2243 GND.n2242 0.152939
R13526 GND.n2244 GND.n2243 0.152939
R13527 GND.n2245 GND.n2244 0.152939
R13528 GND.n2246 GND.n2245 0.152939
R13529 GND.n2247 GND.n2246 0.152939
R13530 GND.n5044 GND.n2660 0.152939
R13531 GND.n5053 GND.n2660 0.152939
R13532 GND.n5054 GND.n5053 0.152939
R13533 GND.n5055 GND.n5054 0.152939
R13534 GND.n5055 GND.n2576 0.152939
R13535 GND.n5068 GND.n2576 0.152939
R13536 GND.n5069 GND.n5068 0.152939
R13537 GND.n5070 GND.n5069 0.152939
R13538 GND.n5070 GND.n2572 0.152939
R13539 GND.n5083 GND.n2572 0.152939
R13540 GND.n5084 GND.n5083 0.152939
R13541 GND.n5085 GND.n5084 0.152939
R13542 GND.n5085 GND.n2568 0.152939
R13543 GND.n5098 GND.n2568 0.152939
R13544 GND.n5099 GND.n5098 0.152939
R13545 GND.n5100 GND.n5099 0.152939
R13546 GND.n5100 GND.n2564 0.152939
R13547 GND.n5113 GND.n2564 0.152939
R13548 GND.n5114 GND.n5113 0.152939
R13549 GND.n5115 GND.n5114 0.152939
R13550 GND.n5116 GND.n5115 0.152939
R13551 GND.n5117 GND.n5116 0.152939
R13552 GND.n5117 GND.n26 0.152939
R13553 GND.n8081 GND.n27 0.152939
R13554 GND.n5138 GND.n27 0.152939
R13555 GND.n5139 GND.n5138 0.152939
R13556 GND.n5140 GND.n5139 0.152939
R13557 GND.n5141 GND.n5140 0.152939
R13558 GND.n5205 GND.n5141 0.152939
R13559 GND.n5206 GND.n5205 0.152939
R13560 GND.n5207 GND.n5206 0.152939
R13561 GND.n5208 GND.n5207 0.152939
R13562 GND.n5212 GND.n5208 0.152939
R13563 GND.n5213 GND.n5212 0.152939
R13564 GND.n5214 GND.n5213 0.152939
R13565 GND.n5215 GND.n5214 0.152939
R13566 GND.n5219 GND.n5215 0.152939
R13567 GND.n5220 GND.n5219 0.152939
R13568 GND.n5221 GND.n5220 0.152939
R13569 GND.n5222 GND.n5221 0.152939
R13570 GND.n5226 GND.n5222 0.152939
R13571 GND.n5227 GND.n5226 0.152939
R13572 GND.n5228 GND.n5227 0.152939
R13573 GND.n5229 GND.n5228 0.152939
R13574 GND.n5230 GND.n5229 0.152939
R13575 GND.n5295 GND.n5230 0.152939
R13576 GND.n5255 GND.n286 0.152939
R13577 GND.n5256 GND.n5255 0.152939
R13578 GND.n5257 GND.n5256 0.152939
R13579 GND.n5257 GND.n5245 0.152939
R13580 GND.n5265 GND.n5245 0.152939
R13581 GND.n5266 GND.n5265 0.152939
R13582 GND.n5267 GND.n5266 0.152939
R13583 GND.n5267 GND.n5241 0.152939
R13584 GND.n5275 GND.n5241 0.152939
R13585 GND.n5276 GND.n5275 0.152939
R13586 GND.n5277 GND.n5276 0.152939
R13587 GND.n5277 GND.n5237 0.152939
R13588 GND.n5285 GND.n5237 0.152939
R13589 GND.n5286 GND.n5285 0.152939
R13590 GND.n5287 GND.n5286 0.152939
R13591 GND.n5287 GND.n5231 0.152939
R13592 GND.n5294 GND.n5231 0.152939
R13593 GND.n8012 GND.n152 0.152939
R13594 GND.n157 GND.n152 0.152939
R13595 GND.n158 GND.n157 0.152939
R13596 GND.n159 GND.n158 0.152939
R13597 GND.n160 GND.n159 0.152939
R13598 GND.n164 GND.n160 0.152939
R13599 GND.n165 GND.n164 0.152939
R13600 GND.n166 GND.n165 0.152939
R13601 GND.n167 GND.n166 0.152939
R13602 GND.n171 GND.n167 0.152939
R13603 GND.n172 GND.n171 0.152939
R13604 GND.n173 GND.n172 0.152939
R13605 GND.n174 GND.n173 0.152939
R13606 GND.n178 GND.n174 0.152939
R13607 GND.n179 GND.n178 0.152939
R13608 GND.n7981 GND.n179 0.152939
R13609 GND.n7981 GND.n7980 0.152939
R13610 GND.n7980 GND.n7979 0.152939
R13611 GND.n7979 GND.n183 0.152939
R13612 GND.n189 GND.n183 0.152939
R13613 GND.n190 GND.n189 0.152939
R13614 GND.n191 GND.n190 0.152939
R13615 GND.n192 GND.n191 0.152939
R13616 GND.n196 GND.n192 0.152939
R13617 GND.n197 GND.n196 0.152939
R13618 GND.n198 GND.n197 0.152939
R13619 GND.n199 GND.n198 0.152939
R13620 GND.n203 GND.n199 0.152939
R13621 GND.n204 GND.n203 0.152939
R13622 GND.n205 GND.n204 0.152939
R13623 GND.n206 GND.n205 0.152939
R13624 GND.n210 GND.n206 0.152939
R13625 GND.n211 GND.n210 0.152939
R13626 GND.n212 GND.n211 0.152939
R13627 GND.n7947 GND.n212 0.152939
R13628 GND.n7947 GND.n7946 0.152939
R13629 GND.n7946 GND.n7945 0.152939
R13630 GND.n7945 GND.n218 0.152939
R13631 GND.n223 GND.n218 0.152939
R13632 GND.n224 GND.n223 0.152939
R13633 GND.n225 GND.n224 0.152939
R13634 GND.n229 GND.n225 0.152939
R13635 GND.n230 GND.n229 0.152939
R13636 GND.n231 GND.n230 0.152939
R13637 GND.n232 GND.n231 0.152939
R13638 GND.n236 GND.n232 0.152939
R13639 GND.n237 GND.n236 0.152939
R13640 GND.n238 GND.n237 0.152939
R13641 GND.n239 GND.n238 0.152939
R13642 GND.n243 GND.n239 0.152939
R13643 GND.n244 GND.n243 0.152939
R13644 GND.n245 GND.n244 0.152939
R13645 GND.n246 GND.n245 0.152939
R13646 GND.n253 GND.n246 0.152939
R13647 GND.n254 GND.n253 0.152939
R13648 GND.n255 GND.n254 0.152939
R13649 GND.n256 GND.n255 0.152939
R13650 GND.n260 GND.n256 0.152939
R13651 GND.n261 GND.n260 0.152939
R13652 GND.n262 GND.n261 0.152939
R13653 GND.n263 GND.n262 0.152939
R13654 GND.n267 GND.n263 0.152939
R13655 GND.n268 GND.n267 0.152939
R13656 GND.n269 GND.n268 0.152939
R13657 GND.n270 GND.n269 0.152939
R13658 GND.n274 GND.n270 0.152939
R13659 GND.n275 GND.n274 0.152939
R13660 GND.n276 GND.n275 0.152939
R13661 GND.n277 GND.n276 0.152939
R13662 GND.n281 GND.n277 0.152939
R13663 GND.n282 GND.n281 0.152939
R13664 GND.n7881 GND.n282 0.152939
R13665 GND.n7881 GND.n7880 0.152939
R13666 GND.n2318 GND.n2317 0.152939
R13667 GND.n2319 GND.n2318 0.152939
R13668 GND.n2320 GND.n2319 0.152939
R13669 GND.n2321 GND.n2320 0.152939
R13670 GND.n2322 GND.n2321 0.152939
R13671 GND.n2323 GND.n2322 0.152939
R13672 GND.n2324 GND.n2323 0.152939
R13673 GND.n2325 GND.n2324 0.152939
R13674 GND.n2326 GND.n2325 0.152939
R13675 GND.n2327 GND.n2326 0.152939
R13676 GND.n2328 GND.n2327 0.152939
R13677 GND.n2329 GND.n2328 0.152939
R13678 GND.n2330 GND.n2329 0.152939
R13679 GND.n2331 GND.n2330 0.152939
R13680 GND.n2332 GND.n2331 0.152939
R13681 GND.n2334 GND.n2332 0.152939
R13682 GND.n2337 GND.n2334 0.152939
R13683 GND.n2338 GND.n2337 0.152939
R13684 GND.n2339 GND.n2338 0.152939
R13685 GND.n2340 GND.n2339 0.152939
R13686 GND.n2341 GND.n2340 0.152939
R13687 GND.n2342 GND.n2341 0.152939
R13688 GND.n2343 GND.n2342 0.152939
R13689 GND.n2344 GND.n2343 0.152939
R13690 GND.n2345 GND.n2344 0.152939
R13691 GND.n2346 GND.n2345 0.152939
R13692 GND.n2347 GND.n2346 0.152939
R13693 GND.n2348 GND.n2347 0.152939
R13694 GND.n2349 GND.n2348 0.152939
R13695 GND.n2350 GND.n2349 0.152939
R13696 GND.n2351 GND.n2350 0.152939
R13697 GND.n2352 GND.n2351 0.152939
R13698 GND.n2353 GND.n2352 0.152939
R13699 GND.n2359 GND.n2358 0.152939
R13700 GND.n2360 GND.n2359 0.152939
R13701 GND.n2361 GND.n2360 0.152939
R13702 GND.n2362 GND.n2361 0.152939
R13703 GND.n2363 GND.n2362 0.152939
R13704 GND.n2364 GND.n2363 0.152939
R13705 GND.n2365 GND.n2364 0.152939
R13706 GND.n2366 GND.n2365 0.152939
R13707 GND.n2367 GND.n2366 0.152939
R13708 GND.n2368 GND.n2367 0.152939
R13709 GND.n2369 GND.n2368 0.152939
R13710 GND.n2370 GND.n2369 0.152939
R13711 GND.n2371 GND.n2370 0.152939
R13712 GND.n2372 GND.n2371 0.152939
R13713 GND.n2373 GND.n2372 0.152939
R13714 GND.n2374 GND.n2373 0.152939
R13715 GND.n2375 GND.n2374 0.152939
R13716 GND.n2378 GND.n2375 0.152939
R13717 GND.n2379 GND.n2378 0.152939
R13718 GND.n2380 GND.n2379 0.152939
R13719 GND.n2381 GND.n2380 0.152939
R13720 GND.n2382 GND.n2381 0.152939
R13721 GND.n2383 GND.n2382 0.152939
R13722 GND.n2384 GND.n2383 0.152939
R13723 GND.n2385 GND.n2384 0.152939
R13724 GND.n2386 GND.n2385 0.152939
R13725 GND.n2387 GND.n2386 0.152939
R13726 GND.n2388 GND.n2387 0.152939
R13727 GND.n2389 GND.n2388 0.152939
R13728 GND.n2390 GND.n2389 0.152939
R13729 GND.n2391 GND.n2390 0.152939
R13730 GND.n2392 GND.n2391 0.152939
R13731 GND.n2393 GND.n2392 0.152939
R13732 GND.n2394 GND.n2393 0.152939
R13733 GND.n5447 GND.n2394 0.152939
R13734 GND.n5447 GND.n5446 0.152939
R13735 GND.n5446 GND.n5445 0.152939
R13736 GND.n2441 GND.n2440 0.152939
R13737 GND.n2442 GND.n2441 0.152939
R13738 GND.n2443 GND.n2442 0.152939
R13739 GND.n2461 GND.n2443 0.152939
R13740 GND.n2462 GND.n2461 0.152939
R13741 GND.n2463 GND.n2462 0.152939
R13742 GND.n2464 GND.n2463 0.152939
R13743 GND.n2482 GND.n2464 0.152939
R13744 GND.n2483 GND.n2482 0.152939
R13745 GND.n2484 GND.n2483 0.152939
R13746 GND.n2485 GND.n2484 0.152939
R13747 GND.n2503 GND.n2485 0.152939
R13748 GND.n2504 GND.n2503 0.152939
R13749 GND.n2505 GND.n2504 0.152939
R13750 GND.n2506 GND.n2505 0.152939
R13751 GND.n2524 GND.n2506 0.152939
R13752 GND.n2525 GND.n2524 0.152939
R13753 GND.n2525 GND.n41 0.152939
R13754 GND.n4027 GND.n3371 0.152939
R13755 GND.n4028 GND.n4027 0.152939
R13756 GND.n4029 GND.n4028 0.152939
R13757 GND.n4030 GND.n4029 0.152939
R13758 GND.n4030 GND.n3342 0.152939
R13759 GND.n4064 GND.n3342 0.152939
R13760 GND.n4065 GND.n4064 0.152939
R13761 GND.n4066 GND.n4065 0.152939
R13762 GND.n4067 GND.n4066 0.152939
R13763 GND.n4067 GND.n3313 0.152939
R13764 GND.n4101 GND.n3313 0.152939
R13765 GND.n4102 GND.n4101 0.152939
R13766 GND.n4103 GND.n4102 0.152939
R13767 GND.n4104 GND.n4103 0.152939
R13768 GND.n4105 GND.n4104 0.152939
R13769 GND.n4108 GND.n4105 0.152939
R13770 GND.n4109 GND.n4108 0.152939
R13771 GND.n4110 GND.n4109 0.152939
R13772 GND.n4111 GND.n4110 0.152939
R13773 GND.n4113 GND.n4111 0.152939
R13774 GND.n4114 GND.n4113 0.152939
R13775 GND.n4114 GND.n3043 0.152939
R13776 GND.n4187 GND.n3043 0.152939
R13777 GND.n4188 GND.n4187 0.152939
R13778 GND.n4189 GND.n4188 0.152939
R13779 GND.n4190 GND.n4189 0.152939
R13780 GND.n4190 GND.n3021 0.152939
R13781 GND.n4219 GND.n3021 0.152939
R13782 GND.n4220 GND.n4219 0.152939
R13783 GND.n4221 GND.n4220 0.152939
R13784 GND.n4222 GND.n4221 0.152939
R13785 GND.n4222 GND.n2998 0.152939
R13786 GND.n4251 GND.n2998 0.152939
R13787 GND.n4252 GND.n4251 0.152939
R13788 GND.n4253 GND.n4252 0.152939
R13789 GND.n4254 GND.n4253 0.152939
R13790 GND.n4254 GND.n2975 0.152939
R13791 GND.n4283 GND.n2975 0.152939
R13792 GND.n4284 GND.n4283 0.152939
R13793 GND.n4285 GND.n4284 0.152939
R13794 GND.n4286 GND.n4285 0.152939
R13795 GND.n4286 GND.n2952 0.152939
R13796 GND.n4315 GND.n2952 0.152939
R13797 GND.n4316 GND.n4315 0.152939
R13798 GND.n4317 GND.n4316 0.152939
R13799 GND.n4318 GND.n4317 0.152939
R13800 GND.n4318 GND.n2929 0.152939
R13801 GND.n4347 GND.n2929 0.152939
R13802 GND.n4348 GND.n4347 0.152939
R13803 GND.n4349 GND.n4348 0.152939
R13804 GND.n4350 GND.n4349 0.152939
R13805 GND.n4350 GND.n2906 0.152939
R13806 GND.n4379 GND.n2906 0.152939
R13807 GND.n4380 GND.n4379 0.152939
R13808 GND.n4381 GND.n4380 0.152939
R13809 GND.n4382 GND.n4381 0.152939
R13810 GND.n4382 GND.n2883 0.152939
R13811 GND.n4411 GND.n2883 0.152939
R13812 GND.n4412 GND.n4411 0.152939
R13813 GND.n4413 GND.n4412 0.152939
R13814 GND.n4414 GND.n4413 0.152939
R13815 GND.n4414 GND.n2860 0.152939
R13816 GND.n4443 GND.n2860 0.152939
R13817 GND.n4444 GND.n4443 0.152939
R13818 GND.n4445 GND.n4444 0.152939
R13819 GND.n4446 GND.n4445 0.152939
R13820 GND.n4446 GND.n2837 0.152939
R13821 GND.n4475 GND.n2837 0.152939
R13822 GND.n4476 GND.n4475 0.152939
R13823 GND.n4477 GND.n4476 0.152939
R13824 GND.n4478 GND.n4477 0.152939
R13825 GND.n4478 GND.n2814 0.152939
R13826 GND.n4507 GND.n2814 0.152939
R13827 GND.n4508 GND.n4507 0.152939
R13828 GND.n4509 GND.n4508 0.152939
R13829 GND.n4510 GND.n4509 0.152939
R13830 GND.n4510 GND.n2791 0.152939
R13831 GND.n4542 GND.n2791 0.152939
R13832 GND.n4543 GND.n4542 0.152939
R13833 GND.n4544 GND.n4543 0.152939
R13834 GND.n4545 GND.n4544 0.152939
R13835 GND.n4546 GND.n4545 0.152939
R13836 GND.n4549 GND.n4546 0.152939
R13837 GND.n4550 GND.n4549 0.152939
R13838 GND.n4551 GND.n4550 0.152939
R13839 GND.n4553 GND.n4551 0.152939
R13840 GND.n4553 GND.n4552 0.152939
R13841 GND.n4552 GND.n1675 0.152939
R13842 GND.n1676 GND.n1675 0.152939
R13843 GND.n1677 GND.n1676 0.152939
R13844 GND.n1710 GND.n1677 0.152939
R13845 GND.n1713 GND.n1710 0.152939
R13846 GND.n1714 GND.n1713 0.152939
R13847 GND.n1715 GND.n1714 0.152939
R13848 GND.n1716 GND.n1715 0.152939
R13849 GND.n1717 GND.n1716 0.152939
R13850 GND.n1754 GND.n1717 0.152939
R13851 GND.n1757 GND.n1754 0.152939
R13852 GND.n1758 GND.n1757 0.152939
R13853 GND.n1759 GND.n1758 0.152939
R13854 GND.n1760 GND.n1759 0.152939
R13855 GND.n1761 GND.n1760 0.152939
R13856 GND.n1776 GND.n1761 0.152939
R13857 GND.n1777 GND.n1776 0.152939
R13858 GND.n1778 GND.n1777 0.152939
R13859 GND.n1779 GND.n1778 0.152939
R13860 GND.n1794 GND.n1779 0.152939
R13861 GND.n1795 GND.n1794 0.152939
R13862 GND.n1796 GND.n1795 0.152939
R13863 GND.n1797 GND.n1796 0.152939
R13864 GND.n1811 GND.n1797 0.152939
R13865 GND.n1812 GND.n1811 0.152939
R13866 GND.n1813 GND.n1812 0.152939
R13867 GND.n1814 GND.n1813 0.152939
R13868 GND.n1828 GND.n1814 0.152939
R13869 GND.n1829 GND.n1828 0.152939
R13870 GND.n1830 GND.n1829 0.152939
R13871 GND.n1831 GND.n1830 0.152939
R13872 GND.n1846 GND.n1831 0.152939
R13873 GND.n1847 GND.n1846 0.152939
R13874 GND.n1848 GND.n1847 0.152939
R13875 GND.n1849 GND.n1848 0.152939
R13876 GND.n1916 GND.n1849 0.152939
R13877 GND.n1917 GND.n1916 0.152939
R13878 GND.n1918 GND.n1917 0.152939
R13879 GND.n1919 GND.n1918 0.152939
R13880 GND.n1942 GND.n1919 0.152939
R13881 GND.n1943 GND.n1942 0.152939
R13882 GND.n1944 GND.n1943 0.152939
R13883 GND.n1945 GND.n1944 0.152939
R13884 GND.n1946 GND.n1945 0.152939
R13885 GND.n1969 GND.n1946 0.152939
R13886 GND.n1970 GND.n1969 0.152939
R13887 GND.n1971 GND.n1970 0.152939
R13888 GND.n1972 GND.n1971 0.152939
R13889 GND.n1973 GND.n1972 0.152939
R13890 GND.n1996 GND.n1973 0.152939
R13891 GND.n1997 GND.n1996 0.152939
R13892 GND.n1998 GND.n1997 0.152939
R13893 GND.n1999 GND.n1998 0.152939
R13894 GND.n2000 GND.n1999 0.152939
R13895 GND.n2022 GND.n2000 0.152939
R13896 GND.n2023 GND.n2022 0.152939
R13897 GND.n2024 GND.n2023 0.152939
R13898 GND.n2025 GND.n2024 0.152939
R13899 GND.n2026 GND.n2025 0.152939
R13900 GND.n2049 GND.n2026 0.152939
R13901 GND.n2050 GND.n2049 0.152939
R13902 GND.n2051 GND.n2050 0.152939
R13903 GND.n2052 GND.n2051 0.152939
R13904 GND.n2053 GND.n2052 0.152939
R13905 GND.n2076 GND.n2053 0.152939
R13906 GND.n2077 GND.n2076 0.152939
R13907 GND.n2078 GND.n2077 0.152939
R13908 GND.n2079 GND.n2078 0.152939
R13909 GND.n2080 GND.n2079 0.152939
R13910 GND.n2103 GND.n2080 0.152939
R13911 GND.n2104 GND.n2103 0.152939
R13912 GND.n2105 GND.n2104 0.152939
R13913 GND.n2106 GND.n2105 0.152939
R13914 GND.n2107 GND.n2106 0.152939
R13915 GND.n2130 GND.n2107 0.152939
R13916 GND.n2131 GND.n2130 0.152939
R13917 GND.n2132 GND.n2131 0.152939
R13918 GND.n2133 GND.n2132 0.152939
R13919 GND.n2134 GND.n2133 0.152939
R13920 GND.n2157 GND.n2134 0.152939
R13921 GND.n2158 GND.n2157 0.152939
R13922 GND.n2159 GND.n2158 0.152939
R13923 GND.n2160 GND.n2159 0.152939
R13924 GND.n2161 GND.n2160 0.152939
R13925 GND.n2183 GND.n2161 0.152939
R13926 GND.n2184 GND.n2183 0.152939
R13927 GND.n2185 GND.n2184 0.152939
R13928 GND.n2186 GND.n2185 0.152939
R13929 GND.n2187 GND.n2186 0.152939
R13930 GND.n2210 GND.n2187 0.152939
R13931 GND.n2211 GND.n2210 0.152939
R13932 GND.n2212 GND.n2211 0.152939
R13933 GND.n2213 GND.n2212 0.152939
R13934 GND.n2214 GND.n2213 0.152939
R13935 GND.n2590 GND.n2214 0.152939
R13936 GND.n2593 GND.n2590 0.152939
R13937 GND.n2594 GND.n2593 0.152939
R13938 GND.n2595 GND.n2594 0.152939
R13939 GND.n2595 GND.n2585 0.152939
R13940 GND.n2601 GND.n2585 0.152939
R13941 GND.n2602 GND.n2601 0.152939
R13942 GND.n2603 GND.n2602 0.152939
R13943 GND.n2603 GND.n2581 0.152939
R13944 GND.n2609 GND.n2581 0.152939
R13945 GND.n2610 GND.n2609 0.152939
R13946 GND.n2611 GND.n2610 0.152939
R13947 GND.n2612 GND.n2611 0.152939
R13948 GND.n2613 GND.n2612 0.152939
R13949 GND.n2616 GND.n2613 0.152939
R13950 GND.n2617 GND.n2616 0.152939
R13951 GND.n2618 GND.n2617 0.152939
R13952 GND.n2619 GND.n2618 0.152939
R13953 GND.n2622 GND.n2619 0.152939
R13954 GND.n2623 GND.n2622 0.152939
R13955 GND.n2624 GND.n2623 0.152939
R13956 GND.n2625 GND.n2624 0.152939
R13957 GND.n2628 GND.n2625 0.152939
R13958 GND.n2629 GND.n2628 0.152939
R13959 GND.n4017 GND.n4016 0.152939
R13960 GND.n4018 GND.n4017 0.152939
R13961 GND.n4019 GND.n4018 0.152939
R13962 GND.n4019 GND.n3353 0.152939
R13963 GND.n4053 GND.n3353 0.152939
R13964 GND.n4054 GND.n4053 0.152939
R13965 GND.n4055 GND.n4054 0.152939
R13966 GND.n4056 GND.n4055 0.152939
R13967 GND.n4056 GND.n3323 0.152939
R13968 GND.n4090 GND.n3323 0.152939
R13969 GND.n4091 GND.n4090 0.152939
R13970 GND.n4092 GND.n4091 0.152939
R13971 GND.n4093 GND.n4092 0.152939
R13972 GND.n4093 GND.n3296 0.152939
R13973 GND.n4145 GND.n3296 0.152939
R13974 GND.n4146 GND.n4145 0.152939
R13975 GND.n4147 GND.n4146 0.152939
R13976 GND.n4147 GND.n1516 0.152939
R13977 GND.n3580 GND.n3523 0.152939
R13978 GND.n3581 GND.n3580 0.152939
R13979 GND.n3582 GND.n3581 0.152939
R13980 GND.n3582 GND.n3574 0.152939
R13981 GND.n3590 GND.n3574 0.152939
R13982 GND.n3591 GND.n3590 0.152939
R13983 GND.n3592 GND.n3591 0.152939
R13984 GND.n3592 GND.n3572 0.152939
R13985 GND.n3600 GND.n3572 0.152939
R13986 GND.n3601 GND.n3600 0.152939
R13987 GND.n3602 GND.n3601 0.152939
R13988 GND.n3602 GND.n3570 0.152939
R13989 GND.n3610 GND.n3570 0.152939
R13990 GND.n3611 GND.n3610 0.152939
R13991 GND.n3612 GND.n3611 0.152939
R13992 GND.n3612 GND.n3568 0.152939
R13993 GND.n3622 GND.n3568 0.152939
R13994 GND.n3623 GND.n3622 0.152939
R13995 GND.n3624 GND.n3623 0.152939
R13996 GND.n3624 GND.n3566 0.152939
R13997 GND.n3632 GND.n3566 0.152939
R13998 GND.n3633 GND.n3632 0.152939
R13999 GND.n3634 GND.n3633 0.152939
R14000 GND.n3634 GND.n3564 0.152939
R14001 GND.n3642 GND.n3564 0.152939
R14002 GND.n3643 GND.n3642 0.152939
R14003 GND.n3644 GND.n3643 0.152939
R14004 GND.n3644 GND.n3562 0.152939
R14005 GND.n3652 GND.n3562 0.152939
R14006 GND.n3653 GND.n3652 0.152939
R14007 GND.n3654 GND.n3653 0.152939
R14008 GND.n3654 GND.n3560 0.152939
R14009 GND.n3662 GND.n3560 0.152939
R14010 GND.n3663 GND.n3662 0.152939
R14011 GND.n3664 GND.n3663 0.152939
R14012 GND.n3664 GND.n3558 0.152939
R14013 GND.n3674 GND.n3558 0.152939
R14014 GND.n3675 GND.n3674 0.152939
R14015 GND.n3676 GND.n3675 0.152939
R14016 GND.n3676 GND.n3556 0.152939
R14017 GND.n3684 GND.n3556 0.152939
R14018 GND.n3685 GND.n3684 0.152939
R14019 GND.n3686 GND.n3685 0.152939
R14020 GND.n3686 GND.n3554 0.152939
R14021 GND.n3694 GND.n3554 0.152939
R14022 GND.n3695 GND.n3694 0.152939
R14023 GND.n3696 GND.n3695 0.152939
R14024 GND.n3696 GND.n3552 0.152939
R14025 GND.n3704 GND.n3552 0.152939
R14026 GND.n3705 GND.n3704 0.152939
R14027 GND.n3706 GND.n3705 0.152939
R14028 GND.n3706 GND.n3550 0.152939
R14029 GND.n3717 GND.n3550 0.152939
R14030 GND.n3718 GND.n3717 0.152939
R14031 GND.n3719 GND.n3718 0.152939
R14032 GND.n3719 GND.n3548 0.152939
R14033 GND.n3727 GND.n3548 0.152939
R14034 GND.n3728 GND.n3727 0.152939
R14035 GND.n3729 GND.n3728 0.152939
R14036 GND.n3729 GND.n3546 0.152939
R14037 GND.n3737 GND.n3546 0.152939
R14038 GND.n3738 GND.n3737 0.152939
R14039 GND.n3739 GND.n3738 0.152939
R14040 GND.n3739 GND.n3544 0.152939
R14041 GND.n3747 GND.n3544 0.152939
R14042 GND.n3748 GND.n3747 0.152939
R14043 GND.n3749 GND.n3748 0.152939
R14044 GND.n3749 GND.n3542 0.152939
R14045 GND.n3757 GND.n3542 0.152939
R14046 GND.n3758 GND.n3757 0.152939
R14047 GND.n3759 GND.n3758 0.152939
R14048 GND.n3759 GND.n3536 0.152939
R14049 GND.n3763 GND.n3536 0.152939
R14050 GND.n3783 GND.n3782 0.152939
R14051 GND.n3784 GND.n3783 0.152939
R14052 GND.n3785 GND.n3784 0.152939
R14053 GND.n3785 GND.n3494 0.152939
R14054 GND.n3819 GND.n3494 0.152939
R14055 GND.n3820 GND.n3819 0.152939
R14056 GND.n3821 GND.n3820 0.152939
R14057 GND.n3822 GND.n3821 0.152939
R14058 GND.n3822 GND.n3465 0.152939
R14059 GND.n3856 GND.n3465 0.152939
R14060 GND.n3857 GND.n3856 0.152939
R14061 GND.n3858 GND.n3857 0.152939
R14062 GND.n3859 GND.n3858 0.152939
R14063 GND.n3859 GND.n3436 0.152939
R14064 GND.n3896 GND.n3436 0.152939
R14065 GND.n3897 GND.n3896 0.152939
R14066 GND.n3899 GND.n3897 0.152939
R14067 GND.n3899 GND.n3898 0.152939
R14068 GND.n6499 GND.n1212 0.152939
R14069 GND.n1217 GND.n1212 0.152939
R14070 GND.n1218 GND.n1217 0.152939
R14071 GND.n1219 GND.n1218 0.152939
R14072 GND.n1220 GND.n1219 0.152939
R14073 GND.n1225 GND.n1220 0.152939
R14074 GND.n1226 GND.n1225 0.152939
R14075 GND.n1227 GND.n1226 0.152939
R14076 GND.n1228 GND.n1227 0.152939
R14077 GND.n1233 GND.n1228 0.152939
R14078 GND.n1234 GND.n1233 0.152939
R14079 GND.n1235 GND.n1234 0.152939
R14080 GND.n1236 GND.n1235 0.152939
R14081 GND.n1241 GND.n1236 0.152939
R14082 GND.n1242 GND.n1241 0.152939
R14083 GND.n1243 GND.n1242 0.152939
R14084 GND.n1244 GND.n1243 0.152939
R14085 GND.n1249 GND.n1244 0.152939
R14086 GND.n1250 GND.n1249 0.152939
R14087 GND.n1251 GND.n1250 0.152939
R14088 GND.n1252 GND.n1251 0.152939
R14089 GND.n1257 GND.n1252 0.152939
R14090 GND.n1258 GND.n1257 0.152939
R14091 GND.n1259 GND.n1258 0.152939
R14092 GND.n1260 GND.n1259 0.152939
R14093 GND.n1265 GND.n1260 0.152939
R14094 GND.n1266 GND.n1265 0.152939
R14095 GND.n1267 GND.n1266 0.152939
R14096 GND.n1268 GND.n1267 0.152939
R14097 GND.n1273 GND.n1268 0.152939
R14098 GND.n1274 GND.n1273 0.152939
R14099 GND.n1275 GND.n1274 0.152939
R14100 GND.n1276 GND.n1275 0.152939
R14101 GND.n1281 GND.n1276 0.152939
R14102 GND.n1282 GND.n1281 0.152939
R14103 GND.n1283 GND.n1282 0.152939
R14104 GND.n1284 GND.n1283 0.152939
R14105 GND.n1289 GND.n1284 0.152939
R14106 GND.n1290 GND.n1289 0.152939
R14107 GND.n1291 GND.n1290 0.152939
R14108 GND.n1292 GND.n1291 0.152939
R14109 GND.n1297 GND.n1292 0.152939
R14110 GND.n1298 GND.n1297 0.152939
R14111 GND.n1299 GND.n1298 0.152939
R14112 GND.n1300 GND.n1299 0.152939
R14113 GND.n1305 GND.n1300 0.152939
R14114 GND.n1306 GND.n1305 0.152939
R14115 GND.n1307 GND.n1306 0.152939
R14116 GND.n1308 GND.n1307 0.152939
R14117 GND.n1313 GND.n1308 0.152939
R14118 GND.n1314 GND.n1313 0.152939
R14119 GND.n1315 GND.n1314 0.152939
R14120 GND.n1316 GND.n1315 0.152939
R14121 GND.n1321 GND.n1316 0.152939
R14122 GND.n1322 GND.n1321 0.152939
R14123 GND.n1323 GND.n1322 0.152939
R14124 GND.n1324 GND.n1323 0.152939
R14125 GND.n3527 GND.n1324 0.152939
R14126 GND.n3528 GND.n3527 0.152939
R14127 GND.n3529 GND.n3528 0.152939
R14128 GND.n3529 GND.n3513 0.152939
R14129 GND.n3793 GND.n3513 0.152939
R14130 GND.n3794 GND.n3793 0.152939
R14131 GND.n3795 GND.n3794 0.152939
R14132 GND.n3796 GND.n3795 0.152939
R14133 GND.n3796 GND.n3483 0.152939
R14134 GND.n3830 GND.n3483 0.152939
R14135 GND.n3831 GND.n3830 0.152939
R14136 GND.n3832 GND.n3831 0.152939
R14137 GND.n3833 GND.n3832 0.152939
R14138 GND.n3833 GND.n3454 0.152939
R14139 GND.n3867 GND.n3454 0.152939
R14140 GND.n3868 GND.n3867 0.152939
R14141 GND.n3869 GND.n3868 0.152939
R14142 GND.n3870 GND.n3869 0.152939
R14143 GND.n3871 GND.n3870 0.152939
R14144 GND.n3872 GND.n3871 0.152939
R14145 GND.n3872 GND.n3402 0.152939
R14146 GND.n3992 GND.n3402 0.152939
R14147 GND.n6628 GND.n1087 0.152939
R14148 GND.n1092 GND.n1087 0.152939
R14149 GND.n1093 GND.n1092 0.152939
R14150 GND.n1094 GND.n1093 0.152939
R14151 GND.n1099 GND.n1094 0.152939
R14152 GND.n1100 GND.n1099 0.152939
R14153 GND.n1101 GND.n1100 0.152939
R14154 GND.n1102 GND.n1101 0.152939
R14155 GND.n1107 GND.n1102 0.152939
R14156 GND.n1108 GND.n1107 0.152939
R14157 GND.n1109 GND.n1108 0.152939
R14158 GND.n1110 GND.n1109 0.152939
R14159 GND.n1115 GND.n1110 0.152939
R14160 GND.n1116 GND.n1115 0.152939
R14161 GND.n1117 GND.n1116 0.152939
R14162 GND.n1118 GND.n1117 0.152939
R14163 GND.n1123 GND.n1118 0.152939
R14164 GND.n1124 GND.n1123 0.152939
R14165 GND.n1125 GND.n1124 0.152939
R14166 GND.n1126 GND.n1125 0.152939
R14167 GND.n1131 GND.n1126 0.152939
R14168 GND.n1132 GND.n1131 0.152939
R14169 GND.n1133 GND.n1132 0.152939
R14170 GND.n1134 GND.n1133 0.152939
R14171 GND.n1139 GND.n1134 0.152939
R14172 GND.n1140 GND.n1139 0.152939
R14173 GND.n1141 GND.n1140 0.152939
R14174 GND.n1142 GND.n1141 0.152939
R14175 GND.n1147 GND.n1142 0.152939
R14176 GND.n1148 GND.n1147 0.152939
R14177 GND.n1149 GND.n1148 0.152939
R14178 GND.n1150 GND.n1149 0.152939
R14179 GND.n1155 GND.n1150 0.152939
R14180 GND.n1156 GND.n1155 0.152939
R14181 GND.n1157 GND.n1156 0.152939
R14182 GND.n1158 GND.n1157 0.152939
R14183 GND.n1163 GND.n1158 0.152939
R14184 GND.n1164 GND.n1163 0.152939
R14185 GND.n1165 GND.n1164 0.152939
R14186 GND.n1166 GND.n1165 0.152939
R14187 GND.n1171 GND.n1166 0.152939
R14188 GND.n1172 GND.n1171 0.152939
R14189 GND.n1173 GND.n1172 0.152939
R14190 GND.n1174 GND.n1173 0.152939
R14191 GND.n1179 GND.n1174 0.152939
R14192 GND.n1180 GND.n1179 0.152939
R14193 GND.n1181 GND.n1180 0.152939
R14194 GND.n1182 GND.n1181 0.152939
R14195 GND.n1187 GND.n1182 0.152939
R14196 GND.n1188 GND.n1187 0.152939
R14197 GND.n1189 GND.n1188 0.152939
R14198 GND.n1190 GND.n1189 0.152939
R14199 GND.n1195 GND.n1190 0.152939
R14200 GND.n1196 GND.n1195 0.152939
R14201 GND.n1197 GND.n1196 0.152939
R14202 GND.n1198 GND.n1197 0.152939
R14203 GND.n1203 GND.n1198 0.152939
R14204 GND.n1204 GND.n1203 0.152939
R14205 GND.n1205 GND.n1204 0.152939
R14206 GND.n1206 GND.n1205 0.152939
R14207 GND.n1211 GND.n1206 0.152939
R14208 GND.n6500 GND.n1211 0.152939
R14209 GND.n6312 GND.n1429 0.152939
R14210 GND.n6308 GND.n1429 0.152939
R14211 GND.n6308 GND.n6307 0.152939
R14212 GND.n6307 GND.n6306 0.152939
R14213 GND.n6306 GND.n1434 0.152939
R14214 GND.n6302 GND.n1434 0.152939
R14215 GND.n6302 GND.n6301 0.152939
R14216 GND.n6301 GND.n6300 0.152939
R14217 GND.n6300 GND.n1439 0.152939
R14218 GND.n6296 GND.n1439 0.152939
R14219 GND.n6296 GND.n6295 0.152939
R14220 GND.n6295 GND.n6294 0.152939
R14221 GND.n6294 GND.n1444 0.152939
R14222 GND.n6290 GND.n1444 0.152939
R14223 GND.n6290 GND.n6289 0.152939
R14224 GND.n6289 GND.n6288 0.152939
R14225 GND.n6288 GND.n1449 0.152939
R14226 GND.n6284 GND.n1449 0.152939
R14227 GND.n6284 GND.n6283 0.152939
R14228 GND.n6283 GND.n6282 0.152939
R14229 GND.n6282 GND.n1454 0.152939
R14230 GND.n6278 GND.n1454 0.152939
R14231 GND.n6278 GND.n6277 0.152939
R14232 GND.n6270 GND.n6269 0.152939
R14233 GND.n6269 GND.n6268 0.152939
R14234 GND.n6268 GND.n1517 0.152939
R14235 GND.n6264 GND.n1517 0.152939
R14236 GND.n6264 GND.n6263 0.152939
R14237 GND.n6263 GND.n6262 0.152939
R14238 GND.n6262 GND.n1523 0.152939
R14239 GND.n6258 GND.n1523 0.152939
R14240 GND.n6258 GND.n6257 0.152939
R14241 GND.n6257 GND.n6256 0.152939
R14242 GND.n6256 GND.n1529 0.152939
R14243 GND.n6252 GND.n1529 0.152939
R14244 GND.n6252 GND.n6251 0.152939
R14245 GND.n6251 GND.n6250 0.152939
R14246 GND.n6250 GND.n1535 0.152939
R14247 GND.n1540 GND.n1535 0.152939
R14248 GND.n6245 GND.n1540 0.152939
R14249 GND.n6245 GND.n6244 0.152939
R14250 GND.n6244 GND.n6243 0.152939
R14251 GND.n6243 GND.n1544 0.152939
R14252 GND.n6239 GND.n1544 0.152939
R14253 GND.n6239 GND.n6238 0.152939
R14254 GND.n6238 GND.n6237 0.152939
R14255 GND.n6237 GND.n1550 0.152939
R14256 GND.n6233 GND.n1550 0.152939
R14257 GND.n6233 GND.n6232 0.152939
R14258 GND.n6232 GND.n6231 0.152939
R14259 GND.n6231 GND.n1556 0.152939
R14260 GND.n6227 GND.n1556 0.152939
R14261 GND.n6227 GND.n6226 0.152939
R14262 GND.n6226 GND.n6225 0.152939
R14263 GND.n6225 GND.n1562 0.152939
R14264 GND.n1566 GND.n1562 0.152939
R14265 GND.n3212 GND.n3211 0.152939
R14266 GND.n3217 GND.n3212 0.152939
R14267 GND.n3218 GND.n3217 0.152939
R14268 GND.n3219 GND.n3218 0.152939
R14269 GND.n3219 GND.n3207 0.152939
R14270 GND.n3225 GND.n3207 0.152939
R14271 GND.n3226 GND.n3225 0.152939
R14272 GND.n3227 GND.n3226 0.152939
R14273 GND.n3227 GND.n3203 0.152939
R14274 GND.n3233 GND.n3203 0.152939
R14275 GND.n3234 GND.n3233 0.152939
R14276 GND.n3235 GND.n3234 0.152939
R14277 GND.n3235 GND.n3199 0.152939
R14278 GND.n3241 GND.n3199 0.152939
R14279 GND.n3242 GND.n3241 0.152939
R14280 GND.n3243 GND.n3242 0.152939
R14281 GND.n3243 GND.n3192 0.152939
R14282 GND.n3249 GND.n3192 0.152939
R14283 GND.n3250 GND.n3249 0.152939
R14284 GND.n3251 GND.n3250 0.152939
R14285 GND.n3251 GND.n3188 0.152939
R14286 GND.n3257 GND.n3188 0.152939
R14287 GND.n3258 GND.n3257 0.152939
R14288 GND.n3259 GND.n3258 0.152939
R14289 GND.n3259 GND.n3184 0.152939
R14290 GND.n3265 GND.n3184 0.152939
R14291 GND.n3266 GND.n3265 0.152939
R14292 GND.n3267 GND.n3266 0.152939
R14293 GND.n3267 GND.n3180 0.152939
R14294 GND.n3273 GND.n3180 0.152939
R14295 GND.n3274 GND.n3273 0.152939
R14296 GND.n3275 GND.n3274 0.152939
R14297 GND.n3275 GND.n3176 0.152939
R14298 GND.n3281 GND.n3176 0.152939
R14299 GND.n3282 GND.n3281 0.152939
R14300 GND.n3283 GND.n3282 0.152939
R14301 GND.n3283 GND.n3168 0.152939
R14302 GND.n6377 GND.n1376 0.152939
R14303 GND.n6377 GND.n6376 0.152939
R14304 GND.n6376 GND.n6375 0.152939
R14305 GND.n6375 GND.n1378 0.152939
R14306 GND.n6371 GND.n1378 0.152939
R14307 GND.n6371 GND.n6370 0.152939
R14308 GND.n6370 GND.n6369 0.152939
R14309 GND.n6369 GND.n1384 0.152939
R14310 GND.n6365 GND.n1384 0.152939
R14311 GND.n6365 GND.n6364 0.152939
R14312 GND.n6364 GND.n6363 0.152939
R14313 GND.n6363 GND.n1390 0.152939
R14314 GND.n6359 GND.n1390 0.152939
R14315 GND.n6359 GND.n6358 0.152939
R14316 GND.n6358 GND.n6357 0.152939
R14317 GND.n6357 GND.n1396 0.152939
R14318 GND.n6350 GND.n1396 0.152939
R14319 GND.n6349 GND.n1399 0.152939
R14320 GND.n6345 GND.n1399 0.152939
R14321 GND.n6345 GND.n6344 0.152939
R14322 GND.n6344 GND.n6343 0.152939
R14323 GND.n6343 GND.n1404 0.152939
R14324 GND.n6339 GND.n1404 0.152939
R14325 GND.n6339 GND.n6338 0.152939
R14326 GND.n6338 GND.n6337 0.152939
R14327 GND.n6337 GND.n1409 0.152939
R14328 GND.n6333 GND.n1409 0.152939
R14329 GND.n6333 GND.n6332 0.152939
R14330 GND.n6332 GND.n6331 0.152939
R14331 GND.n6331 GND.n1414 0.152939
R14332 GND.n6327 GND.n1414 0.152939
R14333 GND.n6327 GND.n6326 0.152939
R14334 GND.n6326 GND.n6325 0.152939
R14335 GND.n6325 GND.n1419 0.152939
R14336 GND.n6321 GND.n1419 0.152939
R14337 GND.n6321 GND.n6320 0.152939
R14338 GND.n6320 GND.n6319 0.152939
R14339 GND.n6319 GND.n1424 0.152939
R14340 GND.n6315 GND.n1424 0.152939
R14341 GND.n6315 GND.n6314 0.152939
R14342 GND.n3993 GND.n3371 0.116354
R14343 GND.n2629 GND.n42 0.116354
R14344 GND.n4160 GND.n4159 0.108732
R14345 GND.n2399 GND.n2247 0.108732
R14346 GND.n8074 GND.n40 0.0767195
R14347 GND.n8074 GND.n41 0.0767195
R14348 GND.n4016 GND.n3382 0.0767195
R14349 GND.n3898 GND.n3382 0.0767195
R14350 GND.n8082 GND.n26 0.0695946
R14351 GND.n8082 GND.n8081 0.0695946
R14352 GND.n6313 GND.n6312 0.0695946
R14353 GND.n6314 GND.n6313 0.0695946
R14354 GND.n5443 GND.n2399 0.063
R14355 GND.n4159 GND.n4158 0.063
R14356 GND.n5443 GND.n5442 0.0534891
R14357 GND.n7879 GND.n7878 0.0534891
R14358 GND.n3775 GND.n3764 0.0534891
R14359 GND.n4158 GND.n4157 0.0534891
R14360 GND.n5043 GND.n2661 0.044054
R14361 GND.n6276 GND.n1459 0.044054
R14362 GND.n5038 GND.n2661 0.0423118
R14363 GND.n3123 GND.n1459 0.0423118
R14364 GND.n5148 GND.n42 0.0370854
R14365 GND.n3993 GND.n3992 0.0370854
R14366 GND.n5442 GND.n2401 0.0344674
R14367 GND.n5047 GND.n2401 0.0344674
R14368 GND.n5047 GND.n2452 0.0344674
R14369 GND.n2453 GND.n2452 0.0344674
R14370 GND.n2454 GND.n2453 0.0344674
R14371 GND.n5062 GND.n2454 0.0344674
R14372 GND.n5062 GND.n2472 0.0344674
R14373 GND.n2473 GND.n2472 0.0344674
R14374 GND.n2474 GND.n2473 0.0344674
R14375 GND.n5077 GND.n2474 0.0344674
R14376 GND.n5077 GND.n2493 0.0344674
R14377 GND.n2494 GND.n2493 0.0344674
R14378 GND.n2495 GND.n2494 0.0344674
R14379 GND.n5092 GND.n2495 0.0344674
R14380 GND.n5092 GND.n2514 0.0344674
R14381 GND.n2515 GND.n2514 0.0344674
R14382 GND.n2516 GND.n2515 0.0344674
R14383 GND.n5107 GND.n2516 0.0344674
R14384 GND.n5107 GND.n2533 0.0344674
R14385 GND.n2534 GND.n2533 0.0344674
R14386 GND.n2535 GND.n2534 0.0344674
R14387 GND.n5127 GND.n2535 0.0344674
R14388 GND.n5128 GND.n5127 0.0344674
R14389 GND.n5132 GND.n5128 0.0344674
R14390 GND.n5132 GND.n2558 0.0344674
R14391 GND.n5358 GND.n2558 0.0344674
R14392 GND.n5358 GND.n2559 0.0344674
R14393 GND.n2559 GND.n57 0.0344674
R14394 GND.n58 GND.n57 0.0344674
R14395 GND.n59 GND.n58 0.0344674
R14396 GND.n5203 GND.n59 0.0344674
R14397 GND.n5203 GND.n77 0.0344674
R14398 GND.n78 GND.n77 0.0344674
R14399 GND.n79 GND.n78 0.0344674
R14400 GND.n5210 GND.n79 0.0344674
R14401 GND.n5210 GND.n98 0.0344674
R14402 GND.n99 GND.n98 0.0344674
R14403 GND.n100 GND.n99 0.0344674
R14404 GND.n5217 GND.n100 0.0344674
R14405 GND.n5217 GND.n119 0.0344674
R14406 GND.n120 GND.n119 0.0344674
R14407 GND.n121 GND.n120 0.0344674
R14408 GND.n5224 GND.n121 0.0344674
R14409 GND.n5224 GND.n140 0.0344674
R14410 GND.n141 GND.n140 0.0344674
R14411 GND.n142 GND.n141 0.0344674
R14412 GND.n7878 GND.n142 0.0344674
R14413 GND.n3775 GND.n3774 0.0344674
R14414 GND.n3774 GND.n3773 0.0344674
R14415 GND.n3773 GND.n3771 0.0344674
R14416 GND.n3771 GND.n3504 0.0344674
R14417 GND.n3813 GND.n3504 0.0344674
R14418 GND.n3813 GND.n3505 0.0344674
R14419 GND.n3809 GND.n3505 0.0344674
R14420 GND.n3809 GND.n3808 0.0344674
R14421 GND.n3808 GND.n3475 0.0344674
R14422 GND.n3850 GND.n3475 0.0344674
R14423 GND.n3850 GND.n3476 0.0344674
R14424 GND.n3846 GND.n3476 0.0344674
R14425 GND.n3846 GND.n3845 0.0344674
R14426 GND.n3845 GND.n3446 0.0344674
R14427 GND.n3890 GND.n3446 0.0344674
R14428 GND.n3890 GND.n3447 0.0344674
R14429 GND.n3886 GND.n3447 0.0344674
R14430 GND.n3886 GND.n3427 0.0344674
R14431 GND.n3907 GND.n3427 0.0344674
R14432 GND.n3907 GND.n3424 0.0344674
R14433 GND.n3978 GND.n3424 0.0344674
R14434 GND.n3978 GND.n3425 0.0344674
R14435 GND.n3974 GND.n3425 0.0344674
R14436 GND.n3974 GND.n3973 0.0344674
R14437 GND.n3973 GND.n3972 0.0344674
R14438 GND.n3972 GND.n3918 0.0344674
R14439 GND.n3926 GND.n3918 0.0344674
R14440 GND.n3926 GND.n3391 0.0344674
R14441 GND.n4010 GND.n3391 0.0344674
R14442 GND.n4010 GND.n3392 0.0344674
R14443 GND.n4006 GND.n3392 0.0344674
R14444 GND.n4006 GND.n4005 0.0344674
R14445 GND.n4005 GND.n3363 0.0344674
R14446 GND.n4047 GND.n3363 0.0344674
R14447 GND.n4047 GND.n3364 0.0344674
R14448 GND.n4043 GND.n3364 0.0344674
R14449 GND.n4043 GND.n4042 0.0344674
R14450 GND.n4042 GND.n3334 0.0344674
R14451 GND.n4084 GND.n3334 0.0344674
R14452 GND.n4084 GND.n3335 0.0344674
R14453 GND.n4080 GND.n3335 0.0344674
R14454 GND.n4080 GND.n4079 0.0344674
R14455 GND.n4079 GND.n3305 0.0344674
R14456 GND.n4139 GND.n3305 0.0344674
R14457 GND.n4139 GND.n3306 0.0344674
R14458 GND.n3306 GND.n3169 0.0344674
R14459 GND.n4157 GND.n3169 0.0344674
R14460 GND.n2249 GND.n2248 0.0343753
R14461 GND.n5036 GND.n5035 0.0343753
R14462 GND.n3167 GND.n3166 0.0343753
R14463 GND.n3127 GND.n3115 0.0343753
R14464 GND.n2407 GND.n2250 0.0272615
R14465 GND.n2408 GND.n2251 0.0272615
R14466 GND.n2409 GND.n2252 0.0272615
R14467 GND.n2410 GND.n2253 0.0272615
R14468 GND.n2411 GND.n2254 0.0272615
R14469 GND.n2412 GND.n2255 0.0272615
R14470 GND.n2413 GND.n2256 0.0272615
R14471 GND.n2414 GND.n2257 0.0272615
R14472 GND.n2415 GND.n2258 0.0272615
R14473 GND.n5593 GND.n2262 0.0272615
R14474 GND.n5592 GND.n2263 0.0272615
R14475 GND.n5028 GND.n2669 0.0272615
R14476 GND.n5029 GND.n2668 0.0272615
R14477 GND.n3163 GND.n3072 0.0272615
R14478 GND.n3162 GND.n3078 0.0272615
R14479 GND.n3159 GND.n3158 0.0272615
R14480 GND.n3155 GND.n3084 0.0272615
R14481 GND.n3154 GND.n3088 0.0272615
R14482 GND.n3151 GND.n3150 0.0272615
R14483 GND.n3147 GND.n3092 0.0272615
R14484 GND.n3146 GND.n3098 0.0272615
R14485 GND.n3143 GND.n3142 0.0272615
R14486 GND.n3136 GND.n3104 0.0272615
R14487 GND.n3135 GND.n3107 0.0272615
R14488 GND.n3132 GND.n3131 0.0272615
R14489 GND.n3128 GND.n3111 0.0272615
R14490 GND.n5037 GND.n5036 0.026584
R14491 GND.n3122 GND.n3115 0.026584
R14492 GND.n2399 GND.n2248 0.0103238
R14493 GND.n4159 GND.n3167 0.0103238
R14494 GND.n5038 GND.n5037 0.00829133
R14495 GND.n3123 GND.n3122 0.00829133
R14496 GND.n2407 GND.n2249 0.00761382
R14497 GND.n2408 GND.n2250 0.00761382
R14498 GND.n2409 GND.n2251 0.00761382
R14499 GND.n2410 GND.n2252 0.00761382
R14500 GND.n2411 GND.n2253 0.00761382
R14501 GND.n2412 GND.n2254 0.00761382
R14502 GND.n2413 GND.n2255 0.00761382
R14503 GND.n2414 GND.n2256 0.00761382
R14504 GND.n2415 GND.n2257 0.00761382
R14505 GND.n2262 GND.n2258 0.00761382
R14506 GND.n5593 GND.n5592 0.00761382
R14507 GND.n2669 GND.n2263 0.00761382
R14508 GND.n5029 GND.n5028 0.00761382
R14509 GND.n5035 GND.n2668 0.00761382
R14510 GND.n3166 GND.n3072 0.00761382
R14511 GND.n3163 GND.n3162 0.00761382
R14512 GND.n3159 GND.n3078 0.00761382
R14513 GND.n3158 GND.n3084 0.00761382
R14514 GND.n3155 GND.n3154 0.00761382
R14515 GND.n3151 GND.n3088 0.00761382
R14516 GND.n3150 GND.n3092 0.00761382
R14517 GND.n3147 GND.n3146 0.00761382
R14518 GND.n3143 GND.n3098 0.00761382
R14519 GND.n3142 GND.n3104 0.00761382
R14520 GND.n3136 GND.n3135 0.00761382
R14521 GND.n3132 GND.n3107 0.00761382
R14522 GND.n3131 GND.n3111 0.00761382
R14523 GND.n3128 GND.n3127 0.00761382
R14524 CS_BIAS.n8 CS_BIAS.n2 161.3
R14525 CS_BIAS.n10 CS_BIAS.n9 161.3
R14526 CS_BIAS.n11 CS_BIAS.n1 161.3
R14527 CS_BIAS.n13 CS_BIAS.n12 161.3
R14528 CS_BIAS.n14 CS_BIAS.n0 161.3
R14529 CS_BIAS.n37 CS_BIAS.n23 161.3
R14530 CS_BIAS.n36 CS_BIAS.n35 161.3
R14531 CS_BIAS.n34 CS_BIAS.n24 161.3
R14532 CS_BIAS.n33 CS_BIAS.n32 161.3
R14533 CS_BIAS.n31 CS_BIAS.n25 161.3
R14534 CS_BIAS.n8 CS_BIAS.n7 118.987
R14535 CS_BIAS.n31 CS_BIAS.n30 118.987
R14536 CS_BIAS.n16 CS_BIAS.n15 69.2143
R14537 CS_BIAS.n39 CS_BIAS.n38 69.2143
R14538 CS_BIAS.n21 CS_BIAS.t20 67.3598
R14539 CS_BIAS.n44 CS_BIAS.t14 67.3598
R14540 CS_BIAS.n42 CS_BIAS.t23 67.3598
R14541 CS_BIAS.n40 CS_BIAS.t15 67.3598
R14542 CS_BIAS.n27 CS_BIAS.t4 67.3598
R14543 CS_BIAS.n19 CS_BIAS.t13 67.3595
R14544 CS_BIAS.n17 CS_BIAS.t21 67.3595
R14545 CS_BIAS.n3 CS_BIAS.t2 67.3595
R14546 CS_BIAS.n19 CS_BIAS.t19 65.6135
R14547 CS_BIAS.n17 CS_BIAS.t12 65.6135
R14548 CS_BIAS.n3 CS_BIAS.t0 65.6135
R14549 CS_BIAS.n21 CS_BIAS.t11 65.6135
R14550 CS_BIAS.n44 CS_BIAS.t8 65.6135
R14551 CS_BIAS.n42 CS_BIAS.t16 65.6135
R14552 CS_BIAS.n40 CS_BIAS.t10 65.6135
R14553 CS_BIAS.n27 CS_BIAS.t6 65.6135
R14554 CS_BIAS.n5 CS_BIAS.n4 62.1308
R14555 CS_BIAS.n28 CS_BIAS.n26 62.1308
R14556 CS_BIAS.n30 CS_BIAS.t18 57.8552
R14557 CS_BIAS.n7 CS_BIAS.t22 57.8549
R14558 CS_BIAS.n15 CS_BIAS.t9 32.5934
R14559 CS_BIAS.n38 CS_BIAS.t17 32.5934
R14560 CS_BIAS.n9 CS_BIAS.n8 32.2376
R14561 CS_BIAS.n32 CS_BIAS.n31 32.2376
R14562 CS_BIAS.n14 CS_BIAS.n13 24.4675
R14563 CS_BIAS.n13 CS_BIAS.n1 24.4675
R14564 CS_BIAS.n9 CS_BIAS.n1 24.4675
R14565 CS_BIAS.n32 CS_BIAS.n24 24.4675
R14566 CS_BIAS.n36 CS_BIAS.n24 24.4675
R14567 CS_BIAS.n37 CS_BIAS.n36 24.4675
R14568 CS_BIAS.n28 CS_BIAS.n27 14.3395
R14569 CS_BIAS.n5 CS_BIAS.n3 14.3395
R14570 CS_BIAS.n15 CS_BIAS.n14 12.968
R14571 CS_BIAS.n38 CS_BIAS.n37 12.968
R14572 CS_BIAS.n46 CS_BIAS.n22 10.7248
R14573 CS_BIAS.n30 CS_BIAS.n29 9.62147
R14574 CS_BIAS.n7 CS_BIAS.n6 9.62138
R14575 CS_BIAS.n6 CS_BIAS.n5 9.503
R14576 CS_BIAS.n29 CS_BIAS.n28 9.503
R14577 CS_BIAS.n18 CS_BIAS.n16 8.80338
R14578 CS_BIAS.n41 CS_BIAS.n39 8.80338
R14579 CS_BIAS.n46 CS_BIAS.n45 7.64156
R14580 CS_BIAS.n4 CS_BIAS.t1 6.70101
R14581 CS_BIAS.n4 CS_BIAS.t3 6.70101
R14582 CS_BIAS.n26 CS_BIAS.t5 6.70101
R14583 CS_BIAS.n26 CS_BIAS.t7 6.70101
R14584 CS_BIAS.n22 CS_BIAS.n21 6.15589
R14585 CS_BIAS.n45 CS_BIAS.n44 6.15589
R14586 CS_BIAS.n43 CS_BIAS.n42 6.15589
R14587 CS_BIAS.n41 CS_BIAS.n40 6.15589
R14588 CS_BIAS.n20 CS_BIAS.n19 6.15588
R14589 CS_BIAS.n18 CS_BIAS.n17 6.15588
R14590 CS_BIAS CS_BIAS.n46 4.87447
R14591 CS_BIAS.n20 CS_BIAS.n18 3.5005
R14592 CS_BIAS.n22 CS_BIAS.n20 3.5005
R14593 CS_BIAS.n43 CS_BIAS.n41 3.5005
R14594 CS_BIAS.n45 CS_BIAS.n43 3.5005
R14595 CS_BIAS.n16 CS_BIAS.n0 0.417535
R14596 CS_BIAS.n39 CS_BIAS.n23 0.417535
R14597 CS_BIAS.n12 CS_BIAS.n0 0.189894
R14598 CS_BIAS.n12 CS_BIAS.n11 0.189894
R14599 CS_BIAS.n11 CS_BIAS.n10 0.189894
R14600 CS_BIAS.n10 CS_BIAS.n2 0.189894
R14601 CS_BIAS.n33 CS_BIAS.n25 0.189894
R14602 CS_BIAS.n34 CS_BIAS.n33 0.189894
R14603 CS_BIAS.n35 CS_BIAS.n34 0.189894
R14604 CS_BIAS.n35 CS_BIAS.n23 0.189894
R14605 CS_BIAS.n6 CS_BIAS.n2 0.0762576
R14606 CS_BIAS.n29 CS_BIAS.n25 0.0762576
R14607 VOUT.n7 VOUT.t24 181.174
R14608 VOUT.n9 VOUT.t17 180.333
R14609 VOUT.n8 VOUT.t25 180.333
R14610 VOUT.n7 VOUT.t19 180.333
R14611 VOUT.n10 VOUT.t18 180.333
R14612 VOUT.n0 VOUT.t21 180.23
R14613 VOUT.n3 VOUT.t23 179.387
R14614 VOUT.n2 VOUT.t22 179.387
R14615 VOUT.n1 VOUT.t20 179.387
R14616 VOUT.n0 VOUT.t16 179.387
R14617 VOUT.n14 VOUT.n12 69.0058
R14618 VOUT.n22 VOUT.n20 69.0058
R14619 VOUT.n18 VOUT.n17 67.6638
R14620 VOUT.n16 VOUT.n15 67.6638
R14621 VOUT.n14 VOUT.n13 67.6638
R14622 VOUT.n26 VOUT.n25 67.6638
R14623 VOUT.n24 VOUT.n23 67.6638
R14624 VOUT.n22 VOUT.n21 67.6638
R14625 VOUT.n19 VOUT.n11 9.52907
R14626 VOUT.n17 VOUT.t12 6.70101
R14627 VOUT.n17 VOUT.t3 6.70101
R14628 VOUT.n15 VOUT.t4 6.70101
R14629 VOUT.n15 VOUT.t10 6.70101
R14630 VOUT.n13 VOUT.t11 6.70101
R14631 VOUT.n13 VOUT.t2 6.70101
R14632 VOUT.n12 VOUT.t14 6.70101
R14633 VOUT.n12 VOUT.t1 6.70101
R14634 VOUT.n25 VOUT.t9 6.70101
R14635 VOUT.n25 VOUT.t15 6.70101
R14636 VOUT.n23 VOUT.t0 6.70101
R14637 VOUT.n23 VOUT.t7 6.70101
R14638 VOUT.n21 VOUT.t8 6.70101
R14639 VOUT.n21 VOUT.t13 6.70101
R14640 VOUT.n20 VOUT.t5 6.70101
R14641 VOUT.n20 VOUT.t6 6.70101
R14642 VOUT.n11 VOUT.n4 5.57564
R14643 VOUT.n28 VOUT.n4 4.87459
R14644 VOUT.n28 VOUT.n27 4.63548
R14645 VOUT.n11 VOUT.n10 4.39182
R14646 VOUT.n4 VOUT.n3 4.39182
R14647 VOUT.n19 VOUT.n18 4.24958
R14648 VOUT.n27 VOUT.n26 4.24958
R14649 VOUT.n27 VOUT.n19 3.82348
R14650 VOUT.n6 VOUT 3.2247
R14651 VOUT.n18 VOUT.n16 1.34245
R14652 VOUT.n16 VOUT.n14 1.34245
R14653 VOUT.n26 VOUT.n24 1.34245
R14654 VOUT.n24 VOUT.n22 1.34245
R14655 VOUT.n10 VOUT.n9 0.842454
R14656 VOUT.n9 VOUT.n8 0.842454
R14657 VOUT.n8 VOUT.n7 0.842454
R14658 VOUT.n3 VOUT.n2 0.842454
R14659 VOUT.n2 VOUT.n1 0.842454
R14660 VOUT.n1 VOUT.n0 0.842454
R14661 VOUT.n6 VOUT.n5 0.372359
R14662 VOUT.n28 VOUT.n6 0.31352
R14663 VOUT.n5 VOUT.t27 0.100127
R14664 VOUT.n5 VOUT.t26 0.0245871
R14665 VOUT VOUT.n28 0.0099
R14666 VN.n2 VN.t0 243.97
R14667 VN.n2 VN.n1 223.454
R14668 VN.n4 VN.n3 223.454
R14669 VN.n6 VN.n5 223.454
R14670 VN.n0 VN.t8 153.089
R14671 VN.n0 VN.t7 136.929
R14672 VN.n1 VN.t1 19.8005
R14673 VN.n1 VN.t4 19.8005
R14674 VN.n3 VN.t2 19.8005
R14675 VN.n3 VN.t6 19.8005
R14676 VN.n5 VN.t3 19.8005
R14677 VN.n5 VN.t5 19.8005
R14678 VN VN.n7 17.5959
R14679 VN.n7 VN.n6 5.40567
R14680 VN.n7 VN.n0 1.188
R14681 VN.n6 VN.n4 0.716017
R14682 VN.n4 VN.n2 0.716017
R14683 a_n11634_10845.n78 a_n11634_10845.n77 28.5533
R14684 a_n11634_10845.n80 a_n11634_10845.n79 21.6125
R14685 a_n11634_10845.n82 a_n11634_10845.n81 28.5533
R14686 a_n11634_10845.n83 a_n11634_10845.n131 161.3
R14687 a_n11634_10845.n84 a_n11634_10845.n83 44.4798
R14688 a_n11634_10845.n86 a_n11634_10845.n85 23.1536
R14689 a_n11634_10845.n88 a_n11634_10845.n87 28.5533
R14690 a_n11634_10845.n89 a_n11634_10845.n104 74.9922
R14691 a_n11634_10845.n132 a_n11634_10845.n104 11.3187
R14692 a_n11634_10845.n103 a_n11634_10845.n89 74.9922
R14693 a_n11634_10845.n91 a_n11634_10845.n90 27.591
R14694 a_n11634_10845.n93 a_n11634_10845.n92 27.7992
R14695 a_n11634_10845.n94 a_n11634_10845.n102 74.9922
R14696 a_n11634_10845.n101 a_n11634_10845.n94 74.9922
R14697 a_n11634_10845.n96 a_n11634_10845.n95 28.5533
R14698 a_n11634_10845.n98 a_n11634_10845.n97 23.3672
R14699 a_n11634_10845.n100 a_n11634_10845.n99 44.4798
R14700 a_n11634_10845.n53 a_n11634_10845.n52 28.5533
R14701 a_n11634_10845.n55 a_n11634_10845.n54 21.6125
R14702 a_n11634_10845.n57 a_n11634_10845.n56 28.5533
R14703 a_n11634_10845.n58 a_n11634_10845.n125 161.3
R14704 a_n11634_10845.n59 a_n11634_10845.n58 44.4798
R14705 a_n11634_10845.n61 a_n11634_10845.n60 23.1536
R14706 a_n11634_10845.n63 a_n11634_10845.n62 28.5533
R14707 a_n11634_10845.n64 a_n11634_10845.n108 74.9922
R14708 a_n11634_10845.n126 a_n11634_10845.n108 11.3187
R14709 a_n11634_10845.n107 a_n11634_10845.n64 74.9922
R14710 a_n11634_10845.n66 a_n11634_10845.n65 27.591
R14711 a_n11634_10845.n68 a_n11634_10845.n67 27.7992
R14712 a_n11634_10845.n69 a_n11634_10845.n106 74.9922
R14713 a_n11634_10845.n105 a_n11634_10845.n69 74.9922
R14714 a_n11634_10845.n71 a_n11634_10845.n70 28.5533
R14715 a_n11634_10845.n73 a_n11634_10845.n72 23.3672
R14716 a_n11634_10845.n75 a_n11634_10845.n74 44.4798
R14717 a_n11634_10845.n28 a_n11634_10845.n27 28.5533
R14718 a_n11634_10845.n30 a_n11634_10845.n29 21.6125
R14719 a_n11634_10845.n32 a_n11634_10845.n31 28.5533
R14720 a_n11634_10845.n33 a_n11634_10845.n149 161.3
R14721 a_n11634_10845.n34 a_n11634_10845.n33 44.4798
R14722 a_n11634_10845.n36 a_n11634_10845.n35 23.1536
R14723 a_n11634_10845.n38 a_n11634_10845.n37 28.5533
R14724 a_n11634_10845.n39 a_n11634_10845.n112 74.9922
R14725 a_n11634_10845.n150 a_n11634_10845.n112 11.3187
R14726 a_n11634_10845.n111 a_n11634_10845.n39 74.9922
R14727 a_n11634_10845.n41 a_n11634_10845.n40 27.591
R14728 a_n11634_10845.n43 a_n11634_10845.n42 27.7992
R14729 a_n11634_10845.n44 a_n11634_10845.n110 74.9922
R14730 a_n11634_10845.n109 a_n11634_10845.n44 74.9922
R14731 a_n11634_10845.n46 a_n11634_10845.n45 28.5533
R14732 a_n11634_10845.n48 a_n11634_10845.n47 23.3672
R14733 a_n11634_10845.n50 a_n11634_10845.n49 44.4798
R14734 a_n11634_10845.n14 a_n11634_10845.n21 44.4798
R14735 a_n11634_10845.n18 a_n11634_10845.n23 27.4881
R14736 a_n11634_10845.n22 a_n11634_10845.n25 27.9045
R14737 a_n11634_10845.n114 a_n11634_10845.n24 74.9922
R14738 a_n11634_10845.n138 a_n11634_10845.t2 156.754
R14739 a_n11634_10845.n119 a_n11634_10845.t4 154.892
R14740 a_n11634_10845.n118 a_n11634_10845.n116 131.358
R14741 a_n11634_10845.n118 a_n11634_10845.n117 129.496
R14742 a_n11634_10845.n138 a_n11634_10845.n137 129.496
R14743 a_n11634_10845.n140 a_n11634_10845.n139 129.496
R14744 a_n11634_10845.t0 a_n11634_10845.n155 97.5754
R14745 a_n11634_10845.n16 a_n11634_10845.n136 75.8453
R14746 a_n11634_10845.n8 a_n11634_10845.n146 77.0535
R14747 a_n11634_10845.n5 a_n11634_10845.n145 77.0535
R14748 a_n11634_10845.n2 a_n11634_10845.n144 77.0535
R14749 a_n11634_10845.n19 a_n11634_10845.n20 51.1079
R14750 a_n11634_10845.n63 a_n11634_10845.n61 114.397
R14751 a_n11634_10845.n88 a_n11634_10845.n86 114.397
R14752 a_n11634_10845.n38 a_n11634_10845.n36 114.397
R14753 a_n11634_10845.n155 a_n11634_10845.t21 67.4583
R14754 a_n11634_10845.n10 a_n11634_10845.n9 0.235669
R14755 a_n11634_10845.n129 a_n11634_10845.n128 54.6972
R14756 a_n11634_10845.n124 a_n11634_10845.n51 54.6972
R14757 a_n11634_10845.n135 a_n11634_10845.n134 54.6972
R14758 a_n11634_10845.n130 a_n11634_10845.n76 54.6972
R14759 a_n11634_10845.n153 a_n11634_10845.n152 54.6972
R14760 a_n11634_10845.n148 a_n11634_10845.n26 54.6972
R14761 a_n11634_10845.n113 a_n11634_10845.n121 54.2104
R14762 a_n11634_10845.n14 a_n11634_10845.n15 0.343823
R14763 a_n11634_10845.n57 a_n11634_10845.n55 99.2359
R14764 a_n11634_10845.n82 a_n11634_10845.n80 99.2359
R14765 a_n11634_10845.n32 a_n11634_10845.n30 99.2359
R14766 a_n11634_10845.n25 a_n11634_10845.n23 139.371
R14767 a_n11634_10845.n68 a_n11634_10845.n66 139.382
R14768 a_n11634_10845.n93 a_n11634_10845.n91 139.382
R14769 a_n11634_10845.n43 a_n11634_10845.n41 139.382
R14770 a_n11634_10845.n117 a_n11634_10845.t6 25.395
R14771 a_n11634_10845.n117 a_n11634_10845.t18 25.395
R14772 a_n11634_10845.n116 a_n11634_10845.t20 25.395
R14773 a_n11634_10845.n116 a_n11634_10845.t8 25.395
R14774 a_n11634_10845.n137 a_n11634_10845.t16 25.395
R14775 a_n11634_10845.n137 a_n11634_10845.t10 25.395
R14776 a_n11634_10845.n139 a_n11634_10845.t12 25.395
R14777 a_n11634_10845.n139 a_n11634_10845.t14 25.395
R14778 a_n11634_10845.n155 a_n11634_10845.n154 24.3555
R14779 a_n11634_10845.n6 a_n11634_10845.n8 1.27042
R14780 a_n11634_10845.n3 a_n11634_10845.n5 1.27042
R14781 a_n11634_10845.n0 a_n11634_10845.n2 1.27042
R14782 a_n11634_10845.n114 a_n11634_10845.n25 65.6956
R14783 a_n11634_10845.n23 a_n11634_10845.n21 76.061
R14784 a_n11634_10845.n20 a_n11634_10845.n15 76.1683
R14785 a_n11634_10845.n75 a_n11634_10845.n73 81.7953
R14786 a_n11634_10845.n73 a_n11634_10845.n71 115.942
R14787 a_n11634_10845.n71 a_n11634_10845.n105 64.8679
R14788 a_n11634_10845.n105 a_n11634_10845.n127 12.2924
R14789 a_n11634_10845.n106 a_n11634_10845.n68 65.8299
R14790 a_n11634_10845.n66 a_n11634_10845.n107 66.0955
R14791 a_n11634_10845.n107 a_n11634_10845.n126 35.6621
R14792 a_n11634_10845.n108 a_n11634_10845.n63 64.8679
R14793 a_n11634_10845.n61 a_n11634_10845.n59 82.2525
R14794 a_n11634_10845.n125 a_n11634_10845.n57 53.5497
R14795 a_n11634_10845.n55 a_n11634_10845.n53 97.3159
R14796 a_n11634_10845.n124 a_n11634_10845.n53 51.6022
R14797 a_n11634_10845.n100 a_n11634_10845.n98 81.7953
R14798 a_n11634_10845.n98 a_n11634_10845.n96 115.942
R14799 a_n11634_10845.n96 a_n11634_10845.n101 64.8679
R14800 a_n11634_10845.n101 a_n11634_10845.n133 12.2924
R14801 a_n11634_10845.n102 a_n11634_10845.n93 65.8299
R14802 a_n11634_10845.n91 a_n11634_10845.n103 66.0955
R14803 a_n11634_10845.n103 a_n11634_10845.n132 35.6621
R14804 a_n11634_10845.n104 a_n11634_10845.n88 64.8679
R14805 a_n11634_10845.n86 a_n11634_10845.n84 82.2525
R14806 a_n11634_10845.n131 a_n11634_10845.n82 53.5497
R14807 a_n11634_10845.n80 a_n11634_10845.n78 97.3159
R14808 a_n11634_10845.n130 a_n11634_10845.n78 51.6022
R14809 a_n11634_10845.n50 a_n11634_10845.n48 81.7953
R14810 a_n11634_10845.n48 a_n11634_10845.n46 115.942
R14811 a_n11634_10845.n46 a_n11634_10845.n109 64.8679
R14812 a_n11634_10845.n109 a_n11634_10845.n151 12.2924
R14813 a_n11634_10845.n110 a_n11634_10845.n43 65.8299
R14814 a_n11634_10845.n41 a_n11634_10845.n111 66.0955
R14815 a_n11634_10845.n111 a_n11634_10845.n150 35.6621
R14816 a_n11634_10845.n112 a_n11634_10845.n38 64.8679
R14817 a_n11634_10845.n36 a_n11634_10845.n34 82.2525
R14818 a_n11634_10845.n149 a_n11634_10845.n32 53.5497
R14819 a_n11634_10845.n30 a_n11634_10845.n28 97.3159
R14820 a_n11634_10845.n148 a_n11634_10845.n28 51.6022
R14821 a_n11634_10845.n19 a_n11634_10845.n143 75.4477
R14822 a_n11634_10845.n17 a_n11634_10845.n9 1.9706
R14823 a_n11634_10845.n127 a_n11634_10845.n106 34.6884
R14824 a_n11634_10845.n59 a_n11634_10845.n123 44.5222
R14825 a_n11634_10845.n133 a_n11634_10845.n102 34.6884
R14826 a_n11634_10845.n84 a_n11634_10845.n122 44.5222
R14827 a_n11634_10845.n151 a_n11634_10845.n110 34.6884
R14828 a_n11634_10845.n34 a_n11634_10845.n115 44.5222
R14829 a_n11634_10845.n6 a_n11634_10845.n7 3.10822
R14830 a_n11634_10845.n3 a_n11634_10845.n4 3.10822
R14831 a_n11634_10845.n0 a_n11634_10845.n1 3.10822
R14832 a_n11634_10845.n114 a_n11634_10845.n121 34.2015
R14833 a_n11634_10845.n128 a_n11634_10845.n75 43.5485
R14834 a_n11634_10845.n134 a_n11634_10845.n100 43.5485
R14835 a_n11634_10845.n152 a_n11634_10845.n50 43.5485
R14836 a_n11634_10845.n142 a_n11634_10845.n135 17.8223
R14837 a_n11634_10845.n26 a_n11634_10845.n147 17.4019
R14838 a_n11634_10845.n141 a_n11634_10845.n9 15.7693
R14839 a_n11634_10845.n51 a_n11634_10845.n120 14.3697
R14840 a_n11634_10845.n16 a_n11634_10845.t15 40.8349
R14841 a_n11634_10845.n17 a_n11634_10845.t11 42.9398
R14842 a_n11634_10845.n17 a_n11634_10845.t13 40.9556
R14843 a_n11634_10845.n136 a_n11634_10845.t9 10.6012
R14844 a_n11634_10845.n10 a_n11634_10845.t1 41.9092
R14845 a_n11634_10845.n7 a_n11634_10845.t37 41.3588
R14846 a_n11634_10845.n8 a_n11634_10845.t27 40.298
R14847 a_n11634_10845.n146 a_n11634_10845.t43 10.6012
R14848 a_n11634_10845.n11 a_n11634_10845.t42 41.8371
R14849 a_n11634_10845.n4 a_n11634_10845.t25 41.3588
R14850 a_n11634_10845.n5 a_n11634_10845.t45 40.298
R14851 a_n11634_10845.n145 a_n11634_10845.t24 10.6012
R14852 a_n11634_10845.n12 a_n11634_10845.t22 41.8371
R14853 a_n11634_10845.n1 a_n11634_10845.t47 41.3588
R14854 a_n11634_10845.n2 a_n11634_10845.t23 40.298
R14855 a_n11634_10845.n144 a_n11634_10845.t44 10.6012
R14856 a_n11634_10845.n13 a_n11634_10845.t26 41.8371
R14857 a_n11634_10845.n121 a_n11634_10845.t39 10.6012
R14858 a_n11634_10845.n143 a_n11634_10845.t33 10.6012
R14859 a_n11634_10845.n15 a_n11634_10845.t36 41.7273
R14860 a_n11634_10845.n126 a_n11634_10845.t5 10.6012
R14861 a_n11634_10845.n128 a_n11634_10845.t19 10.6012
R14862 a_n11634_10845.n127 a_n11634_10845.t7 10.6012
R14863 a_n11634_10845.n123 a_n11634_10845.t17 10.6012
R14864 a_n11634_10845.n124 a_n11634_10845.t3 10.6012
R14865 a_n11634_10845.n132 a_n11634_10845.t30 10.6012
R14866 a_n11634_10845.n134 a_n11634_10845.t28 10.6012
R14867 a_n11634_10845.n133 a_n11634_10845.t32 10.6012
R14868 a_n11634_10845.n122 a_n11634_10845.t35 10.6012
R14869 a_n11634_10845.n130 a_n11634_10845.t29 10.6012
R14870 a_n11634_10845.n150 a_n11634_10845.t46 10.6012
R14871 a_n11634_10845.n152 a_n11634_10845.t38 10.6012
R14872 a_n11634_10845.n151 a_n11634_10845.t41 10.6012
R14873 a_n11634_10845.n115 a_n11634_10845.t34 10.6012
R14874 a_n11634_10845.n148 a_n11634_10845.t31 10.6012
R14875 a_n11634_10845.n76 a_n11634_10845.n129 10.0381
R14876 a_n11634_10845.n120 a_n11634_10845.n119 9.32064
R14877 a_n11634_10845.n141 a_n11634_10845.n140 8.8403
R14878 a_n11634_10845.n113 a_n11634_10845.n142 8.60452
R14879 a_n11634_10845.n147 a_n11634_10845.n6 8.60452
R14880 a_n11634_10845.n154 a_n11634_10845.n153 5.83179
R14881 a_n11634_10845.n4 a_n11634_10845.n0 5.37591
R14882 a_n11634_10845.n154 a_n11634_10845.n9 4.16891
R14883 a_n11634_10845.n147 a_n11634_10845.n120 3.45315
R14884 a_n11634_10845.n1 a_n11634_10845.n14 3.87591
R14885 a_n11634_10845.n7 a_n11634_10845.n3 3.87591
R14886 a_n11634_10845.n119 a_n11634_10845.n118 1.86257
R14887 a_n11634_10845.n140 a_n11634_10845.n138 1.86257
R14888 a_n11634_10845.n142 a_n11634_10845.n141 1.63308
R14889 a_n11634_10845.n10 a_n11634_10845.n136 52.641
R14890 a_n11634_10845.n125 a_n11634_10845.n123 0.974237
R14891 a_n11634_10845.n131 a_n11634_10845.n122 0.974237
R14892 a_n11634_10845.n149 a_n11634_10845.n115 0.974237
R14893 a_n11634_10845.n77 a_n11634_10845.n76 0.881933
R14894 a_n11634_10845.n52 a_n11634_10845.n51 0.881933
R14895 a_n11634_10845.n27 a_n11634_10845.n26 0.881933
R14896 a_n11634_10845.n99 a_n11634_10845.n97 0.758076
R14897 a_n11634_10845.n97 a_n11634_10845.n95 0.758076
R14898 a_n11634_10845.n95 a_n11634_10845.n94 0.758076
R14899 a_n11634_10845.n94 a_n11634_10845.n92 0.758076
R14900 a_n11634_10845.n92 a_n11634_10845.n90 0.758076
R14901 a_n11634_10845.n90 a_n11634_10845.n89 0.758076
R14902 a_n11634_10845.n89 a_n11634_10845.n87 0.758076
R14903 a_n11634_10845.n87 a_n11634_10845.n85 0.758076
R14904 a_n11634_10845.n85 a_n11634_10845.n83 0.758076
R14905 a_n11634_10845.n83 a_n11634_10845.n81 0.758076
R14906 a_n11634_10845.n81 a_n11634_10845.n79 0.758076
R14907 a_n11634_10845.n79 a_n11634_10845.n77 0.758076
R14908 a_n11634_10845.n74 a_n11634_10845.n72 0.758076
R14909 a_n11634_10845.n72 a_n11634_10845.n70 0.758076
R14910 a_n11634_10845.n70 a_n11634_10845.n69 0.758076
R14911 a_n11634_10845.n69 a_n11634_10845.n67 0.758076
R14912 a_n11634_10845.n67 a_n11634_10845.n65 0.758076
R14913 a_n11634_10845.n65 a_n11634_10845.n64 0.758076
R14914 a_n11634_10845.n64 a_n11634_10845.n62 0.758076
R14915 a_n11634_10845.n62 a_n11634_10845.n60 0.758076
R14916 a_n11634_10845.n60 a_n11634_10845.n58 0.758076
R14917 a_n11634_10845.n58 a_n11634_10845.n56 0.758076
R14918 a_n11634_10845.n56 a_n11634_10845.n54 0.758076
R14919 a_n11634_10845.n54 a_n11634_10845.n52 0.758076
R14920 a_n11634_10845.n49 a_n11634_10845.n47 0.758076
R14921 a_n11634_10845.n47 a_n11634_10845.n45 0.758076
R14922 a_n11634_10845.n45 a_n11634_10845.n44 0.758076
R14923 a_n11634_10845.n44 a_n11634_10845.n42 0.758076
R14924 a_n11634_10845.n42 a_n11634_10845.n40 0.758076
R14925 a_n11634_10845.n40 a_n11634_10845.n39 0.758076
R14926 a_n11634_10845.n39 a_n11634_10845.n37 0.758076
R14927 a_n11634_10845.n37 a_n11634_10845.n35 0.758076
R14928 a_n11634_10845.n35 a_n11634_10845.n33 0.758076
R14929 a_n11634_10845.n33 a_n11634_10845.n31 0.758076
R14930 a_n11634_10845.n31 a_n11634_10845.n29 0.758076
R14931 a_n11634_10845.n29 a_n11634_10845.n27 0.758076
R14932 a_n11634_10845.n18 a_n11634_10845.n22 0.758076
R14933 a_n11634_10845.n22 a_n11634_10845.n24 0.568682
R14934 a_n11634_10845.n135 a_n11634_10845.n99 0.503145
R14935 a_n11634_10845.n129 a_n11634_10845.n74 0.503145
R14936 a_n11634_10845.n153 a_n11634_10845.n49 0.503145
R14937 a_n11634_10845.n24 a_n11634_10845.n113 0.503145
R14938 a_n11634_10845.n11 a_n11634_10845.n146 52.1509
R14939 a_n11634_10845.n12 a_n11634_10845.n145 52.1509
R14940 a_n11634_10845.n13 a_n11634_10845.n144 52.1509
R14941 a_n11634_10845.n143 a_n11634_10845.n21 21.6394
R14942 a_n11634_10845.n20 a_n11634_10845.t40 11.0881
R14943 a_n11634_10845.n9 a_n11634_10845.n16 4.14275
R14944 a_n11634_10845.n14 a_n11634_10845.n18 3.78838
R14945 a_n11634_10845.n6 a_n11634_10845.n11 2.96445
R14946 a_n11634_10845.n3 a_n11634_10845.n12 2.96445
R14947 a_n11634_10845.n0 a_n11634_10845.n13 2.96445
R14948 a_n11634_10845.n14 a_n11634_10845.n19 2.9529
R14949 a_n11778_11043.n2 a_n11778_11043.t7 176.341
R14950 a_n11778_11043.n3 a_n11778_11043.t8 175.29
R14951 a_n11778_11043.n0 a_n11778_11043.t13 156.754
R14952 a_n11778_11043.n1 a_n11778_11043.t14 154.892
R14953 a_n11778_11043.n0 a_n11778_11043.t0 154.892
R14954 a_n11778_11043.n0 a_n11778_11043.t16 154.892
R14955 a_n11778_11043.n2 a_n11778_11043.n4 149.084
R14956 a_n11778_11043.n3 a_n11778_11043.n6 149.084
R14957 a_n11778_11043.n3 a_n11778_11043.n5 149.084
R14958 a_n11778_11043.n10 a_n11778_11043.n2 149.084
R14959 a_n11778_11043.n1 a_n11778_11043.n8 129.496
R14960 a_n11778_11043.n0 a_n11778_11043.n7 129.496
R14961 a_n11778_11043.n4 a_n11778_11043.t9 25.395
R14962 a_n11778_11043.n4 a_n11778_11043.t11 25.395
R14963 a_n11778_11043.n8 a_n11778_11043.t15 25.395
R14964 a_n11778_11043.n8 a_n11778_11043.t2 25.395
R14965 a_n11778_11043.n7 a_n11778_11043.t1 25.395
R14966 a_n11778_11043.n7 a_n11778_11043.t17 25.395
R14967 a_n11778_11043.n6 a_n11778_11043.t6 25.395
R14968 a_n11778_11043.n6 a_n11778_11043.t5 25.395
R14969 a_n11778_11043.n5 a_n11778_11043.t10 25.395
R14970 a_n11778_11043.n5 a_n11778_11043.t4 25.395
R14971 a_n11778_11043.n10 a_n11778_11043.t3 25.395
R14972 a_n11778_11043.t12 a_n11778_11043.n10 25.395
R14973 a_n11778_11043.n9 a_n11778_11043.n3 19.251
R14974 a_n11778_11043.n2 a_n11778_11043.n9 14.4902
R14975 a_n11778_11043.n1 a_n11778_11043.n0 6.03498
R14976 a_n11778_11043.n9 a_n11778_11043.n1 5.8403
R14977 VDD.n4076 VDD.n95 455.123
R14978 VDD.n4484 VDD.n4259 455.123
R14979 VDD.n4380 VDD.n4367 455.123
R14980 VDD.n127 VDD.n93 455.123
R14981 VDD.n1803 VDD.n1233 455.123
R14982 VDD.n1806 VDD.n1805 455.123
R14983 VDD.n1586 VDD.n1373 455.123
R14984 VDD.n1588 VDD.n1371 455.123
R14985 VDD.n3924 VDD.n190 276.586
R14986 VDD.n3890 VDD.n187 276.586
R14987 VDD.n3388 VDD.n2910 276.586
R14988 VDD.n3423 VDD.n633 276.586
R14989 VDD.n2858 VDD.n670 276.586
R14990 VDD.n2824 VDD.n2823 276.586
R14991 VDD.n1933 VDD.n1103 276.586
R14992 VDD.n2387 VDD.n1101 276.586
R14993 VDD.n3869 VDD.n188 276.586
R14994 VDD.n3927 VDD.n3926 276.586
R14995 VDD.n3152 VDD.n3151 276.586
R14996 VDD.n3427 VDD.n637 276.586
R14997 VDD.n2901 VDD.n659 276.586
R14998 VDD.n2865 VDD.n658 276.586
R14999 VDD.n1117 VDD.n1104 276.586
R15000 VDD.n2385 VDD.n1105 276.586
R15001 VDD.n1376 VDD.t6 263.938
R15002 VDD.n1390 VDD.t58 263.938
R15003 VDD.n1407 VDD.t3 263.938
R15004 VDD.n1421 VDD.t9 263.938
R15005 VDD.n1438 VDD.t16 263.938
R15006 VDD.n1142 VDD.t90 263.938
R15007 VDD.n1225 VDD.t34 263.938
R15008 VDD.n1202 VDD.t75 263.938
R15009 VDD.n1182 VDD.t72 263.938
R15010 VDD.n1161 VDD.t84 263.938
R15011 VDD.n4363 VDD.t44 263.938
R15012 VDD.n4342 VDD.t87 263.938
R15013 VDD.n4322 VDD.t54 263.938
R15014 VDD.n4301 VDD.t60 263.938
R15015 VDD.n4278 VDD.t66 263.938
R15016 VDD.n137 VDD.t48 263.938
R15017 VDD.n159 VDD.t27 263.938
R15018 VDD.n3944 VDD.t13 263.938
R15019 VDD.n4033 VDD.t38 263.938
R15020 VDD.n3964 VDD.t64 263.938
R15021 VDD.n1114 VDD.t24 261.899
R15022 VDD.n662 VDD.t30 261.899
R15023 VDD.n1134 VDD.t82 261.899
R15024 VDD.n672 VDD.t40 261.899
R15025 VDD.n3117 VDD.t79 261.899
R15026 VDD.n201 VDD.t69 261.899
R15027 VDD.n2921 VDD.t52 261.899
R15028 VDD.n177 VDD.t19 261.899
R15029 VDD.t147 VDD.t112 237.65
R15030 VDD.t105 VDD.t134 237.65
R15031 VDD.n1146 VDD.t147 229.379
R15032 VDD.n4074 VDD.t134 229.379
R15033 VDD.n1376 VDD.t4 210.637
R15034 VDD.n1390 VDD.t56 210.637
R15035 VDD.n1407 VDD.t0 210.637
R15036 VDD.n1421 VDD.t7 210.637
R15037 VDD.n1438 VDD.t14 210.637
R15038 VDD.n1142 VDD.t89 210.637
R15039 VDD.n1225 VDD.t32 210.637
R15040 VDD.n1202 VDD.t74 210.637
R15041 VDD.n1182 VDD.t71 210.637
R15042 VDD.n1161 VDD.t83 210.637
R15043 VDD.n4363 VDD.t42 210.637
R15044 VDD.n4342 VDD.t86 210.637
R15045 VDD.n4322 VDD.t53 210.637
R15046 VDD.n4301 VDD.t59 210.637
R15047 VDD.n4278 VDD.t65 210.637
R15048 VDD.n137 VDD.t46 210.637
R15049 VDD.n159 VDD.t25 210.637
R15050 VDD.n3944 VDD.t10 210.637
R15051 VDD.n4033 VDD.t36 210.637
R15052 VDD.n3964 VDD.t62 210.637
R15053 VDD.n1114 VDD.t21 210.595
R15054 VDD.n662 VDD.t28 210.595
R15055 VDD.n1134 VDD.t80 210.595
R15056 VDD.n672 VDD.t39 210.595
R15057 VDD.n3117 VDD.t77 210.595
R15058 VDD.n201 VDD.t68 210.595
R15059 VDD.n2921 VDD.t49 210.595
R15060 VDD.n177 VDD.t17 210.595
R15061 VDD.n3871 VDD.n188 185
R15062 VDD.n3925 VDD.n188 185
R15063 VDD.n3873 VDD.n3872 185
R15064 VDD.n3872 VDD.n186 185
R15065 VDD.n3874 VDD.n211 185
R15066 VDD.n3884 VDD.n211 185
R15067 VDD.n3875 VDD.n219 185
R15068 VDD.n219 VDD.n209 185
R15069 VDD.n3877 VDD.n3876 185
R15070 VDD.n3878 VDD.n3877 185
R15071 VDD.n3849 VDD.n218 185
R15072 VDD.n218 VDD.n215 185
R15073 VDD.n3848 VDD.n3847 185
R15074 VDD.n3847 VDD.n3846 185
R15075 VDD.n221 VDD.n220 185
R15076 VDD.n222 VDD.n221 185
R15077 VDD.n3839 VDD.n3838 185
R15078 VDD.n3840 VDD.n3839 185
R15079 VDD.n3837 VDD.n230 185
R15080 VDD.n236 VDD.n230 185
R15081 VDD.n3836 VDD.n3835 185
R15082 VDD.n3835 VDD.n3834 185
R15083 VDD.n232 VDD.n231 185
R15084 VDD.n233 VDD.n232 185
R15085 VDD.n3827 VDD.n3826 185
R15086 VDD.n3828 VDD.n3827 185
R15087 VDD.n3825 VDD.n243 185
R15088 VDD.n243 VDD.n240 185
R15089 VDD.n3824 VDD.n3823 185
R15090 VDD.n3823 VDD.n3822 185
R15091 VDD.n245 VDD.n244 185
R15092 VDD.n246 VDD.n245 185
R15093 VDD.n3815 VDD.n3814 185
R15094 VDD.n3816 VDD.n3815 185
R15095 VDD.n3813 VDD.n255 185
R15096 VDD.n255 VDD.n252 185
R15097 VDD.n3812 VDD.n3811 185
R15098 VDD.n3811 VDD.n3810 185
R15099 VDD.n257 VDD.n256 185
R15100 VDD.n258 VDD.n257 185
R15101 VDD.n3803 VDD.n3802 185
R15102 VDD.n3804 VDD.n3803 185
R15103 VDD.n3801 VDD.n267 185
R15104 VDD.n267 VDD.n264 185
R15105 VDD.n3800 VDD.n3799 185
R15106 VDD.n3799 VDD.n3798 185
R15107 VDD.n269 VDD.n268 185
R15108 VDD.n270 VDD.n269 185
R15109 VDD.n3791 VDD.n3790 185
R15110 VDD.n3792 VDD.n3791 185
R15111 VDD.n3789 VDD.n279 185
R15112 VDD.n279 VDD.n276 185
R15113 VDD.n3788 VDD.n3787 185
R15114 VDD.n3787 VDD.n3786 185
R15115 VDD.n281 VDD.n280 185
R15116 VDD.n282 VDD.n281 185
R15117 VDD.n3779 VDD.n3778 185
R15118 VDD.n3780 VDD.n3779 185
R15119 VDD.n3777 VDD.n291 185
R15120 VDD.n291 VDD.n288 185
R15121 VDD.n3776 VDD.n3775 185
R15122 VDD.n3775 VDD.n3774 185
R15123 VDD.n293 VDD.n292 185
R15124 VDD.n294 VDD.n293 185
R15125 VDD.n3767 VDD.n3766 185
R15126 VDD.n3768 VDD.n3767 185
R15127 VDD.n3765 VDD.n303 185
R15128 VDD.n303 VDD.n300 185
R15129 VDD.n3764 VDD.n3763 185
R15130 VDD.n3763 VDD.n3762 185
R15131 VDD.n305 VDD.n304 185
R15132 VDD.n314 VDD.n305 185
R15133 VDD.n3755 VDD.n3754 185
R15134 VDD.n3756 VDD.n3755 185
R15135 VDD.n3753 VDD.n315 185
R15136 VDD.n315 VDD.n311 185
R15137 VDD.n3752 VDD.n3751 185
R15138 VDD.n3751 VDD.n3750 185
R15139 VDD.n317 VDD.n316 185
R15140 VDD.n318 VDD.n317 185
R15141 VDD.n3743 VDD.n3742 185
R15142 VDD.n3744 VDD.n3743 185
R15143 VDD.n3741 VDD.n327 185
R15144 VDD.n327 VDD.n324 185
R15145 VDD.n3740 VDD.n3739 185
R15146 VDD.n3739 VDD.n3738 185
R15147 VDD.n329 VDD.n328 185
R15148 VDD.n330 VDD.n329 185
R15149 VDD.n3731 VDD.n3730 185
R15150 VDD.n3732 VDD.n3731 185
R15151 VDD.n3729 VDD.n339 185
R15152 VDD.n339 VDD.n336 185
R15153 VDD.n3728 VDD.n3727 185
R15154 VDD.n3727 VDD.n3726 185
R15155 VDD.n341 VDD.n340 185
R15156 VDD.n350 VDD.n341 185
R15157 VDD.n3719 VDD.n3718 185
R15158 VDD.n3720 VDD.n3719 185
R15159 VDD.n3717 VDD.n351 185
R15160 VDD.n351 VDD.n347 185
R15161 VDD.n3716 VDD.n3715 185
R15162 VDD.n3715 VDD.n3714 185
R15163 VDD.n353 VDD.n352 185
R15164 VDD.n354 VDD.n353 185
R15165 VDD.n3707 VDD.n3706 185
R15166 VDD.n3708 VDD.n3707 185
R15167 VDD.n3705 VDD.n363 185
R15168 VDD.n363 VDD.n360 185
R15169 VDD.n3704 VDD.n3703 185
R15170 VDD.n3703 VDD.n3702 185
R15171 VDD.n365 VDD.n364 185
R15172 VDD.n366 VDD.n365 185
R15173 VDD.n3695 VDD.n3694 185
R15174 VDD.n3696 VDD.n3695 185
R15175 VDD.n3693 VDD.n375 185
R15176 VDD.n375 VDD.n372 185
R15177 VDD.n3692 VDD.n3691 185
R15178 VDD.n3691 VDD.n3690 185
R15179 VDD.n377 VDD.n376 185
R15180 VDD.n378 VDD.n377 185
R15181 VDD.n3683 VDD.n3682 185
R15182 VDD.n3684 VDD.n3683 185
R15183 VDD.n3681 VDD.n387 185
R15184 VDD.n387 VDD.n384 185
R15185 VDD.n3680 VDD.n3679 185
R15186 VDD.n3679 VDD.n3678 185
R15187 VDD.n389 VDD.n388 185
R15188 VDD.n390 VDD.n389 185
R15189 VDD.n3671 VDD.n3670 185
R15190 VDD.n3672 VDD.n3671 185
R15191 VDD.n3669 VDD.n399 185
R15192 VDD.n399 VDD.n396 185
R15193 VDD.n3668 VDD.n3667 185
R15194 VDD.n3667 VDD.n3666 185
R15195 VDD.n401 VDD.n400 185
R15196 VDD.n402 VDD.n401 185
R15197 VDD.n3659 VDD.n3658 185
R15198 VDD.n3660 VDD.n3659 185
R15199 VDD.n3657 VDD.n411 185
R15200 VDD.n411 VDD.n408 185
R15201 VDD.n3656 VDD.n3655 185
R15202 VDD.n3655 VDD.n3654 185
R15203 VDD.n413 VDD.n412 185
R15204 VDD.n414 VDD.n413 185
R15205 VDD.n3647 VDD.n3646 185
R15206 VDD.n3648 VDD.n3647 185
R15207 VDD.n3645 VDD.n422 185
R15208 VDD.n427 VDD.n422 185
R15209 VDD.n3644 VDD.n3643 185
R15210 VDD.n3643 VDD.n3642 185
R15211 VDD.n424 VDD.n423 185
R15212 VDD.t132 VDD.n424 185
R15213 VDD.n3635 VDD.n3634 185
R15214 VDD.n3636 VDD.n3635 185
R15215 VDD.n3633 VDD.n434 185
R15216 VDD.n434 VDD.n431 185
R15217 VDD.n3632 VDD.n3631 185
R15218 VDD.n3631 VDD.n3630 185
R15219 VDD.n436 VDD.n435 185
R15220 VDD.n437 VDD.n436 185
R15221 VDD.n3623 VDD.n3622 185
R15222 VDD.n3624 VDD.n3623 185
R15223 VDD.n3621 VDD.n446 185
R15224 VDD.n446 VDD.n443 185
R15225 VDD.n3620 VDD.n3619 185
R15226 VDD.n3619 VDD.n3618 185
R15227 VDD.n448 VDD.n447 185
R15228 VDD.n449 VDD.n448 185
R15229 VDD.n3611 VDD.n3610 185
R15230 VDD.n3612 VDD.n3611 185
R15231 VDD.n3609 VDD.n458 185
R15232 VDD.n458 VDD.n455 185
R15233 VDD.n3608 VDD.n3607 185
R15234 VDD.n3607 VDD.n3606 185
R15235 VDD.n460 VDD.n459 185
R15236 VDD.n461 VDD.n460 185
R15237 VDD.n3599 VDD.n3598 185
R15238 VDD.n3600 VDD.n3599 185
R15239 VDD.n3597 VDD.n470 185
R15240 VDD.n470 VDD.n467 185
R15241 VDD.n3596 VDD.n3595 185
R15242 VDD.n3595 VDD.n3594 185
R15243 VDD.n472 VDD.n471 185
R15244 VDD.n473 VDD.n472 185
R15245 VDD.n3587 VDD.n3586 185
R15246 VDD.n3588 VDD.n3587 185
R15247 VDD.n3585 VDD.n482 185
R15248 VDD.n482 VDD.n479 185
R15249 VDD.n3584 VDD.n3583 185
R15250 VDD.n3583 VDD.n3582 185
R15251 VDD.n484 VDD.n483 185
R15252 VDD.n493 VDD.n484 185
R15253 VDD.n3575 VDD.n3574 185
R15254 VDD.n3576 VDD.n3575 185
R15255 VDD.n3573 VDD.n494 185
R15256 VDD.n494 VDD.n490 185
R15257 VDD.n3572 VDD.n3571 185
R15258 VDD.n3571 VDD.n3570 185
R15259 VDD.n496 VDD.n495 185
R15260 VDD.n497 VDD.n496 185
R15261 VDD.n3563 VDD.n3562 185
R15262 VDD.n3564 VDD.n3563 185
R15263 VDD.n3561 VDD.n506 185
R15264 VDD.n506 VDD.n503 185
R15265 VDD.n3560 VDD.n3559 185
R15266 VDD.n3559 VDD.n3558 185
R15267 VDD.n508 VDD.n507 185
R15268 VDD.n509 VDD.n508 185
R15269 VDD.n3551 VDD.n3550 185
R15270 VDD.n3552 VDD.n3551 185
R15271 VDD.n3549 VDD.n518 185
R15272 VDD.n518 VDD.n515 185
R15273 VDD.n3548 VDD.n3547 185
R15274 VDD.n3547 VDD.n3546 185
R15275 VDD.n520 VDD.n519 185
R15276 VDD.n521 VDD.n520 185
R15277 VDD.n3539 VDD.n3538 185
R15278 VDD.n3540 VDD.n3539 185
R15279 VDD.n3537 VDD.n530 185
R15280 VDD.n530 VDD.n527 185
R15281 VDD.n3536 VDD.n3535 185
R15282 VDD.n3535 VDD.n3534 185
R15283 VDD.n532 VDD.n531 185
R15284 VDD.n541 VDD.n532 185
R15285 VDD.n3527 VDD.n3526 185
R15286 VDD.n3528 VDD.n3527 185
R15287 VDD.n3525 VDD.n542 185
R15288 VDD.n542 VDD.n538 185
R15289 VDD.n3524 VDD.n3523 185
R15290 VDD.n3523 VDD.n3522 185
R15291 VDD.n544 VDD.n543 185
R15292 VDD.n545 VDD.n544 185
R15293 VDD.n3515 VDD.n3514 185
R15294 VDD.n3516 VDD.n3515 185
R15295 VDD.n3513 VDD.n554 185
R15296 VDD.n554 VDD.n551 185
R15297 VDD.n3512 VDD.n3511 185
R15298 VDD.n3511 VDD.n3510 185
R15299 VDD.n556 VDD.n555 185
R15300 VDD.n557 VDD.n556 185
R15301 VDD.n3503 VDD.n3502 185
R15302 VDD.n3504 VDD.n3503 185
R15303 VDD.n3501 VDD.n566 185
R15304 VDD.n566 VDD.n563 185
R15305 VDD.n3500 VDD.n3499 185
R15306 VDD.n3499 VDD.n3498 185
R15307 VDD.n568 VDD.n567 185
R15308 VDD.n569 VDD.n568 185
R15309 VDD.n3491 VDD.n3490 185
R15310 VDD.n3492 VDD.n3491 185
R15311 VDD.n3489 VDD.n578 185
R15312 VDD.n578 VDD.n575 185
R15313 VDD.n3488 VDD.n3487 185
R15314 VDD.n3487 VDD.n3486 185
R15315 VDD.n580 VDD.n579 185
R15316 VDD.n581 VDD.n580 185
R15317 VDD.n3479 VDD.n3478 185
R15318 VDD.n3480 VDD.n3479 185
R15319 VDD.n3477 VDD.n590 185
R15320 VDD.n590 VDD.n587 185
R15321 VDD.n3476 VDD.n3475 185
R15322 VDD.n3475 VDD.n3474 185
R15323 VDD.n592 VDD.n591 185
R15324 VDD.n593 VDD.n592 185
R15325 VDD.n3467 VDD.n3466 185
R15326 VDD.n3468 VDD.n3467 185
R15327 VDD.n3465 VDD.n601 185
R15328 VDD.n3369 VDD.n601 185
R15329 VDD.n3464 VDD.n3463 185
R15330 VDD.n3463 VDD.n3462 185
R15331 VDD.n603 VDD.n602 185
R15332 VDD.n604 VDD.n603 185
R15333 VDD.n3455 VDD.n3454 185
R15334 VDD.n3456 VDD.n3455 185
R15335 VDD.n3453 VDD.n613 185
R15336 VDD.n613 VDD.n610 185
R15337 VDD.n3452 VDD.n3451 185
R15338 VDD.n3451 VDD.n3450 185
R15339 VDD.n615 VDD.n614 185
R15340 VDD.n616 VDD.n615 185
R15341 VDD.n3443 VDD.n3442 185
R15342 VDD.n3444 VDD.n3443 185
R15343 VDD.n3441 VDD.n625 185
R15344 VDD.n625 VDD.n622 185
R15345 VDD.n3440 VDD.n3439 185
R15346 VDD.n3439 VDD.n3438 185
R15347 VDD.n627 VDD.n626 185
R15348 VDD.n628 VDD.n627 185
R15349 VDD.n3431 VDD.n3430 185
R15350 VDD.n3432 VDD.n3431 185
R15351 VDD.n3429 VDD.n637 185
R15352 VDD.n637 VDD.n634 185
R15353 VDD.n3428 VDD.n3427 185
R15354 VDD.n639 VDD.n638 185
R15355 VDD.n3121 VDD.n3120 185
R15356 VDD.n3123 VDD.n3122 185
R15357 VDD.n3125 VDD.n3124 185
R15358 VDD.n3127 VDD.n3126 185
R15359 VDD.n3129 VDD.n3128 185
R15360 VDD.n3131 VDD.n3130 185
R15361 VDD.n3133 VDD.n3132 185
R15362 VDD.n3135 VDD.n3134 185
R15363 VDD.n3137 VDD.n3136 185
R15364 VDD.n3139 VDD.n3138 185
R15365 VDD.n3141 VDD.n3140 185
R15366 VDD.n3143 VDD.n3142 185
R15367 VDD.n3145 VDD.n3144 185
R15368 VDD.n3147 VDD.n3146 185
R15369 VDD.n3149 VDD.n3148 185
R15370 VDD.n3151 VDD.n3150 185
R15371 VDD.n3928 VDD.n3927 185
R15372 VDD.n3929 VDD.n182 185
R15373 VDD.n3931 VDD.n3930 185
R15374 VDD.n3933 VDD.n181 185
R15375 VDD.n3935 VDD.n3934 185
R15376 VDD.n3936 VDD.n176 185
R15377 VDD.n3938 VDD.n3937 185
R15378 VDD.n3940 VDD.n173 185
R15379 VDD.n3942 VDD.n3941 185
R15380 VDD.n3855 VDD.n172 185
R15381 VDD.n3857 VDD.n3856 185
R15382 VDD.n3859 VDD.n3853 185
R15383 VDD.n3861 VDD.n3860 185
R15384 VDD.n3862 VDD.n3852 185
R15385 VDD.n3864 VDD.n3863 185
R15386 VDD.n3866 VDD.n3851 185
R15387 VDD.n3867 VDD.n3850 185
R15388 VDD.n3870 VDD.n3869 185
R15389 VDD.n3926 VDD.n183 185
R15390 VDD.n3926 VDD.n3925 185
R15391 VDD.n3170 VDD.n185 185
R15392 VDD.n186 VDD.n185 185
R15393 VDD.n3171 VDD.n210 185
R15394 VDD.n3884 VDD.n210 185
R15395 VDD.n3173 VDD.n3172 185
R15396 VDD.n3172 VDD.n209 185
R15397 VDD.n3174 VDD.n217 185
R15398 VDD.n3878 VDD.n217 185
R15399 VDD.n3176 VDD.n3175 185
R15400 VDD.n3175 VDD.n215 185
R15401 VDD.n3177 VDD.n224 185
R15402 VDD.n3846 VDD.n224 185
R15403 VDD.n3179 VDD.n3178 185
R15404 VDD.n3178 VDD.n222 185
R15405 VDD.n3180 VDD.n229 185
R15406 VDD.n3840 VDD.n229 185
R15407 VDD.n3182 VDD.n3181 185
R15408 VDD.n3181 VDD.n236 185
R15409 VDD.n3183 VDD.n235 185
R15410 VDD.n3834 VDD.n235 185
R15411 VDD.n3185 VDD.n3184 185
R15412 VDD.n3184 VDD.n233 185
R15413 VDD.n3186 VDD.n242 185
R15414 VDD.n3828 VDD.n242 185
R15415 VDD.n3188 VDD.n3187 185
R15416 VDD.n3187 VDD.n240 185
R15417 VDD.n3189 VDD.n248 185
R15418 VDD.n3822 VDD.n248 185
R15419 VDD.n3191 VDD.n3190 185
R15420 VDD.n3190 VDD.n246 185
R15421 VDD.n3192 VDD.n254 185
R15422 VDD.n3816 VDD.n254 185
R15423 VDD.n3194 VDD.n3193 185
R15424 VDD.n3193 VDD.n252 185
R15425 VDD.n3195 VDD.n260 185
R15426 VDD.n3810 VDD.n260 185
R15427 VDD.n3197 VDD.n3196 185
R15428 VDD.n3196 VDD.n258 185
R15429 VDD.n3198 VDD.n266 185
R15430 VDD.n3804 VDD.n266 185
R15431 VDD.n3200 VDD.n3199 185
R15432 VDD.n3199 VDD.n264 185
R15433 VDD.n3201 VDD.n272 185
R15434 VDD.n3798 VDD.n272 185
R15435 VDD.n3203 VDD.n3202 185
R15436 VDD.n3202 VDD.n270 185
R15437 VDD.n3204 VDD.n278 185
R15438 VDD.n3792 VDD.n278 185
R15439 VDD.n3206 VDD.n3205 185
R15440 VDD.n3205 VDD.n276 185
R15441 VDD.n3207 VDD.n284 185
R15442 VDD.n3786 VDD.n284 185
R15443 VDD.n3209 VDD.n3208 185
R15444 VDD.n3208 VDD.n282 185
R15445 VDD.n3210 VDD.n290 185
R15446 VDD.n3780 VDD.n290 185
R15447 VDD.n3212 VDD.n3211 185
R15448 VDD.n3211 VDD.n288 185
R15449 VDD.n3213 VDD.n296 185
R15450 VDD.n3774 VDD.n296 185
R15451 VDD.n3215 VDD.n3214 185
R15452 VDD.n3214 VDD.n294 185
R15453 VDD.n3216 VDD.n302 185
R15454 VDD.n3768 VDD.n302 185
R15455 VDD.n3218 VDD.n3217 185
R15456 VDD.n3217 VDD.n300 185
R15457 VDD.n3219 VDD.n307 185
R15458 VDD.n3762 VDD.n307 185
R15459 VDD.n3221 VDD.n3220 185
R15460 VDD.n3220 VDD.n314 185
R15461 VDD.n3222 VDD.n313 185
R15462 VDD.n3756 VDD.n313 185
R15463 VDD.n3224 VDD.n3223 185
R15464 VDD.n3223 VDD.n311 185
R15465 VDD.n3225 VDD.n320 185
R15466 VDD.n3750 VDD.n320 185
R15467 VDD.n3227 VDD.n3226 185
R15468 VDD.n3226 VDD.n318 185
R15469 VDD.n3228 VDD.n326 185
R15470 VDD.n3744 VDD.n326 185
R15471 VDD.n3230 VDD.n3229 185
R15472 VDD.n3229 VDD.n324 185
R15473 VDD.n3231 VDD.n332 185
R15474 VDD.n3738 VDD.n332 185
R15475 VDD.n3233 VDD.n3232 185
R15476 VDD.n3232 VDD.n330 185
R15477 VDD.n3234 VDD.n338 185
R15478 VDD.n3732 VDD.n338 185
R15479 VDD.n3236 VDD.n3235 185
R15480 VDD.n3235 VDD.n336 185
R15481 VDD.n3237 VDD.n343 185
R15482 VDD.n3726 VDD.n343 185
R15483 VDD.n3239 VDD.n3238 185
R15484 VDD.n3238 VDD.n350 185
R15485 VDD.n3240 VDD.n349 185
R15486 VDD.n3720 VDD.n349 185
R15487 VDD.n3242 VDD.n3241 185
R15488 VDD.n3241 VDD.n347 185
R15489 VDD.n3243 VDD.n356 185
R15490 VDD.n3714 VDD.n356 185
R15491 VDD.n3245 VDD.n3244 185
R15492 VDD.n3244 VDD.n354 185
R15493 VDD.n3246 VDD.n362 185
R15494 VDD.n3708 VDD.n362 185
R15495 VDD.n3248 VDD.n3247 185
R15496 VDD.n3247 VDD.n360 185
R15497 VDD.n3249 VDD.n368 185
R15498 VDD.n3702 VDD.n368 185
R15499 VDD.n3251 VDD.n3250 185
R15500 VDD.n3250 VDD.n366 185
R15501 VDD.n3252 VDD.n374 185
R15502 VDD.n3696 VDD.n374 185
R15503 VDD.n3254 VDD.n3253 185
R15504 VDD.n3253 VDD.n372 185
R15505 VDD.n3255 VDD.n380 185
R15506 VDD.n3690 VDD.n380 185
R15507 VDD.n3257 VDD.n3256 185
R15508 VDD.n3256 VDD.n378 185
R15509 VDD.n3258 VDD.n386 185
R15510 VDD.n3684 VDD.n386 185
R15511 VDD.n3260 VDD.n3259 185
R15512 VDD.n3259 VDD.n384 185
R15513 VDD.n3261 VDD.n392 185
R15514 VDD.n3678 VDD.n392 185
R15515 VDD.n3263 VDD.n3262 185
R15516 VDD.n3262 VDD.n390 185
R15517 VDD.n3264 VDD.n398 185
R15518 VDD.n3672 VDD.n398 185
R15519 VDD.n3266 VDD.n3265 185
R15520 VDD.n3265 VDD.n396 185
R15521 VDD.n3267 VDD.n404 185
R15522 VDD.n3666 VDD.n404 185
R15523 VDD.n3269 VDD.n3268 185
R15524 VDD.n3268 VDD.n402 185
R15525 VDD.n3270 VDD.n410 185
R15526 VDD.n3660 VDD.n410 185
R15527 VDD.n3272 VDD.n3271 185
R15528 VDD.n3271 VDD.n408 185
R15529 VDD.n3273 VDD.n416 185
R15530 VDD.n3654 VDD.n416 185
R15531 VDD.n3275 VDD.n3274 185
R15532 VDD.n3274 VDD.n414 185
R15533 VDD.n3276 VDD.n421 185
R15534 VDD.n3648 VDD.n421 185
R15535 VDD.n3278 VDD.n3277 185
R15536 VDD.n3277 VDD.n427 185
R15537 VDD.n3279 VDD.n426 185
R15538 VDD.n3642 VDD.n426 185
R15539 VDD.n3281 VDD.n3280 185
R15540 VDD.n3280 VDD.t132 185
R15541 VDD.n3282 VDD.n433 185
R15542 VDD.n3636 VDD.n433 185
R15543 VDD.n3284 VDD.n3283 185
R15544 VDD.n3283 VDD.n431 185
R15545 VDD.n3285 VDD.n439 185
R15546 VDD.n3630 VDD.n439 185
R15547 VDD.n3287 VDD.n3286 185
R15548 VDD.n3286 VDD.n437 185
R15549 VDD.n3288 VDD.n445 185
R15550 VDD.n3624 VDD.n445 185
R15551 VDD.n3290 VDD.n3289 185
R15552 VDD.n3289 VDD.n443 185
R15553 VDD.n3291 VDD.n451 185
R15554 VDD.n3618 VDD.n451 185
R15555 VDD.n3293 VDD.n3292 185
R15556 VDD.n3292 VDD.n449 185
R15557 VDD.n3294 VDD.n457 185
R15558 VDD.n3612 VDD.n457 185
R15559 VDD.n3296 VDD.n3295 185
R15560 VDD.n3295 VDD.n455 185
R15561 VDD.n3297 VDD.n463 185
R15562 VDD.n3606 VDD.n463 185
R15563 VDD.n3299 VDD.n3298 185
R15564 VDD.n3298 VDD.n461 185
R15565 VDD.n3300 VDD.n469 185
R15566 VDD.n3600 VDD.n469 185
R15567 VDD.n3302 VDD.n3301 185
R15568 VDD.n3301 VDD.n467 185
R15569 VDD.n3303 VDD.n475 185
R15570 VDD.n3594 VDD.n475 185
R15571 VDD.n3305 VDD.n3304 185
R15572 VDD.n3304 VDD.n473 185
R15573 VDD.n3306 VDD.n481 185
R15574 VDD.n3588 VDD.n481 185
R15575 VDD.n3308 VDD.n3307 185
R15576 VDD.n3307 VDD.n479 185
R15577 VDD.n3309 VDD.n486 185
R15578 VDD.n3582 VDD.n486 185
R15579 VDD.n3311 VDD.n3310 185
R15580 VDD.n3310 VDD.n493 185
R15581 VDD.n3312 VDD.n492 185
R15582 VDD.n3576 VDD.n492 185
R15583 VDD.n3314 VDD.n3313 185
R15584 VDD.n3313 VDD.n490 185
R15585 VDD.n3315 VDD.n499 185
R15586 VDD.n3570 VDD.n499 185
R15587 VDD.n3317 VDD.n3316 185
R15588 VDD.n3316 VDD.n497 185
R15589 VDD.n3318 VDD.n505 185
R15590 VDD.n3564 VDD.n505 185
R15591 VDD.n3320 VDD.n3319 185
R15592 VDD.n3319 VDD.n503 185
R15593 VDD.n3321 VDD.n511 185
R15594 VDD.n3558 VDD.n511 185
R15595 VDD.n3323 VDD.n3322 185
R15596 VDD.n3322 VDD.n509 185
R15597 VDD.n3324 VDD.n517 185
R15598 VDD.n3552 VDD.n517 185
R15599 VDD.n3326 VDD.n3325 185
R15600 VDD.n3325 VDD.n515 185
R15601 VDD.n3327 VDD.n523 185
R15602 VDD.n3546 VDD.n523 185
R15603 VDD.n3329 VDD.n3328 185
R15604 VDD.n3328 VDD.n521 185
R15605 VDD.n3330 VDD.n529 185
R15606 VDD.n3540 VDD.n529 185
R15607 VDD.n3332 VDD.n3331 185
R15608 VDD.n3331 VDD.n527 185
R15609 VDD.n3333 VDD.n534 185
R15610 VDD.n3534 VDD.n534 185
R15611 VDD.n3335 VDD.n3334 185
R15612 VDD.n3334 VDD.n541 185
R15613 VDD.n3336 VDD.n540 185
R15614 VDD.n3528 VDD.n540 185
R15615 VDD.n3338 VDD.n3337 185
R15616 VDD.n3337 VDD.n538 185
R15617 VDD.n3339 VDD.n547 185
R15618 VDD.n3522 VDD.n547 185
R15619 VDD.n3341 VDD.n3340 185
R15620 VDD.n3340 VDD.n545 185
R15621 VDD.n3342 VDD.n553 185
R15622 VDD.n3516 VDD.n553 185
R15623 VDD.n3344 VDD.n3343 185
R15624 VDD.n3343 VDD.n551 185
R15625 VDD.n3345 VDD.n559 185
R15626 VDD.n3510 VDD.n559 185
R15627 VDD.n3347 VDD.n3346 185
R15628 VDD.n3346 VDD.n557 185
R15629 VDD.n3348 VDD.n565 185
R15630 VDD.n3504 VDD.n565 185
R15631 VDD.n3350 VDD.n3349 185
R15632 VDD.n3349 VDD.n563 185
R15633 VDD.n3351 VDD.n571 185
R15634 VDD.n3498 VDD.n571 185
R15635 VDD.n3353 VDD.n3352 185
R15636 VDD.n3352 VDD.n569 185
R15637 VDD.n3354 VDD.n577 185
R15638 VDD.n3492 VDD.n577 185
R15639 VDD.n3356 VDD.n3355 185
R15640 VDD.n3355 VDD.n575 185
R15641 VDD.n3357 VDD.n583 185
R15642 VDD.n3486 VDD.n583 185
R15643 VDD.n3359 VDD.n3358 185
R15644 VDD.n3358 VDD.n581 185
R15645 VDD.n3360 VDD.n589 185
R15646 VDD.n3480 VDD.n589 185
R15647 VDD.n3362 VDD.n3361 185
R15648 VDD.n3361 VDD.n587 185
R15649 VDD.n3363 VDD.n595 185
R15650 VDD.n3474 VDD.n595 185
R15651 VDD.n3365 VDD.n3364 185
R15652 VDD.n3364 VDD.n593 185
R15653 VDD.n3366 VDD.n600 185
R15654 VDD.n3468 VDD.n600 185
R15655 VDD.n3368 VDD.n3367 185
R15656 VDD.n3369 VDD.n3368 185
R15657 VDD.n3169 VDD.n606 185
R15658 VDD.n3462 VDD.n606 185
R15659 VDD.n3168 VDD.n3167 185
R15660 VDD.n3167 VDD.n604 185
R15661 VDD.n3166 VDD.n612 185
R15662 VDD.n3456 VDD.n612 185
R15663 VDD.n3165 VDD.n3164 185
R15664 VDD.n3164 VDD.n610 185
R15665 VDD.n3163 VDD.n618 185
R15666 VDD.n3450 VDD.n618 185
R15667 VDD.n3162 VDD.n3161 185
R15668 VDD.n3161 VDD.n616 185
R15669 VDD.n3160 VDD.n624 185
R15670 VDD.n3444 VDD.n624 185
R15671 VDD.n3159 VDD.n3158 185
R15672 VDD.n3158 VDD.n622 185
R15673 VDD.n3157 VDD.n630 185
R15674 VDD.n3438 VDD.n630 185
R15675 VDD.n3156 VDD.n3155 185
R15676 VDD.n3155 VDD.n628 185
R15677 VDD.n3154 VDD.n636 185
R15678 VDD.n3432 VDD.n636 185
R15679 VDD.n3153 VDD.n3152 185
R15680 VDD.n3152 VDD.n634 185
R15681 VDD.n2860 VDD.n670 185
R15682 VDD.n670 VDD.n640 185
R15683 VDD.n2862 VDD.n2861 185
R15684 VDD.n2863 VDD.n2862 185
R15685 VDD.n671 VDD.n669 185
R15686 VDD.n669 VDD.n666 185
R15687 VDD.n2816 VDD.n2815 185
R15688 VDD.n2817 VDD.n2816 185
R15689 VDD.n2814 VDD.n680 185
R15690 VDD.n680 VDD.n677 185
R15691 VDD.n2813 VDD.n2812 185
R15692 VDD.n2812 VDD.n2811 185
R15693 VDD.n682 VDD.n681 185
R15694 VDD.n683 VDD.n682 185
R15695 VDD.n2799 VDD.n2798 185
R15696 VDD.n2800 VDD.n2799 185
R15697 VDD.n2797 VDD.n693 185
R15698 VDD.n693 VDD.n690 185
R15699 VDD.n2796 VDD.n2795 185
R15700 VDD.n2795 VDD.n2794 185
R15701 VDD.n695 VDD.n694 185
R15702 VDD.n696 VDD.n695 185
R15703 VDD.n2787 VDD.n2786 185
R15704 VDD.n2788 VDD.n2787 185
R15705 VDD.n2785 VDD.n704 185
R15706 VDD.n2147 VDD.n704 185
R15707 VDD.n2784 VDD.n2783 185
R15708 VDD.n2783 VDD.n2782 185
R15709 VDD.n706 VDD.n705 185
R15710 VDD.n707 VDD.n706 185
R15711 VDD.n2775 VDD.n2774 185
R15712 VDD.n2776 VDD.n2775 185
R15713 VDD.n2773 VDD.n716 185
R15714 VDD.n716 VDD.n713 185
R15715 VDD.n2772 VDD.n2771 185
R15716 VDD.n2771 VDD.n2770 185
R15717 VDD.n718 VDD.n717 185
R15718 VDD.n719 VDD.n718 185
R15719 VDD.n2763 VDD.n2762 185
R15720 VDD.n2764 VDD.n2763 185
R15721 VDD.n2761 VDD.n728 185
R15722 VDD.n728 VDD.n725 185
R15723 VDD.n2760 VDD.n2759 185
R15724 VDD.n2759 VDD.n2758 185
R15725 VDD.n730 VDD.n729 185
R15726 VDD.n731 VDD.n730 185
R15727 VDD.n2751 VDD.n2750 185
R15728 VDD.n2752 VDD.n2751 185
R15729 VDD.n2749 VDD.n740 185
R15730 VDD.n740 VDD.n737 185
R15731 VDD.n2748 VDD.n2747 185
R15732 VDD.n2747 VDD.n2746 185
R15733 VDD.n742 VDD.n741 185
R15734 VDD.n743 VDD.n742 185
R15735 VDD.n2739 VDD.n2738 185
R15736 VDD.n2740 VDD.n2739 185
R15737 VDD.n2737 VDD.n752 185
R15738 VDD.n752 VDD.n749 185
R15739 VDD.n2736 VDD.n2735 185
R15740 VDD.n2735 VDD.n2734 185
R15741 VDD.n754 VDD.n753 185
R15742 VDD.n755 VDD.n754 185
R15743 VDD.n2727 VDD.n2726 185
R15744 VDD.n2728 VDD.n2727 185
R15745 VDD.n2725 VDD.n763 185
R15746 VDD.n769 VDD.n763 185
R15747 VDD.n2724 VDD.n2723 185
R15748 VDD.n2723 VDD.n2722 185
R15749 VDD.n765 VDD.n764 185
R15750 VDD.n766 VDD.n765 185
R15751 VDD.n2715 VDD.n2714 185
R15752 VDD.n2716 VDD.n2715 185
R15753 VDD.n2713 VDD.n776 185
R15754 VDD.n776 VDD.n773 185
R15755 VDD.n2712 VDD.n2711 185
R15756 VDD.n2711 VDD.n2710 185
R15757 VDD.n778 VDD.n777 185
R15758 VDD.n779 VDD.n778 185
R15759 VDD.n2703 VDD.n2702 185
R15760 VDD.n2704 VDD.n2703 185
R15761 VDD.n2701 VDD.n788 185
R15762 VDD.n788 VDD.n785 185
R15763 VDD.n2700 VDD.n2699 185
R15764 VDD.n2699 VDD.n2698 185
R15765 VDD.n790 VDD.n789 185
R15766 VDD.n791 VDD.n790 185
R15767 VDD.n2691 VDD.n2690 185
R15768 VDD.n2692 VDD.n2691 185
R15769 VDD.n2689 VDD.n800 185
R15770 VDD.n800 VDD.n797 185
R15771 VDD.n2688 VDD.n2687 185
R15772 VDD.n2687 VDD.n2686 185
R15773 VDD.n802 VDD.n801 185
R15774 VDD.n803 VDD.n802 185
R15775 VDD.n2679 VDD.n2678 185
R15776 VDD.n2680 VDD.n2679 185
R15777 VDD.n2677 VDD.n812 185
R15778 VDD.n812 VDD.n809 185
R15779 VDD.n2676 VDD.n2675 185
R15780 VDD.n2675 VDD.n2674 185
R15781 VDD.n814 VDD.n813 185
R15782 VDD.n815 VDD.n814 185
R15783 VDD.n2667 VDD.n2666 185
R15784 VDD.n2668 VDD.n2667 185
R15785 VDD.n2665 VDD.n824 185
R15786 VDD.n824 VDD.n821 185
R15787 VDD.n2664 VDD.n2663 185
R15788 VDD.n2663 VDD.n2662 185
R15789 VDD.n826 VDD.n825 185
R15790 VDD.n835 VDD.n826 185
R15791 VDD.n2655 VDD.n2654 185
R15792 VDD.n2656 VDD.n2655 185
R15793 VDD.n2653 VDD.n836 185
R15794 VDD.n836 VDD.n832 185
R15795 VDD.n2652 VDD.n2651 185
R15796 VDD.n2651 VDD.n2650 185
R15797 VDD.n838 VDD.n837 185
R15798 VDD.n839 VDD.n838 185
R15799 VDD.n2643 VDD.n2642 185
R15800 VDD.n2644 VDD.n2643 185
R15801 VDD.n2641 VDD.n848 185
R15802 VDD.n848 VDD.n845 185
R15803 VDD.n2640 VDD.n2639 185
R15804 VDD.n2639 VDD.n2638 185
R15805 VDD.n850 VDD.n849 185
R15806 VDD.n851 VDD.n850 185
R15807 VDD.n2631 VDD.n2630 185
R15808 VDD.n2632 VDD.n2631 185
R15809 VDD.n2629 VDD.n860 185
R15810 VDD.n860 VDD.n857 185
R15811 VDD.n2628 VDD.n2627 185
R15812 VDD.n2627 VDD.n2626 185
R15813 VDD.n862 VDD.n861 185
R15814 VDD.n863 VDD.n862 185
R15815 VDD.n2619 VDD.n2618 185
R15816 VDD.n2620 VDD.n2619 185
R15817 VDD.n2617 VDD.n872 185
R15818 VDD.n872 VDD.n869 185
R15819 VDD.n2616 VDD.n2615 185
R15820 VDD.n2615 VDD.n2614 185
R15821 VDD.n874 VDD.n873 185
R15822 VDD.t92 VDD.n874 185
R15823 VDD.n2607 VDD.n2606 185
R15824 VDD.n2608 VDD.n2607 185
R15825 VDD.n2605 VDD.n883 185
R15826 VDD.n883 VDD.n880 185
R15827 VDD.n2604 VDD.n2603 185
R15828 VDD.n2603 VDD.n2602 185
R15829 VDD.n885 VDD.n884 185
R15830 VDD.n886 VDD.n885 185
R15831 VDD.n2595 VDD.n2594 185
R15832 VDD.n2596 VDD.n2595 185
R15833 VDD.n2593 VDD.n895 185
R15834 VDD.n895 VDD.n892 185
R15835 VDD.n2592 VDD.n2591 185
R15836 VDD.n2591 VDD.n2590 185
R15837 VDD.n897 VDD.n896 185
R15838 VDD.n898 VDD.n897 185
R15839 VDD.n2583 VDD.n2582 185
R15840 VDD.n2584 VDD.n2583 185
R15841 VDD.n2581 VDD.n907 185
R15842 VDD.n907 VDD.n904 185
R15843 VDD.n2580 VDD.n2579 185
R15844 VDD.n2579 VDD.n2578 185
R15845 VDD.n909 VDD.n908 185
R15846 VDD.n910 VDD.n909 185
R15847 VDD.n2571 VDD.n2570 185
R15848 VDD.n2572 VDD.n2571 185
R15849 VDD.n2569 VDD.n919 185
R15850 VDD.n919 VDD.n916 185
R15851 VDD.n2568 VDD.n2567 185
R15852 VDD.n2567 VDD.n2566 185
R15853 VDD.n921 VDD.n920 185
R15854 VDD.n922 VDD.n921 185
R15855 VDD.n2559 VDD.n2558 185
R15856 VDD.n2560 VDD.n2559 185
R15857 VDD.n2557 VDD.n931 185
R15858 VDD.n931 VDD.n928 185
R15859 VDD.n2556 VDD.n2555 185
R15860 VDD.n2555 VDD.n2554 185
R15861 VDD.n933 VDD.n932 185
R15862 VDD.n934 VDD.n933 185
R15863 VDD.n2547 VDD.n2546 185
R15864 VDD.n2548 VDD.n2547 185
R15865 VDD.n2545 VDD.n942 185
R15866 VDD.n948 VDD.n942 185
R15867 VDD.n2544 VDD.n2543 185
R15868 VDD.n2543 VDD.n2542 185
R15869 VDD.n944 VDD.n943 185
R15870 VDD.n945 VDD.n944 185
R15871 VDD.n2535 VDD.n2534 185
R15872 VDD.n2536 VDD.n2535 185
R15873 VDD.n2533 VDD.n955 185
R15874 VDD.n955 VDD.n952 185
R15875 VDD.n2532 VDD.n2531 185
R15876 VDD.n2531 VDD.n2530 185
R15877 VDD.n957 VDD.n956 185
R15878 VDD.n958 VDD.n957 185
R15879 VDD.n2523 VDD.n2522 185
R15880 VDD.n2524 VDD.n2523 185
R15881 VDD.n2521 VDD.n967 185
R15882 VDD.n967 VDD.n964 185
R15883 VDD.n2520 VDD.n2519 185
R15884 VDD.n2519 VDD.n2518 185
R15885 VDD.n969 VDD.n968 185
R15886 VDD.n970 VDD.n969 185
R15887 VDD.n2511 VDD.n2510 185
R15888 VDD.n2512 VDD.n2511 185
R15889 VDD.n2509 VDD.n979 185
R15890 VDD.n979 VDD.n976 185
R15891 VDD.n2508 VDD.n2507 185
R15892 VDD.n2507 VDD.n2506 185
R15893 VDD.n981 VDD.n980 185
R15894 VDD.n982 VDD.n981 185
R15895 VDD.n2499 VDD.n2498 185
R15896 VDD.n2500 VDD.n2499 185
R15897 VDD.n2497 VDD.n991 185
R15898 VDD.n991 VDD.n988 185
R15899 VDD.n2496 VDD.n2495 185
R15900 VDD.n2495 VDD.n2494 185
R15901 VDD.n993 VDD.n992 185
R15902 VDD.n994 VDD.n993 185
R15903 VDD.n2487 VDD.n2486 185
R15904 VDD.n2488 VDD.n2487 185
R15905 VDD.n2485 VDD.n1003 185
R15906 VDD.n1003 VDD.n1000 185
R15907 VDD.n2484 VDD.n2483 185
R15908 VDD.n2483 VDD.n2482 185
R15909 VDD.n1005 VDD.n1004 185
R15910 VDD.n1006 VDD.n1005 185
R15911 VDD.n2475 VDD.n2474 185
R15912 VDD.n2476 VDD.n2475 185
R15913 VDD.n2473 VDD.n1015 185
R15914 VDD.n1015 VDD.n1012 185
R15915 VDD.n2472 VDD.n2471 185
R15916 VDD.n2471 VDD.n2470 185
R15917 VDD.n1017 VDD.n1016 185
R15918 VDD.n1026 VDD.n1017 185
R15919 VDD.n2463 VDD.n2462 185
R15920 VDD.n2464 VDD.n2463 185
R15921 VDD.n2461 VDD.n1027 185
R15922 VDD.n1027 VDD.n1023 185
R15923 VDD.n2460 VDD.n2459 185
R15924 VDD.n2459 VDD.n2458 185
R15925 VDD.n1029 VDD.n1028 185
R15926 VDD.n1030 VDD.n1029 185
R15927 VDD.n2451 VDD.n2450 185
R15928 VDD.n2452 VDD.n2451 185
R15929 VDD.n2449 VDD.n1039 185
R15930 VDD.n1039 VDD.n1036 185
R15931 VDD.n2448 VDD.n2447 185
R15932 VDD.n2447 VDD.n2446 185
R15933 VDD.n1041 VDD.n1040 185
R15934 VDD.n1042 VDD.n1041 185
R15935 VDD.n2439 VDD.n2438 185
R15936 VDD.n2440 VDD.n2439 185
R15937 VDD.n2437 VDD.n1051 185
R15938 VDD.n1051 VDD.n1048 185
R15939 VDD.n2436 VDD.n2435 185
R15940 VDD.n2435 VDD.n2434 185
R15941 VDD.n1053 VDD.n1052 185
R15942 VDD.n1054 VDD.n1053 185
R15943 VDD.n2427 VDD.n2426 185
R15944 VDD.n2428 VDD.n2427 185
R15945 VDD.n2425 VDD.n1063 185
R15946 VDD.n1063 VDD.n1060 185
R15947 VDD.n2424 VDD.n2423 185
R15948 VDD.n2423 VDD.n2422 185
R15949 VDD.n1065 VDD.n1064 185
R15950 VDD.n1074 VDD.n1065 185
R15951 VDD.n2415 VDD.n2414 185
R15952 VDD.n2416 VDD.n2415 185
R15953 VDD.n2413 VDD.n1075 185
R15954 VDD.n1075 VDD.n1071 185
R15955 VDD.n2412 VDD.n2411 185
R15956 VDD.n2411 VDD.n2410 185
R15957 VDD.n1077 VDD.n1076 185
R15958 VDD.n1078 VDD.n1077 185
R15959 VDD.n2403 VDD.n2402 185
R15960 VDD.n2404 VDD.n2403 185
R15961 VDD.n2401 VDD.n1087 185
R15962 VDD.n1087 VDD.n1084 185
R15963 VDD.n2400 VDD.n2399 185
R15964 VDD.n2399 VDD.n2398 185
R15965 VDD.n1089 VDD.n1088 185
R15966 VDD.n1090 VDD.n1089 185
R15967 VDD.n2391 VDD.n2390 185
R15968 VDD.n2392 VDD.n2391 185
R15969 VDD.n2389 VDD.n1099 185
R15970 VDD.n1099 VDD.n1096 185
R15971 VDD.n2388 VDD.n2387 185
R15972 VDD.n2387 VDD.n2386 185
R15973 VDD.n1101 VDD.n1100 185
R15974 VDD.n1902 VDD.n1901 185
R15975 VDD.n1903 VDD.n1899 185
R15976 VDD.n1899 VDD.n1102 185
R15977 VDD.n1905 VDD.n1904 185
R15978 VDD.n1907 VDD.n1898 185
R15979 VDD.n1910 VDD.n1909 185
R15980 VDD.n1911 VDD.n1897 185
R15981 VDD.n1913 VDD.n1912 185
R15982 VDD.n1915 VDD.n1896 185
R15983 VDD.n1918 VDD.n1917 185
R15984 VDD.n1919 VDD.n1137 185
R15985 VDD.n1921 VDD.n1920 185
R15986 VDD.n1923 VDD.n1136 185
R15987 VDD.n1926 VDD.n1925 185
R15988 VDD.n1928 VDD.n1133 185
R15989 VDD.n1930 VDD.n1929 185
R15990 VDD.n1932 VDD.n1132 185
R15991 VDD.n1934 VDD.n1933 185
R15992 VDD.n1933 VDD.n1102 185
R15993 VDD.n2825 VDD.n2824 185
R15994 VDD.n2827 VDD.n2826 185
R15995 VDD.n2829 VDD.n2828 185
R15996 VDD.n2831 VDD.n2830 185
R15997 VDD.n2833 VDD.n2832 185
R15998 VDD.n2835 VDD.n2834 185
R15999 VDD.n2837 VDD.n2836 185
R16000 VDD.n2839 VDD.n2838 185
R16001 VDD.n2841 VDD.n2840 185
R16002 VDD.n2843 VDD.n2842 185
R16003 VDD.n2845 VDD.n2844 185
R16004 VDD.n2847 VDD.n2846 185
R16005 VDD.n2849 VDD.n2848 185
R16006 VDD.n2851 VDD.n2850 185
R16007 VDD.n2853 VDD.n2852 185
R16008 VDD.n2855 VDD.n2854 185
R16009 VDD.n2857 VDD.n2856 185
R16010 VDD.n2859 VDD.n2858 185
R16011 VDD.n2823 VDD.n2822 185
R16012 VDD.n2823 VDD.n640 185
R16013 VDD.n2821 VDD.n667 185
R16014 VDD.n2863 VDD.n667 185
R16015 VDD.n2820 VDD.n2819 185
R16016 VDD.n2819 VDD.n666 185
R16017 VDD.n2818 VDD.n675 185
R16018 VDD.n2818 VDD.n2817 185
R16019 VDD.n2134 VDD.n676 185
R16020 VDD.n677 VDD.n676 185
R16021 VDD.n2135 VDD.n684 185
R16022 VDD.n2811 VDD.n684 185
R16023 VDD.n2137 VDD.n2136 185
R16024 VDD.n2136 VDD.n683 185
R16025 VDD.n2138 VDD.n691 185
R16026 VDD.n2800 VDD.n691 185
R16027 VDD.n2140 VDD.n2139 185
R16028 VDD.n2139 VDD.n690 185
R16029 VDD.n2141 VDD.n697 185
R16030 VDD.n2794 VDD.n697 185
R16031 VDD.n2143 VDD.n2142 185
R16032 VDD.n2142 VDD.n696 185
R16033 VDD.n2144 VDD.n702 185
R16034 VDD.n2788 VDD.n702 185
R16035 VDD.n2146 VDD.n2145 185
R16036 VDD.n2147 VDD.n2146 185
R16037 VDD.n2133 VDD.n708 185
R16038 VDD.n2782 VDD.n708 185
R16039 VDD.n2132 VDD.n2131 185
R16040 VDD.n2131 VDD.n707 185
R16041 VDD.n2130 VDD.n714 185
R16042 VDD.n2776 VDD.n714 185
R16043 VDD.n2129 VDD.n2128 185
R16044 VDD.n2128 VDD.n713 185
R16045 VDD.n2127 VDD.n720 185
R16046 VDD.n2770 VDD.n720 185
R16047 VDD.n2126 VDD.n2125 185
R16048 VDD.n2125 VDD.n719 185
R16049 VDD.n2124 VDD.n726 185
R16050 VDD.n2764 VDD.n726 185
R16051 VDD.n2123 VDD.n2122 185
R16052 VDD.n2122 VDD.n725 185
R16053 VDD.n2121 VDD.n732 185
R16054 VDD.n2758 VDD.n732 185
R16055 VDD.n2120 VDD.n2119 185
R16056 VDD.n2119 VDD.n731 185
R16057 VDD.n2118 VDD.n738 185
R16058 VDD.n2752 VDD.n738 185
R16059 VDD.n2117 VDD.n2116 185
R16060 VDD.n2116 VDD.n737 185
R16061 VDD.n2115 VDD.n744 185
R16062 VDD.n2746 VDD.n744 185
R16063 VDD.n2114 VDD.n2113 185
R16064 VDD.n2113 VDD.n743 185
R16065 VDD.n2112 VDD.n750 185
R16066 VDD.n2740 VDD.n750 185
R16067 VDD.n2111 VDD.n2110 185
R16068 VDD.n2110 VDD.n749 185
R16069 VDD.n2109 VDD.n756 185
R16070 VDD.n2734 VDD.n756 185
R16071 VDD.n2108 VDD.n2107 185
R16072 VDD.n2107 VDD.n755 185
R16073 VDD.n2106 VDD.n761 185
R16074 VDD.n2728 VDD.n761 185
R16075 VDD.n2105 VDD.n2104 185
R16076 VDD.n2104 VDD.n769 185
R16077 VDD.n2103 VDD.n767 185
R16078 VDD.n2722 VDD.n767 185
R16079 VDD.n2102 VDD.n2101 185
R16080 VDD.n2101 VDD.n766 185
R16081 VDD.n2100 VDD.n774 185
R16082 VDD.n2716 VDD.n774 185
R16083 VDD.n2099 VDD.n2098 185
R16084 VDD.n2098 VDD.n773 185
R16085 VDD.n2097 VDD.n780 185
R16086 VDD.n2710 VDD.n780 185
R16087 VDD.n2096 VDD.n2095 185
R16088 VDD.n2095 VDD.n779 185
R16089 VDD.n2094 VDD.n786 185
R16090 VDD.n2704 VDD.n786 185
R16091 VDD.n2093 VDD.n2092 185
R16092 VDD.n2092 VDD.n785 185
R16093 VDD.n2091 VDD.n792 185
R16094 VDD.n2698 VDD.n792 185
R16095 VDD.n2090 VDD.n2089 185
R16096 VDD.n2089 VDD.n791 185
R16097 VDD.n2088 VDD.n798 185
R16098 VDD.n2692 VDD.n798 185
R16099 VDD.n2087 VDD.n2086 185
R16100 VDD.n2086 VDD.n797 185
R16101 VDD.n2085 VDD.n804 185
R16102 VDD.n2686 VDD.n804 185
R16103 VDD.n2084 VDD.n2083 185
R16104 VDD.n2083 VDD.n803 185
R16105 VDD.n2082 VDD.n810 185
R16106 VDD.n2680 VDD.n810 185
R16107 VDD.n2081 VDD.n2080 185
R16108 VDD.n2080 VDD.n809 185
R16109 VDD.n2079 VDD.n816 185
R16110 VDD.n2674 VDD.n816 185
R16111 VDD.n2078 VDD.n2077 185
R16112 VDD.n2077 VDD.n815 185
R16113 VDD.n2076 VDD.n822 185
R16114 VDD.n2668 VDD.n822 185
R16115 VDD.n2075 VDD.n2074 185
R16116 VDD.n2074 VDD.n821 185
R16117 VDD.n2073 VDD.n827 185
R16118 VDD.n2662 VDD.n827 185
R16119 VDD.n2072 VDD.n2071 185
R16120 VDD.n2071 VDD.n835 185
R16121 VDD.n2070 VDD.n833 185
R16122 VDD.n2656 VDD.n833 185
R16123 VDD.n2069 VDD.n2068 185
R16124 VDD.n2068 VDD.n832 185
R16125 VDD.n2067 VDD.n840 185
R16126 VDD.n2650 VDD.n840 185
R16127 VDD.n2066 VDD.n2065 185
R16128 VDD.n2065 VDD.n839 185
R16129 VDD.n2064 VDD.n846 185
R16130 VDD.n2644 VDD.n846 185
R16131 VDD.n2063 VDD.n2062 185
R16132 VDD.n2062 VDD.n845 185
R16133 VDD.n2061 VDD.n852 185
R16134 VDD.n2638 VDD.n852 185
R16135 VDD.n2060 VDD.n2059 185
R16136 VDD.n2059 VDD.n851 185
R16137 VDD.n2058 VDD.n858 185
R16138 VDD.n2632 VDD.n858 185
R16139 VDD.n2057 VDD.n2056 185
R16140 VDD.n2056 VDD.n857 185
R16141 VDD.n2055 VDD.n864 185
R16142 VDD.n2626 VDD.n864 185
R16143 VDD.n2054 VDD.n2053 185
R16144 VDD.n2053 VDD.n863 185
R16145 VDD.n2052 VDD.n870 185
R16146 VDD.n2620 VDD.n870 185
R16147 VDD.n2051 VDD.n2050 185
R16148 VDD.n2050 VDD.n869 185
R16149 VDD.n2049 VDD.n875 185
R16150 VDD.n2614 VDD.n875 185
R16151 VDD.n2048 VDD.n2047 185
R16152 VDD.n2047 VDD.t92 185
R16153 VDD.n2046 VDD.n881 185
R16154 VDD.n2608 VDD.n881 185
R16155 VDD.n2045 VDD.n2044 185
R16156 VDD.n2044 VDD.n880 185
R16157 VDD.n2043 VDD.n887 185
R16158 VDD.n2602 VDD.n887 185
R16159 VDD.n2042 VDD.n2041 185
R16160 VDD.n2041 VDD.n886 185
R16161 VDD.n2040 VDD.n893 185
R16162 VDD.n2596 VDD.n893 185
R16163 VDD.n2039 VDD.n2038 185
R16164 VDD.n2038 VDD.n892 185
R16165 VDD.n2037 VDD.n899 185
R16166 VDD.n2590 VDD.n899 185
R16167 VDD.n2036 VDD.n2035 185
R16168 VDD.n2035 VDD.n898 185
R16169 VDD.n2034 VDD.n905 185
R16170 VDD.n2584 VDD.n905 185
R16171 VDD.n2033 VDD.n2032 185
R16172 VDD.n2032 VDD.n904 185
R16173 VDD.n2031 VDD.n911 185
R16174 VDD.n2578 VDD.n911 185
R16175 VDD.n2030 VDD.n2029 185
R16176 VDD.n2029 VDD.n910 185
R16177 VDD.n2028 VDD.n917 185
R16178 VDD.n2572 VDD.n917 185
R16179 VDD.n2027 VDD.n2026 185
R16180 VDD.n2026 VDD.n916 185
R16181 VDD.n2025 VDD.n923 185
R16182 VDD.n2566 VDD.n923 185
R16183 VDD.n2024 VDD.n2023 185
R16184 VDD.n2023 VDD.n922 185
R16185 VDD.n2022 VDD.n929 185
R16186 VDD.n2560 VDD.n929 185
R16187 VDD.n2021 VDD.n2020 185
R16188 VDD.n2020 VDD.n928 185
R16189 VDD.n2019 VDD.n935 185
R16190 VDD.n2554 VDD.n935 185
R16191 VDD.n2018 VDD.n2017 185
R16192 VDD.n2017 VDD.n934 185
R16193 VDD.n2016 VDD.n940 185
R16194 VDD.n2548 VDD.n940 185
R16195 VDD.n2015 VDD.n2014 185
R16196 VDD.n2014 VDD.n948 185
R16197 VDD.n2013 VDD.n946 185
R16198 VDD.n2542 VDD.n946 185
R16199 VDD.n2012 VDD.n2011 185
R16200 VDD.n2011 VDD.n945 185
R16201 VDD.n2010 VDD.n953 185
R16202 VDD.n2536 VDD.n953 185
R16203 VDD.n2009 VDD.n2008 185
R16204 VDD.n2008 VDD.n952 185
R16205 VDD.n2007 VDD.n959 185
R16206 VDD.n2530 VDD.n959 185
R16207 VDD.n2006 VDD.n2005 185
R16208 VDD.n2005 VDD.n958 185
R16209 VDD.n2004 VDD.n965 185
R16210 VDD.n2524 VDD.n965 185
R16211 VDD.n2003 VDD.n2002 185
R16212 VDD.n2002 VDD.n964 185
R16213 VDD.n2001 VDD.n971 185
R16214 VDD.n2518 VDD.n971 185
R16215 VDD.n2000 VDD.n1999 185
R16216 VDD.n1999 VDD.n970 185
R16217 VDD.n1998 VDD.n977 185
R16218 VDD.n2512 VDD.n977 185
R16219 VDD.n1997 VDD.n1996 185
R16220 VDD.n1996 VDD.n976 185
R16221 VDD.n1995 VDD.n983 185
R16222 VDD.n2506 VDD.n983 185
R16223 VDD.n1994 VDD.n1993 185
R16224 VDD.n1993 VDD.n982 185
R16225 VDD.n1992 VDD.n989 185
R16226 VDD.n2500 VDD.n989 185
R16227 VDD.n1991 VDD.n1990 185
R16228 VDD.n1990 VDD.n988 185
R16229 VDD.n1989 VDD.n995 185
R16230 VDD.n2494 VDD.n995 185
R16231 VDD.n1988 VDD.n1987 185
R16232 VDD.n1987 VDD.n994 185
R16233 VDD.n1986 VDD.n1001 185
R16234 VDD.n2488 VDD.n1001 185
R16235 VDD.n1985 VDD.n1984 185
R16236 VDD.n1984 VDD.n1000 185
R16237 VDD.n1983 VDD.n1007 185
R16238 VDD.n2482 VDD.n1007 185
R16239 VDD.n1982 VDD.n1981 185
R16240 VDD.n1981 VDD.n1006 185
R16241 VDD.n1980 VDD.n1013 185
R16242 VDD.n2476 VDD.n1013 185
R16243 VDD.n1979 VDD.n1978 185
R16244 VDD.n1978 VDD.n1012 185
R16245 VDD.n1977 VDD.n1018 185
R16246 VDD.n2470 VDD.n1018 185
R16247 VDD.n1976 VDD.n1975 185
R16248 VDD.n1975 VDD.n1026 185
R16249 VDD.n1974 VDD.n1024 185
R16250 VDD.n2464 VDD.n1024 185
R16251 VDD.n1973 VDD.n1972 185
R16252 VDD.n1972 VDD.n1023 185
R16253 VDD.n1971 VDD.n1031 185
R16254 VDD.n2458 VDD.n1031 185
R16255 VDD.n1970 VDD.n1969 185
R16256 VDD.n1969 VDD.n1030 185
R16257 VDD.n1968 VDD.n1037 185
R16258 VDD.n2452 VDD.n1037 185
R16259 VDD.n1967 VDD.n1966 185
R16260 VDD.n1966 VDD.n1036 185
R16261 VDD.n1965 VDD.n1043 185
R16262 VDD.n2446 VDD.n1043 185
R16263 VDD.n1964 VDD.n1963 185
R16264 VDD.n1963 VDD.n1042 185
R16265 VDD.n1962 VDD.n1049 185
R16266 VDD.n2440 VDD.n1049 185
R16267 VDD.n1961 VDD.n1960 185
R16268 VDD.n1960 VDD.n1048 185
R16269 VDD.n1959 VDD.n1055 185
R16270 VDD.n2434 VDD.n1055 185
R16271 VDD.n1958 VDD.n1957 185
R16272 VDD.n1957 VDD.n1054 185
R16273 VDD.n1956 VDD.n1061 185
R16274 VDD.n2428 VDD.n1061 185
R16275 VDD.n1955 VDD.n1954 185
R16276 VDD.n1954 VDD.n1060 185
R16277 VDD.n1953 VDD.n1066 185
R16278 VDD.n2422 VDD.n1066 185
R16279 VDD.n1952 VDD.n1951 185
R16280 VDD.n1951 VDD.n1074 185
R16281 VDD.n1950 VDD.n1072 185
R16282 VDD.n2416 VDD.n1072 185
R16283 VDD.n1949 VDD.n1948 185
R16284 VDD.n1948 VDD.n1071 185
R16285 VDD.n1947 VDD.n1079 185
R16286 VDD.n2410 VDD.n1079 185
R16287 VDD.n1946 VDD.n1945 185
R16288 VDD.n1945 VDD.n1078 185
R16289 VDD.n1944 VDD.n1085 185
R16290 VDD.n2404 VDD.n1085 185
R16291 VDD.n1943 VDD.n1942 185
R16292 VDD.n1942 VDD.n1084 185
R16293 VDD.n1941 VDD.n1091 185
R16294 VDD.n2398 VDD.n1091 185
R16295 VDD.n1940 VDD.n1939 185
R16296 VDD.n1939 VDD.n1090 185
R16297 VDD.n1938 VDD.n1097 185
R16298 VDD.n2392 VDD.n1097 185
R16299 VDD.n1937 VDD.n1936 185
R16300 VDD.n1936 VDD.n1096 185
R16301 VDD.n1935 VDD.n1103 185
R16302 VDD.n2386 VDD.n1103 185
R16303 VDD.n3924 VDD.n3923 185
R16304 VDD.n3925 VDD.n3924 185
R16305 VDD.n191 VDD.n189 185
R16306 VDD.n189 VDD.n186 185
R16307 VDD.n3883 VDD.n3882 185
R16308 VDD.n3884 VDD.n3883 185
R16309 VDD.n3881 VDD.n212 185
R16310 VDD.n212 VDD.n209 185
R16311 VDD.n3880 VDD.n3879 185
R16312 VDD.n3879 VDD.n3878 185
R16313 VDD.n214 VDD.n213 185
R16314 VDD.n215 VDD.n214 185
R16315 VDD.n3845 VDD.n3844 185
R16316 VDD.n3846 VDD.n3845 185
R16317 VDD.n3843 VDD.n225 185
R16318 VDD.n225 VDD.n222 185
R16319 VDD.n3842 VDD.n3841 185
R16320 VDD.n3841 VDD.n3840 185
R16321 VDD.n227 VDD.n226 185
R16322 VDD.n236 VDD.n227 185
R16323 VDD.n3833 VDD.n3832 185
R16324 VDD.n3834 VDD.n3833 185
R16325 VDD.n3831 VDD.n237 185
R16326 VDD.n237 VDD.n233 185
R16327 VDD.n3830 VDD.n3829 185
R16328 VDD.n3829 VDD.n3828 185
R16329 VDD.n239 VDD.n238 185
R16330 VDD.n240 VDD.n239 185
R16331 VDD.n3821 VDD.n3820 185
R16332 VDD.n3822 VDD.n3821 185
R16333 VDD.n3819 VDD.n249 185
R16334 VDD.n249 VDD.n246 185
R16335 VDD.n3818 VDD.n3817 185
R16336 VDD.n3817 VDD.n3816 185
R16337 VDD.n251 VDD.n250 185
R16338 VDD.n252 VDD.n251 185
R16339 VDD.n3809 VDD.n3808 185
R16340 VDD.n3810 VDD.n3809 185
R16341 VDD.n3807 VDD.n261 185
R16342 VDD.n261 VDD.n258 185
R16343 VDD.n3806 VDD.n3805 185
R16344 VDD.n3805 VDD.n3804 185
R16345 VDD.n263 VDD.n262 185
R16346 VDD.n264 VDD.n263 185
R16347 VDD.n3797 VDD.n3796 185
R16348 VDD.n3798 VDD.n3797 185
R16349 VDD.n3795 VDD.n273 185
R16350 VDD.n273 VDD.n270 185
R16351 VDD.n3794 VDD.n3793 185
R16352 VDD.n3793 VDD.n3792 185
R16353 VDD.n275 VDD.n274 185
R16354 VDD.n276 VDD.n275 185
R16355 VDD.n3785 VDD.n3784 185
R16356 VDD.n3786 VDD.n3785 185
R16357 VDD.n3783 VDD.n285 185
R16358 VDD.n285 VDD.n282 185
R16359 VDD.n3782 VDD.n3781 185
R16360 VDD.n3781 VDD.n3780 185
R16361 VDD.n287 VDD.n286 185
R16362 VDD.n288 VDD.n287 185
R16363 VDD.n3773 VDD.n3772 185
R16364 VDD.n3774 VDD.n3773 185
R16365 VDD.n3771 VDD.n297 185
R16366 VDD.n297 VDD.n294 185
R16367 VDD.n3770 VDD.n3769 185
R16368 VDD.n3769 VDD.n3768 185
R16369 VDD.n299 VDD.n298 185
R16370 VDD.n300 VDD.n299 185
R16371 VDD.n3761 VDD.n3760 185
R16372 VDD.n3762 VDD.n3761 185
R16373 VDD.n3759 VDD.n308 185
R16374 VDD.n314 VDD.n308 185
R16375 VDD.n3758 VDD.n3757 185
R16376 VDD.n3757 VDD.n3756 185
R16377 VDD.n310 VDD.n309 185
R16378 VDD.n311 VDD.n310 185
R16379 VDD.n3749 VDD.n3748 185
R16380 VDD.n3750 VDD.n3749 185
R16381 VDD.n3747 VDD.n321 185
R16382 VDD.n321 VDD.n318 185
R16383 VDD.n3746 VDD.n3745 185
R16384 VDD.n3745 VDD.n3744 185
R16385 VDD.n323 VDD.n322 185
R16386 VDD.n324 VDD.n323 185
R16387 VDD.n3737 VDD.n3736 185
R16388 VDD.n3738 VDD.n3737 185
R16389 VDD.n3735 VDD.n333 185
R16390 VDD.n333 VDD.n330 185
R16391 VDD.n3734 VDD.n3733 185
R16392 VDD.n3733 VDD.n3732 185
R16393 VDD.n335 VDD.n334 185
R16394 VDD.n336 VDD.n335 185
R16395 VDD.n3725 VDD.n3724 185
R16396 VDD.n3726 VDD.n3725 185
R16397 VDD.n3723 VDD.n344 185
R16398 VDD.n350 VDD.n344 185
R16399 VDD.n3722 VDD.n3721 185
R16400 VDD.n3721 VDD.n3720 185
R16401 VDD.n346 VDD.n345 185
R16402 VDD.n347 VDD.n346 185
R16403 VDD.n3713 VDD.n3712 185
R16404 VDD.n3714 VDD.n3713 185
R16405 VDD.n3711 VDD.n357 185
R16406 VDD.n357 VDD.n354 185
R16407 VDD.n3710 VDD.n3709 185
R16408 VDD.n3709 VDD.n3708 185
R16409 VDD.n359 VDD.n358 185
R16410 VDD.n360 VDD.n359 185
R16411 VDD.n3701 VDD.n3700 185
R16412 VDD.n3702 VDD.n3701 185
R16413 VDD.n3699 VDD.n369 185
R16414 VDD.n369 VDD.n366 185
R16415 VDD.n3698 VDD.n3697 185
R16416 VDD.n3697 VDD.n3696 185
R16417 VDD.n371 VDD.n370 185
R16418 VDD.n372 VDD.n371 185
R16419 VDD.n3689 VDD.n3688 185
R16420 VDD.n3690 VDD.n3689 185
R16421 VDD.n3687 VDD.n381 185
R16422 VDD.n381 VDD.n378 185
R16423 VDD.n3686 VDD.n3685 185
R16424 VDD.n3685 VDD.n3684 185
R16425 VDD.n383 VDD.n382 185
R16426 VDD.n384 VDD.n383 185
R16427 VDD.n3677 VDD.n3676 185
R16428 VDD.n3678 VDD.n3677 185
R16429 VDD.n3675 VDD.n393 185
R16430 VDD.n393 VDD.n390 185
R16431 VDD.n3674 VDD.n3673 185
R16432 VDD.n3673 VDD.n3672 185
R16433 VDD.n395 VDD.n394 185
R16434 VDD.n396 VDD.n395 185
R16435 VDD.n3665 VDD.n3664 185
R16436 VDD.n3666 VDD.n3665 185
R16437 VDD.n3663 VDD.n405 185
R16438 VDD.n405 VDD.n402 185
R16439 VDD.n3662 VDD.n3661 185
R16440 VDD.n3661 VDD.n3660 185
R16441 VDD.n407 VDD.n406 185
R16442 VDD.n408 VDD.n407 185
R16443 VDD.n3653 VDD.n3652 185
R16444 VDD.n3654 VDD.n3653 185
R16445 VDD.n3651 VDD.n417 185
R16446 VDD.n417 VDD.n414 185
R16447 VDD.n3650 VDD.n3649 185
R16448 VDD.n3649 VDD.n3648 185
R16449 VDD.n419 VDD.n418 185
R16450 VDD.n427 VDD.n419 185
R16451 VDD.n3641 VDD.n3640 185
R16452 VDD.n3642 VDD.n3641 185
R16453 VDD.n3639 VDD.n428 185
R16454 VDD.n428 VDD.t132 185
R16455 VDD.n3638 VDD.n3637 185
R16456 VDD.n3637 VDD.n3636 185
R16457 VDD.n430 VDD.n429 185
R16458 VDD.n431 VDD.n430 185
R16459 VDD.n3629 VDD.n3628 185
R16460 VDD.n3630 VDD.n3629 185
R16461 VDD.n3627 VDD.n440 185
R16462 VDD.n440 VDD.n437 185
R16463 VDD.n3626 VDD.n3625 185
R16464 VDD.n3625 VDD.n3624 185
R16465 VDD.n442 VDD.n441 185
R16466 VDD.n443 VDD.n442 185
R16467 VDD.n3617 VDD.n3616 185
R16468 VDD.n3618 VDD.n3617 185
R16469 VDD.n3615 VDD.n452 185
R16470 VDD.n452 VDD.n449 185
R16471 VDD.n3614 VDD.n3613 185
R16472 VDD.n3613 VDD.n3612 185
R16473 VDD.n454 VDD.n453 185
R16474 VDD.n455 VDD.n454 185
R16475 VDD.n3605 VDD.n3604 185
R16476 VDD.n3606 VDD.n3605 185
R16477 VDD.n3603 VDD.n464 185
R16478 VDD.n464 VDD.n461 185
R16479 VDD.n3602 VDD.n3601 185
R16480 VDD.n3601 VDD.n3600 185
R16481 VDD.n466 VDD.n465 185
R16482 VDD.n467 VDD.n466 185
R16483 VDD.n3593 VDD.n3592 185
R16484 VDD.n3594 VDD.n3593 185
R16485 VDD.n3591 VDD.n476 185
R16486 VDD.n476 VDD.n473 185
R16487 VDD.n3590 VDD.n3589 185
R16488 VDD.n3589 VDD.n3588 185
R16489 VDD.n478 VDD.n477 185
R16490 VDD.n479 VDD.n478 185
R16491 VDD.n3581 VDD.n3580 185
R16492 VDD.n3582 VDD.n3581 185
R16493 VDD.n3579 VDD.n487 185
R16494 VDD.n493 VDD.n487 185
R16495 VDD.n3578 VDD.n3577 185
R16496 VDD.n3577 VDD.n3576 185
R16497 VDD.n489 VDD.n488 185
R16498 VDD.n490 VDD.n489 185
R16499 VDD.n3569 VDD.n3568 185
R16500 VDD.n3570 VDD.n3569 185
R16501 VDD.n3567 VDD.n500 185
R16502 VDD.n500 VDD.n497 185
R16503 VDD.n3566 VDD.n3565 185
R16504 VDD.n3565 VDD.n3564 185
R16505 VDD.n502 VDD.n501 185
R16506 VDD.n503 VDD.n502 185
R16507 VDD.n3557 VDD.n3556 185
R16508 VDD.n3558 VDD.n3557 185
R16509 VDD.n3555 VDD.n512 185
R16510 VDD.n512 VDD.n509 185
R16511 VDD.n3554 VDD.n3553 185
R16512 VDD.n3553 VDD.n3552 185
R16513 VDD.n514 VDD.n513 185
R16514 VDD.n515 VDD.n514 185
R16515 VDD.n3545 VDD.n3544 185
R16516 VDD.n3546 VDD.n3545 185
R16517 VDD.n3543 VDD.n524 185
R16518 VDD.n524 VDD.n521 185
R16519 VDD.n3542 VDD.n3541 185
R16520 VDD.n3541 VDD.n3540 185
R16521 VDD.n526 VDD.n525 185
R16522 VDD.n527 VDD.n526 185
R16523 VDD.n3533 VDD.n3532 185
R16524 VDD.n3534 VDD.n3533 185
R16525 VDD.n3531 VDD.n535 185
R16526 VDD.n541 VDD.n535 185
R16527 VDD.n3530 VDD.n3529 185
R16528 VDD.n3529 VDD.n3528 185
R16529 VDD.n537 VDD.n536 185
R16530 VDD.n538 VDD.n537 185
R16531 VDD.n3521 VDD.n3520 185
R16532 VDD.n3522 VDD.n3521 185
R16533 VDD.n3519 VDD.n548 185
R16534 VDD.n548 VDD.n545 185
R16535 VDD.n3518 VDD.n3517 185
R16536 VDD.n3517 VDD.n3516 185
R16537 VDD.n550 VDD.n549 185
R16538 VDD.n551 VDD.n550 185
R16539 VDD.n3509 VDD.n3508 185
R16540 VDD.n3510 VDD.n3509 185
R16541 VDD.n3507 VDD.n560 185
R16542 VDD.n560 VDD.n557 185
R16543 VDD.n3506 VDD.n3505 185
R16544 VDD.n3505 VDD.n3504 185
R16545 VDD.n562 VDD.n561 185
R16546 VDD.n563 VDD.n562 185
R16547 VDD.n3497 VDD.n3496 185
R16548 VDD.n3498 VDD.n3497 185
R16549 VDD.n3495 VDD.n572 185
R16550 VDD.n572 VDD.n569 185
R16551 VDD.n3494 VDD.n3493 185
R16552 VDD.n3493 VDD.n3492 185
R16553 VDD.n574 VDD.n573 185
R16554 VDD.n575 VDD.n574 185
R16555 VDD.n3485 VDD.n3484 185
R16556 VDD.n3486 VDD.n3485 185
R16557 VDD.n3483 VDD.n584 185
R16558 VDD.n584 VDD.n581 185
R16559 VDD.n3482 VDD.n3481 185
R16560 VDD.n3481 VDD.n3480 185
R16561 VDD.n586 VDD.n585 185
R16562 VDD.n587 VDD.n586 185
R16563 VDD.n3473 VDD.n3472 185
R16564 VDD.n3474 VDD.n3473 185
R16565 VDD.n3471 VDD.n596 185
R16566 VDD.n596 VDD.n593 185
R16567 VDD.n3470 VDD.n3469 185
R16568 VDD.n3469 VDD.n3468 185
R16569 VDD.n598 VDD.n597 185
R16570 VDD.n3369 VDD.n598 185
R16571 VDD.n3461 VDD.n3460 185
R16572 VDD.n3462 VDD.n3461 185
R16573 VDD.n3459 VDD.n607 185
R16574 VDD.n607 VDD.n604 185
R16575 VDD.n3458 VDD.n3457 185
R16576 VDD.n3457 VDD.n3456 185
R16577 VDD.n609 VDD.n608 185
R16578 VDD.n610 VDD.n609 185
R16579 VDD.n3449 VDD.n3448 185
R16580 VDD.n3450 VDD.n3449 185
R16581 VDD.n3447 VDD.n619 185
R16582 VDD.n619 VDD.n616 185
R16583 VDD.n3446 VDD.n3445 185
R16584 VDD.n3445 VDD.n3444 185
R16585 VDD.n621 VDD.n620 185
R16586 VDD.n622 VDD.n621 185
R16587 VDD.n3437 VDD.n3436 185
R16588 VDD.n3438 VDD.n3437 185
R16589 VDD.n3435 VDD.n631 185
R16590 VDD.n631 VDD.n628 185
R16591 VDD.n3434 VDD.n3433 185
R16592 VDD.n3433 VDD.n3432 185
R16593 VDD.n633 VDD.n632 185
R16594 VDD.n634 VDD.n633 185
R16595 VDD.n3423 VDD.n3422 185
R16596 VDD.n3421 VDD.n2920 185
R16597 VDD.n3420 VDD.n2919 185
R16598 VDD.n3425 VDD.n2919 185
R16599 VDD.n3419 VDD.n3418 185
R16600 VDD.n3417 VDD.n3416 185
R16601 VDD.n3415 VDD.n3414 185
R16602 VDD.n3413 VDD.n3412 185
R16603 VDD.n3411 VDD.n3410 185
R16604 VDD.n3409 VDD.n3408 185
R16605 VDD.n3407 VDD.n3406 185
R16606 VDD.n3405 VDD.n3404 185
R16607 VDD.n3403 VDD.n3402 185
R16608 VDD.n3401 VDD.n3400 185
R16609 VDD.n3399 VDD.n3398 185
R16610 VDD.n3396 VDD.n3395 185
R16611 VDD.n3394 VDD.n3393 185
R16612 VDD.n3392 VDD.n3391 185
R16613 VDD.n3390 VDD.n2910 185
R16614 VDD.n3425 VDD.n2910 185
R16615 VDD.n3891 VDD.n3890 185
R16616 VDD.n3892 VDD.n206 185
R16617 VDD.n3894 VDD.n3893 185
R16618 VDD.n3896 VDD.n205 185
R16619 VDD.n3898 VDD.n3897 185
R16620 VDD.n3899 VDD.n200 185
R16621 VDD.n3901 VDD.n3900 185
R16622 VDD.n3903 VDD.n198 185
R16623 VDD.n3905 VDD.n3904 185
R16624 VDD.n3908 VDD.n197 185
R16625 VDD.n3910 VDD.n3909 185
R16626 VDD.n3912 VDD.n195 185
R16627 VDD.n3914 VDD.n3913 185
R16628 VDD.n3915 VDD.n194 185
R16629 VDD.n3917 VDD.n3916 185
R16630 VDD.n3919 VDD.n192 185
R16631 VDD.n3921 VDD.n3920 185
R16632 VDD.n3922 VDD.n190 185
R16633 VDD.n3888 VDD.n187 185
R16634 VDD.n3925 VDD.n187 185
R16635 VDD.n3887 VDD.n3886 185
R16636 VDD.n3886 VDD.n186 185
R16637 VDD.n3885 VDD.n207 185
R16638 VDD.n3885 VDD.n3884 185
R16639 VDD.n2923 VDD.n208 185
R16640 VDD.n209 VDD.n208 185
R16641 VDD.n2924 VDD.n216 185
R16642 VDD.n3878 VDD.n216 185
R16643 VDD.n2926 VDD.n2925 185
R16644 VDD.n2925 VDD.n215 185
R16645 VDD.n2927 VDD.n223 185
R16646 VDD.n3846 VDD.n223 185
R16647 VDD.n2929 VDD.n2928 185
R16648 VDD.n2928 VDD.n222 185
R16649 VDD.n2930 VDD.n228 185
R16650 VDD.n3840 VDD.n228 185
R16651 VDD.n2932 VDD.n2931 185
R16652 VDD.n2931 VDD.n236 185
R16653 VDD.n2933 VDD.n234 185
R16654 VDD.n3834 VDD.n234 185
R16655 VDD.n2935 VDD.n2934 185
R16656 VDD.n2934 VDD.n233 185
R16657 VDD.n2936 VDD.n241 185
R16658 VDD.n3828 VDD.n241 185
R16659 VDD.n2938 VDD.n2937 185
R16660 VDD.n2937 VDD.n240 185
R16661 VDD.n2939 VDD.n247 185
R16662 VDD.n3822 VDD.n247 185
R16663 VDD.n2941 VDD.n2940 185
R16664 VDD.n2940 VDD.n246 185
R16665 VDD.n2942 VDD.n253 185
R16666 VDD.n3816 VDD.n253 185
R16667 VDD.n2944 VDD.n2943 185
R16668 VDD.n2943 VDD.n252 185
R16669 VDD.n2945 VDD.n259 185
R16670 VDD.n3810 VDD.n259 185
R16671 VDD.n2947 VDD.n2946 185
R16672 VDD.n2946 VDD.n258 185
R16673 VDD.n2948 VDD.n265 185
R16674 VDD.n3804 VDD.n265 185
R16675 VDD.n2950 VDD.n2949 185
R16676 VDD.n2949 VDD.n264 185
R16677 VDD.n2951 VDD.n271 185
R16678 VDD.n3798 VDD.n271 185
R16679 VDD.n2953 VDD.n2952 185
R16680 VDD.n2952 VDD.n270 185
R16681 VDD.n2954 VDD.n277 185
R16682 VDD.n3792 VDD.n277 185
R16683 VDD.n2956 VDD.n2955 185
R16684 VDD.n2955 VDD.n276 185
R16685 VDD.n2957 VDD.n283 185
R16686 VDD.n3786 VDD.n283 185
R16687 VDD.n2959 VDD.n2958 185
R16688 VDD.n2958 VDD.n282 185
R16689 VDD.n2960 VDD.n289 185
R16690 VDD.n3780 VDD.n289 185
R16691 VDD.n2962 VDD.n2961 185
R16692 VDD.n2961 VDD.n288 185
R16693 VDD.n2963 VDD.n295 185
R16694 VDD.n3774 VDD.n295 185
R16695 VDD.n2965 VDD.n2964 185
R16696 VDD.n2964 VDD.n294 185
R16697 VDD.n2966 VDD.n301 185
R16698 VDD.n3768 VDD.n301 185
R16699 VDD.n2968 VDD.n2967 185
R16700 VDD.n2967 VDD.n300 185
R16701 VDD.n2969 VDD.n306 185
R16702 VDD.n3762 VDD.n306 185
R16703 VDD.n2971 VDD.n2970 185
R16704 VDD.n2970 VDD.n314 185
R16705 VDD.n2972 VDD.n312 185
R16706 VDD.n3756 VDD.n312 185
R16707 VDD.n2974 VDD.n2973 185
R16708 VDD.n2973 VDD.n311 185
R16709 VDD.n2975 VDD.n319 185
R16710 VDD.n3750 VDD.n319 185
R16711 VDD.n2977 VDD.n2976 185
R16712 VDD.n2976 VDD.n318 185
R16713 VDD.n2978 VDD.n325 185
R16714 VDD.n3744 VDD.n325 185
R16715 VDD.n2980 VDD.n2979 185
R16716 VDD.n2979 VDD.n324 185
R16717 VDD.n2981 VDD.n331 185
R16718 VDD.n3738 VDD.n331 185
R16719 VDD.n2983 VDD.n2982 185
R16720 VDD.n2982 VDD.n330 185
R16721 VDD.n2984 VDD.n337 185
R16722 VDD.n3732 VDD.n337 185
R16723 VDD.n2986 VDD.n2985 185
R16724 VDD.n2985 VDD.n336 185
R16725 VDD.n2987 VDD.n342 185
R16726 VDD.n3726 VDD.n342 185
R16727 VDD.n2989 VDD.n2988 185
R16728 VDD.n2988 VDD.n350 185
R16729 VDD.n2990 VDD.n348 185
R16730 VDD.n3720 VDD.n348 185
R16731 VDD.n2992 VDD.n2991 185
R16732 VDD.n2991 VDD.n347 185
R16733 VDD.n2993 VDD.n355 185
R16734 VDD.n3714 VDD.n355 185
R16735 VDD.n2995 VDD.n2994 185
R16736 VDD.n2994 VDD.n354 185
R16737 VDD.n2996 VDD.n361 185
R16738 VDD.n3708 VDD.n361 185
R16739 VDD.n2998 VDD.n2997 185
R16740 VDD.n2997 VDD.n360 185
R16741 VDD.n2999 VDD.n367 185
R16742 VDD.n3702 VDD.n367 185
R16743 VDD.n3001 VDD.n3000 185
R16744 VDD.n3000 VDD.n366 185
R16745 VDD.n3002 VDD.n373 185
R16746 VDD.n3696 VDD.n373 185
R16747 VDD.n3004 VDD.n3003 185
R16748 VDD.n3003 VDD.n372 185
R16749 VDD.n3005 VDD.n379 185
R16750 VDD.n3690 VDD.n379 185
R16751 VDD.n3007 VDD.n3006 185
R16752 VDD.n3006 VDD.n378 185
R16753 VDD.n3008 VDD.n385 185
R16754 VDD.n3684 VDD.n385 185
R16755 VDD.n3010 VDD.n3009 185
R16756 VDD.n3009 VDD.n384 185
R16757 VDD.n3011 VDD.n391 185
R16758 VDD.n3678 VDD.n391 185
R16759 VDD.n3013 VDD.n3012 185
R16760 VDD.n3012 VDD.n390 185
R16761 VDD.n3014 VDD.n397 185
R16762 VDD.n3672 VDD.n397 185
R16763 VDD.n3016 VDD.n3015 185
R16764 VDD.n3015 VDD.n396 185
R16765 VDD.n3017 VDD.n403 185
R16766 VDD.n3666 VDD.n403 185
R16767 VDD.n3019 VDD.n3018 185
R16768 VDD.n3018 VDD.n402 185
R16769 VDD.n3020 VDD.n409 185
R16770 VDD.n3660 VDD.n409 185
R16771 VDD.n3022 VDD.n3021 185
R16772 VDD.n3021 VDD.n408 185
R16773 VDD.n3023 VDD.n415 185
R16774 VDD.n3654 VDD.n415 185
R16775 VDD.n3025 VDD.n3024 185
R16776 VDD.n3024 VDD.n414 185
R16777 VDD.n3026 VDD.n420 185
R16778 VDD.n3648 VDD.n420 185
R16779 VDD.n3028 VDD.n3027 185
R16780 VDD.n3027 VDD.n427 185
R16781 VDD.n3029 VDD.n425 185
R16782 VDD.n3642 VDD.n425 185
R16783 VDD.n3031 VDD.n3030 185
R16784 VDD.n3030 VDD.t132 185
R16785 VDD.n3032 VDD.n432 185
R16786 VDD.n3636 VDD.n432 185
R16787 VDD.n3034 VDD.n3033 185
R16788 VDD.n3033 VDD.n431 185
R16789 VDD.n3035 VDD.n438 185
R16790 VDD.n3630 VDD.n438 185
R16791 VDD.n3037 VDD.n3036 185
R16792 VDD.n3036 VDD.n437 185
R16793 VDD.n3038 VDD.n444 185
R16794 VDD.n3624 VDD.n444 185
R16795 VDD.n3040 VDD.n3039 185
R16796 VDD.n3039 VDD.n443 185
R16797 VDD.n3041 VDD.n450 185
R16798 VDD.n3618 VDD.n450 185
R16799 VDD.n3043 VDD.n3042 185
R16800 VDD.n3042 VDD.n449 185
R16801 VDD.n3044 VDD.n456 185
R16802 VDD.n3612 VDD.n456 185
R16803 VDD.n3046 VDD.n3045 185
R16804 VDD.n3045 VDD.n455 185
R16805 VDD.n3047 VDD.n462 185
R16806 VDD.n3606 VDD.n462 185
R16807 VDD.n3049 VDD.n3048 185
R16808 VDD.n3048 VDD.n461 185
R16809 VDD.n3050 VDD.n468 185
R16810 VDD.n3600 VDD.n468 185
R16811 VDD.n3052 VDD.n3051 185
R16812 VDD.n3051 VDD.n467 185
R16813 VDD.n3053 VDD.n474 185
R16814 VDD.n3594 VDD.n474 185
R16815 VDD.n3055 VDD.n3054 185
R16816 VDD.n3054 VDD.n473 185
R16817 VDD.n3056 VDD.n480 185
R16818 VDD.n3588 VDD.n480 185
R16819 VDD.n3058 VDD.n3057 185
R16820 VDD.n3057 VDD.n479 185
R16821 VDD.n3059 VDD.n485 185
R16822 VDD.n3582 VDD.n485 185
R16823 VDD.n3061 VDD.n3060 185
R16824 VDD.n3060 VDD.n493 185
R16825 VDD.n3062 VDD.n491 185
R16826 VDD.n3576 VDD.n491 185
R16827 VDD.n3064 VDD.n3063 185
R16828 VDD.n3063 VDD.n490 185
R16829 VDD.n3065 VDD.n498 185
R16830 VDD.n3570 VDD.n498 185
R16831 VDD.n3067 VDD.n3066 185
R16832 VDD.n3066 VDD.n497 185
R16833 VDD.n3068 VDD.n504 185
R16834 VDD.n3564 VDD.n504 185
R16835 VDD.n3070 VDD.n3069 185
R16836 VDD.n3069 VDD.n503 185
R16837 VDD.n3071 VDD.n510 185
R16838 VDD.n3558 VDD.n510 185
R16839 VDD.n3073 VDD.n3072 185
R16840 VDD.n3072 VDD.n509 185
R16841 VDD.n3074 VDD.n516 185
R16842 VDD.n3552 VDD.n516 185
R16843 VDD.n3076 VDD.n3075 185
R16844 VDD.n3075 VDD.n515 185
R16845 VDD.n3077 VDD.n522 185
R16846 VDD.n3546 VDD.n522 185
R16847 VDD.n3079 VDD.n3078 185
R16848 VDD.n3078 VDD.n521 185
R16849 VDD.n3080 VDD.n528 185
R16850 VDD.n3540 VDD.n528 185
R16851 VDD.n3082 VDD.n3081 185
R16852 VDD.n3081 VDD.n527 185
R16853 VDD.n3083 VDD.n533 185
R16854 VDD.n3534 VDD.n533 185
R16855 VDD.n3085 VDD.n3084 185
R16856 VDD.n3084 VDD.n541 185
R16857 VDD.n3086 VDD.n539 185
R16858 VDD.n3528 VDD.n539 185
R16859 VDD.n3088 VDD.n3087 185
R16860 VDD.n3087 VDD.n538 185
R16861 VDD.n3089 VDD.n546 185
R16862 VDD.n3522 VDD.n546 185
R16863 VDD.n3091 VDD.n3090 185
R16864 VDD.n3090 VDD.n545 185
R16865 VDD.n3092 VDD.n552 185
R16866 VDD.n3516 VDD.n552 185
R16867 VDD.n3094 VDD.n3093 185
R16868 VDD.n3093 VDD.n551 185
R16869 VDD.n3095 VDD.n558 185
R16870 VDD.n3510 VDD.n558 185
R16871 VDD.n3097 VDD.n3096 185
R16872 VDD.n3096 VDD.n557 185
R16873 VDD.n3098 VDD.n564 185
R16874 VDD.n3504 VDD.n564 185
R16875 VDD.n3100 VDD.n3099 185
R16876 VDD.n3099 VDD.n563 185
R16877 VDD.n3101 VDD.n570 185
R16878 VDD.n3498 VDD.n570 185
R16879 VDD.n3103 VDD.n3102 185
R16880 VDD.n3102 VDD.n569 185
R16881 VDD.n3104 VDD.n576 185
R16882 VDD.n3492 VDD.n576 185
R16883 VDD.n3106 VDD.n3105 185
R16884 VDD.n3105 VDD.n575 185
R16885 VDD.n3107 VDD.n582 185
R16886 VDD.n3486 VDD.n582 185
R16887 VDD.n3109 VDD.n3108 185
R16888 VDD.n3108 VDD.n581 185
R16889 VDD.n3110 VDD.n588 185
R16890 VDD.n3480 VDD.n588 185
R16891 VDD.n3112 VDD.n3111 185
R16892 VDD.n3111 VDD.n587 185
R16893 VDD.n3113 VDD.n594 185
R16894 VDD.n3474 VDD.n594 185
R16895 VDD.n3115 VDD.n3114 185
R16896 VDD.n3114 VDD.n593 185
R16897 VDD.n3116 VDD.n599 185
R16898 VDD.n3468 VDD.n599 185
R16899 VDD.n3371 VDD.n3370 185
R16900 VDD.n3370 VDD.n3369 185
R16901 VDD.n3372 VDD.n605 185
R16902 VDD.n3462 VDD.n605 185
R16903 VDD.n3374 VDD.n3373 185
R16904 VDD.n3373 VDD.n604 185
R16905 VDD.n3375 VDD.n611 185
R16906 VDD.n3456 VDD.n611 185
R16907 VDD.n3377 VDD.n3376 185
R16908 VDD.n3376 VDD.n610 185
R16909 VDD.n3378 VDD.n617 185
R16910 VDD.n3450 VDD.n617 185
R16911 VDD.n3380 VDD.n3379 185
R16912 VDD.n3379 VDD.n616 185
R16913 VDD.n3381 VDD.n623 185
R16914 VDD.n3444 VDD.n623 185
R16915 VDD.n3383 VDD.n3382 185
R16916 VDD.n3382 VDD.n622 185
R16917 VDD.n3384 VDD.n629 185
R16918 VDD.n3438 VDD.n629 185
R16919 VDD.n3386 VDD.n3385 185
R16920 VDD.n3385 VDD.n628 185
R16921 VDD.n3387 VDD.n635 185
R16922 VDD.n3432 VDD.n635 185
R16923 VDD.n3389 VDD.n3388 185
R16924 VDD.n3388 VDD.n634 185
R16925 VDD.n1803 VDD.n1802 185
R16926 VDD.n1804 VDD.n1803 185
R16927 VDD.n1234 VDD.n1232 185
R16928 VDD.n1232 VDD.n1231 185
R16929 VDD.n1767 VDD.n1766 185
R16930 VDD.n1766 VDD.n1765 185
R16931 VDD.n1237 VDD.n1236 185
R16932 VDD.n1238 VDD.n1237 185
R16933 VDD.n1754 VDD.n1753 185
R16934 VDD.n1755 VDD.n1754 185
R16935 VDD.n1247 VDD.n1246 185
R16936 VDD.n1246 VDD.n1245 185
R16937 VDD.n1749 VDD.n1748 185
R16938 VDD.n1748 VDD.n1747 185
R16939 VDD.n1250 VDD.n1249 185
R16940 VDD.t33 VDD.n1250 185
R16941 VDD.n1738 VDD.n1737 185
R16942 VDD.n1739 VDD.n1738 185
R16943 VDD.n1258 VDD.n1257 185
R16944 VDD.n1257 VDD.n1256 185
R16945 VDD.n1733 VDD.n1732 185
R16946 VDD.n1732 VDD.n1731 185
R16947 VDD.n1261 VDD.n1260 185
R16948 VDD.n1262 VDD.n1261 185
R16949 VDD.n1722 VDD.n1721 185
R16950 VDD.n1723 VDD.n1722 185
R16951 VDD.n1270 VDD.n1269 185
R16952 VDD.n1269 VDD.n1268 185
R16953 VDD.n1717 VDD.n1716 185
R16954 VDD.n1716 VDD.n1715 185
R16955 VDD.n1273 VDD.n1272 185
R16956 VDD.n1274 VDD.n1273 185
R16957 VDD.n1706 VDD.n1705 185
R16958 VDD.n1707 VDD.n1706 185
R16959 VDD.n1282 VDD.n1281 185
R16960 VDD.n1281 VDD.n1280 185
R16961 VDD.n1701 VDD.n1700 185
R16962 VDD.n1700 VDD.n1699 185
R16963 VDD.n1285 VDD.n1284 185
R16964 VDD.n1286 VDD.n1285 185
R16965 VDD.n1690 VDD.n1689 185
R16966 VDD.n1691 VDD.n1690 185
R16967 VDD.n1294 VDD.n1293 185
R16968 VDD.n1293 VDD.n1292 185
R16969 VDD.n1685 VDD.n1684 185
R16970 VDD.n1684 VDD.n1683 185
R16971 VDD.n1302 VDD.n1301 185
R16972 VDD.t135 VDD.n1302 185
R16973 VDD.n1674 VDD.n1673 185
R16974 VDD.n1675 VDD.n1674 185
R16975 VDD.n1310 VDD.n1309 185
R16976 VDD.n1309 VDD.n1308 185
R16977 VDD.n1669 VDD.n1668 185
R16978 VDD.n1668 VDD.n1667 185
R16979 VDD.n1313 VDD.n1312 185
R16980 VDD.n1314 VDD.n1313 185
R16981 VDD.n1658 VDD.n1657 185
R16982 VDD.n1659 VDD.n1658 185
R16983 VDD.n1322 VDD.n1321 185
R16984 VDD.n1321 VDD.n1320 185
R16985 VDD.n1653 VDD.n1652 185
R16986 VDD.n1652 VDD.n1651 185
R16987 VDD.n1325 VDD.n1324 185
R16988 VDD.n1326 VDD.n1325 185
R16989 VDD.n1642 VDD.n1641 185
R16990 VDD.n1643 VDD.n1642 185
R16991 VDD.n1334 VDD.n1333 185
R16992 VDD.n1333 VDD.n1332 185
R16993 VDD.n1637 VDD.n1636 185
R16994 VDD.n1636 VDD.n1635 185
R16995 VDD.n1337 VDD.n1336 185
R16996 VDD.n1338 VDD.n1337 185
R16997 VDD.n1626 VDD.n1625 185
R16998 VDD.n1627 VDD.n1626 185
R16999 VDD.n1346 VDD.n1345 185
R17000 VDD.n1345 VDD.n1344 185
R17001 VDD.n1621 VDD.n1620 185
R17002 VDD.n1620 VDD.n1619 185
R17003 VDD.n1349 VDD.n1348 185
R17004 VDD.t1 VDD.n1349 185
R17005 VDD.n1610 VDD.n1609 185
R17006 VDD.n1611 VDD.n1610 185
R17007 VDD.n1357 VDD.n1356 185
R17008 VDD.n1356 VDD.n1355 185
R17009 VDD.n1605 VDD.n1604 185
R17010 VDD.n1604 VDD.n1603 185
R17011 VDD.n1360 VDD.n1359 185
R17012 VDD.n1361 VDD.n1360 185
R17013 VDD.n1594 VDD.n1593 185
R17014 VDD.n1595 VDD.n1594 185
R17015 VDD.n1369 VDD.n1368 185
R17016 VDD.n1368 VDD.n1367 185
R17017 VDD.n1589 VDD.n1588 185
R17018 VDD.n1588 VDD.n1587 185
R17019 VDD.n1446 VDD.n1371 185
R17020 VDD.n1450 VDD.n1448 185
R17021 VDD.n1451 VDD.n1445 185
R17022 VDD.n1451 VDD.n1372 185
R17023 VDD.n1454 VDD.n1453 185
R17024 VDD.n1443 VDD.n1442 185
R17025 VDD.n1461 VDD.n1460 185
R17026 VDD.n1463 VDD.n1441 185
R17027 VDD.n1464 VDD.n1440 185
R17028 VDD.n1467 VDD.n1466 185
R17029 VDD.n1468 VDD.n1437 185
R17030 VDD.n1434 VDD.n1433 185
R17031 VDD.n1473 VDD.n1472 185
R17032 VDD.n1475 VDD.n1432 185
R17033 VDD.n1478 VDD.n1477 185
R17034 VDD.n1430 VDD.n1429 185
R17035 VDD.n1484 VDD.n1483 185
R17036 VDD.n1486 VDD.n1428 185
R17037 VDD.n1487 VDD.n1425 185
R17038 VDD.n1490 VDD.n1489 185
R17039 VDD.n1427 VDD.n1423 185
R17040 VDD.n1494 VDD.n1419 185
R17041 VDD.n1496 VDD.n1495 185
R17042 VDD.n1498 VDD.n1418 185
R17043 VDD.n1501 VDD.n1500 185
R17044 VDD.n1416 VDD.n1415 185
R17045 VDD.n1506 VDD.n1505 185
R17046 VDD.n1508 VDD.n1414 185
R17047 VDD.n1511 VDD.n1510 185
R17048 VDD.n1412 VDD.n1411 185
R17049 VDD.n1518 VDD.n1517 185
R17050 VDD.n1520 VDD.n1410 185
R17051 VDD.n1521 VDD.n1409 185
R17052 VDD.n1524 VDD.n1523 185
R17053 VDD.n1525 VDD.n1406 185
R17054 VDD.n1403 VDD.n1402 185
R17055 VDD.n1530 VDD.n1529 185
R17056 VDD.n1532 VDD.n1401 185
R17057 VDD.n1535 VDD.n1534 185
R17058 VDD.n1399 VDD.n1398 185
R17059 VDD.n1540 VDD.n1539 185
R17060 VDD.n1542 VDD.n1397 185
R17061 VDD.n1545 VDD.n1544 185
R17062 VDD.n1395 VDD.n1394 185
R17063 VDD.n1550 VDD.n1549 185
R17064 VDD.n1552 VDD.n1393 185
R17065 VDD.n1555 VDD.n1554 185
R17066 VDD.n1388 VDD.n1387 185
R17067 VDD.n1560 VDD.n1559 185
R17068 VDD.n1562 VDD.n1386 185
R17069 VDD.n1565 VDD.n1564 185
R17070 VDD.n1384 VDD.n1383 185
R17071 VDD.n1570 VDD.n1569 185
R17072 VDD.n1572 VDD.n1382 185
R17073 VDD.n1576 VDD.n1575 185
R17074 VDD.n1573 VDD.n1378 185
R17075 VDD.n1580 VDD.n1380 185
R17076 VDD.n1581 VDD.n1375 185
R17077 VDD.n1582 VDD.n1373 185
R17078 VDD.n1373 VDD.n1372 185
R17079 VDD.n1806 VDD.n1224 185
R17080 VDD.n1809 VDD.n1808 185
R17081 VDD.n1228 VDD.n1222 185
R17082 VDD.n1813 VDD.n1221 185
R17083 VDD.n1814 VDD.n1220 185
R17084 VDD.n1815 VDD.n1218 185
R17085 VDD.n1217 VDD.n1214 185
R17086 VDD.n1819 VDD.n1213 185
R17087 VDD.n1820 VDD.n1212 185
R17088 VDD.n1821 VDD.n1210 185
R17089 VDD.n1209 VDD.n1206 185
R17090 VDD.n1205 VDD.n1201 185
R17091 VDD.n1826 VDD.n1825 185
R17092 VDD.n1828 VDD.n1199 185
R17093 VDD.n1830 VDD.n1829 185
R17094 VDD.n1831 VDD.n1194 185
R17095 VDD.n1833 VDD.n1832 185
R17096 VDD.n1835 VDD.n1192 185
R17097 VDD.n1837 VDD.n1836 185
R17098 VDD.n1838 VDD.n1188 185
R17099 VDD.n1840 VDD.n1839 185
R17100 VDD.n1842 VDD.n1186 185
R17101 VDD.n1844 VDD.n1843 185
R17102 VDD.n1181 VDD.n1180 185
R17103 VDD.n1849 VDD.n1848 185
R17104 VDD.n1851 VDD.n1178 185
R17105 VDD.n1853 VDD.n1852 185
R17106 VDD.n1854 VDD.n1173 185
R17107 VDD.n1856 VDD.n1855 185
R17108 VDD.n1858 VDD.n1171 185
R17109 VDD.n1860 VDD.n1859 185
R17110 VDD.n1861 VDD.n1167 185
R17111 VDD.n1863 VDD.n1862 185
R17112 VDD.n1865 VDD.n1165 185
R17113 VDD.n1867 VDD.n1866 185
R17114 VDD.n1160 VDD.n1159 185
R17115 VDD.n1872 VDD.n1871 185
R17116 VDD.n1874 VDD.n1157 185
R17117 VDD.n1876 VDD.n1875 185
R17118 VDD.n1877 VDD.n1152 185
R17119 VDD.n1879 VDD.n1878 185
R17120 VDD.n1881 VDD.n1150 185
R17121 VDD.n1883 VDD.n1882 185
R17122 VDD.n1884 VDD.n1148 185
R17123 VDD.n1886 VDD.n1885 185
R17124 VDD.n1888 VDD.n1147 185
R17125 VDD.n1889 VDD.n1141 185
R17126 VDD.n1892 VDD.n1891 185
R17127 VDD.n1145 VDD.n1144 185
R17128 VDD.n1786 VDD.n1783 185
R17129 VDD.n1788 VDD.n1787 185
R17130 VDD.n1789 VDD.n1776 185
R17131 VDD.n1791 VDD.n1790 185
R17132 VDD.n1793 VDD.n1775 185
R17133 VDD.n1794 VDD.n1774 185
R17134 VDD.n1797 VDD.n1796 185
R17135 VDD.n1798 VDD.n1772 185
R17136 VDD.n1799 VDD.n1233 185
R17137 VDD.n1805 VDD.n1230 185
R17138 VDD.n1805 VDD.n1804 185
R17139 VDD.n1241 VDD.n1229 185
R17140 VDD.n1231 VDD.n1229 185
R17141 VDD.n1764 VDD.n1763 185
R17142 VDD.n1765 VDD.n1764 185
R17143 VDD.n1240 VDD.n1239 185
R17144 VDD.n1239 VDD.n1238 185
R17145 VDD.n1757 VDD.n1756 185
R17146 VDD.n1756 VDD.n1755 185
R17147 VDD.n1244 VDD.n1243 185
R17148 VDD.n1245 VDD.n1244 185
R17149 VDD.n1746 VDD.n1745 185
R17150 VDD.n1747 VDD.n1746 185
R17151 VDD.n1252 VDD.n1251 185
R17152 VDD.n1251 VDD.t33 185
R17153 VDD.n1741 VDD.n1740 185
R17154 VDD.n1740 VDD.n1739 185
R17155 VDD.n1255 VDD.n1254 185
R17156 VDD.n1256 VDD.n1255 185
R17157 VDD.n1730 VDD.n1729 185
R17158 VDD.n1731 VDD.n1730 185
R17159 VDD.n1264 VDD.n1263 185
R17160 VDD.n1263 VDD.n1262 185
R17161 VDD.n1725 VDD.n1724 185
R17162 VDD.n1724 VDD.n1723 185
R17163 VDD.n1267 VDD.n1266 185
R17164 VDD.n1268 VDD.n1267 185
R17165 VDD.n1714 VDD.n1713 185
R17166 VDD.n1715 VDD.n1714 185
R17167 VDD.n1276 VDD.n1275 185
R17168 VDD.n1275 VDD.n1274 185
R17169 VDD.n1709 VDD.n1708 185
R17170 VDD.n1708 VDD.n1707 185
R17171 VDD.n1279 VDD.n1278 185
R17172 VDD.n1280 VDD.n1279 185
R17173 VDD.n1698 VDD.n1697 185
R17174 VDD.n1699 VDD.n1698 185
R17175 VDD.n1288 VDD.n1287 185
R17176 VDD.n1287 VDD.n1286 185
R17177 VDD.n1693 VDD.n1692 185
R17178 VDD.n1692 VDD.n1691 185
R17179 VDD.n1291 VDD.n1290 185
R17180 VDD.n1292 VDD.n1291 185
R17181 VDD.n1682 VDD.n1681 185
R17182 VDD.n1683 VDD.n1682 185
R17183 VDD.n1304 VDD.n1303 185
R17184 VDD.n1303 VDD.t135 185
R17185 VDD.n1677 VDD.n1676 185
R17186 VDD.n1676 VDD.n1675 185
R17187 VDD.n1307 VDD.n1306 185
R17188 VDD.n1308 VDD.n1307 185
R17189 VDD.n1666 VDD.n1665 185
R17190 VDD.n1667 VDD.n1666 185
R17191 VDD.n1316 VDD.n1315 185
R17192 VDD.n1315 VDD.n1314 185
R17193 VDD.n1661 VDD.n1660 185
R17194 VDD.n1660 VDD.n1659 185
R17195 VDD.n1319 VDD.n1318 185
R17196 VDD.n1320 VDD.n1319 185
R17197 VDD.n1650 VDD.n1649 185
R17198 VDD.n1651 VDD.n1650 185
R17199 VDD.n1328 VDD.n1327 185
R17200 VDD.n1327 VDD.n1326 185
R17201 VDD.n1645 VDD.n1644 185
R17202 VDD.n1644 VDD.n1643 185
R17203 VDD.n1331 VDD.n1330 185
R17204 VDD.n1332 VDD.n1331 185
R17205 VDD.n1634 VDD.n1633 185
R17206 VDD.n1635 VDD.n1634 185
R17207 VDD.n1340 VDD.n1339 185
R17208 VDD.n1339 VDD.n1338 185
R17209 VDD.n1629 VDD.n1628 185
R17210 VDD.n1628 VDD.n1627 185
R17211 VDD.n1343 VDD.n1342 185
R17212 VDD.n1344 VDD.n1343 185
R17213 VDD.n1618 VDD.n1617 185
R17214 VDD.n1619 VDD.n1618 185
R17215 VDD.n1351 VDD.n1350 185
R17216 VDD.n1350 VDD.t1 185
R17217 VDD.n1613 VDD.n1612 185
R17218 VDD.n1612 VDD.n1611 185
R17219 VDD.n1354 VDD.n1353 185
R17220 VDD.n1355 VDD.n1354 185
R17221 VDD.n1602 VDD.n1601 185
R17222 VDD.n1603 VDD.n1602 185
R17223 VDD.n1363 VDD.n1362 185
R17224 VDD.n1362 VDD.n1361 185
R17225 VDD.n1597 VDD.n1596 185
R17226 VDD.n1596 VDD.n1595 185
R17227 VDD.n1366 VDD.n1365 185
R17228 VDD.n1367 VDD.n1366 185
R17229 VDD.n1586 VDD.n1585 185
R17230 VDD.n1587 VDD.n1586 185
R17231 VDD.n4077 VDD.n4076 185
R17232 VDD.n99 VDD.n98 185
R17233 VDD.n4073 VDD.n4072 185
R17234 VDD.n4074 VDD.n4073 185
R17235 VDD.n4071 VDD.n128 185
R17236 VDD.n4070 VDD.n4069 185
R17237 VDD.n4068 VDD.n4067 185
R17238 VDD.n4066 VDD.n4065 185
R17239 VDD.n4064 VDD.n4063 185
R17240 VDD.n4062 VDD.n4061 185
R17241 VDD.n4060 VDD.n4059 185
R17242 VDD.n4058 VDD.n4057 185
R17243 VDD.n4056 VDD.n4055 185
R17244 VDD.n4054 VDD.n4053 185
R17245 VDD.n4052 VDD.n4051 185
R17246 VDD.n4050 VDD.n4049 185
R17247 VDD.n4048 VDD.n4047 185
R17248 VDD.n4046 VDD.n4045 185
R17249 VDD.n4044 VDD.n4043 185
R17250 VDD.n4042 VDD.n4041 185
R17251 VDD.n4040 VDD.n4039 185
R17252 VDD.n4038 VDD.n4037 185
R17253 VDD.n4036 VDD.n4035 185
R17254 VDD.n4027 VDD.n148 185
R17255 VDD.n4029 VDD.n4028 185
R17256 VDD.n4026 VDD.n4025 185
R17257 VDD.n4024 VDD.n4023 185
R17258 VDD.n4022 VDD.n4021 185
R17259 VDD.n4020 VDD.n4019 185
R17260 VDD.n4018 VDD.n4017 185
R17261 VDD.n4016 VDD.n4015 185
R17262 VDD.n4014 VDD.n4013 185
R17263 VDD.n4012 VDD.n4011 185
R17264 VDD.n4010 VDD.n4009 185
R17265 VDD.n4008 VDD.n4007 185
R17266 VDD.n4006 VDD.n4005 185
R17267 VDD.n4004 VDD.n4003 185
R17268 VDD.n4002 VDD.n4001 185
R17269 VDD.n4000 VDD.n3999 185
R17270 VDD.n3998 VDD.n3997 185
R17271 VDD.n3996 VDD.n3995 185
R17272 VDD.n3994 VDD.n3993 185
R17273 VDD.n3992 VDD.n3991 185
R17274 VDD.n3990 VDD.n3989 185
R17275 VDD.n3988 VDD.n3987 185
R17276 VDD.n3947 VDD.n170 185
R17277 VDD.n3949 VDD.n3948 185
R17278 VDD.n3951 VDD.n3950 185
R17279 VDD.n3983 VDD.n3952 185
R17280 VDD.n3982 VDD.n3981 185
R17281 VDD.n3980 VDD.n3979 185
R17282 VDD.n3978 VDD.n3977 185
R17283 VDD.n3976 VDD.n3975 185
R17284 VDD.n3974 VDD.n3973 185
R17285 VDD.n3972 VDD.n3971 185
R17286 VDD.n3970 VDD.n3969 185
R17287 VDD.n3968 VDD.n3967 185
R17288 VDD.n3966 VDD.n3961 185
R17289 VDD.n3960 VDD.n127 185
R17290 VDD.n4074 VDD.n127 185
R17291 VDD.n4380 VDD.n4379 185
R17292 VDD.n4382 VDD.n4365 185
R17293 VDD.n4384 VDD.n4383 185
R17294 VDD.n4385 VDD.n4358 185
R17295 VDD.n4387 VDD.n4386 185
R17296 VDD.n4389 VDD.n4356 185
R17297 VDD.n4391 VDD.n4390 185
R17298 VDD.n4392 VDD.n4351 185
R17299 VDD.n4394 VDD.n4393 185
R17300 VDD.n4396 VDD.n4349 185
R17301 VDD.n4398 VDD.n4397 185
R17302 VDD.n4399 VDD.n4341 185
R17303 VDD.n4401 VDD.n4400 185
R17304 VDD.n4403 VDD.n4339 185
R17305 VDD.n4405 VDD.n4404 185
R17306 VDD.n4406 VDD.n4334 185
R17307 VDD.n4408 VDD.n4407 185
R17308 VDD.n4410 VDD.n4332 185
R17309 VDD.n4412 VDD.n4411 185
R17310 VDD.n4413 VDD.n4328 185
R17311 VDD.n4415 VDD.n4414 185
R17312 VDD.n4417 VDD.n4326 185
R17313 VDD.n4419 VDD.n4418 185
R17314 VDD.n4321 VDD.n4320 185
R17315 VDD.n4424 VDD.n4423 185
R17316 VDD.n4426 VDD.n4318 185
R17317 VDD.n4428 VDD.n4427 185
R17318 VDD.n4429 VDD.n4313 185
R17319 VDD.n4431 VDD.n4430 185
R17320 VDD.n4433 VDD.n4311 185
R17321 VDD.n4435 VDD.n4434 185
R17322 VDD.n4436 VDD.n4307 185
R17323 VDD.n4438 VDD.n4437 185
R17324 VDD.n4440 VDD.n4305 185
R17325 VDD.n4442 VDD.n4441 185
R17326 VDD.n4300 VDD.n4299 185
R17327 VDD.n4447 VDD.n4446 185
R17328 VDD.n4449 VDD.n4297 185
R17329 VDD.n4451 VDD.n4450 185
R17330 VDD.n4452 VDD.n4292 185
R17331 VDD.n4454 VDD.n4453 185
R17332 VDD.n4456 VDD.n4290 185
R17333 VDD.n4458 VDD.n4457 185
R17334 VDD.n4459 VDD.n4286 185
R17335 VDD.n4461 VDD.n4460 185
R17336 VDD.n4463 VDD.n4283 185
R17337 VDD.n4465 VDD.n4464 185
R17338 VDD.n4284 VDD.n4277 185
R17339 VDD.n4469 VDD.n4281 185
R17340 VDD.n4470 VDD.n4273 185
R17341 VDD.n4472 VDD.n4471 185
R17342 VDD.n4474 VDD.n4271 185
R17343 VDD.n4476 VDD.n4475 185
R17344 VDD.n4477 VDD.n4266 185
R17345 VDD.n4479 VDD.n4478 185
R17346 VDD.n4481 VDD.n4265 185
R17347 VDD.n4482 VDD.n4263 185
R17348 VDD.n4485 VDD.n4484 185
R17349 VDD.n4376 VDD.n4367 185
R17350 VDD.n4367 VDD.n4258 185
R17351 VDD.n4375 VDD.n4257 185
R17352 VDD.n4491 VDD.n4257 185
R17353 VDD.n4374 VDD.n4256 185
R17354 VDD.n4492 VDD.n4256 185
R17355 VDD.n4370 VDD.n4255 185
R17356 VDD.n4493 VDD.n4255 185
R17357 VDD.n4246 VDD.n4245 185
R17358 VDD.n4247 VDD.n4246 185
R17359 VDD.n4501 VDD.n4500 185
R17360 VDD.n4500 VDD.n4499 185
R17361 VDD.n4502 VDD.n4214 185
R17362 VDD.n4214 VDD.n4212 185
R17363 VDD.n4504 VDD.n4503 185
R17364 VDD.t43 VDD.n4504 185
R17365 VDD.n4215 VDD.n4213 185
R17366 VDD.n4213 VDD.n4204 185
R17367 VDD.n4239 VDD.n4203 185
R17368 VDD.n4510 VDD.n4203 185
R17369 VDD.n4238 VDD.n4202 185
R17370 VDD.n4511 VDD.n4202 185
R17371 VDD.n4237 VDD.n4201 185
R17372 VDD.n4512 VDD.n4201 185
R17373 VDD.n4218 VDD.n4217 185
R17374 VDD.n4217 VDD.n4193 185
R17375 VDD.n4233 VDD.n4192 185
R17376 VDD.n4518 VDD.n4192 185
R17377 VDD.n4232 VDD.n4191 185
R17378 VDD.n4519 VDD.n4191 185
R17379 VDD.n4231 VDD.n4190 185
R17380 VDD.n4520 VDD.n4190 185
R17381 VDD.n4221 VDD.n4220 185
R17382 VDD.n4220 VDD.n4182 185
R17383 VDD.n4227 VDD.n4181 185
R17384 VDD.n4526 VDD.n4181 185
R17385 VDD.n4226 VDD.n4180 185
R17386 VDD.n4527 VDD.n4180 185
R17387 VDD.n4225 VDD.n4179 185
R17388 VDD.n4528 VDD.n4179 185
R17389 VDD.n4171 VDD.n4170 185
R17390 VDD.n4172 VDD.n4171 185
R17391 VDD.n4536 VDD.n4535 185
R17392 VDD.n4535 VDD.n4534 185
R17393 VDD.n4537 VDD.n29 185
R17394 VDD.n29 VDD.n27 185
R17395 VDD.n4539 VDD.n4538 185
R17396 VDD.t137 VDD.n4539 185
R17397 VDD.n30 VDD.n28 185
R17398 VDD.n28 VDD.n26 185
R17399 VDD.n4164 VDD.n4163 185
R17400 VDD.n4163 VDD.n4162 185
R17401 VDD.n33 VDD.n32 185
R17402 VDD.n34 VDD.n33 185
R17403 VDD.n4153 VDD.n4152 185
R17404 VDD.n4154 VDD.n4153 185
R17405 VDD.n42 VDD.n41 185
R17406 VDD.n41 VDD.n40 185
R17407 VDD.n4148 VDD.n4147 185
R17408 VDD.n4147 VDD.n4146 185
R17409 VDD.n45 VDD.n44 185
R17410 VDD.n46 VDD.n45 185
R17411 VDD.n4137 VDD.n4136 185
R17412 VDD.n4138 VDD.n4137 185
R17413 VDD.n54 VDD.n53 185
R17414 VDD.n53 VDD.n52 185
R17415 VDD.n4132 VDD.n4131 185
R17416 VDD.n4131 VDD.n4130 185
R17417 VDD.n57 VDD.n56 185
R17418 VDD.n58 VDD.n57 185
R17419 VDD.n4121 VDD.n4120 185
R17420 VDD.n4122 VDD.n4121 185
R17421 VDD.n66 VDD.n65 185
R17422 VDD.n65 VDD.n64 185
R17423 VDD.n4116 VDD.n4115 185
R17424 VDD.n4115 VDD.n4114 185
R17425 VDD.n69 VDD.n68 185
R17426 VDD.n70 VDD.n69 185
R17427 VDD.n4106 VDD.n4105 185
R17428 VDD.t11 VDD.n4106 185
R17429 VDD.n78 VDD.n77 185
R17430 VDD.n77 VDD.n76 185
R17431 VDD.n4101 VDD.n4100 185
R17432 VDD.n4100 VDD.n4099 185
R17433 VDD.n81 VDD.n80 185
R17434 VDD.n82 VDD.n81 185
R17435 VDD.n4090 VDD.n4089 185
R17436 VDD.n4091 VDD.n4090 185
R17437 VDD.n90 VDD.n89 185
R17438 VDD.n89 VDD.n88 185
R17439 VDD.n4085 VDD.n4084 185
R17440 VDD.n4084 VDD.n4083 185
R17441 VDD.n93 VDD.n92 185
R17442 VDD.n94 VDD.n93 185
R17443 VDD.n96 VDD.n95 185
R17444 VDD.n95 VDD.n94 185
R17445 VDD.n4082 VDD.n4081 185
R17446 VDD.n4083 VDD.n4082 185
R17447 VDD.n87 VDD.n86 185
R17448 VDD.n88 VDD.n87 185
R17449 VDD.n4093 VDD.n4092 185
R17450 VDD.n4092 VDD.n4091 185
R17451 VDD.n84 VDD.n83 185
R17452 VDD.n83 VDD.n82 185
R17453 VDD.n4098 VDD.n4097 185
R17454 VDD.n4099 VDD.n4098 185
R17455 VDD.n75 VDD.n74 185
R17456 VDD.n76 VDD.n75 185
R17457 VDD.n4108 VDD.n4107 185
R17458 VDD.n4107 VDD.t11 185
R17459 VDD.n72 VDD.n71 185
R17460 VDD.n71 VDD.n70 185
R17461 VDD.n4113 VDD.n4112 185
R17462 VDD.n4114 VDD.n4113 185
R17463 VDD.n63 VDD.n62 185
R17464 VDD.n64 VDD.n63 185
R17465 VDD.n4124 VDD.n4123 185
R17466 VDD.n4123 VDD.n4122 185
R17467 VDD.n60 VDD.n59 185
R17468 VDD.n59 VDD.n58 185
R17469 VDD.n4129 VDD.n4128 185
R17470 VDD.n4130 VDD.n4129 185
R17471 VDD.n51 VDD.n50 185
R17472 VDD.n52 VDD.n51 185
R17473 VDD.n4140 VDD.n4139 185
R17474 VDD.n4139 VDD.n4138 185
R17475 VDD.n48 VDD.n47 185
R17476 VDD.n47 VDD.n46 185
R17477 VDD.n4145 VDD.n4144 185
R17478 VDD.n4146 VDD.n4145 185
R17479 VDD.n39 VDD.n38 185
R17480 VDD.n40 VDD.n39 185
R17481 VDD.n4156 VDD.n4155 185
R17482 VDD.n4155 VDD.n4154 185
R17483 VDD.n36 VDD.n35 185
R17484 VDD.n35 VDD.n34 185
R17485 VDD.n4161 VDD.n4160 185
R17486 VDD.n4162 VDD.n4161 185
R17487 VDD.n24 VDD.n22 185
R17488 VDD.n26 VDD.n24 185
R17489 VDD.n4541 VDD.n4540 185
R17490 VDD.n4540 VDD.t137 185
R17491 VDD.n25 VDD.n23 185
R17492 VDD.n27 VDD.n25 185
R17493 VDD.n4533 VDD.n4532 185
R17494 VDD.n4534 VDD.n4533 185
R17495 VDD.n4531 VDD.n4173 185
R17496 VDD.n4173 VDD.n4172 185
R17497 VDD.n4530 VDD.n4529 185
R17498 VDD.n4529 VDD.n4528 185
R17499 VDD.n4178 VDD.n4177 185
R17500 VDD.n4527 VDD.n4178 185
R17501 VDD.n4525 VDD.n4524 185
R17502 VDD.n4526 VDD.n4525 185
R17503 VDD.n4523 VDD.n4183 185
R17504 VDD.n4183 VDD.n4182 185
R17505 VDD.n4522 VDD.n4521 185
R17506 VDD.n4521 VDD.n4520 185
R17507 VDD.n4189 VDD.n4188 185
R17508 VDD.n4519 VDD.n4189 185
R17509 VDD.n4517 VDD.n4516 185
R17510 VDD.n4518 VDD.n4517 185
R17511 VDD.n4515 VDD.n4194 185
R17512 VDD.n4194 VDD.n4193 185
R17513 VDD.n4514 VDD.n4513 185
R17514 VDD.n4513 VDD.n4512 185
R17515 VDD.n4200 VDD.n4199 185
R17516 VDD.n4511 VDD.n4200 185
R17517 VDD.n4509 VDD.n4508 185
R17518 VDD.n4510 VDD.n4509 185
R17519 VDD.n4507 VDD.n4205 185
R17520 VDD.n4205 VDD.n4204 185
R17521 VDD.n4506 VDD.n4505 185
R17522 VDD.n4505 VDD.t43 185
R17523 VDD.n4211 VDD.n4210 185
R17524 VDD.n4212 VDD.n4211 185
R17525 VDD.n4498 VDD.n4497 185
R17526 VDD.n4499 VDD.n4498 185
R17527 VDD.n4496 VDD.n4248 185
R17528 VDD.n4248 VDD.n4247 185
R17529 VDD.n4495 VDD.n4494 185
R17530 VDD.n4494 VDD.n4493 185
R17531 VDD.n4254 VDD.n4253 185
R17532 VDD.n4492 VDD.n4254 185
R17533 VDD.n4490 VDD.n4489 185
R17534 VDD.n4491 VDD.n4490 185
R17535 VDD.n4488 VDD.n4259 185
R17536 VDD.n4259 VDD.n4258 185
R17537 VDD.n661 VDD.n659 185
R17538 VDD.n659 VDD.n640 185
R17539 VDD.n2804 VDD.n668 185
R17540 VDD.n2863 VDD.n668 185
R17541 VDD.n2806 VDD.n2805 185
R17542 VDD.n2805 VDD.n666 185
R17543 VDD.n2807 VDD.n679 185
R17544 VDD.n2817 VDD.n679 185
R17545 VDD.n2808 VDD.n687 185
R17546 VDD.n687 VDD.n677 185
R17547 VDD.n2810 VDD.n2809 185
R17548 VDD.n2811 VDD.n2810 185
R17549 VDD.n2803 VDD.n686 185
R17550 VDD.n686 VDD.n683 185
R17551 VDD.n2802 VDD.n2801 185
R17552 VDD.n2801 VDD.n2800 185
R17553 VDD.n689 VDD.n688 185
R17554 VDD.n690 VDD.n689 185
R17555 VDD.n2793 VDD.n2792 185
R17556 VDD.n2794 VDD.n2793 185
R17557 VDD.n2791 VDD.n699 185
R17558 VDD.n699 VDD.n696 185
R17559 VDD.n2790 VDD.n2789 185
R17560 VDD.n2789 VDD.n2788 185
R17561 VDD.n701 VDD.n700 185
R17562 VDD.n2147 VDD.n701 185
R17563 VDD.n2781 VDD.n2780 185
R17564 VDD.n2782 VDD.n2781 185
R17565 VDD.n2779 VDD.n710 185
R17566 VDD.n710 VDD.n707 185
R17567 VDD.n2778 VDD.n2777 185
R17568 VDD.n2777 VDD.n2776 185
R17569 VDD.n712 VDD.n711 185
R17570 VDD.n713 VDD.n712 185
R17571 VDD.n2769 VDD.n2768 185
R17572 VDD.n2770 VDD.n2769 185
R17573 VDD.n2767 VDD.n722 185
R17574 VDD.n722 VDD.n719 185
R17575 VDD.n2766 VDD.n2765 185
R17576 VDD.n2765 VDD.n2764 185
R17577 VDD.n724 VDD.n723 185
R17578 VDD.n725 VDD.n724 185
R17579 VDD.n2757 VDD.n2756 185
R17580 VDD.n2758 VDD.n2757 185
R17581 VDD.n2755 VDD.n734 185
R17582 VDD.n734 VDD.n731 185
R17583 VDD.n2754 VDD.n2753 185
R17584 VDD.n2753 VDD.n2752 185
R17585 VDD.n736 VDD.n735 185
R17586 VDD.n737 VDD.n736 185
R17587 VDD.n2745 VDD.n2744 185
R17588 VDD.n2746 VDD.n2745 185
R17589 VDD.n2743 VDD.n746 185
R17590 VDD.n746 VDD.n743 185
R17591 VDD.n2742 VDD.n2741 185
R17592 VDD.n2741 VDD.n2740 185
R17593 VDD.n748 VDD.n747 185
R17594 VDD.n749 VDD.n748 185
R17595 VDD.n2733 VDD.n2732 185
R17596 VDD.n2734 VDD.n2733 185
R17597 VDD.n2731 VDD.n758 185
R17598 VDD.n758 VDD.n755 185
R17599 VDD.n2730 VDD.n2729 185
R17600 VDD.n2729 VDD.n2728 185
R17601 VDD.n760 VDD.n759 185
R17602 VDD.n769 VDD.n760 185
R17603 VDD.n2721 VDD.n2720 185
R17604 VDD.n2722 VDD.n2721 185
R17605 VDD.n2719 VDD.n770 185
R17606 VDD.n770 VDD.n766 185
R17607 VDD.n2718 VDD.n2717 185
R17608 VDD.n2717 VDD.n2716 185
R17609 VDD.n772 VDD.n771 185
R17610 VDD.n773 VDD.n772 185
R17611 VDD.n2709 VDD.n2708 185
R17612 VDD.n2710 VDD.n2709 185
R17613 VDD.n2707 VDD.n782 185
R17614 VDD.n782 VDD.n779 185
R17615 VDD.n2706 VDD.n2705 185
R17616 VDD.n2705 VDD.n2704 185
R17617 VDD.n784 VDD.n783 185
R17618 VDD.n785 VDD.n784 185
R17619 VDD.n2697 VDD.n2696 185
R17620 VDD.n2698 VDD.n2697 185
R17621 VDD.n2695 VDD.n794 185
R17622 VDD.n794 VDD.n791 185
R17623 VDD.n2694 VDD.n2693 185
R17624 VDD.n2693 VDD.n2692 185
R17625 VDD.n796 VDD.n795 185
R17626 VDD.n797 VDD.n796 185
R17627 VDD.n2685 VDD.n2684 185
R17628 VDD.n2686 VDD.n2685 185
R17629 VDD.n2683 VDD.n806 185
R17630 VDD.n806 VDD.n803 185
R17631 VDD.n2682 VDD.n2681 185
R17632 VDD.n2681 VDD.n2680 185
R17633 VDD.n808 VDD.n807 185
R17634 VDD.n809 VDD.n808 185
R17635 VDD.n2673 VDD.n2672 185
R17636 VDD.n2674 VDD.n2673 185
R17637 VDD.n2671 VDD.n818 185
R17638 VDD.n818 VDD.n815 185
R17639 VDD.n2670 VDD.n2669 185
R17640 VDD.n2669 VDD.n2668 185
R17641 VDD.n820 VDD.n819 185
R17642 VDD.n821 VDD.n820 185
R17643 VDD.n2661 VDD.n2660 185
R17644 VDD.n2662 VDD.n2661 185
R17645 VDD.n2659 VDD.n829 185
R17646 VDD.n835 VDD.n829 185
R17647 VDD.n2658 VDD.n2657 185
R17648 VDD.n2657 VDD.n2656 185
R17649 VDD.n831 VDD.n830 185
R17650 VDD.n832 VDD.n831 185
R17651 VDD.n2649 VDD.n2648 185
R17652 VDD.n2650 VDD.n2649 185
R17653 VDD.n2647 VDD.n842 185
R17654 VDD.n842 VDD.n839 185
R17655 VDD.n2646 VDD.n2645 185
R17656 VDD.n2645 VDD.n2644 185
R17657 VDD.n844 VDD.n843 185
R17658 VDD.n845 VDD.n844 185
R17659 VDD.n2637 VDD.n2636 185
R17660 VDD.n2638 VDD.n2637 185
R17661 VDD.n2635 VDD.n854 185
R17662 VDD.n854 VDD.n851 185
R17663 VDD.n2634 VDD.n2633 185
R17664 VDD.n2633 VDD.n2632 185
R17665 VDD.n856 VDD.n855 185
R17666 VDD.n857 VDD.n856 185
R17667 VDD.n2625 VDD.n2624 185
R17668 VDD.n2626 VDD.n2625 185
R17669 VDD.n2623 VDD.n866 185
R17670 VDD.n866 VDD.n863 185
R17671 VDD.n2622 VDD.n2621 185
R17672 VDD.n2621 VDD.n2620 185
R17673 VDD.n868 VDD.n867 185
R17674 VDD.n869 VDD.n868 185
R17675 VDD.n2613 VDD.n2612 185
R17676 VDD.n2614 VDD.n2613 185
R17677 VDD.n2611 VDD.n877 185
R17678 VDD.n877 VDD.t92 185
R17679 VDD.n2610 VDD.n2609 185
R17680 VDD.n2609 VDD.n2608 185
R17681 VDD.n879 VDD.n878 185
R17682 VDD.n880 VDD.n879 185
R17683 VDD.n2601 VDD.n2600 185
R17684 VDD.n2602 VDD.n2601 185
R17685 VDD.n2599 VDD.n889 185
R17686 VDD.n889 VDD.n886 185
R17687 VDD.n2598 VDD.n2597 185
R17688 VDD.n2597 VDD.n2596 185
R17689 VDD.n891 VDD.n890 185
R17690 VDD.n892 VDD.n891 185
R17691 VDD.n2589 VDD.n2588 185
R17692 VDD.n2590 VDD.n2589 185
R17693 VDD.n2587 VDD.n901 185
R17694 VDD.n901 VDD.n898 185
R17695 VDD.n2586 VDD.n2585 185
R17696 VDD.n2585 VDD.n2584 185
R17697 VDD.n903 VDD.n902 185
R17698 VDD.n904 VDD.n903 185
R17699 VDD.n2577 VDD.n2576 185
R17700 VDD.n2578 VDD.n2577 185
R17701 VDD.n2575 VDD.n913 185
R17702 VDD.n913 VDD.n910 185
R17703 VDD.n2574 VDD.n2573 185
R17704 VDD.n2573 VDD.n2572 185
R17705 VDD.n915 VDD.n914 185
R17706 VDD.n916 VDD.n915 185
R17707 VDD.n2565 VDD.n2564 185
R17708 VDD.n2566 VDD.n2565 185
R17709 VDD.n2563 VDD.n925 185
R17710 VDD.n925 VDD.n922 185
R17711 VDD.n2562 VDD.n2561 185
R17712 VDD.n2561 VDD.n2560 185
R17713 VDD.n927 VDD.n926 185
R17714 VDD.n928 VDD.n927 185
R17715 VDD.n2553 VDD.n2552 185
R17716 VDD.n2554 VDD.n2553 185
R17717 VDD.n2551 VDD.n937 185
R17718 VDD.n937 VDD.n934 185
R17719 VDD.n2550 VDD.n2549 185
R17720 VDD.n2549 VDD.n2548 185
R17721 VDD.n939 VDD.n938 185
R17722 VDD.n948 VDD.n939 185
R17723 VDD.n2541 VDD.n2540 185
R17724 VDD.n2542 VDD.n2541 185
R17725 VDD.n2539 VDD.n949 185
R17726 VDD.n949 VDD.n945 185
R17727 VDD.n2538 VDD.n2537 185
R17728 VDD.n2537 VDD.n2536 185
R17729 VDD.n951 VDD.n950 185
R17730 VDD.n952 VDD.n951 185
R17731 VDD.n2529 VDD.n2528 185
R17732 VDD.n2530 VDD.n2529 185
R17733 VDD.n2527 VDD.n961 185
R17734 VDD.n961 VDD.n958 185
R17735 VDD.n2526 VDD.n2525 185
R17736 VDD.n2525 VDD.n2524 185
R17737 VDD.n963 VDD.n962 185
R17738 VDD.n964 VDD.n963 185
R17739 VDD.n2517 VDD.n2516 185
R17740 VDD.n2518 VDD.n2517 185
R17741 VDD.n2515 VDD.n973 185
R17742 VDD.n973 VDD.n970 185
R17743 VDD.n2514 VDD.n2513 185
R17744 VDD.n2513 VDD.n2512 185
R17745 VDD.n975 VDD.n974 185
R17746 VDD.n976 VDD.n975 185
R17747 VDD.n2505 VDD.n2504 185
R17748 VDD.n2506 VDD.n2505 185
R17749 VDD.n2503 VDD.n985 185
R17750 VDD.n985 VDD.n982 185
R17751 VDD.n2502 VDD.n2501 185
R17752 VDD.n2501 VDD.n2500 185
R17753 VDD.n987 VDD.n986 185
R17754 VDD.n988 VDD.n987 185
R17755 VDD.n2493 VDD.n2492 185
R17756 VDD.n2494 VDD.n2493 185
R17757 VDD.n2491 VDD.n997 185
R17758 VDD.n997 VDD.n994 185
R17759 VDD.n2490 VDD.n2489 185
R17760 VDD.n2489 VDD.n2488 185
R17761 VDD.n999 VDD.n998 185
R17762 VDD.n1000 VDD.n999 185
R17763 VDD.n2481 VDD.n2480 185
R17764 VDD.n2482 VDD.n2481 185
R17765 VDD.n2479 VDD.n1009 185
R17766 VDD.n1009 VDD.n1006 185
R17767 VDD.n2478 VDD.n2477 185
R17768 VDD.n2477 VDD.n2476 185
R17769 VDD.n1011 VDD.n1010 185
R17770 VDD.n1012 VDD.n1011 185
R17771 VDD.n2469 VDD.n2468 185
R17772 VDD.n2470 VDD.n2469 185
R17773 VDD.n2467 VDD.n1020 185
R17774 VDD.n1026 VDD.n1020 185
R17775 VDD.n2466 VDD.n2465 185
R17776 VDD.n2465 VDD.n2464 185
R17777 VDD.n1022 VDD.n1021 185
R17778 VDD.n1023 VDD.n1022 185
R17779 VDD.n2457 VDD.n2456 185
R17780 VDD.n2458 VDD.n2457 185
R17781 VDD.n2455 VDD.n1033 185
R17782 VDD.n1033 VDD.n1030 185
R17783 VDD.n2454 VDD.n2453 185
R17784 VDD.n2453 VDD.n2452 185
R17785 VDD.n1035 VDD.n1034 185
R17786 VDD.n1036 VDD.n1035 185
R17787 VDD.n2445 VDD.n2444 185
R17788 VDD.n2446 VDD.n2445 185
R17789 VDD.n2443 VDD.n1045 185
R17790 VDD.n1045 VDD.n1042 185
R17791 VDD.n2442 VDD.n2441 185
R17792 VDD.n2441 VDD.n2440 185
R17793 VDD.n1047 VDD.n1046 185
R17794 VDD.n1048 VDD.n1047 185
R17795 VDD.n2433 VDD.n2432 185
R17796 VDD.n2434 VDD.n2433 185
R17797 VDD.n2431 VDD.n1057 185
R17798 VDD.n1057 VDD.n1054 185
R17799 VDD.n2430 VDD.n2429 185
R17800 VDD.n2429 VDD.n2428 185
R17801 VDD.n1059 VDD.n1058 185
R17802 VDD.n1060 VDD.n1059 185
R17803 VDD.n2421 VDD.n2420 185
R17804 VDD.n2422 VDD.n2421 185
R17805 VDD.n2419 VDD.n1068 185
R17806 VDD.n1074 VDD.n1068 185
R17807 VDD.n2418 VDD.n2417 185
R17808 VDD.n2417 VDD.n2416 185
R17809 VDD.n1070 VDD.n1069 185
R17810 VDD.n1071 VDD.n1070 185
R17811 VDD.n2409 VDD.n2408 185
R17812 VDD.n2410 VDD.n2409 185
R17813 VDD.n2407 VDD.n1081 185
R17814 VDD.n1081 VDD.n1078 185
R17815 VDD.n2406 VDD.n2405 185
R17816 VDD.n2405 VDD.n2404 185
R17817 VDD.n1083 VDD.n1082 185
R17818 VDD.n1084 VDD.n1083 185
R17819 VDD.n2397 VDD.n2396 185
R17820 VDD.n2398 VDD.n2397 185
R17821 VDD.n2395 VDD.n1093 185
R17822 VDD.n1093 VDD.n1090 185
R17823 VDD.n2394 VDD.n2393 185
R17824 VDD.n2393 VDD.n2392 185
R17825 VDD.n1095 VDD.n1094 185
R17826 VDD.n1096 VDD.n1095 185
R17827 VDD.n2385 VDD.n2384 185
R17828 VDD.n2386 VDD.n2385 185
R17829 VDD.n2867 VDD.n658 185
R17830 VDD.n2902 VDD.n658 185
R17831 VDD.n2869 VDD.n2868 185
R17832 VDD.n2871 VDD.n2870 185
R17833 VDD.n2873 VDD.n2872 185
R17834 VDD.n2876 VDD.n2875 185
R17835 VDD.n2878 VDD.n2877 185
R17836 VDD.n2880 VDD.n2879 185
R17837 VDD.n2882 VDD.n2881 185
R17838 VDD.n2884 VDD.n2883 185
R17839 VDD.n2886 VDD.n2885 185
R17840 VDD.n2888 VDD.n2887 185
R17841 VDD.n2890 VDD.n2889 185
R17842 VDD.n2892 VDD.n2891 185
R17843 VDD.n2894 VDD.n2893 185
R17844 VDD.n2896 VDD.n2895 185
R17845 VDD.n2898 VDD.n2897 185
R17846 VDD.n2899 VDD.n660 185
R17847 VDD.n2901 VDD.n2900 185
R17848 VDD.n2902 VDD.n2901 185
R17849 VDD.n2866 VDD.n2865 185
R17850 VDD.n2865 VDD.n640 185
R17851 VDD.n2864 VDD.n664 185
R17852 VDD.n2864 VDD.n2863 185
R17853 VDD.n1118 VDD.n665 185
R17854 VDD.n666 VDD.n665 185
R17855 VDD.n1119 VDD.n678 185
R17856 VDD.n2817 VDD.n678 185
R17857 VDD.n1121 VDD.n1120 185
R17858 VDD.n1120 VDD.n677 185
R17859 VDD.n1122 VDD.n685 185
R17860 VDD.n2811 VDD.n685 185
R17861 VDD.n1124 VDD.n1123 185
R17862 VDD.n1123 VDD.n683 185
R17863 VDD.n1125 VDD.n692 185
R17864 VDD.n2800 VDD.n692 185
R17865 VDD.n1127 VDD.n1126 185
R17866 VDD.n1126 VDD.n690 185
R17867 VDD.n1128 VDD.n698 185
R17868 VDD.n2794 VDD.n698 185
R17869 VDD.n1130 VDD.n1129 185
R17870 VDD.n1129 VDD.n696 185
R17871 VDD.n1131 VDD.n703 185
R17872 VDD.n2788 VDD.n703 185
R17873 VDD.n2149 VDD.n2148 185
R17874 VDD.n2148 VDD.n2147 185
R17875 VDD.n2150 VDD.n709 185
R17876 VDD.n2782 VDD.n709 185
R17877 VDD.n2152 VDD.n2151 185
R17878 VDD.n2151 VDD.n707 185
R17879 VDD.n2153 VDD.n715 185
R17880 VDD.n2776 VDD.n715 185
R17881 VDD.n2155 VDD.n2154 185
R17882 VDD.n2154 VDD.n713 185
R17883 VDD.n2156 VDD.n721 185
R17884 VDD.n2770 VDD.n721 185
R17885 VDD.n2158 VDD.n2157 185
R17886 VDD.n2157 VDD.n719 185
R17887 VDD.n2159 VDD.n727 185
R17888 VDD.n2764 VDD.n727 185
R17889 VDD.n2161 VDD.n2160 185
R17890 VDD.n2160 VDD.n725 185
R17891 VDD.n2162 VDD.n733 185
R17892 VDD.n2758 VDD.n733 185
R17893 VDD.n2164 VDD.n2163 185
R17894 VDD.n2163 VDD.n731 185
R17895 VDD.n2165 VDD.n739 185
R17896 VDD.n2752 VDD.n739 185
R17897 VDD.n2167 VDD.n2166 185
R17898 VDD.n2166 VDD.n737 185
R17899 VDD.n2168 VDD.n745 185
R17900 VDD.n2746 VDD.n745 185
R17901 VDD.n2170 VDD.n2169 185
R17902 VDD.n2169 VDD.n743 185
R17903 VDD.n2171 VDD.n751 185
R17904 VDD.n2740 VDD.n751 185
R17905 VDD.n2173 VDD.n2172 185
R17906 VDD.n2172 VDD.n749 185
R17907 VDD.n2174 VDD.n757 185
R17908 VDD.n2734 VDD.n757 185
R17909 VDD.n2176 VDD.n2175 185
R17910 VDD.n2175 VDD.n755 185
R17911 VDD.n2177 VDD.n762 185
R17912 VDD.n2728 VDD.n762 185
R17913 VDD.n2179 VDD.n2178 185
R17914 VDD.n2178 VDD.n769 185
R17915 VDD.n2180 VDD.n768 185
R17916 VDD.n2722 VDD.n768 185
R17917 VDD.n2182 VDD.n2181 185
R17918 VDD.n2181 VDD.n766 185
R17919 VDD.n2183 VDD.n775 185
R17920 VDD.n2716 VDD.n775 185
R17921 VDD.n2185 VDD.n2184 185
R17922 VDD.n2184 VDD.n773 185
R17923 VDD.n2186 VDD.n781 185
R17924 VDD.n2710 VDD.n781 185
R17925 VDD.n2188 VDD.n2187 185
R17926 VDD.n2187 VDD.n779 185
R17927 VDD.n2189 VDD.n787 185
R17928 VDD.n2704 VDD.n787 185
R17929 VDD.n2191 VDD.n2190 185
R17930 VDD.n2190 VDD.n785 185
R17931 VDD.n2192 VDD.n793 185
R17932 VDD.n2698 VDD.n793 185
R17933 VDD.n2194 VDD.n2193 185
R17934 VDD.n2193 VDD.n791 185
R17935 VDD.n2195 VDD.n799 185
R17936 VDD.n2692 VDD.n799 185
R17937 VDD.n2197 VDD.n2196 185
R17938 VDD.n2196 VDD.n797 185
R17939 VDD.n2198 VDD.n805 185
R17940 VDD.n2686 VDD.n805 185
R17941 VDD.n2200 VDD.n2199 185
R17942 VDD.n2199 VDD.n803 185
R17943 VDD.n2201 VDD.n811 185
R17944 VDD.n2680 VDD.n811 185
R17945 VDD.n2203 VDD.n2202 185
R17946 VDD.n2202 VDD.n809 185
R17947 VDD.n2204 VDD.n817 185
R17948 VDD.n2674 VDD.n817 185
R17949 VDD.n2206 VDD.n2205 185
R17950 VDD.n2205 VDD.n815 185
R17951 VDD.n2207 VDD.n823 185
R17952 VDD.n2668 VDD.n823 185
R17953 VDD.n2209 VDD.n2208 185
R17954 VDD.n2208 VDD.n821 185
R17955 VDD.n2210 VDD.n828 185
R17956 VDD.n2662 VDD.n828 185
R17957 VDD.n2212 VDD.n2211 185
R17958 VDD.n2211 VDD.n835 185
R17959 VDD.n2213 VDD.n834 185
R17960 VDD.n2656 VDD.n834 185
R17961 VDD.n2215 VDD.n2214 185
R17962 VDD.n2214 VDD.n832 185
R17963 VDD.n2216 VDD.n841 185
R17964 VDD.n2650 VDD.n841 185
R17965 VDD.n2218 VDD.n2217 185
R17966 VDD.n2217 VDD.n839 185
R17967 VDD.n2219 VDD.n847 185
R17968 VDD.n2644 VDD.n847 185
R17969 VDD.n2221 VDD.n2220 185
R17970 VDD.n2220 VDD.n845 185
R17971 VDD.n2222 VDD.n853 185
R17972 VDD.n2638 VDD.n853 185
R17973 VDD.n2224 VDD.n2223 185
R17974 VDD.n2223 VDD.n851 185
R17975 VDD.n2225 VDD.n859 185
R17976 VDD.n2632 VDD.n859 185
R17977 VDD.n2227 VDD.n2226 185
R17978 VDD.n2226 VDD.n857 185
R17979 VDD.n2228 VDD.n865 185
R17980 VDD.n2626 VDD.n865 185
R17981 VDD.n2230 VDD.n2229 185
R17982 VDD.n2229 VDD.n863 185
R17983 VDD.n2231 VDD.n871 185
R17984 VDD.n2620 VDD.n871 185
R17985 VDD.n2233 VDD.n2232 185
R17986 VDD.n2232 VDD.n869 185
R17987 VDD.n2234 VDD.n876 185
R17988 VDD.n2614 VDD.n876 185
R17989 VDD.n2236 VDD.n2235 185
R17990 VDD.n2235 VDD.t92 185
R17991 VDD.n2237 VDD.n882 185
R17992 VDD.n2608 VDD.n882 185
R17993 VDD.n2239 VDD.n2238 185
R17994 VDD.n2238 VDD.n880 185
R17995 VDD.n2240 VDD.n888 185
R17996 VDD.n2602 VDD.n888 185
R17997 VDD.n2242 VDD.n2241 185
R17998 VDD.n2241 VDD.n886 185
R17999 VDD.n2243 VDD.n894 185
R18000 VDD.n2596 VDD.n894 185
R18001 VDD.n2245 VDD.n2244 185
R18002 VDD.n2244 VDD.n892 185
R18003 VDD.n2246 VDD.n900 185
R18004 VDD.n2590 VDD.n900 185
R18005 VDD.n2248 VDD.n2247 185
R18006 VDD.n2247 VDD.n898 185
R18007 VDD.n2249 VDD.n906 185
R18008 VDD.n2584 VDD.n906 185
R18009 VDD.n2251 VDD.n2250 185
R18010 VDD.n2250 VDD.n904 185
R18011 VDD.n2252 VDD.n912 185
R18012 VDD.n2578 VDD.n912 185
R18013 VDD.n2254 VDD.n2253 185
R18014 VDD.n2253 VDD.n910 185
R18015 VDD.n2255 VDD.n918 185
R18016 VDD.n2572 VDD.n918 185
R18017 VDD.n2257 VDD.n2256 185
R18018 VDD.n2256 VDD.n916 185
R18019 VDD.n2258 VDD.n924 185
R18020 VDD.n2566 VDD.n924 185
R18021 VDD.n2260 VDD.n2259 185
R18022 VDD.n2259 VDD.n922 185
R18023 VDD.n2261 VDD.n930 185
R18024 VDD.n2560 VDD.n930 185
R18025 VDD.n2263 VDD.n2262 185
R18026 VDD.n2262 VDD.n928 185
R18027 VDD.n2264 VDD.n936 185
R18028 VDD.n2554 VDD.n936 185
R18029 VDD.n2266 VDD.n2265 185
R18030 VDD.n2265 VDD.n934 185
R18031 VDD.n2267 VDD.n941 185
R18032 VDD.n2548 VDD.n941 185
R18033 VDD.n2269 VDD.n2268 185
R18034 VDD.n2268 VDD.n948 185
R18035 VDD.n2270 VDD.n947 185
R18036 VDD.n2542 VDD.n947 185
R18037 VDD.n2272 VDD.n2271 185
R18038 VDD.n2271 VDD.n945 185
R18039 VDD.n2273 VDD.n954 185
R18040 VDD.n2536 VDD.n954 185
R18041 VDD.n2275 VDD.n2274 185
R18042 VDD.n2274 VDD.n952 185
R18043 VDD.n2276 VDD.n960 185
R18044 VDD.n2530 VDD.n960 185
R18045 VDD.n2278 VDD.n2277 185
R18046 VDD.n2277 VDD.n958 185
R18047 VDD.n2279 VDD.n966 185
R18048 VDD.n2524 VDD.n966 185
R18049 VDD.n2281 VDD.n2280 185
R18050 VDD.n2280 VDD.n964 185
R18051 VDD.n2282 VDD.n972 185
R18052 VDD.n2518 VDD.n972 185
R18053 VDD.n2284 VDD.n2283 185
R18054 VDD.n2283 VDD.n970 185
R18055 VDD.n2285 VDD.n978 185
R18056 VDD.n2512 VDD.n978 185
R18057 VDD.n2287 VDD.n2286 185
R18058 VDD.n2286 VDD.n976 185
R18059 VDD.n2288 VDD.n984 185
R18060 VDD.n2506 VDD.n984 185
R18061 VDD.n2290 VDD.n2289 185
R18062 VDD.n2289 VDD.n982 185
R18063 VDD.n2291 VDD.n990 185
R18064 VDD.n2500 VDD.n990 185
R18065 VDD.n2293 VDD.n2292 185
R18066 VDD.n2292 VDD.n988 185
R18067 VDD.n2294 VDD.n996 185
R18068 VDD.n2494 VDD.n996 185
R18069 VDD.n2296 VDD.n2295 185
R18070 VDD.n2295 VDD.n994 185
R18071 VDD.n2297 VDD.n1002 185
R18072 VDD.n2488 VDD.n1002 185
R18073 VDD.n2299 VDD.n2298 185
R18074 VDD.n2298 VDD.n1000 185
R18075 VDD.n2300 VDD.n1008 185
R18076 VDD.n2482 VDD.n1008 185
R18077 VDD.n2302 VDD.n2301 185
R18078 VDD.n2301 VDD.n1006 185
R18079 VDD.n2303 VDD.n1014 185
R18080 VDD.n2476 VDD.n1014 185
R18081 VDD.n2305 VDD.n2304 185
R18082 VDD.n2304 VDD.n1012 185
R18083 VDD.n2306 VDD.n1019 185
R18084 VDD.n2470 VDD.n1019 185
R18085 VDD.n2308 VDD.n2307 185
R18086 VDD.n2307 VDD.n1026 185
R18087 VDD.n2309 VDD.n1025 185
R18088 VDD.n2464 VDD.n1025 185
R18089 VDD.n2311 VDD.n2310 185
R18090 VDD.n2310 VDD.n1023 185
R18091 VDD.n2312 VDD.n1032 185
R18092 VDD.n2458 VDD.n1032 185
R18093 VDD.n2314 VDD.n2313 185
R18094 VDD.n2313 VDD.n1030 185
R18095 VDD.n2315 VDD.n1038 185
R18096 VDD.n2452 VDD.n1038 185
R18097 VDD.n2317 VDD.n2316 185
R18098 VDD.n2316 VDD.n1036 185
R18099 VDD.n2318 VDD.n1044 185
R18100 VDD.n2446 VDD.n1044 185
R18101 VDD.n2320 VDD.n2319 185
R18102 VDD.n2319 VDD.n1042 185
R18103 VDD.n2321 VDD.n1050 185
R18104 VDD.n2440 VDD.n1050 185
R18105 VDD.n2323 VDD.n2322 185
R18106 VDD.n2322 VDD.n1048 185
R18107 VDD.n2324 VDD.n1056 185
R18108 VDD.n2434 VDD.n1056 185
R18109 VDD.n2326 VDD.n2325 185
R18110 VDD.n2325 VDD.n1054 185
R18111 VDD.n2327 VDD.n1062 185
R18112 VDD.n2428 VDD.n1062 185
R18113 VDD.n2329 VDD.n2328 185
R18114 VDD.n2328 VDD.n1060 185
R18115 VDD.n2330 VDD.n1067 185
R18116 VDD.n2422 VDD.n1067 185
R18117 VDD.n2332 VDD.n2331 185
R18118 VDD.n2331 VDD.n1074 185
R18119 VDD.n2333 VDD.n1073 185
R18120 VDD.n2416 VDD.n1073 185
R18121 VDD.n2335 VDD.n2334 185
R18122 VDD.n2334 VDD.n1071 185
R18123 VDD.n2336 VDD.n1080 185
R18124 VDD.n2410 VDD.n1080 185
R18125 VDD.n2338 VDD.n2337 185
R18126 VDD.n2337 VDD.n1078 185
R18127 VDD.n2339 VDD.n1086 185
R18128 VDD.n2404 VDD.n1086 185
R18129 VDD.n2341 VDD.n2340 185
R18130 VDD.n2340 VDD.n1084 185
R18131 VDD.n2342 VDD.n1092 185
R18132 VDD.n2398 VDD.n1092 185
R18133 VDD.n2344 VDD.n2343 185
R18134 VDD.n2343 VDD.n1090 185
R18135 VDD.n2345 VDD.n1098 185
R18136 VDD.n2392 VDD.n1098 185
R18137 VDD.n2347 VDD.n2346 185
R18138 VDD.n2346 VDD.n1096 185
R18139 VDD.n2348 VDD.n1104 185
R18140 VDD.n2386 VDD.n1104 185
R18141 VDD.n2383 VDD.n1105 185
R18142 VDD.n1105 VDD.n1102 185
R18143 VDD.n2382 VDD.n2381 185
R18144 VDD.n2379 VDD.n1106 185
R18145 VDD.n2378 VDD.n2377 185
R18146 VDD.n2376 VDD.n2375 185
R18147 VDD.n2374 VDD.n1108 185
R18148 VDD.n2372 VDD.n2371 185
R18149 VDD.n2370 VDD.n1109 185
R18150 VDD.n2369 VDD.n2368 185
R18151 VDD.n2366 VDD.n2365 185
R18152 VDD.n2364 VDD.n2363 185
R18153 VDD.n2362 VDD.n1112 185
R18154 VDD.n2360 VDD.n2359 185
R18155 VDD.n2358 VDD.n1113 185
R18156 VDD.n2356 VDD.n2355 185
R18157 VDD.n2353 VDD.n1116 185
R18158 VDD.n2351 VDD.n2350 185
R18159 VDD.n2349 VDD.n1117 185
R18160 VDD.n1117 VDD.n1102 185
R18161 VDD.n1295 VDD.t142 161.415
R18162 VDD.n1298 VDD.t144 160.572
R18163 VDD.n1297 VDD.t143 160.572
R18164 VDD.n1296 VDD.t141 160.572
R18165 VDD.n1295 VDD.t136 160.572
R18166 VDD.n16 VDD.t145 160.47
R18167 VDD.n19 VDD.t139 159.627
R18168 VDD.n18 VDD.t138 159.627
R18169 VDD.n17 VDD.t146 159.627
R18170 VDD.n16 VDD.t140 159.627
R18171 VDD.n9 VDD.n7 150.946
R18172 VDD.n2 VDD.n0 150.946
R18173 VDD.n1377 VDD.t5 149.125
R18174 VDD.n1391 VDD.t57 149.125
R18175 VDD.n1408 VDD.t2 149.125
R18176 VDD.n1422 VDD.t8 149.125
R18177 VDD.n1439 VDD.t15 149.125
R18178 VDD.n1143 VDD.t91 149.125
R18179 VDD.n1226 VDD.t35 149.125
R18180 VDD.n1203 VDD.t76 149.125
R18181 VDD.n1183 VDD.t73 149.125
R18182 VDD.n1162 VDD.t85 149.125
R18183 VDD.n4364 VDD.t45 149.125
R18184 VDD.n4343 VDD.t88 149.125
R18185 VDD.n4323 VDD.t55 149.125
R18186 VDD.n4302 VDD.t61 149.125
R18187 VDD.n4279 VDD.t67 149.125
R18188 VDD.n138 VDD.t47 149.125
R18189 VDD.n160 VDD.t26 149.125
R18190 VDD.n3945 VDD.t12 149.125
R18191 VDD.n4034 VDD.t37 149.125
R18192 VDD.n3965 VDD.t63 149.125
R18193 VDD.n9 VDD.n8 149.084
R18194 VDD.n11 VDD.n10 149.084
R18195 VDD.n13 VDD.n12 149.084
R18196 VDD.n6 VDD.n5 149.084
R18197 VDD.n4 VDD.n3 149.084
R18198 VDD.n2 VDD.n1 149.084
R18199 VDD.n1115 VDD.t23 149.028
R18200 VDD.n663 VDD.t31 149.028
R18201 VDD.n1135 VDD.t81 149.028
R18202 VDD.n673 VDD.t41 149.028
R18203 VDD.n3118 VDD.t78 149.028
R18204 VDD.n202 VDD.t70 149.028
R18205 VDD.n2922 VDD.t51 149.028
R18206 VDD.n178 VDD.t20 149.028
R18207 VDD.n4082 VDD.n95 146.341
R18208 VDD.n4082 VDD.n87 146.341
R18209 VDD.n4092 VDD.n87 146.341
R18210 VDD.n4092 VDD.n83 146.341
R18211 VDD.n4098 VDD.n83 146.341
R18212 VDD.n4098 VDD.n75 146.341
R18213 VDD.n4107 VDD.n75 146.341
R18214 VDD.n4107 VDD.n71 146.341
R18215 VDD.n4113 VDD.n71 146.341
R18216 VDD.n4113 VDD.n63 146.341
R18217 VDD.n4123 VDD.n63 146.341
R18218 VDD.n4123 VDD.n59 146.341
R18219 VDD.n4129 VDD.n59 146.341
R18220 VDD.n4129 VDD.n51 146.341
R18221 VDD.n4139 VDD.n51 146.341
R18222 VDD.n4139 VDD.n47 146.341
R18223 VDD.n4145 VDD.n47 146.341
R18224 VDD.n4145 VDD.n39 146.341
R18225 VDD.n4155 VDD.n39 146.341
R18226 VDD.n4155 VDD.n35 146.341
R18227 VDD.n4161 VDD.n35 146.341
R18228 VDD.n4161 VDD.n24 146.341
R18229 VDD.n4540 VDD.n24 146.341
R18230 VDD.n4540 VDD.n25 146.341
R18231 VDD.n4533 VDD.n25 146.341
R18232 VDD.n4533 VDD.n4173 146.341
R18233 VDD.n4529 VDD.n4173 146.341
R18234 VDD.n4529 VDD.n4178 146.341
R18235 VDD.n4525 VDD.n4178 146.341
R18236 VDD.n4525 VDD.n4183 146.341
R18237 VDD.n4521 VDD.n4183 146.341
R18238 VDD.n4521 VDD.n4189 146.341
R18239 VDD.n4517 VDD.n4189 146.341
R18240 VDD.n4517 VDD.n4194 146.341
R18241 VDD.n4513 VDD.n4194 146.341
R18242 VDD.n4513 VDD.n4200 146.341
R18243 VDD.n4509 VDD.n4200 146.341
R18244 VDD.n4509 VDD.n4205 146.341
R18245 VDD.n4505 VDD.n4205 146.341
R18246 VDD.n4505 VDD.n4211 146.341
R18247 VDD.n4498 VDD.n4211 146.341
R18248 VDD.n4498 VDD.n4248 146.341
R18249 VDD.n4494 VDD.n4248 146.341
R18250 VDD.n4494 VDD.n4254 146.341
R18251 VDD.n4490 VDD.n4254 146.341
R18252 VDD.n4490 VDD.n4259 146.341
R18253 VDD.n4482 VDD.n4481 146.341
R18254 VDD.n4479 VDD.n4266 146.341
R18255 VDD.n4475 VDD.n4474 146.341
R18256 VDD.n4472 VDD.n4273 146.341
R18257 VDD.n4284 VDD.n4281 146.341
R18258 VDD.n4464 VDD.n4463 146.341
R18259 VDD.n4461 VDD.n4286 146.341
R18260 VDD.n4457 VDD.n4456 146.341
R18261 VDD.n4454 VDD.n4292 146.341
R18262 VDD.n4450 VDD.n4449 146.341
R18263 VDD.n4447 VDD.n4299 146.341
R18264 VDD.n4441 VDD.n4440 146.341
R18265 VDD.n4438 VDD.n4307 146.341
R18266 VDD.n4434 VDD.n4433 146.341
R18267 VDD.n4431 VDD.n4313 146.341
R18268 VDD.n4427 VDD.n4426 146.341
R18269 VDD.n4424 VDD.n4320 146.341
R18270 VDD.n4418 VDD.n4417 146.341
R18271 VDD.n4415 VDD.n4328 146.341
R18272 VDD.n4411 VDD.n4410 146.341
R18273 VDD.n4408 VDD.n4334 146.341
R18274 VDD.n4404 VDD.n4403 146.341
R18275 VDD.n4401 VDD.n4341 146.341
R18276 VDD.n4397 VDD.n4396 146.341
R18277 VDD.n4394 VDD.n4351 146.341
R18278 VDD.n4390 VDD.n4389 146.341
R18279 VDD.n4387 VDD.n4358 146.341
R18280 VDD.n4383 VDD.n4382 146.341
R18281 VDD.n4084 VDD.n93 146.341
R18282 VDD.n4084 VDD.n89 146.341
R18283 VDD.n4090 VDD.n89 146.341
R18284 VDD.n4090 VDD.n81 146.341
R18285 VDD.n4100 VDD.n81 146.341
R18286 VDD.n4100 VDD.n77 146.341
R18287 VDD.n4106 VDD.n77 146.341
R18288 VDD.n4106 VDD.n69 146.341
R18289 VDD.n4115 VDD.n69 146.341
R18290 VDD.n4115 VDD.n65 146.341
R18291 VDD.n4121 VDD.n65 146.341
R18292 VDD.n4121 VDD.n57 146.341
R18293 VDD.n4131 VDD.n57 146.341
R18294 VDD.n4131 VDD.n53 146.341
R18295 VDD.n4137 VDD.n53 146.341
R18296 VDD.n4137 VDD.n45 146.341
R18297 VDD.n4147 VDD.n45 146.341
R18298 VDD.n4147 VDD.n41 146.341
R18299 VDD.n4153 VDD.n41 146.341
R18300 VDD.n4153 VDD.n33 146.341
R18301 VDD.n4163 VDD.n33 146.341
R18302 VDD.n4163 VDD.n28 146.341
R18303 VDD.n4539 VDD.n28 146.341
R18304 VDD.n4539 VDD.n29 146.341
R18305 VDD.n4535 VDD.n29 146.341
R18306 VDD.n4535 VDD.n4171 146.341
R18307 VDD.n4179 VDD.n4171 146.341
R18308 VDD.n4180 VDD.n4179 146.341
R18309 VDD.n4181 VDD.n4180 146.341
R18310 VDD.n4220 VDD.n4181 146.341
R18311 VDD.n4220 VDD.n4190 146.341
R18312 VDD.n4191 VDD.n4190 146.341
R18313 VDD.n4192 VDD.n4191 146.341
R18314 VDD.n4217 VDD.n4192 146.341
R18315 VDD.n4217 VDD.n4201 146.341
R18316 VDD.n4202 VDD.n4201 146.341
R18317 VDD.n4203 VDD.n4202 146.341
R18318 VDD.n4213 VDD.n4203 146.341
R18319 VDD.n4504 VDD.n4213 146.341
R18320 VDD.n4504 VDD.n4214 146.341
R18321 VDD.n4500 VDD.n4214 146.341
R18322 VDD.n4500 VDD.n4246 146.341
R18323 VDD.n4255 VDD.n4246 146.341
R18324 VDD.n4256 VDD.n4255 146.341
R18325 VDD.n4257 VDD.n4256 146.341
R18326 VDD.n4367 VDD.n4257 146.341
R18327 VDD.n4073 VDD.n99 146.341
R18328 VDD.n4073 VDD.n128 146.341
R18329 VDD.n4069 VDD.n4068 146.341
R18330 VDD.n4065 VDD.n4064 146.341
R18331 VDD.n4061 VDD.n4060 146.341
R18332 VDD.n4057 VDD.n4056 146.341
R18333 VDD.n4053 VDD.n4052 146.341
R18334 VDD.n4049 VDD.n4048 146.341
R18335 VDD.n4045 VDD.n4044 146.341
R18336 VDD.n4041 VDD.n4040 146.341
R18337 VDD.n4037 VDD.n4036 146.341
R18338 VDD.n4028 VDD.n4027 146.341
R18339 VDD.n4025 VDD.n4024 146.341
R18340 VDD.n4021 VDD.n4020 146.341
R18341 VDD.n4017 VDD.n4016 146.341
R18342 VDD.n4013 VDD.n4012 146.341
R18343 VDD.n4009 VDD.n4008 146.341
R18344 VDD.n4005 VDD.n4004 146.341
R18345 VDD.n4001 VDD.n4000 146.341
R18346 VDD.n3997 VDD.n3996 146.341
R18347 VDD.n3993 VDD.n3992 146.341
R18348 VDD.n3989 VDD.n3988 146.341
R18349 VDD.n3948 VDD.n3947 146.341
R18350 VDD.n3952 VDD.n3951 146.341
R18351 VDD.n3981 VDD.n3980 146.341
R18352 VDD.n3977 VDD.n3976 146.341
R18353 VDD.n3973 VDD.n3972 146.341
R18354 VDD.n3969 VDD.n3968 146.341
R18355 VDD.n3961 VDD.n127 146.341
R18356 VDD.n1796 VDD.n1772 146.341
R18357 VDD.n1794 VDD.n1793 146.341
R18358 VDD.n1791 VDD.n1776 146.341
R18359 VDD.n1787 VDD.n1786 146.341
R18360 VDD.n1891 VDD.n1145 146.341
R18361 VDD.n1889 VDD.n1888 146.341
R18362 VDD.n1886 VDD.n1148 146.341
R18363 VDD.n1882 VDD.n1881 146.341
R18364 VDD.n1879 VDD.n1152 146.341
R18365 VDD.n1875 VDD.n1874 146.341
R18366 VDD.n1872 VDD.n1159 146.341
R18367 VDD.n1866 VDD.n1865 146.341
R18368 VDD.n1863 VDD.n1167 146.341
R18369 VDD.n1859 VDD.n1858 146.341
R18370 VDD.n1856 VDD.n1173 146.341
R18371 VDD.n1852 VDD.n1851 146.341
R18372 VDD.n1849 VDD.n1180 146.341
R18373 VDD.n1843 VDD.n1842 146.341
R18374 VDD.n1840 VDD.n1188 146.341
R18375 VDD.n1836 VDD.n1835 146.341
R18376 VDD.n1833 VDD.n1194 146.341
R18377 VDD.n1829 VDD.n1828 146.341
R18378 VDD.n1826 VDD.n1201 146.341
R18379 VDD.n1210 VDD.n1209 146.341
R18380 VDD.n1213 VDD.n1212 146.341
R18381 VDD.n1218 VDD.n1217 146.341
R18382 VDD.n1221 VDD.n1220 146.341
R18383 VDD.n1808 VDD.n1228 146.341
R18384 VDD.n1586 VDD.n1366 146.341
R18385 VDD.n1596 VDD.n1366 146.341
R18386 VDD.n1596 VDD.n1362 146.341
R18387 VDD.n1602 VDD.n1362 146.341
R18388 VDD.n1602 VDD.n1354 146.341
R18389 VDD.n1612 VDD.n1354 146.341
R18390 VDD.n1612 VDD.n1350 146.341
R18391 VDD.n1618 VDD.n1350 146.341
R18392 VDD.n1618 VDD.n1343 146.341
R18393 VDD.n1628 VDD.n1343 146.341
R18394 VDD.n1628 VDD.n1339 146.341
R18395 VDD.n1634 VDD.n1339 146.341
R18396 VDD.n1634 VDD.n1331 146.341
R18397 VDD.n1644 VDD.n1331 146.341
R18398 VDD.n1644 VDD.n1327 146.341
R18399 VDD.n1650 VDD.n1327 146.341
R18400 VDD.n1650 VDD.n1319 146.341
R18401 VDD.n1660 VDD.n1319 146.341
R18402 VDD.n1660 VDD.n1315 146.341
R18403 VDD.n1666 VDD.n1315 146.341
R18404 VDD.n1666 VDD.n1307 146.341
R18405 VDD.n1676 VDD.n1307 146.341
R18406 VDD.n1676 VDD.n1303 146.341
R18407 VDD.n1682 VDD.n1303 146.341
R18408 VDD.n1682 VDD.n1291 146.341
R18409 VDD.n1692 VDD.n1291 146.341
R18410 VDD.n1692 VDD.n1287 146.341
R18411 VDD.n1698 VDD.n1287 146.341
R18412 VDD.n1698 VDD.n1279 146.341
R18413 VDD.n1708 VDD.n1279 146.341
R18414 VDD.n1708 VDD.n1275 146.341
R18415 VDD.n1714 VDD.n1275 146.341
R18416 VDD.n1714 VDD.n1267 146.341
R18417 VDD.n1724 VDD.n1267 146.341
R18418 VDD.n1724 VDD.n1263 146.341
R18419 VDD.n1730 VDD.n1263 146.341
R18420 VDD.n1730 VDD.n1255 146.341
R18421 VDD.n1740 VDD.n1255 146.341
R18422 VDD.n1740 VDD.n1251 146.341
R18423 VDD.n1746 VDD.n1251 146.341
R18424 VDD.n1746 VDD.n1244 146.341
R18425 VDD.n1756 VDD.n1244 146.341
R18426 VDD.n1756 VDD.n1239 146.341
R18427 VDD.n1764 VDD.n1239 146.341
R18428 VDD.n1764 VDD.n1229 146.341
R18429 VDD.n1805 VDD.n1229 146.341
R18430 VDD.n1451 VDD.n1450 146.341
R18431 VDD.n1453 VDD.n1451 146.341
R18432 VDD.n1461 VDD.n1442 146.341
R18433 VDD.n1464 VDD.n1463 146.341
R18434 VDD.n1466 VDD.n1437 146.341
R18435 VDD.n1473 VDD.n1433 146.341
R18436 VDD.n1477 VDD.n1475 146.341
R18437 VDD.n1484 VDD.n1429 146.341
R18438 VDD.n1487 VDD.n1486 146.341
R18439 VDD.n1489 VDD.n1427 146.341
R18440 VDD.n1496 VDD.n1419 146.341
R18441 VDD.n1500 VDD.n1498 146.341
R18442 VDD.n1506 VDD.n1415 146.341
R18443 VDD.n1510 VDD.n1508 146.341
R18444 VDD.n1518 VDD.n1411 146.341
R18445 VDD.n1521 VDD.n1520 146.341
R18446 VDD.n1523 VDD.n1406 146.341
R18447 VDD.n1530 VDD.n1402 146.341
R18448 VDD.n1534 VDD.n1532 146.341
R18449 VDD.n1540 VDD.n1398 146.341
R18450 VDD.n1544 VDD.n1542 146.341
R18451 VDD.n1550 VDD.n1394 146.341
R18452 VDD.n1554 VDD.n1552 146.341
R18453 VDD.n1560 VDD.n1387 146.341
R18454 VDD.n1564 VDD.n1562 146.341
R18455 VDD.n1570 VDD.n1383 146.341
R18456 VDD.n1575 VDD.n1572 146.341
R18457 VDD.n1573 VDD.n1380 146.341
R18458 VDD.n1375 VDD.n1373 146.341
R18459 VDD.n1588 VDD.n1368 146.341
R18460 VDD.n1594 VDD.n1368 146.341
R18461 VDD.n1594 VDD.n1360 146.341
R18462 VDD.n1604 VDD.n1360 146.341
R18463 VDD.n1604 VDD.n1356 146.341
R18464 VDD.n1610 VDD.n1356 146.341
R18465 VDD.n1610 VDD.n1349 146.341
R18466 VDD.n1620 VDD.n1349 146.341
R18467 VDD.n1620 VDD.n1345 146.341
R18468 VDD.n1626 VDD.n1345 146.341
R18469 VDD.n1626 VDD.n1337 146.341
R18470 VDD.n1636 VDD.n1337 146.341
R18471 VDD.n1636 VDD.n1333 146.341
R18472 VDD.n1642 VDD.n1333 146.341
R18473 VDD.n1642 VDD.n1325 146.341
R18474 VDD.n1652 VDD.n1325 146.341
R18475 VDD.n1652 VDD.n1321 146.341
R18476 VDD.n1658 VDD.n1321 146.341
R18477 VDD.n1658 VDD.n1313 146.341
R18478 VDD.n1668 VDD.n1313 146.341
R18479 VDD.n1668 VDD.n1309 146.341
R18480 VDD.n1674 VDD.n1309 146.341
R18481 VDD.n1674 VDD.n1302 146.341
R18482 VDD.n1684 VDD.n1302 146.341
R18483 VDD.n1684 VDD.n1293 146.341
R18484 VDD.n1690 VDD.n1293 146.341
R18485 VDD.n1690 VDD.n1285 146.341
R18486 VDD.n1700 VDD.n1285 146.341
R18487 VDD.n1700 VDD.n1281 146.341
R18488 VDD.n1706 VDD.n1281 146.341
R18489 VDD.n1706 VDD.n1273 146.341
R18490 VDD.n1716 VDD.n1273 146.341
R18491 VDD.n1716 VDD.n1269 146.341
R18492 VDD.n1722 VDD.n1269 146.341
R18493 VDD.n1722 VDD.n1261 146.341
R18494 VDD.n1732 VDD.n1261 146.341
R18495 VDD.n1732 VDD.n1257 146.341
R18496 VDD.n1738 VDD.n1257 146.341
R18497 VDD.n1738 VDD.n1250 146.341
R18498 VDD.n1748 VDD.n1250 146.341
R18499 VDD.n1748 VDD.n1246 146.341
R18500 VDD.n1754 VDD.n1246 146.341
R18501 VDD.n1754 VDD.n1237 146.341
R18502 VDD.n1766 VDD.n1237 146.341
R18503 VDD.n1766 VDD.n1232 146.341
R18504 VDD.n1803 VDD.n1232 146.341
R18505 VDD.n1377 VDD.n1376 114.812
R18506 VDD.n1391 VDD.n1390 114.812
R18507 VDD.n1408 VDD.n1407 114.812
R18508 VDD.n1422 VDD.n1421 114.812
R18509 VDD.n1439 VDD.n1438 114.812
R18510 VDD.n1143 VDD.n1142 114.812
R18511 VDD.n1226 VDD.n1225 114.812
R18512 VDD.n1203 VDD.n1202 114.812
R18513 VDD.n1183 VDD.n1182 114.812
R18514 VDD.n1162 VDD.n1161 114.812
R18515 VDD.n4364 VDD.n4363 114.812
R18516 VDD.n4343 VDD.n4342 114.812
R18517 VDD.n4323 VDD.n4322 114.812
R18518 VDD.n4302 VDD.n4301 114.812
R18519 VDD.n4279 VDD.n4278 114.812
R18520 VDD.n138 VDD.n137 114.812
R18521 VDD.n160 VDD.n159 114.812
R18522 VDD.n3945 VDD.n3944 114.812
R18523 VDD.n4034 VDD.n4033 114.812
R18524 VDD.n3965 VDD.n3964 114.812
R18525 VDD.n1115 VDD.n1114 112.874
R18526 VDD.n663 VDD.n662 112.874
R18527 VDD.n1135 VDD.n1134 112.874
R18528 VDD.n673 VDD.n672 112.874
R18529 VDD.n3118 VDD.n3117 112.874
R18530 VDD.n202 VDD.n201 112.874
R18531 VDD.n2922 VDD.n2921 112.874
R18532 VDD.n178 VDD.n177 112.874
R18533 VDD.n3425 VDD.n2902 109.2
R18534 VDD.n3920 VDD.n3919 99.5127
R18535 VDD.n3917 VDD.n194 99.5127
R18536 VDD.n3913 VDD.n3912 99.5127
R18537 VDD.n3910 VDD.n197 99.5127
R18538 VDD.n3904 VDD.n3903 99.5127
R18539 VDD.n3901 VDD.n200 99.5127
R18540 VDD.n3897 VDD.n3896 99.5127
R18541 VDD.n3894 VDD.n206 99.5127
R18542 VDD.n3388 VDD.n635 99.5127
R18543 VDD.n3385 VDD.n635 99.5127
R18544 VDD.n3385 VDD.n629 99.5127
R18545 VDD.n3382 VDD.n629 99.5127
R18546 VDD.n3382 VDD.n623 99.5127
R18547 VDD.n3379 VDD.n623 99.5127
R18548 VDD.n3379 VDD.n617 99.5127
R18549 VDD.n3376 VDD.n617 99.5127
R18550 VDD.n3376 VDD.n611 99.5127
R18551 VDD.n3373 VDD.n611 99.5127
R18552 VDD.n3373 VDD.n605 99.5127
R18553 VDD.n3370 VDD.n605 99.5127
R18554 VDD.n3370 VDD.n599 99.5127
R18555 VDD.n3114 VDD.n599 99.5127
R18556 VDD.n3114 VDD.n594 99.5127
R18557 VDD.n3111 VDD.n594 99.5127
R18558 VDD.n3111 VDD.n588 99.5127
R18559 VDD.n3108 VDD.n588 99.5127
R18560 VDD.n3108 VDD.n582 99.5127
R18561 VDD.n3105 VDD.n582 99.5127
R18562 VDD.n3105 VDD.n576 99.5127
R18563 VDD.n3102 VDD.n576 99.5127
R18564 VDD.n3102 VDD.n570 99.5127
R18565 VDD.n3099 VDD.n570 99.5127
R18566 VDD.n3099 VDD.n564 99.5127
R18567 VDD.n3096 VDD.n564 99.5127
R18568 VDD.n3096 VDD.n558 99.5127
R18569 VDD.n3093 VDD.n558 99.5127
R18570 VDD.n3093 VDD.n552 99.5127
R18571 VDD.n3090 VDD.n552 99.5127
R18572 VDD.n3090 VDD.n546 99.5127
R18573 VDD.n3087 VDD.n546 99.5127
R18574 VDD.n3087 VDD.n539 99.5127
R18575 VDD.n3084 VDD.n539 99.5127
R18576 VDD.n3084 VDD.n533 99.5127
R18577 VDD.n3081 VDD.n533 99.5127
R18578 VDD.n3081 VDD.n528 99.5127
R18579 VDD.n3078 VDD.n528 99.5127
R18580 VDD.n3078 VDD.n522 99.5127
R18581 VDD.n3075 VDD.n522 99.5127
R18582 VDD.n3075 VDD.n516 99.5127
R18583 VDD.n3072 VDD.n516 99.5127
R18584 VDD.n3072 VDD.n510 99.5127
R18585 VDD.n3069 VDD.n510 99.5127
R18586 VDD.n3069 VDD.n504 99.5127
R18587 VDD.n3066 VDD.n504 99.5127
R18588 VDD.n3066 VDD.n498 99.5127
R18589 VDD.n3063 VDD.n498 99.5127
R18590 VDD.n3063 VDD.n491 99.5127
R18591 VDD.n3060 VDD.n491 99.5127
R18592 VDD.n3060 VDD.n485 99.5127
R18593 VDD.n3057 VDD.n485 99.5127
R18594 VDD.n3057 VDD.n480 99.5127
R18595 VDD.n3054 VDD.n480 99.5127
R18596 VDD.n3054 VDD.n474 99.5127
R18597 VDD.n3051 VDD.n474 99.5127
R18598 VDD.n3051 VDD.n468 99.5127
R18599 VDD.n3048 VDD.n468 99.5127
R18600 VDD.n3048 VDD.n462 99.5127
R18601 VDD.n3045 VDD.n462 99.5127
R18602 VDD.n3045 VDD.n456 99.5127
R18603 VDD.n3042 VDD.n456 99.5127
R18604 VDD.n3042 VDD.n450 99.5127
R18605 VDD.n3039 VDD.n450 99.5127
R18606 VDD.n3039 VDD.n444 99.5127
R18607 VDD.n3036 VDD.n444 99.5127
R18608 VDD.n3036 VDD.n438 99.5127
R18609 VDD.n3033 VDD.n438 99.5127
R18610 VDD.n3033 VDD.n432 99.5127
R18611 VDD.n3030 VDD.n432 99.5127
R18612 VDD.n3030 VDD.n425 99.5127
R18613 VDD.n3027 VDD.n425 99.5127
R18614 VDD.n3027 VDD.n420 99.5127
R18615 VDD.n3024 VDD.n420 99.5127
R18616 VDD.n3024 VDD.n415 99.5127
R18617 VDD.n3021 VDD.n415 99.5127
R18618 VDD.n3021 VDD.n409 99.5127
R18619 VDD.n3018 VDD.n409 99.5127
R18620 VDD.n3018 VDD.n403 99.5127
R18621 VDD.n3015 VDD.n403 99.5127
R18622 VDD.n3015 VDD.n397 99.5127
R18623 VDD.n3012 VDD.n397 99.5127
R18624 VDD.n3012 VDD.n391 99.5127
R18625 VDD.n3009 VDD.n391 99.5127
R18626 VDD.n3009 VDD.n385 99.5127
R18627 VDD.n3006 VDD.n385 99.5127
R18628 VDD.n3006 VDD.n379 99.5127
R18629 VDD.n3003 VDD.n379 99.5127
R18630 VDD.n3003 VDD.n373 99.5127
R18631 VDD.n3000 VDD.n373 99.5127
R18632 VDD.n3000 VDD.n367 99.5127
R18633 VDD.n2997 VDD.n367 99.5127
R18634 VDD.n2997 VDD.n361 99.5127
R18635 VDD.n2994 VDD.n361 99.5127
R18636 VDD.n2994 VDD.n355 99.5127
R18637 VDD.n2991 VDD.n355 99.5127
R18638 VDD.n2991 VDD.n348 99.5127
R18639 VDD.n2988 VDD.n348 99.5127
R18640 VDD.n2988 VDD.n342 99.5127
R18641 VDD.n2985 VDD.n342 99.5127
R18642 VDD.n2985 VDD.n337 99.5127
R18643 VDD.n2982 VDD.n337 99.5127
R18644 VDD.n2982 VDD.n331 99.5127
R18645 VDD.n2979 VDD.n331 99.5127
R18646 VDD.n2979 VDD.n325 99.5127
R18647 VDD.n2976 VDD.n325 99.5127
R18648 VDD.n2976 VDD.n319 99.5127
R18649 VDD.n2973 VDD.n319 99.5127
R18650 VDD.n2973 VDD.n312 99.5127
R18651 VDD.n2970 VDD.n312 99.5127
R18652 VDD.n2970 VDD.n306 99.5127
R18653 VDD.n2967 VDD.n306 99.5127
R18654 VDD.n2967 VDD.n301 99.5127
R18655 VDD.n2964 VDD.n301 99.5127
R18656 VDD.n2964 VDD.n295 99.5127
R18657 VDD.n2961 VDD.n295 99.5127
R18658 VDD.n2961 VDD.n289 99.5127
R18659 VDD.n2958 VDD.n289 99.5127
R18660 VDD.n2958 VDD.n283 99.5127
R18661 VDD.n2955 VDD.n283 99.5127
R18662 VDD.n2955 VDD.n277 99.5127
R18663 VDD.n2952 VDD.n277 99.5127
R18664 VDD.n2952 VDD.n271 99.5127
R18665 VDD.n2949 VDD.n271 99.5127
R18666 VDD.n2949 VDD.n265 99.5127
R18667 VDD.n2946 VDD.n265 99.5127
R18668 VDD.n2946 VDD.n259 99.5127
R18669 VDD.n2943 VDD.n259 99.5127
R18670 VDD.n2943 VDD.n253 99.5127
R18671 VDD.n2940 VDD.n253 99.5127
R18672 VDD.n2940 VDD.n247 99.5127
R18673 VDD.n2937 VDD.n247 99.5127
R18674 VDD.n2937 VDD.n241 99.5127
R18675 VDD.n2934 VDD.n241 99.5127
R18676 VDD.n2934 VDD.n234 99.5127
R18677 VDD.n2931 VDD.n234 99.5127
R18678 VDD.n2931 VDD.n228 99.5127
R18679 VDD.n2928 VDD.n228 99.5127
R18680 VDD.n2928 VDD.n223 99.5127
R18681 VDD.n2925 VDD.n223 99.5127
R18682 VDD.n2925 VDD.n216 99.5127
R18683 VDD.n216 VDD.n208 99.5127
R18684 VDD.n3885 VDD.n208 99.5127
R18685 VDD.n3886 VDD.n3885 99.5127
R18686 VDD.n3886 VDD.n187 99.5127
R18687 VDD.n2920 VDD.n2919 99.5127
R18688 VDD.n3418 VDD.n2919 99.5127
R18689 VDD.n3416 VDD.n3415 99.5127
R18690 VDD.n3412 VDD.n3411 99.5127
R18691 VDD.n3408 VDD.n3407 99.5127
R18692 VDD.n3404 VDD.n3403 99.5127
R18693 VDD.n3400 VDD.n3399 99.5127
R18694 VDD.n3395 VDD.n3394 99.5127
R18695 VDD.n3391 VDD.n2910 99.5127
R18696 VDD.n3433 VDD.n633 99.5127
R18697 VDD.n3433 VDD.n631 99.5127
R18698 VDD.n3437 VDD.n631 99.5127
R18699 VDD.n3437 VDD.n621 99.5127
R18700 VDD.n3445 VDD.n621 99.5127
R18701 VDD.n3445 VDD.n619 99.5127
R18702 VDD.n3449 VDD.n619 99.5127
R18703 VDD.n3449 VDD.n609 99.5127
R18704 VDD.n3457 VDD.n609 99.5127
R18705 VDD.n3457 VDD.n607 99.5127
R18706 VDD.n3461 VDD.n607 99.5127
R18707 VDD.n3461 VDD.n598 99.5127
R18708 VDD.n3469 VDD.n598 99.5127
R18709 VDD.n3469 VDD.n596 99.5127
R18710 VDD.n3473 VDD.n596 99.5127
R18711 VDD.n3473 VDD.n586 99.5127
R18712 VDD.n3481 VDD.n586 99.5127
R18713 VDD.n3481 VDD.n584 99.5127
R18714 VDD.n3485 VDD.n584 99.5127
R18715 VDD.n3485 VDD.n574 99.5127
R18716 VDD.n3493 VDD.n574 99.5127
R18717 VDD.n3493 VDD.n572 99.5127
R18718 VDD.n3497 VDD.n572 99.5127
R18719 VDD.n3497 VDD.n562 99.5127
R18720 VDD.n3505 VDD.n562 99.5127
R18721 VDD.n3505 VDD.n560 99.5127
R18722 VDD.n3509 VDD.n560 99.5127
R18723 VDD.n3509 VDD.n550 99.5127
R18724 VDD.n3517 VDD.n550 99.5127
R18725 VDD.n3517 VDD.n548 99.5127
R18726 VDD.n3521 VDD.n548 99.5127
R18727 VDD.n3521 VDD.n537 99.5127
R18728 VDD.n3529 VDD.n537 99.5127
R18729 VDD.n3529 VDD.n535 99.5127
R18730 VDD.n3533 VDD.n535 99.5127
R18731 VDD.n3533 VDD.n526 99.5127
R18732 VDD.n3541 VDD.n526 99.5127
R18733 VDD.n3541 VDD.n524 99.5127
R18734 VDD.n3545 VDD.n524 99.5127
R18735 VDD.n3545 VDD.n514 99.5127
R18736 VDD.n3553 VDD.n514 99.5127
R18737 VDD.n3553 VDD.n512 99.5127
R18738 VDD.n3557 VDD.n512 99.5127
R18739 VDD.n3557 VDD.n502 99.5127
R18740 VDD.n3565 VDD.n502 99.5127
R18741 VDD.n3565 VDD.n500 99.5127
R18742 VDD.n3569 VDD.n500 99.5127
R18743 VDD.n3569 VDD.n489 99.5127
R18744 VDD.n3577 VDD.n489 99.5127
R18745 VDD.n3577 VDD.n487 99.5127
R18746 VDD.n3581 VDD.n487 99.5127
R18747 VDD.n3581 VDD.n478 99.5127
R18748 VDD.n3589 VDD.n478 99.5127
R18749 VDD.n3589 VDD.n476 99.5127
R18750 VDD.n3593 VDD.n476 99.5127
R18751 VDD.n3593 VDD.n466 99.5127
R18752 VDD.n3601 VDD.n466 99.5127
R18753 VDD.n3601 VDD.n464 99.5127
R18754 VDD.n3605 VDD.n464 99.5127
R18755 VDD.n3605 VDD.n454 99.5127
R18756 VDD.n3613 VDD.n454 99.5127
R18757 VDD.n3613 VDD.n452 99.5127
R18758 VDD.n3617 VDD.n452 99.5127
R18759 VDD.n3617 VDD.n442 99.5127
R18760 VDD.n3625 VDD.n442 99.5127
R18761 VDD.n3625 VDD.n440 99.5127
R18762 VDD.n3629 VDD.n440 99.5127
R18763 VDD.n3629 VDD.n430 99.5127
R18764 VDD.n3637 VDD.n430 99.5127
R18765 VDD.n3637 VDD.n428 99.5127
R18766 VDD.n3641 VDD.n428 99.5127
R18767 VDD.n3641 VDD.n419 99.5127
R18768 VDD.n3649 VDD.n419 99.5127
R18769 VDD.n3649 VDD.n417 99.5127
R18770 VDD.n3653 VDD.n417 99.5127
R18771 VDD.n3653 VDD.n407 99.5127
R18772 VDD.n3661 VDD.n407 99.5127
R18773 VDD.n3661 VDD.n405 99.5127
R18774 VDD.n3665 VDD.n405 99.5127
R18775 VDD.n3665 VDD.n395 99.5127
R18776 VDD.n3673 VDD.n395 99.5127
R18777 VDD.n3673 VDD.n393 99.5127
R18778 VDD.n3677 VDD.n393 99.5127
R18779 VDD.n3677 VDD.n383 99.5127
R18780 VDD.n3685 VDD.n383 99.5127
R18781 VDD.n3685 VDD.n381 99.5127
R18782 VDD.n3689 VDD.n381 99.5127
R18783 VDD.n3689 VDD.n371 99.5127
R18784 VDD.n3697 VDD.n371 99.5127
R18785 VDD.n3697 VDD.n369 99.5127
R18786 VDD.n3701 VDD.n369 99.5127
R18787 VDD.n3701 VDD.n359 99.5127
R18788 VDD.n3709 VDD.n359 99.5127
R18789 VDD.n3709 VDD.n357 99.5127
R18790 VDD.n3713 VDD.n357 99.5127
R18791 VDD.n3713 VDD.n346 99.5127
R18792 VDD.n3721 VDD.n346 99.5127
R18793 VDD.n3721 VDD.n344 99.5127
R18794 VDD.n3725 VDD.n344 99.5127
R18795 VDD.n3725 VDD.n335 99.5127
R18796 VDD.n3733 VDD.n335 99.5127
R18797 VDD.n3733 VDD.n333 99.5127
R18798 VDD.n3737 VDD.n333 99.5127
R18799 VDD.n3737 VDD.n323 99.5127
R18800 VDD.n3745 VDD.n323 99.5127
R18801 VDD.n3745 VDD.n321 99.5127
R18802 VDD.n3749 VDD.n321 99.5127
R18803 VDD.n3749 VDD.n310 99.5127
R18804 VDD.n3757 VDD.n310 99.5127
R18805 VDD.n3757 VDD.n308 99.5127
R18806 VDD.n3761 VDD.n308 99.5127
R18807 VDD.n3761 VDD.n299 99.5127
R18808 VDD.n3769 VDD.n299 99.5127
R18809 VDD.n3769 VDD.n297 99.5127
R18810 VDD.n3773 VDD.n297 99.5127
R18811 VDD.n3773 VDD.n287 99.5127
R18812 VDD.n3781 VDD.n287 99.5127
R18813 VDD.n3781 VDD.n285 99.5127
R18814 VDD.n3785 VDD.n285 99.5127
R18815 VDD.n3785 VDD.n275 99.5127
R18816 VDD.n3793 VDD.n275 99.5127
R18817 VDD.n3793 VDD.n273 99.5127
R18818 VDD.n3797 VDD.n273 99.5127
R18819 VDD.n3797 VDD.n263 99.5127
R18820 VDD.n3805 VDD.n263 99.5127
R18821 VDD.n3805 VDD.n261 99.5127
R18822 VDD.n3809 VDD.n261 99.5127
R18823 VDD.n3809 VDD.n251 99.5127
R18824 VDD.n3817 VDD.n251 99.5127
R18825 VDD.n3817 VDD.n249 99.5127
R18826 VDD.n3821 VDD.n249 99.5127
R18827 VDD.n3821 VDD.n239 99.5127
R18828 VDD.n3829 VDD.n239 99.5127
R18829 VDD.n3829 VDD.n237 99.5127
R18830 VDD.n3833 VDD.n237 99.5127
R18831 VDD.n3833 VDD.n227 99.5127
R18832 VDD.n3841 VDD.n227 99.5127
R18833 VDD.n3841 VDD.n225 99.5127
R18834 VDD.n3845 VDD.n225 99.5127
R18835 VDD.n3845 VDD.n214 99.5127
R18836 VDD.n3879 VDD.n214 99.5127
R18837 VDD.n3879 VDD.n212 99.5127
R18838 VDD.n3883 VDD.n212 99.5127
R18839 VDD.n3883 VDD.n189 99.5127
R18840 VDD.n3924 VDD.n189 99.5127
R18841 VDD.n2856 VDD.n2855 99.5127
R18842 VDD.n2852 VDD.n2851 99.5127
R18843 VDD.n2848 VDD.n2847 99.5127
R18844 VDD.n2844 VDD.n2843 99.5127
R18845 VDD.n2840 VDD.n2839 99.5127
R18846 VDD.n2836 VDD.n2835 99.5127
R18847 VDD.n2832 VDD.n2831 99.5127
R18848 VDD.n2828 VDD.n2827 99.5127
R18849 VDD.n1936 VDD.n1103 99.5127
R18850 VDD.n1936 VDD.n1097 99.5127
R18851 VDD.n1939 VDD.n1097 99.5127
R18852 VDD.n1939 VDD.n1091 99.5127
R18853 VDD.n1942 VDD.n1091 99.5127
R18854 VDD.n1942 VDD.n1085 99.5127
R18855 VDD.n1945 VDD.n1085 99.5127
R18856 VDD.n1945 VDD.n1079 99.5127
R18857 VDD.n1948 VDD.n1079 99.5127
R18858 VDD.n1948 VDD.n1072 99.5127
R18859 VDD.n1951 VDD.n1072 99.5127
R18860 VDD.n1951 VDD.n1066 99.5127
R18861 VDD.n1954 VDD.n1066 99.5127
R18862 VDD.n1954 VDD.n1061 99.5127
R18863 VDD.n1957 VDD.n1061 99.5127
R18864 VDD.n1957 VDD.n1055 99.5127
R18865 VDD.n1960 VDD.n1055 99.5127
R18866 VDD.n1960 VDD.n1049 99.5127
R18867 VDD.n1963 VDD.n1049 99.5127
R18868 VDD.n1963 VDD.n1043 99.5127
R18869 VDD.n1966 VDD.n1043 99.5127
R18870 VDD.n1966 VDD.n1037 99.5127
R18871 VDD.n1969 VDD.n1037 99.5127
R18872 VDD.n1969 VDD.n1031 99.5127
R18873 VDD.n1972 VDD.n1031 99.5127
R18874 VDD.n1972 VDD.n1024 99.5127
R18875 VDD.n1975 VDD.n1024 99.5127
R18876 VDD.n1975 VDD.n1018 99.5127
R18877 VDD.n1978 VDD.n1018 99.5127
R18878 VDD.n1978 VDD.n1013 99.5127
R18879 VDD.n1981 VDD.n1013 99.5127
R18880 VDD.n1981 VDD.n1007 99.5127
R18881 VDD.n1984 VDD.n1007 99.5127
R18882 VDD.n1984 VDD.n1001 99.5127
R18883 VDD.n1987 VDD.n1001 99.5127
R18884 VDD.n1987 VDD.n995 99.5127
R18885 VDD.n1990 VDD.n995 99.5127
R18886 VDD.n1990 VDD.n989 99.5127
R18887 VDD.n1993 VDD.n989 99.5127
R18888 VDD.n1993 VDD.n983 99.5127
R18889 VDD.n1996 VDD.n983 99.5127
R18890 VDD.n1996 VDD.n977 99.5127
R18891 VDD.n1999 VDD.n977 99.5127
R18892 VDD.n1999 VDD.n971 99.5127
R18893 VDD.n2002 VDD.n971 99.5127
R18894 VDD.n2002 VDD.n965 99.5127
R18895 VDD.n2005 VDD.n965 99.5127
R18896 VDD.n2005 VDD.n959 99.5127
R18897 VDD.n2008 VDD.n959 99.5127
R18898 VDD.n2008 VDD.n953 99.5127
R18899 VDD.n2011 VDD.n953 99.5127
R18900 VDD.n2011 VDD.n946 99.5127
R18901 VDD.n2014 VDD.n946 99.5127
R18902 VDD.n2014 VDD.n940 99.5127
R18903 VDD.n2017 VDD.n940 99.5127
R18904 VDD.n2017 VDD.n935 99.5127
R18905 VDD.n2020 VDD.n935 99.5127
R18906 VDD.n2020 VDD.n929 99.5127
R18907 VDD.n2023 VDD.n929 99.5127
R18908 VDD.n2023 VDD.n923 99.5127
R18909 VDD.n2026 VDD.n923 99.5127
R18910 VDD.n2026 VDD.n917 99.5127
R18911 VDD.n2029 VDD.n917 99.5127
R18912 VDD.n2029 VDD.n911 99.5127
R18913 VDD.n2032 VDD.n911 99.5127
R18914 VDD.n2032 VDD.n905 99.5127
R18915 VDD.n2035 VDD.n905 99.5127
R18916 VDD.n2035 VDD.n899 99.5127
R18917 VDD.n2038 VDD.n899 99.5127
R18918 VDD.n2038 VDD.n893 99.5127
R18919 VDD.n2041 VDD.n893 99.5127
R18920 VDD.n2041 VDD.n887 99.5127
R18921 VDD.n2044 VDD.n887 99.5127
R18922 VDD.n2044 VDD.n881 99.5127
R18923 VDD.n2047 VDD.n881 99.5127
R18924 VDD.n2047 VDD.n875 99.5127
R18925 VDD.n2050 VDD.n875 99.5127
R18926 VDD.n2050 VDD.n870 99.5127
R18927 VDD.n2053 VDD.n870 99.5127
R18928 VDD.n2053 VDD.n864 99.5127
R18929 VDD.n2056 VDD.n864 99.5127
R18930 VDD.n2056 VDD.n858 99.5127
R18931 VDD.n2059 VDD.n858 99.5127
R18932 VDD.n2059 VDD.n852 99.5127
R18933 VDD.n2062 VDD.n852 99.5127
R18934 VDD.n2062 VDD.n846 99.5127
R18935 VDD.n2065 VDD.n846 99.5127
R18936 VDD.n2065 VDD.n840 99.5127
R18937 VDD.n2068 VDD.n840 99.5127
R18938 VDD.n2068 VDD.n833 99.5127
R18939 VDD.n2071 VDD.n833 99.5127
R18940 VDD.n2071 VDD.n827 99.5127
R18941 VDD.n2074 VDD.n827 99.5127
R18942 VDD.n2074 VDD.n822 99.5127
R18943 VDD.n2077 VDD.n822 99.5127
R18944 VDD.n2077 VDD.n816 99.5127
R18945 VDD.n2080 VDD.n816 99.5127
R18946 VDD.n2080 VDD.n810 99.5127
R18947 VDD.n2083 VDD.n810 99.5127
R18948 VDD.n2083 VDD.n804 99.5127
R18949 VDD.n2086 VDD.n804 99.5127
R18950 VDD.n2086 VDD.n798 99.5127
R18951 VDD.n2089 VDD.n798 99.5127
R18952 VDD.n2089 VDD.n792 99.5127
R18953 VDD.n2092 VDD.n792 99.5127
R18954 VDD.n2092 VDD.n786 99.5127
R18955 VDD.n2095 VDD.n786 99.5127
R18956 VDD.n2095 VDD.n780 99.5127
R18957 VDD.n2098 VDD.n780 99.5127
R18958 VDD.n2098 VDD.n774 99.5127
R18959 VDD.n2101 VDD.n774 99.5127
R18960 VDD.n2101 VDD.n767 99.5127
R18961 VDD.n2104 VDD.n767 99.5127
R18962 VDD.n2104 VDD.n761 99.5127
R18963 VDD.n2107 VDD.n761 99.5127
R18964 VDD.n2107 VDD.n756 99.5127
R18965 VDD.n2110 VDD.n756 99.5127
R18966 VDD.n2110 VDD.n750 99.5127
R18967 VDD.n2113 VDD.n750 99.5127
R18968 VDD.n2113 VDD.n744 99.5127
R18969 VDD.n2116 VDD.n744 99.5127
R18970 VDD.n2116 VDD.n738 99.5127
R18971 VDD.n2119 VDD.n738 99.5127
R18972 VDD.n2119 VDD.n732 99.5127
R18973 VDD.n2122 VDD.n732 99.5127
R18974 VDD.n2122 VDD.n726 99.5127
R18975 VDD.n2125 VDD.n726 99.5127
R18976 VDD.n2125 VDD.n720 99.5127
R18977 VDD.n2128 VDD.n720 99.5127
R18978 VDD.n2128 VDD.n714 99.5127
R18979 VDD.n2131 VDD.n714 99.5127
R18980 VDD.n2131 VDD.n708 99.5127
R18981 VDD.n2146 VDD.n708 99.5127
R18982 VDD.n2146 VDD.n702 99.5127
R18983 VDD.n2142 VDD.n702 99.5127
R18984 VDD.n2142 VDD.n697 99.5127
R18985 VDD.n2139 VDD.n697 99.5127
R18986 VDD.n2139 VDD.n691 99.5127
R18987 VDD.n2136 VDD.n691 99.5127
R18988 VDD.n2136 VDD.n684 99.5127
R18989 VDD.n684 VDD.n676 99.5127
R18990 VDD.n2818 VDD.n676 99.5127
R18991 VDD.n2819 VDD.n2818 99.5127
R18992 VDD.n2819 VDD.n667 99.5127
R18993 VDD.n2823 VDD.n667 99.5127
R18994 VDD.n1901 VDD.n1899 99.5127
R18995 VDD.n1905 VDD.n1899 99.5127
R18996 VDD.n1909 VDD.n1907 99.5127
R18997 VDD.n1913 VDD.n1897 99.5127
R18998 VDD.n1917 VDD.n1915 99.5127
R18999 VDD.n1921 VDD.n1137 99.5127
R19000 VDD.n1925 VDD.n1923 99.5127
R19001 VDD.n1930 VDD.n1133 99.5127
R19002 VDD.n1933 VDD.n1932 99.5127
R19003 VDD.n2387 VDD.n1099 99.5127
R19004 VDD.n2391 VDD.n1099 99.5127
R19005 VDD.n2391 VDD.n1089 99.5127
R19006 VDD.n2399 VDD.n1089 99.5127
R19007 VDD.n2399 VDD.n1087 99.5127
R19008 VDD.n2403 VDD.n1087 99.5127
R19009 VDD.n2403 VDD.n1077 99.5127
R19010 VDD.n2411 VDD.n1077 99.5127
R19011 VDD.n2411 VDD.n1075 99.5127
R19012 VDD.n2415 VDD.n1075 99.5127
R19013 VDD.n2415 VDD.n1065 99.5127
R19014 VDD.n2423 VDD.n1065 99.5127
R19015 VDD.n2423 VDD.n1063 99.5127
R19016 VDD.n2427 VDD.n1063 99.5127
R19017 VDD.n2427 VDD.n1053 99.5127
R19018 VDD.n2435 VDD.n1053 99.5127
R19019 VDD.n2435 VDD.n1051 99.5127
R19020 VDD.n2439 VDD.n1051 99.5127
R19021 VDD.n2439 VDD.n1041 99.5127
R19022 VDD.n2447 VDD.n1041 99.5127
R19023 VDD.n2447 VDD.n1039 99.5127
R19024 VDD.n2451 VDD.n1039 99.5127
R19025 VDD.n2451 VDD.n1029 99.5127
R19026 VDD.n2459 VDD.n1029 99.5127
R19027 VDD.n2459 VDD.n1027 99.5127
R19028 VDD.n2463 VDD.n1027 99.5127
R19029 VDD.n2463 VDD.n1017 99.5127
R19030 VDD.n2471 VDD.n1017 99.5127
R19031 VDD.n2471 VDD.n1015 99.5127
R19032 VDD.n2475 VDD.n1015 99.5127
R19033 VDD.n2475 VDD.n1005 99.5127
R19034 VDD.n2483 VDD.n1005 99.5127
R19035 VDD.n2483 VDD.n1003 99.5127
R19036 VDD.n2487 VDD.n1003 99.5127
R19037 VDD.n2487 VDD.n993 99.5127
R19038 VDD.n2495 VDD.n993 99.5127
R19039 VDD.n2495 VDD.n991 99.5127
R19040 VDD.n2499 VDD.n991 99.5127
R19041 VDD.n2499 VDD.n981 99.5127
R19042 VDD.n2507 VDD.n981 99.5127
R19043 VDD.n2507 VDD.n979 99.5127
R19044 VDD.n2511 VDD.n979 99.5127
R19045 VDD.n2511 VDD.n969 99.5127
R19046 VDD.n2519 VDD.n969 99.5127
R19047 VDD.n2519 VDD.n967 99.5127
R19048 VDD.n2523 VDD.n967 99.5127
R19049 VDD.n2523 VDD.n957 99.5127
R19050 VDD.n2531 VDD.n957 99.5127
R19051 VDD.n2531 VDD.n955 99.5127
R19052 VDD.n2535 VDD.n955 99.5127
R19053 VDD.n2535 VDD.n944 99.5127
R19054 VDD.n2543 VDD.n944 99.5127
R19055 VDD.n2543 VDD.n942 99.5127
R19056 VDD.n2547 VDD.n942 99.5127
R19057 VDD.n2547 VDD.n933 99.5127
R19058 VDD.n2555 VDD.n933 99.5127
R19059 VDD.n2555 VDD.n931 99.5127
R19060 VDD.n2559 VDD.n931 99.5127
R19061 VDD.n2559 VDD.n921 99.5127
R19062 VDD.n2567 VDD.n921 99.5127
R19063 VDD.n2567 VDD.n919 99.5127
R19064 VDD.n2571 VDD.n919 99.5127
R19065 VDD.n2571 VDD.n909 99.5127
R19066 VDD.n2579 VDD.n909 99.5127
R19067 VDD.n2579 VDD.n907 99.5127
R19068 VDD.n2583 VDD.n907 99.5127
R19069 VDD.n2583 VDD.n897 99.5127
R19070 VDD.n2591 VDD.n897 99.5127
R19071 VDD.n2591 VDD.n895 99.5127
R19072 VDD.n2595 VDD.n895 99.5127
R19073 VDD.n2595 VDD.n885 99.5127
R19074 VDD.n2603 VDD.n885 99.5127
R19075 VDD.n2603 VDD.n883 99.5127
R19076 VDD.n2607 VDD.n883 99.5127
R19077 VDD.n2607 VDD.n874 99.5127
R19078 VDD.n2615 VDD.n874 99.5127
R19079 VDD.n2615 VDD.n872 99.5127
R19080 VDD.n2619 VDD.n872 99.5127
R19081 VDD.n2619 VDD.n862 99.5127
R19082 VDD.n2627 VDD.n862 99.5127
R19083 VDD.n2627 VDD.n860 99.5127
R19084 VDD.n2631 VDD.n860 99.5127
R19085 VDD.n2631 VDD.n850 99.5127
R19086 VDD.n2639 VDD.n850 99.5127
R19087 VDD.n2639 VDD.n848 99.5127
R19088 VDD.n2643 VDD.n848 99.5127
R19089 VDD.n2643 VDD.n838 99.5127
R19090 VDD.n2651 VDD.n838 99.5127
R19091 VDD.n2651 VDD.n836 99.5127
R19092 VDD.n2655 VDD.n836 99.5127
R19093 VDD.n2655 VDD.n826 99.5127
R19094 VDD.n2663 VDD.n826 99.5127
R19095 VDD.n2663 VDD.n824 99.5127
R19096 VDD.n2667 VDD.n824 99.5127
R19097 VDD.n2667 VDD.n814 99.5127
R19098 VDD.n2675 VDD.n814 99.5127
R19099 VDD.n2675 VDD.n812 99.5127
R19100 VDD.n2679 VDD.n812 99.5127
R19101 VDD.n2679 VDD.n802 99.5127
R19102 VDD.n2687 VDD.n802 99.5127
R19103 VDD.n2687 VDD.n800 99.5127
R19104 VDD.n2691 VDD.n800 99.5127
R19105 VDD.n2691 VDD.n790 99.5127
R19106 VDD.n2699 VDD.n790 99.5127
R19107 VDD.n2699 VDD.n788 99.5127
R19108 VDD.n2703 VDD.n788 99.5127
R19109 VDD.n2703 VDD.n778 99.5127
R19110 VDD.n2711 VDD.n778 99.5127
R19111 VDD.n2711 VDD.n776 99.5127
R19112 VDD.n2715 VDD.n776 99.5127
R19113 VDD.n2715 VDD.n765 99.5127
R19114 VDD.n2723 VDD.n765 99.5127
R19115 VDD.n2723 VDD.n763 99.5127
R19116 VDD.n2727 VDD.n763 99.5127
R19117 VDD.n2727 VDD.n754 99.5127
R19118 VDD.n2735 VDD.n754 99.5127
R19119 VDD.n2735 VDD.n752 99.5127
R19120 VDD.n2739 VDD.n752 99.5127
R19121 VDD.n2739 VDD.n742 99.5127
R19122 VDD.n2747 VDD.n742 99.5127
R19123 VDD.n2747 VDD.n740 99.5127
R19124 VDD.n2751 VDD.n740 99.5127
R19125 VDD.n2751 VDD.n730 99.5127
R19126 VDD.n2759 VDD.n730 99.5127
R19127 VDD.n2759 VDD.n728 99.5127
R19128 VDD.n2763 VDD.n728 99.5127
R19129 VDD.n2763 VDD.n718 99.5127
R19130 VDD.n2771 VDD.n718 99.5127
R19131 VDD.n2771 VDD.n716 99.5127
R19132 VDD.n2775 VDD.n716 99.5127
R19133 VDD.n2775 VDD.n706 99.5127
R19134 VDD.n2783 VDD.n706 99.5127
R19135 VDD.n2783 VDD.n704 99.5127
R19136 VDD.n2787 VDD.n704 99.5127
R19137 VDD.n2787 VDD.n695 99.5127
R19138 VDD.n2795 VDD.n695 99.5127
R19139 VDD.n2795 VDD.n693 99.5127
R19140 VDD.n2799 VDD.n693 99.5127
R19141 VDD.n2799 VDD.n682 99.5127
R19142 VDD.n2812 VDD.n682 99.5127
R19143 VDD.n2812 VDD.n680 99.5127
R19144 VDD.n2816 VDD.n680 99.5127
R19145 VDD.n2816 VDD.n669 99.5127
R19146 VDD.n2862 VDD.n669 99.5127
R19147 VDD.n2862 VDD.n670 99.5127
R19148 VDD.n3867 VDD.n3866 99.5127
R19149 VDD.n3864 VDD.n3852 99.5127
R19150 VDD.n3860 VDD.n3859 99.5127
R19151 VDD.n3857 VDD.n3855 99.5127
R19152 VDD.n3941 VDD.n3940 99.5127
R19153 VDD.n3938 VDD.n176 99.5127
R19154 VDD.n3934 VDD.n3933 99.5127
R19155 VDD.n3931 VDD.n182 99.5127
R19156 VDD.n3152 VDD.n636 99.5127
R19157 VDD.n3155 VDD.n636 99.5127
R19158 VDD.n3155 VDD.n630 99.5127
R19159 VDD.n3158 VDD.n630 99.5127
R19160 VDD.n3158 VDD.n624 99.5127
R19161 VDD.n3161 VDD.n624 99.5127
R19162 VDD.n3161 VDD.n618 99.5127
R19163 VDD.n3164 VDD.n618 99.5127
R19164 VDD.n3164 VDD.n612 99.5127
R19165 VDD.n3167 VDD.n612 99.5127
R19166 VDD.n3167 VDD.n606 99.5127
R19167 VDD.n3368 VDD.n606 99.5127
R19168 VDD.n3368 VDD.n600 99.5127
R19169 VDD.n3364 VDD.n600 99.5127
R19170 VDD.n3364 VDD.n595 99.5127
R19171 VDD.n3361 VDD.n595 99.5127
R19172 VDD.n3361 VDD.n589 99.5127
R19173 VDD.n3358 VDD.n589 99.5127
R19174 VDD.n3358 VDD.n583 99.5127
R19175 VDD.n3355 VDD.n583 99.5127
R19176 VDD.n3355 VDD.n577 99.5127
R19177 VDD.n3352 VDD.n577 99.5127
R19178 VDD.n3352 VDD.n571 99.5127
R19179 VDD.n3349 VDD.n571 99.5127
R19180 VDD.n3349 VDD.n565 99.5127
R19181 VDD.n3346 VDD.n565 99.5127
R19182 VDD.n3346 VDD.n559 99.5127
R19183 VDD.n3343 VDD.n559 99.5127
R19184 VDD.n3343 VDD.n553 99.5127
R19185 VDD.n3340 VDD.n553 99.5127
R19186 VDD.n3340 VDD.n547 99.5127
R19187 VDD.n3337 VDD.n547 99.5127
R19188 VDD.n3337 VDD.n540 99.5127
R19189 VDD.n3334 VDD.n540 99.5127
R19190 VDD.n3334 VDD.n534 99.5127
R19191 VDD.n3331 VDD.n534 99.5127
R19192 VDD.n3331 VDD.n529 99.5127
R19193 VDD.n3328 VDD.n529 99.5127
R19194 VDD.n3328 VDD.n523 99.5127
R19195 VDD.n3325 VDD.n523 99.5127
R19196 VDD.n3325 VDD.n517 99.5127
R19197 VDD.n3322 VDD.n517 99.5127
R19198 VDD.n3322 VDD.n511 99.5127
R19199 VDD.n3319 VDD.n511 99.5127
R19200 VDD.n3319 VDD.n505 99.5127
R19201 VDD.n3316 VDD.n505 99.5127
R19202 VDD.n3316 VDD.n499 99.5127
R19203 VDD.n3313 VDD.n499 99.5127
R19204 VDD.n3313 VDD.n492 99.5127
R19205 VDD.n3310 VDD.n492 99.5127
R19206 VDD.n3310 VDD.n486 99.5127
R19207 VDD.n3307 VDD.n486 99.5127
R19208 VDD.n3307 VDD.n481 99.5127
R19209 VDD.n3304 VDD.n481 99.5127
R19210 VDD.n3304 VDD.n475 99.5127
R19211 VDD.n3301 VDD.n475 99.5127
R19212 VDD.n3301 VDD.n469 99.5127
R19213 VDD.n3298 VDD.n469 99.5127
R19214 VDD.n3298 VDD.n463 99.5127
R19215 VDD.n3295 VDD.n463 99.5127
R19216 VDD.n3295 VDD.n457 99.5127
R19217 VDD.n3292 VDD.n457 99.5127
R19218 VDD.n3292 VDD.n451 99.5127
R19219 VDD.n3289 VDD.n451 99.5127
R19220 VDD.n3289 VDD.n445 99.5127
R19221 VDD.n3286 VDD.n445 99.5127
R19222 VDD.n3286 VDD.n439 99.5127
R19223 VDD.n3283 VDD.n439 99.5127
R19224 VDD.n3283 VDD.n433 99.5127
R19225 VDD.n3280 VDD.n433 99.5127
R19226 VDD.n3280 VDD.n426 99.5127
R19227 VDD.n3277 VDD.n426 99.5127
R19228 VDD.n3277 VDD.n421 99.5127
R19229 VDD.n3274 VDD.n421 99.5127
R19230 VDD.n3274 VDD.n416 99.5127
R19231 VDD.n3271 VDD.n416 99.5127
R19232 VDD.n3271 VDD.n410 99.5127
R19233 VDD.n3268 VDD.n410 99.5127
R19234 VDD.n3268 VDD.n404 99.5127
R19235 VDD.n3265 VDD.n404 99.5127
R19236 VDD.n3265 VDD.n398 99.5127
R19237 VDD.n3262 VDD.n398 99.5127
R19238 VDD.n3262 VDD.n392 99.5127
R19239 VDD.n3259 VDD.n392 99.5127
R19240 VDD.n3259 VDD.n386 99.5127
R19241 VDD.n3256 VDD.n386 99.5127
R19242 VDD.n3256 VDD.n380 99.5127
R19243 VDD.n3253 VDD.n380 99.5127
R19244 VDD.n3253 VDD.n374 99.5127
R19245 VDD.n3250 VDD.n374 99.5127
R19246 VDD.n3250 VDD.n368 99.5127
R19247 VDD.n3247 VDD.n368 99.5127
R19248 VDD.n3247 VDD.n362 99.5127
R19249 VDD.n3244 VDD.n362 99.5127
R19250 VDD.n3244 VDD.n356 99.5127
R19251 VDD.n3241 VDD.n356 99.5127
R19252 VDD.n3241 VDD.n349 99.5127
R19253 VDD.n3238 VDD.n349 99.5127
R19254 VDD.n3238 VDD.n343 99.5127
R19255 VDD.n3235 VDD.n343 99.5127
R19256 VDD.n3235 VDD.n338 99.5127
R19257 VDD.n3232 VDD.n338 99.5127
R19258 VDD.n3232 VDD.n332 99.5127
R19259 VDD.n3229 VDD.n332 99.5127
R19260 VDD.n3229 VDD.n326 99.5127
R19261 VDD.n3226 VDD.n326 99.5127
R19262 VDD.n3226 VDD.n320 99.5127
R19263 VDD.n3223 VDD.n320 99.5127
R19264 VDD.n3223 VDD.n313 99.5127
R19265 VDD.n3220 VDD.n313 99.5127
R19266 VDD.n3220 VDD.n307 99.5127
R19267 VDD.n3217 VDD.n307 99.5127
R19268 VDD.n3217 VDD.n302 99.5127
R19269 VDD.n3214 VDD.n302 99.5127
R19270 VDD.n3214 VDD.n296 99.5127
R19271 VDD.n3211 VDD.n296 99.5127
R19272 VDD.n3211 VDD.n290 99.5127
R19273 VDD.n3208 VDD.n290 99.5127
R19274 VDD.n3208 VDD.n284 99.5127
R19275 VDD.n3205 VDD.n284 99.5127
R19276 VDD.n3205 VDD.n278 99.5127
R19277 VDD.n3202 VDD.n278 99.5127
R19278 VDD.n3202 VDD.n272 99.5127
R19279 VDD.n3199 VDD.n272 99.5127
R19280 VDD.n3199 VDD.n266 99.5127
R19281 VDD.n3196 VDD.n266 99.5127
R19282 VDD.n3196 VDD.n260 99.5127
R19283 VDD.n3193 VDD.n260 99.5127
R19284 VDD.n3193 VDD.n254 99.5127
R19285 VDD.n3190 VDD.n254 99.5127
R19286 VDD.n3190 VDD.n248 99.5127
R19287 VDD.n3187 VDD.n248 99.5127
R19288 VDD.n3187 VDD.n242 99.5127
R19289 VDD.n3184 VDD.n242 99.5127
R19290 VDD.n3184 VDD.n235 99.5127
R19291 VDD.n3181 VDD.n235 99.5127
R19292 VDD.n3181 VDD.n229 99.5127
R19293 VDD.n3178 VDD.n229 99.5127
R19294 VDD.n3178 VDD.n224 99.5127
R19295 VDD.n3175 VDD.n224 99.5127
R19296 VDD.n3175 VDD.n217 99.5127
R19297 VDD.n3172 VDD.n217 99.5127
R19298 VDD.n3172 VDD.n210 99.5127
R19299 VDD.n210 VDD.n185 99.5127
R19300 VDD.n3926 VDD.n185 99.5127
R19301 VDD.n3120 VDD.n639 99.5127
R19302 VDD.n3124 VDD.n3123 99.5127
R19303 VDD.n3128 VDD.n3127 99.5127
R19304 VDD.n3132 VDD.n3131 99.5127
R19305 VDD.n3136 VDD.n3135 99.5127
R19306 VDD.n3140 VDD.n3139 99.5127
R19307 VDD.n3144 VDD.n3143 99.5127
R19308 VDD.n3148 VDD.n3147 99.5127
R19309 VDD.n3431 VDD.n637 99.5127
R19310 VDD.n3431 VDD.n627 99.5127
R19311 VDD.n3439 VDD.n627 99.5127
R19312 VDD.n3439 VDD.n625 99.5127
R19313 VDD.n3443 VDD.n625 99.5127
R19314 VDD.n3443 VDD.n615 99.5127
R19315 VDD.n3451 VDD.n615 99.5127
R19316 VDD.n3451 VDD.n613 99.5127
R19317 VDD.n3455 VDD.n613 99.5127
R19318 VDD.n3455 VDD.n603 99.5127
R19319 VDD.n3463 VDD.n603 99.5127
R19320 VDD.n3463 VDD.n601 99.5127
R19321 VDD.n3467 VDD.n601 99.5127
R19322 VDD.n3467 VDD.n592 99.5127
R19323 VDD.n3475 VDD.n592 99.5127
R19324 VDD.n3475 VDD.n590 99.5127
R19325 VDD.n3479 VDD.n590 99.5127
R19326 VDD.n3479 VDD.n580 99.5127
R19327 VDD.n3487 VDD.n580 99.5127
R19328 VDD.n3487 VDD.n578 99.5127
R19329 VDD.n3491 VDD.n578 99.5127
R19330 VDD.n3491 VDD.n568 99.5127
R19331 VDD.n3499 VDD.n568 99.5127
R19332 VDD.n3499 VDD.n566 99.5127
R19333 VDD.n3503 VDD.n566 99.5127
R19334 VDD.n3503 VDD.n556 99.5127
R19335 VDD.n3511 VDD.n556 99.5127
R19336 VDD.n3511 VDD.n554 99.5127
R19337 VDD.n3515 VDD.n554 99.5127
R19338 VDD.n3515 VDD.n544 99.5127
R19339 VDD.n3523 VDD.n544 99.5127
R19340 VDD.n3523 VDD.n542 99.5127
R19341 VDD.n3527 VDD.n542 99.5127
R19342 VDD.n3527 VDD.n532 99.5127
R19343 VDD.n3535 VDD.n532 99.5127
R19344 VDD.n3535 VDD.n530 99.5127
R19345 VDD.n3539 VDD.n530 99.5127
R19346 VDD.n3539 VDD.n520 99.5127
R19347 VDD.n3547 VDD.n520 99.5127
R19348 VDD.n3547 VDD.n518 99.5127
R19349 VDD.n3551 VDD.n518 99.5127
R19350 VDD.n3551 VDD.n508 99.5127
R19351 VDD.n3559 VDD.n508 99.5127
R19352 VDD.n3559 VDD.n506 99.5127
R19353 VDD.n3563 VDD.n506 99.5127
R19354 VDD.n3563 VDD.n496 99.5127
R19355 VDD.n3571 VDD.n496 99.5127
R19356 VDD.n3571 VDD.n494 99.5127
R19357 VDD.n3575 VDD.n494 99.5127
R19358 VDD.n3575 VDD.n484 99.5127
R19359 VDD.n3583 VDD.n484 99.5127
R19360 VDD.n3583 VDD.n482 99.5127
R19361 VDD.n3587 VDD.n482 99.5127
R19362 VDD.n3587 VDD.n472 99.5127
R19363 VDD.n3595 VDD.n472 99.5127
R19364 VDD.n3595 VDD.n470 99.5127
R19365 VDD.n3599 VDD.n470 99.5127
R19366 VDD.n3599 VDD.n460 99.5127
R19367 VDD.n3607 VDD.n460 99.5127
R19368 VDD.n3607 VDD.n458 99.5127
R19369 VDD.n3611 VDD.n458 99.5127
R19370 VDD.n3611 VDD.n448 99.5127
R19371 VDD.n3619 VDD.n448 99.5127
R19372 VDD.n3619 VDD.n446 99.5127
R19373 VDD.n3623 VDD.n446 99.5127
R19374 VDD.n3623 VDD.n436 99.5127
R19375 VDD.n3631 VDD.n436 99.5127
R19376 VDD.n3631 VDD.n434 99.5127
R19377 VDD.n3635 VDD.n434 99.5127
R19378 VDD.n3635 VDD.n424 99.5127
R19379 VDD.n3643 VDD.n424 99.5127
R19380 VDD.n3643 VDD.n422 99.5127
R19381 VDD.n3647 VDD.n422 99.5127
R19382 VDD.n3647 VDD.n413 99.5127
R19383 VDD.n3655 VDD.n413 99.5127
R19384 VDD.n3655 VDD.n411 99.5127
R19385 VDD.n3659 VDD.n411 99.5127
R19386 VDD.n3659 VDD.n401 99.5127
R19387 VDD.n3667 VDD.n401 99.5127
R19388 VDD.n3667 VDD.n399 99.5127
R19389 VDD.n3671 VDD.n399 99.5127
R19390 VDD.n3671 VDD.n389 99.5127
R19391 VDD.n3679 VDD.n389 99.5127
R19392 VDD.n3679 VDD.n387 99.5127
R19393 VDD.n3683 VDD.n387 99.5127
R19394 VDD.n3683 VDD.n377 99.5127
R19395 VDD.n3691 VDD.n377 99.5127
R19396 VDD.n3691 VDD.n375 99.5127
R19397 VDD.n3695 VDD.n375 99.5127
R19398 VDD.n3695 VDD.n365 99.5127
R19399 VDD.n3703 VDD.n365 99.5127
R19400 VDD.n3703 VDD.n363 99.5127
R19401 VDD.n3707 VDD.n363 99.5127
R19402 VDD.n3707 VDD.n353 99.5127
R19403 VDD.n3715 VDD.n353 99.5127
R19404 VDD.n3715 VDD.n351 99.5127
R19405 VDD.n3719 VDD.n351 99.5127
R19406 VDD.n3719 VDD.n341 99.5127
R19407 VDD.n3727 VDD.n341 99.5127
R19408 VDD.n3727 VDD.n339 99.5127
R19409 VDD.n3731 VDD.n339 99.5127
R19410 VDD.n3731 VDD.n329 99.5127
R19411 VDD.n3739 VDD.n329 99.5127
R19412 VDD.n3739 VDD.n327 99.5127
R19413 VDD.n3743 VDD.n327 99.5127
R19414 VDD.n3743 VDD.n317 99.5127
R19415 VDD.n3751 VDD.n317 99.5127
R19416 VDD.n3751 VDD.n315 99.5127
R19417 VDD.n3755 VDD.n315 99.5127
R19418 VDD.n3755 VDD.n305 99.5127
R19419 VDD.n3763 VDD.n305 99.5127
R19420 VDD.n3763 VDD.n303 99.5127
R19421 VDD.n3767 VDD.n303 99.5127
R19422 VDD.n3767 VDD.n293 99.5127
R19423 VDD.n3775 VDD.n293 99.5127
R19424 VDD.n3775 VDD.n291 99.5127
R19425 VDD.n3779 VDD.n291 99.5127
R19426 VDD.n3779 VDD.n281 99.5127
R19427 VDD.n3787 VDD.n281 99.5127
R19428 VDD.n3787 VDD.n279 99.5127
R19429 VDD.n3791 VDD.n279 99.5127
R19430 VDD.n3791 VDD.n269 99.5127
R19431 VDD.n3799 VDD.n269 99.5127
R19432 VDD.n3799 VDD.n267 99.5127
R19433 VDD.n3803 VDD.n267 99.5127
R19434 VDD.n3803 VDD.n257 99.5127
R19435 VDD.n3811 VDD.n257 99.5127
R19436 VDD.n3811 VDD.n255 99.5127
R19437 VDD.n3815 VDD.n255 99.5127
R19438 VDD.n3815 VDD.n245 99.5127
R19439 VDD.n3823 VDD.n245 99.5127
R19440 VDD.n3823 VDD.n243 99.5127
R19441 VDD.n3827 VDD.n243 99.5127
R19442 VDD.n3827 VDD.n232 99.5127
R19443 VDD.n3835 VDD.n232 99.5127
R19444 VDD.n3835 VDD.n230 99.5127
R19445 VDD.n3839 VDD.n230 99.5127
R19446 VDD.n3839 VDD.n221 99.5127
R19447 VDD.n3847 VDD.n221 99.5127
R19448 VDD.n3847 VDD.n218 99.5127
R19449 VDD.n3877 VDD.n218 99.5127
R19450 VDD.n3877 VDD.n219 99.5127
R19451 VDD.n219 VDD.n211 99.5127
R19452 VDD.n3872 VDD.n211 99.5127
R19453 VDD.n3872 VDD.n188 99.5127
R19454 VDD.n2901 VDD.n660 99.5127
R19455 VDD.n2897 VDD.n2896 99.5127
R19456 VDD.n2893 VDD.n2892 99.5127
R19457 VDD.n2889 VDD.n2888 99.5127
R19458 VDD.n2885 VDD.n2884 99.5127
R19459 VDD.n2881 VDD.n2880 99.5127
R19460 VDD.n2877 VDD.n2876 99.5127
R19461 VDD.n2872 VDD.n2871 99.5127
R19462 VDD.n2868 VDD.n658 99.5127
R19463 VDD.n2346 VDD.n1104 99.5127
R19464 VDD.n2346 VDD.n1098 99.5127
R19465 VDD.n2343 VDD.n1098 99.5127
R19466 VDD.n2343 VDD.n1092 99.5127
R19467 VDD.n2340 VDD.n1092 99.5127
R19468 VDD.n2340 VDD.n1086 99.5127
R19469 VDD.n2337 VDD.n1086 99.5127
R19470 VDD.n2337 VDD.n1080 99.5127
R19471 VDD.n2334 VDD.n1080 99.5127
R19472 VDD.n2334 VDD.n1073 99.5127
R19473 VDD.n2331 VDD.n1073 99.5127
R19474 VDD.n2331 VDD.n1067 99.5127
R19475 VDD.n2328 VDD.n1067 99.5127
R19476 VDD.n2328 VDD.n1062 99.5127
R19477 VDD.n2325 VDD.n1062 99.5127
R19478 VDD.n2325 VDD.n1056 99.5127
R19479 VDD.n2322 VDD.n1056 99.5127
R19480 VDD.n2322 VDD.n1050 99.5127
R19481 VDD.n2319 VDD.n1050 99.5127
R19482 VDD.n2319 VDD.n1044 99.5127
R19483 VDD.n2316 VDD.n1044 99.5127
R19484 VDD.n2316 VDD.n1038 99.5127
R19485 VDD.n2313 VDD.n1038 99.5127
R19486 VDD.n2313 VDD.n1032 99.5127
R19487 VDD.n2310 VDD.n1032 99.5127
R19488 VDD.n2310 VDD.n1025 99.5127
R19489 VDD.n2307 VDD.n1025 99.5127
R19490 VDD.n2307 VDD.n1019 99.5127
R19491 VDD.n2304 VDD.n1019 99.5127
R19492 VDD.n2304 VDD.n1014 99.5127
R19493 VDD.n2301 VDD.n1014 99.5127
R19494 VDD.n2301 VDD.n1008 99.5127
R19495 VDD.n2298 VDD.n1008 99.5127
R19496 VDD.n2298 VDD.n1002 99.5127
R19497 VDD.n2295 VDD.n1002 99.5127
R19498 VDD.n2295 VDD.n996 99.5127
R19499 VDD.n2292 VDD.n996 99.5127
R19500 VDD.n2292 VDD.n990 99.5127
R19501 VDD.n2289 VDD.n990 99.5127
R19502 VDD.n2289 VDD.n984 99.5127
R19503 VDD.n2286 VDD.n984 99.5127
R19504 VDD.n2286 VDD.n978 99.5127
R19505 VDD.n2283 VDD.n978 99.5127
R19506 VDD.n2283 VDD.n972 99.5127
R19507 VDD.n2280 VDD.n972 99.5127
R19508 VDD.n2280 VDD.n966 99.5127
R19509 VDD.n2277 VDD.n966 99.5127
R19510 VDD.n2277 VDD.n960 99.5127
R19511 VDD.n2274 VDD.n960 99.5127
R19512 VDD.n2274 VDD.n954 99.5127
R19513 VDD.n2271 VDD.n954 99.5127
R19514 VDD.n2271 VDD.n947 99.5127
R19515 VDD.n2268 VDD.n947 99.5127
R19516 VDD.n2268 VDD.n941 99.5127
R19517 VDD.n2265 VDD.n941 99.5127
R19518 VDD.n2265 VDD.n936 99.5127
R19519 VDD.n2262 VDD.n936 99.5127
R19520 VDD.n2262 VDD.n930 99.5127
R19521 VDD.n2259 VDD.n930 99.5127
R19522 VDD.n2259 VDD.n924 99.5127
R19523 VDD.n2256 VDD.n924 99.5127
R19524 VDD.n2256 VDD.n918 99.5127
R19525 VDD.n2253 VDD.n918 99.5127
R19526 VDD.n2253 VDD.n912 99.5127
R19527 VDD.n2250 VDD.n912 99.5127
R19528 VDD.n2250 VDD.n906 99.5127
R19529 VDD.n2247 VDD.n906 99.5127
R19530 VDD.n2247 VDD.n900 99.5127
R19531 VDD.n2244 VDD.n900 99.5127
R19532 VDD.n2244 VDD.n894 99.5127
R19533 VDD.n2241 VDD.n894 99.5127
R19534 VDD.n2241 VDD.n888 99.5127
R19535 VDD.n2238 VDD.n888 99.5127
R19536 VDD.n2238 VDD.n882 99.5127
R19537 VDD.n2235 VDD.n882 99.5127
R19538 VDD.n2235 VDD.n876 99.5127
R19539 VDD.n2232 VDD.n876 99.5127
R19540 VDD.n2232 VDD.n871 99.5127
R19541 VDD.n2229 VDD.n871 99.5127
R19542 VDD.n2229 VDD.n865 99.5127
R19543 VDD.n2226 VDD.n865 99.5127
R19544 VDD.n2226 VDD.n859 99.5127
R19545 VDD.n2223 VDD.n859 99.5127
R19546 VDD.n2223 VDD.n853 99.5127
R19547 VDD.n2220 VDD.n853 99.5127
R19548 VDD.n2220 VDD.n847 99.5127
R19549 VDD.n2217 VDD.n847 99.5127
R19550 VDD.n2217 VDD.n841 99.5127
R19551 VDD.n2214 VDD.n841 99.5127
R19552 VDD.n2214 VDD.n834 99.5127
R19553 VDD.n2211 VDD.n834 99.5127
R19554 VDD.n2211 VDD.n828 99.5127
R19555 VDD.n2208 VDD.n828 99.5127
R19556 VDD.n2208 VDD.n823 99.5127
R19557 VDD.n2205 VDD.n823 99.5127
R19558 VDD.n2205 VDD.n817 99.5127
R19559 VDD.n2202 VDD.n817 99.5127
R19560 VDD.n2202 VDD.n811 99.5127
R19561 VDD.n2199 VDD.n811 99.5127
R19562 VDD.n2199 VDD.n805 99.5127
R19563 VDD.n2196 VDD.n805 99.5127
R19564 VDD.n2196 VDD.n799 99.5127
R19565 VDD.n2193 VDD.n799 99.5127
R19566 VDD.n2193 VDD.n793 99.5127
R19567 VDD.n2190 VDD.n793 99.5127
R19568 VDD.n2190 VDD.n787 99.5127
R19569 VDD.n2187 VDD.n787 99.5127
R19570 VDD.n2187 VDD.n781 99.5127
R19571 VDD.n2184 VDD.n781 99.5127
R19572 VDD.n2184 VDD.n775 99.5127
R19573 VDD.n2181 VDD.n775 99.5127
R19574 VDD.n2181 VDD.n768 99.5127
R19575 VDD.n2178 VDD.n768 99.5127
R19576 VDD.n2178 VDD.n762 99.5127
R19577 VDD.n2175 VDD.n762 99.5127
R19578 VDD.n2175 VDD.n757 99.5127
R19579 VDD.n2172 VDD.n757 99.5127
R19580 VDD.n2172 VDD.n751 99.5127
R19581 VDD.n2169 VDD.n751 99.5127
R19582 VDD.n2169 VDD.n745 99.5127
R19583 VDD.n2166 VDD.n745 99.5127
R19584 VDD.n2166 VDD.n739 99.5127
R19585 VDD.n2163 VDD.n739 99.5127
R19586 VDD.n2163 VDD.n733 99.5127
R19587 VDD.n2160 VDD.n733 99.5127
R19588 VDD.n2160 VDD.n727 99.5127
R19589 VDD.n2157 VDD.n727 99.5127
R19590 VDD.n2157 VDD.n721 99.5127
R19591 VDD.n2154 VDD.n721 99.5127
R19592 VDD.n2154 VDD.n715 99.5127
R19593 VDD.n2151 VDD.n715 99.5127
R19594 VDD.n2151 VDD.n709 99.5127
R19595 VDD.n2148 VDD.n709 99.5127
R19596 VDD.n2148 VDD.n703 99.5127
R19597 VDD.n1129 VDD.n703 99.5127
R19598 VDD.n1129 VDD.n698 99.5127
R19599 VDD.n1126 VDD.n698 99.5127
R19600 VDD.n1126 VDD.n692 99.5127
R19601 VDD.n1123 VDD.n692 99.5127
R19602 VDD.n1123 VDD.n685 99.5127
R19603 VDD.n1120 VDD.n685 99.5127
R19604 VDD.n1120 VDD.n678 99.5127
R19605 VDD.n678 VDD.n665 99.5127
R19606 VDD.n2864 VDD.n665 99.5127
R19607 VDD.n2865 VDD.n2864 99.5127
R19608 VDD.n2381 VDD.n1105 99.5127
R19609 VDD.n2379 VDD.n2378 99.5127
R19610 VDD.n2375 VDD.n2374 99.5127
R19611 VDD.n2372 VDD.n1109 99.5127
R19612 VDD.n2368 VDD.n2366 99.5127
R19613 VDD.n2363 VDD.n2362 99.5127
R19614 VDD.n2360 VDD.n1113 99.5127
R19615 VDD.n2355 VDD.n2353 99.5127
R19616 VDD.n2351 VDD.n1117 99.5127
R19617 VDD.n2385 VDD.n1095 99.5127
R19618 VDD.n2393 VDD.n1095 99.5127
R19619 VDD.n2393 VDD.n1093 99.5127
R19620 VDD.n2397 VDD.n1093 99.5127
R19621 VDD.n2397 VDD.n1083 99.5127
R19622 VDD.n2405 VDD.n1083 99.5127
R19623 VDD.n2405 VDD.n1081 99.5127
R19624 VDD.n2409 VDD.n1081 99.5127
R19625 VDD.n2409 VDD.n1070 99.5127
R19626 VDD.n2417 VDD.n1070 99.5127
R19627 VDD.n2417 VDD.n1068 99.5127
R19628 VDD.n2421 VDD.n1068 99.5127
R19629 VDD.n2421 VDD.n1059 99.5127
R19630 VDD.n2429 VDD.n1059 99.5127
R19631 VDD.n2429 VDD.n1057 99.5127
R19632 VDD.n2433 VDD.n1057 99.5127
R19633 VDD.n2433 VDD.n1047 99.5127
R19634 VDD.n2441 VDD.n1047 99.5127
R19635 VDD.n2441 VDD.n1045 99.5127
R19636 VDD.n2445 VDD.n1045 99.5127
R19637 VDD.n2445 VDD.n1035 99.5127
R19638 VDD.n2453 VDD.n1035 99.5127
R19639 VDD.n2453 VDD.n1033 99.5127
R19640 VDD.n2457 VDD.n1033 99.5127
R19641 VDD.n2457 VDD.n1022 99.5127
R19642 VDD.n2465 VDD.n1022 99.5127
R19643 VDD.n2465 VDD.n1020 99.5127
R19644 VDD.n2469 VDD.n1020 99.5127
R19645 VDD.n2469 VDD.n1011 99.5127
R19646 VDD.n2477 VDD.n1011 99.5127
R19647 VDD.n2477 VDD.n1009 99.5127
R19648 VDD.n2481 VDD.n1009 99.5127
R19649 VDD.n2481 VDD.n999 99.5127
R19650 VDD.n2489 VDD.n999 99.5127
R19651 VDD.n2489 VDD.n997 99.5127
R19652 VDD.n2493 VDD.n997 99.5127
R19653 VDD.n2493 VDD.n987 99.5127
R19654 VDD.n2501 VDD.n987 99.5127
R19655 VDD.n2501 VDD.n985 99.5127
R19656 VDD.n2505 VDD.n985 99.5127
R19657 VDD.n2505 VDD.n975 99.5127
R19658 VDD.n2513 VDD.n975 99.5127
R19659 VDD.n2513 VDD.n973 99.5127
R19660 VDD.n2517 VDD.n973 99.5127
R19661 VDD.n2517 VDD.n963 99.5127
R19662 VDD.n2525 VDD.n963 99.5127
R19663 VDD.n2525 VDD.n961 99.5127
R19664 VDD.n2529 VDD.n961 99.5127
R19665 VDD.n2529 VDD.n951 99.5127
R19666 VDD.n2537 VDD.n951 99.5127
R19667 VDD.n2537 VDD.n949 99.5127
R19668 VDD.n2541 VDD.n949 99.5127
R19669 VDD.n2541 VDD.n939 99.5127
R19670 VDD.n2549 VDD.n939 99.5127
R19671 VDD.n2549 VDD.n937 99.5127
R19672 VDD.n2553 VDD.n937 99.5127
R19673 VDD.n2553 VDD.n927 99.5127
R19674 VDD.n2561 VDD.n927 99.5127
R19675 VDD.n2561 VDD.n925 99.5127
R19676 VDD.n2565 VDD.n925 99.5127
R19677 VDD.n2565 VDD.n915 99.5127
R19678 VDD.n2573 VDD.n915 99.5127
R19679 VDD.n2573 VDD.n913 99.5127
R19680 VDD.n2577 VDD.n913 99.5127
R19681 VDD.n2577 VDD.n903 99.5127
R19682 VDD.n2585 VDD.n903 99.5127
R19683 VDD.n2585 VDD.n901 99.5127
R19684 VDD.n2589 VDD.n901 99.5127
R19685 VDD.n2589 VDD.n891 99.5127
R19686 VDD.n2597 VDD.n891 99.5127
R19687 VDD.n2597 VDD.n889 99.5127
R19688 VDD.n2601 VDD.n889 99.5127
R19689 VDD.n2601 VDD.n879 99.5127
R19690 VDD.n2609 VDD.n879 99.5127
R19691 VDD.n2609 VDD.n877 99.5127
R19692 VDD.n2613 VDD.n877 99.5127
R19693 VDD.n2613 VDD.n868 99.5127
R19694 VDD.n2621 VDD.n868 99.5127
R19695 VDD.n2621 VDD.n866 99.5127
R19696 VDD.n2625 VDD.n866 99.5127
R19697 VDD.n2625 VDD.n856 99.5127
R19698 VDD.n2633 VDD.n856 99.5127
R19699 VDD.n2633 VDD.n854 99.5127
R19700 VDD.n2637 VDD.n854 99.5127
R19701 VDD.n2637 VDD.n844 99.5127
R19702 VDD.n2645 VDD.n844 99.5127
R19703 VDD.n2645 VDD.n842 99.5127
R19704 VDD.n2649 VDD.n842 99.5127
R19705 VDD.n2649 VDD.n831 99.5127
R19706 VDD.n2657 VDD.n831 99.5127
R19707 VDD.n2657 VDD.n829 99.5127
R19708 VDD.n2661 VDD.n829 99.5127
R19709 VDD.n2661 VDD.n820 99.5127
R19710 VDD.n2669 VDD.n820 99.5127
R19711 VDD.n2669 VDD.n818 99.5127
R19712 VDD.n2673 VDD.n818 99.5127
R19713 VDD.n2673 VDD.n808 99.5127
R19714 VDD.n2681 VDD.n808 99.5127
R19715 VDD.n2681 VDD.n806 99.5127
R19716 VDD.n2685 VDD.n806 99.5127
R19717 VDD.n2685 VDD.n796 99.5127
R19718 VDD.n2693 VDD.n796 99.5127
R19719 VDD.n2693 VDD.n794 99.5127
R19720 VDD.n2697 VDD.n794 99.5127
R19721 VDD.n2697 VDD.n784 99.5127
R19722 VDD.n2705 VDD.n784 99.5127
R19723 VDD.n2705 VDD.n782 99.5127
R19724 VDD.n2709 VDD.n782 99.5127
R19725 VDD.n2709 VDD.n772 99.5127
R19726 VDD.n2717 VDD.n772 99.5127
R19727 VDD.n2717 VDD.n770 99.5127
R19728 VDD.n2721 VDD.n770 99.5127
R19729 VDD.n2721 VDD.n760 99.5127
R19730 VDD.n2729 VDD.n760 99.5127
R19731 VDD.n2729 VDD.n758 99.5127
R19732 VDD.n2733 VDD.n758 99.5127
R19733 VDD.n2733 VDD.n748 99.5127
R19734 VDD.n2741 VDD.n748 99.5127
R19735 VDD.n2741 VDD.n746 99.5127
R19736 VDD.n2745 VDD.n746 99.5127
R19737 VDD.n2745 VDD.n736 99.5127
R19738 VDD.n2753 VDD.n736 99.5127
R19739 VDD.n2753 VDD.n734 99.5127
R19740 VDD.n2757 VDD.n734 99.5127
R19741 VDD.n2757 VDD.n724 99.5127
R19742 VDD.n2765 VDD.n724 99.5127
R19743 VDD.n2765 VDD.n722 99.5127
R19744 VDD.n2769 VDD.n722 99.5127
R19745 VDD.n2769 VDD.n712 99.5127
R19746 VDD.n2777 VDD.n712 99.5127
R19747 VDD.n2777 VDD.n710 99.5127
R19748 VDD.n2781 VDD.n710 99.5127
R19749 VDD.n2781 VDD.n701 99.5127
R19750 VDD.n2789 VDD.n701 99.5127
R19751 VDD.n2789 VDD.n699 99.5127
R19752 VDD.n2793 VDD.n699 99.5127
R19753 VDD.n2793 VDD.n689 99.5127
R19754 VDD.n2801 VDD.n689 99.5127
R19755 VDD.n2801 VDD.n686 99.5127
R19756 VDD.n2810 VDD.n686 99.5127
R19757 VDD.n2810 VDD.n687 99.5127
R19758 VDD.n687 VDD.n679 99.5127
R19759 VDD.n2805 VDD.n679 99.5127
R19760 VDD.n2805 VDD.n668 99.5127
R19761 VDD.n668 VDD.n659 99.5127
R19762 VDD.t112 VDD.n1102 88.2921
R19763 VDD.n175 VDD.t105 88.2921
R19764 VDD.n3426 VDD.n3425 72.8958
R19765 VDD.n3425 VDD.n2918 72.8958
R19766 VDD.n3425 VDD.n2917 72.8958
R19767 VDD.n3425 VDD.n2916 72.8958
R19768 VDD.n3425 VDD.n2915 72.8958
R19769 VDD.n3425 VDD.n2914 72.8958
R19770 VDD.n3425 VDD.n2913 72.8958
R19771 VDD.n3425 VDD.n2912 72.8958
R19772 VDD.n3425 VDD.n2911 72.8958
R19773 VDD.n184 VDD.n175 72.8958
R19774 VDD.n3932 VDD.n175 72.8958
R19775 VDD.n180 VDD.n175 72.8958
R19776 VDD.n3939 VDD.n175 72.8958
R19777 VDD.n175 VDD.n174 72.8958
R19778 VDD.n3858 VDD.n175 72.8958
R19779 VDD.n3854 VDD.n175 72.8958
R19780 VDD.n3865 VDD.n175 72.8958
R19781 VDD.n3868 VDD.n175 72.8958
R19782 VDD.n1900 VDD.n1102 72.8958
R19783 VDD.n1906 VDD.n1102 72.8958
R19784 VDD.n1908 VDD.n1102 72.8958
R19785 VDD.n1914 VDD.n1102 72.8958
R19786 VDD.n1916 VDD.n1102 72.8958
R19787 VDD.n1922 VDD.n1102 72.8958
R19788 VDD.n1924 VDD.n1102 72.8958
R19789 VDD.n1931 VDD.n1102 72.8958
R19790 VDD.n2902 VDD.n649 72.8958
R19791 VDD.n2902 VDD.n648 72.8958
R19792 VDD.n2902 VDD.n647 72.8958
R19793 VDD.n2902 VDD.n646 72.8958
R19794 VDD.n2902 VDD.n645 72.8958
R19795 VDD.n2902 VDD.n644 72.8958
R19796 VDD.n2902 VDD.n643 72.8958
R19797 VDD.n2902 VDD.n642 72.8958
R19798 VDD.n2902 VDD.n641 72.8958
R19799 VDD.n3425 VDD.n3424 72.8958
R19800 VDD.n3425 VDD.n2903 72.8958
R19801 VDD.n3425 VDD.n2904 72.8958
R19802 VDD.n3425 VDD.n2905 72.8958
R19803 VDD.n3425 VDD.n2906 72.8958
R19804 VDD.n3425 VDD.n2907 72.8958
R19805 VDD.n3425 VDD.n2908 72.8958
R19806 VDD.n3425 VDD.n2909 72.8958
R19807 VDD.n3889 VDD.n175 72.8958
R19808 VDD.n3895 VDD.n175 72.8958
R19809 VDD.n204 VDD.n175 72.8958
R19810 VDD.n3902 VDD.n175 72.8958
R19811 VDD.n199 VDD.n175 72.8958
R19812 VDD.n3911 VDD.n175 72.8958
R19813 VDD.n196 VDD.n175 72.8958
R19814 VDD.n3918 VDD.n175 72.8958
R19815 VDD.n193 VDD.n175 72.8958
R19816 VDD.n2902 VDD.n657 72.8958
R19817 VDD.n2902 VDD.n656 72.8958
R19818 VDD.n2902 VDD.n655 72.8958
R19819 VDD.n2902 VDD.n654 72.8958
R19820 VDD.n2902 VDD.n653 72.8958
R19821 VDD.n2902 VDD.n652 72.8958
R19822 VDD.n2902 VDD.n651 72.8958
R19823 VDD.n2902 VDD.n650 72.8958
R19824 VDD.n2380 VDD.n1102 72.8958
R19825 VDD.n1107 VDD.n1102 72.8958
R19826 VDD.n2373 VDD.n1102 72.8958
R19827 VDD.n2367 VDD.n1102 72.8958
R19828 VDD.n1111 VDD.n1102 72.8958
R19829 VDD.n2361 VDD.n1102 72.8958
R19830 VDD.n2354 VDD.n1102 72.8958
R19831 VDD.n2352 VDD.n1102 72.8958
R19832 VDD.n1449 VDD.n1372 66.2847
R19833 VDD.n1452 VDD.n1372 66.2847
R19834 VDD.n1462 VDD.n1372 66.2847
R19835 VDD.n1465 VDD.n1372 66.2847
R19836 VDD.n1436 VDD.n1372 66.2847
R19837 VDD.n1474 VDD.n1372 66.2847
R19838 VDD.n1476 VDD.n1372 66.2847
R19839 VDD.n1485 VDD.n1372 66.2847
R19840 VDD.n1488 VDD.n1372 66.2847
R19841 VDD.n1426 VDD.n1372 66.2847
R19842 VDD.n1497 VDD.n1372 66.2847
R19843 VDD.n1499 VDD.n1372 66.2847
R19844 VDD.n1507 VDD.n1372 66.2847
R19845 VDD.n1509 VDD.n1372 66.2847
R19846 VDD.n1519 VDD.n1372 66.2847
R19847 VDD.n1522 VDD.n1372 66.2847
R19848 VDD.n1405 VDD.n1372 66.2847
R19849 VDD.n1531 VDD.n1372 66.2847
R19850 VDD.n1533 VDD.n1372 66.2847
R19851 VDD.n1541 VDD.n1372 66.2847
R19852 VDD.n1543 VDD.n1372 66.2847
R19853 VDD.n1551 VDD.n1372 66.2847
R19854 VDD.n1553 VDD.n1372 66.2847
R19855 VDD.n1561 VDD.n1372 66.2847
R19856 VDD.n1563 VDD.n1372 66.2847
R19857 VDD.n1571 VDD.n1372 66.2847
R19858 VDD.n1574 VDD.n1372 66.2847
R19859 VDD.n1379 VDD.n1372 66.2847
R19860 VDD.n1807 VDD.n1146 66.2847
R19861 VDD.n1227 VDD.n1146 66.2847
R19862 VDD.n1219 VDD.n1146 66.2847
R19863 VDD.n1216 VDD.n1146 66.2847
R19864 VDD.n1211 VDD.n1146 66.2847
R19865 VDD.n1208 VDD.n1146 66.2847
R19866 VDD.n1827 VDD.n1146 66.2847
R19867 VDD.n1200 VDD.n1146 66.2847
R19868 VDD.n1834 VDD.n1146 66.2847
R19869 VDD.n1193 VDD.n1146 66.2847
R19870 VDD.n1841 VDD.n1146 66.2847
R19871 VDD.n1187 VDD.n1146 66.2847
R19872 VDD.n1850 VDD.n1146 66.2847
R19873 VDD.n1179 VDD.n1146 66.2847
R19874 VDD.n1857 VDD.n1146 66.2847
R19875 VDD.n1172 VDD.n1146 66.2847
R19876 VDD.n1864 VDD.n1146 66.2847
R19877 VDD.n1166 VDD.n1146 66.2847
R19878 VDD.n1873 VDD.n1146 66.2847
R19879 VDD.n1158 VDD.n1146 66.2847
R19880 VDD.n1880 VDD.n1146 66.2847
R19881 VDD.n1151 VDD.n1146 66.2847
R19882 VDD.n1887 VDD.n1146 66.2847
R19883 VDD.n1890 VDD.n1146 66.2847
R19884 VDD.n1785 VDD.n1146 66.2847
R19885 VDD.n1784 VDD.n1146 66.2847
R19886 VDD.n1792 VDD.n1146 66.2847
R19887 VDD.n1795 VDD.n1146 66.2847
R19888 VDD.n1771 VDD.n1146 66.2847
R19889 VDD.n4075 VDD.n4074 66.2847
R19890 VDD.n4074 VDD.n100 66.2847
R19891 VDD.n4074 VDD.n101 66.2847
R19892 VDD.n4074 VDD.n102 66.2847
R19893 VDD.n4074 VDD.n103 66.2847
R19894 VDD.n4074 VDD.n104 66.2847
R19895 VDD.n4074 VDD.n105 66.2847
R19896 VDD.n4074 VDD.n106 66.2847
R19897 VDD.n4074 VDD.n107 66.2847
R19898 VDD.n4074 VDD.n108 66.2847
R19899 VDD.n4074 VDD.n109 66.2847
R19900 VDD.n4074 VDD.n110 66.2847
R19901 VDD.n4074 VDD.n111 66.2847
R19902 VDD.n4074 VDD.n112 66.2847
R19903 VDD.n4074 VDD.n113 66.2847
R19904 VDD.n4074 VDD.n114 66.2847
R19905 VDD.n4074 VDD.n115 66.2847
R19906 VDD.n4074 VDD.n116 66.2847
R19907 VDD.n4074 VDD.n117 66.2847
R19908 VDD.n4074 VDD.n118 66.2847
R19909 VDD.n4074 VDD.n119 66.2847
R19910 VDD.n4074 VDD.n120 66.2847
R19911 VDD.n4074 VDD.n121 66.2847
R19912 VDD.n4074 VDD.n122 66.2847
R19913 VDD.n4074 VDD.n123 66.2847
R19914 VDD.n4074 VDD.n124 66.2847
R19915 VDD.n4074 VDD.n125 66.2847
R19916 VDD.n4074 VDD.n126 66.2847
R19917 VDD.n4381 VDD.n4264 66.2847
R19918 VDD.n4366 VDD.n4264 66.2847
R19919 VDD.n4388 VDD.n4264 66.2847
R19920 VDD.n4357 VDD.n4264 66.2847
R19921 VDD.n4395 VDD.n4264 66.2847
R19922 VDD.n4350 VDD.n4264 66.2847
R19923 VDD.n4402 VDD.n4264 66.2847
R19924 VDD.n4340 VDD.n4264 66.2847
R19925 VDD.n4409 VDD.n4264 66.2847
R19926 VDD.n4333 VDD.n4264 66.2847
R19927 VDD.n4416 VDD.n4264 66.2847
R19928 VDD.n4327 VDD.n4264 66.2847
R19929 VDD.n4425 VDD.n4264 66.2847
R19930 VDD.n4319 VDD.n4264 66.2847
R19931 VDD.n4432 VDD.n4264 66.2847
R19932 VDD.n4312 VDD.n4264 66.2847
R19933 VDD.n4439 VDD.n4264 66.2847
R19934 VDD.n4306 VDD.n4264 66.2847
R19935 VDD.n4448 VDD.n4264 66.2847
R19936 VDD.n4298 VDD.n4264 66.2847
R19937 VDD.n4455 VDD.n4264 66.2847
R19938 VDD.n4291 VDD.n4264 66.2847
R19939 VDD.n4462 VDD.n4264 66.2847
R19940 VDD.n4285 VDD.n4264 66.2847
R19941 VDD.n4280 VDD.n4264 66.2847
R19942 VDD.n4473 VDD.n4264 66.2847
R19943 VDD.n4272 VDD.n4264 66.2847
R19944 VDD.n4480 VDD.n4264 66.2847
R19945 VDD.n4483 VDD.n4264 66.2847
R19946 VDD.n4483 VDD.n4482 52.4337
R19947 VDD.n4480 VDD.n4479 52.4337
R19948 VDD.n4475 VDD.n4272 52.4337
R19949 VDD.n4473 VDD.n4472 52.4337
R19950 VDD.n4281 VDD.n4280 52.4337
R19951 VDD.n4464 VDD.n4285 52.4337
R19952 VDD.n4462 VDD.n4461 52.4337
R19953 VDD.n4457 VDD.n4291 52.4337
R19954 VDD.n4455 VDD.n4454 52.4337
R19955 VDD.n4450 VDD.n4298 52.4337
R19956 VDD.n4448 VDD.n4447 52.4337
R19957 VDD.n4441 VDD.n4306 52.4337
R19958 VDD.n4439 VDD.n4438 52.4337
R19959 VDD.n4434 VDD.n4312 52.4337
R19960 VDD.n4432 VDD.n4431 52.4337
R19961 VDD.n4427 VDD.n4319 52.4337
R19962 VDD.n4425 VDD.n4424 52.4337
R19963 VDD.n4418 VDD.n4327 52.4337
R19964 VDD.n4416 VDD.n4415 52.4337
R19965 VDD.n4411 VDD.n4333 52.4337
R19966 VDD.n4409 VDD.n4408 52.4337
R19967 VDD.n4404 VDD.n4340 52.4337
R19968 VDD.n4402 VDD.n4401 52.4337
R19969 VDD.n4397 VDD.n4350 52.4337
R19970 VDD.n4395 VDD.n4394 52.4337
R19971 VDD.n4390 VDD.n4357 52.4337
R19972 VDD.n4388 VDD.n4387 52.4337
R19973 VDD.n4383 VDD.n4366 52.4337
R19974 VDD.n4381 VDD.n4380 52.4337
R19975 VDD.n4076 VDD.n4075 52.4337
R19976 VDD.n128 VDD.n100 52.4337
R19977 VDD.n4068 VDD.n101 52.4337
R19978 VDD.n4064 VDD.n102 52.4337
R19979 VDD.n4060 VDD.n103 52.4337
R19980 VDD.n4056 VDD.n104 52.4337
R19981 VDD.n4052 VDD.n105 52.4337
R19982 VDD.n4048 VDD.n106 52.4337
R19983 VDD.n4044 VDD.n107 52.4337
R19984 VDD.n4040 VDD.n108 52.4337
R19985 VDD.n4036 VDD.n109 52.4337
R19986 VDD.n4028 VDD.n110 52.4337
R19987 VDD.n4024 VDD.n111 52.4337
R19988 VDD.n4020 VDD.n112 52.4337
R19989 VDD.n4016 VDD.n113 52.4337
R19990 VDD.n4012 VDD.n114 52.4337
R19991 VDD.n4008 VDD.n115 52.4337
R19992 VDD.n4004 VDD.n116 52.4337
R19993 VDD.n4000 VDD.n117 52.4337
R19994 VDD.n3996 VDD.n118 52.4337
R19995 VDD.n3992 VDD.n119 52.4337
R19996 VDD.n3988 VDD.n120 52.4337
R19997 VDD.n3948 VDD.n121 52.4337
R19998 VDD.n3952 VDD.n122 52.4337
R19999 VDD.n3980 VDD.n123 52.4337
R20000 VDD.n3976 VDD.n124 52.4337
R20001 VDD.n3972 VDD.n125 52.4337
R20002 VDD.n3968 VDD.n126 52.4337
R20003 VDD.n1772 VDD.n1771 52.4337
R20004 VDD.n1795 VDD.n1794 52.4337
R20005 VDD.n1792 VDD.n1791 52.4337
R20006 VDD.n1787 VDD.n1784 52.4337
R20007 VDD.n1785 VDD.n1145 52.4337
R20008 VDD.n1890 VDD.n1889 52.4337
R20009 VDD.n1887 VDD.n1886 52.4337
R20010 VDD.n1882 VDD.n1151 52.4337
R20011 VDD.n1880 VDD.n1879 52.4337
R20012 VDD.n1875 VDD.n1158 52.4337
R20013 VDD.n1873 VDD.n1872 52.4337
R20014 VDD.n1866 VDD.n1166 52.4337
R20015 VDD.n1864 VDD.n1863 52.4337
R20016 VDD.n1859 VDD.n1172 52.4337
R20017 VDD.n1857 VDD.n1856 52.4337
R20018 VDD.n1852 VDD.n1179 52.4337
R20019 VDD.n1850 VDD.n1849 52.4337
R20020 VDD.n1843 VDD.n1187 52.4337
R20021 VDD.n1841 VDD.n1840 52.4337
R20022 VDD.n1836 VDD.n1193 52.4337
R20023 VDD.n1834 VDD.n1833 52.4337
R20024 VDD.n1829 VDD.n1200 52.4337
R20025 VDD.n1827 VDD.n1826 52.4337
R20026 VDD.n1209 VDD.n1208 52.4337
R20027 VDD.n1212 VDD.n1211 52.4337
R20028 VDD.n1217 VDD.n1216 52.4337
R20029 VDD.n1220 VDD.n1219 52.4337
R20030 VDD.n1228 VDD.n1227 52.4337
R20031 VDD.n1807 VDD.n1806 52.4337
R20032 VDD.n1449 VDD.n1371 52.4337
R20033 VDD.n1453 VDD.n1452 52.4337
R20034 VDD.n1462 VDD.n1461 52.4337
R20035 VDD.n1465 VDD.n1464 52.4337
R20036 VDD.n1437 VDD.n1436 52.4337
R20037 VDD.n1474 VDD.n1473 52.4337
R20038 VDD.n1477 VDD.n1476 52.4337
R20039 VDD.n1485 VDD.n1484 52.4337
R20040 VDD.n1488 VDD.n1487 52.4337
R20041 VDD.n1427 VDD.n1426 52.4337
R20042 VDD.n1497 VDD.n1496 52.4337
R20043 VDD.n1500 VDD.n1499 52.4337
R20044 VDD.n1507 VDD.n1506 52.4337
R20045 VDD.n1510 VDD.n1509 52.4337
R20046 VDD.n1519 VDD.n1518 52.4337
R20047 VDD.n1522 VDD.n1521 52.4337
R20048 VDD.n1406 VDD.n1405 52.4337
R20049 VDD.n1531 VDD.n1530 52.4337
R20050 VDD.n1534 VDD.n1533 52.4337
R20051 VDD.n1541 VDD.n1540 52.4337
R20052 VDD.n1544 VDD.n1543 52.4337
R20053 VDD.n1551 VDD.n1550 52.4337
R20054 VDD.n1554 VDD.n1553 52.4337
R20055 VDD.n1561 VDD.n1560 52.4337
R20056 VDD.n1564 VDD.n1563 52.4337
R20057 VDD.n1571 VDD.n1570 52.4337
R20058 VDD.n1575 VDD.n1574 52.4337
R20059 VDD.n1380 VDD.n1379 52.4337
R20060 VDD.n1450 VDD.n1449 52.4337
R20061 VDD.n1452 VDD.n1442 52.4337
R20062 VDD.n1463 VDD.n1462 52.4337
R20063 VDD.n1466 VDD.n1465 52.4337
R20064 VDD.n1436 VDD.n1433 52.4337
R20065 VDD.n1475 VDD.n1474 52.4337
R20066 VDD.n1476 VDD.n1429 52.4337
R20067 VDD.n1486 VDD.n1485 52.4337
R20068 VDD.n1489 VDD.n1488 52.4337
R20069 VDD.n1426 VDD.n1419 52.4337
R20070 VDD.n1498 VDD.n1497 52.4337
R20071 VDD.n1499 VDD.n1415 52.4337
R20072 VDD.n1508 VDD.n1507 52.4337
R20073 VDD.n1509 VDD.n1411 52.4337
R20074 VDD.n1520 VDD.n1519 52.4337
R20075 VDD.n1523 VDD.n1522 52.4337
R20076 VDD.n1405 VDD.n1402 52.4337
R20077 VDD.n1532 VDD.n1531 52.4337
R20078 VDD.n1533 VDD.n1398 52.4337
R20079 VDD.n1542 VDD.n1541 52.4337
R20080 VDD.n1543 VDD.n1394 52.4337
R20081 VDD.n1552 VDD.n1551 52.4337
R20082 VDD.n1553 VDD.n1387 52.4337
R20083 VDD.n1562 VDD.n1561 52.4337
R20084 VDD.n1563 VDD.n1383 52.4337
R20085 VDD.n1572 VDD.n1571 52.4337
R20086 VDD.n1574 VDD.n1573 52.4337
R20087 VDD.n1379 VDD.n1375 52.4337
R20088 VDD.n1808 VDD.n1807 52.4337
R20089 VDD.n1227 VDD.n1221 52.4337
R20090 VDD.n1219 VDD.n1218 52.4337
R20091 VDD.n1216 VDD.n1213 52.4337
R20092 VDD.n1211 VDD.n1210 52.4337
R20093 VDD.n1208 VDD.n1201 52.4337
R20094 VDD.n1828 VDD.n1827 52.4337
R20095 VDD.n1200 VDD.n1194 52.4337
R20096 VDD.n1835 VDD.n1834 52.4337
R20097 VDD.n1193 VDD.n1188 52.4337
R20098 VDD.n1842 VDD.n1841 52.4337
R20099 VDD.n1187 VDD.n1180 52.4337
R20100 VDD.n1851 VDD.n1850 52.4337
R20101 VDD.n1179 VDD.n1173 52.4337
R20102 VDD.n1858 VDD.n1857 52.4337
R20103 VDD.n1172 VDD.n1167 52.4337
R20104 VDD.n1865 VDD.n1864 52.4337
R20105 VDD.n1166 VDD.n1159 52.4337
R20106 VDD.n1874 VDD.n1873 52.4337
R20107 VDD.n1158 VDD.n1152 52.4337
R20108 VDD.n1881 VDD.n1880 52.4337
R20109 VDD.n1151 VDD.n1148 52.4337
R20110 VDD.n1888 VDD.n1887 52.4337
R20111 VDD.n1891 VDD.n1890 52.4337
R20112 VDD.n1786 VDD.n1785 52.4337
R20113 VDD.n1784 VDD.n1776 52.4337
R20114 VDD.n1793 VDD.n1792 52.4337
R20115 VDD.n1796 VDD.n1795 52.4337
R20116 VDD.n1771 VDD.n1233 52.4337
R20117 VDD.n4075 VDD.n99 52.4337
R20118 VDD.n4069 VDD.n100 52.4337
R20119 VDD.n4065 VDD.n101 52.4337
R20120 VDD.n4061 VDD.n102 52.4337
R20121 VDD.n4057 VDD.n103 52.4337
R20122 VDD.n4053 VDD.n104 52.4337
R20123 VDD.n4049 VDD.n105 52.4337
R20124 VDD.n4045 VDD.n106 52.4337
R20125 VDD.n4041 VDD.n107 52.4337
R20126 VDD.n4037 VDD.n108 52.4337
R20127 VDD.n4027 VDD.n109 52.4337
R20128 VDD.n4025 VDD.n110 52.4337
R20129 VDD.n4021 VDD.n111 52.4337
R20130 VDD.n4017 VDD.n112 52.4337
R20131 VDD.n4013 VDD.n113 52.4337
R20132 VDD.n4009 VDD.n114 52.4337
R20133 VDD.n4005 VDD.n115 52.4337
R20134 VDD.n4001 VDD.n116 52.4337
R20135 VDD.n3997 VDD.n117 52.4337
R20136 VDD.n3993 VDD.n118 52.4337
R20137 VDD.n3989 VDD.n119 52.4337
R20138 VDD.n3947 VDD.n120 52.4337
R20139 VDD.n3951 VDD.n121 52.4337
R20140 VDD.n3981 VDD.n122 52.4337
R20141 VDD.n3977 VDD.n123 52.4337
R20142 VDD.n3973 VDD.n124 52.4337
R20143 VDD.n3969 VDD.n125 52.4337
R20144 VDD.n3961 VDD.n126 52.4337
R20145 VDD.n4382 VDD.n4381 52.4337
R20146 VDD.n4366 VDD.n4358 52.4337
R20147 VDD.n4389 VDD.n4388 52.4337
R20148 VDD.n4357 VDD.n4351 52.4337
R20149 VDD.n4396 VDD.n4395 52.4337
R20150 VDD.n4350 VDD.n4341 52.4337
R20151 VDD.n4403 VDD.n4402 52.4337
R20152 VDD.n4340 VDD.n4334 52.4337
R20153 VDD.n4410 VDD.n4409 52.4337
R20154 VDD.n4333 VDD.n4328 52.4337
R20155 VDD.n4417 VDD.n4416 52.4337
R20156 VDD.n4327 VDD.n4320 52.4337
R20157 VDD.n4426 VDD.n4425 52.4337
R20158 VDD.n4319 VDD.n4313 52.4337
R20159 VDD.n4433 VDD.n4432 52.4337
R20160 VDD.n4312 VDD.n4307 52.4337
R20161 VDD.n4440 VDD.n4439 52.4337
R20162 VDD.n4306 VDD.n4299 52.4337
R20163 VDD.n4449 VDD.n4448 52.4337
R20164 VDD.n4298 VDD.n4292 52.4337
R20165 VDD.n4456 VDD.n4455 52.4337
R20166 VDD.n4291 VDD.n4286 52.4337
R20167 VDD.n4463 VDD.n4462 52.4337
R20168 VDD.n4285 VDD.n4284 52.4337
R20169 VDD.n4280 VDD.n4273 52.4337
R20170 VDD.n4474 VDD.n4473 52.4337
R20171 VDD.n4272 VDD.n4266 52.4337
R20172 VDD.n4481 VDD.n4480 52.4337
R20173 VDD.n4484 VDD.n4483 52.4337
R20174 VDD.n3920 VDD.n193 39.2114
R20175 VDD.n3918 VDD.n3917 39.2114
R20176 VDD.n3913 VDD.n196 39.2114
R20177 VDD.n3911 VDD.n3910 39.2114
R20178 VDD.n3904 VDD.n199 39.2114
R20179 VDD.n3902 VDD.n3901 39.2114
R20180 VDD.n3897 VDD.n204 39.2114
R20181 VDD.n3895 VDD.n3894 39.2114
R20182 VDD.n3890 VDD.n3889 39.2114
R20183 VDD.n3424 VDD.n3423 39.2114
R20184 VDD.n3418 VDD.n2903 39.2114
R20185 VDD.n3415 VDD.n2904 39.2114
R20186 VDD.n3411 VDD.n2905 39.2114
R20187 VDD.n3407 VDD.n2906 39.2114
R20188 VDD.n3403 VDD.n2907 39.2114
R20189 VDD.n3399 VDD.n2908 39.2114
R20190 VDD.n3394 VDD.n2909 39.2114
R20191 VDD.n2856 VDD.n641 39.2114
R20192 VDD.n2852 VDD.n642 39.2114
R20193 VDD.n2848 VDD.n643 39.2114
R20194 VDD.n2844 VDD.n644 39.2114
R20195 VDD.n2840 VDD.n645 39.2114
R20196 VDD.n2836 VDD.n646 39.2114
R20197 VDD.n2832 VDD.n647 39.2114
R20198 VDD.n2828 VDD.n648 39.2114
R20199 VDD.n2824 VDD.n649 39.2114
R20200 VDD.n1900 VDD.n1101 39.2114
R20201 VDD.n1906 VDD.n1905 39.2114
R20202 VDD.n1909 VDD.n1908 39.2114
R20203 VDD.n1914 VDD.n1913 39.2114
R20204 VDD.n1917 VDD.n1916 39.2114
R20205 VDD.n1922 VDD.n1921 39.2114
R20206 VDD.n1925 VDD.n1924 39.2114
R20207 VDD.n1931 VDD.n1930 39.2114
R20208 VDD.n3868 VDD.n3867 39.2114
R20209 VDD.n3865 VDD.n3864 39.2114
R20210 VDD.n3860 VDD.n3854 39.2114
R20211 VDD.n3858 VDD.n3857 39.2114
R20212 VDD.n3941 VDD.n174 39.2114
R20213 VDD.n3939 VDD.n3938 39.2114
R20214 VDD.n3934 VDD.n180 39.2114
R20215 VDD.n3932 VDD.n3931 39.2114
R20216 VDD.n3927 VDD.n184 39.2114
R20217 VDD.n3427 VDD.n3426 39.2114
R20218 VDD.n3120 VDD.n2918 39.2114
R20219 VDD.n3124 VDD.n2917 39.2114
R20220 VDD.n3128 VDD.n2916 39.2114
R20221 VDD.n3132 VDD.n2915 39.2114
R20222 VDD.n3136 VDD.n2914 39.2114
R20223 VDD.n3140 VDD.n2913 39.2114
R20224 VDD.n3144 VDD.n2912 39.2114
R20225 VDD.n3148 VDD.n2911 39.2114
R20226 VDD.n3426 VDD.n639 39.2114
R20227 VDD.n3123 VDD.n2918 39.2114
R20228 VDD.n3127 VDD.n2917 39.2114
R20229 VDD.n3131 VDD.n2916 39.2114
R20230 VDD.n3135 VDD.n2915 39.2114
R20231 VDD.n3139 VDD.n2914 39.2114
R20232 VDD.n3143 VDD.n2913 39.2114
R20233 VDD.n3147 VDD.n2912 39.2114
R20234 VDD.n3151 VDD.n2911 39.2114
R20235 VDD.n184 VDD.n182 39.2114
R20236 VDD.n3933 VDD.n3932 39.2114
R20237 VDD.n180 VDD.n176 39.2114
R20238 VDD.n3940 VDD.n3939 39.2114
R20239 VDD.n3855 VDD.n174 39.2114
R20240 VDD.n3859 VDD.n3858 39.2114
R20241 VDD.n3854 VDD.n3852 39.2114
R20242 VDD.n3866 VDD.n3865 39.2114
R20243 VDD.n3869 VDD.n3868 39.2114
R20244 VDD.n1901 VDD.n1900 39.2114
R20245 VDD.n1907 VDD.n1906 39.2114
R20246 VDD.n1908 VDD.n1897 39.2114
R20247 VDD.n1915 VDD.n1914 39.2114
R20248 VDD.n1916 VDD.n1137 39.2114
R20249 VDD.n1923 VDD.n1922 39.2114
R20250 VDD.n1924 VDD.n1133 39.2114
R20251 VDD.n1932 VDD.n1931 39.2114
R20252 VDD.n2827 VDD.n649 39.2114
R20253 VDD.n2831 VDD.n648 39.2114
R20254 VDD.n2835 VDD.n647 39.2114
R20255 VDD.n2839 VDD.n646 39.2114
R20256 VDD.n2843 VDD.n645 39.2114
R20257 VDD.n2847 VDD.n644 39.2114
R20258 VDD.n2851 VDD.n643 39.2114
R20259 VDD.n2855 VDD.n642 39.2114
R20260 VDD.n2858 VDD.n641 39.2114
R20261 VDD.n3424 VDD.n2920 39.2114
R20262 VDD.n3416 VDD.n2903 39.2114
R20263 VDD.n3412 VDD.n2904 39.2114
R20264 VDD.n3408 VDD.n2905 39.2114
R20265 VDD.n3404 VDD.n2906 39.2114
R20266 VDD.n3400 VDD.n2907 39.2114
R20267 VDD.n3395 VDD.n2908 39.2114
R20268 VDD.n3391 VDD.n2909 39.2114
R20269 VDD.n3889 VDD.n206 39.2114
R20270 VDD.n3896 VDD.n3895 39.2114
R20271 VDD.n204 VDD.n200 39.2114
R20272 VDD.n3903 VDD.n3902 39.2114
R20273 VDD.n199 VDD.n197 39.2114
R20274 VDD.n3912 VDD.n3911 39.2114
R20275 VDD.n196 VDD.n194 39.2114
R20276 VDD.n3919 VDD.n3918 39.2114
R20277 VDD.n193 VDD.n190 39.2114
R20278 VDD.n660 VDD.n650 39.2114
R20279 VDD.n2896 VDD.n651 39.2114
R20280 VDD.n2892 VDD.n652 39.2114
R20281 VDD.n2888 VDD.n653 39.2114
R20282 VDD.n2884 VDD.n654 39.2114
R20283 VDD.n2880 VDD.n655 39.2114
R20284 VDD.n2876 VDD.n656 39.2114
R20285 VDD.n2871 VDD.n657 39.2114
R20286 VDD.n2381 VDD.n2380 39.2114
R20287 VDD.n2378 VDD.n1107 39.2114
R20288 VDD.n2374 VDD.n2373 39.2114
R20289 VDD.n2367 VDD.n1109 39.2114
R20290 VDD.n2366 VDD.n1111 39.2114
R20291 VDD.n2362 VDD.n2361 39.2114
R20292 VDD.n2354 VDD.n1113 39.2114
R20293 VDD.n2353 VDD.n2352 39.2114
R20294 VDD.n2868 VDD.n657 39.2114
R20295 VDD.n2872 VDD.n656 39.2114
R20296 VDD.n2877 VDD.n655 39.2114
R20297 VDD.n2881 VDD.n654 39.2114
R20298 VDD.n2885 VDD.n653 39.2114
R20299 VDD.n2889 VDD.n652 39.2114
R20300 VDD.n2893 VDD.n651 39.2114
R20301 VDD.n2897 VDD.n650 39.2114
R20302 VDD.n2380 VDD.n2379 39.2114
R20303 VDD.n2375 VDD.n1107 39.2114
R20304 VDD.n2373 VDD.n2372 39.2114
R20305 VDD.n2368 VDD.n2367 39.2114
R20306 VDD.n2363 VDD.n1111 39.2114
R20307 VDD.n2361 VDD.n2360 39.2114
R20308 VDD.n2355 VDD.n2354 39.2114
R20309 VDD.n2352 VDD.n2351 39.2114
R20310 VDD.n1581 VDD.n1377 30.8369
R20311 VDD.n1392 VDD.n1391 30.8369
R20312 VDD.n1525 VDD.n1408 30.8369
R20313 VDD.n1495 VDD.n1422 30.8369
R20314 VDD.n1468 VDD.n1439 30.8369
R20315 VDD.n1144 VDD.n1143 30.8369
R20316 VDD.n1809 VDD.n1226 30.8369
R20317 VDD.n1204 VDD.n1203 30.8369
R20318 VDD.n1848 VDD.n1183 30.8369
R20319 VDD.n1871 VDD.n1162 30.8369
R20320 VDD.n4365 VDD.n4364 30.8369
R20321 VDD.n4344 VDD.n4343 30.8369
R20322 VDD.n4423 VDD.n4323 30.8369
R20323 VDD.n4446 VDD.n4302 30.8369
R20324 VDD.n4469 VDD.n4279 30.8369
R20325 VDD.n4059 VDD.n138 30.8369
R20326 VDD.n4007 VDD.n160 30.8369
R20327 VDD.n3946 VDD.n3945 30.8369
R20328 VDD.n4035 VDD.n4034 30.8369
R20329 VDD.n3966 VDD.n3965 30.8369
R20330 VDD.n2825 VDD.n2822 29.5029
R20331 VDD.n3891 VDD.n3888 29.5029
R20332 VDD.n3928 VDD.n183 29.5029
R20333 VDD.n2867 VDD.n2866 29.5029
R20334 VDD.n2860 VDD.n2859 29.5029
R20335 VDD.n1935 VDD.n1934 29.5029
R20336 VDD.n2388 VDD.n1100 29.5029
R20337 VDD.n3390 VDD.n3389 29.5029
R20338 VDD.n3422 VDD.n632 29.5029
R20339 VDD.n3923 VDD.n3922 29.5029
R20340 VDD.n3871 VDD.n3870 29.5029
R20341 VDD.n3153 VDD.n3150 29.5029
R20342 VDD.n3429 VDD.n3428 29.5029
R20343 VDD.n2384 VDD.n2383 29.5029
R20344 VDD.n2900 VDD.n661 29.5029
R20345 VDD.n2349 VDD.n2348 29.5029
R20346 VDD.n1587 VDD.n1372 27.5258
R20347 VDD.n1804 VDD.n1146 27.5258
R20348 VDD.n4074 VDD.n94 27.5258
R20349 VDD.n4264 VDD.n4258 27.5258
R20350 VDD.n7 VDD.t102 25.395
R20351 VDD.n7 VDD.t106 25.395
R20352 VDD.n8 VDD.t116 25.395
R20353 VDD.n8 VDD.t123 25.395
R20354 VDD.n10 VDD.t131 25.395
R20355 VDD.n10 VDD.t133 25.395
R20356 VDD.n12 VDD.t129 25.395
R20357 VDD.n12 VDD.t96 25.395
R20358 VDD.n5 VDD.t98 25.395
R20359 VDD.n5 VDD.t125 25.395
R20360 VDD.n3 VDD.t93 25.395
R20361 VDD.n3 VDD.t127 25.395
R20362 VDD.n1 VDD.t110 25.395
R20363 VDD.n1 VDD.t100 25.395
R20364 VDD.n0 VDD.t113 25.395
R20365 VDD.n0 VDD.t118 25.395
R20366 VDD.n2357 VDD.n1115 24.049
R20367 VDD.n2874 VDD.n663 24.049
R20368 VDD.n1927 VDD.n1135 24.049
R20369 VDD.n674 VDD.n673 24.049
R20370 VDD.n3119 VDD.n3118 24.049
R20371 VDD.n203 VDD.n202 24.049
R20372 VDD.n3397 VDD.n2922 24.049
R20373 VDD.n179 VDD.n178 24.049
R20374 VDD.n1585 VDD.n1365 19.3944
R20375 VDD.n1597 VDD.n1365 19.3944
R20376 VDD.n1597 VDD.n1363 19.3944
R20377 VDD.n1601 VDD.n1363 19.3944
R20378 VDD.n1601 VDD.n1353 19.3944
R20379 VDD.n1613 VDD.n1353 19.3944
R20380 VDD.n1613 VDD.n1351 19.3944
R20381 VDD.n1617 VDD.n1351 19.3944
R20382 VDD.n1617 VDD.n1342 19.3944
R20383 VDD.n1629 VDD.n1342 19.3944
R20384 VDD.n1629 VDD.n1340 19.3944
R20385 VDD.n1633 VDD.n1340 19.3944
R20386 VDD.n1633 VDD.n1330 19.3944
R20387 VDD.n1645 VDD.n1330 19.3944
R20388 VDD.n1645 VDD.n1328 19.3944
R20389 VDD.n1649 VDD.n1328 19.3944
R20390 VDD.n1649 VDD.n1318 19.3944
R20391 VDD.n1661 VDD.n1318 19.3944
R20392 VDD.n1661 VDD.n1316 19.3944
R20393 VDD.n1665 VDD.n1316 19.3944
R20394 VDD.n1665 VDD.n1306 19.3944
R20395 VDD.n1677 VDD.n1306 19.3944
R20396 VDD.n1677 VDD.n1304 19.3944
R20397 VDD.n1681 VDD.n1304 19.3944
R20398 VDD.n1681 VDD.n1290 19.3944
R20399 VDD.n1693 VDD.n1290 19.3944
R20400 VDD.n1693 VDD.n1288 19.3944
R20401 VDD.n1697 VDD.n1288 19.3944
R20402 VDD.n1697 VDD.n1278 19.3944
R20403 VDD.n1709 VDD.n1278 19.3944
R20404 VDD.n1709 VDD.n1276 19.3944
R20405 VDD.n1713 VDD.n1276 19.3944
R20406 VDD.n1713 VDD.n1266 19.3944
R20407 VDD.n1725 VDD.n1266 19.3944
R20408 VDD.n1725 VDD.n1264 19.3944
R20409 VDD.n1729 VDD.n1264 19.3944
R20410 VDD.n1729 VDD.n1254 19.3944
R20411 VDD.n1741 VDD.n1254 19.3944
R20412 VDD.n1741 VDD.n1252 19.3944
R20413 VDD.n1745 VDD.n1252 19.3944
R20414 VDD.n1745 VDD.n1243 19.3944
R20415 VDD.n1757 VDD.n1243 19.3944
R20416 VDD.n1757 VDD.n1240 19.3944
R20417 VDD.n1763 VDD.n1240 19.3944
R20418 VDD.n1763 VDD.n1241 19.3944
R20419 VDD.n1241 VDD.n1230 19.3944
R20420 VDD.n1555 VDD.n1388 19.3944
R20421 VDD.n1559 VDD.n1388 19.3944
R20422 VDD.n1559 VDD.n1386 19.3944
R20423 VDD.n1565 VDD.n1386 19.3944
R20424 VDD.n1565 VDD.n1384 19.3944
R20425 VDD.n1569 VDD.n1384 19.3944
R20426 VDD.n1569 VDD.n1382 19.3944
R20427 VDD.n1576 VDD.n1382 19.3944
R20428 VDD.n1576 VDD.n1378 19.3944
R20429 VDD.n1580 VDD.n1378 19.3944
R20430 VDD.n1529 VDD.n1403 19.3944
R20431 VDD.n1529 VDD.n1401 19.3944
R20432 VDD.n1535 VDD.n1401 19.3944
R20433 VDD.n1535 VDD.n1399 19.3944
R20434 VDD.n1539 VDD.n1399 19.3944
R20435 VDD.n1539 VDD.n1397 19.3944
R20436 VDD.n1545 VDD.n1397 19.3944
R20437 VDD.n1545 VDD.n1395 19.3944
R20438 VDD.n1549 VDD.n1395 19.3944
R20439 VDD.n1549 VDD.n1393 19.3944
R20440 VDD.n1501 VDD.n1418 19.3944
R20441 VDD.n1501 VDD.n1416 19.3944
R20442 VDD.n1505 VDD.n1416 19.3944
R20443 VDD.n1505 VDD.n1414 19.3944
R20444 VDD.n1511 VDD.n1414 19.3944
R20445 VDD.n1511 VDD.n1412 19.3944
R20446 VDD.n1517 VDD.n1412 19.3944
R20447 VDD.n1517 VDD.n1410 19.3944
R20448 VDD.n1410 VDD.n1409 19.3944
R20449 VDD.n1524 VDD.n1409 19.3944
R20450 VDD.n1472 VDD.n1434 19.3944
R20451 VDD.n1472 VDD.n1432 19.3944
R20452 VDD.n1478 VDD.n1432 19.3944
R20453 VDD.n1478 VDD.n1430 19.3944
R20454 VDD.n1483 VDD.n1430 19.3944
R20455 VDD.n1483 VDD.n1428 19.3944
R20456 VDD.n1428 VDD.n1425 19.3944
R20457 VDD.n1490 VDD.n1425 19.3944
R20458 VDD.n1490 VDD.n1423 19.3944
R20459 VDD.n1494 VDD.n1423 19.3944
R20460 VDD.n1448 VDD.n1446 19.3944
R20461 VDD.n1448 VDD.n1445 19.3944
R20462 VDD.n1454 VDD.n1445 19.3944
R20463 VDD.n1454 VDD.n1443 19.3944
R20464 VDD.n1460 VDD.n1443 19.3944
R20465 VDD.n1460 VDD.n1441 19.3944
R20466 VDD.n1441 VDD.n1440 19.3944
R20467 VDD.n1467 VDD.n1440 19.3944
R20468 VDD.n1799 VDD.n1798 19.3944
R20469 VDD.n1798 VDD.n1797 19.3944
R20470 VDD.n1797 VDD.n1774 19.3944
R20471 VDD.n1775 VDD.n1774 19.3944
R20472 VDD.n1790 VDD.n1775 19.3944
R20473 VDD.n1790 VDD.n1789 19.3944
R20474 VDD.n1789 VDD.n1788 19.3944
R20475 VDD.n1788 VDD.n1783 19.3944
R20476 VDD.n1589 VDD.n1369 19.3944
R20477 VDD.n1593 VDD.n1369 19.3944
R20478 VDD.n1593 VDD.n1359 19.3944
R20479 VDD.n1605 VDD.n1359 19.3944
R20480 VDD.n1605 VDD.n1357 19.3944
R20481 VDD.n1609 VDD.n1357 19.3944
R20482 VDD.n1609 VDD.n1348 19.3944
R20483 VDD.n1621 VDD.n1348 19.3944
R20484 VDD.n1621 VDD.n1346 19.3944
R20485 VDD.n1625 VDD.n1346 19.3944
R20486 VDD.n1625 VDD.n1336 19.3944
R20487 VDD.n1637 VDD.n1336 19.3944
R20488 VDD.n1637 VDD.n1334 19.3944
R20489 VDD.n1641 VDD.n1334 19.3944
R20490 VDD.n1641 VDD.n1324 19.3944
R20491 VDD.n1653 VDD.n1324 19.3944
R20492 VDD.n1653 VDD.n1322 19.3944
R20493 VDD.n1657 VDD.n1322 19.3944
R20494 VDD.n1657 VDD.n1312 19.3944
R20495 VDD.n1669 VDD.n1312 19.3944
R20496 VDD.n1669 VDD.n1310 19.3944
R20497 VDD.n1673 VDD.n1310 19.3944
R20498 VDD.n1673 VDD.n1301 19.3944
R20499 VDD.n1685 VDD.n1301 19.3944
R20500 VDD.n1685 VDD.n1294 19.3944
R20501 VDD.n1689 VDD.n1294 19.3944
R20502 VDD.n1689 VDD.n1284 19.3944
R20503 VDD.n1701 VDD.n1284 19.3944
R20504 VDD.n1701 VDD.n1282 19.3944
R20505 VDD.n1705 VDD.n1282 19.3944
R20506 VDD.n1705 VDD.n1272 19.3944
R20507 VDD.n1717 VDD.n1272 19.3944
R20508 VDD.n1717 VDD.n1270 19.3944
R20509 VDD.n1721 VDD.n1270 19.3944
R20510 VDD.n1721 VDD.n1260 19.3944
R20511 VDD.n1733 VDD.n1260 19.3944
R20512 VDD.n1733 VDD.n1258 19.3944
R20513 VDD.n1737 VDD.n1258 19.3944
R20514 VDD.n1737 VDD.n1249 19.3944
R20515 VDD.n1749 VDD.n1249 19.3944
R20516 VDD.n1749 VDD.n1247 19.3944
R20517 VDD.n1753 VDD.n1247 19.3944
R20518 VDD.n1753 VDD.n1236 19.3944
R20519 VDD.n1767 VDD.n1236 19.3944
R20520 VDD.n1767 VDD.n1234 19.3944
R20521 VDD.n1802 VDD.n1234 19.3944
R20522 VDD.n1206 VDD.n1205 19.3944
R20523 VDD.n1821 VDD.n1206 19.3944
R20524 VDD.n1821 VDD.n1820 19.3944
R20525 VDD.n1820 VDD.n1819 19.3944
R20526 VDD.n1819 VDD.n1214 19.3944
R20527 VDD.n1815 VDD.n1214 19.3944
R20528 VDD.n1815 VDD.n1814 19.3944
R20529 VDD.n1814 VDD.n1813 19.3944
R20530 VDD.n1813 VDD.n1222 19.3944
R20531 VDD.n1844 VDD.n1181 19.3944
R20532 VDD.n1844 VDD.n1186 19.3944
R20533 VDD.n1839 VDD.n1186 19.3944
R20534 VDD.n1839 VDD.n1838 19.3944
R20535 VDD.n1838 VDD.n1837 19.3944
R20536 VDD.n1837 VDD.n1192 19.3944
R20537 VDD.n1832 VDD.n1192 19.3944
R20538 VDD.n1832 VDD.n1831 19.3944
R20539 VDD.n1831 VDD.n1830 19.3944
R20540 VDD.n1830 VDD.n1199 19.3944
R20541 VDD.n1867 VDD.n1160 19.3944
R20542 VDD.n1867 VDD.n1165 19.3944
R20543 VDD.n1862 VDD.n1165 19.3944
R20544 VDD.n1862 VDD.n1861 19.3944
R20545 VDD.n1861 VDD.n1860 19.3944
R20546 VDD.n1860 VDD.n1171 19.3944
R20547 VDD.n1855 VDD.n1171 19.3944
R20548 VDD.n1855 VDD.n1854 19.3944
R20549 VDD.n1854 VDD.n1853 19.3944
R20550 VDD.n1853 VDD.n1178 19.3944
R20551 VDD.n1147 VDD.n1141 19.3944
R20552 VDD.n1885 VDD.n1884 19.3944
R20553 VDD.n1884 VDD.n1883 19.3944
R20554 VDD.n1883 VDD.n1150 19.3944
R20555 VDD.n1878 VDD.n1150 19.3944
R20556 VDD.n1878 VDD.n1877 19.3944
R20557 VDD.n1877 VDD.n1876 19.3944
R20558 VDD.n1876 VDD.n1157 19.3944
R20559 VDD.n4085 VDD.n92 19.3944
R20560 VDD.n4085 VDD.n90 19.3944
R20561 VDD.n4089 VDD.n90 19.3944
R20562 VDD.n4089 VDD.n80 19.3944
R20563 VDD.n4101 VDD.n80 19.3944
R20564 VDD.n4101 VDD.n78 19.3944
R20565 VDD.n4105 VDD.n78 19.3944
R20566 VDD.n4105 VDD.n68 19.3944
R20567 VDD.n4116 VDD.n68 19.3944
R20568 VDD.n4116 VDD.n66 19.3944
R20569 VDD.n4120 VDD.n66 19.3944
R20570 VDD.n4120 VDD.n56 19.3944
R20571 VDD.n4132 VDD.n56 19.3944
R20572 VDD.n4132 VDD.n54 19.3944
R20573 VDD.n4136 VDD.n54 19.3944
R20574 VDD.n4136 VDD.n44 19.3944
R20575 VDD.n4148 VDD.n44 19.3944
R20576 VDD.n4148 VDD.n42 19.3944
R20577 VDD.n4152 VDD.n42 19.3944
R20578 VDD.n4152 VDD.n32 19.3944
R20579 VDD.n4164 VDD.n32 19.3944
R20580 VDD.n4164 VDD.n30 19.3944
R20581 VDD.n4538 VDD.n30 19.3944
R20582 VDD.n4538 VDD.n4537 19.3944
R20583 VDD.n4537 VDD.n4536 19.3944
R20584 VDD.n4536 VDD.n4170 19.3944
R20585 VDD.n4225 VDD.n4170 19.3944
R20586 VDD.n4226 VDD.n4225 19.3944
R20587 VDD.n4227 VDD.n4226 19.3944
R20588 VDD.n4227 VDD.n4221 19.3944
R20589 VDD.n4231 VDD.n4221 19.3944
R20590 VDD.n4232 VDD.n4231 19.3944
R20591 VDD.n4233 VDD.n4232 19.3944
R20592 VDD.n4233 VDD.n4218 19.3944
R20593 VDD.n4237 VDD.n4218 19.3944
R20594 VDD.n4238 VDD.n4237 19.3944
R20595 VDD.n4239 VDD.n4238 19.3944
R20596 VDD.n4239 VDD.n4215 19.3944
R20597 VDD.n4503 VDD.n4215 19.3944
R20598 VDD.n4503 VDD.n4502 19.3944
R20599 VDD.n4502 VDD.n4501 19.3944
R20600 VDD.n4501 VDD.n4245 19.3944
R20601 VDD.n4370 VDD.n4245 19.3944
R20602 VDD.n4374 VDD.n4370 19.3944
R20603 VDD.n4375 VDD.n4374 19.3944
R20604 VDD.n4376 VDD.n4375 19.3944
R20605 VDD.n4400 VDD.n4399 19.3944
R20606 VDD.n4399 VDD.n4398 19.3944
R20607 VDD.n4398 VDD.n4349 19.3944
R20608 VDD.n4393 VDD.n4349 19.3944
R20609 VDD.n4393 VDD.n4392 19.3944
R20610 VDD.n4392 VDD.n4391 19.3944
R20611 VDD.n4391 VDD.n4356 19.3944
R20612 VDD.n4386 VDD.n4356 19.3944
R20613 VDD.n4386 VDD.n4385 19.3944
R20614 VDD.n4385 VDD.n4384 19.3944
R20615 VDD.n4419 VDD.n4321 19.3944
R20616 VDD.n4419 VDD.n4326 19.3944
R20617 VDD.n4414 VDD.n4326 19.3944
R20618 VDD.n4414 VDD.n4413 19.3944
R20619 VDD.n4413 VDD.n4412 19.3944
R20620 VDD.n4412 VDD.n4332 19.3944
R20621 VDD.n4407 VDD.n4332 19.3944
R20622 VDD.n4407 VDD.n4406 19.3944
R20623 VDD.n4406 VDD.n4405 19.3944
R20624 VDD.n4405 VDD.n4339 19.3944
R20625 VDD.n4442 VDD.n4300 19.3944
R20626 VDD.n4442 VDD.n4305 19.3944
R20627 VDD.n4437 VDD.n4305 19.3944
R20628 VDD.n4437 VDD.n4436 19.3944
R20629 VDD.n4436 VDD.n4435 19.3944
R20630 VDD.n4435 VDD.n4311 19.3944
R20631 VDD.n4430 VDD.n4311 19.3944
R20632 VDD.n4430 VDD.n4429 19.3944
R20633 VDD.n4429 VDD.n4428 19.3944
R20634 VDD.n4428 VDD.n4318 19.3944
R20635 VDD.n4465 VDD.n4277 19.3944
R20636 VDD.n4465 VDD.n4283 19.3944
R20637 VDD.n4460 VDD.n4283 19.3944
R20638 VDD.n4460 VDD.n4459 19.3944
R20639 VDD.n4459 VDD.n4458 19.3944
R20640 VDD.n4458 VDD.n4290 19.3944
R20641 VDD.n4453 VDD.n4290 19.3944
R20642 VDD.n4453 VDD.n4452 19.3944
R20643 VDD.n4452 VDD.n4451 19.3944
R20644 VDD.n4451 VDD.n4297 19.3944
R20645 VDD.n4485 VDD.n4263 19.3944
R20646 VDD.n4265 VDD.n4263 19.3944
R20647 VDD.n4478 VDD.n4265 19.3944
R20648 VDD.n4478 VDD.n4477 19.3944
R20649 VDD.n4477 VDD.n4476 19.3944
R20650 VDD.n4476 VDD.n4271 19.3944
R20651 VDD.n4471 VDD.n4271 19.3944
R20652 VDD.n4471 VDD.n4470 19.3944
R20653 VDD.n4081 VDD.n96 19.3944
R20654 VDD.n4081 VDD.n86 19.3944
R20655 VDD.n4093 VDD.n86 19.3944
R20656 VDD.n4093 VDD.n84 19.3944
R20657 VDD.n4097 VDD.n84 19.3944
R20658 VDD.n4097 VDD.n74 19.3944
R20659 VDD.n4108 VDD.n74 19.3944
R20660 VDD.n4108 VDD.n72 19.3944
R20661 VDD.n4112 VDD.n72 19.3944
R20662 VDD.n4112 VDD.n62 19.3944
R20663 VDD.n4124 VDD.n62 19.3944
R20664 VDD.n4124 VDD.n60 19.3944
R20665 VDD.n4128 VDD.n60 19.3944
R20666 VDD.n4128 VDD.n50 19.3944
R20667 VDD.n4140 VDD.n50 19.3944
R20668 VDD.n4140 VDD.n48 19.3944
R20669 VDD.n4144 VDD.n48 19.3944
R20670 VDD.n4144 VDD.n38 19.3944
R20671 VDD.n4156 VDD.n38 19.3944
R20672 VDD.n4156 VDD.n36 19.3944
R20673 VDD.n4160 VDD.n36 19.3944
R20674 VDD.n4160 VDD.n22 19.3944
R20675 VDD.n4541 VDD.n22 19.3944
R20676 VDD.n4541 VDD.n23 19.3944
R20677 VDD.n4532 VDD.n23 19.3944
R20678 VDD.n4532 VDD.n4531 19.3944
R20679 VDD.n4531 VDD.n4530 19.3944
R20680 VDD.n4530 VDD.n4177 19.3944
R20681 VDD.n4524 VDD.n4177 19.3944
R20682 VDD.n4524 VDD.n4523 19.3944
R20683 VDD.n4523 VDD.n4522 19.3944
R20684 VDD.n4522 VDD.n4188 19.3944
R20685 VDD.n4516 VDD.n4188 19.3944
R20686 VDD.n4516 VDD.n4515 19.3944
R20687 VDD.n4515 VDD.n4514 19.3944
R20688 VDD.n4514 VDD.n4199 19.3944
R20689 VDD.n4508 VDD.n4199 19.3944
R20690 VDD.n4508 VDD.n4507 19.3944
R20691 VDD.n4507 VDD.n4506 19.3944
R20692 VDD.n4506 VDD.n4210 19.3944
R20693 VDD.n4497 VDD.n4210 19.3944
R20694 VDD.n4497 VDD.n4496 19.3944
R20695 VDD.n4496 VDD.n4495 19.3944
R20696 VDD.n4495 VDD.n4253 19.3944
R20697 VDD.n4489 VDD.n4253 19.3944
R20698 VDD.n4489 VDD.n4488 19.3944
R20699 VDD.n4077 VDD.n98 19.3944
R20700 VDD.n4072 VDD.n98 19.3944
R20701 VDD.n4072 VDD.n4071 19.3944
R20702 VDD.n4071 VDD.n4070 19.3944
R20703 VDD.n4070 VDD.n4067 19.3944
R20704 VDD.n4067 VDD.n4066 19.3944
R20705 VDD.n4066 VDD.n4063 19.3944
R20706 VDD.n4063 VDD.n4062 19.3944
R20707 VDD.n4029 VDD.n148 19.3944
R20708 VDD.n4029 VDD.n4026 19.3944
R20709 VDD.n4026 VDD.n4023 19.3944
R20710 VDD.n4023 VDD.n4022 19.3944
R20711 VDD.n4022 VDD.n4019 19.3944
R20712 VDD.n4019 VDD.n4018 19.3944
R20713 VDD.n4018 VDD.n4015 19.3944
R20714 VDD.n4015 VDD.n4014 19.3944
R20715 VDD.n4014 VDD.n4011 19.3944
R20716 VDD.n4011 VDD.n4010 19.3944
R20717 VDD.n4006 VDD.n4003 19.3944
R20718 VDD.n4003 VDD.n4002 19.3944
R20719 VDD.n4002 VDD.n3999 19.3944
R20720 VDD.n3999 VDD.n3998 19.3944
R20721 VDD.n3998 VDD.n3995 19.3944
R20722 VDD.n3995 VDD.n3994 19.3944
R20723 VDD.n3994 VDD.n3991 19.3944
R20724 VDD.n3991 VDD.n3990 19.3944
R20725 VDD.n3990 VDD.n3987 19.3944
R20726 VDD.n3987 VDD.n170 19.3944
R20727 VDD.n4055 VDD.n4054 19.3944
R20728 VDD.n4051 VDD.n4050 19.3944
R20729 VDD.n4050 VDD.n4047 19.3944
R20730 VDD.n4047 VDD.n4046 19.3944
R20731 VDD.n4046 VDD.n4043 19.3944
R20732 VDD.n4043 VDD.n4042 19.3944
R20733 VDD.n4042 VDD.n4039 19.3944
R20734 VDD.n4039 VDD.n4038 19.3944
R20735 VDD.n3950 VDD.n3949 19.3944
R20736 VDD.n3983 VDD.n3982 19.3944
R20737 VDD.n3982 VDD.n3979 19.3944
R20738 VDD.n3979 VDD.n3978 19.3944
R20739 VDD.n3978 VDD.n3975 19.3944
R20740 VDD.n3975 VDD.n3974 19.3944
R20741 VDD.n3974 VDD.n3971 19.3944
R20742 VDD.n3971 VDD.n3970 19.3944
R20743 VDD.n3970 VDD.n3967 19.3944
R20744 VDD.n1525 VDD.n1403 18.8126
R20745 VDD.n1848 VDD.n1181 18.8126
R20746 VDD.n4423 VDD.n4321 18.8126
R20747 VDD.n4007 VDD.n4006 18.8126
R20748 VDD.n2386 VDD.n1102 18.2003
R20749 VDD.n2902 VDD.n640 18.2003
R20750 VDD.n3425 VDD.n634 18.2003
R20751 VDD.n3925 VDD.n175 18.2003
R20752 VDD.n1468 VDD.n1467 18.0369
R20753 VDD.n1783 VDD.n1144 18.0369
R20754 VDD.n4470 VDD.n4469 18.0369
R20755 VDD.n4062 VDD.n4059 18.0369
R20756 VDD.n1581 VDD.n1580 15.7096
R20757 VDD.n1809 VDD.n1222 15.7096
R20758 VDD.n4384 VDD.n4365 15.7096
R20759 VDD.n3967 VDD.n3966 15.7096
R20760 VDD.n1587 VDD.n1367 15.0417
R20761 VDD.n1595 VDD.n1367 15.0417
R20762 VDD.n1595 VDD.n1361 15.0417
R20763 VDD.n1603 VDD.n1361 15.0417
R20764 VDD.n1603 VDD.n1355 15.0417
R20765 VDD.n1611 VDD.n1355 15.0417
R20766 VDD.n1611 VDD.t1 15.0417
R20767 VDD.n1619 VDD.t1 15.0417
R20768 VDD.n1619 VDD.n1344 15.0417
R20769 VDD.n1627 VDD.n1344 15.0417
R20770 VDD.n1627 VDD.n1338 15.0417
R20771 VDD.n1635 VDD.n1338 15.0417
R20772 VDD.n1635 VDD.n1332 15.0417
R20773 VDD.n1643 VDD.n1332 15.0417
R20774 VDD.n1643 VDD.n1326 15.0417
R20775 VDD.n1651 VDD.n1326 15.0417
R20776 VDD.n1651 VDD.n1320 15.0417
R20777 VDD.n1659 VDD.n1320 15.0417
R20778 VDD.n1659 VDD.n1314 15.0417
R20779 VDD.n1667 VDD.n1314 15.0417
R20780 VDD.n1667 VDD.n1308 15.0417
R20781 VDD.n1675 VDD.n1308 15.0417
R20782 VDD.n1675 VDD.t135 15.0417
R20783 VDD.n1683 VDD.t135 15.0417
R20784 VDD.n1683 VDD.n1292 15.0417
R20785 VDD.n1691 VDD.n1292 15.0417
R20786 VDD.n1691 VDD.n1286 15.0417
R20787 VDD.n1699 VDD.n1286 15.0417
R20788 VDD.n1699 VDD.n1280 15.0417
R20789 VDD.n1707 VDD.n1280 15.0417
R20790 VDD.n1707 VDD.n1274 15.0417
R20791 VDD.n1715 VDD.n1274 15.0417
R20792 VDD.n1715 VDD.n1268 15.0417
R20793 VDD.n1723 VDD.n1268 15.0417
R20794 VDD.n1723 VDD.n1262 15.0417
R20795 VDD.n1731 VDD.n1262 15.0417
R20796 VDD.n1731 VDD.n1256 15.0417
R20797 VDD.n1739 VDD.n1256 15.0417
R20798 VDD.n1739 VDD.t33 15.0417
R20799 VDD.n1747 VDD.t33 15.0417
R20800 VDD.n1747 VDD.n1245 15.0417
R20801 VDD.n1755 VDD.n1245 15.0417
R20802 VDD.n1755 VDD.n1238 15.0417
R20803 VDD.n1765 VDD.n1238 15.0417
R20804 VDD.n1765 VDD.n1231 15.0417
R20805 VDD.n1804 VDD.n1231 15.0417
R20806 VDD.n4083 VDD.n94 15.0417
R20807 VDD.n4083 VDD.n88 15.0417
R20808 VDD.n4091 VDD.n88 15.0417
R20809 VDD.n4091 VDD.n82 15.0417
R20810 VDD.n4099 VDD.n82 15.0417
R20811 VDD.n4099 VDD.n76 15.0417
R20812 VDD.t11 VDD.n76 15.0417
R20813 VDD.t11 VDD.n70 15.0417
R20814 VDD.n4114 VDD.n70 15.0417
R20815 VDD.n4114 VDD.n64 15.0417
R20816 VDD.n4122 VDD.n64 15.0417
R20817 VDD.n4122 VDD.n58 15.0417
R20818 VDD.n4130 VDD.n58 15.0417
R20819 VDD.n4130 VDD.n52 15.0417
R20820 VDD.n4138 VDD.n52 15.0417
R20821 VDD.n4138 VDD.n46 15.0417
R20822 VDD.n4146 VDD.n46 15.0417
R20823 VDD.n4146 VDD.n40 15.0417
R20824 VDD.n4154 VDD.n40 15.0417
R20825 VDD.n4154 VDD.n34 15.0417
R20826 VDD.n4162 VDD.n34 15.0417
R20827 VDD.n4162 VDD.n26 15.0417
R20828 VDD.t137 VDD.n26 15.0417
R20829 VDD.t137 VDD.n27 15.0417
R20830 VDD.n4534 VDD.n27 15.0417
R20831 VDD.n4534 VDD.n4172 15.0417
R20832 VDD.n4528 VDD.n4172 15.0417
R20833 VDD.n4528 VDD.n4527 15.0417
R20834 VDD.n4527 VDD.n4526 15.0417
R20835 VDD.n4526 VDD.n4182 15.0417
R20836 VDD.n4520 VDD.n4182 15.0417
R20837 VDD.n4520 VDD.n4519 15.0417
R20838 VDD.n4519 VDD.n4518 15.0417
R20839 VDD.n4518 VDD.n4193 15.0417
R20840 VDD.n4512 VDD.n4193 15.0417
R20841 VDD.n4512 VDD.n4511 15.0417
R20842 VDD.n4511 VDD.n4510 15.0417
R20843 VDD.n4510 VDD.n4204 15.0417
R20844 VDD.t43 VDD.n4204 15.0417
R20845 VDD.t43 VDD.n4212 15.0417
R20846 VDD.n4499 VDD.n4212 15.0417
R20847 VDD.n4499 VDD.n4247 15.0417
R20848 VDD.n4493 VDD.n4247 15.0417
R20849 VDD.n4493 VDD.n4492 15.0417
R20850 VDD.n4492 VDD.n4491 15.0417
R20851 VDD.n4491 VDD.n4258 15.0417
R20852 VDD.n1495 VDD.n1418 13.3823
R20853 VDD.n1871 VDD.n1160 13.3823
R20854 VDD.n4446 VDD.n4300 13.3823
R20855 VDD.n4035 VDD.n148 13.3823
R20856 VDD.n1495 VDD.n1494 12.6066
R20857 VDD.n1871 VDD.n1157 12.6066
R20858 VDD.n4446 VDD.n4297 12.6066
R20859 VDD.n4038 VDD.n4035 12.6066
R20860 VDD.n2859 VDD.n2857 10.6151
R20861 VDD.n2857 VDD.n2854 10.6151
R20862 VDD.n2854 VDD.n2853 10.6151
R20863 VDD.n2853 VDD.n2850 10.6151
R20864 VDD.n2850 VDD.n2849 10.6151
R20865 VDD.n2849 VDD.n2846 10.6151
R20866 VDD.n2846 VDD.n2845 10.6151
R20867 VDD.n2845 VDD.n2842 10.6151
R20868 VDD.n2842 VDD.n2841 10.6151
R20869 VDD.n2841 VDD.n2838 10.6151
R20870 VDD.n2838 VDD.n2837 10.6151
R20871 VDD.n2837 VDD.n2834 10.6151
R20872 VDD.n2834 VDD.n2833 10.6151
R20873 VDD.n2830 VDD.n2829 10.6151
R20874 VDD.n2829 VDD.n2826 10.6151
R20875 VDD.n2826 VDD.n2825 10.6151
R20876 VDD.n1937 VDD.n1935 10.6151
R20877 VDD.n1938 VDD.n1937 10.6151
R20878 VDD.n1940 VDD.n1938 10.6151
R20879 VDD.n1941 VDD.n1940 10.6151
R20880 VDD.n1943 VDD.n1941 10.6151
R20881 VDD.n1944 VDD.n1943 10.6151
R20882 VDD.n1946 VDD.n1944 10.6151
R20883 VDD.n1947 VDD.n1946 10.6151
R20884 VDD.n1949 VDD.n1947 10.6151
R20885 VDD.n1950 VDD.n1949 10.6151
R20886 VDD.n1952 VDD.n1950 10.6151
R20887 VDD.n1953 VDD.n1952 10.6151
R20888 VDD.n1955 VDD.n1953 10.6151
R20889 VDD.n1956 VDD.n1955 10.6151
R20890 VDD.n1958 VDD.n1956 10.6151
R20891 VDD.n1959 VDD.n1958 10.6151
R20892 VDD.n1961 VDD.n1959 10.6151
R20893 VDD.n1962 VDD.n1961 10.6151
R20894 VDD.n1964 VDD.n1962 10.6151
R20895 VDD.n1965 VDD.n1964 10.6151
R20896 VDD.n1967 VDD.n1965 10.6151
R20897 VDD.n1968 VDD.n1967 10.6151
R20898 VDD.n1970 VDD.n1968 10.6151
R20899 VDD.n1971 VDD.n1970 10.6151
R20900 VDD.n1973 VDD.n1971 10.6151
R20901 VDD.n1974 VDD.n1973 10.6151
R20902 VDD.n1976 VDD.n1974 10.6151
R20903 VDD.n1977 VDD.n1976 10.6151
R20904 VDD.n1979 VDD.n1977 10.6151
R20905 VDD.n1980 VDD.n1979 10.6151
R20906 VDD.n1982 VDD.n1980 10.6151
R20907 VDD.n1983 VDD.n1982 10.6151
R20908 VDD.n1985 VDD.n1983 10.6151
R20909 VDD.n1986 VDD.n1985 10.6151
R20910 VDD.n1988 VDD.n1986 10.6151
R20911 VDD.n1989 VDD.n1988 10.6151
R20912 VDD.n1991 VDD.n1989 10.6151
R20913 VDD.n1992 VDD.n1991 10.6151
R20914 VDD.n1994 VDD.n1992 10.6151
R20915 VDD.n1995 VDD.n1994 10.6151
R20916 VDD.n1997 VDD.n1995 10.6151
R20917 VDD.n1998 VDD.n1997 10.6151
R20918 VDD.n2000 VDD.n1998 10.6151
R20919 VDD.n2001 VDD.n2000 10.6151
R20920 VDD.n2003 VDD.n2001 10.6151
R20921 VDD.n2004 VDD.n2003 10.6151
R20922 VDD.n2006 VDD.n2004 10.6151
R20923 VDD.n2007 VDD.n2006 10.6151
R20924 VDD.n2009 VDD.n2007 10.6151
R20925 VDD.n2010 VDD.n2009 10.6151
R20926 VDD.n2012 VDD.n2010 10.6151
R20927 VDD.n2013 VDD.n2012 10.6151
R20928 VDD.n2015 VDD.n2013 10.6151
R20929 VDD.n2016 VDD.n2015 10.6151
R20930 VDD.n2018 VDD.n2016 10.6151
R20931 VDD.n2019 VDD.n2018 10.6151
R20932 VDD.n2021 VDD.n2019 10.6151
R20933 VDD.n2022 VDD.n2021 10.6151
R20934 VDD.n2024 VDD.n2022 10.6151
R20935 VDD.n2025 VDD.n2024 10.6151
R20936 VDD.n2027 VDD.n2025 10.6151
R20937 VDD.n2028 VDD.n2027 10.6151
R20938 VDD.n2030 VDD.n2028 10.6151
R20939 VDD.n2031 VDD.n2030 10.6151
R20940 VDD.n2033 VDD.n2031 10.6151
R20941 VDD.n2034 VDD.n2033 10.6151
R20942 VDD.n2036 VDD.n2034 10.6151
R20943 VDD.n2037 VDD.n2036 10.6151
R20944 VDD.n2039 VDD.n2037 10.6151
R20945 VDD.n2040 VDD.n2039 10.6151
R20946 VDD.n2042 VDD.n2040 10.6151
R20947 VDD.n2043 VDD.n2042 10.6151
R20948 VDD.n2045 VDD.n2043 10.6151
R20949 VDD.n2046 VDD.n2045 10.6151
R20950 VDD.n2048 VDD.n2046 10.6151
R20951 VDD.n2049 VDD.n2048 10.6151
R20952 VDD.n2051 VDD.n2049 10.6151
R20953 VDD.n2052 VDD.n2051 10.6151
R20954 VDD.n2054 VDD.n2052 10.6151
R20955 VDD.n2055 VDD.n2054 10.6151
R20956 VDD.n2057 VDD.n2055 10.6151
R20957 VDD.n2058 VDD.n2057 10.6151
R20958 VDD.n2060 VDD.n2058 10.6151
R20959 VDD.n2061 VDD.n2060 10.6151
R20960 VDD.n2063 VDD.n2061 10.6151
R20961 VDD.n2064 VDD.n2063 10.6151
R20962 VDD.n2066 VDD.n2064 10.6151
R20963 VDD.n2067 VDD.n2066 10.6151
R20964 VDD.n2069 VDD.n2067 10.6151
R20965 VDD.n2070 VDD.n2069 10.6151
R20966 VDD.n2072 VDD.n2070 10.6151
R20967 VDD.n2073 VDD.n2072 10.6151
R20968 VDD.n2075 VDD.n2073 10.6151
R20969 VDD.n2076 VDD.n2075 10.6151
R20970 VDD.n2078 VDD.n2076 10.6151
R20971 VDD.n2079 VDD.n2078 10.6151
R20972 VDD.n2081 VDD.n2079 10.6151
R20973 VDD.n2082 VDD.n2081 10.6151
R20974 VDD.n2084 VDD.n2082 10.6151
R20975 VDD.n2085 VDD.n2084 10.6151
R20976 VDD.n2087 VDD.n2085 10.6151
R20977 VDD.n2088 VDD.n2087 10.6151
R20978 VDD.n2090 VDD.n2088 10.6151
R20979 VDD.n2091 VDD.n2090 10.6151
R20980 VDD.n2093 VDD.n2091 10.6151
R20981 VDD.n2094 VDD.n2093 10.6151
R20982 VDD.n2096 VDD.n2094 10.6151
R20983 VDD.n2097 VDD.n2096 10.6151
R20984 VDD.n2099 VDD.n2097 10.6151
R20985 VDD.n2100 VDD.n2099 10.6151
R20986 VDD.n2102 VDD.n2100 10.6151
R20987 VDD.n2103 VDD.n2102 10.6151
R20988 VDD.n2105 VDD.n2103 10.6151
R20989 VDD.n2106 VDD.n2105 10.6151
R20990 VDD.n2108 VDD.n2106 10.6151
R20991 VDD.n2109 VDD.n2108 10.6151
R20992 VDD.n2111 VDD.n2109 10.6151
R20993 VDD.n2112 VDD.n2111 10.6151
R20994 VDD.n2114 VDD.n2112 10.6151
R20995 VDD.n2115 VDD.n2114 10.6151
R20996 VDD.n2117 VDD.n2115 10.6151
R20997 VDD.n2118 VDD.n2117 10.6151
R20998 VDD.n2120 VDD.n2118 10.6151
R20999 VDD.n2121 VDD.n2120 10.6151
R21000 VDD.n2123 VDD.n2121 10.6151
R21001 VDD.n2124 VDD.n2123 10.6151
R21002 VDD.n2126 VDD.n2124 10.6151
R21003 VDD.n2127 VDD.n2126 10.6151
R21004 VDD.n2129 VDD.n2127 10.6151
R21005 VDD.n2130 VDD.n2129 10.6151
R21006 VDD.n2132 VDD.n2130 10.6151
R21007 VDD.n2133 VDD.n2132 10.6151
R21008 VDD.n2145 VDD.n2133 10.6151
R21009 VDD.n2145 VDD.n2144 10.6151
R21010 VDD.n2144 VDD.n2143 10.6151
R21011 VDD.n2143 VDD.n2141 10.6151
R21012 VDD.n2141 VDD.n2140 10.6151
R21013 VDD.n2140 VDD.n2138 10.6151
R21014 VDD.n2138 VDD.n2137 10.6151
R21015 VDD.n2137 VDD.n2135 10.6151
R21016 VDD.n2135 VDD.n2134 10.6151
R21017 VDD.n2134 VDD.n675 10.6151
R21018 VDD.n2820 VDD.n675 10.6151
R21019 VDD.n2821 VDD.n2820 10.6151
R21020 VDD.n2822 VDD.n2821 10.6151
R21021 VDD.n1902 VDD.n1100 10.6151
R21022 VDD.n1903 VDD.n1902 10.6151
R21023 VDD.n1904 VDD.n1903 10.6151
R21024 VDD.n1904 VDD.n1898 10.6151
R21025 VDD.n1910 VDD.n1898 10.6151
R21026 VDD.n1911 VDD.n1910 10.6151
R21027 VDD.n1912 VDD.n1911 10.6151
R21028 VDD.n1912 VDD.n1896 10.6151
R21029 VDD.n1919 VDD.n1918 10.6151
R21030 VDD.n1920 VDD.n1919 10.6151
R21031 VDD.n1920 VDD.n1136 10.6151
R21032 VDD.n1926 VDD.n1136 10.6151
R21033 VDD.n1929 VDD.n1928 10.6151
R21034 VDD.n1929 VDD.n1132 10.6151
R21035 VDD.n1934 VDD.n1132 10.6151
R21036 VDD.n2389 VDD.n2388 10.6151
R21037 VDD.n2390 VDD.n2389 10.6151
R21038 VDD.n2390 VDD.n1088 10.6151
R21039 VDD.n2400 VDD.n1088 10.6151
R21040 VDD.n2401 VDD.n2400 10.6151
R21041 VDD.n2402 VDD.n2401 10.6151
R21042 VDD.n2402 VDD.n1076 10.6151
R21043 VDD.n2412 VDD.n1076 10.6151
R21044 VDD.n2413 VDD.n2412 10.6151
R21045 VDD.n2414 VDD.n2413 10.6151
R21046 VDD.n2414 VDD.n1064 10.6151
R21047 VDD.n2424 VDD.n1064 10.6151
R21048 VDD.n2425 VDD.n2424 10.6151
R21049 VDD.n2426 VDD.n2425 10.6151
R21050 VDD.n2426 VDD.n1052 10.6151
R21051 VDD.n2436 VDD.n1052 10.6151
R21052 VDD.n2437 VDD.n2436 10.6151
R21053 VDD.n2438 VDD.n2437 10.6151
R21054 VDD.n2438 VDD.n1040 10.6151
R21055 VDD.n2448 VDD.n1040 10.6151
R21056 VDD.n2449 VDD.n2448 10.6151
R21057 VDD.n2450 VDD.n2449 10.6151
R21058 VDD.n2450 VDD.n1028 10.6151
R21059 VDD.n2460 VDD.n1028 10.6151
R21060 VDD.n2461 VDD.n2460 10.6151
R21061 VDD.n2462 VDD.n2461 10.6151
R21062 VDD.n2462 VDD.n1016 10.6151
R21063 VDD.n2472 VDD.n1016 10.6151
R21064 VDD.n2473 VDD.n2472 10.6151
R21065 VDD.n2474 VDD.n2473 10.6151
R21066 VDD.n2474 VDD.n1004 10.6151
R21067 VDD.n2484 VDD.n1004 10.6151
R21068 VDD.n2485 VDD.n2484 10.6151
R21069 VDD.n2486 VDD.n2485 10.6151
R21070 VDD.n2486 VDD.n992 10.6151
R21071 VDD.n2496 VDD.n992 10.6151
R21072 VDD.n2497 VDD.n2496 10.6151
R21073 VDD.n2498 VDD.n2497 10.6151
R21074 VDD.n2498 VDD.n980 10.6151
R21075 VDD.n2508 VDD.n980 10.6151
R21076 VDD.n2509 VDD.n2508 10.6151
R21077 VDD.n2510 VDD.n2509 10.6151
R21078 VDD.n2510 VDD.n968 10.6151
R21079 VDD.n2520 VDD.n968 10.6151
R21080 VDD.n2521 VDD.n2520 10.6151
R21081 VDD.n2522 VDD.n2521 10.6151
R21082 VDD.n2522 VDD.n956 10.6151
R21083 VDD.n2532 VDD.n956 10.6151
R21084 VDD.n2533 VDD.n2532 10.6151
R21085 VDD.n2534 VDD.n2533 10.6151
R21086 VDD.n2534 VDD.n943 10.6151
R21087 VDD.n2544 VDD.n943 10.6151
R21088 VDD.n2545 VDD.n2544 10.6151
R21089 VDD.n2546 VDD.n2545 10.6151
R21090 VDD.n2546 VDD.n932 10.6151
R21091 VDD.n2556 VDD.n932 10.6151
R21092 VDD.n2557 VDD.n2556 10.6151
R21093 VDD.n2558 VDD.n2557 10.6151
R21094 VDD.n2558 VDD.n920 10.6151
R21095 VDD.n2568 VDD.n920 10.6151
R21096 VDD.n2569 VDD.n2568 10.6151
R21097 VDD.n2570 VDD.n2569 10.6151
R21098 VDD.n2570 VDD.n908 10.6151
R21099 VDD.n2580 VDD.n908 10.6151
R21100 VDD.n2581 VDD.n2580 10.6151
R21101 VDD.n2582 VDD.n2581 10.6151
R21102 VDD.n2582 VDD.n896 10.6151
R21103 VDD.n2592 VDD.n896 10.6151
R21104 VDD.n2593 VDD.n2592 10.6151
R21105 VDD.n2594 VDD.n2593 10.6151
R21106 VDD.n2594 VDD.n884 10.6151
R21107 VDD.n2604 VDD.n884 10.6151
R21108 VDD.n2605 VDD.n2604 10.6151
R21109 VDD.n2606 VDD.n2605 10.6151
R21110 VDD.n2606 VDD.n873 10.6151
R21111 VDD.n2616 VDD.n873 10.6151
R21112 VDD.n2617 VDD.n2616 10.6151
R21113 VDD.n2618 VDD.n2617 10.6151
R21114 VDD.n2618 VDD.n861 10.6151
R21115 VDD.n2628 VDD.n861 10.6151
R21116 VDD.n2629 VDD.n2628 10.6151
R21117 VDD.n2630 VDD.n2629 10.6151
R21118 VDD.n2630 VDD.n849 10.6151
R21119 VDD.n2640 VDD.n849 10.6151
R21120 VDD.n2641 VDD.n2640 10.6151
R21121 VDD.n2642 VDD.n2641 10.6151
R21122 VDD.n2642 VDD.n837 10.6151
R21123 VDD.n2652 VDD.n837 10.6151
R21124 VDD.n2653 VDD.n2652 10.6151
R21125 VDD.n2654 VDD.n2653 10.6151
R21126 VDD.n2654 VDD.n825 10.6151
R21127 VDD.n2664 VDD.n825 10.6151
R21128 VDD.n2665 VDD.n2664 10.6151
R21129 VDD.n2666 VDD.n2665 10.6151
R21130 VDD.n2666 VDD.n813 10.6151
R21131 VDD.n2676 VDD.n813 10.6151
R21132 VDD.n2677 VDD.n2676 10.6151
R21133 VDD.n2678 VDD.n2677 10.6151
R21134 VDD.n2678 VDD.n801 10.6151
R21135 VDD.n2688 VDD.n801 10.6151
R21136 VDD.n2689 VDD.n2688 10.6151
R21137 VDD.n2690 VDD.n2689 10.6151
R21138 VDD.n2690 VDD.n789 10.6151
R21139 VDD.n2700 VDD.n789 10.6151
R21140 VDD.n2701 VDD.n2700 10.6151
R21141 VDD.n2702 VDD.n2701 10.6151
R21142 VDD.n2702 VDD.n777 10.6151
R21143 VDD.n2712 VDD.n777 10.6151
R21144 VDD.n2713 VDD.n2712 10.6151
R21145 VDD.n2714 VDD.n2713 10.6151
R21146 VDD.n2714 VDD.n764 10.6151
R21147 VDD.n2724 VDD.n764 10.6151
R21148 VDD.n2725 VDD.n2724 10.6151
R21149 VDD.n2726 VDD.n2725 10.6151
R21150 VDD.n2726 VDD.n753 10.6151
R21151 VDD.n2736 VDD.n753 10.6151
R21152 VDD.n2737 VDD.n2736 10.6151
R21153 VDD.n2738 VDD.n2737 10.6151
R21154 VDD.n2738 VDD.n741 10.6151
R21155 VDD.n2748 VDD.n741 10.6151
R21156 VDD.n2749 VDD.n2748 10.6151
R21157 VDD.n2750 VDD.n2749 10.6151
R21158 VDD.n2750 VDD.n729 10.6151
R21159 VDD.n2760 VDD.n729 10.6151
R21160 VDD.n2761 VDD.n2760 10.6151
R21161 VDD.n2762 VDD.n2761 10.6151
R21162 VDD.n2762 VDD.n717 10.6151
R21163 VDD.n2772 VDD.n717 10.6151
R21164 VDD.n2773 VDD.n2772 10.6151
R21165 VDD.n2774 VDD.n2773 10.6151
R21166 VDD.n2774 VDD.n705 10.6151
R21167 VDD.n2784 VDD.n705 10.6151
R21168 VDD.n2785 VDD.n2784 10.6151
R21169 VDD.n2786 VDD.n2785 10.6151
R21170 VDD.n2786 VDD.n694 10.6151
R21171 VDD.n2796 VDD.n694 10.6151
R21172 VDD.n2797 VDD.n2796 10.6151
R21173 VDD.n2798 VDD.n2797 10.6151
R21174 VDD.n2798 VDD.n681 10.6151
R21175 VDD.n2813 VDD.n681 10.6151
R21176 VDD.n2814 VDD.n2813 10.6151
R21177 VDD.n2815 VDD.n2814 10.6151
R21178 VDD.n2815 VDD.n671 10.6151
R21179 VDD.n2861 VDD.n671 10.6151
R21180 VDD.n2861 VDD.n2860 10.6151
R21181 VDD.n3389 VDD.n3387 10.6151
R21182 VDD.n3387 VDD.n3386 10.6151
R21183 VDD.n3386 VDD.n3384 10.6151
R21184 VDD.n3384 VDD.n3383 10.6151
R21185 VDD.n3383 VDD.n3381 10.6151
R21186 VDD.n3381 VDD.n3380 10.6151
R21187 VDD.n3380 VDD.n3378 10.6151
R21188 VDD.n3378 VDD.n3377 10.6151
R21189 VDD.n3377 VDD.n3375 10.6151
R21190 VDD.n3375 VDD.n3374 10.6151
R21191 VDD.n3374 VDD.n3372 10.6151
R21192 VDD.n3372 VDD.n3371 10.6151
R21193 VDD.n3371 VDD.n3116 10.6151
R21194 VDD.n3116 VDD.n3115 10.6151
R21195 VDD.n3115 VDD.n3113 10.6151
R21196 VDD.n3113 VDD.n3112 10.6151
R21197 VDD.n3112 VDD.n3110 10.6151
R21198 VDD.n3110 VDD.n3109 10.6151
R21199 VDD.n3109 VDD.n3107 10.6151
R21200 VDD.n3107 VDD.n3106 10.6151
R21201 VDD.n3106 VDD.n3104 10.6151
R21202 VDD.n3104 VDD.n3103 10.6151
R21203 VDD.n3103 VDD.n3101 10.6151
R21204 VDD.n3101 VDD.n3100 10.6151
R21205 VDD.n3100 VDD.n3098 10.6151
R21206 VDD.n3098 VDD.n3097 10.6151
R21207 VDD.n3097 VDD.n3095 10.6151
R21208 VDD.n3095 VDD.n3094 10.6151
R21209 VDD.n3094 VDD.n3092 10.6151
R21210 VDD.n3092 VDD.n3091 10.6151
R21211 VDD.n3091 VDD.n3089 10.6151
R21212 VDD.n3089 VDD.n3088 10.6151
R21213 VDD.n3088 VDD.n3086 10.6151
R21214 VDD.n3086 VDD.n3085 10.6151
R21215 VDD.n3085 VDD.n3083 10.6151
R21216 VDD.n3083 VDD.n3082 10.6151
R21217 VDD.n3082 VDD.n3080 10.6151
R21218 VDD.n3080 VDD.n3079 10.6151
R21219 VDD.n3079 VDD.n3077 10.6151
R21220 VDD.n3077 VDD.n3076 10.6151
R21221 VDD.n3076 VDD.n3074 10.6151
R21222 VDD.n3074 VDD.n3073 10.6151
R21223 VDD.n3073 VDD.n3071 10.6151
R21224 VDD.n3071 VDD.n3070 10.6151
R21225 VDD.n3070 VDD.n3068 10.6151
R21226 VDD.n3068 VDD.n3067 10.6151
R21227 VDD.n3067 VDD.n3065 10.6151
R21228 VDD.n3065 VDD.n3064 10.6151
R21229 VDD.n3064 VDD.n3062 10.6151
R21230 VDD.n3062 VDD.n3061 10.6151
R21231 VDD.n3061 VDD.n3059 10.6151
R21232 VDD.n3059 VDD.n3058 10.6151
R21233 VDD.n3058 VDD.n3056 10.6151
R21234 VDD.n3056 VDD.n3055 10.6151
R21235 VDD.n3055 VDD.n3053 10.6151
R21236 VDD.n3053 VDD.n3052 10.6151
R21237 VDD.n3052 VDD.n3050 10.6151
R21238 VDD.n3050 VDD.n3049 10.6151
R21239 VDD.n3049 VDD.n3047 10.6151
R21240 VDD.n3047 VDD.n3046 10.6151
R21241 VDD.n3046 VDD.n3044 10.6151
R21242 VDD.n3044 VDD.n3043 10.6151
R21243 VDD.n3043 VDD.n3041 10.6151
R21244 VDD.n3041 VDD.n3040 10.6151
R21245 VDD.n3040 VDD.n3038 10.6151
R21246 VDD.n3038 VDD.n3037 10.6151
R21247 VDD.n3037 VDD.n3035 10.6151
R21248 VDD.n3035 VDD.n3034 10.6151
R21249 VDD.n3034 VDD.n3032 10.6151
R21250 VDD.n3032 VDD.n3031 10.6151
R21251 VDD.n3031 VDD.n3029 10.6151
R21252 VDD.n3029 VDD.n3028 10.6151
R21253 VDD.n3028 VDD.n3026 10.6151
R21254 VDD.n3026 VDD.n3025 10.6151
R21255 VDD.n3025 VDD.n3023 10.6151
R21256 VDD.n3023 VDD.n3022 10.6151
R21257 VDD.n3022 VDD.n3020 10.6151
R21258 VDD.n3020 VDD.n3019 10.6151
R21259 VDD.n3019 VDD.n3017 10.6151
R21260 VDD.n3017 VDD.n3016 10.6151
R21261 VDD.n3016 VDD.n3014 10.6151
R21262 VDD.n3014 VDD.n3013 10.6151
R21263 VDD.n3013 VDD.n3011 10.6151
R21264 VDD.n3011 VDD.n3010 10.6151
R21265 VDD.n3010 VDD.n3008 10.6151
R21266 VDD.n3008 VDD.n3007 10.6151
R21267 VDD.n3007 VDD.n3005 10.6151
R21268 VDD.n3005 VDD.n3004 10.6151
R21269 VDD.n3004 VDD.n3002 10.6151
R21270 VDD.n3002 VDD.n3001 10.6151
R21271 VDD.n3001 VDD.n2999 10.6151
R21272 VDD.n2999 VDD.n2998 10.6151
R21273 VDD.n2998 VDD.n2996 10.6151
R21274 VDD.n2996 VDD.n2995 10.6151
R21275 VDD.n2995 VDD.n2993 10.6151
R21276 VDD.n2993 VDD.n2992 10.6151
R21277 VDD.n2992 VDD.n2990 10.6151
R21278 VDD.n2990 VDD.n2989 10.6151
R21279 VDD.n2989 VDD.n2987 10.6151
R21280 VDD.n2987 VDD.n2986 10.6151
R21281 VDD.n2986 VDD.n2984 10.6151
R21282 VDD.n2984 VDD.n2983 10.6151
R21283 VDD.n2983 VDD.n2981 10.6151
R21284 VDD.n2981 VDD.n2980 10.6151
R21285 VDD.n2980 VDD.n2978 10.6151
R21286 VDD.n2978 VDD.n2977 10.6151
R21287 VDD.n2977 VDD.n2975 10.6151
R21288 VDD.n2975 VDD.n2974 10.6151
R21289 VDD.n2974 VDD.n2972 10.6151
R21290 VDD.n2972 VDD.n2971 10.6151
R21291 VDD.n2971 VDD.n2969 10.6151
R21292 VDD.n2969 VDD.n2968 10.6151
R21293 VDD.n2968 VDD.n2966 10.6151
R21294 VDD.n2966 VDD.n2965 10.6151
R21295 VDD.n2965 VDD.n2963 10.6151
R21296 VDD.n2963 VDD.n2962 10.6151
R21297 VDD.n2962 VDD.n2960 10.6151
R21298 VDD.n2960 VDD.n2959 10.6151
R21299 VDD.n2959 VDD.n2957 10.6151
R21300 VDD.n2957 VDD.n2956 10.6151
R21301 VDD.n2956 VDD.n2954 10.6151
R21302 VDD.n2954 VDD.n2953 10.6151
R21303 VDD.n2953 VDD.n2951 10.6151
R21304 VDD.n2951 VDD.n2950 10.6151
R21305 VDD.n2950 VDD.n2948 10.6151
R21306 VDD.n2948 VDD.n2947 10.6151
R21307 VDD.n2947 VDD.n2945 10.6151
R21308 VDD.n2945 VDD.n2944 10.6151
R21309 VDD.n2944 VDD.n2942 10.6151
R21310 VDD.n2942 VDD.n2941 10.6151
R21311 VDD.n2941 VDD.n2939 10.6151
R21312 VDD.n2939 VDD.n2938 10.6151
R21313 VDD.n2938 VDD.n2936 10.6151
R21314 VDD.n2936 VDD.n2935 10.6151
R21315 VDD.n2935 VDD.n2933 10.6151
R21316 VDD.n2933 VDD.n2932 10.6151
R21317 VDD.n2932 VDD.n2930 10.6151
R21318 VDD.n2930 VDD.n2929 10.6151
R21319 VDD.n2929 VDD.n2927 10.6151
R21320 VDD.n2927 VDD.n2926 10.6151
R21321 VDD.n2926 VDD.n2924 10.6151
R21322 VDD.n2924 VDD.n2923 10.6151
R21323 VDD.n2923 VDD.n207 10.6151
R21324 VDD.n3887 VDD.n207 10.6151
R21325 VDD.n3888 VDD.n3887 10.6151
R21326 VDD.n3422 VDD.n3421 10.6151
R21327 VDD.n3421 VDD.n3420 10.6151
R21328 VDD.n3420 VDD.n3419 10.6151
R21329 VDD.n3419 VDD.n3417 10.6151
R21330 VDD.n3417 VDD.n3414 10.6151
R21331 VDD.n3414 VDD.n3413 10.6151
R21332 VDD.n3413 VDD.n3410 10.6151
R21333 VDD.n3410 VDD.n3409 10.6151
R21334 VDD.n3409 VDD.n3406 10.6151
R21335 VDD.n3406 VDD.n3405 10.6151
R21336 VDD.n3405 VDD.n3402 10.6151
R21337 VDD.n3402 VDD.n3401 10.6151
R21338 VDD.n3401 VDD.n3398 10.6151
R21339 VDD.n3396 VDD.n3393 10.6151
R21340 VDD.n3393 VDD.n3392 10.6151
R21341 VDD.n3392 VDD.n3390 10.6151
R21342 VDD.n3434 VDD.n632 10.6151
R21343 VDD.n3435 VDD.n3434 10.6151
R21344 VDD.n3436 VDD.n3435 10.6151
R21345 VDD.n3436 VDD.n620 10.6151
R21346 VDD.n3446 VDD.n620 10.6151
R21347 VDD.n3447 VDD.n3446 10.6151
R21348 VDD.n3448 VDD.n3447 10.6151
R21349 VDD.n3448 VDD.n608 10.6151
R21350 VDD.n3458 VDD.n608 10.6151
R21351 VDD.n3459 VDD.n3458 10.6151
R21352 VDD.n3460 VDD.n3459 10.6151
R21353 VDD.n3460 VDD.n597 10.6151
R21354 VDD.n3470 VDD.n597 10.6151
R21355 VDD.n3471 VDD.n3470 10.6151
R21356 VDD.n3472 VDD.n3471 10.6151
R21357 VDD.n3472 VDD.n585 10.6151
R21358 VDD.n3482 VDD.n585 10.6151
R21359 VDD.n3483 VDD.n3482 10.6151
R21360 VDD.n3484 VDD.n3483 10.6151
R21361 VDD.n3484 VDD.n573 10.6151
R21362 VDD.n3494 VDD.n573 10.6151
R21363 VDD.n3495 VDD.n3494 10.6151
R21364 VDD.n3496 VDD.n3495 10.6151
R21365 VDD.n3496 VDD.n561 10.6151
R21366 VDD.n3506 VDD.n561 10.6151
R21367 VDD.n3507 VDD.n3506 10.6151
R21368 VDD.n3508 VDD.n3507 10.6151
R21369 VDD.n3508 VDD.n549 10.6151
R21370 VDD.n3518 VDD.n549 10.6151
R21371 VDD.n3519 VDD.n3518 10.6151
R21372 VDD.n3520 VDD.n3519 10.6151
R21373 VDD.n3520 VDD.n536 10.6151
R21374 VDD.n3530 VDD.n536 10.6151
R21375 VDD.n3531 VDD.n3530 10.6151
R21376 VDD.n3532 VDD.n3531 10.6151
R21377 VDD.n3532 VDD.n525 10.6151
R21378 VDD.n3542 VDD.n525 10.6151
R21379 VDD.n3543 VDD.n3542 10.6151
R21380 VDD.n3544 VDD.n3543 10.6151
R21381 VDD.n3544 VDD.n513 10.6151
R21382 VDD.n3554 VDD.n513 10.6151
R21383 VDD.n3555 VDD.n3554 10.6151
R21384 VDD.n3556 VDD.n3555 10.6151
R21385 VDD.n3556 VDD.n501 10.6151
R21386 VDD.n3566 VDD.n501 10.6151
R21387 VDD.n3567 VDD.n3566 10.6151
R21388 VDD.n3568 VDD.n3567 10.6151
R21389 VDD.n3568 VDD.n488 10.6151
R21390 VDD.n3578 VDD.n488 10.6151
R21391 VDD.n3579 VDD.n3578 10.6151
R21392 VDD.n3580 VDD.n3579 10.6151
R21393 VDD.n3580 VDD.n477 10.6151
R21394 VDD.n3590 VDD.n477 10.6151
R21395 VDD.n3591 VDD.n3590 10.6151
R21396 VDD.n3592 VDD.n3591 10.6151
R21397 VDD.n3592 VDD.n465 10.6151
R21398 VDD.n3602 VDD.n465 10.6151
R21399 VDD.n3603 VDD.n3602 10.6151
R21400 VDD.n3604 VDD.n3603 10.6151
R21401 VDD.n3604 VDD.n453 10.6151
R21402 VDD.n3614 VDD.n453 10.6151
R21403 VDD.n3615 VDD.n3614 10.6151
R21404 VDD.n3616 VDD.n3615 10.6151
R21405 VDD.n3616 VDD.n441 10.6151
R21406 VDD.n3626 VDD.n441 10.6151
R21407 VDD.n3627 VDD.n3626 10.6151
R21408 VDD.n3628 VDD.n3627 10.6151
R21409 VDD.n3628 VDD.n429 10.6151
R21410 VDD.n3638 VDD.n429 10.6151
R21411 VDD.n3639 VDD.n3638 10.6151
R21412 VDD.n3640 VDD.n3639 10.6151
R21413 VDD.n3640 VDD.n418 10.6151
R21414 VDD.n3650 VDD.n418 10.6151
R21415 VDD.n3651 VDD.n3650 10.6151
R21416 VDD.n3652 VDD.n3651 10.6151
R21417 VDD.n3652 VDD.n406 10.6151
R21418 VDD.n3662 VDD.n406 10.6151
R21419 VDD.n3663 VDD.n3662 10.6151
R21420 VDD.n3664 VDD.n3663 10.6151
R21421 VDD.n3664 VDD.n394 10.6151
R21422 VDD.n3674 VDD.n394 10.6151
R21423 VDD.n3675 VDD.n3674 10.6151
R21424 VDD.n3676 VDD.n3675 10.6151
R21425 VDD.n3676 VDD.n382 10.6151
R21426 VDD.n3686 VDD.n382 10.6151
R21427 VDD.n3687 VDD.n3686 10.6151
R21428 VDD.n3688 VDD.n3687 10.6151
R21429 VDD.n3688 VDD.n370 10.6151
R21430 VDD.n3698 VDD.n370 10.6151
R21431 VDD.n3699 VDD.n3698 10.6151
R21432 VDD.n3700 VDD.n3699 10.6151
R21433 VDD.n3700 VDD.n358 10.6151
R21434 VDD.n3710 VDD.n358 10.6151
R21435 VDD.n3711 VDD.n3710 10.6151
R21436 VDD.n3712 VDD.n3711 10.6151
R21437 VDD.n3712 VDD.n345 10.6151
R21438 VDD.n3722 VDD.n345 10.6151
R21439 VDD.n3723 VDD.n3722 10.6151
R21440 VDD.n3724 VDD.n3723 10.6151
R21441 VDD.n3724 VDD.n334 10.6151
R21442 VDD.n3734 VDD.n334 10.6151
R21443 VDD.n3735 VDD.n3734 10.6151
R21444 VDD.n3736 VDD.n3735 10.6151
R21445 VDD.n3736 VDD.n322 10.6151
R21446 VDD.n3746 VDD.n322 10.6151
R21447 VDD.n3747 VDD.n3746 10.6151
R21448 VDD.n3748 VDD.n3747 10.6151
R21449 VDD.n3748 VDD.n309 10.6151
R21450 VDD.n3758 VDD.n309 10.6151
R21451 VDD.n3759 VDD.n3758 10.6151
R21452 VDD.n3760 VDD.n3759 10.6151
R21453 VDD.n3760 VDD.n298 10.6151
R21454 VDD.n3770 VDD.n298 10.6151
R21455 VDD.n3771 VDD.n3770 10.6151
R21456 VDD.n3772 VDD.n3771 10.6151
R21457 VDD.n3772 VDD.n286 10.6151
R21458 VDD.n3782 VDD.n286 10.6151
R21459 VDD.n3783 VDD.n3782 10.6151
R21460 VDD.n3784 VDD.n3783 10.6151
R21461 VDD.n3784 VDD.n274 10.6151
R21462 VDD.n3794 VDD.n274 10.6151
R21463 VDD.n3795 VDD.n3794 10.6151
R21464 VDD.n3796 VDD.n3795 10.6151
R21465 VDD.n3796 VDD.n262 10.6151
R21466 VDD.n3806 VDD.n262 10.6151
R21467 VDD.n3807 VDD.n3806 10.6151
R21468 VDD.n3808 VDD.n3807 10.6151
R21469 VDD.n3808 VDD.n250 10.6151
R21470 VDD.n3818 VDD.n250 10.6151
R21471 VDD.n3819 VDD.n3818 10.6151
R21472 VDD.n3820 VDD.n3819 10.6151
R21473 VDD.n3820 VDD.n238 10.6151
R21474 VDD.n3830 VDD.n238 10.6151
R21475 VDD.n3831 VDD.n3830 10.6151
R21476 VDD.n3832 VDD.n3831 10.6151
R21477 VDD.n3832 VDD.n226 10.6151
R21478 VDD.n3842 VDD.n226 10.6151
R21479 VDD.n3843 VDD.n3842 10.6151
R21480 VDD.n3844 VDD.n3843 10.6151
R21481 VDD.n3844 VDD.n213 10.6151
R21482 VDD.n3880 VDD.n213 10.6151
R21483 VDD.n3881 VDD.n3880 10.6151
R21484 VDD.n3882 VDD.n3881 10.6151
R21485 VDD.n3882 VDD.n191 10.6151
R21486 VDD.n3923 VDD.n191 10.6151
R21487 VDD.n3922 VDD.n3921 10.6151
R21488 VDD.n3921 VDD.n192 10.6151
R21489 VDD.n3916 VDD.n192 10.6151
R21490 VDD.n3916 VDD.n3915 10.6151
R21491 VDD.n3915 VDD.n3914 10.6151
R21492 VDD.n3914 VDD.n195 10.6151
R21493 VDD.n3909 VDD.n195 10.6151
R21494 VDD.n3909 VDD.n3908 10.6151
R21495 VDD.n3905 VDD.n198 10.6151
R21496 VDD.n3900 VDD.n198 10.6151
R21497 VDD.n3900 VDD.n3899 10.6151
R21498 VDD.n3899 VDD.n3898 10.6151
R21499 VDD.n3893 VDD.n205 10.6151
R21500 VDD.n3893 VDD.n3892 10.6151
R21501 VDD.n3892 VDD.n3891 10.6151
R21502 VDD.n3870 VDD.n3850 10.6151
R21503 VDD.n3851 VDD.n3850 10.6151
R21504 VDD.n3863 VDD.n3851 10.6151
R21505 VDD.n3863 VDD.n3862 10.6151
R21506 VDD.n3862 VDD.n3861 10.6151
R21507 VDD.n3861 VDD.n3853 10.6151
R21508 VDD.n3856 VDD.n3853 10.6151
R21509 VDD.n3856 VDD.n172 10.6151
R21510 VDD.n3942 VDD.n173 10.6151
R21511 VDD.n3937 VDD.n173 10.6151
R21512 VDD.n3937 VDD.n3936 10.6151
R21513 VDD.n3936 VDD.n3935 10.6151
R21514 VDD.n3930 VDD.n181 10.6151
R21515 VDD.n3930 VDD.n3929 10.6151
R21516 VDD.n3929 VDD.n3928 10.6151
R21517 VDD.n3154 VDD.n3153 10.6151
R21518 VDD.n3156 VDD.n3154 10.6151
R21519 VDD.n3157 VDD.n3156 10.6151
R21520 VDD.n3159 VDD.n3157 10.6151
R21521 VDD.n3160 VDD.n3159 10.6151
R21522 VDD.n3162 VDD.n3160 10.6151
R21523 VDD.n3163 VDD.n3162 10.6151
R21524 VDD.n3165 VDD.n3163 10.6151
R21525 VDD.n3166 VDD.n3165 10.6151
R21526 VDD.n3168 VDD.n3166 10.6151
R21527 VDD.n3169 VDD.n3168 10.6151
R21528 VDD.n3367 VDD.n3169 10.6151
R21529 VDD.n3367 VDD.n3366 10.6151
R21530 VDD.n3366 VDD.n3365 10.6151
R21531 VDD.n3365 VDD.n3363 10.6151
R21532 VDD.n3363 VDD.n3362 10.6151
R21533 VDD.n3362 VDD.n3360 10.6151
R21534 VDD.n3360 VDD.n3359 10.6151
R21535 VDD.n3359 VDD.n3357 10.6151
R21536 VDD.n3357 VDD.n3356 10.6151
R21537 VDD.n3356 VDD.n3354 10.6151
R21538 VDD.n3354 VDD.n3353 10.6151
R21539 VDD.n3353 VDD.n3351 10.6151
R21540 VDD.n3351 VDD.n3350 10.6151
R21541 VDD.n3350 VDD.n3348 10.6151
R21542 VDD.n3348 VDD.n3347 10.6151
R21543 VDD.n3347 VDD.n3345 10.6151
R21544 VDD.n3345 VDD.n3344 10.6151
R21545 VDD.n3344 VDD.n3342 10.6151
R21546 VDD.n3342 VDD.n3341 10.6151
R21547 VDD.n3341 VDD.n3339 10.6151
R21548 VDD.n3339 VDD.n3338 10.6151
R21549 VDD.n3338 VDD.n3336 10.6151
R21550 VDD.n3336 VDD.n3335 10.6151
R21551 VDD.n3335 VDD.n3333 10.6151
R21552 VDD.n3333 VDD.n3332 10.6151
R21553 VDD.n3332 VDD.n3330 10.6151
R21554 VDD.n3330 VDD.n3329 10.6151
R21555 VDD.n3329 VDD.n3327 10.6151
R21556 VDD.n3327 VDD.n3326 10.6151
R21557 VDD.n3326 VDD.n3324 10.6151
R21558 VDD.n3324 VDD.n3323 10.6151
R21559 VDD.n3323 VDD.n3321 10.6151
R21560 VDD.n3321 VDD.n3320 10.6151
R21561 VDD.n3320 VDD.n3318 10.6151
R21562 VDD.n3318 VDD.n3317 10.6151
R21563 VDD.n3317 VDD.n3315 10.6151
R21564 VDD.n3315 VDD.n3314 10.6151
R21565 VDD.n3314 VDD.n3312 10.6151
R21566 VDD.n3312 VDD.n3311 10.6151
R21567 VDD.n3311 VDD.n3309 10.6151
R21568 VDD.n3309 VDD.n3308 10.6151
R21569 VDD.n3308 VDD.n3306 10.6151
R21570 VDD.n3306 VDD.n3305 10.6151
R21571 VDD.n3305 VDD.n3303 10.6151
R21572 VDD.n3303 VDD.n3302 10.6151
R21573 VDD.n3302 VDD.n3300 10.6151
R21574 VDD.n3300 VDD.n3299 10.6151
R21575 VDD.n3299 VDD.n3297 10.6151
R21576 VDD.n3297 VDD.n3296 10.6151
R21577 VDD.n3296 VDD.n3294 10.6151
R21578 VDD.n3294 VDD.n3293 10.6151
R21579 VDD.n3293 VDD.n3291 10.6151
R21580 VDD.n3291 VDD.n3290 10.6151
R21581 VDD.n3290 VDD.n3288 10.6151
R21582 VDD.n3288 VDD.n3287 10.6151
R21583 VDD.n3287 VDD.n3285 10.6151
R21584 VDD.n3285 VDD.n3284 10.6151
R21585 VDD.n3284 VDD.n3282 10.6151
R21586 VDD.n3282 VDD.n3281 10.6151
R21587 VDD.n3281 VDD.n3279 10.6151
R21588 VDD.n3279 VDD.n3278 10.6151
R21589 VDD.n3278 VDD.n3276 10.6151
R21590 VDD.n3276 VDD.n3275 10.6151
R21591 VDD.n3275 VDD.n3273 10.6151
R21592 VDD.n3273 VDD.n3272 10.6151
R21593 VDD.n3272 VDD.n3270 10.6151
R21594 VDD.n3270 VDD.n3269 10.6151
R21595 VDD.n3269 VDD.n3267 10.6151
R21596 VDD.n3267 VDD.n3266 10.6151
R21597 VDD.n3266 VDD.n3264 10.6151
R21598 VDD.n3264 VDD.n3263 10.6151
R21599 VDD.n3263 VDD.n3261 10.6151
R21600 VDD.n3261 VDD.n3260 10.6151
R21601 VDD.n3260 VDD.n3258 10.6151
R21602 VDD.n3258 VDD.n3257 10.6151
R21603 VDD.n3257 VDD.n3255 10.6151
R21604 VDD.n3255 VDD.n3254 10.6151
R21605 VDD.n3254 VDD.n3252 10.6151
R21606 VDD.n3252 VDD.n3251 10.6151
R21607 VDD.n3251 VDD.n3249 10.6151
R21608 VDD.n3249 VDD.n3248 10.6151
R21609 VDD.n3248 VDD.n3246 10.6151
R21610 VDD.n3246 VDD.n3245 10.6151
R21611 VDD.n3245 VDD.n3243 10.6151
R21612 VDD.n3243 VDD.n3242 10.6151
R21613 VDD.n3242 VDD.n3240 10.6151
R21614 VDD.n3240 VDD.n3239 10.6151
R21615 VDD.n3239 VDD.n3237 10.6151
R21616 VDD.n3237 VDD.n3236 10.6151
R21617 VDD.n3236 VDD.n3234 10.6151
R21618 VDD.n3234 VDD.n3233 10.6151
R21619 VDD.n3233 VDD.n3231 10.6151
R21620 VDD.n3231 VDD.n3230 10.6151
R21621 VDD.n3230 VDD.n3228 10.6151
R21622 VDD.n3228 VDD.n3227 10.6151
R21623 VDD.n3227 VDD.n3225 10.6151
R21624 VDD.n3225 VDD.n3224 10.6151
R21625 VDD.n3224 VDD.n3222 10.6151
R21626 VDD.n3222 VDD.n3221 10.6151
R21627 VDD.n3221 VDD.n3219 10.6151
R21628 VDD.n3219 VDD.n3218 10.6151
R21629 VDD.n3218 VDD.n3216 10.6151
R21630 VDD.n3216 VDD.n3215 10.6151
R21631 VDD.n3215 VDD.n3213 10.6151
R21632 VDD.n3213 VDD.n3212 10.6151
R21633 VDD.n3212 VDD.n3210 10.6151
R21634 VDD.n3210 VDD.n3209 10.6151
R21635 VDD.n3209 VDD.n3207 10.6151
R21636 VDD.n3207 VDD.n3206 10.6151
R21637 VDD.n3206 VDD.n3204 10.6151
R21638 VDD.n3204 VDD.n3203 10.6151
R21639 VDD.n3203 VDD.n3201 10.6151
R21640 VDD.n3201 VDD.n3200 10.6151
R21641 VDD.n3200 VDD.n3198 10.6151
R21642 VDD.n3198 VDD.n3197 10.6151
R21643 VDD.n3197 VDD.n3195 10.6151
R21644 VDD.n3195 VDD.n3194 10.6151
R21645 VDD.n3194 VDD.n3192 10.6151
R21646 VDD.n3192 VDD.n3191 10.6151
R21647 VDD.n3191 VDD.n3189 10.6151
R21648 VDD.n3189 VDD.n3188 10.6151
R21649 VDD.n3188 VDD.n3186 10.6151
R21650 VDD.n3186 VDD.n3185 10.6151
R21651 VDD.n3185 VDD.n3183 10.6151
R21652 VDD.n3183 VDD.n3182 10.6151
R21653 VDD.n3182 VDD.n3180 10.6151
R21654 VDD.n3180 VDD.n3179 10.6151
R21655 VDD.n3179 VDD.n3177 10.6151
R21656 VDD.n3177 VDD.n3176 10.6151
R21657 VDD.n3176 VDD.n3174 10.6151
R21658 VDD.n3174 VDD.n3173 10.6151
R21659 VDD.n3173 VDD.n3171 10.6151
R21660 VDD.n3171 VDD.n3170 10.6151
R21661 VDD.n3170 VDD.n183 10.6151
R21662 VDD.n3428 VDD.n638 10.6151
R21663 VDD.n3121 VDD.n638 10.6151
R21664 VDD.n3122 VDD.n3121 10.6151
R21665 VDD.n3125 VDD.n3122 10.6151
R21666 VDD.n3126 VDD.n3125 10.6151
R21667 VDD.n3129 VDD.n3126 10.6151
R21668 VDD.n3130 VDD.n3129 10.6151
R21669 VDD.n3133 VDD.n3130 10.6151
R21670 VDD.n3134 VDD.n3133 10.6151
R21671 VDD.n3137 VDD.n3134 10.6151
R21672 VDD.n3138 VDD.n3137 10.6151
R21673 VDD.n3141 VDD.n3138 10.6151
R21674 VDD.n3142 VDD.n3141 10.6151
R21675 VDD.n3146 VDD.n3145 10.6151
R21676 VDD.n3149 VDD.n3146 10.6151
R21677 VDD.n3150 VDD.n3149 10.6151
R21678 VDD.n3430 VDD.n3429 10.6151
R21679 VDD.n3430 VDD.n626 10.6151
R21680 VDD.n3440 VDD.n626 10.6151
R21681 VDD.n3441 VDD.n3440 10.6151
R21682 VDD.n3442 VDD.n3441 10.6151
R21683 VDD.n3442 VDD.n614 10.6151
R21684 VDD.n3452 VDD.n614 10.6151
R21685 VDD.n3453 VDD.n3452 10.6151
R21686 VDD.n3454 VDD.n3453 10.6151
R21687 VDD.n3454 VDD.n602 10.6151
R21688 VDD.n3464 VDD.n602 10.6151
R21689 VDD.n3465 VDD.n3464 10.6151
R21690 VDD.n3466 VDD.n3465 10.6151
R21691 VDD.n3466 VDD.n591 10.6151
R21692 VDD.n3476 VDD.n591 10.6151
R21693 VDD.n3477 VDD.n3476 10.6151
R21694 VDD.n3478 VDD.n3477 10.6151
R21695 VDD.n3478 VDD.n579 10.6151
R21696 VDD.n3488 VDD.n579 10.6151
R21697 VDD.n3489 VDD.n3488 10.6151
R21698 VDD.n3490 VDD.n3489 10.6151
R21699 VDD.n3490 VDD.n567 10.6151
R21700 VDD.n3500 VDD.n567 10.6151
R21701 VDD.n3501 VDD.n3500 10.6151
R21702 VDD.n3502 VDD.n3501 10.6151
R21703 VDD.n3502 VDD.n555 10.6151
R21704 VDD.n3512 VDD.n555 10.6151
R21705 VDD.n3513 VDD.n3512 10.6151
R21706 VDD.n3514 VDD.n3513 10.6151
R21707 VDD.n3514 VDD.n543 10.6151
R21708 VDD.n3524 VDD.n543 10.6151
R21709 VDD.n3525 VDD.n3524 10.6151
R21710 VDD.n3526 VDD.n3525 10.6151
R21711 VDD.n3526 VDD.n531 10.6151
R21712 VDD.n3536 VDD.n531 10.6151
R21713 VDD.n3537 VDD.n3536 10.6151
R21714 VDD.n3538 VDD.n3537 10.6151
R21715 VDD.n3538 VDD.n519 10.6151
R21716 VDD.n3548 VDD.n519 10.6151
R21717 VDD.n3549 VDD.n3548 10.6151
R21718 VDD.n3550 VDD.n3549 10.6151
R21719 VDD.n3550 VDD.n507 10.6151
R21720 VDD.n3560 VDD.n507 10.6151
R21721 VDD.n3561 VDD.n3560 10.6151
R21722 VDD.n3562 VDD.n3561 10.6151
R21723 VDD.n3562 VDD.n495 10.6151
R21724 VDD.n3572 VDD.n495 10.6151
R21725 VDD.n3573 VDD.n3572 10.6151
R21726 VDD.n3574 VDD.n3573 10.6151
R21727 VDD.n3574 VDD.n483 10.6151
R21728 VDD.n3584 VDD.n483 10.6151
R21729 VDD.n3585 VDD.n3584 10.6151
R21730 VDD.n3586 VDD.n3585 10.6151
R21731 VDD.n3586 VDD.n471 10.6151
R21732 VDD.n3596 VDD.n471 10.6151
R21733 VDD.n3597 VDD.n3596 10.6151
R21734 VDD.n3598 VDD.n3597 10.6151
R21735 VDD.n3598 VDD.n459 10.6151
R21736 VDD.n3608 VDD.n459 10.6151
R21737 VDD.n3609 VDD.n3608 10.6151
R21738 VDD.n3610 VDD.n3609 10.6151
R21739 VDD.n3610 VDD.n447 10.6151
R21740 VDD.n3620 VDD.n447 10.6151
R21741 VDD.n3621 VDD.n3620 10.6151
R21742 VDD.n3622 VDD.n3621 10.6151
R21743 VDD.n3622 VDD.n435 10.6151
R21744 VDD.n3632 VDD.n435 10.6151
R21745 VDD.n3633 VDD.n3632 10.6151
R21746 VDD.n3634 VDD.n3633 10.6151
R21747 VDD.n3634 VDD.n423 10.6151
R21748 VDD.n3644 VDD.n423 10.6151
R21749 VDD.n3645 VDD.n3644 10.6151
R21750 VDD.n3646 VDD.n3645 10.6151
R21751 VDD.n3646 VDD.n412 10.6151
R21752 VDD.n3656 VDD.n412 10.6151
R21753 VDD.n3657 VDD.n3656 10.6151
R21754 VDD.n3658 VDD.n3657 10.6151
R21755 VDD.n3658 VDD.n400 10.6151
R21756 VDD.n3668 VDD.n400 10.6151
R21757 VDD.n3669 VDD.n3668 10.6151
R21758 VDD.n3670 VDD.n3669 10.6151
R21759 VDD.n3670 VDD.n388 10.6151
R21760 VDD.n3680 VDD.n388 10.6151
R21761 VDD.n3681 VDD.n3680 10.6151
R21762 VDD.n3682 VDD.n3681 10.6151
R21763 VDD.n3682 VDD.n376 10.6151
R21764 VDD.n3692 VDD.n376 10.6151
R21765 VDD.n3693 VDD.n3692 10.6151
R21766 VDD.n3694 VDD.n3693 10.6151
R21767 VDD.n3694 VDD.n364 10.6151
R21768 VDD.n3704 VDD.n364 10.6151
R21769 VDD.n3705 VDD.n3704 10.6151
R21770 VDD.n3706 VDD.n3705 10.6151
R21771 VDD.n3706 VDD.n352 10.6151
R21772 VDD.n3716 VDD.n352 10.6151
R21773 VDD.n3717 VDD.n3716 10.6151
R21774 VDD.n3718 VDD.n3717 10.6151
R21775 VDD.n3718 VDD.n340 10.6151
R21776 VDD.n3728 VDD.n340 10.6151
R21777 VDD.n3729 VDD.n3728 10.6151
R21778 VDD.n3730 VDD.n3729 10.6151
R21779 VDD.n3730 VDD.n328 10.6151
R21780 VDD.n3740 VDD.n328 10.6151
R21781 VDD.n3741 VDD.n3740 10.6151
R21782 VDD.n3742 VDD.n3741 10.6151
R21783 VDD.n3742 VDD.n316 10.6151
R21784 VDD.n3752 VDD.n316 10.6151
R21785 VDD.n3753 VDD.n3752 10.6151
R21786 VDD.n3754 VDD.n3753 10.6151
R21787 VDD.n3754 VDD.n304 10.6151
R21788 VDD.n3764 VDD.n304 10.6151
R21789 VDD.n3765 VDD.n3764 10.6151
R21790 VDD.n3766 VDD.n3765 10.6151
R21791 VDD.n3766 VDD.n292 10.6151
R21792 VDD.n3776 VDD.n292 10.6151
R21793 VDD.n3777 VDD.n3776 10.6151
R21794 VDD.n3778 VDD.n3777 10.6151
R21795 VDD.n3778 VDD.n280 10.6151
R21796 VDD.n3788 VDD.n280 10.6151
R21797 VDD.n3789 VDD.n3788 10.6151
R21798 VDD.n3790 VDD.n3789 10.6151
R21799 VDD.n3790 VDD.n268 10.6151
R21800 VDD.n3800 VDD.n268 10.6151
R21801 VDD.n3801 VDD.n3800 10.6151
R21802 VDD.n3802 VDD.n3801 10.6151
R21803 VDD.n3802 VDD.n256 10.6151
R21804 VDD.n3812 VDD.n256 10.6151
R21805 VDD.n3813 VDD.n3812 10.6151
R21806 VDD.n3814 VDD.n3813 10.6151
R21807 VDD.n3814 VDD.n244 10.6151
R21808 VDD.n3824 VDD.n244 10.6151
R21809 VDD.n3825 VDD.n3824 10.6151
R21810 VDD.n3826 VDD.n3825 10.6151
R21811 VDD.n3826 VDD.n231 10.6151
R21812 VDD.n3836 VDD.n231 10.6151
R21813 VDD.n3837 VDD.n3836 10.6151
R21814 VDD.n3838 VDD.n3837 10.6151
R21815 VDD.n3838 VDD.n220 10.6151
R21816 VDD.n3848 VDD.n220 10.6151
R21817 VDD.n3849 VDD.n3848 10.6151
R21818 VDD.n3876 VDD.n3849 10.6151
R21819 VDD.n3876 VDD.n3875 10.6151
R21820 VDD.n3875 VDD.n3874 10.6151
R21821 VDD.n3874 VDD.n3873 10.6151
R21822 VDD.n3873 VDD.n3871 10.6151
R21823 VDD.n2384 VDD.n1094 10.6151
R21824 VDD.n2394 VDD.n1094 10.6151
R21825 VDD.n2395 VDD.n2394 10.6151
R21826 VDD.n2396 VDD.n2395 10.6151
R21827 VDD.n2396 VDD.n1082 10.6151
R21828 VDD.n2406 VDD.n1082 10.6151
R21829 VDD.n2407 VDD.n2406 10.6151
R21830 VDD.n2408 VDD.n2407 10.6151
R21831 VDD.n2408 VDD.n1069 10.6151
R21832 VDD.n2418 VDD.n1069 10.6151
R21833 VDD.n2419 VDD.n2418 10.6151
R21834 VDD.n2420 VDD.n2419 10.6151
R21835 VDD.n2420 VDD.n1058 10.6151
R21836 VDD.n2430 VDD.n1058 10.6151
R21837 VDD.n2431 VDD.n2430 10.6151
R21838 VDD.n2432 VDD.n2431 10.6151
R21839 VDD.n2432 VDD.n1046 10.6151
R21840 VDD.n2442 VDD.n1046 10.6151
R21841 VDD.n2443 VDD.n2442 10.6151
R21842 VDD.n2444 VDD.n2443 10.6151
R21843 VDD.n2444 VDD.n1034 10.6151
R21844 VDD.n2454 VDD.n1034 10.6151
R21845 VDD.n2455 VDD.n2454 10.6151
R21846 VDD.n2456 VDD.n2455 10.6151
R21847 VDD.n2456 VDD.n1021 10.6151
R21848 VDD.n2466 VDD.n1021 10.6151
R21849 VDD.n2467 VDD.n2466 10.6151
R21850 VDD.n2468 VDD.n2467 10.6151
R21851 VDD.n2468 VDD.n1010 10.6151
R21852 VDD.n2478 VDD.n1010 10.6151
R21853 VDD.n2479 VDD.n2478 10.6151
R21854 VDD.n2480 VDD.n2479 10.6151
R21855 VDD.n2480 VDD.n998 10.6151
R21856 VDD.n2490 VDD.n998 10.6151
R21857 VDD.n2491 VDD.n2490 10.6151
R21858 VDD.n2492 VDD.n2491 10.6151
R21859 VDD.n2492 VDD.n986 10.6151
R21860 VDD.n2502 VDD.n986 10.6151
R21861 VDD.n2503 VDD.n2502 10.6151
R21862 VDD.n2504 VDD.n2503 10.6151
R21863 VDD.n2504 VDD.n974 10.6151
R21864 VDD.n2514 VDD.n974 10.6151
R21865 VDD.n2515 VDD.n2514 10.6151
R21866 VDD.n2516 VDD.n2515 10.6151
R21867 VDD.n2516 VDD.n962 10.6151
R21868 VDD.n2526 VDD.n962 10.6151
R21869 VDD.n2527 VDD.n2526 10.6151
R21870 VDD.n2528 VDD.n2527 10.6151
R21871 VDD.n2528 VDD.n950 10.6151
R21872 VDD.n2538 VDD.n950 10.6151
R21873 VDD.n2539 VDD.n2538 10.6151
R21874 VDD.n2540 VDD.n2539 10.6151
R21875 VDD.n2540 VDD.n938 10.6151
R21876 VDD.n2550 VDD.n938 10.6151
R21877 VDD.n2551 VDD.n2550 10.6151
R21878 VDD.n2552 VDD.n2551 10.6151
R21879 VDD.n2552 VDD.n926 10.6151
R21880 VDD.n2562 VDD.n926 10.6151
R21881 VDD.n2563 VDD.n2562 10.6151
R21882 VDD.n2564 VDD.n2563 10.6151
R21883 VDD.n2564 VDD.n914 10.6151
R21884 VDD.n2574 VDD.n914 10.6151
R21885 VDD.n2575 VDD.n2574 10.6151
R21886 VDD.n2576 VDD.n2575 10.6151
R21887 VDD.n2576 VDD.n902 10.6151
R21888 VDD.n2586 VDD.n902 10.6151
R21889 VDD.n2587 VDD.n2586 10.6151
R21890 VDD.n2588 VDD.n2587 10.6151
R21891 VDD.n2588 VDD.n890 10.6151
R21892 VDD.n2598 VDD.n890 10.6151
R21893 VDD.n2599 VDD.n2598 10.6151
R21894 VDD.n2600 VDD.n2599 10.6151
R21895 VDD.n2600 VDD.n878 10.6151
R21896 VDD.n2610 VDD.n878 10.6151
R21897 VDD.n2611 VDD.n2610 10.6151
R21898 VDD.n2612 VDD.n2611 10.6151
R21899 VDD.n2612 VDD.n867 10.6151
R21900 VDD.n2622 VDD.n867 10.6151
R21901 VDD.n2623 VDD.n2622 10.6151
R21902 VDD.n2624 VDD.n2623 10.6151
R21903 VDD.n2624 VDD.n855 10.6151
R21904 VDD.n2634 VDD.n855 10.6151
R21905 VDD.n2635 VDD.n2634 10.6151
R21906 VDD.n2636 VDD.n2635 10.6151
R21907 VDD.n2636 VDD.n843 10.6151
R21908 VDD.n2646 VDD.n843 10.6151
R21909 VDD.n2647 VDD.n2646 10.6151
R21910 VDD.n2648 VDD.n2647 10.6151
R21911 VDD.n2648 VDD.n830 10.6151
R21912 VDD.n2658 VDD.n830 10.6151
R21913 VDD.n2659 VDD.n2658 10.6151
R21914 VDD.n2660 VDD.n2659 10.6151
R21915 VDD.n2660 VDD.n819 10.6151
R21916 VDD.n2670 VDD.n819 10.6151
R21917 VDD.n2671 VDD.n2670 10.6151
R21918 VDD.n2672 VDD.n2671 10.6151
R21919 VDD.n2672 VDD.n807 10.6151
R21920 VDD.n2682 VDD.n807 10.6151
R21921 VDD.n2683 VDD.n2682 10.6151
R21922 VDD.n2684 VDD.n2683 10.6151
R21923 VDD.n2684 VDD.n795 10.6151
R21924 VDD.n2694 VDD.n795 10.6151
R21925 VDD.n2695 VDD.n2694 10.6151
R21926 VDD.n2696 VDD.n2695 10.6151
R21927 VDD.n2696 VDD.n783 10.6151
R21928 VDD.n2706 VDD.n783 10.6151
R21929 VDD.n2707 VDD.n2706 10.6151
R21930 VDD.n2708 VDD.n2707 10.6151
R21931 VDD.n2708 VDD.n771 10.6151
R21932 VDD.n2718 VDD.n771 10.6151
R21933 VDD.n2719 VDD.n2718 10.6151
R21934 VDD.n2720 VDD.n2719 10.6151
R21935 VDD.n2720 VDD.n759 10.6151
R21936 VDD.n2730 VDD.n759 10.6151
R21937 VDD.n2731 VDD.n2730 10.6151
R21938 VDD.n2732 VDD.n2731 10.6151
R21939 VDD.n2732 VDD.n747 10.6151
R21940 VDD.n2742 VDD.n747 10.6151
R21941 VDD.n2743 VDD.n2742 10.6151
R21942 VDD.n2744 VDD.n2743 10.6151
R21943 VDD.n2744 VDD.n735 10.6151
R21944 VDD.n2754 VDD.n735 10.6151
R21945 VDD.n2755 VDD.n2754 10.6151
R21946 VDD.n2756 VDD.n2755 10.6151
R21947 VDD.n2756 VDD.n723 10.6151
R21948 VDD.n2766 VDD.n723 10.6151
R21949 VDD.n2767 VDD.n2766 10.6151
R21950 VDD.n2768 VDD.n2767 10.6151
R21951 VDD.n2768 VDD.n711 10.6151
R21952 VDD.n2778 VDD.n711 10.6151
R21953 VDD.n2779 VDD.n2778 10.6151
R21954 VDD.n2780 VDD.n2779 10.6151
R21955 VDD.n2780 VDD.n700 10.6151
R21956 VDD.n2790 VDD.n700 10.6151
R21957 VDD.n2791 VDD.n2790 10.6151
R21958 VDD.n2792 VDD.n2791 10.6151
R21959 VDD.n2792 VDD.n688 10.6151
R21960 VDD.n2802 VDD.n688 10.6151
R21961 VDD.n2803 VDD.n2802 10.6151
R21962 VDD.n2809 VDD.n2803 10.6151
R21963 VDD.n2809 VDD.n2808 10.6151
R21964 VDD.n2808 VDD.n2807 10.6151
R21965 VDD.n2807 VDD.n2806 10.6151
R21966 VDD.n2806 VDD.n2804 10.6151
R21967 VDD.n2804 VDD.n661 10.6151
R21968 VDD.n2900 VDD.n2899 10.6151
R21969 VDD.n2899 VDD.n2898 10.6151
R21970 VDD.n2898 VDD.n2895 10.6151
R21971 VDD.n2895 VDD.n2894 10.6151
R21972 VDD.n2894 VDD.n2891 10.6151
R21973 VDD.n2891 VDD.n2890 10.6151
R21974 VDD.n2890 VDD.n2887 10.6151
R21975 VDD.n2887 VDD.n2886 10.6151
R21976 VDD.n2886 VDD.n2883 10.6151
R21977 VDD.n2883 VDD.n2882 10.6151
R21978 VDD.n2882 VDD.n2879 10.6151
R21979 VDD.n2879 VDD.n2878 10.6151
R21980 VDD.n2878 VDD.n2875 10.6151
R21981 VDD.n2873 VDD.n2870 10.6151
R21982 VDD.n2870 VDD.n2869 10.6151
R21983 VDD.n2869 VDD.n2867 10.6151
R21984 VDD.n2348 VDD.n2347 10.6151
R21985 VDD.n2347 VDD.n2345 10.6151
R21986 VDD.n2345 VDD.n2344 10.6151
R21987 VDD.n2344 VDD.n2342 10.6151
R21988 VDD.n2342 VDD.n2341 10.6151
R21989 VDD.n2341 VDD.n2339 10.6151
R21990 VDD.n2339 VDD.n2338 10.6151
R21991 VDD.n2338 VDD.n2336 10.6151
R21992 VDD.n2336 VDD.n2335 10.6151
R21993 VDD.n2335 VDD.n2333 10.6151
R21994 VDD.n2333 VDD.n2332 10.6151
R21995 VDD.n2332 VDD.n2330 10.6151
R21996 VDD.n2330 VDD.n2329 10.6151
R21997 VDD.n2329 VDD.n2327 10.6151
R21998 VDD.n2327 VDD.n2326 10.6151
R21999 VDD.n2326 VDD.n2324 10.6151
R22000 VDD.n2324 VDD.n2323 10.6151
R22001 VDD.n2323 VDD.n2321 10.6151
R22002 VDD.n2321 VDD.n2320 10.6151
R22003 VDD.n2320 VDD.n2318 10.6151
R22004 VDD.n2318 VDD.n2317 10.6151
R22005 VDD.n2317 VDD.n2315 10.6151
R22006 VDD.n2315 VDD.n2314 10.6151
R22007 VDD.n2314 VDD.n2312 10.6151
R22008 VDD.n2312 VDD.n2311 10.6151
R22009 VDD.n2311 VDD.n2309 10.6151
R22010 VDD.n2309 VDD.n2308 10.6151
R22011 VDD.n2308 VDD.n2306 10.6151
R22012 VDD.n2306 VDD.n2305 10.6151
R22013 VDD.n2305 VDD.n2303 10.6151
R22014 VDD.n2303 VDD.n2302 10.6151
R22015 VDD.n2302 VDD.n2300 10.6151
R22016 VDD.n2300 VDD.n2299 10.6151
R22017 VDD.n2299 VDD.n2297 10.6151
R22018 VDD.n2297 VDD.n2296 10.6151
R22019 VDD.n2296 VDD.n2294 10.6151
R22020 VDD.n2294 VDD.n2293 10.6151
R22021 VDD.n2293 VDD.n2291 10.6151
R22022 VDD.n2291 VDD.n2290 10.6151
R22023 VDD.n2290 VDD.n2288 10.6151
R22024 VDD.n2288 VDD.n2287 10.6151
R22025 VDD.n2287 VDD.n2285 10.6151
R22026 VDD.n2285 VDD.n2284 10.6151
R22027 VDD.n2284 VDD.n2282 10.6151
R22028 VDD.n2282 VDD.n2281 10.6151
R22029 VDD.n2281 VDD.n2279 10.6151
R22030 VDD.n2279 VDD.n2278 10.6151
R22031 VDD.n2278 VDD.n2276 10.6151
R22032 VDD.n2276 VDD.n2275 10.6151
R22033 VDD.n2275 VDD.n2273 10.6151
R22034 VDD.n2273 VDD.n2272 10.6151
R22035 VDD.n2272 VDD.n2270 10.6151
R22036 VDD.n2270 VDD.n2269 10.6151
R22037 VDD.n2269 VDD.n2267 10.6151
R22038 VDD.n2267 VDD.n2266 10.6151
R22039 VDD.n2266 VDD.n2264 10.6151
R22040 VDD.n2264 VDD.n2263 10.6151
R22041 VDD.n2263 VDD.n2261 10.6151
R22042 VDD.n2261 VDD.n2260 10.6151
R22043 VDD.n2260 VDD.n2258 10.6151
R22044 VDD.n2258 VDD.n2257 10.6151
R22045 VDD.n2257 VDD.n2255 10.6151
R22046 VDD.n2255 VDD.n2254 10.6151
R22047 VDD.n2254 VDD.n2252 10.6151
R22048 VDD.n2252 VDD.n2251 10.6151
R22049 VDD.n2251 VDD.n2249 10.6151
R22050 VDD.n2249 VDD.n2248 10.6151
R22051 VDD.n2248 VDD.n2246 10.6151
R22052 VDD.n2246 VDD.n2245 10.6151
R22053 VDD.n2245 VDD.n2243 10.6151
R22054 VDD.n2243 VDD.n2242 10.6151
R22055 VDD.n2242 VDD.n2240 10.6151
R22056 VDD.n2240 VDD.n2239 10.6151
R22057 VDD.n2239 VDD.n2237 10.6151
R22058 VDD.n2237 VDD.n2236 10.6151
R22059 VDD.n2236 VDD.n2234 10.6151
R22060 VDD.n2234 VDD.n2233 10.6151
R22061 VDD.n2233 VDD.n2231 10.6151
R22062 VDD.n2231 VDD.n2230 10.6151
R22063 VDD.n2230 VDD.n2228 10.6151
R22064 VDD.n2228 VDD.n2227 10.6151
R22065 VDD.n2227 VDD.n2225 10.6151
R22066 VDD.n2225 VDD.n2224 10.6151
R22067 VDD.n2224 VDD.n2222 10.6151
R22068 VDD.n2222 VDD.n2221 10.6151
R22069 VDD.n2221 VDD.n2219 10.6151
R22070 VDD.n2219 VDD.n2218 10.6151
R22071 VDD.n2218 VDD.n2216 10.6151
R22072 VDD.n2216 VDD.n2215 10.6151
R22073 VDD.n2215 VDD.n2213 10.6151
R22074 VDD.n2213 VDD.n2212 10.6151
R22075 VDD.n2212 VDD.n2210 10.6151
R22076 VDD.n2210 VDD.n2209 10.6151
R22077 VDD.n2209 VDD.n2207 10.6151
R22078 VDD.n2207 VDD.n2206 10.6151
R22079 VDD.n2206 VDD.n2204 10.6151
R22080 VDD.n2204 VDD.n2203 10.6151
R22081 VDD.n2203 VDD.n2201 10.6151
R22082 VDD.n2201 VDD.n2200 10.6151
R22083 VDD.n2200 VDD.n2198 10.6151
R22084 VDD.n2198 VDD.n2197 10.6151
R22085 VDD.n2197 VDD.n2195 10.6151
R22086 VDD.n2195 VDD.n2194 10.6151
R22087 VDD.n2194 VDD.n2192 10.6151
R22088 VDD.n2192 VDD.n2191 10.6151
R22089 VDD.n2191 VDD.n2189 10.6151
R22090 VDD.n2189 VDD.n2188 10.6151
R22091 VDD.n2188 VDD.n2186 10.6151
R22092 VDD.n2186 VDD.n2185 10.6151
R22093 VDD.n2185 VDD.n2183 10.6151
R22094 VDD.n2183 VDD.n2182 10.6151
R22095 VDD.n2182 VDD.n2180 10.6151
R22096 VDD.n2180 VDD.n2179 10.6151
R22097 VDD.n2179 VDD.n2177 10.6151
R22098 VDD.n2177 VDD.n2176 10.6151
R22099 VDD.n2176 VDD.n2174 10.6151
R22100 VDD.n2174 VDD.n2173 10.6151
R22101 VDD.n2173 VDD.n2171 10.6151
R22102 VDD.n2171 VDD.n2170 10.6151
R22103 VDD.n2170 VDD.n2168 10.6151
R22104 VDD.n2168 VDD.n2167 10.6151
R22105 VDD.n2167 VDD.n2165 10.6151
R22106 VDD.n2165 VDD.n2164 10.6151
R22107 VDD.n2164 VDD.n2162 10.6151
R22108 VDD.n2162 VDD.n2161 10.6151
R22109 VDD.n2161 VDD.n2159 10.6151
R22110 VDD.n2159 VDD.n2158 10.6151
R22111 VDD.n2158 VDD.n2156 10.6151
R22112 VDD.n2156 VDD.n2155 10.6151
R22113 VDD.n2155 VDD.n2153 10.6151
R22114 VDD.n2153 VDD.n2152 10.6151
R22115 VDD.n2152 VDD.n2150 10.6151
R22116 VDD.n2150 VDD.n2149 10.6151
R22117 VDD.n2149 VDD.n1131 10.6151
R22118 VDD.n1131 VDD.n1130 10.6151
R22119 VDD.n1130 VDD.n1128 10.6151
R22120 VDD.n1128 VDD.n1127 10.6151
R22121 VDD.n1127 VDD.n1125 10.6151
R22122 VDD.n1125 VDD.n1124 10.6151
R22123 VDD.n1124 VDD.n1122 10.6151
R22124 VDD.n1122 VDD.n1121 10.6151
R22125 VDD.n1121 VDD.n1119 10.6151
R22126 VDD.n1119 VDD.n1118 10.6151
R22127 VDD.n1118 VDD.n664 10.6151
R22128 VDD.n2866 VDD.n664 10.6151
R22129 VDD.n2383 VDD.n2382 10.6151
R22130 VDD.n2382 VDD.n1106 10.6151
R22131 VDD.n2377 VDD.n1106 10.6151
R22132 VDD.n2377 VDD.n2376 10.6151
R22133 VDD.n2376 VDD.n1108 10.6151
R22134 VDD.n2371 VDD.n1108 10.6151
R22135 VDD.n2371 VDD.n2370 10.6151
R22136 VDD.n2370 VDD.n2369 10.6151
R22137 VDD.n2365 VDD.n2364 10.6151
R22138 VDD.n2364 VDD.n1112 10.6151
R22139 VDD.n2359 VDD.n1112 10.6151
R22140 VDD.n2359 VDD.n2358 10.6151
R22141 VDD.n2356 VDD.n1116 10.6151
R22142 VDD.n2350 VDD.n1116 10.6151
R22143 VDD.n2350 VDD.n2349 10.6151
R22144 VDD.n1895 VDD.n1894 10.4414
R22145 VDD.n3907 VDD.n3906 10.4414
R22146 VDD.n3985 VDD.n3943 10.4414
R22147 VDD.n1823 VDD.n1110 10.4414
R22148 VDD.n1582 VDD.n1581 10.2793
R22149 VDD.n1809 VDD.n1224 10.2793
R22150 VDD.n3966 VDD.n3960 10.2793
R22151 VDD.n4379 VDD.n4365 10.2793
R22152 VDD.n2386 VDD.n1096 10.2285
R22153 VDD.n2392 VDD.n1096 10.2285
R22154 VDD.n2392 VDD.n1090 10.2285
R22155 VDD.n2398 VDD.n1090 10.2285
R22156 VDD.n2398 VDD.n1084 10.2285
R22157 VDD.n2404 VDD.n1084 10.2285
R22158 VDD.n2404 VDD.n1078 10.2285
R22159 VDD.n2410 VDD.n1078 10.2285
R22160 VDD.n2416 VDD.n1071 10.2285
R22161 VDD.n2416 VDD.n1074 10.2285
R22162 VDD.n2422 VDD.n1060 10.2285
R22163 VDD.n2428 VDD.n1060 10.2285
R22164 VDD.n2428 VDD.n1054 10.2285
R22165 VDD.n2434 VDD.n1054 10.2285
R22166 VDD.n2434 VDD.n1048 10.2285
R22167 VDD.n2440 VDD.n1048 10.2285
R22168 VDD.n2440 VDD.n1042 10.2285
R22169 VDD.n2446 VDD.n1042 10.2285
R22170 VDD.n2446 VDD.n1036 10.2285
R22171 VDD.n2452 VDD.n1036 10.2285
R22172 VDD.n2452 VDD.n1030 10.2285
R22173 VDD.n2458 VDD.n1030 10.2285
R22174 VDD.n2458 VDD.n1023 10.2285
R22175 VDD.n2464 VDD.n1023 10.2285
R22176 VDD.n2464 VDD.n1026 10.2285
R22177 VDD.n2470 VDD.n1012 10.2285
R22178 VDD.n2476 VDD.n1012 10.2285
R22179 VDD.n2476 VDD.n1006 10.2285
R22180 VDD.n2482 VDD.n1006 10.2285
R22181 VDD.n2482 VDD.n1000 10.2285
R22182 VDD.n2488 VDD.n1000 10.2285
R22183 VDD.n2494 VDD.n994 10.2285
R22184 VDD.n2494 VDD.n988 10.2285
R22185 VDD.n2500 VDD.n988 10.2285
R22186 VDD.n2500 VDD.n982 10.2285
R22187 VDD.n2506 VDD.n982 10.2285
R22188 VDD.n2506 VDD.n976 10.2285
R22189 VDD.n2512 VDD.n976 10.2285
R22190 VDD.n2512 VDD.n970 10.2285
R22191 VDD.n2518 VDD.n970 10.2285
R22192 VDD.n2518 VDD.n964 10.2285
R22193 VDD.n2524 VDD.n964 10.2285
R22194 VDD.n2530 VDD.n958 10.2285
R22195 VDD.n2530 VDD.n952 10.2285
R22196 VDD.n2536 VDD.n952 10.2285
R22197 VDD.n2536 VDD.n945 10.2285
R22198 VDD.n2542 VDD.n945 10.2285
R22199 VDD.n2542 VDD.n948 10.2285
R22200 VDD.n2548 VDD.n934 10.2285
R22201 VDD.n2554 VDD.n934 10.2285
R22202 VDD.n2554 VDD.n928 10.2285
R22203 VDD.n2560 VDD.n928 10.2285
R22204 VDD.n2560 VDD.n922 10.2285
R22205 VDD.n2566 VDD.n922 10.2285
R22206 VDD.n2566 VDD.n916 10.2285
R22207 VDD.n2572 VDD.n916 10.2285
R22208 VDD.n2572 VDD.n910 10.2285
R22209 VDD.n2578 VDD.n910 10.2285
R22210 VDD.n2578 VDD.n904 10.2285
R22211 VDD.n2584 VDD.n904 10.2285
R22212 VDD.n2584 VDD.n898 10.2285
R22213 VDD.n2590 VDD.n898 10.2285
R22214 VDD.n2590 VDD.n892 10.2285
R22215 VDD.n2596 VDD.n892 10.2285
R22216 VDD.n2596 VDD.n886 10.2285
R22217 VDD.n2602 VDD.n886 10.2285
R22218 VDD.n2608 VDD.n880 10.2285
R22219 VDD.n2608 VDD.t92 10.2285
R22220 VDD.n2614 VDD.t92 10.2285
R22221 VDD.n2614 VDD.n869 10.2285
R22222 VDD.n2620 VDD.n869 10.2285
R22223 VDD.n2620 VDD.n863 10.2285
R22224 VDD.n2626 VDD.n863 10.2285
R22225 VDD.n2626 VDD.n857 10.2285
R22226 VDD.n2632 VDD.n857 10.2285
R22227 VDD.n2632 VDD.n851 10.2285
R22228 VDD.n2638 VDD.n851 10.2285
R22229 VDD.n2638 VDD.n845 10.2285
R22230 VDD.n2644 VDD.n845 10.2285
R22231 VDD.n2644 VDD.n839 10.2285
R22232 VDD.n2650 VDD.n839 10.2285
R22233 VDD.n2650 VDD.n832 10.2285
R22234 VDD.n2656 VDD.n832 10.2285
R22235 VDD.n2656 VDD.n835 10.2285
R22236 VDD.n2662 VDD.n821 10.2285
R22237 VDD.n2668 VDD.n821 10.2285
R22238 VDD.n2674 VDD.n815 10.2285
R22239 VDD.n2674 VDD.n809 10.2285
R22240 VDD.n2680 VDD.n809 10.2285
R22241 VDD.n2680 VDD.n803 10.2285
R22242 VDD.n2686 VDD.n803 10.2285
R22243 VDD.n2686 VDD.n797 10.2285
R22244 VDD.n2692 VDD.n797 10.2285
R22245 VDD.n2692 VDD.n791 10.2285
R22246 VDD.n2698 VDD.n791 10.2285
R22247 VDD.n2698 VDD.n785 10.2285
R22248 VDD.n2704 VDD.n785 10.2285
R22249 VDD.n2704 VDD.n779 10.2285
R22250 VDD.n2710 VDD.n779 10.2285
R22251 VDD.n2710 VDD.n773 10.2285
R22252 VDD.n2716 VDD.n773 10.2285
R22253 VDD.n2722 VDD.n766 10.2285
R22254 VDD.n2722 VDD.n769 10.2285
R22255 VDD.n2728 VDD.n755 10.2285
R22256 VDD.n2734 VDD.n755 10.2285
R22257 VDD.n2734 VDD.n749 10.2285
R22258 VDD.n2740 VDD.n749 10.2285
R22259 VDD.n2740 VDD.n743 10.2285
R22260 VDD.n2746 VDD.n743 10.2285
R22261 VDD.n2746 VDD.n737 10.2285
R22262 VDD.n2752 VDD.n737 10.2285
R22263 VDD.n2752 VDD.n731 10.2285
R22264 VDD.n2758 VDD.n731 10.2285
R22265 VDD.n2758 VDD.n725 10.2285
R22266 VDD.n2764 VDD.n725 10.2285
R22267 VDD.n2764 VDD.n719 10.2285
R22268 VDD.n2770 VDD.n719 10.2285
R22269 VDD.n2770 VDD.n713 10.2285
R22270 VDD.n2776 VDD.n713 10.2285
R22271 VDD.n2776 VDD.n707 10.2285
R22272 VDD.n2782 VDD.n707 10.2285
R22273 VDD.n2788 VDD.n696 10.2285
R22274 VDD.n2794 VDD.n696 10.2285
R22275 VDD.n2794 VDD.n690 10.2285
R22276 VDD.n2800 VDD.n690 10.2285
R22277 VDD.n2800 VDD.n683 10.2285
R22278 VDD.n2811 VDD.n683 10.2285
R22279 VDD.n2811 VDD.n677 10.2285
R22280 VDD.n2817 VDD.n677 10.2285
R22281 VDD.n2817 VDD.n666 10.2285
R22282 VDD.n2863 VDD.n666 10.2285
R22283 VDD.n2863 VDD.n640 10.2285
R22284 VDD.n3432 VDD.n634 10.2285
R22285 VDD.n3432 VDD.n628 10.2285
R22286 VDD.n3438 VDD.n628 10.2285
R22287 VDD.n3438 VDD.n622 10.2285
R22288 VDD.n3444 VDD.n622 10.2285
R22289 VDD.n3444 VDD.n616 10.2285
R22290 VDD.n3450 VDD.n616 10.2285
R22291 VDD.n3450 VDD.n610 10.2285
R22292 VDD.n3456 VDD.n610 10.2285
R22293 VDD.n3456 VDD.n604 10.2285
R22294 VDD.n3462 VDD.n604 10.2285
R22295 VDD.n3468 VDD.n593 10.2285
R22296 VDD.n3474 VDD.n593 10.2285
R22297 VDD.n3474 VDD.n587 10.2285
R22298 VDD.n3480 VDD.n587 10.2285
R22299 VDD.n3480 VDD.n581 10.2285
R22300 VDD.n3486 VDD.n581 10.2285
R22301 VDD.n3486 VDD.n575 10.2285
R22302 VDD.n3492 VDD.n575 10.2285
R22303 VDD.n3492 VDD.n569 10.2285
R22304 VDD.n3498 VDD.n569 10.2285
R22305 VDD.n3498 VDD.n563 10.2285
R22306 VDD.n3504 VDD.n563 10.2285
R22307 VDD.n3504 VDD.n557 10.2285
R22308 VDD.n3510 VDD.n557 10.2285
R22309 VDD.n3510 VDD.n551 10.2285
R22310 VDD.n3516 VDD.n551 10.2285
R22311 VDD.n3516 VDD.n545 10.2285
R22312 VDD.n3522 VDD.n545 10.2285
R22313 VDD.n3528 VDD.n538 10.2285
R22314 VDD.n3528 VDD.n541 10.2285
R22315 VDD.n3534 VDD.n527 10.2285
R22316 VDD.n3540 VDD.n527 10.2285
R22317 VDD.n3540 VDD.n521 10.2285
R22318 VDD.n3546 VDD.n521 10.2285
R22319 VDD.n3546 VDD.n515 10.2285
R22320 VDD.n3552 VDD.n515 10.2285
R22321 VDD.n3552 VDD.n509 10.2285
R22322 VDD.n3558 VDD.n509 10.2285
R22323 VDD.n3558 VDD.n503 10.2285
R22324 VDD.n3564 VDD.n503 10.2285
R22325 VDD.n3564 VDD.n497 10.2285
R22326 VDD.n3570 VDD.n497 10.2285
R22327 VDD.n3570 VDD.n490 10.2285
R22328 VDD.n3576 VDD.n490 10.2285
R22329 VDD.n3576 VDD.n493 10.2285
R22330 VDD.n3582 VDD.n479 10.2285
R22331 VDD.n3588 VDD.n479 10.2285
R22332 VDD.n3594 VDD.n473 10.2285
R22333 VDD.n3594 VDD.n467 10.2285
R22334 VDD.n3600 VDD.n467 10.2285
R22335 VDD.n3600 VDD.n461 10.2285
R22336 VDD.n3606 VDD.n461 10.2285
R22337 VDD.n3606 VDD.n455 10.2285
R22338 VDD.n3612 VDD.n455 10.2285
R22339 VDD.n3612 VDD.n449 10.2285
R22340 VDD.n3618 VDD.n449 10.2285
R22341 VDD.n3618 VDD.n443 10.2285
R22342 VDD.n3624 VDD.n443 10.2285
R22343 VDD.n3624 VDD.n437 10.2285
R22344 VDD.n3630 VDD.n437 10.2285
R22345 VDD.n3630 VDD.n431 10.2285
R22346 VDD.n3636 VDD.n431 10.2285
R22347 VDD.n3636 VDD.t132 10.2285
R22348 VDD.n3642 VDD.t132 10.2285
R22349 VDD.n3642 VDD.n427 10.2285
R22350 VDD.n3648 VDD.n414 10.2285
R22351 VDD.n3654 VDD.n414 10.2285
R22352 VDD.n3654 VDD.n408 10.2285
R22353 VDD.n3660 VDD.n408 10.2285
R22354 VDD.n3660 VDD.n402 10.2285
R22355 VDD.n3666 VDD.n402 10.2285
R22356 VDD.n3666 VDD.n396 10.2285
R22357 VDD.n3672 VDD.n396 10.2285
R22358 VDD.n3672 VDD.n390 10.2285
R22359 VDD.n3678 VDD.n390 10.2285
R22360 VDD.n3678 VDD.n384 10.2285
R22361 VDD.n3684 VDD.n384 10.2285
R22362 VDD.n3684 VDD.n378 10.2285
R22363 VDD.n3690 VDD.n378 10.2285
R22364 VDD.n3690 VDD.n372 10.2285
R22365 VDD.n3696 VDD.n372 10.2285
R22366 VDD.n3696 VDD.n366 10.2285
R22367 VDD.n3702 VDD.n366 10.2285
R22368 VDD.n3708 VDD.n360 10.2285
R22369 VDD.n3708 VDD.n354 10.2285
R22370 VDD.n3714 VDD.n354 10.2285
R22371 VDD.n3714 VDD.n347 10.2285
R22372 VDD.n3720 VDD.n347 10.2285
R22373 VDD.n3720 VDD.n350 10.2285
R22374 VDD.n3726 VDD.n336 10.2285
R22375 VDD.n3732 VDD.n336 10.2285
R22376 VDD.n3732 VDD.n330 10.2285
R22377 VDD.n3738 VDD.n330 10.2285
R22378 VDD.n3738 VDD.n324 10.2285
R22379 VDD.n3744 VDD.n324 10.2285
R22380 VDD.n3744 VDD.n318 10.2285
R22381 VDD.n3750 VDD.n318 10.2285
R22382 VDD.n3750 VDD.n311 10.2285
R22383 VDD.n3756 VDD.n311 10.2285
R22384 VDD.n3756 VDD.n314 10.2285
R22385 VDD.n3762 VDD.n300 10.2285
R22386 VDD.n3768 VDD.n300 10.2285
R22387 VDD.n3768 VDD.n294 10.2285
R22388 VDD.n3774 VDD.n294 10.2285
R22389 VDD.n3774 VDD.n288 10.2285
R22390 VDD.n3780 VDD.n288 10.2285
R22391 VDD.n3786 VDD.n282 10.2285
R22392 VDD.n3786 VDD.n276 10.2285
R22393 VDD.n3792 VDD.n276 10.2285
R22394 VDD.n3792 VDD.n270 10.2285
R22395 VDD.n3798 VDD.n270 10.2285
R22396 VDD.n3798 VDD.n264 10.2285
R22397 VDD.n3804 VDD.n264 10.2285
R22398 VDD.n3804 VDD.n258 10.2285
R22399 VDD.n3810 VDD.n258 10.2285
R22400 VDD.n3810 VDD.n252 10.2285
R22401 VDD.n3816 VDD.n252 10.2285
R22402 VDD.n3816 VDD.n246 10.2285
R22403 VDD.n3822 VDD.n246 10.2285
R22404 VDD.n3822 VDD.n240 10.2285
R22405 VDD.n3828 VDD.n240 10.2285
R22406 VDD.n3834 VDD.n233 10.2285
R22407 VDD.n3834 VDD.n236 10.2285
R22408 VDD.n3840 VDD.n222 10.2285
R22409 VDD.n3846 VDD.n222 10.2285
R22410 VDD.n3846 VDD.n215 10.2285
R22411 VDD.n3878 VDD.n215 10.2285
R22412 VDD.n3878 VDD.n209 10.2285
R22413 VDD.n3884 VDD.n209 10.2285
R22414 VDD.n3884 VDD.n186 10.2285
R22415 VDD.n3925 VDD.n186 10.2285
R22416 VDD.t126 VDD.n815 9.62685
R22417 VDD.n493 VDD.t130 9.62685
R22418 VDD.n1686 VDD.n1685 9.3005
R22419 VDD.n1687 VDD.n1294 9.3005
R22420 VDD.n1689 VDD.n1688 9.3005
R22421 VDD.n1284 VDD.n1283 9.3005
R22422 VDD.n1702 VDD.n1701 9.3005
R22423 VDD.n1703 VDD.n1282 9.3005
R22424 VDD.n1705 VDD.n1704 9.3005
R22425 VDD.n1272 VDD.n1271 9.3005
R22426 VDD.n1718 VDD.n1717 9.3005
R22427 VDD.n1719 VDD.n1270 9.3005
R22428 VDD.n1721 VDD.n1720 9.3005
R22429 VDD.n1260 VDD.n1259 9.3005
R22430 VDD.n1734 VDD.n1733 9.3005
R22431 VDD.n1735 VDD.n1258 9.3005
R22432 VDD.n1737 VDD.n1736 9.3005
R22433 VDD.n1249 VDD.n1248 9.3005
R22434 VDD.n1750 VDD.n1749 9.3005
R22435 VDD.n1751 VDD.n1247 9.3005
R22436 VDD.n1753 VDD.n1752 9.3005
R22437 VDD.n1236 VDD.n1235 9.3005
R22438 VDD.n1768 VDD.n1767 9.3005
R22439 VDD.n1769 VDD.n1234 9.3005
R22440 VDD.n1802 VDD.n1801 9.3005
R22441 VDD.n1798 VDD.n1770 9.3005
R22442 VDD.n1797 VDD.n1773 9.3005
R22443 VDD.n1777 VDD.n1774 9.3005
R22444 VDD.n1778 VDD.n1775 9.3005
R22445 VDD.n1790 VDD.n1779 9.3005
R22446 VDD.n1789 VDD.n1780 9.3005
R22447 VDD.n1788 VDD.n1781 9.3005
R22448 VDD.n1783 VDD.n1782 9.3005
R22449 VDD.n1800 VDD.n1799 9.3005
R22450 VDD.n1144 VDD.n1138 9.3005
R22451 VDD.n1869 VDD.n1160 9.3005
R22452 VDD.n1868 VDD.n1867 9.3005
R22453 VDD.n1165 VDD.n1164 9.3005
R22454 VDD.n1862 VDD.n1168 9.3005
R22455 VDD.n1861 VDD.n1169 9.3005
R22456 VDD.n1860 VDD.n1170 9.3005
R22457 VDD.n1174 VDD.n1171 9.3005
R22458 VDD.n1855 VDD.n1175 9.3005
R22459 VDD.n1854 VDD.n1176 9.3005
R22460 VDD.n1853 VDD.n1177 9.3005
R22461 VDD.n1184 VDD.n1178 9.3005
R22462 VDD.n1848 VDD.n1847 9.3005
R22463 VDD.n1846 VDD.n1181 9.3005
R22464 VDD.n1845 VDD.n1844 9.3005
R22465 VDD.n1186 VDD.n1185 9.3005
R22466 VDD.n1839 VDD.n1189 9.3005
R22467 VDD.n1838 VDD.n1190 9.3005
R22468 VDD.n1837 VDD.n1191 9.3005
R22469 VDD.n1195 VDD.n1192 9.3005
R22470 VDD.n1832 VDD.n1196 9.3005
R22471 VDD.n1831 VDD.n1197 9.3005
R22472 VDD.n1830 VDD.n1198 9.3005
R22473 VDD.n1871 VDD.n1870 9.3005
R22474 VDD.n1884 VDD.n1139 9.3005
R22475 VDD.n1883 VDD.n1149 9.3005
R22476 VDD.n1153 VDD.n1150 9.3005
R22477 VDD.n1878 VDD.n1154 9.3005
R22478 VDD.n1877 VDD.n1155 9.3005
R22479 VDD.n1876 VDD.n1156 9.3005
R22480 VDD.n1163 VDD.n1157 9.3005
R22481 VDD.n3987 VDD.n3986 9.3005
R22482 VDD.n3990 VDD.n169 9.3005
R22483 VDD.n3991 VDD.n168 9.3005
R22484 VDD.n3994 VDD.n167 9.3005
R22485 VDD.n3995 VDD.n166 9.3005
R22486 VDD.n3998 VDD.n165 9.3005
R22487 VDD.n3999 VDD.n164 9.3005
R22488 VDD.n4002 VDD.n163 9.3005
R22489 VDD.n4003 VDD.n162 9.3005
R22490 VDD.n4006 VDD.n161 9.3005
R22491 VDD.n4007 VDD.n158 9.3005
R22492 VDD.n4010 VDD.n157 9.3005
R22493 VDD.n4011 VDD.n156 9.3005
R22494 VDD.n4014 VDD.n155 9.3005
R22495 VDD.n4015 VDD.n154 9.3005
R22496 VDD.n4018 VDD.n153 9.3005
R22497 VDD.n4019 VDD.n152 9.3005
R22498 VDD.n4022 VDD.n151 9.3005
R22499 VDD.n4023 VDD.n150 9.3005
R22500 VDD.n4026 VDD.n149 9.3005
R22501 VDD.n4030 VDD.n4029 9.3005
R22502 VDD.n4031 VDD.n148 9.3005
R22503 VDD.n4035 VDD.n4032 9.3005
R22504 VDD.n4038 VDD.n147 9.3005
R22505 VDD.n4039 VDD.n146 9.3005
R22506 VDD.n4042 VDD.n145 9.3005
R22507 VDD.n4043 VDD.n144 9.3005
R22508 VDD.n4046 VDD.n143 9.3005
R22509 VDD.n4047 VDD.n142 9.3005
R22510 VDD.n4050 VDD.n141 9.3005
R22511 VDD.n4062 VDD.n135 9.3005
R22512 VDD.n4063 VDD.n134 9.3005
R22513 VDD.n4066 VDD.n133 9.3005
R22514 VDD.n4067 VDD.n132 9.3005
R22515 VDD.n4070 VDD.n131 9.3005
R22516 VDD.n4071 VDD.n130 9.3005
R22517 VDD.n4072 VDD.n129 9.3005
R22518 VDD.n98 VDD.n97 9.3005
R22519 VDD.n4078 VDD.n4077 9.3005
R22520 VDD.n4059 VDD.n136 9.3005
R22521 VDD.n4079 VDD.n96 9.3005
R22522 VDD.n4081 VDD.n4080 9.3005
R22523 VDD.n86 VDD.n85 9.3005
R22524 VDD.n4094 VDD.n4093 9.3005
R22525 VDD.n4095 VDD.n84 9.3005
R22526 VDD.n4097 VDD.n4096 9.3005
R22527 VDD.n74 VDD.n73 9.3005
R22528 VDD.n4109 VDD.n4108 9.3005
R22529 VDD.n4110 VDD.n72 9.3005
R22530 VDD.n4112 VDD.n4111 9.3005
R22531 VDD.n62 VDD.n61 9.3005
R22532 VDD.n4125 VDD.n4124 9.3005
R22533 VDD.n4126 VDD.n60 9.3005
R22534 VDD.n4128 VDD.n4127 9.3005
R22535 VDD.n50 VDD.n49 9.3005
R22536 VDD.n4141 VDD.n4140 9.3005
R22537 VDD.n4142 VDD.n48 9.3005
R22538 VDD.n4144 VDD.n4143 9.3005
R22539 VDD.n38 VDD.n37 9.3005
R22540 VDD.n4157 VDD.n4156 9.3005
R22541 VDD.n4158 VDD.n36 9.3005
R22542 VDD.n4160 VDD.n4159 9.3005
R22543 VDD.n22 VDD.n20 9.3005
R22544 VDD.n4542 VDD.n4541 9.3005
R22545 VDD.n23 VDD.n21 9.3005
R22546 VDD.n4532 VDD.n4174 9.3005
R22547 VDD.n4531 VDD.n4175 9.3005
R22548 VDD.n4530 VDD.n4176 9.3005
R22549 VDD.n4184 VDD.n4177 9.3005
R22550 VDD.n4524 VDD.n4185 9.3005
R22551 VDD.n4523 VDD.n4186 9.3005
R22552 VDD.n4522 VDD.n4187 9.3005
R22553 VDD.n4195 VDD.n4188 9.3005
R22554 VDD.n4516 VDD.n4196 9.3005
R22555 VDD.n4515 VDD.n4197 9.3005
R22556 VDD.n4514 VDD.n4198 9.3005
R22557 VDD.n4206 VDD.n4199 9.3005
R22558 VDD.n4508 VDD.n4207 9.3005
R22559 VDD.n4507 VDD.n4208 9.3005
R22560 VDD.n4506 VDD.n4209 9.3005
R22561 VDD.n4249 VDD.n4210 9.3005
R22562 VDD.n4497 VDD.n4250 9.3005
R22563 VDD.n4496 VDD.n4251 9.3005
R22564 VDD.n4495 VDD.n4252 9.3005
R22565 VDD.n4260 VDD.n4253 9.3005
R22566 VDD.n4489 VDD.n4261 9.3005
R22567 VDD.n4488 VDD.n4487 9.3005
R22568 VDD.n4263 VDD.n4262 9.3005
R22569 VDD.n4267 VDD.n4265 9.3005
R22570 VDD.n4478 VDD.n4268 9.3005
R22571 VDD.n4477 VDD.n4269 9.3005
R22572 VDD.n4476 VDD.n4270 9.3005
R22573 VDD.n4274 VDD.n4271 9.3005
R22574 VDD.n4471 VDD.n4275 9.3005
R22575 VDD.n4470 VDD.n4276 9.3005
R22576 VDD.n4469 VDD.n4468 9.3005
R22577 VDD.n4467 VDD.n4277 9.3005
R22578 VDD.n4466 VDD.n4465 9.3005
R22579 VDD.n4283 VDD.n4282 9.3005
R22580 VDD.n4460 VDD.n4287 9.3005
R22581 VDD.n4459 VDD.n4288 9.3005
R22582 VDD.n4458 VDD.n4289 9.3005
R22583 VDD.n4293 VDD.n4290 9.3005
R22584 VDD.n4453 VDD.n4294 9.3005
R22585 VDD.n4452 VDD.n4295 9.3005
R22586 VDD.n4451 VDD.n4296 9.3005
R22587 VDD.n4303 VDD.n4297 9.3005
R22588 VDD.n4446 VDD.n4445 9.3005
R22589 VDD.n4444 VDD.n4300 9.3005
R22590 VDD.n4443 VDD.n4442 9.3005
R22591 VDD.n4305 VDD.n4304 9.3005
R22592 VDD.n4437 VDD.n4308 9.3005
R22593 VDD.n4436 VDD.n4309 9.3005
R22594 VDD.n4435 VDD.n4310 9.3005
R22595 VDD.n4314 VDD.n4311 9.3005
R22596 VDD.n4430 VDD.n4315 9.3005
R22597 VDD.n4429 VDD.n4316 9.3005
R22598 VDD.n4428 VDD.n4317 9.3005
R22599 VDD.n4324 VDD.n4318 9.3005
R22600 VDD.n4423 VDD.n4422 9.3005
R22601 VDD.n4421 VDD.n4321 9.3005
R22602 VDD.n4420 VDD.n4419 9.3005
R22603 VDD.n4326 VDD.n4325 9.3005
R22604 VDD.n4414 VDD.n4329 9.3005
R22605 VDD.n4413 VDD.n4330 9.3005
R22606 VDD.n4412 VDD.n4331 9.3005
R22607 VDD.n4335 VDD.n4332 9.3005
R22608 VDD.n4407 VDD.n4336 9.3005
R22609 VDD.n4406 VDD.n4337 9.3005
R22610 VDD.n4405 VDD.n4338 9.3005
R22611 VDD.n4345 VDD.n4339 9.3005
R22612 VDD.n4400 VDD.n4346 9.3005
R22613 VDD.n4399 VDD.n4347 9.3005
R22614 VDD.n4398 VDD.n4348 9.3005
R22615 VDD.n4352 VDD.n4349 9.3005
R22616 VDD.n4393 VDD.n4353 9.3005
R22617 VDD.n4392 VDD.n4354 9.3005
R22618 VDD.n4391 VDD.n4355 9.3005
R22619 VDD.n4359 VDD.n4356 9.3005
R22620 VDD.n4386 VDD.n4360 9.3005
R22621 VDD.n4385 VDD.n4361 9.3005
R22622 VDD.n4384 VDD.n4362 9.3005
R22623 VDD.n4368 VDD.n4365 9.3005
R22624 VDD.n4379 VDD.n4378 9.3005
R22625 VDD.n4486 VDD.n4485 9.3005
R22626 VDD.n4086 VDD.n4085 9.3005
R22627 VDD.n4087 VDD.n90 9.3005
R22628 VDD.n4089 VDD.n4088 9.3005
R22629 VDD.n80 VDD.n79 9.3005
R22630 VDD.n4102 VDD.n4101 9.3005
R22631 VDD.n4103 VDD.n78 9.3005
R22632 VDD.n4105 VDD.n4104 9.3005
R22633 VDD.n68 VDD.n67 9.3005
R22634 VDD.n4117 VDD.n4116 9.3005
R22635 VDD.n4118 VDD.n66 9.3005
R22636 VDD.n4120 VDD.n4119 9.3005
R22637 VDD.n56 VDD.n55 9.3005
R22638 VDD.n4133 VDD.n4132 9.3005
R22639 VDD.n4134 VDD.n54 9.3005
R22640 VDD.n4136 VDD.n4135 9.3005
R22641 VDD.n44 VDD.n43 9.3005
R22642 VDD.n4149 VDD.n4148 9.3005
R22643 VDD.n4150 VDD.n42 9.3005
R22644 VDD.n4152 VDD.n4151 9.3005
R22645 VDD.n32 VDD.n31 9.3005
R22646 VDD.n4165 VDD.n4164 9.3005
R22647 VDD.n4166 VDD.n30 9.3005
R22648 VDD.n4538 VDD.n4167 9.3005
R22649 VDD.n4537 VDD.n4168 9.3005
R22650 VDD.n4536 VDD.n4169 9.3005
R22651 VDD.n4223 VDD.n4170 9.3005
R22652 VDD.n4225 VDD.n4224 9.3005
R22653 VDD.n4226 VDD.n4222 9.3005
R22654 VDD.n4228 VDD.n4227 9.3005
R22655 VDD.n4229 VDD.n4221 9.3005
R22656 VDD.n4231 VDD.n4230 9.3005
R22657 VDD.n4232 VDD.n4219 9.3005
R22658 VDD.n4234 VDD.n4233 9.3005
R22659 VDD.n4235 VDD.n4218 9.3005
R22660 VDD.n4237 VDD.n4236 9.3005
R22661 VDD.n4238 VDD.n4216 9.3005
R22662 VDD.n4240 VDD.n4239 9.3005
R22663 VDD.n4241 VDD.n4215 9.3005
R22664 VDD.n4503 VDD.n4242 9.3005
R22665 VDD.n4502 VDD.n4243 9.3005
R22666 VDD.n4501 VDD.n4244 9.3005
R22667 VDD.n4371 VDD.n4245 9.3005
R22668 VDD.n4372 VDD.n4370 9.3005
R22669 VDD.n4374 VDD.n4373 9.3005
R22670 VDD.n4375 VDD.n4369 9.3005
R22671 VDD.n4377 VDD.n4376 9.3005
R22672 VDD.n92 VDD.n91 9.3005
R22673 VDD.n3962 VDD.n3960 9.3005
R22674 VDD.n3966 VDD.n3963 9.3005
R22675 VDD.n3967 VDD.n3959 9.3005
R22676 VDD.n3970 VDD.n3958 9.3005
R22677 VDD.n3971 VDD.n3957 9.3005
R22678 VDD.n3974 VDD.n3956 9.3005
R22679 VDD.n3975 VDD.n3955 9.3005
R22680 VDD.n3978 VDD.n3954 9.3005
R22681 VDD.n3979 VDD.n3953 9.3005
R22682 VDD.n3982 VDD.n171 9.3005
R22683 VDD.n3985 VDD.n3949 9.3005
R22684 VDD.n3985 VDD.n170 9.3005
R22685 VDD.n1823 VDD.n1199 9.3005
R22686 VDD.n1823 VDD.n1206 9.3005
R22687 VDD.n1822 VDD.n1821 9.3005
R22688 VDD.n1820 VDD.n1207 9.3005
R22689 VDD.n1819 VDD.n1818 9.3005
R22690 VDD.n1817 VDD.n1214 9.3005
R22691 VDD.n1816 VDD.n1815 9.3005
R22692 VDD.n1814 VDD.n1215 9.3005
R22693 VDD.n1813 VDD.n1812 9.3005
R22694 VDD.n1811 VDD.n1222 9.3005
R22695 VDD.n1810 VDD.n1809 9.3005
R22696 VDD.n1224 VDD.n1223 9.3005
R22697 VDD.n1365 VDD.n1364 9.3005
R22698 VDD.n1598 VDD.n1597 9.3005
R22699 VDD.n1599 VDD.n1363 9.3005
R22700 VDD.n1601 VDD.n1600 9.3005
R22701 VDD.n1353 VDD.n1352 9.3005
R22702 VDD.n1614 VDD.n1613 9.3005
R22703 VDD.n1615 VDD.n1351 9.3005
R22704 VDD.n1617 VDD.n1616 9.3005
R22705 VDD.n1342 VDD.n1341 9.3005
R22706 VDD.n1630 VDD.n1629 9.3005
R22707 VDD.n1631 VDD.n1340 9.3005
R22708 VDD.n1633 VDD.n1632 9.3005
R22709 VDD.n1330 VDD.n1329 9.3005
R22710 VDD.n1646 VDD.n1645 9.3005
R22711 VDD.n1647 VDD.n1328 9.3005
R22712 VDD.n1649 VDD.n1648 9.3005
R22713 VDD.n1318 VDD.n1317 9.3005
R22714 VDD.n1662 VDD.n1661 9.3005
R22715 VDD.n1663 VDD.n1316 9.3005
R22716 VDD.n1665 VDD.n1664 9.3005
R22717 VDD.n1306 VDD.n1305 9.3005
R22718 VDD.n1678 VDD.n1677 9.3005
R22719 VDD.n1679 VDD.n1304 9.3005
R22720 VDD.n1681 VDD.n1680 9.3005
R22721 VDD.n1290 VDD.n1289 9.3005
R22722 VDD.n1694 VDD.n1693 9.3005
R22723 VDD.n1695 VDD.n1288 9.3005
R22724 VDD.n1697 VDD.n1696 9.3005
R22725 VDD.n1278 VDD.n1277 9.3005
R22726 VDD.n1710 VDD.n1709 9.3005
R22727 VDD.n1711 VDD.n1276 9.3005
R22728 VDD.n1713 VDD.n1712 9.3005
R22729 VDD.n1266 VDD.n1265 9.3005
R22730 VDD.n1726 VDD.n1725 9.3005
R22731 VDD.n1727 VDD.n1264 9.3005
R22732 VDD.n1729 VDD.n1728 9.3005
R22733 VDD.n1254 VDD.n1253 9.3005
R22734 VDD.n1742 VDD.n1741 9.3005
R22735 VDD.n1743 VDD.n1252 9.3005
R22736 VDD.n1745 VDD.n1744 9.3005
R22737 VDD.n1243 VDD.n1242 9.3005
R22738 VDD.n1758 VDD.n1757 9.3005
R22739 VDD.n1759 VDD.n1240 9.3005
R22740 VDD.n1763 VDD.n1762 9.3005
R22741 VDD.n1761 VDD.n1241 9.3005
R22742 VDD.n1760 VDD.n1230 9.3005
R22743 VDD.n1585 VDD.n1584 9.3005
R22744 VDD.n1580 VDD.n1579 9.3005
R22745 VDD.n1578 VDD.n1378 9.3005
R22746 VDD.n1577 VDD.n1576 9.3005
R22747 VDD.n1382 VDD.n1381 9.3005
R22748 VDD.n1569 VDD.n1568 9.3005
R22749 VDD.n1567 VDD.n1384 9.3005
R22750 VDD.n1566 VDD.n1565 9.3005
R22751 VDD.n1386 VDD.n1385 9.3005
R22752 VDD.n1559 VDD.n1558 9.3005
R22753 VDD.n1557 VDD.n1388 9.3005
R22754 VDD.n1556 VDD.n1555 9.3005
R22755 VDD.n1393 VDD.n1389 9.3005
R22756 VDD.n1549 VDD.n1548 9.3005
R22757 VDD.n1547 VDD.n1395 9.3005
R22758 VDD.n1546 VDD.n1545 9.3005
R22759 VDD.n1397 VDD.n1396 9.3005
R22760 VDD.n1539 VDD.n1538 9.3005
R22761 VDD.n1537 VDD.n1399 9.3005
R22762 VDD.n1536 VDD.n1535 9.3005
R22763 VDD.n1401 VDD.n1400 9.3005
R22764 VDD.n1529 VDD.n1528 9.3005
R22765 VDD.n1527 VDD.n1403 9.3005
R22766 VDD.n1526 VDD.n1525 9.3005
R22767 VDD.n1524 VDD.n1404 9.3005
R22768 VDD.n1514 VDD.n1409 9.3005
R22769 VDD.n1515 VDD.n1410 9.3005
R22770 VDD.n1517 VDD.n1516 9.3005
R22771 VDD.n1513 VDD.n1412 9.3005
R22772 VDD.n1512 VDD.n1511 9.3005
R22773 VDD.n1414 VDD.n1413 9.3005
R22774 VDD.n1505 VDD.n1504 9.3005
R22775 VDD.n1503 VDD.n1416 9.3005
R22776 VDD.n1502 VDD.n1501 9.3005
R22777 VDD.n1418 VDD.n1417 9.3005
R22778 VDD.n1495 VDD.n1420 9.3005
R22779 VDD.n1494 VDD.n1493 9.3005
R22780 VDD.n1492 VDD.n1423 9.3005
R22781 VDD.n1491 VDD.n1490 9.3005
R22782 VDD.n1425 VDD.n1424 9.3005
R22783 VDD.n1481 VDD.n1428 9.3005
R22784 VDD.n1483 VDD.n1482 9.3005
R22785 VDD.n1480 VDD.n1430 9.3005
R22786 VDD.n1479 VDD.n1478 9.3005
R22787 VDD.n1432 VDD.n1431 9.3005
R22788 VDD.n1472 VDD.n1471 9.3005
R22789 VDD.n1470 VDD.n1434 9.3005
R22790 VDD.n1467 VDD.n1435 9.3005
R22791 VDD.n1457 VDD.n1440 9.3005
R22792 VDD.n1458 VDD.n1441 9.3005
R22793 VDD.n1460 VDD.n1459 9.3005
R22794 VDD.n1456 VDD.n1443 9.3005
R22795 VDD.n1455 VDD.n1454 9.3005
R22796 VDD.n1445 VDD.n1444 9.3005
R22797 VDD.n1448 VDD.n1447 9.3005
R22798 VDD.n1446 VDD.n1370 9.3005
R22799 VDD.n1469 VDD.n1468 9.3005
R22800 VDD.n1581 VDD.n1374 9.3005
R22801 VDD.n1583 VDD.n1582 9.3005
R22802 VDD.n1591 VDD.n1369 9.3005
R22803 VDD.n1593 VDD.n1592 9.3005
R22804 VDD.n1359 VDD.n1358 9.3005
R22805 VDD.n1606 VDD.n1605 9.3005
R22806 VDD.n1607 VDD.n1357 9.3005
R22807 VDD.n1609 VDD.n1608 9.3005
R22808 VDD.n1348 VDD.n1347 9.3005
R22809 VDD.n1622 VDD.n1621 9.3005
R22810 VDD.n1623 VDD.n1346 9.3005
R22811 VDD.n1625 VDD.n1624 9.3005
R22812 VDD.n1336 VDD.n1335 9.3005
R22813 VDD.n1638 VDD.n1637 9.3005
R22814 VDD.n1639 VDD.n1334 9.3005
R22815 VDD.n1641 VDD.n1640 9.3005
R22816 VDD.n1324 VDD.n1323 9.3005
R22817 VDD.n1654 VDD.n1653 9.3005
R22818 VDD.n1655 VDD.n1322 9.3005
R22819 VDD.n1657 VDD.n1656 9.3005
R22820 VDD.n1312 VDD.n1311 9.3005
R22821 VDD.n1670 VDD.n1669 9.3005
R22822 VDD.n1671 VDD.n1310 9.3005
R22823 VDD.n1673 VDD.n1672 9.3005
R22824 VDD.n1590 VDD.n1589 9.3005
R22825 VDD.n1301 VDD.n1300 9.3005
R22826 VDD.n2728 VDD.t97 9.0252
R22827 VDD.n3522 VDD.t95 9.0252
R22828 VDD.n2422 VDD.t22 8.72438
R22829 VDD.n2147 VDD.t29 8.72438
R22830 VDD.n3369 VDD.t50 8.72438
R22831 VDD.n3828 VDD.t18 8.72438
R22832 VDD.n2147 VDD.t124 8.42355
R22833 VDD.n3369 VDD.t128 8.42355
R22834 VDD.n15 VDD.n14 8.357
R22835 VDD.n4543 VDD.n4542 8.07375
R22836 VDD.n1300 VDD.n1299 8.07375
R22837 VDD.n1468 VDD.n1434 7.95202
R22838 VDD.n1892 VDD.n1144 7.95202
R22839 VDD.n4469 VDD.n4277 7.95202
R22840 VDD.n4059 VDD.n4058 7.95202
R22841 VDD.n2524 VDD.t99 7.82191
R22842 VDD.n3726 VDD.t115 7.82191
R22843 VDD.n1026 VDD.t109 7.22026
R22844 VDD.t122 VDD.n282 7.22026
R22845 VDD.n1525 VDD.n1524 7.17626
R22846 VDD.n1848 VDD.n1178 7.17626
R22847 VDD.n4423 VDD.n4318 7.17626
R22848 VDD.n4010 VDD.n4007 7.17626
R22849 VDD.n2410 VDD.t117 6.61861
R22850 VDD.n3840 VDD.t101 6.61861
R22851 VDD.t121 VDD.n994 6.31779
R22852 VDD.n2716 VDD.t108 6.31779
R22853 VDD.n3534 VDD.t114 6.31779
R22854 VDD.n314 VDD.t120 6.31779
R22855 VDD.n2548 VDD.t119 5.71614
R22856 VDD.n835 VDD.t111 5.71614
R22857 VDD.t107 VDD.n473 5.71614
R22858 VDD.n3702 VDD.t103 5.71614
R22859 VDD.n2830 VDD.n674 5.46391
R22860 VDD.n1928 VDD.n1927 5.46391
R22861 VDD.n3397 VDD.n3396 5.46391
R22862 VDD.n205 VDD.n203 5.46391
R22863 VDD.n181 VDD.n179 5.46391
R22864 VDD.n3145 VDD.n3119 5.46391
R22865 VDD.n2874 VDD.n2873 5.46391
R22866 VDD.n2357 VDD.n2356 5.46391
R22867 VDD.n1896 VDD.n1895 5.30782
R22868 VDD.n1918 VDD.n1895 5.30782
R22869 VDD.n3908 VDD.n3907 5.30782
R22870 VDD.n3907 VDD.n3905 5.30782
R22871 VDD.n3943 VDD.n172 5.30782
R22872 VDD.n3943 VDD.n3942 5.30782
R22873 VDD.n2369 VDD.n1110 5.30782
R22874 VDD.n2365 VDD.n1110 5.30782
R22875 VDD.n2833 VDD.n674 5.15172
R22876 VDD.n1927 VDD.n1926 5.15172
R22877 VDD.n3398 VDD.n3397 5.15172
R22878 VDD.n3898 VDD.n203 5.15172
R22879 VDD.n3935 VDD.n179 5.15172
R22880 VDD.n3142 VDD.n3119 5.15172
R22881 VDD.n2875 VDD.n2874 5.15172
R22882 VDD.n2358 VDD.n2357 5.15172
R22883 VDD.n2602 VDD.t104 5.1145
R22884 VDD.t104 VDD.n880 5.1145
R22885 VDD.n427 VDD.t94 5.1145
R22886 VDD.n3648 VDD.t94 5.1145
R22887 VDD.n1555 VDD.n1392 4.84898
R22888 VDD.n1825 VDD.n1204 4.84898
R22889 VDD.n4400 VDD.n4344 4.84898
R22890 VDD.n3949 VDD.n3946 4.84898
R22891 VDD.n1825 VDD.n1824 4.74817
R22892 VDD.n1893 VDD.n1892 4.74817
R22893 VDD.n1147 VDD.n1140 4.74817
R22894 VDD.n1893 VDD.n1141 4.74817
R22895 VDD.n1885 VDD.n1140 4.74817
R22896 VDD.n4058 VDD.n139 4.74817
R22897 VDD.n4051 VDD.n140 4.74817
R22898 VDD.n4054 VDD.n140 4.74817
R22899 VDD.n4055 VDD.n139 4.74817
R22900 VDD.n3984 VDD.n3983 4.74817
R22901 VDD.n3984 VDD.n3950 4.74817
R22902 VDD.n1824 VDD.n1205 4.74817
R22903 VDD.n948 VDD.t119 4.51285
R22904 VDD.n2662 VDD.t111 4.51285
R22905 VDD.n3588 VDD.t107 4.51285
R22906 VDD.t103 VDD.n360 4.51285
R22907 VDD.n4543 VDD.n19 4.17173
R22908 VDD.n1299 VDD.n1298 4.17173
R22909 VDD.n2488 VDD.t121 3.9112
R22910 VDD.t108 VDD.n766 3.9112
R22911 VDD.n541 VDD.t114 3.9112
R22912 VDD.n3762 VDD.t120 3.9112
R22913 VDD.t117 VDD.n1071 3.61038
R22914 VDD.n236 VDD.t101 3.61038
R22915 VDD.n2470 VDD.t109 3.00873
R22916 VDD.n3780 VDD.t122 3.00873
R22917 VDD.n1299 VDD.n15 2.56827
R22918 VDD VDD.n4543 2.56043
R22919 VDD.t99 VDD.n958 2.40709
R22920 VDD.n350 VDD.t115 2.40709
R22921 VDD.n4 VDD.n2 2.31084
R22922 VDD.n11 VDD.n9 2.31084
R22923 VDD.n1894 VDD.n1893 2.27742
R22924 VDD.n1894 VDD.n1140 2.27742
R22925 VDD.n3906 VDD.n140 2.27742
R22926 VDD.n3906 VDD.n139 2.27742
R22927 VDD.n3985 VDD.n3984 2.27742
R22928 VDD.n1824 VDD.n1823 2.27742
R22929 VDD.n6 VDD.n4 1.86257
R22930 VDD.n13 VDD.n11 1.86257
R22931 VDD.n2782 VDD.t124 1.80544
R22932 VDD.n3468 VDD.t128 1.80544
R22933 VDD.n1393 VDD.n1392 1.74595
R22934 VDD.n1204 VDD.n1199 1.74595
R22935 VDD.n4344 VDD.n4339 1.74595
R22936 VDD.n3946 VDD.n170 1.74595
R22937 VDD.n1074 VDD.t22 1.50462
R22938 VDD.n2788 VDD.t29 1.50462
R22939 VDD.n3462 VDD.t50 1.50462
R22940 VDD.t18 VDD.n233 1.50462
R22941 VDD.n14 VDD.n6 1.44016
R22942 VDD.n14 VDD.n13 1.44016
R22943 VDD.n769 VDD.t97 1.20379
R22944 VDD.t95 VDD.n538 1.20379
R22945 VDD.n19 VDD.n18 0.842454
R22946 VDD.n18 VDD.n17 0.842454
R22947 VDD.n17 VDD.n16 0.842454
R22948 VDD.n1298 VDD.n1297 0.842454
R22949 VDD.n1297 VDD.n1296 0.842454
R22950 VDD.n1296 VDD.n1295 0.842454
R22951 VDD.n2668 VDD.t126 0.602147
R22952 VDD.n3582 VDD.t130 0.602147
R22953 VDD.n1801 VDD.n1800 0.474585
R22954 VDD.n4079 VDD.n4078 0.474585
R22955 VDD.n4487 VDD.n4486 0.474585
R22956 VDD.n4378 VDD.n4377 0.474585
R22957 VDD.n3962 VDD.n91 0.474585
R22958 VDD.n1760 VDD.n1223 0.474585
R22959 VDD.n1584 VDD.n1583 0.474585
R22960 VDD.n1590 VDD.n1370 0.474585
R22961 VDD.n1687 VDD.n1686 0.152939
R22962 VDD.n1688 VDD.n1687 0.152939
R22963 VDD.n1688 VDD.n1283 0.152939
R22964 VDD.n1702 VDD.n1283 0.152939
R22965 VDD.n1703 VDD.n1702 0.152939
R22966 VDD.n1704 VDD.n1703 0.152939
R22967 VDD.n1704 VDD.n1271 0.152939
R22968 VDD.n1718 VDD.n1271 0.152939
R22969 VDD.n1719 VDD.n1718 0.152939
R22970 VDD.n1720 VDD.n1719 0.152939
R22971 VDD.n1720 VDD.n1259 0.152939
R22972 VDD.n1734 VDD.n1259 0.152939
R22973 VDD.n1735 VDD.n1734 0.152939
R22974 VDD.n1736 VDD.n1735 0.152939
R22975 VDD.n1736 VDD.n1248 0.152939
R22976 VDD.n1750 VDD.n1248 0.152939
R22977 VDD.n1751 VDD.n1750 0.152939
R22978 VDD.n1752 VDD.n1751 0.152939
R22979 VDD.n1752 VDD.n1235 0.152939
R22980 VDD.n1768 VDD.n1235 0.152939
R22981 VDD.n1769 VDD.n1768 0.152939
R22982 VDD.n1801 VDD.n1769 0.152939
R22983 VDD.n1800 VDD.n1770 0.152939
R22984 VDD.n1773 VDD.n1770 0.152939
R22985 VDD.n1777 VDD.n1773 0.152939
R22986 VDD.n1778 VDD.n1777 0.152939
R22987 VDD.n1779 VDD.n1778 0.152939
R22988 VDD.n1780 VDD.n1779 0.152939
R22989 VDD.n1781 VDD.n1780 0.152939
R22990 VDD.n1782 VDD.n1781 0.152939
R22991 VDD.n1782 VDD.n1138 0.152939
R22992 VDD.n1149 VDD.n1139 0.152939
R22993 VDD.n1153 VDD.n1149 0.152939
R22994 VDD.n1154 VDD.n1153 0.152939
R22995 VDD.n1155 VDD.n1154 0.152939
R22996 VDD.n1156 VDD.n1155 0.152939
R22997 VDD.n1163 VDD.n1156 0.152939
R22998 VDD.n1870 VDD.n1163 0.152939
R22999 VDD.n1870 VDD.n1869 0.152939
R23000 VDD.n1869 VDD.n1868 0.152939
R23001 VDD.n1868 VDD.n1164 0.152939
R23002 VDD.n1168 VDD.n1164 0.152939
R23003 VDD.n1169 VDD.n1168 0.152939
R23004 VDD.n1170 VDD.n1169 0.152939
R23005 VDD.n1174 VDD.n1170 0.152939
R23006 VDD.n1175 VDD.n1174 0.152939
R23007 VDD.n1176 VDD.n1175 0.152939
R23008 VDD.n1177 VDD.n1176 0.152939
R23009 VDD.n1184 VDD.n1177 0.152939
R23010 VDD.n1847 VDD.n1184 0.152939
R23011 VDD.n1847 VDD.n1846 0.152939
R23012 VDD.n1846 VDD.n1845 0.152939
R23013 VDD.n1845 VDD.n1185 0.152939
R23014 VDD.n1189 VDD.n1185 0.152939
R23015 VDD.n1190 VDD.n1189 0.152939
R23016 VDD.n1191 VDD.n1190 0.152939
R23017 VDD.n1195 VDD.n1191 0.152939
R23018 VDD.n1196 VDD.n1195 0.152939
R23019 VDD.n1197 VDD.n1196 0.152939
R23020 VDD.n1198 VDD.n1197 0.152939
R23021 VDD.n142 VDD.n141 0.152939
R23022 VDD.n143 VDD.n142 0.152939
R23023 VDD.n144 VDD.n143 0.152939
R23024 VDD.n145 VDD.n144 0.152939
R23025 VDD.n146 VDD.n145 0.152939
R23026 VDD.n147 VDD.n146 0.152939
R23027 VDD.n4032 VDD.n147 0.152939
R23028 VDD.n4032 VDD.n4031 0.152939
R23029 VDD.n4031 VDD.n4030 0.152939
R23030 VDD.n4030 VDD.n149 0.152939
R23031 VDD.n150 VDD.n149 0.152939
R23032 VDD.n151 VDD.n150 0.152939
R23033 VDD.n152 VDD.n151 0.152939
R23034 VDD.n153 VDD.n152 0.152939
R23035 VDD.n154 VDD.n153 0.152939
R23036 VDD.n155 VDD.n154 0.152939
R23037 VDD.n156 VDD.n155 0.152939
R23038 VDD.n157 VDD.n156 0.152939
R23039 VDD.n158 VDD.n157 0.152939
R23040 VDD.n161 VDD.n158 0.152939
R23041 VDD.n162 VDD.n161 0.152939
R23042 VDD.n163 VDD.n162 0.152939
R23043 VDD.n164 VDD.n163 0.152939
R23044 VDD.n165 VDD.n164 0.152939
R23045 VDD.n166 VDD.n165 0.152939
R23046 VDD.n167 VDD.n166 0.152939
R23047 VDD.n168 VDD.n167 0.152939
R23048 VDD.n169 VDD.n168 0.152939
R23049 VDD.n3986 VDD.n169 0.152939
R23050 VDD.n4078 VDD.n97 0.152939
R23051 VDD.n129 VDD.n97 0.152939
R23052 VDD.n130 VDD.n129 0.152939
R23053 VDD.n131 VDD.n130 0.152939
R23054 VDD.n132 VDD.n131 0.152939
R23055 VDD.n133 VDD.n132 0.152939
R23056 VDD.n134 VDD.n133 0.152939
R23057 VDD.n135 VDD.n134 0.152939
R23058 VDD.n136 VDD.n135 0.152939
R23059 VDD.n4080 VDD.n4079 0.152939
R23060 VDD.n4080 VDD.n85 0.152939
R23061 VDD.n4094 VDD.n85 0.152939
R23062 VDD.n4095 VDD.n4094 0.152939
R23063 VDD.n4096 VDD.n4095 0.152939
R23064 VDD.n4096 VDD.n73 0.152939
R23065 VDD.n4109 VDD.n73 0.152939
R23066 VDD.n4110 VDD.n4109 0.152939
R23067 VDD.n4111 VDD.n4110 0.152939
R23068 VDD.n4111 VDD.n61 0.152939
R23069 VDD.n4125 VDD.n61 0.152939
R23070 VDD.n4126 VDD.n4125 0.152939
R23071 VDD.n4127 VDD.n4126 0.152939
R23072 VDD.n4127 VDD.n49 0.152939
R23073 VDD.n4141 VDD.n49 0.152939
R23074 VDD.n4142 VDD.n4141 0.152939
R23075 VDD.n4143 VDD.n4142 0.152939
R23076 VDD.n4143 VDD.n37 0.152939
R23077 VDD.n4157 VDD.n37 0.152939
R23078 VDD.n4158 VDD.n4157 0.152939
R23079 VDD.n4159 VDD.n4158 0.152939
R23080 VDD.n4159 VDD.n20 0.152939
R23081 VDD.n4174 VDD.n21 0.152939
R23082 VDD.n4175 VDD.n4174 0.152939
R23083 VDD.n4176 VDD.n4175 0.152939
R23084 VDD.n4184 VDD.n4176 0.152939
R23085 VDD.n4185 VDD.n4184 0.152939
R23086 VDD.n4186 VDD.n4185 0.152939
R23087 VDD.n4187 VDD.n4186 0.152939
R23088 VDD.n4195 VDD.n4187 0.152939
R23089 VDD.n4196 VDD.n4195 0.152939
R23090 VDD.n4197 VDD.n4196 0.152939
R23091 VDD.n4198 VDD.n4197 0.152939
R23092 VDD.n4206 VDD.n4198 0.152939
R23093 VDD.n4207 VDD.n4206 0.152939
R23094 VDD.n4208 VDD.n4207 0.152939
R23095 VDD.n4209 VDD.n4208 0.152939
R23096 VDD.n4249 VDD.n4209 0.152939
R23097 VDD.n4250 VDD.n4249 0.152939
R23098 VDD.n4251 VDD.n4250 0.152939
R23099 VDD.n4252 VDD.n4251 0.152939
R23100 VDD.n4260 VDD.n4252 0.152939
R23101 VDD.n4261 VDD.n4260 0.152939
R23102 VDD.n4487 VDD.n4261 0.152939
R23103 VDD.n4486 VDD.n4262 0.152939
R23104 VDD.n4267 VDD.n4262 0.152939
R23105 VDD.n4268 VDD.n4267 0.152939
R23106 VDD.n4269 VDD.n4268 0.152939
R23107 VDD.n4270 VDD.n4269 0.152939
R23108 VDD.n4274 VDD.n4270 0.152939
R23109 VDD.n4275 VDD.n4274 0.152939
R23110 VDD.n4276 VDD.n4275 0.152939
R23111 VDD.n4468 VDD.n4276 0.152939
R23112 VDD.n4468 VDD.n4467 0.152939
R23113 VDD.n4467 VDD.n4466 0.152939
R23114 VDD.n4466 VDD.n4282 0.152939
R23115 VDD.n4287 VDD.n4282 0.152939
R23116 VDD.n4288 VDD.n4287 0.152939
R23117 VDD.n4289 VDD.n4288 0.152939
R23118 VDD.n4293 VDD.n4289 0.152939
R23119 VDD.n4294 VDD.n4293 0.152939
R23120 VDD.n4295 VDD.n4294 0.152939
R23121 VDD.n4296 VDD.n4295 0.152939
R23122 VDD.n4303 VDD.n4296 0.152939
R23123 VDD.n4445 VDD.n4303 0.152939
R23124 VDD.n4445 VDD.n4444 0.152939
R23125 VDD.n4444 VDD.n4443 0.152939
R23126 VDD.n4443 VDD.n4304 0.152939
R23127 VDD.n4308 VDD.n4304 0.152939
R23128 VDD.n4309 VDD.n4308 0.152939
R23129 VDD.n4310 VDD.n4309 0.152939
R23130 VDD.n4314 VDD.n4310 0.152939
R23131 VDD.n4315 VDD.n4314 0.152939
R23132 VDD.n4316 VDD.n4315 0.152939
R23133 VDD.n4317 VDD.n4316 0.152939
R23134 VDD.n4324 VDD.n4317 0.152939
R23135 VDD.n4422 VDD.n4324 0.152939
R23136 VDD.n4422 VDD.n4421 0.152939
R23137 VDD.n4421 VDD.n4420 0.152939
R23138 VDD.n4420 VDD.n4325 0.152939
R23139 VDD.n4329 VDD.n4325 0.152939
R23140 VDD.n4330 VDD.n4329 0.152939
R23141 VDD.n4331 VDD.n4330 0.152939
R23142 VDD.n4335 VDD.n4331 0.152939
R23143 VDD.n4336 VDD.n4335 0.152939
R23144 VDD.n4337 VDD.n4336 0.152939
R23145 VDD.n4338 VDD.n4337 0.152939
R23146 VDD.n4345 VDD.n4338 0.152939
R23147 VDD.n4346 VDD.n4345 0.152939
R23148 VDD.n4347 VDD.n4346 0.152939
R23149 VDD.n4348 VDD.n4347 0.152939
R23150 VDD.n4352 VDD.n4348 0.152939
R23151 VDD.n4353 VDD.n4352 0.152939
R23152 VDD.n4354 VDD.n4353 0.152939
R23153 VDD.n4355 VDD.n4354 0.152939
R23154 VDD.n4359 VDD.n4355 0.152939
R23155 VDD.n4360 VDD.n4359 0.152939
R23156 VDD.n4361 VDD.n4360 0.152939
R23157 VDD.n4362 VDD.n4361 0.152939
R23158 VDD.n4368 VDD.n4362 0.152939
R23159 VDD.n4378 VDD.n4368 0.152939
R23160 VDD.n4086 VDD.n91 0.152939
R23161 VDD.n4087 VDD.n4086 0.152939
R23162 VDD.n4088 VDD.n4087 0.152939
R23163 VDD.n4088 VDD.n79 0.152939
R23164 VDD.n4102 VDD.n79 0.152939
R23165 VDD.n4103 VDD.n4102 0.152939
R23166 VDD.n4104 VDD.n4103 0.152939
R23167 VDD.n4104 VDD.n67 0.152939
R23168 VDD.n4117 VDD.n67 0.152939
R23169 VDD.n4118 VDD.n4117 0.152939
R23170 VDD.n4119 VDD.n4118 0.152939
R23171 VDD.n4119 VDD.n55 0.152939
R23172 VDD.n4133 VDD.n55 0.152939
R23173 VDD.n4134 VDD.n4133 0.152939
R23174 VDD.n4135 VDD.n4134 0.152939
R23175 VDD.n4135 VDD.n43 0.152939
R23176 VDD.n4149 VDD.n43 0.152939
R23177 VDD.n4150 VDD.n4149 0.152939
R23178 VDD.n4151 VDD.n4150 0.152939
R23179 VDD.n4151 VDD.n31 0.152939
R23180 VDD.n4165 VDD.n31 0.152939
R23181 VDD.n4166 VDD.n4165 0.152939
R23182 VDD.n4167 VDD.n4166 0.152939
R23183 VDD.n4168 VDD.n4167 0.152939
R23184 VDD.n4169 VDD.n4168 0.152939
R23185 VDD.n4223 VDD.n4169 0.152939
R23186 VDD.n4224 VDD.n4223 0.152939
R23187 VDD.n4224 VDD.n4222 0.152939
R23188 VDD.n4228 VDD.n4222 0.152939
R23189 VDD.n4229 VDD.n4228 0.152939
R23190 VDD.n4230 VDD.n4229 0.152939
R23191 VDD.n4230 VDD.n4219 0.152939
R23192 VDD.n4234 VDD.n4219 0.152939
R23193 VDD.n4235 VDD.n4234 0.152939
R23194 VDD.n4236 VDD.n4235 0.152939
R23195 VDD.n4236 VDD.n4216 0.152939
R23196 VDD.n4240 VDD.n4216 0.152939
R23197 VDD.n4241 VDD.n4240 0.152939
R23198 VDD.n4242 VDD.n4241 0.152939
R23199 VDD.n4243 VDD.n4242 0.152939
R23200 VDD.n4244 VDD.n4243 0.152939
R23201 VDD.n4371 VDD.n4244 0.152939
R23202 VDD.n4372 VDD.n4371 0.152939
R23203 VDD.n4373 VDD.n4372 0.152939
R23204 VDD.n4373 VDD.n4369 0.152939
R23205 VDD.n4377 VDD.n4369 0.152939
R23206 VDD.n3953 VDD.n171 0.152939
R23207 VDD.n3954 VDD.n3953 0.152939
R23208 VDD.n3955 VDD.n3954 0.152939
R23209 VDD.n3956 VDD.n3955 0.152939
R23210 VDD.n3957 VDD.n3956 0.152939
R23211 VDD.n3958 VDD.n3957 0.152939
R23212 VDD.n3959 VDD.n3958 0.152939
R23213 VDD.n3963 VDD.n3959 0.152939
R23214 VDD.n3963 VDD.n3962 0.152939
R23215 VDD.n1822 VDD.n1207 0.152939
R23216 VDD.n1818 VDD.n1207 0.152939
R23217 VDD.n1818 VDD.n1817 0.152939
R23218 VDD.n1817 VDD.n1816 0.152939
R23219 VDD.n1816 VDD.n1215 0.152939
R23220 VDD.n1812 VDD.n1215 0.152939
R23221 VDD.n1812 VDD.n1811 0.152939
R23222 VDD.n1811 VDD.n1810 0.152939
R23223 VDD.n1810 VDD.n1223 0.152939
R23224 VDD.n1584 VDD.n1364 0.152939
R23225 VDD.n1598 VDD.n1364 0.152939
R23226 VDD.n1599 VDD.n1598 0.152939
R23227 VDD.n1600 VDD.n1599 0.152939
R23228 VDD.n1600 VDD.n1352 0.152939
R23229 VDD.n1614 VDD.n1352 0.152939
R23230 VDD.n1615 VDD.n1614 0.152939
R23231 VDD.n1616 VDD.n1615 0.152939
R23232 VDD.n1616 VDD.n1341 0.152939
R23233 VDD.n1630 VDD.n1341 0.152939
R23234 VDD.n1631 VDD.n1630 0.152939
R23235 VDD.n1632 VDD.n1631 0.152939
R23236 VDD.n1632 VDD.n1329 0.152939
R23237 VDD.n1646 VDD.n1329 0.152939
R23238 VDD.n1647 VDD.n1646 0.152939
R23239 VDD.n1648 VDD.n1647 0.152939
R23240 VDD.n1648 VDD.n1317 0.152939
R23241 VDD.n1662 VDD.n1317 0.152939
R23242 VDD.n1663 VDD.n1662 0.152939
R23243 VDD.n1664 VDD.n1663 0.152939
R23244 VDD.n1664 VDD.n1305 0.152939
R23245 VDD.n1678 VDD.n1305 0.152939
R23246 VDD.n1679 VDD.n1678 0.152939
R23247 VDD.n1680 VDD.n1679 0.152939
R23248 VDD.n1680 VDD.n1289 0.152939
R23249 VDD.n1694 VDD.n1289 0.152939
R23250 VDD.n1695 VDD.n1694 0.152939
R23251 VDD.n1696 VDD.n1695 0.152939
R23252 VDD.n1696 VDD.n1277 0.152939
R23253 VDD.n1710 VDD.n1277 0.152939
R23254 VDD.n1711 VDD.n1710 0.152939
R23255 VDD.n1712 VDD.n1711 0.152939
R23256 VDD.n1712 VDD.n1265 0.152939
R23257 VDD.n1726 VDD.n1265 0.152939
R23258 VDD.n1727 VDD.n1726 0.152939
R23259 VDD.n1728 VDD.n1727 0.152939
R23260 VDD.n1728 VDD.n1253 0.152939
R23261 VDD.n1742 VDD.n1253 0.152939
R23262 VDD.n1743 VDD.n1742 0.152939
R23263 VDD.n1744 VDD.n1743 0.152939
R23264 VDD.n1744 VDD.n1242 0.152939
R23265 VDD.n1758 VDD.n1242 0.152939
R23266 VDD.n1759 VDD.n1758 0.152939
R23267 VDD.n1762 VDD.n1759 0.152939
R23268 VDD.n1762 VDD.n1761 0.152939
R23269 VDD.n1761 VDD.n1760 0.152939
R23270 VDD.n1447 VDD.n1370 0.152939
R23271 VDD.n1447 VDD.n1444 0.152939
R23272 VDD.n1455 VDD.n1444 0.152939
R23273 VDD.n1456 VDD.n1455 0.152939
R23274 VDD.n1459 VDD.n1456 0.152939
R23275 VDD.n1459 VDD.n1458 0.152939
R23276 VDD.n1458 VDD.n1457 0.152939
R23277 VDD.n1457 VDD.n1435 0.152939
R23278 VDD.n1469 VDD.n1435 0.152939
R23279 VDD.n1470 VDD.n1469 0.152939
R23280 VDD.n1471 VDD.n1470 0.152939
R23281 VDD.n1471 VDD.n1431 0.152939
R23282 VDD.n1479 VDD.n1431 0.152939
R23283 VDD.n1480 VDD.n1479 0.152939
R23284 VDD.n1482 VDD.n1480 0.152939
R23285 VDD.n1482 VDD.n1481 0.152939
R23286 VDD.n1481 VDD.n1424 0.152939
R23287 VDD.n1491 VDD.n1424 0.152939
R23288 VDD.n1492 VDD.n1491 0.152939
R23289 VDD.n1493 VDD.n1492 0.152939
R23290 VDD.n1493 VDD.n1420 0.152939
R23291 VDD.n1420 VDD.n1417 0.152939
R23292 VDD.n1502 VDD.n1417 0.152939
R23293 VDD.n1503 VDD.n1502 0.152939
R23294 VDD.n1504 VDD.n1503 0.152939
R23295 VDD.n1504 VDD.n1413 0.152939
R23296 VDD.n1512 VDD.n1413 0.152939
R23297 VDD.n1513 VDD.n1512 0.152939
R23298 VDD.n1516 VDD.n1513 0.152939
R23299 VDD.n1516 VDD.n1515 0.152939
R23300 VDD.n1515 VDD.n1514 0.152939
R23301 VDD.n1514 VDD.n1404 0.152939
R23302 VDD.n1526 VDD.n1404 0.152939
R23303 VDD.n1527 VDD.n1526 0.152939
R23304 VDD.n1528 VDD.n1527 0.152939
R23305 VDD.n1528 VDD.n1400 0.152939
R23306 VDD.n1536 VDD.n1400 0.152939
R23307 VDD.n1537 VDD.n1536 0.152939
R23308 VDD.n1538 VDD.n1537 0.152939
R23309 VDD.n1538 VDD.n1396 0.152939
R23310 VDD.n1546 VDD.n1396 0.152939
R23311 VDD.n1547 VDD.n1546 0.152939
R23312 VDD.n1548 VDD.n1547 0.152939
R23313 VDD.n1548 VDD.n1389 0.152939
R23314 VDD.n1556 VDD.n1389 0.152939
R23315 VDD.n1557 VDD.n1556 0.152939
R23316 VDD.n1558 VDD.n1557 0.152939
R23317 VDD.n1558 VDD.n1385 0.152939
R23318 VDD.n1566 VDD.n1385 0.152939
R23319 VDD.n1567 VDD.n1566 0.152939
R23320 VDD.n1568 VDD.n1567 0.152939
R23321 VDD.n1568 VDD.n1381 0.152939
R23322 VDD.n1577 VDD.n1381 0.152939
R23323 VDD.n1578 VDD.n1577 0.152939
R23324 VDD.n1579 VDD.n1578 0.152939
R23325 VDD.n1579 VDD.n1374 0.152939
R23326 VDD.n1583 VDD.n1374 0.152939
R23327 VDD.n1591 VDD.n1590 0.152939
R23328 VDD.n1592 VDD.n1591 0.152939
R23329 VDD.n1592 VDD.n1358 0.152939
R23330 VDD.n1606 VDD.n1358 0.152939
R23331 VDD.n1607 VDD.n1606 0.152939
R23332 VDD.n1608 VDD.n1607 0.152939
R23333 VDD.n1608 VDD.n1347 0.152939
R23334 VDD.n1622 VDD.n1347 0.152939
R23335 VDD.n1623 VDD.n1622 0.152939
R23336 VDD.n1624 VDD.n1623 0.152939
R23337 VDD.n1624 VDD.n1335 0.152939
R23338 VDD.n1638 VDD.n1335 0.152939
R23339 VDD.n1639 VDD.n1638 0.152939
R23340 VDD.n1640 VDD.n1639 0.152939
R23341 VDD.n1640 VDD.n1323 0.152939
R23342 VDD.n1654 VDD.n1323 0.152939
R23343 VDD.n1655 VDD.n1654 0.152939
R23344 VDD.n1656 VDD.n1655 0.152939
R23345 VDD.n1656 VDD.n1311 0.152939
R23346 VDD.n1670 VDD.n1311 0.152939
R23347 VDD.n1671 VDD.n1670 0.152939
R23348 VDD.n1672 VDD.n1671 0.152939
R23349 VDD.n1686 VDD.n1300 0.145814
R23350 VDD.n4542 VDD.n20 0.145814
R23351 VDD.n4542 VDD.n21 0.145814
R23352 VDD.n1672 VDD.n1300 0.145814
R23353 VDD.n1894 VDD.n1139 0.110256
R23354 VDD.n1823 VDD.n1198 0.110256
R23355 VDD.n3906 VDD.n141 0.110256
R23356 VDD.n3986 VDD.n3985 0.110256
R23357 VDD.n1894 VDD.n1138 0.0431829
R23358 VDD.n3906 VDD.n136 0.0431829
R23359 VDD.n3985 VDD.n171 0.0431829
R23360 VDD.n1823 VDD.n1822 0.0431829
R23361 VDD VDD.n15 0.00833333
R23362 a_n8732_9422.n0 a_n8732_9422.t7 156.754
R23363 a_n8732_9422.n2 a_n8732_9422.t13 156.754
R23364 a_n8732_9422.n1 a_n8732_9422.t11 156.754
R23365 a_n8732_9422.n0 a_n8732_9422.t1 154.892
R23366 a_n8732_9422.n0 a_n8732_9422.t5 154.892
R23367 a_n8732_9422.n3 a_n8732_9422.t4 154.892
R23368 a_n8732_9422.n0 a_n8732_9422.n10 129.496
R23369 a_n8732_9422.n1 a_n8732_9422.n4 129.496
R23370 a_n8732_9422.n1 a_n8732_9422.n5 129.496
R23371 a_n8732_9422.n2 a_n8732_9422.n7 129.496
R23372 a_n8732_9422.n2 a_n8732_9422.n8 129.496
R23373 a_n8732_9422.n11 a_n8732_9422.n0 129.496
R23374 a_n8732_9422.n9 a_n8732_9422.n2 29.8996
R23375 a_n8732_9422.n10 a_n8732_9422.t6 25.395
R23376 a_n8732_9422.n10 a_n8732_9422.t3 25.395
R23377 a_n8732_9422.n4 a_n8732_9422.t12 25.395
R23378 a_n8732_9422.n4 a_n8732_9422.t15 25.395
R23379 a_n8732_9422.n5 a_n8732_9422.t10 25.395
R23380 a_n8732_9422.n5 a_n8732_9422.t18 25.395
R23381 a_n8732_9422.n7 a_n8732_9422.t9 25.395
R23382 a_n8732_9422.n7 a_n8732_9422.t14 25.395
R23383 a_n8732_9422.n8 a_n8732_9422.t16 25.395
R23384 a_n8732_9422.n8 a_n8732_9422.t17 25.395
R23385 a_n8732_9422.t8 a_n8732_9422.n11 25.395
R23386 a_n8732_9422.n11 a_n8732_9422.t2 25.395
R23387 a_n8732_9422.n6 a_n8732_9422.t0 12.3901
R23388 a_n8732_9422.n6 a_n8732_9422.n1 10.8216
R23389 a_n8732_9422.n0 a_n8732_9422.n3 6.03498
R23390 a_n8732_9422.n3 a_n8732_9422.n9 5.8403
R23391 a_n8732_9422.n9 a_n8732_9422.n6 3.45315
R23392 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t1 98.5576
R23393 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t5 97.0364
R23394 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t7 97.0364
R23395 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t3 97.0364
R23396 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t0 51.0487
R23397 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t9 50.2711
R23398 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t4 46.484
R23399 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t6 46.484
R23400 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t2 46.484
R23401 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.t10 45.7068
R23402 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t11 45.7068
R23403 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t8 45.7068
R23404 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 7.0929
R23405 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 4.84777
R23406 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n3 4.57865
R23407 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 4.56629
R23408 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n4 4.56629
R23409 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 4.56605
R23410 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 3.27913
R23411 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 1.52182
R23412 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 1.52182
R23413 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n0 0.996727
R23414 DIFFPAIR_BIAS DIFFPAIR_BIAS.n10 0.942375
R23415 a_n3337_n4072.n0 a_n3337_n4072.t0 166.048
R23416 a_n3337_n4072.n0 a_n3337_n4072.t2 165.242
R23417 a_n3337_n4072.n0 a_n3337_n4072.t1 164.528
R23418 a_n3337_n4072.t3 a_n3337_n4072.n0 164.528
R23419 a_n3337_n4072.n1 a_n3337_n4072.t7 47.8704
R23420 a_n3337_n4072.n2 a_n3337_n4072.t4 47.8702
R23421 a_n3337_n4072.n2 a_n3337_n4072.t5 47.8702
R23422 a_n3337_n4072.n1 a_n3337_n4072.t6 47.8702
R23423 a_n3337_n4072.n0 a_n3337_n4072.n1 6.4942
R23424 a_n3337_n4072.n0 a_n3337_n4072.n2 3.80629
R23425 VP.n6 VP.t6 243.255
R23426 VP.n3 VP.n1 224.169
R23427 VP.n5 VP.n4 223.454
R23428 VP.n3 VP.n2 223.454
R23429 VP.n0 VP.t7 153.304
R23430 VP.n0 VP.t8 137.145
R23431 VP.n4 VP.t0 19.8005
R23432 VP.n4 VP.t3 19.8005
R23433 VP.n2 VP.t5 19.8005
R23434 VP.n2 VP.t1 19.8005
R23435 VP.n1 VP.t4 19.8005
R23436 VP.n1 VP.t2 19.8005
R23437 VP VP.n7 15.2825
R23438 VP.n7 VP.n6 4.80222
R23439 VP.n7 VP.n0 0.972091
R23440 VP.n5 VP.n3 0.716017
R23441 VP.n6 VP.n5 0.716017
R23442 a_n17232_8522.n5 a_n17232_8522.t2 176.341
R23443 a_n17232_8522.n3 a_n17232_8522.t9 174.48
R23444 a_n17232_8522.n2 a_n17232_8522.n0 150.946
R23445 a_n17232_8522.n7 a_n17232_8522.n6 149.084
R23446 a_n17232_8522.n5 a_n17232_8522.n4 149.084
R23447 a_n17232_8522.n2 a_n17232_8522.n1 149.084
R23448 a_n17232_8522.t11 a_n17232_8522.n19 98.7471
R23449 a_n17232_8522.n19 a_n17232_8522.t10 67.6717
R23450 a_n17232_8522.n13 a_n17232_8522.t19 49.4355
R23451 a_n17232_8522.n9 a_n17232_8522.t14 49.4355
R23452 a_n17232_8522.n12 a_n17232_8522.t16 47.2537
R23453 a_n17232_8522.n11 a_n17232_8522.t21 47.2537
R23454 a_n17232_8522.n10 a_n17232_8522.t17 47.2537
R23455 a_n17232_8522.n9 a_n17232_8522.t15 47.2537
R23456 a_n17232_8522.n16 a_n17232_8522.t13 47.252
R23457 a_n17232_8522.n15 a_n17232_8522.t18 47.252
R23458 a_n17232_8522.n14 a_n17232_8522.t12 47.252
R23459 a_n17232_8522.n13 a_n17232_8522.t20 47.252
R23460 a_n17232_8522.n8 a_n17232_8522.n3 31.6281
R23461 a_n17232_8522.n8 a_n17232_8522.n7 25.4057
R23462 a_n17232_8522.n6 a_n17232_8522.t4 25.395
R23463 a_n17232_8522.n6 a_n17232_8522.t6 25.395
R23464 a_n17232_8522.n4 a_n17232_8522.t1 25.395
R23465 a_n17232_8522.n4 a_n17232_8522.t0 25.395
R23466 a_n17232_8522.n0 a_n17232_8522.t3 25.395
R23467 a_n17232_8522.n0 a_n17232_8522.t8 25.395
R23468 a_n17232_8522.n1 a_n17232_8522.t5 25.395
R23469 a_n17232_8522.n1 a_n17232_8522.t7 25.395
R23470 a_n17232_8522.n19 a_n17232_8522.n18 12.4268
R23471 a_n17232_8522.n18 a_n17232_8522.n8 11.6469
R23472 a_n17232_8522.n17 a_n17232_8522.n12 7.11248
R23473 a_n17232_8522.n17 a_n17232_8522.n16 6.97492
R23474 a_n17232_8522.n18 a_n17232_8522.n17 3.4105
R23475 a_n17232_8522.n14 a_n17232_8522.n13 2.18232
R23476 a_n17232_8522.n15 a_n17232_8522.n14 2.18232
R23477 a_n17232_8522.n16 a_n17232_8522.n15 2.18232
R23478 a_n17232_8522.n10 a_n17232_8522.n9 2.18232
R23479 a_n17232_8522.n11 a_n17232_8522.n10 2.18232
R23480 a_n17232_8522.n12 a_n17232_8522.n11 2.18232
R23481 a_n17232_8522.n7 a_n17232_8522.n5 1.86257
R23482 a_n17232_8522.n3 a_n17232_8522.n2 1.86257
C0 VDD VOUT 38.1964f
C1 VOUT CS_BIAS 22.718401f
C2 a_n13358_11043# VDD 1.91085f
C3 VDD VN 0.243578f
C4 VOUT VP 5.34203f
C5 VOUT VN 0.992027f
C6 CS_BIAS VP 0.326881f
C7 CS_BIAS VN 0.246305f
C8 VP VN 11.676001f
C9 a_11906_11043# VDD 1.91081f
C10 DIFFPAIR_BIAS GND 60.296528f
C11 VN GND 29.812737f
C12 VP GND 28.29834f
C13 CS_BIAS GND 95.08453f
C14 VOUT GND 74.30639f
C15 VDD GND 0.767362p
C16 a_11906_11043# GND 0.744974f
C17 a_n13358_11043# GND 0.744829f
C18 a_n17232_8522.t3 GND 0.054205f
C19 a_n17232_8522.t8 GND 0.054205f
C20 a_n17232_8522.n0 GND 0.259827f
C21 a_n17232_8522.t5 GND 0.054205f
C22 a_n17232_8522.t7 GND 0.054205f
C23 a_n17232_8522.n1 GND 0.237774f
C24 a_n17232_8522.n2 GND 3.53714f
C25 a_n17232_8522.t9 GND 0.32053f
C26 a_n17232_8522.n3 GND 5.70516f
C27 a_n17232_8522.t2 GND 0.332247f
C28 a_n17232_8522.t1 GND 0.054205f
C29 a_n17232_8522.t0 GND 0.054205f
C30 a_n17232_8522.n4 GND 0.237774f
C31 a_n17232_8522.n5 GND 2.86938f
C32 a_n17232_8522.t4 GND 0.054205f
C33 a_n17232_8522.t6 GND 0.054205f
C34 a_n17232_8522.n6 GND 0.237774f
C35 a_n17232_8522.n7 GND 5.90408f
C36 a_n17232_8522.n8 GND 14.028799f
C37 a_n17232_8522.t14 GND 1.97493f
C38 a_n17232_8522.t15 GND 1.92775f
C39 a_n17232_8522.n9 GND 2.20567f
C40 a_n17232_8522.t17 GND 1.92775f
C41 a_n17232_8522.n10 GND 1.18391f
C42 a_n17232_8522.t21 GND 1.92775f
C43 a_n17232_8522.n11 GND 1.18391f
C44 a_n17232_8522.t16 GND 1.92775f
C45 a_n17232_8522.n12 GND 4.25358f
C46 a_n17232_8522.t19 GND 1.97493f
C47 a_n17232_8522.t20 GND 1.9277f
C48 a_n17232_8522.n13 GND 2.20572f
C49 a_n17232_8522.t12 GND 1.9277f
C50 a_n17232_8522.n14 GND 1.18396f
C51 a_n17232_8522.t18 GND 1.9277f
C52 a_n17232_8522.n15 GND 1.18396f
C53 a_n17232_8522.t13 GND 1.9277f
C54 a_n17232_8522.n16 GND 4.00631f
C55 a_n17232_8522.n17 GND 25.3281f
C56 a_n17232_8522.n18 GND 3.41886f
C57 a_n17232_8522.t10 GND 1.33622f
C58 a_n17232_8522.n19 GND 4.24366f
C59 a_n17232_8522.t11 GND 1.99025f
C60 VP.t8 GND 0.998586f
C61 VP.t7 GND 1.10422f
C62 VP.n0 GND 1.96366f
C63 VP.t4 GND 0.005486f
C64 VP.t2 GND 0.005486f
C65 VP.n1 GND 0.01804f
C66 VP.t5 GND 0.005486f
C67 VP.t1 GND 0.005486f
C68 VP.n2 GND 0.017793f
C69 VP.n3 GND 0.151857f
C70 VP.t0 GND 0.005486f
C71 VP.t3 GND 0.005486f
C72 VP.n4 GND 0.017793f
C73 VP.n5 GND 0.074654f
C74 VP.t6 GND 0.030536f
C75 VP.n6 GND 0.082867f
C76 VP.n7 GND 2.70293f
C77 a_n3337_n4072.n0 GND 5.50326f
C78 a_n3337_n4072.n1 GND 1.36774f
C79 a_n3337_n4072.n2 GND 1.19949f
C80 a_n3337_n4072.t0 GND 0.467519f
C81 a_n3337_n4072.t1 GND 0.460965f
C82 a_n3337_n4072.t6 GND 0.49325f
C83 a_n3337_n4072.t7 GND 0.493252f
C84 a_n3337_n4072.t5 GND 0.49325f
C85 a_n3337_n4072.t4 GND 0.49325f
C86 a_n3337_n4072.t2 GND 0.46706f
C87 a_n3337_n4072.t3 GND 0.460965f
C88 DIFFPAIR_BIAS.t8 GND 0.123363f
C89 DIFFPAIR_BIAS.t9 GND 0.131866f
C90 DIFFPAIR_BIAS.n0 GND 0.154206f
C91 DIFFPAIR_BIAS.t10 GND 0.123363f
C92 DIFFPAIR_BIAS.t11 GND 0.123363f
C93 DIFFPAIR_BIAS.t1 GND 0.03384f
C94 DIFFPAIR_BIAS.t5 GND 0.032286f
C95 DIFFPAIR_BIAS.n1 GND 0.20625f
C96 DIFFPAIR_BIAS.t7 GND 0.032286f
C97 DIFFPAIR_BIAS.n2 GND 0.1071f
C98 DIFFPAIR_BIAS.t3 GND 0.032286f
C99 DIFFPAIR_BIAS.n3 GND 0.115886f
C100 DIFFPAIR_BIAS.t2 GND 0.12106f
C101 DIFFPAIR_BIAS.t6 GND 0.12106f
C102 DIFFPAIR_BIAS.t4 GND 0.12106f
C103 DIFFPAIR_BIAS.t0 GND 0.127843f
C104 DIFFPAIR_BIAS.n4 GND 0.154091f
C105 DIFFPAIR_BIAS.n5 GND 0.085007f
C106 DIFFPAIR_BIAS.n6 GND 0.086891f
C107 DIFFPAIR_BIAS.n7 GND 0.083941f
C108 DIFFPAIR_BIAS.n8 GND 0.079859f
C109 DIFFPAIR_BIAS.n9 GND 0.081719f
C110 DIFFPAIR_BIAS.n10 GND 0.041244f
C111 a_n8732_9422.n0 GND 7.22253f
C112 a_n8732_9422.n1 GND 6.63884f
C113 a_n8732_9422.n2 GND 9.05216f
C114 a_n8732_9422.n3 GND 2.06304f
C115 a_n8732_9422.t0 GND 48.452602f
C116 a_n8732_9422.t11 GND 0.297649f
C117 a_n8732_9422.t12 GND 0.056093f
C118 a_n8732_9422.t15 GND 0.056093f
C119 a_n8732_9422.n4 GND 0.19671f
C120 a_n8732_9422.t10 GND 0.056093f
C121 a_n8732_9422.t18 GND 0.056093f
C122 a_n8732_9422.n5 GND 0.19671f
C123 a_n8732_9422.n6 GND 4.76386f
C124 a_n8732_9422.t13 GND 0.29765f
C125 a_n8732_9422.t9 GND 0.056093f
C126 a_n8732_9422.t14 GND 0.056093f
C127 a_n8732_9422.n7 GND 0.19671f
C128 a_n8732_9422.t16 GND 0.056093f
C129 a_n8732_9422.t17 GND 0.056093f
C130 a_n8732_9422.n8 GND 0.19671f
C131 a_n8732_9422.n9 GND 5.80721f
C132 a_n8732_9422.t4 GND 0.284501f
C133 a_n8732_9422.t6 GND 0.056093f
C134 a_n8732_9422.t3 GND 0.056093f
C135 a_n8732_9422.n10 GND 0.19671f
C136 a_n8732_9422.t5 GND 0.284501f
C137 a_n8732_9422.t1 GND 0.284501f
C138 a_n8732_9422.t7 GND 0.29765f
C139 a_n8732_9422.t2 GND 0.056093f
C140 a_n8732_9422.n11 GND 0.19671f
C141 a_n8732_9422.t8 GND 0.056093f
C142 VDD.t113 GND 0.012667f
C143 VDD.t118 GND 0.012667f
C144 VDD.n0 GND 0.06072f
C145 VDD.t110 GND 0.012667f
C146 VDD.t100 GND 0.012667f
C147 VDD.n1 GND 0.055566f
C148 VDD.n2 GND 0.867308f
C149 VDD.t93 GND 0.012667f
C150 VDD.t127 GND 0.012667f
C151 VDD.n3 GND 0.055566f
C152 VDD.n4 GND 0.45469f
C153 VDD.t98 GND 0.012667f
C154 VDD.t125 GND 0.012667f
C155 VDD.n5 GND 0.055566f
C156 VDD.n6 GND 0.375636f
C157 VDD.t102 GND 0.012667f
C158 VDD.t106 GND 0.012667f
C159 VDD.n7 GND 0.06072f
C160 VDD.t116 GND 0.012667f
C161 VDD.t123 GND 0.012667f
C162 VDD.n8 GND 0.055566f
C163 VDD.n9 GND 0.867308f
C164 VDD.t131 GND 0.012667f
C165 VDD.t133 GND 0.012667f
C166 VDD.n10 GND 0.055566f
C167 VDD.n11 GND 0.45469f
C168 VDD.t129 GND 0.012667f
C169 VDD.t96 GND 0.012667f
C170 VDD.n12 GND 0.055566f
C171 VDD.n13 GND 0.375636f
C172 VDD.n14 GND 0.285011f
C173 VDD.n15 GND 2.69436f
C174 VDD.t145 GND 0.070193f
C175 VDD.t140 GND 0.068332f
C176 VDD.n16 GND 0.778374f
C177 VDD.t146 GND 0.068332f
C178 VDD.n17 GND 0.425535f
C179 VDD.t138 GND 0.068332f
C180 VDD.n18 GND 0.425535f
C181 VDD.t139 GND 0.068332f
C182 VDD.n19 GND 0.507397f
C183 VDD.n20 GND 0.006127f
C184 VDD.n21 GND 0.006127f
C185 VDD.n22 GND 0.004948f
C186 VDD.n23 GND 0.004948f
C187 VDD.n24 GND 0.006148f
C188 VDD.n25 GND 0.006148f
C189 VDD.n26 GND 0.473529f
C190 VDD.n27 GND 0.473529f
C191 VDD.n28 GND 0.006148f
C192 VDD.n29 GND 0.006148f
C193 VDD.n30 GND 0.004948f
C194 VDD.n31 GND 0.006148f
C195 VDD.n32 GND 0.004948f
C196 VDD.n33 GND 0.006148f
C197 VDD.n34 GND 0.473529f
C198 VDD.n35 GND 0.006148f
C199 VDD.n36 GND 0.004948f
C200 VDD.n37 GND 0.006148f
C201 VDD.n38 GND 0.004948f
C202 VDD.n39 GND 0.006148f
C203 VDD.n40 GND 0.473529f
C204 VDD.n41 GND 0.006148f
C205 VDD.n42 GND 0.004948f
C206 VDD.n43 GND 0.006148f
C207 VDD.n44 GND 0.004948f
C208 VDD.n45 GND 0.006148f
C209 VDD.n46 GND 0.473529f
C210 VDD.n47 GND 0.006148f
C211 VDD.n48 GND 0.004948f
C212 VDD.n49 GND 0.006148f
C213 VDD.n50 GND 0.004948f
C214 VDD.n51 GND 0.006148f
C215 VDD.n52 GND 0.473529f
C216 VDD.n53 GND 0.006148f
C217 VDD.n54 GND 0.004948f
C218 VDD.n55 GND 0.006148f
C219 VDD.n56 GND 0.004948f
C220 VDD.n57 GND 0.006148f
C221 VDD.n58 GND 0.473529f
C222 VDD.n59 GND 0.006148f
C223 VDD.n60 GND 0.004948f
C224 VDD.n61 GND 0.006148f
C225 VDD.n62 GND 0.004948f
C226 VDD.n63 GND 0.006148f
C227 VDD.n64 GND 0.473529f
C228 VDD.n65 GND 0.006148f
C229 VDD.n66 GND 0.004948f
C230 VDD.n67 GND 0.006148f
C231 VDD.n68 GND 0.004948f
C232 VDD.n69 GND 0.006148f
C233 VDD.n70 GND 0.473529f
C234 VDD.n71 GND 0.006148f
C235 VDD.n72 GND 0.004948f
C236 VDD.n73 GND 0.006148f
C237 VDD.n74 GND 0.004948f
C238 VDD.n75 GND 0.006148f
C239 VDD.n76 GND 0.473529f
C240 VDD.n77 GND 0.006148f
C241 VDD.n78 GND 0.004948f
C242 VDD.n79 GND 0.006148f
C243 VDD.n80 GND 0.004948f
C244 VDD.n81 GND 0.006148f
C245 VDD.n82 GND 0.473529f
C246 VDD.n83 GND 0.006148f
C247 VDD.n84 GND 0.004948f
C248 VDD.n85 GND 0.006148f
C249 VDD.n86 GND 0.004948f
C250 VDD.n87 GND 0.006148f
C251 VDD.n88 GND 0.473529f
C252 VDD.n89 GND 0.006148f
C253 VDD.n90 GND 0.004948f
C254 VDD.n91 GND 0.013671f
C255 VDD.n92 GND 0.004107f
C256 VDD.n93 GND 0.013671f
C257 VDD.n94 GND 0.670043f
C258 VDD.n95 GND 0.013671f
C259 VDD.n96 GND 0.004107f
C260 VDD.n97 GND 0.006148f
C261 VDD.n98 GND 0.004948f
C262 VDD.n99 GND 0.006148f
C263 VDD.t134 GND 7.35153f
C264 VDD.n127 GND 0.014117f
C265 VDD.n128 GND 0.006148f
C266 VDD.n129 GND 0.006148f
C267 VDD.n130 GND 0.006148f
C268 VDD.n131 GND 0.006148f
C269 VDD.n132 GND 0.006148f
C270 VDD.n133 GND 0.006148f
C271 VDD.n134 GND 0.006148f
C272 VDD.n135 GND 0.006148f
C273 VDD.n136 GND 0.003935f
C274 VDD.t48 GND 0.085164f
C275 VDD.t46 GND 0.430073f
C276 VDD.n137 GND 0.075426f
C277 VDD.t47 GND 0.053191f
C278 VDD.n138 GND 0.077435f
C279 VDD.n141 GND 0.005287f
C280 VDD.n142 GND 0.006148f
C281 VDD.n143 GND 0.006148f
C282 VDD.n144 GND 0.006148f
C283 VDD.n145 GND 0.006148f
C284 VDD.n146 GND 0.006148f
C285 VDD.n147 GND 0.006148f
C286 VDD.n148 GND 0.004181f
C287 VDD.n149 GND 0.006148f
C288 VDD.n150 GND 0.006148f
C289 VDD.n151 GND 0.006148f
C290 VDD.n152 GND 0.006148f
C291 VDD.n153 GND 0.006148f
C292 VDD.n154 GND 0.006148f
C293 VDD.n155 GND 0.006148f
C294 VDD.n156 GND 0.006148f
C295 VDD.n157 GND 0.006148f
C296 VDD.n158 GND 0.006148f
C297 VDD.t27 GND 0.085164f
C298 VDD.t25 GND 0.430073f
C299 VDD.n159 GND 0.075426f
C300 VDD.t26 GND 0.053191f
C301 VDD.n160 GND 0.077435f
C302 VDD.n161 GND 0.006148f
C303 VDD.n162 GND 0.006148f
C304 VDD.n163 GND 0.006148f
C305 VDD.n164 GND 0.006148f
C306 VDD.n165 GND 0.006148f
C307 VDD.n166 GND 0.006148f
C308 VDD.n167 GND 0.006148f
C309 VDD.n168 GND 0.006148f
C310 VDD.n169 GND 0.006148f
C311 VDD.n170 GND 0.002697f
C312 VDD.n171 GND 0.003935f
C313 VDD.n172 GND 0.003135f
C314 VDD.n173 GND 0.00418f
C315 VDD.t105 GND 5.13068f
C316 VDD.n175 GND 1.67629f
C317 VDD.n176 GND 0.00418f
C318 VDD.t19 GND 0.089111f
C319 VDD.t17 GND 0.44554f
C320 VDD.n177 GND 0.076053f
C321 VDD.t20 GND 0.056759f
C322 VDD.n178 GND 0.078134f
C323 VDD.n179 GND 0.005158f
C324 VDD.n181 GND 0.003166f
C325 VDD.n182 GND 0.00418f
C326 VDD.n183 GND 0.009354f
C327 VDD.n185 GND 0.00418f
C328 VDD.n186 GND 0.322f
C329 VDD.n187 GND 0.008807f
C330 VDD.n188 GND 0.008807f
C331 VDD.n189 GND 0.00418f
C332 VDD.n190 GND 0.009514f
C333 VDD.n191 GND 0.00418f
C334 VDD.n192 GND 0.00418f
C335 VDD.n194 GND 0.00418f
C336 VDD.n195 GND 0.00418f
C337 VDD.n197 GND 0.00418f
C338 VDD.n198 GND 0.00418f
C339 VDD.n200 GND 0.00418f
C340 VDD.t69 GND 0.089111f
C341 VDD.t68 GND 0.44554f
C342 VDD.n201 GND 0.076053f
C343 VDD.t70 GND 0.056759f
C344 VDD.n202 GND 0.078134f
C345 VDD.n203 GND 0.005158f
C346 VDD.n205 GND 0.003166f
C347 VDD.n206 GND 0.00418f
C348 VDD.n207 GND 0.00418f
C349 VDD.n208 GND 0.00418f
C350 VDD.n209 GND 0.322f
C351 VDD.n210 GND 0.00418f
C352 VDD.n211 GND 0.00418f
C353 VDD.n212 GND 0.00418f
C354 VDD.n213 GND 0.00418f
C355 VDD.n214 GND 0.00418f
C356 VDD.n215 GND 0.322f
C357 VDD.n216 GND 0.00418f
C358 VDD.n217 GND 0.00418f
C359 VDD.n218 GND 0.00418f
C360 VDD.n219 GND 0.00418f
C361 VDD.n220 GND 0.00418f
C362 VDD.n221 GND 0.00418f
C363 VDD.n222 GND 0.322f
C364 VDD.n223 GND 0.00418f
C365 VDD.n224 GND 0.00418f
C366 VDD.n225 GND 0.00418f
C367 VDD.n226 GND 0.00418f
C368 VDD.n227 GND 0.00418f
C369 VDD.t101 GND 0.161f
C370 VDD.n228 GND 0.00418f
C371 VDD.n229 GND 0.00418f
C372 VDD.n230 GND 0.00418f
C373 VDD.n231 GND 0.00418f
C374 VDD.n232 GND 0.00418f
C375 VDD.n233 GND 0.184676f
C376 VDD.n234 GND 0.00418f
C377 VDD.n235 GND 0.00418f
C378 VDD.n236 GND 0.217823f
C379 VDD.n237 GND 0.00418f
C380 VDD.n238 GND 0.00418f
C381 VDD.n239 GND 0.00418f
C382 VDD.n240 GND 0.322f
C383 VDD.n241 GND 0.00418f
C384 VDD.n242 GND 0.00418f
C385 VDD.t18 GND 0.161f
C386 VDD.n243 GND 0.00418f
C387 VDD.n244 GND 0.00418f
C388 VDD.n245 GND 0.00418f
C389 VDD.n246 GND 0.322f
C390 VDD.n247 GND 0.00418f
C391 VDD.n248 GND 0.00418f
C392 VDD.n249 GND 0.00418f
C393 VDD.n250 GND 0.00418f
C394 VDD.n251 GND 0.00418f
C395 VDD.n252 GND 0.322f
C396 VDD.n253 GND 0.00418f
C397 VDD.n254 GND 0.00418f
C398 VDD.n255 GND 0.00418f
C399 VDD.n256 GND 0.00418f
C400 VDD.n257 GND 0.00418f
C401 VDD.n258 GND 0.322f
C402 VDD.n259 GND 0.00418f
C403 VDD.n260 GND 0.00418f
C404 VDD.n261 GND 0.00418f
C405 VDD.n262 GND 0.00418f
C406 VDD.n263 GND 0.00418f
C407 VDD.n264 GND 0.322f
C408 VDD.n265 GND 0.00418f
C409 VDD.n266 GND 0.00418f
C410 VDD.n267 GND 0.00418f
C411 VDD.n268 GND 0.00418f
C412 VDD.n269 GND 0.00418f
C413 VDD.n270 GND 0.322f
C414 VDD.n271 GND 0.00418f
C415 VDD.n272 GND 0.00418f
C416 VDD.n273 GND 0.00418f
C417 VDD.n274 GND 0.00418f
C418 VDD.n275 GND 0.00418f
C419 VDD.n276 GND 0.322f
C420 VDD.n277 GND 0.00418f
C421 VDD.n278 GND 0.00418f
C422 VDD.n279 GND 0.00418f
C423 VDD.n280 GND 0.00418f
C424 VDD.n281 GND 0.00418f
C425 VDD.n282 GND 0.274647f
C426 VDD.n283 GND 0.00418f
C427 VDD.n284 GND 0.00418f
C428 VDD.n285 GND 0.00418f
C429 VDD.n286 GND 0.00418f
C430 VDD.n287 GND 0.00418f
C431 VDD.n288 GND 0.322f
C432 VDD.n289 GND 0.00418f
C433 VDD.n290 GND 0.00418f
C434 VDD.t122 GND 0.161f
C435 VDD.n291 GND 0.00418f
C436 VDD.n292 GND 0.00418f
C437 VDD.n293 GND 0.00418f
C438 VDD.n294 GND 0.322f
C439 VDD.n295 GND 0.00418f
C440 VDD.n296 GND 0.00418f
C441 VDD.n297 GND 0.00418f
C442 VDD.n298 GND 0.00418f
C443 VDD.n299 GND 0.00418f
C444 VDD.n300 GND 0.322f
C445 VDD.n301 GND 0.00418f
C446 VDD.n302 GND 0.00418f
C447 VDD.n303 GND 0.00418f
C448 VDD.n304 GND 0.00418f
C449 VDD.n305 GND 0.00418f
C450 VDD.t120 GND 0.161f
C451 VDD.n306 GND 0.00418f
C452 VDD.n307 GND 0.00418f
C453 VDD.n308 GND 0.00418f
C454 VDD.n309 GND 0.00418f
C455 VDD.n310 GND 0.00418f
C456 VDD.n311 GND 0.322f
C457 VDD.n312 GND 0.00418f
C458 VDD.n313 GND 0.00418f
C459 VDD.n314 GND 0.260441f
C460 VDD.n315 GND 0.00418f
C461 VDD.n316 GND 0.00418f
C462 VDD.n317 GND 0.00418f
C463 VDD.n318 GND 0.322f
C464 VDD.n319 GND 0.00418f
C465 VDD.n320 GND 0.00418f
C466 VDD.n321 GND 0.00418f
C467 VDD.n322 GND 0.00418f
C468 VDD.n323 GND 0.00418f
C469 VDD.n324 GND 0.322f
C470 VDD.n325 GND 0.00418f
C471 VDD.n326 GND 0.00418f
C472 VDD.n327 GND 0.00418f
C473 VDD.n328 GND 0.00418f
C474 VDD.n329 GND 0.00418f
C475 VDD.n330 GND 0.322f
C476 VDD.n331 GND 0.00418f
C477 VDD.n332 GND 0.00418f
C478 VDD.n333 GND 0.00418f
C479 VDD.n334 GND 0.00418f
C480 VDD.n335 GND 0.00418f
C481 VDD.n336 GND 0.322f
C482 VDD.n337 GND 0.00418f
C483 VDD.n338 GND 0.00418f
C484 VDD.n339 GND 0.00418f
C485 VDD.n340 GND 0.00418f
C486 VDD.n341 GND 0.00418f
C487 VDD.t115 GND 0.161f
C488 VDD.n342 GND 0.00418f
C489 VDD.n343 GND 0.00418f
C490 VDD.n344 GND 0.00418f
C491 VDD.n345 GND 0.00418f
C492 VDD.n346 GND 0.00418f
C493 VDD.n347 GND 0.322f
C494 VDD.n348 GND 0.00418f
C495 VDD.n349 GND 0.00418f
C496 VDD.n350 GND 0.198882f
C497 VDD.n351 GND 0.00418f
C498 VDD.n352 GND 0.00418f
C499 VDD.n353 GND 0.00418f
C500 VDD.n354 GND 0.322f
C501 VDD.n355 GND 0.00418f
C502 VDD.n356 GND 0.00418f
C503 VDD.n357 GND 0.00418f
C504 VDD.n358 GND 0.00418f
C505 VDD.n359 GND 0.00418f
C506 VDD.n360 GND 0.232029f
C507 VDD.n361 GND 0.00418f
C508 VDD.n362 GND 0.00418f
C509 VDD.n363 GND 0.00418f
C510 VDD.n364 GND 0.00418f
C511 VDD.n365 GND 0.00418f
C512 VDD.n366 GND 0.322f
C513 VDD.n367 GND 0.00418f
C514 VDD.n368 GND 0.00418f
C515 VDD.t103 GND 0.161f
C516 VDD.n369 GND 0.00418f
C517 VDD.n370 GND 0.00418f
C518 VDD.n371 GND 0.00418f
C519 VDD.n372 GND 0.322f
C520 VDD.n373 GND 0.00418f
C521 VDD.n374 GND 0.00418f
C522 VDD.n375 GND 0.00418f
C523 VDD.n376 GND 0.00418f
C524 VDD.n377 GND 0.00418f
C525 VDD.n378 GND 0.322f
C526 VDD.n379 GND 0.00418f
C527 VDD.n380 GND 0.00418f
C528 VDD.n381 GND 0.00418f
C529 VDD.n382 GND 0.00418f
C530 VDD.n383 GND 0.00418f
C531 VDD.n384 GND 0.322f
C532 VDD.n385 GND 0.00418f
C533 VDD.n386 GND 0.00418f
C534 VDD.n387 GND 0.00418f
C535 VDD.n388 GND 0.00418f
C536 VDD.n389 GND 0.00418f
C537 VDD.n390 GND 0.322f
C538 VDD.n391 GND 0.00418f
C539 VDD.n392 GND 0.00418f
C540 VDD.n393 GND 0.00418f
C541 VDD.n394 GND 0.00418f
C542 VDD.n395 GND 0.00418f
C543 VDD.n396 GND 0.322f
C544 VDD.n397 GND 0.00418f
C545 VDD.n398 GND 0.00418f
C546 VDD.n399 GND 0.00418f
C547 VDD.n400 GND 0.00418f
C548 VDD.n401 GND 0.00418f
C549 VDD.n402 GND 0.322f
C550 VDD.n403 GND 0.00418f
C551 VDD.n404 GND 0.00418f
C552 VDD.n405 GND 0.00418f
C553 VDD.n406 GND 0.00418f
C554 VDD.n407 GND 0.00418f
C555 VDD.n408 GND 0.322f
C556 VDD.n409 GND 0.00418f
C557 VDD.n410 GND 0.00418f
C558 VDD.n411 GND 0.00418f
C559 VDD.n412 GND 0.00418f
C560 VDD.n413 GND 0.00418f
C561 VDD.n414 GND 0.322f
C562 VDD.n415 GND 0.00418f
C563 VDD.n416 GND 0.00418f
C564 VDD.n417 GND 0.00418f
C565 VDD.n418 GND 0.00418f
C566 VDD.n419 GND 0.00418f
C567 VDD.t94 GND 0.161f
C568 VDD.n420 GND 0.00418f
C569 VDD.n421 GND 0.00418f
C570 VDD.n422 GND 0.00418f
C571 VDD.n423 GND 0.00418f
C572 VDD.n424 GND 0.00418f
C573 VDD.t132 GND 0.322f
C574 VDD.n425 GND 0.00418f
C575 VDD.n426 GND 0.00418f
C576 VDD.n427 GND 0.2415f
C577 VDD.n428 GND 0.00418f
C578 VDD.n429 GND 0.00418f
C579 VDD.n430 GND 0.00418f
C580 VDD.n431 GND 0.322f
C581 VDD.n432 GND 0.00418f
C582 VDD.n433 GND 0.00418f
C583 VDD.n434 GND 0.00418f
C584 VDD.n435 GND 0.00418f
C585 VDD.n436 GND 0.00418f
C586 VDD.n437 GND 0.322f
C587 VDD.n438 GND 0.00418f
C588 VDD.n439 GND 0.00418f
C589 VDD.n440 GND 0.00418f
C590 VDD.n441 GND 0.00418f
C591 VDD.n442 GND 0.00418f
C592 VDD.n443 GND 0.322f
C593 VDD.n444 GND 0.00418f
C594 VDD.n445 GND 0.00418f
C595 VDD.n446 GND 0.00418f
C596 VDD.n447 GND 0.00418f
C597 VDD.n448 GND 0.00418f
C598 VDD.n449 GND 0.322f
C599 VDD.n450 GND 0.00418f
C600 VDD.n451 GND 0.00418f
C601 VDD.n452 GND 0.00418f
C602 VDD.n453 GND 0.00418f
C603 VDD.n454 GND 0.00418f
C604 VDD.n455 GND 0.322f
C605 VDD.n456 GND 0.00418f
C606 VDD.n457 GND 0.00418f
C607 VDD.n458 GND 0.00418f
C608 VDD.n459 GND 0.00418f
C609 VDD.n460 GND 0.00418f
C610 VDD.n461 GND 0.322f
C611 VDD.n462 GND 0.00418f
C612 VDD.n463 GND 0.00418f
C613 VDD.n464 GND 0.00418f
C614 VDD.n465 GND 0.00418f
C615 VDD.n466 GND 0.00418f
C616 VDD.n467 GND 0.322f
C617 VDD.n468 GND 0.00418f
C618 VDD.n469 GND 0.00418f
C619 VDD.n470 GND 0.00418f
C620 VDD.n471 GND 0.00418f
C621 VDD.n472 GND 0.00418f
C622 VDD.n473 GND 0.25097f
C623 VDD.n474 GND 0.00418f
C624 VDD.n475 GND 0.00418f
C625 VDD.n476 GND 0.00418f
C626 VDD.n477 GND 0.00418f
C627 VDD.n478 GND 0.00418f
C628 VDD.n479 GND 0.322f
C629 VDD.n480 GND 0.00418f
C630 VDD.n481 GND 0.00418f
C631 VDD.t107 GND 0.161f
C632 VDD.n482 GND 0.00418f
C633 VDD.n483 GND 0.00418f
C634 VDD.n484 GND 0.00418f
C635 VDD.t130 GND 0.161f
C636 VDD.n485 GND 0.00418f
C637 VDD.n486 GND 0.00418f
C638 VDD.n487 GND 0.00418f
C639 VDD.n488 GND 0.00418f
C640 VDD.n489 GND 0.00418f
C641 VDD.n490 GND 0.322f
C642 VDD.n491 GND 0.00418f
C643 VDD.n492 GND 0.00418f
C644 VDD.n493 GND 0.312529f
C645 VDD.n494 GND 0.00418f
C646 VDD.n495 GND 0.00418f
C647 VDD.n496 GND 0.00418f
C648 VDD.n497 GND 0.322f
C649 VDD.n498 GND 0.00418f
C650 VDD.n499 GND 0.00418f
C651 VDD.n500 GND 0.00418f
C652 VDD.n501 GND 0.00418f
C653 VDD.n502 GND 0.00418f
C654 VDD.n503 GND 0.322f
C655 VDD.n504 GND 0.00418f
C656 VDD.n505 GND 0.00418f
C657 VDD.n506 GND 0.00418f
C658 VDD.n507 GND 0.00418f
C659 VDD.n508 GND 0.00418f
C660 VDD.n509 GND 0.322f
C661 VDD.n510 GND 0.00418f
C662 VDD.n511 GND 0.00418f
C663 VDD.n512 GND 0.00418f
C664 VDD.n513 GND 0.00418f
C665 VDD.n514 GND 0.00418f
C666 VDD.n515 GND 0.322f
C667 VDD.n516 GND 0.00418f
C668 VDD.n517 GND 0.00418f
C669 VDD.n518 GND 0.00418f
C670 VDD.n519 GND 0.00418f
C671 VDD.n520 GND 0.00418f
C672 VDD.n521 GND 0.322f
C673 VDD.n522 GND 0.00418f
C674 VDD.n523 GND 0.00418f
C675 VDD.n524 GND 0.00418f
C676 VDD.n525 GND 0.00418f
C677 VDD.n526 GND 0.00418f
C678 VDD.n527 GND 0.322f
C679 VDD.n528 GND 0.00418f
C680 VDD.n529 GND 0.00418f
C681 VDD.n530 GND 0.00418f
C682 VDD.n531 GND 0.00418f
C683 VDD.n532 GND 0.00418f
C684 VDD.t114 GND 0.161f
C685 VDD.n533 GND 0.00418f
C686 VDD.n534 GND 0.00418f
C687 VDD.n535 GND 0.00418f
C688 VDD.n536 GND 0.00418f
C689 VDD.n537 GND 0.00418f
C690 VDD.n538 GND 0.179941f
C691 VDD.n539 GND 0.00418f
C692 VDD.n540 GND 0.00418f
C693 VDD.n541 GND 0.222559f
C694 VDD.n542 GND 0.00418f
C695 VDD.n543 GND 0.00418f
C696 VDD.n544 GND 0.00418f
C697 VDD.n545 GND 0.322f
C698 VDD.n546 GND 0.00418f
C699 VDD.n547 GND 0.00418f
C700 VDD.t95 GND 0.161f
C701 VDD.n548 GND 0.00418f
C702 VDD.n549 GND 0.00418f
C703 VDD.n550 GND 0.00418f
C704 VDD.n551 GND 0.322f
C705 VDD.n552 GND 0.00418f
C706 VDD.n553 GND 0.00418f
C707 VDD.n554 GND 0.00418f
C708 VDD.n555 GND 0.00418f
C709 VDD.n556 GND 0.00418f
C710 VDD.n557 GND 0.322f
C711 VDD.n558 GND 0.00418f
C712 VDD.n559 GND 0.00418f
C713 VDD.n560 GND 0.00418f
C714 VDD.n561 GND 0.00418f
C715 VDD.n562 GND 0.00418f
C716 VDD.n563 GND 0.322f
C717 VDD.n564 GND 0.00418f
C718 VDD.n565 GND 0.00418f
C719 VDD.n566 GND 0.00418f
C720 VDD.n567 GND 0.00418f
C721 VDD.n568 GND 0.00418f
C722 VDD.n569 GND 0.322f
C723 VDD.n570 GND 0.00418f
C724 VDD.n571 GND 0.00418f
C725 VDD.n572 GND 0.00418f
C726 VDD.n573 GND 0.00418f
C727 VDD.n574 GND 0.00418f
C728 VDD.n575 GND 0.322f
C729 VDD.n576 GND 0.00418f
C730 VDD.n577 GND 0.00418f
C731 VDD.n578 GND 0.00418f
C732 VDD.n579 GND 0.00418f
C733 VDD.n580 GND 0.00418f
C734 VDD.n581 GND 0.322f
C735 VDD.n582 GND 0.00418f
C736 VDD.n583 GND 0.00418f
C737 VDD.n584 GND 0.00418f
C738 VDD.n585 GND 0.00418f
C739 VDD.n586 GND 0.00418f
C740 VDD.n587 GND 0.322f
C741 VDD.n588 GND 0.00418f
C742 VDD.n589 GND 0.00418f
C743 VDD.n590 GND 0.00418f
C744 VDD.n591 GND 0.00418f
C745 VDD.n592 GND 0.00418f
C746 VDD.n593 GND 0.322f
C747 VDD.n594 GND 0.00418f
C748 VDD.n595 GND 0.00418f
C749 VDD.n596 GND 0.00418f
C750 VDD.n597 GND 0.00418f
C751 VDD.n598 GND 0.00418f
C752 VDD.t128 GND 0.161f
C753 VDD.n599 GND 0.00418f
C754 VDD.n600 GND 0.00418f
C755 VDD.n601 GND 0.00418f
C756 VDD.n602 GND 0.00418f
C757 VDD.n603 GND 0.00418f
C758 VDD.n604 GND 0.322f
C759 VDD.n605 GND 0.00418f
C760 VDD.n606 GND 0.00418f
C761 VDD.t50 GND 0.161f
C762 VDD.n607 GND 0.00418f
C763 VDD.n608 GND 0.00418f
C764 VDD.n609 GND 0.00418f
C765 VDD.n610 GND 0.322f
C766 VDD.n611 GND 0.00418f
C767 VDD.n612 GND 0.00418f
C768 VDD.n613 GND 0.00418f
C769 VDD.n614 GND 0.00418f
C770 VDD.n615 GND 0.00418f
C771 VDD.n616 GND 0.322f
C772 VDD.n617 GND 0.00418f
C773 VDD.n618 GND 0.00418f
C774 VDD.n619 GND 0.00418f
C775 VDD.n620 GND 0.00418f
C776 VDD.n621 GND 0.00418f
C777 VDD.n622 GND 0.322f
C778 VDD.n623 GND 0.00418f
C779 VDD.n624 GND 0.00418f
C780 VDD.n625 GND 0.00418f
C781 VDD.n626 GND 0.00418f
C782 VDD.n627 GND 0.00418f
C783 VDD.n628 GND 0.322f
C784 VDD.n629 GND 0.00418f
C785 VDD.n630 GND 0.00418f
C786 VDD.n631 GND 0.00418f
C787 VDD.n632 GND 0.008807f
C788 VDD.n633 GND 0.008807f
C789 VDD.n634 GND 0.447485f
C790 VDD.n635 GND 0.00418f
C791 VDD.n636 GND 0.00418f
C792 VDD.n637 GND 0.008807f
C793 VDD.n638 GND 0.00418f
C794 VDD.n639 GND 0.00418f
C795 VDD.n640 GND 0.447485f
C796 VDD.n658 GND 0.009514f
C797 VDD.n659 GND 0.008807f
C798 VDD.n660 GND 0.00418f
C799 VDD.n661 GND 0.008807f
C800 VDD.t30 GND 0.089111f
C801 VDD.t28 GND 0.44554f
C802 VDD.n662 GND 0.076053f
C803 VDD.t31 GND 0.056759f
C804 VDD.n663 GND 0.078134f
C805 VDD.n664 GND 0.00418f
C806 VDD.n665 GND 0.00418f
C807 VDD.n666 GND 0.322f
C808 VDD.n667 GND 0.00418f
C809 VDD.n668 GND 0.00418f
C810 VDD.n669 GND 0.00418f
C811 VDD.n670 GND 0.008807f
C812 VDD.n671 GND 0.00418f
C813 VDD.t40 GND 0.089111f
C814 VDD.t39 GND 0.44554f
C815 VDD.n672 GND 0.076053f
C816 VDD.t41 GND 0.056759f
C817 VDD.n673 GND 0.078134f
C818 VDD.n674 GND 0.005158f
C819 VDD.n675 GND 0.00418f
C820 VDD.n676 GND 0.00418f
C821 VDD.n677 GND 0.322f
C822 VDD.n678 GND 0.00418f
C823 VDD.n679 GND 0.00418f
C824 VDD.n680 GND 0.00418f
C825 VDD.n681 GND 0.00418f
C826 VDD.n682 GND 0.00418f
C827 VDD.n683 GND 0.322f
C828 VDD.n684 GND 0.00418f
C829 VDD.n685 GND 0.00418f
C830 VDD.n686 GND 0.00418f
C831 VDD.n687 GND 0.00418f
C832 VDD.n688 GND 0.00418f
C833 VDD.n689 GND 0.00418f
C834 VDD.n690 GND 0.322f
C835 VDD.n691 GND 0.00418f
C836 VDD.n692 GND 0.00418f
C837 VDD.n693 GND 0.00418f
C838 VDD.n694 GND 0.00418f
C839 VDD.n695 GND 0.00418f
C840 VDD.n696 GND 0.322f
C841 VDD.n697 GND 0.00418f
C842 VDD.n698 GND 0.00418f
C843 VDD.n699 GND 0.00418f
C844 VDD.n700 GND 0.00418f
C845 VDD.n701 GND 0.00418f
C846 VDD.t29 GND 0.161f
C847 VDD.n702 GND 0.00418f
C848 VDD.n703 GND 0.00418f
C849 VDD.n704 GND 0.00418f
C850 VDD.n705 GND 0.00418f
C851 VDD.n706 GND 0.00418f
C852 VDD.n707 GND 0.322f
C853 VDD.n708 GND 0.00418f
C854 VDD.n709 GND 0.00418f
C855 VDD.t124 GND 0.161f
C856 VDD.n710 GND 0.00418f
C857 VDD.n711 GND 0.00418f
C858 VDD.n712 GND 0.00418f
C859 VDD.n713 GND 0.322f
C860 VDD.n714 GND 0.00418f
C861 VDD.n715 GND 0.00418f
C862 VDD.n716 GND 0.00418f
C863 VDD.n717 GND 0.00418f
C864 VDD.n718 GND 0.00418f
C865 VDD.n719 GND 0.322f
C866 VDD.n720 GND 0.00418f
C867 VDD.n721 GND 0.00418f
C868 VDD.n722 GND 0.00418f
C869 VDD.n723 GND 0.00418f
C870 VDD.n724 GND 0.00418f
C871 VDD.n725 GND 0.322f
C872 VDD.n726 GND 0.00418f
C873 VDD.n727 GND 0.00418f
C874 VDD.n728 GND 0.00418f
C875 VDD.n729 GND 0.00418f
C876 VDD.n730 GND 0.00418f
C877 VDD.n731 GND 0.322f
C878 VDD.n732 GND 0.00418f
C879 VDD.n733 GND 0.00418f
C880 VDD.n734 GND 0.00418f
C881 VDD.n735 GND 0.00418f
C882 VDD.n736 GND 0.00418f
C883 VDD.n737 GND 0.322f
C884 VDD.n738 GND 0.00418f
C885 VDD.n739 GND 0.00418f
C886 VDD.n740 GND 0.00418f
C887 VDD.n741 GND 0.00418f
C888 VDD.n742 GND 0.00418f
C889 VDD.n743 GND 0.322f
C890 VDD.n744 GND 0.00418f
C891 VDD.n745 GND 0.00418f
C892 VDD.n746 GND 0.00418f
C893 VDD.n747 GND 0.00418f
C894 VDD.n748 GND 0.00418f
C895 VDD.n749 GND 0.322f
C896 VDD.n750 GND 0.00418f
C897 VDD.n751 GND 0.00418f
C898 VDD.n752 GND 0.00418f
C899 VDD.n753 GND 0.00418f
C900 VDD.n754 GND 0.00418f
C901 VDD.n755 GND 0.322f
C902 VDD.n756 GND 0.00418f
C903 VDD.n757 GND 0.00418f
C904 VDD.n758 GND 0.00418f
C905 VDD.n759 GND 0.00418f
C906 VDD.n760 GND 0.00418f
C907 VDD.t97 GND 0.161f
C908 VDD.n761 GND 0.00418f
C909 VDD.n762 GND 0.00418f
C910 VDD.n763 GND 0.00418f
C911 VDD.n764 GND 0.00418f
C912 VDD.n765 GND 0.00418f
C913 VDD.n766 GND 0.222559f
C914 VDD.n767 GND 0.00418f
C915 VDD.n768 GND 0.00418f
C916 VDD.n769 GND 0.179941f
C917 VDD.n770 GND 0.00418f
C918 VDD.n771 GND 0.00418f
C919 VDD.n772 GND 0.00418f
C920 VDD.n773 GND 0.322f
C921 VDD.n774 GND 0.00418f
C922 VDD.n775 GND 0.00418f
C923 VDD.t108 GND 0.161f
C924 VDD.n776 GND 0.00418f
C925 VDD.n777 GND 0.00418f
C926 VDD.n778 GND 0.00418f
C927 VDD.n779 GND 0.322f
C928 VDD.n780 GND 0.00418f
C929 VDD.n781 GND 0.00418f
C930 VDD.n782 GND 0.00418f
C931 VDD.n783 GND 0.00418f
C932 VDD.n784 GND 0.00418f
C933 VDD.n785 GND 0.322f
C934 VDD.n786 GND 0.00418f
C935 VDD.n787 GND 0.00418f
C936 VDD.n788 GND 0.00418f
C937 VDD.n789 GND 0.00418f
C938 VDD.n790 GND 0.00418f
C939 VDD.n791 GND 0.322f
C940 VDD.n792 GND 0.00418f
C941 VDD.n793 GND 0.00418f
C942 VDD.n794 GND 0.00418f
C943 VDD.n795 GND 0.00418f
C944 VDD.n796 GND 0.00418f
C945 VDD.n797 GND 0.322f
C946 VDD.n798 GND 0.00418f
C947 VDD.n799 GND 0.00418f
C948 VDD.n800 GND 0.00418f
C949 VDD.n801 GND 0.00418f
C950 VDD.n802 GND 0.00418f
C951 VDD.n803 GND 0.322f
C952 VDD.n804 GND 0.00418f
C953 VDD.n805 GND 0.00418f
C954 VDD.n806 GND 0.00418f
C955 VDD.n807 GND 0.00418f
C956 VDD.n808 GND 0.00418f
C957 VDD.n809 GND 0.322f
C958 VDD.n810 GND 0.00418f
C959 VDD.n811 GND 0.00418f
C960 VDD.n812 GND 0.00418f
C961 VDD.n813 GND 0.00418f
C962 VDD.n814 GND 0.00418f
C963 VDD.n815 GND 0.312529f
C964 VDD.n816 GND 0.00418f
C965 VDD.n817 GND 0.00418f
C966 VDD.n818 GND 0.00418f
C967 VDD.n819 GND 0.00418f
C968 VDD.n820 GND 0.00418f
C969 VDD.n821 GND 0.322f
C970 VDD.n822 GND 0.00418f
C971 VDD.n823 GND 0.00418f
C972 VDD.t126 GND 0.161f
C973 VDD.n824 GND 0.00418f
C974 VDD.n825 GND 0.00418f
C975 VDD.n826 GND 0.00418f
C976 VDD.t111 GND 0.161f
C977 VDD.n827 GND 0.00418f
C978 VDD.n828 GND 0.00418f
C979 VDD.n829 GND 0.00418f
C980 VDD.n830 GND 0.00418f
C981 VDD.n831 GND 0.00418f
C982 VDD.n832 GND 0.322f
C983 VDD.n833 GND 0.00418f
C984 VDD.n834 GND 0.00418f
C985 VDD.n835 GND 0.25097f
C986 VDD.n836 GND 0.00418f
C987 VDD.n837 GND 0.00418f
C988 VDD.n838 GND 0.00418f
C989 VDD.n839 GND 0.322f
C990 VDD.n840 GND 0.00418f
C991 VDD.n841 GND 0.00418f
C992 VDD.n842 GND 0.00418f
C993 VDD.n843 GND 0.00418f
C994 VDD.n844 GND 0.00418f
C995 VDD.n845 GND 0.322f
C996 VDD.n846 GND 0.00418f
C997 VDD.n847 GND 0.00418f
C998 VDD.n848 GND 0.00418f
C999 VDD.n849 GND 0.00418f
C1000 VDD.n850 GND 0.00418f
C1001 VDD.n851 GND 0.322f
C1002 VDD.n852 GND 0.00418f
C1003 VDD.n853 GND 0.00418f
C1004 VDD.n854 GND 0.00418f
C1005 VDD.n855 GND 0.00418f
C1006 VDD.n856 GND 0.00418f
C1007 VDD.n857 GND 0.322f
C1008 VDD.n858 GND 0.00418f
C1009 VDD.n859 GND 0.00418f
C1010 VDD.n860 GND 0.00418f
C1011 VDD.n861 GND 0.00418f
C1012 VDD.n862 GND 0.00418f
C1013 VDD.n863 GND 0.322f
C1014 VDD.n864 GND 0.00418f
C1015 VDD.n865 GND 0.00418f
C1016 VDD.n866 GND 0.00418f
C1017 VDD.n867 GND 0.00418f
C1018 VDD.n868 GND 0.00418f
C1019 VDD.n869 GND 0.322f
C1020 VDD.n870 GND 0.00418f
C1021 VDD.n871 GND 0.00418f
C1022 VDD.n872 GND 0.00418f
C1023 VDD.n873 GND 0.00418f
C1024 VDD.n874 GND 0.00418f
C1025 VDD.t92 GND 0.322f
C1026 VDD.n875 GND 0.00418f
C1027 VDD.n876 GND 0.00418f
C1028 VDD.n877 GND 0.00418f
C1029 VDD.n878 GND 0.00418f
C1030 VDD.n879 GND 0.00418f
C1031 VDD.n880 GND 0.2415f
C1032 VDD.n881 GND 0.00418f
C1033 VDD.n882 GND 0.00418f
C1034 VDD.n883 GND 0.00418f
C1035 VDD.n884 GND 0.00418f
C1036 VDD.n885 GND 0.00418f
C1037 VDD.n886 GND 0.322f
C1038 VDD.n887 GND 0.00418f
C1039 VDD.n888 GND 0.00418f
C1040 VDD.t104 GND 0.161f
C1041 VDD.n889 GND 0.00418f
C1042 VDD.n890 GND 0.00418f
C1043 VDD.n891 GND 0.00418f
C1044 VDD.n892 GND 0.322f
C1045 VDD.n893 GND 0.00418f
C1046 VDD.n894 GND 0.00418f
C1047 VDD.n895 GND 0.00418f
C1048 VDD.n896 GND 0.00418f
C1049 VDD.n897 GND 0.00418f
C1050 VDD.n898 GND 0.322f
C1051 VDD.n899 GND 0.00418f
C1052 VDD.n900 GND 0.00418f
C1053 VDD.n901 GND 0.00418f
C1054 VDD.n902 GND 0.00418f
C1055 VDD.n903 GND 0.00418f
C1056 VDD.n904 GND 0.322f
C1057 VDD.n905 GND 0.00418f
C1058 VDD.n906 GND 0.00418f
C1059 VDD.n907 GND 0.00418f
C1060 VDD.n908 GND 0.00418f
C1061 VDD.n909 GND 0.00418f
C1062 VDD.n910 GND 0.322f
C1063 VDD.n911 GND 0.00418f
C1064 VDD.n912 GND 0.00418f
C1065 VDD.n913 GND 0.00418f
C1066 VDD.n914 GND 0.00418f
C1067 VDD.n915 GND 0.00418f
C1068 VDD.n916 GND 0.322f
C1069 VDD.n917 GND 0.00418f
C1070 VDD.n918 GND 0.00418f
C1071 VDD.n919 GND 0.00418f
C1072 VDD.n920 GND 0.00418f
C1073 VDD.n921 GND 0.00418f
C1074 VDD.n922 GND 0.322f
C1075 VDD.n923 GND 0.00418f
C1076 VDD.n924 GND 0.00418f
C1077 VDD.n925 GND 0.00418f
C1078 VDD.n926 GND 0.00418f
C1079 VDD.n927 GND 0.00418f
C1080 VDD.n928 GND 0.322f
C1081 VDD.n929 GND 0.00418f
C1082 VDD.n930 GND 0.00418f
C1083 VDD.n931 GND 0.00418f
C1084 VDD.n932 GND 0.00418f
C1085 VDD.n933 GND 0.00418f
C1086 VDD.n934 GND 0.322f
C1087 VDD.n935 GND 0.00418f
C1088 VDD.n936 GND 0.00418f
C1089 VDD.n937 GND 0.00418f
C1090 VDD.n938 GND 0.00418f
C1091 VDD.n939 GND 0.00418f
C1092 VDD.t119 GND 0.161f
C1093 VDD.n940 GND 0.00418f
C1094 VDD.n941 GND 0.00418f
C1095 VDD.n942 GND 0.00418f
C1096 VDD.n943 GND 0.00418f
C1097 VDD.n944 GND 0.00418f
C1098 VDD.n945 GND 0.322f
C1099 VDD.n946 GND 0.00418f
C1100 VDD.n947 GND 0.00418f
C1101 VDD.n948 GND 0.232029f
C1102 VDD.n949 GND 0.00418f
C1103 VDD.n950 GND 0.00418f
C1104 VDD.n951 GND 0.00418f
C1105 VDD.n952 GND 0.322f
C1106 VDD.n953 GND 0.00418f
C1107 VDD.n954 GND 0.00418f
C1108 VDD.n955 GND 0.00418f
C1109 VDD.n956 GND 0.00418f
C1110 VDD.n957 GND 0.00418f
C1111 VDD.n958 GND 0.198882f
C1112 VDD.n959 GND 0.00418f
C1113 VDD.n960 GND 0.00418f
C1114 VDD.n961 GND 0.00418f
C1115 VDD.n962 GND 0.00418f
C1116 VDD.n963 GND 0.00418f
C1117 VDD.n964 GND 0.322f
C1118 VDD.n965 GND 0.00418f
C1119 VDD.n966 GND 0.00418f
C1120 VDD.t99 GND 0.161f
C1121 VDD.n967 GND 0.00418f
C1122 VDD.n968 GND 0.00418f
C1123 VDD.n969 GND 0.00418f
C1124 VDD.n970 GND 0.322f
C1125 VDD.n971 GND 0.00418f
C1126 VDD.n972 GND 0.00418f
C1127 VDD.n973 GND 0.00418f
C1128 VDD.n974 GND 0.00418f
C1129 VDD.n975 GND 0.00418f
C1130 VDD.n976 GND 0.322f
C1131 VDD.n977 GND 0.00418f
C1132 VDD.n978 GND 0.00418f
C1133 VDD.n979 GND 0.00418f
C1134 VDD.n980 GND 0.00418f
C1135 VDD.n981 GND 0.00418f
C1136 VDD.n982 GND 0.322f
C1137 VDD.n983 GND 0.00418f
C1138 VDD.n984 GND 0.00418f
C1139 VDD.n985 GND 0.00418f
C1140 VDD.n986 GND 0.00418f
C1141 VDD.n987 GND 0.00418f
C1142 VDD.n988 GND 0.322f
C1143 VDD.n989 GND 0.00418f
C1144 VDD.n990 GND 0.00418f
C1145 VDD.n991 GND 0.00418f
C1146 VDD.n992 GND 0.00418f
C1147 VDD.n993 GND 0.00418f
C1148 VDD.n994 GND 0.260441f
C1149 VDD.n995 GND 0.00418f
C1150 VDD.n996 GND 0.00418f
C1151 VDD.n997 GND 0.00418f
C1152 VDD.n998 GND 0.00418f
C1153 VDD.n999 GND 0.00418f
C1154 VDD.n1000 GND 0.322f
C1155 VDD.n1001 GND 0.00418f
C1156 VDD.n1002 GND 0.00418f
C1157 VDD.t121 GND 0.161f
C1158 VDD.n1003 GND 0.00418f
C1159 VDD.n1004 GND 0.00418f
C1160 VDD.n1005 GND 0.00418f
C1161 VDD.n1006 GND 0.322f
C1162 VDD.n1007 GND 0.00418f
C1163 VDD.n1008 GND 0.00418f
C1164 VDD.n1009 GND 0.00418f
C1165 VDD.n1010 GND 0.00418f
C1166 VDD.n1011 GND 0.00418f
C1167 VDD.n1012 GND 0.322f
C1168 VDD.n1013 GND 0.00418f
C1169 VDD.n1014 GND 0.00418f
C1170 VDD.n1015 GND 0.00418f
C1171 VDD.n1016 GND 0.00418f
C1172 VDD.n1017 GND 0.00418f
C1173 VDD.t109 GND 0.161f
C1174 VDD.n1018 GND 0.00418f
C1175 VDD.n1019 GND 0.00418f
C1176 VDD.n1020 GND 0.00418f
C1177 VDD.n1021 GND 0.00418f
C1178 VDD.n1022 GND 0.00418f
C1179 VDD.n1023 GND 0.322f
C1180 VDD.n1024 GND 0.00418f
C1181 VDD.n1025 GND 0.00418f
C1182 VDD.n1026 GND 0.274647f
C1183 VDD.n1027 GND 0.00418f
C1184 VDD.n1028 GND 0.00418f
C1185 VDD.n1029 GND 0.00418f
C1186 VDD.n1030 GND 0.322f
C1187 VDD.n1031 GND 0.00418f
C1188 VDD.n1032 GND 0.00418f
C1189 VDD.n1033 GND 0.00418f
C1190 VDD.n1034 GND 0.00418f
C1191 VDD.n1035 GND 0.00418f
C1192 VDD.n1036 GND 0.322f
C1193 VDD.n1037 GND 0.00418f
C1194 VDD.n1038 GND 0.00418f
C1195 VDD.n1039 GND 0.00418f
C1196 VDD.n1040 GND 0.00418f
C1197 VDD.n1041 GND 0.00418f
C1198 VDD.n1042 GND 0.322f
C1199 VDD.n1043 GND 0.00418f
C1200 VDD.n1044 GND 0.00418f
C1201 VDD.n1045 GND 0.00418f
C1202 VDD.n1046 GND 0.00418f
C1203 VDD.n1047 GND 0.00418f
C1204 VDD.n1048 GND 0.322f
C1205 VDD.n1049 GND 0.00418f
C1206 VDD.n1050 GND 0.00418f
C1207 VDD.n1051 GND 0.00418f
C1208 VDD.n1052 GND 0.00418f
C1209 VDD.n1053 GND 0.00418f
C1210 VDD.n1054 GND 0.322f
C1211 VDD.n1055 GND 0.00418f
C1212 VDD.n1056 GND 0.00418f
C1213 VDD.n1057 GND 0.00418f
C1214 VDD.n1058 GND 0.00418f
C1215 VDD.n1059 GND 0.00418f
C1216 VDD.n1060 GND 0.322f
C1217 VDD.n1061 GND 0.00418f
C1218 VDD.n1062 GND 0.00418f
C1219 VDD.n1063 GND 0.00418f
C1220 VDD.n1064 GND 0.00418f
C1221 VDD.n1065 GND 0.00418f
C1222 VDD.t22 GND 0.161f
C1223 VDD.n1066 GND 0.00418f
C1224 VDD.n1067 GND 0.00418f
C1225 VDD.n1068 GND 0.00418f
C1226 VDD.n1069 GND 0.00418f
C1227 VDD.n1070 GND 0.00418f
C1228 VDD.n1071 GND 0.217823f
C1229 VDD.n1072 GND 0.00418f
C1230 VDD.n1073 GND 0.00418f
C1231 VDD.n1074 GND 0.184676f
C1232 VDD.n1075 GND 0.00418f
C1233 VDD.n1076 GND 0.00418f
C1234 VDD.n1077 GND 0.00418f
C1235 VDD.n1078 GND 0.322f
C1236 VDD.n1079 GND 0.00418f
C1237 VDD.n1080 GND 0.00418f
C1238 VDD.t117 GND 0.161f
C1239 VDD.n1081 GND 0.00418f
C1240 VDD.n1082 GND 0.00418f
C1241 VDD.n1083 GND 0.00418f
C1242 VDD.n1084 GND 0.322f
C1243 VDD.n1085 GND 0.00418f
C1244 VDD.n1086 GND 0.00418f
C1245 VDD.n1087 GND 0.00418f
C1246 VDD.n1088 GND 0.00418f
C1247 VDD.n1089 GND 0.00418f
C1248 VDD.n1090 GND 0.322f
C1249 VDD.n1091 GND 0.00418f
C1250 VDD.n1092 GND 0.00418f
C1251 VDD.n1093 GND 0.00418f
C1252 VDD.n1094 GND 0.00418f
C1253 VDD.n1095 GND 0.00418f
C1254 VDD.n1096 GND 0.322f
C1255 VDD.n1097 GND 0.00418f
C1256 VDD.n1098 GND 0.00418f
C1257 VDD.n1099 GND 0.00418f
C1258 VDD.n1100 GND 0.009514f
C1259 VDD.n1101 GND 0.009514f
C1260 VDD.n1102 GND 1.67629f
C1261 VDD.n1103 GND 0.008807f
C1262 VDD.n1104 GND 0.008807f
C1263 VDD.n1105 GND 0.009514f
C1264 VDD.n1106 GND 0.00418f
C1265 VDD.n1108 GND 0.00418f
C1266 VDD.n1109 GND 0.00418f
C1267 VDD.n1110 GND 0.063036f
C1268 VDD.n1112 GND 0.00418f
C1269 VDD.n1113 GND 0.00418f
C1270 VDD.t24 GND 0.089111f
C1271 VDD.t21 GND 0.44554f
C1272 VDD.n1114 GND 0.076053f
C1273 VDD.t23 GND 0.056759f
C1274 VDD.n1115 GND 0.078134f
C1275 VDD.n1116 GND 0.00418f
C1276 VDD.n1117 GND 0.009514f
C1277 VDD.n1118 GND 0.00418f
C1278 VDD.n1119 GND 0.00418f
C1279 VDD.n1120 GND 0.00418f
C1280 VDD.n1121 GND 0.00418f
C1281 VDD.n1122 GND 0.00418f
C1282 VDD.n1123 GND 0.00418f
C1283 VDD.n1124 GND 0.00418f
C1284 VDD.n1125 GND 0.00418f
C1285 VDD.n1126 GND 0.00418f
C1286 VDD.n1127 GND 0.00418f
C1287 VDD.n1128 GND 0.00418f
C1288 VDD.n1129 GND 0.00418f
C1289 VDD.n1130 GND 0.00418f
C1290 VDD.n1131 GND 0.00418f
C1291 VDD.n1132 GND 0.00418f
C1292 VDD.n1133 GND 0.00418f
C1293 VDD.t82 GND 0.089111f
C1294 VDD.t80 GND 0.44554f
C1295 VDD.n1134 GND 0.076053f
C1296 VDD.t81 GND 0.056759f
C1297 VDD.n1135 GND 0.078134f
C1298 VDD.n1136 GND 0.00418f
C1299 VDD.n1137 GND 0.00418f
C1300 VDD.n1138 GND 0.003935f
C1301 VDD.n1139 GND 0.005287f
C1302 VDD.n1141 GND 0.004948f
C1303 VDD.t90 GND 0.085164f
C1304 VDD.t89 GND 0.430073f
C1305 VDD.n1142 GND 0.075426f
C1306 VDD.t91 GND 0.053191f
C1307 VDD.n1143 GND 0.077435f
C1308 VDD.n1144 GND 0.009278f
C1309 VDD.n1145 GND 0.006148f
C1310 VDD.t112 GND 5.13068f
C1311 VDD.t147 GND 7.35153f
C1312 VDD.n1146 GND 4.04394f
C1313 VDD.n1147 GND 0.004948f
C1314 VDD.n1148 GND 0.006148f
C1315 VDD.n1149 GND 0.006148f
C1316 VDD.n1150 GND 0.004948f
C1317 VDD.n1152 GND 0.006148f
C1318 VDD.n1153 GND 0.006148f
C1319 VDD.n1154 GND 0.006148f
C1320 VDD.n1155 GND 0.006148f
C1321 VDD.n1156 GND 0.006148f
C1322 VDD.n1157 GND 0.004082f
C1323 VDD.n1159 GND 0.006148f
C1324 VDD.n1160 GND 0.004181f
C1325 VDD.t84 GND 0.085164f
C1326 VDD.t83 GND 0.430073f
C1327 VDD.n1161 GND 0.075426f
C1328 VDD.t85 GND 0.053191f
C1329 VDD.n1162 GND 0.077435f
C1330 VDD.n1163 GND 0.006148f
C1331 VDD.n1164 GND 0.006148f
C1332 VDD.n1165 GND 0.004948f
C1333 VDD.n1167 GND 0.006148f
C1334 VDD.n1168 GND 0.006148f
C1335 VDD.n1169 GND 0.006148f
C1336 VDD.n1170 GND 0.006148f
C1337 VDD.n1171 GND 0.004948f
C1338 VDD.n1173 GND 0.006148f
C1339 VDD.n1174 GND 0.006148f
C1340 VDD.n1175 GND 0.006148f
C1341 VDD.n1176 GND 0.006148f
C1342 VDD.n1177 GND 0.006148f
C1343 VDD.n1178 GND 0.00339f
C1344 VDD.n1180 GND 0.006148f
C1345 VDD.n1181 GND 0.004874f
C1346 VDD.t72 GND 0.085164f
C1347 VDD.t71 GND 0.430073f
C1348 VDD.n1182 GND 0.075426f
C1349 VDD.t73 GND 0.053191f
C1350 VDD.n1183 GND 0.077435f
C1351 VDD.n1184 GND 0.006148f
C1352 VDD.n1185 GND 0.006148f
C1353 VDD.n1186 GND 0.004948f
C1354 VDD.n1188 GND 0.006148f
C1355 VDD.n1189 GND 0.006148f
C1356 VDD.n1190 GND 0.006148f
C1357 VDD.n1191 GND 0.006148f
C1358 VDD.n1192 GND 0.004948f
C1359 VDD.n1194 GND 0.006148f
C1360 VDD.n1195 GND 0.006148f
C1361 VDD.n1196 GND 0.006148f
C1362 VDD.n1197 GND 0.006148f
C1363 VDD.n1198 GND 0.005287f
C1364 VDD.n1199 GND 0.002697f
C1365 VDD.n1201 GND 0.006148f
C1366 VDD.t75 GND 0.085164f
C1367 VDD.t74 GND 0.430073f
C1368 VDD.n1202 GND 0.075426f
C1369 VDD.t76 GND 0.053191f
C1370 VDD.n1203 GND 0.077435f
C1371 VDD.n1204 GND 0.006804f
C1372 VDD.n1205 GND 0.004948f
C1373 VDD.n1206 GND 0.004948f
C1374 VDD.n1207 GND 0.006148f
C1375 VDD.n1209 GND 0.006148f
C1376 VDD.n1210 GND 0.006148f
C1377 VDD.n1212 GND 0.006148f
C1378 VDD.n1213 GND 0.006148f
C1379 VDD.n1214 GND 0.004948f
C1380 VDD.n1215 GND 0.006148f
C1381 VDD.n1217 GND 0.006148f
C1382 VDD.n1218 GND 0.006148f
C1383 VDD.n1220 GND 0.006148f
C1384 VDD.n1221 GND 0.006148f
C1385 VDD.n1222 GND 0.004478f
C1386 VDD.n1223 GND 0.014117f
C1387 VDD.n1224 GND 0.002944f
C1388 VDD.t34 GND 0.085164f
C1389 VDD.t32 GND 0.430073f
C1390 VDD.n1225 GND 0.075426f
C1391 VDD.t35 GND 0.053191f
C1392 VDD.n1226 GND 0.077435f
C1393 VDD.n1228 GND 0.006148f
C1394 VDD.n1229 GND 0.006148f
C1395 VDD.n1230 GND 0.004107f
C1396 VDD.n1231 GND 0.473529f
C1397 VDD.n1232 GND 0.006148f
C1398 VDD.n1233 GND 0.014117f
C1399 VDD.n1234 GND 0.004948f
C1400 VDD.n1235 GND 0.006148f
C1401 VDD.n1236 GND 0.004948f
C1402 VDD.n1237 GND 0.006148f
C1403 VDD.n1238 GND 0.473529f
C1404 VDD.n1239 GND 0.006148f
C1405 VDD.n1240 GND 0.004948f
C1406 VDD.n1241 GND 0.004948f
C1407 VDD.n1242 GND 0.006148f
C1408 VDD.n1243 GND 0.004948f
C1409 VDD.n1244 GND 0.006148f
C1410 VDD.n1245 GND 0.473529f
C1411 VDD.n1246 GND 0.006148f
C1412 VDD.n1247 GND 0.004948f
C1413 VDD.n1248 GND 0.006148f
C1414 VDD.n1249 GND 0.004948f
C1415 VDD.n1250 GND 0.006148f
C1416 VDD.t33 GND 0.473529f
C1417 VDD.n1251 GND 0.006148f
C1418 VDD.n1252 GND 0.004948f
C1419 VDD.n1253 GND 0.006148f
C1420 VDD.n1254 GND 0.004948f
C1421 VDD.n1255 GND 0.006148f
C1422 VDD.n1256 GND 0.473529f
C1423 VDD.n1257 GND 0.006148f
C1424 VDD.n1258 GND 0.004948f
C1425 VDD.n1259 GND 0.006148f
C1426 VDD.n1260 GND 0.004948f
C1427 VDD.n1261 GND 0.006148f
C1428 VDD.n1262 GND 0.473529f
C1429 VDD.n1263 GND 0.006148f
C1430 VDD.n1264 GND 0.004948f
C1431 VDD.n1265 GND 0.006148f
C1432 VDD.n1266 GND 0.004948f
C1433 VDD.n1267 GND 0.006148f
C1434 VDD.n1268 GND 0.473529f
C1435 VDD.n1269 GND 0.006148f
C1436 VDD.n1270 GND 0.004948f
C1437 VDD.n1271 GND 0.006148f
C1438 VDD.n1272 GND 0.004948f
C1439 VDD.n1273 GND 0.006148f
C1440 VDD.n1274 GND 0.473529f
C1441 VDD.n1275 GND 0.006148f
C1442 VDD.n1276 GND 0.004948f
C1443 VDD.n1277 GND 0.006148f
C1444 VDD.n1278 GND 0.004948f
C1445 VDD.n1279 GND 0.006148f
C1446 VDD.n1280 GND 0.473529f
C1447 VDD.n1281 GND 0.006148f
C1448 VDD.n1282 GND 0.004948f
C1449 VDD.n1283 GND 0.006148f
C1450 VDD.n1284 GND 0.004948f
C1451 VDD.n1285 GND 0.006148f
C1452 VDD.n1286 GND 0.473529f
C1453 VDD.n1287 GND 0.006148f
C1454 VDD.n1288 GND 0.004948f
C1455 VDD.n1289 GND 0.006148f
C1456 VDD.n1290 GND 0.004948f
C1457 VDD.n1291 GND 0.006148f
C1458 VDD.n1292 GND 0.473529f
C1459 VDD.n1293 GND 0.006148f
C1460 VDD.n1294 GND 0.004948f
C1461 VDD.t142 GND 0.071097f
C1462 VDD.t136 GND 0.069252f
C1463 VDD.n1295 GND 0.776551f
C1464 VDD.t141 GND 0.069252f
C1465 VDD.n1296 GND 0.424616f
C1466 VDD.t143 GND 0.069252f
C1467 VDD.n1297 GND 0.424616f
C1468 VDD.t144 GND 0.069252f
C1469 VDD.n1298 GND 0.506478f
C1470 VDD.n1299 GND 2.23977f
C1471 VDD.n1300 GND 0.136126f
C1472 VDD.n1301 GND 0.004948f
C1473 VDD.n1302 GND 0.006148f
C1474 VDD.t135 GND 0.473529f
C1475 VDD.n1303 GND 0.006148f
C1476 VDD.n1304 GND 0.004948f
C1477 VDD.n1305 GND 0.006148f
C1478 VDD.n1306 GND 0.004948f
C1479 VDD.n1307 GND 0.006148f
C1480 VDD.n1308 GND 0.473529f
C1481 VDD.n1309 GND 0.006148f
C1482 VDD.n1310 GND 0.004948f
C1483 VDD.n1311 GND 0.006148f
C1484 VDD.n1312 GND 0.004948f
C1485 VDD.n1313 GND 0.006148f
C1486 VDD.n1314 GND 0.473529f
C1487 VDD.n1315 GND 0.006148f
C1488 VDD.n1316 GND 0.004948f
C1489 VDD.n1317 GND 0.006148f
C1490 VDD.n1318 GND 0.004948f
C1491 VDD.n1319 GND 0.006148f
C1492 VDD.n1320 GND 0.473529f
C1493 VDD.n1321 GND 0.006148f
C1494 VDD.n1322 GND 0.004948f
C1495 VDD.n1323 GND 0.006148f
C1496 VDD.n1324 GND 0.004948f
C1497 VDD.n1325 GND 0.006148f
C1498 VDD.n1326 GND 0.473529f
C1499 VDD.n1327 GND 0.006148f
C1500 VDD.n1328 GND 0.004948f
C1501 VDD.n1329 GND 0.006148f
C1502 VDD.n1330 GND 0.004948f
C1503 VDD.n1331 GND 0.006148f
C1504 VDD.n1332 GND 0.473529f
C1505 VDD.n1333 GND 0.006148f
C1506 VDD.n1334 GND 0.004948f
C1507 VDD.n1335 GND 0.006148f
C1508 VDD.n1336 GND 0.004948f
C1509 VDD.n1337 GND 0.006148f
C1510 VDD.n1338 GND 0.473529f
C1511 VDD.n1339 GND 0.006148f
C1512 VDD.n1340 GND 0.004948f
C1513 VDD.n1341 GND 0.006148f
C1514 VDD.n1342 GND 0.004948f
C1515 VDD.n1343 GND 0.006148f
C1516 VDD.n1344 GND 0.473529f
C1517 VDD.n1345 GND 0.006148f
C1518 VDD.n1346 GND 0.004948f
C1519 VDD.n1347 GND 0.006148f
C1520 VDD.n1348 GND 0.004948f
C1521 VDD.n1349 GND 0.006148f
C1522 VDD.t1 GND 0.473529f
C1523 VDD.n1350 GND 0.006148f
C1524 VDD.n1351 GND 0.004948f
C1525 VDD.n1352 GND 0.006148f
C1526 VDD.n1353 GND 0.004948f
C1527 VDD.n1354 GND 0.006148f
C1528 VDD.n1355 GND 0.473529f
C1529 VDD.n1356 GND 0.006148f
C1530 VDD.n1357 GND 0.004948f
C1531 VDD.n1358 GND 0.006148f
C1532 VDD.n1359 GND 0.004948f
C1533 VDD.n1360 GND 0.006148f
C1534 VDD.n1361 GND 0.473529f
C1535 VDD.n1362 GND 0.006148f
C1536 VDD.n1363 GND 0.004948f
C1537 VDD.n1364 GND 0.006148f
C1538 VDD.n1365 GND 0.004948f
C1539 VDD.n1366 GND 0.006148f
C1540 VDD.n1367 GND 0.473529f
C1541 VDD.n1368 GND 0.006148f
C1542 VDD.n1369 GND 0.004948f
C1543 VDD.n1370 GND 0.014117f
C1544 VDD.n1371 GND 0.014117f
C1545 VDD.n1372 GND 1.09148f
C1546 VDD.n1373 GND 0.014117f
C1547 VDD.n1374 GND 0.006148f
C1548 VDD.n1375 GND 0.006148f
C1549 VDD.t6 GND 0.085164f
C1550 VDD.t4 GND 0.430073f
C1551 VDD.n1376 GND 0.075426f
C1552 VDD.t5 GND 0.053191f
C1553 VDD.n1377 GND 0.077435f
C1554 VDD.n1378 GND 0.004948f
C1555 VDD.n1380 GND 0.006148f
C1556 VDD.n1381 GND 0.006148f
C1557 VDD.n1382 GND 0.004948f
C1558 VDD.n1383 GND 0.006148f
C1559 VDD.n1384 GND 0.004948f
C1560 VDD.n1385 GND 0.006148f
C1561 VDD.n1386 GND 0.004948f
C1562 VDD.n1387 GND 0.006148f
C1563 VDD.n1388 GND 0.004948f
C1564 VDD.n1389 GND 0.006148f
C1565 VDD.t58 GND 0.085164f
C1566 VDD.t56 GND 0.430073f
C1567 VDD.n1390 GND 0.075426f
C1568 VDD.t57 GND 0.053191f
C1569 VDD.n1391 GND 0.077435f
C1570 VDD.n1392 GND 0.006804f
C1571 VDD.n1393 GND 0.002697f
C1572 VDD.n1394 GND 0.006148f
C1573 VDD.n1395 GND 0.004948f
C1574 VDD.n1396 GND 0.006148f
C1575 VDD.n1397 GND 0.004948f
C1576 VDD.n1398 GND 0.006148f
C1577 VDD.n1399 GND 0.004948f
C1578 VDD.n1400 GND 0.006148f
C1579 VDD.n1401 GND 0.004948f
C1580 VDD.n1402 GND 0.006148f
C1581 VDD.n1403 GND 0.004874f
C1582 VDD.n1404 GND 0.006148f
C1583 VDD.n1406 GND 0.006148f
C1584 VDD.t3 GND 0.085164f
C1585 VDD.t0 GND 0.430073f
C1586 VDD.n1407 GND 0.075426f
C1587 VDD.t2 GND 0.053191f
C1588 VDD.n1408 GND 0.077435f
C1589 VDD.n1409 GND 0.004948f
C1590 VDD.n1410 GND 0.004948f
C1591 VDD.n1411 GND 0.006148f
C1592 VDD.n1412 GND 0.004948f
C1593 VDD.n1413 GND 0.006148f
C1594 VDD.n1414 GND 0.004948f
C1595 VDD.n1415 GND 0.006148f
C1596 VDD.n1416 GND 0.004948f
C1597 VDD.n1417 GND 0.006148f
C1598 VDD.n1418 GND 0.004181f
C1599 VDD.n1419 GND 0.006148f
C1600 VDD.n1420 GND 0.006148f
C1601 VDD.t9 GND 0.085164f
C1602 VDD.t7 GND 0.430073f
C1603 VDD.n1421 GND 0.075426f
C1604 VDD.t8 GND 0.053191f
C1605 VDD.n1422 GND 0.077435f
C1606 VDD.n1423 GND 0.004948f
C1607 VDD.n1424 GND 0.006148f
C1608 VDD.n1425 GND 0.004948f
C1609 VDD.n1427 GND 0.006148f
C1610 VDD.n1428 GND 0.004948f
C1611 VDD.n1429 GND 0.006148f
C1612 VDD.n1430 GND 0.004948f
C1613 VDD.n1431 GND 0.006148f
C1614 VDD.n1432 GND 0.004948f
C1615 VDD.n1433 GND 0.006148f
C1616 VDD.n1434 GND 0.003488f
C1617 VDD.n1435 GND 0.006148f
C1618 VDD.n1437 GND 0.006148f
C1619 VDD.t16 GND 0.085164f
C1620 VDD.t14 GND 0.430073f
C1621 VDD.n1438 GND 0.075426f
C1622 VDD.t15 GND 0.053191f
C1623 VDD.n1439 GND 0.077435f
C1624 VDD.n1440 GND 0.004948f
C1625 VDD.n1441 GND 0.004948f
C1626 VDD.n1442 GND 0.006148f
C1627 VDD.n1443 GND 0.004948f
C1628 VDD.n1444 GND 0.006148f
C1629 VDD.n1445 GND 0.004948f
C1630 VDD.n1446 GND 0.004107f
C1631 VDD.n1447 GND 0.006148f
C1632 VDD.n1448 GND 0.004948f
C1633 VDD.n1450 GND 0.006148f
C1634 VDD.n1451 GND 0.006148f
C1635 VDD.n1453 GND 0.006148f
C1636 VDD.n1454 GND 0.004948f
C1637 VDD.n1455 GND 0.006148f
C1638 VDD.n1456 GND 0.006148f
C1639 VDD.n1457 GND 0.006148f
C1640 VDD.n1458 GND 0.006148f
C1641 VDD.n1459 GND 0.006148f
C1642 VDD.n1460 GND 0.004948f
C1643 VDD.n1461 GND 0.006148f
C1644 VDD.n1463 GND 0.006148f
C1645 VDD.n1464 GND 0.006148f
C1646 VDD.n1466 GND 0.006148f
C1647 VDD.n1467 GND 0.004775f
C1648 VDD.n1468 GND 0.009278f
C1649 VDD.n1469 GND 0.006148f
C1650 VDD.n1470 GND 0.006148f
C1651 VDD.n1471 GND 0.006148f
C1652 VDD.n1472 GND 0.004948f
C1653 VDD.n1473 GND 0.006148f
C1654 VDD.n1475 GND 0.006148f
C1655 VDD.n1477 GND 0.006148f
C1656 VDD.n1478 GND 0.004948f
C1657 VDD.n1479 GND 0.006148f
C1658 VDD.n1480 GND 0.006148f
C1659 VDD.n1481 GND 0.006148f
C1660 VDD.n1482 GND 0.006148f
C1661 VDD.n1483 GND 0.004948f
C1662 VDD.n1484 GND 0.006148f
C1663 VDD.n1486 GND 0.006148f
C1664 VDD.n1487 GND 0.006148f
C1665 VDD.n1489 GND 0.006148f
C1666 VDD.n1490 GND 0.004948f
C1667 VDD.n1491 GND 0.006148f
C1668 VDD.n1492 GND 0.006148f
C1669 VDD.n1493 GND 0.006148f
C1670 VDD.n1494 GND 0.004082f
C1671 VDD.n1495 GND 0.009278f
C1672 VDD.n1496 GND 0.006148f
C1673 VDD.n1498 GND 0.006148f
C1674 VDD.n1500 GND 0.006148f
C1675 VDD.n1501 GND 0.004948f
C1676 VDD.n1502 GND 0.006148f
C1677 VDD.n1503 GND 0.006148f
C1678 VDD.n1504 GND 0.006148f
C1679 VDD.n1505 GND 0.004948f
C1680 VDD.n1506 GND 0.006148f
C1681 VDD.n1508 GND 0.006148f
C1682 VDD.n1510 GND 0.006148f
C1683 VDD.n1511 GND 0.004948f
C1684 VDD.n1512 GND 0.006148f
C1685 VDD.n1513 GND 0.006148f
C1686 VDD.n1514 GND 0.006148f
C1687 VDD.n1515 GND 0.006148f
C1688 VDD.n1516 GND 0.006148f
C1689 VDD.n1517 GND 0.004948f
C1690 VDD.n1518 GND 0.006148f
C1691 VDD.n1520 GND 0.006148f
C1692 VDD.n1521 GND 0.006148f
C1693 VDD.n1523 GND 0.006148f
C1694 VDD.n1524 GND 0.00339f
C1695 VDD.n1525 GND 0.009278f
C1696 VDD.n1526 GND 0.006148f
C1697 VDD.n1527 GND 0.006148f
C1698 VDD.n1528 GND 0.006148f
C1699 VDD.n1529 GND 0.004948f
C1700 VDD.n1530 GND 0.006148f
C1701 VDD.n1532 GND 0.006148f
C1702 VDD.n1534 GND 0.006148f
C1703 VDD.n1535 GND 0.004948f
C1704 VDD.n1536 GND 0.006148f
C1705 VDD.n1537 GND 0.006148f
C1706 VDD.n1538 GND 0.006148f
C1707 VDD.n1539 GND 0.004948f
C1708 VDD.n1540 GND 0.006148f
C1709 VDD.n1542 GND 0.006148f
C1710 VDD.n1544 GND 0.006148f
C1711 VDD.n1545 GND 0.004948f
C1712 VDD.n1546 GND 0.006148f
C1713 VDD.n1547 GND 0.006148f
C1714 VDD.n1548 GND 0.006148f
C1715 VDD.n1549 GND 0.004948f
C1716 VDD.n1550 GND 0.006148f
C1717 VDD.n1552 GND 0.006148f
C1718 VDD.n1554 GND 0.006148f
C1719 VDD.n1555 GND 0.003093f
C1720 VDD.n1556 GND 0.006148f
C1721 VDD.n1557 GND 0.006148f
C1722 VDD.n1558 GND 0.006148f
C1723 VDD.n1559 GND 0.004948f
C1724 VDD.n1560 GND 0.006148f
C1725 VDD.n1562 GND 0.006148f
C1726 VDD.n1564 GND 0.006148f
C1727 VDD.n1565 GND 0.004948f
C1728 VDD.n1566 GND 0.006148f
C1729 VDD.n1567 GND 0.006148f
C1730 VDD.n1568 GND 0.006148f
C1731 VDD.n1569 GND 0.004948f
C1732 VDD.n1570 GND 0.006148f
C1733 VDD.n1572 GND 0.006148f
C1734 VDD.n1573 GND 0.006148f
C1735 VDD.n1575 GND 0.006148f
C1736 VDD.n1576 GND 0.004948f
C1737 VDD.n1577 GND 0.006148f
C1738 VDD.n1578 GND 0.006148f
C1739 VDD.n1579 GND 0.006148f
C1740 VDD.n1580 GND 0.004478f
C1741 VDD.n1581 GND 0.009278f
C1742 VDD.n1582 GND 0.002944f
C1743 VDD.n1583 GND 0.014117f
C1744 VDD.n1584 GND 0.013671f
C1745 VDD.n1585 GND 0.004107f
C1746 VDD.n1586 GND 0.013671f
C1747 VDD.n1587 GND 0.670043f
C1748 VDD.n1588 GND 0.013671f
C1749 VDD.n1589 GND 0.004107f
C1750 VDD.n1590 GND 0.013671f
C1751 VDD.n1591 GND 0.006148f
C1752 VDD.n1592 GND 0.006148f
C1753 VDD.n1593 GND 0.004948f
C1754 VDD.n1594 GND 0.006148f
C1755 VDD.n1595 GND 0.473529f
C1756 VDD.n1596 GND 0.006148f
C1757 VDD.n1597 GND 0.004948f
C1758 VDD.n1598 GND 0.006148f
C1759 VDD.n1599 GND 0.006148f
C1760 VDD.n1600 GND 0.006148f
C1761 VDD.n1601 GND 0.004948f
C1762 VDD.n1602 GND 0.006148f
C1763 VDD.n1603 GND 0.473529f
C1764 VDD.n1604 GND 0.006148f
C1765 VDD.n1605 GND 0.004948f
C1766 VDD.n1606 GND 0.006148f
C1767 VDD.n1607 GND 0.006148f
C1768 VDD.n1608 GND 0.006148f
C1769 VDD.n1609 GND 0.004948f
C1770 VDD.n1610 GND 0.006148f
C1771 VDD.n1611 GND 0.473529f
C1772 VDD.n1612 GND 0.006148f
C1773 VDD.n1613 GND 0.004948f
C1774 VDD.n1614 GND 0.006148f
C1775 VDD.n1615 GND 0.006148f
C1776 VDD.n1616 GND 0.006148f
C1777 VDD.n1617 GND 0.004948f
C1778 VDD.n1618 GND 0.006148f
C1779 VDD.n1619 GND 0.473529f
C1780 VDD.n1620 GND 0.006148f
C1781 VDD.n1621 GND 0.004948f
C1782 VDD.n1622 GND 0.006148f
C1783 VDD.n1623 GND 0.006148f
C1784 VDD.n1624 GND 0.006148f
C1785 VDD.n1625 GND 0.004948f
C1786 VDD.n1626 GND 0.006148f
C1787 VDD.n1627 GND 0.473529f
C1788 VDD.n1628 GND 0.006148f
C1789 VDD.n1629 GND 0.004948f
C1790 VDD.n1630 GND 0.006148f
C1791 VDD.n1631 GND 0.006148f
C1792 VDD.n1632 GND 0.006148f
C1793 VDD.n1633 GND 0.004948f
C1794 VDD.n1634 GND 0.006148f
C1795 VDD.n1635 GND 0.473529f
C1796 VDD.n1636 GND 0.006148f
C1797 VDD.n1637 GND 0.004948f
C1798 VDD.n1638 GND 0.006148f
C1799 VDD.n1639 GND 0.006148f
C1800 VDD.n1640 GND 0.006148f
C1801 VDD.n1641 GND 0.004948f
C1802 VDD.n1642 GND 0.006148f
C1803 VDD.n1643 GND 0.473529f
C1804 VDD.n1644 GND 0.006148f
C1805 VDD.n1645 GND 0.004948f
C1806 VDD.n1646 GND 0.006148f
C1807 VDD.n1647 GND 0.006148f
C1808 VDD.n1648 GND 0.006148f
C1809 VDD.n1649 GND 0.004948f
C1810 VDD.n1650 GND 0.006148f
C1811 VDD.n1651 GND 0.473529f
C1812 VDD.n1652 GND 0.006148f
C1813 VDD.n1653 GND 0.004948f
C1814 VDD.n1654 GND 0.006148f
C1815 VDD.n1655 GND 0.006148f
C1816 VDD.n1656 GND 0.006148f
C1817 VDD.n1657 GND 0.004948f
C1818 VDD.n1658 GND 0.006148f
C1819 VDD.n1659 GND 0.473529f
C1820 VDD.n1660 GND 0.006148f
C1821 VDD.n1661 GND 0.004948f
C1822 VDD.n1662 GND 0.006148f
C1823 VDD.n1663 GND 0.006148f
C1824 VDD.n1664 GND 0.006148f
C1825 VDD.n1665 GND 0.004948f
C1826 VDD.n1666 GND 0.006148f
C1827 VDD.n1667 GND 0.473529f
C1828 VDD.n1668 GND 0.006148f
C1829 VDD.n1669 GND 0.004948f
C1830 VDD.n1670 GND 0.006148f
C1831 VDD.n1671 GND 0.006148f
C1832 VDD.n1672 GND 0.006127f
C1833 VDD.n1673 GND 0.004948f
C1834 VDD.n1674 GND 0.006148f
C1835 VDD.n1675 GND 0.473529f
C1836 VDD.n1676 GND 0.006148f
C1837 VDD.n1677 GND 0.004948f
C1838 VDD.n1678 GND 0.006148f
C1839 VDD.n1679 GND 0.006148f
C1840 VDD.n1680 GND 0.006148f
C1841 VDD.n1681 GND 0.004948f
C1842 VDD.n1682 GND 0.006148f
C1843 VDD.n1683 GND 0.473529f
C1844 VDD.n1684 GND 0.006148f
C1845 VDD.n1685 GND 0.004948f
C1846 VDD.n1686 GND 0.006127f
C1847 VDD.n1687 GND 0.006148f
C1848 VDD.n1688 GND 0.006148f
C1849 VDD.n1689 GND 0.004948f
C1850 VDD.n1690 GND 0.006148f
C1851 VDD.n1691 GND 0.473529f
C1852 VDD.n1692 GND 0.006148f
C1853 VDD.n1693 GND 0.004948f
C1854 VDD.n1694 GND 0.006148f
C1855 VDD.n1695 GND 0.006148f
C1856 VDD.n1696 GND 0.006148f
C1857 VDD.n1697 GND 0.004948f
C1858 VDD.n1698 GND 0.006148f
C1859 VDD.n1699 GND 0.473529f
C1860 VDD.n1700 GND 0.006148f
C1861 VDD.n1701 GND 0.004948f
C1862 VDD.n1702 GND 0.006148f
C1863 VDD.n1703 GND 0.006148f
C1864 VDD.n1704 GND 0.006148f
C1865 VDD.n1705 GND 0.004948f
C1866 VDD.n1706 GND 0.006148f
C1867 VDD.n1707 GND 0.473529f
C1868 VDD.n1708 GND 0.006148f
C1869 VDD.n1709 GND 0.004948f
C1870 VDD.n1710 GND 0.006148f
C1871 VDD.n1711 GND 0.006148f
C1872 VDD.n1712 GND 0.006148f
C1873 VDD.n1713 GND 0.004948f
C1874 VDD.n1714 GND 0.006148f
C1875 VDD.n1715 GND 0.473529f
C1876 VDD.n1716 GND 0.006148f
C1877 VDD.n1717 GND 0.004948f
C1878 VDD.n1718 GND 0.006148f
C1879 VDD.n1719 GND 0.006148f
C1880 VDD.n1720 GND 0.006148f
C1881 VDD.n1721 GND 0.004948f
C1882 VDD.n1722 GND 0.006148f
C1883 VDD.n1723 GND 0.473529f
C1884 VDD.n1724 GND 0.006148f
C1885 VDD.n1725 GND 0.004948f
C1886 VDD.n1726 GND 0.006148f
C1887 VDD.n1727 GND 0.006148f
C1888 VDD.n1728 GND 0.006148f
C1889 VDD.n1729 GND 0.004948f
C1890 VDD.n1730 GND 0.006148f
C1891 VDD.n1731 GND 0.473529f
C1892 VDD.n1732 GND 0.006148f
C1893 VDD.n1733 GND 0.004948f
C1894 VDD.n1734 GND 0.006148f
C1895 VDD.n1735 GND 0.006148f
C1896 VDD.n1736 GND 0.006148f
C1897 VDD.n1737 GND 0.004948f
C1898 VDD.n1738 GND 0.006148f
C1899 VDD.n1739 GND 0.473529f
C1900 VDD.n1740 GND 0.006148f
C1901 VDD.n1741 GND 0.004948f
C1902 VDD.n1742 GND 0.006148f
C1903 VDD.n1743 GND 0.006148f
C1904 VDD.n1744 GND 0.006148f
C1905 VDD.n1745 GND 0.004948f
C1906 VDD.n1746 GND 0.006148f
C1907 VDD.n1747 GND 0.473529f
C1908 VDD.n1748 GND 0.006148f
C1909 VDD.n1749 GND 0.004948f
C1910 VDD.n1750 GND 0.006148f
C1911 VDD.n1751 GND 0.006148f
C1912 VDD.n1752 GND 0.006148f
C1913 VDD.n1753 GND 0.004948f
C1914 VDD.n1754 GND 0.006148f
C1915 VDD.n1755 GND 0.473529f
C1916 VDD.n1756 GND 0.006148f
C1917 VDD.n1757 GND 0.004948f
C1918 VDD.n1758 GND 0.006148f
C1919 VDD.n1759 GND 0.006148f
C1920 VDD.n1760 GND 0.013671f
C1921 VDD.n1761 GND 0.006148f
C1922 VDD.n1762 GND 0.006148f
C1923 VDD.n1763 GND 0.004948f
C1924 VDD.n1764 GND 0.006148f
C1925 VDD.n1765 GND 0.473529f
C1926 VDD.n1766 GND 0.006148f
C1927 VDD.n1767 GND 0.004948f
C1928 VDD.n1768 GND 0.006148f
C1929 VDD.n1769 GND 0.006148f
C1930 VDD.n1770 GND 0.006148f
C1931 VDD.n1772 GND 0.006148f
C1932 VDD.n1773 GND 0.006148f
C1933 VDD.n1774 GND 0.004948f
C1934 VDD.n1775 GND 0.004948f
C1935 VDD.n1776 GND 0.006148f
C1936 VDD.n1777 GND 0.006148f
C1937 VDD.n1778 GND 0.006148f
C1938 VDD.n1779 GND 0.006148f
C1939 VDD.n1780 GND 0.006148f
C1940 VDD.n1781 GND 0.006148f
C1941 VDD.n1782 GND 0.006148f
C1942 VDD.n1783 GND 0.004775f
C1943 VDD.n1786 GND 0.006148f
C1944 VDD.n1787 GND 0.006148f
C1945 VDD.n1788 GND 0.004948f
C1946 VDD.n1789 GND 0.004948f
C1947 VDD.n1790 GND 0.004948f
C1948 VDD.n1791 GND 0.006148f
C1949 VDD.n1793 GND 0.006148f
C1950 VDD.n1794 GND 0.006148f
C1951 VDD.n1796 GND 0.006148f
C1952 VDD.n1797 GND 0.004948f
C1953 VDD.n1798 GND 0.004948f
C1954 VDD.n1799 GND 0.004107f
C1955 VDD.n1800 GND 0.014117f
C1956 VDD.n1801 GND 0.013671f
C1957 VDD.n1802 GND 0.004107f
C1958 VDD.n1803 GND 0.013671f
C1959 VDD.n1804 GND 0.670043f
C1960 VDD.n1805 GND 0.013671f
C1961 VDD.n1806 GND 0.014117f
C1962 VDD.n1808 GND 0.006148f
C1963 VDD.n1809 GND 0.009278f
C1964 VDD.n1810 GND 0.006148f
C1965 VDD.n1811 GND 0.006148f
C1966 VDD.n1812 GND 0.006148f
C1967 VDD.n1813 GND 0.004948f
C1968 VDD.n1814 GND 0.004948f
C1969 VDD.n1815 GND 0.004948f
C1970 VDD.n1816 GND 0.006148f
C1971 VDD.n1817 GND 0.006148f
C1972 VDD.n1818 GND 0.006148f
C1973 VDD.n1819 GND 0.004948f
C1974 VDD.n1820 GND 0.004948f
C1975 VDD.n1821 GND 0.004948f
C1976 VDD.n1822 GND 0.003935f
C1977 VDD.n1823 GND 1.04933f
C1978 VDD.n1825 GND 0.003093f
C1979 VDD.n1826 GND 0.006148f
C1980 VDD.n1828 GND 0.006148f
C1981 VDD.n1829 GND 0.006148f
C1982 VDD.n1830 GND 0.004948f
C1983 VDD.n1831 GND 0.004948f
C1984 VDD.n1832 GND 0.004948f
C1985 VDD.n1833 GND 0.006148f
C1986 VDD.n1835 GND 0.006148f
C1987 VDD.n1836 GND 0.006148f
C1988 VDD.n1837 GND 0.004948f
C1989 VDD.n1838 GND 0.004948f
C1990 VDD.n1839 GND 0.004948f
C1991 VDD.n1840 GND 0.006148f
C1992 VDD.n1842 GND 0.006148f
C1993 VDD.n1843 GND 0.006148f
C1994 VDD.n1844 GND 0.004948f
C1995 VDD.n1845 GND 0.006148f
C1996 VDD.n1846 GND 0.006148f
C1997 VDD.n1847 GND 0.006148f
C1998 VDD.n1848 GND 0.009278f
C1999 VDD.n1849 GND 0.006148f
C2000 VDD.n1851 GND 0.006148f
C2001 VDD.n1852 GND 0.006148f
C2002 VDD.n1853 GND 0.004948f
C2003 VDD.n1854 GND 0.004948f
C2004 VDD.n1855 GND 0.004948f
C2005 VDD.n1856 GND 0.006148f
C2006 VDD.n1858 GND 0.006148f
C2007 VDD.n1859 GND 0.006148f
C2008 VDD.n1860 GND 0.004948f
C2009 VDD.n1861 GND 0.004948f
C2010 VDD.n1862 GND 0.004948f
C2011 VDD.n1863 GND 0.006148f
C2012 VDD.n1865 GND 0.006148f
C2013 VDD.n1866 GND 0.006148f
C2014 VDD.n1867 GND 0.004948f
C2015 VDD.n1868 GND 0.006148f
C2016 VDD.n1869 GND 0.006148f
C2017 VDD.n1870 GND 0.006148f
C2018 VDD.n1871 GND 0.009278f
C2019 VDD.n1872 GND 0.006148f
C2020 VDD.n1874 GND 0.006148f
C2021 VDD.n1875 GND 0.006148f
C2022 VDD.n1876 GND 0.004948f
C2023 VDD.n1877 GND 0.004948f
C2024 VDD.n1878 GND 0.004948f
C2025 VDD.n1879 GND 0.006148f
C2026 VDD.n1881 GND 0.006148f
C2027 VDD.n1882 GND 0.006148f
C2028 VDD.n1883 GND 0.004948f
C2029 VDD.n1884 GND 0.004948f
C2030 VDD.n1885 GND 0.004948f
C2031 VDD.n1886 GND 0.006148f
C2032 VDD.n1888 GND 0.006148f
C2033 VDD.n1889 GND 0.006148f
C2034 VDD.n1891 GND 0.006148f
C2035 VDD.n1892 GND 0.003488f
C2036 VDD.n1894 GND 1.04933f
C2037 VDD.n1895 GND 0.063036f
C2038 VDD.n1896 GND 0.003135f
C2039 VDD.n1897 GND 0.00418f
C2040 VDD.n1898 GND 0.00418f
C2041 VDD.n1899 GND 0.00418f
C2042 VDD.n1901 GND 0.00418f
C2043 VDD.n1902 GND 0.00418f
C2044 VDD.n1903 GND 0.00418f
C2045 VDD.n1904 GND 0.00418f
C2046 VDD.n1905 GND 0.00418f
C2047 VDD.n1907 GND 0.00418f
C2048 VDD.n1909 GND 0.00418f
C2049 VDD.n1910 GND 0.00418f
C2050 VDD.n1911 GND 0.00418f
C2051 VDD.n1912 GND 0.00418f
C2052 VDD.n1913 GND 0.00418f
C2053 VDD.n1915 GND 0.00418f
C2054 VDD.n1917 GND 0.00418f
C2055 VDD.n1918 GND 0.003135f
C2056 VDD.n1919 GND 0.00418f
C2057 VDD.n1920 GND 0.00418f
C2058 VDD.n1921 GND 0.00418f
C2059 VDD.n1923 GND 0.00418f
C2060 VDD.n1925 GND 0.00418f
C2061 VDD.n1926 GND 0.003105f
C2062 VDD.n1927 GND 0.005158f
C2063 VDD.n1928 GND 0.003166f
C2064 VDD.n1929 GND 0.00418f
C2065 VDD.n1930 GND 0.00418f
C2066 VDD.n1932 GND 0.00418f
C2067 VDD.n1933 GND 0.009514f
C2068 VDD.n1934 GND 0.009514f
C2069 VDD.n1935 GND 0.008807f
C2070 VDD.n1936 GND 0.00418f
C2071 VDD.n1937 GND 0.00418f
C2072 VDD.n1938 GND 0.00418f
C2073 VDD.n1939 GND 0.00418f
C2074 VDD.n1940 GND 0.00418f
C2075 VDD.n1941 GND 0.00418f
C2076 VDD.n1942 GND 0.00418f
C2077 VDD.n1943 GND 0.00418f
C2078 VDD.n1944 GND 0.00418f
C2079 VDD.n1945 GND 0.00418f
C2080 VDD.n1946 GND 0.00418f
C2081 VDD.n1947 GND 0.00418f
C2082 VDD.n1948 GND 0.00418f
C2083 VDD.n1949 GND 0.00418f
C2084 VDD.n1950 GND 0.00418f
C2085 VDD.n1951 GND 0.00418f
C2086 VDD.n1952 GND 0.00418f
C2087 VDD.n1953 GND 0.00418f
C2088 VDD.n1954 GND 0.00418f
C2089 VDD.n1955 GND 0.00418f
C2090 VDD.n1956 GND 0.00418f
C2091 VDD.n1957 GND 0.00418f
C2092 VDD.n1958 GND 0.00418f
C2093 VDD.n1959 GND 0.00418f
C2094 VDD.n1960 GND 0.00418f
C2095 VDD.n1961 GND 0.00418f
C2096 VDD.n1962 GND 0.00418f
C2097 VDD.n1963 GND 0.00418f
C2098 VDD.n1964 GND 0.00418f
C2099 VDD.n1965 GND 0.00418f
C2100 VDD.n1966 GND 0.00418f
C2101 VDD.n1967 GND 0.00418f
C2102 VDD.n1968 GND 0.00418f
C2103 VDD.n1969 GND 0.00418f
C2104 VDD.n1970 GND 0.00418f
C2105 VDD.n1971 GND 0.00418f
C2106 VDD.n1972 GND 0.00418f
C2107 VDD.n1973 GND 0.00418f
C2108 VDD.n1974 GND 0.00418f
C2109 VDD.n1975 GND 0.00418f
C2110 VDD.n1976 GND 0.00418f
C2111 VDD.n1977 GND 0.00418f
C2112 VDD.n1978 GND 0.00418f
C2113 VDD.n1979 GND 0.00418f
C2114 VDD.n1980 GND 0.00418f
C2115 VDD.n1981 GND 0.00418f
C2116 VDD.n1982 GND 0.00418f
C2117 VDD.n1983 GND 0.00418f
C2118 VDD.n1984 GND 0.00418f
C2119 VDD.n1985 GND 0.00418f
C2120 VDD.n1986 GND 0.00418f
C2121 VDD.n1987 GND 0.00418f
C2122 VDD.n1988 GND 0.00418f
C2123 VDD.n1989 GND 0.00418f
C2124 VDD.n1990 GND 0.00418f
C2125 VDD.n1991 GND 0.00418f
C2126 VDD.n1992 GND 0.00418f
C2127 VDD.n1993 GND 0.00418f
C2128 VDD.n1994 GND 0.00418f
C2129 VDD.n1995 GND 0.00418f
C2130 VDD.n1996 GND 0.00418f
C2131 VDD.n1997 GND 0.00418f
C2132 VDD.n1998 GND 0.00418f
C2133 VDD.n1999 GND 0.00418f
C2134 VDD.n2000 GND 0.00418f
C2135 VDD.n2001 GND 0.00418f
C2136 VDD.n2002 GND 0.00418f
C2137 VDD.n2003 GND 0.00418f
C2138 VDD.n2004 GND 0.00418f
C2139 VDD.n2005 GND 0.00418f
C2140 VDD.n2006 GND 0.00418f
C2141 VDD.n2007 GND 0.00418f
C2142 VDD.n2008 GND 0.00418f
C2143 VDD.n2009 GND 0.00418f
C2144 VDD.n2010 GND 0.00418f
C2145 VDD.n2011 GND 0.00418f
C2146 VDD.n2012 GND 0.00418f
C2147 VDD.n2013 GND 0.00418f
C2148 VDD.n2014 GND 0.00418f
C2149 VDD.n2015 GND 0.00418f
C2150 VDD.n2016 GND 0.00418f
C2151 VDD.n2017 GND 0.00418f
C2152 VDD.n2018 GND 0.00418f
C2153 VDD.n2019 GND 0.00418f
C2154 VDD.n2020 GND 0.00418f
C2155 VDD.n2021 GND 0.00418f
C2156 VDD.n2022 GND 0.00418f
C2157 VDD.n2023 GND 0.00418f
C2158 VDD.n2024 GND 0.00418f
C2159 VDD.n2025 GND 0.00418f
C2160 VDD.n2026 GND 0.00418f
C2161 VDD.n2027 GND 0.00418f
C2162 VDD.n2028 GND 0.00418f
C2163 VDD.n2029 GND 0.00418f
C2164 VDD.n2030 GND 0.00418f
C2165 VDD.n2031 GND 0.00418f
C2166 VDD.n2032 GND 0.00418f
C2167 VDD.n2033 GND 0.00418f
C2168 VDD.n2034 GND 0.00418f
C2169 VDD.n2035 GND 0.00418f
C2170 VDD.n2036 GND 0.00418f
C2171 VDD.n2037 GND 0.00418f
C2172 VDD.n2038 GND 0.00418f
C2173 VDD.n2039 GND 0.00418f
C2174 VDD.n2040 GND 0.00418f
C2175 VDD.n2041 GND 0.00418f
C2176 VDD.n2042 GND 0.00418f
C2177 VDD.n2043 GND 0.00418f
C2178 VDD.n2044 GND 0.00418f
C2179 VDD.n2045 GND 0.00418f
C2180 VDD.n2046 GND 0.00418f
C2181 VDD.n2047 GND 0.00418f
C2182 VDD.n2048 GND 0.00418f
C2183 VDD.n2049 GND 0.00418f
C2184 VDD.n2050 GND 0.00418f
C2185 VDD.n2051 GND 0.00418f
C2186 VDD.n2052 GND 0.00418f
C2187 VDD.n2053 GND 0.00418f
C2188 VDD.n2054 GND 0.00418f
C2189 VDD.n2055 GND 0.00418f
C2190 VDD.n2056 GND 0.00418f
C2191 VDD.n2057 GND 0.00418f
C2192 VDD.n2058 GND 0.00418f
C2193 VDD.n2059 GND 0.00418f
C2194 VDD.n2060 GND 0.00418f
C2195 VDD.n2061 GND 0.00418f
C2196 VDD.n2062 GND 0.00418f
C2197 VDD.n2063 GND 0.00418f
C2198 VDD.n2064 GND 0.00418f
C2199 VDD.n2065 GND 0.00418f
C2200 VDD.n2066 GND 0.00418f
C2201 VDD.n2067 GND 0.00418f
C2202 VDD.n2068 GND 0.00418f
C2203 VDD.n2069 GND 0.00418f
C2204 VDD.n2070 GND 0.00418f
C2205 VDD.n2071 GND 0.00418f
C2206 VDD.n2072 GND 0.00418f
C2207 VDD.n2073 GND 0.00418f
C2208 VDD.n2074 GND 0.00418f
C2209 VDD.n2075 GND 0.00418f
C2210 VDD.n2076 GND 0.00418f
C2211 VDD.n2077 GND 0.00418f
C2212 VDD.n2078 GND 0.00418f
C2213 VDD.n2079 GND 0.00418f
C2214 VDD.n2080 GND 0.00418f
C2215 VDD.n2081 GND 0.00418f
C2216 VDD.n2082 GND 0.00418f
C2217 VDD.n2083 GND 0.00418f
C2218 VDD.n2084 GND 0.00418f
C2219 VDD.n2085 GND 0.00418f
C2220 VDD.n2086 GND 0.00418f
C2221 VDD.n2087 GND 0.00418f
C2222 VDD.n2088 GND 0.00418f
C2223 VDD.n2089 GND 0.00418f
C2224 VDD.n2090 GND 0.00418f
C2225 VDD.n2091 GND 0.00418f
C2226 VDD.n2092 GND 0.00418f
C2227 VDD.n2093 GND 0.00418f
C2228 VDD.n2094 GND 0.00418f
C2229 VDD.n2095 GND 0.00418f
C2230 VDD.n2096 GND 0.00418f
C2231 VDD.n2097 GND 0.00418f
C2232 VDD.n2098 GND 0.00418f
C2233 VDD.n2099 GND 0.00418f
C2234 VDD.n2100 GND 0.00418f
C2235 VDD.n2101 GND 0.00418f
C2236 VDD.n2102 GND 0.00418f
C2237 VDD.n2103 GND 0.00418f
C2238 VDD.n2104 GND 0.00418f
C2239 VDD.n2105 GND 0.00418f
C2240 VDD.n2106 GND 0.00418f
C2241 VDD.n2107 GND 0.00418f
C2242 VDD.n2108 GND 0.00418f
C2243 VDD.n2109 GND 0.00418f
C2244 VDD.n2110 GND 0.00418f
C2245 VDD.n2111 GND 0.00418f
C2246 VDD.n2112 GND 0.00418f
C2247 VDD.n2113 GND 0.00418f
C2248 VDD.n2114 GND 0.00418f
C2249 VDD.n2115 GND 0.00418f
C2250 VDD.n2116 GND 0.00418f
C2251 VDD.n2117 GND 0.00418f
C2252 VDD.n2118 GND 0.00418f
C2253 VDD.n2119 GND 0.00418f
C2254 VDD.n2120 GND 0.00418f
C2255 VDD.n2121 GND 0.00418f
C2256 VDD.n2122 GND 0.00418f
C2257 VDD.n2123 GND 0.00418f
C2258 VDD.n2124 GND 0.00418f
C2259 VDD.n2125 GND 0.00418f
C2260 VDD.n2126 GND 0.00418f
C2261 VDD.n2127 GND 0.00418f
C2262 VDD.n2128 GND 0.00418f
C2263 VDD.n2129 GND 0.00418f
C2264 VDD.n2130 GND 0.00418f
C2265 VDD.n2131 GND 0.00418f
C2266 VDD.n2132 GND 0.00418f
C2267 VDD.n2133 GND 0.00418f
C2268 VDD.n2134 GND 0.00418f
C2269 VDD.n2135 GND 0.00418f
C2270 VDD.n2136 GND 0.00418f
C2271 VDD.n2137 GND 0.00418f
C2272 VDD.n2138 GND 0.00418f
C2273 VDD.n2139 GND 0.00418f
C2274 VDD.n2140 GND 0.00418f
C2275 VDD.n2141 GND 0.00418f
C2276 VDD.n2142 GND 0.00418f
C2277 VDD.n2143 GND 0.00418f
C2278 VDD.n2144 GND 0.00418f
C2279 VDD.n2145 GND 0.00418f
C2280 VDD.n2146 GND 0.00418f
C2281 VDD.n2147 GND 0.269911f
C2282 VDD.n2148 GND 0.00418f
C2283 VDD.n2149 GND 0.00418f
C2284 VDD.n2150 GND 0.00418f
C2285 VDD.n2151 GND 0.00418f
C2286 VDD.n2152 GND 0.00418f
C2287 VDD.n2153 GND 0.00418f
C2288 VDD.n2154 GND 0.00418f
C2289 VDD.n2155 GND 0.00418f
C2290 VDD.n2156 GND 0.00418f
C2291 VDD.n2157 GND 0.00418f
C2292 VDD.n2158 GND 0.00418f
C2293 VDD.n2159 GND 0.00418f
C2294 VDD.n2160 GND 0.00418f
C2295 VDD.n2161 GND 0.00418f
C2296 VDD.n2162 GND 0.00418f
C2297 VDD.n2163 GND 0.00418f
C2298 VDD.n2164 GND 0.00418f
C2299 VDD.n2165 GND 0.00418f
C2300 VDD.n2166 GND 0.00418f
C2301 VDD.n2167 GND 0.00418f
C2302 VDD.n2168 GND 0.00418f
C2303 VDD.n2169 GND 0.00418f
C2304 VDD.n2170 GND 0.00418f
C2305 VDD.n2171 GND 0.00418f
C2306 VDD.n2172 GND 0.00418f
C2307 VDD.n2173 GND 0.00418f
C2308 VDD.n2174 GND 0.00418f
C2309 VDD.n2175 GND 0.00418f
C2310 VDD.n2176 GND 0.00418f
C2311 VDD.n2177 GND 0.00418f
C2312 VDD.n2178 GND 0.00418f
C2313 VDD.n2179 GND 0.00418f
C2314 VDD.n2180 GND 0.00418f
C2315 VDD.n2181 GND 0.00418f
C2316 VDD.n2182 GND 0.00418f
C2317 VDD.n2183 GND 0.00418f
C2318 VDD.n2184 GND 0.00418f
C2319 VDD.n2185 GND 0.00418f
C2320 VDD.n2186 GND 0.00418f
C2321 VDD.n2187 GND 0.00418f
C2322 VDD.n2188 GND 0.00418f
C2323 VDD.n2189 GND 0.00418f
C2324 VDD.n2190 GND 0.00418f
C2325 VDD.n2191 GND 0.00418f
C2326 VDD.n2192 GND 0.00418f
C2327 VDD.n2193 GND 0.00418f
C2328 VDD.n2194 GND 0.00418f
C2329 VDD.n2195 GND 0.00418f
C2330 VDD.n2196 GND 0.00418f
C2331 VDD.n2197 GND 0.00418f
C2332 VDD.n2198 GND 0.00418f
C2333 VDD.n2199 GND 0.00418f
C2334 VDD.n2200 GND 0.00418f
C2335 VDD.n2201 GND 0.00418f
C2336 VDD.n2202 GND 0.00418f
C2337 VDD.n2203 GND 0.00418f
C2338 VDD.n2204 GND 0.00418f
C2339 VDD.n2205 GND 0.00418f
C2340 VDD.n2206 GND 0.00418f
C2341 VDD.n2207 GND 0.00418f
C2342 VDD.n2208 GND 0.00418f
C2343 VDD.n2209 GND 0.00418f
C2344 VDD.n2210 GND 0.00418f
C2345 VDD.n2211 GND 0.00418f
C2346 VDD.n2212 GND 0.00418f
C2347 VDD.n2213 GND 0.00418f
C2348 VDD.n2214 GND 0.00418f
C2349 VDD.n2215 GND 0.00418f
C2350 VDD.n2216 GND 0.00418f
C2351 VDD.n2217 GND 0.00418f
C2352 VDD.n2218 GND 0.00418f
C2353 VDD.n2219 GND 0.00418f
C2354 VDD.n2220 GND 0.00418f
C2355 VDD.n2221 GND 0.00418f
C2356 VDD.n2222 GND 0.00418f
C2357 VDD.n2223 GND 0.00418f
C2358 VDD.n2224 GND 0.00418f
C2359 VDD.n2225 GND 0.00418f
C2360 VDD.n2226 GND 0.00418f
C2361 VDD.n2227 GND 0.00418f
C2362 VDD.n2228 GND 0.00418f
C2363 VDD.n2229 GND 0.00418f
C2364 VDD.n2230 GND 0.00418f
C2365 VDD.n2231 GND 0.00418f
C2366 VDD.n2232 GND 0.00418f
C2367 VDD.n2233 GND 0.00418f
C2368 VDD.n2234 GND 0.00418f
C2369 VDD.n2235 GND 0.00418f
C2370 VDD.n2236 GND 0.00418f
C2371 VDD.n2237 GND 0.00418f
C2372 VDD.n2238 GND 0.00418f
C2373 VDD.n2239 GND 0.00418f
C2374 VDD.n2240 GND 0.00418f
C2375 VDD.n2241 GND 0.00418f
C2376 VDD.n2242 GND 0.00418f
C2377 VDD.n2243 GND 0.00418f
C2378 VDD.n2244 GND 0.00418f
C2379 VDD.n2245 GND 0.00418f
C2380 VDD.n2246 GND 0.00418f
C2381 VDD.n2247 GND 0.00418f
C2382 VDD.n2248 GND 0.00418f
C2383 VDD.n2249 GND 0.00418f
C2384 VDD.n2250 GND 0.00418f
C2385 VDD.n2251 GND 0.00418f
C2386 VDD.n2252 GND 0.00418f
C2387 VDD.n2253 GND 0.00418f
C2388 VDD.n2254 GND 0.00418f
C2389 VDD.n2255 GND 0.00418f
C2390 VDD.n2256 GND 0.00418f
C2391 VDD.n2257 GND 0.00418f
C2392 VDD.n2258 GND 0.00418f
C2393 VDD.n2259 GND 0.00418f
C2394 VDD.n2260 GND 0.00418f
C2395 VDD.n2261 GND 0.00418f
C2396 VDD.n2262 GND 0.00418f
C2397 VDD.n2263 GND 0.00418f
C2398 VDD.n2264 GND 0.00418f
C2399 VDD.n2265 GND 0.00418f
C2400 VDD.n2266 GND 0.00418f
C2401 VDD.n2267 GND 0.00418f
C2402 VDD.n2268 GND 0.00418f
C2403 VDD.n2269 GND 0.00418f
C2404 VDD.n2270 GND 0.00418f
C2405 VDD.n2271 GND 0.00418f
C2406 VDD.n2272 GND 0.00418f
C2407 VDD.n2273 GND 0.00418f
C2408 VDD.n2274 GND 0.00418f
C2409 VDD.n2275 GND 0.00418f
C2410 VDD.n2276 GND 0.00418f
C2411 VDD.n2277 GND 0.00418f
C2412 VDD.n2278 GND 0.00418f
C2413 VDD.n2279 GND 0.00418f
C2414 VDD.n2280 GND 0.00418f
C2415 VDD.n2281 GND 0.00418f
C2416 VDD.n2282 GND 0.00418f
C2417 VDD.n2283 GND 0.00418f
C2418 VDD.n2284 GND 0.00418f
C2419 VDD.n2285 GND 0.00418f
C2420 VDD.n2286 GND 0.00418f
C2421 VDD.n2287 GND 0.00418f
C2422 VDD.n2288 GND 0.00418f
C2423 VDD.n2289 GND 0.00418f
C2424 VDD.n2290 GND 0.00418f
C2425 VDD.n2291 GND 0.00418f
C2426 VDD.n2292 GND 0.00418f
C2427 VDD.n2293 GND 0.00418f
C2428 VDD.n2294 GND 0.00418f
C2429 VDD.n2295 GND 0.00418f
C2430 VDD.n2296 GND 0.00418f
C2431 VDD.n2297 GND 0.00418f
C2432 VDD.n2298 GND 0.00418f
C2433 VDD.n2299 GND 0.00418f
C2434 VDD.n2300 GND 0.00418f
C2435 VDD.n2301 GND 0.00418f
C2436 VDD.n2302 GND 0.00418f
C2437 VDD.n2303 GND 0.00418f
C2438 VDD.n2304 GND 0.00418f
C2439 VDD.n2305 GND 0.00418f
C2440 VDD.n2306 GND 0.00418f
C2441 VDD.n2307 GND 0.00418f
C2442 VDD.n2308 GND 0.00418f
C2443 VDD.n2309 GND 0.00418f
C2444 VDD.n2310 GND 0.00418f
C2445 VDD.n2311 GND 0.00418f
C2446 VDD.n2312 GND 0.00418f
C2447 VDD.n2313 GND 0.00418f
C2448 VDD.n2314 GND 0.00418f
C2449 VDD.n2315 GND 0.00418f
C2450 VDD.n2316 GND 0.00418f
C2451 VDD.n2317 GND 0.00418f
C2452 VDD.n2318 GND 0.00418f
C2453 VDD.n2319 GND 0.00418f
C2454 VDD.n2320 GND 0.00418f
C2455 VDD.n2321 GND 0.00418f
C2456 VDD.n2322 GND 0.00418f
C2457 VDD.n2323 GND 0.00418f
C2458 VDD.n2324 GND 0.00418f
C2459 VDD.n2325 GND 0.00418f
C2460 VDD.n2326 GND 0.00418f
C2461 VDD.n2327 GND 0.00418f
C2462 VDD.n2328 GND 0.00418f
C2463 VDD.n2329 GND 0.00418f
C2464 VDD.n2330 GND 0.00418f
C2465 VDD.n2331 GND 0.00418f
C2466 VDD.n2332 GND 0.00418f
C2467 VDD.n2333 GND 0.00418f
C2468 VDD.n2334 GND 0.00418f
C2469 VDD.n2335 GND 0.00418f
C2470 VDD.n2336 GND 0.00418f
C2471 VDD.n2337 GND 0.00418f
C2472 VDD.n2338 GND 0.00418f
C2473 VDD.n2339 GND 0.00418f
C2474 VDD.n2340 GND 0.00418f
C2475 VDD.n2341 GND 0.00418f
C2476 VDD.n2342 GND 0.00418f
C2477 VDD.n2343 GND 0.00418f
C2478 VDD.n2344 GND 0.00418f
C2479 VDD.n2345 GND 0.00418f
C2480 VDD.n2346 GND 0.00418f
C2481 VDD.n2347 GND 0.00418f
C2482 VDD.n2348 GND 0.008807f
C2483 VDD.n2349 GND 0.009514f
C2484 VDD.n2350 GND 0.00418f
C2485 VDD.n2351 GND 0.00418f
C2486 VDD.n2353 GND 0.00418f
C2487 VDD.n2355 GND 0.00418f
C2488 VDD.n2356 GND 0.003166f
C2489 VDD.n2357 GND 0.005158f
C2490 VDD.n2358 GND 0.003105f
C2491 VDD.n2359 GND 0.00418f
C2492 VDD.n2360 GND 0.00418f
C2493 VDD.n2362 GND 0.00418f
C2494 VDD.n2363 GND 0.00418f
C2495 VDD.n2364 GND 0.00418f
C2496 VDD.n2365 GND 0.003135f
C2497 VDD.n2366 GND 0.00418f
C2498 VDD.n2368 GND 0.00418f
C2499 VDD.n2369 GND 0.003135f
C2500 VDD.n2370 GND 0.00418f
C2501 VDD.n2371 GND 0.00418f
C2502 VDD.n2372 GND 0.00418f
C2503 VDD.n2374 GND 0.00418f
C2504 VDD.n2375 GND 0.00418f
C2505 VDD.n2376 GND 0.00418f
C2506 VDD.n2377 GND 0.00418f
C2507 VDD.n2378 GND 0.00418f
C2508 VDD.n2379 GND 0.00418f
C2509 VDD.n2381 GND 0.00418f
C2510 VDD.n2382 GND 0.00418f
C2511 VDD.n2383 GND 0.009514f
C2512 VDD.n2384 GND 0.008807f
C2513 VDD.n2385 GND 0.008807f
C2514 VDD.n2386 GND 0.447485f
C2515 VDD.n2387 GND 0.008807f
C2516 VDD.n2388 GND 0.008807f
C2517 VDD.n2389 GND 0.00418f
C2518 VDD.n2390 GND 0.00418f
C2519 VDD.n2391 GND 0.00418f
C2520 VDD.n2392 GND 0.322f
C2521 VDD.n2393 GND 0.00418f
C2522 VDD.n2394 GND 0.00418f
C2523 VDD.n2395 GND 0.00418f
C2524 VDD.n2396 GND 0.00418f
C2525 VDD.n2397 GND 0.00418f
C2526 VDD.n2398 GND 0.322f
C2527 VDD.n2399 GND 0.00418f
C2528 VDD.n2400 GND 0.00418f
C2529 VDD.n2401 GND 0.00418f
C2530 VDD.n2402 GND 0.00418f
C2531 VDD.n2403 GND 0.00418f
C2532 VDD.n2404 GND 0.322f
C2533 VDD.n2405 GND 0.00418f
C2534 VDD.n2406 GND 0.00418f
C2535 VDD.n2407 GND 0.00418f
C2536 VDD.n2408 GND 0.00418f
C2537 VDD.n2409 GND 0.00418f
C2538 VDD.n2410 GND 0.265176f
C2539 VDD.n2411 GND 0.00418f
C2540 VDD.n2412 GND 0.00418f
C2541 VDD.n2413 GND 0.00418f
C2542 VDD.n2414 GND 0.00418f
C2543 VDD.n2415 GND 0.00418f
C2544 VDD.n2416 GND 0.322f
C2545 VDD.n2417 GND 0.00418f
C2546 VDD.n2418 GND 0.00418f
C2547 VDD.n2419 GND 0.00418f
C2548 VDD.n2420 GND 0.00418f
C2549 VDD.n2421 GND 0.00418f
C2550 VDD.n2422 GND 0.298323f
C2551 VDD.n2423 GND 0.00418f
C2552 VDD.n2424 GND 0.00418f
C2553 VDD.n2425 GND 0.00418f
C2554 VDD.n2426 GND 0.00418f
C2555 VDD.n2427 GND 0.00418f
C2556 VDD.n2428 GND 0.322f
C2557 VDD.n2429 GND 0.00418f
C2558 VDD.n2430 GND 0.00418f
C2559 VDD.n2431 GND 0.00418f
C2560 VDD.n2432 GND 0.00418f
C2561 VDD.n2433 GND 0.00418f
C2562 VDD.n2434 GND 0.322f
C2563 VDD.n2435 GND 0.00418f
C2564 VDD.n2436 GND 0.00418f
C2565 VDD.n2437 GND 0.00418f
C2566 VDD.n2438 GND 0.00418f
C2567 VDD.n2439 GND 0.00418f
C2568 VDD.n2440 GND 0.322f
C2569 VDD.n2441 GND 0.00418f
C2570 VDD.n2442 GND 0.00418f
C2571 VDD.n2443 GND 0.00418f
C2572 VDD.n2444 GND 0.00418f
C2573 VDD.n2445 GND 0.00418f
C2574 VDD.n2446 GND 0.322f
C2575 VDD.n2447 GND 0.00418f
C2576 VDD.n2448 GND 0.00418f
C2577 VDD.n2449 GND 0.00418f
C2578 VDD.n2450 GND 0.00418f
C2579 VDD.n2451 GND 0.00418f
C2580 VDD.n2452 GND 0.322f
C2581 VDD.n2453 GND 0.00418f
C2582 VDD.n2454 GND 0.00418f
C2583 VDD.n2455 GND 0.00418f
C2584 VDD.n2456 GND 0.00418f
C2585 VDD.n2457 GND 0.00418f
C2586 VDD.n2458 GND 0.322f
C2587 VDD.n2459 GND 0.00418f
C2588 VDD.n2460 GND 0.00418f
C2589 VDD.n2461 GND 0.00418f
C2590 VDD.n2462 GND 0.00418f
C2591 VDD.n2463 GND 0.00418f
C2592 VDD.n2464 GND 0.322f
C2593 VDD.n2465 GND 0.00418f
C2594 VDD.n2466 GND 0.00418f
C2595 VDD.n2467 GND 0.00418f
C2596 VDD.n2468 GND 0.00418f
C2597 VDD.n2469 GND 0.00418f
C2598 VDD.n2470 GND 0.208353f
C2599 VDD.n2471 GND 0.00418f
C2600 VDD.n2472 GND 0.00418f
C2601 VDD.n2473 GND 0.00418f
C2602 VDD.n2474 GND 0.00418f
C2603 VDD.n2475 GND 0.00418f
C2604 VDD.n2476 GND 0.322f
C2605 VDD.n2477 GND 0.00418f
C2606 VDD.n2478 GND 0.00418f
C2607 VDD.n2479 GND 0.00418f
C2608 VDD.n2480 GND 0.00418f
C2609 VDD.n2481 GND 0.00418f
C2610 VDD.n2482 GND 0.322f
C2611 VDD.n2483 GND 0.00418f
C2612 VDD.n2484 GND 0.00418f
C2613 VDD.n2485 GND 0.00418f
C2614 VDD.n2486 GND 0.00418f
C2615 VDD.n2487 GND 0.00418f
C2616 VDD.n2488 GND 0.222559f
C2617 VDD.n2489 GND 0.00418f
C2618 VDD.n2490 GND 0.00418f
C2619 VDD.n2491 GND 0.00418f
C2620 VDD.n2492 GND 0.00418f
C2621 VDD.n2493 GND 0.00418f
C2622 VDD.n2494 GND 0.322f
C2623 VDD.n2495 GND 0.00418f
C2624 VDD.n2496 GND 0.00418f
C2625 VDD.n2497 GND 0.00418f
C2626 VDD.n2498 GND 0.00418f
C2627 VDD.n2499 GND 0.00418f
C2628 VDD.n2500 GND 0.322f
C2629 VDD.n2501 GND 0.00418f
C2630 VDD.n2502 GND 0.00418f
C2631 VDD.n2503 GND 0.00418f
C2632 VDD.n2504 GND 0.00418f
C2633 VDD.n2505 GND 0.00418f
C2634 VDD.n2506 GND 0.322f
C2635 VDD.n2507 GND 0.00418f
C2636 VDD.n2508 GND 0.00418f
C2637 VDD.n2509 GND 0.00418f
C2638 VDD.n2510 GND 0.00418f
C2639 VDD.n2511 GND 0.00418f
C2640 VDD.n2512 GND 0.322f
C2641 VDD.n2513 GND 0.00418f
C2642 VDD.n2514 GND 0.00418f
C2643 VDD.n2515 GND 0.00418f
C2644 VDD.n2516 GND 0.00418f
C2645 VDD.n2517 GND 0.00418f
C2646 VDD.n2518 GND 0.322f
C2647 VDD.n2519 GND 0.00418f
C2648 VDD.n2520 GND 0.00418f
C2649 VDD.n2521 GND 0.00418f
C2650 VDD.n2522 GND 0.00418f
C2651 VDD.n2523 GND 0.00418f
C2652 VDD.n2524 GND 0.284117f
C2653 VDD.n2525 GND 0.00418f
C2654 VDD.n2526 GND 0.00418f
C2655 VDD.n2527 GND 0.00418f
C2656 VDD.n2528 GND 0.00418f
C2657 VDD.n2529 GND 0.00418f
C2658 VDD.n2530 GND 0.322f
C2659 VDD.n2531 GND 0.00418f
C2660 VDD.n2532 GND 0.00418f
C2661 VDD.n2533 GND 0.00418f
C2662 VDD.n2534 GND 0.00418f
C2663 VDD.n2535 GND 0.00418f
C2664 VDD.n2536 GND 0.322f
C2665 VDD.n2537 GND 0.00418f
C2666 VDD.n2538 GND 0.00418f
C2667 VDD.n2539 GND 0.00418f
C2668 VDD.n2540 GND 0.00418f
C2669 VDD.n2541 GND 0.00418f
C2670 VDD.n2542 GND 0.322f
C2671 VDD.n2543 GND 0.00418f
C2672 VDD.n2544 GND 0.00418f
C2673 VDD.n2545 GND 0.00418f
C2674 VDD.n2546 GND 0.00418f
C2675 VDD.n2547 GND 0.00418f
C2676 VDD.n2548 GND 0.25097f
C2677 VDD.n2549 GND 0.00418f
C2678 VDD.n2550 GND 0.00418f
C2679 VDD.n2551 GND 0.00418f
C2680 VDD.n2552 GND 0.00418f
C2681 VDD.n2553 GND 0.00418f
C2682 VDD.n2554 GND 0.322f
C2683 VDD.n2555 GND 0.00418f
C2684 VDD.n2556 GND 0.00418f
C2685 VDD.n2557 GND 0.00418f
C2686 VDD.n2558 GND 0.00418f
C2687 VDD.n2559 GND 0.00418f
C2688 VDD.n2560 GND 0.322f
C2689 VDD.n2561 GND 0.00418f
C2690 VDD.n2562 GND 0.00418f
C2691 VDD.n2563 GND 0.00418f
C2692 VDD.n2564 GND 0.00418f
C2693 VDD.n2565 GND 0.00418f
C2694 VDD.n2566 GND 0.322f
C2695 VDD.n2567 GND 0.00418f
C2696 VDD.n2568 GND 0.00418f
C2697 VDD.n2569 GND 0.00418f
C2698 VDD.n2570 GND 0.00418f
C2699 VDD.n2571 GND 0.00418f
C2700 VDD.n2572 GND 0.322f
C2701 VDD.n2573 GND 0.00418f
C2702 VDD.n2574 GND 0.00418f
C2703 VDD.n2575 GND 0.00418f
C2704 VDD.n2576 GND 0.00418f
C2705 VDD.n2577 GND 0.00418f
C2706 VDD.n2578 GND 0.322f
C2707 VDD.n2579 GND 0.00418f
C2708 VDD.n2580 GND 0.00418f
C2709 VDD.n2581 GND 0.00418f
C2710 VDD.n2582 GND 0.00418f
C2711 VDD.n2583 GND 0.00418f
C2712 VDD.n2584 GND 0.322f
C2713 VDD.n2585 GND 0.00418f
C2714 VDD.n2586 GND 0.00418f
C2715 VDD.n2587 GND 0.00418f
C2716 VDD.n2588 GND 0.00418f
C2717 VDD.n2589 GND 0.00418f
C2718 VDD.n2590 GND 0.322f
C2719 VDD.n2591 GND 0.00418f
C2720 VDD.n2592 GND 0.00418f
C2721 VDD.n2593 GND 0.00418f
C2722 VDD.n2594 GND 0.00418f
C2723 VDD.n2595 GND 0.00418f
C2724 VDD.n2596 GND 0.322f
C2725 VDD.n2597 GND 0.00418f
C2726 VDD.n2598 GND 0.00418f
C2727 VDD.n2599 GND 0.00418f
C2728 VDD.n2600 GND 0.00418f
C2729 VDD.n2601 GND 0.00418f
C2730 VDD.n2602 GND 0.2415f
C2731 VDD.n2603 GND 0.00418f
C2732 VDD.n2604 GND 0.00418f
C2733 VDD.n2605 GND 0.00418f
C2734 VDD.n2606 GND 0.00418f
C2735 VDD.n2607 GND 0.00418f
C2736 VDD.n2608 GND 0.322f
C2737 VDD.n2609 GND 0.00418f
C2738 VDD.n2610 GND 0.00418f
C2739 VDD.n2611 GND 0.00418f
C2740 VDD.n2612 GND 0.00418f
C2741 VDD.n2613 GND 0.00418f
C2742 VDD.n2614 GND 0.322f
C2743 VDD.n2615 GND 0.00418f
C2744 VDD.n2616 GND 0.00418f
C2745 VDD.n2617 GND 0.00418f
C2746 VDD.n2618 GND 0.00418f
C2747 VDD.n2619 GND 0.00418f
C2748 VDD.n2620 GND 0.322f
C2749 VDD.n2621 GND 0.00418f
C2750 VDD.n2622 GND 0.00418f
C2751 VDD.n2623 GND 0.00418f
C2752 VDD.n2624 GND 0.00418f
C2753 VDD.n2625 GND 0.00418f
C2754 VDD.n2626 GND 0.322f
C2755 VDD.n2627 GND 0.00418f
C2756 VDD.n2628 GND 0.00418f
C2757 VDD.n2629 GND 0.00418f
C2758 VDD.n2630 GND 0.00418f
C2759 VDD.n2631 GND 0.00418f
C2760 VDD.n2632 GND 0.322f
C2761 VDD.n2633 GND 0.00418f
C2762 VDD.n2634 GND 0.00418f
C2763 VDD.n2635 GND 0.00418f
C2764 VDD.n2636 GND 0.00418f
C2765 VDD.n2637 GND 0.00418f
C2766 VDD.n2638 GND 0.322f
C2767 VDD.n2639 GND 0.00418f
C2768 VDD.n2640 GND 0.00418f
C2769 VDD.n2641 GND 0.00418f
C2770 VDD.n2642 GND 0.00418f
C2771 VDD.n2643 GND 0.00418f
C2772 VDD.n2644 GND 0.322f
C2773 VDD.n2645 GND 0.00418f
C2774 VDD.n2646 GND 0.00418f
C2775 VDD.n2647 GND 0.00418f
C2776 VDD.n2648 GND 0.00418f
C2777 VDD.n2649 GND 0.00418f
C2778 VDD.n2650 GND 0.322f
C2779 VDD.n2651 GND 0.00418f
C2780 VDD.n2652 GND 0.00418f
C2781 VDD.n2653 GND 0.00418f
C2782 VDD.n2654 GND 0.00418f
C2783 VDD.n2655 GND 0.00418f
C2784 VDD.n2656 GND 0.322f
C2785 VDD.n2657 GND 0.00418f
C2786 VDD.n2658 GND 0.00418f
C2787 VDD.n2659 GND 0.00418f
C2788 VDD.n2660 GND 0.00418f
C2789 VDD.n2661 GND 0.00418f
C2790 VDD.n2662 GND 0.232029f
C2791 VDD.n2663 GND 0.00418f
C2792 VDD.n2664 GND 0.00418f
C2793 VDD.n2665 GND 0.00418f
C2794 VDD.n2666 GND 0.00418f
C2795 VDD.n2667 GND 0.00418f
C2796 VDD.n2668 GND 0.17047f
C2797 VDD.n2669 GND 0.00418f
C2798 VDD.n2670 GND 0.00418f
C2799 VDD.n2671 GND 0.00418f
C2800 VDD.n2672 GND 0.00418f
C2801 VDD.n2673 GND 0.00418f
C2802 VDD.n2674 GND 0.322f
C2803 VDD.n2675 GND 0.00418f
C2804 VDD.n2676 GND 0.00418f
C2805 VDD.n2677 GND 0.00418f
C2806 VDD.n2678 GND 0.00418f
C2807 VDD.n2679 GND 0.00418f
C2808 VDD.n2680 GND 0.322f
C2809 VDD.n2681 GND 0.00418f
C2810 VDD.n2682 GND 0.00418f
C2811 VDD.n2683 GND 0.00418f
C2812 VDD.n2684 GND 0.00418f
C2813 VDD.n2685 GND 0.00418f
C2814 VDD.n2686 GND 0.322f
C2815 VDD.n2687 GND 0.00418f
C2816 VDD.n2688 GND 0.00418f
C2817 VDD.n2689 GND 0.00418f
C2818 VDD.n2690 GND 0.00418f
C2819 VDD.n2691 GND 0.00418f
C2820 VDD.n2692 GND 0.322f
C2821 VDD.n2693 GND 0.00418f
C2822 VDD.n2694 GND 0.00418f
C2823 VDD.n2695 GND 0.00418f
C2824 VDD.n2696 GND 0.00418f
C2825 VDD.n2697 GND 0.00418f
C2826 VDD.n2698 GND 0.322f
C2827 VDD.n2699 GND 0.00418f
C2828 VDD.n2700 GND 0.00418f
C2829 VDD.n2701 GND 0.00418f
C2830 VDD.n2702 GND 0.00418f
C2831 VDD.n2703 GND 0.00418f
C2832 VDD.n2704 GND 0.322f
C2833 VDD.n2705 GND 0.00418f
C2834 VDD.n2706 GND 0.00418f
C2835 VDD.n2707 GND 0.00418f
C2836 VDD.n2708 GND 0.00418f
C2837 VDD.n2709 GND 0.00418f
C2838 VDD.n2710 GND 0.322f
C2839 VDD.n2711 GND 0.00418f
C2840 VDD.n2712 GND 0.00418f
C2841 VDD.n2713 GND 0.00418f
C2842 VDD.n2714 GND 0.00418f
C2843 VDD.n2715 GND 0.00418f
C2844 VDD.n2716 GND 0.260441f
C2845 VDD.n2717 GND 0.00418f
C2846 VDD.n2718 GND 0.00418f
C2847 VDD.n2719 GND 0.00418f
C2848 VDD.n2720 GND 0.00418f
C2849 VDD.n2721 GND 0.00418f
C2850 VDD.n2722 GND 0.322f
C2851 VDD.n2723 GND 0.00418f
C2852 VDD.n2724 GND 0.00418f
C2853 VDD.n2725 GND 0.00418f
C2854 VDD.n2726 GND 0.00418f
C2855 VDD.n2727 GND 0.00418f
C2856 VDD.n2728 GND 0.303058f
C2857 VDD.n2729 GND 0.00418f
C2858 VDD.n2730 GND 0.00418f
C2859 VDD.n2731 GND 0.00418f
C2860 VDD.n2732 GND 0.00418f
C2861 VDD.n2733 GND 0.00418f
C2862 VDD.n2734 GND 0.322f
C2863 VDD.n2735 GND 0.00418f
C2864 VDD.n2736 GND 0.00418f
C2865 VDD.n2737 GND 0.00418f
C2866 VDD.n2738 GND 0.00418f
C2867 VDD.n2739 GND 0.00418f
C2868 VDD.n2740 GND 0.322f
C2869 VDD.n2741 GND 0.00418f
C2870 VDD.n2742 GND 0.00418f
C2871 VDD.n2743 GND 0.00418f
C2872 VDD.n2744 GND 0.00418f
C2873 VDD.n2745 GND 0.00418f
C2874 VDD.n2746 GND 0.322f
C2875 VDD.n2747 GND 0.00418f
C2876 VDD.n2748 GND 0.00418f
C2877 VDD.n2749 GND 0.00418f
C2878 VDD.n2750 GND 0.00418f
C2879 VDD.n2751 GND 0.00418f
C2880 VDD.n2752 GND 0.322f
C2881 VDD.n2753 GND 0.00418f
C2882 VDD.n2754 GND 0.00418f
C2883 VDD.n2755 GND 0.00418f
C2884 VDD.n2756 GND 0.00418f
C2885 VDD.n2757 GND 0.00418f
C2886 VDD.n2758 GND 0.322f
C2887 VDD.n2759 GND 0.00418f
C2888 VDD.n2760 GND 0.00418f
C2889 VDD.n2761 GND 0.00418f
C2890 VDD.n2762 GND 0.00418f
C2891 VDD.n2763 GND 0.00418f
C2892 VDD.n2764 GND 0.322f
C2893 VDD.n2765 GND 0.00418f
C2894 VDD.n2766 GND 0.00418f
C2895 VDD.n2767 GND 0.00418f
C2896 VDD.n2768 GND 0.00418f
C2897 VDD.n2769 GND 0.00418f
C2898 VDD.n2770 GND 0.322f
C2899 VDD.n2771 GND 0.00418f
C2900 VDD.n2772 GND 0.00418f
C2901 VDD.n2773 GND 0.00418f
C2902 VDD.n2774 GND 0.00418f
C2903 VDD.n2775 GND 0.00418f
C2904 VDD.n2776 GND 0.322f
C2905 VDD.n2777 GND 0.00418f
C2906 VDD.n2778 GND 0.00418f
C2907 VDD.n2779 GND 0.00418f
C2908 VDD.n2780 GND 0.00418f
C2909 VDD.n2781 GND 0.00418f
C2910 VDD.n2782 GND 0.189411f
C2911 VDD.n2783 GND 0.00418f
C2912 VDD.n2784 GND 0.00418f
C2913 VDD.n2785 GND 0.00418f
C2914 VDD.n2786 GND 0.00418f
C2915 VDD.n2787 GND 0.00418f
C2916 VDD.n2788 GND 0.184676f
C2917 VDD.n2789 GND 0.00418f
C2918 VDD.n2790 GND 0.00418f
C2919 VDD.n2791 GND 0.00418f
C2920 VDD.n2792 GND 0.00418f
C2921 VDD.n2793 GND 0.00418f
C2922 VDD.n2794 GND 0.322f
C2923 VDD.n2795 GND 0.00418f
C2924 VDD.n2796 GND 0.00418f
C2925 VDD.n2797 GND 0.00418f
C2926 VDD.n2798 GND 0.00418f
C2927 VDD.n2799 GND 0.00418f
C2928 VDD.n2800 GND 0.322f
C2929 VDD.n2801 GND 0.00418f
C2930 VDD.n2802 GND 0.00418f
C2931 VDD.n2803 GND 0.00418f
C2932 VDD.n2804 GND 0.00418f
C2933 VDD.n2805 GND 0.00418f
C2934 VDD.n2806 GND 0.00418f
C2935 VDD.n2807 GND 0.00418f
C2936 VDD.n2808 GND 0.00418f
C2937 VDD.n2809 GND 0.00418f
C2938 VDD.n2810 GND 0.00418f
C2939 VDD.n2811 GND 0.322f
C2940 VDD.n2812 GND 0.00418f
C2941 VDD.n2813 GND 0.00418f
C2942 VDD.n2814 GND 0.00418f
C2943 VDD.n2815 GND 0.00418f
C2944 VDD.n2816 GND 0.00418f
C2945 VDD.n2817 GND 0.322f
C2946 VDD.n2818 GND 0.00418f
C2947 VDD.n2819 GND 0.00418f
C2948 VDD.n2820 GND 0.00418f
C2949 VDD.n2821 GND 0.00418f
C2950 VDD.n2822 GND 0.009354f
C2951 VDD.n2823 GND 0.008807f
C2952 VDD.n2824 GND 0.009514f
C2953 VDD.n2825 GND 0.008967f
C2954 VDD.n2826 GND 0.00418f
C2955 VDD.n2827 GND 0.00418f
C2956 VDD.n2828 GND 0.00418f
C2957 VDD.n2829 GND 0.00418f
C2958 VDD.n2830 GND 0.003166f
C2959 VDD.n2831 GND 0.00418f
C2960 VDD.n2832 GND 0.00418f
C2961 VDD.n2833 GND 0.003105f
C2962 VDD.n2834 GND 0.00418f
C2963 VDD.n2835 GND 0.00418f
C2964 VDD.n2836 GND 0.00418f
C2965 VDD.n2837 GND 0.00418f
C2966 VDD.n2838 GND 0.00418f
C2967 VDD.n2839 GND 0.00418f
C2968 VDD.n2840 GND 0.00418f
C2969 VDD.n2841 GND 0.00418f
C2970 VDD.n2842 GND 0.00418f
C2971 VDD.n2843 GND 0.00418f
C2972 VDD.n2844 GND 0.00418f
C2973 VDD.n2845 GND 0.00418f
C2974 VDD.n2846 GND 0.00418f
C2975 VDD.n2847 GND 0.00418f
C2976 VDD.n2848 GND 0.00418f
C2977 VDD.n2849 GND 0.00418f
C2978 VDD.n2850 GND 0.00418f
C2979 VDD.n2851 GND 0.00418f
C2980 VDD.n2852 GND 0.00418f
C2981 VDD.n2853 GND 0.00418f
C2982 VDD.n2854 GND 0.00418f
C2983 VDD.n2855 GND 0.00418f
C2984 VDD.n2856 GND 0.00418f
C2985 VDD.n2857 GND 0.00418f
C2986 VDD.n2858 GND 0.009514f
C2987 VDD.n2859 GND 0.009514f
C2988 VDD.n2860 GND 0.008807f
C2989 VDD.n2861 GND 0.00418f
C2990 VDD.n2862 GND 0.00418f
C2991 VDD.n2863 GND 0.322f
C2992 VDD.n2864 GND 0.00418f
C2993 VDD.n2865 GND 0.008807f
C2994 VDD.n2866 GND 0.009354f
C2995 VDD.n2867 GND 0.008967f
C2996 VDD.n2868 GND 0.00418f
C2997 VDD.n2869 GND 0.00418f
C2998 VDD.n2870 GND 0.00418f
C2999 VDD.n2871 GND 0.00418f
C3000 VDD.n2872 GND 0.00418f
C3001 VDD.n2873 GND 0.003166f
C3002 VDD.n2874 GND 0.005158f
C3003 VDD.n2875 GND 0.003105f
C3004 VDD.n2876 GND 0.00418f
C3005 VDD.n2877 GND 0.00418f
C3006 VDD.n2878 GND 0.00418f
C3007 VDD.n2879 GND 0.00418f
C3008 VDD.n2880 GND 0.00418f
C3009 VDD.n2881 GND 0.00418f
C3010 VDD.n2882 GND 0.00418f
C3011 VDD.n2883 GND 0.00418f
C3012 VDD.n2884 GND 0.00418f
C3013 VDD.n2885 GND 0.00418f
C3014 VDD.n2886 GND 0.00418f
C3015 VDD.n2887 GND 0.00418f
C3016 VDD.n2888 GND 0.00418f
C3017 VDD.n2889 GND 0.00418f
C3018 VDD.n2890 GND 0.00418f
C3019 VDD.n2891 GND 0.00418f
C3020 VDD.n2892 GND 0.00418f
C3021 VDD.n2893 GND 0.00418f
C3022 VDD.n2894 GND 0.00418f
C3023 VDD.n2895 GND 0.00418f
C3024 VDD.n2896 GND 0.00418f
C3025 VDD.n2897 GND 0.00418f
C3026 VDD.n2898 GND 0.00418f
C3027 VDD.n2899 GND 0.00418f
C3028 VDD.n2900 GND 0.009514f
C3029 VDD.n2901 GND 0.009514f
C3030 VDD.n2902 GND 2.00539f
C3031 VDD.n2910 GND 0.009514f
C3032 VDD.n2919 GND 0.00418f
C3033 VDD.n2920 GND 0.00418f
C3034 VDD.t52 GND 0.089111f
C3035 VDD.t49 GND 0.44554f
C3036 VDD.n2921 GND 0.076053f
C3037 VDD.t51 GND 0.056759f
C3038 VDD.n2922 GND 0.078134f
C3039 VDD.n2923 GND 0.00418f
C3040 VDD.n2924 GND 0.00418f
C3041 VDD.n2925 GND 0.00418f
C3042 VDD.n2926 GND 0.00418f
C3043 VDD.n2927 GND 0.00418f
C3044 VDD.n2928 GND 0.00418f
C3045 VDD.n2929 GND 0.00418f
C3046 VDD.n2930 GND 0.00418f
C3047 VDD.n2931 GND 0.00418f
C3048 VDD.n2932 GND 0.00418f
C3049 VDD.n2933 GND 0.00418f
C3050 VDD.n2934 GND 0.00418f
C3051 VDD.n2935 GND 0.00418f
C3052 VDD.n2936 GND 0.00418f
C3053 VDD.n2937 GND 0.00418f
C3054 VDD.n2938 GND 0.00418f
C3055 VDD.n2939 GND 0.00418f
C3056 VDD.n2940 GND 0.00418f
C3057 VDD.n2941 GND 0.00418f
C3058 VDD.n2942 GND 0.00418f
C3059 VDD.n2943 GND 0.00418f
C3060 VDD.n2944 GND 0.00418f
C3061 VDD.n2945 GND 0.00418f
C3062 VDD.n2946 GND 0.00418f
C3063 VDD.n2947 GND 0.00418f
C3064 VDD.n2948 GND 0.00418f
C3065 VDD.n2949 GND 0.00418f
C3066 VDD.n2950 GND 0.00418f
C3067 VDD.n2951 GND 0.00418f
C3068 VDD.n2952 GND 0.00418f
C3069 VDD.n2953 GND 0.00418f
C3070 VDD.n2954 GND 0.00418f
C3071 VDD.n2955 GND 0.00418f
C3072 VDD.n2956 GND 0.00418f
C3073 VDD.n2957 GND 0.00418f
C3074 VDD.n2958 GND 0.00418f
C3075 VDD.n2959 GND 0.00418f
C3076 VDD.n2960 GND 0.00418f
C3077 VDD.n2961 GND 0.00418f
C3078 VDD.n2962 GND 0.00418f
C3079 VDD.n2963 GND 0.00418f
C3080 VDD.n2964 GND 0.00418f
C3081 VDD.n2965 GND 0.00418f
C3082 VDD.n2966 GND 0.00418f
C3083 VDD.n2967 GND 0.00418f
C3084 VDD.n2968 GND 0.00418f
C3085 VDD.n2969 GND 0.00418f
C3086 VDD.n2970 GND 0.00418f
C3087 VDD.n2971 GND 0.00418f
C3088 VDD.n2972 GND 0.00418f
C3089 VDD.n2973 GND 0.00418f
C3090 VDD.n2974 GND 0.00418f
C3091 VDD.n2975 GND 0.00418f
C3092 VDD.n2976 GND 0.00418f
C3093 VDD.n2977 GND 0.00418f
C3094 VDD.n2978 GND 0.00418f
C3095 VDD.n2979 GND 0.00418f
C3096 VDD.n2980 GND 0.00418f
C3097 VDD.n2981 GND 0.00418f
C3098 VDD.n2982 GND 0.00418f
C3099 VDD.n2983 GND 0.00418f
C3100 VDD.n2984 GND 0.00418f
C3101 VDD.n2985 GND 0.00418f
C3102 VDD.n2986 GND 0.00418f
C3103 VDD.n2987 GND 0.00418f
C3104 VDD.n2988 GND 0.00418f
C3105 VDD.n2989 GND 0.00418f
C3106 VDD.n2990 GND 0.00418f
C3107 VDD.n2991 GND 0.00418f
C3108 VDD.n2992 GND 0.00418f
C3109 VDD.n2993 GND 0.00418f
C3110 VDD.n2994 GND 0.00418f
C3111 VDD.n2995 GND 0.00418f
C3112 VDD.n2996 GND 0.00418f
C3113 VDD.n2997 GND 0.00418f
C3114 VDD.n2998 GND 0.00418f
C3115 VDD.n2999 GND 0.00418f
C3116 VDD.n3000 GND 0.00418f
C3117 VDD.n3001 GND 0.00418f
C3118 VDD.n3002 GND 0.00418f
C3119 VDD.n3003 GND 0.00418f
C3120 VDD.n3004 GND 0.00418f
C3121 VDD.n3005 GND 0.00418f
C3122 VDD.n3006 GND 0.00418f
C3123 VDD.n3007 GND 0.00418f
C3124 VDD.n3008 GND 0.00418f
C3125 VDD.n3009 GND 0.00418f
C3126 VDD.n3010 GND 0.00418f
C3127 VDD.n3011 GND 0.00418f
C3128 VDD.n3012 GND 0.00418f
C3129 VDD.n3013 GND 0.00418f
C3130 VDD.n3014 GND 0.00418f
C3131 VDD.n3015 GND 0.00418f
C3132 VDD.n3016 GND 0.00418f
C3133 VDD.n3017 GND 0.00418f
C3134 VDD.n3018 GND 0.00418f
C3135 VDD.n3019 GND 0.00418f
C3136 VDD.n3020 GND 0.00418f
C3137 VDD.n3021 GND 0.00418f
C3138 VDD.n3022 GND 0.00418f
C3139 VDD.n3023 GND 0.00418f
C3140 VDD.n3024 GND 0.00418f
C3141 VDD.n3025 GND 0.00418f
C3142 VDD.n3026 GND 0.00418f
C3143 VDD.n3027 GND 0.00418f
C3144 VDD.n3028 GND 0.00418f
C3145 VDD.n3029 GND 0.00418f
C3146 VDD.n3030 GND 0.00418f
C3147 VDD.n3031 GND 0.00418f
C3148 VDD.n3032 GND 0.00418f
C3149 VDD.n3033 GND 0.00418f
C3150 VDD.n3034 GND 0.00418f
C3151 VDD.n3035 GND 0.00418f
C3152 VDD.n3036 GND 0.00418f
C3153 VDD.n3037 GND 0.00418f
C3154 VDD.n3038 GND 0.00418f
C3155 VDD.n3039 GND 0.00418f
C3156 VDD.n3040 GND 0.00418f
C3157 VDD.n3041 GND 0.00418f
C3158 VDD.n3042 GND 0.00418f
C3159 VDD.n3043 GND 0.00418f
C3160 VDD.n3044 GND 0.00418f
C3161 VDD.n3045 GND 0.00418f
C3162 VDD.n3046 GND 0.00418f
C3163 VDD.n3047 GND 0.00418f
C3164 VDD.n3048 GND 0.00418f
C3165 VDD.n3049 GND 0.00418f
C3166 VDD.n3050 GND 0.00418f
C3167 VDD.n3051 GND 0.00418f
C3168 VDD.n3052 GND 0.00418f
C3169 VDD.n3053 GND 0.00418f
C3170 VDD.n3054 GND 0.00418f
C3171 VDD.n3055 GND 0.00418f
C3172 VDD.n3056 GND 0.00418f
C3173 VDD.n3057 GND 0.00418f
C3174 VDD.n3058 GND 0.00418f
C3175 VDD.n3059 GND 0.00418f
C3176 VDD.n3060 GND 0.00418f
C3177 VDD.n3061 GND 0.00418f
C3178 VDD.n3062 GND 0.00418f
C3179 VDD.n3063 GND 0.00418f
C3180 VDD.n3064 GND 0.00418f
C3181 VDD.n3065 GND 0.00418f
C3182 VDD.n3066 GND 0.00418f
C3183 VDD.n3067 GND 0.00418f
C3184 VDD.n3068 GND 0.00418f
C3185 VDD.n3069 GND 0.00418f
C3186 VDD.n3070 GND 0.00418f
C3187 VDD.n3071 GND 0.00418f
C3188 VDD.n3072 GND 0.00418f
C3189 VDD.n3073 GND 0.00418f
C3190 VDD.n3074 GND 0.00418f
C3191 VDD.n3075 GND 0.00418f
C3192 VDD.n3076 GND 0.00418f
C3193 VDD.n3077 GND 0.00418f
C3194 VDD.n3078 GND 0.00418f
C3195 VDD.n3079 GND 0.00418f
C3196 VDD.n3080 GND 0.00418f
C3197 VDD.n3081 GND 0.00418f
C3198 VDD.n3082 GND 0.00418f
C3199 VDD.n3083 GND 0.00418f
C3200 VDD.n3084 GND 0.00418f
C3201 VDD.n3085 GND 0.00418f
C3202 VDD.n3086 GND 0.00418f
C3203 VDD.n3087 GND 0.00418f
C3204 VDD.n3088 GND 0.00418f
C3205 VDD.n3089 GND 0.00418f
C3206 VDD.n3090 GND 0.00418f
C3207 VDD.n3091 GND 0.00418f
C3208 VDD.n3092 GND 0.00418f
C3209 VDD.n3093 GND 0.00418f
C3210 VDD.n3094 GND 0.00418f
C3211 VDD.n3095 GND 0.00418f
C3212 VDD.n3096 GND 0.00418f
C3213 VDD.n3097 GND 0.00418f
C3214 VDD.n3098 GND 0.00418f
C3215 VDD.n3099 GND 0.00418f
C3216 VDD.n3100 GND 0.00418f
C3217 VDD.n3101 GND 0.00418f
C3218 VDD.n3102 GND 0.00418f
C3219 VDD.n3103 GND 0.00418f
C3220 VDD.n3104 GND 0.00418f
C3221 VDD.n3105 GND 0.00418f
C3222 VDD.n3106 GND 0.00418f
C3223 VDD.n3107 GND 0.00418f
C3224 VDD.n3108 GND 0.00418f
C3225 VDD.n3109 GND 0.00418f
C3226 VDD.n3110 GND 0.00418f
C3227 VDD.n3111 GND 0.00418f
C3228 VDD.n3112 GND 0.00418f
C3229 VDD.n3113 GND 0.00418f
C3230 VDD.n3114 GND 0.00418f
C3231 VDD.n3115 GND 0.00418f
C3232 VDD.n3116 GND 0.00418f
C3233 VDD.t79 GND 0.089111f
C3234 VDD.t77 GND 0.44554f
C3235 VDD.n3117 GND 0.076053f
C3236 VDD.t78 GND 0.056759f
C3237 VDD.n3118 GND 0.078134f
C3238 VDD.n3119 GND 0.005158f
C3239 VDD.n3120 GND 0.00418f
C3240 VDD.n3121 GND 0.00418f
C3241 VDD.n3122 GND 0.00418f
C3242 VDD.n3123 GND 0.00418f
C3243 VDD.n3124 GND 0.00418f
C3244 VDD.n3125 GND 0.00418f
C3245 VDD.n3126 GND 0.00418f
C3246 VDD.n3127 GND 0.00418f
C3247 VDD.n3128 GND 0.00418f
C3248 VDD.n3129 GND 0.00418f
C3249 VDD.n3130 GND 0.00418f
C3250 VDD.n3131 GND 0.00418f
C3251 VDD.n3132 GND 0.00418f
C3252 VDD.n3133 GND 0.00418f
C3253 VDD.n3134 GND 0.00418f
C3254 VDD.n3135 GND 0.00418f
C3255 VDD.n3136 GND 0.00418f
C3256 VDD.n3137 GND 0.00418f
C3257 VDD.n3138 GND 0.00418f
C3258 VDD.n3139 GND 0.00418f
C3259 VDD.n3140 GND 0.00418f
C3260 VDD.n3141 GND 0.00418f
C3261 VDD.n3142 GND 0.003105f
C3262 VDD.n3143 GND 0.00418f
C3263 VDD.n3144 GND 0.00418f
C3264 VDD.n3145 GND 0.003166f
C3265 VDD.n3146 GND 0.00418f
C3266 VDD.n3147 GND 0.00418f
C3267 VDD.n3148 GND 0.00418f
C3268 VDD.n3149 GND 0.00418f
C3269 VDD.n3150 GND 0.009514f
C3270 VDD.n3151 GND 0.009514f
C3271 VDD.n3152 GND 0.008807f
C3272 VDD.n3153 GND 0.008807f
C3273 VDD.n3154 GND 0.00418f
C3274 VDD.n3155 GND 0.00418f
C3275 VDD.n3156 GND 0.00418f
C3276 VDD.n3157 GND 0.00418f
C3277 VDD.n3158 GND 0.00418f
C3278 VDD.n3159 GND 0.00418f
C3279 VDD.n3160 GND 0.00418f
C3280 VDD.n3161 GND 0.00418f
C3281 VDD.n3162 GND 0.00418f
C3282 VDD.n3163 GND 0.00418f
C3283 VDD.n3164 GND 0.00418f
C3284 VDD.n3165 GND 0.00418f
C3285 VDD.n3166 GND 0.00418f
C3286 VDD.n3167 GND 0.00418f
C3287 VDD.n3168 GND 0.00418f
C3288 VDD.n3169 GND 0.00418f
C3289 VDD.n3170 GND 0.00418f
C3290 VDD.n3171 GND 0.00418f
C3291 VDD.n3172 GND 0.00418f
C3292 VDD.n3173 GND 0.00418f
C3293 VDD.n3174 GND 0.00418f
C3294 VDD.n3175 GND 0.00418f
C3295 VDD.n3176 GND 0.00418f
C3296 VDD.n3177 GND 0.00418f
C3297 VDD.n3178 GND 0.00418f
C3298 VDD.n3179 GND 0.00418f
C3299 VDD.n3180 GND 0.00418f
C3300 VDD.n3181 GND 0.00418f
C3301 VDD.n3182 GND 0.00418f
C3302 VDD.n3183 GND 0.00418f
C3303 VDD.n3184 GND 0.00418f
C3304 VDD.n3185 GND 0.00418f
C3305 VDD.n3186 GND 0.00418f
C3306 VDD.n3187 GND 0.00418f
C3307 VDD.n3188 GND 0.00418f
C3308 VDD.n3189 GND 0.00418f
C3309 VDD.n3190 GND 0.00418f
C3310 VDD.n3191 GND 0.00418f
C3311 VDD.n3192 GND 0.00418f
C3312 VDD.n3193 GND 0.00418f
C3313 VDD.n3194 GND 0.00418f
C3314 VDD.n3195 GND 0.00418f
C3315 VDD.n3196 GND 0.00418f
C3316 VDD.n3197 GND 0.00418f
C3317 VDD.n3198 GND 0.00418f
C3318 VDD.n3199 GND 0.00418f
C3319 VDD.n3200 GND 0.00418f
C3320 VDD.n3201 GND 0.00418f
C3321 VDD.n3202 GND 0.00418f
C3322 VDD.n3203 GND 0.00418f
C3323 VDD.n3204 GND 0.00418f
C3324 VDD.n3205 GND 0.00418f
C3325 VDD.n3206 GND 0.00418f
C3326 VDD.n3207 GND 0.00418f
C3327 VDD.n3208 GND 0.00418f
C3328 VDD.n3209 GND 0.00418f
C3329 VDD.n3210 GND 0.00418f
C3330 VDD.n3211 GND 0.00418f
C3331 VDD.n3212 GND 0.00418f
C3332 VDD.n3213 GND 0.00418f
C3333 VDD.n3214 GND 0.00418f
C3334 VDD.n3215 GND 0.00418f
C3335 VDD.n3216 GND 0.00418f
C3336 VDD.n3217 GND 0.00418f
C3337 VDD.n3218 GND 0.00418f
C3338 VDD.n3219 GND 0.00418f
C3339 VDD.n3220 GND 0.00418f
C3340 VDD.n3221 GND 0.00418f
C3341 VDD.n3222 GND 0.00418f
C3342 VDD.n3223 GND 0.00418f
C3343 VDD.n3224 GND 0.00418f
C3344 VDD.n3225 GND 0.00418f
C3345 VDD.n3226 GND 0.00418f
C3346 VDD.n3227 GND 0.00418f
C3347 VDD.n3228 GND 0.00418f
C3348 VDD.n3229 GND 0.00418f
C3349 VDD.n3230 GND 0.00418f
C3350 VDD.n3231 GND 0.00418f
C3351 VDD.n3232 GND 0.00418f
C3352 VDD.n3233 GND 0.00418f
C3353 VDD.n3234 GND 0.00418f
C3354 VDD.n3235 GND 0.00418f
C3355 VDD.n3236 GND 0.00418f
C3356 VDD.n3237 GND 0.00418f
C3357 VDD.n3238 GND 0.00418f
C3358 VDD.n3239 GND 0.00418f
C3359 VDD.n3240 GND 0.00418f
C3360 VDD.n3241 GND 0.00418f
C3361 VDD.n3242 GND 0.00418f
C3362 VDD.n3243 GND 0.00418f
C3363 VDD.n3244 GND 0.00418f
C3364 VDD.n3245 GND 0.00418f
C3365 VDD.n3246 GND 0.00418f
C3366 VDD.n3247 GND 0.00418f
C3367 VDD.n3248 GND 0.00418f
C3368 VDD.n3249 GND 0.00418f
C3369 VDD.n3250 GND 0.00418f
C3370 VDD.n3251 GND 0.00418f
C3371 VDD.n3252 GND 0.00418f
C3372 VDD.n3253 GND 0.00418f
C3373 VDD.n3254 GND 0.00418f
C3374 VDD.n3255 GND 0.00418f
C3375 VDD.n3256 GND 0.00418f
C3376 VDD.n3257 GND 0.00418f
C3377 VDD.n3258 GND 0.00418f
C3378 VDD.n3259 GND 0.00418f
C3379 VDD.n3260 GND 0.00418f
C3380 VDD.n3261 GND 0.00418f
C3381 VDD.n3262 GND 0.00418f
C3382 VDD.n3263 GND 0.00418f
C3383 VDD.n3264 GND 0.00418f
C3384 VDD.n3265 GND 0.00418f
C3385 VDD.n3266 GND 0.00418f
C3386 VDD.n3267 GND 0.00418f
C3387 VDD.n3268 GND 0.00418f
C3388 VDD.n3269 GND 0.00418f
C3389 VDD.n3270 GND 0.00418f
C3390 VDD.n3271 GND 0.00418f
C3391 VDD.n3272 GND 0.00418f
C3392 VDD.n3273 GND 0.00418f
C3393 VDD.n3274 GND 0.00418f
C3394 VDD.n3275 GND 0.00418f
C3395 VDD.n3276 GND 0.00418f
C3396 VDD.n3277 GND 0.00418f
C3397 VDD.n3278 GND 0.00418f
C3398 VDD.n3279 GND 0.00418f
C3399 VDD.n3280 GND 0.00418f
C3400 VDD.n3281 GND 0.00418f
C3401 VDD.n3282 GND 0.00418f
C3402 VDD.n3283 GND 0.00418f
C3403 VDD.n3284 GND 0.00418f
C3404 VDD.n3285 GND 0.00418f
C3405 VDD.n3286 GND 0.00418f
C3406 VDD.n3287 GND 0.00418f
C3407 VDD.n3288 GND 0.00418f
C3408 VDD.n3289 GND 0.00418f
C3409 VDD.n3290 GND 0.00418f
C3410 VDD.n3291 GND 0.00418f
C3411 VDD.n3292 GND 0.00418f
C3412 VDD.n3293 GND 0.00418f
C3413 VDD.n3294 GND 0.00418f
C3414 VDD.n3295 GND 0.00418f
C3415 VDD.n3296 GND 0.00418f
C3416 VDD.n3297 GND 0.00418f
C3417 VDD.n3298 GND 0.00418f
C3418 VDD.n3299 GND 0.00418f
C3419 VDD.n3300 GND 0.00418f
C3420 VDD.n3301 GND 0.00418f
C3421 VDD.n3302 GND 0.00418f
C3422 VDD.n3303 GND 0.00418f
C3423 VDD.n3304 GND 0.00418f
C3424 VDD.n3305 GND 0.00418f
C3425 VDD.n3306 GND 0.00418f
C3426 VDD.n3307 GND 0.00418f
C3427 VDD.n3308 GND 0.00418f
C3428 VDD.n3309 GND 0.00418f
C3429 VDD.n3310 GND 0.00418f
C3430 VDD.n3311 GND 0.00418f
C3431 VDD.n3312 GND 0.00418f
C3432 VDD.n3313 GND 0.00418f
C3433 VDD.n3314 GND 0.00418f
C3434 VDD.n3315 GND 0.00418f
C3435 VDD.n3316 GND 0.00418f
C3436 VDD.n3317 GND 0.00418f
C3437 VDD.n3318 GND 0.00418f
C3438 VDD.n3319 GND 0.00418f
C3439 VDD.n3320 GND 0.00418f
C3440 VDD.n3321 GND 0.00418f
C3441 VDD.n3322 GND 0.00418f
C3442 VDD.n3323 GND 0.00418f
C3443 VDD.n3324 GND 0.00418f
C3444 VDD.n3325 GND 0.00418f
C3445 VDD.n3326 GND 0.00418f
C3446 VDD.n3327 GND 0.00418f
C3447 VDD.n3328 GND 0.00418f
C3448 VDD.n3329 GND 0.00418f
C3449 VDD.n3330 GND 0.00418f
C3450 VDD.n3331 GND 0.00418f
C3451 VDD.n3332 GND 0.00418f
C3452 VDD.n3333 GND 0.00418f
C3453 VDD.n3334 GND 0.00418f
C3454 VDD.n3335 GND 0.00418f
C3455 VDD.n3336 GND 0.00418f
C3456 VDD.n3337 GND 0.00418f
C3457 VDD.n3338 GND 0.00418f
C3458 VDD.n3339 GND 0.00418f
C3459 VDD.n3340 GND 0.00418f
C3460 VDD.n3341 GND 0.00418f
C3461 VDD.n3342 GND 0.00418f
C3462 VDD.n3343 GND 0.00418f
C3463 VDD.n3344 GND 0.00418f
C3464 VDD.n3345 GND 0.00418f
C3465 VDD.n3346 GND 0.00418f
C3466 VDD.n3347 GND 0.00418f
C3467 VDD.n3348 GND 0.00418f
C3468 VDD.n3349 GND 0.00418f
C3469 VDD.n3350 GND 0.00418f
C3470 VDD.n3351 GND 0.00418f
C3471 VDD.n3352 GND 0.00418f
C3472 VDD.n3353 GND 0.00418f
C3473 VDD.n3354 GND 0.00418f
C3474 VDD.n3355 GND 0.00418f
C3475 VDD.n3356 GND 0.00418f
C3476 VDD.n3357 GND 0.00418f
C3477 VDD.n3358 GND 0.00418f
C3478 VDD.n3359 GND 0.00418f
C3479 VDD.n3360 GND 0.00418f
C3480 VDD.n3361 GND 0.00418f
C3481 VDD.n3362 GND 0.00418f
C3482 VDD.n3363 GND 0.00418f
C3483 VDD.n3364 GND 0.00418f
C3484 VDD.n3365 GND 0.00418f
C3485 VDD.n3366 GND 0.00418f
C3486 VDD.n3367 GND 0.00418f
C3487 VDD.n3368 GND 0.00418f
C3488 VDD.n3369 GND 0.269911f
C3489 VDD.n3370 GND 0.00418f
C3490 VDD.n3371 GND 0.00418f
C3491 VDD.n3372 GND 0.00418f
C3492 VDD.n3373 GND 0.00418f
C3493 VDD.n3374 GND 0.00418f
C3494 VDD.n3375 GND 0.00418f
C3495 VDD.n3376 GND 0.00418f
C3496 VDD.n3377 GND 0.00418f
C3497 VDD.n3378 GND 0.00418f
C3498 VDD.n3379 GND 0.00418f
C3499 VDD.n3380 GND 0.00418f
C3500 VDD.n3381 GND 0.00418f
C3501 VDD.n3382 GND 0.00418f
C3502 VDD.n3383 GND 0.00418f
C3503 VDD.n3384 GND 0.00418f
C3504 VDD.n3385 GND 0.00418f
C3505 VDD.n3386 GND 0.00418f
C3506 VDD.n3387 GND 0.00418f
C3507 VDD.n3388 GND 0.008807f
C3508 VDD.n3389 GND 0.008807f
C3509 VDD.n3390 GND 0.009514f
C3510 VDD.n3391 GND 0.00418f
C3511 VDD.n3392 GND 0.00418f
C3512 VDD.n3393 GND 0.00418f
C3513 VDD.n3394 GND 0.00418f
C3514 VDD.n3395 GND 0.00418f
C3515 VDD.n3396 GND 0.003166f
C3516 VDD.n3397 GND 0.005158f
C3517 VDD.n3398 GND 0.003105f
C3518 VDD.n3399 GND 0.00418f
C3519 VDD.n3400 GND 0.00418f
C3520 VDD.n3401 GND 0.00418f
C3521 VDD.n3402 GND 0.00418f
C3522 VDD.n3403 GND 0.00418f
C3523 VDD.n3404 GND 0.00418f
C3524 VDD.n3405 GND 0.00418f
C3525 VDD.n3406 GND 0.00418f
C3526 VDD.n3407 GND 0.00418f
C3527 VDD.n3408 GND 0.00418f
C3528 VDD.n3409 GND 0.00418f
C3529 VDD.n3410 GND 0.00418f
C3530 VDD.n3411 GND 0.00418f
C3531 VDD.n3412 GND 0.00418f
C3532 VDD.n3413 GND 0.00418f
C3533 VDD.n3414 GND 0.00418f
C3534 VDD.n3415 GND 0.00418f
C3535 VDD.n3416 GND 0.00418f
C3536 VDD.n3417 GND 0.00418f
C3537 VDD.n3418 GND 0.00418f
C3538 VDD.n3419 GND 0.00418f
C3539 VDD.n3420 GND 0.00418f
C3540 VDD.n3421 GND 0.00418f
C3541 VDD.n3422 GND 0.009514f
C3542 VDD.n3423 GND 0.009514f
C3543 VDD.n3425 GND 2.00539f
C3544 VDD.n3427 GND 0.009514f
C3545 VDD.n3428 GND 0.009514f
C3546 VDD.n3429 GND 0.008807f
C3547 VDD.n3430 GND 0.00418f
C3548 VDD.n3431 GND 0.00418f
C3549 VDD.n3432 GND 0.322f
C3550 VDD.n3433 GND 0.00418f
C3551 VDD.n3434 GND 0.00418f
C3552 VDD.n3435 GND 0.00418f
C3553 VDD.n3436 GND 0.00418f
C3554 VDD.n3437 GND 0.00418f
C3555 VDD.n3438 GND 0.322f
C3556 VDD.n3439 GND 0.00418f
C3557 VDD.n3440 GND 0.00418f
C3558 VDD.n3441 GND 0.00418f
C3559 VDD.n3442 GND 0.00418f
C3560 VDD.n3443 GND 0.00418f
C3561 VDD.n3444 GND 0.322f
C3562 VDD.n3445 GND 0.00418f
C3563 VDD.n3446 GND 0.00418f
C3564 VDD.n3447 GND 0.00418f
C3565 VDD.n3448 GND 0.00418f
C3566 VDD.n3449 GND 0.00418f
C3567 VDD.n3450 GND 0.322f
C3568 VDD.n3451 GND 0.00418f
C3569 VDD.n3452 GND 0.00418f
C3570 VDD.n3453 GND 0.00418f
C3571 VDD.n3454 GND 0.00418f
C3572 VDD.n3455 GND 0.00418f
C3573 VDD.n3456 GND 0.322f
C3574 VDD.n3457 GND 0.00418f
C3575 VDD.n3458 GND 0.00418f
C3576 VDD.n3459 GND 0.00418f
C3577 VDD.n3460 GND 0.00418f
C3578 VDD.n3461 GND 0.00418f
C3579 VDD.n3462 GND 0.184676f
C3580 VDD.n3463 GND 0.00418f
C3581 VDD.n3464 GND 0.00418f
C3582 VDD.n3465 GND 0.00418f
C3583 VDD.n3466 GND 0.00418f
C3584 VDD.n3467 GND 0.00418f
C3585 VDD.n3468 GND 0.189411f
C3586 VDD.n3469 GND 0.00418f
C3587 VDD.n3470 GND 0.00418f
C3588 VDD.n3471 GND 0.00418f
C3589 VDD.n3472 GND 0.00418f
C3590 VDD.n3473 GND 0.00418f
C3591 VDD.n3474 GND 0.322f
C3592 VDD.n3475 GND 0.00418f
C3593 VDD.n3476 GND 0.00418f
C3594 VDD.n3477 GND 0.00418f
C3595 VDD.n3478 GND 0.00418f
C3596 VDD.n3479 GND 0.00418f
C3597 VDD.n3480 GND 0.322f
C3598 VDD.n3481 GND 0.00418f
C3599 VDD.n3482 GND 0.00418f
C3600 VDD.n3483 GND 0.00418f
C3601 VDD.n3484 GND 0.00418f
C3602 VDD.n3485 GND 0.00418f
C3603 VDD.n3486 GND 0.322f
C3604 VDD.n3487 GND 0.00418f
C3605 VDD.n3488 GND 0.00418f
C3606 VDD.n3489 GND 0.00418f
C3607 VDD.n3490 GND 0.00418f
C3608 VDD.n3491 GND 0.00418f
C3609 VDD.n3492 GND 0.322f
C3610 VDD.n3493 GND 0.00418f
C3611 VDD.n3494 GND 0.00418f
C3612 VDD.n3495 GND 0.00418f
C3613 VDD.n3496 GND 0.00418f
C3614 VDD.n3497 GND 0.00418f
C3615 VDD.n3498 GND 0.322f
C3616 VDD.n3499 GND 0.00418f
C3617 VDD.n3500 GND 0.00418f
C3618 VDD.n3501 GND 0.00418f
C3619 VDD.n3502 GND 0.00418f
C3620 VDD.n3503 GND 0.00418f
C3621 VDD.n3504 GND 0.322f
C3622 VDD.n3505 GND 0.00418f
C3623 VDD.n3506 GND 0.00418f
C3624 VDD.n3507 GND 0.00418f
C3625 VDD.n3508 GND 0.00418f
C3626 VDD.n3509 GND 0.00418f
C3627 VDD.n3510 GND 0.322f
C3628 VDD.n3511 GND 0.00418f
C3629 VDD.n3512 GND 0.00418f
C3630 VDD.n3513 GND 0.00418f
C3631 VDD.n3514 GND 0.00418f
C3632 VDD.n3515 GND 0.00418f
C3633 VDD.n3516 GND 0.322f
C3634 VDD.n3517 GND 0.00418f
C3635 VDD.n3518 GND 0.00418f
C3636 VDD.n3519 GND 0.00418f
C3637 VDD.n3520 GND 0.00418f
C3638 VDD.n3521 GND 0.00418f
C3639 VDD.n3522 GND 0.303058f
C3640 VDD.n3523 GND 0.00418f
C3641 VDD.n3524 GND 0.00418f
C3642 VDD.n3525 GND 0.00418f
C3643 VDD.n3526 GND 0.00418f
C3644 VDD.n3527 GND 0.00418f
C3645 VDD.n3528 GND 0.322f
C3646 VDD.n3529 GND 0.00418f
C3647 VDD.n3530 GND 0.00418f
C3648 VDD.n3531 GND 0.00418f
C3649 VDD.n3532 GND 0.00418f
C3650 VDD.n3533 GND 0.00418f
C3651 VDD.n3534 GND 0.260441f
C3652 VDD.n3535 GND 0.00418f
C3653 VDD.n3536 GND 0.00418f
C3654 VDD.n3537 GND 0.00418f
C3655 VDD.n3538 GND 0.00418f
C3656 VDD.n3539 GND 0.00418f
C3657 VDD.n3540 GND 0.322f
C3658 VDD.n3541 GND 0.00418f
C3659 VDD.n3542 GND 0.00418f
C3660 VDD.n3543 GND 0.00418f
C3661 VDD.n3544 GND 0.00418f
C3662 VDD.n3545 GND 0.00418f
C3663 VDD.n3546 GND 0.322f
C3664 VDD.n3547 GND 0.00418f
C3665 VDD.n3548 GND 0.00418f
C3666 VDD.n3549 GND 0.00418f
C3667 VDD.n3550 GND 0.00418f
C3668 VDD.n3551 GND 0.00418f
C3669 VDD.n3552 GND 0.322f
C3670 VDD.n3553 GND 0.00418f
C3671 VDD.n3554 GND 0.00418f
C3672 VDD.n3555 GND 0.00418f
C3673 VDD.n3556 GND 0.00418f
C3674 VDD.n3557 GND 0.00418f
C3675 VDD.n3558 GND 0.322f
C3676 VDD.n3559 GND 0.00418f
C3677 VDD.n3560 GND 0.00418f
C3678 VDD.n3561 GND 0.00418f
C3679 VDD.n3562 GND 0.00418f
C3680 VDD.n3563 GND 0.00418f
C3681 VDD.n3564 GND 0.322f
C3682 VDD.n3565 GND 0.00418f
C3683 VDD.n3566 GND 0.00418f
C3684 VDD.n3567 GND 0.00418f
C3685 VDD.n3568 GND 0.00418f
C3686 VDD.n3569 GND 0.00418f
C3687 VDD.n3570 GND 0.322f
C3688 VDD.n3571 GND 0.00418f
C3689 VDD.n3572 GND 0.00418f
C3690 VDD.n3573 GND 0.00418f
C3691 VDD.n3574 GND 0.00418f
C3692 VDD.n3575 GND 0.00418f
C3693 VDD.n3576 GND 0.322f
C3694 VDD.n3577 GND 0.00418f
C3695 VDD.n3578 GND 0.00418f
C3696 VDD.n3579 GND 0.00418f
C3697 VDD.n3580 GND 0.00418f
C3698 VDD.n3581 GND 0.00418f
C3699 VDD.n3582 GND 0.17047f
C3700 VDD.n3583 GND 0.00418f
C3701 VDD.n3584 GND 0.00418f
C3702 VDD.n3585 GND 0.00418f
C3703 VDD.n3586 GND 0.00418f
C3704 VDD.n3587 GND 0.00418f
C3705 VDD.n3588 GND 0.232029f
C3706 VDD.n3589 GND 0.00418f
C3707 VDD.n3590 GND 0.00418f
C3708 VDD.n3591 GND 0.00418f
C3709 VDD.n3592 GND 0.00418f
C3710 VDD.n3593 GND 0.00418f
C3711 VDD.n3594 GND 0.322f
C3712 VDD.n3595 GND 0.00418f
C3713 VDD.n3596 GND 0.00418f
C3714 VDD.n3597 GND 0.00418f
C3715 VDD.n3598 GND 0.00418f
C3716 VDD.n3599 GND 0.00418f
C3717 VDD.n3600 GND 0.322f
C3718 VDD.n3601 GND 0.00418f
C3719 VDD.n3602 GND 0.00418f
C3720 VDD.n3603 GND 0.00418f
C3721 VDD.n3604 GND 0.00418f
C3722 VDD.n3605 GND 0.00418f
C3723 VDD.n3606 GND 0.322f
C3724 VDD.n3607 GND 0.00418f
C3725 VDD.n3608 GND 0.00418f
C3726 VDD.n3609 GND 0.00418f
C3727 VDD.n3610 GND 0.00418f
C3728 VDD.n3611 GND 0.00418f
C3729 VDD.n3612 GND 0.322f
C3730 VDD.n3613 GND 0.00418f
C3731 VDD.n3614 GND 0.00418f
C3732 VDD.n3615 GND 0.00418f
C3733 VDD.n3616 GND 0.00418f
C3734 VDD.n3617 GND 0.00418f
C3735 VDD.n3618 GND 0.322f
C3736 VDD.n3619 GND 0.00418f
C3737 VDD.n3620 GND 0.00418f
C3738 VDD.n3621 GND 0.00418f
C3739 VDD.n3622 GND 0.00418f
C3740 VDD.n3623 GND 0.00418f
C3741 VDD.n3624 GND 0.322f
C3742 VDD.n3625 GND 0.00418f
C3743 VDD.n3626 GND 0.00418f
C3744 VDD.n3627 GND 0.00418f
C3745 VDD.n3628 GND 0.00418f
C3746 VDD.n3629 GND 0.00418f
C3747 VDD.n3630 GND 0.322f
C3748 VDD.n3631 GND 0.00418f
C3749 VDD.n3632 GND 0.00418f
C3750 VDD.n3633 GND 0.00418f
C3751 VDD.n3634 GND 0.00418f
C3752 VDD.n3635 GND 0.00418f
C3753 VDD.n3636 GND 0.322f
C3754 VDD.n3637 GND 0.00418f
C3755 VDD.n3638 GND 0.00418f
C3756 VDD.n3639 GND 0.00418f
C3757 VDD.n3640 GND 0.00418f
C3758 VDD.n3641 GND 0.00418f
C3759 VDD.n3642 GND 0.322f
C3760 VDD.n3643 GND 0.00418f
C3761 VDD.n3644 GND 0.00418f
C3762 VDD.n3645 GND 0.00418f
C3763 VDD.n3646 GND 0.00418f
C3764 VDD.n3647 GND 0.00418f
C3765 VDD.n3648 GND 0.2415f
C3766 VDD.n3649 GND 0.00418f
C3767 VDD.n3650 GND 0.00418f
C3768 VDD.n3651 GND 0.00418f
C3769 VDD.n3652 GND 0.00418f
C3770 VDD.n3653 GND 0.00418f
C3771 VDD.n3654 GND 0.322f
C3772 VDD.n3655 GND 0.00418f
C3773 VDD.n3656 GND 0.00418f
C3774 VDD.n3657 GND 0.00418f
C3775 VDD.n3658 GND 0.00418f
C3776 VDD.n3659 GND 0.00418f
C3777 VDD.n3660 GND 0.322f
C3778 VDD.n3661 GND 0.00418f
C3779 VDD.n3662 GND 0.00418f
C3780 VDD.n3663 GND 0.00418f
C3781 VDD.n3664 GND 0.00418f
C3782 VDD.n3665 GND 0.00418f
C3783 VDD.n3666 GND 0.322f
C3784 VDD.n3667 GND 0.00418f
C3785 VDD.n3668 GND 0.00418f
C3786 VDD.n3669 GND 0.00418f
C3787 VDD.n3670 GND 0.00418f
C3788 VDD.n3671 GND 0.00418f
C3789 VDD.n3672 GND 0.322f
C3790 VDD.n3673 GND 0.00418f
C3791 VDD.n3674 GND 0.00418f
C3792 VDD.n3675 GND 0.00418f
C3793 VDD.n3676 GND 0.00418f
C3794 VDD.n3677 GND 0.00418f
C3795 VDD.n3678 GND 0.322f
C3796 VDD.n3679 GND 0.00418f
C3797 VDD.n3680 GND 0.00418f
C3798 VDD.n3681 GND 0.00418f
C3799 VDD.n3682 GND 0.00418f
C3800 VDD.n3683 GND 0.00418f
C3801 VDD.n3684 GND 0.322f
C3802 VDD.n3685 GND 0.00418f
C3803 VDD.n3686 GND 0.00418f
C3804 VDD.n3687 GND 0.00418f
C3805 VDD.n3688 GND 0.00418f
C3806 VDD.n3689 GND 0.00418f
C3807 VDD.n3690 GND 0.322f
C3808 VDD.n3691 GND 0.00418f
C3809 VDD.n3692 GND 0.00418f
C3810 VDD.n3693 GND 0.00418f
C3811 VDD.n3694 GND 0.00418f
C3812 VDD.n3695 GND 0.00418f
C3813 VDD.n3696 GND 0.322f
C3814 VDD.n3697 GND 0.00418f
C3815 VDD.n3698 GND 0.00418f
C3816 VDD.n3699 GND 0.00418f
C3817 VDD.n3700 GND 0.00418f
C3818 VDD.n3701 GND 0.00418f
C3819 VDD.n3702 GND 0.25097f
C3820 VDD.n3703 GND 0.00418f
C3821 VDD.n3704 GND 0.00418f
C3822 VDD.n3705 GND 0.00418f
C3823 VDD.n3706 GND 0.00418f
C3824 VDD.n3707 GND 0.00418f
C3825 VDD.n3708 GND 0.322f
C3826 VDD.n3709 GND 0.00418f
C3827 VDD.n3710 GND 0.00418f
C3828 VDD.n3711 GND 0.00418f
C3829 VDD.n3712 GND 0.00418f
C3830 VDD.n3713 GND 0.00418f
C3831 VDD.n3714 GND 0.322f
C3832 VDD.n3715 GND 0.00418f
C3833 VDD.n3716 GND 0.00418f
C3834 VDD.n3717 GND 0.00418f
C3835 VDD.n3718 GND 0.00418f
C3836 VDD.n3719 GND 0.00418f
C3837 VDD.n3720 GND 0.322f
C3838 VDD.n3721 GND 0.00418f
C3839 VDD.n3722 GND 0.00418f
C3840 VDD.n3723 GND 0.00418f
C3841 VDD.n3724 GND 0.00418f
C3842 VDD.n3725 GND 0.00418f
C3843 VDD.n3726 GND 0.284117f
C3844 VDD.n3727 GND 0.00418f
C3845 VDD.n3728 GND 0.00418f
C3846 VDD.n3729 GND 0.00418f
C3847 VDD.n3730 GND 0.00418f
C3848 VDD.n3731 GND 0.00418f
C3849 VDD.n3732 GND 0.322f
C3850 VDD.n3733 GND 0.00418f
C3851 VDD.n3734 GND 0.00418f
C3852 VDD.n3735 GND 0.00418f
C3853 VDD.n3736 GND 0.00418f
C3854 VDD.n3737 GND 0.00418f
C3855 VDD.n3738 GND 0.322f
C3856 VDD.n3739 GND 0.00418f
C3857 VDD.n3740 GND 0.00418f
C3858 VDD.n3741 GND 0.00418f
C3859 VDD.n3742 GND 0.00418f
C3860 VDD.n3743 GND 0.00418f
C3861 VDD.n3744 GND 0.322f
C3862 VDD.n3745 GND 0.00418f
C3863 VDD.n3746 GND 0.00418f
C3864 VDD.n3747 GND 0.00418f
C3865 VDD.n3748 GND 0.00418f
C3866 VDD.n3749 GND 0.00418f
C3867 VDD.n3750 GND 0.322f
C3868 VDD.n3751 GND 0.00418f
C3869 VDD.n3752 GND 0.00418f
C3870 VDD.n3753 GND 0.00418f
C3871 VDD.n3754 GND 0.00418f
C3872 VDD.n3755 GND 0.00418f
C3873 VDD.n3756 GND 0.322f
C3874 VDD.n3757 GND 0.00418f
C3875 VDD.n3758 GND 0.00418f
C3876 VDD.n3759 GND 0.00418f
C3877 VDD.n3760 GND 0.00418f
C3878 VDD.n3761 GND 0.00418f
C3879 VDD.n3762 GND 0.222559f
C3880 VDD.n3763 GND 0.00418f
C3881 VDD.n3764 GND 0.00418f
C3882 VDD.n3765 GND 0.00418f
C3883 VDD.n3766 GND 0.00418f
C3884 VDD.n3767 GND 0.00418f
C3885 VDD.n3768 GND 0.322f
C3886 VDD.n3769 GND 0.00418f
C3887 VDD.n3770 GND 0.00418f
C3888 VDD.n3771 GND 0.00418f
C3889 VDD.n3772 GND 0.00418f
C3890 VDD.n3773 GND 0.00418f
C3891 VDD.n3774 GND 0.322f
C3892 VDD.n3775 GND 0.00418f
C3893 VDD.n3776 GND 0.00418f
C3894 VDD.n3777 GND 0.00418f
C3895 VDD.n3778 GND 0.00418f
C3896 VDD.n3779 GND 0.00418f
C3897 VDD.n3780 GND 0.208353f
C3898 VDD.n3781 GND 0.00418f
C3899 VDD.n3782 GND 0.00418f
C3900 VDD.n3783 GND 0.00418f
C3901 VDD.n3784 GND 0.00418f
C3902 VDD.n3785 GND 0.00418f
C3903 VDD.n3786 GND 0.322f
C3904 VDD.n3787 GND 0.00418f
C3905 VDD.n3788 GND 0.00418f
C3906 VDD.n3789 GND 0.00418f
C3907 VDD.n3790 GND 0.00418f
C3908 VDD.n3791 GND 0.00418f
C3909 VDD.n3792 GND 0.322f
C3910 VDD.n3793 GND 0.00418f
C3911 VDD.n3794 GND 0.00418f
C3912 VDD.n3795 GND 0.00418f
C3913 VDD.n3796 GND 0.00418f
C3914 VDD.n3797 GND 0.00418f
C3915 VDD.n3798 GND 0.322f
C3916 VDD.n3799 GND 0.00418f
C3917 VDD.n3800 GND 0.00418f
C3918 VDD.n3801 GND 0.00418f
C3919 VDD.n3802 GND 0.00418f
C3920 VDD.n3803 GND 0.00418f
C3921 VDD.n3804 GND 0.322f
C3922 VDD.n3805 GND 0.00418f
C3923 VDD.n3806 GND 0.00418f
C3924 VDD.n3807 GND 0.00418f
C3925 VDD.n3808 GND 0.00418f
C3926 VDD.n3809 GND 0.00418f
C3927 VDD.n3810 GND 0.322f
C3928 VDD.n3811 GND 0.00418f
C3929 VDD.n3812 GND 0.00418f
C3930 VDD.n3813 GND 0.00418f
C3931 VDD.n3814 GND 0.00418f
C3932 VDD.n3815 GND 0.00418f
C3933 VDD.n3816 GND 0.322f
C3934 VDD.n3817 GND 0.00418f
C3935 VDD.n3818 GND 0.00418f
C3936 VDD.n3819 GND 0.00418f
C3937 VDD.n3820 GND 0.00418f
C3938 VDD.n3821 GND 0.00418f
C3939 VDD.n3822 GND 0.322f
C3940 VDD.n3823 GND 0.00418f
C3941 VDD.n3824 GND 0.00418f
C3942 VDD.n3825 GND 0.00418f
C3943 VDD.n3826 GND 0.00418f
C3944 VDD.n3827 GND 0.00418f
C3945 VDD.n3828 GND 0.298323f
C3946 VDD.n3829 GND 0.00418f
C3947 VDD.n3830 GND 0.00418f
C3948 VDD.n3831 GND 0.00418f
C3949 VDD.n3832 GND 0.00418f
C3950 VDD.n3833 GND 0.00418f
C3951 VDD.n3834 GND 0.322f
C3952 VDD.n3835 GND 0.00418f
C3953 VDD.n3836 GND 0.00418f
C3954 VDD.n3837 GND 0.00418f
C3955 VDD.n3838 GND 0.00418f
C3956 VDD.n3839 GND 0.00418f
C3957 VDD.n3840 GND 0.265176f
C3958 VDD.n3841 GND 0.00418f
C3959 VDD.n3842 GND 0.00418f
C3960 VDD.n3843 GND 0.00418f
C3961 VDD.n3844 GND 0.00418f
C3962 VDD.n3845 GND 0.00418f
C3963 VDD.n3846 GND 0.322f
C3964 VDD.n3847 GND 0.00418f
C3965 VDD.n3848 GND 0.00418f
C3966 VDD.n3849 GND 0.00418f
C3967 VDD.n3850 GND 0.00418f
C3968 VDD.n3851 GND 0.00418f
C3969 VDD.n3852 GND 0.00418f
C3970 VDD.n3853 GND 0.00418f
C3971 VDD.n3855 GND 0.00418f
C3972 VDD.n3856 GND 0.00418f
C3973 VDD.n3857 GND 0.00418f
C3974 VDD.n3859 GND 0.00418f
C3975 VDD.n3860 GND 0.00418f
C3976 VDD.n3861 GND 0.00418f
C3977 VDD.n3862 GND 0.00418f
C3978 VDD.n3863 GND 0.00418f
C3979 VDD.n3864 GND 0.00418f
C3980 VDD.n3866 GND 0.00418f
C3981 VDD.n3867 GND 0.00418f
C3982 VDD.n3869 GND 0.009514f
C3983 VDD.n3870 GND 0.009514f
C3984 VDD.n3871 GND 0.008807f
C3985 VDD.n3872 GND 0.00418f
C3986 VDD.n3873 GND 0.00418f
C3987 VDD.n3874 GND 0.00418f
C3988 VDD.n3875 GND 0.00418f
C3989 VDD.n3876 GND 0.00418f
C3990 VDD.n3877 GND 0.00418f
C3991 VDD.n3878 GND 0.322f
C3992 VDD.n3879 GND 0.00418f
C3993 VDD.n3880 GND 0.00418f
C3994 VDD.n3881 GND 0.00418f
C3995 VDD.n3882 GND 0.00418f
C3996 VDD.n3883 GND 0.00418f
C3997 VDD.n3884 GND 0.322f
C3998 VDD.n3885 GND 0.00418f
C3999 VDD.n3886 GND 0.00418f
C4000 VDD.n3887 GND 0.00418f
C4001 VDD.n3888 GND 0.009354f
C4002 VDD.n3890 GND 0.009514f
C4003 VDD.n3891 GND 0.008967f
C4004 VDD.n3892 GND 0.00418f
C4005 VDD.n3893 GND 0.00418f
C4006 VDD.n3894 GND 0.00418f
C4007 VDD.n3896 GND 0.00418f
C4008 VDD.n3897 GND 0.00418f
C4009 VDD.n3898 GND 0.003105f
C4010 VDD.n3899 GND 0.00418f
C4011 VDD.n3900 GND 0.00418f
C4012 VDD.n3901 GND 0.00418f
C4013 VDD.n3903 GND 0.00418f
C4014 VDD.n3904 GND 0.00418f
C4015 VDD.n3905 GND 0.003135f
C4016 VDD.n3906 GND 1.05157f
C4017 VDD.n3907 GND 0.06079f
C4018 VDD.n3908 GND 0.003135f
C4019 VDD.n3909 GND 0.00418f
C4020 VDD.n3910 GND 0.00418f
C4021 VDD.n3912 GND 0.00418f
C4022 VDD.n3913 GND 0.00418f
C4023 VDD.n3914 GND 0.00418f
C4024 VDD.n3915 GND 0.00418f
C4025 VDD.n3916 GND 0.00418f
C4026 VDD.n3917 GND 0.00418f
C4027 VDD.n3919 GND 0.00418f
C4028 VDD.n3920 GND 0.00418f
C4029 VDD.n3921 GND 0.00418f
C4030 VDD.n3922 GND 0.009514f
C4031 VDD.n3923 GND 0.008807f
C4032 VDD.n3924 GND 0.008807f
C4033 VDD.n3925 GND 0.447485f
C4034 VDD.n3926 GND 0.008807f
C4035 VDD.n3927 GND 0.009514f
C4036 VDD.n3928 GND 0.008967f
C4037 VDD.n3929 GND 0.00418f
C4038 VDD.n3930 GND 0.00418f
C4039 VDD.n3931 GND 0.00418f
C4040 VDD.n3933 GND 0.00418f
C4041 VDD.n3934 GND 0.00418f
C4042 VDD.n3935 GND 0.003105f
C4043 VDD.n3936 GND 0.00418f
C4044 VDD.n3937 GND 0.00418f
C4045 VDD.n3938 GND 0.00418f
C4046 VDD.n3940 GND 0.00418f
C4047 VDD.n3941 GND 0.00418f
C4048 VDD.n3942 GND 0.003135f
C4049 VDD.n3943 GND 0.06079f
C4050 VDD.t13 GND 0.085164f
C4051 VDD.t10 GND 0.430073f
C4052 VDD.n3944 GND 0.075426f
C4053 VDD.t12 GND 0.053191f
C4054 VDD.n3945 GND 0.077435f
C4055 VDD.n3946 GND 0.006804f
C4056 VDD.n3947 GND 0.006148f
C4057 VDD.n3948 GND 0.006148f
C4058 VDD.n3949 GND 0.003093f
C4059 VDD.n3950 GND 0.004948f
C4060 VDD.n3951 GND 0.006148f
C4061 VDD.n3952 GND 0.006148f
C4062 VDD.n3953 GND 0.006148f
C4063 VDD.n3954 GND 0.006148f
C4064 VDD.n3955 GND 0.006148f
C4065 VDD.n3956 GND 0.006148f
C4066 VDD.n3957 GND 0.006148f
C4067 VDD.n3958 GND 0.006148f
C4068 VDD.n3959 GND 0.006148f
C4069 VDD.n3960 GND 0.002944f
C4070 VDD.n3961 GND 0.006148f
C4071 VDD.n3962 GND 0.014117f
C4072 VDD.n3963 GND 0.006148f
C4073 VDD.t64 GND 0.085164f
C4074 VDD.t62 GND 0.430073f
C4075 VDD.n3964 GND 0.075426f
C4076 VDD.t63 GND 0.053191f
C4077 VDD.n3965 GND 0.077435f
C4078 VDD.n3966 GND 0.009278f
C4079 VDD.n3967 GND 0.004478f
C4080 VDD.n3968 GND 0.006148f
C4081 VDD.n3969 GND 0.006148f
C4082 VDD.n3970 GND 0.004948f
C4083 VDD.n3971 GND 0.004948f
C4084 VDD.n3972 GND 0.006148f
C4085 VDD.n3973 GND 0.006148f
C4086 VDD.n3974 GND 0.004948f
C4087 VDD.n3975 GND 0.004948f
C4088 VDD.n3976 GND 0.006148f
C4089 VDD.n3977 GND 0.006148f
C4090 VDD.n3978 GND 0.004948f
C4091 VDD.n3979 GND 0.004948f
C4092 VDD.n3980 GND 0.006148f
C4093 VDD.n3981 GND 0.006148f
C4094 VDD.n3982 GND 0.004948f
C4095 VDD.n3983 GND 0.004948f
C4096 VDD.n3985 GND 1.05157f
C4097 VDD.n3986 GND 0.005287f
C4098 VDD.n3987 GND 0.004948f
C4099 VDD.n3988 GND 0.006148f
C4100 VDD.n3989 GND 0.006148f
C4101 VDD.n3990 GND 0.004948f
C4102 VDD.n3991 GND 0.004948f
C4103 VDD.n3992 GND 0.006148f
C4104 VDD.n3993 GND 0.006148f
C4105 VDD.n3994 GND 0.004948f
C4106 VDD.n3995 GND 0.004948f
C4107 VDD.n3996 GND 0.006148f
C4108 VDD.n3997 GND 0.006148f
C4109 VDD.n3998 GND 0.004948f
C4110 VDD.n3999 GND 0.004948f
C4111 VDD.n4000 GND 0.006148f
C4112 VDD.n4001 GND 0.006148f
C4113 VDD.n4002 GND 0.004948f
C4114 VDD.n4003 GND 0.004948f
C4115 VDD.n4004 GND 0.006148f
C4116 VDD.n4005 GND 0.006148f
C4117 VDD.n4006 GND 0.004874f
C4118 VDD.n4007 GND 0.009278f
C4119 VDD.n4008 GND 0.006148f
C4120 VDD.n4009 GND 0.006148f
C4121 VDD.n4010 GND 0.00339f
C4122 VDD.n4011 GND 0.004948f
C4123 VDD.n4012 GND 0.006148f
C4124 VDD.n4013 GND 0.006148f
C4125 VDD.n4014 GND 0.004948f
C4126 VDD.n4015 GND 0.004948f
C4127 VDD.n4016 GND 0.006148f
C4128 VDD.n4017 GND 0.006148f
C4129 VDD.n4018 GND 0.004948f
C4130 VDD.n4019 GND 0.004948f
C4131 VDD.n4020 GND 0.006148f
C4132 VDD.n4021 GND 0.006148f
C4133 VDD.n4022 GND 0.004948f
C4134 VDD.n4023 GND 0.004948f
C4135 VDD.n4024 GND 0.006148f
C4136 VDD.n4025 GND 0.006148f
C4137 VDD.n4026 GND 0.004948f
C4138 VDD.n4027 GND 0.006148f
C4139 VDD.n4028 GND 0.006148f
C4140 VDD.n4029 GND 0.004948f
C4141 VDD.n4030 GND 0.006148f
C4142 VDD.n4031 GND 0.006148f
C4143 VDD.n4032 GND 0.006148f
C4144 VDD.t38 GND 0.085164f
C4145 VDD.t36 GND 0.430073f
C4146 VDD.n4033 GND 0.075426f
C4147 VDD.t37 GND 0.053191f
C4148 VDD.n4034 GND 0.077435f
C4149 VDD.n4035 GND 0.009278f
C4150 VDD.n4036 GND 0.006148f
C4151 VDD.n4037 GND 0.006148f
C4152 VDD.n4038 GND 0.004082f
C4153 VDD.n4039 GND 0.004948f
C4154 VDD.n4040 GND 0.006148f
C4155 VDD.n4041 GND 0.006148f
C4156 VDD.n4042 GND 0.004948f
C4157 VDD.n4043 GND 0.004948f
C4158 VDD.n4044 GND 0.006148f
C4159 VDD.n4045 GND 0.006148f
C4160 VDD.n4046 GND 0.004948f
C4161 VDD.n4047 GND 0.004948f
C4162 VDD.n4048 GND 0.006148f
C4163 VDD.n4049 GND 0.006148f
C4164 VDD.n4050 GND 0.004948f
C4165 VDD.n4051 GND 0.004948f
C4166 VDD.n4052 GND 0.006148f
C4167 VDD.n4053 GND 0.006148f
C4168 VDD.n4054 GND 0.004948f
C4169 VDD.n4055 GND 0.004948f
C4170 VDD.n4056 GND 0.006148f
C4171 VDD.n4057 GND 0.006148f
C4172 VDD.n4058 GND 0.003488f
C4173 VDD.n4059 GND 0.009278f
C4174 VDD.n4060 GND 0.006148f
C4175 VDD.n4061 GND 0.006148f
C4176 VDD.n4062 GND 0.004775f
C4177 VDD.n4063 GND 0.004948f
C4178 VDD.n4064 GND 0.006148f
C4179 VDD.n4065 GND 0.006148f
C4180 VDD.n4066 GND 0.004948f
C4181 VDD.n4067 GND 0.004948f
C4182 VDD.n4068 GND 0.006148f
C4183 VDD.n4069 GND 0.006148f
C4184 VDD.n4070 GND 0.004948f
C4185 VDD.n4071 GND 0.004948f
C4186 VDD.n4072 GND 0.004948f
C4187 VDD.n4073 GND 0.006148f
C4188 VDD.n4074 GND 4.04394f
C4189 VDD.n4076 GND 0.014117f
C4190 VDD.n4077 GND 0.004107f
C4191 VDD.n4078 GND 0.014117f
C4192 VDD.n4079 GND 0.013671f
C4193 VDD.n4080 GND 0.006148f
C4194 VDD.n4081 GND 0.004948f
C4195 VDD.n4082 GND 0.006148f
C4196 VDD.n4083 GND 0.473529f
C4197 VDD.n4084 GND 0.006148f
C4198 VDD.n4085 GND 0.004948f
C4199 VDD.n4086 GND 0.006148f
C4200 VDD.n4087 GND 0.006148f
C4201 VDD.n4088 GND 0.006148f
C4202 VDD.n4089 GND 0.004948f
C4203 VDD.n4090 GND 0.006148f
C4204 VDD.n4091 GND 0.473529f
C4205 VDD.n4092 GND 0.006148f
C4206 VDD.n4093 GND 0.004948f
C4207 VDD.n4094 GND 0.006148f
C4208 VDD.n4095 GND 0.006148f
C4209 VDD.n4096 GND 0.006148f
C4210 VDD.n4097 GND 0.004948f
C4211 VDD.n4098 GND 0.006148f
C4212 VDD.n4099 GND 0.473529f
C4213 VDD.n4100 GND 0.006148f
C4214 VDD.n4101 GND 0.004948f
C4215 VDD.n4102 GND 0.006148f
C4216 VDD.n4103 GND 0.006148f
C4217 VDD.n4104 GND 0.006148f
C4218 VDD.n4105 GND 0.004948f
C4219 VDD.n4106 GND 0.006148f
C4220 VDD.t11 GND 0.473529f
C4221 VDD.n4107 GND 0.006148f
C4222 VDD.n4108 GND 0.004948f
C4223 VDD.n4109 GND 0.006148f
C4224 VDD.n4110 GND 0.006148f
C4225 VDD.n4111 GND 0.006148f
C4226 VDD.n4112 GND 0.004948f
C4227 VDD.n4113 GND 0.006148f
C4228 VDD.n4114 GND 0.473529f
C4229 VDD.n4115 GND 0.006148f
C4230 VDD.n4116 GND 0.004948f
C4231 VDD.n4117 GND 0.006148f
C4232 VDD.n4118 GND 0.006148f
C4233 VDD.n4119 GND 0.006148f
C4234 VDD.n4120 GND 0.004948f
C4235 VDD.n4121 GND 0.006148f
C4236 VDD.n4122 GND 0.473529f
C4237 VDD.n4123 GND 0.006148f
C4238 VDD.n4124 GND 0.004948f
C4239 VDD.n4125 GND 0.006148f
C4240 VDD.n4126 GND 0.006148f
C4241 VDD.n4127 GND 0.006148f
C4242 VDD.n4128 GND 0.004948f
C4243 VDD.n4129 GND 0.006148f
C4244 VDD.n4130 GND 0.473529f
C4245 VDD.n4131 GND 0.006148f
C4246 VDD.n4132 GND 0.004948f
C4247 VDD.n4133 GND 0.006148f
C4248 VDD.n4134 GND 0.006148f
C4249 VDD.n4135 GND 0.006148f
C4250 VDD.n4136 GND 0.004948f
C4251 VDD.n4137 GND 0.006148f
C4252 VDD.n4138 GND 0.473529f
C4253 VDD.n4139 GND 0.006148f
C4254 VDD.n4140 GND 0.004948f
C4255 VDD.n4141 GND 0.006148f
C4256 VDD.n4142 GND 0.006148f
C4257 VDD.n4143 GND 0.006148f
C4258 VDD.n4144 GND 0.004948f
C4259 VDD.n4145 GND 0.006148f
C4260 VDD.n4146 GND 0.473529f
C4261 VDD.n4147 GND 0.006148f
C4262 VDD.n4148 GND 0.004948f
C4263 VDD.n4149 GND 0.006148f
C4264 VDD.n4150 GND 0.006148f
C4265 VDD.n4151 GND 0.006148f
C4266 VDD.n4152 GND 0.004948f
C4267 VDD.n4153 GND 0.006148f
C4268 VDD.n4154 GND 0.473529f
C4269 VDD.n4155 GND 0.006148f
C4270 VDD.n4156 GND 0.004948f
C4271 VDD.n4157 GND 0.006148f
C4272 VDD.n4158 GND 0.006148f
C4273 VDD.n4159 GND 0.006148f
C4274 VDD.n4160 GND 0.004948f
C4275 VDD.n4161 GND 0.006148f
C4276 VDD.n4162 GND 0.473529f
C4277 VDD.n4163 GND 0.006148f
C4278 VDD.n4164 GND 0.004948f
C4279 VDD.n4165 GND 0.006148f
C4280 VDD.n4166 GND 0.006148f
C4281 VDD.n4167 GND 0.006148f
C4282 VDD.n4168 GND 0.006148f
C4283 VDD.n4169 GND 0.006148f
C4284 VDD.n4170 GND 0.004948f
C4285 VDD.n4171 GND 0.006148f
C4286 VDD.n4172 GND 0.473529f
C4287 VDD.n4173 GND 0.006148f
C4288 VDD.n4174 GND 0.006148f
C4289 VDD.n4175 GND 0.006148f
C4290 VDD.n4176 GND 0.006148f
C4291 VDD.n4177 GND 0.004948f
C4292 VDD.n4178 GND 0.006148f
C4293 VDD.n4179 GND 0.006148f
C4294 VDD.n4180 GND 0.006148f
C4295 VDD.n4181 GND 0.006148f
C4296 VDD.n4182 GND 0.473529f
C4297 VDD.n4183 GND 0.006148f
C4298 VDD.n4184 GND 0.006148f
C4299 VDD.n4185 GND 0.006148f
C4300 VDD.n4186 GND 0.006148f
C4301 VDD.n4187 GND 0.006148f
C4302 VDD.n4188 GND 0.004948f
C4303 VDD.n4189 GND 0.006148f
C4304 VDD.n4190 GND 0.006148f
C4305 VDD.n4191 GND 0.006148f
C4306 VDD.n4192 GND 0.006148f
C4307 VDD.n4193 GND 0.473529f
C4308 VDD.n4194 GND 0.006148f
C4309 VDD.n4195 GND 0.006148f
C4310 VDD.n4196 GND 0.006148f
C4311 VDD.n4197 GND 0.006148f
C4312 VDD.n4198 GND 0.006148f
C4313 VDD.n4199 GND 0.004948f
C4314 VDD.n4200 GND 0.006148f
C4315 VDD.n4201 GND 0.006148f
C4316 VDD.n4202 GND 0.006148f
C4317 VDD.n4203 GND 0.006148f
C4318 VDD.n4204 GND 0.473529f
C4319 VDD.n4205 GND 0.006148f
C4320 VDD.n4206 GND 0.006148f
C4321 VDD.n4207 GND 0.006148f
C4322 VDD.n4208 GND 0.006148f
C4323 VDD.n4209 GND 0.006148f
C4324 VDD.n4210 GND 0.004948f
C4325 VDD.n4211 GND 0.006148f
C4326 VDD.n4212 GND 0.473529f
C4327 VDD.n4213 GND 0.006148f
C4328 VDD.n4214 GND 0.006148f
C4329 VDD.n4215 GND 0.004948f
C4330 VDD.n4216 GND 0.006148f
C4331 VDD.n4217 GND 0.006148f
C4332 VDD.n4218 GND 0.004948f
C4333 VDD.n4219 GND 0.006148f
C4334 VDD.n4220 GND 0.006148f
C4335 VDD.n4221 GND 0.004948f
C4336 VDD.n4222 GND 0.006148f
C4337 VDD.n4223 GND 0.006148f
C4338 VDD.n4224 GND 0.006148f
C4339 VDD.n4225 GND 0.004948f
C4340 VDD.n4226 GND 0.004948f
C4341 VDD.n4227 GND 0.004948f
C4342 VDD.n4228 GND 0.006148f
C4343 VDD.n4229 GND 0.006148f
C4344 VDD.n4230 GND 0.006148f
C4345 VDD.n4231 GND 0.004948f
C4346 VDD.n4232 GND 0.004948f
C4347 VDD.n4233 GND 0.004948f
C4348 VDD.n4234 GND 0.006148f
C4349 VDD.n4235 GND 0.006148f
C4350 VDD.n4236 GND 0.006148f
C4351 VDD.n4237 GND 0.004948f
C4352 VDD.n4238 GND 0.004948f
C4353 VDD.n4239 GND 0.004948f
C4354 VDD.n4240 GND 0.006148f
C4355 VDD.n4241 GND 0.006148f
C4356 VDD.n4242 GND 0.006148f
C4357 VDD.n4243 GND 0.006148f
C4358 VDD.n4244 GND 0.006148f
C4359 VDD.n4245 GND 0.004948f
C4360 VDD.n4246 GND 0.006148f
C4361 VDD.n4247 GND 0.473529f
C4362 VDD.n4248 GND 0.006148f
C4363 VDD.n4249 GND 0.006148f
C4364 VDD.n4250 GND 0.006148f
C4365 VDD.n4251 GND 0.006148f
C4366 VDD.n4252 GND 0.006148f
C4367 VDD.n4253 GND 0.004948f
C4368 VDD.n4254 GND 0.006148f
C4369 VDD.n4255 GND 0.006148f
C4370 VDD.n4256 GND 0.006148f
C4371 VDD.n4257 GND 0.006148f
C4372 VDD.n4258 GND 0.670043f
C4373 VDD.n4259 GND 0.013671f
C4374 VDD.n4260 GND 0.006148f
C4375 VDD.n4261 GND 0.006148f
C4376 VDD.n4262 GND 0.006148f
C4377 VDD.n4263 GND 0.004948f
C4378 VDD.n4264 GND 1.09148f
C4379 VDD.n4265 GND 0.004948f
C4380 VDD.n4266 GND 0.006148f
C4381 VDD.n4267 GND 0.006148f
C4382 VDD.n4268 GND 0.006148f
C4383 VDD.n4269 GND 0.006148f
C4384 VDD.n4270 GND 0.006148f
C4385 VDD.n4271 GND 0.004948f
C4386 VDD.n4273 GND 0.006148f
C4387 VDD.n4274 GND 0.006148f
C4388 VDD.n4275 GND 0.006148f
C4389 VDD.n4276 GND 0.006148f
C4390 VDD.n4277 GND 0.003488f
C4391 VDD.t66 GND 0.085164f
C4392 VDD.t65 GND 0.430073f
C4393 VDD.n4278 GND 0.075426f
C4394 VDD.t67 GND 0.053191f
C4395 VDD.n4279 GND 0.077435f
C4396 VDD.n4281 GND 0.006148f
C4397 VDD.n4282 GND 0.006148f
C4398 VDD.n4283 GND 0.004948f
C4399 VDD.n4284 GND 0.006148f
C4400 VDD.n4286 GND 0.006148f
C4401 VDD.n4287 GND 0.006148f
C4402 VDD.n4288 GND 0.006148f
C4403 VDD.n4289 GND 0.006148f
C4404 VDD.n4290 GND 0.004948f
C4405 VDD.n4292 GND 0.006148f
C4406 VDD.n4293 GND 0.006148f
C4407 VDD.n4294 GND 0.006148f
C4408 VDD.n4295 GND 0.006148f
C4409 VDD.n4296 GND 0.006148f
C4410 VDD.n4297 GND 0.004082f
C4411 VDD.n4299 GND 0.006148f
C4412 VDD.n4300 GND 0.004181f
C4413 VDD.t60 GND 0.085164f
C4414 VDD.t59 GND 0.430073f
C4415 VDD.n4301 GND 0.075426f
C4416 VDD.t61 GND 0.053191f
C4417 VDD.n4302 GND 0.077435f
C4418 VDD.n4303 GND 0.006148f
C4419 VDD.n4304 GND 0.006148f
C4420 VDD.n4305 GND 0.004948f
C4421 VDD.n4307 GND 0.006148f
C4422 VDD.n4308 GND 0.006148f
C4423 VDD.n4309 GND 0.006148f
C4424 VDD.n4310 GND 0.006148f
C4425 VDD.n4311 GND 0.004948f
C4426 VDD.n4313 GND 0.006148f
C4427 VDD.n4314 GND 0.006148f
C4428 VDD.n4315 GND 0.006148f
C4429 VDD.n4316 GND 0.006148f
C4430 VDD.n4317 GND 0.006148f
C4431 VDD.n4318 GND 0.00339f
C4432 VDD.n4320 GND 0.006148f
C4433 VDD.n4321 GND 0.004874f
C4434 VDD.t54 GND 0.085164f
C4435 VDD.t53 GND 0.430073f
C4436 VDD.n4322 GND 0.075426f
C4437 VDD.t55 GND 0.053191f
C4438 VDD.n4323 GND 0.077435f
C4439 VDD.n4324 GND 0.006148f
C4440 VDD.n4325 GND 0.006148f
C4441 VDD.n4326 GND 0.004948f
C4442 VDD.n4328 GND 0.006148f
C4443 VDD.n4329 GND 0.006148f
C4444 VDD.n4330 GND 0.006148f
C4445 VDD.n4331 GND 0.006148f
C4446 VDD.n4332 GND 0.004948f
C4447 VDD.n4334 GND 0.006148f
C4448 VDD.n4335 GND 0.006148f
C4449 VDD.n4336 GND 0.006148f
C4450 VDD.n4337 GND 0.006148f
C4451 VDD.n4338 GND 0.006148f
C4452 VDD.n4339 GND 0.002697f
C4453 VDD.n4341 GND 0.006148f
C4454 VDD.t87 GND 0.085164f
C4455 VDD.t86 GND 0.430073f
C4456 VDD.n4342 GND 0.075426f
C4457 VDD.t88 GND 0.053191f
C4458 VDD.n4343 GND 0.077435f
C4459 VDD.n4344 GND 0.006804f
C4460 VDD.n4345 GND 0.006148f
C4461 VDD.n4346 GND 0.006148f
C4462 VDD.n4347 GND 0.006148f
C4463 VDD.n4348 GND 0.006148f
C4464 VDD.n4349 GND 0.004948f
C4465 VDD.n4351 GND 0.006148f
C4466 VDD.n4352 GND 0.006148f
C4467 VDD.n4353 GND 0.006148f
C4468 VDD.n4354 GND 0.006148f
C4469 VDD.n4355 GND 0.006148f
C4470 VDD.n4356 GND 0.004948f
C4471 VDD.n4358 GND 0.006148f
C4472 VDD.n4359 GND 0.006148f
C4473 VDD.n4360 GND 0.006148f
C4474 VDD.n4361 GND 0.006148f
C4475 VDD.n4362 GND 0.006148f
C4476 VDD.t44 GND 0.085164f
C4477 VDD.t42 GND 0.430073f
C4478 VDD.n4363 GND 0.075426f
C4479 VDD.t45 GND 0.053191f
C4480 VDD.n4364 GND 0.077435f
C4481 VDD.n4365 GND 0.009278f
C4482 VDD.n4367 GND 0.013671f
C4483 VDD.n4368 GND 0.006148f
C4484 VDD.n4369 GND 0.006148f
C4485 VDD.n4370 GND 0.004948f
C4486 VDD.n4371 GND 0.006148f
C4487 VDD.n4372 GND 0.006148f
C4488 VDD.n4373 GND 0.006148f
C4489 VDD.n4374 GND 0.004948f
C4490 VDD.n4375 GND 0.004948f
C4491 VDD.n4376 GND 0.004107f
C4492 VDD.n4377 GND 0.013671f
C4493 VDD.n4378 GND 0.014117f
C4494 VDD.n4379 GND 0.002944f
C4495 VDD.n4380 GND 0.014117f
C4496 VDD.n4382 GND 0.006148f
C4497 VDD.n4383 GND 0.006148f
C4498 VDD.n4384 GND 0.004478f
C4499 VDD.n4385 GND 0.004948f
C4500 VDD.n4386 GND 0.004948f
C4501 VDD.n4387 GND 0.006148f
C4502 VDD.n4389 GND 0.006148f
C4503 VDD.n4390 GND 0.006148f
C4504 VDD.n4391 GND 0.004948f
C4505 VDD.n4392 GND 0.004948f
C4506 VDD.n4393 GND 0.004948f
C4507 VDD.n4394 GND 0.006148f
C4508 VDD.n4396 GND 0.006148f
C4509 VDD.n4397 GND 0.006148f
C4510 VDD.n4398 GND 0.004948f
C4511 VDD.n4399 GND 0.004948f
C4512 VDD.n4400 GND 0.003093f
C4513 VDD.n4401 GND 0.006148f
C4514 VDD.n4403 GND 0.006148f
C4515 VDD.n4404 GND 0.006148f
C4516 VDD.n4405 GND 0.004948f
C4517 VDD.n4406 GND 0.004948f
C4518 VDD.n4407 GND 0.004948f
C4519 VDD.n4408 GND 0.006148f
C4520 VDD.n4410 GND 0.006148f
C4521 VDD.n4411 GND 0.006148f
C4522 VDD.n4412 GND 0.004948f
C4523 VDD.n4413 GND 0.004948f
C4524 VDD.n4414 GND 0.004948f
C4525 VDD.n4415 GND 0.006148f
C4526 VDD.n4417 GND 0.006148f
C4527 VDD.n4418 GND 0.006148f
C4528 VDD.n4419 GND 0.004948f
C4529 VDD.n4420 GND 0.006148f
C4530 VDD.n4421 GND 0.006148f
C4531 VDD.n4422 GND 0.006148f
C4532 VDD.n4423 GND 0.009278f
C4533 VDD.n4424 GND 0.006148f
C4534 VDD.n4426 GND 0.006148f
C4535 VDD.n4427 GND 0.006148f
C4536 VDD.n4428 GND 0.004948f
C4537 VDD.n4429 GND 0.004948f
C4538 VDD.n4430 GND 0.004948f
C4539 VDD.n4431 GND 0.006148f
C4540 VDD.n4433 GND 0.006148f
C4541 VDD.n4434 GND 0.006148f
C4542 VDD.n4435 GND 0.004948f
C4543 VDD.n4436 GND 0.004948f
C4544 VDD.n4437 GND 0.004948f
C4545 VDD.n4438 GND 0.006148f
C4546 VDD.n4440 GND 0.006148f
C4547 VDD.n4441 GND 0.006148f
C4548 VDD.n4442 GND 0.004948f
C4549 VDD.n4443 GND 0.006148f
C4550 VDD.n4444 GND 0.006148f
C4551 VDD.n4445 GND 0.006148f
C4552 VDD.n4446 GND 0.009278f
C4553 VDD.n4447 GND 0.006148f
C4554 VDD.n4449 GND 0.006148f
C4555 VDD.n4450 GND 0.006148f
C4556 VDD.n4451 GND 0.004948f
C4557 VDD.n4452 GND 0.004948f
C4558 VDD.n4453 GND 0.004948f
C4559 VDD.n4454 GND 0.006148f
C4560 VDD.n4456 GND 0.006148f
C4561 VDD.n4457 GND 0.006148f
C4562 VDD.n4458 GND 0.004948f
C4563 VDD.n4459 GND 0.004948f
C4564 VDD.n4460 GND 0.004948f
C4565 VDD.n4461 GND 0.006148f
C4566 VDD.n4463 GND 0.006148f
C4567 VDD.n4464 GND 0.006148f
C4568 VDD.n4465 GND 0.004948f
C4569 VDD.n4466 GND 0.006148f
C4570 VDD.n4467 GND 0.006148f
C4571 VDD.n4468 GND 0.006148f
C4572 VDD.n4469 GND 0.009278f
C4573 VDD.n4470 GND 0.004775f
C4574 VDD.n4471 GND 0.004948f
C4575 VDD.n4472 GND 0.006148f
C4576 VDD.n4474 GND 0.006148f
C4577 VDD.n4475 GND 0.006148f
C4578 VDD.n4476 GND 0.004948f
C4579 VDD.n4477 GND 0.004948f
C4580 VDD.n4478 GND 0.004948f
C4581 VDD.n4479 GND 0.006148f
C4582 VDD.n4481 GND 0.006148f
C4583 VDD.n4482 GND 0.006148f
C4584 VDD.n4484 GND 0.014117f
C4585 VDD.n4485 GND 0.004107f
C4586 VDD.n4486 GND 0.014117f
C4587 VDD.n4487 GND 0.013671f
C4588 VDD.n4488 GND 0.004107f
C4589 VDD.n4489 GND 0.004948f
C4590 VDD.n4490 GND 0.006148f
C4591 VDD.n4491 GND 0.473529f
C4592 VDD.n4492 GND 0.473529f
C4593 VDD.n4493 GND 0.473529f
C4594 VDD.n4494 GND 0.006148f
C4595 VDD.n4495 GND 0.004948f
C4596 VDD.n4496 GND 0.004948f
C4597 VDD.n4497 GND 0.004948f
C4598 VDD.n4498 GND 0.006148f
C4599 VDD.n4499 GND 0.473529f
C4600 VDD.n4500 GND 0.006148f
C4601 VDD.n4501 GND 0.004948f
C4602 VDD.n4502 GND 0.004948f
C4603 VDD.n4503 GND 0.004948f
C4604 VDD.n4504 GND 0.006148f
C4605 VDD.t43 GND 0.473529f
C4606 VDD.n4505 GND 0.006148f
C4607 VDD.n4506 GND 0.004948f
C4608 VDD.n4507 GND 0.004948f
C4609 VDD.n4508 GND 0.004948f
C4610 VDD.n4509 GND 0.006148f
C4611 VDD.n4510 GND 0.473529f
C4612 VDD.n4511 GND 0.473529f
C4613 VDD.n4512 GND 0.473529f
C4614 VDD.n4513 GND 0.006148f
C4615 VDD.n4514 GND 0.004948f
C4616 VDD.n4515 GND 0.004948f
C4617 VDD.n4516 GND 0.004948f
C4618 VDD.n4517 GND 0.006148f
C4619 VDD.n4518 GND 0.473529f
C4620 VDD.n4519 GND 0.473529f
C4621 VDD.n4520 GND 0.473529f
C4622 VDD.n4521 GND 0.006148f
C4623 VDD.n4522 GND 0.004948f
C4624 VDD.n4523 GND 0.004948f
C4625 VDD.n4524 GND 0.004948f
C4626 VDD.n4525 GND 0.006148f
C4627 VDD.n4526 GND 0.473529f
C4628 VDD.n4527 GND 0.473529f
C4629 VDD.n4528 GND 0.473529f
C4630 VDD.n4529 GND 0.006148f
C4631 VDD.n4530 GND 0.004948f
C4632 VDD.n4531 GND 0.004948f
C4633 VDD.n4532 GND 0.004948f
C4634 VDD.n4533 GND 0.006148f
C4635 VDD.n4534 GND 0.473529f
C4636 VDD.n4535 GND 0.006148f
C4637 VDD.n4536 GND 0.004948f
C4638 VDD.n4537 GND 0.004948f
C4639 VDD.n4538 GND 0.004948f
C4640 VDD.n4539 GND 0.006148f
C4641 VDD.t137 GND 0.473529f
C4642 VDD.n4540 GND 0.006148f
C4643 VDD.n4541 GND 0.004948f
C4644 VDD.n4542 GND 0.136126f
C4645 VDD.n4543 GND 2.23369f
C4646 a_n11778_11043.n0 GND 8.1951f
C4647 a_n11778_11043.n1 GND 5.822741f
C4648 a_n11778_11043.n2 GND 10.6975f
C4649 a_n11778_11043.n3 GND 23.8866f
C4650 a_n11778_11043.t3 GND 0.084679f
C4651 a_n11778_11043.t7 GND 0.519037f
C4652 a_n11778_11043.t9 GND 0.084679f
C4653 a_n11778_11043.t11 GND 0.084679f
C4654 a_n11778_11043.n4 GND 0.371451f
C4655 a_n11778_11043.t8 GND 0.515678f
C4656 a_n11778_11043.t10 GND 0.084679f
C4657 a_n11778_11043.t4 GND 0.084679f
C4658 a_n11778_11043.n5 GND 0.371451f
C4659 a_n11778_11043.t6 GND 0.084679f
C4660 a_n11778_11043.t5 GND 0.084679f
C4661 a_n11778_11043.n6 GND 0.371451f
C4662 a_n11778_11043.t13 GND 0.449343f
C4663 a_n11778_11043.t1 GND 0.084679f
C4664 a_n11778_11043.t17 GND 0.084679f
C4665 a_n11778_11043.n7 GND 0.29696f
C4666 a_n11778_11043.t16 GND 0.429493f
C4667 a_n11778_11043.t0 GND 0.429493f
C4668 a_n11778_11043.t15 GND 0.084679f
C4669 a_n11778_11043.t2 GND 0.084679f
C4670 a_n11778_11043.n8 GND 0.29696f
C4671 a_n11778_11043.t14 GND 0.429493f
C4672 a_n11778_11043.n9 GND 6.62972f
C4673 a_n11778_11043.n10 GND 0.371451f
C4674 a_n11778_11043.t12 GND 0.084679f
C4675 a_n11634_10845.n0 GND 2.63336f
C4676 a_n11634_10845.n1 GND 0.781531f
C4677 a_n11634_10845.n2 GND 0.741219f
C4678 a_n11634_10845.n3 GND 2.5623f
C4679 a_n11634_10845.n4 GND 0.898863f
C4680 a_n11634_10845.n5 GND 0.741219f
C4681 a_n11634_10845.n6 GND 2.6261f
C4682 a_n11634_10845.n7 GND 0.781531f
C4683 a_n11634_10845.n8 GND 0.741219f
C4684 a_n11634_10845.n9 GND 4.33195f
C4685 a_n11634_10845.n10 GND 0.745268f
C4686 a_n11634_10845.n11 GND 0.745323f
C4687 a_n11634_10845.n12 GND 0.745323f
C4688 a_n11634_10845.n13 GND 0.745323f
C4689 a_n11634_10845.n14 GND 1.77899f
C4690 a_n11634_10845.n15 GND 0.745592f
C4691 a_n11634_10845.n16 GND 0.737552f
C4692 a_n11634_10845.n17 GND 0.941867f
C4693 a_n11634_10845.n18 GND 0.154323f
C4694 a_n11634_10845.n19 GND 0.519444f
C4695 a_n11634_10845.n20 GND 0.894419f
C4696 a_n11634_10845.n21 GND 0.145734f
C4697 a_n11634_10845.n22 GND 0.154323f
C4698 a_n11634_10845.n23 GND 0.233664f
C4699 a_n11634_10845.n24 GND 0.128061f
C4700 a_n11634_10845.n25 GND 0.216253f
C4701 a_n11634_10845.n26 GND 1.24679f
C4702 a_n11634_10845.n27 GND 0.205222f
C4703 a_n11634_10845.n28 GND 0.233647f
C4704 a_n11634_10845.n29 GND 0.154323f
C4705 a_n11634_10845.n30 GND 0.203044f
C4706 a_n11634_10845.n31 GND 0.154323f
C4707 a_n11634_10845.n32 GND 0.236952f
C4708 a_n11634_10845.n33 GND 0.154323f
C4709 a_n11634_10845.n34 GND 0.203556f
C4710 a_n11634_10845.n35 GND 0.154323f
C4711 a_n11634_10845.n36 GND 0.196824f
C4712 a_n11634_10845.n37 GND 0.154323f
C4713 a_n11634_10845.n38 GND 0.245908f
C4714 a_n11634_10845.n39 GND 0.154323f
C4715 a_n11634_10845.n40 GND 0.154323f
C4716 a_n11634_10845.n41 GND 0.213214f
C4717 a_n11634_10845.n42 GND 0.154323f
C4718 a_n11634_10845.n43 GND 0.215228f
C4719 a_n11634_10845.n44 GND 0.154323f
C4720 a_n11634_10845.n45 GND 0.154323f
C4721 a_n11634_10845.n46 GND 0.24523f
C4722 a_n11634_10845.n47 GND 0.154323f
C4723 a_n11634_10845.n48 GND 0.198013f
C4724 a_n11634_10845.n49 GND 0.166642f
C4725 a_n11634_10845.n50 GND 0.201314f
C4726 a_n11634_10845.n51 GND 1.13455f
C4727 a_n11634_10845.n52 GND 0.205222f
C4728 a_n11634_10845.n53 GND 0.233647f
C4729 a_n11634_10845.n54 GND 0.154323f
C4730 a_n11634_10845.n55 GND 0.203044f
C4731 a_n11634_10845.n56 GND 0.154323f
C4732 a_n11634_10845.n57 GND 0.236952f
C4733 a_n11634_10845.n58 GND 0.154323f
C4734 a_n11634_10845.n59 GND 0.203556f
C4735 a_n11634_10845.n60 GND 0.154323f
C4736 a_n11634_10845.n61 GND 0.196824f
C4737 a_n11634_10845.n62 GND 0.154323f
C4738 a_n11634_10845.n63 GND 0.245908f
C4739 a_n11634_10845.n64 GND 0.154323f
C4740 a_n11634_10845.n65 GND 0.154323f
C4741 a_n11634_10845.n66 GND 0.213214f
C4742 a_n11634_10845.n67 GND 0.154323f
C4743 a_n11634_10845.n68 GND 0.215228f
C4744 a_n11634_10845.n69 GND 0.154323f
C4745 a_n11634_10845.n70 GND 0.154323f
C4746 a_n11634_10845.n71 GND 0.24523f
C4747 a_n11634_10845.n72 GND 0.154323f
C4748 a_n11634_10845.n73 GND 0.198013f
C4749 a_n11634_10845.n74 GND 0.166642f
C4750 a_n11634_10845.n75 GND 0.201314f
C4751 a_n11634_10845.n76 GND 0.952463f
C4752 a_n11634_10845.n77 GND 0.205222f
C4753 a_n11634_10845.n78 GND 0.233647f
C4754 a_n11634_10845.n79 GND 0.154323f
C4755 a_n11634_10845.n80 GND 0.203044f
C4756 a_n11634_10845.n81 GND 0.154323f
C4757 a_n11634_10845.n82 GND 0.236952f
C4758 a_n11634_10845.n83 GND 0.154323f
C4759 a_n11634_10845.n84 GND 0.203556f
C4760 a_n11634_10845.n85 GND 0.154323f
C4761 a_n11634_10845.n86 GND 0.196824f
C4762 a_n11634_10845.n87 GND 0.154323f
C4763 a_n11634_10845.n88 GND 0.245908f
C4764 a_n11634_10845.n89 GND 0.154323f
C4765 a_n11634_10845.n90 GND 0.154323f
C4766 a_n11634_10845.n91 GND 0.213214f
C4767 a_n11634_10845.n92 GND 0.154323f
C4768 a_n11634_10845.n93 GND 0.215228f
C4769 a_n11634_10845.n94 GND 0.154323f
C4770 a_n11634_10845.n95 GND 0.154323f
C4771 a_n11634_10845.n96 GND 0.24523f
C4772 a_n11634_10845.n97 GND 0.154323f
C4773 a_n11634_10845.n98 GND 0.198013f
C4774 a_n11634_10845.n99 GND 0.166642f
C4775 a_n11634_10845.n100 GND 0.201314f
C4776 a_n11634_10845.n101 GND 0.115132f
C4777 a_n11634_10845.n102 GND 0.163032f
C4778 a_n11634_10845.n103 GND 0.165436f
C4779 a_n11634_10845.n104 GND 0.11212f
C4780 a_n11634_10845.n105 GND 0.115132f
C4781 a_n11634_10845.n106 GND 0.163032f
C4782 a_n11634_10845.n107 GND 0.165436f
C4783 a_n11634_10845.n108 GND 0.11212f
C4784 a_n11634_10845.n109 GND 0.115132f
C4785 a_n11634_10845.n110 GND 0.163032f
C4786 a_n11634_10845.n111 GND 0.165436f
C4787 a_n11634_10845.n112 GND 0.11212f
C4788 a_n11634_10845.n113 GND 0.711626f
C4789 a_n11634_10845.n114 GND 0.161808f
C4790 a_n11634_10845.t38 GND 1.40117f
C4791 a_n11634_10845.t41 GND 1.40117f
C4792 a_n11634_10845.t46 GND 1.40117f
C4793 a_n11634_10845.t34 GND 1.40117f
C4794 a_n11634_10845.n115 GND 0.617205f
C4795 a_n11634_10845.t20 GND 0.060894f
C4796 a_n11634_10845.t8 GND 0.060894f
C4797 a_n11634_10845.n116 GND 0.241413f
C4798 a_n11634_10845.t6 GND 0.060894f
C4799 a_n11634_10845.t18 GND 0.060894f
C4800 a_n11634_10845.n117 GND 0.213548f
C4801 a_n11634_10845.n118 GND 3.88546f
C4802 a_n11634_10845.t4 GND 0.308853f
C4803 a_n11634_10845.n119 GND 3.64128f
C4804 a_n11634_10845.n120 GND 1.37723f
C4805 a_n11634_10845.t42 GND 2.07467f
C4806 a_n11634_10845.t43 GND 1.40117f
C4807 a_n11634_10845.t27 GND 2.05279f
C4808 a_n11634_10845.t37 GND 2.07142f
C4809 a_n11634_10845.t22 GND 2.07467f
C4810 a_n11634_10845.t24 GND 1.40117f
C4811 a_n11634_10845.t45 GND 2.05279f
C4812 a_n11634_10845.t25 GND 2.07142f
C4813 a_n11634_10845.t26 GND 2.07467f
C4814 a_n11634_10845.t44 GND 1.40117f
C4815 a_n11634_10845.t23 GND 2.05279f
C4816 a_n11634_10845.t47 GND 2.07142f
C4817 a_n11634_10845.t36 GND 2.07271f
C4818 a_n11634_10845.t40 GND 1.40117f
C4819 a_n11634_10845.t33 GND 1.40117f
C4820 a_n11634_10845.t39 GND 1.40117f
C4821 a_n11634_10845.n121 GND 0.781702f
C4822 a_n11634_10845.t28 GND 1.40117f
C4823 a_n11634_10845.t32 GND 1.40117f
C4824 a_n11634_10845.t30 GND 1.40117f
C4825 a_n11634_10845.t35 GND 1.40117f
C4826 a_n11634_10845.n122 GND 0.617205f
C4827 a_n11634_10845.t19 GND 1.40117f
C4828 a_n11634_10845.t7 GND 1.40117f
C4829 a_n11634_10845.t5 GND 1.40117f
C4830 a_n11634_10845.t17 GND 1.40117f
C4831 a_n11634_10845.n123 GND 0.617205f
C4832 a_n11634_10845.t3 GND 1.40117f
C4833 a_n11634_10845.n124 GND 0.821535f
C4834 a_n11634_10845.n125 GND 0.101565f
C4835 a_n11634_10845.n126 GND 0.632175f
C4836 a_n11634_10845.n127 GND 0.630769f
C4837 a_n11634_10845.n128 GND 0.802054f
C4838 a_n11634_10845.n129 GND 0.952463f
C4839 a_n11634_10845.t29 GND 1.40117f
C4840 a_n11634_10845.n130 GND 0.821535f
C4841 a_n11634_10845.n131 GND 0.101565f
C4842 a_n11634_10845.n132 GND 0.632175f
C4843 a_n11634_10845.n133 GND 0.630769f
C4844 a_n11634_10845.n134 GND 0.802054f
C4845 a_n11634_10845.n135 GND 1.26446f
C4846 a_n11634_10845.t11 GND 2.10019f
C4847 a_n11634_10845.t13 GND 2.07098f
C4848 a_n11634_10845.t15 GND 2.06556f
C4849 a_n11634_10845.t9 GND 1.40117f
C4850 a_n11634_10845.n136 GND 0.901537f
C4851 a_n11634_10845.t1 GND 2.07443f
C4852 a_n11634_10845.t2 GND 0.323128f
C4853 a_n11634_10845.t16 GND 0.060894f
C4854 a_n11634_10845.t10 GND 0.060894f
C4855 a_n11634_10845.n137 GND 0.213548f
C4856 a_n11634_10845.n138 GND 3.13495f
C4857 a_n11634_10845.t12 GND 0.060894f
C4858 a_n11634_10845.t14 GND 0.060894f
C4859 a_n11634_10845.n139 GND 0.213548f
C4860 a_n11634_10845.n140 GND 4.00004f
C4861 a_n11634_10845.n141 GND 1.62044f
C4862 a_n11634_10845.n142 GND 1.00416f
C4863 a_n11634_10845.n143 GND 0.774188f
C4864 a_n11634_10845.n144 GND 0.90535f
C4865 a_n11634_10845.n145 GND 0.90535f
C4866 a_n11634_10845.n146 GND 0.90535f
C4867 a_n11634_10845.n147 GND 1.08331f
C4868 a_n11634_10845.t31 GND 1.40117f
C4869 a_n11634_10845.n148 GND 0.821535f
C4870 a_n11634_10845.n149 GND 0.101565f
C4871 a_n11634_10845.n150 GND 0.632175f
C4872 a_n11634_10845.n151 GND 0.630769f
C4873 a_n11634_10845.n152 GND 0.802054f
C4874 a_n11634_10845.n153 GND 0.670294f
C4875 a_n11634_10845.n154 GND 2.91651f
C4876 a_n11634_10845.t21 GND 1.49956f
C4877 a_n11634_10845.n155 GND 6.6241f
C4878 a_n11634_10845.t0 GND 2.19692f
C4879 VN.t7 GND 0.72163f
C4880 VN.t8 GND 0.797313f
C4881 VN.n0 GND 1.40982f
C4882 VN.t0 GND 0.02223f
C4883 VN.t1 GND 0.00397f
C4884 VN.t4 GND 0.00397f
C4885 VN.n1 GND 0.012875f
C4886 VN.n2 GND 0.099946f
C4887 VN.t2 GND 0.00397f
C4888 VN.t6 GND 0.00397f
C4889 VN.n3 GND 0.012875f
C4890 VN.n4 GND 0.054017f
C4891 VN.t3 GND 0.00397f
C4892 VN.t5 GND 0.00397f
C4893 VN.n5 GND 0.012875f
C4894 VN.n6 GND 0.075021f
C4895 VN.n7 GND 2.53743f
C4896 VOUT.t21 GND 0.151585f
C4897 VOUT.t16 GND 0.148129f
C4898 VOUT.n0 GND 1.60866f
C4899 VOUT.t20 GND 0.148129f
C4900 VOUT.n1 GND 0.872357f
C4901 VOUT.t22 GND 0.148129f
C4902 VOUT.n2 GND 0.872357f
C4903 VOUT.t23 GND 0.148129f
C4904 VOUT.n3 GND 1.10744f
C4905 VOUT.n4 GND 9.12822f
C4906 VOUT.t27 GND 14.550901f
C4907 VOUT.t26 GND 9.06784f
C4908 VOUT.n5 GND 10.1378f
C4909 VOUT.n6 GND 1.95321f
C4910 VOUT.t24 GND 0.153182f
C4911 VOUT.t19 GND 0.149752f
C4912 VOUT.n7 GND 1.60544f
C4913 VOUT.t25 GND 0.149752f
C4914 VOUT.n8 GND 0.870734f
C4915 VOUT.t17 GND 0.149752f
C4916 VOUT.n9 GND 0.870734f
C4917 VOUT.t18 GND 0.149751f
C4918 VOUT.n10 GND 1.10581f
C4919 VOUT.n11 GND 11.733299f
C4920 VOUT.t14 GND 0.054741f
C4921 VOUT.t1 GND 0.054741f
C4922 VOUT.n12 GND 0.461237f
C4923 VOUT.t11 GND 0.054741f
C4924 VOUT.t2 GND 0.054741f
C4925 VOUT.n13 GND 0.443815f
C4926 VOUT.n14 GND 1.99188f
C4927 VOUT.t4 GND 0.054741f
C4928 VOUT.t10 GND 0.054741f
C4929 VOUT.n15 GND 0.443815f
C4930 VOUT.n16 GND 1.11344f
C4931 VOUT.t12 GND 0.054741f
C4932 VOUT.t3 GND 0.054741f
C4933 VOUT.n17 GND 0.443815f
C4934 VOUT.n18 GND 1.22704f
C4935 VOUT.n19 GND 10.819f
C4936 VOUT.t5 GND 0.054741f
C4937 VOUT.t6 GND 0.054741f
C4938 VOUT.n20 GND 0.461237f
C4939 VOUT.t8 GND 0.054741f
C4940 VOUT.t13 GND 0.054741f
C4941 VOUT.n21 GND 0.443815f
C4942 VOUT.n22 GND 1.99188f
C4943 VOUT.t0 GND 0.054741f
C4944 VOUT.t7 GND 0.054741f
C4945 VOUT.n23 GND 0.443815f
C4946 VOUT.n24 GND 1.11344f
C4947 VOUT.t9 GND 0.054741f
C4948 VOUT.t15 GND 0.054741f
C4949 VOUT.n25 GND 0.443815f
C4950 VOUT.n26 GND 1.22704f
C4951 VOUT.n27 GND 8.08887f
C4952 VOUT.n28 GND 5.415411f
C4953 CS_BIAS.n0 GND 0.01048f
C4954 CS_BIAS.t9 GND 0.380517f
C4955 CS_BIAS.n1 GND 0.010384f
C4956 CS_BIAS.n2 GND 0.004867f
C4957 CS_BIAS.t22 GND 0.457855f
C4958 CS_BIAS.t0 GND 0.473155f
C4959 CS_BIAS.t2 GND 0.477977f
C4960 CS_BIAS.n3 GND 0.412925f
C4961 CS_BIAS.t1 GND 0.020302f
C4962 CS_BIAS.t3 GND 0.020302f
C4963 CS_BIAS.n4 GND 0.144034f
C4964 CS_BIAS.n5 GND 0.307233f
C4965 CS_BIAS.n6 GND 0.10353f
C4966 CS_BIAS.n7 GND 0.12723f
C4967 CS_BIAS.n8 GND 0.011244f
C4968 CS_BIAS.n9 GND 0.011224f
C4969 CS_BIAS.n10 GND 0.005572f
C4970 CS_BIAS.n11 GND 0.005572f
C4971 CS_BIAS.n12 GND 0.005572f
C4972 CS_BIAS.n13 GND 0.010384f
C4973 CS_BIAS.n14 GND 0.007974f
C4974 CS_BIAS.n15 GND 0.163111f
C4975 CS_BIAS.n16 GND 0.058356f
C4976 CS_BIAS.t12 GND 0.473155f
C4977 CS_BIAS.t21 GND 0.477977f
C4978 CS_BIAS.n17 GND 0.359136f
C4979 CS_BIAS.n18 GND 0.10397f
C4980 CS_BIAS.t19 GND 0.473155f
C4981 CS_BIAS.t13 GND 0.477977f
C4982 CS_BIAS.n19 GND 0.359136f
C4983 CS_BIAS.n20 GND 0.081791f
C4984 CS_BIAS.t20 GND 0.477977f
C4985 CS_BIAS.t11 GND 0.473155f
C4986 CS_BIAS.n21 GND 0.359135f
C4987 CS_BIAS.n22 GND 0.587844f
C4988 CS_BIAS.n23 GND 0.01048f
C4989 CS_BIAS.t17 GND 0.380517f
C4990 CS_BIAS.n24 GND 0.010384f
C4991 CS_BIAS.n25 GND 0.004867f
C4992 CS_BIAS.t18 GND 0.457856f
C4993 CS_BIAS.t5 GND 0.020302f
C4994 CS_BIAS.t7 GND 0.020302f
C4995 CS_BIAS.n26 GND 0.144034f
C4996 CS_BIAS.t4 GND 0.477977f
C4997 CS_BIAS.t6 GND 0.473155f
C4998 CS_BIAS.n27 GND 0.412924f
C4999 CS_BIAS.n28 GND 0.307233f
C5000 CS_BIAS.n29 GND 0.103529f
C5001 CS_BIAS.n30 GND 0.12723f
C5002 CS_BIAS.n31 GND 0.011244f
C5003 CS_BIAS.n32 GND 0.011224f
C5004 CS_BIAS.n33 GND 0.005572f
C5005 CS_BIAS.n34 GND 0.005572f
C5006 CS_BIAS.n35 GND 0.005572f
C5007 CS_BIAS.n36 GND 0.010384f
C5008 CS_BIAS.n37 GND 0.007974f
C5009 CS_BIAS.n38 GND 0.163111f
C5010 CS_BIAS.n39 GND 0.058356f
C5011 CS_BIAS.t15 GND 0.477977f
C5012 CS_BIAS.t10 GND 0.473155f
C5013 CS_BIAS.n40 GND 0.359135f
C5014 CS_BIAS.n41 GND 0.10397f
C5015 CS_BIAS.t23 GND 0.477977f
C5016 CS_BIAS.t16 GND 0.473155f
C5017 CS_BIAS.n42 GND 0.359135f
C5018 CS_BIAS.n43 GND 0.081791f
C5019 CS_BIAS.t14 GND 0.477977f
C5020 CS_BIAS.t8 GND 0.473155f
C5021 CS_BIAS.n44 GND 0.359135f
C5022 CS_BIAS.n45 GND 0.126031f
C5023 CS_BIAS.n46 GND 4.56507f
.ends

