* NGSPICE file created from diff_pair_sample_1470.ext - technology: sky130A

.subckt diff_pair_sample_1470 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X1 VTAIL.t4 VP.t0 VDD1.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X2 VDD2.t2 VN.t1 VTAIL.t18 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0.9207 ps=5.91 w=5.58 l=1.84
X3 VDD1.t8 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X4 VTAIL.t17 VN.t2 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X5 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0 ps=0 w=5.58 l=1.84
X6 VDD2.t8 VN.t3 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0 ps=0 w=5.58 l=1.84
X8 VTAIL.t3 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X9 VDD1.t6 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0.9207 ps=5.91 w=5.58 l=1.84
X10 VTAIL.t15 VN.t4 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X11 VDD2.t5 VN.t5 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X12 VTAIL.t7 VP.t4 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X13 VTAIL.t13 VN.t6 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X14 VDD1.t4 VP.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=2.1762 ps=11.94 w=5.58 l=1.84
X15 VDD1.t3 VP.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=2.1762 ps=11.94 w=5.58 l=1.84
X16 VDD2.t3 VN.t7 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=2.1762 ps=11.94 w=5.58 l=1.84
X17 VTAIL.t9 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X18 VDD2.t7 VN.t8 VTAIL.t11 B.t8 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=2.1762 ps=11.94 w=5.58 l=1.84
X19 VDD1.t1 VP.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0.9207 ps=5.91 w=5.58 l=1.84
X20 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0 ps=0 w=5.58 l=1.84
X21 VDD2.t0 VN.t9 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0.9207 ps=5.91 w=5.58 l=1.84
X22 VDD1.t0 VP.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=5.91 as=0.9207 ps=5.91 w=5.58 l=1.84
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1762 pd=11.94 as=0 ps=0 w=5.58 l=1.84
R0 VN.n31 VN.n30 181.465
R1 VN.n63 VN.n62 181.465
R2 VN.n61 VN.n32 161.3
R3 VN.n60 VN.n59 161.3
R4 VN.n58 VN.n33 161.3
R5 VN.n57 VN.n56 161.3
R6 VN.n55 VN.n34 161.3
R7 VN.n53 VN.n52 161.3
R8 VN.n51 VN.n35 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n36 161.3
R11 VN.n46 VN.n45 161.3
R12 VN.n44 VN.n37 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n41 VN.n38 161.3
R15 VN.n29 VN.n0 161.3
R16 VN.n28 VN.n27 161.3
R17 VN.n26 VN.n1 161.3
R18 VN.n25 VN.n24 161.3
R19 VN.n23 VN.n2 161.3
R20 VN.n21 VN.n20 161.3
R21 VN.n19 VN.n3 161.3
R22 VN.n18 VN.n17 161.3
R23 VN.n16 VN.n4 161.3
R24 VN.n14 VN.n13 161.3
R25 VN.n12 VN.n5 161.3
R26 VN.n11 VN.n10 161.3
R27 VN.n9 VN.n6 161.3
R28 VN.n7 VN.t1 107.987
R29 VN.n39 VN.t7 107.987
R30 VN.n8 VN.t6 73.0864
R31 VN.n15 VN.t3 73.0864
R32 VN.n22 VN.t0 73.0864
R33 VN.n30 VN.t8 73.0864
R34 VN.n40 VN.t4 73.0864
R35 VN.n47 VN.t5 73.0864
R36 VN.n54 VN.t2 73.0864
R37 VN.n62 VN.t9 73.0864
R38 VN.n10 VN.n5 56.5617
R39 VN.n17 VN.n3 56.5617
R40 VN.n42 VN.n37 56.5617
R41 VN.n49 VN.n35 56.5617
R42 VN.n8 VN.n7 48.9423
R43 VN.n40 VN.n39 48.9423
R44 VN VN.n63 44.4228
R45 VN.n28 VN.n1 41.0614
R46 VN.n60 VN.n33 41.0614
R47 VN.n24 VN.n1 40.0926
R48 VN.n56 VN.n33 40.0926
R49 VN.n10 VN.n9 24.5923
R50 VN.n14 VN.n5 24.5923
R51 VN.n17 VN.n16 24.5923
R52 VN.n21 VN.n3 24.5923
R53 VN.n24 VN.n23 24.5923
R54 VN.n29 VN.n28 24.5923
R55 VN.n42 VN.n41 24.5923
R56 VN.n49 VN.n48 24.5923
R57 VN.n46 VN.n37 24.5923
R58 VN.n56 VN.n55 24.5923
R59 VN.n53 VN.n35 24.5923
R60 VN.n61 VN.n60 24.5923
R61 VN.n9 VN.n8 20.6576
R62 VN.n22 VN.n21 20.6576
R63 VN.n41 VN.n40 20.6576
R64 VN.n54 VN.n53 20.6576
R65 VN.n15 VN.n14 12.2964
R66 VN.n16 VN.n15 12.2964
R67 VN.n48 VN.n47 12.2964
R68 VN.n47 VN.n46 12.2964
R69 VN.n39 VN.n38 12.2243
R70 VN.n7 VN.n6 12.2243
R71 VN.n30 VN.n29 4.42703
R72 VN.n62 VN.n61 4.42703
R73 VN.n23 VN.n22 3.93519
R74 VN.n55 VN.n54 3.93519
R75 VN.n63 VN.n32 0.189894
R76 VN.n59 VN.n32 0.189894
R77 VN.n59 VN.n58 0.189894
R78 VN.n58 VN.n57 0.189894
R79 VN.n57 VN.n34 0.189894
R80 VN.n52 VN.n34 0.189894
R81 VN.n52 VN.n51 0.189894
R82 VN.n51 VN.n50 0.189894
R83 VN.n50 VN.n36 0.189894
R84 VN.n45 VN.n36 0.189894
R85 VN.n45 VN.n44 0.189894
R86 VN.n44 VN.n43 0.189894
R87 VN.n43 VN.n38 0.189894
R88 VN.n11 VN.n6 0.189894
R89 VN.n12 VN.n11 0.189894
R90 VN.n13 VN.n12 0.189894
R91 VN.n13 VN.n4 0.189894
R92 VN.n18 VN.n4 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n20 VN.n19 0.189894
R95 VN.n20 VN.n2 0.189894
R96 VN.n25 VN.n2 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n27 VN.n26 0.189894
R99 VN.n27 VN.n0 0.189894
R100 VN.n31 VN.n0 0.189894
R101 VN VN.n31 0.0516364
R102 VDD2.n1 VDD2.t2 72.1252
R103 VDD2.n4 VDD2.t0 70.2548
R104 VDD2.n3 VDD2.n2 68.0538
R105 VDD2 VDD2.n7 68.0511
R106 VDD2.n6 VDD2.n5 66.7064
R107 VDD2.n1 VDD2.n0 66.7062
R108 VDD2.n4 VDD2.n3 37.4114
R109 VDD2.n7 VDD2.t1 3.54889
R110 VDD2.n7 VDD2.t3 3.54889
R111 VDD2.n5 VDD2.t9 3.54889
R112 VDD2.n5 VDD2.t5 3.54889
R113 VDD2.n2 VDD2.t4 3.54889
R114 VDD2.n2 VDD2.t7 3.54889
R115 VDD2.n0 VDD2.t6 3.54889
R116 VDD2.n0 VDD2.t8 3.54889
R117 VDD2.n6 VDD2.n4 1.87119
R118 VDD2 VDD2.n6 0.526362
R119 VDD2.n3 VDD2.n1 0.412826
R120 VTAIL.n11 VTAIL.t12 53.576
R121 VTAIL.n17 VTAIL.t11 53.5758
R122 VTAIL.n2 VTAIL.t0 53.5758
R123 VTAIL.n16 VTAIL.t8 53.5758
R124 VTAIL.n15 VTAIL.n14 50.0276
R125 VTAIL.n13 VTAIL.n12 50.0276
R126 VTAIL.n10 VTAIL.n9 50.0276
R127 VTAIL.n8 VTAIL.n7 50.0276
R128 VTAIL.n19 VTAIL.n18 50.0274
R129 VTAIL.n1 VTAIL.n0 50.0274
R130 VTAIL.n4 VTAIL.n3 50.0274
R131 VTAIL.n6 VTAIL.n5 50.0274
R132 VTAIL.n8 VTAIL.n6 20.9186
R133 VTAIL.n17 VTAIL.n16 19.0479
R134 VTAIL.n18 VTAIL.t16 3.54889
R135 VTAIL.n18 VTAIL.t19 3.54889
R136 VTAIL.n0 VTAIL.t18 3.54889
R137 VTAIL.n0 VTAIL.t13 3.54889
R138 VTAIL.n3 VTAIL.t6 3.54889
R139 VTAIL.n3 VTAIL.t3 3.54889
R140 VTAIL.n5 VTAIL.t5 3.54889
R141 VTAIL.n5 VTAIL.t9 3.54889
R142 VTAIL.n14 VTAIL.t1 3.54889
R143 VTAIL.n14 VTAIL.t4 3.54889
R144 VTAIL.n12 VTAIL.t2 3.54889
R145 VTAIL.n12 VTAIL.t7 3.54889
R146 VTAIL.n9 VTAIL.t14 3.54889
R147 VTAIL.n9 VTAIL.t15 3.54889
R148 VTAIL.n7 VTAIL.t10 3.54889
R149 VTAIL.n7 VTAIL.t17 3.54889
R150 VTAIL.n10 VTAIL.n8 1.87119
R151 VTAIL.n11 VTAIL.n10 1.87119
R152 VTAIL.n15 VTAIL.n13 1.87119
R153 VTAIL.n16 VTAIL.n15 1.87119
R154 VTAIL.n6 VTAIL.n4 1.87119
R155 VTAIL.n4 VTAIL.n2 1.87119
R156 VTAIL.n19 VTAIL.n17 1.87119
R157 VTAIL VTAIL.n1 1.46171
R158 VTAIL.n13 VTAIL.n11 1.40567
R159 VTAIL.n2 VTAIL.n1 1.40567
R160 VTAIL VTAIL.n19 0.409983
R161 B.n551 B.n550 585
R162 B.n551 B.n86 585
R163 B.n554 B.n553 585
R164 B.n555 B.n118 585
R165 B.n557 B.n556 585
R166 B.n559 B.n117 585
R167 B.n562 B.n561 585
R168 B.n563 B.n116 585
R169 B.n565 B.n564 585
R170 B.n567 B.n115 585
R171 B.n570 B.n569 585
R172 B.n571 B.n114 585
R173 B.n573 B.n572 585
R174 B.n575 B.n113 585
R175 B.n578 B.n577 585
R176 B.n579 B.n112 585
R177 B.n581 B.n580 585
R178 B.n583 B.n111 585
R179 B.n586 B.n585 585
R180 B.n587 B.n110 585
R181 B.n589 B.n588 585
R182 B.n591 B.n109 585
R183 B.n594 B.n593 585
R184 B.n595 B.n106 585
R185 B.n598 B.n597 585
R186 B.n600 B.n105 585
R187 B.n603 B.n602 585
R188 B.n604 B.n104 585
R189 B.n606 B.n605 585
R190 B.n608 B.n103 585
R191 B.n611 B.n610 585
R192 B.n612 B.n99 585
R193 B.n614 B.n613 585
R194 B.n616 B.n98 585
R195 B.n619 B.n618 585
R196 B.n620 B.n97 585
R197 B.n622 B.n621 585
R198 B.n624 B.n96 585
R199 B.n627 B.n626 585
R200 B.n628 B.n95 585
R201 B.n630 B.n629 585
R202 B.n632 B.n94 585
R203 B.n635 B.n634 585
R204 B.n636 B.n93 585
R205 B.n638 B.n637 585
R206 B.n640 B.n92 585
R207 B.n643 B.n642 585
R208 B.n644 B.n91 585
R209 B.n646 B.n645 585
R210 B.n648 B.n90 585
R211 B.n651 B.n650 585
R212 B.n652 B.n89 585
R213 B.n654 B.n653 585
R214 B.n656 B.n88 585
R215 B.n659 B.n658 585
R216 B.n660 B.n87 585
R217 B.n549 B.n85 585
R218 B.n663 B.n85 585
R219 B.n548 B.n84 585
R220 B.n664 B.n84 585
R221 B.n547 B.n83 585
R222 B.n665 B.n83 585
R223 B.n546 B.n545 585
R224 B.n545 B.n79 585
R225 B.n544 B.n78 585
R226 B.n671 B.n78 585
R227 B.n543 B.n77 585
R228 B.n672 B.n77 585
R229 B.n542 B.n76 585
R230 B.n673 B.n76 585
R231 B.n541 B.n540 585
R232 B.n540 B.n72 585
R233 B.n539 B.n71 585
R234 B.n679 B.n71 585
R235 B.n538 B.n70 585
R236 B.n680 B.n70 585
R237 B.n537 B.n69 585
R238 B.n681 B.n69 585
R239 B.n536 B.n535 585
R240 B.n535 B.n65 585
R241 B.n534 B.n64 585
R242 B.n687 B.n64 585
R243 B.n533 B.n63 585
R244 B.n688 B.n63 585
R245 B.n532 B.n62 585
R246 B.n689 B.n62 585
R247 B.n531 B.n530 585
R248 B.n530 B.n58 585
R249 B.n529 B.n57 585
R250 B.n695 B.n57 585
R251 B.n528 B.n56 585
R252 B.n696 B.n56 585
R253 B.n527 B.n55 585
R254 B.n697 B.n55 585
R255 B.n526 B.n525 585
R256 B.n525 B.n51 585
R257 B.n524 B.n50 585
R258 B.n703 B.n50 585
R259 B.n523 B.n49 585
R260 B.n704 B.n49 585
R261 B.n522 B.n48 585
R262 B.n705 B.n48 585
R263 B.n521 B.n520 585
R264 B.n520 B.n44 585
R265 B.n519 B.n43 585
R266 B.n711 B.n43 585
R267 B.n518 B.n42 585
R268 B.n712 B.n42 585
R269 B.n517 B.n41 585
R270 B.n713 B.n41 585
R271 B.n516 B.n515 585
R272 B.n515 B.n37 585
R273 B.n514 B.n36 585
R274 B.n719 B.n36 585
R275 B.n513 B.n35 585
R276 B.n720 B.n35 585
R277 B.n512 B.n34 585
R278 B.n721 B.n34 585
R279 B.n511 B.n510 585
R280 B.n510 B.n30 585
R281 B.n509 B.n29 585
R282 B.n727 B.n29 585
R283 B.n508 B.n28 585
R284 B.n728 B.n28 585
R285 B.n507 B.n27 585
R286 B.n729 B.n27 585
R287 B.n506 B.n505 585
R288 B.n505 B.n26 585
R289 B.n504 B.n22 585
R290 B.n735 B.n22 585
R291 B.n503 B.n21 585
R292 B.n736 B.n21 585
R293 B.n502 B.n20 585
R294 B.n737 B.n20 585
R295 B.n501 B.n500 585
R296 B.n500 B.n16 585
R297 B.n499 B.n15 585
R298 B.n743 B.n15 585
R299 B.n498 B.n14 585
R300 B.n744 B.n14 585
R301 B.n497 B.n13 585
R302 B.n745 B.n13 585
R303 B.n496 B.n495 585
R304 B.n495 B.n12 585
R305 B.n494 B.n493 585
R306 B.n494 B.n8 585
R307 B.n492 B.n7 585
R308 B.n752 B.n7 585
R309 B.n491 B.n6 585
R310 B.n753 B.n6 585
R311 B.n490 B.n5 585
R312 B.n754 B.n5 585
R313 B.n489 B.n488 585
R314 B.n488 B.n4 585
R315 B.n487 B.n119 585
R316 B.n487 B.n486 585
R317 B.n477 B.n120 585
R318 B.n121 B.n120 585
R319 B.n479 B.n478 585
R320 B.n480 B.n479 585
R321 B.n476 B.n125 585
R322 B.n129 B.n125 585
R323 B.n475 B.n474 585
R324 B.n474 B.n473 585
R325 B.n127 B.n126 585
R326 B.n128 B.n127 585
R327 B.n466 B.n465 585
R328 B.n467 B.n466 585
R329 B.n464 B.n134 585
R330 B.n134 B.n133 585
R331 B.n463 B.n462 585
R332 B.n462 B.n461 585
R333 B.n136 B.n135 585
R334 B.n454 B.n136 585
R335 B.n453 B.n452 585
R336 B.n455 B.n453 585
R337 B.n451 B.n141 585
R338 B.n141 B.n140 585
R339 B.n450 B.n449 585
R340 B.n449 B.n448 585
R341 B.n143 B.n142 585
R342 B.n144 B.n143 585
R343 B.n441 B.n440 585
R344 B.n442 B.n441 585
R345 B.n439 B.n149 585
R346 B.n149 B.n148 585
R347 B.n438 B.n437 585
R348 B.n437 B.n436 585
R349 B.n151 B.n150 585
R350 B.n152 B.n151 585
R351 B.n429 B.n428 585
R352 B.n430 B.n429 585
R353 B.n427 B.n157 585
R354 B.n157 B.n156 585
R355 B.n426 B.n425 585
R356 B.n425 B.n424 585
R357 B.n159 B.n158 585
R358 B.n160 B.n159 585
R359 B.n417 B.n416 585
R360 B.n418 B.n417 585
R361 B.n415 B.n165 585
R362 B.n165 B.n164 585
R363 B.n414 B.n413 585
R364 B.n413 B.n412 585
R365 B.n167 B.n166 585
R366 B.n168 B.n167 585
R367 B.n405 B.n404 585
R368 B.n406 B.n405 585
R369 B.n403 B.n173 585
R370 B.n173 B.n172 585
R371 B.n402 B.n401 585
R372 B.n401 B.n400 585
R373 B.n175 B.n174 585
R374 B.n176 B.n175 585
R375 B.n393 B.n392 585
R376 B.n394 B.n393 585
R377 B.n391 B.n181 585
R378 B.n181 B.n180 585
R379 B.n390 B.n389 585
R380 B.n389 B.n388 585
R381 B.n183 B.n182 585
R382 B.n184 B.n183 585
R383 B.n381 B.n380 585
R384 B.n382 B.n381 585
R385 B.n379 B.n189 585
R386 B.n189 B.n188 585
R387 B.n378 B.n377 585
R388 B.n377 B.n376 585
R389 B.n191 B.n190 585
R390 B.n192 B.n191 585
R391 B.n369 B.n368 585
R392 B.n370 B.n369 585
R393 B.n367 B.n197 585
R394 B.n197 B.n196 585
R395 B.n366 B.n365 585
R396 B.n365 B.n364 585
R397 B.n199 B.n198 585
R398 B.n200 B.n199 585
R399 B.n357 B.n356 585
R400 B.n358 B.n357 585
R401 B.n355 B.n205 585
R402 B.n205 B.n204 585
R403 B.n354 B.n353 585
R404 B.n353 B.n352 585
R405 B.n349 B.n209 585
R406 B.n348 B.n347 585
R407 B.n345 B.n210 585
R408 B.n345 B.n208 585
R409 B.n344 B.n343 585
R410 B.n342 B.n341 585
R411 B.n340 B.n212 585
R412 B.n338 B.n337 585
R413 B.n336 B.n213 585
R414 B.n335 B.n334 585
R415 B.n332 B.n214 585
R416 B.n330 B.n329 585
R417 B.n328 B.n215 585
R418 B.n327 B.n326 585
R419 B.n324 B.n216 585
R420 B.n322 B.n321 585
R421 B.n320 B.n217 585
R422 B.n319 B.n318 585
R423 B.n316 B.n218 585
R424 B.n314 B.n313 585
R425 B.n312 B.n219 585
R426 B.n311 B.n310 585
R427 B.n308 B.n220 585
R428 B.n306 B.n305 585
R429 B.n303 B.n221 585
R430 B.n302 B.n301 585
R431 B.n299 B.n224 585
R432 B.n297 B.n296 585
R433 B.n295 B.n225 585
R434 B.n294 B.n293 585
R435 B.n291 B.n226 585
R436 B.n289 B.n288 585
R437 B.n287 B.n227 585
R438 B.n285 B.n284 585
R439 B.n282 B.n230 585
R440 B.n280 B.n279 585
R441 B.n278 B.n231 585
R442 B.n277 B.n276 585
R443 B.n274 B.n232 585
R444 B.n272 B.n271 585
R445 B.n270 B.n233 585
R446 B.n269 B.n268 585
R447 B.n266 B.n234 585
R448 B.n264 B.n263 585
R449 B.n262 B.n235 585
R450 B.n261 B.n260 585
R451 B.n258 B.n236 585
R452 B.n256 B.n255 585
R453 B.n254 B.n237 585
R454 B.n253 B.n252 585
R455 B.n250 B.n238 585
R456 B.n248 B.n247 585
R457 B.n246 B.n239 585
R458 B.n245 B.n244 585
R459 B.n242 B.n240 585
R460 B.n207 B.n206 585
R461 B.n351 B.n350 585
R462 B.n352 B.n351 585
R463 B.n203 B.n202 585
R464 B.n204 B.n203 585
R465 B.n360 B.n359 585
R466 B.n359 B.n358 585
R467 B.n361 B.n201 585
R468 B.n201 B.n200 585
R469 B.n363 B.n362 585
R470 B.n364 B.n363 585
R471 B.n195 B.n194 585
R472 B.n196 B.n195 585
R473 B.n372 B.n371 585
R474 B.n371 B.n370 585
R475 B.n373 B.n193 585
R476 B.n193 B.n192 585
R477 B.n375 B.n374 585
R478 B.n376 B.n375 585
R479 B.n187 B.n186 585
R480 B.n188 B.n187 585
R481 B.n384 B.n383 585
R482 B.n383 B.n382 585
R483 B.n385 B.n185 585
R484 B.n185 B.n184 585
R485 B.n387 B.n386 585
R486 B.n388 B.n387 585
R487 B.n179 B.n178 585
R488 B.n180 B.n179 585
R489 B.n396 B.n395 585
R490 B.n395 B.n394 585
R491 B.n397 B.n177 585
R492 B.n177 B.n176 585
R493 B.n399 B.n398 585
R494 B.n400 B.n399 585
R495 B.n171 B.n170 585
R496 B.n172 B.n171 585
R497 B.n408 B.n407 585
R498 B.n407 B.n406 585
R499 B.n409 B.n169 585
R500 B.n169 B.n168 585
R501 B.n411 B.n410 585
R502 B.n412 B.n411 585
R503 B.n163 B.n162 585
R504 B.n164 B.n163 585
R505 B.n420 B.n419 585
R506 B.n419 B.n418 585
R507 B.n421 B.n161 585
R508 B.n161 B.n160 585
R509 B.n423 B.n422 585
R510 B.n424 B.n423 585
R511 B.n155 B.n154 585
R512 B.n156 B.n155 585
R513 B.n432 B.n431 585
R514 B.n431 B.n430 585
R515 B.n433 B.n153 585
R516 B.n153 B.n152 585
R517 B.n435 B.n434 585
R518 B.n436 B.n435 585
R519 B.n147 B.n146 585
R520 B.n148 B.n147 585
R521 B.n444 B.n443 585
R522 B.n443 B.n442 585
R523 B.n445 B.n145 585
R524 B.n145 B.n144 585
R525 B.n447 B.n446 585
R526 B.n448 B.n447 585
R527 B.n139 B.n138 585
R528 B.n140 B.n139 585
R529 B.n457 B.n456 585
R530 B.n456 B.n455 585
R531 B.n458 B.n137 585
R532 B.n454 B.n137 585
R533 B.n460 B.n459 585
R534 B.n461 B.n460 585
R535 B.n132 B.n131 585
R536 B.n133 B.n132 585
R537 B.n469 B.n468 585
R538 B.n468 B.n467 585
R539 B.n470 B.n130 585
R540 B.n130 B.n128 585
R541 B.n472 B.n471 585
R542 B.n473 B.n472 585
R543 B.n124 B.n123 585
R544 B.n129 B.n124 585
R545 B.n482 B.n481 585
R546 B.n481 B.n480 585
R547 B.n483 B.n122 585
R548 B.n122 B.n121 585
R549 B.n485 B.n484 585
R550 B.n486 B.n485 585
R551 B.n3 B.n0 585
R552 B.n4 B.n3 585
R553 B.n751 B.n1 585
R554 B.n752 B.n751 585
R555 B.n750 B.n749 585
R556 B.n750 B.n8 585
R557 B.n748 B.n9 585
R558 B.n12 B.n9 585
R559 B.n747 B.n746 585
R560 B.n746 B.n745 585
R561 B.n11 B.n10 585
R562 B.n744 B.n11 585
R563 B.n742 B.n741 585
R564 B.n743 B.n742 585
R565 B.n740 B.n17 585
R566 B.n17 B.n16 585
R567 B.n739 B.n738 585
R568 B.n738 B.n737 585
R569 B.n19 B.n18 585
R570 B.n736 B.n19 585
R571 B.n734 B.n733 585
R572 B.n735 B.n734 585
R573 B.n732 B.n23 585
R574 B.n26 B.n23 585
R575 B.n731 B.n730 585
R576 B.n730 B.n729 585
R577 B.n25 B.n24 585
R578 B.n728 B.n25 585
R579 B.n726 B.n725 585
R580 B.n727 B.n726 585
R581 B.n724 B.n31 585
R582 B.n31 B.n30 585
R583 B.n723 B.n722 585
R584 B.n722 B.n721 585
R585 B.n33 B.n32 585
R586 B.n720 B.n33 585
R587 B.n718 B.n717 585
R588 B.n719 B.n718 585
R589 B.n716 B.n38 585
R590 B.n38 B.n37 585
R591 B.n715 B.n714 585
R592 B.n714 B.n713 585
R593 B.n40 B.n39 585
R594 B.n712 B.n40 585
R595 B.n710 B.n709 585
R596 B.n711 B.n710 585
R597 B.n708 B.n45 585
R598 B.n45 B.n44 585
R599 B.n707 B.n706 585
R600 B.n706 B.n705 585
R601 B.n47 B.n46 585
R602 B.n704 B.n47 585
R603 B.n702 B.n701 585
R604 B.n703 B.n702 585
R605 B.n700 B.n52 585
R606 B.n52 B.n51 585
R607 B.n699 B.n698 585
R608 B.n698 B.n697 585
R609 B.n54 B.n53 585
R610 B.n696 B.n54 585
R611 B.n694 B.n693 585
R612 B.n695 B.n694 585
R613 B.n692 B.n59 585
R614 B.n59 B.n58 585
R615 B.n691 B.n690 585
R616 B.n690 B.n689 585
R617 B.n61 B.n60 585
R618 B.n688 B.n61 585
R619 B.n686 B.n685 585
R620 B.n687 B.n686 585
R621 B.n684 B.n66 585
R622 B.n66 B.n65 585
R623 B.n683 B.n682 585
R624 B.n682 B.n681 585
R625 B.n68 B.n67 585
R626 B.n680 B.n68 585
R627 B.n678 B.n677 585
R628 B.n679 B.n678 585
R629 B.n676 B.n73 585
R630 B.n73 B.n72 585
R631 B.n675 B.n674 585
R632 B.n674 B.n673 585
R633 B.n75 B.n74 585
R634 B.n672 B.n75 585
R635 B.n670 B.n669 585
R636 B.n671 B.n670 585
R637 B.n668 B.n80 585
R638 B.n80 B.n79 585
R639 B.n667 B.n666 585
R640 B.n666 B.n665 585
R641 B.n82 B.n81 585
R642 B.n664 B.n82 585
R643 B.n662 B.n661 585
R644 B.n663 B.n662 585
R645 B.n755 B.n754 585
R646 B.n753 B.n2 585
R647 B.n662 B.n87 487.695
R648 B.n551 B.n85 487.695
R649 B.n353 B.n207 487.695
R650 B.n351 B.n209 487.695
R651 B.n100 B.t14 279.601
R652 B.n107 B.t18 279.601
R653 B.n228 B.t10 279.601
R654 B.n222 B.t21 279.601
R655 B.n552 B.n86 256.663
R656 B.n558 B.n86 256.663
R657 B.n560 B.n86 256.663
R658 B.n566 B.n86 256.663
R659 B.n568 B.n86 256.663
R660 B.n574 B.n86 256.663
R661 B.n576 B.n86 256.663
R662 B.n582 B.n86 256.663
R663 B.n584 B.n86 256.663
R664 B.n590 B.n86 256.663
R665 B.n592 B.n86 256.663
R666 B.n599 B.n86 256.663
R667 B.n601 B.n86 256.663
R668 B.n607 B.n86 256.663
R669 B.n609 B.n86 256.663
R670 B.n615 B.n86 256.663
R671 B.n617 B.n86 256.663
R672 B.n623 B.n86 256.663
R673 B.n625 B.n86 256.663
R674 B.n631 B.n86 256.663
R675 B.n633 B.n86 256.663
R676 B.n639 B.n86 256.663
R677 B.n641 B.n86 256.663
R678 B.n647 B.n86 256.663
R679 B.n649 B.n86 256.663
R680 B.n655 B.n86 256.663
R681 B.n657 B.n86 256.663
R682 B.n346 B.n208 256.663
R683 B.n211 B.n208 256.663
R684 B.n339 B.n208 256.663
R685 B.n333 B.n208 256.663
R686 B.n331 B.n208 256.663
R687 B.n325 B.n208 256.663
R688 B.n323 B.n208 256.663
R689 B.n317 B.n208 256.663
R690 B.n315 B.n208 256.663
R691 B.n309 B.n208 256.663
R692 B.n307 B.n208 256.663
R693 B.n300 B.n208 256.663
R694 B.n298 B.n208 256.663
R695 B.n292 B.n208 256.663
R696 B.n290 B.n208 256.663
R697 B.n283 B.n208 256.663
R698 B.n281 B.n208 256.663
R699 B.n275 B.n208 256.663
R700 B.n273 B.n208 256.663
R701 B.n267 B.n208 256.663
R702 B.n265 B.n208 256.663
R703 B.n259 B.n208 256.663
R704 B.n257 B.n208 256.663
R705 B.n251 B.n208 256.663
R706 B.n249 B.n208 256.663
R707 B.n243 B.n208 256.663
R708 B.n241 B.n208 256.663
R709 B.n757 B.n756 256.663
R710 B.n658 B.n656 163.367
R711 B.n654 B.n89 163.367
R712 B.n650 B.n648 163.367
R713 B.n646 B.n91 163.367
R714 B.n642 B.n640 163.367
R715 B.n638 B.n93 163.367
R716 B.n634 B.n632 163.367
R717 B.n630 B.n95 163.367
R718 B.n626 B.n624 163.367
R719 B.n622 B.n97 163.367
R720 B.n618 B.n616 163.367
R721 B.n614 B.n99 163.367
R722 B.n610 B.n608 163.367
R723 B.n606 B.n104 163.367
R724 B.n602 B.n600 163.367
R725 B.n598 B.n106 163.367
R726 B.n593 B.n591 163.367
R727 B.n589 B.n110 163.367
R728 B.n585 B.n583 163.367
R729 B.n581 B.n112 163.367
R730 B.n577 B.n575 163.367
R731 B.n573 B.n114 163.367
R732 B.n569 B.n567 163.367
R733 B.n565 B.n116 163.367
R734 B.n561 B.n559 163.367
R735 B.n557 B.n118 163.367
R736 B.n553 B.n551 163.367
R737 B.n353 B.n205 163.367
R738 B.n357 B.n205 163.367
R739 B.n357 B.n199 163.367
R740 B.n365 B.n199 163.367
R741 B.n365 B.n197 163.367
R742 B.n369 B.n197 163.367
R743 B.n369 B.n191 163.367
R744 B.n377 B.n191 163.367
R745 B.n377 B.n189 163.367
R746 B.n381 B.n189 163.367
R747 B.n381 B.n183 163.367
R748 B.n389 B.n183 163.367
R749 B.n389 B.n181 163.367
R750 B.n393 B.n181 163.367
R751 B.n393 B.n175 163.367
R752 B.n401 B.n175 163.367
R753 B.n401 B.n173 163.367
R754 B.n405 B.n173 163.367
R755 B.n405 B.n167 163.367
R756 B.n413 B.n167 163.367
R757 B.n413 B.n165 163.367
R758 B.n417 B.n165 163.367
R759 B.n417 B.n159 163.367
R760 B.n425 B.n159 163.367
R761 B.n425 B.n157 163.367
R762 B.n429 B.n157 163.367
R763 B.n429 B.n151 163.367
R764 B.n437 B.n151 163.367
R765 B.n437 B.n149 163.367
R766 B.n441 B.n149 163.367
R767 B.n441 B.n143 163.367
R768 B.n449 B.n143 163.367
R769 B.n449 B.n141 163.367
R770 B.n453 B.n141 163.367
R771 B.n453 B.n136 163.367
R772 B.n462 B.n136 163.367
R773 B.n462 B.n134 163.367
R774 B.n466 B.n134 163.367
R775 B.n466 B.n127 163.367
R776 B.n474 B.n127 163.367
R777 B.n474 B.n125 163.367
R778 B.n479 B.n125 163.367
R779 B.n479 B.n120 163.367
R780 B.n487 B.n120 163.367
R781 B.n488 B.n487 163.367
R782 B.n488 B.n5 163.367
R783 B.n6 B.n5 163.367
R784 B.n7 B.n6 163.367
R785 B.n494 B.n7 163.367
R786 B.n495 B.n494 163.367
R787 B.n495 B.n13 163.367
R788 B.n14 B.n13 163.367
R789 B.n15 B.n14 163.367
R790 B.n500 B.n15 163.367
R791 B.n500 B.n20 163.367
R792 B.n21 B.n20 163.367
R793 B.n22 B.n21 163.367
R794 B.n505 B.n22 163.367
R795 B.n505 B.n27 163.367
R796 B.n28 B.n27 163.367
R797 B.n29 B.n28 163.367
R798 B.n510 B.n29 163.367
R799 B.n510 B.n34 163.367
R800 B.n35 B.n34 163.367
R801 B.n36 B.n35 163.367
R802 B.n515 B.n36 163.367
R803 B.n515 B.n41 163.367
R804 B.n42 B.n41 163.367
R805 B.n43 B.n42 163.367
R806 B.n520 B.n43 163.367
R807 B.n520 B.n48 163.367
R808 B.n49 B.n48 163.367
R809 B.n50 B.n49 163.367
R810 B.n525 B.n50 163.367
R811 B.n525 B.n55 163.367
R812 B.n56 B.n55 163.367
R813 B.n57 B.n56 163.367
R814 B.n530 B.n57 163.367
R815 B.n530 B.n62 163.367
R816 B.n63 B.n62 163.367
R817 B.n64 B.n63 163.367
R818 B.n535 B.n64 163.367
R819 B.n535 B.n69 163.367
R820 B.n70 B.n69 163.367
R821 B.n71 B.n70 163.367
R822 B.n540 B.n71 163.367
R823 B.n540 B.n76 163.367
R824 B.n77 B.n76 163.367
R825 B.n78 B.n77 163.367
R826 B.n545 B.n78 163.367
R827 B.n545 B.n83 163.367
R828 B.n84 B.n83 163.367
R829 B.n85 B.n84 163.367
R830 B.n347 B.n345 163.367
R831 B.n345 B.n344 163.367
R832 B.n341 B.n340 163.367
R833 B.n338 B.n213 163.367
R834 B.n334 B.n332 163.367
R835 B.n330 B.n215 163.367
R836 B.n326 B.n324 163.367
R837 B.n322 B.n217 163.367
R838 B.n318 B.n316 163.367
R839 B.n314 B.n219 163.367
R840 B.n310 B.n308 163.367
R841 B.n306 B.n221 163.367
R842 B.n301 B.n299 163.367
R843 B.n297 B.n225 163.367
R844 B.n293 B.n291 163.367
R845 B.n289 B.n227 163.367
R846 B.n284 B.n282 163.367
R847 B.n280 B.n231 163.367
R848 B.n276 B.n274 163.367
R849 B.n272 B.n233 163.367
R850 B.n268 B.n266 163.367
R851 B.n264 B.n235 163.367
R852 B.n260 B.n258 163.367
R853 B.n256 B.n237 163.367
R854 B.n252 B.n250 163.367
R855 B.n248 B.n239 163.367
R856 B.n244 B.n242 163.367
R857 B.n351 B.n203 163.367
R858 B.n359 B.n203 163.367
R859 B.n359 B.n201 163.367
R860 B.n363 B.n201 163.367
R861 B.n363 B.n195 163.367
R862 B.n371 B.n195 163.367
R863 B.n371 B.n193 163.367
R864 B.n375 B.n193 163.367
R865 B.n375 B.n187 163.367
R866 B.n383 B.n187 163.367
R867 B.n383 B.n185 163.367
R868 B.n387 B.n185 163.367
R869 B.n387 B.n179 163.367
R870 B.n395 B.n179 163.367
R871 B.n395 B.n177 163.367
R872 B.n399 B.n177 163.367
R873 B.n399 B.n171 163.367
R874 B.n407 B.n171 163.367
R875 B.n407 B.n169 163.367
R876 B.n411 B.n169 163.367
R877 B.n411 B.n163 163.367
R878 B.n419 B.n163 163.367
R879 B.n419 B.n161 163.367
R880 B.n423 B.n161 163.367
R881 B.n423 B.n155 163.367
R882 B.n431 B.n155 163.367
R883 B.n431 B.n153 163.367
R884 B.n435 B.n153 163.367
R885 B.n435 B.n147 163.367
R886 B.n443 B.n147 163.367
R887 B.n443 B.n145 163.367
R888 B.n447 B.n145 163.367
R889 B.n447 B.n139 163.367
R890 B.n456 B.n139 163.367
R891 B.n456 B.n137 163.367
R892 B.n460 B.n137 163.367
R893 B.n460 B.n132 163.367
R894 B.n468 B.n132 163.367
R895 B.n468 B.n130 163.367
R896 B.n472 B.n130 163.367
R897 B.n472 B.n124 163.367
R898 B.n481 B.n124 163.367
R899 B.n481 B.n122 163.367
R900 B.n485 B.n122 163.367
R901 B.n485 B.n3 163.367
R902 B.n755 B.n3 163.367
R903 B.n751 B.n2 163.367
R904 B.n751 B.n750 163.367
R905 B.n750 B.n9 163.367
R906 B.n746 B.n9 163.367
R907 B.n746 B.n11 163.367
R908 B.n742 B.n11 163.367
R909 B.n742 B.n17 163.367
R910 B.n738 B.n17 163.367
R911 B.n738 B.n19 163.367
R912 B.n734 B.n19 163.367
R913 B.n734 B.n23 163.367
R914 B.n730 B.n23 163.367
R915 B.n730 B.n25 163.367
R916 B.n726 B.n25 163.367
R917 B.n726 B.n31 163.367
R918 B.n722 B.n31 163.367
R919 B.n722 B.n33 163.367
R920 B.n718 B.n33 163.367
R921 B.n718 B.n38 163.367
R922 B.n714 B.n38 163.367
R923 B.n714 B.n40 163.367
R924 B.n710 B.n40 163.367
R925 B.n710 B.n45 163.367
R926 B.n706 B.n45 163.367
R927 B.n706 B.n47 163.367
R928 B.n702 B.n47 163.367
R929 B.n702 B.n52 163.367
R930 B.n698 B.n52 163.367
R931 B.n698 B.n54 163.367
R932 B.n694 B.n54 163.367
R933 B.n694 B.n59 163.367
R934 B.n690 B.n59 163.367
R935 B.n690 B.n61 163.367
R936 B.n686 B.n61 163.367
R937 B.n686 B.n66 163.367
R938 B.n682 B.n66 163.367
R939 B.n682 B.n68 163.367
R940 B.n678 B.n68 163.367
R941 B.n678 B.n73 163.367
R942 B.n674 B.n73 163.367
R943 B.n674 B.n75 163.367
R944 B.n670 B.n75 163.367
R945 B.n670 B.n80 163.367
R946 B.n666 B.n80 163.367
R947 B.n666 B.n82 163.367
R948 B.n662 B.n82 163.367
R949 B.n352 B.n208 118.564
R950 B.n663 B.n86 118.564
R951 B.n107 B.t19 114.513
R952 B.n228 B.t13 114.513
R953 B.n100 B.t16 114.507
R954 B.n222 B.t23 114.507
R955 B.n108 B.t20 72.4279
R956 B.n229 B.t12 72.4279
R957 B.n101 B.t17 72.4221
R958 B.n223 B.t22 72.4221
R959 B.n657 B.n87 71.676
R960 B.n656 B.n655 71.676
R961 B.n649 B.n89 71.676
R962 B.n648 B.n647 71.676
R963 B.n641 B.n91 71.676
R964 B.n640 B.n639 71.676
R965 B.n633 B.n93 71.676
R966 B.n632 B.n631 71.676
R967 B.n625 B.n95 71.676
R968 B.n624 B.n623 71.676
R969 B.n617 B.n97 71.676
R970 B.n616 B.n615 71.676
R971 B.n609 B.n99 71.676
R972 B.n608 B.n607 71.676
R973 B.n601 B.n104 71.676
R974 B.n600 B.n599 71.676
R975 B.n592 B.n106 71.676
R976 B.n591 B.n590 71.676
R977 B.n584 B.n110 71.676
R978 B.n583 B.n582 71.676
R979 B.n576 B.n112 71.676
R980 B.n575 B.n574 71.676
R981 B.n568 B.n114 71.676
R982 B.n567 B.n566 71.676
R983 B.n560 B.n116 71.676
R984 B.n559 B.n558 71.676
R985 B.n552 B.n118 71.676
R986 B.n553 B.n552 71.676
R987 B.n558 B.n557 71.676
R988 B.n561 B.n560 71.676
R989 B.n566 B.n565 71.676
R990 B.n569 B.n568 71.676
R991 B.n574 B.n573 71.676
R992 B.n577 B.n576 71.676
R993 B.n582 B.n581 71.676
R994 B.n585 B.n584 71.676
R995 B.n590 B.n589 71.676
R996 B.n593 B.n592 71.676
R997 B.n599 B.n598 71.676
R998 B.n602 B.n601 71.676
R999 B.n607 B.n606 71.676
R1000 B.n610 B.n609 71.676
R1001 B.n615 B.n614 71.676
R1002 B.n618 B.n617 71.676
R1003 B.n623 B.n622 71.676
R1004 B.n626 B.n625 71.676
R1005 B.n631 B.n630 71.676
R1006 B.n634 B.n633 71.676
R1007 B.n639 B.n638 71.676
R1008 B.n642 B.n641 71.676
R1009 B.n647 B.n646 71.676
R1010 B.n650 B.n649 71.676
R1011 B.n655 B.n654 71.676
R1012 B.n658 B.n657 71.676
R1013 B.n346 B.n209 71.676
R1014 B.n344 B.n211 71.676
R1015 B.n340 B.n339 71.676
R1016 B.n333 B.n213 71.676
R1017 B.n332 B.n331 71.676
R1018 B.n325 B.n215 71.676
R1019 B.n324 B.n323 71.676
R1020 B.n317 B.n217 71.676
R1021 B.n316 B.n315 71.676
R1022 B.n309 B.n219 71.676
R1023 B.n308 B.n307 71.676
R1024 B.n300 B.n221 71.676
R1025 B.n299 B.n298 71.676
R1026 B.n292 B.n225 71.676
R1027 B.n291 B.n290 71.676
R1028 B.n283 B.n227 71.676
R1029 B.n282 B.n281 71.676
R1030 B.n275 B.n231 71.676
R1031 B.n274 B.n273 71.676
R1032 B.n267 B.n233 71.676
R1033 B.n266 B.n265 71.676
R1034 B.n259 B.n235 71.676
R1035 B.n258 B.n257 71.676
R1036 B.n251 B.n237 71.676
R1037 B.n250 B.n249 71.676
R1038 B.n243 B.n239 71.676
R1039 B.n242 B.n241 71.676
R1040 B.n347 B.n346 71.676
R1041 B.n341 B.n211 71.676
R1042 B.n339 B.n338 71.676
R1043 B.n334 B.n333 71.676
R1044 B.n331 B.n330 71.676
R1045 B.n326 B.n325 71.676
R1046 B.n323 B.n322 71.676
R1047 B.n318 B.n317 71.676
R1048 B.n315 B.n314 71.676
R1049 B.n310 B.n309 71.676
R1050 B.n307 B.n306 71.676
R1051 B.n301 B.n300 71.676
R1052 B.n298 B.n297 71.676
R1053 B.n293 B.n292 71.676
R1054 B.n290 B.n289 71.676
R1055 B.n284 B.n283 71.676
R1056 B.n281 B.n280 71.676
R1057 B.n276 B.n275 71.676
R1058 B.n273 B.n272 71.676
R1059 B.n268 B.n267 71.676
R1060 B.n265 B.n264 71.676
R1061 B.n260 B.n259 71.676
R1062 B.n257 B.n256 71.676
R1063 B.n252 B.n251 71.676
R1064 B.n249 B.n248 71.676
R1065 B.n244 B.n243 71.676
R1066 B.n241 B.n207 71.676
R1067 B.n756 B.n755 71.676
R1068 B.n756 B.n2 71.676
R1069 B.n352 B.n204 68.9088
R1070 B.n358 B.n204 68.9088
R1071 B.n358 B.n200 68.9088
R1072 B.n364 B.n200 68.9088
R1073 B.n364 B.n196 68.9088
R1074 B.n370 B.n196 68.9088
R1075 B.n376 B.n192 68.9088
R1076 B.n376 B.n188 68.9088
R1077 B.n382 B.n188 68.9088
R1078 B.n382 B.n184 68.9088
R1079 B.n388 B.n184 68.9088
R1080 B.n388 B.n180 68.9088
R1081 B.n394 B.n180 68.9088
R1082 B.n394 B.n176 68.9088
R1083 B.n400 B.n176 68.9088
R1084 B.n406 B.n172 68.9088
R1085 B.n406 B.n168 68.9088
R1086 B.n412 B.n168 68.9088
R1087 B.n412 B.n164 68.9088
R1088 B.n418 B.n164 68.9088
R1089 B.n424 B.n160 68.9088
R1090 B.n424 B.n156 68.9088
R1091 B.n430 B.n156 68.9088
R1092 B.n430 B.n152 68.9088
R1093 B.n436 B.n152 68.9088
R1094 B.n442 B.n148 68.9088
R1095 B.n442 B.n144 68.9088
R1096 B.n448 B.n144 68.9088
R1097 B.n448 B.n140 68.9088
R1098 B.n455 B.n140 68.9088
R1099 B.n455 B.n454 68.9088
R1100 B.n461 B.n133 68.9088
R1101 B.n467 B.n133 68.9088
R1102 B.n467 B.n128 68.9088
R1103 B.n473 B.n128 68.9088
R1104 B.n473 B.n129 68.9088
R1105 B.n480 B.n121 68.9088
R1106 B.n486 B.n121 68.9088
R1107 B.n486 B.n4 68.9088
R1108 B.n754 B.n4 68.9088
R1109 B.n754 B.n753 68.9088
R1110 B.n753 B.n752 68.9088
R1111 B.n752 B.n8 68.9088
R1112 B.n12 B.n8 68.9088
R1113 B.n745 B.n12 68.9088
R1114 B.n744 B.n743 68.9088
R1115 B.n743 B.n16 68.9088
R1116 B.n737 B.n16 68.9088
R1117 B.n737 B.n736 68.9088
R1118 B.n736 B.n735 68.9088
R1119 B.n729 B.n26 68.9088
R1120 B.n729 B.n728 68.9088
R1121 B.n728 B.n727 68.9088
R1122 B.n727 B.n30 68.9088
R1123 B.n721 B.n30 68.9088
R1124 B.n721 B.n720 68.9088
R1125 B.n719 B.n37 68.9088
R1126 B.n713 B.n37 68.9088
R1127 B.n713 B.n712 68.9088
R1128 B.n712 B.n711 68.9088
R1129 B.n711 B.n44 68.9088
R1130 B.n705 B.n704 68.9088
R1131 B.n704 B.n703 68.9088
R1132 B.n703 B.n51 68.9088
R1133 B.n697 B.n51 68.9088
R1134 B.n697 B.n696 68.9088
R1135 B.n695 B.n58 68.9088
R1136 B.n689 B.n58 68.9088
R1137 B.n689 B.n688 68.9088
R1138 B.n688 B.n687 68.9088
R1139 B.n687 B.n65 68.9088
R1140 B.n681 B.n65 68.9088
R1141 B.n681 B.n680 68.9088
R1142 B.n680 B.n679 68.9088
R1143 B.n679 B.n72 68.9088
R1144 B.n673 B.n672 68.9088
R1145 B.n672 B.n671 68.9088
R1146 B.n671 B.n79 68.9088
R1147 B.n665 B.n79 68.9088
R1148 B.n665 B.n664 68.9088
R1149 B.n664 B.n663 68.9088
R1150 B.n436 B.t6 64.8554
R1151 B.t1 B.n719 64.8554
R1152 B.n102 B.n101 59.5399
R1153 B.n596 B.n108 59.5399
R1154 B.n286 B.n229 59.5399
R1155 B.n304 B.n223 59.5399
R1156 B.t5 B.n172 56.7485
R1157 B.n696 B.t8 56.7485
R1158 B.n129 B.t0 48.6417
R1159 B.t2 B.n744 48.6417
R1160 B.n461 B.t3 46.615
R1161 B.n735 B.t7 46.615
R1162 B.n101 B.n100 42.0853
R1163 B.n108 B.n107 42.0853
R1164 B.n229 B.n228 42.0853
R1165 B.n223 B.n222 42.0853
R1166 B.n370 B.t11 40.5348
R1167 B.n673 B.t15 40.5348
R1168 B.n418 B.t9 38.5081
R1169 B.n705 B.t4 38.5081
R1170 B.n350 B.n349 31.6883
R1171 B.n354 B.n206 31.6883
R1172 B.n550 B.n549 31.6883
R1173 B.n661 B.n660 31.6883
R1174 B.t9 B.n160 30.4012
R1175 B.t4 B.n44 30.4012
R1176 B.t11 B.n192 28.3745
R1177 B.t15 B.n72 28.3745
R1178 B.n454 B.t3 22.2944
R1179 B.n26 B.t7 22.2944
R1180 B.n480 B.t0 20.2677
R1181 B.n745 B.t2 20.2677
R1182 B B.n757 18.0485
R1183 B.n400 B.t5 12.1608
R1184 B.t8 B.n695 12.1608
R1185 B.n350 B.n202 10.6151
R1186 B.n360 B.n202 10.6151
R1187 B.n361 B.n360 10.6151
R1188 B.n362 B.n361 10.6151
R1189 B.n362 B.n194 10.6151
R1190 B.n372 B.n194 10.6151
R1191 B.n373 B.n372 10.6151
R1192 B.n374 B.n373 10.6151
R1193 B.n374 B.n186 10.6151
R1194 B.n384 B.n186 10.6151
R1195 B.n385 B.n384 10.6151
R1196 B.n386 B.n385 10.6151
R1197 B.n386 B.n178 10.6151
R1198 B.n396 B.n178 10.6151
R1199 B.n397 B.n396 10.6151
R1200 B.n398 B.n397 10.6151
R1201 B.n398 B.n170 10.6151
R1202 B.n408 B.n170 10.6151
R1203 B.n409 B.n408 10.6151
R1204 B.n410 B.n409 10.6151
R1205 B.n410 B.n162 10.6151
R1206 B.n420 B.n162 10.6151
R1207 B.n421 B.n420 10.6151
R1208 B.n422 B.n421 10.6151
R1209 B.n422 B.n154 10.6151
R1210 B.n432 B.n154 10.6151
R1211 B.n433 B.n432 10.6151
R1212 B.n434 B.n433 10.6151
R1213 B.n434 B.n146 10.6151
R1214 B.n444 B.n146 10.6151
R1215 B.n445 B.n444 10.6151
R1216 B.n446 B.n445 10.6151
R1217 B.n446 B.n138 10.6151
R1218 B.n457 B.n138 10.6151
R1219 B.n458 B.n457 10.6151
R1220 B.n459 B.n458 10.6151
R1221 B.n459 B.n131 10.6151
R1222 B.n469 B.n131 10.6151
R1223 B.n470 B.n469 10.6151
R1224 B.n471 B.n470 10.6151
R1225 B.n471 B.n123 10.6151
R1226 B.n482 B.n123 10.6151
R1227 B.n483 B.n482 10.6151
R1228 B.n484 B.n483 10.6151
R1229 B.n484 B.n0 10.6151
R1230 B.n349 B.n348 10.6151
R1231 B.n348 B.n210 10.6151
R1232 B.n343 B.n210 10.6151
R1233 B.n343 B.n342 10.6151
R1234 B.n342 B.n212 10.6151
R1235 B.n337 B.n212 10.6151
R1236 B.n337 B.n336 10.6151
R1237 B.n336 B.n335 10.6151
R1238 B.n335 B.n214 10.6151
R1239 B.n329 B.n214 10.6151
R1240 B.n329 B.n328 10.6151
R1241 B.n328 B.n327 10.6151
R1242 B.n327 B.n216 10.6151
R1243 B.n321 B.n216 10.6151
R1244 B.n321 B.n320 10.6151
R1245 B.n320 B.n319 10.6151
R1246 B.n319 B.n218 10.6151
R1247 B.n313 B.n218 10.6151
R1248 B.n313 B.n312 10.6151
R1249 B.n312 B.n311 10.6151
R1250 B.n311 B.n220 10.6151
R1251 B.n305 B.n220 10.6151
R1252 B.n303 B.n302 10.6151
R1253 B.n302 B.n224 10.6151
R1254 B.n296 B.n224 10.6151
R1255 B.n296 B.n295 10.6151
R1256 B.n295 B.n294 10.6151
R1257 B.n294 B.n226 10.6151
R1258 B.n288 B.n226 10.6151
R1259 B.n288 B.n287 10.6151
R1260 B.n285 B.n230 10.6151
R1261 B.n279 B.n230 10.6151
R1262 B.n279 B.n278 10.6151
R1263 B.n278 B.n277 10.6151
R1264 B.n277 B.n232 10.6151
R1265 B.n271 B.n232 10.6151
R1266 B.n271 B.n270 10.6151
R1267 B.n270 B.n269 10.6151
R1268 B.n269 B.n234 10.6151
R1269 B.n263 B.n234 10.6151
R1270 B.n263 B.n262 10.6151
R1271 B.n262 B.n261 10.6151
R1272 B.n261 B.n236 10.6151
R1273 B.n255 B.n236 10.6151
R1274 B.n255 B.n254 10.6151
R1275 B.n254 B.n253 10.6151
R1276 B.n253 B.n238 10.6151
R1277 B.n247 B.n238 10.6151
R1278 B.n247 B.n246 10.6151
R1279 B.n246 B.n245 10.6151
R1280 B.n245 B.n240 10.6151
R1281 B.n240 B.n206 10.6151
R1282 B.n355 B.n354 10.6151
R1283 B.n356 B.n355 10.6151
R1284 B.n356 B.n198 10.6151
R1285 B.n366 B.n198 10.6151
R1286 B.n367 B.n366 10.6151
R1287 B.n368 B.n367 10.6151
R1288 B.n368 B.n190 10.6151
R1289 B.n378 B.n190 10.6151
R1290 B.n379 B.n378 10.6151
R1291 B.n380 B.n379 10.6151
R1292 B.n380 B.n182 10.6151
R1293 B.n390 B.n182 10.6151
R1294 B.n391 B.n390 10.6151
R1295 B.n392 B.n391 10.6151
R1296 B.n392 B.n174 10.6151
R1297 B.n402 B.n174 10.6151
R1298 B.n403 B.n402 10.6151
R1299 B.n404 B.n403 10.6151
R1300 B.n404 B.n166 10.6151
R1301 B.n414 B.n166 10.6151
R1302 B.n415 B.n414 10.6151
R1303 B.n416 B.n415 10.6151
R1304 B.n416 B.n158 10.6151
R1305 B.n426 B.n158 10.6151
R1306 B.n427 B.n426 10.6151
R1307 B.n428 B.n427 10.6151
R1308 B.n428 B.n150 10.6151
R1309 B.n438 B.n150 10.6151
R1310 B.n439 B.n438 10.6151
R1311 B.n440 B.n439 10.6151
R1312 B.n440 B.n142 10.6151
R1313 B.n450 B.n142 10.6151
R1314 B.n451 B.n450 10.6151
R1315 B.n452 B.n451 10.6151
R1316 B.n452 B.n135 10.6151
R1317 B.n463 B.n135 10.6151
R1318 B.n464 B.n463 10.6151
R1319 B.n465 B.n464 10.6151
R1320 B.n465 B.n126 10.6151
R1321 B.n475 B.n126 10.6151
R1322 B.n476 B.n475 10.6151
R1323 B.n478 B.n476 10.6151
R1324 B.n478 B.n477 10.6151
R1325 B.n477 B.n119 10.6151
R1326 B.n489 B.n119 10.6151
R1327 B.n490 B.n489 10.6151
R1328 B.n491 B.n490 10.6151
R1329 B.n492 B.n491 10.6151
R1330 B.n493 B.n492 10.6151
R1331 B.n496 B.n493 10.6151
R1332 B.n497 B.n496 10.6151
R1333 B.n498 B.n497 10.6151
R1334 B.n499 B.n498 10.6151
R1335 B.n501 B.n499 10.6151
R1336 B.n502 B.n501 10.6151
R1337 B.n503 B.n502 10.6151
R1338 B.n504 B.n503 10.6151
R1339 B.n506 B.n504 10.6151
R1340 B.n507 B.n506 10.6151
R1341 B.n508 B.n507 10.6151
R1342 B.n509 B.n508 10.6151
R1343 B.n511 B.n509 10.6151
R1344 B.n512 B.n511 10.6151
R1345 B.n513 B.n512 10.6151
R1346 B.n514 B.n513 10.6151
R1347 B.n516 B.n514 10.6151
R1348 B.n517 B.n516 10.6151
R1349 B.n518 B.n517 10.6151
R1350 B.n519 B.n518 10.6151
R1351 B.n521 B.n519 10.6151
R1352 B.n522 B.n521 10.6151
R1353 B.n523 B.n522 10.6151
R1354 B.n524 B.n523 10.6151
R1355 B.n526 B.n524 10.6151
R1356 B.n527 B.n526 10.6151
R1357 B.n528 B.n527 10.6151
R1358 B.n529 B.n528 10.6151
R1359 B.n531 B.n529 10.6151
R1360 B.n532 B.n531 10.6151
R1361 B.n533 B.n532 10.6151
R1362 B.n534 B.n533 10.6151
R1363 B.n536 B.n534 10.6151
R1364 B.n537 B.n536 10.6151
R1365 B.n538 B.n537 10.6151
R1366 B.n539 B.n538 10.6151
R1367 B.n541 B.n539 10.6151
R1368 B.n542 B.n541 10.6151
R1369 B.n543 B.n542 10.6151
R1370 B.n544 B.n543 10.6151
R1371 B.n546 B.n544 10.6151
R1372 B.n547 B.n546 10.6151
R1373 B.n548 B.n547 10.6151
R1374 B.n549 B.n548 10.6151
R1375 B.n749 B.n1 10.6151
R1376 B.n749 B.n748 10.6151
R1377 B.n748 B.n747 10.6151
R1378 B.n747 B.n10 10.6151
R1379 B.n741 B.n10 10.6151
R1380 B.n741 B.n740 10.6151
R1381 B.n740 B.n739 10.6151
R1382 B.n739 B.n18 10.6151
R1383 B.n733 B.n18 10.6151
R1384 B.n733 B.n732 10.6151
R1385 B.n732 B.n731 10.6151
R1386 B.n731 B.n24 10.6151
R1387 B.n725 B.n24 10.6151
R1388 B.n725 B.n724 10.6151
R1389 B.n724 B.n723 10.6151
R1390 B.n723 B.n32 10.6151
R1391 B.n717 B.n32 10.6151
R1392 B.n717 B.n716 10.6151
R1393 B.n716 B.n715 10.6151
R1394 B.n715 B.n39 10.6151
R1395 B.n709 B.n39 10.6151
R1396 B.n709 B.n708 10.6151
R1397 B.n708 B.n707 10.6151
R1398 B.n707 B.n46 10.6151
R1399 B.n701 B.n46 10.6151
R1400 B.n701 B.n700 10.6151
R1401 B.n700 B.n699 10.6151
R1402 B.n699 B.n53 10.6151
R1403 B.n693 B.n53 10.6151
R1404 B.n693 B.n692 10.6151
R1405 B.n692 B.n691 10.6151
R1406 B.n691 B.n60 10.6151
R1407 B.n685 B.n60 10.6151
R1408 B.n685 B.n684 10.6151
R1409 B.n684 B.n683 10.6151
R1410 B.n683 B.n67 10.6151
R1411 B.n677 B.n67 10.6151
R1412 B.n677 B.n676 10.6151
R1413 B.n676 B.n675 10.6151
R1414 B.n675 B.n74 10.6151
R1415 B.n669 B.n74 10.6151
R1416 B.n669 B.n668 10.6151
R1417 B.n668 B.n667 10.6151
R1418 B.n667 B.n81 10.6151
R1419 B.n661 B.n81 10.6151
R1420 B.n660 B.n659 10.6151
R1421 B.n659 B.n88 10.6151
R1422 B.n653 B.n88 10.6151
R1423 B.n653 B.n652 10.6151
R1424 B.n652 B.n651 10.6151
R1425 B.n651 B.n90 10.6151
R1426 B.n645 B.n90 10.6151
R1427 B.n645 B.n644 10.6151
R1428 B.n644 B.n643 10.6151
R1429 B.n643 B.n92 10.6151
R1430 B.n637 B.n92 10.6151
R1431 B.n637 B.n636 10.6151
R1432 B.n636 B.n635 10.6151
R1433 B.n635 B.n94 10.6151
R1434 B.n629 B.n94 10.6151
R1435 B.n629 B.n628 10.6151
R1436 B.n628 B.n627 10.6151
R1437 B.n627 B.n96 10.6151
R1438 B.n621 B.n96 10.6151
R1439 B.n621 B.n620 10.6151
R1440 B.n620 B.n619 10.6151
R1441 B.n619 B.n98 10.6151
R1442 B.n613 B.n612 10.6151
R1443 B.n612 B.n611 10.6151
R1444 B.n611 B.n103 10.6151
R1445 B.n605 B.n103 10.6151
R1446 B.n605 B.n604 10.6151
R1447 B.n604 B.n603 10.6151
R1448 B.n603 B.n105 10.6151
R1449 B.n597 B.n105 10.6151
R1450 B.n595 B.n594 10.6151
R1451 B.n594 B.n109 10.6151
R1452 B.n588 B.n109 10.6151
R1453 B.n588 B.n587 10.6151
R1454 B.n587 B.n586 10.6151
R1455 B.n586 B.n111 10.6151
R1456 B.n580 B.n111 10.6151
R1457 B.n580 B.n579 10.6151
R1458 B.n579 B.n578 10.6151
R1459 B.n578 B.n113 10.6151
R1460 B.n572 B.n113 10.6151
R1461 B.n572 B.n571 10.6151
R1462 B.n571 B.n570 10.6151
R1463 B.n570 B.n115 10.6151
R1464 B.n564 B.n115 10.6151
R1465 B.n564 B.n563 10.6151
R1466 B.n563 B.n562 10.6151
R1467 B.n562 B.n117 10.6151
R1468 B.n556 B.n117 10.6151
R1469 B.n556 B.n555 10.6151
R1470 B.n555 B.n554 10.6151
R1471 B.n554 B.n550 10.6151
R1472 B.n757 B.n0 8.11757
R1473 B.n757 B.n1 8.11757
R1474 B.n304 B.n303 6.5566
R1475 B.n287 B.n286 6.5566
R1476 B.n613 B.n102 6.5566
R1477 B.n597 B.n596 6.5566
R1478 B.n305 B.n304 4.05904
R1479 B.n286 B.n285 4.05904
R1480 B.n102 B.n98 4.05904
R1481 B.n596 B.n595 4.05904
R1482 B.t6 B.n148 4.05393
R1483 B.n720 B.t1 4.05393
R1484 VP.n42 VP.n9 181.465
R1485 VP.n74 VP.n73 181.465
R1486 VP.n41 VP.n40 181.465
R1487 VP.n19 VP.n16 161.3
R1488 VP.n21 VP.n20 161.3
R1489 VP.n22 VP.n15 161.3
R1490 VP.n24 VP.n23 161.3
R1491 VP.n26 VP.n14 161.3
R1492 VP.n28 VP.n27 161.3
R1493 VP.n29 VP.n13 161.3
R1494 VP.n31 VP.n30 161.3
R1495 VP.n33 VP.n12 161.3
R1496 VP.n35 VP.n34 161.3
R1497 VP.n36 VP.n11 161.3
R1498 VP.n38 VP.n37 161.3
R1499 VP.n39 VP.n10 161.3
R1500 VP.n72 VP.n0 161.3
R1501 VP.n71 VP.n70 161.3
R1502 VP.n69 VP.n1 161.3
R1503 VP.n68 VP.n67 161.3
R1504 VP.n66 VP.n2 161.3
R1505 VP.n64 VP.n63 161.3
R1506 VP.n62 VP.n3 161.3
R1507 VP.n61 VP.n60 161.3
R1508 VP.n59 VP.n4 161.3
R1509 VP.n57 VP.n56 161.3
R1510 VP.n55 VP.n5 161.3
R1511 VP.n54 VP.n53 161.3
R1512 VP.n52 VP.n6 161.3
R1513 VP.n50 VP.n49 161.3
R1514 VP.n48 VP.n7 161.3
R1515 VP.n47 VP.n46 161.3
R1516 VP.n45 VP.n8 161.3
R1517 VP.n44 VP.n43 161.3
R1518 VP.n17 VP.t8 107.987
R1519 VP.n9 VP.t3 73.0864
R1520 VP.n51 VP.t7 73.0864
R1521 VP.n58 VP.t9 73.0864
R1522 VP.n65 VP.t2 73.0864
R1523 VP.n73 VP.t6 73.0864
R1524 VP.n40 VP.t5 73.0864
R1525 VP.n32 VP.t0 73.0864
R1526 VP.n25 VP.t1 73.0864
R1527 VP.n18 VP.t4 73.0864
R1528 VP.n53 VP.n5 56.5617
R1529 VP.n60 VP.n3 56.5617
R1530 VP.n27 VP.n13 56.5617
R1531 VP.n20 VP.n15 56.5617
R1532 VP.n18 VP.n17 48.9423
R1533 VP.n42 VP.n41 44.0422
R1534 VP.n46 VP.n45 41.0614
R1535 VP.n71 VP.n1 41.0614
R1536 VP.n38 VP.n11 41.0614
R1537 VP.n46 VP.n7 40.0926
R1538 VP.n67 VP.n1 40.0926
R1539 VP.n34 VP.n11 40.0926
R1540 VP.n45 VP.n44 24.5923
R1541 VP.n50 VP.n7 24.5923
R1542 VP.n53 VP.n52 24.5923
R1543 VP.n57 VP.n5 24.5923
R1544 VP.n60 VP.n59 24.5923
R1545 VP.n64 VP.n3 24.5923
R1546 VP.n67 VP.n66 24.5923
R1547 VP.n72 VP.n71 24.5923
R1548 VP.n39 VP.n38 24.5923
R1549 VP.n31 VP.n13 24.5923
R1550 VP.n34 VP.n33 24.5923
R1551 VP.n24 VP.n15 24.5923
R1552 VP.n27 VP.n26 24.5923
R1553 VP.n20 VP.n19 24.5923
R1554 VP.n52 VP.n51 20.6576
R1555 VP.n65 VP.n64 20.6576
R1556 VP.n32 VP.n31 20.6576
R1557 VP.n19 VP.n18 20.6576
R1558 VP.n58 VP.n57 12.2964
R1559 VP.n59 VP.n58 12.2964
R1560 VP.n25 VP.n24 12.2964
R1561 VP.n26 VP.n25 12.2964
R1562 VP.n17 VP.n16 12.2243
R1563 VP.n44 VP.n9 4.42703
R1564 VP.n73 VP.n72 4.42703
R1565 VP.n40 VP.n39 4.42703
R1566 VP.n51 VP.n50 3.93519
R1567 VP.n66 VP.n65 3.93519
R1568 VP.n33 VP.n32 3.93519
R1569 VP.n21 VP.n16 0.189894
R1570 VP.n22 VP.n21 0.189894
R1571 VP.n23 VP.n22 0.189894
R1572 VP.n23 VP.n14 0.189894
R1573 VP.n28 VP.n14 0.189894
R1574 VP.n29 VP.n28 0.189894
R1575 VP.n30 VP.n29 0.189894
R1576 VP.n30 VP.n12 0.189894
R1577 VP.n35 VP.n12 0.189894
R1578 VP.n36 VP.n35 0.189894
R1579 VP.n37 VP.n36 0.189894
R1580 VP.n37 VP.n10 0.189894
R1581 VP.n41 VP.n10 0.189894
R1582 VP.n43 VP.n42 0.189894
R1583 VP.n43 VP.n8 0.189894
R1584 VP.n47 VP.n8 0.189894
R1585 VP.n48 VP.n47 0.189894
R1586 VP.n49 VP.n48 0.189894
R1587 VP.n49 VP.n6 0.189894
R1588 VP.n54 VP.n6 0.189894
R1589 VP.n55 VP.n54 0.189894
R1590 VP.n56 VP.n55 0.189894
R1591 VP.n56 VP.n4 0.189894
R1592 VP.n61 VP.n4 0.189894
R1593 VP.n62 VP.n61 0.189894
R1594 VP.n63 VP.n62 0.189894
R1595 VP.n63 VP.n2 0.189894
R1596 VP.n68 VP.n2 0.189894
R1597 VP.n69 VP.n68 0.189894
R1598 VP.n70 VP.n69 0.189894
R1599 VP.n70 VP.n0 0.189894
R1600 VP.n74 VP.n0 0.189894
R1601 VP VP.n74 0.0516364
R1602 VDD1.n1 VDD1.t1 72.1255
R1603 VDD1.n3 VDD1.t6 72.1252
R1604 VDD1.n5 VDD1.n4 68.0538
R1605 VDD1.n1 VDD1.n0 66.7064
R1606 VDD1.n7 VDD1.n6 66.7062
R1607 VDD1.n3 VDD1.n2 66.7062
R1608 VDD1.n7 VDD1.n5 38.9298
R1609 VDD1.n6 VDD1.t9 3.54889
R1610 VDD1.n6 VDD1.t4 3.54889
R1611 VDD1.n0 VDD1.t5 3.54889
R1612 VDD1.n0 VDD1.t8 3.54889
R1613 VDD1.n4 VDD1.t7 3.54889
R1614 VDD1.n4 VDD1.t3 3.54889
R1615 VDD1.n2 VDD1.t2 3.54889
R1616 VDD1.n2 VDD1.t0 3.54889
R1617 VDD1 VDD1.n7 1.34533
R1618 VDD1 VDD1.n1 0.526362
R1619 VDD1.n5 VDD1.n3 0.412826
C0 VN VTAIL 5.59174f
C1 VP VDD1 5.17405f
C2 VP VTAIL 5.60597f
C3 VN VDD2 4.84216f
C4 VP VDD2 0.486215f
C5 VTAIL VDD1 6.99299f
C6 VDD2 VDD1 1.67796f
C7 VTAIL VDD2 7.03983f
C8 VP VN 6.081759f
C9 VN VDD1 0.151801f
C10 VDD2 B 5.157974f
C11 VDD1 B 5.141833f
C12 VTAIL B 4.763389f
C13 VN B 13.849641f
C14 VP B 12.380272f
C15 VDD1.t1 B 1.07936f
C16 VDD1.t5 B 0.101992f
C17 VDD1.t8 B 0.101992f
C18 VDD1.n0 B 0.842628f
C19 VDD1.n1 B 0.74217f
C20 VDD1.t6 B 1.07936f
C21 VDD1.t2 B 0.101992f
C22 VDD1.t0 B 0.101992f
C23 VDD1.n2 B 0.842624f
C24 VDD1.n3 B 0.735015f
C25 VDD1.t7 B 0.101992f
C26 VDD1.t3 B 0.101992f
C27 VDD1.n4 B 0.851264f
C28 VDD1.n5 B 2.05139f
C29 VDD1.t9 B 0.101992f
C30 VDD1.t4 B 0.101992f
C31 VDD1.n6 B 0.842624f
C32 VDD1.n7 B 2.1782f
C33 VP.n0 B 0.02982f
C34 VP.t6 B 0.806776f
C35 VP.n1 B 0.024094f
C36 VP.n2 B 0.02982f
C37 VP.t2 B 0.806776f
C38 VP.n3 B 0.036335f
C39 VP.n4 B 0.02982f
C40 VP.t9 B 0.806776f
C41 VP.n5 B 0.050361f
C42 VP.n6 B 0.02982f
C43 VP.t7 B 0.806776f
C44 VP.n7 B 0.059098f
C45 VP.n8 B 0.02982f
C46 VP.t3 B 0.806776f
C47 VP.n9 B 0.383333f
C48 VP.n10 B 0.02982f
C49 VP.t5 B 0.806776f
C50 VP.n11 B 0.024094f
C51 VP.n12 B 0.02982f
C52 VP.t0 B 0.806776f
C53 VP.n13 B 0.036335f
C54 VP.n14 B 0.02982f
C55 VP.t1 B 0.806776f
C56 VP.n15 B 0.050361f
C57 VP.n16 B 0.220877f
C58 VP.t4 B 0.806776f
C59 VP.t8 B 0.9543f
C60 VP.n17 B 0.373093f
C61 VP.n18 B 0.389481f
C62 VP.n19 B 0.050931f
C63 VP.n20 B 0.036335f
C64 VP.n21 B 0.02982f
C65 VP.n22 B 0.02982f
C66 VP.n23 B 0.02982f
C67 VP.n24 B 0.041649f
C68 VP.n25 B 0.31331f
C69 VP.n26 B 0.041649f
C70 VP.n27 B 0.050361f
C71 VP.n28 B 0.02982f
C72 VP.n29 B 0.02982f
C73 VP.n30 B 0.02982f
C74 VP.n31 B 0.050931f
C75 VP.n32 B 0.31331f
C76 VP.n33 B 0.032367f
C77 VP.n34 B 0.059098f
C78 VP.n35 B 0.02982f
C79 VP.n36 B 0.02982f
C80 VP.n37 B 0.02982f
C81 VP.n38 B 0.058803f
C82 VP.n39 B 0.032913f
C83 VP.n40 B 0.383333f
C84 VP.n41 B 1.33932f
C85 VP.n42 B 1.36373f
C86 VP.n43 B 0.02982f
C87 VP.n44 B 0.032913f
C88 VP.n45 B 0.058803f
C89 VP.n46 B 0.024094f
C90 VP.n47 B 0.02982f
C91 VP.n48 B 0.02982f
C92 VP.n49 B 0.02982f
C93 VP.n50 B 0.032367f
C94 VP.n51 B 0.31331f
C95 VP.n52 B 0.050931f
C96 VP.n53 B 0.036335f
C97 VP.n54 B 0.02982f
C98 VP.n55 B 0.02982f
C99 VP.n56 B 0.02982f
C100 VP.n57 B 0.041649f
C101 VP.n58 B 0.31331f
C102 VP.n59 B 0.041649f
C103 VP.n60 B 0.050361f
C104 VP.n61 B 0.02982f
C105 VP.n62 B 0.02982f
C106 VP.n63 B 0.02982f
C107 VP.n64 B 0.050931f
C108 VP.n65 B 0.31331f
C109 VP.n66 B 0.032367f
C110 VP.n67 B 0.059098f
C111 VP.n68 B 0.02982f
C112 VP.n69 B 0.02982f
C113 VP.n70 B 0.02982f
C114 VP.n71 B 0.058803f
C115 VP.n72 B 0.032913f
C116 VP.n73 B 0.383333f
C117 VP.n74 B 0.031864f
C118 VTAIL.t18 B 0.122998f
C119 VTAIL.t13 B 0.122998f
C120 VTAIL.n0 B 0.942878f
C121 VTAIL.n1 B 0.518165f
C122 VTAIL.t0 B 1.20181f
C123 VTAIL.n2 B 0.631489f
C124 VTAIL.t6 B 0.122998f
C125 VTAIL.t3 B 0.122998f
C126 VTAIL.n3 B 0.942878f
C127 VTAIL.n4 B 0.596811f
C128 VTAIL.t5 B 0.122998f
C129 VTAIL.t9 B 0.122998f
C130 VTAIL.n5 B 0.942878f
C131 VTAIL.n6 B 1.57621f
C132 VTAIL.t10 B 0.122998f
C133 VTAIL.t17 B 0.122998f
C134 VTAIL.n7 B 0.942883f
C135 VTAIL.n8 B 1.57621f
C136 VTAIL.t14 B 0.122998f
C137 VTAIL.t15 B 0.122998f
C138 VTAIL.n9 B 0.942883f
C139 VTAIL.n10 B 0.596805f
C140 VTAIL.t12 B 1.20181f
C141 VTAIL.n11 B 0.631484f
C142 VTAIL.t2 B 0.122998f
C143 VTAIL.t7 B 0.122998f
C144 VTAIL.n12 B 0.942883f
C145 VTAIL.n13 B 0.554964f
C146 VTAIL.t1 B 0.122998f
C147 VTAIL.t4 B 0.122998f
C148 VTAIL.n14 B 0.942883f
C149 VTAIL.n15 B 0.596805f
C150 VTAIL.t8 B 1.20181f
C151 VTAIL.n16 B 1.48459f
C152 VTAIL.t11 B 1.20181f
C153 VTAIL.n17 B 1.48459f
C154 VTAIL.t16 B 0.122998f
C155 VTAIL.t19 B 0.122998f
C156 VTAIL.n18 B 0.942878f
C157 VTAIL.n19 B 0.465476f
C158 VDD2.t2 B 1.05133f
C159 VDD2.t6 B 0.099344f
C160 VDD2.t8 B 0.099344f
C161 VDD2.n0 B 0.820745f
C162 VDD2.n1 B 0.71593f
C163 VDD2.t4 B 0.099344f
C164 VDD2.t7 B 0.099344f
C165 VDD2.n2 B 0.82916f
C166 VDD2.n3 B 1.9075f
C167 VDD2.t0 B 1.04156f
C168 VDD2.n4 B 2.08154f
C169 VDD2.t9 B 0.099344f
C170 VDD2.t5 B 0.099344f
C171 VDD2.n5 B 0.820748f
C172 VDD2.n6 B 0.355826f
C173 VDD2.t1 B 0.099344f
C174 VDD2.t3 B 0.099344f
C175 VDD2.n7 B 0.82913f
C176 VN.n0 B 0.029042f
C177 VN.t8 B 0.785732f
C178 VN.n1 B 0.023466f
C179 VN.n2 B 0.029042f
C180 VN.t0 B 0.785732f
C181 VN.n3 B 0.035388f
C182 VN.n4 B 0.029042f
C183 VN.t3 B 0.785732f
C184 VN.n5 B 0.049047f
C185 VN.n6 B 0.215116f
C186 VN.t6 B 0.785732f
C187 VN.t1 B 0.929408f
C188 VN.n7 B 0.363361f
C189 VN.n8 B 0.379321f
C190 VN.n9 B 0.049602f
C191 VN.n10 B 0.035388f
C192 VN.n11 B 0.029042f
C193 VN.n12 B 0.029042f
C194 VN.n13 B 0.029042f
C195 VN.n14 B 0.040563f
C196 VN.n15 B 0.305138f
C197 VN.n16 B 0.040563f
C198 VN.n17 B 0.049047f
C199 VN.n18 B 0.029042f
C200 VN.n19 B 0.029042f
C201 VN.n20 B 0.029042f
C202 VN.n21 B 0.049602f
C203 VN.n22 B 0.305138f
C204 VN.n23 B 0.031523f
C205 VN.n24 B 0.057557f
C206 VN.n25 B 0.029042f
C207 VN.n26 B 0.029042f
C208 VN.n27 B 0.029042f
C209 VN.n28 B 0.057269f
C210 VN.n29 B 0.032055f
C211 VN.n30 B 0.373334f
C212 VN.n31 B 0.031032f
C213 VN.n32 B 0.029042f
C214 VN.t9 B 0.785732f
C215 VN.n33 B 0.023466f
C216 VN.n34 B 0.029042f
C217 VN.t2 B 0.785732f
C218 VN.n35 B 0.035388f
C219 VN.n36 B 0.029042f
C220 VN.t5 B 0.785732f
C221 VN.n37 B 0.049047f
C222 VN.n38 B 0.215116f
C223 VN.t4 B 0.785732f
C224 VN.t7 B 0.929408f
C225 VN.n39 B 0.363361f
C226 VN.n40 B 0.379321f
C227 VN.n41 B 0.049602f
C228 VN.n42 B 0.035388f
C229 VN.n43 B 0.029042f
C230 VN.n44 B 0.029042f
C231 VN.n45 B 0.029042f
C232 VN.n46 B 0.040563f
C233 VN.n47 B 0.305138f
C234 VN.n48 B 0.040563f
C235 VN.n49 B 0.049047f
C236 VN.n50 B 0.029042f
C237 VN.n51 B 0.029042f
C238 VN.n52 B 0.029042f
C239 VN.n53 B 0.049602f
C240 VN.n54 B 0.305138f
C241 VN.n55 B 0.031523f
C242 VN.n56 B 0.057557f
C243 VN.n57 B 0.029042f
C244 VN.n58 B 0.029042f
C245 VN.n59 B 0.029042f
C246 VN.n60 B 0.057269f
C247 VN.n61 B 0.032055f
C248 VN.n62 B 0.373334f
C249 VN.n63 B 1.3234f
.ends

