* NGSPICE file created from diff_pair_sample_0971.ext - technology: sky130A

.subckt diff_pair_sample_0971 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=3.64
X1 VDD1.t3 VP.t0 VTAIL.t1 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=3.64
X2 B.t11 B.t9 B.t10 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=3.64
X3 VTAIL.t0 VP.t1 VDD1.t2 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=3.64
X4 B.t8 B.t6 B.t7 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=3.64
X5 VTAIL.t2 VP.t2 VDD1.t1 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=3.64
X6 VDD2.t2 VN.t1 VTAIL.t6 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=3.64
X7 B.t5 B.t3 B.t4 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=3.64
X8 VDD2.t1 VN.t2 VTAIL.t5 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=3.64
X9 VDD1.t0 VP.t3 VTAIL.t3 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=3.64
X10 B.t2 B.t0 B.t1 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=3.64
X11 VTAIL.t4 VN.t3 VDD2.t3 w_n3352_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=3.64
R0 VN.n1 VN.t1 54.1564
R1 VN.n0 VN.t3 54.1564
R2 VN.n0 VN.t2 52.9026
R3 VN.n1 VN.t0 52.9026
R4 VN VN.n1 44.9491
R5 VN VN.n0 2.05897
R6 VDD2.n2 VDD2.n0 177.065
R7 VDD2.n2 VDD2.n1 140.591
R8 VDD2.n1 VDD2.t0 11.2479
R9 VDD2.n1 VDD2.t2 11.2479
R10 VDD2.n0 VDD2.t3 11.2479
R11 VDD2.n0 VDD2.t1 11.2479
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t0 135.161
R14 VTAIL.n4 VTAIL.t6 135.161
R15 VTAIL.n3 VTAIL.t7 135.161
R16 VTAIL.n6 VTAIL.t3 135.16
R17 VTAIL.n7 VTAIL.t5 135.16
R18 VTAIL.n0 VTAIL.t4 135.16
R19 VTAIL.n1 VTAIL.t1 135.16
R20 VTAIL.n2 VTAIL.t2 135.16
R21 VTAIL.n7 VTAIL.n6 18.2807
R22 VTAIL.n3 VTAIL.n2 18.2807
R23 VTAIL.n4 VTAIL.n3 3.42291
R24 VTAIL.n6 VTAIL.n5 3.42291
R25 VTAIL.n2 VTAIL.n1 3.42291
R26 VTAIL VTAIL.n0 1.7699
R27 VTAIL VTAIL.n7 1.65352
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 VP.n19 VP.n18 161.3
R31 VP.n17 VP.n1 161.3
R32 VP.n16 VP.n15 161.3
R33 VP.n14 VP.n2 161.3
R34 VP.n13 VP.n12 161.3
R35 VP.n11 VP.n3 161.3
R36 VP.n10 VP.n9 161.3
R37 VP.n8 VP.n4 161.3
R38 VP.n7 VP.n6 78.5679
R39 VP.n20 VP.n0 78.5679
R40 VP.n12 VP.n2 56.5193
R41 VP.n5 VP.t1 54.1562
R42 VP.n5 VP.t3 52.9026
R43 VP.n7 VP.n5 44.7838
R44 VP.n10 VP.n4 24.4675
R45 VP.n11 VP.n10 24.4675
R46 VP.n12 VP.n11 24.4675
R47 VP.n16 VP.n2 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n6 VP.t2 19.1348
R51 VP.n0 VP.t0 19.1348
R52 VP.n6 VP.n4 11.5
R53 VP.n18 VP.n0 11.5
R54 VP.n8 VP.n7 0.354971
R55 VP.n20 VP.n19 0.354971
R56 VP VP.n20 0.26696
R57 VP.n9 VP.n8 0.189894
R58 VP.n9 VP.n3 0.189894
R59 VP.n13 VP.n3 0.189894
R60 VP.n14 VP.n13 0.189894
R61 VP.n15 VP.n14 0.189894
R62 VP.n15 VP.n1 0.189894
R63 VP.n19 VP.n1 0.189894
R64 VDD1 VDD1.n1 177.589
R65 VDD1 VDD1.n0 140.649
R66 VDD1.n0 VDD1.t2 11.2479
R67 VDD1.n0 VDD1.t0 11.2479
R68 VDD1.n1 VDD1.t1 11.2479
R69 VDD1.n1 VDD1.t3 11.2479
R70 B.n390 B.n389 585
R71 B.n391 B.n46 585
R72 B.n393 B.n392 585
R73 B.n394 B.n45 585
R74 B.n396 B.n395 585
R75 B.n397 B.n44 585
R76 B.n399 B.n398 585
R77 B.n400 B.n43 585
R78 B.n402 B.n401 585
R79 B.n403 B.n42 585
R80 B.n405 B.n404 585
R81 B.n406 B.n41 585
R82 B.n408 B.n407 585
R83 B.n409 B.n40 585
R84 B.n411 B.n410 585
R85 B.n413 B.n37 585
R86 B.n415 B.n414 585
R87 B.n416 B.n36 585
R88 B.n418 B.n417 585
R89 B.n419 B.n35 585
R90 B.n421 B.n420 585
R91 B.n422 B.n34 585
R92 B.n424 B.n423 585
R93 B.n425 B.n31 585
R94 B.n428 B.n427 585
R95 B.n429 B.n30 585
R96 B.n431 B.n430 585
R97 B.n432 B.n29 585
R98 B.n434 B.n433 585
R99 B.n435 B.n28 585
R100 B.n437 B.n436 585
R101 B.n438 B.n27 585
R102 B.n440 B.n439 585
R103 B.n441 B.n26 585
R104 B.n443 B.n442 585
R105 B.n444 B.n25 585
R106 B.n446 B.n445 585
R107 B.n447 B.n24 585
R108 B.n449 B.n448 585
R109 B.n388 B.n47 585
R110 B.n387 B.n386 585
R111 B.n385 B.n48 585
R112 B.n384 B.n383 585
R113 B.n382 B.n49 585
R114 B.n381 B.n380 585
R115 B.n379 B.n50 585
R116 B.n378 B.n377 585
R117 B.n376 B.n51 585
R118 B.n375 B.n374 585
R119 B.n373 B.n52 585
R120 B.n372 B.n371 585
R121 B.n370 B.n53 585
R122 B.n369 B.n368 585
R123 B.n367 B.n54 585
R124 B.n366 B.n365 585
R125 B.n364 B.n55 585
R126 B.n363 B.n362 585
R127 B.n361 B.n56 585
R128 B.n360 B.n359 585
R129 B.n358 B.n57 585
R130 B.n357 B.n356 585
R131 B.n355 B.n58 585
R132 B.n354 B.n353 585
R133 B.n352 B.n59 585
R134 B.n351 B.n350 585
R135 B.n349 B.n60 585
R136 B.n348 B.n347 585
R137 B.n346 B.n61 585
R138 B.n345 B.n344 585
R139 B.n343 B.n62 585
R140 B.n342 B.n341 585
R141 B.n340 B.n63 585
R142 B.n339 B.n338 585
R143 B.n337 B.n64 585
R144 B.n336 B.n335 585
R145 B.n334 B.n65 585
R146 B.n333 B.n332 585
R147 B.n331 B.n66 585
R148 B.n330 B.n329 585
R149 B.n328 B.n67 585
R150 B.n327 B.n326 585
R151 B.n325 B.n68 585
R152 B.n324 B.n323 585
R153 B.n322 B.n69 585
R154 B.n321 B.n320 585
R155 B.n319 B.n70 585
R156 B.n318 B.n317 585
R157 B.n316 B.n71 585
R158 B.n315 B.n314 585
R159 B.n313 B.n72 585
R160 B.n312 B.n311 585
R161 B.n310 B.n73 585
R162 B.n309 B.n308 585
R163 B.n307 B.n74 585
R164 B.n306 B.n305 585
R165 B.n304 B.n75 585
R166 B.n303 B.n302 585
R167 B.n301 B.n76 585
R168 B.n300 B.n299 585
R169 B.n298 B.n77 585
R170 B.n297 B.n296 585
R171 B.n295 B.n78 585
R172 B.n294 B.n293 585
R173 B.n292 B.n79 585
R174 B.n291 B.n290 585
R175 B.n289 B.n80 585
R176 B.n288 B.n287 585
R177 B.n286 B.n81 585
R178 B.n285 B.n284 585
R179 B.n283 B.n82 585
R180 B.n282 B.n281 585
R181 B.n280 B.n83 585
R182 B.n279 B.n278 585
R183 B.n277 B.n84 585
R184 B.n276 B.n275 585
R185 B.n274 B.n85 585
R186 B.n273 B.n272 585
R187 B.n271 B.n86 585
R188 B.n270 B.n269 585
R189 B.n268 B.n87 585
R190 B.n267 B.n266 585
R191 B.n265 B.n88 585
R192 B.n264 B.n263 585
R193 B.n262 B.n89 585
R194 B.n261 B.n260 585
R195 B.n259 B.n90 585
R196 B.n199 B.n114 585
R197 B.n201 B.n200 585
R198 B.n202 B.n113 585
R199 B.n204 B.n203 585
R200 B.n205 B.n112 585
R201 B.n207 B.n206 585
R202 B.n208 B.n111 585
R203 B.n210 B.n209 585
R204 B.n211 B.n110 585
R205 B.n213 B.n212 585
R206 B.n214 B.n109 585
R207 B.n216 B.n215 585
R208 B.n217 B.n108 585
R209 B.n219 B.n218 585
R210 B.n220 B.n105 585
R211 B.n223 B.n222 585
R212 B.n224 B.n104 585
R213 B.n226 B.n225 585
R214 B.n227 B.n103 585
R215 B.n229 B.n228 585
R216 B.n230 B.n102 585
R217 B.n232 B.n231 585
R218 B.n233 B.n101 585
R219 B.n235 B.n234 585
R220 B.n237 B.n236 585
R221 B.n238 B.n97 585
R222 B.n240 B.n239 585
R223 B.n241 B.n96 585
R224 B.n243 B.n242 585
R225 B.n244 B.n95 585
R226 B.n246 B.n245 585
R227 B.n247 B.n94 585
R228 B.n249 B.n248 585
R229 B.n250 B.n93 585
R230 B.n252 B.n251 585
R231 B.n253 B.n92 585
R232 B.n255 B.n254 585
R233 B.n256 B.n91 585
R234 B.n258 B.n257 585
R235 B.n198 B.n197 585
R236 B.n196 B.n115 585
R237 B.n195 B.n194 585
R238 B.n193 B.n116 585
R239 B.n192 B.n191 585
R240 B.n190 B.n117 585
R241 B.n189 B.n188 585
R242 B.n187 B.n118 585
R243 B.n186 B.n185 585
R244 B.n184 B.n119 585
R245 B.n183 B.n182 585
R246 B.n181 B.n120 585
R247 B.n180 B.n179 585
R248 B.n178 B.n121 585
R249 B.n177 B.n176 585
R250 B.n175 B.n122 585
R251 B.n174 B.n173 585
R252 B.n172 B.n123 585
R253 B.n171 B.n170 585
R254 B.n169 B.n124 585
R255 B.n168 B.n167 585
R256 B.n166 B.n125 585
R257 B.n165 B.n164 585
R258 B.n163 B.n126 585
R259 B.n162 B.n161 585
R260 B.n160 B.n127 585
R261 B.n159 B.n158 585
R262 B.n157 B.n128 585
R263 B.n156 B.n155 585
R264 B.n154 B.n129 585
R265 B.n153 B.n152 585
R266 B.n151 B.n130 585
R267 B.n150 B.n149 585
R268 B.n148 B.n131 585
R269 B.n147 B.n146 585
R270 B.n145 B.n132 585
R271 B.n144 B.n143 585
R272 B.n142 B.n133 585
R273 B.n141 B.n140 585
R274 B.n139 B.n134 585
R275 B.n138 B.n137 585
R276 B.n136 B.n135 585
R277 B.n2 B.n0 585
R278 B.n513 B.n1 585
R279 B.n512 B.n511 585
R280 B.n510 B.n3 585
R281 B.n509 B.n508 585
R282 B.n507 B.n4 585
R283 B.n506 B.n505 585
R284 B.n504 B.n5 585
R285 B.n503 B.n502 585
R286 B.n501 B.n6 585
R287 B.n500 B.n499 585
R288 B.n498 B.n7 585
R289 B.n497 B.n496 585
R290 B.n495 B.n8 585
R291 B.n494 B.n493 585
R292 B.n492 B.n9 585
R293 B.n491 B.n490 585
R294 B.n489 B.n10 585
R295 B.n488 B.n487 585
R296 B.n486 B.n11 585
R297 B.n485 B.n484 585
R298 B.n483 B.n12 585
R299 B.n482 B.n481 585
R300 B.n480 B.n13 585
R301 B.n479 B.n478 585
R302 B.n477 B.n14 585
R303 B.n476 B.n475 585
R304 B.n474 B.n15 585
R305 B.n473 B.n472 585
R306 B.n471 B.n16 585
R307 B.n470 B.n469 585
R308 B.n468 B.n17 585
R309 B.n467 B.n466 585
R310 B.n465 B.n18 585
R311 B.n464 B.n463 585
R312 B.n462 B.n19 585
R313 B.n461 B.n460 585
R314 B.n459 B.n20 585
R315 B.n458 B.n457 585
R316 B.n456 B.n21 585
R317 B.n455 B.n454 585
R318 B.n453 B.n22 585
R319 B.n452 B.n451 585
R320 B.n450 B.n23 585
R321 B.n515 B.n514 585
R322 B.n199 B.n198 540.549
R323 B.n448 B.n23 540.549
R324 B.n259 B.n258 540.549
R325 B.n390 B.n47 540.549
R326 B.n98 B.t9 228.35
R327 B.n106 B.t6 228.35
R328 B.n32 B.t3 228.35
R329 B.n38 B.t0 228.35
R330 B.n98 B.t11 220.495
R331 B.n38 B.t1 220.495
R332 B.n106 B.t8 220.494
R333 B.n32 B.t4 220.494
R334 B.n198 B.n115 163.367
R335 B.n194 B.n115 163.367
R336 B.n194 B.n193 163.367
R337 B.n193 B.n192 163.367
R338 B.n192 B.n117 163.367
R339 B.n188 B.n117 163.367
R340 B.n188 B.n187 163.367
R341 B.n187 B.n186 163.367
R342 B.n186 B.n119 163.367
R343 B.n182 B.n119 163.367
R344 B.n182 B.n181 163.367
R345 B.n181 B.n180 163.367
R346 B.n180 B.n121 163.367
R347 B.n176 B.n121 163.367
R348 B.n176 B.n175 163.367
R349 B.n175 B.n174 163.367
R350 B.n174 B.n123 163.367
R351 B.n170 B.n123 163.367
R352 B.n170 B.n169 163.367
R353 B.n169 B.n168 163.367
R354 B.n168 B.n125 163.367
R355 B.n164 B.n125 163.367
R356 B.n164 B.n163 163.367
R357 B.n163 B.n162 163.367
R358 B.n162 B.n127 163.367
R359 B.n158 B.n127 163.367
R360 B.n158 B.n157 163.367
R361 B.n157 B.n156 163.367
R362 B.n156 B.n129 163.367
R363 B.n152 B.n129 163.367
R364 B.n152 B.n151 163.367
R365 B.n151 B.n150 163.367
R366 B.n150 B.n131 163.367
R367 B.n146 B.n131 163.367
R368 B.n146 B.n145 163.367
R369 B.n145 B.n144 163.367
R370 B.n144 B.n133 163.367
R371 B.n140 B.n133 163.367
R372 B.n140 B.n139 163.367
R373 B.n139 B.n138 163.367
R374 B.n138 B.n135 163.367
R375 B.n135 B.n2 163.367
R376 B.n514 B.n2 163.367
R377 B.n514 B.n513 163.367
R378 B.n513 B.n512 163.367
R379 B.n512 B.n3 163.367
R380 B.n508 B.n3 163.367
R381 B.n508 B.n507 163.367
R382 B.n507 B.n506 163.367
R383 B.n506 B.n5 163.367
R384 B.n502 B.n5 163.367
R385 B.n502 B.n501 163.367
R386 B.n501 B.n500 163.367
R387 B.n500 B.n7 163.367
R388 B.n496 B.n7 163.367
R389 B.n496 B.n495 163.367
R390 B.n495 B.n494 163.367
R391 B.n494 B.n9 163.367
R392 B.n490 B.n9 163.367
R393 B.n490 B.n489 163.367
R394 B.n489 B.n488 163.367
R395 B.n488 B.n11 163.367
R396 B.n484 B.n11 163.367
R397 B.n484 B.n483 163.367
R398 B.n483 B.n482 163.367
R399 B.n482 B.n13 163.367
R400 B.n478 B.n13 163.367
R401 B.n478 B.n477 163.367
R402 B.n477 B.n476 163.367
R403 B.n476 B.n15 163.367
R404 B.n472 B.n15 163.367
R405 B.n472 B.n471 163.367
R406 B.n471 B.n470 163.367
R407 B.n470 B.n17 163.367
R408 B.n466 B.n17 163.367
R409 B.n466 B.n465 163.367
R410 B.n465 B.n464 163.367
R411 B.n464 B.n19 163.367
R412 B.n460 B.n19 163.367
R413 B.n460 B.n459 163.367
R414 B.n459 B.n458 163.367
R415 B.n458 B.n21 163.367
R416 B.n454 B.n21 163.367
R417 B.n454 B.n453 163.367
R418 B.n453 B.n452 163.367
R419 B.n452 B.n23 163.367
R420 B.n200 B.n199 163.367
R421 B.n200 B.n113 163.367
R422 B.n204 B.n113 163.367
R423 B.n205 B.n204 163.367
R424 B.n206 B.n205 163.367
R425 B.n206 B.n111 163.367
R426 B.n210 B.n111 163.367
R427 B.n211 B.n210 163.367
R428 B.n212 B.n211 163.367
R429 B.n212 B.n109 163.367
R430 B.n216 B.n109 163.367
R431 B.n217 B.n216 163.367
R432 B.n218 B.n217 163.367
R433 B.n218 B.n105 163.367
R434 B.n223 B.n105 163.367
R435 B.n224 B.n223 163.367
R436 B.n225 B.n224 163.367
R437 B.n225 B.n103 163.367
R438 B.n229 B.n103 163.367
R439 B.n230 B.n229 163.367
R440 B.n231 B.n230 163.367
R441 B.n231 B.n101 163.367
R442 B.n235 B.n101 163.367
R443 B.n236 B.n235 163.367
R444 B.n236 B.n97 163.367
R445 B.n240 B.n97 163.367
R446 B.n241 B.n240 163.367
R447 B.n242 B.n241 163.367
R448 B.n242 B.n95 163.367
R449 B.n246 B.n95 163.367
R450 B.n247 B.n246 163.367
R451 B.n248 B.n247 163.367
R452 B.n248 B.n93 163.367
R453 B.n252 B.n93 163.367
R454 B.n253 B.n252 163.367
R455 B.n254 B.n253 163.367
R456 B.n254 B.n91 163.367
R457 B.n258 B.n91 163.367
R458 B.n260 B.n259 163.367
R459 B.n260 B.n89 163.367
R460 B.n264 B.n89 163.367
R461 B.n265 B.n264 163.367
R462 B.n266 B.n265 163.367
R463 B.n266 B.n87 163.367
R464 B.n270 B.n87 163.367
R465 B.n271 B.n270 163.367
R466 B.n272 B.n271 163.367
R467 B.n272 B.n85 163.367
R468 B.n276 B.n85 163.367
R469 B.n277 B.n276 163.367
R470 B.n278 B.n277 163.367
R471 B.n278 B.n83 163.367
R472 B.n282 B.n83 163.367
R473 B.n283 B.n282 163.367
R474 B.n284 B.n283 163.367
R475 B.n284 B.n81 163.367
R476 B.n288 B.n81 163.367
R477 B.n289 B.n288 163.367
R478 B.n290 B.n289 163.367
R479 B.n290 B.n79 163.367
R480 B.n294 B.n79 163.367
R481 B.n295 B.n294 163.367
R482 B.n296 B.n295 163.367
R483 B.n296 B.n77 163.367
R484 B.n300 B.n77 163.367
R485 B.n301 B.n300 163.367
R486 B.n302 B.n301 163.367
R487 B.n302 B.n75 163.367
R488 B.n306 B.n75 163.367
R489 B.n307 B.n306 163.367
R490 B.n308 B.n307 163.367
R491 B.n308 B.n73 163.367
R492 B.n312 B.n73 163.367
R493 B.n313 B.n312 163.367
R494 B.n314 B.n313 163.367
R495 B.n314 B.n71 163.367
R496 B.n318 B.n71 163.367
R497 B.n319 B.n318 163.367
R498 B.n320 B.n319 163.367
R499 B.n320 B.n69 163.367
R500 B.n324 B.n69 163.367
R501 B.n325 B.n324 163.367
R502 B.n326 B.n325 163.367
R503 B.n326 B.n67 163.367
R504 B.n330 B.n67 163.367
R505 B.n331 B.n330 163.367
R506 B.n332 B.n331 163.367
R507 B.n332 B.n65 163.367
R508 B.n336 B.n65 163.367
R509 B.n337 B.n336 163.367
R510 B.n338 B.n337 163.367
R511 B.n338 B.n63 163.367
R512 B.n342 B.n63 163.367
R513 B.n343 B.n342 163.367
R514 B.n344 B.n343 163.367
R515 B.n344 B.n61 163.367
R516 B.n348 B.n61 163.367
R517 B.n349 B.n348 163.367
R518 B.n350 B.n349 163.367
R519 B.n350 B.n59 163.367
R520 B.n354 B.n59 163.367
R521 B.n355 B.n354 163.367
R522 B.n356 B.n355 163.367
R523 B.n356 B.n57 163.367
R524 B.n360 B.n57 163.367
R525 B.n361 B.n360 163.367
R526 B.n362 B.n361 163.367
R527 B.n362 B.n55 163.367
R528 B.n366 B.n55 163.367
R529 B.n367 B.n366 163.367
R530 B.n368 B.n367 163.367
R531 B.n368 B.n53 163.367
R532 B.n372 B.n53 163.367
R533 B.n373 B.n372 163.367
R534 B.n374 B.n373 163.367
R535 B.n374 B.n51 163.367
R536 B.n378 B.n51 163.367
R537 B.n379 B.n378 163.367
R538 B.n380 B.n379 163.367
R539 B.n380 B.n49 163.367
R540 B.n384 B.n49 163.367
R541 B.n385 B.n384 163.367
R542 B.n386 B.n385 163.367
R543 B.n386 B.n47 163.367
R544 B.n448 B.n447 163.367
R545 B.n447 B.n446 163.367
R546 B.n446 B.n25 163.367
R547 B.n442 B.n25 163.367
R548 B.n442 B.n441 163.367
R549 B.n441 B.n440 163.367
R550 B.n440 B.n27 163.367
R551 B.n436 B.n27 163.367
R552 B.n436 B.n435 163.367
R553 B.n435 B.n434 163.367
R554 B.n434 B.n29 163.367
R555 B.n430 B.n29 163.367
R556 B.n430 B.n429 163.367
R557 B.n429 B.n428 163.367
R558 B.n428 B.n31 163.367
R559 B.n423 B.n31 163.367
R560 B.n423 B.n422 163.367
R561 B.n422 B.n421 163.367
R562 B.n421 B.n35 163.367
R563 B.n417 B.n35 163.367
R564 B.n417 B.n416 163.367
R565 B.n416 B.n415 163.367
R566 B.n415 B.n37 163.367
R567 B.n410 B.n37 163.367
R568 B.n410 B.n409 163.367
R569 B.n409 B.n408 163.367
R570 B.n408 B.n41 163.367
R571 B.n404 B.n41 163.367
R572 B.n404 B.n403 163.367
R573 B.n403 B.n402 163.367
R574 B.n402 B.n43 163.367
R575 B.n398 B.n43 163.367
R576 B.n398 B.n397 163.367
R577 B.n397 B.n396 163.367
R578 B.n396 B.n45 163.367
R579 B.n392 B.n45 163.367
R580 B.n392 B.n391 163.367
R581 B.n391 B.n390 163.367
R582 B.n99 B.t10 143.501
R583 B.n39 B.t2 143.501
R584 B.n107 B.t7 143.5
R585 B.n33 B.t5 143.5
R586 B.n99 B.n98 76.9944
R587 B.n107 B.n106 76.9944
R588 B.n33 B.n32 76.9944
R589 B.n39 B.n38 76.9944
R590 B.n100 B.n99 59.5399
R591 B.n221 B.n107 59.5399
R592 B.n426 B.n33 59.5399
R593 B.n412 B.n39 59.5399
R594 B.n450 B.n449 35.1225
R595 B.n389 B.n388 35.1225
R596 B.n257 B.n90 35.1225
R597 B.n197 B.n114 35.1225
R598 B B.n515 18.0485
R599 B.n449 B.n24 10.6151
R600 B.n445 B.n24 10.6151
R601 B.n445 B.n444 10.6151
R602 B.n444 B.n443 10.6151
R603 B.n443 B.n26 10.6151
R604 B.n439 B.n26 10.6151
R605 B.n439 B.n438 10.6151
R606 B.n438 B.n437 10.6151
R607 B.n437 B.n28 10.6151
R608 B.n433 B.n28 10.6151
R609 B.n433 B.n432 10.6151
R610 B.n432 B.n431 10.6151
R611 B.n431 B.n30 10.6151
R612 B.n427 B.n30 10.6151
R613 B.n425 B.n424 10.6151
R614 B.n424 B.n34 10.6151
R615 B.n420 B.n34 10.6151
R616 B.n420 B.n419 10.6151
R617 B.n419 B.n418 10.6151
R618 B.n418 B.n36 10.6151
R619 B.n414 B.n36 10.6151
R620 B.n414 B.n413 10.6151
R621 B.n411 B.n40 10.6151
R622 B.n407 B.n40 10.6151
R623 B.n407 B.n406 10.6151
R624 B.n406 B.n405 10.6151
R625 B.n405 B.n42 10.6151
R626 B.n401 B.n42 10.6151
R627 B.n401 B.n400 10.6151
R628 B.n400 B.n399 10.6151
R629 B.n399 B.n44 10.6151
R630 B.n395 B.n44 10.6151
R631 B.n395 B.n394 10.6151
R632 B.n394 B.n393 10.6151
R633 B.n393 B.n46 10.6151
R634 B.n389 B.n46 10.6151
R635 B.n261 B.n90 10.6151
R636 B.n262 B.n261 10.6151
R637 B.n263 B.n262 10.6151
R638 B.n263 B.n88 10.6151
R639 B.n267 B.n88 10.6151
R640 B.n268 B.n267 10.6151
R641 B.n269 B.n268 10.6151
R642 B.n269 B.n86 10.6151
R643 B.n273 B.n86 10.6151
R644 B.n274 B.n273 10.6151
R645 B.n275 B.n274 10.6151
R646 B.n275 B.n84 10.6151
R647 B.n279 B.n84 10.6151
R648 B.n280 B.n279 10.6151
R649 B.n281 B.n280 10.6151
R650 B.n281 B.n82 10.6151
R651 B.n285 B.n82 10.6151
R652 B.n286 B.n285 10.6151
R653 B.n287 B.n286 10.6151
R654 B.n287 B.n80 10.6151
R655 B.n291 B.n80 10.6151
R656 B.n292 B.n291 10.6151
R657 B.n293 B.n292 10.6151
R658 B.n293 B.n78 10.6151
R659 B.n297 B.n78 10.6151
R660 B.n298 B.n297 10.6151
R661 B.n299 B.n298 10.6151
R662 B.n299 B.n76 10.6151
R663 B.n303 B.n76 10.6151
R664 B.n304 B.n303 10.6151
R665 B.n305 B.n304 10.6151
R666 B.n305 B.n74 10.6151
R667 B.n309 B.n74 10.6151
R668 B.n310 B.n309 10.6151
R669 B.n311 B.n310 10.6151
R670 B.n311 B.n72 10.6151
R671 B.n315 B.n72 10.6151
R672 B.n316 B.n315 10.6151
R673 B.n317 B.n316 10.6151
R674 B.n317 B.n70 10.6151
R675 B.n321 B.n70 10.6151
R676 B.n322 B.n321 10.6151
R677 B.n323 B.n322 10.6151
R678 B.n323 B.n68 10.6151
R679 B.n327 B.n68 10.6151
R680 B.n328 B.n327 10.6151
R681 B.n329 B.n328 10.6151
R682 B.n329 B.n66 10.6151
R683 B.n333 B.n66 10.6151
R684 B.n334 B.n333 10.6151
R685 B.n335 B.n334 10.6151
R686 B.n335 B.n64 10.6151
R687 B.n339 B.n64 10.6151
R688 B.n340 B.n339 10.6151
R689 B.n341 B.n340 10.6151
R690 B.n341 B.n62 10.6151
R691 B.n345 B.n62 10.6151
R692 B.n346 B.n345 10.6151
R693 B.n347 B.n346 10.6151
R694 B.n347 B.n60 10.6151
R695 B.n351 B.n60 10.6151
R696 B.n352 B.n351 10.6151
R697 B.n353 B.n352 10.6151
R698 B.n353 B.n58 10.6151
R699 B.n357 B.n58 10.6151
R700 B.n358 B.n357 10.6151
R701 B.n359 B.n358 10.6151
R702 B.n359 B.n56 10.6151
R703 B.n363 B.n56 10.6151
R704 B.n364 B.n363 10.6151
R705 B.n365 B.n364 10.6151
R706 B.n365 B.n54 10.6151
R707 B.n369 B.n54 10.6151
R708 B.n370 B.n369 10.6151
R709 B.n371 B.n370 10.6151
R710 B.n371 B.n52 10.6151
R711 B.n375 B.n52 10.6151
R712 B.n376 B.n375 10.6151
R713 B.n377 B.n376 10.6151
R714 B.n377 B.n50 10.6151
R715 B.n381 B.n50 10.6151
R716 B.n382 B.n381 10.6151
R717 B.n383 B.n382 10.6151
R718 B.n383 B.n48 10.6151
R719 B.n387 B.n48 10.6151
R720 B.n388 B.n387 10.6151
R721 B.n201 B.n114 10.6151
R722 B.n202 B.n201 10.6151
R723 B.n203 B.n202 10.6151
R724 B.n203 B.n112 10.6151
R725 B.n207 B.n112 10.6151
R726 B.n208 B.n207 10.6151
R727 B.n209 B.n208 10.6151
R728 B.n209 B.n110 10.6151
R729 B.n213 B.n110 10.6151
R730 B.n214 B.n213 10.6151
R731 B.n215 B.n214 10.6151
R732 B.n215 B.n108 10.6151
R733 B.n219 B.n108 10.6151
R734 B.n220 B.n219 10.6151
R735 B.n222 B.n104 10.6151
R736 B.n226 B.n104 10.6151
R737 B.n227 B.n226 10.6151
R738 B.n228 B.n227 10.6151
R739 B.n228 B.n102 10.6151
R740 B.n232 B.n102 10.6151
R741 B.n233 B.n232 10.6151
R742 B.n234 B.n233 10.6151
R743 B.n238 B.n237 10.6151
R744 B.n239 B.n238 10.6151
R745 B.n239 B.n96 10.6151
R746 B.n243 B.n96 10.6151
R747 B.n244 B.n243 10.6151
R748 B.n245 B.n244 10.6151
R749 B.n245 B.n94 10.6151
R750 B.n249 B.n94 10.6151
R751 B.n250 B.n249 10.6151
R752 B.n251 B.n250 10.6151
R753 B.n251 B.n92 10.6151
R754 B.n255 B.n92 10.6151
R755 B.n256 B.n255 10.6151
R756 B.n257 B.n256 10.6151
R757 B.n197 B.n196 10.6151
R758 B.n196 B.n195 10.6151
R759 B.n195 B.n116 10.6151
R760 B.n191 B.n116 10.6151
R761 B.n191 B.n190 10.6151
R762 B.n190 B.n189 10.6151
R763 B.n189 B.n118 10.6151
R764 B.n185 B.n118 10.6151
R765 B.n185 B.n184 10.6151
R766 B.n184 B.n183 10.6151
R767 B.n183 B.n120 10.6151
R768 B.n179 B.n120 10.6151
R769 B.n179 B.n178 10.6151
R770 B.n178 B.n177 10.6151
R771 B.n177 B.n122 10.6151
R772 B.n173 B.n122 10.6151
R773 B.n173 B.n172 10.6151
R774 B.n172 B.n171 10.6151
R775 B.n171 B.n124 10.6151
R776 B.n167 B.n124 10.6151
R777 B.n167 B.n166 10.6151
R778 B.n166 B.n165 10.6151
R779 B.n165 B.n126 10.6151
R780 B.n161 B.n126 10.6151
R781 B.n161 B.n160 10.6151
R782 B.n160 B.n159 10.6151
R783 B.n159 B.n128 10.6151
R784 B.n155 B.n128 10.6151
R785 B.n155 B.n154 10.6151
R786 B.n154 B.n153 10.6151
R787 B.n153 B.n130 10.6151
R788 B.n149 B.n130 10.6151
R789 B.n149 B.n148 10.6151
R790 B.n148 B.n147 10.6151
R791 B.n147 B.n132 10.6151
R792 B.n143 B.n132 10.6151
R793 B.n143 B.n142 10.6151
R794 B.n142 B.n141 10.6151
R795 B.n141 B.n134 10.6151
R796 B.n137 B.n134 10.6151
R797 B.n137 B.n136 10.6151
R798 B.n136 B.n0 10.6151
R799 B.n511 B.n1 10.6151
R800 B.n511 B.n510 10.6151
R801 B.n510 B.n509 10.6151
R802 B.n509 B.n4 10.6151
R803 B.n505 B.n4 10.6151
R804 B.n505 B.n504 10.6151
R805 B.n504 B.n503 10.6151
R806 B.n503 B.n6 10.6151
R807 B.n499 B.n6 10.6151
R808 B.n499 B.n498 10.6151
R809 B.n498 B.n497 10.6151
R810 B.n497 B.n8 10.6151
R811 B.n493 B.n8 10.6151
R812 B.n493 B.n492 10.6151
R813 B.n492 B.n491 10.6151
R814 B.n491 B.n10 10.6151
R815 B.n487 B.n10 10.6151
R816 B.n487 B.n486 10.6151
R817 B.n486 B.n485 10.6151
R818 B.n485 B.n12 10.6151
R819 B.n481 B.n12 10.6151
R820 B.n481 B.n480 10.6151
R821 B.n480 B.n479 10.6151
R822 B.n479 B.n14 10.6151
R823 B.n475 B.n14 10.6151
R824 B.n475 B.n474 10.6151
R825 B.n474 B.n473 10.6151
R826 B.n473 B.n16 10.6151
R827 B.n469 B.n16 10.6151
R828 B.n469 B.n468 10.6151
R829 B.n468 B.n467 10.6151
R830 B.n467 B.n18 10.6151
R831 B.n463 B.n18 10.6151
R832 B.n463 B.n462 10.6151
R833 B.n462 B.n461 10.6151
R834 B.n461 B.n20 10.6151
R835 B.n457 B.n20 10.6151
R836 B.n457 B.n456 10.6151
R837 B.n456 B.n455 10.6151
R838 B.n455 B.n22 10.6151
R839 B.n451 B.n22 10.6151
R840 B.n451 B.n450 10.6151
R841 B.n426 B.n425 6.5566
R842 B.n413 B.n412 6.5566
R843 B.n222 B.n221 6.5566
R844 B.n234 B.n100 6.5566
R845 B.n427 B.n426 4.05904
R846 B.n412 B.n411 4.05904
R847 B.n221 B.n220 4.05904
R848 B.n237 B.n100 4.05904
R849 B.n515 B.n0 2.81026
R850 B.n515 B.n1 2.81026
C0 B VDD1 1.20009f
C1 VN VDD1 0.155073f
C2 B VN 1.188f
C3 VDD1 VDD2 1.27811f
C4 VP w_n3352_n1546# 6.11895f
C5 VTAIL VDD1 3.76699f
C6 B VDD2 1.26975f
C7 VN VDD2 1.45704f
C8 VTAIL B 2.14471f
C9 VTAIL VN 2.17726f
C10 VTAIL VDD2 3.82817f
C11 VDD1 w_n3352_n1546# 1.40277f
C12 VP VDD1 1.76644f
C13 B w_n3352_n1546# 8.01265f
C14 VN w_n3352_n1546# 5.68792f
C15 VP B 1.91183f
C16 VP VN 5.25734f
C17 VDD2 w_n3352_n1546# 1.48128f
C18 VP VDD2 0.466335f
C19 VTAIL w_n3352_n1546# 1.99151f
C20 VP VTAIL 2.19136f
C21 VDD2 VSUBS 0.823983f
C22 VDD1 VSUBS 3.96801f
C23 VTAIL VSUBS 0.658043f
C24 VN VSUBS 6.0518f
C25 VP VSUBS 2.304541f
C26 B VSUBS 4.153059f
C27 w_n3352_n1546# VSUBS 65.6858f
C28 B.n0 VSUBS 0.006312f
C29 B.n1 VSUBS 0.006312f
C30 B.n2 VSUBS 0.009981f
C31 B.n3 VSUBS 0.009981f
C32 B.n4 VSUBS 0.009981f
C33 B.n5 VSUBS 0.009981f
C34 B.n6 VSUBS 0.009981f
C35 B.n7 VSUBS 0.009981f
C36 B.n8 VSUBS 0.009981f
C37 B.n9 VSUBS 0.009981f
C38 B.n10 VSUBS 0.009981f
C39 B.n11 VSUBS 0.009981f
C40 B.n12 VSUBS 0.009981f
C41 B.n13 VSUBS 0.009981f
C42 B.n14 VSUBS 0.009981f
C43 B.n15 VSUBS 0.009981f
C44 B.n16 VSUBS 0.009981f
C45 B.n17 VSUBS 0.009981f
C46 B.n18 VSUBS 0.009981f
C47 B.n19 VSUBS 0.009981f
C48 B.n20 VSUBS 0.009981f
C49 B.n21 VSUBS 0.009981f
C50 B.n22 VSUBS 0.009981f
C51 B.n23 VSUBS 0.023964f
C52 B.n24 VSUBS 0.009981f
C53 B.n25 VSUBS 0.009981f
C54 B.n26 VSUBS 0.009981f
C55 B.n27 VSUBS 0.009981f
C56 B.n28 VSUBS 0.009981f
C57 B.n29 VSUBS 0.009981f
C58 B.n30 VSUBS 0.009981f
C59 B.n31 VSUBS 0.009981f
C60 B.t5 VSUBS 0.098117f
C61 B.t4 VSUBS 0.127493f
C62 B.t3 VSUBS 0.736001f
C63 B.n32 VSUBS 0.126663f
C64 B.n33 VSUBS 0.098363f
C65 B.n34 VSUBS 0.009981f
C66 B.n35 VSUBS 0.009981f
C67 B.n36 VSUBS 0.009981f
C68 B.n37 VSUBS 0.009981f
C69 B.t2 VSUBS 0.098117f
C70 B.t1 VSUBS 0.127493f
C71 B.t0 VSUBS 0.736001f
C72 B.n38 VSUBS 0.126663f
C73 B.n39 VSUBS 0.098363f
C74 B.n40 VSUBS 0.009981f
C75 B.n41 VSUBS 0.009981f
C76 B.n42 VSUBS 0.009981f
C77 B.n43 VSUBS 0.009981f
C78 B.n44 VSUBS 0.009981f
C79 B.n45 VSUBS 0.009981f
C80 B.n46 VSUBS 0.009981f
C81 B.n47 VSUBS 0.023964f
C82 B.n48 VSUBS 0.009981f
C83 B.n49 VSUBS 0.009981f
C84 B.n50 VSUBS 0.009981f
C85 B.n51 VSUBS 0.009981f
C86 B.n52 VSUBS 0.009981f
C87 B.n53 VSUBS 0.009981f
C88 B.n54 VSUBS 0.009981f
C89 B.n55 VSUBS 0.009981f
C90 B.n56 VSUBS 0.009981f
C91 B.n57 VSUBS 0.009981f
C92 B.n58 VSUBS 0.009981f
C93 B.n59 VSUBS 0.009981f
C94 B.n60 VSUBS 0.009981f
C95 B.n61 VSUBS 0.009981f
C96 B.n62 VSUBS 0.009981f
C97 B.n63 VSUBS 0.009981f
C98 B.n64 VSUBS 0.009981f
C99 B.n65 VSUBS 0.009981f
C100 B.n66 VSUBS 0.009981f
C101 B.n67 VSUBS 0.009981f
C102 B.n68 VSUBS 0.009981f
C103 B.n69 VSUBS 0.009981f
C104 B.n70 VSUBS 0.009981f
C105 B.n71 VSUBS 0.009981f
C106 B.n72 VSUBS 0.009981f
C107 B.n73 VSUBS 0.009981f
C108 B.n74 VSUBS 0.009981f
C109 B.n75 VSUBS 0.009981f
C110 B.n76 VSUBS 0.009981f
C111 B.n77 VSUBS 0.009981f
C112 B.n78 VSUBS 0.009981f
C113 B.n79 VSUBS 0.009981f
C114 B.n80 VSUBS 0.009981f
C115 B.n81 VSUBS 0.009981f
C116 B.n82 VSUBS 0.009981f
C117 B.n83 VSUBS 0.009981f
C118 B.n84 VSUBS 0.009981f
C119 B.n85 VSUBS 0.009981f
C120 B.n86 VSUBS 0.009981f
C121 B.n87 VSUBS 0.009981f
C122 B.n88 VSUBS 0.009981f
C123 B.n89 VSUBS 0.009981f
C124 B.n90 VSUBS 0.023964f
C125 B.n91 VSUBS 0.009981f
C126 B.n92 VSUBS 0.009981f
C127 B.n93 VSUBS 0.009981f
C128 B.n94 VSUBS 0.009981f
C129 B.n95 VSUBS 0.009981f
C130 B.n96 VSUBS 0.009981f
C131 B.n97 VSUBS 0.009981f
C132 B.t10 VSUBS 0.098117f
C133 B.t11 VSUBS 0.127493f
C134 B.t9 VSUBS 0.736001f
C135 B.n98 VSUBS 0.126663f
C136 B.n99 VSUBS 0.098363f
C137 B.n100 VSUBS 0.023125f
C138 B.n101 VSUBS 0.009981f
C139 B.n102 VSUBS 0.009981f
C140 B.n103 VSUBS 0.009981f
C141 B.n104 VSUBS 0.009981f
C142 B.n105 VSUBS 0.009981f
C143 B.t7 VSUBS 0.098117f
C144 B.t8 VSUBS 0.127493f
C145 B.t6 VSUBS 0.736001f
C146 B.n106 VSUBS 0.126663f
C147 B.n107 VSUBS 0.098363f
C148 B.n108 VSUBS 0.009981f
C149 B.n109 VSUBS 0.009981f
C150 B.n110 VSUBS 0.009981f
C151 B.n111 VSUBS 0.009981f
C152 B.n112 VSUBS 0.009981f
C153 B.n113 VSUBS 0.009981f
C154 B.n114 VSUBS 0.025061f
C155 B.n115 VSUBS 0.009981f
C156 B.n116 VSUBS 0.009981f
C157 B.n117 VSUBS 0.009981f
C158 B.n118 VSUBS 0.009981f
C159 B.n119 VSUBS 0.009981f
C160 B.n120 VSUBS 0.009981f
C161 B.n121 VSUBS 0.009981f
C162 B.n122 VSUBS 0.009981f
C163 B.n123 VSUBS 0.009981f
C164 B.n124 VSUBS 0.009981f
C165 B.n125 VSUBS 0.009981f
C166 B.n126 VSUBS 0.009981f
C167 B.n127 VSUBS 0.009981f
C168 B.n128 VSUBS 0.009981f
C169 B.n129 VSUBS 0.009981f
C170 B.n130 VSUBS 0.009981f
C171 B.n131 VSUBS 0.009981f
C172 B.n132 VSUBS 0.009981f
C173 B.n133 VSUBS 0.009981f
C174 B.n134 VSUBS 0.009981f
C175 B.n135 VSUBS 0.009981f
C176 B.n136 VSUBS 0.009981f
C177 B.n137 VSUBS 0.009981f
C178 B.n138 VSUBS 0.009981f
C179 B.n139 VSUBS 0.009981f
C180 B.n140 VSUBS 0.009981f
C181 B.n141 VSUBS 0.009981f
C182 B.n142 VSUBS 0.009981f
C183 B.n143 VSUBS 0.009981f
C184 B.n144 VSUBS 0.009981f
C185 B.n145 VSUBS 0.009981f
C186 B.n146 VSUBS 0.009981f
C187 B.n147 VSUBS 0.009981f
C188 B.n148 VSUBS 0.009981f
C189 B.n149 VSUBS 0.009981f
C190 B.n150 VSUBS 0.009981f
C191 B.n151 VSUBS 0.009981f
C192 B.n152 VSUBS 0.009981f
C193 B.n153 VSUBS 0.009981f
C194 B.n154 VSUBS 0.009981f
C195 B.n155 VSUBS 0.009981f
C196 B.n156 VSUBS 0.009981f
C197 B.n157 VSUBS 0.009981f
C198 B.n158 VSUBS 0.009981f
C199 B.n159 VSUBS 0.009981f
C200 B.n160 VSUBS 0.009981f
C201 B.n161 VSUBS 0.009981f
C202 B.n162 VSUBS 0.009981f
C203 B.n163 VSUBS 0.009981f
C204 B.n164 VSUBS 0.009981f
C205 B.n165 VSUBS 0.009981f
C206 B.n166 VSUBS 0.009981f
C207 B.n167 VSUBS 0.009981f
C208 B.n168 VSUBS 0.009981f
C209 B.n169 VSUBS 0.009981f
C210 B.n170 VSUBS 0.009981f
C211 B.n171 VSUBS 0.009981f
C212 B.n172 VSUBS 0.009981f
C213 B.n173 VSUBS 0.009981f
C214 B.n174 VSUBS 0.009981f
C215 B.n175 VSUBS 0.009981f
C216 B.n176 VSUBS 0.009981f
C217 B.n177 VSUBS 0.009981f
C218 B.n178 VSUBS 0.009981f
C219 B.n179 VSUBS 0.009981f
C220 B.n180 VSUBS 0.009981f
C221 B.n181 VSUBS 0.009981f
C222 B.n182 VSUBS 0.009981f
C223 B.n183 VSUBS 0.009981f
C224 B.n184 VSUBS 0.009981f
C225 B.n185 VSUBS 0.009981f
C226 B.n186 VSUBS 0.009981f
C227 B.n187 VSUBS 0.009981f
C228 B.n188 VSUBS 0.009981f
C229 B.n189 VSUBS 0.009981f
C230 B.n190 VSUBS 0.009981f
C231 B.n191 VSUBS 0.009981f
C232 B.n192 VSUBS 0.009981f
C233 B.n193 VSUBS 0.009981f
C234 B.n194 VSUBS 0.009981f
C235 B.n195 VSUBS 0.009981f
C236 B.n196 VSUBS 0.009981f
C237 B.n197 VSUBS 0.023964f
C238 B.n198 VSUBS 0.023964f
C239 B.n199 VSUBS 0.025061f
C240 B.n200 VSUBS 0.009981f
C241 B.n201 VSUBS 0.009981f
C242 B.n202 VSUBS 0.009981f
C243 B.n203 VSUBS 0.009981f
C244 B.n204 VSUBS 0.009981f
C245 B.n205 VSUBS 0.009981f
C246 B.n206 VSUBS 0.009981f
C247 B.n207 VSUBS 0.009981f
C248 B.n208 VSUBS 0.009981f
C249 B.n209 VSUBS 0.009981f
C250 B.n210 VSUBS 0.009981f
C251 B.n211 VSUBS 0.009981f
C252 B.n212 VSUBS 0.009981f
C253 B.n213 VSUBS 0.009981f
C254 B.n214 VSUBS 0.009981f
C255 B.n215 VSUBS 0.009981f
C256 B.n216 VSUBS 0.009981f
C257 B.n217 VSUBS 0.009981f
C258 B.n218 VSUBS 0.009981f
C259 B.n219 VSUBS 0.009981f
C260 B.n220 VSUBS 0.006899f
C261 B.n221 VSUBS 0.023125f
C262 B.n222 VSUBS 0.008073f
C263 B.n223 VSUBS 0.009981f
C264 B.n224 VSUBS 0.009981f
C265 B.n225 VSUBS 0.009981f
C266 B.n226 VSUBS 0.009981f
C267 B.n227 VSUBS 0.009981f
C268 B.n228 VSUBS 0.009981f
C269 B.n229 VSUBS 0.009981f
C270 B.n230 VSUBS 0.009981f
C271 B.n231 VSUBS 0.009981f
C272 B.n232 VSUBS 0.009981f
C273 B.n233 VSUBS 0.009981f
C274 B.n234 VSUBS 0.008073f
C275 B.n235 VSUBS 0.009981f
C276 B.n236 VSUBS 0.009981f
C277 B.n237 VSUBS 0.006899f
C278 B.n238 VSUBS 0.009981f
C279 B.n239 VSUBS 0.009981f
C280 B.n240 VSUBS 0.009981f
C281 B.n241 VSUBS 0.009981f
C282 B.n242 VSUBS 0.009981f
C283 B.n243 VSUBS 0.009981f
C284 B.n244 VSUBS 0.009981f
C285 B.n245 VSUBS 0.009981f
C286 B.n246 VSUBS 0.009981f
C287 B.n247 VSUBS 0.009981f
C288 B.n248 VSUBS 0.009981f
C289 B.n249 VSUBS 0.009981f
C290 B.n250 VSUBS 0.009981f
C291 B.n251 VSUBS 0.009981f
C292 B.n252 VSUBS 0.009981f
C293 B.n253 VSUBS 0.009981f
C294 B.n254 VSUBS 0.009981f
C295 B.n255 VSUBS 0.009981f
C296 B.n256 VSUBS 0.009981f
C297 B.n257 VSUBS 0.025061f
C298 B.n258 VSUBS 0.025061f
C299 B.n259 VSUBS 0.023964f
C300 B.n260 VSUBS 0.009981f
C301 B.n261 VSUBS 0.009981f
C302 B.n262 VSUBS 0.009981f
C303 B.n263 VSUBS 0.009981f
C304 B.n264 VSUBS 0.009981f
C305 B.n265 VSUBS 0.009981f
C306 B.n266 VSUBS 0.009981f
C307 B.n267 VSUBS 0.009981f
C308 B.n268 VSUBS 0.009981f
C309 B.n269 VSUBS 0.009981f
C310 B.n270 VSUBS 0.009981f
C311 B.n271 VSUBS 0.009981f
C312 B.n272 VSUBS 0.009981f
C313 B.n273 VSUBS 0.009981f
C314 B.n274 VSUBS 0.009981f
C315 B.n275 VSUBS 0.009981f
C316 B.n276 VSUBS 0.009981f
C317 B.n277 VSUBS 0.009981f
C318 B.n278 VSUBS 0.009981f
C319 B.n279 VSUBS 0.009981f
C320 B.n280 VSUBS 0.009981f
C321 B.n281 VSUBS 0.009981f
C322 B.n282 VSUBS 0.009981f
C323 B.n283 VSUBS 0.009981f
C324 B.n284 VSUBS 0.009981f
C325 B.n285 VSUBS 0.009981f
C326 B.n286 VSUBS 0.009981f
C327 B.n287 VSUBS 0.009981f
C328 B.n288 VSUBS 0.009981f
C329 B.n289 VSUBS 0.009981f
C330 B.n290 VSUBS 0.009981f
C331 B.n291 VSUBS 0.009981f
C332 B.n292 VSUBS 0.009981f
C333 B.n293 VSUBS 0.009981f
C334 B.n294 VSUBS 0.009981f
C335 B.n295 VSUBS 0.009981f
C336 B.n296 VSUBS 0.009981f
C337 B.n297 VSUBS 0.009981f
C338 B.n298 VSUBS 0.009981f
C339 B.n299 VSUBS 0.009981f
C340 B.n300 VSUBS 0.009981f
C341 B.n301 VSUBS 0.009981f
C342 B.n302 VSUBS 0.009981f
C343 B.n303 VSUBS 0.009981f
C344 B.n304 VSUBS 0.009981f
C345 B.n305 VSUBS 0.009981f
C346 B.n306 VSUBS 0.009981f
C347 B.n307 VSUBS 0.009981f
C348 B.n308 VSUBS 0.009981f
C349 B.n309 VSUBS 0.009981f
C350 B.n310 VSUBS 0.009981f
C351 B.n311 VSUBS 0.009981f
C352 B.n312 VSUBS 0.009981f
C353 B.n313 VSUBS 0.009981f
C354 B.n314 VSUBS 0.009981f
C355 B.n315 VSUBS 0.009981f
C356 B.n316 VSUBS 0.009981f
C357 B.n317 VSUBS 0.009981f
C358 B.n318 VSUBS 0.009981f
C359 B.n319 VSUBS 0.009981f
C360 B.n320 VSUBS 0.009981f
C361 B.n321 VSUBS 0.009981f
C362 B.n322 VSUBS 0.009981f
C363 B.n323 VSUBS 0.009981f
C364 B.n324 VSUBS 0.009981f
C365 B.n325 VSUBS 0.009981f
C366 B.n326 VSUBS 0.009981f
C367 B.n327 VSUBS 0.009981f
C368 B.n328 VSUBS 0.009981f
C369 B.n329 VSUBS 0.009981f
C370 B.n330 VSUBS 0.009981f
C371 B.n331 VSUBS 0.009981f
C372 B.n332 VSUBS 0.009981f
C373 B.n333 VSUBS 0.009981f
C374 B.n334 VSUBS 0.009981f
C375 B.n335 VSUBS 0.009981f
C376 B.n336 VSUBS 0.009981f
C377 B.n337 VSUBS 0.009981f
C378 B.n338 VSUBS 0.009981f
C379 B.n339 VSUBS 0.009981f
C380 B.n340 VSUBS 0.009981f
C381 B.n341 VSUBS 0.009981f
C382 B.n342 VSUBS 0.009981f
C383 B.n343 VSUBS 0.009981f
C384 B.n344 VSUBS 0.009981f
C385 B.n345 VSUBS 0.009981f
C386 B.n346 VSUBS 0.009981f
C387 B.n347 VSUBS 0.009981f
C388 B.n348 VSUBS 0.009981f
C389 B.n349 VSUBS 0.009981f
C390 B.n350 VSUBS 0.009981f
C391 B.n351 VSUBS 0.009981f
C392 B.n352 VSUBS 0.009981f
C393 B.n353 VSUBS 0.009981f
C394 B.n354 VSUBS 0.009981f
C395 B.n355 VSUBS 0.009981f
C396 B.n356 VSUBS 0.009981f
C397 B.n357 VSUBS 0.009981f
C398 B.n358 VSUBS 0.009981f
C399 B.n359 VSUBS 0.009981f
C400 B.n360 VSUBS 0.009981f
C401 B.n361 VSUBS 0.009981f
C402 B.n362 VSUBS 0.009981f
C403 B.n363 VSUBS 0.009981f
C404 B.n364 VSUBS 0.009981f
C405 B.n365 VSUBS 0.009981f
C406 B.n366 VSUBS 0.009981f
C407 B.n367 VSUBS 0.009981f
C408 B.n368 VSUBS 0.009981f
C409 B.n369 VSUBS 0.009981f
C410 B.n370 VSUBS 0.009981f
C411 B.n371 VSUBS 0.009981f
C412 B.n372 VSUBS 0.009981f
C413 B.n373 VSUBS 0.009981f
C414 B.n374 VSUBS 0.009981f
C415 B.n375 VSUBS 0.009981f
C416 B.n376 VSUBS 0.009981f
C417 B.n377 VSUBS 0.009981f
C418 B.n378 VSUBS 0.009981f
C419 B.n379 VSUBS 0.009981f
C420 B.n380 VSUBS 0.009981f
C421 B.n381 VSUBS 0.009981f
C422 B.n382 VSUBS 0.009981f
C423 B.n383 VSUBS 0.009981f
C424 B.n384 VSUBS 0.009981f
C425 B.n385 VSUBS 0.009981f
C426 B.n386 VSUBS 0.009981f
C427 B.n387 VSUBS 0.009981f
C428 B.n388 VSUBS 0.025061f
C429 B.n389 VSUBS 0.023964f
C430 B.n390 VSUBS 0.025061f
C431 B.n391 VSUBS 0.009981f
C432 B.n392 VSUBS 0.009981f
C433 B.n393 VSUBS 0.009981f
C434 B.n394 VSUBS 0.009981f
C435 B.n395 VSUBS 0.009981f
C436 B.n396 VSUBS 0.009981f
C437 B.n397 VSUBS 0.009981f
C438 B.n398 VSUBS 0.009981f
C439 B.n399 VSUBS 0.009981f
C440 B.n400 VSUBS 0.009981f
C441 B.n401 VSUBS 0.009981f
C442 B.n402 VSUBS 0.009981f
C443 B.n403 VSUBS 0.009981f
C444 B.n404 VSUBS 0.009981f
C445 B.n405 VSUBS 0.009981f
C446 B.n406 VSUBS 0.009981f
C447 B.n407 VSUBS 0.009981f
C448 B.n408 VSUBS 0.009981f
C449 B.n409 VSUBS 0.009981f
C450 B.n410 VSUBS 0.009981f
C451 B.n411 VSUBS 0.006899f
C452 B.n412 VSUBS 0.023125f
C453 B.n413 VSUBS 0.008073f
C454 B.n414 VSUBS 0.009981f
C455 B.n415 VSUBS 0.009981f
C456 B.n416 VSUBS 0.009981f
C457 B.n417 VSUBS 0.009981f
C458 B.n418 VSUBS 0.009981f
C459 B.n419 VSUBS 0.009981f
C460 B.n420 VSUBS 0.009981f
C461 B.n421 VSUBS 0.009981f
C462 B.n422 VSUBS 0.009981f
C463 B.n423 VSUBS 0.009981f
C464 B.n424 VSUBS 0.009981f
C465 B.n425 VSUBS 0.008073f
C466 B.n426 VSUBS 0.023125f
C467 B.n427 VSUBS 0.006899f
C468 B.n428 VSUBS 0.009981f
C469 B.n429 VSUBS 0.009981f
C470 B.n430 VSUBS 0.009981f
C471 B.n431 VSUBS 0.009981f
C472 B.n432 VSUBS 0.009981f
C473 B.n433 VSUBS 0.009981f
C474 B.n434 VSUBS 0.009981f
C475 B.n435 VSUBS 0.009981f
C476 B.n436 VSUBS 0.009981f
C477 B.n437 VSUBS 0.009981f
C478 B.n438 VSUBS 0.009981f
C479 B.n439 VSUBS 0.009981f
C480 B.n440 VSUBS 0.009981f
C481 B.n441 VSUBS 0.009981f
C482 B.n442 VSUBS 0.009981f
C483 B.n443 VSUBS 0.009981f
C484 B.n444 VSUBS 0.009981f
C485 B.n445 VSUBS 0.009981f
C486 B.n446 VSUBS 0.009981f
C487 B.n447 VSUBS 0.009981f
C488 B.n448 VSUBS 0.025061f
C489 B.n449 VSUBS 0.025061f
C490 B.n450 VSUBS 0.023964f
C491 B.n451 VSUBS 0.009981f
C492 B.n452 VSUBS 0.009981f
C493 B.n453 VSUBS 0.009981f
C494 B.n454 VSUBS 0.009981f
C495 B.n455 VSUBS 0.009981f
C496 B.n456 VSUBS 0.009981f
C497 B.n457 VSUBS 0.009981f
C498 B.n458 VSUBS 0.009981f
C499 B.n459 VSUBS 0.009981f
C500 B.n460 VSUBS 0.009981f
C501 B.n461 VSUBS 0.009981f
C502 B.n462 VSUBS 0.009981f
C503 B.n463 VSUBS 0.009981f
C504 B.n464 VSUBS 0.009981f
C505 B.n465 VSUBS 0.009981f
C506 B.n466 VSUBS 0.009981f
C507 B.n467 VSUBS 0.009981f
C508 B.n468 VSUBS 0.009981f
C509 B.n469 VSUBS 0.009981f
C510 B.n470 VSUBS 0.009981f
C511 B.n471 VSUBS 0.009981f
C512 B.n472 VSUBS 0.009981f
C513 B.n473 VSUBS 0.009981f
C514 B.n474 VSUBS 0.009981f
C515 B.n475 VSUBS 0.009981f
C516 B.n476 VSUBS 0.009981f
C517 B.n477 VSUBS 0.009981f
C518 B.n478 VSUBS 0.009981f
C519 B.n479 VSUBS 0.009981f
C520 B.n480 VSUBS 0.009981f
C521 B.n481 VSUBS 0.009981f
C522 B.n482 VSUBS 0.009981f
C523 B.n483 VSUBS 0.009981f
C524 B.n484 VSUBS 0.009981f
C525 B.n485 VSUBS 0.009981f
C526 B.n486 VSUBS 0.009981f
C527 B.n487 VSUBS 0.009981f
C528 B.n488 VSUBS 0.009981f
C529 B.n489 VSUBS 0.009981f
C530 B.n490 VSUBS 0.009981f
C531 B.n491 VSUBS 0.009981f
C532 B.n492 VSUBS 0.009981f
C533 B.n493 VSUBS 0.009981f
C534 B.n494 VSUBS 0.009981f
C535 B.n495 VSUBS 0.009981f
C536 B.n496 VSUBS 0.009981f
C537 B.n497 VSUBS 0.009981f
C538 B.n498 VSUBS 0.009981f
C539 B.n499 VSUBS 0.009981f
C540 B.n500 VSUBS 0.009981f
C541 B.n501 VSUBS 0.009981f
C542 B.n502 VSUBS 0.009981f
C543 B.n503 VSUBS 0.009981f
C544 B.n504 VSUBS 0.009981f
C545 B.n505 VSUBS 0.009981f
C546 B.n506 VSUBS 0.009981f
C547 B.n507 VSUBS 0.009981f
C548 B.n508 VSUBS 0.009981f
C549 B.n509 VSUBS 0.009981f
C550 B.n510 VSUBS 0.009981f
C551 B.n511 VSUBS 0.009981f
C552 B.n512 VSUBS 0.009981f
C553 B.n513 VSUBS 0.009981f
C554 B.n514 VSUBS 0.009981f
C555 B.n515 VSUBS 0.022601f
C556 VDD1.t2 VSUBS 0.047623f
C557 VDD1.t0 VSUBS 0.047623f
C558 VDD1.n0 VSUBS 0.246579f
C559 VDD1.t1 VSUBS 0.047623f
C560 VDD1.t3 VSUBS 0.047623f
C561 VDD1.n1 VSUBS 0.458026f
C562 VP.t0 VSUBS 1.14168f
C563 VP.n0 VSUBS 0.649676f
C564 VP.n1 VSUBS 0.043775f
C565 VP.n2 VSUBS 0.063904f
C566 VP.n3 VSUBS 0.043775f
C567 VP.n4 VSUBS 0.060236f
C568 VP.t1 VSUBS 1.67422f
C569 VP.t3 VSUBS 1.65477f
C570 VP.n5 VSUBS 3.35245f
C571 VP.t2 VSUBS 1.14168f
C572 VP.n6 VSUBS 0.649676f
C573 VP.n7 VSUBS 2.1406f
C574 VP.n8 VSUBS 0.070652f
C575 VP.n9 VSUBS 0.043775f
C576 VP.n10 VSUBS 0.081586f
C577 VP.n11 VSUBS 0.081586f
C578 VP.n12 VSUBS 0.063904f
C579 VP.n13 VSUBS 0.043775f
C580 VP.n14 VSUBS 0.043775f
C581 VP.n15 VSUBS 0.043775f
C582 VP.n16 VSUBS 0.081586f
C583 VP.n17 VSUBS 0.081586f
C584 VP.n18 VSUBS 0.060236f
C585 VP.n19 VSUBS 0.070652f
C586 VP.n20 VSUBS 0.117946f
C587 VTAIL.t4 VSUBS 0.468505f
C588 VTAIL.n0 VSUBS 0.650886f
C589 VTAIL.t1 VSUBS 0.468505f
C590 VTAIL.n1 VSUBS 0.814868f
C591 VTAIL.t2 VSUBS 0.468505f
C592 VTAIL.n2 VSUBS 1.77312f
C593 VTAIL.t7 VSUBS 0.468506f
C594 VTAIL.n3 VSUBS 1.77312f
C595 VTAIL.t6 VSUBS 0.468506f
C596 VTAIL.n4 VSUBS 0.814867f
C597 VTAIL.t0 VSUBS 0.468506f
C598 VTAIL.n5 VSUBS 0.814867f
C599 VTAIL.t3 VSUBS 0.468505f
C600 VTAIL.n6 VSUBS 1.77312f
C601 VTAIL.t5 VSUBS 0.468505f
C602 VTAIL.n7 VSUBS 1.59759f
C603 VDD2.t3 VSUBS 0.048608f
C604 VDD2.t1 VSUBS 0.048608f
C605 VDD2.n0 VSUBS 0.456284f
C606 VDD2.t0 VSUBS 0.048608f
C607 VDD2.t2 VSUBS 0.048608f
C608 VDD2.n1 VSUBS 0.251468f
C609 VDD2.n2 VSUBS 2.65852f
C610 VN.t2 VSUBS 1.59887f
C611 VN.t3 VSUBS 1.61766f
C612 VN.n0 VSUBS 0.992767f
C613 VN.t1 VSUBS 1.61766f
C614 VN.t0 VSUBS 1.59887f
C615 VN.n1 VSUBS 3.25707f
.ends

