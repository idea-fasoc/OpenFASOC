* NGSPICE file created from diff_pair_sample_1287.ext - technology: sky130A

.subckt diff_pair_sample_1287 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=1.62
X2 VTAIL.t10 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=1.14345 ps=7.26 w=6.93 l=1.62
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=1.62
X4 VTAIL.t3 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=1.14345 ps=7.26 w=6.93 l=1.62
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=1.62
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=1.62
X7 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X8 VDD2.t5 VN.t2 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=2.7027 ps=14.64 w=6.93 l=1.62
X9 VTAIL.t12 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X10 VDD2.t3 VN.t4 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X11 VTAIL.t7 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X12 VDD2.t2 VN.t5 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=2.7027 ps=14.64 w=6.93 l=1.62
X13 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=1.14345 ps=7.26 w=6.93 l=1.62
X14 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X15 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=2.7027 ps=14.64 w=6.93 l=1.62
X16 VDD1.t1 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
X17 VTAIL.t14 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=1.14345 ps=7.26 w=6.93 l=1.62
X18 VDD1.t0 VP.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=2.7027 ps=14.64 w=6.93 l=1.62
X19 VTAIL.t9 VN.t7 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.14345 pd=7.26 as=1.14345 ps=7.26 w=6.93 l=1.62
R0 VN.n20 VN.n19 177.204
R1 VN.n41 VN.n40 177.204
R2 VN.n39 VN.n21 161.3
R3 VN.n38 VN.n37 161.3
R4 VN.n36 VN.n22 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n32 VN.n23 161.3
R7 VN.n31 VN.n30 161.3
R8 VN.n29 VN.n24 161.3
R9 VN.n28 VN.n27 161.3
R10 VN.n18 VN.n0 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n1 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n11 VN.n2 161.3
R15 VN.n10 VN.n9 161.3
R16 VN.n8 VN.n3 161.3
R17 VN.n7 VN.n6 161.3
R18 VN.n4 VN.t1 136.07
R19 VN.n25 VN.t2 136.07
R20 VN.n5 VN.t0 103.094
R21 VN.n12 VN.t7 103.094
R22 VN.n19 VN.t5 103.094
R23 VN.n26 VN.t3 103.094
R24 VN.n33 VN.t4 103.094
R25 VN.n40 VN.t6 103.094
R26 VN.n10 VN.n3 56.5193
R27 VN.n17 VN.n1 56.5193
R28 VN.n31 VN.n24 56.5193
R29 VN.n38 VN.n22 56.5193
R30 VN.n5 VN.n4 55.22
R31 VN.n26 VN.n25 55.22
R32 VN VN.n41 42.7827
R33 VN.n6 VN.n3 24.4675
R34 VN.n11 VN.n10 24.4675
R35 VN.n13 VN.n1 24.4675
R36 VN.n18 VN.n17 24.4675
R37 VN.n27 VN.n24 24.4675
R38 VN.n34 VN.n22 24.4675
R39 VN.n32 VN.n31 24.4675
R40 VN.n39 VN.n38 24.4675
R41 VN.n28 VN.n25 17.9267
R42 VN.n7 VN.n4 17.9267
R43 VN.n13 VN.n12 13.4574
R44 VN.n34 VN.n33 13.4574
R45 VN.n6 VN.n5 11.0107
R46 VN.n12 VN.n11 11.0107
R47 VN.n27 VN.n26 11.0107
R48 VN.n33 VN.n32 11.0107
R49 VN.n19 VN.n18 8.56395
R50 VN.n40 VN.n39 8.56395
R51 VN.n41 VN.n21 0.189894
R52 VN.n37 VN.n21 0.189894
R53 VN.n37 VN.n36 0.189894
R54 VN.n36 VN.n35 0.189894
R55 VN.n35 VN.n23 0.189894
R56 VN.n30 VN.n23 0.189894
R57 VN.n30 VN.n29 0.189894
R58 VN.n29 VN.n28 0.189894
R59 VN.n8 VN.n7 0.189894
R60 VN.n9 VN.n8 0.189894
R61 VN.n9 VN.n2 0.189894
R62 VN.n14 VN.n2 0.189894
R63 VN.n15 VN.n14 0.189894
R64 VN.n16 VN.n15 0.189894
R65 VN.n16 VN.n0 0.189894
R66 VN.n20 VN.n0 0.189894
R67 VN VN.n20 0.0516364
R68 VTAIL.n11 VTAIL.t0 55.271
R69 VTAIL.n10 VTAIL.t8 55.271
R70 VTAIL.n7 VTAIL.t14 55.271
R71 VTAIL.n15 VTAIL.t11 55.2709
R72 VTAIL.n2 VTAIL.t10 55.2709
R73 VTAIL.n3 VTAIL.t2 55.2709
R74 VTAIL.n6 VTAIL.t3 55.2709
R75 VTAIL.n14 VTAIL.t6 55.2709
R76 VTAIL.n13 VTAIL.n12 52.4139
R77 VTAIL.n9 VTAIL.n8 52.4139
R78 VTAIL.n1 VTAIL.n0 52.4128
R79 VTAIL.n5 VTAIL.n4 52.4128
R80 VTAIL.n15 VTAIL.n14 20.0221
R81 VTAIL.n7 VTAIL.n6 20.0221
R82 VTAIL.n0 VTAIL.t15 2.85764
R83 VTAIL.n0 VTAIL.t9 2.85764
R84 VTAIL.n4 VTAIL.t5 2.85764
R85 VTAIL.n4 VTAIL.t7 2.85764
R86 VTAIL.n12 VTAIL.t4 2.85764
R87 VTAIL.n12 VTAIL.t1 2.85764
R88 VTAIL.n8 VTAIL.t13 2.85764
R89 VTAIL.n8 VTAIL.t12 2.85764
R90 VTAIL.n9 VTAIL.n7 1.68153
R91 VTAIL.n10 VTAIL.n9 1.68153
R92 VTAIL.n13 VTAIL.n11 1.68153
R93 VTAIL.n14 VTAIL.n13 1.68153
R94 VTAIL.n6 VTAIL.n5 1.68153
R95 VTAIL.n5 VTAIL.n3 1.68153
R96 VTAIL.n2 VTAIL.n1 1.68153
R97 VTAIL VTAIL.n15 1.62334
R98 VTAIL.n11 VTAIL.n10 0.470328
R99 VTAIL.n3 VTAIL.n2 0.470328
R100 VTAIL VTAIL.n1 0.0586897
R101 VDD2.n2 VDD2.n1 69.8767
R102 VDD2.n2 VDD2.n0 69.8767
R103 VDD2 VDD2.n5 69.8749
R104 VDD2.n4 VDD2.n3 69.0926
R105 VDD2.n4 VDD2.n2 37.2541
R106 VDD2.n5 VDD2.t4 2.85764
R107 VDD2.n5 VDD2.t5 2.85764
R108 VDD2.n3 VDD2.t1 2.85764
R109 VDD2.n3 VDD2.t3 2.85764
R110 VDD2.n1 VDD2.t0 2.85764
R111 VDD2.n1 VDD2.t2 2.85764
R112 VDD2.n0 VDD2.t6 2.85764
R113 VDD2.n0 VDD2.t7 2.85764
R114 VDD2 VDD2.n4 0.899207
R115 B.n625 B.n624 585
R116 B.n626 B.n625 585
R117 B.n230 B.n101 585
R118 B.n229 B.n228 585
R119 B.n227 B.n226 585
R120 B.n225 B.n224 585
R121 B.n223 B.n222 585
R122 B.n221 B.n220 585
R123 B.n219 B.n218 585
R124 B.n217 B.n216 585
R125 B.n215 B.n214 585
R126 B.n213 B.n212 585
R127 B.n211 B.n210 585
R128 B.n209 B.n208 585
R129 B.n207 B.n206 585
R130 B.n205 B.n204 585
R131 B.n203 B.n202 585
R132 B.n201 B.n200 585
R133 B.n199 B.n198 585
R134 B.n197 B.n196 585
R135 B.n195 B.n194 585
R136 B.n193 B.n192 585
R137 B.n191 B.n190 585
R138 B.n189 B.n188 585
R139 B.n187 B.n186 585
R140 B.n185 B.n184 585
R141 B.n183 B.n182 585
R142 B.n181 B.n180 585
R143 B.n179 B.n178 585
R144 B.n177 B.n176 585
R145 B.n175 B.n174 585
R146 B.n173 B.n172 585
R147 B.n171 B.n170 585
R148 B.n169 B.n168 585
R149 B.n167 B.n166 585
R150 B.n165 B.n164 585
R151 B.n163 B.n162 585
R152 B.n160 B.n159 585
R153 B.n158 B.n157 585
R154 B.n156 B.n155 585
R155 B.n154 B.n153 585
R156 B.n152 B.n151 585
R157 B.n150 B.n149 585
R158 B.n148 B.n147 585
R159 B.n146 B.n145 585
R160 B.n144 B.n143 585
R161 B.n142 B.n141 585
R162 B.n140 B.n139 585
R163 B.n138 B.n137 585
R164 B.n136 B.n135 585
R165 B.n134 B.n133 585
R166 B.n132 B.n131 585
R167 B.n130 B.n129 585
R168 B.n128 B.n127 585
R169 B.n126 B.n125 585
R170 B.n124 B.n123 585
R171 B.n122 B.n121 585
R172 B.n120 B.n119 585
R173 B.n118 B.n117 585
R174 B.n116 B.n115 585
R175 B.n114 B.n113 585
R176 B.n112 B.n111 585
R177 B.n110 B.n109 585
R178 B.n108 B.n107 585
R179 B.n623 B.n69 585
R180 B.n627 B.n69 585
R181 B.n622 B.n68 585
R182 B.n628 B.n68 585
R183 B.n621 B.n620 585
R184 B.n620 B.n64 585
R185 B.n619 B.n63 585
R186 B.n634 B.n63 585
R187 B.n618 B.n62 585
R188 B.n635 B.n62 585
R189 B.n617 B.n61 585
R190 B.n636 B.n61 585
R191 B.n616 B.n615 585
R192 B.n615 B.n60 585
R193 B.n614 B.n56 585
R194 B.n642 B.n56 585
R195 B.n613 B.n55 585
R196 B.n643 B.n55 585
R197 B.n612 B.n54 585
R198 B.n644 B.n54 585
R199 B.n611 B.n610 585
R200 B.n610 B.n50 585
R201 B.n609 B.n49 585
R202 B.n650 B.n49 585
R203 B.n608 B.n48 585
R204 B.n651 B.n48 585
R205 B.n607 B.n47 585
R206 B.n652 B.n47 585
R207 B.n606 B.n605 585
R208 B.n605 B.n43 585
R209 B.n604 B.n42 585
R210 B.n658 B.n42 585
R211 B.n603 B.n41 585
R212 B.n659 B.n41 585
R213 B.n602 B.n40 585
R214 B.n660 B.n40 585
R215 B.n601 B.n600 585
R216 B.n600 B.n36 585
R217 B.n599 B.n35 585
R218 B.n666 B.n35 585
R219 B.n598 B.n34 585
R220 B.n667 B.n34 585
R221 B.n597 B.n33 585
R222 B.n668 B.n33 585
R223 B.n596 B.n595 585
R224 B.n595 B.n29 585
R225 B.n594 B.n28 585
R226 B.n674 B.n28 585
R227 B.n593 B.n27 585
R228 B.n675 B.n27 585
R229 B.n592 B.n26 585
R230 B.n676 B.n26 585
R231 B.n591 B.n590 585
R232 B.n590 B.n25 585
R233 B.n589 B.n21 585
R234 B.n682 B.n21 585
R235 B.n588 B.n20 585
R236 B.n683 B.n20 585
R237 B.n587 B.n19 585
R238 B.n684 B.n19 585
R239 B.n586 B.n585 585
R240 B.n585 B.n15 585
R241 B.n584 B.n14 585
R242 B.n690 B.n14 585
R243 B.n583 B.n13 585
R244 B.n691 B.n13 585
R245 B.n582 B.n12 585
R246 B.n692 B.n12 585
R247 B.n581 B.n580 585
R248 B.n580 B.n8 585
R249 B.n579 B.n7 585
R250 B.n698 B.n7 585
R251 B.n578 B.n6 585
R252 B.n699 B.n6 585
R253 B.n577 B.n5 585
R254 B.n700 B.n5 585
R255 B.n576 B.n575 585
R256 B.n575 B.n4 585
R257 B.n574 B.n231 585
R258 B.n574 B.n573 585
R259 B.n564 B.n232 585
R260 B.n233 B.n232 585
R261 B.n566 B.n565 585
R262 B.n567 B.n566 585
R263 B.n563 B.n237 585
R264 B.n241 B.n237 585
R265 B.n562 B.n561 585
R266 B.n561 B.n560 585
R267 B.n239 B.n238 585
R268 B.n240 B.n239 585
R269 B.n553 B.n552 585
R270 B.n554 B.n553 585
R271 B.n551 B.n246 585
R272 B.n246 B.n245 585
R273 B.n550 B.n549 585
R274 B.n549 B.n548 585
R275 B.n248 B.n247 585
R276 B.n541 B.n248 585
R277 B.n540 B.n539 585
R278 B.n542 B.n540 585
R279 B.n538 B.n253 585
R280 B.n253 B.n252 585
R281 B.n537 B.n536 585
R282 B.n536 B.n535 585
R283 B.n255 B.n254 585
R284 B.n256 B.n255 585
R285 B.n528 B.n527 585
R286 B.n529 B.n528 585
R287 B.n526 B.n261 585
R288 B.n261 B.n260 585
R289 B.n525 B.n524 585
R290 B.n524 B.n523 585
R291 B.n263 B.n262 585
R292 B.n264 B.n263 585
R293 B.n516 B.n515 585
R294 B.n517 B.n516 585
R295 B.n514 B.n269 585
R296 B.n269 B.n268 585
R297 B.n513 B.n512 585
R298 B.n512 B.n511 585
R299 B.n271 B.n270 585
R300 B.n272 B.n271 585
R301 B.n504 B.n503 585
R302 B.n505 B.n504 585
R303 B.n502 B.n277 585
R304 B.n277 B.n276 585
R305 B.n501 B.n500 585
R306 B.n500 B.n499 585
R307 B.n279 B.n278 585
R308 B.n280 B.n279 585
R309 B.n492 B.n491 585
R310 B.n493 B.n492 585
R311 B.n490 B.n285 585
R312 B.n285 B.n284 585
R313 B.n489 B.n488 585
R314 B.n488 B.n487 585
R315 B.n287 B.n286 585
R316 B.n480 B.n287 585
R317 B.n479 B.n478 585
R318 B.n481 B.n479 585
R319 B.n477 B.n292 585
R320 B.n292 B.n291 585
R321 B.n476 B.n475 585
R322 B.n475 B.n474 585
R323 B.n294 B.n293 585
R324 B.n295 B.n294 585
R325 B.n467 B.n466 585
R326 B.n468 B.n467 585
R327 B.n465 B.n300 585
R328 B.n300 B.n299 585
R329 B.n459 B.n458 585
R330 B.n457 B.n333 585
R331 B.n456 B.n332 585
R332 B.n461 B.n332 585
R333 B.n455 B.n454 585
R334 B.n453 B.n452 585
R335 B.n451 B.n450 585
R336 B.n449 B.n448 585
R337 B.n447 B.n446 585
R338 B.n445 B.n444 585
R339 B.n443 B.n442 585
R340 B.n441 B.n440 585
R341 B.n439 B.n438 585
R342 B.n437 B.n436 585
R343 B.n435 B.n434 585
R344 B.n433 B.n432 585
R345 B.n431 B.n430 585
R346 B.n429 B.n428 585
R347 B.n427 B.n426 585
R348 B.n425 B.n424 585
R349 B.n423 B.n422 585
R350 B.n421 B.n420 585
R351 B.n419 B.n418 585
R352 B.n417 B.n416 585
R353 B.n415 B.n414 585
R354 B.n413 B.n412 585
R355 B.n411 B.n410 585
R356 B.n409 B.n408 585
R357 B.n407 B.n406 585
R358 B.n405 B.n404 585
R359 B.n403 B.n402 585
R360 B.n401 B.n400 585
R361 B.n399 B.n398 585
R362 B.n397 B.n396 585
R363 B.n395 B.n394 585
R364 B.n393 B.n392 585
R365 B.n391 B.n390 585
R366 B.n388 B.n387 585
R367 B.n386 B.n385 585
R368 B.n384 B.n383 585
R369 B.n382 B.n381 585
R370 B.n380 B.n379 585
R371 B.n378 B.n377 585
R372 B.n376 B.n375 585
R373 B.n374 B.n373 585
R374 B.n372 B.n371 585
R375 B.n370 B.n369 585
R376 B.n368 B.n367 585
R377 B.n366 B.n365 585
R378 B.n364 B.n363 585
R379 B.n362 B.n361 585
R380 B.n360 B.n359 585
R381 B.n358 B.n357 585
R382 B.n356 B.n355 585
R383 B.n354 B.n353 585
R384 B.n352 B.n351 585
R385 B.n350 B.n349 585
R386 B.n348 B.n347 585
R387 B.n346 B.n345 585
R388 B.n344 B.n343 585
R389 B.n342 B.n341 585
R390 B.n340 B.n339 585
R391 B.n302 B.n301 585
R392 B.n464 B.n463 585
R393 B.n298 B.n297 585
R394 B.n299 B.n298 585
R395 B.n470 B.n469 585
R396 B.n469 B.n468 585
R397 B.n471 B.n296 585
R398 B.n296 B.n295 585
R399 B.n473 B.n472 585
R400 B.n474 B.n473 585
R401 B.n290 B.n289 585
R402 B.n291 B.n290 585
R403 B.n483 B.n482 585
R404 B.n482 B.n481 585
R405 B.n484 B.n288 585
R406 B.n480 B.n288 585
R407 B.n486 B.n485 585
R408 B.n487 B.n486 585
R409 B.n283 B.n282 585
R410 B.n284 B.n283 585
R411 B.n495 B.n494 585
R412 B.n494 B.n493 585
R413 B.n496 B.n281 585
R414 B.n281 B.n280 585
R415 B.n498 B.n497 585
R416 B.n499 B.n498 585
R417 B.n275 B.n274 585
R418 B.n276 B.n275 585
R419 B.n507 B.n506 585
R420 B.n506 B.n505 585
R421 B.n508 B.n273 585
R422 B.n273 B.n272 585
R423 B.n510 B.n509 585
R424 B.n511 B.n510 585
R425 B.n267 B.n266 585
R426 B.n268 B.n267 585
R427 B.n519 B.n518 585
R428 B.n518 B.n517 585
R429 B.n520 B.n265 585
R430 B.n265 B.n264 585
R431 B.n522 B.n521 585
R432 B.n523 B.n522 585
R433 B.n259 B.n258 585
R434 B.n260 B.n259 585
R435 B.n531 B.n530 585
R436 B.n530 B.n529 585
R437 B.n532 B.n257 585
R438 B.n257 B.n256 585
R439 B.n534 B.n533 585
R440 B.n535 B.n534 585
R441 B.n251 B.n250 585
R442 B.n252 B.n251 585
R443 B.n544 B.n543 585
R444 B.n543 B.n542 585
R445 B.n545 B.n249 585
R446 B.n541 B.n249 585
R447 B.n547 B.n546 585
R448 B.n548 B.n547 585
R449 B.n244 B.n243 585
R450 B.n245 B.n244 585
R451 B.n556 B.n555 585
R452 B.n555 B.n554 585
R453 B.n557 B.n242 585
R454 B.n242 B.n240 585
R455 B.n559 B.n558 585
R456 B.n560 B.n559 585
R457 B.n236 B.n235 585
R458 B.n241 B.n236 585
R459 B.n569 B.n568 585
R460 B.n568 B.n567 585
R461 B.n570 B.n234 585
R462 B.n234 B.n233 585
R463 B.n572 B.n571 585
R464 B.n573 B.n572 585
R465 B.n2 B.n0 585
R466 B.n4 B.n2 585
R467 B.n3 B.n1 585
R468 B.n699 B.n3 585
R469 B.n697 B.n696 585
R470 B.n698 B.n697 585
R471 B.n695 B.n9 585
R472 B.n9 B.n8 585
R473 B.n694 B.n693 585
R474 B.n693 B.n692 585
R475 B.n11 B.n10 585
R476 B.n691 B.n11 585
R477 B.n689 B.n688 585
R478 B.n690 B.n689 585
R479 B.n687 B.n16 585
R480 B.n16 B.n15 585
R481 B.n686 B.n685 585
R482 B.n685 B.n684 585
R483 B.n18 B.n17 585
R484 B.n683 B.n18 585
R485 B.n681 B.n680 585
R486 B.n682 B.n681 585
R487 B.n679 B.n22 585
R488 B.n25 B.n22 585
R489 B.n678 B.n677 585
R490 B.n677 B.n676 585
R491 B.n24 B.n23 585
R492 B.n675 B.n24 585
R493 B.n673 B.n672 585
R494 B.n674 B.n673 585
R495 B.n671 B.n30 585
R496 B.n30 B.n29 585
R497 B.n670 B.n669 585
R498 B.n669 B.n668 585
R499 B.n32 B.n31 585
R500 B.n667 B.n32 585
R501 B.n665 B.n664 585
R502 B.n666 B.n665 585
R503 B.n663 B.n37 585
R504 B.n37 B.n36 585
R505 B.n662 B.n661 585
R506 B.n661 B.n660 585
R507 B.n39 B.n38 585
R508 B.n659 B.n39 585
R509 B.n657 B.n656 585
R510 B.n658 B.n657 585
R511 B.n655 B.n44 585
R512 B.n44 B.n43 585
R513 B.n654 B.n653 585
R514 B.n653 B.n652 585
R515 B.n46 B.n45 585
R516 B.n651 B.n46 585
R517 B.n649 B.n648 585
R518 B.n650 B.n649 585
R519 B.n647 B.n51 585
R520 B.n51 B.n50 585
R521 B.n646 B.n645 585
R522 B.n645 B.n644 585
R523 B.n53 B.n52 585
R524 B.n643 B.n53 585
R525 B.n641 B.n640 585
R526 B.n642 B.n641 585
R527 B.n639 B.n57 585
R528 B.n60 B.n57 585
R529 B.n638 B.n637 585
R530 B.n637 B.n636 585
R531 B.n59 B.n58 585
R532 B.n635 B.n59 585
R533 B.n633 B.n632 585
R534 B.n634 B.n633 585
R535 B.n631 B.n65 585
R536 B.n65 B.n64 585
R537 B.n630 B.n629 585
R538 B.n629 B.n628 585
R539 B.n67 B.n66 585
R540 B.n627 B.n67 585
R541 B.n702 B.n701 585
R542 B.n701 B.n700 585
R543 B.n459 B.n298 463.671
R544 B.n107 B.n67 463.671
R545 B.n463 B.n300 463.671
R546 B.n625 B.n69 463.671
R547 B.n337 B.t19 308.954
R548 B.n334 B.t12 308.954
R549 B.n105 B.t16 308.954
R550 B.n102 B.t8 308.954
R551 B.n626 B.n100 256.663
R552 B.n626 B.n99 256.663
R553 B.n626 B.n98 256.663
R554 B.n626 B.n97 256.663
R555 B.n626 B.n96 256.663
R556 B.n626 B.n95 256.663
R557 B.n626 B.n94 256.663
R558 B.n626 B.n93 256.663
R559 B.n626 B.n92 256.663
R560 B.n626 B.n91 256.663
R561 B.n626 B.n90 256.663
R562 B.n626 B.n89 256.663
R563 B.n626 B.n88 256.663
R564 B.n626 B.n87 256.663
R565 B.n626 B.n86 256.663
R566 B.n626 B.n85 256.663
R567 B.n626 B.n84 256.663
R568 B.n626 B.n83 256.663
R569 B.n626 B.n82 256.663
R570 B.n626 B.n81 256.663
R571 B.n626 B.n80 256.663
R572 B.n626 B.n79 256.663
R573 B.n626 B.n78 256.663
R574 B.n626 B.n77 256.663
R575 B.n626 B.n76 256.663
R576 B.n626 B.n75 256.663
R577 B.n626 B.n74 256.663
R578 B.n626 B.n73 256.663
R579 B.n626 B.n72 256.663
R580 B.n626 B.n71 256.663
R581 B.n626 B.n70 256.663
R582 B.n461 B.n460 256.663
R583 B.n461 B.n303 256.663
R584 B.n461 B.n304 256.663
R585 B.n461 B.n305 256.663
R586 B.n461 B.n306 256.663
R587 B.n461 B.n307 256.663
R588 B.n461 B.n308 256.663
R589 B.n461 B.n309 256.663
R590 B.n461 B.n310 256.663
R591 B.n461 B.n311 256.663
R592 B.n461 B.n312 256.663
R593 B.n461 B.n313 256.663
R594 B.n461 B.n314 256.663
R595 B.n461 B.n315 256.663
R596 B.n461 B.n316 256.663
R597 B.n461 B.n317 256.663
R598 B.n461 B.n318 256.663
R599 B.n461 B.n319 256.663
R600 B.n461 B.n320 256.663
R601 B.n461 B.n321 256.663
R602 B.n461 B.n322 256.663
R603 B.n461 B.n323 256.663
R604 B.n461 B.n324 256.663
R605 B.n461 B.n325 256.663
R606 B.n461 B.n326 256.663
R607 B.n461 B.n327 256.663
R608 B.n461 B.n328 256.663
R609 B.n461 B.n329 256.663
R610 B.n461 B.n330 256.663
R611 B.n461 B.n331 256.663
R612 B.n462 B.n461 256.663
R613 B.n469 B.n298 163.367
R614 B.n469 B.n296 163.367
R615 B.n473 B.n296 163.367
R616 B.n473 B.n290 163.367
R617 B.n482 B.n290 163.367
R618 B.n482 B.n288 163.367
R619 B.n486 B.n288 163.367
R620 B.n486 B.n283 163.367
R621 B.n494 B.n283 163.367
R622 B.n494 B.n281 163.367
R623 B.n498 B.n281 163.367
R624 B.n498 B.n275 163.367
R625 B.n506 B.n275 163.367
R626 B.n506 B.n273 163.367
R627 B.n510 B.n273 163.367
R628 B.n510 B.n267 163.367
R629 B.n518 B.n267 163.367
R630 B.n518 B.n265 163.367
R631 B.n522 B.n265 163.367
R632 B.n522 B.n259 163.367
R633 B.n530 B.n259 163.367
R634 B.n530 B.n257 163.367
R635 B.n534 B.n257 163.367
R636 B.n534 B.n251 163.367
R637 B.n543 B.n251 163.367
R638 B.n543 B.n249 163.367
R639 B.n547 B.n249 163.367
R640 B.n547 B.n244 163.367
R641 B.n555 B.n244 163.367
R642 B.n555 B.n242 163.367
R643 B.n559 B.n242 163.367
R644 B.n559 B.n236 163.367
R645 B.n568 B.n236 163.367
R646 B.n568 B.n234 163.367
R647 B.n572 B.n234 163.367
R648 B.n572 B.n2 163.367
R649 B.n701 B.n2 163.367
R650 B.n701 B.n3 163.367
R651 B.n697 B.n3 163.367
R652 B.n697 B.n9 163.367
R653 B.n693 B.n9 163.367
R654 B.n693 B.n11 163.367
R655 B.n689 B.n11 163.367
R656 B.n689 B.n16 163.367
R657 B.n685 B.n16 163.367
R658 B.n685 B.n18 163.367
R659 B.n681 B.n18 163.367
R660 B.n681 B.n22 163.367
R661 B.n677 B.n22 163.367
R662 B.n677 B.n24 163.367
R663 B.n673 B.n24 163.367
R664 B.n673 B.n30 163.367
R665 B.n669 B.n30 163.367
R666 B.n669 B.n32 163.367
R667 B.n665 B.n32 163.367
R668 B.n665 B.n37 163.367
R669 B.n661 B.n37 163.367
R670 B.n661 B.n39 163.367
R671 B.n657 B.n39 163.367
R672 B.n657 B.n44 163.367
R673 B.n653 B.n44 163.367
R674 B.n653 B.n46 163.367
R675 B.n649 B.n46 163.367
R676 B.n649 B.n51 163.367
R677 B.n645 B.n51 163.367
R678 B.n645 B.n53 163.367
R679 B.n641 B.n53 163.367
R680 B.n641 B.n57 163.367
R681 B.n637 B.n57 163.367
R682 B.n637 B.n59 163.367
R683 B.n633 B.n59 163.367
R684 B.n633 B.n65 163.367
R685 B.n629 B.n65 163.367
R686 B.n629 B.n67 163.367
R687 B.n333 B.n332 163.367
R688 B.n454 B.n332 163.367
R689 B.n452 B.n451 163.367
R690 B.n448 B.n447 163.367
R691 B.n444 B.n443 163.367
R692 B.n440 B.n439 163.367
R693 B.n436 B.n435 163.367
R694 B.n432 B.n431 163.367
R695 B.n428 B.n427 163.367
R696 B.n424 B.n423 163.367
R697 B.n420 B.n419 163.367
R698 B.n416 B.n415 163.367
R699 B.n412 B.n411 163.367
R700 B.n408 B.n407 163.367
R701 B.n404 B.n403 163.367
R702 B.n400 B.n399 163.367
R703 B.n396 B.n395 163.367
R704 B.n392 B.n391 163.367
R705 B.n387 B.n386 163.367
R706 B.n383 B.n382 163.367
R707 B.n379 B.n378 163.367
R708 B.n375 B.n374 163.367
R709 B.n371 B.n370 163.367
R710 B.n367 B.n366 163.367
R711 B.n363 B.n362 163.367
R712 B.n359 B.n358 163.367
R713 B.n355 B.n354 163.367
R714 B.n351 B.n350 163.367
R715 B.n347 B.n346 163.367
R716 B.n343 B.n342 163.367
R717 B.n339 B.n302 163.367
R718 B.n467 B.n300 163.367
R719 B.n467 B.n294 163.367
R720 B.n475 B.n294 163.367
R721 B.n475 B.n292 163.367
R722 B.n479 B.n292 163.367
R723 B.n479 B.n287 163.367
R724 B.n488 B.n287 163.367
R725 B.n488 B.n285 163.367
R726 B.n492 B.n285 163.367
R727 B.n492 B.n279 163.367
R728 B.n500 B.n279 163.367
R729 B.n500 B.n277 163.367
R730 B.n504 B.n277 163.367
R731 B.n504 B.n271 163.367
R732 B.n512 B.n271 163.367
R733 B.n512 B.n269 163.367
R734 B.n516 B.n269 163.367
R735 B.n516 B.n263 163.367
R736 B.n524 B.n263 163.367
R737 B.n524 B.n261 163.367
R738 B.n528 B.n261 163.367
R739 B.n528 B.n255 163.367
R740 B.n536 B.n255 163.367
R741 B.n536 B.n253 163.367
R742 B.n540 B.n253 163.367
R743 B.n540 B.n248 163.367
R744 B.n549 B.n248 163.367
R745 B.n549 B.n246 163.367
R746 B.n553 B.n246 163.367
R747 B.n553 B.n239 163.367
R748 B.n561 B.n239 163.367
R749 B.n561 B.n237 163.367
R750 B.n566 B.n237 163.367
R751 B.n566 B.n232 163.367
R752 B.n574 B.n232 163.367
R753 B.n575 B.n574 163.367
R754 B.n575 B.n5 163.367
R755 B.n6 B.n5 163.367
R756 B.n7 B.n6 163.367
R757 B.n580 B.n7 163.367
R758 B.n580 B.n12 163.367
R759 B.n13 B.n12 163.367
R760 B.n14 B.n13 163.367
R761 B.n585 B.n14 163.367
R762 B.n585 B.n19 163.367
R763 B.n20 B.n19 163.367
R764 B.n21 B.n20 163.367
R765 B.n590 B.n21 163.367
R766 B.n590 B.n26 163.367
R767 B.n27 B.n26 163.367
R768 B.n28 B.n27 163.367
R769 B.n595 B.n28 163.367
R770 B.n595 B.n33 163.367
R771 B.n34 B.n33 163.367
R772 B.n35 B.n34 163.367
R773 B.n600 B.n35 163.367
R774 B.n600 B.n40 163.367
R775 B.n41 B.n40 163.367
R776 B.n42 B.n41 163.367
R777 B.n605 B.n42 163.367
R778 B.n605 B.n47 163.367
R779 B.n48 B.n47 163.367
R780 B.n49 B.n48 163.367
R781 B.n610 B.n49 163.367
R782 B.n610 B.n54 163.367
R783 B.n55 B.n54 163.367
R784 B.n56 B.n55 163.367
R785 B.n615 B.n56 163.367
R786 B.n615 B.n61 163.367
R787 B.n62 B.n61 163.367
R788 B.n63 B.n62 163.367
R789 B.n620 B.n63 163.367
R790 B.n620 B.n68 163.367
R791 B.n69 B.n68 163.367
R792 B.n111 B.n110 163.367
R793 B.n115 B.n114 163.367
R794 B.n119 B.n118 163.367
R795 B.n123 B.n122 163.367
R796 B.n127 B.n126 163.367
R797 B.n131 B.n130 163.367
R798 B.n135 B.n134 163.367
R799 B.n139 B.n138 163.367
R800 B.n143 B.n142 163.367
R801 B.n147 B.n146 163.367
R802 B.n151 B.n150 163.367
R803 B.n155 B.n154 163.367
R804 B.n159 B.n158 163.367
R805 B.n164 B.n163 163.367
R806 B.n168 B.n167 163.367
R807 B.n172 B.n171 163.367
R808 B.n176 B.n175 163.367
R809 B.n180 B.n179 163.367
R810 B.n184 B.n183 163.367
R811 B.n188 B.n187 163.367
R812 B.n192 B.n191 163.367
R813 B.n196 B.n195 163.367
R814 B.n200 B.n199 163.367
R815 B.n204 B.n203 163.367
R816 B.n208 B.n207 163.367
R817 B.n212 B.n211 163.367
R818 B.n216 B.n215 163.367
R819 B.n220 B.n219 163.367
R820 B.n224 B.n223 163.367
R821 B.n228 B.n227 163.367
R822 B.n625 B.n101 163.367
R823 B.n337 B.t21 109.332
R824 B.n102 B.t10 109.332
R825 B.n334 B.t15 109.326
R826 B.n105 B.t17 109.326
R827 B.n461 B.n299 98.2389
R828 B.n627 B.n626 98.2389
R829 B.n460 B.n459 71.676
R830 B.n454 B.n303 71.676
R831 B.n451 B.n304 71.676
R832 B.n447 B.n305 71.676
R833 B.n443 B.n306 71.676
R834 B.n439 B.n307 71.676
R835 B.n435 B.n308 71.676
R836 B.n431 B.n309 71.676
R837 B.n427 B.n310 71.676
R838 B.n423 B.n311 71.676
R839 B.n419 B.n312 71.676
R840 B.n415 B.n313 71.676
R841 B.n411 B.n314 71.676
R842 B.n407 B.n315 71.676
R843 B.n403 B.n316 71.676
R844 B.n399 B.n317 71.676
R845 B.n395 B.n318 71.676
R846 B.n391 B.n319 71.676
R847 B.n386 B.n320 71.676
R848 B.n382 B.n321 71.676
R849 B.n378 B.n322 71.676
R850 B.n374 B.n323 71.676
R851 B.n370 B.n324 71.676
R852 B.n366 B.n325 71.676
R853 B.n362 B.n326 71.676
R854 B.n358 B.n327 71.676
R855 B.n354 B.n328 71.676
R856 B.n350 B.n329 71.676
R857 B.n346 B.n330 71.676
R858 B.n342 B.n331 71.676
R859 B.n462 B.n302 71.676
R860 B.n107 B.n70 71.676
R861 B.n111 B.n71 71.676
R862 B.n115 B.n72 71.676
R863 B.n119 B.n73 71.676
R864 B.n123 B.n74 71.676
R865 B.n127 B.n75 71.676
R866 B.n131 B.n76 71.676
R867 B.n135 B.n77 71.676
R868 B.n139 B.n78 71.676
R869 B.n143 B.n79 71.676
R870 B.n147 B.n80 71.676
R871 B.n151 B.n81 71.676
R872 B.n155 B.n82 71.676
R873 B.n159 B.n83 71.676
R874 B.n164 B.n84 71.676
R875 B.n168 B.n85 71.676
R876 B.n172 B.n86 71.676
R877 B.n176 B.n87 71.676
R878 B.n180 B.n88 71.676
R879 B.n184 B.n89 71.676
R880 B.n188 B.n90 71.676
R881 B.n192 B.n91 71.676
R882 B.n196 B.n92 71.676
R883 B.n200 B.n93 71.676
R884 B.n204 B.n94 71.676
R885 B.n208 B.n95 71.676
R886 B.n212 B.n96 71.676
R887 B.n216 B.n97 71.676
R888 B.n220 B.n98 71.676
R889 B.n224 B.n99 71.676
R890 B.n228 B.n100 71.676
R891 B.n101 B.n100 71.676
R892 B.n227 B.n99 71.676
R893 B.n223 B.n98 71.676
R894 B.n219 B.n97 71.676
R895 B.n215 B.n96 71.676
R896 B.n211 B.n95 71.676
R897 B.n207 B.n94 71.676
R898 B.n203 B.n93 71.676
R899 B.n199 B.n92 71.676
R900 B.n195 B.n91 71.676
R901 B.n191 B.n90 71.676
R902 B.n187 B.n89 71.676
R903 B.n183 B.n88 71.676
R904 B.n179 B.n87 71.676
R905 B.n175 B.n86 71.676
R906 B.n171 B.n85 71.676
R907 B.n167 B.n84 71.676
R908 B.n163 B.n83 71.676
R909 B.n158 B.n82 71.676
R910 B.n154 B.n81 71.676
R911 B.n150 B.n80 71.676
R912 B.n146 B.n79 71.676
R913 B.n142 B.n78 71.676
R914 B.n138 B.n77 71.676
R915 B.n134 B.n76 71.676
R916 B.n130 B.n75 71.676
R917 B.n126 B.n74 71.676
R918 B.n122 B.n73 71.676
R919 B.n118 B.n72 71.676
R920 B.n114 B.n71 71.676
R921 B.n110 B.n70 71.676
R922 B.n460 B.n333 71.676
R923 B.n452 B.n303 71.676
R924 B.n448 B.n304 71.676
R925 B.n444 B.n305 71.676
R926 B.n440 B.n306 71.676
R927 B.n436 B.n307 71.676
R928 B.n432 B.n308 71.676
R929 B.n428 B.n309 71.676
R930 B.n424 B.n310 71.676
R931 B.n420 B.n311 71.676
R932 B.n416 B.n312 71.676
R933 B.n412 B.n313 71.676
R934 B.n408 B.n314 71.676
R935 B.n404 B.n315 71.676
R936 B.n400 B.n316 71.676
R937 B.n396 B.n317 71.676
R938 B.n392 B.n318 71.676
R939 B.n387 B.n319 71.676
R940 B.n383 B.n320 71.676
R941 B.n379 B.n321 71.676
R942 B.n375 B.n322 71.676
R943 B.n371 B.n323 71.676
R944 B.n367 B.n324 71.676
R945 B.n363 B.n325 71.676
R946 B.n359 B.n326 71.676
R947 B.n355 B.n327 71.676
R948 B.n351 B.n328 71.676
R949 B.n347 B.n329 71.676
R950 B.n343 B.n330 71.676
R951 B.n339 B.n331 71.676
R952 B.n463 B.n462 71.676
R953 B.n338 B.t20 71.5148
R954 B.n103 B.t11 71.5148
R955 B.n335 B.t14 71.507
R956 B.n106 B.t18 71.507
R957 B.n468 B.n299 61.2869
R958 B.n468 B.n295 61.2869
R959 B.n474 B.n295 61.2869
R960 B.n474 B.n291 61.2869
R961 B.n481 B.n291 61.2869
R962 B.n481 B.n480 61.2869
R963 B.n487 B.n284 61.2869
R964 B.n493 B.n284 61.2869
R965 B.n493 B.n280 61.2869
R966 B.n499 B.n280 61.2869
R967 B.n499 B.n276 61.2869
R968 B.n505 B.n276 61.2869
R969 B.n505 B.n272 61.2869
R970 B.n511 B.n272 61.2869
R971 B.n517 B.n268 61.2869
R972 B.n517 B.n264 61.2869
R973 B.n523 B.n264 61.2869
R974 B.n523 B.n260 61.2869
R975 B.n529 B.n260 61.2869
R976 B.n535 B.n256 61.2869
R977 B.n535 B.n252 61.2869
R978 B.n542 B.n252 61.2869
R979 B.n542 B.n541 61.2869
R980 B.n548 B.n245 61.2869
R981 B.n554 B.n245 61.2869
R982 B.n554 B.n240 61.2869
R983 B.n560 B.n240 61.2869
R984 B.n560 B.n241 61.2869
R985 B.n567 B.n233 61.2869
R986 B.n573 B.n233 61.2869
R987 B.n573 B.n4 61.2869
R988 B.n700 B.n4 61.2869
R989 B.n700 B.n699 61.2869
R990 B.n699 B.n698 61.2869
R991 B.n698 B.n8 61.2869
R992 B.n692 B.n8 61.2869
R993 B.n691 B.n690 61.2869
R994 B.n690 B.n15 61.2869
R995 B.n684 B.n15 61.2869
R996 B.n684 B.n683 61.2869
R997 B.n683 B.n682 61.2869
R998 B.n676 B.n25 61.2869
R999 B.n676 B.n675 61.2869
R1000 B.n675 B.n674 61.2869
R1001 B.n674 B.n29 61.2869
R1002 B.n668 B.n667 61.2869
R1003 B.n667 B.n666 61.2869
R1004 B.n666 B.n36 61.2869
R1005 B.n660 B.n36 61.2869
R1006 B.n660 B.n659 61.2869
R1007 B.n658 B.n43 61.2869
R1008 B.n652 B.n43 61.2869
R1009 B.n652 B.n651 61.2869
R1010 B.n651 B.n650 61.2869
R1011 B.n650 B.n50 61.2869
R1012 B.n644 B.n50 61.2869
R1013 B.n644 B.n643 61.2869
R1014 B.n643 B.n642 61.2869
R1015 B.n636 B.n60 61.2869
R1016 B.n636 B.n635 61.2869
R1017 B.n635 B.n634 61.2869
R1018 B.n634 B.n64 61.2869
R1019 B.n628 B.n64 61.2869
R1020 B.n628 B.n627 61.2869
R1021 B.n389 B.n338 59.5399
R1022 B.n336 B.n335 59.5399
R1023 B.n161 B.n106 59.5399
R1024 B.n104 B.n103 59.5399
R1025 B.t5 B.n256 57.6818
R1026 B.t1 B.n29 57.6818
R1027 B.n541 B.t7 48.6691
R1028 B.n25 B.t4 48.6691
R1029 B.t3 B.n268 41.4589
R1030 B.n659 B.t6 41.4589
R1031 B.n487 B.t13 37.8538
R1032 B.n642 B.t9 37.8538
R1033 B.n338 B.n337 37.8187
R1034 B.n335 B.n334 37.8187
R1035 B.n106 B.n105 37.8187
R1036 B.n103 B.n102 37.8187
R1037 B.n241 B.t2 32.4462
R1038 B.t0 B.n691 32.4462
R1039 B.n108 B.n66 30.1273
R1040 B.n465 B.n464 30.1273
R1041 B.n458 B.n297 30.1273
R1042 B.n624 B.n623 30.1273
R1043 B.n567 B.t2 28.8411
R1044 B.n692 B.t0 28.8411
R1045 B.n480 B.t13 23.4335
R1046 B.n60 B.t9 23.4335
R1047 B.n511 B.t3 19.8284
R1048 B.t6 B.n658 19.8284
R1049 B B.n702 18.0485
R1050 B.n548 B.t7 12.6183
R1051 B.n682 B.t4 12.6183
R1052 B.n109 B.n108 10.6151
R1053 B.n112 B.n109 10.6151
R1054 B.n113 B.n112 10.6151
R1055 B.n116 B.n113 10.6151
R1056 B.n117 B.n116 10.6151
R1057 B.n120 B.n117 10.6151
R1058 B.n121 B.n120 10.6151
R1059 B.n124 B.n121 10.6151
R1060 B.n125 B.n124 10.6151
R1061 B.n128 B.n125 10.6151
R1062 B.n129 B.n128 10.6151
R1063 B.n132 B.n129 10.6151
R1064 B.n133 B.n132 10.6151
R1065 B.n136 B.n133 10.6151
R1066 B.n137 B.n136 10.6151
R1067 B.n140 B.n137 10.6151
R1068 B.n141 B.n140 10.6151
R1069 B.n144 B.n141 10.6151
R1070 B.n145 B.n144 10.6151
R1071 B.n148 B.n145 10.6151
R1072 B.n149 B.n148 10.6151
R1073 B.n152 B.n149 10.6151
R1074 B.n153 B.n152 10.6151
R1075 B.n156 B.n153 10.6151
R1076 B.n157 B.n156 10.6151
R1077 B.n160 B.n157 10.6151
R1078 B.n165 B.n162 10.6151
R1079 B.n166 B.n165 10.6151
R1080 B.n169 B.n166 10.6151
R1081 B.n170 B.n169 10.6151
R1082 B.n173 B.n170 10.6151
R1083 B.n174 B.n173 10.6151
R1084 B.n177 B.n174 10.6151
R1085 B.n178 B.n177 10.6151
R1086 B.n182 B.n181 10.6151
R1087 B.n185 B.n182 10.6151
R1088 B.n186 B.n185 10.6151
R1089 B.n189 B.n186 10.6151
R1090 B.n190 B.n189 10.6151
R1091 B.n193 B.n190 10.6151
R1092 B.n194 B.n193 10.6151
R1093 B.n197 B.n194 10.6151
R1094 B.n198 B.n197 10.6151
R1095 B.n201 B.n198 10.6151
R1096 B.n202 B.n201 10.6151
R1097 B.n205 B.n202 10.6151
R1098 B.n206 B.n205 10.6151
R1099 B.n209 B.n206 10.6151
R1100 B.n210 B.n209 10.6151
R1101 B.n213 B.n210 10.6151
R1102 B.n214 B.n213 10.6151
R1103 B.n217 B.n214 10.6151
R1104 B.n218 B.n217 10.6151
R1105 B.n221 B.n218 10.6151
R1106 B.n222 B.n221 10.6151
R1107 B.n225 B.n222 10.6151
R1108 B.n226 B.n225 10.6151
R1109 B.n229 B.n226 10.6151
R1110 B.n230 B.n229 10.6151
R1111 B.n624 B.n230 10.6151
R1112 B.n466 B.n465 10.6151
R1113 B.n466 B.n293 10.6151
R1114 B.n476 B.n293 10.6151
R1115 B.n477 B.n476 10.6151
R1116 B.n478 B.n477 10.6151
R1117 B.n478 B.n286 10.6151
R1118 B.n489 B.n286 10.6151
R1119 B.n490 B.n489 10.6151
R1120 B.n491 B.n490 10.6151
R1121 B.n491 B.n278 10.6151
R1122 B.n501 B.n278 10.6151
R1123 B.n502 B.n501 10.6151
R1124 B.n503 B.n502 10.6151
R1125 B.n503 B.n270 10.6151
R1126 B.n513 B.n270 10.6151
R1127 B.n514 B.n513 10.6151
R1128 B.n515 B.n514 10.6151
R1129 B.n515 B.n262 10.6151
R1130 B.n525 B.n262 10.6151
R1131 B.n526 B.n525 10.6151
R1132 B.n527 B.n526 10.6151
R1133 B.n527 B.n254 10.6151
R1134 B.n537 B.n254 10.6151
R1135 B.n538 B.n537 10.6151
R1136 B.n539 B.n538 10.6151
R1137 B.n539 B.n247 10.6151
R1138 B.n550 B.n247 10.6151
R1139 B.n551 B.n550 10.6151
R1140 B.n552 B.n551 10.6151
R1141 B.n552 B.n238 10.6151
R1142 B.n562 B.n238 10.6151
R1143 B.n563 B.n562 10.6151
R1144 B.n565 B.n563 10.6151
R1145 B.n565 B.n564 10.6151
R1146 B.n564 B.n231 10.6151
R1147 B.n576 B.n231 10.6151
R1148 B.n577 B.n576 10.6151
R1149 B.n578 B.n577 10.6151
R1150 B.n579 B.n578 10.6151
R1151 B.n581 B.n579 10.6151
R1152 B.n582 B.n581 10.6151
R1153 B.n583 B.n582 10.6151
R1154 B.n584 B.n583 10.6151
R1155 B.n586 B.n584 10.6151
R1156 B.n587 B.n586 10.6151
R1157 B.n588 B.n587 10.6151
R1158 B.n589 B.n588 10.6151
R1159 B.n591 B.n589 10.6151
R1160 B.n592 B.n591 10.6151
R1161 B.n593 B.n592 10.6151
R1162 B.n594 B.n593 10.6151
R1163 B.n596 B.n594 10.6151
R1164 B.n597 B.n596 10.6151
R1165 B.n598 B.n597 10.6151
R1166 B.n599 B.n598 10.6151
R1167 B.n601 B.n599 10.6151
R1168 B.n602 B.n601 10.6151
R1169 B.n603 B.n602 10.6151
R1170 B.n604 B.n603 10.6151
R1171 B.n606 B.n604 10.6151
R1172 B.n607 B.n606 10.6151
R1173 B.n608 B.n607 10.6151
R1174 B.n609 B.n608 10.6151
R1175 B.n611 B.n609 10.6151
R1176 B.n612 B.n611 10.6151
R1177 B.n613 B.n612 10.6151
R1178 B.n614 B.n613 10.6151
R1179 B.n616 B.n614 10.6151
R1180 B.n617 B.n616 10.6151
R1181 B.n618 B.n617 10.6151
R1182 B.n619 B.n618 10.6151
R1183 B.n621 B.n619 10.6151
R1184 B.n622 B.n621 10.6151
R1185 B.n623 B.n622 10.6151
R1186 B.n458 B.n457 10.6151
R1187 B.n457 B.n456 10.6151
R1188 B.n456 B.n455 10.6151
R1189 B.n455 B.n453 10.6151
R1190 B.n453 B.n450 10.6151
R1191 B.n450 B.n449 10.6151
R1192 B.n449 B.n446 10.6151
R1193 B.n446 B.n445 10.6151
R1194 B.n445 B.n442 10.6151
R1195 B.n442 B.n441 10.6151
R1196 B.n441 B.n438 10.6151
R1197 B.n438 B.n437 10.6151
R1198 B.n437 B.n434 10.6151
R1199 B.n434 B.n433 10.6151
R1200 B.n433 B.n430 10.6151
R1201 B.n430 B.n429 10.6151
R1202 B.n429 B.n426 10.6151
R1203 B.n426 B.n425 10.6151
R1204 B.n425 B.n422 10.6151
R1205 B.n422 B.n421 10.6151
R1206 B.n421 B.n418 10.6151
R1207 B.n418 B.n417 10.6151
R1208 B.n417 B.n414 10.6151
R1209 B.n414 B.n413 10.6151
R1210 B.n413 B.n410 10.6151
R1211 B.n410 B.n409 10.6151
R1212 B.n406 B.n405 10.6151
R1213 B.n405 B.n402 10.6151
R1214 B.n402 B.n401 10.6151
R1215 B.n401 B.n398 10.6151
R1216 B.n398 B.n397 10.6151
R1217 B.n397 B.n394 10.6151
R1218 B.n394 B.n393 10.6151
R1219 B.n393 B.n390 10.6151
R1220 B.n388 B.n385 10.6151
R1221 B.n385 B.n384 10.6151
R1222 B.n384 B.n381 10.6151
R1223 B.n381 B.n380 10.6151
R1224 B.n380 B.n377 10.6151
R1225 B.n377 B.n376 10.6151
R1226 B.n376 B.n373 10.6151
R1227 B.n373 B.n372 10.6151
R1228 B.n372 B.n369 10.6151
R1229 B.n369 B.n368 10.6151
R1230 B.n368 B.n365 10.6151
R1231 B.n365 B.n364 10.6151
R1232 B.n364 B.n361 10.6151
R1233 B.n361 B.n360 10.6151
R1234 B.n360 B.n357 10.6151
R1235 B.n357 B.n356 10.6151
R1236 B.n356 B.n353 10.6151
R1237 B.n353 B.n352 10.6151
R1238 B.n352 B.n349 10.6151
R1239 B.n349 B.n348 10.6151
R1240 B.n348 B.n345 10.6151
R1241 B.n345 B.n344 10.6151
R1242 B.n344 B.n341 10.6151
R1243 B.n341 B.n340 10.6151
R1244 B.n340 B.n301 10.6151
R1245 B.n464 B.n301 10.6151
R1246 B.n470 B.n297 10.6151
R1247 B.n471 B.n470 10.6151
R1248 B.n472 B.n471 10.6151
R1249 B.n472 B.n289 10.6151
R1250 B.n483 B.n289 10.6151
R1251 B.n484 B.n483 10.6151
R1252 B.n485 B.n484 10.6151
R1253 B.n485 B.n282 10.6151
R1254 B.n495 B.n282 10.6151
R1255 B.n496 B.n495 10.6151
R1256 B.n497 B.n496 10.6151
R1257 B.n497 B.n274 10.6151
R1258 B.n507 B.n274 10.6151
R1259 B.n508 B.n507 10.6151
R1260 B.n509 B.n508 10.6151
R1261 B.n509 B.n266 10.6151
R1262 B.n519 B.n266 10.6151
R1263 B.n520 B.n519 10.6151
R1264 B.n521 B.n520 10.6151
R1265 B.n521 B.n258 10.6151
R1266 B.n531 B.n258 10.6151
R1267 B.n532 B.n531 10.6151
R1268 B.n533 B.n532 10.6151
R1269 B.n533 B.n250 10.6151
R1270 B.n544 B.n250 10.6151
R1271 B.n545 B.n544 10.6151
R1272 B.n546 B.n545 10.6151
R1273 B.n546 B.n243 10.6151
R1274 B.n556 B.n243 10.6151
R1275 B.n557 B.n556 10.6151
R1276 B.n558 B.n557 10.6151
R1277 B.n558 B.n235 10.6151
R1278 B.n569 B.n235 10.6151
R1279 B.n570 B.n569 10.6151
R1280 B.n571 B.n570 10.6151
R1281 B.n571 B.n0 10.6151
R1282 B.n696 B.n1 10.6151
R1283 B.n696 B.n695 10.6151
R1284 B.n695 B.n694 10.6151
R1285 B.n694 B.n10 10.6151
R1286 B.n688 B.n10 10.6151
R1287 B.n688 B.n687 10.6151
R1288 B.n687 B.n686 10.6151
R1289 B.n686 B.n17 10.6151
R1290 B.n680 B.n17 10.6151
R1291 B.n680 B.n679 10.6151
R1292 B.n679 B.n678 10.6151
R1293 B.n678 B.n23 10.6151
R1294 B.n672 B.n23 10.6151
R1295 B.n672 B.n671 10.6151
R1296 B.n671 B.n670 10.6151
R1297 B.n670 B.n31 10.6151
R1298 B.n664 B.n31 10.6151
R1299 B.n664 B.n663 10.6151
R1300 B.n663 B.n662 10.6151
R1301 B.n662 B.n38 10.6151
R1302 B.n656 B.n38 10.6151
R1303 B.n656 B.n655 10.6151
R1304 B.n655 B.n654 10.6151
R1305 B.n654 B.n45 10.6151
R1306 B.n648 B.n45 10.6151
R1307 B.n648 B.n647 10.6151
R1308 B.n647 B.n646 10.6151
R1309 B.n646 B.n52 10.6151
R1310 B.n640 B.n52 10.6151
R1311 B.n640 B.n639 10.6151
R1312 B.n639 B.n638 10.6151
R1313 B.n638 B.n58 10.6151
R1314 B.n632 B.n58 10.6151
R1315 B.n632 B.n631 10.6151
R1316 B.n631 B.n630 10.6151
R1317 B.n630 B.n66 10.6151
R1318 B.n162 B.n161 6.5566
R1319 B.n178 B.n104 6.5566
R1320 B.n406 B.n336 6.5566
R1321 B.n390 B.n389 6.5566
R1322 B.n161 B.n160 4.05904
R1323 B.n181 B.n104 4.05904
R1324 B.n409 B.n336 4.05904
R1325 B.n389 B.n388 4.05904
R1326 B.n529 B.t5 3.60558
R1327 B.n668 B.t1 3.60558
R1328 B.n702 B.n0 2.81026
R1329 B.n702 B.n1 2.81026
R1330 VP.n28 VP.n27 177.204
R1331 VP.n50 VP.n49 177.204
R1332 VP.n26 VP.n25 177.204
R1333 VP.n13 VP.n12 161.3
R1334 VP.n14 VP.n9 161.3
R1335 VP.n16 VP.n15 161.3
R1336 VP.n17 VP.n8 161.3
R1337 VP.n20 VP.n19 161.3
R1338 VP.n21 VP.n7 161.3
R1339 VP.n23 VP.n22 161.3
R1340 VP.n24 VP.n6 161.3
R1341 VP.n48 VP.n0 161.3
R1342 VP.n47 VP.n46 161.3
R1343 VP.n45 VP.n1 161.3
R1344 VP.n44 VP.n43 161.3
R1345 VP.n41 VP.n2 161.3
R1346 VP.n40 VP.n39 161.3
R1347 VP.n38 VP.n3 161.3
R1348 VP.n37 VP.n36 161.3
R1349 VP.n34 VP.n4 161.3
R1350 VP.n33 VP.n32 161.3
R1351 VP.n31 VP.n5 161.3
R1352 VP.n30 VP.n29 161.3
R1353 VP.n10 VP.t3 136.07
R1354 VP.n28 VP.t0 103.094
R1355 VP.n35 VP.t1 103.094
R1356 VP.n42 VP.t2 103.094
R1357 VP.n49 VP.t5 103.094
R1358 VP.n25 VP.t7 103.094
R1359 VP.n18 VP.t4 103.094
R1360 VP.n11 VP.t6 103.094
R1361 VP.n33 VP.n5 56.5193
R1362 VP.n40 VP.n3 56.5193
R1363 VP.n47 VP.n1 56.5193
R1364 VP.n23 VP.n7 56.5193
R1365 VP.n16 VP.n9 56.5193
R1366 VP.n11 VP.n10 55.22
R1367 VP.n27 VP.n26 42.402
R1368 VP.n29 VP.n5 24.4675
R1369 VP.n34 VP.n33 24.4675
R1370 VP.n36 VP.n3 24.4675
R1371 VP.n41 VP.n40 24.4675
R1372 VP.n43 VP.n1 24.4675
R1373 VP.n48 VP.n47 24.4675
R1374 VP.n24 VP.n23 24.4675
R1375 VP.n17 VP.n16 24.4675
R1376 VP.n19 VP.n7 24.4675
R1377 VP.n12 VP.n9 24.4675
R1378 VP.n13 VP.n10 17.9267
R1379 VP.n35 VP.n34 13.4574
R1380 VP.n43 VP.n42 13.4574
R1381 VP.n19 VP.n18 13.4574
R1382 VP.n36 VP.n35 11.0107
R1383 VP.n42 VP.n41 11.0107
R1384 VP.n18 VP.n17 11.0107
R1385 VP.n12 VP.n11 11.0107
R1386 VP.n29 VP.n28 8.56395
R1387 VP.n49 VP.n48 8.56395
R1388 VP.n25 VP.n24 8.56395
R1389 VP.n14 VP.n13 0.189894
R1390 VP.n15 VP.n14 0.189894
R1391 VP.n15 VP.n8 0.189894
R1392 VP.n20 VP.n8 0.189894
R1393 VP.n21 VP.n20 0.189894
R1394 VP.n22 VP.n21 0.189894
R1395 VP.n22 VP.n6 0.189894
R1396 VP.n26 VP.n6 0.189894
R1397 VP.n30 VP.n27 0.189894
R1398 VP.n31 VP.n30 0.189894
R1399 VP.n32 VP.n31 0.189894
R1400 VP.n32 VP.n4 0.189894
R1401 VP.n37 VP.n4 0.189894
R1402 VP.n38 VP.n37 0.189894
R1403 VP.n39 VP.n38 0.189894
R1404 VP.n39 VP.n2 0.189894
R1405 VP.n44 VP.n2 0.189894
R1406 VP.n45 VP.n44 0.189894
R1407 VP.n46 VP.n45 0.189894
R1408 VP.n46 VP.n0 0.189894
R1409 VP.n50 VP.n0 0.189894
R1410 VP VP.n50 0.0516364
R1411 VDD1 VDD1.n0 69.9914
R1412 VDD1.n3 VDD1.n2 69.8767
R1413 VDD1.n3 VDD1.n1 69.8767
R1414 VDD1.n5 VDD1.n4 69.0925
R1415 VDD1.n5 VDD1.n3 37.8371
R1416 VDD1.n4 VDD1.t3 2.85764
R1417 VDD1.n4 VDD1.t0 2.85764
R1418 VDD1.n0 VDD1.t4 2.85764
R1419 VDD1.n0 VDD1.t1 2.85764
R1420 VDD1.n2 VDD1.t5 2.85764
R1421 VDD1.n2 VDD1.t2 2.85764
R1422 VDD1.n1 VDD1.t7 2.85764
R1423 VDD1.n1 VDD1.t6 2.85764
R1424 VDD1 VDD1.n5 0.782828
C0 VTAIL VP 5.05869f
C1 VDD2 VP 0.415461f
C2 VDD1 VP 4.90875f
C3 VTAIL VN 5.04459f
C4 VDD2 VN 4.64422f
C5 VTAIL VDD2 6.14761f
C6 VDD1 VN 0.150029f
C7 VTAIL VDD1 6.09977f
C8 VDD2 VDD1 1.26816f
C9 VP VN 5.523951f
C10 VDD2 B 4.003497f
C11 VDD1 B 4.341407f
C12 VTAIL B 6.529171f
C13 VN B 11.21228f
C14 VP B 9.757092f
C15 VDD1.t4 B 0.136858f
C16 VDD1.t1 B 0.136858f
C17 VDD1.n0 B 1.17621f
C18 VDD1.t7 B 0.136858f
C19 VDD1.t6 B 0.136858f
C20 VDD1.n1 B 1.17545f
C21 VDD1.t5 B 0.136858f
C22 VDD1.t2 B 0.136858f
C23 VDD1.n2 B 1.17545f
C24 VDD1.n3 B 2.43102f
C25 VDD1.t3 B 0.136858f
C26 VDD1.t0 B 0.136858f
C27 VDD1.n4 B 1.1709f
C28 VDD1.n5 B 2.23334f
C29 VP.n0 B 0.03192f
C30 VP.t5 B 0.955977f
C31 VP.n1 B 0.04215f
C32 VP.n2 B 0.03192f
C33 VP.t2 B 0.955977f
C34 VP.n3 B 0.046598f
C35 VP.n4 B 0.03192f
C36 VP.t1 B 0.955977f
C37 VP.n5 B 0.051045f
C38 VP.n6 B 0.03192f
C39 VP.t7 B 0.955977f
C40 VP.n7 B 0.04215f
C41 VP.n8 B 0.03192f
C42 VP.t4 B 0.955977f
C43 VP.n9 B 0.046598f
C44 VP.t3 B 1.07614f
C45 VP.n10 B 0.435939f
C46 VP.t6 B 0.955977f
C47 VP.n11 B 0.425423f
C48 VP.n12 B 0.043336f
C49 VP.n13 B 0.204196f
C50 VP.n14 B 0.03192f
C51 VP.n15 B 0.03192f
C52 VP.n16 B 0.046598f
C53 VP.n17 B 0.043336f
C54 VP.n18 B 0.364129f
C55 VP.n19 B 0.046273f
C56 VP.n20 B 0.03192f
C57 VP.n21 B 0.03192f
C58 VP.n22 B 0.03192f
C59 VP.n23 B 0.051045f
C60 VP.n24 B 0.040399f
C61 VP.n25 B 0.434054f
C62 VP.n26 B 1.34548f
C63 VP.n27 B 1.37254f
C64 VP.t0 B 0.955977f
C65 VP.n28 B 0.434054f
C66 VP.n29 B 0.040399f
C67 VP.n30 B 0.03192f
C68 VP.n31 B 0.03192f
C69 VP.n32 B 0.03192f
C70 VP.n33 B 0.04215f
C71 VP.n34 B 0.046273f
C72 VP.n35 B 0.364129f
C73 VP.n36 B 0.043336f
C74 VP.n37 B 0.03192f
C75 VP.n38 B 0.03192f
C76 VP.n39 B 0.03192f
C77 VP.n40 B 0.046598f
C78 VP.n41 B 0.043336f
C79 VP.n42 B 0.364129f
C80 VP.n43 B 0.046273f
C81 VP.n44 B 0.03192f
C82 VP.n45 B 0.03192f
C83 VP.n46 B 0.03192f
C84 VP.n47 B 0.051045f
C85 VP.n48 B 0.040399f
C86 VP.n49 B 0.434054f
C87 VP.n50 B 0.031631f
C88 VDD2.t6 B 0.134252f
C89 VDD2.t7 B 0.134252f
C90 VDD2.n0 B 1.15306f
C91 VDD2.t0 B 0.134252f
C92 VDD2.t2 B 0.134252f
C93 VDD2.n1 B 1.15306f
C94 VDD2.n2 B 2.3329f
C95 VDD2.t1 B 0.134252f
C96 VDD2.t3 B 0.134252f
C97 VDD2.n3 B 1.14861f
C98 VDD2.n4 B 2.16129f
C99 VDD2.t4 B 0.134252f
C100 VDD2.t5 B 0.134252f
C101 VDD2.n5 B 1.15303f
C102 VTAIL.t15 B 0.116469f
C103 VTAIL.t9 B 0.116469f
C104 VTAIL.n0 B 0.944964f
C105 VTAIL.n1 B 0.30765f
C106 VTAIL.t10 B 1.20335f
C107 VTAIL.n2 B 0.395111f
C108 VTAIL.t2 B 1.20335f
C109 VTAIL.n3 B 0.395111f
C110 VTAIL.t5 B 0.116469f
C111 VTAIL.t7 B 0.116469f
C112 VTAIL.n4 B 0.944964f
C113 VTAIL.n5 B 0.418862f
C114 VTAIL.t3 B 1.20335f
C115 VTAIL.n6 B 1.17642f
C116 VTAIL.t14 B 1.20336f
C117 VTAIL.n7 B 1.17641f
C118 VTAIL.t13 B 0.116469f
C119 VTAIL.t12 B 0.116469f
C120 VTAIL.n8 B 0.944971f
C121 VTAIL.n9 B 0.418856f
C122 VTAIL.t8 B 1.20336f
C123 VTAIL.n10 B 0.395101f
C124 VTAIL.t0 B 1.20336f
C125 VTAIL.n11 B 0.395101f
C126 VTAIL.t4 B 0.116469f
C127 VTAIL.t1 B 0.116469f
C128 VTAIL.n12 B 0.944971f
C129 VTAIL.n13 B 0.418856f
C130 VTAIL.t6 B 1.20335f
C131 VTAIL.n14 B 1.17642f
C132 VTAIL.t11 B 1.20335f
C133 VTAIL.n15 B 1.17243f
C134 VN.n0 B 0.031007f
C135 VN.t5 B 0.928619f
C136 VN.n1 B 0.040944f
C137 VN.n2 B 0.031007f
C138 VN.t7 B 0.928619f
C139 VN.n3 B 0.045264f
C140 VN.t1 B 1.04534f
C141 VN.n4 B 0.423463f
C142 VN.t0 B 0.928619f
C143 VN.n5 B 0.413248f
C144 VN.n6 B 0.042096f
C145 VN.n7 B 0.198353f
C146 VN.n8 B 0.031007f
C147 VN.n9 B 0.031007f
C148 VN.n10 B 0.045264f
C149 VN.n11 B 0.042096f
C150 VN.n12 B 0.353709f
C151 VN.n13 B 0.044949f
C152 VN.n14 B 0.031007f
C153 VN.n15 B 0.031007f
C154 VN.n16 B 0.031007f
C155 VN.n17 B 0.049585f
C156 VN.n18 B 0.039242f
C157 VN.n19 B 0.421632f
C158 VN.n20 B 0.030726f
C159 VN.n21 B 0.031007f
C160 VN.t6 B 0.928619f
C161 VN.n22 B 0.040944f
C162 VN.n23 B 0.031007f
C163 VN.t4 B 0.928619f
C164 VN.n24 B 0.045264f
C165 VN.t2 B 1.04534f
C166 VN.n25 B 0.423463f
C167 VN.t3 B 0.928619f
C168 VN.n26 B 0.413248f
C169 VN.n27 B 0.042096f
C170 VN.n28 B 0.198353f
C171 VN.n29 B 0.031007f
C172 VN.n30 B 0.031007f
C173 VN.n31 B 0.045264f
C174 VN.n32 B 0.042096f
C175 VN.n33 B 0.353709f
C176 VN.n34 B 0.044949f
C177 VN.n35 B 0.031007f
C178 VN.n36 B 0.031007f
C179 VN.n37 B 0.031007f
C180 VN.n38 B 0.049585f
C181 VN.n39 B 0.039242f
C182 VN.n40 B 0.421632f
C183 VN.n41 B 1.32732f
.ends

