* NGSPICE file created from diff_pair_sample_1409.ext - technology: sky130A

.subckt diff_pair_sample_1409 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=0 ps=0 w=11.06 l=2.92
X1 B.t8 B.t6 B.t7 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=0 ps=0 w=11.06 l=2.92
X2 B.t5 B.t3 B.t4 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=0 ps=0 w=11.06 l=2.92
X3 VTAIL.t7 VN.t0 VDD2.t2 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=1.8249 ps=11.39 w=11.06 l=2.92
X4 VDD2.t1 VN.t1 VTAIL.t6 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=1.8249 pd=11.39 as=4.3134 ps=22.9 w=11.06 l=2.92
X5 VDD1.t3 VP.t0 VTAIL.t3 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=1.8249 pd=11.39 as=4.3134 ps=22.9 w=11.06 l=2.92
X6 VTAIL.t5 VN.t2 VDD2.t3 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=1.8249 ps=11.39 w=11.06 l=2.92
X7 VDD1.t2 VP.t1 VTAIL.t2 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=1.8249 pd=11.39 as=4.3134 ps=22.9 w=11.06 l=2.92
X8 VDD2.t0 VN.t3 VTAIL.t4 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=1.8249 pd=11.39 as=4.3134 ps=22.9 w=11.06 l=2.92
X9 VTAIL.t1 VP.t2 VDD1.t1 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=1.8249 ps=11.39 w=11.06 l=2.92
X10 VTAIL.t0 VP.t3 VDD1.t0 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=1.8249 ps=11.39 w=11.06 l=2.92
X11 B.t2 B.t0 B.t1 w_n2920_n3180# sky130_fd_pr__pfet_01v8 ad=4.3134 pd=22.9 as=0 ps=0 w=11.06 l=2.92
R0 B.n471 B.n68 585
R1 B.n473 B.n472 585
R2 B.n474 B.n67 585
R3 B.n476 B.n475 585
R4 B.n477 B.n66 585
R5 B.n479 B.n478 585
R6 B.n480 B.n65 585
R7 B.n482 B.n481 585
R8 B.n483 B.n64 585
R9 B.n485 B.n484 585
R10 B.n486 B.n63 585
R11 B.n488 B.n487 585
R12 B.n489 B.n62 585
R13 B.n491 B.n490 585
R14 B.n492 B.n61 585
R15 B.n494 B.n493 585
R16 B.n495 B.n60 585
R17 B.n497 B.n496 585
R18 B.n498 B.n59 585
R19 B.n500 B.n499 585
R20 B.n501 B.n58 585
R21 B.n503 B.n502 585
R22 B.n504 B.n57 585
R23 B.n506 B.n505 585
R24 B.n507 B.n56 585
R25 B.n509 B.n508 585
R26 B.n510 B.n55 585
R27 B.n512 B.n511 585
R28 B.n513 B.n54 585
R29 B.n515 B.n514 585
R30 B.n516 B.n53 585
R31 B.n518 B.n517 585
R32 B.n519 B.n52 585
R33 B.n521 B.n520 585
R34 B.n522 B.n51 585
R35 B.n524 B.n523 585
R36 B.n525 B.n50 585
R37 B.n527 B.n526 585
R38 B.n528 B.n47 585
R39 B.n531 B.n530 585
R40 B.n532 B.n46 585
R41 B.n534 B.n533 585
R42 B.n535 B.n45 585
R43 B.n537 B.n536 585
R44 B.n538 B.n44 585
R45 B.n540 B.n539 585
R46 B.n541 B.n43 585
R47 B.n543 B.n542 585
R48 B.n545 B.n544 585
R49 B.n546 B.n39 585
R50 B.n548 B.n547 585
R51 B.n549 B.n38 585
R52 B.n551 B.n550 585
R53 B.n552 B.n37 585
R54 B.n554 B.n553 585
R55 B.n555 B.n36 585
R56 B.n557 B.n556 585
R57 B.n558 B.n35 585
R58 B.n560 B.n559 585
R59 B.n561 B.n34 585
R60 B.n563 B.n562 585
R61 B.n564 B.n33 585
R62 B.n566 B.n565 585
R63 B.n567 B.n32 585
R64 B.n569 B.n568 585
R65 B.n570 B.n31 585
R66 B.n572 B.n571 585
R67 B.n573 B.n30 585
R68 B.n575 B.n574 585
R69 B.n576 B.n29 585
R70 B.n578 B.n577 585
R71 B.n579 B.n28 585
R72 B.n581 B.n580 585
R73 B.n582 B.n27 585
R74 B.n584 B.n583 585
R75 B.n585 B.n26 585
R76 B.n587 B.n586 585
R77 B.n588 B.n25 585
R78 B.n590 B.n589 585
R79 B.n591 B.n24 585
R80 B.n593 B.n592 585
R81 B.n594 B.n23 585
R82 B.n596 B.n595 585
R83 B.n597 B.n22 585
R84 B.n599 B.n598 585
R85 B.n600 B.n21 585
R86 B.n602 B.n601 585
R87 B.n470 B.n469 585
R88 B.n468 B.n69 585
R89 B.n467 B.n466 585
R90 B.n465 B.n70 585
R91 B.n464 B.n463 585
R92 B.n462 B.n71 585
R93 B.n461 B.n460 585
R94 B.n459 B.n72 585
R95 B.n458 B.n457 585
R96 B.n456 B.n73 585
R97 B.n455 B.n454 585
R98 B.n453 B.n74 585
R99 B.n452 B.n451 585
R100 B.n450 B.n75 585
R101 B.n449 B.n448 585
R102 B.n447 B.n76 585
R103 B.n446 B.n445 585
R104 B.n444 B.n77 585
R105 B.n443 B.n442 585
R106 B.n441 B.n78 585
R107 B.n440 B.n439 585
R108 B.n438 B.n79 585
R109 B.n437 B.n436 585
R110 B.n435 B.n80 585
R111 B.n434 B.n433 585
R112 B.n432 B.n81 585
R113 B.n431 B.n430 585
R114 B.n429 B.n82 585
R115 B.n428 B.n427 585
R116 B.n426 B.n83 585
R117 B.n425 B.n424 585
R118 B.n423 B.n84 585
R119 B.n422 B.n421 585
R120 B.n420 B.n85 585
R121 B.n419 B.n418 585
R122 B.n417 B.n86 585
R123 B.n416 B.n415 585
R124 B.n414 B.n87 585
R125 B.n413 B.n412 585
R126 B.n411 B.n88 585
R127 B.n410 B.n409 585
R128 B.n408 B.n89 585
R129 B.n407 B.n406 585
R130 B.n405 B.n90 585
R131 B.n404 B.n403 585
R132 B.n402 B.n91 585
R133 B.n401 B.n400 585
R134 B.n399 B.n92 585
R135 B.n398 B.n397 585
R136 B.n396 B.n93 585
R137 B.n395 B.n394 585
R138 B.n393 B.n94 585
R139 B.n392 B.n391 585
R140 B.n390 B.n95 585
R141 B.n389 B.n388 585
R142 B.n387 B.n96 585
R143 B.n386 B.n385 585
R144 B.n384 B.n97 585
R145 B.n383 B.n382 585
R146 B.n381 B.n98 585
R147 B.n380 B.n379 585
R148 B.n378 B.n99 585
R149 B.n377 B.n376 585
R150 B.n375 B.n100 585
R151 B.n374 B.n373 585
R152 B.n372 B.n101 585
R153 B.n371 B.n370 585
R154 B.n369 B.n102 585
R155 B.n368 B.n367 585
R156 B.n366 B.n103 585
R157 B.n365 B.n364 585
R158 B.n363 B.n104 585
R159 B.n362 B.n361 585
R160 B.n360 B.n105 585
R161 B.n359 B.n358 585
R162 B.n227 B.n226 585
R163 B.n228 B.n153 585
R164 B.n230 B.n229 585
R165 B.n231 B.n152 585
R166 B.n233 B.n232 585
R167 B.n234 B.n151 585
R168 B.n236 B.n235 585
R169 B.n237 B.n150 585
R170 B.n239 B.n238 585
R171 B.n240 B.n149 585
R172 B.n242 B.n241 585
R173 B.n243 B.n148 585
R174 B.n245 B.n244 585
R175 B.n246 B.n147 585
R176 B.n248 B.n247 585
R177 B.n249 B.n146 585
R178 B.n251 B.n250 585
R179 B.n252 B.n145 585
R180 B.n254 B.n253 585
R181 B.n255 B.n144 585
R182 B.n257 B.n256 585
R183 B.n258 B.n143 585
R184 B.n260 B.n259 585
R185 B.n261 B.n142 585
R186 B.n263 B.n262 585
R187 B.n264 B.n141 585
R188 B.n266 B.n265 585
R189 B.n267 B.n140 585
R190 B.n269 B.n268 585
R191 B.n270 B.n139 585
R192 B.n272 B.n271 585
R193 B.n273 B.n138 585
R194 B.n275 B.n274 585
R195 B.n276 B.n137 585
R196 B.n278 B.n277 585
R197 B.n279 B.n136 585
R198 B.n281 B.n280 585
R199 B.n282 B.n135 585
R200 B.n284 B.n283 585
R201 B.n286 B.n285 585
R202 B.n287 B.n131 585
R203 B.n289 B.n288 585
R204 B.n290 B.n130 585
R205 B.n292 B.n291 585
R206 B.n293 B.n129 585
R207 B.n295 B.n294 585
R208 B.n296 B.n128 585
R209 B.n298 B.n297 585
R210 B.n300 B.n125 585
R211 B.n302 B.n301 585
R212 B.n303 B.n124 585
R213 B.n305 B.n304 585
R214 B.n306 B.n123 585
R215 B.n308 B.n307 585
R216 B.n309 B.n122 585
R217 B.n311 B.n310 585
R218 B.n312 B.n121 585
R219 B.n314 B.n313 585
R220 B.n315 B.n120 585
R221 B.n317 B.n316 585
R222 B.n318 B.n119 585
R223 B.n320 B.n319 585
R224 B.n321 B.n118 585
R225 B.n323 B.n322 585
R226 B.n324 B.n117 585
R227 B.n326 B.n325 585
R228 B.n327 B.n116 585
R229 B.n329 B.n328 585
R230 B.n330 B.n115 585
R231 B.n332 B.n331 585
R232 B.n333 B.n114 585
R233 B.n335 B.n334 585
R234 B.n336 B.n113 585
R235 B.n338 B.n337 585
R236 B.n339 B.n112 585
R237 B.n341 B.n340 585
R238 B.n342 B.n111 585
R239 B.n344 B.n343 585
R240 B.n345 B.n110 585
R241 B.n347 B.n346 585
R242 B.n348 B.n109 585
R243 B.n350 B.n349 585
R244 B.n351 B.n108 585
R245 B.n353 B.n352 585
R246 B.n354 B.n107 585
R247 B.n356 B.n355 585
R248 B.n357 B.n106 585
R249 B.n225 B.n154 585
R250 B.n224 B.n223 585
R251 B.n222 B.n155 585
R252 B.n221 B.n220 585
R253 B.n219 B.n156 585
R254 B.n218 B.n217 585
R255 B.n216 B.n157 585
R256 B.n215 B.n214 585
R257 B.n213 B.n158 585
R258 B.n212 B.n211 585
R259 B.n210 B.n159 585
R260 B.n209 B.n208 585
R261 B.n207 B.n160 585
R262 B.n206 B.n205 585
R263 B.n204 B.n161 585
R264 B.n203 B.n202 585
R265 B.n201 B.n162 585
R266 B.n200 B.n199 585
R267 B.n198 B.n163 585
R268 B.n197 B.n196 585
R269 B.n195 B.n164 585
R270 B.n194 B.n193 585
R271 B.n192 B.n165 585
R272 B.n191 B.n190 585
R273 B.n189 B.n166 585
R274 B.n188 B.n187 585
R275 B.n186 B.n167 585
R276 B.n185 B.n184 585
R277 B.n183 B.n168 585
R278 B.n182 B.n181 585
R279 B.n180 B.n169 585
R280 B.n179 B.n178 585
R281 B.n177 B.n170 585
R282 B.n176 B.n175 585
R283 B.n174 B.n171 585
R284 B.n173 B.n172 585
R285 B.n2 B.n0 585
R286 B.n657 B.n1 585
R287 B.n656 B.n655 585
R288 B.n654 B.n3 585
R289 B.n653 B.n652 585
R290 B.n651 B.n4 585
R291 B.n650 B.n649 585
R292 B.n648 B.n5 585
R293 B.n647 B.n646 585
R294 B.n645 B.n6 585
R295 B.n644 B.n643 585
R296 B.n642 B.n7 585
R297 B.n641 B.n640 585
R298 B.n639 B.n8 585
R299 B.n638 B.n637 585
R300 B.n636 B.n9 585
R301 B.n635 B.n634 585
R302 B.n633 B.n10 585
R303 B.n632 B.n631 585
R304 B.n630 B.n11 585
R305 B.n629 B.n628 585
R306 B.n627 B.n12 585
R307 B.n626 B.n625 585
R308 B.n624 B.n13 585
R309 B.n623 B.n622 585
R310 B.n621 B.n14 585
R311 B.n620 B.n619 585
R312 B.n618 B.n15 585
R313 B.n617 B.n616 585
R314 B.n615 B.n16 585
R315 B.n614 B.n613 585
R316 B.n612 B.n17 585
R317 B.n611 B.n610 585
R318 B.n609 B.n18 585
R319 B.n608 B.n607 585
R320 B.n606 B.n19 585
R321 B.n605 B.n604 585
R322 B.n603 B.n20 585
R323 B.n659 B.n658 585
R324 B.n226 B.n225 487.695
R325 B.n603 B.n602 487.695
R326 B.n358 B.n357 487.695
R327 B.n471 B.n470 487.695
R328 B.n126 B.t0 299.767
R329 B.n132 B.t3 299.767
R330 B.n40 B.t9 299.767
R331 B.n48 B.t6 299.767
R332 B.n126 B.t2 173.864
R333 B.n48 B.t7 173.864
R334 B.n132 B.t5 173.851
R335 B.n40 B.t10 173.851
R336 B.n225 B.n224 163.367
R337 B.n224 B.n155 163.367
R338 B.n220 B.n155 163.367
R339 B.n220 B.n219 163.367
R340 B.n219 B.n218 163.367
R341 B.n218 B.n157 163.367
R342 B.n214 B.n157 163.367
R343 B.n214 B.n213 163.367
R344 B.n213 B.n212 163.367
R345 B.n212 B.n159 163.367
R346 B.n208 B.n159 163.367
R347 B.n208 B.n207 163.367
R348 B.n207 B.n206 163.367
R349 B.n206 B.n161 163.367
R350 B.n202 B.n161 163.367
R351 B.n202 B.n201 163.367
R352 B.n201 B.n200 163.367
R353 B.n200 B.n163 163.367
R354 B.n196 B.n163 163.367
R355 B.n196 B.n195 163.367
R356 B.n195 B.n194 163.367
R357 B.n194 B.n165 163.367
R358 B.n190 B.n165 163.367
R359 B.n190 B.n189 163.367
R360 B.n189 B.n188 163.367
R361 B.n188 B.n167 163.367
R362 B.n184 B.n167 163.367
R363 B.n184 B.n183 163.367
R364 B.n183 B.n182 163.367
R365 B.n182 B.n169 163.367
R366 B.n178 B.n169 163.367
R367 B.n178 B.n177 163.367
R368 B.n177 B.n176 163.367
R369 B.n176 B.n171 163.367
R370 B.n172 B.n171 163.367
R371 B.n172 B.n2 163.367
R372 B.n658 B.n2 163.367
R373 B.n658 B.n657 163.367
R374 B.n657 B.n656 163.367
R375 B.n656 B.n3 163.367
R376 B.n652 B.n3 163.367
R377 B.n652 B.n651 163.367
R378 B.n651 B.n650 163.367
R379 B.n650 B.n5 163.367
R380 B.n646 B.n5 163.367
R381 B.n646 B.n645 163.367
R382 B.n645 B.n644 163.367
R383 B.n644 B.n7 163.367
R384 B.n640 B.n7 163.367
R385 B.n640 B.n639 163.367
R386 B.n639 B.n638 163.367
R387 B.n638 B.n9 163.367
R388 B.n634 B.n9 163.367
R389 B.n634 B.n633 163.367
R390 B.n633 B.n632 163.367
R391 B.n632 B.n11 163.367
R392 B.n628 B.n11 163.367
R393 B.n628 B.n627 163.367
R394 B.n627 B.n626 163.367
R395 B.n626 B.n13 163.367
R396 B.n622 B.n13 163.367
R397 B.n622 B.n621 163.367
R398 B.n621 B.n620 163.367
R399 B.n620 B.n15 163.367
R400 B.n616 B.n15 163.367
R401 B.n616 B.n615 163.367
R402 B.n615 B.n614 163.367
R403 B.n614 B.n17 163.367
R404 B.n610 B.n17 163.367
R405 B.n610 B.n609 163.367
R406 B.n609 B.n608 163.367
R407 B.n608 B.n19 163.367
R408 B.n604 B.n19 163.367
R409 B.n604 B.n603 163.367
R410 B.n226 B.n153 163.367
R411 B.n230 B.n153 163.367
R412 B.n231 B.n230 163.367
R413 B.n232 B.n231 163.367
R414 B.n232 B.n151 163.367
R415 B.n236 B.n151 163.367
R416 B.n237 B.n236 163.367
R417 B.n238 B.n237 163.367
R418 B.n238 B.n149 163.367
R419 B.n242 B.n149 163.367
R420 B.n243 B.n242 163.367
R421 B.n244 B.n243 163.367
R422 B.n244 B.n147 163.367
R423 B.n248 B.n147 163.367
R424 B.n249 B.n248 163.367
R425 B.n250 B.n249 163.367
R426 B.n250 B.n145 163.367
R427 B.n254 B.n145 163.367
R428 B.n255 B.n254 163.367
R429 B.n256 B.n255 163.367
R430 B.n256 B.n143 163.367
R431 B.n260 B.n143 163.367
R432 B.n261 B.n260 163.367
R433 B.n262 B.n261 163.367
R434 B.n262 B.n141 163.367
R435 B.n266 B.n141 163.367
R436 B.n267 B.n266 163.367
R437 B.n268 B.n267 163.367
R438 B.n268 B.n139 163.367
R439 B.n272 B.n139 163.367
R440 B.n273 B.n272 163.367
R441 B.n274 B.n273 163.367
R442 B.n274 B.n137 163.367
R443 B.n278 B.n137 163.367
R444 B.n279 B.n278 163.367
R445 B.n280 B.n279 163.367
R446 B.n280 B.n135 163.367
R447 B.n284 B.n135 163.367
R448 B.n285 B.n284 163.367
R449 B.n285 B.n131 163.367
R450 B.n289 B.n131 163.367
R451 B.n290 B.n289 163.367
R452 B.n291 B.n290 163.367
R453 B.n291 B.n129 163.367
R454 B.n295 B.n129 163.367
R455 B.n296 B.n295 163.367
R456 B.n297 B.n296 163.367
R457 B.n297 B.n125 163.367
R458 B.n302 B.n125 163.367
R459 B.n303 B.n302 163.367
R460 B.n304 B.n303 163.367
R461 B.n304 B.n123 163.367
R462 B.n308 B.n123 163.367
R463 B.n309 B.n308 163.367
R464 B.n310 B.n309 163.367
R465 B.n310 B.n121 163.367
R466 B.n314 B.n121 163.367
R467 B.n315 B.n314 163.367
R468 B.n316 B.n315 163.367
R469 B.n316 B.n119 163.367
R470 B.n320 B.n119 163.367
R471 B.n321 B.n320 163.367
R472 B.n322 B.n321 163.367
R473 B.n322 B.n117 163.367
R474 B.n326 B.n117 163.367
R475 B.n327 B.n326 163.367
R476 B.n328 B.n327 163.367
R477 B.n328 B.n115 163.367
R478 B.n332 B.n115 163.367
R479 B.n333 B.n332 163.367
R480 B.n334 B.n333 163.367
R481 B.n334 B.n113 163.367
R482 B.n338 B.n113 163.367
R483 B.n339 B.n338 163.367
R484 B.n340 B.n339 163.367
R485 B.n340 B.n111 163.367
R486 B.n344 B.n111 163.367
R487 B.n345 B.n344 163.367
R488 B.n346 B.n345 163.367
R489 B.n346 B.n109 163.367
R490 B.n350 B.n109 163.367
R491 B.n351 B.n350 163.367
R492 B.n352 B.n351 163.367
R493 B.n352 B.n107 163.367
R494 B.n356 B.n107 163.367
R495 B.n357 B.n356 163.367
R496 B.n358 B.n105 163.367
R497 B.n362 B.n105 163.367
R498 B.n363 B.n362 163.367
R499 B.n364 B.n363 163.367
R500 B.n364 B.n103 163.367
R501 B.n368 B.n103 163.367
R502 B.n369 B.n368 163.367
R503 B.n370 B.n369 163.367
R504 B.n370 B.n101 163.367
R505 B.n374 B.n101 163.367
R506 B.n375 B.n374 163.367
R507 B.n376 B.n375 163.367
R508 B.n376 B.n99 163.367
R509 B.n380 B.n99 163.367
R510 B.n381 B.n380 163.367
R511 B.n382 B.n381 163.367
R512 B.n382 B.n97 163.367
R513 B.n386 B.n97 163.367
R514 B.n387 B.n386 163.367
R515 B.n388 B.n387 163.367
R516 B.n388 B.n95 163.367
R517 B.n392 B.n95 163.367
R518 B.n393 B.n392 163.367
R519 B.n394 B.n393 163.367
R520 B.n394 B.n93 163.367
R521 B.n398 B.n93 163.367
R522 B.n399 B.n398 163.367
R523 B.n400 B.n399 163.367
R524 B.n400 B.n91 163.367
R525 B.n404 B.n91 163.367
R526 B.n405 B.n404 163.367
R527 B.n406 B.n405 163.367
R528 B.n406 B.n89 163.367
R529 B.n410 B.n89 163.367
R530 B.n411 B.n410 163.367
R531 B.n412 B.n411 163.367
R532 B.n412 B.n87 163.367
R533 B.n416 B.n87 163.367
R534 B.n417 B.n416 163.367
R535 B.n418 B.n417 163.367
R536 B.n418 B.n85 163.367
R537 B.n422 B.n85 163.367
R538 B.n423 B.n422 163.367
R539 B.n424 B.n423 163.367
R540 B.n424 B.n83 163.367
R541 B.n428 B.n83 163.367
R542 B.n429 B.n428 163.367
R543 B.n430 B.n429 163.367
R544 B.n430 B.n81 163.367
R545 B.n434 B.n81 163.367
R546 B.n435 B.n434 163.367
R547 B.n436 B.n435 163.367
R548 B.n436 B.n79 163.367
R549 B.n440 B.n79 163.367
R550 B.n441 B.n440 163.367
R551 B.n442 B.n441 163.367
R552 B.n442 B.n77 163.367
R553 B.n446 B.n77 163.367
R554 B.n447 B.n446 163.367
R555 B.n448 B.n447 163.367
R556 B.n448 B.n75 163.367
R557 B.n452 B.n75 163.367
R558 B.n453 B.n452 163.367
R559 B.n454 B.n453 163.367
R560 B.n454 B.n73 163.367
R561 B.n458 B.n73 163.367
R562 B.n459 B.n458 163.367
R563 B.n460 B.n459 163.367
R564 B.n460 B.n71 163.367
R565 B.n464 B.n71 163.367
R566 B.n465 B.n464 163.367
R567 B.n466 B.n465 163.367
R568 B.n466 B.n69 163.367
R569 B.n470 B.n69 163.367
R570 B.n602 B.n21 163.367
R571 B.n598 B.n21 163.367
R572 B.n598 B.n597 163.367
R573 B.n597 B.n596 163.367
R574 B.n596 B.n23 163.367
R575 B.n592 B.n23 163.367
R576 B.n592 B.n591 163.367
R577 B.n591 B.n590 163.367
R578 B.n590 B.n25 163.367
R579 B.n586 B.n25 163.367
R580 B.n586 B.n585 163.367
R581 B.n585 B.n584 163.367
R582 B.n584 B.n27 163.367
R583 B.n580 B.n27 163.367
R584 B.n580 B.n579 163.367
R585 B.n579 B.n578 163.367
R586 B.n578 B.n29 163.367
R587 B.n574 B.n29 163.367
R588 B.n574 B.n573 163.367
R589 B.n573 B.n572 163.367
R590 B.n572 B.n31 163.367
R591 B.n568 B.n31 163.367
R592 B.n568 B.n567 163.367
R593 B.n567 B.n566 163.367
R594 B.n566 B.n33 163.367
R595 B.n562 B.n33 163.367
R596 B.n562 B.n561 163.367
R597 B.n561 B.n560 163.367
R598 B.n560 B.n35 163.367
R599 B.n556 B.n35 163.367
R600 B.n556 B.n555 163.367
R601 B.n555 B.n554 163.367
R602 B.n554 B.n37 163.367
R603 B.n550 B.n37 163.367
R604 B.n550 B.n549 163.367
R605 B.n549 B.n548 163.367
R606 B.n548 B.n39 163.367
R607 B.n544 B.n39 163.367
R608 B.n544 B.n543 163.367
R609 B.n543 B.n43 163.367
R610 B.n539 B.n43 163.367
R611 B.n539 B.n538 163.367
R612 B.n538 B.n537 163.367
R613 B.n537 B.n45 163.367
R614 B.n533 B.n45 163.367
R615 B.n533 B.n532 163.367
R616 B.n532 B.n531 163.367
R617 B.n531 B.n47 163.367
R618 B.n526 B.n47 163.367
R619 B.n526 B.n525 163.367
R620 B.n525 B.n524 163.367
R621 B.n524 B.n51 163.367
R622 B.n520 B.n51 163.367
R623 B.n520 B.n519 163.367
R624 B.n519 B.n518 163.367
R625 B.n518 B.n53 163.367
R626 B.n514 B.n53 163.367
R627 B.n514 B.n513 163.367
R628 B.n513 B.n512 163.367
R629 B.n512 B.n55 163.367
R630 B.n508 B.n55 163.367
R631 B.n508 B.n507 163.367
R632 B.n507 B.n506 163.367
R633 B.n506 B.n57 163.367
R634 B.n502 B.n57 163.367
R635 B.n502 B.n501 163.367
R636 B.n501 B.n500 163.367
R637 B.n500 B.n59 163.367
R638 B.n496 B.n59 163.367
R639 B.n496 B.n495 163.367
R640 B.n495 B.n494 163.367
R641 B.n494 B.n61 163.367
R642 B.n490 B.n61 163.367
R643 B.n490 B.n489 163.367
R644 B.n489 B.n488 163.367
R645 B.n488 B.n63 163.367
R646 B.n484 B.n63 163.367
R647 B.n484 B.n483 163.367
R648 B.n483 B.n482 163.367
R649 B.n482 B.n65 163.367
R650 B.n478 B.n65 163.367
R651 B.n478 B.n477 163.367
R652 B.n477 B.n476 163.367
R653 B.n476 B.n67 163.367
R654 B.n472 B.n67 163.367
R655 B.n472 B.n471 163.367
R656 B.n127 B.t1 110.834
R657 B.n49 B.t8 110.834
R658 B.n133 B.t4 110.82
R659 B.n41 B.t11 110.82
R660 B.n127 B.n126 63.0308
R661 B.n133 B.n132 63.0308
R662 B.n41 B.n40 63.0308
R663 B.n49 B.n48 63.0308
R664 B.n299 B.n127 59.5399
R665 B.n134 B.n133 59.5399
R666 B.n42 B.n41 59.5399
R667 B.n529 B.n49 59.5399
R668 B.n601 B.n20 31.6883
R669 B.n469 B.n68 31.6883
R670 B.n359 B.n106 31.6883
R671 B.n227 B.n154 31.6883
R672 B B.n659 18.0485
R673 B.n601 B.n600 10.6151
R674 B.n600 B.n599 10.6151
R675 B.n599 B.n22 10.6151
R676 B.n595 B.n22 10.6151
R677 B.n595 B.n594 10.6151
R678 B.n594 B.n593 10.6151
R679 B.n593 B.n24 10.6151
R680 B.n589 B.n24 10.6151
R681 B.n589 B.n588 10.6151
R682 B.n588 B.n587 10.6151
R683 B.n587 B.n26 10.6151
R684 B.n583 B.n26 10.6151
R685 B.n583 B.n582 10.6151
R686 B.n582 B.n581 10.6151
R687 B.n581 B.n28 10.6151
R688 B.n577 B.n28 10.6151
R689 B.n577 B.n576 10.6151
R690 B.n576 B.n575 10.6151
R691 B.n575 B.n30 10.6151
R692 B.n571 B.n30 10.6151
R693 B.n571 B.n570 10.6151
R694 B.n570 B.n569 10.6151
R695 B.n569 B.n32 10.6151
R696 B.n565 B.n32 10.6151
R697 B.n565 B.n564 10.6151
R698 B.n564 B.n563 10.6151
R699 B.n563 B.n34 10.6151
R700 B.n559 B.n34 10.6151
R701 B.n559 B.n558 10.6151
R702 B.n558 B.n557 10.6151
R703 B.n557 B.n36 10.6151
R704 B.n553 B.n36 10.6151
R705 B.n553 B.n552 10.6151
R706 B.n552 B.n551 10.6151
R707 B.n551 B.n38 10.6151
R708 B.n547 B.n38 10.6151
R709 B.n547 B.n546 10.6151
R710 B.n546 B.n545 10.6151
R711 B.n542 B.n541 10.6151
R712 B.n541 B.n540 10.6151
R713 B.n540 B.n44 10.6151
R714 B.n536 B.n44 10.6151
R715 B.n536 B.n535 10.6151
R716 B.n535 B.n534 10.6151
R717 B.n534 B.n46 10.6151
R718 B.n530 B.n46 10.6151
R719 B.n528 B.n527 10.6151
R720 B.n527 B.n50 10.6151
R721 B.n523 B.n50 10.6151
R722 B.n523 B.n522 10.6151
R723 B.n522 B.n521 10.6151
R724 B.n521 B.n52 10.6151
R725 B.n517 B.n52 10.6151
R726 B.n517 B.n516 10.6151
R727 B.n516 B.n515 10.6151
R728 B.n515 B.n54 10.6151
R729 B.n511 B.n54 10.6151
R730 B.n511 B.n510 10.6151
R731 B.n510 B.n509 10.6151
R732 B.n509 B.n56 10.6151
R733 B.n505 B.n56 10.6151
R734 B.n505 B.n504 10.6151
R735 B.n504 B.n503 10.6151
R736 B.n503 B.n58 10.6151
R737 B.n499 B.n58 10.6151
R738 B.n499 B.n498 10.6151
R739 B.n498 B.n497 10.6151
R740 B.n497 B.n60 10.6151
R741 B.n493 B.n60 10.6151
R742 B.n493 B.n492 10.6151
R743 B.n492 B.n491 10.6151
R744 B.n491 B.n62 10.6151
R745 B.n487 B.n62 10.6151
R746 B.n487 B.n486 10.6151
R747 B.n486 B.n485 10.6151
R748 B.n485 B.n64 10.6151
R749 B.n481 B.n64 10.6151
R750 B.n481 B.n480 10.6151
R751 B.n480 B.n479 10.6151
R752 B.n479 B.n66 10.6151
R753 B.n475 B.n66 10.6151
R754 B.n475 B.n474 10.6151
R755 B.n474 B.n473 10.6151
R756 B.n473 B.n68 10.6151
R757 B.n360 B.n359 10.6151
R758 B.n361 B.n360 10.6151
R759 B.n361 B.n104 10.6151
R760 B.n365 B.n104 10.6151
R761 B.n366 B.n365 10.6151
R762 B.n367 B.n366 10.6151
R763 B.n367 B.n102 10.6151
R764 B.n371 B.n102 10.6151
R765 B.n372 B.n371 10.6151
R766 B.n373 B.n372 10.6151
R767 B.n373 B.n100 10.6151
R768 B.n377 B.n100 10.6151
R769 B.n378 B.n377 10.6151
R770 B.n379 B.n378 10.6151
R771 B.n379 B.n98 10.6151
R772 B.n383 B.n98 10.6151
R773 B.n384 B.n383 10.6151
R774 B.n385 B.n384 10.6151
R775 B.n385 B.n96 10.6151
R776 B.n389 B.n96 10.6151
R777 B.n390 B.n389 10.6151
R778 B.n391 B.n390 10.6151
R779 B.n391 B.n94 10.6151
R780 B.n395 B.n94 10.6151
R781 B.n396 B.n395 10.6151
R782 B.n397 B.n396 10.6151
R783 B.n397 B.n92 10.6151
R784 B.n401 B.n92 10.6151
R785 B.n402 B.n401 10.6151
R786 B.n403 B.n402 10.6151
R787 B.n403 B.n90 10.6151
R788 B.n407 B.n90 10.6151
R789 B.n408 B.n407 10.6151
R790 B.n409 B.n408 10.6151
R791 B.n409 B.n88 10.6151
R792 B.n413 B.n88 10.6151
R793 B.n414 B.n413 10.6151
R794 B.n415 B.n414 10.6151
R795 B.n415 B.n86 10.6151
R796 B.n419 B.n86 10.6151
R797 B.n420 B.n419 10.6151
R798 B.n421 B.n420 10.6151
R799 B.n421 B.n84 10.6151
R800 B.n425 B.n84 10.6151
R801 B.n426 B.n425 10.6151
R802 B.n427 B.n426 10.6151
R803 B.n427 B.n82 10.6151
R804 B.n431 B.n82 10.6151
R805 B.n432 B.n431 10.6151
R806 B.n433 B.n432 10.6151
R807 B.n433 B.n80 10.6151
R808 B.n437 B.n80 10.6151
R809 B.n438 B.n437 10.6151
R810 B.n439 B.n438 10.6151
R811 B.n439 B.n78 10.6151
R812 B.n443 B.n78 10.6151
R813 B.n444 B.n443 10.6151
R814 B.n445 B.n444 10.6151
R815 B.n445 B.n76 10.6151
R816 B.n449 B.n76 10.6151
R817 B.n450 B.n449 10.6151
R818 B.n451 B.n450 10.6151
R819 B.n451 B.n74 10.6151
R820 B.n455 B.n74 10.6151
R821 B.n456 B.n455 10.6151
R822 B.n457 B.n456 10.6151
R823 B.n457 B.n72 10.6151
R824 B.n461 B.n72 10.6151
R825 B.n462 B.n461 10.6151
R826 B.n463 B.n462 10.6151
R827 B.n463 B.n70 10.6151
R828 B.n467 B.n70 10.6151
R829 B.n468 B.n467 10.6151
R830 B.n469 B.n468 10.6151
R831 B.n228 B.n227 10.6151
R832 B.n229 B.n228 10.6151
R833 B.n229 B.n152 10.6151
R834 B.n233 B.n152 10.6151
R835 B.n234 B.n233 10.6151
R836 B.n235 B.n234 10.6151
R837 B.n235 B.n150 10.6151
R838 B.n239 B.n150 10.6151
R839 B.n240 B.n239 10.6151
R840 B.n241 B.n240 10.6151
R841 B.n241 B.n148 10.6151
R842 B.n245 B.n148 10.6151
R843 B.n246 B.n245 10.6151
R844 B.n247 B.n246 10.6151
R845 B.n247 B.n146 10.6151
R846 B.n251 B.n146 10.6151
R847 B.n252 B.n251 10.6151
R848 B.n253 B.n252 10.6151
R849 B.n253 B.n144 10.6151
R850 B.n257 B.n144 10.6151
R851 B.n258 B.n257 10.6151
R852 B.n259 B.n258 10.6151
R853 B.n259 B.n142 10.6151
R854 B.n263 B.n142 10.6151
R855 B.n264 B.n263 10.6151
R856 B.n265 B.n264 10.6151
R857 B.n265 B.n140 10.6151
R858 B.n269 B.n140 10.6151
R859 B.n270 B.n269 10.6151
R860 B.n271 B.n270 10.6151
R861 B.n271 B.n138 10.6151
R862 B.n275 B.n138 10.6151
R863 B.n276 B.n275 10.6151
R864 B.n277 B.n276 10.6151
R865 B.n277 B.n136 10.6151
R866 B.n281 B.n136 10.6151
R867 B.n282 B.n281 10.6151
R868 B.n283 B.n282 10.6151
R869 B.n287 B.n286 10.6151
R870 B.n288 B.n287 10.6151
R871 B.n288 B.n130 10.6151
R872 B.n292 B.n130 10.6151
R873 B.n293 B.n292 10.6151
R874 B.n294 B.n293 10.6151
R875 B.n294 B.n128 10.6151
R876 B.n298 B.n128 10.6151
R877 B.n301 B.n300 10.6151
R878 B.n301 B.n124 10.6151
R879 B.n305 B.n124 10.6151
R880 B.n306 B.n305 10.6151
R881 B.n307 B.n306 10.6151
R882 B.n307 B.n122 10.6151
R883 B.n311 B.n122 10.6151
R884 B.n312 B.n311 10.6151
R885 B.n313 B.n312 10.6151
R886 B.n313 B.n120 10.6151
R887 B.n317 B.n120 10.6151
R888 B.n318 B.n317 10.6151
R889 B.n319 B.n318 10.6151
R890 B.n319 B.n118 10.6151
R891 B.n323 B.n118 10.6151
R892 B.n324 B.n323 10.6151
R893 B.n325 B.n324 10.6151
R894 B.n325 B.n116 10.6151
R895 B.n329 B.n116 10.6151
R896 B.n330 B.n329 10.6151
R897 B.n331 B.n330 10.6151
R898 B.n331 B.n114 10.6151
R899 B.n335 B.n114 10.6151
R900 B.n336 B.n335 10.6151
R901 B.n337 B.n336 10.6151
R902 B.n337 B.n112 10.6151
R903 B.n341 B.n112 10.6151
R904 B.n342 B.n341 10.6151
R905 B.n343 B.n342 10.6151
R906 B.n343 B.n110 10.6151
R907 B.n347 B.n110 10.6151
R908 B.n348 B.n347 10.6151
R909 B.n349 B.n348 10.6151
R910 B.n349 B.n108 10.6151
R911 B.n353 B.n108 10.6151
R912 B.n354 B.n353 10.6151
R913 B.n355 B.n354 10.6151
R914 B.n355 B.n106 10.6151
R915 B.n223 B.n154 10.6151
R916 B.n223 B.n222 10.6151
R917 B.n222 B.n221 10.6151
R918 B.n221 B.n156 10.6151
R919 B.n217 B.n156 10.6151
R920 B.n217 B.n216 10.6151
R921 B.n216 B.n215 10.6151
R922 B.n215 B.n158 10.6151
R923 B.n211 B.n158 10.6151
R924 B.n211 B.n210 10.6151
R925 B.n210 B.n209 10.6151
R926 B.n209 B.n160 10.6151
R927 B.n205 B.n160 10.6151
R928 B.n205 B.n204 10.6151
R929 B.n204 B.n203 10.6151
R930 B.n203 B.n162 10.6151
R931 B.n199 B.n162 10.6151
R932 B.n199 B.n198 10.6151
R933 B.n198 B.n197 10.6151
R934 B.n197 B.n164 10.6151
R935 B.n193 B.n164 10.6151
R936 B.n193 B.n192 10.6151
R937 B.n192 B.n191 10.6151
R938 B.n191 B.n166 10.6151
R939 B.n187 B.n166 10.6151
R940 B.n187 B.n186 10.6151
R941 B.n186 B.n185 10.6151
R942 B.n185 B.n168 10.6151
R943 B.n181 B.n168 10.6151
R944 B.n181 B.n180 10.6151
R945 B.n180 B.n179 10.6151
R946 B.n179 B.n170 10.6151
R947 B.n175 B.n170 10.6151
R948 B.n175 B.n174 10.6151
R949 B.n174 B.n173 10.6151
R950 B.n173 B.n0 10.6151
R951 B.n655 B.n1 10.6151
R952 B.n655 B.n654 10.6151
R953 B.n654 B.n653 10.6151
R954 B.n653 B.n4 10.6151
R955 B.n649 B.n4 10.6151
R956 B.n649 B.n648 10.6151
R957 B.n648 B.n647 10.6151
R958 B.n647 B.n6 10.6151
R959 B.n643 B.n6 10.6151
R960 B.n643 B.n642 10.6151
R961 B.n642 B.n641 10.6151
R962 B.n641 B.n8 10.6151
R963 B.n637 B.n8 10.6151
R964 B.n637 B.n636 10.6151
R965 B.n636 B.n635 10.6151
R966 B.n635 B.n10 10.6151
R967 B.n631 B.n10 10.6151
R968 B.n631 B.n630 10.6151
R969 B.n630 B.n629 10.6151
R970 B.n629 B.n12 10.6151
R971 B.n625 B.n12 10.6151
R972 B.n625 B.n624 10.6151
R973 B.n624 B.n623 10.6151
R974 B.n623 B.n14 10.6151
R975 B.n619 B.n14 10.6151
R976 B.n619 B.n618 10.6151
R977 B.n618 B.n617 10.6151
R978 B.n617 B.n16 10.6151
R979 B.n613 B.n16 10.6151
R980 B.n613 B.n612 10.6151
R981 B.n612 B.n611 10.6151
R982 B.n611 B.n18 10.6151
R983 B.n607 B.n18 10.6151
R984 B.n607 B.n606 10.6151
R985 B.n606 B.n605 10.6151
R986 B.n605 B.n20 10.6151
R987 B.n542 B.n42 6.5566
R988 B.n530 B.n529 6.5566
R989 B.n286 B.n134 6.5566
R990 B.n299 B.n298 6.5566
R991 B.n545 B.n42 4.05904
R992 B.n529 B.n528 4.05904
R993 B.n283 B.n134 4.05904
R994 B.n300 B.n299 4.05904
R995 B.n659 B.n0 2.81026
R996 B.n659 B.n1 2.81026
R997 VN.n1 VN.t1 125.532
R998 VN.n0 VN.t2 125.532
R999 VN.n0 VN.t3 124.561
R1000 VN.n1 VN.t0 124.561
R1001 VN VN.n1 49.8961
R1002 VN VN.n0 3.16503
R1003 VDD2.n2 VDD2.n0 117.347
R1004 VDD2.n2 VDD2.n1 75.6927
R1005 VDD2.n1 VDD2.t2 2.93947
R1006 VDD2.n1 VDD2.t1 2.93947
R1007 VDD2.n0 VDD2.t3 2.93947
R1008 VDD2.n0 VDD2.t0 2.93947
R1009 VDD2 VDD2.n2 0.0586897
R1010 VTAIL.n5 VTAIL.t0 61.953
R1011 VTAIL.n4 VTAIL.t6 61.953
R1012 VTAIL.n3 VTAIL.t7 61.953
R1013 VTAIL.n7 VTAIL.t4 61.9529
R1014 VTAIL.n0 VTAIL.t5 61.9529
R1015 VTAIL.n1 VTAIL.t3 61.9529
R1016 VTAIL.n2 VTAIL.t1 61.9529
R1017 VTAIL.n6 VTAIL.t2 61.9529
R1018 VTAIL.n7 VTAIL.n6 24.7031
R1019 VTAIL.n3 VTAIL.n2 24.7031
R1020 VTAIL.n4 VTAIL.n3 2.80222
R1021 VTAIL.n6 VTAIL.n5 2.80222
R1022 VTAIL.n2 VTAIL.n1 2.80222
R1023 VTAIL VTAIL.n0 1.45955
R1024 VTAIL VTAIL.n7 1.34317
R1025 VTAIL.n5 VTAIL.n4 0.470328
R1026 VTAIL.n1 VTAIL.n0 0.470328
R1027 VP.n15 VP.n14 161.3
R1028 VP.n13 VP.n1 161.3
R1029 VP.n12 VP.n11 161.3
R1030 VP.n10 VP.n2 161.3
R1031 VP.n9 VP.n8 161.3
R1032 VP.n7 VP.n3 161.3
R1033 VP.n4 VP.t3 125.532
R1034 VP.n4 VP.t1 124.561
R1035 VP.n6 VP.t2 91.2834
R1036 VP.n0 VP.t0 91.2834
R1037 VP.n6 VP.n5 71.6334
R1038 VP.n16 VP.n0 71.6334
R1039 VP.n12 VP.n2 56.4773
R1040 VP.n5 VP.n4 49.7306
R1041 VP.n8 VP.n7 24.3439
R1042 VP.n8 VP.n2 24.3439
R1043 VP.n13 VP.n12 24.3439
R1044 VP.n14 VP.n13 24.3439
R1045 VP.n7 VP.n6 18.2581
R1046 VP.n14 VP.n0 18.2581
R1047 VP.n5 VP.n3 0.355081
R1048 VP.n16 VP.n15 0.355081
R1049 VP VP.n16 0.26685
R1050 VP.n9 VP.n3 0.189894
R1051 VP.n10 VP.n9 0.189894
R1052 VP.n11 VP.n10 0.189894
R1053 VP.n11 VP.n1 0.189894
R1054 VP.n15 VP.n1 0.189894
R1055 VDD1 VDD1.n1 117.871
R1056 VDD1 VDD1.n0 75.7509
R1057 VDD1.n0 VDD1.t0 2.93947
R1058 VDD1.n0 VDD1.t2 2.93947
R1059 VDD1.n1 VDD1.t1 2.93947
R1060 VDD1.n1 VDD1.t3 2.93947
C0 VDD1 VTAIL 5.25571f
C1 w_n2920_n3180# VN 5.00173f
C2 VP w_n2920_n3180# 5.37792f
C3 VTAIL B 4.77186f
C4 w_n2920_n3180# VDD2 1.55448f
C5 VDD1 w_n2920_n3180# 1.49127f
C6 VP VN 6.25622f
C7 VDD2 VN 4.48717f
C8 VP VDD2 0.414474f
C9 VDD1 VN 0.149096f
C10 w_n2920_n3180# B 9.3758f
C11 VDD1 VP 4.75173f
C12 VDD1 VDD2 1.10274f
C13 B VN 1.15436f
C14 w_n2920_n3180# VTAIL 3.77366f
C15 VP B 1.78012f
C16 B VDD2 1.34988f
C17 VTAIL VN 4.49293f
C18 VP VTAIL 4.50704f
C19 VDD1 B 1.29242f
C20 VTAIL VDD2 5.31206f
C21 VDD2 VSUBS 0.977687f
C22 VDD1 VSUBS 5.84581f
C23 VTAIL VSUBS 1.210846f
C24 VN VSUBS 5.60931f
C25 VP VSUBS 2.430732f
C26 B VSUBS 4.472743f
C27 w_n2920_n3180# VSUBS 0.114476p
C28 VDD1.t0 VSUBS 0.240982f
C29 VDD1.t2 VSUBS 0.240982f
C30 VDD1.n0 VSUBS 1.85552f
C31 VDD1.t1 VSUBS 0.240982f
C32 VDD1.t3 VSUBS 0.240982f
C33 VDD1.n1 VSUBS 2.57495f
C34 VP.t0 VSUBS 2.89688f
C35 VP.n0 VSUBS 1.15065f
C36 VP.n1 VSUBS 0.033002f
C37 VP.n2 VSUBS 0.048387f
C38 VP.n3 VSUBS 0.053273f
C39 VP.t2 VSUBS 2.89688f
C40 VP.t3 VSUBS 3.2396f
C41 VP.t1 VSUBS 3.23008f
C42 VP.n4 VSUBS 3.89962f
C43 VP.n5 VSUBS 1.83768f
C44 VP.n6 VSUBS 1.15065f
C45 VP.n7 VSUBS 0.054186f
C46 VP.n8 VSUBS 0.061816f
C47 VP.n9 VSUBS 0.033002f
C48 VP.n10 VSUBS 0.033002f
C49 VP.n11 VSUBS 0.033002f
C50 VP.n12 VSUBS 0.048387f
C51 VP.n13 VSUBS 0.061816f
C52 VP.n14 VSUBS 0.054186f
C53 VP.n15 VSUBS 0.053273f
C54 VP.n16 VSUBS 0.070179f
C55 VTAIL.t5 VSUBS 2.00559f
C56 VTAIL.n0 VSUBS 0.782498f
C57 VTAIL.t3 VSUBS 2.00559f
C58 VTAIL.n1 VSUBS 0.887939f
C59 VTAIL.t1 VSUBS 2.00559f
C60 VTAIL.n2 VSUBS 2.15088f
C61 VTAIL.t7 VSUBS 2.00561f
C62 VTAIL.n3 VSUBS 2.15086f
C63 VTAIL.t6 VSUBS 2.00561f
C64 VTAIL.n4 VSUBS 0.887925f
C65 VTAIL.t0 VSUBS 2.00561f
C66 VTAIL.n5 VSUBS 0.887925f
C67 VTAIL.t2 VSUBS 2.00559f
C68 VTAIL.n6 VSUBS 2.15088f
C69 VTAIL.t4 VSUBS 2.00559f
C70 VTAIL.n7 VSUBS 2.0363f
C71 VDD2.t3 VSUBS 0.236206f
C72 VDD2.t0 VSUBS 0.236206f
C73 VDD2.n0 VSUBS 2.49918f
C74 VDD2.t2 VSUBS 0.236206f
C75 VDD2.t1 VSUBS 0.236206f
C76 VDD2.n1 VSUBS 1.81816f
C77 VDD2.n2 VSUBS 4.28803f
C78 VN.t3 VSUBS 3.11552f
C79 VN.t2 VSUBS 3.12471f
C80 VN.n0 VSUBS 1.95365f
C81 VN.t1 VSUBS 3.12471f
C82 VN.t0 VSUBS 3.11552f
C83 VN.n1 VSUBS 3.77427f
C84 B.n0 VSUBS 0.004258f
C85 B.n1 VSUBS 0.004258f
C86 B.n2 VSUBS 0.006733f
C87 B.n3 VSUBS 0.006733f
C88 B.n4 VSUBS 0.006733f
C89 B.n5 VSUBS 0.006733f
C90 B.n6 VSUBS 0.006733f
C91 B.n7 VSUBS 0.006733f
C92 B.n8 VSUBS 0.006733f
C93 B.n9 VSUBS 0.006733f
C94 B.n10 VSUBS 0.006733f
C95 B.n11 VSUBS 0.006733f
C96 B.n12 VSUBS 0.006733f
C97 B.n13 VSUBS 0.006733f
C98 B.n14 VSUBS 0.006733f
C99 B.n15 VSUBS 0.006733f
C100 B.n16 VSUBS 0.006733f
C101 B.n17 VSUBS 0.006733f
C102 B.n18 VSUBS 0.006733f
C103 B.n19 VSUBS 0.006733f
C104 B.n20 VSUBS 0.015297f
C105 B.n21 VSUBS 0.006733f
C106 B.n22 VSUBS 0.006733f
C107 B.n23 VSUBS 0.006733f
C108 B.n24 VSUBS 0.006733f
C109 B.n25 VSUBS 0.006733f
C110 B.n26 VSUBS 0.006733f
C111 B.n27 VSUBS 0.006733f
C112 B.n28 VSUBS 0.006733f
C113 B.n29 VSUBS 0.006733f
C114 B.n30 VSUBS 0.006733f
C115 B.n31 VSUBS 0.006733f
C116 B.n32 VSUBS 0.006733f
C117 B.n33 VSUBS 0.006733f
C118 B.n34 VSUBS 0.006733f
C119 B.n35 VSUBS 0.006733f
C120 B.n36 VSUBS 0.006733f
C121 B.n37 VSUBS 0.006733f
C122 B.n38 VSUBS 0.006733f
C123 B.n39 VSUBS 0.006733f
C124 B.t11 VSUBS 0.343546f
C125 B.t10 VSUBS 0.365538f
C126 B.t9 VSUBS 1.43263f
C127 B.n40 VSUBS 0.197118f
C128 B.n41 VSUBS 0.070262f
C129 B.n42 VSUBS 0.0156f
C130 B.n43 VSUBS 0.006733f
C131 B.n44 VSUBS 0.006733f
C132 B.n45 VSUBS 0.006733f
C133 B.n46 VSUBS 0.006733f
C134 B.n47 VSUBS 0.006733f
C135 B.t8 VSUBS 0.34354f
C136 B.t7 VSUBS 0.365533f
C137 B.t6 VSUBS 1.43263f
C138 B.n48 VSUBS 0.197123f
C139 B.n49 VSUBS 0.070268f
C140 B.n50 VSUBS 0.006733f
C141 B.n51 VSUBS 0.006733f
C142 B.n52 VSUBS 0.006733f
C143 B.n53 VSUBS 0.006733f
C144 B.n54 VSUBS 0.006733f
C145 B.n55 VSUBS 0.006733f
C146 B.n56 VSUBS 0.006733f
C147 B.n57 VSUBS 0.006733f
C148 B.n58 VSUBS 0.006733f
C149 B.n59 VSUBS 0.006733f
C150 B.n60 VSUBS 0.006733f
C151 B.n61 VSUBS 0.006733f
C152 B.n62 VSUBS 0.006733f
C153 B.n63 VSUBS 0.006733f
C154 B.n64 VSUBS 0.006733f
C155 B.n65 VSUBS 0.006733f
C156 B.n66 VSUBS 0.006733f
C157 B.n67 VSUBS 0.006733f
C158 B.n68 VSUBS 0.014777f
C159 B.n69 VSUBS 0.006733f
C160 B.n70 VSUBS 0.006733f
C161 B.n71 VSUBS 0.006733f
C162 B.n72 VSUBS 0.006733f
C163 B.n73 VSUBS 0.006733f
C164 B.n74 VSUBS 0.006733f
C165 B.n75 VSUBS 0.006733f
C166 B.n76 VSUBS 0.006733f
C167 B.n77 VSUBS 0.006733f
C168 B.n78 VSUBS 0.006733f
C169 B.n79 VSUBS 0.006733f
C170 B.n80 VSUBS 0.006733f
C171 B.n81 VSUBS 0.006733f
C172 B.n82 VSUBS 0.006733f
C173 B.n83 VSUBS 0.006733f
C174 B.n84 VSUBS 0.006733f
C175 B.n85 VSUBS 0.006733f
C176 B.n86 VSUBS 0.006733f
C177 B.n87 VSUBS 0.006733f
C178 B.n88 VSUBS 0.006733f
C179 B.n89 VSUBS 0.006733f
C180 B.n90 VSUBS 0.006733f
C181 B.n91 VSUBS 0.006733f
C182 B.n92 VSUBS 0.006733f
C183 B.n93 VSUBS 0.006733f
C184 B.n94 VSUBS 0.006733f
C185 B.n95 VSUBS 0.006733f
C186 B.n96 VSUBS 0.006733f
C187 B.n97 VSUBS 0.006733f
C188 B.n98 VSUBS 0.006733f
C189 B.n99 VSUBS 0.006733f
C190 B.n100 VSUBS 0.006733f
C191 B.n101 VSUBS 0.006733f
C192 B.n102 VSUBS 0.006733f
C193 B.n103 VSUBS 0.006733f
C194 B.n104 VSUBS 0.006733f
C195 B.n105 VSUBS 0.006733f
C196 B.n106 VSUBS 0.015597f
C197 B.n107 VSUBS 0.006733f
C198 B.n108 VSUBS 0.006733f
C199 B.n109 VSUBS 0.006733f
C200 B.n110 VSUBS 0.006733f
C201 B.n111 VSUBS 0.006733f
C202 B.n112 VSUBS 0.006733f
C203 B.n113 VSUBS 0.006733f
C204 B.n114 VSUBS 0.006733f
C205 B.n115 VSUBS 0.006733f
C206 B.n116 VSUBS 0.006733f
C207 B.n117 VSUBS 0.006733f
C208 B.n118 VSUBS 0.006733f
C209 B.n119 VSUBS 0.006733f
C210 B.n120 VSUBS 0.006733f
C211 B.n121 VSUBS 0.006733f
C212 B.n122 VSUBS 0.006733f
C213 B.n123 VSUBS 0.006733f
C214 B.n124 VSUBS 0.006733f
C215 B.n125 VSUBS 0.006733f
C216 B.t1 VSUBS 0.34354f
C217 B.t2 VSUBS 0.365533f
C218 B.t0 VSUBS 1.43263f
C219 B.n126 VSUBS 0.197123f
C220 B.n127 VSUBS 0.070268f
C221 B.n128 VSUBS 0.006733f
C222 B.n129 VSUBS 0.006733f
C223 B.n130 VSUBS 0.006733f
C224 B.n131 VSUBS 0.006733f
C225 B.t4 VSUBS 0.343546f
C226 B.t5 VSUBS 0.365538f
C227 B.t3 VSUBS 1.43263f
C228 B.n132 VSUBS 0.197118f
C229 B.n133 VSUBS 0.070262f
C230 B.n134 VSUBS 0.0156f
C231 B.n135 VSUBS 0.006733f
C232 B.n136 VSUBS 0.006733f
C233 B.n137 VSUBS 0.006733f
C234 B.n138 VSUBS 0.006733f
C235 B.n139 VSUBS 0.006733f
C236 B.n140 VSUBS 0.006733f
C237 B.n141 VSUBS 0.006733f
C238 B.n142 VSUBS 0.006733f
C239 B.n143 VSUBS 0.006733f
C240 B.n144 VSUBS 0.006733f
C241 B.n145 VSUBS 0.006733f
C242 B.n146 VSUBS 0.006733f
C243 B.n147 VSUBS 0.006733f
C244 B.n148 VSUBS 0.006733f
C245 B.n149 VSUBS 0.006733f
C246 B.n150 VSUBS 0.006733f
C247 B.n151 VSUBS 0.006733f
C248 B.n152 VSUBS 0.006733f
C249 B.n153 VSUBS 0.006733f
C250 B.n154 VSUBS 0.015297f
C251 B.n155 VSUBS 0.006733f
C252 B.n156 VSUBS 0.006733f
C253 B.n157 VSUBS 0.006733f
C254 B.n158 VSUBS 0.006733f
C255 B.n159 VSUBS 0.006733f
C256 B.n160 VSUBS 0.006733f
C257 B.n161 VSUBS 0.006733f
C258 B.n162 VSUBS 0.006733f
C259 B.n163 VSUBS 0.006733f
C260 B.n164 VSUBS 0.006733f
C261 B.n165 VSUBS 0.006733f
C262 B.n166 VSUBS 0.006733f
C263 B.n167 VSUBS 0.006733f
C264 B.n168 VSUBS 0.006733f
C265 B.n169 VSUBS 0.006733f
C266 B.n170 VSUBS 0.006733f
C267 B.n171 VSUBS 0.006733f
C268 B.n172 VSUBS 0.006733f
C269 B.n173 VSUBS 0.006733f
C270 B.n174 VSUBS 0.006733f
C271 B.n175 VSUBS 0.006733f
C272 B.n176 VSUBS 0.006733f
C273 B.n177 VSUBS 0.006733f
C274 B.n178 VSUBS 0.006733f
C275 B.n179 VSUBS 0.006733f
C276 B.n180 VSUBS 0.006733f
C277 B.n181 VSUBS 0.006733f
C278 B.n182 VSUBS 0.006733f
C279 B.n183 VSUBS 0.006733f
C280 B.n184 VSUBS 0.006733f
C281 B.n185 VSUBS 0.006733f
C282 B.n186 VSUBS 0.006733f
C283 B.n187 VSUBS 0.006733f
C284 B.n188 VSUBS 0.006733f
C285 B.n189 VSUBS 0.006733f
C286 B.n190 VSUBS 0.006733f
C287 B.n191 VSUBS 0.006733f
C288 B.n192 VSUBS 0.006733f
C289 B.n193 VSUBS 0.006733f
C290 B.n194 VSUBS 0.006733f
C291 B.n195 VSUBS 0.006733f
C292 B.n196 VSUBS 0.006733f
C293 B.n197 VSUBS 0.006733f
C294 B.n198 VSUBS 0.006733f
C295 B.n199 VSUBS 0.006733f
C296 B.n200 VSUBS 0.006733f
C297 B.n201 VSUBS 0.006733f
C298 B.n202 VSUBS 0.006733f
C299 B.n203 VSUBS 0.006733f
C300 B.n204 VSUBS 0.006733f
C301 B.n205 VSUBS 0.006733f
C302 B.n206 VSUBS 0.006733f
C303 B.n207 VSUBS 0.006733f
C304 B.n208 VSUBS 0.006733f
C305 B.n209 VSUBS 0.006733f
C306 B.n210 VSUBS 0.006733f
C307 B.n211 VSUBS 0.006733f
C308 B.n212 VSUBS 0.006733f
C309 B.n213 VSUBS 0.006733f
C310 B.n214 VSUBS 0.006733f
C311 B.n215 VSUBS 0.006733f
C312 B.n216 VSUBS 0.006733f
C313 B.n217 VSUBS 0.006733f
C314 B.n218 VSUBS 0.006733f
C315 B.n219 VSUBS 0.006733f
C316 B.n220 VSUBS 0.006733f
C317 B.n221 VSUBS 0.006733f
C318 B.n222 VSUBS 0.006733f
C319 B.n223 VSUBS 0.006733f
C320 B.n224 VSUBS 0.006733f
C321 B.n225 VSUBS 0.015297f
C322 B.n226 VSUBS 0.015597f
C323 B.n227 VSUBS 0.015597f
C324 B.n228 VSUBS 0.006733f
C325 B.n229 VSUBS 0.006733f
C326 B.n230 VSUBS 0.006733f
C327 B.n231 VSUBS 0.006733f
C328 B.n232 VSUBS 0.006733f
C329 B.n233 VSUBS 0.006733f
C330 B.n234 VSUBS 0.006733f
C331 B.n235 VSUBS 0.006733f
C332 B.n236 VSUBS 0.006733f
C333 B.n237 VSUBS 0.006733f
C334 B.n238 VSUBS 0.006733f
C335 B.n239 VSUBS 0.006733f
C336 B.n240 VSUBS 0.006733f
C337 B.n241 VSUBS 0.006733f
C338 B.n242 VSUBS 0.006733f
C339 B.n243 VSUBS 0.006733f
C340 B.n244 VSUBS 0.006733f
C341 B.n245 VSUBS 0.006733f
C342 B.n246 VSUBS 0.006733f
C343 B.n247 VSUBS 0.006733f
C344 B.n248 VSUBS 0.006733f
C345 B.n249 VSUBS 0.006733f
C346 B.n250 VSUBS 0.006733f
C347 B.n251 VSUBS 0.006733f
C348 B.n252 VSUBS 0.006733f
C349 B.n253 VSUBS 0.006733f
C350 B.n254 VSUBS 0.006733f
C351 B.n255 VSUBS 0.006733f
C352 B.n256 VSUBS 0.006733f
C353 B.n257 VSUBS 0.006733f
C354 B.n258 VSUBS 0.006733f
C355 B.n259 VSUBS 0.006733f
C356 B.n260 VSUBS 0.006733f
C357 B.n261 VSUBS 0.006733f
C358 B.n262 VSUBS 0.006733f
C359 B.n263 VSUBS 0.006733f
C360 B.n264 VSUBS 0.006733f
C361 B.n265 VSUBS 0.006733f
C362 B.n266 VSUBS 0.006733f
C363 B.n267 VSUBS 0.006733f
C364 B.n268 VSUBS 0.006733f
C365 B.n269 VSUBS 0.006733f
C366 B.n270 VSUBS 0.006733f
C367 B.n271 VSUBS 0.006733f
C368 B.n272 VSUBS 0.006733f
C369 B.n273 VSUBS 0.006733f
C370 B.n274 VSUBS 0.006733f
C371 B.n275 VSUBS 0.006733f
C372 B.n276 VSUBS 0.006733f
C373 B.n277 VSUBS 0.006733f
C374 B.n278 VSUBS 0.006733f
C375 B.n279 VSUBS 0.006733f
C376 B.n280 VSUBS 0.006733f
C377 B.n281 VSUBS 0.006733f
C378 B.n282 VSUBS 0.006733f
C379 B.n283 VSUBS 0.004654f
C380 B.n284 VSUBS 0.006733f
C381 B.n285 VSUBS 0.006733f
C382 B.n286 VSUBS 0.005446f
C383 B.n287 VSUBS 0.006733f
C384 B.n288 VSUBS 0.006733f
C385 B.n289 VSUBS 0.006733f
C386 B.n290 VSUBS 0.006733f
C387 B.n291 VSUBS 0.006733f
C388 B.n292 VSUBS 0.006733f
C389 B.n293 VSUBS 0.006733f
C390 B.n294 VSUBS 0.006733f
C391 B.n295 VSUBS 0.006733f
C392 B.n296 VSUBS 0.006733f
C393 B.n297 VSUBS 0.006733f
C394 B.n298 VSUBS 0.005446f
C395 B.n299 VSUBS 0.0156f
C396 B.n300 VSUBS 0.004654f
C397 B.n301 VSUBS 0.006733f
C398 B.n302 VSUBS 0.006733f
C399 B.n303 VSUBS 0.006733f
C400 B.n304 VSUBS 0.006733f
C401 B.n305 VSUBS 0.006733f
C402 B.n306 VSUBS 0.006733f
C403 B.n307 VSUBS 0.006733f
C404 B.n308 VSUBS 0.006733f
C405 B.n309 VSUBS 0.006733f
C406 B.n310 VSUBS 0.006733f
C407 B.n311 VSUBS 0.006733f
C408 B.n312 VSUBS 0.006733f
C409 B.n313 VSUBS 0.006733f
C410 B.n314 VSUBS 0.006733f
C411 B.n315 VSUBS 0.006733f
C412 B.n316 VSUBS 0.006733f
C413 B.n317 VSUBS 0.006733f
C414 B.n318 VSUBS 0.006733f
C415 B.n319 VSUBS 0.006733f
C416 B.n320 VSUBS 0.006733f
C417 B.n321 VSUBS 0.006733f
C418 B.n322 VSUBS 0.006733f
C419 B.n323 VSUBS 0.006733f
C420 B.n324 VSUBS 0.006733f
C421 B.n325 VSUBS 0.006733f
C422 B.n326 VSUBS 0.006733f
C423 B.n327 VSUBS 0.006733f
C424 B.n328 VSUBS 0.006733f
C425 B.n329 VSUBS 0.006733f
C426 B.n330 VSUBS 0.006733f
C427 B.n331 VSUBS 0.006733f
C428 B.n332 VSUBS 0.006733f
C429 B.n333 VSUBS 0.006733f
C430 B.n334 VSUBS 0.006733f
C431 B.n335 VSUBS 0.006733f
C432 B.n336 VSUBS 0.006733f
C433 B.n337 VSUBS 0.006733f
C434 B.n338 VSUBS 0.006733f
C435 B.n339 VSUBS 0.006733f
C436 B.n340 VSUBS 0.006733f
C437 B.n341 VSUBS 0.006733f
C438 B.n342 VSUBS 0.006733f
C439 B.n343 VSUBS 0.006733f
C440 B.n344 VSUBS 0.006733f
C441 B.n345 VSUBS 0.006733f
C442 B.n346 VSUBS 0.006733f
C443 B.n347 VSUBS 0.006733f
C444 B.n348 VSUBS 0.006733f
C445 B.n349 VSUBS 0.006733f
C446 B.n350 VSUBS 0.006733f
C447 B.n351 VSUBS 0.006733f
C448 B.n352 VSUBS 0.006733f
C449 B.n353 VSUBS 0.006733f
C450 B.n354 VSUBS 0.006733f
C451 B.n355 VSUBS 0.006733f
C452 B.n356 VSUBS 0.006733f
C453 B.n357 VSUBS 0.015597f
C454 B.n358 VSUBS 0.015297f
C455 B.n359 VSUBS 0.015297f
C456 B.n360 VSUBS 0.006733f
C457 B.n361 VSUBS 0.006733f
C458 B.n362 VSUBS 0.006733f
C459 B.n363 VSUBS 0.006733f
C460 B.n364 VSUBS 0.006733f
C461 B.n365 VSUBS 0.006733f
C462 B.n366 VSUBS 0.006733f
C463 B.n367 VSUBS 0.006733f
C464 B.n368 VSUBS 0.006733f
C465 B.n369 VSUBS 0.006733f
C466 B.n370 VSUBS 0.006733f
C467 B.n371 VSUBS 0.006733f
C468 B.n372 VSUBS 0.006733f
C469 B.n373 VSUBS 0.006733f
C470 B.n374 VSUBS 0.006733f
C471 B.n375 VSUBS 0.006733f
C472 B.n376 VSUBS 0.006733f
C473 B.n377 VSUBS 0.006733f
C474 B.n378 VSUBS 0.006733f
C475 B.n379 VSUBS 0.006733f
C476 B.n380 VSUBS 0.006733f
C477 B.n381 VSUBS 0.006733f
C478 B.n382 VSUBS 0.006733f
C479 B.n383 VSUBS 0.006733f
C480 B.n384 VSUBS 0.006733f
C481 B.n385 VSUBS 0.006733f
C482 B.n386 VSUBS 0.006733f
C483 B.n387 VSUBS 0.006733f
C484 B.n388 VSUBS 0.006733f
C485 B.n389 VSUBS 0.006733f
C486 B.n390 VSUBS 0.006733f
C487 B.n391 VSUBS 0.006733f
C488 B.n392 VSUBS 0.006733f
C489 B.n393 VSUBS 0.006733f
C490 B.n394 VSUBS 0.006733f
C491 B.n395 VSUBS 0.006733f
C492 B.n396 VSUBS 0.006733f
C493 B.n397 VSUBS 0.006733f
C494 B.n398 VSUBS 0.006733f
C495 B.n399 VSUBS 0.006733f
C496 B.n400 VSUBS 0.006733f
C497 B.n401 VSUBS 0.006733f
C498 B.n402 VSUBS 0.006733f
C499 B.n403 VSUBS 0.006733f
C500 B.n404 VSUBS 0.006733f
C501 B.n405 VSUBS 0.006733f
C502 B.n406 VSUBS 0.006733f
C503 B.n407 VSUBS 0.006733f
C504 B.n408 VSUBS 0.006733f
C505 B.n409 VSUBS 0.006733f
C506 B.n410 VSUBS 0.006733f
C507 B.n411 VSUBS 0.006733f
C508 B.n412 VSUBS 0.006733f
C509 B.n413 VSUBS 0.006733f
C510 B.n414 VSUBS 0.006733f
C511 B.n415 VSUBS 0.006733f
C512 B.n416 VSUBS 0.006733f
C513 B.n417 VSUBS 0.006733f
C514 B.n418 VSUBS 0.006733f
C515 B.n419 VSUBS 0.006733f
C516 B.n420 VSUBS 0.006733f
C517 B.n421 VSUBS 0.006733f
C518 B.n422 VSUBS 0.006733f
C519 B.n423 VSUBS 0.006733f
C520 B.n424 VSUBS 0.006733f
C521 B.n425 VSUBS 0.006733f
C522 B.n426 VSUBS 0.006733f
C523 B.n427 VSUBS 0.006733f
C524 B.n428 VSUBS 0.006733f
C525 B.n429 VSUBS 0.006733f
C526 B.n430 VSUBS 0.006733f
C527 B.n431 VSUBS 0.006733f
C528 B.n432 VSUBS 0.006733f
C529 B.n433 VSUBS 0.006733f
C530 B.n434 VSUBS 0.006733f
C531 B.n435 VSUBS 0.006733f
C532 B.n436 VSUBS 0.006733f
C533 B.n437 VSUBS 0.006733f
C534 B.n438 VSUBS 0.006733f
C535 B.n439 VSUBS 0.006733f
C536 B.n440 VSUBS 0.006733f
C537 B.n441 VSUBS 0.006733f
C538 B.n442 VSUBS 0.006733f
C539 B.n443 VSUBS 0.006733f
C540 B.n444 VSUBS 0.006733f
C541 B.n445 VSUBS 0.006733f
C542 B.n446 VSUBS 0.006733f
C543 B.n447 VSUBS 0.006733f
C544 B.n448 VSUBS 0.006733f
C545 B.n449 VSUBS 0.006733f
C546 B.n450 VSUBS 0.006733f
C547 B.n451 VSUBS 0.006733f
C548 B.n452 VSUBS 0.006733f
C549 B.n453 VSUBS 0.006733f
C550 B.n454 VSUBS 0.006733f
C551 B.n455 VSUBS 0.006733f
C552 B.n456 VSUBS 0.006733f
C553 B.n457 VSUBS 0.006733f
C554 B.n458 VSUBS 0.006733f
C555 B.n459 VSUBS 0.006733f
C556 B.n460 VSUBS 0.006733f
C557 B.n461 VSUBS 0.006733f
C558 B.n462 VSUBS 0.006733f
C559 B.n463 VSUBS 0.006733f
C560 B.n464 VSUBS 0.006733f
C561 B.n465 VSUBS 0.006733f
C562 B.n466 VSUBS 0.006733f
C563 B.n467 VSUBS 0.006733f
C564 B.n468 VSUBS 0.006733f
C565 B.n469 VSUBS 0.016117f
C566 B.n470 VSUBS 0.015297f
C567 B.n471 VSUBS 0.015597f
C568 B.n472 VSUBS 0.006733f
C569 B.n473 VSUBS 0.006733f
C570 B.n474 VSUBS 0.006733f
C571 B.n475 VSUBS 0.006733f
C572 B.n476 VSUBS 0.006733f
C573 B.n477 VSUBS 0.006733f
C574 B.n478 VSUBS 0.006733f
C575 B.n479 VSUBS 0.006733f
C576 B.n480 VSUBS 0.006733f
C577 B.n481 VSUBS 0.006733f
C578 B.n482 VSUBS 0.006733f
C579 B.n483 VSUBS 0.006733f
C580 B.n484 VSUBS 0.006733f
C581 B.n485 VSUBS 0.006733f
C582 B.n486 VSUBS 0.006733f
C583 B.n487 VSUBS 0.006733f
C584 B.n488 VSUBS 0.006733f
C585 B.n489 VSUBS 0.006733f
C586 B.n490 VSUBS 0.006733f
C587 B.n491 VSUBS 0.006733f
C588 B.n492 VSUBS 0.006733f
C589 B.n493 VSUBS 0.006733f
C590 B.n494 VSUBS 0.006733f
C591 B.n495 VSUBS 0.006733f
C592 B.n496 VSUBS 0.006733f
C593 B.n497 VSUBS 0.006733f
C594 B.n498 VSUBS 0.006733f
C595 B.n499 VSUBS 0.006733f
C596 B.n500 VSUBS 0.006733f
C597 B.n501 VSUBS 0.006733f
C598 B.n502 VSUBS 0.006733f
C599 B.n503 VSUBS 0.006733f
C600 B.n504 VSUBS 0.006733f
C601 B.n505 VSUBS 0.006733f
C602 B.n506 VSUBS 0.006733f
C603 B.n507 VSUBS 0.006733f
C604 B.n508 VSUBS 0.006733f
C605 B.n509 VSUBS 0.006733f
C606 B.n510 VSUBS 0.006733f
C607 B.n511 VSUBS 0.006733f
C608 B.n512 VSUBS 0.006733f
C609 B.n513 VSUBS 0.006733f
C610 B.n514 VSUBS 0.006733f
C611 B.n515 VSUBS 0.006733f
C612 B.n516 VSUBS 0.006733f
C613 B.n517 VSUBS 0.006733f
C614 B.n518 VSUBS 0.006733f
C615 B.n519 VSUBS 0.006733f
C616 B.n520 VSUBS 0.006733f
C617 B.n521 VSUBS 0.006733f
C618 B.n522 VSUBS 0.006733f
C619 B.n523 VSUBS 0.006733f
C620 B.n524 VSUBS 0.006733f
C621 B.n525 VSUBS 0.006733f
C622 B.n526 VSUBS 0.006733f
C623 B.n527 VSUBS 0.006733f
C624 B.n528 VSUBS 0.004654f
C625 B.n529 VSUBS 0.0156f
C626 B.n530 VSUBS 0.005446f
C627 B.n531 VSUBS 0.006733f
C628 B.n532 VSUBS 0.006733f
C629 B.n533 VSUBS 0.006733f
C630 B.n534 VSUBS 0.006733f
C631 B.n535 VSUBS 0.006733f
C632 B.n536 VSUBS 0.006733f
C633 B.n537 VSUBS 0.006733f
C634 B.n538 VSUBS 0.006733f
C635 B.n539 VSUBS 0.006733f
C636 B.n540 VSUBS 0.006733f
C637 B.n541 VSUBS 0.006733f
C638 B.n542 VSUBS 0.005446f
C639 B.n543 VSUBS 0.006733f
C640 B.n544 VSUBS 0.006733f
C641 B.n545 VSUBS 0.004654f
C642 B.n546 VSUBS 0.006733f
C643 B.n547 VSUBS 0.006733f
C644 B.n548 VSUBS 0.006733f
C645 B.n549 VSUBS 0.006733f
C646 B.n550 VSUBS 0.006733f
C647 B.n551 VSUBS 0.006733f
C648 B.n552 VSUBS 0.006733f
C649 B.n553 VSUBS 0.006733f
C650 B.n554 VSUBS 0.006733f
C651 B.n555 VSUBS 0.006733f
C652 B.n556 VSUBS 0.006733f
C653 B.n557 VSUBS 0.006733f
C654 B.n558 VSUBS 0.006733f
C655 B.n559 VSUBS 0.006733f
C656 B.n560 VSUBS 0.006733f
C657 B.n561 VSUBS 0.006733f
C658 B.n562 VSUBS 0.006733f
C659 B.n563 VSUBS 0.006733f
C660 B.n564 VSUBS 0.006733f
C661 B.n565 VSUBS 0.006733f
C662 B.n566 VSUBS 0.006733f
C663 B.n567 VSUBS 0.006733f
C664 B.n568 VSUBS 0.006733f
C665 B.n569 VSUBS 0.006733f
C666 B.n570 VSUBS 0.006733f
C667 B.n571 VSUBS 0.006733f
C668 B.n572 VSUBS 0.006733f
C669 B.n573 VSUBS 0.006733f
C670 B.n574 VSUBS 0.006733f
C671 B.n575 VSUBS 0.006733f
C672 B.n576 VSUBS 0.006733f
C673 B.n577 VSUBS 0.006733f
C674 B.n578 VSUBS 0.006733f
C675 B.n579 VSUBS 0.006733f
C676 B.n580 VSUBS 0.006733f
C677 B.n581 VSUBS 0.006733f
C678 B.n582 VSUBS 0.006733f
C679 B.n583 VSUBS 0.006733f
C680 B.n584 VSUBS 0.006733f
C681 B.n585 VSUBS 0.006733f
C682 B.n586 VSUBS 0.006733f
C683 B.n587 VSUBS 0.006733f
C684 B.n588 VSUBS 0.006733f
C685 B.n589 VSUBS 0.006733f
C686 B.n590 VSUBS 0.006733f
C687 B.n591 VSUBS 0.006733f
C688 B.n592 VSUBS 0.006733f
C689 B.n593 VSUBS 0.006733f
C690 B.n594 VSUBS 0.006733f
C691 B.n595 VSUBS 0.006733f
C692 B.n596 VSUBS 0.006733f
C693 B.n597 VSUBS 0.006733f
C694 B.n598 VSUBS 0.006733f
C695 B.n599 VSUBS 0.006733f
C696 B.n600 VSUBS 0.006733f
C697 B.n601 VSUBS 0.015597f
C698 B.n602 VSUBS 0.015597f
C699 B.n603 VSUBS 0.015297f
C700 B.n604 VSUBS 0.006733f
C701 B.n605 VSUBS 0.006733f
C702 B.n606 VSUBS 0.006733f
C703 B.n607 VSUBS 0.006733f
C704 B.n608 VSUBS 0.006733f
C705 B.n609 VSUBS 0.006733f
C706 B.n610 VSUBS 0.006733f
C707 B.n611 VSUBS 0.006733f
C708 B.n612 VSUBS 0.006733f
C709 B.n613 VSUBS 0.006733f
C710 B.n614 VSUBS 0.006733f
C711 B.n615 VSUBS 0.006733f
C712 B.n616 VSUBS 0.006733f
C713 B.n617 VSUBS 0.006733f
C714 B.n618 VSUBS 0.006733f
C715 B.n619 VSUBS 0.006733f
C716 B.n620 VSUBS 0.006733f
C717 B.n621 VSUBS 0.006733f
C718 B.n622 VSUBS 0.006733f
C719 B.n623 VSUBS 0.006733f
C720 B.n624 VSUBS 0.006733f
C721 B.n625 VSUBS 0.006733f
C722 B.n626 VSUBS 0.006733f
C723 B.n627 VSUBS 0.006733f
C724 B.n628 VSUBS 0.006733f
C725 B.n629 VSUBS 0.006733f
C726 B.n630 VSUBS 0.006733f
C727 B.n631 VSUBS 0.006733f
C728 B.n632 VSUBS 0.006733f
C729 B.n633 VSUBS 0.006733f
C730 B.n634 VSUBS 0.006733f
C731 B.n635 VSUBS 0.006733f
C732 B.n636 VSUBS 0.006733f
C733 B.n637 VSUBS 0.006733f
C734 B.n638 VSUBS 0.006733f
C735 B.n639 VSUBS 0.006733f
C736 B.n640 VSUBS 0.006733f
C737 B.n641 VSUBS 0.006733f
C738 B.n642 VSUBS 0.006733f
C739 B.n643 VSUBS 0.006733f
C740 B.n644 VSUBS 0.006733f
C741 B.n645 VSUBS 0.006733f
C742 B.n646 VSUBS 0.006733f
C743 B.n647 VSUBS 0.006733f
C744 B.n648 VSUBS 0.006733f
C745 B.n649 VSUBS 0.006733f
C746 B.n650 VSUBS 0.006733f
C747 B.n651 VSUBS 0.006733f
C748 B.n652 VSUBS 0.006733f
C749 B.n653 VSUBS 0.006733f
C750 B.n654 VSUBS 0.006733f
C751 B.n655 VSUBS 0.006733f
C752 B.n656 VSUBS 0.006733f
C753 B.n657 VSUBS 0.006733f
C754 B.n658 VSUBS 0.006733f
C755 B.n659 VSUBS 0.015247f
.ends

