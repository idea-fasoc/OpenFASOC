* NGSPICE file created from diff_pair_sample_0407.ext - technology: sky130A

.subckt diff_pair_sample_0407 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=3.24225 ps=19.98 w=19.65 l=0.66
X1 VDD2.t4 VN.t1 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=7.6635 ps=40.08 w=19.65 l=0.66
X2 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=7.6635 ps=40.08 w=19.65 l=0.66
X3 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=3.24225 ps=19.98 w=19.65 l=0.66
X4 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=0 ps=0 w=19.65 l=0.66
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=0 ps=0 w=19.65 l=0.66
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=0 ps=0 w=19.65 l=0.66
X7 VTAIL.t3 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=3.24225 ps=19.98 w=19.65 l=0.66
X8 VTAIL.t0 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=3.24225 ps=19.98 w=19.65 l=0.66
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=0 ps=0 w=19.65 l=0.66
X10 VDD2.t2 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=7.6635 ps=40.08 w=19.65 l=0.66
X11 VTAIL.t8 VN.t4 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=3.24225 ps=19.98 w=19.65 l=0.66
X12 VDD2.t0 VN.t5 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=3.24225 ps=19.98 w=19.65 l=0.66
X13 VDD1.t2 VP.t3 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6635 pd=40.08 as=3.24225 ps=19.98 w=19.65 l=0.66
X14 VTAIL.t10 VP.t4 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=3.24225 ps=19.98 w=19.65 l=0.66
X15 VDD1.t0 VP.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=3.24225 pd=19.98 as=7.6635 ps=40.08 w=19.65 l=0.66
R0 VN.n1 VN.t0 798.202
R1 VN.n7 VN.t3 798.202
R2 VN.n2 VN.t2 777.409
R3 VN.n4 VN.t1 777.409
R4 VN.n8 VN.t4 777.409
R5 VN.n10 VN.t5 777.409
R6 VN.n5 VN.n4 161.3
R7 VN.n11 VN.n10 161.3
R8 VN.n9 VN.n6 161.3
R9 VN.n3 VN.n0 161.3
R10 VN VN.n11 47.1804
R11 VN.n7 VN.n6 44.8515
R12 VN.n1 VN.n0 44.8515
R13 VN.n3 VN.n2 24.8308
R14 VN.n9 VN.n8 24.8308
R15 VN.n4 VN.n3 23.3702
R16 VN.n10 VN.n9 23.3702
R17 VN.n2 VN.n1 21.148
R18 VN.n8 VN.n7 21.148
R19 VN.n11 VN.n6 0.189894
R20 VN.n5 VN.n0 0.189894
R21 VN VN.n5 0.0516364
R22 VTAIL.n442 VTAIL.n338 289.615
R23 VTAIL.n106 VTAIL.n2 289.615
R24 VTAIL.n332 VTAIL.n228 289.615
R25 VTAIL.n220 VTAIL.n116 289.615
R26 VTAIL.n375 VTAIL.n374 185
R27 VTAIL.n377 VTAIL.n376 185
R28 VTAIL.n370 VTAIL.n369 185
R29 VTAIL.n383 VTAIL.n382 185
R30 VTAIL.n385 VTAIL.n384 185
R31 VTAIL.n366 VTAIL.n365 185
R32 VTAIL.n391 VTAIL.n390 185
R33 VTAIL.n393 VTAIL.n392 185
R34 VTAIL.n362 VTAIL.n361 185
R35 VTAIL.n399 VTAIL.n398 185
R36 VTAIL.n401 VTAIL.n400 185
R37 VTAIL.n358 VTAIL.n357 185
R38 VTAIL.n407 VTAIL.n406 185
R39 VTAIL.n409 VTAIL.n408 185
R40 VTAIL.n354 VTAIL.n353 185
R41 VTAIL.n416 VTAIL.n415 185
R42 VTAIL.n417 VTAIL.n352 185
R43 VTAIL.n419 VTAIL.n418 185
R44 VTAIL.n350 VTAIL.n349 185
R45 VTAIL.n425 VTAIL.n424 185
R46 VTAIL.n427 VTAIL.n426 185
R47 VTAIL.n346 VTAIL.n345 185
R48 VTAIL.n433 VTAIL.n432 185
R49 VTAIL.n435 VTAIL.n434 185
R50 VTAIL.n342 VTAIL.n341 185
R51 VTAIL.n441 VTAIL.n440 185
R52 VTAIL.n443 VTAIL.n442 185
R53 VTAIL.n39 VTAIL.n38 185
R54 VTAIL.n41 VTAIL.n40 185
R55 VTAIL.n34 VTAIL.n33 185
R56 VTAIL.n47 VTAIL.n46 185
R57 VTAIL.n49 VTAIL.n48 185
R58 VTAIL.n30 VTAIL.n29 185
R59 VTAIL.n55 VTAIL.n54 185
R60 VTAIL.n57 VTAIL.n56 185
R61 VTAIL.n26 VTAIL.n25 185
R62 VTAIL.n63 VTAIL.n62 185
R63 VTAIL.n65 VTAIL.n64 185
R64 VTAIL.n22 VTAIL.n21 185
R65 VTAIL.n71 VTAIL.n70 185
R66 VTAIL.n73 VTAIL.n72 185
R67 VTAIL.n18 VTAIL.n17 185
R68 VTAIL.n80 VTAIL.n79 185
R69 VTAIL.n81 VTAIL.n16 185
R70 VTAIL.n83 VTAIL.n82 185
R71 VTAIL.n14 VTAIL.n13 185
R72 VTAIL.n89 VTAIL.n88 185
R73 VTAIL.n91 VTAIL.n90 185
R74 VTAIL.n10 VTAIL.n9 185
R75 VTAIL.n97 VTAIL.n96 185
R76 VTAIL.n99 VTAIL.n98 185
R77 VTAIL.n6 VTAIL.n5 185
R78 VTAIL.n105 VTAIL.n104 185
R79 VTAIL.n107 VTAIL.n106 185
R80 VTAIL.n333 VTAIL.n332 185
R81 VTAIL.n331 VTAIL.n330 185
R82 VTAIL.n232 VTAIL.n231 185
R83 VTAIL.n325 VTAIL.n324 185
R84 VTAIL.n323 VTAIL.n322 185
R85 VTAIL.n236 VTAIL.n235 185
R86 VTAIL.n317 VTAIL.n316 185
R87 VTAIL.n315 VTAIL.n314 185
R88 VTAIL.n240 VTAIL.n239 185
R89 VTAIL.n244 VTAIL.n242 185
R90 VTAIL.n309 VTAIL.n308 185
R91 VTAIL.n307 VTAIL.n306 185
R92 VTAIL.n246 VTAIL.n245 185
R93 VTAIL.n301 VTAIL.n300 185
R94 VTAIL.n299 VTAIL.n298 185
R95 VTAIL.n250 VTAIL.n249 185
R96 VTAIL.n293 VTAIL.n292 185
R97 VTAIL.n291 VTAIL.n290 185
R98 VTAIL.n254 VTAIL.n253 185
R99 VTAIL.n285 VTAIL.n284 185
R100 VTAIL.n283 VTAIL.n282 185
R101 VTAIL.n258 VTAIL.n257 185
R102 VTAIL.n277 VTAIL.n276 185
R103 VTAIL.n275 VTAIL.n274 185
R104 VTAIL.n262 VTAIL.n261 185
R105 VTAIL.n269 VTAIL.n268 185
R106 VTAIL.n267 VTAIL.n266 185
R107 VTAIL.n221 VTAIL.n220 185
R108 VTAIL.n219 VTAIL.n218 185
R109 VTAIL.n120 VTAIL.n119 185
R110 VTAIL.n213 VTAIL.n212 185
R111 VTAIL.n211 VTAIL.n210 185
R112 VTAIL.n124 VTAIL.n123 185
R113 VTAIL.n205 VTAIL.n204 185
R114 VTAIL.n203 VTAIL.n202 185
R115 VTAIL.n128 VTAIL.n127 185
R116 VTAIL.n132 VTAIL.n130 185
R117 VTAIL.n197 VTAIL.n196 185
R118 VTAIL.n195 VTAIL.n194 185
R119 VTAIL.n134 VTAIL.n133 185
R120 VTAIL.n189 VTAIL.n188 185
R121 VTAIL.n187 VTAIL.n186 185
R122 VTAIL.n138 VTAIL.n137 185
R123 VTAIL.n181 VTAIL.n180 185
R124 VTAIL.n179 VTAIL.n178 185
R125 VTAIL.n142 VTAIL.n141 185
R126 VTAIL.n173 VTAIL.n172 185
R127 VTAIL.n171 VTAIL.n170 185
R128 VTAIL.n146 VTAIL.n145 185
R129 VTAIL.n165 VTAIL.n164 185
R130 VTAIL.n163 VTAIL.n162 185
R131 VTAIL.n150 VTAIL.n149 185
R132 VTAIL.n157 VTAIL.n156 185
R133 VTAIL.n155 VTAIL.n154 185
R134 VTAIL.n373 VTAIL.t7 147.659
R135 VTAIL.n37 VTAIL.t2 147.659
R136 VTAIL.n265 VTAIL.t9 147.659
R137 VTAIL.n153 VTAIL.t6 147.659
R138 VTAIL.n376 VTAIL.n375 104.615
R139 VTAIL.n376 VTAIL.n369 104.615
R140 VTAIL.n383 VTAIL.n369 104.615
R141 VTAIL.n384 VTAIL.n383 104.615
R142 VTAIL.n384 VTAIL.n365 104.615
R143 VTAIL.n391 VTAIL.n365 104.615
R144 VTAIL.n392 VTAIL.n391 104.615
R145 VTAIL.n392 VTAIL.n361 104.615
R146 VTAIL.n399 VTAIL.n361 104.615
R147 VTAIL.n400 VTAIL.n399 104.615
R148 VTAIL.n400 VTAIL.n357 104.615
R149 VTAIL.n407 VTAIL.n357 104.615
R150 VTAIL.n408 VTAIL.n407 104.615
R151 VTAIL.n408 VTAIL.n353 104.615
R152 VTAIL.n416 VTAIL.n353 104.615
R153 VTAIL.n417 VTAIL.n416 104.615
R154 VTAIL.n418 VTAIL.n417 104.615
R155 VTAIL.n418 VTAIL.n349 104.615
R156 VTAIL.n425 VTAIL.n349 104.615
R157 VTAIL.n426 VTAIL.n425 104.615
R158 VTAIL.n426 VTAIL.n345 104.615
R159 VTAIL.n433 VTAIL.n345 104.615
R160 VTAIL.n434 VTAIL.n433 104.615
R161 VTAIL.n434 VTAIL.n341 104.615
R162 VTAIL.n441 VTAIL.n341 104.615
R163 VTAIL.n442 VTAIL.n441 104.615
R164 VTAIL.n40 VTAIL.n39 104.615
R165 VTAIL.n40 VTAIL.n33 104.615
R166 VTAIL.n47 VTAIL.n33 104.615
R167 VTAIL.n48 VTAIL.n47 104.615
R168 VTAIL.n48 VTAIL.n29 104.615
R169 VTAIL.n55 VTAIL.n29 104.615
R170 VTAIL.n56 VTAIL.n55 104.615
R171 VTAIL.n56 VTAIL.n25 104.615
R172 VTAIL.n63 VTAIL.n25 104.615
R173 VTAIL.n64 VTAIL.n63 104.615
R174 VTAIL.n64 VTAIL.n21 104.615
R175 VTAIL.n71 VTAIL.n21 104.615
R176 VTAIL.n72 VTAIL.n71 104.615
R177 VTAIL.n72 VTAIL.n17 104.615
R178 VTAIL.n80 VTAIL.n17 104.615
R179 VTAIL.n81 VTAIL.n80 104.615
R180 VTAIL.n82 VTAIL.n81 104.615
R181 VTAIL.n82 VTAIL.n13 104.615
R182 VTAIL.n89 VTAIL.n13 104.615
R183 VTAIL.n90 VTAIL.n89 104.615
R184 VTAIL.n90 VTAIL.n9 104.615
R185 VTAIL.n97 VTAIL.n9 104.615
R186 VTAIL.n98 VTAIL.n97 104.615
R187 VTAIL.n98 VTAIL.n5 104.615
R188 VTAIL.n105 VTAIL.n5 104.615
R189 VTAIL.n106 VTAIL.n105 104.615
R190 VTAIL.n332 VTAIL.n331 104.615
R191 VTAIL.n331 VTAIL.n231 104.615
R192 VTAIL.n324 VTAIL.n231 104.615
R193 VTAIL.n324 VTAIL.n323 104.615
R194 VTAIL.n323 VTAIL.n235 104.615
R195 VTAIL.n316 VTAIL.n235 104.615
R196 VTAIL.n316 VTAIL.n315 104.615
R197 VTAIL.n315 VTAIL.n239 104.615
R198 VTAIL.n244 VTAIL.n239 104.615
R199 VTAIL.n308 VTAIL.n244 104.615
R200 VTAIL.n308 VTAIL.n307 104.615
R201 VTAIL.n307 VTAIL.n245 104.615
R202 VTAIL.n300 VTAIL.n245 104.615
R203 VTAIL.n300 VTAIL.n299 104.615
R204 VTAIL.n299 VTAIL.n249 104.615
R205 VTAIL.n292 VTAIL.n249 104.615
R206 VTAIL.n292 VTAIL.n291 104.615
R207 VTAIL.n291 VTAIL.n253 104.615
R208 VTAIL.n284 VTAIL.n253 104.615
R209 VTAIL.n284 VTAIL.n283 104.615
R210 VTAIL.n283 VTAIL.n257 104.615
R211 VTAIL.n276 VTAIL.n257 104.615
R212 VTAIL.n276 VTAIL.n275 104.615
R213 VTAIL.n275 VTAIL.n261 104.615
R214 VTAIL.n268 VTAIL.n261 104.615
R215 VTAIL.n268 VTAIL.n267 104.615
R216 VTAIL.n220 VTAIL.n219 104.615
R217 VTAIL.n219 VTAIL.n119 104.615
R218 VTAIL.n212 VTAIL.n119 104.615
R219 VTAIL.n212 VTAIL.n211 104.615
R220 VTAIL.n211 VTAIL.n123 104.615
R221 VTAIL.n204 VTAIL.n123 104.615
R222 VTAIL.n204 VTAIL.n203 104.615
R223 VTAIL.n203 VTAIL.n127 104.615
R224 VTAIL.n132 VTAIL.n127 104.615
R225 VTAIL.n196 VTAIL.n132 104.615
R226 VTAIL.n196 VTAIL.n195 104.615
R227 VTAIL.n195 VTAIL.n133 104.615
R228 VTAIL.n188 VTAIL.n133 104.615
R229 VTAIL.n188 VTAIL.n187 104.615
R230 VTAIL.n187 VTAIL.n137 104.615
R231 VTAIL.n180 VTAIL.n137 104.615
R232 VTAIL.n180 VTAIL.n179 104.615
R233 VTAIL.n179 VTAIL.n141 104.615
R234 VTAIL.n172 VTAIL.n141 104.615
R235 VTAIL.n172 VTAIL.n171 104.615
R236 VTAIL.n171 VTAIL.n145 104.615
R237 VTAIL.n164 VTAIL.n145 104.615
R238 VTAIL.n164 VTAIL.n163 104.615
R239 VTAIL.n163 VTAIL.n149 104.615
R240 VTAIL.n156 VTAIL.n149 104.615
R241 VTAIL.n156 VTAIL.n155 104.615
R242 VTAIL.n375 VTAIL.t7 52.3082
R243 VTAIL.n39 VTAIL.t2 52.3082
R244 VTAIL.n267 VTAIL.t9 52.3082
R245 VTAIL.n155 VTAIL.t6 52.3082
R246 VTAIL.n227 VTAIL.n226 43.3415
R247 VTAIL.n115 VTAIL.n114 43.3415
R248 VTAIL.n1 VTAIL.n0 43.3414
R249 VTAIL.n113 VTAIL.n112 43.3414
R250 VTAIL.n447 VTAIL.n446 31.6035
R251 VTAIL.n111 VTAIL.n110 31.6035
R252 VTAIL.n337 VTAIL.n336 31.6035
R253 VTAIL.n225 VTAIL.n224 31.6035
R254 VTAIL.n115 VTAIL.n113 31.0134
R255 VTAIL.n447 VTAIL.n337 30.16
R256 VTAIL.n374 VTAIL.n373 15.6677
R257 VTAIL.n38 VTAIL.n37 15.6677
R258 VTAIL.n266 VTAIL.n265 15.6677
R259 VTAIL.n154 VTAIL.n153 15.6677
R260 VTAIL.n419 VTAIL.n350 13.1884
R261 VTAIL.n83 VTAIL.n14 13.1884
R262 VTAIL.n242 VTAIL.n240 13.1884
R263 VTAIL.n130 VTAIL.n128 13.1884
R264 VTAIL.n377 VTAIL.n372 12.8005
R265 VTAIL.n420 VTAIL.n352 12.8005
R266 VTAIL.n424 VTAIL.n423 12.8005
R267 VTAIL.n41 VTAIL.n36 12.8005
R268 VTAIL.n84 VTAIL.n16 12.8005
R269 VTAIL.n88 VTAIL.n87 12.8005
R270 VTAIL.n314 VTAIL.n313 12.8005
R271 VTAIL.n310 VTAIL.n309 12.8005
R272 VTAIL.n269 VTAIL.n264 12.8005
R273 VTAIL.n202 VTAIL.n201 12.8005
R274 VTAIL.n198 VTAIL.n197 12.8005
R275 VTAIL.n157 VTAIL.n152 12.8005
R276 VTAIL.n378 VTAIL.n370 12.0247
R277 VTAIL.n415 VTAIL.n414 12.0247
R278 VTAIL.n427 VTAIL.n348 12.0247
R279 VTAIL.n42 VTAIL.n34 12.0247
R280 VTAIL.n79 VTAIL.n78 12.0247
R281 VTAIL.n91 VTAIL.n12 12.0247
R282 VTAIL.n317 VTAIL.n238 12.0247
R283 VTAIL.n306 VTAIL.n243 12.0247
R284 VTAIL.n270 VTAIL.n262 12.0247
R285 VTAIL.n205 VTAIL.n126 12.0247
R286 VTAIL.n194 VTAIL.n131 12.0247
R287 VTAIL.n158 VTAIL.n150 12.0247
R288 VTAIL.n382 VTAIL.n381 11.249
R289 VTAIL.n413 VTAIL.n354 11.249
R290 VTAIL.n428 VTAIL.n346 11.249
R291 VTAIL.n46 VTAIL.n45 11.249
R292 VTAIL.n77 VTAIL.n18 11.249
R293 VTAIL.n92 VTAIL.n10 11.249
R294 VTAIL.n318 VTAIL.n236 11.249
R295 VTAIL.n305 VTAIL.n246 11.249
R296 VTAIL.n274 VTAIL.n273 11.249
R297 VTAIL.n206 VTAIL.n124 11.249
R298 VTAIL.n193 VTAIL.n134 11.249
R299 VTAIL.n162 VTAIL.n161 11.249
R300 VTAIL.n385 VTAIL.n368 10.4732
R301 VTAIL.n410 VTAIL.n409 10.4732
R302 VTAIL.n432 VTAIL.n431 10.4732
R303 VTAIL.n49 VTAIL.n32 10.4732
R304 VTAIL.n74 VTAIL.n73 10.4732
R305 VTAIL.n96 VTAIL.n95 10.4732
R306 VTAIL.n322 VTAIL.n321 10.4732
R307 VTAIL.n302 VTAIL.n301 10.4732
R308 VTAIL.n277 VTAIL.n260 10.4732
R309 VTAIL.n210 VTAIL.n209 10.4732
R310 VTAIL.n190 VTAIL.n189 10.4732
R311 VTAIL.n165 VTAIL.n148 10.4732
R312 VTAIL.n386 VTAIL.n366 9.69747
R313 VTAIL.n406 VTAIL.n356 9.69747
R314 VTAIL.n435 VTAIL.n344 9.69747
R315 VTAIL.n50 VTAIL.n30 9.69747
R316 VTAIL.n70 VTAIL.n20 9.69747
R317 VTAIL.n99 VTAIL.n8 9.69747
R318 VTAIL.n325 VTAIL.n234 9.69747
R319 VTAIL.n298 VTAIL.n248 9.69747
R320 VTAIL.n278 VTAIL.n258 9.69747
R321 VTAIL.n213 VTAIL.n122 9.69747
R322 VTAIL.n186 VTAIL.n136 9.69747
R323 VTAIL.n166 VTAIL.n146 9.69747
R324 VTAIL.n446 VTAIL.n445 9.45567
R325 VTAIL.n110 VTAIL.n109 9.45567
R326 VTAIL.n336 VTAIL.n335 9.45567
R327 VTAIL.n224 VTAIL.n223 9.45567
R328 VTAIL.n445 VTAIL.n444 9.3005
R329 VTAIL.n439 VTAIL.n438 9.3005
R330 VTAIL.n437 VTAIL.n436 9.3005
R331 VTAIL.n344 VTAIL.n343 9.3005
R332 VTAIL.n431 VTAIL.n430 9.3005
R333 VTAIL.n429 VTAIL.n428 9.3005
R334 VTAIL.n348 VTAIL.n347 9.3005
R335 VTAIL.n423 VTAIL.n422 9.3005
R336 VTAIL.n395 VTAIL.n394 9.3005
R337 VTAIL.n364 VTAIL.n363 9.3005
R338 VTAIL.n389 VTAIL.n388 9.3005
R339 VTAIL.n387 VTAIL.n386 9.3005
R340 VTAIL.n368 VTAIL.n367 9.3005
R341 VTAIL.n381 VTAIL.n380 9.3005
R342 VTAIL.n379 VTAIL.n378 9.3005
R343 VTAIL.n372 VTAIL.n371 9.3005
R344 VTAIL.n397 VTAIL.n396 9.3005
R345 VTAIL.n360 VTAIL.n359 9.3005
R346 VTAIL.n403 VTAIL.n402 9.3005
R347 VTAIL.n405 VTAIL.n404 9.3005
R348 VTAIL.n356 VTAIL.n355 9.3005
R349 VTAIL.n411 VTAIL.n410 9.3005
R350 VTAIL.n413 VTAIL.n412 9.3005
R351 VTAIL.n414 VTAIL.n351 9.3005
R352 VTAIL.n421 VTAIL.n420 9.3005
R353 VTAIL.n340 VTAIL.n339 9.3005
R354 VTAIL.n109 VTAIL.n108 9.3005
R355 VTAIL.n103 VTAIL.n102 9.3005
R356 VTAIL.n101 VTAIL.n100 9.3005
R357 VTAIL.n8 VTAIL.n7 9.3005
R358 VTAIL.n95 VTAIL.n94 9.3005
R359 VTAIL.n93 VTAIL.n92 9.3005
R360 VTAIL.n12 VTAIL.n11 9.3005
R361 VTAIL.n87 VTAIL.n86 9.3005
R362 VTAIL.n59 VTAIL.n58 9.3005
R363 VTAIL.n28 VTAIL.n27 9.3005
R364 VTAIL.n53 VTAIL.n52 9.3005
R365 VTAIL.n51 VTAIL.n50 9.3005
R366 VTAIL.n32 VTAIL.n31 9.3005
R367 VTAIL.n45 VTAIL.n44 9.3005
R368 VTAIL.n43 VTAIL.n42 9.3005
R369 VTAIL.n36 VTAIL.n35 9.3005
R370 VTAIL.n61 VTAIL.n60 9.3005
R371 VTAIL.n24 VTAIL.n23 9.3005
R372 VTAIL.n67 VTAIL.n66 9.3005
R373 VTAIL.n69 VTAIL.n68 9.3005
R374 VTAIL.n20 VTAIL.n19 9.3005
R375 VTAIL.n75 VTAIL.n74 9.3005
R376 VTAIL.n77 VTAIL.n76 9.3005
R377 VTAIL.n78 VTAIL.n15 9.3005
R378 VTAIL.n85 VTAIL.n84 9.3005
R379 VTAIL.n4 VTAIL.n3 9.3005
R380 VTAIL.n252 VTAIL.n251 9.3005
R381 VTAIL.n295 VTAIL.n294 9.3005
R382 VTAIL.n297 VTAIL.n296 9.3005
R383 VTAIL.n248 VTAIL.n247 9.3005
R384 VTAIL.n303 VTAIL.n302 9.3005
R385 VTAIL.n305 VTAIL.n304 9.3005
R386 VTAIL.n243 VTAIL.n241 9.3005
R387 VTAIL.n311 VTAIL.n310 9.3005
R388 VTAIL.n335 VTAIL.n334 9.3005
R389 VTAIL.n230 VTAIL.n229 9.3005
R390 VTAIL.n329 VTAIL.n328 9.3005
R391 VTAIL.n327 VTAIL.n326 9.3005
R392 VTAIL.n234 VTAIL.n233 9.3005
R393 VTAIL.n321 VTAIL.n320 9.3005
R394 VTAIL.n319 VTAIL.n318 9.3005
R395 VTAIL.n238 VTAIL.n237 9.3005
R396 VTAIL.n313 VTAIL.n312 9.3005
R397 VTAIL.n289 VTAIL.n288 9.3005
R398 VTAIL.n287 VTAIL.n286 9.3005
R399 VTAIL.n256 VTAIL.n255 9.3005
R400 VTAIL.n281 VTAIL.n280 9.3005
R401 VTAIL.n279 VTAIL.n278 9.3005
R402 VTAIL.n260 VTAIL.n259 9.3005
R403 VTAIL.n273 VTAIL.n272 9.3005
R404 VTAIL.n271 VTAIL.n270 9.3005
R405 VTAIL.n264 VTAIL.n263 9.3005
R406 VTAIL.n140 VTAIL.n139 9.3005
R407 VTAIL.n183 VTAIL.n182 9.3005
R408 VTAIL.n185 VTAIL.n184 9.3005
R409 VTAIL.n136 VTAIL.n135 9.3005
R410 VTAIL.n191 VTAIL.n190 9.3005
R411 VTAIL.n193 VTAIL.n192 9.3005
R412 VTAIL.n131 VTAIL.n129 9.3005
R413 VTAIL.n199 VTAIL.n198 9.3005
R414 VTAIL.n223 VTAIL.n222 9.3005
R415 VTAIL.n118 VTAIL.n117 9.3005
R416 VTAIL.n217 VTAIL.n216 9.3005
R417 VTAIL.n215 VTAIL.n214 9.3005
R418 VTAIL.n122 VTAIL.n121 9.3005
R419 VTAIL.n209 VTAIL.n208 9.3005
R420 VTAIL.n207 VTAIL.n206 9.3005
R421 VTAIL.n126 VTAIL.n125 9.3005
R422 VTAIL.n201 VTAIL.n200 9.3005
R423 VTAIL.n177 VTAIL.n176 9.3005
R424 VTAIL.n175 VTAIL.n174 9.3005
R425 VTAIL.n144 VTAIL.n143 9.3005
R426 VTAIL.n169 VTAIL.n168 9.3005
R427 VTAIL.n167 VTAIL.n166 9.3005
R428 VTAIL.n148 VTAIL.n147 9.3005
R429 VTAIL.n161 VTAIL.n160 9.3005
R430 VTAIL.n159 VTAIL.n158 9.3005
R431 VTAIL.n152 VTAIL.n151 9.3005
R432 VTAIL.n390 VTAIL.n389 8.92171
R433 VTAIL.n405 VTAIL.n358 8.92171
R434 VTAIL.n436 VTAIL.n342 8.92171
R435 VTAIL.n54 VTAIL.n53 8.92171
R436 VTAIL.n69 VTAIL.n22 8.92171
R437 VTAIL.n100 VTAIL.n6 8.92171
R438 VTAIL.n326 VTAIL.n232 8.92171
R439 VTAIL.n297 VTAIL.n250 8.92171
R440 VTAIL.n282 VTAIL.n281 8.92171
R441 VTAIL.n214 VTAIL.n120 8.92171
R442 VTAIL.n185 VTAIL.n138 8.92171
R443 VTAIL.n170 VTAIL.n169 8.92171
R444 VTAIL.n393 VTAIL.n364 8.14595
R445 VTAIL.n402 VTAIL.n401 8.14595
R446 VTAIL.n440 VTAIL.n439 8.14595
R447 VTAIL.n57 VTAIL.n28 8.14595
R448 VTAIL.n66 VTAIL.n65 8.14595
R449 VTAIL.n104 VTAIL.n103 8.14595
R450 VTAIL.n330 VTAIL.n329 8.14595
R451 VTAIL.n294 VTAIL.n293 8.14595
R452 VTAIL.n285 VTAIL.n256 8.14595
R453 VTAIL.n218 VTAIL.n217 8.14595
R454 VTAIL.n182 VTAIL.n181 8.14595
R455 VTAIL.n173 VTAIL.n144 8.14595
R456 VTAIL.n394 VTAIL.n362 7.3702
R457 VTAIL.n398 VTAIL.n360 7.3702
R458 VTAIL.n443 VTAIL.n340 7.3702
R459 VTAIL.n446 VTAIL.n338 7.3702
R460 VTAIL.n58 VTAIL.n26 7.3702
R461 VTAIL.n62 VTAIL.n24 7.3702
R462 VTAIL.n107 VTAIL.n4 7.3702
R463 VTAIL.n110 VTAIL.n2 7.3702
R464 VTAIL.n336 VTAIL.n228 7.3702
R465 VTAIL.n333 VTAIL.n230 7.3702
R466 VTAIL.n290 VTAIL.n252 7.3702
R467 VTAIL.n286 VTAIL.n254 7.3702
R468 VTAIL.n224 VTAIL.n116 7.3702
R469 VTAIL.n221 VTAIL.n118 7.3702
R470 VTAIL.n178 VTAIL.n140 7.3702
R471 VTAIL.n174 VTAIL.n142 7.3702
R472 VTAIL.n397 VTAIL.n362 6.59444
R473 VTAIL.n398 VTAIL.n397 6.59444
R474 VTAIL.n444 VTAIL.n443 6.59444
R475 VTAIL.n444 VTAIL.n338 6.59444
R476 VTAIL.n61 VTAIL.n26 6.59444
R477 VTAIL.n62 VTAIL.n61 6.59444
R478 VTAIL.n108 VTAIL.n107 6.59444
R479 VTAIL.n108 VTAIL.n2 6.59444
R480 VTAIL.n334 VTAIL.n228 6.59444
R481 VTAIL.n334 VTAIL.n333 6.59444
R482 VTAIL.n290 VTAIL.n289 6.59444
R483 VTAIL.n289 VTAIL.n254 6.59444
R484 VTAIL.n222 VTAIL.n116 6.59444
R485 VTAIL.n222 VTAIL.n221 6.59444
R486 VTAIL.n178 VTAIL.n177 6.59444
R487 VTAIL.n177 VTAIL.n142 6.59444
R488 VTAIL.n394 VTAIL.n393 5.81868
R489 VTAIL.n401 VTAIL.n360 5.81868
R490 VTAIL.n440 VTAIL.n340 5.81868
R491 VTAIL.n58 VTAIL.n57 5.81868
R492 VTAIL.n65 VTAIL.n24 5.81868
R493 VTAIL.n104 VTAIL.n4 5.81868
R494 VTAIL.n330 VTAIL.n230 5.81868
R495 VTAIL.n293 VTAIL.n252 5.81868
R496 VTAIL.n286 VTAIL.n285 5.81868
R497 VTAIL.n218 VTAIL.n118 5.81868
R498 VTAIL.n181 VTAIL.n140 5.81868
R499 VTAIL.n174 VTAIL.n173 5.81868
R500 VTAIL.n390 VTAIL.n364 5.04292
R501 VTAIL.n402 VTAIL.n358 5.04292
R502 VTAIL.n439 VTAIL.n342 5.04292
R503 VTAIL.n54 VTAIL.n28 5.04292
R504 VTAIL.n66 VTAIL.n22 5.04292
R505 VTAIL.n103 VTAIL.n6 5.04292
R506 VTAIL.n329 VTAIL.n232 5.04292
R507 VTAIL.n294 VTAIL.n250 5.04292
R508 VTAIL.n282 VTAIL.n256 5.04292
R509 VTAIL.n217 VTAIL.n120 5.04292
R510 VTAIL.n182 VTAIL.n138 5.04292
R511 VTAIL.n170 VTAIL.n144 5.04292
R512 VTAIL.n373 VTAIL.n371 4.38563
R513 VTAIL.n37 VTAIL.n35 4.38563
R514 VTAIL.n265 VTAIL.n263 4.38563
R515 VTAIL.n153 VTAIL.n151 4.38563
R516 VTAIL.n389 VTAIL.n366 4.26717
R517 VTAIL.n406 VTAIL.n405 4.26717
R518 VTAIL.n436 VTAIL.n435 4.26717
R519 VTAIL.n53 VTAIL.n30 4.26717
R520 VTAIL.n70 VTAIL.n69 4.26717
R521 VTAIL.n100 VTAIL.n99 4.26717
R522 VTAIL.n326 VTAIL.n325 4.26717
R523 VTAIL.n298 VTAIL.n297 4.26717
R524 VTAIL.n281 VTAIL.n258 4.26717
R525 VTAIL.n214 VTAIL.n213 4.26717
R526 VTAIL.n186 VTAIL.n185 4.26717
R527 VTAIL.n169 VTAIL.n146 4.26717
R528 VTAIL.n386 VTAIL.n385 3.49141
R529 VTAIL.n409 VTAIL.n356 3.49141
R530 VTAIL.n432 VTAIL.n344 3.49141
R531 VTAIL.n50 VTAIL.n49 3.49141
R532 VTAIL.n73 VTAIL.n20 3.49141
R533 VTAIL.n96 VTAIL.n8 3.49141
R534 VTAIL.n322 VTAIL.n234 3.49141
R535 VTAIL.n301 VTAIL.n248 3.49141
R536 VTAIL.n278 VTAIL.n277 3.49141
R537 VTAIL.n210 VTAIL.n122 3.49141
R538 VTAIL.n189 VTAIL.n136 3.49141
R539 VTAIL.n166 VTAIL.n165 3.49141
R540 VTAIL.n382 VTAIL.n368 2.71565
R541 VTAIL.n410 VTAIL.n354 2.71565
R542 VTAIL.n431 VTAIL.n346 2.71565
R543 VTAIL.n46 VTAIL.n32 2.71565
R544 VTAIL.n74 VTAIL.n18 2.71565
R545 VTAIL.n95 VTAIL.n10 2.71565
R546 VTAIL.n321 VTAIL.n236 2.71565
R547 VTAIL.n302 VTAIL.n246 2.71565
R548 VTAIL.n274 VTAIL.n260 2.71565
R549 VTAIL.n209 VTAIL.n124 2.71565
R550 VTAIL.n190 VTAIL.n134 2.71565
R551 VTAIL.n162 VTAIL.n148 2.71565
R552 VTAIL.n381 VTAIL.n370 1.93989
R553 VTAIL.n415 VTAIL.n413 1.93989
R554 VTAIL.n428 VTAIL.n427 1.93989
R555 VTAIL.n45 VTAIL.n34 1.93989
R556 VTAIL.n79 VTAIL.n77 1.93989
R557 VTAIL.n92 VTAIL.n91 1.93989
R558 VTAIL.n318 VTAIL.n317 1.93989
R559 VTAIL.n306 VTAIL.n305 1.93989
R560 VTAIL.n273 VTAIL.n262 1.93989
R561 VTAIL.n206 VTAIL.n205 1.93989
R562 VTAIL.n194 VTAIL.n193 1.93989
R563 VTAIL.n161 VTAIL.n150 1.93989
R564 VTAIL.n378 VTAIL.n377 1.16414
R565 VTAIL.n414 VTAIL.n352 1.16414
R566 VTAIL.n424 VTAIL.n348 1.16414
R567 VTAIL.n42 VTAIL.n41 1.16414
R568 VTAIL.n78 VTAIL.n16 1.16414
R569 VTAIL.n88 VTAIL.n12 1.16414
R570 VTAIL.n314 VTAIL.n238 1.16414
R571 VTAIL.n309 VTAIL.n243 1.16414
R572 VTAIL.n270 VTAIL.n269 1.16414
R573 VTAIL.n202 VTAIL.n126 1.16414
R574 VTAIL.n197 VTAIL.n131 1.16414
R575 VTAIL.n158 VTAIL.n157 1.16414
R576 VTAIL.n0 VTAIL.t4 1.00813
R577 VTAIL.n0 VTAIL.t3 1.00813
R578 VTAIL.n112 VTAIL.t1 1.00813
R579 VTAIL.n112 VTAIL.t0 1.00813
R580 VTAIL.n226 VTAIL.t11 1.00813
R581 VTAIL.n226 VTAIL.t10 1.00813
R582 VTAIL.n114 VTAIL.t5 1.00813
R583 VTAIL.n114 VTAIL.t8 1.00813
R584 VTAIL.n227 VTAIL.n225 0.897052
R585 VTAIL.n111 VTAIL.n1 0.897052
R586 VTAIL.n225 VTAIL.n115 0.853948
R587 VTAIL.n337 VTAIL.n227 0.853948
R588 VTAIL.n113 VTAIL.n111 0.853948
R589 VTAIL VTAIL.n447 0.582397
R590 VTAIL.n374 VTAIL.n372 0.388379
R591 VTAIL.n420 VTAIL.n419 0.388379
R592 VTAIL.n423 VTAIL.n350 0.388379
R593 VTAIL.n38 VTAIL.n36 0.388379
R594 VTAIL.n84 VTAIL.n83 0.388379
R595 VTAIL.n87 VTAIL.n14 0.388379
R596 VTAIL.n313 VTAIL.n240 0.388379
R597 VTAIL.n310 VTAIL.n242 0.388379
R598 VTAIL.n266 VTAIL.n264 0.388379
R599 VTAIL.n201 VTAIL.n128 0.388379
R600 VTAIL.n198 VTAIL.n130 0.388379
R601 VTAIL.n154 VTAIL.n152 0.388379
R602 VTAIL VTAIL.n1 0.272052
R603 VTAIL.n379 VTAIL.n371 0.155672
R604 VTAIL.n380 VTAIL.n379 0.155672
R605 VTAIL.n380 VTAIL.n367 0.155672
R606 VTAIL.n387 VTAIL.n367 0.155672
R607 VTAIL.n388 VTAIL.n387 0.155672
R608 VTAIL.n388 VTAIL.n363 0.155672
R609 VTAIL.n395 VTAIL.n363 0.155672
R610 VTAIL.n396 VTAIL.n395 0.155672
R611 VTAIL.n396 VTAIL.n359 0.155672
R612 VTAIL.n403 VTAIL.n359 0.155672
R613 VTAIL.n404 VTAIL.n403 0.155672
R614 VTAIL.n404 VTAIL.n355 0.155672
R615 VTAIL.n411 VTAIL.n355 0.155672
R616 VTAIL.n412 VTAIL.n411 0.155672
R617 VTAIL.n412 VTAIL.n351 0.155672
R618 VTAIL.n421 VTAIL.n351 0.155672
R619 VTAIL.n422 VTAIL.n421 0.155672
R620 VTAIL.n422 VTAIL.n347 0.155672
R621 VTAIL.n429 VTAIL.n347 0.155672
R622 VTAIL.n430 VTAIL.n429 0.155672
R623 VTAIL.n430 VTAIL.n343 0.155672
R624 VTAIL.n437 VTAIL.n343 0.155672
R625 VTAIL.n438 VTAIL.n437 0.155672
R626 VTAIL.n438 VTAIL.n339 0.155672
R627 VTAIL.n445 VTAIL.n339 0.155672
R628 VTAIL.n43 VTAIL.n35 0.155672
R629 VTAIL.n44 VTAIL.n43 0.155672
R630 VTAIL.n44 VTAIL.n31 0.155672
R631 VTAIL.n51 VTAIL.n31 0.155672
R632 VTAIL.n52 VTAIL.n51 0.155672
R633 VTAIL.n52 VTAIL.n27 0.155672
R634 VTAIL.n59 VTAIL.n27 0.155672
R635 VTAIL.n60 VTAIL.n59 0.155672
R636 VTAIL.n60 VTAIL.n23 0.155672
R637 VTAIL.n67 VTAIL.n23 0.155672
R638 VTAIL.n68 VTAIL.n67 0.155672
R639 VTAIL.n68 VTAIL.n19 0.155672
R640 VTAIL.n75 VTAIL.n19 0.155672
R641 VTAIL.n76 VTAIL.n75 0.155672
R642 VTAIL.n76 VTAIL.n15 0.155672
R643 VTAIL.n85 VTAIL.n15 0.155672
R644 VTAIL.n86 VTAIL.n85 0.155672
R645 VTAIL.n86 VTAIL.n11 0.155672
R646 VTAIL.n93 VTAIL.n11 0.155672
R647 VTAIL.n94 VTAIL.n93 0.155672
R648 VTAIL.n94 VTAIL.n7 0.155672
R649 VTAIL.n101 VTAIL.n7 0.155672
R650 VTAIL.n102 VTAIL.n101 0.155672
R651 VTAIL.n102 VTAIL.n3 0.155672
R652 VTAIL.n109 VTAIL.n3 0.155672
R653 VTAIL.n335 VTAIL.n229 0.155672
R654 VTAIL.n328 VTAIL.n229 0.155672
R655 VTAIL.n328 VTAIL.n327 0.155672
R656 VTAIL.n327 VTAIL.n233 0.155672
R657 VTAIL.n320 VTAIL.n233 0.155672
R658 VTAIL.n320 VTAIL.n319 0.155672
R659 VTAIL.n319 VTAIL.n237 0.155672
R660 VTAIL.n312 VTAIL.n237 0.155672
R661 VTAIL.n312 VTAIL.n311 0.155672
R662 VTAIL.n311 VTAIL.n241 0.155672
R663 VTAIL.n304 VTAIL.n241 0.155672
R664 VTAIL.n304 VTAIL.n303 0.155672
R665 VTAIL.n303 VTAIL.n247 0.155672
R666 VTAIL.n296 VTAIL.n247 0.155672
R667 VTAIL.n296 VTAIL.n295 0.155672
R668 VTAIL.n295 VTAIL.n251 0.155672
R669 VTAIL.n288 VTAIL.n251 0.155672
R670 VTAIL.n288 VTAIL.n287 0.155672
R671 VTAIL.n287 VTAIL.n255 0.155672
R672 VTAIL.n280 VTAIL.n255 0.155672
R673 VTAIL.n280 VTAIL.n279 0.155672
R674 VTAIL.n279 VTAIL.n259 0.155672
R675 VTAIL.n272 VTAIL.n259 0.155672
R676 VTAIL.n272 VTAIL.n271 0.155672
R677 VTAIL.n271 VTAIL.n263 0.155672
R678 VTAIL.n223 VTAIL.n117 0.155672
R679 VTAIL.n216 VTAIL.n117 0.155672
R680 VTAIL.n216 VTAIL.n215 0.155672
R681 VTAIL.n215 VTAIL.n121 0.155672
R682 VTAIL.n208 VTAIL.n121 0.155672
R683 VTAIL.n208 VTAIL.n207 0.155672
R684 VTAIL.n207 VTAIL.n125 0.155672
R685 VTAIL.n200 VTAIL.n125 0.155672
R686 VTAIL.n200 VTAIL.n199 0.155672
R687 VTAIL.n199 VTAIL.n129 0.155672
R688 VTAIL.n192 VTAIL.n129 0.155672
R689 VTAIL.n192 VTAIL.n191 0.155672
R690 VTAIL.n191 VTAIL.n135 0.155672
R691 VTAIL.n184 VTAIL.n135 0.155672
R692 VTAIL.n184 VTAIL.n183 0.155672
R693 VTAIL.n183 VTAIL.n139 0.155672
R694 VTAIL.n176 VTAIL.n139 0.155672
R695 VTAIL.n176 VTAIL.n175 0.155672
R696 VTAIL.n175 VTAIL.n143 0.155672
R697 VTAIL.n168 VTAIL.n143 0.155672
R698 VTAIL.n168 VTAIL.n167 0.155672
R699 VTAIL.n167 VTAIL.n147 0.155672
R700 VTAIL.n160 VTAIL.n147 0.155672
R701 VTAIL.n160 VTAIL.n159 0.155672
R702 VTAIL.n159 VTAIL.n151 0.155672
R703 VDD2.n215 VDD2.n111 289.615
R704 VDD2.n104 VDD2.n0 289.615
R705 VDD2.n216 VDD2.n215 185
R706 VDD2.n214 VDD2.n213 185
R707 VDD2.n115 VDD2.n114 185
R708 VDD2.n208 VDD2.n207 185
R709 VDD2.n206 VDD2.n205 185
R710 VDD2.n119 VDD2.n118 185
R711 VDD2.n200 VDD2.n199 185
R712 VDD2.n198 VDD2.n197 185
R713 VDD2.n123 VDD2.n122 185
R714 VDD2.n127 VDD2.n125 185
R715 VDD2.n192 VDD2.n191 185
R716 VDD2.n190 VDD2.n189 185
R717 VDD2.n129 VDD2.n128 185
R718 VDD2.n184 VDD2.n183 185
R719 VDD2.n182 VDD2.n181 185
R720 VDD2.n133 VDD2.n132 185
R721 VDD2.n176 VDD2.n175 185
R722 VDD2.n174 VDD2.n173 185
R723 VDD2.n137 VDD2.n136 185
R724 VDD2.n168 VDD2.n167 185
R725 VDD2.n166 VDD2.n165 185
R726 VDD2.n141 VDD2.n140 185
R727 VDD2.n160 VDD2.n159 185
R728 VDD2.n158 VDD2.n157 185
R729 VDD2.n145 VDD2.n144 185
R730 VDD2.n152 VDD2.n151 185
R731 VDD2.n150 VDD2.n149 185
R732 VDD2.n37 VDD2.n36 185
R733 VDD2.n39 VDD2.n38 185
R734 VDD2.n32 VDD2.n31 185
R735 VDD2.n45 VDD2.n44 185
R736 VDD2.n47 VDD2.n46 185
R737 VDD2.n28 VDD2.n27 185
R738 VDD2.n53 VDD2.n52 185
R739 VDD2.n55 VDD2.n54 185
R740 VDD2.n24 VDD2.n23 185
R741 VDD2.n61 VDD2.n60 185
R742 VDD2.n63 VDD2.n62 185
R743 VDD2.n20 VDD2.n19 185
R744 VDD2.n69 VDD2.n68 185
R745 VDD2.n71 VDD2.n70 185
R746 VDD2.n16 VDD2.n15 185
R747 VDD2.n78 VDD2.n77 185
R748 VDD2.n79 VDD2.n14 185
R749 VDD2.n81 VDD2.n80 185
R750 VDD2.n12 VDD2.n11 185
R751 VDD2.n87 VDD2.n86 185
R752 VDD2.n89 VDD2.n88 185
R753 VDD2.n8 VDD2.n7 185
R754 VDD2.n95 VDD2.n94 185
R755 VDD2.n97 VDD2.n96 185
R756 VDD2.n4 VDD2.n3 185
R757 VDD2.n103 VDD2.n102 185
R758 VDD2.n105 VDD2.n104 185
R759 VDD2.n148 VDD2.t0 147.659
R760 VDD2.n35 VDD2.t5 147.659
R761 VDD2.n215 VDD2.n214 104.615
R762 VDD2.n214 VDD2.n114 104.615
R763 VDD2.n207 VDD2.n114 104.615
R764 VDD2.n207 VDD2.n206 104.615
R765 VDD2.n206 VDD2.n118 104.615
R766 VDD2.n199 VDD2.n118 104.615
R767 VDD2.n199 VDD2.n198 104.615
R768 VDD2.n198 VDD2.n122 104.615
R769 VDD2.n127 VDD2.n122 104.615
R770 VDD2.n191 VDD2.n127 104.615
R771 VDD2.n191 VDD2.n190 104.615
R772 VDD2.n190 VDD2.n128 104.615
R773 VDD2.n183 VDD2.n128 104.615
R774 VDD2.n183 VDD2.n182 104.615
R775 VDD2.n182 VDD2.n132 104.615
R776 VDD2.n175 VDD2.n132 104.615
R777 VDD2.n175 VDD2.n174 104.615
R778 VDD2.n174 VDD2.n136 104.615
R779 VDD2.n167 VDD2.n136 104.615
R780 VDD2.n167 VDD2.n166 104.615
R781 VDD2.n166 VDD2.n140 104.615
R782 VDD2.n159 VDD2.n140 104.615
R783 VDD2.n159 VDD2.n158 104.615
R784 VDD2.n158 VDD2.n144 104.615
R785 VDD2.n151 VDD2.n144 104.615
R786 VDD2.n151 VDD2.n150 104.615
R787 VDD2.n38 VDD2.n37 104.615
R788 VDD2.n38 VDD2.n31 104.615
R789 VDD2.n45 VDD2.n31 104.615
R790 VDD2.n46 VDD2.n45 104.615
R791 VDD2.n46 VDD2.n27 104.615
R792 VDD2.n53 VDD2.n27 104.615
R793 VDD2.n54 VDD2.n53 104.615
R794 VDD2.n54 VDD2.n23 104.615
R795 VDD2.n61 VDD2.n23 104.615
R796 VDD2.n62 VDD2.n61 104.615
R797 VDD2.n62 VDD2.n19 104.615
R798 VDD2.n69 VDD2.n19 104.615
R799 VDD2.n70 VDD2.n69 104.615
R800 VDD2.n70 VDD2.n15 104.615
R801 VDD2.n78 VDD2.n15 104.615
R802 VDD2.n79 VDD2.n78 104.615
R803 VDD2.n80 VDD2.n79 104.615
R804 VDD2.n80 VDD2.n11 104.615
R805 VDD2.n87 VDD2.n11 104.615
R806 VDD2.n88 VDD2.n87 104.615
R807 VDD2.n88 VDD2.n7 104.615
R808 VDD2.n95 VDD2.n7 104.615
R809 VDD2.n96 VDD2.n95 104.615
R810 VDD2.n96 VDD2.n3 104.615
R811 VDD2.n103 VDD2.n3 104.615
R812 VDD2.n104 VDD2.n103 104.615
R813 VDD2.n110 VDD2.n109 60.1782
R814 VDD2 VDD2.n221 60.1753
R815 VDD2.n150 VDD2.t0 52.3082
R816 VDD2.n37 VDD2.t5 52.3082
R817 VDD2.n110 VDD2.n108 48.8671
R818 VDD2.n220 VDD2.n219 48.2823
R819 VDD2.n220 VDD2.n110 43.4287
R820 VDD2.n149 VDD2.n148 15.6677
R821 VDD2.n36 VDD2.n35 15.6677
R822 VDD2.n125 VDD2.n123 13.1884
R823 VDD2.n81 VDD2.n12 13.1884
R824 VDD2.n197 VDD2.n196 12.8005
R825 VDD2.n193 VDD2.n192 12.8005
R826 VDD2.n152 VDD2.n147 12.8005
R827 VDD2.n39 VDD2.n34 12.8005
R828 VDD2.n82 VDD2.n14 12.8005
R829 VDD2.n86 VDD2.n85 12.8005
R830 VDD2.n200 VDD2.n121 12.0247
R831 VDD2.n189 VDD2.n126 12.0247
R832 VDD2.n153 VDD2.n145 12.0247
R833 VDD2.n40 VDD2.n32 12.0247
R834 VDD2.n77 VDD2.n76 12.0247
R835 VDD2.n89 VDD2.n10 12.0247
R836 VDD2.n201 VDD2.n119 11.249
R837 VDD2.n188 VDD2.n129 11.249
R838 VDD2.n157 VDD2.n156 11.249
R839 VDD2.n44 VDD2.n43 11.249
R840 VDD2.n75 VDD2.n16 11.249
R841 VDD2.n90 VDD2.n8 11.249
R842 VDD2.n205 VDD2.n204 10.4732
R843 VDD2.n185 VDD2.n184 10.4732
R844 VDD2.n160 VDD2.n143 10.4732
R845 VDD2.n47 VDD2.n30 10.4732
R846 VDD2.n72 VDD2.n71 10.4732
R847 VDD2.n94 VDD2.n93 10.4732
R848 VDD2.n208 VDD2.n117 9.69747
R849 VDD2.n181 VDD2.n131 9.69747
R850 VDD2.n161 VDD2.n141 9.69747
R851 VDD2.n48 VDD2.n28 9.69747
R852 VDD2.n68 VDD2.n18 9.69747
R853 VDD2.n97 VDD2.n6 9.69747
R854 VDD2.n219 VDD2.n218 9.45567
R855 VDD2.n108 VDD2.n107 9.45567
R856 VDD2.n135 VDD2.n134 9.3005
R857 VDD2.n178 VDD2.n177 9.3005
R858 VDD2.n180 VDD2.n179 9.3005
R859 VDD2.n131 VDD2.n130 9.3005
R860 VDD2.n186 VDD2.n185 9.3005
R861 VDD2.n188 VDD2.n187 9.3005
R862 VDD2.n126 VDD2.n124 9.3005
R863 VDD2.n194 VDD2.n193 9.3005
R864 VDD2.n218 VDD2.n217 9.3005
R865 VDD2.n113 VDD2.n112 9.3005
R866 VDD2.n212 VDD2.n211 9.3005
R867 VDD2.n210 VDD2.n209 9.3005
R868 VDD2.n117 VDD2.n116 9.3005
R869 VDD2.n204 VDD2.n203 9.3005
R870 VDD2.n202 VDD2.n201 9.3005
R871 VDD2.n121 VDD2.n120 9.3005
R872 VDD2.n196 VDD2.n195 9.3005
R873 VDD2.n172 VDD2.n171 9.3005
R874 VDD2.n170 VDD2.n169 9.3005
R875 VDD2.n139 VDD2.n138 9.3005
R876 VDD2.n164 VDD2.n163 9.3005
R877 VDD2.n162 VDD2.n161 9.3005
R878 VDD2.n143 VDD2.n142 9.3005
R879 VDD2.n156 VDD2.n155 9.3005
R880 VDD2.n154 VDD2.n153 9.3005
R881 VDD2.n147 VDD2.n146 9.3005
R882 VDD2.n107 VDD2.n106 9.3005
R883 VDD2.n101 VDD2.n100 9.3005
R884 VDD2.n99 VDD2.n98 9.3005
R885 VDD2.n6 VDD2.n5 9.3005
R886 VDD2.n93 VDD2.n92 9.3005
R887 VDD2.n91 VDD2.n90 9.3005
R888 VDD2.n10 VDD2.n9 9.3005
R889 VDD2.n85 VDD2.n84 9.3005
R890 VDD2.n57 VDD2.n56 9.3005
R891 VDD2.n26 VDD2.n25 9.3005
R892 VDD2.n51 VDD2.n50 9.3005
R893 VDD2.n49 VDD2.n48 9.3005
R894 VDD2.n30 VDD2.n29 9.3005
R895 VDD2.n43 VDD2.n42 9.3005
R896 VDD2.n41 VDD2.n40 9.3005
R897 VDD2.n34 VDD2.n33 9.3005
R898 VDD2.n59 VDD2.n58 9.3005
R899 VDD2.n22 VDD2.n21 9.3005
R900 VDD2.n65 VDD2.n64 9.3005
R901 VDD2.n67 VDD2.n66 9.3005
R902 VDD2.n18 VDD2.n17 9.3005
R903 VDD2.n73 VDD2.n72 9.3005
R904 VDD2.n75 VDD2.n74 9.3005
R905 VDD2.n76 VDD2.n13 9.3005
R906 VDD2.n83 VDD2.n82 9.3005
R907 VDD2.n2 VDD2.n1 9.3005
R908 VDD2.n209 VDD2.n115 8.92171
R909 VDD2.n180 VDD2.n133 8.92171
R910 VDD2.n165 VDD2.n164 8.92171
R911 VDD2.n52 VDD2.n51 8.92171
R912 VDD2.n67 VDD2.n20 8.92171
R913 VDD2.n98 VDD2.n4 8.92171
R914 VDD2.n213 VDD2.n212 8.14595
R915 VDD2.n177 VDD2.n176 8.14595
R916 VDD2.n168 VDD2.n139 8.14595
R917 VDD2.n55 VDD2.n26 8.14595
R918 VDD2.n64 VDD2.n63 8.14595
R919 VDD2.n102 VDD2.n101 8.14595
R920 VDD2.n219 VDD2.n111 7.3702
R921 VDD2.n216 VDD2.n113 7.3702
R922 VDD2.n173 VDD2.n135 7.3702
R923 VDD2.n169 VDD2.n137 7.3702
R924 VDD2.n56 VDD2.n24 7.3702
R925 VDD2.n60 VDD2.n22 7.3702
R926 VDD2.n105 VDD2.n2 7.3702
R927 VDD2.n108 VDD2.n0 7.3702
R928 VDD2.n217 VDD2.n111 6.59444
R929 VDD2.n217 VDD2.n216 6.59444
R930 VDD2.n173 VDD2.n172 6.59444
R931 VDD2.n172 VDD2.n137 6.59444
R932 VDD2.n59 VDD2.n24 6.59444
R933 VDD2.n60 VDD2.n59 6.59444
R934 VDD2.n106 VDD2.n105 6.59444
R935 VDD2.n106 VDD2.n0 6.59444
R936 VDD2.n213 VDD2.n113 5.81868
R937 VDD2.n176 VDD2.n135 5.81868
R938 VDD2.n169 VDD2.n168 5.81868
R939 VDD2.n56 VDD2.n55 5.81868
R940 VDD2.n63 VDD2.n22 5.81868
R941 VDD2.n102 VDD2.n2 5.81868
R942 VDD2.n212 VDD2.n115 5.04292
R943 VDD2.n177 VDD2.n133 5.04292
R944 VDD2.n165 VDD2.n139 5.04292
R945 VDD2.n52 VDD2.n26 5.04292
R946 VDD2.n64 VDD2.n20 5.04292
R947 VDD2.n101 VDD2.n4 5.04292
R948 VDD2.n148 VDD2.n146 4.38563
R949 VDD2.n35 VDD2.n33 4.38563
R950 VDD2.n209 VDD2.n208 4.26717
R951 VDD2.n181 VDD2.n180 4.26717
R952 VDD2.n164 VDD2.n141 4.26717
R953 VDD2.n51 VDD2.n28 4.26717
R954 VDD2.n68 VDD2.n67 4.26717
R955 VDD2.n98 VDD2.n97 4.26717
R956 VDD2.n205 VDD2.n117 3.49141
R957 VDD2.n184 VDD2.n131 3.49141
R958 VDD2.n161 VDD2.n160 3.49141
R959 VDD2.n48 VDD2.n47 3.49141
R960 VDD2.n71 VDD2.n18 3.49141
R961 VDD2.n94 VDD2.n6 3.49141
R962 VDD2.n204 VDD2.n119 2.71565
R963 VDD2.n185 VDD2.n129 2.71565
R964 VDD2.n157 VDD2.n143 2.71565
R965 VDD2.n44 VDD2.n30 2.71565
R966 VDD2.n72 VDD2.n16 2.71565
R967 VDD2.n93 VDD2.n8 2.71565
R968 VDD2.n201 VDD2.n200 1.93989
R969 VDD2.n189 VDD2.n188 1.93989
R970 VDD2.n156 VDD2.n145 1.93989
R971 VDD2.n43 VDD2.n32 1.93989
R972 VDD2.n77 VDD2.n75 1.93989
R973 VDD2.n90 VDD2.n89 1.93989
R974 VDD2.n197 VDD2.n121 1.16414
R975 VDD2.n192 VDD2.n126 1.16414
R976 VDD2.n153 VDD2.n152 1.16414
R977 VDD2.n40 VDD2.n39 1.16414
R978 VDD2.n76 VDD2.n14 1.16414
R979 VDD2.n86 VDD2.n10 1.16414
R980 VDD2.n221 VDD2.t1 1.00813
R981 VDD2.n221 VDD2.t2 1.00813
R982 VDD2.n109 VDD2.t3 1.00813
R983 VDD2.n109 VDD2.t4 1.00813
R984 VDD2 VDD2.n220 0.698776
R985 VDD2.n196 VDD2.n123 0.388379
R986 VDD2.n193 VDD2.n125 0.388379
R987 VDD2.n149 VDD2.n147 0.388379
R988 VDD2.n36 VDD2.n34 0.388379
R989 VDD2.n82 VDD2.n81 0.388379
R990 VDD2.n85 VDD2.n12 0.388379
R991 VDD2.n218 VDD2.n112 0.155672
R992 VDD2.n211 VDD2.n112 0.155672
R993 VDD2.n211 VDD2.n210 0.155672
R994 VDD2.n210 VDD2.n116 0.155672
R995 VDD2.n203 VDD2.n116 0.155672
R996 VDD2.n203 VDD2.n202 0.155672
R997 VDD2.n202 VDD2.n120 0.155672
R998 VDD2.n195 VDD2.n120 0.155672
R999 VDD2.n195 VDD2.n194 0.155672
R1000 VDD2.n194 VDD2.n124 0.155672
R1001 VDD2.n187 VDD2.n124 0.155672
R1002 VDD2.n187 VDD2.n186 0.155672
R1003 VDD2.n186 VDD2.n130 0.155672
R1004 VDD2.n179 VDD2.n130 0.155672
R1005 VDD2.n179 VDD2.n178 0.155672
R1006 VDD2.n178 VDD2.n134 0.155672
R1007 VDD2.n171 VDD2.n134 0.155672
R1008 VDD2.n171 VDD2.n170 0.155672
R1009 VDD2.n170 VDD2.n138 0.155672
R1010 VDD2.n163 VDD2.n138 0.155672
R1011 VDD2.n163 VDD2.n162 0.155672
R1012 VDD2.n162 VDD2.n142 0.155672
R1013 VDD2.n155 VDD2.n142 0.155672
R1014 VDD2.n155 VDD2.n154 0.155672
R1015 VDD2.n154 VDD2.n146 0.155672
R1016 VDD2.n41 VDD2.n33 0.155672
R1017 VDD2.n42 VDD2.n41 0.155672
R1018 VDD2.n42 VDD2.n29 0.155672
R1019 VDD2.n49 VDD2.n29 0.155672
R1020 VDD2.n50 VDD2.n49 0.155672
R1021 VDD2.n50 VDD2.n25 0.155672
R1022 VDD2.n57 VDD2.n25 0.155672
R1023 VDD2.n58 VDD2.n57 0.155672
R1024 VDD2.n58 VDD2.n21 0.155672
R1025 VDD2.n65 VDD2.n21 0.155672
R1026 VDD2.n66 VDD2.n65 0.155672
R1027 VDD2.n66 VDD2.n17 0.155672
R1028 VDD2.n73 VDD2.n17 0.155672
R1029 VDD2.n74 VDD2.n73 0.155672
R1030 VDD2.n74 VDD2.n13 0.155672
R1031 VDD2.n83 VDD2.n13 0.155672
R1032 VDD2.n84 VDD2.n83 0.155672
R1033 VDD2.n84 VDD2.n9 0.155672
R1034 VDD2.n91 VDD2.n9 0.155672
R1035 VDD2.n92 VDD2.n91 0.155672
R1036 VDD2.n92 VDD2.n5 0.155672
R1037 VDD2.n99 VDD2.n5 0.155672
R1038 VDD2.n100 VDD2.n99 0.155672
R1039 VDD2.n100 VDD2.n1 0.155672
R1040 VDD2.n107 VDD2.n1 0.155672
R1041 B.n113 B.t14 921.01
R1042 B.n110 B.t10 921.01
R1043 B.n492 B.t6 921.01
R1044 B.n490 B.t17 921.01
R1045 B.n855 B.n854 585
R1046 B.n384 B.n108 585
R1047 B.n383 B.n382 585
R1048 B.n381 B.n380 585
R1049 B.n379 B.n378 585
R1050 B.n377 B.n376 585
R1051 B.n375 B.n374 585
R1052 B.n373 B.n372 585
R1053 B.n371 B.n370 585
R1054 B.n369 B.n368 585
R1055 B.n367 B.n366 585
R1056 B.n365 B.n364 585
R1057 B.n363 B.n362 585
R1058 B.n361 B.n360 585
R1059 B.n359 B.n358 585
R1060 B.n357 B.n356 585
R1061 B.n355 B.n354 585
R1062 B.n353 B.n352 585
R1063 B.n351 B.n350 585
R1064 B.n349 B.n348 585
R1065 B.n347 B.n346 585
R1066 B.n345 B.n344 585
R1067 B.n343 B.n342 585
R1068 B.n341 B.n340 585
R1069 B.n339 B.n338 585
R1070 B.n337 B.n336 585
R1071 B.n335 B.n334 585
R1072 B.n333 B.n332 585
R1073 B.n331 B.n330 585
R1074 B.n329 B.n328 585
R1075 B.n327 B.n326 585
R1076 B.n325 B.n324 585
R1077 B.n323 B.n322 585
R1078 B.n321 B.n320 585
R1079 B.n319 B.n318 585
R1080 B.n317 B.n316 585
R1081 B.n315 B.n314 585
R1082 B.n313 B.n312 585
R1083 B.n311 B.n310 585
R1084 B.n309 B.n308 585
R1085 B.n307 B.n306 585
R1086 B.n305 B.n304 585
R1087 B.n303 B.n302 585
R1088 B.n301 B.n300 585
R1089 B.n299 B.n298 585
R1090 B.n297 B.n296 585
R1091 B.n295 B.n294 585
R1092 B.n293 B.n292 585
R1093 B.n291 B.n290 585
R1094 B.n289 B.n288 585
R1095 B.n287 B.n286 585
R1096 B.n285 B.n284 585
R1097 B.n283 B.n282 585
R1098 B.n281 B.n280 585
R1099 B.n279 B.n278 585
R1100 B.n277 B.n276 585
R1101 B.n275 B.n274 585
R1102 B.n273 B.n272 585
R1103 B.n271 B.n270 585
R1104 B.n269 B.n268 585
R1105 B.n267 B.n266 585
R1106 B.n265 B.n264 585
R1107 B.n263 B.n262 585
R1108 B.n261 B.n260 585
R1109 B.n259 B.n258 585
R1110 B.n257 B.n256 585
R1111 B.n255 B.n254 585
R1112 B.n253 B.n252 585
R1113 B.n251 B.n250 585
R1114 B.n249 B.n248 585
R1115 B.n247 B.n246 585
R1116 B.n245 B.n244 585
R1117 B.n243 B.n242 585
R1118 B.n241 B.n240 585
R1119 B.n239 B.n238 585
R1120 B.n237 B.n236 585
R1121 B.n235 B.n234 585
R1122 B.n233 B.n232 585
R1123 B.n231 B.n230 585
R1124 B.n229 B.n228 585
R1125 B.n227 B.n226 585
R1126 B.n225 B.n224 585
R1127 B.n223 B.n222 585
R1128 B.n221 B.n220 585
R1129 B.n219 B.n218 585
R1130 B.n217 B.n216 585
R1131 B.n215 B.n214 585
R1132 B.n213 B.n212 585
R1133 B.n211 B.n210 585
R1134 B.n209 B.n208 585
R1135 B.n207 B.n206 585
R1136 B.n205 B.n204 585
R1137 B.n203 B.n202 585
R1138 B.n201 B.n200 585
R1139 B.n199 B.n198 585
R1140 B.n197 B.n196 585
R1141 B.n195 B.n194 585
R1142 B.n193 B.n192 585
R1143 B.n191 B.n190 585
R1144 B.n189 B.n188 585
R1145 B.n187 B.n186 585
R1146 B.n185 B.n184 585
R1147 B.n183 B.n182 585
R1148 B.n181 B.n180 585
R1149 B.n179 B.n178 585
R1150 B.n177 B.n176 585
R1151 B.n175 B.n174 585
R1152 B.n173 B.n172 585
R1153 B.n171 B.n170 585
R1154 B.n169 B.n168 585
R1155 B.n167 B.n166 585
R1156 B.n165 B.n164 585
R1157 B.n163 B.n162 585
R1158 B.n161 B.n160 585
R1159 B.n159 B.n158 585
R1160 B.n157 B.n156 585
R1161 B.n155 B.n154 585
R1162 B.n153 B.n152 585
R1163 B.n151 B.n150 585
R1164 B.n149 B.n148 585
R1165 B.n147 B.n146 585
R1166 B.n145 B.n144 585
R1167 B.n143 B.n142 585
R1168 B.n141 B.n140 585
R1169 B.n139 B.n138 585
R1170 B.n137 B.n136 585
R1171 B.n135 B.n134 585
R1172 B.n133 B.n132 585
R1173 B.n131 B.n130 585
R1174 B.n129 B.n128 585
R1175 B.n127 B.n126 585
R1176 B.n125 B.n124 585
R1177 B.n123 B.n122 585
R1178 B.n121 B.n120 585
R1179 B.n119 B.n118 585
R1180 B.n117 B.n116 585
R1181 B.n40 B.n39 585
R1182 B.n860 B.n859 585
R1183 B.n853 B.n109 585
R1184 B.n109 B.n37 585
R1185 B.n852 B.n36 585
R1186 B.n864 B.n36 585
R1187 B.n851 B.n35 585
R1188 B.n865 B.n35 585
R1189 B.n850 B.n34 585
R1190 B.n866 B.n34 585
R1191 B.n849 B.n848 585
R1192 B.n848 B.n33 585
R1193 B.n847 B.n29 585
R1194 B.n872 B.n29 585
R1195 B.n846 B.n28 585
R1196 B.n873 B.n28 585
R1197 B.n845 B.n27 585
R1198 B.n874 B.n27 585
R1199 B.n844 B.n843 585
R1200 B.n843 B.n23 585
R1201 B.n842 B.n22 585
R1202 B.n880 B.n22 585
R1203 B.n841 B.n21 585
R1204 B.n881 B.n21 585
R1205 B.n840 B.n20 585
R1206 B.n882 B.n20 585
R1207 B.n839 B.n838 585
R1208 B.n838 B.n16 585
R1209 B.n837 B.n15 585
R1210 B.n888 B.n15 585
R1211 B.n836 B.n14 585
R1212 B.n889 B.n14 585
R1213 B.n835 B.n13 585
R1214 B.n890 B.n13 585
R1215 B.n834 B.n833 585
R1216 B.n833 B.n12 585
R1217 B.n832 B.n831 585
R1218 B.n832 B.n8 585
R1219 B.n830 B.n7 585
R1220 B.n897 B.n7 585
R1221 B.n829 B.n6 585
R1222 B.n898 B.n6 585
R1223 B.n828 B.n5 585
R1224 B.n899 B.n5 585
R1225 B.n827 B.n826 585
R1226 B.n826 B.n4 585
R1227 B.n825 B.n385 585
R1228 B.n825 B.n824 585
R1229 B.n814 B.n386 585
R1230 B.n817 B.n386 585
R1231 B.n816 B.n815 585
R1232 B.n818 B.n816 585
R1233 B.n813 B.n391 585
R1234 B.n391 B.n390 585
R1235 B.n812 B.n811 585
R1236 B.n811 B.n810 585
R1237 B.n393 B.n392 585
R1238 B.n394 B.n393 585
R1239 B.n803 B.n802 585
R1240 B.n804 B.n803 585
R1241 B.n801 B.n398 585
R1242 B.n402 B.n398 585
R1243 B.n800 B.n799 585
R1244 B.n799 B.n798 585
R1245 B.n400 B.n399 585
R1246 B.n401 B.n400 585
R1247 B.n791 B.n790 585
R1248 B.n792 B.n791 585
R1249 B.n789 B.n407 585
R1250 B.n407 B.n406 585
R1251 B.n788 B.n787 585
R1252 B.n787 B.n786 585
R1253 B.n409 B.n408 585
R1254 B.n779 B.n409 585
R1255 B.n778 B.n777 585
R1256 B.n780 B.n778 585
R1257 B.n776 B.n414 585
R1258 B.n414 B.n413 585
R1259 B.n775 B.n774 585
R1260 B.n774 B.n773 585
R1261 B.n416 B.n415 585
R1262 B.n417 B.n416 585
R1263 B.n769 B.n768 585
R1264 B.n420 B.n419 585
R1265 B.n765 B.n764 585
R1266 B.n766 B.n765 585
R1267 B.n763 B.n489 585
R1268 B.n762 B.n761 585
R1269 B.n760 B.n759 585
R1270 B.n758 B.n757 585
R1271 B.n756 B.n755 585
R1272 B.n754 B.n753 585
R1273 B.n752 B.n751 585
R1274 B.n750 B.n749 585
R1275 B.n748 B.n747 585
R1276 B.n746 B.n745 585
R1277 B.n744 B.n743 585
R1278 B.n742 B.n741 585
R1279 B.n740 B.n739 585
R1280 B.n738 B.n737 585
R1281 B.n736 B.n735 585
R1282 B.n734 B.n733 585
R1283 B.n732 B.n731 585
R1284 B.n730 B.n729 585
R1285 B.n728 B.n727 585
R1286 B.n726 B.n725 585
R1287 B.n724 B.n723 585
R1288 B.n722 B.n721 585
R1289 B.n720 B.n719 585
R1290 B.n718 B.n717 585
R1291 B.n716 B.n715 585
R1292 B.n714 B.n713 585
R1293 B.n712 B.n711 585
R1294 B.n710 B.n709 585
R1295 B.n708 B.n707 585
R1296 B.n706 B.n705 585
R1297 B.n704 B.n703 585
R1298 B.n702 B.n701 585
R1299 B.n700 B.n699 585
R1300 B.n698 B.n697 585
R1301 B.n696 B.n695 585
R1302 B.n694 B.n693 585
R1303 B.n692 B.n691 585
R1304 B.n690 B.n689 585
R1305 B.n688 B.n687 585
R1306 B.n686 B.n685 585
R1307 B.n684 B.n683 585
R1308 B.n682 B.n681 585
R1309 B.n680 B.n679 585
R1310 B.n678 B.n677 585
R1311 B.n676 B.n675 585
R1312 B.n674 B.n673 585
R1313 B.n672 B.n671 585
R1314 B.n670 B.n669 585
R1315 B.n668 B.n667 585
R1316 B.n666 B.n665 585
R1317 B.n664 B.n663 585
R1318 B.n662 B.n661 585
R1319 B.n660 B.n659 585
R1320 B.n658 B.n657 585
R1321 B.n656 B.n655 585
R1322 B.n654 B.n653 585
R1323 B.n652 B.n651 585
R1324 B.n650 B.n649 585
R1325 B.n648 B.n647 585
R1326 B.n646 B.n645 585
R1327 B.n644 B.n643 585
R1328 B.n641 B.n640 585
R1329 B.n639 B.n638 585
R1330 B.n637 B.n636 585
R1331 B.n635 B.n634 585
R1332 B.n633 B.n632 585
R1333 B.n631 B.n630 585
R1334 B.n629 B.n628 585
R1335 B.n627 B.n626 585
R1336 B.n625 B.n624 585
R1337 B.n623 B.n622 585
R1338 B.n620 B.n619 585
R1339 B.n618 B.n617 585
R1340 B.n616 B.n615 585
R1341 B.n614 B.n613 585
R1342 B.n612 B.n611 585
R1343 B.n610 B.n609 585
R1344 B.n608 B.n607 585
R1345 B.n606 B.n605 585
R1346 B.n604 B.n603 585
R1347 B.n602 B.n601 585
R1348 B.n600 B.n599 585
R1349 B.n598 B.n597 585
R1350 B.n596 B.n595 585
R1351 B.n594 B.n593 585
R1352 B.n592 B.n591 585
R1353 B.n590 B.n589 585
R1354 B.n588 B.n587 585
R1355 B.n586 B.n585 585
R1356 B.n584 B.n583 585
R1357 B.n582 B.n581 585
R1358 B.n580 B.n579 585
R1359 B.n578 B.n577 585
R1360 B.n576 B.n575 585
R1361 B.n574 B.n573 585
R1362 B.n572 B.n571 585
R1363 B.n570 B.n569 585
R1364 B.n568 B.n567 585
R1365 B.n566 B.n565 585
R1366 B.n564 B.n563 585
R1367 B.n562 B.n561 585
R1368 B.n560 B.n559 585
R1369 B.n558 B.n557 585
R1370 B.n556 B.n555 585
R1371 B.n554 B.n553 585
R1372 B.n552 B.n551 585
R1373 B.n550 B.n549 585
R1374 B.n548 B.n547 585
R1375 B.n546 B.n545 585
R1376 B.n544 B.n543 585
R1377 B.n542 B.n541 585
R1378 B.n540 B.n539 585
R1379 B.n538 B.n537 585
R1380 B.n536 B.n535 585
R1381 B.n534 B.n533 585
R1382 B.n532 B.n531 585
R1383 B.n530 B.n529 585
R1384 B.n528 B.n527 585
R1385 B.n526 B.n525 585
R1386 B.n524 B.n523 585
R1387 B.n522 B.n521 585
R1388 B.n520 B.n519 585
R1389 B.n518 B.n517 585
R1390 B.n516 B.n515 585
R1391 B.n514 B.n513 585
R1392 B.n512 B.n511 585
R1393 B.n510 B.n509 585
R1394 B.n508 B.n507 585
R1395 B.n506 B.n505 585
R1396 B.n504 B.n503 585
R1397 B.n502 B.n501 585
R1398 B.n500 B.n499 585
R1399 B.n498 B.n497 585
R1400 B.n496 B.n495 585
R1401 B.n494 B.n488 585
R1402 B.n766 B.n488 585
R1403 B.n770 B.n418 585
R1404 B.n418 B.n417 585
R1405 B.n772 B.n771 585
R1406 B.n773 B.n772 585
R1407 B.n412 B.n411 585
R1408 B.n413 B.n412 585
R1409 B.n782 B.n781 585
R1410 B.n781 B.n780 585
R1411 B.n783 B.n410 585
R1412 B.n779 B.n410 585
R1413 B.n785 B.n784 585
R1414 B.n786 B.n785 585
R1415 B.n405 B.n404 585
R1416 B.n406 B.n405 585
R1417 B.n794 B.n793 585
R1418 B.n793 B.n792 585
R1419 B.n795 B.n403 585
R1420 B.n403 B.n401 585
R1421 B.n797 B.n796 585
R1422 B.n798 B.n797 585
R1423 B.n397 B.n396 585
R1424 B.n402 B.n397 585
R1425 B.n806 B.n805 585
R1426 B.n805 B.n804 585
R1427 B.n807 B.n395 585
R1428 B.n395 B.n394 585
R1429 B.n809 B.n808 585
R1430 B.n810 B.n809 585
R1431 B.n389 B.n388 585
R1432 B.n390 B.n389 585
R1433 B.n820 B.n819 585
R1434 B.n819 B.n818 585
R1435 B.n821 B.n387 585
R1436 B.n817 B.n387 585
R1437 B.n823 B.n822 585
R1438 B.n824 B.n823 585
R1439 B.n3 B.n0 585
R1440 B.n4 B.n3 585
R1441 B.n896 B.n1 585
R1442 B.n897 B.n896 585
R1443 B.n895 B.n894 585
R1444 B.n895 B.n8 585
R1445 B.n893 B.n9 585
R1446 B.n12 B.n9 585
R1447 B.n892 B.n891 585
R1448 B.n891 B.n890 585
R1449 B.n11 B.n10 585
R1450 B.n889 B.n11 585
R1451 B.n887 B.n886 585
R1452 B.n888 B.n887 585
R1453 B.n885 B.n17 585
R1454 B.n17 B.n16 585
R1455 B.n884 B.n883 585
R1456 B.n883 B.n882 585
R1457 B.n19 B.n18 585
R1458 B.n881 B.n19 585
R1459 B.n879 B.n878 585
R1460 B.n880 B.n879 585
R1461 B.n877 B.n24 585
R1462 B.n24 B.n23 585
R1463 B.n876 B.n875 585
R1464 B.n875 B.n874 585
R1465 B.n26 B.n25 585
R1466 B.n873 B.n26 585
R1467 B.n871 B.n870 585
R1468 B.n872 B.n871 585
R1469 B.n869 B.n30 585
R1470 B.n33 B.n30 585
R1471 B.n868 B.n867 585
R1472 B.n867 B.n866 585
R1473 B.n32 B.n31 585
R1474 B.n865 B.n32 585
R1475 B.n863 B.n862 585
R1476 B.n864 B.n863 585
R1477 B.n861 B.n38 585
R1478 B.n38 B.n37 585
R1479 B.n900 B.n899 585
R1480 B.n898 B.n2 585
R1481 B.n859 B.n38 526.135
R1482 B.n855 B.n109 526.135
R1483 B.n488 B.n416 526.135
R1484 B.n768 B.n418 526.135
R1485 B.n110 B.t12 433.341
R1486 B.n492 B.t9 433.341
R1487 B.n113 B.t15 433.341
R1488 B.n490 B.t19 433.341
R1489 B.n111 B.t13 414.142
R1490 B.n493 B.t8 414.142
R1491 B.n114 B.t16 414.142
R1492 B.n491 B.t18 414.142
R1493 B.n857 B.n856 256.663
R1494 B.n857 B.n107 256.663
R1495 B.n857 B.n106 256.663
R1496 B.n857 B.n105 256.663
R1497 B.n857 B.n104 256.663
R1498 B.n857 B.n103 256.663
R1499 B.n857 B.n102 256.663
R1500 B.n857 B.n101 256.663
R1501 B.n857 B.n100 256.663
R1502 B.n857 B.n99 256.663
R1503 B.n857 B.n98 256.663
R1504 B.n857 B.n97 256.663
R1505 B.n857 B.n96 256.663
R1506 B.n857 B.n95 256.663
R1507 B.n857 B.n94 256.663
R1508 B.n857 B.n93 256.663
R1509 B.n857 B.n92 256.663
R1510 B.n857 B.n91 256.663
R1511 B.n857 B.n90 256.663
R1512 B.n857 B.n89 256.663
R1513 B.n857 B.n88 256.663
R1514 B.n857 B.n87 256.663
R1515 B.n857 B.n86 256.663
R1516 B.n857 B.n85 256.663
R1517 B.n857 B.n84 256.663
R1518 B.n857 B.n83 256.663
R1519 B.n857 B.n82 256.663
R1520 B.n857 B.n81 256.663
R1521 B.n857 B.n80 256.663
R1522 B.n857 B.n79 256.663
R1523 B.n857 B.n78 256.663
R1524 B.n857 B.n77 256.663
R1525 B.n857 B.n76 256.663
R1526 B.n857 B.n75 256.663
R1527 B.n857 B.n74 256.663
R1528 B.n857 B.n73 256.663
R1529 B.n857 B.n72 256.663
R1530 B.n857 B.n71 256.663
R1531 B.n857 B.n70 256.663
R1532 B.n857 B.n69 256.663
R1533 B.n857 B.n68 256.663
R1534 B.n857 B.n67 256.663
R1535 B.n857 B.n66 256.663
R1536 B.n857 B.n65 256.663
R1537 B.n857 B.n64 256.663
R1538 B.n857 B.n63 256.663
R1539 B.n857 B.n62 256.663
R1540 B.n857 B.n61 256.663
R1541 B.n857 B.n60 256.663
R1542 B.n857 B.n59 256.663
R1543 B.n857 B.n58 256.663
R1544 B.n857 B.n57 256.663
R1545 B.n857 B.n56 256.663
R1546 B.n857 B.n55 256.663
R1547 B.n857 B.n54 256.663
R1548 B.n857 B.n53 256.663
R1549 B.n857 B.n52 256.663
R1550 B.n857 B.n51 256.663
R1551 B.n857 B.n50 256.663
R1552 B.n857 B.n49 256.663
R1553 B.n857 B.n48 256.663
R1554 B.n857 B.n47 256.663
R1555 B.n857 B.n46 256.663
R1556 B.n857 B.n45 256.663
R1557 B.n857 B.n44 256.663
R1558 B.n857 B.n43 256.663
R1559 B.n857 B.n42 256.663
R1560 B.n857 B.n41 256.663
R1561 B.n858 B.n857 256.663
R1562 B.n767 B.n766 256.663
R1563 B.n766 B.n421 256.663
R1564 B.n766 B.n422 256.663
R1565 B.n766 B.n423 256.663
R1566 B.n766 B.n424 256.663
R1567 B.n766 B.n425 256.663
R1568 B.n766 B.n426 256.663
R1569 B.n766 B.n427 256.663
R1570 B.n766 B.n428 256.663
R1571 B.n766 B.n429 256.663
R1572 B.n766 B.n430 256.663
R1573 B.n766 B.n431 256.663
R1574 B.n766 B.n432 256.663
R1575 B.n766 B.n433 256.663
R1576 B.n766 B.n434 256.663
R1577 B.n766 B.n435 256.663
R1578 B.n766 B.n436 256.663
R1579 B.n766 B.n437 256.663
R1580 B.n766 B.n438 256.663
R1581 B.n766 B.n439 256.663
R1582 B.n766 B.n440 256.663
R1583 B.n766 B.n441 256.663
R1584 B.n766 B.n442 256.663
R1585 B.n766 B.n443 256.663
R1586 B.n766 B.n444 256.663
R1587 B.n766 B.n445 256.663
R1588 B.n766 B.n446 256.663
R1589 B.n766 B.n447 256.663
R1590 B.n766 B.n448 256.663
R1591 B.n766 B.n449 256.663
R1592 B.n766 B.n450 256.663
R1593 B.n766 B.n451 256.663
R1594 B.n766 B.n452 256.663
R1595 B.n766 B.n453 256.663
R1596 B.n766 B.n454 256.663
R1597 B.n766 B.n455 256.663
R1598 B.n766 B.n456 256.663
R1599 B.n766 B.n457 256.663
R1600 B.n766 B.n458 256.663
R1601 B.n766 B.n459 256.663
R1602 B.n766 B.n460 256.663
R1603 B.n766 B.n461 256.663
R1604 B.n766 B.n462 256.663
R1605 B.n766 B.n463 256.663
R1606 B.n766 B.n464 256.663
R1607 B.n766 B.n465 256.663
R1608 B.n766 B.n466 256.663
R1609 B.n766 B.n467 256.663
R1610 B.n766 B.n468 256.663
R1611 B.n766 B.n469 256.663
R1612 B.n766 B.n470 256.663
R1613 B.n766 B.n471 256.663
R1614 B.n766 B.n472 256.663
R1615 B.n766 B.n473 256.663
R1616 B.n766 B.n474 256.663
R1617 B.n766 B.n475 256.663
R1618 B.n766 B.n476 256.663
R1619 B.n766 B.n477 256.663
R1620 B.n766 B.n478 256.663
R1621 B.n766 B.n479 256.663
R1622 B.n766 B.n480 256.663
R1623 B.n766 B.n481 256.663
R1624 B.n766 B.n482 256.663
R1625 B.n766 B.n483 256.663
R1626 B.n766 B.n484 256.663
R1627 B.n766 B.n485 256.663
R1628 B.n766 B.n486 256.663
R1629 B.n766 B.n487 256.663
R1630 B.n902 B.n901 256.663
R1631 B.n116 B.n40 163.367
R1632 B.n120 B.n119 163.367
R1633 B.n124 B.n123 163.367
R1634 B.n128 B.n127 163.367
R1635 B.n132 B.n131 163.367
R1636 B.n136 B.n135 163.367
R1637 B.n140 B.n139 163.367
R1638 B.n144 B.n143 163.367
R1639 B.n148 B.n147 163.367
R1640 B.n152 B.n151 163.367
R1641 B.n156 B.n155 163.367
R1642 B.n160 B.n159 163.367
R1643 B.n164 B.n163 163.367
R1644 B.n168 B.n167 163.367
R1645 B.n172 B.n171 163.367
R1646 B.n176 B.n175 163.367
R1647 B.n180 B.n179 163.367
R1648 B.n184 B.n183 163.367
R1649 B.n188 B.n187 163.367
R1650 B.n192 B.n191 163.367
R1651 B.n196 B.n195 163.367
R1652 B.n200 B.n199 163.367
R1653 B.n204 B.n203 163.367
R1654 B.n208 B.n207 163.367
R1655 B.n212 B.n211 163.367
R1656 B.n216 B.n215 163.367
R1657 B.n220 B.n219 163.367
R1658 B.n224 B.n223 163.367
R1659 B.n228 B.n227 163.367
R1660 B.n232 B.n231 163.367
R1661 B.n236 B.n235 163.367
R1662 B.n240 B.n239 163.367
R1663 B.n244 B.n243 163.367
R1664 B.n248 B.n247 163.367
R1665 B.n252 B.n251 163.367
R1666 B.n256 B.n255 163.367
R1667 B.n260 B.n259 163.367
R1668 B.n264 B.n263 163.367
R1669 B.n268 B.n267 163.367
R1670 B.n272 B.n271 163.367
R1671 B.n276 B.n275 163.367
R1672 B.n280 B.n279 163.367
R1673 B.n284 B.n283 163.367
R1674 B.n288 B.n287 163.367
R1675 B.n292 B.n291 163.367
R1676 B.n296 B.n295 163.367
R1677 B.n300 B.n299 163.367
R1678 B.n304 B.n303 163.367
R1679 B.n308 B.n307 163.367
R1680 B.n312 B.n311 163.367
R1681 B.n316 B.n315 163.367
R1682 B.n320 B.n319 163.367
R1683 B.n324 B.n323 163.367
R1684 B.n328 B.n327 163.367
R1685 B.n332 B.n331 163.367
R1686 B.n336 B.n335 163.367
R1687 B.n340 B.n339 163.367
R1688 B.n344 B.n343 163.367
R1689 B.n348 B.n347 163.367
R1690 B.n352 B.n351 163.367
R1691 B.n356 B.n355 163.367
R1692 B.n360 B.n359 163.367
R1693 B.n364 B.n363 163.367
R1694 B.n368 B.n367 163.367
R1695 B.n372 B.n371 163.367
R1696 B.n376 B.n375 163.367
R1697 B.n380 B.n379 163.367
R1698 B.n382 B.n108 163.367
R1699 B.n774 B.n416 163.367
R1700 B.n774 B.n414 163.367
R1701 B.n778 B.n414 163.367
R1702 B.n778 B.n409 163.367
R1703 B.n787 B.n409 163.367
R1704 B.n787 B.n407 163.367
R1705 B.n791 B.n407 163.367
R1706 B.n791 B.n400 163.367
R1707 B.n799 B.n400 163.367
R1708 B.n799 B.n398 163.367
R1709 B.n803 B.n398 163.367
R1710 B.n803 B.n393 163.367
R1711 B.n811 B.n393 163.367
R1712 B.n811 B.n391 163.367
R1713 B.n816 B.n391 163.367
R1714 B.n816 B.n386 163.367
R1715 B.n825 B.n386 163.367
R1716 B.n826 B.n825 163.367
R1717 B.n826 B.n5 163.367
R1718 B.n6 B.n5 163.367
R1719 B.n7 B.n6 163.367
R1720 B.n832 B.n7 163.367
R1721 B.n833 B.n832 163.367
R1722 B.n833 B.n13 163.367
R1723 B.n14 B.n13 163.367
R1724 B.n15 B.n14 163.367
R1725 B.n838 B.n15 163.367
R1726 B.n838 B.n20 163.367
R1727 B.n21 B.n20 163.367
R1728 B.n22 B.n21 163.367
R1729 B.n843 B.n22 163.367
R1730 B.n843 B.n27 163.367
R1731 B.n28 B.n27 163.367
R1732 B.n29 B.n28 163.367
R1733 B.n848 B.n29 163.367
R1734 B.n848 B.n34 163.367
R1735 B.n35 B.n34 163.367
R1736 B.n36 B.n35 163.367
R1737 B.n109 B.n36 163.367
R1738 B.n765 B.n420 163.367
R1739 B.n765 B.n489 163.367
R1740 B.n761 B.n760 163.367
R1741 B.n757 B.n756 163.367
R1742 B.n753 B.n752 163.367
R1743 B.n749 B.n748 163.367
R1744 B.n745 B.n744 163.367
R1745 B.n741 B.n740 163.367
R1746 B.n737 B.n736 163.367
R1747 B.n733 B.n732 163.367
R1748 B.n729 B.n728 163.367
R1749 B.n725 B.n724 163.367
R1750 B.n721 B.n720 163.367
R1751 B.n717 B.n716 163.367
R1752 B.n713 B.n712 163.367
R1753 B.n709 B.n708 163.367
R1754 B.n705 B.n704 163.367
R1755 B.n701 B.n700 163.367
R1756 B.n697 B.n696 163.367
R1757 B.n693 B.n692 163.367
R1758 B.n689 B.n688 163.367
R1759 B.n685 B.n684 163.367
R1760 B.n681 B.n680 163.367
R1761 B.n677 B.n676 163.367
R1762 B.n673 B.n672 163.367
R1763 B.n669 B.n668 163.367
R1764 B.n665 B.n664 163.367
R1765 B.n661 B.n660 163.367
R1766 B.n657 B.n656 163.367
R1767 B.n653 B.n652 163.367
R1768 B.n649 B.n648 163.367
R1769 B.n645 B.n644 163.367
R1770 B.n640 B.n639 163.367
R1771 B.n636 B.n635 163.367
R1772 B.n632 B.n631 163.367
R1773 B.n628 B.n627 163.367
R1774 B.n624 B.n623 163.367
R1775 B.n619 B.n618 163.367
R1776 B.n615 B.n614 163.367
R1777 B.n611 B.n610 163.367
R1778 B.n607 B.n606 163.367
R1779 B.n603 B.n602 163.367
R1780 B.n599 B.n598 163.367
R1781 B.n595 B.n594 163.367
R1782 B.n591 B.n590 163.367
R1783 B.n587 B.n586 163.367
R1784 B.n583 B.n582 163.367
R1785 B.n579 B.n578 163.367
R1786 B.n575 B.n574 163.367
R1787 B.n571 B.n570 163.367
R1788 B.n567 B.n566 163.367
R1789 B.n563 B.n562 163.367
R1790 B.n559 B.n558 163.367
R1791 B.n555 B.n554 163.367
R1792 B.n551 B.n550 163.367
R1793 B.n547 B.n546 163.367
R1794 B.n543 B.n542 163.367
R1795 B.n539 B.n538 163.367
R1796 B.n535 B.n534 163.367
R1797 B.n531 B.n530 163.367
R1798 B.n527 B.n526 163.367
R1799 B.n523 B.n522 163.367
R1800 B.n519 B.n518 163.367
R1801 B.n515 B.n514 163.367
R1802 B.n511 B.n510 163.367
R1803 B.n507 B.n506 163.367
R1804 B.n503 B.n502 163.367
R1805 B.n499 B.n498 163.367
R1806 B.n495 B.n488 163.367
R1807 B.n772 B.n418 163.367
R1808 B.n772 B.n412 163.367
R1809 B.n781 B.n412 163.367
R1810 B.n781 B.n410 163.367
R1811 B.n785 B.n410 163.367
R1812 B.n785 B.n405 163.367
R1813 B.n793 B.n405 163.367
R1814 B.n793 B.n403 163.367
R1815 B.n797 B.n403 163.367
R1816 B.n797 B.n397 163.367
R1817 B.n805 B.n397 163.367
R1818 B.n805 B.n395 163.367
R1819 B.n809 B.n395 163.367
R1820 B.n809 B.n389 163.367
R1821 B.n819 B.n389 163.367
R1822 B.n819 B.n387 163.367
R1823 B.n823 B.n387 163.367
R1824 B.n823 B.n3 163.367
R1825 B.n900 B.n3 163.367
R1826 B.n896 B.n2 163.367
R1827 B.n896 B.n895 163.367
R1828 B.n895 B.n9 163.367
R1829 B.n891 B.n9 163.367
R1830 B.n891 B.n11 163.367
R1831 B.n887 B.n11 163.367
R1832 B.n887 B.n17 163.367
R1833 B.n883 B.n17 163.367
R1834 B.n883 B.n19 163.367
R1835 B.n879 B.n19 163.367
R1836 B.n879 B.n24 163.367
R1837 B.n875 B.n24 163.367
R1838 B.n875 B.n26 163.367
R1839 B.n871 B.n26 163.367
R1840 B.n871 B.n30 163.367
R1841 B.n867 B.n30 163.367
R1842 B.n867 B.n32 163.367
R1843 B.n863 B.n32 163.367
R1844 B.n863 B.n38 163.367
R1845 B.n859 B.n858 71.676
R1846 B.n116 B.n41 71.676
R1847 B.n120 B.n42 71.676
R1848 B.n124 B.n43 71.676
R1849 B.n128 B.n44 71.676
R1850 B.n132 B.n45 71.676
R1851 B.n136 B.n46 71.676
R1852 B.n140 B.n47 71.676
R1853 B.n144 B.n48 71.676
R1854 B.n148 B.n49 71.676
R1855 B.n152 B.n50 71.676
R1856 B.n156 B.n51 71.676
R1857 B.n160 B.n52 71.676
R1858 B.n164 B.n53 71.676
R1859 B.n168 B.n54 71.676
R1860 B.n172 B.n55 71.676
R1861 B.n176 B.n56 71.676
R1862 B.n180 B.n57 71.676
R1863 B.n184 B.n58 71.676
R1864 B.n188 B.n59 71.676
R1865 B.n192 B.n60 71.676
R1866 B.n196 B.n61 71.676
R1867 B.n200 B.n62 71.676
R1868 B.n204 B.n63 71.676
R1869 B.n208 B.n64 71.676
R1870 B.n212 B.n65 71.676
R1871 B.n216 B.n66 71.676
R1872 B.n220 B.n67 71.676
R1873 B.n224 B.n68 71.676
R1874 B.n228 B.n69 71.676
R1875 B.n232 B.n70 71.676
R1876 B.n236 B.n71 71.676
R1877 B.n240 B.n72 71.676
R1878 B.n244 B.n73 71.676
R1879 B.n248 B.n74 71.676
R1880 B.n252 B.n75 71.676
R1881 B.n256 B.n76 71.676
R1882 B.n260 B.n77 71.676
R1883 B.n264 B.n78 71.676
R1884 B.n268 B.n79 71.676
R1885 B.n272 B.n80 71.676
R1886 B.n276 B.n81 71.676
R1887 B.n280 B.n82 71.676
R1888 B.n284 B.n83 71.676
R1889 B.n288 B.n84 71.676
R1890 B.n292 B.n85 71.676
R1891 B.n296 B.n86 71.676
R1892 B.n300 B.n87 71.676
R1893 B.n304 B.n88 71.676
R1894 B.n308 B.n89 71.676
R1895 B.n312 B.n90 71.676
R1896 B.n316 B.n91 71.676
R1897 B.n320 B.n92 71.676
R1898 B.n324 B.n93 71.676
R1899 B.n328 B.n94 71.676
R1900 B.n332 B.n95 71.676
R1901 B.n336 B.n96 71.676
R1902 B.n340 B.n97 71.676
R1903 B.n344 B.n98 71.676
R1904 B.n348 B.n99 71.676
R1905 B.n352 B.n100 71.676
R1906 B.n356 B.n101 71.676
R1907 B.n360 B.n102 71.676
R1908 B.n364 B.n103 71.676
R1909 B.n368 B.n104 71.676
R1910 B.n372 B.n105 71.676
R1911 B.n376 B.n106 71.676
R1912 B.n380 B.n107 71.676
R1913 B.n856 B.n108 71.676
R1914 B.n856 B.n855 71.676
R1915 B.n382 B.n107 71.676
R1916 B.n379 B.n106 71.676
R1917 B.n375 B.n105 71.676
R1918 B.n371 B.n104 71.676
R1919 B.n367 B.n103 71.676
R1920 B.n363 B.n102 71.676
R1921 B.n359 B.n101 71.676
R1922 B.n355 B.n100 71.676
R1923 B.n351 B.n99 71.676
R1924 B.n347 B.n98 71.676
R1925 B.n343 B.n97 71.676
R1926 B.n339 B.n96 71.676
R1927 B.n335 B.n95 71.676
R1928 B.n331 B.n94 71.676
R1929 B.n327 B.n93 71.676
R1930 B.n323 B.n92 71.676
R1931 B.n319 B.n91 71.676
R1932 B.n315 B.n90 71.676
R1933 B.n311 B.n89 71.676
R1934 B.n307 B.n88 71.676
R1935 B.n303 B.n87 71.676
R1936 B.n299 B.n86 71.676
R1937 B.n295 B.n85 71.676
R1938 B.n291 B.n84 71.676
R1939 B.n287 B.n83 71.676
R1940 B.n283 B.n82 71.676
R1941 B.n279 B.n81 71.676
R1942 B.n275 B.n80 71.676
R1943 B.n271 B.n79 71.676
R1944 B.n267 B.n78 71.676
R1945 B.n263 B.n77 71.676
R1946 B.n259 B.n76 71.676
R1947 B.n255 B.n75 71.676
R1948 B.n251 B.n74 71.676
R1949 B.n247 B.n73 71.676
R1950 B.n243 B.n72 71.676
R1951 B.n239 B.n71 71.676
R1952 B.n235 B.n70 71.676
R1953 B.n231 B.n69 71.676
R1954 B.n227 B.n68 71.676
R1955 B.n223 B.n67 71.676
R1956 B.n219 B.n66 71.676
R1957 B.n215 B.n65 71.676
R1958 B.n211 B.n64 71.676
R1959 B.n207 B.n63 71.676
R1960 B.n203 B.n62 71.676
R1961 B.n199 B.n61 71.676
R1962 B.n195 B.n60 71.676
R1963 B.n191 B.n59 71.676
R1964 B.n187 B.n58 71.676
R1965 B.n183 B.n57 71.676
R1966 B.n179 B.n56 71.676
R1967 B.n175 B.n55 71.676
R1968 B.n171 B.n54 71.676
R1969 B.n167 B.n53 71.676
R1970 B.n163 B.n52 71.676
R1971 B.n159 B.n51 71.676
R1972 B.n155 B.n50 71.676
R1973 B.n151 B.n49 71.676
R1974 B.n147 B.n48 71.676
R1975 B.n143 B.n47 71.676
R1976 B.n139 B.n46 71.676
R1977 B.n135 B.n45 71.676
R1978 B.n131 B.n44 71.676
R1979 B.n127 B.n43 71.676
R1980 B.n123 B.n42 71.676
R1981 B.n119 B.n41 71.676
R1982 B.n858 B.n40 71.676
R1983 B.n768 B.n767 71.676
R1984 B.n489 B.n421 71.676
R1985 B.n760 B.n422 71.676
R1986 B.n756 B.n423 71.676
R1987 B.n752 B.n424 71.676
R1988 B.n748 B.n425 71.676
R1989 B.n744 B.n426 71.676
R1990 B.n740 B.n427 71.676
R1991 B.n736 B.n428 71.676
R1992 B.n732 B.n429 71.676
R1993 B.n728 B.n430 71.676
R1994 B.n724 B.n431 71.676
R1995 B.n720 B.n432 71.676
R1996 B.n716 B.n433 71.676
R1997 B.n712 B.n434 71.676
R1998 B.n708 B.n435 71.676
R1999 B.n704 B.n436 71.676
R2000 B.n700 B.n437 71.676
R2001 B.n696 B.n438 71.676
R2002 B.n692 B.n439 71.676
R2003 B.n688 B.n440 71.676
R2004 B.n684 B.n441 71.676
R2005 B.n680 B.n442 71.676
R2006 B.n676 B.n443 71.676
R2007 B.n672 B.n444 71.676
R2008 B.n668 B.n445 71.676
R2009 B.n664 B.n446 71.676
R2010 B.n660 B.n447 71.676
R2011 B.n656 B.n448 71.676
R2012 B.n652 B.n449 71.676
R2013 B.n648 B.n450 71.676
R2014 B.n644 B.n451 71.676
R2015 B.n639 B.n452 71.676
R2016 B.n635 B.n453 71.676
R2017 B.n631 B.n454 71.676
R2018 B.n627 B.n455 71.676
R2019 B.n623 B.n456 71.676
R2020 B.n618 B.n457 71.676
R2021 B.n614 B.n458 71.676
R2022 B.n610 B.n459 71.676
R2023 B.n606 B.n460 71.676
R2024 B.n602 B.n461 71.676
R2025 B.n598 B.n462 71.676
R2026 B.n594 B.n463 71.676
R2027 B.n590 B.n464 71.676
R2028 B.n586 B.n465 71.676
R2029 B.n582 B.n466 71.676
R2030 B.n578 B.n467 71.676
R2031 B.n574 B.n468 71.676
R2032 B.n570 B.n469 71.676
R2033 B.n566 B.n470 71.676
R2034 B.n562 B.n471 71.676
R2035 B.n558 B.n472 71.676
R2036 B.n554 B.n473 71.676
R2037 B.n550 B.n474 71.676
R2038 B.n546 B.n475 71.676
R2039 B.n542 B.n476 71.676
R2040 B.n538 B.n477 71.676
R2041 B.n534 B.n478 71.676
R2042 B.n530 B.n479 71.676
R2043 B.n526 B.n480 71.676
R2044 B.n522 B.n481 71.676
R2045 B.n518 B.n482 71.676
R2046 B.n514 B.n483 71.676
R2047 B.n510 B.n484 71.676
R2048 B.n506 B.n485 71.676
R2049 B.n502 B.n486 71.676
R2050 B.n498 B.n487 71.676
R2051 B.n767 B.n420 71.676
R2052 B.n761 B.n421 71.676
R2053 B.n757 B.n422 71.676
R2054 B.n753 B.n423 71.676
R2055 B.n749 B.n424 71.676
R2056 B.n745 B.n425 71.676
R2057 B.n741 B.n426 71.676
R2058 B.n737 B.n427 71.676
R2059 B.n733 B.n428 71.676
R2060 B.n729 B.n429 71.676
R2061 B.n725 B.n430 71.676
R2062 B.n721 B.n431 71.676
R2063 B.n717 B.n432 71.676
R2064 B.n713 B.n433 71.676
R2065 B.n709 B.n434 71.676
R2066 B.n705 B.n435 71.676
R2067 B.n701 B.n436 71.676
R2068 B.n697 B.n437 71.676
R2069 B.n693 B.n438 71.676
R2070 B.n689 B.n439 71.676
R2071 B.n685 B.n440 71.676
R2072 B.n681 B.n441 71.676
R2073 B.n677 B.n442 71.676
R2074 B.n673 B.n443 71.676
R2075 B.n669 B.n444 71.676
R2076 B.n665 B.n445 71.676
R2077 B.n661 B.n446 71.676
R2078 B.n657 B.n447 71.676
R2079 B.n653 B.n448 71.676
R2080 B.n649 B.n449 71.676
R2081 B.n645 B.n450 71.676
R2082 B.n640 B.n451 71.676
R2083 B.n636 B.n452 71.676
R2084 B.n632 B.n453 71.676
R2085 B.n628 B.n454 71.676
R2086 B.n624 B.n455 71.676
R2087 B.n619 B.n456 71.676
R2088 B.n615 B.n457 71.676
R2089 B.n611 B.n458 71.676
R2090 B.n607 B.n459 71.676
R2091 B.n603 B.n460 71.676
R2092 B.n599 B.n461 71.676
R2093 B.n595 B.n462 71.676
R2094 B.n591 B.n463 71.676
R2095 B.n587 B.n464 71.676
R2096 B.n583 B.n465 71.676
R2097 B.n579 B.n466 71.676
R2098 B.n575 B.n467 71.676
R2099 B.n571 B.n468 71.676
R2100 B.n567 B.n469 71.676
R2101 B.n563 B.n470 71.676
R2102 B.n559 B.n471 71.676
R2103 B.n555 B.n472 71.676
R2104 B.n551 B.n473 71.676
R2105 B.n547 B.n474 71.676
R2106 B.n543 B.n475 71.676
R2107 B.n539 B.n476 71.676
R2108 B.n535 B.n477 71.676
R2109 B.n531 B.n478 71.676
R2110 B.n527 B.n479 71.676
R2111 B.n523 B.n480 71.676
R2112 B.n519 B.n481 71.676
R2113 B.n515 B.n482 71.676
R2114 B.n511 B.n483 71.676
R2115 B.n507 B.n484 71.676
R2116 B.n503 B.n485 71.676
R2117 B.n499 B.n486 71.676
R2118 B.n495 B.n487 71.676
R2119 B.n901 B.n900 71.676
R2120 B.n901 B.n2 71.676
R2121 B.n766 B.n417 62.2272
R2122 B.n857 B.n37 62.2272
R2123 B.n115 B.n114 59.5399
R2124 B.n112 B.n111 59.5399
R2125 B.n621 B.n493 59.5399
R2126 B.n642 B.n491 59.5399
R2127 B.n770 B.n769 34.1859
R2128 B.n494 B.n415 34.1859
R2129 B.n854 B.n853 34.1859
R2130 B.n861 B.n860 34.1859
R2131 B.n773 B.n417 30.0105
R2132 B.n773 B.n413 30.0105
R2133 B.n780 B.n413 30.0105
R2134 B.n780 B.n779 30.0105
R2135 B.n786 B.n406 30.0105
R2136 B.n792 B.n406 30.0105
R2137 B.n792 B.n401 30.0105
R2138 B.n798 B.n401 30.0105
R2139 B.n798 B.n402 30.0105
R2140 B.n804 B.n394 30.0105
R2141 B.n810 B.n394 30.0105
R2142 B.n818 B.n390 30.0105
R2143 B.n818 B.n817 30.0105
R2144 B.n824 B.n4 30.0105
R2145 B.n899 B.n4 30.0105
R2146 B.n899 B.n898 30.0105
R2147 B.n898 B.n897 30.0105
R2148 B.n897 B.n8 30.0105
R2149 B.n890 B.n12 30.0105
R2150 B.n890 B.n889 30.0105
R2151 B.n888 B.n16 30.0105
R2152 B.n882 B.n16 30.0105
R2153 B.n881 B.n880 30.0105
R2154 B.n880 B.n23 30.0105
R2155 B.n874 B.n23 30.0105
R2156 B.n874 B.n873 30.0105
R2157 B.n873 B.n872 30.0105
R2158 B.n866 B.n33 30.0105
R2159 B.n866 B.n865 30.0105
R2160 B.n865 B.n864 30.0105
R2161 B.n864 B.n37 30.0105
R2162 B.n114 B.n113 19.2005
R2163 B.n111 B.n110 19.2005
R2164 B.n493 B.n492 19.2005
R2165 B.n491 B.n490 19.2005
R2166 B.n402 B.t1 18.5361
R2167 B.t4 B.n881 18.5361
R2168 B B.n902 18.0485
R2169 B.n824 B.t2 16.7708
R2170 B.t5 B.n8 16.7708
R2171 B.n810 B.t0 15.8882
R2172 B.t3 B.n888 15.8882
R2173 B.n779 B.t7 15.0055
R2174 B.n786 B.t7 15.0055
R2175 B.n872 B.t11 15.0055
R2176 B.n33 B.t11 15.0055
R2177 B.t0 B.n390 14.1229
R2178 B.n889 B.t3 14.1229
R2179 B.n817 B.t2 13.2402
R2180 B.n12 B.t5 13.2402
R2181 B.n804 B.t1 11.4749
R2182 B.n882 B.t4 11.4749
R2183 B.n771 B.n770 10.6151
R2184 B.n771 B.n411 10.6151
R2185 B.n782 B.n411 10.6151
R2186 B.n783 B.n782 10.6151
R2187 B.n784 B.n783 10.6151
R2188 B.n784 B.n404 10.6151
R2189 B.n794 B.n404 10.6151
R2190 B.n795 B.n794 10.6151
R2191 B.n796 B.n795 10.6151
R2192 B.n796 B.n396 10.6151
R2193 B.n806 B.n396 10.6151
R2194 B.n807 B.n806 10.6151
R2195 B.n808 B.n807 10.6151
R2196 B.n808 B.n388 10.6151
R2197 B.n820 B.n388 10.6151
R2198 B.n821 B.n820 10.6151
R2199 B.n822 B.n821 10.6151
R2200 B.n822 B.n0 10.6151
R2201 B.n769 B.n419 10.6151
R2202 B.n764 B.n419 10.6151
R2203 B.n764 B.n763 10.6151
R2204 B.n763 B.n762 10.6151
R2205 B.n762 B.n759 10.6151
R2206 B.n759 B.n758 10.6151
R2207 B.n758 B.n755 10.6151
R2208 B.n755 B.n754 10.6151
R2209 B.n754 B.n751 10.6151
R2210 B.n751 B.n750 10.6151
R2211 B.n750 B.n747 10.6151
R2212 B.n747 B.n746 10.6151
R2213 B.n746 B.n743 10.6151
R2214 B.n743 B.n742 10.6151
R2215 B.n742 B.n739 10.6151
R2216 B.n739 B.n738 10.6151
R2217 B.n738 B.n735 10.6151
R2218 B.n735 B.n734 10.6151
R2219 B.n734 B.n731 10.6151
R2220 B.n731 B.n730 10.6151
R2221 B.n730 B.n727 10.6151
R2222 B.n727 B.n726 10.6151
R2223 B.n726 B.n723 10.6151
R2224 B.n723 B.n722 10.6151
R2225 B.n722 B.n719 10.6151
R2226 B.n719 B.n718 10.6151
R2227 B.n718 B.n715 10.6151
R2228 B.n715 B.n714 10.6151
R2229 B.n714 B.n711 10.6151
R2230 B.n711 B.n710 10.6151
R2231 B.n710 B.n707 10.6151
R2232 B.n707 B.n706 10.6151
R2233 B.n706 B.n703 10.6151
R2234 B.n703 B.n702 10.6151
R2235 B.n702 B.n699 10.6151
R2236 B.n699 B.n698 10.6151
R2237 B.n698 B.n695 10.6151
R2238 B.n695 B.n694 10.6151
R2239 B.n694 B.n691 10.6151
R2240 B.n691 B.n690 10.6151
R2241 B.n690 B.n687 10.6151
R2242 B.n687 B.n686 10.6151
R2243 B.n686 B.n683 10.6151
R2244 B.n683 B.n682 10.6151
R2245 B.n682 B.n679 10.6151
R2246 B.n679 B.n678 10.6151
R2247 B.n678 B.n675 10.6151
R2248 B.n675 B.n674 10.6151
R2249 B.n674 B.n671 10.6151
R2250 B.n671 B.n670 10.6151
R2251 B.n670 B.n667 10.6151
R2252 B.n667 B.n666 10.6151
R2253 B.n666 B.n663 10.6151
R2254 B.n663 B.n662 10.6151
R2255 B.n662 B.n659 10.6151
R2256 B.n659 B.n658 10.6151
R2257 B.n658 B.n655 10.6151
R2258 B.n655 B.n654 10.6151
R2259 B.n654 B.n651 10.6151
R2260 B.n651 B.n650 10.6151
R2261 B.n650 B.n647 10.6151
R2262 B.n647 B.n646 10.6151
R2263 B.n646 B.n643 10.6151
R2264 B.n641 B.n638 10.6151
R2265 B.n638 B.n637 10.6151
R2266 B.n637 B.n634 10.6151
R2267 B.n634 B.n633 10.6151
R2268 B.n633 B.n630 10.6151
R2269 B.n630 B.n629 10.6151
R2270 B.n629 B.n626 10.6151
R2271 B.n626 B.n625 10.6151
R2272 B.n625 B.n622 10.6151
R2273 B.n620 B.n617 10.6151
R2274 B.n617 B.n616 10.6151
R2275 B.n616 B.n613 10.6151
R2276 B.n613 B.n612 10.6151
R2277 B.n612 B.n609 10.6151
R2278 B.n609 B.n608 10.6151
R2279 B.n608 B.n605 10.6151
R2280 B.n605 B.n604 10.6151
R2281 B.n604 B.n601 10.6151
R2282 B.n601 B.n600 10.6151
R2283 B.n600 B.n597 10.6151
R2284 B.n597 B.n596 10.6151
R2285 B.n596 B.n593 10.6151
R2286 B.n593 B.n592 10.6151
R2287 B.n592 B.n589 10.6151
R2288 B.n589 B.n588 10.6151
R2289 B.n588 B.n585 10.6151
R2290 B.n585 B.n584 10.6151
R2291 B.n584 B.n581 10.6151
R2292 B.n581 B.n580 10.6151
R2293 B.n580 B.n577 10.6151
R2294 B.n577 B.n576 10.6151
R2295 B.n576 B.n573 10.6151
R2296 B.n573 B.n572 10.6151
R2297 B.n572 B.n569 10.6151
R2298 B.n569 B.n568 10.6151
R2299 B.n568 B.n565 10.6151
R2300 B.n565 B.n564 10.6151
R2301 B.n564 B.n561 10.6151
R2302 B.n561 B.n560 10.6151
R2303 B.n560 B.n557 10.6151
R2304 B.n557 B.n556 10.6151
R2305 B.n556 B.n553 10.6151
R2306 B.n553 B.n552 10.6151
R2307 B.n552 B.n549 10.6151
R2308 B.n549 B.n548 10.6151
R2309 B.n548 B.n545 10.6151
R2310 B.n545 B.n544 10.6151
R2311 B.n544 B.n541 10.6151
R2312 B.n541 B.n540 10.6151
R2313 B.n540 B.n537 10.6151
R2314 B.n537 B.n536 10.6151
R2315 B.n536 B.n533 10.6151
R2316 B.n533 B.n532 10.6151
R2317 B.n532 B.n529 10.6151
R2318 B.n529 B.n528 10.6151
R2319 B.n528 B.n525 10.6151
R2320 B.n525 B.n524 10.6151
R2321 B.n524 B.n521 10.6151
R2322 B.n521 B.n520 10.6151
R2323 B.n520 B.n517 10.6151
R2324 B.n517 B.n516 10.6151
R2325 B.n516 B.n513 10.6151
R2326 B.n513 B.n512 10.6151
R2327 B.n512 B.n509 10.6151
R2328 B.n509 B.n508 10.6151
R2329 B.n508 B.n505 10.6151
R2330 B.n505 B.n504 10.6151
R2331 B.n504 B.n501 10.6151
R2332 B.n501 B.n500 10.6151
R2333 B.n500 B.n497 10.6151
R2334 B.n497 B.n496 10.6151
R2335 B.n496 B.n494 10.6151
R2336 B.n775 B.n415 10.6151
R2337 B.n776 B.n775 10.6151
R2338 B.n777 B.n776 10.6151
R2339 B.n777 B.n408 10.6151
R2340 B.n788 B.n408 10.6151
R2341 B.n789 B.n788 10.6151
R2342 B.n790 B.n789 10.6151
R2343 B.n790 B.n399 10.6151
R2344 B.n800 B.n399 10.6151
R2345 B.n801 B.n800 10.6151
R2346 B.n802 B.n801 10.6151
R2347 B.n802 B.n392 10.6151
R2348 B.n812 B.n392 10.6151
R2349 B.n813 B.n812 10.6151
R2350 B.n815 B.n813 10.6151
R2351 B.n815 B.n814 10.6151
R2352 B.n814 B.n385 10.6151
R2353 B.n827 B.n385 10.6151
R2354 B.n828 B.n827 10.6151
R2355 B.n829 B.n828 10.6151
R2356 B.n830 B.n829 10.6151
R2357 B.n831 B.n830 10.6151
R2358 B.n834 B.n831 10.6151
R2359 B.n835 B.n834 10.6151
R2360 B.n836 B.n835 10.6151
R2361 B.n837 B.n836 10.6151
R2362 B.n839 B.n837 10.6151
R2363 B.n840 B.n839 10.6151
R2364 B.n841 B.n840 10.6151
R2365 B.n842 B.n841 10.6151
R2366 B.n844 B.n842 10.6151
R2367 B.n845 B.n844 10.6151
R2368 B.n846 B.n845 10.6151
R2369 B.n847 B.n846 10.6151
R2370 B.n849 B.n847 10.6151
R2371 B.n850 B.n849 10.6151
R2372 B.n851 B.n850 10.6151
R2373 B.n852 B.n851 10.6151
R2374 B.n853 B.n852 10.6151
R2375 B.n894 B.n1 10.6151
R2376 B.n894 B.n893 10.6151
R2377 B.n893 B.n892 10.6151
R2378 B.n892 B.n10 10.6151
R2379 B.n886 B.n10 10.6151
R2380 B.n886 B.n885 10.6151
R2381 B.n885 B.n884 10.6151
R2382 B.n884 B.n18 10.6151
R2383 B.n878 B.n18 10.6151
R2384 B.n878 B.n877 10.6151
R2385 B.n877 B.n876 10.6151
R2386 B.n876 B.n25 10.6151
R2387 B.n870 B.n25 10.6151
R2388 B.n870 B.n869 10.6151
R2389 B.n869 B.n868 10.6151
R2390 B.n868 B.n31 10.6151
R2391 B.n862 B.n31 10.6151
R2392 B.n862 B.n861 10.6151
R2393 B.n860 B.n39 10.6151
R2394 B.n117 B.n39 10.6151
R2395 B.n118 B.n117 10.6151
R2396 B.n121 B.n118 10.6151
R2397 B.n122 B.n121 10.6151
R2398 B.n125 B.n122 10.6151
R2399 B.n126 B.n125 10.6151
R2400 B.n129 B.n126 10.6151
R2401 B.n130 B.n129 10.6151
R2402 B.n133 B.n130 10.6151
R2403 B.n134 B.n133 10.6151
R2404 B.n137 B.n134 10.6151
R2405 B.n138 B.n137 10.6151
R2406 B.n141 B.n138 10.6151
R2407 B.n142 B.n141 10.6151
R2408 B.n145 B.n142 10.6151
R2409 B.n146 B.n145 10.6151
R2410 B.n149 B.n146 10.6151
R2411 B.n150 B.n149 10.6151
R2412 B.n153 B.n150 10.6151
R2413 B.n154 B.n153 10.6151
R2414 B.n157 B.n154 10.6151
R2415 B.n158 B.n157 10.6151
R2416 B.n161 B.n158 10.6151
R2417 B.n162 B.n161 10.6151
R2418 B.n165 B.n162 10.6151
R2419 B.n166 B.n165 10.6151
R2420 B.n169 B.n166 10.6151
R2421 B.n170 B.n169 10.6151
R2422 B.n173 B.n170 10.6151
R2423 B.n174 B.n173 10.6151
R2424 B.n177 B.n174 10.6151
R2425 B.n178 B.n177 10.6151
R2426 B.n181 B.n178 10.6151
R2427 B.n182 B.n181 10.6151
R2428 B.n185 B.n182 10.6151
R2429 B.n186 B.n185 10.6151
R2430 B.n189 B.n186 10.6151
R2431 B.n190 B.n189 10.6151
R2432 B.n193 B.n190 10.6151
R2433 B.n194 B.n193 10.6151
R2434 B.n197 B.n194 10.6151
R2435 B.n198 B.n197 10.6151
R2436 B.n201 B.n198 10.6151
R2437 B.n202 B.n201 10.6151
R2438 B.n205 B.n202 10.6151
R2439 B.n206 B.n205 10.6151
R2440 B.n209 B.n206 10.6151
R2441 B.n210 B.n209 10.6151
R2442 B.n213 B.n210 10.6151
R2443 B.n214 B.n213 10.6151
R2444 B.n217 B.n214 10.6151
R2445 B.n218 B.n217 10.6151
R2446 B.n221 B.n218 10.6151
R2447 B.n222 B.n221 10.6151
R2448 B.n225 B.n222 10.6151
R2449 B.n226 B.n225 10.6151
R2450 B.n229 B.n226 10.6151
R2451 B.n230 B.n229 10.6151
R2452 B.n233 B.n230 10.6151
R2453 B.n234 B.n233 10.6151
R2454 B.n237 B.n234 10.6151
R2455 B.n238 B.n237 10.6151
R2456 B.n242 B.n241 10.6151
R2457 B.n245 B.n242 10.6151
R2458 B.n246 B.n245 10.6151
R2459 B.n249 B.n246 10.6151
R2460 B.n250 B.n249 10.6151
R2461 B.n253 B.n250 10.6151
R2462 B.n254 B.n253 10.6151
R2463 B.n257 B.n254 10.6151
R2464 B.n258 B.n257 10.6151
R2465 B.n262 B.n261 10.6151
R2466 B.n265 B.n262 10.6151
R2467 B.n266 B.n265 10.6151
R2468 B.n269 B.n266 10.6151
R2469 B.n270 B.n269 10.6151
R2470 B.n273 B.n270 10.6151
R2471 B.n274 B.n273 10.6151
R2472 B.n277 B.n274 10.6151
R2473 B.n278 B.n277 10.6151
R2474 B.n281 B.n278 10.6151
R2475 B.n282 B.n281 10.6151
R2476 B.n285 B.n282 10.6151
R2477 B.n286 B.n285 10.6151
R2478 B.n289 B.n286 10.6151
R2479 B.n290 B.n289 10.6151
R2480 B.n293 B.n290 10.6151
R2481 B.n294 B.n293 10.6151
R2482 B.n297 B.n294 10.6151
R2483 B.n298 B.n297 10.6151
R2484 B.n301 B.n298 10.6151
R2485 B.n302 B.n301 10.6151
R2486 B.n305 B.n302 10.6151
R2487 B.n306 B.n305 10.6151
R2488 B.n309 B.n306 10.6151
R2489 B.n310 B.n309 10.6151
R2490 B.n313 B.n310 10.6151
R2491 B.n314 B.n313 10.6151
R2492 B.n317 B.n314 10.6151
R2493 B.n318 B.n317 10.6151
R2494 B.n321 B.n318 10.6151
R2495 B.n322 B.n321 10.6151
R2496 B.n325 B.n322 10.6151
R2497 B.n326 B.n325 10.6151
R2498 B.n329 B.n326 10.6151
R2499 B.n330 B.n329 10.6151
R2500 B.n333 B.n330 10.6151
R2501 B.n334 B.n333 10.6151
R2502 B.n337 B.n334 10.6151
R2503 B.n338 B.n337 10.6151
R2504 B.n341 B.n338 10.6151
R2505 B.n342 B.n341 10.6151
R2506 B.n345 B.n342 10.6151
R2507 B.n346 B.n345 10.6151
R2508 B.n349 B.n346 10.6151
R2509 B.n350 B.n349 10.6151
R2510 B.n353 B.n350 10.6151
R2511 B.n354 B.n353 10.6151
R2512 B.n357 B.n354 10.6151
R2513 B.n358 B.n357 10.6151
R2514 B.n361 B.n358 10.6151
R2515 B.n362 B.n361 10.6151
R2516 B.n365 B.n362 10.6151
R2517 B.n366 B.n365 10.6151
R2518 B.n369 B.n366 10.6151
R2519 B.n370 B.n369 10.6151
R2520 B.n373 B.n370 10.6151
R2521 B.n374 B.n373 10.6151
R2522 B.n377 B.n374 10.6151
R2523 B.n378 B.n377 10.6151
R2524 B.n381 B.n378 10.6151
R2525 B.n383 B.n381 10.6151
R2526 B.n384 B.n383 10.6151
R2527 B.n854 B.n384 10.6151
R2528 B.n643 B.n642 9.36635
R2529 B.n621 B.n620 9.36635
R2530 B.n238 B.n115 9.36635
R2531 B.n261 B.n112 9.36635
R2532 B.n902 B.n0 8.11757
R2533 B.n902 B.n1 8.11757
R2534 B.n642 B.n641 1.24928
R2535 B.n622 B.n621 1.24928
R2536 B.n241 B.n115 1.24928
R2537 B.n258 B.n112 1.24928
R2538 VP.n3 VP.t3 798.202
R2539 VP.n8 VP.t1 777.409
R2540 VP.n12 VP.t2 777.409
R2541 VP.n14 VP.t0 777.409
R2542 VP.n6 VP.t5 777.409
R2543 VP.n4 VP.t4 777.409
R2544 VP.n15 VP.n14 161.3
R2545 VP.n5 VP.n2 161.3
R2546 VP.n7 VP.n6 161.3
R2547 VP.n13 VP.n0 161.3
R2548 VP.n12 VP.n11 161.3
R2549 VP.n10 VP.n1 161.3
R2550 VP.n9 VP.n8 161.3
R2551 VP.n9 VP.n7 46.7997
R2552 VP.n3 VP.n2 44.8515
R2553 VP.n12 VP.n1 24.8308
R2554 VP.n13 VP.n12 24.8308
R2555 VP.n5 VP.n4 24.8308
R2556 VP.n8 VP.n1 23.3702
R2557 VP.n14 VP.n13 23.3702
R2558 VP.n6 VP.n5 23.3702
R2559 VP.n4 VP.n3 21.148
R2560 VP.n7 VP.n2 0.189894
R2561 VP.n10 VP.n9 0.189894
R2562 VP.n11 VP.n10 0.189894
R2563 VP.n11 VP.n0 0.189894
R2564 VP.n15 VP.n0 0.189894
R2565 VP VP.n15 0.0516364
R2566 VDD1.n104 VDD1.n0 289.615
R2567 VDD1.n213 VDD1.n109 289.615
R2568 VDD1.n105 VDD1.n104 185
R2569 VDD1.n103 VDD1.n102 185
R2570 VDD1.n4 VDD1.n3 185
R2571 VDD1.n97 VDD1.n96 185
R2572 VDD1.n95 VDD1.n94 185
R2573 VDD1.n8 VDD1.n7 185
R2574 VDD1.n89 VDD1.n88 185
R2575 VDD1.n87 VDD1.n86 185
R2576 VDD1.n12 VDD1.n11 185
R2577 VDD1.n16 VDD1.n14 185
R2578 VDD1.n81 VDD1.n80 185
R2579 VDD1.n79 VDD1.n78 185
R2580 VDD1.n18 VDD1.n17 185
R2581 VDD1.n73 VDD1.n72 185
R2582 VDD1.n71 VDD1.n70 185
R2583 VDD1.n22 VDD1.n21 185
R2584 VDD1.n65 VDD1.n64 185
R2585 VDD1.n63 VDD1.n62 185
R2586 VDD1.n26 VDD1.n25 185
R2587 VDD1.n57 VDD1.n56 185
R2588 VDD1.n55 VDD1.n54 185
R2589 VDD1.n30 VDD1.n29 185
R2590 VDD1.n49 VDD1.n48 185
R2591 VDD1.n47 VDD1.n46 185
R2592 VDD1.n34 VDD1.n33 185
R2593 VDD1.n41 VDD1.n40 185
R2594 VDD1.n39 VDD1.n38 185
R2595 VDD1.n146 VDD1.n145 185
R2596 VDD1.n148 VDD1.n147 185
R2597 VDD1.n141 VDD1.n140 185
R2598 VDD1.n154 VDD1.n153 185
R2599 VDD1.n156 VDD1.n155 185
R2600 VDD1.n137 VDD1.n136 185
R2601 VDD1.n162 VDD1.n161 185
R2602 VDD1.n164 VDD1.n163 185
R2603 VDD1.n133 VDD1.n132 185
R2604 VDD1.n170 VDD1.n169 185
R2605 VDD1.n172 VDD1.n171 185
R2606 VDD1.n129 VDD1.n128 185
R2607 VDD1.n178 VDD1.n177 185
R2608 VDD1.n180 VDD1.n179 185
R2609 VDD1.n125 VDD1.n124 185
R2610 VDD1.n187 VDD1.n186 185
R2611 VDD1.n188 VDD1.n123 185
R2612 VDD1.n190 VDD1.n189 185
R2613 VDD1.n121 VDD1.n120 185
R2614 VDD1.n196 VDD1.n195 185
R2615 VDD1.n198 VDD1.n197 185
R2616 VDD1.n117 VDD1.n116 185
R2617 VDD1.n204 VDD1.n203 185
R2618 VDD1.n206 VDD1.n205 185
R2619 VDD1.n113 VDD1.n112 185
R2620 VDD1.n212 VDD1.n211 185
R2621 VDD1.n214 VDD1.n213 185
R2622 VDD1.n37 VDD1.t2 147.659
R2623 VDD1.n144 VDD1.t4 147.659
R2624 VDD1.n104 VDD1.n103 104.615
R2625 VDD1.n103 VDD1.n3 104.615
R2626 VDD1.n96 VDD1.n3 104.615
R2627 VDD1.n96 VDD1.n95 104.615
R2628 VDD1.n95 VDD1.n7 104.615
R2629 VDD1.n88 VDD1.n7 104.615
R2630 VDD1.n88 VDD1.n87 104.615
R2631 VDD1.n87 VDD1.n11 104.615
R2632 VDD1.n16 VDD1.n11 104.615
R2633 VDD1.n80 VDD1.n16 104.615
R2634 VDD1.n80 VDD1.n79 104.615
R2635 VDD1.n79 VDD1.n17 104.615
R2636 VDD1.n72 VDD1.n17 104.615
R2637 VDD1.n72 VDD1.n71 104.615
R2638 VDD1.n71 VDD1.n21 104.615
R2639 VDD1.n64 VDD1.n21 104.615
R2640 VDD1.n64 VDD1.n63 104.615
R2641 VDD1.n63 VDD1.n25 104.615
R2642 VDD1.n56 VDD1.n25 104.615
R2643 VDD1.n56 VDD1.n55 104.615
R2644 VDD1.n55 VDD1.n29 104.615
R2645 VDD1.n48 VDD1.n29 104.615
R2646 VDD1.n48 VDD1.n47 104.615
R2647 VDD1.n47 VDD1.n33 104.615
R2648 VDD1.n40 VDD1.n33 104.615
R2649 VDD1.n40 VDD1.n39 104.615
R2650 VDD1.n147 VDD1.n146 104.615
R2651 VDD1.n147 VDD1.n140 104.615
R2652 VDD1.n154 VDD1.n140 104.615
R2653 VDD1.n155 VDD1.n154 104.615
R2654 VDD1.n155 VDD1.n136 104.615
R2655 VDD1.n162 VDD1.n136 104.615
R2656 VDD1.n163 VDD1.n162 104.615
R2657 VDD1.n163 VDD1.n132 104.615
R2658 VDD1.n170 VDD1.n132 104.615
R2659 VDD1.n171 VDD1.n170 104.615
R2660 VDD1.n171 VDD1.n128 104.615
R2661 VDD1.n178 VDD1.n128 104.615
R2662 VDD1.n179 VDD1.n178 104.615
R2663 VDD1.n179 VDD1.n124 104.615
R2664 VDD1.n187 VDD1.n124 104.615
R2665 VDD1.n188 VDD1.n187 104.615
R2666 VDD1.n189 VDD1.n188 104.615
R2667 VDD1.n189 VDD1.n120 104.615
R2668 VDD1.n196 VDD1.n120 104.615
R2669 VDD1.n197 VDD1.n196 104.615
R2670 VDD1.n197 VDD1.n116 104.615
R2671 VDD1.n204 VDD1.n116 104.615
R2672 VDD1.n205 VDD1.n204 104.615
R2673 VDD1.n205 VDD1.n112 104.615
R2674 VDD1.n212 VDD1.n112 104.615
R2675 VDD1.n213 VDD1.n212 104.615
R2676 VDD1.n219 VDD1.n218 60.1782
R2677 VDD1.n221 VDD1.n220 60.0202
R2678 VDD1.n39 VDD1.t2 52.3082
R2679 VDD1.n146 VDD1.t4 52.3082
R2680 VDD1 VDD1.n108 48.9806
R2681 VDD1.n219 VDD1.n217 48.8671
R2682 VDD1.n221 VDD1.n219 44.4384
R2683 VDD1.n38 VDD1.n37 15.6677
R2684 VDD1.n145 VDD1.n144 15.6677
R2685 VDD1.n14 VDD1.n12 13.1884
R2686 VDD1.n190 VDD1.n121 13.1884
R2687 VDD1.n86 VDD1.n85 12.8005
R2688 VDD1.n82 VDD1.n81 12.8005
R2689 VDD1.n41 VDD1.n36 12.8005
R2690 VDD1.n148 VDD1.n143 12.8005
R2691 VDD1.n191 VDD1.n123 12.8005
R2692 VDD1.n195 VDD1.n194 12.8005
R2693 VDD1.n89 VDD1.n10 12.0247
R2694 VDD1.n78 VDD1.n15 12.0247
R2695 VDD1.n42 VDD1.n34 12.0247
R2696 VDD1.n149 VDD1.n141 12.0247
R2697 VDD1.n186 VDD1.n185 12.0247
R2698 VDD1.n198 VDD1.n119 12.0247
R2699 VDD1.n90 VDD1.n8 11.249
R2700 VDD1.n77 VDD1.n18 11.249
R2701 VDD1.n46 VDD1.n45 11.249
R2702 VDD1.n153 VDD1.n152 11.249
R2703 VDD1.n184 VDD1.n125 11.249
R2704 VDD1.n199 VDD1.n117 11.249
R2705 VDD1.n94 VDD1.n93 10.4732
R2706 VDD1.n74 VDD1.n73 10.4732
R2707 VDD1.n49 VDD1.n32 10.4732
R2708 VDD1.n156 VDD1.n139 10.4732
R2709 VDD1.n181 VDD1.n180 10.4732
R2710 VDD1.n203 VDD1.n202 10.4732
R2711 VDD1.n97 VDD1.n6 9.69747
R2712 VDD1.n70 VDD1.n20 9.69747
R2713 VDD1.n50 VDD1.n30 9.69747
R2714 VDD1.n157 VDD1.n137 9.69747
R2715 VDD1.n177 VDD1.n127 9.69747
R2716 VDD1.n206 VDD1.n115 9.69747
R2717 VDD1.n108 VDD1.n107 9.45567
R2718 VDD1.n217 VDD1.n216 9.45567
R2719 VDD1.n24 VDD1.n23 9.3005
R2720 VDD1.n67 VDD1.n66 9.3005
R2721 VDD1.n69 VDD1.n68 9.3005
R2722 VDD1.n20 VDD1.n19 9.3005
R2723 VDD1.n75 VDD1.n74 9.3005
R2724 VDD1.n77 VDD1.n76 9.3005
R2725 VDD1.n15 VDD1.n13 9.3005
R2726 VDD1.n83 VDD1.n82 9.3005
R2727 VDD1.n107 VDD1.n106 9.3005
R2728 VDD1.n2 VDD1.n1 9.3005
R2729 VDD1.n101 VDD1.n100 9.3005
R2730 VDD1.n99 VDD1.n98 9.3005
R2731 VDD1.n6 VDD1.n5 9.3005
R2732 VDD1.n93 VDD1.n92 9.3005
R2733 VDD1.n91 VDD1.n90 9.3005
R2734 VDD1.n10 VDD1.n9 9.3005
R2735 VDD1.n85 VDD1.n84 9.3005
R2736 VDD1.n61 VDD1.n60 9.3005
R2737 VDD1.n59 VDD1.n58 9.3005
R2738 VDD1.n28 VDD1.n27 9.3005
R2739 VDD1.n53 VDD1.n52 9.3005
R2740 VDD1.n51 VDD1.n50 9.3005
R2741 VDD1.n32 VDD1.n31 9.3005
R2742 VDD1.n45 VDD1.n44 9.3005
R2743 VDD1.n43 VDD1.n42 9.3005
R2744 VDD1.n36 VDD1.n35 9.3005
R2745 VDD1.n216 VDD1.n215 9.3005
R2746 VDD1.n210 VDD1.n209 9.3005
R2747 VDD1.n208 VDD1.n207 9.3005
R2748 VDD1.n115 VDD1.n114 9.3005
R2749 VDD1.n202 VDD1.n201 9.3005
R2750 VDD1.n200 VDD1.n199 9.3005
R2751 VDD1.n119 VDD1.n118 9.3005
R2752 VDD1.n194 VDD1.n193 9.3005
R2753 VDD1.n166 VDD1.n165 9.3005
R2754 VDD1.n135 VDD1.n134 9.3005
R2755 VDD1.n160 VDD1.n159 9.3005
R2756 VDD1.n158 VDD1.n157 9.3005
R2757 VDD1.n139 VDD1.n138 9.3005
R2758 VDD1.n152 VDD1.n151 9.3005
R2759 VDD1.n150 VDD1.n149 9.3005
R2760 VDD1.n143 VDD1.n142 9.3005
R2761 VDD1.n168 VDD1.n167 9.3005
R2762 VDD1.n131 VDD1.n130 9.3005
R2763 VDD1.n174 VDD1.n173 9.3005
R2764 VDD1.n176 VDD1.n175 9.3005
R2765 VDD1.n127 VDD1.n126 9.3005
R2766 VDD1.n182 VDD1.n181 9.3005
R2767 VDD1.n184 VDD1.n183 9.3005
R2768 VDD1.n185 VDD1.n122 9.3005
R2769 VDD1.n192 VDD1.n191 9.3005
R2770 VDD1.n111 VDD1.n110 9.3005
R2771 VDD1.n98 VDD1.n4 8.92171
R2772 VDD1.n69 VDD1.n22 8.92171
R2773 VDD1.n54 VDD1.n53 8.92171
R2774 VDD1.n161 VDD1.n160 8.92171
R2775 VDD1.n176 VDD1.n129 8.92171
R2776 VDD1.n207 VDD1.n113 8.92171
R2777 VDD1.n102 VDD1.n101 8.14595
R2778 VDD1.n66 VDD1.n65 8.14595
R2779 VDD1.n57 VDD1.n28 8.14595
R2780 VDD1.n164 VDD1.n135 8.14595
R2781 VDD1.n173 VDD1.n172 8.14595
R2782 VDD1.n211 VDD1.n210 8.14595
R2783 VDD1.n108 VDD1.n0 7.3702
R2784 VDD1.n105 VDD1.n2 7.3702
R2785 VDD1.n62 VDD1.n24 7.3702
R2786 VDD1.n58 VDD1.n26 7.3702
R2787 VDD1.n165 VDD1.n133 7.3702
R2788 VDD1.n169 VDD1.n131 7.3702
R2789 VDD1.n214 VDD1.n111 7.3702
R2790 VDD1.n217 VDD1.n109 7.3702
R2791 VDD1.n106 VDD1.n0 6.59444
R2792 VDD1.n106 VDD1.n105 6.59444
R2793 VDD1.n62 VDD1.n61 6.59444
R2794 VDD1.n61 VDD1.n26 6.59444
R2795 VDD1.n168 VDD1.n133 6.59444
R2796 VDD1.n169 VDD1.n168 6.59444
R2797 VDD1.n215 VDD1.n214 6.59444
R2798 VDD1.n215 VDD1.n109 6.59444
R2799 VDD1.n102 VDD1.n2 5.81868
R2800 VDD1.n65 VDD1.n24 5.81868
R2801 VDD1.n58 VDD1.n57 5.81868
R2802 VDD1.n165 VDD1.n164 5.81868
R2803 VDD1.n172 VDD1.n131 5.81868
R2804 VDD1.n211 VDD1.n111 5.81868
R2805 VDD1.n101 VDD1.n4 5.04292
R2806 VDD1.n66 VDD1.n22 5.04292
R2807 VDD1.n54 VDD1.n28 5.04292
R2808 VDD1.n161 VDD1.n135 5.04292
R2809 VDD1.n173 VDD1.n129 5.04292
R2810 VDD1.n210 VDD1.n113 5.04292
R2811 VDD1.n37 VDD1.n35 4.38563
R2812 VDD1.n144 VDD1.n142 4.38563
R2813 VDD1.n98 VDD1.n97 4.26717
R2814 VDD1.n70 VDD1.n69 4.26717
R2815 VDD1.n53 VDD1.n30 4.26717
R2816 VDD1.n160 VDD1.n137 4.26717
R2817 VDD1.n177 VDD1.n176 4.26717
R2818 VDD1.n207 VDD1.n206 4.26717
R2819 VDD1.n94 VDD1.n6 3.49141
R2820 VDD1.n73 VDD1.n20 3.49141
R2821 VDD1.n50 VDD1.n49 3.49141
R2822 VDD1.n157 VDD1.n156 3.49141
R2823 VDD1.n180 VDD1.n127 3.49141
R2824 VDD1.n203 VDD1.n115 3.49141
R2825 VDD1.n93 VDD1.n8 2.71565
R2826 VDD1.n74 VDD1.n18 2.71565
R2827 VDD1.n46 VDD1.n32 2.71565
R2828 VDD1.n153 VDD1.n139 2.71565
R2829 VDD1.n181 VDD1.n125 2.71565
R2830 VDD1.n202 VDD1.n117 2.71565
R2831 VDD1.n90 VDD1.n89 1.93989
R2832 VDD1.n78 VDD1.n77 1.93989
R2833 VDD1.n45 VDD1.n34 1.93989
R2834 VDD1.n152 VDD1.n141 1.93989
R2835 VDD1.n186 VDD1.n184 1.93989
R2836 VDD1.n199 VDD1.n198 1.93989
R2837 VDD1.n86 VDD1.n10 1.16414
R2838 VDD1.n81 VDD1.n15 1.16414
R2839 VDD1.n42 VDD1.n41 1.16414
R2840 VDD1.n149 VDD1.n148 1.16414
R2841 VDD1.n185 VDD1.n123 1.16414
R2842 VDD1.n195 VDD1.n119 1.16414
R2843 VDD1.n220 VDD1.t1 1.00813
R2844 VDD1.n220 VDD1.t0 1.00813
R2845 VDD1.n218 VDD1.t3 1.00813
R2846 VDD1.n218 VDD1.t5 1.00813
R2847 VDD1.n85 VDD1.n12 0.388379
R2848 VDD1.n82 VDD1.n14 0.388379
R2849 VDD1.n38 VDD1.n36 0.388379
R2850 VDD1.n145 VDD1.n143 0.388379
R2851 VDD1.n191 VDD1.n190 0.388379
R2852 VDD1.n194 VDD1.n121 0.388379
R2853 VDD1.n107 VDD1.n1 0.155672
R2854 VDD1.n100 VDD1.n1 0.155672
R2855 VDD1.n100 VDD1.n99 0.155672
R2856 VDD1.n99 VDD1.n5 0.155672
R2857 VDD1.n92 VDD1.n5 0.155672
R2858 VDD1.n92 VDD1.n91 0.155672
R2859 VDD1.n91 VDD1.n9 0.155672
R2860 VDD1.n84 VDD1.n9 0.155672
R2861 VDD1.n84 VDD1.n83 0.155672
R2862 VDD1.n83 VDD1.n13 0.155672
R2863 VDD1.n76 VDD1.n13 0.155672
R2864 VDD1.n76 VDD1.n75 0.155672
R2865 VDD1.n75 VDD1.n19 0.155672
R2866 VDD1.n68 VDD1.n19 0.155672
R2867 VDD1.n68 VDD1.n67 0.155672
R2868 VDD1.n67 VDD1.n23 0.155672
R2869 VDD1.n60 VDD1.n23 0.155672
R2870 VDD1.n60 VDD1.n59 0.155672
R2871 VDD1.n59 VDD1.n27 0.155672
R2872 VDD1.n52 VDD1.n27 0.155672
R2873 VDD1.n52 VDD1.n51 0.155672
R2874 VDD1.n51 VDD1.n31 0.155672
R2875 VDD1.n44 VDD1.n31 0.155672
R2876 VDD1.n44 VDD1.n43 0.155672
R2877 VDD1.n43 VDD1.n35 0.155672
R2878 VDD1.n150 VDD1.n142 0.155672
R2879 VDD1.n151 VDD1.n150 0.155672
R2880 VDD1.n151 VDD1.n138 0.155672
R2881 VDD1.n158 VDD1.n138 0.155672
R2882 VDD1.n159 VDD1.n158 0.155672
R2883 VDD1.n159 VDD1.n134 0.155672
R2884 VDD1.n166 VDD1.n134 0.155672
R2885 VDD1.n167 VDD1.n166 0.155672
R2886 VDD1.n167 VDD1.n130 0.155672
R2887 VDD1.n174 VDD1.n130 0.155672
R2888 VDD1.n175 VDD1.n174 0.155672
R2889 VDD1.n175 VDD1.n126 0.155672
R2890 VDD1.n182 VDD1.n126 0.155672
R2891 VDD1.n183 VDD1.n182 0.155672
R2892 VDD1.n183 VDD1.n122 0.155672
R2893 VDD1.n192 VDD1.n122 0.155672
R2894 VDD1.n193 VDD1.n192 0.155672
R2895 VDD1.n193 VDD1.n118 0.155672
R2896 VDD1.n200 VDD1.n118 0.155672
R2897 VDD1.n201 VDD1.n200 0.155672
R2898 VDD1.n201 VDD1.n114 0.155672
R2899 VDD1.n208 VDD1.n114 0.155672
R2900 VDD1.n209 VDD1.n208 0.155672
R2901 VDD1.n209 VDD1.n110 0.155672
R2902 VDD1.n216 VDD1.n110 0.155672
R2903 VDD1 VDD1.n221 0.155672
C0 VN VDD2 6.69264f
C1 VTAIL VDD2 15.482201f
C2 VP VDD2 0.295202f
C3 VDD1 VDD2 0.696995f
C4 VN VTAIL 6.05736f
C5 VP VN 6.46173f
C6 VN VDD1 0.147852f
C7 VP VTAIL 6.07231f
C8 VTAIL VDD1 15.4529f
C9 VP VDD1 6.83272f
C10 VDD2 B 5.833871f
C11 VDD1 B 5.843071f
C12 VTAIL B 9.138285f
C13 VN B 8.59822f
C14 VP B 6.167877f
C15 VDD1.n0 B 0.033997f
C16 VDD1.n1 B 0.02362f
C17 VDD1.n2 B 0.012692f
C18 VDD1.n3 B 0.03f
C19 VDD1.n4 B 0.013439f
C20 VDD1.n5 B 0.02362f
C21 VDD1.n6 B 0.012692f
C22 VDD1.n7 B 0.03f
C23 VDD1.n8 B 0.013439f
C24 VDD1.n9 B 0.02362f
C25 VDD1.n10 B 0.012692f
C26 VDD1.n11 B 0.03f
C27 VDD1.n12 B 0.013066f
C28 VDD1.n13 B 0.02362f
C29 VDD1.n14 B 0.013066f
C30 VDD1.n15 B 0.012692f
C31 VDD1.n16 B 0.03f
C32 VDD1.n17 B 0.03f
C33 VDD1.n18 B 0.013439f
C34 VDD1.n19 B 0.02362f
C35 VDD1.n20 B 0.012692f
C36 VDD1.n21 B 0.03f
C37 VDD1.n22 B 0.013439f
C38 VDD1.n23 B 0.02362f
C39 VDD1.n24 B 0.012692f
C40 VDD1.n25 B 0.03f
C41 VDD1.n26 B 0.013439f
C42 VDD1.n27 B 0.02362f
C43 VDD1.n28 B 0.012692f
C44 VDD1.n29 B 0.03f
C45 VDD1.n30 B 0.013439f
C46 VDD1.n31 B 0.02362f
C47 VDD1.n32 B 0.012692f
C48 VDD1.n33 B 0.03f
C49 VDD1.n34 B 0.013439f
C50 VDD1.n35 B 2.04013f
C51 VDD1.n36 B 0.012692f
C52 VDD1.t2 B 0.049844f
C53 VDD1.n37 B 0.181594f
C54 VDD1.n38 B 0.017722f
C55 VDD1.n39 B 0.0225f
C56 VDD1.n40 B 0.03f
C57 VDD1.n41 B 0.013439f
C58 VDD1.n42 B 0.012692f
C59 VDD1.n43 B 0.02362f
C60 VDD1.n44 B 0.02362f
C61 VDD1.n45 B 0.012692f
C62 VDD1.n46 B 0.013439f
C63 VDD1.n47 B 0.03f
C64 VDD1.n48 B 0.03f
C65 VDD1.n49 B 0.013439f
C66 VDD1.n50 B 0.012692f
C67 VDD1.n51 B 0.02362f
C68 VDD1.n52 B 0.02362f
C69 VDD1.n53 B 0.012692f
C70 VDD1.n54 B 0.013439f
C71 VDD1.n55 B 0.03f
C72 VDD1.n56 B 0.03f
C73 VDD1.n57 B 0.013439f
C74 VDD1.n58 B 0.012692f
C75 VDD1.n59 B 0.02362f
C76 VDD1.n60 B 0.02362f
C77 VDD1.n61 B 0.012692f
C78 VDD1.n62 B 0.013439f
C79 VDD1.n63 B 0.03f
C80 VDD1.n64 B 0.03f
C81 VDD1.n65 B 0.013439f
C82 VDD1.n66 B 0.012692f
C83 VDD1.n67 B 0.02362f
C84 VDD1.n68 B 0.02362f
C85 VDD1.n69 B 0.012692f
C86 VDD1.n70 B 0.013439f
C87 VDD1.n71 B 0.03f
C88 VDD1.n72 B 0.03f
C89 VDD1.n73 B 0.013439f
C90 VDD1.n74 B 0.012692f
C91 VDD1.n75 B 0.02362f
C92 VDD1.n76 B 0.02362f
C93 VDD1.n77 B 0.012692f
C94 VDD1.n78 B 0.013439f
C95 VDD1.n79 B 0.03f
C96 VDD1.n80 B 0.03f
C97 VDD1.n81 B 0.013439f
C98 VDD1.n82 B 0.012692f
C99 VDD1.n83 B 0.02362f
C100 VDD1.n84 B 0.02362f
C101 VDD1.n85 B 0.012692f
C102 VDD1.n86 B 0.013439f
C103 VDD1.n87 B 0.03f
C104 VDD1.n88 B 0.03f
C105 VDD1.n89 B 0.013439f
C106 VDD1.n90 B 0.012692f
C107 VDD1.n91 B 0.02362f
C108 VDD1.n92 B 0.02362f
C109 VDD1.n93 B 0.012692f
C110 VDD1.n94 B 0.013439f
C111 VDD1.n95 B 0.03f
C112 VDD1.n96 B 0.03f
C113 VDD1.n97 B 0.013439f
C114 VDD1.n98 B 0.012692f
C115 VDD1.n99 B 0.02362f
C116 VDD1.n100 B 0.02362f
C117 VDD1.n101 B 0.012692f
C118 VDD1.n102 B 0.013439f
C119 VDD1.n103 B 0.03f
C120 VDD1.n104 B 0.066355f
C121 VDD1.n105 B 0.013439f
C122 VDD1.n106 B 0.012692f
C123 VDD1.n107 B 0.053629f
C124 VDD1.n108 B 0.054958f
C125 VDD1.n109 B 0.033997f
C126 VDD1.n110 B 0.02362f
C127 VDD1.n111 B 0.012692f
C128 VDD1.n112 B 0.03f
C129 VDD1.n113 B 0.013439f
C130 VDD1.n114 B 0.02362f
C131 VDD1.n115 B 0.012692f
C132 VDD1.n116 B 0.03f
C133 VDD1.n117 B 0.013439f
C134 VDD1.n118 B 0.02362f
C135 VDD1.n119 B 0.012692f
C136 VDD1.n120 B 0.03f
C137 VDD1.n121 B 0.013066f
C138 VDD1.n122 B 0.02362f
C139 VDD1.n123 B 0.013439f
C140 VDD1.n124 B 0.03f
C141 VDD1.n125 B 0.013439f
C142 VDD1.n126 B 0.02362f
C143 VDD1.n127 B 0.012692f
C144 VDD1.n128 B 0.03f
C145 VDD1.n129 B 0.013439f
C146 VDD1.n130 B 0.02362f
C147 VDD1.n131 B 0.012692f
C148 VDD1.n132 B 0.03f
C149 VDD1.n133 B 0.013439f
C150 VDD1.n134 B 0.02362f
C151 VDD1.n135 B 0.012692f
C152 VDD1.n136 B 0.03f
C153 VDD1.n137 B 0.013439f
C154 VDD1.n138 B 0.02362f
C155 VDD1.n139 B 0.012692f
C156 VDD1.n140 B 0.03f
C157 VDD1.n141 B 0.013439f
C158 VDD1.n142 B 2.04013f
C159 VDD1.n143 B 0.012692f
C160 VDD1.t4 B 0.049844f
C161 VDD1.n144 B 0.181594f
C162 VDD1.n145 B 0.017722f
C163 VDD1.n146 B 0.0225f
C164 VDD1.n147 B 0.03f
C165 VDD1.n148 B 0.013439f
C166 VDD1.n149 B 0.012692f
C167 VDD1.n150 B 0.02362f
C168 VDD1.n151 B 0.02362f
C169 VDD1.n152 B 0.012692f
C170 VDD1.n153 B 0.013439f
C171 VDD1.n154 B 0.03f
C172 VDD1.n155 B 0.03f
C173 VDD1.n156 B 0.013439f
C174 VDD1.n157 B 0.012692f
C175 VDD1.n158 B 0.02362f
C176 VDD1.n159 B 0.02362f
C177 VDD1.n160 B 0.012692f
C178 VDD1.n161 B 0.013439f
C179 VDD1.n162 B 0.03f
C180 VDD1.n163 B 0.03f
C181 VDD1.n164 B 0.013439f
C182 VDD1.n165 B 0.012692f
C183 VDD1.n166 B 0.02362f
C184 VDD1.n167 B 0.02362f
C185 VDD1.n168 B 0.012692f
C186 VDD1.n169 B 0.013439f
C187 VDD1.n170 B 0.03f
C188 VDD1.n171 B 0.03f
C189 VDD1.n172 B 0.013439f
C190 VDD1.n173 B 0.012692f
C191 VDD1.n174 B 0.02362f
C192 VDD1.n175 B 0.02362f
C193 VDD1.n176 B 0.012692f
C194 VDD1.n177 B 0.013439f
C195 VDD1.n178 B 0.03f
C196 VDD1.n179 B 0.03f
C197 VDD1.n180 B 0.013439f
C198 VDD1.n181 B 0.012692f
C199 VDD1.n182 B 0.02362f
C200 VDD1.n183 B 0.02362f
C201 VDD1.n184 B 0.012692f
C202 VDD1.n185 B 0.012692f
C203 VDD1.n186 B 0.013439f
C204 VDD1.n187 B 0.03f
C205 VDD1.n188 B 0.03f
C206 VDD1.n189 B 0.03f
C207 VDD1.n190 B 0.013066f
C208 VDD1.n191 B 0.012692f
C209 VDD1.n192 B 0.02362f
C210 VDD1.n193 B 0.02362f
C211 VDD1.n194 B 0.012692f
C212 VDD1.n195 B 0.013439f
C213 VDD1.n196 B 0.03f
C214 VDD1.n197 B 0.03f
C215 VDD1.n198 B 0.013439f
C216 VDD1.n199 B 0.012692f
C217 VDD1.n200 B 0.02362f
C218 VDD1.n201 B 0.02362f
C219 VDD1.n202 B 0.012692f
C220 VDD1.n203 B 0.013439f
C221 VDD1.n204 B 0.03f
C222 VDD1.n205 B 0.03f
C223 VDD1.n206 B 0.013439f
C224 VDD1.n207 B 0.012692f
C225 VDD1.n208 B 0.02362f
C226 VDD1.n209 B 0.02362f
C227 VDD1.n210 B 0.012692f
C228 VDD1.n211 B 0.013439f
C229 VDD1.n212 B 0.03f
C230 VDD1.n213 B 0.066355f
C231 VDD1.n214 B 0.013439f
C232 VDD1.n215 B 0.012692f
C233 VDD1.n216 B 0.053629f
C234 VDD1.n217 B 0.054641f
C235 VDD1.t3 B 0.366774f
C236 VDD1.t5 B 0.366774f
C237 VDD1.n218 B 3.352f
C238 VDD1.n219 B 2.25959f
C239 VDD1.t1 B 0.366774f
C240 VDD1.t0 B 0.366774f
C241 VDD1.n220 B 3.35124f
C242 VDD1.n221 B 2.67617f
C243 VP.n0 B 0.047236f
C244 VP.n1 B 0.010719f
C245 VP.n2 B 0.192098f
C246 VP.t5 B 1.73543f
C247 VP.t4 B 1.73543f
C248 VP.t3 B 1.75233f
C249 VP.n3 B 0.636486f
C250 VP.n4 B 0.653523f
C251 VP.n5 B 0.010719f
C252 VP.n6 B 0.645013f
C253 VP.n7 B 2.32084f
C254 VP.t1 B 1.73543f
C255 VP.n8 B 0.645013f
C256 VP.n9 B 2.35712f
C257 VP.n10 B 0.047236f
C258 VP.n11 B 0.047236f
C259 VP.t2 B 1.73543f
C260 VP.n12 B 0.650255f
C261 VP.n13 B 0.010719f
C262 VP.t0 B 1.73543f
C263 VP.n14 B 0.645013f
C264 VP.n15 B 0.036606f
C265 VDD2.n0 B 0.033978f
C266 VDD2.n1 B 0.023607f
C267 VDD2.n2 B 0.012685f
C268 VDD2.n3 B 0.029983f
C269 VDD2.n4 B 0.013431f
C270 VDD2.n5 B 0.023607f
C271 VDD2.n6 B 0.012685f
C272 VDD2.n7 B 0.029983f
C273 VDD2.n8 B 0.013431f
C274 VDD2.n9 B 0.023607f
C275 VDD2.n10 B 0.012685f
C276 VDD2.n11 B 0.029983f
C277 VDD2.n12 B 0.013058f
C278 VDD2.n13 B 0.023607f
C279 VDD2.n14 B 0.013431f
C280 VDD2.n15 B 0.029983f
C281 VDD2.n16 B 0.013431f
C282 VDD2.n17 B 0.023607f
C283 VDD2.n18 B 0.012685f
C284 VDD2.n19 B 0.029983f
C285 VDD2.n20 B 0.013431f
C286 VDD2.n21 B 0.023607f
C287 VDD2.n22 B 0.012685f
C288 VDD2.n23 B 0.029983f
C289 VDD2.n24 B 0.013431f
C290 VDD2.n25 B 0.023607f
C291 VDD2.n26 B 0.012685f
C292 VDD2.n27 B 0.029983f
C293 VDD2.n28 B 0.013431f
C294 VDD2.n29 B 0.023607f
C295 VDD2.n30 B 0.012685f
C296 VDD2.n31 B 0.029983f
C297 VDD2.n32 B 0.013431f
C298 VDD2.n33 B 2.03896f
C299 VDD2.n34 B 0.012685f
C300 VDD2.t5 B 0.049815f
C301 VDD2.n35 B 0.181489f
C302 VDD2.n36 B 0.017712f
C303 VDD2.n37 B 0.022487f
C304 VDD2.n38 B 0.029983f
C305 VDD2.n39 B 0.013431f
C306 VDD2.n40 B 0.012685f
C307 VDD2.n41 B 0.023607f
C308 VDD2.n42 B 0.023607f
C309 VDD2.n43 B 0.012685f
C310 VDD2.n44 B 0.013431f
C311 VDD2.n45 B 0.029983f
C312 VDD2.n46 B 0.029983f
C313 VDD2.n47 B 0.013431f
C314 VDD2.n48 B 0.012685f
C315 VDD2.n49 B 0.023607f
C316 VDD2.n50 B 0.023607f
C317 VDD2.n51 B 0.012685f
C318 VDD2.n52 B 0.013431f
C319 VDD2.n53 B 0.029983f
C320 VDD2.n54 B 0.029983f
C321 VDD2.n55 B 0.013431f
C322 VDD2.n56 B 0.012685f
C323 VDD2.n57 B 0.023607f
C324 VDD2.n58 B 0.023607f
C325 VDD2.n59 B 0.012685f
C326 VDD2.n60 B 0.013431f
C327 VDD2.n61 B 0.029983f
C328 VDD2.n62 B 0.029983f
C329 VDD2.n63 B 0.013431f
C330 VDD2.n64 B 0.012685f
C331 VDD2.n65 B 0.023607f
C332 VDD2.n66 B 0.023607f
C333 VDD2.n67 B 0.012685f
C334 VDD2.n68 B 0.013431f
C335 VDD2.n69 B 0.029983f
C336 VDD2.n70 B 0.029983f
C337 VDD2.n71 B 0.013431f
C338 VDD2.n72 B 0.012685f
C339 VDD2.n73 B 0.023607f
C340 VDD2.n74 B 0.023607f
C341 VDD2.n75 B 0.012685f
C342 VDD2.n76 B 0.012685f
C343 VDD2.n77 B 0.013431f
C344 VDD2.n78 B 0.029983f
C345 VDD2.n79 B 0.029983f
C346 VDD2.n80 B 0.029983f
C347 VDD2.n81 B 0.013058f
C348 VDD2.n82 B 0.012685f
C349 VDD2.n83 B 0.023607f
C350 VDD2.n84 B 0.023607f
C351 VDD2.n85 B 0.012685f
C352 VDD2.n86 B 0.013431f
C353 VDD2.n87 B 0.029983f
C354 VDD2.n88 B 0.029983f
C355 VDD2.n89 B 0.013431f
C356 VDD2.n90 B 0.012685f
C357 VDD2.n91 B 0.023607f
C358 VDD2.n92 B 0.023607f
C359 VDD2.n93 B 0.012685f
C360 VDD2.n94 B 0.013431f
C361 VDD2.n95 B 0.029983f
C362 VDD2.n96 B 0.029983f
C363 VDD2.n97 B 0.013431f
C364 VDD2.n98 B 0.012685f
C365 VDD2.n99 B 0.023607f
C366 VDD2.n100 B 0.023607f
C367 VDD2.n101 B 0.012685f
C368 VDD2.n102 B 0.013431f
C369 VDD2.n103 B 0.029983f
C370 VDD2.n104 B 0.066317f
C371 VDD2.n105 B 0.013431f
C372 VDD2.n106 B 0.012685f
C373 VDD2.n107 B 0.053598f
C374 VDD2.n108 B 0.05461f
C375 VDD2.t3 B 0.366564f
C376 VDD2.t4 B 0.366564f
C377 VDD2.n109 B 3.35008f
C378 VDD2.n110 B 2.18464f
C379 VDD2.n111 B 0.033978f
C380 VDD2.n112 B 0.023607f
C381 VDD2.n113 B 0.012685f
C382 VDD2.n114 B 0.029983f
C383 VDD2.n115 B 0.013431f
C384 VDD2.n116 B 0.023607f
C385 VDD2.n117 B 0.012685f
C386 VDD2.n118 B 0.029983f
C387 VDD2.n119 B 0.013431f
C388 VDD2.n120 B 0.023607f
C389 VDD2.n121 B 0.012685f
C390 VDD2.n122 B 0.029983f
C391 VDD2.n123 B 0.013058f
C392 VDD2.n124 B 0.023607f
C393 VDD2.n125 B 0.013058f
C394 VDD2.n126 B 0.012685f
C395 VDD2.n127 B 0.029983f
C396 VDD2.n128 B 0.029983f
C397 VDD2.n129 B 0.013431f
C398 VDD2.n130 B 0.023607f
C399 VDD2.n131 B 0.012685f
C400 VDD2.n132 B 0.029983f
C401 VDD2.n133 B 0.013431f
C402 VDD2.n134 B 0.023607f
C403 VDD2.n135 B 0.012685f
C404 VDD2.n136 B 0.029983f
C405 VDD2.n137 B 0.013431f
C406 VDD2.n138 B 0.023607f
C407 VDD2.n139 B 0.012685f
C408 VDD2.n140 B 0.029983f
C409 VDD2.n141 B 0.013431f
C410 VDD2.n142 B 0.023607f
C411 VDD2.n143 B 0.012685f
C412 VDD2.n144 B 0.029983f
C413 VDD2.n145 B 0.013431f
C414 VDD2.n146 B 2.03896f
C415 VDD2.n147 B 0.012685f
C416 VDD2.t0 B 0.049815f
C417 VDD2.n148 B 0.181489f
C418 VDD2.n149 B 0.017712f
C419 VDD2.n150 B 0.022487f
C420 VDD2.n151 B 0.029983f
C421 VDD2.n152 B 0.013431f
C422 VDD2.n153 B 0.012685f
C423 VDD2.n154 B 0.023607f
C424 VDD2.n155 B 0.023607f
C425 VDD2.n156 B 0.012685f
C426 VDD2.n157 B 0.013431f
C427 VDD2.n158 B 0.029983f
C428 VDD2.n159 B 0.029983f
C429 VDD2.n160 B 0.013431f
C430 VDD2.n161 B 0.012685f
C431 VDD2.n162 B 0.023607f
C432 VDD2.n163 B 0.023607f
C433 VDD2.n164 B 0.012685f
C434 VDD2.n165 B 0.013431f
C435 VDD2.n166 B 0.029983f
C436 VDD2.n167 B 0.029983f
C437 VDD2.n168 B 0.013431f
C438 VDD2.n169 B 0.012685f
C439 VDD2.n170 B 0.023607f
C440 VDD2.n171 B 0.023607f
C441 VDD2.n172 B 0.012685f
C442 VDD2.n173 B 0.013431f
C443 VDD2.n174 B 0.029983f
C444 VDD2.n175 B 0.029983f
C445 VDD2.n176 B 0.013431f
C446 VDD2.n177 B 0.012685f
C447 VDD2.n178 B 0.023607f
C448 VDD2.n179 B 0.023607f
C449 VDD2.n180 B 0.012685f
C450 VDD2.n181 B 0.013431f
C451 VDD2.n182 B 0.029983f
C452 VDD2.n183 B 0.029983f
C453 VDD2.n184 B 0.013431f
C454 VDD2.n185 B 0.012685f
C455 VDD2.n186 B 0.023607f
C456 VDD2.n187 B 0.023607f
C457 VDD2.n188 B 0.012685f
C458 VDD2.n189 B 0.013431f
C459 VDD2.n190 B 0.029983f
C460 VDD2.n191 B 0.029983f
C461 VDD2.n192 B 0.013431f
C462 VDD2.n193 B 0.012685f
C463 VDD2.n194 B 0.023607f
C464 VDD2.n195 B 0.023607f
C465 VDD2.n196 B 0.012685f
C466 VDD2.n197 B 0.013431f
C467 VDD2.n198 B 0.029983f
C468 VDD2.n199 B 0.029983f
C469 VDD2.n200 B 0.013431f
C470 VDD2.n201 B 0.012685f
C471 VDD2.n202 B 0.023607f
C472 VDD2.n203 B 0.023607f
C473 VDD2.n204 B 0.012685f
C474 VDD2.n205 B 0.013431f
C475 VDD2.n206 B 0.029983f
C476 VDD2.n207 B 0.029983f
C477 VDD2.n208 B 0.013431f
C478 VDD2.n209 B 0.012685f
C479 VDD2.n210 B 0.023607f
C480 VDD2.n211 B 0.023607f
C481 VDD2.n212 B 0.012685f
C482 VDD2.n213 B 0.013431f
C483 VDD2.n214 B 0.029983f
C484 VDD2.n215 B 0.066317f
C485 VDD2.n216 B 0.013431f
C486 VDD2.n217 B 0.012685f
C487 VDD2.n218 B 0.053598f
C488 VDD2.n219 B 0.053529f
C489 VDD2.n220 B 2.47423f
C490 VDD2.t1 B 0.366564f
C491 VDD2.t2 B 0.366564f
C492 VDD2.n221 B 3.35005f
C493 VTAIL.t4 B 0.371056f
C494 VTAIL.t3 B 0.371056f
C495 VTAIL.n0 B 3.31473f
C496 VTAIL.n1 B 0.334191f
C497 VTAIL.n2 B 0.034394f
C498 VTAIL.n3 B 0.023896f
C499 VTAIL.n4 B 0.012841f
C500 VTAIL.n5 B 0.030351f
C501 VTAIL.n6 B 0.013596f
C502 VTAIL.n7 B 0.023896f
C503 VTAIL.n8 B 0.012841f
C504 VTAIL.n9 B 0.030351f
C505 VTAIL.n10 B 0.013596f
C506 VTAIL.n11 B 0.023896f
C507 VTAIL.n12 B 0.012841f
C508 VTAIL.n13 B 0.030351f
C509 VTAIL.n14 B 0.013218f
C510 VTAIL.n15 B 0.023896f
C511 VTAIL.n16 B 0.013596f
C512 VTAIL.n17 B 0.030351f
C513 VTAIL.n18 B 0.013596f
C514 VTAIL.n19 B 0.023896f
C515 VTAIL.n20 B 0.012841f
C516 VTAIL.n21 B 0.030351f
C517 VTAIL.n22 B 0.013596f
C518 VTAIL.n23 B 0.023896f
C519 VTAIL.n24 B 0.012841f
C520 VTAIL.n25 B 0.030351f
C521 VTAIL.n26 B 0.013596f
C522 VTAIL.n27 B 0.023896f
C523 VTAIL.n28 B 0.012841f
C524 VTAIL.n29 B 0.030351f
C525 VTAIL.n30 B 0.013596f
C526 VTAIL.n31 B 0.023896f
C527 VTAIL.n32 B 0.012841f
C528 VTAIL.n33 B 0.030351f
C529 VTAIL.n34 B 0.013596f
C530 VTAIL.n35 B 2.06395f
C531 VTAIL.n36 B 0.012841f
C532 VTAIL.t2 B 0.050426f
C533 VTAIL.n37 B 0.183714f
C534 VTAIL.n38 B 0.017929f
C535 VTAIL.n39 B 0.022763f
C536 VTAIL.n40 B 0.030351f
C537 VTAIL.n41 B 0.013596f
C538 VTAIL.n42 B 0.012841f
C539 VTAIL.n43 B 0.023896f
C540 VTAIL.n44 B 0.023896f
C541 VTAIL.n45 B 0.012841f
C542 VTAIL.n46 B 0.013596f
C543 VTAIL.n47 B 0.030351f
C544 VTAIL.n48 B 0.030351f
C545 VTAIL.n49 B 0.013596f
C546 VTAIL.n50 B 0.012841f
C547 VTAIL.n51 B 0.023896f
C548 VTAIL.n52 B 0.023896f
C549 VTAIL.n53 B 0.012841f
C550 VTAIL.n54 B 0.013596f
C551 VTAIL.n55 B 0.030351f
C552 VTAIL.n56 B 0.030351f
C553 VTAIL.n57 B 0.013596f
C554 VTAIL.n58 B 0.012841f
C555 VTAIL.n59 B 0.023896f
C556 VTAIL.n60 B 0.023896f
C557 VTAIL.n61 B 0.012841f
C558 VTAIL.n62 B 0.013596f
C559 VTAIL.n63 B 0.030351f
C560 VTAIL.n64 B 0.030351f
C561 VTAIL.n65 B 0.013596f
C562 VTAIL.n66 B 0.012841f
C563 VTAIL.n67 B 0.023896f
C564 VTAIL.n68 B 0.023896f
C565 VTAIL.n69 B 0.012841f
C566 VTAIL.n70 B 0.013596f
C567 VTAIL.n71 B 0.030351f
C568 VTAIL.n72 B 0.030351f
C569 VTAIL.n73 B 0.013596f
C570 VTAIL.n74 B 0.012841f
C571 VTAIL.n75 B 0.023896f
C572 VTAIL.n76 B 0.023896f
C573 VTAIL.n77 B 0.012841f
C574 VTAIL.n78 B 0.012841f
C575 VTAIL.n79 B 0.013596f
C576 VTAIL.n80 B 0.030351f
C577 VTAIL.n81 B 0.030351f
C578 VTAIL.n82 B 0.030351f
C579 VTAIL.n83 B 0.013218f
C580 VTAIL.n84 B 0.012841f
C581 VTAIL.n85 B 0.023896f
C582 VTAIL.n86 B 0.023896f
C583 VTAIL.n87 B 0.012841f
C584 VTAIL.n88 B 0.013596f
C585 VTAIL.n89 B 0.030351f
C586 VTAIL.n90 B 0.030351f
C587 VTAIL.n91 B 0.013596f
C588 VTAIL.n92 B 0.012841f
C589 VTAIL.n93 B 0.023896f
C590 VTAIL.n94 B 0.023896f
C591 VTAIL.n95 B 0.012841f
C592 VTAIL.n96 B 0.013596f
C593 VTAIL.n97 B 0.030351f
C594 VTAIL.n98 B 0.030351f
C595 VTAIL.n99 B 0.013596f
C596 VTAIL.n100 B 0.012841f
C597 VTAIL.n101 B 0.023896f
C598 VTAIL.n102 B 0.023896f
C599 VTAIL.n103 B 0.012841f
C600 VTAIL.n104 B 0.013596f
C601 VTAIL.n105 B 0.030351f
C602 VTAIL.n106 B 0.067129f
C603 VTAIL.n107 B 0.013596f
C604 VTAIL.n108 B 0.012841f
C605 VTAIL.n109 B 0.054255f
C606 VTAIL.n110 B 0.037678f
C607 VTAIL.n111 B 0.154603f
C608 VTAIL.t1 B 0.371056f
C609 VTAIL.t0 B 0.371056f
C610 VTAIL.n112 B 3.31473f
C611 VTAIL.n113 B 2.07031f
C612 VTAIL.t5 B 0.371056f
C613 VTAIL.t8 B 0.371056f
C614 VTAIL.n114 B 3.31475f
C615 VTAIL.n115 B 2.07029f
C616 VTAIL.n116 B 0.034394f
C617 VTAIL.n117 B 0.023896f
C618 VTAIL.n118 B 0.012841f
C619 VTAIL.n119 B 0.030351f
C620 VTAIL.n120 B 0.013596f
C621 VTAIL.n121 B 0.023896f
C622 VTAIL.n122 B 0.012841f
C623 VTAIL.n123 B 0.030351f
C624 VTAIL.n124 B 0.013596f
C625 VTAIL.n125 B 0.023896f
C626 VTAIL.n126 B 0.012841f
C627 VTAIL.n127 B 0.030351f
C628 VTAIL.n128 B 0.013218f
C629 VTAIL.n129 B 0.023896f
C630 VTAIL.n130 B 0.013218f
C631 VTAIL.n131 B 0.012841f
C632 VTAIL.n132 B 0.030351f
C633 VTAIL.n133 B 0.030351f
C634 VTAIL.n134 B 0.013596f
C635 VTAIL.n135 B 0.023896f
C636 VTAIL.n136 B 0.012841f
C637 VTAIL.n137 B 0.030351f
C638 VTAIL.n138 B 0.013596f
C639 VTAIL.n139 B 0.023896f
C640 VTAIL.n140 B 0.012841f
C641 VTAIL.n141 B 0.030351f
C642 VTAIL.n142 B 0.013596f
C643 VTAIL.n143 B 0.023896f
C644 VTAIL.n144 B 0.012841f
C645 VTAIL.n145 B 0.030351f
C646 VTAIL.n146 B 0.013596f
C647 VTAIL.n147 B 0.023896f
C648 VTAIL.n148 B 0.012841f
C649 VTAIL.n149 B 0.030351f
C650 VTAIL.n150 B 0.013596f
C651 VTAIL.n151 B 2.06395f
C652 VTAIL.n152 B 0.012841f
C653 VTAIL.t6 B 0.050426f
C654 VTAIL.n153 B 0.183714f
C655 VTAIL.n154 B 0.017929f
C656 VTAIL.n155 B 0.022763f
C657 VTAIL.n156 B 0.030351f
C658 VTAIL.n157 B 0.013596f
C659 VTAIL.n158 B 0.012841f
C660 VTAIL.n159 B 0.023896f
C661 VTAIL.n160 B 0.023896f
C662 VTAIL.n161 B 0.012841f
C663 VTAIL.n162 B 0.013596f
C664 VTAIL.n163 B 0.030351f
C665 VTAIL.n164 B 0.030351f
C666 VTAIL.n165 B 0.013596f
C667 VTAIL.n166 B 0.012841f
C668 VTAIL.n167 B 0.023896f
C669 VTAIL.n168 B 0.023896f
C670 VTAIL.n169 B 0.012841f
C671 VTAIL.n170 B 0.013596f
C672 VTAIL.n171 B 0.030351f
C673 VTAIL.n172 B 0.030351f
C674 VTAIL.n173 B 0.013596f
C675 VTAIL.n174 B 0.012841f
C676 VTAIL.n175 B 0.023896f
C677 VTAIL.n176 B 0.023896f
C678 VTAIL.n177 B 0.012841f
C679 VTAIL.n178 B 0.013596f
C680 VTAIL.n179 B 0.030351f
C681 VTAIL.n180 B 0.030351f
C682 VTAIL.n181 B 0.013596f
C683 VTAIL.n182 B 0.012841f
C684 VTAIL.n183 B 0.023896f
C685 VTAIL.n184 B 0.023896f
C686 VTAIL.n185 B 0.012841f
C687 VTAIL.n186 B 0.013596f
C688 VTAIL.n187 B 0.030351f
C689 VTAIL.n188 B 0.030351f
C690 VTAIL.n189 B 0.013596f
C691 VTAIL.n190 B 0.012841f
C692 VTAIL.n191 B 0.023896f
C693 VTAIL.n192 B 0.023896f
C694 VTAIL.n193 B 0.012841f
C695 VTAIL.n194 B 0.013596f
C696 VTAIL.n195 B 0.030351f
C697 VTAIL.n196 B 0.030351f
C698 VTAIL.n197 B 0.013596f
C699 VTAIL.n198 B 0.012841f
C700 VTAIL.n199 B 0.023896f
C701 VTAIL.n200 B 0.023896f
C702 VTAIL.n201 B 0.012841f
C703 VTAIL.n202 B 0.013596f
C704 VTAIL.n203 B 0.030351f
C705 VTAIL.n204 B 0.030351f
C706 VTAIL.n205 B 0.013596f
C707 VTAIL.n206 B 0.012841f
C708 VTAIL.n207 B 0.023896f
C709 VTAIL.n208 B 0.023896f
C710 VTAIL.n209 B 0.012841f
C711 VTAIL.n210 B 0.013596f
C712 VTAIL.n211 B 0.030351f
C713 VTAIL.n212 B 0.030351f
C714 VTAIL.n213 B 0.013596f
C715 VTAIL.n214 B 0.012841f
C716 VTAIL.n215 B 0.023896f
C717 VTAIL.n216 B 0.023896f
C718 VTAIL.n217 B 0.012841f
C719 VTAIL.n218 B 0.013596f
C720 VTAIL.n219 B 0.030351f
C721 VTAIL.n220 B 0.067129f
C722 VTAIL.n221 B 0.013596f
C723 VTAIL.n222 B 0.012841f
C724 VTAIL.n223 B 0.054255f
C725 VTAIL.n224 B 0.037678f
C726 VTAIL.n225 B 0.154603f
C727 VTAIL.t11 B 0.371056f
C728 VTAIL.t10 B 0.371056f
C729 VTAIL.n226 B 3.31475f
C730 VTAIL.n227 B 0.378982f
C731 VTAIL.n228 B 0.034394f
C732 VTAIL.n229 B 0.023896f
C733 VTAIL.n230 B 0.012841f
C734 VTAIL.n231 B 0.030351f
C735 VTAIL.n232 B 0.013596f
C736 VTAIL.n233 B 0.023896f
C737 VTAIL.n234 B 0.012841f
C738 VTAIL.n235 B 0.030351f
C739 VTAIL.n236 B 0.013596f
C740 VTAIL.n237 B 0.023896f
C741 VTAIL.n238 B 0.012841f
C742 VTAIL.n239 B 0.030351f
C743 VTAIL.n240 B 0.013218f
C744 VTAIL.n241 B 0.023896f
C745 VTAIL.n242 B 0.013218f
C746 VTAIL.n243 B 0.012841f
C747 VTAIL.n244 B 0.030351f
C748 VTAIL.n245 B 0.030351f
C749 VTAIL.n246 B 0.013596f
C750 VTAIL.n247 B 0.023896f
C751 VTAIL.n248 B 0.012841f
C752 VTAIL.n249 B 0.030351f
C753 VTAIL.n250 B 0.013596f
C754 VTAIL.n251 B 0.023896f
C755 VTAIL.n252 B 0.012841f
C756 VTAIL.n253 B 0.030351f
C757 VTAIL.n254 B 0.013596f
C758 VTAIL.n255 B 0.023896f
C759 VTAIL.n256 B 0.012841f
C760 VTAIL.n257 B 0.030351f
C761 VTAIL.n258 B 0.013596f
C762 VTAIL.n259 B 0.023896f
C763 VTAIL.n260 B 0.012841f
C764 VTAIL.n261 B 0.030351f
C765 VTAIL.n262 B 0.013596f
C766 VTAIL.n263 B 2.06395f
C767 VTAIL.n264 B 0.012841f
C768 VTAIL.t9 B 0.050426f
C769 VTAIL.n265 B 0.183714f
C770 VTAIL.n266 B 0.017929f
C771 VTAIL.n267 B 0.022763f
C772 VTAIL.n268 B 0.030351f
C773 VTAIL.n269 B 0.013596f
C774 VTAIL.n270 B 0.012841f
C775 VTAIL.n271 B 0.023896f
C776 VTAIL.n272 B 0.023896f
C777 VTAIL.n273 B 0.012841f
C778 VTAIL.n274 B 0.013596f
C779 VTAIL.n275 B 0.030351f
C780 VTAIL.n276 B 0.030351f
C781 VTAIL.n277 B 0.013596f
C782 VTAIL.n278 B 0.012841f
C783 VTAIL.n279 B 0.023896f
C784 VTAIL.n280 B 0.023896f
C785 VTAIL.n281 B 0.012841f
C786 VTAIL.n282 B 0.013596f
C787 VTAIL.n283 B 0.030351f
C788 VTAIL.n284 B 0.030351f
C789 VTAIL.n285 B 0.013596f
C790 VTAIL.n286 B 0.012841f
C791 VTAIL.n287 B 0.023896f
C792 VTAIL.n288 B 0.023896f
C793 VTAIL.n289 B 0.012841f
C794 VTAIL.n290 B 0.013596f
C795 VTAIL.n291 B 0.030351f
C796 VTAIL.n292 B 0.030351f
C797 VTAIL.n293 B 0.013596f
C798 VTAIL.n294 B 0.012841f
C799 VTAIL.n295 B 0.023896f
C800 VTAIL.n296 B 0.023896f
C801 VTAIL.n297 B 0.012841f
C802 VTAIL.n298 B 0.013596f
C803 VTAIL.n299 B 0.030351f
C804 VTAIL.n300 B 0.030351f
C805 VTAIL.n301 B 0.013596f
C806 VTAIL.n302 B 0.012841f
C807 VTAIL.n303 B 0.023896f
C808 VTAIL.n304 B 0.023896f
C809 VTAIL.n305 B 0.012841f
C810 VTAIL.n306 B 0.013596f
C811 VTAIL.n307 B 0.030351f
C812 VTAIL.n308 B 0.030351f
C813 VTAIL.n309 B 0.013596f
C814 VTAIL.n310 B 0.012841f
C815 VTAIL.n311 B 0.023896f
C816 VTAIL.n312 B 0.023896f
C817 VTAIL.n313 B 0.012841f
C818 VTAIL.n314 B 0.013596f
C819 VTAIL.n315 B 0.030351f
C820 VTAIL.n316 B 0.030351f
C821 VTAIL.n317 B 0.013596f
C822 VTAIL.n318 B 0.012841f
C823 VTAIL.n319 B 0.023896f
C824 VTAIL.n320 B 0.023896f
C825 VTAIL.n321 B 0.012841f
C826 VTAIL.n322 B 0.013596f
C827 VTAIL.n323 B 0.030351f
C828 VTAIL.n324 B 0.030351f
C829 VTAIL.n325 B 0.013596f
C830 VTAIL.n326 B 0.012841f
C831 VTAIL.n327 B 0.023896f
C832 VTAIL.n328 B 0.023896f
C833 VTAIL.n329 B 0.012841f
C834 VTAIL.n330 B 0.013596f
C835 VTAIL.n331 B 0.030351f
C836 VTAIL.n332 B 0.067129f
C837 VTAIL.n333 B 0.013596f
C838 VTAIL.n334 B 0.012841f
C839 VTAIL.n335 B 0.054255f
C840 VTAIL.n336 B 0.037678f
C841 VTAIL.n337 B 1.7802f
C842 VTAIL.n338 B 0.034394f
C843 VTAIL.n339 B 0.023896f
C844 VTAIL.n340 B 0.012841f
C845 VTAIL.n341 B 0.030351f
C846 VTAIL.n342 B 0.013596f
C847 VTAIL.n343 B 0.023896f
C848 VTAIL.n344 B 0.012841f
C849 VTAIL.n345 B 0.030351f
C850 VTAIL.n346 B 0.013596f
C851 VTAIL.n347 B 0.023896f
C852 VTAIL.n348 B 0.012841f
C853 VTAIL.n349 B 0.030351f
C854 VTAIL.n350 B 0.013218f
C855 VTAIL.n351 B 0.023896f
C856 VTAIL.n352 B 0.013596f
C857 VTAIL.n353 B 0.030351f
C858 VTAIL.n354 B 0.013596f
C859 VTAIL.n355 B 0.023896f
C860 VTAIL.n356 B 0.012841f
C861 VTAIL.n357 B 0.030351f
C862 VTAIL.n358 B 0.013596f
C863 VTAIL.n359 B 0.023896f
C864 VTAIL.n360 B 0.012841f
C865 VTAIL.n361 B 0.030351f
C866 VTAIL.n362 B 0.013596f
C867 VTAIL.n363 B 0.023896f
C868 VTAIL.n364 B 0.012841f
C869 VTAIL.n365 B 0.030351f
C870 VTAIL.n366 B 0.013596f
C871 VTAIL.n367 B 0.023896f
C872 VTAIL.n368 B 0.012841f
C873 VTAIL.n369 B 0.030351f
C874 VTAIL.n370 B 0.013596f
C875 VTAIL.n371 B 2.06395f
C876 VTAIL.n372 B 0.012841f
C877 VTAIL.t7 B 0.050426f
C878 VTAIL.n373 B 0.183714f
C879 VTAIL.n374 B 0.017929f
C880 VTAIL.n375 B 0.022763f
C881 VTAIL.n376 B 0.030351f
C882 VTAIL.n377 B 0.013596f
C883 VTAIL.n378 B 0.012841f
C884 VTAIL.n379 B 0.023896f
C885 VTAIL.n380 B 0.023896f
C886 VTAIL.n381 B 0.012841f
C887 VTAIL.n382 B 0.013596f
C888 VTAIL.n383 B 0.030351f
C889 VTAIL.n384 B 0.030351f
C890 VTAIL.n385 B 0.013596f
C891 VTAIL.n386 B 0.012841f
C892 VTAIL.n387 B 0.023896f
C893 VTAIL.n388 B 0.023896f
C894 VTAIL.n389 B 0.012841f
C895 VTAIL.n390 B 0.013596f
C896 VTAIL.n391 B 0.030351f
C897 VTAIL.n392 B 0.030351f
C898 VTAIL.n393 B 0.013596f
C899 VTAIL.n394 B 0.012841f
C900 VTAIL.n395 B 0.023896f
C901 VTAIL.n396 B 0.023896f
C902 VTAIL.n397 B 0.012841f
C903 VTAIL.n398 B 0.013596f
C904 VTAIL.n399 B 0.030351f
C905 VTAIL.n400 B 0.030351f
C906 VTAIL.n401 B 0.013596f
C907 VTAIL.n402 B 0.012841f
C908 VTAIL.n403 B 0.023896f
C909 VTAIL.n404 B 0.023896f
C910 VTAIL.n405 B 0.012841f
C911 VTAIL.n406 B 0.013596f
C912 VTAIL.n407 B 0.030351f
C913 VTAIL.n408 B 0.030351f
C914 VTAIL.n409 B 0.013596f
C915 VTAIL.n410 B 0.012841f
C916 VTAIL.n411 B 0.023896f
C917 VTAIL.n412 B 0.023896f
C918 VTAIL.n413 B 0.012841f
C919 VTAIL.n414 B 0.012841f
C920 VTAIL.n415 B 0.013596f
C921 VTAIL.n416 B 0.030351f
C922 VTAIL.n417 B 0.030351f
C923 VTAIL.n418 B 0.030351f
C924 VTAIL.n419 B 0.013218f
C925 VTAIL.n420 B 0.012841f
C926 VTAIL.n421 B 0.023896f
C927 VTAIL.n422 B 0.023896f
C928 VTAIL.n423 B 0.012841f
C929 VTAIL.n424 B 0.013596f
C930 VTAIL.n425 B 0.030351f
C931 VTAIL.n426 B 0.030351f
C932 VTAIL.n427 B 0.013596f
C933 VTAIL.n428 B 0.012841f
C934 VTAIL.n429 B 0.023896f
C935 VTAIL.n430 B 0.023896f
C936 VTAIL.n431 B 0.012841f
C937 VTAIL.n432 B 0.013596f
C938 VTAIL.n433 B 0.030351f
C939 VTAIL.n434 B 0.030351f
C940 VTAIL.n435 B 0.013596f
C941 VTAIL.n436 B 0.012841f
C942 VTAIL.n437 B 0.023896f
C943 VTAIL.n438 B 0.023896f
C944 VTAIL.n439 B 0.012841f
C945 VTAIL.n440 B 0.013596f
C946 VTAIL.n441 B 0.030351f
C947 VTAIL.n442 B 0.067129f
C948 VTAIL.n443 B 0.013596f
C949 VTAIL.n444 B 0.012841f
C950 VTAIL.n445 B 0.054255f
C951 VTAIL.n446 B 0.037678f
C952 VTAIL.n447 B 1.75929f
C953 VN.n0 B 0.190456f
C954 VN.t0 B 1.73735f
C955 VN.n1 B 0.631045f
C956 VN.t2 B 1.72059f
C957 VN.n2 B 0.647937f
C958 VN.n3 B 0.010627f
C959 VN.t1 B 1.72059f
C960 VN.n4 B 0.6395f
C961 VN.n5 B 0.036293f
C962 VN.n6 B 0.190456f
C963 VN.t3 B 1.73735f
C964 VN.n7 B 0.631045f
C965 VN.t4 B 1.72059f
C966 VN.n8 B 0.647937f
C967 VN.n9 B 0.010627f
C968 VN.t5 B 1.72059f
C969 VN.n10 B 0.6395f
C970 VN.n11 B 2.33155f
.ends

