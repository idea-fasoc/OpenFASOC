* NGSPICE file created from diff_pair_sample_0297.ext - technology: sky130A

.subckt diff_pair_sample_0297 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=3.3969 ps=18.2 w=8.71 l=2.31
X1 VDD1.t4 VP.t1 VTAIL.t7 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=1.43715 ps=9.04 w=8.71 l=2.31
X2 VDD2.t5 VN.t0 VTAIL.t4 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=1.43715 ps=9.04 w=8.71 l=2.31
X3 VDD2.t4 VN.t1 VTAIL.t3 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=3.3969 ps=18.2 w=8.71 l=2.31
X4 VDD2.t3 VN.t2 VTAIL.t11 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=1.43715 ps=9.04 w=8.71 l=2.31
X5 VDD2.t2 VN.t3 VTAIL.t2 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=3.3969 ps=18.2 w=8.71 l=2.31
X6 VTAIL.t10 VP.t2 VDD1.t3 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=1.43715 ps=9.04 w=8.71 l=2.31
X7 B.t11 B.t9 B.t10 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=0 ps=0 w=8.71 l=2.31
X8 VTAIL.t5 VP.t3 VDD1.t2 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=1.43715 ps=9.04 w=8.71 l=2.31
X9 B.t8 B.t6 B.t7 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=0 ps=0 w=8.71 l=2.31
X10 VTAIL.t1 VN.t4 VDD2.t1 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=1.43715 ps=9.04 w=8.71 l=2.31
X11 VTAIL.t0 VN.t5 VDD2.t0 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=1.43715 ps=9.04 w=8.71 l=2.31
X12 B.t5 B.t3 B.t4 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=0 ps=0 w=8.71 l=2.31
X13 B.t2 B.t0 B.t1 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=0 ps=0 w=8.71 l=2.31
X14 VDD1.t1 VP.t4 VTAIL.t6 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=1.43715 pd=9.04 as=3.3969 ps=18.2 w=8.71 l=2.31
X15 VDD1.t0 VP.t5 VTAIL.t9 w_n3082_n2710# sky130_fd_pr__pfet_01v8 ad=3.3969 pd=18.2 as=1.43715 ps=9.04 w=8.71 l=2.31
R0 VP.n11 VP.n8 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n7 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n6 161.3
R5 VP.n36 VP.n0 161.3
R6 VP.n35 VP.n34 161.3
R7 VP.n33 VP.n1 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n30 VP.n2 161.3
R10 VP.n28 VP.n27 161.3
R11 VP.n26 VP.n3 161.3
R12 VP.n25 VP.n24 161.3
R13 VP.n23 VP.n4 161.3
R14 VP.n22 VP.n21 161.3
R15 VP.n9 VP.t1 124.624
R16 VP.n20 VP.n5 91.6722
R17 VP.n38 VP.n37 91.6722
R18 VP.n19 VP.n18 91.6722
R19 VP.n5 VP.t5 90.8711
R20 VP.n29 VP.t2 90.8711
R21 VP.n37 VP.t0 90.8711
R22 VP.n18 VP.t4 90.8711
R23 VP.n10 VP.t3 90.8711
R24 VP.n10 VP.n9 59.2346
R25 VP.n24 VP.n23 47.2923
R26 VP.n35 VP.n1 47.2923
R27 VP.n16 VP.n7 47.2923
R28 VP.n20 VP.n19 45.1359
R29 VP.n24 VP.n3 33.6945
R30 VP.n31 VP.n1 33.6945
R31 VP.n12 VP.n7 33.6945
R32 VP.n23 VP.n22 24.4675
R33 VP.n28 VP.n3 24.4675
R34 VP.n31 VP.n30 24.4675
R35 VP.n36 VP.n35 24.4675
R36 VP.n17 VP.n16 24.4675
R37 VP.n12 VP.n11 24.4675
R38 VP.n22 VP.n5 19.0848
R39 VP.n37 VP.n36 19.0848
R40 VP.n18 VP.n17 19.0848
R41 VP.n29 VP.n28 12.234
R42 VP.n30 VP.n29 12.234
R43 VP.n11 VP.n10 12.234
R44 VP.n9 VP.n8 9.06133
R45 VP.n19 VP.n6 0.278367
R46 VP.n21 VP.n20 0.278367
R47 VP.n38 VP.n0 0.278367
R48 VP.n13 VP.n8 0.189894
R49 VP.n14 VP.n13 0.189894
R50 VP.n15 VP.n14 0.189894
R51 VP.n15 VP.n6 0.189894
R52 VP.n21 VP.n4 0.189894
R53 VP.n25 VP.n4 0.189894
R54 VP.n26 VP.n25 0.189894
R55 VP.n27 VP.n26 0.189894
R56 VP.n27 VP.n2 0.189894
R57 VP.n32 VP.n2 0.189894
R58 VP.n33 VP.n32 0.189894
R59 VP.n34 VP.n33 0.189894
R60 VP.n34 VP.n0 0.189894
R61 VP VP.n38 0.153454
R62 VTAIL.n186 VTAIL.n146 756.745
R63 VTAIL.n42 VTAIL.n2 756.745
R64 VTAIL.n140 VTAIL.n100 756.745
R65 VTAIL.n92 VTAIL.n52 756.745
R66 VTAIL.n161 VTAIL.n160 585
R67 VTAIL.n158 VTAIL.n157 585
R68 VTAIL.n167 VTAIL.n166 585
R69 VTAIL.n169 VTAIL.n168 585
R70 VTAIL.n154 VTAIL.n153 585
R71 VTAIL.n175 VTAIL.n174 585
R72 VTAIL.n178 VTAIL.n177 585
R73 VTAIL.n176 VTAIL.n150 585
R74 VTAIL.n183 VTAIL.n149 585
R75 VTAIL.n185 VTAIL.n184 585
R76 VTAIL.n187 VTAIL.n186 585
R77 VTAIL.n17 VTAIL.n16 585
R78 VTAIL.n14 VTAIL.n13 585
R79 VTAIL.n23 VTAIL.n22 585
R80 VTAIL.n25 VTAIL.n24 585
R81 VTAIL.n10 VTAIL.n9 585
R82 VTAIL.n31 VTAIL.n30 585
R83 VTAIL.n34 VTAIL.n33 585
R84 VTAIL.n32 VTAIL.n6 585
R85 VTAIL.n39 VTAIL.n5 585
R86 VTAIL.n41 VTAIL.n40 585
R87 VTAIL.n43 VTAIL.n42 585
R88 VTAIL.n141 VTAIL.n140 585
R89 VTAIL.n139 VTAIL.n138 585
R90 VTAIL.n137 VTAIL.n103 585
R91 VTAIL.n107 VTAIL.n104 585
R92 VTAIL.n132 VTAIL.n131 585
R93 VTAIL.n130 VTAIL.n129 585
R94 VTAIL.n109 VTAIL.n108 585
R95 VTAIL.n124 VTAIL.n123 585
R96 VTAIL.n122 VTAIL.n121 585
R97 VTAIL.n113 VTAIL.n112 585
R98 VTAIL.n116 VTAIL.n115 585
R99 VTAIL.n93 VTAIL.n92 585
R100 VTAIL.n91 VTAIL.n90 585
R101 VTAIL.n89 VTAIL.n55 585
R102 VTAIL.n59 VTAIL.n56 585
R103 VTAIL.n84 VTAIL.n83 585
R104 VTAIL.n82 VTAIL.n81 585
R105 VTAIL.n61 VTAIL.n60 585
R106 VTAIL.n76 VTAIL.n75 585
R107 VTAIL.n74 VTAIL.n73 585
R108 VTAIL.n65 VTAIL.n64 585
R109 VTAIL.n68 VTAIL.n67 585
R110 VTAIL.t6 VTAIL.n114 329.039
R111 VTAIL.t2 VTAIL.n66 329.039
R112 VTAIL.t3 VTAIL.n159 329.038
R113 VTAIL.t8 VTAIL.n15 329.038
R114 VTAIL.n160 VTAIL.n157 171.744
R115 VTAIL.n167 VTAIL.n157 171.744
R116 VTAIL.n168 VTAIL.n167 171.744
R117 VTAIL.n168 VTAIL.n153 171.744
R118 VTAIL.n175 VTAIL.n153 171.744
R119 VTAIL.n177 VTAIL.n175 171.744
R120 VTAIL.n177 VTAIL.n176 171.744
R121 VTAIL.n176 VTAIL.n149 171.744
R122 VTAIL.n185 VTAIL.n149 171.744
R123 VTAIL.n186 VTAIL.n185 171.744
R124 VTAIL.n16 VTAIL.n13 171.744
R125 VTAIL.n23 VTAIL.n13 171.744
R126 VTAIL.n24 VTAIL.n23 171.744
R127 VTAIL.n24 VTAIL.n9 171.744
R128 VTAIL.n31 VTAIL.n9 171.744
R129 VTAIL.n33 VTAIL.n31 171.744
R130 VTAIL.n33 VTAIL.n32 171.744
R131 VTAIL.n32 VTAIL.n5 171.744
R132 VTAIL.n41 VTAIL.n5 171.744
R133 VTAIL.n42 VTAIL.n41 171.744
R134 VTAIL.n140 VTAIL.n139 171.744
R135 VTAIL.n139 VTAIL.n103 171.744
R136 VTAIL.n107 VTAIL.n103 171.744
R137 VTAIL.n131 VTAIL.n107 171.744
R138 VTAIL.n131 VTAIL.n130 171.744
R139 VTAIL.n130 VTAIL.n108 171.744
R140 VTAIL.n123 VTAIL.n108 171.744
R141 VTAIL.n123 VTAIL.n122 171.744
R142 VTAIL.n122 VTAIL.n112 171.744
R143 VTAIL.n115 VTAIL.n112 171.744
R144 VTAIL.n92 VTAIL.n91 171.744
R145 VTAIL.n91 VTAIL.n55 171.744
R146 VTAIL.n59 VTAIL.n55 171.744
R147 VTAIL.n83 VTAIL.n59 171.744
R148 VTAIL.n83 VTAIL.n82 171.744
R149 VTAIL.n82 VTAIL.n60 171.744
R150 VTAIL.n75 VTAIL.n60 171.744
R151 VTAIL.n75 VTAIL.n74 171.744
R152 VTAIL.n74 VTAIL.n64 171.744
R153 VTAIL.n67 VTAIL.n64 171.744
R154 VTAIL.n160 VTAIL.t3 85.8723
R155 VTAIL.n16 VTAIL.t8 85.8723
R156 VTAIL.n115 VTAIL.t6 85.8723
R157 VTAIL.n67 VTAIL.t2 85.8723
R158 VTAIL.n99 VTAIL.n98 67.3103
R159 VTAIL.n51 VTAIL.n50 67.3103
R160 VTAIL.n1 VTAIL.n0 67.3102
R161 VTAIL.n49 VTAIL.n48 67.3102
R162 VTAIL.n191 VTAIL.n190 35.8702
R163 VTAIL.n47 VTAIL.n46 35.8702
R164 VTAIL.n145 VTAIL.n144 35.8702
R165 VTAIL.n97 VTAIL.n96 35.8702
R166 VTAIL.n51 VTAIL.n49 24.4272
R167 VTAIL.n191 VTAIL.n145 22.1514
R168 VTAIL.n184 VTAIL.n183 13.1884
R169 VTAIL.n40 VTAIL.n39 13.1884
R170 VTAIL.n138 VTAIL.n137 13.1884
R171 VTAIL.n90 VTAIL.n89 13.1884
R172 VTAIL.n182 VTAIL.n150 12.8005
R173 VTAIL.n187 VTAIL.n148 12.8005
R174 VTAIL.n38 VTAIL.n6 12.8005
R175 VTAIL.n43 VTAIL.n4 12.8005
R176 VTAIL.n141 VTAIL.n102 12.8005
R177 VTAIL.n136 VTAIL.n104 12.8005
R178 VTAIL.n93 VTAIL.n54 12.8005
R179 VTAIL.n88 VTAIL.n56 12.8005
R180 VTAIL.n179 VTAIL.n178 12.0247
R181 VTAIL.n188 VTAIL.n146 12.0247
R182 VTAIL.n35 VTAIL.n34 12.0247
R183 VTAIL.n44 VTAIL.n2 12.0247
R184 VTAIL.n142 VTAIL.n100 12.0247
R185 VTAIL.n133 VTAIL.n132 12.0247
R186 VTAIL.n94 VTAIL.n52 12.0247
R187 VTAIL.n85 VTAIL.n84 12.0247
R188 VTAIL.n174 VTAIL.n152 11.249
R189 VTAIL.n30 VTAIL.n8 11.249
R190 VTAIL.n129 VTAIL.n106 11.249
R191 VTAIL.n81 VTAIL.n58 11.249
R192 VTAIL.n161 VTAIL.n159 10.7239
R193 VTAIL.n17 VTAIL.n15 10.7239
R194 VTAIL.n116 VTAIL.n114 10.7239
R195 VTAIL.n68 VTAIL.n66 10.7239
R196 VTAIL.n173 VTAIL.n154 10.4732
R197 VTAIL.n29 VTAIL.n10 10.4732
R198 VTAIL.n128 VTAIL.n109 10.4732
R199 VTAIL.n80 VTAIL.n61 10.4732
R200 VTAIL.n170 VTAIL.n169 9.69747
R201 VTAIL.n26 VTAIL.n25 9.69747
R202 VTAIL.n125 VTAIL.n124 9.69747
R203 VTAIL.n77 VTAIL.n76 9.69747
R204 VTAIL.n190 VTAIL.n189 9.45567
R205 VTAIL.n46 VTAIL.n45 9.45567
R206 VTAIL.n144 VTAIL.n143 9.45567
R207 VTAIL.n96 VTAIL.n95 9.45567
R208 VTAIL.n189 VTAIL.n188 9.3005
R209 VTAIL.n148 VTAIL.n147 9.3005
R210 VTAIL.n163 VTAIL.n162 9.3005
R211 VTAIL.n165 VTAIL.n164 9.3005
R212 VTAIL.n156 VTAIL.n155 9.3005
R213 VTAIL.n171 VTAIL.n170 9.3005
R214 VTAIL.n173 VTAIL.n172 9.3005
R215 VTAIL.n152 VTAIL.n151 9.3005
R216 VTAIL.n180 VTAIL.n179 9.3005
R217 VTAIL.n182 VTAIL.n181 9.3005
R218 VTAIL.n45 VTAIL.n44 9.3005
R219 VTAIL.n4 VTAIL.n3 9.3005
R220 VTAIL.n19 VTAIL.n18 9.3005
R221 VTAIL.n21 VTAIL.n20 9.3005
R222 VTAIL.n12 VTAIL.n11 9.3005
R223 VTAIL.n27 VTAIL.n26 9.3005
R224 VTAIL.n29 VTAIL.n28 9.3005
R225 VTAIL.n8 VTAIL.n7 9.3005
R226 VTAIL.n36 VTAIL.n35 9.3005
R227 VTAIL.n38 VTAIL.n37 9.3005
R228 VTAIL.n118 VTAIL.n117 9.3005
R229 VTAIL.n120 VTAIL.n119 9.3005
R230 VTAIL.n111 VTAIL.n110 9.3005
R231 VTAIL.n126 VTAIL.n125 9.3005
R232 VTAIL.n128 VTAIL.n127 9.3005
R233 VTAIL.n106 VTAIL.n105 9.3005
R234 VTAIL.n134 VTAIL.n133 9.3005
R235 VTAIL.n136 VTAIL.n135 9.3005
R236 VTAIL.n143 VTAIL.n142 9.3005
R237 VTAIL.n102 VTAIL.n101 9.3005
R238 VTAIL.n70 VTAIL.n69 9.3005
R239 VTAIL.n72 VTAIL.n71 9.3005
R240 VTAIL.n63 VTAIL.n62 9.3005
R241 VTAIL.n78 VTAIL.n77 9.3005
R242 VTAIL.n80 VTAIL.n79 9.3005
R243 VTAIL.n58 VTAIL.n57 9.3005
R244 VTAIL.n86 VTAIL.n85 9.3005
R245 VTAIL.n88 VTAIL.n87 9.3005
R246 VTAIL.n95 VTAIL.n94 9.3005
R247 VTAIL.n54 VTAIL.n53 9.3005
R248 VTAIL.n166 VTAIL.n156 8.92171
R249 VTAIL.n22 VTAIL.n12 8.92171
R250 VTAIL.n121 VTAIL.n111 8.92171
R251 VTAIL.n73 VTAIL.n63 8.92171
R252 VTAIL.n165 VTAIL.n158 8.14595
R253 VTAIL.n21 VTAIL.n14 8.14595
R254 VTAIL.n120 VTAIL.n113 8.14595
R255 VTAIL.n72 VTAIL.n65 8.14595
R256 VTAIL.n162 VTAIL.n161 7.3702
R257 VTAIL.n18 VTAIL.n17 7.3702
R258 VTAIL.n117 VTAIL.n116 7.3702
R259 VTAIL.n69 VTAIL.n68 7.3702
R260 VTAIL.n162 VTAIL.n158 5.81868
R261 VTAIL.n18 VTAIL.n14 5.81868
R262 VTAIL.n117 VTAIL.n113 5.81868
R263 VTAIL.n69 VTAIL.n65 5.81868
R264 VTAIL.n166 VTAIL.n165 5.04292
R265 VTAIL.n22 VTAIL.n21 5.04292
R266 VTAIL.n121 VTAIL.n120 5.04292
R267 VTAIL.n73 VTAIL.n72 5.04292
R268 VTAIL.n169 VTAIL.n156 4.26717
R269 VTAIL.n25 VTAIL.n12 4.26717
R270 VTAIL.n124 VTAIL.n111 4.26717
R271 VTAIL.n76 VTAIL.n63 4.26717
R272 VTAIL.n0 VTAIL.t4 3.73242
R273 VTAIL.n0 VTAIL.t1 3.73242
R274 VTAIL.n48 VTAIL.t9 3.73242
R275 VTAIL.n48 VTAIL.t10 3.73242
R276 VTAIL.n98 VTAIL.t7 3.73242
R277 VTAIL.n98 VTAIL.t5 3.73242
R278 VTAIL.n50 VTAIL.t11 3.73242
R279 VTAIL.n50 VTAIL.t0 3.73242
R280 VTAIL.n170 VTAIL.n154 3.49141
R281 VTAIL.n26 VTAIL.n10 3.49141
R282 VTAIL.n125 VTAIL.n109 3.49141
R283 VTAIL.n77 VTAIL.n61 3.49141
R284 VTAIL.n174 VTAIL.n173 2.71565
R285 VTAIL.n30 VTAIL.n29 2.71565
R286 VTAIL.n129 VTAIL.n128 2.71565
R287 VTAIL.n81 VTAIL.n80 2.71565
R288 VTAIL.n163 VTAIL.n159 2.41285
R289 VTAIL.n19 VTAIL.n15 2.41285
R290 VTAIL.n118 VTAIL.n114 2.41285
R291 VTAIL.n70 VTAIL.n66 2.41285
R292 VTAIL.n97 VTAIL.n51 2.27636
R293 VTAIL.n145 VTAIL.n99 2.27636
R294 VTAIL.n49 VTAIL.n47 2.27636
R295 VTAIL.n178 VTAIL.n152 1.93989
R296 VTAIL.n190 VTAIL.n146 1.93989
R297 VTAIL.n34 VTAIL.n8 1.93989
R298 VTAIL.n46 VTAIL.n2 1.93989
R299 VTAIL.n144 VTAIL.n100 1.93989
R300 VTAIL.n132 VTAIL.n106 1.93989
R301 VTAIL.n96 VTAIL.n52 1.93989
R302 VTAIL.n84 VTAIL.n58 1.93989
R303 VTAIL VTAIL.n191 1.64921
R304 VTAIL.n99 VTAIL.n97 1.60826
R305 VTAIL.n47 VTAIL.n1 1.60826
R306 VTAIL.n179 VTAIL.n150 1.16414
R307 VTAIL.n188 VTAIL.n187 1.16414
R308 VTAIL.n35 VTAIL.n6 1.16414
R309 VTAIL.n44 VTAIL.n43 1.16414
R310 VTAIL.n142 VTAIL.n141 1.16414
R311 VTAIL.n133 VTAIL.n104 1.16414
R312 VTAIL.n94 VTAIL.n93 1.16414
R313 VTAIL.n85 VTAIL.n56 1.16414
R314 VTAIL VTAIL.n1 0.627655
R315 VTAIL.n183 VTAIL.n182 0.388379
R316 VTAIL.n184 VTAIL.n148 0.388379
R317 VTAIL.n39 VTAIL.n38 0.388379
R318 VTAIL.n40 VTAIL.n4 0.388379
R319 VTAIL.n138 VTAIL.n102 0.388379
R320 VTAIL.n137 VTAIL.n136 0.388379
R321 VTAIL.n90 VTAIL.n54 0.388379
R322 VTAIL.n89 VTAIL.n88 0.388379
R323 VTAIL.n164 VTAIL.n163 0.155672
R324 VTAIL.n164 VTAIL.n155 0.155672
R325 VTAIL.n171 VTAIL.n155 0.155672
R326 VTAIL.n172 VTAIL.n171 0.155672
R327 VTAIL.n172 VTAIL.n151 0.155672
R328 VTAIL.n180 VTAIL.n151 0.155672
R329 VTAIL.n181 VTAIL.n180 0.155672
R330 VTAIL.n181 VTAIL.n147 0.155672
R331 VTAIL.n189 VTAIL.n147 0.155672
R332 VTAIL.n20 VTAIL.n19 0.155672
R333 VTAIL.n20 VTAIL.n11 0.155672
R334 VTAIL.n27 VTAIL.n11 0.155672
R335 VTAIL.n28 VTAIL.n27 0.155672
R336 VTAIL.n28 VTAIL.n7 0.155672
R337 VTAIL.n36 VTAIL.n7 0.155672
R338 VTAIL.n37 VTAIL.n36 0.155672
R339 VTAIL.n37 VTAIL.n3 0.155672
R340 VTAIL.n45 VTAIL.n3 0.155672
R341 VTAIL.n143 VTAIL.n101 0.155672
R342 VTAIL.n135 VTAIL.n101 0.155672
R343 VTAIL.n135 VTAIL.n134 0.155672
R344 VTAIL.n134 VTAIL.n105 0.155672
R345 VTAIL.n127 VTAIL.n105 0.155672
R346 VTAIL.n127 VTAIL.n126 0.155672
R347 VTAIL.n126 VTAIL.n110 0.155672
R348 VTAIL.n119 VTAIL.n110 0.155672
R349 VTAIL.n119 VTAIL.n118 0.155672
R350 VTAIL.n95 VTAIL.n53 0.155672
R351 VTAIL.n87 VTAIL.n53 0.155672
R352 VTAIL.n87 VTAIL.n86 0.155672
R353 VTAIL.n86 VTAIL.n57 0.155672
R354 VTAIL.n79 VTAIL.n57 0.155672
R355 VTAIL.n79 VTAIL.n78 0.155672
R356 VTAIL.n78 VTAIL.n62 0.155672
R357 VTAIL.n71 VTAIL.n62 0.155672
R358 VTAIL.n71 VTAIL.n70 0.155672
R359 VDD1.n40 VDD1.n0 756.745
R360 VDD1.n85 VDD1.n45 756.745
R361 VDD1.n41 VDD1.n40 585
R362 VDD1.n39 VDD1.n38 585
R363 VDD1.n37 VDD1.n3 585
R364 VDD1.n7 VDD1.n4 585
R365 VDD1.n32 VDD1.n31 585
R366 VDD1.n30 VDD1.n29 585
R367 VDD1.n9 VDD1.n8 585
R368 VDD1.n24 VDD1.n23 585
R369 VDD1.n22 VDD1.n21 585
R370 VDD1.n13 VDD1.n12 585
R371 VDD1.n16 VDD1.n15 585
R372 VDD1.n60 VDD1.n59 585
R373 VDD1.n57 VDD1.n56 585
R374 VDD1.n66 VDD1.n65 585
R375 VDD1.n68 VDD1.n67 585
R376 VDD1.n53 VDD1.n52 585
R377 VDD1.n74 VDD1.n73 585
R378 VDD1.n77 VDD1.n76 585
R379 VDD1.n75 VDD1.n49 585
R380 VDD1.n82 VDD1.n48 585
R381 VDD1.n84 VDD1.n83 585
R382 VDD1.n86 VDD1.n85 585
R383 VDD1.t4 VDD1.n14 329.039
R384 VDD1.t0 VDD1.n58 329.038
R385 VDD1.n40 VDD1.n39 171.744
R386 VDD1.n39 VDD1.n3 171.744
R387 VDD1.n7 VDD1.n3 171.744
R388 VDD1.n31 VDD1.n7 171.744
R389 VDD1.n31 VDD1.n30 171.744
R390 VDD1.n30 VDD1.n8 171.744
R391 VDD1.n23 VDD1.n8 171.744
R392 VDD1.n23 VDD1.n22 171.744
R393 VDD1.n22 VDD1.n12 171.744
R394 VDD1.n15 VDD1.n12 171.744
R395 VDD1.n59 VDD1.n56 171.744
R396 VDD1.n66 VDD1.n56 171.744
R397 VDD1.n67 VDD1.n66 171.744
R398 VDD1.n67 VDD1.n52 171.744
R399 VDD1.n74 VDD1.n52 171.744
R400 VDD1.n76 VDD1.n74 171.744
R401 VDD1.n76 VDD1.n75 171.744
R402 VDD1.n75 VDD1.n48 171.744
R403 VDD1.n84 VDD1.n48 171.744
R404 VDD1.n85 VDD1.n84 171.744
R405 VDD1.n15 VDD1.t4 85.8723
R406 VDD1.n59 VDD1.t0 85.8723
R407 VDD1.n91 VDD1.n90 84.5026
R408 VDD1.n93 VDD1.n92 83.9889
R409 VDD1 VDD1.n44 54.3141
R410 VDD1.n91 VDD1.n89 54.2005
R411 VDD1.n93 VDD1.n91 40.3414
R412 VDD1.n38 VDD1.n37 13.1884
R413 VDD1.n83 VDD1.n82 13.1884
R414 VDD1.n41 VDD1.n2 12.8005
R415 VDD1.n36 VDD1.n4 12.8005
R416 VDD1.n81 VDD1.n49 12.8005
R417 VDD1.n86 VDD1.n47 12.8005
R418 VDD1.n42 VDD1.n0 12.0247
R419 VDD1.n33 VDD1.n32 12.0247
R420 VDD1.n78 VDD1.n77 12.0247
R421 VDD1.n87 VDD1.n45 12.0247
R422 VDD1.n29 VDD1.n6 11.249
R423 VDD1.n73 VDD1.n51 11.249
R424 VDD1.n16 VDD1.n14 10.7239
R425 VDD1.n60 VDD1.n58 10.7239
R426 VDD1.n28 VDD1.n9 10.4732
R427 VDD1.n72 VDD1.n53 10.4732
R428 VDD1.n25 VDD1.n24 9.69747
R429 VDD1.n69 VDD1.n68 9.69747
R430 VDD1.n44 VDD1.n43 9.45567
R431 VDD1.n89 VDD1.n88 9.45567
R432 VDD1.n18 VDD1.n17 9.3005
R433 VDD1.n20 VDD1.n19 9.3005
R434 VDD1.n11 VDD1.n10 9.3005
R435 VDD1.n26 VDD1.n25 9.3005
R436 VDD1.n28 VDD1.n27 9.3005
R437 VDD1.n6 VDD1.n5 9.3005
R438 VDD1.n34 VDD1.n33 9.3005
R439 VDD1.n36 VDD1.n35 9.3005
R440 VDD1.n43 VDD1.n42 9.3005
R441 VDD1.n2 VDD1.n1 9.3005
R442 VDD1.n88 VDD1.n87 9.3005
R443 VDD1.n47 VDD1.n46 9.3005
R444 VDD1.n62 VDD1.n61 9.3005
R445 VDD1.n64 VDD1.n63 9.3005
R446 VDD1.n55 VDD1.n54 9.3005
R447 VDD1.n70 VDD1.n69 9.3005
R448 VDD1.n72 VDD1.n71 9.3005
R449 VDD1.n51 VDD1.n50 9.3005
R450 VDD1.n79 VDD1.n78 9.3005
R451 VDD1.n81 VDD1.n80 9.3005
R452 VDD1.n21 VDD1.n11 8.92171
R453 VDD1.n65 VDD1.n55 8.92171
R454 VDD1.n20 VDD1.n13 8.14595
R455 VDD1.n64 VDD1.n57 8.14595
R456 VDD1.n17 VDD1.n16 7.3702
R457 VDD1.n61 VDD1.n60 7.3702
R458 VDD1.n17 VDD1.n13 5.81868
R459 VDD1.n61 VDD1.n57 5.81868
R460 VDD1.n21 VDD1.n20 5.04292
R461 VDD1.n65 VDD1.n64 5.04292
R462 VDD1.n24 VDD1.n11 4.26717
R463 VDD1.n68 VDD1.n55 4.26717
R464 VDD1.n92 VDD1.t2 3.73242
R465 VDD1.n92 VDD1.t1 3.73242
R466 VDD1.n90 VDD1.t3 3.73242
R467 VDD1.n90 VDD1.t5 3.73242
R468 VDD1.n25 VDD1.n9 3.49141
R469 VDD1.n69 VDD1.n53 3.49141
R470 VDD1.n29 VDD1.n28 2.71565
R471 VDD1.n73 VDD1.n72 2.71565
R472 VDD1.n18 VDD1.n14 2.41285
R473 VDD1.n62 VDD1.n58 2.41285
R474 VDD1.n44 VDD1.n0 1.93989
R475 VDD1.n32 VDD1.n6 1.93989
R476 VDD1.n77 VDD1.n51 1.93989
R477 VDD1.n89 VDD1.n45 1.93989
R478 VDD1.n42 VDD1.n41 1.16414
R479 VDD1.n33 VDD1.n4 1.16414
R480 VDD1.n78 VDD1.n49 1.16414
R481 VDD1.n87 VDD1.n86 1.16414
R482 VDD1 VDD1.n93 0.511276
R483 VDD1.n38 VDD1.n2 0.388379
R484 VDD1.n37 VDD1.n36 0.388379
R485 VDD1.n82 VDD1.n81 0.388379
R486 VDD1.n83 VDD1.n47 0.388379
R487 VDD1.n43 VDD1.n1 0.155672
R488 VDD1.n35 VDD1.n1 0.155672
R489 VDD1.n35 VDD1.n34 0.155672
R490 VDD1.n34 VDD1.n5 0.155672
R491 VDD1.n27 VDD1.n5 0.155672
R492 VDD1.n27 VDD1.n26 0.155672
R493 VDD1.n26 VDD1.n10 0.155672
R494 VDD1.n19 VDD1.n10 0.155672
R495 VDD1.n19 VDD1.n18 0.155672
R496 VDD1.n63 VDD1.n62 0.155672
R497 VDD1.n63 VDD1.n54 0.155672
R498 VDD1.n70 VDD1.n54 0.155672
R499 VDD1.n71 VDD1.n70 0.155672
R500 VDD1.n71 VDD1.n50 0.155672
R501 VDD1.n79 VDD1.n50 0.155672
R502 VDD1.n80 VDD1.n79 0.155672
R503 VDD1.n80 VDD1.n46 0.155672
R504 VDD1.n88 VDD1.n46 0.155672
R505 VN.n25 VN.n14 161.3
R506 VN.n24 VN.n23 161.3
R507 VN.n22 VN.n15 161.3
R508 VN.n21 VN.n20 161.3
R509 VN.n19 VN.n16 161.3
R510 VN.n11 VN.n0 161.3
R511 VN.n10 VN.n9 161.3
R512 VN.n8 VN.n1 161.3
R513 VN.n7 VN.n6 161.3
R514 VN.n5 VN.n2 161.3
R515 VN.n3 VN.t0 124.624
R516 VN.n17 VN.t3 124.624
R517 VN.n13 VN.n12 91.6722
R518 VN.n27 VN.n26 91.6722
R519 VN.n4 VN.t4 90.8711
R520 VN.n12 VN.t1 90.8711
R521 VN.n18 VN.t5 90.8711
R522 VN.n26 VN.t2 90.8711
R523 VN.n4 VN.n3 59.2346
R524 VN.n18 VN.n17 59.2346
R525 VN.n10 VN.n1 47.2923
R526 VN.n24 VN.n15 47.2923
R527 VN VN.n27 45.4148
R528 VN.n6 VN.n1 33.6945
R529 VN.n20 VN.n15 33.6945
R530 VN.n6 VN.n5 24.4675
R531 VN.n11 VN.n10 24.4675
R532 VN.n20 VN.n19 24.4675
R533 VN.n25 VN.n24 24.4675
R534 VN.n12 VN.n11 19.0848
R535 VN.n26 VN.n25 19.0848
R536 VN.n5 VN.n4 12.234
R537 VN.n19 VN.n18 12.234
R538 VN.n17 VN.n16 9.06133
R539 VN.n3 VN.n2 9.06133
R540 VN.n27 VN.n14 0.278367
R541 VN.n13 VN.n0 0.278367
R542 VN.n23 VN.n14 0.189894
R543 VN.n23 VN.n22 0.189894
R544 VN.n22 VN.n21 0.189894
R545 VN.n21 VN.n16 0.189894
R546 VN.n7 VN.n2 0.189894
R547 VN.n8 VN.n7 0.189894
R548 VN.n9 VN.n8 0.189894
R549 VN.n9 VN.n0 0.189894
R550 VN VN.n13 0.153454
R551 VDD2.n87 VDD2.n47 756.745
R552 VDD2.n40 VDD2.n0 756.745
R553 VDD2.n88 VDD2.n87 585
R554 VDD2.n86 VDD2.n85 585
R555 VDD2.n84 VDD2.n50 585
R556 VDD2.n54 VDD2.n51 585
R557 VDD2.n79 VDD2.n78 585
R558 VDD2.n77 VDD2.n76 585
R559 VDD2.n56 VDD2.n55 585
R560 VDD2.n71 VDD2.n70 585
R561 VDD2.n69 VDD2.n68 585
R562 VDD2.n60 VDD2.n59 585
R563 VDD2.n63 VDD2.n62 585
R564 VDD2.n15 VDD2.n14 585
R565 VDD2.n12 VDD2.n11 585
R566 VDD2.n21 VDD2.n20 585
R567 VDD2.n23 VDD2.n22 585
R568 VDD2.n8 VDD2.n7 585
R569 VDD2.n29 VDD2.n28 585
R570 VDD2.n32 VDD2.n31 585
R571 VDD2.n30 VDD2.n4 585
R572 VDD2.n37 VDD2.n3 585
R573 VDD2.n39 VDD2.n38 585
R574 VDD2.n41 VDD2.n40 585
R575 VDD2.t3 VDD2.n61 329.039
R576 VDD2.t5 VDD2.n13 329.038
R577 VDD2.n87 VDD2.n86 171.744
R578 VDD2.n86 VDD2.n50 171.744
R579 VDD2.n54 VDD2.n50 171.744
R580 VDD2.n78 VDD2.n54 171.744
R581 VDD2.n78 VDD2.n77 171.744
R582 VDD2.n77 VDD2.n55 171.744
R583 VDD2.n70 VDD2.n55 171.744
R584 VDD2.n70 VDD2.n69 171.744
R585 VDD2.n69 VDD2.n59 171.744
R586 VDD2.n62 VDD2.n59 171.744
R587 VDD2.n14 VDD2.n11 171.744
R588 VDD2.n21 VDD2.n11 171.744
R589 VDD2.n22 VDD2.n21 171.744
R590 VDD2.n22 VDD2.n7 171.744
R591 VDD2.n29 VDD2.n7 171.744
R592 VDD2.n31 VDD2.n29 171.744
R593 VDD2.n31 VDD2.n30 171.744
R594 VDD2.n30 VDD2.n3 171.744
R595 VDD2.n39 VDD2.n3 171.744
R596 VDD2.n40 VDD2.n39 171.744
R597 VDD2.n62 VDD2.t3 85.8723
R598 VDD2.n14 VDD2.t5 85.8723
R599 VDD2.n46 VDD2.n45 84.5026
R600 VDD2 VDD2.n93 84.4997
R601 VDD2.n46 VDD2.n44 54.2005
R602 VDD2.n92 VDD2.n91 52.549
R603 VDD2.n92 VDD2.n46 38.6205
R604 VDD2.n85 VDD2.n84 13.1884
R605 VDD2.n38 VDD2.n37 13.1884
R606 VDD2.n88 VDD2.n49 12.8005
R607 VDD2.n83 VDD2.n51 12.8005
R608 VDD2.n36 VDD2.n4 12.8005
R609 VDD2.n41 VDD2.n2 12.8005
R610 VDD2.n89 VDD2.n47 12.0247
R611 VDD2.n80 VDD2.n79 12.0247
R612 VDD2.n33 VDD2.n32 12.0247
R613 VDD2.n42 VDD2.n0 12.0247
R614 VDD2.n76 VDD2.n53 11.249
R615 VDD2.n28 VDD2.n6 11.249
R616 VDD2.n63 VDD2.n61 10.7239
R617 VDD2.n15 VDD2.n13 10.7239
R618 VDD2.n75 VDD2.n56 10.4732
R619 VDD2.n27 VDD2.n8 10.4732
R620 VDD2.n72 VDD2.n71 9.69747
R621 VDD2.n24 VDD2.n23 9.69747
R622 VDD2.n91 VDD2.n90 9.45567
R623 VDD2.n44 VDD2.n43 9.45567
R624 VDD2.n65 VDD2.n64 9.3005
R625 VDD2.n67 VDD2.n66 9.3005
R626 VDD2.n58 VDD2.n57 9.3005
R627 VDD2.n73 VDD2.n72 9.3005
R628 VDD2.n75 VDD2.n74 9.3005
R629 VDD2.n53 VDD2.n52 9.3005
R630 VDD2.n81 VDD2.n80 9.3005
R631 VDD2.n83 VDD2.n82 9.3005
R632 VDD2.n90 VDD2.n89 9.3005
R633 VDD2.n49 VDD2.n48 9.3005
R634 VDD2.n43 VDD2.n42 9.3005
R635 VDD2.n2 VDD2.n1 9.3005
R636 VDD2.n17 VDD2.n16 9.3005
R637 VDD2.n19 VDD2.n18 9.3005
R638 VDD2.n10 VDD2.n9 9.3005
R639 VDD2.n25 VDD2.n24 9.3005
R640 VDD2.n27 VDD2.n26 9.3005
R641 VDD2.n6 VDD2.n5 9.3005
R642 VDD2.n34 VDD2.n33 9.3005
R643 VDD2.n36 VDD2.n35 9.3005
R644 VDD2.n68 VDD2.n58 8.92171
R645 VDD2.n20 VDD2.n10 8.92171
R646 VDD2.n67 VDD2.n60 8.14595
R647 VDD2.n19 VDD2.n12 8.14595
R648 VDD2.n64 VDD2.n63 7.3702
R649 VDD2.n16 VDD2.n15 7.3702
R650 VDD2.n64 VDD2.n60 5.81868
R651 VDD2.n16 VDD2.n12 5.81868
R652 VDD2.n68 VDD2.n67 5.04292
R653 VDD2.n20 VDD2.n19 5.04292
R654 VDD2.n71 VDD2.n58 4.26717
R655 VDD2.n23 VDD2.n10 4.26717
R656 VDD2.n93 VDD2.t0 3.73242
R657 VDD2.n93 VDD2.t2 3.73242
R658 VDD2.n45 VDD2.t1 3.73242
R659 VDD2.n45 VDD2.t4 3.73242
R660 VDD2.n72 VDD2.n56 3.49141
R661 VDD2.n24 VDD2.n8 3.49141
R662 VDD2.n76 VDD2.n75 2.71565
R663 VDD2.n28 VDD2.n27 2.71565
R664 VDD2.n65 VDD2.n61 2.41285
R665 VDD2.n17 VDD2.n13 2.41285
R666 VDD2.n91 VDD2.n47 1.93989
R667 VDD2.n79 VDD2.n53 1.93989
R668 VDD2.n32 VDD2.n6 1.93989
R669 VDD2.n44 VDD2.n0 1.93989
R670 VDD2 VDD2.n92 1.76559
R671 VDD2.n89 VDD2.n88 1.16414
R672 VDD2.n80 VDD2.n51 1.16414
R673 VDD2.n33 VDD2.n4 1.16414
R674 VDD2.n42 VDD2.n41 1.16414
R675 VDD2.n85 VDD2.n49 0.388379
R676 VDD2.n84 VDD2.n83 0.388379
R677 VDD2.n37 VDD2.n36 0.388379
R678 VDD2.n38 VDD2.n2 0.388379
R679 VDD2.n90 VDD2.n48 0.155672
R680 VDD2.n82 VDD2.n48 0.155672
R681 VDD2.n82 VDD2.n81 0.155672
R682 VDD2.n81 VDD2.n52 0.155672
R683 VDD2.n74 VDD2.n52 0.155672
R684 VDD2.n74 VDD2.n73 0.155672
R685 VDD2.n73 VDD2.n57 0.155672
R686 VDD2.n66 VDD2.n57 0.155672
R687 VDD2.n66 VDD2.n65 0.155672
R688 VDD2.n18 VDD2.n17 0.155672
R689 VDD2.n18 VDD2.n9 0.155672
R690 VDD2.n25 VDD2.n9 0.155672
R691 VDD2.n26 VDD2.n25 0.155672
R692 VDD2.n26 VDD2.n5 0.155672
R693 VDD2.n34 VDD2.n5 0.155672
R694 VDD2.n35 VDD2.n34 0.155672
R695 VDD2.n35 VDD2.n1 0.155672
R696 VDD2.n43 VDD2.n1 0.155672
R697 B.n449 B.n62 585
R698 B.n451 B.n450 585
R699 B.n452 B.n61 585
R700 B.n454 B.n453 585
R701 B.n455 B.n60 585
R702 B.n457 B.n456 585
R703 B.n458 B.n59 585
R704 B.n460 B.n459 585
R705 B.n461 B.n58 585
R706 B.n463 B.n462 585
R707 B.n464 B.n57 585
R708 B.n466 B.n465 585
R709 B.n467 B.n56 585
R710 B.n469 B.n468 585
R711 B.n470 B.n55 585
R712 B.n472 B.n471 585
R713 B.n473 B.n54 585
R714 B.n475 B.n474 585
R715 B.n476 B.n53 585
R716 B.n478 B.n477 585
R717 B.n479 B.n52 585
R718 B.n481 B.n480 585
R719 B.n482 B.n51 585
R720 B.n484 B.n483 585
R721 B.n485 B.n50 585
R722 B.n487 B.n486 585
R723 B.n488 B.n49 585
R724 B.n490 B.n489 585
R725 B.n491 B.n48 585
R726 B.n493 B.n492 585
R727 B.n494 B.n47 585
R728 B.n496 B.n495 585
R729 B.n498 B.n497 585
R730 B.n499 B.n43 585
R731 B.n501 B.n500 585
R732 B.n502 B.n42 585
R733 B.n504 B.n503 585
R734 B.n505 B.n41 585
R735 B.n507 B.n506 585
R736 B.n508 B.n40 585
R737 B.n510 B.n509 585
R738 B.n512 B.n37 585
R739 B.n514 B.n513 585
R740 B.n515 B.n36 585
R741 B.n517 B.n516 585
R742 B.n518 B.n35 585
R743 B.n520 B.n519 585
R744 B.n521 B.n34 585
R745 B.n523 B.n522 585
R746 B.n524 B.n33 585
R747 B.n526 B.n525 585
R748 B.n527 B.n32 585
R749 B.n529 B.n528 585
R750 B.n530 B.n31 585
R751 B.n532 B.n531 585
R752 B.n533 B.n30 585
R753 B.n535 B.n534 585
R754 B.n536 B.n29 585
R755 B.n538 B.n537 585
R756 B.n539 B.n28 585
R757 B.n541 B.n540 585
R758 B.n542 B.n27 585
R759 B.n544 B.n543 585
R760 B.n545 B.n26 585
R761 B.n547 B.n546 585
R762 B.n548 B.n25 585
R763 B.n550 B.n549 585
R764 B.n551 B.n24 585
R765 B.n553 B.n552 585
R766 B.n554 B.n23 585
R767 B.n556 B.n555 585
R768 B.n557 B.n22 585
R769 B.n559 B.n558 585
R770 B.n448 B.n447 585
R771 B.n446 B.n63 585
R772 B.n445 B.n444 585
R773 B.n443 B.n64 585
R774 B.n442 B.n441 585
R775 B.n440 B.n65 585
R776 B.n439 B.n438 585
R777 B.n437 B.n66 585
R778 B.n436 B.n435 585
R779 B.n434 B.n67 585
R780 B.n433 B.n432 585
R781 B.n431 B.n68 585
R782 B.n430 B.n429 585
R783 B.n428 B.n69 585
R784 B.n427 B.n426 585
R785 B.n425 B.n70 585
R786 B.n424 B.n423 585
R787 B.n422 B.n71 585
R788 B.n421 B.n420 585
R789 B.n419 B.n72 585
R790 B.n418 B.n417 585
R791 B.n416 B.n73 585
R792 B.n415 B.n414 585
R793 B.n413 B.n74 585
R794 B.n412 B.n411 585
R795 B.n410 B.n75 585
R796 B.n409 B.n408 585
R797 B.n407 B.n76 585
R798 B.n406 B.n405 585
R799 B.n404 B.n77 585
R800 B.n403 B.n402 585
R801 B.n401 B.n78 585
R802 B.n400 B.n399 585
R803 B.n398 B.n79 585
R804 B.n397 B.n396 585
R805 B.n395 B.n80 585
R806 B.n394 B.n393 585
R807 B.n392 B.n81 585
R808 B.n391 B.n390 585
R809 B.n389 B.n82 585
R810 B.n388 B.n387 585
R811 B.n386 B.n83 585
R812 B.n385 B.n384 585
R813 B.n383 B.n84 585
R814 B.n382 B.n381 585
R815 B.n380 B.n85 585
R816 B.n379 B.n378 585
R817 B.n377 B.n86 585
R818 B.n376 B.n375 585
R819 B.n374 B.n87 585
R820 B.n373 B.n372 585
R821 B.n371 B.n88 585
R822 B.n370 B.n369 585
R823 B.n368 B.n89 585
R824 B.n367 B.n366 585
R825 B.n365 B.n90 585
R826 B.n364 B.n363 585
R827 B.n362 B.n91 585
R828 B.n361 B.n360 585
R829 B.n359 B.n92 585
R830 B.n358 B.n357 585
R831 B.n356 B.n93 585
R832 B.n355 B.n354 585
R833 B.n353 B.n94 585
R834 B.n352 B.n351 585
R835 B.n350 B.n95 585
R836 B.n349 B.n348 585
R837 B.n347 B.n96 585
R838 B.n346 B.n345 585
R839 B.n344 B.n97 585
R840 B.n343 B.n342 585
R841 B.n341 B.n98 585
R842 B.n340 B.n339 585
R843 B.n338 B.n99 585
R844 B.n337 B.n336 585
R845 B.n335 B.n100 585
R846 B.n334 B.n333 585
R847 B.n332 B.n101 585
R848 B.n331 B.n330 585
R849 B.n220 B.n219 585
R850 B.n221 B.n142 585
R851 B.n223 B.n222 585
R852 B.n224 B.n141 585
R853 B.n226 B.n225 585
R854 B.n227 B.n140 585
R855 B.n229 B.n228 585
R856 B.n230 B.n139 585
R857 B.n232 B.n231 585
R858 B.n233 B.n138 585
R859 B.n235 B.n234 585
R860 B.n236 B.n137 585
R861 B.n238 B.n237 585
R862 B.n239 B.n136 585
R863 B.n241 B.n240 585
R864 B.n242 B.n135 585
R865 B.n244 B.n243 585
R866 B.n245 B.n134 585
R867 B.n247 B.n246 585
R868 B.n248 B.n133 585
R869 B.n250 B.n249 585
R870 B.n251 B.n132 585
R871 B.n253 B.n252 585
R872 B.n254 B.n131 585
R873 B.n256 B.n255 585
R874 B.n257 B.n130 585
R875 B.n259 B.n258 585
R876 B.n260 B.n129 585
R877 B.n262 B.n261 585
R878 B.n263 B.n128 585
R879 B.n265 B.n264 585
R880 B.n266 B.n125 585
R881 B.n269 B.n268 585
R882 B.n270 B.n124 585
R883 B.n272 B.n271 585
R884 B.n273 B.n123 585
R885 B.n275 B.n274 585
R886 B.n276 B.n122 585
R887 B.n278 B.n277 585
R888 B.n279 B.n121 585
R889 B.n281 B.n280 585
R890 B.n283 B.n282 585
R891 B.n284 B.n117 585
R892 B.n286 B.n285 585
R893 B.n287 B.n116 585
R894 B.n289 B.n288 585
R895 B.n290 B.n115 585
R896 B.n292 B.n291 585
R897 B.n293 B.n114 585
R898 B.n295 B.n294 585
R899 B.n296 B.n113 585
R900 B.n298 B.n297 585
R901 B.n299 B.n112 585
R902 B.n301 B.n300 585
R903 B.n302 B.n111 585
R904 B.n304 B.n303 585
R905 B.n305 B.n110 585
R906 B.n307 B.n306 585
R907 B.n308 B.n109 585
R908 B.n310 B.n309 585
R909 B.n311 B.n108 585
R910 B.n313 B.n312 585
R911 B.n314 B.n107 585
R912 B.n316 B.n315 585
R913 B.n317 B.n106 585
R914 B.n319 B.n318 585
R915 B.n320 B.n105 585
R916 B.n322 B.n321 585
R917 B.n323 B.n104 585
R918 B.n325 B.n324 585
R919 B.n326 B.n103 585
R920 B.n328 B.n327 585
R921 B.n329 B.n102 585
R922 B.n218 B.n143 585
R923 B.n217 B.n216 585
R924 B.n215 B.n144 585
R925 B.n214 B.n213 585
R926 B.n212 B.n145 585
R927 B.n211 B.n210 585
R928 B.n209 B.n146 585
R929 B.n208 B.n207 585
R930 B.n206 B.n147 585
R931 B.n205 B.n204 585
R932 B.n203 B.n148 585
R933 B.n202 B.n201 585
R934 B.n200 B.n149 585
R935 B.n199 B.n198 585
R936 B.n197 B.n150 585
R937 B.n196 B.n195 585
R938 B.n194 B.n151 585
R939 B.n193 B.n192 585
R940 B.n191 B.n152 585
R941 B.n190 B.n189 585
R942 B.n188 B.n153 585
R943 B.n187 B.n186 585
R944 B.n185 B.n154 585
R945 B.n184 B.n183 585
R946 B.n182 B.n155 585
R947 B.n181 B.n180 585
R948 B.n179 B.n156 585
R949 B.n178 B.n177 585
R950 B.n176 B.n157 585
R951 B.n175 B.n174 585
R952 B.n173 B.n158 585
R953 B.n172 B.n171 585
R954 B.n170 B.n159 585
R955 B.n169 B.n168 585
R956 B.n167 B.n160 585
R957 B.n166 B.n165 585
R958 B.n164 B.n161 585
R959 B.n163 B.n162 585
R960 B.n2 B.n0 585
R961 B.n617 B.n1 585
R962 B.n616 B.n615 585
R963 B.n614 B.n3 585
R964 B.n613 B.n612 585
R965 B.n611 B.n4 585
R966 B.n610 B.n609 585
R967 B.n608 B.n5 585
R968 B.n607 B.n606 585
R969 B.n605 B.n6 585
R970 B.n604 B.n603 585
R971 B.n602 B.n7 585
R972 B.n601 B.n600 585
R973 B.n599 B.n8 585
R974 B.n598 B.n597 585
R975 B.n596 B.n9 585
R976 B.n595 B.n594 585
R977 B.n593 B.n10 585
R978 B.n592 B.n591 585
R979 B.n590 B.n11 585
R980 B.n589 B.n588 585
R981 B.n587 B.n12 585
R982 B.n586 B.n585 585
R983 B.n584 B.n13 585
R984 B.n583 B.n582 585
R985 B.n581 B.n14 585
R986 B.n580 B.n579 585
R987 B.n578 B.n15 585
R988 B.n577 B.n576 585
R989 B.n575 B.n16 585
R990 B.n574 B.n573 585
R991 B.n572 B.n17 585
R992 B.n571 B.n570 585
R993 B.n569 B.n18 585
R994 B.n568 B.n567 585
R995 B.n566 B.n19 585
R996 B.n565 B.n564 585
R997 B.n563 B.n20 585
R998 B.n562 B.n561 585
R999 B.n560 B.n21 585
R1000 B.n619 B.n618 585
R1001 B.n220 B.n143 564.573
R1002 B.n558 B.n21 564.573
R1003 B.n330 B.n329 564.573
R1004 B.n449 B.n448 564.573
R1005 B.n118 B.t8 367.676
R1006 B.n44 B.t1 367.676
R1007 B.n126 B.t11 367.676
R1008 B.n38 B.t4 367.676
R1009 B.n119 B.t7 316.476
R1010 B.n45 B.t2 316.476
R1011 B.n127 B.t10 316.476
R1012 B.n39 B.t5 316.476
R1013 B.n118 B.t6 298.433
R1014 B.n126 B.t9 298.433
R1015 B.n38 B.t3 298.433
R1016 B.n44 B.t0 298.433
R1017 B.n216 B.n143 163.367
R1018 B.n216 B.n215 163.367
R1019 B.n215 B.n214 163.367
R1020 B.n214 B.n145 163.367
R1021 B.n210 B.n145 163.367
R1022 B.n210 B.n209 163.367
R1023 B.n209 B.n208 163.367
R1024 B.n208 B.n147 163.367
R1025 B.n204 B.n147 163.367
R1026 B.n204 B.n203 163.367
R1027 B.n203 B.n202 163.367
R1028 B.n202 B.n149 163.367
R1029 B.n198 B.n149 163.367
R1030 B.n198 B.n197 163.367
R1031 B.n197 B.n196 163.367
R1032 B.n196 B.n151 163.367
R1033 B.n192 B.n151 163.367
R1034 B.n192 B.n191 163.367
R1035 B.n191 B.n190 163.367
R1036 B.n190 B.n153 163.367
R1037 B.n186 B.n153 163.367
R1038 B.n186 B.n185 163.367
R1039 B.n185 B.n184 163.367
R1040 B.n184 B.n155 163.367
R1041 B.n180 B.n155 163.367
R1042 B.n180 B.n179 163.367
R1043 B.n179 B.n178 163.367
R1044 B.n178 B.n157 163.367
R1045 B.n174 B.n157 163.367
R1046 B.n174 B.n173 163.367
R1047 B.n173 B.n172 163.367
R1048 B.n172 B.n159 163.367
R1049 B.n168 B.n159 163.367
R1050 B.n168 B.n167 163.367
R1051 B.n167 B.n166 163.367
R1052 B.n166 B.n161 163.367
R1053 B.n162 B.n161 163.367
R1054 B.n162 B.n2 163.367
R1055 B.n618 B.n2 163.367
R1056 B.n618 B.n617 163.367
R1057 B.n617 B.n616 163.367
R1058 B.n616 B.n3 163.367
R1059 B.n612 B.n3 163.367
R1060 B.n612 B.n611 163.367
R1061 B.n611 B.n610 163.367
R1062 B.n610 B.n5 163.367
R1063 B.n606 B.n5 163.367
R1064 B.n606 B.n605 163.367
R1065 B.n605 B.n604 163.367
R1066 B.n604 B.n7 163.367
R1067 B.n600 B.n7 163.367
R1068 B.n600 B.n599 163.367
R1069 B.n599 B.n598 163.367
R1070 B.n598 B.n9 163.367
R1071 B.n594 B.n9 163.367
R1072 B.n594 B.n593 163.367
R1073 B.n593 B.n592 163.367
R1074 B.n592 B.n11 163.367
R1075 B.n588 B.n11 163.367
R1076 B.n588 B.n587 163.367
R1077 B.n587 B.n586 163.367
R1078 B.n586 B.n13 163.367
R1079 B.n582 B.n13 163.367
R1080 B.n582 B.n581 163.367
R1081 B.n581 B.n580 163.367
R1082 B.n580 B.n15 163.367
R1083 B.n576 B.n15 163.367
R1084 B.n576 B.n575 163.367
R1085 B.n575 B.n574 163.367
R1086 B.n574 B.n17 163.367
R1087 B.n570 B.n17 163.367
R1088 B.n570 B.n569 163.367
R1089 B.n569 B.n568 163.367
R1090 B.n568 B.n19 163.367
R1091 B.n564 B.n19 163.367
R1092 B.n564 B.n563 163.367
R1093 B.n563 B.n562 163.367
R1094 B.n562 B.n21 163.367
R1095 B.n221 B.n220 163.367
R1096 B.n222 B.n221 163.367
R1097 B.n222 B.n141 163.367
R1098 B.n226 B.n141 163.367
R1099 B.n227 B.n226 163.367
R1100 B.n228 B.n227 163.367
R1101 B.n228 B.n139 163.367
R1102 B.n232 B.n139 163.367
R1103 B.n233 B.n232 163.367
R1104 B.n234 B.n233 163.367
R1105 B.n234 B.n137 163.367
R1106 B.n238 B.n137 163.367
R1107 B.n239 B.n238 163.367
R1108 B.n240 B.n239 163.367
R1109 B.n240 B.n135 163.367
R1110 B.n244 B.n135 163.367
R1111 B.n245 B.n244 163.367
R1112 B.n246 B.n245 163.367
R1113 B.n246 B.n133 163.367
R1114 B.n250 B.n133 163.367
R1115 B.n251 B.n250 163.367
R1116 B.n252 B.n251 163.367
R1117 B.n252 B.n131 163.367
R1118 B.n256 B.n131 163.367
R1119 B.n257 B.n256 163.367
R1120 B.n258 B.n257 163.367
R1121 B.n258 B.n129 163.367
R1122 B.n262 B.n129 163.367
R1123 B.n263 B.n262 163.367
R1124 B.n264 B.n263 163.367
R1125 B.n264 B.n125 163.367
R1126 B.n269 B.n125 163.367
R1127 B.n270 B.n269 163.367
R1128 B.n271 B.n270 163.367
R1129 B.n271 B.n123 163.367
R1130 B.n275 B.n123 163.367
R1131 B.n276 B.n275 163.367
R1132 B.n277 B.n276 163.367
R1133 B.n277 B.n121 163.367
R1134 B.n281 B.n121 163.367
R1135 B.n282 B.n281 163.367
R1136 B.n282 B.n117 163.367
R1137 B.n286 B.n117 163.367
R1138 B.n287 B.n286 163.367
R1139 B.n288 B.n287 163.367
R1140 B.n288 B.n115 163.367
R1141 B.n292 B.n115 163.367
R1142 B.n293 B.n292 163.367
R1143 B.n294 B.n293 163.367
R1144 B.n294 B.n113 163.367
R1145 B.n298 B.n113 163.367
R1146 B.n299 B.n298 163.367
R1147 B.n300 B.n299 163.367
R1148 B.n300 B.n111 163.367
R1149 B.n304 B.n111 163.367
R1150 B.n305 B.n304 163.367
R1151 B.n306 B.n305 163.367
R1152 B.n306 B.n109 163.367
R1153 B.n310 B.n109 163.367
R1154 B.n311 B.n310 163.367
R1155 B.n312 B.n311 163.367
R1156 B.n312 B.n107 163.367
R1157 B.n316 B.n107 163.367
R1158 B.n317 B.n316 163.367
R1159 B.n318 B.n317 163.367
R1160 B.n318 B.n105 163.367
R1161 B.n322 B.n105 163.367
R1162 B.n323 B.n322 163.367
R1163 B.n324 B.n323 163.367
R1164 B.n324 B.n103 163.367
R1165 B.n328 B.n103 163.367
R1166 B.n329 B.n328 163.367
R1167 B.n330 B.n101 163.367
R1168 B.n334 B.n101 163.367
R1169 B.n335 B.n334 163.367
R1170 B.n336 B.n335 163.367
R1171 B.n336 B.n99 163.367
R1172 B.n340 B.n99 163.367
R1173 B.n341 B.n340 163.367
R1174 B.n342 B.n341 163.367
R1175 B.n342 B.n97 163.367
R1176 B.n346 B.n97 163.367
R1177 B.n347 B.n346 163.367
R1178 B.n348 B.n347 163.367
R1179 B.n348 B.n95 163.367
R1180 B.n352 B.n95 163.367
R1181 B.n353 B.n352 163.367
R1182 B.n354 B.n353 163.367
R1183 B.n354 B.n93 163.367
R1184 B.n358 B.n93 163.367
R1185 B.n359 B.n358 163.367
R1186 B.n360 B.n359 163.367
R1187 B.n360 B.n91 163.367
R1188 B.n364 B.n91 163.367
R1189 B.n365 B.n364 163.367
R1190 B.n366 B.n365 163.367
R1191 B.n366 B.n89 163.367
R1192 B.n370 B.n89 163.367
R1193 B.n371 B.n370 163.367
R1194 B.n372 B.n371 163.367
R1195 B.n372 B.n87 163.367
R1196 B.n376 B.n87 163.367
R1197 B.n377 B.n376 163.367
R1198 B.n378 B.n377 163.367
R1199 B.n378 B.n85 163.367
R1200 B.n382 B.n85 163.367
R1201 B.n383 B.n382 163.367
R1202 B.n384 B.n383 163.367
R1203 B.n384 B.n83 163.367
R1204 B.n388 B.n83 163.367
R1205 B.n389 B.n388 163.367
R1206 B.n390 B.n389 163.367
R1207 B.n390 B.n81 163.367
R1208 B.n394 B.n81 163.367
R1209 B.n395 B.n394 163.367
R1210 B.n396 B.n395 163.367
R1211 B.n396 B.n79 163.367
R1212 B.n400 B.n79 163.367
R1213 B.n401 B.n400 163.367
R1214 B.n402 B.n401 163.367
R1215 B.n402 B.n77 163.367
R1216 B.n406 B.n77 163.367
R1217 B.n407 B.n406 163.367
R1218 B.n408 B.n407 163.367
R1219 B.n408 B.n75 163.367
R1220 B.n412 B.n75 163.367
R1221 B.n413 B.n412 163.367
R1222 B.n414 B.n413 163.367
R1223 B.n414 B.n73 163.367
R1224 B.n418 B.n73 163.367
R1225 B.n419 B.n418 163.367
R1226 B.n420 B.n419 163.367
R1227 B.n420 B.n71 163.367
R1228 B.n424 B.n71 163.367
R1229 B.n425 B.n424 163.367
R1230 B.n426 B.n425 163.367
R1231 B.n426 B.n69 163.367
R1232 B.n430 B.n69 163.367
R1233 B.n431 B.n430 163.367
R1234 B.n432 B.n431 163.367
R1235 B.n432 B.n67 163.367
R1236 B.n436 B.n67 163.367
R1237 B.n437 B.n436 163.367
R1238 B.n438 B.n437 163.367
R1239 B.n438 B.n65 163.367
R1240 B.n442 B.n65 163.367
R1241 B.n443 B.n442 163.367
R1242 B.n444 B.n443 163.367
R1243 B.n444 B.n63 163.367
R1244 B.n448 B.n63 163.367
R1245 B.n558 B.n557 163.367
R1246 B.n557 B.n556 163.367
R1247 B.n556 B.n23 163.367
R1248 B.n552 B.n23 163.367
R1249 B.n552 B.n551 163.367
R1250 B.n551 B.n550 163.367
R1251 B.n550 B.n25 163.367
R1252 B.n546 B.n25 163.367
R1253 B.n546 B.n545 163.367
R1254 B.n545 B.n544 163.367
R1255 B.n544 B.n27 163.367
R1256 B.n540 B.n27 163.367
R1257 B.n540 B.n539 163.367
R1258 B.n539 B.n538 163.367
R1259 B.n538 B.n29 163.367
R1260 B.n534 B.n29 163.367
R1261 B.n534 B.n533 163.367
R1262 B.n533 B.n532 163.367
R1263 B.n532 B.n31 163.367
R1264 B.n528 B.n31 163.367
R1265 B.n528 B.n527 163.367
R1266 B.n527 B.n526 163.367
R1267 B.n526 B.n33 163.367
R1268 B.n522 B.n33 163.367
R1269 B.n522 B.n521 163.367
R1270 B.n521 B.n520 163.367
R1271 B.n520 B.n35 163.367
R1272 B.n516 B.n35 163.367
R1273 B.n516 B.n515 163.367
R1274 B.n515 B.n514 163.367
R1275 B.n514 B.n37 163.367
R1276 B.n509 B.n37 163.367
R1277 B.n509 B.n508 163.367
R1278 B.n508 B.n507 163.367
R1279 B.n507 B.n41 163.367
R1280 B.n503 B.n41 163.367
R1281 B.n503 B.n502 163.367
R1282 B.n502 B.n501 163.367
R1283 B.n501 B.n43 163.367
R1284 B.n497 B.n43 163.367
R1285 B.n497 B.n496 163.367
R1286 B.n496 B.n47 163.367
R1287 B.n492 B.n47 163.367
R1288 B.n492 B.n491 163.367
R1289 B.n491 B.n490 163.367
R1290 B.n490 B.n49 163.367
R1291 B.n486 B.n49 163.367
R1292 B.n486 B.n485 163.367
R1293 B.n485 B.n484 163.367
R1294 B.n484 B.n51 163.367
R1295 B.n480 B.n51 163.367
R1296 B.n480 B.n479 163.367
R1297 B.n479 B.n478 163.367
R1298 B.n478 B.n53 163.367
R1299 B.n474 B.n53 163.367
R1300 B.n474 B.n473 163.367
R1301 B.n473 B.n472 163.367
R1302 B.n472 B.n55 163.367
R1303 B.n468 B.n55 163.367
R1304 B.n468 B.n467 163.367
R1305 B.n467 B.n466 163.367
R1306 B.n466 B.n57 163.367
R1307 B.n462 B.n57 163.367
R1308 B.n462 B.n461 163.367
R1309 B.n461 B.n460 163.367
R1310 B.n460 B.n59 163.367
R1311 B.n456 B.n59 163.367
R1312 B.n456 B.n455 163.367
R1313 B.n455 B.n454 163.367
R1314 B.n454 B.n61 163.367
R1315 B.n450 B.n61 163.367
R1316 B.n450 B.n449 163.367
R1317 B.n120 B.n119 59.5399
R1318 B.n267 B.n127 59.5399
R1319 B.n511 B.n39 59.5399
R1320 B.n46 B.n45 59.5399
R1321 B.n119 B.n118 51.2005
R1322 B.n127 B.n126 51.2005
R1323 B.n39 B.n38 51.2005
R1324 B.n45 B.n44 51.2005
R1325 B.n560 B.n559 36.6834
R1326 B.n447 B.n62 36.6834
R1327 B.n331 B.n102 36.6834
R1328 B.n219 B.n218 36.6834
R1329 B B.n619 18.0485
R1330 B.n559 B.n22 10.6151
R1331 B.n555 B.n22 10.6151
R1332 B.n555 B.n554 10.6151
R1333 B.n554 B.n553 10.6151
R1334 B.n553 B.n24 10.6151
R1335 B.n549 B.n24 10.6151
R1336 B.n549 B.n548 10.6151
R1337 B.n548 B.n547 10.6151
R1338 B.n547 B.n26 10.6151
R1339 B.n543 B.n26 10.6151
R1340 B.n543 B.n542 10.6151
R1341 B.n542 B.n541 10.6151
R1342 B.n541 B.n28 10.6151
R1343 B.n537 B.n28 10.6151
R1344 B.n537 B.n536 10.6151
R1345 B.n536 B.n535 10.6151
R1346 B.n535 B.n30 10.6151
R1347 B.n531 B.n30 10.6151
R1348 B.n531 B.n530 10.6151
R1349 B.n530 B.n529 10.6151
R1350 B.n529 B.n32 10.6151
R1351 B.n525 B.n32 10.6151
R1352 B.n525 B.n524 10.6151
R1353 B.n524 B.n523 10.6151
R1354 B.n523 B.n34 10.6151
R1355 B.n519 B.n34 10.6151
R1356 B.n519 B.n518 10.6151
R1357 B.n518 B.n517 10.6151
R1358 B.n517 B.n36 10.6151
R1359 B.n513 B.n36 10.6151
R1360 B.n513 B.n512 10.6151
R1361 B.n510 B.n40 10.6151
R1362 B.n506 B.n40 10.6151
R1363 B.n506 B.n505 10.6151
R1364 B.n505 B.n504 10.6151
R1365 B.n504 B.n42 10.6151
R1366 B.n500 B.n42 10.6151
R1367 B.n500 B.n499 10.6151
R1368 B.n499 B.n498 10.6151
R1369 B.n495 B.n494 10.6151
R1370 B.n494 B.n493 10.6151
R1371 B.n493 B.n48 10.6151
R1372 B.n489 B.n48 10.6151
R1373 B.n489 B.n488 10.6151
R1374 B.n488 B.n487 10.6151
R1375 B.n487 B.n50 10.6151
R1376 B.n483 B.n50 10.6151
R1377 B.n483 B.n482 10.6151
R1378 B.n482 B.n481 10.6151
R1379 B.n481 B.n52 10.6151
R1380 B.n477 B.n52 10.6151
R1381 B.n477 B.n476 10.6151
R1382 B.n476 B.n475 10.6151
R1383 B.n475 B.n54 10.6151
R1384 B.n471 B.n54 10.6151
R1385 B.n471 B.n470 10.6151
R1386 B.n470 B.n469 10.6151
R1387 B.n469 B.n56 10.6151
R1388 B.n465 B.n56 10.6151
R1389 B.n465 B.n464 10.6151
R1390 B.n464 B.n463 10.6151
R1391 B.n463 B.n58 10.6151
R1392 B.n459 B.n58 10.6151
R1393 B.n459 B.n458 10.6151
R1394 B.n458 B.n457 10.6151
R1395 B.n457 B.n60 10.6151
R1396 B.n453 B.n60 10.6151
R1397 B.n453 B.n452 10.6151
R1398 B.n452 B.n451 10.6151
R1399 B.n451 B.n62 10.6151
R1400 B.n332 B.n331 10.6151
R1401 B.n333 B.n332 10.6151
R1402 B.n333 B.n100 10.6151
R1403 B.n337 B.n100 10.6151
R1404 B.n338 B.n337 10.6151
R1405 B.n339 B.n338 10.6151
R1406 B.n339 B.n98 10.6151
R1407 B.n343 B.n98 10.6151
R1408 B.n344 B.n343 10.6151
R1409 B.n345 B.n344 10.6151
R1410 B.n345 B.n96 10.6151
R1411 B.n349 B.n96 10.6151
R1412 B.n350 B.n349 10.6151
R1413 B.n351 B.n350 10.6151
R1414 B.n351 B.n94 10.6151
R1415 B.n355 B.n94 10.6151
R1416 B.n356 B.n355 10.6151
R1417 B.n357 B.n356 10.6151
R1418 B.n357 B.n92 10.6151
R1419 B.n361 B.n92 10.6151
R1420 B.n362 B.n361 10.6151
R1421 B.n363 B.n362 10.6151
R1422 B.n363 B.n90 10.6151
R1423 B.n367 B.n90 10.6151
R1424 B.n368 B.n367 10.6151
R1425 B.n369 B.n368 10.6151
R1426 B.n369 B.n88 10.6151
R1427 B.n373 B.n88 10.6151
R1428 B.n374 B.n373 10.6151
R1429 B.n375 B.n374 10.6151
R1430 B.n375 B.n86 10.6151
R1431 B.n379 B.n86 10.6151
R1432 B.n380 B.n379 10.6151
R1433 B.n381 B.n380 10.6151
R1434 B.n381 B.n84 10.6151
R1435 B.n385 B.n84 10.6151
R1436 B.n386 B.n385 10.6151
R1437 B.n387 B.n386 10.6151
R1438 B.n387 B.n82 10.6151
R1439 B.n391 B.n82 10.6151
R1440 B.n392 B.n391 10.6151
R1441 B.n393 B.n392 10.6151
R1442 B.n393 B.n80 10.6151
R1443 B.n397 B.n80 10.6151
R1444 B.n398 B.n397 10.6151
R1445 B.n399 B.n398 10.6151
R1446 B.n399 B.n78 10.6151
R1447 B.n403 B.n78 10.6151
R1448 B.n404 B.n403 10.6151
R1449 B.n405 B.n404 10.6151
R1450 B.n405 B.n76 10.6151
R1451 B.n409 B.n76 10.6151
R1452 B.n410 B.n409 10.6151
R1453 B.n411 B.n410 10.6151
R1454 B.n411 B.n74 10.6151
R1455 B.n415 B.n74 10.6151
R1456 B.n416 B.n415 10.6151
R1457 B.n417 B.n416 10.6151
R1458 B.n417 B.n72 10.6151
R1459 B.n421 B.n72 10.6151
R1460 B.n422 B.n421 10.6151
R1461 B.n423 B.n422 10.6151
R1462 B.n423 B.n70 10.6151
R1463 B.n427 B.n70 10.6151
R1464 B.n428 B.n427 10.6151
R1465 B.n429 B.n428 10.6151
R1466 B.n429 B.n68 10.6151
R1467 B.n433 B.n68 10.6151
R1468 B.n434 B.n433 10.6151
R1469 B.n435 B.n434 10.6151
R1470 B.n435 B.n66 10.6151
R1471 B.n439 B.n66 10.6151
R1472 B.n440 B.n439 10.6151
R1473 B.n441 B.n440 10.6151
R1474 B.n441 B.n64 10.6151
R1475 B.n445 B.n64 10.6151
R1476 B.n446 B.n445 10.6151
R1477 B.n447 B.n446 10.6151
R1478 B.n219 B.n142 10.6151
R1479 B.n223 B.n142 10.6151
R1480 B.n224 B.n223 10.6151
R1481 B.n225 B.n224 10.6151
R1482 B.n225 B.n140 10.6151
R1483 B.n229 B.n140 10.6151
R1484 B.n230 B.n229 10.6151
R1485 B.n231 B.n230 10.6151
R1486 B.n231 B.n138 10.6151
R1487 B.n235 B.n138 10.6151
R1488 B.n236 B.n235 10.6151
R1489 B.n237 B.n236 10.6151
R1490 B.n237 B.n136 10.6151
R1491 B.n241 B.n136 10.6151
R1492 B.n242 B.n241 10.6151
R1493 B.n243 B.n242 10.6151
R1494 B.n243 B.n134 10.6151
R1495 B.n247 B.n134 10.6151
R1496 B.n248 B.n247 10.6151
R1497 B.n249 B.n248 10.6151
R1498 B.n249 B.n132 10.6151
R1499 B.n253 B.n132 10.6151
R1500 B.n254 B.n253 10.6151
R1501 B.n255 B.n254 10.6151
R1502 B.n255 B.n130 10.6151
R1503 B.n259 B.n130 10.6151
R1504 B.n260 B.n259 10.6151
R1505 B.n261 B.n260 10.6151
R1506 B.n261 B.n128 10.6151
R1507 B.n265 B.n128 10.6151
R1508 B.n266 B.n265 10.6151
R1509 B.n268 B.n124 10.6151
R1510 B.n272 B.n124 10.6151
R1511 B.n273 B.n272 10.6151
R1512 B.n274 B.n273 10.6151
R1513 B.n274 B.n122 10.6151
R1514 B.n278 B.n122 10.6151
R1515 B.n279 B.n278 10.6151
R1516 B.n280 B.n279 10.6151
R1517 B.n284 B.n283 10.6151
R1518 B.n285 B.n284 10.6151
R1519 B.n285 B.n116 10.6151
R1520 B.n289 B.n116 10.6151
R1521 B.n290 B.n289 10.6151
R1522 B.n291 B.n290 10.6151
R1523 B.n291 B.n114 10.6151
R1524 B.n295 B.n114 10.6151
R1525 B.n296 B.n295 10.6151
R1526 B.n297 B.n296 10.6151
R1527 B.n297 B.n112 10.6151
R1528 B.n301 B.n112 10.6151
R1529 B.n302 B.n301 10.6151
R1530 B.n303 B.n302 10.6151
R1531 B.n303 B.n110 10.6151
R1532 B.n307 B.n110 10.6151
R1533 B.n308 B.n307 10.6151
R1534 B.n309 B.n308 10.6151
R1535 B.n309 B.n108 10.6151
R1536 B.n313 B.n108 10.6151
R1537 B.n314 B.n313 10.6151
R1538 B.n315 B.n314 10.6151
R1539 B.n315 B.n106 10.6151
R1540 B.n319 B.n106 10.6151
R1541 B.n320 B.n319 10.6151
R1542 B.n321 B.n320 10.6151
R1543 B.n321 B.n104 10.6151
R1544 B.n325 B.n104 10.6151
R1545 B.n326 B.n325 10.6151
R1546 B.n327 B.n326 10.6151
R1547 B.n327 B.n102 10.6151
R1548 B.n218 B.n217 10.6151
R1549 B.n217 B.n144 10.6151
R1550 B.n213 B.n144 10.6151
R1551 B.n213 B.n212 10.6151
R1552 B.n212 B.n211 10.6151
R1553 B.n211 B.n146 10.6151
R1554 B.n207 B.n146 10.6151
R1555 B.n207 B.n206 10.6151
R1556 B.n206 B.n205 10.6151
R1557 B.n205 B.n148 10.6151
R1558 B.n201 B.n148 10.6151
R1559 B.n201 B.n200 10.6151
R1560 B.n200 B.n199 10.6151
R1561 B.n199 B.n150 10.6151
R1562 B.n195 B.n150 10.6151
R1563 B.n195 B.n194 10.6151
R1564 B.n194 B.n193 10.6151
R1565 B.n193 B.n152 10.6151
R1566 B.n189 B.n152 10.6151
R1567 B.n189 B.n188 10.6151
R1568 B.n188 B.n187 10.6151
R1569 B.n187 B.n154 10.6151
R1570 B.n183 B.n154 10.6151
R1571 B.n183 B.n182 10.6151
R1572 B.n182 B.n181 10.6151
R1573 B.n181 B.n156 10.6151
R1574 B.n177 B.n156 10.6151
R1575 B.n177 B.n176 10.6151
R1576 B.n176 B.n175 10.6151
R1577 B.n175 B.n158 10.6151
R1578 B.n171 B.n158 10.6151
R1579 B.n171 B.n170 10.6151
R1580 B.n170 B.n169 10.6151
R1581 B.n169 B.n160 10.6151
R1582 B.n165 B.n160 10.6151
R1583 B.n165 B.n164 10.6151
R1584 B.n164 B.n163 10.6151
R1585 B.n163 B.n0 10.6151
R1586 B.n615 B.n1 10.6151
R1587 B.n615 B.n614 10.6151
R1588 B.n614 B.n613 10.6151
R1589 B.n613 B.n4 10.6151
R1590 B.n609 B.n4 10.6151
R1591 B.n609 B.n608 10.6151
R1592 B.n608 B.n607 10.6151
R1593 B.n607 B.n6 10.6151
R1594 B.n603 B.n6 10.6151
R1595 B.n603 B.n602 10.6151
R1596 B.n602 B.n601 10.6151
R1597 B.n601 B.n8 10.6151
R1598 B.n597 B.n8 10.6151
R1599 B.n597 B.n596 10.6151
R1600 B.n596 B.n595 10.6151
R1601 B.n595 B.n10 10.6151
R1602 B.n591 B.n10 10.6151
R1603 B.n591 B.n590 10.6151
R1604 B.n590 B.n589 10.6151
R1605 B.n589 B.n12 10.6151
R1606 B.n585 B.n12 10.6151
R1607 B.n585 B.n584 10.6151
R1608 B.n584 B.n583 10.6151
R1609 B.n583 B.n14 10.6151
R1610 B.n579 B.n14 10.6151
R1611 B.n579 B.n578 10.6151
R1612 B.n578 B.n577 10.6151
R1613 B.n577 B.n16 10.6151
R1614 B.n573 B.n16 10.6151
R1615 B.n573 B.n572 10.6151
R1616 B.n572 B.n571 10.6151
R1617 B.n571 B.n18 10.6151
R1618 B.n567 B.n18 10.6151
R1619 B.n567 B.n566 10.6151
R1620 B.n566 B.n565 10.6151
R1621 B.n565 B.n20 10.6151
R1622 B.n561 B.n20 10.6151
R1623 B.n561 B.n560 10.6151
R1624 B.n511 B.n510 6.5566
R1625 B.n498 B.n46 6.5566
R1626 B.n268 B.n267 6.5566
R1627 B.n280 B.n120 6.5566
R1628 B.n512 B.n511 4.05904
R1629 B.n495 B.n46 4.05904
R1630 B.n267 B.n266 4.05904
R1631 B.n283 B.n120 4.05904
R1632 B.n619 B.n0 2.81026
R1633 B.n619 B.n1 2.81026
C0 B VP 1.72978f
C1 VP w_n3082_n2710# 6.09933f
C2 VP VTAIL 5.11757f
C3 VDD2 B 1.82598f
C4 B VDD1 1.75884f
C5 VDD2 w_n3082_n2710# 2.06572f
C6 VDD1 w_n3082_n2710# 1.98987f
C7 VDD2 VTAIL 6.50165f
C8 VDD1 VTAIL 6.45224f
C9 VDD2 VP 0.433362f
C10 VP VDD1 5.151f
C11 VDD2 VDD1 1.29294f
C12 B VN 1.06732f
C13 w_n3082_n2710# VN 5.70168f
C14 VTAIL VN 5.10332f
C15 VP VN 6.03287f
C16 B w_n3082_n2710# 8.35295f
C17 VDD2 VN 4.87053f
C18 VDD1 VN 0.150243f
C19 B VTAIL 2.85095f
C20 w_n3082_n2710# VTAIL 2.48627f
C21 VDD2 VSUBS 1.618983f
C22 VDD1 VSUBS 1.550346f
C23 VTAIL VSUBS 1.019517f
C24 VN VSUBS 5.448319f
C25 VP VSUBS 2.596189f
C26 B VSUBS 4.069706f
C27 w_n3082_n2710# VSUBS 0.103444p
C28 B.n0 VSUBS 0.00441f
C29 B.n1 VSUBS 0.00441f
C30 B.n2 VSUBS 0.006973f
C31 B.n3 VSUBS 0.006973f
C32 B.n4 VSUBS 0.006973f
C33 B.n5 VSUBS 0.006973f
C34 B.n6 VSUBS 0.006973f
C35 B.n7 VSUBS 0.006973f
C36 B.n8 VSUBS 0.006973f
C37 B.n9 VSUBS 0.006973f
C38 B.n10 VSUBS 0.006973f
C39 B.n11 VSUBS 0.006973f
C40 B.n12 VSUBS 0.006973f
C41 B.n13 VSUBS 0.006973f
C42 B.n14 VSUBS 0.006973f
C43 B.n15 VSUBS 0.006973f
C44 B.n16 VSUBS 0.006973f
C45 B.n17 VSUBS 0.006973f
C46 B.n18 VSUBS 0.006973f
C47 B.n19 VSUBS 0.006973f
C48 B.n20 VSUBS 0.006973f
C49 B.n21 VSUBS 0.017325f
C50 B.n22 VSUBS 0.006973f
C51 B.n23 VSUBS 0.006973f
C52 B.n24 VSUBS 0.006973f
C53 B.n25 VSUBS 0.006973f
C54 B.n26 VSUBS 0.006973f
C55 B.n27 VSUBS 0.006973f
C56 B.n28 VSUBS 0.006973f
C57 B.n29 VSUBS 0.006973f
C58 B.n30 VSUBS 0.006973f
C59 B.n31 VSUBS 0.006973f
C60 B.n32 VSUBS 0.006973f
C61 B.n33 VSUBS 0.006973f
C62 B.n34 VSUBS 0.006973f
C63 B.n35 VSUBS 0.006973f
C64 B.n36 VSUBS 0.006973f
C65 B.n37 VSUBS 0.006973f
C66 B.t5 VSUBS 0.140332f
C67 B.t4 VSUBS 0.166947f
C68 B.t3 VSUBS 0.923488f
C69 B.n38 VSUBS 0.274752f
C70 B.n39 VSUBS 0.201072f
C71 B.n40 VSUBS 0.006973f
C72 B.n41 VSUBS 0.006973f
C73 B.n42 VSUBS 0.006973f
C74 B.n43 VSUBS 0.006973f
C75 B.t2 VSUBS 0.140334f
C76 B.t1 VSUBS 0.166949f
C77 B.t0 VSUBS 0.923488f
C78 B.n44 VSUBS 0.27475f
C79 B.n45 VSUBS 0.20107f
C80 B.n46 VSUBS 0.016157f
C81 B.n47 VSUBS 0.006973f
C82 B.n48 VSUBS 0.006973f
C83 B.n49 VSUBS 0.006973f
C84 B.n50 VSUBS 0.006973f
C85 B.n51 VSUBS 0.006973f
C86 B.n52 VSUBS 0.006973f
C87 B.n53 VSUBS 0.006973f
C88 B.n54 VSUBS 0.006973f
C89 B.n55 VSUBS 0.006973f
C90 B.n56 VSUBS 0.006973f
C91 B.n57 VSUBS 0.006973f
C92 B.n58 VSUBS 0.006973f
C93 B.n59 VSUBS 0.006973f
C94 B.n60 VSUBS 0.006973f
C95 B.n61 VSUBS 0.006973f
C96 B.n62 VSUBS 0.017218f
C97 B.n63 VSUBS 0.006973f
C98 B.n64 VSUBS 0.006973f
C99 B.n65 VSUBS 0.006973f
C100 B.n66 VSUBS 0.006973f
C101 B.n67 VSUBS 0.006973f
C102 B.n68 VSUBS 0.006973f
C103 B.n69 VSUBS 0.006973f
C104 B.n70 VSUBS 0.006973f
C105 B.n71 VSUBS 0.006973f
C106 B.n72 VSUBS 0.006973f
C107 B.n73 VSUBS 0.006973f
C108 B.n74 VSUBS 0.006973f
C109 B.n75 VSUBS 0.006973f
C110 B.n76 VSUBS 0.006973f
C111 B.n77 VSUBS 0.006973f
C112 B.n78 VSUBS 0.006973f
C113 B.n79 VSUBS 0.006973f
C114 B.n80 VSUBS 0.006973f
C115 B.n81 VSUBS 0.006973f
C116 B.n82 VSUBS 0.006973f
C117 B.n83 VSUBS 0.006973f
C118 B.n84 VSUBS 0.006973f
C119 B.n85 VSUBS 0.006973f
C120 B.n86 VSUBS 0.006973f
C121 B.n87 VSUBS 0.006973f
C122 B.n88 VSUBS 0.006973f
C123 B.n89 VSUBS 0.006973f
C124 B.n90 VSUBS 0.006973f
C125 B.n91 VSUBS 0.006973f
C126 B.n92 VSUBS 0.006973f
C127 B.n93 VSUBS 0.006973f
C128 B.n94 VSUBS 0.006973f
C129 B.n95 VSUBS 0.006973f
C130 B.n96 VSUBS 0.006973f
C131 B.n97 VSUBS 0.006973f
C132 B.n98 VSUBS 0.006973f
C133 B.n99 VSUBS 0.006973f
C134 B.n100 VSUBS 0.006973f
C135 B.n101 VSUBS 0.006973f
C136 B.n102 VSUBS 0.017952f
C137 B.n103 VSUBS 0.006973f
C138 B.n104 VSUBS 0.006973f
C139 B.n105 VSUBS 0.006973f
C140 B.n106 VSUBS 0.006973f
C141 B.n107 VSUBS 0.006973f
C142 B.n108 VSUBS 0.006973f
C143 B.n109 VSUBS 0.006973f
C144 B.n110 VSUBS 0.006973f
C145 B.n111 VSUBS 0.006973f
C146 B.n112 VSUBS 0.006973f
C147 B.n113 VSUBS 0.006973f
C148 B.n114 VSUBS 0.006973f
C149 B.n115 VSUBS 0.006973f
C150 B.n116 VSUBS 0.006973f
C151 B.n117 VSUBS 0.006973f
C152 B.t7 VSUBS 0.140334f
C153 B.t8 VSUBS 0.166949f
C154 B.t6 VSUBS 0.923488f
C155 B.n118 VSUBS 0.27475f
C156 B.n119 VSUBS 0.20107f
C157 B.n120 VSUBS 0.016157f
C158 B.n121 VSUBS 0.006973f
C159 B.n122 VSUBS 0.006973f
C160 B.n123 VSUBS 0.006973f
C161 B.n124 VSUBS 0.006973f
C162 B.n125 VSUBS 0.006973f
C163 B.t10 VSUBS 0.140332f
C164 B.t11 VSUBS 0.166947f
C165 B.t9 VSUBS 0.923488f
C166 B.n126 VSUBS 0.274752f
C167 B.n127 VSUBS 0.201072f
C168 B.n128 VSUBS 0.006973f
C169 B.n129 VSUBS 0.006973f
C170 B.n130 VSUBS 0.006973f
C171 B.n131 VSUBS 0.006973f
C172 B.n132 VSUBS 0.006973f
C173 B.n133 VSUBS 0.006973f
C174 B.n134 VSUBS 0.006973f
C175 B.n135 VSUBS 0.006973f
C176 B.n136 VSUBS 0.006973f
C177 B.n137 VSUBS 0.006973f
C178 B.n138 VSUBS 0.006973f
C179 B.n139 VSUBS 0.006973f
C180 B.n140 VSUBS 0.006973f
C181 B.n141 VSUBS 0.006973f
C182 B.n142 VSUBS 0.006973f
C183 B.n143 VSUBS 0.017325f
C184 B.n144 VSUBS 0.006973f
C185 B.n145 VSUBS 0.006973f
C186 B.n146 VSUBS 0.006973f
C187 B.n147 VSUBS 0.006973f
C188 B.n148 VSUBS 0.006973f
C189 B.n149 VSUBS 0.006973f
C190 B.n150 VSUBS 0.006973f
C191 B.n151 VSUBS 0.006973f
C192 B.n152 VSUBS 0.006973f
C193 B.n153 VSUBS 0.006973f
C194 B.n154 VSUBS 0.006973f
C195 B.n155 VSUBS 0.006973f
C196 B.n156 VSUBS 0.006973f
C197 B.n157 VSUBS 0.006973f
C198 B.n158 VSUBS 0.006973f
C199 B.n159 VSUBS 0.006973f
C200 B.n160 VSUBS 0.006973f
C201 B.n161 VSUBS 0.006973f
C202 B.n162 VSUBS 0.006973f
C203 B.n163 VSUBS 0.006973f
C204 B.n164 VSUBS 0.006973f
C205 B.n165 VSUBS 0.006973f
C206 B.n166 VSUBS 0.006973f
C207 B.n167 VSUBS 0.006973f
C208 B.n168 VSUBS 0.006973f
C209 B.n169 VSUBS 0.006973f
C210 B.n170 VSUBS 0.006973f
C211 B.n171 VSUBS 0.006973f
C212 B.n172 VSUBS 0.006973f
C213 B.n173 VSUBS 0.006973f
C214 B.n174 VSUBS 0.006973f
C215 B.n175 VSUBS 0.006973f
C216 B.n176 VSUBS 0.006973f
C217 B.n177 VSUBS 0.006973f
C218 B.n178 VSUBS 0.006973f
C219 B.n179 VSUBS 0.006973f
C220 B.n180 VSUBS 0.006973f
C221 B.n181 VSUBS 0.006973f
C222 B.n182 VSUBS 0.006973f
C223 B.n183 VSUBS 0.006973f
C224 B.n184 VSUBS 0.006973f
C225 B.n185 VSUBS 0.006973f
C226 B.n186 VSUBS 0.006973f
C227 B.n187 VSUBS 0.006973f
C228 B.n188 VSUBS 0.006973f
C229 B.n189 VSUBS 0.006973f
C230 B.n190 VSUBS 0.006973f
C231 B.n191 VSUBS 0.006973f
C232 B.n192 VSUBS 0.006973f
C233 B.n193 VSUBS 0.006973f
C234 B.n194 VSUBS 0.006973f
C235 B.n195 VSUBS 0.006973f
C236 B.n196 VSUBS 0.006973f
C237 B.n197 VSUBS 0.006973f
C238 B.n198 VSUBS 0.006973f
C239 B.n199 VSUBS 0.006973f
C240 B.n200 VSUBS 0.006973f
C241 B.n201 VSUBS 0.006973f
C242 B.n202 VSUBS 0.006973f
C243 B.n203 VSUBS 0.006973f
C244 B.n204 VSUBS 0.006973f
C245 B.n205 VSUBS 0.006973f
C246 B.n206 VSUBS 0.006973f
C247 B.n207 VSUBS 0.006973f
C248 B.n208 VSUBS 0.006973f
C249 B.n209 VSUBS 0.006973f
C250 B.n210 VSUBS 0.006973f
C251 B.n211 VSUBS 0.006973f
C252 B.n212 VSUBS 0.006973f
C253 B.n213 VSUBS 0.006973f
C254 B.n214 VSUBS 0.006973f
C255 B.n215 VSUBS 0.006973f
C256 B.n216 VSUBS 0.006973f
C257 B.n217 VSUBS 0.006973f
C258 B.n218 VSUBS 0.017325f
C259 B.n219 VSUBS 0.017952f
C260 B.n220 VSUBS 0.017952f
C261 B.n221 VSUBS 0.006973f
C262 B.n222 VSUBS 0.006973f
C263 B.n223 VSUBS 0.006973f
C264 B.n224 VSUBS 0.006973f
C265 B.n225 VSUBS 0.006973f
C266 B.n226 VSUBS 0.006973f
C267 B.n227 VSUBS 0.006973f
C268 B.n228 VSUBS 0.006973f
C269 B.n229 VSUBS 0.006973f
C270 B.n230 VSUBS 0.006973f
C271 B.n231 VSUBS 0.006973f
C272 B.n232 VSUBS 0.006973f
C273 B.n233 VSUBS 0.006973f
C274 B.n234 VSUBS 0.006973f
C275 B.n235 VSUBS 0.006973f
C276 B.n236 VSUBS 0.006973f
C277 B.n237 VSUBS 0.006973f
C278 B.n238 VSUBS 0.006973f
C279 B.n239 VSUBS 0.006973f
C280 B.n240 VSUBS 0.006973f
C281 B.n241 VSUBS 0.006973f
C282 B.n242 VSUBS 0.006973f
C283 B.n243 VSUBS 0.006973f
C284 B.n244 VSUBS 0.006973f
C285 B.n245 VSUBS 0.006973f
C286 B.n246 VSUBS 0.006973f
C287 B.n247 VSUBS 0.006973f
C288 B.n248 VSUBS 0.006973f
C289 B.n249 VSUBS 0.006973f
C290 B.n250 VSUBS 0.006973f
C291 B.n251 VSUBS 0.006973f
C292 B.n252 VSUBS 0.006973f
C293 B.n253 VSUBS 0.006973f
C294 B.n254 VSUBS 0.006973f
C295 B.n255 VSUBS 0.006973f
C296 B.n256 VSUBS 0.006973f
C297 B.n257 VSUBS 0.006973f
C298 B.n258 VSUBS 0.006973f
C299 B.n259 VSUBS 0.006973f
C300 B.n260 VSUBS 0.006973f
C301 B.n261 VSUBS 0.006973f
C302 B.n262 VSUBS 0.006973f
C303 B.n263 VSUBS 0.006973f
C304 B.n264 VSUBS 0.006973f
C305 B.n265 VSUBS 0.006973f
C306 B.n266 VSUBS 0.00482f
C307 B.n267 VSUBS 0.016157f
C308 B.n268 VSUBS 0.00564f
C309 B.n269 VSUBS 0.006973f
C310 B.n270 VSUBS 0.006973f
C311 B.n271 VSUBS 0.006973f
C312 B.n272 VSUBS 0.006973f
C313 B.n273 VSUBS 0.006973f
C314 B.n274 VSUBS 0.006973f
C315 B.n275 VSUBS 0.006973f
C316 B.n276 VSUBS 0.006973f
C317 B.n277 VSUBS 0.006973f
C318 B.n278 VSUBS 0.006973f
C319 B.n279 VSUBS 0.006973f
C320 B.n280 VSUBS 0.00564f
C321 B.n281 VSUBS 0.006973f
C322 B.n282 VSUBS 0.006973f
C323 B.n283 VSUBS 0.00482f
C324 B.n284 VSUBS 0.006973f
C325 B.n285 VSUBS 0.006973f
C326 B.n286 VSUBS 0.006973f
C327 B.n287 VSUBS 0.006973f
C328 B.n288 VSUBS 0.006973f
C329 B.n289 VSUBS 0.006973f
C330 B.n290 VSUBS 0.006973f
C331 B.n291 VSUBS 0.006973f
C332 B.n292 VSUBS 0.006973f
C333 B.n293 VSUBS 0.006973f
C334 B.n294 VSUBS 0.006973f
C335 B.n295 VSUBS 0.006973f
C336 B.n296 VSUBS 0.006973f
C337 B.n297 VSUBS 0.006973f
C338 B.n298 VSUBS 0.006973f
C339 B.n299 VSUBS 0.006973f
C340 B.n300 VSUBS 0.006973f
C341 B.n301 VSUBS 0.006973f
C342 B.n302 VSUBS 0.006973f
C343 B.n303 VSUBS 0.006973f
C344 B.n304 VSUBS 0.006973f
C345 B.n305 VSUBS 0.006973f
C346 B.n306 VSUBS 0.006973f
C347 B.n307 VSUBS 0.006973f
C348 B.n308 VSUBS 0.006973f
C349 B.n309 VSUBS 0.006973f
C350 B.n310 VSUBS 0.006973f
C351 B.n311 VSUBS 0.006973f
C352 B.n312 VSUBS 0.006973f
C353 B.n313 VSUBS 0.006973f
C354 B.n314 VSUBS 0.006973f
C355 B.n315 VSUBS 0.006973f
C356 B.n316 VSUBS 0.006973f
C357 B.n317 VSUBS 0.006973f
C358 B.n318 VSUBS 0.006973f
C359 B.n319 VSUBS 0.006973f
C360 B.n320 VSUBS 0.006973f
C361 B.n321 VSUBS 0.006973f
C362 B.n322 VSUBS 0.006973f
C363 B.n323 VSUBS 0.006973f
C364 B.n324 VSUBS 0.006973f
C365 B.n325 VSUBS 0.006973f
C366 B.n326 VSUBS 0.006973f
C367 B.n327 VSUBS 0.006973f
C368 B.n328 VSUBS 0.006973f
C369 B.n329 VSUBS 0.017952f
C370 B.n330 VSUBS 0.017325f
C371 B.n331 VSUBS 0.017325f
C372 B.n332 VSUBS 0.006973f
C373 B.n333 VSUBS 0.006973f
C374 B.n334 VSUBS 0.006973f
C375 B.n335 VSUBS 0.006973f
C376 B.n336 VSUBS 0.006973f
C377 B.n337 VSUBS 0.006973f
C378 B.n338 VSUBS 0.006973f
C379 B.n339 VSUBS 0.006973f
C380 B.n340 VSUBS 0.006973f
C381 B.n341 VSUBS 0.006973f
C382 B.n342 VSUBS 0.006973f
C383 B.n343 VSUBS 0.006973f
C384 B.n344 VSUBS 0.006973f
C385 B.n345 VSUBS 0.006973f
C386 B.n346 VSUBS 0.006973f
C387 B.n347 VSUBS 0.006973f
C388 B.n348 VSUBS 0.006973f
C389 B.n349 VSUBS 0.006973f
C390 B.n350 VSUBS 0.006973f
C391 B.n351 VSUBS 0.006973f
C392 B.n352 VSUBS 0.006973f
C393 B.n353 VSUBS 0.006973f
C394 B.n354 VSUBS 0.006973f
C395 B.n355 VSUBS 0.006973f
C396 B.n356 VSUBS 0.006973f
C397 B.n357 VSUBS 0.006973f
C398 B.n358 VSUBS 0.006973f
C399 B.n359 VSUBS 0.006973f
C400 B.n360 VSUBS 0.006973f
C401 B.n361 VSUBS 0.006973f
C402 B.n362 VSUBS 0.006973f
C403 B.n363 VSUBS 0.006973f
C404 B.n364 VSUBS 0.006973f
C405 B.n365 VSUBS 0.006973f
C406 B.n366 VSUBS 0.006973f
C407 B.n367 VSUBS 0.006973f
C408 B.n368 VSUBS 0.006973f
C409 B.n369 VSUBS 0.006973f
C410 B.n370 VSUBS 0.006973f
C411 B.n371 VSUBS 0.006973f
C412 B.n372 VSUBS 0.006973f
C413 B.n373 VSUBS 0.006973f
C414 B.n374 VSUBS 0.006973f
C415 B.n375 VSUBS 0.006973f
C416 B.n376 VSUBS 0.006973f
C417 B.n377 VSUBS 0.006973f
C418 B.n378 VSUBS 0.006973f
C419 B.n379 VSUBS 0.006973f
C420 B.n380 VSUBS 0.006973f
C421 B.n381 VSUBS 0.006973f
C422 B.n382 VSUBS 0.006973f
C423 B.n383 VSUBS 0.006973f
C424 B.n384 VSUBS 0.006973f
C425 B.n385 VSUBS 0.006973f
C426 B.n386 VSUBS 0.006973f
C427 B.n387 VSUBS 0.006973f
C428 B.n388 VSUBS 0.006973f
C429 B.n389 VSUBS 0.006973f
C430 B.n390 VSUBS 0.006973f
C431 B.n391 VSUBS 0.006973f
C432 B.n392 VSUBS 0.006973f
C433 B.n393 VSUBS 0.006973f
C434 B.n394 VSUBS 0.006973f
C435 B.n395 VSUBS 0.006973f
C436 B.n396 VSUBS 0.006973f
C437 B.n397 VSUBS 0.006973f
C438 B.n398 VSUBS 0.006973f
C439 B.n399 VSUBS 0.006973f
C440 B.n400 VSUBS 0.006973f
C441 B.n401 VSUBS 0.006973f
C442 B.n402 VSUBS 0.006973f
C443 B.n403 VSUBS 0.006973f
C444 B.n404 VSUBS 0.006973f
C445 B.n405 VSUBS 0.006973f
C446 B.n406 VSUBS 0.006973f
C447 B.n407 VSUBS 0.006973f
C448 B.n408 VSUBS 0.006973f
C449 B.n409 VSUBS 0.006973f
C450 B.n410 VSUBS 0.006973f
C451 B.n411 VSUBS 0.006973f
C452 B.n412 VSUBS 0.006973f
C453 B.n413 VSUBS 0.006973f
C454 B.n414 VSUBS 0.006973f
C455 B.n415 VSUBS 0.006973f
C456 B.n416 VSUBS 0.006973f
C457 B.n417 VSUBS 0.006973f
C458 B.n418 VSUBS 0.006973f
C459 B.n419 VSUBS 0.006973f
C460 B.n420 VSUBS 0.006973f
C461 B.n421 VSUBS 0.006973f
C462 B.n422 VSUBS 0.006973f
C463 B.n423 VSUBS 0.006973f
C464 B.n424 VSUBS 0.006973f
C465 B.n425 VSUBS 0.006973f
C466 B.n426 VSUBS 0.006973f
C467 B.n427 VSUBS 0.006973f
C468 B.n428 VSUBS 0.006973f
C469 B.n429 VSUBS 0.006973f
C470 B.n430 VSUBS 0.006973f
C471 B.n431 VSUBS 0.006973f
C472 B.n432 VSUBS 0.006973f
C473 B.n433 VSUBS 0.006973f
C474 B.n434 VSUBS 0.006973f
C475 B.n435 VSUBS 0.006973f
C476 B.n436 VSUBS 0.006973f
C477 B.n437 VSUBS 0.006973f
C478 B.n438 VSUBS 0.006973f
C479 B.n439 VSUBS 0.006973f
C480 B.n440 VSUBS 0.006973f
C481 B.n441 VSUBS 0.006973f
C482 B.n442 VSUBS 0.006973f
C483 B.n443 VSUBS 0.006973f
C484 B.n444 VSUBS 0.006973f
C485 B.n445 VSUBS 0.006973f
C486 B.n446 VSUBS 0.006973f
C487 B.n447 VSUBS 0.018059f
C488 B.n448 VSUBS 0.017325f
C489 B.n449 VSUBS 0.017952f
C490 B.n450 VSUBS 0.006973f
C491 B.n451 VSUBS 0.006973f
C492 B.n452 VSUBS 0.006973f
C493 B.n453 VSUBS 0.006973f
C494 B.n454 VSUBS 0.006973f
C495 B.n455 VSUBS 0.006973f
C496 B.n456 VSUBS 0.006973f
C497 B.n457 VSUBS 0.006973f
C498 B.n458 VSUBS 0.006973f
C499 B.n459 VSUBS 0.006973f
C500 B.n460 VSUBS 0.006973f
C501 B.n461 VSUBS 0.006973f
C502 B.n462 VSUBS 0.006973f
C503 B.n463 VSUBS 0.006973f
C504 B.n464 VSUBS 0.006973f
C505 B.n465 VSUBS 0.006973f
C506 B.n466 VSUBS 0.006973f
C507 B.n467 VSUBS 0.006973f
C508 B.n468 VSUBS 0.006973f
C509 B.n469 VSUBS 0.006973f
C510 B.n470 VSUBS 0.006973f
C511 B.n471 VSUBS 0.006973f
C512 B.n472 VSUBS 0.006973f
C513 B.n473 VSUBS 0.006973f
C514 B.n474 VSUBS 0.006973f
C515 B.n475 VSUBS 0.006973f
C516 B.n476 VSUBS 0.006973f
C517 B.n477 VSUBS 0.006973f
C518 B.n478 VSUBS 0.006973f
C519 B.n479 VSUBS 0.006973f
C520 B.n480 VSUBS 0.006973f
C521 B.n481 VSUBS 0.006973f
C522 B.n482 VSUBS 0.006973f
C523 B.n483 VSUBS 0.006973f
C524 B.n484 VSUBS 0.006973f
C525 B.n485 VSUBS 0.006973f
C526 B.n486 VSUBS 0.006973f
C527 B.n487 VSUBS 0.006973f
C528 B.n488 VSUBS 0.006973f
C529 B.n489 VSUBS 0.006973f
C530 B.n490 VSUBS 0.006973f
C531 B.n491 VSUBS 0.006973f
C532 B.n492 VSUBS 0.006973f
C533 B.n493 VSUBS 0.006973f
C534 B.n494 VSUBS 0.006973f
C535 B.n495 VSUBS 0.00482f
C536 B.n496 VSUBS 0.006973f
C537 B.n497 VSUBS 0.006973f
C538 B.n498 VSUBS 0.00564f
C539 B.n499 VSUBS 0.006973f
C540 B.n500 VSUBS 0.006973f
C541 B.n501 VSUBS 0.006973f
C542 B.n502 VSUBS 0.006973f
C543 B.n503 VSUBS 0.006973f
C544 B.n504 VSUBS 0.006973f
C545 B.n505 VSUBS 0.006973f
C546 B.n506 VSUBS 0.006973f
C547 B.n507 VSUBS 0.006973f
C548 B.n508 VSUBS 0.006973f
C549 B.n509 VSUBS 0.006973f
C550 B.n510 VSUBS 0.00564f
C551 B.n511 VSUBS 0.016157f
C552 B.n512 VSUBS 0.00482f
C553 B.n513 VSUBS 0.006973f
C554 B.n514 VSUBS 0.006973f
C555 B.n515 VSUBS 0.006973f
C556 B.n516 VSUBS 0.006973f
C557 B.n517 VSUBS 0.006973f
C558 B.n518 VSUBS 0.006973f
C559 B.n519 VSUBS 0.006973f
C560 B.n520 VSUBS 0.006973f
C561 B.n521 VSUBS 0.006973f
C562 B.n522 VSUBS 0.006973f
C563 B.n523 VSUBS 0.006973f
C564 B.n524 VSUBS 0.006973f
C565 B.n525 VSUBS 0.006973f
C566 B.n526 VSUBS 0.006973f
C567 B.n527 VSUBS 0.006973f
C568 B.n528 VSUBS 0.006973f
C569 B.n529 VSUBS 0.006973f
C570 B.n530 VSUBS 0.006973f
C571 B.n531 VSUBS 0.006973f
C572 B.n532 VSUBS 0.006973f
C573 B.n533 VSUBS 0.006973f
C574 B.n534 VSUBS 0.006973f
C575 B.n535 VSUBS 0.006973f
C576 B.n536 VSUBS 0.006973f
C577 B.n537 VSUBS 0.006973f
C578 B.n538 VSUBS 0.006973f
C579 B.n539 VSUBS 0.006973f
C580 B.n540 VSUBS 0.006973f
C581 B.n541 VSUBS 0.006973f
C582 B.n542 VSUBS 0.006973f
C583 B.n543 VSUBS 0.006973f
C584 B.n544 VSUBS 0.006973f
C585 B.n545 VSUBS 0.006973f
C586 B.n546 VSUBS 0.006973f
C587 B.n547 VSUBS 0.006973f
C588 B.n548 VSUBS 0.006973f
C589 B.n549 VSUBS 0.006973f
C590 B.n550 VSUBS 0.006973f
C591 B.n551 VSUBS 0.006973f
C592 B.n552 VSUBS 0.006973f
C593 B.n553 VSUBS 0.006973f
C594 B.n554 VSUBS 0.006973f
C595 B.n555 VSUBS 0.006973f
C596 B.n556 VSUBS 0.006973f
C597 B.n557 VSUBS 0.006973f
C598 B.n558 VSUBS 0.017952f
C599 B.n559 VSUBS 0.017952f
C600 B.n560 VSUBS 0.017325f
C601 B.n561 VSUBS 0.006973f
C602 B.n562 VSUBS 0.006973f
C603 B.n563 VSUBS 0.006973f
C604 B.n564 VSUBS 0.006973f
C605 B.n565 VSUBS 0.006973f
C606 B.n566 VSUBS 0.006973f
C607 B.n567 VSUBS 0.006973f
C608 B.n568 VSUBS 0.006973f
C609 B.n569 VSUBS 0.006973f
C610 B.n570 VSUBS 0.006973f
C611 B.n571 VSUBS 0.006973f
C612 B.n572 VSUBS 0.006973f
C613 B.n573 VSUBS 0.006973f
C614 B.n574 VSUBS 0.006973f
C615 B.n575 VSUBS 0.006973f
C616 B.n576 VSUBS 0.006973f
C617 B.n577 VSUBS 0.006973f
C618 B.n578 VSUBS 0.006973f
C619 B.n579 VSUBS 0.006973f
C620 B.n580 VSUBS 0.006973f
C621 B.n581 VSUBS 0.006973f
C622 B.n582 VSUBS 0.006973f
C623 B.n583 VSUBS 0.006973f
C624 B.n584 VSUBS 0.006973f
C625 B.n585 VSUBS 0.006973f
C626 B.n586 VSUBS 0.006973f
C627 B.n587 VSUBS 0.006973f
C628 B.n588 VSUBS 0.006973f
C629 B.n589 VSUBS 0.006973f
C630 B.n590 VSUBS 0.006973f
C631 B.n591 VSUBS 0.006973f
C632 B.n592 VSUBS 0.006973f
C633 B.n593 VSUBS 0.006973f
C634 B.n594 VSUBS 0.006973f
C635 B.n595 VSUBS 0.006973f
C636 B.n596 VSUBS 0.006973f
C637 B.n597 VSUBS 0.006973f
C638 B.n598 VSUBS 0.006973f
C639 B.n599 VSUBS 0.006973f
C640 B.n600 VSUBS 0.006973f
C641 B.n601 VSUBS 0.006973f
C642 B.n602 VSUBS 0.006973f
C643 B.n603 VSUBS 0.006973f
C644 B.n604 VSUBS 0.006973f
C645 B.n605 VSUBS 0.006973f
C646 B.n606 VSUBS 0.006973f
C647 B.n607 VSUBS 0.006973f
C648 B.n608 VSUBS 0.006973f
C649 B.n609 VSUBS 0.006973f
C650 B.n610 VSUBS 0.006973f
C651 B.n611 VSUBS 0.006973f
C652 B.n612 VSUBS 0.006973f
C653 B.n613 VSUBS 0.006973f
C654 B.n614 VSUBS 0.006973f
C655 B.n615 VSUBS 0.006973f
C656 B.n616 VSUBS 0.006973f
C657 B.n617 VSUBS 0.006973f
C658 B.n618 VSUBS 0.006973f
C659 B.n619 VSUBS 0.01579f
C660 VDD2.n0 VSUBS 0.027976f
C661 VDD2.n1 VSUBS 0.025658f
C662 VDD2.n2 VSUBS 0.013787f
C663 VDD2.n3 VSUBS 0.032588f
C664 VDD2.n4 VSUBS 0.014598f
C665 VDD2.n5 VSUBS 0.025658f
C666 VDD2.n6 VSUBS 0.013787f
C667 VDD2.n7 VSUBS 0.032588f
C668 VDD2.n8 VSUBS 0.014598f
C669 VDD2.n9 VSUBS 0.025658f
C670 VDD2.n10 VSUBS 0.013787f
C671 VDD2.n11 VSUBS 0.032588f
C672 VDD2.n12 VSUBS 0.014598f
C673 VDD2.n13 VSUBS 0.163971f
C674 VDD2.t5 VSUBS 0.070021f
C675 VDD2.n14 VSUBS 0.024441f
C676 VDD2.n15 VSUBS 0.024515f
C677 VDD2.n16 VSUBS 0.013787f
C678 VDD2.n17 VSUBS 0.890628f
C679 VDD2.n18 VSUBS 0.025658f
C680 VDD2.n19 VSUBS 0.013787f
C681 VDD2.n20 VSUBS 0.014598f
C682 VDD2.n21 VSUBS 0.032588f
C683 VDD2.n22 VSUBS 0.032588f
C684 VDD2.n23 VSUBS 0.014598f
C685 VDD2.n24 VSUBS 0.013787f
C686 VDD2.n25 VSUBS 0.025658f
C687 VDD2.n26 VSUBS 0.025658f
C688 VDD2.n27 VSUBS 0.013787f
C689 VDD2.n28 VSUBS 0.014598f
C690 VDD2.n29 VSUBS 0.032588f
C691 VDD2.n30 VSUBS 0.032588f
C692 VDD2.n31 VSUBS 0.032588f
C693 VDD2.n32 VSUBS 0.014598f
C694 VDD2.n33 VSUBS 0.013787f
C695 VDD2.n34 VSUBS 0.025658f
C696 VDD2.n35 VSUBS 0.025658f
C697 VDD2.n36 VSUBS 0.013787f
C698 VDD2.n37 VSUBS 0.014193f
C699 VDD2.n38 VSUBS 0.014193f
C700 VDD2.n39 VSUBS 0.032588f
C701 VDD2.n40 VSUBS 0.078157f
C702 VDD2.n41 VSUBS 0.014598f
C703 VDD2.n42 VSUBS 0.013787f
C704 VDD2.n43 VSUBS 0.065967f
C705 VDD2.n44 VSUBS 0.06293f
C706 VDD2.t1 VSUBS 0.1766f
C707 VDD2.t4 VSUBS 0.1766f
C708 VDD2.n45 VSUBS 1.3101f
C709 VDD2.n46 VSUBS 2.64614f
C710 VDD2.n47 VSUBS 0.027976f
C711 VDD2.n48 VSUBS 0.025658f
C712 VDD2.n49 VSUBS 0.013787f
C713 VDD2.n50 VSUBS 0.032588f
C714 VDD2.n51 VSUBS 0.014598f
C715 VDD2.n52 VSUBS 0.025658f
C716 VDD2.n53 VSUBS 0.013787f
C717 VDD2.n54 VSUBS 0.032588f
C718 VDD2.n55 VSUBS 0.032588f
C719 VDD2.n56 VSUBS 0.014598f
C720 VDD2.n57 VSUBS 0.025658f
C721 VDD2.n58 VSUBS 0.013787f
C722 VDD2.n59 VSUBS 0.032588f
C723 VDD2.n60 VSUBS 0.014598f
C724 VDD2.n61 VSUBS 0.163971f
C725 VDD2.t3 VSUBS 0.070021f
C726 VDD2.n62 VSUBS 0.024441f
C727 VDD2.n63 VSUBS 0.024515f
C728 VDD2.n64 VSUBS 0.013787f
C729 VDD2.n65 VSUBS 0.890628f
C730 VDD2.n66 VSUBS 0.025658f
C731 VDD2.n67 VSUBS 0.013787f
C732 VDD2.n68 VSUBS 0.014598f
C733 VDD2.n69 VSUBS 0.032588f
C734 VDD2.n70 VSUBS 0.032588f
C735 VDD2.n71 VSUBS 0.014598f
C736 VDD2.n72 VSUBS 0.013787f
C737 VDD2.n73 VSUBS 0.025658f
C738 VDD2.n74 VSUBS 0.025658f
C739 VDD2.n75 VSUBS 0.013787f
C740 VDD2.n76 VSUBS 0.014598f
C741 VDD2.n77 VSUBS 0.032588f
C742 VDD2.n78 VSUBS 0.032588f
C743 VDD2.n79 VSUBS 0.014598f
C744 VDD2.n80 VSUBS 0.013787f
C745 VDD2.n81 VSUBS 0.025658f
C746 VDD2.n82 VSUBS 0.025658f
C747 VDD2.n83 VSUBS 0.013787f
C748 VDD2.n84 VSUBS 0.014193f
C749 VDD2.n85 VSUBS 0.014193f
C750 VDD2.n86 VSUBS 0.032588f
C751 VDD2.n87 VSUBS 0.078157f
C752 VDD2.n88 VSUBS 0.014598f
C753 VDD2.n89 VSUBS 0.013787f
C754 VDD2.n90 VSUBS 0.065967f
C755 VDD2.n91 VSUBS 0.057137f
C756 VDD2.n92 VSUBS 2.28819f
C757 VDD2.t0 VSUBS 0.1766f
C758 VDD2.t2 VSUBS 0.1766f
C759 VDD2.n93 VSUBS 1.31007f
C760 VN.n0 VSUBS 0.046707f
C761 VN.t1 VSUBS 1.92114f
C762 VN.n1 VSUBS 0.030934f
C763 VN.n2 VSUBS 0.305063f
C764 VN.t4 VSUBS 1.92114f
C765 VN.t0 VSUBS 2.16552f
C766 VN.n3 VSUBS 0.77436f
C767 VN.n4 VSUBS 0.792562f
C768 VN.n5 VSUBS 0.049728f
C769 VN.n6 VSUBS 0.07156f
C770 VN.n7 VSUBS 0.035427f
C771 VN.n8 VSUBS 0.035427f
C772 VN.n9 VSUBS 0.035427f
C773 VN.n10 VSUBS 0.066968f
C774 VN.n11 VSUBS 0.058856f
C775 VN.n12 VSUBS 0.822081f
C776 VN.n13 VSUBS 0.045638f
C777 VN.n14 VSUBS 0.046707f
C778 VN.t2 VSUBS 1.92114f
C779 VN.n15 VSUBS 0.030934f
C780 VN.n16 VSUBS 0.305063f
C781 VN.t5 VSUBS 1.92114f
C782 VN.t3 VSUBS 2.16552f
C783 VN.n17 VSUBS 0.77436f
C784 VN.n18 VSUBS 0.792562f
C785 VN.n19 VSUBS 0.049728f
C786 VN.n20 VSUBS 0.07156f
C787 VN.n21 VSUBS 0.035427f
C788 VN.n22 VSUBS 0.035427f
C789 VN.n23 VSUBS 0.035427f
C790 VN.n24 VSUBS 0.066968f
C791 VN.n25 VSUBS 0.058856f
C792 VN.n26 VSUBS 0.822081f
C793 VN.n27 VSUBS 1.69744f
C794 VDD1.n0 VSUBS 0.024077f
C795 VDD1.n1 VSUBS 0.022082f
C796 VDD1.n2 VSUBS 0.011866f
C797 VDD1.n3 VSUBS 0.028046f
C798 VDD1.n4 VSUBS 0.012564f
C799 VDD1.n5 VSUBS 0.022082f
C800 VDD1.n6 VSUBS 0.011866f
C801 VDD1.n7 VSUBS 0.028046f
C802 VDD1.n8 VSUBS 0.028046f
C803 VDD1.n9 VSUBS 0.012564f
C804 VDD1.n10 VSUBS 0.022082f
C805 VDD1.n11 VSUBS 0.011866f
C806 VDD1.n12 VSUBS 0.028046f
C807 VDD1.n13 VSUBS 0.012564f
C808 VDD1.n14 VSUBS 0.141117f
C809 VDD1.t4 VSUBS 0.060262f
C810 VDD1.n15 VSUBS 0.021035f
C811 VDD1.n16 VSUBS 0.021098f
C812 VDD1.n17 VSUBS 0.011866f
C813 VDD1.n18 VSUBS 0.766497f
C814 VDD1.n19 VSUBS 0.022082f
C815 VDD1.n20 VSUBS 0.011866f
C816 VDD1.n21 VSUBS 0.012564f
C817 VDD1.n22 VSUBS 0.028046f
C818 VDD1.n23 VSUBS 0.028046f
C819 VDD1.n24 VSUBS 0.012564f
C820 VDD1.n25 VSUBS 0.011866f
C821 VDD1.n26 VSUBS 0.022082f
C822 VDD1.n27 VSUBS 0.022082f
C823 VDD1.n28 VSUBS 0.011866f
C824 VDD1.n29 VSUBS 0.012564f
C825 VDD1.n30 VSUBS 0.028046f
C826 VDD1.n31 VSUBS 0.028046f
C827 VDD1.n32 VSUBS 0.012564f
C828 VDD1.n33 VSUBS 0.011866f
C829 VDD1.n34 VSUBS 0.022082f
C830 VDD1.n35 VSUBS 0.022082f
C831 VDD1.n36 VSUBS 0.011866f
C832 VDD1.n37 VSUBS 0.012215f
C833 VDD1.n38 VSUBS 0.012215f
C834 VDD1.n39 VSUBS 0.028046f
C835 VDD1.n40 VSUBS 0.067264f
C836 VDD1.n41 VSUBS 0.012564f
C837 VDD1.n42 VSUBS 0.011866f
C838 VDD1.n43 VSUBS 0.056772f
C839 VDD1.n44 VSUBS 0.054743f
C840 VDD1.n45 VSUBS 0.024077f
C841 VDD1.n46 VSUBS 0.022082f
C842 VDD1.n47 VSUBS 0.011866f
C843 VDD1.n48 VSUBS 0.028046f
C844 VDD1.n49 VSUBS 0.012564f
C845 VDD1.n50 VSUBS 0.022082f
C846 VDD1.n51 VSUBS 0.011866f
C847 VDD1.n52 VSUBS 0.028046f
C848 VDD1.n53 VSUBS 0.012564f
C849 VDD1.n54 VSUBS 0.022082f
C850 VDD1.n55 VSUBS 0.011866f
C851 VDD1.n56 VSUBS 0.028046f
C852 VDD1.n57 VSUBS 0.012564f
C853 VDD1.n58 VSUBS 0.141117f
C854 VDD1.t0 VSUBS 0.060262f
C855 VDD1.n59 VSUBS 0.021035f
C856 VDD1.n60 VSUBS 0.021098f
C857 VDD1.n61 VSUBS 0.011866f
C858 VDD1.n62 VSUBS 0.766497f
C859 VDD1.n63 VSUBS 0.022082f
C860 VDD1.n64 VSUBS 0.011866f
C861 VDD1.n65 VSUBS 0.012564f
C862 VDD1.n66 VSUBS 0.028046f
C863 VDD1.n67 VSUBS 0.028046f
C864 VDD1.n68 VSUBS 0.012564f
C865 VDD1.n69 VSUBS 0.011866f
C866 VDD1.n70 VSUBS 0.022082f
C867 VDD1.n71 VSUBS 0.022082f
C868 VDD1.n72 VSUBS 0.011866f
C869 VDD1.n73 VSUBS 0.012564f
C870 VDD1.n74 VSUBS 0.028046f
C871 VDD1.n75 VSUBS 0.028046f
C872 VDD1.n76 VSUBS 0.028046f
C873 VDD1.n77 VSUBS 0.012564f
C874 VDD1.n78 VSUBS 0.011866f
C875 VDD1.n79 VSUBS 0.022082f
C876 VDD1.n80 VSUBS 0.022082f
C877 VDD1.n81 VSUBS 0.011866f
C878 VDD1.n82 VSUBS 0.012215f
C879 VDD1.n83 VSUBS 0.012215f
C880 VDD1.n84 VSUBS 0.028046f
C881 VDD1.n85 VSUBS 0.067264f
C882 VDD1.n86 VSUBS 0.012564f
C883 VDD1.n87 VSUBS 0.011866f
C884 VDD1.n88 VSUBS 0.056772f
C885 VDD1.n89 VSUBS 0.054159f
C886 VDD1.t3 VSUBS 0.151987f
C887 VDD1.t5 VSUBS 0.151987f
C888 VDD1.n90 VSUBS 1.12751f
C889 VDD1.n91 VSUBS 2.37801f
C890 VDD1.t2 VSUBS 0.151987f
C891 VDD1.t1 VSUBS 0.151987f
C892 VDD1.n92 VSUBS 1.12394f
C893 VDD1.n93 VSUBS 2.36435f
C894 VTAIL.t4 VSUBS 0.209847f
C895 VTAIL.t1 VSUBS 0.209847f
C896 VTAIL.n0 VSUBS 1.42379f
C897 VTAIL.n1 VSUBS 0.828636f
C898 VTAIL.n2 VSUBS 0.033243f
C899 VTAIL.n3 VSUBS 0.030488f
C900 VTAIL.n4 VSUBS 0.016383f
C901 VTAIL.n5 VSUBS 0.038724f
C902 VTAIL.n6 VSUBS 0.017347f
C903 VTAIL.n7 VSUBS 0.030488f
C904 VTAIL.n8 VSUBS 0.016383f
C905 VTAIL.n9 VSUBS 0.038724f
C906 VTAIL.n10 VSUBS 0.017347f
C907 VTAIL.n11 VSUBS 0.030488f
C908 VTAIL.n12 VSUBS 0.016383f
C909 VTAIL.n13 VSUBS 0.038724f
C910 VTAIL.n14 VSUBS 0.017347f
C911 VTAIL.n15 VSUBS 0.19484f
C912 VTAIL.t8 VSUBS 0.083203f
C913 VTAIL.n16 VSUBS 0.029043f
C914 VTAIL.n17 VSUBS 0.02913f
C915 VTAIL.n18 VSUBS 0.016383f
C916 VTAIL.n19 VSUBS 1.0583f
C917 VTAIL.n20 VSUBS 0.030488f
C918 VTAIL.n21 VSUBS 0.016383f
C919 VTAIL.n22 VSUBS 0.017347f
C920 VTAIL.n23 VSUBS 0.038724f
C921 VTAIL.n24 VSUBS 0.038724f
C922 VTAIL.n25 VSUBS 0.017347f
C923 VTAIL.n26 VSUBS 0.016383f
C924 VTAIL.n27 VSUBS 0.030488f
C925 VTAIL.n28 VSUBS 0.030488f
C926 VTAIL.n29 VSUBS 0.016383f
C927 VTAIL.n30 VSUBS 0.017347f
C928 VTAIL.n31 VSUBS 0.038724f
C929 VTAIL.n32 VSUBS 0.038724f
C930 VTAIL.n33 VSUBS 0.038724f
C931 VTAIL.n34 VSUBS 0.017347f
C932 VTAIL.n35 VSUBS 0.016383f
C933 VTAIL.n36 VSUBS 0.030488f
C934 VTAIL.n37 VSUBS 0.030488f
C935 VTAIL.n38 VSUBS 0.016383f
C936 VTAIL.n39 VSUBS 0.016865f
C937 VTAIL.n40 VSUBS 0.016865f
C938 VTAIL.n41 VSUBS 0.038724f
C939 VTAIL.n42 VSUBS 0.092871f
C940 VTAIL.n43 VSUBS 0.017347f
C941 VTAIL.n44 VSUBS 0.016383f
C942 VTAIL.n45 VSUBS 0.078385f
C943 VTAIL.n46 VSUBS 0.046897f
C944 VTAIL.n47 VSUBS 0.412042f
C945 VTAIL.t9 VSUBS 0.209847f
C946 VTAIL.t10 VSUBS 0.209847f
C947 VTAIL.n48 VSUBS 1.42379f
C948 VTAIL.n49 VSUBS 2.43161f
C949 VTAIL.t11 VSUBS 0.209847f
C950 VTAIL.t0 VSUBS 0.209847f
C951 VTAIL.n50 VSUBS 1.4238f
C952 VTAIL.n51 VSUBS 2.4316f
C953 VTAIL.n52 VSUBS 0.033243f
C954 VTAIL.n53 VSUBS 0.030488f
C955 VTAIL.n54 VSUBS 0.016383f
C956 VTAIL.n55 VSUBS 0.038724f
C957 VTAIL.n56 VSUBS 0.017347f
C958 VTAIL.n57 VSUBS 0.030488f
C959 VTAIL.n58 VSUBS 0.016383f
C960 VTAIL.n59 VSUBS 0.038724f
C961 VTAIL.n60 VSUBS 0.038724f
C962 VTAIL.n61 VSUBS 0.017347f
C963 VTAIL.n62 VSUBS 0.030488f
C964 VTAIL.n63 VSUBS 0.016383f
C965 VTAIL.n64 VSUBS 0.038724f
C966 VTAIL.n65 VSUBS 0.017347f
C967 VTAIL.n66 VSUBS 0.19484f
C968 VTAIL.t2 VSUBS 0.083203f
C969 VTAIL.n67 VSUBS 0.029043f
C970 VTAIL.n68 VSUBS 0.02913f
C971 VTAIL.n69 VSUBS 0.016383f
C972 VTAIL.n70 VSUBS 1.0583f
C973 VTAIL.n71 VSUBS 0.030488f
C974 VTAIL.n72 VSUBS 0.016383f
C975 VTAIL.n73 VSUBS 0.017347f
C976 VTAIL.n74 VSUBS 0.038724f
C977 VTAIL.n75 VSUBS 0.038724f
C978 VTAIL.n76 VSUBS 0.017347f
C979 VTAIL.n77 VSUBS 0.016383f
C980 VTAIL.n78 VSUBS 0.030488f
C981 VTAIL.n79 VSUBS 0.030488f
C982 VTAIL.n80 VSUBS 0.016383f
C983 VTAIL.n81 VSUBS 0.017347f
C984 VTAIL.n82 VSUBS 0.038724f
C985 VTAIL.n83 VSUBS 0.038724f
C986 VTAIL.n84 VSUBS 0.017347f
C987 VTAIL.n85 VSUBS 0.016383f
C988 VTAIL.n86 VSUBS 0.030488f
C989 VTAIL.n87 VSUBS 0.030488f
C990 VTAIL.n88 VSUBS 0.016383f
C991 VTAIL.n89 VSUBS 0.016865f
C992 VTAIL.n90 VSUBS 0.016865f
C993 VTAIL.n91 VSUBS 0.038724f
C994 VTAIL.n92 VSUBS 0.092871f
C995 VTAIL.n93 VSUBS 0.017347f
C996 VTAIL.n94 VSUBS 0.016383f
C997 VTAIL.n95 VSUBS 0.078385f
C998 VTAIL.n96 VSUBS 0.046897f
C999 VTAIL.n97 VSUBS 0.412042f
C1000 VTAIL.t7 VSUBS 0.209847f
C1001 VTAIL.t5 VSUBS 0.209847f
C1002 VTAIL.n98 VSUBS 1.4238f
C1003 VTAIL.n99 VSUBS 0.990595f
C1004 VTAIL.n100 VSUBS 0.033243f
C1005 VTAIL.n101 VSUBS 0.030488f
C1006 VTAIL.n102 VSUBS 0.016383f
C1007 VTAIL.n103 VSUBS 0.038724f
C1008 VTAIL.n104 VSUBS 0.017347f
C1009 VTAIL.n105 VSUBS 0.030488f
C1010 VTAIL.n106 VSUBS 0.016383f
C1011 VTAIL.n107 VSUBS 0.038724f
C1012 VTAIL.n108 VSUBS 0.038724f
C1013 VTAIL.n109 VSUBS 0.017347f
C1014 VTAIL.n110 VSUBS 0.030488f
C1015 VTAIL.n111 VSUBS 0.016383f
C1016 VTAIL.n112 VSUBS 0.038724f
C1017 VTAIL.n113 VSUBS 0.017347f
C1018 VTAIL.n114 VSUBS 0.19484f
C1019 VTAIL.t6 VSUBS 0.083203f
C1020 VTAIL.n115 VSUBS 0.029043f
C1021 VTAIL.n116 VSUBS 0.02913f
C1022 VTAIL.n117 VSUBS 0.016383f
C1023 VTAIL.n118 VSUBS 1.0583f
C1024 VTAIL.n119 VSUBS 0.030488f
C1025 VTAIL.n120 VSUBS 0.016383f
C1026 VTAIL.n121 VSUBS 0.017347f
C1027 VTAIL.n122 VSUBS 0.038724f
C1028 VTAIL.n123 VSUBS 0.038724f
C1029 VTAIL.n124 VSUBS 0.017347f
C1030 VTAIL.n125 VSUBS 0.016383f
C1031 VTAIL.n126 VSUBS 0.030488f
C1032 VTAIL.n127 VSUBS 0.030488f
C1033 VTAIL.n128 VSUBS 0.016383f
C1034 VTAIL.n129 VSUBS 0.017347f
C1035 VTAIL.n130 VSUBS 0.038724f
C1036 VTAIL.n131 VSUBS 0.038724f
C1037 VTAIL.n132 VSUBS 0.017347f
C1038 VTAIL.n133 VSUBS 0.016383f
C1039 VTAIL.n134 VSUBS 0.030488f
C1040 VTAIL.n135 VSUBS 0.030488f
C1041 VTAIL.n136 VSUBS 0.016383f
C1042 VTAIL.n137 VSUBS 0.016865f
C1043 VTAIL.n138 VSUBS 0.016865f
C1044 VTAIL.n139 VSUBS 0.038724f
C1045 VTAIL.n140 VSUBS 0.092871f
C1046 VTAIL.n141 VSUBS 0.017347f
C1047 VTAIL.n142 VSUBS 0.016383f
C1048 VTAIL.n143 VSUBS 0.078385f
C1049 VTAIL.n144 VSUBS 0.046897f
C1050 VTAIL.n145 VSUBS 1.62947f
C1051 VTAIL.n146 VSUBS 0.033243f
C1052 VTAIL.n147 VSUBS 0.030488f
C1053 VTAIL.n148 VSUBS 0.016383f
C1054 VTAIL.n149 VSUBS 0.038724f
C1055 VTAIL.n150 VSUBS 0.017347f
C1056 VTAIL.n151 VSUBS 0.030488f
C1057 VTAIL.n152 VSUBS 0.016383f
C1058 VTAIL.n153 VSUBS 0.038724f
C1059 VTAIL.n154 VSUBS 0.017347f
C1060 VTAIL.n155 VSUBS 0.030488f
C1061 VTAIL.n156 VSUBS 0.016383f
C1062 VTAIL.n157 VSUBS 0.038724f
C1063 VTAIL.n158 VSUBS 0.017347f
C1064 VTAIL.n159 VSUBS 0.19484f
C1065 VTAIL.t3 VSUBS 0.083203f
C1066 VTAIL.n160 VSUBS 0.029043f
C1067 VTAIL.n161 VSUBS 0.02913f
C1068 VTAIL.n162 VSUBS 0.016383f
C1069 VTAIL.n163 VSUBS 1.0583f
C1070 VTAIL.n164 VSUBS 0.030488f
C1071 VTAIL.n165 VSUBS 0.016383f
C1072 VTAIL.n166 VSUBS 0.017347f
C1073 VTAIL.n167 VSUBS 0.038724f
C1074 VTAIL.n168 VSUBS 0.038724f
C1075 VTAIL.n169 VSUBS 0.017347f
C1076 VTAIL.n170 VSUBS 0.016383f
C1077 VTAIL.n171 VSUBS 0.030488f
C1078 VTAIL.n172 VSUBS 0.030488f
C1079 VTAIL.n173 VSUBS 0.016383f
C1080 VTAIL.n174 VSUBS 0.017347f
C1081 VTAIL.n175 VSUBS 0.038724f
C1082 VTAIL.n176 VSUBS 0.038724f
C1083 VTAIL.n177 VSUBS 0.038724f
C1084 VTAIL.n178 VSUBS 0.017347f
C1085 VTAIL.n179 VSUBS 0.016383f
C1086 VTAIL.n180 VSUBS 0.030488f
C1087 VTAIL.n181 VSUBS 0.030488f
C1088 VTAIL.n182 VSUBS 0.016383f
C1089 VTAIL.n183 VSUBS 0.016865f
C1090 VTAIL.n184 VSUBS 0.016865f
C1091 VTAIL.n185 VSUBS 0.038724f
C1092 VTAIL.n186 VSUBS 0.092871f
C1093 VTAIL.n187 VSUBS 0.017347f
C1094 VTAIL.n188 VSUBS 0.016383f
C1095 VTAIL.n189 VSUBS 0.078385f
C1096 VTAIL.n190 VSUBS 0.046897f
C1097 VTAIL.n191 VSUBS 1.56785f
C1098 VP.n0 VSUBS 0.048325f
C1099 VP.t0 VSUBS 1.98768f
C1100 VP.n1 VSUBS 0.032005f
C1101 VP.n2 VSUBS 0.036654f
C1102 VP.t2 VSUBS 1.98768f
C1103 VP.n3 VSUBS 0.074038f
C1104 VP.n4 VSUBS 0.036654f
C1105 VP.t5 VSUBS 1.98768f
C1106 VP.n5 VSUBS 0.850552f
C1107 VP.n6 VSUBS 0.048325f
C1108 VP.t4 VSUBS 1.98768f
C1109 VP.n7 VSUBS 0.032005f
C1110 VP.n8 VSUBS 0.315628f
C1111 VP.t3 VSUBS 1.98768f
C1112 VP.t1 VSUBS 2.24052f
C1113 VP.n9 VSUBS 0.801178f
C1114 VP.n10 VSUBS 0.820011f
C1115 VP.n11 VSUBS 0.05145f
C1116 VP.n12 VSUBS 0.074038f
C1117 VP.n13 VSUBS 0.036654f
C1118 VP.n14 VSUBS 0.036654f
C1119 VP.n15 VSUBS 0.036654f
C1120 VP.n16 VSUBS 0.069288f
C1121 VP.n17 VSUBS 0.060894f
C1122 VP.n18 VSUBS 0.850552f
C1123 VP.n19 VSUBS 1.7362f
C1124 VP.n20 VSUBS 1.76539f
C1125 VP.n21 VSUBS 0.048325f
C1126 VP.n22 VSUBS 0.060894f
C1127 VP.n23 VSUBS 0.069288f
C1128 VP.n24 VSUBS 0.032005f
C1129 VP.n25 VSUBS 0.036654f
C1130 VP.n26 VSUBS 0.036654f
C1131 VP.n27 VSUBS 0.036654f
C1132 VP.n28 VSUBS 0.05145f
C1133 VP.n29 VSUBS 0.722651f
C1134 VP.n30 VSUBS 0.05145f
C1135 VP.n31 VSUBS 0.074038f
C1136 VP.n32 VSUBS 0.036654f
C1137 VP.n33 VSUBS 0.036654f
C1138 VP.n34 VSUBS 0.036654f
C1139 VP.n35 VSUBS 0.069288f
C1140 VP.n36 VSUBS 0.060894f
C1141 VP.n37 VSUBS 0.850552f
C1142 VP.n38 VSUBS 0.047219f
.ends

