* NGSPICE file created from diff_pair_sample_0555.ext - technology: sky130A

.subckt diff_pair_sample_0555 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=3.06
X1 VTAIL.t7 VN.t0 VDD2.t9 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X2 VTAIL.t19 VN.t1 VDD2.t8 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X3 VTAIL.t15 VP.t1 VDD1.t8 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X4 VDD2.t7 VN.t2 VTAIL.t4 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=3.06
X5 VDD2.t6 VN.t3 VTAIL.t5 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=3.06
X6 VDD1.t7 VP.t2 VTAIL.t9 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=3.06
X7 VTAIL.t13 VP.t3 VDD1.t6 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X8 B.t11 B.t9 B.t10 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=3.06
X9 VDD2.t5 VN.t4 VTAIL.t18 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=3.06
X10 VDD2.t4 VN.t5 VTAIL.t2 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X11 VDD1.t5 VP.t4 VTAIL.t11 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X12 VTAIL.t0 VN.t6 VDD2.t3 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X13 B.t8 B.t6 B.t7 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=3.06
X14 VDD1.t4 VP.t5 VTAIL.t16 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X15 B.t5 B.t3 B.t4 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=3.06
X16 VTAIL.t8 VP.t6 VDD1.t3 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X17 VDD1.t2 VP.t7 VTAIL.t14 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=3.06
X18 B.t2 B.t0 B.t1 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0 ps=0 w=4.48 l=3.06
X19 VDD2.t2 VN.t7 VTAIL.t6 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X20 VDD2.t1 VN.t8 VTAIL.t3 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=1.7472 pd=9.74 as=0.7392 ps=4.81 w=4.48 l=3.06
X21 VTAIL.t17 VP.t8 VDD1.t1 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
X22 VDD1.t0 VP.t9 VTAIL.t10 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=1.7472 ps=9.74 w=4.48 l=3.06
X23 VTAIL.t1 VN.t9 VDD2.t0 w_n5038_n1864# sky130_fd_pr__pfet_01v8 ad=0.7392 pd=4.81 as=0.7392 ps=4.81 w=4.48 l=3.06
R0 VP.n29 VP.n28 161.3
R1 VP.n30 VP.n25 161.3
R2 VP.n32 VP.n31 161.3
R3 VP.n33 VP.n24 161.3
R4 VP.n35 VP.n34 161.3
R5 VP.n36 VP.n23 161.3
R6 VP.n38 VP.n37 161.3
R7 VP.n39 VP.n22 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n42 VP.n21 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n45 VP.n20 161.3
R12 VP.n47 VP.n46 161.3
R13 VP.n49 VP.n48 161.3
R14 VP.n50 VP.n18 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n17 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n16 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n94 VP.n93 161.3
R27 VP.n92 VP.n91 161.3
R28 VP.n90 VP.n5 161.3
R29 VP.n89 VP.n88 161.3
R30 VP.n87 VP.n6 161.3
R31 VP.n86 VP.n85 161.3
R32 VP.n84 VP.n7 161.3
R33 VP.n83 VP.n82 161.3
R34 VP.n81 VP.n8 161.3
R35 VP.n80 VP.n79 161.3
R36 VP.n78 VP.n9 161.3
R37 VP.n77 VP.n76 161.3
R38 VP.n75 VP.n10 161.3
R39 VP.n74 VP.n73 161.3
R40 VP.n71 VP.n11 161.3
R41 VP.n70 VP.n69 161.3
R42 VP.n68 VP.n12 161.3
R43 VP.n67 VP.n66 161.3
R44 VP.n65 VP.n13 161.3
R45 VP.n64 VP.n63 161.3
R46 VP.n62 VP.n14 161.3
R47 VP.n61 VP.n60 76.4741
R48 VP.n104 VP.n0 76.4741
R49 VP.n59 VP.n15 76.4741
R50 VP.n26 VP.t7 68.2829
R51 VP.n78 VP.n77 56.5617
R52 VP.n89 VP.n6 56.5617
R53 VP.n44 VP.n21 56.5617
R54 VP.n33 VP.n32 56.5617
R55 VP.n27 VP.n26 55.0126
R56 VP.n61 VP.n59 49.9579
R57 VP.n66 VP.n65 48.8116
R58 VP.n100 VP.n2 48.8116
R59 VP.n55 VP.n17 48.8116
R60 VP.n83 VP.t5 35.2842
R61 VP.n60 VP.t2 35.2842
R62 VP.n72 VP.t8 35.2842
R63 VP.n4 VP.t3 35.2842
R64 VP.n0 VP.t9 35.2842
R65 VP.n38 VP.t4 35.2842
R66 VP.n15 VP.t0 35.2842
R67 VP.n19 VP.t1 35.2842
R68 VP.n27 VP.t6 35.2842
R69 VP.n66 VP.n12 32.3425
R70 VP.n96 VP.n2 32.3425
R71 VP.n51 VP.n17 32.3425
R72 VP.n64 VP.n14 24.5923
R73 VP.n65 VP.n64 24.5923
R74 VP.n70 VP.n12 24.5923
R75 VP.n71 VP.n70 24.5923
R76 VP.n73 VP.n10 24.5923
R77 VP.n77 VP.n10 24.5923
R78 VP.n79 VP.n78 24.5923
R79 VP.n79 VP.n8 24.5923
R80 VP.n83 VP.n8 24.5923
R81 VP.n84 VP.n83 24.5923
R82 VP.n85 VP.n84 24.5923
R83 VP.n85 VP.n6 24.5923
R84 VP.n90 VP.n89 24.5923
R85 VP.n91 VP.n90 24.5923
R86 VP.n95 VP.n94 24.5923
R87 VP.n96 VP.n95 24.5923
R88 VP.n101 VP.n100 24.5923
R89 VP.n102 VP.n101 24.5923
R90 VP.n56 VP.n55 24.5923
R91 VP.n57 VP.n56 24.5923
R92 VP.n45 VP.n44 24.5923
R93 VP.n46 VP.n45 24.5923
R94 VP.n50 VP.n49 24.5923
R95 VP.n51 VP.n50 24.5923
R96 VP.n34 VP.n33 24.5923
R97 VP.n34 VP.n23 24.5923
R98 VP.n38 VP.n23 24.5923
R99 VP.n39 VP.n38 24.5923
R100 VP.n40 VP.n39 24.5923
R101 VP.n40 VP.n21 24.5923
R102 VP.n28 VP.n25 24.5923
R103 VP.n32 VP.n25 24.5923
R104 VP.n73 VP.n72 19.1821
R105 VP.n91 VP.n4 19.1821
R106 VP.n46 VP.n19 19.1821
R107 VP.n28 VP.n27 19.1821
R108 VP.n60 VP.n14 13.7719
R109 VP.n102 VP.n0 13.7719
R110 VP.n57 VP.n15 13.7719
R111 VP.n72 VP.n71 5.4107
R112 VP.n94 VP.n4 5.4107
R113 VP.n49 VP.n19 5.4107
R114 VP.n29 VP.n26 4.192
R115 VP.n59 VP.n58 0.354861
R116 VP.n62 VP.n61 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n30 VP.n29 0.189894
R120 VP.n31 VP.n30 0.189894
R121 VP.n31 VP.n24 0.189894
R122 VP.n35 VP.n24 0.189894
R123 VP.n36 VP.n35 0.189894
R124 VP.n37 VP.n36 0.189894
R125 VP.n37 VP.n22 0.189894
R126 VP.n41 VP.n22 0.189894
R127 VP.n42 VP.n41 0.189894
R128 VP.n43 VP.n42 0.189894
R129 VP.n43 VP.n20 0.189894
R130 VP.n47 VP.n20 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n18 0.189894
R133 VP.n52 VP.n18 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n16 0.189894
R137 VP.n58 VP.n16 0.189894
R138 VP.n63 VP.n62 0.189894
R139 VP.n63 VP.n13 0.189894
R140 VP.n67 VP.n13 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n69 VP.n68 0.189894
R143 VP.n69 VP.n11 0.189894
R144 VP.n74 VP.n11 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n76 VP.n75 0.189894
R147 VP.n76 VP.n9 0.189894
R148 VP.n80 VP.n9 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n82 VP.n81 0.189894
R151 VP.n82 VP.n7 0.189894
R152 VP.n86 VP.n7 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n88 VP.n87 0.189894
R155 VP.n88 VP.n5 0.189894
R156 VP.n92 VP.n5 0.189894
R157 VP.n93 VP.n92 0.189894
R158 VP.n93 VP.n3 0.189894
R159 VP.n97 VP.n3 0.189894
R160 VP.n98 VP.n97 0.189894
R161 VP.n99 VP.n98 0.189894
R162 VP.n99 VP.n1 0.189894
R163 VP.n103 VP.n1 0.189894
R164 VTAIL.n104 VTAIL.n86 756.745
R165 VTAIL.n20 VTAIL.n2 756.745
R166 VTAIL.n80 VTAIL.n62 756.745
R167 VTAIL.n52 VTAIL.n34 756.745
R168 VTAIL.n95 VTAIL.n94 585
R169 VTAIL.n97 VTAIL.n96 585
R170 VTAIL.n90 VTAIL.n89 585
R171 VTAIL.n103 VTAIL.n102 585
R172 VTAIL.n105 VTAIL.n104 585
R173 VTAIL.n11 VTAIL.n10 585
R174 VTAIL.n13 VTAIL.n12 585
R175 VTAIL.n6 VTAIL.n5 585
R176 VTAIL.n19 VTAIL.n18 585
R177 VTAIL.n21 VTAIL.n20 585
R178 VTAIL.n81 VTAIL.n80 585
R179 VTAIL.n79 VTAIL.n78 585
R180 VTAIL.n66 VTAIL.n65 585
R181 VTAIL.n73 VTAIL.n72 585
R182 VTAIL.n71 VTAIL.n70 585
R183 VTAIL.n53 VTAIL.n52 585
R184 VTAIL.n51 VTAIL.n50 585
R185 VTAIL.n38 VTAIL.n37 585
R186 VTAIL.n45 VTAIL.n44 585
R187 VTAIL.n43 VTAIL.n42 585
R188 VTAIL.n93 VTAIL.t4 328.587
R189 VTAIL.n9 VTAIL.t10 328.587
R190 VTAIL.n69 VTAIL.t12 328.587
R191 VTAIL.n41 VTAIL.t18 328.587
R192 VTAIL.n96 VTAIL.n95 171.744
R193 VTAIL.n96 VTAIL.n89 171.744
R194 VTAIL.n103 VTAIL.n89 171.744
R195 VTAIL.n104 VTAIL.n103 171.744
R196 VTAIL.n12 VTAIL.n11 171.744
R197 VTAIL.n12 VTAIL.n5 171.744
R198 VTAIL.n19 VTAIL.n5 171.744
R199 VTAIL.n20 VTAIL.n19 171.744
R200 VTAIL.n80 VTAIL.n79 171.744
R201 VTAIL.n79 VTAIL.n65 171.744
R202 VTAIL.n72 VTAIL.n65 171.744
R203 VTAIL.n72 VTAIL.n71 171.744
R204 VTAIL.n52 VTAIL.n51 171.744
R205 VTAIL.n51 VTAIL.n37 171.744
R206 VTAIL.n44 VTAIL.n37 171.744
R207 VTAIL.n44 VTAIL.n43 171.744
R208 VTAIL.n95 VTAIL.t4 85.8723
R209 VTAIL.n11 VTAIL.t10 85.8723
R210 VTAIL.n71 VTAIL.t12 85.8723
R211 VTAIL.n43 VTAIL.t18 85.8723
R212 VTAIL.n61 VTAIL.n60 85.8495
R213 VTAIL.n59 VTAIL.n58 85.8495
R214 VTAIL.n33 VTAIL.n32 85.8495
R215 VTAIL.n31 VTAIL.n30 85.8495
R216 VTAIL.n111 VTAIL.n110 85.8494
R217 VTAIL.n1 VTAIL.n0 85.8494
R218 VTAIL.n27 VTAIL.n26 85.8494
R219 VTAIL.n29 VTAIL.n28 85.8494
R220 VTAIL.n109 VTAIL.n108 30.6338
R221 VTAIL.n25 VTAIL.n24 30.6338
R222 VTAIL.n85 VTAIL.n84 30.6338
R223 VTAIL.n57 VTAIL.n56 30.6338
R224 VTAIL.n31 VTAIL.n29 22.0738
R225 VTAIL.n109 VTAIL.n85 19.1514
R226 VTAIL.n94 VTAIL.n93 16.3651
R227 VTAIL.n10 VTAIL.n9 16.3651
R228 VTAIL.n70 VTAIL.n69 16.3651
R229 VTAIL.n42 VTAIL.n41 16.3651
R230 VTAIL.n97 VTAIL.n92 12.8005
R231 VTAIL.n13 VTAIL.n8 12.8005
R232 VTAIL.n73 VTAIL.n68 12.8005
R233 VTAIL.n45 VTAIL.n40 12.8005
R234 VTAIL.n98 VTAIL.n90 12.0247
R235 VTAIL.n14 VTAIL.n6 12.0247
R236 VTAIL.n74 VTAIL.n66 12.0247
R237 VTAIL.n46 VTAIL.n38 12.0247
R238 VTAIL.n102 VTAIL.n101 11.249
R239 VTAIL.n18 VTAIL.n17 11.249
R240 VTAIL.n78 VTAIL.n77 11.249
R241 VTAIL.n50 VTAIL.n49 11.249
R242 VTAIL.n105 VTAIL.n88 10.4732
R243 VTAIL.n21 VTAIL.n4 10.4732
R244 VTAIL.n81 VTAIL.n64 10.4732
R245 VTAIL.n53 VTAIL.n36 10.4732
R246 VTAIL.n106 VTAIL.n86 9.69747
R247 VTAIL.n22 VTAIL.n2 9.69747
R248 VTAIL.n82 VTAIL.n62 9.69747
R249 VTAIL.n54 VTAIL.n34 9.69747
R250 VTAIL.n108 VTAIL.n107 9.45567
R251 VTAIL.n24 VTAIL.n23 9.45567
R252 VTAIL.n84 VTAIL.n83 9.45567
R253 VTAIL.n56 VTAIL.n55 9.45567
R254 VTAIL.n107 VTAIL.n106 9.3005
R255 VTAIL.n88 VTAIL.n87 9.3005
R256 VTAIL.n101 VTAIL.n100 9.3005
R257 VTAIL.n99 VTAIL.n98 9.3005
R258 VTAIL.n92 VTAIL.n91 9.3005
R259 VTAIL.n23 VTAIL.n22 9.3005
R260 VTAIL.n4 VTAIL.n3 9.3005
R261 VTAIL.n17 VTAIL.n16 9.3005
R262 VTAIL.n15 VTAIL.n14 9.3005
R263 VTAIL.n8 VTAIL.n7 9.3005
R264 VTAIL.n83 VTAIL.n82 9.3005
R265 VTAIL.n64 VTAIL.n63 9.3005
R266 VTAIL.n77 VTAIL.n76 9.3005
R267 VTAIL.n75 VTAIL.n74 9.3005
R268 VTAIL.n68 VTAIL.n67 9.3005
R269 VTAIL.n55 VTAIL.n54 9.3005
R270 VTAIL.n36 VTAIL.n35 9.3005
R271 VTAIL.n49 VTAIL.n48 9.3005
R272 VTAIL.n47 VTAIL.n46 9.3005
R273 VTAIL.n40 VTAIL.n39 9.3005
R274 VTAIL.n110 VTAIL.t6 7.25608
R275 VTAIL.n110 VTAIL.t1 7.25608
R276 VTAIL.n0 VTAIL.t3 7.25608
R277 VTAIL.n0 VTAIL.t19 7.25608
R278 VTAIL.n26 VTAIL.t16 7.25608
R279 VTAIL.n26 VTAIL.t13 7.25608
R280 VTAIL.n28 VTAIL.t9 7.25608
R281 VTAIL.n28 VTAIL.t17 7.25608
R282 VTAIL.n60 VTAIL.t11 7.25608
R283 VTAIL.n60 VTAIL.t15 7.25608
R284 VTAIL.n58 VTAIL.t14 7.25608
R285 VTAIL.n58 VTAIL.t8 7.25608
R286 VTAIL.n32 VTAIL.t2 7.25608
R287 VTAIL.n32 VTAIL.t0 7.25608
R288 VTAIL.n30 VTAIL.t5 7.25608
R289 VTAIL.n30 VTAIL.t7 7.25608
R290 VTAIL.n108 VTAIL.n86 4.26717
R291 VTAIL.n24 VTAIL.n2 4.26717
R292 VTAIL.n84 VTAIL.n62 4.26717
R293 VTAIL.n56 VTAIL.n34 4.26717
R294 VTAIL.n93 VTAIL.n91 3.73474
R295 VTAIL.n9 VTAIL.n7 3.73474
R296 VTAIL.n69 VTAIL.n67 3.73474
R297 VTAIL.n41 VTAIL.n39 3.73474
R298 VTAIL.n106 VTAIL.n105 3.49141
R299 VTAIL.n22 VTAIL.n21 3.49141
R300 VTAIL.n82 VTAIL.n81 3.49141
R301 VTAIL.n54 VTAIL.n53 3.49141
R302 VTAIL.n33 VTAIL.n31 2.92291
R303 VTAIL.n57 VTAIL.n33 2.92291
R304 VTAIL.n61 VTAIL.n59 2.92291
R305 VTAIL.n85 VTAIL.n61 2.92291
R306 VTAIL.n29 VTAIL.n27 2.92291
R307 VTAIL.n27 VTAIL.n25 2.92291
R308 VTAIL.n111 VTAIL.n109 2.92291
R309 VTAIL.n102 VTAIL.n88 2.71565
R310 VTAIL.n18 VTAIL.n4 2.71565
R311 VTAIL.n78 VTAIL.n64 2.71565
R312 VTAIL.n50 VTAIL.n36 2.71565
R313 VTAIL VTAIL.n1 2.2505
R314 VTAIL.n101 VTAIL.n90 1.93989
R315 VTAIL.n17 VTAIL.n6 1.93989
R316 VTAIL.n77 VTAIL.n66 1.93989
R317 VTAIL.n49 VTAIL.n38 1.93989
R318 VTAIL.n59 VTAIL.n57 1.93153
R319 VTAIL.n25 VTAIL.n1 1.93153
R320 VTAIL.n98 VTAIL.n97 1.16414
R321 VTAIL.n14 VTAIL.n13 1.16414
R322 VTAIL.n74 VTAIL.n73 1.16414
R323 VTAIL.n46 VTAIL.n45 1.16414
R324 VTAIL VTAIL.n111 0.672914
R325 VTAIL.n94 VTAIL.n92 0.388379
R326 VTAIL.n10 VTAIL.n8 0.388379
R327 VTAIL.n70 VTAIL.n68 0.388379
R328 VTAIL.n42 VTAIL.n40 0.388379
R329 VTAIL.n99 VTAIL.n91 0.155672
R330 VTAIL.n100 VTAIL.n99 0.155672
R331 VTAIL.n100 VTAIL.n87 0.155672
R332 VTAIL.n107 VTAIL.n87 0.155672
R333 VTAIL.n15 VTAIL.n7 0.155672
R334 VTAIL.n16 VTAIL.n15 0.155672
R335 VTAIL.n16 VTAIL.n3 0.155672
R336 VTAIL.n23 VTAIL.n3 0.155672
R337 VTAIL.n83 VTAIL.n63 0.155672
R338 VTAIL.n76 VTAIL.n63 0.155672
R339 VTAIL.n76 VTAIL.n75 0.155672
R340 VTAIL.n75 VTAIL.n67 0.155672
R341 VTAIL.n55 VTAIL.n35 0.155672
R342 VTAIL.n48 VTAIL.n35 0.155672
R343 VTAIL.n48 VTAIL.n47 0.155672
R344 VTAIL.n47 VTAIL.n39 0.155672
R345 VDD1.n18 VDD1.n0 756.745
R346 VDD1.n43 VDD1.n25 756.745
R347 VDD1.n19 VDD1.n18 585
R348 VDD1.n17 VDD1.n16 585
R349 VDD1.n4 VDD1.n3 585
R350 VDD1.n11 VDD1.n10 585
R351 VDD1.n9 VDD1.n8 585
R352 VDD1.n34 VDD1.n33 585
R353 VDD1.n36 VDD1.n35 585
R354 VDD1.n29 VDD1.n28 585
R355 VDD1.n42 VDD1.n41 585
R356 VDD1.n44 VDD1.n43 585
R357 VDD1.n7 VDD1.t2 328.587
R358 VDD1.n32 VDD1.t7 328.587
R359 VDD1.n18 VDD1.n17 171.744
R360 VDD1.n17 VDD1.n3 171.744
R361 VDD1.n10 VDD1.n3 171.744
R362 VDD1.n10 VDD1.n9 171.744
R363 VDD1.n35 VDD1.n34 171.744
R364 VDD1.n35 VDD1.n28 171.744
R365 VDD1.n42 VDD1.n28 171.744
R366 VDD1.n43 VDD1.n42 171.744
R367 VDD1.n51 VDD1.n50 104.665
R368 VDD1.n24 VDD1.n23 102.528
R369 VDD1.n53 VDD1.n52 102.528
R370 VDD1.n49 VDD1.n48 102.528
R371 VDD1.n9 VDD1.t2 85.8723
R372 VDD1.n34 VDD1.t7 85.8723
R373 VDD1.n24 VDD1.n22 50.235
R374 VDD1.n49 VDD1.n47 50.235
R375 VDD1.n53 VDD1.n51 43.503
R376 VDD1.n8 VDD1.n7 16.3651
R377 VDD1.n33 VDD1.n32 16.3651
R378 VDD1.n11 VDD1.n6 12.8005
R379 VDD1.n36 VDD1.n31 12.8005
R380 VDD1.n12 VDD1.n4 12.0247
R381 VDD1.n37 VDD1.n29 12.0247
R382 VDD1.n16 VDD1.n15 11.249
R383 VDD1.n41 VDD1.n40 11.249
R384 VDD1.n19 VDD1.n2 10.4732
R385 VDD1.n44 VDD1.n27 10.4732
R386 VDD1.n20 VDD1.n0 9.69747
R387 VDD1.n45 VDD1.n25 9.69747
R388 VDD1.n22 VDD1.n21 9.45567
R389 VDD1.n47 VDD1.n46 9.45567
R390 VDD1.n21 VDD1.n20 9.3005
R391 VDD1.n2 VDD1.n1 9.3005
R392 VDD1.n15 VDD1.n14 9.3005
R393 VDD1.n13 VDD1.n12 9.3005
R394 VDD1.n6 VDD1.n5 9.3005
R395 VDD1.n46 VDD1.n45 9.3005
R396 VDD1.n27 VDD1.n26 9.3005
R397 VDD1.n40 VDD1.n39 9.3005
R398 VDD1.n38 VDD1.n37 9.3005
R399 VDD1.n31 VDD1.n30 9.3005
R400 VDD1.n52 VDD1.t8 7.25608
R401 VDD1.n52 VDD1.t9 7.25608
R402 VDD1.n23 VDD1.t3 7.25608
R403 VDD1.n23 VDD1.t5 7.25608
R404 VDD1.n50 VDD1.t6 7.25608
R405 VDD1.n50 VDD1.t0 7.25608
R406 VDD1.n48 VDD1.t1 7.25608
R407 VDD1.n48 VDD1.t4 7.25608
R408 VDD1.n22 VDD1.n0 4.26717
R409 VDD1.n47 VDD1.n25 4.26717
R410 VDD1.n7 VDD1.n5 3.73474
R411 VDD1.n32 VDD1.n30 3.73474
R412 VDD1.n20 VDD1.n19 3.49141
R413 VDD1.n45 VDD1.n44 3.49141
R414 VDD1.n16 VDD1.n2 2.71565
R415 VDD1.n41 VDD1.n27 2.71565
R416 VDD1 VDD1.n53 2.13412
R417 VDD1.n15 VDD1.n4 1.93989
R418 VDD1.n40 VDD1.n29 1.93989
R419 VDD1.n12 VDD1.n11 1.16414
R420 VDD1.n37 VDD1.n36 1.16414
R421 VDD1 VDD1.n24 0.789293
R422 VDD1.n51 VDD1.n49 0.675757
R423 VDD1.n8 VDD1.n6 0.388379
R424 VDD1.n33 VDD1.n31 0.388379
R425 VDD1.n21 VDD1.n1 0.155672
R426 VDD1.n14 VDD1.n1 0.155672
R427 VDD1.n14 VDD1.n13 0.155672
R428 VDD1.n13 VDD1.n5 0.155672
R429 VDD1.n38 VDD1.n30 0.155672
R430 VDD1.n39 VDD1.n38 0.155672
R431 VDD1.n39 VDD1.n26 0.155672
R432 VDD1.n46 VDD1.n26 0.155672
R433 VN.n88 VN.n87 161.3
R434 VN.n86 VN.n46 161.3
R435 VN.n85 VN.n84 161.3
R436 VN.n83 VN.n47 161.3
R437 VN.n82 VN.n81 161.3
R438 VN.n80 VN.n48 161.3
R439 VN.n79 VN.n78 161.3
R440 VN.n77 VN.n76 161.3
R441 VN.n75 VN.n50 161.3
R442 VN.n74 VN.n73 161.3
R443 VN.n72 VN.n51 161.3
R444 VN.n71 VN.n70 161.3
R445 VN.n69 VN.n52 161.3
R446 VN.n68 VN.n67 161.3
R447 VN.n66 VN.n53 161.3
R448 VN.n65 VN.n64 161.3
R449 VN.n63 VN.n54 161.3
R450 VN.n62 VN.n61 161.3
R451 VN.n60 VN.n55 161.3
R452 VN.n59 VN.n58 161.3
R453 VN.n43 VN.n42 161.3
R454 VN.n41 VN.n1 161.3
R455 VN.n40 VN.n39 161.3
R456 VN.n38 VN.n2 161.3
R457 VN.n37 VN.n36 161.3
R458 VN.n35 VN.n3 161.3
R459 VN.n34 VN.n33 161.3
R460 VN.n32 VN.n31 161.3
R461 VN.n30 VN.n5 161.3
R462 VN.n29 VN.n28 161.3
R463 VN.n27 VN.n6 161.3
R464 VN.n26 VN.n25 161.3
R465 VN.n24 VN.n7 161.3
R466 VN.n23 VN.n22 161.3
R467 VN.n21 VN.n8 161.3
R468 VN.n20 VN.n19 161.3
R469 VN.n18 VN.n9 161.3
R470 VN.n17 VN.n16 161.3
R471 VN.n15 VN.n10 161.3
R472 VN.n14 VN.n13 161.3
R473 VN.n44 VN.n0 76.4741
R474 VN.n89 VN.n45 76.4741
R475 VN.n56 VN.t4 68.2831
R476 VN.n11 VN.t8 68.2831
R477 VN.n18 VN.n17 56.5617
R478 VN.n29 VN.n6 56.5617
R479 VN.n63 VN.n62 56.5617
R480 VN.n74 VN.n51 56.5617
R481 VN.n12 VN.n11 55.0126
R482 VN.n57 VN.n56 55.0126
R483 VN VN.n89 50.1231
R484 VN.n40 VN.n2 48.8116
R485 VN.n85 VN.n47 48.8116
R486 VN.n23 VN.t7 35.2842
R487 VN.n12 VN.t1 35.2842
R488 VN.n4 VN.t9 35.2842
R489 VN.n0 VN.t2 35.2842
R490 VN.n68 VN.t5 35.2842
R491 VN.n57 VN.t6 35.2842
R492 VN.n49 VN.t0 35.2842
R493 VN.n45 VN.t3 35.2842
R494 VN.n36 VN.n2 32.3425
R495 VN.n81 VN.n47 32.3425
R496 VN.n13 VN.n10 24.5923
R497 VN.n17 VN.n10 24.5923
R498 VN.n19 VN.n18 24.5923
R499 VN.n19 VN.n8 24.5923
R500 VN.n23 VN.n8 24.5923
R501 VN.n24 VN.n23 24.5923
R502 VN.n25 VN.n24 24.5923
R503 VN.n25 VN.n6 24.5923
R504 VN.n30 VN.n29 24.5923
R505 VN.n31 VN.n30 24.5923
R506 VN.n35 VN.n34 24.5923
R507 VN.n36 VN.n35 24.5923
R508 VN.n41 VN.n40 24.5923
R509 VN.n42 VN.n41 24.5923
R510 VN.n62 VN.n55 24.5923
R511 VN.n58 VN.n55 24.5923
R512 VN.n70 VN.n51 24.5923
R513 VN.n70 VN.n69 24.5923
R514 VN.n69 VN.n68 24.5923
R515 VN.n68 VN.n53 24.5923
R516 VN.n64 VN.n53 24.5923
R517 VN.n64 VN.n63 24.5923
R518 VN.n81 VN.n80 24.5923
R519 VN.n80 VN.n79 24.5923
R520 VN.n76 VN.n75 24.5923
R521 VN.n75 VN.n74 24.5923
R522 VN.n87 VN.n86 24.5923
R523 VN.n86 VN.n85 24.5923
R524 VN.n13 VN.n12 19.1821
R525 VN.n31 VN.n4 19.1821
R526 VN.n58 VN.n57 19.1821
R527 VN.n76 VN.n49 19.1821
R528 VN.n42 VN.n0 13.7719
R529 VN.n87 VN.n45 13.7719
R530 VN.n34 VN.n4 5.4107
R531 VN.n79 VN.n49 5.4107
R532 VN.n59 VN.n56 4.19202
R533 VN.n14 VN.n11 4.19202
R534 VN.n89 VN.n88 0.354861
R535 VN.n44 VN.n43 0.354861
R536 VN VN.n44 0.267071
R537 VN.n88 VN.n46 0.189894
R538 VN.n84 VN.n46 0.189894
R539 VN.n84 VN.n83 0.189894
R540 VN.n83 VN.n82 0.189894
R541 VN.n82 VN.n48 0.189894
R542 VN.n78 VN.n48 0.189894
R543 VN.n78 VN.n77 0.189894
R544 VN.n77 VN.n50 0.189894
R545 VN.n73 VN.n50 0.189894
R546 VN.n73 VN.n72 0.189894
R547 VN.n72 VN.n71 0.189894
R548 VN.n71 VN.n52 0.189894
R549 VN.n67 VN.n52 0.189894
R550 VN.n67 VN.n66 0.189894
R551 VN.n66 VN.n65 0.189894
R552 VN.n65 VN.n54 0.189894
R553 VN.n61 VN.n54 0.189894
R554 VN.n61 VN.n60 0.189894
R555 VN.n60 VN.n59 0.189894
R556 VN.n15 VN.n14 0.189894
R557 VN.n16 VN.n15 0.189894
R558 VN.n16 VN.n9 0.189894
R559 VN.n20 VN.n9 0.189894
R560 VN.n21 VN.n20 0.189894
R561 VN.n22 VN.n21 0.189894
R562 VN.n22 VN.n7 0.189894
R563 VN.n26 VN.n7 0.189894
R564 VN.n27 VN.n26 0.189894
R565 VN.n28 VN.n27 0.189894
R566 VN.n28 VN.n5 0.189894
R567 VN.n32 VN.n5 0.189894
R568 VN.n33 VN.n32 0.189894
R569 VN.n33 VN.n3 0.189894
R570 VN.n37 VN.n3 0.189894
R571 VN.n38 VN.n37 0.189894
R572 VN.n39 VN.n38 0.189894
R573 VN.n39 VN.n1 0.189894
R574 VN.n43 VN.n1 0.189894
R575 VDD2.n45 VDD2.n27 756.745
R576 VDD2.n18 VDD2.n0 756.745
R577 VDD2.n46 VDD2.n45 585
R578 VDD2.n44 VDD2.n43 585
R579 VDD2.n31 VDD2.n30 585
R580 VDD2.n38 VDD2.n37 585
R581 VDD2.n36 VDD2.n35 585
R582 VDD2.n9 VDD2.n8 585
R583 VDD2.n11 VDD2.n10 585
R584 VDD2.n4 VDD2.n3 585
R585 VDD2.n17 VDD2.n16 585
R586 VDD2.n19 VDD2.n18 585
R587 VDD2.n34 VDD2.t6 328.587
R588 VDD2.n7 VDD2.t1 328.587
R589 VDD2.n45 VDD2.n44 171.744
R590 VDD2.n44 VDD2.n30 171.744
R591 VDD2.n37 VDD2.n30 171.744
R592 VDD2.n37 VDD2.n36 171.744
R593 VDD2.n10 VDD2.n9 171.744
R594 VDD2.n10 VDD2.n3 171.744
R595 VDD2.n17 VDD2.n3 171.744
R596 VDD2.n18 VDD2.n17 171.744
R597 VDD2.n26 VDD2.n25 104.665
R598 VDD2 VDD2.n53 104.662
R599 VDD2.n52 VDD2.n51 102.528
R600 VDD2.n24 VDD2.n23 102.528
R601 VDD2.n36 VDD2.t6 85.8723
R602 VDD2.n9 VDD2.t1 85.8723
R603 VDD2.n24 VDD2.n22 50.235
R604 VDD2.n50 VDD2.n49 47.3126
R605 VDD2.n50 VDD2.n26 41.4588
R606 VDD2.n35 VDD2.n34 16.3651
R607 VDD2.n8 VDD2.n7 16.3651
R608 VDD2.n38 VDD2.n33 12.8005
R609 VDD2.n11 VDD2.n6 12.8005
R610 VDD2.n39 VDD2.n31 12.0247
R611 VDD2.n12 VDD2.n4 12.0247
R612 VDD2.n43 VDD2.n42 11.249
R613 VDD2.n16 VDD2.n15 11.249
R614 VDD2.n46 VDD2.n29 10.4732
R615 VDD2.n19 VDD2.n2 10.4732
R616 VDD2.n47 VDD2.n27 9.69747
R617 VDD2.n20 VDD2.n0 9.69747
R618 VDD2.n49 VDD2.n48 9.45567
R619 VDD2.n22 VDD2.n21 9.45567
R620 VDD2.n48 VDD2.n47 9.3005
R621 VDD2.n29 VDD2.n28 9.3005
R622 VDD2.n42 VDD2.n41 9.3005
R623 VDD2.n40 VDD2.n39 9.3005
R624 VDD2.n33 VDD2.n32 9.3005
R625 VDD2.n21 VDD2.n20 9.3005
R626 VDD2.n2 VDD2.n1 9.3005
R627 VDD2.n15 VDD2.n14 9.3005
R628 VDD2.n13 VDD2.n12 9.3005
R629 VDD2.n6 VDD2.n5 9.3005
R630 VDD2.n53 VDD2.t3 7.25608
R631 VDD2.n53 VDD2.t5 7.25608
R632 VDD2.n51 VDD2.t9 7.25608
R633 VDD2.n51 VDD2.t4 7.25608
R634 VDD2.n25 VDD2.t0 7.25608
R635 VDD2.n25 VDD2.t7 7.25608
R636 VDD2.n23 VDD2.t8 7.25608
R637 VDD2.n23 VDD2.t2 7.25608
R638 VDD2.n49 VDD2.n27 4.26717
R639 VDD2.n22 VDD2.n0 4.26717
R640 VDD2.n34 VDD2.n32 3.73474
R641 VDD2.n7 VDD2.n5 3.73474
R642 VDD2.n47 VDD2.n46 3.49141
R643 VDD2.n20 VDD2.n19 3.49141
R644 VDD2.n52 VDD2.n50 2.92291
R645 VDD2.n43 VDD2.n29 2.71565
R646 VDD2.n16 VDD2.n2 2.71565
R647 VDD2.n42 VDD2.n31 1.93989
R648 VDD2.n15 VDD2.n4 1.93989
R649 VDD2.n39 VDD2.n38 1.16414
R650 VDD2.n12 VDD2.n11 1.16414
R651 VDD2 VDD2.n52 0.789293
R652 VDD2.n26 VDD2.n24 0.675757
R653 VDD2.n35 VDD2.n33 0.388379
R654 VDD2.n8 VDD2.n6 0.388379
R655 VDD2.n48 VDD2.n28 0.155672
R656 VDD2.n41 VDD2.n28 0.155672
R657 VDD2.n41 VDD2.n40 0.155672
R658 VDD2.n40 VDD2.n32 0.155672
R659 VDD2.n13 VDD2.n5 0.155672
R660 VDD2.n14 VDD2.n13 0.155672
R661 VDD2.n14 VDD2.n1 0.155672
R662 VDD2.n21 VDD2.n1 0.155672
R663 B.n578 B.n577 585
R664 B.n579 B.n64 585
R665 B.n581 B.n580 585
R666 B.n582 B.n63 585
R667 B.n584 B.n583 585
R668 B.n585 B.n62 585
R669 B.n587 B.n586 585
R670 B.n588 B.n61 585
R671 B.n590 B.n589 585
R672 B.n591 B.n60 585
R673 B.n593 B.n592 585
R674 B.n594 B.n59 585
R675 B.n596 B.n595 585
R676 B.n597 B.n58 585
R677 B.n599 B.n598 585
R678 B.n600 B.n57 585
R679 B.n602 B.n601 585
R680 B.n603 B.n56 585
R681 B.n605 B.n604 585
R682 B.n606 B.n53 585
R683 B.n609 B.n608 585
R684 B.n610 B.n52 585
R685 B.n612 B.n611 585
R686 B.n613 B.n51 585
R687 B.n615 B.n614 585
R688 B.n616 B.n50 585
R689 B.n618 B.n617 585
R690 B.n619 B.n49 585
R691 B.n621 B.n620 585
R692 B.n623 B.n622 585
R693 B.n624 B.n45 585
R694 B.n626 B.n625 585
R695 B.n627 B.n44 585
R696 B.n629 B.n628 585
R697 B.n630 B.n43 585
R698 B.n632 B.n631 585
R699 B.n633 B.n42 585
R700 B.n635 B.n634 585
R701 B.n636 B.n41 585
R702 B.n638 B.n637 585
R703 B.n639 B.n40 585
R704 B.n641 B.n640 585
R705 B.n642 B.n39 585
R706 B.n644 B.n643 585
R707 B.n645 B.n38 585
R708 B.n647 B.n646 585
R709 B.n648 B.n37 585
R710 B.n650 B.n649 585
R711 B.n651 B.n36 585
R712 B.n576 B.n65 585
R713 B.n575 B.n574 585
R714 B.n573 B.n66 585
R715 B.n572 B.n571 585
R716 B.n570 B.n67 585
R717 B.n569 B.n568 585
R718 B.n567 B.n68 585
R719 B.n566 B.n565 585
R720 B.n564 B.n69 585
R721 B.n563 B.n562 585
R722 B.n561 B.n70 585
R723 B.n560 B.n559 585
R724 B.n558 B.n71 585
R725 B.n557 B.n556 585
R726 B.n555 B.n72 585
R727 B.n554 B.n553 585
R728 B.n552 B.n73 585
R729 B.n551 B.n550 585
R730 B.n549 B.n74 585
R731 B.n548 B.n547 585
R732 B.n546 B.n75 585
R733 B.n545 B.n544 585
R734 B.n543 B.n76 585
R735 B.n542 B.n541 585
R736 B.n540 B.n77 585
R737 B.n539 B.n538 585
R738 B.n537 B.n78 585
R739 B.n536 B.n535 585
R740 B.n534 B.n79 585
R741 B.n533 B.n532 585
R742 B.n531 B.n80 585
R743 B.n530 B.n529 585
R744 B.n528 B.n81 585
R745 B.n527 B.n526 585
R746 B.n525 B.n82 585
R747 B.n524 B.n523 585
R748 B.n522 B.n83 585
R749 B.n521 B.n520 585
R750 B.n519 B.n84 585
R751 B.n518 B.n517 585
R752 B.n516 B.n85 585
R753 B.n515 B.n514 585
R754 B.n513 B.n86 585
R755 B.n512 B.n511 585
R756 B.n510 B.n87 585
R757 B.n509 B.n508 585
R758 B.n507 B.n88 585
R759 B.n506 B.n505 585
R760 B.n504 B.n89 585
R761 B.n503 B.n502 585
R762 B.n501 B.n90 585
R763 B.n500 B.n499 585
R764 B.n498 B.n91 585
R765 B.n497 B.n496 585
R766 B.n495 B.n92 585
R767 B.n494 B.n493 585
R768 B.n492 B.n93 585
R769 B.n491 B.n490 585
R770 B.n489 B.n94 585
R771 B.n488 B.n487 585
R772 B.n486 B.n95 585
R773 B.n485 B.n484 585
R774 B.n483 B.n96 585
R775 B.n482 B.n481 585
R776 B.n480 B.n97 585
R777 B.n479 B.n478 585
R778 B.n477 B.n98 585
R779 B.n476 B.n475 585
R780 B.n474 B.n99 585
R781 B.n473 B.n472 585
R782 B.n471 B.n100 585
R783 B.n470 B.n469 585
R784 B.n468 B.n101 585
R785 B.n467 B.n466 585
R786 B.n465 B.n102 585
R787 B.n464 B.n463 585
R788 B.n462 B.n103 585
R789 B.n461 B.n460 585
R790 B.n459 B.n104 585
R791 B.n458 B.n457 585
R792 B.n456 B.n105 585
R793 B.n455 B.n454 585
R794 B.n453 B.n106 585
R795 B.n452 B.n451 585
R796 B.n450 B.n107 585
R797 B.n449 B.n448 585
R798 B.n447 B.n108 585
R799 B.n446 B.n445 585
R800 B.n444 B.n109 585
R801 B.n443 B.n442 585
R802 B.n441 B.n110 585
R803 B.n440 B.n439 585
R804 B.n438 B.n111 585
R805 B.n437 B.n436 585
R806 B.n435 B.n112 585
R807 B.n434 B.n433 585
R808 B.n432 B.n113 585
R809 B.n431 B.n430 585
R810 B.n429 B.n114 585
R811 B.n428 B.n427 585
R812 B.n426 B.n115 585
R813 B.n425 B.n424 585
R814 B.n423 B.n116 585
R815 B.n422 B.n421 585
R816 B.n420 B.n117 585
R817 B.n419 B.n418 585
R818 B.n417 B.n118 585
R819 B.n416 B.n415 585
R820 B.n414 B.n119 585
R821 B.n413 B.n412 585
R822 B.n411 B.n120 585
R823 B.n410 B.n409 585
R824 B.n408 B.n121 585
R825 B.n407 B.n406 585
R826 B.n405 B.n122 585
R827 B.n404 B.n403 585
R828 B.n402 B.n123 585
R829 B.n401 B.n400 585
R830 B.n399 B.n124 585
R831 B.n398 B.n397 585
R832 B.n396 B.n125 585
R833 B.n395 B.n394 585
R834 B.n393 B.n126 585
R835 B.n392 B.n391 585
R836 B.n390 B.n127 585
R837 B.n389 B.n388 585
R838 B.n387 B.n128 585
R839 B.n386 B.n385 585
R840 B.n384 B.n129 585
R841 B.n383 B.n382 585
R842 B.n381 B.n130 585
R843 B.n380 B.n379 585
R844 B.n378 B.n131 585
R845 B.n377 B.n376 585
R846 B.n375 B.n132 585
R847 B.n374 B.n373 585
R848 B.n372 B.n133 585
R849 B.n297 B.n162 585
R850 B.n299 B.n298 585
R851 B.n300 B.n161 585
R852 B.n302 B.n301 585
R853 B.n303 B.n160 585
R854 B.n305 B.n304 585
R855 B.n306 B.n159 585
R856 B.n308 B.n307 585
R857 B.n309 B.n158 585
R858 B.n311 B.n310 585
R859 B.n312 B.n157 585
R860 B.n314 B.n313 585
R861 B.n315 B.n156 585
R862 B.n317 B.n316 585
R863 B.n318 B.n155 585
R864 B.n320 B.n319 585
R865 B.n321 B.n154 585
R866 B.n323 B.n322 585
R867 B.n324 B.n153 585
R868 B.n326 B.n325 585
R869 B.n328 B.n327 585
R870 B.n329 B.n149 585
R871 B.n331 B.n330 585
R872 B.n332 B.n148 585
R873 B.n334 B.n333 585
R874 B.n335 B.n147 585
R875 B.n337 B.n336 585
R876 B.n338 B.n146 585
R877 B.n340 B.n339 585
R878 B.n342 B.n143 585
R879 B.n344 B.n343 585
R880 B.n345 B.n142 585
R881 B.n347 B.n346 585
R882 B.n348 B.n141 585
R883 B.n350 B.n349 585
R884 B.n351 B.n140 585
R885 B.n353 B.n352 585
R886 B.n354 B.n139 585
R887 B.n356 B.n355 585
R888 B.n357 B.n138 585
R889 B.n359 B.n358 585
R890 B.n360 B.n137 585
R891 B.n362 B.n361 585
R892 B.n363 B.n136 585
R893 B.n365 B.n364 585
R894 B.n366 B.n135 585
R895 B.n368 B.n367 585
R896 B.n369 B.n134 585
R897 B.n371 B.n370 585
R898 B.n296 B.n295 585
R899 B.n294 B.n163 585
R900 B.n293 B.n292 585
R901 B.n291 B.n164 585
R902 B.n290 B.n289 585
R903 B.n288 B.n165 585
R904 B.n287 B.n286 585
R905 B.n285 B.n166 585
R906 B.n284 B.n283 585
R907 B.n282 B.n167 585
R908 B.n281 B.n280 585
R909 B.n279 B.n168 585
R910 B.n278 B.n277 585
R911 B.n276 B.n169 585
R912 B.n275 B.n274 585
R913 B.n273 B.n170 585
R914 B.n272 B.n271 585
R915 B.n270 B.n171 585
R916 B.n269 B.n268 585
R917 B.n267 B.n172 585
R918 B.n266 B.n265 585
R919 B.n264 B.n173 585
R920 B.n263 B.n262 585
R921 B.n261 B.n174 585
R922 B.n260 B.n259 585
R923 B.n258 B.n175 585
R924 B.n257 B.n256 585
R925 B.n255 B.n176 585
R926 B.n254 B.n253 585
R927 B.n252 B.n177 585
R928 B.n251 B.n250 585
R929 B.n249 B.n178 585
R930 B.n248 B.n247 585
R931 B.n246 B.n179 585
R932 B.n245 B.n244 585
R933 B.n243 B.n180 585
R934 B.n242 B.n241 585
R935 B.n240 B.n181 585
R936 B.n239 B.n238 585
R937 B.n237 B.n182 585
R938 B.n236 B.n235 585
R939 B.n234 B.n183 585
R940 B.n233 B.n232 585
R941 B.n231 B.n184 585
R942 B.n230 B.n229 585
R943 B.n228 B.n185 585
R944 B.n227 B.n226 585
R945 B.n225 B.n186 585
R946 B.n224 B.n223 585
R947 B.n222 B.n187 585
R948 B.n221 B.n220 585
R949 B.n219 B.n188 585
R950 B.n218 B.n217 585
R951 B.n216 B.n189 585
R952 B.n215 B.n214 585
R953 B.n213 B.n190 585
R954 B.n212 B.n211 585
R955 B.n210 B.n191 585
R956 B.n209 B.n208 585
R957 B.n207 B.n192 585
R958 B.n206 B.n205 585
R959 B.n204 B.n193 585
R960 B.n203 B.n202 585
R961 B.n201 B.n194 585
R962 B.n200 B.n199 585
R963 B.n198 B.n195 585
R964 B.n197 B.n196 585
R965 B.n2 B.n0 585
R966 B.n753 B.n1 585
R967 B.n752 B.n751 585
R968 B.n750 B.n3 585
R969 B.n749 B.n748 585
R970 B.n747 B.n4 585
R971 B.n746 B.n745 585
R972 B.n744 B.n5 585
R973 B.n743 B.n742 585
R974 B.n741 B.n6 585
R975 B.n740 B.n739 585
R976 B.n738 B.n7 585
R977 B.n737 B.n736 585
R978 B.n735 B.n8 585
R979 B.n734 B.n733 585
R980 B.n732 B.n9 585
R981 B.n731 B.n730 585
R982 B.n729 B.n10 585
R983 B.n728 B.n727 585
R984 B.n726 B.n11 585
R985 B.n725 B.n724 585
R986 B.n723 B.n12 585
R987 B.n722 B.n721 585
R988 B.n720 B.n13 585
R989 B.n719 B.n718 585
R990 B.n717 B.n14 585
R991 B.n716 B.n715 585
R992 B.n714 B.n15 585
R993 B.n713 B.n712 585
R994 B.n711 B.n16 585
R995 B.n710 B.n709 585
R996 B.n708 B.n17 585
R997 B.n707 B.n706 585
R998 B.n705 B.n18 585
R999 B.n704 B.n703 585
R1000 B.n702 B.n19 585
R1001 B.n701 B.n700 585
R1002 B.n699 B.n20 585
R1003 B.n698 B.n697 585
R1004 B.n696 B.n21 585
R1005 B.n695 B.n694 585
R1006 B.n693 B.n22 585
R1007 B.n692 B.n691 585
R1008 B.n690 B.n23 585
R1009 B.n689 B.n688 585
R1010 B.n687 B.n24 585
R1011 B.n686 B.n685 585
R1012 B.n684 B.n25 585
R1013 B.n683 B.n682 585
R1014 B.n681 B.n26 585
R1015 B.n680 B.n679 585
R1016 B.n678 B.n27 585
R1017 B.n677 B.n676 585
R1018 B.n675 B.n28 585
R1019 B.n674 B.n673 585
R1020 B.n672 B.n29 585
R1021 B.n671 B.n670 585
R1022 B.n669 B.n30 585
R1023 B.n668 B.n667 585
R1024 B.n666 B.n31 585
R1025 B.n665 B.n664 585
R1026 B.n663 B.n32 585
R1027 B.n662 B.n661 585
R1028 B.n660 B.n33 585
R1029 B.n659 B.n658 585
R1030 B.n657 B.n34 585
R1031 B.n656 B.n655 585
R1032 B.n654 B.n35 585
R1033 B.n653 B.n652 585
R1034 B.n755 B.n754 585
R1035 B.n297 B.n296 454.062
R1036 B.n652 B.n651 454.062
R1037 B.n370 B.n133 454.062
R1038 B.n578 B.n65 454.062
R1039 B.n144 B.t5 307.762
R1040 B.n54 B.t7 307.762
R1041 B.n150 B.t2 307.762
R1042 B.n46 B.t10 307.762
R1043 B.n144 B.t3 243.934
R1044 B.n150 B.t0 243.934
R1045 B.n46 B.t9 243.934
R1046 B.n54 B.t6 243.934
R1047 B.n145 B.t4 242.018
R1048 B.n55 B.t8 242.018
R1049 B.n151 B.t1 242.018
R1050 B.n47 B.t11 242.018
R1051 B.n296 B.n163 163.367
R1052 B.n292 B.n163 163.367
R1053 B.n292 B.n291 163.367
R1054 B.n291 B.n290 163.367
R1055 B.n290 B.n165 163.367
R1056 B.n286 B.n165 163.367
R1057 B.n286 B.n285 163.367
R1058 B.n285 B.n284 163.367
R1059 B.n284 B.n167 163.367
R1060 B.n280 B.n167 163.367
R1061 B.n280 B.n279 163.367
R1062 B.n279 B.n278 163.367
R1063 B.n278 B.n169 163.367
R1064 B.n274 B.n169 163.367
R1065 B.n274 B.n273 163.367
R1066 B.n273 B.n272 163.367
R1067 B.n272 B.n171 163.367
R1068 B.n268 B.n171 163.367
R1069 B.n268 B.n267 163.367
R1070 B.n267 B.n266 163.367
R1071 B.n266 B.n173 163.367
R1072 B.n262 B.n173 163.367
R1073 B.n262 B.n261 163.367
R1074 B.n261 B.n260 163.367
R1075 B.n260 B.n175 163.367
R1076 B.n256 B.n175 163.367
R1077 B.n256 B.n255 163.367
R1078 B.n255 B.n254 163.367
R1079 B.n254 B.n177 163.367
R1080 B.n250 B.n177 163.367
R1081 B.n250 B.n249 163.367
R1082 B.n249 B.n248 163.367
R1083 B.n248 B.n179 163.367
R1084 B.n244 B.n179 163.367
R1085 B.n244 B.n243 163.367
R1086 B.n243 B.n242 163.367
R1087 B.n242 B.n181 163.367
R1088 B.n238 B.n181 163.367
R1089 B.n238 B.n237 163.367
R1090 B.n237 B.n236 163.367
R1091 B.n236 B.n183 163.367
R1092 B.n232 B.n183 163.367
R1093 B.n232 B.n231 163.367
R1094 B.n231 B.n230 163.367
R1095 B.n230 B.n185 163.367
R1096 B.n226 B.n185 163.367
R1097 B.n226 B.n225 163.367
R1098 B.n225 B.n224 163.367
R1099 B.n224 B.n187 163.367
R1100 B.n220 B.n187 163.367
R1101 B.n220 B.n219 163.367
R1102 B.n219 B.n218 163.367
R1103 B.n218 B.n189 163.367
R1104 B.n214 B.n189 163.367
R1105 B.n214 B.n213 163.367
R1106 B.n213 B.n212 163.367
R1107 B.n212 B.n191 163.367
R1108 B.n208 B.n191 163.367
R1109 B.n208 B.n207 163.367
R1110 B.n207 B.n206 163.367
R1111 B.n206 B.n193 163.367
R1112 B.n202 B.n193 163.367
R1113 B.n202 B.n201 163.367
R1114 B.n201 B.n200 163.367
R1115 B.n200 B.n195 163.367
R1116 B.n196 B.n195 163.367
R1117 B.n196 B.n2 163.367
R1118 B.n754 B.n2 163.367
R1119 B.n754 B.n753 163.367
R1120 B.n753 B.n752 163.367
R1121 B.n752 B.n3 163.367
R1122 B.n748 B.n3 163.367
R1123 B.n748 B.n747 163.367
R1124 B.n747 B.n746 163.367
R1125 B.n746 B.n5 163.367
R1126 B.n742 B.n5 163.367
R1127 B.n742 B.n741 163.367
R1128 B.n741 B.n740 163.367
R1129 B.n740 B.n7 163.367
R1130 B.n736 B.n7 163.367
R1131 B.n736 B.n735 163.367
R1132 B.n735 B.n734 163.367
R1133 B.n734 B.n9 163.367
R1134 B.n730 B.n9 163.367
R1135 B.n730 B.n729 163.367
R1136 B.n729 B.n728 163.367
R1137 B.n728 B.n11 163.367
R1138 B.n724 B.n11 163.367
R1139 B.n724 B.n723 163.367
R1140 B.n723 B.n722 163.367
R1141 B.n722 B.n13 163.367
R1142 B.n718 B.n13 163.367
R1143 B.n718 B.n717 163.367
R1144 B.n717 B.n716 163.367
R1145 B.n716 B.n15 163.367
R1146 B.n712 B.n15 163.367
R1147 B.n712 B.n711 163.367
R1148 B.n711 B.n710 163.367
R1149 B.n710 B.n17 163.367
R1150 B.n706 B.n17 163.367
R1151 B.n706 B.n705 163.367
R1152 B.n705 B.n704 163.367
R1153 B.n704 B.n19 163.367
R1154 B.n700 B.n19 163.367
R1155 B.n700 B.n699 163.367
R1156 B.n699 B.n698 163.367
R1157 B.n698 B.n21 163.367
R1158 B.n694 B.n21 163.367
R1159 B.n694 B.n693 163.367
R1160 B.n693 B.n692 163.367
R1161 B.n692 B.n23 163.367
R1162 B.n688 B.n23 163.367
R1163 B.n688 B.n687 163.367
R1164 B.n687 B.n686 163.367
R1165 B.n686 B.n25 163.367
R1166 B.n682 B.n25 163.367
R1167 B.n682 B.n681 163.367
R1168 B.n681 B.n680 163.367
R1169 B.n680 B.n27 163.367
R1170 B.n676 B.n27 163.367
R1171 B.n676 B.n675 163.367
R1172 B.n675 B.n674 163.367
R1173 B.n674 B.n29 163.367
R1174 B.n670 B.n29 163.367
R1175 B.n670 B.n669 163.367
R1176 B.n669 B.n668 163.367
R1177 B.n668 B.n31 163.367
R1178 B.n664 B.n31 163.367
R1179 B.n664 B.n663 163.367
R1180 B.n663 B.n662 163.367
R1181 B.n662 B.n33 163.367
R1182 B.n658 B.n33 163.367
R1183 B.n658 B.n657 163.367
R1184 B.n657 B.n656 163.367
R1185 B.n656 B.n35 163.367
R1186 B.n652 B.n35 163.367
R1187 B.n298 B.n297 163.367
R1188 B.n298 B.n161 163.367
R1189 B.n302 B.n161 163.367
R1190 B.n303 B.n302 163.367
R1191 B.n304 B.n303 163.367
R1192 B.n304 B.n159 163.367
R1193 B.n308 B.n159 163.367
R1194 B.n309 B.n308 163.367
R1195 B.n310 B.n309 163.367
R1196 B.n310 B.n157 163.367
R1197 B.n314 B.n157 163.367
R1198 B.n315 B.n314 163.367
R1199 B.n316 B.n315 163.367
R1200 B.n316 B.n155 163.367
R1201 B.n320 B.n155 163.367
R1202 B.n321 B.n320 163.367
R1203 B.n322 B.n321 163.367
R1204 B.n322 B.n153 163.367
R1205 B.n326 B.n153 163.367
R1206 B.n327 B.n326 163.367
R1207 B.n327 B.n149 163.367
R1208 B.n331 B.n149 163.367
R1209 B.n332 B.n331 163.367
R1210 B.n333 B.n332 163.367
R1211 B.n333 B.n147 163.367
R1212 B.n337 B.n147 163.367
R1213 B.n338 B.n337 163.367
R1214 B.n339 B.n338 163.367
R1215 B.n339 B.n143 163.367
R1216 B.n344 B.n143 163.367
R1217 B.n345 B.n344 163.367
R1218 B.n346 B.n345 163.367
R1219 B.n346 B.n141 163.367
R1220 B.n350 B.n141 163.367
R1221 B.n351 B.n350 163.367
R1222 B.n352 B.n351 163.367
R1223 B.n352 B.n139 163.367
R1224 B.n356 B.n139 163.367
R1225 B.n357 B.n356 163.367
R1226 B.n358 B.n357 163.367
R1227 B.n358 B.n137 163.367
R1228 B.n362 B.n137 163.367
R1229 B.n363 B.n362 163.367
R1230 B.n364 B.n363 163.367
R1231 B.n364 B.n135 163.367
R1232 B.n368 B.n135 163.367
R1233 B.n369 B.n368 163.367
R1234 B.n370 B.n369 163.367
R1235 B.n374 B.n133 163.367
R1236 B.n375 B.n374 163.367
R1237 B.n376 B.n375 163.367
R1238 B.n376 B.n131 163.367
R1239 B.n380 B.n131 163.367
R1240 B.n381 B.n380 163.367
R1241 B.n382 B.n381 163.367
R1242 B.n382 B.n129 163.367
R1243 B.n386 B.n129 163.367
R1244 B.n387 B.n386 163.367
R1245 B.n388 B.n387 163.367
R1246 B.n388 B.n127 163.367
R1247 B.n392 B.n127 163.367
R1248 B.n393 B.n392 163.367
R1249 B.n394 B.n393 163.367
R1250 B.n394 B.n125 163.367
R1251 B.n398 B.n125 163.367
R1252 B.n399 B.n398 163.367
R1253 B.n400 B.n399 163.367
R1254 B.n400 B.n123 163.367
R1255 B.n404 B.n123 163.367
R1256 B.n405 B.n404 163.367
R1257 B.n406 B.n405 163.367
R1258 B.n406 B.n121 163.367
R1259 B.n410 B.n121 163.367
R1260 B.n411 B.n410 163.367
R1261 B.n412 B.n411 163.367
R1262 B.n412 B.n119 163.367
R1263 B.n416 B.n119 163.367
R1264 B.n417 B.n416 163.367
R1265 B.n418 B.n417 163.367
R1266 B.n418 B.n117 163.367
R1267 B.n422 B.n117 163.367
R1268 B.n423 B.n422 163.367
R1269 B.n424 B.n423 163.367
R1270 B.n424 B.n115 163.367
R1271 B.n428 B.n115 163.367
R1272 B.n429 B.n428 163.367
R1273 B.n430 B.n429 163.367
R1274 B.n430 B.n113 163.367
R1275 B.n434 B.n113 163.367
R1276 B.n435 B.n434 163.367
R1277 B.n436 B.n435 163.367
R1278 B.n436 B.n111 163.367
R1279 B.n440 B.n111 163.367
R1280 B.n441 B.n440 163.367
R1281 B.n442 B.n441 163.367
R1282 B.n442 B.n109 163.367
R1283 B.n446 B.n109 163.367
R1284 B.n447 B.n446 163.367
R1285 B.n448 B.n447 163.367
R1286 B.n448 B.n107 163.367
R1287 B.n452 B.n107 163.367
R1288 B.n453 B.n452 163.367
R1289 B.n454 B.n453 163.367
R1290 B.n454 B.n105 163.367
R1291 B.n458 B.n105 163.367
R1292 B.n459 B.n458 163.367
R1293 B.n460 B.n459 163.367
R1294 B.n460 B.n103 163.367
R1295 B.n464 B.n103 163.367
R1296 B.n465 B.n464 163.367
R1297 B.n466 B.n465 163.367
R1298 B.n466 B.n101 163.367
R1299 B.n470 B.n101 163.367
R1300 B.n471 B.n470 163.367
R1301 B.n472 B.n471 163.367
R1302 B.n472 B.n99 163.367
R1303 B.n476 B.n99 163.367
R1304 B.n477 B.n476 163.367
R1305 B.n478 B.n477 163.367
R1306 B.n478 B.n97 163.367
R1307 B.n482 B.n97 163.367
R1308 B.n483 B.n482 163.367
R1309 B.n484 B.n483 163.367
R1310 B.n484 B.n95 163.367
R1311 B.n488 B.n95 163.367
R1312 B.n489 B.n488 163.367
R1313 B.n490 B.n489 163.367
R1314 B.n490 B.n93 163.367
R1315 B.n494 B.n93 163.367
R1316 B.n495 B.n494 163.367
R1317 B.n496 B.n495 163.367
R1318 B.n496 B.n91 163.367
R1319 B.n500 B.n91 163.367
R1320 B.n501 B.n500 163.367
R1321 B.n502 B.n501 163.367
R1322 B.n502 B.n89 163.367
R1323 B.n506 B.n89 163.367
R1324 B.n507 B.n506 163.367
R1325 B.n508 B.n507 163.367
R1326 B.n508 B.n87 163.367
R1327 B.n512 B.n87 163.367
R1328 B.n513 B.n512 163.367
R1329 B.n514 B.n513 163.367
R1330 B.n514 B.n85 163.367
R1331 B.n518 B.n85 163.367
R1332 B.n519 B.n518 163.367
R1333 B.n520 B.n519 163.367
R1334 B.n520 B.n83 163.367
R1335 B.n524 B.n83 163.367
R1336 B.n525 B.n524 163.367
R1337 B.n526 B.n525 163.367
R1338 B.n526 B.n81 163.367
R1339 B.n530 B.n81 163.367
R1340 B.n531 B.n530 163.367
R1341 B.n532 B.n531 163.367
R1342 B.n532 B.n79 163.367
R1343 B.n536 B.n79 163.367
R1344 B.n537 B.n536 163.367
R1345 B.n538 B.n537 163.367
R1346 B.n538 B.n77 163.367
R1347 B.n542 B.n77 163.367
R1348 B.n543 B.n542 163.367
R1349 B.n544 B.n543 163.367
R1350 B.n544 B.n75 163.367
R1351 B.n548 B.n75 163.367
R1352 B.n549 B.n548 163.367
R1353 B.n550 B.n549 163.367
R1354 B.n550 B.n73 163.367
R1355 B.n554 B.n73 163.367
R1356 B.n555 B.n554 163.367
R1357 B.n556 B.n555 163.367
R1358 B.n556 B.n71 163.367
R1359 B.n560 B.n71 163.367
R1360 B.n561 B.n560 163.367
R1361 B.n562 B.n561 163.367
R1362 B.n562 B.n69 163.367
R1363 B.n566 B.n69 163.367
R1364 B.n567 B.n566 163.367
R1365 B.n568 B.n567 163.367
R1366 B.n568 B.n67 163.367
R1367 B.n572 B.n67 163.367
R1368 B.n573 B.n572 163.367
R1369 B.n574 B.n573 163.367
R1370 B.n574 B.n65 163.367
R1371 B.n651 B.n650 163.367
R1372 B.n650 B.n37 163.367
R1373 B.n646 B.n37 163.367
R1374 B.n646 B.n645 163.367
R1375 B.n645 B.n644 163.367
R1376 B.n644 B.n39 163.367
R1377 B.n640 B.n39 163.367
R1378 B.n640 B.n639 163.367
R1379 B.n639 B.n638 163.367
R1380 B.n638 B.n41 163.367
R1381 B.n634 B.n41 163.367
R1382 B.n634 B.n633 163.367
R1383 B.n633 B.n632 163.367
R1384 B.n632 B.n43 163.367
R1385 B.n628 B.n43 163.367
R1386 B.n628 B.n627 163.367
R1387 B.n627 B.n626 163.367
R1388 B.n626 B.n45 163.367
R1389 B.n622 B.n45 163.367
R1390 B.n622 B.n621 163.367
R1391 B.n621 B.n49 163.367
R1392 B.n617 B.n49 163.367
R1393 B.n617 B.n616 163.367
R1394 B.n616 B.n615 163.367
R1395 B.n615 B.n51 163.367
R1396 B.n611 B.n51 163.367
R1397 B.n611 B.n610 163.367
R1398 B.n610 B.n609 163.367
R1399 B.n609 B.n53 163.367
R1400 B.n604 B.n53 163.367
R1401 B.n604 B.n603 163.367
R1402 B.n603 B.n602 163.367
R1403 B.n602 B.n57 163.367
R1404 B.n598 B.n57 163.367
R1405 B.n598 B.n597 163.367
R1406 B.n597 B.n596 163.367
R1407 B.n596 B.n59 163.367
R1408 B.n592 B.n59 163.367
R1409 B.n592 B.n591 163.367
R1410 B.n591 B.n590 163.367
R1411 B.n590 B.n61 163.367
R1412 B.n586 B.n61 163.367
R1413 B.n586 B.n585 163.367
R1414 B.n585 B.n584 163.367
R1415 B.n584 B.n63 163.367
R1416 B.n580 B.n63 163.367
R1417 B.n580 B.n579 163.367
R1418 B.n579 B.n578 163.367
R1419 B.n145 B.n144 65.746
R1420 B.n151 B.n150 65.746
R1421 B.n47 B.n46 65.746
R1422 B.n55 B.n54 65.746
R1423 B.n341 B.n145 59.5399
R1424 B.n152 B.n151 59.5399
R1425 B.n48 B.n47 59.5399
R1426 B.n607 B.n55 59.5399
R1427 B.n577 B.n576 29.5029
R1428 B.n653 B.n36 29.5029
R1429 B.n372 B.n371 29.5029
R1430 B.n295 B.n162 29.5029
R1431 B B.n755 18.0485
R1432 B.n649 B.n36 10.6151
R1433 B.n649 B.n648 10.6151
R1434 B.n648 B.n647 10.6151
R1435 B.n647 B.n38 10.6151
R1436 B.n643 B.n38 10.6151
R1437 B.n643 B.n642 10.6151
R1438 B.n642 B.n641 10.6151
R1439 B.n641 B.n40 10.6151
R1440 B.n637 B.n40 10.6151
R1441 B.n637 B.n636 10.6151
R1442 B.n636 B.n635 10.6151
R1443 B.n635 B.n42 10.6151
R1444 B.n631 B.n42 10.6151
R1445 B.n631 B.n630 10.6151
R1446 B.n630 B.n629 10.6151
R1447 B.n629 B.n44 10.6151
R1448 B.n625 B.n44 10.6151
R1449 B.n625 B.n624 10.6151
R1450 B.n624 B.n623 10.6151
R1451 B.n620 B.n619 10.6151
R1452 B.n619 B.n618 10.6151
R1453 B.n618 B.n50 10.6151
R1454 B.n614 B.n50 10.6151
R1455 B.n614 B.n613 10.6151
R1456 B.n613 B.n612 10.6151
R1457 B.n612 B.n52 10.6151
R1458 B.n608 B.n52 10.6151
R1459 B.n606 B.n605 10.6151
R1460 B.n605 B.n56 10.6151
R1461 B.n601 B.n56 10.6151
R1462 B.n601 B.n600 10.6151
R1463 B.n600 B.n599 10.6151
R1464 B.n599 B.n58 10.6151
R1465 B.n595 B.n58 10.6151
R1466 B.n595 B.n594 10.6151
R1467 B.n594 B.n593 10.6151
R1468 B.n593 B.n60 10.6151
R1469 B.n589 B.n60 10.6151
R1470 B.n589 B.n588 10.6151
R1471 B.n588 B.n587 10.6151
R1472 B.n587 B.n62 10.6151
R1473 B.n583 B.n62 10.6151
R1474 B.n583 B.n582 10.6151
R1475 B.n582 B.n581 10.6151
R1476 B.n581 B.n64 10.6151
R1477 B.n577 B.n64 10.6151
R1478 B.n373 B.n372 10.6151
R1479 B.n373 B.n132 10.6151
R1480 B.n377 B.n132 10.6151
R1481 B.n378 B.n377 10.6151
R1482 B.n379 B.n378 10.6151
R1483 B.n379 B.n130 10.6151
R1484 B.n383 B.n130 10.6151
R1485 B.n384 B.n383 10.6151
R1486 B.n385 B.n384 10.6151
R1487 B.n385 B.n128 10.6151
R1488 B.n389 B.n128 10.6151
R1489 B.n390 B.n389 10.6151
R1490 B.n391 B.n390 10.6151
R1491 B.n391 B.n126 10.6151
R1492 B.n395 B.n126 10.6151
R1493 B.n396 B.n395 10.6151
R1494 B.n397 B.n396 10.6151
R1495 B.n397 B.n124 10.6151
R1496 B.n401 B.n124 10.6151
R1497 B.n402 B.n401 10.6151
R1498 B.n403 B.n402 10.6151
R1499 B.n403 B.n122 10.6151
R1500 B.n407 B.n122 10.6151
R1501 B.n408 B.n407 10.6151
R1502 B.n409 B.n408 10.6151
R1503 B.n409 B.n120 10.6151
R1504 B.n413 B.n120 10.6151
R1505 B.n414 B.n413 10.6151
R1506 B.n415 B.n414 10.6151
R1507 B.n415 B.n118 10.6151
R1508 B.n419 B.n118 10.6151
R1509 B.n420 B.n419 10.6151
R1510 B.n421 B.n420 10.6151
R1511 B.n421 B.n116 10.6151
R1512 B.n425 B.n116 10.6151
R1513 B.n426 B.n425 10.6151
R1514 B.n427 B.n426 10.6151
R1515 B.n427 B.n114 10.6151
R1516 B.n431 B.n114 10.6151
R1517 B.n432 B.n431 10.6151
R1518 B.n433 B.n432 10.6151
R1519 B.n433 B.n112 10.6151
R1520 B.n437 B.n112 10.6151
R1521 B.n438 B.n437 10.6151
R1522 B.n439 B.n438 10.6151
R1523 B.n439 B.n110 10.6151
R1524 B.n443 B.n110 10.6151
R1525 B.n444 B.n443 10.6151
R1526 B.n445 B.n444 10.6151
R1527 B.n445 B.n108 10.6151
R1528 B.n449 B.n108 10.6151
R1529 B.n450 B.n449 10.6151
R1530 B.n451 B.n450 10.6151
R1531 B.n451 B.n106 10.6151
R1532 B.n455 B.n106 10.6151
R1533 B.n456 B.n455 10.6151
R1534 B.n457 B.n456 10.6151
R1535 B.n457 B.n104 10.6151
R1536 B.n461 B.n104 10.6151
R1537 B.n462 B.n461 10.6151
R1538 B.n463 B.n462 10.6151
R1539 B.n463 B.n102 10.6151
R1540 B.n467 B.n102 10.6151
R1541 B.n468 B.n467 10.6151
R1542 B.n469 B.n468 10.6151
R1543 B.n469 B.n100 10.6151
R1544 B.n473 B.n100 10.6151
R1545 B.n474 B.n473 10.6151
R1546 B.n475 B.n474 10.6151
R1547 B.n475 B.n98 10.6151
R1548 B.n479 B.n98 10.6151
R1549 B.n480 B.n479 10.6151
R1550 B.n481 B.n480 10.6151
R1551 B.n481 B.n96 10.6151
R1552 B.n485 B.n96 10.6151
R1553 B.n486 B.n485 10.6151
R1554 B.n487 B.n486 10.6151
R1555 B.n487 B.n94 10.6151
R1556 B.n491 B.n94 10.6151
R1557 B.n492 B.n491 10.6151
R1558 B.n493 B.n492 10.6151
R1559 B.n493 B.n92 10.6151
R1560 B.n497 B.n92 10.6151
R1561 B.n498 B.n497 10.6151
R1562 B.n499 B.n498 10.6151
R1563 B.n499 B.n90 10.6151
R1564 B.n503 B.n90 10.6151
R1565 B.n504 B.n503 10.6151
R1566 B.n505 B.n504 10.6151
R1567 B.n505 B.n88 10.6151
R1568 B.n509 B.n88 10.6151
R1569 B.n510 B.n509 10.6151
R1570 B.n511 B.n510 10.6151
R1571 B.n511 B.n86 10.6151
R1572 B.n515 B.n86 10.6151
R1573 B.n516 B.n515 10.6151
R1574 B.n517 B.n516 10.6151
R1575 B.n517 B.n84 10.6151
R1576 B.n521 B.n84 10.6151
R1577 B.n522 B.n521 10.6151
R1578 B.n523 B.n522 10.6151
R1579 B.n523 B.n82 10.6151
R1580 B.n527 B.n82 10.6151
R1581 B.n528 B.n527 10.6151
R1582 B.n529 B.n528 10.6151
R1583 B.n529 B.n80 10.6151
R1584 B.n533 B.n80 10.6151
R1585 B.n534 B.n533 10.6151
R1586 B.n535 B.n534 10.6151
R1587 B.n535 B.n78 10.6151
R1588 B.n539 B.n78 10.6151
R1589 B.n540 B.n539 10.6151
R1590 B.n541 B.n540 10.6151
R1591 B.n541 B.n76 10.6151
R1592 B.n545 B.n76 10.6151
R1593 B.n546 B.n545 10.6151
R1594 B.n547 B.n546 10.6151
R1595 B.n547 B.n74 10.6151
R1596 B.n551 B.n74 10.6151
R1597 B.n552 B.n551 10.6151
R1598 B.n553 B.n552 10.6151
R1599 B.n553 B.n72 10.6151
R1600 B.n557 B.n72 10.6151
R1601 B.n558 B.n557 10.6151
R1602 B.n559 B.n558 10.6151
R1603 B.n559 B.n70 10.6151
R1604 B.n563 B.n70 10.6151
R1605 B.n564 B.n563 10.6151
R1606 B.n565 B.n564 10.6151
R1607 B.n565 B.n68 10.6151
R1608 B.n569 B.n68 10.6151
R1609 B.n570 B.n569 10.6151
R1610 B.n571 B.n570 10.6151
R1611 B.n571 B.n66 10.6151
R1612 B.n575 B.n66 10.6151
R1613 B.n576 B.n575 10.6151
R1614 B.n299 B.n162 10.6151
R1615 B.n300 B.n299 10.6151
R1616 B.n301 B.n300 10.6151
R1617 B.n301 B.n160 10.6151
R1618 B.n305 B.n160 10.6151
R1619 B.n306 B.n305 10.6151
R1620 B.n307 B.n306 10.6151
R1621 B.n307 B.n158 10.6151
R1622 B.n311 B.n158 10.6151
R1623 B.n312 B.n311 10.6151
R1624 B.n313 B.n312 10.6151
R1625 B.n313 B.n156 10.6151
R1626 B.n317 B.n156 10.6151
R1627 B.n318 B.n317 10.6151
R1628 B.n319 B.n318 10.6151
R1629 B.n319 B.n154 10.6151
R1630 B.n323 B.n154 10.6151
R1631 B.n324 B.n323 10.6151
R1632 B.n325 B.n324 10.6151
R1633 B.n329 B.n328 10.6151
R1634 B.n330 B.n329 10.6151
R1635 B.n330 B.n148 10.6151
R1636 B.n334 B.n148 10.6151
R1637 B.n335 B.n334 10.6151
R1638 B.n336 B.n335 10.6151
R1639 B.n336 B.n146 10.6151
R1640 B.n340 B.n146 10.6151
R1641 B.n343 B.n342 10.6151
R1642 B.n343 B.n142 10.6151
R1643 B.n347 B.n142 10.6151
R1644 B.n348 B.n347 10.6151
R1645 B.n349 B.n348 10.6151
R1646 B.n349 B.n140 10.6151
R1647 B.n353 B.n140 10.6151
R1648 B.n354 B.n353 10.6151
R1649 B.n355 B.n354 10.6151
R1650 B.n355 B.n138 10.6151
R1651 B.n359 B.n138 10.6151
R1652 B.n360 B.n359 10.6151
R1653 B.n361 B.n360 10.6151
R1654 B.n361 B.n136 10.6151
R1655 B.n365 B.n136 10.6151
R1656 B.n366 B.n365 10.6151
R1657 B.n367 B.n366 10.6151
R1658 B.n367 B.n134 10.6151
R1659 B.n371 B.n134 10.6151
R1660 B.n295 B.n294 10.6151
R1661 B.n294 B.n293 10.6151
R1662 B.n293 B.n164 10.6151
R1663 B.n289 B.n164 10.6151
R1664 B.n289 B.n288 10.6151
R1665 B.n288 B.n287 10.6151
R1666 B.n287 B.n166 10.6151
R1667 B.n283 B.n166 10.6151
R1668 B.n283 B.n282 10.6151
R1669 B.n282 B.n281 10.6151
R1670 B.n281 B.n168 10.6151
R1671 B.n277 B.n168 10.6151
R1672 B.n277 B.n276 10.6151
R1673 B.n276 B.n275 10.6151
R1674 B.n275 B.n170 10.6151
R1675 B.n271 B.n170 10.6151
R1676 B.n271 B.n270 10.6151
R1677 B.n270 B.n269 10.6151
R1678 B.n269 B.n172 10.6151
R1679 B.n265 B.n172 10.6151
R1680 B.n265 B.n264 10.6151
R1681 B.n264 B.n263 10.6151
R1682 B.n263 B.n174 10.6151
R1683 B.n259 B.n174 10.6151
R1684 B.n259 B.n258 10.6151
R1685 B.n258 B.n257 10.6151
R1686 B.n257 B.n176 10.6151
R1687 B.n253 B.n176 10.6151
R1688 B.n253 B.n252 10.6151
R1689 B.n252 B.n251 10.6151
R1690 B.n251 B.n178 10.6151
R1691 B.n247 B.n178 10.6151
R1692 B.n247 B.n246 10.6151
R1693 B.n246 B.n245 10.6151
R1694 B.n245 B.n180 10.6151
R1695 B.n241 B.n180 10.6151
R1696 B.n241 B.n240 10.6151
R1697 B.n240 B.n239 10.6151
R1698 B.n239 B.n182 10.6151
R1699 B.n235 B.n182 10.6151
R1700 B.n235 B.n234 10.6151
R1701 B.n234 B.n233 10.6151
R1702 B.n233 B.n184 10.6151
R1703 B.n229 B.n184 10.6151
R1704 B.n229 B.n228 10.6151
R1705 B.n228 B.n227 10.6151
R1706 B.n227 B.n186 10.6151
R1707 B.n223 B.n186 10.6151
R1708 B.n223 B.n222 10.6151
R1709 B.n222 B.n221 10.6151
R1710 B.n221 B.n188 10.6151
R1711 B.n217 B.n188 10.6151
R1712 B.n217 B.n216 10.6151
R1713 B.n216 B.n215 10.6151
R1714 B.n215 B.n190 10.6151
R1715 B.n211 B.n190 10.6151
R1716 B.n211 B.n210 10.6151
R1717 B.n210 B.n209 10.6151
R1718 B.n209 B.n192 10.6151
R1719 B.n205 B.n192 10.6151
R1720 B.n205 B.n204 10.6151
R1721 B.n204 B.n203 10.6151
R1722 B.n203 B.n194 10.6151
R1723 B.n199 B.n194 10.6151
R1724 B.n199 B.n198 10.6151
R1725 B.n198 B.n197 10.6151
R1726 B.n197 B.n0 10.6151
R1727 B.n751 B.n1 10.6151
R1728 B.n751 B.n750 10.6151
R1729 B.n750 B.n749 10.6151
R1730 B.n749 B.n4 10.6151
R1731 B.n745 B.n4 10.6151
R1732 B.n745 B.n744 10.6151
R1733 B.n744 B.n743 10.6151
R1734 B.n743 B.n6 10.6151
R1735 B.n739 B.n6 10.6151
R1736 B.n739 B.n738 10.6151
R1737 B.n738 B.n737 10.6151
R1738 B.n737 B.n8 10.6151
R1739 B.n733 B.n8 10.6151
R1740 B.n733 B.n732 10.6151
R1741 B.n732 B.n731 10.6151
R1742 B.n731 B.n10 10.6151
R1743 B.n727 B.n10 10.6151
R1744 B.n727 B.n726 10.6151
R1745 B.n726 B.n725 10.6151
R1746 B.n725 B.n12 10.6151
R1747 B.n721 B.n12 10.6151
R1748 B.n721 B.n720 10.6151
R1749 B.n720 B.n719 10.6151
R1750 B.n719 B.n14 10.6151
R1751 B.n715 B.n14 10.6151
R1752 B.n715 B.n714 10.6151
R1753 B.n714 B.n713 10.6151
R1754 B.n713 B.n16 10.6151
R1755 B.n709 B.n16 10.6151
R1756 B.n709 B.n708 10.6151
R1757 B.n708 B.n707 10.6151
R1758 B.n707 B.n18 10.6151
R1759 B.n703 B.n18 10.6151
R1760 B.n703 B.n702 10.6151
R1761 B.n702 B.n701 10.6151
R1762 B.n701 B.n20 10.6151
R1763 B.n697 B.n20 10.6151
R1764 B.n697 B.n696 10.6151
R1765 B.n696 B.n695 10.6151
R1766 B.n695 B.n22 10.6151
R1767 B.n691 B.n22 10.6151
R1768 B.n691 B.n690 10.6151
R1769 B.n690 B.n689 10.6151
R1770 B.n689 B.n24 10.6151
R1771 B.n685 B.n24 10.6151
R1772 B.n685 B.n684 10.6151
R1773 B.n684 B.n683 10.6151
R1774 B.n683 B.n26 10.6151
R1775 B.n679 B.n26 10.6151
R1776 B.n679 B.n678 10.6151
R1777 B.n678 B.n677 10.6151
R1778 B.n677 B.n28 10.6151
R1779 B.n673 B.n28 10.6151
R1780 B.n673 B.n672 10.6151
R1781 B.n672 B.n671 10.6151
R1782 B.n671 B.n30 10.6151
R1783 B.n667 B.n30 10.6151
R1784 B.n667 B.n666 10.6151
R1785 B.n666 B.n665 10.6151
R1786 B.n665 B.n32 10.6151
R1787 B.n661 B.n32 10.6151
R1788 B.n661 B.n660 10.6151
R1789 B.n660 B.n659 10.6151
R1790 B.n659 B.n34 10.6151
R1791 B.n655 B.n34 10.6151
R1792 B.n655 B.n654 10.6151
R1793 B.n654 B.n653 10.6151
R1794 B.n620 B.n48 6.5566
R1795 B.n608 B.n607 6.5566
R1796 B.n328 B.n152 6.5566
R1797 B.n341 B.n340 6.5566
R1798 B.n623 B.n48 4.05904
R1799 B.n607 B.n606 4.05904
R1800 B.n325 B.n152 4.05904
R1801 B.n342 B.n341 4.05904
R1802 B.n755 B.n0 2.81026
R1803 B.n755 B.n1 2.81026
C0 VN B 1.36576f
C1 VN VDD1 0.158819f
C2 VTAIL VN 5.88735f
C3 B VDD2 2.19576f
C4 VDD1 VDD2 2.47335f
C5 VTAIL VDD2 7.40095f
C6 VN w_n5038_n1864# 10.794499f
C7 w_n5038_n1864# VDD2 2.61148f
C8 VDD1 B 2.05978f
C9 VTAIL B 2.14738f
C10 VTAIL VDD1 7.345f
C11 B w_n5038_n1864# 9.232889f
C12 VDD1 w_n5038_n1864# 2.44434f
C13 VTAIL w_n5038_n1864# 2.22867f
C14 VN VP 7.687109f
C15 VP VDD2 0.646784f
C16 B VP 2.47354f
C17 VDD1 VP 4.92425f
C18 VN VDD2 4.43982f
C19 VTAIL VP 5.90151f
C20 w_n5038_n1864# VP 11.4515f
C21 VDD2 VSUBS 2.253178f
C22 VDD1 VSUBS 1.98081f
C23 VTAIL VSUBS 0.693713f
C24 VN VSUBS 8.20449f
C25 VP VSUBS 4.202816f
C26 B VSUBS 4.977523f
C27 w_n5038_n1864# VSUBS 0.11795p
C28 B.n0 VSUBS 0.008179f
C29 B.n1 VSUBS 0.008179f
C30 B.n2 VSUBS 0.012934f
C31 B.n3 VSUBS 0.012934f
C32 B.n4 VSUBS 0.012934f
C33 B.n5 VSUBS 0.012934f
C34 B.n6 VSUBS 0.012934f
C35 B.n7 VSUBS 0.012934f
C36 B.n8 VSUBS 0.012934f
C37 B.n9 VSUBS 0.012934f
C38 B.n10 VSUBS 0.012934f
C39 B.n11 VSUBS 0.012934f
C40 B.n12 VSUBS 0.012934f
C41 B.n13 VSUBS 0.012934f
C42 B.n14 VSUBS 0.012934f
C43 B.n15 VSUBS 0.012934f
C44 B.n16 VSUBS 0.012934f
C45 B.n17 VSUBS 0.012934f
C46 B.n18 VSUBS 0.012934f
C47 B.n19 VSUBS 0.012934f
C48 B.n20 VSUBS 0.012934f
C49 B.n21 VSUBS 0.012934f
C50 B.n22 VSUBS 0.012934f
C51 B.n23 VSUBS 0.012934f
C52 B.n24 VSUBS 0.012934f
C53 B.n25 VSUBS 0.012934f
C54 B.n26 VSUBS 0.012934f
C55 B.n27 VSUBS 0.012934f
C56 B.n28 VSUBS 0.012934f
C57 B.n29 VSUBS 0.012934f
C58 B.n30 VSUBS 0.012934f
C59 B.n31 VSUBS 0.012934f
C60 B.n32 VSUBS 0.012934f
C61 B.n33 VSUBS 0.012934f
C62 B.n34 VSUBS 0.012934f
C63 B.n35 VSUBS 0.012934f
C64 B.n36 VSUBS 0.029352f
C65 B.n37 VSUBS 0.012934f
C66 B.n38 VSUBS 0.012934f
C67 B.n39 VSUBS 0.012934f
C68 B.n40 VSUBS 0.012934f
C69 B.n41 VSUBS 0.012934f
C70 B.n42 VSUBS 0.012934f
C71 B.n43 VSUBS 0.012934f
C72 B.n44 VSUBS 0.012934f
C73 B.n45 VSUBS 0.012934f
C74 B.t11 VSUBS 0.118989f
C75 B.t10 VSUBS 0.165763f
C76 B.t9 VSUBS 1.22085f
C77 B.n46 VSUBS 0.285308f
C78 B.n47 VSUBS 0.237402f
C79 B.n48 VSUBS 0.029967f
C80 B.n49 VSUBS 0.012934f
C81 B.n50 VSUBS 0.012934f
C82 B.n51 VSUBS 0.012934f
C83 B.n52 VSUBS 0.012934f
C84 B.n53 VSUBS 0.012934f
C85 B.t8 VSUBS 0.118992f
C86 B.t7 VSUBS 0.165765f
C87 B.t6 VSUBS 1.22085f
C88 B.n54 VSUBS 0.285306f
C89 B.n55 VSUBS 0.2374f
C90 B.n56 VSUBS 0.012934f
C91 B.n57 VSUBS 0.012934f
C92 B.n58 VSUBS 0.012934f
C93 B.n59 VSUBS 0.012934f
C94 B.n60 VSUBS 0.012934f
C95 B.n61 VSUBS 0.012934f
C96 B.n62 VSUBS 0.012934f
C97 B.n63 VSUBS 0.012934f
C98 B.n64 VSUBS 0.012934f
C99 B.n65 VSUBS 0.02733f
C100 B.n66 VSUBS 0.012934f
C101 B.n67 VSUBS 0.012934f
C102 B.n68 VSUBS 0.012934f
C103 B.n69 VSUBS 0.012934f
C104 B.n70 VSUBS 0.012934f
C105 B.n71 VSUBS 0.012934f
C106 B.n72 VSUBS 0.012934f
C107 B.n73 VSUBS 0.012934f
C108 B.n74 VSUBS 0.012934f
C109 B.n75 VSUBS 0.012934f
C110 B.n76 VSUBS 0.012934f
C111 B.n77 VSUBS 0.012934f
C112 B.n78 VSUBS 0.012934f
C113 B.n79 VSUBS 0.012934f
C114 B.n80 VSUBS 0.012934f
C115 B.n81 VSUBS 0.012934f
C116 B.n82 VSUBS 0.012934f
C117 B.n83 VSUBS 0.012934f
C118 B.n84 VSUBS 0.012934f
C119 B.n85 VSUBS 0.012934f
C120 B.n86 VSUBS 0.012934f
C121 B.n87 VSUBS 0.012934f
C122 B.n88 VSUBS 0.012934f
C123 B.n89 VSUBS 0.012934f
C124 B.n90 VSUBS 0.012934f
C125 B.n91 VSUBS 0.012934f
C126 B.n92 VSUBS 0.012934f
C127 B.n93 VSUBS 0.012934f
C128 B.n94 VSUBS 0.012934f
C129 B.n95 VSUBS 0.012934f
C130 B.n96 VSUBS 0.012934f
C131 B.n97 VSUBS 0.012934f
C132 B.n98 VSUBS 0.012934f
C133 B.n99 VSUBS 0.012934f
C134 B.n100 VSUBS 0.012934f
C135 B.n101 VSUBS 0.012934f
C136 B.n102 VSUBS 0.012934f
C137 B.n103 VSUBS 0.012934f
C138 B.n104 VSUBS 0.012934f
C139 B.n105 VSUBS 0.012934f
C140 B.n106 VSUBS 0.012934f
C141 B.n107 VSUBS 0.012934f
C142 B.n108 VSUBS 0.012934f
C143 B.n109 VSUBS 0.012934f
C144 B.n110 VSUBS 0.012934f
C145 B.n111 VSUBS 0.012934f
C146 B.n112 VSUBS 0.012934f
C147 B.n113 VSUBS 0.012934f
C148 B.n114 VSUBS 0.012934f
C149 B.n115 VSUBS 0.012934f
C150 B.n116 VSUBS 0.012934f
C151 B.n117 VSUBS 0.012934f
C152 B.n118 VSUBS 0.012934f
C153 B.n119 VSUBS 0.012934f
C154 B.n120 VSUBS 0.012934f
C155 B.n121 VSUBS 0.012934f
C156 B.n122 VSUBS 0.012934f
C157 B.n123 VSUBS 0.012934f
C158 B.n124 VSUBS 0.012934f
C159 B.n125 VSUBS 0.012934f
C160 B.n126 VSUBS 0.012934f
C161 B.n127 VSUBS 0.012934f
C162 B.n128 VSUBS 0.012934f
C163 B.n129 VSUBS 0.012934f
C164 B.n130 VSUBS 0.012934f
C165 B.n131 VSUBS 0.012934f
C166 B.n132 VSUBS 0.012934f
C167 B.n133 VSUBS 0.02733f
C168 B.n134 VSUBS 0.012934f
C169 B.n135 VSUBS 0.012934f
C170 B.n136 VSUBS 0.012934f
C171 B.n137 VSUBS 0.012934f
C172 B.n138 VSUBS 0.012934f
C173 B.n139 VSUBS 0.012934f
C174 B.n140 VSUBS 0.012934f
C175 B.n141 VSUBS 0.012934f
C176 B.n142 VSUBS 0.012934f
C177 B.n143 VSUBS 0.012934f
C178 B.t4 VSUBS 0.118992f
C179 B.t5 VSUBS 0.165765f
C180 B.t3 VSUBS 1.22085f
C181 B.n144 VSUBS 0.285306f
C182 B.n145 VSUBS 0.2374f
C183 B.n146 VSUBS 0.012934f
C184 B.n147 VSUBS 0.012934f
C185 B.n148 VSUBS 0.012934f
C186 B.n149 VSUBS 0.012934f
C187 B.t1 VSUBS 0.118989f
C188 B.t2 VSUBS 0.165763f
C189 B.t0 VSUBS 1.22085f
C190 B.n150 VSUBS 0.285308f
C191 B.n151 VSUBS 0.237402f
C192 B.n152 VSUBS 0.029967f
C193 B.n153 VSUBS 0.012934f
C194 B.n154 VSUBS 0.012934f
C195 B.n155 VSUBS 0.012934f
C196 B.n156 VSUBS 0.012934f
C197 B.n157 VSUBS 0.012934f
C198 B.n158 VSUBS 0.012934f
C199 B.n159 VSUBS 0.012934f
C200 B.n160 VSUBS 0.012934f
C201 B.n161 VSUBS 0.012934f
C202 B.n162 VSUBS 0.029352f
C203 B.n163 VSUBS 0.012934f
C204 B.n164 VSUBS 0.012934f
C205 B.n165 VSUBS 0.012934f
C206 B.n166 VSUBS 0.012934f
C207 B.n167 VSUBS 0.012934f
C208 B.n168 VSUBS 0.012934f
C209 B.n169 VSUBS 0.012934f
C210 B.n170 VSUBS 0.012934f
C211 B.n171 VSUBS 0.012934f
C212 B.n172 VSUBS 0.012934f
C213 B.n173 VSUBS 0.012934f
C214 B.n174 VSUBS 0.012934f
C215 B.n175 VSUBS 0.012934f
C216 B.n176 VSUBS 0.012934f
C217 B.n177 VSUBS 0.012934f
C218 B.n178 VSUBS 0.012934f
C219 B.n179 VSUBS 0.012934f
C220 B.n180 VSUBS 0.012934f
C221 B.n181 VSUBS 0.012934f
C222 B.n182 VSUBS 0.012934f
C223 B.n183 VSUBS 0.012934f
C224 B.n184 VSUBS 0.012934f
C225 B.n185 VSUBS 0.012934f
C226 B.n186 VSUBS 0.012934f
C227 B.n187 VSUBS 0.012934f
C228 B.n188 VSUBS 0.012934f
C229 B.n189 VSUBS 0.012934f
C230 B.n190 VSUBS 0.012934f
C231 B.n191 VSUBS 0.012934f
C232 B.n192 VSUBS 0.012934f
C233 B.n193 VSUBS 0.012934f
C234 B.n194 VSUBS 0.012934f
C235 B.n195 VSUBS 0.012934f
C236 B.n196 VSUBS 0.012934f
C237 B.n197 VSUBS 0.012934f
C238 B.n198 VSUBS 0.012934f
C239 B.n199 VSUBS 0.012934f
C240 B.n200 VSUBS 0.012934f
C241 B.n201 VSUBS 0.012934f
C242 B.n202 VSUBS 0.012934f
C243 B.n203 VSUBS 0.012934f
C244 B.n204 VSUBS 0.012934f
C245 B.n205 VSUBS 0.012934f
C246 B.n206 VSUBS 0.012934f
C247 B.n207 VSUBS 0.012934f
C248 B.n208 VSUBS 0.012934f
C249 B.n209 VSUBS 0.012934f
C250 B.n210 VSUBS 0.012934f
C251 B.n211 VSUBS 0.012934f
C252 B.n212 VSUBS 0.012934f
C253 B.n213 VSUBS 0.012934f
C254 B.n214 VSUBS 0.012934f
C255 B.n215 VSUBS 0.012934f
C256 B.n216 VSUBS 0.012934f
C257 B.n217 VSUBS 0.012934f
C258 B.n218 VSUBS 0.012934f
C259 B.n219 VSUBS 0.012934f
C260 B.n220 VSUBS 0.012934f
C261 B.n221 VSUBS 0.012934f
C262 B.n222 VSUBS 0.012934f
C263 B.n223 VSUBS 0.012934f
C264 B.n224 VSUBS 0.012934f
C265 B.n225 VSUBS 0.012934f
C266 B.n226 VSUBS 0.012934f
C267 B.n227 VSUBS 0.012934f
C268 B.n228 VSUBS 0.012934f
C269 B.n229 VSUBS 0.012934f
C270 B.n230 VSUBS 0.012934f
C271 B.n231 VSUBS 0.012934f
C272 B.n232 VSUBS 0.012934f
C273 B.n233 VSUBS 0.012934f
C274 B.n234 VSUBS 0.012934f
C275 B.n235 VSUBS 0.012934f
C276 B.n236 VSUBS 0.012934f
C277 B.n237 VSUBS 0.012934f
C278 B.n238 VSUBS 0.012934f
C279 B.n239 VSUBS 0.012934f
C280 B.n240 VSUBS 0.012934f
C281 B.n241 VSUBS 0.012934f
C282 B.n242 VSUBS 0.012934f
C283 B.n243 VSUBS 0.012934f
C284 B.n244 VSUBS 0.012934f
C285 B.n245 VSUBS 0.012934f
C286 B.n246 VSUBS 0.012934f
C287 B.n247 VSUBS 0.012934f
C288 B.n248 VSUBS 0.012934f
C289 B.n249 VSUBS 0.012934f
C290 B.n250 VSUBS 0.012934f
C291 B.n251 VSUBS 0.012934f
C292 B.n252 VSUBS 0.012934f
C293 B.n253 VSUBS 0.012934f
C294 B.n254 VSUBS 0.012934f
C295 B.n255 VSUBS 0.012934f
C296 B.n256 VSUBS 0.012934f
C297 B.n257 VSUBS 0.012934f
C298 B.n258 VSUBS 0.012934f
C299 B.n259 VSUBS 0.012934f
C300 B.n260 VSUBS 0.012934f
C301 B.n261 VSUBS 0.012934f
C302 B.n262 VSUBS 0.012934f
C303 B.n263 VSUBS 0.012934f
C304 B.n264 VSUBS 0.012934f
C305 B.n265 VSUBS 0.012934f
C306 B.n266 VSUBS 0.012934f
C307 B.n267 VSUBS 0.012934f
C308 B.n268 VSUBS 0.012934f
C309 B.n269 VSUBS 0.012934f
C310 B.n270 VSUBS 0.012934f
C311 B.n271 VSUBS 0.012934f
C312 B.n272 VSUBS 0.012934f
C313 B.n273 VSUBS 0.012934f
C314 B.n274 VSUBS 0.012934f
C315 B.n275 VSUBS 0.012934f
C316 B.n276 VSUBS 0.012934f
C317 B.n277 VSUBS 0.012934f
C318 B.n278 VSUBS 0.012934f
C319 B.n279 VSUBS 0.012934f
C320 B.n280 VSUBS 0.012934f
C321 B.n281 VSUBS 0.012934f
C322 B.n282 VSUBS 0.012934f
C323 B.n283 VSUBS 0.012934f
C324 B.n284 VSUBS 0.012934f
C325 B.n285 VSUBS 0.012934f
C326 B.n286 VSUBS 0.012934f
C327 B.n287 VSUBS 0.012934f
C328 B.n288 VSUBS 0.012934f
C329 B.n289 VSUBS 0.012934f
C330 B.n290 VSUBS 0.012934f
C331 B.n291 VSUBS 0.012934f
C332 B.n292 VSUBS 0.012934f
C333 B.n293 VSUBS 0.012934f
C334 B.n294 VSUBS 0.012934f
C335 B.n295 VSUBS 0.02733f
C336 B.n296 VSUBS 0.02733f
C337 B.n297 VSUBS 0.029352f
C338 B.n298 VSUBS 0.012934f
C339 B.n299 VSUBS 0.012934f
C340 B.n300 VSUBS 0.012934f
C341 B.n301 VSUBS 0.012934f
C342 B.n302 VSUBS 0.012934f
C343 B.n303 VSUBS 0.012934f
C344 B.n304 VSUBS 0.012934f
C345 B.n305 VSUBS 0.012934f
C346 B.n306 VSUBS 0.012934f
C347 B.n307 VSUBS 0.012934f
C348 B.n308 VSUBS 0.012934f
C349 B.n309 VSUBS 0.012934f
C350 B.n310 VSUBS 0.012934f
C351 B.n311 VSUBS 0.012934f
C352 B.n312 VSUBS 0.012934f
C353 B.n313 VSUBS 0.012934f
C354 B.n314 VSUBS 0.012934f
C355 B.n315 VSUBS 0.012934f
C356 B.n316 VSUBS 0.012934f
C357 B.n317 VSUBS 0.012934f
C358 B.n318 VSUBS 0.012934f
C359 B.n319 VSUBS 0.012934f
C360 B.n320 VSUBS 0.012934f
C361 B.n321 VSUBS 0.012934f
C362 B.n322 VSUBS 0.012934f
C363 B.n323 VSUBS 0.012934f
C364 B.n324 VSUBS 0.012934f
C365 B.n325 VSUBS 0.00894f
C366 B.n326 VSUBS 0.012934f
C367 B.n327 VSUBS 0.012934f
C368 B.n328 VSUBS 0.010462f
C369 B.n329 VSUBS 0.012934f
C370 B.n330 VSUBS 0.012934f
C371 B.n331 VSUBS 0.012934f
C372 B.n332 VSUBS 0.012934f
C373 B.n333 VSUBS 0.012934f
C374 B.n334 VSUBS 0.012934f
C375 B.n335 VSUBS 0.012934f
C376 B.n336 VSUBS 0.012934f
C377 B.n337 VSUBS 0.012934f
C378 B.n338 VSUBS 0.012934f
C379 B.n339 VSUBS 0.012934f
C380 B.n340 VSUBS 0.010462f
C381 B.n341 VSUBS 0.029967f
C382 B.n342 VSUBS 0.00894f
C383 B.n343 VSUBS 0.012934f
C384 B.n344 VSUBS 0.012934f
C385 B.n345 VSUBS 0.012934f
C386 B.n346 VSUBS 0.012934f
C387 B.n347 VSUBS 0.012934f
C388 B.n348 VSUBS 0.012934f
C389 B.n349 VSUBS 0.012934f
C390 B.n350 VSUBS 0.012934f
C391 B.n351 VSUBS 0.012934f
C392 B.n352 VSUBS 0.012934f
C393 B.n353 VSUBS 0.012934f
C394 B.n354 VSUBS 0.012934f
C395 B.n355 VSUBS 0.012934f
C396 B.n356 VSUBS 0.012934f
C397 B.n357 VSUBS 0.012934f
C398 B.n358 VSUBS 0.012934f
C399 B.n359 VSUBS 0.012934f
C400 B.n360 VSUBS 0.012934f
C401 B.n361 VSUBS 0.012934f
C402 B.n362 VSUBS 0.012934f
C403 B.n363 VSUBS 0.012934f
C404 B.n364 VSUBS 0.012934f
C405 B.n365 VSUBS 0.012934f
C406 B.n366 VSUBS 0.012934f
C407 B.n367 VSUBS 0.012934f
C408 B.n368 VSUBS 0.012934f
C409 B.n369 VSUBS 0.012934f
C410 B.n370 VSUBS 0.029352f
C411 B.n371 VSUBS 0.029352f
C412 B.n372 VSUBS 0.02733f
C413 B.n373 VSUBS 0.012934f
C414 B.n374 VSUBS 0.012934f
C415 B.n375 VSUBS 0.012934f
C416 B.n376 VSUBS 0.012934f
C417 B.n377 VSUBS 0.012934f
C418 B.n378 VSUBS 0.012934f
C419 B.n379 VSUBS 0.012934f
C420 B.n380 VSUBS 0.012934f
C421 B.n381 VSUBS 0.012934f
C422 B.n382 VSUBS 0.012934f
C423 B.n383 VSUBS 0.012934f
C424 B.n384 VSUBS 0.012934f
C425 B.n385 VSUBS 0.012934f
C426 B.n386 VSUBS 0.012934f
C427 B.n387 VSUBS 0.012934f
C428 B.n388 VSUBS 0.012934f
C429 B.n389 VSUBS 0.012934f
C430 B.n390 VSUBS 0.012934f
C431 B.n391 VSUBS 0.012934f
C432 B.n392 VSUBS 0.012934f
C433 B.n393 VSUBS 0.012934f
C434 B.n394 VSUBS 0.012934f
C435 B.n395 VSUBS 0.012934f
C436 B.n396 VSUBS 0.012934f
C437 B.n397 VSUBS 0.012934f
C438 B.n398 VSUBS 0.012934f
C439 B.n399 VSUBS 0.012934f
C440 B.n400 VSUBS 0.012934f
C441 B.n401 VSUBS 0.012934f
C442 B.n402 VSUBS 0.012934f
C443 B.n403 VSUBS 0.012934f
C444 B.n404 VSUBS 0.012934f
C445 B.n405 VSUBS 0.012934f
C446 B.n406 VSUBS 0.012934f
C447 B.n407 VSUBS 0.012934f
C448 B.n408 VSUBS 0.012934f
C449 B.n409 VSUBS 0.012934f
C450 B.n410 VSUBS 0.012934f
C451 B.n411 VSUBS 0.012934f
C452 B.n412 VSUBS 0.012934f
C453 B.n413 VSUBS 0.012934f
C454 B.n414 VSUBS 0.012934f
C455 B.n415 VSUBS 0.012934f
C456 B.n416 VSUBS 0.012934f
C457 B.n417 VSUBS 0.012934f
C458 B.n418 VSUBS 0.012934f
C459 B.n419 VSUBS 0.012934f
C460 B.n420 VSUBS 0.012934f
C461 B.n421 VSUBS 0.012934f
C462 B.n422 VSUBS 0.012934f
C463 B.n423 VSUBS 0.012934f
C464 B.n424 VSUBS 0.012934f
C465 B.n425 VSUBS 0.012934f
C466 B.n426 VSUBS 0.012934f
C467 B.n427 VSUBS 0.012934f
C468 B.n428 VSUBS 0.012934f
C469 B.n429 VSUBS 0.012934f
C470 B.n430 VSUBS 0.012934f
C471 B.n431 VSUBS 0.012934f
C472 B.n432 VSUBS 0.012934f
C473 B.n433 VSUBS 0.012934f
C474 B.n434 VSUBS 0.012934f
C475 B.n435 VSUBS 0.012934f
C476 B.n436 VSUBS 0.012934f
C477 B.n437 VSUBS 0.012934f
C478 B.n438 VSUBS 0.012934f
C479 B.n439 VSUBS 0.012934f
C480 B.n440 VSUBS 0.012934f
C481 B.n441 VSUBS 0.012934f
C482 B.n442 VSUBS 0.012934f
C483 B.n443 VSUBS 0.012934f
C484 B.n444 VSUBS 0.012934f
C485 B.n445 VSUBS 0.012934f
C486 B.n446 VSUBS 0.012934f
C487 B.n447 VSUBS 0.012934f
C488 B.n448 VSUBS 0.012934f
C489 B.n449 VSUBS 0.012934f
C490 B.n450 VSUBS 0.012934f
C491 B.n451 VSUBS 0.012934f
C492 B.n452 VSUBS 0.012934f
C493 B.n453 VSUBS 0.012934f
C494 B.n454 VSUBS 0.012934f
C495 B.n455 VSUBS 0.012934f
C496 B.n456 VSUBS 0.012934f
C497 B.n457 VSUBS 0.012934f
C498 B.n458 VSUBS 0.012934f
C499 B.n459 VSUBS 0.012934f
C500 B.n460 VSUBS 0.012934f
C501 B.n461 VSUBS 0.012934f
C502 B.n462 VSUBS 0.012934f
C503 B.n463 VSUBS 0.012934f
C504 B.n464 VSUBS 0.012934f
C505 B.n465 VSUBS 0.012934f
C506 B.n466 VSUBS 0.012934f
C507 B.n467 VSUBS 0.012934f
C508 B.n468 VSUBS 0.012934f
C509 B.n469 VSUBS 0.012934f
C510 B.n470 VSUBS 0.012934f
C511 B.n471 VSUBS 0.012934f
C512 B.n472 VSUBS 0.012934f
C513 B.n473 VSUBS 0.012934f
C514 B.n474 VSUBS 0.012934f
C515 B.n475 VSUBS 0.012934f
C516 B.n476 VSUBS 0.012934f
C517 B.n477 VSUBS 0.012934f
C518 B.n478 VSUBS 0.012934f
C519 B.n479 VSUBS 0.012934f
C520 B.n480 VSUBS 0.012934f
C521 B.n481 VSUBS 0.012934f
C522 B.n482 VSUBS 0.012934f
C523 B.n483 VSUBS 0.012934f
C524 B.n484 VSUBS 0.012934f
C525 B.n485 VSUBS 0.012934f
C526 B.n486 VSUBS 0.012934f
C527 B.n487 VSUBS 0.012934f
C528 B.n488 VSUBS 0.012934f
C529 B.n489 VSUBS 0.012934f
C530 B.n490 VSUBS 0.012934f
C531 B.n491 VSUBS 0.012934f
C532 B.n492 VSUBS 0.012934f
C533 B.n493 VSUBS 0.012934f
C534 B.n494 VSUBS 0.012934f
C535 B.n495 VSUBS 0.012934f
C536 B.n496 VSUBS 0.012934f
C537 B.n497 VSUBS 0.012934f
C538 B.n498 VSUBS 0.012934f
C539 B.n499 VSUBS 0.012934f
C540 B.n500 VSUBS 0.012934f
C541 B.n501 VSUBS 0.012934f
C542 B.n502 VSUBS 0.012934f
C543 B.n503 VSUBS 0.012934f
C544 B.n504 VSUBS 0.012934f
C545 B.n505 VSUBS 0.012934f
C546 B.n506 VSUBS 0.012934f
C547 B.n507 VSUBS 0.012934f
C548 B.n508 VSUBS 0.012934f
C549 B.n509 VSUBS 0.012934f
C550 B.n510 VSUBS 0.012934f
C551 B.n511 VSUBS 0.012934f
C552 B.n512 VSUBS 0.012934f
C553 B.n513 VSUBS 0.012934f
C554 B.n514 VSUBS 0.012934f
C555 B.n515 VSUBS 0.012934f
C556 B.n516 VSUBS 0.012934f
C557 B.n517 VSUBS 0.012934f
C558 B.n518 VSUBS 0.012934f
C559 B.n519 VSUBS 0.012934f
C560 B.n520 VSUBS 0.012934f
C561 B.n521 VSUBS 0.012934f
C562 B.n522 VSUBS 0.012934f
C563 B.n523 VSUBS 0.012934f
C564 B.n524 VSUBS 0.012934f
C565 B.n525 VSUBS 0.012934f
C566 B.n526 VSUBS 0.012934f
C567 B.n527 VSUBS 0.012934f
C568 B.n528 VSUBS 0.012934f
C569 B.n529 VSUBS 0.012934f
C570 B.n530 VSUBS 0.012934f
C571 B.n531 VSUBS 0.012934f
C572 B.n532 VSUBS 0.012934f
C573 B.n533 VSUBS 0.012934f
C574 B.n534 VSUBS 0.012934f
C575 B.n535 VSUBS 0.012934f
C576 B.n536 VSUBS 0.012934f
C577 B.n537 VSUBS 0.012934f
C578 B.n538 VSUBS 0.012934f
C579 B.n539 VSUBS 0.012934f
C580 B.n540 VSUBS 0.012934f
C581 B.n541 VSUBS 0.012934f
C582 B.n542 VSUBS 0.012934f
C583 B.n543 VSUBS 0.012934f
C584 B.n544 VSUBS 0.012934f
C585 B.n545 VSUBS 0.012934f
C586 B.n546 VSUBS 0.012934f
C587 B.n547 VSUBS 0.012934f
C588 B.n548 VSUBS 0.012934f
C589 B.n549 VSUBS 0.012934f
C590 B.n550 VSUBS 0.012934f
C591 B.n551 VSUBS 0.012934f
C592 B.n552 VSUBS 0.012934f
C593 B.n553 VSUBS 0.012934f
C594 B.n554 VSUBS 0.012934f
C595 B.n555 VSUBS 0.012934f
C596 B.n556 VSUBS 0.012934f
C597 B.n557 VSUBS 0.012934f
C598 B.n558 VSUBS 0.012934f
C599 B.n559 VSUBS 0.012934f
C600 B.n560 VSUBS 0.012934f
C601 B.n561 VSUBS 0.012934f
C602 B.n562 VSUBS 0.012934f
C603 B.n563 VSUBS 0.012934f
C604 B.n564 VSUBS 0.012934f
C605 B.n565 VSUBS 0.012934f
C606 B.n566 VSUBS 0.012934f
C607 B.n567 VSUBS 0.012934f
C608 B.n568 VSUBS 0.012934f
C609 B.n569 VSUBS 0.012934f
C610 B.n570 VSUBS 0.012934f
C611 B.n571 VSUBS 0.012934f
C612 B.n572 VSUBS 0.012934f
C613 B.n573 VSUBS 0.012934f
C614 B.n574 VSUBS 0.012934f
C615 B.n575 VSUBS 0.012934f
C616 B.n576 VSUBS 0.029022f
C617 B.n577 VSUBS 0.02766f
C618 B.n578 VSUBS 0.029352f
C619 B.n579 VSUBS 0.012934f
C620 B.n580 VSUBS 0.012934f
C621 B.n581 VSUBS 0.012934f
C622 B.n582 VSUBS 0.012934f
C623 B.n583 VSUBS 0.012934f
C624 B.n584 VSUBS 0.012934f
C625 B.n585 VSUBS 0.012934f
C626 B.n586 VSUBS 0.012934f
C627 B.n587 VSUBS 0.012934f
C628 B.n588 VSUBS 0.012934f
C629 B.n589 VSUBS 0.012934f
C630 B.n590 VSUBS 0.012934f
C631 B.n591 VSUBS 0.012934f
C632 B.n592 VSUBS 0.012934f
C633 B.n593 VSUBS 0.012934f
C634 B.n594 VSUBS 0.012934f
C635 B.n595 VSUBS 0.012934f
C636 B.n596 VSUBS 0.012934f
C637 B.n597 VSUBS 0.012934f
C638 B.n598 VSUBS 0.012934f
C639 B.n599 VSUBS 0.012934f
C640 B.n600 VSUBS 0.012934f
C641 B.n601 VSUBS 0.012934f
C642 B.n602 VSUBS 0.012934f
C643 B.n603 VSUBS 0.012934f
C644 B.n604 VSUBS 0.012934f
C645 B.n605 VSUBS 0.012934f
C646 B.n606 VSUBS 0.00894f
C647 B.n607 VSUBS 0.029967f
C648 B.n608 VSUBS 0.010462f
C649 B.n609 VSUBS 0.012934f
C650 B.n610 VSUBS 0.012934f
C651 B.n611 VSUBS 0.012934f
C652 B.n612 VSUBS 0.012934f
C653 B.n613 VSUBS 0.012934f
C654 B.n614 VSUBS 0.012934f
C655 B.n615 VSUBS 0.012934f
C656 B.n616 VSUBS 0.012934f
C657 B.n617 VSUBS 0.012934f
C658 B.n618 VSUBS 0.012934f
C659 B.n619 VSUBS 0.012934f
C660 B.n620 VSUBS 0.010462f
C661 B.n621 VSUBS 0.012934f
C662 B.n622 VSUBS 0.012934f
C663 B.n623 VSUBS 0.00894f
C664 B.n624 VSUBS 0.012934f
C665 B.n625 VSUBS 0.012934f
C666 B.n626 VSUBS 0.012934f
C667 B.n627 VSUBS 0.012934f
C668 B.n628 VSUBS 0.012934f
C669 B.n629 VSUBS 0.012934f
C670 B.n630 VSUBS 0.012934f
C671 B.n631 VSUBS 0.012934f
C672 B.n632 VSUBS 0.012934f
C673 B.n633 VSUBS 0.012934f
C674 B.n634 VSUBS 0.012934f
C675 B.n635 VSUBS 0.012934f
C676 B.n636 VSUBS 0.012934f
C677 B.n637 VSUBS 0.012934f
C678 B.n638 VSUBS 0.012934f
C679 B.n639 VSUBS 0.012934f
C680 B.n640 VSUBS 0.012934f
C681 B.n641 VSUBS 0.012934f
C682 B.n642 VSUBS 0.012934f
C683 B.n643 VSUBS 0.012934f
C684 B.n644 VSUBS 0.012934f
C685 B.n645 VSUBS 0.012934f
C686 B.n646 VSUBS 0.012934f
C687 B.n647 VSUBS 0.012934f
C688 B.n648 VSUBS 0.012934f
C689 B.n649 VSUBS 0.012934f
C690 B.n650 VSUBS 0.012934f
C691 B.n651 VSUBS 0.029352f
C692 B.n652 VSUBS 0.02733f
C693 B.n653 VSUBS 0.02733f
C694 B.n654 VSUBS 0.012934f
C695 B.n655 VSUBS 0.012934f
C696 B.n656 VSUBS 0.012934f
C697 B.n657 VSUBS 0.012934f
C698 B.n658 VSUBS 0.012934f
C699 B.n659 VSUBS 0.012934f
C700 B.n660 VSUBS 0.012934f
C701 B.n661 VSUBS 0.012934f
C702 B.n662 VSUBS 0.012934f
C703 B.n663 VSUBS 0.012934f
C704 B.n664 VSUBS 0.012934f
C705 B.n665 VSUBS 0.012934f
C706 B.n666 VSUBS 0.012934f
C707 B.n667 VSUBS 0.012934f
C708 B.n668 VSUBS 0.012934f
C709 B.n669 VSUBS 0.012934f
C710 B.n670 VSUBS 0.012934f
C711 B.n671 VSUBS 0.012934f
C712 B.n672 VSUBS 0.012934f
C713 B.n673 VSUBS 0.012934f
C714 B.n674 VSUBS 0.012934f
C715 B.n675 VSUBS 0.012934f
C716 B.n676 VSUBS 0.012934f
C717 B.n677 VSUBS 0.012934f
C718 B.n678 VSUBS 0.012934f
C719 B.n679 VSUBS 0.012934f
C720 B.n680 VSUBS 0.012934f
C721 B.n681 VSUBS 0.012934f
C722 B.n682 VSUBS 0.012934f
C723 B.n683 VSUBS 0.012934f
C724 B.n684 VSUBS 0.012934f
C725 B.n685 VSUBS 0.012934f
C726 B.n686 VSUBS 0.012934f
C727 B.n687 VSUBS 0.012934f
C728 B.n688 VSUBS 0.012934f
C729 B.n689 VSUBS 0.012934f
C730 B.n690 VSUBS 0.012934f
C731 B.n691 VSUBS 0.012934f
C732 B.n692 VSUBS 0.012934f
C733 B.n693 VSUBS 0.012934f
C734 B.n694 VSUBS 0.012934f
C735 B.n695 VSUBS 0.012934f
C736 B.n696 VSUBS 0.012934f
C737 B.n697 VSUBS 0.012934f
C738 B.n698 VSUBS 0.012934f
C739 B.n699 VSUBS 0.012934f
C740 B.n700 VSUBS 0.012934f
C741 B.n701 VSUBS 0.012934f
C742 B.n702 VSUBS 0.012934f
C743 B.n703 VSUBS 0.012934f
C744 B.n704 VSUBS 0.012934f
C745 B.n705 VSUBS 0.012934f
C746 B.n706 VSUBS 0.012934f
C747 B.n707 VSUBS 0.012934f
C748 B.n708 VSUBS 0.012934f
C749 B.n709 VSUBS 0.012934f
C750 B.n710 VSUBS 0.012934f
C751 B.n711 VSUBS 0.012934f
C752 B.n712 VSUBS 0.012934f
C753 B.n713 VSUBS 0.012934f
C754 B.n714 VSUBS 0.012934f
C755 B.n715 VSUBS 0.012934f
C756 B.n716 VSUBS 0.012934f
C757 B.n717 VSUBS 0.012934f
C758 B.n718 VSUBS 0.012934f
C759 B.n719 VSUBS 0.012934f
C760 B.n720 VSUBS 0.012934f
C761 B.n721 VSUBS 0.012934f
C762 B.n722 VSUBS 0.012934f
C763 B.n723 VSUBS 0.012934f
C764 B.n724 VSUBS 0.012934f
C765 B.n725 VSUBS 0.012934f
C766 B.n726 VSUBS 0.012934f
C767 B.n727 VSUBS 0.012934f
C768 B.n728 VSUBS 0.012934f
C769 B.n729 VSUBS 0.012934f
C770 B.n730 VSUBS 0.012934f
C771 B.n731 VSUBS 0.012934f
C772 B.n732 VSUBS 0.012934f
C773 B.n733 VSUBS 0.012934f
C774 B.n734 VSUBS 0.012934f
C775 B.n735 VSUBS 0.012934f
C776 B.n736 VSUBS 0.012934f
C777 B.n737 VSUBS 0.012934f
C778 B.n738 VSUBS 0.012934f
C779 B.n739 VSUBS 0.012934f
C780 B.n740 VSUBS 0.012934f
C781 B.n741 VSUBS 0.012934f
C782 B.n742 VSUBS 0.012934f
C783 B.n743 VSUBS 0.012934f
C784 B.n744 VSUBS 0.012934f
C785 B.n745 VSUBS 0.012934f
C786 B.n746 VSUBS 0.012934f
C787 B.n747 VSUBS 0.012934f
C788 B.n748 VSUBS 0.012934f
C789 B.n749 VSUBS 0.012934f
C790 B.n750 VSUBS 0.012934f
C791 B.n751 VSUBS 0.012934f
C792 B.n752 VSUBS 0.012934f
C793 B.n753 VSUBS 0.012934f
C794 B.n754 VSUBS 0.012934f
C795 B.n755 VSUBS 0.029288f
C796 VDD2.n0 VSUBS 0.037541f
C797 VDD2.n1 VSUBS 0.036562f
C798 VDD2.n2 VSUBS 0.019646f
C799 VDD2.n3 VSUBS 0.046437f
C800 VDD2.n4 VSUBS 0.020802f
C801 VDD2.n5 VSUBS 0.585139f
C802 VDD2.n6 VSUBS 0.019646f
C803 VDD2.t1 VSUBS 0.100377f
C804 VDD2.n7 VSUBS 0.145767f
C805 VDD2.n8 VSUBS 0.029419f
C806 VDD2.n9 VSUBS 0.034828f
C807 VDD2.n10 VSUBS 0.046437f
C808 VDD2.n11 VSUBS 0.020802f
C809 VDD2.n12 VSUBS 0.019646f
C810 VDD2.n13 VSUBS 0.036562f
C811 VDD2.n14 VSUBS 0.036562f
C812 VDD2.n15 VSUBS 0.019646f
C813 VDD2.n16 VSUBS 0.020802f
C814 VDD2.n17 VSUBS 0.046437f
C815 VDD2.n18 VSUBS 0.103452f
C816 VDD2.n19 VSUBS 0.020802f
C817 VDD2.n20 VSUBS 0.019646f
C818 VDD2.n21 VSUBS 0.080514f
C819 VDD2.n22 VSUBS 0.100772f
C820 VDD2.t8 VSUBS 0.129436f
C821 VDD2.t2 VSUBS 0.129436f
C822 VDD2.n23 VSUBS 0.78422f
C823 VDD2.n24 VSUBS 1.35392f
C824 VDD2.t0 VSUBS 0.129436f
C825 VDD2.t7 VSUBS 0.129436f
C826 VDD2.n25 VSUBS 0.807725f
C827 VDD2.n26 VSUBS 4.17568f
C828 VDD2.n27 VSUBS 0.037541f
C829 VDD2.n28 VSUBS 0.036562f
C830 VDD2.n29 VSUBS 0.019646f
C831 VDD2.n30 VSUBS 0.046437f
C832 VDD2.n31 VSUBS 0.020802f
C833 VDD2.n32 VSUBS 0.585139f
C834 VDD2.n33 VSUBS 0.019646f
C835 VDD2.t6 VSUBS 0.100377f
C836 VDD2.n34 VSUBS 0.145767f
C837 VDD2.n35 VSUBS 0.029419f
C838 VDD2.n36 VSUBS 0.034828f
C839 VDD2.n37 VSUBS 0.046437f
C840 VDD2.n38 VSUBS 0.020802f
C841 VDD2.n39 VSUBS 0.019646f
C842 VDD2.n40 VSUBS 0.036562f
C843 VDD2.n41 VSUBS 0.036562f
C844 VDD2.n42 VSUBS 0.019646f
C845 VDD2.n43 VSUBS 0.020802f
C846 VDD2.n44 VSUBS 0.046437f
C847 VDD2.n45 VSUBS 0.103452f
C848 VDD2.n46 VSUBS 0.020802f
C849 VDD2.n47 VSUBS 0.019646f
C850 VDD2.n48 VSUBS 0.080514f
C851 VDD2.n49 VSUBS 0.07678f
C852 VDD2.n50 VSUBS 3.62931f
C853 VDD2.t9 VSUBS 0.129436f
C854 VDD2.t4 VSUBS 0.129436f
C855 VDD2.n51 VSUBS 0.784224f
C856 VDD2.n52 VSUBS 0.977627f
C857 VDD2.t3 VSUBS 0.129436f
C858 VDD2.t5 VSUBS 0.129436f
C859 VDD2.n53 VSUBS 0.80768f
C860 VN.t2 VSUBS 1.32319f
C861 VN.n0 VSUBS 0.644293f
C862 VN.n1 VSUBS 0.03721f
C863 VN.n2 VSUBS 0.033628f
C864 VN.n3 VSUBS 0.03721f
C865 VN.t9 VSUBS 1.32319f
C866 VN.n4 VSUBS 0.510582f
C867 VN.n5 VSUBS 0.03721f
C868 VN.n6 VSUBS 0.048428f
C869 VN.n7 VSUBS 0.03721f
C870 VN.t7 VSUBS 1.32319f
C871 VN.n8 VSUBS 0.069003f
C872 VN.n9 VSUBS 0.03721f
C873 VN.n10 VSUBS 0.069003f
C874 VN.t8 VSUBS 1.69168f
C875 VN.n11 VSUBS 0.606429f
C876 VN.t1 VSUBS 1.32319f
C877 VN.n12 VSUBS 0.639475f
C878 VN.n13 VSUBS 0.061508f
C879 VN.n14 VSUBS 0.426571f
C880 VN.n15 VSUBS 0.03721f
C881 VN.n16 VSUBS 0.03721f
C882 VN.n17 VSUBS 0.059753f
C883 VN.n18 VSUBS 0.048428f
C884 VN.n19 VSUBS 0.069003f
C885 VN.n20 VSUBS 0.03721f
C886 VN.n21 VSUBS 0.03721f
C887 VN.n22 VSUBS 0.03721f
C888 VN.n23 VSUBS 0.54552f
C889 VN.n24 VSUBS 0.069003f
C890 VN.n25 VSUBS 0.069003f
C891 VN.n26 VSUBS 0.03721f
C892 VN.n27 VSUBS 0.03721f
C893 VN.n28 VSUBS 0.03721f
C894 VN.n29 VSUBS 0.059753f
C895 VN.n30 VSUBS 0.069003f
C896 VN.n31 VSUBS 0.061508f
C897 VN.n32 VSUBS 0.03721f
C898 VN.n33 VSUBS 0.03721f
C899 VN.n34 VSUBS 0.042432f
C900 VN.n35 VSUBS 0.069003f
C901 VN.n36 VSUBS 0.074553f
C902 VN.n37 VSUBS 0.03721f
C903 VN.n38 VSUBS 0.03721f
C904 VN.n39 VSUBS 0.03721f
C905 VN.n40 VSUBS 0.069003f
C906 VN.n41 VSUBS 0.069003f
C907 VN.n42 VSUBS 0.054014f
C908 VN.n43 VSUBS 0.060047f
C909 VN.n44 VSUBS 0.087605f
C910 VN.t3 VSUBS 1.32319f
C911 VN.n45 VSUBS 0.644293f
C912 VN.n46 VSUBS 0.03721f
C913 VN.n47 VSUBS 0.033628f
C914 VN.n48 VSUBS 0.03721f
C915 VN.t0 VSUBS 1.32319f
C916 VN.n49 VSUBS 0.510582f
C917 VN.n50 VSUBS 0.03721f
C918 VN.n51 VSUBS 0.048428f
C919 VN.n52 VSUBS 0.03721f
C920 VN.t5 VSUBS 1.32319f
C921 VN.n53 VSUBS 0.069003f
C922 VN.n54 VSUBS 0.03721f
C923 VN.n55 VSUBS 0.069003f
C924 VN.t4 VSUBS 1.69168f
C925 VN.n56 VSUBS 0.606429f
C926 VN.t6 VSUBS 1.32319f
C927 VN.n57 VSUBS 0.639475f
C928 VN.n58 VSUBS 0.061508f
C929 VN.n59 VSUBS 0.426571f
C930 VN.n60 VSUBS 0.03721f
C931 VN.n61 VSUBS 0.03721f
C932 VN.n62 VSUBS 0.059753f
C933 VN.n63 VSUBS 0.048428f
C934 VN.n64 VSUBS 0.069003f
C935 VN.n65 VSUBS 0.03721f
C936 VN.n66 VSUBS 0.03721f
C937 VN.n67 VSUBS 0.03721f
C938 VN.n68 VSUBS 0.54552f
C939 VN.n69 VSUBS 0.069003f
C940 VN.n70 VSUBS 0.069003f
C941 VN.n71 VSUBS 0.03721f
C942 VN.n72 VSUBS 0.03721f
C943 VN.n73 VSUBS 0.03721f
C944 VN.n74 VSUBS 0.059753f
C945 VN.n75 VSUBS 0.069003f
C946 VN.n76 VSUBS 0.061508f
C947 VN.n77 VSUBS 0.03721f
C948 VN.n78 VSUBS 0.03721f
C949 VN.n79 VSUBS 0.042432f
C950 VN.n80 VSUBS 0.069003f
C951 VN.n81 VSUBS 0.074553f
C952 VN.n82 VSUBS 0.03721f
C953 VN.n83 VSUBS 0.03721f
C954 VN.n84 VSUBS 0.03721f
C955 VN.n85 VSUBS 0.069003f
C956 VN.n86 VSUBS 0.069003f
C957 VN.n87 VSUBS 0.054014f
C958 VN.n88 VSUBS 0.060047f
C959 VN.n89 VSUBS 2.12351f
C960 VDD1.n0 VSUBS 0.037472f
C961 VDD1.n1 VSUBS 0.036495f
C962 VDD1.n2 VSUBS 0.019611f
C963 VDD1.n3 VSUBS 0.046353f
C964 VDD1.n4 VSUBS 0.020764f
C965 VDD1.n5 VSUBS 0.584073f
C966 VDD1.n6 VSUBS 0.019611f
C967 VDD1.t2 VSUBS 0.100194f
C968 VDD1.n7 VSUBS 0.145501f
C969 VDD1.n8 VSUBS 0.029365f
C970 VDD1.n9 VSUBS 0.034764f
C971 VDD1.n10 VSUBS 0.046353f
C972 VDD1.n11 VSUBS 0.020764f
C973 VDD1.n12 VSUBS 0.019611f
C974 VDD1.n13 VSUBS 0.036495f
C975 VDD1.n14 VSUBS 0.036495f
C976 VDD1.n15 VSUBS 0.019611f
C977 VDD1.n16 VSUBS 0.020764f
C978 VDD1.n17 VSUBS 0.046353f
C979 VDD1.n18 VSUBS 0.103264f
C980 VDD1.n19 VSUBS 0.020764f
C981 VDD1.n20 VSUBS 0.019611f
C982 VDD1.n21 VSUBS 0.080368f
C983 VDD1.n22 VSUBS 0.100588f
C984 VDD1.t3 VSUBS 0.1292f
C985 VDD1.t5 VSUBS 0.1292f
C986 VDD1.n23 VSUBS 0.782795f
C987 VDD1.n24 VSUBS 1.36355f
C988 VDD1.n25 VSUBS 0.037472f
C989 VDD1.n26 VSUBS 0.036495f
C990 VDD1.n27 VSUBS 0.019611f
C991 VDD1.n28 VSUBS 0.046353f
C992 VDD1.n29 VSUBS 0.020764f
C993 VDD1.n30 VSUBS 0.584073f
C994 VDD1.n31 VSUBS 0.019611f
C995 VDD1.t7 VSUBS 0.100194f
C996 VDD1.n32 VSUBS 0.145501f
C997 VDD1.n33 VSUBS 0.029365f
C998 VDD1.n34 VSUBS 0.034764f
C999 VDD1.n35 VSUBS 0.046353f
C1000 VDD1.n36 VSUBS 0.020764f
C1001 VDD1.n37 VSUBS 0.019611f
C1002 VDD1.n38 VSUBS 0.036495f
C1003 VDD1.n39 VSUBS 0.036495f
C1004 VDD1.n40 VSUBS 0.019611f
C1005 VDD1.n41 VSUBS 0.020764f
C1006 VDD1.n42 VSUBS 0.046353f
C1007 VDD1.n43 VSUBS 0.103264f
C1008 VDD1.n44 VSUBS 0.020764f
C1009 VDD1.n45 VSUBS 0.019611f
C1010 VDD1.n46 VSUBS 0.080368f
C1011 VDD1.n47 VSUBS 0.100588f
C1012 VDD1.t1 VSUBS 0.1292f
C1013 VDD1.t4 VSUBS 0.1292f
C1014 VDD1.n48 VSUBS 0.782791f
C1015 VDD1.n49 VSUBS 1.35146f
C1016 VDD1.t6 VSUBS 0.1292f
C1017 VDD1.t0 VSUBS 0.1292f
C1018 VDD1.n50 VSUBS 0.806254f
C1019 VDD1.n51 VSUBS 4.35895f
C1020 VDD1.t8 VSUBS 0.1292f
C1021 VDD1.t9 VSUBS 0.1292f
C1022 VDD1.n52 VSUBS 0.782791f
C1023 VDD1.n53 VSUBS 4.30366f
C1024 VTAIL.t3 VSUBS 0.128298f
C1025 VTAIL.t19 VSUBS 0.128298f
C1026 VTAIL.n0 VSUBS 0.674597f
C1027 VTAIL.n1 VSUBS 1.07737f
C1028 VTAIL.n2 VSUBS 0.037211f
C1029 VTAIL.n3 VSUBS 0.03624f
C1030 VTAIL.n4 VSUBS 0.019474f
C1031 VTAIL.n5 VSUBS 0.046029f
C1032 VTAIL.n6 VSUBS 0.020619f
C1033 VTAIL.n7 VSUBS 0.579995f
C1034 VTAIL.n8 VSUBS 0.019474f
C1035 VTAIL.t10 VSUBS 0.099495f
C1036 VTAIL.n9 VSUBS 0.144485f
C1037 VTAIL.n10 VSUBS 0.02916f
C1038 VTAIL.n11 VSUBS 0.034522f
C1039 VTAIL.n12 VSUBS 0.046029f
C1040 VTAIL.n13 VSUBS 0.020619f
C1041 VTAIL.n14 VSUBS 0.019474f
C1042 VTAIL.n15 VSUBS 0.03624f
C1043 VTAIL.n16 VSUBS 0.03624f
C1044 VTAIL.n17 VSUBS 0.019474f
C1045 VTAIL.n18 VSUBS 0.020619f
C1046 VTAIL.n19 VSUBS 0.046029f
C1047 VTAIL.n20 VSUBS 0.102543f
C1048 VTAIL.n21 VSUBS 0.020619f
C1049 VTAIL.n22 VSUBS 0.019474f
C1050 VTAIL.n23 VSUBS 0.079807f
C1051 VTAIL.n24 VSUBS 0.051049f
C1052 VTAIL.n25 VSUBS 0.595474f
C1053 VTAIL.t16 VSUBS 0.128298f
C1054 VTAIL.t13 VSUBS 0.128298f
C1055 VTAIL.n26 VSUBS 0.674597f
C1056 VTAIL.n27 VSUBS 1.27166f
C1057 VTAIL.t9 VSUBS 0.128298f
C1058 VTAIL.t17 VSUBS 0.128298f
C1059 VTAIL.n28 VSUBS 0.674597f
C1060 VTAIL.n29 VSUBS 2.55619f
C1061 VTAIL.t5 VSUBS 0.128298f
C1062 VTAIL.t7 VSUBS 0.128298f
C1063 VTAIL.n30 VSUBS 0.674602f
C1064 VTAIL.n31 VSUBS 2.55618f
C1065 VTAIL.t2 VSUBS 0.128298f
C1066 VTAIL.t0 VSUBS 0.128298f
C1067 VTAIL.n32 VSUBS 0.674602f
C1068 VTAIL.n33 VSUBS 1.27166f
C1069 VTAIL.n34 VSUBS 0.037211f
C1070 VTAIL.n35 VSUBS 0.03624f
C1071 VTAIL.n36 VSUBS 0.019474f
C1072 VTAIL.n37 VSUBS 0.046029f
C1073 VTAIL.n38 VSUBS 0.020619f
C1074 VTAIL.n39 VSUBS 0.579995f
C1075 VTAIL.n40 VSUBS 0.019474f
C1076 VTAIL.t18 VSUBS 0.099495f
C1077 VTAIL.n41 VSUBS 0.144485f
C1078 VTAIL.n42 VSUBS 0.02916f
C1079 VTAIL.n43 VSUBS 0.034522f
C1080 VTAIL.n44 VSUBS 0.046029f
C1081 VTAIL.n45 VSUBS 0.020619f
C1082 VTAIL.n46 VSUBS 0.019474f
C1083 VTAIL.n47 VSUBS 0.03624f
C1084 VTAIL.n48 VSUBS 0.03624f
C1085 VTAIL.n49 VSUBS 0.019474f
C1086 VTAIL.n50 VSUBS 0.020619f
C1087 VTAIL.n51 VSUBS 0.046029f
C1088 VTAIL.n52 VSUBS 0.102543f
C1089 VTAIL.n53 VSUBS 0.020619f
C1090 VTAIL.n54 VSUBS 0.019474f
C1091 VTAIL.n55 VSUBS 0.079807f
C1092 VTAIL.n56 VSUBS 0.051049f
C1093 VTAIL.n57 VSUBS 0.595474f
C1094 VTAIL.t14 VSUBS 0.128298f
C1095 VTAIL.t8 VSUBS 0.128298f
C1096 VTAIL.n58 VSUBS 0.674602f
C1097 VTAIL.n59 VSUBS 1.15589f
C1098 VTAIL.t11 VSUBS 0.128298f
C1099 VTAIL.t15 VSUBS 0.128298f
C1100 VTAIL.n60 VSUBS 0.674602f
C1101 VTAIL.n61 VSUBS 1.27166f
C1102 VTAIL.n62 VSUBS 0.037211f
C1103 VTAIL.n63 VSUBS 0.03624f
C1104 VTAIL.n64 VSUBS 0.019474f
C1105 VTAIL.n65 VSUBS 0.046029f
C1106 VTAIL.n66 VSUBS 0.020619f
C1107 VTAIL.n67 VSUBS 0.579995f
C1108 VTAIL.n68 VSUBS 0.019474f
C1109 VTAIL.t12 VSUBS 0.099495f
C1110 VTAIL.n69 VSUBS 0.144485f
C1111 VTAIL.n70 VSUBS 0.02916f
C1112 VTAIL.n71 VSUBS 0.034522f
C1113 VTAIL.n72 VSUBS 0.046029f
C1114 VTAIL.n73 VSUBS 0.020619f
C1115 VTAIL.n74 VSUBS 0.019474f
C1116 VTAIL.n75 VSUBS 0.03624f
C1117 VTAIL.n76 VSUBS 0.03624f
C1118 VTAIL.n77 VSUBS 0.019474f
C1119 VTAIL.n78 VSUBS 0.020619f
C1120 VTAIL.n79 VSUBS 0.046029f
C1121 VTAIL.n80 VSUBS 0.102543f
C1122 VTAIL.n81 VSUBS 0.020619f
C1123 VTAIL.n82 VSUBS 0.019474f
C1124 VTAIL.n83 VSUBS 0.079807f
C1125 VTAIL.n84 VSUBS 0.051049f
C1126 VTAIL.n85 VSUBS 1.65451f
C1127 VTAIL.n86 VSUBS 0.037211f
C1128 VTAIL.n87 VSUBS 0.03624f
C1129 VTAIL.n88 VSUBS 0.019474f
C1130 VTAIL.n89 VSUBS 0.046029f
C1131 VTAIL.n90 VSUBS 0.020619f
C1132 VTAIL.n91 VSUBS 0.579995f
C1133 VTAIL.n92 VSUBS 0.019474f
C1134 VTAIL.t4 VSUBS 0.099495f
C1135 VTAIL.n93 VSUBS 0.144485f
C1136 VTAIL.n94 VSUBS 0.02916f
C1137 VTAIL.n95 VSUBS 0.034522f
C1138 VTAIL.n96 VSUBS 0.046029f
C1139 VTAIL.n97 VSUBS 0.020619f
C1140 VTAIL.n98 VSUBS 0.019474f
C1141 VTAIL.n99 VSUBS 0.03624f
C1142 VTAIL.n100 VSUBS 0.03624f
C1143 VTAIL.n101 VSUBS 0.019474f
C1144 VTAIL.n102 VSUBS 0.020619f
C1145 VTAIL.n103 VSUBS 0.046029f
C1146 VTAIL.n104 VSUBS 0.102543f
C1147 VTAIL.n105 VSUBS 0.020619f
C1148 VTAIL.n106 VSUBS 0.019474f
C1149 VTAIL.n107 VSUBS 0.079807f
C1150 VTAIL.n108 VSUBS 0.051049f
C1151 VTAIL.n109 VSUBS 1.65451f
C1152 VTAIL.t6 VSUBS 0.128298f
C1153 VTAIL.t1 VSUBS 0.128298f
C1154 VTAIL.n110 VSUBS 0.674597f
C1155 VTAIL.n111 VSUBS 1.00892f
C1156 VP.t9 VSUBS 1.4959f
C1157 VP.n0 VSUBS 0.728389f
C1158 VP.n1 VSUBS 0.042067f
C1159 VP.n2 VSUBS 0.038017f
C1160 VP.n3 VSUBS 0.042067f
C1161 VP.t3 VSUBS 1.4959f
C1162 VP.n4 VSUBS 0.577226f
C1163 VP.n5 VSUBS 0.042067f
C1164 VP.n6 VSUBS 0.054749f
C1165 VP.n7 VSUBS 0.042067f
C1166 VP.t5 VSUBS 1.4959f
C1167 VP.n8 VSUBS 0.078009f
C1168 VP.n9 VSUBS 0.042067f
C1169 VP.n10 VSUBS 0.078009f
C1170 VP.n11 VSUBS 0.042067f
C1171 VP.t8 VSUBS 1.4959f
C1172 VP.n12 VSUBS 0.084284f
C1173 VP.n13 VSUBS 0.042067f
C1174 VP.n14 VSUBS 0.061064f
C1175 VP.t0 VSUBS 1.4959f
C1176 VP.n15 VSUBS 0.728389f
C1177 VP.n16 VSUBS 0.042067f
C1178 VP.n17 VSUBS 0.038017f
C1179 VP.n18 VSUBS 0.042067f
C1180 VP.t1 VSUBS 1.4959f
C1181 VP.n19 VSUBS 0.577226f
C1182 VP.n20 VSUBS 0.042067f
C1183 VP.n21 VSUBS 0.054749f
C1184 VP.n22 VSUBS 0.042067f
C1185 VP.t4 VSUBS 1.4959f
C1186 VP.n23 VSUBS 0.078009f
C1187 VP.n24 VSUBS 0.042067f
C1188 VP.n25 VSUBS 0.078009f
C1189 VP.t7 VSUBS 1.91248f
C1190 VP.n26 VSUBS 0.685585f
C1191 VP.t6 VSUBS 1.4959f
C1192 VP.n27 VSUBS 0.722943f
C1193 VP.n28 VSUBS 0.069537f
C1194 VP.n29 VSUBS 0.482251f
C1195 VP.n30 VSUBS 0.042067f
C1196 VP.n31 VSUBS 0.042067f
C1197 VP.n32 VSUBS 0.067552f
C1198 VP.n33 VSUBS 0.054749f
C1199 VP.n34 VSUBS 0.078009f
C1200 VP.n35 VSUBS 0.042067f
C1201 VP.n36 VSUBS 0.042067f
C1202 VP.n37 VSUBS 0.042067f
C1203 VP.n38 VSUBS 0.616724f
C1204 VP.n39 VSUBS 0.078009f
C1205 VP.n40 VSUBS 0.078009f
C1206 VP.n41 VSUBS 0.042067f
C1207 VP.n42 VSUBS 0.042067f
C1208 VP.n43 VSUBS 0.042067f
C1209 VP.n44 VSUBS 0.067552f
C1210 VP.n45 VSUBS 0.078009f
C1211 VP.n46 VSUBS 0.069537f
C1212 VP.n47 VSUBS 0.042067f
C1213 VP.n48 VSUBS 0.042067f
C1214 VP.n49 VSUBS 0.04797f
C1215 VP.n50 VSUBS 0.078009f
C1216 VP.n51 VSUBS 0.084284f
C1217 VP.n52 VSUBS 0.042067f
C1218 VP.n53 VSUBS 0.042067f
C1219 VP.n54 VSUBS 0.042067f
C1220 VP.n55 VSUBS 0.078009f
C1221 VP.n56 VSUBS 0.078009f
C1222 VP.n57 VSUBS 0.061064f
C1223 VP.n58 VSUBS 0.067884f
C1224 VP.n59 VSUBS 2.38345f
C1225 VP.t2 VSUBS 1.4959f
C1226 VP.n60 VSUBS 0.728389f
C1227 VP.n61 VSUBS 2.41381f
C1228 VP.n62 VSUBS 0.067884f
C1229 VP.n63 VSUBS 0.042067f
C1230 VP.n64 VSUBS 0.078009f
C1231 VP.n65 VSUBS 0.078009f
C1232 VP.n66 VSUBS 0.038017f
C1233 VP.n67 VSUBS 0.042067f
C1234 VP.n68 VSUBS 0.042067f
C1235 VP.n69 VSUBS 0.042067f
C1236 VP.n70 VSUBS 0.078009f
C1237 VP.n71 VSUBS 0.04797f
C1238 VP.n72 VSUBS 0.577226f
C1239 VP.n73 VSUBS 0.069537f
C1240 VP.n74 VSUBS 0.042067f
C1241 VP.n75 VSUBS 0.042067f
C1242 VP.n76 VSUBS 0.042067f
C1243 VP.n77 VSUBS 0.067552f
C1244 VP.n78 VSUBS 0.054749f
C1245 VP.n79 VSUBS 0.078009f
C1246 VP.n80 VSUBS 0.042067f
C1247 VP.n81 VSUBS 0.042067f
C1248 VP.n82 VSUBS 0.042067f
C1249 VP.n83 VSUBS 0.616724f
C1250 VP.n84 VSUBS 0.078009f
C1251 VP.n85 VSUBS 0.078009f
C1252 VP.n86 VSUBS 0.042067f
C1253 VP.n87 VSUBS 0.042067f
C1254 VP.n88 VSUBS 0.042067f
C1255 VP.n89 VSUBS 0.067552f
C1256 VP.n90 VSUBS 0.078009f
C1257 VP.n91 VSUBS 0.069537f
C1258 VP.n92 VSUBS 0.042067f
C1259 VP.n93 VSUBS 0.042067f
C1260 VP.n94 VSUBS 0.04797f
C1261 VP.n95 VSUBS 0.078009f
C1262 VP.n96 VSUBS 0.084284f
C1263 VP.n97 VSUBS 0.042067f
C1264 VP.n98 VSUBS 0.042067f
C1265 VP.n99 VSUBS 0.042067f
C1266 VP.n100 VSUBS 0.078009f
C1267 VP.n101 VSUBS 0.078009f
C1268 VP.n102 VSUBS 0.061064f
C1269 VP.n103 VSUBS 0.067884f
C1270 VP.n104 VSUBS 0.09904f
.ends

