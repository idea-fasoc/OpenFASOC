* NGSPICE file created from diff_pair_sample_1730.ext - technology: sky130A

.subckt diff_pair_sample_1730 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=0 ps=0 w=18.73 l=2.55
X1 B.t8 B.t6 B.t7 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=0 ps=0 w=18.73 l=2.55
X2 VDD2.t1 VN.t0 VTAIL.t2 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=7.3047 ps=38.24 w=18.73 l=2.55
X3 VDD2.t0 VN.t1 VTAIL.t3 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=7.3047 ps=38.24 w=18.73 l=2.55
X4 B.t5 B.t3 B.t4 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=0 ps=0 w=18.73 l=2.55
X5 VDD1.t1 VP.t0 VTAIL.t1 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=7.3047 ps=38.24 w=18.73 l=2.55
X6 VDD1.t0 VP.t1 VTAIL.t0 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=7.3047 ps=38.24 w=18.73 l=2.55
X7 B.t2 B.t0 B.t1 w_n2122_n4714# sky130_fd_pr__pfet_01v8 ad=7.3047 pd=38.24 as=0 ps=0 w=18.73 l=2.55
R0 B.n506 B.n505 585
R1 B.n507 B.n84 585
R2 B.n509 B.n508 585
R3 B.n510 B.n83 585
R4 B.n512 B.n511 585
R5 B.n513 B.n82 585
R6 B.n515 B.n514 585
R7 B.n516 B.n81 585
R8 B.n518 B.n517 585
R9 B.n519 B.n80 585
R10 B.n521 B.n520 585
R11 B.n522 B.n79 585
R12 B.n524 B.n523 585
R13 B.n525 B.n78 585
R14 B.n527 B.n526 585
R15 B.n528 B.n77 585
R16 B.n530 B.n529 585
R17 B.n531 B.n76 585
R18 B.n533 B.n532 585
R19 B.n534 B.n75 585
R20 B.n536 B.n535 585
R21 B.n537 B.n74 585
R22 B.n539 B.n538 585
R23 B.n540 B.n73 585
R24 B.n542 B.n541 585
R25 B.n543 B.n72 585
R26 B.n545 B.n544 585
R27 B.n546 B.n71 585
R28 B.n548 B.n547 585
R29 B.n549 B.n70 585
R30 B.n551 B.n550 585
R31 B.n552 B.n69 585
R32 B.n554 B.n553 585
R33 B.n555 B.n68 585
R34 B.n557 B.n556 585
R35 B.n558 B.n67 585
R36 B.n560 B.n559 585
R37 B.n561 B.n66 585
R38 B.n563 B.n562 585
R39 B.n564 B.n65 585
R40 B.n566 B.n565 585
R41 B.n567 B.n64 585
R42 B.n569 B.n568 585
R43 B.n570 B.n63 585
R44 B.n572 B.n571 585
R45 B.n573 B.n62 585
R46 B.n575 B.n574 585
R47 B.n576 B.n61 585
R48 B.n578 B.n577 585
R49 B.n579 B.n60 585
R50 B.n581 B.n580 585
R51 B.n582 B.n59 585
R52 B.n584 B.n583 585
R53 B.n585 B.n58 585
R54 B.n587 B.n586 585
R55 B.n588 B.n57 585
R56 B.n590 B.n589 585
R57 B.n591 B.n56 585
R58 B.n593 B.n592 585
R59 B.n594 B.n55 585
R60 B.n596 B.n595 585
R61 B.n598 B.n597 585
R62 B.n599 B.n51 585
R63 B.n601 B.n600 585
R64 B.n602 B.n50 585
R65 B.n604 B.n603 585
R66 B.n605 B.n49 585
R67 B.n607 B.n606 585
R68 B.n608 B.n48 585
R69 B.n610 B.n609 585
R70 B.n611 B.n45 585
R71 B.n614 B.n613 585
R72 B.n615 B.n44 585
R73 B.n617 B.n616 585
R74 B.n618 B.n43 585
R75 B.n620 B.n619 585
R76 B.n621 B.n42 585
R77 B.n623 B.n622 585
R78 B.n624 B.n41 585
R79 B.n626 B.n625 585
R80 B.n627 B.n40 585
R81 B.n629 B.n628 585
R82 B.n630 B.n39 585
R83 B.n632 B.n631 585
R84 B.n633 B.n38 585
R85 B.n635 B.n634 585
R86 B.n636 B.n37 585
R87 B.n638 B.n637 585
R88 B.n639 B.n36 585
R89 B.n641 B.n640 585
R90 B.n642 B.n35 585
R91 B.n644 B.n643 585
R92 B.n645 B.n34 585
R93 B.n647 B.n646 585
R94 B.n648 B.n33 585
R95 B.n650 B.n649 585
R96 B.n651 B.n32 585
R97 B.n653 B.n652 585
R98 B.n654 B.n31 585
R99 B.n656 B.n655 585
R100 B.n657 B.n30 585
R101 B.n659 B.n658 585
R102 B.n660 B.n29 585
R103 B.n662 B.n661 585
R104 B.n663 B.n28 585
R105 B.n665 B.n664 585
R106 B.n666 B.n27 585
R107 B.n668 B.n667 585
R108 B.n669 B.n26 585
R109 B.n671 B.n670 585
R110 B.n672 B.n25 585
R111 B.n674 B.n673 585
R112 B.n675 B.n24 585
R113 B.n677 B.n676 585
R114 B.n678 B.n23 585
R115 B.n680 B.n679 585
R116 B.n681 B.n22 585
R117 B.n683 B.n682 585
R118 B.n684 B.n21 585
R119 B.n686 B.n685 585
R120 B.n687 B.n20 585
R121 B.n689 B.n688 585
R122 B.n690 B.n19 585
R123 B.n692 B.n691 585
R124 B.n693 B.n18 585
R125 B.n695 B.n694 585
R126 B.n696 B.n17 585
R127 B.n698 B.n697 585
R128 B.n699 B.n16 585
R129 B.n701 B.n700 585
R130 B.n702 B.n15 585
R131 B.n704 B.n703 585
R132 B.n504 B.n85 585
R133 B.n503 B.n502 585
R134 B.n501 B.n86 585
R135 B.n500 B.n499 585
R136 B.n498 B.n87 585
R137 B.n497 B.n496 585
R138 B.n495 B.n88 585
R139 B.n494 B.n493 585
R140 B.n492 B.n89 585
R141 B.n491 B.n490 585
R142 B.n489 B.n90 585
R143 B.n488 B.n487 585
R144 B.n486 B.n91 585
R145 B.n485 B.n484 585
R146 B.n483 B.n92 585
R147 B.n482 B.n481 585
R148 B.n480 B.n93 585
R149 B.n479 B.n478 585
R150 B.n477 B.n94 585
R151 B.n476 B.n475 585
R152 B.n474 B.n95 585
R153 B.n473 B.n472 585
R154 B.n471 B.n96 585
R155 B.n470 B.n469 585
R156 B.n468 B.n97 585
R157 B.n467 B.n466 585
R158 B.n465 B.n98 585
R159 B.n464 B.n463 585
R160 B.n462 B.n99 585
R161 B.n461 B.n460 585
R162 B.n459 B.n100 585
R163 B.n458 B.n457 585
R164 B.n456 B.n101 585
R165 B.n455 B.n454 585
R166 B.n453 B.n102 585
R167 B.n452 B.n451 585
R168 B.n450 B.n103 585
R169 B.n449 B.n448 585
R170 B.n447 B.n104 585
R171 B.n446 B.n445 585
R172 B.n444 B.n105 585
R173 B.n443 B.n442 585
R174 B.n441 B.n106 585
R175 B.n440 B.n439 585
R176 B.n438 B.n107 585
R177 B.n437 B.n436 585
R178 B.n435 B.n108 585
R179 B.n434 B.n433 585
R180 B.n432 B.n109 585
R181 B.n431 B.n430 585
R182 B.n429 B.n110 585
R183 B.n230 B.n229 585
R184 B.n231 B.n180 585
R185 B.n233 B.n232 585
R186 B.n234 B.n179 585
R187 B.n236 B.n235 585
R188 B.n237 B.n178 585
R189 B.n239 B.n238 585
R190 B.n240 B.n177 585
R191 B.n242 B.n241 585
R192 B.n243 B.n176 585
R193 B.n245 B.n244 585
R194 B.n246 B.n175 585
R195 B.n248 B.n247 585
R196 B.n249 B.n174 585
R197 B.n251 B.n250 585
R198 B.n252 B.n173 585
R199 B.n254 B.n253 585
R200 B.n255 B.n172 585
R201 B.n257 B.n256 585
R202 B.n258 B.n171 585
R203 B.n260 B.n259 585
R204 B.n261 B.n170 585
R205 B.n263 B.n262 585
R206 B.n264 B.n169 585
R207 B.n266 B.n265 585
R208 B.n267 B.n168 585
R209 B.n269 B.n268 585
R210 B.n270 B.n167 585
R211 B.n272 B.n271 585
R212 B.n273 B.n166 585
R213 B.n275 B.n274 585
R214 B.n276 B.n165 585
R215 B.n278 B.n277 585
R216 B.n279 B.n164 585
R217 B.n281 B.n280 585
R218 B.n282 B.n163 585
R219 B.n284 B.n283 585
R220 B.n285 B.n162 585
R221 B.n287 B.n286 585
R222 B.n288 B.n161 585
R223 B.n290 B.n289 585
R224 B.n291 B.n160 585
R225 B.n293 B.n292 585
R226 B.n294 B.n159 585
R227 B.n296 B.n295 585
R228 B.n297 B.n158 585
R229 B.n299 B.n298 585
R230 B.n300 B.n157 585
R231 B.n302 B.n301 585
R232 B.n303 B.n156 585
R233 B.n305 B.n304 585
R234 B.n306 B.n155 585
R235 B.n308 B.n307 585
R236 B.n309 B.n154 585
R237 B.n311 B.n310 585
R238 B.n312 B.n153 585
R239 B.n314 B.n313 585
R240 B.n315 B.n152 585
R241 B.n317 B.n316 585
R242 B.n318 B.n151 585
R243 B.n320 B.n319 585
R244 B.n322 B.n321 585
R245 B.n323 B.n147 585
R246 B.n325 B.n324 585
R247 B.n326 B.n146 585
R248 B.n328 B.n327 585
R249 B.n329 B.n145 585
R250 B.n331 B.n330 585
R251 B.n332 B.n144 585
R252 B.n334 B.n333 585
R253 B.n335 B.n141 585
R254 B.n338 B.n337 585
R255 B.n339 B.n140 585
R256 B.n341 B.n340 585
R257 B.n342 B.n139 585
R258 B.n344 B.n343 585
R259 B.n345 B.n138 585
R260 B.n347 B.n346 585
R261 B.n348 B.n137 585
R262 B.n350 B.n349 585
R263 B.n351 B.n136 585
R264 B.n353 B.n352 585
R265 B.n354 B.n135 585
R266 B.n356 B.n355 585
R267 B.n357 B.n134 585
R268 B.n359 B.n358 585
R269 B.n360 B.n133 585
R270 B.n362 B.n361 585
R271 B.n363 B.n132 585
R272 B.n365 B.n364 585
R273 B.n366 B.n131 585
R274 B.n368 B.n367 585
R275 B.n369 B.n130 585
R276 B.n371 B.n370 585
R277 B.n372 B.n129 585
R278 B.n374 B.n373 585
R279 B.n375 B.n128 585
R280 B.n377 B.n376 585
R281 B.n378 B.n127 585
R282 B.n380 B.n379 585
R283 B.n381 B.n126 585
R284 B.n383 B.n382 585
R285 B.n384 B.n125 585
R286 B.n386 B.n385 585
R287 B.n387 B.n124 585
R288 B.n389 B.n388 585
R289 B.n390 B.n123 585
R290 B.n392 B.n391 585
R291 B.n393 B.n122 585
R292 B.n395 B.n394 585
R293 B.n396 B.n121 585
R294 B.n398 B.n397 585
R295 B.n399 B.n120 585
R296 B.n401 B.n400 585
R297 B.n402 B.n119 585
R298 B.n404 B.n403 585
R299 B.n405 B.n118 585
R300 B.n407 B.n406 585
R301 B.n408 B.n117 585
R302 B.n410 B.n409 585
R303 B.n411 B.n116 585
R304 B.n413 B.n412 585
R305 B.n414 B.n115 585
R306 B.n416 B.n415 585
R307 B.n417 B.n114 585
R308 B.n419 B.n418 585
R309 B.n420 B.n113 585
R310 B.n422 B.n421 585
R311 B.n423 B.n112 585
R312 B.n425 B.n424 585
R313 B.n426 B.n111 585
R314 B.n428 B.n427 585
R315 B.n228 B.n181 585
R316 B.n227 B.n226 585
R317 B.n225 B.n182 585
R318 B.n224 B.n223 585
R319 B.n222 B.n183 585
R320 B.n221 B.n220 585
R321 B.n219 B.n184 585
R322 B.n218 B.n217 585
R323 B.n216 B.n185 585
R324 B.n215 B.n214 585
R325 B.n213 B.n186 585
R326 B.n212 B.n211 585
R327 B.n210 B.n187 585
R328 B.n209 B.n208 585
R329 B.n207 B.n188 585
R330 B.n206 B.n205 585
R331 B.n204 B.n189 585
R332 B.n203 B.n202 585
R333 B.n201 B.n190 585
R334 B.n200 B.n199 585
R335 B.n198 B.n191 585
R336 B.n197 B.n196 585
R337 B.n195 B.n192 585
R338 B.n194 B.n193 585
R339 B.n2 B.n0 585
R340 B.n741 B.n1 585
R341 B.n740 B.n739 585
R342 B.n738 B.n3 585
R343 B.n737 B.n736 585
R344 B.n735 B.n4 585
R345 B.n734 B.n733 585
R346 B.n732 B.n5 585
R347 B.n731 B.n730 585
R348 B.n729 B.n6 585
R349 B.n728 B.n727 585
R350 B.n726 B.n7 585
R351 B.n725 B.n724 585
R352 B.n723 B.n8 585
R353 B.n722 B.n721 585
R354 B.n720 B.n9 585
R355 B.n719 B.n718 585
R356 B.n717 B.n10 585
R357 B.n716 B.n715 585
R358 B.n714 B.n11 585
R359 B.n713 B.n712 585
R360 B.n711 B.n12 585
R361 B.n710 B.n709 585
R362 B.n708 B.n13 585
R363 B.n707 B.n706 585
R364 B.n705 B.n14 585
R365 B.n743 B.n742 585
R366 B.n142 B.t2 552.506
R367 B.n52 B.t4 552.506
R368 B.n148 B.t11 552.506
R369 B.n46 B.t7 552.506
R370 B.n230 B.n181 540.549
R371 B.n705 B.n704 540.549
R372 B.n429 B.n428 540.549
R373 B.n506 B.n85 540.549
R374 B.n143 B.t1 496.652
R375 B.n53 B.t5 496.652
R376 B.n149 B.t10 496.652
R377 B.n47 B.t8 496.652
R378 B.n142 B.t0 384.988
R379 B.n148 B.t9 384.988
R380 B.n46 B.t6 384.988
R381 B.n52 B.t3 384.988
R382 B.n226 B.n181 163.367
R383 B.n226 B.n225 163.367
R384 B.n225 B.n224 163.367
R385 B.n224 B.n183 163.367
R386 B.n220 B.n183 163.367
R387 B.n220 B.n219 163.367
R388 B.n219 B.n218 163.367
R389 B.n218 B.n185 163.367
R390 B.n214 B.n185 163.367
R391 B.n214 B.n213 163.367
R392 B.n213 B.n212 163.367
R393 B.n212 B.n187 163.367
R394 B.n208 B.n187 163.367
R395 B.n208 B.n207 163.367
R396 B.n207 B.n206 163.367
R397 B.n206 B.n189 163.367
R398 B.n202 B.n189 163.367
R399 B.n202 B.n201 163.367
R400 B.n201 B.n200 163.367
R401 B.n200 B.n191 163.367
R402 B.n196 B.n191 163.367
R403 B.n196 B.n195 163.367
R404 B.n195 B.n194 163.367
R405 B.n194 B.n2 163.367
R406 B.n742 B.n2 163.367
R407 B.n742 B.n741 163.367
R408 B.n741 B.n740 163.367
R409 B.n740 B.n3 163.367
R410 B.n736 B.n3 163.367
R411 B.n736 B.n735 163.367
R412 B.n735 B.n734 163.367
R413 B.n734 B.n5 163.367
R414 B.n730 B.n5 163.367
R415 B.n730 B.n729 163.367
R416 B.n729 B.n728 163.367
R417 B.n728 B.n7 163.367
R418 B.n724 B.n7 163.367
R419 B.n724 B.n723 163.367
R420 B.n723 B.n722 163.367
R421 B.n722 B.n9 163.367
R422 B.n718 B.n9 163.367
R423 B.n718 B.n717 163.367
R424 B.n717 B.n716 163.367
R425 B.n716 B.n11 163.367
R426 B.n712 B.n11 163.367
R427 B.n712 B.n711 163.367
R428 B.n711 B.n710 163.367
R429 B.n710 B.n13 163.367
R430 B.n706 B.n13 163.367
R431 B.n706 B.n705 163.367
R432 B.n231 B.n230 163.367
R433 B.n232 B.n231 163.367
R434 B.n232 B.n179 163.367
R435 B.n236 B.n179 163.367
R436 B.n237 B.n236 163.367
R437 B.n238 B.n237 163.367
R438 B.n238 B.n177 163.367
R439 B.n242 B.n177 163.367
R440 B.n243 B.n242 163.367
R441 B.n244 B.n243 163.367
R442 B.n244 B.n175 163.367
R443 B.n248 B.n175 163.367
R444 B.n249 B.n248 163.367
R445 B.n250 B.n249 163.367
R446 B.n250 B.n173 163.367
R447 B.n254 B.n173 163.367
R448 B.n255 B.n254 163.367
R449 B.n256 B.n255 163.367
R450 B.n256 B.n171 163.367
R451 B.n260 B.n171 163.367
R452 B.n261 B.n260 163.367
R453 B.n262 B.n261 163.367
R454 B.n262 B.n169 163.367
R455 B.n266 B.n169 163.367
R456 B.n267 B.n266 163.367
R457 B.n268 B.n267 163.367
R458 B.n268 B.n167 163.367
R459 B.n272 B.n167 163.367
R460 B.n273 B.n272 163.367
R461 B.n274 B.n273 163.367
R462 B.n274 B.n165 163.367
R463 B.n278 B.n165 163.367
R464 B.n279 B.n278 163.367
R465 B.n280 B.n279 163.367
R466 B.n280 B.n163 163.367
R467 B.n284 B.n163 163.367
R468 B.n285 B.n284 163.367
R469 B.n286 B.n285 163.367
R470 B.n286 B.n161 163.367
R471 B.n290 B.n161 163.367
R472 B.n291 B.n290 163.367
R473 B.n292 B.n291 163.367
R474 B.n292 B.n159 163.367
R475 B.n296 B.n159 163.367
R476 B.n297 B.n296 163.367
R477 B.n298 B.n297 163.367
R478 B.n298 B.n157 163.367
R479 B.n302 B.n157 163.367
R480 B.n303 B.n302 163.367
R481 B.n304 B.n303 163.367
R482 B.n304 B.n155 163.367
R483 B.n308 B.n155 163.367
R484 B.n309 B.n308 163.367
R485 B.n310 B.n309 163.367
R486 B.n310 B.n153 163.367
R487 B.n314 B.n153 163.367
R488 B.n315 B.n314 163.367
R489 B.n316 B.n315 163.367
R490 B.n316 B.n151 163.367
R491 B.n320 B.n151 163.367
R492 B.n321 B.n320 163.367
R493 B.n321 B.n147 163.367
R494 B.n325 B.n147 163.367
R495 B.n326 B.n325 163.367
R496 B.n327 B.n326 163.367
R497 B.n327 B.n145 163.367
R498 B.n331 B.n145 163.367
R499 B.n332 B.n331 163.367
R500 B.n333 B.n332 163.367
R501 B.n333 B.n141 163.367
R502 B.n338 B.n141 163.367
R503 B.n339 B.n338 163.367
R504 B.n340 B.n339 163.367
R505 B.n340 B.n139 163.367
R506 B.n344 B.n139 163.367
R507 B.n345 B.n344 163.367
R508 B.n346 B.n345 163.367
R509 B.n346 B.n137 163.367
R510 B.n350 B.n137 163.367
R511 B.n351 B.n350 163.367
R512 B.n352 B.n351 163.367
R513 B.n352 B.n135 163.367
R514 B.n356 B.n135 163.367
R515 B.n357 B.n356 163.367
R516 B.n358 B.n357 163.367
R517 B.n358 B.n133 163.367
R518 B.n362 B.n133 163.367
R519 B.n363 B.n362 163.367
R520 B.n364 B.n363 163.367
R521 B.n364 B.n131 163.367
R522 B.n368 B.n131 163.367
R523 B.n369 B.n368 163.367
R524 B.n370 B.n369 163.367
R525 B.n370 B.n129 163.367
R526 B.n374 B.n129 163.367
R527 B.n375 B.n374 163.367
R528 B.n376 B.n375 163.367
R529 B.n376 B.n127 163.367
R530 B.n380 B.n127 163.367
R531 B.n381 B.n380 163.367
R532 B.n382 B.n381 163.367
R533 B.n382 B.n125 163.367
R534 B.n386 B.n125 163.367
R535 B.n387 B.n386 163.367
R536 B.n388 B.n387 163.367
R537 B.n388 B.n123 163.367
R538 B.n392 B.n123 163.367
R539 B.n393 B.n392 163.367
R540 B.n394 B.n393 163.367
R541 B.n394 B.n121 163.367
R542 B.n398 B.n121 163.367
R543 B.n399 B.n398 163.367
R544 B.n400 B.n399 163.367
R545 B.n400 B.n119 163.367
R546 B.n404 B.n119 163.367
R547 B.n405 B.n404 163.367
R548 B.n406 B.n405 163.367
R549 B.n406 B.n117 163.367
R550 B.n410 B.n117 163.367
R551 B.n411 B.n410 163.367
R552 B.n412 B.n411 163.367
R553 B.n412 B.n115 163.367
R554 B.n416 B.n115 163.367
R555 B.n417 B.n416 163.367
R556 B.n418 B.n417 163.367
R557 B.n418 B.n113 163.367
R558 B.n422 B.n113 163.367
R559 B.n423 B.n422 163.367
R560 B.n424 B.n423 163.367
R561 B.n424 B.n111 163.367
R562 B.n428 B.n111 163.367
R563 B.n430 B.n429 163.367
R564 B.n430 B.n109 163.367
R565 B.n434 B.n109 163.367
R566 B.n435 B.n434 163.367
R567 B.n436 B.n435 163.367
R568 B.n436 B.n107 163.367
R569 B.n440 B.n107 163.367
R570 B.n441 B.n440 163.367
R571 B.n442 B.n441 163.367
R572 B.n442 B.n105 163.367
R573 B.n446 B.n105 163.367
R574 B.n447 B.n446 163.367
R575 B.n448 B.n447 163.367
R576 B.n448 B.n103 163.367
R577 B.n452 B.n103 163.367
R578 B.n453 B.n452 163.367
R579 B.n454 B.n453 163.367
R580 B.n454 B.n101 163.367
R581 B.n458 B.n101 163.367
R582 B.n459 B.n458 163.367
R583 B.n460 B.n459 163.367
R584 B.n460 B.n99 163.367
R585 B.n464 B.n99 163.367
R586 B.n465 B.n464 163.367
R587 B.n466 B.n465 163.367
R588 B.n466 B.n97 163.367
R589 B.n470 B.n97 163.367
R590 B.n471 B.n470 163.367
R591 B.n472 B.n471 163.367
R592 B.n472 B.n95 163.367
R593 B.n476 B.n95 163.367
R594 B.n477 B.n476 163.367
R595 B.n478 B.n477 163.367
R596 B.n478 B.n93 163.367
R597 B.n482 B.n93 163.367
R598 B.n483 B.n482 163.367
R599 B.n484 B.n483 163.367
R600 B.n484 B.n91 163.367
R601 B.n488 B.n91 163.367
R602 B.n489 B.n488 163.367
R603 B.n490 B.n489 163.367
R604 B.n490 B.n89 163.367
R605 B.n494 B.n89 163.367
R606 B.n495 B.n494 163.367
R607 B.n496 B.n495 163.367
R608 B.n496 B.n87 163.367
R609 B.n500 B.n87 163.367
R610 B.n501 B.n500 163.367
R611 B.n502 B.n501 163.367
R612 B.n502 B.n85 163.367
R613 B.n704 B.n15 163.367
R614 B.n700 B.n15 163.367
R615 B.n700 B.n699 163.367
R616 B.n699 B.n698 163.367
R617 B.n698 B.n17 163.367
R618 B.n694 B.n17 163.367
R619 B.n694 B.n693 163.367
R620 B.n693 B.n692 163.367
R621 B.n692 B.n19 163.367
R622 B.n688 B.n19 163.367
R623 B.n688 B.n687 163.367
R624 B.n687 B.n686 163.367
R625 B.n686 B.n21 163.367
R626 B.n682 B.n21 163.367
R627 B.n682 B.n681 163.367
R628 B.n681 B.n680 163.367
R629 B.n680 B.n23 163.367
R630 B.n676 B.n23 163.367
R631 B.n676 B.n675 163.367
R632 B.n675 B.n674 163.367
R633 B.n674 B.n25 163.367
R634 B.n670 B.n25 163.367
R635 B.n670 B.n669 163.367
R636 B.n669 B.n668 163.367
R637 B.n668 B.n27 163.367
R638 B.n664 B.n27 163.367
R639 B.n664 B.n663 163.367
R640 B.n663 B.n662 163.367
R641 B.n662 B.n29 163.367
R642 B.n658 B.n29 163.367
R643 B.n658 B.n657 163.367
R644 B.n657 B.n656 163.367
R645 B.n656 B.n31 163.367
R646 B.n652 B.n31 163.367
R647 B.n652 B.n651 163.367
R648 B.n651 B.n650 163.367
R649 B.n650 B.n33 163.367
R650 B.n646 B.n33 163.367
R651 B.n646 B.n645 163.367
R652 B.n645 B.n644 163.367
R653 B.n644 B.n35 163.367
R654 B.n640 B.n35 163.367
R655 B.n640 B.n639 163.367
R656 B.n639 B.n638 163.367
R657 B.n638 B.n37 163.367
R658 B.n634 B.n37 163.367
R659 B.n634 B.n633 163.367
R660 B.n633 B.n632 163.367
R661 B.n632 B.n39 163.367
R662 B.n628 B.n39 163.367
R663 B.n628 B.n627 163.367
R664 B.n627 B.n626 163.367
R665 B.n626 B.n41 163.367
R666 B.n622 B.n41 163.367
R667 B.n622 B.n621 163.367
R668 B.n621 B.n620 163.367
R669 B.n620 B.n43 163.367
R670 B.n616 B.n43 163.367
R671 B.n616 B.n615 163.367
R672 B.n615 B.n614 163.367
R673 B.n614 B.n45 163.367
R674 B.n609 B.n45 163.367
R675 B.n609 B.n608 163.367
R676 B.n608 B.n607 163.367
R677 B.n607 B.n49 163.367
R678 B.n603 B.n49 163.367
R679 B.n603 B.n602 163.367
R680 B.n602 B.n601 163.367
R681 B.n601 B.n51 163.367
R682 B.n597 B.n51 163.367
R683 B.n597 B.n596 163.367
R684 B.n596 B.n55 163.367
R685 B.n592 B.n55 163.367
R686 B.n592 B.n591 163.367
R687 B.n591 B.n590 163.367
R688 B.n590 B.n57 163.367
R689 B.n586 B.n57 163.367
R690 B.n586 B.n585 163.367
R691 B.n585 B.n584 163.367
R692 B.n584 B.n59 163.367
R693 B.n580 B.n59 163.367
R694 B.n580 B.n579 163.367
R695 B.n579 B.n578 163.367
R696 B.n578 B.n61 163.367
R697 B.n574 B.n61 163.367
R698 B.n574 B.n573 163.367
R699 B.n573 B.n572 163.367
R700 B.n572 B.n63 163.367
R701 B.n568 B.n63 163.367
R702 B.n568 B.n567 163.367
R703 B.n567 B.n566 163.367
R704 B.n566 B.n65 163.367
R705 B.n562 B.n65 163.367
R706 B.n562 B.n561 163.367
R707 B.n561 B.n560 163.367
R708 B.n560 B.n67 163.367
R709 B.n556 B.n67 163.367
R710 B.n556 B.n555 163.367
R711 B.n555 B.n554 163.367
R712 B.n554 B.n69 163.367
R713 B.n550 B.n69 163.367
R714 B.n550 B.n549 163.367
R715 B.n549 B.n548 163.367
R716 B.n548 B.n71 163.367
R717 B.n544 B.n71 163.367
R718 B.n544 B.n543 163.367
R719 B.n543 B.n542 163.367
R720 B.n542 B.n73 163.367
R721 B.n538 B.n73 163.367
R722 B.n538 B.n537 163.367
R723 B.n537 B.n536 163.367
R724 B.n536 B.n75 163.367
R725 B.n532 B.n75 163.367
R726 B.n532 B.n531 163.367
R727 B.n531 B.n530 163.367
R728 B.n530 B.n77 163.367
R729 B.n526 B.n77 163.367
R730 B.n526 B.n525 163.367
R731 B.n525 B.n524 163.367
R732 B.n524 B.n79 163.367
R733 B.n520 B.n79 163.367
R734 B.n520 B.n519 163.367
R735 B.n519 B.n518 163.367
R736 B.n518 B.n81 163.367
R737 B.n514 B.n81 163.367
R738 B.n514 B.n513 163.367
R739 B.n513 B.n512 163.367
R740 B.n512 B.n83 163.367
R741 B.n508 B.n83 163.367
R742 B.n508 B.n507 163.367
R743 B.n507 B.n506 163.367
R744 B.n336 B.n143 59.5399
R745 B.n150 B.n149 59.5399
R746 B.n612 B.n47 59.5399
R747 B.n54 B.n53 59.5399
R748 B.n143 B.n142 55.855
R749 B.n149 B.n148 55.855
R750 B.n47 B.n46 55.855
R751 B.n53 B.n52 55.855
R752 B.n703 B.n14 35.1225
R753 B.n505 B.n504 35.1225
R754 B.n427 B.n110 35.1225
R755 B.n229 B.n228 35.1225
R756 B B.n743 18.0485
R757 B.n703 B.n702 10.6151
R758 B.n702 B.n701 10.6151
R759 B.n701 B.n16 10.6151
R760 B.n697 B.n16 10.6151
R761 B.n697 B.n696 10.6151
R762 B.n696 B.n695 10.6151
R763 B.n695 B.n18 10.6151
R764 B.n691 B.n18 10.6151
R765 B.n691 B.n690 10.6151
R766 B.n690 B.n689 10.6151
R767 B.n689 B.n20 10.6151
R768 B.n685 B.n20 10.6151
R769 B.n685 B.n684 10.6151
R770 B.n684 B.n683 10.6151
R771 B.n683 B.n22 10.6151
R772 B.n679 B.n22 10.6151
R773 B.n679 B.n678 10.6151
R774 B.n678 B.n677 10.6151
R775 B.n677 B.n24 10.6151
R776 B.n673 B.n24 10.6151
R777 B.n673 B.n672 10.6151
R778 B.n672 B.n671 10.6151
R779 B.n671 B.n26 10.6151
R780 B.n667 B.n26 10.6151
R781 B.n667 B.n666 10.6151
R782 B.n666 B.n665 10.6151
R783 B.n665 B.n28 10.6151
R784 B.n661 B.n28 10.6151
R785 B.n661 B.n660 10.6151
R786 B.n660 B.n659 10.6151
R787 B.n659 B.n30 10.6151
R788 B.n655 B.n30 10.6151
R789 B.n655 B.n654 10.6151
R790 B.n654 B.n653 10.6151
R791 B.n653 B.n32 10.6151
R792 B.n649 B.n32 10.6151
R793 B.n649 B.n648 10.6151
R794 B.n648 B.n647 10.6151
R795 B.n647 B.n34 10.6151
R796 B.n643 B.n34 10.6151
R797 B.n643 B.n642 10.6151
R798 B.n642 B.n641 10.6151
R799 B.n641 B.n36 10.6151
R800 B.n637 B.n36 10.6151
R801 B.n637 B.n636 10.6151
R802 B.n636 B.n635 10.6151
R803 B.n635 B.n38 10.6151
R804 B.n631 B.n38 10.6151
R805 B.n631 B.n630 10.6151
R806 B.n630 B.n629 10.6151
R807 B.n629 B.n40 10.6151
R808 B.n625 B.n40 10.6151
R809 B.n625 B.n624 10.6151
R810 B.n624 B.n623 10.6151
R811 B.n623 B.n42 10.6151
R812 B.n619 B.n42 10.6151
R813 B.n619 B.n618 10.6151
R814 B.n618 B.n617 10.6151
R815 B.n617 B.n44 10.6151
R816 B.n613 B.n44 10.6151
R817 B.n611 B.n610 10.6151
R818 B.n610 B.n48 10.6151
R819 B.n606 B.n48 10.6151
R820 B.n606 B.n605 10.6151
R821 B.n605 B.n604 10.6151
R822 B.n604 B.n50 10.6151
R823 B.n600 B.n50 10.6151
R824 B.n600 B.n599 10.6151
R825 B.n599 B.n598 10.6151
R826 B.n595 B.n594 10.6151
R827 B.n594 B.n593 10.6151
R828 B.n593 B.n56 10.6151
R829 B.n589 B.n56 10.6151
R830 B.n589 B.n588 10.6151
R831 B.n588 B.n587 10.6151
R832 B.n587 B.n58 10.6151
R833 B.n583 B.n58 10.6151
R834 B.n583 B.n582 10.6151
R835 B.n582 B.n581 10.6151
R836 B.n581 B.n60 10.6151
R837 B.n577 B.n60 10.6151
R838 B.n577 B.n576 10.6151
R839 B.n576 B.n575 10.6151
R840 B.n575 B.n62 10.6151
R841 B.n571 B.n62 10.6151
R842 B.n571 B.n570 10.6151
R843 B.n570 B.n569 10.6151
R844 B.n569 B.n64 10.6151
R845 B.n565 B.n64 10.6151
R846 B.n565 B.n564 10.6151
R847 B.n564 B.n563 10.6151
R848 B.n563 B.n66 10.6151
R849 B.n559 B.n66 10.6151
R850 B.n559 B.n558 10.6151
R851 B.n558 B.n557 10.6151
R852 B.n557 B.n68 10.6151
R853 B.n553 B.n68 10.6151
R854 B.n553 B.n552 10.6151
R855 B.n552 B.n551 10.6151
R856 B.n551 B.n70 10.6151
R857 B.n547 B.n70 10.6151
R858 B.n547 B.n546 10.6151
R859 B.n546 B.n545 10.6151
R860 B.n545 B.n72 10.6151
R861 B.n541 B.n72 10.6151
R862 B.n541 B.n540 10.6151
R863 B.n540 B.n539 10.6151
R864 B.n539 B.n74 10.6151
R865 B.n535 B.n74 10.6151
R866 B.n535 B.n534 10.6151
R867 B.n534 B.n533 10.6151
R868 B.n533 B.n76 10.6151
R869 B.n529 B.n76 10.6151
R870 B.n529 B.n528 10.6151
R871 B.n528 B.n527 10.6151
R872 B.n527 B.n78 10.6151
R873 B.n523 B.n78 10.6151
R874 B.n523 B.n522 10.6151
R875 B.n522 B.n521 10.6151
R876 B.n521 B.n80 10.6151
R877 B.n517 B.n80 10.6151
R878 B.n517 B.n516 10.6151
R879 B.n516 B.n515 10.6151
R880 B.n515 B.n82 10.6151
R881 B.n511 B.n82 10.6151
R882 B.n511 B.n510 10.6151
R883 B.n510 B.n509 10.6151
R884 B.n509 B.n84 10.6151
R885 B.n505 B.n84 10.6151
R886 B.n431 B.n110 10.6151
R887 B.n432 B.n431 10.6151
R888 B.n433 B.n432 10.6151
R889 B.n433 B.n108 10.6151
R890 B.n437 B.n108 10.6151
R891 B.n438 B.n437 10.6151
R892 B.n439 B.n438 10.6151
R893 B.n439 B.n106 10.6151
R894 B.n443 B.n106 10.6151
R895 B.n444 B.n443 10.6151
R896 B.n445 B.n444 10.6151
R897 B.n445 B.n104 10.6151
R898 B.n449 B.n104 10.6151
R899 B.n450 B.n449 10.6151
R900 B.n451 B.n450 10.6151
R901 B.n451 B.n102 10.6151
R902 B.n455 B.n102 10.6151
R903 B.n456 B.n455 10.6151
R904 B.n457 B.n456 10.6151
R905 B.n457 B.n100 10.6151
R906 B.n461 B.n100 10.6151
R907 B.n462 B.n461 10.6151
R908 B.n463 B.n462 10.6151
R909 B.n463 B.n98 10.6151
R910 B.n467 B.n98 10.6151
R911 B.n468 B.n467 10.6151
R912 B.n469 B.n468 10.6151
R913 B.n469 B.n96 10.6151
R914 B.n473 B.n96 10.6151
R915 B.n474 B.n473 10.6151
R916 B.n475 B.n474 10.6151
R917 B.n475 B.n94 10.6151
R918 B.n479 B.n94 10.6151
R919 B.n480 B.n479 10.6151
R920 B.n481 B.n480 10.6151
R921 B.n481 B.n92 10.6151
R922 B.n485 B.n92 10.6151
R923 B.n486 B.n485 10.6151
R924 B.n487 B.n486 10.6151
R925 B.n487 B.n90 10.6151
R926 B.n491 B.n90 10.6151
R927 B.n492 B.n491 10.6151
R928 B.n493 B.n492 10.6151
R929 B.n493 B.n88 10.6151
R930 B.n497 B.n88 10.6151
R931 B.n498 B.n497 10.6151
R932 B.n499 B.n498 10.6151
R933 B.n499 B.n86 10.6151
R934 B.n503 B.n86 10.6151
R935 B.n504 B.n503 10.6151
R936 B.n229 B.n180 10.6151
R937 B.n233 B.n180 10.6151
R938 B.n234 B.n233 10.6151
R939 B.n235 B.n234 10.6151
R940 B.n235 B.n178 10.6151
R941 B.n239 B.n178 10.6151
R942 B.n240 B.n239 10.6151
R943 B.n241 B.n240 10.6151
R944 B.n241 B.n176 10.6151
R945 B.n245 B.n176 10.6151
R946 B.n246 B.n245 10.6151
R947 B.n247 B.n246 10.6151
R948 B.n247 B.n174 10.6151
R949 B.n251 B.n174 10.6151
R950 B.n252 B.n251 10.6151
R951 B.n253 B.n252 10.6151
R952 B.n253 B.n172 10.6151
R953 B.n257 B.n172 10.6151
R954 B.n258 B.n257 10.6151
R955 B.n259 B.n258 10.6151
R956 B.n259 B.n170 10.6151
R957 B.n263 B.n170 10.6151
R958 B.n264 B.n263 10.6151
R959 B.n265 B.n264 10.6151
R960 B.n265 B.n168 10.6151
R961 B.n269 B.n168 10.6151
R962 B.n270 B.n269 10.6151
R963 B.n271 B.n270 10.6151
R964 B.n271 B.n166 10.6151
R965 B.n275 B.n166 10.6151
R966 B.n276 B.n275 10.6151
R967 B.n277 B.n276 10.6151
R968 B.n277 B.n164 10.6151
R969 B.n281 B.n164 10.6151
R970 B.n282 B.n281 10.6151
R971 B.n283 B.n282 10.6151
R972 B.n283 B.n162 10.6151
R973 B.n287 B.n162 10.6151
R974 B.n288 B.n287 10.6151
R975 B.n289 B.n288 10.6151
R976 B.n289 B.n160 10.6151
R977 B.n293 B.n160 10.6151
R978 B.n294 B.n293 10.6151
R979 B.n295 B.n294 10.6151
R980 B.n295 B.n158 10.6151
R981 B.n299 B.n158 10.6151
R982 B.n300 B.n299 10.6151
R983 B.n301 B.n300 10.6151
R984 B.n301 B.n156 10.6151
R985 B.n305 B.n156 10.6151
R986 B.n306 B.n305 10.6151
R987 B.n307 B.n306 10.6151
R988 B.n307 B.n154 10.6151
R989 B.n311 B.n154 10.6151
R990 B.n312 B.n311 10.6151
R991 B.n313 B.n312 10.6151
R992 B.n313 B.n152 10.6151
R993 B.n317 B.n152 10.6151
R994 B.n318 B.n317 10.6151
R995 B.n319 B.n318 10.6151
R996 B.n323 B.n322 10.6151
R997 B.n324 B.n323 10.6151
R998 B.n324 B.n146 10.6151
R999 B.n328 B.n146 10.6151
R1000 B.n329 B.n328 10.6151
R1001 B.n330 B.n329 10.6151
R1002 B.n330 B.n144 10.6151
R1003 B.n334 B.n144 10.6151
R1004 B.n335 B.n334 10.6151
R1005 B.n337 B.n140 10.6151
R1006 B.n341 B.n140 10.6151
R1007 B.n342 B.n341 10.6151
R1008 B.n343 B.n342 10.6151
R1009 B.n343 B.n138 10.6151
R1010 B.n347 B.n138 10.6151
R1011 B.n348 B.n347 10.6151
R1012 B.n349 B.n348 10.6151
R1013 B.n349 B.n136 10.6151
R1014 B.n353 B.n136 10.6151
R1015 B.n354 B.n353 10.6151
R1016 B.n355 B.n354 10.6151
R1017 B.n355 B.n134 10.6151
R1018 B.n359 B.n134 10.6151
R1019 B.n360 B.n359 10.6151
R1020 B.n361 B.n360 10.6151
R1021 B.n361 B.n132 10.6151
R1022 B.n365 B.n132 10.6151
R1023 B.n366 B.n365 10.6151
R1024 B.n367 B.n366 10.6151
R1025 B.n367 B.n130 10.6151
R1026 B.n371 B.n130 10.6151
R1027 B.n372 B.n371 10.6151
R1028 B.n373 B.n372 10.6151
R1029 B.n373 B.n128 10.6151
R1030 B.n377 B.n128 10.6151
R1031 B.n378 B.n377 10.6151
R1032 B.n379 B.n378 10.6151
R1033 B.n379 B.n126 10.6151
R1034 B.n383 B.n126 10.6151
R1035 B.n384 B.n383 10.6151
R1036 B.n385 B.n384 10.6151
R1037 B.n385 B.n124 10.6151
R1038 B.n389 B.n124 10.6151
R1039 B.n390 B.n389 10.6151
R1040 B.n391 B.n390 10.6151
R1041 B.n391 B.n122 10.6151
R1042 B.n395 B.n122 10.6151
R1043 B.n396 B.n395 10.6151
R1044 B.n397 B.n396 10.6151
R1045 B.n397 B.n120 10.6151
R1046 B.n401 B.n120 10.6151
R1047 B.n402 B.n401 10.6151
R1048 B.n403 B.n402 10.6151
R1049 B.n403 B.n118 10.6151
R1050 B.n407 B.n118 10.6151
R1051 B.n408 B.n407 10.6151
R1052 B.n409 B.n408 10.6151
R1053 B.n409 B.n116 10.6151
R1054 B.n413 B.n116 10.6151
R1055 B.n414 B.n413 10.6151
R1056 B.n415 B.n414 10.6151
R1057 B.n415 B.n114 10.6151
R1058 B.n419 B.n114 10.6151
R1059 B.n420 B.n419 10.6151
R1060 B.n421 B.n420 10.6151
R1061 B.n421 B.n112 10.6151
R1062 B.n425 B.n112 10.6151
R1063 B.n426 B.n425 10.6151
R1064 B.n427 B.n426 10.6151
R1065 B.n228 B.n227 10.6151
R1066 B.n227 B.n182 10.6151
R1067 B.n223 B.n182 10.6151
R1068 B.n223 B.n222 10.6151
R1069 B.n222 B.n221 10.6151
R1070 B.n221 B.n184 10.6151
R1071 B.n217 B.n184 10.6151
R1072 B.n217 B.n216 10.6151
R1073 B.n216 B.n215 10.6151
R1074 B.n215 B.n186 10.6151
R1075 B.n211 B.n186 10.6151
R1076 B.n211 B.n210 10.6151
R1077 B.n210 B.n209 10.6151
R1078 B.n209 B.n188 10.6151
R1079 B.n205 B.n188 10.6151
R1080 B.n205 B.n204 10.6151
R1081 B.n204 B.n203 10.6151
R1082 B.n203 B.n190 10.6151
R1083 B.n199 B.n190 10.6151
R1084 B.n199 B.n198 10.6151
R1085 B.n198 B.n197 10.6151
R1086 B.n197 B.n192 10.6151
R1087 B.n193 B.n192 10.6151
R1088 B.n193 B.n0 10.6151
R1089 B.n739 B.n1 10.6151
R1090 B.n739 B.n738 10.6151
R1091 B.n738 B.n737 10.6151
R1092 B.n737 B.n4 10.6151
R1093 B.n733 B.n4 10.6151
R1094 B.n733 B.n732 10.6151
R1095 B.n732 B.n731 10.6151
R1096 B.n731 B.n6 10.6151
R1097 B.n727 B.n6 10.6151
R1098 B.n727 B.n726 10.6151
R1099 B.n726 B.n725 10.6151
R1100 B.n725 B.n8 10.6151
R1101 B.n721 B.n8 10.6151
R1102 B.n721 B.n720 10.6151
R1103 B.n720 B.n719 10.6151
R1104 B.n719 B.n10 10.6151
R1105 B.n715 B.n10 10.6151
R1106 B.n715 B.n714 10.6151
R1107 B.n714 B.n713 10.6151
R1108 B.n713 B.n12 10.6151
R1109 B.n709 B.n12 10.6151
R1110 B.n709 B.n708 10.6151
R1111 B.n708 B.n707 10.6151
R1112 B.n707 B.n14 10.6151
R1113 B.n613 B.n612 9.36635
R1114 B.n595 B.n54 9.36635
R1115 B.n319 B.n150 9.36635
R1116 B.n337 B.n336 9.36635
R1117 B.n743 B.n0 2.81026
R1118 B.n743 B.n1 2.81026
R1119 B.n612 B.n611 1.24928
R1120 B.n598 B.n54 1.24928
R1121 B.n322 B.n150 1.24928
R1122 B.n336 B.n335 1.24928
R1123 VN VN.t1 275.906
R1124 VN VN.t0 226.524
R1125 VTAIL.n414 VTAIL.n413 756.745
R1126 VTAIL.n102 VTAIL.n101 756.745
R1127 VTAIL.n310 VTAIL.n309 756.745
R1128 VTAIL.n206 VTAIL.n205 756.745
R1129 VTAIL.n347 VTAIL.n346 585
R1130 VTAIL.n349 VTAIL.n348 585
R1131 VTAIL.n342 VTAIL.n341 585
R1132 VTAIL.n355 VTAIL.n354 585
R1133 VTAIL.n357 VTAIL.n356 585
R1134 VTAIL.n338 VTAIL.n337 585
R1135 VTAIL.n364 VTAIL.n363 585
R1136 VTAIL.n365 VTAIL.n336 585
R1137 VTAIL.n367 VTAIL.n366 585
R1138 VTAIL.n334 VTAIL.n333 585
R1139 VTAIL.n373 VTAIL.n372 585
R1140 VTAIL.n375 VTAIL.n374 585
R1141 VTAIL.n330 VTAIL.n329 585
R1142 VTAIL.n381 VTAIL.n380 585
R1143 VTAIL.n383 VTAIL.n382 585
R1144 VTAIL.n326 VTAIL.n325 585
R1145 VTAIL.n389 VTAIL.n388 585
R1146 VTAIL.n391 VTAIL.n390 585
R1147 VTAIL.n322 VTAIL.n321 585
R1148 VTAIL.n397 VTAIL.n396 585
R1149 VTAIL.n399 VTAIL.n398 585
R1150 VTAIL.n318 VTAIL.n317 585
R1151 VTAIL.n405 VTAIL.n404 585
R1152 VTAIL.n407 VTAIL.n406 585
R1153 VTAIL.n314 VTAIL.n313 585
R1154 VTAIL.n413 VTAIL.n412 585
R1155 VTAIL.n35 VTAIL.n34 585
R1156 VTAIL.n37 VTAIL.n36 585
R1157 VTAIL.n30 VTAIL.n29 585
R1158 VTAIL.n43 VTAIL.n42 585
R1159 VTAIL.n45 VTAIL.n44 585
R1160 VTAIL.n26 VTAIL.n25 585
R1161 VTAIL.n52 VTAIL.n51 585
R1162 VTAIL.n53 VTAIL.n24 585
R1163 VTAIL.n55 VTAIL.n54 585
R1164 VTAIL.n22 VTAIL.n21 585
R1165 VTAIL.n61 VTAIL.n60 585
R1166 VTAIL.n63 VTAIL.n62 585
R1167 VTAIL.n18 VTAIL.n17 585
R1168 VTAIL.n69 VTAIL.n68 585
R1169 VTAIL.n71 VTAIL.n70 585
R1170 VTAIL.n14 VTAIL.n13 585
R1171 VTAIL.n77 VTAIL.n76 585
R1172 VTAIL.n79 VTAIL.n78 585
R1173 VTAIL.n10 VTAIL.n9 585
R1174 VTAIL.n85 VTAIL.n84 585
R1175 VTAIL.n87 VTAIL.n86 585
R1176 VTAIL.n6 VTAIL.n5 585
R1177 VTAIL.n93 VTAIL.n92 585
R1178 VTAIL.n95 VTAIL.n94 585
R1179 VTAIL.n2 VTAIL.n1 585
R1180 VTAIL.n101 VTAIL.n100 585
R1181 VTAIL.n309 VTAIL.n308 585
R1182 VTAIL.n210 VTAIL.n209 585
R1183 VTAIL.n303 VTAIL.n302 585
R1184 VTAIL.n301 VTAIL.n300 585
R1185 VTAIL.n214 VTAIL.n213 585
R1186 VTAIL.n295 VTAIL.n294 585
R1187 VTAIL.n293 VTAIL.n292 585
R1188 VTAIL.n218 VTAIL.n217 585
R1189 VTAIL.n287 VTAIL.n286 585
R1190 VTAIL.n285 VTAIL.n284 585
R1191 VTAIL.n222 VTAIL.n221 585
R1192 VTAIL.n279 VTAIL.n278 585
R1193 VTAIL.n277 VTAIL.n276 585
R1194 VTAIL.n226 VTAIL.n225 585
R1195 VTAIL.n271 VTAIL.n270 585
R1196 VTAIL.n269 VTAIL.n268 585
R1197 VTAIL.n230 VTAIL.n229 585
R1198 VTAIL.n234 VTAIL.n232 585
R1199 VTAIL.n263 VTAIL.n262 585
R1200 VTAIL.n261 VTAIL.n260 585
R1201 VTAIL.n236 VTAIL.n235 585
R1202 VTAIL.n255 VTAIL.n254 585
R1203 VTAIL.n253 VTAIL.n252 585
R1204 VTAIL.n240 VTAIL.n239 585
R1205 VTAIL.n247 VTAIL.n246 585
R1206 VTAIL.n245 VTAIL.n244 585
R1207 VTAIL.n205 VTAIL.n204 585
R1208 VTAIL.n106 VTAIL.n105 585
R1209 VTAIL.n199 VTAIL.n198 585
R1210 VTAIL.n197 VTAIL.n196 585
R1211 VTAIL.n110 VTAIL.n109 585
R1212 VTAIL.n191 VTAIL.n190 585
R1213 VTAIL.n189 VTAIL.n188 585
R1214 VTAIL.n114 VTAIL.n113 585
R1215 VTAIL.n183 VTAIL.n182 585
R1216 VTAIL.n181 VTAIL.n180 585
R1217 VTAIL.n118 VTAIL.n117 585
R1218 VTAIL.n175 VTAIL.n174 585
R1219 VTAIL.n173 VTAIL.n172 585
R1220 VTAIL.n122 VTAIL.n121 585
R1221 VTAIL.n167 VTAIL.n166 585
R1222 VTAIL.n165 VTAIL.n164 585
R1223 VTAIL.n126 VTAIL.n125 585
R1224 VTAIL.n130 VTAIL.n128 585
R1225 VTAIL.n159 VTAIL.n158 585
R1226 VTAIL.n157 VTAIL.n156 585
R1227 VTAIL.n132 VTAIL.n131 585
R1228 VTAIL.n151 VTAIL.n150 585
R1229 VTAIL.n149 VTAIL.n148 585
R1230 VTAIL.n136 VTAIL.n135 585
R1231 VTAIL.n143 VTAIL.n142 585
R1232 VTAIL.n141 VTAIL.n140 585
R1233 VTAIL.n345 VTAIL.t2 329.036
R1234 VTAIL.n33 VTAIL.t0 329.036
R1235 VTAIL.n243 VTAIL.t1 329.036
R1236 VTAIL.n139 VTAIL.t3 329.036
R1237 VTAIL.n348 VTAIL.n347 171.744
R1238 VTAIL.n348 VTAIL.n341 171.744
R1239 VTAIL.n355 VTAIL.n341 171.744
R1240 VTAIL.n356 VTAIL.n355 171.744
R1241 VTAIL.n356 VTAIL.n337 171.744
R1242 VTAIL.n364 VTAIL.n337 171.744
R1243 VTAIL.n365 VTAIL.n364 171.744
R1244 VTAIL.n366 VTAIL.n365 171.744
R1245 VTAIL.n366 VTAIL.n333 171.744
R1246 VTAIL.n373 VTAIL.n333 171.744
R1247 VTAIL.n374 VTAIL.n373 171.744
R1248 VTAIL.n374 VTAIL.n329 171.744
R1249 VTAIL.n381 VTAIL.n329 171.744
R1250 VTAIL.n382 VTAIL.n381 171.744
R1251 VTAIL.n382 VTAIL.n325 171.744
R1252 VTAIL.n389 VTAIL.n325 171.744
R1253 VTAIL.n390 VTAIL.n389 171.744
R1254 VTAIL.n390 VTAIL.n321 171.744
R1255 VTAIL.n397 VTAIL.n321 171.744
R1256 VTAIL.n398 VTAIL.n397 171.744
R1257 VTAIL.n398 VTAIL.n317 171.744
R1258 VTAIL.n405 VTAIL.n317 171.744
R1259 VTAIL.n406 VTAIL.n405 171.744
R1260 VTAIL.n406 VTAIL.n313 171.744
R1261 VTAIL.n413 VTAIL.n313 171.744
R1262 VTAIL.n36 VTAIL.n35 171.744
R1263 VTAIL.n36 VTAIL.n29 171.744
R1264 VTAIL.n43 VTAIL.n29 171.744
R1265 VTAIL.n44 VTAIL.n43 171.744
R1266 VTAIL.n44 VTAIL.n25 171.744
R1267 VTAIL.n52 VTAIL.n25 171.744
R1268 VTAIL.n53 VTAIL.n52 171.744
R1269 VTAIL.n54 VTAIL.n53 171.744
R1270 VTAIL.n54 VTAIL.n21 171.744
R1271 VTAIL.n61 VTAIL.n21 171.744
R1272 VTAIL.n62 VTAIL.n61 171.744
R1273 VTAIL.n62 VTAIL.n17 171.744
R1274 VTAIL.n69 VTAIL.n17 171.744
R1275 VTAIL.n70 VTAIL.n69 171.744
R1276 VTAIL.n70 VTAIL.n13 171.744
R1277 VTAIL.n77 VTAIL.n13 171.744
R1278 VTAIL.n78 VTAIL.n77 171.744
R1279 VTAIL.n78 VTAIL.n9 171.744
R1280 VTAIL.n85 VTAIL.n9 171.744
R1281 VTAIL.n86 VTAIL.n85 171.744
R1282 VTAIL.n86 VTAIL.n5 171.744
R1283 VTAIL.n93 VTAIL.n5 171.744
R1284 VTAIL.n94 VTAIL.n93 171.744
R1285 VTAIL.n94 VTAIL.n1 171.744
R1286 VTAIL.n101 VTAIL.n1 171.744
R1287 VTAIL.n309 VTAIL.n209 171.744
R1288 VTAIL.n302 VTAIL.n209 171.744
R1289 VTAIL.n302 VTAIL.n301 171.744
R1290 VTAIL.n301 VTAIL.n213 171.744
R1291 VTAIL.n294 VTAIL.n213 171.744
R1292 VTAIL.n294 VTAIL.n293 171.744
R1293 VTAIL.n293 VTAIL.n217 171.744
R1294 VTAIL.n286 VTAIL.n217 171.744
R1295 VTAIL.n286 VTAIL.n285 171.744
R1296 VTAIL.n285 VTAIL.n221 171.744
R1297 VTAIL.n278 VTAIL.n221 171.744
R1298 VTAIL.n278 VTAIL.n277 171.744
R1299 VTAIL.n277 VTAIL.n225 171.744
R1300 VTAIL.n270 VTAIL.n225 171.744
R1301 VTAIL.n270 VTAIL.n269 171.744
R1302 VTAIL.n269 VTAIL.n229 171.744
R1303 VTAIL.n234 VTAIL.n229 171.744
R1304 VTAIL.n262 VTAIL.n234 171.744
R1305 VTAIL.n262 VTAIL.n261 171.744
R1306 VTAIL.n261 VTAIL.n235 171.744
R1307 VTAIL.n254 VTAIL.n235 171.744
R1308 VTAIL.n254 VTAIL.n253 171.744
R1309 VTAIL.n253 VTAIL.n239 171.744
R1310 VTAIL.n246 VTAIL.n239 171.744
R1311 VTAIL.n246 VTAIL.n245 171.744
R1312 VTAIL.n205 VTAIL.n105 171.744
R1313 VTAIL.n198 VTAIL.n105 171.744
R1314 VTAIL.n198 VTAIL.n197 171.744
R1315 VTAIL.n197 VTAIL.n109 171.744
R1316 VTAIL.n190 VTAIL.n109 171.744
R1317 VTAIL.n190 VTAIL.n189 171.744
R1318 VTAIL.n189 VTAIL.n113 171.744
R1319 VTAIL.n182 VTAIL.n113 171.744
R1320 VTAIL.n182 VTAIL.n181 171.744
R1321 VTAIL.n181 VTAIL.n117 171.744
R1322 VTAIL.n174 VTAIL.n117 171.744
R1323 VTAIL.n174 VTAIL.n173 171.744
R1324 VTAIL.n173 VTAIL.n121 171.744
R1325 VTAIL.n166 VTAIL.n121 171.744
R1326 VTAIL.n166 VTAIL.n165 171.744
R1327 VTAIL.n165 VTAIL.n125 171.744
R1328 VTAIL.n130 VTAIL.n125 171.744
R1329 VTAIL.n158 VTAIL.n130 171.744
R1330 VTAIL.n158 VTAIL.n157 171.744
R1331 VTAIL.n157 VTAIL.n131 171.744
R1332 VTAIL.n150 VTAIL.n131 171.744
R1333 VTAIL.n150 VTAIL.n149 171.744
R1334 VTAIL.n149 VTAIL.n135 171.744
R1335 VTAIL.n142 VTAIL.n135 171.744
R1336 VTAIL.n142 VTAIL.n141 171.744
R1337 VTAIL.n347 VTAIL.t2 85.8723
R1338 VTAIL.n35 VTAIL.t0 85.8723
R1339 VTAIL.n245 VTAIL.t1 85.8723
R1340 VTAIL.n141 VTAIL.t3 85.8723
R1341 VTAIL.n415 VTAIL.n414 34.3187
R1342 VTAIL.n103 VTAIL.n102 34.3187
R1343 VTAIL.n311 VTAIL.n310 34.3187
R1344 VTAIL.n207 VTAIL.n206 34.3187
R1345 VTAIL.n207 VTAIL.n103 33.479
R1346 VTAIL.n415 VTAIL.n311 30.9962
R1347 VTAIL.n367 VTAIL.n334 13.1884
R1348 VTAIL.n55 VTAIL.n22 13.1884
R1349 VTAIL.n232 VTAIL.n230 13.1884
R1350 VTAIL.n128 VTAIL.n126 13.1884
R1351 VTAIL.n368 VTAIL.n336 12.8005
R1352 VTAIL.n372 VTAIL.n371 12.8005
R1353 VTAIL.n412 VTAIL.n312 12.8005
R1354 VTAIL.n56 VTAIL.n24 12.8005
R1355 VTAIL.n60 VTAIL.n59 12.8005
R1356 VTAIL.n100 VTAIL.n0 12.8005
R1357 VTAIL.n308 VTAIL.n208 12.8005
R1358 VTAIL.n268 VTAIL.n267 12.8005
R1359 VTAIL.n264 VTAIL.n263 12.8005
R1360 VTAIL.n204 VTAIL.n104 12.8005
R1361 VTAIL.n164 VTAIL.n163 12.8005
R1362 VTAIL.n160 VTAIL.n159 12.8005
R1363 VTAIL.n363 VTAIL.n362 12.0247
R1364 VTAIL.n375 VTAIL.n332 12.0247
R1365 VTAIL.n411 VTAIL.n314 12.0247
R1366 VTAIL.n51 VTAIL.n50 12.0247
R1367 VTAIL.n63 VTAIL.n20 12.0247
R1368 VTAIL.n99 VTAIL.n2 12.0247
R1369 VTAIL.n307 VTAIL.n210 12.0247
R1370 VTAIL.n271 VTAIL.n228 12.0247
R1371 VTAIL.n260 VTAIL.n233 12.0247
R1372 VTAIL.n203 VTAIL.n106 12.0247
R1373 VTAIL.n167 VTAIL.n124 12.0247
R1374 VTAIL.n156 VTAIL.n129 12.0247
R1375 VTAIL.n361 VTAIL.n338 11.249
R1376 VTAIL.n376 VTAIL.n330 11.249
R1377 VTAIL.n408 VTAIL.n407 11.249
R1378 VTAIL.n49 VTAIL.n26 11.249
R1379 VTAIL.n64 VTAIL.n18 11.249
R1380 VTAIL.n96 VTAIL.n95 11.249
R1381 VTAIL.n304 VTAIL.n303 11.249
R1382 VTAIL.n272 VTAIL.n226 11.249
R1383 VTAIL.n259 VTAIL.n236 11.249
R1384 VTAIL.n200 VTAIL.n199 11.249
R1385 VTAIL.n168 VTAIL.n122 11.249
R1386 VTAIL.n155 VTAIL.n132 11.249
R1387 VTAIL.n346 VTAIL.n345 10.7239
R1388 VTAIL.n34 VTAIL.n33 10.7239
R1389 VTAIL.n244 VTAIL.n243 10.7239
R1390 VTAIL.n140 VTAIL.n139 10.7239
R1391 VTAIL.n358 VTAIL.n357 10.4732
R1392 VTAIL.n380 VTAIL.n379 10.4732
R1393 VTAIL.n404 VTAIL.n316 10.4732
R1394 VTAIL.n46 VTAIL.n45 10.4732
R1395 VTAIL.n68 VTAIL.n67 10.4732
R1396 VTAIL.n92 VTAIL.n4 10.4732
R1397 VTAIL.n300 VTAIL.n212 10.4732
R1398 VTAIL.n276 VTAIL.n275 10.4732
R1399 VTAIL.n256 VTAIL.n255 10.4732
R1400 VTAIL.n196 VTAIL.n108 10.4732
R1401 VTAIL.n172 VTAIL.n171 10.4732
R1402 VTAIL.n152 VTAIL.n151 10.4732
R1403 VTAIL.n354 VTAIL.n340 9.69747
R1404 VTAIL.n383 VTAIL.n328 9.69747
R1405 VTAIL.n403 VTAIL.n318 9.69747
R1406 VTAIL.n42 VTAIL.n28 9.69747
R1407 VTAIL.n71 VTAIL.n16 9.69747
R1408 VTAIL.n91 VTAIL.n6 9.69747
R1409 VTAIL.n299 VTAIL.n214 9.69747
R1410 VTAIL.n279 VTAIL.n224 9.69747
R1411 VTAIL.n252 VTAIL.n238 9.69747
R1412 VTAIL.n195 VTAIL.n110 9.69747
R1413 VTAIL.n175 VTAIL.n120 9.69747
R1414 VTAIL.n148 VTAIL.n134 9.69747
R1415 VTAIL.n410 VTAIL.n312 9.45567
R1416 VTAIL.n98 VTAIL.n0 9.45567
R1417 VTAIL.n306 VTAIL.n208 9.45567
R1418 VTAIL.n202 VTAIL.n104 9.45567
R1419 VTAIL.n393 VTAIL.n392 9.3005
R1420 VTAIL.n395 VTAIL.n394 9.3005
R1421 VTAIL.n320 VTAIL.n319 9.3005
R1422 VTAIL.n401 VTAIL.n400 9.3005
R1423 VTAIL.n403 VTAIL.n402 9.3005
R1424 VTAIL.n316 VTAIL.n315 9.3005
R1425 VTAIL.n409 VTAIL.n408 9.3005
R1426 VTAIL.n411 VTAIL.n410 9.3005
R1427 VTAIL.n387 VTAIL.n386 9.3005
R1428 VTAIL.n385 VTAIL.n384 9.3005
R1429 VTAIL.n328 VTAIL.n327 9.3005
R1430 VTAIL.n379 VTAIL.n378 9.3005
R1431 VTAIL.n377 VTAIL.n376 9.3005
R1432 VTAIL.n332 VTAIL.n331 9.3005
R1433 VTAIL.n371 VTAIL.n370 9.3005
R1434 VTAIL.n344 VTAIL.n343 9.3005
R1435 VTAIL.n351 VTAIL.n350 9.3005
R1436 VTAIL.n353 VTAIL.n352 9.3005
R1437 VTAIL.n340 VTAIL.n339 9.3005
R1438 VTAIL.n359 VTAIL.n358 9.3005
R1439 VTAIL.n361 VTAIL.n360 9.3005
R1440 VTAIL.n362 VTAIL.n335 9.3005
R1441 VTAIL.n369 VTAIL.n368 9.3005
R1442 VTAIL.n324 VTAIL.n323 9.3005
R1443 VTAIL.n81 VTAIL.n80 9.3005
R1444 VTAIL.n83 VTAIL.n82 9.3005
R1445 VTAIL.n8 VTAIL.n7 9.3005
R1446 VTAIL.n89 VTAIL.n88 9.3005
R1447 VTAIL.n91 VTAIL.n90 9.3005
R1448 VTAIL.n4 VTAIL.n3 9.3005
R1449 VTAIL.n97 VTAIL.n96 9.3005
R1450 VTAIL.n99 VTAIL.n98 9.3005
R1451 VTAIL.n75 VTAIL.n74 9.3005
R1452 VTAIL.n73 VTAIL.n72 9.3005
R1453 VTAIL.n16 VTAIL.n15 9.3005
R1454 VTAIL.n67 VTAIL.n66 9.3005
R1455 VTAIL.n65 VTAIL.n64 9.3005
R1456 VTAIL.n20 VTAIL.n19 9.3005
R1457 VTAIL.n59 VTAIL.n58 9.3005
R1458 VTAIL.n32 VTAIL.n31 9.3005
R1459 VTAIL.n39 VTAIL.n38 9.3005
R1460 VTAIL.n41 VTAIL.n40 9.3005
R1461 VTAIL.n28 VTAIL.n27 9.3005
R1462 VTAIL.n47 VTAIL.n46 9.3005
R1463 VTAIL.n49 VTAIL.n48 9.3005
R1464 VTAIL.n50 VTAIL.n23 9.3005
R1465 VTAIL.n57 VTAIL.n56 9.3005
R1466 VTAIL.n12 VTAIL.n11 9.3005
R1467 VTAIL.n307 VTAIL.n306 9.3005
R1468 VTAIL.n305 VTAIL.n304 9.3005
R1469 VTAIL.n212 VTAIL.n211 9.3005
R1470 VTAIL.n299 VTAIL.n298 9.3005
R1471 VTAIL.n297 VTAIL.n296 9.3005
R1472 VTAIL.n216 VTAIL.n215 9.3005
R1473 VTAIL.n291 VTAIL.n290 9.3005
R1474 VTAIL.n289 VTAIL.n288 9.3005
R1475 VTAIL.n220 VTAIL.n219 9.3005
R1476 VTAIL.n283 VTAIL.n282 9.3005
R1477 VTAIL.n281 VTAIL.n280 9.3005
R1478 VTAIL.n224 VTAIL.n223 9.3005
R1479 VTAIL.n275 VTAIL.n274 9.3005
R1480 VTAIL.n273 VTAIL.n272 9.3005
R1481 VTAIL.n228 VTAIL.n227 9.3005
R1482 VTAIL.n267 VTAIL.n266 9.3005
R1483 VTAIL.n265 VTAIL.n264 9.3005
R1484 VTAIL.n233 VTAIL.n231 9.3005
R1485 VTAIL.n259 VTAIL.n258 9.3005
R1486 VTAIL.n257 VTAIL.n256 9.3005
R1487 VTAIL.n238 VTAIL.n237 9.3005
R1488 VTAIL.n251 VTAIL.n250 9.3005
R1489 VTAIL.n249 VTAIL.n248 9.3005
R1490 VTAIL.n242 VTAIL.n241 9.3005
R1491 VTAIL.n138 VTAIL.n137 9.3005
R1492 VTAIL.n145 VTAIL.n144 9.3005
R1493 VTAIL.n147 VTAIL.n146 9.3005
R1494 VTAIL.n134 VTAIL.n133 9.3005
R1495 VTAIL.n153 VTAIL.n152 9.3005
R1496 VTAIL.n155 VTAIL.n154 9.3005
R1497 VTAIL.n129 VTAIL.n127 9.3005
R1498 VTAIL.n161 VTAIL.n160 9.3005
R1499 VTAIL.n187 VTAIL.n186 9.3005
R1500 VTAIL.n112 VTAIL.n111 9.3005
R1501 VTAIL.n193 VTAIL.n192 9.3005
R1502 VTAIL.n195 VTAIL.n194 9.3005
R1503 VTAIL.n108 VTAIL.n107 9.3005
R1504 VTAIL.n201 VTAIL.n200 9.3005
R1505 VTAIL.n203 VTAIL.n202 9.3005
R1506 VTAIL.n185 VTAIL.n184 9.3005
R1507 VTAIL.n116 VTAIL.n115 9.3005
R1508 VTAIL.n179 VTAIL.n178 9.3005
R1509 VTAIL.n177 VTAIL.n176 9.3005
R1510 VTAIL.n120 VTAIL.n119 9.3005
R1511 VTAIL.n171 VTAIL.n170 9.3005
R1512 VTAIL.n169 VTAIL.n168 9.3005
R1513 VTAIL.n124 VTAIL.n123 9.3005
R1514 VTAIL.n163 VTAIL.n162 9.3005
R1515 VTAIL.n353 VTAIL.n342 8.92171
R1516 VTAIL.n384 VTAIL.n326 8.92171
R1517 VTAIL.n400 VTAIL.n399 8.92171
R1518 VTAIL.n41 VTAIL.n30 8.92171
R1519 VTAIL.n72 VTAIL.n14 8.92171
R1520 VTAIL.n88 VTAIL.n87 8.92171
R1521 VTAIL.n296 VTAIL.n295 8.92171
R1522 VTAIL.n280 VTAIL.n222 8.92171
R1523 VTAIL.n251 VTAIL.n240 8.92171
R1524 VTAIL.n192 VTAIL.n191 8.92171
R1525 VTAIL.n176 VTAIL.n118 8.92171
R1526 VTAIL.n147 VTAIL.n136 8.92171
R1527 VTAIL.n350 VTAIL.n349 8.14595
R1528 VTAIL.n388 VTAIL.n387 8.14595
R1529 VTAIL.n396 VTAIL.n320 8.14595
R1530 VTAIL.n38 VTAIL.n37 8.14595
R1531 VTAIL.n76 VTAIL.n75 8.14595
R1532 VTAIL.n84 VTAIL.n8 8.14595
R1533 VTAIL.n292 VTAIL.n216 8.14595
R1534 VTAIL.n284 VTAIL.n283 8.14595
R1535 VTAIL.n248 VTAIL.n247 8.14595
R1536 VTAIL.n188 VTAIL.n112 8.14595
R1537 VTAIL.n180 VTAIL.n179 8.14595
R1538 VTAIL.n144 VTAIL.n143 8.14595
R1539 VTAIL.n346 VTAIL.n344 7.3702
R1540 VTAIL.n391 VTAIL.n324 7.3702
R1541 VTAIL.n395 VTAIL.n322 7.3702
R1542 VTAIL.n34 VTAIL.n32 7.3702
R1543 VTAIL.n79 VTAIL.n12 7.3702
R1544 VTAIL.n83 VTAIL.n10 7.3702
R1545 VTAIL.n291 VTAIL.n218 7.3702
R1546 VTAIL.n287 VTAIL.n220 7.3702
R1547 VTAIL.n244 VTAIL.n242 7.3702
R1548 VTAIL.n187 VTAIL.n114 7.3702
R1549 VTAIL.n183 VTAIL.n116 7.3702
R1550 VTAIL.n140 VTAIL.n138 7.3702
R1551 VTAIL.n392 VTAIL.n391 6.59444
R1552 VTAIL.n392 VTAIL.n322 6.59444
R1553 VTAIL.n80 VTAIL.n79 6.59444
R1554 VTAIL.n80 VTAIL.n10 6.59444
R1555 VTAIL.n288 VTAIL.n218 6.59444
R1556 VTAIL.n288 VTAIL.n287 6.59444
R1557 VTAIL.n184 VTAIL.n114 6.59444
R1558 VTAIL.n184 VTAIL.n183 6.59444
R1559 VTAIL.n349 VTAIL.n344 5.81868
R1560 VTAIL.n388 VTAIL.n324 5.81868
R1561 VTAIL.n396 VTAIL.n395 5.81868
R1562 VTAIL.n37 VTAIL.n32 5.81868
R1563 VTAIL.n76 VTAIL.n12 5.81868
R1564 VTAIL.n84 VTAIL.n83 5.81868
R1565 VTAIL.n292 VTAIL.n291 5.81868
R1566 VTAIL.n284 VTAIL.n220 5.81868
R1567 VTAIL.n247 VTAIL.n242 5.81868
R1568 VTAIL.n188 VTAIL.n187 5.81868
R1569 VTAIL.n180 VTAIL.n116 5.81868
R1570 VTAIL.n143 VTAIL.n138 5.81868
R1571 VTAIL.n350 VTAIL.n342 5.04292
R1572 VTAIL.n387 VTAIL.n326 5.04292
R1573 VTAIL.n399 VTAIL.n320 5.04292
R1574 VTAIL.n38 VTAIL.n30 5.04292
R1575 VTAIL.n75 VTAIL.n14 5.04292
R1576 VTAIL.n87 VTAIL.n8 5.04292
R1577 VTAIL.n295 VTAIL.n216 5.04292
R1578 VTAIL.n283 VTAIL.n222 5.04292
R1579 VTAIL.n248 VTAIL.n240 5.04292
R1580 VTAIL.n191 VTAIL.n112 5.04292
R1581 VTAIL.n179 VTAIL.n118 5.04292
R1582 VTAIL.n144 VTAIL.n136 5.04292
R1583 VTAIL.n354 VTAIL.n353 4.26717
R1584 VTAIL.n384 VTAIL.n383 4.26717
R1585 VTAIL.n400 VTAIL.n318 4.26717
R1586 VTAIL.n42 VTAIL.n41 4.26717
R1587 VTAIL.n72 VTAIL.n71 4.26717
R1588 VTAIL.n88 VTAIL.n6 4.26717
R1589 VTAIL.n296 VTAIL.n214 4.26717
R1590 VTAIL.n280 VTAIL.n279 4.26717
R1591 VTAIL.n252 VTAIL.n251 4.26717
R1592 VTAIL.n192 VTAIL.n110 4.26717
R1593 VTAIL.n176 VTAIL.n175 4.26717
R1594 VTAIL.n148 VTAIL.n147 4.26717
R1595 VTAIL.n357 VTAIL.n340 3.49141
R1596 VTAIL.n380 VTAIL.n328 3.49141
R1597 VTAIL.n404 VTAIL.n403 3.49141
R1598 VTAIL.n45 VTAIL.n28 3.49141
R1599 VTAIL.n68 VTAIL.n16 3.49141
R1600 VTAIL.n92 VTAIL.n91 3.49141
R1601 VTAIL.n300 VTAIL.n299 3.49141
R1602 VTAIL.n276 VTAIL.n224 3.49141
R1603 VTAIL.n255 VTAIL.n238 3.49141
R1604 VTAIL.n196 VTAIL.n195 3.49141
R1605 VTAIL.n172 VTAIL.n120 3.49141
R1606 VTAIL.n151 VTAIL.n134 3.49141
R1607 VTAIL.n358 VTAIL.n338 2.71565
R1608 VTAIL.n379 VTAIL.n330 2.71565
R1609 VTAIL.n407 VTAIL.n316 2.71565
R1610 VTAIL.n46 VTAIL.n26 2.71565
R1611 VTAIL.n67 VTAIL.n18 2.71565
R1612 VTAIL.n95 VTAIL.n4 2.71565
R1613 VTAIL.n303 VTAIL.n212 2.71565
R1614 VTAIL.n275 VTAIL.n226 2.71565
R1615 VTAIL.n256 VTAIL.n236 2.71565
R1616 VTAIL.n199 VTAIL.n108 2.71565
R1617 VTAIL.n171 VTAIL.n122 2.71565
R1618 VTAIL.n152 VTAIL.n132 2.71565
R1619 VTAIL.n243 VTAIL.n241 2.41282
R1620 VTAIL.n139 VTAIL.n137 2.41282
R1621 VTAIL.n345 VTAIL.n343 2.41282
R1622 VTAIL.n33 VTAIL.n31 2.41282
R1623 VTAIL.n363 VTAIL.n361 1.93989
R1624 VTAIL.n376 VTAIL.n375 1.93989
R1625 VTAIL.n408 VTAIL.n314 1.93989
R1626 VTAIL.n51 VTAIL.n49 1.93989
R1627 VTAIL.n64 VTAIL.n63 1.93989
R1628 VTAIL.n96 VTAIL.n2 1.93989
R1629 VTAIL.n304 VTAIL.n210 1.93989
R1630 VTAIL.n272 VTAIL.n271 1.93989
R1631 VTAIL.n260 VTAIL.n259 1.93989
R1632 VTAIL.n200 VTAIL.n106 1.93989
R1633 VTAIL.n168 VTAIL.n167 1.93989
R1634 VTAIL.n156 VTAIL.n155 1.93989
R1635 VTAIL.n311 VTAIL.n207 1.71171
R1636 VTAIL.n362 VTAIL.n336 1.16414
R1637 VTAIL.n372 VTAIL.n332 1.16414
R1638 VTAIL.n412 VTAIL.n411 1.16414
R1639 VTAIL.n50 VTAIL.n24 1.16414
R1640 VTAIL.n60 VTAIL.n20 1.16414
R1641 VTAIL.n100 VTAIL.n99 1.16414
R1642 VTAIL.n308 VTAIL.n307 1.16414
R1643 VTAIL.n268 VTAIL.n228 1.16414
R1644 VTAIL.n263 VTAIL.n233 1.16414
R1645 VTAIL.n204 VTAIL.n203 1.16414
R1646 VTAIL.n164 VTAIL.n124 1.16414
R1647 VTAIL.n159 VTAIL.n129 1.16414
R1648 VTAIL VTAIL.n103 1.14921
R1649 VTAIL VTAIL.n415 0.563
R1650 VTAIL.n368 VTAIL.n367 0.388379
R1651 VTAIL.n371 VTAIL.n334 0.388379
R1652 VTAIL.n414 VTAIL.n312 0.388379
R1653 VTAIL.n56 VTAIL.n55 0.388379
R1654 VTAIL.n59 VTAIL.n22 0.388379
R1655 VTAIL.n102 VTAIL.n0 0.388379
R1656 VTAIL.n310 VTAIL.n208 0.388379
R1657 VTAIL.n267 VTAIL.n230 0.388379
R1658 VTAIL.n264 VTAIL.n232 0.388379
R1659 VTAIL.n206 VTAIL.n104 0.388379
R1660 VTAIL.n163 VTAIL.n126 0.388379
R1661 VTAIL.n160 VTAIL.n128 0.388379
R1662 VTAIL.n351 VTAIL.n343 0.155672
R1663 VTAIL.n352 VTAIL.n351 0.155672
R1664 VTAIL.n352 VTAIL.n339 0.155672
R1665 VTAIL.n359 VTAIL.n339 0.155672
R1666 VTAIL.n360 VTAIL.n359 0.155672
R1667 VTAIL.n360 VTAIL.n335 0.155672
R1668 VTAIL.n369 VTAIL.n335 0.155672
R1669 VTAIL.n370 VTAIL.n369 0.155672
R1670 VTAIL.n370 VTAIL.n331 0.155672
R1671 VTAIL.n377 VTAIL.n331 0.155672
R1672 VTAIL.n378 VTAIL.n377 0.155672
R1673 VTAIL.n378 VTAIL.n327 0.155672
R1674 VTAIL.n385 VTAIL.n327 0.155672
R1675 VTAIL.n386 VTAIL.n385 0.155672
R1676 VTAIL.n386 VTAIL.n323 0.155672
R1677 VTAIL.n393 VTAIL.n323 0.155672
R1678 VTAIL.n394 VTAIL.n393 0.155672
R1679 VTAIL.n394 VTAIL.n319 0.155672
R1680 VTAIL.n401 VTAIL.n319 0.155672
R1681 VTAIL.n402 VTAIL.n401 0.155672
R1682 VTAIL.n402 VTAIL.n315 0.155672
R1683 VTAIL.n409 VTAIL.n315 0.155672
R1684 VTAIL.n410 VTAIL.n409 0.155672
R1685 VTAIL.n39 VTAIL.n31 0.155672
R1686 VTAIL.n40 VTAIL.n39 0.155672
R1687 VTAIL.n40 VTAIL.n27 0.155672
R1688 VTAIL.n47 VTAIL.n27 0.155672
R1689 VTAIL.n48 VTAIL.n47 0.155672
R1690 VTAIL.n48 VTAIL.n23 0.155672
R1691 VTAIL.n57 VTAIL.n23 0.155672
R1692 VTAIL.n58 VTAIL.n57 0.155672
R1693 VTAIL.n58 VTAIL.n19 0.155672
R1694 VTAIL.n65 VTAIL.n19 0.155672
R1695 VTAIL.n66 VTAIL.n65 0.155672
R1696 VTAIL.n66 VTAIL.n15 0.155672
R1697 VTAIL.n73 VTAIL.n15 0.155672
R1698 VTAIL.n74 VTAIL.n73 0.155672
R1699 VTAIL.n74 VTAIL.n11 0.155672
R1700 VTAIL.n81 VTAIL.n11 0.155672
R1701 VTAIL.n82 VTAIL.n81 0.155672
R1702 VTAIL.n82 VTAIL.n7 0.155672
R1703 VTAIL.n89 VTAIL.n7 0.155672
R1704 VTAIL.n90 VTAIL.n89 0.155672
R1705 VTAIL.n90 VTAIL.n3 0.155672
R1706 VTAIL.n97 VTAIL.n3 0.155672
R1707 VTAIL.n98 VTAIL.n97 0.155672
R1708 VTAIL.n306 VTAIL.n305 0.155672
R1709 VTAIL.n305 VTAIL.n211 0.155672
R1710 VTAIL.n298 VTAIL.n211 0.155672
R1711 VTAIL.n298 VTAIL.n297 0.155672
R1712 VTAIL.n297 VTAIL.n215 0.155672
R1713 VTAIL.n290 VTAIL.n215 0.155672
R1714 VTAIL.n290 VTAIL.n289 0.155672
R1715 VTAIL.n289 VTAIL.n219 0.155672
R1716 VTAIL.n282 VTAIL.n219 0.155672
R1717 VTAIL.n282 VTAIL.n281 0.155672
R1718 VTAIL.n281 VTAIL.n223 0.155672
R1719 VTAIL.n274 VTAIL.n223 0.155672
R1720 VTAIL.n274 VTAIL.n273 0.155672
R1721 VTAIL.n273 VTAIL.n227 0.155672
R1722 VTAIL.n266 VTAIL.n227 0.155672
R1723 VTAIL.n266 VTAIL.n265 0.155672
R1724 VTAIL.n265 VTAIL.n231 0.155672
R1725 VTAIL.n258 VTAIL.n231 0.155672
R1726 VTAIL.n258 VTAIL.n257 0.155672
R1727 VTAIL.n257 VTAIL.n237 0.155672
R1728 VTAIL.n250 VTAIL.n237 0.155672
R1729 VTAIL.n250 VTAIL.n249 0.155672
R1730 VTAIL.n249 VTAIL.n241 0.155672
R1731 VTAIL.n202 VTAIL.n201 0.155672
R1732 VTAIL.n201 VTAIL.n107 0.155672
R1733 VTAIL.n194 VTAIL.n107 0.155672
R1734 VTAIL.n194 VTAIL.n193 0.155672
R1735 VTAIL.n193 VTAIL.n111 0.155672
R1736 VTAIL.n186 VTAIL.n111 0.155672
R1737 VTAIL.n186 VTAIL.n185 0.155672
R1738 VTAIL.n185 VTAIL.n115 0.155672
R1739 VTAIL.n178 VTAIL.n115 0.155672
R1740 VTAIL.n178 VTAIL.n177 0.155672
R1741 VTAIL.n177 VTAIL.n119 0.155672
R1742 VTAIL.n170 VTAIL.n119 0.155672
R1743 VTAIL.n170 VTAIL.n169 0.155672
R1744 VTAIL.n169 VTAIL.n123 0.155672
R1745 VTAIL.n162 VTAIL.n123 0.155672
R1746 VTAIL.n162 VTAIL.n161 0.155672
R1747 VTAIL.n161 VTAIL.n127 0.155672
R1748 VTAIL.n154 VTAIL.n127 0.155672
R1749 VTAIL.n154 VTAIL.n153 0.155672
R1750 VTAIL.n153 VTAIL.n133 0.155672
R1751 VTAIL.n146 VTAIL.n133 0.155672
R1752 VTAIL.n146 VTAIL.n145 0.155672
R1753 VTAIL.n145 VTAIL.n137 0.155672
R1754 VDD2.n205 VDD2.n204 756.745
R1755 VDD2.n102 VDD2.n101 756.745
R1756 VDD2.n204 VDD2.n203 585
R1757 VDD2.n105 VDD2.n104 585
R1758 VDD2.n198 VDD2.n197 585
R1759 VDD2.n196 VDD2.n195 585
R1760 VDD2.n109 VDD2.n108 585
R1761 VDD2.n190 VDD2.n189 585
R1762 VDD2.n188 VDD2.n187 585
R1763 VDD2.n113 VDD2.n112 585
R1764 VDD2.n182 VDD2.n181 585
R1765 VDD2.n180 VDD2.n179 585
R1766 VDD2.n117 VDD2.n116 585
R1767 VDD2.n174 VDD2.n173 585
R1768 VDD2.n172 VDD2.n171 585
R1769 VDD2.n121 VDD2.n120 585
R1770 VDD2.n166 VDD2.n165 585
R1771 VDD2.n164 VDD2.n163 585
R1772 VDD2.n125 VDD2.n124 585
R1773 VDD2.n129 VDD2.n127 585
R1774 VDD2.n158 VDD2.n157 585
R1775 VDD2.n156 VDD2.n155 585
R1776 VDD2.n131 VDD2.n130 585
R1777 VDD2.n150 VDD2.n149 585
R1778 VDD2.n148 VDD2.n147 585
R1779 VDD2.n135 VDD2.n134 585
R1780 VDD2.n142 VDD2.n141 585
R1781 VDD2.n140 VDD2.n139 585
R1782 VDD2.n35 VDD2.n34 585
R1783 VDD2.n37 VDD2.n36 585
R1784 VDD2.n30 VDD2.n29 585
R1785 VDD2.n43 VDD2.n42 585
R1786 VDD2.n45 VDD2.n44 585
R1787 VDD2.n26 VDD2.n25 585
R1788 VDD2.n52 VDD2.n51 585
R1789 VDD2.n53 VDD2.n24 585
R1790 VDD2.n55 VDD2.n54 585
R1791 VDD2.n22 VDD2.n21 585
R1792 VDD2.n61 VDD2.n60 585
R1793 VDD2.n63 VDD2.n62 585
R1794 VDD2.n18 VDD2.n17 585
R1795 VDD2.n69 VDD2.n68 585
R1796 VDD2.n71 VDD2.n70 585
R1797 VDD2.n14 VDD2.n13 585
R1798 VDD2.n77 VDD2.n76 585
R1799 VDD2.n79 VDD2.n78 585
R1800 VDD2.n10 VDD2.n9 585
R1801 VDD2.n85 VDD2.n84 585
R1802 VDD2.n87 VDD2.n86 585
R1803 VDD2.n6 VDD2.n5 585
R1804 VDD2.n93 VDD2.n92 585
R1805 VDD2.n95 VDD2.n94 585
R1806 VDD2.n2 VDD2.n1 585
R1807 VDD2.n101 VDD2.n100 585
R1808 VDD2.n138 VDD2.t0 329.036
R1809 VDD2.n33 VDD2.t1 329.036
R1810 VDD2.n204 VDD2.n104 171.744
R1811 VDD2.n197 VDD2.n104 171.744
R1812 VDD2.n197 VDD2.n196 171.744
R1813 VDD2.n196 VDD2.n108 171.744
R1814 VDD2.n189 VDD2.n108 171.744
R1815 VDD2.n189 VDD2.n188 171.744
R1816 VDD2.n188 VDD2.n112 171.744
R1817 VDD2.n181 VDD2.n112 171.744
R1818 VDD2.n181 VDD2.n180 171.744
R1819 VDD2.n180 VDD2.n116 171.744
R1820 VDD2.n173 VDD2.n116 171.744
R1821 VDD2.n173 VDD2.n172 171.744
R1822 VDD2.n172 VDD2.n120 171.744
R1823 VDD2.n165 VDD2.n120 171.744
R1824 VDD2.n165 VDD2.n164 171.744
R1825 VDD2.n164 VDD2.n124 171.744
R1826 VDD2.n129 VDD2.n124 171.744
R1827 VDD2.n157 VDD2.n129 171.744
R1828 VDD2.n157 VDD2.n156 171.744
R1829 VDD2.n156 VDD2.n130 171.744
R1830 VDD2.n149 VDD2.n130 171.744
R1831 VDD2.n149 VDD2.n148 171.744
R1832 VDD2.n148 VDD2.n134 171.744
R1833 VDD2.n141 VDD2.n134 171.744
R1834 VDD2.n141 VDD2.n140 171.744
R1835 VDD2.n36 VDD2.n35 171.744
R1836 VDD2.n36 VDD2.n29 171.744
R1837 VDD2.n43 VDD2.n29 171.744
R1838 VDD2.n44 VDD2.n43 171.744
R1839 VDD2.n44 VDD2.n25 171.744
R1840 VDD2.n52 VDD2.n25 171.744
R1841 VDD2.n53 VDD2.n52 171.744
R1842 VDD2.n54 VDD2.n53 171.744
R1843 VDD2.n54 VDD2.n21 171.744
R1844 VDD2.n61 VDD2.n21 171.744
R1845 VDD2.n62 VDD2.n61 171.744
R1846 VDD2.n62 VDD2.n17 171.744
R1847 VDD2.n69 VDD2.n17 171.744
R1848 VDD2.n70 VDD2.n69 171.744
R1849 VDD2.n70 VDD2.n13 171.744
R1850 VDD2.n77 VDD2.n13 171.744
R1851 VDD2.n78 VDD2.n77 171.744
R1852 VDD2.n78 VDD2.n9 171.744
R1853 VDD2.n85 VDD2.n9 171.744
R1854 VDD2.n86 VDD2.n85 171.744
R1855 VDD2.n86 VDD2.n5 171.744
R1856 VDD2.n93 VDD2.n5 171.744
R1857 VDD2.n94 VDD2.n93 171.744
R1858 VDD2.n94 VDD2.n1 171.744
R1859 VDD2.n101 VDD2.n1 171.744
R1860 VDD2.n206 VDD2.n102 95.769
R1861 VDD2.n140 VDD2.t0 85.8723
R1862 VDD2.n35 VDD2.t1 85.8723
R1863 VDD2.n206 VDD2.n205 50.9975
R1864 VDD2.n127 VDD2.n125 13.1884
R1865 VDD2.n55 VDD2.n22 13.1884
R1866 VDD2.n203 VDD2.n103 12.8005
R1867 VDD2.n163 VDD2.n162 12.8005
R1868 VDD2.n159 VDD2.n158 12.8005
R1869 VDD2.n56 VDD2.n24 12.8005
R1870 VDD2.n60 VDD2.n59 12.8005
R1871 VDD2.n100 VDD2.n0 12.8005
R1872 VDD2.n202 VDD2.n105 12.0247
R1873 VDD2.n166 VDD2.n123 12.0247
R1874 VDD2.n155 VDD2.n128 12.0247
R1875 VDD2.n51 VDD2.n50 12.0247
R1876 VDD2.n63 VDD2.n20 12.0247
R1877 VDD2.n99 VDD2.n2 12.0247
R1878 VDD2.n199 VDD2.n198 11.249
R1879 VDD2.n167 VDD2.n121 11.249
R1880 VDD2.n154 VDD2.n131 11.249
R1881 VDD2.n49 VDD2.n26 11.249
R1882 VDD2.n64 VDD2.n18 11.249
R1883 VDD2.n96 VDD2.n95 11.249
R1884 VDD2.n139 VDD2.n138 10.7239
R1885 VDD2.n34 VDD2.n33 10.7239
R1886 VDD2.n195 VDD2.n107 10.4732
R1887 VDD2.n171 VDD2.n170 10.4732
R1888 VDD2.n151 VDD2.n150 10.4732
R1889 VDD2.n46 VDD2.n45 10.4732
R1890 VDD2.n68 VDD2.n67 10.4732
R1891 VDD2.n92 VDD2.n4 10.4732
R1892 VDD2.n194 VDD2.n109 9.69747
R1893 VDD2.n174 VDD2.n119 9.69747
R1894 VDD2.n147 VDD2.n133 9.69747
R1895 VDD2.n42 VDD2.n28 9.69747
R1896 VDD2.n71 VDD2.n16 9.69747
R1897 VDD2.n91 VDD2.n6 9.69747
R1898 VDD2.n201 VDD2.n103 9.45567
R1899 VDD2.n98 VDD2.n0 9.45567
R1900 VDD2.n202 VDD2.n201 9.3005
R1901 VDD2.n200 VDD2.n199 9.3005
R1902 VDD2.n107 VDD2.n106 9.3005
R1903 VDD2.n194 VDD2.n193 9.3005
R1904 VDD2.n192 VDD2.n191 9.3005
R1905 VDD2.n111 VDD2.n110 9.3005
R1906 VDD2.n186 VDD2.n185 9.3005
R1907 VDD2.n184 VDD2.n183 9.3005
R1908 VDD2.n115 VDD2.n114 9.3005
R1909 VDD2.n178 VDD2.n177 9.3005
R1910 VDD2.n176 VDD2.n175 9.3005
R1911 VDD2.n119 VDD2.n118 9.3005
R1912 VDD2.n170 VDD2.n169 9.3005
R1913 VDD2.n168 VDD2.n167 9.3005
R1914 VDD2.n123 VDD2.n122 9.3005
R1915 VDD2.n162 VDD2.n161 9.3005
R1916 VDD2.n160 VDD2.n159 9.3005
R1917 VDD2.n128 VDD2.n126 9.3005
R1918 VDD2.n154 VDD2.n153 9.3005
R1919 VDD2.n152 VDD2.n151 9.3005
R1920 VDD2.n133 VDD2.n132 9.3005
R1921 VDD2.n146 VDD2.n145 9.3005
R1922 VDD2.n144 VDD2.n143 9.3005
R1923 VDD2.n137 VDD2.n136 9.3005
R1924 VDD2.n81 VDD2.n80 9.3005
R1925 VDD2.n83 VDD2.n82 9.3005
R1926 VDD2.n8 VDD2.n7 9.3005
R1927 VDD2.n89 VDD2.n88 9.3005
R1928 VDD2.n91 VDD2.n90 9.3005
R1929 VDD2.n4 VDD2.n3 9.3005
R1930 VDD2.n97 VDD2.n96 9.3005
R1931 VDD2.n99 VDD2.n98 9.3005
R1932 VDD2.n75 VDD2.n74 9.3005
R1933 VDD2.n73 VDD2.n72 9.3005
R1934 VDD2.n16 VDD2.n15 9.3005
R1935 VDD2.n67 VDD2.n66 9.3005
R1936 VDD2.n65 VDD2.n64 9.3005
R1937 VDD2.n20 VDD2.n19 9.3005
R1938 VDD2.n59 VDD2.n58 9.3005
R1939 VDD2.n32 VDD2.n31 9.3005
R1940 VDD2.n39 VDD2.n38 9.3005
R1941 VDD2.n41 VDD2.n40 9.3005
R1942 VDD2.n28 VDD2.n27 9.3005
R1943 VDD2.n47 VDD2.n46 9.3005
R1944 VDD2.n49 VDD2.n48 9.3005
R1945 VDD2.n50 VDD2.n23 9.3005
R1946 VDD2.n57 VDD2.n56 9.3005
R1947 VDD2.n12 VDD2.n11 9.3005
R1948 VDD2.n191 VDD2.n190 8.92171
R1949 VDD2.n175 VDD2.n117 8.92171
R1950 VDD2.n146 VDD2.n135 8.92171
R1951 VDD2.n41 VDD2.n30 8.92171
R1952 VDD2.n72 VDD2.n14 8.92171
R1953 VDD2.n88 VDD2.n87 8.92171
R1954 VDD2.n187 VDD2.n111 8.14595
R1955 VDD2.n179 VDD2.n178 8.14595
R1956 VDD2.n143 VDD2.n142 8.14595
R1957 VDD2.n38 VDD2.n37 8.14595
R1958 VDD2.n76 VDD2.n75 8.14595
R1959 VDD2.n84 VDD2.n8 8.14595
R1960 VDD2.n186 VDD2.n113 7.3702
R1961 VDD2.n182 VDD2.n115 7.3702
R1962 VDD2.n139 VDD2.n137 7.3702
R1963 VDD2.n34 VDD2.n32 7.3702
R1964 VDD2.n79 VDD2.n12 7.3702
R1965 VDD2.n83 VDD2.n10 7.3702
R1966 VDD2.n183 VDD2.n113 6.59444
R1967 VDD2.n183 VDD2.n182 6.59444
R1968 VDD2.n80 VDD2.n79 6.59444
R1969 VDD2.n80 VDD2.n10 6.59444
R1970 VDD2.n187 VDD2.n186 5.81868
R1971 VDD2.n179 VDD2.n115 5.81868
R1972 VDD2.n142 VDD2.n137 5.81868
R1973 VDD2.n37 VDD2.n32 5.81868
R1974 VDD2.n76 VDD2.n12 5.81868
R1975 VDD2.n84 VDD2.n83 5.81868
R1976 VDD2.n190 VDD2.n111 5.04292
R1977 VDD2.n178 VDD2.n117 5.04292
R1978 VDD2.n143 VDD2.n135 5.04292
R1979 VDD2.n38 VDD2.n30 5.04292
R1980 VDD2.n75 VDD2.n14 5.04292
R1981 VDD2.n87 VDD2.n8 5.04292
R1982 VDD2.n191 VDD2.n109 4.26717
R1983 VDD2.n175 VDD2.n174 4.26717
R1984 VDD2.n147 VDD2.n146 4.26717
R1985 VDD2.n42 VDD2.n41 4.26717
R1986 VDD2.n72 VDD2.n71 4.26717
R1987 VDD2.n88 VDD2.n6 4.26717
R1988 VDD2.n195 VDD2.n194 3.49141
R1989 VDD2.n171 VDD2.n119 3.49141
R1990 VDD2.n150 VDD2.n133 3.49141
R1991 VDD2.n45 VDD2.n28 3.49141
R1992 VDD2.n68 VDD2.n16 3.49141
R1993 VDD2.n92 VDD2.n91 3.49141
R1994 VDD2.n198 VDD2.n107 2.71565
R1995 VDD2.n170 VDD2.n121 2.71565
R1996 VDD2.n151 VDD2.n131 2.71565
R1997 VDD2.n46 VDD2.n26 2.71565
R1998 VDD2.n67 VDD2.n18 2.71565
R1999 VDD2.n95 VDD2.n4 2.71565
R2000 VDD2.n138 VDD2.n136 2.41282
R2001 VDD2.n33 VDD2.n31 2.41282
R2002 VDD2.n199 VDD2.n105 1.93989
R2003 VDD2.n167 VDD2.n166 1.93989
R2004 VDD2.n155 VDD2.n154 1.93989
R2005 VDD2.n51 VDD2.n49 1.93989
R2006 VDD2.n64 VDD2.n63 1.93989
R2007 VDD2.n96 VDD2.n2 1.93989
R2008 VDD2.n203 VDD2.n202 1.16414
R2009 VDD2.n163 VDD2.n123 1.16414
R2010 VDD2.n158 VDD2.n128 1.16414
R2011 VDD2.n50 VDD2.n24 1.16414
R2012 VDD2.n60 VDD2.n20 1.16414
R2013 VDD2.n100 VDD2.n99 1.16414
R2014 VDD2 VDD2.n206 0.679379
R2015 VDD2.n205 VDD2.n103 0.388379
R2016 VDD2.n162 VDD2.n125 0.388379
R2017 VDD2.n159 VDD2.n127 0.388379
R2018 VDD2.n56 VDD2.n55 0.388379
R2019 VDD2.n59 VDD2.n22 0.388379
R2020 VDD2.n102 VDD2.n0 0.388379
R2021 VDD2.n201 VDD2.n200 0.155672
R2022 VDD2.n200 VDD2.n106 0.155672
R2023 VDD2.n193 VDD2.n106 0.155672
R2024 VDD2.n193 VDD2.n192 0.155672
R2025 VDD2.n192 VDD2.n110 0.155672
R2026 VDD2.n185 VDD2.n110 0.155672
R2027 VDD2.n185 VDD2.n184 0.155672
R2028 VDD2.n184 VDD2.n114 0.155672
R2029 VDD2.n177 VDD2.n114 0.155672
R2030 VDD2.n177 VDD2.n176 0.155672
R2031 VDD2.n176 VDD2.n118 0.155672
R2032 VDD2.n169 VDD2.n118 0.155672
R2033 VDD2.n169 VDD2.n168 0.155672
R2034 VDD2.n168 VDD2.n122 0.155672
R2035 VDD2.n161 VDD2.n122 0.155672
R2036 VDD2.n161 VDD2.n160 0.155672
R2037 VDD2.n160 VDD2.n126 0.155672
R2038 VDD2.n153 VDD2.n126 0.155672
R2039 VDD2.n153 VDD2.n152 0.155672
R2040 VDD2.n152 VDD2.n132 0.155672
R2041 VDD2.n145 VDD2.n132 0.155672
R2042 VDD2.n145 VDD2.n144 0.155672
R2043 VDD2.n144 VDD2.n136 0.155672
R2044 VDD2.n39 VDD2.n31 0.155672
R2045 VDD2.n40 VDD2.n39 0.155672
R2046 VDD2.n40 VDD2.n27 0.155672
R2047 VDD2.n47 VDD2.n27 0.155672
R2048 VDD2.n48 VDD2.n47 0.155672
R2049 VDD2.n48 VDD2.n23 0.155672
R2050 VDD2.n57 VDD2.n23 0.155672
R2051 VDD2.n58 VDD2.n57 0.155672
R2052 VDD2.n58 VDD2.n19 0.155672
R2053 VDD2.n65 VDD2.n19 0.155672
R2054 VDD2.n66 VDD2.n65 0.155672
R2055 VDD2.n66 VDD2.n15 0.155672
R2056 VDD2.n73 VDD2.n15 0.155672
R2057 VDD2.n74 VDD2.n73 0.155672
R2058 VDD2.n74 VDD2.n11 0.155672
R2059 VDD2.n81 VDD2.n11 0.155672
R2060 VDD2.n82 VDD2.n81 0.155672
R2061 VDD2.n82 VDD2.n7 0.155672
R2062 VDD2.n89 VDD2.n7 0.155672
R2063 VDD2.n90 VDD2.n89 0.155672
R2064 VDD2.n90 VDD2.n3 0.155672
R2065 VDD2.n97 VDD2.n3 0.155672
R2066 VDD2.n98 VDD2.n97 0.155672
R2067 VP.n0 VP.t0 275.81
R2068 VP.n0 VP.t1 226.188
R2069 VP VP.n0 0.336784
R2070 VDD1.n102 VDD1.n101 756.745
R2071 VDD1.n205 VDD1.n204 756.745
R2072 VDD1.n101 VDD1.n100 585
R2073 VDD1.n2 VDD1.n1 585
R2074 VDD1.n95 VDD1.n94 585
R2075 VDD1.n93 VDD1.n92 585
R2076 VDD1.n6 VDD1.n5 585
R2077 VDD1.n87 VDD1.n86 585
R2078 VDD1.n85 VDD1.n84 585
R2079 VDD1.n10 VDD1.n9 585
R2080 VDD1.n79 VDD1.n78 585
R2081 VDD1.n77 VDD1.n76 585
R2082 VDD1.n14 VDD1.n13 585
R2083 VDD1.n71 VDD1.n70 585
R2084 VDD1.n69 VDD1.n68 585
R2085 VDD1.n18 VDD1.n17 585
R2086 VDD1.n63 VDD1.n62 585
R2087 VDD1.n61 VDD1.n60 585
R2088 VDD1.n22 VDD1.n21 585
R2089 VDD1.n26 VDD1.n24 585
R2090 VDD1.n55 VDD1.n54 585
R2091 VDD1.n53 VDD1.n52 585
R2092 VDD1.n28 VDD1.n27 585
R2093 VDD1.n47 VDD1.n46 585
R2094 VDD1.n45 VDD1.n44 585
R2095 VDD1.n32 VDD1.n31 585
R2096 VDD1.n39 VDD1.n38 585
R2097 VDD1.n37 VDD1.n36 585
R2098 VDD1.n138 VDD1.n137 585
R2099 VDD1.n140 VDD1.n139 585
R2100 VDD1.n133 VDD1.n132 585
R2101 VDD1.n146 VDD1.n145 585
R2102 VDD1.n148 VDD1.n147 585
R2103 VDD1.n129 VDD1.n128 585
R2104 VDD1.n155 VDD1.n154 585
R2105 VDD1.n156 VDD1.n127 585
R2106 VDD1.n158 VDD1.n157 585
R2107 VDD1.n125 VDD1.n124 585
R2108 VDD1.n164 VDD1.n163 585
R2109 VDD1.n166 VDD1.n165 585
R2110 VDD1.n121 VDD1.n120 585
R2111 VDD1.n172 VDD1.n171 585
R2112 VDD1.n174 VDD1.n173 585
R2113 VDD1.n117 VDD1.n116 585
R2114 VDD1.n180 VDD1.n179 585
R2115 VDD1.n182 VDD1.n181 585
R2116 VDD1.n113 VDD1.n112 585
R2117 VDD1.n188 VDD1.n187 585
R2118 VDD1.n190 VDD1.n189 585
R2119 VDD1.n109 VDD1.n108 585
R2120 VDD1.n196 VDD1.n195 585
R2121 VDD1.n198 VDD1.n197 585
R2122 VDD1.n105 VDD1.n104 585
R2123 VDD1.n204 VDD1.n203 585
R2124 VDD1.n35 VDD1.t1 329.036
R2125 VDD1.n136 VDD1.t0 329.036
R2126 VDD1.n101 VDD1.n1 171.744
R2127 VDD1.n94 VDD1.n1 171.744
R2128 VDD1.n94 VDD1.n93 171.744
R2129 VDD1.n93 VDD1.n5 171.744
R2130 VDD1.n86 VDD1.n5 171.744
R2131 VDD1.n86 VDD1.n85 171.744
R2132 VDD1.n85 VDD1.n9 171.744
R2133 VDD1.n78 VDD1.n9 171.744
R2134 VDD1.n78 VDD1.n77 171.744
R2135 VDD1.n77 VDD1.n13 171.744
R2136 VDD1.n70 VDD1.n13 171.744
R2137 VDD1.n70 VDD1.n69 171.744
R2138 VDD1.n69 VDD1.n17 171.744
R2139 VDD1.n62 VDD1.n17 171.744
R2140 VDD1.n62 VDD1.n61 171.744
R2141 VDD1.n61 VDD1.n21 171.744
R2142 VDD1.n26 VDD1.n21 171.744
R2143 VDD1.n54 VDD1.n26 171.744
R2144 VDD1.n54 VDD1.n53 171.744
R2145 VDD1.n53 VDD1.n27 171.744
R2146 VDD1.n46 VDD1.n27 171.744
R2147 VDD1.n46 VDD1.n45 171.744
R2148 VDD1.n45 VDD1.n31 171.744
R2149 VDD1.n38 VDD1.n31 171.744
R2150 VDD1.n38 VDD1.n37 171.744
R2151 VDD1.n139 VDD1.n138 171.744
R2152 VDD1.n139 VDD1.n132 171.744
R2153 VDD1.n146 VDD1.n132 171.744
R2154 VDD1.n147 VDD1.n146 171.744
R2155 VDD1.n147 VDD1.n128 171.744
R2156 VDD1.n155 VDD1.n128 171.744
R2157 VDD1.n156 VDD1.n155 171.744
R2158 VDD1.n157 VDD1.n156 171.744
R2159 VDD1.n157 VDD1.n124 171.744
R2160 VDD1.n164 VDD1.n124 171.744
R2161 VDD1.n165 VDD1.n164 171.744
R2162 VDD1.n165 VDD1.n120 171.744
R2163 VDD1.n172 VDD1.n120 171.744
R2164 VDD1.n173 VDD1.n172 171.744
R2165 VDD1.n173 VDD1.n116 171.744
R2166 VDD1.n180 VDD1.n116 171.744
R2167 VDD1.n181 VDD1.n180 171.744
R2168 VDD1.n181 VDD1.n112 171.744
R2169 VDD1.n188 VDD1.n112 171.744
R2170 VDD1.n189 VDD1.n188 171.744
R2171 VDD1.n189 VDD1.n108 171.744
R2172 VDD1.n196 VDD1.n108 171.744
R2173 VDD1.n197 VDD1.n196 171.744
R2174 VDD1.n197 VDD1.n104 171.744
R2175 VDD1.n204 VDD1.n104 171.744
R2176 VDD1 VDD1.n205 96.9145
R2177 VDD1.n37 VDD1.t1 85.8723
R2178 VDD1.n138 VDD1.t0 85.8723
R2179 VDD1 VDD1.n102 51.6763
R2180 VDD1.n24 VDD1.n22 13.1884
R2181 VDD1.n158 VDD1.n125 13.1884
R2182 VDD1.n100 VDD1.n0 12.8005
R2183 VDD1.n60 VDD1.n59 12.8005
R2184 VDD1.n56 VDD1.n55 12.8005
R2185 VDD1.n159 VDD1.n127 12.8005
R2186 VDD1.n163 VDD1.n162 12.8005
R2187 VDD1.n203 VDD1.n103 12.8005
R2188 VDD1.n99 VDD1.n2 12.0247
R2189 VDD1.n63 VDD1.n20 12.0247
R2190 VDD1.n52 VDD1.n25 12.0247
R2191 VDD1.n154 VDD1.n153 12.0247
R2192 VDD1.n166 VDD1.n123 12.0247
R2193 VDD1.n202 VDD1.n105 12.0247
R2194 VDD1.n96 VDD1.n95 11.249
R2195 VDD1.n64 VDD1.n18 11.249
R2196 VDD1.n51 VDD1.n28 11.249
R2197 VDD1.n152 VDD1.n129 11.249
R2198 VDD1.n167 VDD1.n121 11.249
R2199 VDD1.n199 VDD1.n198 11.249
R2200 VDD1.n36 VDD1.n35 10.7239
R2201 VDD1.n137 VDD1.n136 10.7239
R2202 VDD1.n92 VDD1.n4 10.4732
R2203 VDD1.n68 VDD1.n67 10.4732
R2204 VDD1.n48 VDD1.n47 10.4732
R2205 VDD1.n149 VDD1.n148 10.4732
R2206 VDD1.n171 VDD1.n170 10.4732
R2207 VDD1.n195 VDD1.n107 10.4732
R2208 VDD1.n91 VDD1.n6 9.69747
R2209 VDD1.n71 VDD1.n16 9.69747
R2210 VDD1.n44 VDD1.n30 9.69747
R2211 VDD1.n145 VDD1.n131 9.69747
R2212 VDD1.n174 VDD1.n119 9.69747
R2213 VDD1.n194 VDD1.n109 9.69747
R2214 VDD1.n98 VDD1.n0 9.45567
R2215 VDD1.n201 VDD1.n103 9.45567
R2216 VDD1.n99 VDD1.n98 9.3005
R2217 VDD1.n97 VDD1.n96 9.3005
R2218 VDD1.n4 VDD1.n3 9.3005
R2219 VDD1.n91 VDD1.n90 9.3005
R2220 VDD1.n89 VDD1.n88 9.3005
R2221 VDD1.n8 VDD1.n7 9.3005
R2222 VDD1.n83 VDD1.n82 9.3005
R2223 VDD1.n81 VDD1.n80 9.3005
R2224 VDD1.n12 VDD1.n11 9.3005
R2225 VDD1.n75 VDD1.n74 9.3005
R2226 VDD1.n73 VDD1.n72 9.3005
R2227 VDD1.n16 VDD1.n15 9.3005
R2228 VDD1.n67 VDD1.n66 9.3005
R2229 VDD1.n65 VDD1.n64 9.3005
R2230 VDD1.n20 VDD1.n19 9.3005
R2231 VDD1.n59 VDD1.n58 9.3005
R2232 VDD1.n57 VDD1.n56 9.3005
R2233 VDD1.n25 VDD1.n23 9.3005
R2234 VDD1.n51 VDD1.n50 9.3005
R2235 VDD1.n49 VDD1.n48 9.3005
R2236 VDD1.n30 VDD1.n29 9.3005
R2237 VDD1.n43 VDD1.n42 9.3005
R2238 VDD1.n41 VDD1.n40 9.3005
R2239 VDD1.n34 VDD1.n33 9.3005
R2240 VDD1.n184 VDD1.n183 9.3005
R2241 VDD1.n186 VDD1.n185 9.3005
R2242 VDD1.n111 VDD1.n110 9.3005
R2243 VDD1.n192 VDD1.n191 9.3005
R2244 VDD1.n194 VDD1.n193 9.3005
R2245 VDD1.n107 VDD1.n106 9.3005
R2246 VDD1.n200 VDD1.n199 9.3005
R2247 VDD1.n202 VDD1.n201 9.3005
R2248 VDD1.n178 VDD1.n177 9.3005
R2249 VDD1.n176 VDD1.n175 9.3005
R2250 VDD1.n119 VDD1.n118 9.3005
R2251 VDD1.n170 VDD1.n169 9.3005
R2252 VDD1.n168 VDD1.n167 9.3005
R2253 VDD1.n123 VDD1.n122 9.3005
R2254 VDD1.n162 VDD1.n161 9.3005
R2255 VDD1.n135 VDD1.n134 9.3005
R2256 VDD1.n142 VDD1.n141 9.3005
R2257 VDD1.n144 VDD1.n143 9.3005
R2258 VDD1.n131 VDD1.n130 9.3005
R2259 VDD1.n150 VDD1.n149 9.3005
R2260 VDD1.n152 VDD1.n151 9.3005
R2261 VDD1.n153 VDD1.n126 9.3005
R2262 VDD1.n160 VDD1.n159 9.3005
R2263 VDD1.n115 VDD1.n114 9.3005
R2264 VDD1.n88 VDD1.n87 8.92171
R2265 VDD1.n72 VDD1.n14 8.92171
R2266 VDD1.n43 VDD1.n32 8.92171
R2267 VDD1.n144 VDD1.n133 8.92171
R2268 VDD1.n175 VDD1.n117 8.92171
R2269 VDD1.n191 VDD1.n190 8.92171
R2270 VDD1.n84 VDD1.n8 8.14595
R2271 VDD1.n76 VDD1.n75 8.14595
R2272 VDD1.n40 VDD1.n39 8.14595
R2273 VDD1.n141 VDD1.n140 8.14595
R2274 VDD1.n179 VDD1.n178 8.14595
R2275 VDD1.n187 VDD1.n111 8.14595
R2276 VDD1.n83 VDD1.n10 7.3702
R2277 VDD1.n79 VDD1.n12 7.3702
R2278 VDD1.n36 VDD1.n34 7.3702
R2279 VDD1.n137 VDD1.n135 7.3702
R2280 VDD1.n182 VDD1.n115 7.3702
R2281 VDD1.n186 VDD1.n113 7.3702
R2282 VDD1.n80 VDD1.n10 6.59444
R2283 VDD1.n80 VDD1.n79 6.59444
R2284 VDD1.n183 VDD1.n182 6.59444
R2285 VDD1.n183 VDD1.n113 6.59444
R2286 VDD1.n84 VDD1.n83 5.81868
R2287 VDD1.n76 VDD1.n12 5.81868
R2288 VDD1.n39 VDD1.n34 5.81868
R2289 VDD1.n140 VDD1.n135 5.81868
R2290 VDD1.n179 VDD1.n115 5.81868
R2291 VDD1.n187 VDD1.n186 5.81868
R2292 VDD1.n87 VDD1.n8 5.04292
R2293 VDD1.n75 VDD1.n14 5.04292
R2294 VDD1.n40 VDD1.n32 5.04292
R2295 VDD1.n141 VDD1.n133 5.04292
R2296 VDD1.n178 VDD1.n117 5.04292
R2297 VDD1.n190 VDD1.n111 5.04292
R2298 VDD1.n88 VDD1.n6 4.26717
R2299 VDD1.n72 VDD1.n71 4.26717
R2300 VDD1.n44 VDD1.n43 4.26717
R2301 VDD1.n145 VDD1.n144 4.26717
R2302 VDD1.n175 VDD1.n174 4.26717
R2303 VDD1.n191 VDD1.n109 4.26717
R2304 VDD1.n92 VDD1.n91 3.49141
R2305 VDD1.n68 VDD1.n16 3.49141
R2306 VDD1.n47 VDD1.n30 3.49141
R2307 VDD1.n148 VDD1.n131 3.49141
R2308 VDD1.n171 VDD1.n119 3.49141
R2309 VDD1.n195 VDD1.n194 3.49141
R2310 VDD1.n95 VDD1.n4 2.71565
R2311 VDD1.n67 VDD1.n18 2.71565
R2312 VDD1.n48 VDD1.n28 2.71565
R2313 VDD1.n149 VDD1.n129 2.71565
R2314 VDD1.n170 VDD1.n121 2.71565
R2315 VDD1.n198 VDD1.n107 2.71565
R2316 VDD1.n35 VDD1.n33 2.41282
R2317 VDD1.n136 VDD1.n134 2.41282
R2318 VDD1.n96 VDD1.n2 1.93989
R2319 VDD1.n64 VDD1.n63 1.93989
R2320 VDD1.n52 VDD1.n51 1.93989
R2321 VDD1.n154 VDD1.n152 1.93989
R2322 VDD1.n167 VDD1.n166 1.93989
R2323 VDD1.n199 VDD1.n105 1.93989
R2324 VDD1.n100 VDD1.n99 1.16414
R2325 VDD1.n60 VDD1.n20 1.16414
R2326 VDD1.n55 VDD1.n25 1.16414
R2327 VDD1.n153 VDD1.n127 1.16414
R2328 VDD1.n163 VDD1.n123 1.16414
R2329 VDD1.n203 VDD1.n202 1.16414
R2330 VDD1.n102 VDD1.n0 0.388379
R2331 VDD1.n59 VDD1.n22 0.388379
R2332 VDD1.n56 VDD1.n24 0.388379
R2333 VDD1.n159 VDD1.n158 0.388379
R2334 VDD1.n162 VDD1.n125 0.388379
R2335 VDD1.n205 VDD1.n103 0.388379
R2336 VDD1.n98 VDD1.n97 0.155672
R2337 VDD1.n97 VDD1.n3 0.155672
R2338 VDD1.n90 VDD1.n3 0.155672
R2339 VDD1.n90 VDD1.n89 0.155672
R2340 VDD1.n89 VDD1.n7 0.155672
R2341 VDD1.n82 VDD1.n7 0.155672
R2342 VDD1.n82 VDD1.n81 0.155672
R2343 VDD1.n81 VDD1.n11 0.155672
R2344 VDD1.n74 VDD1.n11 0.155672
R2345 VDD1.n74 VDD1.n73 0.155672
R2346 VDD1.n73 VDD1.n15 0.155672
R2347 VDD1.n66 VDD1.n15 0.155672
R2348 VDD1.n66 VDD1.n65 0.155672
R2349 VDD1.n65 VDD1.n19 0.155672
R2350 VDD1.n58 VDD1.n19 0.155672
R2351 VDD1.n58 VDD1.n57 0.155672
R2352 VDD1.n57 VDD1.n23 0.155672
R2353 VDD1.n50 VDD1.n23 0.155672
R2354 VDD1.n50 VDD1.n49 0.155672
R2355 VDD1.n49 VDD1.n29 0.155672
R2356 VDD1.n42 VDD1.n29 0.155672
R2357 VDD1.n42 VDD1.n41 0.155672
R2358 VDD1.n41 VDD1.n33 0.155672
R2359 VDD1.n142 VDD1.n134 0.155672
R2360 VDD1.n143 VDD1.n142 0.155672
R2361 VDD1.n143 VDD1.n130 0.155672
R2362 VDD1.n150 VDD1.n130 0.155672
R2363 VDD1.n151 VDD1.n150 0.155672
R2364 VDD1.n151 VDD1.n126 0.155672
R2365 VDD1.n160 VDD1.n126 0.155672
R2366 VDD1.n161 VDD1.n160 0.155672
R2367 VDD1.n161 VDD1.n122 0.155672
R2368 VDD1.n168 VDD1.n122 0.155672
R2369 VDD1.n169 VDD1.n168 0.155672
R2370 VDD1.n169 VDD1.n118 0.155672
R2371 VDD1.n176 VDD1.n118 0.155672
R2372 VDD1.n177 VDD1.n176 0.155672
R2373 VDD1.n177 VDD1.n114 0.155672
R2374 VDD1.n184 VDD1.n114 0.155672
R2375 VDD1.n185 VDD1.n184 0.155672
R2376 VDD1.n185 VDD1.n110 0.155672
R2377 VDD1.n192 VDD1.n110 0.155672
R2378 VDD1.n193 VDD1.n192 0.155672
R2379 VDD1.n193 VDD1.n106 0.155672
R2380 VDD1.n200 VDD1.n106 0.155672
R2381 VDD1.n201 VDD1.n200 0.155672
C0 VTAIL B 5.13989f
C1 B VP 1.56451f
C2 VTAIL VP 3.55934f
C3 VN B 1.1205f
C4 VN VTAIL 3.54494f
C5 VDD1 VDD2 0.66939f
C6 VN VP 6.67583f
C7 w_n2122_n4714# VDD1 2.2433f
C8 w_n2122_n4714# VDD2 2.26856f
C9 VDD1 B 2.2298f
C10 VDD1 VTAIL 6.84419f
C11 VDD1 VP 4.36676f
C12 VDD2 B 2.25943f
C13 VDD2 VTAIL 6.89282f
C14 VDD1 VN 0.148099f
C15 VDD2 VP 0.331513f
C16 VDD2 VN 4.1871f
C17 w_n2122_n4714# B 10.6419f
C18 w_n2122_n4714# VTAIL 3.70365f
C19 w_n2122_n4714# VP 3.31952f
C20 w_n2122_n4714# VN 3.04933f
C21 VDD2 VSUBS 1.144512f
C22 VDD1 VSUBS 5.61533f
C23 VTAIL VSUBS 1.262126f
C24 VN VSUBS 9.178479f
C25 VP VSUBS 1.912326f
C26 B VSUBS 4.44262f
C27 w_n2122_n4714# VSUBS 0.122253p
C28 VDD1.n0 VSUBS 0.015647f
C29 VDD1.n1 VSUBS 0.03535f
C30 VDD1.n2 VSUBS 0.015835f
C31 VDD1.n3 VSUBS 0.027832f
C32 VDD1.n4 VSUBS 0.014956f
C33 VDD1.n5 VSUBS 0.03535f
C34 VDD1.n6 VSUBS 0.015835f
C35 VDD1.n7 VSUBS 0.027832f
C36 VDD1.n8 VSUBS 0.014956f
C37 VDD1.n9 VSUBS 0.03535f
C38 VDD1.n10 VSUBS 0.015835f
C39 VDD1.n11 VSUBS 0.027832f
C40 VDD1.n12 VSUBS 0.014956f
C41 VDD1.n13 VSUBS 0.03535f
C42 VDD1.n14 VSUBS 0.015835f
C43 VDD1.n15 VSUBS 0.027832f
C44 VDD1.n16 VSUBS 0.014956f
C45 VDD1.n17 VSUBS 0.03535f
C46 VDD1.n18 VSUBS 0.015835f
C47 VDD1.n19 VSUBS 0.027832f
C48 VDD1.n20 VSUBS 0.014956f
C49 VDD1.n21 VSUBS 0.03535f
C50 VDD1.n22 VSUBS 0.015396f
C51 VDD1.n23 VSUBS 0.027832f
C52 VDD1.n24 VSUBS 0.015396f
C53 VDD1.n25 VSUBS 0.014956f
C54 VDD1.n26 VSUBS 0.03535f
C55 VDD1.n27 VSUBS 0.03535f
C56 VDD1.n28 VSUBS 0.015835f
C57 VDD1.n29 VSUBS 0.027832f
C58 VDD1.n30 VSUBS 0.014956f
C59 VDD1.n31 VSUBS 0.03535f
C60 VDD1.n32 VSUBS 0.015835f
C61 VDD1.n33 VSUBS 2.18819f
C62 VDD1.n34 VSUBS 0.014956f
C63 VDD1.t1 VSUBS 0.076807f
C64 VDD1.n35 VSUBS 0.303885f
C65 VDD1.n36 VSUBS 0.026592f
C66 VDD1.n37 VSUBS 0.026512f
C67 VDD1.n38 VSUBS 0.03535f
C68 VDD1.n39 VSUBS 0.015835f
C69 VDD1.n40 VSUBS 0.014956f
C70 VDD1.n41 VSUBS 0.027832f
C71 VDD1.n42 VSUBS 0.027832f
C72 VDD1.n43 VSUBS 0.014956f
C73 VDD1.n44 VSUBS 0.015835f
C74 VDD1.n45 VSUBS 0.03535f
C75 VDD1.n46 VSUBS 0.03535f
C76 VDD1.n47 VSUBS 0.015835f
C77 VDD1.n48 VSUBS 0.014956f
C78 VDD1.n49 VSUBS 0.027832f
C79 VDD1.n50 VSUBS 0.027832f
C80 VDD1.n51 VSUBS 0.014956f
C81 VDD1.n52 VSUBS 0.015835f
C82 VDD1.n53 VSUBS 0.03535f
C83 VDD1.n54 VSUBS 0.03535f
C84 VDD1.n55 VSUBS 0.015835f
C85 VDD1.n56 VSUBS 0.014956f
C86 VDD1.n57 VSUBS 0.027832f
C87 VDD1.n58 VSUBS 0.027832f
C88 VDD1.n59 VSUBS 0.014956f
C89 VDD1.n60 VSUBS 0.015835f
C90 VDD1.n61 VSUBS 0.03535f
C91 VDD1.n62 VSUBS 0.03535f
C92 VDD1.n63 VSUBS 0.015835f
C93 VDD1.n64 VSUBS 0.014956f
C94 VDD1.n65 VSUBS 0.027832f
C95 VDD1.n66 VSUBS 0.027832f
C96 VDD1.n67 VSUBS 0.014956f
C97 VDD1.n68 VSUBS 0.015835f
C98 VDD1.n69 VSUBS 0.03535f
C99 VDD1.n70 VSUBS 0.03535f
C100 VDD1.n71 VSUBS 0.015835f
C101 VDD1.n72 VSUBS 0.014956f
C102 VDD1.n73 VSUBS 0.027832f
C103 VDD1.n74 VSUBS 0.027832f
C104 VDD1.n75 VSUBS 0.014956f
C105 VDD1.n76 VSUBS 0.015835f
C106 VDD1.n77 VSUBS 0.03535f
C107 VDD1.n78 VSUBS 0.03535f
C108 VDD1.n79 VSUBS 0.015835f
C109 VDD1.n80 VSUBS 0.014956f
C110 VDD1.n81 VSUBS 0.027832f
C111 VDD1.n82 VSUBS 0.027832f
C112 VDD1.n83 VSUBS 0.014956f
C113 VDD1.n84 VSUBS 0.015835f
C114 VDD1.n85 VSUBS 0.03535f
C115 VDD1.n86 VSUBS 0.03535f
C116 VDD1.n87 VSUBS 0.015835f
C117 VDD1.n88 VSUBS 0.014956f
C118 VDD1.n89 VSUBS 0.027832f
C119 VDD1.n90 VSUBS 0.027832f
C120 VDD1.n91 VSUBS 0.014956f
C121 VDD1.n92 VSUBS 0.015835f
C122 VDD1.n93 VSUBS 0.03535f
C123 VDD1.n94 VSUBS 0.03535f
C124 VDD1.n95 VSUBS 0.015835f
C125 VDD1.n96 VSUBS 0.014956f
C126 VDD1.n97 VSUBS 0.027832f
C127 VDD1.n98 VSUBS 0.069275f
C128 VDD1.n99 VSUBS 0.014956f
C129 VDD1.n100 VSUBS 0.015835f
C130 VDD1.n101 VSUBS 0.077546f
C131 VDD1.n102 VSUBS 0.071636f
C132 VDD1.n103 VSUBS 0.015647f
C133 VDD1.n104 VSUBS 0.03535f
C134 VDD1.n105 VSUBS 0.015835f
C135 VDD1.n106 VSUBS 0.027832f
C136 VDD1.n107 VSUBS 0.014956f
C137 VDD1.n108 VSUBS 0.03535f
C138 VDD1.n109 VSUBS 0.015835f
C139 VDD1.n110 VSUBS 0.027832f
C140 VDD1.n111 VSUBS 0.014956f
C141 VDD1.n112 VSUBS 0.03535f
C142 VDD1.n113 VSUBS 0.015835f
C143 VDD1.n114 VSUBS 0.027832f
C144 VDD1.n115 VSUBS 0.014956f
C145 VDD1.n116 VSUBS 0.03535f
C146 VDD1.n117 VSUBS 0.015835f
C147 VDD1.n118 VSUBS 0.027832f
C148 VDD1.n119 VSUBS 0.014956f
C149 VDD1.n120 VSUBS 0.03535f
C150 VDD1.n121 VSUBS 0.015835f
C151 VDD1.n122 VSUBS 0.027832f
C152 VDD1.n123 VSUBS 0.014956f
C153 VDD1.n124 VSUBS 0.03535f
C154 VDD1.n125 VSUBS 0.015396f
C155 VDD1.n126 VSUBS 0.027832f
C156 VDD1.n127 VSUBS 0.015835f
C157 VDD1.n128 VSUBS 0.03535f
C158 VDD1.n129 VSUBS 0.015835f
C159 VDD1.n130 VSUBS 0.027832f
C160 VDD1.n131 VSUBS 0.014956f
C161 VDD1.n132 VSUBS 0.03535f
C162 VDD1.n133 VSUBS 0.015835f
C163 VDD1.n134 VSUBS 2.18819f
C164 VDD1.n135 VSUBS 0.014956f
C165 VDD1.t0 VSUBS 0.076807f
C166 VDD1.n136 VSUBS 0.303885f
C167 VDD1.n137 VSUBS 0.026592f
C168 VDD1.n138 VSUBS 0.026512f
C169 VDD1.n139 VSUBS 0.03535f
C170 VDD1.n140 VSUBS 0.015835f
C171 VDD1.n141 VSUBS 0.014956f
C172 VDD1.n142 VSUBS 0.027832f
C173 VDD1.n143 VSUBS 0.027832f
C174 VDD1.n144 VSUBS 0.014956f
C175 VDD1.n145 VSUBS 0.015835f
C176 VDD1.n146 VSUBS 0.03535f
C177 VDD1.n147 VSUBS 0.03535f
C178 VDD1.n148 VSUBS 0.015835f
C179 VDD1.n149 VSUBS 0.014956f
C180 VDD1.n150 VSUBS 0.027832f
C181 VDD1.n151 VSUBS 0.027832f
C182 VDD1.n152 VSUBS 0.014956f
C183 VDD1.n153 VSUBS 0.014956f
C184 VDD1.n154 VSUBS 0.015835f
C185 VDD1.n155 VSUBS 0.03535f
C186 VDD1.n156 VSUBS 0.03535f
C187 VDD1.n157 VSUBS 0.03535f
C188 VDD1.n158 VSUBS 0.015396f
C189 VDD1.n159 VSUBS 0.014956f
C190 VDD1.n160 VSUBS 0.027832f
C191 VDD1.n161 VSUBS 0.027832f
C192 VDD1.n162 VSUBS 0.014956f
C193 VDD1.n163 VSUBS 0.015835f
C194 VDD1.n164 VSUBS 0.03535f
C195 VDD1.n165 VSUBS 0.03535f
C196 VDD1.n166 VSUBS 0.015835f
C197 VDD1.n167 VSUBS 0.014956f
C198 VDD1.n168 VSUBS 0.027832f
C199 VDD1.n169 VSUBS 0.027832f
C200 VDD1.n170 VSUBS 0.014956f
C201 VDD1.n171 VSUBS 0.015835f
C202 VDD1.n172 VSUBS 0.03535f
C203 VDD1.n173 VSUBS 0.03535f
C204 VDD1.n174 VSUBS 0.015835f
C205 VDD1.n175 VSUBS 0.014956f
C206 VDD1.n176 VSUBS 0.027832f
C207 VDD1.n177 VSUBS 0.027832f
C208 VDD1.n178 VSUBS 0.014956f
C209 VDD1.n179 VSUBS 0.015835f
C210 VDD1.n180 VSUBS 0.03535f
C211 VDD1.n181 VSUBS 0.03535f
C212 VDD1.n182 VSUBS 0.015835f
C213 VDD1.n183 VSUBS 0.014956f
C214 VDD1.n184 VSUBS 0.027832f
C215 VDD1.n185 VSUBS 0.027832f
C216 VDD1.n186 VSUBS 0.014956f
C217 VDD1.n187 VSUBS 0.015835f
C218 VDD1.n188 VSUBS 0.03535f
C219 VDD1.n189 VSUBS 0.03535f
C220 VDD1.n190 VSUBS 0.015835f
C221 VDD1.n191 VSUBS 0.014956f
C222 VDD1.n192 VSUBS 0.027832f
C223 VDD1.n193 VSUBS 0.027832f
C224 VDD1.n194 VSUBS 0.014956f
C225 VDD1.n195 VSUBS 0.015835f
C226 VDD1.n196 VSUBS 0.03535f
C227 VDD1.n197 VSUBS 0.03535f
C228 VDD1.n198 VSUBS 0.015835f
C229 VDD1.n199 VSUBS 0.014956f
C230 VDD1.n200 VSUBS 0.027832f
C231 VDD1.n201 VSUBS 0.069275f
C232 VDD1.n202 VSUBS 0.014956f
C233 VDD1.n203 VSUBS 0.015835f
C234 VDD1.n204 VSUBS 0.077546f
C235 VDD1.n205 VSUBS 1.14072f
C236 VP.t0 VSUBS 5.97209f
C237 VP.t1 VSUBS 5.31075f
C238 VP.n0 VSUBS 6.62974f
C239 VDD2.n0 VSUBS 0.015852f
C240 VDD2.n1 VSUBS 0.035812f
C241 VDD2.n2 VSUBS 0.016043f
C242 VDD2.n3 VSUBS 0.028196f
C243 VDD2.n4 VSUBS 0.015151f
C244 VDD2.n5 VSUBS 0.035812f
C245 VDD2.n6 VSUBS 0.016043f
C246 VDD2.n7 VSUBS 0.028196f
C247 VDD2.n8 VSUBS 0.015151f
C248 VDD2.n9 VSUBS 0.035812f
C249 VDD2.n10 VSUBS 0.016043f
C250 VDD2.n11 VSUBS 0.028196f
C251 VDD2.n12 VSUBS 0.015151f
C252 VDD2.n13 VSUBS 0.035812f
C253 VDD2.n14 VSUBS 0.016043f
C254 VDD2.n15 VSUBS 0.028196f
C255 VDD2.n16 VSUBS 0.015151f
C256 VDD2.n17 VSUBS 0.035812f
C257 VDD2.n18 VSUBS 0.016043f
C258 VDD2.n19 VSUBS 0.028196f
C259 VDD2.n20 VSUBS 0.015151f
C260 VDD2.n21 VSUBS 0.035812f
C261 VDD2.n22 VSUBS 0.015597f
C262 VDD2.n23 VSUBS 0.028196f
C263 VDD2.n24 VSUBS 0.016043f
C264 VDD2.n25 VSUBS 0.035812f
C265 VDD2.n26 VSUBS 0.016043f
C266 VDD2.n27 VSUBS 0.028196f
C267 VDD2.n28 VSUBS 0.015151f
C268 VDD2.n29 VSUBS 0.035812f
C269 VDD2.n30 VSUBS 0.016043f
C270 VDD2.n31 VSUBS 2.21683f
C271 VDD2.n32 VSUBS 0.015151f
C272 VDD2.t1 VSUBS 0.077812f
C273 VDD2.n33 VSUBS 0.307862f
C274 VDD2.n34 VSUBS 0.02694f
C275 VDD2.n35 VSUBS 0.026859f
C276 VDD2.n36 VSUBS 0.035812f
C277 VDD2.n37 VSUBS 0.016043f
C278 VDD2.n38 VSUBS 0.015151f
C279 VDD2.n39 VSUBS 0.028196f
C280 VDD2.n40 VSUBS 0.028196f
C281 VDD2.n41 VSUBS 0.015151f
C282 VDD2.n42 VSUBS 0.016043f
C283 VDD2.n43 VSUBS 0.035812f
C284 VDD2.n44 VSUBS 0.035812f
C285 VDD2.n45 VSUBS 0.016043f
C286 VDD2.n46 VSUBS 0.015151f
C287 VDD2.n47 VSUBS 0.028196f
C288 VDD2.n48 VSUBS 0.028196f
C289 VDD2.n49 VSUBS 0.015151f
C290 VDD2.n50 VSUBS 0.015151f
C291 VDD2.n51 VSUBS 0.016043f
C292 VDD2.n52 VSUBS 0.035812f
C293 VDD2.n53 VSUBS 0.035812f
C294 VDD2.n54 VSUBS 0.035812f
C295 VDD2.n55 VSUBS 0.015597f
C296 VDD2.n56 VSUBS 0.015151f
C297 VDD2.n57 VSUBS 0.028196f
C298 VDD2.n58 VSUBS 0.028196f
C299 VDD2.n59 VSUBS 0.015151f
C300 VDD2.n60 VSUBS 0.016043f
C301 VDD2.n61 VSUBS 0.035812f
C302 VDD2.n62 VSUBS 0.035812f
C303 VDD2.n63 VSUBS 0.016043f
C304 VDD2.n64 VSUBS 0.015151f
C305 VDD2.n65 VSUBS 0.028196f
C306 VDD2.n66 VSUBS 0.028196f
C307 VDD2.n67 VSUBS 0.015151f
C308 VDD2.n68 VSUBS 0.016043f
C309 VDD2.n69 VSUBS 0.035812f
C310 VDD2.n70 VSUBS 0.035812f
C311 VDD2.n71 VSUBS 0.016043f
C312 VDD2.n72 VSUBS 0.015151f
C313 VDD2.n73 VSUBS 0.028196f
C314 VDD2.n74 VSUBS 0.028196f
C315 VDD2.n75 VSUBS 0.015151f
C316 VDD2.n76 VSUBS 0.016043f
C317 VDD2.n77 VSUBS 0.035812f
C318 VDD2.n78 VSUBS 0.035812f
C319 VDD2.n79 VSUBS 0.016043f
C320 VDD2.n80 VSUBS 0.015151f
C321 VDD2.n81 VSUBS 0.028196f
C322 VDD2.n82 VSUBS 0.028196f
C323 VDD2.n83 VSUBS 0.015151f
C324 VDD2.n84 VSUBS 0.016043f
C325 VDD2.n85 VSUBS 0.035812f
C326 VDD2.n86 VSUBS 0.035812f
C327 VDD2.n87 VSUBS 0.016043f
C328 VDD2.n88 VSUBS 0.015151f
C329 VDD2.n89 VSUBS 0.028196f
C330 VDD2.n90 VSUBS 0.028196f
C331 VDD2.n91 VSUBS 0.015151f
C332 VDD2.n92 VSUBS 0.016043f
C333 VDD2.n93 VSUBS 0.035812f
C334 VDD2.n94 VSUBS 0.035812f
C335 VDD2.n95 VSUBS 0.016043f
C336 VDD2.n96 VSUBS 0.015151f
C337 VDD2.n97 VSUBS 0.028196f
C338 VDD2.n98 VSUBS 0.070182f
C339 VDD2.n99 VSUBS 0.015151f
C340 VDD2.n100 VSUBS 0.016043f
C341 VDD2.n101 VSUBS 0.078561f
C342 VDD2.n102 VSUBS 1.09602f
C343 VDD2.n103 VSUBS 0.015852f
C344 VDD2.n104 VSUBS 0.035812f
C345 VDD2.n105 VSUBS 0.016043f
C346 VDD2.n106 VSUBS 0.028196f
C347 VDD2.n107 VSUBS 0.015151f
C348 VDD2.n108 VSUBS 0.035812f
C349 VDD2.n109 VSUBS 0.016043f
C350 VDD2.n110 VSUBS 0.028196f
C351 VDD2.n111 VSUBS 0.015151f
C352 VDD2.n112 VSUBS 0.035812f
C353 VDD2.n113 VSUBS 0.016043f
C354 VDD2.n114 VSUBS 0.028196f
C355 VDD2.n115 VSUBS 0.015151f
C356 VDD2.n116 VSUBS 0.035812f
C357 VDD2.n117 VSUBS 0.016043f
C358 VDD2.n118 VSUBS 0.028196f
C359 VDD2.n119 VSUBS 0.015151f
C360 VDD2.n120 VSUBS 0.035812f
C361 VDD2.n121 VSUBS 0.016043f
C362 VDD2.n122 VSUBS 0.028196f
C363 VDD2.n123 VSUBS 0.015151f
C364 VDD2.n124 VSUBS 0.035812f
C365 VDD2.n125 VSUBS 0.015597f
C366 VDD2.n126 VSUBS 0.028196f
C367 VDD2.n127 VSUBS 0.015597f
C368 VDD2.n128 VSUBS 0.015151f
C369 VDD2.n129 VSUBS 0.035812f
C370 VDD2.n130 VSUBS 0.035812f
C371 VDD2.n131 VSUBS 0.016043f
C372 VDD2.n132 VSUBS 0.028196f
C373 VDD2.n133 VSUBS 0.015151f
C374 VDD2.n134 VSUBS 0.035812f
C375 VDD2.n135 VSUBS 0.016043f
C376 VDD2.n136 VSUBS 2.21683f
C377 VDD2.n137 VSUBS 0.015151f
C378 VDD2.t0 VSUBS 0.077812f
C379 VDD2.n138 VSUBS 0.307862f
C380 VDD2.n139 VSUBS 0.02694f
C381 VDD2.n140 VSUBS 0.026859f
C382 VDD2.n141 VSUBS 0.035812f
C383 VDD2.n142 VSUBS 0.016043f
C384 VDD2.n143 VSUBS 0.015151f
C385 VDD2.n144 VSUBS 0.028196f
C386 VDD2.n145 VSUBS 0.028196f
C387 VDD2.n146 VSUBS 0.015151f
C388 VDD2.n147 VSUBS 0.016043f
C389 VDD2.n148 VSUBS 0.035812f
C390 VDD2.n149 VSUBS 0.035812f
C391 VDD2.n150 VSUBS 0.016043f
C392 VDD2.n151 VSUBS 0.015151f
C393 VDD2.n152 VSUBS 0.028196f
C394 VDD2.n153 VSUBS 0.028196f
C395 VDD2.n154 VSUBS 0.015151f
C396 VDD2.n155 VSUBS 0.016043f
C397 VDD2.n156 VSUBS 0.035812f
C398 VDD2.n157 VSUBS 0.035812f
C399 VDD2.n158 VSUBS 0.016043f
C400 VDD2.n159 VSUBS 0.015151f
C401 VDD2.n160 VSUBS 0.028196f
C402 VDD2.n161 VSUBS 0.028196f
C403 VDD2.n162 VSUBS 0.015151f
C404 VDD2.n163 VSUBS 0.016043f
C405 VDD2.n164 VSUBS 0.035812f
C406 VDD2.n165 VSUBS 0.035812f
C407 VDD2.n166 VSUBS 0.016043f
C408 VDD2.n167 VSUBS 0.015151f
C409 VDD2.n168 VSUBS 0.028196f
C410 VDD2.n169 VSUBS 0.028196f
C411 VDD2.n170 VSUBS 0.015151f
C412 VDD2.n171 VSUBS 0.016043f
C413 VDD2.n172 VSUBS 0.035812f
C414 VDD2.n173 VSUBS 0.035812f
C415 VDD2.n174 VSUBS 0.016043f
C416 VDD2.n175 VSUBS 0.015151f
C417 VDD2.n176 VSUBS 0.028196f
C418 VDD2.n177 VSUBS 0.028196f
C419 VDD2.n178 VSUBS 0.015151f
C420 VDD2.n179 VSUBS 0.016043f
C421 VDD2.n180 VSUBS 0.035812f
C422 VDD2.n181 VSUBS 0.035812f
C423 VDD2.n182 VSUBS 0.016043f
C424 VDD2.n183 VSUBS 0.015151f
C425 VDD2.n184 VSUBS 0.028196f
C426 VDD2.n185 VSUBS 0.028196f
C427 VDD2.n186 VSUBS 0.015151f
C428 VDD2.n187 VSUBS 0.016043f
C429 VDD2.n188 VSUBS 0.035812f
C430 VDD2.n189 VSUBS 0.035812f
C431 VDD2.n190 VSUBS 0.016043f
C432 VDD2.n191 VSUBS 0.015151f
C433 VDD2.n192 VSUBS 0.028196f
C434 VDD2.n193 VSUBS 0.028196f
C435 VDD2.n194 VSUBS 0.015151f
C436 VDD2.n195 VSUBS 0.016043f
C437 VDD2.n196 VSUBS 0.035812f
C438 VDD2.n197 VSUBS 0.035812f
C439 VDD2.n198 VSUBS 0.016043f
C440 VDD2.n199 VSUBS 0.015151f
C441 VDD2.n200 VSUBS 0.028196f
C442 VDD2.n201 VSUBS 0.070182f
C443 VDD2.n202 VSUBS 0.015151f
C444 VDD2.n203 VSUBS 0.016043f
C445 VDD2.n204 VSUBS 0.078561f
C446 VDD2.n205 VSUBS 0.071018f
C447 VDD2.n206 VSUBS 4.22868f
C448 VTAIL.n0 VSUBS 0.015669f
C449 VTAIL.n1 VSUBS 0.035399f
C450 VTAIL.n2 VSUBS 0.015858f
C451 VTAIL.n3 VSUBS 0.027871f
C452 VTAIL.n4 VSUBS 0.014977f
C453 VTAIL.n5 VSUBS 0.035399f
C454 VTAIL.n6 VSUBS 0.015858f
C455 VTAIL.n7 VSUBS 0.027871f
C456 VTAIL.n8 VSUBS 0.014977f
C457 VTAIL.n9 VSUBS 0.035399f
C458 VTAIL.n10 VSUBS 0.015858f
C459 VTAIL.n11 VSUBS 0.027871f
C460 VTAIL.n12 VSUBS 0.014977f
C461 VTAIL.n13 VSUBS 0.035399f
C462 VTAIL.n14 VSUBS 0.015858f
C463 VTAIL.n15 VSUBS 0.027871f
C464 VTAIL.n16 VSUBS 0.014977f
C465 VTAIL.n17 VSUBS 0.035399f
C466 VTAIL.n18 VSUBS 0.015858f
C467 VTAIL.n19 VSUBS 0.027871f
C468 VTAIL.n20 VSUBS 0.014977f
C469 VTAIL.n21 VSUBS 0.035399f
C470 VTAIL.n22 VSUBS 0.015417f
C471 VTAIL.n23 VSUBS 0.027871f
C472 VTAIL.n24 VSUBS 0.015858f
C473 VTAIL.n25 VSUBS 0.035399f
C474 VTAIL.n26 VSUBS 0.015858f
C475 VTAIL.n27 VSUBS 0.027871f
C476 VTAIL.n28 VSUBS 0.014977f
C477 VTAIL.n29 VSUBS 0.035399f
C478 VTAIL.n30 VSUBS 0.015858f
C479 VTAIL.n31 VSUBS 2.19124f
C480 VTAIL.n32 VSUBS 0.014977f
C481 VTAIL.t0 VSUBS 0.076914f
C482 VTAIL.n33 VSUBS 0.304309f
C483 VTAIL.n34 VSUBS 0.026629f
C484 VTAIL.n35 VSUBS 0.026549f
C485 VTAIL.n36 VSUBS 0.035399f
C486 VTAIL.n37 VSUBS 0.015858f
C487 VTAIL.n38 VSUBS 0.014977f
C488 VTAIL.n39 VSUBS 0.027871f
C489 VTAIL.n40 VSUBS 0.027871f
C490 VTAIL.n41 VSUBS 0.014977f
C491 VTAIL.n42 VSUBS 0.015858f
C492 VTAIL.n43 VSUBS 0.035399f
C493 VTAIL.n44 VSUBS 0.035399f
C494 VTAIL.n45 VSUBS 0.015858f
C495 VTAIL.n46 VSUBS 0.014977f
C496 VTAIL.n47 VSUBS 0.027871f
C497 VTAIL.n48 VSUBS 0.027871f
C498 VTAIL.n49 VSUBS 0.014977f
C499 VTAIL.n50 VSUBS 0.014977f
C500 VTAIL.n51 VSUBS 0.015858f
C501 VTAIL.n52 VSUBS 0.035399f
C502 VTAIL.n53 VSUBS 0.035399f
C503 VTAIL.n54 VSUBS 0.035399f
C504 VTAIL.n55 VSUBS 0.015417f
C505 VTAIL.n56 VSUBS 0.014977f
C506 VTAIL.n57 VSUBS 0.027871f
C507 VTAIL.n58 VSUBS 0.027871f
C508 VTAIL.n59 VSUBS 0.014977f
C509 VTAIL.n60 VSUBS 0.015858f
C510 VTAIL.n61 VSUBS 0.035399f
C511 VTAIL.n62 VSUBS 0.035399f
C512 VTAIL.n63 VSUBS 0.015858f
C513 VTAIL.n64 VSUBS 0.014977f
C514 VTAIL.n65 VSUBS 0.027871f
C515 VTAIL.n66 VSUBS 0.027871f
C516 VTAIL.n67 VSUBS 0.014977f
C517 VTAIL.n68 VSUBS 0.015858f
C518 VTAIL.n69 VSUBS 0.035399f
C519 VTAIL.n70 VSUBS 0.035399f
C520 VTAIL.n71 VSUBS 0.015858f
C521 VTAIL.n72 VSUBS 0.014977f
C522 VTAIL.n73 VSUBS 0.027871f
C523 VTAIL.n74 VSUBS 0.027871f
C524 VTAIL.n75 VSUBS 0.014977f
C525 VTAIL.n76 VSUBS 0.015858f
C526 VTAIL.n77 VSUBS 0.035399f
C527 VTAIL.n78 VSUBS 0.035399f
C528 VTAIL.n79 VSUBS 0.015858f
C529 VTAIL.n80 VSUBS 0.014977f
C530 VTAIL.n81 VSUBS 0.027871f
C531 VTAIL.n82 VSUBS 0.027871f
C532 VTAIL.n83 VSUBS 0.014977f
C533 VTAIL.n84 VSUBS 0.015858f
C534 VTAIL.n85 VSUBS 0.035399f
C535 VTAIL.n86 VSUBS 0.035399f
C536 VTAIL.n87 VSUBS 0.015858f
C537 VTAIL.n88 VSUBS 0.014977f
C538 VTAIL.n89 VSUBS 0.027871f
C539 VTAIL.n90 VSUBS 0.027871f
C540 VTAIL.n91 VSUBS 0.014977f
C541 VTAIL.n92 VSUBS 0.015858f
C542 VTAIL.n93 VSUBS 0.035399f
C543 VTAIL.n94 VSUBS 0.035399f
C544 VTAIL.n95 VSUBS 0.015858f
C545 VTAIL.n96 VSUBS 0.014977f
C546 VTAIL.n97 VSUBS 0.027871f
C547 VTAIL.n98 VSUBS 0.069372f
C548 VTAIL.n99 VSUBS 0.014977f
C549 VTAIL.n100 VSUBS 0.015858f
C550 VTAIL.n101 VSUBS 0.077654f
C551 VTAIL.n102 VSUBS 0.050986f
C552 VTAIL.n103 VSUBS 2.40391f
C553 VTAIL.n104 VSUBS 0.015669f
C554 VTAIL.n105 VSUBS 0.035399f
C555 VTAIL.n106 VSUBS 0.015858f
C556 VTAIL.n107 VSUBS 0.027871f
C557 VTAIL.n108 VSUBS 0.014977f
C558 VTAIL.n109 VSUBS 0.035399f
C559 VTAIL.n110 VSUBS 0.015858f
C560 VTAIL.n111 VSUBS 0.027871f
C561 VTAIL.n112 VSUBS 0.014977f
C562 VTAIL.n113 VSUBS 0.035399f
C563 VTAIL.n114 VSUBS 0.015858f
C564 VTAIL.n115 VSUBS 0.027871f
C565 VTAIL.n116 VSUBS 0.014977f
C566 VTAIL.n117 VSUBS 0.035399f
C567 VTAIL.n118 VSUBS 0.015858f
C568 VTAIL.n119 VSUBS 0.027871f
C569 VTAIL.n120 VSUBS 0.014977f
C570 VTAIL.n121 VSUBS 0.035399f
C571 VTAIL.n122 VSUBS 0.015858f
C572 VTAIL.n123 VSUBS 0.027871f
C573 VTAIL.n124 VSUBS 0.014977f
C574 VTAIL.n125 VSUBS 0.035399f
C575 VTAIL.n126 VSUBS 0.015417f
C576 VTAIL.n127 VSUBS 0.027871f
C577 VTAIL.n128 VSUBS 0.015417f
C578 VTAIL.n129 VSUBS 0.014977f
C579 VTAIL.n130 VSUBS 0.035399f
C580 VTAIL.n131 VSUBS 0.035399f
C581 VTAIL.n132 VSUBS 0.015858f
C582 VTAIL.n133 VSUBS 0.027871f
C583 VTAIL.n134 VSUBS 0.014977f
C584 VTAIL.n135 VSUBS 0.035399f
C585 VTAIL.n136 VSUBS 0.015858f
C586 VTAIL.n137 VSUBS 2.19124f
C587 VTAIL.n138 VSUBS 0.014977f
C588 VTAIL.t3 VSUBS 0.076914f
C589 VTAIL.n139 VSUBS 0.304309f
C590 VTAIL.n140 VSUBS 0.026629f
C591 VTAIL.n141 VSUBS 0.026549f
C592 VTAIL.n142 VSUBS 0.035399f
C593 VTAIL.n143 VSUBS 0.015858f
C594 VTAIL.n144 VSUBS 0.014977f
C595 VTAIL.n145 VSUBS 0.027871f
C596 VTAIL.n146 VSUBS 0.027871f
C597 VTAIL.n147 VSUBS 0.014977f
C598 VTAIL.n148 VSUBS 0.015858f
C599 VTAIL.n149 VSUBS 0.035399f
C600 VTAIL.n150 VSUBS 0.035399f
C601 VTAIL.n151 VSUBS 0.015858f
C602 VTAIL.n152 VSUBS 0.014977f
C603 VTAIL.n153 VSUBS 0.027871f
C604 VTAIL.n154 VSUBS 0.027871f
C605 VTAIL.n155 VSUBS 0.014977f
C606 VTAIL.n156 VSUBS 0.015858f
C607 VTAIL.n157 VSUBS 0.035399f
C608 VTAIL.n158 VSUBS 0.035399f
C609 VTAIL.n159 VSUBS 0.015858f
C610 VTAIL.n160 VSUBS 0.014977f
C611 VTAIL.n161 VSUBS 0.027871f
C612 VTAIL.n162 VSUBS 0.027871f
C613 VTAIL.n163 VSUBS 0.014977f
C614 VTAIL.n164 VSUBS 0.015858f
C615 VTAIL.n165 VSUBS 0.035399f
C616 VTAIL.n166 VSUBS 0.035399f
C617 VTAIL.n167 VSUBS 0.015858f
C618 VTAIL.n168 VSUBS 0.014977f
C619 VTAIL.n169 VSUBS 0.027871f
C620 VTAIL.n170 VSUBS 0.027871f
C621 VTAIL.n171 VSUBS 0.014977f
C622 VTAIL.n172 VSUBS 0.015858f
C623 VTAIL.n173 VSUBS 0.035399f
C624 VTAIL.n174 VSUBS 0.035399f
C625 VTAIL.n175 VSUBS 0.015858f
C626 VTAIL.n176 VSUBS 0.014977f
C627 VTAIL.n177 VSUBS 0.027871f
C628 VTAIL.n178 VSUBS 0.027871f
C629 VTAIL.n179 VSUBS 0.014977f
C630 VTAIL.n180 VSUBS 0.015858f
C631 VTAIL.n181 VSUBS 0.035399f
C632 VTAIL.n182 VSUBS 0.035399f
C633 VTAIL.n183 VSUBS 0.015858f
C634 VTAIL.n184 VSUBS 0.014977f
C635 VTAIL.n185 VSUBS 0.027871f
C636 VTAIL.n186 VSUBS 0.027871f
C637 VTAIL.n187 VSUBS 0.014977f
C638 VTAIL.n188 VSUBS 0.015858f
C639 VTAIL.n189 VSUBS 0.035399f
C640 VTAIL.n190 VSUBS 0.035399f
C641 VTAIL.n191 VSUBS 0.015858f
C642 VTAIL.n192 VSUBS 0.014977f
C643 VTAIL.n193 VSUBS 0.027871f
C644 VTAIL.n194 VSUBS 0.027871f
C645 VTAIL.n195 VSUBS 0.014977f
C646 VTAIL.n196 VSUBS 0.015858f
C647 VTAIL.n197 VSUBS 0.035399f
C648 VTAIL.n198 VSUBS 0.035399f
C649 VTAIL.n199 VSUBS 0.015858f
C650 VTAIL.n200 VSUBS 0.014977f
C651 VTAIL.n201 VSUBS 0.027871f
C652 VTAIL.n202 VSUBS 0.069372f
C653 VTAIL.n203 VSUBS 0.014977f
C654 VTAIL.n204 VSUBS 0.015858f
C655 VTAIL.n205 VSUBS 0.077654f
C656 VTAIL.n206 VSUBS 0.050986f
C657 VTAIL.n207 VSUBS 2.45443f
C658 VTAIL.n208 VSUBS 0.015669f
C659 VTAIL.n209 VSUBS 0.035399f
C660 VTAIL.n210 VSUBS 0.015858f
C661 VTAIL.n211 VSUBS 0.027871f
C662 VTAIL.n212 VSUBS 0.014977f
C663 VTAIL.n213 VSUBS 0.035399f
C664 VTAIL.n214 VSUBS 0.015858f
C665 VTAIL.n215 VSUBS 0.027871f
C666 VTAIL.n216 VSUBS 0.014977f
C667 VTAIL.n217 VSUBS 0.035399f
C668 VTAIL.n218 VSUBS 0.015858f
C669 VTAIL.n219 VSUBS 0.027871f
C670 VTAIL.n220 VSUBS 0.014977f
C671 VTAIL.n221 VSUBS 0.035399f
C672 VTAIL.n222 VSUBS 0.015858f
C673 VTAIL.n223 VSUBS 0.027871f
C674 VTAIL.n224 VSUBS 0.014977f
C675 VTAIL.n225 VSUBS 0.035399f
C676 VTAIL.n226 VSUBS 0.015858f
C677 VTAIL.n227 VSUBS 0.027871f
C678 VTAIL.n228 VSUBS 0.014977f
C679 VTAIL.n229 VSUBS 0.035399f
C680 VTAIL.n230 VSUBS 0.015417f
C681 VTAIL.n231 VSUBS 0.027871f
C682 VTAIL.n232 VSUBS 0.015417f
C683 VTAIL.n233 VSUBS 0.014977f
C684 VTAIL.n234 VSUBS 0.035399f
C685 VTAIL.n235 VSUBS 0.035399f
C686 VTAIL.n236 VSUBS 0.015858f
C687 VTAIL.n237 VSUBS 0.027871f
C688 VTAIL.n238 VSUBS 0.014977f
C689 VTAIL.n239 VSUBS 0.035399f
C690 VTAIL.n240 VSUBS 0.015858f
C691 VTAIL.n241 VSUBS 2.19124f
C692 VTAIL.n242 VSUBS 0.014977f
C693 VTAIL.t1 VSUBS 0.076914f
C694 VTAIL.n243 VSUBS 0.304309f
C695 VTAIL.n244 VSUBS 0.026629f
C696 VTAIL.n245 VSUBS 0.026549f
C697 VTAIL.n246 VSUBS 0.035399f
C698 VTAIL.n247 VSUBS 0.015858f
C699 VTAIL.n248 VSUBS 0.014977f
C700 VTAIL.n249 VSUBS 0.027871f
C701 VTAIL.n250 VSUBS 0.027871f
C702 VTAIL.n251 VSUBS 0.014977f
C703 VTAIL.n252 VSUBS 0.015858f
C704 VTAIL.n253 VSUBS 0.035399f
C705 VTAIL.n254 VSUBS 0.035399f
C706 VTAIL.n255 VSUBS 0.015858f
C707 VTAIL.n256 VSUBS 0.014977f
C708 VTAIL.n257 VSUBS 0.027871f
C709 VTAIL.n258 VSUBS 0.027871f
C710 VTAIL.n259 VSUBS 0.014977f
C711 VTAIL.n260 VSUBS 0.015858f
C712 VTAIL.n261 VSUBS 0.035399f
C713 VTAIL.n262 VSUBS 0.035399f
C714 VTAIL.n263 VSUBS 0.015858f
C715 VTAIL.n264 VSUBS 0.014977f
C716 VTAIL.n265 VSUBS 0.027871f
C717 VTAIL.n266 VSUBS 0.027871f
C718 VTAIL.n267 VSUBS 0.014977f
C719 VTAIL.n268 VSUBS 0.015858f
C720 VTAIL.n269 VSUBS 0.035399f
C721 VTAIL.n270 VSUBS 0.035399f
C722 VTAIL.n271 VSUBS 0.015858f
C723 VTAIL.n272 VSUBS 0.014977f
C724 VTAIL.n273 VSUBS 0.027871f
C725 VTAIL.n274 VSUBS 0.027871f
C726 VTAIL.n275 VSUBS 0.014977f
C727 VTAIL.n276 VSUBS 0.015858f
C728 VTAIL.n277 VSUBS 0.035399f
C729 VTAIL.n278 VSUBS 0.035399f
C730 VTAIL.n279 VSUBS 0.015858f
C731 VTAIL.n280 VSUBS 0.014977f
C732 VTAIL.n281 VSUBS 0.027871f
C733 VTAIL.n282 VSUBS 0.027871f
C734 VTAIL.n283 VSUBS 0.014977f
C735 VTAIL.n284 VSUBS 0.015858f
C736 VTAIL.n285 VSUBS 0.035399f
C737 VTAIL.n286 VSUBS 0.035399f
C738 VTAIL.n287 VSUBS 0.015858f
C739 VTAIL.n288 VSUBS 0.014977f
C740 VTAIL.n289 VSUBS 0.027871f
C741 VTAIL.n290 VSUBS 0.027871f
C742 VTAIL.n291 VSUBS 0.014977f
C743 VTAIL.n292 VSUBS 0.015858f
C744 VTAIL.n293 VSUBS 0.035399f
C745 VTAIL.n294 VSUBS 0.035399f
C746 VTAIL.n295 VSUBS 0.015858f
C747 VTAIL.n296 VSUBS 0.014977f
C748 VTAIL.n297 VSUBS 0.027871f
C749 VTAIL.n298 VSUBS 0.027871f
C750 VTAIL.n299 VSUBS 0.014977f
C751 VTAIL.n300 VSUBS 0.015858f
C752 VTAIL.n301 VSUBS 0.035399f
C753 VTAIL.n302 VSUBS 0.035399f
C754 VTAIL.n303 VSUBS 0.015858f
C755 VTAIL.n304 VSUBS 0.014977f
C756 VTAIL.n305 VSUBS 0.027871f
C757 VTAIL.n306 VSUBS 0.069372f
C758 VTAIL.n307 VSUBS 0.014977f
C759 VTAIL.n308 VSUBS 0.015858f
C760 VTAIL.n309 VSUBS 0.077654f
C761 VTAIL.n310 VSUBS 0.050986f
C762 VTAIL.n311 VSUBS 2.23146f
C763 VTAIL.n312 VSUBS 0.015669f
C764 VTAIL.n313 VSUBS 0.035399f
C765 VTAIL.n314 VSUBS 0.015858f
C766 VTAIL.n315 VSUBS 0.027871f
C767 VTAIL.n316 VSUBS 0.014977f
C768 VTAIL.n317 VSUBS 0.035399f
C769 VTAIL.n318 VSUBS 0.015858f
C770 VTAIL.n319 VSUBS 0.027871f
C771 VTAIL.n320 VSUBS 0.014977f
C772 VTAIL.n321 VSUBS 0.035399f
C773 VTAIL.n322 VSUBS 0.015858f
C774 VTAIL.n323 VSUBS 0.027871f
C775 VTAIL.n324 VSUBS 0.014977f
C776 VTAIL.n325 VSUBS 0.035399f
C777 VTAIL.n326 VSUBS 0.015858f
C778 VTAIL.n327 VSUBS 0.027871f
C779 VTAIL.n328 VSUBS 0.014977f
C780 VTAIL.n329 VSUBS 0.035399f
C781 VTAIL.n330 VSUBS 0.015858f
C782 VTAIL.n331 VSUBS 0.027871f
C783 VTAIL.n332 VSUBS 0.014977f
C784 VTAIL.n333 VSUBS 0.035399f
C785 VTAIL.n334 VSUBS 0.015417f
C786 VTAIL.n335 VSUBS 0.027871f
C787 VTAIL.n336 VSUBS 0.015858f
C788 VTAIL.n337 VSUBS 0.035399f
C789 VTAIL.n338 VSUBS 0.015858f
C790 VTAIL.n339 VSUBS 0.027871f
C791 VTAIL.n340 VSUBS 0.014977f
C792 VTAIL.n341 VSUBS 0.035399f
C793 VTAIL.n342 VSUBS 0.015858f
C794 VTAIL.n343 VSUBS 2.19124f
C795 VTAIL.n344 VSUBS 0.014977f
C796 VTAIL.t2 VSUBS 0.076914f
C797 VTAIL.n345 VSUBS 0.304309f
C798 VTAIL.n346 VSUBS 0.026629f
C799 VTAIL.n347 VSUBS 0.026549f
C800 VTAIL.n348 VSUBS 0.035399f
C801 VTAIL.n349 VSUBS 0.015858f
C802 VTAIL.n350 VSUBS 0.014977f
C803 VTAIL.n351 VSUBS 0.027871f
C804 VTAIL.n352 VSUBS 0.027871f
C805 VTAIL.n353 VSUBS 0.014977f
C806 VTAIL.n354 VSUBS 0.015858f
C807 VTAIL.n355 VSUBS 0.035399f
C808 VTAIL.n356 VSUBS 0.035399f
C809 VTAIL.n357 VSUBS 0.015858f
C810 VTAIL.n358 VSUBS 0.014977f
C811 VTAIL.n359 VSUBS 0.027871f
C812 VTAIL.n360 VSUBS 0.027871f
C813 VTAIL.n361 VSUBS 0.014977f
C814 VTAIL.n362 VSUBS 0.014977f
C815 VTAIL.n363 VSUBS 0.015858f
C816 VTAIL.n364 VSUBS 0.035399f
C817 VTAIL.n365 VSUBS 0.035399f
C818 VTAIL.n366 VSUBS 0.035399f
C819 VTAIL.n367 VSUBS 0.015417f
C820 VTAIL.n368 VSUBS 0.014977f
C821 VTAIL.n369 VSUBS 0.027871f
C822 VTAIL.n370 VSUBS 0.027871f
C823 VTAIL.n371 VSUBS 0.014977f
C824 VTAIL.n372 VSUBS 0.015858f
C825 VTAIL.n373 VSUBS 0.035399f
C826 VTAIL.n374 VSUBS 0.035399f
C827 VTAIL.n375 VSUBS 0.015858f
C828 VTAIL.n376 VSUBS 0.014977f
C829 VTAIL.n377 VSUBS 0.027871f
C830 VTAIL.n378 VSUBS 0.027871f
C831 VTAIL.n379 VSUBS 0.014977f
C832 VTAIL.n380 VSUBS 0.015858f
C833 VTAIL.n381 VSUBS 0.035399f
C834 VTAIL.n382 VSUBS 0.035399f
C835 VTAIL.n383 VSUBS 0.015858f
C836 VTAIL.n384 VSUBS 0.014977f
C837 VTAIL.n385 VSUBS 0.027871f
C838 VTAIL.n386 VSUBS 0.027871f
C839 VTAIL.n387 VSUBS 0.014977f
C840 VTAIL.n388 VSUBS 0.015858f
C841 VTAIL.n389 VSUBS 0.035399f
C842 VTAIL.n390 VSUBS 0.035399f
C843 VTAIL.n391 VSUBS 0.015858f
C844 VTAIL.n392 VSUBS 0.014977f
C845 VTAIL.n393 VSUBS 0.027871f
C846 VTAIL.n394 VSUBS 0.027871f
C847 VTAIL.n395 VSUBS 0.014977f
C848 VTAIL.n396 VSUBS 0.015858f
C849 VTAIL.n397 VSUBS 0.035399f
C850 VTAIL.n398 VSUBS 0.035399f
C851 VTAIL.n399 VSUBS 0.015858f
C852 VTAIL.n400 VSUBS 0.014977f
C853 VTAIL.n401 VSUBS 0.027871f
C854 VTAIL.n402 VSUBS 0.027871f
C855 VTAIL.n403 VSUBS 0.014977f
C856 VTAIL.n404 VSUBS 0.015858f
C857 VTAIL.n405 VSUBS 0.035399f
C858 VTAIL.n406 VSUBS 0.035399f
C859 VTAIL.n407 VSUBS 0.015858f
C860 VTAIL.n408 VSUBS 0.014977f
C861 VTAIL.n409 VSUBS 0.027871f
C862 VTAIL.n410 VSUBS 0.069372f
C863 VTAIL.n411 VSUBS 0.014977f
C864 VTAIL.n412 VSUBS 0.015858f
C865 VTAIL.n413 VSUBS 0.077654f
C866 VTAIL.n414 VSUBS 0.050986f
C867 VTAIL.n415 VSUBS 2.1283f
C868 VN.t0 VSUBS 5.12126f
C869 VN.t1 VSUBS 5.75946f
C870 B.n0 VSUBS 0.004326f
C871 B.n1 VSUBS 0.004326f
C872 B.n2 VSUBS 0.006841f
C873 B.n3 VSUBS 0.006841f
C874 B.n4 VSUBS 0.006841f
C875 B.n5 VSUBS 0.006841f
C876 B.n6 VSUBS 0.006841f
C877 B.n7 VSUBS 0.006841f
C878 B.n8 VSUBS 0.006841f
C879 B.n9 VSUBS 0.006841f
C880 B.n10 VSUBS 0.006841f
C881 B.n11 VSUBS 0.006841f
C882 B.n12 VSUBS 0.006841f
C883 B.n13 VSUBS 0.006841f
C884 B.n14 VSUBS 0.016535f
C885 B.n15 VSUBS 0.006841f
C886 B.n16 VSUBS 0.006841f
C887 B.n17 VSUBS 0.006841f
C888 B.n18 VSUBS 0.006841f
C889 B.n19 VSUBS 0.006841f
C890 B.n20 VSUBS 0.006841f
C891 B.n21 VSUBS 0.006841f
C892 B.n22 VSUBS 0.006841f
C893 B.n23 VSUBS 0.006841f
C894 B.n24 VSUBS 0.006841f
C895 B.n25 VSUBS 0.006841f
C896 B.n26 VSUBS 0.006841f
C897 B.n27 VSUBS 0.006841f
C898 B.n28 VSUBS 0.006841f
C899 B.n29 VSUBS 0.006841f
C900 B.n30 VSUBS 0.006841f
C901 B.n31 VSUBS 0.006841f
C902 B.n32 VSUBS 0.006841f
C903 B.n33 VSUBS 0.006841f
C904 B.n34 VSUBS 0.006841f
C905 B.n35 VSUBS 0.006841f
C906 B.n36 VSUBS 0.006841f
C907 B.n37 VSUBS 0.006841f
C908 B.n38 VSUBS 0.006841f
C909 B.n39 VSUBS 0.006841f
C910 B.n40 VSUBS 0.006841f
C911 B.n41 VSUBS 0.006841f
C912 B.n42 VSUBS 0.006841f
C913 B.n43 VSUBS 0.006841f
C914 B.n44 VSUBS 0.006841f
C915 B.n45 VSUBS 0.006841f
C916 B.t8 VSUBS 0.360218f
C917 B.t7 VSUBS 0.392566f
C918 B.t6 VSUBS 2.0619f
C919 B.n46 VSUBS 0.598316f
C920 B.n47 VSUBS 0.329734f
C921 B.n48 VSUBS 0.006841f
C922 B.n49 VSUBS 0.006841f
C923 B.n50 VSUBS 0.006841f
C924 B.n51 VSUBS 0.006841f
C925 B.t5 VSUBS 0.360222f
C926 B.t4 VSUBS 0.392569f
C927 B.t3 VSUBS 2.0619f
C928 B.n52 VSUBS 0.598313f
C929 B.n53 VSUBS 0.329731f
C930 B.n54 VSUBS 0.01585f
C931 B.n55 VSUBS 0.006841f
C932 B.n56 VSUBS 0.006841f
C933 B.n57 VSUBS 0.006841f
C934 B.n58 VSUBS 0.006841f
C935 B.n59 VSUBS 0.006841f
C936 B.n60 VSUBS 0.006841f
C937 B.n61 VSUBS 0.006841f
C938 B.n62 VSUBS 0.006841f
C939 B.n63 VSUBS 0.006841f
C940 B.n64 VSUBS 0.006841f
C941 B.n65 VSUBS 0.006841f
C942 B.n66 VSUBS 0.006841f
C943 B.n67 VSUBS 0.006841f
C944 B.n68 VSUBS 0.006841f
C945 B.n69 VSUBS 0.006841f
C946 B.n70 VSUBS 0.006841f
C947 B.n71 VSUBS 0.006841f
C948 B.n72 VSUBS 0.006841f
C949 B.n73 VSUBS 0.006841f
C950 B.n74 VSUBS 0.006841f
C951 B.n75 VSUBS 0.006841f
C952 B.n76 VSUBS 0.006841f
C953 B.n77 VSUBS 0.006841f
C954 B.n78 VSUBS 0.006841f
C955 B.n79 VSUBS 0.006841f
C956 B.n80 VSUBS 0.006841f
C957 B.n81 VSUBS 0.006841f
C958 B.n82 VSUBS 0.006841f
C959 B.n83 VSUBS 0.006841f
C960 B.n84 VSUBS 0.006841f
C961 B.n85 VSUBS 0.016535f
C962 B.n86 VSUBS 0.006841f
C963 B.n87 VSUBS 0.006841f
C964 B.n88 VSUBS 0.006841f
C965 B.n89 VSUBS 0.006841f
C966 B.n90 VSUBS 0.006841f
C967 B.n91 VSUBS 0.006841f
C968 B.n92 VSUBS 0.006841f
C969 B.n93 VSUBS 0.006841f
C970 B.n94 VSUBS 0.006841f
C971 B.n95 VSUBS 0.006841f
C972 B.n96 VSUBS 0.006841f
C973 B.n97 VSUBS 0.006841f
C974 B.n98 VSUBS 0.006841f
C975 B.n99 VSUBS 0.006841f
C976 B.n100 VSUBS 0.006841f
C977 B.n101 VSUBS 0.006841f
C978 B.n102 VSUBS 0.006841f
C979 B.n103 VSUBS 0.006841f
C980 B.n104 VSUBS 0.006841f
C981 B.n105 VSUBS 0.006841f
C982 B.n106 VSUBS 0.006841f
C983 B.n107 VSUBS 0.006841f
C984 B.n108 VSUBS 0.006841f
C985 B.n109 VSUBS 0.006841f
C986 B.n110 VSUBS 0.016535f
C987 B.n111 VSUBS 0.006841f
C988 B.n112 VSUBS 0.006841f
C989 B.n113 VSUBS 0.006841f
C990 B.n114 VSUBS 0.006841f
C991 B.n115 VSUBS 0.006841f
C992 B.n116 VSUBS 0.006841f
C993 B.n117 VSUBS 0.006841f
C994 B.n118 VSUBS 0.006841f
C995 B.n119 VSUBS 0.006841f
C996 B.n120 VSUBS 0.006841f
C997 B.n121 VSUBS 0.006841f
C998 B.n122 VSUBS 0.006841f
C999 B.n123 VSUBS 0.006841f
C1000 B.n124 VSUBS 0.006841f
C1001 B.n125 VSUBS 0.006841f
C1002 B.n126 VSUBS 0.006841f
C1003 B.n127 VSUBS 0.006841f
C1004 B.n128 VSUBS 0.006841f
C1005 B.n129 VSUBS 0.006841f
C1006 B.n130 VSUBS 0.006841f
C1007 B.n131 VSUBS 0.006841f
C1008 B.n132 VSUBS 0.006841f
C1009 B.n133 VSUBS 0.006841f
C1010 B.n134 VSUBS 0.006841f
C1011 B.n135 VSUBS 0.006841f
C1012 B.n136 VSUBS 0.006841f
C1013 B.n137 VSUBS 0.006841f
C1014 B.n138 VSUBS 0.006841f
C1015 B.n139 VSUBS 0.006841f
C1016 B.n140 VSUBS 0.006841f
C1017 B.n141 VSUBS 0.006841f
C1018 B.t1 VSUBS 0.360222f
C1019 B.t2 VSUBS 0.392569f
C1020 B.t0 VSUBS 2.0619f
C1021 B.n142 VSUBS 0.598313f
C1022 B.n143 VSUBS 0.329731f
C1023 B.n144 VSUBS 0.006841f
C1024 B.n145 VSUBS 0.006841f
C1025 B.n146 VSUBS 0.006841f
C1026 B.n147 VSUBS 0.006841f
C1027 B.t10 VSUBS 0.360218f
C1028 B.t11 VSUBS 0.392566f
C1029 B.t9 VSUBS 2.0619f
C1030 B.n148 VSUBS 0.598316f
C1031 B.n149 VSUBS 0.329734f
C1032 B.n150 VSUBS 0.01585f
C1033 B.n151 VSUBS 0.006841f
C1034 B.n152 VSUBS 0.006841f
C1035 B.n153 VSUBS 0.006841f
C1036 B.n154 VSUBS 0.006841f
C1037 B.n155 VSUBS 0.006841f
C1038 B.n156 VSUBS 0.006841f
C1039 B.n157 VSUBS 0.006841f
C1040 B.n158 VSUBS 0.006841f
C1041 B.n159 VSUBS 0.006841f
C1042 B.n160 VSUBS 0.006841f
C1043 B.n161 VSUBS 0.006841f
C1044 B.n162 VSUBS 0.006841f
C1045 B.n163 VSUBS 0.006841f
C1046 B.n164 VSUBS 0.006841f
C1047 B.n165 VSUBS 0.006841f
C1048 B.n166 VSUBS 0.006841f
C1049 B.n167 VSUBS 0.006841f
C1050 B.n168 VSUBS 0.006841f
C1051 B.n169 VSUBS 0.006841f
C1052 B.n170 VSUBS 0.006841f
C1053 B.n171 VSUBS 0.006841f
C1054 B.n172 VSUBS 0.006841f
C1055 B.n173 VSUBS 0.006841f
C1056 B.n174 VSUBS 0.006841f
C1057 B.n175 VSUBS 0.006841f
C1058 B.n176 VSUBS 0.006841f
C1059 B.n177 VSUBS 0.006841f
C1060 B.n178 VSUBS 0.006841f
C1061 B.n179 VSUBS 0.006841f
C1062 B.n180 VSUBS 0.006841f
C1063 B.n181 VSUBS 0.016535f
C1064 B.n182 VSUBS 0.006841f
C1065 B.n183 VSUBS 0.006841f
C1066 B.n184 VSUBS 0.006841f
C1067 B.n185 VSUBS 0.006841f
C1068 B.n186 VSUBS 0.006841f
C1069 B.n187 VSUBS 0.006841f
C1070 B.n188 VSUBS 0.006841f
C1071 B.n189 VSUBS 0.006841f
C1072 B.n190 VSUBS 0.006841f
C1073 B.n191 VSUBS 0.006841f
C1074 B.n192 VSUBS 0.006841f
C1075 B.n193 VSUBS 0.006841f
C1076 B.n194 VSUBS 0.006841f
C1077 B.n195 VSUBS 0.006841f
C1078 B.n196 VSUBS 0.006841f
C1079 B.n197 VSUBS 0.006841f
C1080 B.n198 VSUBS 0.006841f
C1081 B.n199 VSUBS 0.006841f
C1082 B.n200 VSUBS 0.006841f
C1083 B.n201 VSUBS 0.006841f
C1084 B.n202 VSUBS 0.006841f
C1085 B.n203 VSUBS 0.006841f
C1086 B.n204 VSUBS 0.006841f
C1087 B.n205 VSUBS 0.006841f
C1088 B.n206 VSUBS 0.006841f
C1089 B.n207 VSUBS 0.006841f
C1090 B.n208 VSUBS 0.006841f
C1091 B.n209 VSUBS 0.006841f
C1092 B.n210 VSUBS 0.006841f
C1093 B.n211 VSUBS 0.006841f
C1094 B.n212 VSUBS 0.006841f
C1095 B.n213 VSUBS 0.006841f
C1096 B.n214 VSUBS 0.006841f
C1097 B.n215 VSUBS 0.006841f
C1098 B.n216 VSUBS 0.006841f
C1099 B.n217 VSUBS 0.006841f
C1100 B.n218 VSUBS 0.006841f
C1101 B.n219 VSUBS 0.006841f
C1102 B.n220 VSUBS 0.006841f
C1103 B.n221 VSUBS 0.006841f
C1104 B.n222 VSUBS 0.006841f
C1105 B.n223 VSUBS 0.006841f
C1106 B.n224 VSUBS 0.006841f
C1107 B.n225 VSUBS 0.006841f
C1108 B.n226 VSUBS 0.006841f
C1109 B.n227 VSUBS 0.006841f
C1110 B.n228 VSUBS 0.016535f
C1111 B.n229 VSUBS 0.017067f
C1112 B.n230 VSUBS 0.017067f
C1113 B.n231 VSUBS 0.006841f
C1114 B.n232 VSUBS 0.006841f
C1115 B.n233 VSUBS 0.006841f
C1116 B.n234 VSUBS 0.006841f
C1117 B.n235 VSUBS 0.006841f
C1118 B.n236 VSUBS 0.006841f
C1119 B.n237 VSUBS 0.006841f
C1120 B.n238 VSUBS 0.006841f
C1121 B.n239 VSUBS 0.006841f
C1122 B.n240 VSUBS 0.006841f
C1123 B.n241 VSUBS 0.006841f
C1124 B.n242 VSUBS 0.006841f
C1125 B.n243 VSUBS 0.006841f
C1126 B.n244 VSUBS 0.006841f
C1127 B.n245 VSUBS 0.006841f
C1128 B.n246 VSUBS 0.006841f
C1129 B.n247 VSUBS 0.006841f
C1130 B.n248 VSUBS 0.006841f
C1131 B.n249 VSUBS 0.006841f
C1132 B.n250 VSUBS 0.006841f
C1133 B.n251 VSUBS 0.006841f
C1134 B.n252 VSUBS 0.006841f
C1135 B.n253 VSUBS 0.006841f
C1136 B.n254 VSUBS 0.006841f
C1137 B.n255 VSUBS 0.006841f
C1138 B.n256 VSUBS 0.006841f
C1139 B.n257 VSUBS 0.006841f
C1140 B.n258 VSUBS 0.006841f
C1141 B.n259 VSUBS 0.006841f
C1142 B.n260 VSUBS 0.006841f
C1143 B.n261 VSUBS 0.006841f
C1144 B.n262 VSUBS 0.006841f
C1145 B.n263 VSUBS 0.006841f
C1146 B.n264 VSUBS 0.006841f
C1147 B.n265 VSUBS 0.006841f
C1148 B.n266 VSUBS 0.006841f
C1149 B.n267 VSUBS 0.006841f
C1150 B.n268 VSUBS 0.006841f
C1151 B.n269 VSUBS 0.006841f
C1152 B.n270 VSUBS 0.006841f
C1153 B.n271 VSUBS 0.006841f
C1154 B.n272 VSUBS 0.006841f
C1155 B.n273 VSUBS 0.006841f
C1156 B.n274 VSUBS 0.006841f
C1157 B.n275 VSUBS 0.006841f
C1158 B.n276 VSUBS 0.006841f
C1159 B.n277 VSUBS 0.006841f
C1160 B.n278 VSUBS 0.006841f
C1161 B.n279 VSUBS 0.006841f
C1162 B.n280 VSUBS 0.006841f
C1163 B.n281 VSUBS 0.006841f
C1164 B.n282 VSUBS 0.006841f
C1165 B.n283 VSUBS 0.006841f
C1166 B.n284 VSUBS 0.006841f
C1167 B.n285 VSUBS 0.006841f
C1168 B.n286 VSUBS 0.006841f
C1169 B.n287 VSUBS 0.006841f
C1170 B.n288 VSUBS 0.006841f
C1171 B.n289 VSUBS 0.006841f
C1172 B.n290 VSUBS 0.006841f
C1173 B.n291 VSUBS 0.006841f
C1174 B.n292 VSUBS 0.006841f
C1175 B.n293 VSUBS 0.006841f
C1176 B.n294 VSUBS 0.006841f
C1177 B.n295 VSUBS 0.006841f
C1178 B.n296 VSUBS 0.006841f
C1179 B.n297 VSUBS 0.006841f
C1180 B.n298 VSUBS 0.006841f
C1181 B.n299 VSUBS 0.006841f
C1182 B.n300 VSUBS 0.006841f
C1183 B.n301 VSUBS 0.006841f
C1184 B.n302 VSUBS 0.006841f
C1185 B.n303 VSUBS 0.006841f
C1186 B.n304 VSUBS 0.006841f
C1187 B.n305 VSUBS 0.006841f
C1188 B.n306 VSUBS 0.006841f
C1189 B.n307 VSUBS 0.006841f
C1190 B.n308 VSUBS 0.006841f
C1191 B.n309 VSUBS 0.006841f
C1192 B.n310 VSUBS 0.006841f
C1193 B.n311 VSUBS 0.006841f
C1194 B.n312 VSUBS 0.006841f
C1195 B.n313 VSUBS 0.006841f
C1196 B.n314 VSUBS 0.006841f
C1197 B.n315 VSUBS 0.006841f
C1198 B.n316 VSUBS 0.006841f
C1199 B.n317 VSUBS 0.006841f
C1200 B.n318 VSUBS 0.006841f
C1201 B.n319 VSUBS 0.006439f
C1202 B.n320 VSUBS 0.006841f
C1203 B.n321 VSUBS 0.006841f
C1204 B.n322 VSUBS 0.003823f
C1205 B.n323 VSUBS 0.006841f
C1206 B.n324 VSUBS 0.006841f
C1207 B.n325 VSUBS 0.006841f
C1208 B.n326 VSUBS 0.006841f
C1209 B.n327 VSUBS 0.006841f
C1210 B.n328 VSUBS 0.006841f
C1211 B.n329 VSUBS 0.006841f
C1212 B.n330 VSUBS 0.006841f
C1213 B.n331 VSUBS 0.006841f
C1214 B.n332 VSUBS 0.006841f
C1215 B.n333 VSUBS 0.006841f
C1216 B.n334 VSUBS 0.006841f
C1217 B.n335 VSUBS 0.003823f
C1218 B.n336 VSUBS 0.01585f
C1219 B.n337 VSUBS 0.006439f
C1220 B.n338 VSUBS 0.006841f
C1221 B.n339 VSUBS 0.006841f
C1222 B.n340 VSUBS 0.006841f
C1223 B.n341 VSUBS 0.006841f
C1224 B.n342 VSUBS 0.006841f
C1225 B.n343 VSUBS 0.006841f
C1226 B.n344 VSUBS 0.006841f
C1227 B.n345 VSUBS 0.006841f
C1228 B.n346 VSUBS 0.006841f
C1229 B.n347 VSUBS 0.006841f
C1230 B.n348 VSUBS 0.006841f
C1231 B.n349 VSUBS 0.006841f
C1232 B.n350 VSUBS 0.006841f
C1233 B.n351 VSUBS 0.006841f
C1234 B.n352 VSUBS 0.006841f
C1235 B.n353 VSUBS 0.006841f
C1236 B.n354 VSUBS 0.006841f
C1237 B.n355 VSUBS 0.006841f
C1238 B.n356 VSUBS 0.006841f
C1239 B.n357 VSUBS 0.006841f
C1240 B.n358 VSUBS 0.006841f
C1241 B.n359 VSUBS 0.006841f
C1242 B.n360 VSUBS 0.006841f
C1243 B.n361 VSUBS 0.006841f
C1244 B.n362 VSUBS 0.006841f
C1245 B.n363 VSUBS 0.006841f
C1246 B.n364 VSUBS 0.006841f
C1247 B.n365 VSUBS 0.006841f
C1248 B.n366 VSUBS 0.006841f
C1249 B.n367 VSUBS 0.006841f
C1250 B.n368 VSUBS 0.006841f
C1251 B.n369 VSUBS 0.006841f
C1252 B.n370 VSUBS 0.006841f
C1253 B.n371 VSUBS 0.006841f
C1254 B.n372 VSUBS 0.006841f
C1255 B.n373 VSUBS 0.006841f
C1256 B.n374 VSUBS 0.006841f
C1257 B.n375 VSUBS 0.006841f
C1258 B.n376 VSUBS 0.006841f
C1259 B.n377 VSUBS 0.006841f
C1260 B.n378 VSUBS 0.006841f
C1261 B.n379 VSUBS 0.006841f
C1262 B.n380 VSUBS 0.006841f
C1263 B.n381 VSUBS 0.006841f
C1264 B.n382 VSUBS 0.006841f
C1265 B.n383 VSUBS 0.006841f
C1266 B.n384 VSUBS 0.006841f
C1267 B.n385 VSUBS 0.006841f
C1268 B.n386 VSUBS 0.006841f
C1269 B.n387 VSUBS 0.006841f
C1270 B.n388 VSUBS 0.006841f
C1271 B.n389 VSUBS 0.006841f
C1272 B.n390 VSUBS 0.006841f
C1273 B.n391 VSUBS 0.006841f
C1274 B.n392 VSUBS 0.006841f
C1275 B.n393 VSUBS 0.006841f
C1276 B.n394 VSUBS 0.006841f
C1277 B.n395 VSUBS 0.006841f
C1278 B.n396 VSUBS 0.006841f
C1279 B.n397 VSUBS 0.006841f
C1280 B.n398 VSUBS 0.006841f
C1281 B.n399 VSUBS 0.006841f
C1282 B.n400 VSUBS 0.006841f
C1283 B.n401 VSUBS 0.006841f
C1284 B.n402 VSUBS 0.006841f
C1285 B.n403 VSUBS 0.006841f
C1286 B.n404 VSUBS 0.006841f
C1287 B.n405 VSUBS 0.006841f
C1288 B.n406 VSUBS 0.006841f
C1289 B.n407 VSUBS 0.006841f
C1290 B.n408 VSUBS 0.006841f
C1291 B.n409 VSUBS 0.006841f
C1292 B.n410 VSUBS 0.006841f
C1293 B.n411 VSUBS 0.006841f
C1294 B.n412 VSUBS 0.006841f
C1295 B.n413 VSUBS 0.006841f
C1296 B.n414 VSUBS 0.006841f
C1297 B.n415 VSUBS 0.006841f
C1298 B.n416 VSUBS 0.006841f
C1299 B.n417 VSUBS 0.006841f
C1300 B.n418 VSUBS 0.006841f
C1301 B.n419 VSUBS 0.006841f
C1302 B.n420 VSUBS 0.006841f
C1303 B.n421 VSUBS 0.006841f
C1304 B.n422 VSUBS 0.006841f
C1305 B.n423 VSUBS 0.006841f
C1306 B.n424 VSUBS 0.006841f
C1307 B.n425 VSUBS 0.006841f
C1308 B.n426 VSUBS 0.006841f
C1309 B.n427 VSUBS 0.017067f
C1310 B.n428 VSUBS 0.017067f
C1311 B.n429 VSUBS 0.016535f
C1312 B.n430 VSUBS 0.006841f
C1313 B.n431 VSUBS 0.006841f
C1314 B.n432 VSUBS 0.006841f
C1315 B.n433 VSUBS 0.006841f
C1316 B.n434 VSUBS 0.006841f
C1317 B.n435 VSUBS 0.006841f
C1318 B.n436 VSUBS 0.006841f
C1319 B.n437 VSUBS 0.006841f
C1320 B.n438 VSUBS 0.006841f
C1321 B.n439 VSUBS 0.006841f
C1322 B.n440 VSUBS 0.006841f
C1323 B.n441 VSUBS 0.006841f
C1324 B.n442 VSUBS 0.006841f
C1325 B.n443 VSUBS 0.006841f
C1326 B.n444 VSUBS 0.006841f
C1327 B.n445 VSUBS 0.006841f
C1328 B.n446 VSUBS 0.006841f
C1329 B.n447 VSUBS 0.006841f
C1330 B.n448 VSUBS 0.006841f
C1331 B.n449 VSUBS 0.006841f
C1332 B.n450 VSUBS 0.006841f
C1333 B.n451 VSUBS 0.006841f
C1334 B.n452 VSUBS 0.006841f
C1335 B.n453 VSUBS 0.006841f
C1336 B.n454 VSUBS 0.006841f
C1337 B.n455 VSUBS 0.006841f
C1338 B.n456 VSUBS 0.006841f
C1339 B.n457 VSUBS 0.006841f
C1340 B.n458 VSUBS 0.006841f
C1341 B.n459 VSUBS 0.006841f
C1342 B.n460 VSUBS 0.006841f
C1343 B.n461 VSUBS 0.006841f
C1344 B.n462 VSUBS 0.006841f
C1345 B.n463 VSUBS 0.006841f
C1346 B.n464 VSUBS 0.006841f
C1347 B.n465 VSUBS 0.006841f
C1348 B.n466 VSUBS 0.006841f
C1349 B.n467 VSUBS 0.006841f
C1350 B.n468 VSUBS 0.006841f
C1351 B.n469 VSUBS 0.006841f
C1352 B.n470 VSUBS 0.006841f
C1353 B.n471 VSUBS 0.006841f
C1354 B.n472 VSUBS 0.006841f
C1355 B.n473 VSUBS 0.006841f
C1356 B.n474 VSUBS 0.006841f
C1357 B.n475 VSUBS 0.006841f
C1358 B.n476 VSUBS 0.006841f
C1359 B.n477 VSUBS 0.006841f
C1360 B.n478 VSUBS 0.006841f
C1361 B.n479 VSUBS 0.006841f
C1362 B.n480 VSUBS 0.006841f
C1363 B.n481 VSUBS 0.006841f
C1364 B.n482 VSUBS 0.006841f
C1365 B.n483 VSUBS 0.006841f
C1366 B.n484 VSUBS 0.006841f
C1367 B.n485 VSUBS 0.006841f
C1368 B.n486 VSUBS 0.006841f
C1369 B.n487 VSUBS 0.006841f
C1370 B.n488 VSUBS 0.006841f
C1371 B.n489 VSUBS 0.006841f
C1372 B.n490 VSUBS 0.006841f
C1373 B.n491 VSUBS 0.006841f
C1374 B.n492 VSUBS 0.006841f
C1375 B.n493 VSUBS 0.006841f
C1376 B.n494 VSUBS 0.006841f
C1377 B.n495 VSUBS 0.006841f
C1378 B.n496 VSUBS 0.006841f
C1379 B.n497 VSUBS 0.006841f
C1380 B.n498 VSUBS 0.006841f
C1381 B.n499 VSUBS 0.006841f
C1382 B.n500 VSUBS 0.006841f
C1383 B.n501 VSUBS 0.006841f
C1384 B.n502 VSUBS 0.006841f
C1385 B.n503 VSUBS 0.006841f
C1386 B.n504 VSUBS 0.017287f
C1387 B.n505 VSUBS 0.016315f
C1388 B.n506 VSUBS 0.017067f
C1389 B.n507 VSUBS 0.006841f
C1390 B.n508 VSUBS 0.006841f
C1391 B.n509 VSUBS 0.006841f
C1392 B.n510 VSUBS 0.006841f
C1393 B.n511 VSUBS 0.006841f
C1394 B.n512 VSUBS 0.006841f
C1395 B.n513 VSUBS 0.006841f
C1396 B.n514 VSUBS 0.006841f
C1397 B.n515 VSUBS 0.006841f
C1398 B.n516 VSUBS 0.006841f
C1399 B.n517 VSUBS 0.006841f
C1400 B.n518 VSUBS 0.006841f
C1401 B.n519 VSUBS 0.006841f
C1402 B.n520 VSUBS 0.006841f
C1403 B.n521 VSUBS 0.006841f
C1404 B.n522 VSUBS 0.006841f
C1405 B.n523 VSUBS 0.006841f
C1406 B.n524 VSUBS 0.006841f
C1407 B.n525 VSUBS 0.006841f
C1408 B.n526 VSUBS 0.006841f
C1409 B.n527 VSUBS 0.006841f
C1410 B.n528 VSUBS 0.006841f
C1411 B.n529 VSUBS 0.006841f
C1412 B.n530 VSUBS 0.006841f
C1413 B.n531 VSUBS 0.006841f
C1414 B.n532 VSUBS 0.006841f
C1415 B.n533 VSUBS 0.006841f
C1416 B.n534 VSUBS 0.006841f
C1417 B.n535 VSUBS 0.006841f
C1418 B.n536 VSUBS 0.006841f
C1419 B.n537 VSUBS 0.006841f
C1420 B.n538 VSUBS 0.006841f
C1421 B.n539 VSUBS 0.006841f
C1422 B.n540 VSUBS 0.006841f
C1423 B.n541 VSUBS 0.006841f
C1424 B.n542 VSUBS 0.006841f
C1425 B.n543 VSUBS 0.006841f
C1426 B.n544 VSUBS 0.006841f
C1427 B.n545 VSUBS 0.006841f
C1428 B.n546 VSUBS 0.006841f
C1429 B.n547 VSUBS 0.006841f
C1430 B.n548 VSUBS 0.006841f
C1431 B.n549 VSUBS 0.006841f
C1432 B.n550 VSUBS 0.006841f
C1433 B.n551 VSUBS 0.006841f
C1434 B.n552 VSUBS 0.006841f
C1435 B.n553 VSUBS 0.006841f
C1436 B.n554 VSUBS 0.006841f
C1437 B.n555 VSUBS 0.006841f
C1438 B.n556 VSUBS 0.006841f
C1439 B.n557 VSUBS 0.006841f
C1440 B.n558 VSUBS 0.006841f
C1441 B.n559 VSUBS 0.006841f
C1442 B.n560 VSUBS 0.006841f
C1443 B.n561 VSUBS 0.006841f
C1444 B.n562 VSUBS 0.006841f
C1445 B.n563 VSUBS 0.006841f
C1446 B.n564 VSUBS 0.006841f
C1447 B.n565 VSUBS 0.006841f
C1448 B.n566 VSUBS 0.006841f
C1449 B.n567 VSUBS 0.006841f
C1450 B.n568 VSUBS 0.006841f
C1451 B.n569 VSUBS 0.006841f
C1452 B.n570 VSUBS 0.006841f
C1453 B.n571 VSUBS 0.006841f
C1454 B.n572 VSUBS 0.006841f
C1455 B.n573 VSUBS 0.006841f
C1456 B.n574 VSUBS 0.006841f
C1457 B.n575 VSUBS 0.006841f
C1458 B.n576 VSUBS 0.006841f
C1459 B.n577 VSUBS 0.006841f
C1460 B.n578 VSUBS 0.006841f
C1461 B.n579 VSUBS 0.006841f
C1462 B.n580 VSUBS 0.006841f
C1463 B.n581 VSUBS 0.006841f
C1464 B.n582 VSUBS 0.006841f
C1465 B.n583 VSUBS 0.006841f
C1466 B.n584 VSUBS 0.006841f
C1467 B.n585 VSUBS 0.006841f
C1468 B.n586 VSUBS 0.006841f
C1469 B.n587 VSUBS 0.006841f
C1470 B.n588 VSUBS 0.006841f
C1471 B.n589 VSUBS 0.006841f
C1472 B.n590 VSUBS 0.006841f
C1473 B.n591 VSUBS 0.006841f
C1474 B.n592 VSUBS 0.006841f
C1475 B.n593 VSUBS 0.006841f
C1476 B.n594 VSUBS 0.006841f
C1477 B.n595 VSUBS 0.006439f
C1478 B.n596 VSUBS 0.006841f
C1479 B.n597 VSUBS 0.006841f
C1480 B.n598 VSUBS 0.003823f
C1481 B.n599 VSUBS 0.006841f
C1482 B.n600 VSUBS 0.006841f
C1483 B.n601 VSUBS 0.006841f
C1484 B.n602 VSUBS 0.006841f
C1485 B.n603 VSUBS 0.006841f
C1486 B.n604 VSUBS 0.006841f
C1487 B.n605 VSUBS 0.006841f
C1488 B.n606 VSUBS 0.006841f
C1489 B.n607 VSUBS 0.006841f
C1490 B.n608 VSUBS 0.006841f
C1491 B.n609 VSUBS 0.006841f
C1492 B.n610 VSUBS 0.006841f
C1493 B.n611 VSUBS 0.003823f
C1494 B.n612 VSUBS 0.01585f
C1495 B.n613 VSUBS 0.006439f
C1496 B.n614 VSUBS 0.006841f
C1497 B.n615 VSUBS 0.006841f
C1498 B.n616 VSUBS 0.006841f
C1499 B.n617 VSUBS 0.006841f
C1500 B.n618 VSUBS 0.006841f
C1501 B.n619 VSUBS 0.006841f
C1502 B.n620 VSUBS 0.006841f
C1503 B.n621 VSUBS 0.006841f
C1504 B.n622 VSUBS 0.006841f
C1505 B.n623 VSUBS 0.006841f
C1506 B.n624 VSUBS 0.006841f
C1507 B.n625 VSUBS 0.006841f
C1508 B.n626 VSUBS 0.006841f
C1509 B.n627 VSUBS 0.006841f
C1510 B.n628 VSUBS 0.006841f
C1511 B.n629 VSUBS 0.006841f
C1512 B.n630 VSUBS 0.006841f
C1513 B.n631 VSUBS 0.006841f
C1514 B.n632 VSUBS 0.006841f
C1515 B.n633 VSUBS 0.006841f
C1516 B.n634 VSUBS 0.006841f
C1517 B.n635 VSUBS 0.006841f
C1518 B.n636 VSUBS 0.006841f
C1519 B.n637 VSUBS 0.006841f
C1520 B.n638 VSUBS 0.006841f
C1521 B.n639 VSUBS 0.006841f
C1522 B.n640 VSUBS 0.006841f
C1523 B.n641 VSUBS 0.006841f
C1524 B.n642 VSUBS 0.006841f
C1525 B.n643 VSUBS 0.006841f
C1526 B.n644 VSUBS 0.006841f
C1527 B.n645 VSUBS 0.006841f
C1528 B.n646 VSUBS 0.006841f
C1529 B.n647 VSUBS 0.006841f
C1530 B.n648 VSUBS 0.006841f
C1531 B.n649 VSUBS 0.006841f
C1532 B.n650 VSUBS 0.006841f
C1533 B.n651 VSUBS 0.006841f
C1534 B.n652 VSUBS 0.006841f
C1535 B.n653 VSUBS 0.006841f
C1536 B.n654 VSUBS 0.006841f
C1537 B.n655 VSUBS 0.006841f
C1538 B.n656 VSUBS 0.006841f
C1539 B.n657 VSUBS 0.006841f
C1540 B.n658 VSUBS 0.006841f
C1541 B.n659 VSUBS 0.006841f
C1542 B.n660 VSUBS 0.006841f
C1543 B.n661 VSUBS 0.006841f
C1544 B.n662 VSUBS 0.006841f
C1545 B.n663 VSUBS 0.006841f
C1546 B.n664 VSUBS 0.006841f
C1547 B.n665 VSUBS 0.006841f
C1548 B.n666 VSUBS 0.006841f
C1549 B.n667 VSUBS 0.006841f
C1550 B.n668 VSUBS 0.006841f
C1551 B.n669 VSUBS 0.006841f
C1552 B.n670 VSUBS 0.006841f
C1553 B.n671 VSUBS 0.006841f
C1554 B.n672 VSUBS 0.006841f
C1555 B.n673 VSUBS 0.006841f
C1556 B.n674 VSUBS 0.006841f
C1557 B.n675 VSUBS 0.006841f
C1558 B.n676 VSUBS 0.006841f
C1559 B.n677 VSUBS 0.006841f
C1560 B.n678 VSUBS 0.006841f
C1561 B.n679 VSUBS 0.006841f
C1562 B.n680 VSUBS 0.006841f
C1563 B.n681 VSUBS 0.006841f
C1564 B.n682 VSUBS 0.006841f
C1565 B.n683 VSUBS 0.006841f
C1566 B.n684 VSUBS 0.006841f
C1567 B.n685 VSUBS 0.006841f
C1568 B.n686 VSUBS 0.006841f
C1569 B.n687 VSUBS 0.006841f
C1570 B.n688 VSUBS 0.006841f
C1571 B.n689 VSUBS 0.006841f
C1572 B.n690 VSUBS 0.006841f
C1573 B.n691 VSUBS 0.006841f
C1574 B.n692 VSUBS 0.006841f
C1575 B.n693 VSUBS 0.006841f
C1576 B.n694 VSUBS 0.006841f
C1577 B.n695 VSUBS 0.006841f
C1578 B.n696 VSUBS 0.006841f
C1579 B.n697 VSUBS 0.006841f
C1580 B.n698 VSUBS 0.006841f
C1581 B.n699 VSUBS 0.006841f
C1582 B.n700 VSUBS 0.006841f
C1583 B.n701 VSUBS 0.006841f
C1584 B.n702 VSUBS 0.006841f
C1585 B.n703 VSUBS 0.017067f
C1586 B.n704 VSUBS 0.017067f
C1587 B.n705 VSUBS 0.016535f
C1588 B.n706 VSUBS 0.006841f
C1589 B.n707 VSUBS 0.006841f
C1590 B.n708 VSUBS 0.006841f
C1591 B.n709 VSUBS 0.006841f
C1592 B.n710 VSUBS 0.006841f
C1593 B.n711 VSUBS 0.006841f
C1594 B.n712 VSUBS 0.006841f
C1595 B.n713 VSUBS 0.006841f
C1596 B.n714 VSUBS 0.006841f
C1597 B.n715 VSUBS 0.006841f
C1598 B.n716 VSUBS 0.006841f
C1599 B.n717 VSUBS 0.006841f
C1600 B.n718 VSUBS 0.006841f
C1601 B.n719 VSUBS 0.006841f
C1602 B.n720 VSUBS 0.006841f
C1603 B.n721 VSUBS 0.006841f
C1604 B.n722 VSUBS 0.006841f
C1605 B.n723 VSUBS 0.006841f
C1606 B.n724 VSUBS 0.006841f
C1607 B.n725 VSUBS 0.006841f
C1608 B.n726 VSUBS 0.006841f
C1609 B.n727 VSUBS 0.006841f
C1610 B.n728 VSUBS 0.006841f
C1611 B.n729 VSUBS 0.006841f
C1612 B.n730 VSUBS 0.006841f
C1613 B.n731 VSUBS 0.006841f
C1614 B.n732 VSUBS 0.006841f
C1615 B.n733 VSUBS 0.006841f
C1616 B.n734 VSUBS 0.006841f
C1617 B.n735 VSUBS 0.006841f
C1618 B.n736 VSUBS 0.006841f
C1619 B.n737 VSUBS 0.006841f
C1620 B.n738 VSUBS 0.006841f
C1621 B.n739 VSUBS 0.006841f
C1622 B.n740 VSUBS 0.006841f
C1623 B.n741 VSUBS 0.006841f
C1624 B.n742 VSUBS 0.006841f
C1625 B.n743 VSUBS 0.015491f
.ends

