* NGSPICE file created from diff_pair_sample_0439.ext - technology: sky130A

.subckt diff_pair_sample_0439 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0.98175 ps=6.28 w=5.95 l=3.75
X1 B.t11 B.t9 B.t10 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0 ps=0 w=5.95 l=3.75
X2 VDD2.t2 VN.t1 VTAIL.t6 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=0.98175 pd=6.28 as=2.3205 ps=12.68 w=5.95 l=3.75
X3 B.t8 B.t6 B.t7 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0 ps=0 w=5.95 l=3.75
X4 VDD1.t3 VP.t0 VTAIL.t3 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=0.98175 pd=6.28 as=2.3205 ps=12.68 w=5.95 l=3.75
X5 B.t5 B.t3 B.t4 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0 ps=0 w=5.95 l=3.75
X6 VDD2.t3 VN.t2 VTAIL.t5 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=0.98175 pd=6.28 as=2.3205 ps=12.68 w=5.95 l=3.75
X7 VDD1.t2 VP.t1 VTAIL.t0 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=0.98175 pd=6.28 as=2.3205 ps=12.68 w=5.95 l=3.75
X8 VTAIL.t4 VN.t3 VDD2.t1 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0.98175 ps=6.28 w=5.95 l=3.75
X9 B.t2 B.t0 B.t1 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0 ps=0 w=5.95 l=3.75
X10 VTAIL.t1 VP.t2 VDD1.t1 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0.98175 ps=6.28 w=5.95 l=3.75
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n3418_n2158# sky130_fd_pr__pfet_01v8 ad=2.3205 pd=12.68 as=0.98175 ps=6.28 w=5.95 l=3.75
R0 VN.n0 VN.t0 71.8585
R1 VN.n1 VN.t1 71.8585
R2 VN.n0 VN.t2 70.5207
R3 VN.n1 VN.t3 70.5207
R4 VN VN.n1 47.3321
R5 VN VN.n0 1.89646
R6 VDD2.n2 VDD2.n0 130.72
R7 VDD2.n2 VDD2.n1 91.3244
R8 VDD2.n1 VDD2.t1 5.46353
R9 VDD2.n1 VDD2.t2 5.46353
R10 VDD2.n0 VDD2.t0 5.46353
R11 VDD2.n0 VDD2.t3 5.46353
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n250 VTAIL.n224 756.745
R14 VTAIL.n26 VTAIL.n0 756.745
R15 VTAIL.n58 VTAIL.n32 756.745
R16 VTAIL.n90 VTAIL.n64 756.745
R17 VTAIL.n218 VTAIL.n192 756.745
R18 VTAIL.n186 VTAIL.n160 756.745
R19 VTAIL.n154 VTAIL.n128 756.745
R20 VTAIL.n122 VTAIL.n96 756.745
R21 VTAIL.n235 VTAIL.n234 585
R22 VTAIL.n232 VTAIL.n231 585
R23 VTAIL.n241 VTAIL.n240 585
R24 VTAIL.n243 VTAIL.n242 585
R25 VTAIL.n228 VTAIL.n227 585
R26 VTAIL.n249 VTAIL.n248 585
R27 VTAIL.n251 VTAIL.n250 585
R28 VTAIL.n11 VTAIL.n10 585
R29 VTAIL.n8 VTAIL.n7 585
R30 VTAIL.n17 VTAIL.n16 585
R31 VTAIL.n19 VTAIL.n18 585
R32 VTAIL.n4 VTAIL.n3 585
R33 VTAIL.n25 VTAIL.n24 585
R34 VTAIL.n27 VTAIL.n26 585
R35 VTAIL.n43 VTAIL.n42 585
R36 VTAIL.n40 VTAIL.n39 585
R37 VTAIL.n49 VTAIL.n48 585
R38 VTAIL.n51 VTAIL.n50 585
R39 VTAIL.n36 VTAIL.n35 585
R40 VTAIL.n57 VTAIL.n56 585
R41 VTAIL.n59 VTAIL.n58 585
R42 VTAIL.n75 VTAIL.n74 585
R43 VTAIL.n72 VTAIL.n71 585
R44 VTAIL.n81 VTAIL.n80 585
R45 VTAIL.n83 VTAIL.n82 585
R46 VTAIL.n68 VTAIL.n67 585
R47 VTAIL.n89 VTAIL.n88 585
R48 VTAIL.n91 VTAIL.n90 585
R49 VTAIL.n219 VTAIL.n218 585
R50 VTAIL.n217 VTAIL.n216 585
R51 VTAIL.n196 VTAIL.n195 585
R52 VTAIL.n211 VTAIL.n210 585
R53 VTAIL.n209 VTAIL.n208 585
R54 VTAIL.n200 VTAIL.n199 585
R55 VTAIL.n203 VTAIL.n202 585
R56 VTAIL.n187 VTAIL.n186 585
R57 VTAIL.n185 VTAIL.n184 585
R58 VTAIL.n164 VTAIL.n163 585
R59 VTAIL.n179 VTAIL.n178 585
R60 VTAIL.n177 VTAIL.n176 585
R61 VTAIL.n168 VTAIL.n167 585
R62 VTAIL.n171 VTAIL.n170 585
R63 VTAIL.n155 VTAIL.n154 585
R64 VTAIL.n153 VTAIL.n152 585
R65 VTAIL.n132 VTAIL.n131 585
R66 VTAIL.n147 VTAIL.n146 585
R67 VTAIL.n145 VTAIL.n144 585
R68 VTAIL.n136 VTAIL.n135 585
R69 VTAIL.n139 VTAIL.n138 585
R70 VTAIL.n123 VTAIL.n122 585
R71 VTAIL.n121 VTAIL.n120 585
R72 VTAIL.n100 VTAIL.n99 585
R73 VTAIL.n115 VTAIL.n114 585
R74 VTAIL.n113 VTAIL.n112 585
R75 VTAIL.n104 VTAIL.n103 585
R76 VTAIL.n107 VTAIL.n106 585
R77 VTAIL.t5 VTAIL.n233 327.601
R78 VTAIL.t7 VTAIL.n9 327.601
R79 VTAIL.t0 VTAIL.n41 327.601
R80 VTAIL.t1 VTAIL.n73 327.601
R81 VTAIL.t3 VTAIL.n201 327.601
R82 VTAIL.t2 VTAIL.n169 327.601
R83 VTAIL.t6 VTAIL.n137 327.601
R84 VTAIL.t4 VTAIL.n105 327.601
R85 VTAIL.n234 VTAIL.n231 171.744
R86 VTAIL.n241 VTAIL.n231 171.744
R87 VTAIL.n242 VTAIL.n241 171.744
R88 VTAIL.n242 VTAIL.n227 171.744
R89 VTAIL.n249 VTAIL.n227 171.744
R90 VTAIL.n250 VTAIL.n249 171.744
R91 VTAIL.n10 VTAIL.n7 171.744
R92 VTAIL.n17 VTAIL.n7 171.744
R93 VTAIL.n18 VTAIL.n17 171.744
R94 VTAIL.n18 VTAIL.n3 171.744
R95 VTAIL.n25 VTAIL.n3 171.744
R96 VTAIL.n26 VTAIL.n25 171.744
R97 VTAIL.n42 VTAIL.n39 171.744
R98 VTAIL.n49 VTAIL.n39 171.744
R99 VTAIL.n50 VTAIL.n49 171.744
R100 VTAIL.n50 VTAIL.n35 171.744
R101 VTAIL.n57 VTAIL.n35 171.744
R102 VTAIL.n58 VTAIL.n57 171.744
R103 VTAIL.n74 VTAIL.n71 171.744
R104 VTAIL.n81 VTAIL.n71 171.744
R105 VTAIL.n82 VTAIL.n81 171.744
R106 VTAIL.n82 VTAIL.n67 171.744
R107 VTAIL.n89 VTAIL.n67 171.744
R108 VTAIL.n90 VTAIL.n89 171.744
R109 VTAIL.n218 VTAIL.n217 171.744
R110 VTAIL.n217 VTAIL.n195 171.744
R111 VTAIL.n210 VTAIL.n195 171.744
R112 VTAIL.n210 VTAIL.n209 171.744
R113 VTAIL.n209 VTAIL.n199 171.744
R114 VTAIL.n202 VTAIL.n199 171.744
R115 VTAIL.n186 VTAIL.n185 171.744
R116 VTAIL.n185 VTAIL.n163 171.744
R117 VTAIL.n178 VTAIL.n163 171.744
R118 VTAIL.n178 VTAIL.n177 171.744
R119 VTAIL.n177 VTAIL.n167 171.744
R120 VTAIL.n170 VTAIL.n167 171.744
R121 VTAIL.n154 VTAIL.n153 171.744
R122 VTAIL.n153 VTAIL.n131 171.744
R123 VTAIL.n146 VTAIL.n131 171.744
R124 VTAIL.n146 VTAIL.n145 171.744
R125 VTAIL.n145 VTAIL.n135 171.744
R126 VTAIL.n138 VTAIL.n135 171.744
R127 VTAIL.n122 VTAIL.n121 171.744
R128 VTAIL.n121 VTAIL.n99 171.744
R129 VTAIL.n114 VTAIL.n99 171.744
R130 VTAIL.n114 VTAIL.n113 171.744
R131 VTAIL.n113 VTAIL.n103 171.744
R132 VTAIL.n106 VTAIL.n103 171.744
R133 VTAIL.n234 VTAIL.t5 85.8723
R134 VTAIL.n10 VTAIL.t7 85.8723
R135 VTAIL.n42 VTAIL.t0 85.8723
R136 VTAIL.n74 VTAIL.t1 85.8723
R137 VTAIL.n202 VTAIL.t3 85.8723
R138 VTAIL.n170 VTAIL.t2 85.8723
R139 VTAIL.n138 VTAIL.t6 85.8723
R140 VTAIL.n106 VTAIL.t4 85.8723
R141 VTAIL.n255 VTAIL.n254 31.2157
R142 VTAIL.n31 VTAIL.n30 31.2157
R143 VTAIL.n63 VTAIL.n62 31.2157
R144 VTAIL.n95 VTAIL.n94 31.2157
R145 VTAIL.n223 VTAIL.n222 31.2157
R146 VTAIL.n191 VTAIL.n190 31.2157
R147 VTAIL.n159 VTAIL.n158 31.2157
R148 VTAIL.n127 VTAIL.n126 31.2157
R149 VTAIL.n255 VTAIL.n223 21.0134
R150 VTAIL.n127 VTAIL.n95 21.0134
R151 VTAIL.n235 VTAIL.n233 16.3865
R152 VTAIL.n11 VTAIL.n9 16.3865
R153 VTAIL.n43 VTAIL.n41 16.3865
R154 VTAIL.n75 VTAIL.n73 16.3865
R155 VTAIL.n203 VTAIL.n201 16.3865
R156 VTAIL.n171 VTAIL.n169 16.3865
R157 VTAIL.n139 VTAIL.n137 16.3865
R158 VTAIL.n107 VTAIL.n105 16.3865
R159 VTAIL.n236 VTAIL.n232 12.8005
R160 VTAIL.n12 VTAIL.n8 12.8005
R161 VTAIL.n44 VTAIL.n40 12.8005
R162 VTAIL.n76 VTAIL.n72 12.8005
R163 VTAIL.n204 VTAIL.n200 12.8005
R164 VTAIL.n172 VTAIL.n168 12.8005
R165 VTAIL.n140 VTAIL.n136 12.8005
R166 VTAIL.n108 VTAIL.n104 12.8005
R167 VTAIL.n240 VTAIL.n239 12.0247
R168 VTAIL.n16 VTAIL.n15 12.0247
R169 VTAIL.n48 VTAIL.n47 12.0247
R170 VTAIL.n80 VTAIL.n79 12.0247
R171 VTAIL.n208 VTAIL.n207 12.0247
R172 VTAIL.n176 VTAIL.n175 12.0247
R173 VTAIL.n144 VTAIL.n143 12.0247
R174 VTAIL.n112 VTAIL.n111 12.0247
R175 VTAIL.n243 VTAIL.n230 11.249
R176 VTAIL.n19 VTAIL.n6 11.249
R177 VTAIL.n51 VTAIL.n38 11.249
R178 VTAIL.n83 VTAIL.n70 11.249
R179 VTAIL.n211 VTAIL.n198 11.249
R180 VTAIL.n179 VTAIL.n166 11.249
R181 VTAIL.n147 VTAIL.n134 11.249
R182 VTAIL.n115 VTAIL.n102 11.249
R183 VTAIL.n244 VTAIL.n228 10.4732
R184 VTAIL.n20 VTAIL.n4 10.4732
R185 VTAIL.n52 VTAIL.n36 10.4732
R186 VTAIL.n84 VTAIL.n68 10.4732
R187 VTAIL.n212 VTAIL.n196 10.4732
R188 VTAIL.n180 VTAIL.n164 10.4732
R189 VTAIL.n148 VTAIL.n132 10.4732
R190 VTAIL.n116 VTAIL.n100 10.4732
R191 VTAIL.n248 VTAIL.n247 9.69747
R192 VTAIL.n24 VTAIL.n23 9.69747
R193 VTAIL.n56 VTAIL.n55 9.69747
R194 VTAIL.n88 VTAIL.n87 9.69747
R195 VTAIL.n216 VTAIL.n215 9.69747
R196 VTAIL.n184 VTAIL.n183 9.69747
R197 VTAIL.n152 VTAIL.n151 9.69747
R198 VTAIL.n120 VTAIL.n119 9.69747
R199 VTAIL.n254 VTAIL.n253 9.45567
R200 VTAIL.n30 VTAIL.n29 9.45567
R201 VTAIL.n62 VTAIL.n61 9.45567
R202 VTAIL.n94 VTAIL.n93 9.45567
R203 VTAIL.n222 VTAIL.n221 9.45567
R204 VTAIL.n190 VTAIL.n189 9.45567
R205 VTAIL.n158 VTAIL.n157 9.45567
R206 VTAIL.n126 VTAIL.n125 9.45567
R207 VTAIL.n253 VTAIL.n252 9.3005
R208 VTAIL.n226 VTAIL.n225 9.3005
R209 VTAIL.n247 VTAIL.n246 9.3005
R210 VTAIL.n245 VTAIL.n244 9.3005
R211 VTAIL.n230 VTAIL.n229 9.3005
R212 VTAIL.n239 VTAIL.n238 9.3005
R213 VTAIL.n237 VTAIL.n236 9.3005
R214 VTAIL.n29 VTAIL.n28 9.3005
R215 VTAIL.n2 VTAIL.n1 9.3005
R216 VTAIL.n23 VTAIL.n22 9.3005
R217 VTAIL.n21 VTAIL.n20 9.3005
R218 VTAIL.n6 VTAIL.n5 9.3005
R219 VTAIL.n15 VTAIL.n14 9.3005
R220 VTAIL.n13 VTAIL.n12 9.3005
R221 VTAIL.n61 VTAIL.n60 9.3005
R222 VTAIL.n34 VTAIL.n33 9.3005
R223 VTAIL.n55 VTAIL.n54 9.3005
R224 VTAIL.n53 VTAIL.n52 9.3005
R225 VTAIL.n38 VTAIL.n37 9.3005
R226 VTAIL.n47 VTAIL.n46 9.3005
R227 VTAIL.n45 VTAIL.n44 9.3005
R228 VTAIL.n93 VTAIL.n92 9.3005
R229 VTAIL.n66 VTAIL.n65 9.3005
R230 VTAIL.n87 VTAIL.n86 9.3005
R231 VTAIL.n85 VTAIL.n84 9.3005
R232 VTAIL.n70 VTAIL.n69 9.3005
R233 VTAIL.n79 VTAIL.n78 9.3005
R234 VTAIL.n77 VTAIL.n76 9.3005
R235 VTAIL.n221 VTAIL.n220 9.3005
R236 VTAIL.n194 VTAIL.n193 9.3005
R237 VTAIL.n215 VTAIL.n214 9.3005
R238 VTAIL.n213 VTAIL.n212 9.3005
R239 VTAIL.n198 VTAIL.n197 9.3005
R240 VTAIL.n207 VTAIL.n206 9.3005
R241 VTAIL.n205 VTAIL.n204 9.3005
R242 VTAIL.n189 VTAIL.n188 9.3005
R243 VTAIL.n162 VTAIL.n161 9.3005
R244 VTAIL.n183 VTAIL.n182 9.3005
R245 VTAIL.n181 VTAIL.n180 9.3005
R246 VTAIL.n166 VTAIL.n165 9.3005
R247 VTAIL.n175 VTAIL.n174 9.3005
R248 VTAIL.n173 VTAIL.n172 9.3005
R249 VTAIL.n157 VTAIL.n156 9.3005
R250 VTAIL.n130 VTAIL.n129 9.3005
R251 VTAIL.n151 VTAIL.n150 9.3005
R252 VTAIL.n149 VTAIL.n148 9.3005
R253 VTAIL.n134 VTAIL.n133 9.3005
R254 VTAIL.n143 VTAIL.n142 9.3005
R255 VTAIL.n141 VTAIL.n140 9.3005
R256 VTAIL.n125 VTAIL.n124 9.3005
R257 VTAIL.n98 VTAIL.n97 9.3005
R258 VTAIL.n119 VTAIL.n118 9.3005
R259 VTAIL.n117 VTAIL.n116 9.3005
R260 VTAIL.n102 VTAIL.n101 9.3005
R261 VTAIL.n111 VTAIL.n110 9.3005
R262 VTAIL.n109 VTAIL.n108 9.3005
R263 VTAIL.n251 VTAIL.n226 8.92171
R264 VTAIL.n27 VTAIL.n2 8.92171
R265 VTAIL.n59 VTAIL.n34 8.92171
R266 VTAIL.n91 VTAIL.n66 8.92171
R267 VTAIL.n219 VTAIL.n194 8.92171
R268 VTAIL.n187 VTAIL.n162 8.92171
R269 VTAIL.n155 VTAIL.n130 8.92171
R270 VTAIL.n123 VTAIL.n98 8.92171
R271 VTAIL.n252 VTAIL.n224 8.14595
R272 VTAIL.n28 VTAIL.n0 8.14595
R273 VTAIL.n60 VTAIL.n32 8.14595
R274 VTAIL.n92 VTAIL.n64 8.14595
R275 VTAIL.n220 VTAIL.n192 8.14595
R276 VTAIL.n188 VTAIL.n160 8.14595
R277 VTAIL.n156 VTAIL.n128 8.14595
R278 VTAIL.n124 VTAIL.n96 8.14595
R279 VTAIL.n254 VTAIL.n224 5.81868
R280 VTAIL.n30 VTAIL.n0 5.81868
R281 VTAIL.n62 VTAIL.n32 5.81868
R282 VTAIL.n94 VTAIL.n64 5.81868
R283 VTAIL.n222 VTAIL.n192 5.81868
R284 VTAIL.n190 VTAIL.n160 5.81868
R285 VTAIL.n158 VTAIL.n128 5.81868
R286 VTAIL.n126 VTAIL.n96 5.81868
R287 VTAIL.n252 VTAIL.n251 5.04292
R288 VTAIL.n28 VTAIL.n27 5.04292
R289 VTAIL.n60 VTAIL.n59 5.04292
R290 VTAIL.n92 VTAIL.n91 5.04292
R291 VTAIL.n220 VTAIL.n219 5.04292
R292 VTAIL.n188 VTAIL.n187 5.04292
R293 VTAIL.n156 VTAIL.n155 5.04292
R294 VTAIL.n124 VTAIL.n123 5.04292
R295 VTAIL.n248 VTAIL.n226 4.26717
R296 VTAIL.n24 VTAIL.n2 4.26717
R297 VTAIL.n56 VTAIL.n34 4.26717
R298 VTAIL.n88 VTAIL.n66 4.26717
R299 VTAIL.n216 VTAIL.n194 4.26717
R300 VTAIL.n184 VTAIL.n162 4.26717
R301 VTAIL.n152 VTAIL.n130 4.26717
R302 VTAIL.n120 VTAIL.n98 4.26717
R303 VTAIL.n205 VTAIL.n201 3.71286
R304 VTAIL.n173 VTAIL.n169 3.71286
R305 VTAIL.n141 VTAIL.n137 3.71286
R306 VTAIL.n109 VTAIL.n105 3.71286
R307 VTAIL.n237 VTAIL.n233 3.71286
R308 VTAIL.n13 VTAIL.n9 3.71286
R309 VTAIL.n45 VTAIL.n41 3.71286
R310 VTAIL.n77 VTAIL.n73 3.71286
R311 VTAIL.n159 VTAIL.n127 3.51774
R312 VTAIL.n223 VTAIL.n191 3.51774
R313 VTAIL.n95 VTAIL.n63 3.51774
R314 VTAIL.n247 VTAIL.n228 3.49141
R315 VTAIL.n23 VTAIL.n4 3.49141
R316 VTAIL.n55 VTAIL.n36 3.49141
R317 VTAIL.n87 VTAIL.n68 3.49141
R318 VTAIL.n215 VTAIL.n196 3.49141
R319 VTAIL.n183 VTAIL.n164 3.49141
R320 VTAIL.n151 VTAIL.n132 3.49141
R321 VTAIL.n119 VTAIL.n100 3.49141
R322 VTAIL.n244 VTAIL.n243 2.71565
R323 VTAIL.n20 VTAIL.n19 2.71565
R324 VTAIL.n52 VTAIL.n51 2.71565
R325 VTAIL.n84 VTAIL.n83 2.71565
R326 VTAIL.n212 VTAIL.n211 2.71565
R327 VTAIL.n180 VTAIL.n179 2.71565
R328 VTAIL.n148 VTAIL.n147 2.71565
R329 VTAIL.n116 VTAIL.n115 2.71565
R330 VTAIL.n240 VTAIL.n230 1.93989
R331 VTAIL.n16 VTAIL.n6 1.93989
R332 VTAIL.n48 VTAIL.n38 1.93989
R333 VTAIL.n80 VTAIL.n70 1.93989
R334 VTAIL.n208 VTAIL.n198 1.93989
R335 VTAIL.n176 VTAIL.n166 1.93989
R336 VTAIL.n144 VTAIL.n134 1.93989
R337 VTAIL.n112 VTAIL.n102 1.93989
R338 VTAIL VTAIL.n31 1.81731
R339 VTAIL VTAIL.n255 1.70093
R340 VTAIL.n239 VTAIL.n232 1.16414
R341 VTAIL.n15 VTAIL.n8 1.16414
R342 VTAIL.n47 VTAIL.n40 1.16414
R343 VTAIL.n79 VTAIL.n72 1.16414
R344 VTAIL.n207 VTAIL.n200 1.16414
R345 VTAIL.n175 VTAIL.n168 1.16414
R346 VTAIL.n143 VTAIL.n136 1.16414
R347 VTAIL.n111 VTAIL.n104 1.16414
R348 VTAIL.n191 VTAIL.n159 0.470328
R349 VTAIL.n63 VTAIL.n31 0.470328
R350 VTAIL.n236 VTAIL.n235 0.388379
R351 VTAIL.n12 VTAIL.n11 0.388379
R352 VTAIL.n44 VTAIL.n43 0.388379
R353 VTAIL.n76 VTAIL.n75 0.388379
R354 VTAIL.n204 VTAIL.n203 0.388379
R355 VTAIL.n172 VTAIL.n171 0.388379
R356 VTAIL.n140 VTAIL.n139 0.388379
R357 VTAIL.n108 VTAIL.n107 0.388379
R358 VTAIL.n238 VTAIL.n237 0.155672
R359 VTAIL.n238 VTAIL.n229 0.155672
R360 VTAIL.n245 VTAIL.n229 0.155672
R361 VTAIL.n246 VTAIL.n245 0.155672
R362 VTAIL.n246 VTAIL.n225 0.155672
R363 VTAIL.n253 VTAIL.n225 0.155672
R364 VTAIL.n14 VTAIL.n13 0.155672
R365 VTAIL.n14 VTAIL.n5 0.155672
R366 VTAIL.n21 VTAIL.n5 0.155672
R367 VTAIL.n22 VTAIL.n21 0.155672
R368 VTAIL.n22 VTAIL.n1 0.155672
R369 VTAIL.n29 VTAIL.n1 0.155672
R370 VTAIL.n46 VTAIL.n45 0.155672
R371 VTAIL.n46 VTAIL.n37 0.155672
R372 VTAIL.n53 VTAIL.n37 0.155672
R373 VTAIL.n54 VTAIL.n53 0.155672
R374 VTAIL.n54 VTAIL.n33 0.155672
R375 VTAIL.n61 VTAIL.n33 0.155672
R376 VTAIL.n78 VTAIL.n77 0.155672
R377 VTAIL.n78 VTAIL.n69 0.155672
R378 VTAIL.n85 VTAIL.n69 0.155672
R379 VTAIL.n86 VTAIL.n85 0.155672
R380 VTAIL.n86 VTAIL.n65 0.155672
R381 VTAIL.n93 VTAIL.n65 0.155672
R382 VTAIL.n221 VTAIL.n193 0.155672
R383 VTAIL.n214 VTAIL.n193 0.155672
R384 VTAIL.n214 VTAIL.n213 0.155672
R385 VTAIL.n213 VTAIL.n197 0.155672
R386 VTAIL.n206 VTAIL.n197 0.155672
R387 VTAIL.n206 VTAIL.n205 0.155672
R388 VTAIL.n189 VTAIL.n161 0.155672
R389 VTAIL.n182 VTAIL.n161 0.155672
R390 VTAIL.n182 VTAIL.n181 0.155672
R391 VTAIL.n181 VTAIL.n165 0.155672
R392 VTAIL.n174 VTAIL.n165 0.155672
R393 VTAIL.n174 VTAIL.n173 0.155672
R394 VTAIL.n157 VTAIL.n129 0.155672
R395 VTAIL.n150 VTAIL.n129 0.155672
R396 VTAIL.n150 VTAIL.n149 0.155672
R397 VTAIL.n149 VTAIL.n133 0.155672
R398 VTAIL.n142 VTAIL.n133 0.155672
R399 VTAIL.n142 VTAIL.n141 0.155672
R400 VTAIL.n125 VTAIL.n97 0.155672
R401 VTAIL.n118 VTAIL.n97 0.155672
R402 VTAIL.n118 VTAIL.n117 0.155672
R403 VTAIL.n117 VTAIL.n101 0.155672
R404 VTAIL.n110 VTAIL.n101 0.155672
R405 VTAIL.n110 VTAIL.n109 0.155672
R406 B.n442 B.n441 585
R407 B.n443 B.n56 585
R408 B.n445 B.n444 585
R409 B.n446 B.n55 585
R410 B.n448 B.n447 585
R411 B.n449 B.n54 585
R412 B.n451 B.n450 585
R413 B.n452 B.n53 585
R414 B.n454 B.n453 585
R415 B.n455 B.n52 585
R416 B.n457 B.n456 585
R417 B.n458 B.n51 585
R418 B.n460 B.n459 585
R419 B.n461 B.n50 585
R420 B.n463 B.n462 585
R421 B.n464 B.n49 585
R422 B.n466 B.n465 585
R423 B.n467 B.n48 585
R424 B.n469 B.n468 585
R425 B.n470 B.n47 585
R426 B.n472 B.n471 585
R427 B.n473 B.n46 585
R428 B.n475 B.n474 585
R429 B.n476 B.n43 585
R430 B.n479 B.n478 585
R431 B.n480 B.n42 585
R432 B.n482 B.n481 585
R433 B.n483 B.n41 585
R434 B.n485 B.n484 585
R435 B.n486 B.n40 585
R436 B.n488 B.n487 585
R437 B.n489 B.n39 585
R438 B.n491 B.n490 585
R439 B.n493 B.n492 585
R440 B.n494 B.n35 585
R441 B.n496 B.n495 585
R442 B.n497 B.n34 585
R443 B.n499 B.n498 585
R444 B.n500 B.n33 585
R445 B.n502 B.n501 585
R446 B.n503 B.n32 585
R447 B.n505 B.n504 585
R448 B.n506 B.n31 585
R449 B.n508 B.n507 585
R450 B.n509 B.n30 585
R451 B.n511 B.n510 585
R452 B.n512 B.n29 585
R453 B.n514 B.n513 585
R454 B.n515 B.n28 585
R455 B.n517 B.n516 585
R456 B.n518 B.n27 585
R457 B.n520 B.n519 585
R458 B.n521 B.n26 585
R459 B.n523 B.n522 585
R460 B.n524 B.n25 585
R461 B.n526 B.n525 585
R462 B.n527 B.n24 585
R463 B.n440 B.n57 585
R464 B.n439 B.n438 585
R465 B.n437 B.n58 585
R466 B.n436 B.n435 585
R467 B.n434 B.n59 585
R468 B.n433 B.n432 585
R469 B.n431 B.n60 585
R470 B.n430 B.n429 585
R471 B.n428 B.n61 585
R472 B.n427 B.n426 585
R473 B.n425 B.n62 585
R474 B.n424 B.n423 585
R475 B.n422 B.n63 585
R476 B.n421 B.n420 585
R477 B.n419 B.n64 585
R478 B.n418 B.n417 585
R479 B.n416 B.n65 585
R480 B.n415 B.n414 585
R481 B.n413 B.n66 585
R482 B.n412 B.n411 585
R483 B.n410 B.n67 585
R484 B.n409 B.n408 585
R485 B.n407 B.n68 585
R486 B.n406 B.n405 585
R487 B.n404 B.n69 585
R488 B.n403 B.n402 585
R489 B.n401 B.n70 585
R490 B.n400 B.n399 585
R491 B.n398 B.n71 585
R492 B.n397 B.n396 585
R493 B.n395 B.n72 585
R494 B.n394 B.n393 585
R495 B.n392 B.n73 585
R496 B.n391 B.n390 585
R497 B.n389 B.n74 585
R498 B.n388 B.n387 585
R499 B.n386 B.n75 585
R500 B.n385 B.n384 585
R501 B.n383 B.n76 585
R502 B.n382 B.n381 585
R503 B.n380 B.n77 585
R504 B.n379 B.n378 585
R505 B.n377 B.n78 585
R506 B.n376 B.n375 585
R507 B.n374 B.n79 585
R508 B.n373 B.n372 585
R509 B.n371 B.n80 585
R510 B.n370 B.n369 585
R511 B.n368 B.n81 585
R512 B.n367 B.n366 585
R513 B.n365 B.n82 585
R514 B.n364 B.n363 585
R515 B.n362 B.n83 585
R516 B.n361 B.n360 585
R517 B.n359 B.n84 585
R518 B.n358 B.n357 585
R519 B.n356 B.n85 585
R520 B.n355 B.n354 585
R521 B.n353 B.n86 585
R522 B.n352 B.n351 585
R523 B.n350 B.n87 585
R524 B.n349 B.n348 585
R525 B.n347 B.n88 585
R526 B.n346 B.n345 585
R527 B.n344 B.n89 585
R528 B.n343 B.n342 585
R529 B.n341 B.n90 585
R530 B.n340 B.n339 585
R531 B.n338 B.n91 585
R532 B.n337 B.n336 585
R533 B.n335 B.n92 585
R534 B.n334 B.n333 585
R535 B.n332 B.n93 585
R536 B.n331 B.n330 585
R537 B.n329 B.n94 585
R538 B.n328 B.n327 585
R539 B.n326 B.n95 585
R540 B.n325 B.n324 585
R541 B.n323 B.n96 585
R542 B.n322 B.n321 585
R543 B.n320 B.n97 585
R544 B.n319 B.n318 585
R545 B.n317 B.n98 585
R546 B.n316 B.n315 585
R547 B.n314 B.n99 585
R548 B.n313 B.n312 585
R549 B.n311 B.n100 585
R550 B.n310 B.n309 585
R551 B.n308 B.n101 585
R552 B.n221 B.n134 585
R553 B.n223 B.n222 585
R554 B.n224 B.n133 585
R555 B.n226 B.n225 585
R556 B.n227 B.n132 585
R557 B.n229 B.n228 585
R558 B.n230 B.n131 585
R559 B.n232 B.n231 585
R560 B.n233 B.n130 585
R561 B.n235 B.n234 585
R562 B.n236 B.n129 585
R563 B.n238 B.n237 585
R564 B.n239 B.n128 585
R565 B.n241 B.n240 585
R566 B.n242 B.n127 585
R567 B.n244 B.n243 585
R568 B.n245 B.n126 585
R569 B.n247 B.n246 585
R570 B.n248 B.n125 585
R571 B.n250 B.n249 585
R572 B.n251 B.n124 585
R573 B.n253 B.n252 585
R574 B.n254 B.n123 585
R575 B.n256 B.n255 585
R576 B.n258 B.n257 585
R577 B.n259 B.n119 585
R578 B.n261 B.n260 585
R579 B.n262 B.n118 585
R580 B.n264 B.n263 585
R581 B.n265 B.n117 585
R582 B.n267 B.n266 585
R583 B.n268 B.n116 585
R584 B.n270 B.n269 585
R585 B.n272 B.n113 585
R586 B.n274 B.n273 585
R587 B.n275 B.n112 585
R588 B.n277 B.n276 585
R589 B.n278 B.n111 585
R590 B.n280 B.n279 585
R591 B.n281 B.n110 585
R592 B.n283 B.n282 585
R593 B.n284 B.n109 585
R594 B.n286 B.n285 585
R595 B.n287 B.n108 585
R596 B.n289 B.n288 585
R597 B.n290 B.n107 585
R598 B.n292 B.n291 585
R599 B.n293 B.n106 585
R600 B.n295 B.n294 585
R601 B.n296 B.n105 585
R602 B.n298 B.n297 585
R603 B.n299 B.n104 585
R604 B.n301 B.n300 585
R605 B.n302 B.n103 585
R606 B.n304 B.n303 585
R607 B.n305 B.n102 585
R608 B.n307 B.n306 585
R609 B.n220 B.n219 585
R610 B.n218 B.n135 585
R611 B.n217 B.n216 585
R612 B.n215 B.n136 585
R613 B.n214 B.n213 585
R614 B.n212 B.n137 585
R615 B.n211 B.n210 585
R616 B.n209 B.n138 585
R617 B.n208 B.n207 585
R618 B.n206 B.n139 585
R619 B.n205 B.n204 585
R620 B.n203 B.n140 585
R621 B.n202 B.n201 585
R622 B.n200 B.n141 585
R623 B.n199 B.n198 585
R624 B.n197 B.n142 585
R625 B.n196 B.n195 585
R626 B.n194 B.n143 585
R627 B.n193 B.n192 585
R628 B.n191 B.n144 585
R629 B.n190 B.n189 585
R630 B.n188 B.n145 585
R631 B.n187 B.n186 585
R632 B.n185 B.n146 585
R633 B.n184 B.n183 585
R634 B.n182 B.n147 585
R635 B.n181 B.n180 585
R636 B.n179 B.n148 585
R637 B.n178 B.n177 585
R638 B.n176 B.n149 585
R639 B.n175 B.n174 585
R640 B.n173 B.n150 585
R641 B.n172 B.n171 585
R642 B.n170 B.n151 585
R643 B.n169 B.n168 585
R644 B.n167 B.n152 585
R645 B.n166 B.n165 585
R646 B.n164 B.n153 585
R647 B.n163 B.n162 585
R648 B.n161 B.n154 585
R649 B.n160 B.n159 585
R650 B.n158 B.n155 585
R651 B.n157 B.n156 585
R652 B.n2 B.n0 585
R653 B.n593 B.n1 585
R654 B.n592 B.n591 585
R655 B.n590 B.n3 585
R656 B.n589 B.n588 585
R657 B.n587 B.n4 585
R658 B.n586 B.n585 585
R659 B.n584 B.n5 585
R660 B.n583 B.n582 585
R661 B.n581 B.n6 585
R662 B.n580 B.n579 585
R663 B.n578 B.n7 585
R664 B.n577 B.n576 585
R665 B.n575 B.n8 585
R666 B.n574 B.n573 585
R667 B.n572 B.n9 585
R668 B.n571 B.n570 585
R669 B.n569 B.n10 585
R670 B.n568 B.n567 585
R671 B.n566 B.n11 585
R672 B.n565 B.n564 585
R673 B.n563 B.n12 585
R674 B.n562 B.n561 585
R675 B.n560 B.n13 585
R676 B.n559 B.n558 585
R677 B.n557 B.n14 585
R678 B.n556 B.n555 585
R679 B.n554 B.n15 585
R680 B.n553 B.n552 585
R681 B.n551 B.n16 585
R682 B.n550 B.n549 585
R683 B.n548 B.n17 585
R684 B.n547 B.n546 585
R685 B.n545 B.n18 585
R686 B.n544 B.n543 585
R687 B.n542 B.n19 585
R688 B.n541 B.n540 585
R689 B.n539 B.n20 585
R690 B.n538 B.n537 585
R691 B.n536 B.n21 585
R692 B.n535 B.n534 585
R693 B.n533 B.n22 585
R694 B.n532 B.n531 585
R695 B.n530 B.n23 585
R696 B.n529 B.n528 585
R697 B.n595 B.n594 585
R698 B.n221 B.n220 535.745
R699 B.n528 B.n527 535.745
R700 B.n306 B.n101 535.745
R701 B.n442 B.n57 535.745
R702 B.n114 B.t5 346.351
R703 B.n44 B.t7 346.351
R704 B.n120 B.t2 346.351
R705 B.n36 B.t10 346.351
R706 B.n115 B.t4 267.224
R707 B.n45 B.t8 267.224
R708 B.n121 B.t1 267.224
R709 B.n37 B.t11 267.224
R710 B.n114 B.t3 247.543
R711 B.n120 B.t0 247.543
R712 B.n36 B.t9 247.543
R713 B.n44 B.t6 247.543
R714 B.n220 B.n135 163.367
R715 B.n216 B.n135 163.367
R716 B.n216 B.n215 163.367
R717 B.n215 B.n214 163.367
R718 B.n214 B.n137 163.367
R719 B.n210 B.n137 163.367
R720 B.n210 B.n209 163.367
R721 B.n209 B.n208 163.367
R722 B.n208 B.n139 163.367
R723 B.n204 B.n139 163.367
R724 B.n204 B.n203 163.367
R725 B.n203 B.n202 163.367
R726 B.n202 B.n141 163.367
R727 B.n198 B.n141 163.367
R728 B.n198 B.n197 163.367
R729 B.n197 B.n196 163.367
R730 B.n196 B.n143 163.367
R731 B.n192 B.n143 163.367
R732 B.n192 B.n191 163.367
R733 B.n191 B.n190 163.367
R734 B.n190 B.n145 163.367
R735 B.n186 B.n145 163.367
R736 B.n186 B.n185 163.367
R737 B.n185 B.n184 163.367
R738 B.n184 B.n147 163.367
R739 B.n180 B.n147 163.367
R740 B.n180 B.n179 163.367
R741 B.n179 B.n178 163.367
R742 B.n178 B.n149 163.367
R743 B.n174 B.n149 163.367
R744 B.n174 B.n173 163.367
R745 B.n173 B.n172 163.367
R746 B.n172 B.n151 163.367
R747 B.n168 B.n151 163.367
R748 B.n168 B.n167 163.367
R749 B.n167 B.n166 163.367
R750 B.n166 B.n153 163.367
R751 B.n162 B.n153 163.367
R752 B.n162 B.n161 163.367
R753 B.n161 B.n160 163.367
R754 B.n160 B.n155 163.367
R755 B.n156 B.n155 163.367
R756 B.n156 B.n2 163.367
R757 B.n594 B.n2 163.367
R758 B.n594 B.n593 163.367
R759 B.n593 B.n592 163.367
R760 B.n592 B.n3 163.367
R761 B.n588 B.n3 163.367
R762 B.n588 B.n587 163.367
R763 B.n587 B.n586 163.367
R764 B.n586 B.n5 163.367
R765 B.n582 B.n5 163.367
R766 B.n582 B.n581 163.367
R767 B.n581 B.n580 163.367
R768 B.n580 B.n7 163.367
R769 B.n576 B.n7 163.367
R770 B.n576 B.n575 163.367
R771 B.n575 B.n574 163.367
R772 B.n574 B.n9 163.367
R773 B.n570 B.n9 163.367
R774 B.n570 B.n569 163.367
R775 B.n569 B.n568 163.367
R776 B.n568 B.n11 163.367
R777 B.n564 B.n11 163.367
R778 B.n564 B.n563 163.367
R779 B.n563 B.n562 163.367
R780 B.n562 B.n13 163.367
R781 B.n558 B.n13 163.367
R782 B.n558 B.n557 163.367
R783 B.n557 B.n556 163.367
R784 B.n556 B.n15 163.367
R785 B.n552 B.n15 163.367
R786 B.n552 B.n551 163.367
R787 B.n551 B.n550 163.367
R788 B.n550 B.n17 163.367
R789 B.n546 B.n17 163.367
R790 B.n546 B.n545 163.367
R791 B.n545 B.n544 163.367
R792 B.n544 B.n19 163.367
R793 B.n540 B.n19 163.367
R794 B.n540 B.n539 163.367
R795 B.n539 B.n538 163.367
R796 B.n538 B.n21 163.367
R797 B.n534 B.n21 163.367
R798 B.n534 B.n533 163.367
R799 B.n533 B.n532 163.367
R800 B.n532 B.n23 163.367
R801 B.n528 B.n23 163.367
R802 B.n222 B.n221 163.367
R803 B.n222 B.n133 163.367
R804 B.n226 B.n133 163.367
R805 B.n227 B.n226 163.367
R806 B.n228 B.n227 163.367
R807 B.n228 B.n131 163.367
R808 B.n232 B.n131 163.367
R809 B.n233 B.n232 163.367
R810 B.n234 B.n233 163.367
R811 B.n234 B.n129 163.367
R812 B.n238 B.n129 163.367
R813 B.n239 B.n238 163.367
R814 B.n240 B.n239 163.367
R815 B.n240 B.n127 163.367
R816 B.n244 B.n127 163.367
R817 B.n245 B.n244 163.367
R818 B.n246 B.n245 163.367
R819 B.n246 B.n125 163.367
R820 B.n250 B.n125 163.367
R821 B.n251 B.n250 163.367
R822 B.n252 B.n251 163.367
R823 B.n252 B.n123 163.367
R824 B.n256 B.n123 163.367
R825 B.n257 B.n256 163.367
R826 B.n257 B.n119 163.367
R827 B.n261 B.n119 163.367
R828 B.n262 B.n261 163.367
R829 B.n263 B.n262 163.367
R830 B.n263 B.n117 163.367
R831 B.n267 B.n117 163.367
R832 B.n268 B.n267 163.367
R833 B.n269 B.n268 163.367
R834 B.n269 B.n113 163.367
R835 B.n274 B.n113 163.367
R836 B.n275 B.n274 163.367
R837 B.n276 B.n275 163.367
R838 B.n276 B.n111 163.367
R839 B.n280 B.n111 163.367
R840 B.n281 B.n280 163.367
R841 B.n282 B.n281 163.367
R842 B.n282 B.n109 163.367
R843 B.n286 B.n109 163.367
R844 B.n287 B.n286 163.367
R845 B.n288 B.n287 163.367
R846 B.n288 B.n107 163.367
R847 B.n292 B.n107 163.367
R848 B.n293 B.n292 163.367
R849 B.n294 B.n293 163.367
R850 B.n294 B.n105 163.367
R851 B.n298 B.n105 163.367
R852 B.n299 B.n298 163.367
R853 B.n300 B.n299 163.367
R854 B.n300 B.n103 163.367
R855 B.n304 B.n103 163.367
R856 B.n305 B.n304 163.367
R857 B.n306 B.n305 163.367
R858 B.n310 B.n101 163.367
R859 B.n311 B.n310 163.367
R860 B.n312 B.n311 163.367
R861 B.n312 B.n99 163.367
R862 B.n316 B.n99 163.367
R863 B.n317 B.n316 163.367
R864 B.n318 B.n317 163.367
R865 B.n318 B.n97 163.367
R866 B.n322 B.n97 163.367
R867 B.n323 B.n322 163.367
R868 B.n324 B.n323 163.367
R869 B.n324 B.n95 163.367
R870 B.n328 B.n95 163.367
R871 B.n329 B.n328 163.367
R872 B.n330 B.n329 163.367
R873 B.n330 B.n93 163.367
R874 B.n334 B.n93 163.367
R875 B.n335 B.n334 163.367
R876 B.n336 B.n335 163.367
R877 B.n336 B.n91 163.367
R878 B.n340 B.n91 163.367
R879 B.n341 B.n340 163.367
R880 B.n342 B.n341 163.367
R881 B.n342 B.n89 163.367
R882 B.n346 B.n89 163.367
R883 B.n347 B.n346 163.367
R884 B.n348 B.n347 163.367
R885 B.n348 B.n87 163.367
R886 B.n352 B.n87 163.367
R887 B.n353 B.n352 163.367
R888 B.n354 B.n353 163.367
R889 B.n354 B.n85 163.367
R890 B.n358 B.n85 163.367
R891 B.n359 B.n358 163.367
R892 B.n360 B.n359 163.367
R893 B.n360 B.n83 163.367
R894 B.n364 B.n83 163.367
R895 B.n365 B.n364 163.367
R896 B.n366 B.n365 163.367
R897 B.n366 B.n81 163.367
R898 B.n370 B.n81 163.367
R899 B.n371 B.n370 163.367
R900 B.n372 B.n371 163.367
R901 B.n372 B.n79 163.367
R902 B.n376 B.n79 163.367
R903 B.n377 B.n376 163.367
R904 B.n378 B.n377 163.367
R905 B.n378 B.n77 163.367
R906 B.n382 B.n77 163.367
R907 B.n383 B.n382 163.367
R908 B.n384 B.n383 163.367
R909 B.n384 B.n75 163.367
R910 B.n388 B.n75 163.367
R911 B.n389 B.n388 163.367
R912 B.n390 B.n389 163.367
R913 B.n390 B.n73 163.367
R914 B.n394 B.n73 163.367
R915 B.n395 B.n394 163.367
R916 B.n396 B.n395 163.367
R917 B.n396 B.n71 163.367
R918 B.n400 B.n71 163.367
R919 B.n401 B.n400 163.367
R920 B.n402 B.n401 163.367
R921 B.n402 B.n69 163.367
R922 B.n406 B.n69 163.367
R923 B.n407 B.n406 163.367
R924 B.n408 B.n407 163.367
R925 B.n408 B.n67 163.367
R926 B.n412 B.n67 163.367
R927 B.n413 B.n412 163.367
R928 B.n414 B.n413 163.367
R929 B.n414 B.n65 163.367
R930 B.n418 B.n65 163.367
R931 B.n419 B.n418 163.367
R932 B.n420 B.n419 163.367
R933 B.n420 B.n63 163.367
R934 B.n424 B.n63 163.367
R935 B.n425 B.n424 163.367
R936 B.n426 B.n425 163.367
R937 B.n426 B.n61 163.367
R938 B.n430 B.n61 163.367
R939 B.n431 B.n430 163.367
R940 B.n432 B.n431 163.367
R941 B.n432 B.n59 163.367
R942 B.n436 B.n59 163.367
R943 B.n437 B.n436 163.367
R944 B.n438 B.n437 163.367
R945 B.n438 B.n57 163.367
R946 B.n527 B.n526 163.367
R947 B.n526 B.n25 163.367
R948 B.n522 B.n25 163.367
R949 B.n522 B.n521 163.367
R950 B.n521 B.n520 163.367
R951 B.n520 B.n27 163.367
R952 B.n516 B.n27 163.367
R953 B.n516 B.n515 163.367
R954 B.n515 B.n514 163.367
R955 B.n514 B.n29 163.367
R956 B.n510 B.n29 163.367
R957 B.n510 B.n509 163.367
R958 B.n509 B.n508 163.367
R959 B.n508 B.n31 163.367
R960 B.n504 B.n31 163.367
R961 B.n504 B.n503 163.367
R962 B.n503 B.n502 163.367
R963 B.n502 B.n33 163.367
R964 B.n498 B.n33 163.367
R965 B.n498 B.n497 163.367
R966 B.n497 B.n496 163.367
R967 B.n496 B.n35 163.367
R968 B.n492 B.n35 163.367
R969 B.n492 B.n491 163.367
R970 B.n491 B.n39 163.367
R971 B.n487 B.n39 163.367
R972 B.n487 B.n486 163.367
R973 B.n486 B.n485 163.367
R974 B.n485 B.n41 163.367
R975 B.n481 B.n41 163.367
R976 B.n481 B.n480 163.367
R977 B.n480 B.n479 163.367
R978 B.n479 B.n43 163.367
R979 B.n474 B.n43 163.367
R980 B.n474 B.n473 163.367
R981 B.n473 B.n472 163.367
R982 B.n472 B.n47 163.367
R983 B.n468 B.n47 163.367
R984 B.n468 B.n467 163.367
R985 B.n467 B.n466 163.367
R986 B.n466 B.n49 163.367
R987 B.n462 B.n49 163.367
R988 B.n462 B.n461 163.367
R989 B.n461 B.n460 163.367
R990 B.n460 B.n51 163.367
R991 B.n456 B.n51 163.367
R992 B.n456 B.n455 163.367
R993 B.n455 B.n454 163.367
R994 B.n454 B.n53 163.367
R995 B.n450 B.n53 163.367
R996 B.n450 B.n449 163.367
R997 B.n449 B.n448 163.367
R998 B.n448 B.n55 163.367
R999 B.n444 B.n55 163.367
R1000 B.n444 B.n443 163.367
R1001 B.n443 B.n442 163.367
R1002 B.n115 B.n114 79.1278
R1003 B.n121 B.n120 79.1278
R1004 B.n37 B.n36 79.1278
R1005 B.n45 B.n44 79.1278
R1006 B.n271 B.n115 59.5399
R1007 B.n122 B.n121 59.5399
R1008 B.n38 B.n37 59.5399
R1009 B.n477 B.n45 59.5399
R1010 B.n529 B.n24 34.8103
R1011 B.n441 B.n440 34.8103
R1012 B.n308 B.n307 34.8103
R1013 B.n219 B.n134 34.8103
R1014 B B.n595 18.0485
R1015 B.n525 B.n24 10.6151
R1016 B.n525 B.n524 10.6151
R1017 B.n524 B.n523 10.6151
R1018 B.n523 B.n26 10.6151
R1019 B.n519 B.n26 10.6151
R1020 B.n519 B.n518 10.6151
R1021 B.n518 B.n517 10.6151
R1022 B.n517 B.n28 10.6151
R1023 B.n513 B.n28 10.6151
R1024 B.n513 B.n512 10.6151
R1025 B.n512 B.n511 10.6151
R1026 B.n511 B.n30 10.6151
R1027 B.n507 B.n30 10.6151
R1028 B.n507 B.n506 10.6151
R1029 B.n506 B.n505 10.6151
R1030 B.n505 B.n32 10.6151
R1031 B.n501 B.n32 10.6151
R1032 B.n501 B.n500 10.6151
R1033 B.n500 B.n499 10.6151
R1034 B.n499 B.n34 10.6151
R1035 B.n495 B.n34 10.6151
R1036 B.n495 B.n494 10.6151
R1037 B.n494 B.n493 10.6151
R1038 B.n490 B.n489 10.6151
R1039 B.n489 B.n488 10.6151
R1040 B.n488 B.n40 10.6151
R1041 B.n484 B.n40 10.6151
R1042 B.n484 B.n483 10.6151
R1043 B.n483 B.n482 10.6151
R1044 B.n482 B.n42 10.6151
R1045 B.n478 B.n42 10.6151
R1046 B.n476 B.n475 10.6151
R1047 B.n475 B.n46 10.6151
R1048 B.n471 B.n46 10.6151
R1049 B.n471 B.n470 10.6151
R1050 B.n470 B.n469 10.6151
R1051 B.n469 B.n48 10.6151
R1052 B.n465 B.n48 10.6151
R1053 B.n465 B.n464 10.6151
R1054 B.n464 B.n463 10.6151
R1055 B.n463 B.n50 10.6151
R1056 B.n459 B.n50 10.6151
R1057 B.n459 B.n458 10.6151
R1058 B.n458 B.n457 10.6151
R1059 B.n457 B.n52 10.6151
R1060 B.n453 B.n52 10.6151
R1061 B.n453 B.n452 10.6151
R1062 B.n452 B.n451 10.6151
R1063 B.n451 B.n54 10.6151
R1064 B.n447 B.n54 10.6151
R1065 B.n447 B.n446 10.6151
R1066 B.n446 B.n445 10.6151
R1067 B.n445 B.n56 10.6151
R1068 B.n441 B.n56 10.6151
R1069 B.n309 B.n308 10.6151
R1070 B.n309 B.n100 10.6151
R1071 B.n313 B.n100 10.6151
R1072 B.n314 B.n313 10.6151
R1073 B.n315 B.n314 10.6151
R1074 B.n315 B.n98 10.6151
R1075 B.n319 B.n98 10.6151
R1076 B.n320 B.n319 10.6151
R1077 B.n321 B.n320 10.6151
R1078 B.n321 B.n96 10.6151
R1079 B.n325 B.n96 10.6151
R1080 B.n326 B.n325 10.6151
R1081 B.n327 B.n326 10.6151
R1082 B.n327 B.n94 10.6151
R1083 B.n331 B.n94 10.6151
R1084 B.n332 B.n331 10.6151
R1085 B.n333 B.n332 10.6151
R1086 B.n333 B.n92 10.6151
R1087 B.n337 B.n92 10.6151
R1088 B.n338 B.n337 10.6151
R1089 B.n339 B.n338 10.6151
R1090 B.n339 B.n90 10.6151
R1091 B.n343 B.n90 10.6151
R1092 B.n344 B.n343 10.6151
R1093 B.n345 B.n344 10.6151
R1094 B.n345 B.n88 10.6151
R1095 B.n349 B.n88 10.6151
R1096 B.n350 B.n349 10.6151
R1097 B.n351 B.n350 10.6151
R1098 B.n351 B.n86 10.6151
R1099 B.n355 B.n86 10.6151
R1100 B.n356 B.n355 10.6151
R1101 B.n357 B.n356 10.6151
R1102 B.n357 B.n84 10.6151
R1103 B.n361 B.n84 10.6151
R1104 B.n362 B.n361 10.6151
R1105 B.n363 B.n362 10.6151
R1106 B.n363 B.n82 10.6151
R1107 B.n367 B.n82 10.6151
R1108 B.n368 B.n367 10.6151
R1109 B.n369 B.n368 10.6151
R1110 B.n369 B.n80 10.6151
R1111 B.n373 B.n80 10.6151
R1112 B.n374 B.n373 10.6151
R1113 B.n375 B.n374 10.6151
R1114 B.n375 B.n78 10.6151
R1115 B.n379 B.n78 10.6151
R1116 B.n380 B.n379 10.6151
R1117 B.n381 B.n380 10.6151
R1118 B.n381 B.n76 10.6151
R1119 B.n385 B.n76 10.6151
R1120 B.n386 B.n385 10.6151
R1121 B.n387 B.n386 10.6151
R1122 B.n387 B.n74 10.6151
R1123 B.n391 B.n74 10.6151
R1124 B.n392 B.n391 10.6151
R1125 B.n393 B.n392 10.6151
R1126 B.n393 B.n72 10.6151
R1127 B.n397 B.n72 10.6151
R1128 B.n398 B.n397 10.6151
R1129 B.n399 B.n398 10.6151
R1130 B.n399 B.n70 10.6151
R1131 B.n403 B.n70 10.6151
R1132 B.n404 B.n403 10.6151
R1133 B.n405 B.n404 10.6151
R1134 B.n405 B.n68 10.6151
R1135 B.n409 B.n68 10.6151
R1136 B.n410 B.n409 10.6151
R1137 B.n411 B.n410 10.6151
R1138 B.n411 B.n66 10.6151
R1139 B.n415 B.n66 10.6151
R1140 B.n416 B.n415 10.6151
R1141 B.n417 B.n416 10.6151
R1142 B.n417 B.n64 10.6151
R1143 B.n421 B.n64 10.6151
R1144 B.n422 B.n421 10.6151
R1145 B.n423 B.n422 10.6151
R1146 B.n423 B.n62 10.6151
R1147 B.n427 B.n62 10.6151
R1148 B.n428 B.n427 10.6151
R1149 B.n429 B.n428 10.6151
R1150 B.n429 B.n60 10.6151
R1151 B.n433 B.n60 10.6151
R1152 B.n434 B.n433 10.6151
R1153 B.n435 B.n434 10.6151
R1154 B.n435 B.n58 10.6151
R1155 B.n439 B.n58 10.6151
R1156 B.n440 B.n439 10.6151
R1157 B.n223 B.n134 10.6151
R1158 B.n224 B.n223 10.6151
R1159 B.n225 B.n224 10.6151
R1160 B.n225 B.n132 10.6151
R1161 B.n229 B.n132 10.6151
R1162 B.n230 B.n229 10.6151
R1163 B.n231 B.n230 10.6151
R1164 B.n231 B.n130 10.6151
R1165 B.n235 B.n130 10.6151
R1166 B.n236 B.n235 10.6151
R1167 B.n237 B.n236 10.6151
R1168 B.n237 B.n128 10.6151
R1169 B.n241 B.n128 10.6151
R1170 B.n242 B.n241 10.6151
R1171 B.n243 B.n242 10.6151
R1172 B.n243 B.n126 10.6151
R1173 B.n247 B.n126 10.6151
R1174 B.n248 B.n247 10.6151
R1175 B.n249 B.n248 10.6151
R1176 B.n249 B.n124 10.6151
R1177 B.n253 B.n124 10.6151
R1178 B.n254 B.n253 10.6151
R1179 B.n255 B.n254 10.6151
R1180 B.n259 B.n258 10.6151
R1181 B.n260 B.n259 10.6151
R1182 B.n260 B.n118 10.6151
R1183 B.n264 B.n118 10.6151
R1184 B.n265 B.n264 10.6151
R1185 B.n266 B.n265 10.6151
R1186 B.n266 B.n116 10.6151
R1187 B.n270 B.n116 10.6151
R1188 B.n273 B.n272 10.6151
R1189 B.n273 B.n112 10.6151
R1190 B.n277 B.n112 10.6151
R1191 B.n278 B.n277 10.6151
R1192 B.n279 B.n278 10.6151
R1193 B.n279 B.n110 10.6151
R1194 B.n283 B.n110 10.6151
R1195 B.n284 B.n283 10.6151
R1196 B.n285 B.n284 10.6151
R1197 B.n285 B.n108 10.6151
R1198 B.n289 B.n108 10.6151
R1199 B.n290 B.n289 10.6151
R1200 B.n291 B.n290 10.6151
R1201 B.n291 B.n106 10.6151
R1202 B.n295 B.n106 10.6151
R1203 B.n296 B.n295 10.6151
R1204 B.n297 B.n296 10.6151
R1205 B.n297 B.n104 10.6151
R1206 B.n301 B.n104 10.6151
R1207 B.n302 B.n301 10.6151
R1208 B.n303 B.n302 10.6151
R1209 B.n303 B.n102 10.6151
R1210 B.n307 B.n102 10.6151
R1211 B.n219 B.n218 10.6151
R1212 B.n218 B.n217 10.6151
R1213 B.n217 B.n136 10.6151
R1214 B.n213 B.n136 10.6151
R1215 B.n213 B.n212 10.6151
R1216 B.n212 B.n211 10.6151
R1217 B.n211 B.n138 10.6151
R1218 B.n207 B.n138 10.6151
R1219 B.n207 B.n206 10.6151
R1220 B.n206 B.n205 10.6151
R1221 B.n205 B.n140 10.6151
R1222 B.n201 B.n140 10.6151
R1223 B.n201 B.n200 10.6151
R1224 B.n200 B.n199 10.6151
R1225 B.n199 B.n142 10.6151
R1226 B.n195 B.n142 10.6151
R1227 B.n195 B.n194 10.6151
R1228 B.n194 B.n193 10.6151
R1229 B.n193 B.n144 10.6151
R1230 B.n189 B.n144 10.6151
R1231 B.n189 B.n188 10.6151
R1232 B.n188 B.n187 10.6151
R1233 B.n187 B.n146 10.6151
R1234 B.n183 B.n146 10.6151
R1235 B.n183 B.n182 10.6151
R1236 B.n182 B.n181 10.6151
R1237 B.n181 B.n148 10.6151
R1238 B.n177 B.n148 10.6151
R1239 B.n177 B.n176 10.6151
R1240 B.n176 B.n175 10.6151
R1241 B.n175 B.n150 10.6151
R1242 B.n171 B.n150 10.6151
R1243 B.n171 B.n170 10.6151
R1244 B.n170 B.n169 10.6151
R1245 B.n169 B.n152 10.6151
R1246 B.n165 B.n152 10.6151
R1247 B.n165 B.n164 10.6151
R1248 B.n164 B.n163 10.6151
R1249 B.n163 B.n154 10.6151
R1250 B.n159 B.n154 10.6151
R1251 B.n159 B.n158 10.6151
R1252 B.n158 B.n157 10.6151
R1253 B.n157 B.n0 10.6151
R1254 B.n591 B.n1 10.6151
R1255 B.n591 B.n590 10.6151
R1256 B.n590 B.n589 10.6151
R1257 B.n589 B.n4 10.6151
R1258 B.n585 B.n4 10.6151
R1259 B.n585 B.n584 10.6151
R1260 B.n584 B.n583 10.6151
R1261 B.n583 B.n6 10.6151
R1262 B.n579 B.n6 10.6151
R1263 B.n579 B.n578 10.6151
R1264 B.n578 B.n577 10.6151
R1265 B.n577 B.n8 10.6151
R1266 B.n573 B.n8 10.6151
R1267 B.n573 B.n572 10.6151
R1268 B.n572 B.n571 10.6151
R1269 B.n571 B.n10 10.6151
R1270 B.n567 B.n10 10.6151
R1271 B.n567 B.n566 10.6151
R1272 B.n566 B.n565 10.6151
R1273 B.n565 B.n12 10.6151
R1274 B.n561 B.n12 10.6151
R1275 B.n561 B.n560 10.6151
R1276 B.n560 B.n559 10.6151
R1277 B.n559 B.n14 10.6151
R1278 B.n555 B.n14 10.6151
R1279 B.n555 B.n554 10.6151
R1280 B.n554 B.n553 10.6151
R1281 B.n553 B.n16 10.6151
R1282 B.n549 B.n16 10.6151
R1283 B.n549 B.n548 10.6151
R1284 B.n548 B.n547 10.6151
R1285 B.n547 B.n18 10.6151
R1286 B.n543 B.n18 10.6151
R1287 B.n543 B.n542 10.6151
R1288 B.n542 B.n541 10.6151
R1289 B.n541 B.n20 10.6151
R1290 B.n537 B.n20 10.6151
R1291 B.n537 B.n536 10.6151
R1292 B.n536 B.n535 10.6151
R1293 B.n535 B.n22 10.6151
R1294 B.n531 B.n22 10.6151
R1295 B.n531 B.n530 10.6151
R1296 B.n530 B.n529 10.6151
R1297 B.n490 B.n38 6.5566
R1298 B.n478 B.n477 6.5566
R1299 B.n258 B.n122 6.5566
R1300 B.n271 B.n270 6.5566
R1301 B.n493 B.n38 4.05904
R1302 B.n477 B.n476 4.05904
R1303 B.n255 B.n122 4.05904
R1304 B.n272 B.n271 4.05904
R1305 B.n595 B.n0 2.81026
R1306 B.n595 B.n1 2.81026
R1307 VP.n21 VP.n20 161.3
R1308 VP.n19 VP.n1 161.3
R1309 VP.n18 VP.n17 161.3
R1310 VP.n16 VP.n2 161.3
R1311 VP.n15 VP.n14 161.3
R1312 VP.n13 VP.n3 161.3
R1313 VP.n12 VP.n11 161.3
R1314 VP.n10 VP.n4 161.3
R1315 VP.n9 VP.n8 161.3
R1316 VP.n7 VP.n6 88.1101
R1317 VP.n22 VP.n0 88.1101
R1318 VP.n5 VP.t3 71.8584
R1319 VP.n5 VP.t0 70.5207
R1320 VP.n6 VP.n5 47.1667
R1321 VP.n14 VP.n13 40.4934
R1322 VP.n14 VP.n2 40.4934
R1323 VP.n7 VP.t2 38.2392
R1324 VP.n0 VP.t1 38.2392
R1325 VP.n8 VP.n4 24.4675
R1326 VP.n12 VP.n4 24.4675
R1327 VP.n13 VP.n12 24.4675
R1328 VP.n18 VP.n2 24.4675
R1329 VP.n19 VP.n18 24.4675
R1330 VP.n20 VP.n19 24.4675
R1331 VP.n8 VP.n7 1.95786
R1332 VP.n20 VP.n0 1.95786
R1333 VP.n9 VP.n6 0.354971
R1334 VP.n22 VP.n21 0.354971
R1335 VP VP.n22 0.26696
R1336 VP.n10 VP.n9 0.189894
R1337 VP.n11 VP.n10 0.189894
R1338 VP.n11 VP.n3 0.189894
R1339 VP.n15 VP.n3 0.189894
R1340 VP.n16 VP.n15 0.189894
R1341 VP.n17 VP.n16 0.189894
R1342 VP.n17 VP.n1 0.189894
R1343 VP.n21 VP.n1 0.189894
R1344 VDD1 VDD1.n1 131.245
R1345 VDD1 VDD1.n0 91.3826
R1346 VDD1.n0 VDD1.t0 5.46353
R1347 VDD1.n0 VDD1.t3 5.46353
R1348 VDD1.n1 VDD1.t1 5.46353
R1349 VDD1.n1 VDD1.t2 5.46353
C0 VDD2 VP 0.467336f
C1 B VP 1.98865f
C2 VDD1 w_n3418_n2158# 1.50279f
C3 VDD2 w_n3418_n2158# 1.58426f
C4 VN VTAIL 3.1849f
C5 B w_n3418_n2158# 8.97924f
C6 VP VN 5.90152f
C7 VDD2 VDD1 1.30463f
C8 VP VTAIL 3.19901f
C9 B VDD1 1.30282f
C10 VN w_n3418_n2158# 5.89792f
C11 VDD2 B 1.374f
C12 w_n3418_n2158# VTAIL 2.69249f
C13 VP w_n3418_n2158# 6.34023f
C14 VDD1 VN 0.149893f
C15 VDD1 VTAIL 4.46501f
C16 VDD2 VN 2.66471f
C17 B VN 1.24932f
C18 VDD1 VP 2.98112f
C19 VDD2 VTAIL 4.52693f
C20 B VTAIL 3.30134f
C21 VDD2 VSUBS 0.995773f
C22 VDD1 VSUBS 5.75501f
C23 VTAIL VSUBS 0.795761f
C24 VN VSUBS 6.03086f
C25 VP VSUBS 2.505085f
C26 B VSUBS 4.755225f
C27 w_n3418_n2158# VSUBS 92.080894f
C28 VDD1.t0 VSUBS 0.13751f
C29 VDD1.t3 VSUBS 0.13751f
C30 VDD1.n0 VSUBS 0.907705f
C31 VDD1.t1 VSUBS 0.13751f
C32 VDD1.t2 VSUBS 0.13751f
C33 VDD1.n1 VSUBS 1.44257f
C34 VP.t1 VSUBS 2.18032f
C35 VP.n0 VSUBS 0.939026f
C36 VP.n1 VSUBS 0.036938f
C37 VP.n2 VSUBS 0.073413f
C38 VP.n3 VSUBS 0.036938f
C39 VP.n4 VSUBS 0.068843f
C40 VP.t3 VSUBS 2.69802f
C41 VP.t0 VSUBS 2.67795f
C42 VP.n5 VSUBS 3.73055f
C43 VP.n6 VSUBS 1.96303f
C44 VP.t2 VSUBS 2.18032f
C45 VP.n7 VSUBS 0.939026f
C46 VP.n8 VSUBS 0.037574f
C47 VP.n9 VSUBS 0.059617f
C48 VP.n10 VSUBS 0.036938f
C49 VP.n11 VSUBS 0.036938f
C50 VP.n12 VSUBS 0.068843f
C51 VP.n13 VSUBS 0.073413f
C52 VP.n14 VSUBS 0.029861f
C53 VP.n15 VSUBS 0.036938f
C54 VP.n16 VSUBS 0.036938f
C55 VP.n17 VSUBS 0.036938f
C56 VP.n18 VSUBS 0.068843f
C57 VP.n19 VSUBS 0.068843f
C58 VP.n20 VSUBS 0.037574f
C59 VP.n21 VSUBS 0.059617f
C60 VP.n22 VSUBS 0.113421f
C61 B.n0 VSUBS 0.004994f
C62 B.n1 VSUBS 0.004994f
C63 B.n2 VSUBS 0.007897f
C64 B.n3 VSUBS 0.007897f
C65 B.n4 VSUBS 0.007897f
C66 B.n5 VSUBS 0.007897f
C67 B.n6 VSUBS 0.007897f
C68 B.n7 VSUBS 0.007897f
C69 B.n8 VSUBS 0.007897f
C70 B.n9 VSUBS 0.007897f
C71 B.n10 VSUBS 0.007897f
C72 B.n11 VSUBS 0.007897f
C73 B.n12 VSUBS 0.007897f
C74 B.n13 VSUBS 0.007897f
C75 B.n14 VSUBS 0.007897f
C76 B.n15 VSUBS 0.007897f
C77 B.n16 VSUBS 0.007897f
C78 B.n17 VSUBS 0.007897f
C79 B.n18 VSUBS 0.007897f
C80 B.n19 VSUBS 0.007897f
C81 B.n20 VSUBS 0.007897f
C82 B.n21 VSUBS 0.007897f
C83 B.n22 VSUBS 0.007897f
C84 B.n23 VSUBS 0.007897f
C85 B.n24 VSUBS 0.019694f
C86 B.n25 VSUBS 0.007897f
C87 B.n26 VSUBS 0.007897f
C88 B.n27 VSUBS 0.007897f
C89 B.n28 VSUBS 0.007897f
C90 B.n29 VSUBS 0.007897f
C91 B.n30 VSUBS 0.007897f
C92 B.n31 VSUBS 0.007897f
C93 B.n32 VSUBS 0.007897f
C94 B.n33 VSUBS 0.007897f
C95 B.n34 VSUBS 0.007897f
C96 B.n35 VSUBS 0.007897f
C97 B.t11 VSUBS 0.099868f
C98 B.t10 VSUBS 0.138626f
C99 B.t9 VSUBS 1.2099f
C100 B.n36 VSUBS 0.229306f
C101 B.n37 VSUBS 0.180913f
C102 B.n38 VSUBS 0.018297f
C103 B.n39 VSUBS 0.007897f
C104 B.n40 VSUBS 0.007897f
C105 B.n41 VSUBS 0.007897f
C106 B.n42 VSUBS 0.007897f
C107 B.n43 VSUBS 0.007897f
C108 B.t8 VSUBS 0.09987f
C109 B.t7 VSUBS 0.138628f
C110 B.t6 VSUBS 1.2099f
C111 B.n44 VSUBS 0.229304f
C112 B.n45 VSUBS 0.180911f
C113 B.n46 VSUBS 0.007897f
C114 B.n47 VSUBS 0.007897f
C115 B.n48 VSUBS 0.007897f
C116 B.n49 VSUBS 0.007897f
C117 B.n50 VSUBS 0.007897f
C118 B.n51 VSUBS 0.007897f
C119 B.n52 VSUBS 0.007897f
C120 B.n53 VSUBS 0.007897f
C121 B.n54 VSUBS 0.007897f
C122 B.n55 VSUBS 0.007897f
C123 B.n56 VSUBS 0.007897f
C124 B.n57 VSUBS 0.018862f
C125 B.n58 VSUBS 0.007897f
C126 B.n59 VSUBS 0.007897f
C127 B.n60 VSUBS 0.007897f
C128 B.n61 VSUBS 0.007897f
C129 B.n62 VSUBS 0.007897f
C130 B.n63 VSUBS 0.007897f
C131 B.n64 VSUBS 0.007897f
C132 B.n65 VSUBS 0.007897f
C133 B.n66 VSUBS 0.007897f
C134 B.n67 VSUBS 0.007897f
C135 B.n68 VSUBS 0.007897f
C136 B.n69 VSUBS 0.007897f
C137 B.n70 VSUBS 0.007897f
C138 B.n71 VSUBS 0.007897f
C139 B.n72 VSUBS 0.007897f
C140 B.n73 VSUBS 0.007897f
C141 B.n74 VSUBS 0.007897f
C142 B.n75 VSUBS 0.007897f
C143 B.n76 VSUBS 0.007897f
C144 B.n77 VSUBS 0.007897f
C145 B.n78 VSUBS 0.007897f
C146 B.n79 VSUBS 0.007897f
C147 B.n80 VSUBS 0.007897f
C148 B.n81 VSUBS 0.007897f
C149 B.n82 VSUBS 0.007897f
C150 B.n83 VSUBS 0.007897f
C151 B.n84 VSUBS 0.007897f
C152 B.n85 VSUBS 0.007897f
C153 B.n86 VSUBS 0.007897f
C154 B.n87 VSUBS 0.007897f
C155 B.n88 VSUBS 0.007897f
C156 B.n89 VSUBS 0.007897f
C157 B.n90 VSUBS 0.007897f
C158 B.n91 VSUBS 0.007897f
C159 B.n92 VSUBS 0.007897f
C160 B.n93 VSUBS 0.007897f
C161 B.n94 VSUBS 0.007897f
C162 B.n95 VSUBS 0.007897f
C163 B.n96 VSUBS 0.007897f
C164 B.n97 VSUBS 0.007897f
C165 B.n98 VSUBS 0.007897f
C166 B.n99 VSUBS 0.007897f
C167 B.n100 VSUBS 0.007897f
C168 B.n101 VSUBS 0.018862f
C169 B.n102 VSUBS 0.007897f
C170 B.n103 VSUBS 0.007897f
C171 B.n104 VSUBS 0.007897f
C172 B.n105 VSUBS 0.007897f
C173 B.n106 VSUBS 0.007897f
C174 B.n107 VSUBS 0.007897f
C175 B.n108 VSUBS 0.007897f
C176 B.n109 VSUBS 0.007897f
C177 B.n110 VSUBS 0.007897f
C178 B.n111 VSUBS 0.007897f
C179 B.n112 VSUBS 0.007897f
C180 B.n113 VSUBS 0.007897f
C181 B.t4 VSUBS 0.09987f
C182 B.t5 VSUBS 0.138628f
C183 B.t3 VSUBS 1.2099f
C184 B.n114 VSUBS 0.229304f
C185 B.n115 VSUBS 0.180911f
C186 B.n116 VSUBS 0.007897f
C187 B.n117 VSUBS 0.007897f
C188 B.n118 VSUBS 0.007897f
C189 B.n119 VSUBS 0.007897f
C190 B.t1 VSUBS 0.099868f
C191 B.t2 VSUBS 0.138626f
C192 B.t0 VSUBS 1.2099f
C193 B.n120 VSUBS 0.229306f
C194 B.n121 VSUBS 0.180913f
C195 B.n122 VSUBS 0.018297f
C196 B.n123 VSUBS 0.007897f
C197 B.n124 VSUBS 0.007897f
C198 B.n125 VSUBS 0.007897f
C199 B.n126 VSUBS 0.007897f
C200 B.n127 VSUBS 0.007897f
C201 B.n128 VSUBS 0.007897f
C202 B.n129 VSUBS 0.007897f
C203 B.n130 VSUBS 0.007897f
C204 B.n131 VSUBS 0.007897f
C205 B.n132 VSUBS 0.007897f
C206 B.n133 VSUBS 0.007897f
C207 B.n134 VSUBS 0.019694f
C208 B.n135 VSUBS 0.007897f
C209 B.n136 VSUBS 0.007897f
C210 B.n137 VSUBS 0.007897f
C211 B.n138 VSUBS 0.007897f
C212 B.n139 VSUBS 0.007897f
C213 B.n140 VSUBS 0.007897f
C214 B.n141 VSUBS 0.007897f
C215 B.n142 VSUBS 0.007897f
C216 B.n143 VSUBS 0.007897f
C217 B.n144 VSUBS 0.007897f
C218 B.n145 VSUBS 0.007897f
C219 B.n146 VSUBS 0.007897f
C220 B.n147 VSUBS 0.007897f
C221 B.n148 VSUBS 0.007897f
C222 B.n149 VSUBS 0.007897f
C223 B.n150 VSUBS 0.007897f
C224 B.n151 VSUBS 0.007897f
C225 B.n152 VSUBS 0.007897f
C226 B.n153 VSUBS 0.007897f
C227 B.n154 VSUBS 0.007897f
C228 B.n155 VSUBS 0.007897f
C229 B.n156 VSUBS 0.007897f
C230 B.n157 VSUBS 0.007897f
C231 B.n158 VSUBS 0.007897f
C232 B.n159 VSUBS 0.007897f
C233 B.n160 VSUBS 0.007897f
C234 B.n161 VSUBS 0.007897f
C235 B.n162 VSUBS 0.007897f
C236 B.n163 VSUBS 0.007897f
C237 B.n164 VSUBS 0.007897f
C238 B.n165 VSUBS 0.007897f
C239 B.n166 VSUBS 0.007897f
C240 B.n167 VSUBS 0.007897f
C241 B.n168 VSUBS 0.007897f
C242 B.n169 VSUBS 0.007897f
C243 B.n170 VSUBS 0.007897f
C244 B.n171 VSUBS 0.007897f
C245 B.n172 VSUBS 0.007897f
C246 B.n173 VSUBS 0.007897f
C247 B.n174 VSUBS 0.007897f
C248 B.n175 VSUBS 0.007897f
C249 B.n176 VSUBS 0.007897f
C250 B.n177 VSUBS 0.007897f
C251 B.n178 VSUBS 0.007897f
C252 B.n179 VSUBS 0.007897f
C253 B.n180 VSUBS 0.007897f
C254 B.n181 VSUBS 0.007897f
C255 B.n182 VSUBS 0.007897f
C256 B.n183 VSUBS 0.007897f
C257 B.n184 VSUBS 0.007897f
C258 B.n185 VSUBS 0.007897f
C259 B.n186 VSUBS 0.007897f
C260 B.n187 VSUBS 0.007897f
C261 B.n188 VSUBS 0.007897f
C262 B.n189 VSUBS 0.007897f
C263 B.n190 VSUBS 0.007897f
C264 B.n191 VSUBS 0.007897f
C265 B.n192 VSUBS 0.007897f
C266 B.n193 VSUBS 0.007897f
C267 B.n194 VSUBS 0.007897f
C268 B.n195 VSUBS 0.007897f
C269 B.n196 VSUBS 0.007897f
C270 B.n197 VSUBS 0.007897f
C271 B.n198 VSUBS 0.007897f
C272 B.n199 VSUBS 0.007897f
C273 B.n200 VSUBS 0.007897f
C274 B.n201 VSUBS 0.007897f
C275 B.n202 VSUBS 0.007897f
C276 B.n203 VSUBS 0.007897f
C277 B.n204 VSUBS 0.007897f
C278 B.n205 VSUBS 0.007897f
C279 B.n206 VSUBS 0.007897f
C280 B.n207 VSUBS 0.007897f
C281 B.n208 VSUBS 0.007897f
C282 B.n209 VSUBS 0.007897f
C283 B.n210 VSUBS 0.007897f
C284 B.n211 VSUBS 0.007897f
C285 B.n212 VSUBS 0.007897f
C286 B.n213 VSUBS 0.007897f
C287 B.n214 VSUBS 0.007897f
C288 B.n215 VSUBS 0.007897f
C289 B.n216 VSUBS 0.007897f
C290 B.n217 VSUBS 0.007897f
C291 B.n218 VSUBS 0.007897f
C292 B.n219 VSUBS 0.018862f
C293 B.n220 VSUBS 0.018862f
C294 B.n221 VSUBS 0.019694f
C295 B.n222 VSUBS 0.007897f
C296 B.n223 VSUBS 0.007897f
C297 B.n224 VSUBS 0.007897f
C298 B.n225 VSUBS 0.007897f
C299 B.n226 VSUBS 0.007897f
C300 B.n227 VSUBS 0.007897f
C301 B.n228 VSUBS 0.007897f
C302 B.n229 VSUBS 0.007897f
C303 B.n230 VSUBS 0.007897f
C304 B.n231 VSUBS 0.007897f
C305 B.n232 VSUBS 0.007897f
C306 B.n233 VSUBS 0.007897f
C307 B.n234 VSUBS 0.007897f
C308 B.n235 VSUBS 0.007897f
C309 B.n236 VSUBS 0.007897f
C310 B.n237 VSUBS 0.007897f
C311 B.n238 VSUBS 0.007897f
C312 B.n239 VSUBS 0.007897f
C313 B.n240 VSUBS 0.007897f
C314 B.n241 VSUBS 0.007897f
C315 B.n242 VSUBS 0.007897f
C316 B.n243 VSUBS 0.007897f
C317 B.n244 VSUBS 0.007897f
C318 B.n245 VSUBS 0.007897f
C319 B.n246 VSUBS 0.007897f
C320 B.n247 VSUBS 0.007897f
C321 B.n248 VSUBS 0.007897f
C322 B.n249 VSUBS 0.007897f
C323 B.n250 VSUBS 0.007897f
C324 B.n251 VSUBS 0.007897f
C325 B.n252 VSUBS 0.007897f
C326 B.n253 VSUBS 0.007897f
C327 B.n254 VSUBS 0.007897f
C328 B.n255 VSUBS 0.005458f
C329 B.n256 VSUBS 0.007897f
C330 B.n257 VSUBS 0.007897f
C331 B.n258 VSUBS 0.006387f
C332 B.n259 VSUBS 0.007897f
C333 B.n260 VSUBS 0.007897f
C334 B.n261 VSUBS 0.007897f
C335 B.n262 VSUBS 0.007897f
C336 B.n263 VSUBS 0.007897f
C337 B.n264 VSUBS 0.007897f
C338 B.n265 VSUBS 0.007897f
C339 B.n266 VSUBS 0.007897f
C340 B.n267 VSUBS 0.007897f
C341 B.n268 VSUBS 0.007897f
C342 B.n269 VSUBS 0.007897f
C343 B.n270 VSUBS 0.006387f
C344 B.n271 VSUBS 0.018297f
C345 B.n272 VSUBS 0.005458f
C346 B.n273 VSUBS 0.007897f
C347 B.n274 VSUBS 0.007897f
C348 B.n275 VSUBS 0.007897f
C349 B.n276 VSUBS 0.007897f
C350 B.n277 VSUBS 0.007897f
C351 B.n278 VSUBS 0.007897f
C352 B.n279 VSUBS 0.007897f
C353 B.n280 VSUBS 0.007897f
C354 B.n281 VSUBS 0.007897f
C355 B.n282 VSUBS 0.007897f
C356 B.n283 VSUBS 0.007897f
C357 B.n284 VSUBS 0.007897f
C358 B.n285 VSUBS 0.007897f
C359 B.n286 VSUBS 0.007897f
C360 B.n287 VSUBS 0.007897f
C361 B.n288 VSUBS 0.007897f
C362 B.n289 VSUBS 0.007897f
C363 B.n290 VSUBS 0.007897f
C364 B.n291 VSUBS 0.007897f
C365 B.n292 VSUBS 0.007897f
C366 B.n293 VSUBS 0.007897f
C367 B.n294 VSUBS 0.007897f
C368 B.n295 VSUBS 0.007897f
C369 B.n296 VSUBS 0.007897f
C370 B.n297 VSUBS 0.007897f
C371 B.n298 VSUBS 0.007897f
C372 B.n299 VSUBS 0.007897f
C373 B.n300 VSUBS 0.007897f
C374 B.n301 VSUBS 0.007897f
C375 B.n302 VSUBS 0.007897f
C376 B.n303 VSUBS 0.007897f
C377 B.n304 VSUBS 0.007897f
C378 B.n305 VSUBS 0.007897f
C379 B.n306 VSUBS 0.019694f
C380 B.n307 VSUBS 0.019694f
C381 B.n308 VSUBS 0.018862f
C382 B.n309 VSUBS 0.007897f
C383 B.n310 VSUBS 0.007897f
C384 B.n311 VSUBS 0.007897f
C385 B.n312 VSUBS 0.007897f
C386 B.n313 VSUBS 0.007897f
C387 B.n314 VSUBS 0.007897f
C388 B.n315 VSUBS 0.007897f
C389 B.n316 VSUBS 0.007897f
C390 B.n317 VSUBS 0.007897f
C391 B.n318 VSUBS 0.007897f
C392 B.n319 VSUBS 0.007897f
C393 B.n320 VSUBS 0.007897f
C394 B.n321 VSUBS 0.007897f
C395 B.n322 VSUBS 0.007897f
C396 B.n323 VSUBS 0.007897f
C397 B.n324 VSUBS 0.007897f
C398 B.n325 VSUBS 0.007897f
C399 B.n326 VSUBS 0.007897f
C400 B.n327 VSUBS 0.007897f
C401 B.n328 VSUBS 0.007897f
C402 B.n329 VSUBS 0.007897f
C403 B.n330 VSUBS 0.007897f
C404 B.n331 VSUBS 0.007897f
C405 B.n332 VSUBS 0.007897f
C406 B.n333 VSUBS 0.007897f
C407 B.n334 VSUBS 0.007897f
C408 B.n335 VSUBS 0.007897f
C409 B.n336 VSUBS 0.007897f
C410 B.n337 VSUBS 0.007897f
C411 B.n338 VSUBS 0.007897f
C412 B.n339 VSUBS 0.007897f
C413 B.n340 VSUBS 0.007897f
C414 B.n341 VSUBS 0.007897f
C415 B.n342 VSUBS 0.007897f
C416 B.n343 VSUBS 0.007897f
C417 B.n344 VSUBS 0.007897f
C418 B.n345 VSUBS 0.007897f
C419 B.n346 VSUBS 0.007897f
C420 B.n347 VSUBS 0.007897f
C421 B.n348 VSUBS 0.007897f
C422 B.n349 VSUBS 0.007897f
C423 B.n350 VSUBS 0.007897f
C424 B.n351 VSUBS 0.007897f
C425 B.n352 VSUBS 0.007897f
C426 B.n353 VSUBS 0.007897f
C427 B.n354 VSUBS 0.007897f
C428 B.n355 VSUBS 0.007897f
C429 B.n356 VSUBS 0.007897f
C430 B.n357 VSUBS 0.007897f
C431 B.n358 VSUBS 0.007897f
C432 B.n359 VSUBS 0.007897f
C433 B.n360 VSUBS 0.007897f
C434 B.n361 VSUBS 0.007897f
C435 B.n362 VSUBS 0.007897f
C436 B.n363 VSUBS 0.007897f
C437 B.n364 VSUBS 0.007897f
C438 B.n365 VSUBS 0.007897f
C439 B.n366 VSUBS 0.007897f
C440 B.n367 VSUBS 0.007897f
C441 B.n368 VSUBS 0.007897f
C442 B.n369 VSUBS 0.007897f
C443 B.n370 VSUBS 0.007897f
C444 B.n371 VSUBS 0.007897f
C445 B.n372 VSUBS 0.007897f
C446 B.n373 VSUBS 0.007897f
C447 B.n374 VSUBS 0.007897f
C448 B.n375 VSUBS 0.007897f
C449 B.n376 VSUBS 0.007897f
C450 B.n377 VSUBS 0.007897f
C451 B.n378 VSUBS 0.007897f
C452 B.n379 VSUBS 0.007897f
C453 B.n380 VSUBS 0.007897f
C454 B.n381 VSUBS 0.007897f
C455 B.n382 VSUBS 0.007897f
C456 B.n383 VSUBS 0.007897f
C457 B.n384 VSUBS 0.007897f
C458 B.n385 VSUBS 0.007897f
C459 B.n386 VSUBS 0.007897f
C460 B.n387 VSUBS 0.007897f
C461 B.n388 VSUBS 0.007897f
C462 B.n389 VSUBS 0.007897f
C463 B.n390 VSUBS 0.007897f
C464 B.n391 VSUBS 0.007897f
C465 B.n392 VSUBS 0.007897f
C466 B.n393 VSUBS 0.007897f
C467 B.n394 VSUBS 0.007897f
C468 B.n395 VSUBS 0.007897f
C469 B.n396 VSUBS 0.007897f
C470 B.n397 VSUBS 0.007897f
C471 B.n398 VSUBS 0.007897f
C472 B.n399 VSUBS 0.007897f
C473 B.n400 VSUBS 0.007897f
C474 B.n401 VSUBS 0.007897f
C475 B.n402 VSUBS 0.007897f
C476 B.n403 VSUBS 0.007897f
C477 B.n404 VSUBS 0.007897f
C478 B.n405 VSUBS 0.007897f
C479 B.n406 VSUBS 0.007897f
C480 B.n407 VSUBS 0.007897f
C481 B.n408 VSUBS 0.007897f
C482 B.n409 VSUBS 0.007897f
C483 B.n410 VSUBS 0.007897f
C484 B.n411 VSUBS 0.007897f
C485 B.n412 VSUBS 0.007897f
C486 B.n413 VSUBS 0.007897f
C487 B.n414 VSUBS 0.007897f
C488 B.n415 VSUBS 0.007897f
C489 B.n416 VSUBS 0.007897f
C490 B.n417 VSUBS 0.007897f
C491 B.n418 VSUBS 0.007897f
C492 B.n419 VSUBS 0.007897f
C493 B.n420 VSUBS 0.007897f
C494 B.n421 VSUBS 0.007897f
C495 B.n422 VSUBS 0.007897f
C496 B.n423 VSUBS 0.007897f
C497 B.n424 VSUBS 0.007897f
C498 B.n425 VSUBS 0.007897f
C499 B.n426 VSUBS 0.007897f
C500 B.n427 VSUBS 0.007897f
C501 B.n428 VSUBS 0.007897f
C502 B.n429 VSUBS 0.007897f
C503 B.n430 VSUBS 0.007897f
C504 B.n431 VSUBS 0.007897f
C505 B.n432 VSUBS 0.007897f
C506 B.n433 VSUBS 0.007897f
C507 B.n434 VSUBS 0.007897f
C508 B.n435 VSUBS 0.007897f
C509 B.n436 VSUBS 0.007897f
C510 B.n437 VSUBS 0.007897f
C511 B.n438 VSUBS 0.007897f
C512 B.n439 VSUBS 0.007897f
C513 B.n440 VSUBS 0.019737f
C514 B.n441 VSUBS 0.018819f
C515 B.n442 VSUBS 0.019694f
C516 B.n443 VSUBS 0.007897f
C517 B.n444 VSUBS 0.007897f
C518 B.n445 VSUBS 0.007897f
C519 B.n446 VSUBS 0.007897f
C520 B.n447 VSUBS 0.007897f
C521 B.n448 VSUBS 0.007897f
C522 B.n449 VSUBS 0.007897f
C523 B.n450 VSUBS 0.007897f
C524 B.n451 VSUBS 0.007897f
C525 B.n452 VSUBS 0.007897f
C526 B.n453 VSUBS 0.007897f
C527 B.n454 VSUBS 0.007897f
C528 B.n455 VSUBS 0.007897f
C529 B.n456 VSUBS 0.007897f
C530 B.n457 VSUBS 0.007897f
C531 B.n458 VSUBS 0.007897f
C532 B.n459 VSUBS 0.007897f
C533 B.n460 VSUBS 0.007897f
C534 B.n461 VSUBS 0.007897f
C535 B.n462 VSUBS 0.007897f
C536 B.n463 VSUBS 0.007897f
C537 B.n464 VSUBS 0.007897f
C538 B.n465 VSUBS 0.007897f
C539 B.n466 VSUBS 0.007897f
C540 B.n467 VSUBS 0.007897f
C541 B.n468 VSUBS 0.007897f
C542 B.n469 VSUBS 0.007897f
C543 B.n470 VSUBS 0.007897f
C544 B.n471 VSUBS 0.007897f
C545 B.n472 VSUBS 0.007897f
C546 B.n473 VSUBS 0.007897f
C547 B.n474 VSUBS 0.007897f
C548 B.n475 VSUBS 0.007897f
C549 B.n476 VSUBS 0.005458f
C550 B.n477 VSUBS 0.018297f
C551 B.n478 VSUBS 0.006387f
C552 B.n479 VSUBS 0.007897f
C553 B.n480 VSUBS 0.007897f
C554 B.n481 VSUBS 0.007897f
C555 B.n482 VSUBS 0.007897f
C556 B.n483 VSUBS 0.007897f
C557 B.n484 VSUBS 0.007897f
C558 B.n485 VSUBS 0.007897f
C559 B.n486 VSUBS 0.007897f
C560 B.n487 VSUBS 0.007897f
C561 B.n488 VSUBS 0.007897f
C562 B.n489 VSUBS 0.007897f
C563 B.n490 VSUBS 0.006387f
C564 B.n491 VSUBS 0.007897f
C565 B.n492 VSUBS 0.007897f
C566 B.n493 VSUBS 0.005458f
C567 B.n494 VSUBS 0.007897f
C568 B.n495 VSUBS 0.007897f
C569 B.n496 VSUBS 0.007897f
C570 B.n497 VSUBS 0.007897f
C571 B.n498 VSUBS 0.007897f
C572 B.n499 VSUBS 0.007897f
C573 B.n500 VSUBS 0.007897f
C574 B.n501 VSUBS 0.007897f
C575 B.n502 VSUBS 0.007897f
C576 B.n503 VSUBS 0.007897f
C577 B.n504 VSUBS 0.007897f
C578 B.n505 VSUBS 0.007897f
C579 B.n506 VSUBS 0.007897f
C580 B.n507 VSUBS 0.007897f
C581 B.n508 VSUBS 0.007897f
C582 B.n509 VSUBS 0.007897f
C583 B.n510 VSUBS 0.007897f
C584 B.n511 VSUBS 0.007897f
C585 B.n512 VSUBS 0.007897f
C586 B.n513 VSUBS 0.007897f
C587 B.n514 VSUBS 0.007897f
C588 B.n515 VSUBS 0.007897f
C589 B.n516 VSUBS 0.007897f
C590 B.n517 VSUBS 0.007897f
C591 B.n518 VSUBS 0.007897f
C592 B.n519 VSUBS 0.007897f
C593 B.n520 VSUBS 0.007897f
C594 B.n521 VSUBS 0.007897f
C595 B.n522 VSUBS 0.007897f
C596 B.n523 VSUBS 0.007897f
C597 B.n524 VSUBS 0.007897f
C598 B.n525 VSUBS 0.007897f
C599 B.n526 VSUBS 0.007897f
C600 B.n527 VSUBS 0.019694f
C601 B.n528 VSUBS 0.018862f
C602 B.n529 VSUBS 0.018862f
C603 B.n530 VSUBS 0.007897f
C604 B.n531 VSUBS 0.007897f
C605 B.n532 VSUBS 0.007897f
C606 B.n533 VSUBS 0.007897f
C607 B.n534 VSUBS 0.007897f
C608 B.n535 VSUBS 0.007897f
C609 B.n536 VSUBS 0.007897f
C610 B.n537 VSUBS 0.007897f
C611 B.n538 VSUBS 0.007897f
C612 B.n539 VSUBS 0.007897f
C613 B.n540 VSUBS 0.007897f
C614 B.n541 VSUBS 0.007897f
C615 B.n542 VSUBS 0.007897f
C616 B.n543 VSUBS 0.007897f
C617 B.n544 VSUBS 0.007897f
C618 B.n545 VSUBS 0.007897f
C619 B.n546 VSUBS 0.007897f
C620 B.n547 VSUBS 0.007897f
C621 B.n548 VSUBS 0.007897f
C622 B.n549 VSUBS 0.007897f
C623 B.n550 VSUBS 0.007897f
C624 B.n551 VSUBS 0.007897f
C625 B.n552 VSUBS 0.007897f
C626 B.n553 VSUBS 0.007897f
C627 B.n554 VSUBS 0.007897f
C628 B.n555 VSUBS 0.007897f
C629 B.n556 VSUBS 0.007897f
C630 B.n557 VSUBS 0.007897f
C631 B.n558 VSUBS 0.007897f
C632 B.n559 VSUBS 0.007897f
C633 B.n560 VSUBS 0.007897f
C634 B.n561 VSUBS 0.007897f
C635 B.n562 VSUBS 0.007897f
C636 B.n563 VSUBS 0.007897f
C637 B.n564 VSUBS 0.007897f
C638 B.n565 VSUBS 0.007897f
C639 B.n566 VSUBS 0.007897f
C640 B.n567 VSUBS 0.007897f
C641 B.n568 VSUBS 0.007897f
C642 B.n569 VSUBS 0.007897f
C643 B.n570 VSUBS 0.007897f
C644 B.n571 VSUBS 0.007897f
C645 B.n572 VSUBS 0.007897f
C646 B.n573 VSUBS 0.007897f
C647 B.n574 VSUBS 0.007897f
C648 B.n575 VSUBS 0.007897f
C649 B.n576 VSUBS 0.007897f
C650 B.n577 VSUBS 0.007897f
C651 B.n578 VSUBS 0.007897f
C652 B.n579 VSUBS 0.007897f
C653 B.n580 VSUBS 0.007897f
C654 B.n581 VSUBS 0.007897f
C655 B.n582 VSUBS 0.007897f
C656 B.n583 VSUBS 0.007897f
C657 B.n584 VSUBS 0.007897f
C658 B.n585 VSUBS 0.007897f
C659 B.n586 VSUBS 0.007897f
C660 B.n587 VSUBS 0.007897f
C661 B.n588 VSUBS 0.007897f
C662 B.n589 VSUBS 0.007897f
C663 B.n590 VSUBS 0.007897f
C664 B.n591 VSUBS 0.007897f
C665 B.n592 VSUBS 0.007897f
C666 B.n593 VSUBS 0.007897f
C667 B.n594 VSUBS 0.007897f
C668 B.n595 VSUBS 0.017882f
C669 VTAIL.n0 VSUBS 0.03136f
C670 VTAIL.n1 VSUBS 0.029216f
C671 VTAIL.n2 VSUBS 0.015699f
C672 VTAIL.n3 VSUBS 0.037107f
C673 VTAIL.n4 VSUBS 0.016623f
C674 VTAIL.n5 VSUBS 0.029216f
C675 VTAIL.n6 VSUBS 0.015699f
C676 VTAIL.n7 VSUBS 0.037107f
C677 VTAIL.n8 VSUBS 0.016623f
C678 VTAIL.n9 VSUBS 0.128667f
C679 VTAIL.t7 VSUBS 0.07954f
C680 VTAIL.n10 VSUBS 0.02783f
C681 VTAIL.n11 VSUBS 0.023593f
C682 VTAIL.n12 VSUBS 0.015699f
C683 VTAIL.n13 VSUBS 0.663714f
C684 VTAIL.n14 VSUBS 0.029216f
C685 VTAIL.n15 VSUBS 0.015699f
C686 VTAIL.n16 VSUBS 0.016623f
C687 VTAIL.n17 VSUBS 0.037107f
C688 VTAIL.n18 VSUBS 0.037107f
C689 VTAIL.n19 VSUBS 0.016623f
C690 VTAIL.n20 VSUBS 0.015699f
C691 VTAIL.n21 VSUBS 0.029216f
C692 VTAIL.n22 VSUBS 0.029216f
C693 VTAIL.n23 VSUBS 0.015699f
C694 VTAIL.n24 VSUBS 0.016623f
C695 VTAIL.n25 VSUBS 0.037107f
C696 VTAIL.n26 VSUBS 0.087307f
C697 VTAIL.n27 VSUBS 0.016623f
C698 VTAIL.n28 VSUBS 0.015699f
C699 VTAIL.n29 VSUBS 0.065535f
C700 VTAIL.n30 VSUBS 0.043732f
C701 VTAIL.n31 VSUBS 0.23909f
C702 VTAIL.n32 VSUBS 0.03136f
C703 VTAIL.n33 VSUBS 0.029216f
C704 VTAIL.n34 VSUBS 0.015699f
C705 VTAIL.n35 VSUBS 0.037107f
C706 VTAIL.n36 VSUBS 0.016623f
C707 VTAIL.n37 VSUBS 0.029216f
C708 VTAIL.n38 VSUBS 0.015699f
C709 VTAIL.n39 VSUBS 0.037107f
C710 VTAIL.n40 VSUBS 0.016623f
C711 VTAIL.n41 VSUBS 0.128667f
C712 VTAIL.t0 VSUBS 0.07954f
C713 VTAIL.n42 VSUBS 0.02783f
C714 VTAIL.n43 VSUBS 0.023593f
C715 VTAIL.n44 VSUBS 0.015699f
C716 VTAIL.n45 VSUBS 0.663714f
C717 VTAIL.n46 VSUBS 0.029216f
C718 VTAIL.n47 VSUBS 0.015699f
C719 VTAIL.n48 VSUBS 0.016623f
C720 VTAIL.n49 VSUBS 0.037107f
C721 VTAIL.n50 VSUBS 0.037107f
C722 VTAIL.n51 VSUBS 0.016623f
C723 VTAIL.n52 VSUBS 0.015699f
C724 VTAIL.n53 VSUBS 0.029216f
C725 VTAIL.n54 VSUBS 0.029216f
C726 VTAIL.n55 VSUBS 0.015699f
C727 VTAIL.n56 VSUBS 0.016623f
C728 VTAIL.n57 VSUBS 0.037107f
C729 VTAIL.n58 VSUBS 0.087307f
C730 VTAIL.n59 VSUBS 0.016623f
C731 VTAIL.n60 VSUBS 0.015699f
C732 VTAIL.n61 VSUBS 0.065535f
C733 VTAIL.n62 VSUBS 0.043732f
C734 VTAIL.n63 VSUBS 0.399168f
C735 VTAIL.n64 VSUBS 0.03136f
C736 VTAIL.n65 VSUBS 0.029216f
C737 VTAIL.n66 VSUBS 0.015699f
C738 VTAIL.n67 VSUBS 0.037107f
C739 VTAIL.n68 VSUBS 0.016623f
C740 VTAIL.n69 VSUBS 0.029216f
C741 VTAIL.n70 VSUBS 0.015699f
C742 VTAIL.n71 VSUBS 0.037107f
C743 VTAIL.n72 VSUBS 0.016623f
C744 VTAIL.n73 VSUBS 0.128667f
C745 VTAIL.t1 VSUBS 0.07954f
C746 VTAIL.n74 VSUBS 0.02783f
C747 VTAIL.n75 VSUBS 0.023593f
C748 VTAIL.n76 VSUBS 0.015699f
C749 VTAIL.n77 VSUBS 0.663714f
C750 VTAIL.n78 VSUBS 0.029216f
C751 VTAIL.n79 VSUBS 0.015699f
C752 VTAIL.n80 VSUBS 0.016623f
C753 VTAIL.n81 VSUBS 0.037107f
C754 VTAIL.n82 VSUBS 0.037107f
C755 VTAIL.n83 VSUBS 0.016623f
C756 VTAIL.n84 VSUBS 0.015699f
C757 VTAIL.n85 VSUBS 0.029216f
C758 VTAIL.n86 VSUBS 0.029216f
C759 VTAIL.n87 VSUBS 0.015699f
C760 VTAIL.n88 VSUBS 0.016623f
C761 VTAIL.n89 VSUBS 0.037107f
C762 VTAIL.n90 VSUBS 0.087307f
C763 VTAIL.n91 VSUBS 0.016623f
C764 VTAIL.n92 VSUBS 0.015699f
C765 VTAIL.n93 VSUBS 0.065535f
C766 VTAIL.n94 VSUBS 0.043732f
C767 VTAIL.n95 VSUBS 1.56578f
C768 VTAIL.n96 VSUBS 0.03136f
C769 VTAIL.n97 VSUBS 0.029216f
C770 VTAIL.n98 VSUBS 0.015699f
C771 VTAIL.n99 VSUBS 0.037107f
C772 VTAIL.n100 VSUBS 0.016623f
C773 VTAIL.n101 VSUBS 0.029216f
C774 VTAIL.n102 VSUBS 0.015699f
C775 VTAIL.n103 VSUBS 0.037107f
C776 VTAIL.n104 VSUBS 0.016623f
C777 VTAIL.n105 VSUBS 0.128667f
C778 VTAIL.t4 VSUBS 0.07954f
C779 VTAIL.n106 VSUBS 0.02783f
C780 VTAIL.n107 VSUBS 0.023593f
C781 VTAIL.n108 VSUBS 0.015699f
C782 VTAIL.n109 VSUBS 0.663714f
C783 VTAIL.n110 VSUBS 0.029216f
C784 VTAIL.n111 VSUBS 0.015699f
C785 VTAIL.n112 VSUBS 0.016623f
C786 VTAIL.n113 VSUBS 0.037107f
C787 VTAIL.n114 VSUBS 0.037107f
C788 VTAIL.n115 VSUBS 0.016623f
C789 VTAIL.n116 VSUBS 0.015699f
C790 VTAIL.n117 VSUBS 0.029216f
C791 VTAIL.n118 VSUBS 0.029216f
C792 VTAIL.n119 VSUBS 0.015699f
C793 VTAIL.n120 VSUBS 0.016623f
C794 VTAIL.n121 VSUBS 0.037107f
C795 VTAIL.n122 VSUBS 0.087307f
C796 VTAIL.n123 VSUBS 0.016623f
C797 VTAIL.n124 VSUBS 0.015699f
C798 VTAIL.n125 VSUBS 0.065535f
C799 VTAIL.n126 VSUBS 0.043732f
C800 VTAIL.n127 VSUBS 1.56578f
C801 VTAIL.n128 VSUBS 0.03136f
C802 VTAIL.n129 VSUBS 0.029216f
C803 VTAIL.n130 VSUBS 0.015699f
C804 VTAIL.n131 VSUBS 0.037107f
C805 VTAIL.n132 VSUBS 0.016623f
C806 VTAIL.n133 VSUBS 0.029216f
C807 VTAIL.n134 VSUBS 0.015699f
C808 VTAIL.n135 VSUBS 0.037107f
C809 VTAIL.n136 VSUBS 0.016623f
C810 VTAIL.n137 VSUBS 0.128667f
C811 VTAIL.t6 VSUBS 0.07954f
C812 VTAIL.n138 VSUBS 0.02783f
C813 VTAIL.n139 VSUBS 0.023593f
C814 VTAIL.n140 VSUBS 0.015699f
C815 VTAIL.n141 VSUBS 0.663714f
C816 VTAIL.n142 VSUBS 0.029216f
C817 VTAIL.n143 VSUBS 0.015699f
C818 VTAIL.n144 VSUBS 0.016623f
C819 VTAIL.n145 VSUBS 0.037107f
C820 VTAIL.n146 VSUBS 0.037107f
C821 VTAIL.n147 VSUBS 0.016623f
C822 VTAIL.n148 VSUBS 0.015699f
C823 VTAIL.n149 VSUBS 0.029216f
C824 VTAIL.n150 VSUBS 0.029216f
C825 VTAIL.n151 VSUBS 0.015699f
C826 VTAIL.n152 VSUBS 0.016623f
C827 VTAIL.n153 VSUBS 0.037107f
C828 VTAIL.n154 VSUBS 0.087307f
C829 VTAIL.n155 VSUBS 0.016623f
C830 VTAIL.n156 VSUBS 0.015699f
C831 VTAIL.n157 VSUBS 0.065535f
C832 VTAIL.n158 VSUBS 0.043732f
C833 VTAIL.n159 VSUBS 0.399168f
C834 VTAIL.n160 VSUBS 0.03136f
C835 VTAIL.n161 VSUBS 0.029216f
C836 VTAIL.n162 VSUBS 0.015699f
C837 VTAIL.n163 VSUBS 0.037107f
C838 VTAIL.n164 VSUBS 0.016623f
C839 VTAIL.n165 VSUBS 0.029216f
C840 VTAIL.n166 VSUBS 0.015699f
C841 VTAIL.n167 VSUBS 0.037107f
C842 VTAIL.n168 VSUBS 0.016623f
C843 VTAIL.n169 VSUBS 0.128667f
C844 VTAIL.t2 VSUBS 0.07954f
C845 VTAIL.n170 VSUBS 0.02783f
C846 VTAIL.n171 VSUBS 0.023593f
C847 VTAIL.n172 VSUBS 0.015699f
C848 VTAIL.n173 VSUBS 0.663714f
C849 VTAIL.n174 VSUBS 0.029216f
C850 VTAIL.n175 VSUBS 0.015699f
C851 VTAIL.n176 VSUBS 0.016623f
C852 VTAIL.n177 VSUBS 0.037107f
C853 VTAIL.n178 VSUBS 0.037107f
C854 VTAIL.n179 VSUBS 0.016623f
C855 VTAIL.n180 VSUBS 0.015699f
C856 VTAIL.n181 VSUBS 0.029216f
C857 VTAIL.n182 VSUBS 0.029216f
C858 VTAIL.n183 VSUBS 0.015699f
C859 VTAIL.n184 VSUBS 0.016623f
C860 VTAIL.n185 VSUBS 0.037107f
C861 VTAIL.n186 VSUBS 0.087307f
C862 VTAIL.n187 VSUBS 0.016623f
C863 VTAIL.n188 VSUBS 0.015699f
C864 VTAIL.n189 VSUBS 0.065535f
C865 VTAIL.n190 VSUBS 0.043732f
C866 VTAIL.n191 VSUBS 0.399168f
C867 VTAIL.n192 VSUBS 0.03136f
C868 VTAIL.n193 VSUBS 0.029216f
C869 VTAIL.n194 VSUBS 0.015699f
C870 VTAIL.n195 VSUBS 0.037107f
C871 VTAIL.n196 VSUBS 0.016623f
C872 VTAIL.n197 VSUBS 0.029216f
C873 VTAIL.n198 VSUBS 0.015699f
C874 VTAIL.n199 VSUBS 0.037107f
C875 VTAIL.n200 VSUBS 0.016623f
C876 VTAIL.n201 VSUBS 0.128667f
C877 VTAIL.t3 VSUBS 0.07954f
C878 VTAIL.n202 VSUBS 0.02783f
C879 VTAIL.n203 VSUBS 0.023593f
C880 VTAIL.n204 VSUBS 0.015699f
C881 VTAIL.n205 VSUBS 0.663714f
C882 VTAIL.n206 VSUBS 0.029216f
C883 VTAIL.n207 VSUBS 0.015699f
C884 VTAIL.n208 VSUBS 0.016623f
C885 VTAIL.n209 VSUBS 0.037107f
C886 VTAIL.n210 VSUBS 0.037107f
C887 VTAIL.n211 VSUBS 0.016623f
C888 VTAIL.n212 VSUBS 0.015699f
C889 VTAIL.n213 VSUBS 0.029216f
C890 VTAIL.n214 VSUBS 0.029216f
C891 VTAIL.n215 VSUBS 0.015699f
C892 VTAIL.n216 VSUBS 0.016623f
C893 VTAIL.n217 VSUBS 0.037107f
C894 VTAIL.n218 VSUBS 0.087307f
C895 VTAIL.n219 VSUBS 0.016623f
C896 VTAIL.n220 VSUBS 0.015699f
C897 VTAIL.n221 VSUBS 0.065535f
C898 VTAIL.n222 VSUBS 0.043732f
C899 VTAIL.n223 VSUBS 1.56578f
C900 VTAIL.n224 VSUBS 0.03136f
C901 VTAIL.n225 VSUBS 0.029216f
C902 VTAIL.n226 VSUBS 0.015699f
C903 VTAIL.n227 VSUBS 0.037107f
C904 VTAIL.n228 VSUBS 0.016623f
C905 VTAIL.n229 VSUBS 0.029216f
C906 VTAIL.n230 VSUBS 0.015699f
C907 VTAIL.n231 VSUBS 0.037107f
C908 VTAIL.n232 VSUBS 0.016623f
C909 VTAIL.n233 VSUBS 0.128667f
C910 VTAIL.t5 VSUBS 0.07954f
C911 VTAIL.n234 VSUBS 0.02783f
C912 VTAIL.n235 VSUBS 0.023593f
C913 VTAIL.n236 VSUBS 0.015699f
C914 VTAIL.n237 VSUBS 0.663714f
C915 VTAIL.n238 VSUBS 0.029216f
C916 VTAIL.n239 VSUBS 0.015699f
C917 VTAIL.n240 VSUBS 0.016623f
C918 VTAIL.n241 VSUBS 0.037107f
C919 VTAIL.n242 VSUBS 0.037107f
C920 VTAIL.n243 VSUBS 0.016623f
C921 VTAIL.n244 VSUBS 0.015699f
C922 VTAIL.n245 VSUBS 0.029216f
C923 VTAIL.n246 VSUBS 0.029216f
C924 VTAIL.n247 VSUBS 0.015699f
C925 VTAIL.n248 VSUBS 0.016623f
C926 VTAIL.n249 VSUBS 0.037107f
C927 VTAIL.n250 VSUBS 0.087307f
C928 VTAIL.n251 VSUBS 0.016623f
C929 VTAIL.n252 VSUBS 0.015699f
C930 VTAIL.n253 VSUBS 0.065535f
C931 VTAIL.n254 VSUBS 0.043732f
C932 VTAIL.n255 VSUBS 1.39475f
C933 VDD2.t0 VSUBS 0.133938f
C934 VDD2.t3 VSUBS 0.133938f
C935 VDD2.n0 VSUBS 1.38322f
C936 VDD2.t1 VSUBS 0.133938f
C937 VDD2.t2 VSUBS 0.133938f
C938 VDD2.n1 VSUBS 0.883619f
C939 VDD2.n2 VSUBS 4.06843f
C940 VN.t2 VSUBS 2.56882f
C941 VN.t0 VSUBS 2.58808f
C942 VN.n0 VSUBS 1.53667f
C943 VN.t3 VSUBS 2.56882f
C944 VN.t1 VSUBS 2.58808f
C945 VN.n1 VSUBS 3.59327f
.ends

