* NGSPICE file created from diff_pair_sample_0978.ext - technology: sky130A

.subckt diff_pair_sample_0978 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=7.7649 ps=40.6 w=19.91 l=0.29
X1 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=7.7649 ps=40.6 w=19.91 l=0.29
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=0 ps=0 w=19.91 l=0.29
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=0 ps=0 w=19.91 l=0.29
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=7.7649 ps=40.6 w=19.91 l=0.29
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=0 ps=0 w=19.91 l=0.29
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=0 ps=0 w=19.91 l=0.29
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7649 pd=40.6 as=7.7649 ps=40.6 w=19.91 l=0.29
R0 VN VN.t0 1993.77
R1 VN VN.t1 1948.91
R2 VTAIL.n1 VTAIL.t2 48.9811
R3 VTAIL.n3 VTAIL.t3 48.9809
R4 VTAIL.n0 VTAIL.t0 48.9809
R5 VTAIL.n2 VTAIL.t1 48.9809
R6 VTAIL.n1 VTAIL.n0 30.6169
R7 VTAIL.n3 VTAIL.n2 30.0824
R8 VTAIL.n2 VTAIL.n1 0.737569
R9 VTAIL VTAIL.n0 0.662138
R10 VTAIL VTAIL.n3 0.075931
R11 VDD2.n0 VDD2.t0 107.57
R12 VDD2.n0 VDD2.t1 65.6597
R13 VDD2 VDD2.n0 0.19231
R14 B.n100 B.t6 1872.24
R15 B.n97 B.t2 1872.24
R16 B.n467 B.t13 1872.24
R17 B.n464 B.t9 1872.24
R18 B.n797 B.n796 585
R19 B.n798 B.n797 585
R20 B.n373 B.n95 585
R21 B.n372 B.n371 585
R22 B.n370 B.n369 585
R23 B.n368 B.n367 585
R24 B.n366 B.n365 585
R25 B.n364 B.n363 585
R26 B.n362 B.n361 585
R27 B.n360 B.n359 585
R28 B.n358 B.n357 585
R29 B.n356 B.n355 585
R30 B.n354 B.n353 585
R31 B.n352 B.n351 585
R32 B.n350 B.n349 585
R33 B.n348 B.n347 585
R34 B.n346 B.n345 585
R35 B.n344 B.n343 585
R36 B.n342 B.n341 585
R37 B.n340 B.n339 585
R38 B.n338 B.n337 585
R39 B.n336 B.n335 585
R40 B.n334 B.n333 585
R41 B.n332 B.n331 585
R42 B.n330 B.n329 585
R43 B.n328 B.n327 585
R44 B.n326 B.n325 585
R45 B.n324 B.n323 585
R46 B.n322 B.n321 585
R47 B.n320 B.n319 585
R48 B.n318 B.n317 585
R49 B.n316 B.n315 585
R50 B.n314 B.n313 585
R51 B.n312 B.n311 585
R52 B.n310 B.n309 585
R53 B.n308 B.n307 585
R54 B.n306 B.n305 585
R55 B.n304 B.n303 585
R56 B.n302 B.n301 585
R57 B.n300 B.n299 585
R58 B.n298 B.n297 585
R59 B.n296 B.n295 585
R60 B.n294 B.n293 585
R61 B.n292 B.n291 585
R62 B.n290 B.n289 585
R63 B.n288 B.n287 585
R64 B.n286 B.n285 585
R65 B.n284 B.n283 585
R66 B.n282 B.n281 585
R67 B.n280 B.n279 585
R68 B.n278 B.n277 585
R69 B.n276 B.n275 585
R70 B.n274 B.n273 585
R71 B.n272 B.n271 585
R72 B.n270 B.n269 585
R73 B.n268 B.n267 585
R74 B.n266 B.n265 585
R75 B.n264 B.n263 585
R76 B.n262 B.n261 585
R77 B.n260 B.n259 585
R78 B.n258 B.n257 585
R79 B.n256 B.n255 585
R80 B.n254 B.n253 585
R81 B.n252 B.n251 585
R82 B.n250 B.n249 585
R83 B.n248 B.n247 585
R84 B.n246 B.n245 585
R85 B.n244 B.n243 585
R86 B.n242 B.n241 585
R87 B.n240 B.n239 585
R88 B.n238 B.n237 585
R89 B.n236 B.n235 585
R90 B.n234 B.n233 585
R91 B.n232 B.n231 585
R92 B.n230 B.n229 585
R93 B.n227 B.n226 585
R94 B.n225 B.n224 585
R95 B.n223 B.n222 585
R96 B.n221 B.n220 585
R97 B.n219 B.n218 585
R98 B.n217 B.n216 585
R99 B.n215 B.n214 585
R100 B.n213 B.n212 585
R101 B.n211 B.n210 585
R102 B.n209 B.n208 585
R103 B.n207 B.n206 585
R104 B.n205 B.n204 585
R105 B.n203 B.n202 585
R106 B.n201 B.n200 585
R107 B.n199 B.n198 585
R108 B.n197 B.n196 585
R109 B.n195 B.n194 585
R110 B.n193 B.n192 585
R111 B.n191 B.n190 585
R112 B.n189 B.n188 585
R113 B.n187 B.n186 585
R114 B.n185 B.n184 585
R115 B.n183 B.n182 585
R116 B.n181 B.n180 585
R117 B.n179 B.n178 585
R118 B.n177 B.n176 585
R119 B.n175 B.n174 585
R120 B.n173 B.n172 585
R121 B.n171 B.n170 585
R122 B.n169 B.n168 585
R123 B.n167 B.n166 585
R124 B.n165 B.n164 585
R125 B.n163 B.n162 585
R126 B.n161 B.n160 585
R127 B.n159 B.n158 585
R128 B.n157 B.n156 585
R129 B.n155 B.n154 585
R130 B.n153 B.n152 585
R131 B.n151 B.n150 585
R132 B.n149 B.n148 585
R133 B.n147 B.n146 585
R134 B.n145 B.n144 585
R135 B.n143 B.n142 585
R136 B.n141 B.n140 585
R137 B.n139 B.n138 585
R138 B.n137 B.n136 585
R139 B.n135 B.n134 585
R140 B.n133 B.n132 585
R141 B.n131 B.n130 585
R142 B.n129 B.n128 585
R143 B.n127 B.n126 585
R144 B.n125 B.n124 585
R145 B.n123 B.n122 585
R146 B.n121 B.n120 585
R147 B.n119 B.n118 585
R148 B.n117 B.n116 585
R149 B.n115 B.n114 585
R150 B.n113 B.n112 585
R151 B.n111 B.n110 585
R152 B.n109 B.n108 585
R153 B.n107 B.n106 585
R154 B.n105 B.n104 585
R155 B.n103 B.n102 585
R156 B.n26 B.n25 585
R157 B.n801 B.n800 585
R158 B.n795 B.n96 585
R159 B.n96 B.n23 585
R160 B.n794 B.n22 585
R161 B.n805 B.n22 585
R162 B.n793 B.n21 585
R163 B.n806 B.n21 585
R164 B.n792 B.n20 585
R165 B.n807 B.n20 585
R166 B.n791 B.n790 585
R167 B.n790 B.n16 585
R168 B.n789 B.n15 585
R169 B.n813 B.n15 585
R170 B.n788 B.n14 585
R171 B.n814 B.n14 585
R172 B.n787 B.n13 585
R173 B.n815 B.n13 585
R174 B.n786 B.n785 585
R175 B.n785 B.n12 585
R176 B.n784 B.n783 585
R177 B.n784 B.n8 585
R178 B.n782 B.n7 585
R179 B.n822 B.n7 585
R180 B.n781 B.n6 585
R181 B.n823 B.n6 585
R182 B.n780 B.n5 585
R183 B.n824 B.n5 585
R184 B.n779 B.n778 585
R185 B.n778 B.n4 585
R186 B.n777 B.n374 585
R187 B.n777 B.n776 585
R188 B.n766 B.n375 585
R189 B.n769 B.n375 585
R190 B.n768 B.n767 585
R191 B.n770 B.n768 585
R192 B.n765 B.n380 585
R193 B.n380 B.n379 585
R194 B.n764 B.n763 585
R195 B.n763 B.n762 585
R196 B.n382 B.n381 585
R197 B.n383 B.n382 585
R198 B.n755 B.n754 585
R199 B.n756 B.n755 585
R200 B.n753 B.n388 585
R201 B.n388 B.n387 585
R202 B.n752 B.n751 585
R203 B.n751 B.n750 585
R204 B.n390 B.n389 585
R205 B.n391 B.n390 585
R206 B.n746 B.n745 585
R207 B.n394 B.n393 585
R208 B.n742 B.n741 585
R209 B.n743 B.n742 585
R210 B.n740 B.n463 585
R211 B.n739 B.n738 585
R212 B.n737 B.n736 585
R213 B.n735 B.n734 585
R214 B.n733 B.n732 585
R215 B.n731 B.n730 585
R216 B.n729 B.n728 585
R217 B.n727 B.n726 585
R218 B.n725 B.n724 585
R219 B.n723 B.n722 585
R220 B.n721 B.n720 585
R221 B.n719 B.n718 585
R222 B.n717 B.n716 585
R223 B.n715 B.n714 585
R224 B.n713 B.n712 585
R225 B.n711 B.n710 585
R226 B.n709 B.n708 585
R227 B.n707 B.n706 585
R228 B.n705 B.n704 585
R229 B.n703 B.n702 585
R230 B.n701 B.n700 585
R231 B.n699 B.n698 585
R232 B.n697 B.n696 585
R233 B.n695 B.n694 585
R234 B.n693 B.n692 585
R235 B.n691 B.n690 585
R236 B.n689 B.n688 585
R237 B.n687 B.n686 585
R238 B.n685 B.n684 585
R239 B.n683 B.n682 585
R240 B.n681 B.n680 585
R241 B.n679 B.n678 585
R242 B.n677 B.n676 585
R243 B.n675 B.n674 585
R244 B.n673 B.n672 585
R245 B.n671 B.n670 585
R246 B.n669 B.n668 585
R247 B.n667 B.n666 585
R248 B.n665 B.n664 585
R249 B.n663 B.n662 585
R250 B.n661 B.n660 585
R251 B.n659 B.n658 585
R252 B.n657 B.n656 585
R253 B.n655 B.n654 585
R254 B.n653 B.n652 585
R255 B.n651 B.n650 585
R256 B.n649 B.n648 585
R257 B.n647 B.n646 585
R258 B.n645 B.n644 585
R259 B.n643 B.n642 585
R260 B.n641 B.n640 585
R261 B.n639 B.n638 585
R262 B.n637 B.n636 585
R263 B.n635 B.n634 585
R264 B.n633 B.n632 585
R265 B.n631 B.n630 585
R266 B.n629 B.n628 585
R267 B.n627 B.n626 585
R268 B.n625 B.n624 585
R269 B.n623 B.n622 585
R270 B.n621 B.n620 585
R271 B.n619 B.n618 585
R272 B.n617 B.n616 585
R273 B.n615 B.n614 585
R274 B.n613 B.n612 585
R275 B.n611 B.n610 585
R276 B.n609 B.n608 585
R277 B.n607 B.n606 585
R278 B.n605 B.n604 585
R279 B.n603 B.n602 585
R280 B.n601 B.n600 585
R281 B.n598 B.n597 585
R282 B.n596 B.n595 585
R283 B.n594 B.n593 585
R284 B.n592 B.n591 585
R285 B.n590 B.n589 585
R286 B.n588 B.n587 585
R287 B.n586 B.n585 585
R288 B.n584 B.n583 585
R289 B.n582 B.n581 585
R290 B.n580 B.n579 585
R291 B.n578 B.n577 585
R292 B.n576 B.n575 585
R293 B.n574 B.n573 585
R294 B.n572 B.n571 585
R295 B.n570 B.n569 585
R296 B.n568 B.n567 585
R297 B.n566 B.n565 585
R298 B.n564 B.n563 585
R299 B.n562 B.n561 585
R300 B.n560 B.n559 585
R301 B.n558 B.n557 585
R302 B.n556 B.n555 585
R303 B.n554 B.n553 585
R304 B.n552 B.n551 585
R305 B.n550 B.n549 585
R306 B.n548 B.n547 585
R307 B.n546 B.n545 585
R308 B.n544 B.n543 585
R309 B.n542 B.n541 585
R310 B.n540 B.n539 585
R311 B.n538 B.n537 585
R312 B.n536 B.n535 585
R313 B.n534 B.n533 585
R314 B.n532 B.n531 585
R315 B.n530 B.n529 585
R316 B.n528 B.n527 585
R317 B.n526 B.n525 585
R318 B.n524 B.n523 585
R319 B.n522 B.n521 585
R320 B.n520 B.n519 585
R321 B.n518 B.n517 585
R322 B.n516 B.n515 585
R323 B.n514 B.n513 585
R324 B.n512 B.n511 585
R325 B.n510 B.n509 585
R326 B.n508 B.n507 585
R327 B.n506 B.n505 585
R328 B.n504 B.n503 585
R329 B.n502 B.n501 585
R330 B.n500 B.n499 585
R331 B.n498 B.n497 585
R332 B.n496 B.n495 585
R333 B.n494 B.n493 585
R334 B.n492 B.n491 585
R335 B.n490 B.n489 585
R336 B.n488 B.n487 585
R337 B.n486 B.n485 585
R338 B.n484 B.n483 585
R339 B.n482 B.n481 585
R340 B.n480 B.n479 585
R341 B.n478 B.n477 585
R342 B.n476 B.n475 585
R343 B.n474 B.n473 585
R344 B.n472 B.n471 585
R345 B.n470 B.n469 585
R346 B.n747 B.n392 585
R347 B.n392 B.n391 585
R348 B.n749 B.n748 585
R349 B.n750 B.n749 585
R350 B.n386 B.n385 585
R351 B.n387 B.n386 585
R352 B.n758 B.n757 585
R353 B.n757 B.n756 585
R354 B.n759 B.n384 585
R355 B.n384 B.n383 585
R356 B.n761 B.n760 585
R357 B.n762 B.n761 585
R358 B.n378 B.n377 585
R359 B.n379 B.n378 585
R360 B.n772 B.n771 585
R361 B.n771 B.n770 585
R362 B.n773 B.n376 585
R363 B.n769 B.n376 585
R364 B.n775 B.n774 585
R365 B.n776 B.n775 585
R366 B.n3 B.n0 585
R367 B.n4 B.n3 585
R368 B.n821 B.n1 585
R369 B.n822 B.n821 585
R370 B.n820 B.n819 585
R371 B.n820 B.n8 585
R372 B.n818 B.n9 585
R373 B.n12 B.n9 585
R374 B.n817 B.n816 585
R375 B.n816 B.n815 585
R376 B.n11 B.n10 585
R377 B.n814 B.n11 585
R378 B.n812 B.n811 585
R379 B.n813 B.n812 585
R380 B.n810 B.n17 585
R381 B.n17 B.n16 585
R382 B.n809 B.n808 585
R383 B.n808 B.n807 585
R384 B.n19 B.n18 585
R385 B.n806 B.n19 585
R386 B.n804 B.n803 585
R387 B.n805 B.n804 585
R388 B.n802 B.n24 585
R389 B.n24 B.n23 585
R390 B.n825 B.n824 585
R391 B.n823 B.n2 585
R392 B.n800 B.n24 578.989
R393 B.n797 B.n96 578.989
R394 B.n469 B.n390 578.989
R395 B.n745 B.n392 578.989
R396 B.n798 B.n94 256.663
R397 B.n798 B.n93 256.663
R398 B.n798 B.n92 256.663
R399 B.n798 B.n91 256.663
R400 B.n798 B.n90 256.663
R401 B.n798 B.n89 256.663
R402 B.n798 B.n88 256.663
R403 B.n798 B.n87 256.663
R404 B.n798 B.n86 256.663
R405 B.n798 B.n85 256.663
R406 B.n798 B.n84 256.663
R407 B.n798 B.n83 256.663
R408 B.n798 B.n82 256.663
R409 B.n798 B.n81 256.663
R410 B.n798 B.n80 256.663
R411 B.n798 B.n79 256.663
R412 B.n798 B.n78 256.663
R413 B.n798 B.n77 256.663
R414 B.n798 B.n76 256.663
R415 B.n798 B.n75 256.663
R416 B.n798 B.n74 256.663
R417 B.n798 B.n73 256.663
R418 B.n798 B.n72 256.663
R419 B.n798 B.n71 256.663
R420 B.n798 B.n70 256.663
R421 B.n798 B.n69 256.663
R422 B.n798 B.n68 256.663
R423 B.n798 B.n67 256.663
R424 B.n798 B.n66 256.663
R425 B.n798 B.n65 256.663
R426 B.n798 B.n64 256.663
R427 B.n798 B.n63 256.663
R428 B.n798 B.n62 256.663
R429 B.n798 B.n61 256.663
R430 B.n798 B.n60 256.663
R431 B.n798 B.n59 256.663
R432 B.n798 B.n58 256.663
R433 B.n798 B.n57 256.663
R434 B.n798 B.n56 256.663
R435 B.n798 B.n55 256.663
R436 B.n798 B.n54 256.663
R437 B.n798 B.n53 256.663
R438 B.n798 B.n52 256.663
R439 B.n798 B.n51 256.663
R440 B.n798 B.n50 256.663
R441 B.n798 B.n49 256.663
R442 B.n798 B.n48 256.663
R443 B.n798 B.n47 256.663
R444 B.n798 B.n46 256.663
R445 B.n798 B.n45 256.663
R446 B.n798 B.n44 256.663
R447 B.n798 B.n43 256.663
R448 B.n798 B.n42 256.663
R449 B.n798 B.n41 256.663
R450 B.n798 B.n40 256.663
R451 B.n798 B.n39 256.663
R452 B.n798 B.n38 256.663
R453 B.n798 B.n37 256.663
R454 B.n798 B.n36 256.663
R455 B.n798 B.n35 256.663
R456 B.n798 B.n34 256.663
R457 B.n798 B.n33 256.663
R458 B.n798 B.n32 256.663
R459 B.n798 B.n31 256.663
R460 B.n798 B.n30 256.663
R461 B.n798 B.n29 256.663
R462 B.n798 B.n28 256.663
R463 B.n798 B.n27 256.663
R464 B.n799 B.n798 256.663
R465 B.n744 B.n743 256.663
R466 B.n743 B.n395 256.663
R467 B.n743 B.n396 256.663
R468 B.n743 B.n397 256.663
R469 B.n743 B.n398 256.663
R470 B.n743 B.n399 256.663
R471 B.n743 B.n400 256.663
R472 B.n743 B.n401 256.663
R473 B.n743 B.n402 256.663
R474 B.n743 B.n403 256.663
R475 B.n743 B.n404 256.663
R476 B.n743 B.n405 256.663
R477 B.n743 B.n406 256.663
R478 B.n743 B.n407 256.663
R479 B.n743 B.n408 256.663
R480 B.n743 B.n409 256.663
R481 B.n743 B.n410 256.663
R482 B.n743 B.n411 256.663
R483 B.n743 B.n412 256.663
R484 B.n743 B.n413 256.663
R485 B.n743 B.n414 256.663
R486 B.n743 B.n415 256.663
R487 B.n743 B.n416 256.663
R488 B.n743 B.n417 256.663
R489 B.n743 B.n418 256.663
R490 B.n743 B.n419 256.663
R491 B.n743 B.n420 256.663
R492 B.n743 B.n421 256.663
R493 B.n743 B.n422 256.663
R494 B.n743 B.n423 256.663
R495 B.n743 B.n424 256.663
R496 B.n743 B.n425 256.663
R497 B.n743 B.n426 256.663
R498 B.n743 B.n427 256.663
R499 B.n743 B.n428 256.663
R500 B.n743 B.n429 256.663
R501 B.n743 B.n430 256.663
R502 B.n743 B.n431 256.663
R503 B.n743 B.n432 256.663
R504 B.n743 B.n433 256.663
R505 B.n743 B.n434 256.663
R506 B.n743 B.n435 256.663
R507 B.n743 B.n436 256.663
R508 B.n743 B.n437 256.663
R509 B.n743 B.n438 256.663
R510 B.n743 B.n439 256.663
R511 B.n743 B.n440 256.663
R512 B.n743 B.n441 256.663
R513 B.n743 B.n442 256.663
R514 B.n743 B.n443 256.663
R515 B.n743 B.n444 256.663
R516 B.n743 B.n445 256.663
R517 B.n743 B.n446 256.663
R518 B.n743 B.n447 256.663
R519 B.n743 B.n448 256.663
R520 B.n743 B.n449 256.663
R521 B.n743 B.n450 256.663
R522 B.n743 B.n451 256.663
R523 B.n743 B.n452 256.663
R524 B.n743 B.n453 256.663
R525 B.n743 B.n454 256.663
R526 B.n743 B.n455 256.663
R527 B.n743 B.n456 256.663
R528 B.n743 B.n457 256.663
R529 B.n743 B.n458 256.663
R530 B.n743 B.n459 256.663
R531 B.n743 B.n460 256.663
R532 B.n743 B.n461 256.663
R533 B.n743 B.n462 256.663
R534 B.n827 B.n826 256.663
R535 B.n102 B.n26 163.367
R536 B.n106 B.n105 163.367
R537 B.n110 B.n109 163.367
R538 B.n114 B.n113 163.367
R539 B.n118 B.n117 163.367
R540 B.n122 B.n121 163.367
R541 B.n126 B.n125 163.367
R542 B.n130 B.n129 163.367
R543 B.n134 B.n133 163.367
R544 B.n138 B.n137 163.367
R545 B.n142 B.n141 163.367
R546 B.n146 B.n145 163.367
R547 B.n150 B.n149 163.367
R548 B.n154 B.n153 163.367
R549 B.n158 B.n157 163.367
R550 B.n162 B.n161 163.367
R551 B.n166 B.n165 163.367
R552 B.n170 B.n169 163.367
R553 B.n174 B.n173 163.367
R554 B.n178 B.n177 163.367
R555 B.n182 B.n181 163.367
R556 B.n186 B.n185 163.367
R557 B.n190 B.n189 163.367
R558 B.n194 B.n193 163.367
R559 B.n198 B.n197 163.367
R560 B.n202 B.n201 163.367
R561 B.n206 B.n205 163.367
R562 B.n210 B.n209 163.367
R563 B.n214 B.n213 163.367
R564 B.n218 B.n217 163.367
R565 B.n222 B.n221 163.367
R566 B.n226 B.n225 163.367
R567 B.n231 B.n230 163.367
R568 B.n235 B.n234 163.367
R569 B.n239 B.n238 163.367
R570 B.n243 B.n242 163.367
R571 B.n247 B.n246 163.367
R572 B.n251 B.n250 163.367
R573 B.n255 B.n254 163.367
R574 B.n259 B.n258 163.367
R575 B.n263 B.n262 163.367
R576 B.n267 B.n266 163.367
R577 B.n271 B.n270 163.367
R578 B.n275 B.n274 163.367
R579 B.n279 B.n278 163.367
R580 B.n283 B.n282 163.367
R581 B.n287 B.n286 163.367
R582 B.n291 B.n290 163.367
R583 B.n295 B.n294 163.367
R584 B.n299 B.n298 163.367
R585 B.n303 B.n302 163.367
R586 B.n307 B.n306 163.367
R587 B.n311 B.n310 163.367
R588 B.n315 B.n314 163.367
R589 B.n319 B.n318 163.367
R590 B.n323 B.n322 163.367
R591 B.n327 B.n326 163.367
R592 B.n331 B.n330 163.367
R593 B.n335 B.n334 163.367
R594 B.n339 B.n338 163.367
R595 B.n343 B.n342 163.367
R596 B.n347 B.n346 163.367
R597 B.n351 B.n350 163.367
R598 B.n355 B.n354 163.367
R599 B.n359 B.n358 163.367
R600 B.n363 B.n362 163.367
R601 B.n367 B.n366 163.367
R602 B.n371 B.n370 163.367
R603 B.n797 B.n95 163.367
R604 B.n751 B.n390 163.367
R605 B.n751 B.n388 163.367
R606 B.n755 B.n388 163.367
R607 B.n755 B.n382 163.367
R608 B.n763 B.n382 163.367
R609 B.n763 B.n380 163.367
R610 B.n768 B.n380 163.367
R611 B.n768 B.n375 163.367
R612 B.n777 B.n375 163.367
R613 B.n778 B.n777 163.367
R614 B.n778 B.n5 163.367
R615 B.n6 B.n5 163.367
R616 B.n7 B.n6 163.367
R617 B.n784 B.n7 163.367
R618 B.n785 B.n784 163.367
R619 B.n785 B.n13 163.367
R620 B.n14 B.n13 163.367
R621 B.n15 B.n14 163.367
R622 B.n790 B.n15 163.367
R623 B.n790 B.n20 163.367
R624 B.n21 B.n20 163.367
R625 B.n22 B.n21 163.367
R626 B.n96 B.n22 163.367
R627 B.n742 B.n394 163.367
R628 B.n742 B.n463 163.367
R629 B.n738 B.n737 163.367
R630 B.n734 B.n733 163.367
R631 B.n730 B.n729 163.367
R632 B.n726 B.n725 163.367
R633 B.n722 B.n721 163.367
R634 B.n718 B.n717 163.367
R635 B.n714 B.n713 163.367
R636 B.n710 B.n709 163.367
R637 B.n706 B.n705 163.367
R638 B.n702 B.n701 163.367
R639 B.n698 B.n697 163.367
R640 B.n694 B.n693 163.367
R641 B.n690 B.n689 163.367
R642 B.n686 B.n685 163.367
R643 B.n682 B.n681 163.367
R644 B.n678 B.n677 163.367
R645 B.n674 B.n673 163.367
R646 B.n670 B.n669 163.367
R647 B.n666 B.n665 163.367
R648 B.n662 B.n661 163.367
R649 B.n658 B.n657 163.367
R650 B.n654 B.n653 163.367
R651 B.n650 B.n649 163.367
R652 B.n646 B.n645 163.367
R653 B.n642 B.n641 163.367
R654 B.n638 B.n637 163.367
R655 B.n634 B.n633 163.367
R656 B.n630 B.n629 163.367
R657 B.n626 B.n625 163.367
R658 B.n622 B.n621 163.367
R659 B.n618 B.n617 163.367
R660 B.n614 B.n613 163.367
R661 B.n610 B.n609 163.367
R662 B.n606 B.n605 163.367
R663 B.n602 B.n601 163.367
R664 B.n597 B.n596 163.367
R665 B.n593 B.n592 163.367
R666 B.n589 B.n588 163.367
R667 B.n585 B.n584 163.367
R668 B.n581 B.n580 163.367
R669 B.n577 B.n576 163.367
R670 B.n573 B.n572 163.367
R671 B.n569 B.n568 163.367
R672 B.n565 B.n564 163.367
R673 B.n561 B.n560 163.367
R674 B.n557 B.n556 163.367
R675 B.n553 B.n552 163.367
R676 B.n549 B.n548 163.367
R677 B.n545 B.n544 163.367
R678 B.n541 B.n540 163.367
R679 B.n537 B.n536 163.367
R680 B.n533 B.n532 163.367
R681 B.n529 B.n528 163.367
R682 B.n525 B.n524 163.367
R683 B.n521 B.n520 163.367
R684 B.n517 B.n516 163.367
R685 B.n513 B.n512 163.367
R686 B.n509 B.n508 163.367
R687 B.n505 B.n504 163.367
R688 B.n501 B.n500 163.367
R689 B.n497 B.n496 163.367
R690 B.n493 B.n492 163.367
R691 B.n489 B.n488 163.367
R692 B.n485 B.n484 163.367
R693 B.n481 B.n480 163.367
R694 B.n477 B.n476 163.367
R695 B.n473 B.n472 163.367
R696 B.n749 B.n392 163.367
R697 B.n749 B.n386 163.367
R698 B.n757 B.n386 163.367
R699 B.n757 B.n384 163.367
R700 B.n761 B.n384 163.367
R701 B.n761 B.n378 163.367
R702 B.n771 B.n378 163.367
R703 B.n771 B.n376 163.367
R704 B.n775 B.n376 163.367
R705 B.n775 B.n3 163.367
R706 B.n825 B.n3 163.367
R707 B.n821 B.n2 163.367
R708 B.n821 B.n820 163.367
R709 B.n820 B.n9 163.367
R710 B.n816 B.n9 163.367
R711 B.n816 B.n11 163.367
R712 B.n812 B.n11 163.367
R713 B.n812 B.n17 163.367
R714 B.n808 B.n17 163.367
R715 B.n808 B.n19 163.367
R716 B.n804 B.n19 163.367
R717 B.n804 B.n24 163.367
R718 B.n97 B.t4 82.855
R719 B.n467 B.t15 82.855
R720 B.n100 B.t7 82.8282
R721 B.n464 B.t12 82.8282
R722 B.n800 B.n799 71.676
R723 B.n102 B.n27 71.676
R724 B.n106 B.n28 71.676
R725 B.n110 B.n29 71.676
R726 B.n114 B.n30 71.676
R727 B.n118 B.n31 71.676
R728 B.n122 B.n32 71.676
R729 B.n126 B.n33 71.676
R730 B.n130 B.n34 71.676
R731 B.n134 B.n35 71.676
R732 B.n138 B.n36 71.676
R733 B.n142 B.n37 71.676
R734 B.n146 B.n38 71.676
R735 B.n150 B.n39 71.676
R736 B.n154 B.n40 71.676
R737 B.n158 B.n41 71.676
R738 B.n162 B.n42 71.676
R739 B.n166 B.n43 71.676
R740 B.n170 B.n44 71.676
R741 B.n174 B.n45 71.676
R742 B.n178 B.n46 71.676
R743 B.n182 B.n47 71.676
R744 B.n186 B.n48 71.676
R745 B.n190 B.n49 71.676
R746 B.n194 B.n50 71.676
R747 B.n198 B.n51 71.676
R748 B.n202 B.n52 71.676
R749 B.n206 B.n53 71.676
R750 B.n210 B.n54 71.676
R751 B.n214 B.n55 71.676
R752 B.n218 B.n56 71.676
R753 B.n222 B.n57 71.676
R754 B.n226 B.n58 71.676
R755 B.n231 B.n59 71.676
R756 B.n235 B.n60 71.676
R757 B.n239 B.n61 71.676
R758 B.n243 B.n62 71.676
R759 B.n247 B.n63 71.676
R760 B.n251 B.n64 71.676
R761 B.n255 B.n65 71.676
R762 B.n259 B.n66 71.676
R763 B.n263 B.n67 71.676
R764 B.n267 B.n68 71.676
R765 B.n271 B.n69 71.676
R766 B.n275 B.n70 71.676
R767 B.n279 B.n71 71.676
R768 B.n283 B.n72 71.676
R769 B.n287 B.n73 71.676
R770 B.n291 B.n74 71.676
R771 B.n295 B.n75 71.676
R772 B.n299 B.n76 71.676
R773 B.n303 B.n77 71.676
R774 B.n307 B.n78 71.676
R775 B.n311 B.n79 71.676
R776 B.n315 B.n80 71.676
R777 B.n319 B.n81 71.676
R778 B.n323 B.n82 71.676
R779 B.n327 B.n83 71.676
R780 B.n331 B.n84 71.676
R781 B.n335 B.n85 71.676
R782 B.n339 B.n86 71.676
R783 B.n343 B.n87 71.676
R784 B.n347 B.n88 71.676
R785 B.n351 B.n89 71.676
R786 B.n355 B.n90 71.676
R787 B.n359 B.n91 71.676
R788 B.n363 B.n92 71.676
R789 B.n367 B.n93 71.676
R790 B.n371 B.n94 71.676
R791 B.n95 B.n94 71.676
R792 B.n370 B.n93 71.676
R793 B.n366 B.n92 71.676
R794 B.n362 B.n91 71.676
R795 B.n358 B.n90 71.676
R796 B.n354 B.n89 71.676
R797 B.n350 B.n88 71.676
R798 B.n346 B.n87 71.676
R799 B.n342 B.n86 71.676
R800 B.n338 B.n85 71.676
R801 B.n334 B.n84 71.676
R802 B.n330 B.n83 71.676
R803 B.n326 B.n82 71.676
R804 B.n322 B.n81 71.676
R805 B.n318 B.n80 71.676
R806 B.n314 B.n79 71.676
R807 B.n310 B.n78 71.676
R808 B.n306 B.n77 71.676
R809 B.n302 B.n76 71.676
R810 B.n298 B.n75 71.676
R811 B.n294 B.n74 71.676
R812 B.n290 B.n73 71.676
R813 B.n286 B.n72 71.676
R814 B.n282 B.n71 71.676
R815 B.n278 B.n70 71.676
R816 B.n274 B.n69 71.676
R817 B.n270 B.n68 71.676
R818 B.n266 B.n67 71.676
R819 B.n262 B.n66 71.676
R820 B.n258 B.n65 71.676
R821 B.n254 B.n64 71.676
R822 B.n250 B.n63 71.676
R823 B.n246 B.n62 71.676
R824 B.n242 B.n61 71.676
R825 B.n238 B.n60 71.676
R826 B.n234 B.n59 71.676
R827 B.n230 B.n58 71.676
R828 B.n225 B.n57 71.676
R829 B.n221 B.n56 71.676
R830 B.n217 B.n55 71.676
R831 B.n213 B.n54 71.676
R832 B.n209 B.n53 71.676
R833 B.n205 B.n52 71.676
R834 B.n201 B.n51 71.676
R835 B.n197 B.n50 71.676
R836 B.n193 B.n49 71.676
R837 B.n189 B.n48 71.676
R838 B.n185 B.n47 71.676
R839 B.n181 B.n46 71.676
R840 B.n177 B.n45 71.676
R841 B.n173 B.n44 71.676
R842 B.n169 B.n43 71.676
R843 B.n165 B.n42 71.676
R844 B.n161 B.n41 71.676
R845 B.n157 B.n40 71.676
R846 B.n153 B.n39 71.676
R847 B.n149 B.n38 71.676
R848 B.n145 B.n37 71.676
R849 B.n141 B.n36 71.676
R850 B.n137 B.n35 71.676
R851 B.n133 B.n34 71.676
R852 B.n129 B.n33 71.676
R853 B.n125 B.n32 71.676
R854 B.n121 B.n31 71.676
R855 B.n117 B.n30 71.676
R856 B.n113 B.n29 71.676
R857 B.n109 B.n28 71.676
R858 B.n105 B.n27 71.676
R859 B.n799 B.n26 71.676
R860 B.n745 B.n744 71.676
R861 B.n463 B.n395 71.676
R862 B.n737 B.n396 71.676
R863 B.n733 B.n397 71.676
R864 B.n729 B.n398 71.676
R865 B.n725 B.n399 71.676
R866 B.n721 B.n400 71.676
R867 B.n717 B.n401 71.676
R868 B.n713 B.n402 71.676
R869 B.n709 B.n403 71.676
R870 B.n705 B.n404 71.676
R871 B.n701 B.n405 71.676
R872 B.n697 B.n406 71.676
R873 B.n693 B.n407 71.676
R874 B.n689 B.n408 71.676
R875 B.n685 B.n409 71.676
R876 B.n681 B.n410 71.676
R877 B.n677 B.n411 71.676
R878 B.n673 B.n412 71.676
R879 B.n669 B.n413 71.676
R880 B.n665 B.n414 71.676
R881 B.n661 B.n415 71.676
R882 B.n657 B.n416 71.676
R883 B.n653 B.n417 71.676
R884 B.n649 B.n418 71.676
R885 B.n645 B.n419 71.676
R886 B.n641 B.n420 71.676
R887 B.n637 B.n421 71.676
R888 B.n633 B.n422 71.676
R889 B.n629 B.n423 71.676
R890 B.n625 B.n424 71.676
R891 B.n621 B.n425 71.676
R892 B.n617 B.n426 71.676
R893 B.n613 B.n427 71.676
R894 B.n609 B.n428 71.676
R895 B.n605 B.n429 71.676
R896 B.n601 B.n430 71.676
R897 B.n596 B.n431 71.676
R898 B.n592 B.n432 71.676
R899 B.n588 B.n433 71.676
R900 B.n584 B.n434 71.676
R901 B.n580 B.n435 71.676
R902 B.n576 B.n436 71.676
R903 B.n572 B.n437 71.676
R904 B.n568 B.n438 71.676
R905 B.n564 B.n439 71.676
R906 B.n560 B.n440 71.676
R907 B.n556 B.n441 71.676
R908 B.n552 B.n442 71.676
R909 B.n548 B.n443 71.676
R910 B.n544 B.n444 71.676
R911 B.n540 B.n445 71.676
R912 B.n536 B.n446 71.676
R913 B.n532 B.n447 71.676
R914 B.n528 B.n448 71.676
R915 B.n524 B.n449 71.676
R916 B.n520 B.n450 71.676
R917 B.n516 B.n451 71.676
R918 B.n512 B.n452 71.676
R919 B.n508 B.n453 71.676
R920 B.n504 B.n454 71.676
R921 B.n500 B.n455 71.676
R922 B.n496 B.n456 71.676
R923 B.n492 B.n457 71.676
R924 B.n488 B.n458 71.676
R925 B.n484 B.n459 71.676
R926 B.n480 B.n460 71.676
R927 B.n476 B.n461 71.676
R928 B.n472 B.n462 71.676
R929 B.n744 B.n394 71.676
R930 B.n738 B.n395 71.676
R931 B.n734 B.n396 71.676
R932 B.n730 B.n397 71.676
R933 B.n726 B.n398 71.676
R934 B.n722 B.n399 71.676
R935 B.n718 B.n400 71.676
R936 B.n714 B.n401 71.676
R937 B.n710 B.n402 71.676
R938 B.n706 B.n403 71.676
R939 B.n702 B.n404 71.676
R940 B.n698 B.n405 71.676
R941 B.n694 B.n406 71.676
R942 B.n690 B.n407 71.676
R943 B.n686 B.n408 71.676
R944 B.n682 B.n409 71.676
R945 B.n678 B.n410 71.676
R946 B.n674 B.n411 71.676
R947 B.n670 B.n412 71.676
R948 B.n666 B.n413 71.676
R949 B.n662 B.n414 71.676
R950 B.n658 B.n415 71.676
R951 B.n654 B.n416 71.676
R952 B.n650 B.n417 71.676
R953 B.n646 B.n418 71.676
R954 B.n642 B.n419 71.676
R955 B.n638 B.n420 71.676
R956 B.n634 B.n421 71.676
R957 B.n630 B.n422 71.676
R958 B.n626 B.n423 71.676
R959 B.n622 B.n424 71.676
R960 B.n618 B.n425 71.676
R961 B.n614 B.n426 71.676
R962 B.n610 B.n427 71.676
R963 B.n606 B.n428 71.676
R964 B.n602 B.n429 71.676
R965 B.n597 B.n430 71.676
R966 B.n593 B.n431 71.676
R967 B.n589 B.n432 71.676
R968 B.n585 B.n433 71.676
R969 B.n581 B.n434 71.676
R970 B.n577 B.n435 71.676
R971 B.n573 B.n436 71.676
R972 B.n569 B.n437 71.676
R973 B.n565 B.n438 71.676
R974 B.n561 B.n439 71.676
R975 B.n557 B.n440 71.676
R976 B.n553 B.n441 71.676
R977 B.n549 B.n442 71.676
R978 B.n545 B.n443 71.676
R979 B.n541 B.n444 71.676
R980 B.n537 B.n445 71.676
R981 B.n533 B.n446 71.676
R982 B.n529 B.n447 71.676
R983 B.n525 B.n448 71.676
R984 B.n521 B.n449 71.676
R985 B.n517 B.n450 71.676
R986 B.n513 B.n451 71.676
R987 B.n509 B.n452 71.676
R988 B.n505 B.n453 71.676
R989 B.n501 B.n454 71.676
R990 B.n497 B.n455 71.676
R991 B.n493 B.n456 71.676
R992 B.n489 B.n457 71.676
R993 B.n485 B.n458 71.676
R994 B.n481 B.n459 71.676
R995 B.n477 B.n460 71.676
R996 B.n473 B.n461 71.676
R997 B.n469 B.n462 71.676
R998 B.n826 B.n825 71.676
R999 B.n826 B.n2 71.676
R1000 B.n98 B.t5 70.8307
R1001 B.n468 B.t14 70.8307
R1002 B.n101 B.t8 70.804
R1003 B.n465 B.t11 70.804
R1004 B.n743 B.n391 61.5359
R1005 B.n798 B.n23 61.5359
R1006 B.n228 B.n101 59.5399
R1007 B.n99 B.n98 59.5399
R1008 B.n599 B.n468 59.5399
R1009 B.n466 B.n465 59.5399
R1010 B.n747 B.n746 37.62
R1011 B.n470 B.n389 37.62
R1012 B.n796 B.n795 37.62
R1013 B.n802 B.n801 37.62
R1014 B.n750 B.n391 29.6772
R1015 B.n750 B.n387 29.6772
R1016 B.n756 B.n387 29.6772
R1017 B.n762 B.n383 29.6772
R1018 B.n762 B.n379 29.6772
R1019 B.n770 B.n379 29.6772
R1020 B.n770 B.n769 29.6772
R1021 B.n776 B.n4 29.6772
R1022 B.n824 B.n4 29.6772
R1023 B.n824 B.n823 29.6772
R1024 B.n823 B.n822 29.6772
R1025 B.n822 B.n8 29.6772
R1026 B.n815 B.n12 29.6772
R1027 B.n815 B.n814 29.6772
R1028 B.n814 B.n813 29.6772
R1029 B.n813 B.n16 29.6772
R1030 B.n807 B.n806 29.6772
R1031 B.n806 B.n805 29.6772
R1032 B.n805 B.n23 29.6772
R1033 B.n769 B.t0 29.2407
R1034 B.n12 B.t1 29.2407
R1035 B.n756 B.t10 28.3679
R1036 B.n807 B.t3 28.3679
R1037 B B.n827 18.0485
R1038 B.n101 B.n100 12.0247
R1039 B.n98 B.n97 12.0247
R1040 B.n468 B.n467 12.0247
R1041 B.n465 B.n464 12.0247
R1042 B.n748 B.n747 10.6151
R1043 B.n748 B.n385 10.6151
R1044 B.n758 B.n385 10.6151
R1045 B.n759 B.n758 10.6151
R1046 B.n760 B.n759 10.6151
R1047 B.n760 B.n377 10.6151
R1048 B.n772 B.n377 10.6151
R1049 B.n773 B.n772 10.6151
R1050 B.n774 B.n773 10.6151
R1051 B.n774 B.n0 10.6151
R1052 B.n746 B.n393 10.6151
R1053 B.n741 B.n393 10.6151
R1054 B.n741 B.n740 10.6151
R1055 B.n740 B.n739 10.6151
R1056 B.n739 B.n736 10.6151
R1057 B.n736 B.n735 10.6151
R1058 B.n735 B.n732 10.6151
R1059 B.n732 B.n731 10.6151
R1060 B.n731 B.n728 10.6151
R1061 B.n728 B.n727 10.6151
R1062 B.n727 B.n724 10.6151
R1063 B.n724 B.n723 10.6151
R1064 B.n723 B.n720 10.6151
R1065 B.n720 B.n719 10.6151
R1066 B.n719 B.n716 10.6151
R1067 B.n716 B.n715 10.6151
R1068 B.n715 B.n712 10.6151
R1069 B.n712 B.n711 10.6151
R1070 B.n711 B.n708 10.6151
R1071 B.n708 B.n707 10.6151
R1072 B.n707 B.n704 10.6151
R1073 B.n704 B.n703 10.6151
R1074 B.n703 B.n700 10.6151
R1075 B.n700 B.n699 10.6151
R1076 B.n699 B.n696 10.6151
R1077 B.n696 B.n695 10.6151
R1078 B.n695 B.n692 10.6151
R1079 B.n692 B.n691 10.6151
R1080 B.n691 B.n688 10.6151
R1081 B.n688 B.n687 10.6151
R1082 B.n687 B.n684 10.6151
R1083 B.n684 B.n683 10.6151
R1084 B.n683 B.n680 10.6151
R1085 B.n680 B.n679 10.6151
R1086 B.n679 B.n676 10.6151
R1087 B.n676 B.n675 10.6151
R1088 B.n675 B.n672 10.6151
R1089 B.n672 B.n671 10.6151
R1090 B.n671 B.n668 10.6151
R1091 B.n668 B.n667 10.6151
R1092 B.n667 B.n664 10.6151
R1093 B.n664 B.n663 10.6151
R1094 B.n663 B.n660 10.6151
R1095 B.n660 B.n659 10.6151
R1096 B.n659 B.n656 10.6151
R1097 B.n656 B.n655 10.6151
R1098 B.n655 B.n652 10.6151
R1099 B.n652 B.n651 10.6151
R1100 B.n651 B.n648 10.6151
R1101 B.n648 B.n647 10.6151
R1102 B.n647 B.n644 10.6151
R1103 B.n644 B.n643 10.6151
R1104 B.n643 B.n640 10.6151
R1105 B.n640 B.n639 10.6151
R1106 B.n639 B.n636 10.6151
R1107 B.n636 B.n635 10.6151
R1108 B.n635 B.n632 10.6151
R1109 B.n632 B.n631 10.6151
R1110 B.n631 B.n628 10.6151
R1111 B.n628 B.n627 10.6151
R1112 B.n627 B.n624 10.6151
R1113 B.n624 B.n623 10.6151
R1114 B.n623 B.n620 10.6151
R1115 B.n620 B.n619 10.6151
R1116 B.n616 B.n615 10.6151
R1117 B.n615 B.n612 10.6151
R1118 B.n612 B.n611 10.6151
R1119 B.n611 B.n608 10.6151
R1120 B.n608 B.n607 10.6151
R1121 B.n607 B.n604 10.6151
R1122 B.n604 B.n603 10.6151
R1123 B.n603 B.n600 10.6151
R1124 B.n598 B.n595 10.6151
R1125 B.n595 B.n594 10.6151
R1126 B.n594 B.n591 10.6151
R1127 B.n591 B.n590 10.6151
R1128 B.n590 B.n587 10.6151
R1129 B.n587 B.n586 10.6151
R1130 B.n586 B.n583 10.6151
R1131 B.n583 B.n582 10.6151
R1132 B.n582 B.n579 10.6151
R1133 B.n579 B.n578 10.6151
R1134 B.n578 B.n575 10.6151
R1135 B.n575 B.n574 10.6151
R1136 B.n574 B.n571 10.6151
R1137 B.n571 B.n570 10.6151
R1138 B.n570 B.n567 10.6151
R1139 B.n567 B.n566 10.6151
R1140 B.n566 B.n563 10.6151
R1141 B.n563 B.n562 10.6151
R1142 B.n562 B.n559 10.6151
R1143 B.n559 B.n558 10.6151
R1144 B.n558 B.n555 10.6151
R1145 B.n555 B.n554 10.6151
R1146 B.n554 B.n551 10.6151
R1147 B.n551 B.n550 10.6151
R1148 B.n550 B.n547 10.6151
R1149 B.n547 B.n546 10.6151
R1150 B.n546 B.n543 10.6151
R1151 B.n543 B.n542 10.6151
R1152 B.n542 B.n539 10.6151
R1153 B.n539 B.n538 10.6151
R1154 B.n538 B.n535 10.6151
R1155 B.n535 B.n534 10.6151
R1156 B.n534 B.n531 10.6151
R1157 B.n531 B.n530 10.6151
R1158 B.n530 B.n527 10.6151
R1159 B.n527 B.n526 10.6151
R1160 B.n526 B.n523 10.6151
R1161 B.n523 B.n522 10.6151
R1162 B.n522 B.n519 10.6151
R1163 B.n519 B.n518 10.6151
R1164 B.n518 B.n515 10.6151
R1165 B.n515 B.n514 10.6151
R1166 B.n514 B.n511 10.6151
R1167 B.n511 B.n510 10.6151
R1168 B.n510 B.n507 10.6151
R1169 B.n507 B.n506 10.6151
R1170 B.n506 B.n503 10.6151
R1171 B.n503 B.n502 10.6151
R1172 B.n502 B.n499 10.6151
R1173 B.n499 B.n498 10.6151
R1174 B.n498 B.n495 10.6151
R1175 B.n495 B.n494 10.6151
R1176 B.n494 B.n491 10.6151
R1177 B.n491 B.n490 10.6151
R1178 B.n490 B.n487 10.6151
R1179 B.n487 B.n486 10.6151
R1180 B.n486 B.n483 10.6151
R1181 B.n483 B.n482 10.6151
R1182 B.n482 B.n479 10.6151
R1183 B.n479 B.n478 10.6151
R1184 B.n478 B.n475 10.6151
R1185 B.n475 B.n474 10.6151
R1186 B.n474 B.n471 10.6151
R1187 B.n471 B.n470 10.6151
R1188 B.n752 B.n389 10.6151
R1189 B.n753 B.n752 10.6151
R1190 B.n754 B.n753 10.6151
R1191 B.n754 B.n381 10.6151
R1192 B.n764 B.n381 10.6151
R1193 B.n765 B.n764 10.6151
R1194 B.n767 B.n765 10.6151
R1195 B.n767 B.n766 10.6151
R1196 B.n766 B.n374 10.6151
R1197 B.n779 B.n374 10.6151
R1198 B.n780 B.n779 10.6151
R1199 B.n781 B.n780 10.6151
R1200 B.n782 B.n781 10.6151
R1201 B.n783 B.n782 10.6151
R1202 B.n786 B.n783 10.6151
R1203 B.n787 B.n786 10.6151
R1204 B.n788 B.n787 10.6151
R1205 B.n789 B.n788 10.6151
R1206 B.n791 B.n789 10.6151
R1207 B.n792 B.n791 10.6151
R1208 B.n793 B.n792 10.6151
R1209 B.n794 B.n793 10.6151
R1210 B.n795 B.n794 10.6151
R1211 B.n819 B.n1 10.6151
R1212 B.n819 B.n818 10.6151
R1213 B.n818 B.n817 10.6151
R1214 B.n817 B.n10 10.6151
R1215 B.n811 B.n10 10.6151
R1216 B.n811 B.n810 10.6151
R1217 B.n810 B.n809 10.6151
R1218 B.n809 B.n18 10.6151
R1219 B.n803 B.n18 10.6151
R1220 B.n803 B.n802 10.6151
R1221 B.n801 B.n25 10.6151
R1222 B.n103 B.n25 10.6151
R1223 B.n104 B.n103 10.6151
R1224 B.n107 B.n104 10.6151
R1225 B.n108 B.n107 10.6151
R1226 B.n111 B.n108 10.6151
R1227 B.n112 B.n111 10.6151
R1228 B.n115 B.n112 10.6151
R1229 B.n116 B.n115 10.6151
R1230 B.n119 B.n116 10.6151
R1231 B.n120 B.n119 10.6151
R1232 B.n123 B.n120 10.6151
R1233 B.n124 B.n123 10.6151
R1234 B.n127 B.n124 10.6151
R1235 B.n128 B.n127 10.6151
R1236 B.n131 B.n128 10.6151
R1237 B.n132 B.n131 10.6151
R1238 B.n135 B.n132 10.6151
R1239 B.n136 B.n135 10.6151
R1240 B.n139 B.n136 10.6151
R1241 B.n140 B.n139 10.6151
R1242 B.n143 B.n140 10.6151
R1243 B.n144 B.n143 10.6151
R1244 B.n147 B.n144 10.6151
R1245 B.n148 B.n147 10.6151
R1246 B.n151 B.n148 10.6151
R1247 B.n152 B.n151 10.6151
R1248 B.n155 B.n152 10.6151
R1249 B.n156 B.n155 10.6151
R1250 B.n159 B.n156 10.6151
R1251 B.n160 B.n159 10.6151
R1252 B.n163 B.n160 10.6151
R1253 B.n164 B.n163 10.6151
R1254 B.n167 B.n164 10.6151
R1255 B.n168 B.n167 10.6151
R1256 B.n171 B.n168 10.6151
R1257 B.n172 B.n171 10.6151
R1258 B.n175 B.n172 10.6151
R1259 B.n176 B.n175 10.6151
R1260 B.n179 B.n176 10.6151
R1261 B.n180 B.n179 10.6151
R1262 B.n183 B.n180 10.6151
R1263 B.n184 B.n183 10.6151
R1264 B.n187 B.n184 10.6151
R1265 B.n188 B.n187 10.6151
R1266 B.n191 B.n188 10.6151
R1267 B.n192 B.n191 10.6151
R1268 B.n195 B.n192 10.6151
R1269 B.n196 B.n195 10.6151
R1270 B.n199 B.n196 10.6151
R1271 B.n200 B.n199 10.6151
R1272 B.n203 B.n200 10.6151
R1273 B.n204 B.n203 10.6151
R1274 B.n207 B.n204 10.6151
R1275 B.n208 B.n207 10.6151
R1276 B.n211 B.n208 10.6151
R1277 B.n212 B.n211 10.6151
R1278 B.n215 B.n212 10.6151
R1279 B.n216 B.n215 10.6151
R1280 B.n219 B.n216 10.6151
R1281 B.n220 B.n219 10.6151
R1282 B.n223 B.n220 10.6151
R1283 B.n224 B.n223 10.6151
R1284 B.n227 B.n224 10.6151
R1285 B.n232 B.n229 10.6151
R1286 B.n233 B.n232 10.6151
R1287 B.n236 B.n233 10.6151
R1288 B.n237 B.n236 10.6151
R1289 B.n240 B.n237 10.6151
R1290 B.n241 B.n240 10.6151
R1291 B.n244 B.n241 10.6151
R1292 B.n245 B.n244 10.6151
R1293 B.n249 B.n248 10.6151
R1294 B.n252 B.n249 10.6151
R1295 B.n253 B.n252 10.6151
R1296 B.n256 B.n253 10.6151
R1297 B.n257 B.n256 10.6151
R1298 B.n260 B.n257 10.6151
R1299 B.n261 B.n260 10.6151
R1300 B.n264 B.n261 10.6151
R1301 B.n265 B.n264 10.6151
R1302 B.n268 B.n265 10.6151
R1303 B.n269 B.n268 10.6151
R1304 B.n272 B.n269 10.6151
R1305 B.n273 B.n272 10.6151
R1306 B.n276 B.n273 10.6151
R1307 B.n277 B.n276 10.6151
R1308 B.n280 B.n277 10.6151
R1309 B.n281 B.n280 10.6151
R1310 B.n284 B.n281 10.6151
R1311 B.n285 B.n284 10.6151
R1312 B.n288 B.n285 10.6151
R1313 B.n289 B.n288 10.6151
R1314 B.n292 B.n289 10.6151
R1315 B.n293 B.n292 10.6151
R1316 B.n296 B.n293 10.6151
R1317 B.n297 B.n296 10.6151
R1318 B.n300 B.n297 10.6151
R1319 B.n301 B.n300 10.6151
R1320 B.n304 B.n301 10.6151
R1321 B.n305 B.n304 10.6151
R1322 B.n308 B.n305 10.6151
R1323 B.n309 B.n308 10.6151
R1324 B.n312 B.n309 10.6151
R1325 B.n313 B.n312 10.6151
R1326 B.n316 B.n313 10.6151
R1327 B.n317 B.n316 10.6151
R1328 B.n320 B.n317 10.6151
R1329 B.n321 B.n320 10.6151
R1330 B.n324 B.n321 10.6151
R1331 B.n325 B.n324 10.6151
R1332 B.n328 B.n325 10.6151
R1333 B.n329 B.n328 10.6151
R1334 B.n332 B.n329 10.6151
R1335 B.n333 B.n332 10.6151
R1336 B.n336 B.n333 10.6151
R1337 B.n337 B.n336 10.6151
R1338 B.n340 B.n337 10.6151
R1339 B.n341 B.n340 10.6151
R1340 B.n344 B.n341 10.6151
R1341 B.n345 B.n344 10.6151
R1342 B.n348 B.n345 10.6151
R1343 B.n349 B.n348 10.6151
R1344 B.n352 B.n349 10.6151
R1345 B.n353 B.n352 10.6151
R1346 B.n356 B.n353 10.6151
R1347 B.n357 B.n356 10.6151
R1348 B.n360 B.n357 10.6151
R1349 B.n361 B.n360 10.6151
R1350 B.n364 B.n361 10.6151
R1351 B.n365 B.n364 10.6151
R1352 B.n368 B.n365 10.6151
R1353 B.n369 B.n368 10.6151
R1354 B.n372 B.n369 10.6151
R1355 B.n373 B.n372 10.6151
R1356 B.n796 B.n373 10.6151
R1357 B.n827 B.n0 8.11757
R1358 B.n827 B.n1 8.11757
R1359 B.n616 B.n466 7.18099
R1360 B.n600 B.n599 7.18099
R1361 B.n229 B.n228 7.18099
R1362 B.n245 B.n99 7.18099
R1363 B.n619 B.n466 3.43465
R1364 B.n599 B.n598 3.43465
R1365 B.n228 B.n227 3.43465
R1366 B.n248 B.n99 3.43465
R1367 B.t10 B.n383 1.30976
R1368 B.t3 B.n16 1.30976
R1369 B.n776 B.t0 0.436921
R1370 B.t1 B.n8 0.436921
R1371 VP.n0 VP.t0 1993.39
R1372 VP.n0 VP.t1 1948.86
R1373 VP VP.n0 0.0516364
R1374 VDD1 VDD1.t0 108.228
R1375 VDD1 VDD1.t1 65.8515
C0 VDD1 VTAIL 10.9263f
C1 VTAIL VN 1.25557f
C2 VDD2 VTAIL 10.949901f
C3 VDD1 VN 0.148396f
C4 VTAIL VP 1.27076f
C5 VDD2 VDD1 0.428737f
C6 VDD2 VN 2.221f
C7 VDD1 VP 2.30371f
C8 VN VP 5.84328f
C9 VDD2 VP 0.23944f
C10 VDD2 B 5.026474f
C11 VDD1 B 8.8757f
C12 VTAIL B 8.38237f
C13 VN B 10.14496f
C14 VP B 4.084732f
C15 VDD1.t1 B 4.33815f
C16 VDD1.t0 B 5.09509f
C17 VP.t0 B 1.0685f
C18 VP.t1 B 1.00091f
C19 VP.n0 B 6.02345f
C20 VDD2.t0 B 5.06167f
C21 VDD2.t1 B 4.33299f
C22 VDD2.n0 B 3.66997f
C23 VTAIL.t0 B 3.68586f
C24 VTAIL.n0 B 1.77672f
C25 VTAIL.t2 B 3.68586f
C26 VTAIL.n1 B 1.78167f
C27 VTAIL.t1 B 3.68586f
C28 VTAIL.n2 B 1.74661f
C29 VTAIL.t3 B 3.68586f
C30 VTAIL.n3 B 1.70321f
C31 VN.t1 B 0.978478f
C32 VN.t0 B 1.04594f
.ends

