* NGSPICE file created from diff_pair_sample_1548.ext - technology: sky130A

.subckt diff_pair_sample_1548 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=2.7621 ps=17.07 w=16.74 l=1.38
X1 VTAIL.t5 VP.t0 VDD1.t7 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=2.7621 ps=17.07 w=16.74 l=1.38
X2 VDD1.t6 VP.t1 VTAIL.t2 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X3 VTAIL.t3 VP.t2 VDD1.t5 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X4 VTAIL.t7 VP.t3 VDD1.t4 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=2.7621 ps=17.07 w=16.74 l=1.38
X5 B.t11 B.t9 B.t10 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=0 ps=0 w=16.74 l=1.38
X6 B.t8 B.t6 B.t7 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=0 ps=0 w=16.74 l=1.38
X7 VDD2.t2 VN.t1 VTAIL.t14 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=6.5286 ps=34.26 w=16.74 l=1.38
X8 VTAIL.t13 VN.t2 VDD2.t5 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=2.7621 ps=17.07 w=16.74 l=1.38
X9 VDD1.t3 VP.t4 VTAIL.t1 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=6.5286 ps=34.26 w=16.74 l=1.38
X10 B.t5 B.t3 B.t4 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=0 ps=0 w=16.74 l=1.38
X11 VDD2.t4 VN.t3 VTAIL.t12 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X12 VDD2.t7 VN.t4 VTAIL.t11 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X13 VTAIL.t4 VP.t5 VDD1.t2 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X14 B.t2 B.t0 B.t1 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=6.5286 pd=34.26 as=0 ps=0 w=16.74 l=1.38
X15 VDD1.t1 VP.t6 VTAIL.t6 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=6.5286 ps=34.26 w=16.74 l=1.38
X16 VDD1.t0 VP.t7 VTAIL.t0 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X17 VTAIL.t10 VN.t5 VDD2.t6 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X18 VTAIL.t9 VN.t6 VDD2.t1 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=2.7621 ps=17.07 w=16.74 l=1.38
X19 VDD2.t0 VN.t7 VTAIL.t8 w_n2680_n4316# sky130_fd_pr__pfet_01v8 ad=2.7621 pd=17.07 as=6.5286 ps=34.26 w=16.74 l=1.38
R0 VN.n5 VN.t2 323.56
R1 VN.n25 VN.t1 323.56
R2 VN.n4 VN.t4 292.344
R3 VN.n10 VN.t5 292.344
R4 VN.n17 VN.t7 292.344
R5 VN.n24 VN.t6 292.344
R6 VN.n22 VN.t3 292.344
R7 VN.n36 VN.t0 292.344
R8 VN.n18 VN.n17 170.399
R9 VN.n37 VN.n36 170.399
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n29 VN.n21 161.3
R15 VN.n28 VN.n27 161.3
R16 VN.n26 VN.n23 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n5 VN.n4 59.9731
R25 VN.n25 VN.n24 59.9731
R26 VN.n9 VN.n8 56.5617
R27 VN.n29 VN.n28 56.5617
R28 VN VN.n37 49.1388
R29 VN.n15 VN.n1 44.4521
R30 VN.n34 VN.n20 44.4521
R31 VN.n16 VN.n15 36.702
R32 VN.n35 VN.n34 36.702
R33 VN.n26 VN.n25 26.618
R34 VN.n6 VN.n5 26.618
R35 VN.n8 VN.n3 24.5923
R36 VN.n11 VN.n9 24.5923
R37 VN.n28 VN.n23 24.5923
R38 VN.n30 VN.n29 24.5923
R39 VN.n10 VN.n1 19.4281
R40 VN.n22 VN.n20 19.4281
R41 VN.n17 VN.n16 15.4934
R42 VN.n36 VN.n35 15.4934
R43 VN.n4 VN.n3 5.16479
R44 VN.n11 VN.n10 5.16479
R45 VN.n24 VN.n23 5.16479
R46 VN.n30 VN.n22 5.16479
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n27 VN.n21 0.189894
R53 VN.n27 VN.n26 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VDD2.n2 VDD2.n1 68.9099
R63 VDD2.n2 VDD2.n0 68.9099
R64 VDD2 VDD2.n5 68.9071
R65 VDD2.n4 VDD2.n3 68.2284
R66 VDD2.n4 VDD2.n2 44.7799
R67 VDD2.n5 VDD2.t1 1.94226
R68 VDD2.n5 VDD2.t2 1.94226
R69 VDD2.n3 VDD2.t3 1.94226
R70 VDD2.n3 VDD2.t4 1.94226
R71 VDD2.n1 VDD2.t6 1.94226
R72 VDD2.n1 VDD2.t0 1.94226
R73 VDD2.n0 VDD2.t5 1.94226
R74 VDD2.n0 VDD2.t7 1.94226
R75 VDD2 VDD2.n4 0.795759
R76 VTAIL.n754 VTAIL.n666 756.745
R77 VTAIL.n90 VTAIL.n2 756.745
R78 VTAIL.n184 VTAIL.n96 756.745
R79 VTAIL.n280 VTAIL.n192 756.745
R80 VTAIL.n660 VTAIL.n572 756.745
R81 VTAIL.n564 VTAIL.n476 756.745
R82 VTAIL.n470 VTAIL.n382 756.745
R83 VTAIL.n374 VTAIL.n286 756.745
R84 VTAIL.n697 VTAIL.n696 585
R85 VTAIL.n694 VTAIL.n693 585
R86 VTAIL.n703 VTAIL.n702 585
R87 VTAIL.n705 VTAIL.n704 585
R88 VTAIL.n690 VTAIL.n689 585
R89 VTAIL.n711 VTAIL.n710 585
R90 VTAIL.n713 VTAIL.n712 585
R91 VTAIL.n686 VTAIL.n685 585
R92 VTAIL.n719 VTAIL.n718 585
R93 VTAIL.n721 VTAIL.n720 585
R94 VTAIL.n682 VTAIL.n681 585
R95 VTAIL.n727 VTAIL.n726 585
R96 VTAIL.n729 VTAIL.n728 585
R97 VTAIL.n678 VTAIL.n677 585
R98 VTAIL.n735 VTAIL.n734 585
R99 VTAIL.n738 VTAIL.n737 585
R100 VTAIL.n736 VTAIL.n674 585
R101 VTAIL.n743 VTAIL.n673 585
R102 VTAIL.n745 VTAIL.n744 585
R103 VTAIL.n747 VTAIL.n746 585
R104 VTAIL.n670 VTAIL.n669 585
R105 VTAIL.n753 VTAIL.n752 585
R106 VTAIL.n755 VTAIL.n754 585
R107 VTAIL.n33 VTAIL.n32 585
R108 VTAIL.n30 VTAIL.n29 585
R109 VTAIL.n39 VTAIL.n38 585
R110 VTAIL.n41 VTAIL.n40 585
R111 VTAIL.n26 VTAIL.n25 585
R112 VTAIL.n47 VTAIL.n46 585
R113 VTAIL.n49 VTAIL.n48 585
R114 VTAIL.n22 VTAIL.n21 585
R115 VTAIL.n55 VTAIL.n54 585
R116 VTAIL.n57 VTAIL.n56 585
R117 VTAIL.n18 VTAIL.n17 585
R118 VTAIL.n63 VTAIL.n62 585
R119 VTAIL.n65 VTAIL.n64 585
R120 VTAIL.n14 VTAIL.n13 585
R121 VTAIL.n71 VTAIL.n70 585
R122 VTAIL.n74 VTAIL.n73 585
R123 VTAIL.n72 VTAIL.n10 585
R124 VTAIL.n79 VTAIL.n9 585
R125 VTAIL.n81 VTAIL.n80 585
R126 VTAIL.n83 VTAIL.n82 585
R127 VTAIL.n6 VTAIL.n5 585
R128 VTAIL.n89 VTAIL.n88 585
R129 VTAIL.n91 VTAIL.n90 585
R130 VTAIL.n127 VTAIL.n126 585
R131 VTAIL.n124 VTAIL.n123 585
R132 VTAIL.n133 VTAIL.n132 585
R133 VTAIL.n135 VTAIL.n134 585
R134 VTAIL.n120 VTAIL.n119 585
R135 VTAIL.n141 VTAIL.n140 585
R136 VTAIL.n143 VTAIL.n142 585
R137 VTAIL.n116 VTAIL.n115 585
R138 VTAIL.n149 VTAIL.n148 585
R139 VTAIL.n151 VTAIL.n150 585
R140 VTAIL.n112 VTAIL.n111 585
R141 VTAIL.n157 VTAIL.n156 585
R142 VTAIL.n159 VTAIL.n158 585
R143 VTAIL.n108 VTAIL.n107 585
R144 VTAIL.n165 VTAIL.n164 585
R145 VTAIL.n168 VTAIL.n167 585
R146 VTAIL.n166 VTAIL.n104 585
R147 VTAIL.n173 VTAIL.n103 585
R148 VTAIL.n175 VTAIL.n174 585
R149 VTAIL.n177 VTAIL.n176 585
R150 VTAIL.n100 VTAIL.n99 585
R151 VTAIL.n183 VTAIL.n182 585
R152 VTAIL.n185 VTAIL.n184 585
R153 VTAIL.n223 VTAIL.n222 585
R154 VTAIL.n220 VTAIL.n219 585
R155 VTAIL.n229 VTAIL.n228 585
R156 VTAIL.n231 VTAIL.n230 585
R157 VTAIL.n216 VTAIL.n215 585
R158 VTAIL.n237 VTAIL.n236 585
R159 VTAIL.n239 VTAIL.n238 585
R160 VTAIL.n212 VTAIL.n211 585
R161 VTAIL.n245 VTAIL.n244 585
R162 VTAIL.n247 VTAIL.n246 585
R163 VTAIL.n208 VTAIL.n207 585
R164 VTAIL.n253 VTAIL.n252 585
R165 VTAIL.n255 VTAIL.n254 585
R166 VTAIL.n204 VTAIL.n203 585
R167 VTAIL.n261 VTAIL.n260 585
R168 VTAIL.n264 VTAIL.n263 585
R169 VTAIL.n262 VTAIL.n200 585
R170 VTAIL.n269 VTAIL.n199 585
R171 VTAIL.n271 VTAIL.n270 585
R172 VTAIL.n273 VTAIL.n272 585
R173 VTAIL.n196 VTAIL.n195 585
R174 VTAIL.n279 VTAIL.n278 585
R175 VTAIL.n281 VTAIL.n280 585
R176 VTAIL.n661 VTAIL.n660 585
R177 VTAIL.n659 VTAIL.n658 585
R178 VTAIL.n576 VTAIL.n575 585
R179 VTAIL.n653 VTAIL.n652 585
R180 VTAIL.n651 VTAIL.n650 585
R181 VTAIL.n649 VTAIL.n579 585
R182 VTAIL.n583 VTAIL.n580 585
R183 VTAIL.n644 VTAIL.n643 585
R184 VTAIL.n642 VTAIL.n641 585
R185 VTAIL.n585 VTAIL.n584 585
R186 VTAIL.n636 VTAIL.n635 585
R187 VTAIL.n634 VTAIL.n633 585
R188 VTAIL.n589 VTAIL.n588 585
R189 VTAIL.n628 VTAIL.n627 585
R190 VTAIL.n626 VTAIL.n625 585
R191 VTAIL.n593 VTAIL.n592 585
R192 VTAIL.n620 VTAIL.n619 585
R193 VTAIL.n618 VTAIL.n617 585
R194 VTAIL.n597 VTAIL.n596 585
R195 VTAIL.n612 VTAIL.n611 585
R196 VTAIL.n610 VTAIL.n609 585
R197 VTAIL.n601 VTAIL.n600 585
R198 VTAIL.n604 VTAIL.n603 585
R199 VTAIL.n565 VTAIL.n564 585
R200 VTAIL.n563 VTAIL.n562 585
R201 VTAIL.n480 VTAIL.n479 585
R202 VTAIL.n557 VTAIL.n556 585
R203 VTAIL.n555 VTAIL.n554 585
R204 VTAIL.n553 VTAIL.n483 585
R205 VTAIL.n487 VTAIL.n484 585
R206 VTAIL.n548 VTAIL.n547 585
R207 VTAIL.n546 VTAIL.n545 585
R208 VTAIL.n489 VTAIL.n488 585
R209 VTAIL.n540 VTAIL.n539 585
R210 VTAIL.n538 VTAIL.n537 585
R211 VTAIL.n493 VTAIL.n492 585
R212 VTAIL.n532 VTAIL.n531 585
R213 VTAIL.n530 VTAIL.n529 585
R214 VTAIL.n497 VTAIL.n496 585
R215 VTAIL.n524 VTAIL.n523 585
R216 VTAIL.n522 VTAIL.n521 585
R217 VTAIL.n501 VTAIL.n500 585
R218 VTAIL.n516 VTAIL.n515 585
R219 VTAIL.n514 VTAIL.n513 585
R220 VTAIL.n505 VTAIL.n504 585
R221 VTAIL.n508 VTAIL.n507 585
R222 VTAIL.n471 VTAIL.n470 585
R223 VTAIL.n469 VTAIL.n468 585
R224 VTAIL.n386 VTAIL.n385 585
R225 VTAIL.n463 VTAIL.n462 585
R226 VTAIL.n461 VTAIL.n460 585
R227 VTAIL.n459 VTAIL.n389 585
R228 VTAIL.n393 VTAIL.n390 585
R229 VTAIL.n454 VTAIL.n453 585
R230 VTAIL.n452 VTAIL.n451 585
R231 VTAIL.n395 VTAIL.n394 585
R232 VTAIL.n446 VTAIL.n445 585
R233 VTAIL.n444 VTAIL.n443 585
R234 VTAIL.n399 VTAIL.n398 585
R235 VTAIL.n438 VTAIL.n437 585
R236 VTAIL.n436 VTAIL.n435 585
R237 VTAIL.n403 VTAIL.n402 585
R238 VTAIL.n430 VTAIL.n429 585
R239 VTAIL.n428 VTAIL.n427 585
R240 VTAIL.n407 VTAIL.n406 585
R241 VTAIL.n422 VTAIL.n421 585
R242 VTAIL.n420 VTAIL.n419 585
R243 VTAIL.n411 VTAIL.n410 585
R244 VTAIL.n414 VTAIL.n413 585
R245 VTAIL.n375 VTAIL.n374 585
R246 VTAIL.n373 VTAIL.n372 585
R247 VTAIL.n290 VTAIL.n289 585
R248 VTAIL.n367 VTAIL.n366 585
R249 VTAIL.n365 VTAIL.n364 585
R250 VTAIL.n363 VTAIL.n293 585
R251 VTAIL.n297 VTAIL.n294 585
R252 VTAIL.n358 VTAIL.n357 585
R253 VTAIL.n356 VTAIL.n355 585
R254 VTAIL.n299 VTAIL.n298 585
R255 VTAIL.n350 VTAIL.n349 585
R256 VTAIL.n348 VTAIL.n347 585
R257 VTAIL.n303 VTAIL.n302 585
R258 VTAIL.n342 VTAIL.n341 585
R259 VTAIL.n340 VTAIL.n339 585
R260 VTAIL.n307 VTAIL.n306 585
R261 VTAIL.n334 VTAIL.n333 585
R262 VTAIL.n332 VTAIL.n331 585
R263 VTAIL.n311 VTAIL.n310 585
R264 VTAIL.n326 VTAIL.n325 585
R265 VTAIL.n324 VTAIL.n323 585
R266 VTAIL.n315 VTAIL.n314 585
R267 VTAIL.n318 VTAIL.n317 585
R268 VTAIL.t6 VTAIL.n602 327.466
R269 VTAIL.t7 VTAIL.n506 327.466
R270 VTAIL.t14 VTAIL.n412 327.466
R271 VTAIL.t15 VTAIL.n316 327.466
R272 VTAIL.t8 VTAIL.n695 327.466
R273 VTAIL.t13 VTAIL.n31 327.466
R274 VTAIL.t1 VTAIL.n125 327.466
R275 VTAIL.t5 VTAIL.n221 327.466
R276 VTAIL.n696 VTAIL.n693 171.744
R277 VTAIL.n703 VTAIL.n693 171.744
R278 VTAIL.n704 VTAIL.n703 171.744
R279 VTAIL.n704 VTAIL.n689 171.744
R280 VTAIL.n711 VTAIL.n689 171.744
R281 VTAIL.n712 VTAIL.n711 171.744
R282 VTAIL.n712 VTAIL.n685 171.744
R283 VTAIL.n719 VTAIL.n685 171.744
R284 VTAIL.n720 VTAIL.n719 171.744
R285 VTAIL.n720 VTAIL.n681 171.744
R286 VTAIL.n727 VTAIL.n681 171.744
R287 VTAIL.n728 VTAIL.n727 171.744
R288 VTAIL.n728 VTAIL.n677 171.744
R289 VTAIL.n735 VTAIL.n677 171.744
R290 VTAIL.n737 VTAIL.n735 171.744
R291 VTAIL.n737 VTAIL.n736 171.744
R292 VTAIL.n736 VTAIL.n673 171.744
R293 VTAIL.n745 VTAIL.n673 171.744
R294 VTAIL.n746 VTAIL.n745 171.744
R295 VTAIL.n746 VTAIL.n669 171.744
R296 VTAIL.n753 VTAIL.n669 171.744
R297 VTAIL.n754 VTAIL.n753 171.744
R298 VTAIL.n32 VTAIL.n29 171.744
R299 VTAIL.n39 VTAIL.n29 171.744
R300 VTAIL.n40 VTAIL.n39 171.744
R301 VTAIL.n40 VTAIL.n25 171.744
R302 VTAIL.n47 VTAIL.n25 171.744
R303 VTAIL.n48 VTAIL.n47 171.744
R304 VTAIL.n48 VTAIL.n21 171.744
R305 VTAIL.n55 VTAIL.n21 171.744
R306 VTAIL.n56 VTAIL.n55 171.744
R307 VTAIL.n56 VTAIL.n17 171.744
R308 VTAIL.n63 VTAIL.n17 171.744
R309 VTAIL.n64 VTAIL.n63 171.744
R310 VTAIL.n64 VTAIL.n13 171.744
R311 VTAIL.n71 VTAIL.n13 171.744
R312 VTAIL.n73 VTAIL.n71 171.744
R313 VTAIL.n73 VTAIL.n72 171.744
R314 VTAIL.n72 VTAIL.n9 171.744
R315 VTAIL.n81 VTAIL.n9 171.744
R316 VTAIL.n82 VTAIL.n81 171.744
R317 VTAIL.n82 VTAIL.n5 171.744
R318 VTAIL.n89 VTAIL.n5 171.744
R319 VTAIL.n90 VTAIL.n89 171.744
R320 VTAIL.n126 VTAIL.n123 171.744
R321 VTAIL.n133 VTAIL.n123 171.744
R322 VTAIL.n134 VTAIL.n133 171.744
R323 VTAIL.n134 VTAIL.n119 171.744
R324 VTAIL.n141 VTAIL.n119 171.744
R325 VTAIL.n142 VTAIL.n141 171.744
R326 VTAIL.n142 VTAIL.n115 171.744
R327 VTAIL.n149 VTAIL.n115 171.744
R328 VTAIL.n150 VTAIL.n149 171.744
R329 VTAIL.n150 VTAIL.n111 171.744
R330 VTAIL.n157 VTAIL.n111 171.744
R331 VTAIL.n158 VTAIL.n157 171.744
R332 VTAIL.n158 VTAIL.n107 171.744
R333 VTAIL.n165 VTAIL.n107 171.744
R334 VTAIL.n167 VTAIL.n165 171.744
R335 VTAIL.n167 VTAIL.n166 171.744
R336 VTAIL.n166 VTAIL.n103 171.744
R337 VTAIL.n175 VTAIL.n103 171.744
R338 VTAIL.n176 VTAIL.n175 171.744
R339 VTAIL.n176 VTAIL.n99 171.744
R340 VTAIL.n183 VTAIL.n99 171.744
R341 VTAIL.n184 VTAIL.n183 171.744
R342 VTAIL.n222 VTAIL.n219 171.744
R343 VTAIL.n229 VTAIL.n219 171.744
R344 VTAIL.n230 VTAIL.n229 171.744
R345 VTAIL.n230 VTAIL.n215 171.744
R346 VTAIL.n237 VTAIL.n215 171.744
R347 VTAIL.n238 VTAIL.n237 171.744
R348 VTAIL.n238 VTAIL.n211 171.744
R349 VTAIL.n245 VTAIL.n211 171.744
R350 VTAIL.n246 VTAIL.n245 171.744
R351 VTAIL.n246 VTAIL.n207 171.744
R352 VTAIL.n253 VTAIL.n207 171.744
R353 VTAIL.n254 VTAIL.n253 171.744
R354 VTAIL.n254 VTAIL.n203 171.744
R355 VTAIL.n261 VTAIL.n203 171.744
R356 VTAIL.n263 VTAIL.n261 171.744
R357 VTAIL.n263 VTAIL.n262 171.744
R358 VTAIL.n262 VTAIL.n199 171.744
R359 VTAIL.n271 VTAIL.n199 171.744
R360 VTAIL.n272 VTAIL.n271 171.744
R361 VTAIL.n272 VTAIL.n195 171.744
R362 VTAIL.n279 VTAIL.n195 171.744
R363 VTAIL.n280 VTAIL.n279 171.744
R364 VTAIL.n660 VTAIL.n659 171.744
R365 VTAIL.n659 VTAIL.n575 171.744
R366 VTAIL.n652 VTAIL.n575 171.744
R367 VTAIL.n652 VTAIL.n651 171.744
R368 VTAIL.n651 VTAIL.n579 171.744
R369 VTAIL.n583 VTAIL.n579 171.744
R370 VTAIL.n643 VTAIL.n583 171.744
R371 VTAIL.n643 VTAIL.n642 171.744
R372 VTAIL.n642 VTAIL.n584 171.744
R373 VTAIL.n635 VTAIL.n584 171.744
R374 VTAIL.n635 VTAIL.n634 171.744
R375 VTAIL.n634 VTAIL.n588 171.744
R376 VTAIL.n627 VTAIL.n588 171.744
R377 VTAIL.n627 VTAIL.n626 171.744
R378 VTAIL.n626 VTAIL.n592 171.744
R379 VTAIL.n619 VTAIL.n592 171.744
R380 VTAIL.n619 VTAIL.n618 171.744
R381 VTAIL.n618 VTAIL.n596 171.744
R382 VTAIL.n611 VTAIL.n596 171.744
R383 VTAIL.n611 VTAIL.n610 171.744
R384 VTAIL.n610 VTAIL.n600 171.744
R385 VTAIL.n603 VTAIL.n600 171.744
R386 VTAIL.n564 VTAIL.n563 171.744
R387 VTAIL.n563 VTAIL.n479 171.744
R388 VTAIL.n556 VTAIL.n479 171.744
R389 VTAIL.n556 VTAIL.n555 171.744
R390 VTAIL.n555 VTAIL.n483 171.744
R391 VTAIL.n487 VTAIL.n483 171.744
R392 VTAIL.n547 VTAIL.n487 171.744
R393 VTAIL.n547 VTAIL.n546 171.744
R394 VTAIL.n546 VTAIL.n488 171.744
R395 VTAIL.n539 VTAIL.n488 171.744
R396 VTAIL.n539 VTAIL.n538 171.744
R397 VTAIL.n538 VTAIL.n492 171.744
R398 VTAIL.n531 VTAIL.n492 171.744
R399 VTAIL.n531 VTAIL.n530 171.744
R400 VTAIL.n530 VTAIL.n496 171.744
R401 VTAIL.n523 VTAIL.n496 171.744
R402 VTAIL.n523 VTAIL.n522 171.744
R403 VTAIL.n522 VTAIL.n500 171.744
R404 VTAIL.n515 VTAIL.n500 171.744
R405 VTAIL.n515 VTAIL.n514 171.744
R406 VTAIL.n514 VTAIL.n504 171.744
R407 VTAIL.n507 VTAIL.n504 171.744
R408 VTAIL.n470 VTAIL.n469 171.744
R409 VTAIL.n469 VTAIL.n385 171.744
R410 VTAIL.n462 VTAIL.n385 171.744
R411 VTAIL.n462 VTAIL.n461 171.744
R412 VTAIL.n461 VTAIL.n389 171.744
R413 VTAIL.n393 VTAIL.n389 171.744
R414 VTAIL.n453 VTAIL.n393 171.744
R415 VTAIL.n453 VTAIL.n452 171.744
R416 VTAIL.n452 VTAIL.n394 171.744
R417 VTAIL.n445 VTAIL.n394 171.744
R418 VTAIL.n445 VTAIL.n444 171.744
R419 VTAIL.n444 VTAIL.n398 171.744
R420 VTAIL.n437 VTAIL.n398 171.744
R421 VTAIL.n437 VTAIL.n436 171.744
R422 VTAIL.n436 VTAIL.n402 171.744
R423 VTAIL.n429 VTAIL.n402 171.744
R424 VTAIL.n429 VTAIL.n428 171.744
R425 VTAIL.n428 VTAIL.n406 171.744
R426 VTAIL.n421 VTAIL.n406 171.744
R427 VTAIL.n421 VTAIL.n420 171.744
R428 VTAIL.n420 VTAIL.n410 171.744
R429 VTAIL.n413 VTAIL.n410 171.744
R430 VTAIL.n374 VTAIL.n373 171.744
R431 VTAIL.n373 VTAIL.n289 171.744
R432 VTAIL.n366 VTAIL.n289 171.744
R433 VTAIL.n366 VTAIL.n365 171.744
R434 VTAIL.n365 VTAIL.n293 171.744
R435 VTAIL.n297 VTAIL.n293 171.744
R436 VTAIL.n357 VTAIL.n297 171.744
R437 VTAIL.n357 VTAIL.n356 171.744
R438 VTAIL.n356 VTAIL.n298 171.744
R439 VTAIL.n349 VTAIL.n298 171.744
R440 VTAIL.n349 VTAIL.n348 171.744
R441 VTAIL.n348 VTAIL.n302 171.744
R442 VTAIL.n341 VTAIL.n302 171.744
R443 VTAIL.n341 VTAIL.n340 171.744
R444 VTAIL.n340 VTAIL.n306 171.744
R445 VTAIL.n333 VTAIL.n306 171.744
R446 VTAIL.n333 VTAIL.n332 171.744
R447 VTAIL.n332 VTAIL.n310 171.744
R448 VTAIL.n325 VTAIL.n310 171.744
R449 VTAIL.n325 VTAIL.n324 171.744
R450 VTAIL.n324 VTAIL.n314 171.744
R451 VTAIL.n317 VTAIL.n314 171.744
R452 VTAIL.n696 VTAIL.t8 85.8723
R453 VTAIL.n32 VTAIL.t13 85.8723
R454 VTAIL.n126 VTAIL.t1 85.8723
R455 VTAIL.n222 VTAIL.t5 85.8723
R456 VTAIL.n603 VTAIL.t6 85.8723
R457 VTAIL.n507 VTAIL.t7 85.8723
R458 VTAIL.n413 VTAIL.t14 85.8723
R459 VTAIL.n317 VTAIL.t15 85.8723
R460 VTAIL.n571 VTAIL.n570 51.5496
R461 VTAIL.n381 VTAIL.n380 51.5496
R462 VTAIL.n1 VTAIL.n0 51.5494
R463 VTAIL.n191 VTAIL.n190 51.5494
R464 VTAIL.n759 VTAIL.n758 31.0217
R465 VTAIL.n95 VTAIL.n94 31.0217
R466 VTAIL.n189 VTAIL.n188 31.0217
R467 VTAIL.n285 VTAIL.n284 31.0217
R468 VTAIL.n665 VTAIL.n664 31.0217
R469 VTAIL.n569 VTAIL.n568 31.0217
R470 VTAIL.n475 VTAIL.n474 31.0217
R471 VTAIL.n379 VTAIL.n378 31.0217
R472 VTAIL.n759 VTAIL.n665 28.2721
R473 VTAIL.n379 VTAIL.n285 28.2721
R474 VTAIL.n697 VTAIL.n695 16.3895
R475 VTAIL.n33 VTAIL.n31 16.3895
R476 VTAIL.n127 VTAIL.n125 16.3895
R477 VTAIL.n223 VTAIL.n221 16.3895
R478 VTAIL.n604 VTAIL.n602 16.3895
R479 VTAIL.n508 VTAIL.n506 16.3895
R480 VTAIL.n414 VTAIL.n412 16.3895
R481 VTAIL.n318 VTAIL.n316 16.3895
R482 VTAIL.n744 VTAIL.n743 13.1884
R483 VTAIL.n80 VTAIL.n79 13.1884
R484 VTAIL.n174 VTAIL.n173 13.1884
R485 VTAIL.n270 VTAIL.n269 13.1884
R486 VTAIL.n650 VTAIL.n649 13.1884
R487 VTAIL.n554 VTAIL.n553 13.1884
R488 VTAIL.n460 VTAIL.n459 13.1884
R489 VTAIL.n364 VTAIL.n363 13.1884
R490 VTAIL.n698 VTAIL.n694 12.8005
R491 VTAIL.n742 VTAIL.n674 12.8005
R492 VTAIL.n747 VTAIL.n672 12.8005
R493 VTAIL.n34 VTAIL.n30 12.8005
R494 VTAIL.n78 VTAIL.n10 12.8005
R495 VTAIL.n83 VTAIL.n8 12.8005
R496 VTAIL.n128 VTAIL.n124 12.8005
R497 VTAIL.n172 VTAIL.n104 12.8005
R498 VTAIL.n177 VTAIL.n102 12.8005
R499 VTAIL.n224 VTAIL.n220 12.8005
R500 VTAIL.n268 VTAIL.n200 12.8005
R501 VTAIL.n273 VTAIL.n198 12.8005
R502 VTAIL.n653 VTAIL.n578 12.8005
R503 VTAIL.n648 VTAIL.n580 12.8005
R504 VTAIL.n605 VTAIL.n601 12.8005
R505 VTAIL.n557 VTAIL.n482 12.8005
R506 VTAIL.n552 VTAIL.n484 12.8005
R507 VTAIL.n509 VTAIL.n505 12.8005
R508 VTAIL.n463 VTAIL.n388 12.8005
R509 VTAIL.n458 VTAIL.n390 12.8005
R510 VTAIL.n415 VTAIL.n411 12.8005
R511 VTAIL.n367 VTAIL.n292 12.8005
R512 VTAIL.n362 VTAIL.n294 12.8005
R513 VTAIL.n319 VTAIL.n315 12.8005
R514 VTAIL.n702 VTAIL.n701 12.0247
R515 VTAIL.n739 VTAIL.n738 12.0247
R516 VTAIL.n748 VTAIL.n670 12.0247
R517 VTAIL.n38 VTAIL.n37 12.0247
R518 VTAIL.n75 VTAIL.n74 12.0247
R519 VTAIL.n84 VTAIL.n6 12.0247
R520 VTAIL.n132 VTAIL.n131 12.0247
R521 VTAIL.n169 VTAIL.n168 12.0247
R522 VTAIL.n178 VTAIL.n100 12.0247
R523 VTAIL.n228 VTAIL.n227 12.0247
R524 VTAIL.n265 VTAIL.n264 12.0247
R525 VTAIL.n274 VTAIL.n196 12.0247
R526 VTAIL.n654 VTAIL.n576 12.0247
R527 VTAIL.n645 VTAIL.n644 12.0247
R528 VTAIL.n609 VTAIL.n608 12.0247
R529 VTAIL.n558 VTAIL.n480 12.0247
R530 VTAIL.n549 VTAIL.n548 12.0247
R531 VTAIL.n513 VTAIL.n512 12.0247
R532 VTAIL.n464 VTAIL.n386 12.0247
R533 VTAIL.n455 VTAIL.n454 12.0247
R534 VTAIL.n419 VTAIL.n418 12.0247
R535 VTAIL.n368 VTAIL.n290 12.0247
R536 VTAIL.n359 VTAIL.n358 12.0247
R537 VTAIL.n323 VTAIL.n322 12.0247
R538 VTAIL.n705 VTAIL.n692 11.249
R539 VTAIL.n734 VTAIL.n676 11.249
R540 VTAIL.n752 VTAIL.n751 11.249
R541 VTAIL.n41 VTAIL.n28 11.249
R542 VTAIL.n70 VTAIL.n12 11.249
R543 VTAIL.n88 VTAIL.n87 11.249
R544 VTAIL.n135 VTAIL.n122 11.249
R545 VTAIL.n164 VTAIL.n106 11.249
R546 VTAIL.n182 VTAIL.n181 11.249
R547 VTAIL.n231 VTAIL.n218 11.249
R548 VTAIL.n260 VTAIL.n202 11.249
R549 VTAIL.n278 VTAIL.n277 11.249
R550 VTAIL.n658 VTAIL.n657 11.249
R551 VTAIL.n641 VTAIL.n582 11.249
R552 VTAIL.n612 VTAIL.n599 11.249
R553 VTAIL.n562 VTAIL.n561 11.249
R554 VTAIL.n545 VTAIL.n486 11.249
R555 VTAIL.n516 VTAIL.n503 11.249
R556 VTAIL.n468 VTAIL.n467 11.249
R557 VTAIL.n451 VTAIL.n392 11.249
R558 VTAIL.n422 VTAIL.n409 11.249
R559 VTAIL.n372 VTAIL.n371 11.249
R560 VTAIL.n355 VTAIL.n296 11.249
R561 VTAIL.n326 VTAIL.n313 11.249
R562 VTAIL.n706 VTAIL.n690 10.4732
R563 VTAIL.n733 VTAIL.n678 10.4732
R564 VTAIL.n755 VTAIL.n668 10.4732
R565 VTAIL.n42 VTAIL.n26 10.4732
R566 VTAIL.n69 VTAIL.n14 10.4732
R567 VTAIL.n91 VTAIL.n4 10.4732
R568 VTAIL.n136 VTAIL.n120 10.4732
R569 VTAIL.n163 VTAIL.n108 10.4732
R570 VTAIL.n185 VTAIL.n98 10.4732
R571 VTAIL.n232 VTAIL.n216 10.4732
R572 VTAIL.n259 VTAIL.n204 10.4732
R573 VTAIL.n281 VTAIL.n194 10.4732
R574 VTAIL.n661 VTAIL.n574 10.4732
R575 VTAIL.n640 VTAIL.n585 10.4732
R576 VTAIL.n613 VTAIL.n597 10.4732
R577 VTAIL.n565 VTAIL.n478 10.4732
R578 VTAIL.n544 VTAIL.n489 10.4732
R579 VTAIL.n517 VTAIL.n501 10.4732
R580 VTAIL.n471 VTAIL.n384 10.4732
R581 VTAIL.n450 VTAIL.n395 10.4732
R582 VTAIL.n423 VTAIL.n407 10.4732
R583 VTAIL.n375 VTAIL.n288 10.4732
R584 VTAIL.n354 VTAIL.n299 10.4732
R585 VTAIL.n327 VTAIL.n311 10.4732
R586 VTAIL.n710 VTAIL.n709 9.69747
R587 VTAIL.n730 VTAIL.n729 9.69747
R588 VTAIL.n756 VTAIL.n666 9.69747
R589 VTAIL.n46 VTAIL.n45 9.69747
R590 VTAIL.n66 VTAIL.n65 9.69747
R591 VTAIL.n92 VTAIL.n2 9.69747
R592 VTAIL.n140 VTAIL.n139 9.69747
R593 VTAIL.n160 VTAIL.n159 9.69747
R594 VTAIL.n186 VTAIL.n96 9.69747
R595 VTAIL.n236 VTAIL.n235 9.69747
R596 VTAIL.n256 VTAIL.n255 9.69747
R597 VTAIL.n282 VTAIL.n192 9.69747
R598 VTAIL.n662 VTAIL.n572 9.69747
R599 VTAIL.n637 VTAIL.n636 9.69747
R600 VTAIL.n617 VTAIL.n616 9.69747
R601 VTAIL.n566 VTAIL.n476 9.69747
R602 VTAIL.n541 VTAIL.n540 9.69747
R603 VTAIL.n521 VTAIL.n520 9.69747
R604 VTAIL.n472 VTAIL.n382 9.69747
R605 VTAIL.n447 VTAIL.n446 9.69747
R606 VTAIL.n427 VTAIL.n426 9.69747
R607 VTAIL.n376 VTAIL.n286 9.69747
R608 VTAIL.n351 VTAIL.n350 9.69747
R609 VTAIL.n331 VTAIL.n330 9.69747
R610 VTAIL.n758 VTAIL.n757 9.45567
R611 VTAIL.n94 VTAIL.n93 9.45567
R612 VTAIL.n188 VTAIL.n187 9.45567
R613 VTAIL.n284 VTAIL.n283 9.45567
R614 VTAIL.n664 VTAIL.n663 9.45567
R615 VTAIL.n568 VTAIL.n567 9.45567
R616 VTAIL.n474 VTAIL.n473 9.45567
R617 VTAIL.n378 VTAIL.n377 9.45567
R618 VTAIL.n757 VTAIL.n756 9.3005
R619 VTAIL.n668 VTAIL.n667 9.3005
R620 VTAIL.n751 VTAIL.n750 9.3005
R621 VTAIL.n749 VTAIL.n748 9.3005
R622 VTAIL.n672 VTAIL.n671 9.3005
R623 VTAIL.n717 VTAIL.n716 9.3005
R624 VTAIL.n715 VTAIL.n714 9.3005
R625 VTAIL.n688 VTAIL.n687 9.3005
R626 VTAIL.n709 VTAIL.n708 9.3005
R627 VTAIL.n707 VTAIL.n706 9.3005
R628 VTAIL.n692 VTAIL.n691 9.3005
R629 VTAIL.n701 VTAIL.n700 9.3005
R630 VTAIL.n699 VTAIL.n698 9.3005
R631 VTAIL.n684 VTAIL.n683 9.3005
R632 VTAIL.n723 VTAIL.n722 9.3005
R633 VTAIL.n725 VTAIL.n724 9.3005
R634 VTAIL.n680 VTAIL.n679 9.3005
R635 VTAIL.n731 VTAIL.n730 9.3005
R636 VTAIL.n733 VTAIL.n732 9.3005
R637 VTAIL.n676 VTAIL.n675 9.3005
R638 VTAIL.n740 VTAIL.n739 9.3005
R639 VTAIL.n742 VTAIL.n741 9.3005
R640 VTAIL.n93 VTAIL.n92 9.3005
R641 VTAIL.n4 VTAIL.n3 9.3005
R642 VTAIL.n87 VTAIL.n86 9.3005
R643 VTAIL.n85 VTAIL.n84 9.3005
R644 VTAIL.n8 VTAIL.n7 9.3005
R645 VTAIL.n53 VTAIL.n52 9.3005
R646 VTAIL.n51 VTAIL.n50 9.3005
R647 VTAIL.n24 VTAIL.n23 9.3005
R648 VTAIL.n45 VTAIL.n44 9.3005
R649 VTAIL.n43 VTAIL.n42 9.3005
R650 VTAIL.n28 VTAIL.n27 9.3005
R651 VTAIL.n37 VTAIL.n36 9.3005
R652 VTAIL.n35 VTAIL.n34 9.3005
R653 VTAIL.n20 VTAIL.n19 9.3005
R654 VTAIL.n59 VTAIL.n58 9.3005
R655 VTAIL.n61 VTAIL.n60 9.3005
R656 VTAIL.n16 VTAIL.n15 9.3005
R657 VTAIL.n67 VTAIL.n66 9.3005
R658 VTAIL.n69 VTAIL.n68 9.3005
R659 VTAIL.n12 VTAIL.n11 9.3005
R660 VTAIL.n76 VTAIL.n75 9.3005
R661 VTAIL.n78 VTAIL.n77 9.3005
R662 VTAIL.n187 VTAIL.n186 9.3005
R663 VTAIL.n98 VTAIL.n97 9.3005
R664 VTAIL.n181 VTAIL.n180 9.3005
R665 VTAIL.n179 VTAIL.n178 9.3005
R666 VTAIL.n102 VTAIL.n101 9.3005
R667 VTAIL.n147 VTAIL.n146 9.3005
R668 VTAIL.n145 VTAIL.n144 9.3005
R669 VTAIL.n118 VTAIL.n117 9.3005
R670 VTAIL.n139 VTAIL.n138 9.3005
R671 VTAIL.n137 VTAIL.n136 9.3005
R672 VTAIL.n122 VTAIL.n121 9.3005
R673 VTAIL.n131 VTAIL.n130 9.3005
R674 VTAIL.n129 VTAIL.n128 9.3005
R675 VTAIL.n114 VTAIL.n113 9.3005
R676 VTAIL.n153 VTAIL.n152 9.3005
R677 VTAIL.n155 VTAIL.n154 9.3005
R678 VTAIL.n110 VTAIL.n109 9.3005
R679 VTAIL.n161 VTAIL.n160 9.3005
R680 VTAIL.n163 VTAIL.n162 9.3005
R681 VTAIL.n106 VTAIL.n105 9.3005
R682 VTAIL.n170 VTAIL.n169 9.3005
R683 VTAIL.n172 VTAIL.n171 9.3005
R684 VTAIL.n283 VTAIL.n282 9.3005
R685 VTAIL.n194 VTAIL.n193 9.3005
R686 VTAIL.n277 VTAIL.n276 9.3005
R687 VTAIL.n275 VTAIL.n274 9.3005
R688 VTAIL.n198 VTAIL.n197 9.3005
R689 VTAIL.n243 VTAIL.n242 9.3005
R690 VTAIL.n241 VTAIL.n240 9.3005
R691 VTAIL.n214 VTAIL.n213 9.3005
R692 VTAIL.n235 VTAIL.n234 9.3005
R693 VTAIL.n233 VTAIL.n232 9.3005
R694 VTAIL.n218 VTAIL.n217 9.3005
R695 VTAIL.n227 VTAIL.n226 9.3005
R696 VTAIL.n225 VTAIL.n224 9.3005
R697 VTAIL.n210 VTAIL.n209 9.3005
R698 VTAIL.n249 VTAIL.n248 9.3005
R699 VTAIL.n251 VTAIL.n250 9.3005
R700 VTAIL.n206 VTAIL.n205 9.3005
R701 VTAIL.n257 VTAIL.n256 9.3005
R702 VTAIL.n259 VTAIL.n258 9.3005
R703 VTAIL.n202 VTAIL.n201 9.3005
R704 VTAIL.n266 VTAIL.n265 9.3005
R705 VTAIL.n268 VTAIL.n267 9.3005
R706 VTAIL.n630 VTAIL.n629 9.3005
R707 VTAIL.n632 VTAIL.n631 9.3005
R708 VTAIL.n587 VTAIL.n586 9.3005
R709 VTAIL.n638 VTAIL.n637 9.3005
R710 VTAIL.n640 VTAIL.n639 9.3005
R711 VTAIL.n582 VTAIL.n581 9.3005
R712 VTAIL.n646 VTAIL.n645 9.3005
R713 VTAIL.n648 VTAIL.n647 9.3005
R714 VTAIL.n663 VTAIL.n662 9.3005
R715 VTAIL.n574 VTAIL.n573 9.3005
R716 VTAIL.n657 VTAIL.n656 9.3005
R717 VTAIL.n655 VTAIL.n654 9.3005
R718 VTAIL.n578 VTAIL.n577 9.3005
R719 VTAIL.n591 VTAIL.n590 9.3005
R720 VTAIL.n624 VTAIL.n623 9.3005
R721 VTAIL.n622 VTAIL.n621 9.3005
R722 VTAIL.n595 VTAIL.n594 9.3005
R723 VTAIL.n616 VTAIL.n615 9.3005
R724 VTAIL.n614 VTAIL.n613 9.3005
R725 VTAIL.n599 VTAIL.n598 9.3005
R726 VTAIL.n608 VTAIL.n607 9.3005
R727 VTAIL.n606 VTAIL.n605 9.3005
R728 VTAIL.n534 VTAIL.n533 9.3005
R729 VTAIL.n536 VTAIL.n535 9.3005
R730 VTAIL.n491 VTAIL.n490 9.3005
R731 VTAIL.n542 VTAIL.n541 9.3005
R732 VTAIL.n544 VTAIL.n543 9.3005
R733 VTAIL.n486 VTAIL.n485 9.3005
R734 VTAIL.n550 VTAIL.n549 9.3005
R735 VTAIL.n552 VTAIL.n551 9.3005
R736 VTAIL.n567 VTAIL.n566 9.3005
R737 VTAIL.n478 VTAIL.n477 9.3005
R738 VTAIL.n561 VTAIL.n560 9.3005
R739 VTAIL.n559 VTAIL.n558 9.3005
R740 VTAIL.n482 VTAIL.n481 9.3005
R741 VTAIL.n495 VTAIL.n494 9.3005
R742 VTAIL.n528 VTAIL.n527 9.3005
R743 VTAIL.n526 VTAIL.n525 9.3005
R744 VTAIL.n499 VTAIL.n498 9.3005
R745 VTAIL.n520 VTAIL.n519 9.3005
R746 VTAIL.n518 VTAIL.n517 9.3005
R747 VTAIL.n503 VTAIL.n502 9.3005
R748 VTAIL.n512 VTAIL.n511 9.3005
R749 VTAIL.n510 VTAIL.n509 9.3005
R750 VTAIL.n440 VTAIL.n439 9.3005
R751 VTAIL.n442 VTAIL.n441 9.3005
R752 VTAIL.n397 VTAIL.n396 9.3005
R753 VTAIL.n448 VTAIL.n447 9.3005
R754 VTAIL.n450 VTAIL.n449 9.3005
R755 VTAIL.n392 VTAIL.n391 9.3005
R756 VTAIL.n456 VTAIL.n455 9.3005
R757 VTAIL.n458 VTAIL.n457 9.3005
R758 VTAIL.n473 VTAIL.n472 9.3005
R759 VTAIL.n384 VTAIL.n383 9.3005
R760 VTAIL.n467 VTAIL.n466 9.3005
R761 VTAIL.n465 VTAIL.n464 9.3005
R762 VTAIL.n388 VTAIL.n387 9.3005
R763 VTAIL.n401 VTAIL.n400 9.3005
R764 VTAIL.n434 VTAIL.n433 9.3005
R765 VTAIL.n432 VTAIL.n431 9.3005
R766 VTAIL.n405 VTAIL.n404 9.3005
R767 VTAIL.n426 VTAIL.n425 9.3005
R768 VTAIL.n424 VTAIL.n423 9.3005
R769 VTAIL.n409 VTAIL.n408 9.3005
R770 VTAIL.n418 VTAIL.n417 9.3005
R771 VTAIL.n416 VTAIL.n415 9.3005
R772 VTAIL.n344 VTAIL.n343 9.3005
R773 VTAIL.n346 VTAIL.n345 9.3005
R774 VTAIL.n301 VTAIL.n300 9.3005
R775 VTAIL.n352 VTAIL.n351 9.3005
R776 VTAIL.n354 VTAIL.n353 9.3005
R777 VTAIL.n296 VTAIL.n295 9.3005
R778 VTAIL.n360 VTAIL.n359 9.3005
R779 VTAIL.n362 VTAIL.n361 9.3005
R780 VTAIL.n377 VTAIL.n376 9.3005
R781 VTAIL.n288 VTAIL.n287 9.3005
R782 VTAIL.n371 VTAIL.n370 9.3005
R783 VTAIL.n369 VTAIL.n368 9.3005
R784 VTAIL.n292 VTAIL.n291 9.3005
R785 VTAIL.n305 VTAIL.n304 9.3005
R786 VTAIL.n338 VTAIL.n337 9.3005
R787 VTAIL.n336 VTAIL.n335 9.3005
R788 VTAIL.n309 VTAIL.n308 9.3005
R789 VTAIL.n330 VTAIL.n329 9.3005
R790 VTAIL.n328 VTAIL.n327 9.3005
R791 VTAIL.n313 VTAIL.n312 9.3005
R792 VTAIL.n322 VTAIL.n321 9.3005
R793 VTAIL.n320 VTAIL.n319 9.3005
R794 VTAIL.n713 VTAIL.n688 8.92171
R795 VTAIL.n726 VTAIL.n680 8.92171
R796 VTAIL.n49 VTAIL.n24 8.92171
R797 VTAIL.n62 VTAIL.n16 8.92171
R798 VTAIL.n143 VTAIL.n118 8.92171
R799 VTAIL.n156 VTAIL.n110 8.92171
R800 VTAIL.n239 VTAIL.n214 8.92171
R801 VTAIL.n252 VTAIL.n206 8.92171
R802 VTAIL.n633 VTAIL.n587 8.92171
R803 VTAIL.n620 VTAIL.n595 8.92171
R804 VTAIL.n537 VTAIL.n491 8.92171
R805 VTAIL.n524 VTAIL.n499 8.92171
R806 VTAIL.n443 VTAIL.n397 8.92171
R807 VTAIL.n430 VTAIL.n405 8.92171
R808 VTAIL.n347 VTAIL.n301 8.92171
R809 VTAIL.n334 VTAIL.n309 8.92171
R810 VTAIL.n714 VTAIL.n686 8.14595
R811 VTAIL.n725 VTAIL.n682 8.14595
R812 VTAIL.n50 VTAIL.n22 8.14595
R813 VTAIL.n61 VTAIL.n18 8.14595
R814 VTAIL.n144 VTAIL.n116 8.14595
R815 VTAIL.n155 VTAIL.n112 8.14595
R816 VTAIL.n240 VTAIL.n212 8.14595
R817 VTAIL.n251 VTAIL.n208 8.14595
R818 VTAIL.n632 VTAIL.n589 8.14595
R819 VTAIL.n621 VTAIL.n593 8.14595
R820 VTAIL.n536 VTAIL.n493 8.14595
R821 VTAIL.n525 VTAIL.n497 8.14595
R822 VTAIL.n442 VTAIL.n399 8.14595
R823 VTAIL.n431 VTAIL.n403 8.14595
R824 VTAIL.n346 VTAIL.n303 8.14595
R825 VTAIL.n335 VTAIL.n307 8.14595
R826 VTAIL.n718 VTAIL.n717 7.3702
R827 VTAIL.n722 VTAIL.n721 7.3702
R828 VTAIL.n54 VTAIL.n53 7.3702
R829 VTAIL.n58 VTAIL.n57 7.3702
R830 VTAIL.n148 VTAIL.n147 7.3702
R831 VTAIL.n152 VTAIL.n151 7.3702
R832 VTAIL.n244 VTAIL.n243 7.3702
R833 VTAIL.n248 VTAIL.n247 7.3702
R834 VTAIL.n629 VTAIL.n628 7.3702
R835 VTAIL.n625 VTAIL.n624 7.3702
R836 VTAIL.n533 VTAIL.n532 7.3702
R837 VTAIL.n529 VTAIL.n528 7.3702
R838 VTAIL.n439 VTAIL.n438 7.3702
R839 VTAIL.n435 VTAIL.n434 7.3702
R840 VTAIL.n343 VTAIL.n342 7.3702
R841 VTAIL.n339 VTAIL.n338 7.3702
R842 VTAIL.n718 VTAIL.n684 6.59444
R843 VTAIL.n721 VTAIL.n684 6.59444
R844 VTAIL.n54 VTAIL.n20 6.59444
R845 VTAIL.n57 VTAIL.n20 6.59444
R846 VTAIL.n148 VTAIL.n114 6.59444
R847 VTAIL.n151 VTAIL.n114 6.59444
R848 VTAIL.n244 VTAIL.n210 6.59444
R849 VTAIL.n247 VTAIL.n210 6.59444
R850 VTAIL.n628 VTAIL.n591 6.59444
R851 VTAIL.n625 VTAIL.n591 6.59444
R852 VTAIL.n532 VTAIL.n495 6.59444
R853 VTAIL.n529 VTAIL.n495 6.59444
R854 VTAIL.n438 VTAIL.n401 6.59444
R855 VTAIL.n435 VTAIL.n401 6.59444
R856 VTAIL.n342 VTAIL.n305 6.59444
R857 VTAIL.n339 VTAIL.n305 6.59444
R858 VTAIL.n717 VTAIL.n686 5.81868
R859 VTAIL.n722 VTAIL.n682 5.81868
R860 VTAIL.n53 VTAIL.n22 5.81868
R861 VTAIL.n58 VTAIL.n18 5.81868
R862 VTAIL.n147 VTAIL.n116 5.81868
R863 VTAIL.n152 VTAIL.n112 5.81868
R864 VTAIL.n243 VTAIL.n212 5.81868
R865 VTAIL.n248 VTAIL.n208 5.81868
R866 VTAIL.n629 VTAIL.n589 5.81868
R867 VTAIL.n624 VTAIL.n593 5.81868
R868 VTAIL.n533 VTAIL.n493 5.81868
R869 VTAIL.n528 VTAIL.n497 5.81868
R870 VTAIL.n439 VTAIL.n399 5.81868
R871 VTAIL.n434 VTAIL.n403 5.81868
R872 VTAIL.n343 VTAIL.n303 5.81868
R873 VTAIL.n338 VTAIL.n307 5.81868
R874 VTAIL.n714 VTAIL.n713 5.04292
R875 VTAIL.n726 VTAIL.n725 5.04292
R876 VTAIL.n50 VTAIL.n49 5.04292
R877 VTAIL.n62 VTAIL.n61 5.04292
R878 VTAIL.n144 VTAIL.n143 5.04292
R879 VTAIL.n156 VTAIL.n155 5.04292
R880 VTAIL.n240 VTAIL.n239 5.04292
R881 VTAIL.n252 VTAIL.n251 5.04292
R882 VTAIL.n633 VTAIL.n632 5.04292
R883 VTAIL.n621 VTAIL.n620 5.04292
R884 VTAIL.n537 VTAIL.n536 5.04292
R885 VTAIL.n525 VTAIL.n524 5.04292
R886 VTAIL.n443 VTAIL.n442 5.04292
R887 VTAIL.n431 VTAIL.n430 5.04292
R888 VTAIL.n347 VTAIL.n346 5.04292
R889 VTAIL.n335 VTAIL.n334 5.04292
R890 VTAIL.n710 VTAIL.n688 4.26717
R891 VTAIL.n729 VTAIL.n680 4.26717
R892 VTAIL.n758 VTAIL.n666 4.26717
R893 VTAIL.n46 VTAIL.n24 4.26717
R894 VTAIL.n65 VTAIL.n16 4.26717
R895 VTAIL.n94 VTAIL.n2 4.26717
R896 VTAIL.n140 VTAIL.n118 4.26717
R897 VTAIL.n159 VTAIL.n110 4.26717
R898 VTAIL.n188 VTAIL.n96 4.26717
R899 VTAIL.n236 VTAIL.n214 4.26717
R900 VTAIL.n255 VTAIL.n206 4.26717
R901 VTAIL.n284 VTAIL.n192 4.26717
R902 VTAIL.n664 VTAIL.n572 4.26717
R903 VTAIL.n636 VTAIL.n587 4.26717
R904 VTAIL.n617 VTAIL.n595 4.26717
R905 VTAIL.n568 VTAIL.n476 4.26717
R906 VTAIL.n540 VTAIL.n491 4.26717
R907 VTAIL.n521 VTAIL.n499 4.26717
R908 VTAIL.n474 VTAIL.n382 4.26717
R909 VTAIL.n446 VTAIL.n397 4.26717
R910 VTAIL.n427 VTAIL.n405 4.26717
R911 VTAIL.n378 VTAIL.n286 4.26717
R912 VTAIL.n350 VTAIL.n301 4.26717
R913 VTAIL.n331 VTAIL.n309 4.26717
R914 VTAIL.n699 VTAIL.n695 3.70982
R915 VTAIL.n35 VTAIL.n31 3.70982
R916 VTAIL.n129 VTAIL.n125 3.70982
R917 VTAIL.n225 VTAIL.n221 3.70982
R918 VTAIL.n606 VTAIL.n602 3.70982
R919 VTAIL.n510 VTAIL.n506 3.70982
R920 VTAIL.n416 VTAIL.n412 3.70982
R921 VTAIL.n320 VTAIL.n316 3.70982
R922 VTAIL.n709 VTAIL.n690 3.49141
R923 VTAIL.n730 VTAIL.n678 3.49141
R924 VTAIL.n756 VTAIL.n755 3.49141
R925 VTAIL.n45 VTAIL.n26 3.49141
R926 VTAIL.n66 VTAIL.n14 3.49141
R927 VTAIL.n92 VTAIL.n91 3.49141
R928 VTAIL.n139 VTAIL.n120 3.49141
R929 VTAIL.n160 VTAIL.n108 3.49141
R930 VTAIL.n186 VTAIL.n185 3.49141
R931 VTAIL.n235 VTAIL.n216 3.49141
R932 VTAIL.n256 VTAIL.n204 3.49141
R933 VTAIL.n282 VTAIL.n281 3.49141
R934 VTAIL.n662 VTAIL.n661 3.49141
R935 VTAIL.n637 VTAIL.n585 3.49141
R936 VTAIL.n616 VTAIL.n597 3.49141
R937 VTAIL.n566 VTAIL.n565 3.49141
R938 VTAIL.n541 VTAIL.n489 3.49141
R939 VTAIL.n520 VTAIL.n501 3.49141
R940 VTAIL.n472 VTAIL.n471 3.49141
R941 VTAIL.n447 VTAIL.n395 3.49141
R942 VTAIL.n426 VTAIL.n407 3.49141
R943 VTAIL.n376 VTAIL.n375 3.49141
R944 VTAIL.n351 VTAIL.n299 3.49141
R945 VTAIL.n330 VTAIL.n311 3.49141
R946 VTAIL.n706 VTAIL.n705 2.71565
R947 VTAIL.n734 VTAIL.n733 2.71565
R948 VTAIL.n752 VTAIL.n668 2.71565
R949 VTAIL.n42 VTAIL.n41 2.71565
R950 VTAIL.n70 VTAIL.n69 2.71565
R951 VTAIL.n88 VTAIL.n4 2.71565
R952 VTAIL.n136 VTAIL.n135 2.71565
R953 VTAIL.n164 VTAIL.n163 2.71565
R954 VTAIL.n182 VTAIL.n98 2.71565
R955 VTAIL.n232 VTAIL.n231 2.71565
R956 VTAIL.n260 VTAIL.n259 2.71565
R957 VTAIL.n278 VTAIL.n194 2.71565
R958 VTAIL.n658 VTAIL.n574 2.71565
R959 VTAIL.n641 VTAIL.n640 2.71565
R960 VTAIL.n613 VTAIL.n612 2.71565
R961 VTAIL.n562 VTAIL.n478 2.71565
R962 VTAIL.n545 VTAIL.n544 2.71565
R963 VTAIL.n517 VTAIL.n516 2.71565
R964 VTAIL.n468 VTAIL.n384 2.71565
R965 VTAIL.n451 VTAIL.n450 2.71565
R966 VTAIL.n423 VTAIL.n422 2.71565
R967 VTAIL.n372 VTAIL.n288 2.71565
R968 VTAIL.n355 VTAIL.n354 2.71565
R969 VTAIL.n327 VTAIL.n326 2.71565
R970 VTAIL.n0 VTAIL.t11 1.94226
R971 VTAIL.n0 VTAIL.t10 1.94226
R972 VTAIL.n190 VTAIL.t2 1.94226
R973 VTAIL.n190 VTAIL.t4 1.94226
R974 VTAIL.n570 VTAIL.t0 1.94226
R975 VTAIL.n570 VTAIL.t3 1.94226
R976 VTAIL.n380 VTAIL.t12 1.94226
R977 VTAIL.n380 VTAIL.t9 1.94226
R978 VTAIL.n702 VTAIL.n692 1.93989
R979 VTAIL.n738 VTAIL.n676 1.93989
R980 VTAIL.n751 VTAIL.n670 1.93989
R981 VTAIL.n38 VTAIL.n28 1.93989
R982 VTAIL.n74 VTAIL.n12 1.93989
R983 VTAIL.n87 VTAIL.n6 1.93989
R984 VTAIL.n132 VTAIL.n122 1.93989
R985 VTAIL.n168 VTAIL.n106 1.93989
R986 VTAIL.n181 VTAIL.n100 1.93989
R987 VTAIL.n228 VTAIL.n218 1.93989
R988 VTAIL.n264 VTAIL.n202 1.93989
R989 VTAIL.n277 VTAIL.n196 1.93989
R990 VTAIL.n657 VTAIL.n576 1.93989
R991 VTAIL.n644 VTAIL.n582 1.93989
R992 VTAIL.n609 VTAIL.n599 1.93989
R993 VTAIL.n561 VTAIL.n480 1.93989
R994 VTAIL.n548 VTAIL.n486 1.93989
R995 VTAIL.n513 VTAIL.n503 1.93989
R996 VTAIL.n467 VTAIL.n386 1.93989
R997 VTAIL.n454 VTAIL.n392 1.93989
R998 VTAIL.n419 VTAIL.n409 1.93989
R999 VTAIL.n371 VTAIL.n290 1.93989
R1000 VTAIL.n358 VTAIL.n296 1.93989
R1001 VTAIL.n323 VTAIL.n313 1.93989
R1002 VTAIL.n381 VTAIL.n379 1.47464
R1003 VTAIL.n475 VTAIL.n381 1.47464
R1004 VTAIL.n571 VTAIL.n569 1.47464
R1005 VTAIL.n665 VTAIL.n571 1.47464
R1006 VTAIL.n285 VTAIL.n191 1.47464
R1007 VTAIL.n191 VTAIL.n189 1.47464
R1008 VTAIL.n95 VTAIL.n1 1.47464
R1009 VTAIL VTAIL.n759 1.41645
R1010 VTAIL.n701 VTAIL.n694 1.16414
R1011 VTAIL.n739 VTAIL.n674 1.16414
R1012 VTAIL.n748 VTAIL.n747 1.16414
R1013 VTAIL.n37 VTAIL.n30 1.16414
R1014 VTAIL.n75 VTAIL.n10 1.16414
R1015 VTAIL.n84 VTAIL.n83 1.16414
R1016 VTAIL.n131 VTAIL.n124 1.16414
R1017 VTAIL.n169 VTAIL.n104 1.16414
R1018 VTAIL.n178 VTAIL.n177 1.16414
R1019 VTAIL.n227 VTAIL.n220 1.16414
R1020 VTAIL.n265 VTAIL.n200 1.16414
R1021 VTAIL.n274 VTAIL.n273 1.16414
R1022 VTAIL.n654 VTAIL.n653 1.16414
R1023 VTAIL.n645 VTAIL.n580 1.16414
R1024 VTAIL.n608 VTAIL.n601 1.16414
R1025 VTAIL.n558 VTAIL.n557 1.16414
R1026 VTAIL.n549 VTAIL.n484 1.16414
R1027 VTAIL.n512 VTAIL.n505 1.16414
R1028 VTAIL.n464 VTAIL.n463 1.16414
R1029 VTAIL.n455 VTAIL.n390 1.16414
R1030 VTAIL.n418 VTAIL.n411 1.16414
R1031 VTAIL.n368 VTAIL.n367 1.16414
R1032 VTAIL.n359 VTAIL.n294 1.16414
R1033 VTAIL.n322 VTAIL.n315 1.16414
R1034 VTAIL.n569 VTAIL.n475 0.470328
R1035 VTAIL.n189 VTAIL.n95 0.470328
R1036 VTAIL.n698 VTAIL.n697 0.388379
R1037 VTAIL.n743 VTAIL.n742 0.388379
R1038 VTAIL.n744 VTAIL.n672 0.388379
R1039 VTAIL.n34 VTAIL.n33 0.388379
R1040 VTAIL.n79 VTAIL.n78 0.388379
R1041 VTAIL.n80 VTAIL.n8 0.388379
R1042 VTAIL.n128 VTAIL.n127 0.388379
R1043 VTAIL.n173 VTAIL.n172 0.388379
R1044 VTAIL.n174 VTAIL.n102 0.388379
R1045 VTAIL.n224 VTAIL.n223 0.388379
R1046 VTAIL.n269 VTAIL.n268 0.388379
R1047 VTAIL.n270 VTAIL.n198 0.388379
R1048 VTAIL.n650 VTAIL.n578 0.388379
R1049 VTAIL.n649 VTAIL.n648 0.388379
R1050 VTAIL.n605 VTAIL.n604 0.388379
R1051 VTAIL.n554 VTAIL.n482 0.388379
R1052 VTAIL.n553 VTAIL.n552 0.388379
R1053 VTAIL.n509 VTAIL.n508 0.388379
R1054 VTAIL.n460 VTAIL.n388 0.388379
R1055 VTAIL.n459 VTAIL.n458 0.388379
R1056 VTAIL.n415 VTAIL.n414 0.388379
R1057 VTAIL.n364 VTAIL.n292 0.388379
R1058 VTAIL.n363 VTAIL.n362 0.388379
R1059 VTAIL.n319 VTAIL.n318 0.388379
R1060 VTAIL.n700 VTAIL.n699 0.155672
R1061 VTAIL.n700 VTAIL.n691 0.155672
R1062 VTAIL.n707 VTAIL.n691 0.155672
R1063 VTAIL.n708 VTAIL.n707 0.155672
R1064 VTAIL.n708 VTAIL.n687 0.155672
R1065 VTAIL.n715 VTAIL.n687 0.155672
R1066 VTAIL.n716 VTAIL.n715 0.155672
R1067 VTAIL.n716 VTAIL.n683 0.155672
R1068 VTAIL.n723 VTAIL.n683 0.155672
R1069 VTAIL.n724 VTAIL.n723 0.155672
R1070 VTAIL.n724 VTAIL.n679 0.155672
R1071 VTAIL.n731 VTAIL.n679 0.155672
R1072 VTAIL.n732 VTAIL.n731 0.155672
R1073 VTAIL.n732 VTAIL.n675 0.155672
R1074 VTAIL.n740 VTAIL.n675 0.155672
R1075 VTAIL.n741 VTAIL.n740 0.155672
R1076 VTAIL.n741 VTAIL.n671 0.155672
R1077 VTAIL.n749 VTAIL.n671 0.155672
R1078 VTAIL.n750 VTAIL.n749 0.155672
R1079 VTAIL.n750 VTAIL.n667 0.155672
R1080 VTAIL.n757 VTAIL.n667 0.155672
R1081 VTAIL.n36 VTAIL.n35 0.155672
R1082 VTAIL.n36 VTAIL.n27 0.155672
R1083 VTAIL.n43 VTAIL.n27 0.155672
R1084 VTAIL.n44 VTAIL.n43 0.155672
R1085 VTAIL.n44 VTAIL.n23 0.155672
R1086 VTAIL.n51 VTAIL.n23 0.155672
R1087 VTAIL.n52 VTAIL.n51 0.155672
R1088 VTAIL.n52 VTAIL.n19 0.155672
R1089 VTAIL.n59 VTAIL.n19 0.155672
R1090 VTAIL.n60 VTAIL.n59 0.155672
R1091 VTAIL.n60 VTAIL.n15 0.155672
R1092 VTAIL.n67 VTAIL.n15 0.155672
R1093 VTAIL.n68 VTAIL.n67 0.155672
R1094 VTAIL.n68 VTAIL.n11 0.155672
R1095 VTAIL.n76 VTAIL.n11 0.155672
R1096 VTAIL.n77 VTAIL.n76 0.155672
R1097 VTAIL.n77 VTAIL.n7 0.155672
R1098 VTAIL.n85 VTAIL.n7 0.155672
R1099 VTAIL.n86 VTAIL.n85 0.155672
R1100 VTAIL.n86 VTAIL.n3 0.155672
R1101 VTAIL.n93 VTAIL.n3 0.155672
R1102 VTAIL.n130 VTAIL.n129 0.155672
R1103 VTAIL.n130 VTAIL.n121 0.155672
R1104 VTAIL.n137 VTAIL.n121 0.155672
R1105 VTAIL.n138 VTAIL.n137 0.155672
R1106 VTAIL.n138 VTAIL.n117 0.155672
R1107 VTAIL.n145 VTAIL.n117 0.155672
R1108 VTAIL.n146 VTAIL.n145 0.155672
R1109 VTAIL.n146 VTAIL.n113 0.155672
R1110 VTAIL.n153 VTAIL.n113 0.155672
R1111 VTAIL.n154 VTAIL.n153 0.155672
R1112 VTAIL.n154 VTAIL.n109 0.155672
R1113 VTAIL.n161 VTAIL.n109 0.155672
R1114 VTAIL.n162 VTAIL.n161 0.155672
R1115 VTAIL.n162 VTAIL.n105 0.155672
R1116 VTAIL.n170 VTAIL.n105 0.155672
R1117 VTAIL.n171 VTAIL.n170 0.155672
R1118 VTAIL.n171 VTAIL.n101 0.155672
R1119 VTAIL.n179 VTAIL.n101 0.155672
R1120 VTAIL.n180 VTAIL.n179 0.155672
R1121 VTAIL.n180 VTAIL.n97 0.155672
R1122 VTAIL.n187 VTAIL.n97 0.155672
R1123 VTAIL.n226 VTAIL.n225 0.155672
R1124 VTAIL.n226 VTAIL.n217 0.155672
R1125 VTAIL.n233 VTAIL.n217 0.155672
R1126 VTAIL.n234 VTAIL.n233 0.155672
R1127 VTAIL.n234 VTAIL.n213 0.155672
R1128 VTAIL.n241 VTAIL.n213 0.155672
R1129 VTAIL.n242 VTAIL.n241 0.155672
R1130 VTAIL.n242 VTAIL.n209 0.155672
R1131 VTAIL.n249 VTAIL.n209 0.155672
R1132 VTAIL.n250 VTAIL.n249 0.155672
R1133 VTAIL.n250 VTAIL.n205 0.155672
R1134 VTAIL.n257 VTAIL.n205 0.155672
R1135 VTAIL.n258 VTAIL.n257 0.155672
R1136 VTAIL.n258 VTAIL.n201 0.155672
R1137 VTAIL.n266 VTAIL.n201 0.155672
R1138 VTAIL.n267 VTAIL.n266 0.155672
R1139 VTAIL.n267 VTAIL.n197 0.155672
R1140 VTAIL.n275 VTAIL.n197 0.155672
R1141 VTAIL.n276 VTAIL.n275 0.155672
R1142 VTAIL.n276 VTAIL.n193 0.155672
R1143 VTAIL.n283 VTAIL.n193 0.155672
R1144 VTAIL.n663 VTAIL.n573 0.155672
R1145 VTAIL.n656 VTAIL.n573 0.155672
R1146 VTAIL.n656 VTAIL.n655 0.155672
R1147 VTAIL.n655 VTAIL.n577 0.155672
R1148 VTAIL.n647 VTAIL.n577 0.155672
R1149 VTAIL.n647 VTAIL.n646 0.155672
R1150 VTAIL.n646 VTAIL.n581 0.155672
R1151 VTAIL.n639 VTAIL.n581 0.155672
R1152 VTAIL.n639 VTAIL.n638 0.155672
R1153 VTAIL.n638 VTAIL.n586 0.155672
R1154 VTAIL.n631 VTAIL.n586 0.155672
R1155 VTAIL.n631 VTAIL.n630 0.155672
R1156 VTAIL.n630 VTAIL.n590 0.155672
R1157 VTAIL.n623 VTAIL.n590 0.155672
R1158 VTAIL.n623 VTAIL.n622 0.155672
R1159 VTAIL.n622 VTAIL.n594 0.155672
R1160 VTAIL.n615 VTAIL.n594 0.155672
R1161 VTAIL.n615 VTAIL.n614 0.155672
R1162 VTAIL.n614 VTAIL.n598 0.155672
R1163 VTAIL.n607 VTAIL.n598 0.155672
R1164 VTAIL.n607 VTAIL.n606 0.155672
R1165 VTAIL.n567 VTAIL.n477 0.155672
R1166 VTAIL.n560 VTAIL.n477 0.155672
R1167 VTAIL.n560 VTAIL.n559 0.155672
R1168 VTAIL.n559 VTAIL.n481 0.155672
R1169 VTAIL.n551 VTAIL.n481 0.155672
R1170 VTAIL.n551 VTAIL.n550 0.155672
R1171 VTAIL.n550 VTAIL.n485 0.155672
R1172 VTAIL.n543 VTAIL.n485 0.155672
R1173 VTAIL.n543 VTAIL.n542 0.155672
R1174 VTAIL.n542 VTAIL.n490 0.155672
R1175 VTAIL.n535 VTAIL.n490 0.155672
R1176 VTAIL.n535 VTAIL.n534 0.155672
R1177 VTAIL.n534 VTAIL.n494 0.155672
R1178 VTAIL.n527 VTAIL.n494 0.155672
R1179 VTAIL.n527 VTAIL.n526 0.155672
R1180 VTAIL.n526 VTAIL.n498 0.155672
R1181 VTAIL.n519 VTAIL.n498 0.155672
R1182 VTAIL.n519 VTAIL.n518 0.155672
R1183 VTAIL.n518 VTAIL.n502 0.155672
R1184 VTAIL.n511 VTAIL.n502 0.155672
R1185 VTAIL.n511 VTAIL.n510 0.155672
R1186 VTAIL.n473 VTAIL.n383 0.155672
R1187 VTAIL.n466 VTAIL.n383 0.155672
R1188 VTAIL.n466 VTAIL.n465 0.155672
R1189 VTAIL.n465 VTAIL.n387 0.155672
R1190 VTAIL.n457 VTAIL.n387 0.155672
R1191 VTAIL.n457 VTAIL.n456 0.155672
R1192 VTAIL.n456 VTAIL.n391 0.155672
R1193 VTAIL.n449 VTAIL.n391 0.155672
R1194 VTAIL.n449 VTAIL.n448 0.155672
R1195 VTAIL.n448 VTAIL.n396 0.155672
R1196 VTAIL.n441 VTAIL.n396 0.155672
R1197 VTAIL.n441 VTAIL.n440 0.155672
R1198 VTAIL.n440 VTAIL.n400 0.155672
R1199 VTAIL.n433 VTAIL.n400 0.155672
R1200 VTAIL.n433 VTAIL.n432 0.155672
R1201 VTAIL.n432 VTAIL.n404 0.155672
R1202 VTAIL.n425 VTAIL.n404 0.155672
R1203 VTAIL.n425 VTAIL.n424 0.155672
R1204 VTAIL.n424 VTAIL.n408 0.155672
R1205 VTAIL.n417 VTAIL.n408 0.155672
R1206 VTAIL.n417 VTAIL.n416 0.155672
R1207 VTAIL.n377 VTAIL.n287 0.155672
R1208 VTAIL.n370 VTAIL.n287 0.155672
R1209 VTAIL.n370 VTAIL.n369 0.155672
R1210 VTAIL.n369 VTAIL.n291 0.155672
R1211 VTAIL.n361 VTAIL.n291 0.155672
R1212 VTAIL.n361 VTAIL.n360 0.155672
R1213 VTAIL.n360 VTAIL.n295 0.155672
R1214 VTAIL.n353 VTAIL.n295 0.155672
R1215 VTAIL.n353 VTAIL.n352 0.155672
R1216 VTAIL.n352 VTAIL.n300 0.155672
R1217 VTAIL.n345 VTAIL.n300 0.155672
R1218 VTAIL.n345 VTAIL.n344 0.155672
R1219 VTAIL.n344 VTAIL.n304 0.155672
R1220 VTAIL.n337 VTAIL.n304 0.155672
R1221 VTAIL.n337 VTAIL.n336 0.155672
R1222 VTAIL.n336 VTAIL.n308 0.155672
R1223 VTAIL.n329 VTAIL.n308 0.155672
R1224 VTAIL.n329 VTAIL.n328 0.155672
R1225 VTAIL.n328 VTAIL.n312 0.155672
R1226 VTAIL.n321 VTAIL.n312 0.155672
R1227 VTAIL.n321 VTAIL.n320 0.155672
R1228 VTAIL VTAIL.n1 0.0586897
R1229 VP.n11 VP.t3 323.56
R1230 VP.n5 VP.t0 292.344
R1231 VP.n29 VP.t1 292.344
R1232 VP.n36 VP.t5 292.344
R1233 VP.n43 VP.t4 292.344
R1234 VP.n23 VP.t6 292.344
R1235 VP.n16 VP.t2 292.344
R1236 VP.n10 VP.t7 292.344
R1237 VP.n25 VP.n5 170.399
R1238 VP.n44 VP.n43 170.399
R1239 VP.n24 VP.n23 170.399
R1240 VP.n12 VP.n9 161.3
R1241 VP.n14 VP.n13 161.3
R1242 VP.n15 VP.n8 161.3
R1243 VP.n18 VP.n17 161.3
R1244 VP.n19 VP.n7 161.3
R1245 VP.n21 VP.n20 161.3
R1246 VP.n22 VP.n6 161.3
R1247 VP.n42 VP.n0 161.3
R1248 VP.n41 VP.n40 161.3
R1249 VP.n39 VP.n1 161.3
R1250 VP.n38 VP.n37 161.3
R1251 VP.n35 VP.n2 161.3
R1252 VP.n34 VP.n33 161.3
R1253 VP.n32 VP.n3 161.3
R1254 VP.n31 VP.n30 161.3
R1255 VP.n28 VP.n4 161.3
R1256 VP.n27 VP.n26 161.3
R1257 VP.n11 VP.n10 59.9731
R1258 VP.n35 VP.n34 56.5617
R1259 VP.n15 VP.n14 56.5617
R1260 VP.n25 VP.n24 48.7581
R1261 VP.n30 VP.n28 44.4521
R1262 VP.n41 VP.n1 44.4521
R1263 VP.n21 VP.n7 44.4521
R1264 VP.n28 VP.n27 36.702
R1265 VP.n42 VP.n41 36.702
R1266 VP.n22 VP.n21 36.702
R1267 VP.n12 VP.n11 26.618
R1268 VP.n34 VP.n3 24.5923
R1269 VP.n37 VP.n35 24.5923
R1270 VP.n17 VP.n15 24.5923
R1271 VP.n14 VP.n9 24.5923
R1272 VP.n30 VP.n29 19.4281
R1273 VP.n36 VP.n1 19.4281
R1274 VP.n16 VP.n7 19.4281
R1275 VP.n27 VP.n5 15.4934
R1276 VP.n43 VP.n42 15.4934
R1277 VP.n23 VP.n22 15.4934
R1278 VP.n29 VP.n3 5.16479
R1279 VP.n37 VP.n36 5.16479
R1280 VP.n17 VP.n16 5.16479
R1281 VP.n10 VP.n9 5.16479
R1282 VP.n13 VP.n12 0.189894
R1283 VP.n13 VP.n8 0.189894
R1284 VP.n18 VP.n8 0.189894
R1285 VP.n19 VP.n18 0.189894
R1286 VP.n20 VP.n19 0.189894
R1287 VP.n20 VP.n6 0.189894
R1288 VP.n24 VP.n6 0.189894
R1289 VP.n26 VP.n25 0.189894
R1290 VP.n26 VP.n4 0.189894
R1291 VP.n31 VP.n4 0.189894
R1292 VP.n32 VP.n31 0.189894
R1293 VP.n33 VP.n32 0.189894
R1294 VP.n33 VP.n2 0.189894
R1295 VP.n38 VP.n2 0.189894
R1296 VP.n39 VP.n38 0.189894
R1297 VP.n40 VP.n39 0.189894
R1298 VP.n40 VP.n0 0.189894
R1299 VP.n44 VP.n0 0.189894
R1300 VP VP.n44 0.0516364
R1301 VDD1 VDD1.n0 69.0237
R1302 VDD1.n3 VDD1.n2 68.9099
R1303 VDD1.n3 VDD1.n1 68.9099
R1304 VDD1.n5 VDD1.n4 68.2282
R1305 VDD1.n5 VDD1.n3 45.363
R1306 VDD1.n4 VDD1.t5 1.94226
R1307 VDD1.n4 VDD1.t1 1.94226
R1308 VDD1.n0 VDD1.t4 1.94226
R1309 VDD1.n0 VDD1.t0 1.94226
R1310 VDD1.n2 VDD1.t2 1.94226
R1311 VDD1.n2 VDD1.t3 1.94226
R1312 VDD1.n1 VDD1.t7 1.94226
R1313 VDD1.n1 VDD1.t6 1.94226
R1314 VDD1 VDD1.n5 0.679379
R1315 B.n531 B.n530 585
R1316 B.n532 B.n83 585
R1317 B.n534 B.n533 585
R1318 B.n535 B.n82 585
R1319 B.n537 B.n536 585
R1320 B.n538 B.n81 585
R1321 B.n540 B.n539 585
R1322 B.n541 B.n80 585
R1323 B.n543 B.n542 585
R1324 B.n544 B.n79 585
R1325 B.n546 B.n545 585
R1326 B.n547 B.n78 585
R1327 B.n549 B.n548 585
R1328 B.n550 B.n77 585
R1329 B.n552 B.n551 585
R1330 B.n553 B.n76 585
R1331 B.n555 B.n554 585
R1332 B.n556 B.n75 585
R1333 B.n558 B.n557 585
R1334 B.n559 B.n74 585
R1335 B.n561 B.n560 585
R1336 B.n562 B.n73 585
R1337 B.n564 B.n563 585
R1338 B.n565 B.n72 585
R1339 B.n567 B.n566 585
R1340 B.n568 B.n71 585
R1341 B.n570 B.n569 585
R1342 B.n571 B.n70 585
R1343 B.n573 B.n572 585
R1344 B.n574 B.n69 585
R1345 B.n576 B.n575 585
R1346 B.n577 B.n68 585
R1347 B.n579 B.n578 585
R1348 B.n580 B.n67 585
R1349 B.n582 B.n581 585
R1350 B.n583 B.n66 585
R1351 B.n585 B.n584 585
R1352 B.n586 B.n65 585
R1353 B.n588 B.n587 585
R1354 B.n589 B.n64 585
R1355 B.n591 B.n590 585
R1356 B.n592 B.n63 585
R1357 B.n594 B.n593 585
R1358 B.n595 B.n62 585
R1359 B.n597 B.n596 585
R1360 B.n598 B.n61 585
R1361 B.n600 B.n599 585
R1362 B.n601 B.n60 585
R1363 B.n603 B.n602 585
R1364 B.n604 B.n59 585
R1365 B.n606 B.n605 585
R1366 B.n607 B.n58 585
R1367 B.n609 B.n608 585
R1368 B.n610 B.n57 585
R1369 B.n612 B.n611 585
R1370 B.n613 B.n54 585
R1371 B.n616 B.n615 585
R1372 B.n617 B.n53 585
R1373 B.n619 B.n618 585
R1374 B.n620 B.n52 585
R1375 B.n622 B.n621 585
R1376 B.n623 B.n51 585
R1377 B.n625 B.n624 585
R1378 B.n626 B.n47 585
R1379 B.n628 B.n627 585
R1380 B.n629 B.n46 585
R1381 B.n631 B.n630 585
R1382 B.n632 B.n45 585
R1383 B.n634 B.n633 585
R1384 B.n635 B.n44 585
R1385 B.n637 B.n636 585
R1386 B.n638 B.n43 585
R1387 B.n640 B.n639 585
R1388 B.n641 B.n42 585
R1389 B.n643 B.n642 585
R1390 B.n644 B.n41 585
R1391 B.n646 B.n645 585
R1392 B.n647 B.n40 585
R1393 B.n649 B.n648 585
R1394 B.n650 B.n39 585
R1395 B.n652 B.n651 585
R1396 B.n653 B.n38 585
R1397 B.n655 B.n654 585
R1398 B.n656 B.n37 585
R1399 B.n658 B.n657 585
R1400 B.n659 B.n36 585
R1401 B.n661 B.n660 585
R1402 B.n662 B.n35 585
R1403 B.n664 B.n663 585
R1404 B.n665 B.n34 585
R1405 B.n667 B.n666 585
R1406 B.n668 B.n33 585
R1407 B.n670 B.n669 585
R1408 B.n671 B.n32 585
R1409 B.n673 B.n672 585
R1410 B.n674 B.n31 585
R1411 B.n676 B.n675 585
R1412 B.n677 B.n30 585
R1413 B.n679 B.n678 585
R1414 B.n680 B.n29 585
R1415 B.n682 B.n681 585
R1416 B.n683 B.n28 585
R1417 B.n685 B.n684 585
R1418 B.n686 B.n27 585
R1419 B.n688 B.n687 585
R1420 B.n689 B.n26 585
R1421 B.n691 B.n690 585
R1422 B.n692 B.n25 585
R1423 B.n694 B.n693 585
R1424 B.n695 B.n24 585
R1425 B.n697 B.n696 585
R1426 B.n698 B.n23 585
R1427 B.n700 B.n699 585
R1428 B.n701 B.n22 585
R1429 B.n703 B.n702 585
R1430 B.n704 B.n21 585
R1431 B.n706 B.n705 585
R1432 B.n707 B.n20 585
R1433 B.n709 B.n708 585
R1434 B.n710 B.n19 585
R1435 B.n712 B.n711 585
R1436 B.n529 B.n84 585
R1437 B.n528 B.n527 585
R1438 B.n526 B.n85 585
R1439 B.n525 B.n524 585
R1440 B.n523 B.n86 585
R1441 B.n522 B.n521 585
R1442 B.n520 B.n87 585
R1443 B.n519 B.n518 585
R1444 B.n517 B.n88 585
R1445 B.n516 B.n515 585
R1446 B.n514 B.n89 585
R1447 B.n513 B.n512 585
R1448 B.n511 B.n90 585
R1449 B.n510 B.n509 585
R1450 B.n508 B.n91 585
R1451 B.n507 B.n506 585
R1452 B.n505 B.n92 585
R1453 B.n504 B.n503 585
R1454 B.n502 B.n93 585
R1455 B.n501 B.n500 585
R1456 B.n499 B.n94 585
R1457 B.n498 B.n497 585
R1458 B.n496 B.n95 585
R1459 B.n495 B.n494 585
R1460 B.n493 B.n96 585
R1461 B.n492 B.n491 585
R1462 B.n490 B.n97 585
R1463 B.n489 B.n488 585
R1464 B.n487 B.n98 585
R1465 B.n486 B.n485 585
R1466 B.n484 B.n99 585
R1467 B.n483 B.n482 585
R1468 B.n481 B.n100 585
R1469 B.n480 B.n479 585
R1470 B.n478 B.n101 585
R1471 B.n477 B.n476 585
R1472 B.n475 B.n102 585
R1473 B.n474 B.n473 585
R1474 B.n472 B.n103 585
R1475 B.n471 B.n470 585
R1476 B.n469 B.n104 585
R1477 B.n468 B.n467 585
R1478 B.n466 B.n105 585
R1479 B.n465 B.n464 585
R1480 B.n463 B.n106 585
R1481 B.n462 B.n461 585
R1482 B.n460 B.n107 585
R1483 B.n459 B.n458 585
R1484 B.n457 B.n108 585
R1485 B.n456 B.n455 585
R1486 B.n454 B.n109 585
R1487 B.n453 B.n452 585
R1488 B.n451 B.n110 585
R1489 B.n450 B.n449 585
R1490 B.n448 B.n111 585
R1491 B.n447 B.n446 585
R1492 B.n445 B.n112 585
R1493 B.n444 B.n443 585
R1494 B.n442 B.n113 585
R1495 B.n441 B.n440 585
R1496 B.n439 B.n114 585
R1497 B.n438 B.n437 585
R1498 B.n436 B.n115 585
R1499 B.n435 B.n434 585
R1500 B.n433 B.n116 585
R1501 B.n432 B.n431 585
R1502 B.n430 B.n117 585
R1503 B.n245 B.n244 585
R1504 B.n246 B.n179 585
R1505 B.n248 B.n247 585
R1506 B.n249 B.n178 585
R1507 B.n251 B.n250 585
R1508 B.n252 B.n177 585
R1509 B.n254 B.n253 585
R1510 B.n255 B.n176 585
R1511 B.n257 B.n256 585
R1512 B.n258 B.n175 585
R1513 B.n260 B.n259 585
R1514 B.n261 B.n174 585
R1515 B.n263 B.n262 585
R1516 B.n264 B.n173 585
R1517 B.n266 B.n265 585
R1518 B.n267 B.n172 585
R1519 B.n269 B.n268 585
R1520 B.n270 B.n171 585
R1521 B.n272 B.n271 585
R1522 B.n273 B.n170 585
R1523 B.n275 B.n274 585
R1524 B.n276 B.n169 585
R1525 B.n278 B.n277 585
R1526 B.n279 B.n168 585
R1527 B.n281 B.n280 585
R1528 B.n282 B.n167 585
R1529 B.n284 B.n283 585
R1530 B.n285 B.n166 585
R1531 B.n287 B.n286 585
R1532 B.n288 B.n165 585
R1533 B.n290 B.n289 585
R1534 B.n291 B.n164 585
R1535 B.n293 B.n292 585
R1536 B.n294 B.n163 585
R1537 B.n296 B.n295 585
R1538 B.n297 B.n162 585
R1539 B.n299 B.n298 585
R1540 B.n300 B.n161 585
R1541 B.n302 B.n301 585
R1542 B.n303 B.n160 585
R1543 B.n305 B.n304 585
R1544 B.n306 B.n159 585
R1545 B.n308 B.n307 585
R1546 B.n309 B.n158 585
R1547 B.n311 B.n310 585
R1548 B.n312 B.n157 585
R1549 B.n314 B.n313 585
R1550 B.n315 B.n156 585
R1551 B.n317 B.n316 585
R1552 B.n318 B.n155 585
R1553 B.n320 B.n319 585
R1554 B.n321 B.n154 585
R1555 B.n323 B.n322 585
R1556 B.n324 B.n153 585
R1557 B.n326 B.n325 585
R1558 B.n327 B.n150 585
R1559 B.n330 B.n329 585
R1560 B.n331 B.n149 585
R1561 B.n333 B.n332 585
R1562 B.n334 B.n148 585
R1563 B.n336 B.n335 585
R1564 B.n337 B.n147 585
R1565 B.n339 B.n338 585
R1566 B.n340 B.n146 585
R1567 B.n345 B.n344 585
R1568 B.n346 B.n145 585
R1569 B.n348 B.n347 585
R1570 B.n349 B.n144 585
R1571 B.n351 B.n350 585
R1572 B.n352 B.n143 585
R1573 B.n354 B.n353 585
R1574 B.n355 B.n142 585
R1575 B.n357 B.n356 585
R1576 B.n358 B.n141 585
R1577 B.n360 B.n359 585
R1578 B.n361 B.n140 585
R1579 B.n363 B.n362 585
R1580 B.n364 B.n139 585
R1581 B.n366 B.n365 585
R1582 B.n367 B.n138 585
R1583 B.n369 B.n368 585
R1584 B.n370 B.n137 585
R1585 B.n372 B.n371 585
R1586 B.n373 B.n136 585
R1587 B.n375 B.n374 585
R1588 B.n376 B.n135 585
R1589 B.n378 B.n377 585
R1590 B.n379 B.n134 585
R1591 B.n381 B.n380 585
R1592 B.n382 B.n133 585
R1593 B.n384 B.n383 585
R1594 B.n385 B.n132 585
R1595 B.n387 B.n386 585
R1596 B.n388 B.n131 585
R1597 B.n390 B.n389 585
R1598 B.n391 B.n130 585
R1599 B.n393 B.n392 585
R1600 B.n394 B.n129 585
R1601 B.n396 B.n395 585
R1602 B.n397 B.n128 585
R1603 B.n399 B.n398 585
R1604 B.n400 B.n127 585
R1605 B.n402 B.n401 585
R1606 B.n403 B.n126 585
R1607 B.n405 B.n404 585
R1608 B.n406 B.n125 585
R1609 B.n408 B.n407 585
R1610 B.n409 B.n124 585
R1611 B.n411 B.n410 585
R1612 B.n412 B.n123 585
R1613 B.n414 B.n413 585
R1614 B.n415 B.n122 585
R1615 B.n417 B.n416 585
R1616 B.n418 B.n121 585
R1617 B.n420 B.n419 585
R1618 B.n421 B.n120 585
R1619 B.n423 B.n422 585
R1620 B.n424 B.n119 585
R1621 B.n426 B.n425 585
R1622 B.n427 B.n118 585
R1623 B.n429 B.n428 585
R1624 B.n243 B.n180 585
R1625 B.n242 B.n241 585
R1626 B.n240 B.n181 585
R1627 B.n239 B.n238 585
R1628 B.n237 B.n182 585
R1629 B.n236 B.n235 585
R1630 B.n234 B.n183 585
R1631 B.n233 B.n232 585
R1632 B.n231 B.n184 585
R1633 B.n230 B.n229 585
R1634 B.n228 B.n185 585
R1635 B.n227 B.n226 585
R1636 B.n225 B.n186 585
R1637 B.n224 B.n223 585
R1638 B.n222 B.n187 585
R1639 B.n221 B.n220 585
R1640 B.n219 B.n188 585
R1641 B.n218 B.n217 585
R1642 B.n216 B.n189 585
R1643 B.n215 B.n214 585
R1644 B.n213 B.n190 585
R1645 B.n212 B.n211 585
R1646 B.n210 B.n191 585
R1647 B.n209 B.n208 585
R1648 B.n207 B.n192 585
R1649 B.n206 B.n205 585
R1650 B.n204 B.n193 585
R1651 B.n203 B.n202 585
R1652 B.n201 B.n194 585
R1653 B.n200 B.n199 585
R1654 B.n198 B.n195 585
R1655 B.n197 B.n196 585
R1656 B.n2 B.n0 585
R1657 B.n761 B.n1 585
R1658 B.n760 B.n759 585
R1659 B.n758 B.n3 585
R1660 B.n757 B.n756 585
R1661 B.n755 B.n4 585
R1662 B.n754 B.n753 585
R1663 B.n752 B.n5 585
R1664 B.n751 B.n750 585
R1665 B.n749 B.n6 585
R1666 B.n748 B.n747 585
R1667 B.n746 B.n7 585
R1668 B.n745 B.n744 585
R1669 B.n743 B.n8 585
R1670 B.n742 B.n741 585
R1671 B.n740 B.n9 585
R1672 B.n739 B.n738 585
R1673 B.n737 B.n10 585
R1674 B.n736 B.n735 585
R1675 B.n734 B.n11 585
R1676 B.n733 B.n732 585
R1677 B.n731 B.n12 585
R1678 B.n730 B.n729 585
R1679 B.n728 B.n13 585
R1680 B.n727 B.n726 585
R1681 B.n725 B.n14 585
R1682 B.n724 B.n723 585
R1683 B.n722 B.n15 585
R1684 B.n721 B.n720 585
R1685 B.n719 B.n16 585
R1686 B.n718 B.n717 585
R1687 B.n716 B.n17 585
R1688 B.n715 B.n714 585
R1689 B.n713 B.n18 585
R1690 B.n763 B.n762 585
R1691 B.n245 B.n180 516.524
R1692 B.n713 B.n712 516.524
R1693 B.n430 B.n429 516.524
R1694 B.n531 B.n84 516.524
R1695 B.n341 B.t3 497.307
R1696 B.n151 B.t6 497.307
R1697 B.n48 B.t0 497.307
R1698 B.n55 B.t9 497.307
R1699 B.n341 B.t5 494.041
R1700 B.n55 B.t10 494.041
R1701 B.n151 B.t8 494.041
R1702 B.n48 B.t1 494.041
R1703 B.n342 B.t4 460.877
R1704 B.n56 B.t11 460.877
R1705 B.n152 B.t7 460.877
R1706 B.n49 B.t2 460.877
R1707 B.n241 B.n180 163.367
R1708 B.n241 B.n240 163.367
R1709 B.n240 B.n239 163.367
R1710 B.n239 B.n182 163.367
R1711 B.n235 B.n182 163.367
R1712 B.n235 B.n234 163.367
R1713 B.n234 B.n233 163.367
R1714 B.n233 B.n184 163.367
R1715 B.n229 B.n184 163.367
R1716 B.n229 B.n228 163.367
R1717 B.n228 B.n227 163.367
R1718 B.n227 B.n186 163.367
R1719 B.n223 B.n186 163.367
R1720 B.n223 B.n222 163.367
R1721 B.n222 B.n221 163.367
R1722 B.n221 B.n188 163.367
R1723 B.n217 B.n188 163.367
R1724 B.n217 B.n216 163.367
R1725 B.n216 B.n215 163.367
R1726 B.n215 B.n190 163.367
R1727 B.n211 B.n190 163.367
R1728 B.n211 B.n210 163.367
R1729 B.n210 B.n209 163.367
R1730 B.n209 B.n192 163.367
R1731 B.n205 B.n192 163.367
R1732 B.n205 B.n204 163.367
R1733 B.n204 B.n203 163.367
R1734 B.n203 B.n194 163.367
R1735 B.n199 B.n194 163.367
R1736 B.n199 B.n198 163.367
R1737 B.n198 B.n197 163.367
R1738 B.n197 B.n2 163.367
R1739 B.n762 B.n2 163.367
R1740 B.n762 B.n761 163.367
R1741 B.n761 B.n760 163.367
R1742 B.n760 B.n3 163.367
R1743 B.n756 B.n3 163.367
R1744 B.n756 B.n755 163.367
R1745 B.n755 B.n754 163.367
R1746 B.n754 B.n5 163.367
R1747 B.n750 B.n5 163.367
R1748 B.n750 B.n749 163.367
R1749 B.n749 B.n748 163.367
R1750 B.n748 B.n7 163.367
R1751 B.n744 B.n7 163.367
R1752 B.n744 B.n743 163.367
R1753 B.n743 B.n742 163.367
R1754 B.n742 B.n9 163.367
R1755 B.n738 B.n9 163.367
R1756 B.n738 B.n737 163.367
R1757 B.n737 B.n736 163.367
R1758 B.n736 B.n11 163.367
R1759 B.n732 B.n11 163.367
R1760 B.n732 B.n731 163.367
R1761 B.n731 B.n730 163.367
R1762 B.n730 B.n13 163.367
R1763 B.n726 B.n13 163.367
R1764 B.n726 B.n725 163.367
R1765 B.n725 B.n724 163.367
R1766 B.n724 B.n15 163.367
R1767 B.n720 B.n15 163.367
R1768 B.n720 B.n719 163.367
R1769 B.n719 B.n718 163.367
R1770 B.n718 B.n17 163.367
R1771 B.n714 B.n17 163.367
R1772 B.n714 B.n713 163.367
R1773 B.n246 B.n245 163.367
R1774 B.n247 B.n246 163.367
R1775 B.n247 B.n178 163.367
R1776 B.n251 B.n178 163.367
R1777 B.n252 B.n251 163.367
R1778 B.n253 B.n252 163.367
R1779 B.n253 B.n176 163.367
R1780 B.n257 B.n176 163.367
R1781 B.n258 B.n257 163.367
R1782 B.n259 B.n258 163.367
R1783 B.n259 B.n174 163.367
R1784 B.n263 B.n174 163.367
R1785 B.n264 B.n263 163.367
R1786 B.n265 B.n264 163.367
R1787 B.n265 B.n172 163.367
R1788 B.n269 B.n172 163.367
R1789 B.n270 B.n269 163.367
R1790 B.n271 B.n270 163.367
R1791 B.n271 B.n170 163.367
R1792 B.n275 B.n170 163.367
R1793 B.n276 B.n275 163.367
R1794 B.n277 B.n276 163.367
R1795 B.n277 B.n168 163.367
R1796 B.n281 B.n168 163.367
R1797 B.n282 B.n281 163.367
R1798 B.n283 B.n282 163.367
R1799 B.n283 B.n166 163.367
R1800 B.n287 B.n166 163.367
R1801 B.n288 B.n287 163.367
R1802 B.n289 B.n288 163.367
R1803 B.n289 B.n164 163.367
R1804 B.n293 B.n164 163.367
R1805 B.n294 B.n293 163.367
R1806 B.n295 B.n294 163.367
R1807 B.n295 B.n162 163.367
R1808 B.n299 B.n162 163.367
R1809 B.n300 B.n299 163.367
R1810 B.n301 B.n300 163.367
R1811 B.n301 B.n160 163.367
R1812 B.n305 B.n160 163.367
R1813 B.n306 B.n305 163.367
R1814 B.n307 B.n306 163.367
R1815 B.n307 B.n158 163.367
R1816 B.n311 B.n158 163.367
R1817 B.n312 B.n311 163.367
R1818 B.n313 B.n312 163.367
R1819 B.n313 B.n156 163.367
R1820 B.n317 B.n156 163.367
R1821 B.n318 B.n317 163.367
R1822 B.n319 B.n318 163.367
R1823 B.n319 B.n154 163.367
R1824 B.n323 B.n154 163.367
R1825 B.n324 B.n323 163.367
R1826 B.n325 B.n324 163.367
R1827 B.n325 B.n150 163.367
R1828 B.n330 B.n150 163.367
R1829 B.n331 B.n330 163.367
R1830 B.n332 B.n331 163.367
R1831 B.n332 B.n148 163.367
R1832 B.n336 B.n148 163.367
R1833 B.n337 B.n336 163.367
R1834 B.n338 B.n337 163.367
R1835 B.n338 B.n146 163.367
R1836 B.n345 B.n146 163.367
R1837 B.n346 B.n345 163.367
R1838 B.n347 B.n346 163.367
R1839 B.n347 B.n144 163.367
R1840 B.n351 B.n144 163.367
R1841 B.n352 B.n351 163.367
R1842 B.n353 B.n352 163.367
R1843 B.n353 B.n142 163.367
R1844 B.n357 B.n142 163.367
R1845 B.n358 B.n357 163.367
R1846 B.n359 B.n358 163.367
R1847 B.n359 B.n140 163.367
R1848 B.n363 B.n140 163.367
R1849 B.n364 B.n363 163.367
R1850 B.n365 B.n364 163.367
R1851 B.n365 B.n138 163.367
R1852 B.n369 B.n138 163.367
R1853 B.n370 B.n369 163.367
R1854 B.n371 B.n370 163.367
R1855 B.n371 B.n136 163.367
R1856 B.n375 B.n136 163.367
R1857 B.n376 B.n375 163.367
R1858 B.n377 B.n376 163.367
R1859 B.n377 B.n134 163.367
R1860 B.n381 B.n134 163.367
R1861 B.n382 B.n381 163.367
R1862 B.n383 B.n382 163.367
R1863 B.n383 B.n132 163.367
R1864 B.n387 B.n132 163.367
R1865 B.n388 B.n387 163.367
R1866 B.n389 B.n388 163.367
R1867 B.n389 B.n130 163.367
R1868 B.n393 B.n130 163.367
R1869 B.n394 B.n393 163.367
R1870 B.n395 B.n394 163.367
R1871 B.n395 B.n128 163.367
R1872 B.n399 B.n128 163.367
R1873 B.n400 B.n399 163.367
R1874 B.n401 B.n400 163.367
R1875 B.n401 B.n126 163.367
R1876 B.n405 B.n126 163.367
R1877 B.n406 B.n405 163.367
R1878 B.n407 B.n406 163.367
R1879 B.n407 B.n124 163.367
R1880 B.n411 B.n124 163.367
R1881 B.n412 B.n411 163.367
R1882 B.n413 B.n412 163.367
R1883 B.n413 B.n122 163.367
R1884 B.n417 B.n122 163.367
R1885 B.n418 B.n417 163.367
R1886 B.n419 B.n418 163.367
R1887 B.n419 B.n120 163.367
R1888 B.n423 B.n120 163.367
R1889 B.n424 B.n423 163.367
R1890 B.n425 B.n424 163.367
R1891 B.n425 B.n118 163.367
R1892 B.n429 B.n118 163.367
R1893 B.n431 B.n430 163.367
R1894 B.n431 B.n116 163.367
R1895 B.n435 B.n116 163.367
R1896 B.n436 B.n435 163.367
R1897 B.n437 B.n436 163.367
R1898 B.n437 B.n114 163.367
R1899 B.n441 B.n114 163.367
R1900 B.n442 B.n441 163.367
R1901 B.n443 B.n442 163.367
R1902 B.n443 B.n112 163.367
R1903 B.n447 B.n112 163.367
R1904 B.n448 B.n447 163.367
R1905 B.n449 B.n448 163.367
R1906 B.n449 B.n110 163.367
R1907 B.n453 B.n110 163.367
R1908 B.n454 B.n453 163.367
R1909 B.n455 B.n454 163.367
R1910 B.n455 B.n108 163.367
R1911 B.n459 B.n108 163.367
R1912 B.n460 B.n459 163.367
R1913 B.n461 B.n460 163.367
R1914 B.n461 B.n106 163.367
R1915 B.n465 B.n106 163.367
R1916 B.n466 B.n465 163.367
R1917 B.n467 B.n466 163.367
R1918 B.n467 B.n104 163.367
R1919 B.n471 B.n104 163.367
R1920 B.n472 B.n471 163.367
R1921 B.n473 B.n472 163.367
R1922 B.n473 B.n102 163.367
R1923 B.n477 B.n102 163.367
R1924 B.n478 B.n477 163.367
R1925 B.n479 B.n478 163.367
R1926 B.n479 B.n100 163.367
R1927 B.n483 B.n100 163.367
R1928 B.n484 B.n483 163.367
R1929 B.n485 B.n484 163.367
R1930 B.n485 B.n98 163.367
R1931 B.n489 B.n98 163.367
R1932 B.n490 B.n489 163.367
R1933 B.n491 B.n490 163.367
R1934 B.n491 B.n96 163.367
R1935 B.n495 B.n96 163.367
R1936 B.n496 B.n495 163.367
R1937 B.n497 B.n496 163.367
R1938 B.n497 B.n94 163.367
R1939 B.n501 B.n94 163.367
R1940 B.n502 B.n501 163.367
R1941 B.n503 B.n502 163.367
R1942 B.n503 B.n92 163.367
R1943 B.n507 B.n92 163.367
R1944 B.n508 B.n507 163.367
R1945 B.n509 B.n508 163.367
R1946 B.n509 B.n90 163.367
R1947 B.n513 B.n90 163.367
R1948 B.n514 B.n513 163.367
R1949 B.n515 B.n514 163.367
R1950 B.n515 B.n88 163.367
R1951 B.n519 B.n88 163.367
R1952 B.n520 B.n519 163.367
R1953 B.n521 B.n520 163.367
R1954 B.n521 B.n86 163.367
R1955 B.n525 B.n86 163.367
R1956 B.n526 B.n525 163.367
R1957 B.n527 B.n526 163.367
R1958 B.n527 B.n84 163.367
R1959 B.n712 B.n19 163.367
R1960 B.n708 B.n19 163.367
R1961 B.n708 B.n707 163.367
R1962 B.n707 B.n706 163.367
R1963 B.n706 B.n21 163.367
R1964 B.n702 B.n21 163.367
R1965 B.n702 B.n701 163.367
R1966 B.n701 B.n700 163.367
R1967 B.n700 B.n23 163.367
R1968 B.n696 B.n23 163.367
R1969 B.n696 B.n695 163.367
R1970 B.n695 B.n694 163.367
R1971 B.n694 B.n25 163.367
R1972 B.n690 B.n25 163.367
R1973 B.n690 B.n689 163.367
R1974 B.n689 B.n688 163.367
R1975 B.n688 B.n27 163.367
R1976 B.n684 B.n27 163.367
R1977 B.n684 B.n683 163.367
R1978 B.n683 B.n682 163.367
R1979 B.n682 B.n29 163.367
R1980 B.n678 B.n29 163.367
R1981 B.n678 B.n677 163.367
R1982 B.n677 B.n676 163.367
R1983 B.n676 B.n31 163.367
R1984 B.n672 B.n31 163.367
R1985 B.n672 B.n671 163.367
R1986 B.n671 B.n670 163.367
R1987 B.n670 B.n33 163.367
R1988 B.n666 B.n33 163.367
R1989 B.n666 B.n665 163.367
R1990 B.n665 B.n664 163.367
R1991 B.n664 B.n35 163.367
R1992 B.n660 B.n35 163.367
R1993 B.n660 B.n659 163.367
R1994 B.n659 B.n658 163.367
R1995 B.n658 B.n37 163.367
R1996 B.n654 B.n37 163.367
R1997 B.n654 B.n653 163.367
R1998 B.n653 B.n652 163.367
R1999 B.n652 B.n39 163.367
R2000 B.n648 B.n39 163.367
R2001 B.n648 B.n647 163.367
R2002 B.n647 B.n646 163.367
R2003 B.n646 B.n41 163.367
R2004 B.n642 B.n41 163.367
R2005 B.n642 B.n641 163.367
R2006 B.n641 B.n640 163.367
R2007 B.n640 B.n43 163.367
R2008 B.n636 B.n43 163.367
R2009 B.n636 B.n635 163.367
R2010 B.n635 B.n634 163.367
R2011 B.n634 B.n45 163.367
R2012 B.n630 B.n45 163.367
R2013 B.n630 B.n629 163.367
R2014 B.n629 B.n628 163.367
R2015 B.n628 B.n47 163.367
R2016 B.n624 B.n47 163.367
R2017 B.n624 B.n623 163.367
R2018 B.n623 B.n622 163.367
R2019 B.n622 B.n52 163.367
R2020 B.n618 B.n52 163.367
R2021 B.n618 B.n617 163.367
R2022 B.n617 B.n616 163.367
R2023 B.n616 B.n54 163.367
R2024 B.n611 B.n54 163.367
R2025 B.n611 B.n610 163.367
R2026 B.n610 B.n609 163.367
R2027 B.n609 B.n58 163.367
R2028 B.n605 B.n58 163.367
R2029 B.n605 B.n604 163.367
R2030 B.n604 B.n603 163.367
R2031 B.n603 B.n60 163.367
R2032 B.n599 B.n60 163.367
R2033 B.n599 B.n598 163.367
R2034 B.n598 B.n597 163.367
R2035 B.n597 B.n62 163.367
R2036 B.n593 B.n62 163.367
R2037 B.n593 B.n592 163.367
R2038 B.n592 B.n591 163.367
R2039 B.n591 B.n64 163.367
R2040 B.n587 B.n64 163.367
R2041 B.n587 B.n586 163.367
R2042 B.n586 B.n585 163.367
R2043 B.n585 B.n66 163.367
R2044 B.n581 B.n66 163.367
R2045 B.n581 B.n580 163.367
R2046 B.n580 B.n579 163.367
R2047 B.n579 B.n68 163.367
R2048 B.n575 B.n68 163.367
R2049 B.n575 B.n574 163.367
R2050 B.n574 B.n573 163.367
R2051 B.n573 B.n70 163.367
R2052 B.n569 B.n70 163.367
R2053 B.n569 B.n568 163.367
R2054 B.n568 B.n567 163.367
R2055 B.n567 B.n72 163.367
R2056 B.n563 B.n72 163.367
R2057 B.n563 B.n562 163.367
R2058 B.n562 B.n561 163.367
R2059 B.n561 B.n74 163.367
R2060 B.n557 B.n74 163.367
R2061 B.n557 B.n556 163.367
R2062 B.n556 B.n555 163.367
R2063 B.n555 B.n76 163.367
R2064 B.n551 B.n76 163.367
R2065 B.n551 B.n550 163.367
R2066 B.n550 B.n549 163.367
R2067 B.n549 B.n78 163.367
R2068 B.n545 B.n78 163.367
R2069 B.n545 B.n544 163.367
R2070 B.n544 B.n543 163.367
R2071 B.n543 B.n80 163.367
R2072 B.n539 B.n80 163.367
R2073 B.n539 B.n538 163.367
R2074 B.n538 B.n537 163.367
R2075 B.n537 B.n82 163.367
R2076 B.n533 B.n82 163.367
R2077 B.n533 B.n532 163.367
R2078 B.n532 B.n531 163.367
R2079 B.n343 B.n342 59.5399
R2080 B.n328 B.n152 59.5399
R2081 B.n50 B.n49 59.5399
R2082 B.n614 B.n56 59.5399
R2083 B.n711 B.n18 33.5615
R2084 B.n530 B.n529 33.5615
R2085 B.n428 B.n117 33.5615
R2086 B.n244 B.n243 33.5615
R2087 B.n342 B.n341 33.1641
R2088 B.n152 B.n151 33.1641
R2089 B.n49 B.n48 33.1641
R2090 B.n56 B.n55 33.1641
R2091 B B.n763 18.0485
R2092 B.n711 B.n710 10.6151
R2093 B.n710 B.n709 10.6151
R2094 B.n709 B.n20 10.6151
R2095 B.n705 B.n20 10.6151
R2096 B.n705 B.n704 10.6151
R2097 B.n704 B.n703 10.6151
R2098 B.n703 B.n22 10.6151
R2099 B.n699 B.n22 10.6151
R2100 B.n699 B.n698 10.6151
R2101 B.n698 B.n697 10.6151
R2102 B.n697 B.n24 10.6151
R2103 B.n693 B.n24 10.6151
R2104 B.n693 B.n692 10.6151
R2105 B.n692 B.n691 10.6151
R2106 B.n691 B.n26 10.6151
R2107 B.n687 B.n26 10.6151
R2108 B.n687 B.n686 10.6151
R2109 B.n686 B.n685 10.6151
R2110 B.n685 B.n28 10.6151
R2111 B.n681 B.n28 10.6151
R2112 B.n681 B.n680 10.6151
R2113 B.n680 B.n679 10.6151
R2114 B.n679 B.n30 10.6151
R2115 B.n675 B.n30 10.6151
R2116 B.n675 B.n674 10.6151
R2117 B.n674 B.n673 10.6151
R2118 B.n673 B.n32 10.6151
R2119 B.n669 B.n32 10.6151
R2120 B.n669 B.n668 10.6151
R2121 B.n668 B.n667 10.6151
R2122 B.n667 B.n34 10.6151
R2123 B.n663 B.n34 10.6151
R2124 B.n663 B.n662 10.6151
R2125 B.n662 B.n661 10.6151
R2126 B.n661 B.n36 10.6151
R2127 B.n657 B.n36 10.6151
R2128 B.n657 B.n656 10.6151
R2129 B.n656 B.n655 10.6151
R2130 B.n655 B.n38 10.6151
R2131 B.n651 B.n38 10.6151
R2132 B.n651 B.n650 10.6151
R2133 B.n650 B.n649 10.6151
R2134 B.n649 B.n40 10.6151
R2135 B.n645 B.n40 10.6151
R2136 B.n645 B.n644 10.6151
R2137 B.n644 B.n643 10.6151
R2138 B.n643 B.n42 10.6151
R2139 B.n639 B.n42 10.6151
R2140 B.n639 B.n638 10.6151
R2141 B.n638 B.n637 10.6151
R2142 B.n637 B.n44 10.6151
R2143 B.n633 B.n44 10.6151
R2144 B.n633 B.n632 10.6151
R2145 B.n632 B.n631 10.6151
R2146 B.n631 B.n46 10.6151
R2147 B.n627 B.n626 10.6151
R2148 B.n626 B.n625 10.6151
R2149 B.n625 B.n51 10.6151
R2150 B.n621 B.n51 10.6151
R2151 B.n621 B.n620 10.6151
R2152 B.n620 B.n619 10.6151
R2153 B.n619 B.n53 10.6151
R2154 B.n615 B.n53 10.6151
R2155 B.n613 B.n612 10.6151
R2156 B.n612 B.n57 10.6151
R2157 B.n608 B.n57 10.6151
R2158 B.n608 B.n607 10.6151
R2159 B.n607 B.n606 10.6151
R2160 B.n606 B.n59 10.6151
R2161 B.n602 B.n59 10.6151
R2162 B.n602 B.n601 10.6151
R2163 B.n601 B.n600 10.6151
R2164 B.n600 B.n61 10.6151
R2165 B.n596 B.n61 10.6151
R2166 B.n596 B.n595 10.6151
R2167 B.n595 B.n594 10.6151
R2168 B.n594 B.n63 10.6151
R2169 B.n590 B.n63 10.6151
R2170 B.n590 B.n589 10.6151
R2171 B.n589 B.n588 10.6151
R2172 B.n588 B.n65 10.6151
R2173 B.n584 B.n65 10.6151
R2174 B.n584 B.n583 10.6151
R2175 B.n583 B.n582 10.6151
R2176 B.n582 B.n67 10.6151
R2177 B.n578 B.n67 10.6151
R2178 B.n578 B.n577 10.6151
R2179 B.n577 B.n576 10.6151
R2180 B.n576 B.n69 10.6151
R2181 B.n572 B.n69 10.6151
R2182 B.n572 B.n571 10.6151
R2183 B.n571 B.n570 10.6151
R2184 B.n570 B.n71 10.6151
R2185 B.n566 B.n71 10.6151
R2186 B.n566 B.n565 10.6151
R2187 B.n565 B.n564 10.6151
R2188 B.n564 B.n73 10.6151
R2189 B.n560 B.n73 10.6151
R2190 B.n560 B.n559 10.6151
R2191 B.n559 B.n558 10.6151
R2192 B.n558 B.n75 10.6151
R2193 B.n554 B.n75 10.6151
R2194 B.n554 B.n553 10.6151
R2195 B.n553 B.n552 10.6151
R2196 B.n552 B.n77 10.6151
R2197 B.n548 B.n77 10.6151
R2198 B.n548 B.n547 10.6151
R2199 B.n547 B.n546 10.6151
R2200 B.n546 B.n79 10.6151
R2201 B.n542 B.n79 10.6151
R2202 B.n542 B.n541 10.6151
R2203 B.n541 B.n540 10.6151
R2204 B.n540 B.n81 10.6151
R2205 B.n536 B.n81 10.6151
R2206 B.n536 B.n535 10.6151
R2207 B.n535 B.n534 10.6151
R2208 B.n534 B.n83 10.6151
R2209 B.n530 B.n83 10.6151
R2210 B.n432 B.n117 10.6151
R2211 B.n433 B.n432 10.6151
R2212 B.n434 B.n433 10.6151
R2213 B.n434 B.n115 10.6151
R2214 B.n438 B.n115 10.6151
R2215 B.n439 B.n438 10.6151
R2216 B.n440 B.n439 10.6151
R2217 B.n440 B.n113 10.6151
R2218 B.n444 B.n113 10.6151
R2219 B.n445 B.n444 10.6151
R2220 B.n446 B.n445 10.6151
R2221 B.n446 B.n111 10.6151
R2222 B.n450 B.n111 10.6151
R2223 B.n451 B.n450 10.6151
R2224 B.n452 B.n451 10.6151
R2225 B.n452 B.n109 10.6151
R2226 B.n456 B.n109 10.6151
R2227 B.n457 B.n456 10.6151
R2228 B.n458 B.n457 10.6151
R2229 B.n458 B.n107 10.6151
R2230 B.n462 B.n107 10.6151
R2231 B.n463 B.n462 10.6151
R2232 B.n464 B.n463 10.6151
R2233 B.n464 B.n105 10.6151
R2234 B.n468 B.n105 10.6151
R2235 B.n469 B.n468 10.6151
R2236 B.n470 B.n469 10.6151
R2237 B.n470 B.n103 10.6151
R2238 B.n474 B.n103 10.6151
R2239 B.n475 B.n474 10.6151
R2240 B.n476 B.n475 10.6151
R2241 B.n476 B.n101 10.6151
R2242 B.n480 B.n101 10.6151
R2243 B.n481 B.n480 10.6151
R2244 B.n482 B.n481 10.6151
R2245 B.n482 B.n99 10.6151
R2246 B.n486 B.n99 10.6151
R2247 B.n487 B.n486 10.6151
R2248 B.n488 B.n487 10.6151
R2249 B.n488 B.n97 10.6151
R2250 B.n492 B.n97 10.6151
R2251 B.n493 B.n492 10.6151
R2252 B.n494 B.n493 10.6151
R2253 B.n494 B.n95 10.6151
R2254 B.n498 B.n95 10.6151
R2255 B.n499 B.n498 10.6151
R2256 B.n500 B.n499 10.6151
R2257 B.n500 B.n93 10.6151
R2258 B.n504 B.n93 10.6151
R2259 B.n505 B.n504 10.6151
R2260 B.n506 B.n505 10.6151
R2261 B.n506 B.n91 10.6151
R2262 B.n510 B.n91 10.6151
R2263 B.n511 B.n510 10.6151
R2264 B.n512 B.n511 10.6151
R2265 B.n512 B.n89 10.6151
R2266 B.n516 B.n89 10.6151
R2267 B.n517 B.n516 10.6151
R2268 B.n518 B.n517 10.6151
R2269 B.n518 B.n87 10.6151
R2270 B.n522 B.n87 10.6151
R2271 B.n523 B.n522 10.6151
R2272 B.n524 B.n523 10.6151
R2273 B.n524 B.n85 10.6151
R2274 B.n528 B.n85 10.6151
R2275 B.n529 B.n528 10.6151
R2276 B.n244 B.n179 10.6151
R2277 B.n248 B.n179 10.6151
R2278 B.n249 B.n248 10.6151
R2279 B.n250 B.n249 10.6151
R2280 B.n250 B.n177 10.6151
R2281 B.n254 B.n177 10.6151
R2282 B.n255 B.n254 10.6151
R2283 B.n256 B.n255 10.6151
R2284 B.n256 B.n175 10.6151
R2285 B.n260 B.n175 10.6151
R2286 B.n261 B.n260 10.6151
R2287 B.n262 B.n261 10.6151
R2288 B.n262 B.n173 10.6151
R2289 B.n266 B.n173 10.6151
R2290 B.n267 B.n266 10.6151
R2291 B.n268 B.n267 10.6151
R2292 B.n268 B.n171 10.6151
R2293 B.n272 B.n171 10.6151
R2294 B.n273 B.n272 10.6151
R2295 B.n274 B.n273 10.6151
R2296 B.n274 B.n169 10.6151
R2297 B.n278 B.n169 10.6151
R2298 B.n279 B.n278 10.6151
R2299 B.n280 B.n279 10.6151
R2300 B.n280 B.n167 10.6151
R2301 B.n284 B.n167 10.6151
R2302 B.n285 B.n284 10.6151
R2303 B.n286 B.n285 10.6151
R2304 B.n286 B.n165 10.6151
R2305 B.n290 B.n165 10.6151
R2306 B.n291 B.n290 10.6151
R2307 B.n292 B.n291 10.6151
R2308 B.n292 B.n163 10.6151
R2309 B.n296 B.n163 10.6151
R2310 B.n297 B.n296 10.6151
R2311 B.n298 B.n297 10.6151
R2312 B.n298 B.n161 10.6151
R2313 B.n302 B.n161 10.6151
R2314 B.n303 B.n302 10.6151
R2315 B.n304 B.n303 10.6151
R2316 B.n304 B.n159 10.6151
R2317 B.n308 B.n159 10.6151
R2318 B.n309 B.n308 10.6151
R2319 B.n310 B.n309 10.6151
R2320 B.n310 B.n157 10.6151
R2321 B.n314 B.n157 10.6151
R2322 B.n315 B.n314 10.6151
R2323 B.n316 B.n315 10.6151
R2324 B.n316 B.n155 10.6151
R2325 B.n320 B.n155 10.6151
R2326 B.n321 B.n320 10.6151
R2327 B.n322 B.n321 10.6151
R2328 B.n322 B.n153 10.6151
R2329 B.n326 B.n153 10.6151
R2330 B.n327 B.n326 10.6151
R2331 B.n329 B.n149 10.6151
R2332 B.n333 B.n149 10.6151
R2333 B.n334 B.n333 10.6151
R2334 B.n335 B.n334 10.6151
R2335 B.n335 B.n147 10.6151
R2336 B.n339 B.n147 10.6151
R2337 B.n340 B.n339 10.6151
R2338 B.n344 B.n340 10.6151
R2339 B.n348 B.n145 10.6151
R2340 B.n349 B.n348 10.6151
R2341 B.n350 B.n349 10.6151
R2342 B.n350 B.n143 10.6151
R2343 B.n354 B.n143 10.6151
R2344 B.n355 B.n354 10.6151
R2345 B.n356 B.n355 10.6151
R2346 B.n356 B.n141 10.6151
R2347 B.n360 B.n141 10.6151
R2348 B.n361 B.n360 10.6151
R2349 B.n362 B.n361 10.6151
R2350 B.n362 B.n139 10.6151
R2351 B.n366 B.n139 10.6151
R2352 B.n367 B.n366 10.6151
R2353 B.n368 B.n367 10.6151
R2354 B.n368 B.n137 10.6151
R2355 B.n372 B.n137 10.6151
R2356 B.n373 B.n372 10.6151
R2357 B.n374 B.n373 10.6151
R2358 B.n374 B.n135 10.6151
R2359 B.n378 B.n135 10.6151
R2360 B.n379 B.n378 10.6151
R2361 B.n380 B.n379 10.6151
R2362 B.n380 B.n133 10.6151
R2363 B.n384 B.n133 10.6151
R2364 B.n385 B.n384 10.6151
R2365 B.n386 B.n385 10.6151
R2366 B.n386 B.n131 10.6151
R2367 B.n390 B.n131 10.6151
R2368 B.n391 B.n390 10.6151
R2369 B.n392 B.n391 10.6151
R2370 B.n392 B.n129 10.6151
R2371 B.n396 B.n129 10.6151
R2372 B.n397 B.n396 10.6151
R2373 B.n398 B.n397 10.6151
R2374 B.n398 B.n127 10.6151
R2375 B.n402 B.n127 10.6151
R2376 B.n403 B.n402 10.6151
R2377 B.n404 B.n403 10.6151
R2378 B.n404 B.n125 10.6151
R2379 B.n408 B.n125 10.6151
R2380 B.n409 B.n408 10.6151
R2381 B.n410 B.n409 10.6151
R2382 B.n410 B.n123 10.6151
R2383 B.n414 B.n123 10.6151
R2384 B.n415 B.n414 10.6151
R2385 B.n416 B.n415 10.6151
R2386 B.n416 B.n121 10.6151
R2387 B.n420 B.n121 10.6151
R2388 B.n421 B.n420 10.6151
R2389 B.n422 B.n421 10.6151
R2390 B.n422 B.n119 10.6151
R2391 B.n426 B.n119 10.6151
R2392 B.n427 B.n426 10.6151
R2393 B.n428 B.n427 10.6151
R2394 B.n243 B.n242 10.6151
R2395 B.n242 B.n181 10.6151
R2396 B.n238 B.n181 10.6151
R2397 B.n238 B.n237 10.6151
R2398 B.n237 B.n236 10.6151
R2399 B.n236 B.n183 10.6151
R2400 B.n232 B.n183 10.6151
R2401 B.n232 B.n231 10.6151
R2402 B.n231 B.n230 10.6151
R2403 B.n230 B.n185 10.6151
R2404 B.n226 B.n185 10.6151
R2405 B.n226 B.n225 10.6151
R2406 B.n225 B.n224 10.6151
R2407 B.n224 B.n187 10.6151
R2408 B.n220 B.n187 10.6151
R2409 B.n220 B.n219 10.6151
R2410 B.n219 B.n218 10.6151
R2411 B.n218 B.n189 10.6151
R2412 B.n214 B.n189 10.6151
R2413 B.n214 B.n213 10.6151
R2414 B.n213 B.n212 10.6151
R2415 B.n212 B.n191 10.6151
R2416 B.n208 B.n191 10.6151
R2417 B.n208 B.n207 10.6151
R2418 B.n207 B.n206 10.6151
R2419 B.n206 B.n193 10.6151
R2420 B.n202 B.n193 10.6151
R2421 B.n202 B.n201 10.6151
R2422 B.n201 B.n200 10.6151
R2423 B.n200 B.n195 10.6151
R2424 B.n196 B.n195 10.6151
R2425 B.n196 B.n0 10.6151
R2426 B.n759 B.n1 10.6151
R2427 B.n759 B.n758 10.6151
R2428 B.n758 B.n757 10.6151
R2429 B.n757 B.n4 10.6151
R2430 B.n753 B.n4 10.6151
R2431 B.n753 B.n752 10.6151
R2432 B.n752 B.n751 10.6151
R2433 B.n751 B.n6 10.6151
R2434 B.n747 B.n6 10.6151
R2435 B.n747 B.n746 10.6151
R2436 B.n746 B.n745 10.6151
R2437 B.n745 B.n8 10.6151
R2438 B.n741 B.n8 10.6151
R2439 B.n741 B.n740 10.6151
R2440 B.n740 B.n739 10.6151
R2441 B.n739 B.n10 10.6151
R2442 B.n735 B.n10 10.6151
R2443 B.n735 B.n734 10.6151
R2444 B.n734 B.n733 10.6151
R2445 B.n733 B.n12 10.6151
R2446 B.n729 B.n12 10.6151
R2447 B.n729 B.n728 10.6151
R2448 B.n728 B.n727 10.6151
R2449 B.n727 B.n14 10.6151
R2450 B.n723 B.n14 10.6151
R2451 B.n723 B.n722 10.6151
R2452 B.n722 B.n721 10.6151
R2453 B.n721 B.n16 10.6151
R2454 B.n717 B.n16 10.6151
R2455 B.n717 B.n716 10.6151
R2456 B.n716 B.n715 10.6151
R2457 B.n715 B.n18 10.6151
R2458 B.n627 B.n50 6.5566
R2459 B.n615 B.n614 6.5566
R2460 B.n329 B.n328 6.5566
R2461 B.n344 B.n343 6.5566
R2462 B.n50 B.n46 4.05904
R2463 B.n614 B.n613 4.05904
R2464 B.n328 B.n327 4.05904
R2465 B.n343 B.n145 4.05904
R2466 B.n763 B.n0 2.81026
R2467 B.n763 B.n1 2.81026
C0 w_n2680_n4316# B 9.57606f
C1 VDD2 VP 0.389788f
C2 VP VDD1 10.353f
C3 w_n2680_n4316# VP 5.53692f
C4 VDD2 VTAIL 10.9972f
C5 VTAIL VDD1 10.951f
C6 B VN 0.99949f
C7 w_n2680_n4316# VTAIL 5.28449f
C8 VP VN 7.04215f
C9 VDD2 VDD1 1.16515f
C10 B VP 1.57019f
C11 w_n2680_n4316# VDD2 1.73433f
C12 w_n2680_n4316# VDD1 1.67085f
C13 VN VTAIL 9.92021f
C14 B VTAIL 5.73588f
C15 VDD2 VN 10.1134f
C16 VN VDD1 0.149461f
C17 VP VTAIL 9.93432f
C18 B VDD2 1.46334f
C19 B VDD1 1.40559f
C20 w_n2680_n4316# VN 5.1926f
C21 VDD2 VSUBS 1.597355f
C22 VDD1 VSUBS 2.028994f
C23 VTAIL VSUBS 1.307578f
C24 VN VSUBS 5.54038f
C25 VP VSUBS 2.505455f
C26 B VSUBS 4.042802f
C27 w_n2680_n4316# VSUBS 0.1416p
C28 B.n0 VSUBS 0.004457f
C29 B.n1 VSUBS 0.004457f
C30 B.n2 VSUBS 0.007049f
C31 B.n3 VSUBS 0.007049f
C32 B.n4 VSUBS 0.007049f
C33 B.n5 VSUBS 0.007049f
C34 B.n6 VSUBS 0.007049f
C35 B.n7 VSUBS 0.007049f
C36 B.n8 VSUBS 0.007049f
C37 B.n9 VSUBS 0.007049f
C38 B.n10 VSUBS 0.007049f
C39 B.n11 VSUBS 0.007049f
C40 B.n12 VSUBS 0.007049f
C41 B.n13 VSUBS 0.007049f
C42 B.n14 VSUBS 0.007049f
C43 B.n15 VSUBS 0.007049f
C44 B.n16 VSUBS 0.007049f
C45 B.n17 VSUBS 0.007049f
C46 B.n18 VSUBS 0.01613f
C47 B.n19 VSUBS 0.007049f
C48 B.n20 VSUBS 0.007049f
C49 B.n21 VSUBS 0.007049f
C50 B.n22 VSUBS 0.007049f
C51 B.n23 VSUBS 0.007049f
C52 B.n24 VSUBS 0.007049f
C53 B.n25 VSUBS 0.007049f
C54 B.n26 VSUBS 0.007049f
C55 B.n27 VSUBS 0.007049f
C56 B.n28 VSUBS 0.007049f
C57 B.n29 VSUBS 0.007049f
C58 B.n30 VSUBS 0.007049f
C59 B.n31 VSUBS 0.007049f
C60 B.n32 VSUBS 0.007049f
C61 B.n33 VSUBS 0.007049f
C62 B.n34 VSUBS 0.007049f
C63 B.n35 VSUBS 0.007049f
C64 B.n36 VSUBS 0.007049f
C65 B.n37 VSUBS 0.007049f
C66 B.n38 VSUBS 0.007049f
C67 B.n39 VSUBS 0.007049f
C68 B.n40 VSUBS 0.007049f
C69 B.n41 VSUBS 0.007049f
C70 B.n42 VSUBS 0.007049f
C71 B.n43 VSUBS 0.007049f
C72 B.n44 VSUBS 0.007049f
C73 B.n45 VSUBS 0.007049f
C74 B.n46 VSUBS 0.004872f
C75 B.n47 VSUBS 0.007049f
C76 B.t2 VSUBS 0.322874f
C77 B.t1 VSUBS 0.343054f
C78 B.t0 VSUBS 0.987744f
C79 B.n48 VSUBS 0.480565f
C80 B.n49 VSUBS 0.310677f
C81 B.n50 VSUBS 0.016331f
C82 B.n51 VSUBS 0.007049f
C83 B.n52 VSUBS 0.007049f
C84 B.n53 VSUBS 0.007049f
C85 B.n54 VSUBS 0.007049f
C86 B.t11 VSUBS 0.322877f
C87 B.t10 VSUBS 0.343057f
C88 B.t9 VSUBS 0.987744f
C89 B.n55 VSUBS 0.480561f
C90 B.n56 VSUBS 0.310674f
C91 B.n57 VSUBS 0.007049f
C92 B.n58 VSUBS 0.007049f
C93 B.n59 VSUBS 0.007049f
C94 B.n60 VSUBS 0.007049f
C95 B.n61 VSUBS 0.007049f
C96 B.n62 VSUBS 0.007049f
C97 B.n63 VSUBS 0.007049f
C98 B.n64 VSUBS 0.007049f
C99 B.n65 VSUBS 0.007049f
C100 B.n66 VSUBS 0.007049f
C101 B.n67 VSUBS 0.007049f
C102 B.n68 VSUBS 0.007049f
C103 B.n69 VSUBS 0.007049f
C104 B.n70 VSUBS 0.007049f
C105 B.n71 VSUBS 0.007049f
C106 B.n72 VSUBS 0.007049f
C107 B.n73 VSUBS 0.007049f
C108 B.n74 VSUBS 0.007049f
C109 B.n75 VSUBS 0.007049f
C110 B.n76 VSUBS 0.007049f
C111 B.n77 VSUBS 0.007049f
C112 B.n78 VSUBS 0.007049f
C113 B.n79 VSUBS 0.007049f
C114 B.n80 VSUBS 0.007049f
C115 B.n81 VSUBS 0.007049f
C116 B.n82 VSUBS 0.007049f
C117 B.n83 VSUBS 0.007049f
C118 B.n84 VSUBS 0.01613f
C119 B.n85 VSUBS 0.007049f
C120 B.n86 VSUBS 0.007049f
C121 B.n87 VSUBS 0.007049f
C122 B.n88 VSUBS 0.007049f
C123 B.n89 VSUBS 0.007049f
C124 B.n90 VSUBS 0.007049f
C125 B.n91 VSUBS 0.007049f
C126 B.n92 VSUBS 0.007049f
C127 B.n93 VSUBS 0.007049f
C128 B.n94 VSUBS 0.007049f
C129 B.n95 VSUBS 0.007049f
C130 B.n96 VSUBS 0.007049f
C131 B.n97 VSUBS 0.007049f
C132 B.n98 VSUBS 0.007049f
C133 B.n99 VSUBS 0.007049f
C134 B.n100 VSUBS 0.007049f
C135 B.n101 VSUBS 0.007049f
C136 B.n102 VSUBS 0.007049f
C137 B.n103 VSUBS 0.007049f
C138 B.n104 VSUBS 0.007049f
C139 B.n105 VSUBS 0.007049f
C140 B.n106 VSUBS 0.007049f
C141 B.n107 VSUBS 0.007049f
C142 B.n108 VSUBS 0.007049f
C143 B.n109 VSUBS 0.007049f
C144 B.n110 VSUBS 0.007049f
C145 B.n111 VSUBS 0.007049f
C146 B.n112 VSUBS 0.007049f
C147 B.n113 VSUBS 0.007049f
C148 B.n114 VSUBS 0.007049f
C149 B.n115 VSUBS 0.007049f
C150 B.n116 VSUBS 0.007049f
C151 B.n117 VSUBS 0.01613f
C152 B.n118 VSUBS 0.007049f
C153 B.n119 VSUBS 0.007049f
C154 B.n120 VSUBS 0.007049f
C155 B.n121 VSUBS 0.007049f
C156 B.n122 VSUBS 0.007049f
C157 B.n123 VSUBS 0.007049f
C158 B.n124 VSUBS 0.007049f
C159 B.n125 VSUBS 0.007049f
C160 B.n126 VSUBS 0.007049f
C161 B.n127 VSUBS 0.007049f
C162 B.n128 VSUBS 0.007049f
C163 B.n129 VSUBS 0.007049f
C164 B.n130 VSUBS 0.007049f
C165 B.n131 VSUBS 0.007049f
C166 B.n132 VSUBS 0.007049f
C167 B.n133 VSUBS 0.007049f
C168 B.n134 VSUBS 0.007049f
C169 B.n135 VSUBS 0.007049f
C170 B.n136 VSUBS 0.007049f
C171 B.n137 VSUBS 0.007049f
C172 B.n138 VSUBS 0.007049f
C173 B.n139 VSUBS 0.007049f
C174 B.n140 VSUBS 0.007049f
C175 B.n141 VSUBS 0.007049f
C176 B.n142 VSUBS 0.007049f
C177 B.n143 VSUBS 0.007049f
C178 B.n144 VSUBS 0.007049f
C179 B.n145 VSUBS 0.004872f
C180 B.n146 VSUBS 0.007049f
C181 B.n147 VSUBS 0.007049f
C182 B.n148 VSUBS 0.007049f
C183 B.n149 VSUBS 0.007049f
C184 B.n150 VSUBS 0.007049f
C185 B.t7 VSUBS 0.322874f
C186 B.t8 VSUBS 0.343054f
C187 B.t6 VSUBS 0.987744f
C188 B.n151 VSUBS 0.480565f
C189 B.n152 VSUBS 0.310677f
C190 B.n153 VSUBS 0.007049f
C191 B.n154 VSUBS 0.007049f
C192 B.n155 VSUBS 0.007049f
C193 B.n156 VSUBS 0.007049f
C194 B.n157 VSUBS 0.007049f
C195 B.n158 VSUBS 0.007049f
C196 B.n159 VSUBS 0.007049f
C197 B.n160 VSUBS 0.007049f
C198 B.n161 VSUBS 0.007049f
C199 B.n162 VSUBS 0.007049f
C200 B.n163 VSUBS 0.007049f
C201 B.n164 VSUBS 0.007049f
C202 B.n165 VSUBS 0.007049f
C203 B.n166 VSUBS 0.007049f
C204 B.n167 VSUBS 0.007049f
C205 B.n168 VSUBS 0.007049f
C206 B.n169 VSUBS 0.007049f
C207 B.n170 VSUBS 0.007049f
C208 B.n171 VSUBS 0.007049f
C209 B.n172 VSUBS 0.007049f
C210 B.n173 VSUBS 0.007049f
C211 B.n174 VSUBS 0.007049f
C212 B.n175 VSUBS 0.007049f
C213 B.n176 VSUBS 0.007049f
C214 B.n177 VSUBS 0.007049f
C215 B.n178 VSUBS 0.007049f
C216 B.n179 VSUBS 0.007049f
C217 B.n180 VSUBS 0.01613f
C218 B.n181 VSUBS 0.007049f
C219 B.n182 VSUBS 0.007049f
C220 B.n183 VSUBS 0.007049f
C221 B.n184 VSUBS 0.007049f
C222 B.n185 VSUBS 0.007049f
C223 B.n186 VSUBS 0.007049f
C224 B.n187 VSUBS 0.007049f
C225 B.n188 VSUBS 0.007049f
C226 B.n189 VSUBS 0.007049f
C227 B.n190 VSUBS 0.007049f
C228 B.n191 VSUBS 0.007049f
C229 B.n192 VSUBS 0.007049f
C230 B.n193 VSUBS 0.007049f
C231 B.n194 VSUBS 0.007049f
C232 B.n195 VSUBS 0.007049f
C233 B.n196 VSUBS 0.007049f
C234 B.n197 VSUBS 0.007049f
C235 B.n198 VSUBS 0.007049f
C236 B.n199 VSUBS 0.007049f
C237 B.n200 VSUBS 0.007049f
C238 B.n201 VSUBS 0.007049f
C239 B.n202 VSUBS 0.007049f
C240 B.n203 VSUBS 0.007049f
C241 B.n204 VSUBS 0.007049f
C242 B.n205 VSUBS 0.007049f
C243 B.n206 VSUBS 0.007049f
C244 B.n207 VSUBS 0.007049f
C245 B.n208 VSUBS 0.007049f
C246 B.n209 VSUBS 0.007049f
C247 B.n210 VSUBS 0.007049f
C248 B.n211 VSUBS 0.007049f
C249 B.n212 VSUBS 0.007049f
C250 B.n213 VSUBS 0.007049f
C251 B.n214 VSUBS 0.007049f
C252 B.n215 VSUBS 0.007049f
C253 B.n216 VSUBS 0.007049f
C254 B.n217 VSUBS 0.007049f
C255 B.n218 VSUBS 0.007049f
C256 B.n219 VSUBS 0.007049f
C257 B.n220 VSUBS 0.007049f
C258 B.n221 VSUBS 0.007049f
C259 B.n222 VSUBS 0.007049f
C260 B.n223 VSUBS 0.007049f
C261 B.n224 VSUBS 0.007049f
C262 B.n225 VSUBS 0.007049f
C263 B.n226 VSUBS 0.007049f
C264 B.n227 VSUBS 0.007049f
C265 B.n228 VSUBS 0.007049f
C266 B.n229 VSUBS 0.007049f
C267 B.n230 VSUBS 0.007049f
C268 B.n231 VSUBS 0.007049f
C269 B.n232 VSUBS 0.007049f
C270 B.n233 VSUBS 0.007049f
C271 B.n234 VSUBS 0.007049f
C272 B.n235 VSUBS 0.007049f
C273 B.n236 VSUBS 0.007049f
C274 B.n237 VSUBS 0.007049f
C275 B.n238 VSUBS 0.007049f
C276 B.n239 VSUBS 0.007049f
C277 B.n240 VSUBS 0.007049f
C278 B.n241 VSUBS 0.007049f
C279 B.n242 VSUBS 0.007049f
C280 B.n243 VSUBS 0.01613f
C281 B.n244 VSUBS 0.017454f
C282 B.n245 VSUBS 0.017454f
C283 B.n246 VSUBS 0.007049f
C284 B.n247 VSUBS 0.007049f
C285 B.n248 VSUBS 0.007049f
C286 B.n249 VSUBS 0.007049f
C287 B.n250 VSUBS 0.007049f
C288 B.n251 VSUBS 0.007049f
C289 B.n252 VSUBS 0.007049f
C290 B.n253 VSUBS 0.007049f
C291 B.n254 VSUBS 0.007049f
C292 B.n255 VSUBS 0.007049f
C293 B.n256 VSUBS 0.007049f
C294 B.n257 VSUBS 0.007049f
C295 B.n258 VSUBS 0.007049f
C296 B.n259 VSUBS 0.007049f
C297 B.n260 VSUBS 0.007049f
C298 B.n261 VSUBS 0.007049f
C299 B.n262 VSUBS 0.007049f
C300 B.n263 VSUBS 0.007049f
C301 B.n264 VSUBS 0.007049f
C302 B.n265 VSUBS 0.007049f
C303 B.n266 VSUBS 0.007049f
C304 B.n267 VSUBS 0.007049f
C305 B.n268 VSUBS 0.007049f
C306 B.n269 VSUBS 0.007049f
C307 B.n270 VSUBS 0.007049f
C308 B.n271 VSUBS 0.007049f
C309 B.n272 VSUBS 0.007049f
C310 B.n273 VSUBS 0.007049f
C311 B.n274 VSUBS 0.007049f
C312 B.n275 VSUBS 0.007049f
C313 B.n276 VSUBS 0.007049f
C314 B.n277 VSUBS 0.007049f
C315 B.n278 VSUBS 0.007049f
C316 B.n279 VSUBS 0.007049f
C317 B.n280 VSUBS 0.007049f
C318 B.n281 VSUBS 0.007049f
C319 B.n282 VSUBS 0.007049f
C320 B.n283 VSUBS 0.007049f
C321 B.n284 VSUBS 0.007049f
C322 B.n285 VSUBS 0.007049f
C323 B.n286 VSUBS 0.007049f
C324 B.n287 VSUBS 0.007049f
C325 B.n288 VSUBS 0.007049f
C326 B.n289 VSUBS 0.007049f
C327 B.n290 VSUBS 0.007049f
C328 B.n291 VSUBS 0.007049f
C329 B.n292 VSUBS 0.007049f
C330 B.n293 VSUBS 0.007049f
C331 B.n294 VSUBS 0.007049f
C332 B.n295 VSUBS 0.007049f
C333 B.n296 VSUBS 0.007049f
C334 B.n297 VSUBS 0.007049f
C335 B.n298 VSUBS 0.007049f
C336 B.n299 VSUBS 0.007049f
C337 B.n300 VSUBS 0.007049f
C338 B.n301 VSUBS 0.007049f
C339 B.n302 VSUBS 0.007049f
C340 B.n303 VSUBS 0.007049f
C341 B.n304 VSUBS 0.007049f
C342 B.n305 VSUBS 0.007049f
C343 B.n306 VSUBS 0.007049f
C344 B.n307 VSUBS 0.007049f
C345 B.n308 VSUBS 0.007049f
C346 B.n309 VSUBS 0.007049f
C347 B.n310 VSUBS 0.007049f
C348 B.n311 VSUBS 0.007049f
C349 B.n312 VSUBS 0.007049f
C350 B.n313 VSUBS 0.007049f
C351 B.n314 VSUBS 0.007049f
C352 B.n315 VSUBS 0.007049f
C353 B.n316 VSUBS 0.007049f
C354 B.n317 VSUBS 0.007049f
C355 B.n318 VSUBS 0.007049f
C356 B.n319 VSUBS 0.007049f
C357 B.n320 VSUBS 0.007049f
C358 B.n321 VSUBS 0.007049f
C359 B.n322 VSUBS 0.007049f
C360 B.n323 VSUBS 0.007049f
C361 B.n324 VSUBS 0.007049f
C362 B.n325 VSUBS 0.007049f
C363 B.n326 VSUBS 0.007049f
C364 B.n327 VSUBS 0.004872f
C365 B.n328 VSUBS 0.016331f
C366 B.n329 VSUBS 0.005701f
C367 B.n330 VSUBS 0.007049f
C368 B.n331 VSUBS 0.007049f
C369 B.n332 VSUBS 0.007049f
C370 B.n333 VSUBS 0.007049f
C371 B.n334 VSUBS 0.007049f
C372 B.n335 VSUBS 0.007049f
C373 B.n336 VSUBS 0.007049f
C374 B.n337 VSUBS 0.007049f
C375 B.n338 VSUBS 0.007049f
C376 B.n339 VSUBS 0.007049f
C377 B.n340 VSUBS 0.007049f
C378 B.t4 VSUBS 0.322877f
C379 B.t5 VSUBS 0.343057f
C380 B.t3 VSUBS 0.987744f
C381 B.n341 VSUBS 0.480561f
C382 B.n342 VSUBS 0.310674f
C383 B.n343 VSUBS 0.016331f
C384 B.n344 VSUBS 0.005701f
C385 B.n345 VSUBS 0.007049f
C386 B.n346 VSUBS 0.007049f
C387 B.n347 VSUBS 0.007049f
C388 B.n348 VSUBS 0.007049f
C389 B.n349 VSUBS 0.007049f
C390 B.n350 VSUBS 0.007049f
C391 B.n351 VSUBS 0.007049f
C392 B.n352 VSUBS 0.007049f
C393 B.n353 VSUBS 0.007049f
C394 B.n354 VSUBS 0.007049f
C395 B.n355 VSUBS 0.007049f
C396 B.n356 VSUBS 0.007049f
C397 B.n357 VSUBS 0.007049f
C398 B.n358 VSUBS 0.007049f
C399 B.n359 VSUBS 0.007049f
C400 B.n360 VSUBS 0.007049f
C401 B.n361 VSUBS 0.007049f
C402 B.n362 VSUBS 0.007049f
C403 B.n363 VSUBS 0.007049f
C404 B.n364 VSUBS 0.007049f
C405 B.n365 VSUBS 0.007049f
C406 B.n366 VSUBS 0.007049f
C407 B.n367 VSUBS 0.007049f
C408 B.n368 VSUBS 0.007049f
C409 B.n369 VSUBS 0.007049f
C410 B.n370 VSUBS 0.007049f
C411 B.n371 VSUBS 0.007049f
C412 B.n372 VSUBS 0.007049f
C413 B.n373 VSUBS 0.007049f
C414 B.n374 VSUBS 0.007049f
C415 B.n375 VSUBS 0.007049f
C416 B.n376 VSUBS 0.007049f
C417 B.n377 VSUBS 0.007049f
C418 B.n378 VSUBS 0.007049f
C419 B.n379 VSUBS 0.007049f
C420 B.n380 VSUBS 0.007049f
C421 B.n381 VSUBS 0.007049f
C422 B.n382 VSUBS 0.007049f
C423 B.n383 VSUBS 0.007049f
C424 B.n384 VSUBS 0.007049f
C425 B.n385 VSUBS 0.007049f
C426 B.n386 VSUBS 0.007049f
C427 B.n387 VSUBS 0.007049f
C428 B.n388 VSUBS 0.007049f
C429 B.n389 VSUBS 0.007049f
C430 B.n390 VSUBS 0.007049f
C431 B.n391 VSUBS 0.007049f
C432 B.n392 VSUBS 0.007049f
C433 B.n393 VSUBS 0.007049f
C434 B.n394 VSUBS 0.007049f
C435 B.n395 VSUBS 0.007049f
C436 B.n396 VSUBS 0.007049f
C437 B.n397 VSUBS 0.007049f
C438 B.n398 VSUBS 0.007049f
C439 B.n399 VSUBS 0.007049f
C440 B.n400 VSUBS 0.007049f
C441 B.n401 VSUBS 0.007049f
C442 B.n402 VSUBS 0.007049f
C443 B.n403 VSUBS 0.007049f
C444 B.n404 VSUBS 0.007049f
C445 B.n405 VSUBS 0.007049f
C446 B.n406 VSUBS 0.007049f
C447 B.n407 VSUBS 0.007049f
C448 B.n408 VSUBS 0.007049f
C449 B.n409 VSUBS 0.007049f
C450 B.n410 VSUBS 0.007049f
C451 B.n411 VSUBS 0.007049f
C452 B.n412 VSUBS 0.007049f
C453 B.n413 VSUBS 0.007049f
C454 B.n414 VSUBS 0.007049f
C455 B.n415 VSUBS 0.007049f
C456 B.n416 VSUBS 0.007049f
C457 B.n417 VSUBS 0.007049f
C458 B.n418 VSUBS 0.007049f
C459 B.n419 VSUBS 0.007049f
C460 B.n420 VSUBS 0.007049f
C461 B.n421 VSUBS 0.007049f
C462 B.n422 VSUBS 0.007049f
C463 B.n423 VSUBS 0.007049f
C464 B.n424 VSUBS 0.007049f
C465 B.n425 VSUBS 0.007049f
C466 B.n426 VSUBS 0.007049f
C467 B.n427 VSUBS 0.007049f
C468 B.n428 VSUBS 0.017454f
C469 B.n429 VSUBS 0.017454f
C470 B.n430 VSUBS 0.01613f
C471 B.n431 VSUBS 0.007049f
C472 B.n432 VSUBS 0.007049f
C473 B.n433 VSUBS 0.007049f
C474 B.n434 VSUBS 0.007049f
C475 B.n435 VSUBS 0.007049f
C476 B.n436 VSUBS 0.007049f
C477 B.n437 VSUBS 0.007049f
C478 B.n438 VSUBS 0.007049f
C479 B.n439 VSUBS 0.007049f
C480 B.n440 VSUBS 0.007049f
C481 B.n441 VSUBS 0.007049f
C482 B.n442 VSUBS 0.007049f
C483 B.n443 VSUBS 0.007049f
C484 B.n444 VSUBS 0.007049f
C485 B.n445 VSUBS 0.007049f
C486 B.n446 VSUBS 0.007049f
C487 B.n447 VSUBS 0.007049f
C488 B.n448 VSUBS 0.007049f
C489 B.n449 VSUBS 0.007049f
C490 B.n450 VSUBS 0.007049f
C491 B.n451 VSUBS 0.007049f
C492 B.n452 VSUBS 0.007049f
C493 B.n453 VSUBS 0.007049f
C494 B.n454 VSUBS 0.007049f
C495 B.n455 VSUBS 0.007049f
C496 B.n456 VSUBS 0.007049f
C497 B.n457 VSUBS 0.007049f
C498 B.n458 VSUBS 0.007049f
C499 B.n459 VSUBS 0.007049f
C500 B.n460 VSUBS 0.007049f
C501 B.n461 VSUBS 0.007049f
C502 B.n462 VSUBS 0.007049f
C503 B.n463 VSUBS 0.007049f
C504 B.n464 VSUBS 0.007049f
C505 B.n465 VSUBS 0.007049f
C506 B.n466 VSUBS 0.007049f
C507 B.n467 VSUBS 0.007049f
C508 B.n468 VSUBS 0.007049f
C509 B.n469 VSUBS 0.007049f
C510 B.n470 VSUBS 0.007049f
C511 B.n471 VSUBS 0.007049f
C512 B.n472 VSUBS 0.007049f
C513 B.n473 VSUBS 0.007049f
C514 B.n474 VSUBS 0.007049f
C515 B.n475 VSUBS 0.007049f
C516 B.n476 VSUBS 0.007049f
C517 B.n477 VSUBS 0.007049f
C518 B.n478 VSUBS 0.007049f
C519 B.n479 VSUBS 0.007049f
C520 B.n480 VSUBS 0.007049f
C521 B.n481 VSUBS 0.007049f
C522 B.n482 VSUBS 0.007049f
C523 B.n483 VSUBS 0.007049f
C524 B.n484 VSUBS 0.007049f
C525 B.n485 VSUBS 0.007049f
C526 B.n486 VSUBS 0.007049f
C527 B.n487 VSUBS 0.007049f
C528 B.n488 VSUBS 0.007049f
C529 B.n489 VSUBS 0.007049f
C530 B.n490 VSUBS 0.007049f
C531 B.n491 VSUBS 0.007049f
C532 B.n492 VSUBS 0.007049f
C533 B.n493 VSUBS 0.007049f
C534 B.n494 VSUBS 0.007049f
C535 B.n495 VSUBS 0.007049f
C536 B.n496 VSUBS 0.007049f
C537 B.n497 VSUBS 0.007049f
C538 B.n498 VSUBS 0.007049f
C539 B.n499 VSUBS 0.007049f
C540 B.n500 VSUBS 0.007049f
C541 B.n501 VSUBS 0.007049f
C542 B.n502 VSUBS 0.007049f
C543 B.n503 VSUBS 0.007049f
C544 B.n504 VSUBS 0.007049f
C545 B.n505 VSUBS 0.007049f
C546 B.n506 VSUBS 0.007049f
C547 B.n507 VSUBS 0.007049f
C548 B.n508 VSUBS 0.007049f
C549 B.n509 VSUBS 0.007049f
C550 B.n510 VSUBS 0.007049f
C551 B.n511 VSUBS 0.007049f
C552 B.n512 VSUBS 0.007049f
C553 B.n513 VSUBS 0.007049f
C554 B.n514 VSUBS 0.007049f
C555 B.n515 VSUBS 0.007049f
C556 B.n516 VSUBS 0.007049f
C557 B.n517 VSUBS 0.007049f
C558 B.n518 VSUBS 0.007049f
C559 B.n519 VSUBS 0.007049f
C560 B.n520 VSUBS 0.007049f
C561 B.n521 VSUBS 0.007049f
C562 B.n522 VSUBS 0.007049f
C563 B.n523 VSUBS 0.007049f
C564 B.n524 VSUBS 0.007049f
C565 B.n525 VSUBS 0.007049f
C566 B.n526 VSUBS 0.007049f
C567 B.n527 VSUBS 0.007049f
C568 B.n528 VSUBS 0.007049f
C569 B.n529 VSUBS 0.016941f
C570 B.n530 VSUBS 0.016644f
C571 B.n531 VSUBS 0.017454f
C572 B.n532 VSUBS 0.007049f
C573 B.n533 VSUBS 0.007049f
C574 B.n534 VSUBS 0.007049f
C575 B.n535 VSUBS 0.007049f
C576 B.n536 VSUBS 0.007049f
C577 B.n537 VSUBS 0.007049f
C578 B.n538 VSUBS 0.007049f
C579 B.n539 VSUBS 0.007049f
C580 B.n540 VSUBS 0.007049f
C581 B.n541 VSUBS 0.007049f
C582 B.n542 VSUBS 0.007049f
C583 B.n543 VSUBS 0.007049f
C584 B.n544 VSUBS 0.007049f
C585 B.n545 VSUBS 0.007049f
C586 B.n546 VSUBS 0.007049f
C587 B.n547 VSUBS 0.007049f
C588 B.n548 VSUBS 0.007049f
C589 B.n549 VSUBS 0.007049f
C590 B.n550 VSUBS 0.007049f
C591 B.n551 VSUBS 0.007049f
C592 B.n552 VSUBS 0.007049f
C593 B.n553 VSUBS 0.007049f
C594 B.n554 VSUBS 0.007049f
C595 B.n555 VSUBS 0.007049f
C596 B.n556 VSUBS 0.007049f
C597 B.n557 VSUBS 0.007049f
C598 B.n558 VSUBS 0.007049f
C599 B.n559 VSUBS 0.007049f
C600 B.n560 VSUBS 0.007049f
C601 B.n561 VSUBS 0.007049f
C602 B.n562 VSUBS 0.007049f
C603 B.n563 VSUBS 0.007049f
C604 B.n564 VSUBS 0.007049f
C605 B.n565 VSUBS 0.007049f
C606 B.n566 VSUBS 0.007049f
C607 B.n567 VSUBS 0.007049f
C608 B.n568 VSUBS 0.007049f
C609 B.n569 VSUBS 0.007049f
C610 B.n570 VSUBS 0.007049f
C611 B.n571 VSUBS 0.007049f
C612 B.n572 VSUBS 0.007049f
C613 B.n573 VSUBS 0.007049f
C614 B.n574 VSUBS 0.007049f
C615 B.n575 VSUBS 0.007049f
C616 B.n576 VSUBS 0.007049f
C617 B.n577 VSUBS 0.007049f
C618 B.n578 VSUBS 0.007049f
C619 B.n579 VSUBS 0.007049f
C620 B.n580 VSUBS 0.007049f
C621 B.n581 VSUBS 0.007049f
C622 B.n582 VSUBS 0.007049f
C623 B.n583 VSUBS 0.007049f
C624 B.n584 VSUBS 0.007049f
C625 B.n585 VSUBS 0.007049f
C626 B.n586 VSUBS 0.007049f
C627 B.n587 VSUBS 0.007049f
C628 B.n588 VSUBS 0.007049f
C629 B.n589 VSUBS 0.007049f
C630 B.n590 VSUBS 0.007049f
C631 B.n591 VSUBS 0.007049f
C632 B.n592 VSUBS 0.007049f
C633 B.n593 VSUBS 0.007049f
C634 B.n594 VSUBS 0.007049f
C635 B.n595 VSUBS 0.007049f
C636 B.n596 VSUBS 0.007049f
C637 B.n597 VSUBS 0.007049f
C638 B.n598 VSUBS 0.007049f
C639 B.n599 VSUBS 0.007049f
C640 B.n600 VSUBS 0.007049f
C641 B.n601 VSUBS 0.007049f
C642 B.n602 VSUBS 0.007049f
C643 B.n603 VSUBS 0.007049f
C644 B.n604 VSUBS 0.007049f
C645 B.n605 VSUBS 0.007049f
C646 B.n606 VSUBS 0.007049f
C647 B.n607 VSUBS 0.007049f
C648 B.n608 VSUBS 0.007049f
C649 B.n609 VSUBS 0.007049f
C650 B.n610 VSUBS 0.007049f
C651 B.n611 VSUBS 0.007049f
C652 B.n612 VSUBS 0.007049f
C653 B.n613 VSUBS 0.004872f
C654 B.n614 VSUBS 0.016331f
C655 B.n615 VSUBS 0.005701f
C656 B.n616 VSUBS 0.007049f
C657 B.n617 VSUBS 0.007049f
C658 B.n618 VSUBS 0.007049f
C659 B.n619 VSUBS 0.007049f
C660 B.n620 VSUBS 0.007049f
C661 B.n621 VSUBS 0.007049f
C662 B.n622 VSUBS 0.007049f
C663 B.n623 VSUBS 0.007049f
C664 B.n624 VSUBS 0.007049f
C665 B.n625 VSUBS 0.007049f
C666 B.n626 VSUBS 0.007049f
C667 B.n627 VSUBS 0.005701f
C668 B.n628 VSUBS 0.007049f
C669 B.n629 VSUBS 0.007049f
C670 B.n630 VSUBS 0.007049f
C671 B.n631 VSUBS 0.007049f
C672 B.n632 VSUBS 0.007049f
C673 B.n633 VSUBS 0.007049f
C674 B.n634 VSUBS 0.007049f
C675 B.n635 VSUBS 0.007049f
C676 B.n636 VSUBS 0.007049f
C677 B.n637 VSUBS 0.007049f
C678 B.n638 VSUBS 0.007049f
C679 B.n639 VSUBS 0.007049f
C680 B.n640 VSUBS 0.007049f
C681 B.n641 VSUBS 0.007049f
C682 B.n642 VSUBS 0.007049f
C683 B.n643 VSUBS 0.007049f
C684 B.n644 VSUBS 0.007049f
C685 B.n645 VSUBS 0.007049f
C686 B.n646 VSUBS 0.007049f
C687 B.n647 VSUBS 0.007049f
C688 B.n648 VSUBS 0.007049f
C689 B.n649 VSUBS 0.007049f
C690 B.n650 VSUBS 0.007049f
C691 B.n651 VSUBS 0.007049f
C692 B.n652 VSUBS 0.007049f
C693 B.n653 VSUBS 0.007049f
C694 B.n654 VSUBS 0.007049f
C695 B.n655 VSUBS 0.007049f
C696 B.n656 VSUBS 0.007049f
C697 B.n657 VSUBS 0.007049f
C698 B.n658 VSUBS 0.007049f
C699 B.n659 VSUBS 0.007049f
C700 B.n660 VSUBS 0.007049f
C701 B.n661 VSUBS 0.007049f
C702 B.n662 VSUBS 0.007049f
C703 B.n663 VSUBS 0.007049f
C704 B.n664 VSUBS 0.007049f
C705 B.n665 VSUBS 0.007049f
C706 B.n666 VSUBS 0.007049f
C707 B.n667 VSUBS 0.007049f
C708 B.n668 VSUBS 0.007049f
C709 B.n669 VSUBS 0.007049f
C710 B.n670 VSUBS 0.007049f
C711 B.n671 VSUBS 0.007049f
C712 B.n672 VSUBS 0.007049f
C713 B.n673 VSUBS 0.007049f
C714 B.n674 VSUBS 0.007049f
C715 B.n675 VSUBS 0.007049f
C716 B.n676 VSUBS 0.007049f
C717 B.n677 VSUBS 0.007049f
C718 B.n678 VSUBS 0.007049f
C719 B.n679 VSUBS 0.007049f
C720 B.n680 VSUBS 0.007049f
C721 B.n681 VSUBS 0.007049f
C722 B.n682 VSUBS 0.007049f
C723 B.n683 VSUBS 0.007049f
C724 B.n684 VSUBS 0.007049f
C725 B.n685 VSUBS 0.007049f
C726 B.n686 VSUBS 0.007049f
C727 B.n687 VSUBS 0.007049f
C728 B.n688 VSUBS 0.007049f
C729 B.n689 VSUBS 0.007049f
C730 B.n690 VSUBS 0.007049f
C731 B.n691 VSUBS 0.007049f
C732 B.n692 VSUBS 0.007049f
C733 B.n693 VSUBS 0.007049f
C734 B.n694 VSUBS 0.007049f
C735 B.n695 VSUBS 0.007049f
C736 B.n696 VSUBS 0.007049f
C737 B.n697 VSUBS 0.007049f
C738 B.n698 VSUBS 0.007049f
C739 B.n699 VSUBS 0.007049f
C740 B.n700 VSUBS 0.007049f
C741 B.n701 VSUBS 0.007049f
C742 B.n702 VSUBS 0.007049f
C743 B.n703 VSUBS 0.007049f
C744 B.n704 VSUBS 0.007049f
C745 B.n705 VSUBS 0.007049f
C746 B.n706 VSUBS 0.007049f
C747 B.n707 VSUBS 0.007049f
C748 B.n708 VSUBS 0.007049f
C749 B.n709 VSUBS 0.007049f
C750 B.n710 VSUBS 0.007049f
C751 B.n711 VSUBS 0.017454f
C752 B.n712 VSUBS 0.017454f
C753 B.n713 VSUBS 0.01613f
C754 B.n714 VSUBS 0.007049f
C755 B.n715 VSUBS 0.007049f
C756 B.n716 VSUBS 0.007049f
C757 B.n717 VSUBS 0.007049f
C758 B.n718 VSUBS 0.007049f
C759 B.n719 VSUBS 0.007049f
C760 B.n720 VSUBS 0.007049f
C761 B.n721 VSUBS 0.007049f
C762 B.n722 VSUBS 0.007049f
C763 B.n723 VSUBS 0.007049f
C764 B.n724 VSUBS 0.007049f
C765 B.n725 VSUBS 0.007049f
C766 B.n726 VSUBS 0.007049f
C767 B.n727 VSUBS 0.007049f
C768 B.n728 VSUBS 0.007049f
C769 B.n729 VSUBS 0.007049f
C770 B.n730 VSUBS 0.007049f
C771 B.n731 VSUBS 0.007049f
C772 B.n732 VSUBS 0.007049f
C773 B.n733 VSUBS 0.007049f
C774 B.n734 VSUBS 0.007049f
C775 B.n735 VSUBS 0.007049f
C776 B.n736 VSUBS 0.007049f
C777 B.n737 VSUBS 0.007049f
C778 B.n738 VSUBS 0.007049f
C779 B.n739 VSUBS 0.007049f
C780 B.n740 VSUBS 0.007049f
C781 B.n741 VSUBS 0.007049f
C782 B.n742 VSUBS 0.007049f
C783 B.n743 VSUBS 0.007049f
C784 B.n744 VSUBS 0.007049f
C785 B.n745 VSUBS 0.007049f
C786 B.n746 VSUBS 0.007049f
C787 B.n747 VSUBS 0.007049f
C788 B.n748 VSUBS 0.007049f
C789 B.n749 VSUBS 0.007049f
C790 B.n750 VSUBS 0.007049f
C791 B.n751 VSUBS 0.007049f
C792 B.n752 VSUBS 0.007049f
C793 B.n753 VSUBS 0.007049f
C794 B.n754 VSUBS 0.007049f
C795 B.n755 VSUBS 0.007049f
C796 B.n756 VSUBS 0.007049f
C797 B.n757 VSUBS 0.007049f
C798 B.n758 VSUBS 0.007049f
C799 B.n759 VSUBS 0.007049f
C800 B.n760 VSUBS 0.007049f
C801 B.n761 VSUBS 0.007049f
C802 B.n762 VSUBS 0.007049f
C803 B.n763 VSUBS 0.015961f
C804 VDD1.t4 VSUBS 0.336585f
C805 VDD1.t0 VSUBS 0.336585f
C806 VDD1.n0 VSUBS 2.77304f
C807 VDD1.t7 VSUBS 0.336585f
C808 VDD1.t6 VSUBS 0.336585f
C809 VDD1.n1 VSUBS 2.7718f
C810 VDD1.t2 VSUBS 0.336585f
C811 VDD1.t3 VSUBS 0.336585f
C812 VDD1.n2 VSUBS 2.7718f
C813 VDD1.n3 VSUBS 3.55009f
C814 VDD1.t5 VSUBS 0.336585f
C815 VDD1.t1 VSUBS 0.336585f
C816 VDD1.n4 VSUBS 2.76497f
C817 VDD1.n5 VSUBS 3.26408f
C818 VP.n0 VSUBS 0.03851f
C819 VP.t4 VSUBS 2.44352f
C820 VP.n1 VSUBS 0.066845f
C821 VP.n2 VSUBS 0.03851f
C822 VP.n3 VSUBS 0.043562f
C823 VP.n4 VSUBS 0.03851f
C824 VP.t0 VSUBS 2.44352f
C825 VP.n5 VSUBS 0.946927f
C826 VP.n6 VSUBS 0.03851f
C827 VP.t6 VSUBS 2.44352f
C828 VP.n7 VSUBS 0.066845f
C829 VP.n8 VSUBS 0.03851f
C830 VP.n9 VSUBS 0.043562f
C831 VP.t3 VSUBS 2.53979f
C832 VP.t7 VSUBS 2.44352f
C833 VP.n10 VSUBS 0.921793f
C834 VP.n11 VSUBS 0.960151f
C835 VP.n12 VSUBS 0.207162f
C836 VP.n13 VSUBS 0.03851f
C837 VP.n14 VSUBS 0.055981f
C838 VP.n15 VSUBS 0.055981f
C839 VP.t2 VSUBS 2.44352f
C840 VP.n16 VSUBS 0.866311f
C841 VP.n17 VSUBS 0.043562f
C842 VP.n18 VSUBS 0.03851f
C843 VP.n19 VSUBS 0.03851f
C844 VP.n20 VSUBS 0.03851f
C845 VP.n21 VSUBS 0.031896f
C846 VP.n22 VSUBS 0.064186f
C847 VP.n23 VSUBS 0.946927f
C848 VP.n24 VSUBS 2.01999f
C849 VP.n25 VSUBS 2.04846f
C850 VP.n26 VSUBS 0.03851f
C851 VP.n27 VSUBS 0.064186f
C852 VP.n28 VSUBS 0.031896f
C853 VP.t1 VSUBS 2.44352f
C854 VP.n29 VSUBS 0.866311f
C855 VP.n30 VSUBS 0.066845f
C856 VP.n31 VSUBS 0.03851f
C857 VP.n32 VSUBS 0.03851f
C858 VP.n33 VSUBS 0.03851f
C859 VP.n34 VSUBS 0.055981f
C860 VP.n35 VSUBS 0.055981f
C861 VP.t5 VSUBS 2.44352f
C862 VP.n36 VSUBS 0.866311f
C863 VP.n37 VSUBS 0.043562f
C864 VP.n38 VSUBS 0.03851f
C865 VP.n39 VSUBS 0.03851f
C866 VP.n40 VSUBS 0.03851f
C867 VP.n41 VSUBS 0.031896f
C868 VP.n42 VSUBS 0.064186f
C869 VP.n43 VSUBS 0.946927f
C870 VP.n44 VSUBS 0.034392f
C871 VTAIL.t11 VSUBS 0.308984f
C872 VTAIL.t10 VSUBS 0.308984f
C873 VTAIL.n0 VSUBS 2.39044f
C874 VTAIL.n1 VSUBS 0.692602f
C875 VTAIL.n2 VSUBS 0.024181f
C876 VTAIL.n3 VSUBS 0.023357f
C877 VTAIL.n4 VSUBS 0.012551f
C878 VTAIL.n5 VSUBS 0.029667f
C879 VTAIL.n6 VSUBS 0.01329f
C880 VTAIL.n7 VSUBS 0.023357f
C881 VTAIL.n8 VSUBS 0.012551f
C882 VTAIL.n9 VSUBS 0.029667f
C883 VTAIL.n10 VSUBS 0.01329f
C884 VTAIL.n11 VSUBS 0.023357f
C885 VTAIL.n12 VSUBS 0.012551f
C886 VTAIL.n13 VSUBS 0.029667f
C887 VTAIL.n14 VSUBS 0.01329f
C888 VTAIL.n15 VSUBS 0.023357f
C889 VTAIL.n16 VSUBS 0.012551f
C890 VTAIL.n17 VSUBS 0.029667f
C891 VTAIL.n18 VSUBS 0.01329f
C892 VTAIL.n19 VSUBS 0.023357f
C893 VTAIL.n20 VSUBS 0.012551f
C894 VTAIL.n21 VSUBS 0.029667f
C895 VTAIL.n22 VSUBS 0.01329f
C896 VTAIL.n23 VSUBS 0.023357f
C897 VTAIL.n24 VSUBS 0.012551f
C898 VTAIL.n25 VSUBS 0.029667f
C899 VTAIL.n26 VSUBS 0.01329f
C900 VTAIL.n27 VSUBS 0.023357f
C901 VTAIL.n28 VSUBS 0.012551f
C902 VTAIL.n29 VSUBS 0.029667f
C903 VTAIL.n30 VSUBS 0.01329f
C904 VTAIL.n31 VSUBS 0.176638f
C905 VTAIL.t13 VSUBS 0.063611f
C906 VTAIL.n32 VSUBS 0.02225f
C907 VTAIL.n33 VSUBS 0.018873f
C908 VTAIL.n34 VSUBS 0.012551f
C909 VTAIL.n35 VSUBS 1.67593f
C910 VTAIL.n36 VSUBS 0.023357f
C911 VTAIL.n37 VSUBS 0.012551f
C912 VTAIL.n38 VSUBS 0.01329f
C913 VTAIL.n39 VSUBS 0.029667f
C914 VTAIL.n40 VSUBS 0.029667f
C915 VTAIL.n41 VSUBS 0.01329f
C916 VTAIL.n42 VSUBS 0.012551f
C917 VTAIL.n43 VSUBS 0.023357f
C918 VTAIL.n44 VSUBS 0.023357f
C919 VTAIL.n45 VSUBS 0.012551f
C920 VTAIL.n46 VSUBS 0.01329f
C921 VTAIL.n47 VSUBS 0.029667f
C922 VTAIL.n48 VSUBS 0.029667f
C923 VTAIL.n49 VSUBS 0.01329f
C924 VTAIL.n50 VSUBS 0.012551f
C925 VTAIL.n51 VSUBS 0.023357f
C926 VTAIL.n52 VSUBS 0.023357f
C927 VTAIL.n53 VSUBS 0.012551f
C928 VTAIL.n54 VSUBS 0.01329f
C929 VTAIL.n55 VSUBS 0.029667f
C930 VTAIL.n56 VSUBS 0.029667f
C931 VTAIL.n57 VSUBS 0.01329f
C932 VTAIL.n58 VSUBS 0.012551f
C933 VTAIL.n59 VSUBS 0.023357f
C934 VTAIL.n60 VSUBS 0.023357f
C935 VTAIL.n61 VSUBS 0.012551f
C936 VTAIL.n62 VSUBS 0.01329f
C937 VTAIL.n63 VSUBS 0.029667f
C938 VTAIL.n64 VSUBS 0.029667f
C939 VTAIL.n65 VSUBS 0.01329f
C940 VTAIL.n66 VSUBS 0.012551f
C941 VTAIL.n67 VSUBS 0.023357f
C942 VTAIL.n68 VSUBS 0.023357f
C943 VTAIL.n69 VSUBS 0.012551f
C944 VTAIL.n70 VSUBS 0.01329f
C945 VTAIL.n71 VSUBS 0.029667f
C946 VTAIL.n72 VSUBS 0.029667f
C947 VTAIL.n73 VSUBS 0.029667f
C948 VTAIL.n74 VSUBS 0.01329f
C949 VTAIL.n75 VSUBS 0.012551f
C950 VTAIL.n76 VSUBS 0.023357f
C951 VTAIL.n77 VSUBS 0.023357f
C952 VTAIL.n78 VSUBS 0.012551f
C953 VTAIL.n79 VSUBS 0.01292f
C954 VTAIL.n80 VSUBS 0.01292f
C955 VTAIL.n81 VSUBS 0.029667f
C956 VTAIL.n82 VSUBS 0.029667f
C957 VTAIL.n83 VSUBS 0.01329f
C958 VTAIL.n84 VSUBS 0.012551f
C959 VTAIL.n85 VSUBS 0.023357f
C960 VTAIL.n86 VSUBS 0.023357f
C961 VTAIL.n87 VSUBS 0.012551f
C962 VTAIL.n88 VSUBS 0.01329f
C963 VTAIL.n89 VSUBS 0.029667f
C964 VTAIL.n90 VSUBS 0.066766f
C965 VTAIL.n91 VSUBS 0.01329f
C966 VTAIL.n92 VSUBS 0.012551f
C967 VTAIL.n93 VSUBS 0.052075f
C968 VTAIL.n94 VSUBS 0.033292f
C969 VTAIL.n95 VSUBS 0.165178f
C970 VTAIL.n96 VSUBS 0.024181f
C971 VTAIL.n97 VSUBS 0.023357f
C972 VTAIL.n98 VSUBS 0.012551f
C973 VTAIL.n99 VSUBS 0.029667f
C974 VTAIL.n100 VSUBS 0.01329f
C975 VTAIL.n101 VSUBS 0.023357f
C976 VTAIL.n102 VSUBS 0.012551f
C977 VTAIL.n103 VSUBS 0.029667f
C978 VTAIL.n104 VSUBS 0.01329f
C979 VTAIL.n105 VSUBS 0.023357f
C980 VTAIL.n106 VSUBS 0.012551f
C981 VTAIL.n107 VSUBS 0.029667f
C982 VTAIL.n108 VSUBS 0.01329f
C983 VTAIL.n109 VSUBS 0.023357f
C984 VTAIL.n110 VSUBS 0.012551f
C985 VTAIL.n111 VSUBS 0.029667f
C986 VTAIL.n112 VSUBS 0.01329f
C987 VTAIL.n113 VSUBS 0.023357f
C988 VTAIL.n114 VSUBS 0.012551f
C989 VTAIL.n115 VSUBS 0.029667f
C990 VTAIL.n116 VSUBS 0.01329f
C991 VTAIL.n117 VSUBS 0.023357f
C992 VTAIL.n118 VSUBS 0.012551f
C993 VTAIL.n119 VSUBS 0.029667f
C994 VTAIL.n120 VSUBS 0.01329f
C995 VTAIL.n121 VSUBS 0.023357f
C996 VTAIL.n122 VSUBS 0.012551f
C997 VTAIL.n123 VSUBS 0.029667f
C998 VTAIL.n124 VSUBS 0.01329f
C999 VTAIL.n125 VSUBS 0.176638f
C1000 VTAIL.t1 VSUBS 0.063611f
C1001 VTAIL.n126 VSUBS 0.02225f
C1002 VTAIL.n127 VSUBS 0.018873f
C1003 VTAIL.n128 VSUBS 0.012551f
C1004 VTAIL.n129 VSUBS 1.67593f
C1005 VTAIL.n130 VSUBS 0.023357f
C1006 VTAIL.n131 VSUBS 0.012551f
C1007 VTAIL.n132 VSUBS 0.01329f
C1008 VTAIL.n133 VSUBS 0.029667f
C1009 VTAIL.n134 VSUBS 0.029667f
C1010 VTAIL.n135 VSUBS 0.01329f
C1011 VTAIL.n136 VSUBS 0.012551f
C1012 VTAIL.n137 VSUBS 0.023357f
C1013 VTAIL.n138 VSUBS 0.023357f
C1014 VTAIL.n139 VSUBS 0.012551f
C1015 VTAIL.n140 VSUBS 0.01329f
C1016 VTAIL.n141 VSUBS 0.029667f
C1017 VTAIL.n142 VSUBS 0.029667f
C1018 VTAIL.n143 VSUBS 0.01329f
C1019 VTAIL.n144 VSUBS 0.012551f
C1020 VTAIL.n145 VSUBS 0.023357f
C1021 VTAIL.n146 VSUBS 0.023357f
C1022 VTAIL.n147 VSUBS 0.012551f
C1023 VTAIL.n148 VSUBS 0.01329f
C1024 VTAIL.n149 VSUBS 0.029667f
C1025 VTAIL.n150 VSUBS 0.029667f
C1026 VTAIL.n151 VSUBS 0.01329f
C1027 VTAIL.n152 VSUBS 0.012551f
C1028 VTAIL.n153 VSUBS 0.023357f
C1029 VTAIL.n154 VSUBS 0.023357f
C1030 VTAIL.n155 VSUBS 0.012551f
C1031 VTAIL.n156 VSUBS 0.01329f
C1032 VTAIL.n157 VSUBS 0.029667f
C1033 VTAIL.n158 VSUBS 0.029667f
C1034 VTAIL.n159 VSUBS 0.01329f
C1035 VTAIL.n160 VSUBS 0.012551f
C1036 VTAIL.n161 VSUBS 0.023357f
C1037 VTAIL.n162 VSUBS 0.023357f
C1038 VTAIL.n163 VSUBS 0.012551f
C1039 VTAIL.n164 VSUBS 0.01329f
C1040 VTAIL.n165 VSUBS 0.029667f
C1041 VTAIL.n166 VSUBS 0.029667f
C1042 VTAIL.n167 VSUBS 0.029667f
C1043 VTAIL.n168 VSUBS 0.01329f
C1044 VTAIL.n169 VSUBS 0.012551f
C1045 VTAIL.n170 VSUBS 0.023357f
C1046 VTAIL.n171 VSUBS 0.023357f
C1047 VTAIL.n172 VSUBS 0.012551f
C1048 VTAIL.n173 VSUBS 0.01292f
C1049 VTAIL.n174 VSUBS 0.01292f
C1050 VTAIL.n175 VSUBS 0.029667f
C1051 VTAIL.n176 VSUBS 0.029667f
C1052 VTAIL.n177 VSUBS 0.01329f
C1053 VTAIL.n178 VSUBS 0.012551f
C1054 VTAIL.n179 VSUBS 0.023357f
C1055 VTAIL.n180 VSUBS 0.023357f
C1056 VTAIL.n181 VSUBS 0.012551f
C1057 VTAIL.n182 VSUBS 0.01329f
C1058 VTAIL.n183 VSUBS 0.029667f
C1059 VTAIL.n184 VSUBS 0.066766f
C1060 VTAIL.n185 VSUBS 0.01329f
C1061 VTAIL.n186 VSUBS 0.012551f
C1062 VTAIL.n187 VSUBS 0.052075f
C1063 VTAIL.n188 VSUBS 0.033292f
C1064 VTAIL.n189 VSUBS 0.165178f
C1065 VTAIL.t2 VSUBS 0.308984f
C1066 VTAIL.t4 VSUBS 0.308984f
C1067 VTAIL.n190 VSUBS 2.39044f
C1068 VTAIL.n191 VSUBS 0.799171f
C1069 VTAIL.n192 VSUBS 0.024181f
C1070 VTAIL.n193 VSUBS 0.023357f
C1071 VTAIL.n194 VSUBS 0.012551f
C1072 VTAIL.n195 VSUBS 0.029667f
C1073 VTAIL.n196 VSUBS 0.01329f
C1074 VTAIL.n197 VSUBS 0.023357f
C1075 VTAIL.n198 VSUBS 0.012551f
C1076 VTAIL.n199 VSUBS 0.029667f
C1077 VTAIL.n200 VSUBS 0.01329f
C1078 VTAIL.n201 VSUBS 0.023357f
C1079 VTAIL.n202 VSUBS 0.012551f
C1080 VTAIL.n203 VSUBS 0.029667f
C1081 VTAIL.n204 VSUBS 0.01329f
C1082 VTAIL.n205 VSUBS 0.023357f
C1083 VTAIL.n206 VSUBS 0.012551f
C1084 VTAIL.n207 VSUBS 0.029667f
C1085 VTAIL.n208 VSUBS 0.01329f
C1086 VTAIL.n209 VSUBS 0.023357f
C1087 VTAIL.n210 VSUBS 0.012551f
C1088 VTAIL.n211 VSUBS 0.029667f
C1089 VTAIL.n212 VSUBS 0.01329f
C1090 VTAIL.n213 VSUBS 0.023357f
C1091 VTAIL.n214 VSUBS 0.012551f
C1092 VTAIL.n215 VSUBS 0.029667f
C1093 VTAIL.n216 VSUBS 0.01329f
C1094 VTAIL.n217 VSUBS 0.023357f
C1095 VTAIL.n218 VSUBS 0.012551f
C1096 VTAIL.n219 VSUBS 0.029667f
C1097 VTAIL.n220 VSUBS 0.01329f
C1098 VTAIL.n221 VSUBS 0.176638f
C1099 VTAIL.t5 VSUBS 0.063611f
C1100 VTAIL.n222 VSUBS 0.02225f
C1101 VTAIL.n223 VSUBS 0.018873f
C1102 VTAIL.n224 VSUBS 0.012551f
C1103 VTAIL.n225 VSUBS 1.67593f
C1104 VTAIL.n226 VSUBS 0.023357f
C1105 VTAIL.n227 VSUBS 0.012551f
C1106 VTAIL.n228 VSUBS 0.01329f
C1107 VTAIL.n229 VSUBS 0.029667f
C1108 VTAIL.n230 VSUBS 0.029667f
C1109 VTAIL.n231 VSUBS 0.01329f
C1110 VTAIL.n232 VSUBS 0.012551f
C1111 VTAIL.n233 VSUBS 0.023357f
C1112 VTAIL.n234 VSUBS 0.023357f
C1113 VTAIL.n235 VSUBS 0.012551f
C1114 VTAIL.n236 VSUBS 0.01329f
C1115 VTAIL.n237 VSUBS 0.029667f
C1116 VTAIL.n238 VSUBS 0.029667f
C1117 VTAIL.n239 VSUBS 0.01329f
C1118 VTAIL.n240 VSUBS 0.012551f
C1119 VTAIL.n241 VSUBS 0.023357f
C1120 VTAIL.n242 VSUBS 0.023357f
C1121 VTAIL.n243 VSUBS 0.012551f
C1122 VTAIL.n244 VSUBS 0.01329f
C1123 VTAIL.n245 VSUBS 0.029667f
C1124 VTAIL.n246 VSUBS 0.029667f
C1125 VTAIL.n247 VSUBS 0.01329f
C1126 VTAIL.n248 VSUBS 0.012551f
C1127 VTAIL.n249 VSUBS 0.023357f
C1128 VTAIL.n250 VSUBS 0.023357f
C1129 VTAIL.n251 VSUBS 0.012551f
C1130 VTAIL.n252 VSUBS 0.01329f
C1131 VTAIL.n253 VSUBS 0.029667f
C1132 VTAIL.n254 VSUBS 0.029667f
C1133 VTAIL.n255 VSUBS 0.01329f
C1134 VTAIL.n256 VSUBS 0.012551f
C1135 VTAIL.n257 VSUBS 0.023357f
C1136 VTAIL.n258 VSUBS 0.023357f
C1137 VTAIL.n259 VSUBS 0.012551f
C1138 VTAIL.n260 VSUBS 0.01329f
C1139 VTAIL.n261 VSUBS 0.029667f
C1140 VTAIL.n262 VSUBS 0.029667f
C1141 VTAIL.n263 VSUBS 0.029667f
C1142 VTAIL.n264 VSUBS 0.01329f
C1143 VTAIL.n265 VSUBS 0.012551f
C1144 VTAIL.n266 VSUBS 0.023357f
C1145 VTAIL.n267 VSUBS 0.023357f
C1146 VTAIL.n268 VSUBS 0.012551f
C1147 VTAIL.n269 VSUBS 0.01292f
C1148 VTAIL.n270 VSUBS 0.01292f
C1149 VTAIL.n271 VSUBS 0.029667f
C1150 VTAIL.n272 VSUBS 0.029667f
C1151 VTAIL.n273 VSUBS 0.01329f
C1152 VTAIL.n274 VSUBS 0.012551f
C1153 VTAIL.n275 VSUBS 0.023357f
C1154 VTAIL.n276 VSUBS 0.023357f
C1155 VTAIL.n277 VSUBS 0.012551f
C1156 VTAIL.n278 VSUBS 0.01329f
C1157 VTAIL.n279 VSUBS 0.029667f
C1158 VTAIL.n280 VSUBS 0.066766f
C1159 VTAIL.n281 VSUBS 0.01329f
C1160 VTAIL.n282 VSUBS 0.012551f
C1161 VTAIL.n283 VSUBS 0.052075f
C1162 VTAIL.n284 VSUBS 0.033292f
C1163 VTAIL.n285 VSUBS 1.64418f
C1164 VTAIL.n286 VSUBS 0.024181f
C1165 VTAIL.n287 VSUBS 0.023357f
C1166 VTAIL.n288 VSUBS 0.012551f
C1167 VTAIL.n289 VSUBS 0.029667f
C1168 VTAIL.n290 VSUBS 0.01329f
C1169 VTAIL.n291 VSUBS 0.023357f
C1170 VTAIL.n292 VSUBS 0.012551f
C1171 VTAIL.n293 VSUBS 0.029667f
C1172 VTAIL.n294 VSUBS 0.01329f
C1173 VTAIL.n295 VSUBS 0.023357f
C1174 VTAIL.n296 VSUBS 0.012551f
C1175 VTAIL.n297 VSUBS 0.029667f
C1176 VTAIL.n298 VSUBS 0.029667f
C1177 VTAIL.n299 VSUBS 0.01329f
C1178 VTAIL.n300 VSUBS 0.023357f
C1179 VTAIL.n301 VSUBS 0.012551f
C1180 VTAIL.n302 VSUBS 0.029667f
C1181 VTAIL.n303 VSUBS 0.01329f
C1182 VTAIL.n304 VSUBS 0.023357f
C1183 VTAIL.n305 VSUBS 0.012551f
C1184 VTAIL.n306 VSUBS 0.029667f
C1185 VTAIL.n307 VSUBS 0.01329f
C1186 VTAIL.n308 VSUBS 0.023357f
C1187 VTAIL.n309 VSUBS 0.012551f
C1188 VTAIL.n310 VSUBS 0.029667f
C1189 VTAIL.n311 VSUBS 0.01329f
C1190 VTAIL.n312 VSUBS 0.023357f
C1191 VTAIL.n313 VSUBS 0.012551f
C1192 VTAIL.n314 VSUBS 0.029667f
C1193 VTAIL.n315 VSUBS 0.01329f
C1194 VTAIL.n316 VSUBS 0.176638f
C1195 VTAIL.t15 VSUBS 0.063611f
C1196 VTAIL.n317 VSUBS 0.02225f
C1197 VTAIL.n318 VSUBS 0.018873f
C1198 VTAIL.n319 VSUBS 0.012551f
C1199 VTAIL.n320 VSUBS 1.67593f
C1200 VTAIL.n321 VSUBS 0.023357f
C1201 VTAIL.n322 VSUBS 0.012551f
C1202 VTAIL.n323 VSUBS 0.01329f
C1203 VTAIL.n324 VSUBS 0.029667f
C1204 VTAIL.n325 VSUBS 0.029667f
C1205 VTAIL.n326 VSUBS 0.01329f
C1206 VTAIL.n327 VSUBS 0.012551f
C1207 VTAIL.n328 VSUBS 0.023357f
C1208 VTAIL.n329 VSUBS 0.023357f
C1209 VTAIL.n330 VSUBS 0.012551f
C1210 VTAIL.n331 VSUBS 0.01329f
C1211 VTAIL.n332 VSUBS 0.029667f
C1212 VTAIL.n333 VSUBS 0.029667f
C1213 VTAIL.n334 VSUBS 0.01329f
C1214 VTAIL.n335 VSUBS 0.012551f
C1215 VTAIL.n336 VSUBS 0.023357f
C1216 VTAIL.n337 VSUBS 0.023357f
C1217 VTAIL.n338 VSUBS 0.012551f
C1218 VTAIL.n339 VSUBS 0.01329f
C1219 VTAIL.n340 VSUBS 0.029667f
C1220 VTAIL.n341 VSUBS 0.029667f
C1221 VTAIL.n342 VSUBS 0.01329f
C1222 VTAIL.n343 VSUBS 0.012551f
C1223 VTAIL.n344 VSUBS 0.023357f
C1224 VTAIL.n345 VSUBS 0.023357f
C1225 VTAIL.n346 VSUBS 0.012551f
C1226 VTAIL.n347 VSUBS 0.01329f
C1227 VTAIL.n348 VSUBS 0.029667f
C1228 VTAIL.n349 VSUBS 0.029667f
C1229 VTAIL.n350 VSUBS 0.01329f
C1230 VTAIL.n351 VSUBS 0.012551f
C1231 VTAIL.n352 VSUBS 0.023357f
C1232 VTAIL.n353 VSUBS 0.023357f
C1233 VTAIL.n354 VSUBS 0.012551f
C1234 VTAIL.n355 VSUBS 0.01329f
C1235 VTAIL.n356 VSUBS 0.029667f
C1236 VTAIL.n357 VSUBS 0.029667f
C1237 VTAIL.n358 VSUBS 0.01329f
C1238 VTAIL.n359 VSUBS 0.012551f
C1239 VTAIL.n360 VSUBS 0.023357f
C1240 VTAIL.n361 VSUBS 0.023357f
C1241 VTAIL.n362 VSUBS 0.012551f
C1242 VTAIL.n363 VSUBS 0.01292f
C1243 VTAIL.n364 VSUBS 0.01292f
C1244 VTAIL.n365 VSUBS 0.029667f
C1245 VTAIL.n366 VSUBS 0.029667f
C1246 VTAIL.n367 VSUBS 0.01329f
C1247 VTAIL.n368 VSUBS 0.012551f
C1248 VTAIL.n369 VSUBS 0.023357f
C1249 VTAIL.n370 VSUBS 0.023357f
C1250 VTAIL.n371 VSUBS 0.012551f
C1251 VTAIL.n372 VSUBS 0.01329f
C1252 VTAIL.n373 VSUBS 0.029667f
C1253 VTAIL.n374 VSUBS 0.066766f
C1254 VTAIL.n375 VSUBS 0.01329f
C1255 VTAIL.n376 VSUBS 0.012551f
C1256 VTAIL.n377 VSUBS 0.052075f
C1257 VTAIL.n378 VSUBS 0.033292f
C1258 VTAIL.n379 VSUBS 1.64418f
C1259 VTAIL.t12 VSUBS 0.308984f
C1260 VTAIL.t9 VSUBS 0.308984f
C1261 VTAIL.n380 VSUBS 2.39046f
C1262 VTAIL.n381 VSUBS 0.799155f
C1263 VTAIL.n382 VSUBS 0.024181f
C1264 VTAIL.n383 VSUBS 0.023357f
C1265 VTAIL.n384 VSUBS 0.012551f
C1266 VTAIL.n385 VSUBS 0.029667f
C1267 VTAIL.n386 VSUBS 0.01329f
C1268 VTAIL.n387 VSUBS 0.023357f
C1269 VTAIL.n388 VSUBS 0.012551f
C1270 VTAIL.n389 VSUBS 0.029667f
C1271 VTAIL.n390 VSUBS 0.01329f
C1272 VTAIL.n391 VSUBS 0.023357f
C1273 VTAIL.n392 VSUBS 0.012551f
C1274 VTAIL.n393 VSUBS 0.029667f
C1275 VTAIL.n394 VSUBS 0.029667f
C1276 VTAIL.n395 VSUBS 0.01329f
C1277 VTAIL.n396 VSUBS 0.023357f
C1278 VTAIL.n397 VSUBS 0.012551f
C1279 VTAIL.n398 VSUBS 0.029667f
C1280 VTAIL.n399 VSUBS 0.01329f
C1281 VTAIL.n400 VSUBS 0.023357f
C1282 VTAIL.n401 VSUBS 0.012551f
C1283 VTAIL.n402 VSUBS 0.029667f
C1284 VTAIL.n403 VSUBS 0.01329f
C1285 VTAIL.n404 VSUBS 0.023357f
C1286 VTAIL.n405 VSUBS 0.012551f
C1287 VTAIL.n406 VSUBS 0.029667f
C1288 VTAIL.n407 VSUBS 0.01329f
C1289 VTAIL.n408 VSUBS 0.023357f
C1290 VTAIL.n409 VSUBS 0.012551f
C1291 VTAIL.n410 VSUBS 0.029667f
C1292 VTAIL.n411 VSUBS 0.01329f
C1293 VTAIL.n412 VSUBS 0.176638f
C1294 VTAIL.t14 VSUBS 0.063611f
C1295 VTAIL.n413 VSUBS 0.02225f
C1296 VTAIL.n414 VSUBS 0.018873f
C1297 VTAIL.n415 VSUBS 0.012551f
C1298 VTAIL.n416 VSUBS 1.67593f
C1299 VTAIL.n417 VSUBS 0.023357f
C1300 VTAIL.n418 VSUBS 0.012551f
C1301 VTAIL.n419 VSUBS 0.01329f
C1302 VTAIL.n420 VSUBS 0.029667f
C1303 VTAIL.n421 VSUBS 0.029667f
C1304 VTAIL.n422 VSUBS 0.01329f
C1305 VTAIL.n423 VSUBS 0.012551f
C1306 VTAIL.n424 VSUBS 0.023357f
C1307 VTAIL.n425 VSUBS 0.023357f
C1308 VTAIL.n426 VSUBS 0.012551f
C1309 VTAIL.n427 VSUBS 0.01329f
C1310 VTAIL.n428 VSUBS 0.029667f
C1311 VTAIL.n429 VSUBS 0.029667f
C1312 VTAIL.n430 VSUBS 0.01329f
C1313 VTAIL.n431 VSUBS 0.012551f
C1314 VTAIL.n432 VSUBS 0.023357f
C1315 VTAIL.n433 VSUBS 0.023357f
C1316 VTAIL.n434 VSUBS 0.012551f
C1317 VTAIL.n435 VSUBS 0.01329f
C1318 VTAIL.n436 VSUBS 0.029667f
C1319 VTAIL.n437 VSUBS 0.029667f
C1320 VTAIL.n438 VSUBS 0.01329f
C1321 VTAIL.n439 VSUBS 0.012551f
C1322 VTAIL.n440 VSUBS 0.023357f
C1323 VTAIL.n441 VSUBS 0.023357f
C1324 VTAIL.n442 VSUBS 0.012551f
C1325 VTAIL.n443 VSUBS 0.01329f
C1326 VTAIL.n444 VSUBS 0.029667f
C1327 VTAIL.n445 VSUBS 0.029667f
C1328 VTAIL.n446 VSUBS 0.01329f
C1329 VTAIL.n447 VSUBS 0.012551f
C1330 VTAIL.n448 VSUBS 0.023357f
C1331 VTAIL.n449 VSUBS 0.023357f
C1332 VTAIL.n450 VSUBS 0.012551f
C1333 VTAIL.n451 VSUBS 0.01329f
C1334 VTAIL.n452 VSUBS 0.029667f
C1335 VTAIL.n453 VSUBS 0.029667f
C1336 VTAIL.n454 VSUBS 0.01329f
C1337 VTAIL.n455 VSUBS 0.012551f
C1338 VTAIL.n456 VSUBS 0.023357f
C1339 VTAIL.n457 VSUBS 0.023357f
C1340 VTAIL.n458 VSUBS 0.012551f
C1341 VTAIL.n459 VSUBS 0.01292f
C1342 VTAIL.n460 VSUBS 0.01292f
C1343 VTAIL.n461 VSUBS 0.029667f
C1344 VTAIL.n462 VSUBS 0.029667f
C1345 VTAIL.n463 VSUBS 0.01329f
C1346 VTAIL.n464 VSUBS 0.012551f
C1347 VTAIL.n465 VSUBS 0.023357f
C1348 VTAIL.n466 VSUBS 0.023357f
C1349 VTAIL.n467 VSUBS 0.012551f
C1350 VTAIL.n468 VSUBS 0.01329f
C1351 VTAIL.n469 VSUBS 0.029667f
C1352 VTAIL.n470 VSUBS 0.066766f
C1353 VTAIL.n471 VSUBS 0.01329f
C1354 VTAIL.n472 VSUBS 0.012551f
C1355 VTAIL.n473 VSUBS 0.052075f
C1356 VTAIL.n474 VSUBS 0.033292f
C1357 VTAIL.n475 VSUBS 0.165178f
C1358 VTAIL.n476 VSUBS 0.024181f
C1359 VTAIL.n477 VSUBS 0.023357f
C1360 VTAIL.n478 VSUBS 0.012551f
C1361 VTAIL.n479 VSUBS 0.029667f
C1362 VTAIL.n480 VSUBS 0.01329f
C1363 VTAIL.n481 VSUBS 0.023357f
C1364 VTAIL.n482 VSUBS 0.012551f
C1365 VTAIL.n483 VSUBS 0.029667f
C1366 VTAIL.n484 VSUBS 0.01329f
C1367 VTAIL.n485 VSUBS 0.023357f
C1368 VTAIL.n486 VSUBS 0.012551f
C1369 VTAIL.n487 VSUBS 0.029667f
C1370 VTAIL.n488 VSUBS 0.029667f
C1371 VTAIL.n489 VSUBS 0.01329f
C1372 VTAIL.n490 VSUBS 0.023357f
C1373 VTAIL.n491 VSUBS 0.012551f
C1374 VTAIL.n492 VSUBS 0.029667f
C1375 VTAIL.n493 VSUBS 0.01329f
C1376 VTAIL.n494 VSUBS 0.023357f
C1377 VTAIL.n495 VSUBS 0.012551f
C1378 VTAIL.n496 VSUBS 0.029667f
C1379 VTAIL.n497 VSUBS 0.01329f
C1380 VTAIL.n498 VSUBS 0.023357f
C1381 VTAIL.n499 VSUBS 0.012551f
C1382 VTAIL.n500 VSUBS 0.029667f
C1383 VTAIL.n501 VSUBS 0.01329f
C1384 VTAIL.n502 VSUBS 0.023357f
C1385 VTAIL.n503 VSUBS 0.012551f
C1386 VTAIL.n504 VSUBS 0.029667f
C1387 VTAIL.n505 VSUBS 0.01329f
C1388 VTAIL.n506 VSUBS 0.176638f
C1389 VTAIL.t7 VSUBS 0.063611f
C1390 VTAIL.n507 VSUBS 0.02225f
C1391 VTAIL.n508 VSUBS 0.018873f
C1392 VTAIL.n509 VSUBS 0.012551f
C1393 VTAIL.n510 VSUBS 1.67593f
C1394 VTAIL.n511 VSUBS 0.023357f
C1395 VTAIL.n512 VSUBS 0.012551f
C1396 VTAIL.n513 VSUBS 0.01329f
C1397 VTAIL.n514 VSUBS 0.029667f
C1398 VTAIL.n515 VSUBS 0.029667f
C1399 VTAIL.n516 VSUBS 0.01329f
C1400 VTAIL.n517 VSUBS 0.012551f
C1401 VTAIL.n518 VSUBS 0.023357f
C1402 VTAIL.n519 VSUBS 0.023357f
C1403 VTAIL.n520 VSUBS 0.012551f
C1404 VTAIL.n521 VSUBS 0.01329f
C1405 VTAIL.n522 VSUBS 0.029667f
C1406 VTAIL.n523 VSUBS 0.029667f
C1407 VTAIL.n524 VSUBS 0.01329f
C1408 VTAIL.n525 VSUBS 0.012551f
C1409 VTAIL.n526 VSUBS 0.023357f
C1410 VTAIL.n527 VSUBS 0.023357f
C1411 VTAIL.n528 VSUBS 0.012551f
C1412 VTAIL.n529 VSUBS 0.01329f
C1413 VTAIL.n530 VSUBS 0.029667f
C1414 VTAIL.n531 VSUBS 0.029667f
C1415 VTAIL.n532 VSUBS 0.01329f
C1416 VTAIL.n533 VSUBS 0.012551f
C1417 VTAIL.n534 VSUBS 0.023357f
C1418 VTAIL.n535 VSUBS 0.023357f
C1419 VTAIL.n536 VSUBS 0.012551f
C1420 VTAIL.n537 VSUBS 0.01329f
C1421 VTAIL.n538 VSUBS 0.029667f
C1422 VTAIL.n539 VSUBS 0.029667f
C1423 VTAIL.n540 VSUBS 0.01329f
C1424 VTAIL.n541 VSUBS 0.012551f
C1425 VTAIL.n542 VSUBS 0.023357f
C1426 VTAIL.n543 VSUBS 0.023357f
C1427 VTAIL.n544 VSUBS 0.012551f
C1428 VTAIL.n545 VSUBS 0.01329f
C1429 VTAIL.n546 VSUBS 0.029667f
C1430 VTAIL.n547 VSUBS 0.029667f
C1431 VTAIL.n548 VSUBS 0.01329f
C1432 VTAIL.n549 VSUBS 0.012551f
C1433 VTAIL.n550 VSUBS 0.023357f
C1434 VTAIL.n551 VSUBS 0.023357f
C1435 VTAIL.n552 VSUBS 0.012551f
C1436 VTAIL.n553 VSUBS 0.01292f
C1437 VTAIL.n554 VSUBS 0.01292f
C1438 VTAIL.n555 VSUBS 0.029667f
C1439 VTAIL.n556 VSUBS 0.029667f
C1440 VTAIL.n557 VSUBS 0.01329f
C1441 VTAIL.n558 VSUBS 0.012551f
C1442 VTAIL.n559 VSUBS 0.023357f
C1443 VTAIL.n560 VSUBS 0.023357f
C1444 VTAIL.n561 VSUBS 0.012551f
C1445 VTAIL.n562 VSUBS 0.01329f
C1446 VTAIL.n563 VSUBS 0.029667f
C1447 VTAIL.n564 VSUBS 0.066766f
C1448 VTAIL.n565 VSUBS 0.01329f
C1449 VTAIL.n566 VSUBS 0.012551f
C1450 VTAIL.n567 VSUBS 0.052075f
C1451 VTAIL.n568 VSUBS 0.033292f
C1452 VTAIL.n569 VSUBS 0.165178f
C1453 VTAIL.t0 VSUBS 0.308984f
C1454 VTAIL.t3 VSUBS 0.308984f
C1455 VTAIL.n570 VSUBS 2.39046f
C1456 VTAIL.n571 VSUBS 0.799155f
C1457 VTAIL.n572 VSUBS 0.024181f
C1458 VTAIL.n573 VSUBS 0.023357f
C1459 VTAIL.n574 VSUBS 0.012551f
C1460 VTAIL.n575 VSUBS 0.029667f
C1461 VTAIL.n576 VSUBS 0.01329f
C1462 VTAIL.n577 VSUBS 0.023357f
C1463 VTAIL.n578 VSUBS 0.012551f
C1464 VTAIL.n579 VSUBS 0.029667f
C1465 VTAIL.n580 VSUBS 0.01329f
C1466 VTAIL.n581 VSUBS 0.023357f
C1467 VTAIL.n582 VSUBS 0.012551f
C1468 VTAIL.n583 VSUBS 0.029667f
C1469 VTAIL.n584 VSUBS 0.029667f
C1470 VTAIL.n585 VSUBS 0.01329f
C1471 VTAIL.n586 VSUBS 0.023357f
C1472 VTAIL.n587 VSUBS 0.012551f
C1473 VTAIL.n588 VSUBS 0.029667f
C1474 VTAIL.n589 VSUBS 0.01329f
C1475 VTAIL.n590 VSUBS 0.023357f
C1476 VTAIL.n591 VSUBS 0.012551f
C1477 VTAIL.n592 VSUBS 0.029667f
C1478 VTAIL.n593 VSUBS 0.01329f
C1479 VTAIL.n594 VSUBS 0.023357f
C1480 VTAIL.n595 VSUBS 0.012551f
C1481 VTAIL.n596 VSUBS 0.029667f
C1482 VTAIL.n597 VSUBS 0.01329f
C1483 VTAIL.n598 VSUBS 0.023357f
C1484 VTAIL.n599 VSUBS 0.012551f
C1485 VTAIL.n600 VSUBS 0.029667f
C1486 VTAIL.n601 VSUBS 0.01329f
C1487 VTAIL.n602 VSUBS 0.176638f
C1488 VTAIL.t6 VSUBS 0.063611f
C1489 VTAIL.n603 VSUBS 0.02225f
C1490 VTAIL.n604 VSUBS 0.018873f
C1491 VTAIL.n605 VSUBS 0.012551f
C1492 VTAIL.n606 VSUBS 1.67593f
C1493 VTAIL.n607 VSUBS 0.023357f
C1494 VTAIL.n608 VSUBS 0.012551f
C1495 VTAIL.n609 VSUBS 0.01329f
C1496 VTAIL.n610 VSUBS 0.029667f
C1497 VTAIL.n611 VSUBS 0.029667f
C1498 VTAIL.n612 VSUBS 0.01329f
C1499 VTAIL.n613 VSUBS 0.012551f
C1500 VTAIL.n614 VSUBS 0.023357f
C1501 VTAIL.n615 VSUBS 0.023357f
C1502 VTAIL.n616 VSUBS 0.012551f
C1503 VTAIL.n617 VSUBS 0.01329f
C1504 VTAIL.n618 VSUBS 0.029667f
C1505 VTAIL.n619 VSUBS 0.029667f
C1506 VTAIL.n620 VSUBS 0.01329f
C1507 VTAIL.n621 VSUBS 0.012551f
C1508 VTAIL.n622 VSUBS 0.023357f
C1509 VTAIL.n623 VSUBS 0.023357f
C1510 VTAIL.n624 VSUBS 0.012551f
C1511 VTAIL.n625 VSUBS 0.01329f
C1512 VTAIL.n626 VSUBS 0.029667f
C1513 VTAIL.n627 VSUBS 0.029667f
C1514 VTAIL.n628 VSUBS 0.01329f
C1515 VTAIL.n629 VSUBS 0.012551f
C1516 VTAIL.n630 VSUBS 0.023357f
C1517 VTAIL.n631 VSUBS 0.023357f
C1518 VTAIL.n632 VSUBS 0.012551f
C1519 VTAIL.n633 VSUBS 0.01329f
C1520 VTAIL.n634 VSUBS 0.029667f
C1521 VTAIL.n635 VSUBS 0.029667f
C1522 VTAIL.n636 VSUBS 0.01329f
C1523 VTAIL.n637 VSUBS 0.012551f
C1524 VTAIL.n638 VSUBS 0.023357f
C1525 VTAIL.n639 VSUBS 0.023357f
C1526 VTAIL.n640 VSUBS 0.012551f
C1527 VTAIL.n641 VSUBS 0.01329f
C1528 VTAIL.n642 VSUBS 0.029667f
C1529 VTAIL.n643 VSUBS 0.029667f
C1530 VTAIL.n644 VSUBS 0.01329f
C1531 VTAIL.n645 VSUBS 0.012551f
C1532 VTAIL.n646 VSUBS 0.023357f
C1533 VTAIL.n647 VSUBS 0.023357f
C1534 VTAIL.n648 VSUBS 0.012551f
C1535 VTAIL.n649 VSUBS 0.01292f
C1536 VTAIL.n650 VSUBS 0.01292f
C1537 VTAIL.n651 VSUBS 0.029667f
C1538 VTAIL.n652 VSUBS 0.029667f
C1539 VTAIL.n653 VSUBS 0.01329f
C1540 VTAIL.n654 VSUBS 0.012551f
C1541 VTAIL.n655 VSUBS 0.023357f
C1542 VTAIL.n656 VSUBS 0.023357f
C1543 VTAIL.n657 VSUBS 0.012551f
C1544 VTAIL.n658 VSUBS 0.01329f
C1545 VTAIL.n659 VSUBS 0.029667f
C1546 VTAIL.n660 VSUBS 0.066766f
C1547 VTAIL.n661 VSUBS 0.01329f
C1548 VTAIL.n662 VSUBS 0.012551f
C1549 VTAIL.n663 VSUBS 0.052075f
C1550 VTAIL.n664 VSUBS 0.033292f
C1551 VTAIL.n665 VSUBS 1.64418f
C1552 VTAIL.n666 VSUBS 0.024181f
C1553 VTAIL.n667 VSUBS 0.023357f
C1554 VTAIL.n668 VSUBS 0.012551f
C1555 VTAIL.n669 VSUBS 0.029667f
C1556 VTAIL.n670 VSUBS 0.01329f
C1557 VTAIL.n671 VSUBS 0.023357f
C1558 VTAIL.n672 VSUBS 0.012551f
C1559 VTAIL.n673 VSUBS 0.029667f
C1560 VTAIL.n674 VSUBS 0.01329f
C1561 VTAIL.n675 VSUBS 0.023357f
C1562 VTAIL.n676 VSUBS 0.012551f
C1563 VTAIL.n677 VSUBS 0.029667f
C1564 VTAIL.n678 VSUBS 0.01329f
C1565 VTAIL.n679 VSUBS 0.023357f
C1566 VTAIL.n680 VSUBS 0.012551f
C1567 VTAIL.n681 VSUBS 0.029667f
C1568 VTAIL.n682 VSUBS 0.01329f
C1569 VTAIL.n683 VSUBS 0.023357f
C1570 VTAIL.n684 VSUBS 0.012551f
C1571 VTAIL.n685 VSUBS 0.029667f
C1572 VTAIL.n686 VSUBS 0.01329f
C1573 VTAIL.n687 VSUBS 0.023357f
C1574 VTAIL.n688 VSUBS 0.012551f
C1575 VTAIL.n689 VSUBS 0.029667f
C1576 VTAIL.n690 VSUBS 0.01329f
C1577 VTAIL.n691 VSUBS 0.023357f
C1578 VTAIL.n692 VSUBS 0.012551f
C1579 VTAIL.n693 VSUBS 0.029667f
C1580 VTAIL.n694 VSUBS 0.01329f
C1581 VTAIL.n695 VSUBS 0.176638f
C1582 VTAIL.t8 VSUBS 0.063611f
C1583 VTAIL.n696 VSUBS 0.02225f
C1584 VTAIL.n697 VSUBS 0.018873f
C1585 VTAIL.n698 VSUBS 0.012551f
C1586 VTAIL.n699 VSUBS 1.67593f
C1587 VTAIL.n700 VSUBS 0.023357f
C1588 VTAIL.n701 VSUBS 0.012551f
C1589 VTAIL.n702 VSUBS 0.01329f
C1590 VTAIL.n703 VSUBS 0.029667f
C1591 VTAIL.n704 VSUBS 0.029667f
C1592 VTAIL.n705 VSUBS 0.01329f
C1593 VTAIL.n706 VSUBS 0.012551f
C1594 VTAIL.n707 VSUBS 0.023357f
C1595 VTAIL.n708 VSUBS 0.023357f
C1596 VTAIL.n709 VSUBS 0.012551f
C1597 VTAIL.n710 VSUBS 0.01329f
C1598 VTAIL.n711 VSUBS 0.029667f
C1599 VTAIL.n712 VSUBS 0.029667f
C1600 VTAIL.n713 VSUBS 0.01329f
C1601 VTAIL.n714 VSUBS 0.012551f
C1602 VTAIL.n715 VSUBS 0.023357f
C1603 VTAIL.n716 VSUBS 0.023357f
C1604 VTAIL.n717 VSUBS 0.012551f
C1605 VTAIL.n718 VSUBS 0.01329f
C1606 VTAIL.n719 VSUBS 0.029667f
C1607 VTAIL.n720 VSUBS 0.029667f
C1608 VTAIL.n721 VSUBS 0.01329f
C1609 VTAIL.n722 VSUBS 0.012551f
C1610 VTAIL.n723 VSUBS 0.023357f
C1611 VTAIL.n724 VSUBS 0.023357f
C1612 VTAIL.n725 VSUBS 0.012551f
C1613 VTAIL.n726 VSUBS 0.01329f
C1614 VTAIL.n727 VSUBS 0.029667f
C1615 VTAIL.n728 VSUBS 0.029667f
C1616 VTAIL.n729 VSUBS 0.01329f
C1617 VTAIL.n730 VSUBS 0.012551f
C1618 VTAIL.n731 VSUBS 0.023357f
C1619 VTAIL.n732 VSUBS 0.023357f
C1620 VTAIL.n733 VSUBS 0.012551f
C1621 VTAIL.n734 VSUBS 0.01329f
C1622 VTAIL.n735 VSUBS 0.029667f
C1623 VTAIL.n736 VSUBS 0.029667f
C1624 VTAIL.n737 VSUBS 0.029667f
C1625 VTAIL.n738 VSUBS 0.01329f
C1626 VTAIL.n739 VSUBS 0.012551f
C1627 VTAIL.n740 VSUBS 0.023357f
C1628 VTAIL.n741 VSUBS 0.023357f
C1629 VTAIL.n742 VSUBS 0.012551f
C1630 VTAIL.n743 VSUBS 0.01292f
C1631 VTAIL.n744 VSUBS 0.01292f
C1632 VTAIL.n745 VSUBS 0.029667f
C1633 VTAIL.n746 VSUBS 0.029667f
C1634 VTAIL.n747 VSUBS 0.01329f
C1635 VTAIL.n748 VSUBS 0.012551f
C1636 VTAIL.n749 VSUBS 0.023357f
C1637 VTAIL.n750 VSUBS 0.023357f
C1638 VTAIL.n751 VSUBS 0.012551f
C1639 VTAIL.n752 VSUBS 0.01329f
C1640 VTAIL.n753 VSUBS 0.029667f
C1641 VTAIL.n754 VSUBS 0.066766f
C1642 VTAIL.n755 VSUBS 0.01329f
C1643 VTAIL.n756 VSUBS 0.012551f
C1644 VTAIL.n757 VSUBS 0.052075f
C1645 VTAIL.n758 VSUBS 0.033292f
C1646 VTAIL.n759 VSUBS 1.6398f
C1647 VDD2.t5 VSUBS 0.333331f
C1648 VDD2.t7 VSUBS 0.333331f
C1649 VDD2.n0 VSUBS 2.745f
C1650 VDD2.t6 VSUBS 0.333331f
C1651 VDD2.t0 VSUBS 0.333331f
C1652 VDD2.n1 VSUBS 2.745f
C1653 VDD2.n2 VSUBS 3.46275f
C1654 VDD2.t3 VSUBS 0.333331f
C1655 VDD2.t4 VSUBS 0.333331f
C1656 VDD2.n3 VSUBS 2.73825f
C1657 VDD2.n4 VSUBS 3.2019f
C1658 VDD2.t1 VSUBS 0.333331f
C1659 VDD2.t2 VSUBS 0.333331f
C1660 VDD2.n5 VSUBS 2.74496f
C1661 VN.n0 VSUBS 0.037744f
C1662 VN.t7 VSUBS 2.39487f
C1663 VN.n1 VSUBS 0.065514f
C1664 VN.n2 VSUBS 0.037744f
C1665 VN.n3 VSUBS 0.042695f
C1666 VN.t2 VSUBS 2.48922f
C1667 VN.t4 VSUBS 2.39487f
C1668 VN.n4 VSUBS 0.90344f
C1669 VN.n5 VSUBS 0.941035f
C1670 VN.n6 VSUBS 0.203037f
C1671 VN.n7 VSUBS 0.037744f
C1672 VN.n8 VSUBS 0.054866f
C1673 VN.n9 VSUBS 0.054866f
C1674 VN.t5 VSUBS 2.39487f
C1675 VN.n10 VSUBS 0.849063f
C1676 VN.n11 VSUBS 0.042695f
C1677 VN.n12 VSUBS 0.037744f
C1678 VN.n13 VSUBS 0.037744f
C1679 VN.n14 VSUBS 0.037744f
C1680 VN.n15 VSUBS 0.031261f
C1681 VN.n16 VSUBS 0.062908f
C1682 VN.n17 VSUBS 0.928073f
C1683 VN.n18 VSUBS 0.033707f
C1684 VN.n19 VSUBS 0.037744f
C1685 VN.t0 VSUBS 2.39487f
C1686 VN.n20 VSUBS 0.065514f
C1687 VN.n21 VSUBS 0.037744f
C1688 VN.t3 VSUBS 2.39487f
C1689 VN.n22 VSUBS 0.849063f
C1690 VN.n23 VSUBS 0.042695f
C1691 VN.t1 VSUBS 2.48922f
C1692 VN.t6 VSUBS 2.39487f
C1693 VN.n24 VSUBS 0.90344f
C1694 VN.n25 VSUBS 0.941035f
C1695 VN.n26 VSUBS 0.203037f
C1696 VN.n27 VSUBS 0.037744f
C1697 VN.n28 VSUBS 0.054866f
C1698 VN.n29 VSUBS 0.054866f
C1699 VN.n30 VSUBS 0.042695f
C1700 VN.n31 VSUBS 0.037744f
C1701 VN.n32 VSUBS 0.037744f
C1702 VN.n33 VSUBS 0.037744f
C1703 VN.n34 VSUBS 0.031261f
C1704 VN.n35 VSUBS 0.062908f
C1705 VN.n36 VSUBS 0.928073f
C1706 VN.n37 VSUBS 2.00434f
.ends

