* NGSPICE file created from diff_pair_sample_0202.ext - technology: sky130A

.subckt diff_pair_sample_0202 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X1 VTAIL.t6 VN.t0 VDD2.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X2 VTAIL.t12 VP.t1 VDD1.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X3 VDD1.t7 VP.t2 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=7.3671 ps=38.56 w=18.89 l=3.79
X4 VTAIL.t13 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X5 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=0 ps=0 w=18.89 l=3.79
X6 VTAIL.t4 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X7 VDD2.t7 VN.t2 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X8 VDD1.t5 VP.t4 VTAIL.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X9 VTAIL.t5 VN.t3 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X10 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=7.3671 ps=38.56 w=18.89 l=3.79
X11 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=0 ps=0 w=18.89 l=3.79
X12 VTAIL.t11 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X13 VDD1.t3 VP.t6 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=3.11685 ps=19.22 w=18.89 l=3.79
X14 VDD1.t2 VP.t7 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=7.3671 ps=38.56 w=18.89 l=3.79
X15 VTAIL.t16 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X16 VDD1.t0 VP.t9 VTAIL.t19 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=3.11685 ps=19.22 w=18.89 l=3.79
X17 VDD2.t4 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=7.3671 ps=38.56 w=18.89 l=3.79
X18 VDD2.t3 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=3.11685 ps=19.22 w=18.89 l=3.79
X19 VDD2.t2 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=3.11685 ps=19.22 w=18.89 l=3.79
X20 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=0 ps=0 w=18.89 l=3.79
X21 VDD2.t1 VN.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3671 pd=38.56 as=0 ps=0 w=18.89 l=3.79
X23 VTAIL.t8 VN.t9 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=3.11685 pd=19.22 as=3.11685 ps=19.22 w=18.89 l=3.79
R0 VP.n31 VP.n30 161.3
R1 VP.n32 VP.n27 161.3
R2 VP.n34 VP.n33 161.3
R3 VP.n35 VP.n26 161.3
R4 VP.n37 VP.n36 161.3
R5 VP.n38 VP.n25 161.3
R6 VP.n40 VP.n39 161.3
R7 VP.n41 VP.n24 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n23 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n22 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n21 161.3
R14 VP.n53 VP.n52 161.3
R15 VP.n54 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n17 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n67 VP.n16 161.3
R24 VP.n122 VP.n0 161.3
R25 VP.n121 VP.n120 161.3
R26 VP.n119 VP.n1 161.3
R27 VP.n118 VP.n117 161.3
R28 VP.n116 VP.n2 161.3
R29 VP.n115 VP.n114 161.3
R30 VP.n113 VP.n3 161.3
R31 VP.n112 VP.n111 161.3
R32 VP.n109 VP.n4 161.3
R33 VP.n108 VP.n107 161.3
R34 VP.n106 VP.n5 161.3
R35 VP.n105 VP.n104 161.3
R36 VP.n103 VP.n6 161.3
R37 VP.n102 VP.n101 161.3
R38 VP.n100 VP.n7 161.3
R39 VP.n99 VP.n98 161.3
R40 VP.n96 VP.n8 161.3
R41 VP.n95 VP.n94 161.3
R42 VP.n93 VP.n9 161.3
R43 VP.n92 VP.n91 161.3
R44 VP.n90 VP.n10 161.3
R45 VP.n89 VP.n88 161.3
R46 VP.n87 VP.n11 161.3
R47 VP.n86 VP.n85 161.3
R48 VP.n83 VP.n12 161.3
R49 VP.n82 VP.n81 161.3
R50 VP.n80 VP.n13 161.3
R51 VP.n79 VP.n78 161.3
R52 VP.n77 VP.n14 161.3
R53 VP.n76 VP.n75 161.3
R54 VP.n74 VP.n15 161.3
R55 VP.n73 VP.n72 161.3
R56 VP.n28 VP.t6 152.219
R57 VP.n71 VP.t9 120.118
R58 VP.n84 VP.t1 120.118
R59 VP.n97 VP.t4 120.118
R60 VP.n110 VP.t3 120.118
R61 VP.n123 VP.t7 120.118
R62 VP.n68 VP.t2 120.118
R63 VP.n55 VP.t8 120.118
R64 VP.n42 VP.t0 120.118
R65 VP.n29 VP.t5 120.118
R66 VP.n70 VP.n69 65.057
R67 VP.n71 VP.n70 58.2041
R68 VP.n124 VP.n123 58.2041
R69 VP.n69 VP.n68 58.2041
R70 VP.n29 VP.n28 56.9469
R71 VP.n91 VP.n90 56.5193
R72 VP.n104 VP.n103 56.5193
R73 VP.n49 VP.n48 56.5193
R74 VP.n36 VP.n35 56.5193
R75 VP.n78 VP.n77 47.2923
R76 VP.n117 VP.n116 47.2923
R77 VP.n62 VP.n61 47.2923
R78 VP.n77 VP.n76 33.6945
R79 VP.n117 VP.n1 33.6945
R80 VP.n62 VP.n17 33.6945
R81 VP.n72 VP.n15 24.4675
R82 VP.n76 VP.n15 24.4675
R83 VP.n78 VP.n13 24.4675
R84 VP.n82 VP.n13 24.4675
R85 VP.n83 VP.n82 24.4675
R86 VP.n85 VP.n11 24.4675
R87 VP.n89 VP.n11 24.4675
R88 VP.n90 VP.n89 24.4675
R89 VP.n91 VP.n9 24.4675
R90 VP.n95 VP.n9 24.4675
R91 VP.n96 VP.n95 24.4675
R92 VP.n98 VP.n7 24.4675
R93 VP.n102 VP.n7 24.4675
R94 VP.n103 VP.n102 24.4675
R95 VP.n104 VP.n5 24.4675
R96 VP.n108 VP.n5 24.4675
R97 VP.n109 VP.n108 24.4675
R98 VP.n111 VP.n3 24.4675
R99 VP.n115 VP.n3 24.4675
R100 VP.n116 VP.n115 24.4675
R101 VP.n121 VP.n1 24.4675
R102 VP.n122 VP.n121 24.4675
R103 VP.n66 VP.n17 24.4675
R104 VP.n67 VP.n66 24.4675
R105 VP.n49 VP.n21 24.4675
R106 VP.n53 VP.n21 24.4675
R107 VP.n54 VP.n53 24.4675
R108 VP.n56 VP.n19 24.4675
R109 VP.n60 VP.n19 24.4675
R110 VP.n61 VP.n60 24.4675
R111 VP.n36 VP.n25 24.4675
R112 VP.n40 VP.n25 24.4675
R113 VP.n41 VP.n40 24.4675
R114 VP.n43 VP.n23 24.4675
R115 VP.n47 VP.n23 24.4675
R116 VP.n48 VP.n47 24.4675
R117 VP.n30 VP.n27 24.4675
R118 VP.n34 VP.n27 24.4675
R119 VP.n35 VP.n34 24.4675
R120 VP.n72 VP.n71 23.9782
R121 VP.n123 VP.n122 23.9782
R122 VP.n68 VP.n67 23.9782
R123 VP.n85 VP.n84 18.1061
R124 VP.n110 VP.n109 18.1061
R125 VP.n55 VP.n54 18.1061
R126 VP.n30 VP.n29 18.1061
R127 VP.n97 VP.n96 12.234
R128 VP.n98 VP.n97 12.234
R129 VP.n42 VP.n41 12.234
R130 VP.n43 VP.n42 12.234
R131 VP.n84 VP.n83 6.36192
R132 VP.n111 VP.n110 6.36192
R133 VP.n56 VP.n55 6.36192
R134 VP.n31 VP.n28 2.54561
R135 VP.n69 VP.n16 0.417535
R136 VP.n73 VP.n70 0.417535
R137 VP.n124 VP.n0 0.417535
R138 VP VP.n124 0.394291
R139 VP.n32 VP.n31 0.189894
R140 VP.n33 VP.n32 0.189894
R141 VP.n33 VP.n26 0.189894
R142 VP.n37 VP.n26 0.189894
R143 VP.n38 VP.n37 0.189894
R144 VP.n39 VP.n38 0.189894
R145 VP.n39 VP.n24 0.189894
R146 VP.n44 VP.n24 0.189894
R147 VP.n45 VP.n44 0.189894
R148 VP.n46 VP.n45 0.189894
R149 VP.n46 VP.n22 0.189894
R150 VP.n50 VP.n22 0.189894
R151 VP.n51 VP.n50 0.189894
R152 VP.n52 VP.n51 0.189894
R153 VP.n52 VP.n20 0.189894
R154 VP.n57 VP.n20 0.189894
R155 VP.n58 VP.n57 0.189894
R156 VP.n59 VP.n58 0.189894
R157 VP.n59 VP.n18 0.189894
R158 VP.n63 VP.n18 0.189894
R159 VP.n64 VP.n63 0.189894
R160 VP.n65 VP.n64 0.189894
R161 VP.n65 VP.n16 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n75 VP.n74 0.189894
R164 VP.n75 VP.n14 0.189894
R165 VP.n79 VP.n14 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n81 VP.n80 0.189894
R168 VP.n81 VP.n12 0.189894
R169 VP.n86 VP.n12 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n88 VP.n87 0.189894
R172 VP.n88 VP.n10 0.189894
R173 VP.n92 VP.n10 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n94 VP.n93 0.189894
R176 VP.n94 VP.n8 0.189894
R177 VP.n99 VP.n8 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n101 VP.n100 0.189894
R180 VP.n101 VP.n6 0.189894
R181 VP.n105 VP.n6 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n107 VP.n106 0.189894
R184 VP.n107 VP.n4 0.189894
R185 VP.n112 VP.n4 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n114 VP.n113 0.189894
R188 VP.n114 VP.n2 0.189894
R189 VP.n118 VP.n2 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n120 VP.n119 0.189894
R192 VP.n120 VP.n0 0.189894
R193 VTAIL.n432 VTAIL.n332 289.615
R194 VTAIL.n102 VTAIL.n2 289.615
R195 VTAIL.n326 VTAIL.n226 289.615
R196 VTAIL.n216 VTAIL.n116 289.615
R197 VTAIL.n367 VTAIL.n366 185
R198 VTAIL.n364 VTAIL.n363 185
R199 VTAIL.n373 VTAIL.n372 185
R200 VTAIL.n375 VTAIL.n374 185
R201 VTAIL.n360 VTAIL.n359 185
R202 VTAIL.n381 VTAIL.n380 185
R203 VTAIL.n383 VTAIL.n382 185
R204 VTAIL.n356 VTAIL.n355 185
R205 VTAIL.n389 VTAIL.n388 185
R206 VTAIL.n391 VTAIL.n390 185
R207 VTAIL.n352 VTAIL.n351 185
R208 VTAIL.n397 VTAIL.n396 185
R209 VTAIL.n399 VTAIL.n398 185
R210 VTAIL.n348 VTAIL.n347 185
R211 VTAIL.n405 VTAIL.n404 185
R212 VTAIL.n408 VTAIL.n407 185
R213 VTAIL.n406 VTAIL.n344 185
R214 VTAIL.n413 VTAIL.n343 185
R215 VTAIL.n415 VTAIL.n414 185
R216 VTAIL.n417 VTAIL.n416 185
R217 VTAIL.n340 VTAIL.n339 185
R218 VTAIL.n423 VTAIL.n422 185
R219 VTAIL.n425 VTAIL.n424 185
R220 VTAIL.n336 VTAIL.n335 185
R221 VTAIL.n431 VTAIL.n430 185
R222 VTAIL.n433 VTAIL.n432 185
R223 VTAIL.n37 VTAIL.n36 185
R224 VTAIL.n34 VTAIL.n33 185
R225 VTAIL.n43 VTAIL.n42 185
R226 VTAIL.n45 VTAIL.n44 185
R227 VTAIL.n30 VTAIL.n29 185
R228 VTAIL.n51 VTAIL.n50 185
R229 VTAIL.n53 VTAIL.n52 185
R230 VTAIL.n26 VTAIL.n25 185
R231 VTAIL.n59 VTAIL.n58 185
R232 VTAIL.n61 VTAIL.n60 185
R233 VTAIL.n22 VTAIL.n21 185
R234 VTAIL.n67 VTAIL.n66 185
R235 VTAIL.n69 VTAIL.n68 185
R236 VTAIL.n18 VTAIL.n17 185
R237 VTAIL.n75 VTAIL.n74 185
R238 VTAIL.n78 VTAIL.n77 185
R239 VTAIL.n76 VTAIL.n14 185
R240 VTAIL.n83 VTAIL.n13 185
R241 VTAIL.n85 VTAIL.n84 185
R242 VTAIL.n87 VTAIL.n86 185
R243 VTAIL.n10 VTAIL.n9 185
R244 VTAIL.n93 VTAIL.n92 185
R245 VTAIL.n95 VTAIL.n94 185
R246 VTAIL.n6 VTAIL.n5 185
R247 VTAIL.n101 VTAIL.n100 185
R248 VTAIL.n103 VTAIL.n102 185
R249 VTAIL.n327 VTAIL.n326 185
R250 VTAIL.n325 VTAIL.n324 185
R251 VTAIL.n230 VTAIL.n229 185
R252 VTAIL.n319 VTAIL.n318 185
R253 VTAIL.n317 VTAIL.n316 185
R254 VTAIL.n234 VTAIL.n233 185
R255 VTAIL.n311 VTAIL.n310 185
R256 VTAIL.n309 VTAIL.n308 185
R257 VTAIL.n307 VTAIL.n237 185
R258 VTAIL.n241 VTAIL.n238 185
R259 VTAIL.n302 VTAIL.n301 185
R260 VTAIL.n300 VTAIL.n299 185
R261 VTAIL.n243 VTAIL.n242 185
R262 VTAIL.n294 VTAIL.n293 185
R263 VTAIL.n292 VTAIL.n291 185
R264 VTAIL.n247 VTAIL.n246 185
R265 VTAIL.n286 VTAIL.n285 185
R266 VTAIL.n284 VTAIL.n283 185
R267 VTAIL.n251 VTAIL.n250 185
R268 VTAIL.n278 VTAIL.n277 185
R269 VTAIL.n276 VTAIL.n275 185
R270 VTAIL.n255 VTAIL.n254 185
R271 VTAIL.n270 VTAIL.n269 185
R272 VTAIL.n268 VTAIL.n267 185
R273 VTAIL.n259 VTAIL.n258 185
R274 VTAIL.n262 VTAIL.n261 185
R275 VTAIL.n217 VTAIL.n216 185
R276 VTAIL.n215 VTAIL.n214 185
R277 VTAIL.n120 VTAIL.n119 185
R278 VTAIL.n209 VTAIL.n208 185
R279 VTAIL.n207 VTAIL.n206 185
R280 VTAIL.n124 VTAIL.n123 185
R281 VTAIL.n201 VTAIL.n200 185
R282 VTAIL.n199 VTAIL.n198 185
R283 VTAIL.n197 VTAIL.n127 185
R284 VTAIL.n131 VTAIL.n128 185
R285 VTAIL.n192 VTAIL.n191 185
R286 VTAIL.n190 VTAIL.n189 185
R287 VTAIL.n133 VTAIL.n132 185
R288 VTAIL.n184 VTAIL.n183 185
R289 VTAIL.n182 VTAIL.n181 185
R290 VTAIL.n137 VTAIL.n136 185
R291 VTAIL.n176 VTAIL.n175 185
R292 VTAIL.n174 VTAIL.n173 185
R293 VTAIL.n141 VTAIL.n140 185
R294 VTAIL.n168 VTAIL.n167 185
R295 VTAIL.n166 VTAIL.n165 185
R296 VTAIL.n145 VTAIL.n144 185
R297 VTAIL.n160 VTAIL.n159 185
R298 VTAIL.n158 VTAIL.n157 185
R299 VTAIL.n149 VTAIL.n148 185
R300 VTAIL.n152 VTAIL.n151 185
R301 VTAIL.t15 VTAIL.n260 147.659
R302 VTAIL.t3 VTAIL.n150 147.659
R303 VTAIL.t0 VTAIL.n365 147.659
R304 VTAIL.t18 VTAIL.n35 147.659
R305 VTAIL.n366 VTAIL.n363 104.615
R306 VTAIL.n373 VTAIL.n363 104.615
R307 VTAIL.n374 VTAIL.n373 104.615
R308 VTAIL.n374 VTAIL.n359 104.615
R309 VTAIL.n381 VTAIL.n359 104.615
R310 VTAIL.n382 VTAIL.n381 104.615
R311 VTAIL.n382 VTAIL.n355 104.615
R312 VTAIL.n389 VTAIL.n355 104.615
R313 VTAIL.n390 VTAIL.n389 104.615
R314 VTAIL.n390 VTAIL.n351 104.615
R315 VTAIL.n397 VTAIL.n351 104.615
R316 VTAIL.n398 VTAIL.n397 104.615
R317 VTAIL.n398 VTAIL.n347 104.615
R318 VTAIL.n405 VTAIL.n347 104.615
R319 VTAIL.n407 VTAIL.n405 104.615
R320 VTAIL.n407 VTAIL.n406 104.615
R321 VTAIL.n406 VTAIL.n343 104.615
R322 VTAIL.n415 VTAIL.n343 104.615
R323 VTAIL.n416 VTAIL.n415 104.615
R324 VTAIL.n416 VTAIL.n339 104.615
R325 VTAIL.n423 VTAIL.n339 104.615
R326 VTAIL.n424 VTAIL.n423 104.615
R327 VTAIL.n424 VTAIL.n335 104.615
R328 VTAIL.n431 VTAIL.n335 104.615
R329 VTAIL.n432 VTAIL.n431 104.615
R330 VTAIL.n36 VTAIL.n33 104.615
R331 VTAIL.n43 VTAIL.n33 104.615
R332 VTAIL.n44 VTAIL.n43 104.615
R333 VTAIL.n44 VTAIL.n29 104.615
R334 VTAIL.n51 VTAIL.n29 104.615
R335 VTAIL.n52 VTAIL.n51 104.615
R336 VTAIL.n52 VTAIL.n25 104.615
R337 VTAIL.n59 VTAIL.n25 104.615
R338 VTAIL.n60 VTAIL.n59 104.615
R339 VTAIL.n60 VTAIL.n21 104.615
R340 VTAIL.n67 VTAIL.n21 104.615
R341 VTAIL.n68 VTAIL.n67 104.615
R342 VTAIL.n68 VTAIL.n17 104.615
R343 VTAIL.n75 VTAIL.n17 104.615
R344 VTAIL.n77 VTAIL.n75 104.615
R345 VTAIL.n77 VTAIL.n76 104.615
R346 VTAIL.n76 VTAIL.n13 104.615
R347 VTAIL.n85 VTAIL.n13 104.615
R348 VTAIL.n86 VTAIL.n85 104.615
R349 VTAIL.n86 VTAIL.n9 104.615
R350 VTAIL.n93 VTAIL.n9 104.615
R351 VTAIL.n94 VTAIL.n93 104.615
R352 VTAIL.n94 VTAIL.n5 104.615
R353 VTAIL.n101 VTAIL.n5 104.615
R354 VTAIL.n102 VTAIL.n101 104.615
R355 VTAIL.n326 VTAIL.n325 104.615
R356 VTAIL.n325 VTAIL.n229 104.615
R357 VTAIL.n318 VTAIL.n229 104.615
R358 VTAIL.n318 VTAIL.n317 104.615
R359 VTAIL.n317 VTAIL.n233 104.615
R360 VTAIL.n310 VTAIL.n233 104.615
R361 VTAIL.n310 VTAIL.n309 104.615
R362 VTAIL.n309 VTAIL.n237 104.615
R363 VTAIL.n241 VTAIL.n237 104.615
R364 VTAIL.n301 VTAIL.n241 104.615
R365 VTAIL.n301 VTAIL.n300 104.615
R366 VTAIL.n300 VTAIL.n242 104.615
R367 VTAIL.n293 VTAIL.n242 104.615
R368 VTAIL.n293 VTAIL.n292 104.615
R369 VTAIL.n292 VTAIL.n246 104.615
R370 VTAIL.n285 VTAIL.n246 104.615
R371 VTAIL.n285 VTAIL.n284 104.615
R372 VTAIL.n284 VTAIL.n250 104.615
R373 VTAIL.n277 VTAIL.n250 104.615
R374 VTAIL.n277 VTAIL.n276 104.615
R375 VTAIL.n276 VTAIL.n254 104.615
R376 VTAIL.n269 VTAIL.n254 104.615
R377 VTAIL.n269 VTAIL.n268 104.615
R378 VTAIL.n268 VTAIL.n258 104.615
R379 VTAIL.n261 VTAIL.n258 104.615
R380 VTAIL.n216 VTAIL.n215 104.615
R381 VTAIL.n215 VTAIL.n119 104.615
R382 VTAIL.n208 VTAIL.n119 104.615
R383 VTAIL.n208 VTAIL.n207 104.615
R384 VTAIL.n207 VTAIL.n123 104.615
R385 VTAIL.n200 VTAIL.n123 104.615
R386 VTAIL.n200 VTAIL.n199 104.615
R387 VTAIL.n199 VTAIL.n127 104.615
R388 VTAIL.n131 VTAIL.n127 104.615
R389 VTAIL.n191 VTAIL.n131 104.615
R390 VTAIL.n191 VTAIL.n190 104.615
R391 VTAIL.n190 VTAIL.n132 104.615
R392 VTAIL.n183 VTAIL.n132 104.615
R393 VTAIL.n183 VTAIL.n182 104.615
R394 VTAIL.n182 VTAIL.n136 104.615
R395 VTAIL.n175 VTAIL.n136 104.615
R396 VTAIL.n175 VTAIL.n174 104.615
R397 VTAIL.n174 VTAIL.n140 104.615
R398 VTAIL.n167 VTAIL.n140 104.615
R399 VTAIL.n167 VTAIL.n166 104.615
R400 VTAIL.n166 VTAIL.n144 104.615
R401 VTAIL.n159 VTAIL.n144 104.615
R402 VTAIL.n159 VTAIL.n158 104.615
R403 VTAIL.n158 VTAIL.n148 104.615
R404 VTAIL.n151 VTAIL.n148 104.615
R405 VTAIL.n366 VTAIL.t0 52.3082
R406 VTAIL.n36 VTAIL.t18 52.3082
R407 VTAIL.n261 VTAIL.t15 52.3082
R408 VTAIL.n151 VTAIL.t3 52.3082
R409 VTAIL.n439 VTAIL.n438 42.5856
R410 VTAIL.n1 VTAIL.n0 42.5856
R411 VTAIL.n109 VTAIL.n108 42.5856
R412 VTAIL.n111 VTAIL.n110 42.5856
R413 VTAIL.n225 VTAIL.n224 42.5856
R414 VTAIL.n223 VTAIL.n222 42.5856
R415 VTAIL.n115 VTAIL.n114 42.5856
R416 VTAIL.n113 VTAIL.n112 42.5856
R417 VTAIL.n113 VTAIL.n111 35.7548
R418 VTAIL.n437 VTAIL.n331 32.2031
R419 VTAIL.n437 VTAIL.n436 30.8278
R420 VTAIL.n107 VTAIL.n106 30.8278
R421 VTAIL.n331 VTAIL.n330 30.8278
R422 VTAIL.n221 VTAIL.n220 30.8278
R423 VTAIL.n367 VTAIL.n365 15.6677
R424 VTAIL.n37 VTAIL.n35 15.6677
R425 VTAIL.n262 VTAIL.n260 15.6677
R426 VTAIL.n152 VTAIL.n150 15.6677
R427 VTAIL.n414 VTAIL.n413 13.1884
R428 VTAIL.n84 VTAIL.n83 13.1884
R429 VTAIL.n308 VTAIL.n307 13.1884
R430 VTAIL.n198 VTAIL.n197 13.1884
R431 VTAIL.n368 VTAIL.n364 12.8005
R432 VTAIL.n412 VTAIL.n344 12.8005
R433 VTAIL.n417 VTAIL.n342 12.8005
R434 VTAIL.n38 VTAIL.n34 12.8005
R435 VTAIL.n82 VTAIL.n14 12.8005
R436 VTAIL.n87 VTAIL.n12 12.8005
R437 VTAIL.n311 VTAIL.n236 12.8005
R438 VTAIL.n306 VTAIL.n238 12.8005
R439 VTAIL.n263 VTAIL.n259 12.8005
R440 VTAIL.n201 VTAIL.n126 12.8005
R441 VTAIL.n196 VTAIL.n128 12.8005
R442 VTAIL.n153 VTAIL.n149 12.8005
R443 VTAIL.n372 VTAIL.n371 12.0247
R444 VTAIL.n409 VTAIL.n408 12.0247
R445 VTAIL.n418 VTAIL.n340 12.0247
R446 VTAIL.n42 VTAIL.n41 12.0247
R447 VTAIL.n79 VTAIL.n78 12.0247
R448 VTAIL.n88 VTAIL.n10 12.0247
R449 VTAIL.n312 VTAIL.n234 12.0247
R450 VTAIL.n303 VTAIL.n302 12.0247
R451 VTAIL.n267 VTAIL.n266 12.0247
R452 VTAIL.n202 VTAIL.n124 12.0247
R453 VTAIL.n193 VTAIL.n192 12.0247
R454 VTAIL.n157 VTAIL.n156 12.0247
R455 VTAIL.n375 VTAIL.n362 11.249
R456 VTAIL.n404 VTAIL.n346 11.249
R457 VTAIL.n422 VTAIL.n421 11.249
R458 VTAIL.n45 VTAIL.n32 11.249
R459 VTAIL.n74 VTAIL.n16 11.249
R460 VTAIL.n92 VTAIL.n91 11.249
R461 VTAIL.n316 VTAIL.n315 11.249
R462 VTAIL.n299 VTAIL.n240 11.249
R463 VTAIL.n270 VTAIL.n257 11.249
R464 VTAIL.n206 VTAIL.n205 11.249
R465 VTAIL.n189 VTAIL.n130 11.249
R466 VTAIL.n160 VTAIL.n147 11.249
R467 VTAIL.n376 VTAIL.n360 10.4732
R468 VTAIL.n403 VTAIL.n348 10.4732
R469 VTAIL.n425 VTAIL.n338 10.4732
R470 VTAIL.n46 VTAIL.n30 10.4732
R471 VTAIL.n73 VTAIL.n18 10.4732
R472 VTAIL.n95 VTAIL.n8 10.4732
R473 VTAIL.n319 VTAIL.n232 10.4732
R474 VTAIL.n298 VTAIL.n243 10.4732
R475 VTAIL.n271 VTAIL.n255 10.4732
R476 VTAIL.n209 VTAIL.n122 10.4732
R477 VTAIL.n188 VTAIL.n133 10.4732
R478 VTAIL.n161 VTAIL.n145 10.4732
R479 VTAIL.n380 VTAIL.n379 9.69747
R480 VTAIL.n400 VTAIL.n399 9.69747
R481 VTAIL.n426 VTAIL.n336 9.69747
R482 VTAIL.n50 VTAIL.n49 9.69747
R483 VTAIL.n70 VTAIL.n69 9.69747
R484 VTAIL.n96 VTAIL.n6 9.69747
R485 VTAIL.n320 VTAIL.n230 9.69747
R486 VTAIL.n295 VTAIL.n294 9.69747
R487 VTAIL.n275 VTAIL.n274 9.69747
R488 VTAIL.n210 VTAIL.n120 9.69747
R489 VTAIL.n185 VTAIL.n184 9.69747
R490 VTAIL.n165 VTAIL.n164 9.69747
R491 VTAIL.n436 VTAIL.n435 9.45567
R492 VTAIL.n106 VTAIL.n105 9.45567
R493 VTAIL.n330 VTAIL.n329 9.45567
R494 VTAIL.n220 VTAIL.n219 9.45567
R495 VTAIL.n334 VTAIL.n333 9.3005
R496 VTAIL.n429 VTAIL.n428 9.3005
R497 VTAIL.n427 VTAIL.n426 9.3005
R498 VTAIL.n338 VTAIL.n337 9.3005
R499 VTAIL.n421 VTAIL.n420 9.3005
R500 VTAIL.n419 VTAIL.n418 9.3005
R501 VTAIL.n342 VTAIL.n341 9.3005
R502 VTAIL.n387 VTAIL.n386 9.3005
R503 VTAIL.n385 VTAIL.n384 9.3005
R504 VTAIL.n358 VTAIL.n357 9.3005
R505 VTAIL.n379 VTAIL.n378 9.3005
R506 VTAIL.n377 VTAIL.n376 9.3005
R507 VTAIL.n362 VTAIL.n361 9.3005
R508 VTAIL.n371 VTAIL.n370 9.3005
R509 VTAIL.n369 VTAIL.n368 9.3005
R510 VTAIL.n354 VTAIL.n353 9.3005
R511 VTAIL.n393 VTAIL.n392 9.3005
R512 VTAIL.n395 VTAIL.n394 9.3005
R513 VTAIL.n350 VTAIL.n349 9.3005
R514 VTAIL.n401 VTAIL.n400 9.3005
R515 VTAIL.n403 VTAIL.n402 9.3005
R516 VTAIL.n346 VTAIL.n345 9.3005
R517 VTAIL.n410 VTAIL.n409 9.3005
R518 VTAIL.n412 VTAIL.n411 9.3005
R519 VTAIL.n435 VTAIL.n434 9.3005
R520 VTAIL.n4 VTAIL.n3 9.3005
R521 VTAIL.n99 VTAIL.n98 9.3005
R522 VTAIL.n97 VTAIL.n96 9.3005
R523 VTAIL.n8 VTAIL.n7 9.3005
R524 VTAIL.n91 VTAIL.n90 9.3005
R525 VTAIL.n89 VTAIL.n88 9.3005
R526 VTAIL.n12 VTAIL.n11 9.3005
R527 VTAIL.n57 VTAIL.n56 9.3005
R528 VTAIL.n55 VTAIL.n54 9.3005
R529 VTAIL.n28 VTAIL.n27 9.3005
R530 VTAIL.n49 VTAIL.n48 9.3005
R531 VTAIL.n47 VTAIL.n46 9.3005
R532 VTAIL.n32 VTAIL.n31 9.3005
R533 VTAIL.n41 VTAIL.n40 9.3005
R534 VTAIL.n39 VTAIL.n38 9.3005
R535 VTAIL.n24 VTAIL.n23 9.3005
R536 VTAIL.n63 VTAIL.n62 9.3005
R537 VTAIL.n65 VTAIL.n64 9.3005
R538 VTAIL.n20 VTAIL.n19 9.3005
R539 VTAIL.n71 VTAIL.n70 9.3005
R540 VTAIL.n73 VTAIL.n72 9.3005
R541 VTAIL.n16 VTAIL.n15 9.3005
R542 VTAIL.n80 VTAIL.n79 9.3005
R543 VTAIL.n82 VTAIL.n81 9.3005
R544 VTAIL.n105 VTAIL.n104 9.3005
R545 VTAIL.n288 VTAIL.n287 9.3005
R546 VTAIL.n290 VTAIL.n289 9.3005
R547 VTAIL.n245 VTAIL.n244 9.3005
R548 VTAIL.n296 VTAIL.n295 9.3005
R549 VTAIL.n298 VTAIL.n297 9.3005
R550 VTAIL.n240 VTAIL.n239 9.3005
R551 VTAIL.n304 VTAIL.n303 9.3005
R552 VTAIL.n306 VTAIL.n305 9.3005
R553 VTAIL.n329 VTAIL.n328 9.3005
R554 VTAIL.n228 VTAIL.n227 9.3005
R555 VTAIL.n323 VTAIL.n322 9.3005
R556 VTAIL.n321 VTAIL.n320 9.3005
R557 VTAIL.n232 VTAIL.n231 9.3005
R558 VTAIL.n315 VTAIL.n314 9.3005
R559 VTAIL.n313 VTAIL.n312 9.3005
R560 VTAIL.n236 VTAIL.n235 9.3005
R561 VTAIL.n249 VTAIL.n248 9.3005
R562 VTAIL.n282 VTAIL.n281 9.3005
R563 VTAIL.n280 VTAIL.n279 9.3005
R564 VTAIL.n253 VTAIL.n252 9.3005
R565 VTAIL.n274 VTAIL.n273 9.3005
R566 VTAIL.n272 VTAIL.n271 9.3005
R567 VTAIL.n257 VTAIL.n256 9.3005
R568 VTAIL.n266 VTAIL.n265 9.3005
R569 VTAIL.n264 VTAIL.n263 9.3005
R570 VTAIL.n178 VTAIL.n177 9.3005
R571 VTAIL.n180 VTAIL.n179 9.3005
R572 VTAIL.n135 VTAIL.n134 9.3005
R573 VTAIL.n186 VTAIL.n185 9.3005
R574 VTAIL.n188 VTAIL.n187 9.3005
R575 VTAIL.n130 VTAIL.n129 9.3005
R576 VTAIL.n194 VTAIL.n193 9.3005
R577 VTAIL.n196 VTAIL.n195 9.3005
R578 VTAIL.n219 VTAIL.n218 9.3005
R579 VTAIL.n118 VTAIL.n117 9.3005
R580 VTAIL.n213 VTAIL.n212 9.3005
R581 VTAIL.n211 VTAIL.n210 9.3005
R582 VTAIL.n122 VTAIL.n121 9.3005
R583 VTAIL.n205 VTAIL.n204 9.3005
R584 VTAIL.n203 VTAIL.n202 9.3005
R585 VTAIL.n126 VTAIL.n125 9.3005
R586 VTAIL.n139 VTAIL.n138 9.3005
R587 VTAIL.n172 VTAIL.n171 9.3005
R588 VTAIL.n170 VTAIL.n169 9.3005
R589 VTAIL.n143 VTAIL.n142 9.3005
R590 VTAIL.n164 VTAIL.n163 9.3005
R591 VTAIL.n162 VTAIL.n161 9.3005
R592 VTAIL.n147 VTAIL.n146 9.3005
R593 VTAIL.n156 VTAIL.n155 9.3005
R594 VTAIL.n154 VTAIL.n153 9.3005
R595 VTAIL.n383 VTAIL.n358 8.92171
R596 VTAIL.n396 VTAIL.n350 8.92171
R597 VTAIL.n430 VTAIL.n429 8.92171
R598 VTAIL.n53 VTAIL.n28 8.92171
R599 VTAIL.n66 VTAIL.n20 8.92171
R600 VTAIL.n100 VTAIL.n99 8.92171
R601 VTAIL.n324 VTAIL.n323 8.92171
R602 VTAIL.n291 VTAIL.n245 8.92171
R603 VTAIL.n278 VTAIL.n253 8.92171
R604 VTAIL.n214 VTAIL.n213 8.92171
R605 VTAIL.n181 VTAIL.n135 8.92171
R606 VTAIL.n168 VTAIL.n143 8.92171
R607 VTAIL.n384 VTAIL.n356 8.14595
R608 VTAIL.n395 VTAIL.n352 8.14595
R609 VTAIL.n433 VTAIL.n334 8.14595
R610 VTAIL.n54 VTAIL.n26 8.14595
R611 VTAIL.n65 VTAIL.n22 8.14595
R612 VTAIL.n103 VTAIL.n4 8.14595
R613 VTAIL.n327 VTAIL.n228 8.14595
R614 VTAIL.n290 VTAIL.n247 8.14595
R615 VTAIL.n279 VTAIL.n251 8.14595
R616 VTAIL.n217 VTAIL.n118 8.14595
R617 VTAIL.n180 VTAIL.n137 8.14595
R618 VTAIL.n169 VTAIL.n141 8.14595
R619 VTAIL.n388 VTAIL.n387 7.3702
R620 VTAIL.n392 VTAIL.n391 7.3702
R621 VTAIL.n434 VTAIL.n332 7.3702
R622 VTAIL.n58 VTAIL.n57 7.3702
R623 VTAIL.n62 VTAIL.n61 7.3702
R624 VTAIL.n104 VTAIL.n2 7.3702
R625 VTAIL.n328 VTAIL.n226 7.3702
R626 VTAIL.n287 VTAIL.n286 7.3702
R627 VTAIL.n283 VTAIL.n282 7.3702
R628 VTAIL.n218 VTAIL.n116 7.3702
R629 VTAIL.n177 VTAIL.n176 7.3702
R630 VTAIL.n173 VTAIL.n172 7.3702
R631 VTAIL.n388 VTAIL.n354 6.59444
R632 VTAIL.n391 VTAIL.n354 6.59444
R633 VTAIL.n436 VTAIL.n332 6.59444
R634 VTAIL.n58 VTAIL.n24 6.59444
R635 VTAIL.n61 VTAIL.n24 6.59444
R636 VTAIL.n106 VTAIL.n2 6.59444
R637 VTAIL.n330 VTAIL.n226 6.59444
R638 VTAIL.n286 VTAIL.n249 6.59444
R639 VTAIL.n283 VTAIL.n249 6.59444
R640 VTAIL.n220 VTAIL.n116 6.59444
R641 VTAIL.n176 VTAIL.n139 6.59444
R642 VTAIL.n173 VTAIL.n139 6.59444
R643 VTAIL.n387 VTAIL.n356 5.81868
R644 VTAIL.n392 VTAIL.n352 5.81868
R645 VTAIL.n434 VTAIL.n433 5.81868
R646 VTAIL.n57 VTAIL.n26 5.81868
R647 VTAIL.n62 VTAIL.n22 5.81868
R648 VTAIL.n104 VTAIL.n103 5.81868
R649 VTAIL.n328 VTAIL.n327 5.81868
R650 VTAIL.n287 VTAIL.n247 5.81868
R651 VTAIL.n282 VTAIL.n251 5.81868
R652 VTAIL.n218 VTAIL.n217 5.81868
R653 VTAIL.n177 VTAIL.n137 5.81868
R654 VTAIL.n172 VTAIL.n141 5.81868
R655 VTAIL.n384 VTAIL.n383 5.04292
R656 VTAIL.n396 VTAIL.n395 5.04292
R657 VTAIL.n430 VTAIL.n334 5.04292
R658 VTAIL.n54 VTAIL.n53 5.04292
R659 VTAIL.n66 VTAIL.n65 5.04292
R660 VTAIL.n100 VTAIL.n4 5.04292
R661 VTAIL.n324 VTAIL.n228 5.04292
R662 VTAIL.n291 VTAIL.n290 5.04292
R663 VTAIL.n279 VTAIL.n278 5.04292
R664 VTAIL.n214 VTAIL.n118 5.04292
R665 VTAIL.n181 VTAIL.n180 5.04292
R666 VTAIL.n169 VTAIL.n168 5.04292
R667 VTAIL.n264 VTAIL.n260 4.38563
R668 VTAIL.n154 VTAIL.n150 4.38563
R669 VTAIL.n369 VTAIL.n365 4.38563
R670 VTAIL.n39 VTAIL.n35 4.38563
R671 VTAIL.n380 VTAIL.n358 4.26717
R672 VTAIL.n399 VTAIL.n350 4.26717
R673 VTAIL.n429 VTAIL.n336 4.26717
R674 VTAIL.n50 VTAIL.n28 4.26717
R675 VTAIL.n69 VTAIL.n20 4.26717
R676 VTAIL.n99 VTAIL.n6 4.26717
R677 VTAIL.n323 VTAIL.n230 4.26717
R678 VTAIL.n294 VTAIL.n245 4.26717
R679 VTAIL.n275 VTAIL.n253 4.26717
R680 VTAIL.n213 VTAIL.n120 4.26717
R681 VTAIL.n184 VTAIL.n135 4.26717
R682 VTAIL.n165 VTAIL.n143 4.26717
R683 VTAIL.n115 VTAIL.n113 3.55222
R684 VTAIL.n221 VTAIL.n115 3.55222
R685 VTAIL.n225 VTAIL.n223 3.55222
R686 VTAIL.n331 VTAIL.n225 3.55222
R687 VTAIL.n111 VTAIL.n109 3.55222
R688 VTAIL.n109 VTAIL.n107 3.55222
R689 VTAIL.n439 VTAIL.n437 3.55222
R690 VTAIL.n379 VTAIL.n360 3.49141
R691 VTAIL.n400 VTAIL.n348 3.49141
R692 VTAIL.n426 VTAIL.n425 3.49141
R693 VTAIL.n49 VTAIL.n30 3.49141
R694 VTAIL.n70 VTAIL.n18 3.49141
R695 VTAIL.n96 VTAIL.n95 3.49141
R696 VTAIL.n320 VTAIL.n319 3.49141
R697 VTAIL.n295 VTAIL.n243 3.49141
R698 VTAIL.n274 VTAIL.n255 3.49141
R699 VTAIL.n210 VTAIL.n209 3.49141
R700 VTAIL.n185 VTAIL.n133 3.49141
R701 VTAIL.n164 VTAIL.n145 3.49141
R702 VTAIL VTAIL.n1 2.72248
R703 VTAIL.n376 VTAIL.n375 2.71565
R704 VTAIL.n404 VTAIL.n403 2.71565
R705 VTAIL.n422 VTAIL.n338 2.71565
R706 VTAIL.n46 VTAIL.n45 2.71565
R707 VTAIL.n74 VTAIL.n73 2.71565
R708 VTAIL.n92 VTAIL.n8 2.71565
R709 VTAIL.n316 VTAIL.n232 2.71565
R710 VTAIL.n299 VTAIL.n298 2.71565
R711 VTAIL.n271 VTAIL.n270 2.71565
R712 VTAIL.n206 VTAIL.n122 2.71565
R713 VTAIL.n189 VTAIL.n188 2.71565
R714 VTAIL.n161 VTAIL.n160 2.71565
R715 VTAIL.n223 VTAIL.n221 2.24619
R716 VTAIL.n107 VTAIL.n1 2.24619
R717 VTAIL.n372 VTAIL.n362 1.93989
R718 VTAIL.n408 VTAIL.n346 1.93989
R719 VTAIL.n421 VTAIL.n340 1.93989
R720 VTAIL.n42 VTAIL.n32 1.93989
R721 VTAIL.n78 VTAIL.n16 1.93989
R722 VTAIL.n91 VTAIL.n10 1.93989
R723 VTAIL.n315 VTAIL.n234 1.93989
R724 VTAIL.n302 VTAIL.n240 1.93989
R725 VTAIL.n267 VTAIL.n257 1.93989
R726 VTAIL.n205 VTAIL.n124 1.93989
R727 VTAIL.n192 VTAIL.n130 1.93989
R728 VTAIL.n157 VTAIL.n147 1.93989
R729 VTAIL.n371 VTAIL.n364 1.16414
R730 VTAIL.n409 VTAIL.n344 1.16414
R731 VTAIL.n418 VTAIL.n417 1.16414
R732 VTAIL.n41 VTAIL.n34 1.16414
R733 VTAIL.n79 VTAIL.n14 1.16414
R734 VTAIL.n88 VTAIL.n87 1.16414
R735 VTAIL.n312 VTAIL.n311 1.16414
R736 VTAIL.n303 VTAIL.n238 1.16414
R737 VTAIL.n266 VTAIL.n259 1.16414
R738 VTAIL.n202 VTAIL.n201 1.16414
R739 VTAIL.n193 VTAIL.n128 1.16414
R740 VTAIL.n156 VTAIL.n149 1.16414
R741 VTAIL.n438 VTAIL.t2 1.04867
R742 VTAIL.n438 VTAIL.t8 1.04867
R743 VTAIL.n0 VTAIL.t7 1.04867
R744 VTAIL.n0 VTAIL.t4 1.04867
R745 VTAIL.n108 VTAIL.t17 1.04867
R746 VTAIL.n108 VTAIL.t13 1.04867
R747 VTAIL.n110 VTAIL.t19 1.04867
R748 VTAIL.n110 VTAIL.t12 1.04867
R749 VTAIL.n224 VTAIL.t10 1.04867
R750 VTAIL.n224 VTAIL.t16 1.04867
R751 VTAIL.n222 VTAIL.t14 1.04867
R752 VTAIL.n222 VTAIL.t11 1.04867
R753 VTAIL.n114 VTAIL.t9 1.04867
R754 VTAIL.n114 VTAIL.t5 1.04867
R755 VTAIL.n112 VTAIL.t1 1.04867
R756 VTAIL.n112 VTAIL.t6 1.04867
R757 VTAIL VTAIL.n439 0.830241
R758 VTAIL.n368 VTAIL.n367 0.388379
R759 VTAIL.n413 VTAIL.n412 0.388379
R760 VTAIL.n414 VTAIL.n342 0.388379
R761 VTAIL.n38 VTAIL.n37 0.388379
R762 VTAIL.n83 VTAIL.n82 0.388379
R763 VTAIL.n84 VTAIL.n12 0.388379
R764 VTAIL.n308 VTAIL.n236 0.388379
R765 VTAIL.n307 VTAIL.n306 0.388379
R766 VTAIL.n263 VTAIL.n262 0.388379
R767 VTAIL.n198 VTAIL.n126 0.388379
R768 VTAIL.n197 VTAIL.n196 0.388379
R769 VTAIL.n153 VTAIL.n152 0.388379
R770 VTAIL.n370 VTAIL.n369 0.155672
R771 VTAIL.n370 VTAIL.n361 0.155672
R772 VTAIL.n377 VTAIL.n361 0.155672
R773 VTAIL.n378 VTAIL.n377 0.155672
R774 VTAIL.n378 VTAIL.n357 0.155672
R775 VTAIL.n385 VTAIL.n357 0.155672
R776 VTAIL.n386 VTAIL.n385 0.155672
R777 VTAIL.n386 VTAIL.n353 0.155672
R778 VTAIL.n393 VTAIL.n353 0.155672
R779 VTAIL.n394 VTAIL.n393 0.155672
R780 VTAIL.n394 VTAIL.n349 0.155672
R781 VTAIL.n401 VTAIL.n349 0.155672
R782 VTAIL.n402 VTAIL.n401 0.155672
R783 VTAIL.n402 VTAIL.n345 0.155672
R784 VTAIL.n410 VTAIL.n345 0.155672
R785 VTAIL.n411 VTAIL.n410 0.155672
R786 VTAIL.n411 VTAIL.n341 0.155672
R787 VTAIL.n419 VTAIL.n341 0.155672
R788 VTAIL.n420 VTAIL.n419 0.155672
R789 VTAIL.n420 VTAIL.n337 0.155672
R790 VTAIL.n427 VTAIL.n337 0.155672
R791 VTAIL.n428 VTAIL.n427 0.155672
R792 VTAIL.n428 VTAIL.n333 0.155672
R793 VTAIL.n435 VTAIL.n333 0.155672
R794 VTAIL.n40 VTAIL.n39 0.155672
R795 VTAIL.n40 VTAIL.n31 0.155672
R796 VTAIL.n47 VTAIL.n31 0.155672
R797 VTAIL.n48 VTAIL.n47 0.155672
R798 VTAIL.n48 VTAIL.n27 0.155672
R799 VTAIL.n55 VTAIL.n27 0.155672
R800 VTAIL.n56 VTAIL.n55 0.155672
R801 VTAIL.n56 VTAIL.n23 0.155672
R802 VTAIL.n63 VTAIL.n23 0.155672
R803 VTAIL.n64 VTAIL.n63 0.155672
R804 VTAIL.n64 VTAIL.n19 0.155672
R805 VTAIL.n71 VTAIL.n19 0.155672
R806 VTAIL.n72 VTAIL.n71 0.155672
R807 VTAIL.n72 VTAIL.n15 0.155672
R808 VTAIL.n80 VTAIL.n15 0.155672
R809 VTAIL.n81 VTAIL.n80 0.155672
R810 VTAIL.n81 VTAIL.n11 0.155672
R811 VTAIL.n89 VTAIL.n11 0.155672
R812 VTAIL.n90 VTAIL.n89 0.155672
R813 VTAIL.n90 VTAIL.n7 0.155672
R814 VTAIL.n97 VTAIL.n7 0.155672
R815 VTAIL.n98 VTAIL.n97 0.155672
R816 VTAIL.n98 VTAIL.n3 0.155672
R817 VTAIL.n105 VTAIL.n3 0.155672
R818 VTAIL.n329 VTAIL.n227 0.155672
R819 VTAIL.n322 VTAIL.n227 0.155672
R820 VTAIL.n322 VTAIL.n321 0.155672
R821 VTAIL.n321 VTAIL.n231 0.155672
R822 VTAIL.n314 VTAIL.n231 0.155672
R823 VTAIL.n314 VTAIL.n313 0.155672
R824 VTAIL.n313 VTAIL.n235 0.155672
R825 VTAIL.n305 VTAIL.n235 0.155672
R826 VTAIL.n305 VTAIL.n304 0.155672
R827 VTAIL.n304 VTAIL.n239 0.155672
R828 VTAIL.n297 VTAIL.n239 0.155672
R829 VTAIL.n297 VTAIL.n296 0.155672
R830 VTAIL.n296 VTAIL.n244 0.155672
R831 VTAIL.n289 VTAIL.n244 0.155672
R832 VTAIL.n289 VTAIL.n288 0.155672
R833 VTAIL.n288 VTAIL.n248 0.155672
R834 VTAIL.n281 VTAIL.n248 0.155672
R835 VTAIL.n281 VTAIL.n280 0.155672
R836 VTAIL.n280 VTAIL.n252 0.155672
R837 VTAIL.n273 VTAIL.n252 0.155672
R838 VTAIL.n273 VTAIL.n272 0.155672
R839 VTAIL.n272 VTAIL.n256 0.155672
R840 VTAIL.n265 VTAIL.n256 0.155672
R841 VTAIL.n265 VTAIL.n264 0.155672
R842 VTAIL.n219 VTAIL.n117 0.155672
R843 VTAIL.n212 VTAIL.n117 0.155672
R844 VTAIL.n212 VTAIL.n211 0.155672
R845 VTAIL.n211 VTAIL.n121 0.155672
R846 VTAIL.n204 VTAIL.n121 0.155672
R847 VTAIL.n204 VTAIL.n203 0.155672
R848 VTAIL.n203 VTAIL.n125 0.155672
R849 VTAIL.n195 VTAIL.n125 0.155672
R850 VTAIL.n195 VTAIL.n194 0.155672
R851 VTAIL.n194 VTAIL.n129 0.155672
R852 VTAIL.n187 VTAIL.n129 0.155672
R853 VTAIL.n187 VTAIL.n186 0.155672
R854 VTAIL.n186 VTAIL.n134 0.155672
R855 VTAIL.n179 VTAIL.n134 0.155672
R856 VTAIL.n179 VTAIL.n178 0.155672
R857 VTAIL.n178 VTAIL.n138 0.155672
R858 VTAIL.n171 VTAIL.n138 0.155672
R859 VTAIL.n171 VTAIL.n170 0.155672
R860 VTAIL.n170 VTAIL.n142 0.155672
R861 VTAIL.n163 VTAIL.n142 0.155672
R862 VTAIL.n163 VTAIL.n162 0.155672
R863 VTAIL.n162 VTAIL.n146 0.155672
R864 VTAIL.n155 VTAIL.n146 0.155672
R865 VTAIL.n155 VTAIL.n154 0.155672
R866 VDD1.n100 VDD1.n0 289.615
R867 VDD1.n207 VDD1.n107 289.615
R868 VDD1.n101 VDD1.n100 185
R869 VDD1.n99 VDD1.n98 185
R870 VDD1.n4 VDD1.n3 185
R871 VDD1.n93 VDD1.n92 185
R872 VDD1.n91 VDD1.n90 185
R873 VDD1.n8 VDD1.n7 185
R874 VDD1.n85 VDD1.n84 185
R875 VDD1.n83 VDD1.n82 185
R876 VDD1.n81 VDD1.n11 185
R877 VDD1.n15 VDD1.n12 185
R878 VDD1.n76 VDD1.n75 185
R879 VDD1.n74 VDD1.n73 185
R880 VDD1.n17 VDD1.n16 185
R881 VDD1.n68 VDD1.n67 185
R882 VDD1.n66 VDD1.n65 185
R883 VDD1.n21 VDD1.n20 185
R884 VDD1.n60 VDD1.n59 185
R885 VDD1.n58 VDD1.n57 185
R886 VDD1.n25 VDD1.n24 185
R887 VDD1.n52 VDD1.n51 185
R888 VDD1.n50 VDD1.n49 185
R889 VDD1.n29 VDD1.n28 185
R890 VDD1.n44 VDD1.n43 185
R891 VDD1.n42 VDD1.n41 185
R892 VDD1.n33 VDD1.n32 185
R893 VDD1.n36 VDD1.n35 185
R894 VDD1.n142 VDD1.n141 185
R895 VDD1.n139 VDD1.n138 185
R896 VDD1.n148 VDD1.n147 185
R897 VDD1.n150 VDD1.n149 185
R898 VDD1.n135 VDD1.n134 185
R899 VDD1.n156 VDD1.n155 185
R900 VDD1.n158 VDD1.n157 185
R901 VDD1.n131 VDD1.n130 185
R902 VDD1.n164 VDD1.n163 185
R903 VDD1.n166 VDD1.n165 185
R904 VDD1.n127 VDD1.n126 185
R905 VDD1.n172 VDD1.n171 185
R906 VDD1.n174 VDD1.n173 185
R907 VDD1.n123 VDD1.n122 185
R908 VDD1.n180 VDD1.n179 185
R909 VDD1.n183 VDD1.n182 185
R910 VDD1.n181 VDD1.n119 185
R911 VDD1.n188 VDD1.n118 185
R912 VDD1.n190 VDD1.n189 185
R913 VDD1.n192 VDD1.n191 185
R914 VDD1.n115 VDD1.n114 185
R915 VDD1.n198 VDD1.n197 185
R916 VDD1.n200 VDD1.n199 185
R917 VDD1.n111 VDD1.n110 185
R918 VDD1.n206 VDD1.n205 185
R919 VDD1.n208 VDD1.n207 185
R920 VDD1.t3 VDD1.n34 147.659
R921 VDD1.t0 VDD1.n140 147.659
R922 VDD1.n100 VDD1.n99 104.615
R923 VDD1.n99 VDD1.n3 104.615
R924 VDD1.n92 VDD1.n3 104.615
R925 VDD1.n92 VDD1.n91 104.615
R926 VDD1.n91 VDD1.n7 104.615
R927 VDD1.n84 VDD1.n7 104.615
R928 VDD1.n84 VDD1.n83 104.615
R929 VDD1.n83 VDD1.n11 104.615
R930 VDD1.n15 VDD1.n11 104.615
R931 VDD1.n75 VDD1.n15 104.615
R932 VDD1.n75 VDD1.n74 104.615
R933 VDD1.n74 VDD1.n16 104.615
R934 VDD1.n67 VDD1.n16 104.615
R935 VDD1.n67 VDD1.n66 104.615
R936 VDD1.n66 VDD1.n20 104.615
R937 VDD1.n59 VDD1.n20 104.615
R938 VDD1.n59 VDD1.n58 104.615
R939 VDD1.n58 VDD1.n24 104.615
R940 VDD1.n51 VDD1.n24 104.615
R941 VDD1.n51 VDD1.n50 104.615
R942 VDD1.n50 VDD1.n28 104.615
R943 VDD1.n43 VDD1.n28 104.615
R944 VDD1.n43 VDD1.n42 104.615
R945 VDD1.n42 VDD1.n32 104.615
R946 VDD1.n35 VDD1.n32 104.615
R947 VDD1.n141 VDD1.n138 104.615
R948 VDD1.n148 VDD1.n138 104.615
R949 VDD1.n149 VDD1.n148 104.615
R950 VDD1.n149 VDD1.n134 104.615
R951 VDD1.n156 VDD1.n134 104.615
R952 VDD1.n157 VDD1.n156 104.615
R953 VDD1.n157 VDD1.n130 104.615
R954 VDD1.n164 VDD1.n130 104.615
R955 VDD1.n165 VDD1.n164 104.615
R956 VDD1.n165 VDD1.n126 104.615
R957 VDD1.n172 VDD1.n126 104.615
R958 VDD1.n173 VDD1.n172 104.615
R959 VDD1.n173 VDD1.n122 104.615
R960 VDD1.n180 VDD1.n122 104.615
R961 VDD1.n182 VDD1.n180 104.615
R962 VDD1.n182 VDD1.n181 104.615
R963 VDD1.n181 VDD1.n118 104.615
R964 VDD1.n190 VDD1.n118 104.615
R965 VDD1.n191 VDD1.n190 104.615
R966 VDD1.n191 VDD1.n114 104.615
R967 VDD1.n198 VDD1.n114 104.615
R968 VDD1.n199 VDD1.n198 104.615
R969 VDD1.n199 VDD1.n110 104.615
R970 VDD1.n206 VDD1.n110 104.615
R971 VDD1.n207 VDD1.n206 104.615
R972 VDD1.n215 VDD1.n214 61.8729
R973 VDD1.n106 VDD1.n105 59.2644
R974 VDD1.n213 VDD1.n212 59.2644
R975 VDD1.n217 VDD1.n216 59.2642
R976 VDD1.n217 VDD1.n215 59.2293
R977 VDD1.n35 VDD1.t3 52.3082
R978 VDD1.n141 VDD1.t0 52.3082
R979 VDD1.n106 VDD1.n104 51.0583
R980 VDD1.n213 VDD1.n211 51.0583
R981 VDD1.n36 VDD1.n34 15.6677
R982 VDD1.n142 VDD1.n140 15.6677
R983 VDD1.n82 VDD1.n81 13.1884
R984 VDD1.n189 VDD1.n188 13.1884
R985 VDD1.n85 VDD1.n10 12.8005
R986 VDD1.n80 VDD1.n12 12.8005
R987 VDD1.n37 VDD1.n33 12.8005
R988 VDD1.n143 VDD1.n139 12.8005
R989 VDD1.n187 VDD1.n119 12.8005
R990 VDD1.n192 VDD1.n117 12.8005
R991 VDD1.n86 VDD1.n8 12.0247
R992 VDD1.n77 VDD1.n76 12.0247
R993 VDD1.n41 VDD1.n40 12.0247
R994 VDD1.n147 VDD1.n146 12.0247
R995 VDD1.n184 VDD1.n183 12.0247
R996 VDD1.n193 VDD1.n115 12.0247
R997 VDD1.n90 VDD1.n89 11.249
R998 VDD1.n73 VDD1.n14 11.249
R999 VDD1.n44 VDD1.n31 11.249
R1000 VDD1.n150 VDD1.n137 11.249
R1001 VDD1.n179 VDD1.n121 11.249
R1002 VDD1.n197 VDD1.n196 11.249
R1003 VDD1.n93 VDD1.n6 10.4732
R1004 VDD1.n72 VDD1.n17 10.4732
R1005 VDD1.n45 VDD1.n29 10.4732
R1006 VDD1.n151 VDD1.n135 10.4732
R1007 VDD1.n178 VDD1.n123 10.4732
R1008 VDD1.n200 VDD1.n113 10.4732
R1009 VDD1.n94 VDD1.n4 9.69747
R1010 VDD1.n69 VDD1.n68 9.69747
R1011 VDD1.n49 VDD1.n48 9.69747
R1012 VDD1.n155 VDD1.n154 9.69747
R1013 VDD1.n175 VDD1.n174 9.69747
R1014 VDD1.n201 VDD1.n111 9.69747
R1015 VDD1.n104 VDD1.n103 9.45567
R1016 VDD1.n211 VDD1.n210 9.45567
R1017 VDD1.n62 VDD1.n61 9.3005
R1018 VDD1.n64 VDD1.n63 9.3005
R1019 VDD1.n19 VDD1.n18 9.3005
R1020 VDD1.n70 VDD1.n69 9.3005
R1021 VDD1.n72 VDD1.n71 9.3005
R1022 VDD1.n14 VDD1.n13 9.3005
R1023 VDD1.n78 VDD1.n77 9.3005
R1024 VDD1.n80 VDD1.n79 9.3005
R1025 VDD1.n103 VDD1.n102 9.3005
R1026 VDD1.n2 VDD1.n1 9.3005
R1027 VDD1.n97 VDD1.n96 9.3005
R1028 VDD1.n95 VDD1.n94 9.3005
R1029 VDD1.n6 VDD1.n5 9.3005
R1030 VDD1.n89 VDD1.n88 9.3005
R1031 VDD1.n87 VDD1.n86 9.3005
R1032 VDD1.n10 VDD1.n9 9.3005
R1033 VDD1.n23 VDD1.n22 9.3005
R1034 VDD1.n56 VDD1.n55 9.3005
R1035 VDD1.n54 VDD1.n53 9.3005
R1036 VDD1.n27 VDD1.n26 9.3005
R1037 VDD1.n48 VDD1.n47 9.3005
R1038 VDD1.n46 VDD1.n45 9.3005
R1039 VDD1.n31 VDD1.n30 9.3005
R1040 VDD1.n40 VDD1.n39 9.3005
R1041 VDD1.n38 VDD1.n37 9.3005
R1042 VDD1.n109 VDD1.n108 9.3005
R1043 VDD1.n204 VDD1.n203 9.3005
R1044 VDD1.n202 VDD1.n201 9.3005
R1045 VDD1.n113 VDD1.n112 9.3005
R1046 VDD1.n196 VDD1.n195 9.3005
R1047 VDD1.n194 VDD1.n193 9.3005
R1048 VDD1.n117 VDD1.n116 9.3005
R1049 VDD1.n162 VDD1.n161 9.3005
R1050 VDD1.n160 VDD1.n159 9.3005
R1051 VDD1.n133 VDD1.n132 9.3005
R1052 VDD1.n154 VDD1.n153 9.3005
R1053 VDD1.n152 VDD1.n151 9.3005
R1054 VDD1.n137 VDD1.n136 9.3005
R1055 VDD1.n146 VDD1.n145 9.3005
R1056 VDD1.n144 VDD1.n143 9.3005
R1057 VDD1.n129 VDD1.n128 9.3005
R1058 VDD1.n168 VDD1.n167 9.3005
R1059 VDD1.n170 VDD1.n169 9.3005
R1060 VDD1.n125 VDD1.n124 9.3005
R1061 VDD1.n176 VDD1.n175 9.3005
R1062 VDD1.n178 VDD1.n177 9.3005
R1063 VDD1.n121 VDD1.n120 9.3005
R1064 VDD1.n185 VDD1.n184 9.3005
R1065 VDD1.n187 VDD1.n186 9.3005
R1066 VDD1.n210 VDD1.n209 9.3005
R1067 VDD1.n98 VDD1.n97 8.92171
R1068 VDD1.n65 VDD1.n19 8.92171
R1069 VDD1.n52 VDD1.n27 8.92171
R1070 VDD1.n158 VDD1.n133 8.92171
R1071 VDD1.n171 VDD1.n125 8.92171
R1072 VDD1.n205 VDD1.n204 8.92171
R1073 VDD1.n101 VDD1.n2 8.14595
R1074 VDD1.n64 VDD1.n21 8.14595
R1075 VDD1.n53 VDD1.n25 8.14595
R1076 VDD1.n159 VDD1.n131 8.14595
R1077 VDD1.n170 VDD1.n127 8.14595
R1078 VDD1.n208 VDD1.n109 8.14595
R1079 VDD1.n102 VDD1.n0 7.3702
R1080 VDD1.n61 VDD1.n60 7.3702
R1081 VDD1.n57 VDD1.n56 7.3702
R1082 VDD1.n163 VDD1.n162 7.3702
R1083 VDD1.n167 VDD1.n166 7.3702
R1084 VDD1.n209 VDD1.n107 7.3702
R1085 VDD1.n104 VDD1.n0 6.59444
R1086 VDD1.n60 VDD1.n23 6.59444
R1087 VDD1.n57 VDD1.n23 6.59444
R1088 VDD1.n163 VDD1.n129 6.59444
R1089 VDD1.n166 VDD1.n129 6.59444
R1090 VDD1.n211 VDD1.n107 6.59444
R1091 VDD1.n102 VDD1.n101 5.81868
R1092 VDD1.n61 VDD1.n21 5.81868
R1093 VDD1.n56 VDD1.n25 5.81868
R1094 VDD1.n162 VDD1.n131 5.81868
R1095 VDD1.n167 VDD1.n127 5.81868
R1096 VDD1.n209 VDD1.n208 5.81868
R1097 VDD1.n98 VDD1.n2 5.04292
R1098 VDD1.n65 VDD1.n64 5.04292
R1099 VDD1.n53 VDD1.n52 5.04292
R1100 VDD1.n159 VDD1.n158 5.04292
R1101 VDD1.n171 VDD1.n170 5.04292
R1102 VDD1.n205 VDD1.n109 5.04292
R1103 VDD1.n38 VDD1.n34 4.38563
R1104 VDD1.n144 VDD1.n140 4.38563
R1105 VDD1.n97 VDD1.n4 4.26717
R1106 VDD1.n68 VDD1.n19 4.26717
R1107 VDD1.n49 VDD1.n27 4.26717
R1108 VDD1.n155 VDD1.n133 4.26717
R1109 VDD1.n174 VDD1.n125 4.26717
R1110 VDD1.n204 VDD1.n111 4.26717
R1111 VDD1.n94 VDD1.n93 3.49141
R1112 VDD1.n69 VDD1.n17 3.49141
R1113 VDD1.n48 VDD1.n29 3.49141
R1114 VDD1.n154 VDD1.n135 3.49141
R1115 VDD1.n175 VDD1.n123 3.49141
R1116 VDD1.n201 VDD1.n200 3.49141
R1117 VDD1.n90 VDD1.n6 2.71565
R1118 VDD1.n73 VDD1.n72 2.71565
R1119 VDD1.n45 VDD1.n44 2.71565
R1120 VDD1.n151 VDD1.n150 2.71565
R1121 VDD1.n179 VDD1.n178 2.71565
R1122 VDD1.n197 VDD1.n113 2.71565
R1123 VDD1 VDD1.n217 2.6061
R1124 VDD1.n89 VDD1.n8 1.93989
R1125 VDD1.n76 VDD1.n14 1.93989
R1126 VDD1.n41 VDD1.n31 1.93989
R1127 VDD1.n147 VDD1.n137 1.93989
R1128 VDD1.n183 VDD1.n121 1.93989
R1129 VDD1.n196 VDD1.n115 1.93989
R1130 VDD1.n86 VDD1.n85 1.16414
R1131 VDD1.n77 VDD1.n12 1.16414
R1132 VDD1.n40 VDD1.n33 1.16414
R1133 VDD1.n146 VDD1.n139 1.16414
R1134 VDD1.n184 VDD1.n119 1.16414
R1135 VDD1.n193 VDD1.n192 1.16414
R1136 VDD1.n216 VDD1.t1 1.04867
R1137 VDD1.n216 VDD1.t7 1.04867
R1138 VDD1.n105 VDD1.t4 1.04867
R1139 VDD1.n105 VDD1.t9 1.04867
R1140 VDD1.n214 VDD1.t6 1.04867
R1141 VDD1.n214 VDD1.t2 1.04867
R1142 VDD1.n212 VDD1.t8 1.04867
R1143 VDD1.n212 VDD1.t5 1.04867
R1144 VDD1 VDD1.n106 0.946621
R1145 VDD1.n215 VDD1.n213 0.833085
R1146 VDD1.n82 VDD1.n10 0.388379
R1147 VDD1.n81 VDD1.n80 0.388379
R1148 VDD1.n37 VDD1.n36 0.388379
R1149 VDD1.n143 VDD1.n142 0.388379
R1150 VDD1.n188 VDD1.n187 0.388379
R1151 VDD1.n189 VDD1.n117 0.388379
R1152 VDD1.n103 VDD1.n1 0.155672
R1153 VDD1.n96 VDD1.n1 0.155672
R1154 VDD1.n96 VDD1.n95 0.155672
R1155 VDD1.n95 VDD1.n5 0.155672
R1156 VDD1.n88 VDD1.n5 0.155672
R1157 VDD1.n88 VDD1.n87 0.155672
R1158 VDD1.n87 VDD1.n9 0.155672
R1159 VDD1.n79 VDD1.n9 0.155672
R1160 VDD1.n79 VDD1.n78 0.155672
R1161 VDD1.n78 VDD1.n13 0.155672
R1162 VDD1.n71 VDD1.n13 0.155672
R1163 VDD1.n71 VDD1.n70 0.155672
R1164 VDD1.n70 VDD1.n18 0.155672
R1165 VDD1.n63 VDD1.n18 0.155672
R1166 VDD1.n63 VDD1.n62 0.155672
R1167 VDD1.n62 VDD1.n22 0.155672
R1168 VDD1.n55 VDD1.n22 0.155672
R1169 VDD1.n55 VDD1.n54 0.155672
R1170 VDD1.n54 VDD1.n26 0.155672
R1171 VDD1.n47 VDD1.n26 0.155672
R1172 VDD1.n47 VDD1.n46 0.155672
R1173 VDD1.n46 VDD1.n30 0.155672
R1174 VDD1.n39 VDD1.n30 0.155672
R1175 VDD1.n39 VDD1.n38 0.155672
R1176 VDD1.n145 VDD1.n144 0.155672
R1177 VDD1.n145 VDD1.n136 0.155672
R1178 VDD1.n152 VDD1.n136 0.155672
R1179 VDD1.n153 VDD1.n152 0.155672
R1180 VDD1.n153 VDD1.n132 0.155672
R1181 VDD1.n160 VDD1.n132 0.155672
R1182 VDD1.n161 VDD1.n160 0.155672
R1183 VDD1.n161 VDD1.n128 0.155672
R1184 VDD1.n168 VDD1.n128 0.155672
R1185 VDD1.n169 VDD1.n168 0.155672
R1186 VDD1.n169 VDD1.n124 0.155672
R1187 VDD1.n176 VDD1.n124 0.155672
R1188 VDD1.n177 VDD1.n176 0.155672
R1189 VDD1.n177 VDD1.n120 0.155672
R1190 VDD1.n185 VDD1.n120 0.155672
R1191 VDD1.n186 VDD1.n185 0.155672
R1192 VDD1.n186 VDD1.n116 0.155672
R1193 VDD1.n194 VDD1.n116 0.155672
R1194 VDD1.n195 VDD1.n194 0.155672
R1195 VDD1.n195 VDD1.n112 0.155672
R1196 VDD1.n202 VDD1.n112 0.155672
R1197 VDD1.n203 VDD1.n202 0.155672
R1198 VDD1.n203 VDD1.n108 0.155672
R1199 VDD1.n210 VDD1.n108 0.155672
R1200 B.n1327 B.n1326 585
R1201 B.n1328 B.n1327 585
R1202 B.n482 B.n213 585
R1203 B.n481 B.n480 585
R1204 B.n479 B.n478 585
R1205 B.n477 B.n476 585
R1206 B.n475 B.n474 585
R1207 B.n473 B.n472 585
R1208 B.n471 B.n470 585
R1209 B.n469 B.n468 585
R1210 B.n467 B.n466 585
R1211 B.n465 B.n464 585
R1212 B.n463 B.n462 585
R1213 B.n461 B.n460 585
R1214 B.n459 B.n458 585
R1215 B.n457 B.n456 585
R1216 B.n455 B.n454 585
R1217 B.n453 B.n452 585
R1218 B.n451 B.n450 585
R1219 B.n449 B.n448 585
R1220 B.n447 B.n446 585
R1221 B.n445 B.n444 585
R1222 B.n443 B.n442 585
R1223 B.n441 B.n440 585
R1224 B.n439 B.n438 585
R1225 B.n437 B.n436 585
R1226 B.n435 B.n434 585
R1227 B.n433 B.n432 585
R1228 B.n431 B.n430 585
R1229 B.n429 B.n428 585
R1230 B.n427 B.n426 585
R1231 B.n425 B.n424 585
R1232 B.n423 B.n422 585
R1233 B.n421 B.n420 585
R1234 B.n419 B.n418 585
R1235 B.n417 B.n416 585
R1236 B.n415 B.n414 585
R1237 B.n413 B.n412 585
R1238 B.n411 B.n410 585
R1239 B.n409 B.n408 585
R1240 B.n407 B.n406 585
R1241 B.n405 B.n404 585
R1242 B.n403 B.n402 585
R1243 B.n401 B.n400 585
R1244 B.n399 B.n398 585
R1245 B.n397 B.n396 585
R1246 B.n395 B.n394 585
R1247 B.n393 B.n392 585
R1248 B.n391 B.n390 585
R1249 B.n389 B.n388 585
R1250 B.n387 B.n386 585
R1251 B.n385 B.n384 585
R1252 B.n383 B.n382 585
R1253 B.n381 B.n380 585
R1254 B.n379 B.n378 585
R1255 B.n377 B.n376 585
R1256 B.n375 B.n374 585
R1257 B.n373 B.n372 585
R1258 B.n371 B.n370 585
R1259 B.n369 B.n368 585
R1260 B.n367 B.n366 585
R1261 B.n365 B.n364 585
R1262 B.n363 B.n362 585
R1263 B.n360 B.n359 585
R1264 B.n358 B.n357 585
R1265 B.n356 B.n355 585
R1266 B.n354 B.n353 585
R1267 B.n352 B.n351 585
R1268 B.n350 B.n349 585
R1269 B.n348 B.n347 585
R1270 B.n346 B.n345 585
R1271 B.n344 B.n343 585
R1272 B.n342 B.n341 585
R1273 B.n340 B.n339 585
R1274 B.n338 B.n337 585
R1275 B.n336 B.n335 585
R1276 B.n334 B.n333 585
R1277 B.n332 B.n331 585
R1278 B.n330 B.n329 585
R1279 B.n328 B.n327 585
R1280 B.n326 B.n325 585
R1281 B.n324 B.n323 585
R1282 B.n322 B.n321 585
R1283 B.n320 B.n319 585
R1284 B.n318 B.n317 585
R1285 B.n316 B.n315 585
R1286 B.n314 B.n313 585
R1287 B.n312 B.n311 585
R1288 B.n310 B.n309 585
R1289 B.n308 B.n307 585
R1290 B.n306 B.n305 585
R1291 B.n304 B.n303 585
R1292 B.n302 B.n301 585
R1293 B.n300 B.n299 585
R1294 B.n298 B.n297 585
R1295 B.n296 B.n295 585
R1296 B.n294 B.n293 585
R1297 B.n292 B.n291 585
R1298 B.n290 B.n289 585
R1299 B.n288 B.n287 585
R1300 B.n286 B.n285 585
R1301 B.n284 B.n283 585
R1302 B.n282 B.n281 585
R1303 B.n280 B.n279 585
R1304 B.n278 B.n277 585
R1305 B.n276 B.n275 585
R1306 B.n274 B.n273 585
R1307 B.n272 B.n271 585
R1308 B.n270 B.n269 585
R1309 B.n268 B.n267 585
R1310 B.n266 B.n265 585
R1311 B.n264 B.n263 585
R1312 B.n262 B.n261 585
R1313 B.n260 B.n259 585
R1314 B.n258 B.n257 585
R1315 B.n256 B.n255 585
R1316 B.n254 B.n253 585
R1317 B.n252 B.n251 585
R1318 B.n250 B.n249 585
R1319 B.n248 B.n247 585
R1320 B.n246 B.n245 585
R1321 B.n244 B.n243 585
R1322 B.n242 B.n241 585
R1323 B.n240 B.n239 585
R1324 B.n238 B.n237 585
R1325 B.n236 B.n235 585
R1326 B.n234 B.n233 585
R1327 B.n232 B.n231 585
R1328 B.n230 B.n229 585
R1329 B.n228 B.n227 585
R1330 B.n226 B.n225 585
R1331 B.n224 B.n223 585
R1332 B.n222 B.n221 585
R1333 B.n220 B.n219 585
R1334 B.n1325 B.n146 585
R1335 B.n1329 B.n146 585
R1336 B.n1324 B.n145 585
R1337 B.n1330 B.n145 585
R1338 B.n1323 B.n1322 585
R1339 B.n1322 B.n141 585
R1340 B.n1321 B.n140 585
R1341 B.n1336 B.n140 585
R1342 B.n1320 B.n139 585
R1343 B.n1337 B.n139 585
R1344 B.n1319 B.n138 585
R1345 B.n1338 B.n138 585
R1346 B.n1318 B.n1317 585
R1347 B.n1317 B.n134 585
R1348 B.n1316 B.n133 585
R1349 B.n1344 B.n133 585
R1350 B.n1315 B.n132 585
R1351 B.n1345 B.n132 585
R1352 B.n1314 B.n131 585
R1353 B.n1346 B.n131 585
R1354 B.n1313 B.n1312 585
R1355 B.n1312 B.n127 585
R1356 B.n1311 B.n126 585
R1357 B.n1352 B.n126 585
R1358 B.n1310 B.n125 585
R1359 B.n1353 B.n125 585
R1360 B.n1309 B.n124 585
R1361 B.n1354 B.n124 585
R1362 B.n1308 B.n1307 585
R1363 B.n1307 B.n120 585
R1364 B.n1306 B.n119 585
R1365 B.n1360 B.n119 585
R1366 B.n1305 B.n118 585
R1367 B.n1361 B.n118 585
R1368 B.n1304 B.n117 585
R1369 B.n1362 B.n117 585
R1370 B.n1303 B.n1302 585
R1371 B.n1302 B.n113 585
R1372 B.n1301 B.n112 585
R1373 B.n1368 B.n112 585
R1374 B.n1300 B.n111 585
R1375 B.n1369 B.n111 585
R1376 B.n1299 B.n110 585
R1377 B.n1370 B.n110 585
R1378 B.n1298 B.n1297 585
R1379 B.n1297 B.n106 585
R1380 B.n1296 B.n105 585
R1381 B.n1376 B.n105 585
R1382 B.n1295 B.n104 585
R1383 B.n1377 B.n104 585
R1384 B.n1294 B.n103 585
R1385 B.n1378 B.n103 585
R1386 B.n1293 B.n1292 585
R1387 B.n1292 B.n99 585
R1388 B.n1291 B.n98 585
R1389 B.n1384 B.n98 585
R1390 B.n1290 B.n97 585
R1391 B.n1385 B.n97 585
R1392 B.n1289 B.n96 585
R1393 B.n1386 B.n96 585
R1394 B.n1288 B.n1287 585
R1395 B.n1287 B.n92 585
R1396 B.n1286 B.n91 585
R1397 B.n1392 B.n91 585
R1398 B.n1285 B.n90 585
R1399 B.n1393 B.n90 585
R1400 B.n1284 B.n89 585
R1401 B.n1394 B.n89 585
R1402 B.n1283 B.n1282 585
R1403 B.n1282 B.n85 585
R1404 B.n1281 B.n84 585
R1405 B.n1400 B.n84 585
R1406 B.n1280 B.n83 585
R1407 B.n1401 B.n83 585
R1408 B.n1279 B.n82 585
R1409 B.n1402 B.n82 585
R1410 B.n1278 B.n1277 585
R1411 B.n1277 B.n78 585
R1412 B.n1276 B.n77 585
R1413 B.n1408 B.n77 585
R1414 B.n1275 B.n76 585
R1415 B.n1409 B.n76 585
R1416 B.n1274 B.n75 585
R1417 B.n1410 B.n75 585
R1418 B.n1273 B.n1272 585
R1419 B.n1272 B.n71 585
R1420 B.n1271 B.n70 585
R1421 B.n1416 B.n70 585
R1422 B.n1270 B.n69 585
R1423 B.n1417 B.n69 585
R1424 B.n1269 B.n68 585
R1425 B.n1418 B.n68 585
R1426 B.n1268 B.n1267 585
R1427 B.n1267 B.n64 585
R1428 B.n1266 B.n63 585
R1429 B.n1424 B.n63 585
R1430 B.n1265 B.n62 585
R1431 B.n1425 B.n62 585
R1432 B.n1264 B.n61 585
R1433 B.n1426 B.n61 585
R1434 B.n1263 B.n1262 585
R1435 B.n1262 B.n57 585
R1436 B.n1261 B.n56 585
R1437 B.n1432 B.n56 585
R1438 B.n1260 B.n55 585
R1439 B.n1433 B.n55 585
R1440 B.n1259 B.n54 585
R1441 B.n1434 B.n54 585
R1442 B.n1258 B.n1257 585
R1443 B.n1257 B.n50 585
R1444 B.n1256 B.n49 585
R1445 B.n1440 B.n49 585
R1446 B.n1255 B.n48 585
R1447 B.n1441 B.n48 585
R1448 B.n1254 B.n47 585
R1449 B.n1442 B.n47 585
R1450 B.n1253 B.n1252 585
R1451 B.n1252 B.n43 585
R1452 B.n1251 B.n42 585
R1453 B.n1448 B.n42 585
R1454 B.n1250 B.n41 585
R1455 B.n1449 B.n41 585
R1456 B.n1249 B.n40 585
R1457 B.n1450 B.n40 585
R1458 B.n1248 B.n1247 585
R1459 B.n1247 B.n36 585
R1460 B.n1246 B.n35 585
R1461 B.n1456 B.n35 585
R1462 B.n1245 B.n34 585
R1463 B.n1457 B.n34 585
R1464 B.n1244 B.n33 585
R1465 B.n1458 B.n33 585
R1466 B.n1243 B.n1242 585
R1467 B.n1242 B.n29 585
R1468 B.n1241 B.n28 585
R1469 B.n1464 B.n28 585
R1470 B.n1240 B.n27 585
R1471 B.n1465 B.n27 585
R1472 B.n1239 B.n26 585
R1473 B.n1466 B.n26 585
R1474 B.n1238 B.n1237 585
R1475 B.n1237 B.n22 585
R1476 B.n1236 B.n21 585
R1477 B.n1472 B.n21 585
R1478 B.n1235 B.n20 585
R1479 B.n1473 B.n20 585
R1480 B.n1234 B.n19 585
R1481 B.n1474 B.n19 585
R1482 B.n1233 B.n1232 585
R1483 B.n1232 B.n15 585
R1484 B.n1231 B.n14 585
R1485 B.n1480 B.n14 585
R1486 B.n1230 B.n13 585
R1487 B.n1481 B.n13 585
R1488 B.n1229 B.n12 585
R1489 B.n1482 B.n12 585
R1490 B.n1228 B.n1227 585
R1491 B.n1227 B.n8 585
R1492 B.n1226 B.n7 585
R1493 B.n1488 B.n7 585
R1494 B.n1225 B.n6 585
R1495 B.n1489 B.n6 585
R1496 B.n1224 B.n5 585
R1497 B.n1490 B.n5 585
R1498 B.n1223 B.n1222 585
R1499 B.n1222 B.n4 585
R1500 B.n1221 B.n483 585
R1501 B.n1221 B.n1220 585
R1502 B.n1211 B.n484 585
R1503 B.n485 B.n484 585
R1504 B.n1213 B.n1212 585
R1505 B.n1214 B.n1213 585
R1506 B.n1210 B.n490 585
R1507 B.n490 B.n489 585
R1508 B.n1209 B.n1208 585
R1509 B.n1208 B.n1207 585
R1510 B.n492 B.n491 585
R1511 B.n493 B.n492 585
R1512 B.n1200 B.n1199 585
R1513 B.n1201 B.n1200 585
R1514 B.n1198 B.n498 585
R1515 B.n498 B.n497 585
R1516 B.n1197 B.n1196 585
R1517 B.n1196 B.n1195 585
R1518 B.n500 B.n499 585
R1519 B.n501 B.n500 585
R1520 B.n1188 B.n1187 585
R1521 B.n1189 B.n1188 585
R1522 B.n1186 B.n506 585
R1523 B.n506 B.n505 585
R1524 B.n1185 B.n1184 585
R1525 B.n1184 B.n1183 585
R1526 B.n508 B.n507 585
R1527 B.n509 B.n508 585
R1528 B.n1176 B.n1175 585
R1529 B.n1177 B.n1176 585
R1530 B.n1174 B.n514 585
R1531 B.n514 B.n513 585
R1532 B.n1173 B.n1172 585
R1533 B.n1172 B.n1171 585
R1534 B.n516 B.n515 585
R1535 B.n517 B.n516 585
R1536 B.n1164 B.n1163 585
R1537 B.n1165 B.n1164 585
R1538 B.n1162 B.n522 585
R1539 B.n522 B.n521 585
R1540 B.n1161 B.n1160 585
R1541 B.n1160 B.n1159 585
R1542 B.n524 B.n523 585
R1543 B.n525 B.n524 585
R1544 B.n1152 B.n1151 585
R1545 B.n1153 B.n1152 585
R1546 B.n1150 B.n530 585
R1547 B.n530 B.n529 585
R1548 B.n1149 B.n1148 585
R1549 B.n1148 B.n1147 585
R1550 B.n532 B.n531 585
R1551 B.n533 B.n532 585
R1552 B.n1140 B.n1139 585
R1553 B.n1141 B.n1140 585
R1554 B.n1138 B.n538 585
R1555 B.n538 B.n537 585
R1556 B.n1137 B.n1136 585
R1557 B.n1136 B.n1135 585
R1558 B.n540 B.n539 585
R1559 B.n541 B.n540 585
R1560 B.n1128 B.n1127 585
R1561 B.n1129 B.n1128 585
R1562 B.n1126 B.n546 585
R1563 B.n546 B.n545 585
R1564 B.n1125 B.n1124 585
R1565 B.n1124 B.n1123 585
R1566 B.n548 B.n547 585
R1567 B.n549 B.n548 585
R1568 B.n1116 B.n1115 585
R1569 B.n1117 B.n1116 585
R1570 B.n1114 B.n554 585
R1571 B.n554 B.n553 585
R1572 B.n1113 B.n1112 585
R1573 B.n1112 B.n1111 585
R1574 B.n556 B.n555 585
R1575 B.n557 B.n556 585
R1576 B.n1104 B.n1103 585
R1577 B.n1105 B.n1104 585
R1578 B.n1102 B.n562 585
R1579 B.n562 B.n561 585
R1580 B.n1101 B.n1100 585
R1581 B.n1100 B.n1099 585
R1582 B.n564 B.n563 585
R1583 B.n565 B.n564 585
R1584 B.n1092 B.n1091 585
R1585 B.n1093 B.n1092 585
R1586 B.n1090 B.n569 585
R1587 B.n573 B.n569 585
R1588 B.n1089 B.n1088 585
R1589 B.n1088 B.n1087 585
R1590 B.n571 B.n570 585
R1591 B.n572 B.n571 585
R1592 B.n1080 B.n1079 585
R1593 B.n1081 B.n1080 585
R1594 B.n1078 B.n578 585
R1595 B.n578 B.n577 585
R1596 B.n1077 B.n1076 585
R1597 B.n1076 B.n1075 585
R1598 B.n580 B.n579 585
R1599 B.n581 B.n580 585
R1600 B.n1068 B.n1067 585
R1601 B.n1069 B.n1068 585
R1602 B.n1066 B.n586 585
R1603 B.n586 B.n585 585
R1604 B.n1065 B.n1064 585
R1605 B.n1064 B.n1063 585
R1606 B.n588 B.n587 585
R1607 B.n589 B.n588 585
R1608 B.n1056 B.n1055 585
R1609 B.n1057 B.n1056 585
R1610 B.n1054 B.n593 585
R1611 B.n597 B.n593 585
R1612 B.n1053 B.n1052 585
R1613 B.n1052 B.n1051 585
R1614 B.n595 B.n594 585
R1615 B.n596 B.n595 585
R1616 B.n1044 B.n1043 585
R1617 B.n1045 B.n1044 585
R1618 B.n1042 B.n602 585
R1619 B.n602 B.n601 585
R1620 B.n1041 B.n1040 585
R1621 B.n1040 B.n1039 585
R1622 B.n604 B.n603 585
R1623 B.n605 B.n604 585
R1624 B.n1032 B.n1031 585
R1625 B.n1033 B.n1032 585
R1626 B.n1030 B.n610 585
R1627 B.n610 B.n609 585
R1628 B.n1029 B.n1028 585
R1629 B.n1028 B.n1027 585
R1630 B.n612 B.n611 585
R1631 B.n613 B.n612 585
R1632 B.n1020 B.n1019 585
R1633 B.n1021 B.n1020 585
R1634 B.n1018 B.n618 585
R1635 B.n618 B.n617 585
R1636 B.n1017 B.n1016 585
R1637 B.n1016 B.n1015 585
R1638 B.n620 B.n619 585
R1639 B.n621 B.n620 585
R1640 B.n1008 B.n1007 585
R1641 B.n1009 B.n1008 585
R1642 B.n1006 B.n626 585
R1643 B.n626 B.n625 585
R1644 B.n1005 B.n1004 585
R1645 B.n1004 B.n1003 585
R1646 B.n628 B.n627 585
R1647 B.n629 B.n628 585
R1648 B.n996 B.n995 585
R1649 B.n997 B.n996 585
R1650 B.n994 B.n634 585
R1651 B.n634 B.n633 585
R1652 B.n993 B.n992 585
R1653 B.n992 B.n991 585
R1654 B.n636 B.n635 585
R1655 B.n637 B.n636 585
R1656 B.n984 B.n983 585
R1657 B.n985 B.n984 585
R1658 B.n982 B.n642 585
R1659 B.n642 B.n641 585
R1660 B.n976 B.n975 585
R1661 B.n974 B.n710 585
R1662 B.n973 B.n709 585
R1663 B.n978 B.n709 585
R1664 B.n972 B.n971 585
R1665 B.n970 B.n969 585
R1666 B.n968 B.n967 585
R1667 B.n966 B.n965 585
R1668 B.n964 B.n963 585
R1669 B.n962 B.n961 585
R1670 B.n960 B.n959 585
R1671 B.n958 B.n957 585
R1672 B.n956 B.n955 585
R1673 B.n954 B.n953 585
R1674 B.n952 B.n951 585
R1675 B.n950 B.n949 585
R1676 B.n948 B.n947 585
R1677 B.n946 B.n945 585
R1678 B.n944 B.n943 585
R1679 B.n942 B.n941 585
R1680 B.n940 B.n939 585
R1681 B.n938 B.n937 585
R1682 B.n936 B.n935 585
R1683 B.n934 B.n933 585
R1684 B.n932 B.n931 585
R1685 B.n930 B.n929 585
R1686 B.n928 B.n927 585
R1687 B.n926 B.n925 585
R1688 B.n924 B.n923 585
R1689 B.n922 B.n921 585
R1690 B.n920 B.n919 585
R1691 B.n918 B.n917 585
R1692 B.n916 B.n915 585
R1693 B.n914 B.n913 585
R1694 B.n912 B.n911 585
R1695 B.n910 B.n909 585
R1696 B.n908 B.n907 585
R1697 B.n906 B.n905 585
R1698 B.n904 B.n903 585
R1699 B.n902 B.n901 585
R1700 B.n900 B.n899 585
R1701 B.n898 B.n897 585
R1702 B.n896 B.n895 585
R1703 B.n894 B.n893 585
R1704 B.n892 B.n891 585
R1705 B.n890 B.n889 585
R1706 B.n888 B.n887 585
R1707 B.n886 B.n885 585
R1708 B.n884 B.n883 585
R1709 B.n882 B.n881 585
R1710 B.n880 B.n879 585
R1711 B.n878 B.n877 585
R1712 B.n876 B.n875 585
R1713 B.n874 B.n873 585
R1714 B.n872 B.n871 585
R1715 B.n870 B.n869 585
R1716 B.n868 B.n867 585
R1717 B.n866 B.n865 585
R1718 B.n864 B.n863 585
R1719 B.n862 B.n861 585
R1720 B.n860 B.n859 585
R1721 B.n858 B.n857 585
R1722 B.n856 B.n855 585
R1723 B.n853 B.n852 585
R1724 B.n851 B.n850 585
R1725 B.n849 B.n848 585
R1726 B.n847 B.n846 585
R1727 B.n845 B.n844 585
R1728 B.n843 B.n842 585
R1729 B.n841 B.n840 585
R1730 B.n839 B.n838 585
R1731 B.n837 B.n836 585
R1732 B.n835 B.n834 585
R1733 B.n833 B.n832 585
R1734 B.n831 B.n830 585
R1735 B.n829 B.n828 585
R1736 B.n827 B.n826 585
R1737 B.n825 B.n824 585
R1738 B.n823 B.n822 585
R1739 B.n821 B.n820 585
R1740 B.n819 B.n818 585
R1741 B.n817 B.n816 585
R1742 B.n815 B.n814 585
R1743 B.n813 B.n812 585
R1744 B.n811 B.n810 585
R1745 B.n809 B.n808 585
R1746 B.n807 B.n806 585
R1747 B.n805 B.n804 585
R1748 B.n803 B.n802 585
R1749 B.n801 B.n800 585
R1750 B.n799 B.n798 585
R1751 B.n797 B.n796 585
R1752 B.n795 B.n794 585
R1753 B.n793 B.n792 585
R1754 B.n791 B.n790 585
R1755 B.n789 B.n788 585
R1756 B.n787 B.n786 585
R1757 B.n785 B.n784 585
R1758 B.n783 B.n782 585
R1759 B.n781 B.n780 585
R1760 B.n779 B.n778 585
R1761 B.n777 B.n776 585
R1762 B.n775 B.n774 585
R1763 B.n773 B.n772 585
R1764 B.n771 B.n770 585
R1765 B.n769 B.n768 585
R1766 B.n767 B.n766 585
R1767 B.n765 B.n764 585
R1768 B.n763 B.n762 585
R1769 B.n761 B.n760 585
R1770 B.n759 B.n758 585
R1771 B.n757 B.n756 585
R1772 B.n755 B.n754 585
R1773 B.n753 B.n752 585
R1774 B.n751 B.n750 585
R1775 B.n749 B.n748 585
R1776 B.n747 B.n746 585
R1777 B.n745 B.n744 585
R1778 B.n743 B.n742 585
R1779 B.n741 B.n740 585
R1780 B.n739 B.n738 585
R1781 B.n737 B.n736 585
R1782 B.n735 B.n734 585
R1783 B.n733 B.n732 585
R1784 B.n731 B.n730 585
R1785 B.n729 B.n728 585
R1786 B.n727 B.n726 585
R1787 B.n725 B.n724 585
R1788 B.n723 B.n722 585
R1789 B.n721 B.n720 585
R1790 B.n719 B.n718 585
R1791 B.n717 B.n716 585
R1792 B.n644 B.n643 585
R1793 B.n981 B.n980 585
R1794 B.n640 B.n639 585
R1795 B.n641 B.n640 585
R1796 B.n987 B.n986 585
R1797 B.n986 B.n985 585
R1798 B.n988 B.n638 585
R1799 B.n638 B.n637 585
R1800 B.n990 B.n989 585
R1801 B.n991 B.n990 585
R1802 B.n632 B.n631 585
R1803 B.n633 B.n632 585
R1804 B.n999 B.n998 585
R1805 B.n998 B.n997 585
R1806 B.n1000 B.n630 585
R1807 B.n630 B.n629 585
R1808 B.n1002 B.n1001 585
R1809 B.n1003 B.n1002 585
R1810 B.n624 B.n623 585
R1811 B.n625 B.n624 585
R1812 B.n1011 B.n1010 585
R1813 B.n1010 B.n1009 585
R1814 B.n1012 B.n622 585
R1815 B.n622 B.n621 585
R1816 B.n1014 B.n1013 585
R1817 B.n1015 B.n1014 585
R1818 B.n616 B.n615 585
R1819 B.n617 B.n616 585
R1820 B.n1023 B.n1022 585
R1821 B.n1022 B.n1021 585
R1822 B.n1024 B.n614 585
R1823 B.n614 B.n613 585
R1824 B.n1026 B.n1025 585
R1825 B.n1027 B.n1026 585
R1826 B.n608 B.n607 585
R1827 B.n609 B.n608 585
R1828 B.n1035 B.n1034 585
R1829 B.n1034 B.n1033 585
R1830 B.n1036 B.n606 585
R1831 B.n606 B.n605 585
R1832 B.n1038 B.n1037 585
R1833 B.n1039 B.n1038 585
R1834 B.n600 B.n599 585
R1835 B.n601 B.n600 585
R1836 B.n1047 B.n1046 585
R1837 B.n1046 B.n1045 585
R1838 B.n1048 B.n598 585
R1839 B.n598 B.n596 585
R1840 B.n1050 B.n1049 585
R1841 B.n1051 B.n1050 585
R1842 B.n592 B.n591 585
R1843 B.n597 B.n592 585
R1844 B.n1059 B.n1058 585
R1845 B.n1058 B.n1057 585
R1846 B.n1060 B.n590 585
R1847 B.n590 B.n589 585
R1848 B.n1062 B.n1061 585
R1849 B.n1063 B.n1062 585
R1850 B.n584 B.n583 585
R1851 B.n585 B.n584 585
R1852 B.n1071 B.n1070 585
R1853 B.n1070 B.n1069 585
R1854 B.n1072 B.n582 585
R1855 B.n582 B.n581 585
R1856 B.n1074 B.n1073 585
R1857 B.n1075 B.n1074 585
R1858 B.n576 B.n575 585
R1859 B.n577 B.n576 585
R1860 B.n1083 B.n1082 585
R1861 B.n1082 B.n1081 585
R1862 B.n1084 B.n574 585
R1863 B.n574 B.n572 585
R1864 B.n1086 B.n1085 585
R1865 B.n1087 B.n1086 585
R1866 B.n568 B.n567 585
R1867 B.n573 B.n568 585
R1868 B.n1095 B.n1094 585
R1869 B.n1094 B.n1093 585
R1870 B.n1096 B.n566 585
R1871 B.n566 B.n565 585
R1872 B.n1098 B.n1097 585
R1873 B.n1099 B.n1098 585
R1874 B.n560 B.n559 585
R1875 B.n561 B.n560 585
R1876 B.n1107 B.n1106 585
R1877 B.n1106 B.n1105 585
R1878 B.n1108 B.n558 585
R1879 B.n558 B.n557 585
R1880 B.n1110 B.n1109 585
R1881 B.n1111 B.n1110 585
R1882 B.n552 B.n551 585
R1883 B.n553 B.n552 585
R1884 B.n1119 B.n1118 585
R1885 B.n1118 B.n1117 585
R1886 B.n1120 B.n550 585
R1887 B.n550 B.n549 585
R1888 B.n1122 B.n1121 585
R1889 B.n1123 B.n1122 585
R1890 B.n544 B.n543 585
R1891 B.n545 B.n544 585
R1892 B.n1131 B.n1130 585
R1893 B.n1130 B.n1129 585
R1894 B.n1132 B.n542 585
R1895 B.n542 B.n541 585
R1896 B.n1134 B.n1133 585
R1897 B.n1135 B.n1134 585
R1898 B.n536 B.n535 585
R1899 B.n537 B.n536 585
R1900 B.n1143 B.n1142 585
R1901 B.n1142 B.n1141 585
R1902 B.n1144 B.n534 585
R1903 B.n534 B.n533 585
R1904 B.n1146 B.n1145 585
R1905 B.n1147 B.n1146 585
R1906 B.n528 B.n527 585
R1907 B.n529 B.n528 585
R1908 B.n1155 B.n1154 585
R1909 B.n1154 B.n1153 585
R1910 B.n1156 B.n526 585
R1911 B.n526 B.n525 585
R1912 B.n1158 B.n1157 585
R1913 B.n1159 B.n1158 585
R1914 B.n520 B.n519 585
R1915 B.n521 B.n520 585
R1916 B.n1167 B.n1166 585
R1917 B.n1166 B.n1165 585
R1918 B.n1168 B.n518 585
R1919 B.n518 B.n517 585
R1920 B.n1170 B.n1169 585
R1921 B.n1171 B.n1170 585
R1922 B.n512 B.n511 585
R1923 B.n513 B.n512 585
R1924 B.n1179 B.n1178 585
R1925 B.n1178 B.n1177 585
R1926 B.n1180 B.n510 585
R1927 B.n510 B.n509 585
R1928 B.n1182 B.n1181 585
R1929 B.n1183 B.n1182 585
R1930 B.n504 B.n503 585
R1931 B.n505 B.n504 585
R1932 B.n1191 B.n1190 585
R1933 B.n1190 B.n1189 585
R1934 B.n1192 B.n502 585
R1935 B.n502 B.n501 585
R1936 B.n1194 B.n1193 585
R1937 B.n1195 B.n1194 585
R1938 B.n496 B.n495 585
R1939 B.n497 B.n496 585
R1940 B.n1203 B.n1202 585
R1941 B.n1202 B.n1201 585
R1942 B.n1204 B.n494 585
R1943 B.n494 B.n493 585
R1944 B.n1206 B.n1205 585
R1945 B.n1207 B.n1206 585
R1946 B.n488 B.n487 585
R1947 B.n489 B.n488 585
R1948 B.n1216 B.n1215 585
R1949 B.n1215 B.n1214 585
R1950 B.n1217 B.n486 585
R1951 B.n486 B.n485 585
R1952 B.n1219 B.n1218 585
R1953 B.n1220 B.n1219 585
R1954 B.n2 B.n0 585
R1955 B.n4 B.n2 585
R1956 B.n3 B.n1 585
R1957 B.n1489 B.n3 585
R1958 B.n1487 B.n1486 585
R1959 B.n1488 B.n1487 585
R1960 B.n1485 B.n9 585
R1961 B.n9 B.n8 585
R1962 B.n1484 B.n1483 585
R1963 B.n1483 B.n1482 585
R1964 B.n11 B.n10 585
R1965 B.n1481 B.n11 585
R1966 B.n1479 B.n1478 585
R1967 B.n1480 B.n1479 585
R1968 B.n1477 B.n16 585
R1969 B.n16 B.n15 585
R1970 B.n1476 B.n1475 585
R1971 B.n1475 B.n1474 585
R1972 B.n18 B.n17 585
R1973 B.n1473 B.n18 585
R1974 B.n1471 B.n1470 585
R1975 B.n1472 B.n1471 585
R1976 B.n1469 B.n23 585
R1977 B.n23 B.n22 585
R1978 B.n1468 B.n1467 585
R1979 B.n1467 B.n1466 585
R1980 B.n25 B.n24 585
R1981 B.n1465 B.n25 585
R1982 B.n1463 B.n1462 585
R1983 B.n1464 B.n1463 585
R1984 B.n1461 B.n30 585
R1985 B.n30 B.n29 585
R1986 B.n1460 B.n1459 585
R1987 B.n1459 B.n1458 585
R1988 B.n32 B.n31 585
R1989 B.n1457 B.n32 585
R1990 B.n1455 B.n1454 585
R1991 B.n1456 B.n1455 585
R1992 B.n1453 B.n37 585
R1993 B.n37 B.n36 585
R1994 B.n1452 B.n1451 585
R1995 B.n1451 B.n1450 585
R1996 B.n39 B.n38 585
R1997 B.n1449 B.n39 585
R1998 B.n1447 B.n1446 585
R1999 B.n1448 B.n1447 585
R2000 B.n1445 B.n44 585
R2001 B.n44 B.n43 585
R2002 B.n1444 B.n1443 585
R2003 B.n1443 B.n1442 585
R2004 B.n46 B.n45 585
R2005 B.n1441 B.n46 585
R2006 B.n1439 B.n1438 585
R2007 B.n1440 B.n1439 585
R2008 B.n1437 B.n51 585
R2009 B.n51 B.n50 585
R2010 B.n1436 B.n1435 585
R2011 B.n1435 B.n1434 585
R2012 B.n53 B.n52 585
R2013 B.n1433 B.n53 585
R2014 B.n1431 B.n1430 585
R2015 B.n1432 B.n1431 585
R2016 B.n1429 B.n58 585
R2017 B.n58 B.n57 585
R2018 B.n1428 B.n1427 585
R2019 B.n1427 B.n1426 585
R2020 B.n60 B.n59 585
R2021 B.n1425 B.n60 585
R2022 B.n1423 B.n1422 585
R2023 B.n1424 B.n1423 585
R2024 B.n1421 B.n65 585
R2025 B.n65 B.n64 585
R2026 B.n1420 B.n1419 585
R2027 B.n1419 B.n1418 585
R2028 B.n67 B.n66 585
R2029 B.n1417 B.n67 585
R2030 B.n1415 B.n1414 585
R2031 B.n1416 B.n1415 585
R2032 B.n1413 B.n72 585
R2033 B.n72 B.n71 585
R2034 B.n1412 B.n1411 585
R2035 B.n1411 B.n1410 585
R2036 B.n74 B.n73 585
R2037 B.n1409 B.n74 585
R2038 B.n1407 B.n1406 585
R2039 B.n1408 B.n1407 585
R2040 B.n1405 B.n79 585
R2041 B.n79 B.n78 585
R2042 B.n1404 B.n1403 585
R2043 B.n1403 B.n1402 585
R2044 B.n81 B.n80 585
R2045 B.n1401 B.n81 585
R2046 B.n1399 B.n1398 585
R2047 B.n1400 B.n1399 585
R2048 B.n1397 B.n86 585
R2049 B.n86 B.n85 585
R2050 B.n1396 B.n1395 585
R2051 B.n1395 B.n1394 585
R2052 B.n88 B.n87 585
R2053 B.n1393 B.n88 585
R2054 B.n1391 B.n1390 585
R2055 B.n1392 B.n1391 585
R2056 B.n1389 B.n93 585
R2057 B.n93 B.n92 585
R2058 B.n1388 B.n1387 585
R2059 B.n1387 B.n1386 585
R2060 B.n95 B.n94 585
R2061 B.n1385 B.n95 585
R2062 B.n1383 B.n1382 585
R2063 B.n1384 B.n1383 585
R2064 B.n1381 B.n100 585
R2065 B.n100 B.n99 585
R2066 B.n1380 B.n1379 585
R2067 B.n1379 B.n1378 585
R2068 B.n102 B.n101 585
R2069 B.n1377 B.n102 585
R2070 B.n1375 B.n1374 585
R2071 B.n1376 B.n1375 585
R2072 B.n1373 B.n107 585
R2073 B.n107 B.n106 585
R2074 B.n1372 B.n1371 585
R2075 B.n1371 B.n1370 585
R2076 B.n109 B.n108 585
R2077 B.n1369 B.n109 585
R2078 B.n1367 B.n1366 585
R2079 B.n1368 B.n1367 585
R2080 B.n1365 B.n114 585
R2081 B.n114 B.n113 585
R2082 B.n1364 B.n1363 585
R2083 B.n1363 B.n1362 585
R2084 B.n116 B.n115 585
R2085 B.n1361 B.n116 585
R2086 B.n1359 B.n1358 585
R2087 B.n1360 B.n1359 585
R2088 B.n1357 B.n121 585
R2089 B.n121 B.n120 585
R2090 B.n1356 B.n1355 585
R2091 B.n1355 B.n1354 585
R2092 B.n123 B.n122 585
R2093 B.n1353 B.n123 585
R2094 B.n1351 B.n1350 585
R2095 B.n1352 B.n1351 585
R2096 B.n1349 B.n128 585
R2097 B.n128 B.n127 585
R2098 B.n1348 B.n1347 585
R2099 B.n1347 B.n1346 585
R2100 B.n130 B.n129 585
R2101 B.n1345 B.n130 585
R2102 B.n1343 B.n1342 585
R2103 B.n1344 B.n1343 585
R2104 B.n1341 B.n135 585
R2105 B.n135 B.n134 585
R2106 B.n1340 B.n1339 585
R2107 B.n1339 B.n1338 585
R2108 B.n137 B.n136 585
R2109 B.n1337 B.n137 585
R2110 B.n1335 B.n1334 585
R2111 B.n1336 B.n1335 585
R2112 B.n1333 B.n142 585
R2113 B.n142 B.n141 585
R2114 B.n1332 B.n1331 585
R2115 B.n1331 B.n1330 585
R2116 B.n144 B.n143 585
R2117 B.n1329 B.n144 585
R2118 B.n1492 B.n1491 585
R2119 B.n1491 B.n1490 585
R2120 B.n976 B.n640 497.305
R2121 B.n219 B.n144 497.305
R2122 B.n980 B.n642 497.305
R2123 B.n1327 B.n146 497.305
R2124 B.n713 B.t13 480.781
R2125 B.n711 B.t16 480.781
R2126 B.n216 B.t19 480.781
R2127 B.n214 B.t22 480.781
R2128 B.n714 B.t12 400.877
R2129 B.n215 B.t23 400.877
R2130 B.n712 B.t15 400.877
R2131 B.n217 B.t20 400.877
R2132 B.n713 B.t10 329.454
R2133 B.n711 B.t14 329.454
R2134 B.n216 B.t17 329.454
R2135 B.n214 B.t21 329.454
R2136 B.n1328 B.n212 256.663
R2137 B.n1328 B.n211 256.663
R2138 B.n1328 B.n210 256.663
R2139 B.n1328 B.n209 256.663
R2140 B.n1328 B.n208 256.663
R2141 B.n1328 B.n207 256.663
R2142 B.n1328 B.n206 256.663
R2143 B.n1328 B.n205 256.663
R2144 B.n1328 B.n204 256.663
R2145 B.n1328 B.n203 256.663
R2146 B.n1328 B.n202 256.663
R2147 B.n1328 B.n201 256.663
R2148 B.n1328 B.n200 256.663
R2149 B.n1328 B.n199 256.663
R2150 B.n1328 B.n198 256.663
R2151 B.n1328 B.n197 256.663
R2152 B.n1328 B.n196 256.663
R2153 B.n1328 B.n195 256.663
R2154 B.n1328 B.n194 256.663
R2155 B.n1328 B.n193 256.663
R2156 B.n1328 B.n192 256.663
R2157 B.n1328 B.n191 256.663
R2158 B.n1328 B.n190 256.663
R2159 B.n1328 B.n189 256.663
R2160 B.n1328 B.n188 256.663
R2161 B.n1328 B.n187 256.663
R2162 B.n1328 B.n186 256.663
R2163 B.n1328 B.n185 256.663
R2164 B.n1328 B.n184 256.663
R2165 B.n1328 B.n183 256.663
R2166 B.n1328 B.n182 256.663
R2167 B.n1328 B.n181 256.663
R2168 B.n1328 B.n180 256.663
R2169 B.n1328 B.n179 256.663
R2170 B.n1328 B.n178 256.663
R2171 B.n1328 B.n177 256.663
R2172 B.n1328 B.n176 256.663
R2173 B.n1328 B.n175 256.663
R2174 B.n1328 B.n174 256.663
R2175 B.n1328 B.n173 256.663
R2176 B.n1328 B.n172 256.663
R2177 B.n1328 B.n171 256.663
R2178 B.n1328 B.n170 256.663
R2179 B.n1328 B.n169 256.663
R2180 B.n1328 B.n168 256.663
R2181 B.n1328 B.n167 256.663
R2182 B.n1328 B.n166 256.663
R2183 B.n1328 B.n165 256.663
R2184 B.n1328 B.n164 256.663
R2185 B.n1328 B.n163 256.663
R2186 B.n1328 B.n162 256.663
R2187 B.n1328 B.n161 256.663
R2188 B.n1328 B.n160 256.663
R2189 B.n1328 B.n159 256.663
R2190 B.n1328 B.n158 256.663
R2191 B.n1328 B.n157 256.663
R2192 B.n1328 B.n156 256.663
R2193 B.n1328 B.n155 256.663
R2194 B.n1328 B.n154 256.663
R2195 B.n1328 B.n153 256.663
R2196 B.n1328 B.n152 256.663
R2197 B.n1328 B.n151 256.663
R2198 B.n1328 B.n150 256.663
R2199 B.n1328 B.n149 256.663
R2200 B.n1328 B.n148 256.663
R2201 B.n1328 B.n147 256.663
R2202 B.n978 B.n977 256.663
R2203 B.n978 B.n645 256.663
R2204 B.n978 B.n646 256.663
R2205 B.n978 B.n647 256.663
R2206 B.n978 B.n648 256.663
R2207 B.n978 B.n649 256.663
R2208 B.n978 B.n650 256.663
R2209 B.n978 B.n651 256.663
R2210 B.n978 B.n652 256.663
R2211 B.n978 B.n653 256.663
R2212 B.n978 B.n654 256.663
R2213 B.n978 B.n655 256.663
R2214 B.n978 B.n656 256.663
R2215 B.n978 B.n657 256.663
R2216 B.n978 B.n658 256.663
R2217 B.n978 B.n659 256.663
R2218 B.n978 B.n660 256.663
R2219 B.n978 B.n661 256.663
R2220 B.n978 B.n662 256.663
R2221 B.n978 B.n663 256.663
R2222 B.n978 B.n664 256.663
R2223 B.n978 B.n665 256.663
R2224 B.n978 B.n666 256.663
R2225 B.n978 B.n667 256.663
R2226 B.n978 B.n668 256.663
R2227 B.n978 B.n669 256.663
R2228 B.n978 B.n670 256.663
R2229 B.n978 B.n671 256.663
R2230 B.n978 B.n672 256.663
R2231 B.n978 B.n673 256.663
R2232 B.n978 B.n674 256.663
R2233 B.n978 B.n675 256.663
R2234 B.n978 B.n676 256.663
R2235 B.n978 B.n677 256.663
R2236 B.n978 B.n678 256.663
R2237 B.n978 B.n679 256.663
R2238 B.n978 B.n680 256.663
R2239 B.n978 B.n681 256.663
R2240 B.n978 B.n682 256.663
R2241 B.n978 B.n683 256.663
R2242 B.n978 B.n684 256.663
R2243 B.n978 B.n685 256.663
R2244 B.n978 B.n686 256.663
R2245 B.n978 B.n687 256.663
R2246 B.n978 B.n688 256.663
R2247 B.n978 B.n689 256.663
R2248 B.n978 B.n690 256.663
R2249 B.n978 B.n691 256.663
R2250 B.n978 B.n692 256.663
R2251 B.n978 B.n693 256.663
R2252 B.n978 B.n694 256.663
R2253 B.n978 B.n695 256.663
R2254 B.n978 B.n696 256.663
R2255 B.n978 B.n697 256.663
R2256 B.n978 B.n698 256.663
R2257 B.n978 B.n699 256.663
R2258 B.n978 B.n700 256.663
R2259 B.n978 B.n701 256.663
R2260 B.n978 B.n702 256.663
R2261 B.n978 B.n703 256.663
R2262 B.n978 B.n704 256.663
R2263 B.n978 B.n705 256.663
R2264 B.n978 B.n706 256.663
R2265 B.n978 B.n707 256.663
R2266 B.n978 B.n708 256.663
R2267 B.n979 B.n978 256.663
R2268 B.n986 B.n640 163.367
R2269 B.n986 B.n638 163.367
R2270 B.n990 B.n638 163.367
R2271 B.n990 B.n632 163.367
R2272 B.n998 B.n632 163.367
R2273 B.n998 B.n630 163.367
R2274 B.n1002 B.n630 163.367
R2275 B.n1002 B.n624 163.367
R2276 B.n1010 B.n624 163.367
R2277 B.n1010 B.n622 163.367
R2278 B.n1014 B.n622 163.367
R2279 B.n1014 B.n616 163.367
R2280 B.n1022 B.n616 163.367
R2281 B.n1022 B.n614 163.367
R2282 B.n1026 B.n614 163.367
R2283 B.n1026 B.n608 163.367
R2284 B.n1034 B.n608 163.367
R2285 B.n1034 B.n606 163.367
R2286 B.n1038 B.n606 163.367
R2287 B.n1038 B.n600 163.367
R2288 B.n1046 B.n600 163.367
R2289 B.n1046 B.n598 163.367
R2290 B.n1050 B.n598 163.367
R2291 B.n1050 B.n592 163.367
R2292 B.n1058 B.n592 163.367
R2293 B.n1058 B.n590 163.367
R2294 B.n1062 B.n590 163.367
R2295 B.n1062 B.n584 163.367
R2296 B.n1070 B.n584 163.367
R2297 B.n1070 B.n582 163.367
R2298 B.n1074 B.n582 163.367
R2299 B.n1074 B.n576 163.367
R2300 B.n1082 B.n576 163.367
R2301 B.n1082 B.n574 163.367
R2302 B.n1086 B.n574 163.367
R2303 B.n1086 B.n568 163.367
R2304 B.n1094 B.n568 163.367
R2305 B.n1094 B.n566 163.367
R2306 B.n1098 B.n566 163.367
R2307 B.n1098 B.n560 163.367
R2308 B.n1106 B.n560 163.367
R2309 B.n1106 B.n558 163.367
R2310 B.n1110 B.n558 163.367
R2311 B.n1110 B.n552 163.367
R2312 B.n1118 B.n552 163.367
R2313 B.n1118 B.n550 163.367
R2314 B.n1122 B.n550 163.367
R2315 B.n1122 B.n544 163.367
R2316 B.n1130 B.n544 163.367
R2317 B.n1130 B.n542 163.367
R2318 B.n1134 B.n542 163.367
R2319 B.n1134 B.n536 163.367
R2320 B.n1142 B.n536 163.367
R2321 B.n1142 B.n534 163.367
R2322 B.n1146 B.n534 163.367
R2323 B.n1146 B.n528 163.367
R2324 B.n1154 B.n528 163.367
R2325 B.n1154 B.n526 163.367
R2326 B.n1158 B.n526 163.367
R2327 B.n1158 B.n520 163.367
R2328 B.n1166 B.n520 163.367
R2329 B.n1166 B.n518 163.367
R2330 B.n1170 B.n518 163.367
R2331 B.n1170 B.n512 163.367
R2332 B.n1178 B.n512 163.367
R2333 B.n1178 B.n510 163.367
R2334 B.n1182 B.n510 163.367
R2335 B.n1182 B.n504 163.367
R2336 B.n1190 B.n504 163.367
R2337 B.n1190 B.n502 163.367
R2338 B.n1194 B.n502 163.367
R2339 B.n1194 B.n496 163.367
R2340 B.n1202 B.n496 163.367
R2341 B.n1202 B.n494 163.367
R2342 B.n1206 B.n494 163.367
R2343 B.n1206 B.n488 163.367
R2344 B.n1215 B.n488 163.367
R2345 B.n1215 B.n486 163.367
R2346 B.n1219 B.n486 163.367
R2347 B.n1219 B.n2 163.367
R2348 B.n1491 B.n2 163.367
R2349 B.n1491 B.n3 163.367
R2350 B.n1487 B.n3 163.367
R2351 B.n1487 B.n9 163.367
R2352 B.n1483 B.n9 163.367
R2353 B.n1483 B.n11 163.367
R2354 B.n1479 B.n11 163.367
R2355 B.n1479 B.n16 163.367
R2356 B.n1475 B.n16 163.367
R2357 B.n1475 B.n18 163.367
R2358 B.n1471 B.n18 163.367
R2359 B.n1471 B.n23 163.367
R2360 B.n1467 B.n23 163.367
R2361 B.n1467 B.n25 163.367
R2362 B.n1463 B.n25 163.367
R2363 B.n1463 B.n30 163.367
R2364 B.n1459 B.n30 163.367
R2365 B.n1459 B.n32 163.367
R2366 B.n1455 B.n32 163.367
R2367 B.n1455 B.n37 163.367
R2368 B.n1451 B.n37 163.367
R2369 B.n1451 B.n39 163.367
R2370 B.n1447 B.n39 163.367
R2371 B.n1447 B.n44 163.367
R2372 B.n1443 B.n44 163.367
R2373 B.n1443 B.n46 163.367
R2374 B.n1439 B.n46 163.367
R2375 B.n1439 B.n51 163.367
R2376 B.n1435 B.n51 163.367
R2377 B.n1435 B.n53 163.367
R2378 B.n1431 B.n53 163.367
R2379 B.n1431 B.n58 163.367
R2380 B.n1427 B.n58 163.367
R2381 B.n1427 B.n60 163.367
R2382 B.n1423 B.n60 163.367
R2383 B.n1423 B.n65 163.367
R2384 B.n1419 B.n65 163.367
R2385 B.n1419 B.n67 163.367
R2386 B.n1415 B.n67 163.367
R2387 B.n1415 B.n72 163.367
R2388 B.n1411 B.n72 163.367
R2389 B.n1411 B.n74 163.367
R2390 B.n1407 B.n74 163.367
R2391 B.n1407 B.n79 163.367
R2392 B.n1403 B.n79 163.367
R2393 B.n1403 B.n81 163.367
R2394 B.n1399 B.n81 163.367
R2395 B.n1399 B.n86 163.367
R2396 B.n1395 B.n86 163.367
R2397 B.n1395 B.n88 163.367
R2398 B.n1391 B.n88 163.367
R2399 B.n1391 B.n93 163.367
R2400 B.n1387 B.n93 163.367
R2401 B.n1387 B.n95 163.367
R2402 B.n1383 B.n95 163.367
R2403 B.n1383 B.n100 163.367
R2404 B.n1379 B.n100 163.367
R2405 B.n1379 B.n102 163.367
R2406 B.n1375 B.n102 163.367
R2407 B.n1375 B.n107 163.367
R2408 B.n1371 B.n107 163.367
R2409 B.n1371 B.n109 163.367
R2410 B.n1367 B.n109 163.367
R2411 B.n1367 B.n114 163.367
R2412 B.n1363 B.n114 163.367
R2413 B.n1363 B.n116 163.367
R2414 B.n1359 B.n116 163.367
R2415 B.n1359 B.n121 163.367
R2416 B.n1355 B.n121 163.367
R2417 B.n1355 B.n123 163.367
R2418 B.n1351 B.n123 163.367
R2419 B.n1351 B.n128 163.367
R2420 B.n1347 B.n128 163.367
R2421 B.n1347 B.n130 163.367
R2422 B.n1343 B.n130 163.367
R2423 B.n1343 B.n135 163.367
R2424 B.n1339 B.n135 163.367
R2425 B.n1339 B.n137 163.367
R2426 B.n1335 B.n137 163.367
R2427 B.n1335 B.n142 163.367
R2428 B.n1331 B.n142 163.367
R2429 B.n1331 B.n144 163.367
R2430 B.n710 B.n709 163.367
R2431 B.n971 B.n709 163.367
R2432 B.n969 B.n968 163.367
R2433 B.n965 B.n964 163.367
R2434 B.n961 B.n960 163.367
R2435 B.n957 B.n956 163.367
R2436 B.n953 B.n952 163.367
R2437 B.n949 B.n948 163.367
R2438 B.n945 B.n944 163.367
R2439 B.n941 B.n940 163.367
R2440 B.n937 B.n936 163.367
R2441 B.n933 B.n932 163.367
R2442 B.n929 B.n928 163.367
R2443 B.n925 B.n924 163.367
R2444 B.n921 B.n920 163.367
R2445 B.n917 B.n916 163.367
R2446 B.n913 B.n912 163.367
R2447 B.n909 B.n908 163.367
R2448 B.n905 B.n904 163.367
R2449 B.n901 B.n900 163.367
R2450 B.n897 B.n896 163.367
R2451 B.n893 B.n892 163.367
R2452 B.n889 B.n888 163.367
R2453 B.n885 B.n884 163.367
R2454 B.n881 B.n880 163.367
R2455 B.n877 B.n876 163.367
R2456 B.n873 B.n872 163.367
R2457 B.n869 B.n868 163.367
R2458 B.n865 B.n864 163.367
R2459 B.n861 B.n860 163.367
R2460 B.n857 B.n856 163.367
R2461 B.n852 B.n851 163.367
R2462 B.n848 B.n847 163.367
R2463 B.n844 B.n843 163.367
R2464 B.n840 B.n839 163.367
R2465 B.n836 B.n835 163.367
R2466 B.n832 B.n831 163.367
R2467 B.n828 B.n827 163.367
R2468 B.n824 B.n823 163.367
R2469 B.n820 B.n819 163.367
R2470 B.n816 B.n815 163.367
R2471 B.n812 B.n811 163.367
R2472 B.n808 B.n807 163.367
R2473 B.n804 B.n803 163.367
R2474 B.n800 B.n799 163.367
R2475 B.n796 B.n795 163.367
R2476 B.n792 B.n791 163.367
R2477 B.n788 B.n787 163.367
R2478 B.n784 B.n783 163.367
R2479 B.n780 B.n779 163.367
R2480 B.n776 B.n775 163.367
R2481 B.n772 B.n771 163.367
R2482 B.n768 B.n767 163.367
R2483 B.n764 B.n763 163.367
R2484 B.n760 B.n759 163.367
R2485 B.n756 B.n755 163.367
R2486 B.n752 B.n751 163.367
R2487 B.n748 B.n747 163.367
R2488 B.n744 B.n743 163.367
R2489 B.n740 B.n739 163.367
R2490 B.n736 B.n735 163.367
R2491 B.n732 B.n731 163.367
R2492 B.n728 B.n727 163.367
R2493 B.n724 B.n723 163.367
R2494 B.n720 B.n719 163.367
R2495 B.n716 B.n644 163.367
R2496 B.n984 B.n642 163.367
R2497 B.n984 B.n636 163.367
R2498 B.n992 B.n636 163.367
R2499 B.n992 B.n634 163.367
R2500 B.n996 B.n634 163.367
R2501 B.n996 B.n628 163.367
R2502 B.n1004 B.n628 163.367
R2503 B.n1004 B.n626 163.367
R2504 B.n1008 B.n626 163.367
R2505 B.n1008 B.n620 163.367
R2506 B.n1016 B.n620 163.367
R2507 B.n1016 B.n618 163.367
R2508 B.n1020 B.n618 163.367
R2509 B.n1020 B.n612 163.367
R2510 B.n1028 B.n612 163.367
R2511 B.n1028 B.n610 163.367
R2512 B.n1032 B.n610 163.367
R2513 B.n1032 B.n604 163.367
R2514 B.n1040 B.n604 163.367
R2515 B.n1040 B.n602 163.367
R2516 B.n1044 B.n602 163.367
R2517 B.n1044 B.n595 163.367
R2518 B.n1052 B.n595 163.367
R2519 B.n1052 B.n593 163.367
R2520 B.n1056 B.n593 163.367
R2521 B.n1056 B.n588 163.367
R2522 B.n1064 B.n588 163.367
R2523 B.n1064 B.n586 163.367
R2524 B.n1068 B.n586 163.367
R2525 B.n1068 B.n580 163.367
R2526 B.n1076 B.n580 163.367
R2527 B.n1076 B.n578 163.367
R2528 B.n1080 B.n578 163.367
R2529 B.n1080 B.n571 163.367
R2530 B.n1088 B.n571 163.367
R2531 B.n1088 B.n569 163.367
R2532 B.n1092 B.n569 163.367
R2533 B.n1092 B.n564 163.367
R2534 B.n1100 B.n564 163.367
R2535 B.n1100 B.n562 163.367
R2536 B.n1104 B.n562 163.367
R2537 B.n1104 B.n556 163.367
R2538 B.n1112 B.n556 163.367
R2539 B.n1112 B.n554 163.367
R2540 B.n1116 B.n554 163.367
R2541 B.n1116 B.n548 163.367
R2542 B.n1124 B.n548 163.367
R2543 B.n1124 B.n546 163.367
R2544 B.n1128 B.n546 163.367
R2545 B.n1128 B.n540 163.367
R2546 B.n1136 B.n540 163.367
R2547 B.n1136 B.n538 163.367
R2548 B.n1140 B.n538 163.367
R2549 B.n1140 B.n532 163.367
R2550 B.n1148 B.n532 163.367
R2551 B.n1148 B.n530 163.367
R2552 B.n1152 B.n530 163.367
R2553 B.n1152 B.n524 163.367
R2554 B.n1160 B.n524 163.367
R2555 B.n1160 B.n522 163.367
R2556 B.n1164 B.n522 163.367
R2557 B.n1164 B.n516 163.367
R2558 B.n1172 B.n516 163.367
R2559 B.n1172 B.n514 163.367
R2560 B.n1176 B.n514 163.367
R2561 B.n1176 B.n508 163.367
R2562 B.n1184 B.n508 163.367
R2563 B.n1184 B.n506 163.367
R2564 B.n1188 B.n506 163.367
R2565 B.n1188 B.n500 163.367
R2566 B.n1196 B.n500 163.367
R2567 B.n1196 B.n498 163.367
R2568 B.n1200 B.n498 163.367
R2569 B.n1200 B.n492 163.367
R2570 B.n1208 B.n492 163.367
R2571 B.n1208 B.n490 163.367
R2572 B.n1213 B.n490 163.367
R2573 B.n1213 B.n484 163.367
R2574 B.n1221 B.n484 163.367
R2575 B.n1222 B.n1221 163.367
R2576 B.n1222 B.n5 163.367
R2577 B.n6 B.n5 163.367
R2578 B.n7 B.n6 163.367
R2579 B.n1227 B.n7 163.367
R2580 B.n1227 B.n12 163.367
R2581 B.n13 B.n12 163.367
R2582 B.n14 B.n13 163.367
R2583 B.n1232 B.n14 163.367
R2584 B.n1232 B.n19 163.367
R2585 B.n20 B.n19 163.367
R2586 B.n21 B.n20 163.367
R2587 B.n1237 B.n21 163.367
R2588 B.n1237 B.n26 163.367
R2589 B.n27 B.n26 163.367
R2590 B.n28 B.n27 163.367
R2591 B.n1242 B.n28 163.367
R2592 B.n1242 B.n33 163.367
R2593 B.n34 B.n33 163.367
R2594 B.n35 B.n34 163.367
R2595 B.n1247 B.n35 163.367
R2596 B.n1247 B.n40 163.367
R2597 B.n41 B.n40 163.367
R2598 B.n42 B.n41 163.367
R2599 B.n1252 B.n42 163.367
R2600 B.n1252 B.n47 163.367
R2601 B.n48 B.n47 163.367
R2602 B.n49 B.n48 163.367
R2603 B.n1257 B.n49 163.367
R2604 B.n1257 B.n54 163.367
R2605 B.n55 B.n54 163.367
R2606 B.n56 B.n55 163.367
R2607 B.n1262 B.n56 163.367
R2608 B.n1262 B.n61 163.367
R2609 B.n62 B.n61 163.367
R2610 B.n63 B.n62 163.367
R2611 B.n1267 B.n63 163.367
R2612 B.n1267 B.n68 163.367
R2613 B.n69 B.n68 163.367
R2614 B.n70 B.n69 163.367
R2615 B.n1272 B.n70 163.367
R2616 B.n1272 B.n75 163.367
R2617 B.n76 B.n75 163.367
R2618 B.n77 B.n76 163.367
R2619 B.n1277 B.n77 163.367
R2620 B.n1277 B.n82 163.367
R2621 B.n83 B.n82 163.367
R2622 B.n84 B.n83 163.367
R2623 B.n1282 B.n84 163.367
R2624 B.n1282 B.n89 163.367
R2625 B.n90 B.n89 163.367
R2626 B.n91 B.n90 163.367
R2627 B.n1287 B.n91 163.367
R2628 B.n1287 B.n96 163.367
R2629 B.n97 B.n96 163.367
R2630 B.n98 B.n97 163.367
R2631 B.n1292 B.n98 163.367
R2632 B.n1292 B.n103 163.367
R2633 B.n104 B.n103 163.367
R2634 B.n105 B.n104 163.367
R2635 B.n1297 B.n105 163.367
R2636 B.n1297 B.n110 163.367
R2637 B.n111 B.n110 163.367
R2638 B.n112 B.n111 163.367
R2639 B.n1302 B.n112 163.367
R2640 B.n1302 B.n117 163.367
R2641 B.n118 B.n117 163.367
R2642 B.n119 B.n118 163.367
R2643 B.n1307 B.n119 163.367
R2644 B.n1307 B.n124 163.367
R2645 B.n125 B.n124 163.367
R2646 B.n126 B.n125 163.367
R2647 B.n1312 B.n126 163.367
R2648 B.n1312 B.n131 163.367
R2649 B.n132 B.n131 163.367
R2650 B.n133 B.n132 163.367
R2651 B.n1317 B.n133 163.367
R2652 B.n1317 B.n138 163.367
R2653 B.n139 B.n138 163.367
R2654 B.n140 B.n139 163.367
R2655 B.n1322 B.n140 163.367
R2656 B.n1322 B.n145 163.367
R2657 B.n146 B.n145 163.367
R2658 B.n223 B.n222 163.367
R2659 B.n227 B.n226 163.367
R2660 B.n231 B.n230 163.367
R2661 B.n235 B.n234 163.367
R2662 B.n239 B.n238 163.367
R2663 B.n243 B.n242 163.367
R2664 B.n247 B.n246 163.367
R2665 B.n251 B.n250 163.367
R2666 B.n255 B.n254 163.367
R2667 B.n259 B.n258 163.367
R2668 B.n263 B.n262 163.367
R2669 B.n267 B.n266 163.367
R2670 B.n271 B.n270 163.367
R2671 B.n275 B.n274 163.367
R2672 B.n279 B.n278 163.367
R2673 B.n283 B.n282 163.367
R2674 B.n287 B.n286 163.367
R2675 B.n291 B.n290 163.367
R2676 B.n295 B.n294 163.367
R2677 B.n299 B.n298 163.367
R2678 B.n303 B.n302 163.367
R2679 B.n307 B.n306 163.367
R2680 B.n311 B.n310 163.367
R2681 B.n315 B.n314 163.367
R2682 B.n319 B.n318 163.367
R2683 B.n323 B.n322 163.367
R2684 B.n327 B.n326 163.367
R2685 B.n331 B.n330 163.367
R2686 B.n335 B.n334 163.367
R2687 B.n339 B.n338 163.367
R2688 B.n343 B.n342 163.367
R2689 B.n347 B.n346 163.367
R2690 B.n351 B.n350 163.367
R2691 B.n355 B.n354 163.367
R2692 B.n359 B.n358 163.367
R2693 B.n364 B.n363 163.367
R2694 B.n368 B.n367 163.367
R2695 B.n372 B.n371 163.367
R2696 B.n376 B.n375 163.367
R2697 B.n380 B.n379 163.367
R2698 B.n384 B.n383 163.367
R2699 B.n388 B.n387 163.367
R2700 B.n392 B.n391 163.367
R2701 B.n396 B.n395 163.367
R2702 B.n400 B.n399 163.367
R2703 B.n404 B.n403 163.367
R2704 B.n408 B.n407 163.367
R2705 B.n412 B.n411 163.367
R2706 B.n416 B.n415 163.367
R2707 B.n420 B.n419 163.367
R2708 B.n424 B.n423 163.367
R2709 B.n428 B.n427 163.367
R2710 B.n432 B.n431 163.367
R2711 B.n436 B.n435 163.367
R2712 B.n440 B.n439 163.367
R2713 B.n444 B.n443 163.367
R2714 B.n448 B.n447 163.367
R2715 B.n452 B.n451 163.367
R2716 B.n456 B.n455 163.367
R2717 B.n460 B.n459 163.367
R2718 B.n464 B.n463 163.367
R2719 B.n468 B.n467 163.367
R2720 B.n472 B.n471 163.367
R2721 B.n476 B.n475 163.367
R2722 B.n480 B.n479 163.367
R2723 B.n1327 B.n213 163.367
R2724 B.n714 B.n713 79.9035
R2725 B.n712 B.n711 79.9035
R2726 B.n217 B.n216 79.9035
R2727 B.n215 B.n214 79.9035
R2728 B.n977 B.n976 71.676
R2729 B.n971 B.n645 71.676
R2730 B.n968 B.n646 71.676
R2731 B.n964 B.n647 71.676
R2732 B.n960 B.n648 71.676
R2733 B.n956 B.n649 71.676
R2734 B.n952 B.n650 71.676
R2735 B.n948 B.n651 71.676
R2736 B.n944 B.n652 71.676
R2737 B.n940 B.n653 71.676
R2738 B.n936 B.n654 71.676
R2739 B.n932 B.n655 71.676
R2740 B.n928 B.n656 71.676
R2741 B.n924 B.n657 71.676
R2742 B.n920 B.n658 71.676
R2743 B.n916 B.n659 71.676
R2744 B.n912 B.n660 71.676
R2745 B.n908 B.n661 71.676
R2746 B.n904 B.n662 71.676
R2747 B.n900 B.n663 71.676
R2748 B.n896 B.n664 71.676
R2749 B.n892 B.n665 71.676
R2750 B.n888 B.n666 71.676
R2751 B.n884 B.n667 71.676
R2752 B.n880 B.n668 71.676
R2753 B.n876 B.n669 71.676
R2754 B.n872 B.n670 71.676
R2755 B.n868 B.n671 71.676
R2756 B.n864 B.n672 71.676
R2757 B.n860 B.n673 71.676
R2758 B.n856 B.n674 71.676
R2759 B.n851 B.n675 71.676
R2760 B.n847 B.n676 71.676
R2761 B.n843 B.n677 71.676
R2762 B.n839 B.n678 71.676
R2763 B.n835 B.n679 71.676
R2764 B.n831 B.n680 71.676
R2765 B.n827 B.n681 71.676
R2766 B.n823 B.n682 71.676
R2767 B.n819 B.n683 71.676
R2768 B.n815 B.n684 71.676
R2769 B.n811 B.n685 71.676
R2770 B.n807 B.n686 71.676
R2771 B.n803 B.n687 71.676
R2772 B.n799 B.n688 71.676
R2773 B.n795 B.n689 71.676
R2774 B.n791 B.n690 71.676
R2775 B.n787 B.n691 71.676
R2776 B.n783 B.n692 71.676
R2777 B.n779 B.n693 71.676
R2778 B.n775 B.n694 71.676
R2779 B.n771 B.n695 71.676
R2780 B.n767 B.n696 71.676
R2781 B.n763 B.n697 71.676
R2782 B.n759 B.n698 71.676
R2783 B.n755 B.n699 71.676
R2784 B.n751 B.n700 71.676
R2785 B.n747 B.n701 71.676
R2786 B.n743 B.n702 71.676
R2787 B.n739 B.n703 71.676
R2788 B.n735 B.n704 71.676
R2789 B.n731 B.n705 71.676
R2790 B.n727 B.n706 71.676
R2791 B.n723 B.n707 71.676
R2792 B.n719 B.n708 71.676
R2793 B.n979 B.n644 71.676
R2794 B.n219 B.n147 71.676
R2795 B.n223 B.n148 71.676
R2796 B.n227 B.n149 71.676
R2797 B.n231 B.n150 71.676
R2798 B.n235 B.n151 71.676
R2799 B.n239 B.n152 71.676
R2800 B.n243 B.n153 71.676
R2801 B.n247 B.n154 71.676
R2802 B.n251 B.n155 71.676
R2803 B.n255 B.n156 71.676
R2804 B.n259 B.n157 71.676
R2805 B.n263 B.n158 71.676
R2806 B.n267 B.n159 71.676
R2807 B.n271 B.n160 71.676
R2808 B.n275 B.n161 71.676
R2809 B.n279 B.n162 71.676
R2810 B.n283 B.n163 71.676
R2811 B.n287 B.n164 71.676
R2812 B.n291 B.n165 71.676
R2813 B.n295 B.n166 71.676
R2814 B.n299 B.n167 71.676
R2815 B.n303 B.n168 71.676
R2816 B.n307 B.n169 71.676
R2817 B.n311 B.n170 71.676
R2818 B.n315 B.n171 71.676
R2819 B.n319 B.n172 71.676
R2820 B.n323 B.n173 71.676
R2821 B.n327 B.n174 71.676
R2822 B.n331 B.n175 71.676
R2823 B.n335 B.n176 71.676
R2824 B.n339 B.n177 71.676
R2825 B.n343 B.n178 71.676
R2826 B.n347 B.n179 71.676
R2827 B.n351 B.n180 71.676
R2828 B.n355 B.n181 71.676
R2829 B.n359 B.n182 71.676
R2830 B.n364 B.n183 71.676
R2831 B.n368 B.n184 71.676
R2832 B.n372 B.n185 71.676
R2833 B.n376 B.n186 71.676
R2834 B.n380 B.n187 71.676
R2835 B.n384 B.n188 71.676
R2836 B.n388 B.n189 71.676
R2837 B.n392 B.n190 71.676
R2838 B.n396 B.n191 71.676
R2839 B.n400 B.n192 71.676
R2840 B.n404 B.n193 71.676
R2841 B.n408 B.n194 71.676
R2842 B.n412 B.n195 71.676
R2843 B.n416 B.n196 71.676
R2844 B.n420 B.n197 71.676
R2845 B.n424 B.n198 71.676
R2846 B.n428 B.n199 71.676
R2847 B.n432 B.n200 71.676
R2848 B.n436 B.n201 71.676
R2849 B.n440 B.n202 71.676
R2850 B.n444 B.n203 71.676
R2851 B.n448 B.n204 71.676
R2852 B.n452 B.n205 71.676
R2853 B.n456 B.n206 71.676
R2854 B.n460 B.n207 71.676
R2855 B.n464 B.n208 71.676
R2856 B.n468 B.n209 71.676
R2857 B.n472 B.n210 71.676
R2858 B.n476 B.n211 71.676
R2859 B.n480 B.n212 71.676
R2860 B.n213 B.n212 71.676
R2861 B.n479 B.n211 71.676
R2862 B.n475 B.n210 71.676
R2863 B.n471 B.n209 71.676
R2864 B.n467 B.n208 71.676
R2865 B.n463 B.n207 71.676
R2866 B.n459 B.n206 71.676
R2867 B.n455 B.n205 71.676
R2868 B.n451 B.n204 71.676
R2869 B.n447 B.n203 71.676
R2870 B.n443 B.n202 71.676
R2871 B.n439 B.n201 71.676
R2872 B.n435 B.n200 71.676
R2873 B.n431 B.n199 71.676
R2874 B.n427 B.n198 71.676
R2875 B.n423 B.n197 71.676
R2876 B.n419 B.n196 71.676
R2877 B.n415 B.n195 71.676
R2878 B.n411 B.n194 71.676
R2879 B.n407 B.n193 71.676
R2880 B.n403 B.n192 71.676
R2881 B.n399 B.n191 71.676
R2882 B.n395 B.n190 71.676
R2883 B.n391 B.n189 71.676
R2884 B.n387 B.n188 71.676
R2885 B.n383 B.n187 71.676
R2886 B.n379 B.n186 71.676
R2887 B.n375 B.n185 71.676
R2888 B.n371 B.n184 71.676
R2889 B.n367 B.n183 71.676
R2890 B.n363 B.n182 71.676
R2891 B.n358 B.n181 71.676
R2892 B.n354 B.n180 71.676
R2893 B.n350 B.n179 71.676
R2894 B.n346 B.n178 71.676
R2895 B.n342 B.n177 71.676
R2896 B.n338 B.n176 71.676
R2897 B.n334 B.n175 71.676
R2898 B.n330 B.n174 71.676
R2899 B.n326 B.n173 71.676
R2900 B.n322 B.n172 71.676
R2901 B.n318 B.n171 71.676
R2902 B.n314 B.n170 71.676
R2903 B.n310 B.n169 71.676
R2904 B.n306 B.n168 71.676
R2905 B.n302 B.n167 71.676
R2906 B.n298 B.n166 71.676
R2907 B.n294 B.n165 71.676
R2908 B.n290 B.n164 71.676
R2909 B.n286 B.n163 71.676
R2910 B.n282 B.n162 71.676
R2911 B.n278 B.n161 71.676
R2912 B.n274 B.n160 71.676
R2913 B.n270 B.n159 71.676
R2914 B.n266 B.n158 71.676
R2915 B.n262 B.n157 71.676
R2916 B.n258 B.n156 71.676
R2917 B.n254 B.n155 71.676
R2918 B.n250 B.n154 71.676
R2919 B.n246 B.n153 71.676
R2920 B.n242 B.n152 71.676
R2921 B.n238 B.n151 71.676
R2922 B.n234 B.n150 71.676
R2923 B.n230 B.n149 71.676
R2924 B.n226 B.n148 71.676
R2925 B.n222 B.n147 71.676
R2926 B.n977 B.n710 71.676
R2927 B.n969 B.n645 71.676
R2928 B.n965 B.n646 71.676
R2929 B.n961 B.n647 71.676
R2930 B.n957 B.n648 71.676
R2931 B.n953 B.n649 71.676
R2932 B.n949 B.n650 71.676
R2933 B.n945 B.n651 71.676
R2934 B.n941 B.n652 71.676
R2935 B.n937 B.n653 71.676
R2936 B.n933 B.n654 71.676
R2937 B.n929 B.n655 71.676
R2938 B.n925 B.n656 71.676
R2939 B.n921 B.n657 71.676
R2940 B.n917 B.n658 71.676
R2941 B.n913 B.n659 71.676
R2942 B.n909 B.n660 71.676
R2943 B.n905 B.n661 71.676
R2944 B.n901 B.n662 71.676
R2945 B.n897 B.n663 71.676
R2946 B.n893 B.n664 71.676
R2947 B.n889 B.n665 71.676
R2948 B.n885 B.n666 71.676
R2949 B.n881 B.n667 71.676
R2950 B.n877 B.n668 71.676
R2951 B.n873 B.n669 71.676
R2952 B.n869 B.n670 71.676
R2953 B.n865 B.n671 71.676
R2954 B.n861 B.n672 71.676
R2955 B.n857 B.n673 71.676
R2956 B.n852 B.n674 71.676
R2957 B.n848 B.n675 71.676
R2958 B.n844 B.n676 71.676
R2959 B.n840 B.n677 71.676
R2960 B.n836 B.n678 71.676
R2961 B.n832 B.n679 71.676
R2962 B.n828 B.n680 71.676
R2963 B.n824 B.n681 71.676
R2964 B.n820 B.n682 71.676
R2965 B.n816 B.n683 71.676
R2966 B.n812 B.n684 71.676
R2967 B.n808 B.n685 71.676
R2968 B.n804 B.n686 71.676
R2969 B.n800 B.n687 71.676
R2970 B.n796 B.n688 71.676
R2971 B.n792 B.n689 71.676
R2972 B.n788 B.n690 71.676
R2973 B.n784 B.n691 71.676
R2974 B.n780 B.n692 71.676
R2975 B.n776 B.n693 71.676
R2976 B.n772 B.n694 71.676
R2977 B.n768 B.n695 71.676
R2978 B.n764 B.n696 71.676
R2979 B.n760 B.n697 71.676
R2980 B.n756 B.n698 71.676
R2981 B.n752 B.n699 71.676
R2982 B.n748 B.n700 71.676
R2983 B.n744 B.n701 71.676
R2984 B.n740 B.n702 71.676
R2985 B.n736 B.n703 71.676
R2986 B.n732 B.n704 71.676
R2987 B.n728 B.n705 71.676
R2988 B.n724 B.n706 71.676
R2989 B.n720 B.n707 71.676
R2990 B.n716 B.n708 71.676
R2991 B.n980 B.n979 71.676
R2992 B.n715 B.n714 59.5399
R2993 B.n854 B.n712 59.5399
R2994 B.n218 B.n217 59.5399
R2995 B.n361 B.n215 59.5399
R2996 B.n978 B.n641 50.5281
R2997 B.n1329 B.n1328 50.5281
R2998 B.n220 B.n143 32.3127
R2999 B.n1326 B.n1325 32.3127
R3000 B.n982 B.n981 32.3127
R3001 B.n975 B.n639 32.3127
R3002 B.n985 B.n641 30.9544
R3003 B.n985 B.n637 30.9544
R3004 B.n991 B.n637 30.9544
R3005 B.n991 B.n633 30.9544
R3006 B.n997 B.n633 30.9544
R3007 B.n997 B.n629 30.9544
R3008 B.n1003 B.n629 30.9544
R3009 B.n1003 B.n625 30.9544
R3010 B.n1009 B.n625 30.9544
R3011 B.n1015 B.n621 30.9544
R3012 B.n1015 B.n617 30.9544
R3013 B.n1021 B.n617 30.9544
R3014 B.n1021 B.n613 30.9544
R3015 B.n1027 B.n613 30.9544
R3016 B.n1027 B.n609 30.9544
R3017 B.n1033 B.n609 30.9544
R3018 B.n1033 B.n605 30.9544
R3019 B.n1039 B.n605 30.9544
R3020 B.n1039 B.n601 30.9544
R3021 B.n1045 B.n601 30.9544
R3022 B.n1045 B.n596 30.9544
R3023 B.n1051 B.n596 30.9544
R3024 B.n1051 B.n597 30.9544
R3025 B.n1057 B.n589 30.9544
R3026 B.n1063 B.n589 30.9544
R3027 B.n1063 B.n585 30.9544
R3028 B.n1069 B.n585 30.9544
R3029 B.n1069 B.n581 30.9544
R3030 B.n1075 B.n581 30.9544
R3031 B.n1075 B.n577 30.9544
R3032 B.n1081 B.n577 30.9544
R3033 B.n1081 B.n572 30.9544
R3034 B.n1087 B.n572 30.9544
R3035 B.n1087 B.n573 30.9544
R3036 B.n1093 B.n565 30.9544
R3037 B.n1099 B.n565 30.9544
R3038 B.n1099 B.n561 30.9544
R3039 B.n1105 B.n561 30.9544
R3040 B.n1105 B.n557 30.9544
R3041 B.n1111 B.n557 30.9544
R3042 B.n1111 B.n553 30.9544
R3043 B.n1117 B.n553 30.9544
R3044 B.n1117 B.n549 30.9544
R3045 B.n1123 B.n549 30.9544
R3046 B.n1123 B.n545 30.9544
R3047 B.n1129 B.n545 30.9544
R3048 B.n1135 B.n541 30.9544
R3049 B.n1135 B.n537 30.9544
R3050 B.n1141 B.n537 30.9544
R3051 B.n1141 B.n533 30.9544
R3052 B.n1147 B.n533 30.9544
R3053 B.n1147 B.n529 30.9544
R3054 B.n1153 B.n529 30.9544
R3055 B.n1153 B.n525 30.9544
R3056 B.n1159 B.n525 30.9544
R3057 B.n1159 B.n521 30.9544
R3058 B.n1165 B.n521 30.9544
R3059 B.n1171 B.n517 30.9544
R3060 B.n1171 B.n513 30.9544
R3061 B.n1177 B.n513 30.9544
R3062 B.n1177 B.n509 30.9544
R3063 B.n1183 B.n509 30.9544
R3064 B.n1183 B.n505 30.9544
R3065 B.n1189 B.n505 30.9544
R3066 B.n1189 B.n501 30.9544
R3067 B.n1195 B.n501 30.9544
R3068 B.n1195 B.n497 30.9544
R3069 B.n1201 B.n497 30.9544
R3070 B.n1207 B.n493 30.9544
R3071 B.n1207 B.n489 30.9544
R3072 B.n1214 B.n489 30.9544
R3073 B.n1214 B.n485 30.9544
R3074 B.n1220 B.n485 30.9544
R3075 B.n1220 B.n4 30.9544
R3076 B.n1490 B.n4 30.9544
R3077 B.n1490 B.n1489 30.9544
R3078 B.n1489 B.n1488 30.9544
R3079 B.n1488 B.n8 30.9544
R3080 B.n1482 B.n8 30.9544
R3081 B.n1482 B.n1481 30.9544
R3082 B.n1481 B.n1480 30.9544
R3083 B.n1480 B.n15 30.9544
R3084 B.n1474 B.n1473 30.9544
R3085 B.n1473 B.n1472 30.9544
R3086 B.n1472 B.n22 30.9544
R3087 B.n1466 B.n22 30.9544
R3088 B.n1466 B.n1465 30.9544
R3089 B.n1465 B.n1464 30.9544
R3090 B.n1464 B.n29 30.9544
R3091 B.n1458 B.n29 30.9544
R3092 B.n1458 B.n1457 30.9544
R3093 B.n1457 B.n1456 30.9544
R3094 B.n1456 B.n36 30.9544
R3095 B.n1450 B.n1449 30.9544
R3096 B.n1449 B.n1448 30.9544
R3097 B.n1448 B.n43 30.9544
R3098 B.n1442 B.n43 30.9544
R3099 B.n1442 B.n1441 30.9544
R3100 B.n1441 B.n1440 30.9544
R3101 B.n1440 B.n50 30.9544
R3102 B.n1434 B.n50 30.9544
R3103 B.n1434 B.n1433 30.9544
R3104 B.n1433 B.n1432 30.9544
R3105 B.n1432 B.n57 30.9544
R3106 B.n1426 B.n1425 30.9544
R3107 B.n1425 B.n1424 30.9544
R3108 B.n1424 B.n64 30.9544
R3109 B.n1418 B.n64 30.9544
R3110 B.n1418 B.n1417 30.9544
R3111 B.n1417 B.n1416 30.9544
R3112 B.n1416 B.n71 30.9544
R3113 B.n1410 B.n71 30.9544
R3114 B.n1410 B.n1409 30.9544
R3115 B.n1409 B.n1408 30.9544
R3116 B.n1408 B.n78 30.9544
R3117 B.n1402 B.n78 30.9544
R3118 B.n1401 B.n1400 30.9544
R3119 B.n1400 B.n85 30.9544
R3120 B.n1394 B.n85 30.9544
R3121 B.n1394 B.n1393 30.9544
R3122 B.n1393 B.n1392 30.9544
R3123 B.n1392 B.n92 30.9544
R3124 B.n1386 B.n92 30.9544
R3125 B.n1386 B.n1385 30.9544
R3126 B.n1385 B.n1384 30.9544
R3127 B.n1384 B.n99 30.9544
R3128 B.n1378 B.n99 30.9544
R3129 B.n1377 B.n1376 30.9544
R3130 B.n1376 B.n106 30.9544
R3131 B.n1370 B.n106 30.9544
R3132 B.n1370 B.n1369 30.9544
R3133 B.n1369 B.n1368 30.9544
R3134 B.n1368 B.n113 30.9544
R3135 B.n1362 B.n113 30.9544
R3136 B.n1362 B.n1361 30.9544
R3137 B.n1361 B.n1360 30.9544
R3138 B.n1360 B.n120 30.9544
R3139 B.n1354 B.n120 30.9544
R3140 B.n1354 B.n1353 30.9544
R3141 B.n1353 B.n1352 30.9544
R3142 B.n1352 B.n127 30.9544
R3143 B.n1346 B.n1345 30.9544
R3144 B.n1345 B.n1344 30.9544
R3145 B.n1344 B.n134 30.9544
R3146 B.n1338 B.n134 30.9544
R3147 B.n1338 B.n1337 30.9544
R3148 B.n1337 B.n1336 30.9544
R3149 B.n1336 B.n141 30.9544
R3150 B.n1330 B.n141 30.9544
R3151 B.n1330 B.n1329 30.9544
R3152 B.n573 B.t6 30.4992
R3153 B.t8 B.n1401 30.4992
R3154 B.t9 B.n541 27.7679
R3155 B.t2 B.n57 27.7679
R3156 B.n597 B.t1 26.8575
R3157 B.t0 B.n1377 26.8575
R3158 B.t5 B.n517 24.1263
R3159 B.t4 B.n36 24.1263
R3160 B.t3 B.n493 20.4847
R3161 B.t7 B.n15 20.4847
R3162 B B.n1492 18.0485
R3163 B.n1009 B.t11 16.843
R3164 B.n1346 B.t18 16.843
R3165 B.t11 B.n621 14.1118
R3166 B.t18 B.n127 14.1118
R3167 B.n221 B.n220 10.6151
R3168 B.n224 B.n221 10.6151
R3169 B.n225 B.n224 10.6151
R3170 B.n228 B.n225 10.6151
R3171 B.n229 B.n228 10.6151
R3172 B.n232 B.n229 10.6151
R3173 B.n233 B.n232 10.6151
R3174 B.n236 B.n233 10.6151
R3175 B.n237 B.n236 10.6151
R3176 B.n240 B.n237 10.6151
R3177 B.n241 B.n240 10.6151
R3178 B.n244 B.n241 10.6151
R3179 B.n245 B.n244 10.6151
R3180 B.n248 B.n245 10.6151
R3181 B.n249 B.n248 10.6151
R3182 B.n252 B.n249 10.6151
R3183 B.n253 B.n252 10.6151
R3184 B.n256 B.n253 10.6151
R3185 B.n257 B.n256 10.6151
R3186 B.n260 B.n257 10.6151
R3187 B.n261 B.n260 10.6151
R3188 B.n264 B.n261 10.6151
R3189 B.n265 B.n264 10.6151
R3190 B.n268 B.n265 10.6151
R3191 B.n269 B.n268 10.6151
R3192 B.n272 B.n269 10.6151
R3193 B.n273 B.n272 10.6151
R3194 B.n276 B.n273 10.6151
R3195 B.n277 B.n276 10.6151
R3196 B.n280 B.n277 10.6151
R3197 B.n281 B.n280 10.6151
R3198 B.n284 B.n281 10.6151
R3199 B.n285 B.n284 10.6151
R3200 B.n288 B.n285 10.6151
R3201 B.n289 B.n288 10.6151
R3202 B.n292 B.n289 10.6151
R3203 B.n293 B.n292 10.6151
R3204 B.n296 B.n293 10.6151
R3205 B.n297 B.n296 10.6151
R3206 B.n300 B.n297 10.6151
R3207 B.n301 B.n300 10.6151
R3208 B.n304 B.n301 10.6151
R3209 B.n305 B.n304 10.6151
R3210 B.n308 B.n305 10.6151
R3211 B.n309 B.n308 10.6151
R3212 B.n312 B.n309 10.6151
R3213 B.n313 B.n312 10.6151
R3214 B.n316 B.n313 10.6151
R3215 B.n317 B.n316 10.6151
R3216 B.n320 B.n317 10.6151
R3217 B.n321 B.n320 10.6151
R3218 B.n324 B.n321 10.6151
R3219 B.n325 B.n324 10.6151
R3220 B.n328 B.n325 10.6151
R3221 B.n329 B.n328 10.6151
R3222 B.n332 B.n329 10.6151
R3223 B.n333 B.n332 10.6151
R3224 B.n336 B.n333 10.6151
R3225 B.n337 B.n336 10.6151
R3226 B.n340 B.n337 10.6151
R3227 B.n341 B.n340 10.6151
R3228 B.n345 B.n344 10.6151
R3229 B.n348 B.n345 10.6151
R3230 B.n349 B.n348 10.6151
R3231 B.n352 B.n349 10.6151
R3232 B.n353 B.n352 10.6151
R3233 B.n356 B.n353 10.6151
R3234 B.n357 B.n356 10.6151
R3235 B.n360 B.n357 10.6151
R3236 B.n365 B.n362 10.6151
R3237 B.n366 B.n365 10.6151
R3238 B.n369 B.n366 10.6151
R3239 B.n370 B.n369 10.6151
R3240 B.n373 B.n370 10.6151
R3241 B.n374 B.n373 10.6151
R3242 B.n377 B.n374 10.6151
R3243 B.n378 B.n377 10.6151
R3244 B.n381 B.n378 10.6151
R3245 B.n382 B.n381 10.6151
R3246 B.n385 B.n382 10.6151
R3247 B.n386 B.n385 10.6151
R3248 B.n389 B.n386 10.6151
R3249 B.n390 B.n389 10.6151
R3250 B.n393 B.n390 10.6151
R3251 B.n394 B.n393 10.6151
R3252 B.n397 B.n394 10.6151
R3253 B.n398 B.n397 10.6151
R3254 B.n401 B.n398 10.6151
R3255 B.n402 B.n401 10.6151
R3256 B.n405 B.n402 10.6151
R3257 B.n406 B.n405 10.6151
R3258 B.n409 B.n406 10.6151
R3259 B.n410 B.n409 10.6151
R3260 B.n413 B.n410 10.6151
R3261 B.n414 B.n413 10.6151
R3262 B.n417 B.n414 10.6151
R3263 B.n418 B.n417 10.6151
R3264 B.n421 B.n418 10.6151
R3265 B.n422 B.n421 10.6151
R3266 B.n425 B.n422 10.6151
R3267 B.n426 B.n425 10.6151
R3268 B.n429 B.n426 10.6151
R3269 B.n430 B.n429 10.6151
R3270 B.n433 B.n430 10.6151
R3271 B.n434 B.n433 10.6151
R3272 B.n437 B.n434 10.6151
R3273 B.n438 B.n437 10.6151
R3274 B.n441 B.n438 10.6151
R3275 B.n442 B.n441 10.6151
R3276 B.n445 B.n442 10.6151
R3277 B.n446 B.n445 10.6151
R3278 B.n449 B.n446 10.6151
R3279 B.n450 B.n449 10.6151
R3280 B.n453 B.n450 10.6151
R3281 B.n454 B.n453 10.6151
R3282 B.n457 B.n454 10.6151
R3283 B.n458 B.n457 10.6151
R3284 B.n461 B.n458 10.6151
R3285 B.n462 B.n461 10.6151
R3286 B.n465 B.n462 10.6151
R3287 B.n466 B.n465 10.6151
R3288 B.n469 B.n466 10.6151
R3289 B.n470 B.n469 10.6151
R3290 B.n473 B.n470 10.6151
R3291 B.n474 B.n473 10.6151
R3292 B.n477 B.n474 10.6151
R3293 B.n478 B.n477 10.6151
R3294 B.n481 B.n478 10.6151
R3295 B.n482 B.n481 10.6151
R3296 B.n1326 B.n482 10.6151
R3297 B.n983 B.n982 10.6151
R3298 B.n983 B.n635 10.6151
R3299 B.n993 B.n635 10.6151
R3300 B.n994 B.n993 10.6151
R3301 B.n995 B.n994 10.6151
R3302 B.n995 B.n627 10.6151
R3303 B.n1005 B.n627 10.6151
R3304 B.n1006 B.n1005 10.6151
R3305 B.n1007 B.n1006 10.6151
R3306 B.n1007 B.n619 10.6151
R3307 B.n1017 B.n619 10.6151
R3308 B.n1018 B.n1017 10.6151
R3309 B.n1019 B.n1018 10.6151
R3310 B.n1019 B.n611 10.6151
R3311 B.n1029 B.n611 10.6151
R3312 B.n1030 B.n1029 10.6151
R3313 B.n1031 B.n1030 10.6151
R3314 B.n1031 B.n603 10.6151
R3315 B.n1041 B.n603 10.6151
R3316 B.n1042 B.n1041 10.6151
R3317 B.n1043 B.n1042 10.6151
R3318 B.n1043 B.n594 10.6151
R3319 B.n1053 B.n594 10.6151
R3320 B.n1054 B.n1053 10.6151
R3321 B.n1055 B.n1054 10.6151
R3322 B.n1055 B.n587 10.6151
R3323 B.n1065 B.n587 10.6151
R3324 B.n1066 B.n1065 10.6151
R3325 B.n1067 B.n1066 10.6151
R3326 B.n1067 B.n579 10.6151
R3327 B.n1077 B.n579 10.6151
R3328 B.n1078 B.n1077 10.6151
R3329 B.n1079 B.n1078 10.6151
R3330 B.n1079 B.n570 10.6151
R3331 B.n1089 B.n570 10.6151
R3332 B.n1090 B.n1089 10.6151
R3333 B.n1091 B.n1090 10.6151
R3334 B.n1091 B.n563 10.6151
R3335 B.n1101 B.n563 10.6151
R3336 B.n1102 B.n1101 10.6151
R3337 B.n1103 B.n1102 10.6151
R3338 B.n1103 B.n555 10.6151
R3339 B.n1113 B.n555 10.6151
R3340 B.n1114 B.n1113 10.6151
R3341 B.n1115 B.n1114 10.6151
R3342 B.n1115 B.n547 10.6151
R3343 B.n1125 B.n547 10.6151
R3344 B.n1126 B.n1125 10.6151
R3345 B.n1127 B.n1126 10.6151
R3346 B.n1127 B.n539 10.6151
R3347 B.n1137 B.n539 10.6151
R3348 B.n1138 B.n1137 10.6151
R3349 B.n1139 B.n1138 10.6151
R3350 B.n1139 B.n531 10.6151
R3351 B.n1149 B.n531 10.6151
R3352 B.n1150 B.n1149 10.6151
R3353 B.n1151 B.n1150 10.6151
R3354 B.n1151 B.n523 10.6151
R3355 B.n1161 B.n523 10.6151
R3356 B.n1162 B.n1161 10.6151
R3357 B.n1163 B.n1162 10.6151
R3358 B.n1163 B.n515 10.6151
R3359 B.n1173 B.n515 10.6151
R3360 B.n1174 B.n1173 10.6151
R3361 B.n1175 B.n1174 10.6151
R3362 B.n1175 B.n507 10.6151
R3363 B.n1185 B.n507 10.6151
R3364 B.n1186 B.n1185 10.6151
R3365 B.n1187 B.n1186 10.6151
R3366 B.n1187 B.n499 10.6151
R3367 B.n1197 B.n499 10.6151
R3368 B.n1198 B.n1197 10.6151
R3369 B.n1199 B.n1198 10.6151
R3370 B.n1199 B.n491 10.6151
R3371 B.n1209 B.n491 10.6151
R3372 B.n1210 B.n1209 10.6151
R3373 B.n1212 B.n1210 10.6151
R3374 B.n1212 B.n1211 10.6151
R3375 B.n1211 B.n483 10.6151
R3376 B.n1223 B.n483 10.6151
R3377 B.n1224 B.n1223 10.6151
R3378 B.n1225 B.n1224 10.6151
R3379 B.n1226 B.n1225 10.6151
R3380 B.n1228 B.n1226 10.6151
R3381 B.n1229 B.n1228 10.6151
R3382 B.n1230 B.n1229 10.6151
R3383 B.n1231 B.n1230 10.6151
R3384 B.n1233 B.n1231 10.6151
R3385 B.n1234 B.n1233 10.6151
R3386 B.n1235 B.n1234 10.6151
R3387 B.n1236 B.n1235 10.6151
R3388 B.n1238 B.n1236 10.6151
R3389 B.n1239 B.n1238 10.6151
R3390 B.n1240 B.n1239 10.6151
R3391 B.n1241 B.n1240 10.6151
R3392 B.n1243 B.n1241 10.6151
R3393 B.n1244 B.n1243 10.6151
R3394 B.n1245 B.n1244 10.6151
R3395 B.n1246 B.n1245 10.6151
R3396 B.n1248 B.n1246 10.6151
R3397 B.n1249 B.n1248 10.6151
R3398 B.n1250 B.n1249 10.6151
R3399 B.n1251 B.n1250 10.6151
R3400 B.n1253 B.n1251 10.6151
R3401 B.n1254 B.n1253 10.6151
R3402 B.n1255 B.n1254 10.6151
R3403 B.n1256 B.n1255 10.6151
R3404 B.n1258 B.n1256 10.6151
R3405 B.n1259 B.n1258 10.6151
R3406 B.n1260 B.n1259 10.6151
R3407 B.n1261 B.n1260 10.6151
R3408 B.n1263 B.n1261 10.6151
R3409 B.n1264 B.n1263 10.6151
R3410 B.n1265 B.n1264 10.6151
R3411 B.n1266 B.n1265 10.6151
R3412 B.n1268 B.n1266 10.6151
R3413 B.n1269 B.n1268 10.6151
R3414 B.n1270 B.n1269 10.6151
R3415 B.n1271 B.n1270 10.6151
R3416 B.n1273 B.n1271 10.6151
R3417 B.n1274 B.n1273 10.6151
R3418 B.n1275 B.n1274 10.6151
R3419 B.n1276 B.n1275 10.6151
R3420 B.n1278 B.n1276 10.6151
R3421 B.n1279 B.n1278 10.6151
R3422 B.n1280 B.n1279 10.6151
R3423 B.n1281 B.n1280 10.6151
R3424 B.n1283 B.n1281 10.6151
R3425 B.n1284 B.n1283 10.6151
R3426 B.n1285 B.n1284 10.6151
R3427 B.n1286 B.n1285 10.6151
R3428 B.n1288 B.n1286 10.6151
R3429 B.n1289 B.n1288 10.6151
R3430 B.n1290 B.n1289 10.6151
R3431 B.n1291 B.n1290 10.6151
R3432 B.n1293 B.n1291 10.6151
R3433 B.n1294 B.n1293 10.6151
R3434 B.n1295 B.n1294 10.6151
R3435 B.n1296 B.n1295 10.6151
R3436 B.n1298 B.n1296 10.6151
R3437 B.n1299 B.n1298 10.6151
R3438 B.n1300 B.n1299 10.6151
R3439 B.n1301 B.n1300 10.6151
R3440 B.n1303 B.n1301 10.6151
R3441 B.n1304 B.n1303 10.6151
R3442 B.n1305 B.n1304 10.6151
R3443 B.n1306 B.n1305 10.6151
R3444 B.n1308 B.n1306 10.6151
R3445 B.n1309 B.n1308 10.6151
R3446 B.n1310 B.n1309 10.6151
R3447 B.n1311 B.n1310 10.6151
R3448 B.n1313 B.n1311 10.6151
R3449 B.n1314 B.n1313 10.6151
R3450 B.n1315 B.n1314 10.6151
R3451 B.n1316 B.n1315 10.6151
R3452 B.n1318 B.n1316 10.6151
R3453 B.n1319 B.n1318 10.6151
R3454 B.n1320 B.n1319 10.6151
R3455 B.n1321 B.n1320 10.6151
R3456 B.n1323 B.n1321 10.6151
R3457 B.n1324 B.n1323 10.6151
R3458 B.n1325 B.n1324 10.6151
R3459 B.n975 B.n974 10.6151
R3460 B.n974 B.n973 10.6151
R3461 B.n973 B.n972 10.6151
R3462 B.n972 B.n970 10.6151
R3463 B.n970 B.n967 10.6151
R3464 B.n967 B.n966 10.6151
R3465 B.n966 B.n963 10.6151
R3466 B.n963 B.n962 10.6151
R3467 B.n962 B.n959 10.6151
R3468 B.n959 B.n958 10.6151
R3469 B.n958 B.n955 10.6151
R3470 B.n955 B.n954 10.6151
R3471 B.n954 B.n951 10.6151
R3472 B.n951 B.n950 10.6151
R3473 B.n950 B.n947 10.6151
R3474 B.n947 B.n946 10.6151
R3475 B.n946 B.n943 10.6151
R3476 B.n943 B.n942 10.6151
R3477 B.n942 B.n939 10.6151
R3478 B.n939 B.n938 10.6151
R3479 B.n938 B.n935 10.6151
R3480 B.n935 B.n934 10.6151
R3481 B.n934 B.n931 10.6151
R3482 B.n931 B.n930 10.6151
R3483 B.n930 B.n927 10.6151
R3484 B.n927 B.n926 10.6151
R3485 B.n926 B.n923 10.6151
R3486 B.n923 B.n922 10.6151
R3487 B.n922 B.n919 10.6151
R3488 B.n919 B.n918 10.6151
R3489 B.n918 B.n915 10.6151
R3490 B.n915 B.n914 10.6151
R3491 B.n914 B.n911 10.6151
R3492 B.n911 B.n910 10.6151
R3493 B.n910 B.n907 10.6151
R3494 B.n907 B.n906 10.6151
R3495 B.n906 B.n903 10.6151
R3496 B.n903 B.n902 10.6151
R3497 B.n902 B.n899 10.6151
R3498 B.n899 B.n898 10.6151
R3499 B.n898 B.n895 10.6151
R3500 B.n895 B.n894 10.6151
R3501 B.n894 B.n891 10.6151
R3502 B.n891 B.n890 10.6151
R3503 B.n890 B.n887 10.6151
R3504 B.n887 B.n886 10.6151
R3505 B.n886 B.n883 10.6151
R3506 B.n883 B.n882 10.6151
R3507 B.n882 B.n879 10.6151
R3508 B.n879 B.n878 10.6151
R3509 B.n878 B.n875 10.6151
R3510 B.n875 B.n874 10.6151
R3511 B.n874 B.n871 10.6151
R3512 B.n871 B.n870 10.6151
R3513 B.n870 B.n867 10.6151
R3514 B.n867 B.n866 10.6151
R3515 B.n866 B.n863 10.6151
R3516 B.n863 B.n862 10.6151
R3517 B.n862 B.n859 10.6151
R3518 B.n859 B.n858 10.6151
R3519 B.n858 B.n855 10.6151
R3520 B.n853 B.n850 10.6151
R3521 B.n850 B.n849 10.6151
R3522 B.n849 B.n846 10.6151
R3523 B.n846 B.n845 10.6151
R3524 B.n845 B.n842 10.6151
R3525 B.n842 B.n841 10.6151
R3526 B.n841 B.n838 10.6151
R3527 B.n838 B.n837 10.6151
R3528 B.n834 B.n833 10.6151
R3529 B.n833 B.n830 10.6151
R3530 B.n830 B.n829 10.6151
R3531 B.n829 B.n826 10.6151
R3532 B.n826 B.n825 10.6151
R3533 B.n825 B.n822 10.6151
R3534 B.n822 B.n821 10.6151
R3535 B.n821 B.n818 10.6151
R3536 B.n818 B.n817 10.6151
R3537 B.n817 B.n814 10.6151
R3538 B.n814 B.n813 10.6151
R3539 B.n813 B.n810 10.6151
R3540 B.n810 B.n809 10.6151
R3541 B.n809 B.n806 10.6151
R3542 B.n806 B.n805 10.6151
R3543 B.n805 B.n802 10.6151
R3544 B.n802 B.n801 10.6151
R3545 B.n801 B.n798 10.6151
R3546 B.n798 B.n797 10.6151
R3547 B.n797 B.n794 10.6151
R3548 B.n794 B.n793 10.6151
R3549 B.n793 B.n790 10.6151
R3550 B.n790 B.n789 10.6151
R3551 B.n789 B.n786 10.6151
R3552 B.n786 B.n785 10.6151
R3553 B.n785 B.n782 10.6151
R3554 B.n782 B.n781 10.6151
R3555 B.n781 B.n778 10.6151
R3556 B.n778 B.n777 10.6151
R3557 B.n777 B.n774 10.6151
R3558 B.n774 B.n773 10.6151
R3559 B.n773 B.n770 10.6151
R3560 B.n770 B.n769 10.6151
R3561 B.n769 B.n766 10.6151
R3562 B.n766 B.n765 10.6151
R3563 B.n765 B.n762 10.6151
R3564 B.n762 B.n761 10.6151
R3565 B.n761 B.n758 10.6151
R3566 B.n758 B.n757 10.6151
R3567 B.n757 B.n754 10.6151
R3568 B.n754 B.n753 10.6151
R3569 B.n753 B.n750 10.6151
R3570 B.n750 B.n749 10.6151
R3571 B.n749 B.n746 10.6151
R3572 B.n746 B.n745 10.6151
R3573 B.n745 B.n742 10.6151
R3574 B.n742 B.n741 10.6151
R3575 B.n741 B.n738 10.6151
R3576 B.n738 B.n737 10.6151
R3577 B.n737 B.n734 10.6151
R3578 B.n734 B.n733 10.6151
R3579 B.n733 B.n730 10.6151
R3580 B.n730 B.n729 10.6151
R3581 B.n729 B.n726 10.6151
R3582 B.n726 B.n725 10.6151
R3583 B.n725 B.n722 10.6151
R3584 B.n722 B.n721 10.6151
R3585 B.n721 B.n718 10.6151
R3586 B.n718 B.n717 10.6151
R3587 B.n717 B.n643 10.6151
R3588 B.n981 B.n643 10.6151
R3589 B.n987 B.n639 10.6151
R3590 B.n988 B.n987 10.6151
R3591 B.n989 B.n988 10.6151
R3592 B.n989 B.n631 10.6151
R3593 B.n999 B.n631 10.6151
R3594 B.n1000 B.n999 10.6151
R3595 B.n1001 B.n1000 10.6151
R3596 B.n1001 B.n623 10.6151
R3597 B.n1011 B.n623 10.6151
R3598 B.n1012 B.n1011 10.6151
R3599 B.n1013 B.n1012 10.6151
R3600 B.n1013 B.n615 10.6151
R3601 B.n1023 B.n615 10.6151
R3602 B.n1024 B.n1023 10.6151
R3603 B.n1025 B.n1024 10.6151
R3604 B.n1025 B.n607 10.6151
R3605 B.n1035 B.n607 10.6151
R3606 B.n1036 B.n1035 10.6151
R3607 B.n1037 B.n1036 10.6151
R3608 B.n1037 B.n599 10.6151
R3609 B.n1047 B.n599 10.6151
R3610 B.n1048 B.n1047 10.6151
R3611 B.n1049 B.n1048 10.6151
R3612 B.n1049 B.n591 10.6151
R3613 B.n1059 B.n591 10.6151
R3614 B.n1060 B.n1059 10.6151
R3615 B.n1061 B.n1060 10.6151
R3616 B.n1061 B.n583 10.6151
R3617 B.n1071 B.n583 10.6151
R3618 B.n1072 B.n1071 10.6151
R3619 B.n1073 B.n1072 10.6151
R3620 B.n1073 B.n575 10.6151
R3621 B.n1083 B.n575 10.6151
R3622 B.n1084 B.n1083 10.6151
R3623 B.n1085 B.n1084 10.6151
R3624 B.n1085 B.n567 10.6151
R3625 B.n1095 B.n567 10.6151
R3626 B.n1096 B.n1095 10.6151
R3627 B.n1097 B.n1096 10.6151
R3628 B.n1097 B.n559 10.6151
R3629 B.n1107 B.n559 10.6151
R3630 B.n1108 B.n1107 10.6151
R3631 B.n1109 B.n1108 10.6151
R3632 B.n1109 B.n551 10.6151
R3633 B.n1119 B.n551 10.6151
R3634 B.n1120 B.n1119 10.6151
R3635 B.n1121 B.n1120 10.6151
R3636 B.n1121 B.n543 10.6151
R3637 B.n1131 B.n543 10.6151
R3638 B.n1132 B.n1131 10.6151
R3639 B.n1133 B.n1132 10.6151
R3640 B.n1133 B.n535 10.6151
R3641 B.n1143 B.n535 10.6151
R3642 B.n1144 B.n1143 10.6151
R3643 B.n1145 B.n1144 10.6151
R3644 B.n1145 B.n527 10.6151
R3645 B.n1155 B.n527 10.6151
R3646 B.n1156 B.n1155 10.6151
R3647 B.n1157 B.n1156 10.6151
R3648 B.n1157 B.n519 10.6151
R3649 B.n1167 B.n519 10.6151
R3650 B.n1168 B.n1167 10.6151
R3651 B.n1169 B.n1168 10.6151
R3652 B.n1169 B.n511 10.6151
R3653 B.n1179 B.n511 10.6151
R3654 B.n1180 B.n1179 10.6151
R3655 B.n1181 B.n1180 10.6151
R3656 B.n1181 B.n503 10.6151
R3657 B.n1191 B.n503 10.6151
R3658 B.n1192 B.n1191 10.6151
R3659 B.n1193 B.n1192 10.6151
R3660 B.n1193 B.n495 10.6151
R3661 B.n1203 B.n495 10.6151
R3662 B.n1204 B.n1203 10.6151
R3663 B.n1205 B.n1204 10.6151
R3664 B.n1205 B.n487 10.6151
R3665 B.n1216 B.n487 10.6151
R3666 B.n1217 B.n1216 10.6151
R3667 B.n1218 B.n1217 10.6151
R3668 B.n1218 B.n0 10.6151
R3669 B.n1486 B.n1 10.6151
R3670 B.n1486 B.n1485 10.6151
R3671 B.n1485 B.n1484 10.6151
R3672 B.n1484 B.n10 10.6151
R3673 B.n1478 B.n10 10.6151
R3674 B.n1478 B.n1477 10.6151
R3675 B.n1477 B.n1476 10.6151
R3676 B.n1476 B.n17 10.6151
R3677 B.n1470 B.n17 10.6151
R3678 B.n1470 B.n1469 10.6151
R3679 B.n1469 B.n1468 10.6151
R3680 B.n1468 B.n24 10.6151
R3681 B.n1462 B.n24 10.6151
R3682 B.n1462 B.n1461 10.6151
R3683 B.n1461 B.n1460 10.6151
R3684 B.n1460 B.n31 10.6151
R3685 B.n1454 B.n31 10.6151
R3686 B.n1454 B.n1453 10.6151
R3687 B.n1453 B.n1452 10.6151
R3688 B.n1452 B.n38 10.6151
R3689 B.n1446 B.n38 10.6151
R3690 B.n1446 B.n1445 10.6151
R3691 B.n1445 B.n1444 10.6151
R3692 B.n1444 B.n45 10.6151
R3693 B.n1438 B.n45 10.6151
R3694 B.n1438 B.n1437 10.6151
R3695 B.n1437 B.n1436 10.6151
R3696 B.n1436 B.n52 10.6151
R3697 B.n1430 B.n52 10.6151
R3698 B.n1430 B.n1429 10.6151
R3699 B.n1429 B.n1428 10.6151
R3700 B.n1428 B.n59 10.6151
R3701 B.n1422 B.n59 10.6151
R3702 B.n1422 B.n1421 10.6151
R3703 B.n1421 B.n1420 10.6151
R3704 B.n1420 B.n66 10.6151
R3705 B.n1414 B.n66 10.6151
R3706 B.n1414 B.n1413 10.6151
R3707 B.n1413 B.n1412 10.6151
R3708 B.n1412 B.n73 10.6151
R3709 B.n1406 B.n73 10.6151
R3710 B.n1406 B.n1405 10.6151
R3711 B.n1405 B.n1404 10.6151
R3712 B.n1404 B.n80 10.6151
R3713 B.n1398 B.n80 10.6151
R3714 B.n1398 B.n1397 10.6151
R3715 B.n1397 B.n1396 10.6151
R3716 B.n1396 B.n87 10.6151
R3717 B.n1390 B.n87 10.6151
R3718 B.n1390 B.n1389 10.6151
R3719 B.n1389 B.n1388 10.6151
R3720 B.n1388 B.n94 10.6151
R3721 B.n1382 B.n94 10.6151
R3722 B.n1382 B.n1381 10.6151
R3723 B.n1381 B.n1380 10.6151
R3724 B.n1380 B.n101 10.6151
R3725 B.n1374 B.n101 10.6151
R3726 B.n1374 B.n1373 10.6151
R3727 B.n1373 B.n1372 10.6151
R3728 B.n1372 B.n108 10.6151
R3729 B.n1366 B.n108 10.6151
R3730 B.n1366 B.n1365 10.6151
R3731 B.n1365 B.n1364 10.6151
R3732 B.n1364 B.n115 10.6151
R3733 B.n1358 B.n115 10.6151
R3734 B.n1358 B.n1357 10.6151
R3735 B.n1357 B.n1356 10.6151
R3736 B.n1356 B.n122 10.6151
R3737 B.n1350 B.n122 10.6151
R3738 B.n1350 B.n1349 10.6151
R3739 B.n1349 B.n1348 10.6151
R3740 B.n1348 B.n129 10.6151
R3741 B.n1342 B.n129 10.6151
R3742 B.n1342 B.n1341 10.6151
R3743 B.n1341 B.n1340 10.6151
R3744 B.n1340 B.n136 10.6151
R3745 B.n1334 B.n136 10.6151
R3746 B.n1334 B.n1333 10.6151
R3747 B.n1333 B.n1332 10.6151
R3748 B.n1332 B.n143 10.6151
R3749 B.n1201 B.t3 10.4702
R3750 B.n1474 B.t7 10.4702
R3751 B.n1165 B.t5 6.82856
R3752 B.n1450 B.t4 6.82856
R3753 B.n344 B.n218 6.5566
R3754 B.n361 B.n360 6.5566
R3755 B.n854 B.n853 6.5566
R3756 B.n837 B.n715 6.5566
R3757 B.n1057 B.t1 4.09733
R3758 B.n1378 B.t0 4.09733
R3759 B.n341 B.n218 4.05904
R3760 B.n362 B.n361 4.05904
R3761 B.n855 B.n854 4.05904
R3762 B.n834 B.n715 4.05904
R3763 B.n1129 B.t9 3.18693
R3764 B.n1426 B.t2 3.18693
R3765 B.n1492 B.n0 2.81026
R3766 B.n1492 B.n1 2.81026
R3767 B.n1093 B.t6 0.455704
R3768 B.n1402 B.t8 0.455704
R3769 VN.n105 VN.n54 161.3
R3770 VN.n104 VN.n103 161.3
R3771 VN.n102 VN.n55 161.3
R3772 VN.n101 VN.n100 161.3
R3773 VN.n99 VN.n56 161.3
R3774 VN.n98 VN.n97 161.3
R3775 VN.n96 VN.n57 161.3
R3776 VN.n95 VN.n94 161.3
R3777 VN.n92 VN.n58 161.3
R3778 VN.n91 VN.n90 161.3
R3779 VN.n89 VN.n59 161.3
R3780 VN.n88 VN.n87 161.3
R3781 VN.n86 VN.n60 161.3
R3782 VN.n85 VN.n84 161.3
R3783 VN.n83 VN.n61 161.3
R3784 VN.n82 VN.n81 161.3
R3785 VN.n79 VN.n62 161.3
R3786 VN.n78 VN.n77 161.3
R3787 VN.n76 VN.n63 161.3
R3788 VN.n75 VN.n74 161.3
R3789 VN.n73 VN.n64 161.3
R3790 VN.n72 VN.n71 161.3
R3791 VN.n70 VN.n65 161.3
R3792 VN.n69 VN.n68 161.3
R3793 VN.n51 VN.n0 161.3
R3794 VN.n50 VN.n49 161.3
R3795 VN.n48 VN.n1 161.3
R3796 VN.n47 VN.n46 161.3
R3797 VN.n45 VN.n2 161.3
R3798 VN.n44 VN.n43 161.3
R3799 VN.n42 VN.n3 161.3
R3800 VN.n41 VN.n40 161.3
R3801 VN.n38 VN.n4 161.3
R3802 VN.n37 VN.n36 161.3
R3803 VN.n35 VN.n5 161.3
R3804 VN.n34 VN.n33 161.3
R3805 VN.n32 VN.n6 161.3
R3806 VN.n31 VN.n30 161.3
R3807 VN.n29 VN.n7 161.3
R3808 VN.n28 VN.n27 161.3
R3809 VN.n25 VN.n8 161.3
R3810 VN.n24 VN.n23 161.3
R3811 VN.n22 VN.n9 161.3
R3812 VN.n21 VN.n20 161.3
R3813 VN.n19 VN.n10 161.3
R3814 VN.n18 VN.n17 161.3
R3815 VN.n16 VN.n11 161.3
R3816 VN.n15 VN.n14 161.3
R3817 VN.n12 VN.t6 152.22
R3818 VN.n66 VN.t5 152.22
R3819 VN.n13 VN.t1 120.118
R3820 VN.n26 VN.t8 120.118
R3821 VN.n39 VN.t9 120.118
R3822 VN.n52 VN.t4 120.118
R3823 VN.n67 VN.t3 120.118
R3824 VN.n80 VN.t2 120.118
R3825 VN.n93 VN.t0 120.118
R3826 VN.n106 VN.t7 120.118
R3827 VN VN.n107 65.0951
R3828 VN.n53 VN.n52 58.2041
R3829 VN.n107 VN.n106 58.2041
R3830 VN.n13 VN.n12 56.9468
R3831 VN.n67 VN.n66 56.9468
R3832 VN.n20 VN.n19 56.5193
R3833 VN.n33 VN.n32 56.5193
R3834 VN.n74 VN.n73 56.5193
R3835 VN.n87 VN.n86 56.5193
R3836 VN.n46 VN.n45 47.2923
R3837 VN.n100 VN.n99 47.2923
R3838 VN.n46 VN.n1 33.6945
R3839 VN.n100 VN.n55 33.6945
R3840 VN.n14 VN.n11 24.4675
R3841 VN.n18 VN.n11 24.4675
R3842 VN.n19 VN.n18 24.4675
R3843 VN.n20 VN.n9 24.4675
R3844 VN.n24 VN.n9 24.4675
R3845 VN.n25 VN.n24 24.4675
R3846 VN.n27 VN.n7 24.4675
R3847 VN.n31 VN.n7 24.4675
R3848 VN.n32 VN.n31 24.4675
R3849 VN.n33 VN.n5 24.4675
R3850 VN.n37 VN.n5 24.4675
R3851 VN.n38 VN.n37 24.4675
R3852 VN.n40 VN.n3 24.4675
R3853 VN.n44 VN.n3 24.4675
R3854 VN.n45 VN.n44 24.4675
R3855 VN.n50 VN.n1 24.4675
R3856 VN.n51 VN.n50 24.4675
R3857 VN.n73 VN.n72 24.4675
R3858 VN.n72 VN.n65 24.4675
R3859 VN.n68 VN.n65 24.4675
R3860 VN.n86 VN.n85 24.4675
R3861 VN.n85 VN.n61 24.4675
R3862 VN.n81 VN.n61 24.4675
R3863 VN.n79 VN.n78 24.4675
R3864 VN.n78 VN.n63 24.4675
R3865 VN.n74 VN.n63 24.4675
R3866 VN.n99 VN.n98 24.4675
R3867 VN.n98 VN.n57 24.4675
R3868 VN.n94 VN.n57 24.4675
R3869 VN.n92 VN.n91 24.4675
R3870 VN.n91 VN.n59 24.4675
R3871 VN.n87 VN.n59 24.4675
R3872 VN.n105 VN.n104 24.4675
R3873 VN.n104 VN.n55 24.4675
R3874 VN.n52 VN.n51 23.9782
R3875 VN.n106 VN.n105 23.9782
R3876 VN.n14 VN.n13 18.1061
R3877 VN.n39 VN.n38 18.1061
R3878 VN.n68 VN.n67 18.1061
R3879 VN.n93 VN.n92 18.1061
R3880 VN.n26 VN.n25 12.234
R3881 VN.n27 VN.n26 12.234
R3882 VN.n81 VN.n80 12.234
R3883 VN.n80 VN.n79 12.234
R3884 VN.n40 VN.n39 6.36192
R3885 VN.n94 VN.n93 6.36192
R3886 VN.n69 VN.n66 2.54564
R3887 VN.n15 VN.n12 2.54564
R3888 VN.n107 VN.n54 0.417535
R3889 VN.n53 VN.n0 0.417535
R3890 VN VN.n53 0.394291
R3891 VN.n103 VN.n54 0.189894
R3892 VN.n103 VN.n102 0.189894
R3893 VN.n102 VN.n101 0.189894
R3894 VN.n101 VN.n56 0.189894
R3895 VN.n97 VN.n56 0.189894
R3896 VN.n97 VN.n96 0.189894
R3897 VN.n96 VN.n95 0.189894
R3898 VN.n95 VN.n58 0.189894
R3899 VN.n90 VN.n58 0.189894
R3900 VN.n90 VN.n89 0.189894
R3901 VN.n89 VN.n88 0.189894
R3902 VN.n88 VN.n60 0.189894
R3903 VN.n84 VN.n60 0.189894
R3904 VN.n84 VN.n83 0.189894
R3905 VN.n83 VN.n82 0.189894
R3906 VN.n82 VN.n62 0.189894
R3907 VN.n77 VN.n62 0.189894
R3908 VN.n77 VN.n76 0.189894
R3909 VN.n76 VN.n75 0.189894
R3910 VN.n75 VN.n64 0.189894
R3911 VN.n71 VN.n64 0.189894
R3912 VN.n71 VN.n70 0.189894
R3913 VN.n70 VN.n69 0.189894
R3914 VN.n16 VN.n15 0.189894
R3915 VN.n17 VN.n16 0.189894
R3916 VN.n17 VN.n10 0.189894
R3917 VN.n21 VN.n10 0.189894
R3918 VN.n22 VN.n21 0.189894
R3919 VN.n23 VN.n22 0.189894
R3920 VN.n23 VN.n8 0.189894
R3921 VN.n28 VN.n8 0.189894
R3922 VN.n29 VN.n28 0.189894
R3923 VN.n30 VN.n29 0.189894
R3924 VN.n30 VN.n6 0.189894
R3925 VN.n34 VN.n6 0.189894
R3926 VN.n35 VN.n34 0.189894
R3927 VN.n36 VN.n35 0.189894
R3928 VN.n36 VN.n4 0.189894
R3929 VN.n41 VN.n4 0.189894
R3930 VN.n42 VN.n41 0.189894
R3931 VN.n43 VN.n42 0.189894
R3932 VN.n43 VN.n2 0.189894
R3933 VN.n47 VN.n2 0.189894
R3934 VN.n48 VN.n47 0.189894
R3935 VN.n49 VN.n48 0.189894
R3936 VN.n49 VN.n0 0.189894
R3937 VDD2.n209 VDD2.n109 289.615
R3938 VDD2.n100 VDD2.n0 289.615
R3939 VDD2.n210 VDD2.n209 185
R3940 VDD2.n208 VDD2.n207 185
R3941 VDD2.n113 VDD2.n112 185
R3942 VDD2.n202 VDD2.n201 185
R3943 VDD2.n200 VDD2.n199 185
R3944 VDD2.n117 VDD2.n116 185
R3945 VDD2.n194 VDD2.n193 185
R3946 VDD2.n192 VDD2.n191 185
R3947 VDD2.n190 VDD2.n120 185
R3948 VDD2.n124 VDD2.n121 185
R3949 VDD2.n185 VDD2.n184 185
R3950 VDD2.n183 VDD2.n182 185
R3951 VDD2.n126 VDD2.n125 185
R3952 VDD2.n177 VDD2.n176 185
R3953 VDD2.n175 VDD2.n174 185
R3954 VDD2.n130 VDD2.n129 185
R3955 VDD2.n169 VDD2.n168 185
R3956 VDD2.n167 VDD2.n166 185
R3957 VDD2.n134 VDD2.n133 185
R3958 VDD2.n161 VDD2.n160 185
R3959 VDD2.n159 VDD2.n158 185
R3960 VDD2.n138 VDD2.n137 185
R3961 VDD2.n153 VDD2.n152 185
R3962 VDD2.n151 VDD2.n150 185
R3963 VDD2.n142 VDD2.n141 185
R3964 VDD2.n145 VDD2.n144 185
R3965 VDD2.n35 VDD2.n34 185
R3966 VDD2.n32 VDD2.n31 185
R3967 VDD2.n41 VDD2.n40 185
R3968 VDD2.n43 VDD2.n42 185
R3969 VDD2.n28 VDD2.n27 185
R3970 VDD2.n49 VDD2.n48 185
R3971 VDD2.n51 VDD2.n50 185
R3972 VDD2.n24 VDD2.n23 185
R3973 VDD2.n57 VDD2.n56 185
R3974 VDD2.n59 VDD2.n58 185
R3975 VDD2.n20 VDD2.n19 185
R3976 VDD2.n65 VDD2.n64 185
R3977 VDD2.n67 VDD2.n66 185
R3978 VDD2.n16 VDD2.n15 185
R3979 VDD2.n73 VDD2.n72 185
R3980 VDD2.n76 VDD2.n75 185
R3981 VDD2.n74 VDD2.n12 185
R3982 VDD2.n81 VDD2.n11 185
R3983 VDD2.n83 VDD2.n82 185
R3984 VDD2.n85 VDD2.n84 185
R3985 VDD2.n8 VDD2.n7 185
R3986 VDD2.n91 VDD2.n90 185
R3987 VDD2.n93 VDD2.n92 185
R3988 VDD2.n4 VDD2.n3 185
R3989 VDD2.n99 VDD2.n98 185
R3990 VDD2.n101 VDD2.n100 185
R3991 VDD2.t2 VDD2.n143 147.659
R3992 VDD2.t3 VDD2.n33 147.659
R3993 VDD2.n209 VDD2.n208 104.615
R3994 VDD2.n208 VDD2.n112 104.615
R3995 VDD2.n201 VDD2.n112 104.615
R3996 VDD2.n201 VDD2.n200 104.615
R3997 VDD2.n200 VDD2.n116 104.615
R3998 VDD2.n193 VDD2.n116 104.615
R3999 VDD2.n193 VDD2.n192 104.615
R4000 VDD2.n192 VDD2.n120 104.615
R4001 VDD2.n124 VDD2.n120 104.615
R4002 VDD2.n184 VDD2.n124 104.615
R4003 VDD2.n184 VDD2.n183 104.615
R4004 VDD2.n183 VDD2.n125 104.615
R4005 VDD2.n176 VDD2.n125 104.615
R4006 VDD2.n176 VDD2.n175 104.615
R4007 VDD2.n175 VDD2.n129 104.615
R4008 VDD2.n168 VDD2.n129 104.615
R4009 VDD2.n168 VDD2.n167 104.615
R4010 VDD2.n167 VDD2.n133 104.615
R4011 VDD2.n160 VDD2.n133 104.615
R4012 VDD2.n160 VDD2.n159 104.615
R4013 VDD2.n159 VDD2.n137 104.615
R4014 VDD2.n152 VDD2.n137 104.615
R4015 VDD2.n152 VDD2.n151 104.615
R4016 VDD2.n151 VDD2.n141 104.615
R4017 VDD2.n144 VDD2.n141 104.615
R4018 VDD2.n34 VDD2.n31 104.615
R4019 VDD2.n41 VDD2.n31 104.615
R4020 VDD2.n42 VDD2.n41 104.615
R4021 VDD2.n42 VDD2.n27 104.615
R4022 VDD2.n49 VDD2.n27 104.615
R4023 VDD2.n50 VDD2.n49 104.615
R4024 VDD2.n50 VDD2.n23 104.615
R4025 VDD2.n57 VDD2.n23 104.615
R4026 VDD2.n58 VDD2.n57 104.615
R4027 VDD2.n58 VDD2.n19 104.615
R4028 VDD2.n65 VDD2.n19 104.615
R4029 VDD2.n66 VDD2.n65 104.615
R4030 VDD2.n66 VDD2.n15 104.615
R4031 VDD2.n73 VDD2.n15 104.615
R4032 VDD2.n75 VDD2.n73 104.615
R4033 VDD2.n75 VDD2.n74 104.615
R4034 VDD2.n74 VDD2.n11 104.615
R4035 VDD2.n83 VDD2.n11 104.615
R4036 VDD2.n84 VDD2.n83 104.615
R4037 VDD2.n84 VDD2.n7 104.615
R4038 VDD2.n91 VDD2.n7 104.615
R4039 VDD2.n92 VDD2.n91 104.615
R4040 VDD2.n92 VDD2.n3 104.615
R4041 VDD2.n99 VDD2.n3 104.615
R4042 VDD2.n100 VDD2.n99 104.615
R4043 VDD2.n108 VDD2.n107 61.8729
R4044 VDD2 VDD2.n217 61.8698
R4045 VDD2.n216 VDD2.n215 59.2644
R4046 VDD2.n106 VDD2.n105 59.2644
R4047 VDD2.n214 VDD2.n108 56.8705
R4048 VDD2.n144 VDD2.t2 52.3082
R4049 VDD2.n34 VDD2.t3 52.3082
R4050 VDD2.n106 VDD2.n104 51.0583
R4051 VDD2.n214 VDD2.n213 47.5066
R4052 VDD2.n145 VDD2.n143 15.6677
R4053 VDD2.n35 VDD2.n33 15.6677
R4054 VDD2.n191 VDD2.n190 13.1884
R4055 VDD2.n82 VDD2.n81 13.1884
R4056 VDD2.n194 VDD2.n119 12.8005
R4057 VDD2.n189 VDD2.n121 12.8005
R4058 VDD2.n146 VDD2.n142 12.8005
R4059 VDD2.n36 VDD2.n32 12.8005
R4060 VDD2.n80 VDD2.n12 12.8005
R4061 VDD2.n85 VDD2.n10 12.8005
R4062 VDD2.n195 VDD2.n117 12.0247
R4063 VDD2.n186 VDD2.n185 12.0247
R4064 VDD2.n150 VDD2.n149 12.0247
R4065 VDD2.n40 VDD2.n39 12.0247
R4066 VDD2.n77 VDD2.n76 12.0247
R4067 VDD2.n86 VDD2.n8 12.0247
R4068 VDD2.n199 VDD2.n198 11.249
R4069 VDD2.n182 VDD2.n123 11.249
R4070 VDD2.n153 VDD2.n140 11.249
R4071 VDD2.n43 VDD2.n30 11.249
R4072 VDD2.n72 VDD2.n14 11.249
R4073 VDD2.n90 VDD2.n89 11.249
R4074 VDD2.n202 VDD2.n115 10.4732
R4075 VDD2.n181 VDD2.n126 10.4732
R4076 VDD2.n154 VDD2.n138 10.4732
R4077 VDD2.n44 VDD2.n28 10.4732
R4078 VDD2.n71 VDD2.n16 10.4732
R4079 VDD2.n93 VDD2.n6 10.4732
R4080 VDD2.n203 VDD2.n113 9.69747
R4081 VDD2.n178 VDD2.n177 9.69747
R4082 VDD2.n158 VDD2.n157 9.69747
R4083 VDD2.n48 VDD2.n47 9.69747
R4084 VDD2.n68 VDD2.n67 9.69747
R4085 VDD2.n94 VDD2.n4 9.69747
R4086 VDD2.n213 VDD2.n212 9.45567
R4087 VDD2.n104 VDD2.n103 9.45567
R4088 VDD2.n171 VDD2.n170 9.3005
R4089 VDD2.n173 VDD2.n172 9.3005
R4090 VDD2.n128 VDD2.n127 9.3005
R4091 VDD2.n179 VDD2.n178 9.3005
R4092 VDD2.n181 VDD2.n180 9.3005
R4093 VDD2.n123 VDD2.n122 9.3005
R4094 VDD2.n187 VDD2.n186 9.3005
R4095 VDD2.n189 VDD2.n188 9.3005
R4096 VDD2.n212 VDD2.n211 9.3005
R4097 VDD2.n111 VDD2.n110 9.3005
R4098 VDD2.n206 VDD2.n205 9.3005
R4099 VDD2.n204 VDD2.n203 9.3005
R4100 VDD2.n115 VDD2.n114 9.3005
R4101 VDD2.n198 VDD2.n197 9.3005
R4102 VDD2.n196 VDD2.n195 9.3005
R4103 VDD2.n119 VDD2.n118 9.3005
R4104 VDD2.n132 VDD2.n131 9.3005
R4105 VDD2.n165 VDD2.n164 9.3005
R4106 VDD2.n163 VDD2.n162 9.3005
R4107 VDD2.n136 VDD2.n135 9.3005
R4108 VDD2.n157 VDD2.n156 9.3005
R4109 VDD2.n155 VDD2.n154 9.3005
R4110 VDD2.n140 VDD2.n139 9.3005
R4111 VDD2.n149 VDD2.n148 9.3005
R4112 VDD2.n147 VDD2.n146 9.3005
R4113 VDD2.n2 VDD2.n1 9.3005
R4114 VDD2.n97 VDD2.n96 9.3005
R4115 VDD2.n95 VDD2.n94 9.3005
R4116 VDD2.n6 VDD2.n5 9.3005
R4117 VDD2.n89 VDD2.n88 9.3005
R4118 VDD2.n87 VDD2.n86 9.3005
R4119 VDD2.n10 VDD2.n9 9.3005
R4120 VDD2.n55 VDD2.n54 9.3005
R4121 VDD2.n53 VDD2.n52 9.3005
R4122 VDD2.n26 VDD2.n25 9.3005
R4123 VDD2.n47 VDD2.n46 9.3005
R4124 VDD2.n45 VDD2.n44 9.3005
R4125 VDD2.n30 VDD2.n29 9.3005
R4126 VDD2.n39 VDD2.n38 9.3005
R4127 VDD2.n37 VDD2.n36 9.3005
R4128 VDD2.n22 VDD2.n21 9.3005
R4129 VDD2.n61 VDD2.n60 9.3005
R4130 VDD2.n63 VDD2.n62 9.3005
R4131 VDD2.n18 VDD2.n17 9.3005
R4132 VDD2.n69 VDD2.n68 9.3005
R4133 VDD2.n71 VDD2.n70 9.3005
R4134 VDD2.n14 VDD2.n13 9.3005
R4135 VDD2.n78 VDD2.n77 9.3005
R4136 VDD2.n80 VDD2.n79 9.3005
R4137 VDD2.n103 VDD2.n102 9.3005
R4138 VDD2.n207 VDD2.n206 8.92171
R4139 VDD2.n174 VDD2.n128 8.92171
R4140 VDD2.n161 VDD2.n136 8.92171
R4141 VDD2.n51 VDD2.n26 8.92171
R4142 VDD2.n64 VDD2.n18 8.92171
R4143 VDD2.n98 VDD2.n97 8.92171
R4144 VDD2.n210 VDD2.n111 8.14595
R4145 VDD2.n173 VDD2.n130 8.14595
R4146 VDD2.n162 VDD2.n134 8.14595
R4147 VDD2.n52 VDD2.n24 8.14595
R4148 VDD2.n63 VDD2.n20 8.14595
R4149 VDD2.n101 VDD2.n2 8.14595
R4150 VDD2.n211 VDD2.n109 7.3702
R4151 VDD2.n170 VDD2.n169 7.3702
R4152 VDD2.n166 VDD2.n165 7.3702
R4153 VDD2.n56 VDD2.n55 7.3702
R4154 VDD2.n60 VDD2.n59 7.3702
R4155 VDD2.n102 VDD2.n0 7.3702
R4156 VDD2.n213 VDD2.n109 6.59444
R4157 VDD2.n169 VDD2.n132 6.59444
R4158 VDD2.n166 VDD2.n132 6.59444
R4159 VDD2.n56 VDD2.n22 6.59444
R4160 VDD2.n59 VDD2.n22 6.59444
R4161 VDD2.n104 VDD2.n0 6.59444
R4162 VDD2.n211 VDD2.n210 5.81868
R4163 VDD2.n170 VDD2.n130 5.81868
R4164 VDD2.n165 VDD2.n134 5.81868
R4165 VDD2.n55 VDD2.n24 5.81868
R4166 VDD2.n60 VDD2.n20 5.81868
R4167 VDD2.n102 VDD2.n101 5.81868
R4168 VDD2.n207 VDD2.n111 5.04292
R4169 VDD2.n174 VDD2.n173 5.04292
R4170 VDD2.n162 VDD2.n161 5.04292
R4171 VDD2.n52 VDD2.n51 5.04292
R4172 VDD2.n64 VDD2.n63 5.04292
R4173 VDD2.n98 VDD2.n2 5.04292
R4174 VDD2.n147 VDD2.n143 4.38563
R4175 VDD2.n37 VDD2.n33 4.38563
R4176 VDD2.n206 VDD2.n113 4.26717
R4177 VDD2.n177 VDD2.n128 4.26717
R4178 VDD2.n158 VDD2.n136 4.26717
R4179 VDD2.n48 VDD2.n26 4.26717
R4180 VDD2.n67 VDD2.n18 4.26717
R4181 VDD2.n97 VDD2.n4 4.26717
R4182 VDD2.n216 VDD2.n214 3.55222
R4183 VDD2.n203 VDD2.n202 3.49141
R4184 VDD2.n178 VDD2.n126 3.49141
R4185 VDD2.n157 VDD2.n138 3.49141
R4186 VDD2.n47 VDD2.n28 3.49141
R4187 VDD2.n68 VDD2.n16 3.49141
R4188 VDD2.n94 VDD2.n93 3.49141
R4189 VDD2.n199 VDD2.n115 2.71565
R4190 VDD2.n182 VDD2.n181 2.71565
R4191 VDD2.n154 VDD2.n153 2.71565
R4192 VDD2.n44 VDD2.n43 2.71565
R4193 VDD2.n72 VDD2.n71 2.71565
R4194 VDD2.n90 VDD2.n6 2.71565
R4195 VDD2.n198 VDD2.n117 1.93989
R4196 VDD2.n185 VDD2.n123 1.93989
R4197 VDD2.n150 VDD2.n140 1.93989
R4198 VDD2.n40 VDD2.n30 1.93989
R4199 VDD2.n76 VDD2.n14 1.93989
R4200 VDD2.n89 VDD2.n8 1.93989
R4201 VDD2.n195 VDD2.n194 1.16414
R4202 VDD2.n186 VDD2.n121 1.16414
R4203 VDD2.n149 VDD2.n142 1.16414
R4204 VDD2.n39 VDD2.n32 1.16414
R4205 VDD2.n77 VDD2.n12 1.16414
R4206 VDD2.n86 VDD2.n85 1.16414
R4207 VDD2.n217 VDD2.t6 1.04867
R4208 VDD2.n217 VDD2.t4 1.04867
R4209 VDD2.n215 VDD2.t9 1.04867
R4210 VDD2.n215 VDD2.t7 1.04867
R4211 VDD2.n107 VDD2.t0 1.04867
R4212 VDD2.n107 VDD2.t5 1.04867
R4213 VDD2.n105 VDD2.t8 1.04867
R4214 VDD2.n105 VDD2.t1 1.04867
R4215 VDD2 VDD2.n216 0.946621
R4216 VDD2.n108 VDD2.n106 0.833085
R4217 VDD2.n191 VDD2.n119 0.388379
R4218 VDD2.n190 VDD2.n189 0.388379
R4219 VDD2.n146 VDD2.n145 0.388379
R4220 VDD2.n36 VDD2.n35 0.388379
R4221 VDD2.n81 VDD2.n80 0.388379
R4222 VDD2.n82 VDD2.n10 0.388379
R4223 VDD2.n212 VDD2.n110 0.155672
R4224 VDD2.n205 VDD2.n110 0.155672
R4225 VDD2.n205 VDD2.n204 0.155672
R4226 VDD2.n204 VDD2.n114 0.155672
R4227 VDD2.n197 VDD2.n114 0.155672
R4228 VDD2.n197 VDD2.n196 0.155672
R4229 VDD2.n196 VDD2.n118 0.155672
R4230 VDD2.n188 VDD2.n118 0.155672
R4231 VDD2.n188 VDD2.n187 0.155672
R4232 VDD2.n187 VDD2.n122 0.155672
R4233 VDD2.n180 VDD2.n122 0.155672
R4234 VDD2.n180 VDD2.n179 0.155672
R4235 VDD2.n179 VDD2.n127 0.155672
R4236 VDD2.n172 VDD2.n127 0.155672
R4237 VDD2.n172 VDD2.n171 0.155672
R4238 VDD2.n171 VDD2.n131 0.155672
R4239 VDD2.n164 VDD2.n131 0.155672
R4240 VDD2.n164 VDD2.n163 0.155672
R4241 VDD2.n163 VDD2.n135 0.155672
R4242 VDD2.n156 VDD2.n135 0.155672
R4243 VDD2.n156 VDD2.n155 0.155672
R4244 VDD2.n155 VDD2.n139 0.155672
R4245 VDD2.n148 VDD2.n139 0.155672
R4246 VDD2.n148 VDD2.n147 0.155672
R4247 VDD2.n38 VDD2.n37 0.155672
R4248 VDD2.n38 VDD2.n29 0.155672
R4249 VDD2.n45 VDD2.n29 0.155672
R4250 VDD2.n46 VDD2.n45 0.155672
R4251 VDD2.n46 VDD2.n25 0.155672
R4252 VDD2.n53 VDD2.n25 0.155672
R4253 VDD2.n54 VDD2.n53 0.155672
R4254 VDD2.n54 VDD2.n21 0.155672
R4255 VDD2.n61 VDD2.n21 0.155672
R4256 VDD2.n62 VDD2.n61 0.155672
R4257 VDD2.n62 VDD2.n17 0.155672
R4258 VDD2.n69 VDD2.n17 0.155672
R4259 VDD2.n70 VDD2.n69 0.155672
R4260 VDD2.n70 VDD2.n13 0.155672
R4261 VDD2.n78 VDD2.n13 0.155672
R4262 VDD2.n79 VDD2.n78 0.155672
R4263 VDD2.n79 VDD2.n9 0.155672
R4264 VDD2.n87 VDD2.n9 0.155672
R4265 VDD2.n88 VDD2.n87 0.155672
R4266 VDD2.n88 VDD2.n5 0.155672
R4267 VDD2.n95 VDD2.n5 0.155672
R4268 VDD2.n96 VDD2.n95 0.155672
R4269 VDD2.n96 VDD2.n1 0.155672
R4270 VDD2.n103 VDD2.n1 0.155672
C0 VN VTAIL 18.403198f
C1 VDD2 VN 17.5818f
C2 VN VP 11.4323f
C3 VN VDD1 0.156084f
C4 VDD2 VTAIL 13.734f
C5 VTAIL VP 18.4183f
C6 VTAIL VDD1 13.6752f
C7 VDD2 VP 0.73508f
C8 VDD2 VDD1 2.95028f
C9 VDD1 VP 18.1566f
C10 VDD2 B 9.776757f
C11 VDD1 B 9.774592f
C12 VTAIL B 11.905766f
C13 VN B 24.36992f
C14 VP B 22.898764f
C15 VDD2.n0 B 0.032877f
C16 VDD2.n1 B 0.023732f
C17 VDD2.n2 B 0.012752f
C18 VDD2.n3 B 0.030142f
C19 VDD2.n4 B 0.013503f
C20 VDD2.n5 B 0.023732f
C21 VDD2.n6 B 0.012752f
C22 VDD2.n7 B 0.030142f
C23 VDD2.n8 B 0.013503f
C24 VDD2.n9 B 0.023732f
C25 VDD2.n10 B 0.012752f
C26 VDD2.n11 B 0.030142f
C27 VDD2.n12 B 0.013503f
C28 VDD2.n13 B 0.023732f
C29 VDD2.n14 B 0.012752f
C30 VDD2.n15 B 0.030142f
C31 VDD2.n16 B 0.013503f
C32 VDD2.n17 B 0.023732f
C33 VDD2.n18 B 0.012752f
C34 VDD2.n19 B 0.030142f
C35 VDD2.n20 B 0.013503f
C36 VDD2.n21 B 0.023732f
C37 VDD2.n22 B 0.012752f
C38 VDD2.n23 B 0.030142f
C39 VDD2.n24 B 0.013503f
C40 VDD2.n25 B 0.023732f
C41 VDD2.n26 B 0.012752f
C42 VDD2.n27 B 0.030142f
C43 VDD2.n28 B 0.013503f
C44 VDD2.n29 B 0.023732f
C45 VDD2.n30 B 0.012752f
C46 VDD2.n31 B 0.030142f
C47 VDD2.n32 B 0.013503f
C48 VDD2.n33 B 0.177929f
C49 VDD2.t3 B 0.050017f
C50 VDD2.n34 B 0.022606f
C51 VDD2.n35 B 0.017806f
C52 VDD2.n36 B 0.012752f
C53 VDD2.n37 B 1.96711f
C54 VDD2.n38 B 0.023732f
C55 VDD2.n39 B 0.012752f
C56 VDD2.n40 B 0.013503f
C57 VDD2.n41 B 0.030142f
C58 VDD2.n42 B 0.030142f
C59 VDD2.n43 B 0.013503f
C60 VDD2.n44 B 0.012752f
C61 VDD2.n45 B 0.023732f
C62 VDD2.n46 B 0.023732f
C63 VDD2.n47 B 0.012752f
C64 VDD2.n48 B 0.013503f
C65 VDD2.n49 B 0.030142f
C66 VDD2.n50 B 0.030142f
C67 VDD2.n51 B 0.013503f
C68 VDD2.n52 B 0.012752f
C69 VDD2.n53 B 0.023732f
C70 VDD2.n54 B 0.023732f
C71 VDD2.n55 B 0.012752f
C72 VDD2.n56 B 0.013503f
C73 VDD2.n57 B 0.030142f
C74 VDD2.n58 B 0.030142f
C75 VDD2.n59 B 0.013503f
C76 VDD2.n60 B 0.012752f
C77 VDD2.n61 B 0.023732f
C78 VDD2.n62 B 0.023732f
C79 VDD2.n63 B 0.012752f
C80 VDD2.n64 B 0.013503f
C81 VDD2.n65 B 0.030142f
C82 VDD2.n66 B 0.030142f
C83 VDD2.n67 B 0.013503f
C84 VDD2.n68 B 0.012752f
C85 VDD2.n69 B 0.023732f
C86 VDD2.n70 B 0.023732f
C87 VDD2.n71 B 0.012752f
C88 VDD2.n72 B 0.013503f
C89 VDD2.n73 B 0.030142f
C90 VDD2.n74 B 0.030142f
C91 VDD2.n75 B 0.030142f
C92 VDD2.n76 B 0.013503f
C93 VDD2.n77 B 0.012752f
C94 VDD2.n78 B 0.023732f
C95 VDD2.n79 B 0.023732f
C96 VDD2.n80 B 0.012752f
C97 VDD2.n81 B 0.013127f
C98 VDD2.n82 B 0.013127f
C99 VDD2.n83 B 0.030142f
C100 VDD2.n84 B 0.030142f
C101 VDD2.n85 B 0.013503f
C102 VDD2.n86 B 0.012752f
C103 VDD2.n87 B 0.023732f
C104 VDD2.n88 B 0.023732f
C105 VDD2.n89 B 0.012752f
C106 VDD2.n90 B 0.013503f
C107 VDD2.n91 B 0.030142f
C108 VDD2.n92 B 0.030142f
C109 VDD2.n93 B 0.013503f
C110 VDD2.n94 B 0.012752f
C111 VDD2.n95 B 0.023732f
C112 VDD2.n96 B 0.023732f
C113 VDD2.n97 B 0.012752f
C114 VDD2.n98 B 0.013503f
C115 VDD2.n99 B 0.030142f
C116 VDD2.n100 B 0.064403f
C117 VDD2.n101 B 0.013503f
C118 VDD2.n102 B 0.012752f
C119 VDD2.n103 B 0.052585f
C120 VDD2.n104 B 0.074264f
C121 VDD2.t8 B 0.354254f
C122 VDD2.t1 B 0.354254f
C123 VDD2.n105 B 3.23111f
C124 VDD2.n106 B 0.829995f
C125 VDD2.t0 B 0.354254f
C126 VDD2.t5 B 0.354254f
C127 VDD2.n107 B 3.25982f
C128 VDD2.n108 B 3.76132f
C129 VDD2.n109 B 0.032877f
C130 VDD2.n110 B 0.023732f
C131 VDD2.n111 B 0.012752f
C132 VDD2.n112 B 0.030142f
C133 VDD2.n113 B 0.013503f
C134 VDD2.n114 B 0.023732f
C135 VDD2.n115 B 0.012752f
C136 VDD2.n116 B 0.030142f
C137 VDD2.n117 B 0.013503f
C138 VDD2.n118 B 0.023732f
C139 VDD2.n119 B 0.012752f
C140 VDD2.n120 B 0.030142f
C141 VDD2.n121 B 0.013503f
C142 VDD2.n122 B 0.023732f
C143 VDD2.n123 B 0.012752f
C144 VDD2.n124 B 0.030142f
C145 VDD2.n125 B 0.030142f
C146 VDD2.n126 B 0.013503f
C147 VDD2.n127 B 0.023732f
C148 VDD2.n128 B 0.012752f
C149 VDD2.n129 B 0.030142f
C150 VDD2.n130 B 0.013503f
C151 VDD2.n131 B 0.023732f
C152 VDD2.n132 B 0.012752f
C153 VDD2.n133 B 0.030142f
C154 VDD2.n134 B 0.013503f
C155 VDD2.n135 B 0.023732f
C156 VDD2.n136 B 0.012752f
C157 VDD2.n137 B 0.030142f
C158 VDD2.n138 B 0.013503f
C159 VDD2.n139 B 0.023732f
C160 VDD2.n140 B 0.012752f
C161 VDD2.n141 B 0.030142f
C162 VDD2.n142 B 0.013503f
C163 VDD2.n143 B 0.177929f
C164 VDD2.t2 B 0.050017f
C165 VDD2.n144 B 0.022606f
C166 VDD2.n145 B 0.017806f
C167 VDD2.n146 B 0.012752f
C168 VDD2.n147 B 1.96711f
C169 VDD2.n148 B 0.023732f
C170 VDD2.n149 B 0.012752f
C171 VDD2.n150 B 0.013503f
C172 VDD2.n151 B 0.030142f
C173 VDD2.n152 B 0.030142f
C174 VDD2.n153 B 0.013503f
C175 VDD2.n154 B 0.012752f
C176 VDD2.n155 B 0.023732f
C177 VDD2.n156 B 0.023732f
C178 VDD2.n157 B 0.012752f
C179 VDD2.n158 B 0.013503f
C180 VDD2.n159 B 0.030142f
C181 VDD2.n160 B 0.030142f
C182 VDD2.n161 B 0.013503f
C183 VDD2.n162 B 0.012752f
C184 VDD2.n163 B 0.023732f
C185 VDD2.n164 B 0.023732f
C186 VDD2.n165 B 0.012752f
C187 VDD2.n166 B 0.013503f
C188 VDD2.n167 B 0.030142f
C189 VDD2.n168 B 0.030142f
C190 VDD2.n169 B 0.013503f
C191 VDD2.n170 B 0.012752f
C192 VDD2.n171 B 0.023732f
C193 VDD2.n172 B 0.023732f
C194 VDD2.n173 B 0.012752f
C195 VDD2.n174 B 0.013503f
C196 VDD2.n175 B 0.030142f
C197 VDD2.n176 B 0.030142f
C198 VDD2.n177 B 0.013503f
C199 VDD2.n178 B 0.012752f
C200 VDD2.n179 B 0.023732f
C201 VDD2.n180 B 0.023732f
C202 VDD2.n181 B 0.012752f
C203 VDD2.n182 B 0.013503f
C204 VDD2.n183 B 0.030142f
C205 VDD2.n184 B 0.030142f
C206 VDD2.n185 B 0.013503f
C207 VDD2.n186 B 0.012752f
C208 VDD2.n187 B 0.023732f
C209 VDD2.n188 B 0.023732f
C210 VDD2.n189 B 0.012752f
C211 VDD2.n190 B 0.013127f
C212 VDD2.n191 B 0.013127f
C213 VDD2.n192 B 0.030142f
C214 VDD2.n193 B 0.030142f
C215 VDD2.n194 B 0.013503f
C216 VDD2.n195 B 0.012752f
C217 VDD2.n196 B 0.023732f
C218 VDD2.n197 B 0.023732f
C219 VDD2.n198 B 0.012752f
C220 VDD2.n199 B 0.013503f
C221 VDD2.n200 B 0.030142f
C222 VDD2.n201 B 0.030142f
C223 VDD2.n202 B 0.013503f
C224 VDD2.n203 B 0.012752f
C225 VDD2.n204 B 0.023732f
C226 VDD2.n205 B 0.023732f
C227 VDD2.n206 B 0.012752f
C228 VDD2.n207 B 0.013503f
C229 VDD2.n208 B 0.030142f
C230 VDD2.n209 B 0.064403f
C231 VDD2.n210 B 0.013503f
C232 VDD2.n211 B 0.012752f
C233 VDD2.n212 B 0.052585f
C234 VDD2.n213 B 0.052283f
C235 VDD2.n214 B 3.67849f
C236 VDD2.t9 B 0.354254f
C237 VDD2.t7 B 0.354254f
C238 VDD2.n215 B 3.23112f
C239 VDD2.n216 B 0.544001f
C240 VDD2.t6 B 0.354254f
C241 VDD2.t4 B 0.354254f
C242 VDD2.n217 B 3.25976f
C243 VN.n0 B 0.02952f
C244 VN.t4 B 3.09314f
C245 VN.n1 B 0.031699f
C246 VN.n2 B 0.015693f
C247 VN.n3 B 0.029249f
C248 VN.n4 B 0.015693f
C249 VN.t9 B 3.09314f
C250 VN.n5 B 0.029249f
C251 VN.n6 B 0.015693f
C252 VN.n7 B 0.029249f
C253 VN.n8 B 0.015693f
C254 VN.t8 B 3.09314f
C255 VN.n9 B 0.029249f
C256 VN.n10 B 0.015693f
C257 VN.n11 B 0.029249f
C258 VN.t6 B 3.34371f
C259 VN.n12 B 1.07826f
C260 VN.t1 B 3.09314f
C261 VN.n13 B 1.12398f
C262 VN.n14 B 0.025494f
C263 VN.n15 B 0.202817f
C264 VN.n16 B 0.015693f
C265 VN.n17 B 0.015693f
C266 VN.n18 B 0.029249f
C267 VN.n19 B 0.020286f
C268 VN.n20 B 0.025534f
C269 VN.n21 B 0.015693f
C270 VN.n22 B 0.015693f
C271 VN.n23 B 0.015693f
C272 VN.n24 B 0.029249f
C273 VN.n25 B 0.022029f
C274 VN.n26 B 1.06401f
C275 VN.n27 B 0.022029f
C276 VN.n28 B 0.015693f
C277 VN.n29 B 0.015693f
C278 VN.n30 B 0.015693f
C279 VN.n31 B 0.029249f
C280 VN.n32 B 0.025534f
C281 VN.n33 B 0.020286f
C282 VN.n34 B 0.015693f
C283 VN.n35 B 0.015693f
C284 VN.n36 B 0.015693f
C285 VN.n37 B 0.029249f
C286 VN.n38 B 0.025494f
C287 VN.n39 B 1.06401f
C288 VN.n40 B 0.018563f
C289 VN.n41 B 0.015693f
C290 VN.n42 B 0.015693f
C291 VN.n43 B 0.015693f
C292 VN.n44 B 0.029249f
C293 VN.n45 B 0.029666f
C294 VN.n46 B 0.013703f
C295 VN.n47 B 0.015693f
C296 VN.n48 B 0.015693f
C297 VN.n49 B 0.015693f
C298 VN.n50 B 0.029249f
C299 VN.n51 B 0.02896f
C300 VN.n52 B 1.13466f
C301 VN.n53 B 0.045391f
C302 VN.n54 B 0.02952f
C303 VN.t7 B 3.09314f
C304 VN.n55 B 0.031699f
C305 VN.n56 B 0.015693f
C306 VN.n57 B 0.029249f
C307 VN.n58 B 0.015693f
C308 VN.t0 B 3.09314f
C309 VN.n59 B 0.029249f
C310 VN.n60 B 0.015693f
C311 VN.n61 B 0.029249f
C312 VN.n62 B 0.015693f
C313 VN.t2 B 3.09314f
C314 VN.n63 B 0.029249f
C315 VN.n64 B 0.015693f
C316 VN.n65 B 0.029249f
C317 VN.t5 B 3.34371f
C318 VN.n66 B 1.07826f
C319 VN.t3 B 3.09314f
C320 VN.n67 B 1.12398f
C321 VN.n68 B 0.025494f
C322 VN.n69 B 0.202817f
C323 VN.n70 B 0.015693f
C324 VN.n71 B 0.015693f
C325 VN.n72 B 0.029249f
C326 VN.n73 B 0.020286f
C327 VN.n74 B 0.025534f
C328 VN.n75 B 0.015693f
C329 VN.n76 B 0.015693f
C330 VN.n77 B 0.015693f
C331 VN.n78 B 0.029249f
C332 VN.n79 B 0.022029f
C333 VN.n80 B 1.06401f
C334 VN.n81 B 0.022029f
C335 VN.n82 B 0.015693f
C336 VN.n83 B 0.015693f
C337 VN.n84 B 0.015693f
C338 VN.n85 B 0.029249f
C339 VN.n86 B 0.025534f
C340 VN.n87 B 0.020286f
C341 VN.n88 B 0.015693f
C342 VN.n89 B 0.015693f
C343 VN.n90 B 0.015693f
C344 VN.n91 B 0.029249f
C345 VN.n92 B 0.025494f
C346 VN.n93 B 1.06401f
C347 VN.n94 B 0.018563f
C348 VN.n95 B 0.015693f
C349 VN.n96 B 0.015693f
C350 VN.n97 B 0.015693f
C351 VN.n98 B 0.029249f
C352 VN.n99 B 0.029666f
C353 VN.n100 B 0.013703f
C354 VN.n101 B 0.015693f
C355 VN.n102 B 0.015693f
C356 VN.n103 B 0.015693f
C357 VN.n104 B 0.029249f
C358 VN.n105 B 0.02896f
C359 VN.n106 B 1.13466f
C360 VN.n107 B 1.29824f
C361 VDD1.n0 B 0.033367f
C362 VDD1.n1 B 0.024085f
C363 VDD1.n2 B 0.012942f
C364 VDD1.n3 B 0.030591f
C365 VDD1.n4 B 0.013704f
C366 VDD1.n5 B 0.024085f
C367 VDD1.n6 B 0.012942f
C368 VDD1.n7 B 0.030591f
C369 VDD1.n8 B 0.013704f
C370 VDD1.n9 B 0.024085f
C371 VDD1.n10 B 0.012942f
C372 VDD1.n11 B 0.030591f
C373 VDD1.n12 B 0.013704f
C374 VDD1.n13 B 0.024085f
C375 VDD1.n14 B 0.012942f
C376 VDD1.n15 B 0.030591f
C377 VDD1.n16 B 0.030591f
C378 VDD1.n17 B 0.013704f
C379 VDD1.n18 B 0.024085f
C380 VDD1.n19 B 0.012942f
C381 VDD1.n20 B 0.030591f
C382 VDD1.n21 B 0.013704f
C383 VDD1.n22 B 0.024085f
C384 VDD1.n23 B 0.012942f
C385 VDD1.n24 B 0.030591f
C386 VDD1.n25 B 0.013704f
C387 VDD1.n26 B 0.024085f
C388 VDD1.n27 B 0.012942f
C389 VDD1.n28 B 0.030591f
C390 VDD1.n29 B 0.013704f
C391 VDD1.n30 B 0.024085f
C392 VDD1.n31 B 0.012942f
C393 VDD1.n32 B 0.030591f
C394 VDD1.n33 B 0.013704f
C395 VDD1.n34 B 0.18058f
C396 VDD1.t3 B 0.050763f
C397 VDD1.n35 B 0.022943f
C398 VDD1.n36 B 0.018071f
C399 VDD1.n37 B 0.012942f
C400 VDD1.n38 B 1.99642f
C401 VDD1.n39 B 0.024085f
C402 VDD1.n40 B 0.012942f
C403 VDD1.n41 B 0.013704f
C404 VDD1.n42 B 0.030591f
C405 VDD1.n43 B 0.030591f
C406 VDD1.n44 B 0.013704f
C407 VDD1.n45 B 0.012942f
C408 VDD1.n46 B 0.024085f
C409 VDD1.n47 B 0.024085f
C410 VDD1.n48 B 0.012942f
C411 VDD1.n49 B 0.013704f
C412 VDD1.n50 B 0.030591f
C413 VDD1.n51 B 0.030591f
C414 VDD1.n52 B 0.013704f
C415 VDD1.n53 B 0.012942f
C416 VDD1.n54 B 0.024085f
C417 VDD1.n55 B 0.024085f
C418 VDD1.n56 B 0.012942f
C419 VDD1.n57 B 0.013704f
C420 VDD1.n58 B 0.030591f
C421 VDD1.n59 B 0.030591f
C422 VDD1.n60 B 0.013704f
C423 VDD1.n61 B 0.012942f
C424 VDD1.n62 B 0.024085f
C425 VDD1.n63 B 0.024085f
C426 VDD1.n64 B 0.012942f
C427 VDD1.n65 B 0.013704f
C428 VDD1.n66 B 0.030591f
C429 VDD1.n67 B 0.030591f
C430 VDD1.n68 B 0.013704f
C431 VDD1.n69 B 0.012942f
C432 VDD1.n70 B 0.024085f
C433 VDD1.n71 B 0.024085f
C434 VDD1.n72 B 0.012942f
C435 VDD1.n73 B 0.013704f
C436 VDD1.n74 B 0.030591f
C437 VDD1.n75 B 0.030591f
C438 VDD1.n76 B 0.013704f
C439 VDD1.n77 B 0.012942f
C440 VDD1.n78 B 0.024085f
C441 VDD1.n79 B 0.024085f
C442 VDD1.n80 B 0.012942f
C443 VDD1.n81 B 0.013323f
C444 VDD1.n82 B 0.013323f
C445 VDD1.n83 B 0.030591f
C446 VDD1.n84 B 0.030591f
C447 VDD1.n85 B 0.013704f
C448 VDD1.n86 B 0.012942f
C449 VDD1.n87 B 0.024085f
C450 VDD1.n88 B 0.024085f
C451 VDD1.n89 B 0.012942f
C452 VDD1.n90 B 0.013704f
C453 VDD1.n91 B 0.030591f
C454 VDD1.n92 B 0.030591f
C455 VDD1.n93 B 0.013704f
C456 VDD1.n94 B 0.012942f
C457 VDD1.n95 B 0.024085f
C458 VDD1.n96 B 0.024085f
C459 VDD1.n97 B 0.012942f
C460 VDD1.n98 B 0.013704f
C461 VDD1.n99 B 0.030591f
C462 VDD1.n100 B 0.065363f
C463 VDD1.n101 B 0.013704f
C464 VDD1.n102 B 0.012942f
C465 VDD1.n103 B 0.053369f
C466 VDD1.n104 B 0.075371f
C467 VDD1.t4 B 0.359532f
C468 VDD1.t9 B 0.359532f
C469 VDD1.n105 B 3.27926f
C470 VDD1.n106 B 0.8505f
C471 VDD1.n107 B 0.033367f
C472 VDD1.n108 B 0.024085f
C473 VDD1.n109 B 0.012942f
C474 VDD1.n110 B 0.030591f
C475 VDD1.n111 B 0.013704f
C476 VDD1.n112 B 0.024085f
C477 VDD1.n113 B 0.012942f
C478 VDD1.n114 B 0.030591f
C479 VDD1.n115 B 0.013704f
C480 VDD1.n116 B 0.024085f
C481 VDD1.n117 B 0.012942f
C482 VDD1.n118 B 0.030591f
C483 VDD1.n119 B 0.013704f
C484 VDD1.n120 B 0.024085f
C485 VDD1.n121 B 0.012942f
C486 VDD1.n122 B 0.030591f
C487 VDD1.n123 B 0.013704f
C488 VDD1.n124 B 0.024085f
C489 VDD1.n125 B 0.012942f
C490 VDD1.n126 B 0.030591f
C491 VDD1.n127 B 0.013704f
C492 VDD1.n128 B 0.024085f
C493 VDD1.n129 B 0.012942f
C494 VDD1.n130 B 0.030591f
C495 VDD1.n131 B 0.013704f
C496 VDD1.n132 B 0.024085f
C497 VDD1.n133 B 0.012942f
C498 VDD1.n134 B 0.030591f
C499 VDD1.n135 B 0.013704f
C500 VDD1.n136 B 0.024085f
C501 VDD1.n137 B 0.012942f
C502 VDD1.n138 B 0.030591f
C503 VDD1.n139 B 0.013704f
C504 VDD1.n140 B 0.18058f
C505 VDD1.t0 B 0.050763f
C506 VDD1.n141 B 0.022943f
C507 VDD1.n142 B 0.018071f
C508 VDD1.n143 B 0.012942f
C509 VDD1.n144 B 1.99642f
C510 VDD1.n145 B 0.024085f
C511 VDD1.n146 B 0.012942f
C512 VDD1.n147 B 0.013704f
C513 VDD1.n148 B 0.030591f
C514 VDD1.n149 B 0.030591f
C515 VDD1.n150 B 0.013704f
C516 VDD1.n151 B 0.012942f
C517 VDD1.n152 B 0.024085f
C518 VDD1.n153 B 0.024085f
C519 VDD1.n154 B 0.012942f
C520 VDD1.n155 B 0.013704f
C521 VDD1.n156 B 0.030591f
C522 VDD1.n157 B 0.030591f
C523 VDD1.n158 B 0.013704f
C524 VDD1.n159 B 0.012942f
C525 VDD1.n160 B 0.024085f
C526 VDD1.n161 B 0.024085f
C527 VDD1.n162 B 0.012942f
C528 VDD1.n163 B 0.013704f
C529 VDD1.n164 B 0.030591f
C530 VDD1.n165 B 0.030591f
C531 VDD1.n166 B 0.013704f
C532 VDD1.n167 B 0.012942f
C533 VDD1.n168 B 0.024085f
C534 VDD1.n169 B 0.024085f
C535 VDD1.n170 B 0.012942f
C536 VDD1.n171 B 0.013704f
C537 VDD1.n172 B 0.030591f
C538 VDD1.n173 B 0.030591f
C539 VDD1.n174 B 0.013704f
C540 VDD1.n175 B 0.012942f
C541 VDD1.n176 B 0.024085f
C542 VDD1.n177 B 0.024085f
C543 VDD1.n178 B 0.012942f
C544 VDD1.n179 B 0.013704f
C545 VDD1.n180 B 0.030591f
C546 VDD1.n181 B 0.030591f
C547 VDD1.n182 B 0.030591f
C548 VDD1.n183 B 0.013704f
C549 VDD1.n184 B 0.012942f
C550 VDD1.n185 B 0.024085f
C551 VDD1.n186 B 0.024085f
C552 VDD1.n187 B 0.012942f
C553 VDD1.n188 B 0.013323f
C554 VDD1.n189 B 0.013323f
C555 VDD1.n190 B 0.030591f
C556 VDD1.n191 B 0.030591f
C557 VDD1.n192 B 0.013704f
C558 VDD1.n193 B 0.012942f
C559 VDD1.n194 B 0.024085f
C560 VDD1.n195 B 0.024085f
C561 VDD1.n196 B 0.012942f
C562 VDD1.n197 B 0.013704f
C563 VDD1.n198 B 0.030591f
C564 VDD1.n199 B 0.030591f
C565 VDD1.n200 B 0.013704f
C566 VDD1.n201 B 0.012942f
C567 VDD1.n202 B 0.024085f
C568 VDD1.n203 B 0.024085f
C569 VDD1.n204 B 0.012942f
C570 VDD1.n205 B 0.013704f
C571 VDD1.n206 B 0.030591f
C572 VDD1.n207 B 0.065363f
C573 VDD1.n208 B 0.013704f
C574 VDD1.n209 B 0.012942f
C575 VDD1.n210 B 0.053369f
C576 VDD1.n211 B 0.075371f
C577 VDD1.t8 B 0.359532f
C578 VDD1.t5 B 0.359532f
C579 VDD1.n212 B 3.27925f
C580 VDD1.n213 B 0.842361f
C581 VDD1.t6 B 0.359532f
C582 VDD1.t2 B 0.359532f
C583 VDD1.n214 B 3.30839f
C584 VDD1.n215 B 3.97411f
C585 VDD1.t1 B 0.359532f
C586 VDD1.t7 B 0.359532f
C587 VDD1.n216 B 3.27925f
C588 VDD1.n217 B 4.03541f
C589 VTAIL.t7 B 0.359563f
C590 VTAIL.t4 B 0.359563f
C591 VTAIL.n0 B 3.2018f
C592 VTAIL.n1 B 0.633612f
C593 VTAIL.n2 B 0.033369f
C594 VTAIL.n3 B 0.024087f
C595 VTAIL.n4 B 0.012943f
C596 VTAIL.n5 B 0.030594f
C597 VTAIL.n6 B 0.013705f
C598 VTAIL.n7 B 0.024087f
C599 VTAIL.n8 B 0.012943f
C600 VTAIL.n9 B 0.030594f
C601 VTAIL.n10 B 0.013705f
C602 VTAIL.n11 B 0.024087f
C603 VTAIL.n12 B 0.012943f
C604 VTAIL.n13 B 0.030594f
C605 VTAIL.n14 B 0.013705f
C606 VTAIL.n15 B 0.024087f
C607 VTAIL.n16 B 0.012943f
C608 VTAIL.n17 B 0.030594f
C609 VTAIL.n18 B 0.013705f
C610 VTAIL.n19 B 0.024087f
C611 VTAIL.n20 B 0.012943f
C612 VTAIL.n21 B 0.030594f
C613 VTAIL.n22 B 0.013705f
C614 VTAIL.n23 B 0.024087f
C615 VTAIL.n24 B 0.012943f
C616 VTAIL.n25 B 0.030594f
C617 VTAIL.n26 B 0.013705f
C618 VTAIL.n27 B 0.024087f
C619 VTAIL.n28 B 0.012943f
C620 VTAIL.n29 B 0.030594f
C621 VTAIL.n30 B 0.013705f
C622 VTAIL.n31 B 0.024087f
C623 VTAIL.n32 B 0.012943f
C624 VTAIL.n33 B 0.030594f
C625 VTAIL.n34 B 0.013705f
C626 VTAIL.n35 B 0.180596f
C627 VTAIL.t18 B 0.050767f
C628 VTAIL.n36 B 0.022945f
C629 VTAIL.n37 B 0.018073f
C630 VTAIL.n38 B 0.012943f
C631 VTAIL.n39 B 1.99659f
C632 VTAIL.n40 B 0.024087f
C633 VTAIL.n41 B 0.012943f
C634 VTAIL.n42 B 0.013705f
C635 VTAIL.n43 B 0.030594f
C636 VTAIL.n44 B 0.030594f
C637 VTAIL.n45 B 0.013705f
C638 VTAIL.n46 B 0.012943f
C639 VTAIL.n47 B 0.024087f
C640 VTAIL.n48 B 0.024087f
C641 VTAIL.n49 B 0.012943f
C642 VTAIL.n50 B 0.013705f
C643 VTAIL.n51 B 0.030594f
C644 VTAIL.n52 B 0.030594f
C645 VTAIL.n53 B 0.013705f
C646 VTAIL.n54 B 0.012943f
C647 VTAIL.n55 B 0.024087f
C648 VTAIL.n56 B 0.024087f
C649 VTAIL.n57 B 0.012943f
C650 VTAIL.n58 B 0.013705f
C651 VTAIL.n59 B 0.030594f
C652 VTAIL.n60 B 0.030594f
C653 VTAIL.n61 B 0.013705f
C654 VTAIL.n62 B 0.012943f
C655 VTAIL.n63 B 0.024087f
C656 VTAIL.n64 B 0.024087f
C657 VTAIL.n65 B 0.012943f
C658 VTAIL.n66 B 0.013705f
C659 VTAIL.n67 B 0.030594f
C660 VTAIL.n68 B 0.030594f
C661 VTAIL.n69 B 0.013705f
C662 VTAIL.n70 B 0.012943f
C663 VTAIL.n71 B 0.024087f
C664 VTAIL.n72 B 0.024087f
C665 VTAIL.n73 B 0.012943f
C666 VTAIL.n74 B 0.013705f
C667 VTAIL.n75 B 0.030594f
C668 VTAIL.n76 B 0.030594f
C669 VTAIL.n77 B 0.030594f
C670 VTAIL.n78 B 0.013705f
C671 VTAIL.n79 B 0.012943f
C672 VTAIL.n80 B 0.024087f
C673 VTAIL.n81 B 0.024087f
C674 VTAIL.n82 B 0.012943f
C675 VTAIL.n83 B 0.013324f
C676 VTAIL.n84 B 0.013324f
C677 VTAIL.n85 B 0.030594f
C678 VTAIL.n86 B 0.030594f
C679 VTAIL.n87 B 0.013705f
C680 VTAIL.n88 B 0.012943f
C681 VTAIL.n89 B 0.024087f
C682 VTAIL.n90 B 0.024087f
C683 VTAIL.n91 B 0.012943f
C684 VTAIL.n92 B 0.013705f
C685 VTAIL.n93 B 0.030594f
C686 VTAIL.n94 B 0.030594f
C687 VTAIL.n95 B 0.013705f
C688 VTAIL.n96 B 0.012943f
C689 VTAIL.n97 B 0.024087f
C690 VTAIL.n98 B 0.024087f
C691 VTAIL.n99 B 0.012943f
C692 VTAIL.n100 B 0.013705f
C693 VTAIL.n101 B 0.030594f
C694 VTAIL.n102 B 0.065368f
C695 VTAIL.n103 B 0.013705f
C696 VTAIL.n104 B 0.012943f
C697 VTAIL.n105 B 0.053373f
C698 VTAIL.n106 B 0.036415f
C699 VTAIL.n107 B 0.469239f
C700 VTAIL.t17 B 0.359563f
C701 VTAIL.t13 B 0.359563f
C702 VTAIL.n108 B 3.2018f
C703 VTAIL.n109 B 0.79938f
C704 VTAIL.t19 B 0.359563f
C705 VTAIL.t12 B 0.359563f
C706 VTAIL.n110 B 3.2018f
C707 VTAIL.n111 B 2.66616f
C708 VTAIL.t1 B 0.359563f
C709 VTAIL.t6 B 0.359563f
C710 VTAIL.n112 B 3.2018f
C711 VTAIL.n113 B 2.66616f
C712 VTAIL.t9 B 0.359563f
C713 VTAIL.t5 B 0.359563f
C714 VTAIL.n114 B 3.2018f
C715 VTAIL.n115 B 0.799378f
C716 VTAIL.n116 B 0.033369f
C717 VTAIL.n117 B 0.024087f
C718 VTAIL.n118 B 0.012943f
C719 VTAIL.n119 B 0.030594f
C720 VTAIL.n120 B 0.013705f
C721 VTAIL.n121 B 0.024087f
C722 VTAIL.n122 B 0.012943f
C723 VTAIL.n123 B 0.030594f
C724 VTAIL.n124 B 0.013705f
C725 VTAIL.n125 B 0.024087f
C726 VTAIL.n126 B 0.012943f
C727 VTAIL.n127 B 0.030594f
C728 VTAIL.n128 B 0.013705f
C729 VTAIL.n129 B 0.024087f
C730 VTAIL.n130 B 0.012943f
C731 VTAIL.n131 B 0.030594f
C732 VTAIL.n132 B 0.030594f
C733 VTAIL.n133 B 0.013705f
C734 VTAIL.n134 B 0.024087f
C735 VTAIL.n135 B 0.012943f
C736 VTAIL.n136 B 0.030594f
C737 VTAIL.n137 B 0.013705f
C738 VTAIL.n138 B 0.024087f
C739 VTAIL.n139 B 0.012943f
C740 VTAIL.n140 B 0.030594f
C741 VTAIL.n141 B 0.013705f
C742 VTAIL.n142 B 0.024087f
C743 VTAIL.n143 B 0.012943f
C744 VTAIL.n144 B 0.030594f
C745 VTAIL.n145 B 0.013705f
C746 VTAIL.n146 B 0.024087f
C747 VTAIL.n147 B 0.012943f
C748 VTAIL.n148 B 0.030594f
C749 VTAIL.n149 B 0.013705f
C750 VTAIL.n150 B 0.180596f
C751 VTAIL.t3 B 0.050767f
C752 VTAIL.n151 B 0.022945f
C753 VTAIL.n152 B 0.018073f
C754 VTAIL.n153 B 0.012943f
C755 VTAIL.n154 B 1.99659f
C756 VTAIL.n155 B 0.024087f
C757 VTAIL.n156 B 0.012943f
C758 VTAIL.n157 B 0.013705f
C759 VTAIL.n158 B 0.030594f
C760 VTAIL.n159 B 0.030594f
C761 VTAIL.n160 B 0.013705f
C762 VTAIL.n161 B 0.012943f
C763 VTAIL.n162 B 0.024087f
C764 VTAIL.n163 B 0.024087f
C765 VTAIL.n164 B 0.012943f
C766 VTAIL.n165 B 0.013705f
C767 VTAIL.n166 B 0.030594f
C768 VTAIL.n167 B 0.030594f
C769 VTAIL.n168 B 0.013705f
C770 VTAIL.n169 B 0.012943f
C771 VTAIL.n170 B 0.024087f
C772 VTAIL.n171 B 0.024087f
C773 VTAIL.n172 B 0.012943f
C774 VTAIL.n173 B 0.013705f
C775 VTAIL.n174 B 0.030594f
C776 VTAIL.n175 B 0.030594f
C777 VTAIL.n176 B 0.013705f
C778 VTAIL.n177 B 0.012943f
C779 VTAIL.n178 B 0.024087f
C780 VTAIL.n179 B 0.024087f
C781 VTAIL.n180 B 0.012943f
C782 VTAIL.n181 B 0.013705f
C783 VTAIL.n182 B 0.030594f
C784 VTAIL.n183 B 0.030594f
C785 VTAIL.n184 B 0.013705f
C786 VTAIL.n185 B 0.012943f
C787 VTAIL.n186 B 0.024087f
C788 VTAIL.n187 B 0.024087f
C789 VTAIL.n188 B 0.012943f
C790 VTAIL.n189 B 0.013705f
C791 VTAIL.n190 B 0.030594f
C792 VTAIL.n191 B 0.030594f
C793 VTAIL.n192 B 0.013705f
C794 VTAIL.n193 B 0.012943f
C795 VTAIL.n194 B 0.024087f
C796 VTAIL.n195 B 0.024087f
C797 VTAIL.n196 B 0.012943f
C798 VTAIL.n197 B 0.013324f
C799 VTAIL.n198 B 0.013324f
C800 VTAIL.n199 B 0.030594f
C801 VTAIL.n200 B 0.030594f
C802 VTAIL.n201 B 0.013705f
C803 VTAIL.n202 B 0.012943f
C804 VTAIL.n203 B 0.024087f
C805 VTAIL.n204 B 0.024087f
C806 VTAIL.n205 B 0.012943f
C807 VTAIL.n206 B 0.013705f
C808 VTAIL.n207 B 0.030594f
C809 VTAIL.n208 B 0.030594f
C810 VTAIL.n209 B 0.013705f
C811 VTAIL.n210 B 0.012943f
C812 VTAIL.n211 B 0.024087f
C813 VTAIL.n212 B 0.024087f
C814 VTAIL.n213 B 0.012943f
C815 VTAIL.n214 B 0.013705f
C816 VTAIL.n215 B 0.030594f
C817 VTAIL.n216 B 0.065368f
C818 VTAIL.n217 B 0.013705f
C819 VTAIL.n218 B 0.012943f
C820 VTAIL.n219 B 0.053373f
C821 VTAIL.n220 B 0.036415f
C822 VTAIL.n221 B 0.469239f
C823 VTAIL.t14 B 0.359563f
C824 VTAIL.t11 B 0.359563f
C825 VTAIL.n222 B 3.2018f
C826 VTAIL.n223 B 0.69801f
C827 VTAIL.t10 B 0.359563f
C828 VTAIL.t16 B 0.359563f
C829 VTAIL.n224 B 3.2018f
C830 VTAIL.n225 B 0.799378f
C831 VTAIL.n226 B 0.033369f
C832 VTAIL.n227 B 0.024087f
C833 VTAIL.n228 B 0.012943f
C834 VTAIL.n229 B 0.030594f
C835 VTAIL.n230 B 0.013705f
C836 VTAIL.n231 B 0.024087f
C837 VTAIL.n232 B 0.012943f
C838 VTAIL.n233 B 0.030594f
C839 VTAIL.n234 B 0.013705f
C840 VTAIL.n235 B 0.024087f
C841 VTAIL.n236 B 0.012943f
C842 VTAIL.n237 B 0.030594f
C843 VTAIL.n238 B 0.013705f
C844 VTAIL.n239 B 0.024087f
C845 VTAIL.n240 B 0.012943f
C846 VTAIL.n241 B 0.030594f
C847 VTAIL.n242 B 0.030594f
C848 VTAIL.n243 B 0.013705f
C849 VTAIL.n244 B 0.024087f
C850 VTAIL.n245 B 0.012943f
C851 VTAIL.n246 B 0.030594f
C852 VTAIL.n247 B 0.013705f
C853 VTAIL.n248 B 0.024087f
C854 VTAIL.n249 B 0.012943f
C855 VTAIL.n250 B 0.030594f
C856 VTAIL.n251 B 0.013705f
C857 VTAIL.n252 B 0.024087f
C858 VTAIL.n253 B 0.012943f
C859 VTAIL.n254 B 0.030594f
C860 VTAIL.n255 B 0.013705f
C861 VTAIL.n256 B 0.024087f
C862 VTAIL.n257 B 0.012943f
C863 VTAIL.n258 B 0.030594f
C864 VTAIL.n259 B 0.013705f
C865 VTAIL.n260 B 0.180596f
C866 VTAIL.t15 B 0.050767f
C867 VTAIL.n261 B 0.022945f
C868 VTAIL.n262 B 0.018073f
C869 VTAIL.n263 B 0.012943f
C870 VTAIL.n264 B 1.99659f
C871 VTAIL.n265 B 0.024087f
C872 VTAIL.n266 B 0.012943f
C873 VTAIL.n267 B 0.013705f
C874 VTAIL.n268 B 0.030594f
C875 VTAIL.n269 B 0.030594f
C876 VTAIL.n270 B 0.013705f
C877 VTAIL.n271 B 0.012943f
C878 VTAIL.n272 B 0.024087f
C879 VTAIL.n273 B 0.024087f
C880 VTAIL.n274 B 0.012943f
C881 VTAIL.n275 B 0.013705f
C882 VTAIL.n276 B 0.030594f
C883 VTAIL.n277 B 0.030594f
C884 VTAIL.n278 B 0.013705f
C885 VTAIL.n279 B 0.012943f
C886 VTAIL.n280 B 0.024087f
C887 VTAIL.n281 B 0.024087f
C888 VTAIL.n282 B 0.012943f
C889 VTAIL.n283 B 0.013705f
C890 VTAIL.n284 B 0.030594f
C891 VTAIL.n285 B 0.030594f
C892 VTAIL.n286 B 0.013705f
C893 VTAIL.n287 B 0.012943f
C894 VTAIL.n288 B 0.024087f
C895 VTAIL.n289 B 0.024087f
C896 VTAIL.n290 B 0.012943f
C897 VTAIL.n291 B 0.013705f
C898 VTAIL.n292 B 0.030594f
C899 VTAIL.n293 B 0.030594f
C900 VTAIL.n294 B 0.013705f
C901 VTAIL.n295 B 0.012943f
C902 VTAIL.n296 B 0.024087f
C903 VTAIL.n297 B 0.024087f
C904 VTAIL.n298 B 0.012943f
C905 VTAIL.n299 B 0.013705f
C906 VTAIL.n300 B 0.030594f
C907 VTAIL.n301 B 0.030594f
C908 VTAIL.n302 B 0.013705f
C909 VTAIL.n303 B 0.012943f
C910 VTAIL.n304 B 0.024087f
C911 VTAIL.n305 B 0.024087f
C912 VTAIL.n306 B 0.012943f
C913 VTAIL.n307 B 0.013324f
C914 VTAIL.n308 B 0.013324f
C915 VTAIL.n309 B 0.030594f
C916 VTAIL.n310 B 0.030594f
C917 VTAIL.n311 B 0.013705f
C918 VTAIL.n312 B 0.012943f
C919 VTAIL.n313 B 0.024087f
C920 VTAIL.n314 B 0.024087f
C921 VTAIL.n315 B 0.012943f
C922 VTAIL.n316 B 0.013705f
C923 VTAIL.n317 B 0.030594f
C924 VTAIL.n318 B 0.030594f
C925 VTAIL.n319 B 0.013705f
C926 VTAIL.n320 B 0.012943f
C927 VTAIL.n321 B 0.024087f
C928 VTAIL.n322 B 0.024087f
C929 VTAIL.n323 B 0.012943f
C930 VTAIL.n324 B 0.013705f
C931 VTAIL.n325 B 0.030594f
C932 VTAIL.n326 B 0.065368f
C933 VTAIL.n327 B 0.013705f
C934 VTAIL.n328 B 0.012943f
C935 VTAIL.n329 B 0.053373f
C936 VTAIL.n330 B 0.036415f
C937 VTAIL.n331 B 2.16172f
C938 VTAIL.n332 B 0.033369f
C939 VTAIL.n333 B 0.024087f
C940 VTAIL.n334 B 0.012943f
C941 VTAIL.n335 B 0.030594f
C942 VTAIL.n336 B 0.013705f
C943 VTAIL.n337 B 0.024087f
C944 VTAIL.n338 B 0.012943f
C945 VTAIL.n339 B 0.030594f
C946 VTAIL.n340 B 0.013705f
C947 VTAIL.n341 B 0.024087f
C948 VTAIL.n342 B 0.012943f
C949 VTAIL.n343 B 0.030594f
C950 VTAIL.n344 B 0.013705f
C951 VTAIL.n345 B 0.024087f
C952 VTAIL.n346 B 0.012943f
C953 VTAIL.n347 B 0.030594f
C954 VTAIL.n348 B 0.013705f
C955 VTAIL.n349 B 0.024087f
C956 VTAIL.n350 B 0.012943f
C957 VTAIL.n351 B 0.030594f
C958 VTAIL.n352 B 0.013705f
C959 VTAIL.n353 B 0.024087f
C960 VTAIL.n354 B 0.012943f
C961 VTAIL.n355 B 0.030594f
C962 VTAIL.n356 B 0.013705f
C963 VTAIL.n357 B 0.024087f
C964 VTAIL.n358 B 0.012943f
C965 VTAIL.n359 B 0.030594f
C966 VTAIL.n360 B 0.013705f
C967 VTAIL.n361 B 0.024087f
C968 VTAIL.n362 B 0.012943f
C969 VTAIL.n363 B 0.030594f
C970 VTAIL.n364 B 0.013705f
C971 VTAIL.n365 B 0.180596f
C972 VTAIL.t0 B 0.050767f
C973 VTAIL.n366 B 0.022945f
C974 VTAIL.n367 B 0.018073f
C975 VTAIL.n368 B 0.012943f
C976 VTAIL.n369 B 1.99659f
C977 VTAIL.n370 B 0.024087f
C978 VTAIL.n371 B 0.012943f
C979 VTAIL.n372 B 0.013705f
C980 VTAIL.n373 B 0.030594f
C981 VTAIL.n374 B 0.030594f
C982 VTAIL.n375 B 0.013705f
C983 VTAIL.n376 B 0.012943f
C984 VTAIL.n377 B 0.024087f
C985 VTAIL.n378 B 0.024087f
C986 VTAIL.n379 B 0.012943f
C987 VTAIL.n380 B 0.013705f
C988 VTAIL.n381 B 0.030594f
C989 VTAIL.n382 B 0.030594f
C990 VTAIL.n383 B 0.013705f
C991 VTAIL.n384 B 0.012943f
C992 VTAIL.n385 B 0.024087f
C993 VTAIL.n386 B 0.024087f
C994 VTAIL.n387 B 0.012943f
C995 VTAIL.n388 B 0.013705f
C996 VTAIL.n389 B 0.030594f
C997 VTAIL.n390 B 0.030594f
C998 VTAIL.n391 B 0.013705f
C999 VTAIL.n392 B 0.012943f
C1000 VTAIL.n393 B 0.024087f
C1001 VTAIL.n394 B 0.024087f
C1002 VTAIL.n395 B 0.012943f
C1003 VTAIL.n396 B 0.013705f
C1004 VTAIL.n397 B 0.030594f
C1005 VTAIL.n398 B 0.030594f
C1006 VTAIL.n399 B 0.013705f
C1007 VTAIL.n400 B 0.012943f
C1008 VTAIL.n401 B 0.024087f
C1009 VTAIL.n402 B 0.024087f
C1010 VTAIL.n403 B 0.012943f
C1011 VTAIL.n404 B 0.013705f
C1012 VTAIL.n405 B 0.030594f
C1013 VTAIL.n406 B 0.030594f
C1014 VTAIL.n407 B 0.030594f
C1015 VTAIL.n408 B 0.013705f
C1016 VTAIL.n409 B 0.012943f
C1017 VTAIL.n410 B 0.024087f
C1018 VTAIL.n411 B 0.024087f
C1019 VTAIL.n412 B 0.012943f
C1020 VTAIL.n413 B 0.013324f
C1021 VTAIL.n414 B 0.013324f
C1022 VTAIL.n415 B 0.030594f
C1023 VTAIL.n416 B 0.030594f
C1024 VTAIL.n417 B 0.013705f
C1025 VTAIL.n418 B 0.012943f
C1026 VTAIL.n419 B 0.024087f
C1027 VTAIL.n420 B 0.024087f
C1028 VTAIL.n421 B 0.012943f
C1029 VTAIL.n422 B 0.013705f
C1030 VTAIL.n423 B 0.030594f
C1031 VTAIL.n424 B 0.030594f
C1032 VTAIL.n425 B 0.013705f
C1033 VTAIL.n426 B 0.012943f
C1034 VTAIL.n427 B 0.024087f
C1035 VTAIL.n428 B 0.024087f
C1036 VTAIL.n429 B 0.012943f
C1037 VTAIL.n430 B 0.013705f
C1038 VTAIL.n431 B 0.030594f
C1039 VTAIL.n432 B 0.065368f
C1040 VTAIL.n433 B 0.013705f
C1041 VTAIL.n434 B 0.012943f
C1042 VTAIL.n435 B 0.053373f
C1043 VTAIL.n436 B 0.036415f
C1044 VTAIL.n437 B 2.16172f
C1045 VTAIL.t2 B 0.359563f
C1046 VTAIL.t8 B 0.359563f
C1047 VTAIL.n438 B 3.2018f
C1048 VTAIL.n439 B 0.588114f
C1049 VP.n0 B 0.029907f
C1050 VP.t7 B 3.13375f
C1051 VP.n1 B 0.032116f
C1052 VP.n2 B 0.015899f
C1053 VP.n3 B 0.029633f
C1054 VP.n4 B 0.015899f
C1055 VP.t3 B 3.13375f
C1056 VP.n5 B 0.029633f
C1057 VP.n6 B 0.015899f
C1058 VP.n7 B 0.029633f
C1059 VP.n8 B 0.015899f
C1060 VP.t4 B 3.13375f
C1061 VP.n9 B 0.029633f
C1062 VP.n10 B 0.015899f
C1063 VP.n11 B 0.029633f
C1064 VP.n12 B 0.015899f
C1065 VP.t1 B 3.13375f
C1066 VP.n13 B 0.029633f
C1067 VP.n14 B 0.015899f
C1068 VP.n15 B 0.029633f
C1069 VP.n16 B 0.029907f
C1070 VP.t2 B 3.13375f
C1071 VP.n17 B 0.032116f
C1072 VP.n18 B 0.015899f
C1073 VP.n19 B 0.029633f
C1074 VP.n20 B 0.015899f
C1075 VP.t8 B 3.13375f
C1076 VP.n21 B 0.029633f
C1077 VP.n22 B 0.015899f
C1078 VP.n23 B 0.029633f
C1079 VP.n24 B 0.015899f
C1080 VP.t0 B 3.13375f
C1081 VP.n25 B 0.029633f
C1082 VP.n26 B 0.015899f
C1083 VP.n27 B 0.029633f
C1084 VP.t6 B 3.38761f
C1085 VP.n28 B 1.09242f
C1086 VP.t5 B 3.13375f
C1087 VP.n29 B 1.13873f
C1088 VP.n30 B 0.025829f
C1089 VP.n31 B 0.20548f
C1090 VP.n32 B 0.015899f
C1091 VP.n33 B 0.015899f
C1092 VP.n34 B 0.029633f
C1093 VP.n35 B 0.020552f
C1094 VP.n36 B 0.025869f
C1095 VP.n37 B 0.015899f
C1096 VP.n38 B 0.015899f
C1097 VP.n39 B 0.015899f
C1098 VP.n40 B 0.029633f
C1099 VP.n41 B 0.022318f
C1100 VP.n42 B 1.07798f
C1101 VP.n43 B 0.022318f
C1102 VP.n44 B 0.015899f
C1103 VP.n45 B 0.015899f
C1104 VP.n46 B 0.015899f
C1105 VP.n47 B 0.029633f
C1106 VP.n48 B 0.025869f
C1107 VP.n49 B 0.020552f
C1108 VP.n50 B 0.015899f
C1109 VP.n51 B 0.015899f
C1110 VP.n52 B 0.015899f
C1111 VP.n53 B 0.029633f
C1112 VP.n54 B 0.025829f
C1113 VP.n55 B 1.07798f
C1114 VP.n56 B 0.018807f
C1115 VP.n57 B 0.015899f
C1116 VP.n58 B 0.015899f
C1117 VP.n59 B 0.015899f
C1118 VP.n60 B 0.029633f
C1119 VP.n61 B 0.030055f
C1120 VP.n62 B 0.013883f
C1121 VP.n63 B 0.015899f
C1122 VP.n64 B 0.015899f
C1123 VP.n65 B 0.015899f
C1124 VP.n66 B 0.029633f
C1125 VP.n67 B 0.02934f
C1126 VP.n68 B 1.14956f
C1127 VP.n69 B 1.31186f
C1128 VP.n70 B 1.32065f
C1129 VP.t9 B 3.13375f
C1130 VP.n71 B 1.14956f
C1131 VP.n72 B 0.02934f
C1132 VP.n73 B 0.029907f
C1133 VP.n74 B 0.015899f
C1134 VP.n75 B 0.015899f
C1135 VP.n76 B 0.032116f
C1136 VP.n77 B 0.013883f
C1137 VP.n78 B 0.030055f
C1138 VP.n79 B 0.015899f
C1139 VP.n80 B 0.015899f
C1140 VP.n81 B 0.015899f
C1141 VP.n82 B 0.029633f
C1142 VP.n83 B 0.018807f
C1143 VP.n84 B 1.07798f
C1144 VP.n85 B 0.025829f
C1145 VP.n86 B 0.015899f
C1146 VP.n87 B 0.015899f
C1147 VP.n88 B 0.015899f
C1148 VP.n89 B 0.029633f
C1149 VP.n90 B 0.020552f
C1150 VP.n91 B 0.025869f
C1151 VP.n92 B 0.015899f
C1152 VP.n93 B 0.015899f
C1153 VP.n94 B 0.015899f
C1154 VP.n95 B 0.029633f
C1155 VP.n96 B 0.022318f
C1156 VP.n97 B 1.07798f
C1157 VP.n98 B 0.022318f
C1158 VP.n99 B 0.015899f
C1159 VP.n100 B 0.015899f
C1160 VP.n101 B 0.015899f
C1161 VP.n102 B 0.029633f
C1162 VP.n103 B 0.025869f
C1163 VP.n104 B 0.020552f
C1164 VP.n105 B 0.015899f
C1165 VP.n106 B 0.015899f
C1166 VP.n107 B 0.015899f
C1167 VP.n108 B 0.029633f
C1168 VP.n109 B 0.025829f
C1169 VP.n110 B 1.07798f
C1170 VP.n111 B 0.018807f
C1171 VP.n112 B 0.015899f
C1172 VP.n113 B 0.015899f
C1173 VP.n114 B 0.015899f
C1174 VP.n115 B 0.029633f
C1175 VP.n116 B 0.030055f
C1176 VP.n117 B 0.013883f
C1177 VP.n118 B 0.015899f
C1178 VP.n119 B 0.015899f
C1179 VP.n120 B 0.015899f
C1180 VP.n121 B 0.029633f
C1181 VP.n122 B 0.02934f
C1182 VP.n123 B 1.14956f
C1183 VP.n124 B 0.045987f
.ends

