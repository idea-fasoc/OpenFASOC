* NGSPICE file created from diff_pair_sample_0190.ext - technology: sky130A

.subckt diff_pair_sample_0190 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t1 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=1.5774 ps=9.89 w=9.56 l=1.81
X1 VDD2.t0 VN.t1 VTAIL.t5 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=1.5774 pd=9.89 as=3.7284 ps=19.9 w=9.56 l=1.81
X2 VDD1.t3 VP.t0 VTAIL.t0 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=1.5774 pd=9.89 as=3.7284 ps=19.9 w=9.56 l=1.81
X3 B.t11 B.t9 B.t10 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=0 ps=0 w=9.56 l=1.81
X4 VDD1.t2 VP.t1 VTAIL.t1 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=1.5774 pd=9.89 as=3.7284 ps=19.9 w=9.56 l=1.81
X5 VDD2.t3 VN.t2 VTAIL.t4 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=1.5774 pd=9.89 as=3.7284 ps=19.9 w=9.56 l=1.81
X6 VTAIL.t7 VP.t2 VDD1.t1 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=1.5774 ps=9.89 w=9.56 l=1.81
X7 VTAIL.t3 VN.t3 VDD2.t2 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=1.5774 ps=9.89 w=9.56 l=1.81
X8 B.t8 B.t6 B.t7 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=0 ps=0 w=9.56 l=1.81
X9 B.t5 B.t3 B.t4 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=0 ps=0 w=9.56 l=1.81
X10 B.t2 B.t0 B.t1 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=0 ps=0 w=9.56 l=1.81
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n2254_n2880# sky130_fd_pr__pfet_01v8 ad=3.7284 pd=19.9 as=1.5774 ps=9.89 w=9.56 l=1.81
R0 VN.n0 VN.t3 163.905
R1 VN.n1 VN.t2 163.905
R2 VN.n0 VN.t1 163.475
R3 VN.n1 VN.t0 163.475
R4 VN VN.n1 51.6507
R5 VN VN.n0 9.31357
R6 VDD2.n2 VDD2.n0 114.535
R7 VDD2.n2 VDD2.n1 77.0444
R8 VDD2.n1 VDD2.t1 3.4006
R9 VDD2.n1 VDD2.t3 3.4006
R10 VDD2.n0 VDD2.t2 3.4006
R11 VDD2.n0 VDD2.t0 3.4006
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t7 63.7659
R14 VTAIL.n4 VTAIL.t4 63.7659
R15 VTAIL.n3 VTAIL.t6 63.7659
R16 VTAIL.n7 VTAIL.t5 63.7658
R17 VTAIL.n0 VTAIL.t3 63.7658
R18 VTAIL.n1 VTAIL.t1 63.7658
R19 VTAIL.n2 VTAIL.t2 63.7658
R20 VTAIL.n6 VTAIL.t0 63.7658
R21 VTAIL.n7 VTAIL.n6 22.4531
R22 VTAIL.n3 VTAIL.n2 22.4531
R23 VTAIL.n4 VTAIL.n3 1.84533
R24 VTAIL.n6 VTAIL.n5 1.84533
R25 VTAIL.n2 VTAIL.n1 1.84533
R26 VTAIL VTAIL.n0 0.981103
R27 VTAIL VTAIL.n7 0.864724
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 VP.n5 VP.n4 182.236
R31 VP.n14 VP.n13 182.236
R32 VP.n3 VP.t2 163.905
R33 VP.n3 VP.t0 163.475
R34 VP.n12 VP.n0 161.3
R35 VP.n11 VP.n10 161.3
R36 VP.n9 VP.n1 161.3
R37 VP.n8 VP.n7 161.3
R38 VP.n6 VP.n2 161.3
R39 VP.n5 VP.t3 127.291
R40 VP.n13 VP.t1 127.291
R41 VP.n4 VP.n3 51.27
R42 VP.n7 VP.n1 40.4106
R43 VP.n11 VP.n1 40.4106
R44 VP.n7 VP.n6 24.3439
R45 VP.n12 VP.n11 24.3439
R46 VP.n6 VP.n5 3.40858
R47 VP.n13 VP.n12 3.40858
R48 VP.n4 VP.n2 0.189894
R49 VP.n8 VP.n2 0.189894
R50 VP.n9 VP.n8 0.189894
R51 VP.n10 VP.n9 0.189894
R52 VP.n10 VP.n0 0.189894
R53 VP.n14 VP.n0 0.189894
R54 VP VP.n14 0.0516364
R55 VDD1 VDD1.n1 115.059
R56 VDD1 VDD1.n0 77.1026
R57 VDD1.n0 VDD1.t1 3.4006
R58 VDD1.n0 VDD1.t3 3.4006
R59 VDD1.n1 VDD1.t0 3.4006
R60 VDD1.n1 VDD1.t2 3.4006
R61 B.n384 B.n59 585
R62 B.n386 B.n385 585
R63 B.n387 B.n58 585
R64 B.n389 B.n388 585
R65 B.n390 B.n57 585
R66 B.n392 B.n391 585
R67 B.n393 B.n56 585
R68 B.n395 B.n394 585
R69 B.n396 B.n55 585
R70 B.n398 B.n397 585
R71 B.n399 B.n54 585
R72 B.n401 B.n400 585
R73 B.n402 B.n53 585
R74 B.n404 B.n403 585
R75 B.n405 B.n52 585
R76 B.n407 B.n406 585
R77 B.n408 B.n51 585
R78 B.n410 B.n409 585
R79 B.n411 B.n50 585
R80 B.n413 B.n412 585
R81 B.n414 B.n49 585
R82 B.n416 B.n415 585
R83 B.n417 B.n48 585
R84 B.n419 B.n418 585
R85 B.n420 B.n47 585
R86 B.n422 B.n421 585
R87 B.n423 B.n46 585
R88 B.n425 B.n424 585
R89 B.n426 B.n45 585
R90 B.n428 B.n427 585
R91 B.n429 B.n44 585
R92 B.n431 B.n430 585
R93 B.n432 B.n43 585
R94 B.n434 B.n433 585
R95 B.n436 B.n40 585
R96 B.n438 B.n437 585
R97 B.n439 B.n39 585
R98 B.n441 B.n440 585
R99 B.n442 B.n38 585
R100 B.n444 B.n443 585
R101 B.n445 B.n37 585
R102 B.n447 B.n446 585
R103 B.n448 B.n33 585
R104 B.n450 B.n449 585
R105 B.n451 B.n32 585
R106 B.n453 B.n452 585
R107 B.n454 B.n31 585
R108 B.n456 B.n455 585
R109 B.n457 B.n30 585
R110 B.n459 B.n458 585
R111 B.n460 B.n29 585
R112 B.n462 B.n461 585
R113 B.n463 B.n28 585
R114 B.n465 B.n464 585
R115 B.n466 B.n27 585
R116 B.n468 B.n467 585
R117 B.n469 B.n26 585
R118 B.n471 B.n470 585
R119 B.n472 B.n25 585
R120 B.n474 B.n473 585
R121 B.n475 B.n24 585
R122 B.n477 B.n476 585
R123 B.n478 B.n23 585
R124 B.n480 B.n479 585
R125 B.n481 B.n22 585
R126 B.n483 B.n482 585
R127 B.n484 B.n21 585
R128 B.n486 B.n485 585
R129 B.n487 B.n20 585
R130 B.n489 B.n488 585
R131 B.n490 B.n19 585
R132 B.n492 B.n491 585
R133 B.n493 B.n18 585
R134 B.n495 B.n494 585
R135 B.n496 B.n17 585
R136 B.n498 B.n497 585
R137 B.n499 B.n16 585
R138 B.n501 B.n500 585
R139 B.n383 B.n382 585
R140 B.n381 B.n60 585
R141 B.n380 B.n379 585
R142 B.n378 B.n61 585
R143 B.n377 B.n376 585
R144 B.n375 B.n62 585
R145 B.n374 B.n373 585
R146 B.n372 B.n63 585
R147 B.n371 B.n370 585
R148 B.n369 B.n64 585
R149 B.n368 B.n367 585
R150 B.n366 B.n65 585
R151 B.n365 B.n364 585
R152 B.n363 B.n66 585
R153 B.n362 B.n361 585
R154 B.n360 B.n67 585
R155 B.n359 B.n358 585
R156 B.n357 B.n68 585
R157 B.n356 B.n355 585
R158 B.n354 B.n69 585
R159 B.n353 B.n352 585
R160 B.n351 B.n70 585
R161 B.n350 B.n349 585
R162 B.n348 B.n71 585
R163 B.n347 B.n346 585
R164 B.n345 B.n72 585
R165 B.n344 B.n343 585
R166 B.n342 B.n73 585
R167 B.n341 B.n340 585
R168 B.n339 B.n74 585
R169 B.n338 B.n337 585
R170 B.n336 B.n75 585
R171 B.n335 B.n334 585
R172 B.n333 B.n76 585
R173 B.n332 B.n331 585
R174 B.n330 B.n77 585
R175 B.n329 B.n328 585
R176 B.n327 B.n78 585
R177 B.n326 B.n325 585
R178 B.n324 B.n79 585
R179 B.n323 B.n322 585
R180 B.n321 B.n80 585
R181 B.n320 B.n319 585
R182 B.n318 B.n81 585
R183 B.n317 B.n316 585
R184 B.n315 B.n82 585
R185 B.n314 B.n313 585
R186 B.n312 B.n83 585
R187 B.n311 B.n310 585
R188 B.n309 B.n84 585
R189 B.n308 B.n307 585
R190 B.n306 B.n85 585
R191 B.n305 B.n304 585
R192 B.n303 B.n86 585
R193 B.n302 B.n301 585
R194 B.n183 B.n130 585
R195 B.n185 B.n184 585
R196 B.n186 B.n129 585
R197 B.n188 B.n187 585
R198 B.n189 B.n128 585
R199 B.n191 B.n190 585
R200 B.n192 B.n127 585
R201 B.n194 B.n193 585
R202 B.n195 B.n126 585
R203 B.n197 B.n196 585
R204 B.n198 B.n125 585
R205 B.n200 B.n199 585
R206 B.n201 B.n124 585
R207 B.n203 B.n202 585
R208 B.n204 B.n123 585
R209 B.n206 B.n205 585
R210 B.n207 B.n122 585
R211 B.n209 B.n208 585
R212 B.n210 B.n121 585
R213 B.n212 B.n211 585
R214 B.n213 B.n120 585
R215 B.n215 B.n214 585
R216 B.n216 B.n119 585
R217 B.n218 B.n217 585
R218 B.n219 B.n118 585
R219 B.n221 B.n220 585
R220 B.n222 B.n117 585
R221 B.n224 B.n223 585
R222 B.n225 B.n116 585
R223 B.n227 B.n226 585
R224 B.n228 B.n115 585
R225 B.n230 B.n229 585
R226 B.n231 B.n114 585
R227 B.n233 B.n232 585
R228 B.n235 B.n234 585
R229 B.n236 B.n110 585
R230 B.n238 B.n237 585
R231 B.n239 B.n109 585
R232 B.n241 B.n240 585
R233 B.n242 B.n108 585
R234 B.n244 B.n243 585
R235 B.n245 B.n107 585
R236 B.n247 B.n246 585
R237 B.n248 B.n104 585
R238 B.n251 B.n250 585
R239 B.n252 B.n103 585
R240 B.n254 B.n253 585
R241 B.n255 B.n102 585
R242 B.n257 B.n256 585
R243 B.n258 B.n101 585
R244 B.n260 B.n259 585
R245 B.n261 B.n100 585
R246 B.n263 B.n262 585
R247 B.n264 B.n99 585
R248 B.n266 B.n265 585
R249 B.n267 B.n98 585
R250 B.n269 B.n268 585
R251 B.n270 B.n97 585
R252 B.n272 B.n271 585
R253 B.n273 B.n96 585
R254 B.n275 B.n274 585
R255 B.n276 B.n95 585
R256 B.n278 B.n277 585
R257 B.n279 B.n94 585
R258 B.n281 B.n280 585
R259 B.n282 B.n93 585
R260 B.n284 B.n283 585
R261 B.n285 B.n92 585
R262 B.n287 B.n286 585
R263 B.n288 B.n91 585
R264 B.n290 B.n289 585
R265 B.n291 B.n90 585
R266 B.n293 B.n292 585
R267 B.n294 B.n89 585
R268 B.n296 B.n295 585
R269 B.n297 B.n88 585
R270 B.n299 B.n298 585
R271 B.n300 B.n87 585
R272 B.n182 B.n181 585
R273 B.n180 B.n131 585
R274 B.n179 B.n178 585
R275 B.n177 B.n132 585
R276 B.n176 B.n175 585
R277 B.n174 B.n133 585
R278 B.n173 B.n172 585
R279 B.n171 B.n134 585
R280 B.n170 B.n169 585
R281 B.n168 B.n135 585
R282 B.n167 B.n166 585
R283 B.n165 B.n136 585
R284 B.n164 B.n163 585
R285 B.n162 B.n137 585
R286 B.n161 B.n160 585
R287 B.n159 B.n138 585
R288 B.n158 B.n157 585
R289 B.n156 B.n139 585
R290 B.n155 B.n154 585
R291 B.n153 B.n140 585
R292 B.n152 B.n151 585
R293 B.n150 B.n141 585
R294 B.n149 B.n148 585
R295 B.n147 B.n142 585
R296 B.n146 B.n145 585
R297 B.n144 B.n143 585
R298 B.n2 B.n0 585
R299 B.n541 B.n1 585
R300 B.n540 B.n539 585
R301 B.n538 B.n3 585
R302 B.n537 B.n536 585
R303 B.n535 B.n4 585
R304 B.n534 B.n533 585
R305 B.n532 B.n5 585
R306 B.n531 B.n530 585
R307 B.n529 B.n6 585
R308 B.n528 B.n527 585
R309 B.n526 B.n7 585
R310 B.n525 B.n524 585
R311 B.n523 B.n8 585
R312 B.n522 B.n521 585
R313 B.n520 B.n9 585
R314 B.n519 B.n518 585
R315 B.n517 B.n10 585
R316 B.n516 B.n515 585
R317 B.n514 B.n11 585
R318 B.n513 B.n512 585
R319 B.n511 B.n12 585
R320 B.n510 B.n509 585
R321 B.n508 B.n13 585
R322 B.n507 B.n506 585
R323 B.n505 B.n14 585
R324 B.n504 B.n503 585
R325 B.n502 B.n15 585
R326 B.n543 B.n542 585
R327 B.n181 B.n130 535.745
R328 B.n500 B.n15 535.745
R329 B.n301 B.n300 535.745
R330 B.n384 B.n383 535.745
R331 B.n105 B.t3 333.724
R332 B.n111 B.t6 333.724
R333 B.n34 B.t9 333.724
R334 B.n41 B.t0 333.724
R335 B.n181 B.n180 163.367
R336 B.n180 B.n179 163.367
R337 B.n179 B.n132 163.367
R338 B.n175 B.n132 163.367
R339 B.n175 B.n174 163.367
R340 B.n174 B.n173 163.367
R341 B.n173 B.n134 163.367
R342 B.n169 B.n134 163.367
R343 B.n169 B.n168 163.367
R344 B.n168 B.n167 163.367
R345 B.n167 B.n136 163.367
R346 B.n163 B.n136 163.367
R347 B.n163 B.n162 163.367
R348 B.n162 B.n161 163.367
R349 B.n161 B.n138 163.367
R350 B.n157 B.n138 163.367
R351 B.n157 B.n156 163.367
R352 B.n156 B.n155 163.367
R353 B.n155 B.n140 163.367
R354 B.n151 B.n140 163.367
R355 B.n151 B.n150 163.367
R356 B.n150 B.n149 163.367
R357 B.n149 B.n142 163.367
R358 B.n145 B.n142 163.367
R359 B.n145 B.n144 163.367
R360 B.n144 B.n2 163.367
R361 B.n542 B.n2 163.367
R362 B.n542 B.n541 163.367
R363 B.n541 B.n540 163.367
R364 B.n540 B.n3 163.367
R365 B.n536 B.n3 163.367
R366 B.n536 B.n535 163.367
R367 B.n535 B.n534 163.367
R368 B.n534 B.n5 163.367
R369 B.n530 B.n5 163.367
R370 B.n530 B.n529 163.367
R371 B.n529 B.n528 163.367
R372 B.n528 B.n7 163.367
R373 B.n524 B.n7 163.367
R374 B.n524 B.n523 163.367
R375 B.n523 B.n522 163.367
R376 B.n522 B.n9 163.367
R377 B.n518 B.n9 163.367
R378 B.n518 B.n517 163.367
R379 B.n517 B.n516 163.367
R380 B.n516 B.n11 163.367
R381 B.n512 B.n11 163.367
R382 B.n512 B.n511 163.367
R383 B.n511 B.n510 163.367
R384 B.n510 B.n13 163.367
R385 B.n506 B.n13 163.367
R386 B.n506 B.n505 163.367
R387 B.n505 B.n504 163.367
R388 B.n504 B.n15 163.367
R389 B.n185 B.n130 163.367
R390 B.n186 B.n185 163.367
R391 B.n187 B.n186 163.367
R392 B.n187 B.n128 163.367
R393 B.n191 B.n128 163.367
R394 B.n192 B.n191 163.367
R395 B.n193 B.n192 163.367
R396 B.n193 B.n126 163.367
R397 B.n197 B.n126 163.367
R398 B.n198 B.n197 163.367
R399 B.n199 B.n198 163.367
R400 B.n199 B.n124 163.367
R401 B.n203 B.n124 163.367
R402 B.n204 B.n203 163.367
R403 B.n205 B.n204 163.367
R404 B.n205 B.n122 163.367
R405 B.n209 B.n122 163.367
R406 B.n210 B.n209 163.367
R407 B.n211 B.n210 163.367
R408 B.n211 B.n120 163.367
R409 B.n215 B.n120 163.367
R410 B.n216 B.n215 163.367
R411 B.n217 B.n216 163.367
R412 B.n217 B.n118 163.367
R413 B.n221 B.n118 163.367
R414 B.n222 B.n221 163.367
R415 B.n223 B.n222 163.367
R416 B.n223 B.n116 163.367
R417 B.n227 B.n116 163.367
R418 B.n228 B.n227 163.367
R419 B.n229 B.n228 163.367
R420 B.n229 B.n114 163.367
R421 B.n233 B.n114 163.367
R422 B.n234 B.n233 163.367
R423 B.n234 B.n110 163.367
R424 B.n238 B.n110 163.367
R425 B.n239 B.n238 163.367
R426 B.n240 B.n239 163.367
R427 B.n240 B.n108 163.367
R428 B.n244 B.n108 163.367
R429 B.n245 B.n244 163.367
R430 B.n246 B.n245 163.367
R431 B.n246 B.n104 163.367
R432 B.n251 B.n104 163.367
R433 B.n252 B.n251 163.367
R434 B.n253 B.n252 163.367
R435 B.n253 B.n102 163.367
R436 B.n257 B.n102 163.367
R437 B.n258 B.n257 163.367
R438 B.n259 B.n258 163.367
R439 B.n259 B.n100 163.367
R440 B.n263 B.n100 163.367
R441 B.n264 B.n263 163.367
R442 B.n265 B.n264 163.367
R443 B.n265 B.n98 163.367
R444 B.n269 B.n98 163.367
R445 B.n270 B.n269 163.367
R446 B.n271 B.n270 163.367
R447 B.n271 B.n96 163.367
R448 B.n275 B.n96 163.367
R449 B.n276 B.n275 163.367
R450 B.n277 B.n276 163.367
R451 B.n277 B.n94 163.367
R452 B.n281 B.n94 163.367
R453 B.n282 B.n281 163.367
R454 B.n283 B.n282 163.367
R455 B.n283 B.n92 163.367
R456 B.n287 B.n92 163.367
R457 B.n288 B.n287 163.367
R458 B.n289 B.n288 163.367
R459 B.n289 B.n90 163.367
R460 B.n293 B.n90 163.367
R461 B.n294 B.n293 163.367
R462 B.n295 B.n294 163.367
R463 B.n295 B.n88 163.367
R464 B.n299 B.n88 163.367
R465 B.n300 B.n299 163.367
R466 B.n301 B.n86 163.367
R467 B.n305 B.n86 163.367
R468 B.n306 B.n305 163.367
R469 B.n307 B.n306 163.367
R470 B.n307 B.n84 163.367
R471 B.n311 B.n84 163.367
R472 B.n312 B.n311 163.367
R473 B.n313 B.n312 163.367
R474 B.n313 B.n82 163.367
R475 B.n317 B.n82 163.367
R476 B.n318 B.n317 163.367
R477 B.n319 B.n318 163.367
R478 B.n319 B.n80 163.367
R479 B.n323 B.n80 163.367
R480 B.n324 B.n323 163.367
R481 B.n325 B.n324 163.367
R482 B.n325 B.n78 163.367
R483 B.n329 B.n78 163.367
R484 B.n330 B.n329 163.367
R485 B.n331 B.n330 163.367
R486 B.n331 B.n76 163.367
R487 B.n335 B.n76 163.367
R488 B.n336 B.n335 163.367
R489 B.n337 B.n336 163.367
R490 B.n337 B.n74 163.367
R491 B.n341 B.n74 163.367
R492 B.n342 B.n341 163.367
R493 B.n343 B.n342 163.367
R494 B.n343 B.n72 163.367
R495 B.n347 B.n72 163.367
R496 B.n348 B.n347 163.367
R497 B.n349 B.n348 163.367
R498 B.n349 B.n70 163.367
R499 B.n353 B.n70 163.367
R500 B.n354 B.n353 163.367
R501 B.n355 B.n354 163.367
R502 B.n355 B.n68 163.367
R503 B.n359 B.n68 163.367
R504 B.n360 B.n359 163.367
R505 B.n361 B.n360 163.367
R506 B.n361 B.n66 163.367
R507 B.n365 B.n66 163.367
R508 B.n366 B.n365 163.367
R509 B.n367 B.n366 163.367
R510 B.n367 B.n64 163.367
R511 B.n371 B.n64 163.367
R512 B.n372 B.n371 163.367
R513 B.n373 B.n372 163.367
R514 B.n373 B.n62 163.367
R515 B.n377 B.n62 163.367
R516 B.n378 B.n377 163.367
R517 B.n379 B.n378 163.367
R518 B.n379 B.n60 163.367
R519 B.n383 B.n60 163.367
R520 B.n500 B.n499 163.367
R521 B.n499 B.n498 163.367
R522 B.n498 B.n17 163.367
R523 B.n494 B.n17 163.367
R524 B.n494 B.n493 163.367
R525 B.n493 B.n492 163.367
R526 B.n492 B.n19 163.367
R527 B.n488 B.n19 163.367
R528 B.n488 B.n487 163.367
R529 B.n487 B.n486 163.367
R530 B.n486 B.n21 163.367
R531 B.n482 B.n21 163.367
R532 B.n482 B.n481 163.367
R533 B.n481 B.n480 163.367
R534 B.n480 B.n23 163.367
R535 B.n476 B.n23 163.367
R536 B.n476 B.n475 163.367
R537 B.n475 B.n474 163.367
R538 B.n474 B.n25 163.367
R539 B.n470 B.n25 163.367
R540 B.n470 B.n469 163.367
R541 B.n469 B.n468 163.367
R542 B.n468 B.n27 163.367
R543 B.n464 B.n27 163.367
R544 B.n464 B.n463 163.367
R545 B.n463 B.n462 163.367
R546 B.n462 B.n29 163.367
R547 B.n458 B.n29 163.367
R548 B.n458 B.n457 163.367
R549 B.n457 B.n456 163.367
R550 B.n456 B.n31 163.367
R551 B.n452 B.n31 163.367
R552 B.n452 B.n451 163.367
R553 B.n451 B.n450 163.367
R554 B.n450 B.n33 163.367
R555 B.n446 B.n33 163.367
R556 B.n446 B.n445 163.367
R557 B.n445 B.n444 163.367
R558 B.n444 B.n38 163.367
R559 B.n440 B.n38 163.367
R560 B.n440 B.n439 163.367
R561 B.n439 B.n438 163.367
R562 B.n438 B.n40 163.367
R563 B.n433 B.n40 163.367
R564 B.n433 B.n432 163.367
R565 B.n432 B.n431 163.367
R566 B.n431 B.n44 163.367
R567 B.n427 B.n44 163.367
R568 B.n427 B.n426 163.367
R569 B.n426 B.n425 163.367
R570 B.n425 B.n46 163.367
R571 B.n421 B.n46 163.367
R572 B.n421 B.n420 163.367
R573 B.n420 B.n419 163.367
R574 B.n419 B.n48 163.367
R575 B.n415 B.n48 163.367
R576 B.n415 B.n414 163.367
R577 B.n414 B.n413 163.367
R578 B.n413 B.n50 163.367
R579 B.n409 B.n50 163.367
R580 B.n409 B.n408 163.367
R581 B.n408 B.n407 163.367
R582 B.n407 B.n52 163.367
R583 B.n403 B.n52 163.367
R584 B.n403 B.n402 163.367
R585 B.n402 B.n401 163.367
R586 B.n401 B.n54 163.367
R587 B.n397 B.n54 163.367
R588 B.n397 B.n396 163.367
R589 B.n396 B.n395 163.367
R590 B.n395 B.n56 163.367
R591 B.n391 B.n56 163.367
R592 B.n391 B.n390 163.367
R593 B.n390 B.n389 163.367
R594 B.n389 B.n58 163.367
R595 B.n385 B.n58 163.367
R596 B.n385 B.n384 163.367
R597 B.n105 B.t5 150.119
R598 B.n41 B.t1 150.119
R599 B.n111 B.t8 150.107
R600 B.n34 B.t10 150.107
R601 B.n106 B.t4 108.615
R602 B.n42 B.t2 108.615
R603 B.n112 B.t7 108.605
R604 B.n35 B.t11 108.605
R605 B.n249 B.n106 59.5399
R606 B.n113 B.n112 59.5399
R607 B.n36 B.n35 59.5399
R608 B.n435 B.n42 59.5399
R609 B.n106 B.n105 41.5035
R610 B.n112 B.n111 41.5035
R611 B.n35 B.n34 41.5035
R612 B.n42 B.n41 41.5035
R613 B.n502 B.n501 34.8103
R614 B.n382 B.n59 34.8103
R615 B.n302 B.n87 34.8103
R616 B.n183 B.n182 34.8103
R617 B B.n543 18.0485
R618 B.n501 B.n16 10.6151
R619 B.n497 B.n16 10.6151
R620 B.n497 B.n496 10.6151
R621 B.n496 B.n495 10.6151
R622 B.n495 B.n18 10.6151
R623 B.n491 B.n18 10.6151
R624 B.n491 B.n490 10.6151
R625 B.n490 B.n489 10.6151
R626 B.n489 B.n20 10.6151
R627 B.n485 B.n20 10.6151
R628 B.n485 B.n484 10.6151
R629 B.n484 B.n483 10.6151
R630 B.n483 B.n22 10.6151
R631 B.n479 B.n22 10.6151
R632 B.n479 B.n478 10.6151
R633 B.n478 B.n477 10.6151
R634 B.n477 B.n24 10.6151
R635 B.n473 B.n24 10.6151
R636 B.n473 B.n472 10.6151
R637 B.n472 B.n471 10.6151
R638 B.n471 B.n26 10.6151
R639 B.n467 B.n26 10.6151
R640 B.n467 B.n466 10.6151
R641 B.n466 B.n465 10.6151
R642 B.n465 B.n28 10.6151
R643 B.n461 B.n28 10.6151
R644 B.n461 B.n460 10.6151
R645 B.n460 B.n459 10.6151
R646 B.n459 B.n30 10.6151
R647 B.n455 B.n30 10.6151
R648 B.n455 B.n454 10.6151
R649 B.n454 B.n453 10.6151
R650 B.n453 B.n32 10.6151
R651 B.n449 B.n448 10.6151
R652 B.n448 B.n447 10.6151
R653 B.n447 B.n37 10.6151
R654 B.n443 B.n37 10.6151
R655 B.n443 B.n442 10.6151
R656 B.n442 B.n441 10.6151
R657 B.n441 B.n39 10.6151
R658 B.n437 B.n39 10.6151
R659 B.n437 B.n436 10.6151
R660 B.n434 B.n43 10.6151
R661 B.n430 B.n43 10.6151
R662 B.n430 B.n429 10.6151
R663 B.n429 B.n428 10.6151
R664 B.n428 B.n45 10.6151
R665 B.n424 B.n45 10.6151
R666 B.n424 B.n423 10.6151
R667 B.n423 B.n422 10.6151
R668 B.n422 B.n47 10.6151
R669 B.n418 B.n47 10.6151
R670 B.n418 B.n417 10.6151
R671 B.n417 B.n416 10.6151
R672 B.n416 B.n49 10.6151
R673 B.n412 B.n49 10.6151
R674 B.n412 B.n411 10.6151
R675 B.n411 B.n410 10.6151
R676 B.n410 B.n51 10.6151
R677 B.n406 B.n51 10.6151
R678 B.n406 B.n405 10.6151
R679 B.n405 B.n404 10.6151
R680 B.n404 B.n53 10.6151
R681 B.n400 B.n53 10.6151
R682 B.n400 B.n399 10.6151
R683 B.n399 B.n398 10.6151
R684 B.n398 B.n55 10.6151
R685 B.n394 B.n55 10.6151
R686 B.n394 B.n393 10.6151
R687 B.n393 B.n392 10.6151
R688 B.n392 B.n57 10.6151
R689 B.n388 B.n57 10.6151
R690 B.n388 B.n387 10.6151
R691 B.n387 B.n386 10.6151
R692 B.n386 B.n59 10.6151
R693 B.n303 B.n302 10.6151
R694 B.n304 B.n303 10.6151
R695 B.n304 B.n85 10.6151
R696 B.n308 B.n85 10.6151
R697 B.n309 B.n308 10.6151
R698 B.n310 B.n309 10.6151
R699 B.n310 B.n83 10.6151
R700 B.n314 B.n83 10.6151
R701 B.n315 B.n314 10.6151
R702 B.n316 B.n315 10.6151
R703 B.n316 B.n81 10.6151
R704 B.n320 B.n81 10.6151
R705 B.n321 B.n320 10.6151
R706 B.n322 B.n321 10.6151
R707 B.n322 B.n79 10.6151
R708 B.n326 B.n79 10.6151
R709 B.n327 B.n326 10.6151
R710 B.n328 B.n327 10.6151
R711 B.n328 B.n77 10.6151
R712 B.n332 B.n77 10.6151
R713 B.n333 B.n332 10.6151
R714 B.n334 B.n333 10.6151
R715 B.n334 B.n75 10.6151
R716 B.n338 B.n75 10.6151
R717 B.n339 B.n338 10.6151
R718 B.n340 B.n339 10.6151
R719 B.n340 B.n73 10.6151
R720 B.n344 B.n73 10.6151
R721 B.n345 B.n344 10.6151
R722 B.n346 B.n345 10.6151
R723 B.n346 B.n71 10.6151
R724 B.n350 B.n71 10.6151
R725 B.n351 B.n350 10.6151
R726 B.n352 B.n351 10.6151
R727 B.n352 B.n69 10.6151
R728 B.n356 B.n69 10.6151
R729 B.n357 B.n356 10.6151
R730 B.n358 B.n357 10.6151
R731 B.n358 B.n67 10.6151
R732 B.n362 B.n67 10.6151
R733 B.n363 B.n362 10.6151
R734 B.n364 B.n363 10.6151
R735 B.n364 B.n65 10.6151
R736 B.n368 B.n65 10.6151
R737 B.n369 B.n368 10.6151
R738 B.n370 B.n369 10.6151
R739 B.n370 B.n63 10.6151
R740 B.n374 B.n63 10.6151
R741 B.n375 B.n374 10.6151
R742 B.n376 B.n375 10.6151
R743 B.n376 B.n61 10.6151
R744 B.n380 B.n61 10.6151
R745 B.n381 B.n380 10.6151
R746 B.n382 B.n381 10.6151
R747 B.n184 B.n183 10.6151
R748 B.n184 B.n129 10.6151
R749 B.n188 B.n129 10.6151
R750 B.n189 B.n188 10.6151
R751 B.n190 B.n189 10.6151
R752 B.n190 B.n127 10.6151
R753 B.n194 B.n127 10.6151
R754 B.n195 B.n194 10.6151
R755 B.n196 B.n195 10.6151
R756 B.n196 B.n125 10.6151
R757 B.n200 B.n125 10.6151
R758 B.n201 B.n200 10.6151
R759 B.n202 B.n201 10.6151
R760 B.n202 B.n123 10.6151
R761 B.n206 B.n123 10.6151
R762 B.n207 B.n206 10.6151
R763 B.n208 B.n207 10.6151
R764 B.n208 B.n121 10.6151
R765 B.n212 B.n121 10.6151
R766 B.n213 B.n212 10.6151
R767 B.n214 B.n213 10.6151
R768 B.n214 B.n119 10.6151
R769 B.n218 B.n119 10.6151
R770 B.n219 B.n218 10.6151
R771 B.n220 B.n219 10.6151
R772 B.n220 B.n117 10.6151
R773 B.n224 B.n117 10.6151
R774 B.n225 B.n224 10.6151
R775 B.n226 B.n225 10.6151
R776 B.n226 B.n115 10.6151
R777 B.n230 B.n115 10.6151
R778 B.n231 B.n230 10.6151
R779 B.n232 B.n231 10.6151
R780 B.n236 B.n235 10.6151
R781 B.n237 B.n236 10.6151
R782 B.n237 B.n109 10.6151
R783 B.n241 B.n109 10.6151
R784 B.n242 B.n241 10.6151
R785 B.n243 B.n242 10.6151
R786 B.n243 B.n107 10.6151
R787 B.n247 B.n107 10.6151
R788 B.n248 B.n247 10.6151
R789 B.n250 B.n103 10.6151
R790 B.n254 B.n103 10.6151
R791 B.n255 B.n254 10.6151
R792 B.n256 B.n255 10.6151
R793 B.n256 B.n101 10.6151
R794 B.n260 B.n101 10.6151
R795 B.n261 B.n260 10.6151
R796 B.n262 B.n261 10.6151
R797 B.n262 B.n99 10.6151
R798 B.n266 B.n99 10.6151
R799 B.n267 B.n266 10.6151
R800 B.n268 B.n267 10.6151
R801 B.n268 B.n97 10.6151
R802 B.n272 B.n97 10.6151
R803 B.n273 B.n272 10.6151
R804 B.n274 B.n273 10.6151
R805 B.n274 B.n95 10.6151
R806 B.n278 B.n95 10.6151
R807 B.n279 B.n278 10.6151
R808 B.n280 B.n279 10.6151
R809 B.n280 B.n93 10.6151
R810 B.n284 B.n93 10.6151
R811 B.n285 B.n284 10.6151
R812 B.n286 B.n285 10.6151
R813 B.n286 B.n91 10.6151
R814 B.n290 B.n91 10.6151
R815 B.n291 B.n290 10.6151
R816 B.n292 B.n291 10.6151
R817 B.n292 B.n89 10.6151
R818 B.n296 B.n89 10.6151
R819 B.n297 B.n296 10.6151
R820 B.n298 B.n297 10.6151
R821 B.n298 B.n87 10.6151
R822 B.n182 B.n131 10.6151
R823 B.n178 B.n131 10.6151
R824 B.n178 B.n177 10.6151
R825 B.n177 B.n176 10.6151
R826 B.n176 B.n133 10.6151
R827 B.n172 B.n133 10.6151
R828 B.n172 B.n171 10.6151
R829 B.n171 B.n170 10.6151
R830 B.n170 B.n135 10.6151
R831 B.n166 B.n135 10.6151
R832 B.n166 B.n165 10.6151
R833 B.n165 B.n164 10.6151
R834 B.n164 B.n137 10.6151
R835 B.n160 B.n137 10.6151
R836 B.n160 B.n159 10.6151
R837 B.n159 B.n158 10.6151
R838 B.n158 B.n139 10.6151
R839 B.n154 B.n139 10.6151
R840 B.n154 B.n153 10.6151
R841 B.n153 B.n152 10.6151
R842 B.n152 B.n141 10.6151
R843 B.n148 B.n141 10.6151
R844 B.n148 B.n147 10.6151
R845 B.n147 B.n146 10.6151
R846 B.n146 B.n143 10.6151
R847 B.n143 B.n0 10.6151
R848 B.n539 B.n1 10.6151
R849 B.n539 B.n538 10.6151
R850 B.n538 B.n537 10.6151
R851 B.n537 B.n4 10.6151
R852 B.n533 B.n4 10.6151
R853 B.n533 B.n532 10.6151
R854 B.n532 B.n531 10.6151
R855 B.n531 B.n6 10.6151
R856 B.n527 B.n6 10.6151
R857 B.n527 B.n526 10.6151
R858 B.n526 B.n525 10.6151
R859 B.n525 B.n8 10.6151
R860 B.n521 B.n8 10.6151
R861 B.n521 B.n520 10.6151
R862 B.n520 B.n519 10.6151
R863 B.n519 B.n10 10.6151
R864 B.n515 B.n10 10.6151
R865 B.n515 B.n514 10.6151
R866 B.n514 B.n513 10.6151
R867 B.n513 B.n12 10.6151
R868 B.n509 B.n12 10.6151
R869 B.n509 B.n508 10.6151
R870 B.n508 B.n507 10.6151
R871 B.n507 B.n14 10.6151
R872 B.n503 B.n14 10.6151
R873 B.n503 B.n502 10.6151
R874 B.n36 B.n32 9.36635
R875 B.n435 B.n434 9.36635
R876 B.n232 B.n113 9.36635
R877 B.n250 B.n249 9.36635
R878 B.n543 B.n0 2.81026
R879 B.n543 B.n1 2.81026
R880 B.n449 B.n36 1.24928
R881 B.n436 B.n435 1.24928
R882 B.n235 B.n113 1.24928
R883 B.n249 B.n248 1.24928
C0 VP VTAIL 3.48509f
C1 VN B 0.92707f
C2 w_n2254_n2880# B 7.589479f
C3 VDD2 VN 3.57088f
C4 VDD2 w_n2254_n2880# 1.26863f
C5 B VDD1 1.0574f
C6 VN VTAIL 3.47098f
C7 w_n2254_n2880# VTAIL 3.40995f
C8 VP VN 5.17239f
C9 VP w_n2254_n2880# 3.91791f
C10 VDD2 VDD1 0.834274f
C11 VTAIL VDD1 4.73884f
C12 VP VDD1 3.76609f
C13 VDD2 B 1.09663f
C14 w_n2254_n2880# VN 3.63015f
C15 B VTAIL 3.79731f
C16 VP B 1.40092f
C17 VN VDD1 0.147774f
C18 VDD2 VTAIL 4.78775f
C19 w_n2254_n2880# VDD1 1.23018f
C20 VP VDD2 0.343524f
C21 VDD2 VSUBS 0.764084f
C22 VDD1 VSUBS 4.959923f
C23 VTAIL VSUBS 0.99564f
C24 VN VSUBS 5.083529f
C25 VP VSUBS 1.76448f
C26 B VSUBS 3.385417f
C27 w_n2254_n2880# VSUBS 80.251396f
C28 B.n0 VSUBS 0.00483f
C29 B.n1 VSUBS 0.00483f
C30 B.n2 VSUBS 0.007638f
C31 B.n3 VSUBS 0.007638f
C32 B.n4 VSUBS 0.007638f
C33 B.n5 VSUBS 0.007638f
C34 B.n6 VSUBS 0.007638f
C35 B.n7 VSUBS 0.007638f
C36 B.n8 VSUBS 0.007638f
C37 B.n9 VSUBS 0.007638f
C38 B.n10 VSUBS 0.007638f
C39 B.n11 VSUBS 0.007638f
C40 B.n12 VSUBS 0.007638f
C41 B.n13 VSUBS 0.007638f
C42 B.n14 VSUBS 0.007638f
C43 B.n15 VSUBS 0.018407f
C44 B.n16 VSUBS 0.007638f
C45 B.n17 VSUBS 0.007638f
C46 B.n18 VSUBS 0.007638f
C47 B.n19 VSUBS 0.007638f
C48 B.n20 VSUBS 0.007638f
C49 B.n21 VSUBS 0.007638f
C50 B.n22 VSUBS 0.007638f
C51 B.n23 VSUBS 0.007638f
C52 B.n24 VSUBS 0.007638f
C53 B.n25 VSUBS 0.007638f
C54 B.n26 VSUBS 0.007638f
C55 B.n27 VSUBS 0.007638f
C56 B.n28 VSUBS 0.007638f
C57 B.n29 VSUBS 0.007638f
C58 B.n30 VSUBS 0.007638f
C59 B.n31 VSUBS 0.007638f
C60 B.n32 VSUBS 0.007188f
C61 B.n33 VSUBS 0.007638f
C62 B.t11 VSUBS 0.330666f
C63 B.t10 VSUBS 0.348261f
C64 B.t9 VSUBS 0.850652f
C65 B.n34 VSUBS 0.168756f
C66 B.n35 VSUBS 0.07453f
C67 B.n36 VSUBS 0.017696f
C68 B.n37 VSUBS 0.007638f
C69 B.n38 VSUBS 0.007638f
C70 B.n39 VSUBS 0.007638f
C71 B.n40 VSUBS 0.007638f
C72 B.t2 VSUBS 0.330662f
C73 B.t1 VSUBS 0.348256f
C74 B.t0 VSUBS 0.850652f
C75 B.n41 VSUBS 0.16876f
C76 B.n42 VSUBS 0.074534f
C77 B.n43 VSUBS 0.007638f
C78 B.n44 VSUBS 0.007638f
C79 B.n45 VSUBS 0.007638f
C80 B.n46 VSUBS 0.007638f
C81 B.n47 VSUBS 0.007638f
C82 B.n48 VSUBS 0.007638f
C83 B.n49 VSUBS 0.007638f
C84 B.n50 VSUBS 0.007638f
C85 B.n51 VSUBS 0.007638f
C86 B.n52 VSUBS 0.007638f
C87 B.n53 VSUBS 0.007638f
C88 B.n54 VSUBS 0.007638f
C89 B.n55 VSUBS 0.007638f
C90 B.n56 VSUBS 0.007638f
C91 B.n57 VSUBS 0.007638f
C92 B.n58 VSUBS 0.007638f
C93 B.n59 VSUBS 0.018036f
C94 B.n60 VSUBS 0.007638f
C95 B.n61 VSUBS 0.007638f
C96 B.n62 VSUBS 0.007638f
C97 B.n63 VSUBS 0.007638f
C98 B.n64 VSUBS 0.007638f
C99 B.n65 VSUBS 0.007638f
C100 B.n66 VSUBS 0.007638f
C101 B.n67 VSUBS 0.007638f
C102 B.n68 VSUBS 0.007638f
C103 B.n69 VSUBS 0.007638f
C104 B.n70 VSUBS 0.007638f
C105 B.n71 VSUBS 0.007638f
C106 B.n72 VSUBS 0.007638f
C107 B.n73 VSUBS 0.007638f
C108 B.n74 VSUBS 0.007638f
C109 B.n75 VSUBS 0.007638f
C110 B.n76 VSUBS 0.007638f
C111 B.n77 VSUBS 0.007638f
C112 B.n78 VSUBS 0.007638f
C113 B.n79 VSUBS 0.007638f
C114 B.n80 VSUBS 0.007638f
C115 B.n81 VSUBS 0.007638f
C116 B.n82 VSUBS 0.007638f
C117 B.n83 VSUBS 0.007638f
C118 B.n84 VSUBS 0.007638f
C119 B.n85 VSUBS 0.007638f
C120 B.n86 VSUBS 0.007638f
C121 B.n87 VSUBS 0.018882f
C122 B.n88 VSUBS 0.007638f
C123 B.n89 VSUBS 0.007638f
C124 B.n90 VSUBS 0.007638f
C125 B.n91 VSUBS 0.007638f
C126 B.n92 VSUBS 0.007638f
C127 B.n93 VSUBS 0.007638f
C128 B.n94 VSUBS 0.007638f
C129 B.n95 VSUBS 0.007638f
C130 B.n96 VSUBS 0.007638f
C131 B.n97 VSUBS 0.007638f
C132 B.n98 VSUBS 0.007638f
C133 B.n99 VSUBS 0.007638f
C134 B.n100 VSUBS 0.007638f
C135 B.n101 VSUBS 0.007638f
C136 B.n102 VSUBS 0.007638f
C137 B.n103 VSUBS 0.007638f
C138 B.n104 VSUBS 0.007638f
C139 B.t4 VSUBS 0.330662f
C140 B.t5 VSUBS 0.348256f
C141 B.t3 VSUBS 0.850652f
C142 B.n105 VSUBS 0.16876f
C143 B.n106 VSUBS 0.074534f
C144 B.n107 VSUBS 0.007638f
C145 B.n108 VSUBS 0.007638f
C146 B.n109 VSUBS 0.007638f
C147 B.n110 VSUBS 0.007638f
C148 B.t7 VSUBS 0.330666f
C149 B.t8 VSUBS 0.348261f
C150 B.t6 VSUBS 0.850652f
C151 B.n111 VSUBS 0.168756f
C152 B.n112 VSUBS 0.07453f
C153 B.n113 VSUBS 0.017696f
C154 B.n114 VSUBS 0.007638f
C155 B.n115 VSUBS 0.007638f
C156 B.n116 VSUBS 0.007638f
C157 B.n117 VSUBS 0.007638f
C158 B.n118 VSUBS 0.007638f
C159 B.n119 VSUBS 0.007638f
C160 B.n120 VSUBS 0.007638f
C161 B.n121 VSUBS 0.007638f
C162 B.n122 VSUBS 0.007638f
C163 B.n123 VSUBS 0.007638f
C164 B.n124 VSUBS 0.007638f
C165 B.n125 VSUBS 0.007638f
C166 B.n126 VSUBS 0.007638f
C167 B.n127 VSUBS 0.007638f
C168 B.n128 VSUBS 0.007638f
C169 B.n129 VSUBS 0.007638f
C170 B.n130 VSUBS 0.018882f
C171 B.n131 VSUBS 0.007638f
C172 B.n132 VSUBS 0.007638f
C173 B.n133 VSUBS 0.007638f
C174 B.n134 VSUBS 0.007638f
C175 B.n135 VSUBS 0.007638f
C176 B.n136 VSUBS 0.007638f
C177 B.n137 VSUBS 0.007638f
C178 B.n138 VSUBS 0.007638f
C179 B.n139 VSUBS 0.007638f
C180 B.n140 VSUBS 0.007638f
C181 B.n141 VSUBS 0.007638f
C182 B.n142 VSUBS 0.007638f
C183 B.n143 VSUBS 0.007638f
C184 B.n144 VSUBS 0.007638f
C185 B.n145 VSUBS 0.007638f
C186 B.n146 VSUBS 0.007638f
C187 B.n147 VSUBS 0.007638f
C188 B.n148 VSUBS 0.007638f
C189 B.n149 VSUBS 0.007638f
C190 B.n150 VSUBS 0.007638f
C191 B.n151 VSUBS 0.007638f
C192 B.n152 VSUBS 0.007638f
C193 B.n153 VSUBS 0.007638f
C194 B.n154 VSUBS 0.007638f
C195 B.n155 VSUBS 0.007638f
C196 B.n156 VSUBS 0.007638f
C197 B.n157 VSUBS 0.007638f
C198 B.n158 VSUBS 0.007638f
C199 B.n159 VSUBS 0.007638f
C200 B.n160 VSUBS 0.007638f
C201 B.n161 VSUBS 0.007638f
C202 B.n162 VSUBS 0.007638f
C203 B.n163 VSUBS 0.007638f
C204 B.n164 VSUBS 0.007638f
C205 B.n165 VSUBS 0.007638f
C206 B.n166 VSUBS 0.007638f
C207 B.n167 VSUBS 0.007638f
C208 B.n168 VSUBS 0.007638f
C209 B.n169 VSUBS 0.007638f
C210 B.n170 VSUBS 0.007638f
C211 B.n171 VSUBS 0.007638f
C212 B.n172 VSUBS 0.007638f
C213 B.n173 VSUBS 0.007638f
C214 B.n174 VSUBS 0.007638f
C215 B.n175 VSUBS 0.007638f
C216 B.n176 VSUBS 0.007638f
C217 B.n177 VSUBS 0.007638f
C218 B.n178 VSUBS 0.007638f
C219 B.n179 VSUBS 0.007638f
C220 B.n180 VSUBS 0.007638f
C221 B.n181 VSUBS 0.018407f
C222 B.n182 VSUBS 0.018407f
C223 B.n183 VSUBS 0.018882f
C224 B.n184 VSUBS 0.007638f
C225 B.n185 VSUBS 0.007638f
C226 B.n186 VSUBS 0.007638f
C227 B.n187 VSUBS 0.007638f
C228 B.n188 VSUBS 0.007638f
C229 B.n189 VSUBS 0.007638f
C230 B.n190 VSUBS 0.007638f
C231 B.n191 VSUBS 0.007638f
C232 B.n192 VSUBS 0.007638f
C233 B.n193 VSUBS 0.007638f
C234 B.n194 VSUBS 0.007638f
C235 B.n195 VSUBS 0.007638f
C236 B.n196 VSUBS 0.007638f
C237 B.n197 VSUBS 0.007638f
C238 B.n198 VSUBS 0.007638f
C239 B.n199 VSUBS 0.007638f
C240 B.n200 VSUBS 0.007638f
C241 B.n201 VSUBS 0.007638f
C242 B.n202 VSUBS 0.007638f
C243 B.n203 VSUBS 0.007638f
C244 B.n204 VSUBS 0.007638f
C245 B.n205 VSUBS 0.007638f
C246 B.n206 VSUBS 0.007638f
C247 B.n207 VSUBS 0.007638f
C248 B.n208 VSUBS 0.007638f
C249 B.n209 VSUBS 0.007638f
C250 B.n210 VSUBS 0.007638f
C251 B.n211 VSUBS 0.007638f
C252 B.n212 VSUBS 0.007638f
C253 B.n213 VSUBS 0.007638f
C254 B.n214 VSUBS 0.007638f
C255 B.n215 VSUBS 0.007638f
C256 B.n216 VSUBS 0.007638f
C257 B.n217 VSUBS 0.007638f
C258 B.n218 VSUBS 0.007638f
C259 B.n219 VSUBS 0.007638f
C260 B.n220 VSUBS 0.007638f
C261 B.n221 VSUBS 0.007638f
C262 B.n222 VSUBS 0.007638f
C263 B.n223 VSUBS 0.007638f
C264 B.n224 VSUBS 0.007638f
C265 B.n225 VSUBS 0.007638f
C266 B.n226 VSUBS 0.007638f
C267 B.n227 VSUBS 0.007638f
C268 B.n228 VSUBS 0.007638f
C269 B.n229 VSUBS 0.007638f
C270 B.n230 VSUBS 0.007638f
C271 B.n231 VSUBS 0.007638f
C272 B.n232 VSUBS 0.007188f
C273 B.n233 VSUBS 0.007638f
C274 B.n234 VSUBS 0.007638f
C275 B.n235 VSUBS 0.004268f
C276 B.n236 VSUBS 0.007638f
C277 B.n237 VSUBS 0.007638f
C278 B.n238 VSUBS 0.007638f
C279 B.n239 VSUBS 0.007638f
C280 B.n240 VSUBS 0.007638f
C281 B.n241 VSUBS 0.007638f
C282 B.n242 VSUBS 0.007638f
C283 B.n243 VSUBS 0.007638f
C284 B.n244 VSUBS 0.007638f
C285 B.n245 VSUBS 0.007638f
C286 B.n246 VSUBS 0.007638f
C287 B.n247 VSUBS 0.007638f
C288 B.n248 VSUBS 0.004268f
C289 B.n249 VSUBS 0.017696f
C290 B.n250 VSUBS 0.007188f
C291 B.n251 VSUBS 0.007638f
C292 B.n252 VSUBS 0.007638f
C293 B.n253 VSUBS 0.007638f
C294 B.n254 VSUBS 0.007638f
C295 B.n255 VSUBS 0.007638f
C296 B.n256 VSUBS 0.007638f
C297 B.n257 VSUBS 0.007638f
C298 B.n258 VSUBS 0.007638f
C299 B.n259 VSUBS 0.007638f
C300 B.n260 VSUBS 0.007638f
C301 B.n261 VSUBS 0.007638f
C302 B.n262 VSUBS 0.007638f
C303 B.n263 VSUBS 0.007638f
C304 B.n264 VSUBS 0.007638f
C305 B.n265 VSUBS 0.007638f
C306 B.n266 VSUBS 0.007638f
C307 B.n267 VSUBS 0.007638f
C308 B.n268 VSUBS 0.007638f
C309 B.n269 VSUBS 0.007638f
C310 B.n270 VSUBS 0.007638f
C311 B.n271 VSUBS 0.007638f
C312 B.n272 VSUBS 0.007638f
C313 B.n273 VSUBS 0.007638f
C314 B.n274 VSUBS 0.007638f
C315 B.n275 VSUBS 0.007638f
C316 B.n276 VSUBS 0.007638f
C317 B.n277 VSUBS 0.007638f
C318 B.n278 VSUBS 0.007638f
C319 B.n279 VSUBS 0.007638f
C320 B.n280 VSUBS 0.007638f
C321 B.n281 VSUBS 0.007638f
C322 B.n282 VSUBS 0.007638f
C323 B.n283 VSUBS 0.007638f
C324 B.n284 VSUBS 0.007638f
C325 B.n285 VSUBS 0.007638f
C326 B.n286 VSUBS 0.007638f
C327 B.n287 VSUBS 0.007638f
C328 B.n288 VSUBS 0.007638f
C329 B.n289 VSUBS 0.007638f
C330 B.n290 VSUBS 0.007638f
C331 B.n291 VSUBS 0.007638f
C332 B.n292 VSUBS 0.007638f
C333 B.n293 VSUBS 0.007638f
C334 B.n294 VSUBS 0.007638f
C335 B.n295 VSUBS 0.007638f
C336 B.n296 VSUBS 0.007638f
C337 B.n297 VSUBS 0.007638f
C338 B.n298 VSUBS 0.007638f
C339 B.n299 VSUBS 0.007638f
C340 B.n300 VSUBS 0.018882f
C341 B.n301 VSUBS 0.018407f
C342 B.n302 VSUBS 0.018407f
C343 B.n303 VSUBS 0.007638f
C344 B.n304 VSUBS 0.007638f
C345 B.n305 VSUBS 0.007638f
C346 B.n306 VSUBS 0.007638f
C347 B.n307 VSUBS 0.007638f
C348 B.n308 VSUBS 0.007638f
C349 B.n309 VSUBS 0.007638f
C350 B.n310 VSUBS 0.007638f
C351 B.n311 VSUBS 0.007638f
C352 B.n312 VSUBS 0.007638f
C353 B.n313 VSUBS 0.007638f
C354 B.n314 VSUBS 0.007638f
C355 B.n315 VSUBS 0.007638f
C356 B.n316 VSUBS 0.007638f
C357 B.n317 VSUBS 0.007638f
C358 B.n318 VSUBS 0.007638f
C359 B.n319 VSUBS 0.007638f
C360 B.n320 VSUBS 0.007638f
C361 B.n321 VSUBS 0.007638f
C362 B.n322 VSUBS 0.007638f
C363 B.n323 VSUBS 0.007638f
C364 B.n324 VSUBS 0.007638f
C365 B.n325 VSUBS 0.007638f
C366 B.n326 VSUBS 0.007638f
C367 B.n327 VSUBS 0.007638f
C368 B.n328 VSUBS 0.007638f
C369 B.n329 VSUBS 0.007638f
C370 B.n330 VSUBS 0.007638f
C371 B.n331 VSUBS 0.007638f
C372 B.n332 VSUBS 0.007638f
C373 B.n333 VSUBS 0.007638f
C374 B.n334 VSUBS 0.007638f
C375 B.n335 VSUBS 0.007638f
C376 B.n336 VSUBS 0.007638f
C377 B.n337 VSUBS 0.007638f
C378 B.n338 VSUBS 0.007638f
C379 B.n339 VSUBS 0.007638f
C380 B.n340 VSUBS 0.007638f
C381 B.n341 VSUBS 0.007638f
C382 B.n342 VSUBS 0.007638f
C383 B.n343 VSUBS 0.007638f
C384 B.n344 VSUBS 0.007638f
C385 B.n345 VSUBS 0.007638f
C386 B.n346 VSUBS 0.007638f
C387 B.n347 VSUBS 0.007638f
C388 B.n348 VSUBS 0.007638f
C389 B.n349 VSUBS 0.007638f
C390 B.n350 VSUBS 0.007638f
C391 B.n351 VSUBS 0.007638f
C392 B.n352 VSUBS 0.007638f
C393 B.n353 VSUBS 0.007638f
C394 B.n354 VSUBS 0.007638f
C395 B.n355 VSUBS 0.007638f
C396 B.n356 VSUBS 0.007638f
C397 B.n357 VSUBS 0.007638f
C398 B.n358 VSUBS 0.007638f
C399 B.n359 VSUBS 0.007638f
C400 B.n360 VSUBS 0.007638f
C401 B.n361 VSUBS 0.007638f
C402 B.n362 VSUBS 0.007638f
C403 B.n363 VSUBS 0.007638f
C404 B.n364 VSUBS 0.007638f
C405 B.n365 VSUBS 0.007638f
C406 B.n366 VSUBS 0.007638f
C407 B.n367 VSUBS 0.007638f
C408 B.n368 VSUBS 0.007638f
C409 B.n369 VSUBS 0.007638f
C410 B.n370 VSUBS 0.007638f
C411 B.n371 VSUBS 0.007638f
C412 B.n372 VSUBS 0.007638f
C413 B.n373 VSUBS 0.007638f
C414 B.n374 VSUBS 0.007638f
C415 B.n375 VSUBS 0.007638f
C416 B.n376 VSUBS 0.007638f
C417 B.n377 VSUBS 0.007638f
C418 B.n378 VSUBS 0.007638f
C419 B.n379 VSUBS 0.007638f
C420 B.n380 VSUBS 0.007638f
C421 B.n381 VSUBS 0.007638f
C422 B.n382 VSUBS 0.019254f
C423 B.n383 VSUBS 0.018407f
C424 B.n384 VSUBS 0.018882f
C425 B.n385 VSUBS 0.007638f
C426 B.n386 VSUBS 0.007638f
C427 B.n387 VSUBS 0.007638f
C428 B.n388 VSUBS 0.007638f
C429 B.n389 VSUBS 0.007638f
C430 B.n390 VSUBS 0.007638f
C431 B.n391 VSUBS 0.007638f
C432 B.n392 VSUBS 0.007638f
C433 B.n393 VSUBS 0.007638f
C434 B.n394 VSUBS 0.007638f
C435 B.n395 VSUBS 0.007638f
C436 B.n396 VSUBS 0.007638f
C437 B.n397 VSUBS 0.007638f
C438 B.n398 VSUBS 0.007638f
C439 B.n399 VSUBS 0.007638f
C440 B.n400 VSUBS 0.007638f
C441 B.n401 VSUBS 0.007638f
C442 B.n402 VSUBS 0.007638f
C443 B.n403 VSUBS 0.007638f
C444 B.n404 VSUBS 0.007638f
C445 B.n405 VSUBS 0.007638f
C446 B.n406 VSUBS 0.007638f
C447 B.n407 VSUBS 0.007638f
C448 B.n408 VSUBS 0.007638f
C449 B.n409 VSUBS 0.007638f
C450 B.n410 VSUBS 0.007638f
C451 B.n411 VSUBS 0.007638f
C452 B.n412 VSUBS 0.007638f
C453 B.n413 VSUBS 0.007638f
C454 B.n414 VSUBS 0.007638f
C455 B.n415 VSUBS 0.007638f
C456 B.n416 VSUBS 0.007638f
C457 B.n417 VSUBS 0.007638f
C458 B.n418 VSUBS 0.007638f
C459 B.n419 VSUBS 0.007638f
C460 B.n420 VSUBS 0.007638f
C461 B.n421 VSUBS 0.007638f
C462 B.n422 VSUBS 0.007638f
C463 B.n423 VSUBS 0.007638f
C464 B.n424 VSUBS 0.007638f
C465 B.n425 VSUBS 0.007638f
C466 B.n426 VSUBS 0.007638f
C467 B.n427 VSUBS 0.007638f
C468 B.n428 VSUBS 0.007638f
C469 B.n429 VSUBS 0.007638f
C470 B.n430 VSUBS 0.007638f
C471 B.n431 VSUBS 0.007638f
C472 B.n432 VSUBS 0.007638f
C473 B.n433 VSUBS 0.007638f
C474 B.n434 VSUBS 0.007188f
C475 B.n435 VSUBS 0.017696f
C476 B.n436 VSUBS 0.004268f
C477 B.n437 VSUBS 0.007638f
C478 B.n438 VSUBS 0.007638f
C479 B.n439 VSUBS 0.007638f
C480 B.n440 VSUBS 0.007638f
C481 B.n441 VSUBS 0.007638f
C482 B.n442 VSUBS 0.007638f
C483 B.n443 VSUBS 0.007638f
C484 B.n444 VSUBS 0.007638f
C485 B.n445 VSUBS 0.007638f
C486 B.n446 VSUBS 0.007638f
C487 B.n447 VSUBS 0.007638f
C488 B.n448 VSUBS 0.007638f
C489 B.n449 VSUBS 0.004268f
C490 B.n450 VSUBS 0.007638f
C491 B.n451 VSUBS 0.007638f
C492 B.n452 VSUBS 0.007638f
C493 B.n453 VSUBS 0.007638f
C494 B.n454 VSUBS 0.007638f
C495 B.n455 VSUBS 0.007638f
C496 B.n456 VSUBS 0.007638f
C497 B.n457 VSUBS 0.007638f
C498 B.n458 VSUBS 0.007638f
C499 B.n459 VSUBS 0.007638f
C500 B.n460 VSUBS 0.007638f
C501 B.n461 VSUBS 0.007638f
C502 B.n462 VSUBS 0.007638f
C503 B.n463 VSUBS 0.007638f
C504 B.n464 VSUBS 0.007638f
C505 B.n465 VSUBS 0.007638f
C506 B.n466 VSUBS 0.007638f
C507 B.n467 VSUBS 0.007638f
C508 B.n468 VSUBS 0.007638f
C509 B.n469 VSUBS 0.007638f
C510 B.n470 VSUBS 0.007638f
C511 B.n471 VSUBS 0.007638f
C512 B.n472 VSUBS 0.007638f
C513 B.n473 VSUBS 0.007638f
C514 B.n474 VSUBS 0.007638f
C515 B.n475 VSUBS 0.007638f
C516 B.n476 VSUBS 0.007638f
C517 B.n477 VSUBS 0.007638f
C518 B.n478 VSUBS 0.007638f
C519 B.n479 VSUBS 0.007638f
C520 B.n480 VSUBS 0.007638f
C521 B.n481 VSUBS 0.007638f
C522 B.n482 VSUBS 0.007638f
C523 B.n483 VSUBS 0.007638f
C524 B.n484 VSUBS 0.007638f
C525 B.n485 VSUBS 0.007638f
C526 B.n486 VSUBS 0.007638f
C527 B.n487 VSUBS 0.007638f
C528 B.n488 VSUBS 0.007638f
C529 B.n489 VSUBS 0.007638f
C530 B.n490 VSUBS 0.007638f
C531 B.n491 VSUBS 0.007638f
C532 B.n492 VSUBS 0.007638f
C533 B.n493 VSUBS 0.007638f
C534 B.n494 VSUBS 0.007638f
C535 B.n495 VSUBS 0.007638f
C536 B.n496 VSUBS 0.007638f
C537 B.n497 VSUBS 0.007638f
C538 B.n498 VSUBS 0.007638f
C539 B.n499 VSUBS 0.007638f
C540 B.n500 VSUBS 0.018882f
C541 B.n501 VSUBS 0.018882f
C542 B.n502 VSUBS 0.018407f
C543 B.n503 VSUBS 0.007638f
C544 B.n504 VSUBS 0.007638f
C545 B.n505 VSUBS 0.007638f
C546 B.n506 VSUBS 0.007638f
C547 B.n507 VSUBS 0.007638f
C548 B.n508 VSUBS 0.007638f
C549 B.n509 VSUBS 0.007638f
C550 B.n510 VSUBS 0.007638f
C551 B.n511 VSUBS 0.007638f
C552 B.n512 VSUBS 0.007638f
C553 B.n513 VSUBS 0.007638f
C554 B.n514 VSUBS 0.007638f
C555 B.n515 VSUBS 0.007638f
C556 B.n516 VSUBS 0.007638f
C557 B.n517 VSUBS 0.007638f
C558 B.n518 VSUBS 0.007638f
C559 B.n519 VSUBS 0.007638f
C560 B.n520 VSUBS 0.007638f
C561 B.n521 VSUBS 0.007638f
C562 B.n522 VSUBS 0.007638f
C563 B.n523 VSUBS 0.007638f
C564 B.n524 VSUBS 0.007638f
C565 B.n525 VSUBS 0.007638f
C566 B.n526 VSUBS 0.007638f
C567 B.n527 VSUBS 0.007638f
C568 B.n528 VSUBS 0.007638f
C569 B.n529 VSUBS 0.007638f
C570 B.n530 VSUBS 0.007638f
C571 B.n531 VSUBS 0.007638f
C572 B.n532 VSUBS 0.007638f
C573 B.n533 VSUBS 0.007638f
C574 B.n534 VSUBS 0.007638f
C575 B.n535 VSUBS 0.007638f
C576 B.n536 VSUBS 0.007638f
C577 B.n537 VSUBS 0.007638f
C578 B.n538 VSUBS 0.007638f
C579 B.n539 VSUBS 0.007638f
C580 B.n540 VSUBS 0.007638f
C581 B.n541 VSUBS 0.007638f
C582 B.n542 VSUBS 0.007638f
C583 B.n543 VSUBS 0.017294f
C584 VDD1.t1 VSUBS 0.203688f
C585 VDD1.t3 VSUBS 0.203688f
C586 VDD1.n0 VSUBS 1.52246f
C587 VDD1.t0 VSUBS 0.203688f
C588 VDD1.t2 VSUBS 0.203688f
C589 VDD1.n1 VSUBS 2.11127f
C590 VP.n0 VSUBS 0.043643f
C591 VP.t1 VSUBS 2.04255f
C592 VP.n1 VSUBS 0.035316f
C593 VP.n2 VSUBS 0.043643f
C594 VP.t3 VSUBS 2.04255f
C595 VP.t2 VSUBS 2.25713f
C596 VP.t0 VSUBS 2.2546f
C597 VP.n3 VSUBS 3.29155f
C598 VP.n4 VSUBS 2.23031f
C599 VP.n5 VSUBS 0.845315f
C600 VP.n6 VSUBS 0.047036f
C601 VP.n7 VSUBS 0.087202f
C602 VP.n8 VSUBS 0.043643f
C603 VP.n9 VSUBS 0.043643f
C604 VP.n10 VSUBS 0.043643f
C605 VP.n11 VSUBS 0.087202f
C606 VP.n12 VSUBS 0.047036f
C607 VP.n13 VSUBS 0.845315f
C608 VP.n14 VSUBS 0.046736f
C609 VTAIL.t3 VSUBS 1.64893f
C610 VTAIL.n0 VSUBS 0.711786f
C611 VTAIL.t1 VSUBS 1.64893f
C612 VTAIL.n1 VSUBS 0.778632f
C613 VTAIL.t2 VSUBS 1.64893f
C614 VTAIL.n2 VSUBS 1.8485f
C615 VTAIL.t6 VSUBS 1.64894f
C616 VTAIL.n3 VSUBS 1.84849f
C617 VTAIL.t4 VSUBS 1.64894f
C618 VTAIL.n4 VSUBS 0.778619f
C619 VTAIL.t7 VSUBS 1.64894f
C620 VTAIL.n5 VSUBS 0.778619f
C621 VTAIL.t0 VSUBS 1.64893f
C622 VTAIL.n6 VSUBS 1.8485f
C623 VTAIL.t5 VSUBS 1.64893f
C624 VTAIL.n7 VSUBS 1.77266f
C625 VDD2.t2 VSUBS 0.203678f
C626 VDD2.t0 VSUBS 0.203678f
C627 VDD2.n0 VSUBS 2.08791f
C628 VDD2.t1 VSUBS 0.203678f
C629 VDD2.t3 VSUBS 0.203678f
C630 VDD2.n1 VSUBS 1.52189f
C631 VDD2.n2 VSUBS 3.80942f
C632 VN.t3 VSUBS 2.18016f
C633 VN.t1 VSUBS 2.17772f
C634 VN.n0 VSUBS 1.52465f
C635 VN.t2 VSUBS 2.18016f
C636 VN.t0 VSUBS 2.17772f
C637 VN.n1 VSUBS 3.20471f
.ends

