* NGSPICE file created from diff_pair_sample_1561.ext - technology: sky130A

.subckt diff_pair_sample_1561 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0.1452 ps=1.21 w=0.88 l=1.73
X1 VTAIL.t6 VN.t1 VDD2.t1 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0.1452 ps=1.21 w=0.88 l=1.73
X2 VDD1.t3 VP.t0 VTAIL.t3 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.1452 pd=1.21 as=0.3432 ps=2.54 w=0.88 l=1.73
X3 VDD2.t3 VN.t2 VTAIL.t5 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.1452 pd=1.21 as=0.3432 ps=2.54 w=0.88 l=1.73
X4 B.t11 B.t9 B.t10 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0 ps=0 w=0.88 l=1.73
X5 VTAIL.t0 VP.t1 VDD1.t2 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0.1452 ps=1.21 w=0.88 l=1.73
X6 VDD2.t2 VN.t3 VTAIL.t4 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.1452 pd=1.21 as=0.3432 ps=2.54 w=0.88 l=1.73
X7 VDD1.t1 VP.t2 VTAIL.t1 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.1452 pd=1.21 as=0.3432 ps=2.54 w=0.88 l=1.73
X8 VTAIL.t2 VP.t3 VDD1.t0 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0.1452 ps=1.21 w=0.88 l=1.73
X9 B.t8 B.t6 B.t7 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0 ps=0 w=0.88 l=1.73
X10 B.t5 B.t3 B.t4 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0 ps=0 w=0.88 l=1.73
X11 B.t2 B.t0 B.t1 w_n2206_n1144# sky130_fd_pr__pfet_01v8 ad=0.3432 pd=2.54 as=0 ps=0 w=0.88 l=1.73
R0 VN.n0 VN.t0 47.8259
R1 VN.n1 VN.t2 47.8259
R2 VN.n0 VN.t3 47.4011
R3 VN.n1 VN.t1 47.4011
R4 VN VN.n1 44.9273
R5 VN VN.n0 9.469
R6 VDD2.n2 VDD2.n0 667.606
R7 VDD2.n2 VDD2.n1 637.806
R8 VDD2.n1 VDD2.t1 36.938
R9 VDD2.n1 VDD2.t3 36.938
R10 VDD2.n0 VDD2.t0 36.938
R11 VDD2.n0 VDD2.t2 36.938
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n6 VTAIL.t3 658.064
R14 VTAIL.n5 VTAIL.t0 658.064
R15 VTAIL.n4 VTAIL.t5 658.064
R16 VTAIL.n3 VTAIL.t6 658.064
R17 VTAIL.n7 VTAIL.t4 658.063
R18 VTAIL.n0 VTAIL.t7 658.063
R19 VTAIL.n1 VTAIL.t1 658.063
R20 VTAIL.n2 VTAIL.t2 658.063
R21 VTAIL.n7 VTAIL.n6 14.9014
R22 VTAIL.n3 VTAIL.n2 14.9014
R23 VTAIL.n4 VTAIL.n3 1.77636
R24 VTAIL.n6 VTAIL.n5 1.77636
R25 VTAIL.n2 VTAIL.n1 1.77636
R26 VTAIL VTAIL.n0 0.946621
R27 VTAIL VTAIL.n7 0.830241
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 VP.n5 VP.n4 184.417
R31 VP.n14 VP.n13 184.417
R32 VP.n12 VP.n0 161.3
R33 VP.n11 VP.n10 161.3
R34 VP.n9 VP.n1 161.3
R35 VP.n8 VP.n7 161.3
R36 VP.n6 VP.n2 161.3
R37 VP.n3 VP.t1 47.8259
R38 VP.n3 VP.t0 47.4011
R39 VP.n4 VP.n3 44.5467
R40 VP.n7 VP.n1 40.577
R41 VP.n11 VP.n1 40.577
R42 VP.n7 VP.n6 24.5923
R43 VP.n12 VP.n11 24.5923
R44 VP.n5 VP.t3 12.2595
R45 VP.n13 VP.t2 12.2595
R46 VP.n6 VP.n5 1.47601
R47 VP.n13 VP.n12 1.47601
R48 VP.n4 VP.n2 0.189894
R49 VP.n8 VP.n2 0.189894
R50 VP.n9 VP.n8 0.189894
R51 VP.n10 VP.n9 0.189894
R52 VP.n10 VP.n0 0.189894
R53 VP.n14 VP.n0 0.189894
R54 VP VP.n14 0.0516364
R55 VDD1 VDD1.n1 668.13
R56 VDD1 VDD1.n0 637.864
R57 VDD1.n0 VDD1.t2 36.938
R58 VDD1.n0 VDD1.t3 36.938
R59 VDD1.n1 VDD1.t0 36.938
R60 VDD1.n1 VDD1.t1 36.938
R61 B.n64 B.t11 688.654
R62 B.n72 B.t8 688.654
R63 B.n20 B.t4 688.654
R64 B.n26 B.t1 688.654
R65 B.n65 B.t10 648.702
R66 B.n73 B.t7 648.702
R67 B.n21 B.t5 648.702
R68 B.n27 B.t2 648.702
R69 B.n250 B.n249 585
R70 B.n251 B.n32 585
R71 B.n253 B.n252 585
R72 B.n254 B.n31 585
R73 B.n256 B.n255 585
R74 B.n257 B.n30 585
R75 B.n259 B.n258 585
R76 B.n260 B.n29 585
R77 B.n262 B.n261 585
R78 B.n264 B.n263 585
R79 B.n265 B.n25 585
R80 B.n267 B.n266 585
R81 B.n268 B.n24 585
R82 B.n270 B.n269 585
R83 B.n271 B.n23 585
R84 B.n273 B.n272 585
R85 B.n274 B.n22 585
R86 B.n276 B.n275 585
R87 B.n278 B.n19 585
R88 B.n280 B.n279 585
R89 B.n281 B.n18 585
R90 B.n283 B.n282 585
R91 B.n284 B.n17 585
R92 B.n286 B.n285 585
R93 B.n287 B.n16 585
R94 B.n289 B.n288 585
R95 B.n290 B.n15 585
R96 B.n248 B.n33 585
R97 B.n247 B.n246 585
R98 B.n245 B.n34 585
R99 B.n244 B.n243 585
R100 B.n242 B.n35 585
R101 B.n241 B.n240 585
R102 B.n239 B.n36 585
R103 B.n238 B.n237 585
R104 B.n236 B.n37 585
R105 B.n235 B.n234 585
R106 B.n233 B.n38 585
R107 B.n232 B.n231 585
R108 B.n230 B.n39 585
R109 B.n229 B.n228 585
R110 B.n227 B.n40 585
R111 B.n226 B.n225 585
R112 B.n224 B.n41 585
R113 B.n223 B.n222 585
R114 B.n221 B.n42 585
R115 B.n220 B.n219 585
R116 B.n218 B.n43 585
R117 B.n217 B.n216 585
R118 B.n215 B.n44 585
R119 B.n214 B.n213 585
R120 B.n212 B.n45 585
R121 B.n211 B.n210 585
R122 B.n209 B.n46 585
R123 B.n208 B.n207 585
R124 B.n206 B.n47 585
R125 B.n205 B.n204 585
R126 B.n203 B.n48 585
R127 B.n202 B.n201 585
R128 B.n200 B.n49 585
R129 B.n199 B.n198 585
R130 B.n197 B.n50 585
R131 B.n196 B.n195 585
R132 B.n194 B.n51 585
R133 B.n193 B.n192 585
R134 B.n191 B.n52 585
R135 B.n190 B.n189 585
R136 B.n188 B.n53 585
R137 B.n187 B.n186 585
R138 B.n185 B.n54 585
R139 B.n184 B.n183 585
R140 B.n182 B.n55 585
R141 B.n181 B.n180 585
R142 B.n179 B.n56 585
R143 B.n178 B.n177 585
R144 B.n176 B.n57 585
R145 B.n175 B.n174 585
R146 B.n173 B.n58 585
R147 B.n172 B.n171 585
R148 B.n170 B.n59 585
R149 B.n128 B.n77 585
R150 B.n130 B.n129 585
R151 B.n131 B.n76 585
R152 B.n133 B.n132 585
R153 B.n134 B.n75 585
R154 B.n136 B.n135 585
R155 B.n137 B.n74 585
R156 B.n139 B.n138 585
R157 B.n140 B.n71 585
R158 B.n143 B.n142 585
R159 B.n144 B.n70 585
R160 B.n146 B.n145 585
R161 B.n147 B.n69 585
R162 B.n149 B.n148 585
R163 B.n150 B.n68 585
R164 B.n152 B.n151 585
R165 B.n153 B.n67 585
R166 B.n155 B.n154 585
R167 B.n157 B.n156 585
R168 B.n158 B.n63 585
R169 B.n160 B.n159 585
R170 B.n161 B.n62 585
R171 B.n163 B.n162 585
R172 B.n164 B.n61 585
R173 B.n166 B.n165 585
R174 B.n167 B.n60 585
R175 B.n169 B.n168 585
R176 B.n127 B.n126 585
R177 B.n125 B.n78 585
R178 B.n124 B.n123 585
R179 B.n122 B.n79 585
R180 B.n121 B.n120 585
R181 B.n119 B.n80 585
R182 B.n118 B.n117 585
R183 B.n116 B.n81 585
R184 B.n115 B.n114 585
R185 B.n113 B.n82 585
R186 B.n112 B.n111 585
R187 B.n110 B.n83 585
R188 B.n109 B.n108 585
R189 B.n107 B.n84 585
R190 B.n106 B.n105 585
R191 B.n104 B.n85 585
R192 B.n103 B.n102 585
R193 B.n101 B.n86 585
R194 B.n100 B.n99 585
R195 B.n98 B.n87 585
R196 B.n97 B.n96 585
R197 B.n95 B.n88 585
R198 B.n94 B.n93 585
R199 B.n92 B.n89 585
R200 B.n91 B.n90 585
R201 B.n2 B.n0 585
R202 B.n329 B.n1 585
R203 B.n328 B.n327 585
R204 B.n326 B.n3 585
R205 B.n325 B.n324 585
R206 B.n323 B.n4 585
R207 B.n322 B.n321 585
R208 B.n320 B.n5 585
R209 B.n319 B.n318 585
R210 B.n317 B.n6 585
R211 B.n316 B.n315 585
R212 B.n314 B.n7 585
R213 B.n313 B.n312 585
R214 B.n311 B.n8 585
R215 B.n310 B.n309 585
R216 B.n308 B.n9 585
R217 B.n307 B.n306 585
R218 B.n305 B.n10 585
R219 B.n304 B.n303 585
R220 B.n302 B.n11 585
R221 B.n301 B.n300 585
R222 B.n299 B.n12 585
R223 B.n298 B.n297 585
R224 B.n296 B.n13 585
R225 B.n295 B.n294 585
R226 B.n293 B.n14 585
R227 B.n292 B.n291 585
R228 B.n331 B.n330 585
R229 B.n126 B.n77 578.989
R230 B.n292 B.n15 578.989
R231 B.n168 B.n59 578.989
R232 B.n250 B.n33 578.989
R233 B.n64 B.t9 207.572
R234 B.n72 B.t6 207.572
R235 B.n20 B.t3 207.572
R236 B.n26 B.t0 207.572
R237 B.n126 B.n125 163.367
R238 B.n125 B.n124 163.367
R239 B.n124 B.n79 163.367
R240 B.n120 B.n79 163.367
R241 B.n120 B.n119 163.367
R242 B.n119 B.n118 163.367
R243 B.n118 B.n81 163.367
R244 B.n114 B.n81 163.367
R245 B.n114 B.n113 163.367
R246 B.n113 B.n112 163.367
R247 B.n112 B.n83 163.367
R248 B.n108 B.n83 163.367
R249 B.n108 B.n107 163.367
R250 B.n107 B.n106 163.367
R251 B.n106 B.n85 163.367
R252 B.n102 B.n85 163.367
R253 B.n102 B.n101 163.367
R254 B.n101 B.n100 163.367
R255 B.n100 B.n87 163.367
R256 B.n96 B.n87 163.367
R257 B.n96 B.n95 163.367
R258 B.n95 B.n94 163.367
R259 B.n94 B.n89 163.367
R260 B.n90 B.n89 163.367
R261 B.n90 B.n2 163.367
R262 B.n330 B.n2 163.367
R263 B.n330 B.n329 163.367
R264 B.n329 B.n328 163.367
R265 B.n328 B.n3 163.367
R266 B.n324 B.n3 163.367
R267 B.n324 B.n323 163.367
R268 B.n323 B.n322 163.367
R269 B.n322 B.n5 163.367
R270 B.n318 B.n5 163.367
R271 B.n318 B.n317 163.367
R272 B.n317 B.n316 163.367
R273 B.n316 B.n7 163.367
R274 B.n312 B.n7 163.367
R275 B.n312 B.n311 163.367
R276 B.n311 B.n310 163.367
R277 B.n310 B.n9 163.367
R278 B.n306 B.n9 163.367
R279 B.n306 B.n305 163.367
R280 B.n305 B.n304 163.367
R281 B.n304 B.n11 163.367
R282 B.n300 B.n11 163.367
R283 B.n300 B.n299 163.367
R284 B.n299 B.n298 163.367
R285 B.n298 B.n13 163.367
R286 B.n294 B.n13 163.367
R287 B.n294 B.n293 163.367
R288 B.n293 B.n292 163.367
R289 B.n130 B.n77 163.367
R290 B.n131 B.n130 163.367
R291 B.n132 B.n131 163.367
R292 B.n132 B.n75 163.367
R293 B.n136 B.n75 163.367
R294 B.n137 B.n136 163.367
R295 B.n138 B.n137 163.367
R296 B.n138 B.n71 163.367
R297 B.n143 B.n71 163.367
R298 B.n144 B.n143 163.367
R299 B.n145 B.n144 163.367
R300 B.n145 B.n69 163.367
R301 B.n149 B.n69 163.367
R302 B.n150 B.n149 163.367
R303 B.n151 B.n150 163.367
R304 B.n151 B.n67 163.367
R305 B.n155 B.n67 163.367
R306 B.n156 B.n155 163.367
R307 B.n156 B.n63 163.367
R308 B.n160 B.n63 163.367
R309 B.n161 B.n160 163.367
R310 B.n162 B.n161 163.367
R311 B.n162 B.n61 163.367
R312 B.n166 B.n61 163.367
R313 B.n167 B.n166 163.367
R314 B.n168 B.n167 163.367
R315 B.n172 B.n59 163.367
R316 B.n173 B.n172 163.367
R317 B.n174 B.n173 163.367
R318 B.n174 B.n57 163.367
R319 B.n178 B.n57 163.367
R320 B.n179 B.n178 163.367
R321 B.n180 B.n179 163.367
R322 B.n180 B.n55 163.367
R323 B.n184 B.n55 163.367
R324 B.n185 B.n184 163.367
R325 B.n186 B.n185 163.367
R326 B.n186 B.n53 163.367
R327 B.n190 B.n53 163.367
R328 B.n191 B.n190 163.367
R329 B.n192 B.n191 163.367
R330 B.n192 B.n51 163.367
R331 B.n196 B.n51 163.367
R332 B.n197 B.n196 163.367
R333 B.n198 B.n197 163.367
R334 B.n198 B.n49 163.367
R335 B.n202 B.n49 163.367
R336 B.n203 B.n202 163.367
R337 B.n204 B.n203 163.367
R338 B.n204 B.n47 163.367
R339 B.n208 B.n47 163.367
R340 B.n209 B.n208 163.367
R341 B.n210 B.n209 163.367
R342 B.n210 B.n45 163.367
R343 B.n214 B.n45 163.367
R344 B.n215 B.n214 163.367
R345 B.n216 B.n215 163.367
R346 B.n216 B.n43 163.367
R347 B.n220 B.n43 163.367
R348 B.n221 B.n220 163.367
R349 B.n222 B.n221 163.367
R350 B.n222 B.n41 163.367
R351 B.n226 B.n41 163.367
R352 B.n227 B.n226 163.367
R353 B.n228 B.n227 163.367
R354 B.n228 B.n39 163.367
R355 B.n232 B.n39 163.367
R356 B.n233 B.n232 163.367
R357 B.n234 B.n233 163.367
R358 B.n234 B.n37 163.367
R359 B.n238 B.n37 163.367
R360 B.n239 B.n238 163.367
R361 B.n240 B.n239 163.367
R362 B.n240 B.n35 163.367
R363 B.n244 B.n35 163.367
R364 B.n245 B.n244 163.367
R365 B.n246 B.n245 163.367
R366 B.n246 B.n33 163.367
R367 B.n288 B.n15 163.367
R368 B.n288 B.n287 163.367
R369 B.n287 B.n286 163.367
R370 B.n286 B.n17 163.367
R371 B.n282 B.n17 163.367
R372 B.n282 B.n281 163.367
R373 B.n281 B.n280 163.367
R374 B.n280 B.n19 163.367
R375 B.n275 B.n19 163.367
R376 B.n275 B.n274 163.367
R377 B.n274 B.n273 163.367
R378 B.n273 B.n23 163.367
R379 B.n269 B.n23 163.367
R380 B.n269 B.n268 163.367
R381 B.n268 B.n267 163.367
R382 B.n267 B.n25 163.367
R383 B.n263 B.n25 163.367
R384 B.n263 B.n262 163.367
R385 B.n262 B.n29 163.367
R386 B.n258 B.n29 163.367
R387 B.n258 B.n257 163.367
R388 B.n257 B.n256 163.367
R389 B.n256 B.n31 163.367
R390 B.n252 B.n31 163.367
R391 B.n252 B.n251 163.367
R392 B.n251 B.n250 163.367
R393 B.n66 B.n65 59.5399
R394 B.n141 B.n73 59.5399
R395 B.n277 B.n21 59.5399
R396 B.n28 B.n27 59.5399
R397 B.n65 B.n64 39.952
R398 B.n73 B.n72 39.952
R399 B.n21 B.n20 39.952
R400 B.n27 B.n26 39.952
R401 B.n291 B.n290 37.62
R402 B.n249 B.n248 37.62
R403 B.n170 B.n169 37.62
R404 B.n128 B.n127 37.62
R405 B B.n331 18.0485
R406 B.n290 B.n289 10.6151
R407 B.n289 B.n16 10.6151
R408 B.n285 B.n16 10.6151
R409 B.n285 B.n284 10.6151
R410 B.n284 B.n283 10.6151
R411 B.n283 B.n18 10.6151
R412 B.n279 B.n18 10.6151
R413 B.n279 B.n278 10.6151
R414 B.n276 B.n22 10.6151
R415 B.n272 B.n22 10.6151
R416 B.n272 B.n271 10.6151
R417 B.n271 B.n270 10.6151
R418 B.n270 B.n24 10.6151
R419 B.n266 B.n24 10.6151
R420 B.n266 B.n265 10.6151
R421 B.n265 B.n264 10.6151
R422 B.n261 B.n260 10.6151
R423 B.n260 B.n259 10.6151
R424 B.n259 B.n30 10.6151
R425 B.n255 B.n30 10.6151
R426 B.n255 B.n254 10.6151
R427 B.n254 B.n253 10.6151
R428 B.n253 B.n32 10.6151
R429 B.n249 B.n32 10.6151
R430 B.n171 B.n170 10.6151
R431 B.n171 B.n58 10.6151
R432 B.n175 B.n58 10.6151
R433 B.n176 B.n175 10.6151
R434 B.n177 B.n176 10.6151
R435 B.n177 B.n56 10.6151
R436 B.n181 B.n56 10.6151
R437 B.n182 B.n181 10.6151
R438 B.n183 B.n182 10.6151
R439 B.n183 B.n54 10.6151
R440 B.n187 B.n54 10.6151
R441 B.n188 B.n187 10.6151
R442 B.n189 B.n188 10.6151
R443 B.n189 B.n52 10.6151
R444 B.n193 B.n52 10.6151
R445 B.n194 B.n193 10.6151
R446 B.n195 B.n194 10.6151
R447 B.n195 B.n50 10.6151
R448 B.n199 B.n50 10.6151
R449 B.n200 B.n199 10.6151
R450 B.n201 B.n200 10.6151
R451 B.n201 B.n48 10.6151
R452 B.n205 B.n48 10.6151
R453 B.n206 B.n205 10.6151
R454 B.n207 B.n206 10.6151
R455 B.n207 B.n46 10.6151
R456 B.n211 B.n46 10.6151
R457 B.n212 B.n211 10.6151
R458 B.n213 B.n212 10.6151
R459 B.n213 B.n44 10.6151
R460 B.n217 B.n44 10.6151
R461 B.n218 B.n217 10.6151
R462 B.n219 B.n218 10.6151
R463 B.n219 B.n42 10.6151
R464 B.n223 B.n42 10.6151
R465 B.n224 B.n223 10.6151
R466 B.n225 B.n224 10.6151
R467 B.n225 B.n40 10.6151
R468 B.n229 B.n40 10.6151
R469 B.n230 B.n229 10.6151
R470 B.n231 B.n230 10.6151
R471 B.n231 B.n38 10.6151
R472 B.n235 B.n38 10.6151
R473 B.n236 B.n235 10.6151
R474 B.n237 B.n236 10.6151
R475 B.n237 B.n36 10.6151
R476 B.n241 B.n36 10.6151
R477 B.n242 B.n241 10.6151
R478 B.n243 B.n242 10.6151
R479 B.n243 B.n34 10.6151
R480 B.n247 B.n34 10.6151
R481 B.n248 B.n247 10.6151
R482 B.n129 B.n128 10.6151
R483 B.n129 B.n76 10.6151
R484 B.n133 B.n76 10.6151
R485 B.n134 B.n133 10.6151
R486 B.n135 B.n134 10.6151
R487 B.n135 B.n74 10.6151
R488 B.n139 B.n74 10.6151
R489 B.n140 B.n139 10.6151
R490 B.n142 B.n70 10.6151
R491 B.n146 B.n70 10.6151
R492 B.n147 B.n146 10.6151
R493 B.n148 B.n147 10.6151
R494 B.n148 B.n68 10.6151
R495 B.n152 B.n68 10.6151
R496 B.n153 B.n152 10.6151
R497 B.n154 B.n153 10.6151
R498 B.n158 B.n157 10.6151
R499 B.n159 B.n158 10.6151
R500 B.n159 B.n62 10.6151
R501 B.n163 B.n62 10.6151
R502 B.n164 B.n163 10.6151
R503 B.n165 B.n164 10.6151
R504 B.n165 B.n60 10.6151
R505 B.n169 B.n60 10.6151
R506 B.n127 B.n78 10.6151
R507 B.n123 B.n78 10.6151
R508 B.n123 B.n122 10.6151
R509 B.n122 B.n121 10.6151
R510 B.n121 B.n80 10.6151
R511 B.n117 B.n80 10.6151
R512 B.n117 B.n116 10.6151
R513 B.n116 B.n115 10.6151
R514 B.n115 B.n82 10.6151
R515 B.n111 B.n82 10.6151
R516 B.n111 B.n110 10.6151
R517 B.n110 B.n109 10.6151
R518 B.n109 B.n84 10.6151
R519 B.n105 B.n84 10.6151
R520 B.n105 B.n104 10.6151
R521 B.n104 B.n103 10.6151
R522 B.n103 B.n86 10.6151
R523 B.n99 B.n86 10.6151
R524 B.n99 B.n98 10.6151
R525 B.n98 B.n97 10.6151
R526 B.n97 B.n88 10.6151
R527 B.n93 B.n88 10.6151
R528 B.n93 B.n92 10.6151
R529 B.n92 B.n91 10.6151
R530 B.n91 B.n0 10.6151
R531 B.n327 B.n1 10.6151
R532 B.n327 B.n326 10.6151
R533 B.n326 B.n325 10.6151
R534 B.n325 B.n4 10.6151
R535 B.n321 B.n4 10.6151
R536 B.n321 B.n320 10.6151
R537 B.n320 B.n319 10.6151
R538 B.n319 B.n6 10.6151
R539 B.n315 B.n6 10.6151
R540 B.n315 B.n314 10.6151
R541 B.n314 B.n313 10.6151
R542 B.n313 B.n8 10.6151
R543 B.n309 B.n8 10.6151
R544 B.n309 B.n308 10.6151
R545 B.n308 B.n307 10.6151
R546 B.n307 B.n10 10.6151
R547 B.n303 B.n10 10.6151
R548 B.n303 B.n302 10.6151
R549 B.n302 B.n301 10.6151
R550 B.n301 B.n12 10.6151
R551 B.n297 B.n12 10.6151
R552 B.n297 B.n296 10.6151
R553 B.n296 B.n295 10.6151
R554 B.n295 B.n14 10.6151
R555 B.n291 B.n14 10.6151
R556 B.n277 B.n276 6.5566
R557 B.n264 B.n28 6.5566
R558 B.n142 B.n141 6.5566
R559 B.n154 B.n66 6.5566
R560 B.n278 B.n277 4.05904
R561 B.n261 B.n28 4.05904
R562 B.n141 B.n140 4.05904
R563 B.n157 B.n66 4.05904
R564 B.n331 B.n0 2.81026
R565 B.n331 B.n1 2.81026
C0 VDD2 VP 0.347647f
C1 VDD1 VN 0.155579f
C2 VP B 1.22812f
C3 VN w_n2206_n1144# 3.33092f
C4 VDD1 VTAIL 2.29748f
C5 VDD2 VN 0.616002f
C6 VTAIL w_n2206_n1144# 1.30094f
C7 VN B 0.766544f
C8 VDD2 VTAIL 2.34585f
C9 VDD1 w_n2206_n1144# 0.971946f
C10 VTAIL B 0.960894f
C11 VN VP 3.51245f
C12 VDD2 VDD1 0.814886f
C13 VTAIL VP 1.10906f
C14 VDD1 B 0.80823f
C15 VDD2 w_n2206_n1144# 1.00746f
C16 B w_n2206_n1144# 5.08476f
C17 VDD1 VP 0.80609f
C18 VDD2 B 0.846674f
C19 VTAIL VN 1.09495f
C20 VP w_n2206_n1144# 3.60414f
C21 VDD2 VSUBS 0.513493f
C22 VDD1 VSUBS 2.812527f
C23 VTAIL VSUBS 0.332783f
C24 VN VSUBS 4.78955f
C25 VP VSUBS 1.268571f
C26 B VSUBS 2.444165f
C27 w_n2206_n1144# VSUBS 32.587f
C28 B.n0 VSUBS 0.006855f
C29 B.n1 VSUBS 0.006855f
C30 B.n2 VSUBS 0.01084f
C31 B.n3 VSUBS 0.01084f
C32 B.n4 VSUBS 0.01084f
C33 B.n5 VSUBS 0.01084f
C34 B.n6 VSUBS 0.01084f
C35 B.n7 VSUBS 0.01084f
C36 B.n8 VSUBS 0.01084f
C37 B.n9 VSUBS 0.01084f
C38 B.n10 VSUBS 0.01084f
C39 B.n11 VSUBS 0.01084f
C40 B.n12 VSUBS 0.01084f
C41 B.n13 VSUBS 0.01084f
C42 B.n14 VSUBS 0.01084f
C43 B.n15 VSUBS 0.028507f
C44 B.n16 VSUBS 0.01084f
C45 B.n17 VSUBS 0.01084f
C46 B.n18 VSUBS 0.01084f
C47 B.n19 VSUBS 0.01084f
C48 B.t5 VSUBS 0.026321f
C49 B.t4 VSUBS 0.029037f
C50 B.t3 VSUBS 0.122008f
C51 B.n20 VSUBS 0.075375f
C52 B.n21 VSUBS 0.062275f
C53 B.n22 VSUBS 0.01084f
C54 B.n23 VSUBS 0.01084f
C55 B.n24 VSUBS 0.01084f
C56 B.n25 VSUBS 0.01084f
C57 B.t2 VSUBS 0.026321f
C58 B.t1 VSUBS 0.029037f
C59 B.t0 VSUBS 0.122008f
C60 B.n26 VSUBS 0.075375f
C61 B.n27 VSUBS 0.062275f
C62 B.n28 VSUBS 0.025115f
C63 B.n29 VSUBS 0.01084f
C64 B.n30 VSUBS 0.01084f
C65 B.n31 VSUBS 0.01084f
C66 B.n32 VSUBS 0.01084f
C67 B.n33 VSUBS 0.027287f
C68 B.n34 VSUBS 0.01084f
C69 B.n35 VSUBS 0.01084f
C70 B.n36 VSUBS 0.01084f
C71 B.n37 VSUBS 0.01084f
C72 B.n38 VSUBS 0.01084f
C73 B.n39 VSUBS 0.01084f
C74 B.n40 VSUBS 0.01084f
C75 B.n41 VSUBS 0.01084f
C76 B.n42 VSUBS 0.01084f
C77 B.n43 VSUBS 0.01084f
C78 B.n44 VSUBS 0.01084f
C79 B.n45 VSUBS 0.01084f
C80 B.n46 VSUBS 0.01084f
C81 B.n47 VSUBS 0.01084f
C82 B.n48 VSUBS 0.01084f
C83 B.n49 VSUBS 0.01084f
C84 B.n50 VSUBS 0.01084f
C85 B.n51 VSUBS 0.01084f
C86 B.n52 VSUBS 0.01084f
C87 B.n53 VSUBS 0.01084f
C88 B.n54 VSUBS 0.01084f
C89 B.n55 VSUBS 0.01084f
C90 B.n56 VSUBS 0.01084f
C91 B.n57 VSUBS 0.01084f
C92 B.n58 VSUBS 0.01084f
C93 B.n59 VSUBS 0.027287f
C94 B.n60 VSUBS 0.01084f
C95 B.n61 VSUBS 0.01084f
C96 B.n62 VSUBS 0.01084f
C97 B.n63 VSUBS 0.01084f
C98 B.t10 VSUBS 0.026321f
C99 B.t11 VSUBS 0.029037f
C100 B.t9 VSUBS 0.122008f
C101 B.n64 VSUBS 0.075375f
C102 B.n65 VSUBS 0.062275f
C103 B.n66 VSUBS 0.025115f
C104 B.n67 VSUBS 0.01084f
C105 B.n68 VSUBS 0.01084f
C106 B.n69 VSUBS 0.01084f
C107 B.n70 VSUBS 0.01084f
C108 B.n71 VSUBS 0.01084f
C109 B.t7 VSUBS 0.026321f
C110 B.t8 VSUBS 0.029037f
C111 B.t6 VSUBS 0.122008f
C112 B.n72 VSUBS 0.075375f
C113 B.n73 VSUBS 0.062275f
C114 B.n74 VSUBS 0.01084f
C115 B.n75 VSUBS 0.01084f
C116 B.n76 VSUBS 0.01084f
C117 B.n77 VSUBS 0.028507f
C118 B.n78 VSUBS 0.01084f
C119 B.n79 VSUBS 0.01084f
C120 B.n80 VSUBS 0.01084f
C121 B.n81 VSUBS 0.01084f
C122 B.n82 VSUBS 0.01084f
C123 B.n83 VSUBS 0.01084f
C124 B.n84 VSUBS 0.01084f
C125 B.n85 VSUBS 0.01084f
C126 B.n86 VSUBS 0.01084f
C127 B.n87 VSUBS 0.01084f
C128 B.n88 VSUBS 0.01084f
C129 B.n89 VSUBS 0.01084f
C130 B.n90 VSUBS 0.01084f
C131 B.n91 VSUBS 0.01084f
C132 B.n92 VSUBS 0.01084f
C133 B.n93 VSUBS 0.01084f
C134 B.n94 VSUBS 0.01084f
C135 B.n95 VSUBS 0.01084f
C136 B.n96 VSUBS 0.01084f
C137 B.n97 VSUBS 0.01084f
C138 B.n98 VSUBS 0.01084f
C139 B.n99 VSUBS 0.01084f
C140 B.n100 VSUBS 0.01084f
C141 B.n101 VSUBS 0.01084f
C142 B.n102 VSUBS 0.01084f
C143 B.n103 VSUBS 0.01084f
C144 B.n104 VSUBS 0.01084f
C145 B.n105 VSUBS 0.01084f
C146 B.n106 VSUBS 0.01084f
C147 B.n107 VSUBS 0.01084f
C148 B.n108 VSUBS 0.01084f
C149 B.n109 VSUBS 0.01084f
C150 B.n110 VSUBS 0.01084f
C151 B.n111 VSUBS 0.01084f
C152 B.n112 VSUBS 0.01084f
C153 B.n113 VSUBS 0.01084f
C154 B.n114 VSUBS 0.01084f
C155 B.n115 VSUBS 0.01084f
C156 B.n116 VSUBS 0.01084f
C157 B.n117 VSUBS 0.01084f
C158 B.n118 VSUBS 0.01084f
C159 B.n119 VSUBS 0.01084f
C160 B.n120 VSUBS 0.01084f
C161 B.n121 VSUBS 0.01084f
C162 B.n122 VSUBS 0.01084f
C163 B.n123 VSUBS 0.01084f
C164 B.n124 VSUBS 0.01084f
C165 B.n125 VSUBS 0.01084f
C166 B.n126 VSUBS 0.027287f
C167 B.n127 VSUBS 0.027287f
C168 B.n128 VSUBS 0.028507f
C169 B.n129 VSUBS 0.01084f
C170 B.n130 VSUBS 0.01084f
C171 B.n131 VSUBS 0.01084f
C172 B.n132 VSUBS 0.01084f
C173 B.n133 VSUBS 0.01084f
C174 B.n134 VSUBS 0.01084f
C175 B.n135 VSUBS 0.01084f
C176 B.n136 VSUBS 0.01084f
C177 B.n137 VSUBS 0.01084f
C178 B.n138 VSUBS 0.01084f
C179 B.n139 VSUBS 0.01084f
C180 B.n140 VSUBS 0.007492f
C181 B.n141 VSUBS 0.025115f
C182 B.n142 VSUBS 0.008768f
C183 B.n143 VSUBS 0.01084f
C184 B.n144 VSUBS 0.01084f
C185 B.n145 VSUBS 0.01084f
C186 B.n146 VSUBS 0.01084f
C187 B.n147 VSUBS 0.01084f
C188 B.n148 VSUBS 0.01084f
C189 B.n149 VSUBS 0.01084f
C190 B.n150 VSUBS 0.01084f
C191 B.n151 VSUBS 0.01084f
C192 B.n152 VSUBS 0.01084f
C193 B.n153 VSUBS 0.01084f
C194 B.n154 VSUBS 0.008768f
C195 B.n155 VSUBS 0.01084f
C196 B.n156 VSUBS 0.01084f
C197 B.n157 VSUBS 0.007492f
C198 B.n158 VSUBS 0.01084f
C199 B.n159 VSUBS 0.01084f
C200 B.n160 VSUBS 0.01084f
C201 B.n161 VSUBS 0.01084f
C202 B.n162 VSUBS 0.01084f
C203 B.n163 VSUBS 0.01084f
C204 B.n164 VSUBS 0.01084f
C205 B.n165 VSUBS 0.01084f
C206 B.n166 VSUBS 0.01084f
C207 B.n167 VSUBS 0.01084f
C208 B.n168 VSUBS 0.028507f
C209 B.n169 VSUBS 0.028507f
C210 B.n170 VSUBS 0.027287f
C211 B.n171 VSUBS 0.01084f
C212 B.n172 VSUBS 0.01084f
C213 B.n173 VSUBS 0.01084f
C214 B.n174 VSUBS 0.01084f
C215 B.n175 VSUBS 0.01084f
C216 B.n176 VSUBS 0.01084f
C217 B.n177 VSUBS 0.01084f
C218 B.n178 VSUBS 0.01084f
C219 B.n179 VSUBS 0.01084f
C220 B.n180 VSUBS 0.01084f
C221 B.n181 VSUBS 0.01084f
C222 B.n182 VSUBS 0.01084f
C223 B.n183 VSUBS 0.01084f
C224 B.n184 VSUBS 0.01084f
C225 B.n185 VSUBS 0.01084f
C226 B.n186 VSUBS 0.01084f
C227 B.n187 VSUBS 0.01084f
C228 B.n188 VSUBS 0.01084f
C229 B.n189 VSUBS 0.01084f
C230 B.n190 VSUBS 0.01084f
C231 B.n191 VSUBS 0.01084f
C232 B.n192 VSUBS 0.01084f
C233 B.n193 VSUBS 0.01084f
C234 B.n194 VSUBS 0.01084f
C235 B.n195 VSUBS 0.01084f
C236 B.n196 VSUBS 0.01084f
C237 B.n197 VSUBS 0.01084f
C238 B.n198 VSUBS 0.01084f
C239 B.n199 VSUBS 0.01084f
C240 B.n200 VSUBS 0.01084f
C241 B.n201 VSUBS 0.01084f
C242 B.n202 VSUBS 0.01084f
C243 B.n203 VSUBS 0.01084f
C244 B.n204 VSUBS 0.01084f
C245 B.n205 VSUBS 0.01084f
C246 B.n206 VSUBS 0.01084f
C247 B.n207 VSUBS 0.01084f
C248 B.n208 VSUBS 0.01084f
C249 B.n209 VSUBS 0.01084f
C250 B.n210 VSUBS 0.01084f
C251 B.n211 VSUBS 0.01084f
C252 B.n212 VSUBS 0.01084f
C253 B.n213 VSUBS 0.01084f
C254 B.n214 VSUBS 0.01084f
C255 B.n215 VSUBS 0.01084f
C256 B.n216 VSUBS 0.01084f
C257 B.n217 VSUBS 0.01084f
C258 B.n218 VSUBS 0.01084f
C259 B.n219 VSUBS 0.01084f
C260 B.n220 VSUBS 0.01084f
C261 B.n221 VSUBS 0.01084f
C262 B.n222 VSUBS 0.01084f
C263 B.n223 VSUBS 0.01084f
C264 B.n224 VSUBS 0.01084f
C265 B.n225 VSUBS 0.01084f
C266 B.n226 VSUBS 0.01084f
C267 B.n227 VSUBS 0.01084f
C268 B.n228 VSUBS 0.01084f
C269 B.n229 VSUBS 0.01084f
C270 B.n230 VSUBS 0.01084f
C271 B.n231 VSUBS 0.01084f
C272 B.n232 VSUBS 0.01084f
C273 B.n233 VSUBS 0.01084f
C274 B.n234 VSUBS 0.01084f
C275 B.n235 VSUBS 0.01084f
C276 B.n236 VSUBS 0.01084f
C277 B.n237 VSUBS 0.01084f
C278 B.n238 VSUBS 0.01084f
C279 B.n239 VSUBS 0.01084f
C280 B.n240 VSUBS 0.01084f
C281 B.n241 VSUBS 0.01084f
C282 B.n242 VSUBS 0.01084f
C283 B.n243 VSUBS 0.01084f
C284 B.n244 VSUBS 0.01084f
C285 B.n245 VSUBS 0.01084f
C286 B.n246 VSUBS 0.01084f
C287 B.n247 VSUBS 0.01084f
C288 B.n248 VSUBS 0.028399f
C289 B.n249 VSUBS 0.027395f
C290 B.n250 VSUBS 0.028507f
C291 B.n251 VSUBS 0.01084f
C292 B.n252 VSUBS 0.01084f
C293 B.n253 VSUBS 0.01084f
C294 B.n254 VSUBS 0.01084f
C295 B.n255 VSUBS 0.01084f
C296 B.n256 VSUBS 0.01084f
C297 B.n257 VSUBS 0.01084f
C298 B.n258 VSUBS 0.01084f
C299 B.n259 VSUBS 0.01084f
C300 B.n260 VSUBS 0.01084f
C301 B.n261 VSUBS 0.007492f
C302 B.n262 VSUBS 0.01084f
C303 B.n263 VSUBS 0.01084f
C304 B.n264 VSUBS 0.008768f
C305 B.n265 VSUBS 0.01084f
C306 B.n266 VSUBS 0.01084f
C307 B.n267 VSUBS 0.01084f
C308 B.n268 VSUBS 0.01084f
C309 B.n269 VSUBS 0.01084f
C310 B.n270 VSUBS 0.01084f
C311 B.n271 VSUBS 0.01084f
C312 B.n272 VSUBS 0.01084f
C313 B.n273 VSUBS 0.01084f
C314 B.n274 VSUBS 0.01084f
C315 B.n275 VSUBS 0.01084f
C316 B.n276 VSUBS 0.008768f
C317 B.n277 VSUBS 0.025115f
C318 B.n278 VSUBS 0.007492f
C319 B.n279 VSUBS 0.01084f
C320 B.n280 VSUBS 0.01084f
C321 B.n281 VSUBS 0.01084f
C322 B.n282 VSUBS 0.01084f
C323 B.n283 VSUBS 0.01084f
C324 B.n284 VSUBS 0.01084f
C325 B.n285 VSUBS 0.01084f
C326 B.n286 VSUBS 0.01084f
C327 B.n287 VSUBS 0.01084f
C328 B.n288 VSUBS 0.01084f
C329 B.n289 VSUBS 0.01084f
C330 B.n290 VSUBS 0.028507f
C331 B.n291 VSUBS 0.027287f
C332 B.n292 VSUBS 0.027287f
C333 B.n293 VSUBS 0.01084f
C334 B.n294 VSUBS 0.01084f
C335 B.n295 VSUBS 0.01084f
C336 B.n296 VSUBS 0.01084f
C337 B.n297 VSUBS 0.01084f
C338 B.n298 VSUBS 0.01084f
C339 B.n299 VSUBS 0.01084f
C340 B.n300 VSUBS 0.01084f
C341 B.n301 VSUBS 0.01084f
C342 B.n302 VSUBS 0.01084f
C343 B.n303 VSUBS 0.01084f
C344 B.n304 VSUBS 0.01084f
C345 B.n305 VSUBS 0.01084f
C346 B.n306 VSUBS 0.01084f
C347 B.n307 VSUBS 0.01084f
C348 B.n308 VSUBS 0.01084f
C349 B.n309 VSUBS 0.01084f
C350 B.n310 VSUBS 0.01084f
C351 B.n311 VSUBS 0.01084f
C352 B.n312 VSUBS 0.01084f
C353 B.n313 VSUBS 0.01084f
C354 B.n314 VSUBS 0.01084f
C355 B.n315 VSUBS 0.01084f
C356 B.n316 VSUBS 0.01084f
C357 B.n317 VSUBS 0.01084f
C358 B.n318 VSUBS 0.01084f
C359 B.n319 VSUBS 0.01084f
C360 B.n320 VSUBS 0.01084f
C361 B.n321 VSUBS 0.01084f
C362 B.n322 VSUBS 0.01084f
C363 B.n323 VSUBS 0.01084f
C364 B.n324 VSUBS 0.01084f
C365 B.n325 VSUBS 0.01084f
C366 B.n326 VSUBS 0.01084f
C367 B.n327 VSUBS 0.01084f
C368 B.n328 VSUBS 0.01084f
C369 B.n329 VSUBS 0.01084f
C370 B.n330 VSUBS 0.01084f
C371 B.n331 VSUBS 0.024546f
C372 VDD1.t2 VSUBS 0.014816f
C373 VDD1.t3 VSUBS 0.014816f
C374 VDD1.n0 VSUBS 0.040046f
C375 VDD1.t0 VSUBS 0.014816f
C376 VDD1.t1 VSUBS 0.014816f
C377 VDD1.n1 VSUBS 0.073722f
C378 VP.n0 VSUBS 0.061115f
C379 VP.t2 VSUBS 0.16198f
C380 VP.n1 VSUBS 0.049361f
C381 VP.n2 VSUBS 0.061115f
C382 VP.t3 VSUBS 0.16198f
C383 VP.t1 VSUBS 0.480652f
C384 VP.t0 VSUBS 0.477109f
C385 VP.n3 VSUBS 2.08835f
C386 VP.n4 VSUBS 2.38708f
C387 VP.n5 VSUBS 0.267439f
C388 VP.n6 VSUBS 0.06074f
C389 VP.n7 VSUBS 0.120827f
C390 VP.n8 VSUBS 0.061115f
C391 VP.n9 VSUBS 0.061115f
C392 VP.n10 VSUBS 0.061115f
C393 VP.n11 VSUBS 0.120827f
C394 VP.n12 VSUBS 0.06074f
C395 VP.n13 VSUBS 0.267439f
C396 VP.n14 VSUBS 0.065215f
C397 VTAIL.t7 VSUBS 0.07274f
C398 VTAIL.n0 VSUBS 0.230375f
C399 VTAIL.t1 VSUBS 0.07274f
C400 VTAIL.n1 VSUBS 0.287201f
C401 VTAIL.t2 VSUBS 0.07274f
C402 VTAIL.n2 VSUBS 0.717319f
C403 VTAIL.t6 VSUBS 0.07274f
C404 VTAIL.n3 VSUBS 0.717319f
C405 VTAIL.t5 VSUBS 0.07274f
C406 VTAIL.n4 VSUBS 0.287201f
C407 VTAIL.t0 VSUBS 0.07274f
C408 VTAIL.n5 VSUBS 0.287201f
C409 VTAIL.t3 VSUBS 0.07274f
C410 VTAIL.n6 VSUBS 0.717319f
C411 VTAIL.t4 VSUBS 0.07274f
C412 VTAIL.n7 VSUBS 0.652522f
C413 VDD2.t0 VSUBS 0.01534f
C414 VDD2.t2 VSUBS 0.01534f
C415 VDD2.n0 VSUBS 0.073739f
C416 VDD2.t1 VSUBS 0.01534f
C417 VDD2.t3 VSUBS 0.01534f
C418 VDD2.n1 VSUBS 0.041438f
C419 VDD2.n2 VSUBS 1.99248f
C420 VN.t0 VSUBS 0.454839f
C421 VN.t3 VSUBS 0.451487f
C422 VN.n0 VSUBS 0.310504f
C423 VN.t2 VSUBS 0.454839f
C424 VN.t1 VSUBS 0.451487f
C425 VN.n1 VSUBS 2.01036f
.ends

