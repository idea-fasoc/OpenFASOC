* NGSPICE file created from diff_pair_sample_1339.ext - technology: sky130A

.subckt diff_pair_sample_1339 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=4.8282 ps=25.54 w=12.38 l=3.92
X1 VDD1.t9 VP.t0 VTAIL.t5 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=2.0427 ps=12.71 w=12.38 l=3.92
X2 VDD1.t8 VP.t1 VTAIL.t7 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=4.8282 ps=25.54 w=12.38 l=3.92
X3 VDD1.t7 VP.t2 VTAIL.t0 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=2.0427 ps=12.71 w=12.38 l=3.92
X4 B.t11 B.t9 B.t10 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=0 ps=0 w=12.38 l=3.92
X5 VTAIL.t6 VP.t3 VDD1.t6 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X6 VDD2.t8 VN.t1 VTAIL.t13 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=4.8282 ps=25.54 w=12.38 l=3.92
X7 VDD2.t7 VN.t2 VTAIL.t14 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X8 VDD2.t6 VN.t3 VTAIL.t15 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=2.0427 ps=12.71 w=12.38 l=3.92
X9 VTAIL.t10 VN.t4 VDD2.t5 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X10 VTAIL.t18 VN.t5 VDD2.t4 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X11 VDD1.t5 VP.t4 VTAIL.t4 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=4.8282 ps=25.54 w=12.38 l=3.92
X12 VTAIL.t2 VP.t5 VDD1.t4 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X13 B.t8 B.t6 B.t7 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=0 ps=0 w=12.38 l=3.92
X14 VDD1.t3 VP.t6 VTAIL.t1 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X15 VTAIL.t17 VN.t6 VDD2.t3 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X16 B.t5 B.t3 B.t4 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=0 ps=0 w=12.38 l=3.92
X17 VTAIL.t12 VN.t7 VDD2.t2 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X18 VDD2.t1 VN.t8 VTAIL.t16 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X19 VTAIL.t9 VP.t7 VDD1.t2 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X20 VTAIL.t8 VP.t8 VDD1.t1 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
X21 VDD2.t0 VN.t9 VTAIL.t19 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=2.0427 ps=12.71 w=12.38 l=3.92
X22 B.t2 B.t0 B.t1 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=4.8282 pd=25.54 as=0 ps=0 w=12.38 l=3.92
X23 VDD1.t0 VP.t9 VTAIL.t3 w_n6070_n3444# sky130_fd_pr__pfet_01v8 ad=2.0427 pd=12.71 as=2.0427 ps=12.71 w=12.38 l=3.92
R0 VN.n107 VN.n55 161.3
R1 VN.n106 VN.n105 161.3
R2 VN.n104 VN.n56 161.3
R3 VN.n103 VN.n102 161.3
R4 VN.n101 VN.n57 161.3
R5 VN.n100 VN.n99 161.3
R6 VN.n98 VN.n58 161.3
R7 VN.n97 VN.n96 161.3
R8 VN.n94 VN.n59 161.3
R9 VN.n93 VN.n92 161.3
R10 VN.n91 VN.n60 161.3
R11 VN.n90 VN.n89 161.3
R12 VN.n88 VN.n61 161.3
R13 VN.n87 VN.n86 161.3
R14 VN.n85 VN.n62 161.3
R15 VN.n84 VN.n83 161.3
R16 VN.n82 VN.n63 161.3
R17 VN.n81 VN.n80 161.3
R18 VN.n79 VN.n64 161.3
R19 VN.n78 VN.n77 161.3
R20 VN.n76 VN.n65 161.3
R21 VN.n75 VN.n74 161.3
R22 VN.n73 VN.n66 161.3
R23 VN.n72 VN.n71 161.3
R24 VN.n70 VN.n67 161.3
R25 VN.n52 VN.n0 161.3
R26 VN.n51 VN.n50 161.3
R27 VN.n49 VN.n1 161.3
R28 VN.n48 VN.n47 161.3
R29 VN.n46 VN.n2 161.3
R30 VN.n45 VN.n44 161.3
R31 VN.n43 VN.n3 161.3
R32 VN.n42 VN.n41 161.3
R33 VN.n39 VN.n4 161.3
R34 VN.n38 VN.n37 161.3
R35 VN.n36 VN.n5 161.3
R36 VN.n35 VN.n34 161.3
R37 VN.n33 VN.n6 161.3
R38 VN.n32 VN.n31 161.3
R39 VN.n30 VN.n7 161.3
R40 VN.n29 VN.n28 161.3
R41 VN.n27 VN.n8 161.3
R42 VN.n26 VN.n25 161.3
R43 VN.n24 VN.n9 161.3
R44 VN.n23 VN.n22 161.3
R45 VN.n21 VN.n10 161.3
R46 VN.n20 VN.n19 161.3
R47 VN.n18 VN.n11 161.3
R48 VN.n17 VN.n16 161.3
R49 VN.n15 VN.n12 161.3
R50 VN.n13 VN.t3 108.032
R51 VN.n68 VN.t1 108.032
R52 VN.n53 VN.t0 76.1122
R53 VN.n27 VN.t8 76.1122
R54 VN.n14 VN.t5 76.1122
R55 VN.n40 VN.t6 76.1122
R56 VN.n108 VN.t9 76.1122
R57 VN.n82 VN.t2 76.1122
R58 VN.n69 VN.t7 76.1122
R59 VN.n95 VN.t4 76.1122
R60 VN.n14 VN.n13 62.7546
R61 VN.n69 VN.n68 62.7546
R62 VN VN.n109 60.9092
R63 VN.n54 VN.n53 57.6421
R64 VN.n109 VN.n108 57.6421
R65 VN.n21 VN.n20 52.5823
R66 VN.n34 VN.n33 52.5823
R67 VN.n47 VN.n46 52.5823
R68 VN.n76 VN.n75 52.5823
R69 VN.n89 VN.n88 52.5823
R70 VN.n102 VN.n101 52.5823
R71 VN.n22 VN.n21 28.2389
R72 VN.n33 VN.n32 28.2389
R73 VN.n47 VN.n1 28.2389
R74 VN.n77 VN.n76 28.2389
R75 VN.n88 VN.n87 28.2389
R76 VN.n102 VN.n56 28.2389
R77 VN.n16 VN.n15 24.3439
R78 VN.n16 VN.n11 24.3439
R79 VN.n20 VN.n11 24.3439
R80 VN.n22 VN.n9 24.3439
R81 VN.n26 VN.n9 24.3439
R82 VN.n27 VN.n26 24.3439
R83 VN.n28 VN.n27 24.3439
R84 VN.n28 VN.n7 24.3439
R85 VN.n32 VN.n7 24.3439
R86 VN.n34 VN.n5 24.3439
R87 VN.n38 VN.n5 24.3439
R88 VN.n39 VN.n38 24.3439
R89 VN.n41 VN.n3 24.3439
R90 VN.n45 VN.n3 24.3439
R91 VN.n46 VN.n45 24.3439
R92 VN.n51 VN.n1 24.3439
R93 VN.n52 VN.n51 24.3439
R94 VN.n53 VN.n52 24.3439
R95 VN.n75 VN.n66 24.3439
R96 VN.n71 VN.n66 24.3439
R97 VN.n71 VN.n70 24.3439
R98 VN.n87 VN.n62 24.3439
R99 VN.n83 VN.n62 24.3439
R100 VN.n83 VN.n82 24.3439
R101 VN.n82 VN.n81 24.3439
R102 VN.n81 VN.n64 24.3439
R103 VN.n77 VN.n64 24.3439
R104 VN.n101 VN.n100 24.3439
R105 VN.n100 VN.n58 24.3439
R106 VN.n96 VN.n58 24.3439
R107 VN.n94 VN.n93 24.3439
R108 VN.n93 VN.n60 24.3439
R109 VN.n89 VN.n60 24.3439
R110 VN.n108 VN.n107 24.3439
R111 VN.n107 VN.n106 24.3439
R112 VN.n106 VN.n56 24.3439
R113 VN.n15 VN.n14 12.1722
R114 VN.n40 VN.n39 12.1722
R115 VN.n41 VN.n40 12.1722
R116 VN.n70 VN.n69 12.1722
R117 VN.n96 VN.n95 12.1722
R118 VN.n95 VN.n94 12.1722
R119 VN.n68 VN.n67 2.54519
R120 VN.n13 VN.n12 2.54519
R121 VN.n109 VN.n55 0.417764
R122 VN.n54 VN.n0 0.417764
R123 VN VN.n54 0.394061
R124 VN.n105 VN.n55 0.189894
R125 VN.n105 VN.n104 0.189894
R126 VN.n104 VN.n103 0.189894
R127 VN.n103 VN.n57 0.189894
R128 VN.n99 VN.n57 0.189894
R129 VN.n99 VN.n98 0.189894
R130 VN.n98 VN.n97 0.189894
R131 VN.n97 VN.n59 0.189894
R132 VN.n92 VN.n59 0.189894
R133 VN.n92 VN.n91 0.189894
R134 VN.n91 VN.n90 0.189894
R135 VN.n90 VN.n61 0.189894
R136 VN.n86 VN.n61 0.189894
R137 VN.n86 VN.n85 0.189894
R138 VN.n85 VN.n84 0.189894
R139 VN.n84 VN.n63 0.189894
R140 VN.n80 VN.n63 0.189894
R141 VN.n80 VN.n79 0.189894
R142 VN.n79 VN.n78 0.189894
R143 VN.n78 VN.n65 0.189894
R144 VN.n74 VN.n65 0.189894
R145 VN.n74 VN.n73 0.189894
R146 VN.n73 VN.n72 0.189894
R147 VN.n72 VN.n67 0.189894
R148 VN.n17 VN.n12 0.189894
R149 VN.n18 VN.n17 0.189894
R150 VN.n19 VN.n18 0.189894
R151 VN.n19 VN.n10 0.189894
R152 VN.n23 VN.n10 0.189894
R153 VN.n24 VN.n23 0.189894
R154 VN.n25 VN.n24 0.189894
R155 VN.n25 VN.n8 0.189894
R156 VN.n29 VN.n8 0.189894
R157 VN.n30 VN.n29 0.189894
R158 VN.n31 VN.n30 0.189894
R159 VN.n31 VN.n6 0.189894
R160 VN.n35 VN.n6 0.189894
R161 VN.n36 VN.n35 0.189894
R162 VN.n37 VN.n36 0.189894
R163 VN.n37 VN.n4 0.189894
R164 VN.n42 VN.n4 0.189894
R165 VN.n43 VN.n42 0.189894
R166 VN.n44 VN.n43 0.189894
R167 VN.n44 VN.n2 0.189894
R168 VN.n48 VN.n2 0.189894
R169 VN.n49 VN.n48 0.189894
R170 VN.n50 VN.n49 0.189894
R171 VN.n50 VN.n0 0.189894
R172 VTAIL.n11 VTAIL.t13 57.4191
R173 VTAIL.n17 VTAIL.t11 57.419
R174 VTAIL.n2 VTAIL.t4 57.419
R175 VTAIL.n16 VTAIL.t7 57.419
R176 VTAIL.n15 VTAIL.n14 54.7936
R177 VTAIL.n13 VTAIL.n12 54.7936
R178 VTAIL.n10 VTAIL.n9 54.7936
R179 VTAIL.n8 VTAIL.n7 54.7936
R180 VTAIL.n19 VTAIL.n18 54.7933
R181 VTAIL.n1 VTAIL.n0 54.7933
R182 VTAIL.n4 VTAIL.n3 54.7933
R183 VTAIL.n6 VTAIL.n5 54.7933
R184 VTAIL.n8 VTAIL.n6 30.3669
R185 VTAIL.n17 VTAIL.n16 26.7031
R186 VTAIL.n10 VTAIL.n8 3.66429
R187 VTAIL.n11 VTAIL.n10 3.66429
R188 VTAIL.n15 VTAIL.n13 3.66429
R189 VTAIL.n16 VTAIL.n15 3.66429
R190 VTAIL.n6 VTAIL.n4 3.66429
R191 VTAIL.n4 VTAIL.n2 3.66429
R192 VTAIL.n19 VTAIL.n17 3.66429
R193 VTAIL VTAIL.n1 2.80653
R194 VTAIL.n18 VTAIL.t16 2.62611
R195 VTAIL.n18 VTAIL.t17 2.62611
R196 VTAIL.n0 VTAIL.t15 2.62611
R197 VTAIL.n0 VTAIL.t18 2.62611
R198 VTAIL.n3 VTAIL.t3 2.62611
R199 VTAIL.n3 VTAIL.t2 2.62611
R200 VTAIL.n5 VTAIL.t5 2.62611
R201 VTAIL.n5 VTAIL.t8 2.62611
R202 VTAIL.n14 VTAIL.t1 2.62611
R203 VTAIL.n14 VTAIL.t9 2.62611
R204 VTAIL.n12 VTAIL.t0 2.62611
R205 VTAIL.n12 VTAIL.t6 2.62611
R206 VTAIL.n9 VTAIL.t14 2.62611
R207 VTAIL.n9 VTAIL.t12 2.62611
R208 VTAIL.n7 VTAIL.t19 2.62611
R209 VTAIL.n7 VTAIL.t10 2.62611
R210 VTAIL.n13 VTAIL.n11 2.30222
R211 VTAIL.n2 VTAIL.n1 2.30222
R212 VTAIL VTAIL.n19 0.858259
R213 VDD2.n1 VDD2.t6 77.7616
R214 VDD2.n3 VDD2.n2 74.1646
R215 VDD2 VDD2.n7 74.1618
R216 VDD2.n4 VDD2.t0 74.0979
R217 VDD2.n6 VDD2.n5 71.4724
R218 VDD2.n1 VDD2.n0 71.4721
R219 VDD2.n4 VDD2.n3 51.7907
R220 VDD2.n6 VDD2.n4 3.66429
R221 VDD2.n7 VDD2.t2 2.62611
R222 VDD2.n7 VDD2.t8 2.62611
R223 VDD2.n5 VDD2.t5 2.62611
R224 VDD2.n5 VDD2.t7 2.62611
R225 VDD2.n2 VDD2.t3 2.62611
R226 VDD2.n2 VDD2.t9 2.62611
R227 VDD2.n0 VDD2.t4 2.62611
R228 VDD2.n0 VDD2.t1 2.62611
R229 VDD2 VDD2.n6 0.974638
R230 VDD2.n3 VDD2.n1 0.861102
R231 VP.n32 VP.n29 161.3
R232 VP.n34 VP.n33 161.3
R233 VP.n35 VP.n28 161.3
R234 VP.n37 VP.n36 161.3
R235 VP.n38 VP.n27 161.3
R236 VP.n40 VP.n39 161.3
R237 VP.n41 VP.n26 161.3
R238 VP.n43 VP.n42 161.3
R239 VP.n44 VP.n25 161.3
R240 VP.n46 VP.n45 161.3
R241 VP.n47 VP.n24 161.3
R242 VP.n49 VP.n48 161.3
R243 VP.n50 VP.n23 161.3
R244 VP.n52 VP.n51 161.3
R245 VP.n53 VP.n22 161.3
R246 VP.n55 VP.n54 161.3
R247 VP.n56 VP.n21 161.3
R248 VP.n59 VP.n58 161.3
R249 VP.n60 VP.n20 161.3
R250 VP.n62 VP.n61 161.3
R251 VP.n63 VP.n19 161.3
R252 VP.n65 VP.n64 161.3
R253 VP.n66 VP.n18 161.3
R254 VP.n68 VP.n67 161.3
R255 VP.n69 VP.n17 161.3
R256 VP.n124 VP.n0 161.3
R257 VP.n123 VP.n122 161.3
R258 VP.n121 VP.n1 161.3
R259 VP.n120 VP.n119 161.3
R260 VP.n118 VP.n2 161.3
R261 VP.n117 VP.n116 161.3
R262 VP.n115 VP.n3 161.3
R263 VP.n114 VP.n113 161.3
R264 VP.n111 VP.n4 161.3
R265 VP.n110 VP.n109 161.3
R266 VP.n108 VP.n5 161.3
R267 VP.n107 VP.n106 161.3
R268 VP.n105 VP.n6 161.3
R269 VP.n104 VP.n103 161.3
R270 VP.n102 VP.n7 161.3
R271 VP.n101 VP.n100 161.3
R272 VP.n99 VP.n8 161.3
R273 VP.n98 VP.n97 161.3
R274 VP.n96 VP.n9 161.3
R275 VP.n95 VP.n94 161.3
R276 VP.n93 VP.n10 161.3
R277 VP.n92 VP.n91 161.3
R278 VP.n90 VP.n11 161.3
R279 VP.n89 VP.n88 161.3
R280 VP.n87 VP.n12 161.3
R281 VP.n85 VP.n84 161.3
R282 VP.n83 VP.n13 161.3
R283 VP.n82 VP.n81 161.3
R284 VP.n80 VP.n14 161.3
R285 VP.n79 VP.n78 161.3
R286 VP.n77 VP.n15 161.3
R287 VP.n76 VP.n75 161.3
R288 VP.n74 VP.n16 161.3
R289 VP.n30 VP.t2 108.031
R290 VP.n125 VP.t4 76.1122
R291 VP.n99 VP.t9 76.1122
R292 VP.n73 VP.t0 76.1122
R293 VP.n86 VP.t8 76.1122
R294 VP.n112 VP.t5 76.1122
R295 VP.n44 VP.t6 76.1122
R296 VP.n70 VP.t1 76.1122
R297 VP.n57 VP.t7 76.1122
R298 VP.n31 VP.t3 76.1122
R299 VP.n31 VP.n30 62.7547
R300 VP.n72 VP.n71 60.871
R301 VP.n73 VP.n72 57.6421
R302 VP.n126 VP.n125 57.6421
R303 VP.n71 VP.n70 57.6421
R304 VP.n80 VP.n79 52.5823
R305 VP.n93 VP.n92 52.5823
R306 VP.n106 VP.n105 52.5823
R307 VP.n119 VP.n118 52.5823
R308 VP.n64 VP.n63 52.5823
R309 VP.n51 VP.n50 52.5823
R310 VP.n38 VP.n37 52.5823
R311 VP.n79 VP.n15 28.2389
R312 VP.n94 VP.n93 28.2389
R313 VP.n105 VP.n104 28.2389
R314 VP.n119 VP.n1 28.2389
R315 VP.n64 VP.n18 28.2389
R316 VP.n50 VP.n49 28.2389
R317 VP.n39 VP.n38 28.2389
R318 VP.n74 VP.n73 24.3439
R319 VP.n75 VP.n74 24.3439
R320 VP.n75 VP.n15 24.3439
R321 VP.n81 VP.n80 24.3439
R322 VP.n81 VP.n13 24.3439
R323 VP.n85 VP.n13 24.3439
R324 VP.n88 VP.n87 24.3439
R325 VP.n88 VP.n11 24.3439
R326 VP.n92 VP.n11 24.3439
R327 VP.n94 VP.n9 24.3439
R328 VP.n98 VP.n9 24.3439
R329 VP.n99 VP.n98 24.3439
R330 VP.n100 VP.n99 24.3439
R331 VP.n100 VP.n7 24.3439
R332 VP.n104 VP.n7 24.3439
R333 VP.n106 VP.n5 24.3439
R334 VP.n110 VP.n5 24.3439
R335 VP.n111 VP.n110 24.3439
R336 VP.n113 VP.n3 24.3439
R337 VP.n117 VP.n3 24.3439
R338 VP.n118 VP.n117 24.3439
R339 VP.n123 VP.n1 24.3439
R340 VP.n124 VP.n123 24.3439
R341 VP.n125 VP.n124 24.3439
R342 VP.n68 VP.n18 24.3439
R343 VP.n69 VP.n68 24.3439
R344 VP.n70 VP.n69 24.3439
R345 VP.n51 VP.n22 24.3439
R346 VP.n55 VP.n22 24.3439
R347 VP.n56 VP.n55 24.3439
R348 VP.n58 VP.n20 24.3439
R349 VP.n62 VP.n20 24.3439
R350 VP.n63 VP.n62 24.3439
R351 VP.n39 VP.n26 24.3439
R352 VP.n43 VP.n26 24.3439
R353 VP.n44 VP.n43 24.3439
R354 VP.n45 VP.n44 24.3439
R355 VP.n45 VP.n24 24.3439
R356 VP.n49 VP.n24 24.3439
R357 VP.n33 VP.n32 24.3439
R358 VP.n33 VP.n28 24.3439
R359 VP.n37 VP.n28 24.3439
R360 VP.n86 VP.n85 12.1722
R361 VP.n87 VP.n86 12.1722
R362 VP.n112 VP.n111 12.1722
R363 VP.n113 VP.n112 12.1722
R364 VP.n57 VP.n56 12.1722
R365 VP.n58 VP.n57 12.1722
R366 VP.n32 VP.n31 12.1722
R367 VP.n30 VP.n29 2.54517
R368 VP.n71 VP.n17 0.417764
R369 VP.n72 VP.n16 0.417764
R370 VP.n126 VP.n0 0.417764
R371 VP VP.n126 0.394061
R372 VP.n34 VP.n29 0.189894
R373 VP.n35 VP.n34 0.189894
R374 VP.n36 VP.n35 0.189894
R375 VP.n36 VP.n27 0.189894
R376 VP.n40 VP.n27 0.189894
R377 VP.n41 VP.n40 0.189894
R378 VP.n42 VP.n41 0.189894
R379 VP.n42 VP.n25 0.189894
R380 VP.n46 VP.n25 0.189894
R381 VP.n47 VP.n46 0.189894
R382 VP.n48 VP.n47 0.189894
R383 VP.n48 VP.n23 0.189894
R384 VP.n52 VP.n23 0.189894
R385 VP.n53 VP.n52 0.189894
R386 VP.n54 VP.n53 0.189894
R387 VP.n54 VP.n21 0.189894
R388 VP.n59 VP.n21 0.189894
R389 VP.n60 VP.n59 0.189894
R390 VP.n61 VP.n60 0.189894
R391 VP.n61 VP.n19 0.189894
R392 VP.n65 VP.n19 0.189894
R393 VP.n66 VP.n65 0.189894
R394 VP.n67 VP.n66 0.189894
R395 VP.n67 VP.n17 0.189894
R396 VP.n76 VP.n16 0.189894
R397 VP.n77 VP.n76 0.189894
R398 VP.n78 VP.n77 0.189894
R399 VP.n78 VP.n14 0.189894
R400 VP.n82 VP.n14 0.189894
R401 VP.n83 VP.n82 0.189894
R402 VP.n84 VP.n83 0.189894
R403 VP.n84 VP.n12 0.189894
R404 VP.n89 VP.n12 0.189894
R405 VP.n90 VP.n89 0.189894
R406 VP.n91 VP.n90 0.189894
R407 VP.n91 VP.n10 0.189894
R408 VP.n95 VP.n10 0.189894
R409 VP.n96 VP.n95 0.189894
R410 VP.n97 VP.n96 0.189894
R411 VP.n97 VP.n8 0.189894
R412 VP.n101 VP.n8 0.189894
R413 VP.n102 VP.n101 0.189894
R414 VP.n103 VP.n102 0.189894
R415 VP.n103 VP.n6 0.189894
R416 VP.n107 VP.n6 0.189894
R417 VP.n108 VP.n107 0.189894
R418 VP.n109 VP.n108 0.189894
R419 VP.n109 VP.n4 0.189894
R420 VP.n114 VP.n4 0.189894
R421 VP.n115 VP.n114 0.189894
R422 VP.n116 VP.n115 0.189894
R423 VP.n116 VP.n2 0.189894
R424 VP.n120 VP.n2 0.189894
R425 VP.n121 VP.n120 0.189894
R426 VP.n122 VP.n121 0.189894
R427 VP.n122 VP.n0 0.189894
R428 VDD1.n1 VDD1.t7 77.7617
R429 VDD1.n3 VDD1.t9 77.7616
R430 VDD1.n5 VDD1.n4 74.1646
R431 VDD1.n1 VDD1.n0 71.4724
R432 VDD1.n7 VDD1.n6 71.4722
R433 VDD1.n3 VDD1.n2 71.4721
R434 VDD1.n7 VDD1.n5 54.2056
R435 VDD1 VDD1.n7 2.69016
R436 VDD1.n6 VDD1.t2 2.62611
R437 VDD1.n6 VDD1.t8 2.62611
R438 VDD1.n0 VDD1.t6 2.62611
R439 VDD1.n0 VDD1.t3 2.62611
R440 VDD1.n4 VDD1.t4 2.62611
R441 VDD1.n4 VDD1.t5 2.62611
R442 VDD1.n2 VDD1.t1 2.62611
R443 VDD1.n2 VDD1.t0 2.62611
R444 VDD1 VDD1.n1 0.974638
R445 VDD1.n5 VDD1.n3 0.861102
R446 B.n790 B.n789 585
R447 B.n791 B.n94 585
R448 B.n793 B.n792 585
R449 B.n794 B.n93 585
R450 B.n796 B.n795 585
R451 B.n797 B.n92 585
R452 B.n799 B.n798 585
R453 B.n800 B.n91 585
R454 B.n802 B.n801 585
R455 B.n803 B.n90 585
R456 B.n805 B.n804 585
R457 B.n806 B.n89 585
R458 B.n808 B.n807 585
R459 B.n809 B.n88 585
R460 B.n811 B.n810 585
R461 B.n812 B.n87 585
R462 B.n814 B.n813 585
R463 B.n815 B.n86 585
R464 B.n817 B.n816 585
R465 B.n818 B.n85 585
R466 B.n820 B.n819 585
R467 B.n821 B.n84 585
R468 B.n823 B.n822 585
R469 B.n824 B.n83 585
R470 B.n826 B.n825 585
R471 B.n827 B.n82 585
R472 B.n829 B.n828 585
R473 B.n830 B.n81 585
R474 B.n832 B.n831 585
R475 B.n833 B.n80 585
R476 B.n835 B.n834 585
R477 B.n836 B.n79 585
R478 B.n838 B.n837 585
R479 B.n839 B.n78 585
R480 B.n841 B.n840 585
R481 B.n842 B.n77 585
R482 B.n844 B.n843 585
R483 B.n845 B.n76 585
R484 B.n847 B.n846 585
R485 B.n848 B.n75 585
R486 B.n850 B.n849 585
R487 B.n851 B.n74 585
R488 B.n853 B.n852 585
R489 B.n855 B.n71 585
R490 B.n857 B.n856 585
R491 B.n858 B.n70 585
R492 B.n860 B.n859 585
R493 B.n861 B.n69 585
R494 B.n863 B.n862 585
R495 B.n864 B.n68 585
R496 B.n866 B.n865 585
R497 B.n867 B.n65 585
R498 B.n870 B.n869 585
R499 B.n871 B.n64 585
R500 B.n873 B.n872 585
R501 B.n874 B.n63 585
R502 B.n876 B.n875 585
R503 B.n877 B.n62 585
R504 B.n879 B.n878 585
R505 B.n880 B.n61 585
R506 B.n882 B.n881 585
R507 B.n883 B.n60 585
R508 B.n885 B.n884 585
R509 B.n886 B.n59 585
R510 B.n888 B.n887 585
R511 B.n889 B.n58 585
R512 B.n891 B.n890 585
R513 B.n892 B.n57 585
R514 B.n894 B.n893 585
R515 B.n895 B.n56 585
R516 B.n897 B.n896 585
R517 B.n898 B.n55 585
R518 B.n900 B.n899 585
R519 B.n901 B.n54 585
R520 B.n903 B.n902 585
R521 B.n904 B.n53 585
R522 B.n906 B.n905 585
R523 B.n907 B.n52 585
R524 B.n909 B.n908 585
R525 B.n910 B.n51 585
R526 B.n912 B.n911 585
R527 B.n913 B.n50 585
R528 B.n915 B.n914 585
R529 B.n916 B.n49 585
R530 B.n918 B.n917 585
R531 B.n919 B.n48 585
R532 B.n921 B.n920 585
R533 B.n922 B.n47 585
R534 B.n924 B.n923 585
R535 B.n925 B.n46 585
R536 B.n927 B.n926 585
R537 B.n928 B.n45 585
R538 B.n930 B.n929 585
R539 B.n931 B.n44 585
R540 B.n933 B.n932 585
R541 B.n788 B.n95 585
R542 B.n787 B.n786 585
R543 B.n785 B.n96 585
R544 B.n784 B.n783 585
R545 B.n782 B.n97 585
R546 B.n781 B.n780 585
R547 B.n779 B.n98 585
R548 B.n778 B.n777 585
R549 B.n776 B.n99 585
R550 B.n775 B.n774 585
R551 B.n773 B.n100 585
R552 B.n772 B.n771 585
R553 B.n770 B.n101 585
R554 B.n769 B.n768 585
R555 B.n767 B.n102 585
R556 B.n766 B.n765 585
R557 B.n764 B.n103 585
R558 B.n763 B.n762 585
R559 B.n761 B.n104 585
R560 B.n760 B.n759 585
R561 B.n758 B.n105 585
R562 B.n757 B.n756 585
R563 B.n755 B.n106 585
R564 B.n754 B.n753 585
R565 B.n752 B.n107 585
R566 B.n751 B.n750 585
R567 B.n749 B.n108 585
R568 B.n748 B.n747 585
R569 B.n746 B.n109 585
R570 B.n745 B.n744 585
R571 B.n743 B.n110 585
R572 B.n742 B.n741 585
R573 B.n740 B.n111 585
R574 B.n739 B.n738 585
R575 B.n737 B.n112 585
R576 B.n736 B.n735 585
R577 B.n734 B.n113 585
R578 B.n733 B.n732 585
R579 B.n731 B.n114 585
R580 B.n730 B.n729 585
R581 B.n728 B.n115 585
R582 B.n727 B.n726 585
R583 B.n725 B.n116 585
R584 B.n724 B.n723 585
R585 B.n722 B.n117 585
R586 B.n721 B.n720 585
R587 B.n719 B.n118 585
R588 B.n718 B.n717 585
R589 B.n716 B.n119 585
R590 B.n715 B.n714 585
R591 B.n713 B.n120 585
R592 B.n712 B.n711 585
R593 B.n710 B.n121 585
R594 B.n709 B.n708 585
R595 B.n707 B.n122 585
R596 B.n706 B.n705 585
R597 B.n704 B.n123 585
R598 B.n703 B.n702 585
R599 B.n701 B.n124 585
R600 B.n700 B.n699 585
R601 B.n698 B.n125 585
R602 B.n697 B.n696 585
R603 B.n695 B.n126 585
R604 B.n694 B.n693 585
R605 B.n692 B.n127 585
R606 B.n691 B.n690 585
R607 B.n689 B.n128 585
R608 B.n688 B.n687 585
R609 B.n686 B.n129 585
R610 B.n685 B.n684 585
R611 B.n683 B.n130 585
R612 B.n682 B.n681 585
R613 B.n680 B.n131 585
R614 B.n679 B.n678 585
R615 B.n677 B.n132 585
R616 B.n676 B.n675 585
R617 B.n674 B.n133 585
R618 B.n673 B.n672 585
R619 B.n671 B.n134 585
R620 B.n670 B.n669 585
R621 B.n668 B.n135 585
R622 B.n667 B.n666 585
R623 B.n665 B.n136 585
R624 B.n664 B.n663 585
R625 B.n662 B.n137 585
R626 B.n661 B.n660 585
R627 B.n659 B.n138 585
R628 B.n658 B.n657 585
R629 B.n656 B.n139 585
R630 B.n655 B.n654 585
R631 B.n653 B.n140 585
R632 B.n652 B.n651 585
R633 B.n650 B.n141 585
R634 B.n649 B.n648 585
R635 B.n647 B.n142 585
R636 B.n646 B.n645 585
R637 B.n644 B.n143 585
R638 B.n643 B.n642 585
R639 B.n641 B.n144 585
R640 B.n640 B.n639 585
R641 B.n638 B.n145 585
R642 B.n637 B.n636 585
R643 B.n635 B.n146 585
R644 B.n634 B.n633 585
R645 B.n632 B.n147 585
R646 B.n631 B.n630 585
R647 B.n629 B.n148 585
R648 B.n628 B.n627 585
R649 B.n626 B.n149 585
R650 B.n625 B.n624 585
R651 B.n623 B.n150 585
R652 B.n622 B.n621 585
R653 B.n620 B.n151 585
R654 B.n619 B.n618 585
R655 B.n617 B.n152 585
R656 B.n616 B.n615 585
R657 B.n614 B.n153 585
R658 B.n613 B.n612 585
R659 B.n611 B.n154 585
R660 B.n610 B.n609 585
R661 B.n608 B.n155 585
R662 B.n607 B.n606 585
R663 B.n605 B.n156 585
R664 B.n604 B.n603 585
R665 B.n602 B.n157 585
R666 B.n601 B.n600 585
R667 B.n599 B.n158 585
R668 B.n598 B.n597 585
R669 B.n596 B.n159 585
R670 B.n595 B.n594 585
R671 B.n593 B.n160 585
R672 B.n592 B.n591 585
R673 B.n590 B.n161 585
R674 B.n589 B.n588 585
R675 B.n587 B.n162 585
R676 B.n586 B.n585 585
R677 B.n584 B.n163 585
R678 B.n583 B.n582 585
R679 B.n581 B.n164 585
R680 B.n580 B.n579 585
R681 B.n578 B.n165 585
R682 B.n577 B.n576 585
R683 B.n575 B.n166 585
R684 B.n574 B.n573 585
R685 B.n572 B.n167 585
R686 B.n571 B.n570 585
R687 B.n569 B.n168 585
R688 B.n568 B.n567 585
R689 B.n566 B.n169 585
R690 B.n565 B.n564 585
R691 B.n563 B.n170 585
R692 B.n562 B.n561 585
R693 B.n560 B.n171 585
R694 B.n559 B.n558 585
R695 B.n557 B.n172 585
R696 B.n556 B.n555 585
R697 B.n554 B.n173 585
R698 B.n553 B.n552 585
R699 B.n551 B.n174 585
R700 B.n550 B.n549 585
R701 B.n548 B.n175 585
R702 B.n547 B.n546 585
R703 B.n545 B.n176 585
R704 B.n544 B.n543 585
R705 B.n542 B.n177 585
R706 B.n541 B.n540 585
R707 B.n539 B.n178 585
R708 B.n395 B.n230 585
R709 B.n397 B.n396 585
R710 B.n398 B.n229 585
R711 B.n400 B.n399 585
R712 B.n401 B.n228 585
R713 B.n403 B.n402 585
R714 B.n404 B.n227 585
R715 B.n406 B.n405 585
R716 B.n407 B.n226 585
R717 B.n409 B.n408 585
R718 B.n410 B.n225 585
R719 B.n412 B.n411 585
R720 B.n413 B.n224 585
R721 B.n415 B.n414 585
R722 B.n416 B.n223 585
R723 B.n418 B.n417 585
R724 B.n419 B.n222 585
R725 B.n421 B.n420 585
R726 B.n422 B.n221 585
R727 B.n424 B.n423 585
R728 B.n425 B.n220 585
R729 B.n427 B.n426 585
R730 B.n428 B.n219 585
R731 B.n430 B.n429 585
R732 B.n431 B.n218 585
R733 B.n433 B.n432 585
R734 B.n434 B.n217 585
R735 B.n436 B.n435 585
R736 B.n437 B.n216 585
R737 B.n439 B.n438 585
R738 B.n440 B.n215 585
R739 B.n442 B.n441 585
R740 B.n443 B.n214 585
R741 B.n445 B.n444 585
R742 B.n446 B.n213 585
R743 B.n448 B.n447 585
R744 B.n449 B.n212 585
R745 B.n451 B.n450 585
R746 B.n452 B.n211 585
R747 B.n454 B.n453 585
R748 B.n455 B.n210 585
R749 B.n457 B.n456 585
R750 B.n458 B.n207 585
R751 B.n461 B.n460 585
R752 B.n462 B.n206 585
R753 B.n464 B.n463 585
R754 B.n465 B.n205 585
R755 B.n467 B.n466 585
R756 B.n468 B.n204 585
R757 B.n470 B.n469 585
R758 B.n471 B.n203 585
R759 B.n473 B.n472 585
R760 B.n475 B.n474 585
R761 B.n476 B.n199 585
R762 B.n478 B.n477 585
R763 B.n479 B.n198 585
R764 B.n481 B.n480 585
R765 B.n482 B.n197 585
R766 B.n484 B.n483 585
R767 B.n485 B.n196 585
R768 B.n487 B.n486 585
R769 B.n488 B.n195 585
R770 B.n490 B.n489 585
R771 B.n491 B.n194 585
R772 B.n493 B.n492 585
R773 B.n494 B.n193 585
R774 B.n496 B.n495 585
R775 B.n497 B.n192 585
R776 B.n499 B.n498 585
R777 B.n500 B.n191 585
R778 B.n502 B.n501 585
R779 B.n503 B.n190 585
R780 B.n505 B.n504 585
R781 B.n506 B.n189 585
R782 B.n508 B.n507 585
R783 B.n509 B.n188 585
R784 B.n511 B.n510 585
R785 B.n512 B.n187 585
R786 B.n514 B.n513 585
R787 B.n515 B.n186 585
R788 B.n517 B.n516 585
R789 B.n518 B.n185 585
R790 B.n520 B.n519 585
R791 B.n521 B.n184 585
R792 B.n523 B.n522 585
R793 B.n524 B.n183 585
R794 B.n526 B.n525 585
R795 B.n527 B.n182 585
R796 B.n529 B.n528 585
R797 B.n530 B.n181 585
R798 B.n532 B.n531 585
R799 B.n533 B.n180 585
R800 B.n535 B.n534 585
R801 B.n536 B.n179 585
R802 B.n538 B.n537 585
R803 B.n394 B.n393 585
R804 B.n392 B.n231 585
R805 B.n391 B.n390 585
R806 B.n389 B.n232 585
R807 B.n388 B.n387 585
R808 B.n386 B.n233 585
R809 B.n385 B.n384 585
R810 B.n383 B.n234 585
R811 B.n382 B.n381 585
R812 B.n380 B.n235 585
R813 B.n379 B.n378 585
R814 B.n377 B.n236 585
R815 B.n376 B.n375 585
R816 B.n374 B.n237 585
R817 B.n373 B.n372 585
R818 B.n371 B.n238 585
R819 B.n370 B.n369 585
R820 B.n368 B.n239 585
R821 B.n367 B.n366 585
R822 B.n365 B.n240 585
R823 B.n364 B.n363 585
R824 B.n362 B.n241 585
R825 B.n361 B.n360 585
R826 B.n359 B.n242 585
R827 B.n358 B.n357 585
R828 B.n356 B.n243 585
R829 B.n355 B.n354 585
R830 B.n353 B.n244 585
R831 B.n352 B.n351 585
R832 B.n350 B.n245 585
R833 B.n349 B.n348 585
R834 B.n347 B.n246 585
R835 B.n346 B.n345 585
R836 B.n344 B.n247 585
R837 B.n343 B.n342 585
R838 B.n341 B.n248 585
R839 B.n340 B.n339 585
R840 B.n338 B.n249 585
R841 B.n337 B.n336 585
R842 B.n335 B.n250 585
R843 B.n334 B.n333 585
R844 B.n332 B.n251 585
R845 B.n331 B.n330 585
R846 B.n329 B.n252 585
R847 B.n328 B.n327 585
R848 B.n326 B.n253 585
R849 B.n325 B.n324 585
R850 B.n323 B.n254 585
R851 B.n322 B.n321 585
R852 B.n320 B.n255 585
R853 B.n319 B.n318 585
R854 B.n317 B.n256 585
R855 B.n316 B.n315 585
R856 B.n314 B.n257 585
R857 B.n313 B.n312 585
R858 B.n311 B.n258 585
R859 B.n310 B.n309 585
R860 B.n308 B.n259 585
R861 B.n307 B.n306 585
R862 B.n305 B.n260 585
R863 B.n304 B.n303 585
R864 B.n302 B.n261 585
R865 B.n301 B.n300 585
R866 B.n299 B.n262 585
R867 B.n298 B.n297 585
R868 B.n296 B.n263 585
R869 B.n295 B.n294 585
R870 B.n293 B.n264 585
R871 B.n292 B.n291 585
R872 B.n290 B.n265 585
R873 B.n289 B.n288 585
R874 B.n287 B.n266 585
R875 B.n286 B.n285 585
R876 B.n284 B.n267 585
R877 B.n283 B.n282 585
R878 B.n281 B.n268 585
R879 B.n280 B.n279 585
R880 B.n278 B.n269 585
R881 B.n277 B.n276 585
R882 B.n275 B.n270 585
R883 B.n274 B.n273 585
R884 B.n272 B.n271 585
R885 B.n2 B.n0 585
R886 B.n1057 B.n1 585
R887 B.n1056 B.n1055 585
R888 B.n1054 B.n3 585
R889 B.n1053 B.n1052 585
R890 B.n1051 B.n4 585
R891 B.n1050 B.n1049 585
R892 B.n1048 B.n5 585
R893 B.n1047 B.n1046 585
R894 B.n1045 B.n6 585
R895 B.n1044 B.n1043 585
R896 B.n1042 B.n7 585
R897 B.n1041 B.n1040 585
R898 B.n1039 B.n8 585
R899 B.n1038 B.n1037 585
R900 B.n1036 B.n9 585
R901 B.n1035 B.n1034 585
R902 B.n1033 B.n10 585
R903 B.n1032 B.n1031 585
R904 B.n1030 B.n11 585
R905 B.n1029 B.n1028 585
R906 B.n1027 B.n12 585
R907 B.n1026 B.n1025 585
R908 B.n1024 B.n13 585
R909 B.n1023 B.n1022 585
R910 B.n1021 B.n14 585
R911 B.n1020 B.n1019 585
R912 B.n1018 B.n15 585
R913 B.n1017 B.n1016 585
R914 B.n1015 B.n16 585
R915 B.n1014 B.n1013 585
R916 B.n1012 B.n17 585
R917 B.n1011 B.n1010 585
R918 B.n1009 B.n18 585
R919 B.n1008 B.n1007 585
R920 B.n1006 B.n19 585
R921 B.n1005 B.n1004 585
R922 B.n1003 B.n20 585
R923 B.n1002 B.n1001 585
R924 B.n1000 B.n21 585
R925 B.n999 B.n998 585
R926 B.n997 B.n22 585
R927 B.n996 B.n995 585
R928 B.n994 B.n23 585
R929 B.n993 B.n992 585
R930 B.n991 B.n24 585
R931 B.n990 B.n989 585
R932 B.n988 B.n25 585
R933 B.n987 B.n986 585
R934 B.n985 B.n26 585
R935 B.n984 B.n983 585
R936 B.n982 B.n27 585
R937 B.n981 B.n980 585
R938 B.n979 B.n28 585
R939 B.n978 B.n977 585
R940 B.n976 B.n29 585
R941 B.n975 B.n974 585
R942 B.n973 B.n30 585
R943 B.n972 B.n971 585
R944 B.n970 B.n31 585
R945 B.n969 B.n968 585
R946 B.n967 B.n32 585
R947 B.n966 B.n965 585
R948 B.n964 B.n33 585
R949 B.n963 B.n962 585
R950 B.n961 B.n34 585
R951 B.n960 B.n959 585
R952 B.n958 B.n35 585
R953 B.n957 B.n956 585
R954 B.n955 B.n36 585
R955 B.n954 B.n953 585
R956 B.n952 B.n37 585
R957 B.n951 B.n950 585
R958 B.n949 B.n38 585
R959 B.n948 B.n947 585
R960 B.n946 B.n39 585
R961 B.n945 B.n944 585
R962 B.n943 B.n40 585
R963 B.n942 B.n941 585
R964 B.n940 B.n41 585
R965 B.n939 B.n938 585
R966 B.n937 B.n42 585
R967 B.n936 B.n935 585
R968 B.n934 B.n43 585
R969 B.n1059 B.n1058 585
R970 B.n395 B.n394 521.33
R971 B.n932 B.n43 521.33
R972 B.n539 B.n538 521.33
R973 B.n790 B.n95 521.33
R974 B.n200 B.t9 285.546
R975 B.n208 B.t6 285.546
R976 B.n66 B.t3 285.546
R977 B.n72 B.t0 285.546
R978 B.n200 B.t11 192.16
R979 B.n72 B.t1 192.16
R980 B.n208 B.t8 192.144
R981 B.n66 B.t4 192.144
R982 B.n394 B.n231 163.367
R983 B.n390 B.n231 163.367
R984 B.n390 B.n389 163.367
R985 B.n389 B.n388 163.367
R986 B.n388 B.n233 163.367
R987 B.n384 B.n233 163.367
R988 B.n384 B.n383 163.367
R989 B.n383 B.n382 163.367
R990 B.n382 B.n235 163.367
R991 B.n378 B.n235 163.367
R992 B.n378 B.n377 163.367
R993 B.n377 B.n376 163.367
R994 B.n376 B.n237 163.367
R995 B.n372 B.n237 163.367
R996 B.n372 B.n371 163.367
R997 B.n371 B.n370 163.367
R998 B.n370 B.n239 163.367
R999 B.n366 B.n239 163.367
R1000 B.n366 B.n365 163.367
R1001 B.n365 B.n364 163.367
R1002 B.n364 B.n241 163.367
R1003 B.n360 B.n241 163.367
R1004 B.n360 B.n359 163.367
R1005 B.n359 B.n358 163.367
R1006 B.n358 B.n243 163.367
R1007 B.n354 B.n243 163.367
R1008 B.n354 B.n353 163.367
R1009 B.n353 B.n352 163.367
R1010 B.n352 B.n245 163.367
R1011 B.n348 B.n245 163.367
R1012 B.n348 B.n347 163.367
R1013 B.n347 B.n346 163.367
R1014 B.n346 B.n247 163.367
R1015 B.n342 B.n247 163.367
R1016 B.n342 B.n341 163.367
R1017 B.n341 B.n340 163.367
R1018 B.n340 B.n249 163.367
R1019 B.n336 B.n249 163.367
R1020 B.n336 B.n335 163.367
R1021 B.n335 B.n334 163.367
R1022 B.n334 B.n251 163.367
R1023 B.n330 B.n251 163.367
R1024 B.n330 B.n329 163.367
R1025 B.n329 B.n328 163.367
R1026 B.n328 B.n253 163.367
R1027 B.n324 B.n253 163.367
R1028 B.n324 B.n323 163.367
R1029 B.n323 B.n322 163.367
R1030 B.n322 B.n255 163.367
R1031 B.n318 B.n255 163.367
R1032 B.n318 B.n317 163.367
R1033 B.n317 B.n316 163.367
R1034 B.n316 B.n257 163.367
R1035 B.n312 B.n257 163.367
R1036 B.n312 B.n311 163.367
R1037 B.n311 B.n310 163.367
R1038 B.n310 B.n259 163.367
R1039 B.n306 B.n259 163.367
R1040 B.n306 B.n305 163.367
R1041 B.n305 B.n304 163.367
R1042 B.n304 B.n261 163.367
R1043 B.n300 B.n261 163.367
R1044 B.n300 B.n299 163.367
R1045 B.n299 B.n298 163.367
R1046 B.n298 B.n263 163.367
R1047 B.n294 B.n263 163.367
R1048 B.n294 B.n293 163.367
R1049 B.n293 B.n292 163.367
R1050 B.n292 B.n265 163.367
R1051 B.n288 B.n265 163.367
R1052 B.n288 B.n287 163.367
R1053 B.n287 B.n286 163.367
R1054 B.n286 B.n267 163.367
R1055 B.n282 B.n267 163.367
R1056 B.n282 B.n281 163.367
R1057 B.n281 B.n280 163.367
R1058 B.n280 B.n269 163.367
R1059 B.n276 B.n269 163.367
R1060 B.n276 B.n275 163.367
R1061 B.n275 B.n274 163.367
R1062 B.n274 B.n271 163.367
R1063 B.n271 B.n2 163.367
R1064 B.n1058 B.n2 163.367
R1065 B.n1058 B.n1057 163.367
R1066 B.n1057 B.n1056 163.367
R1067 B.n1056 B.n3 163.367
R1068 B.n1052 B.n3 163.367
R1069 B.n1052 B.n1051 163.367
R1070 B.n1051 B.n1050 163.367
R1071 B.n1050 B.n5 163.367
R1072 B.n1046 B.n5 163.367
R1073 B.n1046 B.n1045 163.367
R1074 B.n1045 B.n1044 163.367
R1075 B.n1044 B.n7 163.367
R1076 B.n1040 B.n7 163.367
R1077 B.n1040 B.n1039 163.367
R1078 B.n1039 B.n1038 163.367
R1079 B.n1038 B.n9 163.367
R1080 B.n1034 B.n9 163.367
R1081 B.n1034 B.n1033 163.367
R1082 B.n1033 B.n1032 163.367
R1083 B.n1032 B.n11 163.367
R1084 B.n1028 B.n11 163.367
R1085 B.n1028 B.n1027 163.367
R1086 B.n1027 B.n1026 163.367
R1087 B.n1026 B.n13 163.367
R1088 B.n1022 B.n13 163.367
R1089 B.n1022 B.n1021 163.367
R1090 B.n1021 B.n1020 163.367
R1091 B.n1020 B.n15 163.367
R1092 B.n1016 B.n15 163.367
R1093 B.n1016 B.n1015 163.367
R1094 B.n1015 B.n1014 163.367
R1095 B.n1014 B.n17 163.367
R1096 B.n1010 B.n17 163.367
R1097 B.n1010 B.n1009 163.367
R1098 B.n1009 B.n1008 163.367
R1099 B.n1008 B.n19 163.367
R1100 B.n1004 B.n19 163.367
R1101 B.n1004 B.n1003 163.367
R1102 B.n1003 B.n1002 163.367
R1103 B.n1002 B.n21 163.367
R1104 B.n998 B.n21 163.367
R1105 B.n998 B.n997 163.367
R1106 B.n997 B.n996 163.367
R1107 B.n996 B.n23 163.367
R1108 B.n992 B.n23 163.367
R1109 B.n992 B.n991 163.367
R1110 B.n991 B.n990 163.367
R1111 B.n990 B.n25 163.367
R1112 B.n986 B.n25 163.367
R1113 B.n986 B.n985 163.367
R1114 B.n985 B.n984 163.367
R1115 B.n984 B.n27 163.367
R1116 B.n980 B.n27 163.367
R1117 B.n980 B.n979 163.367
R1118 B.n979 B.n978 163.367
R1119 B.n978 B.n29 163.367
R1120 B.n974 B.n29 163.367
R1121 B.n974 B.n973 163.367
R1122 B.n973 B.n972 163.367
R1123 B.n972 B.n31 163.367
R1124 B.n968 B.n31 163.367
R1125 B.n968 B.n967 163.367
R1126 B.n967 B.n966 163.367
R1127 B.n966 B.n33 163.367
R1128 B.n962 B.n33 163.367
R1129 B.n962 B.n961 163.367
R1130 B.n961 B.n960 163.367
R1131 B.n960 B.n35 163.367
R1132 B.n956 B.n35 163.367
R1133 B.n956 B.n955 163.367
R1134 B.n955 B.n954 163.367
R1135 B.n954 B.n37 163.367
R1136 B.n950 B.n37 163.367
R1137 B.n950 B.n949 163.367
R1138 B.n949 B.n948 163.367
R1139 B.n948 B.n39 163.367
R1140 B.n944 B.n39 163.367
R1141 B.n944 B.n943 163.367
R1142 B.n943 B.n942 163.367
R1143 B.n942 B.n41 163.367
R1144 B.n938 B.n41 163.367
R1145 B.n938 B.n937 163.367
R1146 B.n937 B.n936 163.367
R1147 B.n936 B.n43 163.367
R1148 B.n396 B.n395 163.367
R1149 B.n396 B.n229 163.367
R1150 B.n400 B.n229 163.367
R1151 B.n401 B.n400 163.367
R1152 B.n402 B.n401 163.367
R1153 B.n402 B.n227 163.367
R1154 B.n406 B.n227 163.367
R1155 B.n407 B.n406 163.367
R1156 B.n408 B.n407 163.367
R1157 B.n408 B.n225 163.367
R1158 B.n412 B.n225 163.367
R1159 B.n413 B.n412 163.367
R1160 B.n414 B.n413 163.367
R1161 B.n414 B.n223 163.367
R1162 B.n418 B.n223 163.367
R1163 B.n419 B.n418 163.367
R1164 B.n420 B.n419 163.367
R1165 B.n420 B.n221 163.367
R1166 B.n424 B.n221 163.367
R1167 B.n425 B.n424 163.367
R1168 B.n426 B.n425 163.367
R1169 B.n426 B.n219 163.367
R1170 B.n430 B.n219 163.367
R1171 B.n431 B.n430 163.367
R1172 B.n432 B.n431 163.367
R1173 B.n432 B.n217 163.367
R1174 B.n436 B.n217 163.367
R1175 B.n437 B.n436 163.367
R1176 B.n438 B.n437 163.367
R1177 B.n438 B.n215 163.367
R1178 B.n442 B.n215 163.367
R1179 B.n443 B.n442 163.367
R1180 B.n444 B.n443 163.367
R1181 B.n444 B.n213 163.367
R1182 B.n448 B.n213 163.367
R1183 B.n449 B.n448 163.367
R1184 B.n450 B.n449 163.367
R1185 B.n450 B.n211 163.367
R1186 B.n454 B.n211 163.367
R1187 B.n455 B.n454 163.367
R1188 B.n456 B.n455 163.367
R1189 B.n456 B.n207 163.367
R1190 B.n461 B.n207 163.367
R1191 B.n462 B.n461 163.367
R1192 B.n463 B.n462 163.367
R1193 B.n463 B.n205 163.367
R1194 B.n467 B.n205 163.367
R1195 B.n468 B.n467 163.367
R1196 B.n469 B.n468 163.367
R1197 B.n469 B.n203 163.367
R1198 B.n473 B.n203 163.367
R1199 B.n474 B.n473 163.367
R1200 B.n474 B.n199 163.367
R1201 B.n478 B.n199 163.367
R1202 B.n479 B.n478 163.367
R1203 B.n480 B.n479 163.367
R1204 B.n480 B.n197 163.367
R1205 B.n484 B.n197 163.367
R1206 B.n485 B.n484 163.367
R1207 B.n486 B.n485 163.367
R1208 B.n486 B.n195 163.367
R1209 B.n490 B.n195 163.367
R1210 B.n491 B.n490 163.367
R1211 B.n492 B.n491 163.367
R1212 B.n492 B.n193 163.367
R1213 B.n496 B.n193 163.367
R1214 B.n497 B.n496 163.367
R1215 B.n498 B.n497 163.367
R1216 B.n498 B.n191 163.367
R1217 B.n502 B.n191 163.367
R1218 B.n503 B.n502 163.367
R1219 B.n504 B.n503 163.367
R1220 B.n504 B.n189 163.367
R1221 B.n508 B.n189 163.367
R1222 B.n509 B.n508 163.367
R1223 B.n510 B.n509 163.367
R1224 B.n510 B.n187 163.367
R1225 B.n514 B.n187 163.367
R1226 B.n515 B.n514 163.367
R1227 B.n516 B.n515 163.367
R1228 B.n516 B.n185 163.367
R1229 B.n520 B.n185 163.367
R1230 B.n521 B.n520 163.367
R1231 B.n522 B.n521 163.367
R1232 B.n522 B.n183 163.367
R1233 B.n526 B.n183 163.367
R1234 B.n527 B.n526 163.367
R1235 B.n528 B.n527 163.367
R1236 B.n528 B.n181 163.367
R1237 B.n532 B.n181 163.367
R1238 B.n533 B.n532 163.367
R1239 B.n534 B.n533 163.367
R1240 B.n534 B.n179 163.367
R1241 B.n538 B.n179 163.367
R1242 B.n540 B.n539 163.367
R1243 B.n540 B.n177 163.367
R1244 B.n544 B.n177 163.367
R1245 B.n545 B.n544 163.367
R1246 B.n546 B.n545 163.367
R1247 B.n546 B.n175 163.367
R1248 B.n550 B.n175 163.367
R1249 B.n551 B.n550 163.367
R1250 B.n552 B.n551 163.367
R1251 B.n552 B.n173 163.367
R1252 B.n556 B.n173 163.367
R1253 B.n557 B.n556 163.367
R1254 B.n558 B.n557 163.367
R1255 B.n558 B.n171 163.367
R1256 B.n562 B.n171 163.367
R1257 B.n563 B.n562 163.367
R1258 B.n564 B.n563 163.367
R1259 B.n564 B.n169 163.367
R1260 B.n568 B.n169 163.367
R1261 B.n569 B.n568 163.367
R1262 B.n570 B.n569 163.367
R1263 B.n570 B.n167 163.367
R1264 B.n574 B.n167 163.367
R1265 B.n575 B.n574 163.367
R1266 B.n576 B.n575 163.367
R1267 B.n576 B.n165 163.367
R1268 B.n580 B.n165 163.367
R1269 B.n581 B.n580 163.367
R1270 B.n582 B.n581 163.367
R1271 B.n582 B.n163 163.367
R1272 B.n586 B.n163 163.367
R1273 B.n587 B.n586 163.367
R1274 B.n588 B.n587 163.367
R1275 B.n588 B.n161 163.367
R1276 B.n592 B.n161 163.367
R1277 B.n593 B.n592 163.367
R1278 B.n594 B.n593 163.367
R1279 B.n594 B.n159 163.367
R1280 B.n598 B.n159 163.367
R1281 B.n599 B.n598 163.367
R1282 B.n600 B.n599 163.367
R1283 B.n600 B.n157 163.367
R1284 B.n604 B.n157 163.367
R1285 B.n605 B.n604 163.367
R1286 B.n606 B.n605 163.367
R1287 B.n606 B.n155 163.367
R1288 B.n610 B.n155 163.367
R1289 B.n611 B.n610 163.367
R1290 B.n612 B.n611 163.367
R1291 B.n612 B.n153 163.367
R1292 B.n616 B.n153 163.367
R1293 B.n617 B.n616 163.367
R1294 B.n618 B.n617 163.367
R1295 B.n618 B.n151 163.367
R1296 B.n622 B.n151 163.367
R1297 B.n623 B.n622 163.367
R1298 B.n624 B.n623 163.367
R1299 B.n624 B.n149 163.367
R1300 B.n628 B.n149 163.367
R1301 B.n629 B.n628 163.367
R1302 B.n630 B.n629 163.367
R1303 B.n630 B.n147 163.367
R1304 B.n634 B.n147 163.367
R1305 B.n635 B.n634 163.367
R1306 B.n636 B.n635 163.367
R1307 B.n636 B.n145 163.367
R1308 B.n640 B.n145 163.367
R1309 B.n641 B.n640 163.367
R1310 B.n642 B.n641 163.367
R1311 B.n642 B.n143 163.367
R1312 B.n646 B.n143 163.367
R1313 B.n647 B.n646 163.367
R1314 B.n648 B.n647 163.367
R1315 B.n648 B.n141 163.367
R1316 B.n652 B.n141 163.367
R1317 B.n653 B.n652 163.367
R1318 B.n654 B.n653 163.367
R1319 B.n654 B.n139 163.367
R1320 B.n658 B.n139 163.367
R1321 B.n659 B.n658 163.367
R1322 B.n660 B.n659 163.367
R1323 B.n660 B.n137 163.367
R1324 B.n664 B.n137 163.367
R1325 B.n665 B.n664 163.367
R1326 B.n666 B.n665 163.367
R1327 B.n666 B.n135 163.367
R1328 B.n670 B.n135 163.367
R1329 B.n671 B.n670 163.367
R1330 B.n672 B.n671 163.367
R1331 B.n672 B.n133 163.367
R1332 B.n676 B.n133 163.367
R1333 B.n677 B.n676 163.367
R1334 B.n678 B.n677 163.367
R1335 B.n678 B.n131 163.367
R1336 B.n682 B.n131 163.367
R1337 B.n683 B.n682 163.367
R1338 B.n684 B.n683 163.367
R1339 B.n684 B.n129 163.367
R1340 B.n688 B.n129 163.367
R1341 B.n689 B.n688 163.367
R1342 B.n690 B.n689 163.367
R1343 B.n690 B.n127 163.367
R1344 B.n694 B.n127 163.367
R1345 B.n695 B.n694 163.367
R1346 B.n696 B.n695 163.367
R1347 B.n696 B.n125 163.367
R1348 B.n700 B.n125 163.367
R1349 B.n701 B.n700 163.367
R1350 B.n702 B.n701 163.367
R1351 B.n702 B.n123 163.367
R1352 B.n706 B.n123 163.367
R1353 B.n707 B.n706 163.367
R1354 B.n708 B.n707 163.367
R1355 B.n708 B.n121 163.367
R1356 B.n712 B.n121 163.367
R1357 B.n713 B.n712 163.367
R1358 B.n714 B.n713 163.367
R1359 B.n714 B.n119 163.367
R1360 B.n718 B.n119 163.367
R1361 B.n719 B.n718 163.367
R1362 B.n720 B.n719 163.367
R1363 B.n720 B.n117 163.367
R1364 B.n724 B.n117 163.367
R1365 B.n725 B.n724 163.367
R1366 B.n726 B.n725 163.367
R1367 B.n726 B.n115 163.367
R1368 B.n730 B.n115 163.367
R1369 B.n731 B.n730 163.367
R1370 B.n732 B.n731 163.367
R1371 B.n732 B.n113 163.367
R1372 B.n736 B.n113 163.367
R1373 B.n737 B.n736 163.367
R1374 B.n738 B.n737 163.367
R1375 B.n738 B.n111 163.367
R1376 B.n742 B.n111 163.367
R1377 B.n743 B.n742 163.367
R1378 B.n744 B.n743 163.367
R1379 B.n744 B.n109 163.367
R1380 B.n748 B.n109 163.367
R1381 B.n749 B.n748 163.367
R1382 B.n750 B.n749 163.367
R1383 B.n750 B.n107 163.367
R1384 B.n754 B.n107 163.367
R1385 B.n755 B.n754 163.367
R1386 B.n756 B.n755 163.367
R1387 B.n756 B.n105 163.367
R1388 B.n760 B.n105 163.367
R1389 B.n761 B.n760 163.367
R1390 B.n762 B.n761 163.367
R1391 B.n762 B.n103 163.367
R1392 B.n766 B.n103 163.367
R1393 B.n767 B.n766 163.367
R1394 B.n768 B.n767 163.367
R1395 B.n768 B.n101 163.367
R1396 B.n772 B.n101 163.367
R1397 B.n773 B.n772 163.367
R1398 B.n774 B.n773 163.367
R1399 B.n774 B.n99 163.367
R1400 B.n778 B.n99 163.367
R1401 B.n779 B.n778 163.367
R1402 B.n780 B.n779 163.367
R1403 B.n780 B.n97 163.367
R1404 B.n784 B.n97 163.367
R1405 B.n785 B.n784 163.367
R1406 B.n786 B.n785 163.367
R1407 B.n786 B.n95 163.367
R1408 B.n932 B.n931 163.367
R1409 B.n931 B.n930 163.367
R1410 B.n930 B.n45 163.367
R1411 B.n926 B.n45 163.367
R1412 B.n926 B.n925 163.367
R1413 B.n925 B.n924 163.367
R1414 B.n924 B.n47 163.367
R1415 B.n920 B.n47 163.367
R1416 B.n920 B.n919 163.367
R1417 B.n919 B.n918 163.367
R1418 B.n918 B.n49 163.367
R1419 B.n914 B.n49 163.367
R1420 B.n914 B.n913 163.367
R1421 B.n913 B.n912 163.367
R1422 B.n912 B.n51 163.367
R1423 B.n908 B.n51 163.367
R1424 B.n908 B.n907 163.367
R1425 B.n907 B.n906 163.367
R1426 B.n906 B.n53 163.367
R1427 B.n902 B.n53 163.367
R1428 B.n902 B.n901 163.367
R1429 B.n901 B.n900 163.367
R1430 B.n900 B.n55 163.367
R1431 B.n896 B.n55 163.367
R1432 B.n896 B.n895 163.367
R1433 B.n895 B.n894 163.367
R1434 B.n894 B.n57 163.367
R1435 B.n890 B.n57 163.367
R1436 B.n890 B.n889 163.367
R1437 B.n889 B.n888 163.367
R1438 B.n888 B.n59 163.367
R1439 B.n884 B.n59 163.367
R1440 B.n884 B.n883 163.367
R1441 B.n883 B.n882 163.367
R1442 B.n882 B.n61 163.367
R1443 B.n878 B.n61 163.367
R1444 B.n878 B.n877 163.367
R1445 B.n877 B.n876 163.367
R1446 B.n876 B.n63 163.367
R1447 B.n872 B.n63 163.367
R1448 B.n872 B.n871 163.367
R1449 B.n871 B.n870 163.367
R1450 B.n870 B.n65 163.367
R1451 B.n865 B.n65 163.367
R1452 B.n865 B.n864 163.367
R1453 B.n864 B.n863 163.367
R1454 B.n863 B.n69 163.367
R1455 B.n859 B.n69 163.367
R1456 B.n859 B.n858 163.367
R1457 B.n858 B.n857 163.367
R1458 B.n857 B.n71 163.367
R1459 B.n852 B.n71 163.367
R1460 B.n852 B.n851 163.367
R1461 B.n851 B.n850 163.367
R1462 B.n850 B.n75 163.367
R1463 B.n846 B.n75 163.367
R1464 B.n846 B.n845 163.367
R1465 B.n845 B.n844 163.367
R1466 B.n844 B.n77 163.367
R1467 B.n840 B.n77 163.367
R1468 B.n840 B.n839 163.367
R1469 B.n839 B.n838 163.367
R1470 B.n838 B.n79 163.367
R1471 B.n834 B.n79 163.367
R1472 B.n834 B.n833 163.367
R1473 B.n833 B.n832 163.367
R1474 B.n832 B.n81 163.367
R1475 B.n828 B.n81 163.367
R1476 B.n828 B.n827 163.367
R1477 B.n827 B.n826 163.367
R1478 B.n826 B.n83 163.367
R1479 B.n822 B.n83 163.367
R1480 B.n822 B.n821 163.367
R1481 B.n821 B.n820 163.367
R1482 B.n820 B.n85 163.367
R1483 B.n816 B.n85 163.367
R1484 B.n816 B.n815 163.367
R1485 B.n815 B.n814 163.367
R1486 B.n814 B.n87 163.367
R1487 B.n810 B.n87 163.367
R1488 B.n810 B.n809 163.367
R1489 B.n809 B.n808 163.367
R1490 B.n808 B.n89 163.367
R1491 B.n804 B.n89 163.367
R1492 B.n804 B.n803 163.367
R1493 B.n803 B.n802 163.367
R1494 B.n802 B.n91 163.367
R1495 B.n798 B.n91 163.367
R1496 B.n798 B.n797 163.367
R1497 B.n797 B.n796 163.367
R1498 B.n796 B.n93 163.367
R1499 B.n792 B.n93 163.367
R1500 B.n792 B.n791 163.367
R1501 B.n791 B.n790 163.367
R1502 B.n201 B.t10 109.736
R1503 B.n73 B.t2 109.736
R1504 B.n209 B.t7 109.721
R1505 B.n67 B.t5 109.721
R1506 B.n201 B.n200 82.4247
R1507 B.n209 B.n208 82.4247
R1508 B.n67 B.n66 82.4247
R1509 B.n73 B.n72 82.4247
R1510 B.n202 B.n201 59.5399
R1511 B.n459 B.n209 59.5399
R1512 B.n868 B.n67 59.5399
R1513 B.n854 B.n73 59.5399
R1514 B.n934 B.n933 33.8737
R1515 B.n789 B.n788 33.8737
R1516 B.n537 B.n178 33.8737
R1517 B.n393 B.n230 33.8737
R1518 B B.n1059 18.0485
R1519 B.n933 B.n44 10.6151
R1520 B.n929 B.n44 10.6151
R1521 B.n929 B.n928 10.6151
R1522 B.n928 B.n927 10.6151
R1523 B.n927 B.n46 10.6151
R1524 B.n923 B.n46 10.6151
R1525 B.n923 B.n922 10.6151
R1526 B.n922 B.n921 10.6151
R1527 B.n921 B.n48 10.6151
R1528 B.n917 B.n48 10.6151
R1529 B.n917 B.n916 10.6151
R1530 B.n916 B.n915 10.6151
R1531 B.n915 B.n50 10.6151
R1532 B.n911 B.n50 10.6151
R1533 B.n911 B.n910 10.6151
R1534 B.n910 B.n909 10.6151
R1535 B.n909 B.n52 10.6151
R1536 B.n905 B.n52 10.6151
R1537 B.n905 B.n904 10.6151
R1538 B.n904 B.n903 10.6151
R1539 B.n903 B.n54 10.6151
R1540 B.n899 B.n54 10.6151
R1541 B.n899 B.n898 10.6151
R1542 B.n898 B.n897 10.6151
R1543 B.n897 B.n56 10.6151
R1544 B.n893 B.n56 10.6151
R1545 B.n893 B.n892 10.6151
R1546 B.n892 B.n891 10.6151
R1547 B.n891 B.n58 10.6151
R1548 B.n887 B.n58 10.6151
R1549 B.n887 B.n886 10.6151
R1550 B.n886 B.n885 10.6151
R1551 B.n885 B.n60 10.6151
R1552 B.n881 B.n60 10.6151
R1553 B.n881 B.n880 10.6151
R1554 B.n880 B.n879 10.6151
R1555 B.n879 B.n62 10.6151
R1556 B.n875 B.n62 10.6151
R1557 B.n875 B.n874 10.6151
R1558 B.n874 B.n873 10.6151
R1559 B.n873 B.n64 10.6151
R1560 B.n869 B.n64 10.6151
R1561 B.n867 B.n866 10.6151
R1562 B.n866 B.n68 10.6151
R1563 B.n862 B.n68 10.6151
R1564 B.n862 B.n861 10.6151
R1565 B.n861 B.n860 10.6151
R1566 B.n860 B.n70 10.6151
R1567 B.n856 B.n70 10.6151
R1568 B.n856 B.n855 10.6151
R1569 B.n853 B.n74 10.6151
R1570 B.n849 B.n74 10.6151
R1571 B.n849 B.n848 10.6151
R1572 B.n848 B.n847 10.6151
R1573 B.n847 B.n76 10.6151
R1574 B.n843 B.n76 10.6151
R1575 B.n843 B.n842 10.6151
R1576 B.n842 B.n841 10.6151
R1577 B.n841 B.n78 10.6151
R1578 B.n837 B.n78 10.6151
R1579 B.n837 B.n836 10.6151
R1580 B.n836 B.n835 10.6151
R1581 B.n835 B.n80 10.6151
R1582 B.n831 B.n80 10.6151
R1583 B.n831 B.n830 10.6151
R1584 B.n830 B.n829 10.6151
R1585 B.n829 B.n82 10.6151
R1586 B.n825 B.n82 10.6151
R1587 B.n825 B.n824 10.6151
R1588 B.n824 B.n823 10.6151
R1589 B.n823 B.n84 10.6151
R1590 B.n819 B.n84 10.6151
R1591 B.n819 B.n818 10.6151
R1592 B.n818 B.n817 10.6151
R1593 B.n817 B.n86 10.6151
R1594 B.n813 B.n86 10.6151
R1595 B.n813 B.n812 10.6151
R1596 B.n812 B.n811 10.6151
R1597 B.n811 B.n88 10.6151
R1598 B.n807 B.n88 10.6151
R1599 B.n807 B.n806 10.6151
R1600 B.n806 B.n805 10.6151
R1601 B.n805 B.n90 10.6151
R1602 B.n801 B.n90 10.6151
R1603 B.n801 B.n800 10.6151
R1604 B.n800 B.n799 10.6151
R1605 B.n799 B.n92 10.6151
R1606 B.n795 B.n92 10.6151
R1607 B.n795 B.n794 10.6151
R1608 B.n794 B.n793 10.6151
R1609 B.n793 B.n94 10.6151
R1610 B.n789 B.n94 10.6151
R1611 B.n541 B.n178 10.6151
R1612 B.n542 B.n541 10.6151
R1613 B.n543 B.n542 10.6151
R1614 B.n543 B.n176 10.6151
R1615 B.n547 B.n176 10.6151
R1616 B.n548 B.n547 10.6151
R1617 B.n549 B.n548 10.6151
R1618 B.n549 B.n174 10.6151
R1619 B.n553 B.n174 10.6151
R1620 B.n554 B.n553 10.6151
R1621 B.n555 B.n554 10.6151
R1622 B.n555 B.n172 10.6151
R1623 B.n559 B.n172 10.6151
R1624 B.n560 B.n559 10.6151
R1625 B.n561 B.n560 10.6151
R1626 B.n561 B.n170 10.6151
R1627 B.n565 B.n170 10.6151
R1628 B.n566 B.n565 10.6151
R1629 B.n567 B.n566 10.6151
R1630 B.n567 B.n168 10.6151
R1631 B.n571 B.n168 10.6151
R1632 B.n572 B.n571 10.6151
R1633 B.n573 B.n572 10.6151
R1634 B.n573 B.n166 10.6151
R1635 B.n577 B.n166 10.6151
R1636 B.n578 B.n577 10.6151
R1637 B.n579 B.n578 10.6151
R1638 B.n579 B.n164 10.6151
R1639 B.n583 B.n164 10.6151
R1640 B.n584 B.n583 10.6151
R1641 B.n585 B.n584 10.6151
R1642 B.n585 B.n162 10.6151
R1643 B.n589 B.n162 10.6151
R1644 B.n590 B.n589 10.6151
R1645 B.n591 B.n590 10.6151
R1646 B.n591 B.n160 10.6151
R1647 B.n595 B.n160 10.6151
R1648 B.n596 B.n595 10.6151
R1649 B.n597 B.n596 10.6151
R1650 B.n597 B.n158 10.6151
R1651 B.n601 B.n158 10.6151
R1652 B.n602 B.n601 10.6151
R1653 B.n603 B.n602 10.6151
R1654 B.n603 B.n156 10.6151
R1655 B.n607 B.n156 10.6151
R1656 B.n608 B.n607 10.6151
R1657 B.n609 B.n608 10.6151
R1658 B.n609 B.n154 10.6151
R1659 B.n613 B.n154 10.6151
R1660 B.n614 B.n613 10.6151
R1661 B.n615 B.n614 10.6151
R1662 B.n615 B.n152 10.6151
R1663 B.n619 B.n152 10.6151
R1664 B.n620 B.n619 10.6151
R1665 B.n621 B.n620 10.6151
R1666 B.n621 B.n150 10.6151
R1667 B.n625 B.n150 10.6151
R1668 B.n626 B.n625 10.6151
R1669 B.n627 B.n626 10.6151
R1670 B.n627 B.n148 10.6151
R1671 B.n631 B.n148 10.6151
R1672 B.n632 B.n631 10.6151
R1673 B.n633 B.n632 10.6151
R1674 B.n633 B.n146 10.6151
R1675 B.n637 B.n146 10.6151
R1676 B.n638 B.n637 10.6151
R1677 B.n639 B.n638 10.6151
R1678 B.n639 B.n144 10.6151
R1679 B.n643 B.n144 10.6151
R1680 B.n644 B.n643 10.6151
R1681 B.n645 B.n644 10.6151
R1682 B.n645 B.n142 10.6151
R1683 B.n649 B.n142 10.6151
R1684 B.n650 B.n649 10.6151
R1685 B.n651 B.n650 10.6151
R1686 B.n651 B.n140 10.6151
R1687 B.n655 B.n140 10.6151
R1688 B.n656 B.n655 10.6151
R1689 B.n657 B.n656 10.6151
R1690 B.n657 B.n138 10.6151
R1691 B.n661 B.n138 10.6151
R1692 B.n662 B.n661 10.6151
R1693 B.n663 B.n662 10.6151
R1694 B.n663 B.n136 10.6151
R1695 B.n667 B.n136 10.6151
R1696 B.n668 B.n667 10.6151
R1697 B.n669 B.n668 10.6151
R1698 B.n669 B.n134 10.6151
R1699 B.n673 B.n134 10.6151
R1700 B.n674 B.n673 10.6151
R1701 B.n675 B.n674 10.6151
R1702 B.n675 B.n132 10.6151
R1703 B.n679 B.n132 10.6151
R1704 B.n680 B.n679 10.6151
R1705 B.n681 B.n680 10.6151
R1706 B.n681 B.n130 10.6151
R1707 B.n685 B.n130 10.6151
R1708 B.n686 B.n685 10.6151
R1709 B.n687 B.n686 10.6151
R1710 B.n687 B.n128 10.6151
R1711 B.n691 B.n128 10.6151
R1712 B.n692 B.n691 10.6151
R1713 B.n693 B.n692 10.6151
R1714 B.n693 B.n126 10.6151
R1715 B.n697 B.n126 10.6151
R1716 B.n698 B.n697 10.6151
R1717 B.n699 B.n698 10.6151
R1718 B.n699 B.n124 10.6151
R1719 B.n703 B.n124 10.6151
R1720 B.n704 B.n703 10.6151
R1721 B.n705 B.n704 10.6151
R1722 B.n705 B.n122 10.6151
R1723 B.n709 B.n122 10.6151
R1724 B.n710 B.n709 10.6151
R1725 B.n711 B.n710 10.6151
R1726 B.n711 B.n120 10.6151
R1727 B.n715 B.n120 10.6151
R1728 B.n716 B.n715 10.6151
R1729 B.n717 B.n716 10.6151
R1730 B.n717 B.n118 10.6151
R1731 B.n721 B.n118 10.6151
R1732 B.n722 B.n721 10.6151
R1733 B.n723 B.n722 10.6151
R1734 B.n723 B.n116 10.6151
R1735 B.n727 B.n116 10.6151
R1736 B.n728 B.n727 10.6151
R1737 B.n729 B.n728 10.6151
R1738 B.n729 B.n114 10.6151
R1739 B.n733 B.n114 10.6151
R1740 B.n734 B.n733 10.6151
R1741 B.n735 B.n734 10.6151
R1742 B.n735 B.n112 10.6151
R1743 B.n739 B.n112 10.6151
R1744 B.n740 B.n739 10.6151
R1745 B.n741 B.n740 10.6151
R1746 B.n741 B.n110 10.6151
R1747 B.n745 B.n110 10.6151
R1748 B.n746 B.n745 10.6151
R1749 B.n747 B.n746 10.6151
R1750 B.n747 B.n108 10.6151
R1751 B.n751 B.n108 10.6151
R1752 B.n752 B.n751 10.6151
R1753 B.n753 B.n752 10.6151
R1754 B.n753 B.n106 10.6151
R1755 B.n757 B.n106 10.6151
R1756 B.n758 B.n757 10.6151
R1757 B.n759 B.n758 10.6151
R1758 B.n759 B.n104 10.6151
R1759 B.n763 B.n104 10.6151
R1760 B.n764 B.n763 10.6151
R1761 B.n765 B.n764 10.6151
R1762 B.n765 B.n102 10.6151
R1763 B.n769 B.n102 10.6151
R1764 B.n770 B.n769 10.6151
R1765 B.n771 B.n770 10.6151
R1766 B.n771 B.n100 10.6151
R1767 B.n775 B.n100 10.6151
R1768 B.n776 B.n775 10.6151
R1769 B.n777 B.n776 10.6151
R1770 B.n777 B.n98 10.6151
R1771 B.n781 B.n98 10.6151
R1772 B.n782 B.n781 10.6151
R1773 B.n783 B.n782 10.6151
R1774 B.n783 B.n96 10.6151
R1775 B.n787 B.n96 10.6151
R1776 B.n788 B.n787 10.6151
R1777 B.n397 B.n230 10.6151
R1778 B.n398 B.n397 10.6151
R1779 B.n399 B.n398 10.6151
R1780 B.n399 B.n228 10.6151
R1781 B.n403 B.n228 10.6151
R1782 B.n404 B.n403 10.6151
R1783 B.n405 B.n404 10.6151
R1784 B.n405 B.n226 10.6151
R1785 B.n409 B.n226 10.6151
R1786 B.n410 B.n409 10.6151
R1787 B.n411 B.n410 10.6151
R1788 B.n411 B.n224 10.6151
R1789 B.n415 B.n224 10.6151
R1790 B.n416 B.n415 10.6151
R1791 B.n417 B.n416 10.6151
R1792 B.n417 B.n222 10.6151
R1793 B.n421 B.n222 10.6151
R1794 B.n422 B.n421 10.6151
R1795 B.n423 B.n422 10.6151
R1796 B.n423 B.n220 10.6151
R1797 B.n427 B.n220 10.6151
R1798 B.n428 B.n427 10.6151
R1799 B.n429 B.n428 10.6151
R1800 B.n429 B.n218 10.6151
R1801 B.n433 B.n218 10.6151
R1802 B.n434 B.n433 10.6151
R1803 B.n435 B.n434 10.6151
R1804 B.n435 B.n216 10.6151
R1805 B.n439 B.n216 10.6151
R1806 B.n440 B.n439 10.6151
R1807 B.n441 B.n440 10.6151
R1808 B.n441 B.n214 10.6151
R1809 B.n445 B.n214 10.6151
R1810 B.n446 B.n445 10.6151
R1811 B.n447 B.n446 10.6151
R1812 B.n447 B.n212 10.6151
R1813 B.n451 B.n212 10.6151
R1814 B.n452 B.n451 10.6151
R1815 B.n453 B.n452 10.6151
R1816 B.n453 B.n210 10.6151
R1817 B.n457 B.n210 10.6151
R1818 B.n458 B.n457 10.6151
R1819 B.n460 B.n206 10.6151
R1820 B.n464 B.n206 10.6151
R1821 B.n465 B.n464 10.6151
R1822 B.n466 B.n465 10.6151
R1823 B.n466 B.n204 10.6151
R1824 B.n470 B.n204 10.6151
R1825 B.n471 B.n470 10.6151
R1826 B.n472 B.n471 10.6151
R1827 B.n476 B.n475 10.6151
R1828 B.n477 B.n476 10.6151
R1829 B.n477 B.n198 10.6151
R1830 B.n481 B.n198 10.6151
R1831 B.n482 B.n481 10.6151
R1832 B.n483 B.n482 10.6151
R1833 B.n483 B.n196 10.6151
R1834 B.n487 B.n196 10.6151
R1835 B.n488 B.n487 10.6151
R1836 B.n489 B.n488 10.6151
R1837 B.n489 B.n194 10.6151
R1838 B.n493 B.n194 10.6151
R1839 B.n494 B.n493 10.6151
R1840 B.n495 B.n494 10.6151
R1841 B.n495 B.n192 10.6151
R1842 B.n499 B.n192 10.6151
R1843 B.n500 B.n499 10.6151
R1844 B.n501 B.n500 10.6151
R1845 B.n501 B.n190 10.6151
R1846 B.n505 B.n190 10.6151
R1847 B.n506 B.n505 10.6151
R1848 B.n507 B.n506 10.6151
R1849 B.n507 B.n188 10.6151
R1850 B.n511 B.n188 10.6151
R1851 B.n512 B.n511 10.6151
R1852 B.n513 B.n512 10.6151
R1853 B.n513 B.n186 10.6151
R1854 B.n517 B.n186 10.6151
R1855 B.n518 B.n517 10.6151
R1856 B.n519 B.n518 10.6151
R1857 B.n519 B.n184 10.6151
R1858 B.n523 B.n184 10.6151
R1859 B.n524 B.n523 10.6151
R1860 B.n525 B.n524 10.6151
R1861 B.n525 B.n182 10.6151
R1862 B.n529 B.n182 10.6151
R1863 B.n530 B.n529 10.6151
R1864 B.n531 B.n530 10.6151
R1865 B.n531 B.n180 10.6151
R1866 B.n535 B.n180 10.6151
R1867 B.n536 B.n535 10.6151
R1868 B.n537 B.n536 10.6151
R1869 B.n393 B.n392 10.6151
R1870 B.n392 B.n391 10.6151
R1871 B.n391 B.n232 10.6151
R1872 B.n387 B.n232 10.6151
R1873 B.n387 B.n386 10.6151
R1874 B.n386 B.n385 10.6151
R1875 B.n385 B.n234 10.6151
R1876 B.n381 B.n234 10.6151
R1877 B.n381 B.n380 10.6151
R1878 B.n380 B.n379 10.6151
R1879 B.n379 B.n236 10.6151
R1880 B.n375 B.n236 10.6151
R1881 B.n375 B.n374 10.6151
R1882 B.n374 B.n373 10.6151
R1883 B.n373 B.n238 10.6151
R1884 B.n369 B.n238 10.6151
R1885 B.n369 B.n368 10.6151
R1886 B.n368 B.n367 10.6151
R1887 B.n367 B.n240 10.6151
R1888 B.n363 B.n240 10.6151
R1889 B.n363 B.n362 10.6151
R1890 B.n362 B.n361 10.6151
R1891 B.n361 B.n242 10.6151
R1892 B.n357 B.n242 10.6151
R1893 B.n357 B.n356 10.6151
R1894 B.n356 B.n355 10.6151
R1895 B.n355 B.n244 10.6151
R1896 B.n351 B.n244 10.6151
R1897 B.n351 B.n350 10.6151
R1898 B.n350 B.n349 10.6151
R1899 B.n349 B.n246 10.6151
R1900 B.n345 B.n246 10.6151
R1901 B.n345 B.n344 10.6151
R1902 B.n344 B.n343 10.6151
R1903 B.n343 B.n248 10.6151
R1904 B.n339 B.n248 10.6151
R1905 B.n339 B.n338 10.6151
R1906 B.n338 B.n337 10.6151
R1907 B.n337 B.n250 10.6151
R1908 B.n333 B.n250 10.6151
R1909 B.n333 B.n332 10.6151
R1910 B.n332 B.n331 10.6151
R1911 B.n331 B.n252 10.6151
R1912 B.n327 B.n252 10.6151
R1913 B.n327 B.n326 10.6151
R1914 B.n326 B.n325 10.6151
R1915 B.n325 B.n254 10.6151
R1916 B.n321 B.n254 10.6151
R1917 B.n321 B.n320 10.6151
R1918 B.n320 B.n319 10.6151
R1919 B.n319 B.n256 10.6151
R1920 B.n315 B.n256 10.6151
R1921 B.n315 B.n314 10.6151
R1922 B.n314 B.n313 10.6151
R1923 B.n313 B.n258 10.6151
R1924 B.n309 B.n258 10.6151
R1925 B.n309 B.n308 10.6151
R1926 B.n308 B.n307 10.6151
R1927 B.n307 B.n260 10.6151
R1928 B.n303 B.n260 10.6151
R1929 B.n303 B.n302 10.6151
R1930 B.n302 B.n301 10.6151
R1931 B.n301 B.n262 10.6151
R1932 B.n297 B.n262 10.6151
R1933 B.n297 B.n296 10.6151
R1934 B.n296 B.n295 10.6151
R1935 B.n295 B.n264 10.6151
R1936 B.n291 B.n264 10.6151
R1937 B.n291 B.n290 10.6151
R1938 B.n290 B.n289 10.6151
R1939 B.n289 B.n266 10.6151
R1940 B.n285 B.n266 10.6151
R1941 B.n285 B.n284 10.6151
R1942 B.n284 B.n283 10.6151
R1943 B.n283 B.n268 10.6151
R1944 B.n279 B.n268 10.6151
R1945 B.n279 B.n278 10.6151
R1946 B.n278 B.n277 10.6151
R1947 B.n277 B.n270 10.6151
R1948 B.n273 B.n270 10.6151
R1949 B.n273 B.n272 10.6151
R1950 B.n272 B.n0 10.6151
R1951 B.n1055 B.n1 10.6151
R1952 B.n1055 B.n1054 10.6151
R1953 B.n1054 B.n1053 10.6151
R1954 B.n1053 B.n4 10.6151
R1955 B.n1049 B.n4 10.6151
R1956 B.n1049 B.n1048 10.6151
R1957 B.n1048 B.n1047 10.6151
R1958 B.n1047 B.n6 10.6151
R1959 B.n1043 B.n6 10.6151
R1960 B.n1043 B.n1042 10.6151
R1961 B.n1042 B.n1041 10.6151
R1962 B.n1041 B.n8 10.6151
R1963 B.n1037 B.n8 10.6151
R1964 B.n1037 B.n1036 10.6151
R1965 B.n1036 B.n1035 10.6151
R1966 B.n1035 B.n10 10.6151
R1967 B.n1031 B.n10 10.6151
R1968 B.n1031 B.n1030 10.6151
R1969 B.n1030 B.n1029 10.6151
R1970 B.n1029 B.n12 10.6151
R1971 B.n1025 B.n12 10.6151
R1972 B.n1025 B.n1024 10.6151
R1973 B.n1024 B.n1023 10.6151
R1974 B.n1023 B.n14 10.6151
R1975 B.n1019 B.n14 10.6151
R1976 B.n1019 B.n1018 10.6151
R1977 B.n1018 B.n1017 10.6151
R1978 B.n1017 B.n16 10.6151
R1979 B.n1013 B.n16 10.6151
R1980 B.n1013 B.n1012 10.6151
R1981 B.n1012 B.n1011 10.6151
R1982 B.n1011 B.n18 10.6151
R1983 B.n1007 B.n18 10.6151
R1984 B.n1007 B.n1006 10.6151
R1985 B.n1006 B.n1005 10.6151
R1986 B.n1005 B.n20 10.6151
R1987 B.n1001 B.n20 10.6151
R1988 B.n1001 B.n1000 10.6151
R1989 B.n1000 B.n999 10.6151
R1990 B.n999 B.n22 10.6151
R1991 B.n995 B.n22 10.6151
R1992 B.n995 B.n994 10.6151
R1993 B.n994 B.n993 10.6151
R1994 B.n993 B.n24 10.6151
R1995 B.n989 B.n24 10.6151
R1996 B.n989 B.n988 10.6151
R1997 B.n988 B.n987 10.6151
R1998 B.n987 B.n26 10.6151
R1999 B.n983 B.n26 10.6151
R2000 B.n983 B.n982 10.6151
R2001 B.n982 B.n981 10.6151
R2002 B.n981 B.n28 10.6151
R2003 B.n977 B.n28 10.6151
R2004 B.n977 B.n976 10.6151
R2005 B.n976 B.n975 10.6151
R2006 B.n975 B.n30 10.6151
R2007 B.n971 B.n30 10.6151
R2008 B.n971 B.n970 10.6151
R2009 B.n970 B.n969 10.6151
R2010 B.n969 B.n32 10.6151
R2011 B.n965 B.n32 10.6151
R2012 B.n965 B.n964 10.6151
R2013 B.n964 B.n963 10.6151
R2014 B.n963 B.n34 10.6151
R2015 B.n959 B.n34 10.6151
R2016 B.n959 B.n958 10.6151
R2017 B.n958 B.n957 10.6151
R2018 B.n957 B.n36 10.6151
R2019 B.n953 B.n36 10.6151
R2020 B.n953 B.n952 10.6151
R2021 B.n952 B.n951 10.6151
R2022 B.n951 B.n38 10.6151
R2023 B.n947 B.n38 10.6151
R2024 B.n947 B.n946 10.6151
R2025 B.n946 B.n945 10.6151
R2026 B.n945 B.n40 10.6151
R2027 B.n941 B.n40 10.6151
R2028 B.n941 B.n940 10.6151
R2029 B.n940 B.n939 10.6151
R2030 B.n939 B.n42 10.6151
R2031 B.n935 B.n42 10.6151
R2032 B.n935 B.n934 10.6151
R2033 B.n868 B.n867 6.5566
R2034 B.n855 B.n854 6.5566
R2035 B.n460 B.n459 6.5566
R2036 B.n472 B.n202 6.5566
R2037 B.n869 B.n868 4.05904
R2038 B.n854 B.n853 4.05904
R2039 B.n459 B.n458 4.05904
R2040 B.n475 B.n202 4.05904
R2041 B.n1059 B.n0 2.81026
R2042 B.n1059 B.n1 2.81026
C0 w_n6070_n3444# VN 13.408599f
C1 VP w_n6070_n3444# 14.2029f
C2 VDD2 VDD1 3.03467f
C3 VDD2 VN 11.765201f
C4 VTAIL VDD1 11.2472f
C5 VP VDD2 0.751043f
C6 VTAIL VN 12.9545f
C7 B w_n6070_n3444# 12.8724f
C8 VTAIL VP 12.9695f
C9 VDD1 VN 0.156068f
C10 VDD2 B 3.19218f
C11 VP VDD1 12.356701f
C12 VTAIL B 4.31387f
C13 VDD2 w_n6070_n3444# 3.52436f
C14 VP VN 10.425301f
C15 VTAIL w_n6070_n3444# 3.45168f
C16 VDD1 B 3.02286f
C17 B VN 1.61869f
C18 VDD1 w_n6070_n3444# 3.3122f
C19 VTAIL VDD2 11.3079f
C20 VP B 2.96173f
C21 VDD2 VSUBS 2.69327f
C22 VDD1 VSUBS 2.533946f
C23 VTAIL VSUBS 1.6334f
C24 VN VSUBS 9.9472f
C25 VP VSUBS 5.954547f
C26 B VSUBS 7.034169f
C27 w_n6070_n3444# VSUBS 0.257198p
C28 B.n0 VSUBS 0.005491f
C29 B.n1 VSUBS 0.005491f
C30 B.n2 VSUBS 0.008683f
C31 B.n3 VSUBS 0.008683f
C32 B.n4 VSUBS 0.008683f
C33 B.n5 VSUBS 0.008683f
C34 B.n6 VSUBS 0.008683f
C35 B.n7 VSUBS 0.008683f
C36 B.n8 VSUBS 0.008683f
C37 B.n9 VSUBS 0.008683f
C38 B.n10 VSUBS 0.008683f
C39 B.n11 VSUBS 0.008683f
C40 B.n12 VSUBS 0.008683f
C41 B.n13 VSUBS 0.008683f
C42 B.n14 VSUBS 0.008683f
C43 B.n15 VSUBS 0.008683f
C44 B.n16 VSUBS 0.008683f
C45 B.n17 VSUBS 0.008683f
C46 B.n18 VSUBS 0.008683f
C47 B.n19 VSUBS 0.008683f
C48 B.n20 VSUBS 0.008683f
C49 B.n21 VSUBS 0.008683f
C50 B.n22 VSUBS 0.008683f
C51 B.n23 VSUBS 0.008683f
C52 B.n24 VSUBS 0.008683f
C53 B.n25 VSUBS 0.008683f
C54 B.n26 VSUBS 0.008683f
C55 B.n27 VSUBS 0.008683f
C56 B.n28 VSUBS 0.008683f
C57 B.n29 VSUBS 0.008683f
C58 B.n30 VSUBS 0.008683f
C59 B.n31 VSUBS 0.008683f
C60 B.n32 VSUBS 0.008683f
C61 B.n33 VSUBS 0.008683f
C62 B.n34 VSUBS 0.008683f
C63 B.n35 VSUBS 0.008683f
C64 B.n36 VSUBS 0.008683f
C65 B.n37 VSUBS 0.008683f
C66 B.n38 VSUBS 0.008683f
C67 B.n39 VSUBS 0.008683f
C68 B.n40 VSUBS 0.008683f
C69 B.n41 VSUBS 0.008683f
C70 B.n42 VSUBS 0.008683f
C71 B.n43 VSUBS 0.020271f
C72 B.n44 VSUBS 0.008683f
C73 B.n45 VSUBS 0.008683f
C74 B.n46 VSUBS 0.008683f
C75 B.n47 VSUBS 0.008683f
C76 B.n48 VSUBS 0.008683f
C77 B.n49 VSUBS 0.008683f
C78 B.n50 VSUBS 0.008683f
C79 B.n51 VSUBS 0.008683f
C80 B.n52 VSUBS 0.008683f
C81 B.n53 VSUBS 0.008683f
C82 B.n54 VSUBS 0.008683f
C83 B.n55 VSUBS 0.008683f
C84 B.n56 VSUBS 0.008683f
C85 B.n57 VSUBS 0.008683f
C86 B.n58 VSUBS 0.008683f
C87 B.n59 VSUBS 0.008683f
C88 B.n60 VSUBS 0.008683f
C89 B.n61 VSUBS 0.008683f
C90 B.n62 VSUBS 0.008683f
C91 B.n63 VSUBS 0.008683f
C92 B.n64 VSUBS 0.008683f
C93 B.n65 VSUBS 0.008683f
C94 B.t5 VSUBS 0.502099f
C95 B.t4 VSUBS 0.537912f
C96 B.t3 VSUBS 2.80786f
C97 B.n66 VSUBS 0.31311f
C98 B.n67 VSUBS 0.095871f
C99 B.n68 VSUBS 0.008683f
C100 B.n69 VSUBS 0.008683f
C101 B.n70 VSUBS 0.008683f
C102 B.n71 VSUBS 0.008683f
C103 B.t2 VSUBS 0.502089f
C104 B.t1 VSUBS 0.537904f
C105 B.t0 VSUBS 2.80786f
C106 B.n72 VSUBS 0.313119f
C107 B.n73 VSUBS 0.095881f
C108 B.n74 VSUBS 0.008683f
C109 B.n75 VSUBS 0.008683f
C110 B.n76 VSUBS 0.008683f
C111 B.n77 VSUBS 0.008683f
C112 B.n78 VSUBS 0.008683f
C113 B.n79 VSUBS 0.008683f
C114 B.n80 VSUBS 0.008683f
C115 B.n81 VSUBS 0.008683f
C116 B.n82 VSUBS 0.008683f
C117 B.n83 VSUBS 0.008683f
C118 B.n84 VSUBS 0.008683f
C119 B.n85 VSUBS 0.008683f
C120 B.n86 VSUBS 0.008683f
C121 B.n87 VSUBS 0.008683f
C122 B.n88 VSUBS 0.008683f
C123 B.n89 VSUBS 0.008683f
C124 B.n90 VSUBS 0.008683f
C125 B.n91 VSUBS 0.008683f
C126 B.n92 VSUBS 0.008683f
C127 B.n93 VSUBS 0.008683f
C128 B.n94 VSUBS 0.008683f
C129 B.n95 VSUBS 0.020271f
C130 B.n96 VSUBS 0.008683f
C131 B.n97 VSUBS 0.008683f
C132 B.n98 VSUBS 0.008683f
C133 B.n99 VSUBS 0.008683f
C134 B.n100 VSUBS 0.008683f
C135 B.n101 VSUBS 0.008683f
C136 B.n102 VSUBS 0.008683f
C137 B.n103 VSUBS 0.008683f
C138 B.n104 VSUBS 0.008683f
C139 B.n105 VSUBS 0.008683f
C140 B.n106 VSUBS 0.008683f
C141 B.n107 VSUBS 0.008683f
C142 B.n108 VSUBS 0.008683f
C143 B.n109 VSUBS 0.008683f
C144 B.n110 VSUBS 0.008683f
C145 B.n111 VSUBS 0.008683f
C146 B.n112 VSUBS 0.008683f
C147 B.n113 VSUBS 0.008683f
C148 B.n114 VSUBS 0.008683f
C149 B.n115 VSUBS 0.008683f
C150 B.n116 VSUBS 0.008683f
C151 B.n117 VSUBS 0.008683f
C152 B.n118 VSUBS 0.008683f
C153 B.n119 VSUBS 0.008683f
C154 B.n120 VSUBS 0.008683f
C155 B.n121 VSUBS 0.008683f
C156 B.n122 VSUBS 0.008683f
C157 B.n123 VSUBS 0.008683f
C158 B.n124 VSUBS 0.008683f
C159 B.n125 VSUBS 0.008683f
C160 B.n126 VSUBS 0.008683f
C161 B.n127 VSUBS 0.008683f
C162 B.n128 VSUBS 0.008683f
C163 B.n129 VSUBS 0.008683f
C164 B.n130 VSUBS 0.008683f
C165 B.n131 VSUBS 0.008683f
C166 B.n132 VSUBS 0.008683f
C167 B.n133 VSUBS 0.008683f
C168 B.n134 VSUBS 0.008683f
C169 B.n135 VSUBS 0.008683f
C170 B.n136 VSUBS 0.008683f
C171 B.n137 VSUBS 0.008683f
C172 B.n138 VSUBS 0.008683f
C173 B.n139 VSUBS 0.008683f
C174 B.n140 VSUBS 0.008683f
C175 B.n141 VSUBS 0.008683f
C176 B.n142 VSUBS 0.008683f
C177 B.n143 VSUBS 0.008683f
C178 B.n144 VSUBS 0.008683f
C179 B.n145 VSUBS 0.008683f
C180 B.n146 VSUBS 0.008683f
C181 B.n147 VSUBS 0.008683f
C182 B.n148 VSUBS 0.008683f
C183 B.n149 VSUBS 0.008683f
C184 B.n150 VSUBS 0.008683f
C185 B.n151 VSUBS 0.008683f
C186 B.n152 VSUBS 0.008683f
C187 B.n153 VSUBS 0.008683f
C188 B.n154 VSUBS 0.008683f
C189 B.n155 VSUBS 0.008683f
C190 B.n156 VSUBS 0.008683f
C191 B.n157 VSUBS 0.008683f
C192 B.n158 VSUBS 0.008683f
C193 B.n159 VSUBS 0.008683f
C194 B.n160 VSUBS 0.008683f
C195 B.n161 VSUBS 0.008683f
C196 B.n162 VSUBS 0.008683f
C197 B.n163 VSUBS 0.008683f
C198 B.n164 VSUBS 0.008683f
C199 B.n165 VSUBS 0.008683f
C200 B.n166 VSUBS 0.008683f
C201 B.n167 VSUBS 0.008683f
C202 B.n168 VSUBS 0.008683f
C203 B.n169 VSUBS 0.008683f
C204 B.n170 VSUBS 0.008683f
C205 B.n171 VSUBS 0.008683f
C206 B.n172 VSUBS 0.008683f
C207 B.n173 VSUBS 0.008683f
C208 B.n174 VSUBS 0.008683f
C209 B.n175 VSUBS 0.008683f
C210 B.n176 VSUBS 0.008683f
C211 B.n177 VSUBS 0.008683f
C212 B.n178 VSUBS 0.020271f
C213 B.n179 VSUBS 0.008683f
C214 B.n180 VSUBS 0.008683f
C215 B.n181 VSUBS 0.008683f
C216 B.n182 VSUBS 0.008683f
C217 B.n183 VSUBS 0.008683f
C218 B.n184 VSUBS 0.008683f
C219 B.n185 VSUBS 0.008683f
C220 B.n186 VSUBS 0.008683f
C221 B.n187 VSUBS 0.008683f
C222 B.n188 VSUBS 0.008683f
C223 B.n189 VSUBS 0.008683f
C224 B.n190 VSUBS 0.008683f
C225 B.n191 VSUBS 0.008683f
C226 B.n192 VSUBS 0.008683f
C227 B.n193 VSUBS 0.008683f
C228 B.n194 VSUBS 0.008683f
C229 B.n195 VSUBS 0.008683f
C230 B.n196 VSUBS 0.008683f
C231 B.n197 VSUBS 0.008683f
C232 B.n198 VSUBS 0.008683f
C233 B.n199 VSUBS 0.008683f
C234 B.t10 VSUBS 0.502089f
C235 B.t11 VSUBS 0.537904f
C236 B.t9 VSUBS 2.80786f
C237 B.n200 VSUBS 0.313119f
C238 B.n201 VSUBS 0.095881f
C239 B.n202 VSUBS 0.020118f
C240 B.n203 VSUBS 0.008683f
C241 B.n204 VSUBS 0.008683f
C242 B.n205 VSUBS 0.008683f
C243 B.n206 VSUBS 0.008683f
C244 B.n207 VSUBS 0.008683f
C245 B.t7 VSUBS 0.502099f
C246 B.t8 VSUBS 0.537912f
C247 B.t6 VSUBS 2.80786f
C248 B.n208 VSUBS 0.31311f
C249 B.n209 VSUBS 0.095871f
C250 B.n210 VSUBS 0.008683f
C251 B.n211 VSUBS 0.008683f
C252 B.n212 VSUBS 0.008683f
C253 B.n213 VSUBS 0.008683f
C254 B.n214 VSUBS 0.008683f
C255 B.n215 VSUBS 0.008683f
C256 B.n216 VSUBS 0.008683f
C257 B.n217 VSUBS 0.008683f
C258 B.n218 VSUBS 0.008683f
C259 B.n219 VSUBS 0.008683f
C260 B.n220 VSUBS 0.008683f
C261 B.n221 VSUBS 0.008683f
C262 B.n222 VSUBS 0.008683f
C263 B.n223 VSUBS 0.008683f
C264 B.n224 VSUBS 0.008683f
C265 B.n225 VSUBS 0.008683f
C266 B.n226 VSUBS 0.008683f
C267 B.n227 VSUBS 0.008683f
C268 B.n228 VSUBS 0.008683f
C269 B.n229 VSUBS 0.008683f
C270 B.n230 VSUBS 0.021357f
C271 B.n231 VSUBS 0.008683f
C272 B.n232 VSUBS 0.008683f
C273 B.n233 VSUBS 0.008683f
C274 B.n234 VSUBS 0.008683f
C275 B.n235 VSUBS 0.008683f
C276 B.n236 VSUBS 0.008683f
C277 B.n237 VSUBS 0.008683f
C278 B.n238 VSUBS 0.008683f
C279 B.n239 VSUBS 0.008683f
C280 B.n240 VSUBS 0.008683f
C281 B.n241 VSUBS 0.008683f
C282 B.n242 VSUBS 0.008683f
C283 B.n243 VSUBS 0.008683f
C284 B.n244 VSUBS 0.008683f
C285 B.n245 VSUBS 0.008683f
C286 B.n246 VSUBS 0.008683f
C287 B.n247 VSUBS 0.008683f
C288 B.n248 VSUBS 0.008683f
C289 B.n249 VSUBS 0.008683f
C290 B.n250 VSUBS 0.008683f
C291 B.n251 VSUBS 0.008683f
C292 B.n252 VSUBS 0.008683f
C293 B.n253 VSUBS 0.008683f
C294 B.n254 VSUBS 0.008683f
C295 B.n255 VSUBS 0.008683f
C296 B.n256 VSUBS 0.008683f
C297 B.n257 VSUBS 0.008683f
C298 B.n258 VSUBS 0.008683f
C299 B.n259 VSUBS 0.008683f
C300 B.n260 VSUBS 0.008683f
C301 B.n261 VSUBS 0.008683f
C302 B.n262 VSUBS 0.008683f
C303 B.n263 VSUBS 0.008683f
C304 B.n264 VSUBS 0.008683f
C305 B.n265 VSUBS 0.008683f
C306 B.n266 VSUBS 0.008683f
C307 B.n267 VSUBS 0.008683f
C308 B.n268 VSUBS 0.008683f
C309 B.n269 VSUBS 0.008683f
C310 B.n270 VSUBS 0.008683f
C311 B.n271 VSUBS 0.008683f
C312 B.n272 VSUBS 0.008683f
C313 B.n273 VSUBS 0.008683f
C314 B.n274 VSUBS 0.008683f
C315 B.n275 VSUBS 0.008683f
C316 B.n276 VSUBS 0.008683f
C317 B.n277 VSUBS 0.008683f
C318 B.n278 VSUBS 0.008683f
C319 B.n279 VSUBS 0.008683f
C320 B.n280 VSUBS 0.008683f
C321 B.n281 VSUBS 0.008683f
C322 B.n282 VSUBS 0.008683f
C323 B.n283 VSUBS 0.008683f
C324 B.n284 VSUBS 0.008683f
C325 B.n285 VSUBS 0.008683f
C326 B.n286 VSUBS 0.008683f
C327 B.n287 VSUBS 0.008683f
C328 B.n288 VSUBS 0.008683f
C329 B.n289 VSUBS 0.008683f
C330 B.n290 VSUBS 0.008683f
C331 B.n291 VSUBS 0.008683f
C332 B.n292 VSUBS 0.008683f
C333 B.n293 VSUBS 0.008683f
C334 B.n294 VSUBS 0.008683f
C335 B.n295 VSUBS 0.008683f
C336 B.n296 VSUBS 0.008683f
C337 B.n297 VSUBS 0.008683f
C338 B.n298 VSUBS 0.008683f
C339 B.n299 VSUBS 0.008683f
C340 B.n300 VSUBS 0.008683f
C341 B.n301 VSUBS 0.008683f
C342 B.n302 VSUBS 0.008683f
C343 B.n303 VSUBS 0.008683f
C344 B.n304 VSUBS 0.008683f
C345 B.n305 VSUBS 0.008683f
C346 B.n306 VSUBS 0.008683f
C347 B.n307 VSUBS 0.008683f
C348 B.n308 VSUBS 0.008683f
C349 B.n309 VSUBS 0.008683f
C350 B.n310 VSUBS 0.008683f
C351 B.n311 VSUBS 0.008683f
C352 B.n312 VSUBS 0.008683f
C353 B.n313 VSUBS 0.008683f
C354 B.n314 VSUBS 0.008683f
C355 B.n315 VSUBS 0.008683f
C356 B.n316 VSUBS 0.008683f
C357 B.n317 VSUBS 0.008683f
C358 B.n318 VSUBS 0.008683f
C359 B.n319 VSUBS 0.008683f
C360 B.n320 VSUBS 0.008683f
C361 B.n321 VSUBS 0.008683f
C362 B.n322 VSUBS 0.008683f
C363 B.n323 VSUBS 0.008683f
C364 B.n324 VSUBS 0.008683f
C365 B.n325 VSUBS 0.008683f
C366 B.n326 VSUBS 0.008683f
C367 B.n327 VSUBS 0.008683f
C368 B.n328 VSUBS 0.008683f
C369 B.n329 VSUBS 0.008683f
C370 B.n330 VSUBS 0.008683f
C371 B.n331 VSUBS 0.008683f
C372 B.n332 VSUBS 0.008683f
C373 B.n333 VSUBS 0.008683f
C374 B.n334 VSUBS 0.008683f
C375 B.n335 VSUBS 0.008683f
C376 B.n336 VSUBS 0.008683f
C377 B.n337 VSUBS 0.008683f
C378 B.n338 VSUBS 0.008683f
C379 B.n339 VSUBS 0.008683f
C380 B.n340 VSUBS 0.008683f
C381 B.n341 VSUBS 0.008683f
C382 B.n342 VSUBS 0.008683f
C383 B.n343 VSUBS 0.008683f
C384 B.n344 VSUBS 0.008683f
C385 B.n345 VSUBS 0.008683f
C386 B.n346 VSUBS 0.008683f
C387 B.n347 VSUBS 0.008683f
C388 B.n348 VSUBS 0.008683f
C389 B.n349 VSUBS 0.008683f
C390 B.n350 VSUBS 0.008683f
C391 B.n351 VSUBS 0.008683f
C392 B.n352 VSUBS 0.008683f
C393 B.n353 VSUBS 0.008683f
C394 B.n354 VSUBS 0.008683f
C395 B.n355 VSUBS 0.008683f
C396 B.n356 VSUBS 0.008683f
C397 B.n357 VSUBS 0.008683f
C398 B.n358 VSUBS 0.008683f
C399 B.n359 VSUBS 0.008683f
C400 B.n360 VSUBS 0.008683f
C401 B.n361 VSUBS 0.008683f
C402 B.n362 VSUBS 0.008683f
C403 B.n363 VSUBS 0.008683f
C404 B.n364 VSUBS 0.008683f
C405 B.n365 VSUBS 0.008683f
C406 B.n366 VSUBS 0.008683f
C407 B.n367 VSUBS 0.008683f
C408 B.n368 VSUBS 0.008683f
C409 B.n369 VSUBS 0.008683f
C410 B.n370 VSUBS 0.008683f
C411 B.n371 VSUBS 0.008683f
C412 B.n372 VSUBS 0.008683f
C413 B.n373 VSUBS 0.008683f
C414 B.n374 VSUBS 0.008683f
C415 B.n375 VSUBS 0.008683f
C416 B.n376 VSUBS 0.008683f
C417 B.n377 VSUBS 0.008683f
C418 B.n378 VSUBS 0.008683f
C419 B.n379 VSUBS 0.008683f
C420 B.n380 VSUBS 0.008683f
C421 B.n381 VSUBS 0.008683f
C422 B.n382 VSUBS 0.008683f
C423 B.n383 VSUBS 0.008683f
C424 B.n384 VSUBS 0.008683f
C425 B.n385 VSUBS 0.008683f
C426 B.n386 VSUBS 0.008683f
C427 B.n387 VSUBS 0.008683f
C428 B.n388 VSUBS 0.008683f
C429 B.n389 VSUBS 0.008683f
C430 B.n390 VSUBS 0.008683f
C431 B.n391 VSUBS 0.008683f
C432 B.n392 VSUBS 0.008683f
C433 B.n393 VSUBS 0.020271f
C434 B.n394 VSUBS 0.020271f
C435 B.n395 VSUBS 0.021357f
C436 B.n396 VSUBS 0.008683f
C437 B.n397 VSUBS 0.008683f
C438 B.n398 VSUBS 0.008683f
C439 B.n399 VSUBS 0.008683f
C440 B.n400 VSUBS 0.008683f
C441 B.n401 VSUBS 0.008683f
C442 B.n402 VSUBS 0.008683f
C443 B.n403 VSUBS 0.008683f
C444 B.n404 VSUBS 0.008683f
C445 B.n405 VSUBS 0.008683f
C446 B.n406 VSUBS 0.008683f
C447 B.n407 VSUBS 0.008683f
C448 B.n408 VSUBS 0.008683f
C449 B.n409 VSUBS 0.008683f
C450 B.n410 VSUBS 0.008683f
C451 B.n411 VSUBS 0.008683f
C452 B.n412 VSUBS 0.008683f
C453 B.n413 VSUBS 0.008683f
C454 B.n414 VSUBS 0.008683f
C455 B.n415 VSUBS 0.008683f
C456 B.n416 VSUBS 0.008683f
C457 B.n417 VSUBS 0.008683f
C458 B.n418 VSUBS 0.008683f
C459 B.n419 VSUBS 0.008683f
C460 B.n420 VSUBS 0.008683f
C461 B.n421 VSUBS 0.008683f
C462 B.n422 VSUBS 0.008683f
C463 B.n423 VSUBS 0.008683f
C464 B.n424 VSUBS 0.008683f
C465 B.n425 VSUBS 0.008683f
C466 B.n426 VSUBS 0.008683f
C467 B.n427 VSUBS 0.008683f
C468 B.n428 VSUBS 0.008683f
C469 B.n429 VSUBS 0.008683f
C470 B.n430 VSUBS 0.008683f
C471 B.n431 VSUBS 0.008683f
C472 B.n432 VSUBS 0.008683f
C473 B.n433 VSUBS 0.008683f
C474 B.n434 VSUBS 0.008683f
C475 B.n435 VSUBS 0.008683f
C476 B.n436 VSUBS 0.008683f
C477 B.n437 VSUBS 0.008683f
C478 B.n438 VSUBS 0.008683f
C479 B.n439 VSUBS 0.008683f
C480 B.n440 VSUBS 0.008683f
C481 B.n441 VSUBS 0.008683f
C482 B.n442 VSUBS 0.008683f
C483 B.n443 VSUBS 0.008683f
C484 B.n444 VSUBS 0.008683f
C485 B.n445 VSUBS 0.008683f
C486 B.n446 VSUBS 0.008683f
C487 B.n447 VSUBS 0.008683f
C488 B.n448 VSUBS 0.008683f
C489 B.n449 VSUBS 0.008683f
C490 B.n450 VSUBS 0.008683f
C491 B.n451 VSUBS 0.008683f
C492 B.n452 VSUBS 0.008683f
C493 B.n453 VSUBS 0.008683f
C494 B.n454 VSUBS 0.008683f
C495 B.n455 VSUBS 0.008683f
C496 B.n456 VSUBS 0.008683f
C497 B.n457 VSUBS 0.008683f
C498 B.n458 VSUBS 0.006001f
C499 B.n459 VSUBS 0.020118f
C500 B.n460 VSUBS 0.007023f
C501 B.n461 VSUBS 0.008683f
C502 B.n462 VSUBS 0.008683f
C503 B.n463 VSUBS 0.008683f
C504 B.n464 VSUBS 0.008683f
C505 B.n465 VSUBS 0.008683f
C506 B.n466 VSUBS 0.008683f
C507 B.n467 VSUBS 0.008683f
C508 B.n468 VSUBS 0.008683f
C509 B.n469 VSUBS 0.008683f
C510 B.n470 VSUBS 0.008683f
C511 B.n471 VSUBS 0.008683f
C512 B.n472 VSUBS 0.007023f
C513 B.n473 VSUBS 0.008683f
C514 B.n474 VSUBS 0.008683f
C515 B.n475 VSUBS 0.006001f
C516 B.n476 VSUBS 0.008683f
C517 B.n477 VSUBS 0.008683f
C518 B.n478 VSUBS 0.008683f
C519 B.n479 VSUBS 0.008683f
C520 B.n480 VSUBS 0.008683f
C521 B.n481 VSUBS 0.008683f
C522 B.n482 VSUBS 0.008683f
C523 B.n483 VSUBS 0.008683f
C524 B.n484 VSUBS 0.008683f
C525 B.n485 VSUBS 0.008683f
C526 B.n486 VSUBS 0.008683f
C527 B.n487 VSUBS 0.008683f
C528 B.n488 VSUBS 0.008683f
C529 B.n489 VSUBS 0.008683f
C530 B.n490 VSUBS 0.008683f
C531 B.n491 VSUBS 0.008683f
C532 B.n492 VSUBS 0.008683f
C533 B.n493 VSUBS 0.008683f
C534 B.n494 VSUBS 0.008683f
C535 B.n495 VSUBS 0.008683f
C536 B.n496 VSUBS 0.008683f
C537 B.n497 VSUBS 0.008683f
C538 B.n498 VSUBS 0.008683f
C539 B.n499 VSUBS 0.008683f
C540 B.n500 VSUBS 0.008683f
C541 B.n501 VSUBS 0.008683f
C542 B.n502 VSUBS 0.008683f
C543 B.n503 VSUBS 0.008683f
C544 B.n504 VSUBS 0.008683f
C545 B.n505 VSUBS 0.008683f
C546 B.n506 VSUBS 0.008683f
C547 B.n507 VSUBS 0.008683f
C548 B.n508 VSUBS 0.008683f
C549 B.n509 VSUBS 0.008683f
C550 B.n510 VSUBS 0.008683f
C551 B.n511 VSUBS 0.008683f
C552 B.n512 VSUBS 0.008683f
C553 B.n513 VSUBS 0.008683f
C554 B.n514 VSUBS 0.008683f
C555 B.n515 VSUBS 0.008683f
C556 B.n516 VSUBS 0.008683f
C557 B.n517 VSUBS 0.008683f
C558 B.n518 VSUBS 0.008683f
C559 B.n519 VSUBS 0.008683f
C560 B.n520 VSUBS 0.008683f
C561 B.n521 VSUBS 0.008683f
C562 B.n522 VSUBS 0.008683f
C563 B.n523 VSUBS 0.008683f
C564 B.n524 VSUBS 0.008683f
C565 B.n525 VSUBS 0.008683f
C566 B.n526 VSUBS 0.008683f
C567 B.n527 VSUBS 0.008683f
C568 B.n528 VSUBS 0.008683f
C569 B.n529 VSUBS 0.008683f
C570 B.n530 VSUBS 0.008683f
C571 B.n531 VSUBS 0.008683f
C572 B.n532 VSUBS 0.008683f
C573 B.n533 VSUBS 0.008683f
C574 B.n534 VSUBS 0.008683f
C575 B.n535 VSUBS 0.008683f
C576 B.n536 VSUBS 0.008683f
C577 B.n537 VSUBS 0.021357f
C578 B.n538 VSUBS 0.021357f
C579 B.n539 VSUBS 0.020271f
C580 B.n540 VSUBS 0.008683f
C581 B.n541 VSUBS 0.008683f
C582 B.n542 VSUBS 0.008683f
C583 B.n543 VSUBS 0.008683f
C584 B.n544 VSUBS 0.008683f
C585 B.n545 VSUBS 0.008683f
C586 B.n546 VSUBS 0.008683f
C587 B.n547 VSUBS 0.008683f
C588 B.n548 VSUBS 0.008683f
C589 B.n549 VSUBS 0.008683f
C590 B.n550 VSUBS 0.008683f
C591 B.n551 VSUBS 0.008683f
C592 B.n552 VSUBS 0.008683f
C593 B.n553 VSUBS 0.008683f
C594 B.n554 VSUBS 0.008683f
C595 B.n555 VSUBS 0.008683f
C596 B.n556 VSUBS 0.008683f
C597 B.n557 VSUBS 0.008683f
C598 B.n558 VSUBS 0.008683f
C599 B.n559 VSUBS 0.008683f
C600 B.n560 VSUBS 0.008683f
C601 B.n561 VSUBS 0.008683f
C602 B.n562 VSUBS 0.008683f
C603 B.n563 VSUBS 0.008683f
C604 B.n564 VSUBS 0.008683f
C605 B.n565 VSUBS 0.008683f
C606 B.n566 VSUBS 0.008683f
C607 B.n567 VSUBS 0.008683f
C608 B.n568 VSUBS 0.008683f
C609 B.n569 VSUBS 0.008683f
C610 B.n570 VSUBS 0.008683f
C611 B.n571 VSUBS 0.008683f
C612 B.n572 VSUBS 0.008683f
C613 B.n573 VSUBS 0.008683f
C614 B.n574 VSUBS 0.008683f
C615 B.n575 VSUBS 0.008683f
C616 B.n576 VSUBS 0.008683f
C617 B.n577 VSUBS 0.008683f
C618 B.n578 VSUBS 0.008683f
C619 B.n579 VSUBS 0.008683f
C620 B.n580 VSUBS 0.008683f
C621 B.n581 VSUBS 0.008683f
C622 B.n582 VSUBS 0.008683f
C623 B.n583 VSUBS 0.008683f
C624 B.n584 VSUBS 0.008683f
C625 B.n585 VSUBS 0.008683f
C626 B.n586 VSUBS 0.008683f
C627 B.n587 VSUBS 0.008683f
C628 B.n588 VSUBS 0.008683f
C629 B.n589 VSUBS 0.008683f
C630 B.n590 VSUBS 0.008683f
C631 B.n591 VSUBS 0.008683f
C632 B.n592 VSUBS 0.008683f
C633 B.n593 VSUBS 0.008683f
C634 B.n594 VSUBS 0.008683f
C635 B.n595 VSUBS 0.008683f
C636 B.n596 VSUBS 0.008683f
C637 B.n597 VSUBS 0.008683f
C638 B.n598 VSUBS 0.008683f
C639 B.n599 VSUBS 0.008683f
C640 B.n600 VSUBS 0.008683f
C641 B.n601 VSUBS 0.008683f
C642 B.n602 VSUBS 0.008683f
C643 B.n603 VSUBS 0.008683f
C644 B.n604 VSUBS 0.008683f
C645 B.n605 VSUBS 0.008683f
C646 B.n606 VSUBS 0.008683f
C647 B.n607 VSUBS 0.008683f
C648 B.n608 VSUBS 0.008683f
C649 B.n609 VSUBS 0.008683f
C650 B.n610 VSUBS 0.008683f
C651 B.n611 VSUBS 0.008683f
C652 B.n612 VSUBS 0.008683f
C653 B.n613 VSUBS 0.008683f
C654 B.n614 VSUBS 0.008683f
C655 B.n615 VSUBS 0.008683f
C656 B.n616 VSUBS 0.008683f
C657 B.n617 VSUBS 0.008683f
C658 B.n618 VSUBS 0.008683f
C659 B.n619 VSUBS 0.008683f
C660 B.n620 VSUBS 0.008683f
C661 B.n621 VSUBS 0.008683f
C662 B.n622 VSUBS 0.008683f
C663 B.n623 VSUBS 0.008683f
C664 B.n624 VSUBS 0.008683f
C665 B.n625 VSUBS 0.008683f
C666 B.n626 VSUBS 0.008683f
C667 B.n627 VSUBS 0.008683f
C668 B.n628 VSUBS 0.008683f
C669 B.n629 VSUBS 0.008683f
C670 B.n630 VSUBS 0.008683f
C671 B.n631 VSUBS 0.008683f
C672 B.n632 VSUBS 0.008683f
C673 B.n633 VSUBS 0.008683f
C674 B.n634 VSUBS 0.008683f
C675 B.n635 VSUBS 0.008683f
C676 B.n636 VSUBS 0.008683f
C677 B.n637 VSUBS 0.008683f
C678 B.n638 VSUBS 0.008683f
C679 B.n639 VSUBS 0.008683f
C680 B.n640 VSUBS 0.008683f
C681 B.n641 VSUBS 0.008683f
C682 B.n642 VSUBS 0.008683f
C683 B.n643 VSUBS 0.008683f
C684 B.n644 VSUBS 0.008683f
C685 B.n645 VSUBS 0.008683f
C686 B.n646 VSUBS 0.008683f
C687 B.n647 VSUBS 0.008683f
C688 B.n648 VSUBS 0.008683f
C689 B.n649 VSUBS 0.008683f
C690 B.n650 VSUBS 0.008683f
C691 B.n651 VSUBS 0.008683f
C692 B.n652 VSUBS 0.008683f
C693 B.n653 VSUBS 0.008683f
C694 B.n654 VSUBS 0.008683f
C695 B.n655 VSUBS 0.008683f
C696 B.n656 VSUBS 0.008683f
C697 B.n657 VSUBS 0.008683f
C698 B.n658 VSUBS 0.008683f
C699 B.n659 VSUBS 0.008683f
C700 B.n660 VSUBS 0.008683f
C701 B.n661 VSUBS 0.008683f
C702 B.n662 VSUBS 0.008683f
C703 B.n663 VSUBS 0.008683f
C704 B.n664 VSUBS 0.008683f
C705 B.n665 VSUBS 0.008683f
C706 B.n666 VSUBS 0.008683f
C707 B.n667 VSUBS 0.008683f
C708 B.n668 VSUBS 0.008683f
C709 B.n669 VSUBS 0.008683f
C710 B.n670 VSUBS 0.008683f
C711 B.n671 VSUBS 0.008683f
C712 B.n672 VSUBS 0.008683f
C713 B.n673 VSUBS 0.008683f
C714 B.n674 VSUBS 0.008683f
C715 B.n675 VSUBS 0.008683f
C716 B.n676 VSUBS 0.008683f
C717 B.n677 VSUBS 0.008683f
C718 B.n678 VSUBS 0.008683f
C719 B.n679 VSUBS 0.008683f
C720 B.n680 VSUBS 0.008683f
C721 B.n681 VSUBS 0.008683f
C722 B.n682 VSUBS 0.008683f
C723 B.n683 VSUBS 0.008683f
C724 B.n684 VSUBS 0.008683f
C725 B.n685 VSUBS 0.008683f
C726 B.n686 VSUBS 0.008683f
C727 B.n687 VSUBS 0.008683f
C728 B.n688 VSUBS 0.008683f
C729 B.n689 VSUBS 0.008683f
C730 B.n690 VSUBS 0.008683f
C731 B.n691 VSUBS 0.008683f
C732 B.n692 VSUBS 0.008683f
C733 B.n693 VSUBS 0.008683f
C734 B.n694 VSUBS 0.008683f
C735 B.n695 VSUBS 0.008683f
C736 B.n696 VSUBS 0.008683f
C737 B.n697 VSUBS 0.008683f
C738 B.n698 VSUBS 0.008683f
C739 B.n699 VSUBS 0.008683f
C740 B.n700 VSUBS 0.008683f
C741 B.n701 VSUBS 0.008683f
C742 B.n702 VSUBS 0.008683f
C743 B.n703 VSUBS 0.008683f
C744 B.n704 VSUBS 0.008683f
C745 B.n705 VSUBS 0.008683f
C746 B.n706 VSUBS 0.008683f
C747 B.n707 VSUBS 0.008683f
C748 B.n708 VSUBS 0.008683f
C749 B.n709 VSUBS 0.008683f
C750 B.n710 VSUBS 0.008683f
C751 B.n711 VSUBS 0.008683f
C752 B.n712 VSUBS 0.008683f
C753 B.n713 VSUBS 0.008683f
C754 B.n714 VSUBS 0.008683f
C755 B.n715 VSUBS 0.008683f
C756 B.n716 VSUBS 0.008683f
C757 B.n717 VSUBS 0.008683f
C758 B.n718 VSUBS 0.008683f
C759 B.n719 VSUBS 0.008683f
C760 B.n720 VSUBS 0.008683f
C761 B.n721 VSUBS 0.008683f
C762 B.n722 VSUBS 0.008683f
C763 B.n723 VSUBS 0.008683f
C764 B.n724 VSUBS 0.008683f
C765 B.n725 VSUBS 0.008683f
C766 B.n726 VSUBS 0.008683f
C767 B.n727 VSUBS 0.008683f
C768 B.n728 VSUBS 0.008683f
C769 B.n729 VSUBS 0.008683f
C770 B.n730 VSUBS 0.008683f
C771 B.n731 VSUBS 0.008683f
C772 B.n732 VSUBS 0.008683f
C773 B.n733 VSUBS 0.008683f
C774 B.n734 VSUBS 0.008683f
C775 B.n735 VSUBS 0.008683f
C776 B.n736 VSUBS 0.008683f
C777 B.n737 VSUBS 0.008683f
C778 B.n738 VSUBS 0.008683f
C779 B.n739 VSUBS 0.008683f
C780 B.n740 VSUBS 0.008683f
C781 B.n741 VSUBS 0.008683f
C782 B.n742 VSUBS 0.008683f
C783 B.n743 VSUBS 0.008683f
C784 B.n744 VSUBS 0.008683f
C785 B.n745 VSUBS 0.008683f
C786 B.n746 VSUBS 0.008683f
C787 B.n747 VSUBS 0.008683f
C788 B.n748 VSUBS 0.008683f
C789 B.n749 VSUBS 0.008683f
C790 B.n750 VSUBS 0.008683f
C791 B.n751 VSUBS 0.008683f
C792 B.n752 VSUBS 0.008683f
C793 B.n753 VSUBS 0.008683f
C794 B.n754 VSUBS 0.008683f
C795 B.n755 VSUBS 0.008683f
C796 B.n756 VSUBS 0.008683f
C797 B.n757 VSUBS 0.008683f
C798 B.n758 VSUBS 0.008683f
C799 B.n759 VSUBS 0.008683f
C800 B.n760 VSUBS 0.008683f
C801 B.n761 VSUBS 0.008683f
C802 B.n762 VSUBS 0.008683f
C803 B.n763 VSUBS 0.008683f
C804 B.n764 VSUBS 0.008683f
C805 B.n765 VSUBS 0.008683f
C806 B.n766 VSUBS 0.008683f
C807 B.n767 VSUBS 0.008683f
C808 B.n768 VSUBS 0.008683f
C809 B.n769 VSUBS 0.008683f
C810 B.n770 VSUBS 0.008683f
C811 B.n771 VSUBS 0.008683f
C812 B.n772 VSUBS 0.008683f
C813 B.n773 VSUBS 0.008683f
C814 B.n774 VSUBS 0.008683f
C815 B.n775 VSUBS 0.008683f
C816 B.n776 VSUBS 0.008683f
C817 B.n777 VSUBS 0.008683f
C818 B.n778 VSUBS 0.008683f
C819 B.n779 VSUBS 0.008683f
C820 B.n780 VSUBS 0.008683f
C821 B.n781 VSUBS 0.008683f
C822 B.n782 VSUBS 0.008683f
C823 B.n783 VSUBS 0.008683f
C824 B.n784 VSUBS 0.008683f
C825 B.n785 VSUBS 0.008683f
C826 B.n786 VSUBS 0.008683f
C827 B.n787 VSUBS 0.008683f
C828 B.n788 VSUBS 0.02126f
C829 B.n789 VSUBS 0.020367f
C830 B.n790 VSUBS 0.021357f
C831 B.n791 VSUBS 0.008683f
C832 B.n792 VSUBS 0.008683f
C833 B.n793 VSUBS 0.008683f
C834 B.n794 VSUBS 0.008683f
C835 B.n795 VSUBS 0.008683f
C836 B.n796 VSUBS 0.008683f
C837 B.n797 VSUBS 0.008683f
C838 B.n798 VSUBS 0.008683f
C839 B.n799 VSUBS 0.008683f
C840 B.n800 VSUBS 0.008683f
C841 B.n801 VSUBS 0.008683f
C842 B.n802 VSUBS 0.008683f
C843 B.n803 VSUBS 0.008683f
C844 B.n804 VSUBS 0.008683f
C845 B.n805 VSUBS 0.008683f
C846 B.n806 VSUBS 0.008683f
C847 B.n807 VSUBS 0.008683f
C848 B.n808 VSUBS 0.008683f
C849 B.n809 VSUBS 0.008683f
C850 B.n810 VSUBS 0.008683f
C851 B.n811 VSUBS 0.008683f
C852 B.n812 VSUBS 0.008683f
C853 B.n813 VSUBS 0.008683f
C854 B.n814 VSUBS 0.008683f
C855 B.n815 VSUBS 0.008683f
C856 B.n816 VSUBS 0.008683f
C857 B.n817 VSUBS 0.008683f
C858 B.n818 VSUBS 0.008683f
C859 B.n819 VSUBS 0.008683f
C860 B.n820 VSUBS 0.008683f
C861 B.n821 VSUBS 0.008683f
C862 B.n822 VSUBS 0.008683f
C863 B.n823 VSUBS 0.008683f
C864 B.n824 VSUBS 0.008683f
C865 B.n825 VSUBS 0.008683f
C866 B.n826 VSUBS 0.008683f
C867 B.n827 VSUBS 0.008683f
C868 B.n828 VSUBS 0.008683f
C869 B.n829 VSUBS 0.008683f
C870 B.n830 VSUBS 0.008683f
C871 B.n831 VSUBS 0.008683f
C872 B.n832 VSUBS 0.008683f
C873 B.n833 VSUBS 0.008683f
C874 B.n834 VSUBS 0.008683f
C875 B.n835 VSUBS 0.008683f
C876 B.n836 VSUBS 0.008683f
C877 B.n837 VSUBS 0.008683f
C878 B.n838 VSUBS 0.008683f
C879 B.n839 VSUBS 0.008683f
C880 B.n840 VSUBS 0.008683f
C881 B.n841 VSUBS 0.008683f
C882 B.n842 VSUBS 0.008683f
C883 B.n843 VSUBS 0.008683f
C884 B.n844 VSUBS 0.008683f
C885 B.n845 VSUBS 0.008683f
C886 B.n846 VSUBS 0.008683f
C887 B.n847 VSUBS 0.008683f
C888 B.n848 VSUBS 0.008683f
C889 B.n849 VSUBS 0.008683f
C890 B.n850 VSUBS 0.008683f
C891 B.n851 VSUBS 0.008683f
C892 B.n852 VSUBS 0.008683f
C893 B.n853 VSUBS 0.006001f
C894 B.n854 VSUBS 0.020118f
C895 B.n855 VSUBS 0.007023f
C896 B.n856 VSUBS 0.008683f
C897 B.n857 VSUBS 0.008683f
C898 B.n858 VSUBS 0.008683f
C899 B.n859 VSUBS 0.008683f
C900 B.n860 VSUBS 0.008683f
C901 B.n861 VSUBS 0.008683f
C902 B.n862 VSUBS 0.008683f
C903 B.n863 VSUBS 0.008683f
C904 B.n864 VSUBS 0.008683f
C905 B.n865 VSUBS 0.008683f
C906 B.n866 VSUBS 0.008683f
C907 B.n867 VSUBS 0.007023f
C908 B.n868 VSUBS 0.020118f
C909 B.n869 VSUBS 0.006001f
C910 B.n870 VSUBS 0.008683f
C911 B.n871 VSUBS 0.008683f
C912 B.n872 VSUBS 0.008683f
C913 B.n873 VSUBS 0.008683f
C914 B.n874 VSUBS 0.008683f
C915 B.n875 VSUBS 0.008683f
C916 B.n876 VSUBS 0.008683f
C917 B.n877 VSUBS 0.008683f
C918 B.n878 VSUBS 0.008683f
C919 B.n879 VSUBS 0.008683f
C920 B.n880 VSUBS 0.008683f
C921 B.n881 VSUBS 0.008683f
C922 B.n882 VSUBS 0.008683f
C923 B.n883 VSUBS 0.008683f
C924 B.n884 VSUBS 0.008683f
C925 B.n885 VSUBS 0.008683f
C926 B.n886 VSUBS 0.008683f
C927 B.n887 VSUBS 0.008683f
C928 B.n888 VSUBS 0.008683f
C929 B.n889 VSUBS 0.008683f
C930 B.n890 VSUBS 0.008683f
C931 B.n891 VSUBS 0.008683f
C932 B.n892 VSUBS 0.008683f
C933 B.n893 VSUBS 0.008683f
C934 B.n894 VSUBS 0.008683f
C935 B.n895 VSUBS 0.008683f
C936 B.n896 VSUBS 0.008683f
C937 B.n897 VSUBS 0.008683f
C938 B.n898 VSUBS 0.008683f
C939 B.n899 VSUBS 0.008683f
C940 B.n900 VSUBS 0.008683f
C941 B.n901 VSUBS 0.008683f
C942 B.n902 VSUBS 0.008683f
C943 B.n903 VSUBS 0.008683f
C944 B.n904 VSUBS 0.008683f
C945 B.n905 VSUBS 0.008683f
C946 B.n906 VSUBS 0.008683f
C947 B.n907 VSUBS 0.008683f
C948 B.n908 VSUBS 0.008683f
C949 B.n909 VSUBS 0.008683f
C950 B.n910 VSUBS 0.008683f
C951 B.n911 VSUBS 0.008683f
C952 B.n912 VSUBS 0.008683f
C953 B.n913 VSUBS 0.008683f
C954 B.n914 VSUBS 0.008683f
C955 B.n915 VSUBS 0.008683f
C956 B.n916 VSUBS 0.008683f
C957 B.n917 VSUBS 0.008683f
C958 B.n918 VSUBS 0.008683f
C959 B.n919 VSUBS 0.008683f
C960 B.n920 VSUBS 0.008683f
C961 B.n921 VSUBS 0.008683f
C962 B.n922 VSUBS 0.008683f
C963 B.n923 VSUBS 0.008683f
C964 B.n924 VSUBS 0.008683f
C965 B.n925 VSUBS 0.008683f
C966 B.n926 VSUBS 0.008683f
C967 B.n927 VSUBS 0.008683f
C968 B.n928 VSUBS 0.008683f
C969 B.n929 VSUBS 0.008683f
C970 B.n930 VSUBS 0.008683f
C971 B.n931 VSUBS 0.008683f
C972 B.n932 VSUBS 0.021357f
C973 B.n933 VSUBS 0.021357f
C974 B.n934 VSUBS 0.020271f
C975 B.n935 VSUBS 0.008683f
C976 B.n936 VSUBS 0.008683f
C977 B.n937 VSUBS 0.008683f
C978 B.n938 VSUBS 0.008683f
C979 B.n939 VSUBS 0.008683f
C980 B.n940 VSUBS 0.008683f
C981 B.n941 VSUBS 0.008683f
C982 B.n942 VSUBS 0.008683f
C983 B.n943 VSUBS 0.008683f
C984 B.n944 VSUBS 0.008683f
C985 B.n945 VSUBS 0.008683f
C986 B.n946 VSUBS 0.008683f
C987 B.n947 VSUBS 0.008683f
C988 B.n948 VSUBS 0.008683f
C989 B.n949 VSUBS 0.008683f
C990 B.n950 VSUBS 0.008683f
C991 B.n951 VSUBS 0.008683f
C992 B.n952 VSUBS 0.008683f
C993 B.n953 VSUBS 0.008683f
C994 B.n954 VSUBS 0.008683f
C995 B.n955 VSUBS 0.008683f
C996 B.n956 VSUBS 0.008683f
C997 B.n957 VSUBS 0.008683f
C998 B.n958 VSUBS 0.008683f
C999 B.n959 VSUBS 0.008683f
C1000 B.n960 VSUBS 0.008683f
C1001 B.n961 VSUBS 0.008683f
C1002 B.n962 VSUBS 0.008683f
C1003 B.n963 VSUBS 0.008683f
C1004 B.n964 VSUBS 0.008683f
C1005 B.n965 VSUBS 0.008683f
C1006 B.n966 VSUBS 0.008683f
C1007 B.n967 VSUBS 0.008683f
C1008 B.n968 VSUBS 0.008683f
C1009 B.n969 VSUBS 0.008683f
C1010 B.n970 VSUBS 0.008683f
C1011 B.n971 VSUBS 0.008683f
C1012 B.n972 VSUBS 0.008683f
C1013 B.n973 VSUBS 0.008683f
C1014 B.n974 VSUBS 0.008683f
C1015 B.n975 VSUBS 0.008683f
C1016 B.n976 VSUBS 0.008683f
C1017 B.n977 VSUBS 0.008683f
C1018 B.n978 VSUBS 0.008683f
C1019 B.n979 VSUBS 0.008683f
C1020 B.n980 VSUBS 0.008683f
C1021 B.n981 VSUBS 0.008683f
C1022 B.n982 VSUBS 0.008683f
C1023 B.n983 VSUBS 0.008683f
C1024 B.n984 VSUBS 0.008683f
C1025 B.n985 VSUBS 0.008683f
C1026 B.n986 VSUBS 0.008683f
C1027 B.n987 VSUBS 0.008683f
C1028 B.n988 VSUBS 0.008683f
C1029 B.n989 VSUBS 0.008683f
C1030 B.n990 VSUBS 0.008683f
C1031 B.n991 VSUBS 0.008683f
C1032 B.n992 VSUBS 0.008683f
C1033 B.n993 VSUBS 0.008683f
C1034 B.n994 VSUBS 0.008683f
C1035 B.n995 VSUBS 0.008683f
C1036 B.n996 VSUBS 0.008683f
C1037 B.n997 VSUBS 0.008683f
C1038 B.n998 VSUBS 0.008683f
C1039 B.n999 VSUBS 0.008683f
C1040 B.n1000 VSUBS 0.008683f
C1041 B.n1001 VSUBS 0.008683f
C1042 B.n1002 VSUBS 0.008683f
C1043 B.n1003 VSUBS 0.008683f
C1044 B.n1004 VSUBS 0.008683f
C1045 B.n1005 VSUBS 0.008683f
C1046 B.n1006 VSUBS 0.008683f
C1047 B.n1007 VSUBS 0.008683f
C1048 B.n1008 VSUBS 0.008683f
C1049 B.n1009 VSUBS 0.008683f
C1050 B.n1010 VSUBS 0.008683f
C1051 B.n1011 VSUBS 0.008683f
C1052 B.n1012 VSUBS 0.008683f
C1053 B.n1013 VSUBS 0.008683f
C1054 B.n1014 VSUBS 0.008683f
C1055 B.n1015 VSUBS 0.008683f
C1056 B.n1016 VSUBS 0.008683f
C1057 B.n1017 VSUBS 0.008683f
C1058 B.n1018 VSUBS 0.008683f
C1059 B.n1019 VSUBS 0.008683f
C1060 B.n1020 VSUBS 0.008683f
C1061 B.n1021 VSUBS 0.008683f
C1062 B.n1022 VSUBS 0.008683f
C1063 B.n1023 VSUBS 0.008683f
C1064 B.n1024 VSUBS 0.008683f
C1065 B.n1025 VSUBS 0.008683f
C1066 B.n1026 VSUBS 0.008683f
C1067 B.n1027 VSUBS 0.008683f
C1068 B.n1028 VSUBS 0.008683f
C1069 B.n1029 VSUBS 0.008683f
C1070 B.n1030 VSUBS 0.008683f
C1071 B.n1031 VSUBS 0.008683f
C1072 B.n1032 VSUBS 0.008683f
C1073 B.n1033 VSUBS 0.008683f
C1074 B.n1034 VSUBS 0.008683f
C1075 B.n1035 VSUBS 0.008683f
C1076 B.n1036 VSUBS 0.008683f
C1077 B.n1037 VSUBS 0.008683f
C1078 B.n1038 VSUBS 0.008683f
C1079 B.n1039 VSUBS 0.008683f
C1080 B.n1040 VSUBS 0.008683f
C1081 B.n1041 VSUBS 0.008683f
C1082 B.n1042 VSUBS 0.008683f
C1083 B.n1043 VSUBS 0.008683f
C1084 B.n1044 VSUBS 0.008683f
C1085 B.n1045 VSUBS 0.008683f
C1086 B.n1046 VSUBS 0.008683f
C1087 B.n1047 VSUBS 0.008683f
C1088 B.n1048 VSUBS 0.008683f
C1089 B.n1049 VSUBS 0.008683f
C1090 B.n1050 VSUBS 0.008683f
C1091 B.n1051 VSUBS 0.008683f
C1092 B.n1052 VSUBS 0.008683f
C1093 B.n1053 VSUBS 0.008683f
C1094 B.n1054 VSUBS 0.008683f
C1095 B.n1055 VSUBS 0.008683f
C1096 B.n1056 VSUBS 0.008683f
C1097 B.n1057 VSUBS 0.008683f
C1098 B.n1058 VSUBS 0.008683f
C1099 B.n1059 VSUBS 0.019661f
C1100 VDD1.t7 VSUBS 3.15739f
C1101 VDD1.t6 VSUBS 0.304512f
C1102 VDD1.t3 VSUBS 0.304512f
C1103 VDD1.n0 VSUBS 2.37892f
C1104 VDD1.n1 VSUBS 2.09272f
C1105 VDD1.t9 VSUBS 3.15738f
C1106 VDD1.t1 VSUBS 0.304512f
C1107 VDD1.t0 VSUBS 0.304512f
C1108 VDD1.n2 VSUBS 2.37891f
C1109 VDD1.n3 VSUBS 2.08219f
C1110 VDD1.t4 VSUBS 0.304512f
C1111 VDD1.t5 VSUBS 0.304512f
C1112 VDD1.n4 VSUBS 2.42422f
C1113 VDD1.n5 VSUBS 5.03621f
C1114 VDD1.t2 VSUBS 0.304512f
C1115 VDD1.t8 VSUBS 0.304512f
C1116 VDD1.n6 VSUBS 2.3789f
C1117 VDD1.n7 VSUBS 5.00959f
C1118 VP.n0 VSUBS 0.046381f
C1119 VP.t4 VSUBS 3.26225f
C1120 VP.n1 VSUBS 0.048814f
C1121 VP.n2 VSUBS 0.02465f
C1122 VP.n3 VSUBS 0.046172f
C1123 VP.n4 VSUBS 0.02465f
C1124 VP.t5 VSUBS 3.26225f
C1125 VP.n5 VSUBS 0.046172f
C1126 VP.n6 VSUBS 0.02465f
C1127 VP.n7 VSUBS 0.046172f
C1128 VP.n8 VSUBS 0.02465f
C1129 VP.t9 VSUBS 3.26225f
C1130 VP.n9 VSUBS 0.046172f
C1131 VP.n10 VSUBS 0.02465f
C1132 VP.n11 VSUBS 0.046172f
C1133 VP.n12 VSUBS 0.02465f
C1134 VP.t8 VSUBS 3.26225f
C1135 VP.n13 VSUBS 0.046172f
C1136 VP.n14 VSUBS 0.02465f
C1137 VP.n15 VSUBS 0.048814f
C1138 VP.n16 VSUBS 0.046381f
C1139 VP.t0 VSUBS 3.26225f
C1140 VP.n17 VSUBS 0.046381f
C1141 VP.t1 VSUBS 3.26225f
C1142 VP.n18 VSUBS 0.048814f
C1143 VP.n19 VSUBS 0.02465f
C1144 VP.n20 VSUBS 0.046172f
C1145 VP.n21 VSUBS 0.02465f
C1146 VP.t7 VSUBS 3.26225f
C1147 VP.n22 VSUBS 0.046172f
C1148 VP.n23 VSUBS 0.02465f
C1149 VP.n24 VSUBS 0.046172f
C1150 VP.n25 VSUBS 0.02465f
C1151 VP.t6 VSUBS 3.26225f
C1152 VP.n26 VSUBS 0.046172f
C1153 VP.n27 VSUBS 0.02465f
C1154 VP.n28 VSUBS 0.046172f
C1155 VP.n29 VSUBS 0.322481f
C1156 VP.t3 VSUBS 3.26225f
C1157 VP.t2 VSUBS 3.65836f
C1158 VP.n30 VSUBS 1.17732f
C1159 VP.n31 VSUBS 1.23049f
C1160 VP.n32 VSUBS 0.034774f
C1161 VP.n33 VSUBS 0.046172f
C1162 VP.n34 VSUBS 0.02465f
C1163 VP.n35 VSUBS 0.02465f
C1164 VP.n36 VSUBS 0.02465f
C1165 VP.n37 VSUBS 0.044214f
C1166 VP.n38 VSUBS 0.025429f
C1167 VP.n39 VSUBS 0.048814f
C1168 VP.n40 VSUBS 0.02465f
C1169 VP.n41 VSUBS 0.02465f
C1170 VP.n42 VSUBS 0.02465f
C1171 VP.n43 VSUBS 0.046172f
C1172 VP.n44 VSUBS 1.16368f
C1173 VP.n45 VSUBS 0.046172f
C1174 VP.n46 VSUBS 0.02465f
C1175 VP.n47 VSUBS 0.02465f
C1176 VP.n48 VSUBS 0.02465f
C1177 VP.n49 VSUBS 0.048814f
C1178 VP.n50 VSUBS 0.025429f
C1179 VP.n51 VSUBS 0.044214f
C1180 VP.n52 VSUBS 0.02465f
C1181 VP.n53 VSUBS 0.02465f
C1182 VP.n54 VSUBS 0.02465f
C1183 VP.n55 VSUBS 0.046172f
C1184 VP.n56 VSUBS 0.034774f
C1185 VP.n57 VSUBS 1.1403f
C1186 VP.n58 VSUBS 0.034774f
C1187 VP.n59 VSUBS 0.02465f
C1188 VP.n60 VSUBS 0.02465f
C1189 VP.n61 VSUBS 0.02465f
C1190 VP.n62 VSUBS 0.046172f
C1191 VP.n63 VSUBS 0.044214f
C1192 VP.n64 VSUBS 0.025429f
C1193 VP.n65 VSUBS 0.02465f
C1194 VP.n66 VSUBS 0.02465f
C1195 VP.n67 VSUBS 0.02465f
C1196 VP.n68 VSUBS 0.046172f
C1197 VP.n69 VSUBS 0.046172f
C1198 VP.n70 VSUBS 1.25588f
C1199 VP.n71 VSUBS 1.86814f
C1200 VP.n72 VSUBS 1.88266f
C1201 VP.n73 VSUBS 1.25588f
C1202 VP.n74 VSUBS 0.046172f
C1203 VP.n75 VSUBS 0.046172f
C1204 VP.n76 VSUBS 0.02465f
C1205 VP.n77 VSUBS 0.02465f
C1206 VP.n78 VSUBS 0.02465f
C1207 VP.n79 VSUBS 0.025429f
C1208 VP.n80 VSUBS 0.044214f
C1209 VP.n81 VSUBS 0.046172f
C1210 VP.n82 VSUBS 0.02465f
C1211 VP.n83 VSUBS 0.02465f
C1212 VP.n84 VSUBS 0.02465f
C1213 VP.n85 VSUBS 0.034774f
C1214 VP.n86 VSUBS 1.1403f
C1215 VP.n87 VSUBS 0.034774f
C1216 VP.n88 VSUBS 0.046172f
C1217 VP.n89 VSUBS 0.02465f
C1218 VP.n90 VSUBS 0.02465f
C1219 VP.n91 VSUBS 0.02465f
C1220 VP.n92 VSUBS 0.044214f
C1221 VP.n93 VSUBS 0.025429f
C1222 VP.n94 VSUBS 0.048814f
C1223 VP.n95 VSUBS 0.02465f
C1224 VP.n96 VSUBS 0.02465f
C1225 VP.n97 VSUBS 0.02465f
C1226 VP.n98 VSUBS 0.046172f
C1227 VP.n99 VSUBS 1.16368f
C1228 VP.n100 VSUBS 0.046172f
C1229 VP.n101 VSUBS 0.02465f
C1230 VP.n102 VSUBS 0.02465f
C1231 VP.n103 VSUBS 0.02465f
C1232 VP.n104 VSUBS 0.048814f
C1233 VP.n105 VSUBS 0.025429f
C1234 VP.n106 VSUBS 0.044214f
C1235 VP.n107 VSUBS 0.02465f
C1236 VP.n108 VSUBS 0.02465f
C1237 VP.n109 VSUBS 0.02465f
C1238 VP.n110 VSUBS 0.046172f
C1239 VP.n111 VSUBS 0.034774f
C1240 VP.n112 VSUBS 1.1403f
C1241 VP.n113 VSUBS 0.034774f
C1242 VP.n114 VSUBS 0.02465f
C1243 VP.n115 VSUBS 0.02465f
C1244 VP.n116 VSUBS 0.02465f
C1245 VP.n117 VSUBS 0.046172f
C1246 VP.n118 VSUBS 0.044214f
C1247 VP.n119 VSUBS 0.025429f
C1248 VP.n120 VSUBS 0.02465f
C1249 VP.n121 VSUBS 0.02465f
C1250 VP.n122 VSUBS 0.02465f
C1251 VP.n123 VSUBS 0.046172f
C1252 VP.n124 VSUBS 0.046172f
C1253 VP.n125 VSUBS 1.25588f
C1254 VP.n126 VSUBS 0.07191f
C1255 VDD2.t6 VSUBS 3.15882f
C1256 VDD2.t4 VSUBS 0.304651f
C1257 VDD2.t1 VSUBS 0.304651f
C1258 VDD2.n0 VSUBS 2.38f
C1259 VDD2.n1 VSUBS 2.08314f
C1260 VDD2.t3 VSUBS 0.304651f
C1261 VDD2.t9 VSUBS 0.304651f
C1262 VDD2.n2 VSUBS 2.42533f
C1263 VDD2.n3 VSUBS 4.83683f
C1264 VDD2.t0 VSUBS 3.10789f
C1265 VDD2.n4 VSUBS 4.93161f
C1266 VDD2.t5 VSUBS 0.304651f
C1267 VDD2.t7 VSUBS 0.304651f
C1268 VDD2.n5 VSUBS 2.38f
C1269 VDD2.n6 VSUBS 1.06342f
C1270 VDD2.t2 VSUBS 0.304651f
C1271 VDD2.t8 VSUBS 0.304651f
C1272 VDD2.n7 VSUBS 2.42526f
C1273 VTAIL.t15 VSUBS 0.293627f
C1274 VTAIL.t18 VSUBS 0.293627f
C1275 VTAIL.n0 VSUBS 2.12015f
C1276 VTAIL.n1 VSUBS 1.20331f
C1277 VTAIL.t4 VSUBS 2.8008f
C1278 VTAIL.n2 VSUBS 1.40641f
C1279 VTAIL.t3 VSUBS 0.293627f
C1280 VTAIL.t2 VSUBS 0.293627f
C1281 VTAIL.n3 VSUBS 2.12015f
C1282 VTAIL.n4 VSUBS 1.41799f
C1283 VTAIL.t5 VSUBS 0.293627f
C1284 VTAIL.t8 VSUBS 0.293627f
C1285 VTAIL.n5 VSUBS 2.12015f
C1286 VTAIL.n6 VSUBS 3.21216f
C1287 VTAIL.t19 VSUBS 0.293627f
C1288 VTAIL.t10 VSUBS 0.293627f
C1289 VTAIL.n7 VSUBS 2.12016f
C1290 VTAIL.n8 VSUBS 3.21215f
C1291 VTAIL.t14 VSUBS 0.293627f
C1292 VTAIL.t12 VSUBS 0.293627f
C1293 VTAIL.n9 VSUBS 2.12016f
C1294 VTAIL.n10 VSUBS 1.41798f
C1295 VTAIL.t13 VSUBS 2.80082f
C1296 VTAIL.n11 VSUBS 1.40639f
C1297 VTAIL.t0 VSUBS 0.293627f
C1298 VTAIL.t6 VSUBS 0.293627f
C1299 VTAIL.n12 VSUBS 2.12016f
C1300 VTAIL.n13 VSUBS 1.28625f
C1301 VTAIL.t1 VSUBS 0.293627f
C1302 VTAIL.t9 VSUBS 0.293627f
C1303 VTAIL.n14 VSUBS 2.12016f
C1304 VTAIL.n15 VSUBS 1.41798f
C1305 VTAIL.t7 VSUBS 2.8008f
C1306 VTAIL.n16 VSUBS 2.97798f
C1307 VTAIL.t11 VSUBS 2.8008f
C1308 VTAIL.n17 VSUBS 2.97798f
C1309 VTAIL.t16 VSUBS 0.293627f
C1310 VTAIL.t17 VSUBS 0.293627f
C1311 VTAIL.n18 VSUBS 2.12015f
C1312 VTAIL.n19 VSUBS 1.14661f
C1313 VN.n0 VSUBS 0.042502f
C1314 VN.t0 VSUBS 2.98946f
C1315 VN.n1 VSUBS 0.044732f
C1316 VN.n2 VSUBS 0.022589f
C1317 VN.n3 VSUBS 0.042312f
C1318 VN.n4 VSUBS 0.022589f
C1319 VN.t6 VSUBS 2.98946f
C1320 VN.n5 VSUBS 0.042312f
C1321 VN.n6 VSUBS 0.022589f
C1322 VN.n7 VSUBS 0.042312f
C1323 VN.n8 VSUBS 0.022589f
C1324 VN.t8 VSUBS 2.98946f
C1325 VN.n9 VSUBS 0.042312f
C1326 VN.n10 VSUBS 0.022589f
C1327 VN.n11 VSUBS 0.042312f
C1328 VN.n12 VSUBS 0.295515f
C1329 VN.t5 VSUBS 2.98946f
C1330 VN.t3 VSUBS 3.35246f
C1331 VN.n13 VSUBS 1.07887f
C1332 VN.n14 VSUBS 1.1276f
C1333 VN.n15 VSUBS 0.031866f
C1334 VN.n16 VSUBS 0.042312f
C1335 VN.n17 VSUBS 0.022589f
C1336 VN.n18 VSUBS 0.022589f
C1337 VN.n19 VSUBS 0.022589f
C1338 VN.n20 VSUBS 0.040516f
C1339 VN.n21 VSUBS 0.023302f
C1340 VN.n22 VSUBS 0.044732f
C1341 VN.n23 VSUBS 0.022589f
C1342 VN.n24 VSUBS 0.022589f
C1343 VN.n25 VSUBS 0.022589f
C1344 VN.n26 VSUBS 0.042312f
C1345 VN.n27 VSUBS 1.06637f
C1346 VN.n28 VSUBS 0.042312f
C1347 VN.n29 VSUBS 0.022589f
C1348 VN.n30 VSUBS 0.022589f
C1349 VN.n31 VSUBS 0.022589f
C1350 VN.n32 VSUBS 0.044732f
C1351 VN.n33 VSUBS 0.023302f
C1352 VN.n34 VSUBS 0.040516f
C1353 VN.n35 VSUBS 0.022589f
C1354 VN.n36 VSUBS 0.022589f
C1355 VN.n37 VSUBS 0.022589f
C1356 VN.n38 VSUBS 0.042312f
C1357 VN.n39 VSUBS 0.031866f
C1358 VN.n40 VSUBS 1.04495f
C1359 VN.n41 VSUBS 0.031866f
C1360 VN.n42 VSUBS 0.022589f
C1361 VN.n43 VSUBS 0.022589f
C1362 VN.n44 VSUBS 0.022589f
C1363 VN.n45 VSUBS 0.042312f
C1364 VN.n46 VSUBS 0.040516f
C1365 VN.n47 VSUBS 0.023302f
C1366 VN.n48 VSUBS 0.022589f
C1367 VN.n49 VSUBS 0.022589f
C1368 VN.n50 VSUBS 0.022589f
C1369 VN.n51 VSUBS 0.042312f
C1370 VN.n52 VSUBS 0.042312f
C1371 VN.n53 VSUBS 1.15087f
C1372 VN.n54 VSUBS 0.065897f
C1373 VN.n55 VSUBS 0.042502f
C1374 VN.t9 VSUBS 2.98946f
C1375 VN.n56 VSUBS 0.044732f
C1376 VN.n57 VSUBS 0.022589f
C1377 VN.n58 VSUBS 0.042312f
C1378 VN.n59 VSUBS 0.022589f
C1379 VN.t4 VSUBS 2.98946f
C1380 VN.n60 VSUBS 0.042312f
C1381 VN.n61 VSUBS 0.022589f
C1382 VN.n62 VSUBS 0.042312f
C1383 VN.n63 VSUBS 0.022589f
C1384 VN.t2 VSUBS 2.98946f
C1385 VN.n64 VSUBS 0.042312f
C1386 VN.n65 VSUBS 0.022589f
C1387 VN.n66 VSUBS 0.042312f
C1388 VN.n67 VSUBS 0.295515f
C1389 VN.t7 VSUBS 2.98946f
C1390 VN.t1 VSUBS 3.35246f
C1391 VN.n68 VSUBS 1.07887f
C1392 VN.n69 VSUBS 1.1276f
C1393 VN.n70 VSUBS 0.031866f
C1394 VN.n71 VSUBS 0.042312f
C1395 VN.n72 VSUBS 0.022589f
C1396 VN.n73 VSUBS 0.022589f
C1397 VN.n74 VSUBS 0.022589f
C1398 VN.n75 VSUBS 0.040516f
C1399 VN.n76 VSUBS 0.023302f
C1400 VN.n77 VSUBS 0.044732f
C1401 VN.n78 VSUBS 0.022589f
C1402 VN.n79 VSUBS 0.022589f
C1403 VN.n80 VSUBS 0.022589f
C1404 VN.n81 VSUBS 0.042312f
C1405 VN.n82 VSUBS 1.06637f
C1406 VN.n83 VSUBS 0.042312f
C1407 VN.n84 VSUBS 0.022589f
C1408 VN.n85 VSUBS 0.022589f
C1409 VN.n86 VSUBS 0.022589f
C1410 VN.n87 VSUBS 0.044732f
C1411 VN.n88 VSUBS 0.023302f
C1412 VN.n89 VSUBS 0.040516f
C1413 VN.n90 VSUBS 0.022589f
C1414 VN.n91 VSUBS 0.022589f
C1415 VN.n92 VSUBS 0.022589f
C1416 VN.n93 VSUBS 0.042312f
C1417 VN.n94 VSUBS 0.031866f
C1418 VN.n95 VSUBS 1.04495f
C1419 VN.n96 VSUBS 0.031866f
C1420 VN.n97 VSUBS 0.022589f
C1421 VN.n98 VSUBS 0.022589f
C1422 VN.n99 VSUBS 0.022589f
C1423 VN.n100 VSUBS 0.042312f
C1424 VN.n101 VSUBS 0.040516f
C1425 VN.n102 VSUBS 0.023302f
C1426 VN.n103 VSUBS 0.022589f
C1427 VN.n104 VSUBS 0.022589f
C1428 VN.n105 VSUBS 0.022589f
C1429 VN.n106 VSUBS 0.042312f
C1430 VN.n107 VSUBS 0.042312f
C1431 VN.n108 VSUBS 1.15087f
C1432 VN.n109 VSUBS 1.71703f
.ends

