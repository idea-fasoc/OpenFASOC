* NGSPICE file created from diff_pair_sample_0188.ext - technology: sky130A

.subckt diff_pair_sample_0188 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=0.94
X1 B.t8 B.t6 B.t7 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=0.94
X2 VTAIL.t6 VN.t0 VDD2.t1 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=0.94
X3 VTAIL.t5 VN.t1 VDD2.t0 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=0.94
X4 VDD2.t3 VN.t2 VTAIL.t4 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=0.94
X5 VTAIL.t7 VP.t0 VDD1.t3 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=0.94
X6 VDD2.t2 VN.t3 VTAIL.t3 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=0.94
X7 VDD1.t2 VP.t1 VTAIL.t2 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=0.94
X8 VTAIL.t1 VP.t2 VDD1.t1 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=0.94
X9 B.t5 B.t3 B.t4 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=0.94
X10 B.t2 B.t0 B.t1 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=0.94
X11 VDD1.t0 VP.t3 VTAIL.t0 w_n1732_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=0.94
R0 B.n327 B.n86 585
R1 B.n326 B.n325 585
R2 B.n324 B.n87 585
R3 B.n323 B.n322 585
R4 B.n321 B.n88 585
R5 B.n320 B.n319 585
R6 B.n318 B.n89 585
R7 B.n317 B.n316 585
R8 B.n315 B.n90 585
R9 B.n314 B.n313 585
R10 B.n312 B.n91 585
R11 B.n311 B.n310 585
R12 B.n309 B.n92 585
R13 B.n308 B.n307 585
R14 B.n306 B.n93 585
R15 B.n305 B.n304 585
R16 B.n303 B.n94 585
R17 B.n302 B.n301 585
R18 B.n300 B.n95 585
R19 B.n299 B.n298 585
R20 B.n297 B.n96 585
R21 B.n296 B.n295 585
R22 B.n294 B.n97 585
R23 B.n293 B.n292 585
R24 B.n291 B.n98 585
R25 B.n290 B.n289 585
R26 B.n288 B.n99 585
R27 B.n287 B.n286 585
R28 B.n285 B.n100 585
R29 B.n284 B.n283 585
R30 B.n282 B.n101 585
R31 B.n281 B.n280 585
R32 B.n279 B.n102 585
R33 B.n278 B.n277 585
R34 B.n276 B.n103 585
R35 B.n275 B.n274 585
R36 B.n273 B.n104 585
R37 B.n272 B.n271 585
R38 B.n270 B.n105 585
R39 B.n269 B.n268 585
R40 B.n267 B.n106 585
R41 B.n266 B.n265 585
R42 B.n264 B.n107 585
R43 B.n263 B.n262 585
R44 B.n261 B.n108 585
R45 B.n260 B.n259 585
R46 B.n255 B.n109 585
R47 B.n254 B.n253 585
R48 B.n252 B.n110 585
R49 B.n251 B.n250 585
R50 B.n249 B.n111 585
R51 B.n248 B.n247 585
R52 B.n246 B.n112 585
R53 B.n245 B.n244 585
R54 B.n243 B.n113 585
R55 B.n241 B.n240 585
R56 B.n239 B.n116 585
R57 B.n238 B.n237 585
R58 B.n236 B.n117 585
R59 B.n235 B.n234 585
R60 B.n233 B.n118 585
R61 B.n232 B.n231 585
R62 B.n230 B.n119 585
R63 B.n229 B.n228 585
R64 B.n227 B.n120 585
R65 B.n226 B.n225 585
R66 B.n224 B.n121 585
R67 B.n223 B.n222 585
R68 B.n221 B.n122 585
R69 B.n220 B.n219 585
R70 B.n218 B.n123 585
R71 B.n217 B.n216 585
R72 B.n215 B.n124 585
R73 B.n214 B.n213 585
R74 B.n212 B.n125 585
R75 B.n211 B.n210 585
R76 B.n209 B.n126 585
R77 B.n208 B.n207 585
R78 B.n206 B.n127 585
R79 B.n205 B.n204 585
R80 B.n203 B.n128 585
R81 B.n202 B.n201 585
R82 B.n200 B.n129 585
R83 B.n199 B.n198 585
R84 B.n197 B.n130 585
R85 B.n196 B.n195 585
R86 B.n194 B.n131 585
R87 B.n193 B.n192 585
R88 B.n191 B.n132 585
R89 B.n190 B.n189 585
R90 B.n188 B.n133 585
R91 B.n187 B.n186 585
R92 B.n185 B.n134 585
R93 B.n184 B.n183 585
R94 B.n182 B.n135 585
R95 B.n181 B.n180 585
R96 B.n179 B.n136 585
R97 B.n178 B.n177 585
R98 B.n176 B.n137 585
R99 B.n175 B.n174 585
R100 B.n329 B.n328 585
R101 B.n330 B.n85 585
R102 B.n332 B.n331 585
R103 B.n333 B.n84 585
R104 B.n335 B.n334 585
R105 B.n336 B.n83 585
R106 B.n338 B.n337 585
R107 B.n339 B.n82 585
R108 B.n341 B.n340 585
R109 B.n342 B.n81 585
R110 B.n344 B.n343 585
R111 B.n345 B.n80 585
R112 B.n347 B.n346 585
R113 B.n348 B.n79 585
R114 B.n350 B.n349 585
R115 B.n351 B.n78 585
R116 B.n353 B.n352 585
R117 B.n354 B.n77 585
R118 B.n356 B.n355 585
R119 B.n357 B.n76 585
R120 B.n359 B.n358 585
R121 B.n360 B.n75 585
R122 B.n362 B.n361 585
R123 B.n363 B.n74 585
R124 B.n365 B.n364 585
R125 B.n366 B.n73 585
R126 B.n368 B.n367 585
R127 B.n369 B.n72 585
R128 B.n371 B.n370 585
R129 B.n372 B.n71 585
R130 B.n374 B.n373 585
R131 B.n375 B.n70 585
R132 B.n377 B.n376 585
R133 B.n378 B.n69 585
R134 B.n380 B.n379 585
R135 B.n381 B.n68 585
R136 B.n383 B.n382 585
R137 B.n384 B.n67 585
R138 B.n386 B.n385 585
R139 B.n387 B.n66 585
R140 B.n539 B.n538 585
R141 B.n537 B.n12 585
R142 B.n536 B.n535 585
R143 B.n534 B.n13 585
R144 B.n533 B.n532 585
R145 B.n531 B.n14 585
R146 B.n530 B.n529 585
R147 B.n528 B.n15 585
R148 B.n527 B.n526 585
R149 B.n525 B.n16 585
R150 B.n524 B.n523 585
R151 B.n522 B.n17 585
R152 B.n521 B.n520 585
R153 B.n519 B.n18 585
R154 B.n518 B.n517 585
R155 B.n516 B.n19 585
R156 B.n515 B.n514 585
R157 B.n513 B.n20 585
R158 B.n512 B.n511 585
R159 B.n510 B.n21 585
R160 B.n509 B.n508 585
R161 B.n507 B.n22 585
R162 B.n506 B.n505 585
R163 B.n504 B.n23 585
R164 B.n503 B.n502 585
R165 B.n501 B.n24 585
R166 B.n500 B.n499 585
R167 B.n498 B.n25 585
R168 B.n497 B.n496 585
R169 B.n495 B.n26 585
R170 B.n494 B.n493 585
R171 B.n492 B.n27 585
R172 B.n491 B.n490 585
R173 B.n489 B.n28 585
R174 B.n488 B.n487 585
R175 B.n486 B.n29 585
R176 B.n485 B.n484 585
R177 B.n483 B.n30 585
R178 B.n482 B.n481 585
R179 B.n480 B.n31 585
R180 B.n479 B.n478 585
R181 B.n477 B.n32 585
R182 B.n476 B.n475 585
R183 B.n474 B.n33 585
R184 B.n473 B.n472 585
R185 B.n471 B.n470 585
R186 B.n469 B.n37 585
R187 B.n468 B.n467 585
R188 B.n466 B.n38 585
R189 B.n465 B.n464 585
R190 B.n463 B.n39 585
R191 B.n462 B.n461 585
R192 B.n460 B.n40 585
R193 B.n459 B.n458 585
R194 B.n457 B.n41 585
R195 B.n455 B.n454 585
R196 B.n453 B.n44 585
R197 B.n452 B.n451 585
R198 B.n450 B.n45 585
R199 B.n449 B.n448 585
R200 B.n447 B.n46 585
R201 B.n446 B.n445 585
R202 B.n444 B.n47 585
R203 B.n443 B.n442 585
R204 B.n441 B.n48 585
R205 B.n440 B.n439 585
R206 B.n438 B.n49 585
R207 B.n437 B.n436 585
R208 B.n435 B.n50 585
R209 B.n434 B.n433 585
R210 B.n432 B.n51 585
R211 B.n431 B.n430 585
R212 B.n429 B.n52 585
R213 B.n428 B.n427 585
R214 B.n426 B.n53 585
R215 B.n425 B.n424 585
R216 B.n423 B.n54 585
R217 B.n422 B.n421 585
R218 B.n420 B.n55 585
R219 B.n419 B.n418 585
R220 B.n417 B.n56 585
R221 B.n416 B.n415 585
R222 B.n414 B.n57 585
R223 B.n413 B.n412 585
R224 B.n411 B.n58 585
R225 B.n410 B.n409 585
R226 B.n408 B.n59 585
R227 B.n407 B.n406 585
R228 B.n405 B.n60 585
R229 B.n404 B.n403 585
R230 B.n402 B.n61 585
R231 B.n401 B.n400 585
R232 B.n399 B.n62 585
R233 B.n398 B.n397 585
R234 B.n396 B.n63 585
R235 B.n395 B.n394 585
R236 B.n393 B.n64 585
R237 B.n392 B.n391 585
R238 B.n390 B.n65 585
R239 B.n389 B.n388 585
R240 B.n540 B.n11 585
R241 B.n542 B.n541 585
R242 B.n543 B.n10 585
R243 B.n545 B.n544 585
R244 B.n546 B.n9 585
R245 B.n548 B.n547 585
R246 B.n549 B.n8 585
R247 B.n551 B.n550 585
R248 B.n552 B.n7 585
R249 B.n554 B.n553 585
R250 B.n555 B.n6 585
R251 B.n557 B.n556 585
R252 B.n558 B.n5 585
R253 B.n560 B.n559 585
R254 B.n561 B.n4 585
R255 B.n563 B.n562 585
R256 B.n564 B.n3 585
R257 B.n566 B.n565 585
R258 B.n567 B.n0 585
R259 B.n2 B.n1 585
R260 B.n148 B.n147 585
R261 B.n149 B.n146 585
R262 B.n151 B.n150 585
R263 B.n152 B.n145 585
R264 B.n154 B.n153 585
R265 B.n155 B.n144 585
R266 B.n157 B.n156 585
R267 B.n158 B.n143 585
R268 B.n160 B.n159 585
R269 B.n161 B.n142 585
R270 B.n163 B.n162 585
R271 B.n164 B.n141 585
R272 B.n166 B.n165 585
R273 B.n167 B.n140 585
R274 B.n169 B.n168 585
R275 B.n170 B.n139 585
R276 B.n172 B.n171 585
R277 B.n173 B.n138 585
R278 B.n114 B.t9 539.644
R279 B.n256 B.t0 539.644
R280 B.n42 B.t6 539.644
R281 B.n34 B.t3 539.644
R282 B.n174 B.n173 434.841
R283 B.n328 B.n327 434.841
R284 B.n388 B.n387 434.841
R285 B.n538 B.n11 434.841
R286 B.n569 B.n568 256.663
R287 B.n568 B.n567 235.042
R288 B.n568 B.n2 235.042
R289 B.n174 B.n137 163.367
R290 B.n178 B.n137 163.367
R291 B.n179 B.n178 163.367
R292 B.n180 B.n179 163.367
R293 B.n180 B.n135 163.367
R294 B.n184 B.n135 163.367
R295 B.n185 B.n184 163.367
R296 B.n186 B.n185 163.367
R297 B.n186 B.n133 163.367
R298 B.n190 B.n133 163.367
R299 B.n191 B.n190 163.367
R300 B.n192 B.n191 163.367
R301 B.n192 B.n131 163.367
R302 B.n196 B.n131 163.367
R303 B.n197 B.n196 163.367
R304 B.n198 B.n197 163.367
R305 B.n198 B.n129 163.367
R306 B.n202 B.n129 163.367
R307 B.n203 B.n202 163.367
R308 B.n204 B.n203 163.367
R309 B.n204 B.n127 163.367
R310 B.n208 B.n127 163.367
R311 B.n209 B.n208 163.367
R312 B.n210 B.n209 163.367
R313 B.n210 B.n125 163.367
R314 B.n214 B.n125 163.367
R315 B.n215 B.n214 163.367
R316 B.n216 B.n215 163.367
R317 B.n216 B.n123 163.367
R318 B.n220 B.n123 163.367
R319 B.n221 B.n220 163.367
R320 B.n222 B.n221 163.367
R321 B.n222 B.n121 163.367
R322 B.n226 B.n121 163.367
R323 B.n227 B.n226 163.367
R324 B.n228 B.n227 163.367
R325 B.n228 B.n119 163.367
R326 B.n232 B.n119 163.367
R327 B.n233 B.n232 163.367
R328 B.n234 B.n233 163.367
R329 B.n234 B.n117 163.367
R330 B.n238 B.n117 163.367
R331 B.n239 B.n238 163.367
R332 B.n240 B.n239 163.367
R333 B.n240 B.n113 163.367
R334 B.n245 B.n113 163.367
R335 B.n246 B.n245 163.367
R336 B.n247 B.n246 163.367
R337 B.n247 B.n111 163.367
R338 B.n251 B.n111 163.367
R339 B.n252 B.n251 163.367
R340 B.n253 B.n252 163.367
R341 B.n253 B.n109 163.367
R342 B.n260 B.n109 163.367
R343 B.n261 B.n260 163.367
R344 B.n262 B.n261 163.367
R345 B.n262 B.n107 163.367
R346 B.n266 B.n107 163.367
R347 B.n267 B.n266 163.367
R348 B.n268 B.n267 163.367
R349 B.n268 B.n105 163.367
R350 B.n272 B.n105 163.367
R351 B.n273 B.n272 163.367
R352 B.n274 B.n273 163.367
R353 B.n274 B.n103 163.367
R354 B.n278 B.n103 163.367
R355 B.n279 B.n278 163.367
R356 B.n280 B.n279 163.367
R357 B.n280 B.n101 163.367
R358 B.n284 B.n101 163.367
R359 B.n285 B.n284 163.367
R360 B.n286 B.n285 163.367
R361 B.n286 B.n99 163.367
R362 B.n290 B.n99 163.367
R363 B.n291 B.n290 163.367
R364 B.n292 B.n291 163.367
R365 B.n292 B.n97 163.367
R366 B.n296 B.n97 163.367
R367 B.n297 B.n296 163.367
R368 B.n298 B.n297 163.367
R369 B.n298 B.n95 163.367
R370 B.n302 B.n95 163.367
R371 B.n303 B.n302 163.367
R372 B.n304 B.n303 163.367
R373 B.n304 B.n93 163.367
R374 B.n308 B.n93 163.367
R375 B.n309 B.n308 163.367
R376 B.n310 B.n309 163.367
R377 B.n310 B.n91 163.367
R378 B.n314 B.n91 163.367
R379 B.n315 B.n314 163.367
R380 B.n316 B.n315 163.367
R381 B.n316 B.n89 163.367
R382 B.n320 B.n89 163.367
R383 B.n321 B.n320 163.367
R384 B.n322 B.n321 163.367
R385 B.n322 B.n87 163.367
R386 B.n326 B.n87 163.367
R387 B.n327 B.n326 163.367
R388 B.n387 B.n386 163.367
R389 B.n386 B.n67 163.367
R390 B.n382 B.n67 163.367
R391 B.n382 B.n381 163.367
R392 B.n381 B.n380 163.367
R393 B.n380 B.n69 163.367
R394 B.n376 B.n69 163.367
R395 B.n376 B.n375 163.367
R396 B.n375 B.n374 163.367
R397 B.n374 B.n71 163.367
R398 B.n370 B.n71 163.367
R399 B.n370 B.n369 163.367
R400 B.n369 B.n368 163.367
R401 B.n368 B.n73 163.367
R402 B.n364 B.n73 163.367
R403 B.n364 B.n363 163.367
R404 B.n363 B.n362 163.367
R405 B.n362 B.n75 163.367
R406 B.n358 B.n75 163.367
R407 B.n358 B.n357 163.367
R408 B.n357 B.n356 163.367
R409 B.n356 B.n77 163.367
R410 B.n352 B.n77 163.367
R411 B.n352 B.n351 163.367
R412 B.n351 B.n350 163.367
R413 B.n350 B.n79 163.367
R414 B.n346 B.n79 163.367
R415 B.n346 B.n345 163.367
R416 B.n345 B.n344 163.367
R417 B.n344 B.n81 163.367
R418 B.n340 B.n81 163.367
R419 B.n340 B.n339 163.367
R420 B.n339 B.n338 163.367
R421 B.n338 B.n83 163.367
R422 B.n334 B.n83 163.367
R423 B.n334 B.n333 163.367
R424 B.n333 B.n332 163.367
R425 B.n332 B.n85 163.367
R426 B.n328 B.n85 163.367
R427 B.n538 B.n537 163.367
R428 B.n537 B.n536 163.367
R429 B.n536 B.n13 163.367
R430 B.n532 B.n13 163.367
R431 B.n532 B.n531 163.367
R432 B.n531 B.n530 163.367
R433 B.n530 B.n15 163.367
R434 B.n526 B.n15 163.367
R435 B.n526 B.n525 163.367
R436 B.n525 B.n524 163.367
R437 B.n524 B.n17 163.367
R438 B.n520 B.n17 163.367
R439 B.n520 B.n519 163.367
R440 B.n519 B.n518 163.367
R441 B.n518 B.n19 163.367
R442 B.n514 B.n19 163.367
R443 B.n514 B.n513 163.367
R444 B.n513 B.n512 163.367
R445 B.n512 B.n21 163.367
R446 B.n508 B.n21 163.367
R447 B.n508 B.n507 163.367
R448 B.n507 B.n506 163.367
R449 B.n506 B.n23 163.367
R450 B.n502 B.n23 163.367
R451 B.n502 B.n501 163.367
R452 B.n501 B.n500 163.367
R453 B.n500 B.n25 163.367
R454 B.n496 B.n25 163.367
R455 B.n496 B.n495 163.367
R456 B.n495 B.n494 163.367
R457 B.n494 B.n27 163.367
R458 B.n490 B.n27 163.367
R459 B.n490 B.n489 163.367
R460 B.n489 B.n488 163.367
R461 B.n488 B.n29 163.367
R462 B.n484 B.n29 163.367
R463 B.n484 B.n483 163.367
R464 B.n483 B.n482 163.367
R465 B.n482 B.n31 163.367
R466 B.n478 B.n31 163.367
R467 B.n478 B.n477 163.367
R468 B.n477 B.n476 163.367
R469 B.n476 B.n33 163.367
R470 B.n472 B.n33 163.367
R471 B.n472 B.n471 163.367
R472 B.n471 B.n37 163.367
R473 B.n467 B.n37 163.367
R474 B.n467 B.n466 163.367
R475 B.n466 B.n465 163.367
R476 B.n465 B.n39 163.367
R477 B.n461 B.n39 163.367
R478 B.n461 B.n460 163.367
R479 B.n460 B.n459 163.367
R480 B.n459 B.n41 163.367
R481 B.n454 B.n41 163.367
R482 B.n454 B.n453 163.367
R483 B.n453 B.n452 163.367
R484 B.n452 B.n45 163.367
R485 B.n448 B.n45 163.367
R486 B.n448 B.n447 163.367
R487 B.n447 B.n446 163.367
R488 B.n446 B.n47 163.367
R489 B.n442 B.n47 163.367
R490 B.n442 B.n441 163.367
R491 B.n441 B.n440 163.367
R492 B.n440 B.n49 163.367
R493 B.n436 B.n49 163.367
R494 B.n436 B.n435 163.367
R495 B.n435 B.n434 163.367
R496 B.n434 B.n51 163.367
R497 B.n430 B.n51 163.367
R498 B.n430 B.n429 163.367
R499 B.n429 B.n428 163.367
R500 B.n428 B.n53 163.367
R501 B.n424 B.n53 163.367
R502 B.n424 B.n423 163.367
R503 B.n423 B.n422 163.367
R504 B.n422 B.n55 163.367
R505 B.n418 B.n55 163.367
R506 B.n418 B.n417 163.367
R507 B.n417 B.n416 163.367
R508 B.n416 B.n57 163.367
R509 B.n412 B.n57 163.367
R510 B.n412 B.n411 163.367
R511 B.n411 B.n410 163.367
R512 B.n410 B.n59 163.367
R513 B.n406 B.n59 163.367
R514 B.n406 B.n405 163.367
R515 B.n405 B.n404 163.367
R516 B.n404 B.n61 163.367
R517 B.n400 B.n61 163.367
R518 B.n400 B.n399 163.367
R519 B.n399 B.n398 163.367
R520 B.n398 B.n63 163.367
R521 B.n394 B.n63 163.367
R522 B.n394 B.n393 163.367
R523 B.n393 B.n392 163.367
R524 B.n392 B.n65 163.367
R525 B.n388 B.n65 163.367
R526 B.n542 B.n11 163.367
R527 B.n543 B.n542 163.367
R528 B.n544 B.n543 163.367
R529 B.n544 B.n9 163.367
R530 B.n548 B.n9 163.367
R531 B.n549 B.n548 163.367
R532 B.n550 B.n549 163.367
R533 B.n550 B.n7 163.367
R534 B.n554 B.n7 163.367
R535 B.n555 B.n554 163.367
R536 B.n556 B.n555 163.367
R537 B.n556 B.n5 163.367
R538 B.n560 B.n5 163.367
R539 B.n561 B.n560 163.367
R540 B.n562 B.n561 163.367
R541 B.n562 B.n3 163.367
R542 B.n566 B.n3 163.367
R543 B.n567 B.n566 163.367
R544 B.n148 B.n2 163.367
R545 B.n149 B.n148 163.367
R546 B.n150 B.n149 163.367
R547 B.n150 B.n145 163.367
R548 B.n154 B.n145 163.367
R549 B.n155 B.n154 163.367
R550 B.n156 B.n155 163.367
R551 B.n156 B.n143 163.367
R552 B.n160 B.n143 163.367
R553 B.n161 B.n160 163.367
R554 B.n162 B.n161 163.367
R555 B.n162 B.n141 163.367
R556 B.n166 B.n141 163.367
R557 B.n167 B.n166 163.367
R558 B.n168 B.n167 163.367
R559 B.n168 B.n139 163.367
R560 B.n172 B.n139 163.367
R561 B.n173 B.n172 163.367
R562 B.n256 B.t1 135.957
R563 B.n42 B.t8 135.957
R564 B.n114 B.t10 135.94
R565 B.n34 B.t5 135.94
R566 B.n257 B.t2 111.326
R567 B.n43 B.t7 111.326
R568 B.n115 B.t11 111.311
R569 B.n35 B.t4 111.311
R570 B.n242 B.n115 59.5399
R571 B.n258 B.n257 59.5399
R572 B.n456 B.n43 59.5399
R573 B.n36 B.n35 59.5399
R574 B.n540 B.n539 28.2542
R575 B.n389 B.n66 28.2542
R576 B.n329 B.n86 28.2542
R577 B.n175 B.n138 28.2542
R578 B.n115 B.n114 24.6308
R579 B.n257 B.n256 24.6308
R580 B.n43 B.n42 24.6308
R581 B.n35 B.n34 24.6308
R582 B B.n569 18.0485
R583 B.n541 B.n540 10.6151
R584 B.n541 B.n10 10.6151
R585 B.n545 B.n10 10.6151
R586 B.n546 B.n545 10.6151
R587 B.n547 B.n546 10.6151
R588 B.n547 B.n8 10.6151
R589 B.n551 B.n8 10.6151
R590 B.n552 B.n551 10.6151
R591 B.n553 B.n552 10.6151
R592 B.n553 B.n6 10.6151
R593 B.n557 B.n6 10.6151
R594 B.n558 B.n557 10.6151
R595 B.n559 B.n558 10.6151
R596 B.n559 B.n4 10.6151
R597 B.n563 B.n4 10.6151
R598 B.n564 B.n563 10.6151
R599 B.n565 B.n564 10.6151
R600 B.n565 B.n0 10.6151
R601 B.n539 B.n12 10.6151
R602 B.n535 B.n12 10.6151
R603 B.n535 B.n534 10.6151
R604 B.n534 B.n533 10.6151
R605 B.n533 B.n14 10.6151
R606 B.n529 B.n14 10.6151
R607 B.n529 B.n528 10.6151
R608 B.n528 B.n527 10.6151
R609 B.n527 B.n16 10.6151
R610 B.n523 B.n16 10.6151
R611 B.n523 B.n522 10.6151
R612 B.n522 B.n521 10.6151
R613 B.n521 B.n18 10.6151
R614 B.n517 B.n18 10.6151
R615 B.n517 B.n516 10.6151
R616 B.n516 B.n515 10.6151
R617 B.n515 B.n20 10.6151
R618 B.n511 B.n20 10.6151
R619 B.n511 B.n510 10.6151
R620 B.n510 B.n509 10.6151
R621 B.n509 B.n22 10.6151
R622 B.n505 B.n22 10.6151
R623 B.n505 B.n504 10.6151
R624 B.n504 B.n503 10.6151
R625 B.n503 B.n24 10.6151
R626 B.n499 B.n24 10.6151
R627 B.n499 B.n498 10.6151
R628 B.n498 B.n497 10.6151
R629 B.n497 B.n26 10.6151
R630 B.n493 B.n26 10.6151
R631 B.n493 B.n492 10.6151
R632 B.n492 B.n491 10.6151
R633 B.n491 B.n28 10.6151
R634 B.n487 B.n28 10.6151
R635 B.n487 B.n486 10.6151
R636 B.n486 B.n485 10.6151
R637 B.n485 B.n30 10.6151
R638 B.n481 B.n30 10.6151
R639 B.n481 B.n480 10.6151
R640 B.n480 B.n479 10.6151
R641 B.n479 B.n32 10.6151
R642 B.n475 B.n32 10.6151
R643 B.n475 B.n474 10.6151
R644 B.n474 B.n473 10.6151
R645 B.n470 B.n469 10.6151
R646 B.n469 B.n468 10.6151
R647 B.n468 B.n38 10.6151
R648 B.n464 B.n38 10.6151
R649 B.n464 B.n463 10.6151
R650 B.n463 B.n462 10.6151
R651 B.n462 B.n40 10.6151
R652 B.n458 B.n40 10.6151
R653 B.n458 B.n457 10.6151
R654 B.n455 B.n44 10.6151
R655 B.n451 B.n44 10.6151
R656 B.n451 B.n450 10.6151
R657 B.n450 B.n449 10.6151
R658 B.n449 B.n46 10.6151
R659 B.n445 B.n46 10.6151
R660 B.n445 B.n444 10.6151
R661 B.n444 B.n443 10.6151
R662 B.n443 B.n48 10.6151
R663 B.n439 B.n48 10.6151
R664 B.n439 B.n438 10.6151
R665 B.n438 B.n437 10.6151
R666 B.n437 B.n50 10.6151
R667 B.n433 B.n50 10.6151
R668 B.n433 B.n432 10.6151
R669 B.n432 B.n431 10.6151
R670 B.n431 B.n52 10.6151
R671 B.n427 B.n52 10.6151
R672 B.n427 B.n426 10.6151
R673 B.n426 B.n425 10.6151
R674 B.n425 B.n54 10.6151
R675 B.n421 B.n54 10.6151
R676 B.n421 B.n420 10.6151
R677 B.n420 B.n419 10.6151
R678 B.n419 B.n56 10.6151
R679 B.n415 B.n56 10.6151
R680 B.n415 B.n414 10.6151
R681 B.n414 B.n413 10.6151
R682 B.n413 B.n58 10.6151
R683 B.n409 B.n58 10.6151
R684 B.n409 B.n408 10.6151
R685 B.n408 B.n407 10.6151
R686 B.n407 B.n60 10.6151
R687 B.n403 B.n60 10.6151
R688 B.n403 B.n402 10.6151
R689 B.n402 B.n401 10.6151
R690 B.n401 B.n62 10.6151
R691 B.n397 B.n62 10.6151
R692 B.n397 B.n396 10.6151
R693 B.n396 B.n395 10.6151
R694 B.n395 B.n64 10.6151
R695 B.n391 B.n64 10.6151
R696 B.n391 B.n390 10.6151
R697 B.n390 B.n389 10.6151
R698 B.n385 B.n66 10.6151
R699 B.n385 B.n384 10.6151
R700 B.n384 B.n383 10.6151
R701 B.n383 B.n68 10.6151
R702 B.n379 B.n68 10.6151
R703 B.n379 B.n378 10.6151
R704 B.n378 B.n377 10.6151
R705 B.n377 B.n70 10.6151
R706 B.n373 B.n70 10.6151
R707 B.n373 B.n372 10.6151
R708 B.n372 B.n371 10.6151
R709 B.n371 B.n72 10.6151
R710 B.n367 B.n72 10.6151
R711 B.n367 B.n366 10.6151
R712 B.n366 B.n365 10.6151
R713 B.n365 B.n74 10.6151
R714 B.n361 B.n74 10.6151
R715 B.n361 B.n360 10.6151
R716 B.n360 B.n359 10.6151
R717 B.n359 B.n76 10.6151
R718 B.n355 B.n76 10.6151
R719 B.n355 B.n354 10.6151
R720 B.n354 B.n353 10.6151
R721 B.n353 B.n78 10.6151
R722 B.n349 B.n78 10.6151
R723 B.n349 B.n348 10.6151
R724 B.n348 B.n347 10.6151
R725 B.n347 B.n80 10.6151
R726 B.n343 B.n80 10.6151
R727 B.n343 B.n342 10.6151
R728 B.n342 B.n341 10.6151
R729 B.n341 B.n82 10.6151
R730 B.n337 B.n82 10.6151
R731 B.n337 B.n336 10.6151
R732 B.n336 B.n335 10.6151
R733 B.n335 B.n84 10.6151
R734 B.n331 B.n84 10.6151
R735 B.n331 B.n330 10.6151
R736 B.n330 B.n329 10.6151
R737 B.n147 B.n1 10.6151
R738 B.n147 B.n146 10.6151
R739 B.n151 B.n146 10.6151
R740 B.n152 B.n151 10.6151
R741 B.n153 B.n152 10.6151
R742 B.n153 B.n144 10.6151
R743 B.n157 B.n144 10.6151
R744 B.n158 B.n157 10.6151
R745 B.n159 B.n158 10.6151
R746 B.n159 B.n142 10.6151
R747 B.n163 B.n142 10.6151
R748 B.n164 B.n163 10.6151
R749 B.n165 B.n164 10.6151
R750 B.n165 B.n140 10.6151
R751 B.n169 B.n140 10.6151
R752 B.n170 B.n169 10.6151
R753 B.n171 B.n170 10.6151
R754 B.n171 B.n138 10.6151
R755 B.n176 B.n175 10.6151
R756 B.n177 B.n176 10.6151
R757 B.n177 B.n136 10.6151
R758 B.n181 B.n136 10.6151
R759 B.n182 B.n181 10.6151
R760 B.n183 B.n182 10.6151
R761 B.n183 B.n134 10.6151
R762 B.n187 B.n134 10.6151
R763 B.n188 B.n187 10.6151
R764 B.n189 B.n188 10.6151
R765 B.n189 B.n132 10.6151
R766 B.n193 B.n132 10.6151
R767 B.n194 B.n193 10.6151
R768 B.n195 B.n194 10.6151
R769 B.n195 B.n130 10.6151
R770 B.n199 B.n130 10.6151
R771 B.n200 B.n199 10.6151
R772 B.n201 B.n200 10.6151
R773 B.n201 B.n128 10.6151
R774 B.n205 B.n128 10.6151
R775 B.n206 B.n205 10.6151
R776 B.n207 B.n206 10.6151
R777 B.n207 B.n126 10.6151
R778 B.n211 B.n126 10.6151
R779 B.n212 B.n211 10.6151
R780 B.n213 B.n212 10.6151
R781 B.n213 B.n124 10.6151
R782 B.n217 B.n124 10.6151
R783 B.n218 B.n217 10.6151
R784 B.n219 B.n218 10.6151
R785 B.n219 B.n122 10.6151
R786 B.n223 B.n122 10.6151
R787 B.n224 B.n223 10.6151
R788 B.n225 B.n224 10.6151
R789 B.n225 B.n120 10.6151
R790 B.n229 B.n120 10.6151
R791 B.n230 B.n229 10.6151
R792 B.n231 B.n230 10.6151
R793 B.n231 B.n118 10.6151
R794 B.n235 B.n118 10.6151
R795 B.n236 B.n235 10.6151
R796 B.n237 B.n236 10.6151
R797 B.n237 B.n116 10.6151
R798 B.n241 B.n116 10.6151
R799 B.n244 B.n243 10.6151
R800 B.n244 B.n112 10.6151
R801 B.n248 B.n112 10.6151
R802 B.n249 B.n248 10.6151
R803 B.n250 B.n249 10.6151
R804 B.n250 B.n110 10.6151
R805 B.n254 B.n110 10.6151
R806 B.n255 B.n254 10.6151
R807 B.n259 B.n255 10.6151
R808 B.n263 B.n108 10.6151
R809 B.n264 B.n263 10.6151
R810 B.n265 B.n264 10.6151
R811 B.n265 B.n106 10.6151
R812 B.n269 B.n106 10.6151
R813 B.n270 B.n269 10.6151
R814 B.n271 B.n270 10.6151
R815 B.n271 B.n104 10.6151
R816 B.n275 B.n104 10.6151
R817 B.n276 B.n275 10.6151
R818 B.n277 B.n276 10.6151
R819 B.n277 B.n102 10.6151
R820 B.n281 B.n102 10.6151
R821 B.n282 B.n281 10.6151
R822 B.n283 B.n282 10.6151
R823 B.n283 B.n100 10.6151
R824 B.n287 B.n100 10.6151
R825 B.n288 B.n287 10.6151
R826 B.n289 B.n288 10.6151
R827 B.n289 B.n98 10.6151
R828 B.n293 B.n98 10.6151
R829 B.n294 B.n293 10.6151
R830 B.n295 B.n294 10.6151
R831 B.n295 B.n96 10.6151
R832 B.n299 B.n96 10.6151
R833 B.n300 B.n299 10.6151
R834 B.n301 B.n300 10.6151
R835 B.n301 B.n94 10.6151
R836 B.n305 B.n94 10.6151
R837 B.n306 B.n305 10.6151
R838 B.n307 B.n306 10.6151
R839 B.n307 B.n92 10.6151
R840 B.n311 B.n92 10.6151
R841 B.n312 B.n311 10.6151
R842 B.n313 B.n312 10.6151
R843 B.n313 B.n90 10.6151
R844 B.n317 B.n90 10.6151
R845 B.n318 B.n317 10.6151
R846 B.n319 B.n318 10.6151
R847 B.n319 B.n88 10.6151
R848 B.n323 B.n88 10.6151
R849 B.n324 B.n323 10.6151
R850 B.n325 B.n324 10.6151
R851 B.n325 B.n86 10.6151
R852 B.n473 B.n36 9.36635
R853 B.n456 B.n455 9.36635
R854 B.n242 B.n241 9.36635
R855 B.n258 B.n108 9.36635
R856 B.n569 B.n0 8.11757
R857 B.n569 B.n1 8.11757
R858 B.n470 B.n36 1.24928
R859 B.n457 B.n456 1.24928
R860 B.n243 B.n242 1.24928
R861 B.n259 B.n258 1.24928
R862 VN.n0 VN.t0 397.798
R863 VN.n1 VN.t3 397.798
R864 VN.n1 VN.t1 397.711
R865 VN.n0 VN.t2 397.711
R866 VN VN.n1 73.5917
R867 VN VN.n0 31.2622
R868 VDD2.n2 VDD2.n0 110.001
R869 VDD2.n2 VDD2.n1 71.6648
R870 VDD2.n1 VDD2.t0 2.47236
R871 VDD2.n1 VDD2.t2 2.47236
R872 VDD2.n0 VDD2.t1 2.47236
R873 VDD2.n0 VDD2.t3 2.47236
R874 VDD2 VDD2.n2 0.0586897
R875 VTAIL.n5 VTAIL.t1 57.4581
R876 VTAIL.n4 VTAIL.t3 57.4581
R877 VTAIL.n3 VTAIL.t5 57.4581
R878 VTAIL.n7 VTAIL.t4 57.4578
R879 VTAIL.n0 VTAIL.t6 57.4578
R880 VTAIL.n1 VTAIL.t0 57.4578
R881 VTAIL.n2 VTAIL.t7 57.4578
R882 VTAIL.n6 VTAIL.t2 57.4578
R883 VTAIL.n7 VTAIL.n6 24.7979
R884 VTAIL.n3 VTAIL.n2 24.7979
R885 VTAIL.n4 VTAIL.n3 1.09533
R886 VTAIL.n6 VTAIL.n5 1.09533
R887 VTAIL.n2 VTAIL.n1 1.09533
R888 VTAIL VTAIL.n0 0.606103
R889 VTAIL VTAIL.n7 0.489724
R890 VTAIL.n5 VTAIL.n4 0.470328
R891 VTAIL.n1 VTAIL.n0 0.470328
R892 VP.n0 VP.t2 397.798
R893 VP.n0 VP.t1 397.711
R894 VP.n2 VP.t0 379.19
R895 VP.n3 VP.t3 379.19
R896 VP.n4 VP.n3 80.6037
R897 VP.n2 VP.n1 80.6037
R898 VP.n1 VP.n0 73.3062
R899 VP.n3 VP.n2 48.2005
R900 VP.n4 VP.n1 0.380177
R901 VP VP.n4 0.146778
R902 VDD1 VDD1.n1 110.525
R903 VDD1 VDD1.n0 71.723
R904 VDD1.n0 VDD1.t1 2.47236
R905 VDD1.n0 VDD1.t2 2.47236
R906 VDD1.n1 VDD1.t3 2.47236
R907 VDD1.n1 VDD1.t0 2.47236
C0 VTAIL VDD2 6.6417f
C1 VTAIL VN 3.49433f
C2 VN VDD2 3.88626f
C3 VDD1 VP 4.02712f
C4 B VP 1.16114f
C5 VDD1 B 0.999711f
C6 w_n1732_n3598# VP 2.87158f
C7 VDD1 w_n1732_n3598# 1.15038f
C8 w_n1732_n3598# B 7.52554f
C9 VTAIL VP 3.50844f
C10 VDD1 VTAIL 6.59862f
C11 VDD2 VP 0.288787f
C12 VDD1 VDD2 0.624375f
C13 VTAIL B 4.32296f
C14 VDD2 B 1.02486f
C15 VN VP 5.21036f
C16 VTAIL w_n1732_n3598# 4.36704f
C17 VDD1 VN 0.14761f
C18 w_n1732_n3598# VDD2 1.16983f
C19 VN B 0.806349f
C20 w_n1732_n3598# VN 2.65312f
C21 VDD2 VSUBS 0.734139f
C22 VDD1 VSUBS 5.133701f
C23 VTAIL VSUBS 0.978833f
C24 VN VSUBS 5.58331f
C25 VP VSUBS 1.480861f
C26 B VSUBS 2.933125f
C27 w_n1732_n3598# VSUBS 76.589f
C28 VDD1.t1 VSUBS 0.28356f
C29 VDD1.t2 VSUBS 0.28356f
C30 VDD1.n0 VSUBS 2.242f
C31 VDD1.t3 VSUBS 0.28356f
C32 VDD1.t0 VSUBS 0.28356f
C33 VDD1.n1 VSUBS 2.95315f
C34 VP.t1 VSUBS 1.95697f
C35 VP.t2 VSUBS 1.95716f
C36 VP.n0 VSUBS 2.83378f
C37 VP.n1 VSUBS 3.38352f
C38 VP.t0 VSUBS 1.92185f
C39 VP.n2 VSUBS 0.754316f
C40 VP.t3 VSUBS 1.92185f
C41 VP.n3 VSUBS 0.754316f
C42 VP.n4 VSUBS 0.069383f
C43 VTAIL.t6 VSUBS 2.2792f
C44 VTAIL.n0 VSUBS 0.707329f
C45 VTAIL.t0 VSUBS 2.2792f
C46 VTAIL.n1 VSUBS 0.743031f
C47 VTAIL.t7 VSUBS 2.2792f
C48 VTAIL.n2 VSUBS 1.92356f
C49 VTAIL.t5 VSUBS 2.27921f
C50 VTAIL.n3 VSUBS 1.92356f
C51 VTAIL.t3 VSUBS 2.27921f
C52 VTAIL.n4 VSUBS 0.743023f
C53 VTAIL.t1 VSUBS 2.27921f
C54 VTAIL.n5 VSUBS 0.743023f
C55 VTAIL.t2 VSUBS 2.2792f
C56 VTAIL.n6 VSUBS 1.92356f
C57 VTAIL.t4 VSUBS 2.2792f
C58 VTAIL.n7 VSUBS 1.87937f
C59 VDD2.t1 VSUBS 0.283582f
C60 VDD2.t3 VSUBS 0.283582f
C61 VDD2.n0 VSUBS 2.92792f
C62 VDD2.t0 VSUBS 0.283582f
C63 VDD2.t2 VSUBS 0.283582f
C64 VDD2.n1 VSUBS 2.24165f
C65 VDD2.n2 VSUBS 4.09396f
C66 VN.t0 VSUBS 1.91012f
C67 VN.t2 VSUBS 1.90994f
C68 VN.n0 VSUBS 1.40501f
C69 VN.t3 VSUBS 1.91012f
C70 VN.t1 VSUBS 1.90994f
C71 VN.n1 VSUBS 2.78681f
C72 B.n0 VSUBS 0.006877f
C73 B.n1 VSUBS 0.006877f
C74 B.n2 VSUBS 0.010171f
C75 B.n3 VSUBS 0.007794f
C76 B.n4 VSUBS 0.007794f
C77 B.n5 VSUBS 0.007794f
C78 B.n6 VSUBS 0.007794f
C79 B.n7 VSUBS 0.007794f
C80 B.n8 VSUBS 0.007794f
C81 B.n9 VSUBS 0.007794f
C82 B.n10 VSUBS 0.007794f
C83 B.n11 VSUBS 0.016088f
C84 B.n12 VSUBS 0.007794f
C85 B.n13 VSUBS 0.007794f
C86 B.n14 VSUBS 0.007794f
C87 B.n15 VSUBS 0.007794f
C88 B.n16 VSUBS 0.007794f
C89 B.n17 VSUBS 0.007794f
C90 B.n18 VSUBS 0.007794f
C91 B.n19 VSUBS 0.007794f
C92 B.n20 VSUBS 0.007794f
C93 B.n21 VSUBS 0.007794f
C94 B.n22 VSUBS 0.007794f
C95 B.n23 VSUBS 0.007794f
C96 B.n24 VSUBS 0.007794f
C97 B.n25 VSUBS 0.007794f
C98 B.n26 VSUBS 0.007794f
C99 B.n27 VSUBS 0.007794f
C100 B.n28 VSUBS 0.007794f
C101 B.n29 VSUBS 0.007794f
C102 B.n30 VSUBS 0.007794f
C103 B.n31 VSUBS 0.007794f
C104 B.n32 VSUBS 0.007794f
C105 B.n33 VSUBS 0.007794f
C106 B.t4 VSUBS 0.481654f
C107 B.t5 VSUBS 0.49275f
C108 B.t3 VSUBS 0.576639f
C109 B.n34 VSUBS 0.182448f
C110 B.n35 VSUBS 0.072359f
C111 B.n36 VSUBS 0.018058f
C112 B.n37 VSUBS 0.007794f
C113 B.n38 VSUBS 0.007794f
C114 B.n39 VSUBS 0.007794f
C115 B.n40 VSUBS 0.007794f
C116 B.n41 VSUBS 0.007794f
C117 B.t7 VSUBS 0.481643f
C118 B.t8 VSUBS 0.49274f
C119 B.t6 VSUBS 0.576639f
C120 B.n42 VSUBS 0.182458f
C121 B.n43 VSUBS 0.07237f
C122 B.n44 VSUBS 0.007794f
C123 B.n45 VSUBS 0.007794f
C124 B.n46 VSUBS 0.007794f
C125 B.n47 VSUBS 0.007794f
C126 B.n48 VSUBS 0.007794f
C127 B.n49 VSUBS 0.007794f
C128 B.n50 VSUBS 0.007794f
C129 B.n51 VSUBS 0.007794f
C130 B.n52 VSUBS 0.007794f
C131 B.n53 VSUBS 0.007794f
C132 B.n54 VSUBS 0.007794f
C133 B.n55 VSUBS 0.007794f
C134 B.n56 VSUBS 0.007794f
C135 B.n57 VSUBS 0.007794f
C136 B.n58 VSUBS 0.007794f
C137 B.n59 VSUBS 0.007794f
C138 B.n60 VSUBS 0.007794f
C139 B.n61 VSUBS 0.007794f
C140 B.n62 VSUBS 0.007794f
C141 B.n63 VSUBS 0.007794f
C142 B.n64 VSUBS 0.007794f
C143 B.n65 VSUBS 0.007794f
C144 B.n66 VSUBS 0.016088f
C145 B.n67 VSUBS 0.007794f
C146 B.n68 VSUBS 0.007794f
C147 B.n69 VSUBS 0.007794f
C148 B.n70 VSUBS 0.007794f
C149 B.n71 VSUBS 0.007794f
C150 B.n72 VSUBS 0.007794f
C151 B.n73 VSUBS 0.007794f
C152 B.n74 VSUBS 0.007794f
C153 B.n75 VSUBS 0.007794f
C154 B.n76 VSUBS 0.007794f
C155 B.n77 VSUBS 0.007794f
C156 B.n78 VSUBS 0.007794f
C157 B.n79 VSUBS 0.007794f
C158 B.n80 VSUBS 0.007794f
C159 B.n81 VSUBS 0.007794f
C160 B.n82 VSUBS 0.007794f
C161 B.n83 VSUBS 0.007794f
C162 B.n84 VSUBS 0.007794f
C163 B.n85 VSUBS 0.007794f
C164 B.n86 VSUBS 0.016088f
C165 B.n87 VSUBS 0.007794f
C166 B.n88 VSUBS 0.007794f
C167 B.n89 VSUBS 0.007794f
C168 B.n90 VSUBS 0.007794f
C169 B.n91 VSUBS 0.007794f
C170 B.n92 VSUBS 0.007794f
C171 B.n93 VSUBS 0.007794f
C172 B.n94 VSUBS 0.007794f
C173 B.n95 VSUBS 0.007794f
C174 B.n96 VSUBS 0.007794f
C175 B.n97 VSUBS 0.007794f
C176 B.n98 VSUBS 0.007794f
C177 B.n99 VSUBS 0.007794f
C178 B.n100 VSUBS 0.007794f
C179 B.n101 VSUBS 0.007794f
C180 B.n102 VSUBS 0.007794f
C181 B.n103 VSUBS 0.007794f
C182 B.n104 VSUBS 0.007794f
C183 B.n105 VSUBS 0.007794f
C184 B.n106 VSUBS 0.007794f
C185 B.n107 VSUBS 0.007794f
C186 B.n108 VSUBS 0.007336f
C187 B.n109 VSUBS 0.007794f
C188 B.n110 VSUBS 0.007794f
C189 B.n111 VSUBS 0.007794f
C190 B.n112 VSUBS 0.007794f
C191 B.n113 VSUBS 0.007794f
C192 B.t11 VSUBS 0.481654f
C193 B.t10 VSUBS 0.49275f
C194 B.t9 VSUBS 0.576639f
C195 B.n114 VSUBS 0.182448f
C196 B.n115 VSUBS 0.072359f
C197 B.n116 VSUBS 0.007794f
C198 B.n117 VSUBS 0.007794f
C199 B.n118 VSUBS 0.007794f
C200 B.n119 VSUBS 0.007794f
C201 B.n120 VSUBS 0.007794f
C202 B.n121 VSUBS 0.007794f
C203 B.n122 VSUBS 0.007794f
C204 B.n123 VSUBS 0.007794f
C205 B.n124 VSUBS 0.007794f
C206 B.n125 VSUBS 0.007794f
C207 B.n126 VSUBS 0.007794f
C208 B.n127 VSUBS 0.007794f
C209 B.n128 VSUBS 0.007794f
C210 B.n129 VSUBS 0.007794f
C211 B.n130 VSUBS 0.007794f
C212 B.n131 VSUBS 0.007794f
C213 B.n132 VSUBS 0.007794f
C214 B.n133 VSUBS 0.007794f
C215 B.n134 VSUBS 0.007794f
C216 B.n135 VSUBS 0.007794f
C217 B.n136 VSUBS 0.007794f
C218 B.n137 VSUBS 0.007794f
C219 B.n138 VSUBS 0.016088f
C220 B.n139 VSUBS 0.007794f
C221 B.n140 VSUBS 0.007794f
C222 B.n141 VSUBS 0.007794f
C223 B.n142 VSUBS 0.007794f
C224 B.n143 VSUBS 0.007794f
C225 B.n144 VSUBS 0.007794f
C226 B.n145 VSUBS 0.007794f
C227 B.n146 VSUBS 0.007794f
C228 B.n147 VSUBS 0.007794f
C229 B.n148 VSUBS 0.007794f
C230 B.n149 VSUBS 0.007794f
C231 B.n150 VSUBS 0.007794f
C232 B.n151 VSUBS 0.007794f
C233 B.n152 VSUBS 0.007794f
C234 B.n153 VSUBS 0.007794f
C235 B.n154 VSUBS 0.007794f
C236 B.n155 VSUBS 0.007794f
C237 B.n156 VSUBS 0.007794f
C238 B.n157 VSUBS 0.007794f
C239 B.n158 VSUBS 0.007794f
C240 B.n159 VSUBS 0.007794f
C241 B.n160 VSUBS 0.007794f
C242 B.n161 VSUBS 0.007794f
C243 B.n162 VSUBS 0.007794f
C244 B.n163 VSUBS 0.007794f
C245 B.n164 VSUBS 0.007794f
C246 B.n165 VSUBS 0.007794f
C247 B.n166 VSUBS 0.007794f
C248 B.n167 VSUBS 0.007794f
C249 B.n168 VSUBS 0.007794f
C250 B.n169 VSUBS 0.007794f
C251 B.n170 VSUBS 0.007794f
C252 B.n171 VSUBS 0.007794f
C253 B.n172 VSUBS 0.007794f
C254 B.n173 VSUBS 0.016088f
C255 B.n174 VSUBS 0.017152f
C256 B.n175 VSUBS 0.017152f
C257 B.n176 VSUBS 0.007794f
C258 B.n177 VSUBS 0.007794f
C259 B.n178 VSUBS 0.007794f
C260 B.n179 VSUBS 0.007794f
C261 B.n180 VSUBS 0.007794f
C262 B.n181 VSUBS 0.007794f
C263 B.n182 VSUBS 0.007794f
C264 B.n183 VSUBS 0.007794f
C265 B.n184 VSUBS 0.007794f
C266 B.n185 VSUBS 0.007794f
C267 B.n186 VSUBS 0.007794f
C268 B.n187 VSUBS 0.007794f
C269 B.n188 VSUBS 0.007794f
C270 B.n189 VSUBS 0.007794f
C271 B.n190 VSUBS 0.007794f
C272 B.n191 VSUBS 0.007794f
C273 B.n192 VSUBS 0.007794f
C274 B.n193 VSUBS 0.007794f
C275 B.n194 VSUBS 0.007794f
C276 B.n195 VSUBS 0.007794f
C277 B.n196 VSUBS 0.007794f
C278 B.n197 VSUBS 0.007794f
C279 B.n198 VSUBS 0.007794f
C280 B.n199 VSUBS 0.007794f
C281 B.n200 VSUBS 0.007794f
C282 B.n201 VSUBS 0.007794f
C283 B.n202 VSUBS 0.007794f
C284 B.n203 VSUBS 0.007794f
C285 B.n204 VSUBS 0.007794f
C286 B.n205 VSUBS 0.007794f
C287 B.n206 VSUBS 0.007794f
C288 B.n207 VSUBS 0.007794f
C289 B.n208 VSUBS 0.007794f
C290 B.n209 VSUBS 0.007794f
C291 B.n210 VSUBS 0.007794f
C292 B.n211 VSUBS 0.007794f
C293 B.n212 VSUBS 0.007794f
C294 B.n213 VSUBS 0.007794f
C295 B.n214 VSUBS 0.007794f
C296 B.n215 VSUBS 0.007794f
C297 B.n216 VSUBS 0.007794f
C298 B.n217 VSUBS 0.007794f
C299 B.n218 VSUBS 0.007794f
C300 B.n219 VSUBS 0.007794f
C301 B.n220 VSUBS 0.007794f
C302 B.n221 VSUBS 0.007794f
C303 B.n222 VSUBS 0.007794f
C304 B.n223 VSUBS 0.007794f
C305 B.n224 VSUBS 0.007794f
C306 B.n225 VSUBS 0.007794f
C307 B.n226 VSUBS 0.007794f
C308 B.n227 VSUBS 0.007794f
C309 B.n228 VSUBS 0.007794f
C310 B.n229 VSUBS 0.007794f
C311 B.n230 VSUBS 0.007794f
C312 B.n231 VSUBS 0.007794f
C313 B.n232 VSUBS 0.007794f
C314 B.n233 VSUBS 0.007794f
C315 B.n234 VSUBS 0.007794f
C316 B.n235 VSUBS 0.007794f
C317 B.n236 VSUBS 0.007794f
C318 B.n237 VSUBS 0.007794f
C319 B.n238 VSUBS 0.007794f
C320 B.n239 VSUBS 0.007794f
C321 B.n240 VSUBS 0.007794f
C322 B.n241 VSUBS 0.007336f
C323 B.n242 VSUBS 0.018058f
C324 B.n243 VSUBS 0.004356f
C325 B.n244 VSUBS 0.007794f
C326 B.n245 VSUBS 0.007794f
C327 B.n246 VSUBS 0.007794f
C328 B.n247 VSUBS 0.007794f
C329 B.n248 VSUBS 0.007794f
C330 B.n249 VSUBS 0.007794f
C331 B.n250 VSUBS 0.007794f
C332 B.n251 VSUBS 0.007794f
C333 B.n252 VSUBS 0.007794f
C334 B.n253 VSUBS 0.007794f
C335 B.n254 VSUBS 0.007794f
C336 B.n255 VSUBS 0.007794f
C337 B.t2 VSUBS 0.481643f
C338 B.t1 VSUBS 0.49274f
C339 B.t0 VSUBS 0.576639f
C340 B.n256 VSUBS 0.182458f
C341 B.n257 VSUBS 0.07237f
C342 B.n258 VSUBS 0.018058f
C343 B.n259 VSUBS 0.004356f
C344 B.n260 VSUBS 0.007794f
C345 B.n261 VSUBS 0.007794f
C346 B.n262 VSUBS 0.007794f
C347 B.n263 VSUBS 0.007794f
C348 B.n264 VSUBS 0.007794f
C349 B.n265 VSUBS 0.007794f
C350 B.n266 VSUBS 0.007794f
C351 B.n267 VSUBS 0.007794f
C352 B.n268 VSUBS 0.007794f
C353 B.n269 VSUBS 0.007794f
C354 B.n270 VSUBS 0.007794f
C355 B.n271 VSUBS 0.007794f
C356 B.n272 VSUBS 0.007794f
C357 B.n273 VSUBS 0.007794f
C358 B.n274 VSUBS 0.007794f
C359 B.n275 VSUBS 0.007794f
C360 B.n276 VSUBS 0.007794f
C361 B.n277 VSUBS 0.007794f
C362 B.n278 VSUBS 0.007794f
C363 B.n279 VSUBS 0.007794f
C364 B.n280 VSUBS 0.007794f
C365 B.n281 VSUBS 0.007794f
C366 B.n282 VSUBS 0.007794f
C367 B.n283 VSUBS 0.007794f
C368 B.n284 VSUBS 0.007794f
C369 B.n285 VSUBS 0.007794f
C370 B.n286 VSUBS 0.007794f
C371 B.n287 VSUBS 0.007794f
C372 B.n288 VSUBS 0.007794f
C373 B.n289 VSUBS 0.007794f
C374 B.n290 VSUBS 0.007794f
C375 B.n291 VSUBS 0.007794f
C376 B.n292 VSUBS 0.007794f
C377 B.n293 VSUBS 0.007794f
C378 B.n294 VSUBS 0.007794f
C379 B.n295 VSUBS 0.007794f
C380 B.n296 VSUBS 0.007794f
C381 B.n297 VSUBS 0.007794f
C382 B.n298 VSUBS 0.007794f
C383 B.n299 VSUBS 0.007794f
C384 B.n300 VSUBS 0.007794f
C385 B.n301 VSUBS 0.007794f
C386 B.n302 VSUBS 0.007794f
C387 B.n303 VSUBS 0.007794f
C388 B.n304 VSUBS 0.007794f
C389 B.n305 VSUBS 0.007794f
C390 B.n306 VSUBS 0.007794f
C391 B.n307 VSUBS 0.007794f
C392 B.n308 VSUBS 0.007794f
C393 B.n309 VSUBS 0.007794f
C394 B.n310 VSUBS 0.007794f
C395 B.n311 VSUBS 0.007794f
C396 B.n312 VSUBS 0.007794f
C397 B.n313 VSUBS 0.007794f
C398 B.n314 VSUBS 0.007794f
C399 B.n315 VSUBS 0.007794f
C400 B.n316 VSUBS 0.007794f
C401 B.n317 VSUBS 0.007794f
C402 B.n318 VSUBS 0.007794f
C403 B.n319 VSUBS 0.007794f
C404 B.n320 VSUBS 0.007794f
C405 B.n321 VSUBS 0.007794f
C406 B.n322 VSUBS 0.007794f
C407 B.n323 VSUBS 0.007794f
C408 B.n324 VSUBS 0.007794f
C409 B.n325 VSUBS 0.007794f
C410 B.n326 VSUBS 0.007794f
C411 B.n327 VSUBS 0.017152f
C412 B.n328 VSUBS 0.016088f
C413 B.n329 VSUBS 0.017152f
C414 B.n330 VSUBS 0.007794f
C415 B.n331 VSUBS 0.007794f
C416 B.n332 VSUBS 0.007794f
C417 B.n333 VSUBS 0.007794f
C418 B.n334 VSUBS 0.007794f
C419 B.n335 VSUBS 0.007794f
C420 B.n336 VSUBS 0.007794f
C421 B.n337 VSUBS 0.007794f
C422 B.n338 VSUBS 0.007794f
C423 B.n339 VSUBS 0.007794f
C424 B.n340 VSUBS 0.007794f
C425 B.n341 VSUBS 0.007794f
C426 B.n342 VSUBS 0.007794f
C427 B.n343 VSUBS 0.007794f
C428 B.n344 VSUBS 0.007794f
C429 B.n345 VSUBS 0.007794f
C430 B.n346 VSUBS 0.007794f
C431 B.n347 VSUBS 0.007794f
C432 B.n348 VSUBS 0.007794f
C433 B.n349 VSUBS 0.007794f
C434 B.n350 VSUBS 0.007794f
C435 B.n351 VSUBS 0.007794f
C436 B.n352 VSUBS 0.007794f
C437 B.n353 VSUBS 0.007794f
C438 B.n354 VSUBS 0.007794f
C439 B.n355 VSUBS 0.007794f
C440 B.n356 VSUBS 0.007794f
C441 B.n357 VSUBS 0.007794f
C442 B.n358 VSUBS 0.007794f
C443 B.n359 VSUBS 0.007794f
C444 B.n360 VSUBS 0.007794f
C445 B.n361 VSUBS 0.007794f
C446 B.n362 VSUBS 0.007794f
C447 B.n363 VSUBS 0.007794f
C448 B.n364 VSUBS 0.007794f
C449 B.n365 VSUBS 0.007794f
C450 B.n366 VSUBS 0.007794f
C451 B.n367 VSUBS 0.007794f
C452 B.n368 VSUBS 0.007794f
C453 B.n369 VSUBS 0.007794f
C454 B.n370 VSUBS 0.007794f
C455 B.n371 VSUBS 0.007794f
C456 B.n372 VSUBS 0.007794f
C457 B.n373 VSUBS 0.007794f
C458 B.n374 VSUBS 0.007794f
C459 B.n375 VSUBS 0.007794f
C460 B.n376 VSUBS 0.007794f
C461 B.n377 VSUBS 0.007794f
C462 B.n378 VSUBS 0.007794f
C463 B.n379 VSUBS 0.007794f
C464 B.n380 VSUBS 0.007794f
C465 B.n381 VSUBS 0.007794f
C466 B.n382 VSUBS 0.007794f
C467 B.n383 VSUBS 0.007794f
C468 B.n384 VSUBS 0.007794f
C469 B.n385 VSUBS 0.007794f
C470 B.n386 VSUBS 0.007794f
C471 B.n387 VSUBS 0.016088f
C472 B.n388 VSUBS 0.017152f
C473 B.n389 VSUBS 0.017152f
C474 B.n390 VSUBS 0.007794f
C475 B.n391 VSUBS 0.007794f
C476 B.n392 VSUBS 0.007794f
C477 B.n393 VSUBS 0.007794f
C478 B.n394 VSUBS 0.007794f
C479 B.n395 VSUBS 0.007794f
C480 B.n396 VSUBS 0.007794f
C481 B.n397 VSUBS 0.007794f
C482 B.n398 VSUBS 0.007794f
C483 B.n399 VSUBS 0.007794f
C484 B.n400 VSUBS 0.007794f
C485 B.n401 VSUBS 0.007794f
C486 B.n402 VSUBS 0.007794f
C487 B.n403 VSUBS 0.007794f
C488 B.n404 VSUBS 0.007794f
C489 B.n405 VSUBS 0.007794f
C490 B.n406 VSUBS 0.007794f
C491 B.n407 VSUBS 0.007794f
C492 B.n408 VSUBS 0.007794f
C493 B.n409 VSUBS 0.007794f
C494 B.n410 VSUBS 0.007794f
C495 B.n411 VSUBS 0.007794f
C496 B.n412 VSUBS 0.007794f
C497 B.n413 VSUBS 0.007794f
C498 B.n414 VSUBS 0.007794f
C499 B.n415 VSUBS 0.007794f
C500 B.n416 VSUBS 0.007794f
C501 B.n417 VSUBS 0.007794f
C502 B.n418 VSUBS 0.007794f
C503 B.n419 VSUBS 0.007794f
C504 B.n420 VSUBS 0.007794f
C505 B.n421 VSUBS 0.007794f
C506 B.n422 VSUBS 0.007794f
C507 B.n423 VSUBS 0.007794f
C508 B.n424 VSUBS 0.007794f
C509 B.n425 VSUBS 0.007794f
C510 B.n426 VSUBS 0.007794f
C511 B.n427 VSUBS 0.007794f
C512 B.n428 VSUBS 0.007794f
C513 B.n429 VSUBS 0.007794f
C514 B.n430 VSUBS 0.007794f
C515 B.n431 VSUBS 0.007794f
C516 B.n432 VSUBS 0.007794f
C517 B.n433 VSUBS 0.007794f
C518 B.n434 VSUBS 0.007794f
C519 B.n435 VSUBS 0.007794f
C520 B.n436 VSUBS 0.007794f
C521 B.n437 VSUBS 0.007794f
C522 B.n438 VSUBS 0.007794f
C523 B.n439 VSUBS 0.007794f
C524 B.n440 VSUBS 0.007794f
C525 B.n441 VSUBS 0.007794f
C526 B.n442 VSUBS 0.007794f
C527 B.n443 VSUBS 0.007794f
C528 B.n444 VSUBS 0.007794f
C529 B.n445 VSUBS 0.007794f
C530 B.n446 VSUBS 0.007794f
C531 B.n447 VSUBS 0.007794f
C532 B.n448 VSUBS 0.007794f
C533 B.n449 VSUBS 0.007794f
C534 B.n450 VSUBS 0.007794f
C535 B.n451 VSUBS 0.007794f
C536 B.n452 VSUBS 0.007794f
C537 B.n453 VSUBS 0.007794f
C538 B.n454 VSUBS 0.007794f
C539 B.n455 VSUBS 0.007336f
C540 B.n456 VSUBS 0.018058f
C541 B.n457 VSUBS 0.004356f
C542 B.n458 VSUBS 0.007794f
C543 B.n459 VSUBS 0.007794f
C544 B.n460 VSUBS 0.007794f
C545 B.n461 VSUBS 0.007794f
C546 B.n462 VSUBS 0.007794f
C547 B.n463 VSUBS 0.007794f
C548 B.n464 VSUBS 0.007794f
C549 B.n465 VSUBS 0.007794f
C550 B.n466 VSUBS 0.007794f
C551 B.n467 VSUBS 0.007794f
C552 B.n468 VSUBS 0.007794f
C553 B.n469 VSUBS 0.007794f
C554 B.n470 VSUBS 0.004356f
C555 B.n471 VSUBS 0.007794f
C556 B.n472 VSUBS 0.007794f
C557 B.n473 VSUBS 0.007336f
C558 B.n474 VSUBS 0.007794f
C559 B.n475 VSUBS 0.007794f
C560 B.n476 VSUBS 0.007794f
C561 B.n477 VSUBS 0.007794f
C562 B.n478 VSUBS 0.007794f
C563 B.n479 VSUBS 0.007794f
C564 B.n480 VSUBS 0.007794f
C565 B.n481 VSUBS 0.007794f
C566 B.n482 VSUBS 0.007794f
C567 B.n483 VSUBS 0.007794f
C568 B.n484 VSUBS 0.007794f
C569 B.n485 VSUBS 0.007794f
C570 B.n486 VSUBS 0.007794f
C571 B.n487 VSUBS 0.007794f
C572 B.n488 VSUBS 0.007794f
C573 B.n489 VSUBS 0.007794f
C574 B.n490 VSUBS 0.007794f
C575 B.n491 VSUBS 0.007794f
C576 B.n492 VSUBS 0.007794f
C577 B.n493 VSUBS 0.007794f
C578 B.n494 VSUBS 0.007794f
C579 B.n495 VSUBS 0.007794f
C580 B.n496 VSUBS 0.007794f
C581 B.n497 VSUBS 0.007794f
C582 B.n498 VSUBS 0.007794f
C583 B.n499 VSUBS 0.007794f
C584 B.n500 VSUBS 0.007794f
C585 B.n501 VSUBS 0.007794f
C586 B.n502 VSUBS 0.007794f
C587 B.n503 VSUBS 0.007794f
C588 B.n504 VSUBS 0.007794f
C589 B.n505 VSUBS 0.007794f
C590 B.n506 VSUBS 0.007794f
C591 B.n507 VSUBS 0.007794f
C592 B.n508 VSUBS 0.007794f
C593 B.n509 VSUBS 0.007794f
C594 B.n510 VSUBS 0.007794f
C595 B.n511 VSUBS 0.007794f
C596 B.n512 VSUBS 0.007794f
C597 B.n513 VSUBS 0.007794f
C598 B.n514 VSUBS 0.007794f
C599 B.n515 VSUBS 0.007794f
C600 B.n516 VSUBS 0.007794f
C601 B.n517 VSUBS 0.007794f
C602 B.n518 VSUBS 0.007794f
C603 B.n519 VSUBS 0.007794f
C604 B.n520 VSUBS 0.007794f
C605 B.n521 VSUBS 0.007794f
C606 B.n522 VSUBS 0.007794f
C607 B.n523 VSUBS 0.007794f
C608 B.n524 VSUBS 0.007794f
C609 B.n525 VSUBS 0.007794f
C610 B.n526 VSUBS 0.007794f
C611 B.n527 VSUBS 0.007794f
C612 B.n528 VSUBS 0.007794f
C613 B.n529 VSUBS 0.007794f
C614 B.n530 VSUBS 0.007794f
C615 B.n531 VSUBS 0.007794f
C616 B.n532 VSUBS 0.007794f
C617 B.n533 VSUBS 0.007794f
C618 B.n534 VSUBS 0.007794f
C619 B.n535 VSUBS 0.007794f
C620 B.n536 VSUBS 0.007794f
C621 B.n537 VSUBS 0.007794f
C622 B.n538 VSUBS 0.017152f
C623 B.n539 VSUBS 0.017152f
C624 B.n540 VSUBS 0.016088f
C625 B.n541 VSUBS 0.007794f
C626 B.n542 VSUBS 0.007794f
C627 B.n543 VSUBS 0.007794f
C628 B.n544 VSUBS 0.007794f
C629 B.n545 VSUBS 0.007794f
C630 B.n546 VSUBS 0.007794f
C631 B.n547 VSUBS 0.007794f
C632 B.n548 VSUBS 0.007794f
C633 B.n549 VSUBS 0.007794f
C634 B.n550 VSUBS 0.007794f
C635 B.n551 VSUBS 0.007794f
C636 B.n552 VSUBS 0.007794f
C637 B.n553 VSUBS 0.007794f
C638 B.n554 VSUBS 0.007794f
C639 B.n555 VSUBS 0.007794f
C640 B.n556 VSUBS 0.007794f
C641 B.n557 VSUBS 0.007794f
C642 B.n558 VSUBS 0.007794f
C643 B.n559 VSUBS 0.007794f
C644 B.n560 VSUBS 0.007794f
C645 B.n561 VSUBS 0.007794f
C646 B.n562 VSUBS 0.007794f
C647 B.n563 VSUBS 0.007794f
C648 B.n564 VSUBS 0.007794f
C649 B.n565 VSUBS 0.007794f
C650 B.n566 VSUBS 0.007794f
C651 B.n567 VSUBS 0.010171f
C652 B.n568 VSUBS 0.010835f
C653 B.n569 VSUBS 0.021546f
.ends

