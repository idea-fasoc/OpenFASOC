* NGSPICE file created from diff_pair_sample_0856.ext - technology: sky130A

.subckt diff_pair_sample_0856 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=0 ps=0 w=11.22 l=0.8
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=0 ps=0 w=11.22 l=0.8
X2 VTAIL.t11 VP.t0 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=1.8513 ps=11.55 w=11.22 l=0.8
X3 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=0 ps=0 w=11.22 l=0.8
X4 VTAIL.t3 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=1.8513 ps=11.55 w=11.22 l=0.8
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=0 ps=0 w=11.22 l=0.8
X6 VDD1.t4 VP.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=1.8513 ps=11.55 w=11.22 l=0.8
X7 VDD2.t4 VN.t1 VTAIL.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=1.8513 ps=11.55 w=11.22 l=0.8
X8 VTAIL.t1 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=1.8513 ps=11.55 w=11.22 l=0.8
X9 VDD2.t2 VN.t3 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=4.3758 ps=23.22 w=11.22 l=0.8
X10 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=4.3758 ps=23.22 w=11.22 l=0.8
X11 VDD1.t0 VP.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=4.3758 ps=23.22 w=11.22 l=0.8
X12 VDD2.t0 VN.t5 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=1.8513 ps=11.55 w=11.22 l=0.8
X13 VDD1.t3 VP.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=4.3758 ps=23.22 w=11.22 l=0.8
X14 VTAIL.t7 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8513 pd=11.55 as=1.8513 ps=11.55 w=11.22 l=0.8
X15 VDD1.t5 VP.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3758 pd=23.22 as=1.8513 ps=11.55 w=11.22 l=0.8
R0 B.n624 B.n623 585
R1 B.n265 B.n86 585
R2 B.n264 B.n263 585
R3 B.n262 B.n261 585
R4 B.n260 B.n259 585
R5 B.n258 B.n257 585
R6 B.n256 B.n255 585
R7 B.n254 B.n253 585
R8 B.n252 B.n251 585
R9 B.n250 B.n249 585
R10 B.n248 B.n247 585
R11 B.n246 B.n245 585
R12 B.n244 B.n243 585
R13 B.n242 B.n241 585
R14 B.n240 B.n239 585
R15 B.n238 B.n237 585
R16 B.n236 B.n235 585
R17 B.n234 B.n233 585
R18 B.n232 B.n231 585
R19 B.n230 B.n229 585
R20 B.n228 B.n227 585
R21 B.n226 B.n225 585
R22 B.n224 B.n223 585
R23 B.n222 B.n221 585
R24 B.n220 B.n219 585
R25 B.n218 B.n217 585
R26 B.n216 B.n215 585
R27 B.n214 B.n213 585
R28 B.n212 B.n211 585
R29 B.n210 B.n209 585
R30 B.n208 B.n207 585
R31 B.n206 B.n205 585
R32 B.n204 B.n203 585
R33 B.n202 B.n201 585
R34 B.n200 B.n199 585
R35 B.n198 B.n197 585
R36 B.n196 B.n195 585
R37 B.n194 B.n193 585
R38 B.n192 B.n191 585
R39 B.n189 B.n188 585
R40 B.n187 B.n186 585
R41 B.n185 B.n184 585
R42 B.n183 B.n182 585
R43 B.n181 B.n180 585
R44 B.n179 B.n178 585
R45 B.n177 B.n176 585
R46 B.n175 B.n174 585
R47 B.n173 B.n172 585
R48 B.n171 B.n170 585
R49 B.n168 B.n167 585
R50 B.n166 B.n165 585
R51 B.n164 B.n163 585
R52 B.n162 B.n161 585
R53 B.n160 B.n159 585
R54 B.n158 B.n157 585
R55 B.n156 B.n155 585
R56 B.n154 B.n153 585
R57 B.n152 B.n151 585
R58 B.n150 B.n149 585
R59 B.n148 B.n147 585
R60 B.n146 B.n145 585
R61 B.n144 B.n143 585
R62 B.n142 B.n141 585
R63 B.n140 B.n139 585
R64 B.n138 B.n137 585
R65 B.n136 B.n135 585
R66 B.n134 B.n133 585
R67 B.n132 B.n131 585
R68 B.n130 B.n129 585
R69 B.n128 B.n127 585
R70 B.n126 B.n125 585
R71 B.n124 B.n123 585
R72 B.n122 B.n121 585
R73 B.n120 B.n119 585
R74 B.n118 B.n117 585
R75 B.n116 B.n115 585
R76 B.n114 B.n113 585
R77 B.n112 B.n111 585
R78 B.n110 B.n109 585
R79 B.n108 B.n107 585
R80 B.n106 B.n105 585
R81 B.n104 B.n103 585
R82 B.n102 B.n101 585
R83 B.n100 B.n99 585
R84 B.n98 B.n97 585
R85 B.n96 B.n95 585
R86 B.n94 B.n93 585
R87 B.n92 B.n91 585
R88 B.n622 B.n42 585
R89 B.n627 B.n42 585
R90 B.n621 B.n41 585
R91 B.n628 B.n41 585
R92 B.n620 B.n619 585
R93 B.n619 B.n37 585
R94 B.n618 B.n36 585
R95 B.n634 B.n36 585
R96 B.n617 B.n35 585
R97 B.n635 B.n35 585
R98 B.n616 B.n34 585
R99 B.n636 B.n34 585
R100 B.n615 B.n614 585
R101 B.n614 B.n30 585
R102 B.n613 B.n29 585
R103 B.n642 B.n29 585
R104 B.n612 B.n28 585
R105 B.n643 B.n28 585
R106 B.n611 B.n27 585
R107 B.n644 B.n27 585
R108 B.n610 B.n609 585
R109 B.n609 B.n23 585
R110 B.n608 B.n22 585
R111 B.n650 B.n22 585
R112 B.n607 B.n21 585
R113 B.n651 B.n21 585
R114 B.n606 B.n20 585
R115 B.n652 B.n20 585
R116 B.n605 B.n604 585
R117 B.n604 B.n19 585
R118 B.n603 B.n15 585
R119 B.n658 B.n15 585
R120 B.n602 B.n14 585
R121 B.n659 B.n14 585
R122 B.n601 B.n13 585
R123 B.n660 B.n13 585
R124 B.n600 B.n599 585
R125 B.n599 B.n12 585
R126 B.n598 B.n597 585
R127 B.n598 B.n8 585
R128 B.n596 B.n7 585
R129 B.n667 B.n7 585
R130 B.n595 B.n6 585
R131 B.n668 B.n6 585
R132 B.n594 B.n5 585
R133 B.n669 B.n5 585
R134 B.n593 B.n592 585
R135 B.n592 B.n4 585
R136 B.n591 B.n266 585
R137 B.n591 B.n590 585
R138 B.n580 B.n267 585
R139 B.n583 B.n267 585
R140 B.n582 B.n581 585
R141 B.n584 B.n582 585
R142 B.n579 B.n272 585
R143 B.n272 B.n271 585
R144 B.n578 B.n577 585
R145 B.n577 B.n576 585
R146 B.n274 B.n273 585
R147 B.n569 B.n274 585
R148 B.n568 B.n567 585
R149 B.n570 B.n568 585
R150 B.n566 B.n279 585
R151 B.n279 B.n278 585
R152 B.n565 B.n564 585
R153 B.n564 B.n563 585
R154 B.n281 B.n280 585
R155 B.n282 B.n281 585
R156 B.n556 B.n555 585
R157 B.n557 B.n556 585
R158 B.n554 B.n287 585
R159 B.n287 B.n286 585
R160 B.n553 B.n552 585
R161 B.n552 B.n551 585
R162 B.n289 B.n288 585
R163 B.n290 B.n289 585
R164 B.n544 B.n543 585
R165 B.n545 B.n544 585
R166 B.n542 B.n295 585
R167 B.n295 B.n294 585
R168 B.n541 B.n540 585
R169 B.n540 B.n539 585
R170 B.n297 B.n296 585
R171 B.n298 B.n297 585
R172 B.n532 B.n531 585
R173 B.n533 B.n532 585
R174 B.n530 B.n303 585
R175 B.n303 B.n302 585
R176 B.n525 B.n524 585
R177 B.n523 B.n349 585
R178 B.n522 B.n348 585
R179 B.n527 B.n348 585
R180 B.n521 B.n520 585
R181 B.n519 B.n518 585
R182 B.n517 B.n516 585
R183 B.n515 B.n514 585
R184 B.n513 B.n512 585
R185 B.n511 B.n510 585
R186 B.n509 B.n508 585
R187 B.n507 B.n506 585
R188 B.n505 B.n504 585
R189 B.n503 B.n502 585
R190 B.n501 B.n500 585
R191 B.n499 B.n498 585
R192 B.n497 B.n496 585
R193 B.n495 B.n494 585
R194 B.n493 B.n492 585
R195 B.n491 B.n490 585
R196 B.n489 B.n488 585
R197 B.n487 B.n486 585
R198 B.n485 B.n484 585
R199 B.n483 B.n482 585
R200 B.n481 B.n480 585
R201 B.n479 B.n478 585
R202 B.n477 B.n476 585
R203 B.n475 B.n474 585
R204 B.n473 B.n472 585
R205 B.n471 B.n470 585
R206 B.n469 B.n468 585
R207 B.n467 B.n466 585
R208 B.n465 B.n464 585
R209 B.n463 B.n462 585
R210 B.n461 B.n460 585
R211 B.n459 B.n458 585
R212 B.n457 B.n456 585
R213 B.n455 B.n454 585
R214 B.n453 B.n452 585
R215 B.n451 B.n450 585
R216 B.n449 B.n448 585
R217 B.n447 B.n446 585
R218 B.n445 B.n444 585
R219 B.n443 B.n442 585
R220 B.n441 B.n440 585
R221 B.n439 B.n438 585
R222 B.n437 B.n436 585
R223 B.n435 B.n434 585
R224 B.n433 B.n432 585
R225 B.n431 B.n430 585
R226 B.n429 B.n428 585
R227 B.n427 B.n426 585
R228 B.n425 B.n424 585
R229 B.n423 B.n422 585
R230 B.n421 B.n420 585
R231 B.n419 B.n418 585
R232 B.n417 B.n416 585
R233 B.n415 B.n414 585
R234 B.n413 B.n412 585
R235 B.n411 B.n410 585
R236 B.n409 B.n408 585
R237 B.n407 B.n406 585
R238 B.n405 B.n404 585
R239 B.n403 B.n402 585
R240 B.n401 B.n400 585
R241 B.n399 B.n398 585
R242 B.n397 B.n396 585
R243 B.n395 B.n394 585
R244 B.n393 B.n392 585
R245 B.n391 B.n390 585
R246 B.n389 B.n388 585
R247 B.n387 B.n386 585
R248 B.n385 B.n384 585
R249 B.n383 B.n382 585
R250 B.n381 B.n380 585
R251 B.n379 B.n378 585
R252 B.n377 B.n376 585
R253 B.n375 B.n374 585
R254 B.n373 B.n372 585
R255 B.n371 B.n370 585
R256 B.n369 B.n368 585
R257 B.n367 B.n366 585
R258 B.n365 B.n364 585
R259 B.n363 B.n362 585
R260 B.n361 B.n360 585
R261 B.n359 B.n358 585
R262 B.n357 B.n356 585
R263 B.n305 B.n304 585
R264 B.n529 B.n528 585
R265 B.n528 B.n527 585
R266 B.n301 B.n300 585
R267 B.n302 B.n301 585
R268 B.n535 B.n534 585
R269 B.n534 B.n533 585
R270 B.n536 B.n299 585
R271 B.n299 B.n298 585
R272 B.n538 B.n537 585
R273 B.n539 B.n538 585
R274 B.n293 B.n292 585
R275 B.n294 B.n293 585
R276 B.n547 B.n546 585
R277 B.n546 B.n545 585
R278 B.n548 B.n291 585
R279 B.n291 B.n290 585
R280 B.n550 B.n549 585
R281 B.n551 B.n550 585
R282 B.n285 B.n284 585
R283 B.n286 B.n285 585
R284 B.n559 B.n558 585
R285 B.n558 B.n557 585
R286 B.n560 B.n283 585
R287 B.n283 B.n282 585
R288 B.n562 B.n561 585
R289 B.n563 B.n562 585
R290 B.n277 B.n276 585
R291 B.n278 B.n277 585
R292 B.n572 B.n571 585
R293 B.n571 B.n570 585
R294 B.n573 B.n275 585
R295 B.n569 B.n275 585
R296 B.n575 B.n574 585
R297 B.n576 B.n575 585
R298 B.n270 B.n269 585
R299 B.n271 B.n270 585
R300 B.n586 B.n585 585
R301 B.n585 B.n584 585
R302 B.n587 B.n268 585
R303 B.n583 B.n268 585
R304 B.n589 B.n588 585
R305 B.n590 B.n589 585
R306 B.n3 B.n0 585
R307 B.n4 B.n3 585
R308 B.n666 B.n1 585
R309 B.n667 B.n666 585
R310 B.n665 B.n664 585
R311 B.n665 B.n8 585
R312 B.n663 B.n9 585
R313 B.n12 B.n9 585
R314 B.n662 B.n661 585
R315 B.n661 B.n660 585
R316 B.n11 B.n10 585
R317 B.n659 B.n11 585
R318 B.n657 B.n656 585
R319 B.n658 B.n657 585
R320 B.n655 B.n16 585
R321 B.n19 B.n16 585
R322 B.n654 B.n653 585
R323 B.n653 B.n652 585
R324 B.n18 B.n17 585
R325 B.n651 B.n18 585
R326 B.n649 B.n648 585
R327 B.n650 B.n649 585
R328 B.n647 B.n24 585
R329 B.n24 B.n23 585
R330 B.n646 B.n645 585
R331 B.n645 B.n644 585
R332 B.n26 B.n25 585
R333 B.n643 B.n26 585
R334 B.n641 B.n640 585
R335 B.n642 B.n641 585
R336 B.n639 B.n31 585
R337 B.n31 B.n30 585
R338 B.n638 B.n637 585
R339 B.n637 B.n636 585
R340 B.n33 B.n32 585
R341 B.n635 B.n33 585
R342 B.n633 B.n632 585
R343 B.n634 B.n633 585
R344 B.n631 B.n38 585
R345 B.n38 B.n37 585
R346 B.n630 B.n629 585
R347 B.n629 B.n628 585
R348 B.n40 B.n39 585
R349 B.n627 B.n40 585
R350 B.n670 B.n669 585
R351 B.n668 B.n2 585
R352 B.n89 B.t10 539.891
R353 B.n87 B.t17 539.891
R354 B.n353 B.t14 539.891
R355 B.n350 B.t6 539.891
R356 B.n91 B.n40 502.111
R357 B.n624 B.n42 502.111
R358 B.n528 B.n303 502.111
R359 B.n525 B.n301 502.111
R360 B.n87 B.t18 290.272
R361 B.n353 B.t16 290.272
R362 B.n89 B.t12 290.272
R363 B.n350 B.t9 290.272
R364 B.n88 B.t19 268.356
R365 B.n354 B.t15 268.356
R366 B.n90 B.t13 268.356
R367 B.n351 B.t8 268.356
R368 B.n626 B.n625 256.663
R369 B.n626 B.n85 256.663
R370 B.n626 B.n84 256.663
R371 B.n626 B.n83 256.663
R372 B.n626 B.n82 256.663
R373 B.n626 B.n81 256.663
R374 B.n626 B.n80 256.663
R375 B.n626 B.n79 256.663
R376 B.n626 B.n78 256.663
R377 B.n626 B.n77 256.663
R378 B.n626 B.n76 256.663
R379 B.n626 B.n75 256.663
R380 B.n626 B.n74 256.663
R381 B.n626 B.n73 256.663
R382 B.n626 B.n72 256.663
R383 B.n626 B.n71 256.663
R384 B.n626 B.n70 256.663
R385 B.n626 B.n69 256.663
R386 B.n626 B.n68 256.663
R387 B.n626 B.n67 256.663
R388 B.n626 B.n66 256.663
R389 B.n626 B.n65 256.663
R390 B.n626 B.n64 256.663
R391 B.n626 B.n63 256.663
R392 B.n626 B.n62 256.663
R393 B.n626 B.n61 256.663
R394 B.n626 B.n60 256.663
R395 B.n626 B.n59 256.663
R396 B.n626 B.n58 256.663
R397 B.n626 B.n57 256.663
R398 B.n626 B.n56 256.663
R399 B.n626 B.n55 256.663
R400 B.n626 B.n54 256.663
R401 B.n626 B.n53 256.663
R402 B.n626 B.n52 256.663
R403 B.n626 B.n51 256.663
R404 B.n626 B.n50 256.663
R405 B.n626 B.n49 256.663
R406 B.n626 B.n48 256.663
R407 B.n626 B.n47 256.663
R408 B.n626 B.n46 256.663
R409 B.n626 B.n45 256.663
R410 B.n626 B.n44 256.663
R411 B.n626 B.n43 256.663
R412 B.n527 B.n526 256.663
R413 B.n527 B.n306 256.663
R414 B.n527 B.n307 256.663
R415 B.n527 B.n308 256.663
R416 B.n527 B.n309 256.663
R417 B.n527 B.n310 256.663
R418 B.n527 B.n311 256.663
R419 B.n527 B.n312 256.663
R420 B.n527 B.n313 256.663
R421 B.n527 B.n314 256.663
R422 B.n527 B.n315 256.663
R423 B.n527 B.n316 256.663
R424 B.n527 B.n317 256.663
R425 B.n527 B.n318 256.663
R426 B.n527 B.n319 256.663
R427 B.n527 B.n320 256.663
R428 B.n527 B.n321 256.663
R429 B.n527 B.n322 256.663
R430 B.n527 B.n323 256.663
R431 B.n527 B.n324 256.663
R432 B.n527 B.n325 256.663
R433 B.n527 B.n326 256.663
R434 B.n527 B.n327 256.663
R435 B.n527 B.n328 256.663
R436 B.n527 B.n329 256.663
R437 B.n527 B.n330 256.663
R438 B.n527 B.n331 256.663
R439 B.n527 B.n332 256.663
R440 B.n527 B.n333 256.663
R441 B.n527 B.n334 256.663
R442 B.n527 B.n335 256.663
R443 B.n527 B.n336 256.663
R444 B.n527 B.n337 256.663
R445 B.n527 B.n338 256.663
R446 B.n527 B.n339 256.663
R447 B.n527 B.n340 256.663
R448 B.n527 B.n341 256.663
R449 B.n527 B.n342 256.663
R450 B.n527 B.n343 256.663
R451 B.n527 B.n344 256.663
R452 B.n527 B.n345 256.663
R453 B.n527 B.n346 256.663
R454 B.n527 B.n347 256.663
R455 B.n672 B.n671 256.663
R456 B.n95 B.n94 163.367
R457 B.n99 B.n98 163.367
R458 B.n103 B.n102 163.367
R459 B.n107 B.n106 163.367
R460 B.n111 B.n110 163.367
R461 B.n115 B.n114 163.367
R462 B.n119 B.n118 163.367
R463 B.n123 B.n122 163.367
R464 B.n127 B.n126 163.367
R465 B.n131 B.n130 163.367
R466 B.n135 B.n134 163.367
R467 B.n139 B.n138 163.367
R468 B.n143 B.n142 163.367
R469 B.n147 B.n146 163.367
R470 B.n151 B.n150 163.367
R471 B.n155 B.n154 163.367
R472 B.n159 B.n158 163.367
R473 B.n163 B.n162 163.367
R474 B.n167 B.n166 163.367
R475 B.n172 B.n171 163.367
R476 B.n176 B.n175 163.367
R477 B.n180 B.n179 163.367
R478 B.n184 B.n183 163.367
R479 B.n188 B.n187 163.367
R480 B.n193 B.n192 163.367
R481 B.n197 B.n196 163.367
R482 B.n201 B.n200 163.367
R483 B.n205 B.n204 163.367
R484 B.n209 B.n208 163.367
R485 B.n213 B.n212 163.367
R486 B.n217 B.n216 163.367
R487 B.n221 B.n220 163.367
R488 B.n225 B.n224 163.367
R489 B.n229 B.n228 163.367
R490 B.n233 B.n232 163.367
R491 B.n237 B.n236 163.367
R492 B.n241 B.n240 163.367
R493 B.n245 B.n244 163.367
R494 B.n249 B.n248 163.367
R495 B.n253 B.n252 163.367
R496 B.n257 B.n256 163.367
R497 B.n261 B.n260 163.367
R498 B.n263 B.n86 163.367
R499 B.n532 B.n303 163.367
R500 B.n532 B.n297 163.367
R501 B.n540 B.n297 163.367
R502 B.n540 B.n295 163.367
R503 B.n544 B.n295 163.367
R504 B.n544 B.n289 163.367
R505 B.n552 B.n289 163.367
R506 B.n552 B.n287 163.367
R507 B.n556 B.n287 163.367
R508 B.n556 B.n281 163.367
R509 B.n564 B.n281 163.367
R510 B.n564 B.n279 163.367
R511 B.n568 B.n279 163.367
R512 B.n568 B.n274 163.367
R513 B.n577 B.n274 163.367
R514 B.n577 B.n272 163.367
R515 B.n582 B.n272 163.367
R516 B.n582 B.n267 163.367
R517 B.n591 B.n267 163.367
R518 B.n592 B.n591 163.367
R519 B.n592 B.n5 163.367
R520 B.n6 B.n5 163.367
R521 B.n7 B.n6 163.367
R522 B.n598 B.n7 163.367
R523 B.n599 B.n598 163.367
R524 B.n599 B.n13 163.367
R525 B.n14 B.n13 163.367
R526 B.n15 B.n14 163.367
R527 B.n604 B.n15 163.367
R528 B.n604 B.n20 163.367
R529 B.n21 B.n20 163.367
R530 B.n22 B.n21 163.367
R531 B.n609 B.n22 163.367
R532 B.n609 B.n27 163.367
R533 B.n28 B.n27 163.367
R534 B.n29 B.n28 163.367
R535 B.n614 B.n29 163.367
R536 B.n614 B.n34 163.367
R537 B.n35 B.n34 163.367
R538 B.n36 B.n35 163.367
R539 B.n619 B.n36 163.367
R540 B.n619 B.n41 163.367
R541 B.n42 B.n41 163.367
R542 B.n349 B.n348 163.367
R543 B.n520 B.n348 163.367
R544 B.n518 B.n517 163.367
R545 B.n514 B.n513 163.367
R546 B.n510 B.n509 163.367
R547 B.n506 B.n505 163.367
R548 B.n502 B.n501 163.367
R549 B.n498 B.n497 163.367
R550 B.n494 B.n493 163.367
R551 B.n490 B.n489 163.367
R552 B.n486 B.n485 163.367
R553 B.n482 B.n481 163.367
R554 B.n478 B.n477 163.367
R555 B.n474 B.n473 163.367
R556 B.n470 B.n469 163.367
R557 B.n466 B.n465 163.367
R558 B.n462 B.n461 163.367
R559 B.n458 B.n457 163.367
R560 B.n454 B.n453 163.367
R561 B.n450 B.n449 163.367
R562 B.n446 B.n445 163.367
R563 B.n442 B.n441 163.367
R564 B.n438 B.n437 163.367
R565 B.n434 B.n433 163.367
R566 B.n430 B.n429 163.367
R567 B.n426 B.n425 163.367
R568 B.n422 B.n421 163.367
R569 B.n418 B.n417 163.367
R570 B.n414 B.n413 163.367
R571 B.n410 B.n409 163.367
R572 B.n406 B.n405 163.367
R573 B.n402 B.n401 163.367
R574 B.n398 B.n397 163.367
R575 B.n394 B.n393 163.367
R576 B.n390 B.n389 163.367
R577 B.n386 B.n385 163.367
R578 B.n382 B.n381 163.367
R579 B.n378 B.n377 163.367
R580 B.n374 B.n373 163.367
R581 B.n370 B.n369 163.367
R582 B.n366 B.n365 163.367
R583 B.n362 B.n361 163.367
R584 B.n358 B.n357 163.367
R585 B.n528 B.n305 163.367
R586 B.n534 B.n301 163.367
R587 B.n534 B.n299 163.367
R588 B.n538 B.n299 163.367
R589 B.n538 B.n293 163.367
R590 B.n546 B.n293 163.367
R591 B.n546 B.n291 163.367
R592 B.n550 B.n291 163.367
R593 B.n550 B.n285 163.367
R594 B.n558 B.n285 163.367
R595 B.n558 B.n283 163.367
R596 B.n562 B.n283 163.367
R597 B.n562 B.n277 163.367
R598 B.n571 B.n277 163.367
R599 B.n571 B.n275 163.367
R600 B.n575 B.n275 163.367
R601 B.n575 B.n270 163.367
R602 B.n585 B.n270 163.367
R603 B.n585 B.n268 163.367
R604 B.n589 B.n268 163.367
R605 B.n589 B.n3 163.367
R606 B.n670 B.n3 163.367
R607 B.n666 B.n2 163.367
R608 B.n666 B.n665 163.367
R609 B.n665 B.n9 163.367
R610 B.n661 B.n9 163.367
R611 B.n661 B.n11 163.367
R612 B.n657 B.n11 163.367
R613 B.n657 B.n16 163.367
R614 B.n653 B.n16 163.367
R615 B.n653 B.n18 163.367
R616 B.n649 B.n18 163.367
R617 B.n649 B.n24 163.367
R618 B.n645 B.n24 163.367
R619 B.n645 B.n26 163.367
R620 B.n641 B.n26 163.367
R621 B.n641 B.n31 163.367
R622 B.n637 B.n31 163.367
R623 B.n637 B.n33 163.367
R624 B.n633 B.n33 163.367
R625 B.n633 B.n38 163.367
R626 B.n629 B.n38 163.367
R627 B.n629 B.n40 163.367
R628 B.n527 B.n302 78.0241
R629 B.n627 B.n626 78.0241
R630 B.n91 B.n43 71.676
R631 B.n95 B.n44 71.676
R632 B.n99 B.n45 71.676
R633 B.n103 B.n46 71.676
R634 B.n107 B.n47 71.676
R635 B.n111 B.n48 71.676
R636 B.n115 B.n49 71.676
R637 B.n119 B.n50 71.676
R638 B.n123 B.n51 71.676
R639 B.n127 B.n52 71.676
R640 B.n131 B.n53 71.676
R641 B.n135 B.n54 71.676
R642 B.n139 B.n55 71.676
R643 B.n143 B.n56 71.676
R644 B.n147 B.n57 71.676
R645 B.n151 B.n58 71.676
R646 B.n155 B.n59 71.676
R647 B.n159 B.n60 71.676
R648 B.n163 B.n61 71.676
R649 B.n167 B.n62 71.676
R650 B.n172 B.n63 71.676
R651 B.n176 B.n64 71.676
R652 B.n180 B.n65 71.676
R653 B.n184 B.n66 71.676
R654 B.n188 B.n67 71.676
R655 B.n193 B.n68 71.676
R656 B.n197 B.n69 71.676
R657 B.n201 B.n70 71.676
R658 B.n205 B.n71 71.676
R659 B.n209 B.n72 71.676
R660 B.n213 B.n73 71.676
R661 B.n217 B.n74 71.676
R662 B.n221 B.n75 71.676
R663 B.n225 B.n76 71.676
R664 B.n229 B.n77 71.676
R665 B.n233 B.n78 71.676
R666 B.n237 B.n79 71.676
R667 B.n241 B.n80 71.676
R668 B.n245 B.n81 71.676
R669 B.n249 B.n82 71.676
R670 B.n253 B.n83 71.676
R671 B.n257 B.n84 71.676
R672 B.n261 B.n85 71.676
R673 B.n625 B.n86 71.676
R674 B.n625 B.n624 71.676
R675 B.n263 B.n85 71.676
R676 B.n260 B.n84 71.676
R677 B.n256 B.n83 71.676
R678 B.n252 B.n82 71.676
R679 B.n248 B.n81 71.676
R680 B.n244 B.n80 71.676
R681 B.n240 B.n79 71.676
R682 B.n236 B.n78 71.676
R683 B.n232 B.n77 71.676
R684 B.n228 B.n76 71.676
R685 B.n224 B.n75 71.676
R686 B.n220 B.n74 71.676
R687 B.n216 B.n73 71.676
R688 B.n212 B.n72 71.676
R689 B.n208 B.n71 71.676
R690 B.n204 B.n70 71.676
R691 B.n200 B.n69 71.676
R692 B.n196 B.n68 71.676
R693 B.n192 B.n67 71.676
R694 B.n187 B.n66 71.676
R695 B.n183 B.n65 71.676
R696 B.n179 B.n64 71.676
R697 B.n175 B.n63 71.676
R698 B.n171 B.n62 71.676
R699 B.n166 B.n61 71.676
R700 B.n162 B.n60 71.676
R701 B.n158 B.n59 71.676
R702 B.n154 B.n58 71.676
R703 B.n150 B.n57 71.676
R704 B.n146 B.n56 71.676
R705 B.n142 B.n55 71.676
R706 B.n138 B.n54 71.676
R707 B.n134 B.n53 71.676
R708 B.n130 B.n52 71.676
R709 B.n126 B.n51 71.676
R710 B.n122 B.n50 71.676
R711 B.n118 B.n49 71.676
R712 B.n114 B.n48 71.676
R713 B.n110 B.n47 71.676
R714 B.n106 B.n46 71.676
R715 B.n102 B.n45 71.676
R716 B.n98 B.n44 71.676
R717 B.n94 B.n43 71.676
R718 B.n526 B.n525 71.676
R719 B.n520 B.n306 71.676
R720 B.n517 B.n307 71.676
R721 B.n513 B.n308 71.676
R722 B.n509 B.n309 71.676
R723 B.n505 B.n310 71.676
R724 B.n501 B.n311 71.676
R725 B.n497 B.n312 71.676
R726 B.n493 B.n313 71.676
R727 B.n489 B.n314 71.676
R728 B.n485 B.n315 71.676
R729 B.n481 B.n316 71.676
R730 B.n477 B.n317 71.676
R731 B.n473 B.n318 71.676
R732 B.n469 B.n319 71.676
R733 B.n465 B.n320 71.676
R734 B.n461 B.n321 71.676
R735 B.n457 B.n322 71.676
R736 B.n453 B.n323 71.676
R737 B.n449 B.n324 71.676
R738 B.n445 B.n325 71.676
R739 B.n441 B.n326 71.676
R740 B.n437 B.n327 71.676
R741 B.n433 B.n328 71.676
R742 B.n429 B.n329 71.676
R743 B.n425 B.n330 71.676
R744 B.n421 B.n331 71.676
R745 B.n417 B.n332 71.676
R746 B.n413 B.n333 71.676
R747 B.n409 B.n334 71.676
R748 B.n405 B.n335 71.676
R749 B.n401 B.n336 71.676
R750 B.n397 B.n337 71.676
R751 B.n393 B.n338 71.676
R752 B.n389 B.n339 71.676
R753 B.n385 B.n340 71.676
R754 B.n381 B.n341 71.676
R755 B.n377 B.n342 71.676
R756 B.n373 B.n343 71.676
R757 B.n369 B.n344 71.676
R758 B.n365 B.n345 71.676
R759 B.n361 B.n346 71.676
R760 B.n357 B.n347 71.676
R761 B.n526 B.n349 71.676
R762 B.n518 B.n306 71.676
R763 B.n514 B.n307 71.676
R764 B.n510 B.n308 71.676
R765 B.n506 B.n309 71.676
R766 B.n502 B.n310 71.676
R767 B.n498 B.n311 71.676
R768 B.n494 B.n312 71.676
R769 B.n490 B.n313 71.676
R770 B.n486 B.n314 71.676
R771 B.n482 B.n315 71.676
R772 B.n478 B.n316 71.676
R773 B.n474 B.n317 71.676
R774 B.n470 B.n318 71.676
R775 B.n466 B.n319 71.676
R776 B.n462 B.n320 71.676
R777 B.n458 B.n321 71.676
R778 B.n454 B.n322 71.676
R779 B.n450 B.n323 71.676
R780 B.n446 B.n324 71.676
R781 B.n442 B.n325 71.676
R782 B.n438 B.n326 71.676
R783 B.n434 B.n327 71.676
R784 B.n430 B.n328 71.676
R785 B.n426 B.n329 71.676
R786 B.n422 B.n330 71.676
R787 B.n418 B.n331 71.676
R788 B.n414 B.n332 71.676
R789 B.n410 B.n333 71.676
R790 B.n406 B.n334 71.676
R791 B.n402 B.n335 71.676
R792 B.n398 B.n336 71.676
R793 B.n394 B.n337 71.676
R794 B.n390 B.n338 71.676
R795 B.n386 B.n339 71.676
R796 B.n382 B.n340 71.676
R797 B.n378 B.n341 71.676
R798 B.n374 B.n342 71.676
R799 B.n370 B.n343 71.676
R800 B.n366 B.n344 71.676
R801 B.n362 B.n345 71.676
R802 B.n358 B.n346 71.676
R803 B.n347 B.n305 71.676
R804 B.n671 B.n670 71.676
R805 B.n671 B.n2 71.676
R806 B.n169 B.n90 59.5399
R807 B.n190 B.n88 59.5399
R808 B.n355 B.n354 59.5399
R809 B.n352 B.n351 59.5399
R810 B.n533 B.n302 45.3476
R811 B.n533 B.n298 45.3476
R812 B.n539 B.n298 45.3476
R813 B.n539 B.n294 45.3476
R814 B.n545 B.n294 45.3476
R815 B.n551 B.n290 45.3476
R816 B.n551 B.n286 45.3476
R817 B.n557 B.n286 45.3476
R818 B.n557 B.n282 45.3476
R819 B.n563 B.n282 45.3476
R820 B.n570 B.n278 45.3476
R821 B.n570 B.n569 45.3476
R822 B.n576 B.n271 45.3476
R823 B.n584 B.n271 45.3476
R824 B.n584 B.n583 45.3476
R825 B.n590 B.n4 45.3476
R826 B.n669 B.n4 45.3476
R827 B.n669 B.n668 45.3476
R828 B.n668 B.n667 45.3476
R829 B.n667 B.n8 45.3476
R830 B.n660 B.n12 45.3476
R831 B.n660 B.n659 45.3476
R832 B.n659 B.n658 45.3476
R833 B.n652 B.n19 45.3476
R834 B.n652 B.n651 45.3476
R835 B.n650 B.n23 45.3476
R836 B.n644 B.n23 45.3476
R837 B.n644 B.n643 45.3476
R838 B.n643 B.n642 45.3476
R839 B.n642 B.n30 45.3476
R840 B.n636 B.n635 45.3476
R841 B.n635 B.n634 45.3476
R842 B.n634 B.n37 45.3476
R843 B.n628 B.n37 45.3476
R844 B.n628 B.n627 45.3476
R845 B.t7 B.n290 42.6801
R846 B.t11 B.n30 42.6801
R847 B.n569 B.t3 41.3464
R848 B.n19 B.t1 41.3464
R849 B.n590 B.t5 34.6777
R850 B.t0 B.n8 34.6777
R851 B.n524 B.n300 32.6249
R852 B.n530 B.n529 32.6249
R853 B.n623 B.n622 32.6249
R854 B.n92 B.n39 32.6249
R855 B.n563 B.t4 26.6752
R856 B.t2 B.n650 26.6752
R857 B.n90 B.n89 21.9157
R858 B.n88 B.n87 21.9157
R859 B.n354 B.n353 21.9157
R860 B.n351 B.n350 21.9157
R861 B.t4 B.n278 18.6728
R862 B.n651 B.t2 18.6728
R863 B B.n672 18.0485
R864 B.n583 B.t5 10.6704
R865 B.n12 B.t0 10.6704
R866 B.n535 B.n300 10.6151
R867 B.n536 B.n535 10.6151
R868 B.n537 B.n536 10.6151
R869 B.n537 B.n292 10.6151
R870 B.n547 B.n292 10.6151
R871 B.n548 B.n547 10.6151
R872 B.n549 B.n548 10.6151
R873 B.n549 B.n284 10.6151
R874 B.n559 B.n284 10.6151
R875 B.n560 B.n559 10.6151
R876 B.n561 B.n560 10.6151
R877 B.n561 B.n276 10.6151
R878 B.n572 B.n276 10.6151
R879 B.n573 B.n572 10.6151
R880 B.n574 B.n573 10.6151
R881 B.n574 B.n269 10.6151
R882 B.n586 B.n269 10.6151
R883 B.n587 B.n586 10.6151
R884 B.n588 B.n587 10.6151
R885 B.n588 B.n0 10.6151
R886 B.n524 B.n523 10.6151
R887 B.n523 B.n522 10.6151
R888 B.n522 B.n521 10.6151
R889 B.n521 B.n519 10.6151
R890 B.n519 B.n516 10.6151
R891 B.n516 B.n515 10.6151
R892 B.n515 B.n512 10.6151
R893 B.n512 B.n511 10.6151
R894 B.n511 B.n508 10.6151
R895 B.n508 B.n507 10.6151
R896 B.n507 B.n504 10.6151
R897 B.n504 B.n503 10.6151
R898 B.n503 B.n500 10.6151
R899 B.n500 B.n499 10.6151
R900 B.n499 B.n496 10.6151
R901 B.n496 B.n495 10.6151
R902 B.n495 B.n492 10.6151
R903 B.n492 B.n491 10.6151
R904 B.n491 B.n488 10.6151
R905 B.n488 B.n487 10.6151
R906 B.n487 B.n484 10.6151
R907 B.n484 B.n483 10.6151
R908 B.n483 B.n480 10.6151
R909 B.n480 B.n479 10.6151
R910 B.n479 B.n476 10.6151
R911 B.n476 B.n475 10.6151
R912 B.n475 B.n472 10.6151
R913 B.n472 B.n471 10.6151
R914 B.n471 B.n468 10.6151
R915 B.n468 B.n467 10.6151
R916 B.n467 B.n464 10.6151
R917 B.n464 B.n463 10.6151
R918 B.n463 B.n460 10.6151
R919 B.n460 B.n459 10.6151
R920 B.n459 B.n456 10.6151
R921 B.n456 B.n455 10.6151
R922 B.n455 B.n452 10.6151
R923 B.n452 B.n451 10.6151
R924 B.n448 B.n447 10.6151
R925 B.n447 B.n444 10.6151
R926 B.n444 B.n443 10.6151
R927 B.n443 B.n440 10.6151
R928 B.n440 B.n439 10.6151
R929 B.n439 B.n436 10.6151
R930 B.n436 B.n435 10.6151
R931 B.n435 B.n432 10.6151
R932 B.n432 B.n431 10.6151
R933 B.n428 B.n427 10.6151
R934 B.n427 B.n424 10.6151
R935 B.n424 B.n423 10.6151
R936 B.n423 B.n420 10.6151
R937 B.n420 B.n419 10.6151
R938 B.n419 B.n416 10.6151
R939 B.n416 B.n415 10.6151
R940 B.n415 B.n412 10.6151
R941 B.n412 B.n411 10.6151
R942 B.n411 B.n408 10.6151
R943 B.n408 B.n407 10.6151
R944 B.n407 B.n404 10.6151
R945 B.n404 B.n403 10.6151
R946 B.n403 B.n400 10.6151
R947 B.n400 B.n399 10.6151
R948 B.n399 B.n396 10.6151
R949 B.n396 B.n395 10.6151
R950 B.n395 B.n392 10.6151
R951 B.n392 B.n391 10.6151
R952 B.n391 B.n388 10.6151
R953 B.n388 B.n387 10.6151
R954 B.n387 B.n384 10.6151
R955 B.n384 B.n383 10.6151
R956 B.n383 B.n380 10.6151
R957 B.n380 B.n379 10.6151
R958 B.n379 B.n376 10.6151
R959 B.n376 B.n375 10.6151
R960 B.n375 B.n372 10.6151
R961 B.n372 B.n371 10.6151
R962 B.n371 B.n368 10.6151
R963 B.n368 B.n367 10.6151
R964 B.n367 B.n364 10.6151
R965 B.n364 B.n363 10.6151
R966 B.n363 B.n360 10.6151
R967 B.n360 B.n359 10.6151
R968 B.n359 B.n356 10.6151
R969 B.n356 B.n304 10.6151
R970 B.n529 B.n304 10.6151
R971 B.n531 B.n530 10.6151
R972 B.n531 B.n296 10.6151
R973 B.n541 B.n296 10.6151
R974 B.n542 B.n541 10.6151
R975 B.n543 B.n542 10.6151
R976 B.n543 B.n288 10.6151
R977 B.n553 B.n288 10.6151
R978 B.n554 B.n553 10.6151
R979 B.n555 B.n554 10.6151
R980 B.n555 B.n280 10.6151
R981 B.n565 B.n280 10.6151
R982 B.n566 B.n565 10.6151
R983 B.n567 B.n566 10.6151
R984 B.n567 B.n273 10.6151
R985 B.n578 B.n273 10.6151
R986 B.n579 B.n578 10.6151
R987 B.n581 B.n579 10.6151
R988 B.n581 B.n580 10.6151
R989 B.n580 B.n266 10.6151
R990 B.n593 B.n266 10.6151
R991 B.n594 B.n593 10.6151
R992 B.n595 B.n594 10.6151
R993 B.n596 B.n595 10.6151
R994 B.n597 B.n596 10.6151
R995 B.n600 B.n597 10.6151
R996 B.n601 B.n600 10.6151
R997 B.n602 B.n601 10.6151
R998 B.n603 B.n602 10.6151
R999 B.n605 B.n603 10.6151
R1000 B.n606 B.n605 10.6151
R1001 B.n607 B.n606 10.6151
R1002 B.n608 B.n607 10.6151
R1003 B.n610 B.n608 10.6151
R1004 B.n611 B.n610 10.6151
R1005 B.n612 B.n611 10.6151
R1006 B.n613 B.n612 10.6151
R1007 B.n615 B.n613 10.6151
R1008 B.n616 B.n615 10.6151
R1009 B.n617 B.n616 10.6151
R1010 B.n618 B.n617 10.6151
R1011 B.n620 B.n618 10.6151
R1012 B.n621 B.n620 10.6151
R1013 B.n622 B.n621 10.6151
R1014 B.n664 B.n1 10.6151
R1015 B.n664 B.n663 10.6151
R1016 B.n663 B.n662 10.6151
R1017 B.n662 B.n10 10.6151
R1018 B.n656 B.n10 10.6151
R1019 B.n656 B.n655 10.6151
R1020 B.n655 B.n654 10.6151
R1021 B.n654 B.n17 10.6151
R1022 B.n648 B.n17 10.6151
R1023 B.n648 B.n647 10.6151
R1024 B.n647 B.n646 10.6151
R1025 B.n646 B.n25 10.6151
R1026 B.n640 B.n25 10.6151
R1027 B.n640 B.n639 10.6151
R1028 B.n639 B.n638 10.6151
R1029 B.n638 B.n32 10.6151
R1030 B.n632 B.n32 10.6151
R1031 B.n632 B.n631 10.6151
R1032 B.n631 B.n630 10.6151
R1033 B.n630 B.n39 10.6151
R1034 B.n93 B.n92 10.6151
R1035 B.n96 B.n93 10.6151
R1036 B.n97 B.n96 10.6151
R1037 B.n100 B.n97 10.6151
R1038 B.n101 B.n100 10.6151
R1039 B.n104 B.n101 10.6151
R1040 B.n105 B.n104 10.6151
R1041 B.n108 B.n105 10.6151
R1042 B.n109 B.n108 10.6151
R1043 B.n112 B.n109 10.6151
R1044 B.n113 B.n112 10.6151
R1045 B.n116 B.n113 10.6151
R1046 B.n117 B.n116 10.6151
R1047 B.n120 B.n117 10.6151
R1048 B.n121 B.n120 10.6151
R1049 B.n124 B.n121 10.6151
R1050 B.n125 B.n124 10.6151
R1051 B.n128 B.n125 10.6151
R1052 B.n129 B.n128 10.6151
R1053 B.n132 B.n129 10.6151
R1054 B.n133 B.n132 10.6151
R1055 B.n136 B.n133 10.6151
R1056 B.n137 B.n136 10.6151
R1057 B.n140 B.n137 10.6151
R1058 B.n141 B.n140 10.6151
R1059 B.n144 B.n141 10.6151
R1060 B.n145 B.n144 10.6151
R1061 B.n148 B.n145 10.6151
R1062 B.n149 B.n148 10.6151
R1063 B.n152 B.n149 10.6151
R1064 B.n153 B.n152 10.6151
R1065 B.n156 B.n153 10.6151
R1066 B.n157 B.n156 10.6151
R1067 B.n160 B.n157 10.6151
R1068 B.n161 B.n160 10.6151
R1069 B.n164 B.n161 10.6151
R1070 B.n165 B.n164 10.6151
R1071 B.n168 B.n165 10.6151
R1072 B.n173 B.n170 10.6151
R1073 B.n174 B.n173 10.6151
R1074 B.n177 B.n174 10.6151
R1075 B.n178 B.n177 10.6151
R1076 B.n181 B.n178 10.6151
R1077 B.n182 B.n181 10.6151
R1078 B.n185 B.n182 10.6151
R1079 B.n186 B.n185 10.6151
R1080 B.n189 B.n186 10.6151
R1081 B.n194 B.n191 10.6151
R1082 B.n195 B.n194 10.6151
R1083 B.n198 B.n195 10.6151
R1084 B.n199 B.n198 10.6151
R1085 B.n202 B.n199 10.6151
R1086 B.n203 B.n202 10.6151
R1087 B.n206 B.n203 10.6151
R1088 B.n207 B.n206 10.6151
R1089 B.n210 B.n207 10.6151
R1090 B.n211 B.n210 10.6151
R1091 B.n214 B.n211 10.6151
R1092 B.n215 B.n214 10.6151
R1093 B.n218 B.n215 10.6151
R1094 B.n219 B.n218 10.6151
R1095 B.n222 B.n219 10.6151
R1096 B.n223 B.n222 10.6151
R1097 B.n226 B.n223 10.6151
R1098 B.n227 B.n226 10.6151
R1099 B.n230 B.n227 10.6151
R1100 B.n231 B.n230 10.6151
R1101 B.n234 B.n231 10.6151
R1102 B.n235 B.n234 10.6151
R1103 B.n238 B.n235 10.6151
R1104 B.n239 B.n238 10.6151
R1105 B.n242 B.n239 10.6151
R1106 B.n243 B.n242 10.6151
R1107 B.n246 B.n243 10.6151
R1108 B.n247 B.n246 10.6151
R1109 B.n250 B.n247 10.6151
R1110 B.n251 B.n250 10.6151
R1111 B.n254 B.n251 10.6151
R1112 B.n255 B.n254 10.6151
R1113 B.n258 B.n255 10.6151
R1114 B.n259 B.n258 10.6151
R1115 B.n262 B.n259 10.6151
R1116 B.n264 B.n262 10.6151
R1117 B.n265 B.n264 10.6151
R1118 B.n623 B.n265 10.6151
R1119 B.n451 B.n352 9.36635
R1120 B.n428 B.n355 9.36635
R1121 B.n169 B.n168 9.36635
R1122 B.n191 B.n190 9.36635
R1123 B.n672 B.n0 8.11757
R1124 B.n672 B.n1 8.11757
R1125 B.n576 B.t3 4.00171
R1126 B.n658 B.t1 4.00171
R1127 B.n545 B.t7 2.66797
R1128 B.n636 B.t11 2.66797
R1129 B.n448 B.n352 1.24928
R1130 B.n431 B.n355 1.24928
R1131 B.n170 B.n169 1.24928
R1132 B.n190 B.n189 1.24928
R1133 VP.n3 VP.t5 411.195
R1134 VP.n8 VP.t1 387.709
R1135 VP.n12 VP.t0 387.709
R1136 VP.n14 VP.t2 387.709
R1137 VP.n6 VP.t3 387.709
R1138 VP.n4 VP.t4 387.709
R1139 VP.n15 VP.n14 161.3
R1140 VP.n5 VP.n2 161.3
R1141 VP.n7 VP.n6 161.3
R1142 VP.n13 VP.n0 161.3
R1143 VP.n12 VP.n11 161.3
R1144 VP.n10 VP.n1 161.3
R1145 VP.n9 VP.n8 161.3
R1146 VP.n3 VP.n2 44.8973
R1147 VP.n9 VP.n7 41.1028
R1148 VP.n8 VP.n1 33.5944
R1149 VP.n14 VP.n13 33.5944
R1150 VP.n6 VP.n5 33.5944
R1151 VP.n4 VP.n3 18.1882
R1152 VP.n12 VP.n1 14.6066
R1153 VP.n13 VP.n12 14.6066
R1154 VP.n5 VP.n4 14.6066
R1155 VP.n7 VP.n2 0.189894
R1156 VP.n10 VP.n9 0.189894
R1157 VP.n11 VP.n10 0.189894
R1158 VP.n11 VP.n0 0.189894
R1159 VP.n15 VP.n0 0.189894
R1160 VP VP.n15 0.0516364
R1161 VDD1.n60 VDD1.n59 289.615
R1162 VDD1.n121 VDD1.n120 289.615
R1163 VDD1.n59 VDD1.n58 185
R1164 VDD1.n2 VDD1.n1 185
R1165 VDD1.n53 VDD1.n52 185
R1166 VDD1.n51 VDD1.n50 185
R1167 VDD1.n6 VDD1.n5 185
R1168 VDD1.n45 VDD1.n44 185
R1169 VDD1.n43 VDD1.n42 185
R1170 VDD1.n10 VDD1.n9 185
R1171 VDD1.n37 VDD1.n36 185
R1172 VDD1.n35 VDD1.n34 185
R1173 VDD1.n14 VDD1.n13 185
R1174 VDD1.n29 VDD1.n28 185
R1175 VDD1.n27 VDD1.n26 185
R1176 VDD1.n18 VDD1.n17 185
R1177 VDD1.n21 VDD1.n20 185
R1178 VDD1.n82 VDD1.n81 185
R1179 VDD1.n79 VDD1.n78 185
R1180 VDD1.n88 VDD1.n87 185
R1181 VDD1.n90 VDD1.n89 185
R1182 VDD1.n75 VDD1.n74 185
R1183 VDD1.n96 VDD1.n95 185
R1184 VDD1.n98 VDD1.n97 185
R1185 VDD1.n71 VDD1.n70 185
R1186 VDD1.n104 VDD1.n103 185
R1187 VDD1.n106 VDD1.n105 185
R1188 VDD1.n67 VDD1.n66 185
R1189 VDD1.n112 VDD1.n111 185
R1190 VDD1.n114 VDD1.n113 185
R1191 VDD1.n63 VDD1.n62 185
R1192 VDD1.n120 VDD1.n119 185
R1193 VDD1.t4 VDD1.n80 147.659
R1194 VDD1.t5 VDD1.n19 147.659
R1195 VDD1.n59 VDD1.n1 104.615
R1196 VDD1.n52 VDD1.n1 104.615
R1197 VDD1.n52 VDD1.n51 104.615
R1198 VDD1.n51 VDD1.n5 104.615
R1199 VDD1.n44 VDD1.n5 104.615
R1200 VDD1.n44 VDD1.n43 104.615
R1201 VDD1.n43 VDD1.n9 104.615
R1202 VDD1.n36 VDD1.n9 104.615
R1203 VDD1.n36 VDD1.n35 104.615
R1204 VDD1.n35 VDD1.n13 104.615
R1205 VDD1.n28 VDD1.n13 104.615
R1206 VDD1.n28 VDD1.n27 104.615
R1207 VDD1.n27 VDD1.n17 104.615
R1208 VDD1.n20 VDD1.n17 104.615
R1209 VDD1.n81 VDD1.n78 104.615
R1210 VDD1.n88 VDD1.n78 104.615
R1211 VDD1.n89 VDD1.n88 104.615
R1212 VDD1.n89 VDD1.n74 104.615
R1213 VDD1.n96 VDD1.n74 104.615
R1214 VDD1.n97 VDD1.n96 104.615
R1215 VDD1.n97 VDD1.n70 104.615
R1216 VDD1.n104 VDD1.n70 104.615
R1217 VDD1.n105 VDD1.n104 104.615
R1218 VDD1.n105 VDD1.n66 104.615
R1219 VDD1.n112 VDD1.n66 104.615
R1220 VDD1.n113 VDD1.n112 104.615
R1221 VDD1.n113 VDD1.n62 104.615
R1222 VDD1.n120 VDD1.n62 104.615
R1223 VDD1.n123 VDD1.n122 65.0635
R1224 VDD1.n125 VDD1.n124 64.8744
R1225 VDD1.n20 VDD1.t5 52.3082
R1226 VDD1.n81 VDD1.t4 52.3082
R1227 VDD1 VDD1.n60 51.2044
R1228 VDD1.n123 VDD1.n121 51.0909
R1229 VDD1.n125 VDD1.n123 37.6237
R1230 VDD1.n21 VDD1.n19 15.6677
R1231 VDD1.n82 VDD1.n80 15.6677
R1232 VDD1.n22 VDD1.n18 12.8005
R1233 VDD1.n83 VDD1.n79 12.8005
R1234 VDD1.n26 VDD1.n25 12.0247
R1235 VDD1.n87 VDD1.n86 12.0247
R1236 VDD1.n58 VDD1.n0 11.249
R1237 VDD1.n29 VDD1.n16 11.249
R1238 VDD1.n90 VDD1.n77 11.249
R1239 VDD1.n119 VDD1.n61 11.249
R1240 VDD1.n57 VDD1.n2 10.4732
R1241 VDD1.n30 VDD1.n14 10.4732
R1242 VDD1.n91 VDD1.n75 10.4732
R1243 VDD1.n118 VDD1.n63 10.4732
R1244 VDD1.n54 VDD1.n53 9.69747
R1245 VDD1.n34 VDD1.n33 9.69747
R1246 VDD1.n95 VDD1.n94 9.69747
R1247 VDD1.n115 VDD1.n114 9.69747
R1248 VDD1.n56 VDD1.n0 9.45567
R1249 VDD1.n117 VDD1.n61 9.45567
R1250 VDD1.n47 VDD1.n46 9.3005
R1251 VDD1.n49 VDD1.n48 9.3005
R1252 VDD1.n4 VDD1.n3 9.3005
R1253 VDD1.n55 VDD1.n54 9.3005
R1254 VDD1.n57 VDD1.n56 9.3005
R1255 VDD1.n8 VDD1.n7 9.3005
R1256 VDD1.n41 VDD1.n40 9.3005
R1257 VDD1.n39 VDD1.n38 9.3005
R1258 VDD1.n12 VDD1.n11 9.3005
R1259 VDD1.n33 VDD1.n32 9.3005
R1260 VDD1.n31 VDD1.n30 9.3005
R1261 VDD1.n16 VDD1.n15 9.3005
R1262 VDD1.n25 VDD1.n24 9.3005
R1263 VDD1.n23 VDD1.n22 9.3005
R1264 VDD1.n69 VDD1.n68 9.3005
R1265 VDD1.n108 VDD1.n107 9.3005
R1266 VDD1.n110 VDD1.n109 9.3005
R1267 VDD1.n65 VDD1.n64 9.3005
R1268 VDD1.n116 VDD1.n115 9.3005
R1269 VDD1.n118 VDD1.n117 9.3005
R1270 VDD1.n100 VDD1.n99 9.3005
R1271 VDD1.n73 VDD1.n72 9.3005
R1272 VDD1.n94 VDD1.n93 9.3005
R1273 VDD1.n92 VDD1.n91 9.3005
R1274 VDD1.n77 VDD1.n76 9.3005
R1275 VDD1.n86 VDD1.n85 9.3005
R1276 VDD1.n84 VDD1.n83 9.3005
R1277 VDD1.n102 VDD1.n101 9.3005
R1278 VDD1.n50 VDD1.n4 8.92171
R1279 VDD1.n37 VDD1.n12 8.92171
R1280 VDD1.n98 VDD1.n73 8.92171
R1281 VDD1.n111 VDD1.n65 8.92171
R1282 VDD1.n49 VDD1.n6 8.14595
R1283 VDD1.n38 VDD1.n10 8.14595
R1284 VDD1.n99 VDD1.n71 8.14595
R1285 VDD1.n110 VDD1.n67 8.14595
R1286 VDD1.n46 VDD1.n45 7.3702
R1287 VDD1.n42 VDD1.n41 7.3702
R1288 VDD1.n103 VDD1.n102 7.3702
R1289 VDD1.n107 VDD1.n106 7.3702
R1290 VDD1.n45 VDD1.n8 6.59444
R1291 VDD1.n42 VDD1.n8 6.59444
R1292 VDD1.n103 VDD1.n69 6.59444
R1293 VDD1.n106 VDD1.n69 6.59444
R1294 VDD1.n46 VDD1.n6 5.81868
R1295 VDD1.n41 VDD1.n10 5.81868
R1296 VDD1.n102 VDD1.n71 5.81868
R1297 VDD1.n107 VDD1.n67 5.81868
R1298 VDD1.n50 VDD1.n49 5.04292
R1299 VDD1.n38 VDD1.n37 5.04292
R1300 VDD1.n99 VDD1.n98 5.04292
R1301 VDD1.n111 VDD1.n110 5.04292
R1302 VDD1.n84 VDD1.n80 4.38563
R1303 VDD1.n23 VDD1.n19 4.38563
R1304 VDD1.n53 VDD1.n4 4.26717
R1305 VDD1.n34 VDD1.n12 4.26717
R1306 VDD1.n95 VDD1.n73 4.26717
R1307 VDD1.n114 VDD1.n65 4.26717
R1308 VDD1.n54 VDD1.n2 3.49141
R1309 VDD1.n33 VDD1.n14 3.49141
R1310 VDD1.n94 VDD1.n75 3.49141
R1311 VDD1.n115 VDD1.n63 3.49141
R1312 VDD1.n58 VDD1.n57 2.71565
R1313 VDD1.n30 VDD1.n29 2.71565
R1314 VDD1.n91 VDD1.n90 2.71565
R1315 VDD1.n119 VDD1.n118 2.71565
R1316 VDD1.n60 VDD1.n0 1.93989
R1317 VDD1.n26 VDD1.n16 1.93989
R1318 VDD1.n87 VDD1.n77 1.93989
R1319 VDD1.n121 VDD1.n61 1.93989
R1320 VDD1.n124 VDD1.t1 1.76521
R1321 VDD1.n124 VDD1.t3 1.76521
R1322 VDD1.n122 VDD1.t2 1.76521
R1323 VDD1.n122 VDD1.t0 1.76521
R1324 VDD1.n25 VDD1.n18 1.16414
R1325 VDD1.n86 VDD1.n79 1.16414
R1326 VDD1.n22 VDD1.n21 0.388379
R1327 VDD1.n83 VDD1.n82 0.388379
R1328 VDD1 VDD1.n125 0.185845
R1329 VDD1.n56 VDD1.n55 0.155672
R1330 VDD1.n55 VDD1.n3 0.155672
R1331 VDD1.n48 VDD1.n3 0.155672
R1332 VDD1.n48 VDD1.n47 0.155672
R1333 VDD1.n47 VDD1.n7 0.155672
R1334 VDD1.n40 VDD1.n7 0.155672
R1335 VDD1.n40 VDD1.n39 0.155672
R1336 VDD1.n39 VDD1.n11 0.155672
R1337 VDD1.n32 VDD1.n11 0.155672
R1338 VDD1.n32 VDD1.n31 0.155672
R1339 VDD1.n31 VDD1.n15 0.155672
R1340 VDD1.n24 VDD1.n15 0.155672
R1341 VDD1.n24 VDD1.n23 0.155672
R1342 VDD1.n85 VDD1.n84 0.155672
R1343 VDD1.n85 VDD1.n76 0.155672
R1344 VDD1.n92 VDD1.n76 0.155672
R1345 VDD1.n93 VDD1.n92 0.155672
R1346 VDD1.n93 VDD1.n72 0.155672
R1347 VDD1.n100 VDD1.n72 0.155672
R1348 VDD1.n101 VDD1.n100 0.155672
R1349 VDD1.n101 VDD1.n68 0.155672
R1350 VDD1.n108 VDD1.n68 0.155672
R1351 VDD1.n109 VDD1.n108 0.155672
R1352 VDD1.n109 VDD1.n64 0.155672
R1353 VDD1.n116 VDD1.n64 0.155672
R1354 VDD1.n117 VDD1.n116 0.155672
R1355 VTAIL.n254 VTAIL.n253 289.615
R1356 VTAIL.n62 VTAIL.n61 289.615
R1357 VTAIL.n192 VTAIL.n191 289.615
R1358 VTAIL.n128 VTAIL.n127 289.615
R1359 VTAIL.n215 VTAIL.n214 185
R1360 VTAIL.n212 VTAIL.n211 185
R1361 VTAIL.n221 VTAIL.n220 185
R1362 VTAIL.n223 VTAIL.n222 185
R1363 VTAIL.n208 VTAIL.n207 185
R1364 VTAIL.n229 VTAIL.n228 185
R1365 VTAIL.n231 VTAIL.n230 185
R1366 VTAIL.n204 VTAIL.n203 185
R1367 VTAIL.n237 VTAIL.n236 185
R1368 VTAIL.n239 VTAIL.n238 185
R1369 VTAIL.n200 VTAIL.n199 185
R1370 VTAIL.n245 VTAIL.n244 185
R1371 VTAIL.n247 VTAIL.n246 185
R1372 VTAIL.n196 VTAIL.n195 185
R1373 VTAIL.n253 VTAIL.n252 185
R1374 VTAIL.n23 VTAIL.n22 185
R1375 VTAIL.n20 VTAIL.n19 185
R1376 VTAIL.n29 VTAIL.n28 185
R1377 VTAIL.n31 VTAIL.n30 185
R1378 VTAIL.n16 VTAIL.n15 185
R1379 VTAIL.n37 VTAIL.n36 185
R1380 VTAIL.n39 VTAIL.n38 185
R1381 VTAIL.n12 VTAIL.n11 185
R1382 VTAIL.n45 VTAIL.n44 185
R1383 VTAIL.n47 VTAIL.n46 185
R1384 VTAIL.n8 VTAIL.n7 185
R1385 VTAIL.n53 VTAIL.n52 185
R1386 VTAIL.n55 VTAIL.n54 185
R1387 VTAIL.n4 VTAIL.n3 185
R1388 VTAIL.n61 VTAIL.n60 185
R1389 VTAIL.n191 VTAIL.n190 185
R1390 VTAIL.n134 VTAIL.n133 185
R1391 VTAIL.n185 VTAIL.n184 185
R1392 VTAIL.n183 VTAIL.n182 185
R1393 VTAIL.n138 VTAIL.n137 185
R1394 VTAIL.n177 VTAIL.n176 185
R1395 VTAIL.n175 VTAIL.n174 185
R1396 VTAIL.n142 VTAIL.n141 185
R1397 VTAIL.n169 VTAIL.n168 185
R1398 VTAIL.n167 VTAIL.n166 185
R1399 VTAIL.n146 VTAIL.n145 185
R1400 VTAIL.n161 VTAIL.n160 185
R1401 VTAIL.n159 VTAIL.n158 185
R1402 VTAIL.n150 VTAIL.n149 185
R1403 VTAIL.n153 VTAIL.n152 185
R1404 VTAIL.n127 VTAIL.n126 185
R1405 VTAIL.n70 VTAIL.n69 185
R1406 VTAIL.n121 VTAIL.n120 185
R1407 VTAIL.n119 VTAIL.n118 185
R1408 VTAIL.n74 VTAIL.n73 185
R1409 VTAIL.n113 VTAIL.n112 185
R1410 VTAIL.n111 VTAIL.n110 185
R1411 VTAIL.n78 VTAIL.n77 185
R1412 VTAIL.n105 VTAIL.n104 185
R1413 VTAIL.n103 VTAIL.n102 185
R1414 VTAIL.n82 VTAIL.n81 185
R1415 VTAIL.n97 VTAIL.n96 185
R1416 VTAIL.n95 VTAIL.n94 185
R1417 VTAIL.n86 VTAIL.n85 185
R1418 VTAIL.n89 VTAIL.n88 185
R1419 VTAIL.t0 VTAIL.n213 147.659
R1420 VTAIL.t9 VTAIL.n21 147.659
R1421 VTAIL.t8 VTAIL.n151 147.659
R1422 VTAIL.t5 VTAIL.n87 147.659
R1423 VTAIL.n214 VTAIL.n211 104.615
R1424 VTAIL.n221 VTAIL.n211 104.615
R1425 VTAIL.n222 VTAIL.n221 104.615
R1426 VTAIL.n222 VTAIL.n207 104.615
R1427 VTAIL.n229 VTAIL.n207 104.615
R1428 VTAIL.n230 VTAIL.n229 104.615
R1429 VTAIL.n230 VTAIL.n203 104.615
R1430 VTAIL.n237 VTAIL.n203 104.615
R1431 VTAIL.n238 VTAIL.n237 104.615
R1432 VTAIL.n238 VTAIL.n199 104.615
R1433 VTAIL.n245 VTAIL.n199 104.615
R1434 VTAIL.n246 VTAIL.n245 104.615
R1435 VTAIL.n246 VTAIL.n195 104.615
R1436 VTAIL.n253 VTAIL.n195 104.615
R1437 VTAIL.n22 VTAIL.n19 104.615
R1438 VTAIL.n29 VTAIL.n19 104.615
R1439 VTAIL.n30 VTAIL.n29 104.615
R1440 VTAIL.n30 VTAIL.n15 104.615
R1441 VTAIL.n37 VTAIL.n15 104.615
R1442 VTAIL.n38 VTAIL.n37 104.615
R1443 VTAIL.n38 VTAIL.n11 104.615
R1444 VTAIL.n45 VTAIL.n11 104.615
R1445 VTAIL.n46 VTAIL.n45 104.615
R1446 VTAIL.n46 VTAIL.n7 104.615
R1447 VTAIL.n53 VTAIL.n7 104.615
R1448 VTAIL.n54 VTAIL.n53 104.615
R1449 VTAIL.n54 VTAIL.n3 104.615
R1450 VTAIL.n61 VTAIL.n3 104.615
R1451 VTAIL.n191 VTAIL.n133 104.615
R1452 VTAIL.n184 VTAIL.n133 104.615
R1453 VTAIL.n184 VTAIL.n183 104.615
R1454 VTAIL.n183 VTAIL.n137 104.615
R1455 VTAIL.n176 VTAIL.n137 104.615
R1456 VTAIL.n176 VTAIL.n175 104.615
R1457 VTAIL.n175 VTAIL.n141 104.615
R1458 VTAIL.n168 VTAIL.n141 104.615
R1459 VTAIL.n168 VTAIL.n167 104.615
R1460 VTAIL.n167 VTAIL.n145 104.615
R1461 VTAIL.n160 VTAIL.n145 104.615
R1462 VTAIL.n160 VTAIL.n159 104.615
R1463 VTAIL.n159 VTAIL.n149 104.615
R1464 VTAIL.n152 VTAIL.n149 104.615
R1465 VTAIL.n127 VTAIL.n69 104.615
R1466 VTAIL.n120 VTAIL.n69 104.615
R1467 VTAIL.n120 VTAIL.n119 104.615
R1468 VTAIL.n119 VTAIL.n73 104.615
R1469 VTAIL.n112 VTAIL.n73 104.615
R1470 VTAIL.n112 VTAIL.n111 104.615
R1471 VTAIL.n111 VTAIL.n77 104.615
R1472 VTAIL.n104 VTAIL.n77 104.615
R1473 VTAIL.n104 VTAIL.n103 104.615
R1474 VTAIL.n103 VTAIL.n81 104.615
R1475 VTAIL.n96 VTAIL.n81 104.615
R1476 VTAIL.n96 VTAIL.n95 104.615
R1477 VTAIL.n95 VTAIL.n85 104.615
R1478 VTAIL.n88 VTAIL.n85 104.615
R1479 VTAIL.n214 VTAIL.t0 52.3082
R1480 VTAIL.n22 VTAIL.t9 52.3082
R1481 VTAIL.n152 VTAIL.t8 52.3082
R1482 VTAIL.n88 VTAIL.t5 52.3082
R1483 VTAIL.n131 VTAIL.n130 48.1967
R1484 VTAIL.n67 VTAIL.n66 48.1967
R1485 VTAIL.n1 VTAIL.n0 48.1965
R1486 VTAIL.n65 VTAIL.n64 48.1965
R1487 VTAIL.n255 VTAIL.n254 33.7369
R1488 VTAIL.n63 VTAIL.n62 33.7369
R1489 VTAIL.n193 VTAIL.n192 33.7369
R1490 VTAIL.n129 VTAIL.n128 33.7369
R1491 VTAIL.n67 VTAIL.n65 23.9876
R1492 VTAIL.n255 VTAIL.n193 23.0134
R1493 VTAIL.n215 VTAIL.n213 15.6677
R1494 VTAIL.n23 VTAIL.n21 15.6677
R1495 VTAIL.n153 VTAIL.n151 15.6677
R1496 VTAIL.n89 VTAIL.n87 15.6677
R1497 VTAIL.n216 VTAIL.n212 12.8005
R1498 VTAIL.n24 VTAIL.n20 12.8005
R1499 VTAIL.n154 VTAIL.n150 12.8005
R1500 VTAIL.n90 VTAIL.n86 12.8005
R1501 VTAIL.n220 VTAIL.n219 12.0247
R1502 VTAIL.n28 VTAIL.n27 12.0247
R1503 VTAIL.n158 VTAIL.n157 12.0247
R1504 VTAIL.n94 VTAIL.n93 12.0247
R1505 VTAIL.n223 VTAIL.n210 11.249
R1506 VTAIL.n252 VTAIL.n194 11.249
R1507 VTAIL.n31 VTAIL.n18 11.249
R1508 VTAIL.n60 VTAIL.n2 11.249
R1509 VTAIL.n190 VTAIL.n132 11.249
R1510 VTAIL.n161 VTAIL.n148 11.249
R1511 VTAIL.n126 VTAIL.n68 11.249
R1512 VTAIL.n97 VTAIL.n84 11.249
R1513 VTAIL.n224 VTAIL.n208 10.4732
R1514 VTAIL.n251 VTAIL.n196 10.4732
R1515 VTAIL.n32 VTAIL.n16 10.4732
R1516 VTAIL.n59 VTAIL.n4 10.4732
R1517 VTAIL.n189 VTAIL.n134 10.4732
R1518 VTAIL.n162 VTAIL.n146 10.4732
R1519 VTAIL.n125 VTAIL.n70 10.4732
R1520 VTAIL.n98 VTAIL.n82 10.4732
R1521 VTAIL.n228 VTAIL.n227 9.69747
R1522 VTAIL.n248 VTAIL.n247 9.69747
R1523 VTAIL.n36 VTAIL.n35 9.69747
R1524 VTAIL.n56 VTAIL.n55 9.69747
R1525 VTAIL.n186 VTAIL.n185 9.69747
R1526 VTAIL.n166 VTAIL.n165 9.69747
R1527 VTAIL.n122 VTAIL.n121 9.69747
R1528 VTAIL.n102 VTAIL.n101 9.69747
R1529 VTAIL.n250 VTAIL.n194 9.45567
R1530 VTAIL.n58 VTAIL.n2 9.45567
R1531 VTAIL.n188 VTAIL.n132 9.45567
R1532 VTAIL.n124 VTAIL.n68 9.45567
R1533 VTAIL.n202 VTAIL.n201 9.3005
R1534 VTAIL.n241 VTAIL.n240 9.3005
R1535 VTAIL.n243 VTAIL.n242 9.3005
R1536 VTAIL.n198 VTAIL.n197 9.3005
R1537 VTAIL.n249 VTAIL.n248 9.3005
R1538 VTAIL.n251 VTAIL.n250 9.3005
R1539 VTAIL.n233 VTAIL.n232 9.3005
R1540 VTAIL.n206 VTAIL.n205 9.3005
R1541 VTAIL.n227 VTAIL.n226 9.3005
R1542 VTAIL.n225 VTAIL.n224 9.3005
R1543 VTAIL.n210 VTAIL.n209 9.3005
R1544 VTAIL.n219 VTAIL.n218 9.3005
R1545 VTAIL.n217 VTAIL.n216 9.3005
R1546 VTAIL.n235 VTAIL.n234 9.3005
R1547 VTAIL.n10 VTAIL.n9 9.3005
R1548 VTAIL.n49 VTAIL.n48 9.3005
R1549 VTAIL.n51 VTAIL.n50 9.3005
R1550 VTAIL.n6 VTAIL.n5 9.3005
R1551 VTAIL.n57 VTAIL.n56 9.3005
R1552 VTAIL.n59 VTAIL.n58 9.3005
R1553 VTAIL.n41 VTAIL.n40 9.3005
R1554 VTAIL.n14 VTAIL.n13 9.3005
R1555 VTAIL.n35 VTAIL.n34 9.3005
R1556 VTAIL.n33 VTAIL.n32 9.3005
R1557 VTAIL.n18 VTAIL.n17 9.3005
R1558 VTAIL.n27 VTAIL.n26 9.3005
R1559 VTAIL.n25 VTAIL.n24 9.3005
R1560 VTAIL.n43 VTAIL.n42 9.3005
R1561 VTAIL.n189 VTAIL.n188 9.3005
R1562 VTAIL.n187 VTAIL.n186 9.3005
R1563 VTAIL.n136 VTAIL.n135 9.3005
R1564 VTAIL.n181 VTAIL.n180 9.3005
R1565 VTAIL.n179 VTAIL.n178 9.3005
R1566 VTAIL.n140 VTAIL.n139 9.3005
R1567 VTAIL.n173 VTAIL.n172 9.3005
R1568 VTAIL.n171 VTAIL.n170 9.3005
R1569 VTAIL.n144 VTAIL.n143 9.3005
R1570 VTAIL.n165 VTAIL.n164 9.3005
R1571 VTAIL.n163 VTAIL.n162 9.3005
R1572 VTAIL.n148 VTAIL.n147 9.3005
R1573 VTAIL.n157 VTAIL.n156 9.3005
R1574 VTAIL.n155 VTAIL.n154 9.3005
R1575 VTAIL.n115 VTAIL.n114 9.3005
R1576 VTAIL.n117 VTAIL.n116 9.3005
R1577 VTAIL.n72 VTAIL.n71 9.3005
R1578 VTAIL.n123 VTAIL.n122 9.3005
R1579 VTAIL.n125 VTAIL.n124 9.3005
R1580 VTAIL.n76 VTAIL.n75 9.3005
R1581 VTAIL.n109 VTAIL.n108 9.3005
R1582 VTAIL.n107 VTAIL.n106 9.3005
R1583 VTAIL.n80 VTAIL.n79 9.3005
R1584 VTAIL.n101 VTAIL.n100 9.3005
R1585 VTAIL.n99 VTAIL.n98 9.3005
R1586 VTAIL.n84 VTAIL.n83 9.3005
R1587 VTAIL.n93 VTAIL.n92 9.3005
R1588 VTAIL.n91 VTAIL.n90 9.3005
R1589 VTAIL.n231 VTAIL.n206 8.92171
R1590 VTAIL.n244 VTAIL.n198 8.92171
R1591 VTAIL.n39 VTAIL.n14 8.92171
R1592 VTAIL.n52 VTAIL.n6 8.92171
R1593 VTAIL.n182 VTAIL.n136 8.92171
R1594 VTAIL.n169 VTAIL.n144 8.92171
R1595 VTAIL.n118 VTAIL.n72 8.92171
R1596 VTAIL.n105 VTAIL.n80 8.92171
R1597 VTAIL.n232 VTAIL.n204 8.14595
R1598 VTAIL.n243 VTAIL.n200 8.14595
R1599 VTAIL.n40 VTAIL.n12 8.14595
R1600 VTAIL.n51 VTAIL.n8 8.14595
R1601 VTAIL.n181 VTAIL.n138 8.14595
R1602 VTAIL.n170 VTAIL.n142 8.14595
R1603 VTAIL.n117 VTAIL.n74 8.14595
R1604 VTAIL.n106 VTAIL.n78 8.14595
R1605 VTAIL.n236 VTAIL.n235 7.3702
R1606 VTAIL.n240 VTAIL.n239 7.3702
R1607 VTAIL.n44 VTAIL.n43 7.3702
R1608 VTAIL.n48 VTAIL.n47 7.3702
R1609 VTAIL.n178 VTAIL.n177 7.3702
R1610 VTAIL.n174 VTAIL.n173 7.3702
R1611 VTAIL.n114 VTAIL.n113 7.3702
R1612 VTAIL.n110 VTAIL.n109 7.3702
R1613 VTAIL.n236 VTAIL.n202 6.59444
R1614 VTAIL.n239 VTAIL.n202 6.59444
R1615 VTAIL.n44 VTAIL.n10 6.59444
R1616 VTAIL.n47 VTAIL.n10 6.59444
R1617 VTAIL.n177 VTAIL.n140 6.59444
R1618 VTAIL.n174 VTAIL.n140 6.59444
R1619 VTAIL.n113 VTAIL.n76 6.59444
R1620 VTAIL.n110 VTAIL.n76 6.59444
R1621 VTAIL.n235 VTAIL.n204 5.81868
R1622 VTAIL.n240 VTAIL.n200 5.81868
R1623 VTAIL.n43 VTAIL.n12 5.81868
R1624 VTAIL.n48 VTAIL.n8 5.81868
R1625 VTAIL.n178 VTAIL.n138 5.81868
R1626 VTAIL.n173 VTAIL.n142 5.81868
R1627 VTAIL.n114 VTAIL.n74 5.81868
R1628 VTAIL.n109 VTAIL.n78 5.81868
R1629 VTAIL.n232 VTAIL.n231 5.04292
R1630 VTAIL.n244 VTAIL.n243 5.04292
R1631 VTAIL.n40 VTAIL.n39 5.04292
R1632 VTAIL.n52 VTAIL.n51 5.04292
R1633 VTAIL.n182 VTAIL.n181 5.04292
R1634 VTAIL.n170 VTAIL.n169 5.04292
R1635 VTAIL.n118 VTAIL.n117 5.04292
R1636 VTAIL.n106 VTAIL.n105 5.04292
R1637 VTAIL.n217 VTAIL.n213 4.38563
R1638 VTAIL.n25 VTAIL.n21 4.38563
R1639 VTAIL.n155 VTAIL.n151 4.38563
R1640 VTAIL.n91 VTAIL.n87 4.38563
R1641 VTAIL.n228 VTAIL.n206 4.26717
R1642 VTAIL.n247 VTAIL.n198 4.26717
R1643 VTAIL.n36 VTAIL.n14 4.26717
R1644 VTAIL.n55 VTAIL.n6 4.26717
R1645 VTAIL.n185 VTAIL.n136 4.26717
R1646 VTAIL.n166 VTAIL.n144 4.26717
R1647 VTAIL.n121 VTAIL.n72 4.26717
R1648 VTAIL.n102 VTAIL.n80 4.26717
R1649 VTAIL.n227 VTAIL.n208 3.49141
R1650 VTAIL.n248 VTAIL.n196 3.49141
R1651 VTAIL.n35 VTAIL.n16 3.49141
R1652 VTAIL.n56 VTAIL.n4 3.49141
R1653 VTAIL.n186 VTAIL.n134 3.49141
R1654 VTAIL.n165 VTAIL.n146 3.49141
R1655 VTAIL.n122 VTAIL.n70 3.49141
R1656 VTAIL.n101 VTAIL.n82 3.49141
R1657 VTAIL.n224 VTAIL.n223 2.71565
R1658 VTAIL.n252 VTAIL.n251 2.71565
R1659 VTAIL.n32 VTAIL.n31 2.71565
R1660 VTAIL.n60 VTAIL.n59 2.71565
R1661 VTAIL.n190 VTAIL.n189 2.71565
R1662 VTAIL.n162 VTAIL.n161 2.71565
R1663 VTAIL.n126 VTAIL.n125 2.71565
R1664 VTAIL.n98 VTAIL.n97 2.71565
R1665 VTAIL.n220 VTAIL.n210 1.93989
R1666 VTAIL.n254 VTAIL.n194 1.93989
R1667 VTAIL.n28 VTAIL.n18 1.93989
R1668 VTAIL.n62 VTAIL.n2 1.93989
R1669 VTAIL.n192 VTAIL.n132 1.93989
R1670 VTAIL.n158 VTAIL.n148 1.93989
R1671 VTAIL.n128 VTAIL.n68 1.93989
R1672 VTAIL.n94 VTAIL.n84 1.93989
R1673 VTAIL.n0 VTAIL.t4 1.76521
R1674 VTAIL.n0 VTAIL.t3 1.76521
R1675 VTAIL.n64 VTAIL.t10 1.76521
R1676 VTAIL.n64 VTAIL.t11 1.76521
R1677 VTAIL.n130 VTAIL.t6 1.76521
R1678 VTAIL.n130 VTAIL.t7 1.76521
R1679 VTAIL.n66 VTAIL.t2 1.76521
R1680 VTAIL.n66 VTAIL.t1 1.76521
R1681 VTAIL.n219 VTAIL.n212 1.16414
R1682 VTAIL.n27 VTAIL.n20 1.16414
R1683 VTAIL.n157 VTAIL.n150 1.16414
R1684 VTAIL.n93 VTAIL.n86 1.16414
R1685 VTAIL.n129 VTAIL.n67 0.974638
R1686 VTAIL.n193 VTAIL.n131 0.974638
R1687 VTAIL.n65 VTAIL.n63 0.974638
R1688 VTAIL.n131 VTAIL.n129 0.957397
R1689 VTAIL.n63 VTAIL.n1 0.957397
R1690 VTAIL VTAIL.n255 0.672914
R1691 VTAIL.n216 VTAIL.n215 0.388379
R1692 VTAIL.n24 VTAIL.n23 0.388379
R1693 VTAIL.n154 VTAIL.n153 0.388379
R1694 VTAIL.n90 VTAIL.n89 0.388379
R1695 VTAIL VTAIL.n1 0.302224
R1696 VTAIL.n218 VTAIL.n217 0.155672
R1697 VTAIL.n218 VTAIL.n209 0.155672
R1698 VTAIL.n225 VTAIL.n209 0.155672
R1699 VTAIL.n226 VTAIL.n225 0.155672
R1700 VTAIL.n226 VTAIL.n205 0.155672
R1701 VTAIL.n233 VTAIL.n205 0.155672
R1702 VTAIL.n234 VTAIL.n233 0.155672
R1703 VTAIL.n234 VTAIL.n201 0.155672
R1704 VTAIL.n241 VTAIL.n201 0.155672
R1705 VTAIL.n242 VTAIL.n241 0.155672
R1706 VTAIL.n242 VTAIL.n197 0.155672
R1707 VTAIL.n249 VTAIL.n197 0.155672
R1708 VTAIL.n250 VTAIL.n249 0.155672
R1709 VTAIL.n26 VTAIL.n25 0.155672
R1710 VTAIL.n26 VTAIL.n17 0.155672
R1711 VTAIL.n33 VTAIL.n17 0.155672
R1712 VTAIL.n34 VTAIL.n33 0.155672
R1713 VTAIL.n34 VTAIL.n13 0.155672
R1714 VTAIL.n41 VTAIL.n13 0.155672
R1715 VTAIL.n42 VTAIL.n41 0.155672
R1716 VTAIL.n42 VTAIL.n9 0.155672
R1717 VTAIL.n49 VTAIL.n9 0.155672
R1718 VTAIL.n50 VTAIL.n49 0.155672
R1719 VTAIL.n50 VTAIL.n5 0.155672
R1720 VTAIL.n57 VTAIL.n5 0.155672
R1721 VTAIL.n58 VTAIL.n57 0.155672
R1722 VTAIL.n188 VTAIL.n187 0.155672
R1723 VTAIL.n187 VTAIL.n135 0.155672
R1724 VTAIL.n180 VTAIL.n135 0.155672
R1725 VTAIL.n180 VTAIL.n179 0.155672
R1726 VTAIL.n179 VTAIL.n139 0.155672
R1727 VTAIL.n172 VTAIL.n139 0.155672
R1728 VTAIL.n172 VTAIL.n171 0.155672
R1729 VTAIL.n171 VTAIL.n143 0.155672
R1730 VTAIL.n164 VTAIL.n143 0.155672
R1731 VTAIL.n164 VTAIL.n163 0.155672
R1732 VTAIL.n163 VTAIL.n147 0.155672
R1733 VTAIL.n156 VTAIL.n147 0.155672
R1734 VTAIL.n156 VTAIL.n155 0.155672
R1735 VTAIL.n124 VTAIL.n123 0.155672
R1736 VTAIL.n123 VTAIL.n71 0.155672
R1737 VTAIL.n116 VTAIL.n71 0.155672
R1738 VTAIL.n116 VTAIL.n115 0.155672
R1739 VTAIL.n115 VTAIL.n75 0.155672
R1740 VTAIL.n108 VTAIL.n75 0.155672
R1741 VTAIL.n108 VTAIL.n107 0.155672
R1742 VTAIL.n107 VTAIL.n79 0.155672
R1743 VTAIL.n100 VTAIL.n79 0.155672
R1744 VTAIL.n100 VTAIL.n99 0.155672
R1745 VTAIL.n99 VTAIL.n83 0.155672
R1746 VTAIL.n92 VTAIL.n83 0.155672
R1747 VTAIL.n92 VTAIL.n91 0.155672
R1748 VN.n1 VN.t5 411.195
R1749 VN.n7 VN.t4 411.195
R1750 VN.n2 VN.t0 387.709
R1751 VN.n4 VN.t3 387.709
R1752 VN.n8 VN.t2 387.709
R1753 VN.n10 VN.t1 387.709
R1754 VN.n5 VN.n4 161.3
R1755 VN.n11 VN.n10 161.3
R1756 VN.n9 VN.n6 161.3
R1757 VN.n3 VN.n0 161.3
R1758 VN.n7 VN.n6 44.8973
R1759 VN.n1 VN.n0 44.8973
R1760 VN VN.n11 41.4835
R1761 VN.n4 VN.n3 33.5944
R1762 VN.n10 VN.n9 33.5944
R1763 VN.n2 VN.n1 18.1882
R1764 VN.n8 VN.n7 18.1882
R1765 VN.n3 VN.n2 14.6066
R1766 VN.n9 VN.n8 14.6066
R1767 VN.n11 VN.n6 0.189894
R1768 VN.n5 VN.n0 0.189894
R1769 VN VN.n5 0.0516364
R1770 VDD2.n123 VDD2.n122 289.615
R1771 VDD2.n60 VDD2.n59 289.615
R1772 VDD2.n122 VDD2.n121 185
R1773 VDD2.n65 VDD2.n64 185
R1774 VDD2.n116 VDD2.n115 185
R1775 VDD2.n114 VDD2.n113 185
R1776 VDD2.n69 VDD2.n68 185
R1777 VDD2.n108 VDD2.n107 185
R1778 VDD2.n106 VDD2.n105 185
R1779 VDD2.n73 VDD2.n72 185
R1780 VDD2.n100 VDD2.n99 185
R1781 VDD2.n98 VDD2.n97 185
R1782 VDD2.n77 VDD2.n76 185
R1783 VDD2.n92 VDD2.n91 185
R1784 VDD2.n90 VDD2.n89 185
R1785 VDD2.n81 VDD2.n80 185
R1786 VDD2.n84 VDD2.n83 185
R1787 VDD2.n21 VDD2.n20 185
R1788 VDD2.n18 VDD2.n17 185
R1789 VDD2.n27 VDD2.n26 185
R1790 VDD2.n29 VDD2.n28 185
R1791 VDD2.n14 VDD2.n13 185
R1792 VDD2.n35 VDD2.n34 185
R1793 VDD2.n37 VDD2.n36 185
R1794 VDD2.n10 VDD2.n9 185
R1795 VDD2.n43 VDD2.n42 185
R1796 VDD2.n45 VDD2.n44 185
R1797 VDD2.n6 VDD2.n5 185
R1798 VDD2.n51 VDD2.n50 185
R1799 VDD2.n53 VDD2.n52 185
R1800 VDD2.n2 VDD2.n1 185
R1801 VDD2.n59 VDD2.n58 185
R1802 VDD2.t0 VDD2.n19 147.659
R1803 VDD2.t4 VDD2.n82 147.659
R1804 VDD2.n122 VDD2.n64 104.615
R1805 VDD2.n115 VDD2.n64 104.615
R1806 VDD2.n115 VDD2.n114 104.615
R1807 VDD2.n114 VDD2.n68 104.615
R1808 VDD2.n107 VDD2.n68 104.615
R1809 VDD2.n107 VDD2.n106 104.615
R1810 VDD2.n106 VDD2.n72 104.615
R1811 VDD2.n99 VDD2.n72 104.615
R1812 VDD2.n99 VDD2.n98 104.615
R1813 VDD2.n98 VDD2.n76 104.615
R1814 VDD2.n91 VDD2.n76 104.615
R1815 VDD2.n91 VDD2.n90 104.615
R1816 VDD2.n90 VDD2.n80 104.615
R1817 VDD2.n83 VDD2.n80 104.615
R1818 VDD2.n20 VDD2.n17 104.615
R1819 VDD2.n27 VDD2.n17 104.615
R1820 VDD2.n28 VDD2.n27 104.615
R1821 VDD2.n28 VDD2.n13 104.615
R1822 VDD2.n35 VDD2.n13 104.615
R1823 VDD2.n36 VDD2.n35 104.615
R1824 VDD2.n36 VDD2.n9 104.615
R1825 VDD2.n43 VDD2.n9 104.615
R1826 VDD2.n44 VDD2.n43 104.615
R1827 VDD2.n44 VDD2.n5 104.615
R1828 VDD2.n51 VDD2.n5 104.615
R1829 VDD2.n52 VDD2.n51 104.615
R1830 VDD2.n52 VDD2.n1 104.615
R1831 VDD2.n59 VDD2.n1 104.615
R1832 VDD2.n62 VDD2.n61 65.0635
R1833 VDD2 VDD2.n125 65.0598
R1834 VDD2.n83 VDD2.t4 52.3082
R1835 VDD2.n20 VDD2.t0 52.3082
R1836 VDD2.n62 VDD2.n60 51.0909
R1837 VDD2.n124 VDD2.n123 50.4157
R1838 VDD2.n124 VDD2.n62 36.5537
R1839 VDD2.n84 VDD2.n82 15.6677
R1840 VDD2.n21 VDD2.n19 15.6677
R1841 VDD2.n85 VDD2.n81 12.8005
R1842 VDD2.n22 VDD2.n18 12.8005
R1843 VDD2.n89 VDD2.n88 12.0247
R1844 VDD2.n26 VDD2.n25 12.0247
R1845 VDD2.n121 VDD2.n63 11.249
R1846 VDD2.n92 VDD2.n79 11.249
R1847 VDD2.n29 VDD2.n16 11.249
R1848 VDD2.n58 VDD2.n0 11.249
R1849 VDD2.n120 VDD2.n65 10.4732
R1850 VDD2.n93 VDD2.n77 10.4732
R1851 VDD2.n30 VDD2.n14 10.4732
R1852 VDD2.n57 VDD2.n2 10.4732
R1853 VDD2.n117 VDD2.n116 9.69747
R1854 VDD2.n97 VDD2.n96 9.69747
R1855 VDD2.n34 VDD2.n33 9.69747
R1856 VDD2.n54 VDD2.n53 9.69747
R1857 VDD2.n119 VDD2.n63 9.45567
R1858 VDD2.n56 VDD2.n0 9.45567
R1859 VDD2.n110 VDD2.n109 9.3005
R1860 VDD2.n112 VDD2.n111 9.3005
R1861 VDD2.n67 VDD2.n66 9.3005
R1862 VDD2.n118 VDD2.n117 9.3005
R1863 VDD2.n120 VDD2.n119 9.3005
R1864 VDD2.n71 VDD2.n70 9.3005
R1865 VDD2.n104 VDD2.n103 9.3005
R1866 VDD2.n102 VDD2.n101 9.3005
R1867 VDD2.n75 VDD2.n74 9.3005
R1868 VDD2.n96 VDD2.n95 9.3005
R1869 VDD2.n94 VDD2.n93 9.3005
R1870 VDD2.n79 VDD2.n78 9.3005
R1871 VDD2.n88 VDD2.n87 9.3005
R1872 VDD2.n86 VDD2.n85 9.3005
R1873 VDD2.n8 VDD2.n7 9.3005
R1874 VDD2.n47 VDD2.n46 9.3005
R1875 VDD2.n49 VDD2.n48 9.3005
R1876 VDD2.n4 VDD2.n3 9.3005
R1877 VDD2.n55 VDD2.n54 9.3005
R1878 VDD2.n57 VDD2.n56 9.3005
R1879 VDD2.n39 VDD2.n38 9.3005
R1880 VDD2.n12 VDD2.n11 9.3005
R1881 VDD2.n33 VDD2.n32 9.3005
R1882 VDD2.n31 VDD2.n30 9.3005
R1883 VDD2.n16 VDD2.n15 9.3005
R1884 VDD2.n25 VDD2.n24 9.3005
R1885 VDD2.n23 VDD2.n22 9.3005
R1886 VDD2.n41 VDD2.n40 9.3005
R1887 VDD2.n113 VDD2.n67 8.92171
R1888 VDD2.n100 VDD2.n75 8.92171
R1889 VDD2.n37 VDD2.n12 8.92171
R1890 VDD2.n50 VDD2.n4 8.92171
R1891 VDD2.n112 VDD2.n69 8.14595
R1892 VDD2.n101 VDD2.n73 8.14595
R1893 VDD2.n38 VDD2.n10 8.14595
R1894 VDD2.n49 VDD2.n6 8.14595
R1895 VDD2.n109 VDD2.n108 7.3702
R1896 VDD2.n105 VDD2.n104 7.3702
R1897 VDD2.n42 VDD2.n41 7.3702
R1898 VDD2.n46 VDD2.n45 7.3702
R1899 VDD2.n108 VDD2.n71 6.59444
R1900 VDD2.n105 VDD2.n71 6.59444
R1901 VDD2.n42 VDD2.n8 6.59444
R1902 VDD2.n45 VDD2.n8 6.59444
R1903 VDD2.n109 VDD2.n69 5.81868
R1904 VDD2.n104 VDD2.n73 5.81868
R1905 VDD2.n41 VDD2.n10 5.81868
R1906 VDD2.n46 VDD2.n6 5.81868
R1907 VDD2.n113 VDD2.n112 5.04292
R1908 VDD2.n101 VDD2.n100 5.04292
R1909 VDD2.n38 VDD2.n37 5.04292
R1910 VDD2.n50 VDD2.n49 5.04292
R1911 VDD2.n23 VDD2.n19 4.38563
R1912 VDD2.n86 VDD2.n82 4.38563
R1913 VDD2.n116 VDD2.n67 4.26717
R1914 VDD2.n97 VDD2.n75 4.26717
R1915 VDD2.n34 VDD2.n12 4.26717
R1916 VDD2.n53 VDD2.n4 4.26717
R1917 VDD2.n117 VDD2.n65 3.49141
R1918 VDD2.n96 VDD2.n77 3.49141
R1919 VDD2.n33 VDD2.n14 3.49141
R1920 VDD2.n54 VDD2.n2 3.49141
R1921 VDD2.n121 VDD2.n120 2.71565
R1922 VDD2.n93 VDD2.n92 2.71565
R1923 VDD2.n30 VDD2.n29 2.71565
R1924 VDD2.n58 VDD2.n57 2.71565
R1925 VDD2.n123 VDD2.n63 1.93989
R1926 VDD2.n89 VDD2.n79 1.93989
R1927 VDD2.n26 VDD2.n16 1.93989
R1928 VDD2.n60 VDD2.n0 1.93989
R1929 VDD2.n125 VDD2.t3 1.76521
R1930 VDD2.n125 VDD2.t1 1.76521
R1931 VDD2.n61 VDD2.t5 1.76521
R1932 VDD2.n61 VDD2.t2 1.76521
R1933 VDD2.n88 VDD2.n81 1.16414
R1934 VDD2.n25 VDD2.n18 1.16414
R1935 VDD2 VDD2.n124 0.789293
R1936 VDD2.n85 VDD2.n84 0.388379
R1937 VDD2.n22 VDD2.n21 0.388379
R1938 VDD2.n119 VDD2.n118 0.155672
R1939 VDD2.n118 VDD2.n66 0.155672
R1940 VDD2.n111 VDD2.n66 0.155672
R1941 VDD2.n111 VDD2.n110 0.155672
R1942 VDD2.n110 VDD2.n70 0.155672
R1943 VDD2.n103 VDD2.n70 0.155672
R1944 VDD2.n103 VDD2.n102 0.155672
R1945 VDD2.n102 VDD2.n74 0.155672
R1946 VDD2.n95 VDD2.n74 0.155672
R1947 VDD2.n95 VDD2.n94 0.155672
R1948 VDD2.n94 VDD2.n78 0.155672
R1949 VDD2.n87 VDD2.n78 0.155672
R1950 VDD2.n87 VDD2.n86 0.155672
R1951 VDD2.n24 VDD2.n23 0.155672
R1952 VDD2.n24 VDD2.n15 0.155672
R1953 VDD2.n31 VDD2.n15 0.155672
R1954 VDD2.n32 VDD2.n31 0.155672
R1955 VDD2.n32 VDD2.n11 0.155672
R1956 VDD2.n39 VDD2.n11 0.155672
R1957 VDD2.n40 VDD2.n39 0.155672
R1958 VDD2.n40 VDD2.n7 0.155672
R1959 VDD2.n47 VDD2.n7 0.155672
R1960 VDD2.n48 VDD2.n47 0.155672
R1961 VDD2.n48 VDD2.n3 0.155672
R1962 VDD2.n55 VDD2.n3 0.155672
R1963 VDD2.n56 VDD2.n55 0.155672
C0 VP VN 5.03274f
C1 VDD2 VN 4.34428f
C2 VTAIL VP 4.10475f
C3 VTAIL VDD2 9.0145f
C4 VDD1 VP 4.49781f
C5 VDD1 VDD2 0.745955f
C6 VDD2 VP 0.305484f
C7 VTAIL VN 4.09021f
C8 VDD1 VN 0.147818f
C9 VTAIL VDD1 8.97897f
C10 VDD2 B 4.41881f
C11 VDD1 B 4.457129f
C12 VTAIL B 6.192194f
C13 VN B 7.87191f
C14 VP B 6.009953f
C15 VDD2.n0 B 0.012876f
C16 VDD2.n1 B 0.029029f
C17 VDD2.n2 B 0.013004f
C18 VDD2.n3 B 0.022856f
C19 VDD2.n4 B 0.012282f
C20 VDD2.n5 B 0.029029f
C21 VDD2.n6 B 0.013004f
C22 VDD2.n7 B 0.022856f
C23 VDD2.n8 B 0.012282f
C24 VDD2.n9 B 0.029029f
C25 VDD2.n10 B 0.013004f
C26 VDD2.n11 B 0.022856f
C27 VDD2.n12 B 0.012282f
C28 VDD2.n13 B 0.029029f
C29 VDD2.n14 B 0.013004f
C30 VDD2.n15 B 0.022856f
C31 VDD2.n16 B 0.012282f
C32 VDD2.n17 B 0.029029f
C33 VDD2.n18 B 0.013004f
C34 VDD2.n19 B 0.127409f
C35 VDD2.t0 B 0.04757f
C36 VDD2.n20 B 0.021772f
C37 VDD2.n21 B 0.017148f
C38 VDD2.n22 B 0.012282f
C39 VDD2.n23 B 1.09107f
C40 VDD2.n24 B 0.022856f
C41 VDD2.n25 B 0.012282f
C42 VDD2.n26 B 0.013004f
C43 VDD2.n27 B 0.029029f
C44 VDD2.n28 B 0.029029f
C45 VDD2.n29 B 0.013004f
C46 VDD2.n30 B 0.012282f
C47 VDD2.n31 B 0.022856f
C48 VDD2.n32 B 0.022856f
C49 VDD2.n33 B 0.012282f
C50 VDD2.n34 B 0.013004f
C51 VDD2.n35 B 0.029029f
C52 VDD2.n36 B 0.029029f
C53 VDD2.n37 B 0.013004f
C54 VDD2.n38 B 0.012282f
C55 VDD2.n39 B 0.022856f
C56 VDD2.n40 B 0.022856f
C57 VDD2.n41 B 0.012282f
C58 VDD2.n42 B 0.013004f
C59 VDD2.n43 B 0.029029f
C60 VDD2.n44 B 0.029029f
C61 VDD2.n45 B 0.013004f
C62 VDD2.n46 B 0.012282f
C63 VDD2.n47 B 0.022856f
C64 VDD2.n48 B 0.022856f
C65 VDD2.n49 B 0.012282f
C66 VDD2.n50 B 0.013004f
C67 VDD2.n51 B 0.029029f
C68 VDD2.n52 B 0.029029f
C69 VDD2.n53 B 0.013004f
C70 VDD2.n54 B 0.012282f
C71 VDD2.n55 B 0.022856f
C72 VDD2.n56 B 0.05845f
C73 VDD2.n57 B 0.012282f
C74 VDD2.n58 B 0.013004f
C75 VDD2.n59 B 0.056844f
C76 VDD2.n60 B 0.065289f
C77 VDD2.t5 B 0.202646f
C78 VDD2.t2 B 0.202646f
C79 VDD2.n61 B 1.80843f
C80 VDD2.n62 B 1.68223f
C81 VDD2.n63 B 0.012876f
C82 VDD2.n64 B 0.029029f
C83 VDD2.n65 B 0.013004f
C84 VDD2.n66 B 0.022856f
C85 VDD2.n67 B 0.012282f
C86 VDD2.n68 B 0.029029f
C87 VDD2.n69 B 0.013004f
C88 VDD2.n70 B 0.022856f
C89 VDD2.n71 B 0.012282f
C90 VDD2.n72 B 0.029029f
C91 VDD2.n73 B 0.013004f
C92 VDD2.n74 B 0.022856f
C93 VDD2.n75 B 0.012282f
C94 VDD2.n76 B 0.029029f
C95 VDD2.n77 B 0.013004f
C96 VDD2.n78 B 0.022856f
C97 VDD2.n79 B 0.012282f
C98 VDD2.n80 B 0.029029f
C99 VDD2.n81 B 0.013004f
C100 VDD2.n82 B 0.127409f
C101 VDD2.t4 B 0.04757f
C102 VDD2.n83 B 0.021772f
C103 VDD2.n84 B 0.017148f
C104 VDD2.n85 B 0.012282f
C105 VDD2.n86 B 1.09107f
C106 VDD2.n87 B 0.022856f
C107 VDD2.n88 B 0.012282f
C108 VDD2.n89 B 0.013004f
C109 VDD2.n90 B 0.029029f
C110 VDD2.n91 B 0.029029f
C111 VDD2.n92 B 0.013004f
C112 VDD2.n93 B 0.012282f
C113 VDD2.n94 B 0.022856f
C114 VDD2.n95 B 0.022856f
C115 VDD2.n96 B 0.012282f
C116 VDD2.n97 B 0.013004f
C117 VDD2.n98 B 0.029029f
C118 VDD2.n99 B 0.029029f
C119 VDD2.n100 B 0.013004f
C120 VDD2.n101 B 0.012282f
C121 VDD2.n102 B 0.022856f
C122 VDD2.n103 B 0.022856f
C123 VDD2.n104 B 0.012282f
C124 VDD2.n105 B 0.013004f
C125 VDD2.n106 B 0.029029f
C126 VDD2.n107 B 0.029029f
C127 VDD2.n108 B 0.013004f
C128 VDD2.n109 B 0.012282f
C129 VDD2.n110 B 0.022856f
C130 VDD2.n111 B 0.022856f
C131 VDD2.n112 B 0.012282f
C132 VDD2.n113 B 0.013004f
C133 VDD2.n114 B 0.029029f
C134 VDD2.n115 B 0.029029f
C135 VDD2.n116 B 0.013004f
C136 VDD2.n117 B 0.012282f
C137 VDD2.n118 B 0.022856f
C138 VDD2.n119 B 0.05845f
C139 VDD2.n120 B 0.012282f
C140 VDD2.n121 B 0.013004f
C141 VDD2.n122 B 0.056844f
C142 VDD2.n123 B 0.064021f
C143 VDD2.n124 B 1.83916f
C144 VDD2.t3 B 0.202646f
C145 VDD2.t1 B 0.202646f
C146 VDD2.n125 B 1.80842f
C147 VN.n0 B 0.18874f
C148 VN.t5 B 1.14505f
C149 VN.n1 B 0.428684f
C150 VN.t0 B 1.11932f
C151 VN.n2 B 0.452858f
C152 VN.n3 B 0.009906f
C153 VN.t3 B 1.11932f
C154 VN.n4 B 0.448613f
C155 VN.n5 B 0.03383f
C156 VN.n6 B 0.18874f
C157 VN.t4 B 1.14505f
C158 VN.n7 B 0.428684f
C159 VN.t2 B 1.11932f
C160 VN.n8 B 0.452858f
C161 VN.n9 B 0.009906f
C162 VN.t1 B 1.11932f
C163 VN.n10 B 0.448613f
C164 VN.n11 B 1.76649f
C165 VTAIL.t4 B 0.21364f
C166 VTAIL.t3 B 0.21364f
C167 VTAIL.n0 B 1.84208f
C168 VTAIL.n1 B 0.31702f
C169 VTAIL.n2 B 0.013574f
C170 VTAIL.n3 B 0.030604f
C171 VTAIL.n4 B 0.01371f
C172 VTAIL.n5 B 0.024096f
C173 VTAIL.n6 B 0.012948f
C174 VTAIL.n7 B 0.030604f
C175 VTAIL.n8 B 0.01371f
C176 VTAIL.n9 B 0.024096f
C177 VTAIL.n10 B 0.012948f
C178 VTAIL.n11 B 0.030604f
C179 VTAIL.n12 B 0.01371f
C180 VTAIL.n13 B 0.024096f
C181 VTAIL.n14 B 0.012948f
C182 VTAIL.n15 B 0.030604f
C183 VTAIL.n16 B 0.01371f
C184 VTAIL.n17 B 0.024096f
C185 VTAIL.n18 B 0.012948f
C186 VTAIL.n19 B 0.030604f
C187 VTAIL.n20 B 0.01371f
C188 VTAIL.n21 B 0.134321f
C189 VTAIL.t9 B 0.05015f
C190 VTAIL.n22 B 0.022953f
C191 VTAIL.n23 B 0.018079f
C192 VTAIL.n24 B 0.012948f
C193 VTAIL.n25 B 1.15026f
C194 VTAIL.n26 B 0.024096f
C195 VTAIL.n27 B 0.012948f
C196 VTAIL.n28 B 0.01371f
C197 VTAIL.n29 B 0.030604f
C198 VTAIL.n30 B 0.030604f
C199 VTAIL.n31 B 0.01371f
C200 VTAIL.n32 B 0.012948f
C201 VTAIL.n33 B 0.024096f
C202 VTAIL.n34 B 0.024096f
C203 VTAIL.n35 B 0.012948f
C204 VTAIL.n36 B 0.01371f
C205 VTAIL.n37 B 0.030604f
C206 VTAIL.n38 B 0.030604f
C207 VTAIL.n39 B 0.01371f
C208 VTAIL.n40 B 0.012948f
C209 VTAIL.n41 B 0.024096f
C210 VTAIL.n42 B 0.024096f
C211 VTAIL.n43 B 0.012948f
C212 VTAIL.n44 B 0.01371f
C213 VTAIL.n45 B 0.030604f
C214 VTAIL.n46 B 0.030604f
C215 VTAIL.n47 B 0.01371f
C216 VTAIL.n48 B 0.012948f
C217 VTAIL.n49 B 0.024096f
C218 VTAIL.n50 B 0.024096f
C219 VTAIL.n51 B 0.012948f
C220 VTAIL.n52 B 0.01371f
C221 VTAIL.n53 B 0.030604f
C222 VTAIL.n54 B 0.030604f
C223 VTAIL.n55 B 0.01371f
C224 VTAIL.n56 B 0.012948f
C225 VTAIL.n57 B 0.024096f
C226 VTAIL.n58 B 0.061621f
C227 VTAIL.n59 B 0.012948f
C228 VTAIL.n60 B 0.01371f
C229 VTAIL.n61 B 0.059928f
C230 VTAIL.n62 B 0.050876f
C231 VTAIL.n63 B 0.171995f
C232 VTAIL.t10 B 0.21364f
C233 VTAIL.t11 B 0.21364f
C234 VTAIL.n64 B 1.84208f
C235 VTAIL.n65 B 1.52449f
C236 VTAIL.t2 B 0.21364f
C237 VTAIL.t1 B 0.21364f
C238 VTAIL.n66 B 1.84209f
C239 VTAIL.n67 B 1.52448f
C240 VTAIL.n68 B 0.013574f
C241 VTAIL.n69 B 0.030604f
C242 VTAIL.n70 B 0.01371f
C243 VTAIL.n71 B 0.024096f
C244 VTAIL.n72 B 0.012948f
C245 VTAIL.n73 B 0.030604f
C246 VTAIL.n74 B 0.01371f
C247 VTAIL.n75 B 0.024096f
C248 VTAIL.n76 B 0.012948f
C249 VTAIL.n77 B 0.030604f
C250 VTAIL.n78 B 0.01371f
C251 VTAIL.n79 B 0.024096f
C252 VTAIL.n80 B 0.012948f
C253 VTAIL.n81 B 0.030604f
C254 VTAIL.n82 B 0.01371f
C255 VTAIL.n83 B 0.024096f
C256 VTAIL.n84 B 0.012948f
C257 VTAIL.n85 B 0.030604f
C258 VTAIL.n86 B 0.01371f
C259 VTAIL.n87 B 0.134321f
C260 VTAIL.t5 B 0.05015f
C261 VTAIL.n88 B 0.022953f
C262 VTAIL.n89 B 0.018079f
C263 VTAIL.n90 B 0.012948f
C264 VTAIL.n91 B 1.15026f
C265 VTAIL.n92 B 0.024096f
C266 VTAIL.n93 B 0.012948f
C267 VTAIL.n94 B 0.01371f
C268 VTAIL.n95 B 0.030604f
C269 VTAIL.n96 B 0.030604f
C270 VTAIL.n97 B 0.01371f
C271 VTAIL.n98 B 0.012948f
C272 VTAIL.n99 B 0.024096f
C273 VTAIL.n100 B 0.024096f
C274 VTAIL.n101 B 0.012948f
C275 VTAIL.n102 B 0.01371f
C276 VTAIL.n103 B 0.030604f
C277 VTAIL.n104 B 0.030604f
C278 VTAIL.n105 B 0.01371f
C279 VTAIL.n106 B 0.012948f
C280 VTAIL.n107 B 0.024096f
C281 VTAIL.n108 B 0.024096f
C282 VTAIL.n109 B 0.012948f
C283 VTAIL.n110 B 0.01371f
C284 VTAIL.n111 B 0.030604f
C285 VTAIL.n112 B 0.030604f
C286 VTAIL.n113 B 0.01371f
C287 VTAIL.n114 B 0.012948f
C288 VTAIL.n115 B 0.024096f
C289 VTAIL.n116 B 0.024096f
C290 VTAIL.n117 B 0.012948f
C291 VTAIL.n118 B 0.01371f
C292 VTAIL.n119 B 0.030604f
C293 VTAIL.n120 B 0.030604f
C294 VTAIL.n121 B 0.01371f
C295 VTAIL.n122 B 0.012948f
C296 VTAIL.n123 B 0.024096f
C297 VTAIL.n124 B 0.061621f
C298 VTAIL.n125 B 0.012948f
C299 VTAIL.n126 B 0.01371f
C300 VTAIL.n127 B 0.059928f
C301 VTAIL.n128 B 0.050876f
C302 VTAIL.n129 B 0.171995f
C303 VTAIL.t6 B 0.21364f
C304 VTAIL.t7 B 0.21364f
C305 VTAIL.n130 B 1.84209f
C306 VTAIL.n131 B 0.369221f
C307 VTAIL.n132 B 0.013574f
C308 VTAIL.n133 B 0.030604f
C309 VTAIL.n134 B 0.01371f
C310 VTAIL.n135 B 0.024096f
C311 VTAIL.n136 B 0.012948f
C312 VTAIL.n137 B 0.030604f
C313 VTAIL.n138 B 0.01371f
C314 VTAIL.n139 B 0.024096f
C315 VTAIL.n140 B 0.012948f
C316 VTAIL.n141 B 0.030604f
C317 VTAIL.n142 B 0.01371f
C318 VTAIL.n143 B 0.024096f
C319 VTAIL.n144 B 0.012948f
C320 VTAIL.n145 B 0.030604f
C321 VTAIL.n146 B 0.01371f
C322 VTAIL.n147 B 0.024096f
C323 VTAIL.n148 B 0.012948f
C324 VTAIL.n149 B 0.030604f
C325 VTAIL.n150 B 0.01371f
C326 VTAIL.n151 B 0.134321f
C327 VTAIL.t8 B 0.05015f
C328 VTAIL.n152 B 0.022953f
C329 VTAIL.n153 B 0.018079f
C330 VTAIL.n154 B 0.012948f
C331 VTAIL.n155 B 1.15026f
C332 VTAIL.n156 B 0.024096f
C333 VTAIL.n157 B 0.012948f
C334 VTAIL.n158 B 0.01371f
C335 VTAIL.n159 B 0.030604f
C336 VTAIL.n160 B 0.030604f
C337 VTAIL.n161 B 0.01371f
C338 VTAIL.n162 B 0.012948f
C339 VTAIL.n163 B 0.024096f
C340 VTAIL.n164 B 0.024096f
C341 VTAIL.n165 B 0.012948f
C342 VTAIL.n166 B 0.01371f
C343 VTAIL.n167 B 0.030604f
C344 VTAIL.n168 B 0.030604f
C345 VTAIL.n169 B 0.01371f
C346 VTAIL.n170 B 0.012948f
C347 VTAIL.n171 B 0.024096f
C348 VTAIL.n172 B 0.024096f
C349 VTAIL.n173 B 0.012948f
C350 VTAIL.n174 B 0.01371f
C351 VTAIL.n175 B 0.030604f
C352 VTAIL.n176 B 0.030604f
C353 VTAIL.n177 B 0.01371f
C354 VTAIL.n178 B 0.012948f
C355 VTAIL.n179 B 0.024096f
C356 VTAIL.n180 B 0.024096f
C357 VTAIL.n181 B 0.012948f
C358 VTAIL.n182 B 0.01371f
C359 VTAIL.n183 B 0.030604f
C360 VTAIL.n184 B 0.030604f
C361 VTAIL.n185 B 0.01371f
C362 VTAIL.n186 B 0.012948f
C363 VTAIL.n187 B 0.024096f
C364 VTAIL.n188 B 0.061621f
C365 VTAIL.n189 B 0.012948f
C366 VTAIL.n190 B 0.01371f
C367 VTAIL.n191 B 0.059928f
C368 VTAIL.n192 B 0.050876f
C369 VTAIL.n193 B 1.25162f
C370 VTAIL.n194 B 0.013574f
C371 VTAIL.n195 B 0.030604f
C372 VTAIL.n196 B 0.01371f
C373 VTAIL.n197 B 0.024096f
C374 VTAIL.n198 B 0.012948f
C375 VTAIL.n199 B 0.030604f
C376 VTAIL.n200 B 0.01371f
C377 VTAIL.n201 B 0.024096f
C378 VTAIL.n202 B 0.012948f
C379 VTAIL.n203 B 0.030604f
C380 VTAIL.n204 B 0.01371f
C381 VTAIL.n205 B 0.024096f
C382 VTAIL.n206 B 0.012948f
C383 VTAIL.n207 B 0.030604f
C384 VTAIL.n208 B 0.01371f
C385 VTAIL.n209 B 0.024096f
C386 VTAIL.n210 B 0.012948f
C387 VTAIL.n211 B 0.030604f
C388 VTAIL.n212 B 0.01371f
C389 VTAIL.n213 B 0.134321f
C390 VTAIL.t0 B 0.05015f
C391 VTAIL.n214 B 0.022953f
C392 VTAIL.n215 B 0.018079f
C393 VTAIL.n216 B 0.012948f
C394 VTAIL.n217 B 1.15026f
C395 VTAIL.n218 B 0.024096f
C396 VTAIL.n219 B 0.012948f
C397 VTAIL.n220 B 0.01371f
C398 VTAIL.n221 B 0.030604f
C399 VTAIL.n222 B 0.030604f
C400 VTAIL.n223 B 0.01371f
C401 VTAIL.n224 B 0.012948f
C402 VTAIL.n225 B 0.024096f
C403 VTAIL.n226 B 0.024096f
C404 VTAIL.n227 B 0.012948f
C405 VTAIL.n228 B 0.01371f
C406 VTAIL.n229 B 0.030604f
C407 VTAIL.n230 B 0.030604f
C408 VTAIL.n231 B 0.01371f
C409 VTAIL.n232 B 0.012948f
C410 VTAIL.n233 B 0.024096f
C411 VTAIL.n234 B 0.024096f
C412 VTAIL.n235 B 0.012948f
C413 VTAIL.n236 B 0.01371f
C414 VTAIL.n237 B 0.030604f
C415 VTAIL.n238 B 0.030604f
C416 VTAIL.n239 B 0.01371f
C417 VTAIL.n240 B 0.012948f
C418 VTAIL.n241 B 0.024096f
C419 VTAIL.n242 B 0.024096f
C420 VTAIL.n243 B 0.012948f
C421 VTAIL.n244 B 0.01371f
C422 VTAIL.n245 B 0.030604f
C423 VTAIL.n246 B 0.030604f
C424 VTAIL.n247 B 0.01371f
C425 VTAIL.n248 B 0.012948f
C426 VTAIL.n249 B 0.024096f
C427 VTAIL.n250 B 0.061621f
C428 VTAIL.n251 B 0.012948f
C429 VTAIL.n252 B 0.01371f
C430 VTAIL.n253 B 0.059928f
C431 VTAIL.n254 B 0.050876f
C432 VTAIL.n255 B 1.2282f
C433 VDD1.n0 B 0.012987f
C434 VDD1.n1 B 0.02928f
C435 VDD1.n2 B 0.013116f
C436 VDD1.n3 B 0.023053f
C437 VDD1.n4 B 0.012388f
C438 VDD1.n5 B 0.02928f
C439 VDD1.n6 B 0.013116f
C440 VDD1.n7 B 0.023053f
C441 VDD1.n8 B 0.012388f
C442 VDD1.n9 B 0.02928f
C443 VDD1.n10 B 0.013116f
C444 VDD1.n11 B 0.023053f
C445 VDD1.n12 B 0.012388f
C446 VDD1.n13 B 0.02928f
C447 VDD1.n14 B 0.013116f
C448 VDD1.n15 B 0.023053f
C449 VDD1.n16 B 0.012388f
C450 VDD1.n17 B 0.02928f
C451 VDD1.n18 B 0.013116f
C452 VDD1.n19 B 0.128509f
C453 VDD1.t5 B 0.04798f
C454 VDD1.n20 B 0.02196f
C455 VDD1.n21 B 0.017296f
C456 VDD1.n22 B 0.012388f
C457 VDD1.n23 B 1.10049f
C458 VDD1.n24 B 0.023053f
C459 VDD1.n25 B 0.012388f
C460 VDD1.n26 B 0.013116f
C461 VDD1.n27 B 0.02928f
C462 VDD1.n28 B 0.02928f
C463 VDD1.n29 B 0.013116f
C464 VDD1.n30 B 0.012388f
C465 VDD1.n31 B 0.023053f
C466 VDD1.n32 B 0.023053f
C467 VDD1.n33 B 0.012388f
C468 VDD1.n34 B 0.013116f
C469 VDD1.n35 B 0.02928f
C470 VDD1.n36 B 0.02928f
C471 VDD1.n37 B 0.013116f
C472 VDD1.n38 B 0.012388f
C473 VDD1.n39 B 0.023053f
C474 VDD1.n40 B 0.023053f
C475 VDD1.n41 B 0.012388f
C476 VDD1.n42 B 0.013116f
C477 VDD1.n43 B 0.02928f
C478 VDD1.n44 B 0.02928f
C479 VDD1.n45 B 0.013116f
C480 VDD1.n46 B 0.012388f
C481 VDD1.n47 B 0.023053f
C482 VDD1.n48 B 0.023053f
C483 VDD1.n49 B 0.012388f
C484 VDD1.n50 B 0.013116f
C485 VDD1.n51 B 0.02928f
C486 VDD1.n52 B 0.02928f
C487 VDD1.n53 B 0.013116f
C488 VDD1.n54 B 0.012388f
C489 VDD1.n55 B 0.023053f
C490 VDD1.n56 B 0.058954f
C491 VDD1.n57 B 0.012388f
C492 VDD1.n58 B 0.013116f
C493 VDD1.n59 B 0.057335f
C494 VDD1.n60 B 0.066182f
C495 VDD1.n61 B 0.012987f
C496 VDD1.n62 B 0.02928f
C497 VDD1.n63 B 0.013116f
C498 VDD1.n64 B 0.023053f
C499 VDD1.n65 B 0.012388f
C500 VDD1.n66 B 0.02928f
C501 VDD1.n67 B 0.013116f
C502 VDD1.n68 B 0.023053f
C503 VDD1.n69 B 0.012388f
C504 VDD1.n70 B 0.02928f
C505 VDD1.n71 B 0.013116f
C506 VDD1.n72 B 0.023053f
C507 VDD1.n73 B 0.012388f
C508 VDD1.n74 B 0.02928f
C509 VDD1.n75 B 0.013116f
C510 VDD1.n76 B 0.023053f
C511 VDD1.n77 B 0.012388f
C512 VDD1.n78 B 0.02928f
C513 VDD1.n79 B 0.013116f
C514 VDD1.n80 B 0.128509f
C515 VDD1.t4 B 0.04798f
C516 VDD1.n81 B 0.02196f
C517 VDD1.n82 B 0.017296f
C518 VDD1.n83 B 0.012388f
C519 VDD1.n84 B 1.10049f
C520 VDD1.n85 B 0.023053f
C521 VDD1.n86 B 0.012388f
C522 VDD1.n87 B 0.013116f
C523 VDD1.n88 B 0.02928f
C524 VDD1.n89 B 0.02928f
C525 VDD1.n90 B 0.013116f
C526 VDD1.n91 B 0.012388f
C527 VDD1.n92 B 0.023053f
C528 VDD1.n93 B 0.023053f
C529 VDD1.n94 B 0.012388f
C530 VDD1.n95 B 0.013116f
C531 VDD1.n96 B 0.02928f
C532 VDD1.n97 B 0.02928f
C533 VDD1.n98 B 0.013116f
C534 VDD1.n99 B 0.012388f
C535 VDD1.n100 B 0.023053f
C536 VDD1.n101 B 0.023053f
C537 VDD1.n102 B 0.012388f
C538 VDD1.n103 B 0.013116f
C539 VDD1.n104 B 0.02928f
C540 VDD1.n105 B 0.02928f
C541 VDD1.n106 B 0.013116f
C542 VDD1.n107 B 0.012388f
C543 VDD1.n108 B 0.023053f
C544 VDD1.n109 B 0.023053f
C545 VDD1.n110 B 0.012388f
C546 VDD1.n111 B 0.013116f
C547 VDD1.n112 B 0.02928f
C548 VDD1.n113 B 0.02928f
C549 VDD1.n114 B 0.013116f
C550 VDD1.n115 B 0.012388f
C551 VDD1.n116 B 0.023053f
C552 VDD1.n117 B 0.058954f
C553 VDD1.n118 B 0.012388f
C554 VDD1.n119 B 0.013116f
C555 VDD1.n120 B 0.057335f
C556 VDD1.n121 B 0.065853f
C557 VDD1.t2 B 0.204396f
C558 VDD1.t0 B 0.204396f
C559 VDD1.n122 B 1.82405f
C560 VDD1.n123 B 1.76975f
C561 VDD1.t1 B 0.204396f
C562 VDD1.t3 B 0.204396f
C563 VDD1.n124 B 1.82325f
C564 VDD1.n125 B 2.03846f
C565 VP.n0 B 0.044509f
C566 VP.n1 B 0.0101f
C567 VP.n2 B 0.192438f
C568 VP.t3 B 1.14125f
C569 VP.t4 B 1.14125f
C570 VP.t5 B 1.16749f
C571 VP.n3 B 0.437084f
C572 VP.n4 B 0.461732f
C573 VP.n5 B 0.0101f
C574 VP.n6 B 0.457403f
C575 VP.n7 B 1.77185f
C576 VP.t1 B 1.14125f
C577 VP.n8 B 0.457403f
C578 VP.n9 B 1.81066f
C579 VP.n10 B 0.044509f
C580 VP.n11 B 0.044509f
C581 VP.t0 B 1.14125f
C582 VP.n12 B 0.45658f
C583 VP.n13 B 0.0101f
C584 VP.t2 B 1.14125f
C585 VP.n14 B 0.457403f
C586 VP.n15 B 0.034493f
.ends

