* NGSPICE file created from diff_pair_sample_0307.ext - technology: sky130A

.subckt diff_pair_sample_0307 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0558 pd=18.85 as=7.2228 ps=37.82 w=18.52 l=1.39
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=0 ps=0 w=18.52 l=1.39
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=0 ps=0 w=18.52 l=1.39
X3 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0558 pd=18.85 as=7.2228 ps=37.82 w=18.52 l=1.39
X4 VTAIL.t7 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=3.0558 ps=18.85 w=18.52 l=1.39
X5 VDD1.t2 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0558 pd=18.85 as=7.2228 ps=37.82 w=18.52 l=1.39
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=0 ps=0 w=18.52 l=1.39
X7 VDD2.t1 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0558 pd=18.85 as=7.2228 ps=37.82 w=18.52 l=1.39
X8 VTAIL.t4 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=3.0558 ps=18.85 w=18.52 l=1.39
X9 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=3.0558 ps=18.85 w=18.52 l=1.39
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=0 ps=0 w=18.52 l=1.39
X11 VTAIL.t3 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=7.2228 pd=37.82 as=3.0558 ps=18.85 w=18.52 l=1.39
R0 VN.n0 VN.t3 359.877
R1 VN.n1 VN.t2 359.877
R2 VN.n0 VN.t0 359.642
R3 VN.n1 VN.t1 359.642
R4 VN VN.n1 65.4262
R5 VN VN.n0 17.5133
R6 VTAIL.n5 VTAIL.t2 43.4728
R7 VTAIL.n4 VTAIL.t5 43.4728
R8 VTAIL.n3 VTAIL.t7 43.4728
R9 VTAIL.n7 VTAIL.t6 43.4727
R10 VTAIL.n0 VTAIL.t4 43.4727
R11 VTAIL.n1 VTAIL.t0 43.4727
R12 VTAIL.n2 VTAIL.t3 43.4727
R13 VTAIL.n6 VTAIL.t1 43.4727
R14 VTAIL.n7 VTAIL.n6 29.8152
R15 VTAIL.n3 VTAIL.n2 29.8152
R16 VTAIL.n4 VTAIL.n3 1.48326
R17 VTAIL.n6 VTAIL.n5 1.48326
R18 VTAIL.n2 VTAIL.n1 1.48326
R19 VTAIL VTAIL.n0 0.800069
R20 VTAIL VTAIL.n7 0.68369
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 103.21
R24 VDD2.n2 VDD2.n1 59.0824
R25 VDD2.n1 VDD2.t2 1.06961
R26 VDD2.n1 VDD2.t1 1.06961
R27 VDD2.n0 VDD2.t0 1.06961
R28 VDD2.n0 VDD2.t3 1.06961
R29 VDD2 VDD2.n2 0.0586897
R30 B.n853 B.n852 585
R31 B.n854 B.n853 585
R32 B.n373 B.n111 585
R33 B.n372 B.n371 585
R34 B.n370 B.n369 585
R35 B.n368 B.n367 585
R36 B.n366 B.n365 585
R37 B.n364 B.n363 585
R38 B.n362 B.n361 585
R39 B.n360 B.n359 585
R40 B.n358 B.n357 585
R41 B.n356 B.n355 585
R42 B.n354 B.n353 585
R43 B.n352 B.n351 585
R44 B.n350 B.n349 585
R45 B.n348 B.n347 585
R46 B.n346 B.n345 585
R47 B.n344 B.n343 585
R48 B.n342 B.n341 585
R49 B.n340 B.n339 585
R50 B.n338 B.n337 585
R51 B.n336 B.n335 585
R52 B.n334 B.n333 585
R53 B.n332 B.n331 585
R54 B.n330 B.n329 585
R55 B.n328 B.n327 585
R56 B.n326 B.n325 585
R57 B.n324 B.n323 585
R58 B.n322 B.n321 585
R59 B.n320 B.n319 585
R60 B.n318 B.n317 585
R61 B.n316 B.n315 585
R62 B.n314 B.n313 585
R63 B.n312 B.n311 585
R64 B.n310 B.n309 585
R65 B.n308 B.n307 585
R66 B.n306 B.n305 585
R67 B.n304 B.n303 585
R68 B.n302 B.n301 585
R69 B.n300 B.n299 585
R70 B.n298 B.n297 585
R71 B.n296 B.n295 585
R72 B.n294 B.n293 585
R73 B.n292 B.n291 585
R74 B.n290 B.n289 585
R75 B.n288 B.n287 585
R76 B.n286 B.n285 585
R77 B.n284 B.n283 585
R78 B.n282 B.n281 585
R79 B.n280 B.n279 585
R80 B.n278 B.n277 585
R81 B.n276 B.n275 585
R82 B.n274 B.n273 585
R83 B.n272 B.n271 585
R84 B.n270 B.n269 585
R85 B.n268 B.n267 585
R86 B.n266 B.n265 585
R87 B.n264 B.n263 585
R88 B.n262 B.n261 585
R89 B.n260 B.n259 585
R90 B.n258 B.n257 585
R91 B.n256 B.n255 585
R92 B.n254 B.n253 585
R93 B.n252 B.n251 585
R94 B.n250 B.n249 585
R95 B.n248 B.n247 585
R96 B.n246 B.n245 585
R97 B.n244 B.n243 585
R98 B.n242 B.n241 585
R99 B.n240 B.n239 585
R100 B.n238 B.n237 585
R101 B.n235 B.n234 585
R102 B.n233 B.n232 585
R103 B.n231 B.n230 585
R104 B.n229 B.n228 585
R105 B.n227 B.n226 585
R106 B.n225 B.n224 585
R107 B.n223 B.n222 585
R108 B.n221 B.n220 585
R109 B.n219 B.n218 585
R110 B.n217 B.n216 585
R111 B.n215 B.n214 585
R112 B.n213 B.n212 585
R113 B.n211 B.n210 585
R114 B.n209 B.n208 585
R115 B.n207 B.n206 585
R116 B.n205 B.n204 585
R117 B.n203 B.n202 585
R118 B.n201 B.n200 585
R119 B.n199 B.n198 585
R120 B.n197 B.n196 585
R121 B.n195 B.n194 585
R122 B.n193 B.n192 585
R123 B.n191 B.n190 585
R124 B.n189 B.n188 585
R125 B.n187 B.n186 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n180 585
R129 B.n179 B.n178 585
R130 B.n177 B.n176 585
R131 B.n175 B.n174 585
R132 B.n173 B.n172 585
R133 B.n171 B.n170 585
R134 B.n169 B.n168 585
R135 B.n167 B.n166 585
R136 B.n165 B.n164 585
R137 B.n163 B.n162 585
R138 B.n161 B.n160 585
R139 B.n159 B.n158 585
R140 B.n157 B.n156 585
R141 B.n155 B.n154 585
R142 B.n153 B.n152 585
R143 B.n151 B.n150 585
R144 B.n149 B.n148 585
R145 B.n147 B.n146 585
R146 B.n145 B.n144 585
R147 B.n143 B.n142 585
R148 B.n141 B.n140 585
R149 B.n139 B.n138 585
R150 B.n137 B.n136 585
R151 B.n135 B.n134 585
R152 B.n133 B.n132 585
R153 B.n131 B.n130 585
R154 B.n129 B.n128 585
R155 B.n127 B.n126 585
R156 B.n125 B.n124 585
R157 B.n123 B.n122 585
R158 B.n121 B.n120 585
R159 B.n119 B.n118 585
R160 B.n46 B.n45 585
R161 B.n857 B.n856 585
R162 B.n851 B.n112 585
R163 B.n112 B.n43 585
R164 B.n850 B.n42 585
R165 B.n861 B.n42 585
R166 B.n849 B.n41 585
R167 B.n862 B.n41 585
R168 B.n848 B.n40 585
R169 B.n863 B.n40 585
R170 B.n847 B.n846 585
R171 B.n846 B.n36 585
R172 B.n845 B.n35 585
R173 B.n869 B.n35 585
R174 B.n844 B.n34 585
R175 B.n870 B.n34 585
R176 B.n843 B.n33 585
R177 B.n871 B.n33 585
R178 B.n842 B.n841 585
R179 B.n841 B.n29 585
R180 B.n840 B.n28 585
R181 B.n877 B.n28 585
R182 B.n839 B.n27 585
R183 B.n878 B.n27 585
R184 B.n838 B.n26 585
R185 B.n879 B.n26 585
R186 B.n837 B.n836 585
R187 B.n836 B.n22 585
R188 B.n835 B.n21 585
R189 B.n885 B.n21 585
R190 B.n834 B.n20 585
R191 B.n886 B.n20 585
R192 B.n833 B.n19 585
R193 B.n887 B.n19 585
R194 B.n832 B.n831 585
R195 B.n831 B.n15 585
R196 B.n830 B.n14 585
R197 B.n893 B.n14 585
R198 B.n829 B.n13 585
R199 B.n894 B.n13 585
R200 B.n828 B.n12 585
R201 B.n895 B.n12 585
R202 B.n827 B.n826 585
R203 B.n826 B.n825 585
R204 B.n824 B.n823 585
R205 B.n824 B.n8 585
R206 B.n822 B.n7 585
R207 B.n902 B.n7 585
R208 B.n821 B.n6 585
R209 B.n903 B.n6 585
R210 B.n820 B.n5 585
R211 B.n904 B.n5 585
R212 B.n819 B.n818 585
R213 B.n818 B.n4 585
R214 B.n817 B.n374 585
R215 B.n817 B.n816 585
R216 B.n807 B.n375 585
R217 B.n376 B.n375 585
R218 B.n809 B.n808 585
R219 B.n810 B.n809 585
R220 B.n806 B.n381 585
R221 B.n381 B.n380 585
R222 B.n805 B.n804 585
R223 B.n804 B.n803 585
R224 B.n383 B.n382 585
R225 B.n384 B.n383 585
R226 B.n796 B.n795 585
R227 B.n797 B.n796 585
R228 B.n794 B.n388 585
R229 B.n392 B.n388 585
R230 B.n793 B.n792 585
R231 B.n792 B.n791 585
R232 B.n390 B.n389 585
R233 B.n391 B.n390 585
R234 B.n784 B.n783 585
R235 B.n785 B.n784 585
R236 B.n782 B.n397 585
R237 B.n397 B.n396 585
R238 B.n781 B.n780 585
R239 B.n780 B.n779 585
R240 B.n399 B.n398 585
R241 B.n400 B.n399 585
R242 B.n772 B.n771 585
R243 B.n773 B.n772 585
R244 B.n770 B.n404 585
R245 B.n408 B.n404 585
R246 B.n769 B.n768 585
R247 B.n768 B.n767 585
R248 B.n406 B.n405 585
R249 B.n407 B.n406 585
R250 B.n760 B.n759 585
R251 B.n761 B.n760 585
R252 B.n758 B.n413 585
R253 B.n413 B.n412 585
R254 B.n757 B.n756 585
R255 B.n756 B.n755 585
R256 B.n415 B.n414 585
R257 B.n416 B.n415 585
R258 B.n751 B.n750 585
R259 B.n419 B.n418 585
R260 B.n747 B.n746 585
R261 B.n748 B.n747 585
R262 B.n745 B.n484 585
R263 B.n744 B.n743 585
R264 B.n742 B.n741 585
R265 B.n740 B.n739 585
R266 B.n738 B.n737 585
R267 B.n736 B.n735 585
R268 B.n734 B.n733 585
R269 B.n732 B.n731 585
R270 B.n730 B.n729 585
R271 B.n728 B.n727 585
R272 B.n726 B.n725 585
R273 B.n724 B.n723 585
R274 B.n722 B.n721 585
R275 B.n720 B.n719 585
R276 B.n718 B.n717 585
R277 B.n716 B.n715 585
R278 B.n714 B.n713 585
R279 B.n712 B.n711 585
R280 B.n710 B.n709 585
R281 B.n708 B.n707 585
R282 B.n706 B.n705 585
R283 B.n704 B.n703 585
R284 B.n702 B.n701 585
R285 B.n700 B.n699 585
R286 B.n698 B.n697 585
R287 B.n696 B.n695 585
R288 B.n694 B.n693 585
R289 B.n692 B.n691 585
R290 B.n690 B.n689 585
R291 B.n688 B.n687 585
R292 B.n686 B.n685 585
R293 B.n684 B.n683 585
R294 B.n682 B.n681 585
R295 B.n680 B.n679 585
R296 B.n678 B.n677 585
R297 B.n676 B.n675 585
R298 B.n674 B.n673 585
R299 B.n672 B.n671 585
R300 B.n670 B.n669 585
R301 B.n668 B.n667 585
R302 B.n666 B.n665 585
R303 B.n664 B.n663 585
R304 B.n662 B.n661 585
R305 B.n660 B.n659 585
R306 B.n658 B.n657 585
R307 B.n656 B.n655 585
R308 B.n654 B.n653 585
R309 B.n652 B.n651 585
R310 B.n650 B.n649 585
R311 B.n648 B.n647 585
R312 B.n646 B.n645 585
R313 B.n644 B.n643 585
R314 B.n642 B.n641 585
R315 B.n640 B.n639 585
R316 B.n638 B.n637 585
R317 B.n636 B.n635 585
R318 B.n634 B.n633 585
R319 B.n632 B.n631 585
R320 B.n630 B.n629 585
R321 B.n628 B.n627 585
R322 B.n626 B.n625 585
R323 B.n624 B.n623 585
R324 B.n622 B.n621 585
R325 B.n620 B.n619 585
R326 B.n618 B.n617 585
R327 B.n616 B.n615 585
R328 B.n614 B.n613 585
R329 B.n611 B.n610 585
R330 B.n609 B.n608 585
R331 B.n607 B.n606 585
R332 B.n605 B.n604 585
R333 B.n603 B.n602 585
R334 B.n601 B.n600 585
R335 B.n599 B.n598 585
R336 B.n597 B.n596 585
R337 B.n595 B.n594 585
R338 B.n593 B.n592 585
R339 B.n591 B.n590 585
R340 B.n589 B.n588 585
R341 B.n587 B.n586 585
R342 B.n585 B.n584 585
R343 B.n583 B.n582 585
R344 B.n581 B.n580 585
R345 B.n579 B.n578 585
R346 B.n577 B.n576 585
R347 B.n575 B.n574 585
R348 B.n573 B.n572 585
R349 B.n571 B.n570 585
R350 B.n569 B.n568 585
R351 B.n567 B.n566 585
R352 B.n565 B.n564 585
R353 B.n563 B.n562 585
R354 B.n561 B.n560 585
R355 B.n559 B.n558 585
R356 B.n557 B.n556 585
R357 B.n555 B.n554 585
R358 B.n553 B.n552 585
R359 B.n551 B.n550 585
R360 B.n549 B.n548 585
R361 B.n547 B.n546 585
R362 B.n545 B.n544 585
R363 B.n543 B.n542 585
R364 B.n541 B.n540 585
R365 B.n539 B.n538 585
R366 B.n537 B.n536 585
R367 B.n535 B.n534 585
R368 B.n533 B.n532 585
R369 B.n531 B.n530 585
R370 B.n529 B.n528 585
R371 B.n527 B.n526 585
R372 B.n525 B.n524 585
R373 B.n523 B.n522 585
R374 B.n521 B.n520 585
R375 B.n519 B.n518 585
R376 B.n517 B.n516 585
R377 B.n515 B.n514 585
R378 B.n513 B.n512 585
R379 B.n511 B.n510 585
R380 B.n509 B.n508 585
R381 B.n507 B.n506 585
R382 B.n505 B.n504 585
R383 B.n503 B.n502 585
R384 B.n501 B.n500 585
R385 B.n499 B.n498 585
R386 B.n497 B.n496 585
R387 B.n495 B.n494 585
R388 B.n493 B.n492 585
R389 B.n491 B.n490 585
R390 B.n752 B.n417 585
R391 B.n417 B.n416 585
R392 B.n754 B.n753 585
R393 B.n755 B.n754 585
R394 B.n411 B.n410 585
R395 B.n412 B.n411 585
R396 B.n763 B.n762 585
R397 B.n762 B.n761 585
R398 B.n764 B.n409 585
R399 B.n409 B.n407 585
R400 B.n766 B.n765 585
R401 B.n767 B.n766 585
R402 B.n403 B.n402 585
R403 B.n408 B.n403 585
R404 B.n775 B.n774 585
R405 B.n774 B.n773 585
R406 B.n776 B.n401 585
R407 B.n401 B.n400 585
R408 B.n778 B.n777 585
R409 B.n779 B.n778 585
R410 B.n395 B.n394 585
R411 B.n396 B.n395 585
R412 B.n787 B.n786 585
R413 B.n786 B.n785 585
R414 B.n788 B.n393 585
R415 B.n393 B.n391 585
R416 B.n790 B.n789 585
R417 B.n791 B.n790 585
R418 B.n387 B.n386 585
R419 B.n392 B.n387 585
R420 B.n799 B.n798 585
R421 B.n798 B.n797 585
R422 B.n800 B.n385 585
R423 B.n385 B.n384 585
R424 B.n802 B.n801 585
R425 B.n803 B.n802 585
R426 B.n379 B.n378 585
R427 B.n380 B.n379 585
R428 B.n812 B.n811 585
R429 B.n811 B.n810 585
R430 B.n813 B.n377 585
R431 B.n377 B.n376 585
R432 B.n815 B.n814 585
R433 B.n816 B.n815 585
R434 B.n3 B.n0 585
R435 B.n4 B.n3 585
R436 B.n901 B.n1 585
R437 B.n902 B.n901 585
R438 B.n900 B.n899 585
R439 B.n900 B.n8 585
R440 B.n898 B.n9 585
R441 B.n825 B.n9 585
R442 B.n897 B.n896 585
R443 B.n896 B.n895 585
R444 B.n11 B.n10 585
R445 B.n894 B.n11 585
R446 B.n892 B.n891 585
R447 B.n893 B.n892 585
R448 B.n890 B.n16 585
R449 B.n16 B.n15 585
R450 B.n889 B.n888 585
R451 B.n888 B.n887 585
R452 B.n18 B.n17 585
R453 B.n886 B.n18 585
R454 B.n884 B.n883 585
R455 B.n885 B.n884 585
R456 B.n882 B.n23 585
R457 B.n23 B.n22 585
R458 B.n881 B.n880 585
R459 B.n880 B.n879 585
R460 B.n25 B.n24 585
R461 B.n878 B.n25 585
R462 B.n876 B.n875 585
R463 B.n877 B.n876 585
R464 B.n874 B.n30 585
R465 B.n30 B.n29 585
R466 B.n873 B.n872 585
R467 B.n872 B.n871 585
R468 B.n32 B.n31 585
R469 B.n870 B.n32 585
R470 B.n868 B.n867 585
R471 B.n869 B.n868 585
R472 B.n866 B.n37 585
R473 B.n37 B.n36 585
R474 B.n865 B.n864 585
R475 B.n864 B.n863 585
R476 B.n39 B.n38 585
R477 B.n862 B.n39 585
R478 B.n860 B.n859 585
R479 B.n861 B.n860 585
R480 B.n858 B.n44 585
R481 B.n44 B.n43 585
R482 B.n905 B.n904 585
R483 B.n903 B.n2 585
R484 B.n116 B.t15 526.107
R485 B.n113 B.t4 526.107
R486 B.n488 B.t8 526.107
R487 B.n485 B.t12 526.107
R488 B.n856 B.n44 478.086
R489 B.n853 B.n112 478.086
R490 B.n490 B.n415 478.086
R491 B.n750 B.n417 478.086
R492 B.n854 B.n110 256.663
R493 B.n854 B.n109 256.663
R494 B.n854 B.n108 256.663
R495 B.n854 B.n107 256.663
R496 B.n854 B.n106 256.663
R497 B.n854 B.n105 256.663
R498 B.n854 B.n104 256.663
R499 B.n854 B.n103 256.663
R500 B.n854 B.n102 256.663
R501 B.n854 B.n101 256.663
R502 B.n854 B.n100 256.663
R503 B.n854 B.n99 256.663
R504 B.n854 B.n98 256.663
R505 B.n854 B.n97 256.663
R506 B.n854 B.n96 256.663
R507 B.n854 B.n95 256.663
R508 B.n854 B.n94 256.663
R509 B.n854 B.n93 256.663
R510 B.n854 B.n92 256.663
R511 B.n854 B.n91 256.663
R512 B.n854 B.n90 256.663
R513 B.n854 B.n89 256.663
R514 B.n854 B.n88 256.663
R515 B.n854 B.n87 256.663
R516 B.n854 B.n86 256.663
R517 B.n854 B.n85 256.663
R518 B.n854 B.n84 256.663
R519 B.n854 B.n83 256.663
R520 B.n854 B.n82 256.663
R521 B.n854 B.n81 256.663
R522 B.n854 B.n80 256.663
R523 B.n854 B.n79 256.663
R524 B.n854 B.n78 256.663
R525 B.n854 B.n77 256.663
R526 B.n854 B.n76 256.663
R527 B.n854 B.n75 256.663
R528 B.n854 B.n74 256.663
R529 B.n854 B.n73 256.663
R530 B.n854 B.n72 256.663
R531 B.n854 B.n71 256.663
R532 B.n854 B.n70 256.663
R533 B.n854 B.n69 256.663
R534 B.n854 B.n68 256.663
R535 B.n854 B.n67 256.663
R536 B.n854 B.n66 256.663
R537 B.n854 B.n65 256.663
R538 B.n854 B.n64 256.663
R539 B.n854 B.n63 256.663
R540 B.n854 B.n62 256.663
R541 B.n854 B.n61 256.663
R542 B.n854 B.n60 256.663
R543 B.n854 B.n59 256.663
R544 B.n854 B.n58 256.663
R545 B.n854 B.n57 256.663
R546 B.n854 B.n56 256.663
R547 B.n854 B.n55 256.663
R548 B.n854 B.n54 256.663
R549 B.n854 B.n53 256.663
R550 B.n854 B.n52 256.663
R551 B.n854 B.n51 256.663
R552 B.n854 B.n50 256.663
R553 B.n854 B.n49 256.663
R554 B.n854 B.n48 256.663
R555 B.n854 B.n47 256.663
R556 B.n855 B.n854 256.663
R557 B.n749 B.n748 256.663
R558 B.n748 B.n420 256.663
R559 B.n748 B.n421 256.663
R560 B.n748 B.n422 256.663
R561 B.n748 B.n423 256.663
R562 B.n748 B.n424 256.663
R563 B.n748 B.n425 256.663
R564 B.n748 B.n426 256.663
R565 B.n748 B.n427 256.663
R566 B.n748 B.n428 256.663
R567 B.n748 B.n429 256.663
R568 B.n748 B.n430 256.663
R569 B.n748 B.n431 256.663
R570 B.n748 B.n432 256.663
R571 B.n748 B.n433 256.663
R572 B.n748 B.n434 256.663
R573 B.n748 B.n435 256.663
R574 B.n748 B.n436 256.663
R575 B.n748 B.n437 256.663
R576 B.n748 B.n438 256.663
R577 B.n748 B.n439 256.663
R578 B.n748 B.n440 256.663
R579 B.n748 B.n441 256.663
R580 B.n748 B.n442 256.663
R581 B.n748 B.n443 256.663
R582 B.n748 B.n444 256.663
R583 B.n748 B.n445 256.663
R584 B.n748 B.n446 256.663
R585 B.n748 B.n447 256.663
R586 B.n748 B.n448 256.663
R587 B.n748 B.n449 256.663
R588 B.n748 B.n450 256.663
R589 B.n748 B.n451 256.663
R590 B.n748 B.n452 256.663
R591 B.n748 B.n453 256.663
R592 B.n748 B.n454 256.663
R593 B.n748 B.n455 256.663
R594 B.n748 B.n456 256.663
R595 B.n748 B.n457 256.663
R596 B.n748 B.n458 256.663
R597 B.n748 B.n459 256.663
R598 B.n748 B.n460 256.663
R599 B.n748 B.n461 256.663
R600 B.n748 B.n462 256.663
R601 B.n748 B.n463 256.663
R602 B.n748 B.n464 256.663
R603 B.n748 B.n465 256.663
R604 B.n748 B.n466 256.663
R605 B.n748 B.n467 256.663
R606 B.n748 B.n468 256.663
R607 B.n748 B.n469 256.663
R608 B.n748 B.n470 256.663
R609 B.n748 B.n471 256.663
R610 B.n748 B.n472 256.663
R611 B.n748 B.n473 256.663
R612 B.n748 B.n474 256.663
R613 B.n748 B.n475 256.663
R614 B.n748 B.n476 256.663
R615 B.n748 B.n477 256.663
R616 B.n748 B.n478 256.663
R617 B.n748 B.n479 256.663
R618 B.n748 B.n480 256.663
R619 B.n748 B.n481 256.663
R620 B.n748 B.n482 256.663
R621 B.n748 B.n483 256.663
R622 B.n907 B.n906 256.663
R623 B.n118 B.n46 163.367
R624 B.n122 B.n121 163.367
R625 B.n126 B.n125 163.367
R626 B.n130 B.n129 163.367
R627 B.n134 B.n133 163.367
R628 B.n138 B.n137 163.367
R629 B.n142 B.n141 163.367
R630 B.n146 B.n145 163.367
R631 B.n150 B.n149 163.367
R632 B.n154 B.n153 163.367
R633 B.n158 B.n157 163.367
R634 B.n162 B.n161 163.367
R635 B.n166 B.n165 163.367
R636 B.n170 B.n169 163.367
R637 B.n174 B.n173 163.367
R638 B.n178 B.n177 163.367
R639 B.n182 B.n181 163.367
R640 B.n186 B.n185 163.367
R641 B.n190 B.n189 163.367
R642 B.n194 B.n193 163.367
R643 B.n198 B.n197 163.367
R644 B.n202 B.n201 163.367
R645 B.n206 B.n205 163.367
R646 B.n210 B.n209 163.367
R647 B.n214 B.n213 163.367
R648 B.n218 B.n217 163.367
R649 B.n222 B.n221 163.367
R650 B.n226 B.n225 163.367
R651 B.n230 B.n229 163.367
R652 B.n234 B.n233 163.367
R653 B.n239 B.n238 163.367
R654 B.n243 B.n242 163.367
R655 B.n247 B.n246 163.367
R656 B.n251 B.n250 163.367
R657 B.n255 B.n254 163.367
R658 B.n259 B.n258 163.367
R659 B.n263 B.n262 163.367
R660 B.n267 B.n266 163.367
R661 B.n271 B.n270 163.367
R662 B.n275 B.n274 163.367
R663 B.n279 B.n278 163.367
R664 B.n283 B.n282 163.367
R665 B.n287 B.n286 163.367
R666 B.n291 B.n290 163.367
R667 B.n295 B.n294 163.367
R668 B.n299 B.n298 163.367
R669 B.n303 B.n302 163.367
R670 B.n307 B.n306 163.367
R671 B.n311 B.n310 163.367
R672 B.n315 B.n314 163.367
R673 B.n319 B.n318 163.367
R674 B.n323 B.n322 163.367
R675 B.n327 B.n326 163.367
R676 B.n331 B.n330 163.367
R677 B.n335 B.n334 163.367
R678 B.n339 B.n338 163.367
R679 B.n343 B.n342 163.367
R680 B.n347 B.n346 163.367
R681 B.n351 B.n350 163.367
R682 B.n355 B.n354 163.367
R683 B.n359 B.n358 163.367
R684 B.n363 B.n362 163.367
R685 B.n367 B.n366 163.367
R686 B.n371 B.n370 163.367
R687 B.n853 B.n111 163.367
R688 B.n756 B.n415 163.367
R689 B.n756 B.n413 163.367
R690 B.n760 B.n413 163.367
R691 B.n760 B.n406 163.367
R692 B.n768 B.n406 163.367
R693 B.n768 B.n404 163.367
R694 B.n772 B.n404 163.367
R695 B.n772 B.n399 163.367
R696 B.n780 B.n399 163.367
R697 B.n780 B.n397 163.367
R698 B.n784 B.n397 163.367
R699 B.n784 B.n390 163.367
R700 B.n792 B.n390 163.367
R701 B.n792 B.n388 163.367
R702 B.n796 B.n388 163.367
R703 B.n796 B.n383 163.367
R704 B.n804 B.n383 163.367
R705 B.n804 B.n381 163.367
R706 B.n809 B.n381 163.367
R707 B.n809 B.n375 163.367
R708 B.n817 B.n375 163.367
R709 B.n818 B.n817 163.367
R710 B.n818 B.n5 163.367
R711 B.n6 B.n5 163.367
R712 B.n7 B.n6 163.367
R713 B.n824 B.n7 163.367
R714 B.n826 B.n824 163.367
R715 B.n826 B.n12 163.367
R716 B.n13 B.n12 163.367
R717 B.n14 B.n13 163.367
R718 B.n831 B.n14 163.367
R719 B.n831 B.n19 163.367
R720 B.n20 B.n19 163.367
R721 B.n21 B.n20 163.367
R722 B.n836 B.n21 163.367
R723 B.n836 B.n26 163.367
R724 B.n27 B.n26 163.367
R725 B.n28 B.n27 163.367
R726 B.n841 B.n28 163.367
R727 B.n841 B.n33 163.367
R728 B.n34 B.n33 163.367
R729 B.n35 B.n34 163.367
R730 B.n846 B.n35 163.367
R731 B.n846 B.n40 163.367
R732 B.n41 B.n40 163.367
R733 B.n42 B.n41 163.367
R734 B.n112 B.n42 163.367
R735 B.n747 B.n419 163.367
R736 B.n747 B.n484 163.367
R737 B.n743 B.n742 163.367
R738 B.n739 B.n738 163.367
R739 B.n735 B.n734 163.367
R740 B.n731 B.n730 163.367
R741 B.n727 B.n726 163.367
R742 B.n723 B.n722 163.367
R743 B.n719 B.n718 163.367
R744 B.n715 B.n714 163.367
R745 B.n711 B.n710 163.367
R746 B.n707 B.n706 163.367
R747 B.n703 B.n702 163.367
R748 B.n699 B.n698 163.367
R749 B.n695 B.n694 163.367
R750 B.n691 B.n690 163.367
R751 B.n687 B.n686 163.367
R752 B.n683 B.n682 163.367
R753 B.n679 B.n678 163.367
R754 B.n675 B.n674 163.367
R755 B.n671 B.n670 163.367
R756 B.n667 B.n666 163.367
R757 B.n663 B.n662 163.367
R758 B.n659 B.n658 163.367
R759 B.n655 B.n654 163.367
R760 B.n651 B.n650 163.367
R761 B.n647 B.n646 163.367
R762 B.n643 B.n642 163.367
R763 B.n639 B.n638 163.367
R764 B.n635 B.n634 163.367
R765 B.n631 B.n630 163.367
R766 B.n627 B.n626 163.367
R767 B.n623 B.n622 163.367
R768 B.n619 B.n618 163.367
R769 B.n615 B.n614 163.367
R770 B.n610 B.n609 163.367
R771 B.n606 B.n605 163.367
R772 B.n602 B.n601 163.367
R773 B.n598 B.n597 163.367
R774 B.n594 B.n593 163.367
R775 B.n590 B.n589 163.367
R776 B.n586 B.n585 163.367
R777 B.n582 B.n581 163.367
R778 B.n578 B.n577 163.367
R779 B.n574 B.n573 163.367
R780 B.n570 B.n569 163.367
R781 B.n566 B.n565 163.367
R782 B.n562 B.n561 163.367
R783 B.n558 B.n557 163.367
R784 B.n554 B.n553 163.367
R785 B.n550 B.n549 163.367
R786 B.n546 B.n545 163.367
R787 B.n542 B.n541 163.367
R788 B.n538 B.n537 163.367
R789 B.n534 B.n533 163.367
R790 B.n530 B.n529 163.367
R791 B.n526 B.n525 163.367
R792 B.n522 B.n521 163.367
R793 B.n518 B.n517 163.367
R794 B.n514 B.n513 163.367
R795 B.n510 B.n509 163.367
R796 B.n506 B.n505 163.367
R797 B.n502 B.n501 163.367
R798 B.n498 B.n497 163.367
R799 B.n494 B.n493 163.367
R800 B.n754 B.n417 163.367
R801 B.n754 B.n411 163.367
R802 B.n762 B.n411 163.367
R803 B.n762 B.n409 163.367
R804 B.n766 B.n409 163.367
R805 B.n766 B.n403 163.367
R806 B.n774 B.n403 163.367
R807 B.n774 B.n401 163.367
R808 B.n778 B.n401 163.367
R809 B.n778 B.n395 163.367
R810 B.n786 B.n395 163.367
R811 B.n786 B.n393 163.367
R812 B.n790 B.n393 163.367
R813 B.n790 B.n387 163.367
R814 B.n798 B.n387 163.367
R815 B.n798 B.n385 163.367
R816 B.n802 B.n385 163.367
R817 B.n802 B.n379 163.367
R818 B.n811 B.n379 163.367
R819 B.n811 B.n377 163.367
R820 B.n815 B.n377 163.367
R821 B.n815 B.n3 163.367
R822 B.n905 B.n3 163.367
R823 B.n901 B.n2 163.367
R824 B.n901 B.n900 163.367
R825 B.n900 B.n9 163.367
R826 B.n896 B.n9 163.367
R827 B.n896 B.n11 163.367
R828 B.n892 B.n11 163.367
R829 B.n892 B.n16 163.367
R830 B.n888 B.n16 163.367
R831 B.n888 B.n18 163.367
R832 B.n884 B.n18 163.367
R833 B.n884 B.n23 163.367
R834 B.n880 B.n23 163.367
R835 B.n880 B.n25 163.367
R836 B.n876 B.n25 163.367
R837 B.n876 B.n30 163.367
R838 B.n872 B.n30 163.367
R839 B.n872 B.n32 163.367
R840 B.n868 B.n32 163.367
R841 B.n868 B.n37 163.367
R842 B.n864 B.n37 163.367
R843 B.n864 B.n39 163.367
R844 B.n860 B.n39 163.367
R845 B.n860 B.n44 163.367
R846 B.n113 B.t6 103.68
R847 B.n488 B.t11 103.68
R848 B.n116 B.t16 103.654
R849 B.n485 B.t14 103.654
R850 B.n856 B.n855 71.676
R851 B.n118 B.n47 71.676
R852 B.n122 B.n48 71.676
R853 B.n126 B.n49 71.676
R854 B.n130 B.n50 71.676
R855 B.n134 B.n51 71.676
R856 B.n138 B.n52 71.676
R857 B.n142 B.n53 71.676
R858 B.n146 B.n54 71.676
R859 B.n150 B.n55 71.676
R860 B.n154 B.n56 71.676
R861 B.n158 B.n57 71.676
R862 B.n162 B.n58 71.676
R863 B.n166 B.n59 71.676
R864 B.n170 B.n60 71.676
R865 B.n174 B.n61 71.676
R866 B.n178 B.n62 71.676
R867 B.n182 B.n63 71.676
R868 B.n186 B.n64 71.676
R869 B.n190 B.n65 71.676
R870 B.n194 B.n66 71.676
R871 B.n198 B.n67 71.676
R872 B.n202 B.n68 71.676
R873 B.n206 B.n69 71.676
R874 B.n210 B.n70 71.676
R875 B.n214 B.n71 71.676
R876 B.n218 B.n72 71.676
R877 B.n222 B.n73 71.676
R878 B.n226 B.n74 71.676
R879 B.n230 B.n75 71.676
R880 B.n234 B.n76 71.676
R881 B.n239 B.n77 71.676
R882 B.n243 B.n78 71.676
R883 B.n247 B.n79 71.676
R884 B.n251 B.n80 71.676
R885 B.n255 B.n81 71.676
R886 B.n259 B.n82 71.676
R887 B.n263 B.n83 71.676
R888 B.n267 B.n84 71.676
R889 B.n271 B.n85 71.676
R890 B.n275 B.n86 71.676
R891 B.n279 B.n87 71.676
R892 B.n283 B.n88 71.676
R893 B.n287 B.n89 71.676
R894 B.n291 B.n90 71.676
R895 B.n295 B.n91 71.676
R896 B.n299 B.n92 71.676
R897 B.n303 B.n93 71.676
R898 B.n307 B.n94 71.676
R899 B.n311 B.n95 71.676
R900 B.n315 B.n96 71.676
R901 B.n319 B.n97 71.676
R902 B.n323 B.n98 71.676
R903 B.n327 B.n99 71.676
R904 B.n331 B.n100 71.676
R905 B.n335 B.n101 71.676
R906 B.n339 B.n102 71.676
R907 B.n343 B.n103 71.676
R908 B.n347 B.n104 71.676
R909 B.n351 B.n105 71.676
R910 B.n355 B.n106 71.676
R911 B.n359 B.n107 71.676
R912 B.n363 B.n108 71.676
R913 B.n367 B.n109 71.676
R914 B.n371 B.n110 71.676
R915 B.n111 B.n110 71.676
R916 B.n370 B.n109 71.676
R917 B.n366 B.n108 71.676
R918 B.n362 B.n107 71.676
R919 B.n358 B.n106 71.676
R920 B.n354 B.n105 71.676
R921 B.n350 B.n104 71.676
R922 B.n346 B.n103 71.676
R923 B.n342 B.n102 71.676
R924 B.n338 B.n101 71.676
R925 B.n334 B.n100 71.676
R926 B.n330 B.n99 71.676
R927 B.n326 B.n98 71.676
R928 B.n322 B.n97 71.676
R929 B.n318 B.n96 71.676
R930 B.n314 B.n95 71.676
R931 B.n310 B.n94 71.676
R932 B.n306 B.n93 71.676
R933 B.n302 B.n92 71.676
R934 B.n298 B.n91 71.676
R935 B.n294 B.n90 71.676
R936 B.n290 B.n89 71.676
R937 B.n286 B.n88 71.676
R938 B.n282 B.n87 71.676
R939 B.n278 B.n86 71.676
R940 B.n274 B.n85 71.676
R941 B.n270 B.n84 71.676
R942 B.n266 B.n83 71.676
R943 B.n262 B.n82 71.676
R944 B.n258 B.n81 71.676
R945 B.n254 B.n80 71.676
R946 B.n250 B.n79 71.676
R947 B.n246 B.n78 71.676
R948 B.n242 B.n77 71.676
R949 B.n238 B.n76 71.676
R950 B.n233 B.n75 71.676
R951 B.n229 B.n74 71.676
R952 B.n225 B.n73 71.676
R953 B.n221 B.n72 71.676
R954 B.n217 B.n71 71.676
R955 B.n213 B.n70 71.676
R956 B.n209 B.n69 71.676
R957 B.n205 B.n68 71.676
R958 B.n201 B.n67 71.676
R959 B.n197 B.n66 71.676
R960 B.n193 B.n65 71.676
R961 B.n189 B.n64 71.676
R962 B.n185 B.n63 71.676
R963 B.n181 B.n62 71.676
R964 B.n177 B.n61 71.676
R965 B.n173 B.n60 71.676
R966 B.n169 B.n59 71.676
R967 B.n165 B.n58 71.676
R968 B.n161 B.n57 71.676
R969 B.n157 B.n56 71.676
R970 B.n153 B.n55 71.676
R971 B.n149 B.n54 71.676
R972 B.n145 B.n53 71.676
R973 B.n141 B.n52 71.676
R974 B.n137 B.n51 71.676
R975 B.n133 B.n50 71.676
R976 B.n129 B.n49 71.676
R977 B.n125 B.n48 71.676
R978 B.n121 B.n47 71.676
R979 B.n855 B.n46 71.676
R980 B.n750 B.n749 71.676
R981 B.n484 B.n420 71.676
R982 B.n742 B.n421 71.676
R983 B.n738 B.n422 71.676
R984 B.n734 B.n423 71.676
R985 B.n730 B.n424 71.676
R986 B.n726 B.n425 71.676
R987 B.n722 B.n426 71.676
R988 B.n718 B.n427 71.676
R989 B.n714 B.n428 71.676
R990 B.n710 B.n429 71.676
R991 B.n706 B.n430 71.676
R992 B.n702 B.n431 71.676
R993 B.n698 B.n432 71.676
R994 B.n694 B.n433 71.676
R995 B.n690 B.n434 71.676
R996 B.n686 B.n435 71.676
R997 B.n682 B.n436 71.676
R998 B.n678 B.n437 71.676
R999 B.n674 B.n438 71.676
R1000 B.n670 B.n439 71.676
R1001 B.n666 B.n440 71.676
R1002 B.n662 B.n441 71.676
R1003 B.n658 B.n442 71.676
R1004 B.n654 B.n443 71.676
R1005 B.n650 B.n444 71.676
R1006 B.n646 B.n445 71.676
R1007 B.n642 B.n446 71.676
R1008 B.n638 B.n447 71.676
R1009 B.n634 B.n448 71.676
R1010 B.n630 B.n449 71.676
R1011 B.n626 B.n450 71.676
R1012 B.n622 B.n451 71.676
R1013 B.n618 B.n452 71.676
R1014 B.n614 B.n453 71.676
R1015 B.n609 B.n454 71.676
R1016 B.n605 B.n455 71.676
R1017 B.n601 B.n456 71.676
R1018 B.n597 B.n457 71.676
R1019 B.n593 B.n458 71.676
R1020 B.n589 B.n459 71.676
R1021 B.n585 B.n460 71.676
R1022 B.n581 B.n461 71.676
R1023 B.n577 B.n462 71.676
R1024 B.n573 B.n463 71.676
R1025 B.n569 B.n464 71.676
R1026 B.n565 B.n465 71.676
R1027 B.n561 B.n466 71.676
R1028 B.n557 B.n467 71.676
R1029 B.n553 B.n468 71.676
R1030 B.n549 B.n469 71.676
R1031 B.n545 B.n470 71.676
R1032 B.n541 B.n471 71.676
R1033 B.n537 B.n472 71.676
R1034 B.n533 B.n473 71.676
R1035 B.n529 B.n474 71.676
R1036 B.n525 B.n475 71.676
R1037 B.n521 B.n476 71.676
R1038 B.n517 B.n477 71.676
R1039 B.n513 B.n478 71.676
R1040 B.n509 B.n479 71.676
R1041 B.n505 B.n480 71.676
R1042 B.n501 B.n481 71.676
R1043 B.n497 B.n482 71.676
R1044 B.n493 B.n483 71.676
R1045 B.n749 B.n419 71.676
R1046 B.n743 B.n420 71.676
R1047 B.n739 B.n421 71.676
R1048 B.n735 B.n422 71.676
R1049 B.n731 B.n423 71.676
R1050 B.n727 B.n424 71.676
R1051 B.n723 B.n425 71.676
R1052 B.n719 B.n426 71.676
R1053 B.n715 B.n427 71.676
R1054 B.n711 B.n428 71.676
R1055 B.n707 B.n429 71.676
R1056 B.n703 B.n430 71.676
R1057 B.n699 B.n431 71.676
R1058 B.n695 B.n432 71.676
R1059 B.n691 B.n433 71.676
R1060 B.n687 B.n434 71.676
R1061 B.n683 B.n435 71.676
R1062 B.n679 B.n436 71.676
R1063 B.n675 B.n437 71.676
R1064 B.n671 B.n438 71.676
R1065 B.n667 B.n439 71.676
R1066 B.n663 B.n440 71.676
R1067 B.n659 B.n441 71.676
R1068 B.n655 B.n442 71.676
R1069 B.n651 B.n443 71.676
R1070 B.n647 B.n444 71.676
R1071 B.n643 B.n445 71.676
R1072 B.n639 B.n446 71.676
R1073 B.n635 B.n447 71.676
R1074 B.n631 B.n448 71.676
R1075 B.n627 B.n449 71.676
R1076 B.n623 B.n450 71.676
R1077 B.n619 B.n451 71.676
R1078 B.n615 B.n452 71.676
R1079 B.n610 B.n453 71.676
R1080 B.n606 B.n454 71.676
R1081 B.n602 B.n455 71.676
R1082 B.n598 B.n456 71.676
R1083 B.n594 B.n457 71.676
R1084 B.n590 B.n458 71.676
R1085 B.n586 B.n459 71.676
R1086 B.n582 B.n460 71.676
R1087 B.n578 B.n461 71.676
R1088 B.n574 B.n462 71.676
R1089 B.n570 B.n463 71.676
R1090 B.n566 B.n464 71.676
R1091 B.n562 B.n465 71.676
R1092 B.n558 B.n466 71.676
R1093 B.n554 B.n467 71.676
R1094 B.n550 B.n468 71.676
R1095 B.n546 B.n469 71.676
R1096 B.n542 B.n470 71.676
R1097 B.n538 B.n471 71.676
R1098 B.n534 B.n472 71.676
R1099 B.n530 B.n473 71.676
R1100 B.n526 B.n474 71.676
R1101 B.n522 B.n475 71.676
R1102 B.n518 B.n476 71.676
R1103 B.n514 B.n477 71.676
R1104 B.n510 B.n478 71.676
R1105 B.n506 B.n479 71.676
R1106 B.n502 B.n480 71.676
R1107 B.n498 B.n481 71.676
R1108 B.n494 B.n482 71.676
R1109 B.n490 B.n483 71.676
R1110 B.n906 B.n905 71.676
R1111 B.n906 B.n2 71.676
R1112 B.n114 B.t7 70.3215
R1113 B.n489 B.t10 70.3215
R1114 B.n117 B.t17 70.2968
R1115 B.n486 B.t13 70.2968
R1116 B.n236 B.n117 59.5399
R1117 B.n115 B.n114 59.5399
R1118 B.n612 B.n489 59.5399
R1119 B.n487 B.n486 59.5399
R1120 B.n748 B.n416 50.3892
R1121 B.n854 B.n43 50.3892
R1122 B.n117 B.n116 33.3581
R1123 B.n114 B.n113 33.3581
R1124 B.n489 B.n488 33.3581
R1125 B.n486 B.n485 33.3581
R1126 B.n755 B.n416 31.4357
R1127 B.n755 B.n412 31.4357
R1128 B.n761 B.n412 31.4357
R1129 B.n761 B.n407 31.4357
R1130 B.n767 B.n407 31.4357
R1131 B.n767 B.n408 31.4357
R1132 B.n773 B.n400 31.4357
R1133 B.n779 B.n400 31.4357
R1134 B.n779 B.n396 31.4357
R1135 B.n785 B.n396 31.4357
R1136 B.n785 B.n391 31.4357
R1137 B.n791 B.n391 31.4357
R1138 B.n791 B.n392 31.4357
R1139 B.n797 B.n384 31.4357
R1140 B.n803 B.n384 31.4357
R1141 B.n803 B.n380 31.4357
R1142 B.n810 B.n380 31.4357
R1143 B.n816 B.n376 31.4357
R1144 B.n816 B.n4 31.4357
R1145 B.n904 B.n4 31.4357
R1146 B.n904 B.n903 31.4357
R1147 B.n903 B.n902 31.4357
R1148 B.n902 B.n8 31.4357
R1149 B.n825 B.n8 31.4357
R1150 B.n895 B.n894 31.4357
R1151 B.n894 B.n893 31.4357
R1152 B.n893 B.n15 31.4357
R1153 B.n887 B.n15 31.4357
R1154 B.n886 B.n885 31.4357
R1155 B.n885 B.n22 31.4357
R1156 B.n879 B.n22 31.4357
R1157 B.n879 B.n878 31.4357
R1158 B.n878 B.n877 31.4357
R1159 B.n877 B.n29 31.4357
R1160 B.n871 B.n29 31.4357
R1161 B.n870 B.n869 31.4357
R1162 B.n869 B.n36 31.4357
R1163 B.n863 B.n36 31.4357
R1164 B.n863 B.n862 31.4357
R1165 B.n862 B.n861 31.4357
R1166 B.n861 B.n43 31.4357
R1167 B.n752 B.n751 31.0639
R1168 B.n491 B.n414 31.0639
R1169 B.n852 B.n851 31.0639
R1170 B.n858 B.n857 31.0639
R1171 B.n773 B.t9 30.0488
R1172 B.n871 B.t5 30.0488
R1173 B.n797 B.t3 21.7278
R1174 B.n887 B.t1 21.7278
R1175 B.t0 B.n376 19.8786
R1176 B.n825 B.t2 19.8786
R1177 B B.n907 18.0485
R1178 B.n810 B.t0 11.5575
R1179 B.n895 B.t2 11.5575
R1180 B.n753 B.n752 10.6151
R1181 B.n753 B.n410 10.6151
R1182 B.n763 B.n410 10.6151
R1183 B.n764 B.n763 10.6151
R1184 B.n765 B.n764 10.6151
R1185 B.n765 B.n402 10.6151
R1186 B.n775 B.n402 10.6151
R1187 B.n776 B.n775 10.6151
R1188 B.n777 B.n776 10.6151
R1189 B.n777 B.n394 10.6151
R1190 B.n787 B.n394 10.6151
R1191 B.n788 B.n787 10.6151
R1192 B.n789 B.n788 10.6151
R1193 B.n789 B.n386 10.6151
R1194 B.n799 B.n386 10.6151
R1195 B.n800 B.n799 10.6151
R1196 B.n801 B.n800 10.6151
R1197 B.n801 B.n378 10.6151
R1198 B.n812 B.n378 10.6151
R1199 B.n813 B.n812 10.6151
R1200 B.n814 B.n813 10.6151
R1201 B.n814 B.n0 10.6151
R1202 B.n751 B.n418 10.6151
R1203 B.n746 B.n418 10.6151
R1204 B.n746 B.n745 10.6151
R1205 B.n745 B.n744 10.6151
R1206 B.n744 B.n741 10.6151
R1207 B.n741 B.n740 10.6151
R1208 B.n740 B.n737 10.6151
R1209 B.n737 B.n736 10.6151
R1210 B.n736 B.n733 10.6151
R1211 B.n733 B.n732 10.6151
R1212 B.n732 B.n729 10.6151
R1213 B.n729 B.n728 10.6151
R1214 B.n728 B.n725 10.6151
R1215 B.n725 B.n724 10.6151
R1216 B.n724 B.n721 10.6151
R1217 B.n721 B.n720 10.6151
R1218 B.n720 B.n717 10.6151
R1219 B.n717 B.n716 10.6151
R1220 B.n716 B.n713 10.6151
R1221 B.n713 B.n712 10.6151
R1222 B.n712 B.n709 10.6151
R1223 B.n709 B.n708 10.6151
R1224 B.n708 B.n705 10.6151
R1225 B.n705 B.n704 10.6151
R1226 B.n704 B.n701 10.6151
R1227 B.n701 B.n700 10.6151
R1228 B.n700 B.n697 10.6151
R1229 B.n697 B.n696 10.6151
R1230 B.n696 B.n693 10.6151
R1231 B.n693 B.n692 10.6151
R1232 B.n692 B.n689 10.6151
R1233 B.n689 B.n688 10.6151
R1234 B.n688 B.n685 10.6151
R1235 B.n685 B.n684 10.6151
R1236 B.n684 B.n681 10.6151
R1237 B.n681 B.n680 10.6151
R1238 B.n680 B.n677 10.6151
R1239 B.n677 B.n676 10.6151
R1240 B.n676 B.n673 10.6151
R1241 B.n673 B.n672 10.6151
R1242 B.n672 B.n669 10.6151
R1243 B.n669 B.n668 10.6151
R1244 B.n668 B.n665 10.6151
R1245 B.n665 B.n664 10.6151
R1246 B.n664 B.n661 10.6151
R1247 B.n661 B.n660 10.6151
R1248 B.n660 B.n657 10.6151
R1249 B.n657 B.n656 10.6151
R1250 B.n656 B.n653 10.6151
R1251 B.n653 B.n652 10.6151
R1252 B.n652 B.n649 10.6151
R1253 B.n649 B.n648 10.6151
R1254 B.n648 B.n645 10.6151
R1255 B.n645 B.n644 10.6151
R1256 B.n644 B.n641 10.6151
R1257 B.n641 B.n640 10.6151
R1258 B.n640 B.n637 10.6151
R1259 B.n637 B.n636 10.6151
R1260 B.n636 B.n633 10.6151
R1261 B.n633 B.n632 10.6151
R1262 B.n629 B.n628 10.6151
R1263 B.n628 B.n625 10.6151
R1264 B.n625 B.n624 10.6151
R1265 B.n624 B.n621 10.6151
R1266 B.n621 B.n620 10.6151
R1267 B.n620 B.n617 10.6151
R1268 B.n617 B.n616 10.6151
R1269 B.n616 B.n613 10.6151
R1270 B.n611 B.n608 10.6151
R1271 B.n608 B.n607 10.6151
R1272 B.n607 B.n604 10.6151
R1273 B.n604 B.n603 10.6151
R1274 B.n603 B.n600 10.6151
R1275 B.n600 B.n599 10.6151
R1276 B.n599 B.n596 10.6151
R1277 B.n596 B.n595 10.6151
R1278 B.n595 B.n592 10.6151
R1279 B.n592 B.n591 10.6151
R1280 B.n591 B.n588 10.6151
R1281 B.n588 B.n587 10.6151
R1282 B.n587 B.n584 10.6151
R1283 B.n584 B.n583 10.6151
R1284 B.n583 B.n580 10.6151
R1285 B.n580 B.n579 10.6151
R1286 B.n579 B.n576 10.6151
R1287 B.n576 B.n575 10.6151
R1288 B.n575 B.n572 10.6151
R1289 B.n572 B.n571 10.6151
R1290 B.n571 B.n568 10.6151
R1291 B.n568 B.n567 10.6151
R1292 B.n567 B.n564 10.6151
R1293 B.n564 B.n563 10.6151
R1294 B.n563 B.n560 10.6151
R1295 B.n560 B.n559 10.6151
R1296 B.n559 B.n556 10.6151
R1297 B.n556 B.n555 10.6151
R1298 B.n555 B.n552 10.6151
R1299 B.n552 B.n551 10.6151
R1300 B.n551 B.n548 10.6151
R1301 B.n548 B.n547 10.6151
R1302 B.n547 B.n544 10.6151
R1303 B.n544 B.n543 10.6151
R1304 B.n543 B.n540 10.6151
R1305 B.n540 B.n539 10.6151
R1306 B.n539 B.n536 10.6151
R1307 B.n536 B.n535 10.6151
R1308 B.n535 B.n532 10.6151
R1309 B.n532 B.n531 10.6151
R1310 B.n531 B.n528 10.6151
R1311 B.n528 B.n527 10.6151
R1312 B.n527 B.n524 10.6151
R1313 B.n524 B.n523 10.6151
R1314 B.n523 B.n520 10.6151
R1315 B.n520 B.n519 10.6151
R1316 B.n519 B.n516 10.6151
R1317 B.n516 B.n515 10.6151
R1318 B.n515 B.n512 10.6151
R1319 B.n512 B.n511 10.6151
R1320 B.n511 B.n508 10.6151
R1321 B.n508 B.n507 10.6151
R1322 B.n507 B.n504 10.6151
R1323 B.n504 B.n503 10.6151
R1324 B.n503 B.n500 10.6151
R1325 B.n500 B.n499 10.6151
R1326 B.n499 B.n496 10.6151
R1327 B.n496 B.n495 10.6151
R1328 B.n495 B.n492 10.6151
R1329 B.n492 B.n491 10.6151
R1330 B.n757 B.n414 10.6151
R1331 B.n758 B.n757 10.6151
R1332 B.n759 B.n758 10.6151
R1333 B.n759 B.n405 10.6151
R1334 B.n769 B.n405 10.6151
R1335 B.n770 B.n769 10.6151
R1336 B.n771 B.n770 10.6151
R1337 B.n771 B.n398 10.6151
R1338 B.n781 B.n398 10.6151
R1339 B.n782 B.n781 10.6151
R1340 B.n783 B.n782 10.6151
R1341 B.n783 B.n389 10.6151
R1342 B.n793 B.n389 10.6151
R1343 B.n794 B.n793 10.6151
R1344 B.n795 B.n794 10.6151
R1345 B.n795 B.n382 10.6151
R1346 B.n805 B.n382 10.6151
R1347 B.n806 B.n805 10.6151
R1348 B.n808 B.n806 10.6151
R1349 B.n808 B.n807 10.6151
R1350 B.n807 B.n374 10.6151
R1351 B.n819 B.n374 10.6151
R1352 B.n820 B.n819 10.6151
R1353 B.n821 B.n820 10.6151
R1354 B.n822 B.n821 10.6151
R1355 B.n823 B.n822 10.6151
R1356 B.n827 B.n823 10.6151
R1357 B.n828 B.n827 10.6151
R1358 B.n829 B.n828 10.6151
R1359 B.n830 B.n829 10.6151
R1360 B.n832 B.n830 10.6151
R1361 B.n833 B.n832 10.6151
R1362 B.n834 B.n833 10.6151
R1363 B.n835 B.n834 10.6151
R1364 B.n837 B.n835 10.6151
R1365 B.n838 B.n837 10.6151
R1366 B.n839 B.n838 10.6151
R1367 B.n840 B.n839 10.6151
R1368 B.n842 B.n840 10.6151
R1369 B.n843 B.n842 10.6151
R1370 B.n844 B.n843 10.6151
R1371 B.n845 B.n844 10.6151
R1372 B.n847 B.n845 10.6151
R1373 B.n848 B.n847 10.6151
R1374 B.n849 B.n848 10.6151
R1375 B.n850 B.n849 10.6151
R1376 B.n851 B.n850 10.6151
R1377 B.n899 B.n1 10.6151
R1378 B.n899 B.n898 10.6151
R1379 B.n898 B.n897 10.6151
R1380 B.n897 B.n10 10.6151
R1381 B.n891 B.n10 10.6151
R1382 B.n891 B.n890 10.6151
R1383 B.n890 B.n889 10.6151
R1384 B.n889 B.n17 10.6151
R1385 B.n883 B.n17 10.6151
R1386 B.n883 B.n882 10.6151
R1387 B.n882 B.n881 10.6151
R1388 B.n881 B.n24 10.6151
R1389 B.n875 B.n24 10.6151
R1390 B.n875 B.n874 10.6151
R1391 B.n874 B.n873 10.6151
R1392 B.n873 B.n31 10.6151
R1393 B.n867 B.n31 10.6151
R1394 B.n867 B.n866 10.6151
R1395 B.n866 B.n865 10.6151
R1396 B.n865 B.n38 10.6151
R1397 B.n859 B.n38 10.6151
R1398 B.n859 B.n858 10.6151
R1399 B.n857 B.n45 10.6151
R1400 B.n119 B.n45 10.6151
R1401 B.n120 B.n119 10.6151
R1402 B.n123 B.n120 10.6151
R1403 B.n124 B.n123 10.6151
R1404 B.n127 B.n124 10.6151
R1405 B.n128 B.n127 10.6151
R1406 B.n131 B.n128 10.6151
R1407 B.n132 B.n131 10.6151
R1408 B.n135 B.n132 10.6151
R1409 B.n136 B.n135 10.6151
R1410 B.n139 B.n136 10.6151
R1411 B.n140 B.n139 10.6151
R1412 B.n143 B.n140 10.6151
R1413 B.n144 B.n143 10.6151
R1414 B.n147 B.n144 10.6151
R1415 B.n148 B.n147 10.6151
R1416 B.n151 B.n148 10.6151
R1417 B.n152 B.n151 10.6151
R1418 B.n155 B.n152 10.6151
R1419 B.n156 B.n155 10.6151
R1420 B.n159 B.n156 10.6151
R1421 B.n160 B.n159 10.6151
R1422 B.n163 B.n160 10.6151
R1423 B.n164 B.n163 10.6151
R1424 B.n167 B.n164 10.6151
R1425 B.n168 B.n167 10.6151
R1426 B.n171 B.n168 10.6151
R1427 B.n172 B.n171 10.6151
R1428 B.n175 B.n172 10.6151
R1429 B.n176 B.n175 10.6151
R1430 B.n179 B.n176 10.6151
R1431 B.n180 B.n179 10.6151
R1432 B.n183 B.n180 10.6151
R1433 B.n184 B.n183 10.6151
R1434 B.n187 B.n184 10.6151
R1435 B.n188 B.n187 10.6151
R1436 B.n191 B.n188 10.6151
R1437 B.n192 B.n191 10.6151
R1438 B.n195 B.n192 10.6151
R1439 B.n196 B.n195 10.6151
R1440 B.n199 B.n196 10.6151
R1441 B.n200 B.n199 10.6151
R1442 B.n203 B.n200 10.6151
R1443 B.n204 B.n203 10.6151
R1444 B.n207 B.n204 10.6151
R1445 B.n208 B.n207 10.6151
R1446 B.n211 B.n208 10.6151
R1447 B.n212 B.n211 10.6151
R1448 B.n215 B.n212 10.6151
R1449 B.n216 B.n215 10.6151
R1450 B.n219 B.n216 10.6151
R1451 B.n220 B.n219 10.6151
R1452 B.n223 B.n220 10.6151
R1453 B.n224 B.n223 10.6151
R1454 B.n227 B.n224 10.6151
R1455 B.n228 B.n227 10.6151
R1456 B.n231 B.n228 10.6151
R1457 B.n232 B.n231 10.6151
R1458 B.n235 B.n232 10.6151
R1459 B.n240 B.n237 10.6151
R1460 B.n241 B.n240 10.6151
R1461 B.n244 B.n241 10.6151
R1462 B.n245 B.n244 10.6151
R1463 B.n248 B.n245 10.6151
R1464 B.n249 B.n248 10.6151
R1465 B.n252 B.n249 10.6151
R1466 B.n253 B.n252 10.6151
R1467 B.n257 B.n256 10.6151
R1468 B.n260 B.n257 10.6151
R1469 B.n261 B.n260 10.6151
R1470 B.n264 B.n261 10.6151
R1471 B.n265 B.n264 10.6151
R1472 B.n268 B.n265 10.6151
R1473 B.n269 B.n268 10.6151
R1474 B.n272 B.n269 10.6151
R1475 B.n273 B.n272 10.6151
R1476 B.n276 B.n273 10.6151
R1477 B.n277 B.n276 10.6151
R1478 B.n280 B.n277 10.6151
R1479 B.n281 B.n280 10.6151
R1480 B.n284 B.n281 10.6151
R1481 B.n285 B.n284 10.6151
R1482 B.n288 B.n285 10.6151
R1483 B.n289 B.n288 10.6151
R1484 B.n292 B.n289 10.6151
R1485 B.n293 B.n292 10.6151
R1486 B.n296 B.n293 10.6151
R1487 B.n297 B.n296 10.6151
R1488 B.n300 B.n297 10.6151
R1489 B.n301 B.n300 10.6151
R1490 B.n304 B.n301 10.6151
R1491 B.n305 B.n304 10.6151
R1492 B.n308 B.n305 10.6151
R1493 B.n309 B.n308 10.6151
R1494 B.n312 B.n309 10.6151
R1495 B.n313 B.n312 10.6151
R1496 B.n316 B.n313 10.6151
R1497 B.n317 B.n316 10.6151
R1498 B.n320 B.n317 10.6151
R1499 B.n321 B.n320 10.6151
R1500 B.n324 B.n321 10.6151
R1501 B.n325 B.n324 10.6151
R1502 B.n328 B.n325 10.6151
R1503 B.n329 B.n328 10.6151
R1504 B.n332 B.n329 10.6151
R1505 B.n333 B.n332 10.6151
R1506 B.n336 B.n333 10.6151
R1507 B.n337 B.n336 10.6151
R1508 B.n340 B.n337 10.6151
R1509 B.n341 B.n340 10.6151
R1510 B.n344 B.n341 10.6151
R1511 B.n345 B.n344 10.6151
R1512 B.n348 B.n345 10.6151
R1513 B.n349 B.n348 10.6151
R1514 B.n352 B.n349 10.6151
R1515 B.n353 B.n352 10.6151
R1516 B.n356 B.n353 10.6151
R1517 B.n357 B.n356 10.6151
R1518 B.n360 B.n357 10.6151
R1519 B.n361 B.n360 10.6151
R1520 B.n364 B.n361 10.6151
R1521 B.n365 B.n364 10.6151
R1522 B.n368 B.n365 10.6151
R1523 B.n369 B.n368 10.6151
R1524 B.n372 B.n369 10.6151
R1525 B.n373 B.n372 10.6151
R1526 B.n852 B.n373 10.6151
R1527 B.n392 B.t3 9.70842
R1528 B.t1 B.n886 9.70842
R1529 B.n907 B.n0 8.11757
R1530 B.n907 B.n1 8.11757
R1531 B.n629 B.n487 6.5566
R1532 B.n613 B.n612 6.5566
R1533 B.n237 B.n236 6.5566
R1534 B.n253 B.n115 6.5566
R1535 B.n632 B.n487 4.05904
R1536 B.n612 B.n611 4.05904
R1537 B.n236 B.n235 4.05904
R1538 B.n256 B.n115 4.05904
R1539 B.n408 B.t9 1.38735
R1540 B.t5 B.n870 1.38735
R1541 VP.n2 VP.t2 359.877
R1542 VP.n2 VP.t1 359.642
R1543 VP.n3 VP.t3 321.103
R1544 VP.n9 VP.t0 321.103
R1545 VP.n4 VP.n3 168.186
R1546 VP.n10 VP.n9 168.186
R1547 VP.n8 VP.n0 161.3
R1548 VP.n7 VP.n6 161.3
R1549 VP.n5 VP.n1 161.3
R1550 VP.n4 VP.n2 65.0455
R1551 VP.n7 VP.n1 40.577
R1552 VP.n8 VP.n7 40.577
R1553 VP.n3 VP.n1 17.7066
R1554 VP.n9 VP.n8 17.7066
R1555 VP.n5 VP.n4 0.189894
R1556 VP.n6 VP.n5 0.189894
R1557 VP.n6 VP.n0 0.189894
R1558 VP.n10 VP.n0 0.189894
R1559 VP VP.n10 0.0516364
R1560 VDD1 VDD1.n1 103.736
R1561 VDD1 VDD1.n0 59.1406
R1562 VDD1.n0 VDD1.t1 1.06961
R1563 VDD1.n0 VDD1.t2 1.06961
R1564 VDD1.n1 VDD1.t0 1.06961
R1565 VDD1.n1 VDD1.t3 1.06961
C0 VTAIL VN 5.60999f
C1 VN VDD2 6.16013f
C2 VTAIL VP 5.62409f
C3 VDD2 VP 0.317461f
C4 VN VDD1 0.148056f
C5 VTAIL VDD2 7.68635f
C6 VP VDD1 6.3291f
C7 VN VP 6.5197f
C8 VTAIL VDD1 7.64025f
C9 VDD2 VDD1 0.730623f
C10 VDD2 B 3.594375f
C11 VDD1 B 8.020861f
C12 VTAIL B 13.125081f
C13 VN B 9.42863f
C14 VP B 6.790532f
C15 VDD1.t1 B 0.389508f
C16 VDD1.t2 B 0.389508f
C17 VDD1.n0 B 3.55004f
C18 VDD1.t0 B 0.389508f
C19 VDD1.t3 B 0.389508f
C20 VDD1.n1 B 4.442f
C21 VP.n0 B 0.035985f
C22 VP.t0 B 2.54938f
C23 VP.n1 B 0.06192f
C24 VP.t2 B 2.66066f
C25 VP.t1 B 2.65998f
C26 VP.n2 B 3.33512f
C27 VP.t3 B 2.54938f
C28 VP.n3 B 0.97811f
C29 VP.n4 B 2.37547f
C30 VP.n5 B 0.035985f
C31 VP.n6 B 0.035985f
C32 VP.n7 B 0.029064f
C33 VP.n8 B 0.06192f
C34 VP.n9 B 0.97811f
C35 VP.n10 B 0.031294f
C36 VDD2.t0 B 0.392282f
C37 VDD2.t3 B 0.392282f
C38 VDD2.n0 B 4.444839f
C39 VDD2.t2 B 0.392282f
C40 VDD2.t1 B 0.392282f
C41 VDD2.n1 B 3.57496f
C42 VDD2.n2 B 4.17724f
C43 VTAIL.t4 B 2.49385f
C44 VTAIL.n0 B 0.27334f
C45 VTAIL.t0 B 2.49385f
C46 VTAIL.n1 B 0.306367f
C47 VTAIL.t3 B 2.49385f
C48 VTAIL.n2 B 1.33094f
C49 VTAIL.t7 B 2.49386f
C50 VTAIL.n3 B 1.33093f
C51 VTAIL.t5 B 2.49386f
C52 VTAIL.n4 B 0.306352f
C53 VTAIL.t2 B 2.49386f
C54 VTAIL.n5 B 0.306352f
C55 VTAIL.t1 B 2.49385f
C56 VTAIL.n6 B 1.33094f
C57 VTAIL.t6 B 2.49385f
C58 VTAIL.n7 B 1.29229f
C59 VN.t3 B 2.63895f
C60 VN.t0 B 2.63827f
C61 VN.n0 B 1.87435f
C62 VN.t2 B 2.63895f
C63 VN.t1 B 2.63827f
C64 VN.n1 B 3.32802f
.ends

