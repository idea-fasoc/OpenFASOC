* NGSPICE file created from diff_pair_sample_1689.ext - technology: sky130A

.subckt diff_pair_sample_1689 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=1.1616 ps=7.37 w=7.04 l=1.88
X1 VTAIL.t5 VP.t0 VDD1.t5 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=1.1616 ps=7.37 w=7.04 l=1.88
X2 VDD2.t4 VN.t1 VTAIL.t6 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=1.1616 ps=7.37 w=7.04 l=1.88
X3 VDD1.t4 VP.t1 VTAIL.t1 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=2.7456 ps=14.86 w=7.04 l=1.88
X4 VDD2.t3 VN.t2 VTAIL.t10 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=2.7456 ps=14.86 w=7.04 l=1.88
X5 B.t11 B.t9 B.t10 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=0 ps=0 w=7.04 l=1.88
X6 VTAIL.t9 VN.t3 VDD2.t2 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=1.1616 ps=7.37 w=7.04 l=1.88
X7 VDD1.t3 VP.t2 VTAIL.t3 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=2.7456 ps=14.86 w=7.04 l=1.88
X8 VDD2.t1 VN.t4 VTAIL.t8 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=2.7456 ps=14.86 w=7.04 l=1.88
X9 VTAIL.t0 VP.t3 VDD1.t2 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=1.1616 ps=7.37 w=7.04 l=1.88
X10 VTAIL.t11 VN.t5 VDD2.t0 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=1.1616 pd=7.37 as=1.1616 ps=7.37 w=7.04 l=1.88
X11 B.t8 B.t6 B.t7 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=0 ps=0 w=7.04 l=1.88
X12 VDD1.t1 VP.t4 VTAIL.t2 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=1.1616 ps=7.37 w=7.04 l=1.88
X13 B.t5 B.t3 B.t4 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=0 ps=0 w=7.04 l=1.88
X14 B.t2 B.t0 B.t1 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=0 ps=0 w=7.04 l=1.88
X15 VDD1.t0 VP.t5 VTAIL.t4 w_n2738_n2376# sky130_fd_pr__pfet_01v8 ad=2.7456 pd=14.86 as=1.1616 ps=7.37 w=7.04 l=1.88
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n2 VN.t1 121.297
R9 VN.n14 VN.t2 121.297
R10 VN.n3 VN.t3 90.2473
R11 VN.n10 VN.t4 90.2473
R12 VN.n15 VN.t5 90.2473
R13 VN.n22 VN.t0 90.2473
R14 VN.n11 VN.n10 88.2837
R15 VN.n23 VN.n22 88.2837
R16 VN.n3 VN.n2 57.9446
R17 VN.n15 VN.n14 57.9446
R18 VN.n8 VN.n1 54.6242
R19 VN.n20 VN.n13 54.6242
R20 VN VN.n23 42.4111
R21 VN.n9 VN.n8 26.5299
R22 VN.n21 VN.n20 26.5299
R23 VN.n4 VN.n1 24.5923
R24 VN.n16 VN.n13 24.5923
R25 VN.n10 VN.n9 22.625
R26 VN.n22 VN.n21 22.625
R27 VN.n17 VN.n14 12.9017
R28 VN.n5 VN.n2 12.9017
R29 VN.n4 VN.n3 12.2964
R30 VN.n16 VN.n15 12.2964
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VTAIL.n7 VTAIL.t10 73.9288
R41 VTAIL.n11 VTAIL.t8 73.9285
R42 VTAIL.n2 VTAIL.t3 73.9285
R43 VTAIL.n10 VTAIL.t1 73.9285
R44 VTAIL.n9 VTAIL.n8 69.3116
R45 VTAIL.n6 VTAIL.n5 69.3116
R46 VTAIL.n1 VTAIL.n0 69.3115
R47 VTAIL.n4 VTAIL.n3 69.3115
R48 VTAIL.n6 VTAIL.n4 22.2462
R49 VTAIL.n11 VTAIL.n10 20.341
R50 VTAIL.n0 VTAIL.t6 4.61769
R51 VTAIL.n0 VTAIL.t9 4.61769
R52 VTAIL.n3 VTAIL.t2 4.61769
R53 VTAIL.n3 VTAIL.t0 4.61769
R54 VTAIL.n8 VTAIL.t4 4.61769
R55 VTAIL.n8 VTAIL.t5 4.61769
R56 VTAIL.n5 VTAIL.t7 4.61769
R57 VTAIL.n5 VTAIL.t11 4.61769
R58 VTAIL.n7 VTAIL.n6 1.90567
R59 VTAIL.n10 VTAIL.n9 1.90567
R60 VTAIL.n4 VTAIL.n2 1.90567
R61 VTAIL.n9 VTAIL.n7 1.42291
R62 VTAIL.n2 VTAIL.n1 1.42291
R63 VTAIL VTAIL.n11 1.37119
R64 VTAIL VTAIL.n1 0.534983
R65 VDD2.n1 VDD2.t4 91.9809
R66 VDD2.n2 VDD2.t5 90.6076
R67 VDD2.n1 VDD2.n0 86.4113
R68 VDD2 VDD2.n3 86.4083
R69 VDD2.n2 VDD2.n1 35.9761
R70 VDD2.n3 VDD2.t0 4.61769
R71 VDD2.n3 VDD2.t3 4.61769
R72 VDD2.n0 VDD2.t2 4.61769
R73 VDD2.n0 VDD2.t1 4.61769
R74 VDD2 VDD2.n2 1.48757
R75 VP.n9 VP.n8 161.3
R76 VP.n10 VP.n5 161.3
R77 VP.n12 VP.n11 161.3
R78 VP.n13 VP.n4 161.3
R79 VP.n30 VP.n0 161.3
R80 VP.n29 VP.n28 161.3
R81 VP.n27 VP.n1 161.3
R82 VP.n26 VP.n25 161.3
R83 VP.n23 VP.n2 161.3
R84 VP.n22 VP.n21 161.3
R85 VP.n20 VP.n3 161.3
R86 VP.n19 VP.n18 161.3
R87 VP.n6 VP.t5 121.297
R88 VP.n17 VP.t4 90.2473
R89 VP.n24 VP.t3 90.2473
R90 VP.n31 VP.t2 90.2473
R91 VP.n14 VP.t1 90.2473
R92 VP.n7 VP.t0 90.2473
R93 VP.n17 VP.n16 88.2837
R94 VP.n32 VP.n31 88.2837
R95 VP.n15 VP.n14 88.2837
R96 VP.n7 VP.n6 57.9446
R97 VP.n22 VP.n3 54.6242
R98 VP.n29 VP.n1 54.6242
R99 VP.n12 VP.n5 54.6242
R100 VP.n16 VP.n15 42.1322
R101 VP.n18 VP.n3 26.5299
R102 VP.n30 VP.n29 26.5299
R103 VP.n13 VP.n12 26.5299
R104 VP.n23 VP.n22 24.5923
R105 VP.n25 VP.n1 24.5923
R106 VP.n8 VP.n5 24.5923
R107 VP.n18 VP.n17 22.625
R108 VP.n31 VP.n30 22.625
R109 VP.n14 VP.n13 22.625
R110 VP.n9 VP.n6 12.9017
R111 VP.n24 VP.n23 12.2964
R112 VP.n25 VP.n24 12.2964
R113 VP.n8 VP.n7 12.2964
R114 VP.n15 VP.n4 0.278335
R115 VP.n19 VP.n16 0.278335
R116 VP.n32 VP.n0 0.278335
R117 VP.n10 VP.n9 0.189894
R118 VP.n11 VP.n10 0.189894
R119 VP.n11 VP.n4 0.189894
R120 VP.n20 VP.n19 0.189894
R121 VP.n21 VP.n20 0.189894
R122 VP.n21 VP.n2 0.189894
R123 VP.n26 VP.n2 0.189894
R124 VP.n27 VP.n26 0.189894
R125 VP.n28 VP.n27 0.189894
R126 VP.n28 VP.n0 0.189894
R127 VP VP.n32 0.153485
R128 VDD1 VDD1.t0 92.0946
R129 VDD1.n1 VDD1.t1 91.9809
R130 VDD1.n1 VDD1.n0 86.4113
R131 VDD1.n3 VDD1.n2 85.9902
R132 VDD1.n3 VDD1.n1 37.5117
R133 VDD1.n2 VDD1.t5 4.61769
R134 VDD1.n2 VDD1.t4 4.61769
R135 VDD1.n0 VDD1.t2 4.61769
R136 VDD1.n0 VDD1.t3 4.61769
R137 VDD1 VDD1.n3 0.418603
R138 B.n395 B.n394 585
R139 B.n396 B.n55 585
R140 B.n398 B.n397 585
R141 B.n399 B.n54 585
R142 B.n401 B.n400 585
R143 B.n402 B.n53 585
R144 B.n404 B.n403 585
R145 B.n405 B.n52 585
R146 B.n407 B.n406 585
R147 B.n408 B.n51 585
R148 B.n410 B.n409 585
R149 B.n411 B.n50 585
R150 B.n413 B.n412 585
R151 B.n414 B.n49 585
R152 B.n416 B.n415 585
R153 B.n417 B.n48 585
R154 B.n419 B.n418 585
R155 B.n420 B.n47 585
R156 B.n422 B.n421 585
R157 B.n423 B.n46 585
R158 B.n425 B.n424 585
R159 B.n426 B.n45 585
R160 B.n428 B.n427 585
R161 B.n429 B.n44 585
R162 B.n431 B.n430 585
R163 B.n432 B.n43 585
R164 B.n434 B.n433 585
R165 B.n436 B.n40 585
R166 B.n438 B.n437 585
R167 B.n439 B.n39 585
R168 B.n441 B.n440 585
R169 B.n442 B.n38 585
R170 B.n444 B.n443 585
R171 B.n445 B.n37 585
R172 B.n447 B.n446 585
R173 B.n448 B.n33 585
R174 B.n450 B.n449 585
R175 B.n451 B.n32 585
R176 B.n453 B.n452 585
R177 B.n454 B.n31 585
R178 B.n456 B.n455 585
R179 B.n457 B.n30 585
R180 B.n459 B.n458 585
R181 B.n460 B.n29 585
R182 B.n462 B.n461 585
R183 B.n463 B.n28 585
R184 B.n465 B.n464 585
R185 B.n466 B.n27 585
R186 B.n468 B.n467 585
R187 B.n469 B.n26 585
R188 B.n471 B.n470 585
R189 B.n472 B.n25 585
R190 B.n474 B.n473 585
R191 B.n475 B.n24 585
R192 B.n477 B.n476 585
R193 B.n478 B.n23 585
R194 B.n480 B.n479 585
R195 B.n481 B.n22 585
R196 B.n483 B.n482 585
R197 B.n484 B.n21 585
R198 B.n486 B.n485 585
R199 B.n487 B.n20 585
R200 B.n489 B.n488 585
R201 B.n490 B.n19 585
R202 B.n393 B.n56 585
R203 B.n392 B.n391 585
R204 B.n390 B.n57 585
R205 B.n389 B.n388 585
R206 B.n387 B.n58 585
R207 B.n386 B.n385 585
R208 B.n384 B.n59 585
R209 B.n383 B.n382 585
R210 B.n381 B.n60 585
R211 B.n380 B.n379 585
R212 B.n378 B.n61 585
R213 B.n377 B.n376 585
R214 B.n375 B.n62 585
R215 B.n374 B.n373 585
R216 B.n372 B.n63 585
R217 B.n371 B.n370 585
R218 B.n369 B.n64 585
R219 B.n368 B.n367 585
R220 B.n366 B.n65 585
R221 B.n365 B.n364 585
R222 B.n363 B.n66 585
R223 B.n362 B.n361 585
R224 B.n360 B.n67 585
R225 B.n359 B.n358 585
R226 B.n357 B.n68 585
R227 B.n356 B.n355 585
R228 B.n354 B.n69 585
R229 B.n353 B.n352 585
R230 B.n351 B.n70 585
R231 B.n350 B.n349 585
R232 B.n348 B.n71 585
R233 B.n347 B.n346 585
R234 B.n345 B.n72 585
R235 B.n344 B.n343 585
R236 B.n342 B.n73 585
R237 B.n341 B.n340 585
R238 B.n339 B.n74 585
R239 B.n338 B.n337 585
R240 B.n336 B.n75 585
R241 B.n335 B.n334 585
R242 B.n333 B.n76 585
R243 B.n332 B.n331 585
R244 B.n330 B.n77 585
R245 B.n329 B.n328 585
R246 B.n327 B.n78 585
R247 B.n326 B.n325 585
R248 B.n324 B.n79 585
R249 B.n323 B.n322 585
R250 B.n321 B.n80 585
R251 B.n320 B.n319 585
R252 B.n318 B.n81 585
R253 B.n317 B.n316 585
R254 B.n315 B.n82 585
R255 B.n314 B.n313 585
R256 B.n312 B.n83 585
R257 B.n311 B.n310 585
R258 B.n309 B.n84 585
R259 B.n308 B.n307 585
R260 B.n306 B.n85 585
R261 B.n305 B.n304 585
R262 B.n303 B.n86 585
R263 B.n302 B.n301 585
R264 B.n300 B.n87 585
R265 B.n299 B.n298 585
R266 B.n297 B.n88 585
R267 B.n296 B.n295 585
R268 B.n294 B.n89 585
R269 B.n293 B.n292 585
R270 B.n291 B.n90 585
R271 B.n194 B.n193 585
R272 B.n195 B.n126 585
R273 B.n197 B.n196 585
R274 B.n198 B.n125 585
R275 B.n200 B.n199 585
R276 B.n201 B.n124 585
R277 B.n203 B.n202 585
R278 B.n204 B.n123 585
R279 B.n206 B.n205 585
R280 B.n207 B.n122 585
R281 B.n209 B.n208 585
R282 B.n210 B.n121 585
R283 B.n212 B.n211 585
R284 B.n213 B.n120 585
R285 B.n215 B.n214 585
R286 B.n216 B.n119 585
R287 B.n218 B.n217 585
R288 B.n219 B.n118 585
R289 B.n221 B.n220 585
R290 B.n222 B.n117 585
R291 B.n224 B.n223 585
R292 B.n225 B.n116 585
R293 B.n227 B.n226 585
R294 B.n228 B.n115 585
R295 B.n230 B.n229 585
R296 B.n231 B.n114 585
R297 B.n233 B.n232 585
R298 B.n235 B.n234 585
R299 B.n236 B.n110 585
R300 B.n238 B.n237 585
R301 B.n239 B.n109 585
R302 B.n241 B.n240 585
R303 B.n242 B.n108 585
R304 B.n244 B.n243 585
R305 B.n245 B.n107 585
R306 B.n247 B.n246 585
R307 B.n248 B.n104 585
R308 B.n251 B.n250 585
R309 B.n252 B.n103 585
R310 B.n254 B.n253 585
R311 B.n255 B.n102 585
R312 B.n257 B.n256 585
R313 B.n258 B.n101 585
R314 B.n260 B.n259 585
R315 B.n261 B.n100 585
R316 B.n263 B.n262 585
R317 B.n264 B.n99 585
R318 B.n266 B.n265 585
R319 B.n267 B.n98 585
R320 B.n269 B.n268 585
R321 B.n270 B.n97 585
R322 B.n272 B.n271 585
R323 B.n273 B.n96 585
R324 B.n275 B.n274 585
R325 B.n276 B.n95 585
R326 B.n278 B.n277 585
R327 B.n279 B.n94 585
R328 B.n281 B.n280 585
R329 B.n282 B.n93 585
R330 B.n284 B.n283 585
R331 B.n285 B.n92 585
R332 B.n287 B.n286 585
R333 B.n288 B.n91 585
R334 B.n290 B.n289 585
R335 B.n192 B.n127 585
R336 B.n191 B.n190 585
R337 B.n189 B.n128 585
R338 B.n188 B.n187 585
R339 B.n186 B.n129 585
R340 B.n185 B.n184 585
R341 B.n183 B.n130 585
R342 B.n182 B.n181 585
R343 B.n180 B.n131 585
R344 B.n179 B.n178 585
R345 B.n177 B.n132 585
R346 B.n176 B.n175 585
R347 B.n174 B.n133 585
R348 B.n173 B.n172 585
R349 B.n171 B.n134 585
R350 B.n170 B.n169 585
R351 B.n168 B.n135 585
R352 B.n167 B.n166 585
R353 B.n165 B.n136 585
R354 B.n164 B.n163 585
R355 B.n162 B.n137 585
R356 B.n161 B.n160 585
R357 B.n159 B.n138 585
R358 B.n158 B.n157 585
R359 B.n156 B.n139 585
R360 B.n155 B.n154 585
R361 B.n153 B.n140 585
R362 B.n152 B.n151 585
R363 B.n150 B.n141 585
R364 B.n149 B.n148 585
R365 B.n147 B.n142 585
R366 B.n146 B.n145 585
R367 B.n144 B.n143 585
R368 B.n2 B.n0 585
R369 B.n541 B.n1 585
R370 B.n540 B.n539 585
R371 B.n538 B.n3 585
R372 B.n537 B.n536 585
R373 B.n535 B.n4 585
R374 B.n534 B.n533 585
R375 B.n532 B.n5 585
R376 B.n531 B.n530 585
R377 B.n529 B.n6 585
R378 B.n528 B.n527 585
R379 B.n526 B.n7 585
R380 B.n525 B.n524 585
R381 B.n523 B.n8 585
R382 B.n522 B.n521 585
R383 B.n520 B.n9 585
R384 B.n519 B.n518 585
R385 B.n517 B.n10 585
R386 B.n516 B.n515 585
R387 B.n514 B.n11 585
R388 B.n513 B.n512 585
R389 B.n511 B.n12 585
R390 B.n510 B.n509 585
R391 B.n508 B.n13 585
R392 B.n507 B.n506 585
R393 B.n505 B.n14 585
R394 B.n504 B.n503 585
R395 B.n502 B.n15 585
R396 B.n501 B.n500 585
R397 B.n499 B.n16 585
R398 B.n498 B.n497 585
R399 B.n496 B.n17 585
R400 B.n495 B.n494 585
R401 B.n493 B.n18 585
R402 B.n492 B.n491 585
R403 B.n543 B.n542 585
R404 B.n193 B.n192 487.695
R405 B.n492 B.n19 487.695
R406 B.n289 B.n90 487.695
R407 B.n395 B.n56 487.695
R408 B.n105 B.t3 296.868
R409 B.n111 B.t6 296.868
R410 B.n34 B.t0 296.868
R411 B.n41 B.t9 296.868
R412 B.n192 B.n191 163.367
R413 B.n191 B.n128 163.367
R414 B.n187 B.n128 163.367
R415 B.n187 B.n186 163.367
R416 B.n186 B.n185 163.367
R417 B.n185 B.n130 163.367
R418 B.n181 B.n130 163.367
R419 B.n181 B.n180 163.367
R420 B.n180 B.n179 163.367
R421 B.n179 B.n132 163.367
R422 B.n175 B.n132 163.367
R423 B.n175 B.n174 163.367
R424 B.n174 B.n173 163.367
R425 B.n173 B.n134 163.367
R426 B.n169 B.n134 163.367
R427 B.n169 B.n168 163.367
R428 B.n168 B.n167 163.367
R429 B.n167 B.n136 163.367
R430 B.n163 B.n136 163.367
R431 B.n163 B.n162 163.367
R432 B.n162 B.n161 163.367
R433 B.n161 B.n138 163.367
R434 B.n157 B.n138 163.367
R435 B.n157 B.n156 163.367
R436 B.n156 B.n155 163.367
R437 B.n155 B.n140 163.367
R438 B.n151 B.n140 163.367
R439 B.n151 B.n150 163.367
R440 B.n150 B.n149 163.367
R441 B.n149 B.n142 163.367
R442 B.n145 B.n142 163.367
R443 B.n145 B.n144 163.367
R444 B.n144 B.n2 163.367
R445 B.n542 B.n2 163.367
R446 B.n542 B.n541 163.367
R447 B.n541 B.n540 163.367
R448 B.n540 B.n3 163.367
R449 B.n536 B.n3 163.367
R450 B.n536 B.n535 163.367
R451 B.n535 B.n534 163.367
R452 B.n534 B.n5 163.367
R453 B.n530 B.n5 163.367
R454 B.n530 B.n529 163.367
R455 B.n529 B.n528 163.367
R456 B.n528 B.n7 163.367
R457 B.n524 B.n7 163.367
R458 B.n524 B.n523 163.367
R459 B.n523 B.n522 163.367
R460 B.n522 B.n9 163.367
R461 B.n518 B.n9 163.367
R462 B.n518 B.n517 163.367
R463 B.n517 B.n516 163.367
R464 B.n516 B.n11 163.367
R465 B.n512 B.n11 163.367
R466 B.n512 B.n511 163.367
R467 B.n511 B.n510 163.367
R468 B.n510 B.n13 163.367
R469 B.n506 B.n13 163.367
R470 B.n506 B.n505 163.367
R471 B.n505 B.n504 163.367
R472 B.n504 B.n15 163.367
R473 B.n500 B.n15 163.367
R474 B.n500 B.n499 163.367
R475 B.n499 B.n498 163.367
R476 B.n498 B.n17 163.367
R477 B.n494 B.n17 163.367
R478 B.n494 B.n493 163.367
R479 B.n493 B.n492 163.367
R480 B.n193 B.n126 163.367
R481 B.n197 B.n126 163.367
R482 B.n198 B.n197 163.367
R483 B.n199 B.n198 163.367
R484 B.n199 B.n124 163.367
R485 B.n203 B.n124 163.367
R486 B.n204 B.n203 163.367
R487 B.n205 B.n204 163.367
R488 B.n205 B.n122 163.367
R489 B.n209 B.n122 163.367
R490 B.n210 B.n209 163.367
R491 B.n211 B.n210 163.367
R492 B.n211 B.n120 163.367
R493 B.n215 B.n120 163.367
R494 B.n216 B.n215 163.367
R495 B.n217 B.n216 163.367
R496 B.n217 B.n118 163.367
R497 B.n221 B.n118 163.367
R498 B.n222 B.n221 163.367
R499 B.n223 B.n222 163.367
R500 B.n223 B.n116 163.367
R501 B.n227 B.n116 163.367
R502 B.n228 B.n227 163.367
R503 B.n229 B.n228 163.367
R504 B.n229 B.n114 163.367
R505 B.n233 B.n114 163.367
R506 B.n234 B.n233 163.367
R507 B.n234 B.n110 163.367
R508 B.n238 B.n110 163.367
R509 B.n239 B.n238 163.367
R510 B.n240 B.n239 163.367
R511 B.n240 B.n108 163.367
R512 B.n244 B.n108 163.367
R513 B.n245 B.n244 163.367
R514 B.n246 B.n245 163.367
R515 B.n246 B.n104 163.367
R516 B.n251 B.n104 163.367
R517 B.n252 B.n251 163.367
R518 B.n253 B.n252 163.367
R519 B.n253 B.n102 163.367
R520 B.n257 B.n102 163.367
R521 B.n258 B.n257 163.367
R522 B.n259 B.n258 163.367
R523 B.n259 B.n100 163.367
R524 B.n263 B.n100 163.367
R525 B.n264 B.n263 163.367
R526 B.n265 B.n264 163.367
R527 B.n265 B.n98 163.367
R528 B.n269 B.n98 163.367
R529 B.n270 B.n269 163.367
R530 B.n271 B.n270 163.367
R531 B.n271 B.n96 163.367
R532 B.n275 B.n96 163.367
R533 B.n276 B.n275 163.367
R534 B.n277 B.n276 163.367
R535 B.n277 B.n94 163.367
R536 B.n281 B.n94 163.367
R537 B.n282 B.n281 163.367
R538 B.n283 B.n282 163.367
R539 B.n283 B.n92 163.367
R540 B.n287 B.n92 163.367
R541 B.n288 B.n287 163.367
R542 B.n289 B.n288 163.367
R543 B.n293 B.n90 163.367
R544 B.n294 B.n293 163.367
R545 B.n295 B.n294 163.367
R546 B.n295 B.n88 163.367
R547 B.n299 B.n88 163.367
R548 B.n300 B.n299 163.367
R549 B.n301 B.n300 163.367
R550 B.n301 B.n86 163.367
R551 B.n305 B.n86 163.367
R552 B.n306 B.n305 163.367
R553 B.n307 B.n306 163.367
R554 B.n307 B.n84 163.367
R555 B.n311 B.n84 163.367
R556 B.n312 B.n311 163.367
R557 B.n313 B.n312 163.367
R558 B.n313 B.n82 163.367
R559 B.n317 B.n82 163.367
R560 B.n318 B.n317 163.367
R561 B.n319 B.n318 163.367
R562 B.n319 B.n80 163.367
R563 B.n323 B.n80 163.367
R564 B.n324 B.n323 163.367
R565 B.n325 B.n324 163.367
R566 B.n325 B.n78 163.367
R567 B.n329 B.n78 163.367
R568 B.n330 B.n329 163.367
R569 B.n331 B.n330 163.367
R570 B.n331 B.n76 163.367
R571 B.n335 B.n76 163.367
R572 B.n336 B.n335 163.367
R573 B.n337 B.n336 163.367
R574 B.n337 B.n74 163.367
R575 B.n341 B.n74 163.367
R576 B.n342 B.n341 163.367
R577 B.n343 B.n342 163.367
R578 B.n343 B.n72 163.367
R579 B.n347 B.n72 163.367
R580 B.n348 B.n347 163.367
R581 B.n349 B.n348 163.367
R582 B.n349 B.n70 163.367
R583 B.n353 B.n70 163.367
R584 B.n354 B.n353 163.367
R585 B.n355 B.n354 163.367
R586 B.n355 B.n68 163.367
R587 B.n359 B.n68 163.367
R588 B.n360 B.n359 163.367
R589 B.n361 B.n360 163.367
R590 B.n361 B.n66 163.367
R591 B.n365 B.n66 163.367
R592 B.n366 B.n365 163.367
R593 B.n367 B.n366 163.367
R594 B.n367 B.n64 163.367
R595 B.n371 B.n64 163.367
R596 B.n372 B.n371 163.367
R597 B.n373 B.n372 163.367
R598 B.n373 B.n62 163.367
R599 B.n377 B.n62 163.367
R600 B.n378 B.n377 163.367
R601 B.n379 B.n378 163.367
R602 B.n379 B.n60 163.367
R603 B.n383 B.n60 163.367
R604 B.n384 B.n383 163.367
R605 B.n385 B.n384 163.367
R606 B.n385 B.n58 163.367
R607 B.n389 B.n58 163.367
R608 B.n390 B.n389 163.367
R609 B.n391 B.n390 163.367
R610 B.n391 B.n56 163.367
R611 B.n488 B.n19 163.367
R612 B.n488 B.n487 163.367
R613 B.n487 B.n486 163.367
R614 B.n486 B.n21 163.367
R615 B.n482 B.n21 163.367
R616 B.n482 B.n481 163.367
R617 B.n481 B.n480 163.367
R618 B.n480 B.n23 163.367
R619 B.n476 B.n23 163.367
R620 B.n476 B.n475 163.367
R621 B.n475 B.n474 163.367
R622 B.n474 B.n25 163.367
R623 B.n470 B.n25 163.367
R624 B.n470 B.n469 163.367
R625 B.n469 B.n468 163.367
R626 B.n468 B.n27 163.367
R627 B.n464 B.n27 163.367
R628 B.n464 B.n463 163.367
R629 B.n463 B.n462 163.367
R630 B.n462 B.n29 163.367
R631 B.n458 B.n29 163.367
R632 B.n458 B.n457 163.367
R633 B.n457 B.n456 163.367
R634 B.n456 B.n31 163.367
R635 B.n452 B.n31 163.367
R636 B.n452 B.n451 163.367
R637 B.n451 B.n450 163.367
R638 B.n450 B.n33 163.367
R639 B.n446 B.n33 163.367
R640 B.n446 B.n445 163.367
R641 B.n445 B.n444 163.367
R642 B.n444 B.n38 163.367
R643 B.n440 B.n38 163.367
R644 B.n440 B.n439 163.367
R645 B.n439 B.n438 163.367
R646 B.n438 B.n40 163.367
R647 B.n433 B.n40 163.367
R648 B.n433 B.n432 163.367
R649 B.n432 B.n431 163.367
R650 B.n431 B.n44 163.367
R651 B.n427 B.n44 163.367
R652 B.n427 B.n426 163.367
R653 B.n426 B.n425 163.367
R654 B.n425 B.n46 163.367
R655 B.n421 B.n46 163.367
R656 B.n421 B.n420 163.367
R657 B.n420 B.n419 163.367
R658 B.n419 B.n48 163.367
R659 B.n415 B.n48 163.367
R660 B.n415 B.n414 163.367
R661 B.n414 B.n413 163.367
R662 B.n413 B.n50 163.367
R663 B.n409 B.n50 163.367
R664 B.n409 B.n408 163.367
R665 B.n408 B.n407 163.367
R666 B.n407 B.n52 163.367
R667 B.n403 B.n52 163.367
R668 B.n403 B.n402 163.367
R669 B.n402 B.n401 163.367
R670 B.n401 B.n54 163.367
R671 B.n397 B.n54 163.367
R672 B.n397 B.n396 163.367
R673 B.n396 B.n395 163.367
R674 B.n105 B.t5 157.106
R675 B.n41 B.t10 157.106
R676 B.n111 B.t8 157.099
R677 B.n34 B.t1 157.099
R678 B.n106 B.t4 114.246
R679 B.n42 B.t11 114.246
R680 B.n112 B.t7 114.237
R681 B.n35 B.t2 114.237
R682 B.n249 B.n106 59.5399
R683 B.n113 B.n112 59.5399
R684 B.n36 B.n35 59.5399
R685 B.n435 B.n42 59.5399
R686 B.n106 B.n105 42.8611
R687 B.n112 B.n111 42.8611
R688 B.n35 B.n34 42.8611
R689 B.n42 B.n41 42.8611
R690 B.n491 B.n490 31.6883
R691 B.n394 B.n393 31.6883
R692 B.n291 B.n290 31.6883
R693 B.n194 B.n127 31.6883
R694 B B.n543 18.0485
R695 B.n490 B.n489 10.6151
R696 B.n489 B.n20 10.6151
R697 B.n485 B.n20 10.6151
R698 B.n485 B.n484 10.6151
R699 B.n484 B.n483 10.6151
R700 B.n483 B.n22 10.6151
R701 B.n479 B.n22 10.6151
R702 B.n479 B.n478 10.6151
R703 B.n478 B.n477 10.6151
R704 B.n477 B.n24 10.6151
R705 B.n473 B.n24 10.6151
R706 B.n473 B.n472 10.6151
R707 B.n472 B.n471 10.6151
R708 B.n471 B.n26 10.6151
R709 B.n467 B.n26 10.6151
R710 B.n467 B.n466 10.6151
R711 B.n466 B.n465 10.6151
R712 B.n465 B.n28 10.6151
R713 B.n461 B.n28 10.6151
R714 B.n461 B.n460 10.6151
R715 B.n460 B.n459 10.6151
R716 B.n459 B.n30 10.6151
R717 B.n455 B.n30 10.6151
R718 B.n455 B.n454 10.6151
R719 B.n454 B.n453 10.6151
R720 B.n453 B.n32 10.6151
R721 B.n449 B.n448 10.6151
R722 B.n448 B.n447 10.6151
R723 B.n447 B.n37 10.6151
R724 B.n443 B.n37 10.6151
R725 B.n443 B.n442 10.6151
R726 B.n442 B.n441 10.6151
R727 B.n441 B.n39 10.6151
R728 B.n437 B.n39 10.6151
R729 B.n437 B.n436 10.6151
R730 B.n434 B.n43 10.6151
R731 B.n430 B.n43 10.6151
R732 B.n430 B.n429 10.6151
R733 B.n429 B.n428 10.6151
R734 B.n428 B.n45 10.6151
R735 B.n424 B.n45 10.6151
R736 B.n424 B.n423 10.6151
R737 B.n423 B.n422 10.6151
R738 B.n422 B.n47 10.6151
R739 B.n418 B.n47 10.6151
R740 B.n418 B.n417 10.6151
R741 B.n417 B.n416 10.6151
R742 B.n416 B.n49 10.6151
R743 B.n412 B.n49 10.6151
R744 B.n412 B.n411 10.6151
R745 B.n411 B.n410 10.6151
R746 B.n410 B.n51 10.6151
R747 B.n406 B.n51 10.6151
R748 B.n406 B.n405 10.6151
R749 B.n405 B.n404 10.6151
R750 B.n404 B.n53 10.6151
R751 B.n400 B.n53 10.6151
R752 B.n400 B.n399 10.6151
R753 B.n399 B.n398 10.6151
R754 B.n398 B.n55 10.6151
R755 B.n394 B.n55 10.6151
R756 B.n292 B.n291 10.6151
R757 B.n292 B.n89 10.6151
R758 B.n296 B.n89 10.6151
R759 B.n297 B.n296 10.6151
R760 B.n298 B.n297 10.6151
R761 B.n298 B.n87 10.6151
R762 B.n302 B.n87 10.6151
R763 B.n303 B.n302 10.6151
R764 B.n304 B.n303 10.6151
R765 B.n304 B.n85 10.6151
R766 B.n308 B.n85 10.6151
R767 B.n309 B.n308 10.6151
R768 B.n310 B.n309 10.6151
R769 B.n310 B.n83 10.6151
R770 B.n314 B.n83 10.6151
R771 B.n315 B.n314 10.6151
R772 B.n316 B.n315 10.6151
R773 B.n316 B.n81 10.6151
R774 B.n320 B.n81 10.6151
R775 B.n321 B.n320 10.6151
R776 B.n322 B.n321 10.6151
R777 B.n322 B.n79 10.6151
R778 B.n326 B.n79 10.6151
R779 B.n327 B.n326 10.6151
R780 B.n328 B.n327 10.6151
R781 B.n328 B.n77 10.6151
R782 B.n332 B.n77 10.6151
R783 B.n333 B.n332 10.6151
R784 B.n334 B.n333 10.6151
R785 B.n334 B.n75 10.6151
R786 B.n338 B.n75 10.6151
R787 B.n339 B.n338 10.6151
R788 B.n340 B.n339 10.6151
R789 B.n340 B.n73 10.6151
R790 B.n344 B.n73 10.6151
R791 B.n345 B.n344 10.6151
R792 B.n346 B.n345 10.6151
R793 B.n346 B.n71 10.6151
R794 B.n350 B.n71 10.6151
R795 B.n351 B.n350 10.6151
R796 B.n352 B.n351 10.6151
R797 B.n352 B.n69 10.6151
R798 B.n356 B.n69 10.6151
R799 B.n357 B.n356 10.6151
R800 B.n358 B.n357 10.6151
R801 B.n358 B.n67 10.6151
R802 B.n362 B.n67 10.6151
R803 B.n363 B.n362 10.6151
R804 B.n364 B.n363 10.6151
R805 B.n364 B.n65 10.6151
R806 B.n368 B.n65 10.6151
R807 B.n369 B.n368 10.6151
R808 B.n370 B.n369 10.6151
R809 B.n370 B.n63 10.6151
R810 B.n374 B.n63 10.6151
R811 B.n375 B.n374 10.6151
R812 B.n376 B.n375 10.6151
R813 B.n376 B.n61 10.6151
R814 B.n380 B.n61 10.6151
R815 B.n381 B.n380 10.6151
R816 B.n382 B.n381 10.6151
R817 B.n382 B.n59 10.6151
R818 B.n386 B.n59 10.6151
R819 B.n387 B.n386 10.6151
R820 B.n388 B.n387 10.6151
R821 B.n388 B.n57 10.6151
R822 B.n392 B.n57 10.6151
R823 B.n393 B.n392 10.6151
R824 B.n195 B.n194 10.6151
R825 B.n196 B.n195 10.6151
R826 B.n196 B.n125 10.6151
R827 B.n200 B.n125 10.6151
R828 B.n201 B.n200 10.6151
R829 B.n202 B.n201 10.6151
R830 B.n202 B.n123 10.6151
R831 B.n206 B.n123 10.6151
R832 B.n207 B.n206 10.6151
R833 B.n208 B.n207 10.6151
R834 B.n208 B.n121 10.6151
R835 B.n212 B.n121 10.6151
R836 B.n213 B.n212 10.6151
R837 B.n214 B.n213 10.6151
R838 B.n214 B.n119 10.6151
R839 B.n218 B.n119 10.6151
R840 B.n219 B.n218 10.6151
R841 B.n220 B.n219 10.6151
R842 B.n220 B.n117 10.6151
R843 B.n224 B.n117 10.6151
R844 B.n225 B.n224 10.6151
R845 B.n226 B.n225 10.6151
R846 B.n226 B.n115 10.6151
R847 B.n230 B.n115 10.6151
R848 B.n231 B.n230 10.6151
R849 B.n232 B.n231 10.6151
R850 B.n236 B.n235 10.6151
R851 B.n237 B.n236 10.6151
R852 B.n237 B.n109 10.6151
R853 B.n241 B.n109 10.6151
R854 B.n242 B.n241 10.6151
R855 B.n243 B.n242 10.6151
R856 B.n243 B.n107 10.6151
R857 B.n247 B.n107 10.6151
R858 B.n248 B.n247 10.6151
R859 B.n250 B.n103 10.6151
R860 B.n254 B.n103 10.6151
R861 B.n255 B.n254 10.6151
R862 B.n256 B.n255 10.6151
R863 B.n256 B.n101 10.6151
R864 B.n260 B.n101 10.6151
R865 B.n261 B.n260 10.6151
R866 B.n262 B.n261 10.6151
R867 B.n262 B.n99 10.6151
R868 B.n266 B.n99 10.6151
R869 B.n267 B.n266 10.6151
R870 B.n268 B.n267 10.6151
R871 B.n268 B.n97 10.6151
R872 B.n272 B.n97 10.6151
R873 B.n273 B.n272 10.6151
R874 B.n274 B.n273 10.6151
R875 B.n274 B.n95 10.6151
R876 B.n278 B.n95 10.6151
R877 B.n279 B.n278 10.6151
R878 B.n280 B.n279 10.6151
R879 B.n280 B.n93 10.6151
R880 B.n284 B.n93 10.6151
R881 B.n285 B.n284 10.6151
R882 B.n286 B.n285 10.6151
R883 B.n286 B.n91 10.6151
R884 B.n290 B.n91 10.6151
R885 B.n190 B.n127 10.6151
R886 B.n190 B.n189 10.6151
R887 B.n189 B.n188 10.6151
R888 B.n188 B.n129 10.6151
R889 B.n184 B.n129 10.6151
R890 B.n184 B.n183 10.6151
R891 B.n183 B.n182 10.6151
R892 B.n182 B.n131 10.6151
R893 B.n178 B.n131 10.6151
R894 B.n178 B.n177 10.6151
R895 B.n177 B.n176 10.6151
R896 B.n176 B.n133 10.6151
R897 B.n172 B.n133 10.6151
R898 B.n172 B.n171 10.6151
R899 B.n171 B.n170 10.6151
R900 B.n170 B.n135 10.6151
R901 B.n166 B.n135 10.6151
R902 B.n166 B.n165 10.6151
R903 B.n165 B.n164 10.6151
R904 B.n164 B.n137 10.6151
R905 B.n160 B.n137 10.6151
R906 B.n160 B.n159 10.6151
R907 B.n159 B.n158 10.6151
R908 B.n158 B.n139 10.6151
R909 B.n154 B.n139 10.6151
R910 B.n154 B.n153 10.6151
R911 B.n153 B.n152 10.6151
R912 B.n152 B.n141 10.6151
R913 B.n148 B.n141 10.6151
R914 B.n148 B.n147 10.6151
R915 B.n147 B.n146 10.6151
R916 B.n146 B.n143 10.6151
R917 B.n143 B.n0 10.6151
R918 B.n539 B.n1 10.6151
R919 B.n539 B.n538 10.6151
R920 B.n538 B.n537 10.6151
R921 B.n537 B.n4 10.6151
R922 B.n533 B.n4 10.6151
R923 B.n533 B.n532 10.6151
R924 B.n532 B.n531 10.6151
R925 B.n531 B.n6 10.6151
R926 B.n527 B.n6 10.6151
R927 B.n527 B.n526 10.6151
R928 B.n526 B.n525 10.6151
R929 B.n525 B.n8 10.6151
R930 B.n521 B.n8 10.6151
R931 B.n521 B.n520 10.6151
R932 B.n520 B.n519 10.6151
R933 B.n519 B.n10 10.6151
R934 B.n515 B.n10 10.6151
R935 B.n515 B.n514 10.6151
R936 B.n514 B.n513 10.6151
R937 B.n513 B.n12 10.6151
R938 B.n509 B.n12 10.6151
R939 B.n509 B.n508 10.6151
R940 B.n508 B.n507 10.6151
R941 B.n507 B.n14 10.6151
R942 B.n503 B.n14 10.6151
R943 B.n503 B.n502 10.6151
R944 B.n502 B.n501 10.6151
R945 B.n501 B.n16 10.6151
R946 B.n497 B.n16 10.6151
R947 B.n497 B.n496 10.6151
R948 B.n496 B.n495 10.6151
R949 B.n495 B.n18 10.6151
R950 B.n491 B.n18 10.6151
R951 B.n36 B.n32 9.36635
R952 B.n435 B.n434 9.36635
R953 B.n232 B.n113 9.36635
R954 B.n250 B.n249 9.36635
R955 B.n543 B.n0 2.81026
R956 B.n543 B.n1 2.81026
R957 B.n449 B.n36 1.24928
R958 B.n436 B.n435 1.24928
R959 B.n235 B.n113 1.24928
R960 B.n249 B.n248 1.24928
C0 VN VDD2 3.82221f
C1 VTAIL B 2.32854f
C2 VDD1 B 1.51667f
C3 VTAIL w_n2738_n2376# 2.21331f
C4 VDD1 w_n2738_n2376# 1.76637f
C5 VTAIL VP 4.14356f
C6 VDD1 VP 4.06693f
C7 VTAIL VDD2 5.75935f
C8 VDD1 VDD2 1.15054f
C9 VN VTAIL 4.1293f
C10 VDD1 VN 0.150115f
C11 VDD1 VTAIL 5.71277f
C12 w_n2738_n2376# B 7.2929f
C13 VP B 1.54351f
C14 VP w_n2738_n2376# 5.26925f
C15 B VDD2 1.57351f
C16 VN B 0.95947f
C17 w_n2738_n2376# VDD2 1.82848f
C18 VP VDD2 0.397201f
C19 VN w_n2738_n2376# 4.91728f
C20 VN VP 5.30615f
C21 VDD2 VSUBS 1.319237f
C22 VDD1 VSUBS 1.726332f
C23 VTAIL VSUBS 0.639446f
C24 VN VSUBS 4.88906f
C25 VP VSUBS 2.08713f
C26 B VSUBS 3.505297f
C27 w_n2738_n2376# VSUBS 80.92429f
C28 B.n0 VSUBS 0.00478f
C29 B.n1 VSUBS 0.00478f
C30 B.n2 VSUBS 0.007559f
C31 B.n3 VSUBS 0.007559f
C32 B.n4 VSUBS 0.007559f
C33 B.n5 VSUBS 0.007559f
C34 B.n6 VSUBS 0.007559f
C35 B.n7 VSUBS 0.007559f
C36 B.n8 VSUBS 0.007559f
C37 B.n9 VSUBS 0.007559f
C38 B.n10 VSUBS 0.007559f
C39 B.n11 VSUBS 0.007559f
C40 B.n12 VSUBS 0.007559f
C41 B.n13 VSUBS 0.007559f
C42 B.n14 VSUBS 0.007559f
C43 B.n15 VSUBS 0.007559f
C44 B.n16 VSUBS 0.007559f
C45 B.n17 VSUBS 0.007559f
C46 B.n18 VSUBS 0.007559f
C47 B.n19 VSUBS 0.018003f
C48 B.n20 VSUBS 0.007559f
C49 B.n21 VSUBS 0.007559f
C50 B.n22 VSUBS 0.007559f
C51 B.n23 VSUBS 0.007559f
C52 B.n24 VSUBS 0.007559f
C53 B.n25 VSUBS 0.007559f
C54 B.n26 VSUBS 0.007559f
C55 B.n27 VSUBS 0.007559f
C56 B.n28 VSUBS 0.007559f
C57 B.n29 VSUBS 0.007559f
C58 B.n30 VSUBS 0.007559f
C59 B.n31 VSUBS 0.007559f
C60 B.n32 VSUBS 0.007114f
C61 B.n33 VSUBS 0.007559f
C62 B.t2 VSUBS 0.229211f
C63 B.t1 VSUBS 0.246385f
C64 B.t0 VSUBS 0.658088f
C65 B.n34 VSUBS 0.131022f
C66 B.n35 VSUBS 0.07373f
C67 B.n36 VSUBS 0.017513f
C68 B.n37 VSUBS 0.007559f
C69 B.n38 VSUBS 0.007559f
C70 B.n39 VSUBS 0.007559f
C71 B.n40 VSUBS 0.007559f
C72 B.t11 VSUBS 0.22921f
C73 B.t10 VSUBS 0.246384f
C74 B.t9 VSUBS 0.658088f
C75 B.n41 VSUBS 0.131024f
C76 B.n42 VSUBS 0.073731f
C77 B.n43 VSUBS 0.007559f
C78 B.n44 VSUBS 0.007559f
C79 B.n45 VSUBS 0.007559f
C80 B.n46 VSUBS 0.007559f
C81 B.n47 VSUBS 0.007559f
C82 B.n48 VSUBS 0.007559f
C83 B.n49 VSUBS 0.007559f
C84 B.n50 VSUBS 0.007559f
C85 B.n51 VSUBS 0.007559f
C86 B.n52 VSUBS 0.007559f
C87 B.n53 VSUBS 0.007559f
C88 B.n54 VSUBS 0.007559f
C89 B.n55 VSUBS 0.007559f
C90 B.n56 VSUBS 0.016678f
C91 B.n57 VSUBS 0.007559f
C92 B.n58 VSUBS 0.007559f
C93 B.n59 VSUBS 0.007559f
C94 B.n60 VSUBS 0.007559f
C95 B.n61 VSUBS 0.007559f
C96 B.n62 VSUBS 0.007559f
C97 B.n63 VSUBS 0.007559f
C98 B.n64 VSUBS 0.007559f
C99 B.n65 VSUBS 0.007559f
C100 B.n66 VSUBS 0.007559f
C101 B.n67 VSUBS 0.007559f
C102 B.n68 VSUBS 0.007559f
C103 B.n69 VSUBS 0.007559f
C104 B.n70 VSUBS 0.007559f
C105 B.n71 VSUBS 0.007559f
C106 B.n72 VSUBS 0.007559f
C107 B.n73 VSUBS 0.007559f
C108 B.n74 VSUBS 0.007559f
C109 B.n75 VSUBS 0.007559f
C110 B.n76 VSUBS 0.007559f
C111 B.n77 VSUBS 0.007559f
C112 B.n78 VSUBS 0.007559f
C113 B.n79 VSUBS 0.007559f
C114 B.n80 VSUBS 0.007559f
C115 B.n81 VSUBS 0.007559f
C116 B.n82 VSUBS 0.007559f
C117 B.n83 VSUBS 0.007559f
C118 B.n84 VSUBS 0.007559f
C119 B.n85 VSUBS 0.007559f
C120 B.n86 VSUBS 0.007559f
C121 B.n87 VSUBS 0.007559f
C122 B.n88 VSUBS 0.007559f
C123 B.n89 VSUBS 0.007559f
C124 B.n90 VSUBS 0.016678f
C125 B.n91 VSUBS 0.007559f
C126 B.n92 VSUBS 0.007559f
C127 B.n93 VSUBS 0.007559f
C128 B.n94 VSUBS 0.007559f
C129 B.n95 VSUBS 0.007559f
C130 B.n96 VSUBS 0.007559f
C131 B.n97 VSUBS 0.007559f
C132 B.n98 VSUBS 0.007559f
C133 B.n99 VSUBS 0.007559f
C134 B.n100 VSUBS 0.007559f
C135 B.n101 VSUBS 0.007559f
C136 B.n102 VSUBS 0.007559f
C137 B.n103 VSUBS 0.007559f
C138 B.n104 VSUBS 0.007559f
C139 B.t4 VSUBS 0.22921f
C140 B.t5 VSUBS 0.246384f
C141 B.t3 VSUBS 0.658088f
C142 B.n105 VSUBS 0.131024f
C143 B.n106 VSUBS 0.073731f
C144 B.n107 VSUBS 0.007559f
C145 B.n108 VSUBS 0.007559f
C146 B.n109 VSUBS 0.007559f
C147 B.n110 VSUBS 0.007559f
C148 B.t7 VSUBS 0.229211f
C149 B.t8 VSUBS 0.246385f
C150 B.t6 VSUBS 0.658088f
C151 B.n111 VSUBS 0.131022f
C152 B.n112 VSUBS 0.07373f
C153 B.n113 VSUBS 0.017513f
C154 B.n114 VSUBS 0.007559f
C155 B.n115 VSUBS 0.007559f
C156 B.n116 VSUBS 0.007559f
C157 B.n117 VSUBS 0.007559f
C158 B.n118 VSUBS 0.007559f
C159 B.n119 VSUBS 0.007559f
C160 B.n120 VSUBS 0.007559f
C161 B.n121 VSUBS 0.007559f
C162 B.n122 VSUBS 0.007559f
C163 B.n123 VSUBS 0.007559f
C164 B.n124 VSUBS 0.007559f
C165 B.n125 VSUBS 0.007559f
C166 B.n126 VSUBS 0.007559f
C167 B.n127 VSUBS 0.016678f
C168 B.n128 VSUBS 0.007559f
C169 B.n129 VSUBS 0.007559f
C170 B.n130 VSUBS 0.007559f
C171 B.n131 VSUBS 0.007559f
C172 B.n132 VSUBS 0.007559f
C173 B.n133 VSUBS 0.007559f
C174 B.n134 VSUBS 0.007559f
C175 B.n135 VSUBS 0.007559f
C176 B.n136 VSUBS 0.007559f
C177 B.n137 VSUBS 0.007559f
C178 B.n138 VSUBS 0.007559f
C179 B.n139 VSUBS 0.007559f
C180 B.n140 VSUBS 0.007559f
C181 B.n141 VSUBS 0.007559f
C182 B.n142 VSUBS 0.007559f
C183 B.n143 VSUBS 0.007559f
C184 B.n144 VSUBS 0.007559f
C185 B.n145 VSUBS 0.007559f
C186 B.n146 VSUBS 0.007559f
C187 B.n147 VSUBS 0.007559f
C188 B.n148 VSUBS 0.007559f
C189 B.n149 VSUBS 0.007559f
C190 B.n150 VSUBS 0.007559f
C191 B.n151 VSUBS 0.007559f
C192 B.n152 VSUBS 0.007559f
C193 B.n153 VSUBS 0.007559f
C194 B.n154 VSUBS 0.007559f
C195 B.n155 VSUBS 0.007559f
C196 B.n156 VSUBS 0.007559f
C197 B.n157 VSUBS 0.007559f
C198 B.n158 VSUBS 0.007559f
C199 B.n159 VSUBS 0.007559f
C200 B.n160 VSUBS 0.007559f
C201 B.n161 VSUBS 0.007559f
C202 B.n162 VSUBS 0.007559f
C203 B.n163 VSUBS 0.007559f
C204 B.n164 VSUBS 0.007559f
C205 B.n165 VSUBS 0.007559f
C206 B.n166 VSUBS 0.007559f
C207 B.n167 VSUBS 0.007559f
C208 B.n168 VSUBS 0.007559f
C209 B.n169 VSUBS 0.007559f
C210 B.n170 VSUBS 0.007559f
C211 B.n171 VSUBS 0.007559f
C212 B.n172 VSUBS 0.007559f
C213 B.n173 VSUBS 0.007559f
C214 B.n174 VSUBS 0.007559f
C215 B.n175 VSUBS 0.007559f
C216 B.n176 VSUBS 0.007559f
C217 B.n177 VSUBS 0.007559f
C218 B.n178 VSUBS 0.007559f
C219 B.n179 VSUBS 0.007559f
C220 B.n180 VSUBS 0.007559f
C221 B.n181 VSUBS 0.007559f
C222 B.n182 VSUBS 0.007559f
C223 B.n183 VSUBS 0.007559f
C224 B.n184 VSUBS 0.007559f
C225 B.n185 VSUBS 0.007559f
C226 B.n186 VSUBS 0.007559f
C227 B.n187 VSUBS 0.007559f
C228 B.n188 VSUBS 0.007559f
C229 B.n189 VSUBS 0.007559f
C230 B.n190 VSUBS 0.007559f
C231 B.n191 VSUBS 0.007559f
C232 B.n192 VSUBS 0.016678f
C233 B.n193 VSUBS 0.018003f
C234 B.n194 VSUBS 0.018003f
C235 B.n195 VSUBS 0.007559f
C236 B.n196 VSUBS 0.007559f
C237 B.n197 VSUBS 0.007559f
C238 B.n198 VSUBS 0.007559f
C239 B.n199 VSUBS 0.007559f
C240 B.n200 VSUBS 0.007559f
C241 B.n201 VSUBS 0.007559f
C242 B.n202 VSUBS 0.007559f
C243 B.n203 VSUBS 0.007559f
C244 B.n204 VSUBS 0.007559f
C245 B.n205 VSUBS 0.007559f
C246 B.n206 VSUBS 0.007559f
C247 B.n207 VSUBS 0.007559f
C248 B.n208 VSUBS 0.007559f
C249 B.n209 VSUBS 0.007559f
C250 B.n210 VSUBS 0.007559f
C251 B.n211 VSUBS 0.007559f
C252 B.n212 VSUBS 0.007559f
C253 B.n213 VSUBS 0.007559f
C254 B.n214 VSUBS 0.007559f
C255 B.n215 VSUBS 0.007559f
C256 B.n216 VSUBS 0.007559f
C257 B.n217 VSUBS 0.007559f
C258 B.n218 VSUBS 0.007559f
C259 B.n219 VSUBS 0.007559f
C260 B.n220 VSUBS 0.007559f
C261 B.n221 VSUBS 0.007559f
C262 B.n222 VSUBS 0.007559f
C263 B.n223 VSUBS 0.007559f
C264 B.n224 VSUBS 0.007559f
C265 B.n225 VSUBS 0.007559f
C266 B.n226 VSUBS 0.007559f
C267 B.n227 VSUBS 0.007559f
C268 B.n228 VSUBS 0.007559f
C269 B.n229 VSUBS 0.007559f
C270 B.n230 VSUBS 0.007559f
C271 B.n231 VSUBS 0.007559f
C272 B.n232 VSUBS 0.007114f
C273 B.n233 VSUBS 0.007559f
C274 B.n234 VSUBS 0.007559f
C275 B.n235 VSUBS 0.004224f
C276 B.n236 VSUBS 0.007559f
C277 B.n237 VSUBS 0.007559f
C278 B.n238 VSUBS 0.007559f
C279 B.n239 VSUBS 0.007559f
C280 B.n240 VSUBS 0.007559f
C281 B.n241 VSUBS 0.007559f
C282 B.n242 VSUBS 0.007559f
C283 B.n243 VSUBS 0.007559f
C284 B.n244 VSUBS 0.007559f
C285 B.n245 VSUBS 0.007559f
C286 B.n246 VSUBS 0.007559f
C287 B.n247 VSUBS 0.007559f
C288 B.n248 VSUBS 0.004224f
C289 B.n249 VSUBS 0.017513f
C290 B.n250 VSUBS 0.007114f
C291 B.n251 VSUBS 0.007559f
C292 B.n252 VSUBS 0.007559f
C293 B.n253 VSUBS 0.007559f
C294 B.n254 VSUBS 0.007559f
C295 B.n255 VSUBS 0.007559f
C296 B.n256 VSUBS 0.007559f
C297 B.n257 VSUBS 0.007559f
C298 B.n258 VSUBS 0.007559f
C299 B.n259 VSUBS 0.007559f
C300 B.n260 VSUBS 0.007559f
C301 B.n261 VSUBS 0.007559f
C302 B.n262 VSUBS 0.007559f
C303 B.n263 VSUBS 0.007559f
C304 B.n264 VSUBS 0.007559f
C305 B.n265 VSUBS 0.007559f
C306 B.n266 VSUBS 0.007559f
C307 B.n267 VSUBS 0.007559f
C308 B.n268 VSUBS 0.007559f
C309 B.n269 VSUBS 0.007559f
C310 B.n270 VSUBS 0.007559f
C311 B.n271 VSUBS 0.007559f
C312 B.n272 VSUBS 0.007559f
C313 B.n273 VSUBS 0.007559f
C314 B.n274 VSUBS 0.007559f
C315 B.n275 VSUBS 0.007559f
C316 B.n276 VSUBS 0.007559f
C317 B.n277 VSUBS 0.007559f
C318 B.n278 VSUBS 0.007559f
C319 B.n279 VSUBS 0.007559f
C320 B.n280 VSUBS 0.007559f
C321 B.n281 VSUBS 0.007559f
C322 B.n282 VSUBS 0.007559f
C323 B.n283 VSUBS 0.007559f
C324 B.n284 VSUBS 0.007559f
C325 B.n285 VSUBS 0.007559f
C326 B.n286 VSUBS 0.007559f
C327 B.n287 VSUBS 0.007559f
C328 B.n288 VSUBS 0.007559f
C329 B.n289 VSUBS 0.018003f
C330 B.n290 VSUBS 0.018003f
C331 B.n291 VSUBS 0.016678f
C332 B.n292 VSUBS 0.007559f
C333 B.n293 VSUBS 0.007559f
C334 B.n294 VSUBS 0.007559f
C335 B.n295 VSUBS 0.007559f
C336 B.n296 VSUBS 0.007559f
C337 B.n297 VSUBS 0.007559f
C338 B.n298 VSUBS 0.007559f
C339 B.n299 VSUBS 0.007559f
C340 B.n300 VSUBS 0.007559f
C341 B.n301 VSUBS 0.007559f
C342 B.n302 VSUBS 0.007559f
C343 B.n303 VSUBS 0.007559f
C344 B.n304 VSUBS 0.007559f
C345 B.n305 VSUBS 0.007559f
C346 B.n306 VSUBS 0.007559f
C347 B.n307 VSUBS 0.007559f
C348 B.n308 VSUBS 0.007559f
C349 B.n309 VSUBS 0.007559f
C350 B.n310 VSUBS 0.007559f
C351 B.n311 VSUBS 0.007559f
C352 B.n312 VSUBS 0.007559f
C353 B.n313 VSUBS 0.007559f
C354 B.n314 VSUBS 0.007559f
C355 B.n315 VSUBS 0.007559f
C356 B.n316 VSUBS 0.007559f
C357 B.n317 VSUBS 0.007559f
C358 B.n318 VSUBS 0.007559f
C359 B.n319 VSUBS 0.007559f
C360 B.n320 VSUBS 0.007559f
C361 B.n321 VSUBS 0.007559f
C362 B.n322 VSUBS 0.007559f
C363 B.n323 VSUBS 0.007559f
C364 B.n324 VSUBS 0.007559f
C365 B.n325 VSUBS 0.007559f
C366 B.n326 VSUBS 0.007559f
C367 B.n327 VSUBS 0.007559f
C368 B.n328 VSUBS 0.007559f
C369 B.n329 VSUBS 0.007559f
C370 B.n330 VSUBS 0.007559f
C371 B.n331 VSUBS 0.007559f
C372 B.n332 VSUBS 0.007559f
C373 B.n333 VSUBS 0.007559f
C374 B.n334 VSUBS 0.007559f
C375 B.n335 VSUBS 0.007559f
C376 B.n336 VSUBS 0.007559f
C377 B.n337 VSUBS 0.007559f
C378 B.n338 VSUBS 0.007559f
C379 B.n339 VSUBS 0.007559f
C380 B.n340 VSUBS 0.007559f
C381 B.n341 VSUBS 0.007559f
C382 B.n342 VSUBS 0.007559f
C383 B.n343 VSUBS 0.007559f
C384 B.n344 VSUBS 0.007559f
C385 B.n345 VSUBS 0.007559f
C386 B.n346 VSUBS 0.007559f
C387 B.n347 VSUBS 0.007559f
C388 B.n348 VSUBS 0.007559f
C389 B.n349 VSUBS 0.007559f
C390 B.n350 VSUBS 0.007559f
C391 B.n351 VSUBS 0.007559f
C392 B.n352 VSUBS 0.007559f
C393 B.n353 VSUBS 0.007559f
C394 B.n354 VSUBS 0.007559f
C395 B.n355 VSUBS 0.007559f
C396 B.n356 VSUBS 0.007559f
C397 B.n357 VSUBS 0.007559f
C398 B.n358 VSUBS 0.007559f
C399 B.n359 VSUBS 0.007559f
C400 B.n360 VSUBS 0.007559f
C401 B.n361 VSUBS 0.007559f
C402 B.n362 VSUBS 0.007559f
C403 B.n363 VSUBS 0.007559f
C404 B.n364 VSUBS 0.007559f
C405 B.n365 VSUBS 0.007559f
C406 B.n366 VSUBS 0.007559f
C407 B.n367 VSUBS 0.007559f
C408 B.n368 VSUBS 0.007559f
C409 B.n369 VSUBS 0.007559f
C410 B.n370 VSUBS 0.007559f
C411 B.n371 VSUBS 0.007559f
C412 B.n372 VSUBS 0.007559f
C413 B.n373 VSUBS 0.007559f
C414 B.n374 VSUBS 0.007559f
C415 B.n375 VSUBS 0.007559f
C416 B.n376 VSUBS 0.007559f
C417 B.n377 VSUBS 0.007559f
C418 B.n378 VSUBS 0.007559f
C419 B.n379 VSUBS 0.007559f
C420 B.n380 VSUBS 0.007559f
C421 B.n381 VSUBS 0.007559f
C422 B.n382 VSUBS 0.007559f
C423 B.n383 VSUBS 0.007559f
C424 B.n384 VSUBS 0.007559f
C425 B.n385 VSUBS 0.007559f
C426 B.n386 VSUBS 0.007559f
C427 B.n387 VSUBS 0.007559f
C428 B.n388 VSUBS 0.007559f
C429 B.n389 VSUBS 0.007559f
C430 B.n390 VSUBS 0.007559f
C431 B.n391 VSUBS 0.007559f
C432 B.n392 VSUBS 0.007559f
C433 B.n393 VSUBS 0.017599f
C434 B.n394 VSUBS 0.017083f
C435 B.n395 VSUBS 0.018003f
C436 B.n396 VSUBS 0.007559f
C437 B.n397 VSUBS 0.007559f
C438 B.n398 VSUBS 0.007559f
C439 B.n399 VSUBS 0.007559f
C440 B.n400 VSUBS 0.007559f
C441 B.n401 VSUBS 0.007559f
C442 B.n402 VSUBS 0.007559f
C443 B.n403 VSUBS 0.007559f
C444 B.n404 VSUBS 0.007559f
C445 B.n405 VSUBS 0.007559f
C446 B.n406 VSUBS 0.007559f
C447 B.n407 VSUBS 0.007559f
C448 B.n408 VSUBS 0.007559f
C449 B.n409 VSUBS 0.007559f
C450 B.n410 VSUBS 0.007559f
C451 B.n411 VSUBS 0.007559f
C452 B.n412 VSUBS 0.007559f
C453 B.n413 VSUBS 0.007559f
C454 B.n414 VSUBS 0.007559f
C455 B.n415 VSUBS 0.007559f
C456 B.n416 VSUBS 0.007559f
C457 B.n417 VSUBS 0.007559f
C458 B.n418 VSUBS 0.007559f
C459 B.n419 VSUBS 0.007559f
C460 B.n420 VSUBS 0.007559f
C461 B.n421 VSUBS 0.007559f
C462 B.n422 VSUBS 0.007559f
C463 B.n423 VSUBS 0.007559f
C464 B.n424 VSUBS 0.007559f
C465 B.n425 VSUBS 0.007559f
C466 B.n426 VSUBS 0.007559f
C467 B.n427 VSUBS 0.007559f
C468 B.n428 VSUBS 0.007559f
C469 B.n429 VSUBS 0.007559f
C470 B.n430 VSUBS 0.007559f
C471 B.n431 VSUBS 0.007559f
C472 B.n432 VSUBS 0.007559f
C473 B.n433 VSUBS 0.007559f
C474 B.n434 VSUBS 0.007114f
C475 B.n435 VSUBS 0.017513f
C476 B.n436 VSUBS 0.004224f
C477 B.n437 VSUBS 0.007559f
C478 B.n438 VSUBS 0.007559f
C479 B.n439 VSUBS 0.007559f
C480 B.n440 VSUBS 0.007559f
C481 B.n441 VSUBS 0.007559f
C482 B.n442 VSUBS 0.007559f
C483 B.n443 VSUBS 0.007559f
C484 B.n444 VSUBS 0.007559f
C485 B.n445 VSUBS 0.007559f
C486 B.n446 VSUBS 0.007559f
C487 B.n447 VSUBS 0.007559f
C488 B.n448 VSUBS 0.007559f
C489 B.n449 VSUBS 0.004224f
C490 B.n450 VSUBS 0.007559f
C491 B.n451 VSUBS 0.007559f
C492 B.n452 VSUBS 0.007559f
C493 B.n453 VSUBS 0.007559f
C494 B.n454 VSUBS 0.007559f
C495 B.n455 VSUBS 0.007559f
C496 B.n456 VSUBS 0.007559f
C497 B.n457 VSUBS 0.007559f
C498 B.n458 VSUBS 0.007559f
C499 B.n459 VSUBS 0.007559f
C500 B.n460 VSUBS 0.007559f
C501 B.n461 VSUBS 0.007559f
C502 B.n462 VSUBS 0.007559f
C503 B.n463 VSUBS 0.007559f
C504 B.n464 VSUBS 0.007559f
C505 B.n465 VSUBS 0.007559f
C506 B.n466 VSUBS 0.007559f
C507 B.n467 VSUBS 0.007559f
C508 B.n468 VSUBS 0.007559f
C509 B.n469 VSUBS 0.007559f
C510 B.n470 VSUBS 0.007559f
C511 B.n471 VSUBS 0.007559f
C512 B.n472 VSUBS 0.007559f
C513 B.n473 VSUBS 0.007559f
C514 B.n474 VSUBS 0.007559f
C515 B.n475 VSUBS 0.007559f
C516 B.n476 VSUBS 0.007559f
C517 B.n477 VSUBS 0.007559f
C518 B.n478 VSUBS 0.007559f
C519 B.n479 VSUBS 0.007559f
C520 B.n480 VSUBS 0.007559f
C521 B.n481 VSUBS 0.007559f
C522 B.n482 VSUBS 0.007559f
C523 B.n483 VSUBS 0.007559f
C524 B.n484 VSUBS 0.007559f
C525 B.n485 VSUBS 0.007559f
C526 B.n486 VSUBS 0.007559f
C527 B.n487 VSUBS 0.007559f
C528 B.n488 VSUBS 0.007559f
C529 B.n489 VSUBS 0.007559f
C530 B.n490 VSUBS 0.018003f
C531 B.n491 VSUBS 0.016678f
C532 B.n492 VSUBS 0.016678f
C533 B.n493 VSUBS 0.007559f
C534 B.n494 VSUBS 0.007559f
C535 B.n495 VSUBS 0.007559f
C536 B.n496 VSUBS 0.007559f
C537 B.n497 VSUBS 0.007559f
C538 B.n498 VSUBS 0.007559f
C539 B.n499 VSUBS 0.007559f
C540 B.n500 VSUBS 0.007559f
C541 B.n501 VSUBS 0.007559f
C542 B.n502 VSUBS 0.007559f
C543 B.n503 VSUBS 0.007559f
C544 B.n504 VSUBS 0.007559f
C545 B.n505 VSUBS 0.007559f
C546 B.n506 VSUBS 0.007559f
C547 B.n507 VSUBS 0.007559f
C548 B.n508 VSUBS 0.007559f
C549 B.n509 VSUBS 0.007559f
C550 B.n510 VSUBS 0.007559f
C551 B.n511 VSUBS 0.007559f
C552 B.n512 VSUBS 0.007559f
C553 B.n513 VSUBS 0.007559f
C554 B.n514 VSUBS 0.007559f
C555 B.n515 VSUBS 0.007559f
C556 B.n516 VSUBS 0.007559f
C557 B.n517 VSUBS 0.007559f
C558 B.n518 VSUBS 0.007559f
C559 B.n519 VSUBS 0.007559f
C560 B.n520 VSUBS 0.007559f
C561 B.n521 VSUBS 0.007559f
C562 B.n522 VSUBS 0.007559f
C563 B.n523 VSUBS 0.007559f
C564 B.n524 VSUBS 0.007559f
C565 B.n525 VSUBS 0.007559f
C566 B.n526 VSUBS 0.007559f
C567 B.n527 VSUBS 0.007559f
C568 B.n528 VSUBS 0.007559f
C569 B.n529 VSUBS 0.007559f
C570 B.n530 VSUBS 0.007559f
C571 B.n531 VSUBS 0.007559f
C572 B.n532 VSUBS 0.007559f
C573 B.n533 VSUBS 0.007559f
C574 B.n534 VSUBS 0.007559f
C575 B.n535 VSUBS 0.007559f
C576 B.n536 VSUBS 0.007559f
C577 B.n537 VSUBS 0.007559f
C578 B.n538 VSUBS 0.007559f
C579 B.n539 VSUBS 0.007559f
C580 B.n540 VSUBS 0.007559f
C581 B.n541 VSUBS 0.007559f
C582 B.n542 VSUBS 0.007559f
C583 B.n543 VSUBS 0.017116f
C584 VDD1.t0 VSUBS 1.13987f
C585 VDD1.t1 VSUBS 1.13909f
C586 VDD1.t2 VSUBS 0.123087f
C587 VDD1.t3 VSUBS 0.123087f
C588 VDD1.n0 VSUBS 0.852162f
C589 VDD1.n1 VSUBS 2.50921f
C590 VDD1.t5 VSUBS 0.123087f
C591 VDD1.t4 VSUBS 0.123087f
C592 VDD1.n2 VSUBS 0.849461f
C593 VDD1.n3 VSUBS 2.1438f
C594 VP.n0 VSUBS 0.056945f
C595 VP.t2 VSUBS 1.52629f
C596 VP.n1 VSUBS 0.074883f
C597 VP.n2 VSUBS 0.043195f
C598 VP.t3 VSUBS 1.52629f
C599 VP.n3 VSUBS 0.048041f
C600 VP.n4 VSUBS 0.056945f
C601 VP.t1 VSUBS 1.52629f
C602 VP.n5 VSUBS 0.074883f
C603 VP.t5 VSUBS 1.72545f
C604 VP.n6 VSUBS 0.677971f
C605 VP.t0 VSUBS 1.52629f
C606 VP.n7 VSUBS 0.672085f
C607 VP.n8 VSUBS 0.060329f
C608 VP.n9 VSUBS 0.318729f
C609 VP.n10 VSUBS 0.043195f
C610 VP.n11 VSUBS 0.043195f
C611 VP.n12 VSUBS 0.048041f
C612 VP.n13 VSUBS 0.079594f
C613 VP.n14 VSUBS 0.704425f
C614 VP.n15 VSUBS 1.8241f
C615 VP.n16 VSUBS 1.86106f
C616 VP.t4 VSUBS 1.52629f
C617 VP.n17 VSUBS 0.704425f
C618 VP.n18 VSUBS 0.079594f
C619 VP.n19 VSUBS 0.056945f
C620 VP.n20 VSUBS 0.043195f
C621 VP.n21 VSUBS 0.043195f
C622 VP.n22 VSUBS 0.074883f
C623 VP.n23 VSUBS 0.060329f
C624 VP.n24 VSUBS 0.573595f
C625 VP.n25 VSUBS 0.060329f
C626 VP.n26 VSUBS 0.043195f
C627 VP.n27 VSUBS 0.043195f
C628 VP.n28 VSUBS 0.043195f
C629 VP.n29 VSUBS 0.048041f
C630 VP.n30 VSUBS 0.079594f
C631 VP.n31 VSUBS 0.704425f
C632 VP.n32 VSUBS 0.048207f
C633 VDD2.t4 VSUBS 1.12522f
C634 VDD2.t2 VSUBS 0.121589f
C635 VDD2.t1 VSUBS 0.121589f
C636 VDD2.n0 VSUBS 0.84179f
C637 VDD2.n1 VSUBS 2.38953f
C638 VDD2.t5 VSUBS 1.11727f
C639 VDD2.n2 VSUBS 2.1207f
C640 VDD2.t0 VSUBS 0.121589f
C641 VDD2.t3 VSUBS 0.121589f
C642 VDD2.n3 VSUBS 0.841764f
C643 VTAIL.t6 VSUBS 0.173718f
C644 VTAIL.t9 VSUBS 0.173718f
C645 VTAIL.n0 VSUBS 1.07193f
C646 VTAIL.n1 VSUBS 0.814934f
C647 VTAIL.t3 VSUBS 1.46001f
C648 VTAIL.n2 VSUBS 1.03854f
C649 VTAIL.t2 VSUBS 0.173718f
C650 VTAIL.t0 VSUBS 0.173718f
C651 VTAIL.n3 VSUBS 1.07193f
C652 VTAIL.n4 VSUBS 2.22793f
C653 VTAIL.t7 VSUBS 0.173718f
C654 VTAIL.t11 VSUBS 0.173718f
C655 VTAIL.n5 VSUBS 1.07193f
C656 VTAIL.n6 VSUBS 2.22793f
C657 VTAIL.t10 VSUBS 1.46002f
C658 VTAIL.n7 VSUBS 1.03853f
C659 VTAIL.t4 VSUBS 0.173718f
C660 VTAIL.t5 VSUBS 0.173718f
C661 VTAIL.n8 VSUBS 1.07193f
C662 VTAIL.n9 VSUBS 0.952845f
C663 VTAIL.t1 VSUBS 1.46001f
C664 VTAIL.n10 VSUBS 2.12193f
C665 VTAIL.t8 VSUBS 1.46001f
C666 VTAIL.n11 VSUBS 2.06815f
C667 VN.n0 VSUBS 0.054648f
C668 VN.t4 VSUBS 1.46473f
C669 VN.n1 VSUBS 0.071863f
C670 VN.t1 VSUBS 1.65585f
C671 VN.n2 VSUBS 0.650626f
C672 VN.t3 VSUBS 1.46473f
C673 VN.n3 VSUBS 0.644978f
C674 VN.n4 VSUBS 0.057896f
C675 VN.n5 VSUBS 0.305873f
C676 VN.n6 VSUBS 0.041453f
C677 VN.n7 VSUBS 0.041453f
C678 VN.n8 VSUBS 0.046103f
C679 VN.n9 VSUBS 0.076384f
C680 VN.n10 VSUBS 0.676013f
C681 VN.n11 VSUBS 0.046263f
C682 VN.n12 VSUBS 0.054648f
C683 VN.t0 VSUBS 1.46473f
C684 VN.n13 VSUBS 0.071863f
C685 VN.t2 VSUBS 1.65585f
C686 VN.n14 VSUBS 0.650626f
C687 VN.t5 VSUBS 1.46473f
C688 VN.n15 VSUBS 0.644978f
C689 VN.n16 VSUBS 0.057896f
C690 VN.n17 VSUBS 0.305873f
C691 VN.n18 VSUBS 0.041453f
C692 VN.n19 VSUBS 0.041453f
C693 VN.n20 VSUBS 0.046103f
C694 VN.n21 VSUBS 0.076384f
C695 VN.n22 VSUBS 0.676013f
C696 VN.n23 VSUBS 1.77346f
.ends

