* NGSPICE file created from diff_pair_sample_0861.ext - technology: sky130A

.subckt diff_pair_sample_0861 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X1 VTAIL.t14 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X2 VTAIL.t2 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=1.8018 ps=11.25 w=10.92 l=0.19
X3 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=0 ps=0 w=10.92 l=0.19
X4 VDD1.t6 VP.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=4.2588 ps=22.62 w=10.92 l=0.19
X5 VDD2.t7 VN.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X6 VDD2.t6 VN.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X7 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X8 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=0 ps=0 w=10.92 l=0.19
X9 VDD1.t4 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=0 ps=0 w=10.92 l=0.19
X11 VDD2.t3 VN.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=4.2588 ps=22.62 w=10.92 l=0.19
X12 VDD2.t2 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=4.2588 ps=22.62 w=10.92 l=0.19
X13 VTAIL.t5 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=1.8018 ps=11.25 w=10.92 l=0.19
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=0 ps=0 w=10.92 l=0.19
X15 VDD1.t2 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=4.2588 ps=22.62 w=10.92 l=0.19
X16 VTAIL.t9 VN.t6 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=1.8018 ps=11.25 w=10.92 l=0.19
X17 VTAIL.t8 VN.t7 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2588 pd=22.62 as=1.8018 ps=11.25 w=10.92 l=0.19
X18 VDD1.t1 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8018 pd=11.25 as=1.8018 ps=11.25 w=10.92 l=0.19
R0 VN.n5 VN.t4 1590.91
R1 VN.n1 VN.t7 1590.91
R2 VN.n12 VN.t6 1590.91
R3 VN.n8 VN.t5 1590.91
R4 VN.n4 VN.t1 1550.01
R5 VN.n2 VN.t2 1550.01
R6 VN.n11 VN.t3 1550.01
R7 VN.n9 VN.t0 1550.01
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN VN.n13 39.2221
R15 VN.n3 VN.n2 37.9763
R16 VN.n4 VN.n3 37.9763
R17 VN.n11 VN.n10 37.9763
R18 VN.n10 VN.n9 37.9763
R19 VN.n2 VN.n1 35.055
R20 VN.n5 VN.n4 35.055
R21 VN.n12 VN.n11 35.055
R22 VN.n9 VN.n8 35.055
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VDD2.n2 VDD2.n1 60.0504
R27 VDD2.n2 VDD2.n0 60.0504
R28 VDD2 VDD2.n5 60.0476
R29 VDD2.n4 VDD2.n3 59.8819
R30 VDD2.n4 VDD2.n2 35.1463
R31 VDD2.n5 VDD2.t0 1.81369
R32 VDD2.n5 VDD2.t2 1.81369
R33 VDD2.n3 VDD2.t5 1.81369
R34 VDD2.n3 VDD2.t6 1.81369
R35 VDD2.n1 VDD2.t4 1.81369
R36 VDD2.n1 VDD2.t3 1.81369
R37 VDD2.n0 VDD2.t1 1.81369
R38 VDD2.n0 VDD2.t7 1.81369
R39 VDD2 VDD2.n4 0.282828
R40 VTAIL.n11 VTAIL.t2 45.0162
R41 VTAIL.n10 VTAIL.t10 45.0162
R42 VTAIL.n7 VTAIL.t9 45.0162
R43 VTAIL.n15 VTAIL.t11 45.0161
R44 VTAIL.n2 VTAIL.t8 45.0161
R45 VTAIL.n3 VTAIL.t4 45.0161
R46 VTAIL.n6 VTAIL.t5 45.0161
R47 VTAIL.n14 VTAIL.t6 45.0161
R48 VTAIL.n13 VTAIL.n12 43.2031
R49 VTAIL.n9 VTAIL.n8 43.2031
R50 VTAIL.n1 VTAIL.n0 43.2028
R51 VTAIL.n5 VTAIL.n4 43.2028
R52 VTAIL.n15 VTAIL.n14 22.2289
R53 VTAIL.n7 VTAIL.n6 22.2289
R54 VTAIL.n0 VTAIL.t13 1.81369
R55 VTAIL.n0 VTAIL.t14 1.81369
R56 VTAIL.n4 VTAIL.t7 1.81369
R57 VTAIL.n4 VTAIL.t1 1.81369
R58 VTAIL.n12 VTAIL.t3 1.81369
R59 VTAIL.n12 VTAIL.t0 1.81369
R60 VTAIL.n8 VTAIL.t12 1.81369
R61 VTAIL.n8 VTAIL.t15 1.81369
R62 VTAIL.n11 VTAIL.n10 0.470328
R63 VTAIL.n3 VTAIL.n2 0.470328
R64 VTAIL.n9 VTAIL.n7 0.448776
R65 VTAIL.n10 VTAIL.n9 0.448776
R66 VTAIL.n13 VTAIL.n11 0.448776
R67 VTAIL.n14 VTAIL.n13 0.448776
R68 VTAIL.n6 VTAIL.n5 0.448776
R69 VTAIL.n5 VTAIL.n3 0.448776
R70 VTAIL.n2 VTAIL.n1 0.448776
R71 VTAIL VTAIL.n15 0.390586
R72 VTAIL VTAIL.n1 0.0586897
R73 B.n80 B.t16 1624.64
R74 B.n77 B.t12 1624.64
R75 B.n326 B.t19 1624.64
R76 B.n324 B.t8 1624.64
R77 B.n566 B.n565 585
R78 B.n251 B.n76 585
R79 B.n250 B.n249 585
R80 B.n248 B.n247 585
R81 B.n246 B.n245 585
R82 B.n244 B.n243 585
R83 B.n242 B.n241 585
R84 B.n240 B.n239 585
R85 B.n238 B.n237 585
R86 B.n236 B.n235 585
R87 B.n234 B.n233 585
R88 B.n232 B.n231 585
R89 B.n230 B.n229 585
R90 B.n228 B.n227 585
R91 B.n226 B.n225 585
R92 B.n224 B.n223 585
R93 B.n222 B.n221 585
R94 B.n220 B.n219 585
R95 B.n218 B.n217 585
R96 B.n216 B.n215 585
R97 B.n214 B.n213 585
R98 B.n212 B.n211 585
R99 B.n210 B.n209 585
R100 B.n208 B.n207 585
R101 B.n206 B.n205 585
R102 B.n204 B.n203 585
R103 B.n202 B.n201 585
R104 B.n200 B.n199 585
R105 B.n198 B.n197 585
R106 B.n196 B.n195 585
R107 B.n194 B.n193 585
R108 B.n192 B.n191 585
R109 B.n190 B.n189 585
R110 B.n188 B.n187 585
R111 B.n186 B.n185 585
R112 B.n184 B.n183 585
R113 B.n182 B.n181 585
R114 B.n180 B.n179 585
R115 B.n178 B.n177 585
R116 B.n176 B.n175 585
R117 B.n174 B.n173 585
R118 B.n172 B.n171 585
R119 B.n170 B.n169 585
R120 B.n168 B.n167 585
R121 B.n166 B.n165 585
R122 B.n164 B.n163 585
R123 B.n162 B.n161 585
R124 B.n160 B.n159 585
R125 B.n158 B.n157 585
R126 B.n156 B.n155 585
R127 B.n154 B.n153 585
R128 B.n152 B.n151 585
R129 B.n150 B.n149 585
R130 B.n148 B.n147 585
R131 B.n146 B.n145 585
R132 B.n144 B.n143 585
R133 B.n142 B.n141 585
R134 B.n140 B.n139 585
R135 B.n138 B.n137 585
R136 B.n136 B.n135 585
R137 B.n134 B.n133 585
R138 B.n132 B.n131 585
R139 B.n130 B.n129 585
R140 B.n128 B.n127 585
R141 B.n126 B.n125 585
R142 B.n124 B.n123 585
R143 B.n122 B.n121 585
R144 B.n120 B.n119 585
R145 B.n118 B.n117 585
R146 B.n116 B.n115 585
R147 B.n114 B.n113 585
R148 B.n112 B.n111 585
R149 B.n110 B.n109 585
R150 B.n108 B.n107 585
R151 B.n106 B.n105 585
R152 B.n104 B.n103 585
R153 B.n102 B.n101 585
R154 B.n100 B.n99 585
R155 B.n98 B.n97 585
R156 B.n96 B.n95 585
R157 B.n94 B.n93 585
R158 B.n92 B.n91 585
R159 B.n90 B.n89 585
R160 B.n88 B.n87 585
R161 B.n86 B.n85 585
R162 B.n84 B.n83 585
R163 B.n564 B.n33 585
R164 B.n569 B.n33 585
R165 B.n563 B.n32 585
R166 B.n570 B.n32 585
R167 B.n562 B.n561 585
R168 B.n561 B.n28 585
R169 B.n560 B.n27 585
R170 B.n576 B.n27 585
R171 B.n559 B.n26 585
R172 B.n577 B.n26 585
R173 B.n558 B.n25 585
R174 B.n578 B.n25 585
R175 B.n557 B.n556 585
R176 B.n556 B.n21 585
R177 B.n555 B.n20 585
R178 B.n584 B.n20 585
R179 B.n554 B.n19 585
R180 B.n585 B.n19 585
R181 B.n553 B.n18 585
R182 B.n586 B.n18 585
R183 B.n552 B.n551 585
R184 B.n551 B.n17 585
R185 B.n550 B.n12 585
R186 B.n592 B.n12 585
R187 B.n549 B.n11 585
R188 B.n593 B.n11 585
R189 B.n548 B.n10 585
R190 B.n594 B.n10 585
R191 B.n547 B.n7 585
R192 B.n597 B.n7 585
R193 B.n546 B.n6 585
R194 B.n598 B.n6 585
R195 B.n545 B.n5 585
R196 B.n599 B.n5 585
R197 B.n544 B.n543 585
R198 B.n543 B.n4 585
R199 B.n542 B.n252 585
R200 B.n542 B.n541 585
R201 B.n532 B.n253 585
R202 B.n254 B.n253 585
R203 B.n534 B.n533 585
R204 B.n535 B.n534 585
R205 B.n531 B.n258 585
R206 B.n261 B.n258 585
R207 B.n530 B.n529 585
R208 B.n529 B.n528 585
R209 B.n260 B.n259 585
R210 B.n521 B.n260 585
R211 B.n520 B.n519 585
R212 B.n522 B.n520 585
R213 B.n518 B.n266 585
R214 B.n266 B.n265 585
R215 B.n517 B.n516 585
R216 B.n516 B.n515 585
R217 B.n268 B.n267 585
R218 B.n269 B.n268 585
R219 B.n508 B.n507 585
R220 B.n509 B.n508 585
R221 B.n506 B.n274 585
R222 B.n274 B.n273 585
R223 B.n505 B.n504 585
R224 B.n504 B.n503 585
R225 B.n276 B.n275 585
R226 B.n277 B.n276 585
R227 B.n499 B.n498 585
R228 B.n280 B.n279 585
R229 B.n495 B.n494 585
R230 B.n496 B.n495 585
R231 B.n493 B.n323 585
R232 B.n492 B.n491 585
R233 B.n490 B.n489 585
R234 B.n488 B.n487 585
R235 B.n486 B.n485 585
R236 B.n484 B.n483 585
R237 B.n482 B.n481 585
R238 B.n480 B.n479 585
R239 B.n478 B.n477 585
R240 B.n476 B.n475 585
R241 B.n474 B.n473 585
R242 B.n472 B.n471 585
R243 B.n470 B.n469 585
R244 B.n468 B.n467 585
R245 B.n466 B.n465 585
R246 B.n464 B.n463 585
R247 B.n462 B.n461 585
R248 B.n460 B.n459 585
R249 B.n458 B.n457 585
R250 B.n456 B.n455 585
R251 B.n454 B.n453 585
R252 B.n452 B.n451 585
R253 B.n450 B.n449 585
R254 B.n448 B.n447 585
R255 B.n446 B.n445 585
R256 B.n444 B.n443 585
R257 B.n442 B.n441 585
R258 B.n440 B.n439 585
R259 B.n438 B.n437 585
R260 B.n436 B.n435 585
R261 B.n434 B.n433 585
R262 B.n432 B.n431 585
R263 B.n430 B.n429 585
R264 B.n428 B.n427 585
R265 B.n426 B.n425 585
R266 B.n423 B.n422 585
R267 B.n421 B.n420 585
R268 B.n419 B.n418 585
R269 B.n417 B.n416 585
R270 B.n415 B.n414 585
R271 B.n413 B.n412 585
R272 B.n411 B.n410 585
R273 B.n409 B.n408 585
R274 B.n407 B.n406 585
R275 B.n405 B.n404 585
R276 B.n402 B.n401 585
R277 B.n400 B.n399 585
R278 B.n398 B.n397 585
R279 B.n396 B.n395 585
R280 B.n394 B.n393 585
R281 B.n392 B.n391 585
R282 B.n390 B.n389 585
R283 B.n388 B.n387 585
R284 B.n386 B.n385 585
R285 B.n384 B.n383 585
R286 B.n382 B.n381 585
R287 B.n380 B.n379 585
R288 B.n378 B.n377 585
R289 B.n376 B.n375 585
R290 B.n374 B.n373 585
R291 B.n372 B.n371 585
R292 B.n370 B.n369 585
R293 B.n368 B.n367 585
R294 B.n366 B.n365 585
R295 B.n364 B.n363 585
R296 B.n362 B.n361 585
R297 B.n360 B.n359 585
R298 B.n358 B.n357 585
R299 B.n356 B.n355 585
R300 B.n354 B.n353 585
R301 B.n352 B.n351 585
R302 B.n350 B.n349 585
R303 B.n348 B.n347 585
R304 B.n346 B.n345 585
R305 B.n344 B.n343 585
R306 B.n342 B.n341 585
R307 B.n340 B.n339 585
R308 B.n338 B.n337 585
R309 B.n336 B.n335 585
R310 B.n334 B.n333 585
R311 B.n332 B.n331 585
R312 B.n330 B.n329 585
R313 B.n328 B.n322 585
R314 B.n496 B.n322 585
R315 B.n500 B.n278 585
R316 B.n278 B.n277 585
R317 B.n502 B.n501 585
R318 B.n503 B.n502 585
R319 B.n272 B.n271 585
R320 B.n273 B.n272 585
R321 B.n511 B.n510 585
R322 B.n510 B.n509 585
R323 B.n512 B.n270 585
R324 B.n270 B.n269 585
R325 B.n514 B.n513 585
R326 B.n515 B.n514 585
R327 B.n264 B.n263 585
R328 B.n265 B.n264 585
R329 B.n524 B.n523 585
R330 B.n523 B.n522 585
R331 B.n525 B.n262 585
R332 B.n521 B.n262 585
R333 B.n527 B.n526 585
R334 B.n528 B.n527 585
R335 B.n257 B.n256 585
R336 B.n261 B.n257 585
R337 B.n537 B.n536 585
R338 B.n536 B.n535 585
R339 B.n538 B.n255 585
R340 B.n255 B.n254 585
R341 B.n540 B.n539 585
R342 B.n541 B.n540 585
R343 B.n3 B.n0 585
R344 B.n4 B.n3 585
R345 B.n596 B.n1 585
R346 B.n597 B.n596 585
R347 B.n595 B.n9 585
R348 B.n595 B.n594 585
R349 B.n14 B.n8 585
R350 B.n593 B.n8 585
R351 B.n591 B.n590 585
R352 B.n592 B.n591 585
R353 B.n589 B.n13 585
R354 B.n17 B.n13 585
R355 B.n588 B.n587 585
R356 B.n587 B.n586 585
R357 B.n16 B.n15 585
R358 B.n585 B.n16 585
R359 B.n583 B.n582 585
R360 B.n584 B.n583 585
R361 B.n581 B.n22 585
R362 B.n22 B.n21 585
R363 B.n580 B.n579 585
R364 B.n579 B.n578 585
R365 B.n24 B.n23 585
R366 B.n577 B.n24 585
R367 B.n575 B.n574 585
R368 B.n576 B.n575 585
R369 B.n573 B.n29 585
R370 B.n29 B.n28 585
R371 B.n572 B.n571 585
R372 B.n571 B.n570 585
R373 B.n31 B.n30 585
R374 B.n569 B.n31 585
R375 B.n600 B.n599 585
R376 B.n598 B.n2 585
R377 B.n83 B.n31 578.989
R378 B.n566 B.n33 578.989
R379 B.n322 B.n276 578.989
R380 B.n498 B.n278 578.989
R381 B.n568 B.n567 256.663
R382 B.n568 B.n75 256.663
R383 B.n568 B.n74 256.663
R384 B.n568 B.n73 256.663
R385 B.n568 B.n72 256.663
R386 B.n568 B.n71 256.663
R387 B.n568 B.n70 256.663
R388 B.n568 B.n69 256.663
R389 B.n568 B.n68 256.663
R390 B.n568 B.n67 256.663
R391 B.n568 B.n66 256.663
R392 B.n568 B.n65 256.663
R393 B.n568 B.n64 256.663
R394 B.n568 B.n63 256.663
R395 B.n568 B.n62 256.663
R396 B.n568 B.n61 256.663
R397 B.n568 B.n60 256.663
R398 B.n568 B.n59 256.663
R399 B.n568 B.n58 256.663
R400 B.n568 B.n57 256.663
R401 B.n568 B.n56 256.663
R402 B.n568 B.n55 256.663
R403 B.n568 B.n54 256.663
R404 B.n568 B.n53 256.663
R405 B.n568 B.n52 256.663
R406 B.n568 B.n51 256.663
R407 B.n568 B.n50 256.663
R408 B.n568 B.n49 256.663
R409 B.n568 B.n48 256.663
R410 B.n568 B.n47 256.663
R411 B.n568 B.n46 256.663
R412 B.n568 B.n45 256.663
R413 B.n568 B.n44 256.663
R414 B.n568 B.n43 256.663
R415 B.n568 B.n42 256.663
R416 B.n568 B.n41 256.663
R417 B.n568 B.n40 256.663
R418 B.n568 B.n39 256.663
R419 B.n568 B.n38 256.663
R420 B.n568 B.n37 256.663
R421 B.n568 B.n36 256.663
R422 B.n568 B.n35 256.663
R423 B.n568 B.n34 256.663
R424 B.n497 B.n496 256.663
R425 B.n496 B.n281 256.663
R426 B.n496 B.n282 256.663
R427 B.n496 B.n283 256.663
R428 B.n496 B.n284 256.663
R429 B.n496 B.n285 256.663
R430 B.n496 B.n286 256.663
R431 B.n496 B.n287 256.663
R432 B.n496 B.n288 256.663
R433 B.n496 B.n289 256.663
R434 B.n496 B.n290 256.663
R435 B.n496 B.n291 256.663
R436 B.n496 B.n292 256.663
R437 B.n496 B.n293 256.663
R438 B.n496 B.n294 256.663
R439 B.n496 B.n295 256.663
R440 B.n496 B.n296 256.663
R441 B.n496 B.n297 256.663
R442 B.n496 B.n298 256.663
R443 B.n496 B.n299 256.663
R444 B.n496 B.n300 256.663
R445 B.n496 B.n301 256.663
R446 B.n496 B.n302 256.663
R447 B.n496 B.n303 256.663
R448 B.n496 B.n304 256.663
R449 B.n496 B.n305 256.663
R450 B.n496 B.n306 256.663
R451 B.n496 B.n307 256.663
R452 B.n496 B.n308 256.663
R453 B.n496 B.n309 256.663
R454 B.n496 B.n310 256.663
R455 B.n496 B.n311 256.663
R456 B.n496 B.n312 256.663
R457 B.n496 B.n313 256.663
R458 B.n496 B.n314 256.663
R459 B.n496 B.n315 256.663
R460 B.n496 B.n316 256.663
R461 B.n496 B.n317 256.663
R462 B.n496 B.n318 256.663
R463 B.n496 B.n319 256.663
R464 B.n496 B.n320 256.663
R465 B.n496 B.n321 256.663
R466 B.n602 B.n601 256.663
R467 B.n87 B.n86 163.367
R468 B.n91 B.n90 163.367
R469 B.n95 B.n94 163.367
R470 B.n99 B.n98 163.367
R471 B.n103 B.n102 163.367
R472 B.n107 B.n106 163.367
R473 B.n111 B.n110 163.367
R474 B.n115 B.n114 163.367
R475 B.n119 B.n118 163.367
R476 B.n123 B.n122 163.367
R477 B.n127 B.n126 163.367
R478 B.n131 B.n130 163.367
R479 B.n135 B.n134 163.367
R480 B.n139 B.n138 163.367
R481 B.n143 B.n142 163.367
R482 B.n147 B.n146 163.367
R483 B.n151 B.n150 163.367
R484 B.n155 B.n154 163.367
R485 B.n159 B.n158 163.367
R486 B.n163 B.n162 163.367
R487 B.n167 B.n166 163.367
R488 B.n171 B.n170 163.367
R489 B.n175 B.n174 163.367
R490 B.n179 B.n178 163.367
R491 B.n183 B.n182 163.367
R492 B.n187 B.n186 163.367
R493 B.n191 B.n190 163.367
R494 B.n195 B.n194 163.367
R495 B.n199 B.n198 163.367
R496 B.n203 B.n202 163.367
R497 B.n207 B.n206 163.367
R498 B.n211 B.n210 163.367
R499 B.n215 B.n214 163.367
R500 B.n219 B.n218 163.367
R501 B.n223 B.n222 163.367
R502 B.n227 B.n226 163.367
R503 B.n231 B.n230 163.367
R504 B.n235 B.n234 163.367
R505 B.n239 B.n238 163.367
R506 B.n243 B.n242 163.367
R507 B.n247 B.n246 163.367
R508 B.n249 B.n76 163.367
R509 B.n504 B.n276 163.367
R510 B.n504 B.n274 163.367
R511 B.n508 B.n274 163.367
R512 B.n508 B.n268 163.367
R513 B.n516 B.n268 163.367
R514 B.n516 B.n266 163.367
R515 B.n520 B.n266 163.367
R516 B.n520 B.n260 163.367
R517 B.n529 B.n260 163.367
R518 B.n529 B.n258 163.367
R519 B.n534 B.n258 163.367
R520 B.n534 B.n253 163.367
R521 B.n542 B.n253 163.367
R522 B.n543 B.n542 163.367
R523 B.n543 B.n5 163.367
R524 B.n6 B.n5 163.367
R525 B.n7 B.n6 163.367
R526 B.n10 B.n7 163.367
R527 B.n11 B.n10 163.367
R528 B.n12 B.n11 163.367
R529 B.n551 B.n12 163.367
R530 B.n551 B.n18 163.367
R531 B.n19 B.n18 163.367
R532 B.n20 B.n19 163.367
R533 B.n556 B.n20 163.367
R534 B.n556 B.n25 163.367
R535 B.n26 B.n25 163.367
R536 B.n27 B.n26 163.367
R537 B.n561 B.n27 163.367
R538 B.n561 B.n32 163.367
R539 B.n33 B.n32 163.367
R540 B.n495 B.n280 163.367
R541 B.n495 B.n323 163.367
R542 B.n491 B.n490 163.367
R543 B.n487 B.n486 163.367
R544 B.n483 B.n482 163.367
R545 B.n479 B.n478 163.367
R546 B.n475 B.n474 163.367
R547 B.n471 B.n470 163.367
R548 B.n467 B.n466 163.367
R549 B.n463 B.n462 163.367
R550 B.n459 B.n458 163.367
R551 B.n455 B.n454 163.367
R552 B.n451 B.n450 163.367
R553 B.n447 B.n446 163.367
R554 B.n443 B.n442 163.367
R555 B.n439 B.n438 163.367
R556 B.n435 B.n434 163.367
R557 B.n431 B.n430 163.367
R558 B.n427 B.n426 163.367
R559 B.n422 B.n421 163.367
R560 B.n418 B.n417 163.367
R561 B.n414 B.n413 163.367
R562 B.n410 B.n409 163.367
R563 B.n406 B.n405 163.367
R564 B.n401 B.n400 163.367
R565 B.n397 B.n396 163.367
R566 B.n393 B.n392 163.367
R567 B.n389 B.n388 163.367
R568 B.n385 B.n384 163.367
R569 B.n381 B.n380 163.367
R570 B.n377 B.n376 163.367
R571 B.n373 B.n372 163.367
R572 B.n369 B.n368 163.367
R573 B.n365 B.n364 163.367
R574 B.n361 B.n360 163.367
R575 B.n357 B.n356 163.367
R576 B.n353 B.n352 163.367
R577 B.n349 B.n348 163.367
R578 B.n345 B.n344 163.367
R579 B.n341 B.n340 163.367
R580 B.n337 B.n336 163.367
R581 B.n333 B.n332 163.367
R582 B.n329 B.n322 163.367
R583 B.n502 B.n278 163.367
R584 B.n502 B.n272 163.367
R585 B.n510 B.n272 163.367
R586 B.n510 B.n270 163.367
R587 B.n514 B.n270 163.367
R588 B.n514 B.n264 163.367
R589 B.n523 B.n264 163.367
R590 B.n523 B.n262 163.367
R591 B.n527 B.n262 163.367
R592 B.n527 B.n257 163.367
R593 B.n536 B.n257 163.367
R594 B.n536 B.n255 163.367
R595 B.n540 B.n255 163.367
R596 B.n540 B.n3 163.367
R597 B.n600 B.n3 163.367
R598 B.n596 B.n2 163.367
R599 B.n596 B.n595 163.367
R600 B.n595 B.n8 163.367
R601 B.n591 B.n8 163.367
R602 B.n591 B.n13 163.367
R603 B.n587 B.n13 163.367
R604 B.n587 B.n16 163.367
R605 B.n583 B.n16 163.367
R606 B.n583 B.n22 163.367
R607 B.n579 B.n22 163.367
R608 B.n579 B.n24 163.367
R609 B.n575 B.n24 163.367
R610 B.n575 B.n29 163.367
R611 B.n571 B.n29 163.367
R612 B.n571 B.n31 163.367
R613 B.n496 B.n277 95.7708
R614 B.n569 B.n568 95.7708
R615 B.n77 B.t14 78.8122
R616 B.n326 B.t21 78.8122
R617 B.n80 B.t17 78.7985
R618 B.n324 B.t11 78.7985
R619 B.n83 B.n34 71.676
R620 B.n87 B.n35 71.676
R621 B.n91 B.n36 71.676
R622 B.n95 B.n37 71.676
R623 B.n99 B.n38 71.676
R624 B.n103 B.n39 71.676
R625 B.n107 B.n40 71.676
R626 B.n111 B.n41 71.676
R627 B.n115 B.n42 71.676
R628 B.n119 B.n43 71.676
R629 B.n123 B.n44 71.676
R630 B.n127 B.n45 71.676
R631 B.n131 B.n46 71.676
R632 B.n135 B.n47 71.676
R633 B.n139 B.n48 71.676
R634 B.n143 B.n49 71.676
R635 B.n147 B.n50 71.676
R636 B.n151 B.n51 71.676
R637 B.n155 B.n52 71.676
R638 B.n159 B.n53 71.676
R639 B.n163 B.n54 71.676
R640 B.n167 B.n55 71.676
R641 B.n171 B.n56 71.676
R642 B.n175 B.n57 71.676
R643 B.n179 B.n58 71.676
R644 B.n183 B.n59 71.676
R645 B.n187 B.n60 71.676
R646 B.n191 B.n61 71.676
R647 B.n195 B.n62 71.676
R648 B.n199 B.n63 71.676
R649 B.n203 B.n64 71.676
R650 B.n207 B.n65 71.676
R651 B.n211 B.n66 71.676
R652 B.n215 B.n67 71.676
R653 B.n219 B.n68 71.676
R654 B.n223 B.n69 71.676
R655 B.n227 B.n70 71.676
R656 B.n231 B.n71 71.676
R657 B.n235 B.n72 71.676
R658 B.n239 B.n73 71.676
R659 B.n243 B.n74 71.676
R660 B.n247 B.n75 71.676
R661 B.n567 B.n76 71.676
R662 B.n567 B.n566 71.676
R663 B.n249 B.n75 71.676
R664 B.n246 B.n74 71.676
R665 B.n242 B.n73 71.676
R666 B.n238 B.n72 71.676
R667 B.n234 B.n71 71.676
R668 B.n230 B.n70 71.676
R669 B.n226 B.n69 71.676
R670 B.n222 B.n68 71.676
R671 B.n218 B.n67 71.676
R672 B.n214 B.n66 71.676
R673 B.n210 B.n65 71.676
R674 B.n206 B.n64 71.676
R675 B.n202 B.n63 71.676
R676 B.n198 B.n62 71.676
R677 B.n194 B.n61 71.676
R678 B.n190 B.n60 71.676
R679 B.n186 B.n59 71.676
R680 B.n182 B.n58 71.676
R681 B.n178 B.n57 71.676
R682 B.n174 B.n56 71.676
R683 B.n170 B.n55 71.676
R684 B.n166 B.n54 71.676
R685 B.n162 B.n53 71.676
R686 B.n158 B.n52 71.676
R687 B.n154 B.n51 71.676
R688 B.n150 B.n50 71.676
R689 B.n146 B.n49 71.676
R690 B.n142 B.n48 71.676
R691 B.n138 B.n47 71.676
R692 B.n134 B.n46 71.676
R693 B.n130 B.n45 71.676
R694 B.n126 B.n44 71.676
R695 B.n122 B.n43 71.676
R696 B.n118 B.n42 71.676
R697 B.n114 B.n41 71.676
R698 B.n110 B.n40 71.676
R699 B.n106 B.n39 71.676
R700 B.n102 B.n38 71.676
R701 B.n98 B.n37 71.676
R702 B.n94 B.n36 71.676
R703 B.n90 B.n35 71.676
R704 B.n86 B.n34 71.676
R705 B.n498 B.n497 71.676
R706 B.n323 B.n281 71.676
R707 B.n490 B.n282 71.676
R708 B.n486 B.n283 71.676
R709 B.n482 B.n284 71.676
R710 B.n478 B.n285 71.676
R711 B.n474 B.n286 71.676
R712 B.n470 B.n287 71.676
R713 B.n466 B.n288 71.676
R714 B.n462 B.n289 71.676
R715 B.n458 B.n290 71.676
R716 B.n454 B.n291 71.676
R717 B.n450 B.n292 71.676
R718 B.n446 B.n293 71.676
R719 B.n442 B.n294 71.676
R720 B.n438 B.n295 71.676
R721 B.n434 B.n296 71.676
R722 B.n430 B.n297 71.676
R723 B.n426 B.n298 71.676
R724 B.n421 B.n299 71.676
R725 B.n417 B.n300 71.676
R726 B.n413 B.n301 71.676
R727 B.n409 B.n302 71.676
R728 B.n405 B.n303 71.676
R729 B.n400 B.n304 71.676
R730 B.n396 B.n305 71.676
R731 B.n392 B.n306 71.676
R732 B.n388 B.n307 71.676
R733 B.n384 B.n308 71.676
R734 B.n380 B.n309 71.676
R735 B.n376 B.n310 71.676
R736 B.n372 B.n311 71.676
R737 B.n368 B.n312 71.676
R738 B.n364 B.n313 71.676
R739 B.n360 B.n314 71.676
R740 B.n356 B.n315 71.676
R741 B.n352 B.n316 71.676
R742 B.n348 B.n317 71.676
R743 B.n344 B.n318 71.676
R744 B.n340 B.n319 71.676
R745 B.n336 B.n320 71.676
R746 B.n332 B.n321 71.676
R747 B.n497 B.n280 71.676
R748 B.n491 B.n281 71.676
R749 B.n487 B.n282 71.676
R750 B.n483 B.n283 71.676
R751 B.n479 B.n284 71.676
R752 B.n475 B.n285 71.676
R753 B.n471 B.n286 71.676
R754 B.n467 B.n287 71.676
R755 B.n463 B.n288 71.676
R756 B.n459 B.n289 71.676
R757 B.n455 B.n290 71.676
R758 B.n451 B.n291 71.676
R759 B.n447 B.n292 71.676
R760 B.n443 B.n293 71.676
R761 B.n439 B.n294 71.676
R762 B.n435 B.n295 71.676
R763 B.n431 B.n296 71.676
R764 B.n427 B.n297 71.676
R765 B.n422 B.n298 71.676
R766 B.n418 B.n299 71.676
R767 B.n414 B.n300 71.676
R768 B.n410 B.n301 71.676
R769 B.n406 B.n302 71.676
R770 B.n401 B.n303 71.676
R771 B.n397 B.n304 71.676
R772 B.n393 B.n305 71.676
R773 B.n389 B.n306 71.676
R774 B.n385 B.n307 71.676
R775 B.n381 B.n308 71.676
R776 B.n377 B.n309 71.676
R777 B.n373 B.n310 71.676
R778 B.n369 B.n311 71.676
R779 B.n365 B.n312 71.676
R780 B.n361 B.n313 71.676
R781 B.n357 B.n314 71.676
R782 B.n353 B.n315 71.676
R783 B.n349 B.n316 71.676
R784 B.n345 B.n317 71.676
R785 B.n341 B.n318 71.676
R786 B.n337 B.n319 71.676
R787 B.n333 B.n320 71.676
R788 B.n329 B.n321 71.676
R789 B.n601 B.n600 71.676
R790 B.n601 B.n2 71.676
R791 B.n78 B.t15 68.7273
R792 B.n327 B.t20 68.7273
R793 B.n81 B.t18 68.7136
R794 B.n325 B.t10 68.7136
R795 B.n82 B.n81 59.5399
R796 B.n79 B.n78 59.5399
R797 B.n403 B.n327 59.5399
R798 B.n424 B.n325 59.5399
R799 B.n503 B.n277 46.1876
R800 B.n503 B.n273 46.1876
R801 B.n509 B.n273 46.1876
R802 B.n515 B.n269 46.1876
R803 B.n515 B.n265 46.1876
R804 B.n522 B.n265 46.1876
R805 B.n522 B.n521 46.1876
R806 B.n528 B.n261 46.1876
R807 B.n541 B.n254 46.1876
R808 B.n599 B.n4 46.1876
R809 B.n599 B.n598 46.1876
R810 B.n598 B.n597 46.1876
R811 B.n594 B.n593 46.1876
R812 B.n586 B.n17 46.1876
R813 B.n585 B.n584 46.1876
R814 B.n584 B.n21 46.1876
R815 B.n578 B.n21 46.1876
R816 B.n578 B.n577 46.1876
R817 B.n576 B.n28 46.1876
R818 B.n570 B.n28 46.1876
R819 B.n570 B.n569 46.1876
R820 B.n535 B.t7 42.7915
R821 B.n592 B.t0 42.7915
R822 B.t4 B.n4 40.0746
R823 B.n597 B.t2 40.0746
R824 B.n500 B.n499 37.62
R825 B.n328 B.n275 37.62
R826 B.n565 B.n564 37.62
R827 B.n84 B.n30 37.62
R828 B.n509 B.t9 37.3577
R829 B.t13 B.n576 37.3577
R830 B.n535 B.t1 27.8486
R831 B.t3 B.n592 27.8486
R832 B.n521 B.t5 25.1317
R833 B.t6 B.n585 25.1317
R834 B.n528 B.t5 21.0564
R835 B.n586 B.t6 21.0564
R836 B.t1 B.n254 18.3395
R837 B.n593 B.t3 18.3395
R838 B B.n602 18.0485
R839 B.n501 B.n500 10.6151
R840 B.n501 B.n271 10.6151
R841 B.n511 B.n271 10.6151
R842 B.n512 B.n511 10.6151
R843 B.n513 B.n512 10.6151
R844 B.n513 B.n263 10.6151
R845 B.n524 B.n263 10.6151
R846 B.n525 B.n524 10.6151
R847 B.n526 B.n525 10.6151
R848 B.n526 B.n256 10.6151
R849 B.n537 B.n256 10.6151
R850 B.n538 B.n537 10.6151
R851 B.n539 B.n538 10.6151
R852 B.n539 B.n0 10.6151
R853 B.n499 B.n279 10.6151
R854 B.n494 B.n279 10.6151
R855 B.n494 B.n493 10.6151
R856 B.n493 B.n492 10.6151
R857 B.n492 B.n489 10.6151
R858 B.n489 B.n488 10.6151
R859 B.n488 B.n485 10.6151
R860 B.n485 B.n484 10.6151
R861 B.n484 B.n481 10.6151
R862 B.n481 B.n480 10.6151
R863 B.n480 B.n477 10.6151
R864 B.n477 B.n476 10.6151
R865 B.n476 B.n473 10.6151
R866 B.n473 B.n472 10.6151
R867 B.n472 B.n469 10.6151
R868 B.n469 B.n468 10.6151
R869 B.n468 B.n465 10.6151
R870 B.n465 B.n464 10.6151
R871 B.n464 B.n461 10.6151
R872 B.n461 B.n460 10.6151
R873 B.n460 B.n457 10.6151
R874 B.n457 B.n456 10.6151
R875 B.n456 B.n453 10.6151
R876 B.n453 B.n452 10.6151
R877 B.n452 B.n449 10.6151
R878 B.n449 B.n448 10.6151
R879 B.n448 B.n445 10.6151
R880 B.n445 B.n444 10.6151
R881 B.n444 B.n441 10.6151
R882 B.n441 B.n440 10.6151
R883 B.n440 B.n437 10.6151
R884 B.n437 B.n436 10.6151
R885 B.n436 B.n433 10.6151
R886 B.n433 B.n432 10.6151
R887 B.n432 B.n429 10.6151
R888 B.n429 B.n428 10.6151
R889 B.n428 B.n425 10.6151
R890 B.n423 B.n420 10.6151
R891 B.n420 B.n419 10.6151
R892 B.n419 B.n416 10.6151
R893 B.n416 B.n415 10.6151
R894 B.n415 B.n412 10.6151
R895 B.n412 B.n411 10.6151
R896 B.n411 B.n408 10.6151
R897 B.n408 B.n407 10.6151
R898 B.n407 B.n404 10.6151
R899 B.n402 B.n399 10.6151
R900 B.n399 B.n398 10.6151
R901 B.n398 B.n395 10.6151
R902 B.n395 B.n394 10.6151
R903 B.n394 B.n391 10.6151
R904 B.n391 B.n390 10.6151
R905 B.n390 B.n387 10.6151
R906 B.n387 B.n386 10.6151
R907 B.n386 B.n383 10.6151
R908 B.n383 B.n382 10.6151
R909 B.n382 B.n379 10.6151
R910 B.n379 B.n378 10.6151
R911 B.n378 B.n375 10.6151
R912 B.n375 B.n374 10.6151
R913 B.n374 B.n371 10.6151
R914 B.n371 B.n370 10.6151
R915 B.n370 B.n367 10.6151
R916 B.n367 B.n366 10.6151
R917 B.n366 B.n363 10.6151
R918 B.n363 B.n362 10.6151
R919 B.n362 B.n359 10.6151
R920 B.n359 B.n358 10.6151
R921 B.n358 B.n355 10.6151
R922 B.n355 B.n354 10.6151
R923 B.n354 B.n351 10.6151
R924 B.n351 B.n350 10.6151
R925 B.n350 B.n347 10.6151
R926 B.n347 B.n346 10.6151
R927 B.n346 B.n343 10.6151
R928 B.n343 B.n342 10.6151
R929 B.n342 B.n339 10.6151
R930 B.n339 B.n338 10.6151
R931 B.n338 B.n335 10.6151
R932 B.n335 B.n334 10.6151
R933 B.n334 B.n331 10.6151
R934 B.n331 B.n330 10.6151
R935 B.n330 B.n328 10.6151
R936 B.n505 B.n275 10.6151
R937 B.n506 B.n505 10.6151
R938 B.n507 B.n506 10.6151
R939 B.n507 B.n267 10.6151
R940 B.n517 B.n267 10.6151
R941 B.n518 B.n517 10.6151
R942 B.n519 B.n518 10.6151
R943 B.n519 B.n259 10.6151
R944 B.n530 B.n259 10.6151
R945 B.n531 B.n530 10.6151
R946 B.n533 B.n531 10.6151
R947 B.n533 B.n532 10.6151
R948 B.n532 B.n252 10.6151
R949 B.n544 B.n252 10.6151
R950 B.n545 B.n544 10.6151
R951 B.n546 B.n545 10.6151
R952 B.n547 B.n546 10.6151
R953 B.n548 B.n547 10.6151
R954 B.n549 B.n548 10.6151
R955 B.n550 B.n549 10.6151
R956 B.n552 B.n550 10.6151
R957 B.n553 B.n552 10.6151
R958 B.n554 B.n553 10.6151
R959 B.n555 B.n554 10.6151
R960 B.n557 B.n555 10.6151
R961 B.n558 B.n557 10.6151
R962 B.n559 B.n558 10.6151
R963 B.n560 B.n559 10.6151
R964 B.n562 B.n560 10.6151
R965 B.n563 B.n562 10.6151
R966 B.n564 B.n563 10.6151
R967 B.n9 B.n1 10.6151
R968 B.n14 B.n9 10.6151
R969 B.n590 B.n14 10.6151
R970 B.n590 B.n589 10.6151
R971 B.n589 B.n588 10.6151
R972 B.n588 B.n15 10.6151
R973 B.n582 B.n15 10.6151
R974 B.n582 B.n581 10.6151
R975 B.n581 B.n580 10.6151
R976 B.n580 B.n23 10.6151
R977 B.n574 B.n23 10.6151
R978 B.n574 B.n573 10.6151
R979 B.n573 B.n572 10.6151
R980 B.n572 B.n30 10.6151
R981 B.n85 B.n84 10.6151
R982 B.n88 B.n85 10.6151
R983 B.n89 B.n88 10.6151
R984 B.n92 B.n89 10.6151
R985 B.n93 B.n92 10.6151
R986 B.n96 B.n93 10.6151
R987 B.n97 B.n96 10.6151
R988 B.n100 B.n97 10.6151
R989 B.n101 B.n100 10.6151
R990 B.n104 B.n101 10.6151
R991 B.n105 B.n104 10.6151
R992 B.n108 B.n105 10.6151
R993 B.n109 B.n108 10.6151
R994 B.n112 B.n109 10.6151
R995 B.n113 B.n112 10.6151
R996 B.n116 B.n113 10.6151
R997 B.n117 B.n116 10.6151
R998 B.n120 B.n117 10.6151
R999 B.n121 B.n120 10.6151
R1000 B.n124 B.n121 10.6151
R1001 B.n125 B.n124 10.6151
R1002 B.n128 B.n125 10.6151
R1003 B.n129 B.n128 10.6151
R1004 B.n132 B.n129 10.6151
R1005 B.n133 B.n132 10.6151
R1006 B.n136 B.n133 10.6151
R1007 B.n137 B.n136 10.6151
R1008 B.n140 B.n137 10.6151
R1009 B.n141 B.n140 10.6151
R1010 B.n144 B.n141 10.6151
R1011 B.n145 B.n144 10.6151
R1012 B.n148 B.n145 10.6151
R1013 B.n149 B.n148 10.6151
R1014 B.n152 B.n149 10.6151
R1015 B.n153 B.n152 10.6151
R1016 B.n156 B.n153 10.6151
R1017 B.n157 B.n156 10.6151
R1018 B.n161 B.n160 10.6151
R1019 B.n164 B.n161 10.6151
R1020 B.n165 B.n164 10.6151
R1021 B.n168 B.n165 10.6151
R1022 B.n169 B.n168 10.6151
R1023 B.n172 B.n169 10.6151
R1024 B.n173 B.n172 10.6151
R1025 B.n176 B.n173 10.6151
R1026 B.n177 B.n176 10.6151
R1027 B.n181 B.n180 10.6151
R1028 B.n184 B.n181 10.6151
R1029 B.n185 B.n184 10.6151
R1030 B.n188 B.n185 10.6151
R1031 B.n189 B.n188 10.6151
R1032 B.n192 B.n189 10.6151
R1033 B.n193 B.n192 10.6151
R1034 B.n196 B.n193 10.6151
R1035 B.n197 B.n196 10.6151
R1036 B.n200 B.n197 10.6151
R1037 B.n201 B.n200 10.6151
R1038 B.n204 B.n201 10.6151
R1039 B.n205 B.n204 10.6151
R1040 B.n208 B.n205 10.6151
R1041 B.n209 B.n208 10.6151
R1042 B.n212 B.n209 10.6151
R1043 B.n213 B.n212 10.6151
R1044 B.n216 B.n213 10.6151
R1045 B.n217 B.n216 10.6151
R1046 B.n220 B.n217 10.6151
R1047 B.n221 B.n220 10.6151
R1048 B.n224 B.n221 10.6151
R1049 B.n225 B.n224 10.6151
R1050 B.n228 B.n225 10.6151
R1051 B.n229 B.n228 10.6151
R1052 B.n232 B.n229 10.6151
R1053 B.n233 B.n232 10.6151
R1054 B.n236 B.n233 10.6151
R1055 B.n237 B.n236 10.6151
R1056 B.n240 B.n237 10.6151
R1057 B.n241 B.n240 10.6151
R1058 B.n244 B.n241 10.6151
R1059 B.n245 B.n244 10.6151
R1060 B.n248 B.n245 10.6151
R1061 B.n250 B.n248 10.6151
R1062 B.n251 B.n250 10.6151
R1063 B.n565 B.n251 10.6151
R1064 B.n81 B.n80 10.0853
R1065 B.n78 B.n77 10.0853
R1066 B.n327 B.n326 10.0853
R1067 B.n325 B.n324 10.0853
R1068 B.n425 B.n424 9.36635
R1069 B.n403 B.n402 9.36635
R1070 B.n157 B.n82 9.36635
R1071 B.n180 B.n79 9.36635
R1072 B.t9 B.n269 8.83039
R1073 B.n577 B.t13 8.83039
R1074 B.n602 B.n0 8.11757
R1075 B.n602 B.n1 8.11757
R1076 B.n541 B.t4 6.1135
R1077 B.n594 B.t2 6.1135
R1078 B.n261 B.t7 3.39661
R1079 B.n17 B.t0 3.39661
R1080 B.n424 B.n423 1.24928
R1081 B.n404 B.n403 1.24928
R1082 B.n160 B.n82 1.24928
R1083 B.n177 B.n79 1.24928
R1084 VP.n13 VP.t5 1590.91
R1085 VP.n9 VP.t4 1590.91
R1086 VP.n2 VP.t0 1590.91
R1087 VP.n6 VP.t1 1590.91
R1088 VP.n12 VP.t2 1550.01
R1089 VP.n10 VP.t6 1550.01
R1090 VP.n3 VP.t3 1550.01
R1091 VP.n5 VP.t7 1550.01
R1092 VP.n2 VP.n1 161.489
R1093 VP.n14 VP.n13 161.3
R1094 VP.n4 VP.n1 161.3
R1095 VP.n7 VP.n6 161.3
R1096 VP.n11 VP.n0 161.3
R1097 VP.n9 VP.n8 161.3
R1098 VP.n8 VP.n7 38.8414
R1099 VP.n11 VP.n10 37.9763
R1100 VP.n12 VP.n11 37.9763
R1101 VP.n4 VP.n3 37.9763
R1102 VP.n5 VP.n4 37.9763
R1103 VP.n10 VP.n9 35.055
R1104 VP.n13 VP.n12 35.055
R1105 VP.n3 VP.n2 35.055
R1106 VP.n6 VP.n5 35.055
R1107 VP.n7 VP.n1 0.189894
R1108 VP.n8 VP.n0 0.189894
R1109 VP.n14 VP.n0 0.189894
R1110 VP VP.n14 0.0516364
R1111 VDD1 VDD1.n0 60.1642
R1112 VDD1.n3 VDD1.n2 60.0504
R1113 VDD1.n3 VDD1.n1 60.0504
R1114 VDD1.n5 VDD1.n4 59.8817
R1115 VDD1.n5 VDD1.n3 35.7293
R1116 VDD1.n4 VDD1.t0 1.81369
R1117 VDD1.n4 VDD1.t6 1.81369
R1118 VDD1.n0 VDD1.t7 1.81369
R1119 VDD1.n0 VDD1.t4 1.81369
R1120 VDD1.n2 VDD1.t5 1.81369
R1121 VDD1.n2 VDD1.t2 1.81369
R1122 VDD1.n1 VDD1.t3 1.81369
R1123 VDD1.n1 VDD1.t1 1.81369
R1124 VDD1 VDD1.n5 0.166448
C0 VDD1 VP 2.45033f
C1 VP VN 4.51428f
C2 VTAIL VDD2 18.3053f
C3 VP VDD2 0.263052f
C4 VDD1 VN 0.147201f
C5 VDD1 VDD2 0.577749f
C6 VN VDD2 2.33465f
C7 VTAIL VP 1.89355f
C8 VTAIL VDD1 18.2671f
C9 VTAIL VN 1.87944f
C10 VDD2 B 2.989168f
C11 VDD1 B 3.159405f
C12 VTAIL B 7.739376f
C13 VN B 6.34759f
C14 VP B 4.560637f
C15 VDD1.t7 B 0.329944f
C16 VDD1.t4 B 0.329944f
C17 VDD1.n0 B 2.92066f
C18 VDD1.t3 B 0.329944f
C19 VDD1.t1 B 0.329944f
C20 VDD1.n1 B 2.91983f
C21 VDD1.t5 B 0.329944f
C22 VDD1.t2 B 0.329944f
C23 VDD1.n2 B 2.91983f
C24 VDD1.n3 B 2.85437f
C25 VDD1.t0 B 0.329944f
C26 VDD1.t6 B 0.329944f
C27 VDD1.n4 B 2.91866f
C28 VDD1.n5 B 3.15036f
C29 VP.n0 B 0.047884f
C30 VP.t2 B 0.280975f
C31 VP.t6 B 0.280975f
C32 VP.t4 B 0.284002f
C33 VP.n1 B 0.103084f
C34 VP.t7 B 0.280975f
C35 VP.t3 B 0.280975f
C36 VP.t0 B 0.284002f
C37 VP.n2 B 0.131246f
C38 VP.n3 B 0.118618f
C39 VP.n4 B 0.016475f
C40 VP.n5 B 0.118618f
C41 VP.t1 B 0.284002f
C42 VP.n6 B 0.131181f
C43 VP.n7 B 1.7286f
C44 VP.n8 B 1.77304f
C45 VP.n9 B 0.131181f
C46 VP.n10 B 0.118618f
C47 VP.n11 B 0.016475f
C48 VP.n12 B 0.118618f
C49 VP.t5 B 0.284002f
C50 VP.n13 B 0.131181f
C51 VP.n14 B 0.037108f
C52 VTAIL.t13 B 0.215224f
C53 VTAIL.t14 B 0.215224f
C54 VTAIL.n0 B 1.82559f
C55 VTAIL.n1 B 0.292573f
C56 VTAIL.t8 B 2.32405f
C57 VTAIL.n2 B 0.414167f
C58 VTAIL.t4 B 2.32405f
C59 VTAIL.n3 B 0.414167f
C60 VTAIL.t7 B 0.215224f
C61 VTAIL.t1 B 0.215224f
C62 VTAIL.n4 B 1.82559f
C63 VTAIL.n5 B 0.323923f
C64 VTAIL.t5 B 2.32405f
C65 VTAIL.n6 B 1.50778f
C66 VTAIL.t9 B 2.32407f
C67 VTAIL.n7 B 1.50776f
C68 VTAIL.t12 B 0.215224f
C69 VTAIL.t15 B 0.215224f
C70 VTAIL.n8 B 1.82559f
C71 VTAIL.n9 B 0.323916f
C72 VTAIL.t10 B 2.32407f
C73 VTAIL.n10 B 0.41415f
C74 VTAIL.t2 B 2.32407f
C75 VTAIL.n11 B 0.41415f
C76 VTAIL.t3 B 0.215224f
C77 VTAIL.t0 B 0.215224f
C78 VTAIL.n12 B 1.82559f
C79 VTAIL.n13 B 0.323916f
C80 VTAIL.t6 B 2.32405f
C81 VTAIL.n14 B 1.50778f
C82 VTAIL.t11 B 2.32405f
C83 VTAIL.n15 B 1.5031f
C84 VDD2.t1 B 0.329005f
C85 VDD2.t7 B 0.329005f
C86 VDD2.n0 B 2.91152f
C87 VDD2.t4 B 0.329005f
C88 VDD2.t3 B 0.329005f
C89 VDD2.n1 B 2.91152f
C90 VDD2.n2 B 2.76414f
C91 VDD2.t5 B 0.329005f
C92 VDD2.t6 B 0.329005f
C93 VDD2.n3 B 2.91036f
C94 VDD2.n4 B 3.09697f
C95 VDD2.t0 B 0.329005f
C96 VDD2.t2 B 0.329005f
C97 VDD2.n5 B 2.91148f
C98 VN.n0 B 0.099185f
C99 VN.t1 B 0.270348f
C100 VN.t2 B 0.270348f
C101 VN.t7 B 0.27326f
C102 VN.n1 B 0.126282f
C103 VN.n2 B 0.114132f
C104 VN.n3 B 0.015852f
C105 VN.n4 B 0.114132f
C106 VN.t4 B 0.27326f
C107 VN.n5 B 0.12622f
C108 VN.n6 B 0.035705f
C109 VN.n7 B 0.099185f
C110 VN.t6 B 0.27326f
C111 VN.t3 B 0.270348f
C112 VN.t0 B 0.270348f
C113 VN.t5 B 0.27326f
C114 VN.n8 B 0.126282f
C115 VN.n9 B 0.114132f
C116 VN.n10 B 0.015852f
C117 VN.n11 B 0.114132f
C118 VN.n12 B 0.12622f
C119 VN.n13 B 1.69362f
.ends

