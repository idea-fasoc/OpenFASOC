* NGSPICE file created from diff_pair_sample_1789.ext - technology: sky130A

.subckt diff_pair_sample_1789 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0.96195 ps=6.16 w=5.83 l=1.94
X1 VDD1.t8 VP.t1 VTAIL.t12 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0.96195 ps=6.16 w=5.83 l=1.94
X2 VTAIL.t15 VP.t2 VDD1.t7 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X3 VDD1.t6 VP.t3 VTAIL.t17 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=2.2737 ps=12.44 w=5.83 l=1.94
X4 B.t11 B.t9 B.t10 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0 ps=0 w=5.83 l=1.94
X5 VDD2.t9 VN.t0 VTAIL.t2 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X6 B.t8 B.t6 B.t7 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0 ps=0 w=5.83 l=1.94
X7 VDD1.t5 VP.t4 VTAIL.t16 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X8 VTAIL.t10 VP.t5 VDD1.t4 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X9 VTAIL.t0 VN.t1 VDD2.t8 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X10 VDD2.t7 VN.t2 VTAIL.t1 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=2.2737 ps=12.44 w=5.83 l=1.94
X11 VDD2.t6 VN.t3 VTAIL.t7 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X12 VDD1.t3 VP.t6 VTAIL.t18 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X13 VTAIL.t3 VN.t4 VDD2.t5 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X14 VTAIL.t8 VN.t5 VDD2.t4 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X15 B.t5 B.t3 B.t4 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0 ps=0 w=5.83 l=1.94
X16 VTAIL.t14 VP.t7 VDD1.t2 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X17 VDD2.t3 VN.t6 VTAIL.t4 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=2.2737 ps=12.44 w=5.83 l=1.94
X18 VTAIL.t9 VP.t8 VDD1.t1 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X19 VTAIL.t5 VN.t7 VDD2.t2 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=0.96195 ps=6.16 w=5.83 l=1.94
X20 VDD2.t1 VN.t8 VTAIL.t6 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0.96195 ps=6.16 w=5.83 l=1.94
X21 VDD1.t0 VP.t9 VTAIL.t13 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=0.96195 pd=6.16 as=2.2737 ps=12.44 w=5.83 l=1.94
X22 B.t2 B.t0 B.t1 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0 ps=0 w=5.83 l=1.94
X23 VDD2.t0 VN.t9 VTAIL.t19 w_n3694_n2134# sky130_fd_pr__pfet_01v8 ad=2.2737 pd=12.44 as=0.96195 ps=6.16 w=5.83 l=1.94
R0 VP.n44 VP.n43 183.81
R1 VP.n76 VP.n75 183.81
R2 VP.n42 VP.n41 183.81
R3 VP.n20 VP.n19 161.3
R4 VP.n21 VP.n16 161.3
R5 VP.n23 VP.n22 161.3
R6 VP.n24 VP.n15 161.3
R7 VP.n26 VP.n25 161.3
R8 VP.n27 VP.n14 161.3
R9 VP.n29 VP.n28 161.3
R10 VP.n30 VP.n13 161.3
R11 VP.n32 VP.n31 161.3
R12 VP.n34 VP.n12 161.3
R13 VP.n36 VP.n35 161.3
R14 VP.n37 VP.n11 161.3
R15 VP.n39 VP.n38 161.3
R16 VP.n40 VP.n10 161.3
R17 VP.n74 VP.n0 161.3
R18 VP.n73 VP.n72 161.3
R19 VP.n71 VP.n1 161.3
R20 VP.n70 VP.n69 161.3
R21 VP.n68 VP.n2 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n64 VP.n3 161.3
R24 VP.n63 VP.n62 161.3
R25 VP.n61 VP.n4 161.3
R26 VP.n60 VP.n59 161.3
R27 VP.n58 VP.n5 161.3
R28 VP.n57 VP.n56 161.3
R29 VP.n55 VP.n6 161.3
R30 VP.n54 VP.n53 161.3
R31 VP.n52 VP.n51 161.3
R32 VP.n50 VP.n8 161.3
R33 VP.n49 VP.n48 161.3
R34 VP.n47 VP.n9 161.3
R35 VP.n46 VP.n45 161.3
R36 VP.n18 VP.t1 105.222
R37 VP.n60 VP.t4 72.4247
R38 VP.n44 VP.t0 72.4247
R39 VP.n7 VP.t7 72.4247
R40 VP.n67 VP.t2 72.4247
R41 VP.n75 VP.t9 72.4247
R42 VP.n26 VP.t6 72.4247
R43 VP.n41 VP.t3 72.4247
R44 VP.n33 VP.t8 72.4247
R45 VP.n17 VP.t5 72.4247
R46 VP.n18 VP.n17 56.8484
R47 VP.n56 VP.n55 53.6055
R48 VP.n62 VP.n3 53.6055
R49 VP.n28 VP.n13 53.6055
R50 VP.n22 VP.n21 53.6055
R51 VP.n50 VP.n49 49.7204
R52 VP.n69 VP.n1 49.7204
R53 VP.n35 VP.n11 49.7204
R54 VP.n43 VP.n42 44.7619
R55 VP.n49 VP.n9 31.2664
R56 VP.n73 VP.n1 31.2664
R57 VP.n39 VP.n11 31.2664
R58 VP.n56 VP.n5 27.3813
R59 VP.n62 VP.n61 27.3813
R60 VP.n28 VP.n27 27.3813
R61 VP.n22 VP.n15 27.3813
R62 VP.n45 VP.n9 24.4675
R63 VP.n51 VP.n50 24.4675
R64 VP.n55 VP.n54 24.4675
R65 VP.n60 VP.n5 24.4675
R66 VP.n61 VP.n60 24.4675
R67 VP.n66 VP.n3 24.4675
R68 VP.n69 VP.n68 24.4675
R69 VP.n74 VP.n73 24.4675
R70 VP.n40 VP.n39 24.4675
R71 VP.n32 VP.n13 24.4675
R72 VP.n35 VP.n34 24.4675
R73 VP.n26 VP.n15 24.4675
R74 VP.n27 VP.n26 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 13.2127
R77 VP.n67 VP.n66 13.2127
R78 VP.n33 VP.n32 13.2127
R79 VP.n20 VP.n17 13.2127
R80 VP.n19 VP.n18 12.4717
R81 VP.n51 VP.n7 11.2553
R82 VP.n68 VP.n67 11.2553
R83 VP.n34 VP.n33 11.2553
R84 VP.n45 VP.n44 1.95786
R85 VP.n75 VP.n74 1.95786
R86 VP.n41 VP.n40 1.95786
R87 VP.n19 VP.n16 0.189894
R88 VP.n23 VP.n16 0.189894
R89 VP.n24 VP.n23 0.189894
R90 VP.n25 VP.n24 0.189894
R91 VP.n25 VP.n14 0.189894
R92 VP.n29 VP.n14 0.189894
R93 VP.n30 VP.n29 0.189894
R94 VP.n31 VP.n30 0.189894
R95 VP.n31 VP.n12 0.189894
R96 VP.n36 VP.n12 0.189894
R97 VP.n37 VP.n36 0.189894
R98 VP.n38 VP.n37 0.189894
R99 VP.n38 VP.n10 0.189894
R100 VP.n42 VP.n10 0.189894
R101 VP.n46 VP.n43 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n48 VP.n47 0.189894
R104 VP.n48 VP.n8 0.189894
R105 VP.n52 VP.n8 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n6 0.189894
R108 VP.n57 VP.n6 0.189894
R109 VP.n58 VP.n57 0.189894
R110 VP.n59 VP.n58 0.189894
R111 VP.n59 VP.n4 0.189894
R112 VP.n63 VP.n4 0.189894
R113 VP.n64 VP.n63 0.189894
R114 VP.n65 VP.n64 0.189894
R115 VP.n65 VP.n2 0.189894
R116 VP.n70 VP.n2 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n72 VP.n71 0.189894
R119 VP.n72 VP.n0 0.189894
R120 VP.n76 VP.n0 0.189894
R121 VP VP.n76 0.0516364
R122 VTAIL.n132 VTAIL.n131 756.745
R123 VTAIL.n30 VTAIL.n29 756.745
R124 VTAIL.n102 VTAIL.n101 756.745
R125 VTAIL.n68 VTAIL.n67 756.745
R126 VTAIL.n115 VTAIL.n114 585
R127 VTAIL.n117 VTAIL.n116 585
R128 VTAIL.n110 VTAIL.n109 585
R129 VTAIL.n123 VTAIL.n122 585
R130 VTAIL.n125 VTAIL.n124 585
R131 VTAIL.n106 VTAIL.n105 585
R132 VTAIL.n131 VTAIL.n130 585
R133 VTAIL.n13 VTAIL.n12 585
R134 VTAIL.n15 VTAIL.n14 585
R135 VTAIL.n8 VTAIL.n7 585
R136 VTAIL.n21 VTAIL.n20 585
R137 VTAIL.n23 VTAIL.n22 585
R138 VTAIL.n4 VTAIL.n3 585
R139 VTAIL.n29 VTAIL.n28 585
R140 VTAIL.n101 VTAIL.n100 585
R141 VTAIL.n76 VTAIL.n75 585
R142 VTAIL.n95 VTAIL.n94 585
R143 VTAIL.n93 VTAIL.n92 585
R144 VTAIL.n80 VTAIL.n79 585
R145 VTAIL.n87 VTAIL.n86 585
R146 VTAIL.n85 VTAIL.n84 585
R147 VTAIL.n67 VTAIL.n66 585
R148 VTAIL.n42 VTAIL.n41 585
R149 VTAIL.n61 VTAIL.n60 585
R150 VTAIL.n59 VTAIL.n58 585
R151 VTAIL.n46 VTAIL.n45 585
R152 VTAIL.n53 VTAIL.n52 585
R153 VTAIL.n51 VTAIL.n50 585
R154 VTAIL.n113 VTAIL.t4 329.175
R155 VTAIL.n11 VTAIL.t13 329.175
R156 VTAIL.n83 VTAIL.t17 329.175
R157 VTAIL.n49 VTAIL.t1 329.175
R158 VTAIL.n116 VTAIL.n115 171.744
R159 VTAIL.n116 VTAIL.n109 171.744
R160 VTAIL.n123 VTAIL.n109 171.744
R161 VTAIL.n124 VTAIL.n123 171.744
R162 VTAIL.n124 VTAIL.n105 171.744
R163 VTAIL.n131 VTAIL.n105 171.744
R164 VTAIL.n14 VTAIL.n13 171.744
R165 VTAIL.n14 VTAIL.n7 171.744
R166 VTAIL.n21 VTAIL.n7 171.744
R167 VTAIL.n22 VTAIL.n21 171.744
R168 VTAIL.n22 VTAIL.n3 171.744
R169 VTAIL.n29 VTAIL.n3 171.744
R170 VTAIL.n101 VTAIL.n75 171.744
R171 VTAIL.n94 VTAIL.n75 171.744
R172 VTAIL.n94 VTAIL.n93 171.744
R173 VTAIL.n93 VTAIL.n79 171.744
R174 VTAIL.n86 VTAIL.n79 171.744
R175 VTAIL.n86 VTAIL.n85 171.744
R176 VTAIL.n67 VTAIL.n41 171.744
R177 VTAIL.n60 VTAIL.n41 171.744
R178 VTAIL.n60 VTAIL.n59 171.744
R179 VTAIL.n59 VTAIL.n45 171.744
R180 VTAIL.n52 VTAIL.n45 171.744
R181 VTAIL.n52 VTAIL.n51 171.744
R182 VTAIL.n115 VTAIL.t4 85.8723
R183 VTAIL.n13 VTAIL.t13 85.8723
R184 VTAIL.n85 VTAIL.t17 85.8723
R185 VTAIL.n51 VTAIL.t1 85.8723
R186 VTAIL.n73 VTAIL.n72 78.6281
R187 VTAIL.n71 VTAIL.n70 78.6281
R188 VTAIL.n39 VTAIL.n38 78.6281
R189 VTAIL.n37 VTAIL.n36 78.6281
R190 VTAIL.n135 VTAIL.n134 78.6271
R191 VTAIL.n1 VTAIL.n0 78.6271
R192 VTAIL.n33 VTAIL.n32 78.6271
R193 VTAIL.n35 VTAIL.n34 78.6271
R194 VTAIL.n133 VTAIL.n132 34.7066
R195 VTAIL.n31 VTAIL.n30 34.7066
R196 VTAIL.n103 VTAIL.n102 34.7066
R197 VTAIL.n69 VTAIL.n68 34.7066
R198 VTAIL.n37 VTAIL.n35 21.3065
R199 VTAIL.n133 VTAIL.n103 19.3496
R200 VTAIL.n130 VTAIL.n104 12.0247
R201 VTAIL.n28 VTAIL.n2 12.0247
R202 VTAIL.n100 VTAIL.n74 12.0247
R203 VTAIL.n66 VTAIL.n40 12.0247
R204 VTAIL.n129 VTAIL.n106 11.249
R205 VTAIL.n27 VTAIL.n4 11.249
R206 VTAIL.n99 VTAIL.n76 11.249
R207 VTAIL.n65 VTAIL.n42 11.249
R208 VTAIL.n114 VTAIL.n113 10.722
R209 VTAIL.n12 VTAIL.n11 10.722
R210 VTAIL.n84 VTAIL.n83 10.722
R211 VTAIL.n50 VTAIL.n49 10.722
R212 VTAIL.n126 VTAIL.n125 10.4732
R213 VTAIL.n24 VTAIL.n23 10.4732
R214 VTAIL.n96 VTAIL.n95 10.4732
R215 VTAIL.n62 VTAIL.n61 10.4732
R216 VTAIL.n122 VTAIL.n108 9.69747
R217 VTAIL.n20 VTAIL.n6 9.69747
R218 VTAIL.n92 VTAIL.n78 9.69747
R219 VTAIL.n58 VTAIL.n44 9.69747
R220 VTAIL.n128 VTAIL.n104 9.45567
R221 VTAIL.n26 VTAIL.n2 9.45567
R222 VTAIL.n98 VTAIL.n74 9.45567
R223 VTAIL.n64 VTAIL.n40 9.45567
R224 VTAIL.n112 VTAIL.n111 9.3005
R225 VTAIL.n119 VTAIL.n118 9.3005
R226 VTAIL.n121 VTAIL.n120 9.3005
R227 VTAIL.n108 VTAIL.n107 9.3005
R228 VTAIL.n127 VTAIL.n126 9.3005
R229 VTAIL.n129 VTAIL.n128 9.3005
R230 VTAIL.n10 VTAIL.n9 9.3005
R231 VTAIL.n17 VTAIL.n16 9.3005
R232 VTAIL.n19 VTAIL.n18 9.3005
R233 VTAIL.n6 VTAIL.n5 9.3005
R234 VTAIL.n25 VTAIL.n24 9.3005
R235 VTAIL.n27 VTAIL.n26 9.3005
R236 VTAIL.n99 VTAIL.n98 9.3005
R237 VTAIL.n97 VTAIL.n96 9.3005
R238 VTAIL.n78 VTAIL.n77 9.3005
R239 VTAIL.n91 VTAIL.n90 9.3005
R240 VTAIL.n89 VTAIL.n88 9.3005
R241 VTAIL.n82 VTAIL.n81 9.3005
R242 VTAIL.n55 VTAIL.n54 9.3005
R243 VTAIL.n57 VTAIL.n56 9.3005
R244 VTAIL.n44 VTAIL.n43 9.3005
R245 VTAIL.n63 VTAIL.n62 9.3005
R246 VTAIL.n65 VTAIL.n64 9.3005
R247 VTAIL.n48 VTAIL.n47 9.3005
R248 VTAIL.n121 VTAIL.n110 8.92171
R249 VTAIL.n19 VTAIL.n8 8.92171
R250 VTAIL.n91 VTAIL.n80 8.92171
R251 VTAIL.n57 VTAIL.n46 8.92171
R252 VTAIL.n118 VTAIL.n117 8.14595
R253 VTAIL.n16 VTAIL.n15 8.14595
R254 VTAIL.n88 VTAIL.n87 8.14595
R255 VTAIL.n54 VTAIL.n53 8.14595
R256 VTAIL.n114 VTAIL.n112 7.3702
R257 VTAIL.n12 VTAIL.n10 7.3702
R258 VTAIL.n84 VTAIL.n82 7.3702
R259 VTAIL.n50 VTAIL.n48 7.3702
R260 VTAIL.n117 VTAIL.n112 5.81868
R261 VTAIL.n15 VTAIL.n10 5.81868
R262 VTAIL.n87 VTAIL.n82 5.81868
R263 VTAIL.n53 VTAIL.n48 5.81868
R264 VTAIL.n134 VTAIL.t7 5.57597
R265 VTAIL.n134 VTAIL.t0 5.57597
R266 VTAIL.n0 VTAIL.t6 5.57597
R267 VTAIL.n0 VTAIL.t5 5.57597
R268 VTAIL.n32 VTAIL.t16 5.57597
R269 VTAIL.n32 VTAIL.t15 5.57597
R270 VTAIL.n34 VTAIL.t11 5.57597
R271 VTAIL.n34 VTAIL.t14 5.57597
R272 VTAIL.n72 VTAIL.t18 5.57597
R273 VTAIL.n72 VTAIL.t9 5.57597
R274 VTAIL.n70 VTAIL.t12 5.57597
R275 VTAIL.n70 VTAIL.t10 5.57597
R276 VTAIL.n38 VTAIL.t2 5.57597
R277 VTAIL.n38 VTAIL.t3 5.57597
R278 VTAIL.n36 VTAIL.t19 5.57597
R279 VTAIL.n36 VTAIL.t8 5.57597
R280 VTAIL.n118 VTAIL.n110 5.04292
R281 VTAIL.n16 VTAIL.n8 5.04292
R282 VTAIL.n88 VTAIL.n80 5.04292
R283 VTAIL.n54 VTAIL.n46 5.04292
R284 VTAIL.n122 VTAIL.n121 4.26717
R285 VTAIL.n20 VTAIL.n19 4.26717
R286 VTAIL.n92 VTAIL.n91 4.26717
R287 VTAIL.n58 VTAIL.n57 4.26717
R288 VTAIL.n125 VTAIL.n108 3.49141
R289 VTAIL.n23 VTAIL.n6 3.49141
R290 VTAIL.n95 VTAIL.n78 3.49141
R291 VTAIL.n61 VTAIL.n44 3.49141
R292 VTAIL.n126 VTAIL.n106 2.71565
R293 VTAIL.n24 VTAIL.n4 2.71565
R294 VTAIL.n96 VTAIL.n76 2.71565
R295 VTAIL.n62 VTAIL.n42 2.71565
R296 VTAIL.n113 VTAIL.n111 2.4147
R297 VTAIL.n11 VTAIL.n9 2.4147
R298 VTAIL.n83 VTAIL.n81 2.4147
R299 VTAIL.n49 VTAIL.n47 2.4147
R300 VTAIL.n39 VTAIL.n37 1.9574
R301 VTAIL.n69 VTAIL.n39 1.9574
R302 VTAIL.n73 VTAIL.n71 1.9574
R303 VTAIL.n103 VTAIL.n73 1.9574
R304 VTAIL.n35 VTAIL.n33 1.9574
R305 VTAIL.n33 VTAIL.n31 1.9574
R306 VTAIL.n135 VTAIL.n133 1.9574
R307 VTAIL.n130 VTAIL.n129 1.93989
R308 VTAIL.n28 VTAIL.n27 1.93989
R309 VTAIL.n100 VTAIL.n99 1.93989
R310 VTAIL.n66 VTAIL.n65 1.93989
R311 VTAIL VTAIL.n1 1.52636
R312 VTAIL.n71 VTAIL.n69 1.44878
R313 VTAIL.n31 VTAIL.n1 1.44878
R314 VTAIL.n132 VTAIL.n104 1.16414
R315 VTAIL.n30 VTAIL.n2 1.16414
R316 VTAIL.n102 VTAIL.n74 1.16414
R317 VTAIL.n68 VTAIL.n40 1.16414
R318 VTAIL VTAIL.n135 0.431534
R319 VTAIL.n119 VTAIL.n111 0.155672
R320 VTAIL.n120 VTAIL.n119 0.155672
R321 VTAIL.n120 VTAIL.n107 0.155672
R322 VTAIL.n127 VTAIL.n107 0.155672
R323 VTAIL.n128 VTAIL.n127 0.155672
R324 VTAIL.n17 VTAIL.n9 0.155672
R325 VTAIL.n18 VTAIL.n17 0.155672
R326 VTAIL.n18 VTAIL.n5 0.155672
R327 VTAIL.n25 VTAIL.n5 0.155672
R328 VTAIL.n26 VTAIL.n25 0.155672
R329 VTAIL.n98 VTAIL.n97 0.155672
R330 VTAIL.n97 VTAIL.n77 0.155672
R331 VTAIL.n90 VTAIL.n77 0.155672
R332 VTAIL.n90 VTAIL.n89 0.155672
R333 VTAIL.n89 VTAIL.n81 0.155672
R334 VTAIL.n64 VTAIL.n63 0.155672
R335 VTAIL.n63 VTAIL.n43 0.155672
R336 VTAIL.n56 VTAIL.n43 0.155672
R337 VTAIL.n56 VTAIL.n55 0.155672
R338 VTAIL.n55 VTAIL.n47 0.155672
R339 VDD1.n28 VDD1.n27 756.745
R340 VDD1.n59 VDD1.n58 756.745
R341 VDD1.n27 VDD1.n26 585
R342 VDD1.n2 VDD1.n1 585
R343 VDD1.n21 VDD1.n20 585
R344 VDD1.n19 VDD1.n18 585
R345 VDD1.n6 VDD1.n5 585
R346 VDD1.n13 VDD1.n12 585
R347 VDD1.n11 VDD1.n10 585
R348 VDD1.n42 VDD1.n41 585
R349 VDD1.n44 VDD1.n43 585
R350 VDD1.n37 VDD1.n36 585
R351 VDD1.n50 VDD1.n49 585
R352 VDD1.n52 VDD1.n51 585
R353 VDD1.n33 VDD1.n32 585
R354 VDD1.n58 VDD1.n57 585
R355 VDD1.n40 VDD1.t9 329.175
R356 VDD1.n9 VDD1.t8 329.175
R357 VDD1.n27 VDD1.n1 171.744
R358 VDD1.n20 VDD1.n1 171.744
R359 VDD1.n20 VDD1.n19 171.744
R360 VDD1.n19 VDD1.n5 171.744
R361 VDD1.n12 VDD1.n5 171.744
R362 VDD1.n12 VDD1.n11 171.744
R363 VDD1.n43 VDD1.n42 171.744
R364 VDD1.n43 VDD1.n36 171.744
R365 VDD1.n50 VDD1.n36 171.744
R366 VDD1.n51 VDD1.n50 171.744
R367 VDD1.n51 VDD1.n32 171.744
R368 VDD1.n58 VDD1.n32 171.744
R369 VDD1.n63 VDD1.n62 96.7182
R370 VDD1.n30 VDD1.n29 95.3069
R371 VDD1.n61 VDD1.n60 95.3059
R372 VDD1.n65 VDD1.n64 95.3057
R373 VDD1.n11 VDD1.t8 85.8723
R374 VDD1.n42 VDD1.t9 85.8723
R375 VDD1.n30 VDD1.n28 53.3422
R376 VDD1.n61 VDD1.n59 53.3422
R377 VDD1.n65 VDD1.n63 39.5979
R378 VDD1.n26 VDD1.n0 12.0247
R379 VDD1.n57 VDD1.n31 12.0247
R380 VDD1.n25 VDD1.n2 11.249
R381 VDD1.n56 VDD1.n33 11.249
R382 VDD1.n41 VDD1.n40 10.722
R383 VDD1.n10 VDD1.n9 10.722
R384 VDD1.n22 VDD1.n21 10.4732
R385 VDD1.n53 VDD1.n52 10.4732
R386 VDD1.n18 VDD1.n4 9.69747
R387 VDD1.n49 VDD1.n35 9.69747
R388 VDD1.n24 VDD1.n0 9.45567
R389 VDD1.n55 VDD1.n31 9.45567
R390 VDD1.n15 VDD1.n14 9.3005
R391 VDD1.n17 VDD1.n16 9.3005
R392 VDD1.n4 VDD1.n3 9.3005
R393 VDD1.n23 VDD1.n22 9.3005
R394 VDD1.n25 VDD1.n24 9.3005
R395 VDD1.n8 VDD1.n7 9.3005
R396 VDD1.n39 VDD1.n38 9.3005
R397 VDD1.n46 VDD1.n45 9.3005
R398 VDD1.n48 VDD1.n47 9.3005
R399 VDD1.n35 VDD1.n34 9.3005
R400 VDD1.n54 VDD1.n53 9.3005
R401 VDD1.n56 VDD1.n55 9.3005
R402 VDD1.n17 VDD1.n6 8.92171
R403 VDD1.n48 VDD1.n37 8.92171
R404 VDD1.n14 VDD1.n13 8.14595
R405 VDD1.n45 VDD1.n44 8.14595
R406 VDD1.n10 VDD1.n8 7.3702
R407 VDD1.n41 VDD1.n39 7.3702
R408 VDD1.n13 VDD1.n8 5.81868
R409 VDD1.n44 VDD1.n39 5.81868
R410 VDD1.n64 VDD1.t1 5.57597
R411 VDD1.n64 VDD1.t6 5.57597
R412 VDD1.n29 VDD1.t4 5.57597
R413 VDD1.n29 VDD1.t3 5.57597
R414 VDD1.n62 VDD1.t7 5.57597
R415 VDD1.n62 VDD1.t0 5.57597
R416 VDD1.n60 VDD1.t2 5.57597
R417 VDD1.n60 VDD1.t5 5.57597
R418 VDD1.n14 VDD1.n6 5.04292
R419 VDD1.n45 VDD1.n37 5.04292
R420 VDD1.n18 VDD1.n17 4.26717
R421 VDD1.n49 VDD1.n48 4.26717
R422 VDD1.n21 VDD1.n4 3.49141
R423 VDD1.n52 VDD1.n35 3.49141
R424 VDD1.n22 VDD1.n2 2.71565
R425 VDD1.n53 VDD1.n33 2.71565
R426 VDD1.n40 VDD1.n38 2.4147
R427 VDD1.n9 VDD1.n7 2.4147
R428 VDD1.n26 VDD1.n25 1.93989
R429 VDD1.n57 VDD1.n56 1.93989
R430 VDD1 VDD1.n65 1.40998
R431 VDD1.n28 VDD1.n0 1.16414
R432 VDD1.n59 VDD1.n31 1.16414
R433 VDD1 VDD1.n30 0.547914
R434 VDD1.n63 VDD1.n61 0.434378
R435 VDD1.n24 VDD1.n23 0.155672
R436 VDD1.n23 VDD1.n3 0.155672
R437 VDD1.n16 VDD1.n3 0.155672
R438 VDD1.n16 VDD1.n15 0.155672
R439 VDD1.n15 VDD1.n7 0.155672
R440 VDD1.n46 VDD1.n38 0.155672
R441 VDD1.n47 VDD1.n46 0.155672
R442 VDD1.n47 VDD1.n34 0.155672
R443 VDD1.n54 VDD1.n34 0.155672
R444 VDD1.n55 VDD1.n54 0.155672
R445 B.n466 B.n465 585
R446 B.n467 B.n58 585
R447 B.n469 B.n468 585
R448 B.n470 B.n57 585
R449 B.n472 B.n471 585
R450 B.n473 B.n56 585
R451 B.n475 B.n474 585
R452 B.n476 B.n55 585
R453 B.n478 B.n477 585
R454 B.n479 B.n54 585
R455 B.n481 B.n480 585
R456 B.n482 B.n53 585
R457 B.n484 B.n483 585
R458 B.n485 B.n52 585
R459 B.n487 B.n486 585
R460 B.n488 B.n51 585
R461 B.n490 B.n489 585
R462 B.n491 B.n50 585
R463 B.n493 B.n492 585
R464 B.n494 B.n49 585
R465 B.n496 B.n495 585
R466 B.n497 B.n45 585
R467 B.n499 B.n498 585
R468 B.n500 B.n44 585
R469 B.n502 B.n501 585
R470 B.n503 B.n43 585
R471 B.n505 B.n504 585
R472 B.n506 B.n42 585
R473 B.n508 B.n507 585
R474 B.n509 B.n41 585
R475 B.n511 B.n510 585
R476 B.n512 B.n40 585
R477 B.n514 B.n513 585
R478 B.n516 B.n37 585
R479 B.n518 B.n517 585
R480 B.n519 B.n36 585
R481 B.n521 B.n520 585
R482 B.n522 B.n35 585
R483 B.n524 B.n523 585
R484 B.n525 B.n34 585
R485 B.n527 B.n526 585
R486 B.n528 B.n33 585
R487 B.n530 B.n529 585
R488 B.n531 B.n32 585
R489 B.n533 B.n532 585
R490 B.n534 B.n31 585
R491 B.n536 B.n535 585
R492 B.n537 B.n30 585
R493 B.n539 B.n538 585
R494 B.n540 B.n29 585
R495 B.n542 B.n541 585
R496 B.n543 B.n28 585
R497 B.n545 B.n544 585
R498 B.n546 B.n27 585
R499 B.n548 B.n547 585
R500 B.n549 B.n26 585
R501 B.n464 B.n59 585
R502 B.n463 B.n462 585
R503 B.n461 B.n60 585
R504 B.n460 B.n459 585
R505 B.n458 B.n61 585
R506 B.n457 B.n456 585
R507 B.n455 B.n62 585
R508 B.n454 B.n453 585
R509 B.n452 B.n63 585
R510 B.n451 B.n450 585
R511 B.n449 B.n64 585
R512 B.n448 B.n447 585
R513 B.n446 B.n65 585
R514 B.n445 B.n444 585
R515 B.n443 B.n66 585
R516 B.n442 B.n441 585
R517 B.n440 B.n67 585
R518 B.n439 B.n438 585
R519 B.n437 B.n68 585
R520 B.n436 B.n435 585
R521 B.n434 B.n69 585
R522 B.n433 B.n432 585
R523 B.n431 B.n70 585
R524 B.n430 B.n429 585
R525 B.n428 B.n71 585
R526 B.n427 B.n426 585
R527 B.n425 B.n72 585
R528 B.n424 B.n423 585
R529 B.n422 B.n73 585
R530 B.n421 B.n420 585
R531 B.n419 B.n74 585
R532 B.n418 B.n417 585
R533 B.n416 B.n75 585
R534 B.n415 B.n414 585
R535 B.n413 B.n76 585
R536 B.n412 B.n411 585
R537 B.n410 B.n77 585
R538 B.n409 B.n408 585
R539 B.n407 B.n78 585
R540 B.n406 B.n405 585
R541 B.n404 B.n79 585
R542 B.n403 B.n402 585
R543 B.n401 B.n80 585
R544 B.n400 B.n399 585
R545 B.n398 B.n81 585
R546 B.n397 B.n396 585
R547 B.n395 B.n82 585
R548 B.n394 B.n393 585
R549 B.n392 B.n83 585
R550 B.n391 B.n390 585
R551 B.n389 B.n84 585
R552 B.n388 B.n387 585
R553 B.n386 B.n85 585
R554 B.n385 B.n384 585
R555 B.n383 B.n86 585
R556 B.n382 B.n381 585
R557 B.n380 B.n87 585
R558 B.n379 B.n378 585
R559 B.n377 B.n88 585
R560 B.n376 B.n375 585
R561 B.n374 B.n89 585
R562 B.n373 B.n372 585
R563 B.n371 B.n90 585
R564 B.n370 B.n369 585
R565 B.n368 B.n91 585
R566 B.n367 B.n366 585
R567 B.n365 B.n92 585
R568 B.n364 B.n363 585
R569 B.n362 B.n93 585
R570 B.n361 B.n360 585
R571 B.n359 B.n94 585
R572 B.n358 B.n357 585
R573 B.n356 B.n95 585
R574 B.n355 B.n354 585
R575 B.n353 B.n96 585
R576 B.n352 B.n351 585
R577 B.n350 B.n97 585
R578 B.n349 B.n348 585
R579 B.n347 B.n98 585
R580 B.n346 B.n345 585
R581 B.n344 B.n99 585
R582 B.n343 B.n342 585
R583 B.n341 B.n100 585
R584 B.n340 B.n339 585
R585 B.n338 B.n101 585
R586 B.n337 B.n336 585
R587 B.n335 B.n102 585
R588 B.n334 B.n333 585
R589 B.n332 B.n103 585
R590 B.n331 B.n330 585
R591 B.n329 B.n104 585
R592 B.n328 B.n327 585
R593 B.n326 B.n105 585
R594 B.n325 B.n324 585
R595 B.n323 B.n106 585
R596 B.n322 B.n321 585
R597 B.n320 B.n107 585
R598 B.n235 B.n234 585
R599 B.n236 B.n139 585
R600 B.n238 B.n237 585
R601 B.n239 B.n138 585
R602 B.n241 B.n240 585
R603 B.n242 B.n137 585
R604 B.n244 B.n243 585
R605 B.n245 B.n136 585
R606 B.n247 B.n246 585
R607 B.n248 B.n135 585
R608 B.n250 B.n249 585
R609 B.n251 B.n134 585
R610 B.n253 B.n252 585
R611 B.n254 B.n133 585
R612 B.n256 B.n255 585
R613 B.n257 B.n132 585
R614 B.n259 B.n258 585
R615 B.n260 B.n131 585
R616 B.n262 B.n261 585
R617 B.n263 B.n130 585
R618 B.n265 B.n264 585
R619 B.n266 B.n129 585
R620 B.n268 B.n267 585
R621 B.n270 B.n126 585
R622 B.n272 B.n271 585
R623 B.n273 B.n125 585
R624 B.n275 B.n274 585
R625 B.n276 B.n124 585
R626 B.n278 B.n277 585
R627 B.n279 B.n123 585
R628 B.n281 B.n280 585
R629 B.n282 B.n122 585
R630 B.n284 B.n283 585
R631 B.n286 B.n285 585
R632 B.n287 B.n118 585
R633 B.n289 B.n288 585
R634 B.n290 B.n117 585
R635 B.n292 B.n291 585
R636 B.n293 B.n116 585
R637 B.n295 B.n294 585
R638 B.n296 B.n115 585
R639 B.n298 B.n297 585
R640 B.n299 B.n114 585
R641 B.n301 B.n300 585
R642 B.n302 B.n113 585
R643 B.n304 B.n303 585
R644 B.n305 B.n112 585
R645 B.n307 B.n306 585
R646 B.n308 B.n111 585
R647 B.n310 B.n309 585
R648 B.n311 B.n110 585
R649 B.n313 B.n312 585
R650 B.n314 B.n109 585
R651 B.n316 B.n315 585
R652 B.n317 B.n108 585
R653 B.n319 B.n318 585
R654 B.n233 B.n140 585
R655 B.n232 B.n231 585
R656 B.n230 B.n141 585
R657 B.n229 B.n228 585
R658 B.n227 B.n142 585
R659 B.n226 B.n225 585
R660 B.n224 B.n143 585
R661 B.n223 B.n222 585
R662 B.n221 B.n144 585
R663 B.n220 B.n219 585
R664 B.n218 B.n145 585
R665 B.n217 B.n216 585
R666 B.n215 B.n146 585
R667 B.n214 B.n213 585
R668 B.n212 B.n147 585
R669 B.n211 B.n210 585
R670 B.n209 B.n148 585
R671 B.n208 B.n207 585
R672 B.n206 B.n149 585
R673 B.n205 B.n204 585
R674 B.n203 B.n150 585
R675 B.n202 B.n201 585
R676 B.n200 B.n151 585
R677 B.n199 B.n198 585
R678 B.n197 B.n152 585
R679 B.n196 B.n195 585
R680 B.n194 B.n153 585
R681 B.n193 B.n192 585
R682 B.n191 B.n154 585
R683 B.n190 B.n189 585
R684 B.n188 B.n155 585
R685 B.n187 B.n186 585
R686 B.n185 B.n156 585
R687 B.n184 B.n183 585
R688 B.n182 B.n157 585
R689 B.n181 B.n180 585
R690 B.n179 B.n158 585
R691 B.n178 B.n177 585
R692 B.n176 B.n159 585
R693 B.n175 B.n174 585
R694 B.n173 B.n160 585
R695 B.n172 B.n171 585
R696 B.n170 B.n161 585
R697 B.n169 B.n168 585
R698 B.n167 B.n162 585
R699 B.n166 B.n165 585
R700 B.n164 B.n163 585
R701 B.n2 B.n0 585
R702 B.n621 B.n1 585
R703 B.n620 B.n619 585
R704 B.n618 B.n3 585
R705 B.n617 B.n616 585
R706 B.n615 B.n4 585
R707 B.n614 B.n613 585
R708 B.n612 B.n5 585
R709 B.n611 B.n610 585
R710 B.n609 B.n6 585
R711 B.n608 B.n607 585
R712 B.n606 B.n7 585
R713 B.n605 B.n604 585
R714 B.n603 B.n8 585
R715 B.n602 B.n601 585
R716 B.n600 B.n9 585
R717 B.n599 B.n598 585
R718 B.n597 B.n10 585
R719 B.n596 B.n595 585
R720 B.n594 B.n11 585
R721 B.n593 B.n592 585
R722 B.n591 B.n12 585
R723 B.n590 B.n589 585
R724 B.n588 B.n13 585
R725 B.n587 B.n586 585
R726 B.n585 B.n14 585
R727 B.n584 B.n583 585
R728 B.n582 B.n15 585
R729 B.n581 B.n580 585
R730 B.n579 B.n16 585
R731 B.n578 B.n577 585
R732 B.n576 B.n17 585
R733 B.n575 B.n574 585
R734 B.n573 B.n18 585
R735 B.n572 B.n571 585
R736 B.n570 B.n19 585
R737 B.n569 B.n568 585
R738 B.n567 B.n20 585
R739 B.n566 B.n565 585
R740 B.n564 B.n21 585
R741 B.n563 B.n562 585
R742 B.n561 B.n22 585
R743 B.n560 B.n559 585
R744 B.n558 B.n23 585
R745 B.n557 B.n556 585
R746 B.n555 B.n24 585
R747 B.n554 B.n553 585
R748 B.n552 B.n25 585
R749 B.n551 B.n550 585
R750 B.n623 B.n622 585
R751 B.n235 B.n140 569.379
R752 B.n550 B.n549 569.379
R753 B.n320 B.n319 569.379
R754 B.n465 B.n464 569.379
R755 B.n119 B.t11 308.921
R756 B.n46 B.t7 308.921
R757 B.n127 B.t5 308.921
R758 B.n38 B.t1 308.921
R759 B.n119 B.t9 279.197
R760 B.n127 B.t3 279.197
R761 B.n38 B.t0 279.197
R762 B.n46 B.t6 279.197
R763 B.n120 B.t10 264.897
R764 B.n47 B.t8 264.897
R765 B.n128 B.t4 264.896
R766 B.n39 B.t2 264.896
R767 B.n231 B.n140 163.367
R768 B.n231 B.n230 163.367
R769 B.n230 B.n229 163.367
R770 B.n229 B.n142 163.367
R771 B.n225 B.n142 163.367
R772 B.n225 B.n224 163.367
R773 B.n224 B.n223 163.367
R774 B.n223 B.n144 163.367
R775 B.n219 B.n144 163.367
R776 B.n219 B.n218 163.367
R777 B.n218 B.n217 163.367
R778 B.n217 B.n146 163.367
R779 B.n213 B.n146 163.367
R780 B.n213 B.n212 163.367
R781 B.n212 B.n211 163.367
R782 B.n211 B.n148 163.367
R783 B.n207 B.n148 163.367
R784 B.n207 B.n206 163.367
R785 B.n206 B.n205 163.367
R786 B.n205 B.n150 163.367
R787 B.n201 B.n150 163.367
R788 B.n201 B.n200 163.367
R789 B.n200 B.n199 163.367
R790 B.n199 B.n152 163.367
R791 B.n195 B.n152 163.367
R792 B.n195 B.n194 163.367
R793 B.n194 B.n193 163.367
R794 B.n193 B.n154 163.367
R795 B.n189 B.n154 163.367
R796 B.n189 B.n188 163.367
R797 B.n188 B.n187 163.367
R798 B.n187 B.n156 163.367
R799 B.n183 B.n156 163.367
R800 B.n183 B.n182 163.367
R801 B.n182 B.n181 163.367
R802 B.n181 B.n158 163.367
R803 B.n177 B.n158 163.367
R804 B.n177 B.n176 163.367
R805 B.n176 B.n175 163.367
R806 B.n175 B.n160 163.367
R807 B.n171 B.n160 163.367
R808 B.n171 B.n170 163.367
R809 B.n170 B.n169 163.367
R810 B.n169 B.n162 163.367
R811 B.n165 B.n162 163.367
R812 B.n165 B.n164 163.367
R813 B.n164 B.n2 163.367
R814 B.n622 B.n2 163.367
R815 B.n622 B.n621 163.367
R816 B.n621 B.n620 163.367
R817 B.n620 B.n3 163.367
R818 B.n616 B.n3 163.367
R819 B.n616 B.n615 163.367
R820 B.n615 B.n614 163.367
R821 B.n614 B.n5 163.367
R822 B.n610 B.n5 163.367
R823 B.n610 B.n609 163.367
R824 B.n609 B.n608 163.367
R825 B.n608 B.n7 163.367
R826 B.n604 B.n7 163.367
R827 B.n604 B.n603 163.367
R828 B.n603 B.n602 163.367
R829 B.n602 B.n9 163.367
R830 B.n598 B.n9 163.367
R831 B.n598 B.n597 163.367
R832 B.n597 B.n596 163.367
R833 B.n596 B.n11 163.367
R834 B.n592 B.n11 163.367
R835 B.n592 B.n591 163.367
R836 B.n591 B.n590 163.367
R837 B.n590 B.n13 163.367
R838 B.n586 B.n13 163.367
R839 B.n586 B.n585 163.367
R840 B.n585 B.n584 163.367
R841 B.n584 B.n15 163.367
R842 B.n580 B.n15 163.367
R843 B.n580 B.n579 163.367
R844 B.n579 B.n578 163.367
R845 B.n578 B.n17 163.367
R846 B.n574 B.n17 163.367
R847 B.n574 B.n573 163.367
R848 B.n573 B.n572 163.367
R849 B.n572 B.n19 163.367
R850 B.n568 B.n19 163.367
R851 B.n568 B.n567 163.367
R852 B.n567 B.n566 163.367
R853 B.n566 B.n21 163.367
R854 B.n562 B.n21 163.367
R855 B.n562 B.n561 163.367
R856 B.n561 B.n560 163.367
R857 B.n560 B.n23 163.367
R858 B.n556 B.n23 163.367
R859 B.n556 B.n555 163.367
R860 B.n555 B.n554 163.367
R861 B.n554 B.n25 163.367
R862 B.n550 B.n25 163.367
R863 B.n236 B.n235 163.367
R864 B.n237 B.n236 163.367
R865 B.n237 B.n138 163.367
R866 B.n241 B.n138 163.367
R867 B.n242 B.n241 163.367
R868 B.n243 B.n242 163.367
R869 B.n243 B.n136 163.367
R870 B.n247 B.n136 163.367
R871 B.n248 B.n247 163.367
R872 B.n249 B.n248 163.367
R873 B.n249 B.n134 163.367
R874 B.n253 B.n134 163.367
R875 B.n254 B.n253 163.367
R876 B.n255 B.n254 163.367
R877 B.n255 B.n132 163.367
R878 B.n259 B.n132 163.367
R879 B.n260 B.n259 163.367
R880 B.n261 B.n260 163.367
R881 B.n261 B.n130 163.367
R882 B.n265 B.n130 163.367
R883 B.n266 B.n265 163.367
R884 B.n267 B.n266 163.367
R885 B.n267 B.n126 163.367
R886 B.n272 B.n126 163.367
R887 B.n273 B.n272 163.367
R888 B.n274 B.n273 163.367
R889 B.n274 B.n124 163.367
R890 B.n278 B.n124 163.367
R891 B.n279 B.n278 163.367
R892 B.n280 B.n279 163.367
R893 B.n280 B.n122 163.367
R894 B.n284 B.n122 163.367
R895 B.n285 B.n284 163.367
R896 B.n285 B.n118 163.367
R897 B.n289 B.n118 163.367
R898 B.n290 B.n289 163.367
R899 B.n291 B.n290 163.367
R900 B.n291 B.n116 163.367
R901 B.n295 B.n116 163.367
R902 B.n296 B.n295 163.367
R903 B.n297 B.n296 163.367
R904 B.n297 B.n114 163.367
R905 B.n301 B.n114 163.367
R906 B.n302 B.n301 163.367
R907 B.n303 B.n302 163.367
R908 B.n303 B.n112 163.367
R909 B.n307 B.n112 163.367
R910 B.n308 B.n307 163.367
R911 B.n309 B.n308 163.367
R912 B.n309 B.n110 163.367
R913 B.n313 B.n110 163.367
R914 B.n314 B.n313 163.367
R915 B.n315 B.n314 163.367
R916 B.n315 B.n108 163.367
R917 B.n319 B.n108 163.367
R918 B.n321 B.n320 163.367
R919 B.n321 B.n106 163.367
R920 B.n325 B.n106 163.367
R921 B.n326 B.n325 163.367
R922 B.n327 B.n326 163.367
R923 B.n327 B.n104 163.367
R924 B.n331 B.n104 163.367
R925 B.n332 B.n331 163.367
R926 B.n333 B.n332 163.367
R927 B.n333 B.n102 163.367
R928 B.n337 B.n102 163.367
R929 B.n338 B.n337 163.367
R930 B.n339 B.n338 163.367
R931 B.n339 B.n100 163.367
R932 B.n343 B.n100 163.367
R933 B.n344 B.n343 163.367
R934 B.n345 B.n344 163.367
R935 B.n345 B.n98 163.367
R936 B.n349 B.n98 163.367
R937 B.n350 B.n349 163.367
R938 B.n351 B.n350 163.367
R939 B.n351 B.n96 163.367
R940 B.n355 B.n96 163.367
R941 B.n356 B.n355 163.367
R942 B.n357 B.n356 163.367
R943 B.n357 B.n94 163.367
R944 B.n361 B.n94 163.367
R945 B.n362 B.n361 163.367
R946 B.n363 B.n362 163.367
R947 B.n363 B.n92 163.367
R948 B.n367 B.n92 163.367
R949 B.n368 B.n367 163.367
R950 B.n369 B.n368 163.367
R951 B.n369 B.n90 163.367
R952 B.n373 B.n90 163.367
R953 B.n374 B.n373 163.367
R954 B.n375 B.n374 163.367
R955 B.n375 B.n88 163.367
R956 B.n379 B.n88 163.367
R957 B.n380 B.n379 163.367
R958 B.n381 B.n380 163.367
R959 B.n381 B.n86 163.367
R960 B.n385 B.n86 163.367
R961 B.n386 B.n385 163.367
R962 B.n387 B.n386 163.367
R963 B.n387 B.n84 163.367
R964 B.n391 B.n84 163.367
R965 B.n392 B.n391 163.367
R966 B.n393 B.n392 163.367
R967 B.n393 B.n82 163.367
R968 B.n397 B.n82 163.367
R969 B.n398 B.n397 163.367
R970 B.n399 B.n398 163.367
R971 B.n399 B.n80 163.367
R972 B.n403 B.n80 163.367
R973 B.n404 B.n403 163.367
R974 B.n405 B.n404 163.367
R975 B.n405 B.n78 163.367
R976 B.n409 B.n78 163.367
R977 B.n410 B.n409 163.367
R978 B.n411 B.n410 163.367
R979 B.n411 B.n76 163.367
R980 B.n415 B.n76 163.367
R981 B.n416 B.n415 163.367
R982 B.n417 B.n416 163.367
R983 B.n417 B.n74 163.367
R984 B.n421 B.n74 163.367
R985 B.n422 B.n421 163.367
R986 B.n423 B.n422 163.367
R987 B.n423 B.n72 163.367
R988 B.n427 B.n72 163.367
R989 B.n428 B.n427 163.367
R990 B.n429 B.n428 163.367
R991 B.n429 B.n70 163.367
R992 B.n433 B.n70 163.367
R993 B.n434 B.n433 163.367
R994 B.n435 B.n434 163.367
R995 B.n435 B.n68 163.367
R996 B.n439 B.n68 163.367
R997 B.n440 B.n439 163.367
R998 B.n441 B.n440 163.367
R999 B.n441 B.n66 163.367
R1000 B.n445 B.n66 163.367
R1001 B.n446 B.n445 163.367
R1002 B.n447 B.n446 163.367
R1003 B.n447 B.n64 163.367
R1004 B.n451 B.n64 163.367
R1005 B.n452 B.n451 163.367
R1006 B.n453 B.n452 163.367
R1007 B.n453 B.n62 163.367
R1008 B.n457 B.n62 163.367
R1009 B.n458 B.n457 163.367
R1010 B.n459 B.n458 163.367
R1011 B.n459 B.n60 163.367
R1012 B.n463 B.n60 163.367
R1013 B.n464 B.n463 163.367
R1014 B.n549 B.n548 163.367
R1015 B.n548 B.n27 163.367
R1016 B.n544 B.n27 163.367
R1017 B.n544 B.n543 163.367
R1018 B.n543 B.n542 163.367
R1019 B.n542 B.n29 163.367
R1020 B.n538 B.n29 163.367
R1021 B.n538 B.n537 163.367
R1022 B.n537 B.n536 163.367
R1023 B.n536 B.n31 163.367
R1024 B.n532 B.n31 163.367
R1025 B.n532 B.n531 163.367
R1026 B.n531 B.n530 163.367
R1027 B.n530 B.n33 163.367
R1028 B.n526 B.n33 163.367
R1029 B.n526 B.n525 163.367
R1030 B.n525 B.n524 163.367
R1031 B.n524 B.n35 163.367
R1032 B.n520 B.n35 163.367
R1033 B.n520 B.n519 163.367
R1034 B.n519 B.n518 163.367
R1035 B.n518 B.n37 163.367
R1036 B.n513 B.n37 163.367
R1037 B.n513 B.n512 163.367
R1038 B.n512 B.n511 163.367
R1039 B.n511 B.n41 163.367
R1040 B.n507 B.n41 163.367
R1041 B.n507 B.n506 163.367
R1042 B.n506 B.n505 163.367
R1043 B.n505 B.n43 163.367
R1044 B.n501 B.n43 163.367
R1045 B.n501 B.n500 163.367
R1046 B.n500 B.n499 163.367
R1047 B.n499 B.n45 163.367
R1048 B.n495 B.n45 163.367
R1049 B.n495 B.n494 163.367
R1050 B.n494 B.n493 163.367
R1051 B.n493 B.n50 163.367
R1052 B.n489 B.n50 163.367
R1053 B.n489 B.n488 163.367
R1054 B.n488 B.n487 163.367
R1055 B.n487 B.n52 163.367
R1056 B.n483 B.n52 163.367
R1057 B.n483 B.n482 163.367
R1058 B.n482 B.n481 163.367
R1059 B.n481 B.n54 163.367
R1060 B.n477 B.n54 163.367
R1061 B.n477 B.n476 163.367
R1062 B.n476 B.n475 163.367
R1063 B.n475 B.n56 163.367
R1064 B.n471 B.n56 163.367
R1065 B.n471 B.n470 163.367
R1066 B.n470 B.n469 163.367
R1067 B.n469 B.n58 163.367
R1068 B.n465 B.n58 163.367
R1069 B.n121 B.n120 59.5399
R1070 B.n269 B.n128 59.5399
R1071 B.n515 B.n39 59.5399
R1072 B.n48 B.n47 59.5399
R1073 B.n120 B.n119 44.0247
R1074 B.n128 B.n127 44.0247
R1075 B.n39 B.n38 44.0247
R1076 B.n47 B.n46 44.0247
R1077 B.n551 B.n26 36.9956
R1078 B.n466 B.n59 36.9956
R1079 B.n318 B.n107 36.9956
R1080 B.n234 B.n233 36.9956
R1081 B B.n623 18.0485
R1082 B.n547 B.n26 10.6151
R1083 B.n547 B.n546 10.6151
R1084 B.n546 B.n545 10.6151
R1085 B.n545 B.n28 10.6151
R1086 B.n541 B.n28 10.6151
R1087 B.n541 B.n540 10.6151
R1088 B.n540 B.n539 10.6151
R1089 B.n539 B.n30 10.6151
R1090 B.n535 B.n30 10.6151
R1091 B.n535 B.n534 10.6151
R1092 B.n534 B.n533 10.6151
R1093 B.n533 B.n32 10.6151
R1094 B.n529 B.n32 10.6151
R1095 B.n529 B.n528 10.6151
R1096 B.n528 B.n527 10.6151
R1097 B.n527 B.n34 10.6151
R1098 B.n523 B.n34 10.6151
R1099 B.n523 B.n522 10.6151
R1100 B.n522 B.n521 10.6151
R1101 B.n521 B.n36 10.6151
R1102 B.n517 B.n36 10.6151
R1103 B.n517 B.n516 10.6151
R1104 B.n514 B.n40 10.6151
R1105 B.n510 B.n40 10.6151
R1106 B.n510 B.n509 10.6151
R1107 B.n509 B.n508 10.6151
R1108 B.n508 B.n42 10.6151
R1109 B.n504 B.n42 10.6151
R1110 B.n504 B.n503 10.6151
R1111 B.n503 B.n502 10.6151
R1112 B.n502 B.n44 10.6151
R1113 B.n498 B.n497 10.6151
R1114 B.n497 B.n496 10.6151
R1115 B.n496 B.n49 10.6151
R1116 B.n492 B.n49 10.6151
R1117 B.n492 B.n491 10.6151
R1118 B.n491 B.n490 10.6151
R1119 B.n490 B.n51 10.6151
R1120 B.n486 B.n51 10.6151
R1121 B.n486 B.n485 10.6151
R1122 B.n485 B.n484 10.6151
R1123 B.n484 B.n53 10.6151
R1124 B.n480 B.n53 10.6151
R1125 B.n480 B.n479 10.6151
R1126 B.n479 B.n478 10.6151
R1127 B.n478 B.n55 10.6151
R1128 B.n474 B.n55 10.6151
R1129 B.n474 B.n473 10.6151
R1130 B.n473 B.n472 10.6151
R1131 B.n472 B.n57 10.6151
R1132 B.n468 B.n57 10.6151
R1133 B.n468 B.n467 10.6151
R1134 B.n467 B.n466 10.6151
R1135 B.n322 B.n107 10.6151
R1136 B.n323 B.n322 10.6151
R1137 B.n324 B.n323 10.6151
R1138 B.n324 B.n105 10.6151
R1139 B.n328 B.n105 10.6151
R1140 B.n329 B.n328 10.6151
R1141 B.n330 B.n329 10.6151
R1142 B.n330 B.n103 10.6151
R1143 B.n334 B.n103 10.6151
R1144 B.n335 B.n334 10.6151
R1145 B.n336 B.n335 10.6151
R1146 B.n336 B.n101 10.6151
R1147 B.n340 B.n101 10.6151
R1148 B.n341 B.n340 10.6151
R1149 B.n342 B.n341 10.6151
R1150 B.n342 B.n99 10.6151
R1151 B.n346 B.n99 10.6151
R1152 B.n347 B.n346 10.6151
R1153 B.n348 B.n347 10.6151
R1154 B.n348 B.n97 10.6151
R1155 B.n352 B.n97 10.6151
R1156 B.n353 B.n352 10.6151
R1157 B.n354 B.n353 10.6151
R1158 B.n354 B.n95 10.6151
R1159 B.n358 B.n95 10.6151
R1160 B.n359 B.n358 10.6151
R1161 B.n360 B.n359 10.6151
R1162 B.n360 B.n93 10.6151
R1163 B.n364 B.n93 10.6151
R1164 B.n365 B.n364 10.6151
R1165 B.n366 B.n365 10.6151
R1166 B.n366 B.n91 10.6151
R1167 B.n370 B.n91 10.6151
R1168 B.n371 B.n370 10.6151
R1169 B.n372 B.n371 10.6151
R1170 B.n372 B.n89 10.6151
R1171 B.n376 B.n89 10.6151
R1172 B.n377 B.n376 10.6151
R1173 B.n378 B.n377 10.6151
R1174 B.n378 B.n87 10.6151
R1175 B.n382 B.n87 10.6151
R1176 B.n383 B.n382 10.6151
R1177 B.n384 B.n383 10.6151
R1178 B.n384 B.n85 10.6151
R1179 B.n388 B.n85 10.6151
R1180 B.n389 B.n388 10.6151
R1181 B.n390 B.n389 10.6151
R1182 B.n390 B.n83 10.6151
R1183 B.n394 B.n83 10.6151
R1184 B.n395 B.n394 10.6151
R1185 B.n396 B.n395 10.6151
R1186 B.n396 B.n81 10.6151
R1187 B.n400 B.n81 10.6151
R1188 B.n401 B.n400 10.6151
R1189 B.n402 B.n401 10.6151
R1190 B.n402 B.n79 10.6151
R1191 B.n406 B.n79 10.6151
R1192 B.n407 B.n406 10.6151
R1193 B.n408 B.n407 10.6151
R1194 B.n408 B.n77 10.6151
R1195 B.n412 B.n77 10.6151
R1196 B.n413 B.n412 10.6151
R1197 B.n414 B.n413 10.6151
R1198 B.n414 B.n75 10.6151
R1199 B.n418 B.n75 10.6151
R1200 B.n419 B.n418 10.6151
R1201 B.n420 B.n419 10.6151
R1202 B.n420 B.n73 10.6151
R1203 B.n424 B.n73 10.6151
R1204 B.n425 B.n424 10.6151
R1205 B.n426 B.n425 10.6151
R1206 B.n426 B.n71 10.6151
R1207 B.n430 B.n71 10.6151
R1208 B.n431 B.n430 10.6151
R1209 B.n432 B.n431 10.6151
R1210 B.n432 B.n69 10.6151
R1211 B.n436 B.n69 10.6151
R1212 B.n437 B.n436 10.6151
R1213 B.n438 B.n437 10.6151
R1214 B.n438 B.n67 10.6151
R1215 B.n442 B.n67 10.6151
R1216 B.n443 B.n442 10.6151
R1217 B.n444 B.n443 10.6151
R1218 B.n444 B.n65 10.6151
R1219 B.n448 B.n65 10.6151
R1220 B.n449 B.n448 10.6151
R1221 B.n450 B.n449 10.6151
R1222 B.n450 B.n63 10.6151
R1223 B.n454 B.n63 10.6151
R1224 B.n455 B.n454 10.6151
R1225 B.n456 B.n455 10.6151
R1226 B.n456 B.n61 10.6151
R1227 B.n460 B.n61 10.6151
R1228 B.n461 B.n460 10.6151
R1229 B.n462 B.n461 10.6151
R1230 B.n462 B.n59 10.6151
R1231 B.n234 B.n139 10.6151
R1232 B.n238 B.n139 10.6151
R1233 B.n239 B.n238 10.6151
R1234 B.n240 B.n239 10.6151
R1235 B.n240 B.n137 10.6151
R1236 B.n244 B.n137 10.6151
R1237 B.n245 B.n244 10.6151
R1238 B.n246 B.n245 10.6151
R1239 B.n246 B.n135 10.6151
R1240 B.n250 B.n135 10.6151
R1241 B.n251 B.n250 10.6151
R1242 B.n252 B.n251 10.6151
R1243 B.n252 B.n133 10.6151
R1244 B.n256 B.n133 10.6151
R1245 B.n257 B.n256 10.6151
R1246 B.n258 B.n257 10.6151
R1247 B.n258 B.n131 10.6151
R1248 B.n262 B.n131 10.6151
R1249 B.n263 B.n262 10.6151
R1250 B.n264 B.n263 10.6151
R1251 B.n264 B.n129 10.6151
R1252 B.n268 B.n129 10.6151
R1253 B.n271 B.n270 10.6151
R1254 B.n271 B.n125 10.6151
R1255 B.n275 B.n125 10.6151
R1256 B.n276 B.n275 10.6151
R1257 B.n277 B.n276 10.6151
R1258 B.n277 B.n123 10.6151
R1259 B.n281 B.n123 10.6151
R1260 B.n282 B.n281 10.6151
R1261 B.n283 B.n282 10.6151
R1262 B.n287 B.n286 10.6151
R1263 B.n288 B.n287 10.6151
R1264 B.n288 B.n117 10.6151
R1265 B.n292 B.n117 10.6151
R1266 B.n293 B.n292 10.6151
R1267 B.n294 B.n293 10.6151
R1268 B.n294 B.n115 10.6151
R1269 B.n298 B.n115 10.6151
R1270 B.n299 B.n298 10.6151
R1271 B.n300 B.n299 10.6151
R1272 B.n300 B.n113 10.6151
R1273 B.n304 B.n113 10.6151
R1274 B.n305 B.n304 10.6151
R1275 B.n306 B.n305 10.6151
R1276 B.n306 B.n111 10.6151
R1277 B.n310 B.n111 10.6151
R1278 B.n311 B.n310 10.6151
R1279 B.n312 B.n311 10.6151
R1280 B.n312 B.n109 10.6151
R1281 B.n316 B.n109 10.6151
R1282 B.n317 B.n316 10.6151
R1283 B.n318 B.n317 10.6151
R1284 B.n233 B.n232 10.6151
R1285 B.n232 B.n141 10.6151
R1286 B.n228 B.n141 10.6151
R1287 B.n228 B.n227 10.6151
R1288 B.n227 B.n226 10.6151
R1289 B.n226 B.n143 10.6151
R1290 B.n222 B.n143 10.6151
R1291 B.n222 B.n221 10.6151
R1292 B.n221 B.n220 10.6151
R1293 B.n220 B.n145 10.6151
R1294 B.n216 B.n145 10.6151
R1295 B.n216 B.n215 10.6151
R1296 B.n215 B.n214 10.6151
R1297 B.n214 B.n147 10.6151
R1298 B.n210 B.n147 10.6151
R1299 B.n210 B.n209 10.6151
R1300 B.n209 B.n208 10.6151
R1301 B.n208 B.n149 10.6151
R1302 B.n204 B.n149 10.6151
R1303 B.n204 B.n203 10.6151
R1304 B.n203 B.n202 10.6151
R1305 B.n202 B.n151 10.6151
R1306 B.n198 B.n151 10.6151
R1307 B.n198 B.n197 10.6151
R1308 B.n197 B.n196 10.6151
R1309 B.n196 B.n153 10.6151
R1310 B.n192 B.n153 10.6151
R1311 B.n192 B.n191 10.6151
R1312 B.n191 B.n190 10.6151
R1313 B.n190 B.n155 10.6151
R1314 B.n186 B.n155 10.6151
R1315 B.n186 B.n185 10.6151
R1316 B.n185 B.n184 10.6151
R1317 B.n184 B.n157 10.6151
R1318 B.n180 B.n157 10.6151
R1319 B.n180 B.n179 10.6151
R1320 B.n179 B.n178 10.6151
R1321 B.n178 B.n159 10.6151
R1322 B.n174 B.n159 10.6151
R1323 B.n174 B.n173 10.6151
R1324 B.n173 B.n172 10.6151
R1325 B.n172 B.n161 10.6151
R1326 B.n168 B.n161 10.6151
R1327 B.n168 B.n167 10.6151
R1328 B.n167 B.n166 10.6151
R1329 B.n166 B.n163 10.6151
R1330 B.n163 B.n0 10.6151
R1331 B.n619 B.n1 10.6151
R1332 B.n619 B.n618 10.6151
R1333 B.n618 B.n617 10.6151
R1334 B.n617 B.n4 10.6151
R1335 B.n613 B.n4 10.6151
R1336 B.n613 B.n612 10.6151
R1337 B.n612 B.n611 10.6151
R1338 B.n611 B.n6 10.6151
R1339 B.n607 B.n6 10.6151
R1340 B.n607 B.n606 10.6151
R1341 B.n606 B.n605 10.6151
R1342 B.n605 B.n8 10.6151
R1343 B.n601 B.n8 10.6151
R1344 B.n601 B.n600 10.6151
R1345 B.n600 B.n599 10.6151
R1346 B.n599 B.n10 10.6151
R1347 B.n595 B.n10 10.6151
R1348 B.n595 B.n594 10.6151
R1349 B.n594 B.n593 10.6151
R1350 B.n593 B.n12 10.6151
R1351 B.n589 B.n12 10.6151
R1352 B.n589 B.n588 10.6151
R1353 B.n588 B.n587 10.6151
R1354 B.n587 B.n14 10.6151
R1355 B.n583 B.n14 10.6151
R1356 B.n583 B.n582 10.6151
R1357 B.n582 B.n581 10.6151
R1358 B.n581 B.n16 10.6151
R1359 B.n577 B.n16 10.6151
R1360 B.n577 B.n576 10.6151
R1361 B.n576 B.n575 10.6151
R1362 B.n575 B.n18 10.6151
R1363 B.n571 B.n18 10.6151
R1364 B.n571 B.n570 10.6151
R1365 B.n570 B.n569 10.6151
R1366 B.n569 B.n20 10.6151
R1367 B.n565 B.n20 10.6151
R1368 B.n565 B.n564 10.6151
R1369 B.n564 B.n563 10.6151
R1370 B.n563 B.n22 10.6151
R1371 B.n559 B.n22 10.6151
R1372 B.n559 B.n558 10.6151
R1373 B.n558 B.n557 10.6151
R1374 B.n557 B.n24 10.6151
R1375 B.n553 B.n24 10.6151
R1376 B.n553 B.n552 10.6151
R1377 B.n552 B.n551 10.6151
R1378 B.n516 B.n515 9.36635
R1379 B.n498 B.n48 9.36635
R1380 B.n269 B.n268 9.36635
R1381 B.n286 B.n121 9.36635
R1382 B.n623 B.n0 2.81026
R1383 B.n623 B.n1 2.81026
R1384 B.n515 B.n514 1.24928
R1385 B.n48 B.n44 1.24928
R1386 B.n270 B.n269 1.24928
R1387 B.n283 B.n121 1.24928
R1388 VN.n32 VN.n31 183.81
R1389 VN.n65 VN.n64 183.81
R1390 VN.n63 VN.n33 161.3
R1391 VN.n62 VN.n61 161.3
R1392 VN.n60 VN.n34 161.3
R1393 VN.n59 VN.n58 161.3
R1394 VN.n57 VN.n35 161.3
R1395 VN.n55 VN.n54 161.3
R1396 VN.n53 VN.n36 161.3
R1397 VN.n52 VN.n51 161.3
R1398 VN.n50 VN.n37 161.3
R1399 VN.n49 VN.n48 161.3
R1400 VN.n47 VN.n38 161.3
R1401 VN.n46 VN.n45 161.3
R1402 VN.n44 VN.n39 161.3
R1403 VN.n43 VN.n42 161.3
R1404 VN.n30 VN.n0 161.3
R1405 VN.n29 VN.n28 161.3
R1406 VN.n27 VN.n1 161.3
R1407 VN.n26 VN.n25 161.3
R1408 VN.n24 VN.n2 161.3
R1409 VN.n22 VN.n21 161.3
R1410 VN.n20 VN.n3 161.3
R1411 VN.n19 VN.n18 161.3
R1412 VN.n17 VN.n4 161.3
R1413 VN.n16 VN.n15 161.3
R1414 VN.n14 VN.n5 161.3
R1415 VN.n13 VN.n12 161.3
R1416 VN.n11 VN.n6 161.3
R1417 VN.n10 VN.n9 161.3
R1418 VN.n8 VN.t8 105.222
R1419 VN.n41 VN.t2 105.222
R1420 VN.n16 VN.t3 72.4247
R1421 VN.n7 VN.t7 72.4247
R1422 VN.n23 VN.t1 72.4247
R1423 VN.n31 VN.t6 72.4247
R1424 VN.n49 VN.t0 72.4247
R1425 VN.n40 VN.t4 72.4247
R1426 VN.n56 VN.t5 72.4247
R1427 VN.n64 VN.t9 72.4247
R1428 VN.n8 VN.n7 56.8484
R1429 VN.n41 VN.n40 56.8484
R1430 VN.n12 VN.n11 53.6055
R1431 VN.n18 VN.n3 53.6055
R1432 VN.n45 VN.n44 53.6055
R1433 VN.n51 VN.n36 53.6055
R1434 VN.n25 VN.n1 49.7204
R1435 VN.n58 VN.n34 49.7204
R1436 VN VN.n65 45.1425
R1437 VN.n29 VN.n1 31.2664
R1438 VN.n62 VN.n34 31.2664
R1439 VN.n12 VN.n5 27.3813
R1440 VN.n18 VN.n17 27.3813
R1441 VN.n45 VN.n38 27.3813
R1442 VN.n51 VN.n50 27.3813
R1443 VN.n11 VN.n10 24.4675
R1444 VN.n16 VN.n5 24.4675
R1445 VN.n17 VN.n16 24.4675
R1446 VN.n22 VN.n3 24.4675
R1447 VN.n25 VN.n24 24.4675
R1448 VN.n30 VN.n29 24.4675
R1449 VN.n44 VN.n43 24.4675
R1450 VN.n50 VN.n49 24.4675
R1451 VN.n49 VN.n38 24.4675
R1452 VN.n58 VN.n57 24.4675
R1453 VN.n55 VN.n36 24.4675
R1454 VN.n63 VN.n62 24.4675
R1455 VN.n10 VN.n7 13.2127
R1456 VN.n23 VN.n22 13.2127
R1457 VN.n43 VN.n40 13.2127
R1458 VN.n56 VN.n55 13.2127
R1459 VN.n42 VN.n41 12.4717
R1460 VN.n9 VN.n8 12.4717
R1461 VN.n24 VN.n23 11.2553
R1462 VN.n57 VN.n56 11.2553
R1463 VN.n31 VN.n30 1.95786
R1464 VN.n64 VN.n63 1.95786
R1465 VN.n65 VN.n33 0.189894
R1466 VN.n61 VN.n33 0.189894
R1467 VN.n61 VN.n60 0.189894
R1468 VN.n60 VN.n59 0.189894
R1469 VN.n59 VN.n35 0.189894
R1470 VN.n54 VN.n35 0.189894
R1471 VN.n54 VN.n53 0.189894
R1472 VN.n53 VN.n52 0.189894
R1473 VN.n52 VN.n37 0.189894
R1474 VN.n48 VN.n37 0.189894
R1475 VN.n48 VN.n47 0.189894
R1476 VN.n47 VN.n46 0.189894
R1477 VN.n46 VN.n39 0.189894
R1478 VN.n42 VN.n39 0.189894
R1479 VN.n9 VN.n6 0.189894
R1480 VN.n13 VN.n6 0.189894
R1481 VN.n14 VN.n13 0.189894
R1482 VN.n15 VN.n14 0.189894
R1483 VN.n15 VN.n4 0.189894
R1484 VN.n19 VN.n4 0.189894
R1485 VN.n20 VN.n19 0.189894
R1486 VN.n21 VN.n20 0.189894
R1487 VN.n21 VN.n2 0.189894
R1488 VN.n26 VN.n2 0.189894
R1489 VN.n27 VN.n26 0.189894
R1490 VN.n28 VN.n27 0.189894
R1491 VN.n28 VN.n0 0.189894
R1492 VN.n32 VN.n0 0.189894
R1493 VN VN.n32 0.0516364
R1494 VDD2.n61 VDD2.n60 756.745
R1495 VDD2.n28 VDD2.n27 756.745
R1496 VDD2.n60 VDD2.n59 585
R1497 VDD2.n35 VDD2.n34 585
R1498 VDD2.n54 VDD2.n53 585
R1499 VDD2.n52 VDD2.n51 585
R1500 VDD2.n39 VDD2.n38 585
R1501 VDD2.n46 VDD2.n45 585
R1502 VDD2.n44 VDD2.n43 585
R1503 VDD2.n11 VDD2.n10 585
R1504 VDD2.n13 VDD2.n12 585
R1505 VDD2.n6 VDD2.n5 585
R1506 VDD2.n19 VDD2.n18 585
R1507 VDD2.n21 VDD2.n20 585
R1508 VDD2.n2 VDD2.n1 585
R1509 VDD2.n27 VDD2.n26 585
R1510 VDD2.n9 VDD2.t1 329.175
R1511 VDD2.n42 VDD2.t0 329.175
R1512 VDD2.n60 VDD2.n34 171.744
R1513 VDD2.n53 VDD2.n34 171.744
R1514 VDD2.n53 VDD2.n52 171.744
R1515 VDD2.n52 VDD2.n38 171.744
R1516 VDD2.n45 VDD2.n38 171.744
R1517 VDD2.n45 VDD2.n44 171.744
R1518 VDD2.n12 VDD2.n11 171.744
R1519 VDD2.n12 VDD2.n5 171.744
R1520 VDD2.n19 VDD2.n5 171.744
R1521 VDD2.n20 VDD2.n19 171.744
R1522 VDD2.n20 VDD2.n1 171.744
R1523 VDD2.n27 VDD2.n1 171.744
R1524 VDD2.n32 VDD2.n31 96.7182
R1525 VDD2 VDD2.n65 96.7152
R1526 VDD2.n64 VDD2.n63 95.3069
R1527 VDD2.n30 VDD2.n29 95.3059
R1528 VDD2.n44 VDD2.t0 85.8723
R1529 VDD2.n11 VDD2.t1 85.8723
R1530 VDD2.n30 VDD2.n28 53.3422
R1531 VDD2.n62 VDD2.n61 51.3853
R1532 VDD2.n62 VDD2.n32 38.0364
R1533 VDD2.n59 VDD2.n33 12.0247
R1534 VDD2.n26 VDD2.n0 12.0247
R1535 VDD2.n58 VDD2.n35 11.249
R1536 VDD2.n25 VDD2.n2 11.249
R1537 VDD2.n10 VDD2.n9 10.722
R1538 VDD2.n43 VDD2.n42 10.722
R1539 VDD2.n55 VDD2.n54 10.4732
R1540 VDD2.n22 VDD2.n21 10.4732
R1541 VDD2.n51 VDD2.n37 9.69747
R1542 VDD2.n18 VDD2.n4 9.69747
R1543 VDD2.n57 VDD2.n33 9.45567
R1544 VDD2.n24 VDD2.n0 9.45567
R1545 VDD2.n48 VDD2.n47 9.3005
R1546 VDD2.n50 VDD2.n49 9.3005
R1547 VDD2.n37 VDD2.n36 9.3005
R1548 VDD2.n56 VDD2.n55 9.3005
R1549 VDD2.n58 VDD2.n57 9.3005
R1550 VDD2.n41 VDD2.n40 9.3005
R1551 VDD2.n8 VDD2.n7 9.3005
R1552 VDD2.n15 VDD2.n14 9.3005
R1553 VDD2.n17 VDD2.n16 9.3005
R1554 VDD2.n4 VDD2.n3 9.3005
R1555 VDD2.n23 VDD2.n22 9.3005
R1556 VDD2.n25 VDD2.n24 9.3005
R1557 VDD2.n50 VDD2.n39 8.92171
R1558 VDD2.n17 VDD2.n6 8.92171
R1559 VDD2.n47 VDD2.n46 8.14595
R1560 VDD2.n14 VDD2.n13 8.14595
R1561 VDD2.n43 VDD2.n41 7.3702
R1562 VDD2.n10 VDD2.n8 7.3702
R1563 VDD2.n46 VDD2.n41 5.81868
R1564 VDD2.n13 VDD2.n8 5.81868
R1565 VDD2.n65 VDD2.t5 5.57597
R1566 VDD2.n65 VDD2.t7 5.57597
R1567 VDD2.n63 VDD2.t4 5.57597
R1568 VDD2.n63 VDD2.t9 5.57597
R1569 VDD2.n31 VDD2.t8 5.57597
R1570 VDD2.n31 VDD2.t3 5.57597
R1571 VDD2.n29 VDD2.t2 5.57597
R1572 VDD2.n29 VDD2.t6 5.57597
R1573 VDD2.n47 VDD2.n39 5.04292
R1574 VDD2.n14 VDD2.n6 5.04292
R1575 VDD2.n51 VDD2.n50 4.26717
R1576 VDD2.n18 VDD2.n17 4.26717
R1577 VDD2.n54 VDD2.n37 3.49141
R1578 VDD2.n21 VDD2.n4 3.49141
R1579 VDD2.n55 VDD2.n35 2.71565
R1580 VDD2.n22 VDD2.n2 2.71565
R1581 VDD2.n9 VDD2.n7 2.4147
R1582 VDD2.n42 VDD2.n40 2.4147
R1583 VDD2.n64 VDD2.n62 1.9574
R1584 VDD2.n59 VDD2.n58 1.93989
R1585 VDD2.n26 VDD2.n25 1.93989
R1586 VDD2.n61 VDD2.n33 1.16414
R1587 VDD2.n28 VDD2.n0 1.16414
R1588 VDD2 VDD2.n64 0.547914
R1589 VDD2.n32 VDD2.n30 0.434378
R1590 VDD2.n57 VDD2.n56 0.155672
R1591 VDD2.n56 VDD2.n36 0.155672
R1592 VDD2.n49 VDD2.n36 0.155672
R1593 VDD2.n49 VDD2.n48 0.155672
R1594 VDD2.n48 VDD2.n40 0.155672
R1595 VDD2.n15 VDD2.n7 0.155672
R1596 VDD2.n16 VDD2.n15 0.155672
R1597 VDD2.n16 VDD2.n3 0.155672
R1598 VDD2.n23 VDD2.n3 0.155672
R1599 VDD2.n24 VDD2.n23 0.155672
C0 w_n3694_n2134# B 7.71628f
C1 VTAIL B 2.11832f
C2 B VP 1.84041f
C3 VTAIL w_n3694_n2134# 2.23604f
C4 VDD1 VN 0.151805f
C5 w_n3694_n2134# VP 8.064981f
C6 VTAIL VP 5.90416f
C7 VDD1 VDD2 1.7438f
C8 B VN 1.03875f
C9 w_n3694_n2134# VN 7.58607f
C10 B VDD2 1.83359f
C11 VTAIL VN 5.88993f
C12 w_n3694_n2134# VDD2 2.21082f
C13 VN VP 6.28105f
C14 VTAIL VDD2 7.21163f
C15 VP VDD2 0.498779f
C16 VDD1 B 1.74134f
C17 w_n3694_n2134# VDD1 2.10151f
C18 VTAIL VDD1 7.16411f
C19 VN VDD2 5.10348f
C20 VDD1 VP 5.44787f
C21 VDD2 VSUBS 1.573035f
C22 VDD1 VSUBS 1.485596f
C23 VTAIL VSUBS 0.601297f
C24 VN VSUBS 6.2932f
C25 VP VSUBS 2.977799f
C26 B VSUBS 4.023697f
C27 w_n3694_n2134# VSUBS 98.4525f
C28 VDD2.n0 VSUBS 0.015008f
C29 VDD2.n1 VSUBS 0.033823f
C30 VDD2.n2 VSUBS 0.015152f
C31 VDD2.n3 VSUBS 0.02663f
C32 VDD2.n4 VSUBS 0.01431f
C33 VDD2.n5 VSUBS 0.033823f
C34 VDD2.n6 VSUBS 0.015152f
C35 VDD2.n7 VSUBS 0.587536f
C36 VDD2.n8 VSUBS 0.01431f
C37 VDD2.t1 VSUBS 0.072863f
C38 VDD2.n9 VSUBS 0.135858f
C39 VDD2.n10 VSUBS 0.025433f
C40 VDD2.n11 VSUBS 0.025367f
C41 VDD2.n12 VSUBS 0.033823f
C42 VDD2.n13 VSUBS 0.015152f
C43 VDD2.n14 VSUBS 0.01431f
C44 VDD2.n15 VSUBS 0.02663f
C45 VDD2.n16 VSUBS 0.02663f
C46 VDD2.n17 VSUBS 0.01431f
C47 VDD2.n18 VSUBS 0.015152f
C48 VDD2.n19 VSUBS 0.033823f
C49 VDD2.n20 VSUBS 0.033823f
C50 VDD2.n21 VSUBS 0.015152f
C51 VDD2.n22 VSUBS 0.01431f
C52 VDD2.n23 VSUBS 0.02663f
C53 VDD2.n24 VSUBS 0.068466f
C54 VDD2.n25 VSUBS 0.01431f
C55 VDD2.n26 VSUBS 0.015152f
C56 VDD2.n27 VSUBS 0.074966f
C57 VDD2.n28 VSUBS 0.076707f
C58 VDD2.t2 VSUBS 0.122685f
C59 VDD2.t6 VSUBS 0.122685f
C60 VDD2.n29 VSUBS 0.825225f
C61 VDD2.n30 VSUBS 0.830237f
C62 VDD2.t8 VSUBS 0.122685f
C63 VDD2.t3 VSUBS 0.122685f
C64 VDD2.n31 VSUBS 0.835596f
C65 VDD2.n32 VSUBS 2.52122f
C66 VDD2.n33 VSUBS 0.015008f
C67 VDD2.n34 VSUBS 0.033823f
C68 VDD2.n35 VSUBS 0.015152f
C69 VDD2.n36 VSUBS 0.02663f
C70 VDD2.n37 VSUBS 0.01431f
C71 VDD2.n38 VSUBS 0.033823f
C72 VDD2.n39 VSUBS 0.015152f
C73 VDD2.n40 VSUBS 0.587536f
C74 VDD2.n41 VSUBS 0.01431f
C75 VDD2.t0 VSUBS 0.072863f
C76 VDD2.n42 VSUBS 0.135858f
C77 VDD2.n43 VSUBS 0.025433f
C78 VDD2.n44 VSUBS 0.025367f
C79 VDD2.n45 VSUBS 0.033823f
C80 VDD2.n46 VSUBS 0.015152f
C81 VDD2.n47 VSUBS 0.01431f
C82 VDD2.n48 VSUBS 0.02663f
C83 VDD2.n49 VSUBS 0.02663f
C84 VDD2.n50 VSUBS 0.01431f
C85 VDD2.n51 VSUBS 0.015152f
C86 VDD2.n52 VSUBS 0.033823f
C87 VDD2.n53 VSUBS 0.033823f
C88 VDD2.n54 VSUBS 0.015152f
C89 VDD2.n55 VSUBS 0.01431f
C90 VDD2.n56 VSUBS 0.02663f
C91 VDD2.n57 VSUBS 0.068466f
C92 VDD2.n58 VSUBS 0.01431f
C93 VDD2.n59 VSUBS 0.015152f
C94 VDD2.n60 VSUBS 0.074966f
C95 VDD2.n61 VSUBS 0.068566f
C96 VDD2.n62 VSUBS 2.29251f
C97 VDD2.t4 VSUBS 0.122685f
C98 VDD2.t9 VSUBS 0.122685f
C99 VDD2.n63 VSUBS 0.825227f
C100 VDD2.n64 VSUBS 0.624792f
C101 VDD2.t5 VSUBS 0.122685f
C102 VDD2.t7 VSUBS 0.122685f
C103 VDD2.n65 VSUBS 0.835563f
C104 VN.n0 VSUBS 0.040515f
C105 VN.t6 VSUBS 1.21076f
C106 VN.n1 VSUBS 0.037708f
C107 VN.n2 VSUBS 0.040515f
C108 VN.t1 VSUBS 1.21076f
C109 VN.n3 VSUBS 0.071457f
C110 VN.n4 VSUBS 0.040515f
C111 VN.t3 VSUBS 1.21076f
C112 VN.n5 VSUBS 0.079001f
C113 VN.n6 VSUBS 0.040515f
C114 VN.t7 VSUBS 1.21076f
C115 VN.n7 VSUBS 0.561565f
C116 VN.t8 VSUBS 1.4188f
C117 VN.n8 VSUBS 0.557388f
C118 VN.n9 VSUBS 0.301975f
C119 VN.n10 VSUBS 0.058361f
C120 VN.n11 VSUBS 0.071457f
C121 VN.n12 VSUBS 0.043349f
C122 VN.n13 VSUBS 0.040515f
C123 VN.n14 VSUBS 0.040515f
C124 VN.n15 VSUBS 0.040515f
C125 VN.n16 VSUBS 0.50357f
C126 VN.n17 VSUBS 0.079001f
C127 VN.n18 VSUBS 0.043349f
C128 VN.n19 VSUBS 0.040515f
C129 VN.n20 VSUBS 0.040515f
C130 VN.n21 VSUBS 0.040515f
C131 VN.n22 VSUBS 0.058361f
C132 VN.n23 VSUBS 0.46534f
C133 VN.n24 VSUBS 0.055379f
C134 VN.n25 VSUBS 0.074752f
C135 VN.n26 VSUBS 0.040515f
C136 VN.n27 VSUBS 0.040515f
C137 VN.n28 VSUBS 0.040515f
C138 VN.n29 VSUBS 0.081346f
C139 VN.n30 VSUBS 0.041212f
C140 VN.n31 VSUBS 0.563008f
C141 VN.n32 VSUBS 0.045027f
C142 VN.n33 VSUBS 0.040515f
C143 VN.t9 VSUBS 1.21076f
C144 VN.n34 VSUBS 0.037708f
C145 VN.n35 VSUBS 0.040515f
C146 VN.t5 VSUBS 1.21076f
C147 VN.n36 VSUBS 0.071457f
C148 VN.n37 VSUBS 0.040515f
C149 VN.t0 VSUBS 1.21076f
C150 VN.n38 VSUBS 0.079001f
C151 VN.n39 VSUBS 0.040515f
C152 VN.t4 VSUBS 1.21076f
C153 VN.n40 VSUBS 0.561565f
C154 VN.t2 VSUBS 1.4188f
C155 VN.n41 VSUBS 0.557388f
C156 VN.n42 VSUBS 0.301975f
C157 VN.n43 VSUBS 0.058361f
C158 VN.n44 VSUBS 0.071457f
C159 VN.n45 VSUBS 0.043349f
C160 VN.n46 VSUBS 0.040515f
C161 VN.n47 VSUBS 0.040515f
C162 VN.n48 VSUBS 0.040515f
C163 VN.n49 VSUBS 0.50357f
C164 VN.n50 VSUBS 0.079001f
C165 VN.n51 VSUBS 0.043349f
C166 VN.n52 VSUBS 0.040515f
C167 VN.n53 VSUBS 0.040515f
C168 VN.n54 VSUBS 0.040515f
C169 VN.n55 VSUBS 0.058361f
C170 VN.n56 VSUBS 0.46534f
C171 VN.n57 VSUBS 0.055379f
C172 VN.n58 VSUBS 0.074752f
C173 VN.n59 VSUBS 0.040515f
C174 VN.n60 VSUBS 0.040515f
C175 VN.n61 VSUBS 0.040515f
C176 VN.n62 VSUBS 0.081346f
C177 VN.n63 VSUBS 0.041212f
C178 VN.n64 VSUBS 0.563008f
C179 VN.n65 VSUBS 1.89566f
C180 B.n0 VSUBS 0.00496f
C181 B.n1 VSUBS 0.00496f
C182 B.n2 VSUBS 0.007844f
C183 B.n3 VSUBS 0.007844f
C184 B.n4 VSUBS 0.007844f
C185 B.n5 VSUBS 0.007844f
C186 B.n6 VSUBS 0.007844f
C187 B.n7 VSUBS 0.007844f
C188 B.n8 VSUBS 0.007844f
C189 B.n9 VSUBS 0.007844f
C190 B.n10 VSUBS 0.007844f
C191 B.n11 VSUBS 0.007844f
C192 B.n12 VSUBS 0.007844f
C193 B.n13 VSUBS 0.007844f
C194 B.n14 VSUBS 0.007844f
C195 B.n15 VSUBS 0.007844f
C196 B.n16 VSUBS 0.007844f
C197 B.n17 VSUBS 0.007844f
C198 B.n18 VSUBS 0.007844f
C199 B.n19 VSUBS 0.007844f
C200 B.n20 VSUBS 0.007844f
C201 B.n21 VSUBS 0.007844f
C202 B.n22 VSUBS 0.007844f
C203 B.n23 VSUBS 0.007844f
C204 B.n24 VSUBS 0.007844f
C205 B.n25 VSUBS 0.007844f
C206 B.n26 VSUBS 0.020285f
C207 B.n27 VSUBS 0.007844f
C208 B.n28 VSUBS 0.007844f
C209 B.n29 VSUBS 0.007844f
C210 B.n30 VSUBS 0.007844f
C211 B.n31 VSUBS 0.007844f
C212 B.n32 VSUBS 0.007844f
C213 B.n33 VSUBS 0.007844f
C214 B.n34 VSUBS 0.007844f
C215 B.n35 VSUBS 0.007844f
C216 B.n36 VSUBS 0.007844f
C217 B.n37 VSUBS 0.007844f
C218 B.t2 VSUBS 0.096595f
C219 B.t1 VSUBS 0.119089f
C220 B.t0 VSUBS 0.591045f
C221 B.n38 VSUBS 0.207916f
C222 B.n39 VSUBS 0.16903f
C223 B.n40 VSUBS 0.007844f
C224 B.n41 VSUBS 0.007844f
C225 B.n42 VSUBS 0.007844f
C226 B.n43 VSUBS 0.007844f
C227 B.n44 VSUBS 0.004383f
C228 B.n45 VSUBS 0.007844f
C229 B.t8 VSUBS 0.096597f
C230 B.t7 VSUBS 0.119091f
C231 B.t6 VSUBS 0.591045f
C232 B.n46 VSUBS 0.207914f
C233 B.n47 VSUBS 0.169028f
C234 B.n48 VSUBS 0.018173f
C235 B.n49 VSUBS 0.007844f
C236 B.n50 VSUBS 0.007844f
C237 B.n51 VSUBS 0.007844f
C238 B.n52 VSUBS 0.007844f
C239 B.n53 VSUBS 0.007844f
C240 B.n54 VSUBS 0.007844f
C241 B.n55 VSUBS 0.007844f
C242 B.n56 VSUBS 0.007844f
C243 B.n57 VSUBS 0.007844f
C244 B.n58 VSUBS 0.007844f
C245 B.n59 VSUBS 0.020445f
C246 B.n60 VSUBS 0.007844f
C247 B.n61 VSUBS 0.007844f
C248 B.n62 VSUBS 0.007844f
C249 B.n63 VSUBS 0.007844f
C250 B.n64 VSUBS 0.007844f
C251 B.n65 VSUBS 0.007844f
C252 B.n66 VSUBS 0.007844f
C253 B.n67 VSUBS 0.007844f
C254 B.n68 VSUBS 0.007844f
C255 B.n69 VSUBS 0.007844f
C256 B.n70 VSUBS 0.007844f
C257 B.n71 VSUBS 0.007844f
C258 B.n72 VSUBS 0.007844f
C259 B.n73 VSUBS 0.007844f
C260 B.n74 VSUBS 0.007844f
C261 B.n75 VSUBS 0.007844f
C262 B.n76 VSUBS 0.007844f
C263 B.n77 VSUBS 0.007844f
C264 B.n78 VSUBS 0.007844f
C265 B.n79 VSUBS 0.007844f
C266 B.n80 VSUBS 0.007844f
C267 B.n81 VSUBS 0.007844f
C268 B.n82 VSUBS 0.007844f
C269 B.n83 VSUBS 0.007844f
C270 B.n84 VSUBS 0.007844f
C271 B.n85 VSUBS 0.007844f
C272 B.n86 VSUBS 0.007844f
C273 B.n87 VSUBS 0.007844f
C274 B.n88 VSUBS 0.007844f
C275 B.n89 VSUBS 0.007844f
C276 B.n90 VSUBS 0.007844f
C277 B.n91 VSUBS 0.007844f
C278 B.n92 VSUBS 0.007844f
C279 B.n93 VSUBS 0.007844f
C280 B.n94 VSUBS 0.007844f
C281 B.n95 VSUBS 0.007844f
C282 B.n96 VSUBS 0.007844f
C283 B.n97 VSUBS 0.007844f
C284 B.n98 VSUBS 0.007844f
C285 B.n99 VSUBS 0.007844f
C286 B.n100 VSUBS 0.007844f
C287 B.n101 VSUBS 0.007844f
C288 B.n102 VSUBS 0.007844f
C289 B.n103 VSUBS 0.007844f
C290 B.n104 VSUBS 0.007844f
C291 B.n105 VSUBS 0.007844f
C292 B.n106 VSUBS 0.007844f
C293 B.n107 VSUBS 0.019626f
C294 B.n108 VSUBS 0.007844f
C295 B.n109 VSUBS 0.007844f
C296 B.n110 VSUBS 0.007844f
C297 B.n111 VSUBS 0.007844f
C298 B.n112 VSUBS 0.007844f
C299 B.n113 VSUBS 0.007844f
C300 B.n114 VSUBS 0.007844f
C301 B.n115 VSUBS 0.007844f
C302 B.n116 VSUBS 0.007844f
C303 B.n117 VSUBS 0.007844f
C304 B.n118 VSUBS 0.007844f
C305 B.t10 VSUBS 0.096597f
C306 B.t11 VSUBS 0.119091f
C307 B.t9 VSUBS 0.591045f
C308 B.n119 VSUBS 0.207914f
C309 B.n120 VSUBS 0.169028f
C310 B.n121 VSUBS 0.018173f
C311 B.n122 VSUBS 0.007844f
C312 B.n123 VSUBS 0.007844f
C313 B.n124 VSUBS 0.007844f
C314 B.n125 VSUBS 0.007844f
C315 B.n126 VSUBS 0.007844f
C316 B.t4 VSUBS 0.096595f
C317 B.t5 VSUBS 0.119089f
C318 B.t3 VSUBS 0.591045f
C319 B.n127 VSUBS 0.207916f
C320 B.n128 VSUBS 0.16903f
C321 B.n129 VSUBS 0.007844f
C322 B.n130 VSUBS 0.007844f
C323 B.n131 VSUBS 0.007844f
C324 B.n132 VSUBS 0.007844f
C325 B.n133 VSUBS 0.007844f
C326 B.n134 VSUBS 0.007844f
C327 B.n135 VSUBS 0.007844f
C328 B.n136 VSUBS 0.007844f
C329 B.n137 VSUBS 0.007844f
C330 B.n138 VSUBS 0.007844f
C331 B.n139 VSUBS 0.007844f
C332 B.n140 VSUBS 0.019626f
C333 B.n141 VSUBS 0.007844f
C334 B.n142 VSUBS 0.007844f
C335 B.n143 VSUBS 0.007844f
C336 B.n144 VSUBS 0.007844f
C337 B.n145 VSUBS 0.007844f
C338 B.n146 VSUBS 0.007844f
C339 B.n147 VSUBS 0.007844f
C340 B.n148 VSUBS 0.007844f
C341 B.n149 VSUBS 0.007844f
C342 B.n150 VSUBS 0.007844f
C343 B.n151 VSUBS 0.007844f
C344 B.n152 VSUBS 0.007844f
C345 B.n153 VSUBS 0.007844f
C346 B.n154 VSUBS 0.007844f
C347 B.n155 VSUBS 0.007844f
C348 B.n156 VSUBS 0.007844f
C349 B.n157 VSUBS 0.007844f
C350 B.n158 VSUBS 0.007844f
C351 B.n159 VSUBS 0.007844f
C352 B.n160 VSUBS 0.007844f
C353 B.n161 VSUBS 0.007844f
C354 B.n162 VSUBS 0.007844f
C355 B.n163 VSUBS 0.007844f
C356 B.n164 VSUBS 0.007844f
C357 B.n165 VSUBS 0.007844f
C358 B.n166 VSUBS 0.007844f
C359 B.n167 VSUBS 0.007844f
C360 B.n168 VSUBS 0.007844f
C361 B.n169 VSUBS 0.007844f
C362 B.n170 VSUBS 0.007844f
C363 B.n171 VSUBS 0.007844f
C364 B.n172 VSUBS 0.007844f
C365 B.n173 VSUBS 0.007844f
C366 B.n174 VSUBS 0.007844f
C367 B.n175 VSUBS 0.007844f
C368 B.n176 VSUBS 0.007844f
C369 B.n177 VSUBS 0.007844f
C370 B.n178 VSUBS 0.007844f
C371 B.n179 VSUBS 0.007844f
C372 B.n180 VSUBS 0.007844f
C373 B.n181 VSUBS 0.007844f
C374 B.n182 VSUBS 0.007844f
C375 B.n183 VSUBS 0.007844f
C376 B.n184 VSUBS 0.007844f
C377 B.n185 VSUBS 0.007844f
C378 B.n186 VSUBS 0.007844f
C379 B.n187 VSUBS 0.007844f
C380 B.n188 VSUBS 0.007844f
C381 B.n189 VSUBS 0.007844f
C382 B.n190 VSUBS 0.007844f
C383 B.n191 VSUBS 0.007844f
C384 B.n192 VSUBS 0.007844f
C385 B.n193 VSUBS 0.007844f
C386 B.n194 VSUBS 0.007844f
C387 B.n195 VSUBS 0.007844f
C388 B.n196 VSUBS 0.007844f
C389 B.n197 VSUBS 0.007844f
C390 B.n198 VSUBS 0.007844f
C391 B.n199 VSUBS 0.007844f
C392 B.n200 VSUBS 0.007844f
C393 B.n201 VSUBS 0.007844f
C394 B.n202 VSUBS 0.007844f
C395 B.n203 VSUBS 0.007844f
C396 B.n204 VSUBS 0.007844f
C397 B.n205 VSUBS 0.007844f
C398 B.n206 VSUBS 0.007844f
C399 B.n207 VSUBS 0.007844f
C400 B.n208 VSUBS 0.007844f
C401 B.n209 VSUBS 0.007844f
C402 B.n210 VSUBS 0.007844f
C403 B.n211 VSUBS 0.007844f
C404 B.n212 VSUBS 0.007844f
C405 B.n213 VSUBS 0.007844f
C406 B.n214 VSUBS 0.007844f
C407 B.n215 VSUBS 0.007844f
C408 B.n216 VSUBS 0.007844f
C409 B.n217 VSUBS 0.007844f
C410 B.n218 VSUBS 0.007844f
C411 B.n219 VSUBS 0.007844f
C412 B.n220 VSUBS 0.007844f
C413 B.n221 VSUBS 0.007844f
C414 B.n222 VSUBS 0.007844f
C415 B.n223 VSUBS 0.007844f
C416 B.n224 VSUBS 0.007844f
C417 B.n225 VSUBS 0.007844f
C418 B.n226 VSUBS 0.007844f
C419 B.n227 VSUBS 0.007844f
C420 B.n228 VSUBS 0.007844f
C421 B.n229 VSUBS 0.007844f
C422 B.n230 VSUBS 0.007844f
C423 B.n231 VSUBS 0.007844f
C424 B.n232 VSUBS 0.007844f
C425 B.n233 VSUBS 0.019626f
C426 B.n234 VSUBS 0.020285f
C427 B.n235 VSUBS 0.020285f
C428 B.n236 VSUBS 0.007844f
C429 B.n237 VSUBS 0.007844f
C430 B.n238 VSUBS 0.007844f
C431 B.n239 VSUBS 0.007844f
C432 B.n240 VSUBS 0.007844f
C433 B.n241 VSUBS 0.007844f
C434 B.n242 VSUBS 0.007844f
C435 B.n243 VSUBS 0.007844f
C436 B.n244 VSUBS 0.007844f
C437 B.n245 VSUBS 0.007844f
C438 B.n246 VSUBS 0.007844f
C439 B.n247 VSUBS 0.007844f
C440 B.n248 VSUBS 0.007844f
C441 B.n249 VSUBS 0.007844f
C442 B.n250 VSUBS 0.007844f
C443 B.n251 VSUBS 0.007844f
C444 B.n252 VSUBS 0.007844f
C445 B.n253 VSUBS 0.007844f
C446 B.n254 VSUBS 0.007844f
C447 B.n255 VSUBS 0.007844f
C448 B.n256 VSUBS 0.007844f
C449 B.n257 VSUBS 0.007844f
C450 B.n258 VSUBS 0.007844f
C451 B.n259 VSUBS 0.007844f
C452 B.n260 VSUBS 0.007844f
C453 B.n261 VSUBS 0.007844f
C454 B.n262 VSUBS 0.007844f
C455 B.n263 VSUBS 0.007844f
C456 B.n264 VSUBS 0.007844f
C457 B.n265 VSUBS 0.007844f
C458 B.n266 VSUBS 0.007844f
C459 B.n267 VSUBS 0.007844f
C460 B.n268 VSUBS 0.007382f
C461 B.n269 VSUBS 0.018173f
C462 B.n270 VSUBS 0.004383f
C463 B.n271 VSUBS 0.007844f
C464 B.n272 VSUBS 0.007844f
C465 B.n273 VSUBS 0.007844f
C466 B.n274 VSUBS 0.007844f
C467 B.n275 VSUBS 0.007844f
C468 B.n276 VSUBS 0.007844f
C469 B.n277 VSUBS 0.007844f
C470 B.n278 VSUBS 0.007844f
C471 B.n279 VSUBS 0.007844f
C472 B.n280 VSUBS 0.007844f
C473 B.n281 VSUBS 0.007844f
C474 B.n282 VSUBS 0.007844f
C475 B.n283 VSUBS 0.004383f
C476 B.n284 VSUBS 0.007844f
C477 B.n285 VSUBS 0.007844f
C478 B.n286 VSUBS 0.007382f
C479 B.n287 VSUBS 0.007844f
C480 B.n288 VSUBS 0.007844f
C481 B.n289 VSUBS 0.007844f
C482 B.n290 VSUBS 0.007844f
C483 B.n291 VSUBS 0.007844f
C484 B.n292 VSUBS 0.007844f
C485 B.n293 VSUBS 0.007844f
C486 B.n294 VSUBS 0.007844f
C487 B.n295 VSUBS 0.007844f
C488 B.n296 VSUBS 0.007844f
C489 B.n297 VSUBS 0.007844f
C490 B.n298 VSUBS 0.007844f
C491 B.n299 VSUBS 0.007844f
C492 B.n300 VSUBS 0.007844f
C493 B.n301 VSUBS 0.007844f
C494 B.n302 VSUBS 0.007844f
C495 B.n303 VSUBS 0.007844f
C496 B.n304 VSUBS 0.007844f
C497 B.n305 VSUBS 0.007844f
C498 B.n306 VSUBS 0.007844f
C499 B.n307 VSUBS 0.007844f
C500 B.n308 VSUBS 0.007844f
C501 B.n309 VSUBS 0.007844f
C502 B.n310 VSUBS 0.007844f
C503 B.n311 VSUBS 0.007844f
C504 B.n312 VSUBS 0.007844f
C505 B.n313 VSUBS 0.007844f
C506 B.n314 VSUBS 0.007844f
C507 B.n315 VSUBS 0.007844f
C508 B.n316 VSUBS 0.007844f
C509 B.n317 VSUBS 0.007844f
C510 B.n318 VSUBS 0.020285f
C511 B.n319 VSUBS 0.020285f
C512 B.n320 VSUBS 0.019626f
C513 B.n321 VSUBS 0.007844f
C514 B.n322 VSUBS 0.007844f
C515 B.n323 VSUBS 0.007844f
C516 B.n324 VSUBS 0.007844f
C517 B.n325 VSUBS 0.007844f
C518 B.n326 VSUBS 0.007844f
C519 B.n327 VSUBS 0.007844f
C520 B.n328 VSUBS 0.007844f
C521 B.n329 VSUBS 0.007844f
C522 B.n330 VSUBS 0.007844f
C523 B.n331 VSUBS 0.007844f
C524 B.n332 VSUBS 0.007844f
C525 B.n333 VSUBS 0.007844f
C526 B.n334 VSUBS 0.007844f
C527 B.n335 VSUBS 0.007844f
C528 B.n336 VSUBS 0.007844f
C529 B.n337 VSUBS 0.007844f
C530 B.n338 VSUBS 0.007844f
C531 B.n339 VSUBS 0.007844f
C532 B.n340 VSUBS 0.007844f
C533 B.n341 VSUBS 0.007844f
C534 B.n342 VSUBS 0.007844f
C535 B.n343 VSUBS 0.007844f
C536 B.n344 VSUBS 0.007844f
C537 B.n345 VSUBS 0.007844f
C538 B.n346 VSUBS 0.007844f
C539 B.n347 VSUBS 0.007844f
C540 B.n348 VSUBS 0.007844f
C541 B.n349 VSUBS 0.007844f
C542 B.n350 VSUBS 0.007844f
C543 B.n351 VSUBS 0.007844f
C544 B.n352 VSUBS 0.007844f
C545 B.n353 VSUBS 0.007844f
C546 B.n354 VSUBS 0.007844f
C547 B.n355 VSUBS 0.007844f
C548 B.n356 VSUBS 0.007844f
C549 B.n357 VSUBS 0.007844f
C550 B.n358 VSUBS 0.007844f
C551 B.n359 VSUBS 0.007844f
C552 B.n360 VSUBS 0.007844f
C553 B.n361 VSUBS 0.007844f
C554 B.n362 VSUBS 0.007844f
C555 B.n363 VSUBS 0.007844f
C556 B.n364 VSUBS 0.007844f
C557 B.n365 VSUBS 0.007844f
C558 B.n366 VSUBS 0.007844f
C559 B.n367 VSUBS 0.007844f
C560 B.n368 VSUBS 0.007844f
C561 B.n369 VSUBS 0.007844f
C562 B.n370 VSUBS 0.007844f
C563 B.n371 VSUBS 0.007844f
C564 B.n372 VSUBS 0.007844f
C565 B.n373 VSUBS 0.007844f
C566 B.n374 VSUBS 0.007844f
C567 B.n375 VSUBS 0.007844f
C568 B.n376 VSUBS 0.007844f
C569 B.n377 VSUBS 0.007844f
C570 B.n378 VSUBS 0.007844f
C571 B.n379 VSUBS 0.007844f
C572 B.n380 VSUBS 0.007844f
C573 B.n381 VSUBS 0.007844f
C574 B.n382 VSUBS 0.007844f
C575 B.n383 VSUBS 0.007844f
C576 B.n384 VSUBS 0.007844f
C577 B.n385 VSUBS 0.007844f
C578 B.n386 VSUBS 0.007844f
C579 B.n387 VSUBS 0.007844f
C580 B.n388 VSUBS 0.007844f
C581 B.n389 VSUBS 0.007844f
C582 B.n390 VSUBS 0.007844f
C583 B.n391 VSUBS 0.007844f
C584 B.n392 VSUBS 0.007844f
C585 B.n393 VSUBS 0.007844f
C586 B.n394 VSUBS 0.007844f
C587 B.n395 VSUBS 0.007844f
C588 B.n396 VSUBS 0.007844f
C589 B.n397 VSUBS 0.007844f
C590 B.n398 VSUBS 0.007844f
C591 B.n399 VSUBS 0.007844f
C592 B.n400 VSUBS 0.007844f
C593 B.n401 VSUBS 0.007844f
C594 B.n402 VSUBS 0.007844f
C595 B.n403 VSUBS 0.007844f
C596 B.n404 VSUBS 0.007844f
C597 B.n405 VSUBS 0.007844f
C598 B.n406 VSUBS 0.007844f
C599 B.n407 VSUBS 0.007844f
C600 B.n408 VSUBS 0.007844f
C601 B.n409 VSUBS 0.007844f
C602 B.n410 VSUBS 0.007844f
C603 B.n411 VSUBS 0.007844f
C604 B.n412 VSUBS 0.007844f
C605 B.n413 VSUBS 0.007844f
C606 B.n414 VSUBS 0.007844f
C607 B.n415 VSUBS 0.007844f
C608 B.n416 VSUBS 0.007844f
C609 B.n417 VSUBS 0.007844f
C610 B.n418 VSUBS 0.007844f
C611 B.n419 VSUBS 0.007844f
C612 B.n420 VSUBS 0.007844f
C613 B.n421 VSUBS 0.007844f
C614 B.n422 VSUBS 0.007844f
C615 B.n423 VSUBS 0.007844f
C616 B.n424 VSUBS 0.007844f
C617 B.n425 VSUBS 0.007844f
C618 B.n426 VSUBS 0.007844f
C619 B.n427 VSUBS 0.007844f
C620 B.n428 VSUBS 0.007844f
C621 B.n429 VSUBS 0.007844f
C622 B.n430 VSUBS 0.007844f
C623 B.n431 VSUBS 0.007844f
C624 B.n432 VSUBS 0.007844f
C625 B.n433 VSUBS 0.007844f
C626 B.n434 VSUBS 0.007844f
C627 B.n435 VSUBS 0.007844f
C628 B.n436 VSUBS 0.007844f
C629 B.n437 VSUBS 0.007844f
C630 B.n438 VSUBS 0.007844f
C631 B.n439 VSUBS 0.007844f
C632 B.n440 VSUBS 0.007844f
C633 B.n441 VSUBS 0.007844f
C634 B.n442 VSUBS 0.007844f
C635 B.n443 VSUBS 0.007844f
C636 B.n444 VSUBS 0.007844f
C637 B.n445 VSUBS 0.007844f
C638 B.n446 VSUBS 0.007844f
C639 B.n447 VSUBS 0.007844f
C640 B.n448 VSUBS 0.007844f
C641 B.n449 VSUBS 0.007844f
C642 B.n450 VSUBS 0.007844f
C643 B.n451 VSUBS 0.007844f
C644 B.n452 VSUBS 0.007844f
C645 B.n453 VSUBS 0.007844f
C646 B.n454 VSUBS 0.007844f
C647 B.n455 VSUBS 0.007844f
C648 B.n456 VSUBS 0.007844f
C649 B.n457 VSUBS 0.007844f
C650 B.n458 VSUBS 0.007844f
C651 B.n459 VSUBS 0.007844f
C652 B.n460 VSUBS 0.007844f
C653 B.n461 VSUBS 0.007844f
C654 B.n462 VSUBS 0.007844f
C655 B.n463 VSUBS 0.007844f
C656 B.n464 VSUBS 0.019626f
C657 B.n465 VSUBS 0.020285f
C658 B.n466 VSUBS 0.019467f
C659 B.n467 VSUBS 0.007844f
C660 B.n468 VSUBS 0.007844f
C661 B.n469 VSUBS 0.007844f
C662 B.n470 VSUBS 0.007844f
C663 B.n471 VSUBS 0.007844f
C664 B.n472 VSUBS 0.007844f
C665 B.n473 VSUBS 0.007844f
C666 B.n474 VSUBS 0.007844f
C667 B.n475 VSUBS 0.007844f
C668 B.n476 VSUBS 0.007844f
C669 B.n477 VSUBS 0.007844f
C670 B.n478 VSUBS 0.007844f
C671 B.n479 VSUBS 0.007844f
C672 B.n480 VSUBS 0.007844f
C673 B.n481 VSUBS 0.007844f
C674 B.n482 VSUBS 0.007844f
C675 B.n483 VSUBS 0.007844f
C676 B.n484 VSUBS 0.007844f
C677 B.n485 VSUBS 0.007844f
C678 B.n486 VSUBS 0.007844f
C679 B.n487 VSUBS 0.007844f
C680 B.n488 VSUBS 0.007844f
C681 B.n489 VSUBS 0.007844f
C682 B.n490 VSUBS 0.007844f
C683 B.n491 VSUBS 0.007844f
C684 B.n492 VSUBS 0.007844f
C685 B.n493 VSUBS 0.007844f
C686 B.n494 VSUBS 0.007844f
C687 B.n495 VSUBS 0.007844f
C688 B.n496 VSUBS 0.007844f
C689 B.n497 VSUBS 0.007844f
C690 B.n498 VSUBS 0.007382f
C691 B.n499 VSUBS 0.007844f
C692 B.n500 VSUBS 0.007844f
C693 B.n501 VSUBS 0.007844f
C694 B.n502 VSUBS 0.007844f
C695 B.n503 VSUBS 0.007844f
C696 B.n504 VSUBS 0.007844f
C697 B.n505 VSUBS 0.007844f
C698 B.n506 VSUBS 0.007844f
C699 B.n507 VSUBS 0.007844f
C700 B.n508 VSUBS 0.007844f
C701 B.n509 VSUBS 0.007844f
C702 B.n510 VSUBS 0.007844f
C703 B.n511 VSUBS 0.007844f
C704 B.n512 VSUBS 0.007844f
C705 B.n513 VSUBS 0.007844f
C706 B.n514 VSUBS 0.004383f
C707 B.n515 VSUBS 0.018173f
C708 B.n516 VSUBS 0.007382f
C709 B.n517 VSUBS 0.007844f
C710 B.n518 VSUBS 0.007844f
C711 B.n519 VSUBS 0.007844f
C712 B.n520 VSUBS 0.007844f
C713 B.n521 VSUBS 0.007844f
C714 B.n522 VSUBS 0.007844f
C715 B.n523 VSUBS 0.007844f
C716 B.n524 VSUBS 0.007844f
C717 B.n525 VSUBS 0.007844f
C718 B.n526 VSUBS 0.007844f
C719 B.n527 VSUBS 0.007844f
C720 B.n528 VSUBS 0.007844f
C721 B.n529 VSUBS 0.007844f
C722 B.n530 VSUBS 0.007844f
C723 B.n531 VSUBS 0.007844f
C724 B.n532 VSUBS 0.007844f
C725 B.n533 VSUBS 0.007844f
C726 B.n534 VSUBS 0.007844f
C727 B.n535 VSUBS 0.007844f
C728 B.n536 VSUBS 0.007844f
C729 B.n537 VSUBS 0.007844f
C730 B.n538 VSUBS 0.007844f
C731 B.n539 VSUBS 0.007844f
C732 B.n540 VSUBS 0.007844f
C733 B.n541 VSUBS 0.007844f
C734 B.n542 VSUBS 0.007844f
C735 B.n543 VSUBS 0.007844f
C736 B.n544 VSUBS 0.007844f
C737 B.n545 VSUBS 0.007844f
C738 B.n546 VSUBS 0.007844f
C739 B.n547 VSUBS 0.007844f
C740 B.n548 VSUBS 0.007844f
C741 B.n549 VSUBS 0.020285f
C742 B.n550 VSUBS 0.019626f
C743 B.n551 VSUBS 0.019626f
C744 B.n552 VSUBS 0.007844f
C745 B.n553 VSUBS 0.007844f
C746 B.n554 VSUBS 0.007844f
C747 B.n555 VSUBS 0.007844f
C748 B.n556 VSUBS 0.007844f
C749 B.n557 VSUBS 0.007844f
C750 B.n558 VSUBS 0.007844f
C751 B.n559 VSUBS 0.007844f
C752 B.n560 VSUBS 0.007844f
C753 B.n561 VSUBS 0.007844f
C754 B.n562 VSUBS 0.007844f
C755 B.n563 VSUBS 0.007844f
C756 B.n564 VSUBS 0.007844f
C757 B.n565 VSUBS 0.007844f
C758 B.n566 VSUBS 0.007844f
C759 B.n567 VSUBS 0.007844f
C760 B.n568 VSUBS 0.007844f
C761 B.n569 VSUBS 0.007844f
C762 B.n570 VSUBS 0.007844f
C763 B.n571 VSUBS 0.007844f
C764 B.n572 VSUBS 0.007844f
C765 B.n573 VSUBS 0.007844f
C766 B.n574 VSUBS 0.007844f
C767 B.n575 VSUBS 0.007844f
C768 B.n576 VSUBS 0.007844f
C769 B.n577 VSUBS 0.007844f
C770 B.n578 VSUBS 0.007844f
C771 B.n579 VSUBS 0.007844f
C772 B.n580 VSUBS 0.007844f
C773 B.n581 VSUBS 0.007844f
C774 B.n582 VSUBS 0.007844f
C775 B.n583 VSUBS 0.007844f
C776 B.n584 VSUBS 0.007844f
C777 B.n585 VSUBS 0.007844f
C778 B.n586 VSUBS 0.007844f
C779 B.n587 VSUBS 0.007844f
C780 B.n588 VSUBS 0.007844f
C781 B.n589 VSUBS 0.007844f
C782 B.n590 VSUBS 0.007844f
C783 B.n591 VSUBS 0.007844f
C784 B.n592 VSUBS 0.007844f
C785 B.n593 VSUBS 0.007844f
C786 B.n594 VSUBS 0.007844f
C787 B.n595 VSUBS 0.007844f
C788 B.n596 VSUBS 0.007844f
C789 B.n597 VSUBS 0.007844f
C790 B.n598 VSUBS 0.007844f
C791 B.n599 VSUBS 0.007844f
C792 B.n600 VSUBS 0.007844f
C793 B.n601 VSUBS 0.007844f
C794 B.n602 VSUBS 0.007844f
C795 B.n603 VSUBS 0.007844f
C796 B.n604 VSUBS 0.007844f
C797 B.n605 VSUBS 0.007844f
C798 B.n606 VSUBS 0.007844f
C799 B.n607 VSUBS 0.007844f
C800 B.n608 VSUBS 0.007844f
C801 B.n609 VSUBS 0.007844f
C802 B.n610 VSUBS 0.007844f
C803 B.n611 VSUBS 0.007844f
C804 B.n612 VSUBS 0.007844f
C805 B.n613 VSUBS 0.007844f
C806 B.n614 VSUBS 0.007844f
C807 B.n615 VSUBS 0.007844f
C808 B.n616 VSUBS 0.007844f
C809 B.n617 VSUBS 0.007844f
C810 B.n618 VSUBS 0.007844f
C811 B.n619 VSUBS 0.007844f
C812 B.n620 VSUBS 0.007844f
C813 B.n621 VSUBS 0.007844f
C814 B.n622 VSUBS 0.007844f
C815 B.n623 VSUBS 0.017761f
C816 VDD1.n0 VSUBS 0.015112f
C817 VDD1.n1 VSUBS 0.034059f
C818 VDD1.n2 VSUBS 0.015257f
C819 VDD1.n3 VSUBS 0.026815f
C820 VDD1.n4 VSUBS 0.014409f
C821 VDD1.n5 VSUBS 0.034059f
C822 VDD1.n6 VSUBS 0.015257f
C823 VDD1.n7 VSUBS 0.591627f
C824 VDD1.n8 VSUBS 0.014409f
C825 VDD1.t8 VSUBS 0.07337f
C826 VDD1.n9 VSUBS 0.136804f
C827 VDD1.n10 VSUBS 0.02561f
C828 VDD1.n11 VSUBS 0.025544f
C829 VDD1.n12 VSUBS 0.034059f
C830 VDD1.n13 VSUBS 0.015257f
C831 VDD1.n14 VSUBS 0.014409f
C832 VDD1.n15 VSUBS 0.026815f
C833 VDD1.n16 VSUBS 0.026815f
C834 VDD1.n17 VSUBS 0.014409f
C835 VDD1.n18 VSUBS 0.015257f
C836 VDD1.n19 VSUBS 0.034059f
C837 VDD1.n20 VSUBS 0.034059f
C838 VDD1.n21 VSUBS 0.015257f
C839 VDD1.n22 VSUBS 0.014409f
C840 VDD1.n23 VSUBS 0.026815f
C841 VDD1.n24 VSUBS 0.068943f
C842 VDD1.n25 VSUBS 0.014409f
C843 VDD1.n26 VSUBS 0.015257f
C844 VDD1.n27 VSUBS 0.075488f
C845 VDD1.n28 VSUBS 0.077241f
C846 VDD1.t4 VSUBS 0.123539f
C847 VDD1.t3 VSUBS 0.123539f
C848 VDD1.n29 VSUBS 0.830973f
C849 VDD1.n30 VSUBS 0.844393f
C850 VDD1.n31 VSUBS 0.015112f
C851 VDD1.n32 VSUBS 0.034059f
C852 VDD1.n33 VSUBS 0.015257f
C853 VDD1.n34 VSUBS 0.026815f
C854 VDD1.n35 VSUBS 0.014409f
C855 VDD1.n36 VSUBS 0.034059f
C856 VDD1.n37 VSUBS 0.015257f
C857 VDD1.n38 VSUBS 0.591627f
C858 VDD1.n39 VSUBS 0.014409f
C859 VDD1.t9 VSUBS 0.07337f
C860 VDD1.n40 VSUBS 0.136804f
C861 VDD1.n41 VSUBS 0.02561f
C862 VDD1.n42 VSUBS 0.025544f
C863 VDD1.n43 VSUBS 0.034059f
C864 VDD1.n44 VSUBS 0.015257f
C865 VDD1.n45 VSUBS 0.014409f
C866 VDD1.n46 VSUBS 0.026815f
C867 VDD1.n47 VSUBS 0.026815f
C868 VDD1.n48 VSUBS 0.014409f
C869 VDD1.n49 VSUBS 0.015257f
C870 VDD1.n50 VSUBS 0.034059f
C871 VDD1.n51 VSUBS 0.034059f
C872 VDD1.n52 VSUBS 0.015257f
C873 VDD1.n53 VSUBS 0.014409f
C874 VDD1.n54 VSUBS 0.026815f
C875 VDD1.n55 VSUBS 0.068943f
C876 VDD1.n56 VSUBS 0.014409f
C877 VDD1.n57 VSUBS 0.015257f
C878 VDD1.n58 VSUBS 0.075488f
C879 VDD1.n59 VSUBS 0.077241f
C880 VDD1.t2 VSUBS 0.123539f
C881 VDD1.t5 VSUBS 0.123539f
C882 VDD1.n60 VSUBS 0.830971f
C883 VDD1.n61 VSUBS 0.836017f
C884 VDD1.t7 VSUBS 0.123539f
C885 VDD1.t0 VSUBS 0.123539f
C886 VDD1.n62 VSUBS 0.841414f
C887 VDD1.n63 VSUBS 2.64952f
C888 VDD1.t1 VSUBS 0.123539f
C889 VDD1.t6 VSUBS 0.123539f
C890 VDD1.n64 VSUBS 0.830968f
C891 VDD1.n65 VSUBS 2.78776f
C892 VTAIL.t6 VSUBS 0.149367f
C893 VTAIL.t5 VSUBS 0.149367f
C894 VTAIL.n0 VSUBS 0.900141f
C895 VTAIL.n1 VSUBS 0.87024f
C896 VTAIL.n2 VSUBS 0.018272f
C897 VTAIL.n3 VSUBS 0.041179f
C898 VTAIL.n4 VSUBS 0.018447f
C899 VTAIL.n5 VSUBS 0.032421f
C900 VTAIL.n6 VSUBS 0.017422f
C901 VTAIL.n7 VSUBS 0.041179f
C902 VTAIL.n8 VSUBS 0.018447f
C903 VTAIL.n9 VSUBS 0.715312f
C904 VTAIL.n10 VSUBS 0.017422f
C905 VTAIL.t13 VSUBS 0.088709f
C906 VTAIL.n11 VSUBS 0.165404f
C907 VTAIL.n12 VSUBS 0.030964f
C908 VTAIL.n13 VSUBS 0.030884f
C909 VTAIL.n14 VSUBS 0.041179f
C910 VTAIL.n15 VSUBS 0.018447f
C911 VTAIL.n16 VSUBS 0.017422f
C912 VTAIL.n17 VSUBS 0.032421f
C913 VTAIL.n18 VSUBS 0.032421f
C914 VTAIL.n19 VSUBS 0.017422f
C915 VTAIL.n20 VSUBS 0.018447f
C916 VTAIL.n21 VSUBS 0.041179f
C917 VTAIL.n22 VSUBS 0.041179f
C918 VTAIL.n23 VSUBS 0.018447f
C919 VTAIL.n24 VSUBS 0.017422f
C920 VTAIL.n25 VSUBS 0.032421f
C921 VTAIL.n26 VSUBS 0.083356f
C922 VTAIL.n27 VSUBS 0.017422f
C923 VTAIL.n28 VSUBS 0.018447f
C924 VTAIL.n29 VSUBS 0.09127f
C925 VTAIL.n30 VSUBS 0.061133f
C926 VTAIL.n31 VSUBS 0.38668f
C927 VTAIL.t16 VSUBS 0.149367f
C928 VTAIL.t15 VSUBS 0.149367f
C929 VTAIL.n32 VSUBS 0.900141f
C930 VTAIL.n33 VSUBS 0.968404f
C931 VTAIL.t11 VSUBS 0.149367f
C932 VTAIL.t14 VSUBS 0.149367f
C933 VTAIL.n34 VSUBS 0.900141f
C934 VTAIL.n35 VSUBS 2.13829f
C935 VTAIL.t19 VSUBS 0.149367f
C936 VTAIL.t8 VSUBS 0.149367f
C937 VTAIL.n36 VSUBS 0.900145f
C938 VTAIL.n37 VSUBS 2.13829f
C939 VTAIL.t2 VSUBS 0.149367f
C940 VTAIL.t3 VSUBS 0.149367f
C941 VTAIL.n38 VSUBS 0.900145f
C942 VTAIL.n39 VSUBS 0.968401f
C943 VTAIL.n40 VSUBS 0.018272f
C944 VTAIL.n41 VSUBS 0.041179f
C945 VTAIL.n42 VSUBS 0.018447f
C946 VTAIL.n43 VSUBS 0.032421f
C947 VTAIL.n44 VSUBS 0.017422f
C948 VTAIL.n45 VSUBS 0.041179f
C949 VTAIL.n46 VSUBS 0.018447f
C950 VTAIL.n47 VSUBS 0.715312f
C951 VTAIL.n48 VSUBS 0.017422f
C952 VTAIL.t1 VSUBS 0.088709f
C953 VTAIL.n49 VSUBS 0.165404f
C954 VTAIL.n50 VSUBS 0.030964f
C955 VTAIL.n51 VSUBS 0.030884f
C956 VTAIL.n52 VSUBS 0.041179f
C957 VTAIL.n53 VSUBS 0.018447f
C958 VTAIL.n54 VSUBS 0.017422f
C959 VTAIL.n55 VSUBS 0.032421f
C960 VTAIL.n56 VSUBS 0.032421f
C961 VTAIL.n57 VSUBS 0.017422f
C962 VTAIL.n58 VSUBS 0.018447f
C963 VTAIL.n59 VSUBS 0.041179f
C964 VTAIL.n60 VSUBS 0.041179f
C965 VTAIL.n61 VSUBS 0.018447f
C966 VTAIL.n62 VSUBS 0.017422f
C967 VTAIL.n63 VSUBS 0.032421f
C968 VTAIL.n64 VSUBS 0.083356f
C969 VTAIL.n65 VSUBS 0.017422f
C970 VTAIL.n66 VSUBS 0.018447f
C971 VTAIL.n67 VSUBS 0.09127f
C972 VTAIL.n68 VSUBS 0.061133f
C973 VTAIL.n69 VSUBS 0.38668f
C974 VTAIL.t12 VSUBS 0.149367f
C975 VTAIL.t10 VSUBS 0.149367f
C976 VTAIL.n70 VSUBS 0.900145f
C977 VTAIL.n71 VSUBS 0.915266f
C978 VTAIL.t18 VSUBS 0.149367f
C979 VTAIL.t9 VSUBS 0.149367f
C980 VTAIL.n72 VSUBS 0.900145f
C981 VTAIL.n73 VSUBS 0.968401f
C982 VTAIL.n74 VSUBS 0.018272f
C983 VTAIL.n75 VSUBS 0.041179f
C984 VTAIL.n76 VSUBS 0.018447f
C985 VTAIL.n77 VSUBS 0.032421f
C986 VTAIL.n78 VSUBS 0.017422f
C987 VTAIL.n79 VSUBS 0.041179f
C988 VTAIL.n80 VSUBS 0.018447f
C989 VTAIL.n81 VSUBS 0.715312f
C990 VTAIL.n82 VSUBS 0.017422f
C991 VTAIL.t17 VSUBS 0.088709f
C992 VTAIL.n83 VSUBS 0.165404f
C993 VTAIL.n84 VSUBS 0.030964f
C994 VTAIL.n85 VSUBS 0.030884f
C995 VTAIL.n86 VSUBS 0.041179f
C996 VTAIL.n87 VSUBS 0.018447f
C997 VTAIL.n88 VSUBS 0.017422f
C998 VTAIL.n89 VSUBS 0.032421f
C999 VTAIL.n90 VSUBS 0.032421f
C1000 VTAIL.n91 VSUBS 0.017422f
C1001 VTAIL.n92 VSUBS 0.018447f
C1002 VTAIL.n93 VSUBS 0.041179f
C1003 VTAIL.n94 VSUBS 0.041179f
C1004 VTAIL.n95 VSUBS 0.018447f
C1005 VTAIL.n96 VSUBS 0.017422f
C1006 VTAIL.n97 VSUBS 0.032421f
C1007 VTAIL.n98 VSUBS 0.083356f
C1008 VTAIL.n99 VSUBS 0.017422f
C1009 VTAIL.n100 VSUBS 0.018447f
C1010 VTAIL.n101 VSUBS 0.09127f
C1011 VTAIL.n102 VSUBS 0.061133f
C1012 VTAIL.n103 VSUBS 1.40527f
C1013 VTAIL.n104 VSUBS 0.018272f
C1014 VTAIL.n105 VSUBS 0.041179f
C1015 VTAIL.n106 VSUBS 0.018447f
C1016 VTAIL.n107 VSUBS 0.032421f
C1017 VTAIL.n108 VSUBS 0.017422f
C1018 VTAIL.n109 VSUBS 0.041179f
C1019 VTAIL.n110 VSUBS 0.018447f
C1020 VTAIL.n111 VSUBS 0.715312f
C1021 VTAIL.n112 VSUBS 0.017422f
C1022 VTAIL.t4 VSUBS 0.088709f
C1023 VTAIL.n113 VSUBS 0.165404f
C1024 VTAIL.n114 VSUBS 0.030964f
C1025 VTAIL.n115 VSUBS 0.030884f
C1026 VTAIL.n116 VSUBS 0.041179f
C1027 VTAIL.n117 VSUBS 0.018447f
C1028 VTAIL.n118 VSUBS 0.017422f
C1029 VTAIL.n119 VSUBS 0.032421f
C1030 VTAIL.n120 VSUBS 0.032421f
C1031 VTAIL.n121 VSUBS 0.017422f
C1032 VTAIL.n122 VSUBS 0.018447f
C1033 VTAIL.n123 VSUBS 0.041179f
C1034 VTAIL.n124 VSUBS 0.041179f
C1035 VTAIL.n125 VSUBS 0.018447f
C1036 VTAIL.n126 VSUBS 0.017422f
C1037 VTAIL.n127 VSUBS 0.032421f
C1038 VTAIL.n128 VSUBS 0.083356f
C1039 VTAIL.n129 VSUBS 0.017422f
C1040 VTAIL.n130 VSUBS 0.018447f
C1041 VTAIL.n131 VSUBS 0.09127f
C1042 VTAIL.n132 VSUBS 0.061133f
C1043 VTAIL.n133 VSUBS 1.40527f
C1044 VTAIL.t7 VSUBS 0.149367f
C1045 VTAIL.t0 VSUBS 0.149367f
C1046 VTAIL.n134 VSUBS 0.900141f
C1047 VTAIL.n135 VSUBS 0.808999f
C1048 VP.n0 VSUBS 0.041912f
C1049 VP.t9 VSUBS 1.25252f
C1050 VP.n1 VSUBS 0.039008f
C1051 VP.n2 VSUBS 0.041912f
C1052 VP.t2 VSUBS 1.25252f
C1053 VP.n3 VSUBS 0.073922f
C1054 VP.n4 VSUBS 0.041912f
C1055 VP.t4 VSUBS 1.25252f
C1056 VP.n5 VSUBS 0.081726f
C1057 VP.n6 VSUBS 0.041912f
C1058 VP.t7 VSUBS 1.25252f
C1059 VP.n7 VSUBS 0.481391f
C1060 VP.n8 VSUBS 0.041912f
C1061 VP.n9 VSUBS 0.084152f
C1062 VP.n10 VSUBS 0.041912f
C1063 VP.t3 VSUBS 1.25252f
C1064 VP.n11 VSUBS 0.039008f
C1065 VP.n12 VSUBS 0.041912f
C1066 VP.t8 VSUBS 1.25252f
C1067 VP.n13 VSUBS 0.073922f
C1068 VP.n14 VSUBS 0.041912f
C1069 VP.t6 VSUBS 1.25252f
C1070 VP.n15 VSUBS 0.081726f
C1071 VP.n16 VSUBS 0.041912f
C1072 VP.t5 VSUBS 1.25252f
C1073 VP.n17 VSUBS 0.580936f
C1074 VP.t1 VSUBS 1.46774f
C1075 VP.n18 VSUBS 0.576615f
C1076 VP.n19 VSUBS 0.312391f
C1077 VP.n20 VSUBS 0.060374f
C1078 VP.n21 VSUBS 0.073922f
C1079 VP.n22 VSUBS 0.044844f
C1080 VP.n23 VSUBS 0.041912f
C1081 VP.n24 VSUBS 0.041912f
C1082 VP.n25 VSUBS 0.041912f
C1083 VP.n26 VSUBS 0.52094f
C1084 VP.n27 VSUBS 0.081726f
C1085 VP.n28 VSUBS 0.044844f
C1086 VP.n29 VSUBS 0.041912f
C1087 VP.n30 VSUBS 0.041912f
C1088 VP.n31 VSUBS 0.041912f
C1089 VP.n32 VSUBS 0.060374f
C1090 VP.n33 VSUBS 0.481391f
C1091 VP.n34 VSUBS 0.057289f
C1092 VP.n35 VSUBS 0.077331f
C1093 VP.n36 VSUBS 0.041912f
C1094 VP.n37 VSUBS 0.041912f
C1095 VP.n38 VSUBS 0.041912f
C1096 VP.n39 VSUBS 0.084152f
C1097 VP.n40 VSUBS 0.042634f
C1098 VP.n41 VSUBS 0.582429f
C1099 VP.n42 VSUBS 1.93364f
C1100 VP.n43 VSUBS 1.9673f
C1101 VP.t0 VSUBS 1.25252f
C1102 VP.n44 VSUBS 0.582429f
C1103 VP.n45 VSUBS 0.042634f
C1104 VP.n46 VSUBS 0.041912f
C1105 VP.n47 VSUBS 0.041912f
C1106 VP.n48 VSUBS 0.041912f
C1107 VP.n49 VSUBS 0.039008f
C1108 VP.n50 VSUBS 0.077331f
C1109 VP.n51 VSUBS 0.057289f
C1110 VP.n52 VSUBS 0.041912f
C1111 VP.n53 VSUBS 0.041912f
C1112 VP.n54 VSUBS 0.060374f
C1113 VP.n55 VSUBS 0.073922f
C1114 VP.n56 VSUBS 0.044844f
C1115 VP.n57 VSUBS 0.041912f
C1116 VP.n58 VSUBS 0.041912f
C1117 VP.n59 VSUBS 0.041912f
C1118 VP.n60 VSUBS 0.52094f
C1119 VP.n61 VSUBS 0.081726f
C1120 VP.n62 VSUBS 0.044844f
C1121 VP.n63 VSUBS 0.041912f
C1122 VP.n64 VSUBS 0.041912f
C1123 VP.n65 VSUBS 0.041912f
C1124 VP.n66 VSUBS 0.060374f
C1125 VP.n67 VSUBS 0.481391f
C1126 VP.n68 VSUBS 0.057289f
C1127 VP.n69 VSUBS 0.077331f
C1128 VP.n70 VSUBS 0.041912f
C1129 VP.n71 VSUBS 0.041912f
C1130 VP.n72 VSUBS 0.041912f
C1131 VP.n73 VSUBS 0.084152f
C1132 VP.n74 VSUBS 0.042634f
C1133 VP.n75 VSUBS 0.582429f
C1134 VP.n76 VSUBS 0.046581f
.ends

