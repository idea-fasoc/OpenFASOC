* NGSPICE file created from diff_pair_sample_1271.ext - technology: sky130A

.subckt diff_pair_sample_1271 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=2.83
X1 VTAIL.t15 VP.t0 VDD1.t6 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X2 VTAIL.t2 VN.t0 VDD2.t7 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X3 B.t8 B.t6 B.t7 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=2.83
X4 VDD1.t0 VP.t1 VTAIL.t14 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X5 VDD2.t6 VN.t1 VTAIL.t5 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X6 VDD2.t5 VN.t2 VTAIL.t7 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=2.83
X7 VTAIL.t6 VN.t3 VDD2.t4 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X8 VTAIL.t4 VN.t4 VDD2.t3 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=2.83
X9 VDD1.t4 VP.t2 VTAIL.t13 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=2.83
X10 VTAIL.t12 VP.t3 VDD1.t1 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=2.83
X11 VDD2.t2 VN.t5 VTAIL.t1 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X12 VTAIL.t11 VP.t4 VDD1.t7 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X13 B.t5 B.t3 B.t4 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=2.83
X14 VDD2.t1 VN.t6 VTAIL.t3 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=2.83
X15 VDD1.t3 VP.t5 VTAIL.t10 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=2.83
X16 VTAIL.t0 VN.t7 VDD2.t0 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=2.83
X17 B.t2 B.t0 B.t1 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=2.83
X18 VDD1.t2 VP.t6 VTAIL.t9 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=2.94195 pd=18.16 as=2.94195 ps=18.16 w=17.83 l=2.83
X19 VTAIL.t8 VP.t7 VDD1.t5 w_n4130_n4534# sky130_fd_pr__pfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=2.83
R0 B.n518 B.n517 585
R1 B.n516 B.n153 585
R2 B.n515 B.n514 585
R3 B.n513 B.n154 585
R4 B.n512 B.n511 585
R5 B.n510 B.n155 585
R6 B.n509 B.n508 585
R7 B.n507 B.n156 585
R8 B.n506 B.n505 585
R9 B.n504 B.n157 585
R10 B.n503 B.n502 585
R11 B.n501 B.n158 585
R12 B.n500 B.n499 585
R13 B.n498 B.n159 585
R14 B.n497 B.n496 585
R15 B.n495 B.n160 585
R16 B.n494 B.n493 585
R17 B.n492 B.n161 585
R18 B.n491 B.n490 585
R19 B.n489 B.n162 585
R20 B.n488 B.n487 585
R21 B.n486 B.n163 585
R22 B.n485 B.n484 585
R23 B.n483 B.n164 585
R24 B.n482 B.n481 585
R25 B.n480 B.n165 585
R26 B.n479 B.n478 585
R27 B.n477 B.n166 585
R28 B.n476 B.n475 585
R29 B.n474 B.n167 585
R30 B.n473 B.n472 585
R31 B.n471 B.n168 585
R32 B.n470 B.n469 585
R33 B.n468 B.n169 585
R34 B.n467 B.n466 585
R35 B.n465 B.n170 585
R36 B.n464 B.n463 585
R37 B.n462 B.n171 585
R38 B.n461 B.n460 585
R39 B.n459 B.n172 585
R40 B.n458 B.n457 585
R41 B.n456 B.n173 585
R42 B.n455 B.n454 585
R43 B.n453 B.n174 585
R44 B.n452 B.n451 585
R45 B.n450 B.n175 585
R46 B.n449 B.n448 585
R47 B.n447 B.n176 585
R48 B.n446 B.n445 585
R49 B.n444 B.n177 585
R50 B.n443 B.n442 585
R51 B.n441 B.n178 585
R52 B.n440 B.n439 585
R53 B.n438 B.n179 585
R54 B.n437 B.n436 585
R55 B.n435 B.n180 585
R56 B.n434 B.n433 585
R57 B.n432 B.n181 585
R58 B.n431 B.n430 585
R59 B.n428 B.n182 585
R60 B.n427 B.n426 585
R61 B.n425 B.n185 585
R62 B.n424 B.n423 585
R63 B.n422 B.n186 585
R64 B.n421 B.n420 585
R65 B.n419 B.n187 585
R66 B.n418 B.n417 585
R67 B.n416 B.n188 585
R68 B.n414 B.n413 585
R69 B.n412 B.n191 585
R70 B.n411 B.n410 585
R71 B.n409 B.n192 585
R72 B.n408 B.n407 585
R73 B.n406 B.n193 585
R74 B.n405 B.n404 585
R75 B.n403 B.n194 585
R76 B.n402 B.n401 585
R77 B.n400 B.n195 585
R78 B.n399 B.n398 585
R79 B.n397 B.n196 585
R80 B.n396 B.n395 585
R81 B.n394 B.n197 585
R82 B.n393 B.n392 585
R83 B.n391 B.n198 585
R84 B.n390 B.n389 585
R85 B.n388 B.n199 585
R86 B.n387 B.n386 585
R87 B.n385 B.n200 585
R88 B.n384 B.n383 585
R89 B.n382 B.n201 585
R90 B.n381 B.n380 585
R91 B.n379 B.n202 585
R92 B.n378 B.n377 585
R93 B.n376 B.n203 585
R94 B.n375 B.n374 585
R95 B.n373 B.n204 585
R96 B.n372 B.n371 585
R97 B.n370 B.n205 585
R98 B.n369 B.n368 585
R99 B.n367 B.n206 585
R100 B.n366 B.n365 585
R101 B.n364 B.n207 585
R102 B.n363 B.n362 585
R103 B.n361 B.n208 585
R104 B.n360 B.n359 585
R105 B.n358 B.n209 585
R106 B.n357 B.n356 585
R107 B.n355 B.n210 585
R108 B.n354 B.n353 585
R109 B.n352 B.n211 585
R110 B.n351 B.n350 585
R111 B.n349 B.n212 585
R112 B.n348 B.n347 585
R113 B.n346 B.n213 585
R114 B.n345 B.n344 585
R115 B.n343 B.n214 585
R116 B.n342 B.n341 585
R117 B.n340 B.n215 585
R118 B.n339 B.n338 585
R119 B.n337 B.n216 585
R120 B.n336 B.n335 585
R121 B.n334 B.n217 585
R122 B.n333 B.n332 585
R123 B.n331 B.n218 585
R124 B.n330 B.n329 585
R125 B.n328 B.n219 585
R126 B.n327 B.n326 585
R127 B.n519 B.n152 585
R128 B.n521 B.n520 585
R129 B.n522 B.n151 585
R130 B.n524 B.n523 585
R131 B.n525 B.n150 585
R132 B.n527 B.n526 585
R133 B.n528 B.n149 585
R134 B.n530 B.n529 585
R135 B.n531 B.n148 585
R136 B.n533 B.n532 585
R137 B.n534 B.n147 585
R138 B.n536 B.n535 585
R139 B.n537 B.n146 585
R140 B.n539 B.n538 585
R141 B.n540 B.n145 585
R142 B.n542 B.n541 585
R143 B.n543 B.n144 585
R144 B.n545 B.n544 585
R145 B.n546 B.n143 585
R146 B.n548 B.n547 585
R147 B.n549 B.n142 585
R148 B.n551 B.n550 585
R149 B.n552 B.n141 585
R150 B.n554 B.n553 585
R151 B.n555 B.n140 585
R152 B.n557 B.n556 585
R153 B.n558 B.n139 585
R154 B.n560 B.n559 585
R155 B.n561 B.n138 585
R156 B.n563 B.n562 585
R157 B.n564 B.n137 585
R158 B.n566 B.n565 585
R159 B.n567 B.n136 585
R160 B.n569 B.n568 585
R161 B.n570 B.n135 585
R162 B.n572 B.n571 585
R163 B.n573 B.n134 585
R164 B.n575 B.n574 585
R165 B.n576 B.n133 585
R166 B.n578 B.n577 585
R167 B.n579 B.n132 585
R168 B.n581 B.n580 585
R169 B.n582 B.n131 585
R170 B.n584 B.n583 585
R171 B.n585 B.n130 585
R172 B.n587 B.n586 585
R173 B.n588 B.n129 585
R174 B.n590 B.n589 585
R175 B.n591 B.n128 585
R176 B.n593 B.n592 585
R177 B.n594 B.n127 585
R178 B.n596 B.n595 585
R179 B.n597 B.n126 585
R180 B.n599 B.n598 585
R181 B.n600 B.n125 585
R182 B.n602 B.n601 585
R183 B.n603 B.n124 585
R184 B.n605 B.n604 585
R185 B.n606 B.n123 585
R186 B.n608 B.n607 585
R187 B.n609 B.n122 585
R188 B.n611 B.n610 585
R189 B.n612 B.n121 585
R190 B.n614 B.n613 585
R191 B.n615 B.n120 585
R192 B.n617 B.n616 585
R193 B.n618 B.n119 585
R194 B.n620 B.n619 585
R195 B.n621 B.n118 585
R196 B.n623 B.n622 585
R197 B.n624 B.n117 585
R198 B.n626 B.n625 585
R199 B.n627 B.n116 585
R200 B.n629 B.n628 585
R201 B.n630 B.n115 585
R202 B.n632 B.n631 585
R203 B.n633 B.n114 585
R204 B.n635 B.n634 585
R205 B.n636 B.n113 585
R206 B.n638 B.n637 585
R207 B.n639 B.n112 585
R208 B.n641 B.n640 585
R209 B.n642 B.n111 585
R210 B.n644 B.n643 585
R211 B.n645 B.n110 585
R212 B.n647 B.n646 585
R213 B.n648 B.n109 585
R214 B.n650 B.n649 585
R215 B.n651 B.n108 585
R216 B.n653 B.n652 585
R217 B.n654 B.n107 585
R218 B.n656 B.n655 585
R219 B.n657 B.n106 585
R220 B.n659 B.n658 585
R221 B.n660 B.n105 585
R222 B.n662 B.n661 585
R223 B.n663 B.n104 585
R224 B.n665 B.n664 585
R225 B.n666 B.n103 585
R226 B.n668 B.n667 585
R227 B.n669 B.n102 585
R228 B.n671 B.n670 585
R229 B.n672 B.n101 585
R230 B.n674 B.n673 585
R231 B.n675 B.n100 585
R232 B.n677 B.n676 585
R233 B.n678 B.n99 585
R234 B.n680 B.n679 585
R235 B.n681 B.n98 585
R236 B.n683 B.n682 585
R237 B.n874 B.n29 585
R238 B.n873 B.n872 585
R239 B.n871 B.n30 585
R240 B.n870 B.n869 585
R241 B.n868 B.n31 585
R242 B.n867 B.n866 585
R243 B.n865 B.n32 585
R244 B.n864 B.n863 585
R245 B.n862 B.n33 585
R246 B.n861 B.n860 585
R247 B.n859 B.n34 585
R248 B.n858 B.n857 585
R249 B.n856 B.n35 585
R250 B.n855 B.n854 585
R251 B.n853 B.n36 585
R252 B.n852 B.n851 585
R253 B.n850 B.n37 585
R254 B.n849 B.n848 585
R255 B.n847 B.n38 585
R256 B.n846 B.n845 585
R257 B.n844 B.n39 585
R258 B.n843 B.n842 585
R259 B.n841 B.n40 585
R260 B.n840 B.n839 585
R261 B.n838 B.n41 585
R262 B.n837 B.n836 585
R263 B.n835 B.n42 585
R264 B.n834 B.n833 585
R265 B.n832 B.n43 585
R266 B.n831 B.n830 585
R267 B.n829 B.n44 585
R268 B.n828 B.n827 585
R269 B.n826 B.n45 585
R270 B.n825 B.n824 585
R271 B.n823 B.n46 585
R272 B.n822 B.n821 585
R273 B.n820 B.n47 585
R274 B.n819 B.n818 585
R275 B.n817 B.n48 585
R276 B.n816 B.n815 585
R277 B.n814 B.n49 585
R278 B.n813 B.n812 585
R279 B.n811 B.n50 585
R280 B.n810 B.n809 585
R281 B.n808 B.n51 585
R282 B.n807 B.n806 585
R283 B.n805 B.n52 585
R284 B.n804 B.n803 585
R285 B.n802 B.n53 585
R286 B.n801 B.n800 585
R287 B.n799 B.n54 585
R288 B.n798 B.n797 585
R289 B.n796 B.n55 585
R290 B.n795 B.n794 585
R291 B.n793 B.n56 585
R292 B.n792 B.n791 585
R293 B.n790 B.n57 585
R294 B.n789 B.n788 585
R295 B.n787 B.n58 585
R296 B.n786 B.n785 585
R297 B.n784 B.n59 585
R298 B.n783 B.n782 585
R299 B.n781 B.n63 585
R300 B.n780 B.n779 585
R301 B.n778 B.n64 585
R302 B.n777 B.n776 585
R303 B.n775 B.n65 585
R304 B.n774 B.n773 585
R305 B.n771 B.n66 585
R306 B.n770 B.n769 585
R307 B.n768 B.n69 585
R308 B.n767 B.n766 585
R309 B.n765 B.n70 585
R310 B.n764 B.n763 585
R311 B.n762 B.n71 585
R312 B.n761 B.n760 585
R313 B.n759 B.n72 585
R314 B.n758 B.n757 585
R315 B.n756 B.n73 585
R316 B.n755 B.n754 585
R317 B.n753 B.n74 585
R318 B.n752 B.n751 585
R319 B.n750 B.n75 585
R320 B.n749 B.n748 585
R321 B.n747 B.n76 585
R322 B.n746 B.n745 585
R323 B.n744 B.n77 585
R324 B.n743 B.n742 585
R325 B.n741 B.n78 585
R326 B.n740 B.n739 585
R327 B.n738 B.n79 585
R328 B.n737 B.n736 585
R329 B.n735 B.n80 585
R330 B.n734 B.n733 585
R331 B.n732 B.n81 585
R332 B.n731 B.n730 585
R333 B.n729 B.n82 585
R334 B.n728 B.n727 585
R335 B.n726 B.n83 585
R336 B.n725 B.n724 585
R337 B.n723 B.n84 585
R338 B.n722 B.n721 585
R339 B.n720 B.n85 585
R340 B.n719 B.n718 585
R341 B.n717 B.n86 585
R342 B.n716 B.n715 585
R343 B.n714 B.n87 585
R344 B.n713 B.n712 585
R345 B.n711 B.n88 585
R346 B.n710 B.n709 585
R347 B.n708 B.n89 585
R348 B.n707 B.n706 585
R349 B.n705 B.n90 585
R350 B.n704 B.n703 585
R351 B.n702 B.n91 585
R352 B.n701 B.n700 585
R353 B.n699 B.n92 585
R354 B.n698 B.n697 585
R355 B.n696 B.n93 585
R356 B.n695 B.n694 585
R357 B.n693 B.n94 585
R358 B.n692 B.n691 585
R359 B.n690 B.n95 585
R360 B.n689 B.n688 585
R361 B.n687 B.n96 585
R362 B.n686 B.n685 585
R363 B.n684 B.n97 585
R364 B.n876 B.n875 585
R365 B.n877 B.n28 585
R366 B.n879 B.n878 585
R367 B.n880 B.n27 585
R368 B.n882 B.n881 585
R369 B.n883 B.n26 585
R370 B.n885 B.n884 585
R371 B.n886 B.n25 585
R372 B.n888 B.n887 585
R373 B.n889 B.n24 585
R374 B.n891 B.n890 585
R375 B.n892 B.n23 585
R376 B.n894 B.n893 585
R377 B.n895 B.n22 585
R378 B.n897 B.n896 585
R379 B.n898 B.n21 585
R380 B.n900 B.n899 585
R381 B.n901 B.n20 585
R382 B.n903 B.n902 585
R383 B.n904 B.n19 585
R384 B.n906 B.n905 585
R385 B.n907 B.n18 585
R386 B.n909 B.n908 585
R387 B.n910 B.n17 585
R388 B.n912 B.n911 585
R389 B.n913 B.n16 585
R390 B.n915 B.n914 585
R391 B.n916 B.n15 585
R392 B.n918 B.n917 585
R393 B.n919 B.n14 585
R394 B.n921 B.n920 585
R395 B.n922 B.n13 585
R396 B.n924 B.n923 585
R397 B.n925 B.n12 585
R398 B.n927 B.n926 585
R399 B.n928 B.n11 585
R400 B.n930 B.n929 585
R401 B.n931 B.n10 585
R402 B.n933 B.n932 585
R403 B.n934 B.n9 585
R404 B.n936 B.n935 585
R405 B.n937 B.n8 585
R406 B.n939 B.n938 585
R407 B.n940 B.n7 585
R408 B.n942 B.n941 585
R409 B.n943 B.n6 585
R410 B.n945 B.n944 585
R411 B.n946 B.n5 585
R412 B.n948 B.n947 585
R413 B.n949 B.n4 585
R414 B.n951 B.n950 585
R415 B.n952 B.n3 585
R416 B.n954 B.n953 585
R417 B.n955 B.n0 585
R418 B.n2 B.n1 585
R419 B.n247 B.n246 585
R420 B.n249 B.n248 585
R421 B.n250 B.n245 585
R422 B.n252 B.n251 585
R423 B.n253 B.n244 585
R424 B.n255 B.n254 585
R425 B.n256 B.n243 585
R426 B.n258 B.n257 585
R427 B.n259 B.n242 585
R428 B.n261 B.n260 585
R429 B.n262 B.n241 585
R430 B.n264 B.n263 585
R431 B.n265 B.n240 585
R432 B.n267 B.n266 585
R433 B.n268 B.n239 585
R434 B.n270 B.n269 585
R435 B.n271 B.n238 585
R436 B.n273 B.n272 585
R437 B.n274 B.n237 585
R438 B.n276 B.n275 585
R439 B.n277 B.n236 585
R440 B.n279 B.n278 585
R441 B.n280 B.n235 585
R442 B.n282 B.n281 585
R443 B.n283 B.n234 585
R444 B.n285 B.n284 585
R445 B.n286 B.n233 585
R446 B.n288 B.n287 585
R447 B.n289 B.n232 585
R448 B.n291 B.n290 585
R449 B.n292 B.n231 585
R450 B.n294 B.n293 585
R451 B.n295 B.n230 585
R452 B.n297 B.n296 585
R453 B.n298 B.n229 585
R454 B.n300 B.n299 585
R455 B.n301 B.n228 585
R456 B.n303 B.n302 585
R457 B.n304 B.n227 585
R458 B.n306 B.n305 585
R459 B.n307 B.n226 585
R460 B.n309 B.n308 585
R461 B.n310 B.n225 585
R462 B.n312 B.n311 585
R463 B.n313 B.n224 585
R464 B.n315 B.n314 585
R465 B.n316 B.n223 585
R466 B.n318 B.n317 585
R467 B.n319 B.n222 585
R468 B.n321 B.n320 585
R469 B.n322 B.n221 585
R470 B.n324 B.n323 585
R471 B.n325 B.n220 585
R472 B.n327 B.n220 521.33
R473 B.n517 B.n152 521.33
R474 B.n684 B.n683 521.33
R475 B.n876 B.n29 521.33
R476 B.n189 B.t0 360.209
R477 B.n183 B.t3 360.209
R478 B.n67 B.t9 360.209
R479 B.n60 B.t6 360.209
R480 B.n957 B.n956 256.663
R481 B.n956 B.n955 235.042
R482 B.n956 B.n2 235.042
R483 B.n183 B.t4 170.415
R484 B.n67 B.t11 170.415
R485 B.n189 B.t1 170.392
R486 B.n60 B.t8 170.392
R487 B.n328 B.n327 163.367
R488 B.n329 B.n328 163.367
R489 B.n329 B.n218 163.367
R490 B.n333 B.n218 163.367
R491 B.n334 B.n333 163.367
R492 B.n335 B.n334 163.367
R493 B.n335 B.n216 163.367
R494 B.n339 B.n216 163.367
R495 B.n340 B.n339 163.367
R496 B.n341 B.n340 163.367
R497 B.n341 B.n214 163.367
R498 B.n345 B.n214 163.367
R499 B.n346 B.n345 163.367
R500 B.n347 B.n346 163.367
R501 B.n347 B.n212 163.367
R502 B.n351 B.n212 163.367
R503 B.n352 B.n351 163.367
R504 B.n353 B.n352 163.367
R505 B.n353 B.n210 163.367
R506 B.n357 B.n210 163.367
R507 B.n358 B.n357 163.367
R508 B.n359 B.n358 163.367
R509 B.n359 B.n208 163.367
R510 B.n363 B.n208 163.367
R511 B.n364 B.n363 163.367
R512 B.n365 B.n364 163.367
R513 B.n365 B.n206 163.367
R514 B.n369 B.n206 163.367
R515 B.n370 B.n369 163.367
R516 B.n371 B.n370 163.367
R517 B.n371 B.n204 163.367
R518 B.n375 B.n204 163.367
R519 B.n376 B.n375 163.367
R520 B.n377 B.n376 163.367
R521 B.n377 B.n202 163.367
R522 B.n381 B.n202 163.367
R523 B.n382 B.n381 163.367
R524 B.n383 B.n382 163.367
R525 B.n383 B.n200 163.367
R526 B.n387 B.n200 163.367
R527 B.n388 B.n387 163.367
R528 B.n389 B.n388 163.367
R529 B.n389 B.n198 163.367
R530 B.n393 B.n198 163.367
R531 B.n394 B.n393 163.367
R532 B.n395 B.n394 163.367
R533 B.n395 B.n196 163.367
R534 B.n399 B.n196 163.367
R535 B.n400 B.n399 163.367
R536 B.n401 B.n400 163.367
R537 B.n401 B.n194 163.367
R538 B.n405 B.n194 163.367
R539 B.n406 B.n405 163.367
R540 B.n407 B.n406 163.367
R541 B.n407 B.n192 163.367
R542 B.n411 B.n192 163.367
R543 B.n412 B.n411 163.367
R544 B.n413 B.n412 163.367
R545 B.n413 B.n188 163.367
R546 B.n418 B.n188 163.367
R547 B.n419 B.n418 163.367
R548 B.n420 B.n419 163.367
R549 B.n420 B.n186 163.367
R550 B.n424 B.n186 163.367
R551 B.n425 B.n424 163.367
R552 B.n426 B.n425 163.367
R553 B.n426 B.n182 163.367
R554 B.n431 B.n182 163.367
R555 B.n432 B.n431 163.367
R556 B.n433 B.n432 163.367
R557 B.n433 B.n180 163.367
R558 B.n437 B.n180 163.367
R559 B.n438 B.n437 163.367
R560 B.n439 B.n438 163.367
R561 B.n439 B.n178 163.367
R562 B.n443 B.n178 163.367
R563 B.n444 B.n443 163.367
R564 B.n445 B.n444 163.367
R565 B.n445 B.n176 163.367
R566 B.n449 B.n176 163.367
R567 B.n450 B.n449 163.367
R568 B.n451 B.n450 163.367
R569 B.n451 B.n174 163.367
R570 B.n455 B.n174 163.367
R571 B.n456 B.n455 163.367
R572 B.n457 B.n456 163.367
R573 B.n457 B.n172 163.367
R574 B.n461 B.n172 163.367
R575 B.n462 B.n461 163.367
R576 B.n463 B.n462 163.367
R577 B.n463 B.n170 163.367
R578 B.n467 B.n170 163.367
R579 B.n468 B.n467 163.367
R580 B.n469 B.n468 163.367
R581 B.n469 B.n168 163.367
R582 B.n473 B.n168 163.367
R583 B.n474 B.n473 163.367
R584 B.n475 B.n474 163.367
R585 B.n475 B.n166 163.367
R586 B.n479 B.n166 163.367
R587 B.n480 B.n479 163.367
R588 B.n481 B.n480 163.367
R589 B.n481 B.n164 163.367
R590 B.n485 B.n164 163.367
R591 B.n486 B.n485 163.367
R592 B.n487 B.n486 163.367
R593 B.n487 B.n162 163.367
R594 B.n491 B.n162 163.367
R595 B.n492 B.n491 163.367
R596 B.n493 B.n492 163.367
R597 B.n493 B.n160 163.367
R598 B.n497 B.n160 163.367
R599 B.n498 B.n497 163.367
R600 B.n499 B.n498 163.367
R601 B.n499 B.n158 163.367
R602 B.n503 B.n158 163.367
R603 B.n504 B.n503 163.367
R604 B.n505 B.n504 163.367
R605 B.n505 B.n156 163.367
R606 B.n509 B.n156 163.367
R607 B.n510 B.n509 163.367
R608 B.n511 B.n510 163.367
R609 B.n511 B.n154 163.367
R610 B.n515 B.n154 163.367
R611 B.n516 B.n515 163.367
R612 B.n517 B.n516 163.367
R613 B.n683 B.n98 163.367
R614 B.n679 B.n98 163.367
R615 B.n679 B.n678 163.367
R616 B.n678 B.n677 163.367
R617 B.n677 B.n100 163.367
R618 B.n673 B.n100 163.367
R619 B.n673 B.n672 163.367
R620 B.n672 B.n671 163.367
R621 B.n671 B.n102 163.367
R622 B.n667 B.n102 163.367
R623 B.n667 B.n666 163.367
R624 B.n666 B.n665 163.367
R625 B.n665 B.n104 163.367
R626 B.n661 B.n104 163.367
R627 B.n661 B.n660 163.367
R628 B.n660 B.n659 163.367
R629 B.n659 B.n106 163.367
R630 B.n655 B.n106 163.367
R631 B.n655 B.n654 163.367
R632 B.n654 B.n653 163.367
R633 B.n653 B.n108 163.367
R634 B.n649 B.n108 163.367
R635 B.n649 B.n648 163.367
R636 B.n648 B.n647 163.367
R637 B.n647 B.n110 163.367
R638 B.n643 B.n110 163.367
R639 B.n643 B.n642 163.367
R640 B.n642 B.n641 163.367
R641 B.n641 B.n112 163.367
R642 B.n637 B.n112 163.367
R643 B.n637 B.n636 163.367
R644 B.n636 B.n635 163.367
R645 B.n635 B.n114 163.367
R646 B.n631 B.n114 163.367
R647 B.n631 B.n630 163.367
R648 B.n630 B.n629 163.367
R649 B.n629 B.n116 163.367
R650 B.n625 B.n116 163.367
R651 B.n625 B.n624 163.367
R652 B.n624 B.n623 163.367
R653 B.n623 B.n118 163.367
R654 B.n619 B.n118 163.367
R655 B.n619 B.n618 163.367
R656 B.n618 B.n617 163.367
R657 B.n617 B.n120 163.367
R658 B.n613 B.n120 163.367
R659 B.n613 B.n612 163.367
R660 B.n612 B.n611 163.367
R661 B.n611 B.n122 163.367
R662 B.n607 B.n122 163.367
R663 B.n607 B.n606 163.367
R664 B.n606 B.n605 163.367
R665 B.n605 B.n124 163.367
R666 B.n601 B.n124 163.367
R667 B.n601 B.n600 163.367
R668 B.n600 B.n599 163.367
R669 B.n599 B.n126 163.367
R670 B.n595 B.n126 163.367
R671 B.n595 B.n594 163.367
R672 B.n594 B.n593 163.367
R673 B.n593 B.n128 163.367
R674 B.n589 B.n128 163.367
R675 B.n589 B.n588 163.367
R676 B.n588 B.n587 163.367
R677 B.n587 B.n130 163.367
R678 B.n583 B.n130 163.367
R679 B.n583 B.n582 163.367
R680 B.n582 B.n581 163.367
R681 B.n581 B.n132 163.367
R682 B.n577 B.n132 163.367
R683 B.n577 B.n576 163.367
R684 B.n576 B.n575 163.367
R685 B.n575 B.n134 163.367
R686 B.n571 B.n134 163.367
R687 B.n571 B.n570 163.367
R688 B.n570 B.n569 163.367
R689 B.n569 B.n136 163.367
R690 B.n565 B.n136 163.367
R691 B.n565 B.n564 163.367
R692 B.n564 B.n563 163.367
R693 B.n563 B.n138 163.367
R694 B.n559 B.n138 163.367
R695 B.n559 B.n558 163.367
R696 B.n558 B.n557 163.367
R697 B.n557 B.n140 163.367
R698 B.n553 B.n140 163.367
R699 B.n553 B.n552 163.367
R700 B.n552 B.n551 163.367
R701 B.n551 B.n142 163.367
R702 B.n547 B.n142 163.367
R703 B.n547 B.n546 163.367
R704 B.n546 B.n545 163.367
R705 B.n545 B.n144 163.367
R706 B.n541 B.n144 163.367
R707 B.n541 B.n540 163.367
R708 B.n540 B.n539 163.367
R709 B.n539 B.n146 163.367
R710 B.n535 B.n146 163.367
R711 B.n535 B.n534 163.367
R712 B.n534 B.n533 163.367
R713 B.n533 B.n148 163.367
R714 B.n529 B.n148 163.367
R715 B.n529 B.n528 163.367
R716 B.n528 B.n527 163.367
R717 B.n527 B.n150 163.367
R718 B.n523 B.n150 163.367
R719 B.n523 B.n522 163.367
R720 B.n522 B.n521 163.367
R721 B.n521 B.n152 163.367
R722 B.n872 B.n29 163.367
R723 B.n872 B.n871 163.367
R724 B.n871 B.n870 163.367
R725 B.n870 B.n31 163.367
R726 B.n866 B.n31 163.367
R727 B.n866 B.n865 163.367
R728 B.n865 B.n864 163.367
R729 B.n864 B.n33 163.367
R730 B.n860 B.n33 163.367
R731 B.n860 B.n859 163.367
R732 B.n859 B.n858 163.367
R733 B.n858 B.n35 163.367
R734 B.n854 B.n35 163.367
R735 B.n854 B.n853 163.367
R736 B.n853 B.n852 163.367
R737 B.n852 B.n37 163.367
R738 B.n848 B.n37 163.367
R739 B.n848 B.n847 163.367
R740 B.n847 B.n846 163.367
R741 B.n846 B.n39 163.367
R742 B.n842 B.n39 163.367
R743 B.n842 B.n841 163.367
R744 B.n841 B.n840 163.367
R745 B.n840 B.n41 163.367
R746 B.n836 B.n41 163.367
R747 B.n836 B.n835 163.367
R748 B.n835 B.n834 163.367
R749 B.n834 B.n43 163.367
R750 B.n830 B.n43 163.367
R751 B.n830 B.n829 163.367
R752 B.n829 B.n828 163.367
R753 B.n828 B.n45 163.367
R754 B.n824 B.n45 163.367
R755 B.n824 B.n823 163.367
R756 B.n823 B.n822 163.367
R757 B.n822 B.n47 163.367
R758 B.n818 B.n47 163.367
R759 B.n818 B.n817 163.367
R760 B.n817 B.n816 163.367
R761 B.n816 B.n49 163.367
R762 B.n812 B.n49 163.367
R763 B.n812 B.n811 163.367
R764 B.n811 B.n810 163.367
R765 B.n810 B.n51 163.367
R766 B.n806 B.n51 163.367
R767 B.n806 B.n805 163.367
R768 B.n805 B.n804 163.367
R769 B.n804 B.n53 163.367
R770 B.n800 B.n53 163.367
R771 B.n800 B.n799 163.367
R772 B.n799 B.n798 163.367
R773 B.n798 B.n55 163.367
R774 B.n794 B.n55 163.367
R775 B.n794 B.n793 163.367
R776 B.n793 B.n792 163.367
R777 B.n792 B.n57 163.367
R778 B.n788 B.n57 163.367
R779 B.n788 B.n787 163.367
R780 B.n787 B.n786 163.367
R781 B.n786 B.n59 163.367
R782 B.n782 B.n59 163.367
R783 B.n782 B.n781 163.367
R784 B.n781 B.n780 163.367
R785 B.n780 B.n64 163.367
R786 B.n776 B.n64 163.367
R787 B.n776 B.n775 163.367
R788 B.n775 B.n774 163.367
R789 B.n774 B.n66 163.367
R790 B.n769 B.n66 163.367
R791 B.n769 B.n768 163.367
R792 B.n768 B.n767 163.367
R793 B.n767 B.n70 163.367
R794 B.n763 B.n70 163.367
R795 B.n763 B.n762 163.367
R796 B.n762 B.n761 163.367
R797 B.n761 B.n72 163.367
R798 B.n757 B.n72 163.367
R799 B.n757 B.n756 163.367
R800 B.n756 B.n755 163.367
R801 B.n755 B.n74 163.367
R802 B.n751 B.n74 163.367
R803 B.n751 B.n750 163.367
R804 B.n750 B.n749 163.367
R805 B.n749 B.n76 163.367
R806 B.n745 B.n76 163.367
R807 B.n745 B.n744 163.367
R808 B.n744 B.n743 163.367
R809 B.n743 B.n78 163.367
R810 B.n739 B.n78 163.367
R811 B.n739 B.n738 163.367
R812 B.n738 B.n737 163.367
R813 B.n737 B.n80 163.367
R814 B.n733 B.n80 163.367
R815 B.n733 B.n732 163.367
R816 B.n732 B.n731 163.367
R817 B.n731 B.n82 163.367
R818 B.n727 B.n82 163.367
R819 B.n727 B.n726 163.367
R820 B.n726 B.n725 163.367
R821 B.n725 B.n84 163.367
R822 B.n721 B.n84 163.367
R823 B.n721 B.n720 163.367
R824 B.n720 B.n719 163.367
R825 B.n719 B.n86 163.367
R826 B.n715 B.n86 163.367
R827 B.n715 B.n714 163.367
R828 B.n714 B.n713 163.367
R829 B.n713 B.n88 163.367
R830 B.n709 B.n88 163.367
R831 B.n709 B.n708 163.367
R832 B.n708 B.n707 163.367
R833 B.n707 B.n90 163.367
R834 B.n703 B.n90 163.367
R835 B.n703 B.n702 163.367
R836 B.n702 B.n701 163.367
R837 B.n701 B.n92 163.367
R838 B.n697 B.n92 163.367
R839 B.n697 B.n696 163.367
R840 B.n696 B.n695 163.367
R841 B.n695 B.n94 163.367
R842 B.n691 B.n94 163.367
R843 B.n691 B.n690 163.367
R844 B.n690 B.n689 163.367
R845 B.n689 B.n96 163.367
R846 B.n685 B.n96 163.367
R847 B.n685 B.n684 163.367
R848 B.n877 B.n876 163.367
R849 B.n878 B.n877 163.367
R850 B.n878 B.n27 163.367
R851 B.n882 B.n27 163.367
R852 B.n883 B.n882 163.367
R853 B.n884 B.n883 163.367
R854 B.n884 B.n25 163.367
R855 B.n888 B.n25 163.367
R856 B.n889 B.n888 163.367
R857 B.n890 B.n889 163.367
R858 B.n890 B.n23 163.367
R859 B.n894 B.n23 163.367
R860 B.n895 B.n894 163.367
R861 B.n896 B.n895 163.367
R862 B.n896 B.n21 163.367
R863 B.n900 B.n21 163.367
R864 B.n901 B.n900 163.367
R865 B.n902 B.n901 163.367
R866 B.n902 B.n19 163.367
R867 B.n906 B.n19 163.367
R868 B.n907 B.n906 163.367
R869 B.n908 B.n907 163.367
R870 B.n908 B.n17 163.367
R871 B.n912 B.n17 163.367
R872 B.n913 B.n912 163.367
R873 B.n914 B.n913 163.367
R874 B.n914 B.n15 163.367
R875 B.n918 B.n15 163.367
R876 B.n919 B.n918 163.367
R877 B.n920 B.n919 163.367
R878 B.n920 B.n13 163.367
R879 B.n924 B.n13 163.367
R880 B.n925 B.n924 163.367
R881 B.n926 B.n925 163.367
R882 B.n926 B.n11 163.367
R883 B.n930 B.n11 163.367
R884 B.n931 B.n930 163.367
R885 B.n932 B.n931 163.367
R886 B.n932 B.n9 163.367
R887 B.n936 B.n9 163.367
R888 B.n937 B.n936 163.367
R889 B.n938 B.n937 163.367
R890 B.n938 B.n7 163.367
R891 B.n942 B.n7 163.367
R892 B.n943 B.n942 163.367
R893 B.n944 B.n943 163.367
R894 B.n944 B.n5 163.367
R895 B.n948 B.n5 163.367
R896 B.n949 B.n948 163.367
R897 B.n950 B.n949 163.367
R898 B.n950 B.n3 163.367
R899 B.n954 B.n3 163.367
R900 B.n955 B.n954 163.367
R901 B.n246 B.n2 163.367
R902 B.n249 B.n246 163.367
R903 B.n250 B.n249 163.367
R904 B.n251 B.n250 163.367
R905 B.n251 B.n244 163.367
R906 B.n255 B.n244 163.367
R907 B.n256 B.n255 163.367
R908 B.n257 B.n256 163.367
R909 B.n257 B.n242 163.367
R910 B.n261 B.n242 163.367
R911 B.n262 B.n261 163.367
R912 B.n263 B.n262 163.367
R913 B.n263 B.n240 163.367
R914 B.n267 B.n240 163.367
R915 B.n268 B.n267 163.367
R916 B.n269 B.n268 163.367
R917 B.n269 B.n238 163.367
R918 B.n273 B.n238 163.367
R919 B.n274 B.n273 163.367
R920 B.n275 B.n274 163.367
R921 B.n275 B.n236 163.367
R922 B.n279 B.n236 163.367
R923 B.n280 B.n279 163.367
R924 B.n281 B.n280 163.367
R925 B.n281 B.n234 163.367
R926 B.n285 B.n234 163.367
R927 B.n286 B.n285 163.367
R928 B.n287 B.n286 163.367
R929 B.n287 B.n232 163.367
R930 B.n291 B.n232 163.367
R931 B.n292 B.n291 163.367
R932 B.n293 B.n292 163.367
R933 B.n293 B.n230 163.367
R934 B.n297 B.n230 163.367
R935 B.n298 B.n297 163.367
R936 B.n299 B.n298 163.367
R937 B.n299 B.n228 163.367
R938 B.n303 B.n228 163.367
R939 B.n304 B.n303 163.367
R940 B.n305 B.n304 163.367
R941 B.n305 B.n226 163.367
R942 B.n309 B.n226 163.367
R943 B.n310 B.n309 163.367
R944 B.n311 B.n310 163.367
R945 B.n311 B.n224 163.367
R946 B.n315 B.n224 163.367
R947 B.n316 B.n315 163.367
R948 B.n317 B.n316 163.367
R949 B.n317 B.n222 163.367
R950 B.n321 B.n222 163.367
R951 B.n322 B.n321 163.367
R952 B.n323 B.n322 163.367
R953 B.n323 B.n220 163.367
R954 B.n184 B.t5 109.13
R955 B.n68 B.t10 109.13
R956 B.n190 B.t2 109.108
R957 B.n61 B.t7 109.108
R958 B.n190 B.n189 61.2853
R959 B.n184 B.n183 61.2853
R960 B.n68 B.n67 61.2853
R961 B.n61 B.n60 61.2853
R962 B.n415 B.n190 59.5399
R963 B.n429 B.n184 59.5399
R964 B.n772 B.n68 59.5399
R965 B.n62 B.n61 59.5399
R966 B.n875 B.n874 33.8737
R967 B.n682 B.n97 33.8737
R968 B.n519 B.n518 33.8737
R969 B.n326 B.n325 33.8737
R970 B B.n957 18.0485
R971 B.n875 B.n28 10.6151
R972 B.n879 B.n28 10.6151
R973 B.n880 B.n879 10.6151
R974 B.n881 B.n880 10.6151
R975 B.n881 B.n26 10.6151
R976 B.n885 B.n26 10.6151
R977 B.n886 B.n885 10.6151
R978 B.n887 B.n886 10.6151
R979 B.n887 B.n24 10.6151
R980 B.n891 B.n24 10.6151
R981 B.n892 B.n891 10.6151
R982 B.n893 B.n892 10.6151
R983 B.n893 B.n22 10.6151
R984 B.n897 B.n22 10.6151
R985 B.n898 B.n897 10.6151
R986 B.n899 B.n898 10.6151
R987 B.n899 B.n20 10.6151
R988 B.n903 B.n20 10.6151
R989 B.n904 B.n903 10.6151
R990 B.n905 B.n904 10.6151
R991 B.n905 B.n18 10.6151
R992 B.n909 B.n18 10.6151
R993 B.n910 B.n909 10.6151
R994 B.n911 B.n910 10.6151
R995 B.n911 B.n16 10.6151
R996 B.n915 B.n16 10.6151
R997 B.n916 B.n915 10.6151
R998 B.n917 B.n916 10.6151
R999 B.n917 B.n14 10.6151
R1000 B.n921 B.n14 10.6151
R1001 B.n922 B.n921 10.6151
R1002 B.n923 B.n922 10.6151
R1003 B.n923 B.n12 10.6151
R1004 B.n927 B.n12 10.6151
R1005 B.n928 B.n927 10.6151
R1006 B.n929 B.n928 10.6151
R1007 B.n929 B.n10 10.6151
R1008 B.n933 B.n10 10.6151
R1009 B.n934 B.n933 10.6151
R1010 B.n935 B.n934 10.6151
R1011 B.n935 B.n8 10.6151
R1012 B.n939 B.n8 10.6151
R1013 B.n940 B.n939 10.6151
R1014 B.n941 B.n940 10.6151
R1015 B.n941 B.n6 10.6151
R1016 B.n945 B.n6 10.6151
R1017 B.n946 B.n945 10.6151
R1018 B.n947 B.n946 10.6151
R1019 B.n947 B.n4 10.6151
R1020 B.n951 B.n4 10.6151
R1021 B.n952 B.n951 10.6151
R1022 B.n953 B.n952 10.6151
R1023 B.n953 B.n0 10.6151
R1024 B.n874 B.n873 10.6151
R1025 B.n873 B.n30 10.6151
R1026 B.n869 B.n30 10.6151
R1027 B.n869 B.n868 10.6151
R1028 B.n868 B.n867 10.6151
R1029 B.n867 B.n32 10.6151
R1030 B.n863 B.n32 10.6151
R1031 B.n863 B.n862 10.6151
R1032 B.n862 B.n861 10.6151
R1033 B.n861 B.n34 10.6151
R1034 B.n857 B.n34 10.6151
R1035 B.n857 B.n856 10.6151
R1036 B.n856 B.n855 10.6151
R1037 B.n855 B.n36 10.6151
R1038 B.n851 B.n36 10.6151
R1039 B.n851 B.n850 10.6151
R1040 B.n850 B.n849 10.6151
R1041 B.n849 B.n38 10.6151
R1042 B.n845 B.n38 10.6151
R1043 B.n845 B.n844 10.6151
R1044 B.n844 B.n843 10.6151
R1045 B.n843 B.n40 10.6151
R1046 B.n839 B.n40 10.6151
R1047 B.n839 B.n838 10.6151
R1048 B.n838 B.n837 10.6151
R1049 B.n837 B.n42 10.6151
R1050 B.n833 B.n42 10.6151
R1051 B.n833 B.n832 10.6151
R1052 B.n832 B.n831 10.6151
R1053 B.n831 B.n44 10.6151
R1054 B.n827 B.n44 10.6151
R1055 B.n827 B.n826 10.6151
R1056 B.n826 B.n825 10.6151
R1057 B.n825 B.n46 10.6151
R1058 B.n821 B.n46 10.6151
R1059 B.n821 B.n820 10.6151
R1060 B.n820 B.n819 10.6151
R1061 B.n819 B.n48 10.6151
R1062 B.n815 B.n48 10.6151
R1063 B.n815 B.n814 10.6151
R1064 B.n814 B.n813 10.6151
R1065 B.n813 B.n50 10.6151
R1066 B.n809 B.n50 10.6151
R1067 B.n809 B.n808 10.6151
R1068 B.n808 B.n807 10.6151
R1069 B.n807 B.n52 10.6151
R1070 B.n803 B.n52 10.6151
R1071 B.n803 B.n802 10.6151
R1072 B.n802 B.n801 10.6151
R1073 B.n801 B.n54 10.6151
R1074 B.n797 B.n54 10.6151
R1075 B.n797 B.n796 10.6151
R1076 B.n796 B.n795 10.6151
R1077 B.n795 B.n56 10.6151
R1078 B.n791 B.n56 10.6151
R1079 B.n791 B.n790 10.6151
R1080 B.n790 B.n789 10.6151
R1081 B.n789 B.n58 10.6151
R1082 B.n785 B.n784 10.6151
R1083 B.n784 B.n783 10.6151
R1084 B.n783 B.n63 10.6151
R1085 B.n779 B.n63 10.6151
R1086 B.n779 B.n778 10.6151
R1087 B.n778 B.n777 10.6151
R1088 B.n777 B.n65 10.6151
R1089 B.n773 B.n65 10.6151
R1090 B.n771 B.n770 10.6151
R1091 B.n770 B.n69 10.6151
R1092 B.n766 B.n69 10.6151
R1093 B.n766 B.n765 10.6151
R1094 B.n765 B.n764 10.6151
R1095 B.n764 B.n71 10.6151
R1096 B.n760 B.n71 10.6151
R1097 B.n760 B.n759 10.6151
R1098 B.n759 B.n758 10.6151
R1099 B.n758 B.n73 10.6151
R1100 B.n754 B.n73 10.6151
R1101 B.n754 B.n753 10.6151
R1102 B.n753 B.n752 10.6151
R1103 B.n752 B.n75 10.6151
R1104 B.n748 B.n75 10.6151
R1105 B.n748 B.n747 10.6151
R1106 B.n747 B.n746 10.6151
R1107 B.n746 B.n77 10.6151
R1108 B.n742 B.n77 10.6151
R1109 B.n742 B.n741 10.6151
R1110 B.n741 B.n740 10.6151
R1111 B.n740 B.n79 10.6151
R1112 B.n736 B.n79 10.6151
R1113 B.n736 B.n735 10.6151
R1114 B.n735 B.n734 10.6151
R1115 B.n734 B.n81 10.6151
R1116 B.n730 B.n81 10.6151
R1117 B.n730 B.n729 10.6151
R1118 B.n729 B.n728 10.6151
R1119 B.n728 B.n83 10.6151
R1120 B.n724 B.n83 10.6151
R1121 B.n724 B.n723 10.6151
R1122 B.n723 B.n722 10.6151
R1123 B.n722 B.n85 10.6151
R1124 B.n718 B.n85 10.6151
R1125 B.n718 B.n717 10.6151
R1126 B.n717 B.n716 10.6151
R1127 B.n716 B.n87 10.6151
R1128 B.n712 B.n87 10.6151
R1129 B.n712 B.n711 10.6151
R1130 B.n711 B.n710 10.6151
R1131 B.n710 B.n89 10.6151
R1132 B.n706 B.n89 10.6151
R1133 B.n706 B.n705 10.6151
R1134 B.n705 B.n704 10.6151
R1135 B.n704 B.n91 10.6151
R1136 B.n700 B.n91 10.6151
R1137 B.n700 B.n699 10.6151
R1138 B.n699 B.n698 10.6151
R1139 B.n698 B.n93 10.6151
R1140 B.n694 B.n93 10.6151
R1141 B.n694 B.n693 10.6151
R1142 B.n693 B.n692 10.6151
R1143 B.n692 B.n95 10.6151
R1144 B.n688 B.n95 10.6151
R1145 B.n688 B.n687 10.6151
R1146 B.n687 B.n686 10.6151
R1147 B.n686 B.n97 10.6151
R1148 B.n682 B.n681 10.6151
R1149 B.n681 B.n680 10.6151
R1150 B.n680 B.n99 10.6151
R1151 B.n676 B.n99 10.6151
R1152 B.n676 B.n675 10.6151
R1153 B.n675 B.n674 10.6151
R1154 B.n674 B.n101 10.6151
R1155 B.n670 B.n101 10.6151
R1156 B.n670 B.n669 10.6151
R1157 B.n669 B.n668 10.6151
R1158 B.n668 B.n103 10.6151
R1159 B.n664 B.n103 10.6151
R1160 B.n664 B.n663 10.6151
R1161 B.n663 B.n662 10.6151
R1162 B.n662 B.n105 10.6151
R1163 B.n658 B.n105 10.6151
R1164 B.n658 B.n657 10.6151
R1165 B.n657 B.n656 10.6151
R1166 B.n656 B.n107 10.6151
R1167 B.n652 B.n107 10.6151
R1168 B.n652 B.n651 10.6151
R1169 B.n651 B.n650 10.6151
R1170 B.n650 B.n109 10.6151
R1171 B.n646 B.n109 10.6151
R1172 B.n646 B.n645 10.6151
R1173 B.n645 B.n644 10.6151
R1174 B.n644 B.n111 10.6151
R1175 B.n640 B.n111 10.6151
R1176 B.n640 B.n639 10.6151
R1177 B.n639 B.n638 10.6151
R1178 B.n638 B.n113 10.6151
R1179 B.n634 B.n113 10.6151
R1180 B.n634 B.n633 10.6151
R1181 B.n633 B.n632 10.6151
R1182 B.n632 B.n115 10.6151
R1183 B.n628 B.n115 10.6151
R1184 B.n628 B.n627 10.6151
R1185 B.n627 B.n626 10.6151
R1186 B.n626 B.n117 10.6151
R1187 B.n622 B.n117 10.6151
R1188 B.n622 B.n621 10.6151
R1189 B.n621 B.n620 10.6151
R1190 B.n620 B.n119 10.6151
R1191 B.n616 B.n119 10.6151
R1192 B.n616 B.n615 10.6151
R1193 B.n615 B.n614 10.6151
R1194 B.n614 B.n121 10.6151
R1195 B.n610 B.n121 10.6151
R1196 B.n610 B.n609 10.6151
R1197 B.n609 B.n608 10.6151
R1198 B.n608 B.n123 10.6151
R1199 B.n604 B.n123 10.6151
R1200 B.n604 B.n603 10.6151
R1201 B.n603 B.n602 10.6151
R1202 B.n602 B.n125 10.6151
R1203 B.n598 B.n125 10.6151
R1204 B.n598 B.n597 10.6151
R1205 B.n597 B.n596 10.6151
R1206 B.n596 B.n127 10.6151
R1207 B.n592 B.n127 10.6151
R1208 B.n592 B.n591 10.6151
R1209 B.n591 B.n590 10.6151
R1210 B.n590 B.n129 10.6151
R1211 B.n586 B.n129 10.6151
R1212 B.n586 B.n585 10.6151
R1213 B.n585 B.n584 10.6151
R1214 B.n584 B.n131 10.6151
R1215 B.n580 B.n131 10.6151
R1216 B.n580 B.n579 10.6151
R1217 B.n579 B.n578 10.6151
R1218 B.n578 B.n133 10.6151
R1219 B.n574 B.n133 10.6151
R1220 B.n574 B.n573 10.6151
R1221 B.n573 B.n572 10.6151
R1222 B.n572 B.n135 10.6151
R1223 B.n568 B.n135 10.6151
R1224 B.n568 B.n567 10.6151
R1225 B.n567 B.n566 10.6151
R1226 B.n566 B.n137 10.6151
R1227 B.n562 B.n137 10.6151
R1228 B.n562 B.n561 10.6151
R1229 B.n561 B.n560 10.6151
R1230 B.n560 B.n139 10.6151
R1231 B.n556 B.n139 10.6151
R1232 B.n556 B.n555 10.6151
R1233 B.n555 B.n554 10.6151
R1234 B.n554 B.n141 10.6151
R1235 B.n550 B.n141 10.6151
R1236 B.n550 B.n549 10.6151
R1237 B.n549 B.n548 10.6151
R1238 B.n548 B.n143 10.6151
R1239 B.n544 B.n143 10.6151
R1240 B.n544 B.n543 10.6151
R1241 B.n543 B.n542 10.6151
R1242 B.n542 B.n145 10.6151
R1243 B.n538 B.n145 10.6151
R1244 B.n538 B.n537 10.6151
R1245 B.n537 B.n536 10.6151
R1246 B.n536 B.n147 10.6151
R1247 B.n532 B.n147 10.6151
R1248 B.n532 B.n531 10.6151
R1249 B.n531 B.n530 10.6151
R1250 B.n530 B.n149 10.6151
R1251 B.n526 B.n149 10.6151
R1252 B.n526 B.n525 10.6151
R1253 B.n525 B.n524 10.6151
R1254 B.n524 B.n151 10.6151
R1255 B.n520 B.n151 10.6151
R1256 B.n520 B.n519 10.6151
R1257 B.n247 B.n1 10.6151
R1258 B.n248 B.n247 10.6151
R1259 B.n248 B.n245 10.6151
R1260 B.n252 B.n245 10.6151
R1261 B.n253 B.n252 10.6151
R1262 B.n254 B.n253 10.6151
R1263 B.n254 B.n243 10.6151
R1264 B.n258 B.n243 10.6151
R1265 B.n259 B.n258 10.6151
R1266 B.n260 B.n259 10.6151
R1267 B.n260 B.n241 10.6151
R1268 B.n264 B.n241 10.6151
R1269 B.n265 B.n264 10.6151
R1270 B.n266 B.n265 10.6151
R1271 B.n266 B.n239 10.6151
R1272 B.n270 B.n239 10.6151
R1273 B.n271 B.n270 10.6151
R1274 B.n272 B.n271 10.6151
R1275 B.n272 B.n237 10.6151
R1276 B.n276 B.n237 10.6151
R1277 B.n277 B.n276 10.6151
R1278 B.n278 B.n277 10.6151
R1279 B.n278 B.n235 10.6151
R1280 B.n282 B.n235 10.6151
R1281 B.n283 B.n282 10.6151
R1282 B.n284 B.n283 10.6151
R1283 B.n284 B.n233 10.6151
R1284 B.n288 B.n233 10.6151
R1285 B.n289 B.n288 10.6151
R1286 B.n290 B.n289 10.6151
R1287 B.n290 B.n231 10.6151
R1288 B.n294 B.n231 10.6151
R1289 B.n295 B.n294 10.6151
R1290 B.n296 B.n295 10.6151
R1291 B.n296 B.n229 10.6151
R1292 B.n300 B.n229 10.6151
R1293 B.n301 B.n300 10.6151
R1294 B.n302 B.n301 10.6151
R1295 B.n302 B.n227 10.6151
R1296 B.n306 B.n227 10.6151
R1297 B.n307 B.n306 10.6151
R1298 B.n308 B.n307 10.6151
R1299 B.n308 B.n225 10.6151
R1300 B.n312 B.n225 10.6151
R1301 B.n313 B.n312 10.6151
R1302 B.n314 B.n313 10.6151
R1303 B.n314 B.n223 10.6151
R1304 B.n318 B.n223 10.6151
R1305 B.n319 B.n318 10.6151
R1306 B.n320 B.n319 10.6151
R1307 B.n320 B.n221 10.6151
R1308 B.n324 B.n221 10.6151
R1309 B.n325 B.n324 10.6151
R1310 B.n326 B.n219 10.6151
R1311 B.n330 B.n219 10.6151
R1312 B.n331 B.n330 10.6151
R1313 B.n332 B.n331 10.6151
R1314 B.n332 B.n217 10.6151
R1315 B.n336 B.n217 10.6151
R1316 B.n337 B.n336 10.6151
R1317 B.n338 B.n337 10.6151
R1318 B.n338 B.n215 10.6151
R1319 B.n342 B.n215 10.6151
R1320 B.n343 B.n342 10.6151
R1321 B.n344 B.n343 10.6151
R1322 B.n344 B.n213 10.6151
R1323 B.n348 B.n213 10.6151
R1324 B.n349 B.n348 10.6151
R1325 B.n350 B.n349 10.6151
R1326 B.n350 B.n211 10.6151
R1327 B.n354 B.n211 10.6151
R1328 B.n355 B.n354 10.6151
R1329 B.n356 B.n355 10.6151
R1330 B.n356 B.n209 10.6151
R1331 B.n360 B.n209 10.6151
R1332 B.n361 B.n360 10.6151
R1333 B.n362 B.n361 10.6151
R1334 B.n362 B.n207 10.6151
R1335 B.n366 B.n207 10.6151
R1336 B.n367 B.n366 10.6151
R1337 B.n368 B.n367 10.6151
R1338 B.n368 B.n205 10.6151
R1339 B.n372 B.n205 10.6151
R1340 B.n373 B.n372 10.6151
R1341 B.n374 B.n373 10.6151
R1342 B.n374 B.n203 10.6151
R1343 B.n378 B.n203 10.6151
R1344 B.n379 B.n378 10.6151
R1345 B.n380 B.n379 10.6151
R1346 B.n380 B.n201 10.6151
R1347 B.n384 B.n201 10.6151
R1348 B.n385 B.n384 10.6151
R1349 B.n386 B.n385 10.6151
R1350 B.n386 B.n199 10.6151
R1351 B.n390 B.n199 10.6151
R1352 B.n391 B.n390 10.6151
R1353 B.n392 B.n391 10.6151
R1354 B.n392 B.n197 10.6151
R1355 B.n396 B.n197 10.6151
R1356 B.n397 B.n396 10.6151
R1357 B.n398 B.n397 10.6151
R1358 B.n398 B.n195 10.6151
R1359 B.n402 B.n195 10.6151
R1360 B.n403 B.n402 10.6151
R1361 B.n404 B.n403 10.6151
R1362 B.n404 B.n193 10.6151
R1363 B.n408 B.n193 10.6151
R1364 B.n409 B.n408 10.6151
R1365 B.n410 B.n409 10.6151
R1366 B.n410 B.n191 10.6151
R1367 B.n414 B.n191 10.6151
R1368 B.n417 B.n416 10.6151
R1369 B.n417 B.n187 10.6151
R1370 B.n421 B.n187 10.6151
R1371 B.n422 B.n421 10.6151
R1372 B.n423 B.n422 10.6151
R1373 B.n423 B.n185 10.6151
R1374 B.n427 B.n185 10.6151
R1375 B.n428 B.n427 10.6151
R1376 B.n430 B.n181 10.6151
R1377 B.n434 B.n181 10.6151
R1378 B.n435 B.n434 10.6151
R1379 B.n436 B.n435 10.6151
R1380 B.n436 B.n179 10.6151
R1381 B.n440 B.n179 10.6151
R1382 B.n441 B.n440 10.6151
R1383 B.n442 B.n441 10.6151
R1384 B.n442 B.n177 10.6151
R1385 B.n446 B.n177 10.6151
R1386 B.n447 B.n446 10.6151
R1387 B.n448 B.n447 10.6151
R1388 B.n448 B.n175 10.6151
R1389 B.n452 B.n175 10.6151
R1390 B.n453 B.n452 10.6151
R1391 B.n454 B.n453 10.6151
R1392 B.n454 B.n173 10.6151
R1393 B.n458 B.n173 10.6151
R1394 B.n459 B.n458 10.6151
R1395 B.n460 B.n459 10.6151
R1396 B.n460 B.n171 10.6151
R1397 B.n464 B.n171 10.6151
R1398 B.n465 B.n464 10.6151
R1399 B.n466 B.n465 10.6151
R1400 B.n466 B.n169 10.6151
R1401 B.n470 B.n169 10.6151
R1402 B.n471 B.n470 10.6151
R1403 B.n472 B.n471 10.6151
R1404 B.n472 B.n167 10.6151
R1405 B.n476 B.n167 10.6151
R1406 B.n477 B.n476 10.6151
R1407 B.n478 B.n477 10.6151
R1408 B.n478 B.n165 10.6151
R1409 B.n482 B.n165 10.6151
R1410 B.n483 B.n482 10.6151
R1411 B.n484 B.n483 10.6151
R1412 B.n484 B.n163 10.6151
R1413 B.n488 B.n163 10.6151
R1414 B.n489 B.n488 10.6151
R1415 B.n490 B.n489 10.6151
R1416 B.n490 B.n161 10.6151
R1417 B.n494 B.n161 10.6151
R1418 B.n495 B.n494 10.6151
R1419 B.n496 B.n495 10.6151
R1420 B.n496 B.n159 10.6151
R1421 B.n500 B.n159 10.6151
R1422 B.n501 B.n500 10.6151
R1423 B.n502 B.n501 10.6151
R1424 B.n502 B.n157 10.6151
R1425 B.n506 B.n157 10.6151
R1426 B.n507 B.n506 10.6151
R1427 B.n508 B.n507 10.6151
R1428 B.n508 B.n155 10.6151
R1429 B.n512 B.n155 10.6151
R1430 B.n513 B.n512 10.6151
R1431 B.n514 B.n513 10.6151
R1432 B.n514 B.n153 10.6151
R1433 B.n518 B.n153 10.6151
R1434 B.n957 B.n0 8.11757
R1435 B.n957 B.n1 8.11757
R1436 B.n785 B.n62 6.5566
R1437 B.n773 B.n772 6.5566
R1438 B.n416 B.n415 6.5566
R1439 B.n429 B.n428 6.5566
R1440 B.n62 B.n58 4.05904
R1441 B.n772 B.n771 4.05904
R1442 B.n415 B.n414 4.05904
R1443 B.n430 B.n429 4.05904
R1444 VP.n18 VP.t3 183.798
R1445 VP.n19 VP.n16 161.3
R1446 VP.n21 VP.n20 161.3
R1447 VP.n22 VP.n15 161.3
R1448 VP.n24 VP.n23 161.3
R1449 VP.n25 VP.n14 161.3
R1450 VP.n27 VP.n26 161.3
R1451 VP.n29 VP.n13 161.3
R1452 VP.n31 VP.n30 161.3
R1453 VP.n32 VP.n12 161.3
R1454 VP.n34 VP.n33 161.3
R1455 VP.n35 VP.n11 161.3
R1456 VP.n37 VP.n36 161.3
R1457 VP.n69 VP.n68 161.3
R1458 VP.n67 VP.n1 161.3
R1459 VP.n66 VP.n65 161.3
R1460 VP.n64 VP.n2 161.3
R1461 VP.n63 VP.n62 161.3
R1462 VP.n61 VP.n3 161.3
R1463 VP.n59 VP.n58 161.3
R1464 VP.n57 VP.n4 161.3
R1465 VP.n56 VP.n55 161.3
R1466 VP.n54 VP.n5 161.3
R1467 VP.n53 VP.n52 161.3
R1468 VP.n51 VP.n6 161.3
R1469 VP.n50 VP.n49 161.3
R1470 VP.n47 VP.n7 161.3
R1471 VP.n46 VP.n45 161.3
R1472 VP.n44 VP.n8 161.3
R1473 VP.n43 VP.n42 161.3
R1474 VP.n41 VP.n9 161.3
R1475 VP.n40 VP.t7 151.839
R1476 VP.n48 VP.t6 151.839
R1477 VP.n60 VP.t4 151.839
R1478 VP.n0 VP.t2 151.839
R1479 VP.n10 VP.t5 151.839
R1480 VP.n28 VP.t0 151.839
R1481 VP.n17 VP.t1 151.839
R1482 VP.n40 VP.n39 66.0897
R1483 VP.n70 VP.n0 66.0897
R1484 VP.n38 VP.n10 66.0897
R1485 VP.n18 VP.n17 57.5527
R1486 VP.n39 VP.n38 56.5296
R1487 VP.n55 VP.n54 56.5193
R1488 VP.n23 VP.n22 56.5193
R1489 VP.n46 VP.n8 49.2348
R1490 VP.n66 VP.n2 49.2348
R1491 VP.n34 VP.n12 49.2348
R1492 VP.n42 VP.n8 31.752
R1493 VP.n67 VP.n66 31.752
R1494 VP.n35 VP.n34 31.752
R1495 VP.n42 VP.n41 24.4675
R1496 VP.n47 VP.n46 24.4675
R1497 VP.n49 VP.n47 24.4675
R1498 VP.n53 VP.n6 24.4675
R1499 VP.n54 VP.n53 24.4675
R1500 VP.n55 VP.n4 24.4675
R1501 VP.n59 VP.n4 24.4675
R1502 VP.n62 VP.n61 24.4675
R1503 VP.n62 VP.n2 24.4675
R1504 VP.n68 VP.n67 24.4675
R1505 VP.n36 VP.n35 24.4675
R1506 VP.n23 VP.n14 24.4675
R1507 VP.n27 VP.n14 24.4675
R1508 VP.n30 VP.n29 24.4675
R1509 VP.n30 VP.n12 24.4675
R1510 VP.n21 VP.n16 24.4675
R1511 VP.n22 VP.n21 24.4675
R1512 VP.n41 VP.n40 23.9782
R1513 VP.n68 VP.n0 23.9782
R1514 VP.n36 VP.n10 23.9782
R1515 VP.n48 VP.n6 16.1487
R1516 VP.n60 VP.n59 16.1487
R1517 VP.n28 VP.n27 16.1487
R1518 VP.n17 VP.n16 16.1487
R1519 VP.n49 VP.n48 8.31928
R1520 VP.n61 VP.n60 8.31928
R1521 VP.n29 VP.n28 8.31928
R1522 VP.n19 VP.n18 5.24057
R1523 VP.n38 VP.n37 0.354971
R1524 VP.n39 VP.n9 0.354971
R1525 VP.n70 VP.n69 0.354971
R1526 VP VP.n70 0.26696
R1527 VP.n20 VP.n19 0.189894
R1528 VP.n20 VP.n15 0.189894
R1529 VP.n24 VP.n15 0.189894
R1530 VP.n25 VP.n24 0.189894
R1531 VP.n26 VP.n25 0.189894
R1532 VP.n26 VP.n13 0.189894
R1533 VP.n31 VP.n13 0.189894
R1534 VP.n32 VP.n31 0.189894
R1535 VP.n33 VP.n32 0.189894
R1536 VP.n33 VP.n11 0.189894
R1537 VP.n37 VP.n11 0.189894
R1538 VP.n43 VP.n9 0.189894
R1539 VP.n44 VP.n43 0.189894
R1540 VP.n45 VP.n44 0.189894
R1541 VP.n45 VP.n7 0.189894
R1542 VP.n50 VP.n7 0.189894
R1543 VP.n51 VP.n50 0.189894
R1544 VP.n52 VP.n51 0.189894
R1545 VP.n52 VP.n5 0.189894
R1546 VP.n56 VP.n5 0.189894
R1547 VP.n57 VP.n56 0.189894
R1548 VP.n58 VP.n57 0.189894
R1549 VP.n58 VP.n3 0.189894
R1550 VP.n63 VP.n3 0.189894
R1551 VP.n64 VP.n63 0.189894
R1552 VP.n65 VP.n64 0.189894
R1553 VP.n65 VP.n1 0.189894
R1554 VP.n69 VP.n1 0.189894
R1555 VDD1 VDD1.n0 69.3013
R1556 VDD1.n3 VDD1.n2 69.1875
R1557 VDD1.n3 VDD1.n1 69.1875
R1558 VDD1.n5 VDD1.n4 67.8808
R1559 VDD1.n5 VDD1.n3 51.9276
R1560 VDD1.n4 VDD1.t6 1.82355
R1561 VDD1.n4 VDD1.t3 1.82355
R1562 VDD1.n0 VDD1.t1 1.82355
R1563 VDD1.n0 VDD1.t0 1.82355
R1564 VDD1.n2 VDD1.t7 1.82355
R1565 VDD1.n2 VDD1.t4 1.82355
R1566 VDD1.n1 VDD1.t5 1.82355
R1567 VDD1.n1 VDD1.t2 1.82355
R1568 VDD1 VDD1.n5 1.30438
R1569 VTAIL.n11 VTAIL.t12 53.0253
R1570 VTAIL.n10 VTAIL.t7 53.0253
R1571 VTAIL.n7 VTAIL.t0 53.0253
R1572 VTAIL.n15 VTAIL.t3 53.025
R1573 VTAIL.n2 VTAIL.t4 53.025
R1574 VTAIL.n3 VTAIL.t13 53.025
R1575 VTAIL.n6 VTAIL.t8 53.025
R1576 VTAIL.n14 VTAIL.t10 53.025
R1577 VTAIL.n13 VTAIL.n12 51.2022
R1578 VTAIL.n9 VTAIL.n8 51.2022
R1579 VTAIL.n1 VTAIL.n0 51.202
R1580 VTAIL.n5 VTAIL.n4 51.202
R1581 VTAIL.n15 VTAIL.n14 30.4617
R1582 VTAIL.n7 VTAIL.n6 30.4617
R1583 VTAIL.n9 VTAIL.n7 2.72464
R1584 VTAIL.n10 VTAIL.n9 2.72464
R1585 VTAIL.n13 VTAIL.n11 2.72464
R1586 VTAIL.n14 VTAIL.n13 2.72464
R1587 VTAIL.n6 VTAIL.n5 2.72464
R1588 VTAIL.n5 VTAIL.n3 2.72464
R1589 VTAIL.n2 VTAIL.n1 2.72464
R1590 VTAIL VTAIL.n15 2.66645
R1591 VTAIL.n0 VTAIL.t1 1.82355
R1592 VTAIL.n0 VTAIL.t6 1.82355
R1593 VTAIL.n4 VTAIL.t9 1.82355
R1594 VTAIL.n4 VTAIL.t11 1.82355
R1595 VTAIL.n12 VTAIL.t14 1.82355
R1596 VTAIL.n12 VTAIL.t15 1.82355
R1597 VTAIL.n8 VTAIL.t5 1.82355
R1598 VTAIL.n8 VTAIL.t2 1.82355
R1599 VTAIL.n11 VTAIL.n10 0.470328
R1600 VTAIL.n3 VTAIL.n2 0.470328
R1601 VTAIL VTAIL.n1 0.0586897
R1602 VN.n37 VN.t2 183.798
R1603 VN.n8 VN.t4 183.798
R1604 VN.n56 VN.n55 161.3
R1605 VN.n54 VN.n30 161.3
R1606 VN.n53 VN.n52 161.3
R1607 VN.n51 VN.n31 161.3
R1608 VN.n50 VN.n49 161.3
R1609 VN.n48 VN.n32 161.3
R1610 VN.n46 VN.n45 161.3
R1611 VN.n44 VN.n33 161.3
R1612 VN.n43 VN.n42 161.3
R1613 VN.n41 VN.n34 161.3
R1614 VN.n40 VN.n39 161.3
R1615 VN.n38 VN.n35 161.3
R1616 VN.n27 VN.n26 161.3
R1617 VN.n25 VN.n1 161.3
R1618 VN.n24 VN.n23 161.3
R1619 VN.n22 VN.n2 161.3
R1620 VN.n21 VN.n20 161.3
R1621 VN.n19 VN.n3 161.3
R1622 VN.n17 VN.n16 161.3
R1623 VN.n15 VN.n4 161.3
R1624 VN.n14 VN.n13 161.3
R1625 VN.n12 VN.n5 161.3
R1626 VN.n11 VN.n10 161.3
R1627 VN.n9 VN.n6 161.3
R1628 VN.n7 VN.t5 151.839
R1629 VN.n18 VN.t3 151.839
R1630 VN.n0 VN.t6 151.839
R1631 VN.n36 VN.t0 151.839
R1632 VN.n47 VN.t1 151.839
R1633 VN.n29 VN.t7 151.839
R1634 VN.n28 VN.n0 66.0897
R1635 VN.n57 VN.n29 66.0897
R1636 VN.n8 VN.n7 57.5527
R1637 VN.n37 VN.n36 57.5527
R1638 VN VN.n57 56.695
R1639 VN.n13 VN.n12 56.5193
R1640 VN.n42 VN.n41 56.5193
R1641 VN.n24 VN.n2 49.2348
R1642 VN.n53 VN.n31 49.2348
R1643 VN.n25 VN.n24 31.752
R1644 VN.n54 VN.n53 31.752
R1645 VN.n11 VN.n6 24.4675
R1646 VN.n12 VN.n11 24.4675
R1647 VN.n13 VN.n4 24.4675
R1648 VN.n17 VN.n4 24.4675
R1649 VN.n20 VN.n19 24.4675
R1650 VN.n20 VN.n2 24.4675
R1651 VN.n26 VN.n25 24.4675
R1652 VN.n41 VN.n40 24.4675
R1653 VN.n40 VN.n35 24.4675
R1654 VN.n49 VN.n31 24.4675
R1655 VN.n49 VN.n48 24.4675
R1656 VN.n46 VN.n33 24.4675
R1657 VN.n42 VN.n33 24.4675
R1658 VN.n55 VN.n54 24.4675
R1659 VN.n26 VN.n0 23.9782
R1660 VN.n55 VN.n29 23.9782
R1661 VN.n7 VN.n6 16.1487
R1662 VN.n18 VN.n17 16.1487
R1663 VN.n36 VN.n35 16.1487
R1664 VN.n47 VN.n46 16.1487
R1665 VN.n19 VN.n18 8.31928
R1666 VN.n48 VN.n47 8.31928
R1667 VN.n38 VN.n37 5.2406
R1668 VN.n9 VN.n8 5.2406
R1669 VN.n57 VN.n56 0.354971
R1670 VN.n28 VN.n27 0.354971
R1671 VN VN.n28 0.26696
R1672 VN.n56 VN.n30 0.189894
R1673 VN.n52 VN.n30 0.189894
R1674 VN.n52 VN.n51 0.189894
R1675 VN.n51 VN.n50 0.189894
R1676 VN.n50 VN.n32 0.189894
R1677 VN.n45 VN.n32 0.189894
R1678 VN.n45 VN.n44 0.189894
R1679 VN.n44 VN.n43 0.189894
R1680 VN.n43 VN.n34 0.189894
R1681 VN.n39 VN.n34 0.189894
R1682 VN.n39 VN.n38 0.189894
R1683 VN.n10 VN.n9 0.189894
R1684 VN.n10 VN.n5 0.189894
R1685 VN.n14 VN.n5 0.189894
R1686 VN.n15 VN.n14 0.189894
R1687 VN.n16 VN.n15 0.189894
R1688 VN.n16 VN.n3 0.189894
R1689 VN.n21 VN.n3 0.189894
R1690 VN.n22 VN.n21 0.189894
R1691 VN.n23 VN.n22 0.189894
R1692 VN.n23 VN.n1 0.189894
R1693 VN.n27 VN.n1 0.189894
R1694 VDD2.n2 VDD2.n1 69.1875
R1695 VDD2.n2 VDD2.n0 69.1875
R1696 VDD2 VDD2.n5 69.1847
R1697 VDD2.n4 VDD2.n3 67.881
R1698 VDD2.n4 VDD2.n2 51.3446
R1699 VDD2.n5 VDD2.t7 1.82355
R1700 VDD2.n5 VDD2.t5 1.82355
R1701 VDD2.n3 VDD2.t0 1.82355
R1702 VDD2.n3 VDD2.t6 1.82355
R1703 VDD2.n1 VDD2.t4 1.82355
R1704 VDD2.n1 VDD2.t1 1.82355
R1705 VDD2.n0 VDD2.t3 1.82355
R1706 VDD2.n0 VDD2.t2 1.82355
R1707 VDD2 VDD2.n4 1.42076
C0 VP w_n4130_n4534# 9.11933f
C1 VDD2 VN 12.9085f
C2 VP B 2.24835f
C3 VN w_n4130_n4534# 8.58249f
C4 VDD2 VDD1 1.89599f
C5 w_n4130_n4534# VDD1 2.18336f
C6 VN B 1.3472f
C7 B VDD1 1.87579f
C8 VDD2 VTAIL 10.0639f
C9 VTAIL w_n4130_n4534# 5.53261f
C10 VN VP 9.025769f
C11 VP VDD1 13.299f
C12 VTAIL B 7.02408f
C13 VN VDD1 0.151975f
C14 VTAIL VP 13.1285f
C15 VTAIL VN 13.1144f
C16 VTAIL VDD1 10.008f
C17 VDD2 w_n4130_n4534# 2.30771f
C18 VDD2 B 1.97906f
C19 B w_n4130_n4534# 12.1025f
C20 VDD2 VP 0.543976f
C21 VDD2 VSUBS 2.10543f
C22 VDD1 VSUBS 2.78966f
C23 VTAIL VSUBS 1.637922f
C24 VN VSUBS 7.279759f
C25 VP VSUBS 4.047893f
C26 B VSUBS 5.754088f
C27 w_n4130_n4534# VSUBS 0.229017p
C28 VDD2.t3 VSUBS 0.376207f
C29 VDD2.t2 VSUBS 0.376207f
C30 VDD2.n0 VSUBS 3.13284f
C31 VDD2.t4 VSUBS 0.376207f
C32 VDD2.t1 VSUBS 0.376207f
C33 VDD2.n1 VSUBS 3.13284f
C34 VDD2.n2 VSUBS 4.651f
C35 VDD2.t0 VSUBS 0.376207f
C36 VDD2.t6 VSUBS 0.376207f
C37 VDD2.n3 VSUBS 3.11604f
C38 VDD2.n4 VSUBS 4.01834f
C39 VDD2.t7 VSUBS 0.376207f
C40 VDD2.t5 VSUBS 0.376207f
C41 VDD2.n5 VSUBS 3.13278f
C42 VN.t6 VSUBS 3.45487f
C43 VN.n0 VSUBS 1.29682f
C44 VN.n1 VSUBS 0.024897f
C45 VN.n2 VSUBS 0.046169f
C46 VN.n3 VSUBS 0.024897f
C47 VN.t3 VSUBS 3.45487f
C48 VN.n4 VSUBS 0.046402f
C49 VN.n5 VSUBS 0.024897f
C50 VN.n6 VSUBS 0.038613f
C51 VN.t5 VSUBS 3.45487f
C52 VN.n7 VSUBS 1.27701f
C53 VN.t4 VSUBS 3.6917f
C54 VN.n8 VSUBS 1.24412f
C55 VN.n9 VSUBS 0.262386f
C56 VN.n10 VSUBS 0.024897f
C57 VN.n11 VSUBS 0.046402f
C58 VN.n12 VSUBS 0.036345f
C59 VN.n13 VSUBS 0.036345f
C60 VN.n14 VSUBS 0.024897f
C61 VN.n15 VSUBS 0.024897f
C62 VN.n16 VSUBS 0.024897f
C63 VN.n17 VSUBS 0.038613f
C64 VN.n18 VSUBS 1.19647f
C65 VN.n19 VSUBS 0.031282f
C66 VN.n20 VSUBS 0.046402f
C67 VN.n21 VSUBS 0.024897f
C68 VN.n22 VSUBS 0.024897f
C69 VN.n23 VSUBS 0.024897f
C70 VN.n24 VSUBS 0.022844f
C71 VN.n25 VSUBS 0.050079f
C72 VN.n26 VSUBS 0.045944f
C73 VN.n27 VSUBS 0.040183f
C74 VN.n28 VSUBS 0.045819f
C75 VN.t7 VSUBS 3.45487f
C76 VN.n29 VSUBS 1.29682f
C77 VN.n30 VSUBS 0.024897f
C78 VN.n31 VSUBS 0.046169f
C79 VN.n32 VSUBS 0.024897f
C80 VN.t1 VSUBS 3.45487f
C81 VN.n33 VSUBS 0.046402f
C82 VN.n34 VSUBS 0.024897f
C83 VN.n35 VSUBS 0.038613f
C84 VN.t2 VSUBS 3.6917f
C85 VN.t0 VSUBS 3.45487f
C86 VN.n36 VSUBS 1.27701f
C87 VN.n37 VSUBS 1.24412f
C88 VN.n38 VSUBS 0.262386f
C89 VN.n39 VSUBS 0.024897f
C90 VN.n40 VSUBS 0.046402f
C91 VN.n41 VSUBS 0.036345f
C92 VN.n42 VSUBS 0.036345f
C93 VN.n43 VSUBS 0.024897f
C94 VN.n44 VSUBS 0.024897f
C95 VN.n45 VSUBS 0.024897f
C96 VN.n46 VSUBS 0.038613f
C97 VN.n47 VSUBS 1.19647f
C98 VN.n48 VSUBS 0.031282f
C99 VN.n49 VSUBS 0.046402f
C100 VN.n50 VSUBS 0.024897f
C101 VN.n51 VSUBS 0.024897f
C102 VN.n52 VSUBS 0.024897f
C103 VN.n53 VSUBS 0.022844f
C104 VN.n54 VSUBS 0.050079f
C105 VN.n55 VSUBS 0.045944f
C106 VN.n56 VSUBS 0.040183f
C107 VN.n57 VSUBS 1.67666f
C108 VTAIL.t1 VSUBS 0.33444f
C109 VTAIL.t6 VSUBS 0.33444f
C110 VTAIL.n0 VSUBS 2.61764f
C111 VTAIL.n1 VSUBS 0.805556f
C112 VTAIL.t4 VSUBS 3.41989f
C113 VTAIL.n2 VSUBS 0.946898f
C114 VTAIL.t13 VSUBS 3.41989f
C115 VTAIL.n3 VSUBS 0.946898f
C116 VTAIL.t9 VSUBS 0.33444f
C117 VTAIL.t11 VSUBS 0.33444f
C118 VTAIL.n4 VSUBS 2.61764f
C119 VTAIL.n5 VSUBS 1.00946f
C120 VTAIL.t8 VSUBS 3.41989f
C121 VTAIL.n6 VSUBS 2.61736f
C122 VTAIL.t0 VSUBS 3.41989f
C123 VTAIL.n7 VSUBS 2.61735f
C124 VTAIL.t5 VSUBS 0.33444f
C125 VTAIL.t2 VSUBS 0.33444f
C126 VTAIL.n8 VSUBS 2.61764f
C127 VTAIL.n9 VSUBS 1.00945f
C128 VTAIL.t7 VSUBS 3.41989f
C129 VTAIL.n10 VSUBS 0.946892f
C130 VTAIL.t12 VSUBS 3.41989f
C131 VTAIL.n11 VSUBS 0.946892f
C132 VTAIL.t14 VSUBS 0.33444f
C133 VTAIL.t15 VSUBS 0.33444f
C134 VTAIL.n12 VSUBS 2.61764f
C135 VTAIL.n13 VSUBS 1.00945f
C136 VTAIL.t10 VSUBS 3.41989f
C137 VTAIL.n14 VSUBS 2.61736f
C138 VTAIL.t3 VSUBS 3.41989f
C139 VTAIL.n15 VSUBS 2.6129f
C140 VDD1.t1 VSUBS 0.377709f
C141 VDD1.t0 VSUBS 0.377709f
C142 VDD1.n0 VSUBS 3.14698f
C143 VDD1.t5 VSUBS 0.377709f
C144 VDD1.t2 VSUBS 0.377709f
C145 VDD1.n1 VSUBS 3.14535f
C146 VDD1.t7 VSUBS 0.377709f
C147 VDD1.t4 VSUBS 0.377709f
C148 VDD1.n2 VSUBS 3.14535f
C149 VDD1.n3 VSUBS 4.72501f
C150 VDD1.t6 VSUBS 0.377709f
C151 VDD1.t3 VSUBS 0.377709f
C152 VDD1.n4 VSUBS 3.12847f
C153 VDD1.n5 VSUBS 4.06791f
C154 VP.t2 VSUBS 3.70348f
C155 VP.n0 VSUBS 1.39014f
C156 VP.n1 VSUBS 0.026689f
C157 VP.n2 VSUBS 0.049492f
C158 VP.n3 VSUBS 0.026689f
C159 VP.t4 VSUBS 3.70348f
C160 VP.n4 VSUBS 0.049741f
C161 VP.n5 VSUBS 0.026689f
C162 VP.n6 VSUBS 0.041392f
C163 VP.n7 VSUBS 0.026689f
C164 VP.n8 VSUBS 0.024487f
C165 VP.n9 VSUBS 0.043075f
C166 VP.t7 VSUBS 3.70348f
C167 VP.t5 VSUBS 3.70348f
C168 VP.n10 VSUBS 1.39014f
C169 VP.n11 VSUBS 0.026689f
C170 VP.n12 VSUBS 0.049492f
C171 VP.n13 VSUBS 0.026689f
C172 VP.t0 VSUBS 3.70348f
C173 VP.n14 VSUBS 0.049741f
C174 VP.n15 VSUBS 0.026689f
C175 VP.n16 VSUBS 0.041392f
C176 VP.t3 VSUBS 3.95736f
C177 VP.t1 VSUBS 3.70348f
C178 VP.n17 VSUBS 1.36891f
C179 VP.n18 VSUBS 1.33365f
C180 VP.n19 VSUBS 0.281268f
C181 VP.n20 VSUBS 0.026689f
C182 VP.n21 VSUBS 0.049741f
C183 VP.n22 VSUBS 0.038961f
C184 VP.n23 VSUBS 0.038961f
C185 VP.n24 VSUBS 0.026689f
C186 VP.n25 VSUBS 0.026689f
C187 VP.n26 VSUBS 0.026689f
C188 VP.n27 VSUBS 0.041392f
C189 VP.n28 VSUBS 1.28257f
C190 VP.n29 VSUBS 0.033533f
C191 VP.n30 VSUBS 0.049741f
C192 VP.n31 VSUBS 0.026689f
C193 VP.n32 VSUBS 0.026689f
C194 VP.n33 VSUBS 0.026689f
C195 VP.n34 VSUBS 0.024487f
C196 VP.n35 VSUBS 0.053683f
C197 VP.n36 VSUBS 0.04925f
C198 VP.n37 VSUBS 0.043075f
C199 VP.n38 VSUBS 1.78683f
C200 VP.n39 VSUBS 1.8038f
C201 VP.n40 VSUBS 1.39014f
C202 VP.n41 VSUBS 0.04925f
C203 VP.n42 VSUBS 0.053683f
C204 VP.n43 VSUBS 0.026689f
C205 VP.n44 VSUBS 0.026689f
C206 VP.n45 VSUBS 0.026689f
C207 VP.n46 VSUBS 0.049492f
C208 VP.n47 VSUBS 0.049741f
C209 VP.t6 VSUBS 3.70348f
C210 VP.n48 VSUBS 1.28257f
C211 VP.n49 VSUBS 0.033533f
C212 VP.n50 VSUBS 0.026689f
C213 VP.n51 VSUBS 0.026689f
C214 VP.n52 VSUBS 0.026689f
C215 VP.n53 VSUBS 0.049741f
C216 VP.n54 VSUBS 0.038961f
C217 VP.n55 VSUBS 0.038961f
C218 VP.n56 VSUBS 0.026689f
C219 VP.n57 VSUBS 0.026689f
C220 VP.n58 VSUBS 0.026689f
C221 VP.n59 VSUBS 0.041392f
C222 VP.n60 VSUBS 1.28257f
C223 VP.n61 VSUBS 0.033533f
C224 VP.n62 VSUBS 0.049741f
C225 VP.n63 VSUBS 0.026689f
C226 VP.n64 VSUBS 0.026689f
C227 VP.n65 VSUBS 0.026689f
C228 VP.n66 VSUBS 0.024487f
C229 VP.n67 VSUBS 0.053683f
C230 VP.n68 VSUBS 0.04925f
C231 VP.n69 VSUBS 0.043075f
C232 VP.n70 VSUBS 0.049117f
C233 B.n0 VSUBS 0.005854f
C234 B.n1 VSUBS 0.005854f
C235 B.n2 VSUBS 0.008657f
C236 B.n3 VSUBS 0.006634f
C237 B.n4 VSUBS 0.006634f
C238 B.n5 VSUBS 0.006634f
C239 B.n6 VSUBS 0.006634f
C240 B.n7 VSUBS 0.006634f
C241 B.n8 VSUBS 0.006634f
C242 B.n9 VSUBS 0.006634f
C243 B.n10 VSUBS 0.006634f
C244 B.n11 VSUBS 0.006634f
C245 B.n12 VSUBS 0.006634f
C246 B.n13 VSUBS 0.006634f
C247 B.n14 VSUBS 0.006634f
C248 B.n15 VSUBS 0.006634f
C249 B.n16 VSUBS 0.006634f
C250 B.n17 VSUBS 0.006634f
C251 B.n18 VSUBS 0.006634f
C252 B.n19 VSUBS 0.006634f
C253 B.n20 VSUBS 0.006634f
C254 B.n21 VSUBS 0.006634f
C255 B.n22 VSUBS 0.006634f
C256 B.n23 VSUBS 0.006634f
C257 B.n24 VSUBS 0.006634f
C258 B.n25 VSUBS 0.006634f
C259 B.n26 VSUBS 0.006634f
C260 B.n27 VSUBS 0.006634f
C261 B.n28 VSUBS 0.006634f
C262 B.n29 VSUBS 0.01628f
C263 B.n30 VSUBS 0.006634f
C264 B.n31 VSUBS 0.006634f
C265 B.n32 VSUBS 0.006634f
C266 B.n33 VSUBS 0.006634f
C267 B.n34 VSUBS 0.006634f
C268 B.n35 VSUBS 0.006634f
C269 B.n36 VSUBS 0.006634f
C270 B.n37 VSUBS 0.006634f
C271 B.n38 VSUBS 0.006634f
C272 B.n39 VSUBS 0.006634f
C273 B.n40 VSUBS 0.006634f
C274 B.n41 VSUBS 0.006634f
C275 B.n42 VSUBS 0.006634f
C276 B.n43 VSUBS 0.006634f
C277 B.n44 VSUBS 0.006634f
C278 B.n45 VSUBS 0.006634f
C279 B.n46 VSUBS 0.006634f
C280 B.n47 VSUBS 0.006634f
C281 B.n48 VSUBS 0.006634f
C282 B.n49 VSUBS 0.006634f
C283 B.n50 VSUBS 0.006634f
C284 B.n51 VSUBS 0.006634f
C285 B.n52 VSUBS 0.006634f
C286 B.n53 VSUBS 0.006634f
C287 B.n54 VSUBS 0.006634f
C288 B.n55 VSUBS 0.006634f
C289 B.n56 VSUBS 0.006634f
C290 B.n57 VSUBS 0.006634f
C291 B.n58 VSUBS 0.004585f
C292 B.n59 VSUBS 0.006634f
C293 B.t7 VSUBS 0.570101f
C294 B.t8 VSUBS 0.591601f
C295 B.t6 VSUBS 2.13595f
C296 B.n60 VSUBS 0.33371f
C297 B.n61 VSUBS 0.069239f
C298 B.n62 VSUBS 0.015371f
C299 B.n63 VSUBS 0.006634f
C300 B.n64 VSUBS 0.006634f
C301 B.n65 VSUBS 0.006634f
C302 B.n66 VSUBS 0.006634f
C303 B.t10 VSUBS 0.57008f
C304 B.t11 VSUBS 0.591585f
C305 B.t9 VSUBS 2.13595f
C306 B.n67 VSUBS 0.333727f
C307 B.n68 VSUBS 0.06926f
C308 B.n69 VSUBS 0.006634f
C309 B.n70 VSUBS 0.006634f
C310 B.n71 VSUBS 0.006634f
C311 B.n72 VSUBS 0.006634f
C312 B.n73 VSUBS 0.006634f
C313 B.n74 VSUBS 0.006634f
C314 B.n75 VSUBS 0.006634f
C315 B.n76 VSUBS 0.006634f
C316 B.n77 VSUBS 0.006634f
C317 B.n78 VSUBS 0.006634f
C318 B.n79 VSUBS 0.006634f
C319 B.n80 VSUBS 0.006634f
C320 B.n81 VSUBS 0.006634f
C321 B.n82 VSUBS 0.006634f
C322 B.n83 VSUBS 0.006634f
C323 B.n84 VSUBS 0.006634f
C324 B.n85 VSUBS 0.006634f
C325 B.n86 VSUBS 0.006634f
C326 B.n87 VSUBS 0.006634f
C327 B.n88 VSUBS 0.006634f
C328 B.n89 VSUBS 0.006634f
C329 B.n90 VSUBS 0.006634f
C330 B.n91 VSUBS 0.006634f
C331 B.n92 VSUBS 0.006634f
C332 B.n93 VSUBS 0.006634f
C333 B.n94 VSUBS 0.006634f
C334 B.n95 VSUBS 0.006634f
C335 B.n96 VSUBS 0.006634f
C336 B.n97 VSUBS 0.01628f
C337 B.n98 VSUBS 0.006634f
C338 B.n99 VSUBS 0.006634f
C339 B.n100 VSUBS 0.006634f
C340 B.n101 VSUBS 0.006634f
C341 B.n102 VSUBS 0.006634f
C342 B.n103 VSUBS 0.006634f
C343 B.n104 VSUBS 0.006634f
C344 B.n105 VSUBS 0.006634f
C345 B.n106 VSUBS 0.006634f
C346 B.n107 VSUBS 0.006634f
C347 B.n108 VSUBS 0.006634f
C348 B.n109 VSUBS 0.006634f
C349 B.n110 VSUBS 0.006634f
C350 B.n111 VSUBS 0.006634f
C351 B.n112 VSUBS 0.006634f
C352 B.n113 VSUBS 0.006634f
C353 B.n114 VSUBS 0.006634f
C354 B.n115 VSUBS 0.006634f
C355 B.n116 VSUBS 0.006634f
C356 B.n117 VSUBS 0.006634f
C357 B.n118 VSUBS 0.006634f
C358 B.n119 VSUBS 0.006634f
C359 B.n120 VSUBS 0.006634f
C360 B.n121 VSUBS 0.006634f
C361 B.n122 VSUBS 0.006634f
C362 B.n123 VSUBS 0.006634f
C363 B.n124 VSUBS 0.006634f
C364 B.n125 VSUBS 0.006634f
C365 B.n126 VSUBS 0.006634f
C366 B.n127 VSUBS 0.006634f
C367 B.n128 VSUBS 0.006634f
C368 B.n129 VSUBS 0.006634f
C369 B.n130 VSUBS 0.006634f
C370 B.n131 VSUBS 0.006634f
C371 B.n132 VSUBS 0.006634f
C372 B.n133 VSUBS 0.006634f
C373 B.n134 VSUBS 0.006634f
C374 B.n135 VSUBS 0.006634f
C375 B.n136 VSUBS 0.006634f
C376 B.n137 VSUBS 0.006634f
C377 B.n138 VSUBS 0.006634f
C378 B.n139 VSUBS 0.006634f
C379 B.n140 VSUBS 0.006634f
C380 B.n141 VSUBS 0.006634f
C381 B.n142 VSUBS 0.006634f
C382 B.n143 VSUBS 0.006634f
C383 B.n144 VSUBS 0.006634f
C384 B.n145 VSUBS 0.006634f
C385 B.n146 VSUBS 0.006634f
C386 B.n147 VSUBS 0.006634f
C387 B.n148 VSUBS 0.006634f
C388 B.n149 VSUBS 0.006634f
C389 B.n150 VSUBS 0.006634f
C390 B.n151 VSUBS 0.006634f
C391 B.n152 VSUBS 0.015525f
C392 B.n153 VSUBS 0.006634f
C393 B.n154 VSUBS 0.006634f
C394 B.n155 VSUBS 0.006634f
C395 B.n156 VSUBS 0.006634f
C396 B.n157 VSUBS 0.006634f
C397 B.n158 VSUBS 0.006634f
C398 B.n159 VSUBS 0.006634f
C399 B.n160 VSUBS 0.006634f
C400 B.n161 VSUBS 0.006634f
C401 B.n162 VSUBS 0.006634f
C402 B.n163 VSUBS 0.006634f
C403 B.n164 VSUBS 0.006634f
C404 B.n165 VSUBS 0.006634f
C405 B.n166 VSUBS 0.006634f
C406 B.n167 VSUBS 0.006634f
C407 B.n168 VSUBS 0.006634f
C408 B.n169 VSUBS 0.006634f
C409 B.n170 VSUBS 0.006634f
C410 B.n171 VSUBS 0.006634f
C411 B.n172 VSUBS 0.006634f
C412 B.n173 VSUBS 0.006634f
C413 B.n174 VSUBS 0.006634f
C414 B.n175 VSUBS 0.006634f
C415 B.n176 VSUBS 0.006634f
C416 B.n177 VSUBS 0.006634f
C417 B.n178 VSUBS 0.006634f
C418 B.n179 VSUBS 0.006634f
C419 B.n180 VSUBS 0.006634f
C420 B.n181 VSUBS 0.006634f
C421 B.n182 VSUBS 0.006634f
C422 B.t5 VSUBS 0.57008f
C423 B.t4 VSUBS 0.591585f
C424 B.t3 VSUBS 2.13595f
C425 B.n183 VSUBS 0.333727f
C426 B.n184 VSUBS 0.06926f
C427 B.n185 VSUBS 0.006634f
C428 B.n186 VSUBS 0.006634f
C429 B.n187 VSUBS 0.006634f
C430 B.n188 VSUBS 0.006634f
C431 B.t2 VSUBS 0.570101f
C432 B.t1 VSUBS 0.591601f
C433 B.t0 VSUBS 2.13595f
C434 B.n189 VSUBS 0.33371f
C435 B.n190 VSUBS 0.069239f
C436 B.n191 VSUBS 0.006634f
C437 B.n192 VSUBS 0.006634f
C438 B.n193 VSUBS 0.006634f
C439 B.n194 VSUBS 0.006634f
C440 B.n195 VSUBS 0.006634f
C441 B.n196 VSUBS 0.006634f
C442 B.n197 VSUBS 0.006634f
C443 B.n198 VSUBS 0.006634f
C444 B.n199 VSUBS 0.006634f
C445 B.n200 VSUBS 0.006634f
C446 B.n201 VSUBS 0.006634f
C447 B.n202 VSUBS 0.006634f
C448 B.n203 VSUBS 0.006634f
C449 B.n204 VSUBS 0.006634f
C450 B.n205 VSUBS 0.006634f
C451 B.n206 VSUBS 0.006634f
C452 B.n207 VSUBS 0.006634f
C453 B.n208 VSUBS 0.006634f
C454 B.n209 VSUBS 0.006634f
C455 B.n210 VSUBS 0.006634f
C456 B.n211 VSUBS 0.006634f
C457 B.n212 VSUBS 0.006634f
C458 B.n213 VSUBS 0.006634f
C459 B.n214 VSUBS 0.006634f
C460 B.n215 VSUBS 0.006634f
C461 B.n216 VSUBS 0.006634f
C462 B.n217 VSUBS 0.006634f
C463 B.n218 VSUBS 0.006634f
C464 B.n219 VSUBS 0.006634f
C465 B.n220 VSUBS 0.015525f
C466 B.n221 VSUBS 0.006634f
C467 B.n222 VSUBS 0.006634f
C468 B.n223 VSUBS 0.006634f
C469 B.n224 VSUBS 0.006634f
C470 B.n225 VSUBS 0.006634f
C471 B.n226 VSUBS 0.006634f
C472 B.n227 VSUBS 0.006634f
C473 B.n228 VSUBS 0.006634f
C474 B.n229 VSUBS 0.006634f
C475 B.n230 VSUBS 0.006634f
C476 B.n231 VSUBS 0.006634f
C477 B.n232 VSUBS 0.006634f
C478 B.n233 VSUBS 0.006634f
C479 B.n234 VSUBS 0.006634f
C480 B.n235 VSUBS 0.006634f
C481 B.n236 VSUBS 0.006634f
C482 B.n237 VSUBS 0.006634f
C483 B.n238 VSUBS 0.006634f
C484 B.n239 VSUBS 0.006634f
C485 B.n240 VSUBS 0.006634f
C486 B.n241 VSUBS 0.006634f
C487 B.n242 VSUBS 0.006634f
C488 B.n243 VSUBS 0.006634f
C489 B.n244 VSUBS 0.006634f
C490 B.n245 VSUBS 0.006634f
C491 B.n246 VSUBS 0.006634f
C492 B.n247 VSUBS 0.006634f
C493 B.n248 VSUBS 0.006634f
C494 B.n249 VSUBS 0.006634f
C495 B.n250 VSUBS 0.006634f
C496 B.n251 VSUBS 0.006634f
C497 B.n252 VSUBS 0.006634f
C498 B.n253 VSUBS 0.006634f
C499 B.n254 VSUBS 0.006634f
C500 B.n255 VSUBS 0.006634f
C501 B.n256 VSUBS 0.006634f
C502 B.n257 VSUBS 0.006634f
C503 B.n258 VSUBS 0.006634f
C504 B.n259 VSUBS 0.006634f
C505 B.n260 VSUBS 0.006634f
C506 B.n261 VSUBS 0.006634f
C507 B.n262 VSUBS 0.006634f
C508 B.n263 VSUBS 0.006634f
C509 B.n264 VSUBS 0.006634f
C510 B.n265 VSUBS 0.006634f
C511 B.n266 VSUBS 0.006634f
C512 B.n267 VSUBS 0.006634f
C513 B.n268 VSUBS 0.006634f
C514 B.n269 VSUBS 0.006634f
C515 B.n270 VSUBS 0.006634f
C516 B.n271 VSUBS 0.006634f
C517 B.n272 VSUBS 0.006634f
C518 B.n273 VSUBS 0.006634f
C519 B.n274 VSUBS 0.006634f
C520 B.n275 VSUBS 0.006634f
C521 B.n276 VSUBS 0.006634f
C522 B.n277 VSUBS 0.006634f
C523 B.n278 VSUBS 0.006634f
C524 B.n279 VSUBS 0.006634f
C525 B.n280 VSUBS 0.006634f
C526 B.n281 VSUBS 0.006634f
C527 B.n282 VSUBS 0.006634f
C528 B.n283 VSUBS 0.006634f
C529 B.n284 VSUBS 0.006634f
C530 B.n285 VSUBS 0.006634f
C531 B.n286 VSUBS 0.006634f
C532 B.n287 VSUBS 0.006634f
C533 B.n288 VSUBS 0.006634f
C534 B.n289 VSUBS 0.006634f
C535 B.n290 VSUBS 0.006634f
C536 B.n291 VSUBS 0.006634f
C537 B.n292 VSUBS 0.006634f
C538 B.n293 VSUBS 0.006634f
C539 B.n294 VSUBS 0.006634f
C540 B.n295 VSUBS 0.006634f
C541 B.n296 VSUBS 0.006634f
C542 B.n297 VSUBS 0.006634f
C543 B.n298 VSUBS 0.006634f
C544 B.n299 VSUBS 0.006634f
C545 B.n300 VSUBS 0.006634f
C546 B.n301 VSUBS 0.006634f
C547 B.n302 VSUBS 0.006634f
C548 B.n303 VSUBS 0.006634f
C549 B.n304 VSUBS 0.006634f
C550 B.n305 VSUBS 0.006634f
C551 B.n306 VSUBS 0.006634f
C552 B.n307 VSUBS 0.006634f
C553 B.n308 VSUBS 0.006634f
C554 B.n309 VSUBS 0.006634f
C555 B.n310 VSUBS 0.006634f
C556 B.n311 VSUBS 0.006634f
C557 B.n312 VSUBS 0.006634f
C558 B.n313 VSUBS 0.006634f
C559 B.n314 VSUBS 0.006634f
C560 B.n315 VSUBS 0.006634f
C561 B.n316 VSUBS 0.006634f
C562 B.n317 VSUBS 0.006634f
C563 B.n318 VSUBS 0.006634f
C564 B.n319 VSUBS 0.006634f
C565 B.n320 VSUBS 0.006634f
C566 B.n321 VSUBS 0.006634f
C567 B.n322 VSUBS 0.006634f
C568 B.n323 VSUBS 0.006634f
C569 B.n324 VSUBS 0.006634f
C570 B.n325 VSUBS 0.015525f
C571 B.n326 VSUBS 0.01628f
C572 B.n327 VSUBS 0.01628f
C573 B.n328 VSUBS 0.006634f
C574 B.n329 VSUBS 0.006634f
C575 B.n330 VSUBS 0.006634f
C576 B.n331 VSUBS 0.006634f
C577 B.n332 VSUBS 0.006634f
C578 B.n333 VSUBS 0.006634f
C579 B.n334 VSUBS 0.006634f
C580 B.n335 VSUBS 0.006634f
C581 B.n336 VSUBS 0.006634f
C582 B.n337 VSUBS 0.006634f
C583 B.n338 VSUBS 0.006634f
C584 B.n339 VSUBS 0.006634f
C585 B.n340 VSUBS 0.006634f
C586 B.n341 VSUBS 0.006634f
C587 B.n342 VSUBS 0.006634f
C588 B.n343 VSUBS 0.006634f
C589 B.n344 VSUBS 0.006634f
C590 B.n345 VSUBS 0.006634f
C591 B.n346 VSUBS 0.006634f
C592 B.n347 VSUBS 0.006634f
C593 B.n348 VSUBS 0.006634f
C594 B.n349 VSUBS 0.006634f
C595 B.n350 VSUBS 0.006634f
C596 B.n351 VSUBS 0.006634f
C597 B.n352 VSUBS 0.006634f
C598 B.n353 VSUBS 0.006634f
C599 B.n354 VSUBS 0.006634f
C600 B.n355 VSUBS 0.006634f
C601 B.n356 VSUBS 0.006634f
C602 B.n357 VSUBS 0.006634f
C603 B.n358 VSUBS 0.006634f
C604 B.n359 VSUBS 0.006634f
C605 B.n360 VSUBS 0.006634f
C606 B.n361 VSUBS 0.006634f
C607 B.n362 VSUBS 0.006634f
C608 B.n363 VSUBS 0.006634f
C609 B.n364 VSUBS 0.006634f
C610 B.n365 VSUBS 0.006634f
C611 B.n366 VSUBS 0.006634f
C612 B.n367 VSUBS 0.006634f
C613 B.n368 VSUBS 0.006634f
C614 B.n369 VSUBS 0.006634f
C615 B.n370 VSUBS 0.006634f
C616 B.n371 VSUBS 0.006634f
C617 B.n372 VSUBS 0.006634f
C618 B.n373 VSUBS 0.006634f
C619 B.n374 VSUBS 0.006634f
C620 B.n375 VSUBS 0.006634f
C621 B.n376 VSUBS 0.006634f
C622 B.n377 VSUBS 0.006634f
C623 B.n378 VSUBS 0.006634f
C624 B.n379 VSUBS 0.006634f
C625 B.n380 VSUBS 0.006634f
C626 B.n381 VSUBS 0.006634f
C627 B.n382 VSUBS 0.006634f
C628 B.n383 VSUBS 0.006634f
C629 B.n384 VSUBS 0.006634f
C630 B.n385 VSUBS 0.006634f
C631 B.n386 VSUBS 0.006634f
C632 B.n387 VSUBS 0.006634f
C633 B.n388 VSUBS 0.006634f
C634 B.n389 VSUBS 0.006634f
C635 B.n390 VSUBS 0.006634f
C636 B.n391 VSUBS 0.006634f
C637 B.n392 VSUBS 0.006634f
C638 B.n393 VSUBS 0.006634f
C639 B.n394 VSUBS 0.006634f
C640 B.n395 VSUBS 0.006634f
C641 B.n396 VSUBS 0.006634f
C642 B.n397 VSUBS 0.006634f
C643 B.n398 VSUBS 0.006634f
C644 B.n399 VSUBS 0.006634f
C645 B.n400 VSUBS 0.006634f
C646 B.n401 VSUBS 0.006634f
C647 B.n402 VSUBS 0.006634f
C648 B.n403 VSUBS 0.006634f
C649 B.n404 VSUBS 0.006634f
C650 B.n405 VSUBS 0.006634f
C651 B.n406 VSUBS 0.006634f
C652 B.n407 VSUBS 0.006634f
C653 B.n408 VSUBS 0.006634f
C654 B.n409 VSUBS 0.006634f
C655 B.n410 VSUBS 0.006634f
C656 B.n411 VSUBS 0.006634f
C657 B.n412 VSUBS 0.006634f
C658 B.n413 VSUBS 0.006634f
C659 B.n414 VSUBS 0.004585f
C660 B.n415 VSUBS 0.015371f
C661 B.n416 VSUBS 0.005366f
C662 B.n417 VSUBS 0.006634f
C663 B.n418 VSUBS 0.006634f
C664 B.n419 VSUBS 0.006634f
C665 B.n420 VSUBS 0.006634f
C666 B.n421 VSUBS 0.006634f
C667 B.n422 VSUBS 0.006634f
C668 B.n423 VSUBS 0.006634f
C669 B.n424 VSUBS 0.006634f
C670 B.n425 VSUBS 0.006634f
C671 B.n426 VSUBS 0.006634f
C672 B.n427 VSUBS 0.006634f
C673 B.n428 VSUBS 0.005366f
C674 B.n429 VSUBS 0.015371f
C675 B.n430 VSUBS 0.004585f
C676 B.n431 VSUBS 0.006634f
C677 B.n432 VSUBS 0.006634f
C678 B.n433 VSUBS 0.006634f
C679 B.n434 VSUBS 0.006634f
C680 B.n435 VSUBS 0.006634f
C681 B.n436 VSUBS 0.006634f
C682 B.n437 VSUBS 0.006634f
C683 B.n438 VSUBS 0.006634f
C684 B.n439 VSUBS 0.006634f
C685 B.n440 VSUBS 0.006634f
C686 B.n441 VSUBS 0.006634f
C687 B.n442 VSUBS 0.006634f
C688 B.n443 VSUBS 0.006634f
C689 B.n444 VSUBS 0.006634f
C690 B.n445 VSUBS 0.006634f
C691 B.n446 VSUBS 0.006634f
C692 B.n447 VSUBS 0.006634f
C693 B.n448 VSUBS 0.006634f
C694 B.n449 VSUBS 0.006634f
C695 B.n450 VSUBS 0.006634f
C696 B.n451 VSUBS 0.006634f
C697 B.n452 VSUBS 0.006634f
C698 B.n453 VSUBS 0.006634f
C699 B.n454 VSUBS 0.006634f
C700 B.n455 VSUBS 0.006634f
C701 B.n456 VSUBS 0.006634f
C702 B.n457 VSUBS 0.006634f
C703 B.n458 VSUBS 0.006634f
C704 B.n459 VSUBS 0.006634f
C705 B.n460 VSUBS 0.006634f
C706 B.n461 VSUBS 0.006634f
C707 B.n462 VSUBS 0.006634f
C708 B.n463 VSUBS 0.006634f
C709 B.n464 VSUBS 0.006634f
C710 B.n465 VSUBS 0.006634f
C711 B.n466 VSUBS 0.006634f
C712 B.n467 VSUBS 0.006634f
C713 B.n468 VSUBS 0.006634f
C714 B.n469 VSUBS 0.006634f
C715 B.n470 VSUBS 0.006634f
C716 B.n471 VSUBS 0.006634f
C717 B.n472 VSUBS 0.006634f
C718 B.n473 VSUBS 0.006634f
C719 B.n474 VSUBS 0.006634f
C720 B.n475 VSUBS 0.006634f
C721 B.n476 VSUBS 0.006634f
C722 B.n477 VSUBS 0.006634f
C723 B.n478 VSUBS 0.006634f
C724 B.n479 VSUBS 0.006634f
C725 B.n480 VSUBS 0.006634f
C726 B.n481 VSUBS 0.006634f
C727 B.n482 VSUBS 0.006634f
C728 B.n483 VSUBS 0.006634f
C729 B.n484 VSUBS 0.006634f
C730 B.n485 VSUBS 0.006634f
C731 B.n486 VSUBS 0.006634f
C732 B.n487 VSUBS 0.006634f
C733 B.n488 VSUBS 0.006634f
C734 B.n489 VSUBS 0.006634f
C735 B.n490 VSUBS 0.006634f
C736 B.n491 VSUBS 0.006634f
C737 B.n492 VSUBS 0.006634f
C738 B.n493 VSUBS 0.006634f
C739 B.n494 VSUBS 0.006634f
C740 B.n495 VSUBS 0.006634f
C741 B.n496 VSUBS 0.006634f
C742 B.n497 VSUBS 0.006634f
C743 B.n498 VSUBS 0.006634f
C744 B.n499 VSUBS 0.006634f
C745 B.n500 VSUBS 0.006634f
C746 B.n501 VSUBS 0.006634f
C747 B.n502 VSUBS 0.006634f
C748 B.n503 VSUBS 0.006634f
C749 B.n504 VSUBS 0.006634f
C750 B.n505 VSUBS 0.006634f
C751 B.n506 VSUBS 0.006634f
C752 B.n507 VSUBS 0.006634f
C753 B.n508 VSUBS 0.006634f
C754 B.n509 VSUBS 0.006634f
C755 B.n510 VSUBS 0.006634f
C756 B.n511 VSUBS 0.006634f
C757 B.n512 VSUBS 0.006634f
C758 B.n513 VSUBS 0.006634f
C759 B.n514 VSUBS 0.006634f
C760 B.n515 VSUBS 0.006634f
C761 B.n516 VSUBS 0.006634f
C762 B.n517 VSUBS 0.01628f
C763 B.n518 VSUBS 0.015525f
C764 B.n519 VSUBS 0.01628f
C765 B.n520 VSUBS 0.006634f
C766 B.n521 VSUBS 0.006634f
C767 B.n522 VSUBS 0.006634f
C768 B.n523 VSUBS 0.006634f
C769 B.n524 VSUBS 0.006634f
C770 B.n525 VSUBS 0.006634f
C771 B.n526 VSUBS 0.006634f
C772 B.n527 VSUBS 0.006634f
C773 B.n528 VSUBS 0.006634f
C774 B.n529 VSUBS 0.006634f
C775 B.n530 VSUBS 0.006634f
C776 B.n531 VSUBS 0.006634f
C777 B.n532 VSUBS 0.006634f
C778 B.n533 VSUBS 0.006634f
C779 B.n534 VSUBS 0.006634f
C780 B.n535 VSUBS 0.006634f
C781 B.n536 VSUBS 0.006634f
C782 B.n537 VSUBS 0.006634f
C783 B.n538 VSUBS 0.006634f
C784 B.n539 VSUBS 0.006634f
C785 B.n540 VSUBS 0.006634f
C786 B.n541 VSUBS 0.006634f
C787 B.n542 VSUBS 0.006634f
C788 B.n543 VSUBS 0.006634f
C789 B.n544 VSUBS 0.006634f
C790 B.n545 VSUBS 0.006634f
C791 B.n546 VSUBS 0.006634f
C792 B.n547 VSUBS 0.006634f
C793 B.n548 VSUBS 0.006634f
C794 B.n549 VSUBS 0.006634f
C795 B.n550 VSUBS 0.006634f
C796 B.n551 VSUBS 0.006634f
C797 B.n552 VSUBS 0.006634f
C798 B.n553 VSUBS 0.006634f
C799 B.n554 VSUBS 0.006634f
C800 B.n555 VSUBS 0.006634f
C801 B.n556 VSUBS 0.006634f
C802 B.n557 VSUBS 0.006634f
C803 B.n558 VSUBS 0.006634f
C804 B.n559 VSUBS 0.006634f
C805 B.n560 VSUBS 0.006634f
C806 B.n561 VSUBS 0.006634f
C807 B.n562 VSUBS 0.006634f
C808 B.n563 VSUBS 0.006634f
C809 B.n564 VSUBS 0.006634f
C810 B.n565 VSUBS 0.006634f
C811 B.n566 VSUBS 0.006634f
C812 B.n567 VSUBS 0.006634f
C813 B.n568 VSUBS 0.006634f
C814 B.n569 VSUBS 0.006634f
C815 B.n570 VSUBS 0.006634f
C816 B.n571 VSUBS 0.006634f
C817 B.n572 VSUBS 0.006634f
C818 B.n573 VSUBS 0.006634f
C819 B.n574 VSUBS 0.006634f
C820 B.n575 VSUBS 0.006634f
C821 B.n576 VSUBS 0.006634f
C822 B.n577 VSUBS 0.006634f
C823 B.n578 VSUBS 0.006634f
C824 B.n579 VSUBS 0.006634f
C825 B.n580 VSUBS 0.006634f
C826 B.n581 VSUBS 0.006634f
C827 B.n582 VSUBS 0.006634f
C828 B.n583 VSUBS 0.006634f
C829 B.n584 VSUBS 0.006634f
C830 B.n585 VSUBS 0.006634f
C831 B.n586 VSUBS 0.006634f
C832 B.n587 VSUBS 0.006634f
C833 B.n588 VSUBS 0.006634f
C834 B.n589 VSUBS 0.006634f
C835 B.n590 VSUBS 0.006634f
C836 B.n591 VSUBS 0.006634f
C837 B.n592 VSUBS 0.006634f
C838 B.n593 VSUBS 0.006634f
C839 B.n594 VSUBS 0.006634f
C840 B.n595 VSUBS 0.006634f
C841 B.n596 VSUBS 0.006634f
C842 B.n597 VSUBS 0.006634f
C843 B.n598 VSUBS 0.006634f
C844 B.n599 VSUBS 0.006634f
C845 B.n600 VSUBS 0.006634f
C846 B.n601 VSUBS 0.006634f
C847 B.n602 VSUBS 0.006634f
C848 B.n603 VSUBS 0.006634f
C849 B.n604 VSUBS 0.006634f
C850 B.n605 VSUBS 0.006634f
C851 B.n606 VSUBS 0.006634f
C852 B.n607 VSUBS 0.006634f
C853 B.n608 VSUBS 0.006634f
C854 B.n609 VSUBS 0.006634f
C855 B.n610 VSUBS 0.006634f
C856 B.n611 VSUBS 0.006634f
C857 B.n612 VSUBS 0.006634f
C858 B.n613 VSUBS 0.006634f
C859 B.n614 VSUBS 0.006634f
C860 B.n615 VSUBS 0.006634f
C861 B.n616 VSUBS 0.006634f
C862 B.n617 VSUBS 0.006634f
C863 B.n618 VSUBS 0.006634f
C864 B.n619 VSUBS 0.006634f
C865 B.n620 VSUBS 0.006634f
C866 B.n621 VSUBS 0.006634f
C867 B.n622 VSUBS 0.006634f
C868 B.n623 VSUBS 0.006634f
C869 B.n624 VSUBS 0.006634f
C870 B.n625 VSUBS 0.006634f
C871 B.n626 VSUBS 0.006634f
C872 B.n627 VSUBS 0.006634f
C873 B.n628 VSUBS 0.006634f
C874 B.n629 VSUBS 0.006634f
C875 B.n630 VSUBS 0.006634f
C876 B.n631 VSUBS 0.006634f
C877 B.n632 VSUBS 0.006634f
C878 B.n633 VSUBS 0.006634f
C879 B.n634 VSUBS 0.006634f
C880 B.n635 VSUBS 0.006634f
C881 B.n636 VSUBS 0.006634f
C882 B.n637 VSUBS 0.006634f
C883 B.n638 VSUBS 0.006634f
C884 B.n639 VSUBS 0.006634f
C885 B.n640 VSUBS 0.006634f
C886 B.n641 VSUBS 0.006634f
C887 B.n642 VSUBS 0.006634f
C888 B.n643 VSUBS 0.006634f
C889 B.n644 VSUBS 0.006634f
C890 B.n645 VSUBS 0.006634f
C891 B.n646 VSUBS 0.006634f
C892 B.n647 VSUBS 0.006634f
C893 B.n648 VSUBS 0.006634f
C894 B.n649 VSUBS 0.006634f
C895 B.n650 VSUBS 0.006634f
C896 B.n651 VSUBS 0.006634f
C897 B.n652 VSUBS 0.006634f
C898 B.n653 VSUBS 0.006634f
C899 B.n654 VSUBS 0.006634f
C900 B.n655 VSUBS 0.006634f
C901 B.n656 VSUBS 0.006634f
C902 B.n657 VSUBS 0.006634f
C903 B.n658 VSUBS 0.006634f
C904 B.n659 VSUBS 0.006634f
C905 B.n660 VSUBS 0.006634f
C906 B.n661 VSUBS 0.006634f
C907 B.n662 VSUBS 0.006634f
C908 B.n663 VSUBS 0.006634f
C909 B.n664 VSUBS 0.006634f
C910 B.n665 VSUBS 0.006634f
C911 B.n666 VSUBS 0.006634f
C912 B.n667 VSUBS 0.006634f
C913 B.n668 VSUBS 0.006634f
C914 B.n669 VSUBS 0.006634f
C915 B.n670 VSUBS 0.006634f
C916 B.n671 VSUBS 0.006634f
C917 B.n672 VSUBS 0.006634f
C918 B.n673 VSUBS 0.006634f
C919 B.n674 VSUBS 0.006634f
C920 B.n675 VSUBS 0.006634f
C921 B.n676 VSUBS 0.006634f
C922 B.n677 VSUBS 0.006634f
C923 B.n678 VSUBS 0.006634f
C924 B.n679 VSUBS 0.006634f
C925 B.n680 VSUBS 0.006634f
C926 B.n681 VSUBS 0.006634f
C927 B.n682 VSUBS 0.015525f
C928 B.n683 VSUBS 0.015525f
C929 B.n684 VSUBS 0.01628f
C930 B.n685 VSUBS 0.006634f
C931 B.n686 VSUBS 0.006634f
C932 B.n687 VSUBS 0.006634f
C933 B.n688 VSUBS 0.006634f
C934 B.n689 VSUBS 0.006634f
C935 B.n690 VSUBS 0.006634f
C936 B.n691 VSUBS 0.006634f
C937 B.n692 VSUBS 0.006634f
C938 B.n693 VSUBS 0.006634f
C939 B.n694 VSUBS 0.006634f
C940 B.n695 VSUBS 0.006634f
C941 B.n696 VSUBS 0.006634f
C942 B.n697 VSUBS 0.006634f
C943 B.n698 VSUBS 0.006634f
C944 B.n699 VSUBS 0.006634f
C945 B.n700 VSUBS 0.006634f
C946 B.n701 VSUBS 0.006634f
C947 B.n702 VSUBS 0.006634f
C948 B.n703 VSUBS 0.006634f
C949 B.n704 VSUBS 0.006634f
C950 B.n705 VSUBS 0.006634f
C951 B.n706 VSUBS 0.006634f
C952 B.n707 VSUBS 0.006634f
C953 B.n708 VSUBS 0.006634f
C954 B.n709 VSUBS 0.006634f
C955 B.n710 VSUBS 0.006634f
C956 B.n711 VSUBS 0.006634f
C957 B.n712 VSUBS 0.006634f
C958 B.n713 VSUBS 0.006634f
C959 B.n714 VSUBS 0.006634f
C960 B.n715 VSUBS 0.006634f
C961 B.n716 VSUBS 0.006634f
C962 B.n717 VSUBS 0.006634f
C963 B.n718 VSUBS 0.006634f
C964 B.n719 VSUBS 0.006634f
C965 B.n720 VSUBS 0.006634f
C966 B.n721 VSUBS 0.006634f
C967 B.n722 VSUBS 0.006634f
C968 B.n723 VSUBS 0.006634f
C969 B.n724 VSUBS 0.006634f
C970 B.n725 VSUBS 0.006634f
C971 B.n726 VSUBS 0.006634f
C972 B.n727 VSUBS 0.006634f
C973 B.n728 VSUBS 0.006634f
C974 B.n729 VSUBS 0.006634f
C975 B.n730 VSUBS 0.006634f
C976 B.n731 VSUBS 0.006634f
C977 B.n732 VSUBS 0.006634f
C978 B.n733 VSUBS 0.006634f
C979 B.n734 VSUBS 0.006634f
C980 B.n735 VSUBS 0.006634f
C981 B.n736 VSUBS 0.006634f
C982 B.n737 VSUBS 0.006634f
C983 B.n738 VSUBS 0.006634f
C984 B.n739 VSUBS 0.006634f
C985 B.n740 VSUBS 0.006634f
C986 B.n741 VSUBS 0.006634f
C987 B.n742 VSUBS 0.006634f
C988 B.n743 VSUBS 0.006634f
C989 B.n744 VSUBS 0.006634f
C990 B.n745 VSUBS 0.006634f
C991 B.n746 VSUBS 0.006634f
C992 B.n747 VSUBS 0.006634f
C993 B.n748 VSUBS 0.006634f
C994 B.n749 VSUBS 0.006634f
C995 B.n750 VSUBS 0.006634f
C996 B.n751 VSUBS 0.006634f
C997 B.n752 VSUBS 0.006634f
C998 B.n753 VSUBS 0.006634f
C999 B.n754 VSUBS 0.006634f
C1000 B.n755 VSUBS 0.006634f
C1001 B.n756 VSUBS 0.006634f
C1002 B.n757 VSUBS 0.006634f
C1003 B.n758 VSUBS 0.006634f
C1004 B.n759 VSUBS 0.006634f
C1005 B.n760 VSUBS 0.006634f
C1006 B.n761 VSUBS 0.006634f
C1007 B.n762 VSUBS 0.006634f
C1008 B.n763 VSUBS 0.006634f
C1009 B.n764 VSUBS 0.006634f
C1010 B.n765 VSUBS 0.006634f
C1011 B.n766 VSUBS 0.006634f
C1012 B.n767 VSUBS 0.006634f
C1013 B.n768 VSUBS 0.006634f
C1014 B.n769 VSUBS 0.006634f
C1015 B.n770 VSUBS 0.006634f
C1016 B.n771 VSUBS 0.004585f
C1017 B.n772 VSUBS 0.015371f
C1018 B.n773 VSUBS 0.005366f
C1019 B.n774 VSUBS 0.006634f
C1020 B.n775 VSUBS 0.006634f
C1021 B.n776 VSUBS 0.006634f
C1022 B.n777 VSUBS 0.006634f
C1023 B.n778 VSUBS 0.006634f
C1024 B.n779 VSUBS 0.006634f
C1025 B.n780 VSUBS 0.006634f
C1026 B.n781 VSUBS 0.006634f
C1027 B.n782 VSUBS 0.006634f
C1028 B.n783 VSUBS 0.006634f
C1029 B.n784 VSUBS 0.006634f
C1030 B.n785 VSUBS 0.005366f
C1031 B.n786 VSUBS 0.006634f
C1032 B.n787 VSUBS 0.006634f
C1033 B.n788 VSUBS 0.006634f
C1034 B.n789 VSUBS 0.006634f
C1035 B.n790 VSUBS 0.006634f
C1036 B.n791 VSUBS 0.006634f
C1037 B.n792 VSUBS 0.006634f
C1038 B.n793 VSUBS 0.006634f
C1039 B.n794 VSUBS 0.006634f
C1040 B.n795 VSUBS 0.006634f
C1041 B.n796 VSUBS 0.006634f
C1042 B.n797 VSUBS 0.006634f
C1043 B.n798 VSUBS 0.006634f
C1044 B.n799 VSUBS 0.006634f
C1045 B.n800 VSUBS 0.006634f
C1046 B.n801 VSUBS 0.006634f
C1047 B.n802 VSUBS 0.006634f
C1048 B.n803 VSUBS 0.006634f
C1049 B.n804 VSUBS 0.006634f
C1050 B.n805 VSUBS 0.006634f
C1051 B.n806 VSUBS 0.006634f
C1052 B.n807 VSUBS 0.006634f
C1053 B.n808 VSUBS 0.006634f
C1054 B.n809 VSUBS 0.006634f
C1055 B.n810 VSUBS 0.006634f
C1056 B.n811 VSUBS 0.006634f
C1057 B.n812 VSUBS 0.006634f
C1058 B.n813 VSUBS 0.006634f
C1059 B.n814 VSUBS 0.006634f
C1060 B.n815 VSUBS 0.006634f
C1061 B.n816 VSUBS 0.006634f
C1062 B.n817 VSUBS 0.006634f
C1063 B.n818 VSUBS 0.006634f
C1064 B.n819 VSUBS 0.006634f
C1065 B.n820 VSUBS 0.006634f
C1066 B.n821 VSUBS 0.006634f
C1067 B.n822 VSUBS 0.006634f
C1068 B.n823 VSUBS 0.006634f
C1069 B.n824 VSUBS 0.006634f
C1070 B.n825 VSUBS 0.006634f
C1071 B.n826 VSUBS 0.006634f
C1072 B.n827 VSUBS 0.006634f
C1073 B.n828 VSUBS 0.006634f
C1074 B.n829 VSUBS 0.006634f
C1075 B.n830 VSUBS 0.006634f
C1076 B.n831 VSUBS 0.006634f
C1077 B.n832 VSUBS 0.006634f
C1078 B.n833 VSUBS 0.006634f
C1079 B.n834 VSUBS 0.006634f
C1080 B.n835 VSUBS 0.006634f
C1081 B.n836 VSUBS 0.006634f
C1082 B.n837 VSUBS 0.006634f
C1083 B.n838 VSUBS 0.006634f
C1084 B.n839 VSUBS 0.006634f
C1085 B.n840 VSUBS 0.006634f
C1086 B.n841 VSUBS 0.006634f
C1087 B.n842 VSUBS 0.006634f
C1088 B.n843 VSUBS 0.006634f
C1089 B.n844 VSUBS 0.006634f
C1090 B.n845 VSUBS 0.006634f
C1091 B.n846 VSUBS 0.006634f
C1092 B.n847 VSUBS 0.006634f
C1093 B.n848 VSUBS 0.006634f
C1094 B.n849 VSUBS 0.006634f
C1095 B.n850 VSUBS 0.006634f
C1096 B.n851 VSUBS 0.006634f
C1097 B.n852 VSUBS 0.006634f
C1098 B.n853 VSUBS 0.006634f
C1099 B.n854 VSUBS 0.006634f
C1100 B.n855 VSUBS 0.006634f
C1101 B.n856 VSUBS 0.006634f
C1102 B.n857 VSUBS 0.006634f
C1103 B.n858 VSUBS 0.006634f
C1104 B.n859 VSUBS 0.006634f
C1105 B.n860 VSUBS 0.006634f
C1106 B.n861 VSUBS 0.006634f
C1107 B.n862 VSUBS 0.006634f
C1108 B.n863 VSUBS 0.006634f
C1109 B.n864 VSUBS 0.006634f
C1110 B.n865 VSUBS 0.006634f
C1111 B.n866 VSUBS 0.006634f
C1112 B.n867 VSUBS 0.006634f
C1113 B.n868 VSUBS 0.006634f
C1114 B.n869 VSUBS 0.006634f
C1115 B.n870 VSUBS 0.006634f
C1116 B.n871 VSUBS 0.006634f
C1117 B.n872 VSUBS 0.006634f
C1118 B.n873 VSUBS 0.006634f
C1119 B.n874 VSUBS 0.01628f
C1120 B.n875 VSUBS 0.015525f
C1121 B.n876 VSUBS 0.015525f
C1122 B.n877 VSUBS 0.006634f
C1123 B.n878 VSUBS 0.006634f
C1124 B.n879 VSUBS 0.006634f
C1125 B.n880 VSUBS 0.006634f
C1126 B.n881 VSUBS 0.006634f
C1127 B.n882 VSUBS 0.006634f
C1128 B.n883 VSUBS 0.006634f
C1129 B.n884 VSUBS 0.006634f
C1130 B.n885 VSUBS 0.006634f
C1131 B.n886 VSUBS 0.006634f
C1132 B.n887 VSUBS 0.006634f
C1133 B.n888 VSUBS 0.006634f
C1134 B.n889 VSUBS 0.006634f
C1135 B.n890 VSUBS 0.006634f
C1136 B.n891 VSUBS 0.006634f
C1137 B.n892 VSUBS 0.006634f
C1138 B.n893 VSUBS 0.006634f
C1139 B.n894 VSUBS 0.006634f
C1140 B.n895 VSUBS 0.006634f
C1141 B.n896 VSUBS 0.006634f
C1142 B.n897 VSUBS 0.006634f
C1143 B.n898 VSUBS 0.006634f
C1144 B.n899 VSUBS 0.006634f
C1145 B.n900 VSUBS 0.006634f
C1146 B.n901 VSUBS 0.006634f
C1147 B.n902 VSUBS 0.006634f
C1148 B.n903 VSUBS 0.006634f
C1149 B.n904 VSUBS 0.006634f
C1150 B.n905 VSUBS 0.006634f
C1151 B.n906 VSUBS 0.006634f
C1152 B.n907 VSUBS 0.006634f
C1153 B.n908 VSUBS 0.006634f
C1154 B.n909 VSUBS 0.006634f
C1155 B.n910 VSUBS 0.006634f
C1156 B.n911 VSUBS 0.006634f
C1157 B.n912 VSUBS 0.006634f
C1158 B.n913 VSUBS 0.006634f
C1159 B.n914 VSUBS 0.006634f
C1160 B.n915 VSUBS 0.006634f
C1161 B.n916 VSUBS 0.006634f
C1162 B.n917 VSUBS 0.006634f
C1163 B.n918 VSUBS 0.006634f
C1164 B.n919 VSUBS 0.006634f
C1165 B.n920 VSUBS 0.006634f
C1166 B.n921 VSUBS 0.006634f
C1167 B.n922 VSUBS 0.006634f
C1168 B.n923 VSUBS 0.006634f
C1169 B.n924 VSUBS 0.006634f
C1170 B.n925 VSUBS 0.006634f
C1171 B.n926 VSUBS 0.006634f
C1172 B.n927 VSUBS 0.006634f
C1173 B.n928 VSUBS 0.006634f
C1174 B.n929 VSUBS 0.006634f
C1175 B.n930 VSUBS 0.006634f
C1176 B.n931 VSUBS 0.006634f
C1177 B.n932 VSUBS 0.006634f
C1178 B.n933 VSUBS 0.006634f
C1179 B.n934 VSUBS 0.006634f
C1180 B.n935 VSUBS 0.006634f
C1181 B.n936 VSUBS 0.006634f
C1182 B.n937 VSUBS 0.006634f
C1183 B.n938 VSUBS 0.006634f
C1184 B.n939 VSUBS 0.006634f
C1185 B.n940 VSUBS 0.006634f
C1186 B.n941 VSUBS 0.006634f
C1187 B.n942 VSUBS 0.006634f
C1188 B.n943 VSUBS 0.006634f
C1189 B.n944 VSUBS 0.006634f
C1190 B.n945 VSUBS 0.006634f
C1191 B.n946 VSUBS 0.006634f
C1192 B.n947 VSUBS 0.006634f
C1193 B.n948 VSUBS 0.006634f
C1194 B.n949 VSUBS 0.006634f
C1195 B.n950 VSUBS 0.006634f
C1196 B.n951 VSUBS 0.006634f
C1197 B.n952 VSUBS 0.006634f
C1198 B.n953 VSUBS 0.006634f
C1199 B.n954 VSUBS 0.006634f
C1200 B.n955 VSUBS 0.008657f
C1201 B.n956 VSUBS 0.009222f
C1202 B.n957 VSUBS 0.018339f
.ends

