* NGSPICE file created from diff_pair_sample_0302.ext - technology: sky130A

.subckt diff_pair_sample_0302 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=1.43
X1 VTAIL.t14 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X2 VDD2.t4 VN.t1 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X3 VTAIL.t12 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=1.43
X4 VTAIL.t3 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=1.43
X5 VDD2.t0 VN.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X6 VTAIL.t1 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=1.43
X7 VTAIL.t2 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X8 VDD1.t4 VP.t3 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X9 VDD1.t3 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=1.43
X10 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=1.43
X11 VTAIL.t10 VN.t4 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=1.43
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=1.43
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=1.43
X14 VDD1.t2 VP.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X15 VDD2.t2 VN.t5 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=1.43
X16 VTAIL.t5 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X17 VTAIL.t8 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=1.43
X18 VDD1.t0 VP.t7 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=1.43
X19 VDD2.t3 VN.t7 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=1.43
R0 B.n548 B.n547 585
R1 B.n548 B.n64 585
R2 B.n551 B.n550 585
R3 B.n552 B.n112 585
R4 B.n554 B.n553 585
R5 B.n556 B.n111 585
R6 B.n559 B.n558 585
R7 B.n560 B.n110 585
R8 B.n562 B.n561 585
R9 B.n564 B.n109 585
R10 B.n567 B.n566 585
R11 B.n568 B.n108 585
R12 B.n570 B.n569 585
R13 B.n572 B.n107 585
R14 B.n575 B.n574 585
R15 B.n576 B.n106 585
R16 B.n578 B.n577 585
R17 B.n580 B.n105 585
R18 B.n583 B.n582 585
R19 B.n584 B.n104 585
R20 B.n586 B.n585 585
R21 B.n588 B.n103 585
R22 B.n591 B.n590 585
R23 B.n592 B.n102 585
R24 B.n594 B.n593 585
R25 B.n596 B.n101 585
R26 B.n599 B.n598 585
R27 B.n600 B.n100 585
R28 B.n602 B.n601 585
R29 B.n604 B.n99 585
R30 B.n607 B.n606 585
R31 B.n608 B.n98 585
R32 B.n610 B.n609 585
R33 B.n612 B.n97 585
R34 B.n615 B.n614 585
R35 B.n616 B.n96 585
R36 B.n618 B.n617 585
R37 B.n620 B.n95 585
R38 B.n623 B.n622 585
R39 B.n624 B.n92 585
R40 B.n627 B.n626 585
R41 B.n629 B.n91 585
R42 B.n632 B.n631 585
R43 B.n633 B.n90 585
R44 B.n635 B.n634 585
R45 B.n637 B.n89 585
R46 B.n640 B.n639 585
R47 B.n641 B.n85 585
R48 B.n643 B.n642 585
R49 B.n645 B.n84 585
R50 B.n648 B.n647 585
R51 B.n649 B.n83 585
R52 B.n651 B.n650 585
R53 B.n653 B.n82 585
R54 B.n656 B.n655 585
R55 B.n657 B.n81 585
R56 B.n659 B.n658 585
R57 B.n661 B.n80 585
R58 B.n664 B.n663 585
R59 B.n665 B.n79 585
R60 B.n667 B.n666 585
R61 B.n669 B.n78 585
R62 B.n672 B.n671 585
R63 B.n673 B.n77 585
R64 B.n675 B.n674 585
R65 B.n677 B.n76 585
R66 B.n680 B.n679 585
R67 B.n681 B.n75 585
R68 B.n683 B.n682 585
R69 B.n685 B.n74 585
R70 B.n688 B.n687 585
R71 B.n689 B.n73 585
R72 B.n691 B.n690 585
R73 B.n693 B.n72 585
R74 B.n696 B.n695 585
R75 B.n697 B.n71 585
R76 B.n699 B.n698 585
R77 B.n701 B.n70 585
R78 B.n704 B.n703 585
R79 B.n705 B.n69 585
R80 B.n707 B.n706 585
R81 B.n709 B.n68 585
R82 B.n712 B.n711 585
R83 B.n713 B.n67 585
R84 B.n715 B.n714 585
R85 B.n717 B.n66 585
R86 B.n720 B.n719 585
R87 B.n721 B.n65 585
R88 B.n546 B.n63 585
R89 B.n724 B.n63 585
R90 B.n545 B.n62 585
R91 B.n725 B.n62 585
R92 B.n544 B.n61 585
R93 B.n726 B.n61 585
R94 B.n543 B.n542 585
R95 B.n542 B.n57 585
R96 B.n541 B.n56 585
R97 B.n732 B.n56 585
R98 B.n540 B.n55 585
R99 B.n733 B.n55 585
R100 B.n539 B.n54 585
R101 B.n734 B.n54 585
R102 B.n538 B.n537 585
R103 B.n537 B.n50 585
R104 B.n536 B.n49 585
R105 B.n740 B.n49 585
R106 B.n535 B.n48 585
R107 B.n741 B.n48 585
R108 B.n534 B.n47 585
R109 B.n742 B.n47 585
R110 B.n533 B.n532 585
R111 B.n532 B.n43 585
R112 B.n531 B.n42 585
R113 B.n748 B.n42 585
R114 B.n530 B.n41 585
R115 B.n749 B.n41 585
R116 B.n529 B.n40 585
R117 B.n750 B.n40 585
R118 B.n528 B.n527 585
R119 B.n527 B.n36 585
R120 B.n526 B.n35 585
R121 B.n756 B.n35 585
R122 B.n525 B.n34 585
R123 B.n757 B.n34 585
R124 B.n524 B.n33 585
R125 B.n758 B.n33 585
R126 B.n523 B.n522 585
R127 B.n522 B.n32 585
R128 B.n521 B.n28 585
R129 B.n764 B.n28 585
R130 B.n520 B.n27 585
R131 B.n765 B.n27 585
R132 B.n519 B.n26 585
R133 B.n766 B.n26 585
R134 B.n518 B.n517 585
R135 B.n517 B.n22 585
R136 B.n516 B.n21 585
R137 B.n772 B.n21 585
R138 B.n515 B.n20 585
R139 B.n773 B.n20 585
R140 B.n514 B.n19 585
R141 B.n774 B.n19 585
R142 B.n513 B.n512 585
R143 B.n512 B.n15 585
R144 B.n511 B.n14 585
R145 B.n780 B.n14 585
R146 B.n510 B.n13 585
R147 B.n781 B.n13 585
R148 B.n509 B.n12 585
R149 B.n782 B.n12 585
R150 B.n508 B.n507 585
R151 B.n507 B.n8 585
R152 B.n506 B.n7 585
R153 B.n788 B.n7 585
R154 B.n505 B.n6 585
R155 B.n789 B.n6 585
R156 B.n504 B.n5 585
R157 B.n790 B.n5 585
R158 B.n503 B.n502 585
R159 B.n502 B.n4 585
R160 B.n501 B.n113 585
R161 B.n501 B.n500 585
R162 B.n491 B.n114 585
R163 B.n115 B.n114 585
R164 B.n493 B.n492 585
R165 B.n494 B.n493 585
R166 B.n490 B.n119 585
R167 B.n123 B.n119 585
R168 B.n489 B.n488 585
R169 B.n488 B.n487 585
R170 B.n121 B.n120 585
R171 B.n122 B.n121 585
R172 B.n480 B.n479 585
R173 B.n481 B.n480 585
R174 B.n478 B.n128 585
R175 B.n128 B.n127 585
R176 B.n477 B.n476 585
R177 B.n476 B.n475 585
R178 B.n130 B.n129 585
R179 B.n131 B.n130 585
R180 B.n468 B.n467 585
R181 B.n469 B.n468 585
R182 B.n466 B.n136 585
R183 B.n136 B.n135 585
R184 B.n465 B.n464 585
R185 B.n464 B.n463 585
R186 B.n138 B.n137 585
R187 B.n456 B.n138 585
R188 B.n455 B.n454 585
R189 B.n457 B.n455 585
R190 B.n453 B.n143 585
R191 B.n143 B.n142 585
R192 B.n452 B.n451 585
R193 B.n451 B.n450 585
R194 B.n145 B.n144 585
R195 B.n146 B.n145 585
R196 B.n443 B.n442 585
R197 B.n444 B.n443 585
R198 B.n441 B.n151 585
R199 B.n151 B.n150 585
R200 B.n440 B.n439 585
R201 B.n439 B.n438 585
R202 B.n153 B.n152 585
R203 B.n154 B.n153 585
R204 B.n431 B.n430 585
R205 B.n432 B.n431 585
R206 B.n429 B.n159 585
R207 B.n159 B.n158 585
R208 B.n428 B.n427 585
R209 B.n427 B.n426 585
R210 B.n161 B.n160 585
R211 B.n162 B.n161 585
R212 B.n419 B.n418 585
R213 B.n420 B.n419 585
R214 B.n417 B.n166 585
R215 B.n170 B.n166 585
R216 B.n416 B.n415 585
R217 B.n415 B.n414 585
R218 B.n168 B.n167 585
R219 B.n169 B.n168 585
R220 B.n407 B.n406 585
R221 B.n408 B.n407 585
R222 B.n405 B.n175 585
R223 B.n175 B.n174 585
R224 B.n404 B.n403 585
R225 B.n403 B.n402 585
R226 B.n399 B.n179 585
R227 B.n398 B.n397 585
R228 B.n395 B.n180 585
R229 B.n395 B.n178 585
R230 B.n394 B.n393 585
R231 B.n392 B.n391 585
R232 B.n390 B.n182 585
R233 B.n388 B.n387 585
R234 B.n386 B.n183 585
R235 B.n385 B.n384 585
R236 B.n382 B.n184 585
R237 B.n380 B.n379 585
R238 B.n378 B.n185 585
R239 B.n377 B.n376 585
R240 B.n374 B.n186 585
R241 B.n372 B.n371 585
R242 B.n370 B.n187 585
R243 B.n369 B.n368 585
R244 B.n366 B.n188 585
R245 B.n364 B.n363 585
R246 B.n362 B.n189 585
R247 B.n361 B.n360 585
R248 B.n358 B.n190 585
R249 B.n356 B.n355 585
R250 B.n354 B.n191 585
R251 B.n353 B.n352 585
R252 B.n350 B.n192 585
R253 B.n348 B.n347 585
R254 B.n346 B.n193 585
R255 B.n345 B.n344 585
R256 B.n342 B.n194 585
R257 B.n340 B.n339 585
R258 B.n338 B.n195 585
R259 B.n337 B.n336 585
R260 B.n334 B.n196 585
R261 B.n332 B.n331 585
R262 B.n330 B.n197 585
R263 B.n329 B.n328 585
R264 B.n326 B.n198 585
R265 B.n324 B.n323 585
R266 B.n321 B.n199 585
R267 B.n320 B.n319 585
R268 B.n317 B.n202 585
R269 B.n315 B.n314 585
R270 B.n313 B.n203 585
R271 B.n312 B.n311 585
R272 B.n309 B.n204 585
R273 B.n307 B.n306 585
R274 B.n305 B.n205 585
R275 B.n303 B.n302 585
R276 B.n300 B.n208 585
R277 B.n298 B.n297 585
R278 B.n296 B.n209 585
R279 B.n295 B.n294 585
R280 B.n292 B.n210 585
R281 B.n290 B.n289 585
R282 B.n288 B.n211 585
R283 B.n287 B.n286 585
R284 B.n284 B.n212 585
R285 B.n282 B.n281 585
R286 B.n280 B.n213 585
R287 B.n279 B.n278 585
R288 B.n276 B.n214 585
R289 B.n274 B.n273 585
R290 B.n272 B.n215 585
R291 B.n271 B.n270 585
R292 B.n268 B.n216 585
R293 B.n266 B.n265 585
R294 B.n264 B.n217 585
R295 B.n263 B.n262 585
R296 B.n260 B.n218 585
R297 B.n258 B.n257 585
R298 B.n256 B.n219 585
R299 B.n255 B.n254 585
R300 B.n252 B.n220 585
R301 B.n250 B.n249 585
R302 B.n248 B.n221 585
R303 B.n247 B.n246 585
R304 B.n244 B.n222 585
R305 B.n242 B.n241 585
R306 B.n240 B.n223 585
R307 B.n239 B.n238 585
R308 B.n236 B.n224 585
R309 B.n234 B.n233 585
R310 B.n232 B.n225 585
R311 B.n231 B.n230 585
R312 B.n228 B.n226 585
R313 B.n177 B.n176 585
R314 B.n401 B.n400 585
R315 B.n402 B.n401 585
R316 B.n173 B.n172 585
R317 B.n174 B.n173 585
R318 B.n410 B.n409 585
R319 B.n409 B.n408 585
R320 B.n411 B.n171 585
R321 B.n171 B.n169 585
R322 B.n413 B.n412 585
R323 B.n414 B.n413 585
R324 B.n165 B.n164 585
R325 B.n170 B.n165 585
R326 B.n422 B.n421 585
R327 B.n421 B.n420 585
R328 B.n423 B.n163 585
R329 B.n163 B.n162 585
R330 B.n425 B.n424 585
R331 B.n426 B.n425 585
R332 B.n157 B.n156 585
R333 B.n158 B.n157 585
R334 B.n434 B.n433 585
R335 B.n433 B.n432 585
R336 B.n435 B.n155 585
R337 B.n155 B.n154 585
R338 B.n437 B.n436 585
R339 B.n438 B.n437 585
R340 B.n149 B.n148 585
R341 B.n150 B.n149 585
R342 B.n446 B.n445 585
R343 B.n445 B.n444 585
R344 B.n447 B.n147 585
R345 B.n147 B.n146 585
R346 B.n449 B.n448 585
R347 B.n450 B.n449 585
R348 B.n141 B.n140 585
R349 B.n142 B.n141 585
R350 B.n459 B.n458 585
R351 B.n458 B.n457 585
R352 B.n460 B.n139 585
R353 B.n456 B.n139 585
R354 B.n462 B.n461 585
R355 B.n463 B.n462 585
R356 B.n134 B.n133 585
R357 B.n135 B.n134 585
R358 B.n471 B.n470 585
R359 B.n470 B.n469 585
R360 B.n472 B.n132 585
R361 B.n132 B.n131 585
R362 B.n474 B.n473 585
R363 B.n475 B.n474 585
R364 B.n126 B.n125 585
R365 B.n127 B.n126 585
R366 B.n483 B.n482 585
R367 B.n482 B.n481 585
R368 B.n484 B.n124 585
R369 B.n124 B.n122 585
R370 B.n486 B.n485 585
R371 B.n487 B.n486 585
R372 B.n118 B.n117 585
R373 B.n123 B.n118 585
R374 B.n496 B.n495 585
R375 B.n495 B.n494 585
R376 B.n497 B.n116 585
R377 B.n116 B.n115 585
R378 B.n499 B.n498 585
R379 B.n500 B.n499 585
R380 B.n2 B.n0 585
R381 B.n4 B.n2 585
R382 B.n3 B.n1 585
R383 B.n789 B.n3 585
R384 B.n787 B.n786 585
R385 B.n788 B.n787 585
R386 B.n785 B.n9 585
R387 B.n9 B.n8 585
R388 B.n784 B.n783 585
R389 B.n783 B.n782 585
R390 B.n11 B.n10 585
R391 B.n781 B.n11 585
R392 B.n779 B.n778 585
R393 B.n780 B.n779 585
R394 B.n777 B.n16 585
R395 B.n16 B.n15 585
R396 B.n776 B.n775 585
R397 B.n775 B.n774 585
R398 B.n18 B.n17 585
R399 B.n773 B.n18 585
R400 B.n771 B.n770 585
R401 B.n772 B.n771 585
R402 B.n769 B.n23 585
R403 B.n23 B.n22 585
R404 B.n768 B.n767 585
R405 B.n767 B.n766 585
R406 B.n25 B.n24 585
R407 B.n765 B.n25 585
R408 B.n763 B.n762 585
R409 B.n764 B.n763 585
R410 B.n761 B.n29 585
R411 B.n32 B.n29 585
R412 B.n760 B.n759 585
R413 B.n759 B.n758 585
R414 B.n31 B.n30 585
R415 B.n757 B.n31 585
R416 B.n755 B.n754 585
R417 B.n756 B.n755 585
R418 B.n753 B.n37 585
R419 B.n37 B.n36 585
R420 B.n752 B.n751 585
R421 B.n751 B.n750 585
R422 B.n39 B.n38 585
R423 B.n749 B.n39 585
R424 B.n747 B.n746 585
R425 B.n748 B.n747 585
R426 B.n745 B.n44 585
R427 B.n44 B.n43 585
R428 B.n744 B.n743 585
R429 B.n743 B.n742 585
R430 B.n46 B.n45 585
R431 B.n741 B.n46 585
R432 B.n739 B.n738 585
R433 B.n740 B.n739 585
R434 B.n737 B.n51 585
R435 B.n51 B.n50 585
R436 B.n736 B.n735 585
R437 B.n735 B.n734 585
R438 B.n53 B.n52 585
R439 B.n733 B.n53 585
R440 B.n731 B.n730 585
R441 B.n732 B.n731 585
R442 B.n729 B.n58 585
R443 B.n58 B.n57 585
R444 B.n728 B.n727 585
R445 B.n727 B.n726 585
R446 B.n60 B.n59 585
R447 B.n725 B.n60 585
R448 B.n723 B.n722 585
R449 B.n724 B.n723 585
R450 B.n792 B.n791 585
R451 B.n791 B.n790 585
R452 B.n401 B.n179 478.086
R453 B.n723 B.n65 478.086
R454 B.n403 B.n177 478.086
R455 B.n548 B.n63 478.086
R456 B.n206 B.t12 390.048
R457 B.n200 B.t16 390.048
R458 B.n86 B.t8 390.048
R459 B.n93 B.t19 390.048
R460 B.n549 B.n64 256.663
R461 B.n555 B.n64 256.663
R462 B.n557 B.n64 256.663
R463 B.n563 B.n64 256.663
R464 B.n565 B.n64 256.663
R465 B.n571 B.n64 256.663
R466 B.n573 B.n64 256.663
R467 B.n579 B.n64 256.663
R468 B.n581 B.n64 256.663
R469 B.n587 B.n64 256.663
R470 B.n589 B.n64 256.663
R471 B.n595 B.n64 256.663
R472 B.n597 B.n64 256.663
R473 B.n603 B.n64 256.663
R474 B.n605 B.n64 256.663
R475 B.n611 B.n64 256.663
R476 B.n613 B.n64 256.663
R477 B.n619 B.n64 256.663
R478 B.n621 B.n64 256.663
R479 B.n628 B.n64 256.663
R480 B.n630 B.n64 256.663
R481 B.n636 B.n64 256.663
R482 B.n638 B.n64 256.663
R483 B.n644 B.n64 256.663
R484 B.n646 B.n64 256.663
R485 B.n652 B.n64 256.663
R486 B.n654 B.n64 256.663
R487 B.n660 B.n64 256.663
R488 B.n662 B.n64 256.663
R489 B.n668 B.n64 256.663
R490 B.n670 B.n64 256.663
R491 B.n676 B.n64 256.663
R492 B.n678 B.n64 256.663
R493 B.n684 B.n64 256.663
R494 B.n686 B.n64 256.663
R495 B.n692 B.n64 256.663
R496 B.n694 B.n64 256.663
R497 B.n700 B.n64 256.663
R498 B.n702 B.n64 256.663
R499 B.n708 B.n64 256.663
R500 B.n710 B.n64 256.663
R501 B.n716 B.n64 256.663
R502 B.n718 B.n64 256.663
R503 B.n396 B.n178 256.663
R504 B.n181 B.n178 256.663
R505 B.n389 B.n178 256.663
R506 B.n383 B.n178 256.663
R507 B.n381 B.n178 256.663
R508 B.n375 B.n178 256.663
R509 B.n373 B.n178 256.663
R510 B.n367 B.n178 256.663
R511 B.n365 B.n178 256.663
R512 B.n359 B.n178 256.663
R513 B.n357 B.n178 256.663
R514 B.n351 B.n178 256.663
R515 B.n349 B.n178 256.663
R516 B.n343 B.n178 256.663
R517 B.n341 B.n178 256.663
R518 B.n335 B.n178 256.663
R519 B.n333 B.n178 256.663
R520 B.n327 B.n178 256.663
R521 B.n325 B.n178 256.663
R522 B.n318 B.n178 256.663
R523 B.n316 B.n178 256.663
R524 B.n310 B.n178 256.663
R525 B.n308 B.n178 256.663
R526 B.n301 B.n178 256.663
R527 B.n299 B.n178 256.663
R528 B.n293 B.n178 256.663
R529 B.n291 B.n178 256.663
R530 B.n285 B.n178 256.663
R531 B.n283 B.n178 256.663
R532 B.n277 B.n178 256.663
R533 B.n275 B.n178 256.663
R534 B.n269 B.n178 256.663
R535 B.n267 B.n178 256.663
R536 B.n261 B.n178 256.663
R537 B.n259 B.n178 256.663
R538 B.n253 B.n178 256.663
R539 B.n251 B.n178 256.663
R540 B.n245 B.n178 256.663
R541 B.n243 B.n178 256.663
R542 B.n237 B.n178 256.663
R543 B.n235 B.n178 256.663
R544 B.n229 B.n178 256.663
R545 B.n227 B.n178 256.663
R546 B.n401 B.n173 163.367
R547 B.n409 B.n173 163.367
R548 B.n409 B.n171 163.367
R549 B.n413 B.n171 163.367
R550 B.n413 B.n165 163.367
R551 B.n421 B.n165 163.367
R552 B.n421 B.n163 163.367
R553 B.n425 B.n163 163.367
R554 B.n425 B.n157 163.367
R555 B.n433 B.n157 163.367
R556 B.n433 B.n155 163.367
R557 B.n437 B.n155 163.367
R558 B.n437 B.n149 163.367
R559 B.n445 B.n149 163.367
R560 B.n445 B.n147 163.367
R561 B.n449 B.n147 163.367
R562 B.n449 B.n141 163.367
R563 B.n458 B.n141 163.367
R564 B.n458 B.n139 163.367
R565 B.n462 B.n139 163.367
R566 B.n462 B.n134 163.367
R567 B.n470 B.n134 163.367
R568 B.n470 B.n132 163.367
R569 B.n474 B.n132 163.367
R570 B.n474 B.n126 163.367
R571 B.n482 B.n126 163.367
R572 B.n482 B.n124 163.367
R573 B.n486 B.n124 163.367
R574 B.n486 B.n118 163.367
R575 B.n495 B.n118 163.367
R576 B.n495 B.n116 163.367
R577 B.n499 B.n116 163.367
R578 B.n499 B.n2 163.367
R579 B.n791 B.n2 163.367
R580 B.n791 B.n3 163.367
R581 B.n787 B.n3 163.367
R582 B.n787 B.n9 163.367
R583 B.n783 B.n9 163.367
R584 B.n783 B.n11 163.367
R585 B.n779 B.n11 163.367
R586 B.n779 B.n16 163.367
R587 B.n775 B.n16 163.367
R588 B.n775 B.n18 163.367
R589 B.n771 B.n18 163.367
R590 B.n771 B.n23 163.367
R591 B.n767 B.n23 163.367
R592 B.n767 B.n25 163.367
R593 B.n763 B.n25 163.367
R594 B.n763 B.n29 163.367
R595 B.n759 B.n29 163.367
R596 B.n759 B.n31 163.367
R597 B.n755 B.n31 163.367
R598 B.n755 B.n37 163.367
R599 B.n751 B.n37 163.367
R600 B.n751 B.n39 163.367
R601 B.n747 B.n39 163.367
R602 B.n747 B.n44 163.367
R603 B.n743 B.n44 163.367
R604 B.n743 B.n46 163.367
R605 B.n739 B.n46 163.367
R606 B.n739 B.n51 163.367
R607 B.n735 B.n51 163.367
R608 B.n735 B.n53 163.367
R609 B.n731 B.n53 163.367
R610 B.n731 B.n58 163.367
R611 B.n727 B.n58 163.367
R612 B.n727 B.n60 163.367
R613 B.n723 B.n60 163.367
R614 B.n397 B.n395 163.367
R615 B.n395 B.n394 163.367
R616 B.n391 B.n390 163.367
R617 B.n388 B.n183 163.367
R618 B.n384 B.n382 163.367
R619 B.n380 B.n185 163.367
R620 B.n376 B.n374 163.367
R621 B.n372 B.n187 163.367
R622 B.n368 B.n366 163.367
R623 B.n364 B.n189 163.367
R624 B.n360 B.n358 163.367
R625 B.n356 B.n191 163.367
R626 B.n352 B.n350 163.367
R627 B.n348 B.n193 163.367
R628 B.n344 B.n342 163.367
R629 B.n340 B.n195 163.367
R630 B.n336 B.n334 163.367
R631 B.n332 B.n197 163.367
R632 B.n328 B.n326 163.367
R633 B.n324 B.n199 163.367
R634 B.n319 B.n317 163.367
R635 B.n315 B.n203 163.367
R636 B.n311 B.n309 163.367
R637 B.n307 B.n205 163.367
R638 B.n302 B.n300 163.367
R639 B.n298 B.n209 163.367
R640 B.n294 B.n292 163.367
R641 B.n290 B.n211 163.367
R642 B.n286 B.n284 163.367
R643 B.n282 B.n213 163.367
R644 B.n278 B.n276 163.367
R645 B.n274 B.n215 163.367
R646 B.n270 B.n268 163.367
R647 B.n266 B.n217 163.367
R648 B.n262 B.n260 163.367
R649 B.n258 B.n219 163.367
R650 B.n254 B.n252 163.367
R651 B.n250 B.n221 163.367
R652 B.n246 B.n244 163.367
R653 B.n242 B.n223 163.367
R654 B.n238 B.n236 163.367
R655 B.n234 B.n225 163.367
R656 B.n230 B.n228 163.367
R657 B.n403 B.n175 163.367
R658 B.n407 B.n175 163.367
R659 B.n407 B.n168 163.367
R660 B.n415 B.n168 163.367
R661 B.n415 B.n166 163.367
R662 B.n419 B.n166 163.367
R663 B.n419 B.n161 163.367
R664 B.n427 B.n161 163.367
R665 B.n427 B.n159 163.367
R666 B.n431 B.n159 163.367
R667 B.n431 B.n153 163.367
R668 B.n439 B.n153 163.367
R669 B.n439 B.n151 163.367
R670 B.n443 B.n151 163.367
R671 B.n443 B.n145 163.367
R672 B.n451 B.n145 163.367
R673 B.n451 B.n143 163.367
R674 B.n455 B.n143 163.367
R675 B.n455 B.n138 163.367
R676 B.n464 B.n138 163.367
R677 B.n464 B.n136 163.367
R678 B.n468 B.n136 163.367
R679 B.n468 B.n130 163.367
R680 B.n476 B.n130 163.367
R681 B.n476 B.n128 163.367
R682 B.n480 B.n128 163.367
R683 B.n480 B.n121 163.367
R684 B.n488 B.n121 163.367
R685 B.n488 B.n119 163.367
R686 B.n493 B.n119 163.367
R687 B.n493 B.n114 163.367
R688 B.n501 B.n114 163.367
R689 B.n502 B.n501 163.367
R690 B.n502 B.n5 163.367
R691 B.n6 B.n5 163.367
R692 B.n7 B.n6 163.367
R693 B.n507 B.n7 163.367
R694 B.n507 B.n12 163.367
R695 B.n13 B.n12 163.367
R696 B.n14 B.n13 163.367
R697 B.n512 B.n14 163.367
R698 B.n512 B.n19 163.367
R699 B.n20 B.n19 163.367
R700 B.n21 B.n20 163.367
R701 B.n517 B.n21 163.367
R702 B.n517 B.n26 163.367
R703 B.n27 B.n26 163.367
R704 B.n28 B.n27 163.367
R705 B.n522 B.n28 163.367
R706 B.n522 B.n33 163.367
R707 B.n34 B.n33 163.367
R708 B.n35 B.n34 163.367
R709 B.n527 B.n35 163.367
R710 B.n527 B.n40 163.367
R711 B.n41 B.n40 163.367
R712 B.n42 B.n41 163.367
R713 B.n532 B.n42 163.367
R714 B.n532 B.n47 163.367
R715 B.n48 B.n47 163.367
R716 B.n49 B.n48 163.367
R717 B.n537 B.n49 163.367
R718 B.n537 B.n54 163.367
R719 B.n55 B.n54 163.367
R720 B.n56 B.n55 163.367
R721 B.n542 B.n56 163.367
R722 B.n542 B.n61 163.367
R723 B.n62 B.n61 163.367
R724 B.n63 B.n62 163.367
R725 B.n719 B.n717 163.367
R726 B.n715 B.n67 163.367
R727 B.n711 B.n709 163.367
R728 B.n707 B.n69 163.367
R729 B.n703 B.n701 163.367
R730 B.n699 B.n71 163.367
R731 B.n695 B.n693 163.367
R732 B.n691 B.n73 163.367
R733 B.n687 B.n685 163.367
R734 B.n683 B.n75 163.367
R735 B.n679 B.n677 163.367
R736 B.n675 B.n77 163.367
R737 B.n671 B.n669 163.367
R738 B.n667 B.n79 163.367
R739 B.n663 B.n661 163.367
R740 B.n659 B.n81 163.367
R741 B.n655 B.n653 163.367
R742 B.n651 B.n83 163.367
R743 B.n647 B.n645 163.367
R744 B.n643 B.n85 163.367
R745 B.n639 B.n637 163.367
R746 B.n635 B.n90 163.367
R747 B.n631 B.n629 163.367
R748 B.n627 B.n92 163.367
R749 B.n622 B.n620 163.367
R750 B.n618 B.n96 163.367
R751 B.n614 B.n612 163.367
R752 B.n610 B.n98 163.367
R753 B.n606 B.n604 163.367
R754 B.n602 B.n100 163.367
R755 B.n598 B.n596 163.367
R756 B.n594 B.n102 163.367
R757 B.n590 B.n588 163.367
R758 B.n586 B.n104 163.367
R759 B.n582 B.n580 163.367
R760 B.n578 B.n106 163.367
R761 B.n574 B.n572 163.367
R762 B.n570 B.n108 163.367
R763 B.n566 B.n564 163.367
R764 B.n562 B.n110 163.367
R765 B.n558 B.n556 163.367
R766 B.n554 B.n112 163.367
R767 B.n550 B.n548 163.367
R768 B.n206 B.t15 103.823
R769 B.n93 B.t20 103.823
R770 B.n200 B.t18 103.808
R771 B.n86 B.t10 103.808
R772 B.n402 B.n178 83.2877
R773 B.n724 B.n64 83.2877
R774 B.n396 B.n179 71.676
R775 B.n394 B.n181 71.676
R776 B.n390 B.n389 71.676
R777 B.n383 B.n183 71.676
R778 B.n382 B.n381 71.676
R779 B.n375 B.n185 71.676
R780 B.n374 B.n373 71.676
R781 B.n367 B.n187 71.676
R782 B.n366 B.n365 71.676
R783 B.n359 B.n189 71.676
R784 B.n358 B.n357 71.676
R785 B.n351 B.n191 71.676
R786 B.n350 B.n349 71.676
R787 B.n343 B.n193 71.676
R788 B.n342 B.n341 71.676
R789 B.n335 B.n195 71.676
R790 B.n334 B.n333 71.676
R791 B.n327 B.n197 71.676
R792 B.n326 B.n325 71.676
R793 B.n318 B.n199 71.676
R794 B.n317 B.n316 71.676
R795 B.n310 B.n203 71.676
R796 B.n309 B.n308 71.676
R797 B.n301 B.n205 71.676
R798 B.n300 B.n299 71.676
R799 B.n293 B.n209 71.676
R800 B.n292 B.n291 71.676
R801 B.n285 B.n211 71.676
R802 B.n284 B.n283 71.676
R803 B.n277 B.n213 71.676
R804 B.n276 B.n275 71.676
R805 B.n269 B.n215 71.676
R806 B.n268 B.n267 71.676
R807 B.n261 B.n217 71.676
R808 B.n260 B.n259 71.676
R809 B.n253 B.n219 71.676
R810 B.n252 B.n251 71.676
R811 B.n245 B.n221 71.676
R812 B.n244 B.n243 71.676
R813 B.n237 B.n223 71.676
R814 B.n236 B.n235 71.676
R815 B.n229 B.n225 71.676
R816 B.n228 B.n227 71.676
R817 B.n718 B.n65 71.676
R818 B.n717 B.n716 71.676
R819 B.n710 B.n67 71.676
R820 B.n709 B.n708 71.676
R821 B.n702 B.n69 71.676
R822 B.n701 B.n700 71.676
R823 B.n694 B.n71 71.676
R824 B.n693 B.n692 71.676
R825 B.n686 B.n73 71.676
R826 B.n685 B.n684 71.676
R827 B.n678 B.n75 71.676
R828 B.n677 B.n676 71.676
R829 B.n670 B.n77 71.676
R830 B.n669 B.n668 71.676
R831 B.n662 B.n79 71.676
R832 B.n661 B.n660 71.676
R833 B.n654 B.n81 71.676
R834 B.n653 B.n652 71.676
R835 B.n646 B.n83 71.676
R836 B.n645 B.n644 71.676
R837 B.n638 B.n85 71.676
R838 B.n637 B.n636 71.676
R839 B.n630 B.n90 71.676
R840 B.n629 B.n628 71.676
R841 B.n621 B.n92 71.676
R842 B.n620 B.n619 71.676
R843 B.n613 B.n96 71.676
R844 B.n612 B.n611 71.676
R845 B.n605 B.n98 71.676
R846 B.n604 B.n603 71.676
R847 B.n597 B.n100 71.676
R848 B.n596 B.n595 71.676
R849 B.n589 B.n102 71.676
R850 B.n588 B.n587 71.676
R851 B.n581 B.n104 71.676
R852 B.n580 B.n579 71.676
R853 B.n573 B.n106 71.676
R854 B.n572 B.n571 71.676
R855 B.n565 B.n108 71.676
R856 B.n564 B.n563 71.676
R857 B.n557 B.n110 71.676
R858 B.n556 B.n555 71.676
R859 B.n549 B.n112 71.676
R860 B.n550 B.n549 71.676
R861 B.n555 B.n554 71.676
R862 B.n558 B.n557 71.676
R863 B.n563 B.n562 71.676
R864 B.n566 B.n565 71.676
R865 B.n571 B.n570 71.676
R866 B.n574 B.n573 71.676
R867 B.n579 B.n578 71.676
R868 B.n582 B.n581 71.676
R869 B.n587 B.n586 71.676
R870 B.n590 B.n589 71.676
R871 B.n595 B.n594 71.676
R872 B.n598 B.n597 71.676
R873 B.n603 B.n602 71.676
R874 B.n606 B.n605 71.676
R875 B.n611 B.n610 71.676
R876 B.n614 B.n613 71.676
R877 B.n619 B.n618 71.676
R878 B.n622 B.n621 71.676
R879 B.n628 B.n627 71.676
R880 B.n631 B.n630 71.676
R881 B.n636 B.n635 71.676
R882 B.n639 B.n638 71.676
R883 B.n644 B.n643 71.676
R884 B.n647 B.n646 71.676
R885 B.n652 B.n651 71.676
R886 B.n655 B.n654 71.676
R887 B.n660 B.n659 71.676
R888 B.n663 B.n662 71.676
R889 B.n668 B.n667 71.676
R890 B.n671 B.n670 71.676
R891 B.n676 B.n675 71.676
R892 B.n679 B.n678 71.676
R893 B.n684 B.n683 71.676
R894 B.n687 B.n686 71.676
R895 B.n692 B.n691 71.676
R896 B.n695 B.n694 71.676
R897 B.n700 B.n699 71.676
R898 B.n703 B.n702 71.676
R899 B.n708 B.n707 71.676
R900 B.n711 B.n710 71.676
R901 B.n716 B.n715 71.676
R902 B.n719 B.n718 71.676
R903 B.n397 B.n396 71.676
R904 B.n391 B.n181 71.676
R905 B.n389 B.n388 71.676
R906 B.n384 B.n383 71.676
R907 B.n381 B.n380 71.676
R908 B.n376 B.n375 71.676
R909 B.n373 B.n372 71.676
R910 B.n368 B.n367 71.676
R911 B.n365 B.n364 71.676
R912 B.n360 B.n359 71.676
R913 B.n357 B.n356 71.676
R914 B.n352 B.n351 71.676
R915 B.n349 B.n348 71.676
R916 B.n344 B.n343 71.676
R917 B.n341 B.n340 71.676
R918 B.n336 B.n335 71.676
R919 B.n333 B.n332 71.676
R920 B.n328 B.n327 71.676
R921 B.n325 B.n324 71.676
R922 B.n319 B.n318 71.676
R923 B.n316 B.n315 71.676
R924 B.n311 B.n310 71.676
R925 B.n308 B.n307 71.676
R926 B.n302 B.n301 71.676
R927 B.n299 B.n298 71.676
R928 B.n294 B.n293 71.676
R929 B.n291 B.n290 71.676
R930 B.n286 B.n285 71.676
R931 B.n283 B.n282 71.676
R932 B.n278 B.n277 71.676
R933 B.n275 B.n274 71.676
R934 B.n270 B.n269 71.676
R935 B.n267 B.n266 71.676
R936 B.n262 B.n261 71.676
R937 B.n259 B.n258 71.676
R938 B.n254 B.n253 71.676
R939 B.n251 B.n250 71.676
R940 B.n246 B.n245 71.676
R941 B.n243 B.n242 71.676
R942 B.n238 B.n237 71.676
R943 B.n235 B.n234 71.676
R944 B.n230 B.n229 71.676
R945 B.n227 B.n177 71.676
R946 B.n207 B.t14 69.6888
R947 B.n94 B.t21 69.6888
R948 B.n201 B.t17 69.675
R949 B.n87 B.t11 69.675
R950 B.n304 B.n207 59.5399
R951 B.n322 B.n201 59.5399
R952 B.n88 B.n87 59.5399
R953 B.n625 B.n94 59.5399
R954 B.n402 B.n174 46.0454
R955 B.n408 B.n174 46.0454
R956 B.n408 B.n169 46.0454
R957 B.n414 B.n169 46.0454
R958 B.n414 B.n170 46.0454
R959 B.n420 B.n162 46.0454
R960 B.n426 B.n162 46.0454
R961 B.n426 B.n158 46.0454
R962 B.n432 B.n158 46.0454
R963 B.n432 B.n154 46.0454
R964 B.n438 B.n154 46.0454
R965 B.n438 B.n150 46.0454
R966 B.n444 B.n150 46.0454
R967 B.n450 B.n146 46.0454
R968 B.n450 B.n142 46.0454
R969 B.n457 B.n142 46.0454
R970 B.n457 B.n456 46.0454
R971 B.n463 B.n135 46.0454
R972 B.n469 B.n135 46.0454
R973 B.n469 B.n131 46.0454
R974 B.n475 B.n131 46.0454
R975 B.n481 B.n127 46.0454
R976 B.n481 B.n122 46.0454
R977 B.n487 B.n122 46.0454
R978 B.n487 B.n123 46.0454
R979 B.n494 B.n115 46.0454
R980 B.n500 B.n115 46.0454
R981 B.n500 B.n4 46.0454
R982 B.n790 B.n4 46.0454
R983 B.n790 B.n789 46.0454
R984 B.n789 B.n788 46.0454
R985 B.n788 B.n8 46.0454
R986 B.n782 B.n8 46.0454
R987 B.n781 B.n780 46.0454
R988 B.n780 B.n15 46.0454
R989 B.n774 B.n15 46.0454
R990 B.n774 B.n773 46.0454
R991 B.n772 B.n22 46.0454
R992 B.n766 B.n22 46.0454
R993 B.n766 B.n765 46.0454
R994 B.n765 B.n764 46.0454
R995 B.n758 B.n32 46.0454
R996 B.n758 B.n757 46.0454
R997 B.n757 B.n756 46.0454
R998 B.n756 B.n36 46.0454
R999 B.n750 B.n749 46.0454
R1000 B.n749 B.n748 46.0454
R1001 B.n748 B.n43 46.0454
R1002 B.n742 B.n43 46.0454
R1003 B.n742 B.n741 46.0454
R1004 B.n741 B.n740 46.0454
R1005 B.n740 B.n50 46.0454
R1006 B.n734 B.n50 46.0454
R1007 B.n733 B.n732 46.0454
R1008 B.n732 B.n57 46.0454
R1009 B.n726 B.n57 46.0454
R1010 B.n726 B.n725 46.0454
R1011 B.n725 B.n724 46.0454
R1012 B.n170 B.t13 41.3055
R1013 B.t9 B.n733 41.3055
R1014 B.n123 B.t0 37.2427
R1015 B.t2 B.n781 37.2427
R1016 B.n207 B.n206 34.1338
R1017 B.n201 B.n200 34.1338
R1018 B.n87 B.n86 34.1338
R1019 B.n94 B.n93 34.1338
R1020 B.t1 B.n146 33.1799
R1021 B.t5 B.n36 33.1799
R1022 B.n722 B.n721 31.0639
R1023 B.n547 B.n546 31.0639
R1024 B.n404 B.n176 31.0639
R1025 B.n400 B.n399 31.0639
R1026 B.n475 B.t3 29.1171
R1027 B.t6 B.n772 29.1171
R1028 B.n463 B.t4 25.0544
R1029 B.n764 B.t7 25.0544
R1030 B.n456 B.t4 20.9916
R1031 B.n32 B.t7 20.9916
R1032 B B.n792 18.0485
R1033 B.t3 B.n127 16.9288
R1034 B.n773 B.t6 16.9288
R1035 B.n444 B.t1 12.866
R1036 B.n750 B.t5 12.866
R1037 B.n721 B.n720 10.6151
R1038 B.n720 B.n66 10.6151
R1039 B.n714 B.n66 10.6151
R1040 B.n714 B.n713 10.6151
R1041 B.n713 B.n712 10.6151
R1042 B.n712 B.n68 10.6151
R1043 B.n706 B.n68 10.6151
R1044 B.n706 B.n705 10.6151
R1045 B.n705 B.n704 10.6151
R1046 B.n704 B.n70 10.6151
R1047 B.n698 B.n70 10.6151
R1048 B.n698 B.n697 10.6151
R1049 B.n697 B.n696 10.6151
R1050 B.n696 B.n72 10.6151
R1051 B.n690 B.n72 10.6151
R1052 B.n690 B.n689 10.6151
R1053 B.n689 B.n688 10.6151
R1054 B.n688 B.n74 10.6151
R1055 B.n682 B.n74 10.6151
R1056 B.n682 B.n681 10.6151
R1057 B.n681 B.n680 10.6151
R1058 B.n680 B.n76 10.6151
R1059 B.n674 B.n76 10.6151
R1060 B.n674 B.n673 10.6151
R1061 B.n673 B.n672 10.6151
R1062 B.n672 B.n78 10.6151
R1063 B.n666 B.n78 10.6151
R1064 B.n666 B.n665 10.6151
R1065 B.n665 B.n664 10.6151
R1066 B.n664 B.n80 10.6151
R1067 B.n658 B.n80 10.6151
R1068 B.n658 B.n657 10.6151
R1069 B.n657 B.n656 10.6151
R1070 B.n656 B.n82 10.6151
R1071 B.n650 B.n82 10.6151
R1072 B.n650 B.n649 10.6151
R1073 B.n649 B.n648 10.6151
R1074 B.n648 B.n84 10.6151
R1075 B.n642 B.n641 10.6151
R1076 B.n641 B.n640 10.6151
R1077 B.n640 B.n89 10.6151
R1078 B.n634 B.n89 10.6151
R1079 B.n634 B.n633 10.6151
R1080 B.n633 B.n632 10.6151
R1081 B.n632 B.n91 10.6151
R1082 B.n626 B.n91 10.6151
R1083 B.n624 B.n623 10.6151
R1084 B.n623 B.n95 10.6151
R1085 B.n617 B.n95 10.6151
R1086 B.n617 B.n616 10.6151
R1087 B.n616 B.n615 10.6151
R1088 B.n615 B.n97 10.6151
R1089 B.n609 B.n97 10.6151
R1090 B.n609 B.n608 10.6151
R1091 B.n608 B.n607 10.6151
R1092 B.n607 B.n99 10.6151
R1093 B.n601 B.n99 10.6151
R1094 B.n601 B.n600 10.6151
R1095 B.n600 B.n599 10.6151
R1096 B.n599 B.n101 10.6151
R1097 B.n593 B.n101 10.6151
R1098 B.n593 B.n592 10.6151
R1099 B.n592 B.n591 10.6151
R1100 B.n591 B.n103 10.6151
R1101 B.n585 B.n103 10.6151
R1102 B.n585 B.n584 10.6151
R1103 B.n584 B.n583 10.6151
R1104 B.n583 B.n105 10.6151
R1105 B.n577 B.n105 10.6151
R1106 B.n577 B.n576 10.6151
R1107 B.n576 B.n575 10.6151
R1108 B.n575 B.n107 10.6151
R1109 B.n569 B.n107 10.6151
R1110 B.n569 B.n568 10.6151
R1111 B.n568 B.n567 10.6151
R1112 B.n567 B.n109 10.6151
R1113 B.n561 B.n109 10.6151
R1114 B.n561 B.n560 10.6151
R1115 B.n560 B.n559 10.6151
R1116 B.n559 B.n111 10.6151
R1117 B.n553 B.n111 10.6151
R1118 B.n553 B.n552 10.6151
R1119 B.n552 B.n551 10.6151
R1120 B.n551 B.n547 10.6151
R1121 B.n405 B.n404 10.6151
R1122 B.n406 B.n405 10.6151
R1123 B.n406 B.n167 10.6151
R1124 B.n416 B.n167 10.6151
R1125 B.n417 B.n416 10.6151
R1126 B.n418 B.n417 10.6151
R1127 B.n418 B.n160 10.6151
R1128 B.n428 B.n160 10.6151
R1129 B.n429 B.n428 10.6151
R1130 B.n430 B.n429 10.6151
R1131 B.n430 B.n152 10.6151
R1132 B.n440 B.n152 10.6151
R1133 B.n441 B.n440 10.6151
R1134 B.n442 B.n441 10.6151
R1135 B.n442 B.n144 10.6151
R1136 B.n452 B.n144 10.6151
R1137 B.n453 B.n452 10.6151
R1138 B.n454 B.n453 10.6151
R1139 B.n454 B.n137 10.6151
R1140 B.n465 B.n137 10.6151
R1141 B.n466 B.n465 10.6151
R1142 B.n467 B.n466 10.6151
R1143 B.n467 B.n129 10.6151
R1144 B.n477 B.n129 10.6151
R1145 B.n478 B.n477 10.6151
R1146 B.n479 B.n478 10.6151
R1147 B.n479 B.n120 10.6151
R1148 B.n489 B.n120 10.6151
R1149 B.n490 B.n489 10.6151
R1150 B.n492 B.n490 10.6151
R1151 B.n492 B.n491 10.6151
R1152 B.n491 B.n113 10.6151
R1153 B.n503 B.n113 10.6151
R1154 B.n504 B.n503 10.6151
R1155 B.n505 B.n504 10.6151
R1156 B.n506 B.n505 10.6151
R1157 B.n508 B.n506 10.6151
R1158 B.n509 B.n508 10.6151
R1159 B.n510 B.n509 10.6151
R1160 B.n511 B.n510 10.6151
R1161 B.n513 B.n511 10.6151
R1162 B.n514 B.n513 10.6151
R1163 B.n515 B.n514 10.6151
R1164 B.n516 B.n515 10.6151
R1165 B.n518 B.n516 10.6151
R1166 B.n519 B.n518 10.6151
R1167 B.n520 B.n519 10.6151
R1168 B.n521 B.n520 10.6151
R1169 B.n523 B.n521 10.6151
R1170 B.n524 B.n523 10.6151
R1171 B.n525 B.n524 10.6151
R1172 B.n526 B.n525 10.6151
R1173 B.n528 B.n526 10.6151
R1174 B.n529 B.n528 10.6151
R1175 B.n530 B.n529 10.6151
R1176 B.n531 B.n530 10.6151
R1177 B.n533 B.n531 10.6151
R1178 B.n534 B.n533 10.6151
R1179 B.n535 B.n534 10.6151
R1180 B.n536 B.n535 10.6151
R1181 B.n538 B.n536 10.6151
R1182 B.n539 B.n538 10.6151
R1183 B.n540 B.n539 10.6151
R1184 B.n541 B.n540 10.6151
R1185 B.n543 B.n541 10.6151
R1186 B.n544 B.n543 10.6151
R1187 B.n545 B.n544 10.6151
R1188 B.n546 B.n545 10.6151
R1189 B.n399 B.n398 10.6151
R1190 B.n398 B.n180 10.6151
R1191 B.n393 B.n180 10.6151
R1192 B.n393 B.n392 10.6151
R1193 B.n392 B.n182 10.6151
R1194 B.n387 B.n182 10.6151
R1195 B.n387 B.n386 10.6151
R1196 B.n386 B.n385 10.6151
R1197 B.n385 B.n184 10.6151
R1198 B.n379 B.n184 10.6151
R1199 B.n379 B.n378 10.6151
R1200 B.n378 B.n377 10.6151
R1201 B.n377 B.n186 10.6151
R1202 B.n371 B.n186 10.6151
R1203 B.n371 B.n370 10.6151
R1204 B.n370 B.n369 10.6151
R1205 B.n369 B.n188 10.6151
R1206 B.n363 B.n188 10.6151
R1207 B.n363 B.n362 10.6151
R1208 B.n362 B.n361 10.6151
R1209 B.n361 B.n190 10.6151
R1210 B.n355 B.n190 10.6151
R1211 B.n355 B.n354 10.6151
R1212 B.n354 B.n353 10.6151
R1213 B.n353 B.n192 10.6151
R1214 B.n347 B.n192 10.6151
R1215 B.n347 B.n346 10.6151
R1216 B.n346 B.n345 10.6151
R1217 B.n345 B.n194 10.6151
R1218 B.n339 B.n194 10.6151
R1219 B.n339 B.n338 10.6151
R1220 B.n338 B.n337 10.6151
R1221 B.n337 B.n196 10.6151
R1222 B.n331 B.n196 10.6151
R1223 B.n331 B.n330 10.6151
R1224 B.n330 B.n329 10.6151
R1225 B.n329 B.n198 10.6151
R1226 B.n323 B.n198 10.6151
R1227 B.n321 B.n320 10.6151
R1228 B.n320 B.n202 10.6151
R1229 B.n314 B.n202 10.6151
R1230 B.n314 B.n313 10.6151
R1231 B.n313 B.n312 10.6151
R1232 B.n312 B.n204 10.6151
R1233 B.n306 B.n204 10.6151
R1234 B.n306 B.n305 10.6151
R1235 B.n303 B.n208 10.6151
R1236 B.n297 B.n208 10.6151
R1237 B.n297 B.n296 10.6151
R1238 B.n296 B.n295 10.6151
R1239 B.n295 B.n210 10.6151
R1240 B.n289 B.n210 10.6151
R1241 B.n289 B.n288 10.6151
R1242 B.n288 B.n287 10.6151
R1243 B.n287 B.n212 10.6151
R1244 B.n281 B.n212 10.6151
R1245 B.n281 B.n280 10.6151
R1246 B.n280 B.n279 10.6151
R1247 B.n279 B.n214 10.6151
R1248 B.n273 B.n214 10.6151
R1249 B.n273 B.n272 10.6151
R1250 B.n272 B.n271 10.6151
R1251 B.n271 B.n216 10.6151
R1252 B.n265 B.n216 10.6151
R1253 B.n265 B.n264 10.6151
R1254 B.n264 B.n263 10.6151
R1255 B.n263 B.n218 10.6151
R1256 B.n257 B.n218 10.6151
R1257 B.n257 B.n256 10.6151
R1258 B.n256 B.n255 10.6151
R1259 B.n255 B.n220 10.6151
R1260 B.n249 B.n220 10.6151
R1261 B.n249 B.n248 10.6151
R1262 B.n248 B.n247 10.6151
R1263 B.n247 B.n222 10.6151
R1264 B.n241 B.n222 10.6151
R1265 B.n241 B.n240 10.6151
R1266 B.n240 B.n239 10.6151
R1267 B.n239 B.n224 10.6151
R1268 B.n233 B.n224 10.6151
R1269 B.n233 B.n232 10.6151
R1270 B.n232 B.n231 10.6151
R1271 B.n231 B.n226 10.6151
R1272 B.n226 B.n176 10.6151
R1273 B.n400 B.n172 10.6151
R1274 B.n410 B.n172 10.6151
R1275 B.n411 B.n410 10.6151
R1276 B.n412 B.n411 10.6151
R1277 B.n412 B.n164 10.6151
R1278 B.n422 B.n164 10.6151
R1279 B.n423 B.n422 10.6151
R1280 B.n424 B.n423 10.6151
R1281 B.n424 B.n156 10.6151
R1282 B.n434 B.n156 10.6151
R1283 B.n435 B.n434 10.6151
R1284 B.n436 B.n435 10.6151
R1285 B.n436 B.n148 10.6151
R1286 B.n446 B.n148 10.6151
R1287 B.n447 B.n446 10.6151
R1288 B.n448 B.n447 10.6151
R1289 B.n448 B.n140 10.6151
R1290 B.n459 B.n140 10.6151
R1291 B.n460 B.n459 10.6151
R1292 B.n461 B.n460 10.6151
R1293 B.n461 B.n133 10.6151
R1294 B.n471 B.n133 10.6151
R1295 B.n472 B.n471 10.6151
R1296 B.n473 B.n472 10.6151
R1297 B.n473 B.n125 10.6151
R1298 B.n483 B.n125 10.6151
R1299 B.n484 B.n483 10.6151
R1300 B.n485 B.n484 10.6151
R1301 B.n485 B.n117 10.6151
R1302 B.n496 B.n117 10.6151
R1303 B.n497 B.n496 10.6151
R1304 B.n498 B.n497 10.6151
R1305 B.n498 B.n0 10.6151
R1306 B.n786 B.n1 10.6151
R1307 B.n786 B.n785 10.6151
R1308 B.n785 B.n784 10.6151
R1309 B.n784 B.n10 10.6151
R1310 B.n778 B.n10 10.6151
R1311 B.n778 B.n777 10.6151
R1312 B.n777 B.n776 10.6151
R1313 B.n776 B.n17 10.6151
R1314 B.n770 B.n17 10.6151
R1315 B.n770 B.n769 10.6151
R1316 B.n769 B.n768 10.6151
R1317 B.n768 B.n24 10.6151
R1318 B.n762 B.n24 10.6151
R1319 B.n762 B.n761 10.6151
R1320 B.n761 B.n760 10.6151
R1321 B.n760 B.n30 10.6151
R1322 B.n754 B.n30 10.6151
R1323 B.n754 B.n753 10.6151
R1324 B.n753 B.n752 10.6151
R1325 B.n752 B.n38 10.6151
R1326 B.n746 B.n38 10.6151
R1327 B.n746 B.n745 10.6151
R1328 B.n745 B.n744 10.6151
R1329 B.n744 B.n45 10.6151
R1330 B.n738 B.n45 10.6151
R1331 B.n738 B.n737 10.6151
R1332 B.n737 B.n736 10.6151
R1333 B.n736 B.n52 10.6151
R1334 B.n730 B.n52 10.6151
R1335 B.n730 B.n729 10.6151
R1336 B.n729 B.n728 10.6151
R1337 B.n728 B.n59 10.6151
R1338 B.n722 B.n59 10.6151
R1339 B.n494 B.t0 8.80321
R1340 B.n782 B.t2 8.80321
R1341 B.n642 B.n88 6.5566
R1342 B.n626 B.n625 6.5566
R1343 B.n322 B.n321 6.5566
R1344 B.n305 B.n304 6.5566
R1345 B.n420 B.t13 4.74042
R1346 B.n734 B.t9 4.74042
R1347 B.n88 B.n84 4.05904
R1348 B.n625 B.n624 4.05904
R1349 B.n323 B.n322 4.05904
R1350 B.n304 B.n303 4.05904
R1351 B.n792 B.n0 2.81026
R1352 B.n792 B.n1 2.81026
R1353 VN.n5 VN.t2 216.931
R1354 VN.n24 VN.t5 216.931
R1355 VN.n4 VN.t1 184.88
R1356 VN.n10 VN.t0 184.88
R1357 VN.n17 VN.t7 184.88
R1358 VN.n23 VN.t6 184.88
R1359 VN.n29 VN.t3 184.88
R1360 VN.n36 VN.t4 184.88
R1361 VN.n18 VN.n17 178.917
R1362 VN.n37 VN.n36 178.917
R1363 VN.n35 VN.n19 161.3
R1364 VN.n34 VN.n33 161.3
R1365 VN.n32 VN.n20 161.3
R1366 VN.n31 VN.n30 161.3
R1367 VN.n28 VN.n21 161.3
R1368 VN.n27 VN.n26 161.3
R1369 VN.n25 VN.n22 161.3
R1370 VN.n16 VN.n0 161.3
R1371 VN.n15 VN.n14 161.3
R1372 VN.n13 VN.n1 161.3
R1373 VN.n12 VN.n11 161.3
R1374 VN.n9 VN.n2 161.3
R1375 VN.n8 VN.n7 161.3
R1376 VN.n6 VN.n3 161.3
R1377 VN.n15 VN.n1 56.5193
R1378 VN.n34 VN.n20 56.5193
R1379 VN.n5 VN.n4 47.4662
R1380 VN.n24 VN.n23 47.4662
R1381 VN VN.n37 44.8812
R1382 VN.n8 VN.n3 40.4934
R1383 VN.n9 VN.n8 40.4934
R1384 VN.n27 VN.n22 40.4934
R1385 VN.n28 VN.n27 40.4934
R1386 VN.n11 VN.n1 24.4675
R1387 VN.n16 VN.n15 24.4675
R1388 VN.n30 VN.n20 24.4675
R1389 VN.n35 VN.n34 24.4675
R1390 VN.n4 VN.n3 18.5954
R1391 VN.n10 VN.n9 18.5954
R1392 VN.n23 VN.n22 18.5954
R1393 VN.n29 VN.n28 18.5954
R1394 VN.n25 VN.n24 18.0957
R1395 VN.n6 VN.n5 18.0957
R1396 VN.n17 VN.n16 6.85126
R1397 VN.n36 VN.n35 6.85126
R1398 VN.n11 VN.n10 5.87258
R1399 VN.n30 VN.n29 5.87258
R1400 VN.n37 VN.n19 0.189894
R1401 VN.n33 VN.n19 0.189894
R1402 VN.n33 VN.n32 0.189894
R1403 VN.n32 VN.n31 0.189894
R1404 VN.n31 VN.n21 0.189894
R1405 VN.n26 VN.n21 0.189894
R1406 VN.n26 VN.n25 0.189894
R1407 VN.n7 VN.n6 0.189894
R1408 VN.n7 VN.n2 0.189894
R1409 VN.n12 VN.n2 0.189894
R1410 VN.n13 VN.n12 0.189894
R1411 VN.n14 VN.n13 0.189894
R1412 VN.n14 VN.n0 0.189894
R1413 VN.n18 VN.n0 0.189894
R1414 VN VN.n18 0.0516364
R1415 VDD2.n2 VDD2.n1 61.5546
R1416 VDD2.n2 VDD2.n0 61.5546
R1417 VDD2 VDD2.n5 61.5518
R1418 VDD2.n4 VDD2.n3 60.8516
R1419 VDD2.n4 VDD2.n2 39.9998
R1420 VDD2.n5 VDD2.t1 1.80542
R1421 VDD2.n5 VDD2.t2 1.80542
R1422 VDD2.n3 VDD2.t6 1.80542
R1423 VDD2.n3 VDD2.t0 1.80542
R1424 VDD2.n1 VDD2.t7 1.80542
R1425 VDD2.n1 VDD2.t3 1.80542
R1426 VDD2.n0 VDD2.t5 1.80542
R1427 VDD2.n0 VDD2.t4 1.80542
R1428 VDD2 VDD2.n4 0.81731
R1429 VTAIL.n11 VTAIL.t3 45.9776
R1430 VTAIL.n10 VTAIL.t9 45.9776
R1431 VTAIL.n7 VTAIL.t10 45.9776
R1432 VTAIL.n15 VTAIL.t7 45.9775
R1433 VTAIL.n2 VTAIL.t12 45.9775
R1434 VTAIL.n3 VTAIL.t0 45.9775
R1435 VTAIL.n6 VTAIL.t1 45.9775
R1436 VTAIL.n14 VTAIL.t15 45.9775
R1437 VTAIL.n13 VTAIL.n12 44.1728
R1438 VTAIL.n9 VTAIL.n8 44.1728
R1439 VTAIL.n1 VTAIL.n0 44.1725
R1440 VTAIL.n5 VTAIL.n4 44.1725
R1441 VTAIL.n15 VTAIL.n14 23.341
R1442 VTAIL.n7 VTAIL.n6 23.341
R1443 VTAIL.n0 VTAIL.t13 1.80542
R1444 VTAIL.n0 VTAIL.t14 1.80542
R1445 VTAIL.n4 VTAIL.t6 1.80542
R1446 VTAIL.n4 VTAIL.t2 1.80542
R1447 VTAIL.n12 VTAIL.t4 1.80542
R1448 VTAIL.n12 VTAIL.t5 1.80542
R1449 VTAIL.n8 VTAIL.t11 1.80542
R1450 VTAIL.n8 VTAIL.t8 1.80542
R1451 VTAIL.n9 VTAIL.n7 1.51774
R1452 VTAIL.n10 VTAIL.n9 1.51774
R1453 VTAIL.n13 VTAIL.n11 1.51774
R1454 VTAIL.n14 VTAIL.n13 1.51774
R1455 VTAIL.n6 VTAIL.n5 1.51774
R1456 VTAIL.n5 VTAIL.n3 1.51774
R1457 VTAIL.n2 VTAIL.n1 1.51774
R1458 VTAIL VTAIL.n15 1.45955
R1459 VTAIL.n11 VTAIL.n10 0.470328
R1460 VTAIL.n3 VTAIL.n2 0.470328
R1461 VTAIL VTAIL.n1 0.0586897
R1462 VP.n11 VP.t0 216.931
R1463 VP.n25 VP.t1 184.88
R1464 VP.n31 VP.t5 184.88
R1465 VP.n38 VP.t2 184.88
R1466 VP.n45 VP.t4 184.88
R1467 VP.n23 VP.t7 184.88
R1468 VP.n16 VP.t6 184.88
R1469 VP.n10 VP.t3 184.88
R1470 VP.n26 VP.n25 178.917
R1471 VP.n46 VP.n45 178.917
R1472 VP.n24 VP.n23 178.917
R1473 VP.n12 VP.n9 161.3
R1474 VP.n14 VP.n13 161.3
R1475 VP.n15 VP.n8 161.3
R1476 VP.n18 VP.n17 161.3
R1477 VP.n19 VP.n7 161.3
R1478 VP.n21 VP.n20 161.3
R1479 VP.n22 VP.n6 161.3
R1480 VP.n44 VP.n0 161.3
R1481 VP.n43 VP.n42 161.3
R1482 VP.n41 VP.n1 161.3
R1483 VP.n40 VP.n39 161.3
R1484 VP.n37 VP.n2 161.3
R1485 VP.n36 VP.n35 161.3
R1486 VP.n34 VP.n3 161.3
R1487 VP.n33 VP.n32 161.3
R1488 VP.n30 VP.n4 161.3
R1489 VP.n29 VP.n28 161.3
R1490 VP.n27 VP.n5 161.3
R1491 VP.n30 VP.n29 56.5193
R1492 VP.n43 VP.n1 56.5193
R1493 VP.n21 VP.n7 56.5193
R1494 VP.n11 VP.n10 47.4662
R1495 VP.n26 VP.n24 44.5005
R1496 VP.n36 VP.n3 40.4934
R1497 VP.n37 VP.n36 40.4934
R1498 VP.n15 VP.n14 40.4934
R1499 VP.n14 VP.n9 40.4934
R1500 VP.n29 VP.n5 24.4675
R1501 VP.n32 VP.n30 24.4675
R1502 VP.n39 VP.n1 24.4675
R1503 VP.n44 VP.n43 24.4675
R1504 VP.n22 VP.n21 24.4675
R1505 VP.n17 VP.n7 24.4675
R1506 VP.n31 VP.n3 18.5954
R1507 VP.n38 VP.n37 18.5954
R1508 VP.n16 VP.n15 18.5954
R1509 VP.n10 VP.n9 18.5954
R1510 VP.n12 VP.n11 18.0957
R1511 VP.n25 VP.n5 6.85126
R1512 VP.n45 VP.n44 6.85126
R1513 VP.n23 VP.n22 6.85126
R1514 VP.n32 VP.n31 5.87258
R1515 VP.n39 VP.n38 5.87258
R1516 VP.n17 VP.n16 5.87258
R1517 VP.n13 VP.n12 0.189894
R1518 VP.n13 VP.n8 0.189894
R1519 VP.n18 VP.n8 0.189894
R1520 VP.n19 VP.n18 0.189894
R1521 VP.n20 VP.n19 0.189894
R1522 VP.n20 VP.n6 0.189894
R1523 VP.n24 VP.n6 0.189894
R1524 VP.n27 VP.n26 0.189894
R1525 VP.n28 VP.n27 0.189894
R1526 VP.n28 VP.n4 0.189894
R1527 VP.n33 VP.n4 0.189894
R1528 VP.n34 VP.n33 0.189894
R1529 VP.n35 VP.n34 0.189894
R1530 VP.n35 VP.n2 0.189894
R1531 VP.n40 VP.n2 0.189894
R1532 VP.n41 VP.n40 0.189894
R1533 VP.n42 VP.n41 0.189894
R1534 VP.n42 VP.n0 0.189894
R1535 VP.n46 VP.n0 0.189894
R1536 VP VP.n46 0.0516364
R1537 VDD1 VDD1.n0 61.6684
R1538 VDD1.n3 VDD1.n2 61.5546
R1539 VDD1.n3 VDD1.n1 61.5546
R1540 VDD1.n5 VDD1.n4 60.8514
R1541 VDD1.n5 VDD1.n3 40.5828
R1542 VDD1.n4 VDD1.t1 1.80542
R1543 VDD1.n4 VDD1.t0 1.80542
R1544 VDD1.n0 VDD1.t7 1.80542
R1545 VDD1.n0 VDD1.t4 1.80542
R1546 VDD1.n2 VDD1.t5 1.80542
R1547 VDD1.n2 VDD1.t3 1.80542
R1548 VDD1.n1 VDD1.t6 1.80542
R1549 VDD1.n1 VDD1.t2 1.80542
R1550 VDD1 VDD1.n5 0.700931
C0 VDD1 VDD2 1.19381f
C1 VN VP 6.04388f
C2 VTAIL VN 6.90882f
C3 VTAIL VP 6.92292f
C4 VN VDD2 6.8396f
C5 VDD1 VN 0.149679f
C6 VP VDD2 0.395237f
C7 VDD1 VP 7.08435f
C8 VTAIL VDD2 8.121119f
C9 VDD1 VTAIL 8.07455f
C10 VDD2 B 4.116332f
C11 VDD1 B 4.431564f
C12 VTAIL B 8.986009f
C13 VN B 11.01837f
C14 VP B 9.424911f
C15 VDD1.t7 B 0.219169f
C16 VDD1.t4 B 0.219169f
C17 VDD1.n0 B 1.94587f
C18 VDD1.t6 B 0.219169f
C19 VDD1.t2 B 0.219169f
C20 VDD1.n1 B 1.94503f
C21 VDD1.t5 B 0.219169f
C22 VDD1.t3 B 0.219169f
C23 VDD1.n2 B 1.94503f
C24 VDD1.n3 B 2.61885f
C25 VDD1.t1 B 0.219169f
C26 VDD1.t0 B 0.219169f
C27 VDD1.n4 B 1.94044f
C28 VDD1.n5 B 2.52363f
C29 VP.n0 B 0.032299f
C30 VP.t4 B 1.37681f
C31 VP.n1 B 0.048051f
C32 VP.n2 B 0.032299f
C33 VP.t2 B 1.37681f
C34 VP.n3 B 0.057061f
C35 VP.n4 B 0.032299f
C36 VP.n5 B 0.038799f
C37 VP.n6 B 0.032299f
C38 VP.t7 B 1.37681f
C39 VP.n7 B 0.048051f
C40 VP.n8 B 0.032299f
C41 VP.t6 B 1.37681f
C42 VP.n9 B 0.057061f
C43 VP.t0 B 1.46869f
C44 VP.t3 B 1.37681f
C45 VP.n10 B 0.568746f
C46 VP.n11 B 0.577509f
C47 VP.n12 B 0.200975f
C48 VP.n13 B 0.032299f
C49 VP.n14 B 0.026111f
C50 VP.n15 B 0.057061f
C51 VP.n16 B 0.503037f
C52 VP.n17 B 0.03761f
C53 VP.n18 B 0.032299f
C54 VP.n19 B 0.032299f
C55 VP.n20 B 0.032299f
C56 VP.n21 B 0.046251f
C57 VP.n22 B 0.038799f
C58 VP.n23 B 0.561059f
C59 VP.n24 B 1.47178f
C60 VP.t1 B 1.37681f
C61 VP.n25 B 0.561059f
C62 VP.n26 B 1.49787f
C63 VP.n27 B 0.032299f
C64 VP.n28 B 0.032299f
C65 VP.n29 B 0.046251f
C66 VP.n30 B 0.048051f
C67 VP.t5 B 1.37681f
C68 VP.n31 B 0.503037f
C69 VP.n32 B 0.03761f
C70 VP.n33 B 0.032299f
C71 VP.n34 B 0.032299f
C72 VP.n35 B 0.032299f
C73 VP.n36 B 0.026111f
C74 VP.n37 B 0.057061f
C75 VP.n38 B 0.503037f
C76 VP.n39 B 0.03761f
C77 VP.n40 B 0.032299f
C78 VP.n41 B 0.032299f
C79 VP.n42 B 0.032299f
C80 VP.n43 B 0.046251f
C81 VP.n44 B 0.038799f
C82 VP.n45 B 0.561059f
C83 VP.n46 B 0.031367f
C84 VTAIL.t13 B 0.168589f
C85 VTAIL.t14 B 0.168589f
C86 VTAIL.n0 B 1.43323f
C87 VTAIL.n1 B 0.292697f
C88 VTAIL.t12 B 1.82532f
C89 VTAIL.n2 B 0.386192f
C90 VTAIL.t0 B 1.82532f
C91 VTAIL.n3 B 0.386192f
C92 VTAIL.t6 B 0.168589f
C93 VTAIL.t2 B 0.168589f
C94 VTAIL.n4 B 1.43323f
C95 VTAIL.n5 B 0.384128f
C96 VTAIL.t1 B 1.82532f
C97 VTAIL.n6 B 1.30862f
C98 VTAIL.t10 B 1.82534f
C99 VTAIL.n7 B 1.30861f
C100 VTAIL.t11 B 0.168589f
C101 VTAIL.t8 B 0.168589f
C102 VTAIL.n8 B 1.43324f
C103 VTAIL.n9 B 0.384124f
C104 VTAIL.t9 B 1.82534f
C105 VTAIL.n10 B 0.38618f
C106 VTAIL.t3 B 1.82534f
C107 VTAIL.n11 B 0.38618f
C108 VTAIL.t4 B 0.168589f
C109 VTAIL.t5 B 0.168589f
C110 VTAIL.n12 B 1.43324f
C111 VTAIL.n13 B 0.384124f
C112 VTAIL.t15 B 1.82532f
C113 VTAIL.n14 B 1.30862f
C114 VTAIL.t7 B 1.82532f
C115 VTAIL.n15 B 1.30497f
C116 VDD2.t5 B 0.216171f
C117 VDD2.t4 B 0.216171f
C118 VDD2.n0 B 1.91842f
C119 VDD2.t7 B 0.216171f
C120 VDD2.t3 B 0.216171f
C121 VDD2.n1 B 1.91842f
C122 VDD2.n2 B 2.53031f
C123 VDD2.t6 B 0.216171f
C124 VDD2.t0 B 0.216171f
C125 VDD2.n3 B 1.9139f
C126 VDD2.n4 B 2.45907f
C127 VDD2.t1 B 0.216171f
C128 VDD2.t2 B 0.216171f
C129 VDD2.n5 B 1.91839f
C130 VN.n0 B 0.031743f
C131 VN.t7 B 1.35308f
C132 VN.n1 B 0.047223f
C133 VN.n2 B 0.031743f
C134 VN.t0 B 1.35308f
C135 VN.n3 B 0.056078f
C136 VN.t2 B 1.44339f
C137 VN.t1 B 1.35308f
C138 VN.n4 B 0.558946f
C139 VN.n5 B 0.567558f
C140 VN.n6 B 0.197512f
C141 VN.n7 B 0.031743f
C142 VN.n8 B 0.025661f
C143 VN.n9 B 0.056078f
C144 VN.n10 B 0.494369f
C145 VN.n11 B 0.036962f
C146 VN.n12 B 0.031743f
C147 VN.n13 B 0.031743f
C148 VN.n14 B 0.031743f
C149 VN.n15 B 0.045454f
C150 VN.n16 B 0.038131f
C151 VN.n17 B 0.551391f
C152 VN.n18 B 0.030827f
C153 VN.n19 B 0.031743f
C154 VN.t4 B 1.35308f
C155 VN.n20 B 0.047223f
C156 VN.n21 B 0.031743f
C157 VN.t3 B 1.35308f
C158 VN.n22 B 0.056078f
C159 VN.t5 B 1.44339f
C160 VN.t6 B 1.35308f
C161 VN.n23 B 0.558946f
C162 VN.n24 B 0.567558f
C163 VN.n25 B 0.197512f
C164 VN.n26 B 0.031743f
C165 VN.n27 B 0.025661f
C166 VN.n28 B 0.056078f
C167 VN.n29 B 0.494369f
C168 VN.n30 B 0.036962f
C169 VN.n31 B 0.031743f
C170 VN.n32 B 0.031743f
C171 VN.n33 B 0.031743f
C172 VN.n34 B 0.045454f
C173 VN.n35 B 0.038131f
C174 VN.n36 B 0.551391f
C175 VN.n37 B 1.46718f
.ends

