* NGSPICE file created from diff_pair_sample_0878.ext - technology: sky130A

.subckt diff_pair_sample_0878 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.38
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.38
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.38
X3 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=3.0264 ps=16.3 w=7.76 l=2.38
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=3.0264 ps=16.3 w=7.76 l=2.38
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=3.0264 ps=16.3 w=7.76 l=2.38
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.38
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0264 pd=16.3 as=3.0264 ps=16.3 w=7.76 l=2.38
R0 B.n544 B.n543 585
R1 B.n218 B.n81 585
R2 B.n217 B.n216 585
R3 B.n215 B.n214 585
R4 B.n213 B.n212 585
R5 B.n211 B.n210 585
R6 B.n209 B.n208 585
R7 B.n207 B.n206 585
R8 B.n205 B.n204 585
R9 B.n203 B.n202 585
R10 B.n201 B.n200 585
R11 B.n199 B.n198 585
R12 B.n197 B.n196 585
R13 B.n195 B.n194 585
R14 B.n193 B.n192 585
R15 B.n191 B.n190 585
R16 B.n189 B.n188 585
R17 B.n187 B.n186 585
R18 B.n185 B.n184 585
R19 B.n183 B.n182 585
R20 B.n181 B.n180 585
R21 B.n179 B.n178 585
R22 B.n177 B.n176 585
R23 B.n175 B.n174 585
R24 B.n173 B.n172 585
R25 B.n171 B.n170 585
R26 B.n169 B.n168 585
R27 B.n167 B.n166 585
R28 B.n165 B.n164 585
R29 B.n162 B.n161 585
R30 B.n160 B.n159 585
R31 B.n158 B.n157 585
R32 B.n156 B.n155 585
R33 B.n154 B.n153 585
R34 B.n152 B.n151 585
R35 B.n150 B.n149 585
R36 B.n148 B.n147 585
R37 B.n146 B.n145 585
R38 B.n144 B.n143 585
R39 B.n141 B.n140 585
R40 B.n139 B.n138 585
R41 B.n137 B.n136 585
R42 B.n135 B.n134 585
R43 B.n133 B.n132 585
R44 B.n131 B.n130 585
R45 B.n129 B.n128 585
R46 B.n127 B.n126 585
R47 B.n125 B.n124 585
R48 B.n123 B.n122 585
R49 B.n121 B.n120 585
R50 B.n119 B.n118 585
R51 B.n117 B.n116 585
R52 B.n115 B.n114 585
R53 B.n113 B.n112 585
R54 B.n111 B.n110 585
R55 B.n109 B.n108 585
R56 B.n107 B.n106 585
R57 B.n105 B.n104 585
R58 B.n103 B.n102 585
R59 B.n101 B.n100 585
R60 B.n99 B.n98 585
R61 B.n97 B.n96 585
R62 B.n95 B.n94 585
R63 B.n93 B.n92 585
R64 B.n91 B.n90 585
R65 B.n89 B.n88 585
R66 B.n87 B.n86 585
R67 B.n46 B.n45 585
R68 B.n542 B.n47 585
R69 B.n547 B.n47 585
R70 B.n541 B.n540 585
R71 B.n540 B.n43 585
R72 B.n539 B.n42 585
R73 B.n553 B.n42 585
R74 B.n538 B.n41 585
R75 B.n554 B.n41 585
R76 B.n537 B.n40 585
R77 B.n555 B.n40 585
R78 B.n536 B.n535 585
R79 B.n535 B.n36 585
R80 B.n534 B.n35 585
R81 B.n561 B.n35 585
R82 B.n533 B.n34 585
R83 B.n562 B.n34 585
R84 B.n532 B.n33 585
R85 B.n563 B.n33 585
R86 B.n531 B.n530 585
R87 B.n530 B.n29 585
R88 B.n529 B.n28 585
R89 B.n569 B.n28 585
R90 B.n528 B.n27 585
R91 B.n570 B.n27 585
R92 B.n527 B.n26 585
R93 B.n571 B.n26 585
R94 B.n526 B.n525 585
R95 B.n525 B.n22 585
R96 B.n524 B.n21 585
R97 B.n577 B.n21 585
R98 B.n523 B.n20 585
R99 B.n578 B.n20 585
R100 B.n522 B.n19 585
R101 B.n579 B.n19 585
R102 B.n521 B.n520 585
R103 B.n520 B.n15 585
R104 B.n519 B.n14 585
R105 B.n585 B.n14 585
R106 B.n518 B.n13 585
R107 B.n586 B.n13 585
R108 B.n517 B.n12 585
R109 B.n587 B.n12 585
R110 B.n516 B.n515 585
R111 B.n515 B.n8 585
R112 B.n514 B.n7 585
R113 B.n593 B.n7 585
R114 B.n513 B.n6 585
R115 B.n594 B.n6 585
R116 B.n512 B.n5 585
R117 B.n595 B.n5 585
R118 B.n511 B.n510 585
R119 B.n510 B.n4 585
R120 B.n509 B.n219 585
R121 B.n509 B.n508 585
R122 B.n499 B.n220 585
R123 B.n221 B.n220 585
R124 B.n501 B.n500 585
R125 B.n502 B.n501 585
R126 B.n498 B.n226 585
R127 B.n226 B.n225 585
R128 B.n497 B.n496 585
R129 B.n496 B.n495 585
R130 B.n228 B.n227 585
R131 B.n229 B.n228 585
R132 B.n488 B.n487 585
R133 B.n489 B.n488 585
R134 B.n486 B.n234 585
R135 B.n234 B.n233 585
R136 B.n485 B.n484 585
R137 B.n484 B.n483 585
R138 B.n236 B.n235 585
R139 B.n237 B.n236 585
R140 B.n476 B.n475 585
R141 B.n477 B.n476 585
R142 B.n474 B.n242 585
R143 B.n242 B.n241 585
R144 B.n473 B.n472 585
R145 B.n472 B.n471 585
R146 B.n244 B.n243 585
R147 B.n245 B.n244 585
R148 B.n464 B.n463 585
R149 B.n465 B.n464 585
R150 B.n462 B.n249 585
R151 B.n253 B.n249 585
R152 B.n461 B.n460 585
R153 B.n460 B.n459 585
R154 B.n251 B.n250 585
R155 B.n252 B.n251 585
R156 B.n452 B.n451 585
R157 B.n453 B.n452 585
R158 B.n450 B.n258 585
R159 B.n258 B.n257 585
R160 B.n449 B.n448 585
R161 B.n448 B.n447 585
R162 B.n260 B.n259 585
R163 B.n261 B.n260 585
R164 B.n440 B.n439 585
R165 B.n441 B.n440 585
R166 B.n264 B.n263 585
R167 B.n307 B.n306 585
R168 B.n308 B.n304 585
R169 B.n304 B.n265 585
R170 B.n310 B.n309 585
R171 B.n312 B.n303 585
R172 B.n315 B.n314 585
R173 B.n316 B.n302 585
R174 B.n318 B.n317 585
R175 B.n320 B.n301 585
R176 B.n323 B.n322 585
R177 B.n324 B.n300 585
R178 B.n326 B.n325 585
R179 B.n328 B.n299 585
R180 B.n331 B.n330 585
R181 B.n332 B.n298 585
R182 B.n334 B.n333 585
R183 B.n336 B.n297 585
R184 B.n339 B.n338 585
R185 B.n340 B.n296 585
R186 B.n342 B.n341 585
R187 B.n344 B.n295 585
R188 B.n347 B.n346 585
R189 B.n348 B.n294 585
R190 B.n350 B.n349 585
R191 B.n352 B.n293 585
R192 B.n355 B.n354 585
R193 B.n356 B.n292 585
R194 B.n358 B.n357 585
R195 B.n360 B.n291 585
R196 B.n363 B.n362 585
R197 B.n364 B.n287 585
R198 B.n366 B.n365 585
R199 B.n368 B.n286 585
R200 B.n371 B.n370 585
R201 B.n372 B.n285 585
R202 B.n374 B.n373 585
R203 B.n376 B.n284 585
R204 B.n379 B.n378 585
R205 B.n380 B.n281 585
R206 B.n383 B.n382 585
R207 B.n385 B.n280 585
R208 B.n388 B.n387 585
R209 B.n389 B.n279 585
R210 B.n391 B.n390 585
R211 B.n393 B.n278 585
R212 B.n396 B.n395 585
R213 B.n397 B.n277 585
R214 B.n399 B.n398 585
R215 B.n401 B.n276 585
R216 B.n404 B.n403 585
R217 B.n405 B.n275 585
R218 B.n407 B.n406 585
R219 B.n409 B.n274 585
R220 B.n412 B.n411 585
R221 B.n413 B.n273 585
R222 B.n415 B.n414 585
R223 B.n417 B.n272 585
R224 B.n420 B.n419 585
R225 B.n421 B.n271 585
R226 B.n423 B.n422 585
R227 B.n425 B.n270 585
R228 B.n428 B.n427 585
R229 B.n429 B.n269 585
R230 B.n431 B.n430 585
R231 B.n433 B.n268 585
R232 B.n434 B.n267 585
R233 B.n437 B.n436 585
R234 B.n438 B.n266 585
R235 B.n266 B.n265 585
R236 B.n443 B.n442 585
R237 B.n442 B.n441 585
R238 B.n444 B.n262 585
R239 B.n262 B.n261 585
R240 B.n446 B.n445 585
R241 B.n447 B.n446 585
R242 B.n256 B.n255 585
R243 B.n257 B.n256 585
R244 B.n455 B.n454 585
R245 B.n454 B.n453 585
R246 B.n456 B.n254 585
R247 B.n254 B.n252 585
R248 B.n458 B.n457 585
R249 B.n459 B.n458 585
R250 B.n248 B.n247 585
R251 B.n253 B.n248 585
R252 B.n467 B.n466 585
R253 B.n466 B.n465 585
R254 B.n468 B.n246 585
R255 B.n246 B.n245 585
R256 B.n470 B.n469 585
R257 B.n471 B.n470 585
R258 B.n240 B.n239 585
R259 B.n241 B.n240 585
R260 B.n479 B.n478 585
R261 B.n478 B.n477 585
R262 B.n480 B.n238 585
R263 B.n238 B.n237 585
R264 B.n482 B.n481 585
R265 B.n483 B.n482 585
R266 B.n232 B.n231 585
R267 B.n233 B.n232 585
R268 B.n491 B.n490 585
R269 B.n490 B.n489 585
R270 B.n492 B.n230 585
R271 B.n230 B.n229 585
R272 B.n494 B.n493 585
R273 B.n495 B.n494 585
R274 B.n224 B.n223 585
R275 B.n225 B.n224 585
R276 B.n504 B.n503 585
R277 B.n503 B.n502 585
R278 B.n505 B.n222 585
R279 B.n222 B.n221 585
R280 B.n507 B.n506 585
R281 B.n508 B.n507 585
R282 B.n2 B.n0 585
R283 B.n4 B.n2 585
R284 B.n3 B.n1 585
R285 B.n594 B.n3 585
R286 B.n592 B.n591 585
R287 B.n593 B.n592 585
R288 B.n590 B.n9 585
R289 B.n9 B.n8 585
R290 B.n589 B.n588 585
R291 B.n588 B.n587 585
R292 B.n11 B.n10 585
R293 B.n586 B.n11 585
R294 B.n584 B.n583 585
R295 B.n585 B.n584 585
R296 B.n582 B.n16 585
R297 B.n16 B.n15 585
R298 B.n581 B.n580 585
R299 B.n580 B.n579 585
R300 B.n18 B.n17 585
R301 B.n578 B.n18 585
R302 B.n576 B.n575 585
R303 B.n577 B.n576 585
R304 B.n574 B.n23 585
R305 B.n23 B.n22 585
R306 B.n573 B.n572 585
R307 B.n572 B.n571 585
R308 B.n25 B.n24 585
R309 B.n570 B.n25 585
R310 B.n568 B.n567 585
R311 B.n569 B.n568 585
R312 B.n566 B.n30 585
R313 B.n30 B.n29 585
R314 B.n565 B.n564 585
R315 B.n564 B.n563 585
R316 B.n32 B.n31 585
R317 B.n562 B.n32 585
R318 B.n560 B.n559 585
R319 B.n561 B.n560 585
R320 B.n558 B.n37 585
R321 B.n37 B.n36 585
R322 B.n557 B.n556 585
R323 B.n556 B.n555 585
R324 B.n39 B.n38 585
R325 B.n554 B.n39 585
R326 B.n552 B.n551 585
R327 B.n553 B.n552 585
R328 B.n550 B.n44 585
R329 B.n44 B.n43 585
R330 B.n549 B.n548 585
R331 B.n548 B.n547 585
R332 B.n597 B.n596 585
R333 B.n596 B.n595 585
R334 B.n442 B.n264 497.305
R335 B.n548 B.n46 497.305
R336 B.n440 B.n266 497.305
R337 B.n544 B.n47 497.305
R338 B.n282 B.t2 286.267
R339 B.n288 B.t6 286.267
R340 B.n84 B.t13 286.267
R341 B.n82 B.t9 286.267
R342 B.n546 B.n545 256.663
R343 B.n546 B.n80 256.663
R344 B.n546 B.n79 256.663
R345 B.n546 B.n78 256.663
R346 B.n546 B.n77 256.663
R347 B.n546 B.n76 256.663
R348 B.n546 B.n75 256.663
R349 B.n546 B.n74 256.663
R350 B.n546 B.n73 256.663
R351 B.n546 B.n72 256.663
R352 B.n546 B.n71 256.663
R353 B.n546 B.n70 256.663
R354 B.n546 B.n69 256.663
R355 B.n546 B.n68 256.663
R356 B.n546 B.n67 256.663
R357 B.n546 B.n66 256.663
R358 B.n546 B.n65 256.663
R359 B.n546 B.n64 256.663
R360 B.n546 B.n63 256.663
R361 B.n546 B.n62 256.663
R362 B.n546 B.n61 256.663
R363 B.n546 B.n60 256.663
R364 B.n546 B.n59 256.663
R365 B.n546 B.n58 256.663
R366 B.n546 B.n57 256.663
R367 B.n546 B.n56 256.663
R368 B.n546 B.n55 256.663
R369 B.n546 B.n54 256.663
R370 B.n546 B.n53 256.663
R371 B.n546 B.n52 256.663
R372 B.n546 B.n51 256.663
R373 B.n546 B.n50 256.663
R374 B.n546 B.n49 256.663
R375 B.n546 B.n48 256.663
R376 B.n305 B.n265 256.663
R377 B.n311 B.n265 256.663
R378 B.n313 B.n265 256.663
R379 B.n319 B.n265 256.663
R380 B.n321 B.n265 256.663
R381 B.n327 B.n265 256.663
R382 B.n329 B.n265 256.663
R383 B.n335 B.n265 256.663
R384 B.n337 B.n265 256.663
R385 B.n343 B.n265 256.663
R386 B.n345 B.n265 256.663
R387 B.n351 B.n265 256.663
R388 B.n353 B.n265 256.663
R389 B.n359 B.n265 256.663
R390 B.n361 B.n265 256.663
R391 B.n367 B.n265 256.663
R392 B.n369 B.n265 256.663
R393 B.n375 B.n265 256.663
R394 B.n377 B.n265 256.663
R395 B.n384 B.n265 256.663
R396 B.n386 B.n265 256.663
R397 B.n392 B.n265 256.663
R398 B.n394 B.n265 256.663
R399 B.n400 B.n265 256.663
R400 B.n402 B.n265 256.663
R401 B.n408 B.n265 256.663
R402 B.n410 B.n265 256.663
R403 B.n416 B.n265 256.663
R404 B.n418 B.n265 256.663
R405 B.n424 B.n265 256.663
R406 B.n426 B.n265 256.663
R407 B.n432 B.n265 256.663
R408 B.n435 B.n265 256.663
R409 B.n442 B.n262 163.367
R410 B.n446 B.n262 163.367
R411 B.n446 B.n256 163.367
R412 B.n454 B.n256 163.367
R413 B.n454 B.n254 163.367
R414 B.n458 B.n254 163.367
R415 B.n458 B.n248 163.367
R416 B.n466 B.n248 163.367
R417 B.n466 B.n246 163.367
R418 B.n470 B.n246 163.367
R419 B.n470 B.n240 163.367
R420 B.n478 B.n240 163.367
R421 B.n478 B.n238 163.367
R422 B.n482 B.n238 163.367
R423 B.n482 B.n232 163.367
R424 B.n490 B.n232 163.367
R425 B.n490 B.n230 163.367
R426 B.n494 B.n230 163.367
R427 B.n494 B.n224 163.367
R428 B.n503 B.n224 163.367
R429 B.n503 B.n222 163.367
R430 B.n507 B.n222 163.367
R431 B.n507 B.n2 163.367
R432 B.n596 B.n2 163.367
R433 B.n596 B.n3 163.367
R434 B.n592 B.n3 163.367
R435 B.n592 B.n9 163.367
R436 B.n588 B.n9 163.367
R437 B.n588 B.n11 163.367
R438 B.n584 B.n11 163.367
R439 B.n584 B.n16 163.367
R440 B.n580 B.n16 163.367
R441 B.n580 B.n18 163.367
R442 B.n576 B.n18 163.367
R443 B.n576 B.n23 163.367
R444 B.n572 B.n23 163.367
R445 B.n572 B.n25 163.367
R446 B.n568 B.n25 163.367
R447 B.n568 B.n30 163.367
R448 B.n564 B.n30 163.367
R449 B.n564 B.n32 163.367
R450 B.n560 B.n32 163.367
R451 B.n560 B.n37 163.367
R452 B.n556 B.n37 163.367
R453 B.n556 B.n39 163.367
R454 B.n552 B.n39 163.367
R455 B.n552 B.n44 163.367
R456 B.n548 B.n44 163.367
R457 B.n306 B.n304 163.367
R458 B.n310 B.n304 163.367
R459 B.n314 B.n312 163.367
R460 B.n318 B.n302 163.367
R461 B.n322 B.n320 163.367
R462 B.n326 B.n300 163.367
R463 B.n330 B.n328 163.367
R464 B.n334 B.n298 163.367
R465 B.n338 B.n336 163.367
R466 B.n342 B.n296 163.367
R467 B.n346 B.n344 163.367
R468 B.n350 B.n294 163.367
R469 B.n354 B.n352 163.367
R470 B.n358 B.n292 163.367
R471 B.n362 B.n360 163.367
R472 B.n366 B.n287 163.367
R473 B.n370 B.n368 163.367
R474 B.n374 B.n285 163.367
R475 B.n378 B.n376 163.367
R476 B.n383 B.n281 163.367
R477 B.n387 B.n385 163.367
R478 B.n391 B.n279 163.367
R479 B.n395 B.n393 163.367
R480 B.n399 B.n277 163.367
R481 B.n403 B.n401 163.367
R482 B.n407 B.n275 163.367
R483 B.n411 B.n409 163.367
R484 B.n415 B.n273 163.367
R485 B.n419 B.n417 163.367
R486 B.n423 B.n271 163.367
R487 B.n427 B.n425 163.367
R488 B.n431 B.n269 163.367
R489 B.n434 B.n433 163.367
R490 B.n436 B.n266 163.367
R491 B.n440 B.n260 163.367
R492 B.n448 B.n260 163.367
R493 B.n448 B.n258 163.367
R494 B.n452 B.n258 163.367
R495 B.n452 B.n251 163.367
R496 B.n460 B.n251 163.367
R497 B.n460 B.n249 163.367
R498 B.n464 B.n249 163.367
R499 B.n464 B.n244 163.367
R500 B.n472 B.n244 163.367
R501 B.n472 B.n242 163.367
R502 B.n476 B.n242 163.367
R503 B.n476 B.n236 163.367
R504 B.n484 B.n236 163.367
R505 B.n484 B.n234 163.367
R506 B.n488 B.n234 163.367
R507 B.n488 B.n228 163.367
R508 B.n496 B.n228 163.367
R509 B.n496 B.n226 163.367
R510 B.n501 B.n226 163.367
R511 B.n501 B.n220 163.367
R512 B.n509 B.n220 163.367
R513 B.n510 B.n509 163.367
R514 B.n510 B.n5 163.367
R515 B.n6 B.n5 163.367
R516 B.n7 B.n6 163.367
R517 B.n515 B.n7 163.367
R518 B.n515 B.n12 163.367
R519 B.n13 B.n12 163.367
R520 B.n14 B.n13 163.367
R521 B.n520 B.n14 163.367
R522 B.n520 B.n19 163.367
R523 B.n20 B.n19 163.367
R524 B.n21 B.n20 163.367
R525 B.n525 B.n21 163.367
R526 B.n525 B.n26 163.367
R527 B.n27 B.n26 163.367
R528 B.n28 B.n27 163.367
R529 B.n530 B.n28 163.367
R530 B.n530 B.n33 163.367
R531 B.n34 B.n33 163.367
R532 B.n35 B.n34 163.367
R533 B.n535 B.n35 163.367
R534 B.n535 B.n40 163.367
R535 B.n41 B.n40 163.367
R536 B.n42 B.n41 163.367
R537 B.n540 B.n42 163.367
R538 B.n540 B.n47 163.367
R539 B.n88 B.n87 163.367
R540 B.n92 B.n91 163.367
R541 B.n96 B.n95 163.367
R542 B.n100 B.n99 163.367
R543 B.n104 B.n103 163.367
R544 B.n108 B.n107 163.367
R545 B.n112 B.n111 163.367
R546 B.n116 B.n115 163.367
R547 B.n120 B.n119 163.367
R548 B.n124 B.n123 163.367
R549 B.n128 B.n127 163.367
R550 B.n132 B.n131 163.367
R551 B.n136 B.n135 163.367
R552 B.n140 B.n139 163.367
R553 B.n145 B.n144 163.367
R554 B.n149 B.n148 163.367
R555 B.n153 B.n152 163.367
R556 B.n157 B.n156 163.367
R557 B.n161 B.n160 163.367
R558 B.n166 B.n165 163.367
R559 B.n170 B.n169 163.367
R560 B.n174 B.n173 163.367
R561 B.n178 B.n177 163.367
R562 B.n182 B.n181 163.367
R563 B.n186 B.n185 163.367
R564 B.n190 B.n189 163.367
R565 B.n194 B.n193 163.367
R566 B.n198 B.n197 163.367
R567 B.n202 B.n201 163.367
R568 B.n206 B.n205 163.367
R569 B.n210 B.n209 163.367
R570 B.n214 B.n213 163.367
R571 B.n216 B.n81 163.367
R572 B.n282 B.t5 126.674
R573 B.n82 B.t11 126.674
R574 B.n288 B.t8 126.665
R575 B.n84 B.t14 126.665
R576 B.n441 B.n265 107.174
R577 B.n547 B.n546 107.174
R578 B.n283 B.t4 74.1166
R579 B.n83 B.t12 74.1166
R580 B.n289 B.t7 74.1079
R581 B.n85 B.t15 74.1079
R582 B.n305 B.n264 71.676
R583 B.n311 B.n310 71.676
R584 B.n314 B.n313 71.676
R585 B.n319 B.n318 71.676
R586 B.n322 B.n321 71.676
R587 B.n327 B.n326 71.676
R588 B.n330 B.n329 71.676
R589 B.n335 B.n334 71.676
R590 B.n338 B.n337 71.676
R591 B.n343 B.n342 71.676
R592 B.n346 B.n345 71.676
R593 B.n351 B.n350 71.676
R594 B.n354 B.n353 71.676
R595 B.n359 B.n358 71.676
R596 B.n362 B.n361 71.676
R597 B.n367 B.n366 71.676
R598 B.n370 B.n369 71.676
R599 B.n375 B.n374 71.676
R600 B.n378 B.n377 71.676
R601 B.n384 B.n383 71.676
R602 B.n387 B.n386 71.676
R603 B.n392 B.n391 71.676
R604 B.n395 B.n394 71.676
R605 B.n400 B.n399 71.676
R606 B.n403 B.n402 71.676
R607 B.n408 B.n407 71.676
R608 B.n411 B.n410 71.676
R609 B.n416 B.n415 71.676
R610 B.n419 B.n418 71.676
R611 B.n424 B.n423 71.676
R612 B.n427 B.n426 71.676
R613 B.n432 B.n431 71.676
R614 B.n435 B.n434 71.676
R615 B.n48 B.n46 71.676
R616 B.n88 B.n49 71.676
R617 B.n92 B.n50 71.676
R618 B.n96 B.n51 71.676
R619 B.n100 B.n52 71.676
R620 B.n104 B.n53 71.676
R621 B.n108 B.n54 71.676
R622 B.n112 B.n55 71.676
R623 B.n116 B.n56 71.676
R624 B.n120 B.n57 71.676
R625 B.n124 B.n58 71.676
R626 B.n128 B.n59 71.676
R627 B.n132 B.n60 71.676
R628 B.n136 B.n61 71.676
R629 B.n140 B.n62 71.676
R630 B.n145 B.n63 71.676
R631 B.n149 B.n64 71.676
R632 B.n153 B.n65 71.676
R633 B.n157 B.n66 71.676
R634 B.n161 B.n67 71.676
R635 B.n166 B.n68 71.676
R636 B.n170 B.n69 71.676
R637 B.n174 B.n70 71.676
R638 B.n178 B.n71 71.676
R639 B.n182 B.n72 71.676
R640 B.n186 B.n73 71.676
R641 B.n190 B.n74 71.676
R642 B.n194 B.n75 71.676
R643 B.n198 B.n76 71.676
R644 B.n202 B.n77 71.676
R645 B.n206 B.n78 71.676
R646 B.n210 B.n79 71.676
R647 B.n214 B.n80 71.676
R648 B.n545 B.n81 71.676
R649 B.n545 B.n544 71.676
R650 B.n216 B.n80 71.676
R651 B.n213 B.n79 71.676
R652 B.n209 B.n78 71.676
R653 B.n205 B.n77 71.676
R654 B.n201 B.n76 71.676
R655 B.n197 B.n75 71.676
R656 B.n193 B.n74 71.676
R657 B.n189 B.n73 71.676
R658 B.n185 B.n72 71.676
R659 B.n181 B.n71 71.676
R660 B.n177 B.n70 71.676
R661 B.n173 B.n69 71.676
R662 B.n169 B.n68 71.676
R663 B.n165 B.n67 71.676
R664 B.n160 B.n66 71.676
R665 B.n156 B.n65 71.676
R666 B.n152 B.n64 71.676
R667 B.n148 B.n63 71.676
R668 B.n144 B.n62 71.676
R669 B.n139 B.n61 71.676
R670 B.n135 B.n60 71.676
R671 B.n131 B.n59 71.676
R672 B.n127 B.n58 71.676
R673 B.n123 B.n57 71.676
R674 B.n119 B.n56 71.676
R675 B.n115 B.n55 71.676
R676 B.n111 B.n54 71.676
R677 B.n107 B.n53 71.676
R678 B.n103 B.n52 71.676
R679 B.n99 B.n51 71.676
R680 B.n95 B.n50 71.676
R681 B.n91 B.n49 71.676
R682 B.n87 B.n48 71.676
R683 B.n306 B.n305 71.676
R684 B.n312 B.n311 71.676
R685 B.n313 B.n302 71.676
R686 B.n320 B.n319 71.676
R687 B.n321 B.n300 71.676
R688 B.n328 B.n327 71.676
R689 B.n329 B.n298 71.676
R690 B.n336 B.n335 71.676
R691 B.n337 B.n296 71.676
R692 B.n344 B.n343 71.676
R693 B.n345 B.n294 71.676
R694 B.n352 B.n351 71.676
R695 B.n353 B.n292 71.676
R696 B.n360 B.n359 71.676
R697 B.n361 B.n287 71.676
R698 B.n368 B.n367 71.676
R699 B.n369 B.n285 71.676
R700 B.n376 B.n375 71.676
R701 B.n377 B.n281 71.676
R702 B.n385 B.n384 71.676
R703 B.n386 B.n279 71.676
R704 B.n393 B.n392 71.676
R705 B.n394 B.n277 71.676
R706 B.n401 B.n400 71.676
R707 B.n402 B.n275 71.676
R708 B.n409 B.n408 71.676
R709 B.n410 B.n273 71.676
R710 B.n417 B.n416 71.676
R711 B.n418 B.n271 71.676
R712 B.n425 B.n424 71.676
R713 B.n426 B.n269 71.676
R714 B.n433 B.n432 71.676
R715 B.n436 B.n435 71.676
R716 B.n381 B.n283 59.5399
R717 B.n290 B.n289 59.5399
R718 B.n142 B.n85 59.5399
R719 B.n163 B.n83 59.5399
R720 B.n441 B.n261 57.3845
R721 B.n447 B.n261 57.3845
R722 B.n447 B.n257 57.3845
R723 B.n453 B.n257 57.3845
R724 B.n453 B.n252 57.3845
R725 B.n459 B.n252 57.3845
R726 B.n459 B.n253 57.3845
R727 B.n465 B.n245 57.3845
R728 B.n471 B.n245 57.3845
R729 B.n471 B.n241 57.3845
R730 B.n477 B.n241 57.3845
R731 B.n477 B.n237 57.3845
R732 B.n483 B.n237 57.3845
R733 B.n483 B.n233 57.3845
R734 B.n489 B.n233 57.3845
R735 B.n489 B.n229 57.3845
R736 B.n495 B.n229 57.3845
R737 B.n502 B.n225 57.3845
R738 B.n502 B.n221 57.3845
R739 B.n508 B.n221 57.3845
R740 B.n508 B.n4 57.3845
R741 B.n595 B.n4 57.3845
R742 B.n595 B.n594 57.3845
R743 B.n594 B.n593 57.3845
R744 B.n593 B.n8 57.3845
R745 B.n587 B.n8 57.3845
R746 B.n587 B.n586 57.3845
R747 B.n585 B.n15 57.3845
R748 B.n579 B.n15 57.3845
R749 B.n579 B.n578 57.3845
R750 B.n578 B.n577 57.3845
R751 B.n577 B.n22 57.3845
R752 B.n571 B.n22 57.3845
R753 B.n571 B.n570 57.3845
R754 B.n570 B.n569 57.3845
R755 B.n569 B.n29 57.3845
R756 B.n563 B.n29 57.3845
R757 B.n562 B.n561 57.3845
R758 B.n561 B.n36 57.3845
R759 B.n555 B.n36 57.3845
R760 B.n555 B.n554 57.3845
R761 B.n554 B.n553 57.3845
R762 B.n553 B.n43 57.3845
R763 B.n547 B.n43 57.3845
R764 B.n283 B.n282 52.5581
R765 B.n289 B.n288 52.5581
R766 B.n85 B.n84 52.5581
R767 B.n83 B.n82 52.5581
R768 B.n465 B.t3 43.8824
R769 B.n563 B.t10 43.8824
R770 B.t0 B.n225 33.7558
R771 B.n586 B.t1 33.7558
R772 B.n549 B.n45 32.3127
R773 B.n543 B.n542 32.3127
R774 B.n439 B.n438 32.3127
R775 B.n443 B.n263 32.3127
R776 B.n495 B.t0 23.6292
R777 B.t1 B.n585 23.6292
R778 B B.n597 18.0485
R779 B.n253 B.t3 13.5026
R780 B.t10 B.n562 13.5026
R781 B.n86 B.n45 10.6151
R782 B.n89 B.n86 10.6151
R783 B.n90 B.n89 10.6151
R784 B.n93 B.n90 10.6151
R785 B.n94 B.n93 10.6151
R786 B.n97 B.n94 10.6151
R787 B.n98 B.n97 10.6151
R788 B.n101 B.n98 10.6151
R789 B.n102 B.n101 10.6151
R790 B.n105 B.n102 10.6151
R791 B.n106 B.n105 10.6151
R792 B.n109 B.n106 10.6151
R793 B.n110 B.n109 10.6151
R794 B.n113 B.n110 10.6151
R795 B.n114 B.n113 10.6151
R796 B.n117 B.n114 10.6151
R797 B.n118 B.n117 10.6151
R798 B.n121 B.n118 10.6151
R799 B.n122 B.n121 10.6151
R800 B.n125 B.n122 10.6151
R801 B.n126 B.n125 10.6151
R802 B.n129 B.n126 10.6151
R803 B.n130 B.n129 10.6151
R804 B.n133 B.n130 10.6151
R805 B.n134 B.n133 10.6151
R806 B.n137 B.n134 10.6151
R807 B.n138 B.n137 10.6151
R808 B.n141 B.n138 10.6151
R809 B.n146 B.n143 10.6151
R810 B.n147 B.n146 10.6151
R811 B.n150 B.n147 10.6151
R812 B.n151 B.n150 10.6151
R813 B.n154 B.n151 10.6151
R814 B.n155 B.n154 10.6151
R815 B.n158 B.n155 10.6151
R816 B.n159 B.n158 10.6151
R817 B.n162 B.n159 10.6151
R818 B.n167 B.n164 10.6151
R819 B.n168 B.n167 10.6151
R820 B.n171 B.n168 10.6151
R821 B.n172 B.n171 10.6151
R822 B.n175 B.n172 10.6151
R823 B.n176 B.n175 10.6151
R824 B.n179 B.n176 10.6151
R825 B.n180 B.n179 10.6151
R826 B.n183 B.n180 10.6151
R827 B.n184 B.n183 10.6151
R828 B.n187 B.n184 10.6151
R829 B.n188 B.n187 10.6151
R830 B.n191 B.n188 10.6151
R831 B.n192 B.n191 10.6151
R832 B.n195 B.n192 10.6151
R833 B.n196 B.n195 10.6151
R834 B.n199 B.n196 10.6151
R835 B.n200 B.n199 10.6151
R836 B.n203 B.n200 10.6151
R837 B.n204 B.n203 10.6151
R838 B.n207 B.n204 10.6151
R839 B.n208 B.n207 10.6151
R840 B.n211 B.n208 10.6151
R841 B.n212 B.n211 10.6151
R842 B.n215 B.n212 10.6151
R843 B.n217 B.n215 10.6151
R844 B.n218 B.n217 10.6151
R845 B.n543 B.n218 10.6151
R846 B.n439 B.n259 10.6151
R847 B.n449 B.n259 10.6151
R848 B.n450 B.n449 10.6151
R849 B.n451 B.n450 10.6151
R850 B.n451 B.n250 10.6151
R851 B.n461 B.n250 10.6151
R852 B.n462 B.n461 10.6151
R853 B.n463 B.n462 10.6151
R854 B.n463 B.n243 10.6151
R855 B.n473 B.n243 10.6151
R856 B.n474 B.n473 10.6151
R857 B.n475 B.n474 10.6151
R858 B.n475 B.n235 10.6151
R859 B.n485 B.n235 10.6151
R860 B.n486 B.n485 10.6151
R861 B.n487 B.n486 10.6151
R862 B.n487 B.n227 10.6151
R863 B.n497 B.n227 10.6151
R864 B.n498 B.n497 10.6151
R865 B.n500 B.n498 10.6151
R866 B.n500 B.n499 10.6151
R867 B.n499 B.n219 10.6151
R868 B.n511 B.n219 10.6151
R869 B.n512 B.n511 10.6151
R870 B.n513 B.n512 10.6151
R871 B.n514 B.n513 10.6151
R872 B.n516 B.n514 10.6151
R873 B.n517 B.n516 10.6151
R874 B.n518 B.n517 10.6151
R875 B.n519 B.n518 10.6151
R876 B.n521 B.n519 10.6151
R877 B.n522 B.n521 10.6151
R878 B.n523 B.n522 10.6151
R879 B.n524 B.n523 10.6151
R880 B.n526 B.n524 10.6151
R881 B.n527 B.n526 10.6151
R882 B.n528 B.n527 10.6151
R883 B.n529 B.n528 10.6151
R884 B.n531 B.n529 10.6151
R885 B.n532 B.n531 10.6151
R886 B.n533 B.n532 10.6151
R887 B.n534 B.n533 10.6151
R888 B.n536 B.n534 10.6151
R889 B.n537 B.n536 10.6151
R890 B.n538 B.n537 10.6151
R891 B.n539 B.n538 10.6151
R892 B.n541 B.n539 10.6151
R893 B.n542 B.n541 10.6151
R894 B.n307 B.n263 10.6151
R895 B.n308 B.n307 10.6151
R896 B.n309 B.n308 10.6151
R897 B.n309 B.n303 10.6151
R898 B.n315 B.n303 10.6151
R899 B.n316 B.n315 10.6151
R900 B.n317 B.n316 10.6151
R901 B.n317 B.n301 10.6151
R902 B.n323 B.n301 10.6151
R903 B.n324 B.n323 10.6151
R904 B.n325 B.n324 10.6151
R905 B.n325 B.n299 10.6151
R906 B.n331 B.n299 10.6151
R907 B.n332 B.n331 10.6151
R908 B.n333 B.n332 10.6151
R909 B.n333 B.n297 10.6151
R910 B.n339 B.n297 10.6151
R911 B.n340 B.n339 10.6151
R912 B.n341 B.n340 10.6151
R913 B.n341 B.n295 10.6151
R914 B.n347 B.n295 10.6151
R915 B.n348 B.n347 10.6151
R916 B.n349 B.n348 10.6151
R917 B.n349 B.n293 10.6151
R918 B.n355 B.n293 10.6151
R919 B.n356 B.n355 10.6151
R920 B.n357 B.n356 10.6151
R921 B.n357 B.n291 10.6151
R922 B.n364 B.n363 10.6151
R923 B.n365 B.n364 10.6151
R924 B.n365 B.n286 10.6151
R925 B.n371 B.n286 10.6151
R926 B.n372 B.n371 10.6151
R927 B.n373 B.n372 10.6151
R928 B.n373 B.n284 10.6151
R929 B.n379 B.n284 10.6151
R930 B.n380 B.n379 10.6151
R931 B.n382 B.n280 10.6151
R932 B.n388 B.n280 10.6151
R933 B.n389 B.n388 10.6151
R934 B.n390 B.n389 10.6151
R935 B.n390 B.n278 10.6151
R936 B.n396 B.n278 10.6151
R937 B.n397 B.n396 10.6151
R938 B.n398 B.n397 10.6151
R939 B.n398 B.n276 10.6151
R940 B.n404 B.n276 10.6151
R941 B.n405 B.n404 10.6151
R942 B.n406 B.n405 10.6151
R943 B.n406 B.n274 10.6151
R944 B.n412 B.n274 10.6151
R945 B.n413 B.n412 10.6151
R946 B.n414 B.n413 10.6151
R947 B.n414 B.n272 10.6151
R948 B.n420 B.n272 10.6151
R949 B.n421 B.n420 10.6151
R950 B.n422 B.n421 10.6151
R951 B.n422 B.n270 10.6151
R952 B.n428 B.n270 10.6151
R953 B.n429 B.n428 10.6151
R954 B.n430 B.n429 10.6151
R955 B.n430 B.n268 10.6151
R956 B.n268 B.n267 10.6151
R957 B.n437 B.n267 10.6151
R958 B.n438 B.n437 10.6151
R959 B.n444 B.n443 10.6151
R960 B.n445 B.n444 10.6151
R961 B.n445 B.n255 10.6151
R962 B.n455 B.n255 10.6151
R963 B.n456 B.n455 10.6151
R964 B.n457 B.n456 10.6151
R965 B.n457 B.n247 10.6151
R966 B.n467 B.n247 10.6151
R967 B.n468 B.n467 10.6151
R968 B.n469 B.n468 10.6151
R969 B.n469 B.n239 10.6151
R970 B.n479 B.n239 10.6151
R971 B.n480 B.n479 10.6151
R972 B.n481 B.n480 10.6151
R973 B.n481 B.n231 10.6151
R974 B.n491 B.n231 10.6151
R975 B.n492 B.n491 10.6151
R976 B.n493 B.n492 10.6151
R977 B.n493 B.n223 10.6151
R978 B.n504 B.n223 10.6151
R979 B.n505 B.n504 10.6151
R980 B.n506 B.n505 10.6151
R981 B.n506 B.n0 10.6151
R982 B.n591 B.n1 10.6151
R983 B.n591 B.n590 10.6151
R984 B.n590 B.n589 10.6151
R985 B.n589 B.n10 10.6151
R986 B.n583 B.n10 10.6151
R987 B.n583 B.n582 10.6151
R988 B.n582 B.n581 10.6151
R989 B.n581 B.n17 10.6151
R990 B.n575 B.n17 10.6151
R991 B.n575 B.n574 10.6151
R992 B.n574 B.n573 10.6151
R993 B.n573 B.n24 10.6151
R994 B.n567 B.n24 10.6151
R995 B.n567 B.n566 10.6151
R996 B.n566 B.n565 10.6151
R997 B.n565 B.n31 10.6151
R998 B.n559 B.n31 10.6151
R999 B.n559 B.n558 10.6151
R1000 B.n558 B.n557 10.6151
R1001 B.n557 B.n38 10.6151
R1002 B.n551 B.n38 10.6151
R1003 B.n551 B.n550 10.6151
R1004 B.n550 B.n549 10.6151
R1005 B.n142 B.n141 9.36635
R1006 B.n164 B.n163 9.36635
R1007 B.n291 B.n290 9.36635
R1008 B.n382 B.n381 9.36635
R1009 B.n597 B.n0 2.81026
R1010 B.n597 B.n1 2.81026
R1011 B.n143 B.n142 1.24928
R1012 B.n163 B.n162 1.24928
R1013 B.n363 B.n290 1.24928
R1014 B.n381 B.n380 1.24928
R1015 VN VN.t1 168.751
R1016 VN VN.t0 128.13
R1017 VTAIL.n2 VTAIL.t1 49.9296
R1018 VTAIL.n1 VTAIL.t2 49.9296
R1019 VTAIL.n3 VTAIL.t3 49.9295
R1020 VTAIL.n0 VTAIL.t0 49.9295
R1021 VTAIL.n1 VTAIL.n0 23.7289
R1022 VTAIL.n3 VTAIL.n2 21.3927
R1023 VTAIL.n2 VTAIL.n1 1.63843
R1024 VTAIL VTAIL.n0 1.11257
R1025 VTAIL VTAIL.n3 0.526362
R1026 VDD2.n0 VDD2.t1 101.629
R1027 VDD2.n0 VDD2.t0 66.6084
R1028 VDD2 VDD2.n0 0.642741
R1029 VP.n0 VP.t1 168.655
R1030 VP.n0 VP.t0 127.793
R1031 VP VP.n0 0.336784
R1032 VDD1 VDD1.t1 102.739
R1033 VDD1 VDD1.t0 67.2506
C0 VDD1 VP 2.03311f
C1 VTAIL VP 1.71088f
C2 VDD1 VTAIL 3.90162f
C3 VDD2 VP 0.323808f
C4 VDD1 VDD2 0.64776f
C5 VN VP 4.56435f
C6 VDD1 VN 0.148355f
C7 VTAIL VDD2 3.95158f
C8 VTAIL VN 1.69664f
C9 VN VDD2 1.85952f
C10 VDD2 B 3.555877f
C11 VDD1 B 6.34558f
C12 VTAIL B 5.533646f
C13 VN B 7.9181f
C14 VP B 5.829003f
C15 VDD1.t0 B 1.38613f
C16 VDD1.t1 B 1.83764f
C17 VP.t1 B 2.04862f
C18 VP.t0 B 1.65244f
C19 VP.n0 B 2.83748f
C20 VDD2.t1 B 1.2403f
C21 VDD2.t0 B 0.950286f
C22 VDD2.n0 B 1.72612f
C23 VTAIL.t0 B 0.977694f
C24 VTAIL.n0 B 1.02924f
C25 VTAIL.t2 B 0.9777f
C26 VTAIL.n1 B 1.05539f
C27 VTAIL.t1 B 0.977699f
C28 VTAIL.n2 B 0.93921f
C29 VTAIL.t3 B 0.977694f
C30 VTAIL.n3 B 0.883911f
C31 VN.t0 B 1.14583f
C32 VN.t1 B 1.42159f
.ends

