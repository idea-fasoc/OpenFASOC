* NGSPICE file created from diff_pair_sample_1450.ext - technology: sky130A

.subckt diff_pair_sample_1450 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=3.9351 ps=20.96 w=10.09 l=0.86
X1 B.t11 B.t9 B.t10 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=0 ps=0 w=10.09 l=0.86
X2 B.t8 B.t6 B.t7 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=0 ps=0 w=10.09 l=0.86
X3 B.t5 B.t3 B.t4 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=0 ps=0 w=10.09 l=0.86
X4 VDD1.t0 VP.t1 VTAIL.t2 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=3.9351 ps=20.96 w=10.09 l=0.86
X5 B.t2 B.t0 B.t1 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=0 ps=0 w=10.09 l=0.86
X6 VDD2.t1 VN.t0 VTAIL.t0 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=3.9351 ps=20.96 w=10.09 l=0.86
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n1446_n2990# sky130_fd_pr__pfet_01v8 ad=3.9351 pd=20.96 as=3.9351 ps=20.96 w=10.09 l=0.86
R0 VP.n0 VP.t0 528.624
R1 VP.n0 VP.t1 490.014
R2 VP VP.n0 0.0516364
R3 VTAIL.n210 VTAIL.n162 756.745
R4 VTAIL.n48 VTAIL.n0 756.745
R5 VTAIL.n156 VTAIL.n108 756.745
R6 VTAIL.n102 VTAIL.n54 756.745
R7 VTAIL.n178 VTAIL.n177 585
R8 VTAIL.n183 VTAIL.n182 585
R9 VTAIL.n185 VTAIL.n184 585
R10 VTAIL.n174 VTAIL.n173 585
R11 VTAIL.n191 VTAIL.n190 585
R12 VTAIL.n193 VTAIL.n192 585
R13 VTAIL.n170 VTAIL.n169 585
R14 VTAIL.n200 VTAIL.n199 585
R15 VTAIL.n201 VTAIL.n168 585
R16 VTAIL.n203 VTAIL.n202 585
R17 VTAIL.n166 VTAIL.n165 585
R18 VTAIL.n209 VTAIL.n208 585
R19 VTAIL.n211 VTAIL.n210 585
R20 VTAIL.n16 VTAIL.n15 585
R21 VTAIL.n21 VTAIL.n20 585
R22 VTAIL.n23 VTAIL.n22 585
R23 VTAIL.n12 VTAIL.n11 585
R24 VTAIL.n29 VTAIL.n28 585
R25 VTAIL.n31 VTAIL.n30 585
R26 VTAIL.n8 VTAIL.n7 585
R27 VTAIL.n38 VTAIL.n37 585
R28 VTAIL.n39 VTAIL.n6 585
R29 VTAIL.n41 VTAIL.n40 585
R30 VTAIL.n4 VTAIL.n3 585
R31 VTAIL.n47 VTAIL.n46 585
R32 VTAIL.n49 VTAIL.n48 585
R33 VTAIL.n157 VTAIL.n156 585
R34 VTAIL.n155 VTAIL.n154 585
R35 VTAIL.n112 VTAIL.n111 585
R36 VTAIL.n149 VTAIL.n148 585
R37 VTAIL.n147 VTAIL.n114 585
R38 VTAIL.n146 VTAIL.n145 585
R39 VTAIL.n117 VTAIL.n115 585
R40 VTAIL.n140 VTAIL.n139 585
R41 VTAIL.n138 VTAIL.n137 585
R42 VTAIL.n121 VTAIL.n120 585
R43 VTAIL.n132 VTAIL.n131 585
R44 VTAIL.n130 VTAIL.n129 585
R45 VTAIL.n125 VTAIL.n124 585
R46 VTAIL.n103 VTAIL.n102 585
R47 VTAIL.n101 VTAIL.n100 585
R48 VTAIL.n58 VTAIL.n57 585
R49 VTAIL.n95 VTAIL.n94 585
R50 VTAIL.n93 VTAIL.n60 585
R51 VTAIL.n92 VTAIL.n91 585
R52 VTAIL.n63 VTAIL.n61 585
R53 VTAIL.n86 VTAIL.n85 585
R54 VTAIL.n84 VTAIL.n83 585
R55 VTAIL.n67 VTAIL.n66 585
R56 VTAIL.n78 VTAIL.n77 585
R57 VTAIL.n76 VTAIL.n75 585
R58 VTAIL.n71 VTAIL.n70 585
R59 VTAIL.n179 VTAIL.t1 329.038
R60 VTAIL.n17 VTAIL.t2 329.038
R61 VTAIL.n126 VTAIL.t3 329.038
R62 VTAIL.n72 VTAIL.t0 329.038
R63 VTAIL.n183 VTAIL.n177 171.744
R64 VTAIL.n184 VTAIL.n183 171.744
R65 VTAIL.n184 VTAIL.n173 171.744
R66 VTAIL.n191 VTAIL.n173 171.744
R67 VTAIL.n192 VTAIL.n191 171.744
R68 VTAIL.n192 VTAIL.n169 171.744
R69 VTAIL.n200 VTAIL.n169 171.744
R70 VTAIL.n201 VTAIL.n200 171.744
R71 VTAIL.n202 VTAIL.n201 171.744
R72 VTAIL.n202 VTAIL.n165 171.744
R73 VTAIL.n209 VTAIL.n165 171.744
R74 VTAIL.n210 VTAIL.n209 171.744
R75 VTAIL.n21 VTAIL.n15 171.744
R76 VTAIL.n22 VTAIL.n21 171.744
R77 VTAIL.n22 VTAIL.n11 171.744
R78 VTAIL.n29 VTAIL.n11 171.744
R79 VTAIL.n30 VTAIL.n29 171.744
R80 VTAIL.n30 VTAIL.n7 171.744
R81 VTAIL.n38 VTAIL.n7 171.744
R82 VTAIL.n39 VTAIL.n38 171.744
R83 VTAIL.n40 VTAIL.n39 171.744
R84 VTAIL.n40 VTAIL.n3 171.744
R85 VTAIL.n47 VTAIL.n3 171.744
R86 VTAIL.n48 VTAIL.n47 171.744
R87 VTAIL.n156 VTAIL.n155 171.744
R88 VTAIL.n155 VTAIL.n111 171.744
R89 VTAIL.n148 VTAIL.n111 171.744
R90 VTAIL.n148 VTAIL.n147 171.744
R91 VTAIL.n147 VTAIL.n146 171.744
R92 VTAIL.n146 VTAIL.n115 171.744
R93 VTAIL.n139 VTAIL.n115 171.744
R94 VTAIL.n139 VTAIL.n138 171.744
R95 VTAIL.n138 VTAIL.n120 171.744
R96 VTAIL.n131 VTAIL.n120 171.744
R97 VTAIL.n131 VTAIL.n130 171.744
R98 VTAIL.n130 VTAIL.n124 171.744
R99 VTAIL.n102 VTAIL.n101 171.744
R100 VTAIL.n101 VTAIL.n57 171.744
R101 VTAIL.n94 VTAIL.n57 171.744
R102 VTAIL.n94 VTAIL.n93 171.744
R103 VTAIL.n93 VTAIL.n92 171.744
R104 VTAIL.n92 VTAIL.n61 171.744
R105 VTAIL.n85 VTAIL.n61 171.744
R106 VTAIL.n85 VTAIL.n84 171.744
R107 VTAIL.n84 VTAIL.n66 171.744
R108 VTAIL.n77 VTAIL.n66 171.744
R109 VTAIL.n77 VTAIL.n76 171.744
R110 VTAIL.n76 VTAIL.n70 171.744
R111 VTAIL.t1 VTAIL.n177 85.8723
R112 VTAIL.t2 VTAIL.n15 85.8723
R113 VTAIL.t3 VTAIL.n124 85.8723
R114 VTAIL.t0 VTAIL.n70 85.8723
R115 VTAIL.n215 VTAIL.n214 34.7066
R116 VTAIL.n53 VTAIL.n52 34.7066
R117 VTAIL.n161 VTAIL.n160 34.7066
R118 VTAIL.n107 VTAIL.n106 34.7066
R119 VTAIL.n107 VTAIL.n53 23.1341
R120 VTAIL.n215 VTAIL.n161 22.1083
R121 VTAIL.n203 VTAIL.n168 13.1884
R122 VTAIL.n41 VTAIL.n6 13.1884
R123 VTAIL.n149 VTAIL.n114 13.1884
R124 VTAIL.n95 VTAIL.n60 13.1884
R125 VTAIL.n199 VTAIL.n198 12.8005
R126 VTAIL.n204 VTAIL.n166 12.8005
R127 VTAIL.n37 VTAIL.n36 12.8005
R128 VTAIL.n42 VTAIL.n4 12.8005
R129 VTAIL.n150 VTAIL.n112 12.8005
R130 VTAIL.n145 VTAIL.n116 12.8005
R131 VTAIL.n96 VTAIL.n58 12.8005
R132 VTAIL.n91 VTAIL.n62 12.8005
R133 VTAIL.n197 VTAIL.n170 12.0247
R134 VTAIL.n208 VTAIL.n207 12.0247
R135 VTAIL.n35 VTAIL.n8 12.0247
R136 VTAIL.n46 VTAIL.n45 12.0247
R137 VTAIL.n154 VTAIL.n153 12.0247
R138 VTAIL.n144 VTAIL.n117 12.0247
R139 VTAIL.n100 VTAIL.n99 12.0247
R140 VTAIL.n90 VTAIL.n63 12.0247
R141 VTAIL.n194 VTAIL.n193 11.249
R142 VTAIL.n211 VTAIL.n164 11.249
R143 VTAIL.n32 VTAIL.n31 11.249
R144 VTAIL.n49 VTAIL.n2 11.249
R145 VTAIL.n157 VTAIL.n110 11.249
R146 VTAIL.n141 VTAIL.n140 11.249
R147 VTAIL.n103 VTAIL.n56 11.249
R148 VTAIL.n87 VTAIL.n86 11.249
R149 VTAIL.n179 VTAIL.n178 10.7239
R150 VTAIL.n17 VTAIL.n16 10.7239
R151 VTAIL.n126 VTAIL.n125 10.7239
R152 VTAIL.n72 VTAIL.n71 10.7239
R153 VTAIL.n190 VTAIL.n172 10.4732
R154 VTAIL.n212 VTAIL.n162 10.4732
R155 VTAIL.n28 VTAIL.n10 10.4732
R156 VTAIL.n50 VTAIL.n0 10.4732
R157 VTAIL.n158 VTAIL.n108 10.4732
R158 VTAIL.n137 VTAIL.n119 10.4732
R159 VTAIL.n104 VTAIL.n54 10.4732
R160 VTAIL.n83 VTAIL.n65 10.4732
R161 VTAIL.n189 VTAIL.n174 9.69747
R162 VTAIL.n27 VTAIL.n12 9.69747
R163 VTAIL.n136 VTAIL.n121 9.69747
R164 VTAIL.n82 VTAIL.n67 9.69747
R165 VTAIL.n214 VTAIL.n213 9.45567
R166 VTAIL.n52 VTAIL.n51 9.45567
R167 VTAIL.n160 VTAIL.n159 9.45567
R168 VTAIL.n106 VTAIL.n105 9.45567
R169 VTAIL.n213 VTAIL.n212 9.3005
R170 VTAIL.n164 VTAIL.n163 9.3005
R171 VTAIL.n207 VTAIL.n206 9.3005
R172 VTAIL.n205 VTAIL.n204 9.3005
R173 VTAIL.n181 VTAIL.n180 9.3005
R174 VTAIL.n176 VTAIL.n175 9.3005
R175 VTAIL.n187 VTAIL.n186 9.3005
R176 VTAIL.n189 VTAIL.n188 9.3005
R177 VTAIL.n172 VTAIL.n171 9.3005
R178 VTAIL.n195 VTAIL.n194 9.3005
R179 VTAIL.n197 VTAIL.n196 9.3005
R180 VTAIL.n198 VTAIL.n167 9.3005
R181 VTAIL.n51 VTAIL.n50 9.3005
R182 VTAIL.n2 VTAIL.n1 9.3005
R183 VTAIL.n45 VTAIL.n44 9.3005
R184 VTAIL.n43 VTAIL.n42 9.3005
R185 VTAIL.n19 VTAIL.n18 9.3005
R186 VTAIL.n14 VTAIL.n13 9.3005
R187 VTAIL.n25 VTAIL.n24 9.3005
R188 VTAIL.n27 VTAIL.n26 9.3005
R189 VTAIL.n10 VTAIL.n9 9.3005
R190 VTAIL.n33 VTAIL.n32 9.3005
R191 VTAIL.n35 VTAIL.n34 9.3005
R192 VTAIL.n36 VTAIL.n5 9.3005
R193 VTAIL.n128 VTAIL.n127 9.3005
R194 VTAIL.n123 VTAIL.n122 9.3005
R195 VTAIL.n134 VTAIL.n133 9.3005
R196 VTAIL.n136 VTAIL.n135 9.3005
R197 VTAIL.n119 VTAIL.n118 9.3005
R198 VTAIL.n142 VTAIL.n141 9.3005
R199 VTAIL.n144 VTAIL.n143 9.3005
R200 VTAIL.n116 VTAIL.n113 9.3005
R201 VTAIL.n159 VTAIL.n158 9.3005
R202 VTAIL.n110 VTAIL.n109 9.3005
R203 VTAIL.n153 VTAIL.n152 9.3005
R204 VTAIL.n151 VTAIL.n150 9.3005
R205 VTAIL.n74 VTAIL.n73 9.3005
R206 VTAIL.n69 VTAIL.n68 9.3005
R207 VTAIL.n80 VTAIL.n79 9.3005
R208 VTAIL.n82 VTAIL.n81 9.3005
R209 VTAIL.n65 VTAIL.n64 9.3005
R210 VTAIL.n88 VTAIL.n87 9.3005
R211 VTAIL.n90 VTAIL.n89 9.3005
R212 VTAIL.n62 VTAIL.n59 9.3005
R213 VTAIL.n105 VTAIL.n104 9.3005
R214 VTAIL.n56 VTAIL.n55 9.3005
R215 VTAIL.n99 VTAIL.n98 9.3005
R216 VTAIL.n97 VTAIL.n96 9.3005
R217 VTAIL.n186 VTAIL.n185 8.92171
R218 VTAIL.n24 VTAIL.n23 8.92171
R219 VTAIL.n133 VTAIL.n132 8.92171
R220 VTAIL.n79 VTAIL.n78 8.92171
R221 VTAIL.n182 VTAIL.n176 8.14595
R222 VTAIL.n20 VTAIL.n14 8.14595
R223 VTAIL.n129 VTAIL.n123 8.14595
R224 VTAIL.n75 VTAIL.n69 8.14595
R225 VTAIL.n181 VTAIL.n178 7.3702
R226 VTAIL.n19 VTAIL.n16 7.3702
R227 VTAIL.n128 VTAIL.n125 7.3702
R228 VTAIL.n74 VTAIL.n71 7.3702
R229 VTAIL.n182 VTAIL.n181 5.81868
R230 VTAIL.n20 VTAIL.n19 5.81868
R231 VTAIL.n129 VTAIL.n128 5.81868
R232 VTAIL.n75 VTAIL.n74 5.81868
R233 VTAIL.n185 VTAIL.n176 5.04292
R234 VTAIL.n23 VTAIL.n14 5.04292
R235 VTAIL.n132 VTAIL.n123 5.04292
R236 VTAIL.n78 VTAIL.n69 5.04292
R237 VTAIL.n186 VTAIL.n174 4.26717
R238 VTAIL.n24 VTAIL.n12 4.26717
R239 VTAIL.n133 VTAIL.n121 4.26717
R240 VTAIL.n79 VTAIL.n67 4.26717
R241 VTAIL.n190 VTAIL.n189 3.49141
R242 VTAIL.n214 VTAIL.n162 3.49141
R243 VTAIL.n28 VTAIL.n27 3.49141
R244 VTAIL.n52 VTAIL.n0 3.49141
R245 VTAIL.n160 VTAIL.n108 3.49141
R246 VTAIL.n137 VTAIL.n136 3.49141
R247 VTAIL.n106 VTAIL.n54 3.49141
R248 VTAIL.n83 VTAIL.n82 3.49141
R249 VTAIL.n193 VTAIL.n172 2.71565
R250 VTAIL.n212 VTAIL.n211 2.71565
R251 VTAIL.n31 VTAIL.n10 2.71565
R252 VTAIL.n50 VTAIL.n49 2.71565
R253 VTAIL.n158 VTAIL.n157 2.71565
R254 VTAIL.n140 VTAIL.n119 2.71565
R255 VTAIL.n104 VTAIL.n103 2.71565
R256 VTAIL.n86 VTAIL.n65 2.71565
R257 VTAIL.n180 VTAIL.n179 2.41283
R258 VTAIL.n18 VTAIL.n17 2.41283
R259 VTAIL.n127 VTAIL.n126 2.41283
R260 VTAIL.n73 VTAIL.n72 2.41283
R261 VTAIL.n194 VTAIL.n170 1.93989
R262 VTAIL.n208 VTAIL.n164 1.93989
R263 VTAIL.n32 VTAIL.n8 1.93989
R264 VTAIL.n46 VTAIL.n2 1.93989
R265 VTAIL.n154 VTAIL.n110 1.93989
R266 VTAIL.n141 VTAIL.n117 1.93989
R267 VTAIL.n100 VTAIL.n56 1.93989
R268 VTAIL.n87 VTAIL.n63 1.93989
R269 VTAIL.n199 VTAIL.n197 1.16414
R270 VTAIL.n207 VTAIL.n166 1.16414
R271 VTAIL.n37 VTAIL.n35 1.16414
R272 VTAIL.n45 VTAIL.n4 1.16414
R273 VTAIL.n153 VTAIL.n112 1.16414
R274 VTAIL.n145 VTAIL.n144 1.16414
R275 VTAIL.n99 VTAIL.n58 1.16414
R276 VTAIL.n91 VTAIL.n90 1.16414
R277 VTAIL.n161 VTAIL.n107 0.983259
R278 VTAIL VTAIL.n53 0.784983
R279 VTAIL.n198 VTAIL.n168 0.388379
R280 VTAIL.n204 VTAIL.n203 0.388379
R281 VTAIL.n36 VTAIL.n6 0.388379
R282 VTAIL.n42 VTAIL.n41 0.388379
R283 VTAIL.n150 VTAIL.n149 0.388379
R284 VTAIL.n116 VTAIL.n114 0.388379
R285 VTAIL.n96 VTAIL.n95 0.388379
R286 VTAIL.n62 VTAIL.n60 0.388379
R287 VTAIL VTAIL.n215 0.198776
R288 VTAIL.n180 VTAIL.n175 0.155672
R289 VTAIL.n187 VTAIL.n175 0.155672
R290 VTAIL.n188 VTAIL.n187 0.155672
R291 VTAIL.n188 VTAIL.n171 0.155672
R292 VTAIL.n195 VTAIL.n171 0.155672
R293 VTAIL.n196 VTAIL.n195 0.155672
R294 VTAIL.n196 VTAIL.n167 0.155672
R295 VTAIL.n205 VTAIL.n167 0.155672
R296 VTAIL.n206 VTAIL.n205 0.155672
R297 VTAIL.n206 VTAIL.n163 0.155672
R298 VTAIL.n213 VTAIL.n163 0.155672
R299 VTAIL.n18 VTAIL.n13 0.155672
R300 VTAIL.n25 VTAIL.n13 0.155672
R301 VTAIL.n26 VTAIL.n25 0.155672
R302 VTAIL.n26 VTAIL.n9 0.155672
R303 VTAIL.n33 VTAIL.n9 0.155672
R304 VTAIL.n34 VTAIL.n33 0.155672
R305 VTAIL.n34 VTAIL.n5 0.155672
R306 VTAIL.n43 VTAIL.n5 0.155672
R307 VTAIL.n44 VTAIL.n43 0.155672
R308 VTAIL.n44 VTAIL.n1 0.155672
R309 VTAIL.n51 VTAIL.n1 0.155672
R310 VTAIL.n159 VTAIL.n109 0.155672
R311 VTAIL.n152 VTAIL.n109 0.155672
R312 VTAIL.n152 VTAIL.n151 0.155672
R313 VTAIL.n151 VTAIL.n113 0.155672
R314 VTAIL.n143 VTAIL.n113 0.155672
R315 VTAIL.n143 VTAIL.n142 0.155672
R316 VTAIL.n142 VTAIL.n118 0.155672
R317 VTAIL.n135 VTAIL.n118 0.155672
R318 VTAIL.n135 VTAIL.n134 0.155672
R319 VTAIL.n134 VTAIL.n122 0.155672
R320 VTAIL.n127 VTAIL.n122 0.155672
R321 VTAIL.n105 VTAIL.n55 0.155672
R322 VTAIL.n98 VTAIL.n55 0.155672
R323 VTAIL.n98 VTAIL.n97 0.155672
R324 VTAIL.n97 VTAIL.n59 0.155672
R325 VTAIL.n89 VTAIL.n59 0.155672
R326 VTAIL.n89 VTAIL.n88 0.155672
R327 VTAIL.n88 VTAIL.n64 0.155672
R328 VTAIL.n81 VTAIL.n64 0.155672
R329 VTAIL.n81 VTAIL.n80 0.155672
R330 VTAIL.n80 VTAIL.n68 0.155672
R331 VTAIL.n73 VTAIL.n68 0.155672
R332 VDD1.n48 VDD1.n0 756.745
R333 VDD1.n101 VDD1.n53 756.745
R334 VDD1.n49 VDD1.n48 585
R335 VDD1.n47 VDD1.n46 585
R336 VDD1.n4 VDD1.n3 585
R337 VDD1.n41 VDD1.n40 585
R338 VDD1.n39 VDD1.n6 585
R339 VDD1.n38 VDD1.n37 585
R340 VDD1.n9 VDD1.n7 585
R341 VDD1.n32 VDD1.n31 585
R342 VDD1.n30 VDD1.n29 585
R343 VDD1.n13 VDD1.n12 585
R344 VDD1.n24 VDD1.n23 585
R345 VDD1.n22 VDD1.n21 585
R346 VDD1.n17 VDD1.n16 585
R347 VDD1.n69 VDD1.n68 585
R348 VDD1.n74 VDD1.n73 585
R349 VDD1.n76 VDD1.n75 585
R350 VDD1.n65 VDD1.n64 585
R351 VDD1.n82 VDD1.n81 585
R352 VDD1.n84 VDD1.n83 585
R353 VDD1.n61 VDD1.n60 585
R354 VDD1.n91 VDD1.n90 585
R355 VDD1.n92 VDD1.n59 585
R356 VDD1.n94 VDD1.n93 585
R357 VDD1.n57 VDD1.n56 585
R358 VDD1.n100 VDD1.n99 585
R359 VDD1.n102 VDD1.n101 585
R360 VDD1.n70 VDD1.t0 329.038
R361 VDD1.n18 VDD1.t1 329.038
R362 VDD1.n48 VDD1.n47 171.744
R363 VDD1.n47 VDD1.n3 171.744
R364 VDD1.n40 VDD1.n3 171.744
R365 VDD1.n40 VDD1.n39 171.744
R366 VDD1.n39 VDD1.n38 171.744
R367 VDD1.n38 VDD1.n7 171.744
R368 VDD1.n31 VDD1.n7 171.744
R369 VDD1.n31 VDD1.n30 171.744
R370 VDD1.n30 VDD1.n12 171.744
R371 VDD1.n23 VDD1.n12 171.744
R372 VDD1.n23 VDD1.n22 171.744
R373 VDD1.n22 VDD1.n16 171.744
R374 VDD1.n74 VDD1.n68 171.744
R375 VDD1.n75 VDD1.n74 171.744
R376 VDD1.n75 VDD1.n64 171.744
R377 VDD1.n82 VDD1.n64 171.744
R378 VDD1.n83 VDD1.n82 171.744
R379 VDD1.n83 VDD1.n60 171.744
R380 VDD1.n91 VDD1.n60 171.744
R381 VDD1.n92 VDD1.n91 171.744
R382 VDD1.n93 VDD1.n92 171.744
R383 VDD1.n93 VDD1.n56 171.744
R384 VDD1.n100 VDD1.n56 171.744
R385 VDD1.n101 VDD1.n100 171.744
R386 VDD1 VDD1.n105 86.5933
R387 VDD1.t1 VDD1.n16 85.8723
R388 VDD1.t0 VDD1.n68 85.8723
R389 VDD1 VDD1.n52 51.7
R390 VDD1.n41 VDD1.n6 13.1884
R391 VDD1.n94 VDD1.n59 13.1884
R392 VDD1.n42 VDD1.n4 12.8005
R393 VDD1.n37 VDD1.n8 12.8005
R394 VDD1.n90 VDD1.n89 12.8005
R395 VDD1.n95 VDD1.n57 12.8005
R396 VDD1.n46 VDD1.n45 12.0247
R397 VDD1.n36 VDD1.n9 12.0247
R398 VDD1.n88 VDD1.n61 12.0247
R399 VDD1.n99 VDD1.n98 12.0247
R400 VDD1.n49 VDD1.n2 11.249
R401 VDD1.n33 VDD1.n32 11.249
R402 VDD1.n85 VDD1.n84 11.249
R403 VDD1.n102 VDD1.n55 11.249
R404 VDD1.n18 VDD1.n17 10.7239
R405 VDD1.n70 VDD1.n69 10.7239
R406 VDD1.n50 VDD1.n0 10.4732
R407 VDD1.n29 VDD1.n11 10.4732
R408 VDD1.n81 VDD1.n63 10.4732
R409 VDD1.n103 VDD1.n53 10.4732
R410 VDD1.n28 VDD1.n13 9.69747
R411 VDD1.n80 VDD1.n65 9.69747
R412 VDD1.n52 VDD1.n51 9.45567
R413 VDD1.n105 VDD1.n104 9.45567
R414 VDD1.n20 VDD1.n19 9.3005
R415 VDD1.n15 VDD1.n14 9.3005
R416 VDD1.n26 VDD1.n25 9.3005
R417 VDD1.n28 VDD1.n27 9.3005
R418 VDD1.n11 VDD1.n10 9.3005
R419 VDD1.n34 VDD1.n33 9.3005
R420 VDD1.n36 VDD1.n35 9.3005
R421 VDD1.n8 VDD1.n5 9.3005
R422 VDD1.n51 VDD1.n50 9.3005
R423 VDD1.n2 VDD1.n1 9.3005
R424 VDD1.n45 VDD1.n44 9.3005
R425 VDD1.n43 VDD1.n42 9.3005
R426 VDD1.n104 VDD1.n103 9.3005
R427 VDD1.n55 VDD1.n54 9.3005
R428 VDD1.n98 VDD1.n97 9.3005
R429 VDD1.n96 VDD1.n95 9.3005
R430 VDD1.n72 VDD1.n71 9.3005
R431 VDD1.n67 VDD1.n66 9.3005
R432 VDD1.n78 VDD1.n77 9.3005
R433 VDD1.n80 VDD1.n79 9.3005
R434 VDD1.n63 VDD1.n62 9.3005
R435 VDD1.n86 VDD1.n85 9.3005
R436 VDD1.n88 VDD1.n87 9.3005
R437 VDD1.n89 VDD1.n58 9.3005
R438 VDD1.n25 VDD1.n24 8.92171
R439 VDD1.n77 VDD1.n76 8.92171
R440 VDD1.n21 VDD1.n15 8.14595
R441 VDD1.n73 VDD1.n67 8.14595
R442 VDD1.n20 VDD1.n17 7.3702
R443 VDD1.n72 VDD1.n69 7.3702
R444 VDD1.n21 VDD1.n20 5.81868
R445 VDD1.n73 VDD1.n72 5.81868
R446 VDD1.n24 VDD1.n15 5.04292
R447 VDD1.n76 VDD1.n67 5.04292
R448 VDD1.n25 VDD1.n13 4.26717
R449 VDD1.n77 VDD1.n65 4.26717
R450 VDD1.n52 VDD1.n0 3.49141
R451 VDD1.n29 VDD1.n28 3.49141
R452 VDD1.n81 VDD1.n80 3.49141
R453 VDD1.n105 VDD1.n53 3.49141
R454 VDD1.n50 VDD1.n49 2.71565
R455 VDD1.n32 VDD1.n11 2.71565
R456 VDD1.n84 VDD1.n63 2.71565
R457 VDD1.n103 VDD1.n102 2.71565
R458 VDD1.n19 VDD1.n18 2.41283
R459 VDD1.n71 VDD1.n70 2.41283
R460 VDD1.n46 VDD1.n2 1.93989
R461 VDD1.n33 VDD1.n9 1.93989
R462 VDD1.n85 VDD1.n61 1.93989
R463 VDD1.n99 VDD1.n55 1.93989
R464 VDD1.n45 VDD1.n4 1.16414
R465 VDD1.n37 VDD1.n36 1.16414
R466 VDD1.n90 VDD1.n88 1.16414
R467 VDD1.n98 VDD1.n57 1.16414
R468 VDD1.n42 VDD1.n41 0.388379
R469 VDD1.n8 VDD1.n6 0.388379
R470 VDD1.n89 VDD1.n59 0.388379
R471 VDD1.n95 VDD1.n94 0.388379
R472 VDD1.n51 VDD1.n1 0.155672
R473 VDD1.n44 VDD1.n1 0.155672
R474 VDD1.n44 VDD1.n43 0.155672
R475 VDD1.n43 VDD1.n5 0.155672
R476 VDD1.n35 VDD1.n5 0.155672
R477 VDD1.n35 VDD1.n34 0.155672
R478 VDD1.n34 VDD1.n10 0.155672
R479 VDD1.n27 VDD1.n10 0.155672
R480 VDD1.n27 VDD1.n26 0.155672
R481 VDD1.n26 VDD1.n14 0.155672
R482 VDD1.n19 VDD1.n14 0.155672
R483 VDD1.n71 VDD1.n66 0.155672
R484 VDD1.n78 VDD1.n66 0.155672
R485 VDD1.n79 VDD1.n78 0.155672
R486 VDD1.n79 VDD1.n62 0.155672
R487 VDD1.n86 VDD1.n62 0.155672
R488 VDD1.n87 VDD1.n86 0.155672
R489 VDD1.n87 VDD1.n58 0.155672
R490 VDD1.n96 VDD1.n58 0.155672
R491 VDD1.n97 VDD1.n96 0.155672
R492 VDD1.n97 VDD1.n54 0.155672
R493 VDD1.n104 VDD1.n54 0.155672
R494 B.n316 B.n55 585
R495 B.n318 B.n317 585
R496 B.n319 B.n54 585
R497 B.n321 B.n320 585
R498 B.n322 B.n53 585
R499 B.n324 B.n323 585
R500 B.n325 B.n52 585
R501 B.n327 B.n326 585
R502 B.n328 B.n51 585
R503 B.n330 B.n329 585
R504 B.n331 B.n50 585
R505 B.n333 B.n332 585
R506 B.n334 B.n49 585
R507 B.n336 B.n335 585
R508 B.n337 B.n48 585
R509 B.n339 B.n338 585
R510 B.n340 B.n47 585
R511 B.n342 B.n341 585
R512 B.n343 B.n46 585
R513 B.n345 B.n344 585
R514 B.n346 B.n45 585
R515 B.n348 B.n347 585
R516 B.n349 B.n44 585
R517 B.n351 B.n350 585
R518 B.n352 B.n43 585
R519 B.n354 B.n353 585
R520 B.n355 B.n42 585
R521 B.n357 B.n356 585
R522 B.n358 B.n41 585
R523 B.n360 B.n359 585
R524 B.n361 B.n40 585
R525 B.n363 B.n362 585
R526 B.n364 B.n39 585
R527 B.n366 B.n365 585
R528 B.n367 B.n35 585
R529 B.n369 B.n368 585
R530 B.n370 B.n34 585
R531 B.n372 B.n371 585
R532 B.n373 B.n33 585
R533 B.n375 B.n374 585
R534 B.n376 B.n32 585
R535 B.n378 B.n377 585
R536 B.n379 B.n31 585
R537 B.n381 B.n380 585
R538 B.n382 B.n30 585
R539 B.n384 B.n383 585
R540 B.n386 B.n27 585
R541 B.n388 B.n387 585
R542 B.n389 B.n26 585
R543 B.n391 B.n390 585
R544 B.n392 B.n25 585
R545 B.n394 B.n393 585
R546 B.n395 B.n24 585
R547 B.n397 B.n396 585
R548 B.n398 B.n23 585
R549 B.n400 B.n399 585
R550 B.n401 B.n22 585
R551 B.n403 B.n402 585
R552 B.n404 B.n21 585
R553 B.n406 B.n405 585
R554 B.n407 B.n20 585
R555 B.n409 B.n408 585
R556 B.n410 B.n19 585
R557 B.n412 B.n411 585
R558 B.n413 B.n18 585
R559 B.n415 B.n414 585
R560 B.n416 B.n17 585
R561 B.n418 B.n417 585
R562 B.n419 B.n16 585
R563 B.n421 B.n420 585
R564 B.n422 B.n15 585
R565 B.n424 B.n423 585
R566 B.n425 B.n14 585
R567 B.n427 B.n426 585
R568 B.n428 B.n13 585
R569 B.n430 B.n429 585
R570 B.n431 B.n12 585
R571 B.n433 B.n432 585
R572 B.n434 B.n11 585
R573 B.n436 B.n435 585
R574 B.n437 B.n10 585
R575 B.n439 B.n438 585
R576 B.n315 B.n314 585
R577 B.n313 B.n56 585
R578 B.n312 B.n311 585
R579 B.n310 B.n57 585
R580 B.n309 B.n308 585
R581 B.n307 B.n58 585
R582 B.n306 B.n305 585
R583 B.n304 B.n59 585
R584 B.n303 B.n302 585
R585 B.n301 B.n60 585
R586 B.n300 B.n299 585
R587 B.n298 B.n61 585
R588 B.n297 B.n296 585
R589 B.n295 B.n62 585
R590 B.n294 B.n293 585
R591 B.n292 B.n63 585
R592 B.n291 B.n290 585
R593 B.n289 B.n64 585
R594 B.n288 B.n287 585
R595 B.n286 B.n65 585
R596 B.n285 B.n284 585
R597 B.n283 B.n66 585
R598 B.n282 B.n281 585
R599 B.n280 B.n67 585
R600 B.n279 B.n278 585
R601 B.n277 B.n68 585
R602 B.n276 B.n275 585
R603 B.n274 B.n69 585
R604 B.n273 B.n272 585
R605 B.n271 B.n70 585
R606 B.n270 B.n269 585
R607 B.n145 B.n116 585
R608 B.n147 B.n146 585
R609 B.n148 B.n115 585
R610 B.n150 B.n149 585
R611 B.n151 B.n114 585
R612 B.n153 B.n152 585
R613 B.n154 B.n113 585
R614 B.n156 B.n155 585
R615 B.n157 B.n112 585
R616 B.n159 B.n158 585
R617 B.n160 B.n111 585
R618 B.n162 B.n161 585
R619 B.n163 B.n110 585
R620 B.n165 B.n164 585
R621 B.n166 B.n109 585
R622 B.n168 B.n167 585
R623 B.n169 B.n108 585
R624 B.n171 B.n170 585
R625 B.n172 B.n107 585
R626 B.n174 B.n173 585
R627 B.n175 B.n106 585
R628 B.n177 B.n176 585
R629 B.n178 B.n105 585
R630 B.n180 B.n179 585
R631 B.n181 B.n104 585
R632 B.n183 B.n182 585
R633 B.n184 B.n103 585
R634 B.n186 B.n185 585
R635 B.n187 B.n102 585
R636 B.n189 B.n188 585
R637 B.n190 B.n101 585
R638 B.n192 B.n191 585
R639 B.n193 B.n100 585
R640 B.n195 B.n194 585
R641 B.n196 B.n99 585
R642 B.n198 B.n197 585
R643 B.n200 B.n96 585
R644 B.n202 B.n201 585
R645 B.n203 B.n95 585
R646 B.n205 B.n204 585
R647 B.n206 B.n94 585
R648 B.n208 B.n207 585
R649 B.n209 B.n93 585
R650 B.n211 B.n210 585
R651 B.n212 B.n92 585
R652 B.n214 B.n213 585
R653 B.n216 B.n215 585
R654 B.n217 B.n88 585
R655 B.n219 B.n218 585
R656 B.n220 B.n87 585
R657 B.n222 B.n221 585
R658 B.n223 B.n86 585
R659 B.n225 B.n224 585
R660 B.n226 B.n85 585
R661 B.n228 B.n227 585
R662 B.n229 B.n84 585
R663 B.n231 B.n230 585
R664 B.n232 B.n83 585
R665 B.n234 B.n233 585
R666 B.n235 B.n82 585
R667 B.n237 B.n236 585
R668 B.n238 B.n81 585
R669 B.n240 B.n239 585
R670 B.n241 B.n80 585
R671 B.n243 B.n242 585
R672 B.n244 B.n79 585
R673 B.n246 B.n245 585
R674 B.n247 B.n78 585
R675 B.n249 B.n248 585
R676 B.n250 B.n77 585
R677 B.n252 B.n251 585
R678 B.n253 B.n76 585
R679 B.n255 B.n254 585
R680 B.n256 B.n75 585
R681 B.n258 B.n257 585
R682 B.n259 B.n74 585
R683 B.n261 B.n260 585
R684 B.n262 B.n73 585
R685 B.n264 B.n263 585
R686 B.n265 B.n72 585
R687 B.n267 B.n266 585
R688 B.n268 B.n71 585
R689 B.n144 B.n143 585
R690 B.n142 B.n117 585
R691 B.n141 B.n140 585
R692 B.n139 B.n118 585
R693 B.n138 B.n137 585
R694 B.n136 B.n119 585
R695 B.n135 B.n134 585
R696 B.n133 B.n120 585
R697 B.n132 B.n131 585
R698 B.n130 B.n121 585
R699 B.n129 B.n128 585
R700 B.n127 B.n122 585
R701 B.n126 B.n125 585
R702 B.n124 B.n123 585
R703 B.n2 B.n0 585
R704 B.n461 B.n1 585
R705 B.n460 B.n459 585
R706 B.n458 B.n3 585
R707 B.n457 B.n456 585
R708 B.n455 B.n4 585
R709 B.n454 B.n453 585
R710 B.n452 B.n5 585
R711 B.n451 B.n450 585
R712 B.n449 B.n6 585
R713 B.n448 B.n447 585
R714 B.n446 B.n7 585
R715 B.n445 B.n444 585
R716 B.n443 B.n8 585
R717 B.n442 B.n441 585
R718 B.n440 B.n9 585
R719 B.n463 B.n462 585
R720 B.n143 B.n116 492.5
R721 B.n438 B.n9 492.5
R722 B.n269 B.n268 492.5
R723 B.n316 B.n315 492.5
R724 B.n89 B.t9 484.627
R725 B.n97 B.t6 484.627
R726 B.n28 B.t0 484.627
R727 B.n36 B.t3 484.627
R728 B.n89 B.t11 364.401
R729 B.n36 B.t4 364.401
R730 B.n97 B.t8 364.401
R731 B.n28 B.t1 364.401
R732 B.n90 B.t10 341.322
R733 B.n37 B.t5 341.322
R734 B.n98 B.t7 341.322
R735 B.n29 B.t2 341.322
R736 B.n143 B.n142 163.367
R737 B.n142 B.n141 163.367
R738 B.n141 B.n118 163.367
R739 B.n137 B.n118 163.367
R740 B.n137 B.n136 163.367
R741 B.n136 B.n135 163.367
R742 B.n135 B.n120 163.367
R743 B.n131 B.n120 163.367
R744 B.n131 B.n130 163.367
R745 B.n130 B.n129 163.367
R746 B.n129 B.n122 163.367
R747 B.n125 B.n122 163.367
R748 B.n125 B.n124 163.367
R749 B.n124 B.n2 163.367
R750 B.n462 B.n2 163.367
R751 B.n462 B.n461 163.367
R752 B.n461 B.n460 163.367
R753 B.n460 B.n3 163.367
R754 B.n456 B.n3 163.367
R755 B.n456 B.n455 163.367
R756 B.n455 B.n454 163.367
R757 B.n454 B.n5 163.367
R758 B.n450 B.n5 163.367
R759 B.n450 B.n449 163.367
R760 B.n449 B.n448 163.367
R761 B.n448 B.n7 163.367
R762 B.n444 B.n7 163.367
R763 B.n444 B.n443 163.367
R764 B.n443 B.n442 163.367
R765 B.n442 B.n9 163.367
R766 B.n147 B.n116 163.367
R767 B.n148 B.n147 163.367
R768 B.n149 B.n148 163.367
R769 B.n149 B.n114 163.367
R770 B.n153 B.n114 163.367
R771 B.n154 B.n153 163.367
R772 B.n155 B.n154 163.367
R773 B.n155 B.n112 163.367
R774 B.n159 B.n112 163.367
R775 B.n160 B.n159 163.367
R776 B.n161 B.n160 163.367
R777 B.n161 B.n110 163.367
R778 B.n165 B.n110 163.367
R779 B.n166 B.n165 163.367
R780 B.n167 B.n166 163.367
R781 B.n167 B.n108 163.367
R782 B.n171 B.n108 163.367
R783 B.n172 B.n171 163.367
R784 B.n173 B.n172 163.367
R785 B.n173 B.n106 163.367
R786 B.n177 B.n106 163.367
R787 B.n178 B.n177 163.367
R788 B.n179 B.n178 163.367
R789 B.n179 B.n104 163.367
R790 B.n183 B.n104 163.367
R791 B.n184 B.n183 163.367
R792 B.n185 B.n184 163.367
R793 B.n185 B.n102 163.367
R794 B.n189 B.n102 163.367
R795 B.n190 B.n189 163.367
R796 B.n191 B.n190 163.367
R797 B.n191 B.n100 163.367
R798 B.n195 B.n100 163.367
R799 B.n196 B.n195 163.367
R800 B.n197 B.n196 163.367
R801 B.n197 B.n96 163.367
R802 B.n202 B.n96 163.367
R803 B.n203 B.n202 163.367
R804 B.n204 B.n203 163.367
R805 B.n204 B.n94 163.367
R806 B.n208 B.n94 163.367
R807 B.n209 B.n208 163.367
R808 B.n210 B.n209 163.367
R809 B.n210 B.n92 163.367
R810 B.n214 B.n92 163.367
R811 B.n215 B.n214 163.367
R812 B.n215 B.n88 163.367
R813 B.n219 B.n88 163.367
R814 B.n220 B.n219 163.367
R815 B.n221 B.n220 163.367
R816 B.n221 B.n86 163.367
R817 B.n225 B.n86 163.367
R818 B.n226 B.n225 163.367
R819 B.n227 B.n226 163.367
R820 B.n227 B.n84 163.367
R821 B.n231 B.n84 163.367
R822 B.n232 B.n231 163.367
R823 B.n233 B.n232 163.367
R824 B.n233 B.n82 163.367
R825 B.n237 B.n82 163.367
R826 B.n238 B.n237 163.367
R827 B.n239 B.n238 163.367
R828 B.n239 B.n80 163.367
R829 B.n243 B.n80 163.367
R830 B.n244 B.n243 163.367
R831 B.n245 B.n244 163.367
R832 B.n245 B.n78 163.367
R833 B.n249 B.n78 163.367
R834 B.n250 B.n249 163.367
R835 B.n251 B.n250 163.367
R836 B.n251 B.n76 163.367
R837 B.n255 B.n76 163.367
R838 B.n256 B.n255 163.367
R839 B.n257 B.n256 163.367
R840 B.n257 B.n74 163.367
R841 B.n261 B.n74 163.367
R842 B.n262 B.n261 163.367
R843 B.n263 B.n262 163.367
R844 B.n263 B.n72 163.367
R845 B.n267 B.n72 163.367
R846 B.n268 B.n267 163.367
R847 B.n269 B.n70 163.367
R848 B.n273 B.n70 163.367
R849 B.n274 B.n273 163.367
R850 B.n275 B.n274 163.367
R851 B.n275 B.n68 163.367
R852 B.n279 B.n68 163.367
R853 B.n280 B.n279 163.367
R854 B.n281 B.n280 163.367
R855 B.n281 B.n66 163.367
R856 B.n285 B.n66 163.367
R857 B.n286 B.n285 163.367
R858 B.n287 B.n286 163.367
R859 B.n287 B.n64 163.367
R860 B.n291 B.n64 163.367
R861 B.n292 B.n291 163.367
R862 B.n293 B.n292 163.367
R863 B.n293 B.n62 163.367
R864 B.n297 B.n62 163.367
R865 B.n298 B.n297 163.367
R866 B.n299 B.n298 163.367
R867 B.n299 B.n60 163.367
R868 B.n303 B.n60 163.367
R869 B.n304 B.n303 163.367
R870 B.n305 B.n304 163.367
R871 B.n305 B.n58 163.367
R872 B.n309 B.n58 163.367
R873 B.n310 B.n309 163.367
R874 B.n311 B.n310 163.367
R875 B.n311 B.n56 163.367
R876 B.n315 B.n56 163.367
R877 B.n438 B.n437 163.367
R878 B.n437 B.n436 163.367
R879 B.n436 B.n11 163.367
R880 B.n432 B.n11 163.367
R881 B.n432 B.n431 163.367
R882 B.n431 B.n430 163.367
R883 B.n430 B.n13 163.367
R884 B.n426 B.n13 163.367
R885 B.n426 B.n425 163.367
R886 B.n425 B.n424 163.367
R887 B.n424 B.n15 163.367
R888 B.n420 B.n15 163.367
R889 B.n420 B.n419 163.367
R890 B.n419 B.n418 163.367
R891 B.n418 B.n17 163.367
R892 B.n414 B.n17 163.367
R893 B.n414 B.n413 163.367
R894 B.n413 B.n412 163.367
R895 B.n412 B.n19 163.367
R896 B.n408 B.n19 163.367
R897 B.n408 B.n407 163.367
R898 B.n407 B.n406 163.367
R899 B.n406 B.n21 163.367
R900 B.n402 B.n21 163.367
R901 B.n402 B.n401 163.367
R902 B.n401 B.n400 163.367
R903 B.n400 B.n23 163.367
R904 B.n396 B.n23 163.367
R905 B.n396 B.n395 163.367
R906 B.n395 B.n394 163.367
R907 B.n394 B.n25 163.367
R908 B.n390 B.n25 163.367
R909 B.n390 B.n389 163.367
R910 B.n389 B.n388 163.367
R911 B.n388 B.n27 163.367
R912 B.n383 B.n27 163.367
R913 B.n383 B.n382 163.367
R914 B.n382 B.n381 163.367
R915 B.n381 B.n31 163.367
R916 B.n377 B.n31 163.367
R917 B.n377 B.n376 163.367
R918 B.n376 B.n375 163.367
R919 B.n375 B.n33 163.367
R920 B.n371 B.n33 163.367
R921 B.n371 B.n370 163.367
R922 B.n370 B.n369 163.367
R923 B.n369 B.n35 163.367
R924 B.n365 B.n35 163.367
R925 B.n365 B.n364 163.367
R926 B.n364 B.n363 163.367
R927 B.n363 B.n40 163.367
R928 B.n359 B.n40 163.367
R929 B.n359 B.n358 163.367
R930 B.n358 B.n357 163.367
R931 B.n357 B.n42 163.367
R932 B.n353 B.n42 163.367
R933 B.n353 B.n352 163.367
R934 B.n352 B.n351 163.367
R935 B.n351 B.n44 163.367
R936 B.n347 B.n44 163.367
R937 B.n347 B.n346 163.367
R938 B.n346 B.n345 163.367
R939 B.n345 B.n46 163.367
R940 B.n341 B.n46 163.367
R941 B.n341 B.n340 163.367
R942 B.n340 B.n339 163.367
R943 B.n339 B.n48 163.367
R944 B.n335 B.n48 163.367
R945 B.n335 B.n334 163.367
R946 B.n334 B.n333 163.367
R947 B.n333 B.n50 163.367
R948 B.n329 B.n50 163.367
R949 B.n329 B.n328 163.367
R950 B.n328 B.n327 163.367
R951 B.n327 B.n52 163.367
R952 B.n323 B.n52 163.367
R953 B.n323 B.n322 163.367
R954 B.n322 B.n321 163.367
R955 B.n321 B.n54 163.367
R956 B.n317 B.n54 163.367
R957 B.n317 B.n316 163.367
R958 B.n91 B.n90 59.5399
R959 B.n199 B.n98 59.5399
R960 B.n385 B.n29 59.5399
R961 B.n38 B.n37 59.5399
R962 B.n440 B.n439 32.0005
R963 B.n314 B.n55 32.0005
R964 B.n270 B.n71 32.0005
R965 B.n145 B.n144 32.0005
R966 B.n90 B.n89 23.0793
R967 B.n98 B.n97 23.0793
R968 B.n29 B.n28 23.0793
R969 B.n37 B.n36 23.0793
R970 B B.n463 18.0485
R971 B.n439 B.n10 10.6151
R972 B.n435 B.n10 10.6151
R973 B.n435 B.n434 10.6151
R974 B.n434 B.n433 10.6151
R975 B.n433 B.n12 10.6151
R976 B.n429 B.n12 10.6151
R977 B.n429 B.n428 10.6151
R978 B.n428 B.n427 10.6151
R979 B.n427 B.n14 10.6151
R980 B.n423 B.n14 10.6151
R981 B.n423 B.n422 10.6151
R982 B.n422 B.n421 10.6151
R983 B.n421 B.n16 10.6151
R984 B.n417 B.n16 10.6151
R985 B.n417 B.n416 10.6151
R986 B.n416 B.n415 10.6151
R987 B.n415 B.n18 10.6151
R988 B.n411 B.n18 10.6151
R989 B.n411 B.n410 10.6151
R990 B.n410 B.n409 10.6151
R991 B.n409 B.n20 10.6151
R992 B.n405 B.n20 10.6151
R993 B.n405 B.n404 10.6151
R994 B.n404 B.n403 10.6151
R995 B.n403 B.n22 10.6151
R996 B.n399 B.n22 10.6151
R997 B.n399 B.n398 10.6151
R998 B.n398 B.n397 10.6151
R999 B.n397 B.n24 10.6151
R1000 B.n393 B.n24 10.6151
R1001 B.n393 B.n392 10.6151
R1002 B.n392 B.n391 10.6151
R1003 B.n391 B.n26 10.6151
R1004 B.n387 B.n26 10.6151
R1005 B.n387 B.n386 10.6151
R1006 B.n384 B.n30 10.6151
R1007 B.n380 B.n30 10.6151
R1008 B.n380 B.n379 10.6151
R1009 B.n379 B.n378 10.6151
R1010 B.n378 B.n32 10.6151
R1011 B.n374 B.n32 10.6151
R1012 B.n374 B.n373 10.6151
R1013 B.n373 B.n372 10.6151
R1014 B.n372 B.n34 10.6151
R1015 B.n368 B.n367 10.6151
R1016 B.n367 B.n366 10.6151
R1017 B.n366 B.n39 10.6151
R1018 B.n362 B.n39 10.6151
R1019 B.n362 B.n361 10.6151
R1020 B.n361 B.n360 10.6151
R1021 B.n360 B.n41 10.6151
R1022 B.n356 B.n41 10.6151
R1023 B.n356 B.n355 10.6151
R1024 B.n355 B.n354 10.6151
R1025 B.n354 B.n43 10.6151
R1026 B.n350 B.n43 10.6151
R1027 B.n350 B.n349 10.6151
R1028 B.n349 B.n348 10.6151
R1029 B.n348 B.n45 10.6151
R1030 B.n344 B.n45 10.6151
R1031 B.n344 B.n343 10.6151
R1032 B.n343 B.n342 10.6151
R1033 B.n342 B.n47 10.6151
R1034 B.n338 B.n47 10.6151
R1035 B.n338 B.n337 10.6151
R1036 B.n337 B.n336 10.6151
R1037 B.n336 B.n49 10.6151
R1038 B.n332 B.n49 10.6151
R1039 B.n332 B.n331 10.6151
R1040 B.n331 B.n330 10.6151
R1041 B.n330 B.n51 10.6151
R1042 B.n326 B.n51 10.6151
R1043 B.n326 B.n325 10.6151
R1044 B.n325 B.n324 10.6151
R1045 B.n324 B.n53 10.6151
R1046 B.n320 B.n53 10.6151
R1047 B.n320 B.n319 10.6151
R1048 B.n319 B.n318 10.6151
R1049 B.n318 B.n55 10.6151
R1050 B.n271 B.n270 10.6151
R1051 B.n272 B.n271 10.6151
R1052 B.n272 B.n69 10.6151
R1053 B.n276 B.n69 10.6151
R1054 B.n277 B.n276 10.6151
R1055 B.n278 B.n277 10.6151
R1056 B.n278 B.n67 10.6151
R1057 B.n282 B.n67 10.6151
R1058 B.n283 B.n282 10.6151
R1059 B.n284 B.n283 10.6151
R1060 B.n284 B.n65 10.6151
R1061 B.n288 B.n65 10.6151
R1062 B.n289 B.n288 10.6151
R1063 B.n290 B.n289 10.6151
R1064 B.n290 B.n63 10.6151
R1065 B.n294 B.n63 10.6151
R1066 B.n295 B.n294 10.6151
R1067 B.n296 B.n295 10.6151
R1068 B.n296 B.n61 10.6151
R1069 B.n300 B.n61 10.6151
R1070 B.n301 B.n300 10.6151
R1071 B.n302 B.n301 10.6151
R1072 B.n302 B.n59 10.6151
R1073 B.n306 B.n59 10.6151
R1074 B.n307 B.n306 10.6151
R1075 B.n308 B.n307 10.6151
R1076 B.n308 B.n57 10.6151
R1077 B.n312 B.n57 10.6151
R1078 B.n313 B.n312 10.6151
R1079 B.n314 B.n313 10.6151
R1080 B.n146 B.n145 10.6151
R1081 B.n146 B.n115 10.6151
R1082 B.n150 B.n115 10.6151
R1083 B.n151 B.n150 10.6151
R1084 B.n152 B.n151 10.6151
R1085 B.n152 B.n113 10.6151
R1086 B.n156 B.n113 10.6151
R1087 B.n157 B.n156 10.6151
R1088 B.n158 B.n157 10.6151
R1089 B.n158 B.n111 10.6151
R1090 B.n162 B.n111 10.6151
R1091 B.n163 B.n162 10.6151
R1092 B.n164 B.n163 10.6151
R1093 B.n164 B.n109 10.6151
R1094 B.n168 B.n109 10.6151
R1095 B.n169 B.n168 10.6151
R1096 B.n170 B.n169 10.6151
R1097 B.n170 B.n107 10.6151
R1098 B.n174 B.n107 10.6151
R1099 B.n175 B.n174 10.6151
R1100 B.n176 B.n175 10.6151
R1101 B.n176 B.n105 10.6151
R1102 B.n180 B.n105 10.6151
R1103 B.n181 B.n180 10.6151
R1104 B.n182 B.n181 10.6151
R1105 B.n182 B.n103 10.6151
R1106 B.n186 B.n103 10.6151
R1107 B.n187 B.n186 10.6151
R1108 B.n188 B.n187 10.6151
R1109 B.n188 B.n101 10.6151
R1110 B.n192 B.n101 10.6151
R1111 B.n193 B.n192 10.6151
R1112 B.n194 B.n193 10.6151
R1113 B.n194 B.n99 10.6151
R1114 B.n198 B.n99 10.6151
R1115 B.n201 B.n200 10.6151
R1116 B.n201 B.n95 10.6151
R1117 B.n205 B.n95 10.6151
R1118 B.n206 B.n205 10.6151
R1119 B.n207 B.n206 10.6151
R1120 B.n207 B.n93 10.6151
R1121 B.n211 B.n93 10.6151
R1122 B.n212 B.n211 10.6151
R1123 B.n213 B.n212 10.6151
R1124 B.n217 B.n216 10.6151
R1125 B.n218 B.n217 10.6151
R1126 B.n218 B.n87 10.6151
R1127 B.n222 B.n87 10.6151
R1128 B.n223 B.n222 10.6151
R1129 B.n224 B.n223 10.6151
R1130 B.n224 B.n85 10.6151
R1131 B.n228 B.n85 10.6151
R1132 B.n229 B.n228 10.6151
R1133 B.n230 B.n229 10.6151
R1134 B.n230 B.n83 10.6151
R1135 B.n234 B.n83 10.6151
R1136 B.n235 B.n234 10.6151
R1137 B.n236 B.n235 10.6151
R1138 B.n236 B.n81 10.6151
R1139 B.n240 B.n81 10.6151
R1140 B.n241 B.n240 10.6151
R1141 B.n242 B.n241 10.6151
R1142 B.n242 B.n79 10.6151
R1143 B.n246 B.n79 10.6151
R1144 B.n247 B.n246 10.6151
R1145 B.n248 B.n247 10.6151
R1146 B.n248 B.n77 10.6151
R1147 B.n252 B.n77 10.6151
R1148 B.n253 B.n252 10.6151
R1149 B.n254 B.n253 10.6151
R1150 B.n254 B.n75 10.6151
R1151 B.n258 B.n75 10.6151
R1152 B.n259 B.n258 10.6151
R1153 B.n260 B.n259 10.6151
R1154 B.n260 B.n73 10.6151
R1155 B.n264 B.n73 10.6151
R1156 B.n265 B.n264 10.6151
R1157 B.n266 B.n265 10.6151
R1158 B.n266 B.n71 10.6151
R1159 B.n144 B.n117 10.6151
R1160 B.n140 B.n117 10.6151
R1161 B.n140 B.n139 10.6151
R1162 B.n139 B.n138 10.6151
R1163 B.n138 B.n119 10.6151
R1164 B.n134 B.n119 10.6151
R1165 B.n134 B.n133 10.6151
R1166 B.n133 B.n132 10.6151
R1167 B.n132 B.n121 10.6151
R1168 B.n128 B.n121 10.6151
R1169 B.n128 B.n127 10.6151
R1170 B.n127 B.n126 10.6151
R1171 B.n126 B.n123 10.6151
R1172 B.n123 B.n0 10.6151
R1173 B.n459 B.n1 10.6151
R1174 B.n459 B.n458 10.6151
R1175 B.n458 B.n457 10.6151
R1176 B.n457 B.n4 10.6151
R1177 B.n453 B.n4 10.6151
R1178 B.n453 B.n452 10.6151
R1179 B.n452 B.n451 10.6151
R1180 B.n451 B.n6 10.6151
R1181 B.n447 B.n6 10.6151
R1182 B.n447 B.n446 10.6151
R1183 B.n446 B.n445 10.6151
R1184 B.n445 B.n8 10.6151
R1185 B.n441 B.n8 10.6151
R1186 B.n441 B.n440 10.6151
R1187 B.n386 B.n385 8.74196
R1188 B.n368 B.n38 8.74196
R1189 B.n199 B.n198 8.74196
R1190 B.n216 B.n91 8.74196
R1191 B.n463 B.n0 2.81026
R1192 B.n463 B.n1 2.81026
R1193 B.n385 B.n384 1.87367
R1194 B.n38 B.n34 1.87367
R1195 B.n200 B.n199 1.87367
R1196 B.n213 B.n91 1.87367
R1197 VN VN.t0 529.004
R1198 VN VN.t1 490.065
R1199 VDD2.n101 VDD2.n53 756.745
R1200 VDD2.n48 VDD2.n0 756.745
R1201 VDD2.n102 VDD2.n101 585
R1202 VDD2.n100 VDD2.n99 585
R1203 VDD2.n57 VDD2.n56 585
R1204 VDD2.n94 VDD2.n93 585
R1205 VDD2.n92 VDD2.n59 585
R1206 VDD2.n91 VDD2.n90 585
R1207 VDD2.n62 VDD2.n60 585
R1208 VDD2.n85 VDD2.n84 585
R1209 VDD2.n83 VDD2.n82 585
R1210 VDD2.n66 VDD2.n65 585
R1211 VDD2.n77 VDD2.n76 585
R1212 VDD2.n75 VDD2.n74 585
R1213 VDD2.n70 VDD2.n69 585
R1214 VDD2.n16 VDD2.n15 585
R1215 VDD2.n21 VDD2.n20 585
R1216 VDD2.n23 VDD2.n22 585
R1217 VDD2.n12 VDD2.n11 585
R1218 VDD2.n29 VDD2.n28 585
R1219 VDD2.n31 VDD2.n30 585
R1220 VDD2.n8 VDD2.n7 585
R1221 VDD2.n38 VDD2.n37 585
R1222 VDD2.n39 VDD2.n6 585
R1223 VDD2.n41 VDD2.n40 585
R1224 VDD2.n4 VDD2.n3 585
R1225 VDD2.n47 VDD2.n46 585
R1226 VDD2.n49 VDD2.n48 585
R1227 VDD2.n17 VDD2.t0 329.038
R1228 VDD2.n71 VDD2.t1 329.038
R1229 VDD2.n101 VDD2.n100 171.744
R1230 VDD2.n100 VDD2.n56 171.744
R1231 VDD2.n93 VDD2.n56 171.744
R1232 VDD2.n93 VDD2.n92 171.744
R1233 VDD2.n92 VDD2.n91 171.744
R1234 VDD2.n91 VDD2.n60 171.744
R1235 VDD2.n84 VDD2.n60 171.744
R1236 VDD2.n84 VDD2.n83 171.744
R1237 VDD2.n83 VDD2.n65 171.744
R1238 VDD2.n76 VDD2.n65 171.744
R1239 VDD2.n76 VDD2.n75 171.744
R1240 VDD2.n75 VDD2.n69 171.744
R1241 VDD2.n21 VDD2.n15 171.744
R1242 VDD2.n22 VDD2.n21 171.744
R1243 VDD2.n22 VDD2.n11 171.744
R1244 VDD2.n29 VDD2.n11 171.744
R1245 VDD2.n30 VDD2.n29 171.744
R1246 VDD2.n30 VDD2.n7 171.744
R1247 VDD2.n38 VDD2.n7 171.744
R1248 VDD2.n39 VDD2.n38 171.744
R1249 VDD2.n40 VDD2.n39 171.744
R1250 VDD2.n40 VDD2.n3 171.744
R1251 VDD2.n47 VDD2.n3 171.744
R1252 VDD2.n48 VDD2.n47 171.744
R1253 VDD2.t1 VDD2.n69 85.8723
R1254 VDD2.t0 VDD2.n15 85.8723
R1255 VDD2.n106 VDD2.n52 85.812
R1256 VDD2.n106 VDD2.n105 51.3853
R1257 VDD2.n94 VDD2.n59 13.1884
R1258 VDD2.n41 VDD2.n6 13.1884
R1259 VDD2.n95 VDD2.n57 12.8005
R1260 VDD2.n90 VDD2.n61 12.8005
R1261 VDD2.n37 VDD2.n36 12.8005
R1262 VDD2.n42 VDD2.n4 12.8005
R1263 VDD2.n99 VDD2.n98 12.0247
R1264 VDD2.n89 VDD2.n62 12.0247
R1265 VDD2.n35 VDD2.n8 12.0247
R1266 VDD2.n46 VDD2.n45 12.0247
R1267 VDD2.n102 VDD2.n55 11.249
R1268 VDD2.n86 VDD2.n85 11.249
R1269 VDD2.n32 VDD2.n31 11.249
R1270 VDD2.n49 VDD2.n2 11.249
R1271 VDD2.n71 VDD2.n70 10.7239
R1272 VDD2.n17 VDD2.n16 10.7239
R1273 VDD2.n103 VDD2.n53 10.4732
R1274 VDD2.n82 VDD2.n64 10.4732
R1275 VDD2.n28 VDD2.n10 10.4732
R1276 VDD2.n50 VDD2.n0 10.4732
R1277 VDD2.n81 VDD2.n66 9.69747
R1278 VDD2.n27 VDD2.n12 9.69747
R1279 VDD2.n105 VDD2.n104 9.45567
R1280 VDD2.n52 VDD2.n51 9.45567
R1281 VDD2.n73 VDD2.n72 9.3005
R1282 VDD2.n68 VDD2.n67 9.3005
R1283 VDD2.n79 VDD2.n78 9.3005
R1284 VDD2.n81 VDD2.n80 9.3005
R1285 VDD2.n64 VDD2.n63 9.3005
R1286 VDD2.n87 VDD2.n86 9.3005
R1287 VDD2.n89 VDD2.n88 9.3005
R1288 VDD2.n61 VDD2.n58 9.3005
R1289 VDD2.n104 VDD2.n103 9.3005
R1290 VDD2.n55 VDD2.n54 9.3005
R1291 VDD2.n98 VDD2.n97 9.3005
R1292 VDD2.n96 VDD2.n95 9.3005
R1293 VDD2.n51 VDD2.n50 9.3005
R1294 VDD2.n2 VDD2.n1 9.3005
R1295 VDD2.n45 VDD2.n44 9.3005
R1296 VDD2.n43 VDD2.n42 9.3005
R1297 VDD2.n19 VDD2.n18 9.3005
R1298 VDD2.n14 VDD2.n13 9.3005
R1299 VDD2.n25 VDD2.n24 9.3005
R1300 VDD2.n27 VDD2.n26 9.3005
R1301 VDD2.n10 VDD2.n9 9.3005
R1302 VDD2.n33 VDD2.n32 9.3005
R1303 VDD2.n35 VDD2.n34 9.3005
R1304 VDD2.n36 VDD2.n5 9.3005
R1305 VDD2.n78 VDD2.n77 8.92171
R1306 VDD2.n24 VDD2.n23 8.92171
R1307 VDD2.n74 VDD2.n68 8.14595
R1308 VDD2.n20 VDD2.n14 8.14595
R1309 VDD2.n73 VDD2.n70 7.3702
R1310 VDD2.n19 VDD2.n16 7.3702
R1311 VDD2.n74 VDD2.n73 5.81868
R1312 VDD2.n20 VDD2.n19 5.81868
R1313 VDD2.n77 VDD2.n68 5.04292
R1314 VDD2.n23 VDD2.n14 5.04292
R1315 VDD2.n78 VDD2.n66 4.26717
R1316 VDD2.n24 VDD2.n12 4.26717
R1317 VDD2.n105 VDD2.n53 3.49141
R1318 VDD2.n82 VDD2.n81 3.49141
R1319 VDD2.n28 VDD2.n27 3.49141
R1320 VDD2.n52 VDD2.n0 3.49141
R1321 VDD2.n103 VDD2.n102 2.71565
R1322 VDD2.n85 VDD2.n64 2.71565
R1323 VDD2.n31 VDD2.n10 2.71565
R1324 VDD2.n50 VDD2.n49 2.71565
R1325 VDD2.n72 VDD2.n71 2.41283
R1326 VDD2.n18 VDD2.n17 2.41283
R1327 VDD2.n99 VDD2.n55 1.93989
R1328 VDD2.n86 VDD2.n62 1.93989
R1329 VDD2.n32 VDD2.n8 1.93989
R1330 VDD2.n46 VDD2.n2 1.93989
R1331 VDD2.n98 VDD2.n57 1.16414
R1332 VDD2.n90 VDD2.n89 1.16414
R1333 VDD2.n37 VDD2.n35 1.16414
R1334 VDD2.n45 VDD2.n4 1.16414
R1335 VDD2.n95 VDD2.n94 0.388379
R1336 VDD2.n61 VDD2.n59 0.388379
R1337 VDD2.n36 VDD2.n6 0.388379
R1338 VDD2.n42 VDD2.n41 0.388379
R1339 VDD2 VDD2.n106 0.315155
R1340 VDD2.n104 VDD2.n54 0.155672
R1341 VDD2.n97 VDD2.n54 0.155672
R1342 VDD2.n97 VDD2.n96 0.155672
R1343 VDD2.n96 VDD2.n58 0.155672
R1344 VDD2.n88 VDD2.n58 0.155672
R1345 VDD2.n88 VDD2.n87 0.155672
R1346 VDD2.n87 VDD2.n63 0.155672
R1347 VDD2.n80 VDD2.n63 0.155672
R1348 VDD2.n80 VDD2.n79 0.155672
R1349 VDD2.n79 VDD2.n67 0.155672
R1350 VDD2.n72 VDD2.n67 0.155672
R1351 VDD2.n18 VDD2.n13 0.155672
R1352 VDD2.n25 VDD2.n13 0.155672
R1353 VDD2.n26 VDD2.n25 0.155672
R1354 VDD2.n26 VDD2.n9 0.155672
R1355 VDD2.n33 VDD2.n9 0.155672
R1356 VDD2.n34 VDD2.n33 0.155672
R1357 VDD2.n34 VDD2.n5 0.155672
R1358 VDD2.n43 VDD2.n5 0.155672
R1359 VDD2.n44 VDD2.n43 0.155672
R1360 VDD2.n44 VDD2.n1 0.155672
R1361 VDD2.n51 VDD2.n1 0.155672
C0 VP VDD1 1.93803f
C1 VDD2 w_n1446_n2990# 1.45552f
C2 VP VN 4.28033f
C3 VDD2 B 1.31913f
C4 VP w_n1446_n2990# 1.98906f
C5 VTAIL VDD1 4.774509f
C6 VP B 1.02225f
C7 VN VTAIL 1.43093f
C8 VN VDD1 0.148662f
C9 w_n1446_n2990# VTAIL 2.57821f
C10 VP VDD2 0.261373f
C11 VTAIL B 2.46359f
C12 w_n1446_n2990# VDD1 1.44925f
C13 VN w_n1446_n2990# 1.80862f
C14 B VDD1 1.3035f
C15 VN B 0.732579f
C16 VDD2 VTAIL 4.811f
C17 w_n1446_n2990# B 6.39755f
C18 VDD2 VDD1 0.477343f
C19 VP VTAIL 1.44542f
C20 VDD2 VN 1.8288f
C21 VDD2 VSUBS 0.680443f
C22 VDD1 VSUBS 2.370862f
C23 VTAIL VSUBS 0.708495f
C24 VN VSUBS 4.15455f
C25 VP VSUBS 1.075414f
C26 B VSUBS 2.452699f
C27 w_n1446_n2990# VSUBS 53.3921f
C28 VDD2.n0 VSUBS 0.01645f
C29 VDD2.n1 VSUBS 0.014971f
C30 VDD2.n2 VSUBS 0.008045f
C31 VDD2.n3 VSUBS 0.019015f
C32 VDD2.n4 VSUBS 0.008518f
C33 VDD2.n5 VSUBS 0.014971f
C34 VDD2.n6 VSUBS 0.008281f
C35 VDD2.n7 VSUBS 0.019015f
C36 VDD2.n8 VSUBS 0.008518f
C37 VDD2.n9 VSUBS 0.014971f
C38 VDD2.n10 VSUBS 0.008045f
C39 VDD2.n11 VSUBS 0.019015f
C40 VDD2.n12 VSUBS 0.008518f
C41 VDD2.n13 VSUBS 0.014971f
C42 VDD2.n14 VSUBS 0.008045f
C43 VDD2.n15 VSUBS 0.014261f
C44 VDD2.n16 VSUBS 0.014304f
C45 VDD2.t0 VSUBS 0.040892f
C46 VDD2.n17 VSUBS 0.104986f
C47 VDD2.n18 VSUBS 0.610242f
C48 VDD2.n19 VSUBS 0.008045f
C49 VDD2.n20 VSUBS 0.008518f
C50 VDD2.n21 VSUBS 0.019015f
C51 VDD2.n22 VSUBS 0.019015f
C52 VDD2.n23 VSUBS 0.008518f
C53 VDD2.n24 VSUBS 0.008045f
C54 VDD2.n25 VSUBS 0.014971f
C55 VDD2.n26 VSUBS 0.014971f
C56 VDD2.n27 VSUBS 0.008045f
C57 VDD2.n28 VSUBS 0.008518f
C58 VDD2.n29 VSUBS 0.019015f
C59 VDD2.n30 VSUBS 0.019015f
C60 VDD2.n31 VSUBS 0.008518f
C61 VDD2.n32 VSUBS 0.008045f
C62 VDD2.n33 VSUBS 0.014971f
C63 VDD2.n34 VSUBS 0.014971f
C64 VDD2.n35 VSUBS 0.008045f
C65 VDD2.n36 VSUBS 0.008045f
C66 VDD2.n37 VSUBS 0.008518f
C67 VDD2.n38 VSUBS 0.019015f
C68 VDD2.n39 VSUBS 0.019015f
C69 VDD2.n40 VSUBS 0.019015f
C70 VDD2.n41 VSUBS 0.008281f
C71 VDD2.n42 VSUBS 0.008045f
C72 VDD2.n43 VSUBS 0.014971f
C73 VDD2.n44 VSUBS 0.014971f
C74 VDD2.n45 VSUBS 0.008045f
C75 VDD2.n46 VSUBS 0.008518f
C76 VDD2.n47 VSUBS 0.019015f
C77 VDD2.n48 VSUBS 0.046035f
C78 VDD2.n49 VSUBS 0.008518f
C79 VDD2.n50 VSUBS 0.008045f
C80 VDD2.n51 VSUBS 0.037263f
C81 VDD2.n52 VSUBS 0.328163f
C82 VDD2.n53 VSUBS 0.01645f
C83 VDD2.n54 VSUBS 0.014971f
C84 VDD2.n55 VSUBS 0.008045f
C85 VDD2.n56 VSUBS 0.019015f
C86 VDD2.n57 VSUBS 0.008518f
C87 VDD2.n58 VSUBS 0.014971f
C88 VDD2.n59 VSUBS 0.008281f
C89 VDD2.n60 VSUBS 0.019015f
C90 VDD2.n61 VSUBS 0.008045f
C91 VDD2.n62 VSUBS 0.008518f
C92 VDD2.n63 VSUBS 0.014971f
C93 VDD2.n64 VSUBS 0.008045f
C94 VDD2.n65 VSUBS 0.019015f
C95 VDD2.n66 VSUBS 0.008518f
C96 VDD2.n67 VSUBS 0.014971f
C97 VDD2.n68 VSUBS 0.008045f
C98 VDD2.n69 VSUBS 0.014261f
C99 VDD2.n70 VSUBS 0.014304f
C100 VDD2.t1 VSUBS 0.040892f
C101 VDD2.n71 VSUBS 0.104986f
C102 VDD2.n72 VSUBS 0.610242f
C103 VDD2.n73 VSUBS 0.008045f
C104 VDD2.n74 VSUBS 0.008518f
C105 VDD2.n75 VSUBS 0.019015f
C106 VDD2.n76 VSUBS 0.019015f
C107 VDD2.n77 VSUBS 0.008518f
C108 VDD2.n78 VSUBS 0.008045f
C109 VDD2.n79 VSUBS 0.014971f
C110 VDD2.n80 VSUBS 0.014971f
C111 VDD2.n81 VSUBS 0.008045f
C112 VDD2.n82 VSUBS 0.008518f
C113 VDD2.n83 VSUBS 0.019015f
C114 VDD2.n84 VSUBS 0.019015f
C115 VDD2.n85 VSUBS 0.008518f
C116 VDD2.n86 VSUBS 0.008045f
C117 VDD2.n87 VSUBS 0.014971f
C118 VDD2.n88 VSUBS 0.014971f
C119 VDD2.n89 VSUBS 0.008045f
C120 VDD2.n90 VSUBS 0.008518f
C121 VDD2.n91 VSUBS 0.019015f
C122 VDD2.n92 VSUBS 0.019015f
C123 VDD2.n93 VSUBS 0.019015f
C124 VDD2.n94 VSUBS 0.008281f
C125 VDD2.n95 VSUBS 0.008045f
C126 VDD2.n96 VSUBS 0.014971f
C127 VDD2.n97 VSUBS 0.014971f
C128 VDD2.n98 VSUBS 0.008045f
C129 VDD2.n99 VSUBS 0.008518f
C130 VDD2.n100 VSUBS 0.019015f
C131 VDD2.n101 VSUBS 0.046035f
C132 VDD2.n102 VSUBS 0.008518f
C133 VDD2.n103 VSUBS 0.008045f
C134 VDD2.n104 VSUBS 0.037263f
C135 VDD2.n105 VSUBS 0.033547f
C136 VDD2.n106 VSUBS 1.5148f
C137 VN.t1 VSUBS 0.840527f
C138 VN.t0 VSUBS 0.935888f
C139 B.n0 VSUBS 0.004786f
C140 B.n1 VSUBS 0.004786f
C141 B.n2 VSUBS 0.007569f
C142 B.n3 VSUBS 0.007569f
C143 B.n4 VSUBS 0.007569f
C144 B.n5 VSUBS 0.007569f
C145 B.n6 VSUBS 0.007569f
C146 B.n7 VSUBS 0.007569f
C147 B.n8 VSUBS 0.007569f
C148 B.n9 VSUBS 0.016841f
C149 B.n10 VSUBS 0.007569f
C150 B.n11 VSUBS 0.007569f
C151 B.n12 VSUBS 0.007569f
C152 B.n13 VSUBS 0.007569f
C153 B.n14 VSUBS 0.007569f
C154 B.n15 VSUBS 0.007569f
C155 B.n16 VSUBS 0.007569f
C156 B.n17 VSUBS 0.007569f
C157 B.n18 VSUBS 0.007569f
C158 B.n19 VSUBS 0.007569f
C159 B.n20 VSUBS 0.007569f
C160 B.n21 VSUBS 0.007569f
C161 B.n22 VSUBS 0.007569f
C162 B.n23 VSUBS 0.007569f
C163 B.n24 VSUBS 0.007569f
C164 B.n25 VSUBS 0.007569f
C165 B.n26 VSUBS 0.007569f
C166 B.n27 VSUBS 0.007569f
C167 B.t2 VSUBS 0.183323f
C168 B.t1 VSUBS 0.197503f
C169 B.t0 VSUBS 0.39742f
C170 B.n28 VSUBS 0.300015f
C171 B.n29 VSUBS 0.234689f
C172 B.n30 VSUBS 0.007569f
C173 B.n31 VSUBS 0.007569f
C174 B.n32 VSUBS 0.007569f
C175 B.n33 VSUBS 0.007569f
C176 B.n34 VSUBS 0.004452f
C177 B.n35 VSUBS 0.007569f
C178 B.t5 VSUBS 0.183325f
C179 B.t4 VSUBS 0.197505f
C180 B.t3 VSUBS 0.39742f
C181 B.n36 VSUBS 0.300012f
C182 B.n37 VSUBS 0.234686f
C183 B.n38 VSUBS 0.017536f
C184 B.n39 VSUBS 0.007569f
C185 B.n40 VSUBS 0.007569f
C186 B.n41 VSUBS 0.007569f
C187 B.n42 VSUBS 0.007569f
C188 B.n43 VSUBS 0.007569f
C189 B.n44 VSUBS 0.007569f
C190 B.n45 VSUBS 0.007569f
C191 B.n46 VSUBS 0.007569f
C192 B.n47 VSUBS 0.007569f
C193 B.n48 VSUBS 0.007569f
C194 B.n49 VSUBS 0.007569f
C195 B.n50 VSUBS 0.007569f
C196 B.n51 VSUBS 0.007569f
C197 B.n52 VSUBS 0.007569f
C198 B.n53 VSUBS 0.007569f
C199 B.n54 VSUBS 0.007569f
C200 B.n55 VSUBS 0.017197f
C201 B.n56 VSUBS 0.007569f
C202 B.n57 VSUBS 0.007569f
C203 B.n58 VSUBS 0.007569f
C204 B.n59 VSUBS 0.007569f
C205 B.n60 VSUBS 0.007569f
C206 B.n61 VSUBS 0.007569f
C207 B.n62 VSUBS 0.007569f
C208 B.n63 VSUBS 0.007569f
C209 B.n64 VSUBS 0.007569f
C210 B.n65 VSUBS 0.007569f
C211 B.n66 VSUBS 0.007569f
C212 B.n67 VSUBS 0.007569f
C213 B.n68 VSUBS 0.007569f
C214 B.n69 VSUBS 0.007569f
C215 B.n70 VSUBS 0.007569f
C216 B.n71 VSUBS 0.01811f
C217 B.n72 VSUBS 0.007569f
C218 B.n73 VSUBS 0.007569f
C219 B.n74 VSUBS 0.007569f
C220 B.n75 VSUBS 0.007569f
C221 B.n76 VSUBS 0.007569f
C222 B.n77 VSUBS 0.007569f
C223 B.n78 VSUBS 0.007569f
C224 B.n79 VSUBS 0.007569f
C225 B.n80 VSUBS 0.007569f
C226 B.n81 VSUBS 0.007569f
C227 B.n82 VSUBS 0.007569f
C228 B.n83 VSUBS 0.007569f
C229 B.n84 VSUBS 0.007569f
C230 B.n85 VSUBS 0.007569f
C231 B.n86 VSUBS 0.007569f
C232 B.n87 VSUBS 0.007569f
C233 B.n88 VSUBS 0.007569f
C234 B.t10 VSUBS 0.183325f
C235 B.t11 VSUBS 0.197505f
C236 B.t9 VSUBS 0.39742f
C237 B.n89 VSUBS 0.300012f
C238 B.n90 VSUBS 0.234686f
C239 B.n91 VSUBS 0.017536f
C240 B.n92 VSUBS 0.007569f
C241 B.n93 VSUBS 0.007569f
C242 B.n94 VSUBS 0.007569f
C243 B.n95 VSUBS 0.007569f
C244 B.n96 VSUBS 0.007569f
C245 B.t7 VSUBS 0.183323f
C246 B.t8 VSUBS 0.197503f
C247 B.t6 VSUBS 0.39742f
C248 B.n97 VSUBS 0.300015f
C249 B.n98 VSUBS 0.234689f
C250 B.n99 VSUBS 0.007569f
C251 B.n100 VSUBS 0.007569f
C252 B.n101 VSUBS 0.007569f
C253 B.n102 VSUBS 0.007569f
C254 B.n103 VSUBS 0.007569f
C255 B.n104 VSUBS 0.007569f
C256 B.n105 VSUBS 0.007569f
C257 B.n106 VSUBS 0.007569f
C258 B.n107 VSUBS 0.007569f
C259 B.n108 VSUBS 0.007569f
C260 B.n109 VSUBS 0.007569f
C261 B.n110 VSUBS 0.007569f
C262 B.n111 VSUBS 0.007569f
C263 B.n112 VSUBS 0.007569f
C264 B.n113 VSUBS 0.007569f
C265 B.n114 VSUBS 0.007569f
C266 B.n115 VSUBS 0.007569f
C267 B.n116 VSUBS 0.01811f
C268 B.n117 VSUBS 0.007569f
C269 B.n118 VSUBS 0.007569f
C270 B.n119 VSUBS 0.007569f
C271 B.n120 VSUBS 0.007569f
C272 B.n121 VSUBS 0.007569f
C273 B.n122 VSUBS 0.007569f
C274 B.n123 VSUBS 0.007569f
C275 B.n124 VSUBS 0.007569f
C276 B.n125 VSUBS 0.007569f
C277 B.n126 VSUBS 0.007569f
C278 B.n127 VSUBS 0.007569f
C279 B.n128 VSUBS 0.007569f
C280 B.n129 VSUBS 0.007569f
C281 B.n130 VSUBS 0.007569f
C282 B.n131 VSUBS 0.007569f
C283 B.n132 VSUBS 0.007569f
C284 B.n133 VSUBS 0.007569f
C285 B.n134 VSUBS 0.007569f
C286 B.n135 VSUBS 0.007569f
C287 B.n136 VSUBS 0.007569f
C288 B.n137 VSUBS 0.007569f
C289 B.n138 VSUBS 0.007569f
C290 B.n139 VSUBS 0.007569f
C291 B.n140 VSUBS 0.007569f
C292 B.n141 VSUBS 0.007569f
C293 B.n142 VSUBS 0.007569f
C294 B.n143 VSUBS 0.016841f
C295 B.n144 VSUBS 0.016841f
C296 B.n145 VSUBS 0.01811f
C297 B.n146 VSUBS 0.007569f
C298 B.n147 VSUBS 0.007569f
C299 B.n148 VSUBS 0.007569f
C300 B.n149 VSUBS 0.007569f
C301 B.n150 VSUBS 0.007569f
C302 B.n151 VSUBS 0.007569f
C303 B.n152 VSUBS 0.007569f
C304 B.n153 VSUBS 0.007569f
C305 B.n154 VSUBS 0.007569f
C306 B.n155 VSUBS 0.007569f
C307 B.n156 VSUBS 0.007569f
C308 B.n157 VSUBS 0.007569f
C309 B.n158 VSUBS 0.007569f
C310 B.n159 VSUBS 0.007569f
C311 B.n160 VSUBS 0.007569f
C312 B.n161 VSUBS 0.007569f
C313 B.n162 VSUBS 0.007569f
C314 B.n163 VSUBS 0.007569f
C315 B.n164 VSUBS 0.007569f
C316 B.n165 VSUBS 0.007569f
C317 B.n166 VSUBS 0.007569f
C318 B.n167 VSUBS 0.007569f
C319 B.n168 VSUBS 0.007569f
C320 B.n169 VSUBS 0.007569f
C321 B.n170 VSUBS 0.007569f
C322 B.n171 VSUBS 0.007569f
C323 B.n172 VSUBS 0.007569f
C324 B.n173 VSUBS 0.007569f
C325 B.n174 VSUBS 0.007569f
C326 B.n175 VSUBS 0.007569f
C327 B.n176 VSUBS 0.007569f
C328 B.n177 VSUBS 0.007569f
C329 B.n178 VSUBS 0.007569f
C330 B.n179 VSUBS 0.007569f
C331 B.n180 VSUBS 0.007569f
C332 B.n181 VSUBS 0.007569f
C333 B.n182 VSUBS 0.007569f
C334 B.n183 VSUBS 0.007569f
C335 B.n184 VSUBS 0.007569f
C336 B.n185 VSUBS 0.007569f
C337 B.n186 VSUBS 0.007569f
C338 B.n187 VSUBS 0.007569f
C339 B.n188 VSUBS 0.007569f
C340 B.n189 VSUBS 0.007569f
C341 B.n190 VSUBS 0.007569f
C342 B.n191 VSUBS 0.007569f
C343 B.n192 VSUBS 0.007569f
C344 B.n193 VSUBS 0.007569f
C345 B.n194 VSUBS 0.007569f
C346 B.n195 VSUBS 0.007569f
C347 B.n196 VSUBS 0.007569f
C348 B.n197 VSUBS 0.007569f
C349 B.n198 VSUBS 0.006901f
C350 B.n199 VSUBS 0.017536f
C351 B.n200 VSUBS 0.004452f
C352 B.n201 VSUBS 0.007569f
C353 B.n202 VSUBS 0.007569f
C354 B.n203 VSUBS 0.007569f
C355 B.n204 VSUBS 0.007569f
C356 B.n205 VSUBS 0.007569f
C357 B.n206 VSUBS 0.007569f
C358 B.n207 VSUBS 0.007569f
C359 B.n208 VSUBS 0.007569f
C360 B.n209 VSUBS 0.007569f
C361 B.n210 VSUBS 0.007569f
C362 B.n211 VSUBS 0.007569f
C363 B.n212 VSUBS 0.007569f
C364 B.n213 VSUBS 0.004452f
C365 B.n214 VSUBS 0.007569f
C366 B.n215 VSUBS 0.007569f
C367 B.n216 VSUBS 0.006901f
C368 B.n217 VSUBS 0.007569f
C369 B.n218 VSUBS 0.007569f
C370 B.n219 VSUBS 0.007569f
C371 B.n220 VSUBS 0.007569f
C372 B.n221 VSUBS 0.007569f
C373 B.n222 VSUBS 0.007569f
C374 B.n223 VSUBS 0.007569f
C375 B.n224 VSUBS 0.007569f
C376 B.n225 VSUBS 0.007569f
C377 B.n226 VSUBS 0.007569f
C378 B.n227 VSUBS 0.007569f
C379 B.n228 VSUBS 0.007569f
C380 B.n229 VSUBS 0.007569f
C381 B.n230 VSUBS 0.007569f
C382 B.n231 VSUBS 0.007569f
C383 B.n232 VSUBS 0.007569f
C384 B.n233 VSUBS 0.007569f
C385 B.n234 VSUBS 0.007569f
C386 B.n235 VSUBS 0.007569f
C387 B.n236 VSUBS 0.007569f
C388 B.n237 VSUBS 0.007569f
C389 B.n238 VSUBS 0.007569f
C390 B.n239 VSUBS 0.007569f
C391 B.n240 VSUBS 0.007569f
C392 B.n241 VSUBS 0.007569f
C393 B.n242 VSUBS 0.007569f
C394 B.n243 VSUBS 0.007569f
C395 B.n244 VSUBS 0.007569f
C396 B.n245 VSUBS 0.007569f
C397 B.n246 VSUBS 0.007569f
C398 B.n247 VSUBS 0.007569f
C399 B.n248 VSUBS 0.007569f
C400 B.n249 VSUBS 0.007569f
C401 B.n250 VSUBS 0.007569f
C402 B.n251 VSUBS 0.007569f
C403 B.n252 VSUBS 0.007569f
C404 B.n253 VSUBS 0.007569f
C405 B.n254 VSUBS 0.007569f
C406 B.n255 VSUBS 0.007569f
C407 B.n256 VSUBS 0.007569f
C408 B.n257 VSUBS 0.007569f
C409 B.n258 VSUBS 0.007569f
C410 B.n259 VSUBS 0.007569f
C411 B.n260 VSUBS 0.007569f
C412 B.n261 VSUBS 0.007569f
C413 B.n262 VSUBS 0.007569f
C414 B.n263 VSUBS 0.007569f
C415 B.n264 VSUBS 0.007569f
C416 B.n265 VSUBS 0.007569f
C417 B.n266 VSUBS 0.007569f
C418 B.n267 VSUBS 0.007569f
C419 B.n268 VSUBS 0.01811f
C420 B.n269 VSUBS 0.016841f
C421 B.n270 VSUBS 0.016841f
C422 B.n271 VSUBS 0.007569f
C423 B.n272 VSUBS 0.007569f
C424 B.n273 VSUBS 0.007569f
C425 B.n274 VSUBS 0.007569f
C426 B.n275 VSUBS 0.007569f
C427 B.n276 VSUBS 0.007569f
C428 B.n277 VSUBS 0.007569f
C429 B.n278 VSUBS 0.007569f
C430 B.n279 VSUBS 0.007569f
C431 B.n280 VSUBS 0.007569f
C432 B.n281 VSUBS 0.007569f
C433 B.n282 VSUBS 0.007569f
C434 B.n283 VSUBS 0.007569f
C435 B.n284 VSUBS 0.007569f
C436 B.n285 VSUBS 0.007569f
C437 B.n286 VSUBS 0.007569f
C438 B.n287 VSUBS 0.007569f
C439 B.n288 VSUBS 0.007569f
C440 B.n289 VSUBS 0.007569f
C441 B.n290 VSUBS 0.007569f
C442 B.n291 VSUBS 0.007569f
C443 B.n292 VSUBS 0.007569f
C444 B.n293 VSUBS 0.007569f
C445 B.n294 VSUBS 0.007569f
C446 B.n295 VSUBS 0.007569f
C447 B.n296 VSUBS 0.007569f
C448 B.n297 VSUBS 0.007569f
C449 B.n298 VSUBS 0.007569f
C450 B.n299 VSUBS 0.007569f
C451 B.n300 VSUBS 0.007569f
C452 B.n301 VSUBS 0.007569f
C453 B.n302 VSUBS 0.007569f
C454 B.n303 VSUBS 0.007569f
C455 B.n304 VSUBS 0.007569f
C456 B.n305 VSUBS 0.007569f
C457 B.n306 VSUBS 0.007569f
C458 B.n307 VSUBS 0.007569f
C459 B.n308 VSUBS 0.007569f
C460 B.n309 VSUBS 0.007569f
C461 B.n310 VSUBS 0.007569f
C462 B.n311 VSUBS 0.007569f
C463 B.n312 VSUBS 0.007569f
C464 B.n313 VSUBS 0.007569f
C465 B.n314 VSUBS 0.017753f
C466 B.n315 VSUBS 0.016841f
C467 B.n316 VSUBS 0.01811f
C468 B.n317 VSUBS 0.007569f
C469 B.n318 VSUBS 0.007569f
C470 B.n319 VSUBS 0.007569f
C471 B.n320 VSUBS 0.007569f
C472 B.n321 VSUBS 0.007569f
C473 B.n322 VSUBS 0.007569f
C474 B.n323 VSUBS 0.007569f
C475 B.n324 VSUBS 0.007569f
C476 B.n325 VSUBS 0.007569f
C477 B.n326 VSUBS 0.007569f
C478 B.n327 VSUBS 0.007569f
C479 B.n328 VSUBS 0.007569f
C480 B.n329 VSUBS 0.007569f
C481 B.n330 VSUBS 0.007569f
C482 B.n331 VSUBS 0.007569f
C483 B.n332 VSUBS 0.007569f
C484 B.n333 VSUBS 0.007569f
C485 B.n334 VSUBS 0.007569f
C486 B.n335 VSUBS 0.007569f
C487 B.n336 VSUBS 0.007569f
C488 B.n337 VSUBS 0.007569f
C489 B.n338 VSUBS 0.007569f
C490 B.n339 VSUBS 0.007569f
C491 B.n340 VSUBS 0.007569f
C492 B.n341 VSUBS 0.007569f
C493 B.n342 VSUBS 0.007569f
C494 B.n343 VSUBS 0.007569f
C495 B.n344 VSUBS 0.007569f
C496 B.n345 VSUBS 0.007569f
C497 B.n346 VSUBS 0.007569f
C498 B.n347 VSUBS 0.007569f
C499 B.n348 VSUBS 0.007569f
C500 B.n349 VSUBS 0.007569f
C501 B.n350 VSUBS 0.007569f
C502 B.n351 VSUBS 0.007569f
C503 B.n352 VSUBS 0.007569f
C504 B.n353 VSUBS 0.007569f
C505 B.n354 VSUBS 0.007569f
C506 B.n355 VSUBS 0.007569f
C507 B.n356 VSUBS 0.007569f
C508 B.n357 VSUBS 0.007569f
C509 B.n358 VSUBS 0.007569f
C510 B.n359 VSUBS 0.007569f
C511 B.n360 VSUBS 0.007569f
C512 B.n361 VSUBS 0.007569f
C513 B.n362 VSUBS 0.007569f
C514 B.n363 VSUBS 0.007569f
C515 B.n364 VSUBS 0.007569f
C516 B.n365 VSUBS 0.007569f
C517 B.n366 VSUBS 0.007569f
C518 B.n367 VSUBS 0.007569f
C519 B.n368 VSUBS 0.006901f
C520 B.n369 VSUBS 0.007569f
C521 B.n370 VSUBS 0.007569f
C522 B.n371 VSUBS 0.007569f
C523 B.n372 VSUBS 0.007569f
C524 B.n373 VSUBS 0.007569f
C525 B.n374 VSUBS 0.007569f
C526 B.n375 VSUBS 0.007569f
C527 B.n376 VSUBS 0.007569f
C528 B.n377 VSUBS 0.007569f
C529 B.n378 VSUBS 0.007569f
C530 B.n379 VSUBS 0.007569f
C531 B.n380 VSUBS 0.007569f
C532 B.n381 VSUBS 0.007569f
C533 B.n382 VSUBS 0.007569f
C534 B.n383 VSUBS 0.007569f
C535 B.n384 VSUBS 0.004452f
C536 B.n385 VSUBS 0.017536f
C537 B.n386 VSUBS 0.006901f
C538 B.n387 VSUBS 0.007569f
C539 B.n388 VSUBS 0.007569f
C540 B.n389 VSUBS 0.007569f
C541 B.n390 VSUBS 0.007569f
C542 B.n391 VSUBS 0.007569f
C543 B.n392 VSUBS 0.007569f
C544 B.n393 VSUBS 0.007569f
C545 B.n394 VSUBS 0.007569f
C546 B.n395 VSUBS 0.007569f
C547 B.n396 VSUBS 0.007569f
C548 B.n397 VSUBS 0.007569f
C549 B.n398 VSUBS 0.007569f
C550 B.n399 VSUBS 0.007569f
C551 B.n400 VSUBS 0.007569f
C552 B.n401 VSUBS 0.007569f
C553 B.n402 VSUBS 0.007569f
C554 B.n403 VSUBS 0.007569f
C555 B.n404 VSUBS 0.007569f
C556 B.n405 VSUBS 0.007569f
C557 B.n406 VSUBS 0.007569f
C558 B.n407 VSUBS 0.007569f
C559 B.n408 VSUBS 0.007569f
C560 B.n409 VSUBS 0.007569f
C561 B.n410 VSUBS 0.007569f
C562 B.n411 VSUBS 0.007569f
C563 B.n412 VSUBS 0.007569f
C564 B.n413 VSUBS 0.007569f
C565 B.n414 VSUBS 0.007569f
C566 B.n415 VSUBS 0.007569f
C567 B.n416 VSUBS 0.007569f
C568 B.n417 VSUBS 0.007569f
C569 B.n418 VSUBS 0.007569f
C570 B.n419 VSUBS 0.007569f
C571 B.n420 VSUBS 0.007569f
C572 B.n421 VSUBS 0.007569f
C573 B.n422 VSUBS 0.007569f
C574 B.n423 VSUBS 0.007569f
C575 B.n424 VSUBS 0.007569f
C576 B.n425 VSUBS 0.007569f
C577 B.n426 VSUBS 0.007569f
C578 B.n427 VSUBS 0.007569f
C579 B.n428 VSUBS 0.007569f
C580 B.n429 VSUBS 0.007569f
C581 B.n430 VSUBS 0.007569f
C582 B.n431 VSUBS 0.007569f
C583 B.n432 VSUBS 0.007569f
C584 B.n433 VSUBS 0.007569f
C585 B.n434 VSUBS 0.007569f
C586 B.n435 VSUBS 0.007569f
C587 B.n436 VSUBS 0.007569f
C588 B.n437 VSUBS 0.007569f
C589 B.n438 VSUBS 0.01811f
C590 B.n439 VSUBS 0.01811f
C591 B.n440 VSUBS 0.016841f
C592 B.n441 VSUBS 0.007569f
C593 B.n442 VSUBS 0.007569f
C594 B.n443 VSUBS 0.007569f
C595 B.n444 VSUBS 0.007569f
C596 B.n445 VSUBS 0.007569f
C597 B.n446 VSUBS 0.007569f
C598 B.n447 VSUBS 0.007569f
C599 B.n448 VSUBS 0.007569f
C600 B.n449 VSUBS 0.007569f
C601 B.n450 VSUBS 0.007569f
C602 B.n451 VSUBS 0.007569f
C603 B.n452 VSUBS 0.007569f
C604 B.n453 VSUBS 0.007569f
C605 B.n454 VSUBS 0.007569f
C606 B.n455 VSUBS 0.007569f
C607 B.n456 VSUBS 0.007569f
C608 B.n457 VSUBS 0.007569f
C609 B.n458 VSUBS 0.007569f
C610 B.n459 VSUBS 0.007569f
C611 B.n460 VSUBS 0.007569f
C612 B.n461 VSUBS 0.007569f
C613 B.n462 VSUBS 0.007569f
C614 B.n463 VSUBS 0.017138f
C615 VDD1.n0 VSUBS 0.016263f
C616 VDD1.n1 VSUBS 0.0148f
C617 VDD1.n2 VSUBS 0.007953f
C618 VDD1.n3 VSUBS 0.018798f
C619 VDD1.n4 VSUBS 0.008421f
C620 VDD1.n5 VSUBS 0.0148f
C621 VDD1.n6 VSUBS 0.008187f
C622 VDD1.n7 VSUBS 0.018798f
C623 VDD1.n8 VSUBS 0.007953f
C624 VDD1.n9 VSUBS 0.008421f
C625 VDD1.n10 VSUBS 0.0148f
C626 VDD1.n11 VSUBS 0.007953f
C627 VDD1.n12 VSUBS 0.018798f
C628 VDD1.n13 VSUBS 0.008421f
C629 VDD1.n14 VSUBS 0.0148f
C630 VDD1.n15 VSUBS 0.007953f
C631 VDD1.n16 VSUBS 0.014098f
C632 VDD1.n17 VSUBS 0.014141f
C633 VDD1.t1 VSUBS 0.040426f
C634 VDD1.n18 VSUBS 0.10379f
C635 VDD1.n19 VSUBS 0.603292f
C636 VDD1.n20 VSUBS 0.007953f
C637 VDD1.n21 VSUBS 0.008421f
C638 VDD1.n22 VSUBS 0.018798f
C639 VDD1.n23 VSUBS 0.018798f
C640 VDD1.n24 VSUBS 0.008421f
C641 VDD1.n25 VSUBS 0.007953f
C642 VDD1.n26 VSUBS 0.0148f
C643 VDD1.n27 VSUBS 0.0148f
C644 VDD1.n28 VSUBS 0.007953f
C645 VDD1.n29 VSUBS 0.008421f
C646 VDD1.n30 VSUBS 0.018798f
C647 VDD1.n31 VSUBS 0.018798f
C648 VDD1.n32 VSUBS 0.008421f
C649 VDD1.n33 VSUBS 0.007953f
C650 VDD1.n34 VSUBS 0.0148f
C651 VDD1.n35 VSUBS 0.0148f
C652 VDD1.n36 VSUBS 0.007953f
C653 VDD1.n37 VSUBS 0.008421f
C654 VDD1.n38 VSUBS 0.018798f
C655 VDD1.n39 VSUBS 0.018798f
C656 VDD1.n40 VSUBS 0.018798f
C657 VDD1.n41 VSUBS 0.008187f
C658 VDD1.n42 VSUBS 0.007953f
C659 VDD1.n43 VSUBS 0.0148f
C660 VDD1.n44 VSUBS 0.0148f
C661 VDD1.n45 VSUBS 0.007953f
C662 VDD1.n46 VSUBS 0.008421f
C663 VDD1.n47 VSUBS 0.018798f
C664 VDD1.n48 VSUBS 0.045511f
C665 VDD1.n49 VSUBS 0.008421f
C666 VDD1.n50 VSUBS 0.007953f
C667 VDD1.n51 VSUBS 0.036838f
C668 VDD1.n52 VSUBS 0.033439f
C669 VDD1.n53 VSUBS 0.016263f
C670 VDD1.n54 VSUBS 0.0148f
C671 VDD1.n55 VSUBS 0.007953f
C672 VDD1.n56 VSUBS 0.018798f
C673 VDD1.n57 VSUBS 0.008421f
C674 VDD1.n58 VSUBS 0.0148f
C675 VDD1.n59 VSUBS 0.008187f
C676 VDD1.n60 VSUBS 0.018798f
C677 VDD1.n61 VSUBS 0.008421f
C678 VDD1.n62 VSUBS 0.0148f
C679 VDD1.n63 VSUBS 0.007953f
C680 VDD1.n64 VSUBS 0.018798f
C681 VDD1.n65 VSUBS 0.008421f
C682 VDD1.n66 VSUBS 0.0148f
C683 VDD1.n67 VSUBS 0.007953f
C684 VDD1.n68 VSUBS 0.014098f
C685 VDD1.n69 VSUBS 0.014141f
C686 VDD1.t0 VSUBS 0.040426f
C687 VDD1.n70 VSUBS 0.10379f
C688 VDD1.n71 VSUBS 0.603292f
C689 VDD1.n72 VSUBS 0.007953f
C690 VDD1.n73 VSUBS 0.008421f
C691 VDD1.n74 VSUBS 0.018798f
C692 VDD1.n75 VSUBS 0.018798f
C693 VDD1.n76 VSUBS 0.008421f
C694 VDD1.n77 VSUBS 0.007953f
C695 VDD1.n78 VSUBS 0.0148f
C696 VDD1.n79 VSUBS 0.0148f
C697 VDD1.n80 VSUBS 0.007953f
C698 VDD1.n81 VSUBS 0.008421f
C699 VDD1.n82 VSUBS 0.018798f
C700 VDD1.n83 VSUBS 0.018798f
C701 VDD1.n84 VSUBS 0.008421f
C702 VDD1.n85 VSUBS 0.007953f
C703 VDD1.n86 VSUBS 0.0148f
C704 VDD1.n87 VSUBS 0.0148f
C705 VDD1.n88 VSUBS 0.007953f
C706 VDD1.n89 VSUBS 0.007953f
C707 VDD1.n90 VSUBS 0.008421f
C708 VDD1.n91 VSUBS 0.018798f
C709 VDD1.n92 VSUBS 0.018798f
C710 VDD1.n93 VSUBS 0.018798f
C711 VDD1.n94 VSUBS 0.008187f
C712 VDD1.n95 VSUBS 0.007953f
C713 VDD1.n96 VSUBS 0.0148f
C714 VDD1.n97 VSUBS 0.0148f
C715 VDD1.n98 VSUBS 0.007953f
C716 VDD1.n99 VSUBS 0.008421f
C717 VDD1.n100 VSUBS 0.018798f
C718 VDD1.n101 VSUBS 0.045511f
C719 VDD1.n102 VSUBS 0.008421f
C720 VDD1.n103 VSUBS 0.007953f
C721 VDD1.n104 VSUBS 0.036838f
C722 VDD1.n105 VSUBS 0.343719f
C723 VTAIL.n0 VSUBS 0.027177f
C724 VTAIL.n1 VSUBS 0.024732f
C725 VTAIL.n2 VSUBS 0.01329f
C726 VTAIL.n3 VSUBS 0.031413f
C727 VTAIL.n4 VSUBS 0.014072f
C728 VTAIL.n5 VSUBS 0.024732f
C729 VTAIL.n6 VSUBS 0.013681f
C730 VTAIL.n7 VSUBS 0.031413f
C731 VTAIL.n8 VSUBS 0.014072f
C732 VTAIL.n9 VSUBS 0.024732f
C733 VTAIL.n10 VSUBS 0.01329f
C734 VTAIL.n11 VSUBS 0.031413f
C735 VTAIL.n12 VSUBS 0.014072f
C736 VTAIL.n13 VSUBS 0.024732f
C737 VTAIL.n14 VSUBS 0.01329f
C738 VTAIL.n15 VSUBS 0.02356f
C739 VTAIL.n16 VSUBS 0.02363f
C740 VTAIL.t2 VSUBS 0.067555f
C741 VTAIL.n17 VSUBS 0.173442f
C742 VTAIL.n18 VSUBS 1.00815f
C743 VTAIL.n19 VSUBS 0.01329f
C744 VTAIL.n20 VSUBS 0.014072f
C745 VTAIL.n21 VSUBS 0.031413f
C746 VTAIL.n22 VSUBS 0.031413f
C747 VTAIL.n23 VSUBS 0.014072f
C748 VTAIL.n24 VSUBS 0.01329f
C749 VTAIL.n25 VSUBS 0.024732f
C750 VTAIL.n26 VSUBS 0.024732f
C751 VTAIL.n27 VSUBS 0.01329f
C752 VTAIL.n28 VSUBS 0.014072f
C753 VTAIL.n29 VSUBS 0.031413f
C754 VTAIL.n30 VSUBS 0.031413f
C755 VTAIL.n31 VSUBS 0.014072f
C756 VTAIL.n32 VSUBS 0.01329f
C757 VTAIL.n33 VSUBS 0.024732f
C758 VTAIL.n34 VSUBS 0.024732f
C759 VTAIL.n35 VSUBS 0.01329f
C760 VTAIL.n36 VSUBS 0.01329f
C761 VTAIL.n37 VSUBS 0.014072f
C762 VTAIL.n38 VSUBS 0.031413f
C763 VTAIL.n39 VSUBS 0.031413f
C764 VTAIL.n40 VSUBS 0.031413f
C765 VTAIL.n41 VSUBS 0.013681f
C766 VTAIL.n42 VSUBS 0.01329f
C767 VTAIL.n43 VSUBS 0.024732f
C768 VTAIL.n44 VSUBS 0.024732f
C769 VTAIL.n45 VSUBS 0.01329f
C770 VTAIL.n46 VSUBS 0.014072f
C771 VTAIL.n47 VSUBS 0.031413f
C772 VTAIL.n48 VSUBS 0.076052f
C773 VTAIL.n49 VSUBS 0.014072f
C774 VTAIL.n50 VSUBS 0.01329f
C775 VTAIL.n51 VSUBS 0.06156f
C776 VTAIL.n52 VSUBS 0.038377f
C777 VTAIL.n53 VSUBS 1.28015f
C778 VTAIL.n54 VSUBS 0.027177f
C779 VTAIL.n55 VSUBS 0.024732f
C780 VTAIL.n56 VSUBS 0.01329f
C781 VTAIL.n57 VSUBS 0.031413f
C782 VTAIL.n58 VSUBS 0.014072f
C783 VTAIL.n59 VSUBS 0.024732f
C784 VTAIL.n60 VSUBS 0.013681f
C785 VTAIL.n61 VSUBS 0.031413f
C786 VTAIL.n62 VSUBS 0.01329f
C787 VTAIL.n63 VSUBS 0.014072f
C788 VTAIL.n64 VSUBS 0.024732f
C789 VTAIL.n65 VSUBS 0.01329f
C790 VTAIL.n66 VSUBS 0.031413f
C791 VTAIL.n67 VSUBS 0.014072f
C792 VTAIL.n68 VSUBS 0.024732f
C793 VTAIL.n69 VSUBS 0.01329f
C794 VTAIL.n70 VSUBS 0.02356f
C795 VTAIL.n71 VSUBS 0.02363f
C796 VTAIL.t0 VSUBS 0.067555f
C797 VTAIL.n72 VSUBS 0.173442f
C798 VTAIL.n73 VSUBS 1.00815f
C799 VTAIL.n74 VSUBS 0.01329f
C800 VTAIL.n75 VSUBS 0.014072f
C801 VTAIL.n76 VSUBS 0.031413f
C802 VTAIL.n77 VSUBS 0.031413f
C803 VTAIL.n78 VSUBS 0.014072f
C804 VTAIL.n79 VSUBS 0.01329f
C805 VTAIL.n80 VSUBS 0.024732f
C806 VTAIL.n81 VSUBS 0.024732f
C807 VTAIL.n82 VSUBS 0.01329f
C808 VTAIL.n83 VSUBS 0.014072f
C809 VTAIL.n84 VSUBS 0.031413f
C810 VTAIL.n85 VSUBS 0.031413f
C811 VTAIL.n86 VSUBS 0.014072f
C812 VTAIL.n87 VSUBS 0.01329f
C813 VTAIL.n88 VSUBS 0.024732f
C814 VTAIL.n89 VSUBS 0.024732f
C815 VTAIL.n90 VSUBS 0.01329f
C816 VTAIL.n91 VSUBS 0.014072f
C817 VTAIL.n92 VSUBS 0.031413f
C818 VTAIL.n93 VSUBS 0.031413f
C819 VTAIL.n94 VSUBS 0.031413f
C820 VTAIL.n95 VSUBS 0.013681f
C821 VTAIL.n96 VSUBS 0.01329f
C822 VTAIL.n97 VSUBS 0.024732f
C823 VTAIL.n98 VSUBS 0.024732f
C824 VTAIL.n99 VSUBS 0.01329f
C825 VTAIL.n100 VSUBS 0.014072f
C826 VTAIL.n101 VSUBS 0.031413f
C827 VTAIL.n102 VSUBS 0.076052f
C828 VTAIL.n103 VSUBS 0.014072f
C829 VTAIL.n104 VSUBS 0.01329f
C830 VTAIL.n105 VSUBS 0.06156f
C831 VTAIL.n106 VSUBS 0.038377f
C832 VTAIL.n107 VSUBS 1.29595f
C833 VTAIL.n108 VSUBS 0.027177f
C834 VTAIL.n109 VSUBS 0.024732f
C835 VTAIL.n110 VSUBS 0.01329f
C836 VTAIL.n111 VSUBS 0.031413f
C837 VTAIL.n112 VSUBS 0.014072f
C838 VTAIL.n113 VSUBS 0.024732f
C839 VTAIL.n114 VSUBS 0.013681f
C840 VTAIL.n115 VSUBS 0.031413f
C841 VTAIL.n116 VSUBS 0.01329f
C842 VTAIL.n117 VSUBS 0.014072f
C843 VTAIL.n118 VSUBS 0.024732f
C844 VTAIL.n119 VSUBS 0.01329f
C845 VTAIL.n120 VSUBS 0.031413f
C846 VTAIL.n121 VSUBS 0.014072f
C847 VTAIL.n122 VSUBS 0.024732f
C848 VTAIL.n123 VSUBS 0.01329f
C849 VTAIL.n124 VSUBS 0.02356f
C850 VTAIL.n125 VSUBS 0.02363f
C851 VTAIL.t3 VSUBS 0.067555f
C852 VTAIL.n126 VSUBS 0.173442f
C853 VTAIL.n127 VSUBS 1.00815f
C854 VTAIL.n128 VSUBS 0.01329f
C855 VTAIL.n129 VSUBS 0.014072f
C856 VTAIL.n130 VSUBS 0.031413f
C857 VTAIL.n131 VSUBS 0.031413f
C858 VTAIL.n132 VSUBS 0.014072f
C859 VTAIL.n133 VSUBS 0.01329f
C860 VTAIL.n134 VSUBS 0.024732f
C861 VTAIL.n135 VSUBS 0.024732f
C862 VTAIL.n136 VSUBS 0.01329f
C863 VTAIL.n137 VSUBS 0.014072f
C864 VTAIL.n138 VSUBS 0.031413f
C865 VTAIL.n139 VSUBS 0.031413f
C866 VTAIL.n140 VSUBS 0.014072f
C867 VTAIL.n141 VSUBS 0.01329f
C868 VTAIL.n142 VSUBS 0.024732f
C869 VTAIL.n143 VSUBS 0.024732f
C870 VTAIL.n144 VSUBS 0.01329f
C871 VTAIL.n145 VSUBS 0.014072f
C872 VTAIL.n146 VSUBS 0.031413f
C873 VTAIL.n147 VSUBS 0.031413f
C874 VTAIL.n148 VSUBS 0.031413f
C875 VTAIL.n149 VSUBS 0.013681f
C876 VTAIL.n150 VSUBS 0.01329f
C877 VTAIL.n151 VSUBS 0.024732f
C878 VTAIL.n152 VSUBS 0.024732f
C879 VTAIL.n153 VSUBS 0.01329f
C880 VTAIL.n154 VSUBS 0.014072f
C881 VTAIL.n155 VSUBS 0.031413f
C882 VTAIL.n156 VSUBS 0.076052f
C883 VTAIL.n157 VSUBS 0.014072f
C884 VTAIL.n158 VSUBS 0.01329f
C885 VTAIL.n159 VSUBS 0.06156f
C886 VTAIL.n160 VSUBS 0.038377f
C887 VTAIL.n161 VSUBS 1.2142f
C888 VTAIL.n162 VSUBS 0.027177f
C889 VTAIL.n163 VSUBS 0.024732f
C890 VTAIL.n164 VSUBS 0.01329f
C891 VTAIL.n165 VSUBS 0.031413f
C892 VTAIL.n166 VSUBS 0.014072f
C893 VTAIL.n167 VSUBS 0.024732f
C894 VTAIL.n168 VSUBS 0.013681f
C895 VTAIL.n169 VSUBS 0.031413f
C896 VTAIL.n170 VSUBS 0.014072f
C897 VTAIL.n171 VSUBS 0.024732f
C898 VTAIL.n172 VSUBS 0.01329f
C899 VTAIL.n173 VSUBS 0.031413f
C900 VTAIL.n174 VSUBS 0.014072f
C901 VTAIL.n175 VSUBS 0.024732f
C902 VTAIL.n176 VSUBS 0.01329f
C903 VTAIL.n177 VSUBS 0.02356f
C904 VTAIL.n178 VSUBS 0.02363f
C905 VTAIL.t1 VSUBS 0.067555f
C906 VTAIL.n179 VSUBS 0.173442f
C907 VTAIL.n180 VSUBS 1.00815f
C908 VTAIL.n181 VSUBS 0.01329f
C909 VTAIL.n182 VSUBS 0.014072f
C910 VTAIL.n183 VSUBS 0.031413f
C911 VTAIL.n184 VSUBS 0.031413f
C912 VTAIL.n185 VSUBS 0.014072f
C913 VTAIL.n186 VSUBS 0.01329f
C914 VTAIL.n187 VSUBS 0.024732f
C915 VTAIL.n188 VSUBS 0.024732f
C916 VTAIL.n189 VSUBS 0.01329f
C917 VTAIL.n190 VSUBS 0.014072f
C918 VTAIL.n191 VSUBS 0.031413f
C919 VTAIL.n192 VSUBS 0.031413f
C920 VTAIL.n193 VSUBS 0.014072f
C921 VTAIL.n194 VSUBS 0.01329f
C922 VTAIL.n195 VSUBS 0.024732f
C923 VTAIL.n196 VSUBS 0.024732f
C924 VTAIL.n197 VSUBS 0.01329f
C925 VTAIL.n198 VSUBS 0.01329f
C926 VTAIL.n199 VSUBS 0.014072f
C927 VTAIL.n200 VSUBS 0.031413f
C928 VTAIL.n201 VSUBS 0.031413f
C929 VTAIL.n202 VSUBS 0.031413f
C930 VTAIL.n203 VSUBS 0.013681f
C931 VTAIL.n204 VSUBS 0.01329f
C932 VTAIL.n205 VSUBS 0.024732f
C933 VTAIL.n206 VSUBS 0.024732f
C934 VTAIL.n207 VSUBS 0.01329f
C935 VTAIL.n208 VSUBS 0.014072f
C936 VTAIL.n209 VSUBS 0.031413f
C937 VTAIL.n210 VSUBS 0.076052f
C938 VTAIL.n211 VSUBS 0.014072f
C939 VTAIL.n212 VSUBS 0.01329f
C940 VTAIL.n213 VSUBS 0.06156f
C941 VTAIL.n214 VSUBS 0.038377f
C942 VTAIL.n215 VSUBS 1.15168f
C943 VP.t0 VSUBS 0.942797f
C944 VP.t1 VSUBS 0.848797f
C945 VP.n0 VSUBS 2.49491f
.ends

