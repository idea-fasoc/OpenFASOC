* NGSPICE file created from diff_pair_sample_0426.ext - technology: sky130A

.subckt diff_pair_sample_0426 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=3.8298 ps=20.42 w=9.82 l=3.16
X1 VDD1.t9 VP.t0 VTAIL.t15 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=1.6203 ps=10.15 w=9.82 l=3.16
X2 VTAIL.t11 VN.t1 VDD2.t8 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X3 VTAIL.t7 VN.t2 VDD2.t7 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X4 VDD2.t6 VN.t3 VTAIL.t8 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=1.6203 ps=10.15 w=9.82 l=3.16
X5 VDD2.t5 VN.t4 VTAIL.t3 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X6 B.t11 B.t9 B.t10 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=0 ps=0 w=9.82 l=3.16
X7 B.t8 B.t6 B.t7 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=0 ps=0 w=9.82 l=3.16
X8 VDD2.t4 VN.t5 VTAIL.t4 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=3.8298 ps=20.42 w=9.82 l=3.16
X9 VTAIL.t14 VP.t1 VDD1.t8 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X10 VDD2.t3 VN.t6 VTAIL.t2 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=1.6203 ps=10.15 w=9.82 l=3.16
X11 VTAIL.t18 VP.t2 VDD1.t7 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X12 VDD1.t6 VP.t3 VTAIL.t0 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=1.6203 ps=10.15 w=9.82 l=3.16
X13 B.t5 B.t3 B.t4 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=0 ps=0 w=9.82 l=3.16
X14 VTAIL.t1 VP.t4 VDD1.t5 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X15 VDD2.t2 VN.t7 VTAIL.t9 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X16 VDD1.t4 VP.t5 VTAIL.t17 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=3.8298 ps=20.42 w=9.82 l=3.16
X17 VTAIL.t12 VP.t6 VDD1.t3 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X18 VDD1.t2 VP.t7 VTAIL.t13 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X19 VDD1.t1 VP.t8 VTAIL.t16 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=3.8298 ps=20.42 w=9.82 l=3.16
X20 B.t2 B.t0 B.t1 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=3.8298 pd=20.42 as=0 ps=0 w=9.82 l=3.16
X21 VDD1.t0 VP.t9 VTAIL.t19 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X22 VTAIL.t6 VN.t8 VDD2.t1 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
X23 VTAIL.t5 VN.t9 VDD2.t0 w_n5158_n2932# sky130_fd_pr__pfet_01v8 ad=1.6203 pd=10.15 as=1.6203 ps=10.15 w=9.82 l=3.16
R0 VN.n94 VN.n93 161.3
R1 VN.n92 VN.n49 161.3
R2 VN.n91 VN.n90 161.3
R3 VN.n89 VN.n50 161.3
R4 VN.n88 VN.n87 161.3
R5 VN.n86 VN.n51 161.3
R6 VN.n85 VN.n84 161.3
R7 VN.n83 VN.n82 161.3
R8 VN.n81 VN.n53 161.3
R9 VN.n80 VN.n79 161.3
R10 VN.n78 VN.n54 161.3
R11 VN.n77 VN.n76 161.3
R12 VN.n75 VN.n55 161.3
R13 VN.n74 VN.n73 161.3
R14 VN.n72 VN.n71 161.3
R15 VN.n70 VN.n57 161.3
R16 VN.n69 VN.n68 161.3
R17 VN.n67 VN.n58 161.3
R18 VN.n66 VN.n65 161.3
R19 VN.n64 VN.n59 161.3
R20 VN.n63 VN.n62 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n1 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n41 VN.n2 161.3
R25 VN.n40 VN.n39 161.3
R26 VN.n38 VN.n3 161.3
R27 VN.n37 VN.n36 161.3
R28 VN.n35 VN.n34 161.3
R29 VN.n33 VN.n5 161.3
R30 VN.n32 VN.n31 161.3
R31 VN.n30 VN.n6 161.3
R32 VN.n29 VN.n28 161.3
R33 VN.n27 VN.n7 161.3
R34 VN.n26 VN.n25 161.3
R35 VN.n24 VN.n23 161.3
R36 VN.n22 VN.n9 161.3
R37 VN.n21 VN.n20 161.3
R38 VN.n19 VN.n10 161.3
R39 VN.n18 VN.n17 161.3
R40 VN.n16 VN.n11 161.3
R41 VN.n15 VN.n14 161.3
R42 VN.n61 VN.t5 107.288
R43 VN.n13 VN.t3 107.288
R44 VN.n47 VN.n0 78.693
R45 VN.n95 VN.n48 78.693
R46 VN.n12 VN.t1 74.8935
R47 VN.n8 VN.t4 74.8935
R48 VN.n4 VN.t2 74.8935
R49 VN.n0 VN.t0 74.8935
R50 VN.n60 VN.t9 74.8935
R51 VN.n56 VN.t7 74.8935
R52 VN.n52 VN.t8 74.8935
R53 VN.n48 VN.t6 74.8935
R54 VN.n13 VN.n12 62.3674
R55 VN.n61 VN.n60 62.3674
R56 VN VN.n95 54.6987
R57 VN.n39 VN.n2 41.8712
R58 VN.n87 VN.n50 41.8712
R59 VN.n21 VN.n10 40.8975
R60 VN.n28 VN.n6 40.8975
R61 VN.n69 VN.n58 40.8975
R62 VN.n76 VN.n54 40.8975
R63 VN.n17 VN.n10 39.9237
R64 VN.n32 VN.n6 39.9237
R65 VN.n65 VN.n58 39.9237
R66 VN.n80 VN.n54 39.9237
R67 VN.n43 VN.n2 38.95
R68 VN.n91 VN.n50 38.95
R69 VN.n16 VN.n15 24.3439
R70 VN.n17 VN.n16 24.3439
R71 VN.n22 VN.n21 24.3439
R72 VN.n23 VN.n22 24.3439
R73 VN.n27 VN.n26 24.3439
R74 VN.n28 VN.n27 24.3439
R75 VN.n33 VN.n32 24.3439
R76 VN.n34 VN.n33 24.3439
R77 VN.n38 VN.n37 24.3439
R78 VN.n39 VN.n38 24.3439
R79 VN.n44 VN.n43 24.3439
R80 VN.n45 VN.n44 24.3439
R81 VN.n65 VN.n64 24.3439
R82 VN.n64 VN.n63 24.3439
R83 VN.n76 VN.n75 24.3439
R84 VN.n75 VN.n74 24.3439
R85 VN.n71 VN.n70 24.3439
R86 VN.n70 VN.n69 24.3439
R87 VN.n87 VN.n86 24.3439
R88 VN.n86 VN.n85 24.3439
R89 VN.n82 VN.n81 24.3439
R90 VN.n81 VN.n80 24.3439
R91 VN.n93 VN.n92 24.3439
R92 VN.n92 VN.n91 24.3439
R93 VN.n37 VN.n4 12.6591
R94 VN.n85 VN.n52 12.6591
R95 VN.n23 VN.n8 12.1722
R96 VN.n26 VN.n8 12.1722
R97 VN.n74 VN.n56 12.1722
R98 VN.n71 VN.n56 12.1722
R99 VN.n15 VN.n12 11.6853
R100 VN.n34 VN.n4 11.6853
R101 VN.n63 VN.n60 11.6853
R102 VN.n82 VN.n52 11.6853
R103 VN.n45 VN.n0 11.1985
R104 VN.n93 VN.n48 11.1985
R105 VN.n62 VN.n61 4.34077
R106 VN.n14 VN.n13 4.34077
R107 VN.n95 VN.n94 0.355081
R108 VN.n47 VN.n46 0.355081
R109 VN VN.n47 0.26685
R110 VN.n94 VN.n49 0.189894
R111 VN.n90 VN.n49 0.189894
R112 VN.n90 VN.n89 0.189894
R113 VN.n89 VN.n88 0.189894
R114 VN.n88 VN.n51 0.189894
R115 VN.n84 VN.n51 0.189894
R116 VN.n84 VN.n83 0.189894
R117 VN.n83 VN.n53 0.189894
R118 VN.n79 VN.n53 0.189894
R119 VN.n79 VN.n78 0.189894
R120 VN.n78 VN.n77 0.189894
R121 VN.n77 VN.n55 0.189894
R122 VN.n73 VN.n55 0.189894
R123 VN.n73 VN.n72 0.189894
R124 VN.n72 VN.n57 0.189894
R125 VN.n68 VN.n57 0.189894
R126 VN.n68 VN.n67 0.189894
R127 VN.n67 VN.n66 0.189894
R128 VN.n66 VN.n59 0.189894
R129 VN.n62 VN.n59 0.189894
R130 VN.n14 VN.n11 0.189894
R131 VN.n18 VN.n11 0.189894
R132 VN.n19 VN.n18 0.189894
R133 VN.n20 VN.n19 0.189894
R134 VN.n20 VN.n9 0.189894
R135 VN.n24 VN.n9 0.189894
R136 VN.n25 VN.n24 0.189894
R137 VN.n25 VN.n7 0.189894
R138 VN.n29 VN.n7 0.189894
R139 VN.n30 VN.n29 0.189894
R140 VN.n31 VN.n30 0.189894
R141 VN.n31 VN.n5 0.189894
R142 VN.n35 VN.n5 0.189894
R143 VN.n36 VN.n35 0.189894
R144 VN.n36 VN.n3 0.189894
R145 VN.n40 VN.n3 0.189894
R146 VN.n41 VN.n40 0.189894
R147 VN.n42 VN.n41 0.189894
R148 VN.n42 VN.n1 0.189894
R149 VN.n46 VN.n1 0.189894
R150 VTAIL.n11 VTAIL.t4 68.7183
R151 VTAIL.n17 VTAIL.t10 68.7182
R152 VTAIL.n2 VTAIL.t16 68.7182
R153 VTAIL.n16 VTAIL.t17 68.7182
R154 VTAIL.n15 VTAIL.n14 65.4083
R155 VTAIL.n13 VTAIL.n12 65.4083
R156 VTAIL.n10 VTAIL.n9 65.4083
R157 VTAIL.n8 VTAIL.n7 65.4083
R158 VTAIL.n19 VTAIL.n18 65.408
R159 VTAIL.n1 VTAIL.n0 65.408
R160 VTAIL.n4 VTAIL.n3 65.408
R161 VTAIL.n6 VTAIL.n5 65.408
R162 VTAIL.n8 VTAIL.n6 26.8496
R163 VTAIL.n17 VTAIL.n16 23.841
R164 VTAIL.n18 VTAIL.t3 3.31058
R165 VTAIL.n18 VTAIL.t7 3.31058
R166 VTAIL.n0 VTAIL.t8 3.31058
R167 VTAIL.n0 VTAIL.t11 3.31058
R168 VTAIL.n3 VTAIL.t13 3.31058
R169 VTAIL.n3 VTAIL.t12 3.31058
R170 VTAIL.n5 VTAIL.t0 3.31058
R171 VTAIL.n5 VTAIL.t1 3.31058
R172 VTAIL.n14 VTAIL.t19 3.31058
R173 VTAIL.n14 VTAIL.t14 3.31058
R174 VTAIL.n12 VTAIL.t15 3.31058
R175 VTAIL.n12 VTAIL.t18 3.31058
R176 VTAIL.n9 VTAIL.t9 3.31058
R177 VTAIL.n9 VTAIL.t5 3.31058
R178 VTAIL.n7 VTAIL.t2 3.31058
R179 VTAIL.n7 VTAIL.t6 3.31058
R180 VTAIL.n10 VTAIL.n8 3.00912
R181 VTAIL.n11 VTAIL.n10 3.00912
R182 VTAIL.n15 VTAIL.n13 3.00912
R183 VTAIL.n16 VTAIL.n15 3.00912
R184 VTAIL.n6 VTAIL.n4 3.00912
R185 VTAIL.n4 VTAIL.n2 3.00912
R186 VTAIL.n19 VTAIL.n17 3.00912
R187 VTAIL VTAIL.n1 2.31516
R188 VTAIL.n13 VTAIL.n11 1.97464
R189 VTAIL.n2 VTAIL.n1 1.97464
R190 VTAIL VTAIL.n19 0.694465
R191 VDD2.n1 VDD2.t6 88.4056
R192 VDD2.n4 VDD2.t3 85.3971
R193 VDD2.n3 VDD2.n2 84.2879
R194 VDD2 VDD2.n7 84.2851
R195 VDD2.n6 VDD2.n5 82.0871
R196 VDD2.n1 VDD2.n0 82.0868
R197 VDD2.n4 VDD2.n3 46.4718
R198 VDD2.n7 VDD2.t0 3.31058
R199 VDD2.n7 VDD2.t4 3.31058
R200 VDD2.n5 VDD2.t1 3.31058
R201 VDD2.n5 VDD2.t2 3.31058
R202 VDD2.n2 VDD2.t7 3.31058
R203 VDD2.n2 VDD2.t9 3.31058
R204 VDD2.n0 VDD2.t8 3.31058
R205 VDD2.n0 VDD2.t5 3.31058
R206 VDD2.n6 VDD2.n4 3.00912
R207 VDD2 VDD2.n6 0.810845
R208 VDD2.n3 VDD2.n1 0.697309
R209 VP.n32 VP.n31 161.3
R210 VP.n33 VP.n28 161.3
R211 VP.n35 VP.n34 161.3
R212 VP.n36 VP.n27 161.3
R213 VP.n38 VP.n37 161.3
R214 VP.n39 VP.n26 161.3
R215 VP.n41 VP.n40 161.3
R216 VP.n43 VP.n42 161.3
R217 VP.n44 VP.n24 161.3
R218 VP.n46 VP.n45 161.3
R219 VP.n47 VP.n23 161.3
R220 VP.n49 VP.n48 161.3
R221 VP.n50 VP.n22 161.3
R222 VP.n52 VP.n51 161.3
R223 VP.n54 VP.n53 161.3
R224 VP.n55 VP.n20 161.3
R225 VP.n57 VP.n56 161.3
R226 VP.n58 VP.n19 161.3
R227 VP.n60 VP.n59 161.3
R228 VP.n61 VP.n18 161.3
R229 VP.n63 VP.n62 161.3
R230 VP.n109 VP.n108 161.3
R231 VP.n107 VP.n1 161.3
R232 VP.n106 VP.n105 161.3
R233 VP.n104 VP.n2 161.3
R234 VP.n103 VP.n102 161.3
R235 VP.n101 VP.n3 161.3
R236 VP.n100 VP.n99 161.3
R237 VP.n98 VP.n97 161.3
R238 VP.n96 VP.n5 161.3
R239 VP.n95 VP.n94 161.3
R240 VP.n93 VP.n6 161.3
R241 VP.n92 VP.n91 161.3
R242 VP.n90 VP.n7 161.3
R243 VP.n89 VP.n88 161.3
R244 VP.n87 VP.n86 161.3
R245 VP.n85 VP.n9 161.3
R246 VP.n84 VP.n83 161.3
R247 VP.n82 VP.n10 161.3
R248 VP.n81 VP.n80 161.3
R249 VP.n79 VP.n11 161.3
R250 VP.n78 VP.n77 161.3
R251 VP.n76 VP.n75 161.3
R252 VP.n74 VP.n13 161.3
R253 VP.n73 VP.n72 161.3
R254 VP.n71 VP.n14 161.3
R255 VP.n70 VP.n69 161.3
R256 VP.n68 VP.n15 161.3
R257 VP.n67 VP.n66 161.3
R258 VP.n30 VP.t0 107.288
R259 VP.n65 VP.n16 78.693
R260 VP.n110 VP.n0 78.693
R261 VP.n64 VP.n17 78.693
R262 VP.n16 VP.t3 74.8935
R263 VP.n12 VP.t4 74.8935
R264 VP.n8 VP.t7 74.8935
R265 VP.n4 VP.t6 74.8935
R266 VP.n0 VP.t8 74.8935
R267 VP.n17 VP.t5 74.8935
R268 VP.n21 VP.t1 74.8935
R269 VP.n25 VP.t9 74.8935
R270 VP.n29 VP.t2 74.8935
R271 VP.n30 VP.n29 62.3674
R272 VP.n65 VP.n64 54.5332
R273 VP.n73 VP.n14 41.8712
R274 VP.n102 VP.n2 41.8712
R275 VP.n56 VP.n19 41.8712
R276 VP.n84 VP.n10 40.8975
R277 VP.n91 VP.n6 40.8975
R278 VP.n45 VP.n23 40.8975
R279 VP.n38 VP.n27 40.8975
R280 VP.n80 VP.n10 39.9237
R281 VP.n95 VP.n6 39.9237
R282 VP.n49 VP.n23 39.9237
R283 VP.n34 VP.n27 39.9237
R284 VP.n69 VP.n14 38.95
R285 VP.n106 VP.n2 38.95
R286 VP.n60 VP.n19 38.95
R287 VP.n68 VP.n67 24.3439
R288 VP.n69 VP.n68 24.3439
R289 VP.n74 VP.n73 24.3439
R290 VP.n75 VP.n74 24.3439
R291 VP.n79 VP.n78 24.3439
R292 VP.n80 VP.n79 24.3439
R293 VP.n85 VP.n84 24.3439
R294 VP.n86 VP.n85 24.3439
R295 VP.n90 VP.n89 24.3439
R296 VP.n91 VP.n90 24.3439
R297 VP.n96 VP.n95 24.3439
R298 VP.n97 VP.n96 24.3439
R299 VP.n101 VP.n100 24.3439
R300 VP.n102 VP.n101 24.3439
R301 VP.n107 VP.n106 24.3439
R302 VP.n108 VP.n107 24.3439
R303 VP.n61 VP.n60 24.3439
R304 VP.n62 VP.n61 24.3439
R305 VP.n50 VP.n49 24.3439
R306 VP.n51 VP.n50 24.3439
R307 VP.n55 VP.n54 24.3439
R308 VP.n56 VP.n55 24.3439
R309 VP.n39 VP.n38 24.3439
R310 VP.n40 VP.n39 24.3439
R311 VP.n44 VP.n43 24.3439
R312 VP.n45 VP.n44 24.3439
R313 VP.n33 VP.n32 24.3439
R314 VP.n34 VP.n33 24.3439
R315 VP.n75 VP.n12 12.6591
R316 VP.n100 VP.n4 12.6591
R317 VP.n54 VP.n21 12.6591
R318 VP.n86 VP.n8 12.1722
R319 VP.n89 VP.n8 12.1722
R320 VP.n40 VP.n25 12.1722
R321 VP.n43 VP.n25 12.1722
R322 VP.n78 VP.n12 11.6853
R323 VP.n97 VP.n4 11.6853
R324 VP.n51 VP.n21 11.6853
R325 VP.n32 VP.n29 11.6853
R326 VP.n67 VP.n16 11.1985
R327 VP.n108 VP.n0 11.1985
R328 VP.n62 VP.n17 11.1985
R329 VP.n31 VP.n30 4.34075
R330 VP.n64 VP.n63 0.355081
R331 VP.n66 VP.n65 0.355081
R332 VP.n110 VP.n109 0.355081
R333 VP VP.n110 0.26685
R334 VP.n31 VP.n28 0.189894
R335 VP.n35 VP.n28 0.189894
R336 VP.n36 VP.n35 0.189894
R337 VP.n37 VP.n36 0.189894
R338 VP.n37 VP.n26 0.189894
R339 VP.n41 VP.n26 0.189894
R340 VP.n42 VP.n41 0.189894
R341 VP.n42 VP.n24 0.189894
R342 VP.n46 VP.n24 0.189894
R343 VP.n47 VP.n46 0.189894
R344 VP.n48 VP.n47 0.189894
R345 VP.n48 VP.n22 0.189894
R346 VP.n52 VP.n22 0.189894
R347 VP.n53 VP.n52 0.189894
R348 VP.n53 VP.n20 0.189894
R349 VP.n57 VP.n20 0.189894
R350 VP.n58 VP.n57 0.189894
R351 VP.n59 VP.n58 0.189894
R352 VP.n59 VP.n18 0.189894
R353 VP.n63 VP.n18 0.189894
R354 VP.n66 VP.n15 0.189894
R355 VP.n70 VP.n15 0.189894
R356 VP.n71 VP.n70 0.189894
R357 VP.n72 VP.n71 0.189894
R358 VP.n72 VP.n13 0.189894
R359 VP.n76 VP.n13 0.189894
R360 VP.n77 VP.n76 0.189894
R361 VP.n77 VP.n11 0.189894
R362 VP.n81 VP.n11 0.189894
R363 VP.n82 VP.n81 0.189894
R364 VP.n83 VP.n82 0.189894
R365 VP.n83 VP.n9 0.189894
R366 VP.n87 VP.n9 0.189894
R367 VP.n88 VP.n87 0.189894
R368 VP.n88 VP.n7 0.189894
R369 VP.n92 VP.n7 0.189894
R370 VP.n93 VP.n92 0.189894
R371 VP.n94 VP.n93 0.189894
R372 VP.n94 VP.n5 0.189894
R373 VP.n98 VP.n5 0.189894
R374 VP.n99 VP.n98 0.189894
R375 VP.n99 VP.n3 0.189894
R376 VP.n103 VP.n3 0.189894
R377 VP.n104 VP.n103 0.189894
R378 VP.n105 VP.n104 0.189894
R379 VP.n105 VP.n1 0.189894
R380 VP.n109 VP.n1 0.189894
R381 VDD1.n1 VDD1.t9 88.4057
R382 VDD1.n3 VDD1.t6 88.4056
R383 VDD1.n5 VDD1.n4 84.2879
R384 VDD1.n1 VDD1.n0 82.0871
R385 VDD1.n7 VDD1.n6 82.0869
R386 VDD1.n3 VDD1.n2 82.0868
R387 VDD1.n7 VDD1.n5 48.5591
R388 VDD1.n6 VDD1.t8 3.31058
R389 VDD1.n6 VDD1.t4 3.31058
R390 VDD1.n0 VDD1.t7 3.31058
R391 VDD1.n0 VDD1.t0 3.31058
R392 VDD1.n4 VDD1.t3 3.31058
R393 VDD1.n4 VDD1.t1 3.31058
R394 VDD1.n2 VDD1.t5 3.31058
R395 VDD1.n2 VDD1.t2 3.31058
R396 VDD1 VDD1.n7 2.19878
R397 VDD1 VDD1.n1 0.810845
R398 VDD1.n5 VDD1.n3 0.697309
R399 B.n452 B.n151 585
R400 B.n451 B.n450 585
R401 B.n449 B.n152 585
R402 B.n448 B.n447 585
R403 B.n446 B.n153 585
R404 B.n445 B.n444 585
R405 B.n443 B.n154 585
R406 B.n442 B.n441 585
R407 B.n440 B.n155 585
R408 B.n439 B.n438 585
R409 B.n437 B.n156 585
R410 B.n436 B.n435 585
R411 B.n434 B.n157 585
R412 B.n433 B.n432 585
R413 B.n431 B.n158 585
R414 B.n430 B.n429 585
R415 B.n428 B.n159 585
R416 B.n427 B.n426 585
R417 B.n425 B.n160 585
R418 B.n424 B.n423 585
R419 B.n422 B.n161 585
R420 B.n421 B.n420 585
R421 B.n419 B.n162 585
R422 B.n418 B.n417 585
R423 B.n416 B.n163 585
R424 B.n415 B.n414 585
R425 B.n413 B.n164 585
R426 B.n412 B.n411 585
R427 B.n410 B.n165 585
R428 B.n409 B.n408 585
R429 B.n407 B.n166 585
R430 B.n406 B.n405 585
R431 B.n404 B.n167 585
R432 B.n403 B.n402 585
R433 B.n401 B.n168 585
R434 B.n400 B.n399 585
R435 B.n395 B.n169 585
R436 B.n394 B.n393 585
R437 B.n392 B.n170 585
R438 B.n391 B.n390 585
R439 B.n389 B.n171 585
R440 B.n388 B.n387 585
R441 B.n386 B.n172 585
R442 B.n385 B.n384 585
R443 B.n383 B.n173 585
R444 B.n381 B.n380 585
R445 B.n379 B.n176 585
R446 B.n378 B.n377 585
R447 B.n376 B.n177 585
R448 B.n375 B.n374 585
R449 B.n373 B.n178 585
R450 B.n372 B.n371 585
R451 B.n370 B.n179 585
R452 B.n369 B.n368 585
R453 B.n367 B.n180 585
R454 B.n366 B.n365 585
R455 B.n364 B.n181 585
R456 B.n363 B.n362 585
R457 B.n361 B.n182 585
R458 B.n360 B.n359 585
R459 B.n358 B.n183 585
R460 B.n357 B.n356 585
R461 B.n355 B.n184 585
R462 B.n354 B.n353 585
R463 B.n352 B.n185 585
R464 B.n351 B.n350 585
R465 B.n349 B.n186 585
R466 B.n348 B.n347 585
R467 B.n346 B.n187 585
R468 B.n345 B.n344 585
R469 B.n343 B.n188 585
R470 B.n342 B.n341 585
R471 B.n340 B.n189 585
R472 B.n339 B.n338 585
R473 B.n337 B.n190 585
R474 B.n336 B.n335 585
R475 B.n334 B.n191 585
R476 B.n333 B.n332 585
R477 B.n331 B.n192 585
R478 B.n330 B.n329 585
R479 B.n454 B.n453 585
R480 B.n455 B.n150 585
R481 B.n457 B.n456 585
R482 B.n458 B.n149 585
R483 B.n460 B.n459 585
R484 B.n461 B.n148 585
R485 B.n463 B.n462 585
R486 B.n464 B.n147 585
R487 B.n466 B.n465 585
R488 B.n467 B.n146 585
R489 B.n469 B.n468 585
R490 B.n470 B.n145 585
R491 B.n472 B.n471 585
R492 B.n473 B.n144 585
R493 B.n475 B.n474 585
R494 B.n476 B.n143 585
R495 B.n478 B.n477 585
R496 B.n479 B.n142 585
R497 B.n481 B.n480 585
R498 B.n482 B.n141 585
R499 B.n484 B.n483 585
R500 B.n485 B.n140 585
R501 B.n487 B.n486 585
R502 B.n488 B.n139 585
R503 B.n490 B.n489 585
R504 B.n491 B.n138 585
R505 B.n493 B.n492 585
R506 B.n494 B.n137 585
R507 B.n496 B.n495 585
R508 B.n497 B.n136 585
R509 B.n499 B.n498 585
R510 B.n500 B.n135 585
R511 B.n502 B.n501 585
R512 B.n503 B.n134 585
R513 B.n505 B.n504 585
R514 B.n506 B.n133 585
R515 B.n508 B.n507 585
R516 B.n509 B.n132 585
R517 B.n511 B.n510 585
R518 B.n512 B.n131 585
R519 B.n514 B.n513 585
R520 B.n515 B.n130 585
R521 B.n517 B.n516 585
R522 B.n518 B.n129 585
R523 B.n520 B.n519 585
R524 B.n521 B.n128 585
R525 B.n523 B.n522 585
R526 B.n524 B.n127 585
R527 B.n526 B.n525 585
R528 B.n527 B.n126 585
R529 B.n529 B.n528 585
R530 B.n530 B.n125 585
R531 B.n532 B.n531 585
R532 B.n533 B.n124 585
R533 B.n535 B.n534 585
R534 B.n536 B.n123 585
R535 B.n538 B.n537 585
R536 B.n539 B.n122 585
R537 B.n541 B.n540 585
R538 B.n542 B.n121 585
R539 B.n544 B.n543 585
R540 B.n545 B.n120 585
R541 B.n547 B.n546 585
R542 B.n548 B.n119 585
R543 B.n550 B.n549 585
R544 B.n551 B.n118 585
R545 B.n553 B.n552 585
R546 B.n554 B.n117 585
R547 B.n556 B.n555 585
R548 B.n557 B.n116 585
R549 B.n559 B.n558 585
R550 B.n560 B.n115 585
R551 B.n562 B.n561 585
R552 B.n563 B.n114 585
R553 B.n565 B.n564 585
R554 B.n566 B.n113 585
R555 B.n568 B.n567 585
R556 B.n569 B.n112 585
R557 B.n571 B.n570 585
R558 B.n572 B.n111 585
R559 B.n574 B.n573 585
R560 B.n575 B.n110 585
R561 B.n577 B.n576 585
R562 B.n578 B.n109 585
R563 B.n580 B.n579 585
R564 B.n581 B.n108 585
R565 B.n583 B.n582 585
R566 B.n584 B.n107 585
R567 B.n586 B.n585 585
R568 B.n587 B.n106 585
R569 B.n589 B.n588 585
R570 B.n590 B.n105 585
R571 B.n592 B.n591 585
R572 B.n593 B.n104 585
R573 B.n595 B.n594 585
R574 B.n596 B.n103 585
R575 B.n598 B.n597 585
R576 B.n599 B.n102 585
R577 B.n601 B.n600 585
R578 B.n602 B.n101 585
R579 B.n604 B.n603 585
R580 B.n605 B.n100 585
R581 B.n607 B.n606 585
R582 B.n608 B.n99 585
R583 B.n610 B.n609 585
R584 B.n611 B.n98 585
R585 B.n613 B.n612 585
R586 B.n614 B.n97 585
R587 B.n616 B.n615 585
R588 B.n617 B.n96 585
R589 B.n619 B.n618 585
R590 B.n620 B.n95 585
R591 B.n622 B.n621 585
R592 B.n623 B.n94 585
R593 B.n625 B.n624 585
R594 B.n626 B.n93 585
R595 B.n628 B.n627 585
R596 B.n629 B.n92 585
R597 B.n631 B.n630 585
R598 B.n632 B.n91 585
R599 B.n634 B.n633 585
R600 B.n635 B.n90 585
R601 B.n637 B.n636 585
R602 B.n638 B.n89 585
R603 B.n640 B.n639 585
R604 B.n641 B.n88 585
R605 B.n643 B.n642 585
R606 B.n644 B.n87 585
R607 B.n646 B.n645 585
R608 B.n647 B.n86 585
R609 B.n649 B.n648 585
R610 B.n650 B.n85 585
R611 B.n652 B.n651 585
R612 B.n653 B.n84 585
R613 B.n655 B.n654 585
R614 B.n656 B.n83 585
R615 B.n658 B.n657 585
R616 B.n659 B.n82 585
R617 B.n661 B.n660 585
R618 B.n662 B.n81 585
R619 B.n784 B.n783 585
R620 B.n782 B.n37 585
R621 B.n781 B.n780 585
R622 B.n779 B.n38 585
R623 B.n778 B.n777 585
R624 B.n776 B.n39 585
R625 B.n775 B.n774 585
R626 B.n773 B.n40 585
R627 B.n772 B.n771 585
R628 B.n770 B.n41 585
R629 B.n769 B.n768 585
R630 B.n767 B.n42 585
R631 B.n766 B.n765 585
R632 B.n764 B.n43 585
R633 B.n763 B.n762 585
R634 B.n761 B.n44 585
R635 B.n760 B.n759 585
R636 B.n758 B.n45 585
R637 B.n757 B.n756 585
R638 B.n755 B.n46 585
R639 B.n754 B.n753 585
R640 B.n752 B.n47 585
R641 B.n751 B.n750 585
R642 B.n749 B.n48 585
R643 B.n748 B.n747 585
R644 B.n746 B.n49 585
R645 B.n745 B.n744 585
R646 B.n743 B.n50 585
R647 B.n742 B.n741 585
R648 B.n740 B.n51 585
R649 B.n739 B.n738 585
R650 B.n737 B.n52 585
R651 B.n736 B.n735 585
R652 B.n734 B.n53 585
R653 B.n733 B.n732 585
R654 B.n731 B.n730 585
R655 B.n729 B.n57 585
R656 B.n728 B.n727 585
R657 B.n726 B.n58 585
R658 B.n725 B.n724 585
R659 B.n723 B.n59 585
R660 B.n722 B.n721 585
R661 B.n720 B.n60 585
R662 B.n719 B.n718 585
R663 B.n717 B.n61 585
R664 B.n715 B.n714 585
R665 B.n713 B.n64 585
R666 B.n712 B.n711 585
R667 B.n710 B.n65 585
R668 B.n709 B.n708 585
R669 B.n707 B.n66 585
R670 B.n706 B.n705 585
R671 B.n704 B.n67 585
R672 B.n703 B.n702 585
R673 B.n701 B.n68 585
R674 B.n700 B.n699 585
R675 B.n698 B.n69 585
R676 B.n697 B.n696 585
R677 B.n695 B.n70 585
R678 B.n694 B.n693 585
R679 B.n692 B.n71 585
R680 B.n691 B.n690 585
R681 B.n689 B.n72 585
R682 B.n688 B.n687 585
R683 B.n686 B.n73 585
R684 B.n685 B.n684 585
R685 B.n683 B.n74 585
R686 B.n682 B.n681 585
R687 B.n680 B.n75 585
R688 B.n679 B.n678 585
R689 B.n677 B.n76 585
R690 B.n676 B.n675 585
R691 B.n674 B.n77 585
R692 B.n673 B.n672 585
R693 B.n671 B.n78 585
R694 B.n670 B.n669 585
R695 B.n668 B.n79 585
R696 B.n667 B.n666 585
R697 B.n665 B.n80 585
R698 B.n664 B.n663 585
R699 B.n785 B.n36 585
R700 B.n787 B.n786 585
R701 B.n788 B.n35 585
R702 B.n790 B.n789 585
R703 B.n791 B.n34 585
R704 B.n793 B.n792 585
R705 B.n794 B.n33 585
R706 B.n796 B.n795 585
R707 B.n797 B.n32 585
R708 B.n799 B.n798 585
R709 B.n800 B.n31 585
R710 B.n802 B.n801 585
R711 B.n803 B.n30 585
R712 B.n805 B.n804 585
R713 B.n806 B.n29 585
R714 B.n808 B.n807 585
R715 B.n809 B.n28 585
R716 B.n811 B.n810 585
R717 B.n812 B.n27 585
R718 B.n814 B.n813 585
R719 B.n815 B.n26 585
R720 B.n817 B.n816 585
R721 B.n818 B.n25 585
R722 B.n820 B.n819 585
R723 B.n821 B.n24 585
R724 B.n823 B.n822 585
R725 B.n824 B.n23 585
R726 B.n826 B.n825 585
R727 B.n827 B.n22 585
R728 B.n829 B.n828 585
R729 B.n830 B.n21 585
R730 B.n832 B.n831 585
R731 B.n833 B.n20 585
R732 B.n835 B.n834 585
R733 B.n836 B.n19 585
R734 B.n838 B.n837 585
R735 B.n839 B.n18 585
R736 B.n841 B.n840 585
R737 B.n842 B.n17 585
R738 B.n844 B.n843 585
R739 B.n845 B.n16 585
R740 B.n847 B.n846 585
R741 B.n848 B.n15 585
R742 B.n850 B.n849 585
R743 B.n851 B.n14 585
R744 B.n853 B.n852 585
R745 B.n854 B.n13 585
R746 B.n856 B.n855 585
R747 B.n857 B.n12 585
R748 B.n859 B.n858 585
R749 B.n860 B.n11 585
R750 B.n862 B.n861 585
R751 B.n863 B.n10 585
R752 B.n865 B.n864 585
R753 B.n866 B.n9 585
R754 B.n868 B.n867 585
R755 B.n869 B.n8 585
R756 B.n871 B.n870 585
R757 B.n872 B.n7 585
R758 B.n874 B.n873 585
R759 B.n875 B.n6 585
R760 B.n877 B.n876 585
R761 B.n878 B.n5 585
R762 B.n880 B.n879 585
R763 B.n881 B.n4 585
R764 B.n883 B.n882 585
R765 B.n884 B.n3 585
R766 B.n886 B.n885 585
R767 B.n887 B.n0 585
R768 B.n2 B.n1 585
R769 B.n228 B.n227 585
R770 B.n229 B.n226 585
R771 B.n231 B.n230 585
R772 B.n232 B.n225 585
R773 B.n234 B.n233 585
R774 B.n235 B.n224 585
R775 B.n237 B.n236 585
R776 B.n238 B.n223 585
R777 B.n240 B.n239 585
R778 B.n241 B.n222 585
R779 B.n243 B.n242 585
R780 B.n244 B.n221 585
R781 B.n246 B.n245 585
R782 B.n247 B.n220 585
R783 B.n249 B.n248 585
R784 B.n250 B.n219 585
R785 B.n252 B.n251 585
R786 B.n253 B.n218 585
R787 B.n255 B.n254 585
R788 B.n256 B.n217 585
R789 B.n258 B.n257 585
R790 B.n259 B.n216 585
R791 B.n261 B.n260 585
R792 B.n262 B.n215 585
R793 B.n264 B.n263 585
R794 B.n265 B.n214 585
R795 B.n267 B.n266 585
R796 B.n268 B.n213 585
R797 B.n270 B.n269 585
R798 B.n271 B.n212 585
R799 B.n273 B.n272 585
R800 B.n274 B.n211 585
R801 B.n276 B.n275 585
R802 B.n277 B.n210 585
R803 B.n279 B.n278 585
R804 B.n280 B.n209 585
R805 B.n282 B.n281 585
R806 B.n283 B.n208 585
R807 B.n285 B.n284 585
R808 B.n286 B.n207 585
R809 B.n288 B.n287 585
R810 B.n289 B.n206 585
R811 B.n291 B.n290 585
R812 B.n292 B.n205 585
R813 B.n294 B.n293 585
R814 B.n295 B.n204 585
R815 B.n297 B.n296 585
R816 B.n298 B.n203 585
R817 B.n300 B.n299 585
R818 B.n301 B.n202 585
R819 B.n303 B.n302 585
R820 B.n304 B.n201 585
R821 B.n306 B.n305 585
R822 B.n307 B.n200 585
R823 B.n309 B.n308 585
R824 B.n310 B.n199 585
R825 B.n312 B.n311 585
R826 B.n313 B.n198 585
R827 B.n315 B.n314 585
R828 B.n316 B.n197 585
R829 B.n318 B.n317 585
R830 B.n319 B.n196 585
R831 B.n321 B.n320 585
R832 B.n322 B.n195 585
R833 B.n324 B.n323 585
R834 B.n325 B.n194 585
R835 B.n327 B.n326 585
R836 B.n328 B.n193 585
R837 B.n330 B.n193 530.939
R838 B.n454 B.n151 530.939
R839 B.n664 B.n81 530.939
R840 B.n785 B.n784 530.939
R841 B.n174 B.t3 283.654
R842 B.n396 B.t0 283.654
R843 B.n62 B.t6 283.654
R844 B.n54 B.t9 283.654
R845 B.n889 B.n888 256.663
R846 B.n888 B.n887 235.042
R847 B.n888 B.n2 235.042
R848 B.n396 B.t1 181.252
R849 B.n62 B.t8 181.252
R850 B.n174 B.t4 181.242
R851 B.n54 B.t11 181.242
R852 B.n331 B.n330 163.367
R853 B.n332 B.n331 163.367
R854 B.n332 B.n191 163.367
R855 B.n336 B.n191 163.367
R856 B.n337 B.n336 163.367
R857 B.n338 B.n337 163.367
R858 B.n338 B.n189 163.367
R859 B.n342 B.n189 163.367
R860 B.n343 B.n342 163.367
R861 B.n344 B.n343 163.367
R862 B.n344 B.n187 163.367
R863 B.n348 B.n187 163.367
R864 B.n349 B.n348 163.367
R865 B.n350 B.n349 163.367
R866 B.n350 B.n185 163.367
R867 B.n354 B.n185 163.367
R868 B.n355 B.n354 163.367
R869 B.n356 B.n355 163.367
R870 B.n356 B.n183 163.367
R871 B.n360 B.n183 163.367
R872 B.n361 B.n360 163.367
R873 B.n362 B.n361 163.367
R874 B.n362 B.n181 163.367
R875 B.n366 B.n181 163.367
R876 B.n367 B.n366 163.367
R877 B.n368 B.n367 163.367
R878 B.n368 B.n179 163.367
R879 B.n372 B.n179 163.367
R880 B.n373 B.n372 163.367
R881 B.n374 B.n373 163.367
R882 B.n374 B.n177 163.367
R883 B.n378 B.n177 163.367
R884 B.n379 B.n378 163.367
R885 B.n380 B.n379 163.367
R886 B.n380 B.n173 163.367
R887 B.n385 B.n173 163.367
R888 B.n386 B.n385 163.367
R889 B.n387 B.n386 163.367
R890 B.n387 B.n171 163.367
R891 B.n391 B.n171 163.367
R892 B.n392 B.n391 163.367
R893 B.n393 B.n392 163.367
R894 B.n393 B.n169 163.367
R895 B.n400 B.n169 163.367
R896 B.n401 B.n400 163.367
R897 B.n402 B.n401 163.367
R898 B.n402 B.n167 163.367
R899 B.n406 B.n167 163.367
R900 B.n407 B.n406 163.367
R901 B.n408 B.n407 163.367
R902 B.n408 B.n165 163.367
R903 B.n412 B.n165 163.367
R904 B.n413 B.n412 163.367
R905 B.n414 B.n413 163.367
R906 B.n414 B.n163 163.367
R907 B.n418 B.n163 163.367
R908 B.n419 B.n418 163.367
R909 B.n420 B.n419 163.367
R910 B.n420 B.n161 163.367
R911 B.n424 B.n161 163.367
R912 B.n425 B.n424 163.367
R913 B.n426 B.n425 163.367
R914 B.n426 B.n159 163.367
R915 B.n430 B.n159 163.367
R916 B.n431 B.n430 163.367
R917 B.n432 B.n431 163.367
R918 B.n432 B.n157 163.367
R919 B.n436 B.n157 163.367
R920 B.n437 B.n436 163.367
R921 B.n438 B.n437 163.367
R922 B.n438 B.n155 163.367
R923 B.n442 B.n155 163.367
R924 B.n443 B.n442 163.367
R925 B.n444 B.n443 163.367
R926 B.n444 B.n153 163.367
R927 B.n448 B.n153 163.367
R928 B.n449 B.n448 163.367
R929 B.n450 B.n449 163.367
R930 B.n450 B.n151 163.367
R931 B.n660 B.n81 163.367
R932 B.n660 B.n659 163.367
R933 B.n659 B.n658 163.367
R934 B.n658 B.n83 163.367
R935 B.n654 B.n83 163.367
R936 B.n654 B.n653 163.367
R937 B.n653 B.n652 163.367
R938 B.n652 B.n85 163.367
R939 B.n648 B.n85 163.367
R940 B.n648 B.n647 163.367
R941 B.n647 B.n646 163.367
R942 B.n646 B.n87 163.367
R943 B.n642 B.n87 163.367
R944 B.n642 B.n641 163.367
R945 B.n641 B.n640 163.367
R946 B.n640 B.n89 163.367
R947 B.n636 B.n89 163.367
R948 B.n636 B.n635 163.367
R949 B.n635 B.n634 163.367
R950 B.n634 B.n91 163.367
R951 B.n630 B.n91 163.367
R952 B.n630 B.n629 163.367
R953 B.n629 B.n628 163.367
R954 B.n628 B.n93 163.367
R955 B.n624 B.n93 163.367
R956 B.n624 B.n623 163.367
R957 B.n623 B.n622 163.367
R958 B.n622 B.n95 163.367
R959 B.n618 B.n95 163.367
R960 B.n618 B.n617 163.367
R961 B.n617 B.n616 163.367
R962 B.n616 B.n97 163.367
R963 B.n612 B.n97 163.367
R964 B.n612 B.n611 163.367
R965 B.n611 B.n610 163.367
R966 B.n610 B.n99 163.367
R967 B.n606 B.n99 163.367
R968 B.n606 B.n605 163.367
R969 B.n605 B.n604 163.367
R970 B.n604 B.n101 163.367
R971 B.n600 B.n101 163.367
R972 B.n600 B.n599 163.367
R973 B.n599 B.n598 163.367
R974 B.n598 B.n103 163.367
R975 B.n594 B.n103 163.367
R976 B.n594 B.n593 163.367
R977 B.n593 B.n592 163.367
R978 B.n592 B.n105 163.367
R979 B.n588 B.n105 163.367
R980 B.n588 B.n587 163.367
R981 B.n587 B.n586 163.367
R982 B.n586 B.n107 163.367
R983 B.n582 B.n107 163.367
R984 B.n582 B.n581 163.367
R985 B.n581 B.n580 163.367
R986 B.n580 B.n109 163.367
R987 B.n576 B.n109 163.367
R988 B.n576 B.n575 163.367
R989 B.n575 B.n574 163.367
R990 B.n574 B.n111 163.367
R991 B.n570 B.n111 163.367
R992 B.n570 B.n569 163.367
R993 B.n569 B.n568 163.367
R994 B.n568 B.n113 163.367
R995 B.n564 B.n113 163.367
R996 B.n564 B.n563 163.367
R997 B.n563 B.n562 163.367
R998 B.n562 B.n115 163.367
R999 B.n558 B.n115 163.367
R1000 B.n558 B.n557 163.367
R1001 B.n557 B.n556 163.367
R1002 B.n556 B.n117 163.367
R1003 B.n552 B.n117 163.367
R1004 B.n552 B.n551 163.367
R1005 B.n551 B.n550 163.367
R1006 B.n550 B.n119 163.367
R1007 B.n546 B.n119 163.367
R1008 B.n546 B.n545 163.367
R1009 B.n545 B.n544 163.367
R1010 B.n544 B.n121 163.367
R1011 B.n540 B.n121 163.367
R1012 B.n540 B.n539 163.367
R1013 B.n539 B.n538 163.367
R1014 B.n538 B.n123 163.367
R1015 B.n534 B.n123 163.367
R1016 B.n534 B.n533 163.367
R1017 B.n533 B.n532 163.367
R1018 B.n532 B.n125 163.367
R1019 B.n528 B.n125 163.367
R1020 B.n528 B.n527 163.367
R1021 B.n527 B.n526 163.367
R1022 B.n526 B.n127 163.367
R1023 B.n522 B.n127 163.367
R1024 B.n522 B.n521 163.367
R1025 B.n521 B.n520 163.367
R1026 B.n520 B.n129 163.367
R1027 B.n516 B.n129 163.367
R1028 B.n516 B.n515 163.367
R1029 B.n515 B.n514 163.367
R1030 B.n514 B.n131 163.367
R1031 B.n510 B.n131 163.367
R1032 B.n510 B.n509 163.367
R1033 B.n509 B.n508 163.367
R1034 B.n508 B.n133 163.367
R1035 B.n504 B.n133 163.367
R1036 B.n504 B.n503 163.367
R1037 B.n503 B.n502 163.367
R1038 B.n502 B.n135 163.367
R1039 B.n498 B.n135 163.367
R1040 B.n498 B.n497 163.367
R1041 B.n497 B.n496 163.367
R1042 B.n496 B.n137 163.367
R1043 B.n492 B.n137 163.367
R1044 B.n492 B.n491 163.367
R1045 B.n491 B.n490 163.367
R1046 B.n490 B.n139 163.367
R1047 B.n486 B.n139 163.367
R1048 B.n486 B.n485 163.367
R1049 B.n485 B.n484 163.367
R1050 B.n484 B.n141 163.367
R1051 B.n480 B.n141 163.367
R1052 B.n480 B.n479 163.367
R1053 B.n479 B.n478 163.367
R1054 B.n478 B.n143 163.367
R1055 B.n474 B.n143 163.367
R1056 B.n474 B.n473 163.367
R1057 B.n473 B.n472 163.367
R1058 B.n472 B.n145 163.367
R1059 B.n468 B.n145 163.367
R1060 B.n468 B.n467 163.367
R1061 B.n467 B.n466 163.367
R1062 B.n466 B.n147 163.367
R1063 B.n462 B.n147 163.367
R1064 B.n462 B.n461 163.367
R1065 B.n461 B.n460 163.367
R1066 B.n460 B.n149 163.367
R1067 B.n456 B.n149 163.367
R1068 B.n456 B.n455 163.367
R1069 B.n455 B.n454 163.367
R1070 B.n784 B.n37 163.367
R1071 B.n780 B.n37 163.367
R1072 B.n780 B.n779 163.367
R1073 B.n779 B.n778 163.367
R1074 B.n778 B.n39 163.367
R1075 B.n774 B.n39 163.367
R1076 B.n774 B.n773 163.367
R1077 B.n773 B.n772 163.367
R1078 B.n772 B.n41 163.367
R1079 B.n768 B.n41 163.367
R1080 B.n768 B.n767 163.367
R1081 B.n767 B.n766 163.367
R1082 B.n766 B.n43 163.367
R1083 B.n762 B.n43 163.367
R1084 B.n762 B.n761 163.367
R1085 B.n761 B.n760 163.367
R1086 B.n760 B.n45 163.367
R1087 B.n756 B.n45 163.367
R1088 B.n756 B.n755 163.367
R1089 B.n755 B.n754 163.367
R1090 B.n754 B.n47 163.367
R1091 B.n750 B.n47 163.367
R1092 B.n750 B.n749 163.367
R1093 B.n749 B.n748 163.367
R1094 B.n748 B.n49 163.367
R1095 B.n744 B.n49 163.367
R1096 B.n744 B.n743 163.367
R1097 B.n743 B.n742 163.367
R1098 B.n742 B.n51 163.367
R1099 B.n738 B.n51 163.367
R1100 B.n738 B.n737 163.367
R1101 B.n737 B.n736 163.367
R1102 B.n736 B.n53 163.367
R1103 B.n732 B.n53 163.367
R1104 B.n732 B.n731 163.367
R1105 B.n731 B.n57 163.367
R1106 B.n727 B.n57 163.367
R1107 B.n727 B.n726 163.367
R1108 B.n726 B.n725 163.367
R1109 B.n725 B.n59 163.367
R1110 B.n721 B.n59 163.367
R1111 B.n721 B.n720 163.367
R1112 B.n720 B.n719 163.367
R1113 B.n719 B.n61 163.367
R1114 B.n714 B.n61 163.367
R1115 B.n714 B.n713 163.367
R1116 B.n713 B.n712 163.367
R1117 B.n712 B.n65 163.367
R1118 B.n708 B.n65 163.367
R1119 B.n708 B.n707 163.367
R1120 B.n707 B.n706 163.367
R1121 B.n706 B.n67 163.367
R1122 B.n702 B.n67 163.367
R1123 B.n702 B.n701 163.367
R1124 B.n701 B.n700 163.367
R1125 B.n700 B.n69 163.367
R1126 B.n696 B.n69 163.367
R1127 B.n696 B.n695 163.367
R1128 B.n695 B.n694 163.367
R1129 B.n694 B.n71 163.367
R1130 B.n690 B.n71 163.367
R1131 B.n690 B.n689 163.367
R1132 B.n689 B.n688 163.367
R1133 B.n688 B.n73 163.367
R1134 B.n684 B.n73 163.367
R1135 B.n684 B.n683 163.367
R1136 B.n683 B.n682 163.367
R1137 B.n682 B.n75 163.367
R1138 B.n678 B.n75 163.367
R1139 B.n678 B.n677 163.367
R1140 B.n677 B.n676 163.367
R1141 B.n676 B.n77 163.367
R1142 B.n672 B.n77 163.367
R1143 B.n672 B.n671 163.367
R1144 B.n671 B.n670 163.367
R1145 B.n670 B.n79 163.367
R1146 B.n666 B.n79 163.367
R1147 B.n666 B.n665 163.367
R1148 B.n665 B.n664 163.367
R1149 B.n786 B.n785 163.367
R1150 B.n786 B.n35 163.367
R1151 B.n790 B.n35 163.367
R1152 B.n791 B.n790 163.367
R1153 B.n792 B.n791 163.367
R1154 B.n792 B.n33 163.367
R1155 B.n796 B.n33 163.367
R1156 B.n797 B.n796 163.367
R1157 B.n798 B.n797 163.367
R1158 B.n798 B.n31 163.367
R1159 B.n802 B.n31 163.367
R1160 B.n803 B.n802 163.367
R1161 B.n804 B.n803 163.367
R1162 B.n804 B.n29 163.367
R1163 B.n808 B.n29 163.367
R1164 B.n809 B.n808 163.367
R1165 B.n810 B.n809 163.367
R1166 B.n810 B.n27 163.367
R1167 B.n814 B.n27 163.367
R1168 B.n815 B.n814 163.367
R1169 B.n816 B.n815 163.367
R1170 B.n816 B.n25 163.367
R1171 B.n820 B.n25 163.367
R1172 B.n821 B.n820 163.367
R1173 B.n822 B.n821 163.367
R1174 B.n822 B.n23 163.367
R1175 B.n826 B.n23 163.367
R1176 B.n827 B.n826 163.367
R1177 B.n828 B.n827 163.367
R1178 B.n828 B.n21 163.367
R1179 B.n832 B.n21 163.367
R1180 B.n833 B.n832 163.367
R1181 B.n834 B.n833 163.367
R1182 B.n834 B.n19 163.367
R1183 B.n838 B.n19 163.367
R1184 B.n839 B.n838 163.367
R1185 B.n840 B.n839 163.367
R1186 B.n840 B.n17 163.367
R1187 B.n844 B.n17 163.367
R1188 B.n845 B.n844 163.367
R1189 B.n846 B.n845 163.367
R1190 B.n846 B.n15 163.367
R1191 B.n850 B.n15 163.367
R1192 B.n851 B.n850 163.367
R1193 B.n852 B.n851 163.367
R1194 B.n852 B.n13 163.367
R1195 B.n856 B.n13 163.367
R1196 B.n857 B.n856 163.367
R1197 B.n858 B.n857 163.367
R1198 B.n858 B.n11 163.367
R1199 B.n862 B.n11 163.367
R1200 B.n863 B.n862 163.367
R1201 B.n864 B.n863 163.367
R1202 B.n864 B.n9 163.367
R1203 B.n868 B.n9 163.367
R1204 B.n869 B.n868 163.367
R1205 B.n870 B.n869 163.367
R1206 B.n870 B.n7 163.367
R1207 B.n874 B.n7 163.367
R1208 B.n875 B.n874 163.367
R1209 B.n876 B.n875 163.367
R1210 B.n876 B.n5 163.367
R1211 B.n880 B.n5 163.367
R1212 B.n881 B.n880 163.367
R1213 B.n882 B.n881 163.367
R1214 B.n882 B.n3 163.367
R1215 B.n886 B.n3 163.367
R1216 B.n887 B.n886 163.367
R1217 B.n228 B.n2 163.367
R1218 B.n229 B.n228 163.367
R1219 B.n230 B.n229 163.367
R1220 B.n230 B.n225 163.367
R1221 B.n234 B.n225 163.367
R1222 B.n235 B.n234 163.367
R1223 B.n236 B.n235 163.367
R1224 B.n236 B.n223 163.367
R1225 B.n240 B.n223 163.367
R1226 B.n241 B.n240 163.367
R1227 B.n242 B.n241 163.367
R1228 B.n242 B.n221 163.367
R1229 B.n246 B.n221 163.367
R1230 B.n247 B.n246 163.367
R1231 B.n248 B.n247 163.367
R1232 B.n248 B.n219 163.367
R1233 B.n252 B.n219 163.367
R1234 B.n253 B.n252 163.367
R1235 B.n254 B.n253 163.367
R1236 B.n254 B.n217 163.367
R1237 B.n258 B.n217 163.367
R1238 B.n259 B.n258 163.367
R1239 B.n260 B.n259 163.367
R1240 B.n260 B.n215 163.367
R1241 B.n264 B.n215 163.367
R1242 B.n265 B.n264 163.367
R1243 B.n266 B.n265 163.367
R1244 B.n266 B.n213 163.367
R1245 B.n270 B.n213 163.367
R1246 B.n271 B.n270 163.367
R1247 B.n272 B.n271 163.367
R1248 B.n272 B.n211 163.367
R1249 B.n276 B.n211 163.367
R1250 B.n277 B.n276 163.367
R1251 B.n278 B.n277 163.367
R1252 B.n278 B.n209 163.367
R1253 B.n282 B.n209 163.367
R1254 B.n283 B.n282 163.367
R1255 B.n284 B.n283 163.367
R1256 B.n284 B.n207 163.367
R1257 B.n288 B.n207 163.367
R1258 B.n289 B.n288 163.367
R1259 B.n290 B.n289 163.367
R1260 B.n290 B.n205 163.367
R1261 B.n294 B.n205 163.367
R1262 B.n295 B.n294 163.367
R1263 B.n296 B.n295 163.367
R1264 B.n296 B.n203 163.367
R1265 B.n300 B.n203 163.367
R1266 B.n301 B.n300 163.367
R1267 B.n302 B.n301 163.367
R1268 B.n302 B.n201 163.367
R1269 B.n306 B.n201 163.367
R1270 B.n307 B.n306 163.367
R1271 B.n308 B.n307 163.367
R1272 B.n308 B.n199 163.367
R1273 B.n312 B.n199 163.367
R1274 B.n313 B.n312 163.367
R1275 B.n314 B.n313 163.367
R1276 B.n314 B.n197 163.367
R1277 B.n318 B.n197 163.367
R1278 B.n319 B.n318 163.367
R1279 B.n320 B.n319 163.367
R1280 B.n320 B.n195 163.367
R1281 B.n324 B.n195 163.367
R1282 B.n325 B.n324 163.367
R1283 B.n326 B.n325 163.367
R1284 B.n326 B.n193 163.367
R1285 B.n397 B.t2 113.567
R1286 B.n63 B.t7 113.567
R1287 B.n175 B.t5 113.556
R1288 B.n55 B.t10 113.556
R1289 B.n175 B.n174 67.6854
R1290 B.n397 B.n396 67.6854
R1291 B.n63 B.n62 67.6854
R1292 B.n55 B.n54 67.6854
R1293 B.n382 B.n175 59.5399
R1294 B.n398 B.n397 59.5399
R1295 B.n716 B.n63 59.5399
R1296 B.n56 B.n55 59.5399
R1297 B.n783 B.n36 34.4981
R1298 B.n663 B.n662 34.4981
R1299 B.n453 B.n452 34.4981
R1300 B.n329 B.n328 34.4981
R1301 B B.n889 18.0485
R1302 B.n787 B.n36 10.6151
R1303 B.n788 B.n787 10.6151
R1304 B.n789 B.n788 10.6151
R1305 B.n789 B.n34 10.6151
R1306 B.n793 B.n34 10.6151
R1307 B.n794 B.n793 10.6151
R1308 B.n795 B.n794 10.6151
R1309 B.n795 B.n32 10.6151
R1310 B.n799 B.n32 10.6151
R1311 B.n800 B.n799 10.6151
R1312 B.n801 B.n800 10.6151
R1313 B.n801 B.n30 10.6151
R1314 B.n805 B.n30 10.6151
R1315 B.n806 B.n805 10.6151
R1316 B.n807 B.n806 10.6151
R1317 B.n807 B.n28 10.6151
R1318 B.n811 B.n28 10.6151
R1319 B.n812 B.n811 10.6151
R1320 B.n813 B.n812 10.6151
R1321 B.n813 B.n26 10.6151
R1322 B.n817 B.n26 10.6151
R1323 B.n818 B.n817 10.6151
R1324 B.n819 B.n818 10.6151
R1325 B.n819 B.n24 10.6151
R1326 B.n823 B.n24 10.6151
R1327 B.n824 B.n823 10.6151
R1328 B.n825 B.n824 10.6151
R1329 B.n825 B.n22 10.6151
R1330 B.n829 B.n22 10.6151
R1331 B.n830 B.n829 10.6151
R1332 B.n831 B.n830 10.6151
R1333 B.n831 B.n20 10.6151
R1334 B.n835 B.n20 10.6151
R1335 B.n836 B.n835 10.6151
R1336 B.n837 B.n836 10.6151
R1337 B.n837 B.n18 10.6151
R1338 B.n841 B.n18 10.6151
R1339 B.n842 B.n841 10.6151
R1340 B.n843 B.n842 10.6151
R1341 B.n843 B.n16 10.6151
R1342 B.n847 B.n16 10.6151
R1343 B.n848 B.n847 10.6151
R1344 B.n849 B.n848 10.6151
R1345 B.n849 B.n14 10.6151
R1346 B.n853 B.n14 10.6151
R1347 B.n854 B.n853 10.6151
R1348 B.n855 B.n854 10.6151
R1349 B.n855 B.n12 10.6151
R1350 B.n859 B.n12 10.6151
R1351 B.n860 B.n859 10.6151
R1352 B.n861 B.n860 10.6151
R1353 B.n861 B.n10 10.6151
R1354 B.n865 B.n10 10.6151
R1355 B.n866 B.n865 10.6151
R1356 B.n867 B.n866 10.6151
R1357 B.n867 B.n8 10.6151
R1358 B.n871 B.n8 10.6151
R1359 B.n872 B.n871 10.6151
R1360 B.n873 B.n872 10.6151
R1361 B.n873 B.n6 10.6151
R1362 B.n877 B.n6 10.6151
R1363 B.n878 B.n877 10.6151
R1364 B.n879 B.n878 10.6151
R1365 B.n879 B.n4 10.6151
R1366 B.n883 B.n4 10.6151
R1367 B.n884 B.n883 10.6151
R1368 B.n885 B.n884 10.6151
R1369 B.n885 B.n0 10.6151
R1370 B.n783 B.n782 10.6151
R1371 B.n782 B.n781 10.6151
R1372 B.n781 B.n38 10.6151
R1373 B.n777 B.n38 10.6151
R1374 B.n777 B.n776 10.6151
R1375 B.n776 B.n775 10.6151
R1376 B.n775 B.n40 10.6151
R1377 B.n771 B.n40 10.6151
R1378 B.n771 B.n770 10.6151
R1379 B.n770 B.n769 10.6151
R1380 B.n769 B.n42 10.6151
R1381 B.n765 B.n42 10.6151
R1382 B.n765 B.n764 10.6151
R1383 B.n764 B.n763 10.6151
R1384 B.n763 B.n44 10.6151
R1385 B.n759 B.n44 10.6151
R1386 B.n759 B.n758 10.6151
R1387 B.n758 B.n757 10.6151
R1388 B.n757 B.n46 10.6151
R1389 B.n753 B.n46 10.6151
R1390 B.n753 B.n752 10.6151
R1391 B.n752 B.n751 10.6151
R1392 B.n751 B.n48 10.6151
R1393 B.n747 B.n48 10.6151
R1394 B.n747 B.n746 10.6151
R1395 B.n746 B.n745 10.6151
R1396 B.n745 B.n50 10.6151
R1397 B.n741 B.n50 10.6151
R1398 B.n741 B.n740 10.6151
R1399 B.n740 B.n739 10.6151
R1400 B.n739 B.n52 10.6151
R1401 B.n735 B.n52 10.6151
R1402 B.n735 B.n734 10.6151
R1403 B.n734 B.n733 10.6151
R1404 B.n730 B.n729 10.6151
R1405 B.n729 B.n728 10.6151
R1406 B.n728 B.n58 10.6151
R1407 B.n724 B.n58 10.6151
R1408 B.n724 B.n723 10.6151
R1409 B.n723 B.n722 10.6151
R1410 B.n722 B.n60 10.6151
R1411 B.n718 B.n60 10.6151
R1412 B.n718 B.n717 10.6151
R1413 B.n715 B.n64 10.6151
R1414 B.n711 B.n64 10.6151
R1415 B.n711 B.n710 10.6151
R1416 B.n710 B.n709 10.6151
R1417 B.n709 B.n66 10.6151
R1418 B.n705 B.n66 10.6151
R1419 B.n705 B.n704 10.6151
R1420 B.n704 B.n703 10.6151
R1421 B.n703 B.n68 10.6151
R1422 B.n699 B.n68 10.6151
R1423 B.n699 B.n698 10.6151
R1424 B.n698 B.n697 10.6151
R1425 B.n697 B.n70 10.6151
R1426 B.n693 B.n70 10.6151
R1427 B.n693 B.n692 10.6151
R1428 B.n692 B.n691 10.6151
R1429 B.n691 B.n72 10.6151
R1430 B.n687 B.n72 10.6151
R1431 B.n687 B.n686 10.6151
R1432 B.n686 B.n685 10.6151
R1433 B.n685 B.n74 10.6151
R1434 B.n681 B.n74 10.6151
R1435 B.n681 B.n680 10.6151
R1436 B.n680 B.n679 10.6151
R1437 B.n679 B.n76 10.6151
R1438 B.n675 B.n76 10.6151
R1439 B.n675 B.n674 10.6151
R1440 B.n674 B.n673 10.6151
R1441 B.n673 B.n78 10.6151
R1442 B.n669 B.n78 10.6151
R1443 B.n669 B.n668 10.6151
R1444 B.n668 B.n667 10.6151
R1445 B.n667 B.n80 10.6151
R1446 B.n663 B.n80 10.6151
R1447 B.n662 B.n661 10.6151
R1448 B.n661 B.n82 10.6151
R1449 B.n657 B.n82 10.6151
R1450 B.n657 B.n656 10.6151
R1451 B.n656 B.n655 10.6151
R1452 B.n655 B.n84 10.6151
R1453 B.n651 B.n84 10.6151
R1454 B.n651 B.n650 10.6151
R1455 B.n650 B.n649 10.6151
R1456 B.n649 B.n86 10.6151
R1457 B.n645 B.n86 10.6151
R1458 B.n645 B.n644 10.6151
R1459 B.n644 B.n643 10.6151
R1460 B.n643 B.n88 10.6151
R1461 B.n639 B.n88 10.6151
R1462 B.n639 B.n638 10.6151
R1463 B.n638 B.n637 10.6151
R1464 B.n637 B.n90 10.6151
R1465 B.n633 B.n90 10.6151
R1466 B.n633 B.n632 10.6151
R1467 B.n632 B.n631 10.6151
R1468 B.n631 B.n92 10.6151
R1469 B.n627 B.n92 10.6151
R1470 B.n627 B.n626 10.6151
R1471 B.n626 B.n625 10.6151
R1472 B.n625 B.n94 10.6151
R1473 B.n621 B.n94 10.6151
R1474 B.n621 B.n620 10.6151
R1475 B.n620 B.n619 10.6151
R1476 B.n619 B.n96 10.6151
R1477 B.n615 B.n96 10.6151
R1478 B.n615 B.n614 10.6151
R1479 B.n614 B.n613 10.6151
R1480 B.n613 B.n98 10.6151
R1481 B.n609 B.n98 10.6151
R1482 B.n609 B.n608 10.6151
R1483 B.n608 B.n607 10.6151
R1484 B.n607 B.n100 10.6151
R1485 B.n603 B.n100 10.6151
R1486 B.n603 B.n602 10.6151
R1487 B.n602 B.n601 10.6151
R1488 B.n601 B.n102 10.6151
R1489 B.n597 B.n102 10.6151
R1490 B.n597 B.n596 10.6151
R1491 B.n596 B.n595 10.6151
R1492 B.n595 B.n104 10.6151
R1493 B.n591 B.n104 10.6151
R1494 B.n591 B.n590 10.6151
R1495 B.n590 B.n589 10.6151
R1496 B.n589 B.n106 10.6151
R1497 B.n585 B.n106 10.6151
R1498 B.n585 B.n584 10.6151
R1499 B.n584 B.n583 10.6151
R1500 B.n583 B.n108 10.6151
R1501 B.n579 B.n108 10.6151
R1502 B.n579 B.n578 10.6151
R1503 B.n578 B.n577 10.6151
R1504 B.n577 B.n110 10.6151
R1505 B.n573 B.n110 10.6151
R1506 B.n573 B.n572 10.6151
R1507 B.n572 B.n571 10.6151
R1508 B.n571 B.n112 10.6151
R1509 B.n567 B.n112 10.6151
R1510 B.n567 B.n566 10.6151
R1511 B.n566 B.n565 10.6151
R1512 B.n565 B.n114 10.6151
R1513 B.n561 B.n114 10.6151
R1514 B.n561 B.n560 10.6151
R1515 B.n560 B.n559 10.6151
R1516 B.n559 B.n116 10.6151
R1517 B.n555 B.n116 10.6151
R1518 B.n555 B.n554 10.6151
R1519 B.n554 B.n553 10.6151
R1520 B.n553 B.n118 10.6151
R1521 B.n549 B.n118 10.6151
R1522 B.n549 B.n548 10.6151
R1523 B.n548 B.n547 10.6151
R1524 B.n547 B.n120 10.6151
R1525 B.n543 B.n120 10.6151
R1526 B.n543 B.n542 10.6151
R1527 B.n542 B.n541 10.6151
R1528 B.n541 B.n122 10.6151
R1529 B.n537 B.n122 10.6151
R1530 B.n537 B.n536 10.6151
R1531 B.n536 B.n535 10.6151
R1532 B.n535 B.n124 10.6151
R1533 B.n531 B.n124 10.6151
R1534 B.n531 B.n530 10.6151
R1535 B.n530 B.n529 10.6151
R1536 B.n529 B.n126 10.6151
R1537 B.n525 B.n126 10.6151
R1538 B.n525 B.n524 10.6151
R1539 B.n524 B.n523 10.6151
R1540 B.n523 B.n128 10.6151
R1541 B.n519 B.n128 10.6151
R1542 B.n519 B.n518 10.6151
R1543 B.n518 B.n517 10.6151
R1544 B.n517 B.n130 10.6151
R1545 B.n513 B.n130 10.6151
R1546 B.n513 B.n512 10.6151
R1547 B.n512 B.n511 10.6151
R1548 B.n511 B.n132 10.6151
R1549 B.n507 B.n132 10.6151
R1550 B.n507 B.n506 10.6151
R1551 B.n506 B.n505 10.6151
R1552 B.n505 B.n134 10.6151
R1553 B.n501 B.n134 10.6151
R1554 B.n501 B.n500 10.6151
R1555 B.n500 B.n499 10.6151
R1556 B.n499 B.n136 10.6151
R1557 B.n495 B.n136 10.6151
R1558 B.n495 B.n494 10.6151
R1559 B.n494 B.n493 10.6151
R1560 B.n493 B.n138 10.6151
R1561 B.n489 B.n138 10.6151
R1562 B.n489 B.n488 10.6151
R1563 B.n488 B.n487 10.6151
R1564 B.n487 B.n140 10.6151
R1565 B.n483 B.n140 10.6151
R1566 B.n483 B.n482 10.6151
R1567 B.n482 B.n481 10.6151
R1568 B.n481 B.n142 10.6151
R1569 B.n477 B.n142 10.6151
R1570 B.n477 B.n476 10.6151
R1571 B.n476 B.n475 10.6151
R1572 B.n475 B.n144 10.6151
R1573 B.n471 B.n144 10.6151
R1574 B.n471 B.n470 10.6151
R1575 B.n470 B.n469 10.6151
R1576 B.n469 B.n146 10.6151
R1577 B.n465 B.n146 10.6151
R1578 B.n465 B.n464 10.6151
R1579 B.n464 B.n463 10.6151
R1580 B.n463 B.n148 10.6151
R1581 B.n459 B.n148 10.6151
R1582 B.n459 B.n458 10.6151
R1583 B.n458 B.n457 10.6151
R1584 B.n457 B.n150 10.6151
R1585 B.n453 B.n150 10.6151
R1586 B.n227 B.n1 10.6151
R1587 B.n227 B.n226 10.6151
R1588 B.n231 B.n226 10.6151
R1589 B.n232 B.n231 10.6151
R1590 B.n233 B.n232 10.6151
R1591 B.n233 B.n224 10.6151
R1592 B.n237 B.n224 10.6151
R1593 B.n238 B.n237 10.6151
R1594 B.n239 B.n238 10.6151
R1595 B.n239 B.n222 10.6151
R1596 B.n243 B.n222 10.6151
R1597 B.n244 B.n243 10.6151
R1598 B.n245 B.n244 10.6151
R1599 B.n245 B.n220 10.6151
R1600 B.n249 B.n220 10.6151
R1601 B.n250 B.n249 10.6151
R1602 B.n251 B.n250 10.6151
R1603 B.n251 B.n218 10.6151
R1604 B.n255 B.n218 10.6151
R1605 B.n256 B.n255 10.6151
R1606 B.n257 B.n256 10.6151
R1607 B.n257 B.n216 10.6151
R1608 B.n261 B.n216 10.6151
R1609 B.n262 B.n261 10.6151
R1610 B.n263 B.n262 10.6151
R1611 B.n263 B.n214 10.6151
R1612 B.n267 B.n214 10.6151
R1613 B.n268 B.n267 10.6151
R1614 B.n269 B.n268 10.6151
R1615 B.n269 B.n212 10.6151
R1616 B.n273 B.n212 10.6151
R1617 B.n274 B.n273 10.6151
R1618 B.n275 B.n274 10.6151
R1619 B.n275 B.n210 10.6151
R1620 B.n279 B.n210 10.6151
R1621 B.n280 B.n279 10.6151
R1622 B.n281 B.n280 10.6151
R1623 B.n281 B.n208 10.6151
R1624 B.n285 B.n208 10.6151
R1625 B.n286 B.n285 10.6151
R1626 B.n287 B.n286 10.6151
R1627 B.n287 B.n206 10.6151
R1628 B.n291 B.n206 10.6151
R1629 B.n292 B.n291 10.6151
R1630 B.n293 B.n292 10.6151
R1631 B.n293 B.n204 10.6151
R1632 B.n297 B.n204 10.6151
R1633 B.n298 B.n297 10.6151
R1634 B.n299 B.n298 10.6151
R1635 B.n299 B.n202 10.6151
R1636 B.n303 B.n202 10.6151
R1637 B.n304 B.n303 10.6151
R1638 B.n305 B.n304 10.6151
R1639 B.n305 B.n200 10.6151
R1640 B.n309 B.n200 10.6151
R1641 B.n310 B.n309 10.6151
R1642 B.n311 B.n310 10.6151
R1643 B.n311 B.n198 10.6151
R1644 B.n315 B.n198 10.6151
R1645 B.n316 B.n315 10.6151
R1646 B.n317 B.n316 10.6151
R1647 B.n317 B.n196 10.6151
R1648 B.n321 B.n196 10.6151
R1649 B.n322 B.n321 10.6151
R1650 B.n323 B.n322 10.6151
R1651 B.n323 B.n194 10.6151
R1652 B.n327 B.n194 10.6151
R1653 B.n328 B.n327 10.6151
R1654 B.n329 B.n192 10.6151
R1655 B.n333 B.n192 10.6151
R1656 B.n334 B.n333 10.6151
R1657 B.n335 B.n334 10.6151
R1658 B.n335 B.n190 10.6151
R1659 B.n339 B.n190 10.6151
R1660 B.n340 B.n339 10.6151
R1661 B.n341 B.n340 10.6151
R1662 B.n341 B.n188 10.6151
R1663 B.n345 B.n188 10.6151
R1664 B.n346 B.n345 10.6151
R1665 B.n347 B.n346 10.6151
R1666 B.n347 B.n186 10.6151
R1667 B.n351 B.n186 10.6151
R1668 B.n352 B.n351 10.6151
R1669 B.n353 B.n352 10.6151
R1670 B.n353 B.n184 10.6151
R1671 B.n357 B.n184 10.6151
R1672 B.n358 B.n357 10.6151
R1673 B.n359 B.n358 10.6151
R1674 B.n359 B.n182 10.6151
R1675 B.n363 B.n182 10.6151
R1676 B.n364 B.n363 10.6151
R1677 B.n365 B.n364 10.6151
R1678 B.n365 B.n180 10.6151
R1679 B.n369 B.n180 10.6151
R1680 B.n370 B.n369 10.6151
R1681 B.n371 B.n370 10.6151
R1682 B.n371 B.n178 10.6151
R1683 B.n375 B.n178 10.6151
R1684 B.n376 B.n375 10.6151
R1685 B.n377 B.n376 10.6151
R1686 B.n377 B.n176 10.6151
R1687 B.n381 B.n176 10.6151
R1688 B.n384 B.n383 10.6151
R1689 B.n384 B.n172 10.6151
R1690 B.n388 B.n172 10.6151
R1691 B.n389 B.n388 10.6151
R1692 B.n390 B.n389 10.6151
R1693 B.n390 B.n170 10.6151
R1694 B.n394 B.n170 10.6151
R1695 B.n395 B.n394 10.6151
R1696 B.n399 B.n395 10.6151
R1697 B.n403 B.n168 10.6151
R1698 B.n404 B.n403 10.6151
R1699 B.n405 B.n404 10.6151
R1700 B.n405 B.n166 10.6151
R1701 B.n409 B.n166 10.6151
R1702 B.n410 B.n409 10.6151
R1703 B.n411 B.n410 10.6151
R1704 B.n411 B.n164 10.6151
R1705 B.n415 B.n164 10.6151
R1706 B.n416 B.n415 10.6151
R1707 B.n417 B.n416 10.6151
R1708 B.n417 B.n162 10.6151
R1709 B.n421 B.n162 10.6151
R1710 B.n422 B.n421 10.6151
R1711 B.n423 B.n422 10.6151
R1712 B.n423 B.n160 10.6151
R1713 B.n427 B.n160 10.6151
R1714 B.n428 B.n427 10.6151
R1715 B.n429 B.n428 10.6151
R1716 B.n429 B.n158 10.6151
R1717 B.n433 B.n158 10.6151
R1718 B.n434 B.n433 10.6151
R1719 B.n435 B.n434 10.6151
R1720 B.n435 B.n156 10.6151
R1721 B.n439 B.n156 10.6151
R1722 B.n440 B.n439 10.6151
R1723 B.n441 B.n440 10.6151
R1724 B.n441 B.n154 10.6151
R1725 B.n445 B.n154 10.6151
R1726 B.n446 B.n445 10.6151
R1727 B.n447 B.n446 10.6151
R1728 B.n447 B.n152 10.6151
R1729 B.n451 B.n152 10.6151
R1730 B.n452 B.n451 10.6151
R1731 B.n733 B.n56 9.36635
R1732 B.n716 B.n715 9.36635
R1733 B.n382 B.n381 9.36635
R1734 B.n398 B.n168 9.36635
R1735 B.n889 B.n0 8.11757
R1736 B.n889 B.n1 8.11757
R1737 B.n730 B.n56 1.24928
R1738 B.n717 B.n716 1.24928
R1739 B.n383 B.n382 1.24928
R1740 B.n399 B.n398 1.24928
C0 VTAIL VP 10.149099f
C1 VDD2 VN 9.15191f
C2 VTAIL VN 10.1349f
C3 VDD1 B 2.52461f
C4 VDD2 VDD1 2.53614f
C5 VTAIL VDD1 9.686231f
C6 w_n5158_n2932# B 10.8773f
C7 w_n5158_n2932# VDD2 3.01786f
C8 w_n5158_n2932# VTAIL 2.97864f
C9 VP VN 8.83389f
C10 VDD2 B 2.66433f
C11 VTAIL B 3.44671f
C12 VDD2 VTAIL 9.74187f
C13 VP VDD1 9.648581f
C14 VDD1 VN 0.153909f
C15 w_n5158_n2932# VP 11.8728f
C16 w_n5158_n2932# VN 11.199599f
C17 VP B 2.53114f
C18 VN B 1.3959f
C19 w_n5158_n2932# VDD1 2.8452f
C20 VDD2 VP 0.654144f
C21 VDD2 VSUBS 2.332974f
C22 VDD1 VSUBS 2.137478f
C23 VTAIL VSUBS 1.36815f
C24 VN VSUBS 8.57477f
C25 VP VSUBS 4.87314f
C26 B VSUBS 5.87788f
C27 w_n5158_n2932# VSUBS 0.186864p
C28 B.n0 VSUBS 0.008598f
C29 B.n1 VSUBS 0.008598f
C30 B.n2 VSUBS 0.012715f
C31 B.n3 VSUBS 0.009744f
C32 B.n4 VSUBS 0.009744f
C33 B.n5 VSUBS 0.009744f
C34 B.n6 VSUBS 0.009744f
C35 B.n7 VSUBS 0.009744f
C36 B.n8 VSUBS 0.009744f
C37 B.n9 VSUBS 0.009744f
C38 B.n10 VSUBS 0.009744f
C39 B.n11 VSUBS 0.009744f
C40 B.n12 VSUBS 0.009744f
C41 B.n13 VSUBS 0.009744f
C42 B.n14 VSUBS 0.009744f
C43 B.n15 VSUBS 0.009744f
C44 B.n16 VSUBS 0.009744f
C45 B.n17 VSUBS 0.009744f
C46 B.n18 VSUBS 0.009744f
C47 B.n19 VSUBS 0.009744f
C48 B.n20 VSUBS 0.009744f
C49 B.n21 VSUBS 0.009744f
C50 B.n22 VSUBS 0.009744f
C51 B.n23 VSUBS 0.009744f
C52 B.n24 VSUBS 0.009744f
C53 B.n25 VSUBS 0.009744f
C54 B.n26 VSUBS 0.009744f
C55 B.n27 VSUBS 0.009744f
C56 B.n28 VSUBS 0.009744f
C57 B.n29 VSUBS 0.009744f
C58 B.n30 VSUBS 0.009744f
C59 B.n31 VSUBS 0.009744f
C60 B.n32 VSUBS 0.009744f
C61 B.n33 VSUBS 0.009744f
C62 B.n34 VSUBS 0.009744f
C63 B.n35 VSUBS 0.009744f
C64 B.n36 VSUBS 0.022939f
C65 B.n37 VSUBS 0.009744f
C66 B.n38 VSUBS 0.009744f
C67 B.n39 VSUBS 0.009744f
C68 B.n40 VSUBS 0.009744f
C69 B.n41 VSUBS 0.009744f
C70 B.n42 VSUBS 0.009744f
C71 B.n43 VSUBS 0.009744f
C72 B.n44 VSUBS 0.009744f
C73 B.n45 VSUBS 0.009744f
C74 B.n46 VSUBS 0.009744f
C75 B.n47 VSUBS 0.009744f
C76 B.n48 VSUBS 0.009744f
C77 B.n49 VSUBS 0.009744f
C78 B.n50 VSUBS 0.009744f
C79 B.n51 VSUBS 0.009744f
C80 B.n52 VSUBS 0.009744f
C81 B.n53 VSUBS 0.009744f
C82 B.t10 VSUBS 0.434859f
C83 B.t11 VSUBS 0.468117f
C84 B.t9 VSUBS 2.01461f
C85 B.n54 VSUBS 0.258116f
C86 B.n55 VSUBS 0.102954f
C87 B.n56 VSUBS 0.022576f
C88 B.n57 VSUBS 0.009744f
C89 B.n58 VSUBS 0.009744f
C90 B.n59 VSUBS 0.009744f
C91 B.n60 VSUBS 0.009744f
C92 B.n61 VSUBS 0.009744f
C93 B.t7 VSUBS 0.434853f
C94 B.t8 VSUBS 0.468112f
C95 B.t6 VSUBS 2.01461f
C96 B.n62 VSUBS 0.258121f
C97 B.n63 VSUBS 0.10296f
C98 B.n64 VSUBS 0.009744f
C99 B.n65 VSUBS 0.009744f
C100 B.n66 VSUBS 0.009744f
C101 B.n67 VSUBS 0.009744f
C102 B.n68 VSUBS 0.009744f
C103 B.n69 VSUBS 0.009744f
C104 B.n70 VSUBS 0.009744f
C105 B.n71 VSUBS 0.009744f
C106 B.n72 VSUBS 0.009744f
C107 B.n73 VSUBS 0.009744f
C108 B.n74 VSUBS 0.009744f
C109 B.n75 VSUBS 0.009744f
C110 B.n76 VSUBS 0.009744f
C111 B.n77 VSUBS 0.009744f
C112 B.n78 VSUBS 0.009744f
C113 B.n79 VSUBS 0.009744f
C114 B.n80 VSUBS 0.009744f
C115 B.n81 VSUBS 0.022939f
C116 B.n82 VSUBS 0.009744f
C117 B.n83 VSUBS 0.009744f
C118 B.n84 VSUBS 0.009744f
C119 B.n85 VSUBS 0.009744f
C120 B.n86 VSUBS 0.009744f
C121 B.n87 VSUBS 0.009744f
C122 B.n88 VSUBS 0.009744f
C123 B.n89 VSUBS 0.009744f
C124 B.n90 VSUBS 0.009744f
C125 B.n91 VSUBS 0.009744f
C126 B.n92 VSUBS 0.009744f
C127 B.n93 VSUBS 0.009744f
C128 B.n94 VSUBS 0.009744f
C129 B.n95 VSUBS 0.009744f
C130 B.n96 VSUBS 0.009744f
C131 B.n97 VSUBS 0.009744f
C132 B.n98 VSUBS 0.009744f
C133 B.n99 VSUBS 0.009744f
C134 B.n100 VSUBS 0.009744f
C135 B.n101 VSUBS 0.009744f
C136 B.n102 VSUBS 0.009744f
C137 B.n103 VSUBS 0.009744f
C138 B.n104 VSUBS 0.009744f
C139 B.n105 VSUBS 0.009744f
C140 B.n106 VSUBS 0.009744f
C141 B.n107 VSUBS 0.009744f
C142 B.n108 VSUBS 0.009744f
C143 B.n109 VSUBS 0.009744f
C144 B.n110 VSUBS 0.009744f
C145 B.n111 VSUBS 0.009744f
C146 B.n112 VSUBS 0.009744f
C147 B.n113 VSUBS 0.009744f
C148 B.n114 VSUBS 0.009744f
C149 B.n115 VSUBS 0.009744f
C150 B.n116 VSUBS 0.009744f
C151 B.n117 VSUBS 0.009744f
C152 B.n118 VSUBS 0.009744f
C153 B.n119 VSUBS 0.009744f
C154 B.n120 VSUBS 0.009744f
C155 B.n121 VSUBS 0.009744f
C156 B.n122 VSUBS 0.009744f
C157 B.n123 VSUBS 0.009744f
C158 B.n124 VSUBS 0.009744f
C159 B.n125 VSUBS 0.009744f
C160 B.n126 VSUBS 0.009744f
C161 B.n127 VSUBS 0.009744f
C162 B.n128 VSUBS 0.009744f
C163 B.n129 VSUBS 0.009744f
C164 B.n130 VSUBS 0.009744f
C165 B.n131 VSUBS 0.009744f
C166 B.n132 VSUBS 0.009744f
C167 B.n133 VSUBS 0.009744f
C168 B.n134 VSUBS 0.009744f
C169 B.n135 VSUBS 0.009744f
C170 B.n136 VSUBS 0.009744f
C171 B.n137 VSUBS 0.009744f
C172 B.n138 VSUBS 0.009744f
C173 B.n139 VSUBS 0.009744f
C174 B.n140 VSUBS 0.009744f
C175 B.n141 VSUBS 0.009744f
C176 B.n142 VSUBS 0.009744f
C177 B.n143 VSUBS 0.009744f
C178 B.n144 VSUBS 0.009744f
C179 B.n145 VSUBS 0.009744f
C180 B.n146 VSUBS 0.009744f
C181 B.n147 VSUBS 0.009744f
C182 B.n148 VSUBS 0.009744f
C183 B.n149 VSUBS 0.009744f
C184 B.n150 VSUBS 0.009744f
C185 B.n151 VSUBS 0.024348f
C186 B.n152 VSUBS 0.009744f
C187 B.n153 VSUBS 0.009744f
C188 B.n154 VSUBS 0.009744f
C189 B.n155 VSUBS 0.009744f
C190 B.n156 VSUBS 0.009744f
C191 B.n157 VSUBS 0.009744f
C192 B.n158 VSUBS 0.009744f
C193 B.n159 VSUBS 0.009744f
C194 B.n160 VSUBS 0.009744f
C195 B.n161 VSUBS 0.009744f
C196 B.n162 VSUBS 0.009744f
C197 B.n163 VSUBS 0.009744f
C198 B.n164 VSUBS 0.009744f
C199 B.n165 VSUBS 0.009744f
C200 B.n166 VSUBS 0.009744f
C201 B.n167 VSUBS 0.009744f
C202 B.n168 VSUBS 0.009171f
C203 B.n169 VSUBS 0.009744f
C204 B.n170 VSUBS 0.009744f
C205 B.n171 VSUBS 0.009744f
C206 B.n172 VSUBS 0.009744f
C207 B.n173 VSUBS 0.009744f
C208 B.t5 VSUBS 0.434859f
C209 B.t4 VSUBS 0.468117f
C210 B.t3 VSUBS 2.01461f
C211 B.n174 VSUBS 0.258116f
C212 B.n175 VSUBS 0.102954f
C213 B.n176 VSUBS 0.009744f
C214 B.n177 VSUBS 0.009744f
C215 B.n178 VSUBS 0.009744f
C216 B.n179 VSUBS 0.009744f
C217 B.n180 VSUBS 0.009744f
C218 B.n181 VSUBS 0.009744f
C219 B.n182 VSUBS 0.009744f
C220 B.n183 VSUBS 0.009744f
C221 B.n184 VSUBS 0.009744f
C222 B.n185 VSUBS 0.009744f
C223 B.n186 VSUBS 0.009744f
C224 B.n187 VSUBS 0.009744f
C225 B.n188 VSUBS 0.009744f
C226 B.n189 VSUBS 0.009744f
C227 B.n190 VSUBS 0.009744f
C228 B.n191 VSUBS 0.009744f
C229 B.n192 VSUBS 0.009744f
C230 B.n193 VSUBS 0.022939f
C231 B.n194 VSUBS 0.009744f
C232 B.n195 VSUBS 0.009744f
C233 B.n196 VSUBS 0.009744f
C234 B.n197 VSUBS 0.009744f
C235 B.n198 VSUBS 0.009744f
C236 B.n199 VSUBS 0.009744f
C237 B.n200 VSUBS 0.009744f
C238 B.n201 VSUBS 0.009744f
C239 B.n202 VSUBS 0.009744f
C240 B.n203 VSUBS 0.009744f
C241 B.n204 VSUBS 0.009744f
C242 B.n205 VSUBS 0.009744f
C243 B.n206 VSUBS 0.009744f
C244 B.n207 VSUBS 0.009744f
C245 B.n208 VSUBS 0.009744f
C246 B.n209 VSUBS 0.009744f
C247 B.n210 VSUBS 0.009744f
C248 B.n211 VSUBS 0.009744f
C249 B.n212 VSUBS 0.009744f
C250 B.n213 VSUBS 0.009744f
C251 B.n214 VSUBS 0.009744f
C252 B.n215 VSUBS 0.009744f
C253 B.n216 VSUBS 0.009744f
C254 B.n217 VSUBS 0.009744f
C255 B.n218 VSUBS 0.009744f
C256 B.n219 VSUBS 0.009744f
C257 B.n220 VSUBS 0.009744f
C258 B.n221 VSUBS 0.009744f
C259 B.n222 VSUBS 0.009744f
C260 B.n223 VSUBS 0.009744f
C261 B.n224 VSUBS 0.009744f
C262 B.n225 VSUBS 0.009744f
C263 B.n226 VSUBS 0.009744f
C264 B.n227 VSUBS 0.009744f
C265 B.n228 VSUBS 0.009744f
C266 B.n229 VSUBS 0.009744f
C267 B.n230 VSUBS 0.009744f
C268 B.n231 VSUBS 0.009744f
C269 B.n232 VSUBS 0.009744f
C270 B.n233 VSUBS 0.009744f
C271 B.n234 VSUBS 0.009744f
C272 B.n235 VSUBS 0.009744f
C273 B.n236 VSUBS 0.009744f
C274 B.n237 VSUBS 0.009744f
C275 B.n238 VSUBS 0.009744f
C276 B.n239 VSUBS 0.009744f
C277 B.n240 VSUBS 0.009744f
C278 B.n241 VSUBS 0.009744f
C279 B.n242 VSUBS 0.009744f
C280 B.n243 VSUBS 0.009744f
C281 B.n244 VSUBS 0.009744f
C282 B.n245 VSUBS 0.009744f
C283 B.n246 VSUBS 0.009744f
C284 B.n247 VSUBS 0.009744f
C285 B.n248 VSUBS 0.009744f
C286 B.n249 VSUBS 0.009744f
C287 B.n250 VSUBS 0.009744f
C288 B.n251 VSUBS 0.009744f
C289 B.n252 VSUBS 0.009744f
C290 B.n253 VSUBS 0.009744f
C291 B.n254 VSUBS 0.009744f
C292 B.n255 VSUBS 0.009744f
C293 B.n256 VSUBS 0.009744f
C294 B.n257 VSUBS 0.009744f
C295 B.n258 VSUBS 0.009744f
C296 B.n259 VSUBS 0.009744f
C297 B.n260 VSUBS 0.009744f
C298 B.n261 VSUBS 0.009744f
C299 B.n262 VSUBS 0.009744f
C300 B.n263 VSUBS 0.009744f
C301 B.n264 VSUBS 0.009744f
C302 B.n265 VSUBS 0.009744f
C303 B.n266 VSUBS 0.009744f
C304 B.n267 VSUBS 0.009744f
C305 B.n268 VSUBS 0.009744f
C306 B.n269 VSUBS 0.009744f
C307 B.n270 VSUBS 0.009744f
C308 B.n271 VSUBS 0.009744f
C309 B.n272 VSUBS 0.009744f
C310 B.n273 VSUBS 0.009744f
C311 B.n274 VSUBS 0.009744f
C312 B.n275 VSUBS 0.009744f
C313 B.n276 VSUBS 0.009744f
C314 B.n277 VSUBS 0.009744f
C315 B.n278 VSUBS 0.009744f
C316 B.n279 VSUBS 0.009744f
C317 B.n280 VSUBS 0.009744f
C318 B.n281 VSUBS 0.009744f
C319 B.n282 VSUBS 0.009744f
C320 B.n283 VSUBS 0.009744f
C321 B.n284 VSUBS 0.009744f
C322 B.n285 VSUBS 0.009744f
C323 B.n286 VSUBS 0.009744f
C324 B.n287 VSUBS 0.009744f
C325 B.n288 VSUBS 0.009744f
C326 B.n289 VSUBS 0.009744f
C327 B.n290 VSUBS 0.009744f
C328 B.n291 VSUBS 0.009744f
C329 B.n292 VSUBS 0.009744f
C330 B.n293 VSUBS 0.009744f
C331 B.n294 VSUBS 0.009744f
C332 B.n295 VSUBS 0.009744f
C333 B.n296 VSUBS 0.009744f
C334 B.n297 VSUBS 0.009744f
C335 B.n298 VSUBS 0.009744f
C336 B.n299 VSUBS 0.009744f
C337 B.n300 VSUBS 0.009744f
C338 B.n301 VSUBS 0.009744f
C339 B.n302 VSUBS 0.009744f
C340 B.n303 VSUBS 0.009744f
C341 B.n304 VSUBS 0.009744f
C342 B.n305 VSUBS 0.009744f
C343 B.n306 VSUBS 0.009744f
C344 B.n307 VSUBS 0.009744f
C345 B.n308 VSUBS 0.009744f
C346 B.n309 VSUBS 0.009744f
C347 B.n310 VSUBS 0.009744f
C348 B.n311 VSUBS 0.009744f
C349 B.n312 VSUBS 0.009744f
C350 B.n313 VSUBS 0.009744f
C351 B.n314 VSUBS 0.009744f
C352 B.n315 VSUBS 0.009744f
C353 B.n316 VSUBS 0.009744f
C354 B.n317 VSUBS 0.009744f
C355 B.n318 VSUBS 0.009744f
C356 B.n319 VSUBS 0.009744f
C357 B.n320 VSUBS 0.009744f
C358 B.n321 VSUBS 0.009744f
C359 B.n322 VSUBS 0.009744f
C360 B.n323 VSUBS 0.009744f
C361 B.n324 VSUBS 0.009744f
C362 B.n325 VSUBS 0.009744f
C363 B.n326 VSUBS 0.009744f
C364 B.n327 VSUBS 0.009744f
C365 B.n328 VSUBS 0.022939f
C366 B.n329 VSUBS 0.024348f
C367 B.n330 VSUBS 0.024348f
C368 B.n331 VSUBS 0.009744f
C369 B.n332 VSUBS 0.009744f
C370 B.n333 VSUBS 0.009744f
C371 B.n334 VSUBS 0.009744f
C372 B.n335 VSUBS 0.009744f
C373 B.n336 VSUBS 0.009744f
C374 B.n337 VSUBS 0.009744f
C375 B.n338 VSUBS 0.009744f
C376 B.n339 VSUBS 0.009744f
C377 B.n340 VSUBS 0.009744f
C378 B.n341 VSUBS 0.009744f
C379 B.n342 VSUBS 0.009744f
C380 B.n343 VSUBS 0.009744f
C381 B.n344 VSUBS 0.009744f
C382 B.n345 VSUBS 0.009744f
C383 B.n346 VSUBS 0.009744f
C384 B.n347 VSUBS 0.009744f
C385 B.n348 VSUBS 0.009744f
C386 B.n349 VSUBS 0.009744f
C387 B.n350 VSUBS 0.009744f
C388 B.n351 VSUBS 0.009744f
C389 B.n352 VSUBS 0.009744f
C390 B.n353 VSUBS 0.009744f
C391 B.n354 VSUBS 0.009744f
C392 B.n355 VSUBS 0.009744f
C393 B.n356 VSUBS 0.009744f
C394 B.n357 VSUBS 0.009744f
C395 B.n358 VSUBS 0.009744f
C396 B.n359 VSUBS 0.009744f
C397 B.n360 VSUBS 0.009744f
C398 B.n361 VSUBS 0.009744f
C399 B.n362 VSUBS 0.009744f
C400 B.n363 VSUBS 0.009744f
C401 B.n364 VSUBS 0.009744f
C402 B.n365 VSUBS 0.009744f
C403 B.n366 VSUBS 0.009744f
C404 B.n367 VSUBS 0.009744f
C405 B.n368 VSUBS 0.009744f
C406 B.n369 VSUBS 0.009744f
C407 B.n370 VSUBS 0.009744f
C408 B.n371 VSUBS 0.009744f
C409 B.n372 VSUBS 0.009744f
C410 B.n373 VSUBS 0.009744f
C411 B.n374 VSUBS 0.009744f
C412 B.n375 VSUBS 0.009744f
C413 B.n376 VSUBS 0.009744f
C414 B.n377 VSUBS 0.009744f
C415 B.n378 VSUBS 0.009744f
C416 B.n379 VSUBS 0.009744f
C417 B.n380 VSUBS 0.009744f
C418 B.n381 VSUBS 0.009171f
C419 B.n382 VSUBS 0.022576f
C420 B.n383 VSUBS 0.005445f
C421 B.n384 VSUBS 0.009744f
C422 B.n385 VSUBS 0.009744f
C423 B.n386 VSUBS 0.009744f
C424 B.n387 VSUBS 0.009744f
C425 B.n388 VSUBS 0.009744f
C426 B.n389 VSUBS 0.009744f
C427 B.n390 VSUBS 0.009744f
C428 B.n391 VSUBS 0.009744f
C429 B.n392 VSUBS 0.009744f
C430 B.n393 VSUBS 0.009744f
C431 B.n394 VSUBS 0.009744f
C432 B.n395 VSUBS 0.009744f
C433 B.t2 VSUBS 0.434853f
C434 B.t1 VSUBS 0.468112f
C435 B.t0 VSUBS 2.01461f
C436 B.n396 VSUBS 0.258121f
C437 B.n397 VSUBS 0.10296f
C438 B.n398 VSUBS 0.022576f
C439 B.n399 VSUBS 0.005445f
C440 B.n400 VSUBS 0.009744f
C441 B.n401 VSUBS 0.009744f
C442 B.n402 VSUBS 0.009744f
C443 B.n403 VSUBS 0.009744f
C444 B.n404 VSUBS 0.009744f
C445 B.n405 VSUBS 0.009744f
C446 B.n406 VSUBS 0.009744f
C447 B.n407 VSUBS 0.009744f
C448 B.n408 VSUBS 0.009744f
C449 B.n409 VSUBS 0.009744f
C450 B.n410 VSUBS 0.009744f
C451 B.n411 VSUBS 0.009744f
C452 B.n412 VSUBS 0.009744f
C453 B.n413 VSUBS 0.009744f
C454 B.n414 VSUBS 0.009744f
C455 B.n415 VSUBS 0.009744f
C456 B.n416 VSUBS 0.009744f
C457 B.n417 VSUBS 0.009744f
C458 B.n418 VSUBS 0.009744f
C459 B.n419 VSUBS 0.009744f
C460 B.n420 VSUBS 0.009744f
C461 B.n421 VSUBS 0.009744f
C462 B.n422 VSUBS 0.009744f
C463 B.n423 VSUBS 0.009744f
C464 B.n424 VSUBS 0.009744f
C465 B.n425 VSUBS 0.009744f
C466 B.n426 VSUBS 0.009744f
C467 B.n427 VSUBS 0.009744f
C468 B.n428 VSUBS 0.009744f
C469 B.n429 VSUBS 0.009744f
C470 B.n430 VSUBS 0.009744f
C471 B.n431 VSUBS 0.009744f
C472 B.n432 VSUBS 0.009744f
C473 B.n433 VSUBS 0.009744f
C474 B.n434 VSUBS 0.009744f
C475 B.n435 VSUBS 0.009744f
C476 B.n436 VSUBS 0.009744f
C477 B.n437 VSUBS 0.009744f
C478 B.n438 VSUBS 0.009744f
C479 B.n439 VSUBS 0.009744f
C480 B.n440 VSUBS 0.009744f
C481 B.n441 VSUBS 0.009744f
C482 B.n442 VSUBS 0.009744f
C483 B.n443 VSUBS 0.009744f
C484 B.n444 VSUBS 0.009744f
C485 B.n445 VSUBS 0.009744f
C486 B.n446 VSUBS 0.009744f
C487 B.n447 VSUBS 0.009744f
C488 B.n448 VSUBS 0.009744f
C489 B.n449 VSUBS 0.009744f
C490 B.n450 VSUBS 0.009744f
C491 B.n451 VSUBS 0.009744f
C492 B.n452 VSUBS 0.023258f
C493 B.n453 VSUBS 0.024029f
C494 B.n454 VSUBS 0.022939f
C495 B.n455 VSUBS 0.009744f
C496 B.n456 VSUBS 0.009744f
C497 B.n457 VSUBS 0.009744f
C498 B.n458 VSUBS 0.009744f
C499 B.n459 VSUBS 0.009744f
C500 B.n460 VSUBS 0.009744f
C501 B.n461 VSUBS 0.009744f
C502 B.n462 VSUBS 0.009744f
C503 B.n463 VSUBS 0.009744f
C504 B.n464 VSUBS 0.009744f
C505 B.n465 VSUBS 0.009744f
C506 B.n466 VSUBS 0.009744f
C507 B.n467 VSUBS 0.009744f
C508 B.n468 VSUBS 0.009744f
C509 B.n469 VSUBS 0.009744f
C510 B.n470 VSUBS 0.009744f
C511 B.n471 VSUBS 0.009744f
C512 B.n472 VSUBS 0.009744f
C513 B.n473 VSUBS 0.009744f
C514 B.n474 VSUBS 0.009744f
C515 B.n475 VSUBS 0.009744f
C516 B.n476 VSUBS 0.009744f
C517 B.n477 VSUBS 0.009744f
C518 B.n478 VSUBS 0.009744f
C519 B.n479 VSUBS 0.009744f
C520 B.n480 VSUBS 0.009744f
C521 B.n481 VSUBS 0.009744f
C522 B.n482 VSUBS 0.009744f
C523 B.n483 VSUBS 0.009744f
C524 B.n484 VSUBS 0.009744f
C525 B.n485 VSUBS 0.009744f
C526 B.n486 VSUBS 0.009744f
C527 B.n487 VSUBS 0.009744f
C528 B.n488 VSUBS 0.009744f
C529 B.n489 VSUBS 0.009744f
C530 B.n490 VSUBS 0.009744f
C531 B.n491 VSUBS 0.009744f
C532 B.n492 VSUBS 0.009744f
C533 B.n493 VSUBS 0.009744f
C534 B.n494 VSUBS 0.009744f
C535 B.n495 VSUBS 0.009744f
C536 B.n496 VSUBS 0.009744f
C537 B.n497 VSUBS 0.009744f
C538 B.n498 VSUBS 0.009744f
C539 B.n499 VSUBS 0.009744f
C540 B.n500 VSUBS 0.009744f
C541 B.n501 VSUBS 0.009744f
C542 B.n502 VSUBS 0.009744f
C543 B.n503 VSUBS 0.009744f
C544 B.n504 VSUBS 0.009744f
C545 B.n505 VSUBS 0.009744f
C546 B.n506 VSUBS 0.009744f
C547 B.n507 VSUBS 0.009744f
C548 B.n508 VSUBS 0.009744f
C549 B.n509 VSUBS 0.009744f
C550 B.n510 VSUBS 0.009744f
C551 B.n511 VSUBS 0.009744f
C552 B.n512 VSUBS 0.009744f
C553 B.n513 VSUBS 0.009744f
C554 B.n514 VSUBS 0.009744f
C555 B.n515 VSUBS 0.009744f
C556 B.n516 VSUBS 0.009744f
C557 B.n517 VSUBS 0.009744f
C558 B.n518 VSUBS 0.009744f
C559 B.n519 VSUBS 0.009744f
C560 B.n520 VSUBS 0.009744f
C561 B.n521 VSUBS 0.009744f
C562 B.n522 VSUBS 0.009744f
C563 B.n523 VSUBS 0.009744f
C564 B.n524 VSUBS 0.009744f
C565 B.n525 VSUBS 0.009744f
C566 B.n526 VSUBS 0.009744f
C567 B.n527 VSUBS 0.009744f
C568 B.n528 VSUBS 0.009744f
C569 B.n529 VSUBS 0.009744f
C570 B.n530 VSUBS 0.009744f
C571 B.n531 VSUBS 0.009744f
C572 B.n532 VSUBS 0.009744f
C573 B.n533 VSUBS 0.009744f
C574 B.n534 VSUBS 0.009744f
C575 B.n535 VSUBS 0.009744f
C576 B.n536 VSUBS 0.009744f
C577 B.n537 VSUBS 0.009744f
C578 B.n538 VSUBS 0.009744f
C579 B.n539 VSUBS 0.009744f
C580 B.n540 VSUBS 0.009744f
C581 B.n541 VSUBS 0.009744f
C582 B.n542 VSUBS 0.009744f
C583 B.n543 VSUBS 0.009744f
C584 B.n544 VSUBS 0.009744f
C585 B.n545 VSUBS 0.009744f
C586 B.n546 VSUBS 0.009744f
C587 B.n547 VSUBS 0.009744f
C588 B.n548 VSUBS 0.009744f
C589 B.n549 VSUBS 0.009744f
C590 B.n550 VSUBS 0.009744f
C591 B.n551 VSUBS 0.009744f
C592 B.n552 VSUBS 0.009744f
C593 B.n553 VSUBS 0.009744f
C594 B.n554 VSUBS 0.009744f
C595 B.n555 VSUBS 0.009744f
C596 B.n556 VSUBS 0.009744f
C597 B.n557 VSUBS 0.009744f
C598 B.n558 VSUBS 0.009744f
C599 B.n559 VSUBS 0.009744f
C600 B.n560 VSUBS 0.009744f
C601 B.n561 VSUBS 0.009744f
C602 B.n562 VSUBS 0.009744f
C603 B.n563 VSUBS 0.009744f
C604 B.n564 VSUBS 0.009744f
C605 B.n565 VSUBS 0.009744f
C606 B.n566 VSUBS 0.009744f
C607 B.n567 VSUBS 0.009744f
C608 B.n568 VSUBS 0.009744f
C609 B.n569 VSUBS 0.009744f
C610 B.n570 VSUBS 0.009744f
C611 B.n571 VSUBS 0.009744f
C612 B.n572 VSUBS 0.009744f
C613 B.n573 VSUBS 0.009744f
C614 B.n574 VSUBS 0.009744f
C615 B.n575 VSUBS 0.009744f
C616 B.n576 VSUBS 0.009744f
C617 B.n577 VSUBS 0.009744f
C618 B.n578 VSUBS 0.009744f
C619 B.n579 VSUBS 0.009744f
C620 B.n580 VSUBS 0.009744f
C621 B.n581 VSUBS 0.009744f
C622 B.n582 VSUBS 0.009744f
C623 B.n583 VSUBS 0.009744f
C624 B.n584 VSUBS 0.009744f
C625 B.n585 VSUBS 0.009744f
C626 B.n586 VSUBS 0.009744f
C627 B.n587 VSUBS 0.009744f
C628 B.n588 VSUBS 0.009744f
C629 B.n589 VSUBS 0.009744f
C630 B.n590 VSUBS 0.009744f
C631 B.n591 VSUBS 0.009744f
C632 B.n592 VSUBS 0.009744f
C633 B.n593 VSUBS 0.009744f
C634 B.n594 VSUBS 0.009744f
C635 B.n595 VSUBS 0.009744f
C636 B.n596 VSUBS 0.009744f
C637 B.n597 VSUBS 0.009744f
C638 B.n598 VSUBS 0.009744f
C639 B.n599 VSUBS 0.009744f
C640 B.n600 VSUBS 0.009744f
C641 B.n601 VSUBS 0.009744f
C642 B.n602 VSUBS 0.009744f
C643 B.n603 VSUBS 0.009744f
C644 B.n604 VSUBS 0.009744f
C645 B.n605 VSUBS 0.009744f
C646 B.n606 VSUBS 0.009744f
C647 B.n607 VSUBS 0.009744f
C648 B.n608 VSUBS 0.009744f
C649 B.n609 VSUBS 0.009744f
C650 B.n610 VSUBS 0.009744f
C651 B.n611 VSUBS 0.009744f
C652 B.n612 VSUBS 0.009744f
C653 B.n613 VSUBS 0.009744f
C654 B.n614 VSUBS 0.009744f
C655 B.n615 VSUBS 0.009744f
C656 B.n616 VSUBS 0.009744f
C657 B.n617 VSUBS 0.009744f
C658 B.n618 VSUBS 0.009744f
C659 B.n619 VSUBS 0.009744f
C660 B.n620 VSUBS 0.009744f
C661 B.n621 VSUBS 0.009744f
C662 B.n622 VSUBS 0.009744f
C663 B.n623 VSUBS 0.009744f
C664 B.n624 VSUBS 0.009744f
C665 B.n625 VSUBS 0.009744f
C666 B.n626 VSUBS 0.009744f
C667 B.n627 VSUBS 0.009744f
C668 B.n628 VSUBS 0.009744f
C669 B.n629 VSUBS 0.009744f
C670 B.n630 VSUBS 0.009744f
C671 B.n631 VSUBS 0.009744f
C672 B.n632 VSUBS 0.009744f
C673 B.n633 VSUBS 0.009744f
C674 B.n634 VSUBS 0.009744f
C675 B.n635 VSUBS 0.009744f
C676 B.n636 VSUBS 0.009744f
C677 B.n637 VSUBS 0.009744f
C678 B.n638 VSUBS 0.009744f
C679 B.n639 VSUBS 0.009744f
C680 B.n640 VSUBS 0.009744f
C681 B.n641 VSUBS 0.009744f
C682 B.n642 VSUBS 0.009744f
C683 B.n643 VSUBS 0.009744f
C684 B.n644 VSUBS 0.009744f
C685 B.n645 VSUBS 0.009744f
C686 B.n646 VSUBS 0.009744f
C687 B.n647 VSUBS 0.009744f
C688 B.n648 VSUBS 0.009744f
C689 B.n649 VSUBS 0.009744f
C690 B.n650 VSUBS 0.009744f
C691 B.n651 VSUBS 0.009744f
C692 B.n652 VSUBS 0.009744f
C693 B.n653 VSUBS 0.009744f
C694 B.n654 VSUBS 0.009744f
C695 B.n655 VSUBS 0.009744f
C696 B.n656 VSUBS 0.009744f
C697 B.n657 VSUBS 0.009744f
C698 B.n658 VSUBS 0.009744f
C699 B.n659 VSUBS 0.009744f
C700 B.n660 VSUBS 0.009744f
C701 B.n661 VSUBS 0.009744f
C702 B.n662 VSUBS 0.022939f
C703 B.n663 VSUBS 0.024348f
C704 B.n664 VSUBS 0.024348f
C705 B.n665 VSUBS 0.009744f
C706 B.n666 VSUBS 0.009744f
C707 B.n667 VSUBS 0.009744f
C708 B.n668 VSUBS 0.009744f
C709 B.n669 VSUBS 0.009744f
C710 B.n670 VSUBS 0.009744f
C711 B.n671 VSUBS 0.009744f
C712 B.n672 VSUBS 0.009744f
C713 B.n673 VSUBS 0.009744f
C714 B.n674 VSUBS 0.009744f
C715 B.n675 VSUBS 0.009744f
C716 B.n676 VSUBS 0.009744f
C717 B.n677 VSUBS 0.009744f
C718 B.n678 VSUBS 0.009744f
C719 B.n679 VSUBS 0.009744f
C720 B.n680 VSUBS 0.009744f
C721 B.n681 VSUBS 0.009744f
C722 B.n682 VSUBS 0.009744f
C723 B.n683 VSUBS 0.009744f
C724 B.n684 VSUBS 0.009744f
C725 B.n685 VSUBS 0.009744f
C726 B.n686 VSUBS 0.009744f
C727 B.n687 VSUBS 0.009744f
C728 B.n688 VSUBS 0.009744f
C729 B.n689 VSUBS 0.009744f
C730 B.n690 VSUBS 0.009744f
C731 B.n691 VSUBS 0.009744f
C732 B.n692 VSUBS 0.009744f
C733 B.n693 VSUBS 0.009744f
C734 B.n694 VSUBS 0.009744f
C735 B.n695 VSUBS 0.009744f
C736 B.n696 VSUBS 0.009744f
C737 B.n697 VSUBS 0.009744f
C738 B.n698 VSUBS 0.009744f
C739 B.n699 VSUBS 0.009744f
C740 B.n700 VSUBS 0.009744f
C741 B.n701 VSUBS 0.009744f
C742 B.n702 VSUBS 0.009744f
C743 B.n703 VSUBS 0.009744f
C744 B.n704 VSUBS 0.009744f
C745 B.n705 VSUBS 0.009744f
C746 B.n706 VSUBS 0.009744f
C747 B.n707 VSUBS 0.009744f
C748 B.n708 VSUBS 0.009744f
C749 B.n709 VSUBS 0.009744f
C750 B.n710 VSUBS 0.009744f
C751 B.n711 VSUBS 0.009744f
C752 B.n712 VSUBS 0.009744f
C753 B.n713 VSUBS 0.009744f
C754 B.n714 VSUBS 0.009744f
C755 B.n715 VSUBS 0.009171f
C756 B.n716 VSUBS 0.022576f
C757 B.n717 VSUBS 0.005445f
C758 B.n718 VSUBS 0.009744f
C759 B.n719 VSUBS 0.009744f
C760 B.n720 VSUBS 0.009744f
C761 B.n721 VSUBS 0.009744f
C762 B.n722 VSUBS 0.009744f
C763 B.n723 VSUBS 0.009744f
C764 B.n724 VSUBS 0.009744f
C765 B.n725 VSUBS 0.009744f
C766 B.n726 VSUBS 0.009744f
C767 B.n727 VSUBS 0.009744f
C768 B.n728 VSUBS 0.009744f
C769 B.n729 VSUBS 0.009744f
C770 B.n730 VSUBS 0.005445f
C771 B.n731 VSUBS 0.009744f
C772 B.n732 VSUBS 0.009744f
C773 B.n733 VSUBS 0.009171f
C774 B.n734 VSUBS 0.009744f
C775 B.n735 VSUBS 0.009744f
C776 B.n736 VSUBS 0.009744f
C777 B.n737 VSUBS 0.009744f
C778 B.n738 VSUBS 0.009744f
C779 B.n739 VSUBS 0.009744f
C780 B.n740 VSUBS 0.009744f
C781 B.n741 VSUBS 0.009744f
C782 B.n742 VSUBS 0.009744f
C783 B.n743 VSUBS 0.009744f
C784 B.n744 VSUBS 0.009744f
C785 B.n745 VSUBS 0.009744f
C786 B.n746 VSUBS 0.009744f
C787 B.n747 VSUBS 0.009744f
C788 B.n748 VSUBS 0.009744f
C789 B.n749 VSUBS 0.009744f
C790 B.n750 VSUBS 0.009744f
C791 B.n751 VSUBS 0.009744f
C792 B.n752 VSUBS 0.009744f
C793 B.n753 VSUBS 0.009744f
C794 B.n754 VSUBS 0.009744f
C795 B.n755 VSUBS 0.009744f
C796 B.n756 VSUBS 0.009744f
C797 B.n757 VSUBS 0.009744f
C798 B.n758 VSUBS 0.009744f
C799 B.n759 VSUBS 0.009744f
C800 B.n760 VSUBS 0.009744f
C801 B.n761 VSUBS 0.009744f
C802 B.n762 VSUBS 0.009744f
C803 B.n763 VSUBS 0.009744f
C804 B.n764 VSUBS 0.009744f
C805 B.n765 VSUBS 0.009744f
C806 B.n766 VSUBS 0.009744f
C807 B.n767 VSUBS 0.009744f
C808 B.n768 VSUBS 0.009744f
C809 B.n769 VSUBS 0.009744f
C810 B.n770 VSUBS 0.009744f
C811 B.n771 VSUBS 0.009744f
C812 B.n772 VSUBS 0.009744f
C813 B.n773 VSUBS 0.009744f
C814 B.n774 VSUBS 0.009744f
C815 B.n775 VSUBS 0.009744f
C816 B.n776 VSUBS 0.009744f
C817 B.n777 VSUBS 0.009744f
C818 B.n778 VSUBS 0.009744f
C819 B.n779 VSUBS 0.009744f
C820 B.n780 VSUBS 0.009744f
C821 B.n781 VSUBS 0.009744f
C822 B.n782 VSUBS 0.009744f
C823 B.n783 VSUBS 0.024348f
C824 B.n784 VSUBS 0.024348f
C825 B.n785 VSUBS 0.022939f
C826 B.n786 VSUBS 0.009744f
C827 B.n787 VSUBS 0.009744f
C828 B.n788 VSUBS 0.009744f
C829 B.n789 VSUBS 0.009744f
C830 B.n790 VSUBS 0.009744f
C831 B.n791 VSUBS 0.009744f
C832 B.n792 VSUBS 0.009744f
C833 B.n793 VSUBS 0.009744f
C834 B.n794 VSUBS 0.009744f
C835 B.n795 VSUBS 0.009744f
C836 B.n796 VSUBS 0.009744f
C837 B.n797 VSUBS 0.009744f
C838 B.n798 VSUBS 0.009744f
C839 B.n799 VSUBS 0.009744f
C840 B.n800 VSUBS 0.009744f
C841 B.n801 VSUBS 0.009744f
C842 B.n802 VSUBS 0.009744f
C843 B.n803 VSUBS 0.009744f
C844 B.n804 VSUBS 0.009744f
C845 B.n805 VSUBS 0.009744f
C846 B.n806 VSUBS 0.009744f
C847 B.n807 VSUBS 0.009744f
C848 B.n808 VSUBS 0.009744f
C849 B.n809 VSUBS 0.009744f
C850 B.n810 VSUBS 0.009744f
C851 B.n811 VSUBS 0.009744f
C852 B.n812 VSUBS 0.009744f
C853 B.n813 VSUBS 0.009744f
C854 B.n814 VSUBS 0.009744f
C855 B.n815 VSUBS 0.009744f
C856 B.n816 VSUBS 0.009744f
C857 B.n817 VSUBS 0.009744f
C858 B.n818 VSUBS 0.009744f
C859 B.n819 VSUBS 0.009744f
C860 B.n820 VSUBS 0.009744f
C861 B.n821 VSUBS 0.009744f
C862 B.n822 VSUBS 0.009744f
C863 B.n823 VSUBS 0.009744f
C864 B.n824 VSUBS 0.009744f
C865 B.n825 VSUBS 0.009744f
C866 B.n826 VSUBS 0.009744f
C867 B.n827 VSUBS 0.009744f
C868 B.n828 VSUBS 0.009744f
C869 B.n829 VSUBS 0.009744f
C870 B.n830 VSUBS 0.009744f
C871 B.n831 VSUBS 0.009744f
C872 B.n832 VSUBS 0.009744f
C873 B.n833 VSUBS 0.009744f
C874 B.n834 VSUBS 0.009744f
C875 B.n835 VSUBS 0.009744f
C876 B.n836 VSUBS 0.009744f
C877 B.n837 VSUBS 0.009744f
C878 B.n838 VSUBS 0.009744f
C879 B.n839 VSUBS 0.009744f
C880 B.n840 VSUBS 0.009744f
C881 B.n841 VSUBS 0.009744f
C882 B.n842 VSUBS 0.009744f
C883 B.n843 VSUBS 0.009744f
C884 B.n844 VSUBS 0.009744f
C885 B.n845 VSUBS 0.009744f
C886 B.n846 VSUBS 0.009744f
C887 B.n847 VSUBS 0.009744f
C888 B.n848 VSUBS 0.009744f
C889 B.n849 VSUBS 0.009744f
C890 B.n850 VSUBS 0.009744f
C891 B.n851 VSUBS 0.009744f
C892 B.n852 VSUBS 0.009744f
C893 B.n853 VSUBS 0.009744f
C894 B.n854 VSUBS 0.009744f
C895 B.n855 VSUBS 0.009744f
C896 B.n856 VSUBS 0.009744f
C897 B.n857 VSUBS 0.009744f
C898 B.n858 VSUBS 0.009744f
C899 B.n859 VSUBS 0.009744f
C900 B.n860 VSUBS 0.009744f
C901 B.n861 VSUBS 0.009744f
C902 B.n862 VSUBS 0.009744f
C903 B.n863 VSUBS 0.009744f
C904 B.n864 VSUBS 0.009744f
C905 B.n865 VSUBS 0.009744f
C906 B.n866 VSUBS 0.009744f
C907 B.n867 VSUBS 0.009744f
C908 B.n868 VSUBS 0.009744f
C909 B.n869 VSUBS 0.009744f
C910 B.n870 VSUBS 0.009744f
C911 B.n871 VSUBS 0.009744f
C912 B.n872 VSUBS 0.009744f
C913 B.n873 VSUBS 0.009744f
C914 B.n874 VSUBS 0.009744f
C915 B.n875 VSUBS 0.009744f
C916 B.n876 VSUBS 0.009744f
C917 B.n877 VSUBS 0.009744f
C918 B.n878 VSUBS 0.009744f
C919 B.n879 VSUBS 0.009744f
C920 B.n880 VSUBS 0.009744f
C921 B.n881 VSUBS 0.009744f
C922 B.n882 VSUBS 0.009744f
C923 B.n883 VSUBS 0.009744f
C924 B.n884 VSUBS 0.009744f
C925 B.n885 VSUBS 0.009744f
C926 B.n886 VSUBS 0.009744f
C927 B.n887 VSUBS 0.012715f
C928 B.n888 VSUBS 0.013545f
C929 B.n889 VSUBS 0.026936f
C930 VDD1.t9 VSUBS 2.46871f
C931 VDD1.t7 VSUBS 0.244853f
C932 VDD1.t0 VSUBS 0.244853f
C933 VDD1.n0 VSUBS 1.8566f
C934 VDD1.n1 VSUBS 1.86953f
C935 VDD1.t6 VSUBS 2.4687f
C936 VDD1.t5 VSUBS 0.244853f
C937 VDD1.t2 VSUBS 0.244853f
C938 VDD1.n2 VSUBS 1.8566f
C939 VDD1.n3 VSUBS 1.85905f
C940 VDD1.t3 VSUBS 0.244853f
C941 VDD1.t1 VSUBS 0.244853f
C942 VDD1.n4 VSUBS 1.88522f
C943 VDD1.n5 VSUBS 4.33247f
C944 VDD1.t8 VSUBS 0.244853f
C945 VDD1.t4 VSUBS 0.244853f
C946 VDD1.n6 VSUBS 1.85659f
C947 VDD1.n7 VSUBS 4.3818f
C948 VP.t8 VSUBS 2.50164f
C949 VP.n0 VSUBS 0.998069f
C950 VP.n1 VSUBS 0.029777f
C951 VP.n2 VSUBS 0.024183f
C952 VP.n3 VSUBS 0.029777f
C953 VP.t6 VSUBS 2.50164f
C954 VP.n4 VSUBS 0.890717f
C955 VP.n5 VSUBS 0.029777f
C956 VP.n6 VSUBS 0.024106f
C957 VP.n7 VSUBS 0.029777f
C958 VP.t7 VSUBS 2.50164f
C959 VP.n8 VSUBS 0.890717f
C960 VP.n9 VSUBS 0.029777f
C961 VP.n10 VSUBS 0.024106f
C962 VP.n11 VSUBS 0.029777f
C963 VP.t4 VSUBS 2.50164f
C964 VP.n12 VSUBS 0.890717f
C965 VP.n13 VSUBS 0.029777f
C966 VP.n14 VSUBS 0.024183f
C967 VP.n15 VSUBS 0.029777f
C968 VP.t3 VSUBS 2.50164f
C969 VP.n16 VSUBS 0.998069f
C970 VP.t5 VSUBS 2.50164f
C971 VP.n17 VSUBS 0.998069f
C972 VP.n18 VSUBS 0.029777f
C973 VP.n19 VSUBS 0.024183f
C974 VP.n20 VSUBS 0.029777f
C975 VP.t1 VSUBS 2.50164f
C976 VP.n21 VSUBS 0.890717f
C977 VP.n22 VSUBS 0.029777f
C978 VP.n23 VSUBS 0.024106f
C979 VP.n24 VSUBS 0.029777f
C980 VP.t9 VSUBS 2.50164f
C981 VP.n25 VSUBS 0.890717f
C982 VP.n26 VSUBS 0.029777f
C983 VP.n27 VSUBS 0.024106f
C984 VP.n28 VSUBS 0.029777f
C985 VP.t2 VSUBS 2.50164f
C986 VP.n29 VSUBS 0.988283f
C987 VP.t0 VSUBS 2.83266f
C988 VP.n30 VSUBS 0.944935f
C989 VP.n31 VSUBS 0.346313f
C990 VP.n32 VSUBS 0.041455f
C991 VP.n33 VSUBS 0.055775f
C992 VP.n34 VSUBS 0.059644f
C993 VP.n35 VSUBS 0.029777f
C994 VP.n36 VSUBS 0.029777f
C995 VP.n37 VSUBS 0.029777f
C996 VP.n38 VSUBS 0.059342f
C997 VP.n39 VSUBS 0.055775f
C998 VP.n40 VSUBS 0.042006f
C999 VP.n41 VSUBS 0.029777f
C1000 VP.n42 VSUBS 0.029777f
C1001 VP.n43 VSUBS 0.042006f
C1002 VP.n44 VSUBS 0.055775f
C1003 VP.n45 VSUBS 0.059342f
C1004 VP.n46 VSUBS 0.029777f
C1005 VP.n47 VSUBS 0.029777f
C1006 VP.n48 VSUBS 0.029777f
C1007 VP.n49 VSUBS 0.059644f
C1008 VP.n50 VSUBS 0.055775f
C1009 VP.n51 VSUBS 0.041455f
C1010 VP.n52 VSUBS 0.029777f
C1011 VP.n53 VSUBS 0.029777f
C1012 VP.n54 VSUBS 0.042557f
C1013 VP.n55 VSUBS 0.055775f
C1014 VP.n56 VSUBS 0.059003f
C1015 VP.n57 VSUBS 0.029777f
C1016 VP.n58 VSUBS 0.029777f
C1017 VP.n59 VSUBS 0.029777f
C1018 VP.n60 VSUBS 0.059906f
C1019 VP.n61 VSUBS 0.055775f
C1020 VP.n62 VSUBS 0.040904f
C1021 VP.n63 VSUBS 0.048067f
C1022 VP.n64 VSUBS 1.91383f
C1023 VP.n65 VSUBS 1.93341f
C1024 VP.n66 VSUBS 0.048067f
C1025 VP.n67 VSUBS 0.040904f
C1026 VP.n68 VSUBS 0.055775f
C1027 VP.n69 VSUBS 0.059906f
C1028 VP.n70 VSUBS 0.029777f
C1029 VP.n71 VSUBS 0.029777f
C1030 VP.n72 VSUBS 0.029777f
C1031 VP.n73 VSUBS 0.059003f
C1032 VP.n74 VSUBS 0.055775f
C1033 VP.n75 VSUBS 0.042557f
C1034 VP.n76 VSUBS 0.029777f
C1035 VP.n77 VSUBS 0.029777f
C1036 VP.n78 VSUBS 0.041455f
C1037 VP.n79 VSUBS 0.055775f
C1038 VP.n80 VSUBS 0.059644f
C1039 VP.n81 VSUBS 0.029777f
C1040 VP.n82 VSUBS 0.029777f
C1041 VP.n83 VSUBS 0.029777f
C1042 VP.n84 VSUBS 0.059342f
C1043 VP.n85 VSUBS 0.055775f
C1044 VP.n86 VSUBS 0.042006f
C1045 VP.n87 VSUBS 0.029777f
C1046 VP.n88 VSUBS 0.029777f
C1047 VP.n89 VSUBS 0.042006f
C1048 VP.n90 VSUBS 0.055775f
C1049 VP.n91 VSUBS 0.059342f
C1050 VP.n92 VSUBS 0.029777f
C1051 VP.n93 VSUBS 0.029777f
C1052 VP.n94 VSUBS 0.029777f
C1053 VP.n95 VSUBS 0.059644f
C1054 VP.n96 VSUBS 0.055775f
C1055 VP.n97 VSUBS 0.041455f
C1056 VP.n98 VSUBS 0.029777f
C1057 VP.n99 VSUBS 0.029777f
C1058 VP.n100 VSUBS 0.042557f
C1059 VP.n101 VSUBS 0.055775f
C1060 VP.n102 VSUBS 0.059003f
C1061 VP.n103 VSUBS 0.029777f
C1062 VP.n104 VSUBS 0.029777f
C1063 VP.n105 VSUBS 0.029777f
C1064 VP.n106 VSUBS 0.059906f
C1065 VP.n107 VSUBS 0.055775f
C1066 VP.n108 VSUBS 0.040904f
C1067 VP.n109 VSUBS 0.048067f
C1068 VP.n110 VSUBS 0.07405f
C1069 VDD2.t6 VSUBS 2.47936f
C1070 VDD2.t8 VSUBS 0.24591f
C1071 VDD2.t5 VSUBS 0.24591f
C1072 VDD2.n0 VSUBS 1.86462f
C1073 VDD2.n1 VSUBS 1.86708f
C1074 VDD2.t7 VSUBS 0.24591f
C1075 VDD2.t9 VSUBS 0.24591f
C1076 VDD2.n2 VSUBS 1.89337f
C1077 VDD2.n3 VSUBS 4.1755f
C1078 VDD2.t3 VSUBS 2.44655f
C1079 VDD2.n4 VSUBS 4.32362f
C1080 VDD2.t1 VSUBS 0.24591f
C1081 VDD2.t2 VSUBS 0.24591f
C1082 VDD2.n5 VSUBS 1.86462f
C1083 VDD2.n6 VSUBS 0.945839f
C1084 VDD2.t0 VSUBS 0.24591f
C1085 VDD2.t4 VSUBS 0.24591f
C1086 VDD2.n7 VSUBS 1.89331f
C1087 VTAIL.t8 VSUBS 0.236201f
C1088 VTAIL.t11 VSUBS 0.236201f
C1089 VTAIL.n0 VSUBS 1.65632f
C1090 VTAIL.n1 VSUBS 1.04788f
C1091 VTAIL.t16 VSUBS 2.20106f
C1092 VTAIL.n2 VSUBS 1.21539f
C1093 VTAIL.t13 VSUBS 0.236201f
C1094 VTAIL.t12 VSUBS 0.236201f
C1095 VTAIL.n3 VSUBS 1.65632f
C1096 VTAIL.n4 VSUBS 1.21741f
C1097 VTAIL.t0 VSUBS 0.236201f
C1098 VTAIL.t1 VSUBS 0.236201f
C1099 VTAIL.n5 VSUBS 1.65632f
C1100 VTAIL.n6 VSUBS 2.75624f
C1101 VTAIL.t2 VSUBS 0.236201f
C1102 VTAIL.t6 VSUBS 0.236201f
C1103 VTAIL.n7 VSUBS 1.65633f
C1104 VTAIL.n8 VSUBS 2.75623f
C1105 VTAIL.t9 VSUBS 0.236201f
C1106 VTAIL.t5 VSUBS 0.236201f
C1107 VTAIL.n9 VSUBS 1.65633f
C1108 VTAIL.n10 VSUBS 1.2174f
C1109 VTAIL.t4 VSUBS 2.20108f
C1110 VTAIL.n11 VSUBS 1.21537f
C1111 VTAIL.t15 VSUBS 0.236201f
C1112 VTAIL.t18 VSUBS 0.236201f
C1113 VTAIL.n12 VSUBS 1.65633f
C1114 VTAIL.n13 VSUBS 1.11594f
C1115 VTAIL.t19 VSUBS 0.236201f
C1116 VTAIL.t14 VSUBS 0.236201f
C1117 VTAIL.n14 VSUBS 1.65633f
C1118 VTAIL.n15 VSUBS 1.2174f
C1119 VTAIL.t17 VSUBS 2.20106f
C1120 VTAIL.n16 VSUBS 2.56059f
C1121 VTAIL.t10 VSUBS 2.20106f
C1122 VTAIL.n17 VSUBS 2.5606f
C1123 VTAIL.t3 VSUBS 0.236201f
C1124 VTAIL.t7 VSUBS 0.236201f
C1125 VTAIL.n18 VSUBS 1.65632f
C1126 VTAIL.n19 VSUBS 0.990391f
C1127 VN.t0 VSUBS 2.28947f
C1128 VN.n0 VSUBS 0.913423f
C1129 VN.n1 VSUBS 0.027252f
C1130 VN.n2 VSUBS 0.022132f
C1131 VN.n3 VSUBS 0.027252f
C1132 VN.t2 VSUBS 2.28947f
C1133 VN.n4 VSUBS 0.815176f
C1134 VN.n5 VSUBS 0.027252f
C1135 VN.n6 VSUBS 0.022062f
C1136 VN.n7 VSUBS 0.027252f
C1137 VN.t4 VSUBS 2.28947f
C1138 VN.n8 VSUBS 0.815176f
C1139 VN.n9 VSUBS 0.027252f
C1140 VN.n10 VSUBS 0.022062f
C1141 VN.n11 VSUBS 0.027252f
C1142 VN.t1 VSUBS 2.28947f
C1143 VN.n12 VSUBS 0.904468f
C1144 VN.t3 VSUBS 2.59243f
C1145 VN.n13 VSUBS 0.864795f
C1146 VN.n14 VSUBS 0.316942f
C1147 VN.n15 VSUBS 0.03794f
C1148 VN.n16 VSUBS 0.051045f
C1149 VN.n17 VSUBS 0.054586f
C1150 VN.n18 VSUBS 0.027252f
C1151 VN.n19 VSUBS 0.027252f
C1152 VN.n20 VSUBS 0.027252f
C1153 VN.n21 VSUBS 0.054309f
C1154 VN.n22 VSUBS 0.051045f
C1155 VN.n23 VSUBS 0.038444f
C1156 VN.n24 VSUBS 0.027252f
C1157 VN.n25 VSUBS 0.027252f
C1158 VN.n26 VSUBS 0.038444f
C1159 VN.n27 VSUBS 0.051045f
C1160 VN.n28 VSUBS 0.054309f
C1161 VN.n29 VSUBS 0.027252f
C1162 VN.n30 VSUBS 0.027252f
C1163 VN.n31 VSUBS 0.027252f
C1164 VN.n32 VSUBS 0.054586f
C1165 VN.n33 VSUBS 0.051045f
C1166 VN.n34 VSUBS 0.03794f
C1167 VN.n35 VSUBS 0.027252f
C1168 VN.n36 VSUBS 0.027252f
C1169 VN.n37 VSUBS 0.038948f
C1170 VN.n38 VSUBS 0.051045f
C1171 VN.n39 VSUBS 0.053999f
C1172 VN.n40 VSUBS 0.027252f
C1173 VN.n41 VSUBS 0.027252f
C1174 VN.n42 VSUBS 0.027252f
C1175 VN.n43 VSUBS 0.054825f
C1176 VN.n44 VSUBS 0.051045f
C1177 VN.n45 VSUBS 0.037436f
C1178 VN.n46 VSUBS 0.043991f
C1179 VN.n47 VSUBS 0.067769f
C1180 VN.t6 VSUBS 2.28947f
C1181 VN.n48 VSUBS 0.913423f
C1182 VN.n49 VSUBS 0.027252f
C1183 VN.n50 VSUBS 0.022132f
C1184 VN.n51 VSUBS 0.027252f
C1185 VN.t8 VSUBS 2.28947f
C1186 VN.n52 VSUBS 0.815176f
C1187 VN.n53 VSUBS 0.027252f
C1188 VN.n54 VSUBS 0.022062f
C1189 VN.n55 VSUBS 0.027252f
C1190 VN.t7 VSUBS 2.28947f
C1191 VN.n56 VSUBS 0.815176f
C1192 VN.n57 VSUBS 0.027252f
C1193 VN.n58 VSUBS 0.022062f
C1194 VN.n59 VSUBS 0.027252f
C1195 VN.t9 VSUBS 2.28947f
C1196 VN.n60 VSUBS 0.904468f
C1197 VN.t5 VSUBS 2.59243f
C1198 VN.n61 VSUBS 0.864795f
C1199 VN.n62 VSUBS 0.316942f
C1200 VN.n63 VSUBS 0.03794f
C1201 VN.n64 VSUBS 0.051045f
C1202 VN.n65 VSUBS 0.054586f
C1203 VN.n66 VSUBS 0.027252f
C1204 VN.n67 VSUBS 0.027252f
C1205 VN.n68 VSUBS 0.027252f
C1206 VN.n69 VSUBS 0.054309f
C1207 VN.n70 VSUBS 0.051045f
C1208 VN.n71 VSUBS 0.038444f
C1209 VN.n72 VSUBS 0.027252f
C1210 VN.n73 VSUBS 0.027252f
C1211 VN.n74 VSUBS 0.038444f
C1212 VN.n75 VSUBS 0.051045f
C1213 VN.n76 VSUBS 0.054309f
C1214 VN.n77 VSUBS 0.027252f
C1215 VN.n78 VSUBS 0.027252f
C1216 VN.n79 VSUBS 0.027252f
C1217 VN.n80 VSUBS 0.054586f
C1218 VN.n81 VSUBS 0.051045f
C1219 VN.n82 VSUBS 0.03794f
C1220 VN.n83 VSUBS 0.027252f
C1221 VN.n84 VSUBS 0.027252f
C1222 VN.n85 VSUBS 0.038948f
C1223 VN.n86 VSUBS 0.051045f
C1224 VN.n87 VSUBS 0.053999f
C1225 VN.n88 VSUBS 0.027252f
C1226 VN.n89 VSUBS 0.027252f
C1227 VN.n90 VSUBS 0.027252f
C1228 VN.n91 VSUBS 0.054825f
C1229 VN.n92 VSUBS 0.051045f
C1230 VN.n93 VSUBS 0.037436f
C1231 VN.n94 VSUBS 0.043991f
C1232 VN.n95 VSUBS 1.76237f
.ends

