* NGSPICE file created from diff_pair_sample_0691.ext - technology: sky130A

.subckt diff_pair_sample_0691 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=1.78
X1 VTAIL.t6 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=1.78
X2 VTAIL.t7 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=1.78
X3 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=1.78
X4 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=1.78
X5 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=1.78
X6 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=1.78
X7 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=1.78
X8 VDD2.t0 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=1.78
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=1.78
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=1.78
X11 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=1.78
R0 VN.n0 VN.t2 105.374
R1 VN.n1 VN.t3 105.374
R2 VN.n0 VN.t0 104.945
R3 VN.n1 VN.t1 104.945
R4 VN VN.n1 48.1909
R5 VN VN.n0 9.34621
R6 VTAIL.n5 VTAIL.t3 60.2615
R7 VTAIL.n4 VTAIL.t4 60.2615
R8 VTAIL.n3 VTAIL.t6 60.2615
R9 VTAIL.n7 VTAIL.t5 60.2614
R10 VTAIL.n0 VTAIL.t7 60.2614
R11 VTAIL.n1 VTAIL.t1 60.2614
R12 VTAIL.n2 VTAIL.t0 60.2614
R13 VTAIL.n6 VTAIL.t2 60.2614
R14 VTAIL.n7 VTAIL.n6 18.5824
R15 VTAIL.n3 VTAIL.n2 18.5824
R16 VTAIL.n4 VTAIL.n3 1.81947
R17 VTAIL.n6 VTAIL.n5 1.81947
R18 VTAIL.n2 VTAIL.n1 1.81947
R19 VTAIL VTAIL.n0 0.968172
R20 VTAIL VTAIL.n7 0.851793
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 106.626
R24 VDD2.n2 VDD2.n1 73.0578
R25 VDD2.n1 VDD2.t2 3.88285
R26 VDD2.n1 VDD2.t0 3.88285
R27 VDD2.n0 VDD2.t1 3.88285
R28 VDD2.n0 VDD2.t3 3.88285
R29 VDD2 VDD2.n2 0.0586897
R30 B.n382 B.n381 585
R31 B.n384 B.n82 585
R32 B.n387 B.n386 585
R33 B.n388 B.n81 585
R34 B.n390 B.n389 585
R35 B.n392 B.n80 585
R36 B.n395 B.n394 585
R37 B.n396 B.n79 585
R38 B.n398 B.n397 585
R39 B.n400 B.n78 585
R40 B.n403 B.n402 585
R41 B.n404 B.n77 585
R42 B.n406 B.n405 585
R43 B.n408 B.n76 585
R44 B.n411 B.n410 585
R45 B.n412 B.n75 585
R46 B.n414 B.n413 585
R47 B.n416 B.n74 585
R48 B.n419 B.n418 585
R49 B.n420 B.n70 585
R50 B.n422 B.n421 585
R51 B.n424 B.n69 585
R52 B.n427 B.n426 585
R53 B.n428 B.n68 585
R54 B.n430 B.n429 585
R55 B.n432 B.n67 585
R56 B.n435 B.n434 585
R57 B.n436 B.n66 585
R58 B.n438 B.n437 585
R59 B.n440 B.n65 585
R60 B.n443 B.n442 585
R61 B.n445 B.n62 585
R62 B.n447 B.n446 585
R63 B.n449 B.n61 585
R64 B.n452 B.n451 585
R65 B.n453 B.n60 585
R66 B.n455 B.n454 585
R67 B.n457 B.n59 585
R68 B.n460 B.n459 585
R69 B.n461 B.n58 585
R70 B.n463 B.n462 585
R71 B.n465 B.n57 585
R72 B.n468 B.n467 585
R73 B.n469 B.n56 585
R74 B.n471 B.n470 585
R75 B.n473 B.n55 585
R76 B.n476 B.n475 585
R77 B.n477 B.n54 585
R78 B.n479 B.n478 585
R79 B.n481 B.n53 585
R80 B.n484 B.n483 585
R81 B.n485 B.n52 585
R82 B.n380 B.n50 585
R83 B.n488 B.n50 585
R84 B.n379 B.n49 585
R85 B.n489 B.n49 585
R86 B.n378 B.n48 585
R87 B.n490 B.n48 585
R88 B.n377 B.n376 585
R89 B.n376 B.n44 585
R90 B.n375 B.n43 585
R91 B.n496 B.n43 585
R92 B.n374 B.n42 585
R93 B.n497 B.n42 585
R94 B.n373 B.n41 585
R95 B.n498 B.n41 585
R96 B.n372 B.n371 585
R97 B.n371 B.n37 585
R98 B.n370 B.n36 585
R99 B.n504 B.n36 585
R100 B.n369 B.n35 585
R101 B.n505 B.n35 585
R102 B.n368 B.n34 585
R103 B.n506 B.n34 585
R104 B.n367 B.n366 585
R105 B.n366 B.n30 585
R106 B.n365 B.n29 585
R107 B.n512 B.n29 585
R108 B.n364 B.n28 585
R109 B.n513 B.n28 585
R110 B.n363 B.n27 585
R111 B.n514 B.n27 585
R112 B.n362 B.n361 585
R113 B.n361 B.n26 585
R114 B.n360 B.n22 585
R115 B.n520 B.n22 585
R116 B.n359 B.n21 585
R117 B.n521 B.n21 585
R118 B.n358 B.n20 585
R119 B.n522 B.n20 585
R120 B.n357 B.n356 585
R121 B.n356 B.n16 585
R122 B.n355 B.n15 585
R123 B.n528 B.n15 585
R124 B.n354 B.n14 585
R125 B.n529 B.n14 585
R126 B.n353 B.n13 585
R127 B.n530 B.n13 585
R128 B.n352 B.n351 585
R129 B.n351 B.n12 585
R130 B.n350 B.n349 585
R131 B.n350 B.n8 585
R132 B.n348 B.n7 585
R133 B.n537 B.n7 585
R134 B.n347 B.n6 585
R135 B.n538 B.n6 585
R136 B.n346 B.n5 585
R137 B.n539 B.n5 585
R138 B.n345 B.n344 585
R139 B.n344 B.n4 585
R140 B.n343 B.n83 585
R141 B.n343 B.n342 585
R142 B.n333 B.n84 585
R143 B.n85 B.n84 585
R144 B.n335 B.n334 585
R145 B.n336 B.n335 585
R146 B.n332 B.n89 585
R147 B.n93 B.n89 585
R148 B.n331 B.n330 585
R149 B.n330 B.n329 585
R150 B.n91 B.n90 585
R151 B.n92 B.n91 585
R152 B.n322 B.n321 585
R153 B.n323 B.n322 585
R154 B.n320 B.n98 585
R155 B.n98 B.n97 585
R156 B.n319 B.n318 585
R157 B.n318 B.n317 585
R158 B.n100 B.n99 585
R159 B.n310 B.n100 585
R160 B.n309 B.n308 585
R161 B.n311 B.n309 585
R162 B.n307 B.n105 585
R163 B.n105 B.n104 585
R164 B.n306 B.n305 585
R165 B.n305 B.n304 585
R166 B.n107 B.n106 585
R167 B.n108 B.n107 585
R168 B.n297 B.n296 585
R169 B.n298 B.n297 585
R170 B.n295 B.n113 585
R171 B.n113 B.n112 585
R172 B.n294 B.n293 585
R173 B.n293 B.n292 585
R174 B.n115 B.n114 585
R175 B.n116 B.n115 585
R176 B.n285 B.n284 585
R177 B.n286 B.n285 585
R178 B.n283 B.n121 585
R179 B.n121 B.n120 585
R180 B.n282 B.n281 585
R181 B.n281 B.n280 585
R182 B.n123 B.n122 585
R183 B.n124 B.n123 585
R184 B.n273 B.n272 585
R185 B.n274 B.n273 585
R186 B.n271 B.n129 585
R187 B.n129 B.n128 585
R188 B.n270 B.n269 585
R189 B.n269 B.n268 585
R190 B.n265 B.n133 585
R191 B.n264 B.n263 585
R192 B.n261 B.n134 585
R193 B.n261 B.n132 585
R194 B.n260 B.n259 585
R195 B.n258 B.n257 585
R196 B.n256 B.n136 585
R197 B.n254 B.n253 585
R198 B.n252 B.n137 585
R199 B.n251 B.n250 585
R200 B.n248 B.n138 585
R201 B.n246 B.n245 585
R202 B.n244 B.n139 585
R203 B.n243 B.n242 585
R204 B.n240 B.n140 585
R205 B.n238 B.n237 585
R206 B.n236 B.n141 585
R207 B.n235 B.n234 585
R208 B.n232 B.n142 585
R209 B.n230 B.n229 585
R210 B.n228 B.n143 585
R211 B.n227 B.n226 585
R212 B.n224 B.n223 585
R213 B.n222 B.n221 585
R214 B.n220 B.n148 585
R215 B.n218 B.n217 585
R216 B.n216 B.n149 585
R217 B.n215 B.n214 585
R218 B.n212 B.n150 585
R219 B.n210 B.n209 585
R220 B.n208 B.n151 585
R221 B.n207 B.n206 585
R222 B.n204 B.n203 585
R223 B.n202 B.n201 585
R224 B.n200 B.n156 585
R225 B.n198 B.n197 585
R226 B.n196 B.n157 585
R227 B.n195 B.n194 585
R228 B.n192 B.n158 585
R229 B.n190 B.n189 585
R230 B.n188 B.n159 585
R231 B.n187 B.n186 585
R232 B.n184 B.n160 585
R233 B.n182 B.n181 585
R234 B.n180 B.n161 585
R235 B.n179 B.n178 585
R236 B.n176 B.n162 585
R237 B.n174 B.n173 585
R238 B.n172 B.n163 585
R239 B.n171 B.n170 585
R240 B.n168 B.n164 585
R241 B.n166 B.n165 585
R242 B.n131 B.n130 585
R243 B.n132 B.n131 585
R244 B.n267 B.n266 585
R245 B.n268 B.n267 585
R246 B.n127 B.n126 585
R247 B.n128 B.n127 585
R248 B.n276 B.n275 585
R249 B.n275 B.n274 585
R250 B.n277 B.n125 585
R251 B.n125 B.n124 585
R252 B.n279 B.n278 585
R253 B.n280 B.n279 585
R254 B.n119 B.n118 585
R255 B.n120 B.n119 585
R256 B.n288 B.n287 585
R257 B.n287 B.n286 585
R258 B.n289 B.n117 585
R259 B.n117 B.n116 585
R260 B.n291 B.n290 585
R261 B.n292 B.n291 585
R262 B.n111 B.n110 585
R263 B.n112 B.n111 585
R264 B.n300 B.n299 585
R265 B.n299 B.n298 585
R266 B.n301 B.n109 585
R267 B.n109 B.n108 585
R268 B.n303 B.n302 585
R269 B.n304 B.n303 585
R270 B.n103 B.n102 585
R271 B.n104 B.n103 585
R272 B.n313 B.n312 585
R273 B.n312 B.n311 585
R274 B.n314 B.n101 585
R275 B.n310 B.n101 585
R276 B.n316 B.n315 585
R277 B.n317 B.n316 585
R278 B.n96 B.n95 585
R279 B.n97 B.n96 585
R280 B.n325 B.n324 585
R281 B.n324 B.n323 585
R282 B.n326 B.n94 585
R283 B.n94 B.n92 585
R284 B.n328 B.n327 585
R285 B.n329 B.n328 585
R286 B.n88 B.n87 585
R287 B.n93 B.n88 585
R288 B.n338 B.n337 585
R289 B.n337 B.n336 585
R290 B.n339 B.n86 585
R291 B.n86 B.n85 585
R292 B.n341 B.n340 585
R293 B.n342 B.n341 585
R294 B.n3 B.n0 585
R295 B.n4 B.n3 585
R296 B.n536 B.n1 585
R297 B.n537 B.n536 585
R298 B.n535 B.n534 585
R299 B.n535 B.n8 585
R300 B.n533 B.n9 585
R301 B.n12 B.n9 585
R302 B.n532 B.n531 585
R303 B.n531 B.n530 585
R304 B.n11 B.n10 585
R305 B.n529 B.n11 585
R306 B.n527 B.n526 585
R307 B.n528 B.n527 585
R308 B.n525 B.n17 585
R309 B.n17 B.n16 585
R310 B.n524 B.n523 585
R311 B.n523 B.n522 585
R312 B.n19 B.n18 585
R313 B.n521 B.n19 585
R314 B.n519 B.n518 585
R315 B.n520 B.n519 585
R316 B.n517 B.n23 585
R317 B.n26 B.n23 585
R318 B.n516 B.n515 585
R319 B.n515 B.n514 585
R320 B.n25 B.n24 585
R321 B.n513 B.n25 585
R322 B.n511 B.n510 585
R323 B.n512 B.n511 585
R324 B.n509 B.n31 585
R325 B.n31 B.n30 585
R326 B.n508 B.n507 585
R327 B.n507 B.n506 585
R328 B.n33 B.n32 585
R329 B.n505 B.n33 585
R330 B.n503 B.n502 585
R331 B.n504 B.n503 585
R332 B.n501 B.n38 585
R333 B.n38 B.n37 585
R334 B.n500 B.n499 585
R335 B.n499 B.n498 585
R336 B.n40 B.n39 585
R337 B.n497 B.n40 585
R338 B.n495 B.n494 585
R339 B.n496 B.n495 585
R340 B.n493 B.n45 585
R341 B.n45 B.n44 585
R342 B.n492 B.n491 585
R343 B.n491 B.n490 585
R344 B.n47 B.n46 585
R345 B.n489 B.n47 585
R346 B.n487 B.n486 585
R347 B.n488 B.n487 585
R348 B.n540 B.n539 585
R349 B.n538 B.n2 585
R350 B.n487 B.n52 554.963
R351 B.n382 B.n50 554.963
R352 B.n269 B.n131 554.963
R353 B.n267 B.n133 554.963
R354 B.n63 B.t15 275.401
R355 B.n71 B.t8 275.401
R356 B.n152 B.t12 275.401
R357 B.n144 B.t4 275.401
R358 B.n383 B.n51 256.663
R359 B.n385 B.n51 256.663
R360 B.n391 B.n51 256.663
R361 B.n393 B.n51 256.663
R362 B.n399 B.n51 256.663
R363 B.n401 B.n51 256.663
R364 B.n407 B.n51 256.663
R365 B.n409 B.n51 256.663
R366 B.n415 B.n51 256.663
R367 B.n417 B.n51 256.663
R368 B.n423 B.n51 256.663
R369 B.n425 B.n51 256.663
R370 B.n431 B.n51 256.663
R371 B.n433 B.n51 256.663
R372 B.n439 B.n51 256.663
R373 B.n441 B.n51 256.663
R374 B.n448 B.n51 256.663
R375 B.n450 B.n51 256.663
R376 B.n456 B.n51 256.663
R377 B.n458 B.n51 256.663
R378 B.n464 B.n51 256.663
R379 B.n466 B.n51 256.663
R380 B.n472 B.n51 256.663
R381 B.n474 B.n51 256.663
R382 B.n480 B.n51 256.663
R383 B.n482 B.n51 256.663
R384 B.n262 B.n132 256.663
R385 B.n135 B.n132 256.663
R386 B.n255 B.n132 256.663
R387 B.n249 B.n132 256.663
R388 B.n247 B.n132 256.663
R389 B.n241 B.n132 256.663
R390 B.n239 B.n132 256.663
R391 B.n233 B.n132 256.663
R392 B.n231 B.n132 256.663
R393 B.n225 B.n132 256.663
R394 B.n147 B.n132 256.663
R395 B.n219 B.n132 256.663
R396 B.n213 B.n132 256.663
R397 B.n211 B.n132 256.663
R398 B.n205 B.n132 256.663
R399 B.n155 B.n132 256.663
R400 B.n199 B.n132 256.663
R401 B.n193 B.n132 256.663
R402 B.n191 B.n132 256.663
R403 B.n185 B.n132 256.663
R404 B.n183 B.n132 256.663
R405 B.n177 B.n132 256.663
R406 B.n175 B.n132 256.663
R407 B.n169 B.n132 256.663
R408 B.n167 B.n132 256.663
R409 B.n542 B.n541 256.663
R410 B.n483 B.n481 163.367
R411 B.n479 B.n54 163.367
R412 B.n475 B.n473 163.367
R413 B.n471 B.n56 163.367
R414 B.n467 B.n465 163.367
R415 B.n463 B.n58 163.367
R416 B.n459 B.n457 163.367
R417 B.n455 B.n60 163.367
R418 B.n451 B.n449 163.367
R419 B.n447 B.n62 163.367
R420 B.n442 B.n440 163.367
R421 B.n438 B.n66 163.367
R422 B.n434 B.n432 163.367
R423 B.n430 B.n68 163.367
R424 B.n426 B.n424 163.367
R425 B.n422 B.n70 163.367
R426 B.n418 B.n416 163.367
R427 B.n414 B.n75 163.367
R428 B.n410 B.n408 163.367
R429 B.n406 B.n77 163.367
R430 B.n402 B.n400 163.367
R431 B.n398 B.n79 163.367
R432 B.n394 B.n392 163.367
R433 B.n390 B.n81 163.367
R434 B.n386 B.n384 163.367
R435 B.n269 B.n129 163.367
R436 B.n273 B.n129 163.367
R437 B.n273 B.n123 163.367
R438 B.n281 B.n123 163.367
R439 B.n281 B.n121 163.367
R440 B.n285 B.n121 163.367
R441 B.n285 B.n115 163.367
R442 B.n293 B.n115 163.367
R443 B.n293 B.n113 163.367
R444 B.n297 B.n113 163.367
R445 B.n297 B.n107 163.367
R446 B.n305 B.n107 163.367
R447 B.n305 B.n105 163.367
R448 B.n309 B.n105 163.367
R449 B.n309 B.n100 163.367
R450 B.n318 B.n100 163.367
R451 B.n318 B.n98 163.367
R452 B.n322 B.n98 163.367
R453 B.n322 B.n91 163.367
R454 B.n330 B.n91 163.367
R455 B.n330 B.n89 163.367
R456 B.n335 B.n89 163.367
R457 B.n335 B.n84 163.367
R458 B.n343 B.n84 163.367
R459 B.n344 B.n343 163.367
R460 B.n344 B.n5 163.367
R461 B.n6 B.n5 163.367
R462 B.n7 B.n6 163.367
R463 B.n350 B.n7 163.367
R464 B.n351 B.n350 163.367
R465 B.n351 B.n13 163.367
R466 B.n14 B.n13 163.367
R467 B.n15 B.n14 163.367
R468 B.n356 B.n15 163.367
R469 B.n356 B.n20 163.367
R470 B.n21 B.n20 163.367
R471 B.n22 B.n21 163.367
R472 B.n361 B.n22 163.367
R473 B.n361 B.n27 163.367
R474 B.n28 B.n27 163.367
R475 B.n29 B.n28 163.367
R476 B.n366 B.n29 163.367
R477 B.n366 B.n34 163.367
R478 B.n35 B.n34 163.367
R479 B.n36 B.n35 163.367
R480 B.n371 B.n36 163.367
R481 B.n371 B.n41 163.367
R482 B.n42 B.n41 163.367
R483 B.n43 B.n42 163.367
R484 B.n376 B.n43 163.367
R485 B.n376 B.n48 163.367
R486 B.n49 B.n48 163.367
R487 B.n50 B.n49 163.367
R488 B.n263 B.n261 163.367
R489 B.n261 B.n260 163.367
R490 B.n257 B.n256 163.367
R491 B.n254 B.n137 163.367
R492 B.n250 B.n248 163.367
R493 B.n246 B.n139 163.367
R494 B.n242 B.n240 163.367
R495 B.n238 B.n141 163.367
R496 B.n234 B.n232 163.367
R497 B.n230 B.n143 163.367
R498 B.n226 B.n224 163.367
R499 B.n221 B.n220 163.367
R500 B.n218 B.n149 163.367
R501 B.n214 B.n212 163.367
R502 B.n210 B.n151 163.367
R503 B.n206 B.n204 163.367
R504 B.n201 B.n200 163.367
R505 B.n198 B.n157 163.367
R506 B.n194 B.n192 163.367
R507 B.n190 B.n159 163.367
R508 B.n186 B.n184 163.367
R509 B.n182 B.n161 163.367
R510 B.n178 B.n176 163.367
R511 B.n174 B.n163 163.367
R512 B.n170 B.n168 163.367
R513 B.n166 B.n131 163.367
R514 B.n267 B.n127 163.367
R515 B.n275 B.n127 163.367
R516 B.n275 B.n125 163.367
R517 B.n279 B.n125 163.367
R518 B.n279 B.n119 163.367
R519 B.n287 B.n119 163.367
R520 B.n287 B.n117 163.367
R521 B.n291 B.n117 163.367
R522 B.n291 B.n111 163.367
R523 B.n299 B.n111 163.367
R524 B.n299 B.n109 163.367
R525 B.n303 B.n109 163.367
R526 B.n303 B.n103 163.367
R527 B.n312 B.n103 163.367
R528 B.n312 B.n101 163.367
R529 B.n316 B.n101 163.367
R530 B.n316 B.n96 163.367
R531 B.n324 B.n96 163.367
R532 B.n324 B.n94 163.367
R533 B.n328 B.n94 163.367
R534 B.n328 B.n88 163.367
R535 B.n337 B.n88 163.367
R536 B.n337 B.n86 163.367
R537 B.n341 B.n86 163.367
R538 B.n341 B.n3 163.367
R539 B.n540 B.n3 163.367
R540 B.n536 B.n2 163.367
R541 B.n536 B.n535 163.367
R542 B.n535 B.n9 163.367
R543 B.n531 B.n9 163.367
R544 B.n531 B.n11 163.367
R545 B.n527 B.n11 163.367
R546 B.n527 B.n17 163.367
R547 B.n523 B.n17 163.367
R548 B.n523 B.n19 163.367
R549 B.n519 B.n19 163.367
R550 B.n519 B.n23 163.367
R551 B.n515 B.n23 163.367
R552 B.n515 B.n25 163.367
R553 B.n511 B.n25 163.367
R554 B.n511 B.n31 163.367
R555 B.n507 B.n31 163.367
R556 B.n507 B.n33 163.367
R557 B.n503 B.n33 163.367
R558 B.n503 B.n38 163.367
R559 B.n499 B.n38 163.367
R560 B.n499 B.n40 163.367
R561 B.n495 B.n40 163.367
R562 B.n495 B.n45 163.367
R563 B.n491 B.n45 163.367
R564 B.n491 B.n47 163.367
R565 B.n487 B.n47 163.367
R566 B.n268 B.n132 147.375
R567 B.n488 B.n51 147.375
R568 B.n71 B.t10 117.626
R569 B.n152 B.t14 117.626
R570 B.n63 B.t16 117.621
R571 B.n144 B.t7 117.621
R572 B.n72 B.t11 76.7042
R573 B.n153 B.t13 76.7042
R574 B.n64 B.t17 76.6994
R575 B.n145 B.t6 76.6994
R576 B.n268 B.n128 72.0969
R577 B.n274 B.n128 72.0969
R578 B.n274 B.n124 72.0969
R579 B.n280 B.n124 72.0969
R580 B.n280 B.n120 72.0969
R581 B.n286 B.n120 72.0969
R582 B.n292 B.n116 72.0969
R583 B.n292 B.n112 72.0969
R584 B.n298 B.n112 72.0969
R585 B.n298 B.n108 72.0969
R586 B.n304 B.n108 72.0969
R587 B.n304 B.n104 72.0969
R588 B.n311 B.n104 72.0969
R589 B.n311 B.n310 72.0969
R590 B.n317 B.n97 72.0969
R591 B.n323 B.n97 72.0969
R592 B.n323 B.n92 72.0969
R593 B.n329 B.n92 72.0969
R594 B.n329 B.n93 72.0969
R595 B.n336 B.n85 72.0969
R596 B.n342 B.n85 72.0969
R597 B.n342 B.n4 72.0969
R598 B.n539 B.n4 72.0969
R599 B.n539 B.n538 72.0969
R600 B.n538 B.n537 72.0969
R601 B.n537 B.n8 72.0969
R602 B.n12 B.n8 72.0969
R603 B.n530 B.n12 72.0969
R604 B.n529 B.n528 72.0969
R605 B.n528 B.n16 72.0969
R606 B.n522 B.n16 72.0969
R607 B.n522 B.n521 72.0969
R608 B.n521 B.n520 72.0969
R609 B.n514 B.n26 72.0969
R610 B.n514 B.n513 72.0969
R611 B.n513 B.n512 72.0969
R612 B.n512 B.n30 72.0969
R613 B.n506 B.n30 72.0969
R614 B.n506 B.n505 72.0969
R615 B.n505 B.n504 72.0969
R616 B.n504 B.n37 72.0969
R617 B.n498 B.n497 72.0969
R618 B.n497 B.n496 72.0969
R619 B.n496 B.n44 72.0969
R620 B.n490 B.n44 72.0969
R621 B.n490 B.n489 72.0969
R622 B.n489 B.n488 72.0969
R623 B.n482 B.n52 71.676
R624 B.n481 B.n480 71.676
R625 B.n474 B.n54 71.676
R626 B.n473 B.n472 71.676
R627 B.n466 B.n56 71.676
R628 B.n465 B.n464 71.676
R629 B.n458 B.n58 71.676
R630 B.n457 B.n456 71.676
R631 B.n450 B.n60 71.676
R632 B.n449 B.n448 71.676
R633 B.n441 B.n62 71.676
R634 B.n440 B.n439 71.676
R635 B.n433 B.n66 71.676
R636 B.n432 B.n431 71.676
R637 B.n425 B.n68 71.676
R638 B.n424 B.n423 71.676
R639 B.n417 B.n70 71.676
R640 B.n416 B.n415 71.676
R641 B.n409 B.n75 71.676
R642 B.n408 B.n407 71.676
R643 B.n401 B.n77 71.676
R644 B.n400 B.n399 71.676
R645 B.n393 B.n79 71.676
R646 B.n392 B.n391 71.676
R647 B.n385 B.n81 71.676
R648 B.n384 B.n383 71.676
R649 B.n383 B.n382 71.676
R650 B.n386 B.n385 71.676
R651 B.n391 B.n390 71.676
R652 B.n394 B.n393 71.676
R653 B.n399 B.n398 71.676
R654 B.n402 B.n401 71.676
R655 B.n407 B.n406 71.676
R656 B.n410 B.n409 71.676
R657 B.n415 B.n414 71.676
R658 B.n418 B.n417 71.676
R659 B.n423 B.n422 71.676
R660 B.n426 B.n425 71.676
R661 B.n431 B.n430 71.676
R662 B.n434 B.n433 71.676
R663 B.n439 B.n438 71.676
R664 B.n442 B.n441 71.676
R665 B.n448 B.n447 71.676
R666 B.n451 B.n450 71.676
R667 B.n456 B.n455 71.676
R668 B.n459 B.n458 71.676
R669 B.n464 B.n463 71.676
R670 B.n467 B.n466 71.676
R671 B.n472 B.n471 71.676
R672 B.n475 B.n474 71.676
R673 B.n480 B.n479 71.676
R674 B.n483 B.n482 71.676
R675 B.n262 B.n133 71.676
R676 B.n260 B.n135 71.676
R677 B.n256 B.n255 71.676
R678 B.n249 B.n137 71.676
R679 B.n248 B.n247 71.676
R680 B.n241 B.n139 71.676
R681 B.n240 B.n239 71.676
R682 B.n233 B.n141 71.676
R683 B.n232 B.n231 71.676
R684 B.n225 B.n143 71.676
R685 B.n224 B.n147 71.676
R686 B.n220 B.n219 71.676
R687 B.n213 B.n149 71.676
R688 B.n212 B.n211 71.676
R689 B.n205 B.n151 71.676
R690 B.n204 B.n155 71.676
R691 B.n200 B.n199 71.676
R692 B.n193 B.n157 71.676
R693 B.n192 B.n191 71.676
R694 B.n185 B.n159 71.676
R695 B.n184 B.n183 71.676
R696 B.n177 B.n161 71.676
R697 B.n176 B.n175 71.676
R698 B.n169 B.n163 71.676
R699 B.n168 B.n167 71.676
R700 B.n263 B.n262 71.676
R701 B.n257 B.n135 71.676
R702 B.n255 B.n254 71.676
R703 B.n250 B.n249 71.676
R704 B.n247 B.n246 71.676
R705 B.n242 B.n241 71.676
R706 B.n239 B.n238 71.676
R707 B.n234 B.n233 71.676
R708 B.n231 B.n230 71.676
R709 B.n226 B.n225 71.676
R710 B.n221 B.n147 71.676
R711 B.n219 B.n218 71.676
R712 B.n214 B.n213 71.676
R713 B.n211 B.n210 71.676
R714 B.n206 B.n205 71.676
R715 B.n201 B.n155 71.676
R716 B.n199 B.n198 71.676
R717 B.n194 B.n193 71.676
R718 B.n191 B.n190 71.676
R719 B.n186 B.n185 71.676
R720 B.n183 B.n182 71.676
R721 B.n178 B.n177 71.676
R722 B.n175 B.n174 71.676
R723 B.n170 B.n169 71.676
R724 B.n167 B.n166 71.676
R725 B.n541 B.n540 71.676
R726 B.n541 B.n2 71.676
R727 B.n444 B.n64 59.5399
R728 B.n73 B.n72 59.5399
R729 B.n154 B.n153 59.5399
R730 B.n146 B.n145 59.5399
R731 B.t5 B.n116 59.374
R732 B.t9 B.n37 59.374
R733 B.n93 B.t1 57.2535
R734 B.t3 B.n529 57.2535
R735 B.n310 B.t0 42.4101
R736 B.n26 B.t2 42.4101
R737 B.n64 B.n63 40.9217
R738 B.n72 B.n71 40.9217
R739 B.n153 B.n152 40.9217
R740 B.n145 B.n144 40.9217
R741 B.n381 B.n380 36.059
R742 B.n266 B.n265 36.059
R743 B.n270 B.n130 36.059
R744 B.n486 B.n485 36.059
R745 B.n317 B.t0 29.6872
R746 B.n520 B.t2 29.6872
R747 B B.n542 18.0485
R748 B.n336 B.t1 14.8439
R749 B.n530 B.t3 14.8439
R750 B.n286 B.t5 12.7234
R751 B.n498 B.t9 12.7234
R752 B.n266 B.n126 10.6151
R753 B.n276 B.n126 10.6151
R754 B.n277 B.n276 10.6151
R755 B.n278 B.n277 10.6151
R756 B.n278 B.n118 10.6151
R757 B.n288 B.n118 10.6151
R758 B.n289 B.n288 10.6151
R759 B.n290 B.n289 10.6151
R760 B.n290 B.n110 10.6151
R761 B.n300 B.n110 10.6151
R762 B.n301 B.n300 10.6151
R763 B.n302 B.n301 10.6151
R764 B.n302 B.n102 10.6151
R765 B.n313 B.n102 10.6151
R766 B.n314 B.n313 10.6151
R767 B.n315 B.n314 10.6151
R768 B.n315 B.n95 10.6151
R769 B.n325 B.n95 10.6151
R770 B.n326 B.n325 10.6151
R771 B.n327 B.n326 10.6151
R772 B.n327 B.n87 10.6151
R773 B.n338 B.n87 10.6151
R774 B.n339 B.n338 10.6151
R775 B.n340 B.n339 10.6151
R776 B.n340 B.n0 10.6151
R777 B.n265 B.n264 10.6151
R778 B.n264 B.n134 10.6151
R779 B.n259 B.n134 10.6151
R780 B.n259 B.n258 10.6151
R781 B.n258 B.n136 10.6151
R782 B.n253 B.n136 10.6151
R783 B.n253 B.n252 10.6151
R784 B.n252 B.n251 10.6151
R785 B.n251 B.n138 10.6151
R786 B.n245 B.n138 10.6151
R787 B.n245 B.n244 10.6151
R788 B.n244 B.n243 10.6151
R789 B.n243 B.n140 10.6151
R790 B.n237 B.n140 10.6151
R791 B.n237 B.n236 10.6151
R792 B.n236 B.n235 10.6151
R793 B.n235 B.n142 10.6151
R794 B.n229 B.n142 10.6151
R795 B.n229 B.n228 10.6151
R796 B.n228 B.n227 10.6151
R797 B.n223 B.n222 10.6151
R798 B.n222 B.n148 10.6151
R799 B.n217 B.n148 10.6151
R800 B.n217 B.n216 10.6151
R801 B.n216 B.n215 10.6151
R802 B.n215 B.n150 10.6151
R803 B.n209 B.n150 10.6151
R804 B.n209 B.n208 10.6151
R805 B.n208 B.n207 10.6151
R806 B.n203 B.n202 10.6151
R807 B.n202 B.n156 10.6151
R808 B.n197 B.n156 10.6151
R809 B.n197 B.n196 10.6151
R810 B.n196 B.n195 10.6151
R811 B.n195 B.n158 10.6151
R812 B.n189 B.n158 10.6151
R813 B.n189 B.n188 10.6151
R814 B.n188 B.n187 10.6151
R815 B.n187 B.n160 10.6151
R816 B.n181 B.n160 10.6151
R817 B.n181 B.n180 10.6151
R818 B.n180 B.n179 10.6151
R819 B.n179 B.n162 10.6151
R820 B.n173 B.n162 10.6151
R821 B.n173 B.n172 10.6151
R822 B.n172 B.n171 10.6151
R823 B.n171 B.n164 10.6151
R824 B.n165 B.n164 10.6151
R825 B.n165 B.n130 10.6151
R826 B.n271 B.n270 10.6151
R827 B.n272 B.n271 10.6151
R828 B.n272 B.n122 10.6151
R829 B.n282 B.n122 10.6151
R830 B.n283 B.n282 10.6151
R831 B.n284 B.n283 10.6151
R832 B.n284 B.n114 10.6151
R833 B.n294 B.n114 10.6151
R834 B.n295 B.n294 10.6151
R835 B.n296 B.n295 10.6151
R836 B.n296 B.n106 10.6151
R837 B.n306 B.n106 10.6151
R838 B.n307 B.n306 10.6151
R839 B.n308 B.n307 10.6151
R840 B.n308 B.n99 10.6151
R841 B.n319 B.n99 10.6151
R842 B.n320 B.n319 10.6151
R843 B.n321 B.n320 10.6151
R844 B.n321 B.n90 10.6151
R845 B.n331 B.n90 10.6151
R846 B.n332 B.n331 10.6151
R847 B.n334 B.n332 10.6151
R848 B.n334 B.n333 10.6151
R849 B.n333 B.n83 10.6151
R850 B.n345 B.n83 10.6151
R851 B.n346 B.n345 10.6151
R852 B.n347 B.n346 10.6151
R853 B.n348 B.n347 10.6151
R854 B.n349 B.n348 10.6151
R855 B.n352 B.n349 10.6151
R856 B.n353 B.n352 10.6151
R857 B.n354 B.n353 10.6151
R858 B.n355 B.n354 10.6151
R859 B.n357 B.n355 10.6151
R860 B.n358 B.n357 10.6151
R861 B.n359 B.n358 10.6151
R862 B.n360 B.n359 10.6151
R863 B.n362 B.n360 10.6151
R864 B.n363 B.n362 10.6151
R865 B.n364 B.n363 10.6151
R866 B.n365 B.n364 10.6151
R867 B.n367 B.n365 10.6151
R868 B.n368 B.n367 10.6151
R869 B.n369 B.n368 10.6151
R870 B.n370 B.n369 10.6151
R871 B.n372 B.n370 10.6151
R872 B.n373 B.n372 10.6151
R873 B.n374 B.n373 10.6151
R874 B.n375 B.n374 10.6151
R875 B.n377 B.n375 10.6151
R876 B.n378 B.n377 10.6151
R877 B.n379 B.n378 10.6151
R878 B.n380 B.n379 10.6151
R879 B.n534 B.n1 10.6151
R880 B.n534 B.n533 10.6151
R881 B.n533 B.n532 10.6151
R882 B.n532 B.n10 10.6151
R883 B.n526 B.n10 10.6151
R884 B.n526 B.n525 10.6151
R885 B.n525 B.n524 10.6151
R886 B.n524 B.n18 10.6151
R887 B.n518 B.n18 10.6151
R888 B.n518 B.n517 10.6151
R889 B.n517 B.n516 10.6151
R890 B.n516 B.n24 10.6151
R891 B.n510 B.n24 10.6151
R892 B.n510 B.n509 10.6151
R893 B.n509 B.n508 10.6151
R894 B.n508 B.n32 10.6151
R895 B.n502 B.n32 10.6151
R896 B.n502 B.n501 10.6151
R897 B.n501 B.n500 10.6151
R898 B.n500 B.n39 10.6151
R899 B.n494 B.n39 10.6151
R900 B.n494 B.n493 10.6151
R901 B.n493 B.n492 10.6151
R902 B.n492 B.n46 10.6151
R903 B.n486 B.n46 10.6151
R904 B.n485 B.n484 10.6151
R905 B.n484 B.n53 10.6151
R906 B.n478 B.n53 10.6151
R907 B.n478 B.n477 10.6151
R908 B.n477 B.n476 10.6151
R909 B.n476 B.n55 10.6151
R910 B.n470 B.n55 10.6151
R911 B.n470 B.n469 10.6151
R912 B.n469 B.n468 10.6151
R913 B.n468 B.n57 10.6151
R914 B.n462 B.n57 10.6151
R915 B.n462 B.n461 10.6151
R916 B.n461 B.n460 10.6151
R917 B.n460 B.n59 10.6151
R918 B.n454 B.n59 10.6151
R919 B.n454 B.n453 10.6151
R920 B.n453 B.n452 10.6151
R921 B.n452 B.n61 10.6151
R922 B.n446 B.n61 10.6151
R923 B.n446 B.n445 10.6151
R924 B.n443 B.n65 10.6151
R925 B.n437 B.n65 10.6151
R926 B.n437 B.n436 10.6151
R927 B.n436 B.n435 10.6151
R928 B.n435 B.n67 10.6151
R929 B.n429 B.n67 10.6151
R930 B.n429 B.n428 10.6151
R931 B.n428 B.n427 10.6151
R932 B.n427 B.n69 10.6151
R933 B.n421 B.n420 10.6151
R934 B.n420 B.n419 10.6151
R935 B.n419 B.n74 10.6151
R936 B.n413 B.n74 10.6151
R937 B.n413 B.n412 10.6151
R938 B.n412 B.n411 10.6151
R939 B.n411 B.n76 10.6151
R940 B.n405 B.n76 10.6151
R941 B.n405 B.n404 10.6151
R942 B.n404 B.n403 10.6151
R943 B.n403 B.n78 10.6151
R944 B.n397 B.n78 10.6151
R945 B.n397 B.n396 10.6151
R946 B.n396 B.n395 10.6151
R947 B.n395 B.n80 10.6151
R948 B.n389 B.n80 10.6151
R949 B.n389 B.n388 10.6151
R950 B.n388 B.n387 10.6151
R951 B.n387 B.n82 10.6151
R952 B.n381 B.n82 10.6151
R953 B.n227 B.n146 9.36635
R954 B.n203 B.n154 9.36635
R955 B.n445 B.n444 9.36635
R956 B.n421 B.n73 9.36635
R957 B.n542 B.n0 8.11757
R958 B.n542 B.n1 8.11757
R959 B.n223 B.n146 1.24928
R960 B.n207 B.n154 1.24928
R961 B.n444 B.n443 1.24928
R962 B.n73 B.n69 1.24928
R963 VP.n5 VP.n4 183.188
R964 VP.n14 VP.n13 183.188
R965 VP.n12 VP.n0 161.3
R966 VP.n11 VP.n10 161.3
R967 VP.n9 VP.n1 161.3
R968 VP.n8 VP.n7 161.3
R969 VP.n6 VP.n2 161.3
R970 VP.n3 VP.t2 105.374
R971 VP.n3 VP.t1 104.945
R972 VP.n5 VP.t3 69.0511
R973 VP.n13 VP.t0 69.0511
R974 VP.n4 VP.n3 47.8102
R975 VP.n7 VP.n1 40.577
R976 VP.n11 VP.n1 40.577
R977 VP.n7 VP.n6 24.5923
R978 VP.n12 VP.n11 24.5923
R979 VP.n6 VP.n5 2.7056
R980 VP.n13 VP.n12 2.7056
R981 VP.n4 VP.n2 0.189894
R982 VP.n8 VP.n2 0.189894
R983 VP.n9 VP.n8 0.189894
R984 VP.n10 VP.n9 0.189894
R985 VP.n10 VP.n0 0.189894
R986 VP.n14 VP.n0 0.189894
R987 VP VP.n14 0.0516364
R988 VDD1 VDD1.n1 107.15
R989 VDD1 VDD1.n0 73.116
R990 VDD1.n0 VDD1.t1 3.88285
R991 VDD1.n0 VDD1.t2 3.88285
R992 VDD1.n1 VDD1.t0 3.88285
R993 VDD1.n1 VDD1.t3 3.88285
C0 VTAIL VDD2 3.54793f
C1 VDD1 VN 0.148415f
C2 VP VN 4.31911f
C3 VDD1 VDD2 0.826815f
C4 VP VDD2 0.346324f
C5 VTAIL VDD1 3.49922f
C6 VTAIL VP 2.23183f
C7 VP VDD1 2.2386f
C8 VN VDD2 2.0453f
C9 VTAIL VN 2.21773f
C10 VDD2 B 2.754925f
C11 VDD1 B 5.89742f
C12 VTAIL B 5.298665f
C13 VN B 8.538641f
C14 VP B 6.598629f
C15 VDD1.t1 B 0.109969f
C16 VDD1.t2 B 0.109969f
C17 VDD1.n0 B 0.89837f
C18 VDD1.t0 B 0.109969f
C19 VDD1.t3 B 0.109969f
C20 VDD1.n1 B 1.29205f
C21 VP.n0 B 0.03613f
C22 VP.t0 B 0.859104f
C23 VP.n1 B 0.029181f
C24 VP.n2 B 0.03613f
C25 VP.t3 B 0.859104f
C26 VP.t2 B 1.03582f
C27 VP.t1 B 1.03373f
C28 VP.n3 B 1.96718f
C29 VP.n4 B 1.62582f
C30 VP.n5 B 0.417978f
C31 VP.n6 B 0.037562f
C32 VP.n7 B 0.07143f
C33 VP.n8 B 0.03613f
C34 VP.n9 B 0.03613f
C35 VP.n10 B 0.03613f
C36 VP.n11 B 0.07143f
C37 VP.n12 B 0.037562f
C38 VP.n13 B 0.417978f
C39 VP.n14 B 0.038652f
C40 VDD2.t1 B 0.108021f
C41 VDD2.t3 B 0.108021f
C42 VDD2.n0 B 1.24791f
C43 VDD2.t2 B 0.108021f
C44 VDD2.t0 B 0.108021f
C45 VDD2.n1 B 0.882143f
C46 VDD2.n2 B 2.775f
C47 VTAIL.t7 B 0.754981f
C48 VTAIL.n0 B 0.307894f
C49 VTAIL.t1 B 0.754981f
C50 VTAIL.n1 B 0.360754f
C51 VTAIL.t0 B 0.754981f
C52 VTAIL.n2 B 0.979284f
C53 VTAIL.t6 B 0.754986f
C54 VTAIL.n3 B 0.979279f
C55 VTAIL.t4 B 0.754986f
C56 VTAIL.n4 B 0.360749f
C57 VTAIL.t3 B 0.754986f
C58 VTAIL.n5 B 0.360749f
C59 VTAIL.t2 B 0.754981f
C60 VTAIL.n6 B 0.979284f
C61 VTAIL.t5 B 0.754981f
C62 VTAIL.n7 B 0.919198f
C63 VN.t2 B 1.00613f
C64 VN.t0 B 1.00411f
C65 VN.n0 B 0.719326f
C66 VN.t3 B 1.00613f
C67 VN.t1 B 1.00411f
C68 VN.n1 B 1.93177f
.ends

