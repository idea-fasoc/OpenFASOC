* NGSPICE file created from diff_pair_sample_1376.ext - technology: sky130A

.subckt diff_pair_sample_1376 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
X1 VTAIL.t0 VP.t0 VDD1.t3 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X2 B.t11 B.t9 B.t10 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X3 VDD1.t2 VP.t1 VTAIL.t3 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
X4 B.t8 B.t6 B.t7 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X5 VDD2.t2 VN.t1 VTAIL.t5 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
X6 VTAIL.t6 VN.t2 VDD2.t1 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X7 VTAIL.t1 VP.t2 VDD1.t1 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X8 VTAIL.t4 VN.t3 VDD2.t0 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X9 B.t5 B.t3 B.t4 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X10 B.t2 B.t0 B.t1 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X11 VDD1.t0 VP.t3 VTAIL.t2 w_n2926_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
R0 VN.n1 VN.t1 112.889
R1 VN.n0 VN.t2 112.889
R2 VN.n0 VN.t0 111.913
R3 VN.n1 VN.t3 111.913
R4 VN VN.n1 48.7434
R5 VN VN.n0 3.12601
R6 VTAIL.n5 VTAIL.t0 63.3851
R7 VTAIL.n4 VTAIL.t5 63.3851
R8 VTAIL.n3 VTAIL.t4 63.3851
R9 VTAIL.n7 VTAIL.t7 63.385
R10 VTAIL.n0 VTAIL.t6 63.385
R11 VTAIL.n1 VTAIL.t2 63.385
R12 VTAIL.n2 VTAIL.t1 63.385
R13 VTAIL.n6 VTAIL.t3 63.385
R14 VTAIL.n7 VTAIL.n6 23.4014
R15 VTAIL.n3 VTAIL.n2 23.4014
R16 VTAIL.n4 VTAIL.n3 2.81084
R17 VTAIL.n6 VTAIL.n5 2.81084
R18 VTAIL.n2 VTAIL.n1 2.81084
R19 VTAIL VTAIL.n0 1.46386
R20 VTAIL VTAIL.n7 1.34748
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 117.026
R24 VDD2.n2 VDD2.n1 76.6566
R25 VDD2.n1 VDD2.t0 3.40773
R26 VDD2.n1 VDD2.t2 3.40773
R27 VDD2.n0 VDD2.t1 3.40773
R28 VDD2.n0 VDD2.t3 3.40773
R29 VDD2 VDD2.n2 0.0586897
R30 VP.n15 VP.n14 161.3
R31 VP.n13 VP.n1 161.3
R32 VP.n12 VP.n11 161.3
R33 VP.n10 VP.n2 161.3
R34 VP.n9 VP.n8 161.3
R35 VP.n7 VP.n3 161.3
R36 VP.n4 VP.t0 112.889
R37 VP.n4 VP.t1 111.913
R38 VP.n6 VP.t2 78.4694
R39 VP.n0 VP.t3 78.4694
R40 VP.n6 VP.n5 71.5558
R41 VP.n16 VP.n0 71.5558
R42 VP.n12 VP.n2 56.5617
R43 VP.n5 VP.n4 48.5782
R44 VP.n8 VP.n7 24.5923
R45 VP.n8 VP.n2 24.5923
R46 VP.n13 VP.n12 24.5923
R47 VP.n14 VP.n13 24.5923
R48 VP.n7 VP.n6 18.6903
R49 VP.n14 VP.n0 18.6903
R50 VP.n5 VP.n3 0.354861
R51 VP.n16 VP.n15 0.354861
R52 VP VP.n16 0.267071
R53 VP.n9 VP.n3 0.189894
R54 VP.n10 VP.n9 0.189894
R55 VP.n11 VP.n10 0.189894
R56 VP.n11 VP.n1 0.189894
R57 VP.n15 VP.n1 0.189894
R58 VDD1 VDD1.n1 117.552
R59 VDD1 VDD1.n0 76.7147
R60 VDD1.n0 VDD1.t3 3.40773
R61 VDD1.n0 VDD1.t2 3.40773
R62 VDD1.n1 VDD1.t1 3.40773
R63 VDD1.n1 VDD1.t0 3.40773
R64 B.n449 B.n64 585
R65 B.n451 B.n450 585
R66 B.n452 B.n63 585
R67 B.n454 B.n453 585
R68 B.n455 B.n62 585
R69 B.n457 B.n456 585
R70 B.n458 B.n61 585
R71 B.n460 B.n459 585
R72 B.n461 B.n60 585
R73 B.n463 B.n462 585
R74 B.n464 B.n59 585
R75 B.n466 B.n465 585
R76 B.n467 B.n58 585
R77 B.n469 B.n468 585
R78 B.n470 B.n57 585
R79 B.n472 B.n471 585
R80 B.n473 B.n56 585
R81 B.n475 B.n474 585
R82 B.n476 B.n55 585
R83 B.n478 B.n477 585
R84 B.n479 B.n54 585
R85 B.n481 B.n480 585
R86 B.n482 B.n53 585
R87 B.n484 B.n483 585
R88 B.n485 B.n52 585
R89 B.n487 B.n486 585
R90 B.n488 B.n51 585
R91 B.n490 B.n489 585
R92 B.n491 B.n50 585
R93 B.n493 B.n492 585
R94 B.n494 B.n49 585
R95 B.n496 B.n495 585
R96 B.n497 B.n45 585
R97 B.n499 B.n498 585
R98 B.n500 B.n44 585
R99 B.n502 B.n501 585
R100 B.n503 B.n43 585
R101 B.n505 B.n504 585
R102 B.n506 B.n42 585
R103 B.n508 B.n507 585
R104 B.n509 B.n41 585
R105 B.n511 B.n510 585
R106 B.n512 B.n40 585
R107 B.n514 B.n513 585
R108 B.n516 B.n37 585
R109 B.n518 B.n517 585
R110 B.n519 B.n36 585
R111 B.n521 B.n520 585
R112 B.n522 B.n35 585
R113 B.n524 B.n523 585
R114 B.n525 B.n34 585
R115 B.n527 B.n526 585
R116 B.n528 B.n33 585
R117 B.n530 B.n529 585
R118 B.n531 B.n32 585
R119 B.n533 B.n532 585
R120 B.n534 B.n31 585
R121 B.n536 B.n535 585
R122 B.n537 B.n30 585
R123 B.n539 B.n538 585
R124 B.n540 B.n29 585
R125 B.n542 B.n541 585
R126 B.n543 B.n28 585
R127 B.n545 B.n544 585
R128 B.n546 B.n27 585
R129 B.n548 B.n547 585
R130 B.n549 B.n26 585
R131 B.n551 B.n550 585
R132 B.n552 B.n25 585
R133 B.n554 B.n553 585
R134 B.n555 B.n24 585
R135 B.n557 B.n556 585
R136 B.n558 B.n23 585
R137 B.n560 B.n559 585
R138 B.n561 B.n22 585
R139 B.n563 B.n562 585
R140 B.n564 B.n21 585
R141 B.n566 B.n565 585
R142 B.n448 B.n447 585
R143 B.n446 B.n65 585
R144 B.n445 B.n444 585
R145 B.n443 B.n66 585
R146 B.n442 B.n441 585
R147 B.n440 B.n67 585
R148 B.n439 B.n438 585
R149 B.n437 B.n68 585
R150 B.n436 B.n435 585
R151 B.n434 B.n69 585
R152 B.n433 B.n432 585
R153 B.n431 B.n70 585
R154 B.n430 B.n429 585
R155 B.n428 B.n71 585
R156 B.n427 B.n426 585
R157 B.n425 B.n72 585
R158 B.n424 B.n423 585
R159 B.n422 B.n73 585
R160 B.n421 B.n420 585
R161 B.n419 B.n74 585
R162 B.n418 B.n417 585
R163 B.n416 B.n75 585
R164 B.n415 B.n414 585
R165 B.n413 B.n76 585
R166 B.n412 B.n411 585
R167 B.n410 B.n77 585
R168 B.n409 B.n408 585
R169 B.n407 B.n78 585
R170 B.n406 B.n405 585
R171 B.n404 B.n79 585
R172 B.n403 B.n402 585
R173 B.n401 B.n80 585
R174 B.n400 B.n399 585
R175 B.n398 B.n81 585
R176 B.n397 B.n396 585
R177 B.n395 B.n82 585
R178 B.n394 B.n393 585
R179 B.n392 B.n83 585
R180 B.n391 B.n390 585
R181 B.n389 B.n84 585
R182 B.n388 B.n387 585
R183 B.n386 B.n85 585
R184 B.n385 B.n384 585
R185 B.n383 B.n86 585
R186 B.n382 B.n381 585
R187 B.n380 B.n87 585
R188 B.n379 B.n378 585
R189 B.n377 B.n88 585
R190 B.n376 B.n375 585
R191 B.n374 B.n89 585
R192 B.n373 B.n372 585
R193 B.n371 B.n90 585
R194 B.n370 B.n369 585
R195 B.n368 B.n91 585
R196 B.n367 B.n366 585
R197 B.n365 B.n92 585
R198 B.n364 B.n363 585
R199 B.n362 B.n93 585
R200 B.n361 B.n360 585
R201 B.n359 B.n94 585
R202 B.n358 B.n357 585
R203 B.n356 B.n95 585
R204 B.n355 B.n354 585
R205 B.n353 B.n96 585
R206 B.n352 B.n351 585
R207 B.n350 B.n97 585
R208 B.n349 B.n348 585
R209 B.n347 B.n98 585
R210 B.n346 B.n345 585
R211 B.n344 B.n99 585
R212 B.n343 B.n342 585
R213 B.n341 B.n100 585
R214 B.n340 B.n339 585
R215 B.n338 B.n101 585
R216 B.n337 B.n336 585
R217 B.n218 B.n145 585
R218 B.n220 B.n219 585
R219 B.n221 B.n144 585
R220 B.n223 B.n222 585
R221 B.n224 B.n143 585
R222 B.n226 B.n225 585
R223 B.n227 B.n142 585
R224 B.n229 B.n228 585
R225 B.n230 B.n141 585
R226 B.n232 B.n231 585
R227 B.n233 B.n140 585
R228 B.n235 B.n234 585
R229 B.n236 B.n139 585
R230 B.n238 B.n237 585
R231 B.n239 B.n138 585
R232 B.n241 B.n240 585
R233 B.n242 B.n137 585
R234 B.n244 B.n243 585
R235 B.n245 B.n136 585
R236 B.n247 B.n246 585
R237 B.n248 B.n135 585
R238 B.n250 B.n249 585
R239 B.n251 B.n134 585
R240 B.n253 B.n252 585
R241 B.n254 B.n133 585
R242 B.n256 B.n255 585
R243 B.n257 B.n132 585
R244 B.n259 B.n258 585
R245 B.n260 B.n131 585
R246 B.n262 B.n261 585
R247 B.n263 B.n130 585
R248 B.n265 B.n264 585
R249 B.n266 B.n129 585
R250 B.n268 B.n267 585
R251 B.n270 B.n126 585
R252 B.n272 B.n271 585
R253 B.n273 B.n125 585
R254 B.n275 B.n274 585
R255 B.n276 B.n124 585
R256 B.n278 B.n277 585
R257 B.n279 B.n123 585
R258 B.n281 B.n280 585
R259 B.n282 B.n122 585
R260 B.n284 B.n283 585
R261 B.n286 B.n285 585
R262 B.n287 B.n118 585
R263 B.n289 B.n288 585
R264 B.n290 B.n117 585
R265 B.n292 B.n291 585
R266 B.n293 B.n116 585
R267 B.n295 B.n294 585
R268 B.n296 B.n115 585
R269 B.n298 B.n297 585
R270 B.n299 B.n114 585
R271 B.n301 B.n300 585
R272 B.n302 B.n113 585
R273 B.n304 B.n303 585
R274 B.n305 B.n112 585
R275 B.n307 B.n306 585
R276 B.n308 B.n111 585
R277 B.n310 B.n309 585
R278 B.n311 B.n110 585
R279 B.n313 B.n312 585
R280 B.n314 B.n109 585
R281 B.n316 B.n315 585
R282 B.n317 B.n108 585
R283 B.n319 B.n318 585
R284 B.n320 B.n107 585
R285 B.n322 B.n321 585
R286 B.n323 B.n106 585
R287 B.n325 B.n324 585
R288 B.n326 B.n105 585
R289 B.n328 B.n327 585
R290 B.n329 B.n104 585
R291 B.n331 B.n330 585
R292 B.n332 B.n103 585
R293 B.n334 B.n333 585
R294 B.n335 B.n102 585
R295 B.n217 B.n216 585
R296 B.n215 B.n146 585
R297 B.n214 B.n213 585
R298 B.n212 B.n147 585
R299 B.n211 B.n210 585
R300 B.n209 B.n148 585
R301 B.n208 B.n207 585
R302 B.n206 B.n149 585
R303 B.n205 B.n204 585
R304 B.n203 B.n150 585
R305 B.n202 B.n201 585
R306 B.n200 B.n151 585
R307 B.n199 B.n198 585
R308 B.n197 B.n152 585
R309 B.n196 B.n195 585
R310 B.n194 B.n153 585
R311 B.n193 B.n192 585
R312 B.n191 B.n154 585
R313 B.n190 B.n189 585
R314 B.n188 B.n155 585
R315 B.n187 B.n186 585
R316 B.n185 B.n156 585
R317 B.n184 B.n183 585
R318 B.n182 B.n157 585
R319 B.n181 B.n180 585
R320 B.n179 B.n158 585
R321 B.n178 B.n177 585
R322 B.n176 B.n159 585
R323 B.n175 B.n174 585
R324 B.n173 B.n160 585
R325 B.n172 B.n171 585
R326 B.n170 B.n161 585
R327 B.n169 B.n168 585
R328 B.n167 B.n162 585
R329 B.n166 B.n165 585
R330 B.n164 B.n163 585
R331 B.n2 B.n0 585
R332 B.n621 B.n1 585
R333 B.n620 B.n619 585
R334 B.n618 B.n3 585
R335 B.n617 B.n616 585
R336 B.n615 B.n4 585
R337 B.n614 B.n613 585
R338 B.n612 B.n5 585
R339 B.n611 B.n610 585
R340 B.n609 B.n6 585
R341 B.n608 B.n607 585
R342 B.n606 B.n7 585
R343 B.n605 B.n604 585
R344 B.n603 B.n8 585
R345 B.n602 B.n601 585
R346 B.n600 B.n9 585
R347 B.n599 B.n598 585
R348 B.n597 B.n10 585
R349 B.n596 B.n595 585
R350 B.n594 B.n11 585
R351 B.n593 B.n592 585
R352 B.n591 B.n12 585
R353 B.n590 B.n589 585
R354 B.n588 B.n13 585
R355 B.n587 B.n586 585
R356 B.n585 B.n14 585
R357 B.n584 B.n583 585
R358 B.n582 B.n15 585
R359 B.n581 B.n580 585
R360 B.n579 B.n16 585
R361 B.n578 B.n577 585
R362 B.n576 B.n17 585
R363 B.n575 B.n574 585
R364 B.n573 B.n18 585
R365 B.n572 B.n571 585
R366 B.n570 B.n19 585
R367 B.n569 B.n568 585
R368 B.n567 B.n20 585
R369 B.n623 B.n622 585
R370 B.n218 B.n217 506.916
R371 B.n567 B.n566 506.916
R372 B.n337 B.n102 506.916
R373 B.n447 B.n64 506.916
R374 B.n119 B.t6 286.966
R375 B.n127 B.t0 286.966
R376 B.n38 B.t9 286.966
R377 B.n46 B.t3 286.966
R378 B.n119 B.t8 171.458
R379 B.n46 B.t4 171.458
R380 B.n127 B.t2 171.447
R381 B.n38 B.t10 171.447
R382 B.n217 B.n146 163.367
R383 B.n213 B.n146 163.367
R384 B.n213 B.n212 163.367
R385 B.n212 B.n211 163.367
R386 B.n211 B.n148 163.367
R387 B.n207 B.n148 163.367
R388 B.n207 B.n206 163.367
R389 B.n206 B.n205 163.367
R390 B.n205 B.n150 163.367
R391 B.n201 B.n150 163.367
R392 B.n201 B.n200 163.367
R393 B.n200 B.n199 163.367
R394 B.n199 B.n152 163.367
R395 B.n195 B.n152 163.367
R396 B.n195 B.n194 163.367
R397 B.n194 B.n193 163.367
R398 B.n193 B.n154 163.367
R399 B.n189 B.n154 163.367
R400 B.n189 B.n188 163.367
R401 B.n188 B.n187 163.367
R402 B.n187 B.n156 163.367
R403 B.n183 B.n156 163.367
R404 B.n183 B.n182 163.367
R405 B.n182 B.n181 163.367
R406 B.n181 B.n158 163.367
R407 B.n177 B.n158 163.367
R408 B.n177 B.n176 163.367
R409 B.n176 B.n175 163.367
R410 B.n175 B.n160 163.367
R411 B.n171 B.n160 163.367
R412 B.n171 B.n170 163.367
R413 B.n170 B.n169 163.367
R414 B.n169 B.n162 163.367
R415 B.n165 B.n162 163.367
R416 B.n165 B.n164 163.367
R417 B.n164 B.n2 163.367
R418 B.n622 B.n2 163.367
R419 B.n622 B.n621 163.367
R420 B.n621 B.n620 163.367
R421 B.n620 B.n3 163.367
R422 B.n616 B.n3 163.367
R423 B.n616 B.n615 163.367
R424 B.n615 B.n614 163.367
R425 B.n614 B.n5 163.367
R426 B.n610 B.n5 163.367
R427 B.n610 B.n609 163.367
R428 B.n609 B.n608 163.367
R429 B.n608 B.n7 163.367
R430 B.n604 B.n7 163.367
R431 B.n604 B.n603 163.367
R432 B.n603 B.n602 163.367
R433 B.n602 B.n9 163.367
R434 B.n598 B.n9 163.367
R435 B.n598 B.n597 163.367
R436 B.n597 B.n596 163.367
R437 B.n596 B.n11 163.367
R438 B.n592 B.n11 163.367
R439 B.n592 B.n591 163.367
R440 B.n591 B.n590 163.367
R441 B.n590 B.n13 163.367
R442 B.n586 B.n13 163.367
R443 B.n586 B.n585 163.367
R444 B.n585 B.n584 163.367
R445 B.n584 B.n15 163.367
R446 B.n580 B.n15 163.367
R447 B.n580 B.n579 163.367
R448 B.n579 B.n578 163.367
R449 B.n578 B.n17 163.367
R450 B.n574 B.n17 163.367
R451 B.n574 B.n573 163.367
R452 B.n573 B.n572 163.367
R453 B.n572 B.n19 163.367
R454 B.n568 B.n19 163.367
R455 B.n568 B.n567 163.367
R456 B.n219 B.n218 163.367
R457 B.n219 B.n144 163.367
R458 B.n223 B.n144 163.367
R459 B.n224 B.n223 163.367
R460 B.n225 B.n224 163.367
R461 B.n225 B.n142 163.367
R462 B.n229 B.n142 163.367
R463 B.n230 B.n229 163.367
R464 B.n231 B.n230 163.367
R465 B.n231 B.n140 163.367
R466 B.n235 B.n140 163.367
R467 B.n236 B.n235 163.367
R468 B.n237 B.n236 163.367
R469 B.n237 B.n138 163.367
R470 B.n241 B.n138 163.367
R471 B.n242 B.n241 163.367
R472 B.n243 B.n242 163.367
R473 B.n243 B.n136 163.367
R474 B.n247 B.n136 163.367
R475 B.n248 B.n247 163.367
R476 B.n249 B.n248 163.367
R477 B.n249 B.n134 163.367
R478 B.n253 B.n134 163.367
R479 B.n254 B.n253 163.367
R480 B.n255 B.n254 163.367
R481 B.n255 B.n132 163.367
R482 B.n259 B.n132 163.367
R483 B.n260 B.n259 163.367
R484 B.n261 B.n260 163.367
R485 B.n261 B.n130 163.367
R486 B.n265 B.n130 163.367
R487 B.n266 B.n265 163.367
R488 B.n267 B.n266 163.367
R489 B.n267 B.n126 163.367
R490 B.n272 B.n126 163.367
R491 B.n273 B.n272 163.367
R492 B.n274 B.n273 163.367
R493 B.n274 B.n124 163.367
R494 B.n278 B.n124 163.367
R495 B.n279 B.n278 163.367
R496 B.n280 B.n279 163.367
R497 B.n280 B.n122 163.367
R498 B.n284 B.n122 163.367
R499 B.n285 B.n284 163.367
R500 B.n285 B.n118 163.367
R501 B.n289 B.n118 163.367
R502 B.n290 B.n289 163.367
R503 B.n291 B.n290 163.367
R504 B.n291 B.n116 163.367
R505 B.n295 B.n116 163.367
R506 B.n296 B.n295 163.367
R507 B.n297 B.n296 163.367
R508 B.n297 B.n114 163.367
R509 B.n301 B.n114 163.367
R510 B.n302 B.n301 163.367
R511 B.n303 B.n302 163.367
R512 B.n303 B.n112 163.367
R513 B.n307 B.n112 163.367
R514 B.n308 B.n307 163.367
R515 B.n309 B.n308 163.367
R516 B.n309 B.n110 163.367
R517 B.n313 B.n110 163.367
R518 B.n314 B.n313 163.367
R519 B.n315 B.n314 163.367
R520 B.n315 B.n108 163.367
R521 B.n319 B.n108 163.367
R522 B.n320 B.n319 163.367
R523 B.n321 B.n320 163.367
R524 B.n321 B.n106 163.367
R525 B.n325 B.n106 163.367
R526 B.n326 B.n325 163.367
R527 B.n327 B.n326 163.367
R528 B.n327 B.n104 163.367
R529 B.n331 B.n104 163.367
R530 B.n332 B.n331 163.367
R531 B.n333 B.n332 163.367
R532 B.n333 B.n102 163.367
R533 B.n338 B.n337 163.367
R534 B.n339 B.n338 163.367
R535 B.n339 B.n100 163.367
R536 B.n343 B.n100 163.367
R537 B.n344 B.n343 163.367
R538 B.n345 B.n344 163.367
R539 B.n345 B.n98 163.367
R540 B.n349 B.n98 163.367
R541 B.n350 B.n349 163.367
R542 B.n351 B.n350 163.367
R543 B.n351 B.n96 163.367
R544 B.n355 B.n96 163.367
R545 B.n356 B.n355 163.367
R546 B.n357 B.n356 163.367
R547 B.n357 B.n94 163.367
R548 B.n361 B.n94 163.367
R549 B.n362 B.n361 163.367
R550 B.n363 B.n362 163.367
R551 B.n363 B.n92 163.367
R552 B.n367 B.n92 163.367
R553 B.n368 B.n367 163.367
R554 B.n369 B.n368 163.367
R555 B.n369 B.n90 163.367
R556 B.n373 B.n90 163.367
R557 B.n374 B.n373 163.367
R558 B.n375 B.n374 163.367
R559 B.n375 B.n88 163.367
R560 B.n379 B.n88 163.367
R561 B.n380 B.n379 163.367
R562 B.n381 B.n380 163.367
R563 B.n381 B.n86 163.367
R564 B.n385 B.n86 163.367
R565 B.n386 B.n385 163.367
R566 B.n387 B.n386 163.367
R567 B.n387 B.n84 163.367
R568 B.n391 B.n84 163.367
R569 B.n392 B.n391 163.367
R570 B.n393 B.n392 163.367
R571 B.n393 B.n82 163.367
R572 B.n397 B.n82 163.367
R573 B.n398 B.n397 163.367
R574 B.n399 B.n398 163.367
R575 B.n399 B.n80 163.367
R576 B.n403 B.n80 163.367
R577 B.n404 B.n403 163.367
R578 B.n405 B.n404 163.367
R579 B.n405 B.n78 163.367
R580 B.n409 B.n78 163.367
R581 B.n410 B.n409 163.367
R582 B.n411 B.n410 163.367
R583 B.n411 B.n76 163.367
R584 B.n415 B.n76 163.367
R585 B.n416 B.n415 163.367
R586 B.n417 B.n416 163.367
R587 B.n417 B.n74 163.367
R588 B.n421 B.n74 163.367
R589 B.n422 B.n421 163.367
R590 B.n423 B.n422 163.367
R591 B.n423 B.n72 163.367
R592 B.n427 B.n72 163.367
R593 B.n428 B.n427 163.367
R594 B.n429 B.n428 163.367
R595 B.n429 B.n70 163.367
R596 B.n433 B.n70 163.367
R597 B.n434 B.n433 163.367
R598 B.n435 B.n434 163.367
R599 B.n435 B.n68 163.367
R600 B.n439 B.n68 163.367
R601 B.n440 B.n439 163.367
R602 B.n441 B.n440 163.367
R603 B.n441 B.n66 163.367
R604 B.n445 B.n66 163.367
R605 B.n446 B.n445 163.367
R606 B.n447 B.n446 163.367
R607 B.n566 B.n21 163.367
R608 B.n562 B.n21 163.367
R609 B.n562 B.n561 163.367
R610 B.n561 B.n560 163.367
R611 B.n560 B.n23 163.367
R612 B.n556 B.n23 163.367
R613 B.n556 B.n555 163.367
R614 B.n555 B.n554 163.367
R615 B.n554 B.n25 163.367
R616 B.n550 B.n25 163.367
R617 B.n550 B.n549 163.367
R618 B.n549 B.n548 163.367
R619 B.n548 B.n27 163.367
R620 B.n544 B.n27 163.367
R621 B.n544 B.n543 163.367
R622 B.n543 B.n542 163.367
R623 B.n542 B.n29 163.367
R624 B.n538 B.n29 163.367
R625 B.n538 B.n537 163.367
R626 B.n537 B.n536 163.367
R627 B.n536 B.n31 163.367
R628 B.n532 B.n31 163.367
R629 B.n532 B.n531 163.367
R630 B.n531 B.n530 163.367
R631 B.n530 B.n33 163.367
R632 B.n526 B.n33 163.367
R633 B.n526 B.n525 163.367
R634 B.n525 B.n524 163.367
R635 B.n524 B.n35 163.367
R636 B.n520 B.n35 163.367
R637 B.n520 B.n519 163.367
R638 B.n519 B.n518 163.367
R639 B.n518 B.n37 163.367
R640 B.n513 B.n37 163.367
R641 B.n513 B.n512 163.367
R642 B.n512 B.n511 163.367
R643 B.n511 B.n41 163.367
R644 B.n507 B.n41 163.367
R645 B.n507 B.n506 163.367
R646 B.n506 B.n505 163.367
R647 B.n505 B.n43 163.367
R648 B.n501 B.n43 163.367
R649 B.n501 B.n500 163.367
R650 B.n500 B.n499 163.367
R651 B.n499 B.n45 163.367
R652 B.n495 B.n45 163.367
R653 B.n495 B.n494 163.367
R654 B.n494 B.n493 163.367
R655 B.n493 B.n50 163.367
R656 B.n489 B.n50 163.367
R657 B.n489 B.n488 163.367
R658 B.n488 B.n487 163.367
R659 B.n487 B.n52 163.367
R660 B.n483 B.n52 163.367
R661 B.n483 B.n482 163.367
R662 B.n482 B.n481 163.367
R663 B.n481 B.n54 163.367
R664 B.n477 B.n54 163.367
R665 B.n477 B.n476 163.367
R666 B.n476 B.n475 163.367
R667 B.n475 B.n56 163.367
R668 B.n471 B.n56 163.367
R669 B.n471 B.n470 163.367
R670 B.n470 B.n469 163.367
R671 B.n469 B.n58 163.367
R672 B.n465 B.n58 163.367
R673 B.n465 B.n464 163.367
R674 B.n464 B.n463 163.367
R675 B.n463 B.n60 163.367
R676 B.n459 B.n60 163.367
R677 B.n459 B.n458 163.367
R678 B.n458 B.n457 163.367
R679 B.n457 B.n62 163.367
R680 B.n453 B.n62 163.367
R681 B.n453 B.n452 163.367
R682 B.n452 B.n451 163.367
R683 B.n451 B.n64 163.367
R684 B.n120 B.t7 108.234
R685 B.n47 B.t5 108.234
R686 B.n128 B.t1 108.224
R687 B.n39 B.t11 108.224
R688 B.n120 B.n119 63.2247
R689 B.n128 B.n127 63.2247
R690 B.n39 B.n38 63.2247
R691 B.n47 B.n46 63.2247
R692 B.n121 B.n120 59.5399
R693 B.n269 B.n128 59.5399
R694 B.n515 B.n39 59.5399
R695 B.n48 B.n47 59.5399
R696 B.n565 B.n20 32.9371
R697 B.n449 B.n448 32.9371
R698 B.n336 B.n335 32.9371
R699 B.n216 B.n145 32.9371
R700 B B.n623 18.0485
R701 B.n565 B.n564 10.6151
R702 B.n564 B.n563 10.6151
R703 B.n563 B.n22 10.6151
R704 B.n559 B.n22 10.6151
R705 B.n559 B.n558 10.6151
R706 B.n558 B.n557 10.6151
R707 B.n557 B.n24 10.6151
R708 B.n553 B.n24 10.6151
R709 B.n553 B.n552 10.6151
R710 B.n552 B.n551 10.6151
R711 B.n551 B.n26 10.6151
R712 B.n547 B.n26 10.6151
R713 B.n547 B.n546 10.6151
R714 B.n546 B.n545 10.6151
R715 B.n545 B.n28 10.6151
R716 B.n541 B.n28 10.6151
R717 B.n541 B.n540 10.6151
R718 B.n540 B.n539 10.6151
R719 B.n539 B.n30 10.6151
R720 B.n535 B.n30 10.6151
R721 B.n535 B.n534 10.6151
R722 B.n534 B.n533 10.6151
R723 B.n533 B.n32 10.6151
R724 B.n529 B.n32 10.6151
R725 B.n529 B.n528 10.6151
R726 B.n528 B.n527 10.6151
R727 B.n527 B.n34 10.6151
R728 B.n523 B.n34 10.6151
R729 B.n523 B.n522 10.6151
R730 B.n522 B.n521 10.6151
R731 B.n521 B.n36 10.6151
R732 B.n517 B.n36 10.6151
R733 B.n517 B.n516 10.6151
R734 B.n514 B.n40 10.6151
R735 B.n510 B.n40 10.6151
R736 B.n510 B.n509 10.6151
R737 B.n509 B.n508 10.6151
R738 B.n508 B.n42 10.6151
R739 B.n504 B.n42 10.6151
R740 B.n504 B.n503 10.6151
R741 B.n503 B.n502 10.6151
R742 B.n502 B.n44 10.6151
R743 B.n498 B.n497 10.6151
R744 B.n497 B.n496 10.6151
R745 B.n496 B.n49 10.6151
R746 B.n492 B.n49 10.6151
R747 B.n492 B.n491 10.6151
R748 B.n491 B.n490 10.6151
R749 B.n490 B.n51 10.6151
R750 B.n486 B.n51 10.6151
R751 B.n486 B.n485 10.6151
R752 B.n485 B.n484 10.6151
R753 B.n484 B.n53 10.6151
R754 B.n480 B.n53 10.6151
R755 B.n480 B.n479 10.6151
R756 B.n479 B.n478 10.6151
R757 B.n478 B.n55 10.6151
R758 B.n474 B.n55 10.6151
R759 B.n474 B.n473 10.6151
R760 B.n473 B.n472 10.6151
R761 B.n472 B.n57 10.6151
R762 B.n468 B.n57 10.6151
R763 B.n468 B.n467 10.6151
R764 B.n467 B.n466 10.6151
R765 B.n466 B.n59 10.6151
R766 B.n462 B.n59 10.6151
R767 B.n462 B.n461 10.6151
R768 B.n461 B.n460 10.6151
R769 B.n460 B.n61 10.6151
R770 B.n456 B.n61 10.6151
R771 B.n456 B.n455 10.6151
R772 B.n455 B.n454 10.6151
R773 B.n454 B.n63 10.6151
R774 B.n450 B.n63 10.6151
R775 B.n450 B.n449 10.6151
R776 B.n336 B.n101 10.6151
R777 B.n340 B.n101 10.6151
R778 B.n341 B.n340 10.6151
R779 B.n342 B.n341 10.6151
R780 B.n342 B.n99 10.6151
R781 B.n346 B.n99 10.6151
R782 B.n347 B.n346 10.6151
R783 B.n348 B.n347 10.6151
R784 B.n348 B.n97 10.6151
R785 B.n352 B.n97 10.6151
R786 B.n353 B.n352 10.6151
R787 B.n354 B.n353 10.6151
R788 B.n354 B.n95 10.6151
R789 B.n358 B.n95 10.6151
R790 B.n359 B.n358 10.6151
R791 B.n360 B.n359 10.6151
R792 B.n360 B.n93 10.6151
R793 B.n364 B.n93 10.6151
R794 B.n365 B.n364 10.6151
R795 B.n366 B.n365 10.6151
R796 B.n366 B.n91 10.6151
R797 B.n370 B.n91 10.6151
R798 B.n371 B.n370 10.6151
R799 B.n372 B.n371 10.6151
R800 B.n372 B.n89 10.6151
R801 B.n376 B.n89 10.6151
R802 B.n377 B.n376 10.6151
R803 B.n378 B.n377 10.6151
R804 B.n378 B.n87 10.6151
R805 B.n382 B.n87 10.6151
R806 B.n383 B.n382 10.6151
R807 B.n384 B.n383 10.6151
R808 B.n384 B.n85 10.6151
R809 B.n388 B.n85 10.6151
R810 B.n389 B.n388 10.6151
R811 B.n390 B.n389 10.6151
R812 B.n390 B.n83 10.6151
R813 B.n394 B.n83 10.6151
R814 B.n395 B.n394 10.6151
R815 B.n396 B.n395 10.6151
R816 B.n396 B.n81 10.6151
R817 B.n400 B.n81 10.6151
R818 B.n401 B.n400 10.6151
R819 B.n402 B.n401 10.6151
R820 B.n402 B.n79 10.6151
R821 B.n406 B.n79 10.6151
R822 B.n407 B.n406 10.6151
R823 B.n408 B.n407 10.6151
R824 B.n408 B.n77 10.6151
R825 B.n412 B.n77 10.6151
R826 B.n413 B.n412 10.6151
R827 B.n414 B.n413 10.6151
R828 B.n414 B.n75 10.6151
R829 B.n418 B.n75 10.6151
R830 B.n419 B.n418 10.6151
R831 B.n420 B.n419 10.6151
R832 B.n420 B.n73 10.6151
R833 B.n424 B.n73 10.6151
R834 B.n425 B.n424 10.6151
R835 B.n426 B.n425 10.6151
R836 B.n426 B.n71 10.6151
R837 B.n430 B.n71 10.6151
R838 B.n431 B.n430 10.6151
R839 B.n432 B.n431 10.6151
R840 B.n432 B.n69 10.6151
R841 B.n436 B.n69 10.6151
R842 B.n437 B.n436 10.6151
R843 B.n438 B.n437 10.6151
R844 B.n438 B.n67 10.6151
R845 B.n442 B.n67 10.6151
R846 B.n443 B.n442 10.6151
R847 B.n444 B.n443 10.6151
R848 B.n444 B.n65 10.6151
R849 B.n448 B.n65 10.6151
R850 B.n220 B.n145 10.6151
R851 B.n221 B.n220 10.6151
R852 B.n222 B.n221 10.6151
R853 B.n222 B.n143 10.6151
R854 B.n226 B.n143 10.6151
R855 B.n227 B.n226 10.6151
R856 B.n228 B.n227 10.6151
R857 B.n228 B.n141 10.6151
R858 B.n232 B.n141 10.6151
R859 B.n233 B.n232 10.6151
R860 B.n234 B.n233 10.6151
R861 B.n234 B.n139 10.6151
R862 B.n238 B.n139 10.6151
R863 B.n239 B.n238 10.6151
R864 B.n240 B.n239 10.6151
R865 B.n240 B.n137 10.6151
R866 B.n244 B.n137 10.6151
R867 B.n245 B.n244 10.6151
R868 B.n246 B.n245 10.6151
R869 B.n246 B.n135 10.6151
R870 B.n250 B.n135 10.6151
R871 B.n251 B.n250 10.6151
R872 B.n252 B.n251 10.6151
R873 B.n252 B.n133 10.6151
R874 B.n256 B.n133 10.6151
R875 B.n257 B.n256 10.6151
R876 B.n258 B.n257 10.6151
R877 B.n258 B.n131 10.6151
R878 B.n262 B.n131 10.6151
R879 B.n263 B.n262 10.6151
R880 B.n264 B.n263 10.6151
R881 B.n264 B.n129 10.6151
R882 B.n268 B.n129 10.6151
R883 B.n271 B.n270 10.6151
R884 B.n271 B.n125 10.6151
R885 B.n275 B.n125 10.6151
R886 B.n276 B.n275 10.6151
R887 B.n277 B.n276 10.6151
R888 B.n277 B.n123 10.6151
R889 B.n281 B.n123 10.6151
R890 B.n282 B.n281 10.6151
R891 B.n283 B.n282 10.6151
R892 B.n287 B.n286 10.6151
R893 B.n288 B.n287 10.6151
R894 B.n288 B.n117 10.6151
R895 B.n292 B.n117 10.6151
R896 B.n293 B.n292 10.6151
R897 B.n294 B.n293 10.6151
R898 B.n294 B.n115 10.6151
R899 B.n298 B.n115 10.6151
R900 B.n299 B.n298 10.6151
R901 B.n300 B.n299 10.6151
R902 B.n300 B.n113 10.6151
R903 B.n304 B.n113 10.6151
R904 B.n305 B.n304 10.6151
R905 B.n306 B.n305 10.6151
R906 B.n306 B.n111 10.6151
R907 B.n310 B.n111 10.6151
R908 B.n311 B.n310 10.6151
R909 B.n312 B.n311 10.6151
R910 B.n312 B.n109 10.6151
R911 B.n316 B.n109 10.6151
R912 B.n317 B.n316 10.6151
R913 B.n318 B.n317 10.6151
R914 B.n318 B.n107 10.6151
R915 B.n322 B.n107 10.6151
R916 B.n323 B.n322 10.6151
R917 B.n324 B.n323 10.6151
R918 B.n324 B.n105 10.6151
R919 B.n328 B.n105 10.6151
R920 B.n329 B.n328 10.6151
R921 B.n330 B.n329 10.6151
R922 B.n330 B.n103 10.6151
R923 B.n334 B.n103 10.6151
R924 B.n335 B.n334 10.6151
R925 B.n216 B.n215 10.6151
R926 B.n215 B.n214 10.6151
R927 B.n214 B.n147 10.6151
R928 B.n210 B.n147 10.6151
R929 B.n210 B.n209 10.6151
R930 B.n209 B.n208 10.6151
R931 B.n208 B.n149 10.6151
R932 B.n204 B.n149 10.6151
R933 B.n204 B.n203 10.6151
R934 B.n203 B.n202 10.6151
R935 B.n202 B.n151 10.6151
R936 B.n198 B.n151 10.6151
R937 B.n198 B.n197 10.6151
R938 B.n197 B.n196 10.6151
R939 B.n196 B.n153 10.6151
R940 B.n192 B.n153 10.6151
R941 B.n192 B.n191 10.6151
R942 B.n191 B.n190 10.6151
R943 B.n190 B.n155 10.6151
R944 B.n186 B.n155 10.6151
R945 B.n186 B.n185 10.6151
R946 B.n185 B.n184 10.6151
R947 B.n184 B.n157 10.6151
R948 B.n180 B.n157 10.6151
R949 B.n180 B.n179 10.6151
R950 B.n179 B.n178 10.6151
R951 B.n178 B.n159 10.6151
R952 B.n174 B.n159 10.6151
R953 B.n174 B.n173 10.6151
R954 B.n173 B.n172 10.6151
R955 B.n172 B.n161 10.6151
R956 B.n168 B.n161 10.6151
R957 B.n168 B.n167 10.6151
R958 B.n167 B.n166 10.6151
R959 B.n166 B.n163 10.6151
R960 B.n163 B.n0 10.6151
R961 B.n619 B.n1 10.6151
R962 B.n619 B.n618 10.6151
R963 B.n618 B.n617 10.6151
R964 B.n617 B.n4 10.6151
R965 B.n613 B.n4 10.6151
R966 B.n613 B.n612 10.6151
R967 B.n612 B.n611 10.6151
R968 B.n611 B.n6 10.6151
R969 B.n607 B.n6 10.6151
R970 B.n607 B.n606 10.6151
R971 B.n606 B.n605 10.6151
R972 B.n605 B.n8 10.6151
R973 B.n601 B.n8 10.6151
R974 B.n601 B.n600 10.6151
R975 B.n600 B.n599 10.6151
R976 B.n599 B.n10 10.6151
R977 B.n595 B.n10 10.6151
R978 B.n595 B.n594 10.6151
R979 B.n594 B.n593 10.6151
R980 B.n593 B.n12 10.6151
R981 B.n589 B.n12 10.6151
R982 B.n589 B.n588 10.6151
R983 B.n588 B.n587 10.6151
R984 B.n587 B.n14 10.6151
R985 B.n583 B.n14 10.6151
R986 B.n583 B.n582 10.6151
R987 B.n582 B.n581 10.6151
R988 B.n581 B.n16 10.6151
R989 B.n577 B.n16 10.6151
R990 B.n577 B.n576 10.6151
R991 B.n576 B.n575 10.6151
R992 B.n575 B.n18 10.6151
R993 B.n571 B.n18 10.6151
R994 B.n571 B.n570 10.6151
R995 B.n570 B.n569 10.6151
R996 B.n569 B.n20 10.6151
R997 B.n516 B.n515 9.36635
R998 B.n498 B.n48 9.36635
R999 B.n269 B.n268 9.36635
R1000 B.n286 B.n121 9.36635
R1001 B.n623 B.n0 2.81026
R1002 B.n623 B.n1 2.81026
R1003 B.n515 B.n514 1.24928
R1004 B.n48 B.n44 1.24928
R1005 B.n270 B.n269 1.24928
R1006 B.n283 B.n121 1.24928
C0 VTAIL VP 4.00607f
C1 VDD1 VP 4.18109f
C2 VDD2 VP 0.415778f
C3 B VP 1.77366f
C4 VP VN 5.97301f
C5 w_n2926_n2876# VP 5.35021f
C6 VDD1 VTAIL 4.91294f
C7 VTAIL VDD2 4.96936f
C8 B VTAIL 4.26799f
C9 VTAIL VN 3.99196f
C10 VDD1 VDD2 1.10531f
C11 w_n2926_n2876# VTAIL 3.43613f
C12 B VDD1 1.25324f
C13 B VDD2 1.31087f
C14 VDD1 VN 0.149772f
C15 VDD2 VN 3.9159f
C16 B VN 1.14653f
C17 VDD1 w_n2926_n2876# 1.45229f
C18 w_n2926_n2876# VDD2 1.51572f
C19 B w_n2926_n2876# 8.961981f
C20 w_n2926_n2876# VN 4.97323f
C21 VDD2 VSUBS 0.943831f
C22 VDD1 VSUBS 5.61401f
C23 VTAIL VSUBS 1.143486f
C24 VN VSUBS 5.588719f
C25 VP VSUBS 2.382771f
C26 B VSUBS 4.353094f
C27 w_n2926_n2876# VSUBS 0.104037p
C28 B.n0 VSUBS 0.004458f
C29 B.n1 VSUBS 0.004458f
C30 B.n2 VSUBS 0.00705f
C31 B.n3 VSUBS 0.00705f
C32 B.n4 VSUBS 0.00705f
C33 B.n5 VSUBS 0.00705f
C34 B.n6 VSUBS 0.00705f
C35 B.n7 VSUBS 0.00705f
C36 B.n8 VSUBS 0.00705f
C37 B.n9 VSUBS 0.00705f
C38 B.n10 VSUBS 0.00705f
C39 B.n11 VSUBS 0.00705f
C40 B.n12 VSUBS 0.00705f
C41 B.n13 VSUBS 0.00705f
C42 B.n14 VSUBS 0.00705f
C43 B.n15 VSUBS 0.00705f
C44 B.n16 VSUBS 0.00705f
C45 B.n17 VSUBS 0.00705f
C46 B.n18 VSUBS 0.00705f
C47 B.n19 VSUBS 0.00705f
C48 B.n20 VSUBS 0.016397f
C49 B.n21 VSUBS 0.00705f
C50 B.n22 VSUBS 0.00705f
C51 B.n23 VSUBS 0.00705f
C52 B.n24 VSUBS 0.00705f
C53 B.n25 VSUBS 0.00705f
C54 B.n26 VSUBS 0.00705f
C55 B.n27 VSUBS 0.00705f
C56 B.n28 VSUBS 0.00705f
C57 B.n29 VSUBS 0.00705f
C58 B.n30 VSUBS 0.00705f
C59 B.n31 VSUBS 0.00705f
C60 B.n32 VSUBS 0.00705f
C61 B.n33 VSUBS 0.00705f
C62 B.n34 VSUBS 0.00705f
C63 B.n35 VSUBS 0.00705f
C64 B.n36 VSUBS 0.00705f
C65 B.n37 VSUBS 0.00705f
C66 B.t11 VSUBS 0.304496f
C67 B.t10 VSUBS 0.327881f
C68 B.t9 VSUBS 1.30929f
C69 B.n38 VSUBS 0.1771f
C70 B.n39 VSUBS 0.073468f
C71 B.n40 VSUBS 0.00705f
C72 B.n41 VSUBS 0.00705f
C73 B.n42 VSUBS 0.00705f
C74 B.n43 VSUBS 0.00705f
C75 B.n44 VSUBS 0.00394f
C76 B.n45 VSUBS 0.00705f
C77 B.t5 VSUBS 0.304492f
C78 B.t4 VSUBS 0.327877f
C79 B.t3 VSUBS 1.30929f
C80 B.n46 VSUBS 0.177104f
C81 B.n47 VSUBS 0.073472f
C82 B.n48 VSUBS 0.016334f
C83 B.n49 VSUBS 0.00705f
C84 B.n50 VSUBS 0.00705f
C85 B.n51 VSUBS 0.00705f
C86 B.n52 VSUBS 0.00705f
C87 B.n53 VSUBS 0.00705f
C88 B.n54 VSUBS 0.00705f
C89 B.n55 VSUBS 0.00705f
C90 B.n56 VSUBS 0.00705f
C91 B.n57 VSUBS 0.00705f
C92 B.n58 VSUBS 0.00705f
C93 B.n59 VSUBS 0.00705f
C94 B.n60 VSUBS 0.00705f
C95 B.n61 VSUBS 0.00705f
C96 B.n62 VSUBS 0.00705f
C97 B.n63 VSUBS 0.00705f
C98 B.n64 VSUBS 0.01678f
C99 B.n65 VSUBS 0.00705f
C100 B.n66 VSUBS 0.00705f
C101 B.n67 VSUBS 0.00705f
C102 B.n68 VSUBS 0.00705f
C103 B.n69 VSUBS 0.00705f
C104 B.n70 VSUBS 0.00705f
C105 B.n71 VSUBS 0.00705f
C106 B.n72 VSUBS 0.00705f
C107 B.n73 VSUBS 0.00705f
C108 B.n74 VSUBS 0.00705f
C109 B.n75 VSUBS 0.00705f
C110 B.n76 VSUBS 0.00705f
C111 B.n77 VSUBS 0.00705f
C112 B.n78 VSUBS 0.00705f
C113 B.n79 VSUBS 0.00705f
C114 B.n80 VSUBS 0.00705f
C115 B.n81 VSUBS 0.00705f
C116 B.n82 VSUBS 0.00705f
C117 B.n83 VSUBS 0.00705f
C118 B.n84 VSUBS 0.00705f
C119 B.n85 VSUBS 0.00705f
C120 B.n86 VSUBS 0.00705f
C121 B.n87 VSUBS 0.00705f
C122 B.n88 VSUBS 0.00705f
C123 B.n89 VSUBS 0.00705f
C124 B.n90 VSUBS 0.00705f
C125 B.n91 VSUBS 0.00705f
C126 B.n92 VSUBS 0.00705f
C127 B.n93 VSUBS 0.00705f
C128 B.n94 VSUBS 0.00705f
C129 B.n95 VSUBS 0.00705f
C130 B.n96 VSUBS 0.00705f
C131 B.n97 VSUBS 0.00705f
C132 B.n98 VSUBS 0.00705f
C133 B.n99 VSUBS 0.00705f
C134 B.n100 VSUBS 0.00705f
C135 B.n101 VSUBS 0.00705f
C136 B.n102 VSUBS 0.01678f
C137 B.n103 VSUBS 0.00705f
C138 B.n104 VSUBS 0.00705f
C139 B.n105 VSUBS 0.00705f
C140 B.n106 VSUBS 0.00705f
C141 B.n107 VSUBS 0.00705f
C142 B.n108 VSUBS 0.00705f
C143 B.n109 VSUBS 0.00705f
C144 B.n110 VSUBS 0.00705f
C145 B.n111 VSUBS 0.00705f
C146 B.n112 VSUBS 0.00705f
C147 B.n113 VSUBS 0.00705f
C148 B.n114 VSUBS 0.00705f
C149 B.n115 VSUBS 0.00705f
C150 B.n116 VSUBS 0.00705f
C151 B.n117 VSUBS 0.00705f
C152 B.n118 VSUBS 0.00705f
C153 B.t7 VSUBS 0.304492f
C154 B.t8 VSUBS 0.327877f
C155 B.t6 VSUBS 1.30929f
C156 B.n119 VSUBS 0.177104f
C157 B.n120 VSUBS 0.073472f
C158 B.n121 VSUBS 0.016334f
C159 B.n122 VSUBS 0.00705f
C160 B.n123 VSUBS 0.00705f
C161 B.n124 VSUBS 0.00705f
C162 B.n125 VSUBS 0.00705f
C163 B.n126 VSUBS 0.00705f
C164 B.t1 VSUBS 0.304496f
C165 B.t2 VSUBS 0.327881f
C166 B.t0 VSUBS 1.30929f
C167 B.n127 VSUBS 0.1771f
C168 B.n128 VSUBS 0.073468f
C169 B.n129 VSUBS 0.00705f
C170 B.n130 VSUBS 0.00705f
C171 B.n131 VSUBS 0.00705f
C172 B.n132 VSUBS 0.00705f
C173 B.n133 VSUBS 0.00705f
C174 B.n134 VSUBS 0.00705f
C175 B.n135 VSUBS 0.00705f
C176 B.n136 VSUBS 0.00705f
C177 B.n137 VSUBS 0.00705f
C178 B.n138 VSUBS 0.00705f
C179 B.n139 VSUBS 0.00705f
C180 B.n140 VSUBS 0.00705f
C181 B.n141 VSUBS 0.00705f
C182 B.n142 VSUBS 0.00705f
C183 B.n143 VSUBS 0.00705f
C184 B.n144 VSUBS 0.00705f
C185 B.n145 VSUBS 0.01678f
C186 B.n146 VSUBS 0.00705f
C187 B.n147 VSUBS 0.00705f
C188 B.n148 VSUBS 0.00705f
C189 B.n149 VSUBS 0.00705f
C190 B.n150 VSUBS 0.00705f
C191 B.n151 VSUBS 0.00705f
C192 B.n152 VSUBS 0.00705f
C193 B.n153 VSUBS 0.00705f
C194 B.n154 VSUBS 0.00705f
C195 B.n155 VSUBS 0.00705f
C196 B.n156 VSUBS 0.00705f
C197 B.n157 VSUBS 0.00705f
C198 B.n158 VSUBS 0.00705f
C199 B.n159 VSUBS 0.00705f
C200 B.n160 VSUBS 0.00705f
C201 B.n161 VSUBS 0.00705f
C202 B.n162 VSUBS 0.00705f
C203 B.n163 VSUBS 0.00705f
C204 B.n164 VSUBS 0.00705f
C205 B.n165 VSUBS 0.00705f
C206 B.n166 VSUBS 0.00705f
C207 B.n167 VSUBS 0.00705f
C208 B.n168 VSUBS 0.00705f
C209 B.n169 VSUBS 0.00705f
C210 B.n170 VSUBS 0.00705f
C211 B.n171 VSUBS 0.00705f
C212 B.n172 VSUBS 0.00705f
C213 B.n173 VSUBS 0.00705f
C214 B.n174 VSUBS 0.00705f
C215 B.n175 VSUBS 0.00705f
C216 B.n176 VSUBS 0.00705f
C217 B.n177 VSUBS 0.00705f
C218 B.n178 VSUBS 0.00705f
C219 B.n179 VSUBS 0.00705f
C220 B.n180 VSUBS 0.00705f
C221 B.n181 VSUBS 0.00705f
C222 B.n182 VSUBS 0.00705f
C223 B.n183 VSUBS 0.00705f
C224 B.n184 VSUBS 0.00705f
C225 B.n185 VSUBS 0.00705f
C226 B.n186 VSUBS 0.00705f
C227 B.n187 VSUBS 0.00705f
C228 B.n188 VSUBS 0.00705f
C229 B.n189 VSUBS 0.00705f
C230 B.n190 VSUBS 0.00705f
C231 B.n191 VSUBS 0.00705f
C232 B.n192 VSUBS 0.00705f
C233 B.n193 VSUBS 0.00705f
C234 B.n194 VSUBS 0.00705f
C235 B.n195 VSUBS 0.00705f
C236 B.n196 VSUBS 0.00705f
C237 B.n197 VSUBS 0.00705f
C238 B.n198 VSUBS 0.00705f
C239 B.n199 VSUBS 0.00705f
C240 B.n200 VSUBS 0.00705f
C241 B.n201 VSUBS 0.00705f
C242 B.n202 VSUBS 0.00705f
C243 B.n203 VSUBS 0.00705f
C244 B.n204 VSUBS 0.00705f
C245 B.n205 VSUBS 0.00705f
C246 B.n206 VSUBS 0.00705f
C247 B.n207 VSUBS 0.00705f
C248 B.n208 VSUBS 0.00705f
C249 B.n209 VSUBS 0.00705f
C250 B.n210 VSUBS 0.00705f
C251 B.n211 VSUBS 0.00705f
C252 B.n212 VSUBS 0.00705f
C253 B.n213 VSUBS 0.00705f
C254 B.n214 VSUBS 0.00705f
C255 B.n215 VSUBS 0.00705f
C256 B.n216 VSUBS 0.016397f
C257 B.n217 VSUBS 0.016397f
C258 B.n218 VSUBS 0.01678f
C259 B.n219 VSUBS 0.00705f
C260 B.n220 VSUBS 0.00705f
C261 B.n221 VSUBS 0.00705f
C262 B.n222 VSUBS 0.00705f
C263 B.n223 VSUBS 0.00705f
C264 B.n224 VSUBS 0.00705f
C265 B.n225 VSUBS 0.00705f
C266 B.n226 VSUBS 0.00705f
C267 B.n227 VSUBS 0.00705f
C268 B.n228 VSUBS 0.00705f
C269 B.n229 VSUBS 0.00705f
C270 B.n230 VSUBS 0.00705f
C271 B.n231 VSUBS 0.00705f
C272 B.n232 VSUBS 0.00705f
C273 B.n233 VSUBS 0.00705f
C274 B.n234 VSUBS 0.00705f
C275 B.n235 VSUBS 0.00705f
C276 B.n236 VSUBS 0.00705f
C277 B.n237 VSUBS 0.00705f
C278 B.n238 VSUBS 0.00705f
C279 B.n239 VSUBS 0.00705f
C280 B.n240 VSUBS 0.00705f
C281 B.n241 VSUBS 0.00705f
C282 B.n242 VSUBS 0.00705f
C283 B.n243 VSUBS 0.00705f
C284 B.n244 VSUBS 0.00705f
C285 B.n245 VSUBS 0.00705f
C286 B.n246 VSUBS 0.00705f
C287 B.n247 VSUBS 0.00705f
C288 B.n248 VSUBS 0.00705f
C289 B.n249 VSUBS 0.00705f
C290 B.n250 VSUBS 0.00705f
C291 B.n251 VSUBS 0.00705f
C292 B.n252 VSUBS 0.00705f
C293 B.n253 VSUBS 0.00705f
C294 B.n254 VSUBS 0.00705f
C295 B.n255 VSUBS 0.00705f
C296 B.n256 VSUBS 0.00705f
C297 B.n257 VSUBS 0.00705f
C298 B.n258 VSUBS 0.00705f
C299 B.n259 VSUBS 0.00705f
C300 B.n260 VSUBS 0.00705f
C301 B.n261 VSUBS 0.00705f
C302 B.n262 VSUBS 0.00705f
C303 B.n263 VSUBS 0.00705f
C304 B.n264 VSUBS 0.00705f
C305 B.n265 VSUBS 0.00705f
C306 B.n266 VSUBS 0.00705f
C307 B.n267 VSUBS 0.00705f
C308 B.n268 VSUBS 0.006635f
C309 B.n269 VSUBS 0.016334f
C310 B.n270 VSUBS 0.00394f
C311 B.n271 VSUBS 0.00705f
C312 B.n272 VSUBS 0.00705f
C313 B.n273 VSUBS 0.00705f
C314 B.n274 VSUBS 0.00705f
C315 B.n275 VSUBS 0.00705f
C316 B.n276 VSUBS 0.00705f
C317 B.n277 VSUBS 0.00705f
C318 B.n278 VSUBS 0.00705f
C319 B.n279 VSUBS 0.00705f
C320 B.n280 VSUBS 0.00705f
C321 B.n281 VSUBS 0.00705f
C322 B.n282 VSUBS 0.00705f
C323 B.n283 VSUBS 0.00394f
C324 B.n284 VSUBS 0.00705f
C325 B.n285 VSUBS 0.00705f
C326 B.n286 VSUBS 0.006635f
C327 B.n287 VSUBS 0.00705f
C328 B.n288 VSUBS 0.00705f
C329 B.n289 VSUBS 0.00705f
C330 B.n290 VSUBS 0.00705f
C331 B.n291 VSUBS 0.00705f
C332 B.n292 VSUBS 0.00705f
C333 B.n293 VSUBS 0.00705f
C334 B.n294 VSUBS 0.00705f
C335 B.n295 VSUBS 0.00705f
C336 B.n296 VSUBS 0.00705f
C337 B.n297 VSUBS 0.00705f
C338 B.n298 VSUBS 0.00705f
C339 B.n299 VSUBS 0.00705f
C340 B.n300 VSUBS 0.00705f
C341 B.n301 VSUBS 0.00705f
C342 B.n302 VSUBS 0.00705f
C343 B.n303 VSUBS 0.00705f
C344 B.n304 VSUBS 0.00705f
C345 B.n305 VSUBS 0.00705f
C346 B.n306 VSUBS 0.00705f
C347 B.n307 VSUBS 0.00705f
C348 B.n308 VSUBS 0.00705f
C349 B.n309 VSUBS 0.00705f
C350 B.n310 VSUBS 0.00705f
C351 B.n311 VSUBS 0.00705f
C352 B.n312 VSUBS 0.00705f
C353 B.n313 VSUBS 0.00705f
C354 B.n314 VSUBS 0.00705f
C355 B.n315 VSUBS 0.00705f
C356 B.n316 VSUBS 0.00705f
C357 B.n317 VSUBS 0.00705f
C358 B.n318 VSUBS 0.00705f
C359 B.n319 VSUBS 0.00705f
C360 B.n320 VSUBS 0.00705f
C361 B.n321 VSUBS 0.00705f
C362 B.n322 VSUBS 0.00705f
C363 B.n323 VSUBS 0.00705f
C364 B.n324 VSUBS 0.00705f
C365 B.n325 VSUBS 0.00705f
C366 B.n326 VSUBS 0.00705f
C367 B.n327 VSUBS 0.00705f
C368 B.n328 VSUBS 0.00705f
C369 B.n329 VSUBS 0.00705f
C370 B.n330 VSUBS 0.00705f
C371 B.n331 VSUBS 0.00705f
C372 B.n332 VSUBS 0.00705f
C373 B.n333 VSUBS 0.00705f
C374 B.n334 VSUBS 0.00705f
C375 B.n335 VSUBS 0.01678f
C376 B.n336 VSUBS 0.016397f
C377 B.n337 VSUBS 0.016397f
C378 B.n338 VSUBS 0.00705f
C379 B.n339 VSUBS 0.00705f
C380 B.n340 VSUBS 0.00705f
C381 B.n341 VSUBS 0.00705f
C382 B.n342 VSUBS 0.00705f
C383 B.n343 VSUBS 0.00705f
C384 B.n344 VSUBS 0.00705f
C385 B.n345 VSUBS 0.00705f
C386 B.n346 VSUBS 0.00705f
C387 B.n347 VSUBS 0.00705f
C388 B.n348 VSUBS 0.00705f
C389 B.n349 VSUBS 0.00705f
C390 B.n350 VSUBS 0.00705f
C391 B.n351 VSUBS 0.00705f
C392 B.n352 VSUBS 0.00705f
C393 B.n353 VSUBS 0.00705f
C394 B.n354 VSUBS 0.00705f
C395 B.n355 VSUBS 0.00705f
C396 B.n356 VSUBS 0.00705f
C397 B.n357 VSUBS 0.00705f
C398 B.n358 VSUBS 0.00705f
C399 B.n359 VSUBS 0.00705f
C400 B.n360 VSUBS 0.00705f
C401 B.n361 VSUBS 0.00705f
C402 B.n362 VSUBS 0.00705f
C403 B.n363 VSUBS 0.00705f
C404 B.n364 VSUBS 0.00705f
C405 B.n365 VSUBS 0.00705f
C406 B.n366 VSUBS 0.00705f
C407 B.n367 VSUBS 0.00705f
C408 B.n368 VSUBS 0.00705f
C409 B.n369 VSUBS 0.00705f
C410 B.n370 VSUBS 0.00705f
C411 B.n371 VSUBS 0.00705f
C412 B.n372 VSUBS 0.00705f
C413 B.n373 VSUBS 0.00705f
C414 B.n374 VSUBS 0.00705f
C415 B.n375 VSUBS 0.00705f
C416 B.n376 VSUBS 0.00705f
C417 B.n377 VSUBS 0.00705f
C418 B.n378 VSUBS 0.00705f
C419 B.n379 VSUBS 0.00705f
C420 B.n380 VSUBS 0.00705f
C421 B.n381 VSUBS 0.00705f
C422 B.n382 VSUBS 0.00705f
C423 B.n383 VSUBS 0.00705f
C424 B.n384 VSUBS 0.00705f
C425 B.n385 VSUBS 0.00705f
C426 B.n386 VSUBS 0.00705f
C427 B.n387 VSUBS 0.00705f
C428 B.n388 VSUBS 0.00705f
C429 B.n389 VSUBS 0.00705f
C430 B.n390 VSUBS 0.00705f
C431 B.n391 VSUBS 0.00705f
C432 B.n392 VSUBS 0.00705f
C433 B.n393 VSUBS 0.00705f
C434 B.n394 VSUBS 0.00705f
C435 B.n395 VSUBS 0.00705f
C436 B.n396 VSUBS 0.00705f
C437 B.n397 VSUBS 0.00705f
C438 B.n398 VSUBS 0.00705f
C439 B.n399 VSUBS 0.00705f
C440 B.n400 VSUBS 0.00705f
C441 B.n401 VSUBS 0.00705f
C442 B.n402 VSUBS 0.00705f
C443 B.n403 VSUBS 0.00705f
C444 B.n404 VSUBS 0.00705f
C445 B.n405 VSUBS 0.00705f
C446 B.n406 VSUBS 0.00705f
C447 B.n407 VSUBS 0.00705f
C448 B.n408 VSUBS 0.00705f
C449 B.n409 VSUBS 0.00705f
C450 B.n410 VSUBS 0.00705f
C451 B.n411 VSUBS 0.00705f
C452 B.n412 VSUBS 0.00705f
C453 B.n413 VSUBS 0.00705f
C454 B.n414 VSUBS 0.00705f
C455 B.n415 VSUBS 0.00705f
C456 B.n416 VSUBS 0.00705f
C457 B.n417 VSUBS 0.00705f
C458 B.n418 VSUBS 0.00705f
C459 B.n419 VSUBS 0.00705f
C460 B.n420 VSUBS 0.00705f
C461 B.n421 VSUBS 0.00705f
C462 B.n422 VSUBS 0.00705f
C463 B.n423 VSUBS 0.00705f
C464 B.n424 VSUBS 0.00705f
C465 B.n425 VSUBS 0.00705f
C466 B.n426 VSUBS 0.00705f
C467 B.n427 VSUBS 0.00705f
C468 B.n428 VSUBS 0.00705f
C469 B.n429 VSUBS 0.00705f
C470 B.n430 VSUBS 0.00705f
C471 B.n431 VSUBS 0.00705f
C472 B.n432 VSUBS 0.00705f
C473 B.n433 VSUBS 0.00705f
C474 B.n434 VSUBS 0.00705f
C475 B.n435 VSUBS 0.00705f
C476 B.n436 VSUBS 0.00705f
C477 B.n437 VSUBS 0.00705f
C478 B.n438 VSUBS 0.00705f
C479 B.n439 VSUBS 0.00705f
C480 B.n440 VSUBS 0.00705f
C481 B.n441 VSUBS 0.00705f
C482 B.n442 VSUBS 0.00705f
C483 B.n443 VSUBS 0.00705f
C484 B.n444 VSUBS 0.00705f
C485 B.n445 VSUBS 0.00705f
C486 B.n446 VSUBS 0.00705f
C487 B.n447 VSUBS 0.016397f
C488 B.n448 VSUBS 0.017223f
C489 B.n449 VSUBS 0.015954f
C490 B.n450 VSUBS 0.00705f
C491 B.n451 VSUBS 0.00705f
C492 B.n452 VSUBS 0.00705f
C493 B.n453 VSUBS 0.00705f
C494 B.n454 VSUBS 0.00705f
C495 B.n455 VSUBS 0.00705f
C496 B.n456 VSUBS 0.00705f
C497 B.n457 VSUBS 0.00705f
C498 B.n458 VSUBS 0.00705f
C499 B.n459 VSUBS 0.00705f
C500 B.n460 VSUBS 0.00705f
C501 B.n461 VSUBS 0.00705f
C502 B.n462 VSUBS 0.00705f
C503 B.n463 VSUBS 0.00705f
C504 B.n464 VSUBS 0.00705f
C505 B.n465 VSUBS 0.00705f
C506 B.n466 VSUBS 0.00705f
C507 B.n467 VSUBS 0.00705f
C508 B.n468 VSUBS 0.00705f
C509 B.n469 VSUBS 0.00705f
C510 B.n470 VSUBS 0.00705f
C511 B.n471 VSUBS 0.00705f
C512 B.n472 VSUBS 0.00705f
C513 B.n473 VSUBS 0.00705f
C514 B.n474 VSUBS 0.00705f
C515 B.n475 VSUBS 0.00705f
C516 B.n476 VSUBS 0.00705f
C517 B.n477 VSUBS 0.00705f
C518 B.n478 VSUBS 0.00705f
C519 B.n479 VSUBS 0.00705f
C520 B.n480 VSUBS 0.00705f
C521 B.n481 VSUBS 0.00705f
C522 B.n482 VSUBS 0.00705f
C523 B.n483 VSUBS 0.00705f
C524 B.n484 VSUBS 0.00705f
C525 B.n485 VSUBS 0.00705f
C526 B.n486 VSUBS 0.00705f
C527 B.n487 VSUBS 0.00705f
C528 B.n488 VSUBS 0.00705f
C529 B.n489 VSUBS 0.00705f
C530 B.n490 VSUBS 0.00705f
C531 B.n491 VSUBS 0.00705f
C532 B.n492 VSUBS 0.00705f
C533 B.n493 VSUBS 0.00705f
C534 B.n494 VSUBS 0.00705f
C535 B.n495 VSUBS 0.00705f
C536 B.n496 VSUBS 0.00705f
C537 B.n497 VSUBS 0.00705f
C538 B.n498 VSUBS 0.006635f
C539 B.n499 VSUBS 0.00705f
C540 B.n500 VSUBS 0.00705f
C541 B.n501 VSUBS 0.00705f
C542 B.n502 VSUBS 0.00705f
C543 B.n503 VSUBS 0.00705f
C544 B.n504 VSUBS 0.00705f
C545 B.n505 VSUBS 0.00705f
C546 B.n506 VSUBS 0.00705f
C547 B.n507 VSUBS 0.00705f
C548 B.n508 VSUBS 0.00705f
C549 B.n509 VSUBS 0.00705f
C550 B.n510 VSUBS 0.00705f
C551 B.n511 VSUBS 0.00705f
C552 B.n512 VSUBS 0.00705f
C553 B.n513 VSUBS 0.00705f
C554 B.n514 VSUBS 0.00394f
C555 B.n515 VSUBS 0.016334f
C556 B.n516 VSUBS 0.006635f
C557 B.n517 VSUBS 0.00705f
C558 B.n518 VSUBS 0.00705f
C559 B.n519 VSUBS 0.00705f
C560 B.n520 VSUBS 0.00705f
C561 B.n521 VSUBS 0.00705f
C562 B.n522 VSUBS 0.00705f
C563 B.n523 VSUBS 0.00705f
C564 B.n524 VSUBS 0.00705f
C565 B.n525 VSUBS 0.00705f
C566 B.n526 VSUBS 0.00705f
C567 B.n527 VSUBS 0.00705f
C568 B.n528 VSUBS 0.00705f
C569 B.n529 VSUBS 0.00705f
C570 B.n530 VSUBS 0.00705f
C571 B.n531 VSUBS 0.00705f
C572 B.n532 VSUBS 0.00705f
C573 B.n533 VSUBS 0.00705f
C574 B.n534 VSUBS 0.00705f
C575 B.n535 VSUBS 0.00705f
C576 B.n536 VSUBS 0.00705f
C577 B.n537 VSUBS 0.00705f
C578 B.n538 VSUBS 0.00705f
C579 B.n539 VSUBS 0.00705f
C580 B.n540 VSUBS 0.00705f
C581 B.n541 VSUBS 0.00705f
C582 B.n542 VSUBS 0.00705f
C583 B.n543 VSUBS 0.00705f
C584 B.n544 VSUBS 0.00705f
C585 B.n545 VSUBS 0.00705f
C586 B.n546 VSUBS 0.00705f
C587 B.n547 VSUBS 0.00705f
C588 B.n548 VSUBS 0.00705f
C589 B.n549 VSUBS 0.00705f
C590 B.n550 VSUBS 0.00705f
C591 B.n551 VSUBS 0.00705f
C592 B.n552 VSUBS 0.00705f
C593 B.n553 VSUBS 0.00705f
C594 B.n554 VSUBS 0.00705f
C595 B.n555 VSUBS 0.00705f
C596 B.n556 VSUBS 0.00705f
C597 B.n557 VSUBS 0.00705f
C598 B.n558 VSUBS 0.00705f
C599 B.n559 VSUBS 0.00705f
C600 B.n560 VSUBS 0.00705f
C601 B.n561 VSUBS 0.00705f
C602 B.n562 VSUBS 0.00705f
C603 B.n563 VSUBS 0.00705f
C604 B.n564 VSUBS 0.00705f
C605 B.n565 VSUBS 0.01678f
C606 B.n566 VSUBS 0.01678f
C607 B.n567 VSUBS 0.016397f
C608 B.n568 VSUBS 0.00705f
C609 B.n569 VSUBS 0.00705f
C610 B.n570 VSUBS 0.00705f
C611 B.n571 VSUBS 0.00705f
C612 B.n572 VSUBS 0.00705f
C613 B.n573 VSUBS 0.00705f
C614 B.n574 VSUBS 0.00705f
C615 B.n575 VSUBS 0.00705f
C616 B.n576 VSUBS 0.00705f
C617 B.n577 VSUBS 0.00705f
C618 B.n578 VSUBS 0.00705f
C619 B.n579 VSUBS 0.00705f
C620 B.n580 VSUBS 0.00705f
C621 B.n581 VSUBS 0.00705f
C622 B.n582 VSUBS 0.00705f
C623 B.n583 VSUBS 0.00705f
C624 B.n584 VSUBS 0.00705f
C625 B.n585 VSUBS 0.00705f
C626 B.n586 VSUBS 0.00705f
C627 B.n587 VSUBS 0.00705f
C628 B.n588 VSUBS 0.00705f
C629 B.n589 VSUBS 0.00705f
C630 B.n590 VSUBS 0.00705f
C631 B.n591 VSUBS 0.00705f
C632 B.n592 VSUBS 0.00705f
C633 B.n593 VSUBS 0.00705f
C634 B.n594 VSUBS 0.00705f
C635 B.n595 VSUBS 0.00705f
C636 B.n596 VSUBS 0.00705f
C637 B.n597 VSUBS 0.00705f
C638 B.n598 VSUBS 0.00705f
C639 B.n599 VSUBS 0.00705f
C640 B.n600 VSUBS 0.00705f
C641 B.n601 VSUBS 0.00705f
C642 B.n602 VSUBS 0.00705f
C643 B.n603 VSUBS 0.00705f
C644 B.n604 VSUBS 0.00705f
C645 B.n605 VSUBS 0.00705f
C646 B.n606 VSUBS 0.00705f
C647 B.n607 VSUBS 0.00705f
C648 B.n608 VSUBS 0.00705f
C649 B.n609 VSUBS 0.00705f
C650 B.n610 VSUBS 0.00705f
C651 B.n611 VSUBS 0.00705f
C652 B.n612 VSUBS 0.00705f
C653 B.n613 VSUBS 0.00705f
C654 B.n614 VSUBS 0.00705f
C655 B.n615 VSUBS 0.00705f
C656 B.n616 VSUBS 0.00705f
C657 B.n617 VSUBS 0.00705f
C658 B.n618 VSUBS 0.00705f
C659 B.n619 VSUBS 0.00705f
C660 B.n620 VSUBS 0.00705f
C661 B.n621 VSUBS 0.00705f
C662 B.n622 VSUBS 0.00705f
C663 B.n623 VSUBS 0.015964f
C664 VDD1.t3 VSUBS 0.207675f
C665 VDD1.t2 VSUBS 0.207675f
C666 VDD1.n0 VSUBS 1.55043f
C667 VDD1.t1 VSUBS 0.207675f
C668 VDD1.t0 VSUBS 0.207675f
C669 VDD1.n1 VSUBS 2.20932f
C670 VP.t3 VSUBS 2.61105f
C671 VP.n0 VSUBS 1.06306f
C672 VP.n1 VSUBS 0.034539f
C673 VP.n2 VSUBS 0.050207f
C674 VP.n3 VSUBS 0.055736f
C675 VP.t2 VSUBS 2.61105f
C676 VP.t0 VSUBS 2.96843f
C677 VP.t1 VSUBS 2.95852f
C678 VP.n4 VSUBS 3.73837f
C679 VP.n5 VSUBS 1.8584f
C680 VP.n6 VSUBS 1.06306f
C681 VP.n7 VSUBS 0.05646f
C682 VP.n8 VSUBS 0.064048f
C683 VP.n9 VSUBS 0.034539f
C684 VP.n10 VSUBS 0.034539f
C685 VP.n11 VSUBS 0.034539f
C686 VP.n12 VSUBS 0.050207f
C687 VP.n13 VSUBS 0.064048f
C688 VP.n14 VSUBS 0.05646f
C689 VP.n15 VSUBS 0.055736f
C690 VP.n16 VSUBS 0.073111f
C691 VDD2.t1 VSUBS 0.205408f
C692 VDD2.t3 VSUBS 0.205408f
C693 VDD2.n0 VSUBS 2.16098f
C694 VDD2.t0 VSUBS 0.205408f
C695 VDD2.t2 VSUBS 0.205408f
C696 VDD2.n1 VSUBS 1.53293f
C697 VDD2.n2 VSUBS 4.13186f
C698 VTAIL.t6 VSUBS 1.71202f
C699 VTAIL.n0 VSUBS 0.783387f
C700 VTAIL.t2 VSUBS 1.71202f
C701 VTAIL.n1 VSUBS 0.892012f
C702 VTAIL.t1 VSUBS 1.71202f
C703 VTAIL.n2 VSUBS 2.08395f
C704 VTAIL.t4 VSUBS 1.71203f
C705 VTAIL.n3 VSUBS 2.08393f
C706 VTAIL.t5 VSUBS 1.71203f
C707 VTAIL.n4 VSUBS 0.891999f
C708 VTAIL.t0 VSUBS 1.71203f
C709 VTAIL.n5 VSUBS 0.891999f
C710 VTAIL.t3 VSUBS 1.71202f
C711 VTAIL.n6 VSUBS 2.08395f
C712 VTAIL.t7 VSUBS 1.71202f
C713 VTAIL.n7 VSUBS 1.96594f
C714 VN.t0 VSUBS 2.84581f
C715 VN.t2 VSUBS 2.85534f
C716 VN.n0 VSUBS 1.76808f
C717 VN.t1 VSUBS 2.85534f
C718 VN.t3 VSUBS 2.84581f
C719 VN.n1 VSUBS 3.60955f
.ends

