* NGSPICE file created from diff_pair_sample_1492.ext - technology: sky130A

.subckt diff_pair_sample_1492 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t19 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=3.8688 ps=20.62 w=9.92 l=3.47
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=3.8688 ps=20.62 w=9.92 l=3.47
X2 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=1.6368 ps=10.25 w=9.92 l=3.47
X3 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=0 ps=0 w=9.92 l=3.47
X4 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=1.6368 ps=10.25 w=9.92 l=3.47
X5 VDD1.t4 VP.t1 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=1.6368 ps=10.25 w=9.92 l=3.47
X6 VDD1.t3 VP.t2 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=3.8688 ps=20.62 w=9.92 l=3.47
X7 VDD1.t2 VP.t3 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=1.6368 ps=10.25 w=9.92 l=3.47
X8 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=0 ps=0 w=9.92 l=3.47
X9 VTAIL.t8 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=1.6368 ps=10.25 w=9.92 l=3.47
X10 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=3.8688 ps=20.62 w=9.92 l=3.47
X11 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=0 ps=0 w=9.92 l=3.47
X12 VTAIL.t7 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=1.6368 ps=10.25 w=9.92 l=3.47
X13 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=1.6368 ps=10.25 w=9.92 l=3.47
X14 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6368 pd=10.25 as=1.6368 ps=10.25 w=9.92 l=3.47
X15 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=3.8688 pd=20.62 as=0 ps=0 w=9.92 l=3.47
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n50 VP.n49 161.3
R8 VP.n48 VP.n1 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n2 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n42 VP.n3 161.3
R13 VP.n41 VP.n40 161.3
R14 VP.n39 VP.n4 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n14 VP.t3 103.058
R23 VP.n27 VP.n8 75.4905
R24 VP.n51 VP.n0 75.4905
R25 VP.n26 VP.n9 75.4905
R26 VP.n4 VP.t4 68.8973
R27 VP.n8 VP.t1 68.8973
R28 VP.n0 VP.t2 68.8973
R29 VP.n13 VP.t5 68.8973
R30 VP.n9 VP.t0 68.8973
R31 VP.n27 VP.n26 50.6662
R32 VP.n14 VP.n13 50.305
R33 VP.n35 VP.n6 50.2647
R34 VP.n43 VP.n2 50.2647
R35 VP.n18 VP.n11 50.2647
R36 VP.n31 VP.n6 30.8893
R37 VP.n47 VP.n2 30.8893
R38 VP.n22 VP.n11 30.8893
R39 VP.n30 VP.n29 24.5923
R40 VP.n31 VP.n30 24.5923
R41 VP.n36 VP.n35 24.5923
R42 VP.n37 VP.n36 24.5923
R43 VP.n37 VP.n4 24.5923
R44 VP.n41 VP.n4 24.5923
R45 VP.n42 VP.n41 24.5923
R46 VP.n43 VP.n42 24.5923
R47 VP.n48 VP.n47 24.5923
R48 VP.n49 VP.n48 24.5923
R49 VP.n23 VP.n22 24.5923
R50 VP.n24 VP.n23 24.5923
R51 VP.n16 VP.n13 24.5923
R52 VP.n17 VP.n16 24.5923
R53 VP.n18 VP.n17 24.5923
R54 VP.n29 VP.n8 14.7556
R55 VP.n49 VP.n0 14.7556
R56 VP.n24 VP.n9 14.7556
R57 VP.n15 VP.n14 2.98131
R58 VP.n26 VP.n25 0.354861
R59 VP.n28 VP.n27 0.354861
R60 VP.n51 VP.n50 0.354861
R61 VP VP.n51 0.267071
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VTAIL.n218 VTAIL.n170 289.615
R83 VTAIL.n50 VTAIL.n2 289.615
R84 VTAIL.n164 VTAIL.n116 289.615
R85 VTAIL.n108 VTAIL.n60 289.615
R86 VTAIL.n186 VTAIL.n185 185
R87 VTAIL.n191 VTAIL.n190 185
R88 VTAIL.n193 VTAIL.n192 185
R89 VTAIL.n182 VTAIL.n181 185
R90 VTAIL.n199 VTAIL.n198 185
R91 VTAIL.n201 VTAIL.n200 185
R92 VTAIL.n178 VTAIL.n177 185
R93 VTAIL.n208 VTAIL.n207 185
R94 VTAIL.n209 VTAIL.n176 185
R95 VTAIL.n211 VTAIL.n210 185
R96 VTAIL.n174 VTAIL.n173 185
R97 VTAIL.n217 VTAIL.n216 185
R98 VTAIL.n219 VTAIL.n218 185
R99 VTAIL.n18 VTAIL.n17 185
R100 VTAIL.n23 VTAIL.n22 185
R101 VTAIL.n25 VTAIL.n24 185
R102 VTAIL.n14 VTAIL.n13 185
R103 VTAIL.n31 VTAIL.n30 185
R104 VTAIL.n33 VTAIL.n32 185
R105 VTAIL.n10 VTAIL.n9 185
R106 VTAIL.n40 VTAIL.n39 185
R107 VTAIL.n41 VTAIL.n8 185
R108 VTAIL.n43 VTAIL.n42 185
R109 VTAIL.n6 VTAIL.n5 185
R110 VTAIL.n49 VTAIL.n48 185
R111 VTAIL.n51 VTAIL.n50 185
R112 VTAIL.n165 VTAIL.n164 185
R113 VTAIL.n163 VTAIL.n162 185
R114 VTAIL.n120 VTAIL.n119 185
R115 VTAIL.n157 VTAIL.n156 185
R116 VTAIL.n155 VTAIL.n122 185
R117 VTAIL.n154 VTAIL.n153 185
R118 VTAIL.n125 VTAIL.n123 185
R119 VTAIL.n148 VTAIL.n147 185
R120 VTAIL.n146 VTAIL.n145 185
R121 VTAIL.n129 VTAIL.n128 185
R122 VTAIL.n140 VTAIL.n139 185
R123 VTAIL.n138 VTAIL.n137 185
R124 VTAIL.n133 VTAIL.n132 185
R125 VTAIL.n109 VTAIL.n108 185
R126 VTAIL.n107 VTAIL.n106 185
R127 VTAIL.n64 VTAIL.n63 185
R128 VTAIL.n101 VTAIL.n100 185
R129 VTAIL.n99 VTAIL.n66 185
R130 VTAIL.n98 VTAIL.n97 185
R131 VTAIL.n69 VTAIL.n67 185
R132 VTAIL.n92 VTAIL.n91 185
R133 VTAIL.n90 VTAIL.n89 185
R134 VTAIL.n73 VTAIL.n72 185
R135 VTAIL.n84 VTAIL.n83 185
R136 VTAIL.n82 VTAIL.n81 185
R137 VTAIL.n77 VTAIL.n76 185
R138 VTAIL.n187 VTAIL.t11 149.524
R139 VTAIL.n19 VTAIL.t10 149.524
R140 VTAIL.n134 VTAIL.t9 149.524
R141 VTAIL.n78 VTAIL.t0 149.524
R142 VTAIL.n191 VTAIL.n185 104.615
R143 VTAIL.n192 VTAIL.n191 104.615
R144 VTAIL.n192 VTAIL.n181 104.615
R145 VTAIL.n199 VTAIL.n181 104.615
R146 VTAIL.n200 VTAIL.n199 104.615
R147 VTAIL.n200 VTAIL.n177 104.615
R148 VTAIL.n208 VTAIL.n177 104.615
R149 VTAIL.n209 VTAIL.n208 104.615
R150 VTAIL.n210 VTAIL.n209 104.615
R151 VTAIL.n210 VTAIL.n173 104.615
R152 VTAIL.n217 VTAIL.n173 104.615
R153 VTAIL.n218 VTAIL.n217 104.615
R154 VTAIL.n23 VTAIL.n17 104.615
R155 VTAIL.n24 VTAIL.n23 104.615
R156 VTAIL.n24 VTAIL.n13 104.615
R157 VTAIL.n31 VTAIL.n13 104.615
R158 VTAIL.n32 VTAIL.n31 104.615
R159 VTAIL.n32 VTAIL.n9 104.615
R160 VTAIL.n40 VTAIL.n9 104.615
R161 VTAIL.n41 VTAIL.n40 104.615
R162 VTAIL.n42 VTAIL.n41 104.615
R163 VTAIL.n42 VTAIL.n5 104.615
R164 VTAIL.n49 VTAIL.n5 104.615
R165 VTAIL.n50 VTAIL.n49 104.615
R166 VTAIL.n164 VTAIL.n163 104.615
R167 VTAIL.n163 VTAIL.n119 104.615
R168 VTAIL.n156 VTAIL.n119 104.615
R169 VTAIL.n156 VTAIL.n155 104.615
R170 VTAIL.n155 VTAIL.n154 104.615
R171 VTAIL.n154 VTAIL.n123 104.615
R172 VTAIL.n147 VTAIL.n123 104.615
R173 VTAIL.n147 VTAIL.n146 104.615
R174 VTAIL.n146 VTAIL.n128 104.615
R175 VTAIL.n139 VTAIL.n128 104.615
R176 VTAIL.n139 VTAIL.n138 104.615
R177 VTAIL.n138 VTAIL.n132 104.615
R178 VTAIL.n108 VTAIL.n107 104.615
R179 VTAIL.n107 VTAIL.n63 104.615
R180 VTAIL.n100 VTAIL.n63 104.615
R181 VTAIL.n100 VTAIL.n99 104.615
R182 VTAIL.n99 VTAIL.n98 104.615
R183 VTAIL.n98 VTAIL.n67 104.615
R184 VTAIL.n91 VTAIL.n67 104.615
R185 VTAIL.n91 VTAIL.n90 104.615
R186 VTAIL.n90 VTAIL.n72 104.615
R187 VTAIL.n83 VTAIL.n72 104.615
R188 VTAIL.n83 VTAIL.n82 104.615
R189 VTAIL.n82 VTAIL.n76 104.615
R190 VTAIL.t11 VTAIL.n185 52.3082
R191 VTAIL.t10 VTAIL.n17 52.3082
R192 VTAIL.t9 VTAIL.n132 52.3082
R193 VTAIL.t0 VTAIL.n76 52.3082
R194 VTAIL.n115 VTAIL.n114 45.1858
R195 VTAIL.n59 VTAIL.n58 45.1858
R196 VTAIL.n1 VTAIL.n0 45.1856
R197 VTAIL.n57 VTAIL.n56 45.1856
R198 VTAIL.n223 VTAIL.n222 31.4096
R199 VTAIL.n55 VTAIL.n54 31.4096
R200 VTAIL.n169 VTAIL.n168 31.4096
R201 VTAIL.n113 VTAIL.n112 31.4096
R202 VTAIL.n59 VTAIL.n57 27.4703
R203 VTAIL.n223 VTAIL.n169 24.1945
R204 VTAIL.n211 VTAIL.n176 13.1884
R205 VTAIL.n43 VTAIL.n8 13.1884
R206 VTAIL.n157 VTAIL.n122 13.1884
R207 VTAIL.n101 VTAIL.n66 13.1884
R208 VTAIL.n207 VTAIL.n206 12.8005
R209 VTAIL.n212 VTAIL.n174 12.8005
R210 VTAIL.n39 VTAIL.n38 12.8005
R211 VTAIL.n44 VTAIL.n6 12.8005
R212 VTAIL.n158 VTAIL.n120 12.8005
R213 VTAIL.n153 VTAIL.n124 12.8005
R214 VTAIL.n102 VTAIL.n64 12.8005
R215 VTAIL.n97 VTAIL.n68 12.8005
R216 VTAIL.n205 VTAIL.n178 12.0247
R217 VTAIL.n216 VTAIL.n215 12.0247
R218 VTAIL.n37 VTAIL.n10 12.0247
R219 VTAIL.n48 VTAIL.n47 12.0247
R220 VTAIL.n162 VTAIL.n161 12.0247
R221 VTAIL.n152 VTAIL.n125 12.0247
R222 VTAIL.n106 VTAIL.n105 12.0247
R223 VTAIL.n96 VTAIL.n69 12.0247
R224 VTAIL.n202 VTAIL.n201 11.249
R225 VTAIL.n219 VTAIL.n172 11.249
R226 VTAIL.n34 VTAIL.n33 11.249
R227 VTAIL.n51 VTAIL.n4 11.249
R228 VTAIL.n165 VTAIL.n118 11.249
R229 VTAIL.n149 VTAIL.n148 11.249
R230 VTAIL.n109 VTAIL.n62 11.249
R231 VTAIL.n93 VTAIL.n92 11.249
R232 VTAIL.n198 VTAIL.n180 10.4732
R233 VTAIL.n220 VTAIL.n170 10.4732
R234 VTAIL.n30 VTAIL.n12 10.4732
R235 VTAIL.n52 VTAIL.n2 10.4732
R236 VTAIL.n166 VTAIL.n116 10.4732
R237 VTAIL.n145 VTAIL.n127 10.4732
R238 VTAIL.n110 VTAIL.n60 10.4732
R239 VTAIL.n89 VTAIL.n71 10.4732
R240 VTAIL.n187 VTAIL.n186 10.2747
R241 VTAIL.n19 VTAIL.n18 10.2747
R242 VTAIL.n134 VTAIL.n133 10.2747
R243 VTAIL.n78 VTAIL.n77 10.2747
R244 VTAIL.n197 VTAIL.n182 9.69747
R245 VTAIL.n29 VTAIL.n14 9.69747
R246 VTAIL.n144 VTAIL.n129 9.69747
R247 VTAIL.n88 VTAIL.n73 9.69747
R248 VTAIL.n222 VTAIL.n221 9.45567
R249 VTAIL.n54 VTAIL.n53 9.45567
R250 VTAIL.n168 VTAIL.n167 9.45567
R251 VTAIL.n112 VTAIL.n111 9.45567
R252 VTAIL.n221 VTAIL.n220 9.3005
R253 VTAIL.n172 VTAIL.n171 9.3005
R254 VTAIL.n215 VTAIL.n214 9.3005
R255 VTAIL.n213 VTAIL.n212 9.3005
R256 VTAIL.n189 VTAIL.n188 9.3005
R257 VTAIL.n184 VTAIL.n183 9.3005
R258 VTAIL.n195 VTAIL.n194 9.3005
R259 VTAIL.n197 VTAIL.n196 9.3005
R260 VTAIL.n180 VTAIL.n179 9.3005
R261 VTAIL.n203 VTAIL.n202 9.3005
R262 VTAIL.n205 VTAIL.n204 9.3005
R263 VTAIL.n206 VTAIL.n175 9.3005
R264 VTAIL.n53 VTAIL.n52 9.3005
R265 VTAIL.n4 VTAIL.n3 9.3005
R266 VTAIL.n47 VTAIL.n46 9.3005
R267 VTAIL.n45 VTAIL.n44 9.3005
R268 VTAIL.n21 VTAIL.n20 9.3005
R269 VTAIL.n16 VTAIL.n15 9.3005
R270 VTAIL.n27 VTAIL.n26 9.3005
R271 VTAIL.n29 VTAIL.n28 9.3005
R272 VTAIL.n12 VTAIL.n11 9.3005
R273 VTAIL.n35 VTAIL.n34 9.3005
R274 VTAIL.n37 VTAIL.n36 9.3005
R275 VTAIL.n38 VTAIL.n7 9.3005
R276 VTAIL.n136 VTAIL.n135 9.3005
R277 VTAIL.n131 VTAIL.n130 9.3005
R278 VTAIL.n142 VTAIL.n141 9.3005
R279 VTAIL.n144 VTAIL.n143 9.3005
R280 VTAIL.n127 VTAIL.n126 9.3005
R281 VTAIL.n150 VTAIL.n149 9.3005
R282 VTAIL.n152 VTAIL.n151 9.3005
R283 VTAIL.n124 VTAIL.n121 9.3005
R284 VTAIL.n167 VTAIL.n166 9.3005
R285 VTAIL.n118 VTAIL.n117 9.3005
R286 VTAIL.n161 VTAIL.n160 9.3005
R287 VTAIL.n159 VTAIL.n158 9.3005
R288 VTAIL.n80 VTAIL.n79 9.3005
R289 VTAIL.n75 VTAIL.n74 9.3005
R290 VTAIL.n86 VTAIL.n85 9.3005
R291 VTAIL.n88 VTAIL.n87 9.3005
R292 VTAIL.n71 VTAIL.n70 9.3005
R293 VTAIL.n94 VTAIL.n93 9.3005
R294 VTAIL.n96 VTAIL.n95 9.3005
R295 VTAIL.n68 VTAIL.n65 9.3005
R296 VTAIL.n111 VTAIL.n110 9.3005
R297 VTAIL.n62 VTAIL.n61 9.3005
R298 VTAIL.n105 VTAIL.n104 9.3005
R299 VTAIL.n103 VTAIL.n102 9.3005
R300 VTAIL.n194 VTAIL.n193 8.92171
R301 VTAIL.n26 VTAIL.n25 8.92171
R302 VTAIL.n141 VTAIL.n140 8.92171
R303 VTAIL.n85 VTAIL.n84 8.92171
R304 VTAIL.n190 VTAIL.n184 8.14595
R305 VTAIL.n22 VTAIL.n16 8.14595
R306 VTAIL.n137 VTAIL.n131 8.14595
R307 VTAIL.n81 VTAIL.n75 8.14595
R308 VTAIL.n189 VTAIL.n186 7.3702
R309 VTAIL.n21 VTAIL.n18 7.3702
R310 VTAIL.n136 VTAIL.n133 7.3702
R311 VTAIL.n80 VTAIL.n77 7.3702
R312 VTAIL.n190 VTAIL.n189 5.81868
R313 VTAIL.n22 VTAIL.n21 5.81868
R314 VTAIL.n137 VTAIL.n136 5.81868
R315 VTAIL.n81 VTAIL.n80 5.81868
R316 VTAIL.n193 VTAIL.n184 5.04292
R317 VTAIL.n25 VTAIL.n16 5.04292
R318 VTAIL.n140 VTAIL.n131 5.04292
R319 VTAIL.n84 VTAIL.n75 5.04292
R320 VTAIL.n194 VTAIL.n182 4.26717
R321 VTAIL.n26 VTAIL.n14 4.26717
R322 VTAIL.n141 VTAIL.n129 4.26717
R323 VTAIL.n85 VTAIL.n73 4.26717
R324 VTAIL.n198 VTAIL.n197 3.49141
R325 VTAIL.n222 VTAIL.n170 3.49141
R326 VTAIL.n30 VTAIL.n29 3.49141
R327 VTAIL.n54 VTAIL.n2 3.49141
R328 VTAIL.n168 VTAIL.n116 3.49141
R329 VTAIL.n145 VTAIL.n144 3.49141
R330 VTAIL.n112 VTAIL.n60 3.49141
R331 VTAIL.n89 VTAIL.n88 3.49141
R332 VTAIL.n113 VTAIL.n59 3.27636
R333 VTAIL.n169 VTAIL.n115 3.27636
R334 VTAIL.n57 VTAIL.n55 3.27636
R335 VTAIL.n188 VTAIL.n187 2.84303
R336 VTAIL.n20 VTAIL.n19 2.84303
R337 VTAIL.n135 VTAIL.n134 2.84303
R338 VTAIL.n79 VTAIL.n78 2.84303
R339 VTAIL.n201 VTAIL.n180 2.71565
R340 VTAIL.n220 VTAIL.n219 2.71565
R341 VTAIL.n33 VTAIL.n12 2.71565
R342 VTAIL.n52 VTAIL.n51 2.71565
R343 VTAIL.n166 VTAIL.n165 2.71565
R344 VTAIL.n148 VTAIL.n127 2.71565
R345 VTAIL.n110 VTAIL.n109 2.71565
R346 VTAIL.n92 VTAIL.n71 2.71565
R347 VTAIL VTAIL.n223 2.39921
R348 VTAIL.n115 VTAIL.n113 2.10826
R349 VTAIL.n55 VTAIL.n1 2.10826
R350 VTAIL.n0 VTAIL.t4 1.99647
R351 VTAIL.n0 VTAIL.t2 1.99647
R352 VTAIL.n56 VTAIL.t5 1.99647
R353 VTAIL.n56 VTAIL.t8 1.99647
R354 VTAIL.n114 VTAIL.t6 1.99647
R355 VTAIL.n114 VTAIL.t7 1.99647
R356 VTAIL.n58 VTAIL.t3 1.99647
R357 VTAIL.n58 VTAIL.t1 1.99647
R358 VTAIL.n202 VTAIL.n178 1.93989
R359 VTAIL.n216 VTAIL.n172 1.93989
R360 VTAIL.n34 VTAIL.n10 1.93989
R361 VTAIL.n48 VTAIL.n4 1.93989
R362 VTAIL.n162 VTAIL.n118 1.93989
R363 VTAIL.n149 VTAIL.n125 1.93989
R364 VTAIL.n106 VTAIL.n62 1.93989
R365 VTAIL.n93 VTAIL.n69 1.93989
R366 VTAIL.n207 VTAIL.n205 1.16414
R367 VTAIL.n215 VTAIL.n174 1.16414
R368 VTAIL.n39 VTAIL.n37 1.16414
R369 VTAIL.n47 VTAIL.n6 1.16414
R370 VTAIL.n161 VTAIL.n120 1.16414
R371 VTAIL.n153 VTAIL.n152 1.16414
R372 VTAIL.n105 VTAIL.n64 1.16414
R373 VTAIL.n97 VTAIL.n96 1.16414
R374 VTAIL VTAIL.n1 0.877655
R375 VTAIL.n206 VTAIL.n176 0.388379
R376 VTAIL.n212 VTAIL.n211 0.388379
R377 VTAIL.n38 VTAIL.n8 0.388379
R378 VTAIL.n44 VTAIL.n43 0.388379
R379 VTAIL.n158 VTAIL.n157 0.388379
R380 VTAIL.n124 VTAIL.n122 0.388379
R381 VTAIL.n102 VTAIL.n101 0.388379
R382 VTAIL.n68 VTAIL.n66 0.388379
R383 VTAIL.n188 VTAIL.n183 0.155672
R384 VTAIL.n195 VTAIL.n183 0.155672
R385 VTAIL.n196 VTAIL.n195 0.155672
R386 VTAIL.n196 VTAIL.n179 0.155672
R387 VTAIL.n203 VTAIL.n179 0.155672
R388 VTAIL.n204 VTAIL.n203 0.155672
R389 VTAIL.n204 VTAIL.n175 0.155672
R390 VTAIL.n213 VTAIL.n175 0.155672
R391 VTAIL.n214 VTAIL.n213 0.155672
R392 VTAIL.n214 VTAIL.n171 0.155672
R393 VTAIL.n221 VTAIL.n171 0.155672
R394 VTAIL.n20 VTAIL.n15 0.155672
R395 VTAIL.n27 VTAIL.n15 0.155672
R396 VTAIL.n28 VTAIL.n27 0.155672
R397 VTAIL.n28 VTAIL.n11 0.155672
R398 VTAIL.n35 VTAIL.n11 0.155672
R399 VTAIL.n36 VTAIL.n35 0.155672
R400 VTAIL.n36 VTAIL.n7 0.155672
R401 VTAIL.n45 VTAIL.n7 0.155672
R402 VTAIL.n46 VTAIL.n45 0.155672
R403 VTAIL.n46 VTAIL.n3 0.155672
R404 VTAIL.n53 VTAIL.n3 0.155672
R405 VTAIL.n167 VTAIL.n117 0.155672
R406 VTAIL.n160 VTAIL.n117 0.155672
R407 VTAIL.n160 VTAIL.n159 0.155672
R408 VTAIL.n159 VTAIL.n121 0.155672
R409 VTAIL.n151 VTAIL.n121 0.155672
R410 VTAIL.n151 VTAIL.n150 0.155672
R411 VTAIL.n150 VTAIL.n126 0.155672
R412 VTAIL.n143 VTAIL.n126 0.155672
R413 VTAIL.n143 VTAIL.n142 0.155672
R414 VTAIL.n142 VTAIL.n130 0.155672
R415 VTAIL.n135 VTAIL.n130 0.155672
R416 VTAIL.n111 VTAIL.n61 0.155672
R417 VTAIL.n104 VTAIL.n61 0.155672
R418 VTAIL.n104 VTAIL.n103 0.155672
R419 VTAIL.n103 VTAIL.n65 0.155672
R420 VTAIL.n95 VTAIL.n65 0.155672
R421 VTAIL.n95 VTAIL.n94 0.155672
R422 VTAIL.n94 VTAIL.n70 0.155672
R423 VTAIL.n87 VTAIL.n70 0.155672
R424 VTAIL.n87 VTAIL.n86 0.155672
R425 VTAIL.n86 VTAIL.n74 0.155672
R426 VTAIL.n79 VTAIL.n74 0.155672
R427 VDD1.n48 VDD1.n0 289.615
R428 VDD1.n101 VDD1.n53 289.615
R429 VDD1.n49 VDD1.n48 185
R430 VDD1.n47 VDD1.n46 185
R431 VDD1.n4 VDD1.n3 185
R432 VDD1.n41 VDD1.n40 185
R433 VDD1.n39 VDD1.n6 185
R434 VDD1.n38 VDD1.n37 185
R435 VDD1.n9 VDD1.n7 185
R436 VDD1.n32 VDD1.n31 185
R437 VDD1.n30 VDD1.n29 185
R438 VDD1.n13 VDD1.n12 185
R439 VDD1.n24 VDD1.n23 185
R440 VDD1.n22 VDD1.n21 185
R441 VDD1.n17 VDD1.n16 185
R442 VDD1.n69 VDD1.n68 185
R443 VDD1.n74 VDD1.n73 185
R444 VDD1.n76 VDD1.n75 185
R445 VDD1.n65 VDD1.n64 185
R446 VDD1.n82 VDD1.n81 185
R447 VDD1.n84 VDD1.n83 185
R448 VDD1.n61 VDD1.n60 185
R449 VDD1.n91 VDD1.n90 185
R450 VDD1.n92 VDD1.n59 185
R451 VDD1.n94 VDD1.n93 185
R452 VDD1.n57 VDD1.n56 185
R453 VDD1.n100 VDD1.n99 185
R454 VDD1.n102 VDD1.n101 185
R455 VDD1.n18 VDD1.t2 149.524
R456 VDD1.n70 VDD1.t4 149.524
R457 VDD1.n48 VDD1.n47 104.615
R458 VDD1.n47 VDD1.n3 104.615
R459 VDD1.n40 VDD1.n3 104.615
R460 VDD1.n40 VDD1.n39 104.615
R461 VDD1.n39 VDD1.n38 104.615
R462 VDD1.n38 VDD1.n7 104.615
R463 VDD1.n31 VDD1.n7 104.615
R464 VDD1.n31 VDD1.n30 104.615
R465 VDD1.n30 VDD1.n12 104.615
R466 VDD1.n23 VDD1.n12 104.615
R467 VDD1.n23 VDD1.n22 104.615
R468 VDD1.n22 VDD1.n16 104.615
R469 VDD1.n74 VDD1.n68 104.615
R470 VDD1.n75 VDD1.n74 104.615
R471 VDD1.n75 VDD1.n64 104.615
R472 VDD1.n82 VDD1.n64 104.615
R473 VDD1.n83 VDD1.n82 104.615
R474 VDD1.n83 VDD1.n60 104.615
R475 VDD1.n91 VDD1.n60 104.615
R476 VDD1.n92 VDD1.n91 104.615
R477 VDD1.n93 VDD1.n92 104.615
R478 VDD1.n93 VDD1.n56 104.615
R479 VDD1.n100 VDD1.n56 104.615
R480 VDD1.n101 VDD1.n100 104.615
R481 VDD1.n107 VDD1.n106 62.628
R482 VDD1.n109 VDD1.n108 61.8644
R483 VDD1.t2 VDD1.n16 52.3082
R484 VDD1.t4 VDD1.n68 52.3082
R485 VDD1 VDD1.n52 50.6035
R486 VDD1.n107 VDD1.n105 50.4899
R487 VDD1.n109 VDD1.n107 45.1345
R488 VDD1.n41 VDD1.n6 13.1884
R489 VDD1.n94 VDD1.n59 13.1884
R490 VDD1.n42 VDD1.n4 12.8005
R491 VDD1.n37 VDD1.n8 12.8005
R492 VDD1.n90 VDD1.n89 12.8005
R493 VDD1.n95 VDD1.n57 12.8005
R494 VDD1.n46 VDD1.n45 12.0247
R495 VDD1.n36 VDD1.n9 12.0247
R496 VDD1.n88 VDD1.n61 12.0247
R497 VDD1.n99 VDD1.n98 12.0247
R498 VDD1.n49 VDD1.n2 11.249
R499 VDD1.n33 VDD1.n32 11.249
R500 VDD1.n85 VDD1.n84 11.249
R501 VDD1.n102 VDD1.n55 11.249
R502 VDD1.n50 VDD1.n0 10.4732
R503 VDD1.n29 VDD1.n11 10.4732
R504 VDD1.n81 VDD1.n63 10.4732
R505 VDD1.n103 VDD1.n53 10.4732
R506 VDD1.n18 VDD1.n17 10.2747
R507 VDD1.n70 VDD1.n69 10.2747
R508 VDD1.n28 VDD1.n13 9.69747
R509 VDD1.n80 VDD1.n65 9.69747
R510 VDD1.n52 VDD1.n51 9.45567
R511 VDD1.n105 VDD1.n104 9.45567
R512 VDD1.n20 VDD1.n19 9.3005
R513 VDD1.n15 VDD1.n14 9.3005
R514 VDD1.n26 VDD1.n25 9.3005
R515 VDD1.n28 VDD1.n27 9.3005
R516 VDD1.n11 VDD1.n10 9.3005
R517 VDD1.n34 VDD1.n33 9.3005
R518 VDD1.n36 VDD1.n35 9.3005
R519 VDD1.n8 VDD1.n5 9.3005
R520 VDD1.n51 VDD1.n50 9.3005
R521 VDD1.n2 VDD1.n1 9.3005
R522 VDD1.n45 VDD1.n44 9.3005
R523 VDD1.n43 VDD1.n42 9.3005
R524 VDD1.n104 VDD1.n103 9.3005
R525 VDD1.n55 VDD1.n54 9.3005
R526 VDD1.n98 VDD1.n97 9.3005
R527 VDD1.n96 VDD1.n95 9.3005
R528 VDD1.n72 VDD1.n71 9.3005
R529 VDD1.n67 VDD1.n66 9.3005
R530 VDD1.n78 VDD1.n77 9.3005
R531 VDD1.n80 VDD1.n79 9.3005
R532 VDD1.n63 VDD1.n62 9.3005
R533 VDD1.n86 VDD1.n85 9.3005
R534 VDD1.n88 VDD1.n87 9.3005
R535 VDD1.n89 VDD1.n58 9.3005
R536 VDD1.n25 VDD1.n24 8.92171
R537 VDD1.n77 VDD1.n76 8.92171
R538 VDD1.n21 VDD1.n15 8.14595
R539 VDD1.n73 VDD1.n67 8.14595
R540 VDD1.n20 VDD1.n17 7.3702
R541 VDD1.n72 VDD1.n69 7.3702
R542 VDD1.n21 VDD1.n20 5.81868
R543 VDD1.n73 VDD1.n72 5.81868
R544 VDD1.n24 VDD1.n15 5.04292
R545 VDD1.n76 VDD1.n67 5.04292
R546 VDD1.n25 VDD1.n13 4.26717
R547 VDD1.n77 VDD1.n65 4.26717
R548 VDD1.n52 VDD1.n0 3.49141
R549 VDD1.n29 VDD1.n28 3.49141
R550 VDD1.n81 VDD1.n80 3.49141
R551 VDD1.n105 VDD1.n53 3.49141
R552 VDD1.n19 VDD1.n18 2.84303
R553 VDD1.n71 VDD1.n70 2.84303
R554 VDD1.n50 VDD1.n49 2.71565
R555 VDD1.n32 VDD1.n11 2.71565
R556 VDD1.n84 VDD1.n63 2.71565
R557 VDD1.n103 VDD1.n102 2.71565
R558 VDD1.n108 VDD1.t0 1.99647
R559 VDD1.n108 VDD1.t5 1.99647
R560 VDD1.n106 VDD1.t1 1.99647
R561 VDD1.n106 VDD1.t3 1.99647
R562 VDD1.n46 VDD1.n2 1.93989
R563 VDD1.n33 VDD1.n9 1.93989
R564 VDD1.n85 VDD1.n61 1.93989
R565 VDD1.n99 VDD1.n55 1.93989
R566 VDD1.n45 VDD1.n4 1.16414
R567 VDD1.n37 VDD1.n36 1.16414
R568 VDD1.n90 VDD1.n88 1.16414
R569 VDD1.n98 VDD1.n57 1.16414
R570 VDD1 VDD1.n109 0.761276
R571 VDD1.n42 VDD1.n41 0.388379
R572 VDD1.n8 VDD1.n6 0.388379
R573 VDD1.n89 VDD1.n59 0.388379
R574 VDD1.n95 VDD1.n94 0.388379
R575 VDD1.n51 VDD1.n1 0.155672
R576 VDD1.n44 VDD1.n1 0.155672
R577 VDD1.n44 VDD1.n43 0.155672
R578 VDD1.n43 VDD1.n5 0.155672
R579 VDD1.n35 VDD1.n5 0.155672
R580 VDD1.n35 VDD1.n34 0.155672
R581 VDD1.n34 VDD1.n10 0.155672
R582 VDD1.n27 VDD1.n10 0.155672
R583 VDD1.n27 VDD1.n26 0.155672
R584 VDD1.n26 VDD1.n14 0.155672
R585 VDD1.n19 VDD1.n14 0.155672
R586 VDD1.n71 VDD1.n66 0.155672
R587 VDD1.n78 VDD1.n66 0.155672
R588 VDD1.n79 VDD1.n78 0.155672
R589 VDD1.n79 VDD1.n62 0.155672
R590 VDD1.n86 VDD1.n62 0.155672
R591 VDD1.n87 VDD1.n86 0.155672
R592 VDD1.n87 VDD1.n58 0.155672
R593 VDD1.n96 VDD1.n58 0.155672
R594 VDD1.n97 VDD1.n96 0.155672
R595 VDD1.n97 VDD1.n54 0.155672
R596 VDD1.n104 VDD1.n54 0.155672
R597 B.n843 B.n842 585
R598 B.n844 B.n843 585
R599 B.n303 B.n138 585
R600 B.n302 B.n301 585
R601 B.n300 B.n299 585
R602 B.n298 B.n297 585
R603 B.n296 B.n295 585
R604 B.n294 B.n293 585
R605 B.n292 B.n291 585
R606 B.n290 B.n289 585
R607 B.n288 B.n287 585
R608 B.n286 B.n285 585
R609 B.n284 B.n283 585
R610 B.n282 B.n281 585
R611 B.n280 B.n279 585
R612 B.n278 B.n277 585
R613 B.n276 B.n275 585
R614 B.n274 B.n273 585
R615 B.n272 B.n271 585
R616 B.n270 B.n269 585
R617 B.n268 B.n267 585
R618 B.n266 B.n265 585
R619 B.n264 B.n263 585
R620 B.n262 B.n261 585
R621 B.n260 B.n259 585
R622 B.n258 B.n257 585
R623 B.n256 B.n255 585
R624 B.n254 B.n253 585
R625 B.n252 B.n251 585
R626 B.n250 B.n249 585
R627 B.n248 B.n247 585
R628 B.n246 B.n245 585
R629 B.n244 B.n243 585
R630 B.n242 B.n241 585
R631 B.n240 B.n239 585
R632 B.n238 B.n237 585
R633 B.n236 B.n235 585
R634 B.n233 B.n232 585
R635 B.n231 B.n230 585
R636 B.n229 B.n228 585
R637 B.n227 B.n226 585
R638 B.n225 B.n224 585
R639 B.n223 B.n222 585
R640 B.n221 B.n220 585
R641 B.n219 B.n218 585
R642 B.n217 B.n216 585
R643 B.n215 B.n214 585
R644 B.n213 B.n212 585
R645 B.n211 B.n210 585
R646 B.n209 B.n208 585
R647 B.n207 B.n206 585
R648 B.n205 B.n204 585
R649 B.n203 B.n202 585
R650 B.n201 B.n200 585
R651 B.n199 B.n198 585
R652 B.n197 B.n196 585
R653 B.n195 B.n194 585
R654 B.n193 B.n192 585
R655 B.n191 B.n190 585
R656 B.n189 B.n188 585
R657 B.n187 B.n186 585
R658 B.n185 B.n184 585
R659 B.n183 B.n182 585
R660 B.n181 B.n180 585
R661 B.n179 B.n178 585
R662 B.n177 B.n176 585
R663 B.n175 B.n174 585
R664 B.n173 B.n172 585
R665 B.n171 B.n170 585
R666 B.n169 B.n168 585
R667 B.n167 B.n166 585
R668 B.n165 B.n164 585
R669 B.n163 B.n162 585
R670 B.n161 B.n160 585
R671 B.n159 B.n158 585
R672 B.n157 B.n156 585
R673 B.n155 B.n154 585
R674 B.n153 B.n152 585
R675 B.n151 B.n150 585
R676 B.n149 B.n148 585
R677 B.n147 B.n146 585
R678 B.n145 B.n144 585
R679 B.n841 B.n97 585
R680 B.n845 B.n97 585
R681 B.n840 B.n96 585
R682 B.n846 B.n96 585
R683 B.n839 B.n838 585
R684 B.n838 B.n92 585
R685 B.n837 B.n91 585
R686 B.n852 B.n91 585
R687 B.n836 B.n90 585
R688 B.n853 B.n90 585
R689 B.n835 B.n89 585
R690 B.n854 B.n89 585
R691 B.n834 B.n833 585
R692 B.n833 B.n85 585
R693 B.n832 B.n84 585
R694 B.n860 B.n84 585
R695 B.n831 B.n83 585
R696 B.n861 B.n83 585
R697 B.n830 B.n82 585
R698 B.n862 B.n82 585
R699 B.n829 B.n828 585
R700 B.n828 B.n78 585
R701 B.n827 B.n77 585
R702 B.n868 B.n77 585
R703 B.n826 B.n76 585
R704 B.n869 B.n76 585
R705 B.n825 B.n75 585
R706 B.n870 B.n75 585
R707 B.n824 B.n823 585
R708 B.n823 B.n71 585
R709 B.n822 B.n70 585
R710 B.n876 B.n70 585
R711 B.n821 B.n69 585
R712 B.n877 B.n69 585
R713 B.n820 B.n68 585
R714 B.n878 B.n68 585
R715 B.n819 B.n818 585
R716 B.n818 B.n64 585
R717 B.n817 B.n63 585
R718 B.n884 B.n63 585
R719 B.n816 B.n62 585
R720 B.n885 B.n62 585
R721 B.n815 B.n61 585
R722 B.n886 B.n61 585
R723 B.n814 B.n813 585
R724 B.n813 B.n57 585
R725 B.n812 B.n56 585
R726 B.n892 B.n56 585
R727 B.n811 B.n55 585
R728 B.n893 B.n55 585
R729 B.n810 B.n54 585
R730 B.n894 B.n54 585
R731 B.n809 B.n808 585
R732 B.n808 B.n50 585
R733 B.n807 B.n49 585
R734 B.n900 B.n49 585
R735 B.n806 B.n48 585
R736 B.n901 B.n48 585
R737 B.n805 B.n47 585
R738 B.n902 B.n47 585
R739 B.n804 B.n803 585
R740 B.n803 B.n43 585
R741 B.n802 B.n42 585
R742 B.n908 B.n42 585
R743 B.n801 B.n41 585
R744 B.n909 B.n41 585
R745 B.n800 B.n40 585
R746 B.n910 B.n40 585
R747 B.n799 B.n798 585
R748 B.n798 B.n39 585
R749 B.n797 B.n35 585
R750 B.n916 B.n35 585
R751 B.n796 B.n34 585
R752 B.n917 B.n34 585
R753 B.n795 B.n33 585
R754 B.n918 B.n33 585
R755 B.n794 B.n793 585
R756 B.n793 B.n29 585
R757 B.n792 B.n28 585
R758 B.n924 B.n28 585
R759 B.n791 B.n27 585
R760 B.n925 B.n27 585
R761 B.n790 B.n26 585
R762 B.n926 B.n26 585
R763 B.n789 B.n788 585
R764 B.n788 B.n22 585
R765 B.n787 B.n21 585
R766 B.n932 B.n21 585
R767 B.n786 B.n20 585
R768 B.n933 B.n20 585
R769 B.n785 B.n19 585
R770 B.n934 B.n19 585
R771 B.n784 B.n783 585
R772 B.n783 B.n15 585
R773 B.n782 B.n14 585
R774 B.n940 B.n14 585
R775 B.n781 B.n13 585
R776 B.n941 B.n13 585
R777 B.n780 B.n12 585
R778 B.n942 B.n12 585
R779 B.n779 B.n778 585
R780 B.n778 B.n8 585
R781 B.n777 B.n7 585
R782 B.n948 B.n7 585
R783 B.n776 B.n6 585
R784 B.n949 B.n6 585
R785 B.n775 B.n5 585
R786 B.n950 B.n5 585
R787 B.n774 B.n773 585
R788 B.n773 B.n4 585
R789 B.n772 B.n304 585
R790 B.n772 B.n771 585
R791 B.n762 B.n305 585
R792 B.n306 B.n305 585
R793 B.n764 B.n763 585
R794 B.n765 B.n764 585
R795 B.n761 B.n311 585
R796 B.n311 B.n310 585
R797 B.n760 B.n759 585
R798 B.n759 B.n758 585
R799 B.n313 B.n312 585
R800 B.n314 B.n313 585
R801 B.n751 B.n750 585
R802 B.n752 B.n751 585
R803 B.n749 B.n319 585
R804 B.n319 B.n318 585
R805 B.n748 B.n747 585
R806 B.n747 B.n746 585
R807 B.n321 B.n320 585
R808 B.n322 B.n321 585
R809 B.n739 B.n738 585
R810 B.n740 B.n739 585
R811 B.n737 B.n327 585
R812 B.n327 B.n326 585
R813 B.n736 B.n735 585
R814 B.n735 B.n734 585
R815 B.n329 B.n328 585
R816 B.n330 B.n329 585
R817 B.n727 B.n726 585
R818 B.n728 B.n727 585
R819 B.n725 B.n335 585
R820 B.n335 B.n334 585
R821 B.n724 B.n723 585
R822 B.n723 B.n722 585
R823 B.n337 B.n336 585
R824 B.n715 B.n337 585
R825 B.n714 B.n713 585
R826 B.n716 B.n714 585
R827 B.n712 B.n342 585
R828 B.n342 B.n341 585
R829 B.n711 B.n710 585
R830 B.n710 B.n709 585
R831 B.n344 B.n343 585
R832 B.n345 B.n344 585
R833 B.n702 B.n701 585
R834 B.n703 B.n702 585
R835 B.n700 B.n350 585
R836 B.n350 B.n349 585
R837 B.n699 B.n698 585
R838 B.n698 B.n697 585
R839 B.n352 B.n351 585
R840 B.n353 B.n352 585
R841 B.n690 B.n689 585
R842 B.n691 B.n690 585
R843 B.n688 B.n358 585
R844 B.n358 B.n357 585
R845 B.n687 B.n686 585
R846 B.n686 B.n685 585
R847 B.n360 B.n359 585
R848 B.n361 B.n360 585
R849 B.n678 B.n677 585
R850 B.n679 B.n678 585
R851 B.n676 B.n366 585
R852 B.n366 B.n365 585
R853 B.n675 B.n674 585
R854 B.n674 B.n673 585
R855 B.n368 B.n367 585
R856 B.n369 B.n368 585
R857 B.n666 B.n665 585
R858 B.n667 B.n666 585
R859 B.n664 B.n374 585
R860 B.n374 B.n373 585
R861 B.n663 B.n662 585
R862 B.n662 B.n661 585
R863 B.n376 B.n375 585
R864 B.n377 B.n376 585
R865 B.n654 B.n653 585
R866 B.n655 B.n654 585
R867 B.n652 B.n382 585
R868 B.n382 B.n381 585
R869 B.n651 B.n650 585
R870 B.n650 B.n649 585
R871 B.n384 B.n383 585
R872 B.n385 B.n384 585
R873 B.n642 B.n641 585
R874 B.n643 B.n642 585
R875 B.n640 B.n390 585
R876 B.n390 B.n389 585
R877 B.n639 B.n638 585
R878 B.n638 B.n637 585
R879 B.n392 B.n391 585
R880 B.n393 B.n392 585
R881 B.n630 B.n629 585
R882 B.n631 B.n630 585
R883 B.n628 B.n398 585
R884 B.n398 B.n397 585
R885 B.n627 B.n626 585
R886 B.n626 B.n625 585
R887 B.n400 B.n399 585
R888 B.n401 B.n400 585
R889 B.n618 B.n617 585
R890 B.n619 B.n618 585
R891 B.n616 B.n406 585
R892 B.n406 B.n405 585
R893 B.n610 B.n609 585
R894 B.n608 B.n448 585
R895 B.n607 B.n447 585
R896 B.n612 B.n447 585
R897 B.n606 B.n605 585
R898 B.n604 B.n603 585
R899 B.n602 B.n601 585
R900 B.n600 B.n599 585
R901 B.n598 B.n597 585
R902 B.n596 B.n595 585
R903 B.n594 B.n593 585
R904 B.n592 B.n591 585
R905 B.n590 B.n589 585
R906 B.n588 B.n587 585
R907 B.n586 B.n585 585
R908 B.n584 B.n583 585
R909 B.n582 B.n581 585
R910 B.n580 B.n579 585
R911 B.n578 B.n577 585
R912 B.n576 B.n575 585
R913 B.n574 B.n573 585
R914 B.n572 B.n571 585
R915 B.n570 B.n569 585
R916 B.n568 B.n567 585
R917 B.n566 B.n565 585
R918 B.n564 B.n563 585
R919 B.n562 B.n561 585
R920 B.n560 B.n559 585
R921 B.n558 B.n557 585
R922 B.n556 B.n555 585
R923 B.n554 B.n553 585
R924 B.n552 B.n551 585
R925 B.n550 B.n549 585
R926 B.n548 B.n547 585
R927 B.n546 B.n545 585
R928 B.n544 B.n543 585
R929 B.n542 B.n541 585
R930 B.n539 B.n538 585
R931 B.n537 B.n536 585
R932 B.n535 B.n534 585
R933 B.n533 B.n532 585
R934 B.n531 B.n530 585
R935 B.n529 B.n528 585
R936 B.n527 B.n526 585
R937 B.n525 B.n524 585
R938 B.n523 B.n522 585
R939 B.n521 B.n520 585
R940 B.n519 B.n518 585
R941 B.n517 B.n516 585
R942 B.n515 B.n514 585
R943 B.n513 B.n512 585
R944 B.n511 B.n510 585
R945 B.n509 B.n508 585
R946 B.n507 B.n506 585
R947 B.n505 B.n504 585
R948 B.n503 B.n502 585
R949 B.n501 B.n500 585
R950 B.n499 B.n498 585
R951 B.n497 B.n496 585
R952 B.n495 B.n494 585
R953 B.n493 B.n492 585
R954 B.n491 B.n490 585
R955 B.n489 B.n488 585
R956 B.n487 B.n486 585
R957 B.n485 B.n484 585
R958 B.n483 B.n482 585
R959 B.n481 B.n480 585
R960 B.n479 B.n478 585
R961 B.n477 B.n476 585
R962 B.n475 B.n474 585
R963 B.n473 B.n472 585
R964 B.n471 B.n470 585
R965 B.n469 B.n468 585
R966 B.n467 B.n466 585
R967 B.n465 B.n464 585
R968 B.n463 B.n462 585
R969 B.n461 B.n460 585
R970 B.n459 B.n458 585
R971 B.n457 B.n456 585
R972 B.n455 B.n454 585
R973 B.n408 B.n407 585
R974 B.n615 B.n614 585
R975 B.n404 B.n403 585
R976 B.n405 B.n404 585
R977 B.n621 B.n620 585
R978 B.n620 B.n619 585
R979 B.n622 B.n402 585
R980 B.n402 B.n401 585
R981 B.n624 B.n623 585
R982 B.n625 B.n624 585
R983 B.n396 B.n395 585
R984 B.n397 B.n396 585
R985 B.n633 B.n632 585
R986 B.n632 B.n631 585
R987 B.n634 B.n394 585
R988 B.n394 B.n393 585
R989 B.n636 B.n635 585
R990 B.n637 B.n636 585
R991 B.n388 B.n387 585
R992 B.n389 B.n388 585
R993 B.n645 B.n644 585
R994 B.n644 B.n643 585
R995 B.n646 B.n386 585
R996 B.n386 B.n385 585
R997 B.n648 B.n647 585
R998 B.n649 B.n648 585
R999 B.n380 B.n379 585
R1000 B.n381 B.n380 585
R1001 B.n657 B.n656 585
R1002 B.n656 B.n655 585
R1003 B.n658 B.n378 585
R1004 B.n378 B.n377 585
R1005 B.n660 B.n659 585
R1006 B.n661 B.n660 585
R1007 B.n372 B.n371 585
R1008 B.n373 B.n372 585
R1009 B.n669 B.n668 585
R1010 B.n668 B.n667 585
R1011 B.n670 B.n370 585
R1012 B.n370 B.n369 585
R1013 B.n672 B.n671 585
R1014 B.n673 B.n672 585
R1015 B.n364 B.n363 585
R1016 B.n365 B.n364 585
R1017 B.n681 B.n680 585
R1018 B.n680 B.n679 585
R1019 B.n682 B.n362 585
R1020 B.n362 B.n361 585
R1021 B.n684 B.n683 585
R1022 B.n685 B.n684 585
R1023 B.n356 B.n355 585
R1024 B.n357 B.n356 585
R1025 B.n693 B.n692 585
R1026 B.n692 B.n691 585
R1027 B.n694 B.n354 585
R1028 B.n354 B.n353 585
R1029 B.n696 B.n695 585
R1030 B.n697 B.n696 585
R1031 B.n348 B.n347 585
R1032 B.n349 B.n348 585
R1033 B.n705 B.n704 585
R1034 B.n704 B.n703 585
R1035 B.n706 B.n346 585
R1036 B.n346 B.n345 585
R1037 B.n708 B.n707 585
R1038 B.n709 B.n708 585
R1039 B.n340 B.n339 585
R1040 B.n341 B.n340 585
R1041 B.n718 B.n717 585
R1042 B.n717 B.n716 585
R1043 B.n719 B.n338 585
R1044 B.n715 B.n338 585
R1045 B.n721 B.n720 585
R1046 B.n722 B.n721 585
R1047 B.n333 B.n332 585
R1048 B.n334 B.n333 585
R1049 B.n730 B.n729 585
R1050 B.n729 B.n728 585
R1051 B.n731 B.n331 585
R1052 B.n331 B.n330 585
R1053 B.n733 B.n732 585
R1054 B.n734 B.n733 585
R1055 B.n325 B.n324 585
R1056 B.n326 B.n325 585
R1057 B.n742 B.n741 585
R1058 B.n741 B.n740 585
R1059 B.n743 B.n323 585
R1060 B.n323 B.n322 585
R1061 B.n745 B.n744 585
R1062 B.n746 B.n745 585
R1063 B.n317 B.n316 585
R1064 B.n318 B.n317 585
R1065 B.n754 B.n753 585
R1066 B.n753 B.n752 585
R1067 B.n755 B.n315 585
R1068 B.n315 B.n314 585
R1069 B.n757 B.n756 585
R1070 B.n758 B.n757 585
R1071 B.n309 B.n308 585
R1072 B.n310 B.n309 585
R1073 B.n767 B.n766 585
R1074 B.n766 B.n765 585
R1075 B.n768 B.n307 585
R1076 B.n307 B.n306 585
R1077 B.n770 B.n769 585
R1078 B.n771 B.n770 585
R1079 B.n2 B.n0 585
R1080 B.n4 B.n2 585
R1081 B.n3 B.n1 585
R1082 B.n949 B.n3 585
R1083 B.n947 B.n946 585
R1084 B.n948 B.n947 585
R1085 B.n945 B.n9 585
R1086 B.n9 B.n8 585
R1087 B.n944 B.n943 585
R1088 B.n943 B.n942 585
R1089 B.n11 B.n10 585
R1090 B.n941 B.n11 585
R1091 B.n939 B.n938 585
R1092 B.n940 B.n939 585
R1093 B.n937 B.n16 585
R1094 B.n16 B.n15 585
R1095 B.n936 B.n935 585
R1096 B.n935 B.n934 585
R1097 B.n18 B.n17 585
R1098 B.n933 B.n18 585
R1099 B.n931 B.n930 585
R1100 B.n932 B.n931 585
R1101 B.n929 B.n23 585
R1102 B.n23 B.n22 585
R1103 B.n928 B.n927 585
R1104 B.n927 B.n926 585
R1105 B.n25 B.n24 585
R1106 B.n925 B.n25 585
R1107 B.n923 B.n922 585
R1108 B.n924 B.n923 585
R1109 B.n921 B.n30 585
R1110 B.n30 B.n29 585
R1111 B.n920 B.n919 585
R1112 B.n919 B.n918 585
R1113 B.n32 B.n31 585
R1114 B.n917 B.n32 585
R1115 B.n915 B.n914 585
R1116 B.n916 B.n915 585
R1117 B.n913 B.n36 585
R1118 B.n39 B.n36 585
R1119 B.n912 B.n911 585
R1120 B.n911 B.n910 585
R1121 B.n38 B.n37 585
R1122 B.n909 B.n38 585
R1123 B.n907 B.n906 585
R1124 B.n908 B.n907 585
R1125 B.n905 B.n44 585
R1126 B.n44 B.n43 585
R1127 B.n904 B.n903 585
R1128 B.n903 B.n902 585
R1129 B.n46 B.n45 585
R1130 B.n901 B.n46 585
R1131 B.n899 B.n898 585
R1132 B.n900 B.n899 585
R1133 B.n897 B.n51 585
R1134 B.n51 B.n50 585
R1135 B.n896 B.n895 585
R1136 B.n895 B.n894 585
R1137 B.n53 B.n52 585
R1138 B.n893 B.n53 585
R1139 B.n891 B.n890 585
R1140 B.n892 B.n891 585
R1141 B.n889 B.n58 585
R1142 B.n58 B.n57 585
R1143 B.n888 B.n887 585
R1144 B.n887 B.n886 585
R1145 B.n60 B.n59 585
R1146 B.n885 B.n60 585
R1147 B.n883 B.n882 585
R1148 B.n884 B.n883 585
R1149 B.n881 B.n65 585
R1150 B.n65 B.n64 585
R1151 B.n880 B.n879 585
R1152 B.n879 B.n878 585
R1153 B.n67 B.n66 585
R1154 B.n877 B.n67 585
R1155 B.n875 B.n874 585
R1156 B.n876 B.n875 585
R1157 B.n873 B.n72 585
R1158 B.n72 B.n71 585
R1159 B.n872 B.n871 585
R1160 B.n871 B.n870 585
R1161 B.n74 B.n73 585
R1162 B.n869 B.n74 585
R1163 B.n867 B.n866 585
R1164 B.n868 B.n867 585
R1165 B.n865 B.n79 585
R1166 B.n79 B.n78 585
R1167 B.n864 B.n863 585
R1168 B.n863 B.n862 585
R1169 B.n81 B.n80 585
R1170 B.n861 B.n81 585
R1171 B.n859 B.n858 585
R1172 B.n860 B.n859 585
R1173 B.n857 B.n86 585
R1174 B.n86 B.n85 585
R1175 B.n856 B.n855 585
R1176 B.n855 B.n854 585
R1177 B.n88 B.n87 585
R1178 B.n853 B.n88 585
R1179 B.n851 B.n850 585
R1180 B.n852 B.n851 585
R1181 B.n849 B.n93 585
R1182 B.n93 B.n92 585
R1183 B.n848 B.n847 585
R1184 B.n847 B.n846 585
R1185 B.n95 B.n94 585
R1186 B.n845 B.n95 585
R1187 B.n952 B.n951 585
R1188 B.n951 B.n950 585
R1189 B.n610 B.n404 434.841
R1190 B.n144 B.n95 434.841
R1191 B.n614 B.n406 434.841
R1192 B.n843 B.n97 434.841
R1193 B.n451 B.t15 319.793
R1194 B.n139 B.t17 319.793
R1195 B.n449 B.t12 319.793
R1196 B.n141 B.t7 319.793
R1197 B.n451 B.t13 277.964
R1198 B.n449 B.t9 277.964
R1199 B.n141 B.t5 277.964
R1200 B.n139 B.t16 277.964
R1201 B.n844 B.n137 256.663
R1202 B.n844 B.n136 256.663
R1203 B.n844 B.n135 256.663
R1204 B.n844 B.n134 256.663
R1205 B.n844 B.n133 256.663
R1206 B.n844 B.n132 256.663
R1207 B.n844 B.n131 256.663
R1208 B.n844 B.n130 256.663
R1209 B.n844 B.n129 256.663
R1210 B.n844 B.n128 256.663
R1211 B.n844 B.n127 256.663
R1212 B.n844 B.n126 256.663
R1213 B.n844 B.n125 256.663
R1214 B.n844 B.n124 256.663
R1215 B.n844 B.n123 256.663
R1216 B.n844 B.n122 256.663
R1217 B.n844 B.n121 256.663
R1218 B.n844 B.n120 256.663
R1219 B.n844 B.n119 256.663
R1220 B.n844 B.n118 256.663
R1221 B.n844 B.n117 256.663
R1222 B.n844 B.n116 256.663
R1223 B.n844 B.n115 256.663
R1224 B.n844 B.n114 256.663
R1225 B.n844 B.n113 256.663
R1226 B.n844 B.n112 256.663
R1227 B.n844 B.n111 256.663
R1228 B.n844 B.n110 256.663
R1229 B.n844 B.n109 256.663
R1230 B.n844 B.n108 256.663
R1231 B.n844 B.n107 256.663
R1232 B.n844 B.n106 256.663
R1233 B.n844 B.n105 256.663
R1234 B.n844 B.n104 256.663
R1235 B.n844 B.n103 256.663
R1236 B.n844 B.n102 256.663
R1237 B.n844 B.n101 256.663
R1238 B.n844 B.n100 256.663
R1239 B.n844 B.n99 256.663
R1240 B.n844 B.n98 256.663
R1241 B.n612 B.n611 256.663
R1242 B.n612 B.n409 256.663
R1243 B.n612 B.n410 256.663
R1244 B.n612 B.n411 256.663
R1245 B.n612 B.n412 256.663
R1246 B.n612 B.n413 256.663
R1247 B.n612 B.n414 256.663
R1248 B.n612 B.n415 256.663
R1249 B.n612 B.n416 256.663
R1250 B.n612 B.n417 256.663
R1251 B.n612 B.n418 256.663
R1252 B.n612 B.n419 256.663
R1253 B.n612 B.n420 256.663
R1254 B.n612 B.n421 256.663
R1255 B.n612 B.n422 256.663
R1256 B.n612 B.n423 256.663
R1257 B.n612 B.n424 256.663
R1258 B.n612 B.n425 256.663
R1259 B.n612 B.n426 256.663
R1260 B.n612 B.n427 256.663
R1261 B.n612 B.n428 256.663
R1262 B.n612 B.n429 256.663
R1263 B.n612 B.n430 256.663
R1264 B.n612 B.n431 256.663
R1265 B.n612 B.n432 256.663
R1266 B.n612 B.n433 256.663
R1267 B.n612 B.n434 256.663
R1268 B.n612 B.n435 256.663
R1269 B.n612 B.n436 256.663
R1270 B.n612 B.n437 256.663
R1271 B.n612 B.n438 256.663
R1272 B.n612 B.n439 256.663
R1273 B.n612 B.n440 256.663
R1274 B.n612 B.n441 256.663
R1275 B.n612 B.n442 256.663
R1276 B.n612 B.n443 256.663
R1277 B.n612 B.n444 256.663
R1278 B.n612 B.n445 256.663
R1279 B.n612 B.n446 256.663
R1280 B.n613 B.n612 256.663
R1281 B.n452 B.t14 246.095
R1282 B.n140 B.t18 246.095
R1283 B.n450 B.t11 246.095
R1284 B.n142 B.t8 246.095
R1285 B.n620 B.n404 163.367
R1286 B.n620 B.n402 163.367
R1287 B.n624 B.n402 163.367
R1288 B.n624 B.n396 163.367
R1289 B.n632 B.n396 163.367
R1290 B.n632 B.n394 163.367
R1291 B.n636 B.n394 163.367
R1292 B.n636 B.n388 163.367
R1293 B.n644 B.n388 163.367
R1294 B.n644 B.n386 163.367
R1295 B.n648 B.n386 163.367
R1296 B.n648 B.n380 163.367
R1297 B.n656 B.n380 163.367
R1298 B.n656 B.n378 163.367
R1299 B.n660 B.n378 163.367
R1300 B.n660 B.n372 163.367
R1301 B.n668 B.n372 163.367
R1302 B.n668 B.n370 163.367
R1303 B.n672 B.n370 163.367
R1304 B.n672 B.n364 163.367
R1305 B.n680 B.n364 163.367
R1306 B.n680 B.n362 163.367
R1307 B.n684 B.n362 163.367
R1308 B.n684 B.n356 163.367
R1309 B.n692 B.n356 163.367
R1310 B.n692 B.n354 163.367
R1311 B.n696 B.n354 163.367
R1312 B.n696 B.n348 163.367
R1313 B.n704 B.n348 163.367
R1314 B.n704 B.n346 163.367
R1315 B.n708 B.n346 163.367
R1316 B.n708 B.n340 163.367
R1317 B.n717 B.n340 163.367
R1318 B.n717 B.n338 163.367
R1319 B.n721 B.n338 163.367
R1320 B.n721 B.n333 163.367
R1321 B.n729 B.n333 163.367
R1322 B.n729 B.n331 163.367
R1323 B.n733 B.n331 163.367
R1324 B.n733 B.n325 163.367
R1325 B.n741 B.n325 163.367
R1326 B.n741 B.n323 163.367
R1327 B.n745 B.n323 163.367
R1328 B.n745 B.n317 163.367
R1329 B.n753 B.n317 163.367
R1330 B.n753 B.n315 163.367
R1331 B.n757 B.n315 163.367
R1332 B.n757 B.n309 163.367
R1333 B.n766 B.n309 163.367
R1334 B.n766 B.n307 163.367
R1335 B.n770 B.n307 163.367
R1336 B.n770 B.n2 163.367
R1337 B.n951 B.n2 163.367
R1338 B.n951 B.n3 163.367
R1339 B.n947 B.n3 163.367
R1340 B.n947 B.n9 163.367
R1341 B.n943 B.n9 163.367
R1342 B.n943 B.n11 163.367
R1343 B.n939 B.n11 163.367
R1344 B.n939 B.n16 163.367
R1345 B.n935 B.n16 163.367
R1346 B.n935 B.n18 163.367
R1347 B.n931 B.n18 163.367
R1348 B.n931 B.n23 163.367
R1349 B.n927 B.n23 163.367
R1350 B.n927 B.n25 163.367
R1351 B.n923 B.n25 163.367
R1352 B.n923 B.n30 163.367
R1353 B.n919 B.n30 163.367
R1354 B.n919 B.n32 163.367
R1355 B.n915 B.n32 163.367
R1356 B.n915 B.n36 163.367
R1357 B.n911 B.n36 163.367
R1358 B.n911 B.n38 163.367
R1359 B.n907 B.n38 163.367
R1360 B.n907 B.n44 163.367
R1361 B.n903 B.n44 163.367
R1362 B.n903 B.n46 163.367
R1363 B.n899 B.n46 163.367
R1364 B.n899 B.n51 163.367
R1365 B.n895 B.n51 163.367
R1366 B.n895 B.n53 163.367
R1367 B.n891 B.n53 163.367
R1368 B.n891 B.n58 163.367
R1369 B.n887 B.n58 163.367
R1370 B.n887 B.n60 163.367
R1371 B.n883 B.n60 163.367
R1372 B.n883 B.n65 163.367
R1373 B.n879 B.n65 163.367
R1374 B.n879 B.n67 163.367
R1375 B.n875 B.n67 163.367
R1376 B.n875 B.n72 163.367
R1377 B.n871 B.n72 163.367
R1378 B.n871 B.n74 163.367
R1379 B.n867 B.n74 163.367
R1380 B.n867 B.n79 163.367
R1381 B.n863 B.n79 163.367
R1382 B.n863 B.n81 163.367
R1383 B.n859 B.n81 163.367
R1384 B.n859 B.n86 163.367
R1385 B.n855 B.n86 163.367
R1386 B.n855 B.n88 163.367
R1387 B.n851 B.n88 163.367
R1388 B.n851 B.n93 163.367
R1389 B.n847 B.n93 163.367
R1390 B.n847 B.n95 163.367
R1391 B.n448 B.n447 163.367
R1392 B.n605 B.n447 163.367
R1393 B.n603 B.n602 163.367
R1394 B.n599 B.n598 163.367
R1395 B.n595 B.n594 163.367
R1396 B.n591 B.n590 163.367
R1397 B.n587 B.n586 163.367
R1398 B.n583 B.n582 163.367
R1399 B.n579 B.n578 163.367
R1400 B.n575 B.n574 163.367
R1401 B.n571 B.n570 163.367
R1402 B.n567 B.n566 163.367
R1403 B.n563 B.n562 163.367
R1404 B.n559 B.n558 163.367
R1405 B.n555 B.n554 163.367
R1406 B.n551 B.n550 163.367
R1407 B.n547 B.n546 163.367
R1408 B.n543 B.n542 163.367
R1409 B.n538 B.n537 163.367
R1410 B.n534 B.n533 163.367
R1411 B.n530 B.n529 163.367
R1412 B.n526 B.n525 163.367
R1413 B.n522 B.n521 163.367
R1414 B.n518 B.n517 163.367
R1415 B.n514 B.n513 163.367
R1416 B.n510 B.n509 163.367
R1417 B.n506 B.n505 163.367
R1418 B.n502 B.n501 163.367
R1419 B.n498 B.n497 163.367
R1420 B.n494 B.n493 163.367
R1421 B.n490 B.n489 163.367
R1422 B.n486 B.n485 163.367
R1423 B.n482 B.n481 163.367
R1424 B.n478 B.n477 163.367
R1425 B.n474 B.n473 163.367
R1426 B.n470 B.n469 163.367
R1427 B.n466 B.n465 163.367
R1428 B.n462 B.n461 163.367
R1429 B.n458 B.n457 163.367
R1430 B.n454 B.n408 163.367
R1431 B.n618 B.n406 163.367
R1432 B.n618 B.n400 163.367
R1433 B.n626 B.n400 163.367
R1434 B.n626 B.n398 163.367
R1435 B.n630 B.n398 163.367
R1436 B.n630 B.n392 163.367
R1437 B.n638 B.n392 163.367
R1438 B.n638 B.n390 163.367
R1439 B.n642 B.n390 163.367
R1440 B.n642 B.n384 163.367
R1441 B.n650 B.n384 163.367
R1442 B.n650 B.n382 163.367
R1443 B.n654 B.n382 163.367
R1444 B.n654 B.n376 163.367
R1445 B.n662 B.n376 163.367
R1446 B.n662 B.n374 163.367
R1447 B.n666 B.n374 163.367
R1448 B.n666 B.n368 163.367
R1449 B.n674 B.n368 163.367
R1450 B.n674 B.n366 163.367
R1451 B.n678 B.n366 163.367
R1452 B.n678 B.n360 163.367
R1453 B.n686 B.n360 163.367
R1454 B.n686 B.n358 163.367
R1455 B.n690 B.n358 163.367
R1456 B.n690 B.n352 163.367
R1457 B.n698 B.n352 163.367
R1458 B.n698 B.n350 163.367
R1459 B.n702 B.n350 163.367
R1460 B.n702 B.n344 163.367
R1461 B.n710 B.n344 163.367
R1462 B.n710 B.n342 163.367
R1463 B.n714 B.n342 163.367
R1464 B.n714 B.n337 163.367
R1465 B.n723 B.n337 163.367
R1466 B.n723 B.n335 163.367
R1467 B.n727 B.n335 163.367
R1468 B.n727 B.n329 163.367
R1469 B.n735 B.n329 163.367
R1470 B.n735 B.n327 163.367
R1471 B.n739 B.n327 163.367
R1472 B.n739 B.n321 163.367
R1473 B.n747 B.n321 163.367
R1474 B.n747 B.n319 163.367
R1475 B.n751 B.n319 163.367
R1476 B.n751 B.n313 163.367
R1477 B.n759 B.n313 163.367
R1478 B.n759 B.n311 163.367
R1479 B.n764 B.n311 163.367
R1480 B.n764 B.n305 163.367
R1481 B.n772 B.n305 163.367
R1482 B.n773 B.n772 163.367
R1483 B.n773 B.n5 163.367
R1484 B.n6 B.n5 163.367
R1485 B.n7 B.n6 163.367
R1486 B.n778 B.n7 163.367
R1487 B.n778 B.n12 163.367
R1488 B.n13 B.n12 163.367
R1489 B.n14 B.n13 163.367
R1490 B.n783 B.n14 163.367
R1491 B.n783 B.n19 163.367
R1492 B.n20 B.n19 163.367
R1493 B.n21 B.n20 163.367
R1494 B.n788 B.n21 163.367
R1495 B.n788 B.n26 163.367
R1496 B.n27 B.n26 163.367
R1497 B.n28 B.n27 163.367
R1498 B.n793 B.n28 163.367
R1499 B.n793 B.n33 163.367
R1500 B.n34 B.n33 163.367
R1501 B.n35 B.n34 163.367
R1502 B.n798 B.n35 163.367
R1503 B.n798 B.n40 163.367
R1504 B.n41 B.n40 163.367
R1505 B.n42 B.n41 163.367
R1506 B.n803 B.n42 163.367
R1507 B.n803 B.n47 163.367
R1508 B.n48 B.n47 163.367
R1509 B.n49 B.n48 163.367
R1510 B.n808 B.n49 163.367
R1511 B.n808 B.n54 163.367
R1512 B.n55 B.n54 163.367
R1513 B.n56 B.n55 163.367
R1514 B.n813 B.n56 163.367
R1515 B.n813 B.n61 163.367
R1516 B.n62 B.n61 163.367
R1517 B.n63 B.n62 163.367
R1518 B.n818 B.n63 163.367
R1519 B.n818 B.n68 163.367
R1520 B.n69 B.n68 163.367
R1521 B.n70 B.n69 163.367
R1522 B.n823 B.n70 163.367
R1523 B.n823 B.n75 163.367
R1524 B.n76 B.n75 163.367
R1525 B.n77 B.n76 163.367
R1526 B.n828 B.n77 163.367
R1527 B.n828 B.n82 163.367
R1528 B.n83 B.n82 163.367
R1529 B.n84 B.n83 163.367
R1530 B.n833 B.n84 163.367
R1531 B.n833 B.n89 163.367
R1532 B.n90 B.n89 163.367
R1533 B.n91 B.n90 163.367
R1534 B.n838 B.n91 163.367
R1535 B.n838 B.n96 163.367
R1536 B.n97 B.n96 163.367
R1537 B.n148 B.n147 163.367
R1538 B.n152 B.n151 163.367
R1539 B.n156 B.n155 163.367
R1540 B.n160 B.n159 163.367
R1541 B.n164 B.n163 163.367
R1542 B.n168 B.n167 163.367
R1543 B.n172 B.n171 163.367
R1544 B.n176 B.n175 163.367
R1545 B.n180 B.n179 163.367
R1546 B.n184 B.n183 163.367
R1547 B.n188 B.n187 163.367
R1548 B.n192 B.n191 163.367
R1549 B.n196 B.n195 163.367
R1550 B.n200 B.n199 163.367
R1551 B.n204 B.n203 163.367
R1552 B.n208 B.n207 163.367
R1553 B.n212 B.n211 163.367
R1554 B.n216 B.n215 163.367
R1555 B.n220 B.n219 163.367
R1556 B.n224 B.n223 163.367
R1557 B.n228 B.n227 163.367
R1558 B.n232 B.n231 163.367
R1559 B.n237 B.n236 163.367
R1560 B.n241 B.n240 163.367
R1561 B.n245 B.n244 163.367
R1562 B.n249 B.n248 163.367
R1563 B.n253 B.n252 163.367
R1564 B.n257 B.n256 163.367
R1565 B.n261 B.n260 163.367
R1566 B.n265 B.n264 163.367
R1567 B.n269 B.n268 163.367
R1568 B.n273 B.n272 163.367
R1569 B.n277 B.n276 163.367
R1570 B.n281 B.n280 163.367
R1571 B.n285 B.n284 163.367
R1572 B.n289 B.n288 163.367
R1573 B.n293 B.n292 163.367
R1574 B.n297 B.n296 163.367
R1575 B.n301 B.n300 163.367
R1576 B.n843 B.n138 163.367
R1577 B.n612 B.n405 80.3559
R1578 B.n845 B.n844 80.3559
R1579 B.n452 B.n451 73.6975
R1580 B.n450 B.n449 73.6975
R1581 B.n142 B.n141 73.6975
R1582 B.n140 B.n139 73.6975
R1583 B.n611 B.n610 71.676
R1584 B.n605 B.n409 71.676
R1585 B.n602 B.n410 71.676
R1586 B.n598 B.n411 71.676
R1587 B.n594 B.n412 71.676
R1588 B.n590 B.n413 71.676
R1589 B.n586 B.n414 71.676
R1590 B.n582 B.n415 71.676
R1591 B.n578 B.n416 71.676
R1592 B.n574 B.n417 71.676
R1593 B.n570 B.n418 71.676
R1594 B.n566 B.n419 71.676
R1595 B.n562 B.n420 71.676
R1596 B.n558 B.n421 71.676
R1597 B.n554 B.n422 71.676
R1598 B.n550 B.n423 71.676
R1599 B.n546 B.n424 71.676
R1600 B.n542 B.n425 71.676
R1601 B.n537 B.n426 71.676
R1602 B.n533 B.n427 71.676
R1603 B.n529 B.n428 71.676
R1604 B.n525 B.n429 71.676
R1605 B.n521 B.n430 71.676
R1606 B.n517 B.n431 71.676
R1607 B.n513 B.n432 71.676
R1608 B.n509 B.n433 71.676
R1609 B.n505 B.n434 71.676
R1610 B.n501 B.n435 71.676
R1611 B.n497 B.n436 71.676
R1612 B.n493 B.n437 71.676
R1613 B.n489 B.n438 71.676
R1614 B.n485 B.n439 71.676
R1615 B.n481 B.n440 71.676
R1616 B.n477 B.n441 71.676
R1617 B.n473 B.n442 71.676
R1618 B.n469 B.n443 71.676
R1619 B.n465 B.n444 71.676
R1620 B.n461 B.n445 71.676
R1621 B.n457 B.n446 71.676
R1622 B.n613 B.n408 71.676
R1623 B.n144 B.n98 71.676
R1624 B.n148 B.n99 71.676
R1625 B.n152 B.n100 71.676
R1626 B.n156 B.n101 71.676
R1627 B.n160 B.n102 71.676
R1628 B.n164 B.n103 71.676
R1629 B.n168 B.n104 71.676
R1630 B.n172 B.n105 71.676
R1631 B.n176 B.n106 71.676
R1632 B.n180 B.n107 71.676
R1633 B.n184 B.n108 71.676
R1634 B.n188 B.n109 71.676
R1635 B.n192 B.n110 71.676
R1636 B.n196 B.n111 71.676
R1637 B.n200 B.n112 71.676
R1638 B.n204 B.n113 71.676
R1639 B.n208 B.n114 71.676
R1640 B.n212 B.n115 71.676
R1641 B.n216 B.n116 71.676
R1642 B.n220 B.n117 71.676
R1643 B.n224 B.n118 71.676
R1644 B.n228 B.n119 71.676
R1645 B.n232 B.n120 71.676
R1646 B.n237 B.n121 71.676
R1647 B.n241 B.n122 71.676
R1648 B.n245 B.n123 71.676
R1649 B.n249 B.n124 71.676
R1650 B.n253 B.n125 71.676
R1651 B.n257 B.n126 71.676
R1652 B.n261 B.n127 71.676
R1653 B.n265 B.n128 71.676
R1654 B.n269 B.n129 71.676
R1655 B.n273 B.n130 71.676
R1656 B.n277 B.n131 71.676
R1657 B.n281 B.n132 71.676
R1658 B.n285 B.n133 71.676
R1659 B.n289 B.n134 71.676
R1660 B.n293 B.n135 71.676
R1661 B.n297 B.n136 71.676
R1662 B.n301 B.n137 71.676
R1663 B.n138 B.n137 71.676
R1664 B.n300 B.n136 71.676
R1665 B.n296 B.n135 71.676
R1666 B.n292 B.n134 71.676
R1667 B.n288 B.n133 71.676
R1668 B.n284 B.n132 71.676
R1669 B.n280 B.n131 71.676
R1670 B.n276 B.n130 71.676
R1671 B.n272 B.n129 71.676
R1672 B.n268 B.n128 71.676
R1673 B.n264 B.n127 71.676
R1674 B.n260 B.n126 71.676
R1675 B.n256 B.n125 71.676
R1676 B.n252 B.n124 71.676
R1677 B.n248 B.n123 71.676
R1678 B.n244 B.n122 71.676
R1679 B.n240 B.n121 71.676
R1680 B.n236 B.n120 71.676
R1681 B.n231 B.n119 71.676
R1682 B.n227 B.n118 71.676
R1683 B.n223 B.n117 71.676
R1684 B.n219 B.n116 71.676
R1685 B.n215 B.n115 71.676
R1686 B.n211 B.n114 71.676
R1687 B.n207 B.n113 71.676
R1688 B.n203 B.n112 71.676
R1689 B.n199 B.n111 71.676
R1690 B.n195 B.n110 71.676
R1691 B.n191 B.n109 71.676
R1692 B.n187 B.n108 71.676
R1693 B.n183 B.n107 71.676
R1694 B.n179 B.n106 71.676
R1695 B.n175 B.n105 71.676
R1696 B.n171 B.n104 71.676
R1697 B.n167 B.n103 71.676
R1698 B.n163 B.n102 71.676
R1699 B.n159 B.n101 71.676
R1700 B.n155 B.n100 71.676
R1701 B.n151 B.n99 71.676
R1702 B.n147 B.n98 71.676
R1703 B.n611 B.n448 71.676
R1704 B.n603 B.n409 71.676
R1705 B.n599 B.n410 71.676
R1706 B.n595 B.n411 71.676
R1707 B.n591 B.n412 71.676
R1708 B.n587 B.n413 71.676
R1709 B.n583 B.n414 71.676
R1710 B.n579 B.n415 71.676
R1711 B.n575 B.n416 71.676
R1712 B.n571 B.n417 71.676
R1713 B.n567 B.n418 71.676
R1714 B.n563 B.n419 71.676
R1715 B.n559 B.n420 71.676
R1716 B.n555 B.n421 71.676
R1717 B.n551 B.n422 71.676
R1718 B.n547 B.n423 71.676
R1719 B.n543 B.n424 71.676
R1720 B.n538 B.n425 71.676
R1721 B.n534 B.n426 71.676
R1722 B.n530 B.n427 71.676
R1723 B.n526 B.n428 71.676
R1724 B.n522 B.n429 71.676
R1725 B.n518 B.n430 71.676
R1726 B.n514 B.n431 71.676
R1727 B.n510 B.n432 71.676
R1728 B.n506 B.n433 71.676
R1729 B.n502 B.n434 71.676
R1730 B.n498 B.n435 71.676
R1731 B.n494 B.n436 71.676
R1732 B.n490 B.n437 71.676
R1733 B.n486 B.n438 71.676
R1734 B.n482 B.n439 71.676
R1735 B.n478 B.n440 71.676
R1736 B.n474 B.n441 71.676
R1737 B.n470 B.n442 71.676
R1738 B.n466 B.n443 71.676
R1739 B.n462 B.n444 71.676
R1740 B.n458 B.n445 71.676
R1741 B.n454 B.n446 71.676
R1742 B.n614 B.n613 71.676
R1743 B.n453 B.n452 59.5399
R1744 B.n540 B.n450 59.5399
R1745 B.n143 B.n142 59.5399
R1746 B.n234 B.n140 59.5399
R1747 B.n619 B.n405 49.2272
R1748 B.n619 B.n401 49.2272
R1749 B.n625 B.n401 49.2272
R1750 B.n625 B.n397 49.2272
R1751 B.n631 B.n397 49.2272
R1752 B.n631 B.n393 49.2272
R1753 B.n637 B.n393 49.2272
R1754 B.n637 B.n389 49.2272
R1755 B.n643 B.n389 49.2272
R1756 B.n649 B.n385 49.2272
R1757 B.n649 B.n381 49.2272
R1758 B.n655 B.n381 49.2272
R1759 B.n655 B.n377 49.2272
R1760 B.n661 B.n377 49.2272
R1761 B.n661 B.n373 49.2272
R1762 B.n667 B.n373 49.2272
R1763 B.n667 B.n369 49.2272
R1764 B.n673 B.n369 49.2272
R1765 B.n673 B.n365 49.2272
R1766 B.n679 B.n365 49.2272
R1767 B.n679 B.n361 49.2272
R1768 B.n685 B.n361 49.2272
R1769 B.n691 B.n357 49.2272
R1770 B.n691 B.n353 49.2272
R1771 B.n697 B.n353 49.2272
R1772 B.n697 B.n349 49.2272
R1773 B.n703 B.n349 49.2272
R1774 B.n703 B.n345 49.2272
R1775 B.n709 B.n345 49.2272
R1776 B.n709 B.n341 49.2272
R1777 B.n716 B.n341 49.2272
R1778 B.n716 B.n715 49.2272
R1779 B.n722 B.n334 49.2272
R1780 B.n728 B.n334 49.2272
R1781 B.n728 B.n330 49.2272
R1782 B.n734 B.n330 49.2272
R1783 B.n734 B.n326 49.2272
R1784 B.n740 B.n326 49.2272
R1785 B.n740 B.n322 49.2272
R1786 B.n746 B.n322 49.2272
R1787 B.n746 B.n318 49.2272
R1788 B.n752 B.n318 49.2272
R1789 B.n758 B.n314 49.2272
R1790 B.n758 B.n310 49.2272
R1791 B.n765 B.n310 49.2272
R1792 B.n765 B.n306 49.2272
R1793 B.n771 B.n306 49.2272
R1794 B.n771 B.n4 49.2272
R1795 B.n950 B.n4 49.2272
R1796 B.n950 B.n949 49.2272
R1797 B.n949 B.n948 49.2272
R1798 B.n948 B.n8 49.2272
R1799 B.n942 B.n8 49.2272
R1800 B.n942 B.n941 49.2272
R1801 B.n941 B.n940 49.2272
R1802 B.n940 B.n15 49.2272
R1803 B.n934 B.n933 49.2272
R1804 B.n933 B.n932 49.2272
R1805 B.n932 B.n22 49.2272
R1806 B.n926 B.n22 49.2272
R1807 B.n926 B.n925 49.2272
R1808 B.n925 B.n924 49.2272
R1809 B.n924 B.n29 49.2272
R1810 B.n918 B.n29 49.2272
R1811 B.n918 B.n917 49.2272
R1812 B.n917 B.n916 49.2272
R1813 B.n910 B.n39 49.2272
R1814 B.n910 B.n909 49.2272
R1815 B.n909 B.n908 49.2272
R1816 B.n908 B.n43 49.2272
R1817 B.n902 B.n43 49.2272
R1818 B.n902 B.n901 49.2272
R1819 B.n901 B.n900 49.2272
R1820 B.n900 B.n50 49.2272
R1821 B.n894 B.n50 49.2272
R1822 B.n894 B.n893 49.2272
R1823 B.n892 B.n57 49.2272
R1824 B.n886 B.n57 49.2272
R1825 B.n886 B.n885 49.2272
R1826 B.n885 B.n884 49.2272
R1827 B.n884 B.n64 49.2272
R1828 B.n878 B.n64 49.2272
R1829 B.n878 B.n877 49.2272
R1830 B.n877 B.n876 49.2272
R1831 B.n876 B.n71 49.2272
R1832 B.n870 B.n71 49.2272
R1833 B.n870 B.n869 49.2272
R1834 B.n869 B.n868 49.2272
R1835 B.n868 B.n78 49.2272
R1836 B.n862 B.n861 49.2272
R1837 B.n861 B.n860 49.2272
R1838 B.n860 B.n85 49.2272
R1839 B.n854 B.n85 49.2272
R1840 B.n854 B.n853 49.2272
R1841 B.n853 B.n852 49.2272
R1842 B.n852 B.n92 49.2272
R1843 B.n846 B.n92 49.2272
R1844 B.n846 B.n845 49.2272
R1845 B.t10 B.n385 45.6076
R1846 B.t6 B.n78 45.6076
R1847 B.n752 B.t0 39.8162
R1848 B.n934 B.t4 39.8162
R1849 B.n715 B.t1 31.1292
R1850 B.n39 B.t2 31.1292
R1851 B.n145 B.n94 28.2542
R1852 B.n842 B.n841 28.2542
R1853 B.n616 B.n615 28.2542
R1854 B.n609 B.n403 28.2542
R1855 B.t3 B.n357 26.7856
R1856 B.n893 B.t19 26.7856
R1857 B.n685 B.t3 22.4421
R1858 B.t19 B.n892 22.4421
R1859 B.n722 B.t1 18.0986
R1860 B.n916 B.t2 18.0986
R1861 B B.n952 18.0485
R1862 B.n146 B.n145 10.6151
R1863 B.n149 B.n146 10.6151
R1864 B.n150 B.n149 10.6151
R1865 B.n153 B.n150 10.6151
R1866 B.n154 B.n153 10.6151
R1867 B.n157 B.n154 10.6151
R1868 B.n158 B.n157 10.6151
R1869 B.n161 B.n158 10.6151
R1870 B.n162 B.n161 10.6151
R1871 B.n165 B.n162 10.6151
R1872 B.n166 B.n165 10.6151
R1873 B.n169 B.n166 10.6151
R1874 B.n170 B.n169 10.6151
R1875 B.n173 B.n170 10.6151
R1876 B.n174 B.n173 10.6151
R1877 B.n177 B.n174 10.6151
R1878 B.n178 B.n177 10.6151
R1879 B.n181 B.n178 10.6151
R1880 B.n182 B.n181 10.6151
R1881 B.n185 B.n182 10.6151
R1882 B.n186 B.n185 10.6151
R1883 B.n189 B.n186 10.6151
R1884 B.n190 B.n189 10.6151
R1885 B.n193 B.n190 10.6151
R1886 B.n194 B.n193 10.6151
R1887 B.n197 B.n194 10.6151
R1888 B.n198 B.n197 10.6151
R1889 B.n201 B.n198 10.6151
R1890 B.n202 B.n201 10.6151
R1891 B.n205 B.n202 10.6151
R1892 B.n206 B.n205 10.6151
R1893 B.n209 B.n206 10.6151
R1894 B.n210 B.n209 10.6151
R1895 B.n213 B.n210 10.6151
R1896 B.n214 B.n213 10.6151
R1897 B.n218 B.n217 10.6151
R1898 B.n221 B.n218 10.6151
R1899 B.n222 B.n221 10.6151
R1900 B.n225 B.n222 10.6151
R1901 B.n226 B.n225 10.6151
R1902 B.n229 B.n226 10.6151
R1903 B.n230 B.n229 10.6151
R1904 B.n233 B.n230 10.6151
R1905 B.n238 B.n235 10.6151
R1906 B.n239 B.n238 10.6151
R1907 B.n242 B.n239 10.6151
R1908 B.n243 B.n242 10.6151
R1909 B.n246 B.n243 10.6151
R1910 B.n247 B.n246 10.6151
R1911 B.n250 B.n247 10.6151
R1912 B.n251 B.n250 10.6151
R1913 B.n254 B.n251 10.6151
R1914 B.n255 B.n254 10.6151
R1915 B.n258 B.n255 10.6151
R1916 B.n259 B.n258 10.6151
R1917 B.n262 B.n259 10.6151
R1918 B.n263 B.n262 10.6151
R1919 B.n266 B.n263 10.6151
R1920 B.n267 B.n266 10.6151
R1921 B.n270 B.n267 10.6151
R1922 B.n271 B.n270 10.6151
R1923 B.n274 B.n271 10.6151
R1924 B.n275 B.n274 10.6151
R1925 B.n278 B.n275 10.6151
R1926 B.n279 B.n278 10.6151
R1927 B.n282 B.n279 10.6151
R1928 B.n283 B.n282 10.6151
R1929 B.n286 B.n283 10.6151
R1930 B.n287 B.n286 10.6151
R1931 B.n290 B.n287 10.6151
R1932 B.n291 B.n290 10.6151
R1933 B.n294 B.n291 10.6151
R1934 B.n295 B.n294 10.6151
R1935 B.n298 B.n295 10.6151
R1936 B.n299 B.n298 10.6151
R1937 B.n302 B.n299 10.6151
R1938 B.n303 B.n302 10.6151
R1939 B.n842 B.n303 10.6151
R1940 B.n617 B.n616 10.6151
R1941 B.n617 B.n399 10.6151
R1942 B.n627 B.n399 10.6151
R1943 B.n628 B.n627 10.6151
R1944 B.n629 B.n628 10.6151
R1945 B.n629 B.n391 10.6151
R1946 B.n639 B.n391 10.6151
R1947 B.n640 B.n639 10.6151
R1948 B.n641 B.n640 10.6151
R1949 B.n641 B.n383 10.6151
R1950 B.n651 B.n383 10.6151
R1951 B.n652 B.n651 10.6151
R1952 B.n653 B.n652 10.6151
R1953 B.n653 B.n375 10.6151
R1954 B.n663 B.n375 10.6151
R1955 B.n664 B.n663 10.6151
R1956 B.n665 B.n664 10.6151
R1957 B.n665 B.n367 10.6151
R1958 B.n675 B.n367 10.6151
R1959 B.n676 B.n675 10.6151
R1960 B.n677 B.n676 10.6151
R1961 B.n677 B.n359 10.6151
R1962 B.n687 B.n359 10.6151
R1963 B.n688 B.n687 10.6151
R1964 B.n689 B.n688 10.6151
R1965 B.n689 B.n351 10.6151
R1966 B.n699 B.n351 10.6151
R1967 B.n700 B.n699 10.6151
R1968 B.n701 B.n700 10.6151
R1969 B.n701 B.n343 10.6151
R1970 B.n711 B.n343 10.6151
R1971 B.n712 B.n711 10.6151
R1972 B.n713 B.n712 10.6151
R1973 B.n713 B.n336 10.6151
R1974 B.n724 B.n336 10.6151
R1975 B.n725 B.n724 10.6151
R1976 B.n726 B.n725 10.6151
R1977 B.n726 B.n328 10.6151
R1978 B.n736 B.n328 10.6151
R1979 B.n737 B.n736 10.6151
R1980 B.n738 B.n737 10.6151
R1981 B.n738 B.n320 10.6151
R1982 B.n748 B.n320 10.6151
R1983 B.n749 B.n748 10.6151
R1984 B.n750 B.n749 10.6151
R1985 B.n750 B.n312 10.6151
R1986 B.n760 B.n312 10.6151
R1987 B.n761 B.n760 10.6151
R1988 B.n763 B.n761 10.6151
R1989 B.n763 B.n762 10.6151
R1990 B.n762 B.n304 10.6151
R1991 B.n774 B.n304 10.6151
R1992 B.n775 B.n774 10.6151
R1993 B.n776 B.n775 10.6151
R1994 B.n777 B.n776 10.6151
R1995 B.n779 B.n777 10.6151
R1996 B.n780 B.n779 10.6151
R1997 B.n781 B.n780 10.6151
R1998 B.n782 B.n781 10.6151
R1999 B.n784 B.n782 10.6151
R2000 B.n785 B.n784 10.6151
R2001 B.n786 B.n785 10.6151
R2002 B.n787 B.n786 10.6151
R2003 B.n789 B.n787 10.6151
R2004 B.n790 B.n789 10.6151
R2005 B.n791 B.n790 10.6151
R2006 B.n792 B.n791 10.6151
R2007 B.n794 B.n792 10.6151
R2008 B.n795 B.n794 10.6151
R2009 B.n796 B.n795 10.6151
R2010 B.n797 B.n796 10.6151
R2011 B.n799 B.n797 10.6151
R2012 B.n800 B.n799 10.6151
R2013 B.n801 B.n800 10.6151
R2014 B.n802 B.n801 10.6151
R2015 B.n804 B.n802 10.6151
R2016 B.n805 B.n804 10.6151
R2017 B.n806 B.n805 10.6151
R2018 B.n807 B.n806 10.6151
R2019 B.n809 B.n807 10.6151
R2020 B.n810 B.n809 10.6151
R2021 B.n811 B.n810 10.6151
R2022 B.n812 B.n811 10.6151
R2023 B.n814 B.n812 10.6151
R2024 B.n815 B.n814 10.6151
R2025 B.n816 B.n815 10.6151
R2026 B.n817 B.n816 10.6151
R2027 B.n819 B.n817 10.6151
R2028 B.n820 B.n819 10.6151
R2029 B.n821 B.n820 10.6151
R2030 B.n822 B.n821 10.6151
R2031 B.n824 B.n822 10.6151
R2032 B.n825 B.n824 10.6151
R2033 B.n826 B.n825 10.6151
R2034 B.n827 B.n826 10.6151
R2035 B.n829 B.n827 10.6151
R2036 B.n830 B.n829 10.6151
R2037 B.n831 B.n830 10.6151
R2038 B.n832 B.n831 10.6151
R2039 B.n834 B.n832 10.6151
R2040 B.n835 B.n834 10.6151
R2041 B.n836 B.n835 10.6151
R2042 B.n837 B.n836 10.6151
R2043 B.n839 B.n837 10.6151
R2044 B.n840 B.n839 10.6151
R2045 B.n841 B.n840 10.6151
R2046 B.n609 B.n608 10.6151
R2047 B.n608 B.n607 10.6151
R2048 B.n607 B.n606 10.6151
R2049 B.n606 B.n604 10.6151
R2050 B.n604 B.n601 10.6151
R2051 B.n601 B.n600 10.6151
R2052 B.n600 B.n597 10.6151
R2053 B.n597 B.n596 10.6151
R2054 B.n596 B.n593 10.6151
R2055 B.n593 B.n592 10.6151
R2056 B.n592 B.n589 10.6151
R2057 B.n589 B.n588 10.6151
R2058 B.n588 B.n585 10.6151
R2059 B.n585 B.n584 10.6151
R2060 B.n584 B.n581 10.6151
R2061 B.n581 B.n580 10.6151
R2062 B.n580 B.n577 10.6151
R2063 B.n577 B.n576 10.6151
R2064 B.n576 B.n573 10.6151
R2065 B.n573 B.n572 10.6151
R2066 B.n572 B.n569 10.6151
R2067 B.n569 B.n568 10.6151
R2068 B.n568 B.n565 10.6151
R2069 B.n565 B.n564 10.6151
R2070 B.n564 B.n561 10.6151
R2071 B.n561 B.n560 10.6151
R2072 B.n560 B.n557 10.6151
R2073 B.n557 B.n556 10.6151
R2074 B.n556 B.n553 10.6151
R2075 B.n553 B.n552 10.6151
R2076 B.n552 B.n549 10.6151
R2077 B.n549 B.n548 10.6151
R2078 B.n548 B.n545 10.6151
R2079 B.n545 B.n544 10.6151
R2080 B.n544 B.n541 10.6151
R2081 B.n539 B.n536 10.6151
R2082 B.n536 B.n535 10.6151
R2083 B.n535 B.n532 10.6151
R2084 B.n532 B.n531 10.6151
R2085 B.n531 B.n528 10.6151
R2086 B.n528 B.n527 10.6151
R2087 B.n527 B.n524 10.6151
R2088 B.n524 B.n523 10.6151
R2089 B.n520 B.n519 10.6151
R2090 B.n519 B.n516 10.6151
R2091 B.n516 B.n515 10.6151
R2092 B.n515 B.n512 10.6151
R2093 B.n512 B.n511 10.6151
R2094 B.n511 B.n508 10.6151
R2095 B.n508 B.n507 10.6151
R2096 B.n507 B.n504 10.6151
R2097 B.n504 B.n503 10.6151
R2098 B.n503 B.n500 10.6151
R2099 B.n500 B.n499 10.6151
R2100 B.n499 B.n496 10.6151
R2101 B.n496 B.n495 10.6151
R2102 B.n495 B.n492 10.6151
R2103 B.n492 B.n491 10.6151
R2104 B.n491 B.n488 10.6151
R2105 B.n488 B.n487 10.6151
R2106 B.n487 B.n484 10.6151
R2107 B.n484 B.n483 10.6151
R2108 B.n483 B.n480 10.6151
R2109 B.n480 B.n479 10.6151
R2110 B.n479 B.n476 10.6151
R2111 B.n476 B.n475 10.6151
R2112 B.n475 B.n472 10.6151
R2113 B.n472 B.n471 10.6151
R2114 B.n471 B.n468 10.6151
R2115 B.n468 B.n467 10.6151
R2116 B.n467 B.n464 10.6151
R2117 B.n464 B.n463 10.6151
R2118 B.n463 B.n460 10.6151
R2119 B.n460 B.n459 10.6151
R2120 B.n459 B.n456 10.6151
R2121 B.n456 B.n455 10.6151
R2122 B.n455 B.n407 10.6151
R2123 B.n615 B.n407 10.6151
R2124 B.n621 B.n403 10.6151
R2125 B.n622 B.n621 10.6151
R2126 B.n623 B.n622 10.6151
R2127 B.n623 B.n395 10.6151
R2128 B.n633 B.n395 10.6151
R2129 B.n634 B.n633 10.6151
R2130 B.n635 B.n634 10.6151
R2131 B.n635 B.n387 10.6151
R2132 B.n645 B.n387 10.6151
R2133 B.n646 B.n645 10.6151
R2134 B.n647 B.n646 10.6151
R2135 B.n647 B.n379 10.6151
R2136 B.n657 B.n379 10.6151
R2137 B.n658 B.n657 10.6151
R2138 B.n659 B.n658 10.6151
R2139 B.n659 B.n371 10.6151
R2140 B.n669 B.n371 10.6151
R2141 B.n670 B.n669 10.6151
R2142 B.n671 B.n670 10.6151
R2143 B.n671 B.n363 10.6151
R2144 B.n681 B.n363 10.6151
R2145 B.n682 B.n681 10.6151
R2146 B.n683 B.n682 10.6151
R2147 B.n683 B.n355 10.6151
R2148 B.n693 B.n355 10.6151
R2149 B.n694 B.n693 10.6151
R2150 B.n695 B.n694 10.6151
R2151 B.n695 B.n347 10.6151
R2152 B.n705 B.n347 10.6151
R2153 B.n706 B.n705 10.6151
R2154 B.n707 B.n706 10.6151
R2155 B.n707 B.n339 10.6151
R2156 B.n718 B.n339 10.6151
R2157 B.n719 B.n718 10.6151
R2158 B.n720 B.n719 10.6151
R2159 B.n720 B.n332 10.6151
R2160 B.n730 B.n332 10.6151
R2161 B.n731 B.n730 10.6151
R2162 B.n732 B.n731 10.6151
R2163 B.n732 B.n324 10.6151
R2164 B.n742 B.n324 10.6151
R2165 B.n743 B.n742 10.6151
R2166 B.n744 B.n743 10.6151
R2167 B.n744 B.n316 10.6151
R2168 B.n754 B.n316 10.6151
R2169 B.n755 B.n754 10.6151
R2170 B.n756 B.n755 10.6151
R2171 B.n756 B.n308 10.6151
R2172 B.n767 B.n308 10.6151
R2173 B.n768 B.n767 10.6151
R2174 B.n769 B.n768 10.6151
R2175 B.n769 B.n0 10.6151
R2176 B.n946 B.n1 10.6151
R2177 B.n946 B.n945 10.6151
R2178 B.n945 B.n944 10.6151
R2179 B.n944 B.n10 10.6151
R2180 B.n938 B.n10 10.6151
R2181 B.n938 B.n937 10.6151
R2182 B.n937 B.n936 10.6151
R2183 B.n936 B.n17 10.6151
R2184 B.n930 B.n17 10.6151
R2185 B.n930 B.n929 10.6151
R2186 B.n929 B.n928 10.6151
R2187 B.n928 B.n24 10.6151
R2188 B.n922 B.n24 10.6151
R2189 B.n922 B.n921 10.6151
R2190 B.n921 B.n920 10.6151
R2191 B.n920 B.n31 10.6151
R2192 B.n914 B.n31 10.6151
R2193 B.n914 B.n913 10.6151
R2194 B.n913 B.n912 10.6151
R2195 B.n912 B.n37 10.6151
R2196 B.n906 B.n37 10.6151
R2197 B.n906 B.n905 10.6151
R2198 B.n905 B.n904 10.6151
R2199 B.n904 B.n45 10.6151
R2200 B.n898 B.n45 10.6151
R2201 B.n898 B.n897 10.6151
R2202 B.n897 B.n896 10.6151
R2203 B.n896 B.n52 10.6151
R2204 B.n890 B.n52 10.6151
R2205 B.n890 B.n889 10.6151
R2206 B.n889 B.n888 10.6151
R2207 B.n888 B.n59 10.6151
R2208 B.n882 B.n59 10.6151
R2209 B.n882 B.n881 10.6151
R2210 B.n881 B.n880 10.6151
R2211 B.n880 B.n66 10.6151
R2212 B.n874 B.n66 10.6151
R2213 B.n874 B.n873 10.6151
R2214 B.n873 B.n872 10.6151
R2215 B.n872 B.n73 10.6151
R2216 B.n866 B.n73 10.6151
R2217 B.n866 B.n865 10.6151
R2218 B.n865 B.n864 10.6151
R2219 B.n864 B.n80 10.6151
R2220 B.n858 B.n80 10.6151
R2221 B.n858 B.n857 10.6151
R2222 B.n857 B.n856 10.6151
R2223 B.n856 B.n87 10.6151
R2224 B.n850 B.n87 10.6151
R2225 B.n850 B.n849 10.6151
R2226 B.n849 B.n848 10.6151
R2227 B.n848 B.n94 10.6151
R2228 B.t0 B.n314 9.41149
R2229 B.t4 B.n15 9.41149
R2230 B.n217 B.n143 6.5566
R2231 B.n234 B.n233 6.5566
R2232 B.n540 B.n539 6.5566
R2233 B.n523 B.n453 6.5566
R2234 B.n214 B.n143 4.05904
R2235 B.n235 B.n234 4.05904
R2236 B.n541 B.n540 4.05904
R2237 B.n520 B.n453 4.05904
R2238 B.n643 B.t10 3.62011
R2239 B.n862 B.t6 3.62011
R2240 B.n952 B.n0 2.81026
R2241 B.n952 B.n1 2.81026
R2242 VN.n34 VN.n33 161.3
R2243 VN.n32 VN.n19 161.3
R2244 VN.n31 VN.n30 161.3
R2245 VN.n29 VN.n20 161.3
R2246 VN.n28 VN.n27 161.3
R2247 VN.n26 VN.n21 161.3
R2248 VN.n25 VN.n24 161.3
R2249 VN.n16 VN.n15 161.3
R2250 VN.n14 VN.n1 161.3
R2251 VN.n13 VN.n12 161.3
R2252 VN.n11 VN.n2 161.3
R2253 VN.n10 VN.n9 161.3
R2254 VN.n8 VN.n3 161.3
R2255 VN.n7 VN.n6 161.3
R2256 VN.n23 VN.t3 103.058
R2257 VN.n5 VN.t1 103.058
R2258 VN.n17 VN.n0 75.4905
R2259 VN.n35 VN.n18 75.4905
R2260 VN.n4 VN.t5 68.8973
R2261 VN.n0 VN.t0 68.8973
R2262 VN.n22 VN.t2 68.8973
R2263 VN.n18 VN.t4 68.8973
R2264 VN VN.n35 50.8315
R2265 VN.n5 VN.n4 50.305
R2266 VN.n23 VN.n22 50.305
R2267 VN.n9 VN.n2 50.2647
R2268 VN.n27 VN.n20 50.2647
R2269 VN.n13 VN.n2 30.8893
R2270 VN.n31 VN.n20 30.8893
R2271 VN.n7 VN.n4 24.5923
R2272 VN.n8 VN.n7 24.5923
R2273 VN.n9 VN.n8 24.5923
R2274 VN.n14 VN.n13 24.5923
R2275 VN.n15 VN.n14 24.5923
R2276 VN.n27 VN.n26 24.5923
R2277 VN.n26 VN.n25 24.5923
R2278 VN.n25 VN.n22 24.5923
R2279 VN.n33 VN.n32 24.5923
R2280 VN.n32 VN.n31 24.5923
R2281 VN.n15 VN.n0 14.7556
R2282 VN.n33 VN.n18 14.7556
R2283 VN.n6 VN.n5 2.98133
R2284 VN.n24 VN.n23 2.98133
R2285 VN.n35 VN.n34 0.354861
R2286 VN.n17 VN.n16 0.354861
R2287 VN VN.n17 0.267071
R2288 VN.n34 VN.n19 0.189894
R2289 VN.n30 VN.n19 0.189894
R2290 VN.n30 VN.n29 0.189894
R2291 VN.n29 VN.n28 0.189894
R2292 VN.n28 VN.n21 0.189894
R2293 VN.n24 VN.n21 0.189894
R2294 VN.n6 VN.n3 0.189894
R2295 VN.n10 VN.n3 0.189894
R2296 VN.n11 VN.n10 0.189894
R2297 VN.n12 VN.n11 0.189894
R2298 VN.n12 VN.n1 0.189894
R2299 VN.n16 VN.n1 0.189894
R2300 VDD2.n103 VDD2.n55 289.615
R2301 VDD2.n48 VDD2.n0 289.615
R2302 VDD2.n104 VDD2.n103 185
R2303 VDD2.n102 VDD2.n101 185
R2304 VDD2.n59 VDD2.n58 185
R2305 VDD2.n96 VDD2.n95 185
R2306 VDD2.n94 VDD2.n61 185
R2307 VDD2.n93 VDD2.n92 185
R2308 VDD2.n64 VDD2.n62 185
R2309 VDD2.n87 VDD2.n86 185
R2310 VDD2.n85 VDD2.n84 185
R2311 VDD2.n68 VDD2.n67 185
R2312 VDD2.n79 VDD2.n78 185
R2313 VDD2.n77 VDD2.n76 185
R2314 VDD2.n72 VDD2.n71 185
R2315 VDD2.n16 VDD2.n15 185
R2316 VDD2.n21 VDD2.n20 185
R2317 VDD2.n23 VDD2.n22 185
R2318 VDD2.n12 VDD2.n11 185
R2319 VDD2.n29 VDD2.n28 185
R2320 VDD2.n31 VDD2.n30 185
R2321 VDD2.n8 VDD2.n7 185
R2322 VDD2.n38 VDD2.n37 185
R2323 VDD2.n39 VDD2.n6 185
R2324 VDD2.n41 VDD2.n40 185
R2325 VDD2.n4 VDD2.n3 185
R2326 VDD2.n47 VDD2.n46 185
R2327 VDD2.n49 VDD2.n48 185
R2328 VDD2.n73 VDD2.t1 149.524
R2329 VDD2.n17 VDD2.t4 149.524
R2330 VDD2.n103 VDD2.n102 104.615
R2331 VDD2.n102 VDD2.n58 104.615
R2332 VDD2.n95 VDD2.n58 104.615
R2333 VDD2.n95 VDD2.n94 104.615
R2334 VDD2.n94 VDD2.n93 104.615
R2335 VDD2.n93 VDD2.n62 104.615
R2336 VDD2.n86 VDD2.n62 104.615
R2337 VDD2.n86 VDD2.n85 104.615
R2338 VDD2.n85 VDD2.n67 104.615
R2339 VDD2.n78 VDD2.n67 104.615
R2340 VDD2.n78 VDD2.n77 104.615
R2341 VDD2.n77 VDD2.n71 104.615
R2342 VDD2.n21 VDD2.n15 104.615
R2343 VDD2.n22 VDD2.n21 104.615
R2344 VDD2.n22 VDD2.n11 104.615
R2345 VDD2.n29 VDD2.n11 104.615
R2346 VDD2.n30 VDD2.n29 104.615
R2347 VDD2.n30 VDD2.n7 104.615
R2348 VDD2.n38 VDD2.n7 104.615
R2349 VDD2.n39 VDD2.n38 104.615
R2350 VDD2.n40 VDD2.n39 104.615
R2351 VDD2.n40 VDD2.n3 104.615
R2352 VDD2.n47 VDD2.n3 104.615
R2353 VDD2.n48 VDD2.n47 104.615
R2354 VDD2.n54 VDD2.n53 62.628
R2355 VDD2 VDD2.n109 62.6252
R2356 VDD2.t1 VDD2.n71 52.3082
R2357 VDD2.t4 VDD2.n15 52.3082
R2358 VDD2.n54 VDD2.n52 50.4899
R2359 VDD2.n108 VDD2.n107 48.0884
R2360 VDD2.n108 VDD2.n54 42.9136
R2361 VDD2.n96 VDD2.n61 13.1884
R2362 VDD2.n41 VDD2.n6 13.1884
R2363 VDD2.n97 VDD2.n59 12.8005
R2364 VDD2.n92 VDD2.n63 12.8005
R2365 VDD2.n37 VDD2.n36 12.8005
R2366 VDD2.n42 VDD2.n4 12.8005
R2367 VDD2.n101 VDD2.n100 12.0247
R2368 VDD2.n91 VDD2.n64 12.0247
R2369 VDD2.n35 VDD2.n8 12.0247
R2370 VDD2.n46 VDD2.n45 12.0247
R2371 VDD2.n104 VDD2.n57 11.249
R2372 VDD2.n88 VDD2.n87 11.249
R2373 VDD2.n32 VDD2.n31 11.249
R2374 VDD2.n49 VDD2.n2 11.249
R2375 VDD2.n105 VDD2.n55 10.4732
R2376 VDD2.n84 VDD2.n66 10.4732
R2377 VDD2.n28 VDD2.n10 10.4732
R2378 VDD2.n50 VDD2.n0 10.4732
R2379 VDD2.n73 VDD2.n72 10.2747
R2380 VDD2.n17 VDD2.n16 10.2747
R2381 VDD2.n83 VDD2.n68 9.69747
R2382 VDD2.n27 VDD2.n12 9.69747
R2383 VDD2.n107 VDD2.n106 9.45567
R2384 VDD2.n52 VDD2.n51 9.45567
R2385 VDD2.n75 VDD2.n74 9.3005
R2386 VDD2.n70 VDD2.n69 9.3005
R2387 VDD2.n81 VDD2.n80 9.3005
R2388 VDD2.n83 VDD2.n82 9.3005
R2389 VDD2.n66 VDD2.n65 9.3005
R2390 VDD2.n89 VDD2.n88 9.3005
R2391 VDD2.n91 VDD2.n90 9.3005
R2392 VDD2.n63 VDD2.n60 9.3005
R2393 VDD2.n106 VDD2.n105 9.3005
R2394 VDD2.n57 VDD2.n56 9.3005
R2395 VDD2.n100 VDD2.n99 9.3005
R2396 VDD2.n98 VDD2.n97 9.3005
R2397 VDD2.n51 VDD2.n50 9.3005
R2398 VDD2.n2 VDD2.n1 9.3005
R2399 VDD2.n45 VDD2.n44 9.3005
R2400 VDD2.n43 VDD2.n42 9.3005
R2401 VDD2.n19 VDD2.n18 9.3005
R2402 VDD2.n14 VDD2.n13 9.3005
R2403 VDD2.n25 VDD2.n24 9.3005
R2404 VDD2.n27 VDD2.n26 9.3005
R2405 VDD2.n10 VDD2.n9 9.3005
R2406 VDD2.n33 VDD2.n32 9.3005
R2407 VDD2.n35 VDD2.n34 9.3005
R2408 VDD2.n36 VDD2.n5 9.3005
R2409 VDD2.n80 VDD2.n79 8.92171
R2410 VDD2.n24 VDD2.n23 8.92171
R2411 VDD2.n76 VDD2.n70 8.14595
R2412 VDD2.n20 VDD2.n14 8.14595
R2413 VDD2.n75 VDD2.n72 7.3702
R2414 VDD2.n19 VDD2.n16 7.3702
R2415 VDD2.n76 VDD2.n75 5.81868
R2416 VDD2.n20 VDD2.n19 5.81868
R2417 VDD2.n79 VDD2.n70 5.04292
R2418 VDD2.n23 VDD2.n14 5.04292
R2419 VDD2.n80 VDD2.n68 4.26717
R2420 VDD2.n24 VDD2.n12 4.26717
R2421 VDD2.n107 VDD2.n55 3.49141
R2422 VDD2.n84 VDD2.n83 3.49141
R2423 VDD2.n28 VDD2.n27 3.49141
R2424 VDD2.n52 VDD2.n0 3.49141
R2425 VDD2.n74 VDD2.n73 2.84303
R2426 VDD2.n18 VDD2.n17 2.84303
R2427 VDD2.n105 VDD2.n104 2.71565
R2428 VDD2.n87 VDD2.n66 2.71565
R2429 VDD2.n31 VDD2.n10 2.71565
R2430 VDD2.n50 VDD2.n49 2.71565
R2431 VDD2 VDD2.n108 2.51559
R2432 VDD2.n109 VDD2.t3 1.99647
R2433 VDD2.n109 VDD2.t2 1.99647
R2434 VDD2.n53 VDD2.t0 1.99647
R2435 VDD2.n53 VDD2.t5 1.99647
R2436 VDD2.n101 VDD2.n57 1.93989
R2437 VDD2.n88 VDD2.n64 1.93989
R2438 VDD2.n32 VDD2.n8 1.93989
R2439 VDD2.n46 VDD2.n2 1.93989
R2440 VDD2.n100 VDD2.n59 1.16414
R2441 VDD2.n92 VDD2.n91 1.16414
R2442 VDD2.n37 VDD2.n35 1.16414
R2443 VDD2.n45 VDD2.n4 1.16414
R2444 VDD2.n97 VDD2.n96 0.388379
R2445 VDD2.n63 VDD2.n61 0.388379
R2446 VDD2.n36 VDD2.n6 0.388379
R2447 VDD2.n42 VDD2.n41 0.388379
R2448 VDD2.n106 VDD2.n56 0.155672
R2449 VDD2.n99 VDD2.n56 0.155672
R2450 VDD2.n99 VDD2.n98 0.155672
R2451 VDD2.n98 VDD2.n60 0.155672
R2452 VDD2.n90 VDD2.n60 0.155672
R2453 VDD2.n90 VDD2.n89 0.155672
R2454 VDD2.n89 VDD2.n65 0.155672
R2455 VDD2.n82 VDD2.n65 0.155672
R2456 VDD2.n82 VDD2.n81 0.155672
R2457 VDD2.n81 VDD2.n69 0.155672
R2458 VDD2.n74 VDD2.n69 0.155672
R2459 VDD2.n18 VDD2.n13 0.155672
R2460 VDD2.n25 VDD2.n13 0.155672
R2461 VDD2.n26 VDD2.n25 0.155672
R2462 VDD2.n26 VDD2.n9 0.155672
R2463 VDD2.n33 VDD2.n9 0.155672
R2464 VDD2.n34 VDD2.n33 0.155672
R2465 VDD2.n34 VDD2.n5 0.155672
R2466 VDD2.n43 VDD2.n5 0.155672
R2467 VDD2.n44 VDD2.n43 0.155672
R2468 VDD2.n44 VDD2.n1 0.155672
R2469 VDD2.n51 VDD2.n1 0.155672
C0 VDD1 VDD2 1.74601f
C1 VN VDD2 5.90266f
C2 VDD1 VP 6.27992f
C3 VP VN 7.37932f
C4 VDD1 VN 0.152232f
C5 VTAIL VDD2 7.38485f
C6 VTAIL VP 6.38343f
C7 VP VDD2 0.532269f
C8 VTAIL VDD1 7.32707f
C9 VTAIL VN 6.36922f
C10 VDD2 B 6.279733f
C11 VDD1 B 6.448449f
C12 VTAIL B 7.527582f
C13 VN B 15.284449f
C14 VP B 14.001151f
C15 VDD2.n0 B 0.0279f
C16 VDD2.n1 B 0.021501f
C17 VDD2.n2 B 0.011554f
C18 VDD2.n3 B 0.027308f
C19 VDD2.n4 B 0.012233f
C20 VDD2.n5 B 0.021501f
C21 VDD2.n6 B 0.011893f
C22 VDD2.n7 B 0.027308f
C23 VDD2.n8 B 0.012233f
C24 VDD2.n9 B 0.021501f
C25 VDD2.n10 B 0.011554f
C26 VDD2.n11 B 0.027308f
C27 VDD2.n12 B 0.012233f
C28 VDD2.n13 B 0.021501f
C29 VDD2.n14 B 0.011554f
C30 VDD2.n15 B 0.020481f
C31 VDD2.n16 B 0.019305f
C32 VDD2.t4 B 0.045882f
C33 VDD2.n17 B 0.13785f
C34 VDD2.n18 B 0.885749f
C35 VDD2.n19 B 0.011554f
C36 VDD2.n20 B 0.012233f
C37 VDD2.n21 B 0.027308f
C38 VDD2.n22 B 0.027308f
C39 VDD2.n23 B 0.012233f
C40 VDD2.n24 B 0.011554f
C41 VDD2.n25 B 0.021501f
C42 VDD2.n26 B 0.021501f
C43 VDD2.n27 B 0.011554f
C44 VDD2.n28 B 0.012233f
C45 VDD2.n29 B 0.027308f
C46 VDD2.n30 B 0.027308f
C47 VDD2.n31 B 0.012233f
C48 VDD2.n32 B 0.011554f
C49 VDD2.n33 B 0.021501f
C50 VDD2.n34 B 0.021501f
C51 VDD2.n35 B 0.011554f
C52 VDD2.n36 B 0.011554f
C53 VDD2.n37 B 0.012233f
C54 VDD2.n38 B 0.027308f
C55 VDD2.n39 B 0.027308f
C56 VDD2.n40 B 0.027308f
C57 VDD2.n41 B 0.011893f
C58 VDD2.n42 B 0.011554f
C59 VDD2.n43 B 0.021501f
C60 VDD2.n44 B 0.021501f
C61 VDD2.n45 B 0.011554f
C62 VDD2.n46 B 0.012233f
C63 VDD2.n47 B 0.027308f
C64 VDD2.n48 B 0.055013f
C65 VDD2.n49 B 0.012233f
C66 VDD2.n50 B 0.011554f
C67 VDD2.n51 B 0.048523f
C68 VDD2.n52 B 0.05504f
C69 VDD2.t0 B 0.168545f
C70 VDD2.t5 B 0.168545f
C71 VDD2.n53 B 1.48823f
C72 VDD2.n54 B 2.51342f
C73 VDD2.n55 B 0.0279f
C74 VDD2.n56 B 0.021501f
C75 VDD2.n57 B 0.011554f
C76 VDD2.n58 B 0.027308f
C77 VDD2.n59 B 0.012233f
C78 VDD2.n60 B 0.021501f
C79 VDD2.n61 B 0.011893f
C80 VDD2.n62 B 0.027308f
C81 VDD2.n63 B 0.011554f
C82 VDD2.n64 B 0.012233f
C83 VDD2.n65 B 0.021501f
C84 VDD2.n66 B 0.011554f
C85 VDD2.n67 B 0.027308f
C86 VDD2.n68 B 0.012233f
C87 VDD2.n69 B 0.021501f
C88 VDD2.n70 B 0.011554f
C89 VDD2.n71 B 0.020481f
C90 VDD2.n72 B 0.019305f
C91 VDD2.t1 B 0.045882f
C92 VDD2.n73 B 0.13785f
C93 VDD2.n74 B 0.885749f
C94 VDD2.n75 B 0.011554f
C95 VDD2.n76 B 0.012233f
C96 VDD2.n77 B 0.027308f
C97 VDD2.n78 B 0.027308f
C98 VDD2.n79 B 0.012233f
C99 VDD2.n80 B 0.011554f
C100 VDD2.n81 B 0.021501f
C101 VDD2.n82 B 0.021501f
C102 VDD2.n83 B 0.011554f
C103 VDD2.n84 B 0.012233f
C104 VDD2.n85 B 0.027308f
C105 VDD2.n86 B 0.027308f
C106 VDD2.n87 B 0.012233f
C107 VDD2.n88 B 0.011554f
C108 VDD2.n89 B 0.021501f
C109 VDD2.n90 B 0.021501f
C110 VDD2.n91 B 0.011554f
C111 VDD2.n92 B 0.012233f
C112 VDD2.n93 B 0.027308f
C113 VDD2.n94 B 0.027308f
C114 VDD2.n95 B 0.027308f
C115 VDD2.n96 B 0.011893f
C116 VDD2.n97 B 0.011554f
C117 VDD2.n98 B 0.021501f
C118 VDD2.n99 B 0.021501f
C119 VDD2.n100 B 0.011554f
C120 VDD2.n101 B 0.012233f
C121 VDD2.n102 B 0.027308f
C122 VDD2.n103 B 0.055013f
C123 VDD2.n104 B 0.012233f
C124 VDD2.n105 B 0.011554f
C125 VDD2.n106 B 0.048523f
C126 VDD2.n107 B 0.045179f
C127 VDD2.n108 B 2.26853f
C128 VDD2.t3 B 0.168545f
C129 VDD2.t2 B 0.168545f
C130 VDD2.n109 B 1.4882f
C131 VN.t0 B 1.86742f
C132 VN.n0 B 0.744427f
C133 VN.n1 B 0.020031f
C134 VN.n2 B 0.018886f
C135 VN.n3 B 0.020031f
C136 VN.t5 B 1.86742f
C137 VN.n4 B 0.741677f
C138 VN.t1 B 2.13727f
C139 VN.n5 B 0.693164f
C140 VN.n6 B 0.244399f
C141 VN.n7 B 0.037146f
C142 VN.n8 B 0.037146f
C143 VN.n9 B 0.036584f
C144 VN.n10 B 0.020031f
C145 VN.n11 B 0.020031f
C146 VN.n12 B 0.020031f
C147 VN.n13 B 0.039912f
C148 VN.n14 B 0.037146f
C149 VN.n15 B 0.029811f
C150 VN.n16 B 0.032325f
C151 VN.n17 B 0.04982f
C152 VN.t4 B 1.86742f
C153 VN.n18 B 0.744427f
C154 VN.n19 B 0.020031f
C155 VN.n20 B 0.018886f
C156 VN.n21 B 0.020031f
C157 VN.t2 B 1.86742f
C158 VN.n22 B 0.741677f
C159 VN.t3 B 2.13727f
C160 VN.n23 B 0.693164f
C161 VN.n24 B 0.244399f
C162 VN.n25 B 0.037146f
C163 VN.n26 B 0.037146f
C164 VN.n27 B 0.036584f
C165 VN.n28 B 0.020031f
C166 VN.n29 B 0.020031f
C167 VN.n30 B 0.020031f
C168 VN.n31 B 0.039912f
C169 VN.n32 B 0.037146f
C170 VN.n33 B 0.029811f
C171 VN.n34 B 0.032325f
C172 VN.n35 B 1.17205f
C173 VDD1.n0 B 0.02836f
C174 VDD1.n1 B 0.021855f
C175 VDD1.n2 B 0.011744f
C176 VDD1.n3 B 0.027758f
C177 VDD1.n4 B 0.012435f
C178 VDD1.n5 B 0.021855f
C179 VDD1.n6 B 0.012089f
C180 VDD1.n7 B 0.027758f
C181 VDD1.n8 B 0.011744f
C182 VDD1.n9 B 0.012435f
C183 VDD1.n10 B 0.021855f
C184 VDD1.n11 B 0.011744f
C185 VDD1.n12 B 0.027758f
C186 VDD1.n13 B 0.012435f
C187 VDD1.n14 B 0.021855f
C188 VDD1.n15 B 0.011744f
C189 VDD1.n16 B 0.020819f
C190 VDD1.n17 B 0.019623f
C191 VDD1.t2 B 0.046639f
C192 VDD1.n18 B 0.140122f
C193 VDD1.n19 B 0.900353f
C194 VDD1.n20 B 0.011744f
C195 VDD1.n21 B 0.012435f
C196 VDD1.n22 B 0.027758f
C197 VDD1.n23 B 0.027758f
C198 VDD1.n24 B 0.012435f
C199 VDD1.n25 B 0.011744f
C200 VDD1.n26 B 0.021855f
C201 VDD1.n27 B 0.021855f
C202 VDD1.n28 B 0.011744f
C203 VDD1.n29 B 0.012435f
C204 VDD1.n30 B 0.027758f
C205 VDD1.n31 B 0.027758f
C206 VDD1.n32 B 0.012435f
C207 VDD1.n33 B 0.011744f
C208 VDD1.n34 B 0.021855f
C209 VDD1.n35 B 0.021855f
C210 VDD1.n36 B 0.011744f
C211 VDD1.n37 B 0.012435f
C212 VDD1.n38 B 0.027758f
C213 VDD1.n39 B 0.027758f
C214 VDD1.n40 B 0.027758f
C215 VDD1.n41 B 0.012089f
C216 VDD1.n42 B 0.011744f
C217 VDD1.n43 B 0.021855f
C218 VDD1.n44 B 0.021855f
C219 VDD1.n45 B 0.011744f
C220 VDD1.n46 B 0.012435f
C221 VDD1.n47 B 0.027758f
C222 VDD1.n48 B 0.05592f
C223 VDD1.n49 B 0.012435f
C224 VDD1.n50 B 0.011744f
C225 VDD1.n51 B 0.049323f
C226 VDD1.n52 B 0.056785f
C227 VDD1.n53 B 0.02836f
C228 VDD1.n54 B 0.021855f
C229 VDD1.n55 B 0.011744f
C230 VDD1.n56 B 0.027758f
C231 VDD1.n57 B 0.012435f
C232 VDD1.n58 B 0.021855f
C233 VDD1.n59 B 0.012089f
C234 VDD1.n60 B 0.027758f
C235 VDD1.n61 B 0.012435f
C236 VDD1.n62 B 0.021855f
C237 VDD1.n63 B 0.011744f
C238 VDD1.n64 B 0.027758f
C239 VDD1.n65 B 0.012435f
C240 VDD1.n66 B 0.021855f
C241 VDD1.n67 B 0.011744f
C242 VDD1.n68 B 0.020819f
C243 VDD1.n69 B 0.019623f
C244 VDD1.t4 B 0.046639f
C245 VDD1.n70 B 0.140122f
C246 VDD1.n71 B 0.900353f
C247 VDD1.n72 B 0.011744f
C248 VDD1.n73 B 0.012435f
C249 VDD1.n74 B 0.027758f
C250 VDD1.n75 B 0.027758f
C251 VDD1.n76 B 0.012435f
C252 VDD1.n77 B 0.011744f
C253 VDD1.n78 B 0.021855f
C254 VDD1.n79 B 0.021855f
C255 VDD1.n80 B 0.011744f
C256 VDD1.n81 B 0.012435f
C257 VDD1.n82 B 0.027758f
C258 VDD1.n83 B 0.027758f
C259 VDD1.n84 B 0.012435f
C260 VDD1.n85 B 0.011744f
C261 VDD1.n86 B 0.021855f
C262 VDD1.n87 B 0.021855f
C263 VDD1.n88 B 0.011744f
C264 VDD1.n89 B 0.011744f
C265 VDD1.n90 B 0.012435f
C266 VDD1.n91 B 0.027758f
C267 VDD1.n92 B 0.027758f
C268 VDD1.n93 B 0.027758f
C269 VDD1.n94 B 0.012089f
C270 VDD1.n95 B 0.011744f
C271 VDD1.n96 B 0.021855f
C272 VDD1.n97 B 0.021855f
C273 VDD1.n98 B 0.011744f
C274 VDD1.n99 B 0.012435f
C275 VDD1.n100 B 0.027758f
C276 VDD1.n101 B 0.05592f
C277 VDD1.n102 B 0.012435f
C278 VDD1.n103 B 0.011744f
C279 VDD1.n104 B 0.049323f
C280 VDD1.n105 B 0.055947f
C281 VDD1.t1 B 0.171324f
C282 VDD1.t3 B 0.171324f
C283 VDD1.n106 B 1.51277f
C284 VDD1.n107 B 2.68181f
C285 VDD1.t0 B 0.171324f
C286 VDD1.t5 B 0.171324f
C287 VDD1.n108 B 1.50701f
C288 VDD1.n109 B 2.51302f
C289 VTAIL.t4 B 0.197064f
C290 VTAIL.t2 B 0.197064f
C291 VTAIL.n0 B 1.65929f
C292 VTAIL.n1 B 0.487387f
C293 VTAIL.n2 B 0.032621f
C294 VTAIL.n3 B 0.025139f
C295 VTAIL.n4 B 0.013508f
C296 VTAIL.n5 B 0.031929f
C297 VTAIL.n6 B 0.014303f
C298 VTAIL.n7 B 0.025139f
C299 VTAIL.n8 B 0.013906f
C300 VTAIL.n9 B 0.031929f
C301 VTAIL.n10 B 0.014303f
C302 VTAIL.n11 B 0.025139f
C303 VTAIL.n12 B 0.013508f
C304 VTAIL.n13 B 0.031929f
C305 VTAIL.n14 B 0.014303f
C306 VTAIL.n15 B 0.025139f
C307 VTAIL.n16 B 0.013508f
C308 VTAIL.n17 B 0.023947f
C309 VTAIL.n18 B 0.022571f
C310 VTAIL.t10 B 0.053646f
C311 VTAIL.n19 B 0.161175f
C312 VTAIL.n20 B 1.03562f
C313 VTAIL.n21 B 0.013508f
C314 VTAIL.n22 B 0.014303f
C315 VTAIL.n23 B 0.031929f
C316 VTAIL.n24 B 0.031929f
C317 VTAIL.n25 B 0.014303f
C318 VTAIL.n26 B 0.013508f
C319 VTAIL.n27 B 0.025139f
C320 VTAIL.n28 B 0.025139f
C321 VTAIL.n29 B 0.013508f
C322 VTAIL.n30 B 0.014303f
C323 VTAIL.n31 B 0.031929f
C324 VTAIL.n32 B 0.031929f
C325 VTAIL.n33 B 0.014303f
C326 VTAIL.n34 B 0.013508f
C327 VTAIL.n35 B 0.025139f
C328 VTAIL.n36 B 0.025139f
C329 VTAIL.n37 B 0.013508f
C330 VTAIL.n38 B 0.013508f
C331 VTAIL.n39 B 0.014303f
C332 VTAIL.n40 B 0.031929f
C333 VTAIL.n41 B 0.031929f
C334 VTAIL.n42 B 0.031929f
C335 VTAIL.n43 B 0.013906f
C336 VTAIL.n44 B 0.013508f
C337 VTAIL.n45 B 0.025139f
C338 VTAIL.n46 B 0.025139f
C339 VTAIL.n47 B 0.013508f
C340 VTAIL.n48 B 0.014303f
C341 VTAIL.n49 B 0.031929f
C342 VTAIL.n50 B 0.064322f
C343 VTAIL.n51 B 0.014303f
C344 VTAIL.n52 B 0.013508f
C345 VTAIL.n53 B 0.056733f
C346 VTAIL.n54 B 0.035455f
C347 VTAIL.n55 B 0.45678f
C348 VTAIL.t5 B 0.197064f
C349 VTAIL.t8 B 0.197064f
C350 VTAIL.n56 B 1.65929f
C351 VTAIL.n57 B 2.07584f
C352 VTAIL.t3 B 0.197064f
C353 VTAIL.t1 B 0.197064f
C354 VTAIL.n58 B 1.6593f
C355 VTAIL.n59 B 2.07583f
C356 VTAIL.n60 B 0.032621f
C357 VTAIL.n61 B 0.025139f
C358 VTAIL.n62 B 0.013508f
C359 VTAIL.n63 B 0.031929f
C360 VTAIL.n64 B 0.014303f
C361 VTAIL.n65 B 0.025139f
C362 VTAIL.n66 B 0.013906f
C363 VTAIL.n67 B 0.031929f
C364 VTAIL.n68 B 0.013508f
C365 VTAIL.n69 B 0.014303f
C366 VTAIL.n70 B 0.025139f
C367 VTAIL.n71 B 0.013508f
C368 VTAIL.n72 B 0.031929f
C369 VTAIL.n73 B 0.014303f
C370 VTAIL.n74 B 0.025139f
C371 VTAIL.n75 B 0.013508f
C372 VTAIL.n76 B 0.023947f
C373 VTAIL.n77 B 0.022571f
C374 VTAIL.t0 B 0.053646f
C375 VTAIL.n78 B 0.161174f
C376 VTAIL.n79 B 1.03562f
C377 VTAIL.n80 B 0.013508f
C378 VTAIL.n81 B 0.014303f
C379 VTAIL.n82 B 0.031929f
C380 VTAIL.n83 B 0.031929f
C381 VTAIL.n84 B 0.014303f
C382 VTAIL.n85 B 0.013508f
C383 VTAIL.n86 B 0.025139f
C384 VTAIL.n87 B 0.025139f
C385 VTAIL.n88 B 0.013508f
C386 VTAIL.n89 B 0.014303f
C387 VTAIL.n90 B 0.031929f
C388 VTAIL.n91 B 0.031929f
C389 VTAIL.n92 B 0.014303f
C390 VTAIL.n93 B 0.013508f
C391 VTAIL.n94 B 0.025139f
C392 VTAIL.n95 B 0.025139f
C393 VTAIL.n96 B 0.013508f
C394 VTAIL.n97 B 0.014303f
C395 VTAIL.n98 B 0.031929f
C396 VTAIL.n99 B 0.031929f
C397 VTAIL.n100 B 0.031929f
C398 VTAIL.n101 B 0.013906f
C399 VTAIL.n102 B 0.013508f
C400 VTAIL.n103 B 0.025139f
C401 VTAIL.n104 B 0.025139f
C402 VTAIL.n105 B 0.013508f
C403 VTAIL.n106 B 0.014303f
C404 VTAIL.n107 B 0.031929f
C405 VTAIL.n108 B 0.064322f
C406 VTAIL.n109 B 0.014303f
C407 VTAIL.n110 B 0.013508f
C408 VTAIL.n111 B 0.056733f
C409 VTAIL.n112 B 0.035455f
C410 VTAIL.n113 B 0.45678f
C411 VTAIL.t6 B 0.197064f
C412 VTAIL.t7 B 0.197064f
C413 VTAIL.n114 B 1.6593f
C414 VTAIL.n115 B 0.681677f
C415 VTAIL.n116 B 0.032621f
C416 VTAIL.n117 B 0.025139f
C417 VTAIL.n118 B 0.013508f
C418 VTAIL.n119 B 0.031929f
C419 VTAIL.n120 B 0.014303f
C420 VTAIL.n121 B 0.025139f
C421 VTAIL.n122 B 0.013906f
C422 VTAIL.n123 B 0.031929f
C423 VTAIL.n124 B 0.013508f
C424 VTAIL.n125 B 0.014303f
C425 VTAIL.n126 B 0.025139f
C426 VTAIL.n127 B 0.013508f
C427 VTAIL.n128 B 0.031929f
C428 VTAIL.n129 B 0.014303f
C429 VTAIL.n130 B 0.025139f
C430 VTAIL.n131 B 0.013508f
C431 VTAIL.n132 B 0.023947f
C432 VTAIL.n133 B 0.022571f
C433 VTAIL.t9 B 0.053646f
C434 VTAIL.n134 B 0.161174f
C435 VTAIL.n135 B 1.03562f
C436 VTAIL.n136 B 0.013508f
C437 VTAIL.n137 B 0.014303f
C438 VTAIL.n138 B 0.031929f
C439 VTAIL.n139 B 0.031929f
C440 VTAIL.n140 B 0.014303f
C441 VTAIL.n141 B 0.013508f
C442 VTAIL.n142 B 0.025139f
C443 VTAIL.n143 B 0.025139f
C444 VTAIL.n144 B 0.013508f
C445 VTAIL.n145 B 0.014303f
C446 VTAIL.n146 B 0.031929f
C447 VTAIL.n147 B 0.031929f
C448 VTAIL.n148 B 0.014303f
C449 VTAIL.n149 B 0.013508f
C450 VTAIL.n150 B 0.025139f
C451 VTAIL.n151 B 0.025139f
C452 VTAIL.n152 B 0.013508f
C453 VTAIL.n153 B 0.014303f
C454 VTAIL.n154 B 0.031929f
C455 VTAIL.n155 B 0.031929f
C456 VTAIL.n156 B 0.031929f
C457 VTAIL.n157 B 0.013906f
C458 VTAIL.n158 B 0.013508f
C459 VTAIL.n159 B 0.025139f
C460 VTAIL.n160 B 0.025139f
C461 VTAIL.n161 B 0.013508f
C462 VTAIL.n162 B 0.014303f
C463 VTAIL.n163 B 0.031929f
C464 VTAIL.n164 B 0.064322f
C465 VTAIL.n165 B 0.014303f
C466 VTAIL.n166 B 0.013508f
C467 VTAIL.n167 B 0.056733f
C468 VTAIL.n168 B 0.035455f
C469 VTAIL.n169 B 1.58559f
C470 VTAIL.n170 B 0.032621f
C471 VTAIL.n171 B 0.025139f
C472 VTAIL.n172 B 0.013508f
C473 VTAIL.n173 B 0.031929f
C474 VTAIL.n174 B 0.014303f
C475 VTAIL.n175 B 0.025139f
C476 VTAIL.n176 B 0.013906f
C477 VTAIL.n177 B 0.031929f
C478 VTAIL.n178 B 0.014303f
C479 VTAIL.n179 B 0.025139f
C480 VTAIL.n180 B 0.013508f
C481 VTAIL.n181 B 0.031929f
C482 VTAIL.n182 B 0.014303f
C483 VTAIL.n183 B 0.025139f
C484 VTAIL.n184 B 0.013508f
C485 VTAIL.n185 B 0.023947f
C486 VTAIL.n186 B 0.022571f
C487 VTAIL.t11 B 0.053646f
C488 VTAIL.n187 B 0.161175f
C489 VTAIL.n188 B 1.03562f
C490 VTAIL.n189 B 0.013508f
C491 VTAIL.n190 B 0.014303f
C492 VTAIL.n191 B 0.031929f
C493 VTAIL.n192 B 0.031929f
C494 VTAIL.n193 B 0.014303f
C495 VTAIL.n194 B 0.013508f
C496 VTAIL.n195 B 0.025139f
C497 VTAIL.n196 B 0.025139f
C498 VTAIL.n197 B 0.013508f
C499 VTAIL.n198 B 0.014303f
C500 VTAIL.n199 B 0.031929f
C501 VTAIL.n200 B 0.031929f
C502 VTAIL.n201 B 0.014303f
C503 VTAIL.n202 B 0.013508f
C504 VTAIL.n203 B 0.025139f
C505 VTAIL.n204 B 0.025139f
C506 VTAIL.n205 B 0.013508f
C507 VTAIL.n206 B 0.013508f
C508 VTAIL.n207 B 0.014303f
C509 VTAIL.n208 B 0.031929f
C510 VTAIL.n209 B 0.031929f
C511 VTAIL.n210 B 0.031929f
C512 VTAIL.n211 B 0.013906f
C513 VTAIL.n212 B 0.013508f
C514 VTAIL.n213 B 0.025139f
C515 VTAIL.n214 B 0.025139f
C516 VTAIL.n215 B 0.013508f
C517 VTAIL.n216 B 0.014303f
C518 VTAIL.n217 B 0.031929f
C519 VTAIL.n218 B 0.064322f
C520 VTAIL.n219 B 0.014303f
C521 VTAIL.n220 B 0.013508f
C522 VTAIL.n221 B 0.056733f
C523 VTAIL.n222 B 0.035455f
C524 VTAIL.n223 B 1.51453f
C525 VP.t2 B 1.90806f
C526 VP.n0 B 0.760629f
C527 VP.n1 B 0.020467f
C528 VP.n2 B 0.019297f
C529 VP.n3 B 0.020467f
C530 VP.t4 B 1.90806f
C531 VP.n4 B 0.69609f
C532 VP.n5 B 0.020467f
C533 VP.n6 B 0.019297f
C534 VP.n7 B 0.020467f
C535 VP.t1 B 1.90806f
C536 VP.n8 B 0.760629f
C537 VP.t0 B 1.90806f
C538 VP.n9 B 0.760629f
C539 VP.n10 B 0.020467f
C540 VP.n11 B 0.019297f
C541 VP.n12 B 0.020467f
C542 VP.t5 B 1.90806f
C543 VP.n13 B 0.75782f
C544 VP.t3 B 2.18379f
C545 VP.n14 B 0.708252f
C546 VP.n15 B 0.249719f
C547 VP.n16 B 0.037954f
C548 VP.n17 B 0.037954f
C549 VP.n18 B 0.03738f
C550 VP.n19 B 0.020467f
C551 VP.n20 B 0.020467f
C552 VP.n21 B 0.020467f
C553 VP.n22 B 0.040781f
C554 VP.n23 B 0.037954f
C555 VP.n24 B 0.030459f
C556 VP.n25 B 0.033028f
C557 VP.n26 B 1.18924f
C558 VP.n27 B 1.2038f
C559 VP.n28 B 0.033028f
C560 VP.n29 B 0.030459f
C561 VP.n30 B 0.037954f
C562 VP.n31 B 0.040781f
C563 VP.n32 B 0.020467f
C564 VP.n33 B 0.020467f
C565 VP.n34 B 0.020467f
C566 VP.n35 B 0.03738f
C567 VP.n36 B 0.037954f
C568 VP.n37 B 0.037954f
C569 VP.n38 B 0.020467f
C570 VP.n39 B 0.020467f
C571 VP.n40 B 0.020467f
C572 VP.n41 B 0.037954f
C573 VP.n42 B 0.037954f
C574 VP.n43 B 0.03738f
C575 VP.n44 B 0.020467f
C576 VP.n45 B 0.020467f
C577 VP.n46 B 0.020467f
C578 VP.n47 B 0.040781f
C579 VP.n48 B 0.037954f
C580 VP.n49 B 0.030459f
C581 VP.n50 B 0.033028f
C582 VP.n51 B 0.050904f
.ends

