* NGSPICE file created from diff_pair_sample_0548.ext - technology: sky130A

.subckt diff_pair_sample_0548 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t0 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=0.4785 ps=3.23 w=2.9 l=2.19
X1 B.t11 B.t9 B.t10 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0 ps=0 w=2.9 l=2.19
X2 VDD1.t5 VP.t0 VTAIL.t3 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=1.131 ps=6.58 w=2.9 l=2.19
X3 VDD2.t3 VN.t1 VTAIL.t10 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=1.131 ps=6.58 w=2.9 l=2.19
X4 VTAIL.t4 VP.t1 VDD1.t4 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=0.4785 ps=3.23 w=2.9 l=2.19
X5 VDD1.t3 VP.t2 VTAIL.t5 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0.4785 ps=3.23 w=2.9 l=2.19
X6 VTAIL.t9 VN.t2 VDD2.t5 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=0.4785 ps=3.23 w=2.9 l=2.19
X7 B.t8 B.t6 B.t7 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0 ps=0 w=2.9 l=2.19
X8 B.t5 B.t3 B.t4 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0 ps=0 w=2.9 l=2.19
X9 VDD1.t2 VP.t3 VTAIL.t0 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=1.131 ps=6.58 w=2.9 l=2.19
X10 VDD1.t1 VP.t4 VTAIL.t1 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0.4785 ps=3.23 w=2.9 l=2.19
X11 VDD2.t1 VN.t3 VTAIL.t8 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=1.131 ps=6.58 w=2.9 l=2.19
X12 B.t2 B.t0 B.t1 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0 ps=0 w=2.9 l=2.19
X13 VTAIL.t2 VP.t5 VDD1.t0 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=0.4785 pd=3.23 as=0.4785 ps=3.23 w=2.9 l=2.19
X14 VDD2.t2 VN.t4 VTAIL.t7 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0.4785 ps=3.23 w=2.9 l=2.19
X15 VDD2.t4 VN.t5 VTAIL.t6 w_n2986_n1548# sky130_fd_pr__pfet_01v8 ad=1.131 pd=6.58 as=0.4785 ps=3.23 w=2.9 l=2.19
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n13 VN.n12 97.6287
R11 VN.n27 VN.n26 97.6287
R12 VN.n3 VN.t5 64.2823
R13 VN.n17 VN.t1 64.2823
R14 VN.n4 VN.n3 59.4178
R15 VN.n18 VN.n17 59.4178
R16 VN.n10 VN.n1 41.5458
R17 VN.n24 VN.n15 41.5458
R18 VN VN.n27 40.4224
R19 VN.n6 VN.n1 39.6083
R20 VN.n20 VN.n15 39.6083
R21 VN.n4 VN.t0 31.9137
R22 VN.n12 VN.t3 31.9137
R23 VN.n18 VN.t2 31.9137
R24 VN.n26 VN.t4 31.9137
R25 VN.n6 VN.n5 24.5923
R26 VN.n11 VN.n10 24.5923
R27 VN.n20 VN.n19 24.5923
R28 VN.n25 VN.n24 24.5923
R29 VN.n12 VN.n11 13.2801
R30 VN.n26 VN.n25 13.2801
R31 VN.n5 VN.n4 12.2964
R32 VN.n19 VN.n18 12.2964
R33 VN.n17 VN.n16 9.60944
R34 VN.n3 VN.n2 9.60944
R35 VN.n27 VN.n14 0.278335
R36 VN.n13 VN.n0 0.278335
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153485
R46 VDD2.n1 VDD2.t4 153.567
R47 VDD2.n2 VDD2.t2 151.994
R48 VDD2.n1 VDD2.n0 141.273
R49 VDD2 VDD2.n3 141.27
R50 VDD2.n2 VDD2.n1 33.2756
R51 VDD2.n3 VDD2.t5 11.2091
R52 VDD2.n3 VDD2.t3 11.2091
R53 VDD2.n0 VDD2.t0 11.2091
R54 VDD2.n0 VDD2.t1 11.2091
R55 VDD2 VDD2.n2 1.688
R56 VTAIL.n7 VTAIL.t10 135.315
R57 VTAIL.n10 VTAIL.t3 135.315
R58 VTAIL.n11 VTAIL.t8 135.315
R59 VTAIL.n2 VTAIL.t0 135.315
R60 VTAIL.n9 VTAIL.n8 124.106
R61 VTAIL.n6 VTAIL.n5 124.106
R62 VTAIL.n1 VTAIL.n0 124.106
R63 VTAIL.n4 VTAIL.n3 124.106
R64 VTAIL.n6 VTAIL.n4 19.2117
R65 VTAIL.n11 VTAIL.n10 17.0393
R66 VTAIL.n0 VTAIL.t6 11.2091
R67 VTAIL.n0 VTAIL.t11 11.2091
R68 VTAIL.n3 VTAIL.t5 11.2091
R69 VTAIL.n3 VTAIL.t4 11.2091
R70 VTAIL.n8 VTAIL.t1 11.2091
R71 VTAIL.n8 VTAIL.t2 11.2091
R72 VTAIL.n5 VTAIL.t7 11.2091
R73 VTAIL.n5 VTAIL.t9 11.2091
R74 VTAIL.n7 VTAIL.n6 2.17291
R75 VTAIL.n10 VTAIL.n9 2.17291
R76 VTAIL.n4 VTAIL.n2 2.17291
R77 VTAIL VTAIL.n11 1.57162
R78 VTAIL.n9 VTAIL.n7 1.55653
R79 VTAIL.n2 VTAIL.n1 1.55653
R80 VTAIL VTAIL.n1 0.601793
R81 B.n238 B.n237 585
R82 B.n236 B.n83 585
R83 B.n235 B.n234 585
R84 B.n233 B.n84 585
R85 B.n232 B.n231 585
R86 B.n230 B.n85 585
R87 B.n229 B.n228 585
R88 B.n227 B.n86 585
R89 B.n226 B.n225 585
R90 B.n224 B.n87 585
R91 B.n223 B.n222 585
R92 B.n221 B.n88 585
R93 B.n220 B.n219 585
R94 B.n218 B.n89 585
R95 B.n217 B.n216 585
R96 B.n215 B.n214 585
R97 B.n213 B.n93 585
R98 B.n212 B.n211 585
R99 B.n210 B.n94 585
R100 B.n209 B.n208 585
R101 B.n207 B.n95 585
R102 B.n206 B.n205 585
R103 B.n204 B.n96 585
R104 B.n203 B.n202 585
R105 B.n200 B.n97 585
R106 B.n199 B.n198 585
R107 B.n197 B.n100 585
R108 B.n196 B.n195 585
R109 B.n194 B.n101 585
R110 B.n193 B.n192 585
R111 B.n191 B.n102 585
R112 B.n190 B.n189 585
R113 B.n188 B.n103 585
R114 B.n187 B.n186 585
R115 B.n185 B.n104 585
R116 B.n184 B.n183 585
R117 B.n182 B.n105 585
R118 B.n181 B.n180 585
R119 B.n179 B.n106 585
R120 B.n239 B.n82 585
R121 B.n241 B.n240 585
R122 B.n242 B.n81 585
R123 B.n244 B.n243 585
R124 B.n245 B.n80 585
R125 B.n247 B.n246 585
R126 B.n248 B.n79 585
R127 B.n250 B.n249 585
R128 B.n251 B.n78 585
R129 B.n253 B.n252 585
R130 B.n254 B.n77 585
R131 B.n256 B.n255 585
R132 B.n257 B.n76 585
R133 B.n259 B.n258 585
R134 B.n260 B.n75 585
R135 B.n262 B.n261 585
R136 B.n263 B.n74 585
R137 B.n265 B.n264 585
R138 B.n266 B.n73 585
R139 B.n268 B.n267 585
R140 B.n269 B.n72 585
R141 B.n271 B.n270 585
R142 B.n272 B.n71 585
R143 B.n274 B.n273 585
R144 B.n275 B.n70 585
R145 B.n277 B.n276 585
R146 B.n278 B.n69 585
R147 B.n280 B.n279 585
R148 B.n281 B.n68 585
R149 B.n283 B.n282 585
R150 B.n284 B.n67 585
R151 B.n286 B.n285 585
R152 B.n287 B.n66 585
R153 B.n289 B.n288 585
R154 B.n290 B.n65 585
R155 B.n292 B.n291 585
R156 B.n293 B.n64 585
R157 B.n295 B.n294 585
R158 B.n296 B.n63 585
R159 B.n298 B.n297 585
R160 B.n299 B.n62 585
R161 B.n301 B.n300 585
R162 B.n302 B.n61 585
R163 B.n304 B.n303 585
R164 B.n305 B.n60 585
R165 B.n307 B.n306 585
R166 B.n308 B.n59 585
R167 B.n310 B.n309 585
R168 B.n311 B.n58 585
R169 B.n313 B.n312 585
R170 B.n314 B.n57 585
R171 B.n316 B.n315 585
R172 B.n317 B.n56 585
R173 B.n319 B.n318 585
R174 B.n320 B.n55 585
R175 B.n322 B.n321 585
R176 B.n323 B.n54 585
R177 B.n325 B.n324 585
R178 B.n326 B.n53 585
R179 B.n328 B.n327 585
R180 B.n329 B.n52 585
R181 B.n331 B.n330 585
R182 B.n332 B.n51 585
R183 B.n334 B.n333 585
R184 B.n335 B.n50 585
R185 B.n337 B.n336 585
R186 B.n338 B.n49 585
R187 B.n340 B.n339 585
R188 B.n341 B.n48 585
R189 B.n343 B.n342 585
R190 B.n344 B.n47 585
R191 B.n346 B.n345 585
R192 B.n347 B.n46 585
R193 B.n349 B.n348 585
R194 B.n350 B.n45 585
R195 B.n352 B.n351 585
R196 B.n412 B.n411 585
R197 B.n410 B.n21 585
R198 B.n409 B.n408 585
R199 B.n407 B.n22 585
R200 B.n406 B.n405 585
R201 B.n404 B.n23 585
R202 B.n403 B.n402 585
R203 B.n401 B.n24 585
R204 B.n400 B.n399 585
R205 B.n398 B.n25 585
R206 B.n397 B.n396 585
R207 B.n395 B.n26 585
R208 B.n394 B.n393 585
R209 B.n392 B.n27 585
R210 B.n391 B.n390 585
R211 B.n389 B.n388 585
R212 B.n387 B.n31 585
R213 B.n386 B.n385 585
R214 B.n384 B.n32 585
R215 B.n383 B.n382 585
R216 B.n381 B.n33 585
R217 B.n380 B.n379 585
R218 B.n378 B.n34 585
R219 B.n377 B.n376 585
R220 B.n374 B.n35 585
R221 B.n373 B.n372 585
R222 B.n371 B.n38 585
R223 B.n370 B.n369 585
R224 B.n368 B.n39 585
R225 B.n367 B.n366 585
R226 B.n365 B.n40 585
R227 B.n364 B.n363 585
R228 B.n362 B.n41 585
R229 B.n361 B.n360 585
R230 B.n359 B.n42 585
R231 B.n358 B.n357 585
R232 B.n356 B.n43 585
R233 B.n355 B.n354 585
R234 B.n353 B.n44 585
R235 B.n413 B.n20 585
R236 B.n415 B.n414 585
R237 B.n416 B.n19 585
R238 B.n418 B.n417 585
R239 B.n419 B.n18 585
R240 B.n421 B.n420 585
R241 B.n422 B.n17 585
R242 B.n424 B.n423 585
R243 B.n425 B.n16 585
R244 B.n427 B.n426 585
R245 B.n428 B.n15 585
R246 B.n430 B.n429 585
R247 B.n431 B.n14 585
R248 B.n433 B.n432 585
R249 B.n434 B.n13 585
R250 B.n436 B.n435 585
R251 B.n437 B.n12 585
R252 B.n439 B.n438 585
R253 B.n440 B.n11 585
R254 B.n442 B.n441 585
R255 B.n443 B.n10 585
R256 B.n445 B.n444 585
R257 B.n446 B.n9 585
R258 B.n448 B.n447 585
R259 B.n449 B.n8 585
R260 B.n451 B.n450 585
R261 B.n452 B.n7 585
R262 B.n454 B.n453 585
R263 B.n455 B.n6 585
R264 B.n457 B.n456 585
R265 B.n458 B.n5 585
R266 B.n460 B.n459 585
R267 B.n461 B.n4 585
R268 B.n463 B.n462 585
R269 B.n464 B.n3 585
R270 B.n466 B.n465 585
R271 B.n467 B.n0 585
R272 B.n2 B.n1 585
R273 B.n125 B.n124 585
R274 B.n127 B.n126 585
R275 B.n128 B.n123 585
R276 B.n130 B.n129 585
R277 B.n131 B.n122 585
R278 B.n133 B.n132 585
R279 B.n134 B.n121 585
R280 B.n136 B.n135 585
R281 B.n137 B.n120 585
R282 B.n139 B.n138 585
R283 B.n140 B.n119 585
R284 B.n142 B.n141 585
R285 B.n143 B.n118 585
R286 B.n145 B.n144 585
R287 B.n146 B.n117 585
R288 B.n148 B.n147 585
R289 B.n149 B.n116 585
R290 B.n151 B.n150 585
R291 B.n152 B.n115 585
R292 B.n154 B.n153 585
R293 B.n155 B.n114 585
R294 B.n157 B.n156 585
R295 B.n158 B.n113 585
R296 B.n160 B.n159 585
R297 B.n161 B.n112 585
R298 B.n163 B.n162 585
R299 B.n164 B.n111 585
R300 B.n166 B.n165 585
R301 B.n167 B.n110 585
R302 B.n169 B.n168 585
R303 B.n170 B.n109 585
R304 B.n172 B.n171 585
R305 B.n173 B.n108 585
R306 B.n175 B.n174 585
R307 B.n176 B.n107 585
R308 B.n178 B.n177 585
R309 B.n179 B.n178 564.573
R310 B.n239 B.n238 564.573
R311 B.n353 B.n352 564.573
R312 B.n413 B.n412 564.573
R313 B.n469 B.n468 256.663
R314 B.n98 B.t0 239.244
R315 B.n90 B.t9 239.244
R316 B.n36 B.t3 239.244
R317 B.n28 B.t6 239.244
R318 B.n468 B.n467 235.042
R319 B.n468 B.n2 235.042
R320 B.n90 B.t10 192.53
R321 B.n36 B.t5 192.53
R322 B.n98 B.t1 192.529
R323 B.n28 B.t8 192.529
R324 B.n180 B.n179 163.367
R325 B.n180 B.n105 163.367
R326 B.n184 B.n105 163.367
R327 B.n185 B.n184 163.367
R328 B.n186 B.n185 163.367
R329 B.n186 B.n103 163.367
R330 B.n190 B.n103 163.367
R331 B.n191 B.n190 163.367
R332 B.n192 B.n191 163.367
R333 B.n192 B.n101 163.367
R334 B.n196 B.n101 163.367
R335 B.n197 B.n196 163.367
R336 B.n198 B.n197 163.367
R337 B.n198 B.n97 163.367
R338 B.n203 B.n97 163.367
R339 B.n204 B.n203 163.367
R340 B.n205 B.n204 163.367
R341 B.n205 B.n95 163.367
R342 B.n209 B.n95 163.367
R343 B.n210 B.n209 163.367
R344 B.n211 B.n210 163.367
R345 B.n211 B.n93 163.367
R346 B.n215 B.n93 163.367
R347 B.n216 B.n215 163.367
R348 B.n216 B.n89 163.367
R349 B.n220 B.n89 163.367
R350 B.n221 B.n220 163.367
R351 B.n222 B.n221 163.367
R352 B.n222 B.n87 163.367
R353 B.n226 B.n87 163.367
R354 B.n227 B.n226 163.367
R355 B.n228 B.n227 163.367
R356 B.n228 B.n85 163.367
R357 B.n232 B.n85 163.367
R358 B.n233 B.n232 163.367
R359 B.n234 B.n233 163.367
R360 B.n234 B.n83 163.367
R361 B.n238 B.n83 163.367
R362 B.n352 B.n45 163.367
R363 B.n348 B.n45 163.367
R364 B.n348 B.n347 163.367
R365 B.n347 B.n346 163.367
R366 B.n346 B.n47 163.367
R367 B.n342 B.n47 163.367
R368 B.n342 B.n341 163.367
R369 B.n341 B.n340 163.367
R370 B.n340 B.n49 163.367
R371 B.n336 B.n49 163.367
R372 B.n336 B.n335 163.367
R373 B.n335 B.n334 163.367
R374 B.n334 B.n51 163.367
R375 B.n330 B.n51 163.367
R376 B.n330 B.n329 163.367
R377 B.n329 B.n328 163.367
R378 B.n328 B.n53 163.367
R379 B.n324 B.n53 163.367
R380 B.n324 B.n323 163.367
R381 B.n323 B.n322 163.367
R382 B.n322 B.n55 163.367
R383 B.n318 B.n55 163.367
R384 B.n318 B.n317 163.367
R385 B.n317 B.n316 163.367
R386 B.n316 B.n57 163.367
R387 B.n312 B.n57 163.367
R388 B.n312 B.n311 163.367
R389 B.n311 B.n310 163.367
R390 B.n310 B.n59 163.367
R391 B.n306 B.n59 163.367
R392 B.n306 B.n305 163.367
R393 B.n305 B.n304 163.367
R394 B.n304 B.n61 163.367
R395 B.n300 B.n61 163.367
R396 B.n300 B.n299 163.367
R397 B.n299 B.n298 163.367
R398 B.n298 B.n63 163.367
R399 B.n294 B.n63 163.367
R400 B.n294 B.n293 163.367
R401 B.n293 B.n292 163.367
R402 B.n292 B.n65 163.367
R403 B.n288 B.n65 163.367
R404 B.n288 B.n287 163.367
R405 B.n287 B.n286 163.367
R406 B.n286 B.n67 163.367
R407 B.n282 B.n67 163.367
R408 B.n282 B.n281 163.367
R409 B.n281 B.n280 163.367
R410 B.n280 B.n69 163.367
R411 B.n276 B.n69 163.367
R412 B.n276 B.n275 163.367
R413 B.n275 B.n274 163.367
R414 B.n274 B.n71 163.367
R415 B.n270 B.n71 163.367
R416 B.n270 B.n269 163.367
R417 B.n269 B.n268 163.367
R418 B.n268 B.n73 163.367
R419 B.n264 B.n73 163.367
R420 B.n264 B.n263 163.367
R421 B.n263 B.n262 163.367
R422 B.n262 B.n75 163.367
R423 B.n258 B.n75 163.367
R424 B.n258 B.n257 163.367
R425 B.n257 B.n256 163.367
R426 B.n256 B.n77 163.367
R427 B.n252 B.n77 163.367
R428 B.n252 B.n251 163.367
R429 B.n251 B.n250 163.367
R430 B.n250 B.n79 163.367
R431 B.n246 B.n79 163.367
R432 B.n246 B.n245 163.367
R433 B.n245 B.n244 163.367
R434 B.n244 B.n81 163.367
R435 B.n240 B.n81 163.367
R436 B.n240 B.n239 163.367
R437 B.n412 B.n21 163.367
R438 B.n408 B.n21 163.367
R439 B.n408 B.n407 163.367
R440 B.n407 B.n406 163.367
R441 B.n406 B.n23 163.367
R442 B.n402 B.n23 163.367
R443 B.n402 B.n401 163.367
R444 B.n401 B.n400 163.367
R445 B.n400 B.n25 163.367
R446 B.n396 B.n25 163.367
R447 B.n396 B.n395 163.367
R448 B.n395 B.n394 163.367
R449 B.n394 B.n27 163.367
R450 B.n390 B.n27 163.367
R451 B.n390 B.n389 163.367
R452 B.n389 B.n31 163.367
R453 B.n385 B.n31 163.367
R454 B.n385 B.n384 163.367
R455 B.n384 B.n383 163.367
R456 B.n383 B.n33 163.367
R457 B.n379 B.n33 163.367
R458 B.n379 B.n378 163.367
R459 B.n378 B.n377 163.367
R460 B.n377 B.n35 163.367
R461 B.n372 B.n35 163.367
R462 B.n372 B.n371 163.367
R463 B.n371 B.n370 163.367
R464 B.n370 B.n39 163.367
R465 B.n366 B.n39 163.367
R466 B.n366 B.n365 163.367
R467 B.n365 B.n364 163.367
R468 B.n364 B.n41 163.367
R469 B.n360 B.n41 163.367
R470 B.n360 B.n359 163.367
R471 B.n359 B.n358 163.367
R472 B.n358 B.n43 163.367
R473 B.n354 B.n43 163.367
R474 B.n354 B.n353 163.367
R475 B.n414 B.n413 163.367
R476 B.n414 B.n19 163.367
R477 B.n418 B.n19 163.367
R478 B.n419 B.n418 163.367
R479 B.n420 B.n419 163.367
R480 B.n420 B.n17 163.367
R481 B.n424 B.n17 163.367
R482 B.n425 B.n424 163.367
R483 B.n426 B.n425 163.367
R484 B.n426 B.n15 163.367
R485 B.n430 B.n15 163.367
R486 B.n431 B.n430 163.367
R487 B.n432 B.n431 163.367
R488 B.n432 B.n13 163.367
R489 B.n436 B.n13 163.367
R490 B.n437 B.n436 163.367
R491 B.n438 B.n437 163.367
R492 B.n438 B.n11 163.367
R493 B.n442 B.n11 163.367
R494 B.n443 B.n442 163.367
R495 B.n444 B.n443 163.367
R496 B.n444 B.n9 163.367
R497 B.n448 B.n9 163.367
R498 B.n449 B.n448 163.367
R499 B.n450 B.n449 163.367
R500 B.n450 B.n7 163.367
R501 B.n454 B.n7 163.367
R502 B.n455 B.n454 163.367
R503 B.n456 B.n455 163.367
R504 B.n456 B.n5 163.367
R505 B.n460 B.n5 163.367
R506 B.n461 B.n460 163.367
R507 B.n462 B.n461 163.367
R508 B.n462 B.n3 163.367
R509 B.n466 B.n3 163.367
R510 B.n467 B.n466 163.367
R511 B.n125 B.n2 163.367
R512 B.n126 B.n125 163.367
R513 B.n126 B.n123 163.367
R514 B.n130 B.n123 163.367
R515 B.n131 B.n130 163.367
R516 B.n132 B.n131 163.367
R517 B.n132 B.n121 163.367
R518 B.n136 B.n121 163.367
R519 B.n137 B.n136 163.367
R520 B.n138 B.n137 163.367
R521 B.n138 B.n119 163.367
R522 B.n142 B.n119 163.367
R523 B.n143 B.n142 163.367
R524 B.n144 B.n143 163.367
R525 B.n144 B.n117 163.367
R526 B.n148 B.n117 163.367
R527 B.n149 B.n148 163.367
R528 B.n150 B.n149 163.367
R529 B.n150 B.n115 163.367
R530 B.n154 B.n115 163.367
R531 B.n155 B.n154 163.367
R532 B.n156 B.n155 163.367
R533 B.n156 B.n113 163.367
R534 B.n160 B.n113 163.367
R535 B.n161 B.n160 163.367
R536 B.n162 B.n161 163.367
R537 B.n162 B.n111 163.367
R538 B.n166 B.n111 163.367
R539 B.n167 B.n166 163.367
R540 B.n168 B.n167 163.367
R541 B.n168 B.n109 163.367
R542 B.n172 B.n109 163.367
R543 B.n173 B.n172 163.367
R544 B.n174 B.n173 163.367
R545 B.n174 B.n107 163.367
R546 B.n178 B.n107 163.367
R547 B.n91 B.t11 143.657
R548 B.n37 B.t4 143.657
R549 B.n99 B.t2 143.655
R550 B.n29 B.t7 143.655
R551 B.n201 B.n99 59.5399
R552 B.n92 B.n91 59.5399
R553 B.n375 B.n37 59.5399
R554 B.n30 B.n29 59.5399
R555 B.n99 B.n98 48.8732
R556 B.n91 B.n90 48.8732
R557 B.n37 B.n36 48.8732
R558 B.n29 B.n28 48.8732
R559 B.n411 B.n20 36.6834
R560 B.n351 B.n44 36.6834
R561 B.n237 B.n82 36.6834
R562 B.n177 B.n106 36.6834
R563 B B.n469 18.0485
R564 B.n415 B.n20 10.6151
R565 B.n416 B.n415 10.6151
R566 B.n417 B.n416 10.6151
R567 B.n417 B.n18 10.6151
R568 B.n421 B.n18 10.6151
R569 B.n422 B.n421 10.6151
R570 B.n423 B.n422 10.6151
R571 B.n423 B.n16 10.6151
R572 B.n427 B.n16 10.6151
R573 B.n428 B.n427 10.6151
R574 B.n429 B.n428 10.6151
R575 B.n429 B.n14 10.6151
R576 B.n433 B.n14 10.6151
R577 B.n434 B.n433 10.6151
R578 B.n435 B.n434 10.6151
R579 B.n435 B.n12 10.6151
R580 B.n439 B.n12 10.6151
R581 B.n440 B.n439 10.6151
R582 B.n441 B.n440 10.6151
R583 B.n441 B.n10 10.6151
R584 B.n445 B.n10 10.6151
R585 B.n446 B.n445 10.6151
R586 B.n447 B.n446 10.6151
R587 B.n447 B.n8 10.6151
R588 B.n451 B.n8 10.6151
R589 B.n452 B.n451 10.6151
R590 B.n453 B.n452 10.6151
R591 B.n453 B.n6 10.6151
R592 B.n457 B.n6 10.6151
R593 B.n458 B.n457 10.6151
R594 B.n459 B.n458 10.6151
R595 B.n459 B.n4 10.6151
R596 B.n463 B.n4 10.6151
R597 B.n464 B.n463 10.6151
R598 B.n465 B.n464 10.6151
R599 B.n465 B.n0 10.6151
R600 B.n411 B.n410 10.6151
R601 B.n410 B.n409 10.6151
R602 B.n409 B.n22 10.6151
R603 B.n405 B.n22 10.6151
R604 B.n405 B.n404 10.6151
R605 B.n404 B.n403 10.6151
R606 B.n403 B.n24 10.6151
R607 B.n399 B.n24 10.6151
R608 B.n399 B.n398 10.6151
R609 B.n398 B.n397 10.6151
R610 B.n397 B.n26 10.6151
R611 B.n393 B.n26 10.6151
R612 B.n393 B.n392 10.6151
R613 B.n392 B.n391 10.6151
R614 B.n388 B.n387 10.6151
R615 B.n387 B.n386 10.6151
R616 B.n386 B.n32 10.6151
R617 B.n382 B.n32 10.6151
R618 B.n382 B.n381 10.6151
R619 B.n381 B.n380 10.6151
R620 B.n380 B.n34 10.6151
R621 B.n376 B.n34 10.6151
R622 B.n374 B.n373 10.6151
R623 B.n373 B.n38 10.6151
R624 B.n369 B.n38 10.6151
R625 B.n369 B.n368 10.6151
R626 B.n368 B.n367 10.6151
R627 B.n367 B.n40 10.6151
R628 B.n363 B.n40 10.6151
R629 B.n363 B.n362 10.6151
R630 B.n362 B.n361 10.6151
R631 B.n361 B.n42 10.6151
R632 B.n357 B.n42 10.6151
R633 B.n357 B.n356 10.6151
R634 B.n356 B.n355 10.6151
R635 B.n355 B.n44 10.6151
R636 B.n351 B.n350 10.6151
R637 B.n350 B.n349 10.6151
R638 B.n349 B.n46 10.6151
R639 B.n345 B.n46 10.6151
R640 B.n345 B.n344 10.6151
R641 B.n344 B.n343 10.6151
R642 B.n343 B.n48 10.6151
R643 B.n339 B.n48 10.6151
R644 B.n339 B.n338 10.6151
R645 B.n338 B.n337 10.6151
R646 B.n337 B.n50 10.6151
R647 B.n333 B.n50 10.6151
R648 B.n333 B.n332 10.6151
R649 B.n332 B.n331 10.6151
R650 B.n331 B.n52 10.6151
R651 B.n327 B.n52 10.6151
R652 B.n327 B.n326 10.6151
R653 B.n326 B.n325 10.6151
R654 B.n325 B.n54 10.6151
R655 B.n321 B.n54 10.6151
R656 B.n321 B.n320 10.6151
R657 B.n320 B.n319 10.6151
R658 B.n319 B.n56 10.6151
R659 B.n315 B.n56 10.6151
R660 B.n315 B.n314 10.6151
R661 B.n314 B.n313 10.6151
R662 B.n313 B.n58 10.6151
R663 B.n309 B.n58 10.6151
R664 B.n309 B.n308 10.6151
R665 B.n308 B.n307 10.6151
R666 B.n307 B.n60 10.6151
R667 B.n303 B.n60 10.6151
R668 B.n303 B.n302 10.6151
R669 B.n302 B.n301 10.6151
R670 B.n301 B.n62 10.6151
R671 B.n297 B.n62 10.6151
R672 B.n297 B.n296 10.6151
R673 B.n296 B.n295 10.6151
R674 B.n295 B.n64 10.6151
R675 B.n291 B.n64 10.6151
R676 B.n291 B.n290 10.6151
R677 B.n290 B.n289 10.6151
R678 B.n289 B.n66 10.6151
R679 B.n285 B.n66 10.6151
R680 B.n285 B.n284 10.6151
R681 B.n284 B.n283 10.6151
R682 B.n283 B.n68 10.6151
R683 B.n279 B.n68 10.6151
R684 B.n279 B.n278 10.6151
R685 B.n278 B.n277 10.6151
R686 B.n277 B.n70 10.6151
R687 B.n273 B.n70 10.6151
R688 B.n273 B.n272 10.6151
R689 B.n272 B.n271 10.6151
R690 B.n271 B.n72 10.6151
R691 B.n267 B.n72 10.6151
R692 B.n267 B.n266 10.6151
R693 B.n266 B.n265 10.6151
R694 B.n265 B.n74 10.6151
R695 B.n261 B.n74 10.6151
R696 B.n261 B.n260 10.6151
R697 B.n260 B.n259 10.6151
R698 B.n259 B.n76 10.6151
R699 B.n255 B.n76 10.6151
R700 B.n255 B.n254 10.6151
R701 B.n254 B.n253 10.6151
R702 B.n253 B.n78 10.6151
R703 B.n249 B.n78 10.6151
R704 B.n249 B.n248 10.6151
R705 B.n248 B.n247 10.6151
R706 B.n247 B.n80 10.6151
R707 B.n243 B.n80 10.6151
R708 B.n243 B.n242 10.6151
R709 B.n242 B.n241 10.6151
R710 B.n241 B.n82 10.6151
R711 B.n124 B.n1 10.6151
R712 B.n127 B.n124 10.6151
R713 B.n128 B.n127 10.6151
R714 B.n129 B.n128 10.6151
R715 B.n129 B.n122 10.6151
R716 B.n133 B.n122 10.6151
R717 B.n134 B.n133 10.6151
R718 B.n135 B.n134 10.6151
R719 B.n135 B.n120 10.6151
R720 B.n139 B.n120 10.6151
R721 B.n140 B.n139 10.6151
R722 B.n141 B.n140 10.6151
R723 B.n141 B.n118 10.6151
R724 B.n145 B.n118 10.6151
R725 B.n146 B.n145 10.6151
R726 B.n147 B.n146 10.6151
R727 B.n147 B.n116 10.6151
R728 B.n151 B.n116 10.6151
R729 B.n152 B.n151 10.6151
R730 B.n153 B.n152 10.6151
R731 B.n153 B.n114 10.6151
R732 B.n157 B.n114 10.6151
R733 B.n158 B.n157 10.6151
R734 B.n159 B.n158 10.6151
R735 B.n159 B.n112 10.6151
R736 B.n163 B.n112 10.6151
R737 B.n164 B.n163 10.6151
R738 B.n165 B.n164 10.6151
R739 B.n165 B.n110 10.6151
R740 B.n169 B.n110 10.6151
R741 B.n170 B.n169 10.6151
R742 B.n171 B.n170 10.6151
R743 B.n171 B.n108 10.6151
R744 B.n175 B.n108 10.6151
R745 B.n176 B.n175 10.6151
R746 B.n177 B.n176 10.6151
R747 B.n181 B.n106 10.6151
R748 B.n182 B.n181 10.6151
R749 B.n183 B.n182 10.6151
R750 B.n183 B.n104 10.6151
R751 B.n187 B.n104 10.6151
R752 B.n188 B.n187 10.6151
R753 B.n189 B.n188 10.6151
R754 B.n189 B.n102 10.6151
R755 B.n193 B.n102 10.6151
R756 B.n194 B.n193 10.6151
R757 B.n195 B.n194 10.6151
R758 B.n195 B.n100 10.6151
R759 B.n199 B.n100 10.6151
R760 B.n200 B.n199 10.6151
R761 B.n202 B.n96 10.6151
R762 B.n206 B.n96 10.6151
R763 B.n207 B.n206 10.6151
R764 B.n208 B.n207 10.6151
R765 B.n208 B.n94 10.6151
R766 B.n212 B.n94 10.6151
R767 B.n213 B.n212 10.6151
R768 B.n214 B.n213 10.6151
R769 B.n218 B.n217 10.6151
R770 B.n219 B.n218 10.6151
R771 B.n219 B.n88 10.6151
R772 B.n223 B.n88 10.6151
R773 B.n224 B.n223 10.6151
R774 B.n225 B.n224 10.6151
R775 B.n225 B.n86 10.6151
R776 B.n229 B.n86 10.6151
R777 B.n230 B.n229 10.6151
R778 B.n231 B.n230 10.6151
R779 B.n231 B.n84 10.6151
R780 B.n235 B.n84 10.6151
R781 B.n236 B.n235 10.6151
R782 B.n237 B.n236 10.6151
R783 B.n469 B.n0 8.11757
R784 B.n469 B.n1 8.11757
R785 B.n388 B.n30 6.5566
R786 B.n376 B.n375 6.5566
R787 B.n202 B.n201 6.5566
R788 B.n214 B.n92 6.5566
R789 B.n391 B.n30 4.05904
R790 B.n375 B.n374 4.05904
R791 B.n201 B.n200 4.05904
R792 B.n217 B.n92 4.05904
R793 VP.n11 VP.n8 161.3
R794 VP.n13 VP.n12 161.3
R795 VP.n14 VP.n7 161.3
R796 VP.n16 VP.n15 161.3
R797 VP.n17 VP.n6 161.3
R798 VP.n36 VP.n0 161.3
R799 VP.n35 VP.n34 161.3
R800 VP.n33 VP.n1 161.3
R801 VP.n32 VP.n31 161.3
R802 VP.n30 VP.n2 161.3
R803 VP.n28 VP.n27 161.3
R804 VP.n26 VP.n3 161.3
R805 VP.n25 VP.n24 161.3
R806 VP.n23 VP.n4 161.3
R807 VP.n22 VP.n21 161.3
R808 VP.n20 VP.n5 97.6287
R809 VP.n38 VP.n37 97.6287
R810 VP.n19 VP.n18 97.6287
R811 VP.n9 VP.t4 64.2823
R812 VP.n10 VP.n9 59.4178
R813 VP.n24 VP.n23 41.5458
R814 VP.n35 VP.n1 41.5458
R815 VP.n16 VP.n7 41.5458
R816 VP.n20 VP.n19 40.1436
R817 VP.n24 VP.n3 39.6083
R818 VP.n31 VP.n1 39.6083
R819 VP.n12 VP.n7 39.6083
R820 VP.n5 VP.t2 31.9137
R821 VP.n29 VP.t1 31.9137
R822 VP.n37 VP.t3 31.9137
R823 VP.n18 VP.t0 31.9137
R824 VP.n10 VP.t5 31.9137
R825 VP.n23 VP.n22 24.5923
R826 VP.n28 VP.n3 24.5923
R827 VP.n31 VP.n30 24.5923
R828 VP.n36 VP.n35 24.5923
R829 VP.n17 VP.n16 24.5923
R830 VP.n12 VP.n11 24.5923
R831 VP.n22 VP.n5 13.2801
R832 VP.n37 VP.n36 13.2801
R833 VP.n18 VP.n17 13.2801
R834 VP.n29 VP.n28 12.2964
R835 VP.n30 VP.n29 12.2964
R836 VP.n11 VP.n10 12.2964
R837 VP.n9 VP.n8 9.60944
R838 VP.n19 VP.n6 0.278335
R839 VP.n21 VP.n20 0.278335
R840 VP.n38 VP.n0 0.278335
R841 VP.n13 VP.n8 0.189894
R842 VP.n14 VP.n13 0.189894
R843 VP.n15 VP.n14 0.189894
R844 VP.n15 VP.n6 0.189894
R845 VP.n21 VP.n4 0.189894
R846 VP.n25 VP.n4 0.189894
R847 VP.n26 VP.n25 0.189894
R848 VP.n27 VP.n26 0.189894
R849 VP.n27 VP.n2 0.189894
R850 VP.n32 VP.n2 0.189894
R851 VP.n33 VP.n32 0.189894
R852 VP.n34 VP.n33 0.189894
R853 VP.n34 VP.n0 0.189894
R854 VP VP.n38 0.153485
R855 VDD1 VDD1.t1 153.681
R856 VDD1.n1 VDD1.t3 153.567
R857 VDD1.n1 VDD1.n0 141.273
R858 VDD1.n3 VDD1.n2 140.786
R859 VDD1.n3 VDD1.n1 34.9449
R860 VDD1.n2 VDD1.t0 11.2091
R861 VDD1.n2 VDD1.t5 11.2091
R862 VDD1.n0 VDD1.t4 11.2091
R863 VDD1.n0 VDD1.t2 11.2091
R864 VDD1 VDD1.n3 0.485414
C0 B VDD1 1.27244f
C1 w_n2986_n1548# VDD1 1.54741f
C2 B VTAIL 1.4884f
C3 w_n2986_n1548# VTAIL 1.61595f
C4 B VP 1.61666f
C5 VP w_n2986_n1548# 5.77173f
C6 VDD2 VDD1 1.24465f
C7 VDD2 VTAIL 4.22258f
C8 VN B 0.976542f
C9 VN w_n2986_n1548# 5.38933f
C10 VDD2 VP 0.428827f
C11 VTAIL VDD1 4.17251f
C12 VDD2 VN 1.86142f
C13 VP VDD1 2.13236f
C14 VP VTAIL 2.51082f
C15 VN VDD1 0.155557f
C16 VN VTAIL 2.49666f
C17 B w_n2986_n1548# 6.580359f
C18 VN VP 4.84826f
C19 VDD2 B 1.33689f
C20 VDD2 w_n2986_n1548# 1.61888f
C21 VDD2 VSUBS 0.998417f
C22 VDD1 VSUBS 1.612975f
C23 VTAIL VSUBS 0.508025f
C24 VN VSUBS 4.99338f
C25 VP VSUBS 2.101475f
C26 B VSUBS 3.26827f
C27 w_n2986_n1548# VSUBS 58.585297f
C28 VDD1.t1 VSUBS 0.392837f
C29 VDD1.t3 VSUBS 0.392428f
C30 VDD1.t4 VSUBS 0.052452f
C31 VDD1.t2 VSUBS 0.052452f
C32 VDD1.n0 VSUBS 0.273296f
C33 VDD1.n1 VSUBS 2.26576f
C34 VDD1.t0 VSUBS 0.052452f
C35 VDD1.t5 VSUBS 0.052452f
C36 VDD1.n2 VSUBS 0.271596f
C37 VDD1.n3 VSUBS 1.89284f
C38 VP.n0 VSUBS 0.070682f
C39 VP.t3 VSUBS 0.844582f
C40 VP.n1 VSUBS 0.043371f
C41 VP.n2 VSUBS 0.053615f
C42 VP.t1 VSUBS 0.844582f
C43 VP.n3 VSUBS 0.106495f
C44 VP.n4 VSUBS 0.053615f
C45 VP.t2 VSUBS 0.844582f
C46 VP.n5 VSUBS 0.525239f
C47 VP.n6 VSUBS 0.070682f
C48 VP.t0 VSUBS 0.844582f
C49 VP.n7 VSUBS 0.043371f
C50 VP.n8 VSUBS 0.455703f
C51 VP.t5 VSUBS 0.844582f
C52 VP.t4 VSUBS 1.17234f
C53 VP.n9 VSUBS 0.485077f
C54 VP.n10 VSUBS 0.504288f
C55 VP.n11 VSUBS 0.074883f
C56 VP.n12 VSUBS 0.106495f
C57 VP.n13 VSUBS 0.053615f
C58 VP.n14 VSUBS 0.053615f
C59 VP.n15 VSUBS 0.053615f
C60 VP.n16 VSUBS 0.105433f
C61 VP.n17 VSUBS 0.076846f
C62 VP.n18 VSUBS 0.525239f
C63 VP.n19 VSUBS 2.10556f
C64 VP.n20 VSUBS 2.15371f
C65 VP.n21 VSUBS 0.070682f
C66 VP.n22 VSUBS 0.076846f
C67 VP.n23 VSUBS 0.105433f
C68 VP.n24 VSUBS 0.043371f
C69 VP.n25 VSUBS 0.053615f
C70 VP.n26 VSUBS 0.053615f
C71 VP.n27 VSUBS 0.053615f
C72 VP.n28 VSUBS 0.074883f
C73 VP.n29 VSUBS 0.367173f
C74 VP.n30 VSUBS 0.074883f
C75 VP.n31 VSUBS 0.106495f
C76 VP.n32 VSUBS 0.053615f
C77 VP.n33 VSUBS 0.053615f
C78 VP.n34 VSUBS 0.053615f
C79 VP.n35 VSUBS 0.105433f
C80 VP.n36 VSUBS 0.076846f
C81 VP.n37 VSUBS 0.525239f
C82 VP.n38 VSUBS 0.076547f
C83 B.n0 VSUBS 0.006965f
C84 B.n1 VSUBS 0.006965f
C85 B.n2 VSUBS 0.0103f
C86 B.n3 VSUBS 0.007893f
C87 B.n4 VSUBS 0.007893f
C88 B.n5 VSUBS 0.007893f
C89 B.n6 VSUBS 0.007893f
C90 B.n7 VSUBS 0.007893f
C91 B.n8 VSUBS 0.007893f
C92 B.n9 VSUBS 0.007893f
C93 B.n10 VSUBS 0.007893f
C94 B.n11 VSUBS 0.007893f
C95 B.n12 VSUBS 0.007893f
C96 B.n13 VSUBS 0.007893f
C97 B.n14 VSUBS 0.007893f
C98 B.n15 VSUBS 0.007893f
C99 B.n16 VSUBS 0.007893f
C100 B.n17 VSUBS 0.007893f
C101 B.n18 VSUBS 0.007893f
C102 B.n19 VSUBS 0.007893f
C103 B.n20 VSUBS 0.01949f
C104 B.n21 VSUBS 0.007893f
C105 B.n22 VSUBS 0.007893f
C106 B.n23 VSUBS 0.007893f
C107 B.n24 VSUBS 0.007893f
C108 B.n25 VSUBS 0.007893f
C109 B.n26 VSUBS 0.007893f
C110 B.n27 VSUBS 0.007893f
C111 B.t7 VSUBS 0.077919f
C112 B.t8 VSUBS 0.093108f
C113 B.t6 VSUBS 0.346926f
C114 B.n28 VSUBS 0.08705f
C115 B.n29 VSUBS 0.071096f
C116 B.n30 VSUBS 0.018288f
C117 B.n31 VSUBS 0.007893f
C118 B.n32 VSUBS 0.007893f
C119 B.n33 VSUBS 0.007893f
C120 B.n34 VSUBS 0.007893f
C121 B.n35 VSUBS 0.007893f
C122 B.t4 VSUBS 0.077919f
C123 B.t5 VSUBS 0.093108f
C124 B.t3 VSUBS 0.346926f
C125 B.n36 VSUBS 0.08705f
C126 B.n37 VSUBS 0.071096f
C127 B.n38 VSUBS 0.007893f
C128 B.n39 VSUBS 0.007893f
C129 B.n40 VSUBS 0.007893f
C130 B.n41 VSUBS 0.007893f
C131 B.n42 VSUBS 0.007893f
C132 B.n43 VSUBS 0.007893f
C133 B.n44 VSUBS 0.020441f
C134 B.n45 VSUBS 0.007893f
C135 B.n46 VSUBS 0.007893f
C136 B.n47 VSUBS 0.007893f
C137 B.n48 VSUBS 0.007893f
C138 B.n49 VSUBS 0.007893f
C139 B.n50 VSUBS 0.007893f
C140 B.n51 VSUBS 0.007893f
C141 B.n52 VSUBS 0.007893f
C142 B.n53 VSUBS 0.007893f
C143 B.n54 VSUBS 0.007893f
C144 B.n55 VSUBS 0.007893f
C145 B.n56 VSUBS 0.007893f
C146 B.n57 VSUBS 0.007893f
C147 B.n58 VSUBS 0.007893f
C148 B.n59 VSUBS 0.007893f
C149 B.n60 VSUBS 0.007893f
C150 B.n61 VSUBS 0.007893f
C151 B.n62 VSUBS 0.007893f
C152 B.n63 VSUBS 0.007893f
C153 B.n64 VSUBS 0.007893f
C154 B.n65 VSUBS 0.007893f
C155 B.n66 VSUBS 0.007893f
C156 B.n67 VSUBS 0.007893f
C157 B.n68 VSUBS 0.007893f
C158 B.n69 VSUBS 0.007893f
C159 B.n70 VSUBS 0.007893f
C160 B.n71 VSUBS 0.007893f
C161 B.n72 VSUBS 0.007893f
C162 B.n73 VSUBS 0.007893f
C163 B.n74 VSUBS 0.007893f
C164 B.n75 VSUBS 0.007893f
C165 B.n76 VSUBS 0.007893f
C166 B.n77 VSUBS 0.007893f
C167 B.n78 VSUBS 0.007893f
C168 B.n79 VSUBS 0.007893f
C169 B.n80 VSUBS 0.007893f
C170 B.n81 VSUBS 0.007893f
C171 B.n82 VSUBS 0.02032f
C172 B.n83 VSUBS 0.007893f
C173 B.n84 VSUBS 0.007893f
C174 B.n85 VSUBS 0.007893f
C175 B.n86 VSUBS 0.007893f
C176 B.n87 VSUBS 0.007893f
C177 B.n88 VSUBS 0.007893f
C178 B.n89 VSUBS 0.007893f
C179 B.t11 VSUBS 0.077919f
C180 B.t10 VSUBS 0.093108f
C181 B.t9 VSUBS 0.346926f
C182 B.n90 VSUBS 0.08705f
C183 B.n91 VSUBS 0.071096f
C184 B.n92 VSUBS 0.018288f
C185 B.n93 VSUBS 0.007893f
C186 B.n94 VSUBS 0.007893f
C187 B.n95 VSUBS 0.007893f
C188 B.n96 VSUBS 0.007893f
C189 B.n97 VSUBS 0.007893f
C190 B.t2 VSUBS 0.077919f
C191 B.t1 VSUBS 0.093108f
C192 B.t0 VSUBS 0.346926f
C193 B.n98 VSUBS 0.08705f
C194 B.n99 VSUBS 0.071096f
C195 B.n100 VSUBS 0.007893f
C196 B.n101 VSUBS 0.007893f
C197 B.n102 VSUBS 0.007893f
C198 B.n103 VSUBS 0.007893f
C199 B.n104 VSUBS 0.007893f
C200 B.n105 VSUBS 0.007893f
C201 B.n106 VSUBS 0.020441f
C202 B.n107 VSUBS 0.007893f
C203 B.n108 VSUBS 0.007893f
C204 B.n109 VSUBS 0.007893f
C205 B.n110 VSUBS 0.007893f
C206 B.n111 VSUBS 0.007893f
C207 B.n112 VSUBS 0.007893f
C208 B.n113 VSUBS 0.007893f
C209 B.n114 VSUBS 0.007893f
C210 B.n115 VSUBS 0.007893f
C211 B.n116 VSUBS 0.007893f
C212 B.n117 VSUBS 0.007893f
C213 B.n118 VSUBS 0.007893f
C214 B.n119 VSUBS 0.007893f
C215 B.n120 VSUBS 0.007893f
C216 B.n121 VSUBS 0.007893f
C217 B.n122 VSUBS 0.007893f
C218 B.n123 VSUBS 0.007893f
C219 B.n124 VSUBS 0.007893f
C220 B.n125 VSUBS 0.007893f
C221 B.n126 VSUBS 0.007893f
C222 B.n127 VSUBS 0.007893f
C223 B.n128 VSUBS 0.007893f
C224 B.n129 VSUBS 0.007893f
C225 B.n130 VSUBS 0.007893f
C226 B.n131 VSUBS 0.007893f
C227 B.n132 VSUBS 0.007893f
C228 B.n133 VSUBS 0.007893f
C229 B.n134 VSUBS 0.007893f
C230 B.n135 VSUBS 0.007893f
C231 B.n136 VSUBS 0.007893f
C232 B.n137 VSUBS 0.007893f
C233 B.n138 VSUBS 0.007893f
C234 B.n139 VSUBS 0.007893f
C235 B.n140 VSUBS 0.007893f
C236 B.n141 VSUBS 0.007893f
C237 B.n142 VSUBS 0.007893f
C238 B.n143 VSUBS 0.007893f
C239 B.n144 VSUBS 0.007893f
C240 B.n145 VSUBS 0.007893f
C241 B.n146 VSUBS 0.007893f
C242 B.n147 VSUBS 0.007893f
C243 B.n148 VSUBS 0.007893f
C244 B.n149 VSUBS 0.007893f
C245 B.n150 VSUBS 0.007893f
C246 B.n151 VSUBS 0.007893f
C247 B.n152 VSUBS 0.007893f
C248 B.n153 VSUBS 0.007893f
C249 B.n154 VSUBS 0.007893f
C250 B.n155 VSUBS 0.007893f
C251 B.n156 VSUBS 0.007893f
C252 B.n157 VSUBS 0.007893f
C253 B.n158 VSUBS 0.007893f
C254 B.n159 VSUBS 0.007893f
C255 B.n160 VSUBS 0.007893f
C256 B.n161 VSUBS 0.007893f
C257 B.n162 VSUBS 0.007893f
C258 B.n163 VSUBS 0.007893f
C259 B.n164 VSUBS 0.007893f
C260 B.n165 VSUBS 0.007893f
C261 B.n166 VSUBS 0.007893f
C262 B.n167 VSUBS 0.007893f
C263 B.n168 VSUBS 0.007893f
C264 B.n169 VSUBS 0.007893f
C265 B.n170 VSUBS 0.007893f
C266 B.n171 VSUBS 0.007893f
C267 B.n172 VSUBS 0.007893f
C268 B.n173 VSUBS 0.007893f
C269 B.n174 VSUBS 0.007893f
C270 B.n175 VSUBS 0.007893f
C271 B.n176 VSUBS 0.007893f
C272 B.n177 VSUBS 0.01949f
C273 B.n178 VSUBS 0.01949f
C274 B.n179 VSUBS 0.020441f
C275 B.n180 VSUBS 0.007893f
C276 B.n181 VSUBS 0.007893f
C277 B.n182 VSUBS 0.007893f
C278 B.n183 VSUBS 0.007893f
C279 B.n184 VSUBS 0.007893f
C280 B.n185 VSUBS 0.007893f
C281 B.n186 VSUBS 0.007893f
C282 B.n187 VSUBS 0.007893f
C283 B.n188 VSUBS 0.007893f
C284 B.n189 VSUBS 0.007893f
C285 B.n190 VSUBS 0.007893f
C286 B.n191 VSUBS 0.007893f
C287 B.n192 VSUBS 0.007893f
C288 B.n193 VSUBS 0.007893f
C289 B.n194 VSUBS 0.007893f
C290 B.n195 VSUBS 0.007893f
C291 B.n196 VSUBS 0.007893f
C292 B.n197 VSUBS 0.007893f
C293 B.n198 VSUBS 0.007893f
C294 B.n199 VSUBS 0.007893f
C295 B.n200 VSUBS 0.005456f
C296 B.n201 VSUBS 0.018288f
C297 B.n202 VSUBS 0.006384f
C298 B.n203 VSUBS 0.007893f
C299 B.n204 VSUBS 0.007893f
C300 B.n205 VSUBS 0.007893f
C301 B.n206 VSUBS 0.007893f
C302 B.n207 VSUBS 0.007893f
C303 B.n208 VSUBS 0.007893f
C304 B.n209 VSUBS 0.007893f
C305 B.n210 VSUBS 0.007893f
C306 B.n211 VSUBS 0.007893f
C307 B.n212 VSUBS 0.007893f
C308 B.n213 VSUBS 0.007893f
C309 B.n214 VSUBS 0.006384f
C310 B.n215 VSUBS 0.007893f
C311 B.n216 VSUBS 0.007893f
C312 B.n217 VSUBS 0.005456f
C313 B.n218 VSUBS 0.007893f
C314 B.n219 VSUBS 0.007893f
C315 B.n220 VSUBS 0.007893f
C316 B.n221 VSUBS 0.007893f
C317 B.n222 VSUBS 0.007893f
C318 B.n223 VSUBS 0.007893f
C319 B.n224 VSUBS 0.007893f
C320 B.n225 VSUBS 0.007893f
C321 B.n226 VSUBS 0.007893f
C322 B.n227 VSUBS 0.007893f
C323 B.n228 VSUBS 0.007893f
C324 B.n229 VSUBS 0.007893f
C325 B.n230 VSUBS 0.007893f
C326 B.n231 VSUBS 0.007893f
C327 B.n232 VSUBS 0.007893f
C328 B.n233 VSUBS 0.007893f
C329 B.n234 VSUBS 0.007893f
C330 B.n235 VSUBS 0.007893f
C331 B.n236 VSUBS 0.007893f
C332 B.n237 VSUBS 0.019611f
C333 B.n238 VSUBS 0.020441f
C334 B.n239 VSUBS 0.01949f
C335 B.n240 VSUBS 0.007893f
C336 B.n241 VSUBS 0.007893f
C337 B.n242 VSUBS 0.007893f
C338 B.n243 VSUBS 0.007893f
C339 B.n244 VSUBS 0.007893f
C340 B.n245 VSUBS 0.007893f
C341 B.n246 VSUBS 0.007893f
C342 B.n247 VSUBS 0.007893f
C343 B.n248 VSUBS 0.007893f
C344 B.n249 VSUBS 0.007893f
C345 B.n250 VSUBS 0.007893f
C346 B.n251 VSUBS 0.007893f
C347 B.n252 VSUBS 0.007893f
C348 B.n253 VSUBS 0.007893f
C349 B.n254 VSUBS 0.007893f
C350 B.n255 VSUBS 0.007893f
C351 B.n256 VSUBS 0.007893f
C352 B.n257 VSUBS 0.007893f
C353 B.n258 VSUBS 0.007893f
C354 B.n259 VSUBS 0.007893f
C355 B.n260 VSUBS 0.007893f
C356 B.n261 VSUBS 0.007893f
C357 B.n262 VSUBS 0.007893f
C358 B.n263 VSUBS 0.007893f
C359 B.n264 VSUBS 0.007893f
C360 B.n265 VSUBS 0.007893f
C361 B.n266 VSUBS 0.007893f
C362 B.n267 VSUBS 0.007893f
C363 B.n268 VSUBS 0.007893f
C364 B.n269 VSUBS 0.007893f
C365 B.n270 VSUBS 0.007893f
C366 B.n271 VSUBS 0.007893f
C367 B.n272 VSUBS 0.007893f
C368 B.n273 VSUBS 0.007893f
C369 B.n274 VSUBS 0.007893f
C370 B.n275 VSUBS 0.007893f
C371 B.n276 VSUBS 0.007893f
C372 B.n277 VSUBS 0.007893f
C373 B.n278 VSUBS 0.007893f
C374 B.n279 VSUBS 0.007893f
C375 B.n280 VSUBS 0.007893f
C376 B.n281 VSUBS 0.007893f
C377 B.n282 VSUBS 0.007893f
C378 B.n283 VSUBS 0.007893f
C379 B.n284 VSUBS 0.007893f
C380 B.n285 VSUBS 0.007893f
C381 B.n286 VSUBS 0.007893f
C382 B.n287 VSUBS 0.007893f
C383 B.n288 VSUBS 0.007893f
C384 B.n289 VSUBS 0.007893f
C385 B.n290 VSUBS 0.007893f
C386 B.n291 VSUBS 0.007893f
C387 B.n292 VSUBS 0.007893f
C388 B.n293 VSUBS 0.007893f
C389 B.n294 VSUBS 0.007893f
C390 B.n295 VSUBS 0.007893f
C391 B.n296 VSUBS 0.007893f
C392 B.n297 VSUBS 0.007893f
C393 B.n298 VSUBS 0.007893f
C394 B.n299 VSUBS 0.007893f
C395 B.n300 VSUBS 0.007893f
C396 B.n301 VSUBS 0.007893f
C397 B.n302 VSUBS 0.007893f
C398 B.n303 VSUBS 0.007893f
C399 B.n304 VSUBS 0.007893f
C400 B.n305 VSUBS 0.007893f
C401 B.n306 VSUBS 0.007893f
C402 B.n307 VSUBS 0.007893f
C403 B.n308 VSUBS 0.007893f
C404 B.n309 VSUBS 0.007893f
C405 B.n310 VSUBS 0.007893f
C406 B.n311 VSUBS 0.007893f
C407 B.n312 VSUBS 0.007893f
C408 B.n313 VSUBS 0.007893f
C409 B.n314 VSUBS 0.007893f
C410 B.n315 VSUBS 0.007893f
C411 B.n316 VSUBS 0.007893f
C412 B.n317 VSUBS 0.007893f
C413 B.n318 VSUBS 0.007893f
C414 B.n319 VSUBS 0.007893f
C415 B.n320 VSUBS 0.007893f
C416 B.n321 VSUBS 0.007893f
C417 B.n322 VSUBS 0.007893f
C418 B.n323 VSUBS 0.007893f
C419 B.n324 VSUBS 0.007893f
C420 B.n325 VSUBS 0.007893f
C421 B.n326 VSUBS 0.007893f
C422 B.n327 VSUBS 0.007893f
C423 B.n328 VSUBS 0.007893f
C424 B.n329 VSUBS 0.007893f
C425 B.n330 VSUBS 0.007893f
C426 B.n331 VSUBS 0.007893f
C427 B.n332 VSUBS 0.007893f
C428 B.n333 VSUBS 0.007893f
C429 B.n334 VSUBS 0.007893f
C430 B.n335 VSUBS 0.007893f
C431 B.n336 VSUBS 0.007893f
C432 B.n337 VSUBS 0.007893f
C433 B.n338 VSUBS 0.007893f
C434 B.n339 VSUBS 0.007893f
C435 B.n340 VSUBS 0.007893f
C436 B.n341 VSUBS 0.007893f
C437 B.n342 VSUBS 0.007893f
C438 B.n343 VSUBS 0.007893f
C439 B.n344 VSUBS 0.007893f
C440 B.n345 VSUBS 0.007893f
C441 B.n346 VSUBS 0.007893f
C442 B.n347 VSUBS 0.007893f
C443 B.n348 VSUBS 0.007893f
C444 B.n349 VSUBS 0.007893f
C445 B.n350 VSUBS 0.007893f
C446 B.n351 VSUBS 0.01949f
C447 B.n352 VSUBS 0.01949f
C448 B.n353 VSUBS 0.020441f
C449 B.n354 VSUBS 0.007893f
C450 B.n355 VSUBS 0.007893f
C451 B.n356 VSUBS 0.007893f
C452 B.n357 VSUBS 0.007893f
C453 B.n358 VSUBS 0.007893f
C454 B.n359 VSUBS 0.007893f
C455 B.n360 VSUBS 0.007893f
C456 B.n361 VSUBS 0.007893f
C457 B.n362 VSUBS 0.007893f
C458 B.n363 VSUBS 0.007893f
C459 B.n364 VSUBS 0.007893f
C460 B.n365 VSUBS 0.007893f
C461 B.n366 VSUBS 0.007893f
C462 B.n367 VSUBS 0.007893f
C463 B.n368 VSUBS 0.007893f
C464 B.n369 VSUBS 0.007893f
C465 B.n370 VSUBS 0.007893f
C466 B.n371 VSUBS 0.007893f
C467 B.n372 VSUBS 0.007893f
C468 B.n373 VSUBS 0.007893f
C469 B.n374 VSUBS 0.005456f
C470 B.n375 VSUBS 0.018288f
C471 B.n376 VSUBS 0.006384f
C472 B.n377 VSUBS 0.007893f
C473 B.n378 VSUBS 0.007893f
C474 B.n379 VSUBS 0.007893f
C475 B.n380 VSUBS 0.007893f
C476 B.n381 VSUBS 0.007893f
C477 B.n382 VSUBS 0.007893f
C478 B.n383 VSUBS 0.007893f
C479 B.n384 VSUBS 0.007893f
C480 B.n385 VSUBS 0.007893f
C481 B.n386 VSUBS 0.007893f
C482 B.n387 VSUBS 0.007893f
C483 B.n388 VSUBS 0.006384f
C484 B.n389 VSUBS 0.007893f
C485 B.n390 VSUBS 0.007893f
C486 B.n391 VSUBS 0.005456f
C487 B.n392 VSUBS 0.007893f
C488 B.n393 VSUBS 0.007893f
C489 B.n394 VSUBS 0.007893f
C490 B.n395 VSUBS 0.007893f
C491 B.n396 VSUBS 0.007893f
C492 B.n397 VSUBS 0.007893f
C493 B.n398 VSUBS 0.007893f
C494 B.n399 VSUBS 0.007893f
C495 B.n400 VSUBS 0.007893f
C496 B.n401 VSUBS 0.007893f
C497 B.n402 VSUBS 0.007893f
C498 B.n403 VSUBS 0.007893f
C499 B.n404 VSUBS 0.007893f
C500 B.n405 VSUBS 0.007893f
C501 B.n406 VSUBS 0.007893f
C502 B.n407 VSUBS 0.007893f
C503 B.n408 VSUBS 0.007893f
C504 B.n409 VSUBS 0.007893f
C505 B.n410 VSUBS 0.007893f
C506 B.n411 VSUBS 0.020441f
C507 B.n412 VSUBS 0.020441f
C508 B.n413 VSUBS 0.01949f
C509 B.n414 VSUBS 0.007893f
C510 B.n415 VSUBS 0.007893f
C511 B.n416 VSUBS 0.007893f
C512 B.n417 VSUBS 0.007893f
C513 B.n418 VSUBS 0.007893f
C514 B.n419 VSUBS 0.007893f
C515 B.n420 VSUBS 0.007893f
C516 B.n421 VSUBS 0.007893f
C517 B.n422 VSUBS 0.007893f
C518 B.n423 VSUBS 0.007893f
C519 B.n424 VSUBS 0.007893f
C520 B.n425 VSUBS 0.007893f
C521 B.n426 VSUBS 0.007893f
C522 B.n427 VSUBS 0.007893f
C523 B.n428 VSUBS 0.007893f
C524 B.n429 VSUBS 0.007893f
C525 B.n430 VSUBS 0.007893f
C526 B.n431 VSUBS 0.007893f
C527 B.n432 VSUBS 0.007893f
C528 B.n433 VSUBS 0.007893f
C529 B.n434 VSUBS 0.007893f
C530 B.n435 VSUBS 0.007893f
C531 B.n436 VSUBS 0.007893f
C532 B.n437 VSUBS 0.007893f
C533 B.n438 VSUBS 0.007893f
C534 B.n439 VSUBS 0.007893f
C535 B.n440 VSUBS 0.007893f
C536 B.n441 VSUBS 0.007893f
C537 B.n442 VSUBS 0.007893f
C538 B.n443 VSUBS 0.007893f
C539 B.n444 VSUBS 0.007893f
C540 B.n445 VSUBS 0.007893f
C541 B.n446 VSUBS 0.007893f
C542 B.n447 VSUBS 0.007893f
C543 B.n448 VSUBS 0.007893f
C544 B.n449 VSUBS 0.007893f
C545 B.n450 VSUBS 0.007893f
C546 B.n451 VSUBS 0.007893f
C547 B.n452 VSUBS 0.007893f
C548 B.n453 VSUBS 0.007893f
C549 B.n454 VSUBS 0.007893f
C550 B.n455 VSUBS 0.007893f
C551 B.n456 VSUBS 0.007893f
C552 B.n457 VSUBS 0.007893f
C553 B.n458 VSUBS 0.007893f
C554 B.n459 VSUBS 0.007893f
C555 B.n460 VSUBS 0.007893f
C556 B.n461 VSUBS 0.007893f
C557 B.n462 VSUBS 0.007893f
C558 B.n463 VSUBS 0.007893f
C559 B.n464 VSUBS 0.007893f
C560 B.n465 VSUBS 0.007893f
C561 B.n466 VSUBS 0.007893f
C562 B.n467 VSUBS 0.0103f
C563 B.n468 VSUBS 0.010972f
C564 B.n469 VSUBS 0.02182f
C565 VTAIL.t6 VSUBS 0.071105f
C566 VTAIL.t11 VSUBS 0.071105f
C567 VTAIL.n0 VSUBS 0.316918f
C568 VTAIL.n1 VSUBS 0.612119f
C569 VTAIL.t0 VSUBS 0.474415f
C570 VTAIL.n2 VSUBS 0.805622f
C571 VTAIL.t5 VSUBS 0.071105f
C572 VTAIL.t4 VSUBS 0.071105f
C573 VTAIL.n3 VSUBS 0.316918f
C574 VTAIL.n4 VSUBS 1.71943f
C575 VTAIL.t7 VSUBS 0.071105f
C576 VTAIL.t9 VSUBS 0.071105f
C577 VTAIL.n5 VSUBS 0.316919f
C578 VTAIL.n6 VSUBS 1.71943f
C579 VTAIL.t10 VSUBS 0.474417f
C580 VTAIL.n7 VSUBS 0.80562f
C581 VTAIL.t1 VSUBS 0.071105f
C582 VTAIL.t2 VSUBS 0.071105f
C583 VTAIL.n8 VSUBS 0.316919f
C584 VTAIL.n9 VSUBS 0.769195f
C585 VTAIL.t3 VSUBS 0.474415f
C586 VTAIL.n10 VSUBS 1.53866f
C587 VTAIL.t8 VSUBS 0.474415f
C588 VTAIL.n11 VSUBS 1.47855f
C589 VDD2.t4 VSUBS 0.265177f
C590 VDD2.t0 VSUBS 0.035444f
C591 VDD2.t1 VSUBS 0.035444f
C592 VDD2.n0 VSUBS 0.184675f
C593 VDD2.n1 VSUBS 1.46614f
C594 VDD2.t2 VSUBS 0.262143f
C595 VDD2.n2 VSUBS 1.25655f
C596 VDD2.t5 VSUBS 0.035444f
C597 VDD2.t3 VSUBS 0.035444f
C598 VDD2.n3 VSUBS 0.184665f
C599 VN.n0 VSUBS 0.058765f
C600 VN.t3 VSUBS 0.702189f
C601 VN.n1 VSUBS 0.036059f
C602 VN.n2 VSUBS 0.378873f
C603 VN.t0 VSUBS 0.702189f
C604 VN.t5 VSUBS 0.974684f
C605 VN.n3 VSUBS 0.403295f
C606 VN.n4 VSUBS 0.419267f
C607 VN.n5 VSUBS 0.062258f
C608 VN.n6 VSUBS 0.088541f
C609 VN.n7 VSUBS 0.044576f
C610 VN.n8 VSUBS 0.044576f
C611 VN.n9 VSUBS 0.044576f
C612 VN.n10 VSUBS 0.087658f
C613 VN.n11 VSUBS 0.06389f
C614 VN.n12 VSUBS 0.436686f
C615 VN.n13 VSUBS 0.063641f
C616 VN.n14 VSUBS 0.058765f
C617 VN.t4 VSUBS 0.702189f
C618 VN.n15 VSUBS 0.036059f
C619 VN.n16 VSUBS 0.378873f
C620 VN.t2 VSUBS 0.702189f
C621 VN.t1 VSUBS 0.974684f
C622 VN.n17 VSUBS 0.403295f
C623 VN.n18 VSUBS 0.419267f
C624 VN.n19 VSUBS 0.062258f
C625 VN.n20 VSUBS 0.088541f
C626 VN.n21 VSUBS 0.044576f
C627 VN.n22 VSUBS 0.044576f
C628 VN.n23 VSUBS 0.044576f
C629 VN.n24 VSUBS 0.087658f
C630 VN.n25 VSUBS 0.06389f
C631 VN.n26 VSUBS 0.436686f
C632 VN.n27 VSUBS 1.77546f
.ends

