* NGSPICE file created from diff_pair_sample_0569.ext - technology: sky130A

.subckt diff_pair_sample_0569 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=1.3884 ps=7.9 w=3.56 l=2.41
X1 VDD1.t5 VP.t0 VTAIL.t1 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0.5874 ps=3.89 w=3.56 l=2.41
X2 VTAIL.t7 VN.t1 VDD2.t4 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=0.5874 ps=3.89 w=3.56 l=2.41
X3 B.t11 B.t9 B.t10 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0 ps=0 w=3.56 l=2.41
X4 VDD2.t3 VN.t2 VTAIL.t6 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=1.3884 ps=7.9 w=3.56 l=2.41
X5 VTAIL.t5 VP.t1 VDD1.t4 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=0.5874 ps=3.89 w=3.56 l=2.41
X6 VDD2.t2 VN.t3 VTAIL.t9 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0.5874 ps=3.89 w=3.56 l=2.41
X7 VTAIL.t8 VN.t4 VDD2.t1 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=0.5874 ps=3.89 w=3.56 l=2.41
X8 VDD1.t3 VP.t2 VTAIL.t3 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=1.3884 ps=7.9 w=3.56 l=2.41
X9 VDD1.t2 VP.t3 VTAIL.t2 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0.5874 ps=3.89 w=3.56 l=2.41
X10 VDD2.t0 VN.t5 VTAIL.t10 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0.5874 ps=3.89 w=3.56 l=2.41
X11 B.t8 B.t6 B.t7 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0 ps=0 w=3.56 l=2.41
X12 B.t5 B.t3 B.t4 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0 ps=0 w=3.56 l=2.41
X13 VTAIL.t4 VP.t4 VDD1.t1 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=0.5874 ps=3.89 w=3.56 l=2.41
X14 B.t2 B.t0 B.t1 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=1.3884 pd=7.9 as=0 ps=0 w=3.56 l=2.41
X15 VDD1.t0 VP.t5 VTAIL.t0 w_n3162_n1680# sky130_fd_pr__pfet_01v8 ad=0.5874 pd=3.89 as=1.3884 ps=7.9 w=3.56 l=2.41
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n13 VN.n12 98.9213
R11 VN.n27 VN.n26 98.9213
R12 VN.n3 VN.t5 69.7532
R13 VN.n17 VN.t2 69.7532
R14 VN.n6 VN.n1 53.0692
R15 VN.n20 VN.n15 53.0692
R16 VN.n4 VN.n3 47.8856
R17 VN.n18 VN.n17 47.8856
R18 VN VN.n27 41.8163
R19 VN.n4 VN.t4 35.6005
R20 VN.n12 VN.t0 35.6005
R21 VN.n18 VN.t1 35.6005
R22 VN.n26 VN.t3 35.6005
R23 VN.n10 VN.n1 27.752
R24 VN.n24 VN.n15 27.752
R25 VN.n5 VN.n4 24.3439
R26 VN.n6 VN.n5 24.3439
R27 VN.n11 VN.n10 24.3439
R28 VN.n20 VN.n19 24.3439
R29 VN.n19 VN.n18 24.3439
R30 VN.n25 VN.n24 24.3439
R31 VN.n12 VN.n11 11.6853
R32 VN.n26 VN.n25 11.6853
R33 VN.n17 VN.n16 6.74271
R34 VN.n3 VN.n2 6.74271
R35 VN.n27 VN.n14 0.278398
R36 VN.n13 VN.n0 0.278398
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153422
R46 VTAIL.n7 VTAIL.t6 113.912
R47 VTAIL.n11 VTAIL.t11 113.912
R48 VTAIL.n2 VTAIL.t0 113.912
R49 VTAIL.n10 VTAIL.t3 113.912
R50 VTAIL.n9 VTAIL.n8 104.781
R51 VTAIL.n6 VTAIL.n5 104.781
R52 VTAIL.n1 VTAIL.n0 104.781
R53 VTAIL.n4 VTAIL.n3 104.781
R54 VTAIL.n6 VTAIL.n4 20.16
R55 VTAIL.n11 VTAIL.n10 17.7979
R56 VTAIL.n0 VTAIL.t10 9.13112
R57 VTAIL.n0 VTAIL.t8 9.13112
R58 VTAIL.n3 VTAIL.t1 9.13112
R59 VTAIL.n3 VTAIL.t4 9.13112
R60 VTAIL.n8 VTAIL.t2 9.13112
R61 VTAIL.n8 VTAIL.t5 9.13112
R62 VTAIL.n5 VTAIL.t9 9.13112
R63 VTAIL.n5 VTAIL.t7 9.13112
R64 VTAIL.n7 VTAIL.n6 2.36257
R65 VTAIL.n10 VTAIL.n9 2.36257
R66 VTAIL.n4 VTAIL.n2 2.36257
R67 VTAIL VTAIL.n11 1.71386
R68 VTAIL.n9 VTAIL.n7 1.65136
R69 VTAIL.n2 VTAIL.n1 1.65136
R70 VTAIL VTAIL.n1 0.649207
R71 VDD2.n1 VDD2.t0 132.306
R72 VDD2.n2 VDD2.t2 130.59
R73 VDD2.n1 VDD2.n0 121.995
R74 VDD2 VDD2.n3 121.993
R75 VDD2.n2 VDD2.n1 34.461
R76 VDD2.n3 VDD2.t4 9.13112
R77 VDD2.n3 VDD2.t3 9.13112
R78 VDD2.n0 VDD2.t1 9.13112
R79 VDD2.n0 VDD2.t5 9.13112
R80 VDD2 VDD2.n2 1.83024
R81 VP.n11 VP.n8 161.3
R82 VP.n13 VP.n12 161.3
R83 VP.n14 VP.n7 161.3
R84 VP.n16 VP.n15 161.3
R85 VP.n17 VP.n6 161.3
R86 VP.n37 VP.n0 161.3
R87 VP.n36 VP.n35 161.3
R88 VP.n34 VP.n1 161.3
R89 VP.n33 VP.n32 161.3
R90 VP.n31 VP.n2 161.3
R91 VP.n30 VP.n29 161.3
R92 VP.n28 VP.n3 161.3
R93 VP.n27 VP.n26 161.3
R94 VP.n25 VP.n4 161.3
R95 VP.n24 VP.n23 161.3
R96 VP.n22 VP.n5 161.3
R97 VP.n21 VP.n20 98.9213
R98 VP.n39 VP.n38 98.9213
R99 VP.n19 VP.n18 98.9213
R100 VP.n9 VP.t3 69.7532
R101 VP.n26 VP.n25 53.0692
R102 VP.n32 VP.n1 53.0692
R103 VP.n12 VP.n7 53.0692
R104 VP.n10 VP.n9 47.8856
R105 VP.n21 VP.n19 41.5374
R106 VP.n30 VP.t4 35.6005
R107 VP.n20 VP.t0 35.6005
R108 VP.n38 VP.t5 35.6005
R109 VP.n10 VP.t1 35.6005
R110 VP.n18 VP.t2 35.6005
R111 VP.n25 VP.n24 27.752
R112 VP.n36 VP.n1 27.752
R113 VP.n16 VP.n7 27.752
R114 VP.n24 VP.n5 24.3439
R115 VP.n26 VP.n3 24.3439
R116 VP.n30 VP.n3 24.3439
R117 VP.n31 VP.n30 24.3439
R118 VP.n32 VP.n31 24.3439
R119 VP.n37 VP.n36 24.3439
R120 VP.n17 VP.n16 24.3439
R121 VP.n11 VP.n10 24.3439
R122 VP.n12 VP.n11 24.3439
R123 VP.n20 VP.n5 11.6853
R124 VP.n38 VP.n37 11.6853
R125 VP.n18 VP.n17 11.6853
R126 VP.n9 VP.n8 6.74271
R127 VP.n19 VP.n6 0.278398
R128 VP.n22 VP.n21 0.278398
R129 VP.n39 VP.n0 0.278398
R130 VP.n13 VP.n8 0.189894
R131 VP.n14 VP.n13 0.189894
R132 VP.n15 VP.n14 0.189894
R133 VP.n15 VP.n6 0.189894
R134 VP.n23 VP.n22 0.189894
R135 VP.n23 VP.n4 0.189894
R136 VP.n27 VP.n4 0.189894
R137 VP.n28 VP.n27 0.189894
R138 VP.n29 VP.n28 0.189894
R139 VP.n29 VP.n2 0.189894
R140 VP.n33 VP.n2 0.189894
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n0 0.189894
R144 VP VP.n39 0.153422
R145 VDD1 VDD1.t2 132.421
R146 VDD1.n1 VDD1.t5 132.306
R147 VDD1.n1 VDD1.n0 121.995
R148 VDD1.n3 VDD1.n2 121.46
R149 VDD1.n3 VDD1.n1 36.225
R150 VDD1.n2 VDD1.t4 9.13112
R151 VDD1.n2 VDD1.t3 9.13112
R152 VDD1.n0 VDD1.t1 9.13112
R153 VDD1.n0 VDD1.t0 9.13112
R154 VDD1 VDD1.n3 0.532828
R155 B.n259 B.n258 585
R156 B.n257 B.n90 585
R157 B.n256 B.n255 585
R158 B.n254 B.n91 585
R159 B.n253 B.n252 585
R160 B.n251 B.n92 585
R161 B.n250 B.n249 585
R162 B.n248 B.n93 585
R163 B.n247 B.n246 585
R164 B.n245 B.n94 585
R165 B.n244 B.n243 585
R166 B.n242 B.n95 585
R167 B.n241 B.n240 585
R168 B.n239 B.n96 585
R169 B.n238 B.n237 585
R170 B.n236 B.n97 585
R171 B.n235 B.n234 585
R172 B.n232 B.n98 585
R173 B.n231 B.n230 585
R174 B.n229 B.n101 585
R175 B.n228 B.n227 585
R176 B.n226 B.n102 585
R177 B.n225 B.n224 585
R178 B.n223 B.n103 585
R179 B.n222 B.n221 585
R180 B.n220 B.n104 585
R181 B.n218 B.n217 585
R182 B.n216 B.n107 585
R183 B.n215 B.n214 585
R184 B.n213 B.n108 585
R185 B.n212 B.n211 585
R186 B.n210 B.n109 585
R187 B.n209 B.n208 585
R188 B.n207 B.n110 585
R189 B.n206 B.n205 585
R190 B.n204 B.n111 585
R191 B.n203 B.n202 585
R192 B.n201 B.n112 585
R193 B.n200 B.n199 585
R194 B.n198 B.n113 585
R195 B.n197 B.n196 585
R196 B.n195 B.n114 585
R197 B.n194 B.n193 585
R198 B.n260 B.n89 585
R199 B.n262 B.n261 585
R200 B.n263 B.n88 585
R201 B.n265 B.n264 585
R202 B.n266 B.n87 585
R203 B.n268 B.n267 585
R204 B.n269 B.n86 585
R205 B.n271 B.n270 585
R206 B.n272 B.n85 585
R207 B.n274 B.n273 585
R208 B.n275 B.n84 585
R209 B.n277 B.n276 585
R210 B.n278 B.n83 585
R211 B.n280 B.n279 585
R212 B.n281 B.n82 585
R213 B.n283 B.n282 585
R214 B.n284 B.n81 585
R215 B.n286 B.n285 585
R216 B.n287 B.n80 585
R217 B.n289 B.n288 585
R218 B.n290 B.n79 585
R219 B.n292 B.n291 585
R220 B.n293 B.n78 585
R221 B.n295 B.n294 585
R222 B.n296 B.n77 585
R223 B.n298 B.n297 585
R224 B.n299 B.n76 585
R225 B.n301 B.n300 585
R226 B.n302 B.n75 585
R227 B.n304 B.n303 585
R228 B.n305 B.n74 585
R229 B.n307 B.n306 585
R230 B.n308 B.n73 585
R231 B.n310 B.n309 585
R232 B.n311 B.n72 585
R233 B.n313 B.n312 585
R234 B.n314 B.n71 585
R235 B.n316 B.n315 585
R236 B.n317 B.n70 585
R237 B.n319 B.n318 585
R238 B.n320 B.n69 585
R239 B.n322 B.n321 585
R240 B.n323 B.n68 585
R241 B.n325 B.n324 585
R242 B.n326 B.n67 585
R243 B.n328 B.n327 585
R244 B.n329 B.n66 585
R245 B.n331 B.n330 585
R246 B.n332 B.n65 585
R247 B.n334 B.n333 585
R248 B.n335 B.n64 585
R249 B.n337 B.n336 585
R250 B.n338 B.n63 585
R251 B.n340 B.n339 585
R252 B.n341 B.n62 585
R253 B.n343 B.n342 585
R254 B.n344 B.n61 585
R255 B.n346 B.n345 585
R256 B.n347 B.n60 585
R257 B.n349 B.n348 585
R258 B.n350 B.n59 585
R259 B.n352 B.n351 585
R260 B.n353 B.n58 585
R261 B.n355 B.n354 585
R262 B.n356 B.n57 585
R263 B.n358 B.n357 585
R264 B.n359 B.n56 585
R265 B.n361 B.n360 585
R266 B.n362 B.n55 585
R267 B.n364 B.n363 585
R268 B.n365 B.n54 585
R269 B.n367 B.n366 585
R270 B.n368 B.n53 585
R271 B.n370 B.n369 585
R272 B.n371 B.n52 585
R273 B.n373 B.n372 585
R274 B.n374 B.n51 585
R275 B.n376 B.n375 585
R276 B.n377 B.n50 585
R277 B.n379 B.n378 585
R278 B.n380 B.n49 585
R279 B.n382 B.n381 585
R280 B.n447 B.n22 585
R281 B.n446 B.n445 585
R282 B.n444 B.n23 585
R283 B.n443 B.n442 585
R284 B.n441 B.n24 585
R285 B.n440 B.n439 585
R286 B.n438 B.n25 585
R287 B.n437 B.n436 585
R288 B.n435 B.n26 585
R289 B.n434 B.n433 585
R290 B.n432 B.n27 585
R291 B.n431 B.n430 585
R292 B.n429 B.n28 585
R293 B.n428 B.n427 585
R294 B.n426 B.n29 585
R295 B.n425 B.n424 585
R296 B.n423 B.n30 585
R297 B.n422 B.n421 585
R298 B.n420 B.n31 585
R299 B.n419 B.n418 585
R300 B.n417 B.n35 585
R301 B.n416 B.n415 585
R302 B.n414 B.n36 585
R303 B.n413 B.n412 585
R304 B.n411 B.n37 585
R305 B.n410 B.n409 585
R306 B.n407 B.n38 585
R307 B.n406 B.n405 585
R308 B.n404 B.n41 585
R309 B.n403 B.n402 585
R310 B.n401 B.n42 585
R311 B.n400 B.n399 585
R312 B.n398 B.n43 585
R313 B.n397 B.n396 585
R314 B.n395 B.n44 585
R315 B.n394 B.n393 585
R316 B.n392 B.n45 585
R317 B.n391 B.n390 585
R318 B.n389 B.n46 585
R319 B.n388 B.n387 585
R320 B.n386 B.n47 585
R321 B.n385 B.n384 585
R322 B.n383 B.n48 585
R323 B.n449 B.n448 585
R324 B.n450 B.n21 585
R325 B.n452 B.n451 585
R326 B.n453 B.n20 585
R327 B.n455 B.n454 585
R328 B.n456 B.n19 585
R329 B.n458 B.n457 585
R330 B.n459 B.n18 585
R331 B.n461 B.n460 585
R332 B.n462 B.n17 585
R333 B.n464 B.n463 585
R334 B.n465 B.n16 585
R335 B.n467 B.n466 585
R336 B.n468 B.n15 585
R337 B.n470 B.n469 585
R338 B.n471 B.n14 585
R339 B.n473 B.n472 585
R340 B.n474 B.n13 585
R341 B.n476 B.n475 585
R342 B.n477 B.n12 585
R343 B.n479 B.n478 585
R344 B.n480 B.n11 585
R345 B.n482 B.n481 585
R346 B.n483 B.n10 585
R347 B.n485 B.n484 585
R348 B.n486 B.n9 585
R349 B.n488 B.n487 585
R350 B.n489 B.n8 585
R351 B.n491 B.n490 585
R352 B.n492 B.n7 585
R353 B.n494 B.n493 585
R354 B.n495 B.n6 585
R355 B.n497 B.n496 585
R356 B.n498 B.n5 585
R357 B.n500 B.n499 585
R358 B.n501 B.n4 585
R359 B.n503 B.n502 585
R360 B.n504 B.n3 585
R361 B.n506 B.n505 585
R362 B.n507 B.n0 585
R363 B.n2 B.n1 585
R364 B.n135 B.n134 585
R365 B.n137 B.n136 585
R366 B.n138 B.n133 585
R367 B.n140 B.n139 585
R368 B.n141 B.n132 585
R369 B.n143 B.n142 585
R370 B.n144 B.n131 585
R371 B.n146 B.n145 585
R372 B.n147 B.n130 585
R373 B.n149 B.n148 585
R374 B.n150 B.n129 585
R375 B.n152 B.n151 585
R376 B.n153 B.n128 585
R377 B.n155 B.n154 585
R378 B.n156 B.n127 585
R379 B.n158 B.n157 585
R380 B.n159 B.n126 585
R381 B.n161 B.n160 585
R382 B.n162 B.n125 585
R383 B.n164 B.n163 585
R384 B.n165 B.n124 585
R385 B.n167 B.n166 585
R386 B.n168 B.n123 585
R387 B.n170 B.n169 585
R388 B.n171 B.n122 585
R389 B.n173 B.n172 585
R390 B.n174 B.n121 585
R391 B.n176 B.n175 585
R392 B.n177 B.n120 585
R393 B.n179 B.n178 585
R394 B.n180 B.n119 585
R395 B.n182 B.n181 585
R396 B.n183 B.n118 585
R397 B.n185 B.n184 585
R398 B.n186 B.n117 585
R399 B.n188 B.n187 585
R400 B.n189 B.n116 585
R401 B.n191 B.n190 585
R402 B.n192 B.n115 585
R403 B.n193 B.n192 487.695
R404 B.n260 B.n259 487.695
R405 B.n381 B.n48 487.695
R406 B.n448 B.n447 487.695
R407 B.n509 B.n508 256.663
R408 B.n99 B.t3 244
R409 B.n39 B.t9 244
R410 B.n105 B.t6 243.655
R411 B.n32 B.t0 243.655
R412 B.n508 B.n507 235.042
R413 B.n508 B.n2 235.042
R414 B.n99 B.t4 182.636
R415 B.n39 B.t11 182.636
R416 B.n105 B.t7 182.632
R417 B.n32 B.t2 182.632
R418 B.n193 B.n114 163.367
R419 B.n197 B.n114 163.367
R420 B.n198 B.n197 163.367
R421 B.n199 B.n198 163.367
R422 B.n199 B.n112 163.367
R423 B.n203 B.n112 163.367
R424 B.n204 B.n203 163.367
R425 B.n205 B.n204 163.367
R426 B.n205 B.n110 163.367
R427 B.n209 B.n110 163.367
R428 B.n210 B.n209 163.367
R429 B.n211 B.n210 163.367
R430 B.n211 B.n108 163.367
R431 B.n215 B.n108 163.367
R432 B.n216 B.n215 163.367
R433 B.n217 B.n216 163.367
R434 B.n217 B.n104 163.367
R435 B.n222 B.n104 163.367
R436 B.n223 B.n222 163.367
R437 B.n224 B.n223 163.367
R438 B.n224 B.n102 163.367
R439 B.n228 B.n102 163.367
R440 B.n229 B.n228 163.367
R441 B.n230 B.n229 163.367
R442 B.n230 B.n98 163.367
R443 B.n235 B.n98 163.367
R444 B.n236 B.n235 163.367
R445 B.n237 B.n236 163.367
R446 B.n237 B.n96 163.367
R447 B.n241 B.n96 163.367
R448 B.n242 B.n241 163.367
R449 B.n243 B.n242 163.367
R450 B.n243 B.n94 163.367
R451 B.n247 B.n94 163.367
R452 B.n248 B.n247 163.367
R453 B.n249 B.n248 163.367
R454 B.n249 B.n92 163.367
R455 B.n253 B.n92 163.367
R456 B.n254 B.n253 163.367
R457 B.n255 B.n254 163.367
R458 B.n255 B.n90 163.367
R459 B.n259 B.n90 163.367
R460 B.n381 B.n380 163.367
R461 B.n380 B.n379 163.367
R462 B.n379 B.n50 163.367
R463 B.n375 B.n50 163.367
R464 B.n375 B.n374 163.367
R465 B.n374 B.n373 163.367
R466 B.n373 B.n52 163.367
R467 B.n369 B.n52 163.367
R468 B.n369 B.n368 163.367
R469 B.n368 B.n367 163.367
R470 B.n367 B.n54 163.367
R471 B.n363 B.n54 163.367
R472 B.n363 B.n362 163.367
R473 B.n362 B.n361 163.367
R474 B.n361 B.n56 163.367
R475 B.n357 B.n56 163.367
R476 B.n357 B.n356 163.367
R477 B.n356 B.n355 163.367
R478 B.n355 B.n58 163.367
R479 B.n351 B.n58 163.367
R480 B.n351 B.n350 163.367
R481 B.n350 B.n349 163.367
R482 B.n349 B.n60 163.367
R483 B.n345 B.n60 163.367
R484 B.n345 B.n344 163.367
R485 B.n344 B.n343 163.367
R486 B.n343 B.n62 163.367
R487 B.n339 B.n62 163.367
R488 B.n339 B.n338 163.367
R489 B.n338 B.n337 163.367
R490 B.n337 B.n64 163.367
R491 B.n333 B.n64 163.367
R492 B.n333 B.n332 163.367
R493 B.n332 B.n331 163.367
R494 B.n331 B.n66 163.367
R495 B.n327 B.n66 163.367
R496 B.n327 B.n326 163.367
R497 B.n326 B.n325 163.367
R498 B.n325 B.n68 163.367
R499 B.n321 B.n68 163.367
R500 B.n321 B.n320 163.367
R501 B.n320 B.n319 163.367
R502 B.n319 B.n70 163.367
R503 B.n315 B.n70 163.367
R504 B.n315 B.n314 163.367
R505 B.n314 B.n313 163.367
R506 B.n313 B.n72 163.367
R507 B.n309 B.n72 163.367
R508 B.n309 B.n308 163.367
R509 B.n308 B.n307 163.367
R510 B.n307 B.n74 163.367
R511 B.n303 B.n74 163.367
R512 B.n303 B.n302 163.367
R513 B.n302 B.n301 163.367
R514 B.n301 B.n76 163.367
R515 B.n297 B.n76 163.367
R516 B.n297 B.n296 163.367
R517 B.n296 B.n295 163.367
R518 B.n295 B.n78 163.367
R519 B.n291 B.n78 163.367
R520 B.n291 B.n290 163.367
R521 B.n290 B.n289 163.367
R522 B.n289 B.n80 163.367
R523 B.n285 B.n80 163.367
R524 B.n285 B.n284 163.367
R525 B.n284 B.n283 163.367
R526 B.n283 B.n82 163.367
R527 B.n279 B.n82 163.367
R528 B.n279 B.n278 163.367
R529 B.n278 B.n277 163.367
R530 B.n277 B.n84 163.367
R531 B.n273 B.n84 163.367
R532 B.n273 B.n272 163.367
R533 B.n272 B.n271 163.367
R534 B.n271 B.n86 163.367
R535 B.n267 B.n86 163.367
R536 B.n267 B.n266 163.367
R537 B.n266 B.n265 163.367
R538 B.n265 B.n88 163.367
R539 B.n261 B.n88 163.367
R540 B.n261 B.n260 163.367
R541 B.n447 B.n446 163.367
R542 B.n446 B.n23 163.367
R543 B.n442 B.n23 163.367
R544 B.n442 B.n441 163.367
R545 B.n441 B.n440 163.367
R546 B.n440 B.n25 163.367
R547 B.n436 B.n25 163.367
R548 B.n436 B.n435 163.367
R549 B.n435 B.n434 163.367
R550 B.n434 B.n27 163.367
R551 B.n430 B.n27 163.367
R552 B.n430 B.n429 163.367
R553 B.n429 B.n428 163.367
R554 B.n428 B.n29 163.367
R555 B.n424 B.n29 163.367
R556 B.n424 B.n423 163.367
R557 B.n423 B.n422 163.367
R558 B.n422 B.n31 163.367
R559 B.n418 B.n31 163.367
R560 B.n418 B.n417 163.367
R561 B.n417 B.n416 163.367
R562 B.n416 B.n36 163.367
R563 B.n412 B.n36 163.367
R564 B.n412 B.n411 163.367
R565 B.n411 B.n410 163.367
R566 B.n410 B.n38 163.367
R567 B.n405 B.n38 163.367
R568 B.n405 B.n404 163.367
R569 B.n404 B.n403 163.367
R570 B.n403 B.n42 163.367
R571 B.n399 B.n42 163.367
R572 B.n399 B.n398 163.367
R573 B.n398 B.n397 163.367
R574 B.n397 B.n44 163.367
R575 B.n393 B.n44 163.367
R576 B.n393 B.n392 163.367
R577 B.n392 B.n391 163.367
R578 B.n391 B.n46 163.367
R579 B.n387 B.n46 163.367
R580 B.n387 B.n386 163.367
R581 B.n386 B.n385 163.367
R582 B.n385 B.n48 163.367
R583 B.n448 B.n21 163.367
R584 B.n452 B.n21 163.367
R585 B.n453 B.n452 163.367
R586 B.n454 B.n453 163.367
R587 B.n454 B.n19 163.367
R588 B.n458 B.n19 163.367
R589 B.n459 B.n458 163.367
R590 B.n460 B.n459 163.367
R591 B.n460 B.n17 163.367
R592 B.n464 B.n17 163.367
R593 B.n465 B.n464 163.367
R594 B.n466 B.n465 163.367
R595 B.n466 B.n15 163.367
R596 B.n470 B.n15 163.367
R597 B.n471 B.n470 163.367
R598 B.n472 B.n471 163.367
R599 B.n472 B.n13 163.367
R600 B.n476 B.n13 163.367
R601 B.n477 B.n476 163.367
R602 B.n478 B.n477 163.367
R603 B.n478 B.n11 163.367
R604 B.n482 B.n11 163.367
R605 B.n483 B.n482 163.367
R606 B.n484 B.n483 163.367
R607 B.n484 B.n9 163.367
R608 B.n488 B.n9 163.367
R609 B.n489 B.n488 163.367
R610 B.n490 B.n489 163.367
R611 B.n490 B.n7 163.367
R612 B.n494 B.n7 163.367
R613 B.n495 B.n494 163.367
R614 B.n496 B.n495 163.367
R615 B.n496 B.n5 163.367
R616 B.n500 B.n5 163.367
R617 B.n501 B.n500 163.367
R618 B.n502 B.n501 163.367
R619 B.n502 B.n3 163.367
R620 B.n506 B.n3 163.367
R621 B.n507 B.n506 163.367
R622 B.n134 B.n2 163.367
R623 B.n137 B.n134 163.367
R624 B.n138 B.n137 163.367
R625 B.n139 B.n138 163.367
R626 B.n139 B.n132 163.367
R627 B.n143 B.n132 163.367
R628 B.n144 B.n143 163.367
R629 B.n145 B.n144 163.367
R630 B.n145 B.n130 163.367
R631 B.n149 B.n130 163.367
R632 B.n150 B.n149 163.367
R633 B.n151 B.n150 163.367
R634 B.n151 B.n128 163.367
R635 B.n155 B.n128 163.367
R636 B.n156 B.n155 163.367
R637 B.n157 B.n156 163.367
R638 B.n157 B.n126 163.367
R639 B.n161 B.n126 163.367
R640 B.n162 B.n161 163.367
R641 B.n163 B.n162 163.367
R642 B.n163 B.n124 163.367
R643 B.n167 B.n124 163.367
R644 B.n168 B.n167 163.367
R645 B.n169 B.n168 163.367
R646 B.n169 B.n122 163.367
R647 B.n173 B.n122 163.367
R648 B.n174 B.n173 163.367
R649 B.n175 B.n174 163.367
R650 B.n175 B.n120 163.367
R651 B.n179 B.n120 163.367
R652 B.n180 B.n179 163.367
R653 B.n181 B.n180 163.367
R654 B.n181 B.n118 163.367
R655 B.n185 B.n118 163.367
R656 B.n186 B.n185 163.367
R657 B.n187 B.n186 163.367
R658 B.n187 B.n116 163.367
R659 B.n191 B.n116 163.367
R660 B.n192 B.n191 163.367
R661 B.n100 B.t5 129.496
R662 B.n40 B.t10 129.496
R663 B.n106 B.t8 129.494
R664 B.n33 B.t1 129.494
R665 B.n219 B.n106 59.5399
R666 B.n233 B.n100 59.5399
R667 B.n408 B.n40 59.5399
R668 B.n34 B.n33 59.5399
R669 B.n106 B.n105 53.1399
R670 B.n100 B.n99 53.1399
R671 B.n40 B.n39 53.1399
R672 B.n33 B.n32 53.1399
R673 B.n449 B.n22 31.6883
R674 B.n383 B.n382 31.6883
R675 B.n258 B.n89 31.6883
R676 B.n194 B.n115 31.6883
R677 B B.n509 18.0485
R678 B.n450 B.n449 10.6151
R679 B.n451 B.n450 10.6151
R680 B.n451 B.n20 10.6151
R681 B.n455 B.n20 10.6151
R682 B.n456 B.n455 10.6151
R683 B.n457 B.n456 10.6151
R684 B.n457 B.n18 10.6151
R685 B.n461 B.n18 10.6151
R686 B.n462 B.n461 10.6151
R687 B.n463 B.n462 10.6151
R688 B.n463 B.n16 10.6151
R689 B.n467 B.n16 10.6151
R690 B.n468 B.n467 10.6151
R691 B.n469 B.n468 10.6151
R692 B.n469 B.n14 10.6151
R693 B.n473 B.n14 10.6151
R694 B.n474 B.n473 10.6151
R695 B.n475 B.n474 10.6151
R696 B.n475 B.n12 10.6151
R697 B.n479 B.n12 10.6151
R698 B.n480 B.n479 10.6151
R699 B.n481 B.n480 10.6151
R700 B.n481 B.n10 10.6151
R701 B.n485 B.n10 10.6151
R702 B.n486 B.n485 10.6151
R703 B.n487 B.n486 10.6151
R704 B.n487 B.n8 10.6151
R705 B.n491 B.n8 10.6151
R706 B.n492 B.n491 10.6151
R707 B.n493 B.n492 10.6151
R708 B.n493 B.n6 10.6151
R709 B.n497 B.n6 10.6151
R710 B.n498 B.n497 10.6151
R711 B.n499 B.n498 10.6151
R712 B.n499 B.n4 10.6151
R713 B.n503 B.n4 10.6151
R714 B.n504 B.n503 10.6151
R715 B.n505 B.n504 10.6151
R716 B.n505 B.n0 10.6151
R717 B.n445 B.n22 10.6151
R718 B.n445 B.n444 10.6151
R719 B.n444 B.n443 10.6151
R720 B.n443 B.n24 10.6151
R721 B.n439 B.n24 10.6151
R722 B.n439 B.n438 10.6151
R723 B.n438 B.n437 10.6151
R724 B.n437 B.n26 10.6151
R725 B.n433 B.n26 10.6151
R726 B.n433 B.n432 10.6151
R727 B.n432 B.n431 10.6151
R728 B.n431 B.n28 10.6151
R729 B.n427 B.n28 10.6151
R730 B.n427 B.n426 10.6151
R731 B.n426 B.n425 10.6151
R732 B.n425 B.n30 10.6151
R733 B.n421 B.n420 10.6151
R734 B.n420 B.n419 10.6151
R735 B.n419 B.n35 10.6151
R736 B.n415 B.n35 10.6151
R737 B.n415 B.n414 10.6151
R738 B.n414 B.n413 10.6151
R739 B.n413 B.n37 10.6151
R740 B.n409 B.n37 10.6151
R741 B.n407 B.n406 10.6151
R742 B.n406 B.n41 10.6151
R743 B.n402 B.n41 10.6151
R744 B.n402 B.n401 10.6151
R745 B.n401 B.n400 10.6151
R746 B.n400 B.n43 10.6151
R747 B.n396 B.n43 10.6151
R748 B.n396 B.n395 10.6151
R749 B.n395 B.n394 10.6151
R750 B.n394 B.n45 10.6151
R751 B.n390 B.n45 10.6151
R752 B.n390 B.n389 10.6151
R753 B.n389 B.n388 10.6151
R754 B.n388 B.n47 10.6151
R755 B.n384 B.n47 10.6151
R756 B.n384 B.n383 10.6151
R757 B.n382 B.n49 10.6151
R758 B.n378 B.n49 10.6151
R759 B.n378 B.n377 10.6151
R760 B.n377 B.n376 10.6151
R761 B.n376 B.n51 10.6151
R762 B.n372 B.n51 10.6151
R763 B.n372 B.n371 10.6151
R764 B.n371 B.n370 10.6151
R765 B.n370 B.n53 10.6151
R766 B.n366 B.n53 10.6151
R767 B.n366 B.n365 10.6151
R768 B.n365 B.n364 10.6151
R769 B.n364 B.n55 10.6151
R770 B.n360 B.n55 10.6151
R771 B.n360 B.n359 10.6151
R772 B.n359 B.n358 10.6151
R773 B.n358 B.n57 10.6151
R774 B.n354 B.n57 10.6151
R775 B.n354 B.n353 10.6151
R776 B.n353 B.n352 10.6151
R777 B.n352 B.n59 10.6151
R778 B.n348 B.n59 10.6151
R779 B.n348 B.n347 10.6151
R780 B.n347 B.n346 10.6151
R781 B.n346 B.n61 10.6151
R782 B.n342 B.n61 10.6151
R783 B.n342 B.n341 10.6151
R784 B.n341 B.n340 10.6151
R785 B.n340 B.n63 10.6151
R786 B.n336 B.n63 10.6151
R787 B.n336 B.n335 10.6151
R788 B.n335 B.n334 10.6151
R789 B.n334 B.n65 10.6151
R790 B.n330 B.n65 10.6151
R791 B.n330 B.n329 10.6151
R792 B.n329 B.n328 10.6151
R793 B.n328 B.n67 10.6151
R794 B.n324 B.n67 10.6151
R795 B.n324 B.n323 10.6151
R796 B.n323 B.n322 10.6151
R797 B.n322 B.n69 10.6151
R798 B.n318 B.n69 10.6151
R799 B.n318 B.n317 10.6151
R800 B.n317 B.n316 10.6151
R801 B.n316 B.n71 10.6151
R802 B.n312 B.n71 10.6151
R803 B.n312 B.n311 10.6151
R804 B.n311 B.n310 10.6151
R805 B.n310 B.n73 10.6151
R806 B.n306 B.n73 10.6151
R807 B.n306 B.n305 10.6151
R808 B.n305 B.n304 10.6151
R809 B.n304 B.n75 10.6151
R810 B.n300 B.n75 10.6151
R811 B.n300 B.n299 10.6151
R812 B.n299 B.n298 10.6151
R813 B.n298 B.n77 10.6151
R814 B.n294 B.n77 10.6151
R815 B.n294 B.n293 10.6151
R816 B.n293 B.n292 10.6151
R817 B.n292 B.n79 10.6151
R818 B.n288 B.n79 10.6151
R819 B.n288 B.n287 10.6151
R820 B.n287 B.n286 10.6151
R821 B.n286 B.n81 10.6151
R822 B.n282 B.n81 10.6151
R823 B.n282 B.n281 10.6151
R824 B.n281 B.n280 10.6151
R825 B.n280 B.n83 10.6151
R826 B.n276 B.n83 10.6151
R827 B.n276 B.n275 10.6151
R828 B.n275 B.n274 10.6151
R829 B.n274 B.n85 10.6151
R830 B.n270 B.n85 10.6151
R831 B.n270 B.n269 10.6151
R832 B.n269 B.n268 10.6151
R833 B.n268 B.n87 10.6151
R834 B.n264 B.n87 10.6151
R835 B.n264 B.n263 10.6151
R836 B.n263 B.n262 10.6151
R837 B.n262 B.n89 10.6151
R838 B.n135 B.n1 10.6151
R839 B.n136 B.n135 10.6151
R840 B.n136 B.n133 10.6151
R841 B.n140 B.n133 10.6151
R842 B.n141 B.n140 10.6151
R843 B.n142 B.n141 10.6151
R844 B.n142 B.n131 10.6151
R845 B.n146 B.n131 10.6151
R846 B.n147 B.n146 10.6151
R847 B.n148 B.n147 10.6151
R848 B.n148 B.n129 10.6151
R849 B.n152 B.n129 10.6151
R850 B.n153 B.n152 10.6151
R851 B.n154 B.n153 10.6151
R852 B.n154 B.n127 10.6151
R853 B.n158 B.n127 10.6151
R854 B.n159 B.n158 10.6151
R855 B.n160 B.n159 10.6151
R856 B.n160 B.n125 10.6151
R857 B.n164 B.n125 10.6151
R858 B.n165 B.n164 10.6151
R859 B.n166 B.n165 10.6151
R860 B.n166 B.n123 10.6151
R861 B.n170 B.n123 10.6151
R862 B.n171 B.n170 10.6151
R863 B.n172 B.n171 10.6151
R864 B.n172 B.n121 10.6151
R865 B.n176 B.n121 10.6151
R866 B.n177 B.n176 10.6151
R867 B.n178 B.n177 10.6151
R868 B.n178 B.n119 10.6151
R869 B.n182 B.n119 10.6151
R870 B.n183 B.n182 10.6151
R871 B.n184 B.n183 10.6151
R872 B.n184 B.n117 10.6151
R873 B.n188 B.n117 10.6151
R874 B.n189 B.n188 10.6151
R875 B.n190 B.n189 10.6151
R876 B.n190 B.n115 10.6151
R877 B.n195 B.n194 10.6151
R878 B.n196 B.n195 10.6151
R879 B.n196 B.n113 10.6151
R880 B.n200 B.n113 10.6151
R881 B.n201 B.n200 10.6151
R882 B.n202 B.n201 10.6151
R883 B.n202 B.n111 10.6151
R884 B.n206 B.n111 10.6151
R885 B.n207 B.n206 10.6151
R886 B.n208 B.n207 10.6151
R887 B.n208 B.n109 10.6151
R888 B.n212 B.n109 10.6151
R889 B.n213 B.n212 10.6151
R890 B.n214 B.n213 10.6151
R891 B.n214 B.n107 10.6151
R892 B.n218 B.n107 10.6151
R893 B.n221 B.n220 10.6151
R894 B.n221 B.n103 10.6151
R895 B.n225 B.n103 10.6151
R896 B.n226 B.n225 10.6151
R897 B.n227 B.n226 10.6151
R898 B.n227 B.n101 10.6151
R899 B.n231 B.n101 10.6151
R900 B.n232 B.n231 10.6151
R901 B.n234 B.n97 10.6151
R902 B.n238 B.n97 10.6151
R903 B.n239 B.n238 10.6151
R904 B.n240 B.n239 10.6151
R905 B.n240 B.n95 10.6151
R906 B.n244 B.n95 10.6151
R907 B.n245 B.n244 10.6151
R908 B.n246 B.n245 10.6151
R909 B.n246 B.n93 10.6151
R910 B.n250 B.n93 10.6151
R911 B.n251 B.n250 10.6151
R912 B.n252 B.n251 10.6151
R913 B.n252 B.n91 10.6151
R914 B.n256 B.n91 10.6151
R915 B.n257 B.n256 10.6151
R916 B.n258 B.n257 10.6151
R917 B.n509 B.n0 8.11757
R918 B.n509 B.n1 8.11757
R919 B.n421 B.n34 6.4005
R920 B.n409 B.n408 6.4005
R921 B.n220 B.n219 6.4005
R922 B.n233 B.n232 6.4005
R923 B.n34 B.n30 4.21513
R924 B.n408 B.n407 4.21513
R925 B.n219 B.n218 4.21513
R926 B.n234 B.n233 4.21513
C0 VDD2 VTAIL 4.60505f
C1 VDD2 VP 0.44639f
C2 VN VTAIL 2.89686f
C3 VN VP 5.19063f
C4 VDD1 VTAIL 4.55359f
C5 VDD1 VP 2.52561f
C6 VTAIL w_n3162_n1680# 1.74506f
C7 B VTAIL 1.70948f
C8 VP w_n3162_n1680# 6.2108f
C9 B VP 1.71817f
C10 VDD2 VN 2.23636f
C11 VDD2 VDD1 1.332f
C12 VDD2 w_n3162_n1680# 1.73245f
C13 VDD2 B 1.44907f
C14 VDD1 VN 0.154779f
C15 VN w_n3162_n1680# 5.80399f
C16 B VN 1.03775f
C17 VDD1 w_n3162_n1680# 1.65384f
C18 VDD1 B 1.37936f
C19 B w_n3162_n1680# 7.079f
C20 VP VTAIL 2.91102f
C21 VDD2 VSUBS 1.27655f
C22 VDD1 VSUBS 1.729916f
C23 VTAIL VSUBS 0.544406f
C24 VN VSUBS 5.424531f
C25 VP VSUBS 2.278203f
C26 B VSUBS 3.523045f
C27 w_n3162_n1680# VSUBS 67.047005f
C28 B.n0 VSUBS 0.006487f
C29 B.n1 VSUBS 0.006487f
C30 B.n2 VSUBS 0.009593f
C31 B.n3 VSUBS 0.007352f
C32 B.n4 VSUBS 0.007352f
C33 B.n5 VSUBS 0.007352f
C34 B.n6 VSUBS 0.007352f
C35 B.n7 VSUBS 0.007352f
C36 B.n8 VSUBS 0.007352f
C37 B.n9 VSUBS 0.007352f
C38 B.n10 VSUBS 0.007352f
C39 B.n11 VSUBS 0.007352f
C40 B.n12 VSUBS 0.007352f
C41 B.n13 VSUBS 0.007352f
C42 B.n14 VSUBS 0.007352f
C43 B.n15 VSUBS 0.007352f
C44 B.n16 VSUBS 0.007352f
C45 B.n17 VSUBS 0.007352f
C46 B.n18 VSUBS 0.007352f
C47 B.n19 VSUBS 0.007352f
C48 B.n20 VSUBS 0.007352f
C49 B.n21 VSUBS 0.007352f
C50 B.n22 VSUBS 0.017116f
C51 B.n23 VSUBS 0.007352f
C52 B.n24 VSUBS 0.007352f
C53 B.n25 VSUBS 0.007352f
C54 B.n26 VSUBS 0.007352f
C55 B.n27 VSUBS 0.007352f
C56 B.n28 VSUBS 0.007352f
C57 B.n29 VSUBS 0.007352f
C58 B.n30 VSUBS 0.005135f
C59 B.n31 VSUBS 0.007352f
C60 B.t1 VSUBS 0.094906f
C61 B.t2 VSUBS 0.112218f
C62 B.t0 VSUBS 0.434265f
C63 B.n32 VSUBS 0.089972f
C64 B.n33 VSUBS 0.069986f
C65 B.n34 VSUBS 0.017033f
C66 B.n35 VSUBS 0.007352f
C67 B.n36 VSUBS 0.007352f
C68 B.n37 VSUBS 0.007352f
C69 B.n38 VSUBS 0.007352f
C70 B.t10 VSUBS 0.094906f
C71 B.t11 VSUBS 0.112218f
C72 B.t9 VSUBS 0.434298f
C73 B.n39 VSUBS 0.089939f
C74 B.n40 VSUBS 0.069986f
C75 B.n41 VSUBS 0.007352f
C76 B.n42 VSUBS 0.007352f
C77 B.n43 VSUBS 0.007352f
C78 B.n44 VSUBS 0.007352f
C79 B.n45 VSUBS 0.007352f
C80 B.n46 VSUBS 0.007352f
C81 B.n47 VSUBS 0.007352f
C82 B.n48 VSUBS 0.017116f
C83 B.n49 VSUBS 0.007352f
C84 B.n50 VSUBS 0.007352f
C85 B.n51 VSUBS 0.007352f
C86 B.n52 VSUBS 0.007352f
C87 B.n53 VSUBS 0.007352f
C88 B.n54 VSUBS 0.007352f
C89 B.n55 VSUBS 0.007352f
C90 B.n56 VSUBS 0.007352f
C91 B.n57 VSUBS 0.007352f
C92 B.n58 VSUBS 0.007352f
C93 B.n59 VSUBS 0.007352f
C94 B.n60 VSUBS 0.007352f
C95 B.n61 VSUBS 0.007352f
C96 B.n62 VSUBS 0.007352f
C97 B.n63 VSUBS 0.007352f
C98 B.n64 VSUBS 0.007352f
C99 B.n65 VSUBS 0.007352f
C100 B.n66 VSUBS 0.007352f
C101 B.n67 VSUBS 0.007352f
C102 B.n68 VSUBS 0.007352f
C103 B.n69 VSUBS 0.007352f
C104 B.n70 VSUBS 0.007352f
C105 B.n71 VSUBS 0.007352f
C106 B.n72 VSUBS 0.007352f
C107 B.n73 VSUBS 0.007352f
C108 B.n74 VSUBS 0.007352f
C109 B.n75 VSUBS 0.007352f
C110 B.n76 VSUBS 0.007352f
C111 B.n77 VSUBS 0.007352f
C112 B.n78 VSUBS 0.007352f
C113 B.n79 VSUBS 0.007352f
C114 B.n80 VSUBS 0.007352f
C115 B.n81 VSUBS 0.007352f
C116 B.n82 VSUBS 0.007352f
C117 B.n83 VSUBS 0.007352f
C118 B.n84 VSUBS 0.007352f
C119 B.n85 VSUBS 0.007352f
C120 B.n86 VSUBS 0.007352f
C121 B.n87 VSUBS 0.007352f
C122 B.n88 VSUBS 0.007352f
C123 B.n89 VSUBS 0.01751f
C124 B.n90 VSUBS 0.007352f
C125 B.n91 VSUBS 0.007352f
C126 B.n92 VSUBS 0.007352f
C127 B.n93 VSUBS 0.007352f
C128 B.n94 VSUBS 0.007352f
C129 B.n95 VSUBS 0.007352f
C130 B.n96 VSUBS 0.007352f
C131 B.n97 VSUBS 0.007352f
C132 B.n98 VSUBS 0.007352f
C133 B.t5 VSUBS 0.094906f
C134 B.t4 VSUBS 0.112218f
C135 B.t3 VSUBS 0.434298f
C136 B.n99 VSUBS 0.089939f
C137 B.n100 VSUBS 0.069986f
C138 B.n101 VSUBS 0.007352f
C139 B.n102 VSUBS 0.007352f
C140 B.n103 VSUBS 0.007352f
C141 B.n104 VSUBS 0.007352f
C142 B.t8 VSUBS 0.094906f
C143 B.t7 VSUBS 0.112218f
C144 B.t6 VSUBS 0.434265f
C145 B.n105 VSUBS 0.089972f
C146 B.n106 VSUBS 0.069986f
C147 B.n107 VSUBS 0.007352f
C148 B.n108 VSUBS 0.007352f
C149 B.n109 VSUBS 0.007352f
C150 B.n110 VSUBS 0.007352f
C151 B.n111 VSUBS 0.007352f
C152 B.n112 VSUBS 0.007352f
C153 B.n113 VSUBS 0.007352f
C154 B.n114 VSUBS 0.007352f
C155 B.n115 VSUBS 0.016614f
C156 B.n116 VSUBS 0.007352f
C157 B.n117 VSUBS 0.007352f
C158 B.n118 VSUBS 0.007352f
C159 B.n119 VSUBS 0.007352f
C160 B.n120 VSUBS 0.007352f
C161 B.n121 VSUBS 0.007352f
C162 B.n122 VSUBS 0.007352f
C163 B.n123 VSUBS 0.007352f
C164 B.n124 VSUBS 0.007352f
C165 B.n125 VSUBS 0.007352f
C166 B.n126 VSUBS 0.007352f
C167 B.n127 VSUBS 0.007352f
C168 B.n128 VSUBS 0.007352f
C169 B.n129 VSUBS 0.007352f
C170 B.n130 VSUBS 0.007352f
C171 B.n131 VSUBS 0.007352f
C172 B.n132 VSUBS 0.007352f
C173 B.n133 VSUBS 0.007352f
C174 B.n134 VSUBS 0.007352f
C175 B.n135 VSUBS 0.007352f
C176 B.n136 VSUBS 0.007352f
C177 B.n137 VSUBS 0.007352f
C178 B.n138 VSUBS 0.007352f
C179 B.n139 VSUBS 0.007352f
C180 B.n140 VSUBS 0.007352f
C181 B.n141 VSUBS 0.007352f
C182 B.n142 VSUBS 0.007352f
C183 B.n143 VSUBS 0.007352f
C184 B.n144 VSUBS 0.007352f
C185 B.n145 VSUBS 0.007352f
C186 B.n146 VSUBS 0.007352f
C187 B.n147 VSUBS 0.007352f
C188 B.n148 VSUBS 0.007352f
C189 B.n149 VSUBS 0.007352f
C190 B.n150 VSUBS 0.007352f
C191 B.n151 VSUBS 0.007352f
C192 B.n152 VSUBS 0.007352f
C193 B.n153 VSUBS 0.007352f
C194 B.n154 VSUBS 0.007352f
C195 B.n155 VSUBS 0.007352f
C196 B.n156 VSUBS 0.007352f
C197 B.n157 VSUBS 0.007352f
C198 B.n158 VSUBS 0.007352f
C199 B.n159 VSUBS 0.007352f
C200 B.n160 VSUBS 0.007352f
C201 B.n161 VSUBS 0.007352f
C202 B.n162 VSUBS 0.007352f
C203 B.n163 VSUBS 0.007352f
C204 B.n164 VSUBS 0.007352f
C205 B.n165 VSUBS 0.007352f
C206 B.n166 VSUBS 0.007352f
C207 B.n167 VSUBS 0.007352f
C208 B.n168 VSUBS 0.007352f
C209 B.n169 VSUBS 0.007352f
C210 B.n170 VSUBS 0.007352f
C211 B.n171 VSUBS 0.007352f
C212 B.n172 VSUBS 0.007352f
C213 B.n173 VSUBS 0.007352f
C214 B.n174 VSUBS 0.007352f
C215 B.n175 VSUBS 0.007352f
C216 B.n176 VSUBS 0.007352f
C217 B.n177 VSUBS 0.007352f
C218 B.n178 VSUBS 0.007352f
C219 B.n179 VSUBS 0.007352f
C220 B.n180 VSUBS 0.007352f
C221 B.n181 VSUBS 0.007352f
C222 B.n182 VSUBS 0.007352f
C223 B.n183 VSUBS 0.007352f
C224 B.n184 VSUBS 0.007352f
C225 B.n185 VSUBS 0.007352f
C226 B.n186 VSUBS 0.007352f
C227 B.n187 VSUBS 0.007352f
C228 B.n188 VSUBS 0.007352f
C229 B.n189 VSUBS 0.007352f
C230 B.n190 VSUBS 0.007352f
C231 B.n191 VSUBS 0.007352f
C232 B.n192 VSUBS 0.016614f
C233 B.n193 VSUBS 0.017116f
C234 B.n194 VSUBS 0.017116f
C235 B.n195 VSUBS 0.007352f
C236 B.n196 VSUBS 0.007352f
C237 B.n197 VSUBS 0.007352f
C238 B.n198 VSUBS 0.007352f
C239 B.n199 VSUBS 0.007352f
C240 B.n200 VSUBS 0.007352f
C241 B.n201 VSUBS 0.007352f
C242 B.n202 VSUBS 0.007352f
C243 B.n203 VSUBS 0.007352f
C244 B.n204 VSUBS 0.007352f
C245 B.n205 VSUBS 0.007352f
C246 B.n206 VSUBS 0.007352f
C247 B.n207 VSUBS 0.007352f
C248 B.n208 VSUBS 0.007352f
C249 B.n209 VSUBS 0.007352f
C250 B.n210 VSUBS 0.007352f
C251 B.n211 VSUBS 0.007352f
C252 B.n212 VSUBS 0.007352f
C253 B.n213 VSUBS 0.007352f
C254 B.n214 VSUBS 0.007352f
C255 B.n215 VSUBS 0.007352f
C256 B.n216 VSUBS 0.007352f
C257 B.n217 VSUBS 0.007352f
C258 B.n218 VSUBS 0.005135f
C259 B.n219 VSUBS 0.017033f
C260 B.n220 VSUBS 0.005892f
C261 B.n221 VSUBS 0.007352f
C262 B.n222 VSUBS 0.007352f
C263 B.n223 VSUBS 0.007352f
C264 B.n224 VSUBS 0.007352f
C265 B.n225 VSUBS 0.007352f
C266 B.n226 VSUBS 0.007352f
C267 B.n227 VSUBS 0.007352f
C268 B.n228 VSUBS 0.007352f
C269 B.n229 VSUBS 0.007352f
C270 B.n230 VSUBS 0.007352f
C271 B.n231 VSUBS 0.007352f
C272 B.n232 VSUBS 0.005892f
C273 B.n233 VSUBS 0.017033f
C274 B.n234 VSUBS 0.005135f
C275 B.n235 VSUBS 0.007352f
C276 B.n236 VSUBS 0.007352f
C277 B.n237 VSUBS 0.007352f
C278 B.n238 VSUBS 0.007352f
C279 B.n239 VSUBS 0.007352f
C280 B.n240 VSUBS 0.007352f
C281 B.n241 VSUBS 0.007352f
C282 B.n242 VSUBS 0.007352f
C283 B.n243 VSUBS 0.007352f
C284 B.n244 VSUBS 0.007352f
C285 B.n245 VSUBS 0.007352f
C286 B.n246 VSUBS 0.007352f
C287 B.n247 VSUBS 0.007352f
C288 B.n248 VSUBS 0.007352f
C289 B.n249 VSUBS 0.007352f
C290 B.n250 VSUBS 0.007352f
C291 B.n251 VSUBS 0.007352f
C292 B.n252 VSUBS 0.007352f
C293 B.n253 VSUBS 0.007352f
C294 B.n254 VSUBS 0.007352f
C295 B.n255 VSUBS 0.007352f
C296 B.n256 VSUBS 0.007352f
C297 B.n257 VSUBS 0.007352f
C298 B.n258 VSUBS 0.016221f
C299 B.n259 VSUBS 0.017116f
C300 B.n260 VSUBS 0.016614f
C301 B.n261 VSUBS 0.007352f
C302 B.n262 VSUBS 0.007352f
C303 B.n263 VSUBS 0.007352f
C304 B.n264 VSUBS 0.007352f
C305 B.n265 VSUBS 0.007352f
C306 B.n266 VSUBS 0.007352f
C307 B.n267 VSUBS 0.007352f
C308 B.n268 VSUBS 0.007352f
C309 B.n269 VSUBS 0.007352f
C310 B.n270 VSUBS 0.007352f
C311 B.n271 VSUBS 0.007352f
C312 B.n272 VSUBS 0.007352f
C313 B.n273 VSUBS 0.007352f
C314 B.n274 VSUBS 0.007352f
C315 B.n275 VSUBS 0.007352f
C316 B.n276 VSUBS 0.007352f
C317 B.n277 VSUBS 0.007352f
C318 B.n278 VSUBS 0.007352f
C319 B.n279 VSUBS 0.007352f
C320 B.n280 VSUBS 0.007352f
C321 B.n281 VSUBS 0.007352f
C322 B.n282 VSUBS 0.007352f
C323 B.n283 VSUBS 0.007352f
C324 B.n284 VSUBS 0.007352f
C325 B.n285 VSUBS 0.007352f
C326 B.n286 VSUBS 0.007352f
C327 B.n287 VSUBS 0.007352f
C328 B.n288 VSUBS 0.007352f
C329 B.n289 VSUBS 0.007352f
C330 B.n290 VSUBS 0.007352f
C331 B.n291 VSUBS 0.007352f
C332 B.n292 VSUBS 0.007352f
C333 B.n293 VSUBS 0.007352f
C334 B.n294 VSUBS 0.007352f
C335 B.n295 VSUBS 0.007352f
C336 B.n296 VSUBS 0.007352f
C337 B.n297 VSUBS 0.007352f
C338 B.n298 VSUBS 0.007352f
C339 B.n299 VSUBS 0.007352f
C340 B.n300 VSUBS 0.007352f
C341 B.n301 VSUBS 0.007352f
C342 B.n302 VSUBS 0.007352f
C343 B.n303 VSUBS 0.007352f
C344 B.n304 VSUBS 0.007352f
C345 B.n305 VSUBS 0.007352f
C346 B.n306 VSUBS 0.007352f
C347 B.n307 VSUBS 0.007352f
C348 B.n308 VSUBS 0.007352f
C349 B.n309 VSUBS 0.007352f
C350 B.n310 VSUBS 0.007352f
C351 B.n311 VSUBS 0.007352f
C352 B.n312 VSUBS 0.007352f
C353 B.n313 VSUBS 0.007352f
C354 B.n314 VSUBS 0.007352f
C355 B.n315 VSUBS 0.007352f
C356 B.n316 VSUBS 0.007352f
C357 B.n317 VSUBS 0.007352f
C358 B.n318 VSUBS 0.007352f
C359 B.n319 VSUBS 0.007352f
C360 B.n320 VSUBS 0.007352f
C361 B.n321 VSUBS 0.007352f
C362 B.n322 VSUBS 0.007352f
C363 B.n323 VSUBS 0.007352f
C364 B.n324 VSUBS 0.007352f
C365 B.n325 VSUBS 0.007352f
C366 B.n326 VSUBS 0.007352f
C367 B.n327 VSUBS 0.007352f
C368 B.n328 VSUBS 0.007352f
C369 B.n329 VSUBS 0.007352f
C370 B.n330 VSUBS 0.007352f
C371 B.n331 VSUBS 0.007352f
C372 B.n332 VSUBS 0.007352f
C373 B.n333 VSUBS 0.007352f
C374 B.n334 VSUBS 0.007352f
C375 B.n335 VSUBS 0.007352f
C376 B.n336 VSUBS 0.007352f
C377 B.n337 VSUBS 0.007352f
C378 B.n338 VSUBS 0.007352f
C379 B.n339 VSUBS 0.007352f
C380 B.n340 VSUBS 0.007352f
C381 B.n341 VSUBS 0.007352f
C382 B.n342 VSUBS 0.007352f
C383 B.n343 VSUBS 0.007352f
C384 B.n344 VSUBS 0.007352f
C385 B.n345 VSUBS 0.007352f
C386 B.n346 VSUBS 0.007352f
C387 B.n347 VSUBS 0.007352f
C388 B.n348 VSUBS 0.007352f
C389 B.n349 VSUBS 0.007352f
C390 B.n350 VSUBS 0.007352f
C391 B.n351 VSUBS 0.007352f
C392 B.n352 VSUBS 0.007352f
C393 B.n353 VSUBS 0.007352f
C394 B.n354 VSUBS 0.007352f
C395 B.n355 VSUBS 0.007352f
C396 B.n356 VSUBS 0.007352f
C397 B.n357 VSUBS 0.007352f
C398 B.n358 VSUBS 0.007352f
C399 B.n359 VSUBS 0.007352f
C400 B.n360 VSUBS 0.007352f
C401 B.n361 VSUBS 0.007352f
C402 B.n362 VSUBS 0.007352f
C403 B.n363 VSUBS 0.007352f
C404 B.n364 VSUBS 0.007352f
C405 B.n365 VSUBS 0.007352f
C406 B.n366 VSUBS 0.007352f
C407 B.n367 VSUBS 0.007352f
C408 B.n368 VSUBS 0.007352f
C409 B.n369 VSUBS 0.007352f
C410 B.n370 VSUBS 0.007352f
C411 B.n371 VSUBS 0.007352f
C412 B.n372 VSUBS 0.007352f
C413 B.n373 VSUBS 0.007352f
C414 B.n374 VSUBS 0.007352f
C415 B.n375 VSUBS 0.007352f
C416 B.n376 VSUBS 0.007352f
C417 B.n377 VSUBS 0.007352f
C418 B.n378 VSUBS 0.007352f
C419 B.n379 VSUBS 0.007352f
C420 B.n380 VSUBS 0.007352f
C421 B.n381 VSUBS 0.016614f
C422 B.n382 VSUBS 0.016614f
C423 B.n383 VSUBS 0.017116f
C424 B.n384 VSUBS 0.007352f
C425 B.n385 VSUBS 0.007352f
C426 B.n386 VSUBS 0.007352f
C427 B.n387 VSUBS 0.007352f
C428 B.n388 VSUBS 0.007352f
C429 B.n389 VSUBS 0.007352f
C430 B.n390 VSUBS 0.007352f
C431 B.n391 VSUBS 0.007352f
C432 B.n392 VSUBS 0.007352f
C433 B.n393 VSUBS 0.007352f
C434 B.n394 VSUBS 0.007352f
C435 B.n395 VSUBS 0.007352f
C436 B.n396 VSUBS 0.007352f
C437 B.n397 VSUBS 0.007352f
C438 B.n398 VSUBS 0.007352f
C439 B.n399 VSUBS 0.007352f
C440 B.n400 VSUBS 0.007352f
C441 B.n401 VSUBS 0.007352f
C442 B.n402 VSUBS 0.007352f
C443 B.n403 VSUBS 0.007352f
C444 B.n404 VSUBS 0.007352f
C445 B.n405 VSUBS 0.007352f
C446 B.n406 VSUBS 0.007352f
C447 B.n407 VSUBS 0.005135f
C448 B.n408 VSUBS 0.017033f
C449 B.n409 VSUBS 0.005892f
C450 B.n410 VSUBS 0.007352f
C451 B.n411 VSUBS 0.007352f
C452 B.n412 VSUBS 0.007352f
C453 B.n413 VSUBS 0.007352f
C454 B.n414 VSUBS 0.007352f
C455 B.n415 VSUBS 0.007352f
C456 B.n416 VSUBS 0.007352f
C457 B.n417 VSUBS 0.007352f
C458 B.n418 VSUBS 0.007352f
C459 B.n419 VSUBS 0.007352f
C460 B.n420 VSUBS 0.007352f
C461 B.n421 VSUBS 0.005892f
C462 B.n422 VSUBS 0.007352f
C463 B.n423 VSUBS 0.007352f
C464 B.n424 VSUBS 0.007352f
C465 B.n425 VSUBS 0.007352f
C466 B.n426 VSUBS 0.007352f
C467 B.n427 VSUBS 0.007352f
C468 B.n428 VSUBS 0.007352f
C469 B.n429 VSUBS 0.007352f
C470 B.n430 VSUBS 0.007352f
C471 B.n431 VSUBS 0.007352f
C472 B.n432 VSUBS 0.007352f
C473 B.n433 VSUBS 0.007352f
C474 B.n434 VSUBS 0.007352f
C475 B.n435 VSUBS 0.007352f
C476 B.n436 VSUBS 0.007352f
C477 B.n437 VSUBS 0.007352f
C478 B.n438 VSUBS 0.007352f
C479 B.n439 VSUBS 0.007352f
C480 B.n440 VSUBS 0.007352f
C481 B.n441 VSUBS 0.007352f
C482 B.n442 VSUBS 0.007352f
C483 B.n443 VSUBS 0.007352f
C484 B.n444 VSUBS 0.007352f
C485 B.n445 VSUBS 0.007352f
C486 B.n446 VSUBS 0.007352f
C487 B.n447 VSUBS 0.017116f
C488 B.n448 VSUBS 0.016614f
C489 B.n449 VSUBS 0.016614f
C490 B.n450 VSUBS 0.007352f
C491 B.n451 VSUBS 0.007352f
C492 B.n452 VSUBS 0.007352f
C493 B.n453 VSUBS 0.007352f
C494 B.n454 VSUBS 0.007352f
C495 B.n455 VSUBS 0.007352f
C496 B.n456 VSUBS 0.007352f
C497 B.n457 VSUBS 0.007352f
C498 B.n458 VSUBS 0.007352f
C499 B.n459 VSUBS 0.007352f
C500 B.n460 VSUBS 0.007352f
C501 B.n461 VSUBS 0.007352f
C502 B.n462 VSUBS 0.007352f
C503 B.n463 VSUBS 0.007352f
C504 B.n464 VSUBS 0.007352f
C505 B.n465 VSUBS 0.007352f
C506 B.n466 VSUBS 0.007352f
C507 B.n467 VSUBS 0.007352f
C508 B.n468 VSUBS 0.007352f
C509 B.n469 VSUBS 0.007352f
C510 B.n470 VSUBS 0.007352f
C511 B.n471 VSUBS 0.007352f
C512 B.n472 VSUBS 0.007352f
C513 B.n473 VSUBS 0.007352f
C514 B.n474 VSUBS 0.007352f
C515 B.n475 VSUBS 0.007352f
C516 B.n476 VSUBS 0.007352f
C517 B.n477 VSUBS 0.007352f
C518 B.n478 VSUBS 0.007352f
C519 B.n479 VSUBS 0.007352f
C520 B.n480 VSUBS 0.007352f
C521 B.n481 VSUBS 0.007352f
C522 B.n482 VSUBS 0.007352f
C523 B.n483 VSUBS 0.007352f
C524 B.n484 VSUBS 0.007352f
C525 B.n485 VSUBS 0.007352f
C526 B.n486 VSUBS 0.007352f
C527 B.n487 VSUBS 0.007352f
C528 B.n488 VSUBS 0.007352f
C529 B.n489 VSUBS 0.007352f
C530 B.n490 VSUBS 0.007352f
C531 B.n491 VSUBS 0.007352f
C532 B.n492 VSUBS 0.007352f
C533 B.n493 VSUBS 0.007352f
C534 B.n494 VSUBS 0.007352f
C535 B.n495 VSUBS 0.007352f
C536 B.n496 VSUBS 0.007352f
C537 B.n497 VSUBS 0.007352f
C538 B.n498 VSUBS 0.007352f
C539 B.n499 VSUBS 0.007352f
C540 B.n500 VSUBS 0.007352f
C541 B.n501 VSUBS 0.007352f
C542 B.n502 VSUBS 0.007352f
C543 B.n503 VSUBS 0.007352f
C544 B.n504 VSUBS 0.007352f
C545 B.n505 VSUBS 0.007352f
C546 B.n506 VSUBS 0.007352f
C547 B.n507 VSUBS 0.009593f
C548 B.n508 VSUBS 0.010219f
C549 B.n509 VSUBS 0.020322f
C550 VDD1.t2 VSUBS 0.508711f
C551 VDD1.t5 VSUBS 0.508194f
C552 VDD1.t1 VSUBS 0.064155f
C553 VDD1.t0 VSUBS 0.064155f
C554 VDD1.n0 VSUBS 0.362286f
C555 VDD1.n1 VSUBS 2.43622f
C556 VDD1.t4 VSUBS 0.064155f
C557 VDD1.t3 VSUBS 0.064155f
C558 VDD1.n2 VSUBS 0.359954f
C559 VDD1.n3 VSUBS 2.01608f
C560 VP.n0 VSUBS 0.064369f
C561 VP.t5 VSUBS 1.06173f
C562 VP.n1 VSUBS 0.051344f
C563 VP.n2 VSUBS 0.04882f
C564 VP.t4 VSUBS 1.06173f
C565 VP.n3 VSUBS 0.091445f
C566 VP.n4 VSUBS 0.04882f
C567 VP.n5 VSUBS 0.067967f
C568 VP.n6 VSUBS 0.064369f
C569 VP.t2 VSUBS 1.06173f
C570 VP.n7 VSUBS 0.051344f
C571 VP.n8 VSUBS 0.462702f
C572 VP.t1 VSUBS 1.06173f
C573 VP.t3 VSUBS 1.41808f
C574 VP.n9 VSUBS 0.5432f
C575 VP.n10 VSUBS 0.598469f
C576 VP.n11 VSUBS 0.091445f
C577 VP.n12 VSUBS 0.087046f
C578 VP.n13 VSUBS 0.04882f
C579 VP.n14 VSUBS 0.04882f
C580 VP.n15 VSUBS 0.04882f
C581 VP.n16 VSUBS 0.096213f
C582 VP.n17 VSUBS 0.067967f
C583 VP.n18 VSUBS 0.593243f
C584 VP.n19 VSUBS 2.03494f
C585 VP.t0 VSUBS 1.06173f
C586 VP.n20 VSUBS 0.593243f
C587 VP.n21 VSUBS 2.07706f
C588 VP.n22 VSUBS 0.064369f
C589 VP.n23 VSUBS 0.04882f
C590 VP.n24 VSUBS 0.096213f
C591 VP.n25 VSUBS 0.051344f
C592 VP.n26 VSUBS 0.087046f
C593 VP.n27 VSUBS 0.04882f
C594 VP.n28 VSUBS 0.04882f
C595 VP.n29 VSUBS 0.04882f
C596 VP.n30 VSUBS 0.482724f
C597 VP.n31 VSUBS 0.091445f
C598 VP.n32 VSUBS 0.087046f
C599 VP.n33 VSUBS 0.04882f
C600 VP.n34 VSUBS 0.04882f
C601 VP.n35 VSUBS 0.04882f
C602 VP.n36 VSUBS 0.096213f
C603 VP.n37 VSUBS 0.067967f
C604 VP.n38 VSUBS 0.593243f
C605 VP.n39 VSUBS 0.074489f
C606 VDD2.t0 VSUBS 0.492565f
C607 VDD2.t1 VSUBS 0.062182f
C608 VDD2.t5 VSUBS 0.062182f
C609 VDD2.n0 VSUBS 0.351144f
C610 VDD2.n1 VSUBS 2.26316f
C611 VDD2.t2 VSUBS 0.486569f
C612 VDD2.n2 VSUBS 1.92664f
C613 VDD2.t4 VSUBS 0.062182f
C614 VDD2.t3 VSUBS 0.062182f
C615 VDD2.n3 VSUBS 0.351127f
C616 VTAIL.t10 VSUBS 0.084642f
C617 VTAIL.t8 VSUBS 0.084642f
C618 VTAIL.n0 VSUBS 0.411024f
C619 VTAIL.n1 VSUBS 0.652964f
C620 VTAIL.t0 VSUBS 0.597201f
C621 VTAIL.n2 VSUBS 0.863737f
C622 VTAIL.t1 VSUBS 0.084642f
C623 VTAIL.t4 VSUBS 0.084642f
C624 VTAIL.n3 VSUBS 0.411024f
C625 VTAIL.n4 VSUBS 1.82325f
C626 VTAIL.t9 VSUBS 0.084642f
C627 VTAIL.t7 VSUBS 0.084642f
C628 VTAIL.n5 VSUBS 0.411026f
C629 VTAIL.n6 VSUBS 1.82325f
C630 VTAIL.t6 VSUBS 0.597204f
C631 VTAIL.n7 VSUBS 0.863734f
C632 VTAIL.t2 VSUBS 0.084642f
C633 VTAIL.t5 VSUBS 0.084642f
C634 VTAIL.n8 VSUBS 0.411026f
C635 VTAIL.n9 VSUBS 0.81907f
C636 VTAIL.t3 VSUBS 0.597201f
C637 VTAIL.n10 VSUBS 1.63892f
C638 VTAIL.t11 VSUBS 0.597201f
C639 VTAIL.n11 VSUBS 1.57603f
C640 VN.n0 VSUBS 0.061435f
C641 VN.t0 VSUBS 1.01335f
C642 VN.n1 VSUBS 0.049004f
C643 VN.n2 VSUBS 0.441618f
C644 VN.t4 VSUBS 1.01335f
C645 VN.t5 VSUBS 1.35347f
C646 VN.n3 VSUBS 0.518449f
C647 VN.n4 VSUBS 0.571199f
C648 VN.n5 VSUBS 0.087278f
C649 VN.n6 VSUBS 0.08308f
C650 VN.n7 VSUBS 0.046596f
C651 VN.n8 VSUBS 0.046596f
C652 VN.n9 VSUBS 0.046596f
C653 VN.n10 VSUBS 0.091829f
C654 VN.n11 VSUBS 0.06487f
C655 VN.n12 VSUBS 0.566211f
C656 VN.n13 VSUBS 0.071095f
C657 VN.n14 VSUBS 0.061435f
C658 VN.t3 VSUBS 1.01335f
C659 VN.n15 VSUBS 0.049004f
C660 VN.n16 VSUBS 0.441618f
C661 VN.t1 VSUBS 1.01335f
C662 VN.t2 VSUBS 1.35347f
C663 VN.n17 VSUBS 0.518449f
C664 VN.n18 VSUBS 0.571199f
C665 VN.n19 VSUBS 0.087278f
C666 VN.n20 VSUBS 0.08308f
C667 VN.n21 VSUBS 0.046596f
C668 VN.n22 VSUBS 0.046596f
C669 VN.n23 VSUBS 0.046596f
C670 VN.n24 VSUBS 0.091829f
C671 VN.n25 VSUBS 0.06487f
C672 VN.n26 VSUBS 0.566211f
C673 VN.n27 VSUBS 1.96806f
.ends

