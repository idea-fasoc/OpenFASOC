* NGSPICE file created from diff_pair_sample_1613.ext - technology: sky130A

.subckt diff_pair_sample_1613 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X1 VDD1.t3 VP.t1 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=1.29
X2 VTAIL.t17 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X3 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=1.29
X4 VDD2.t9 VN.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=1.29
X5 VDD1.t0 VP.t3 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=1.29
X6 VDD2.t8 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X7 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=1.29
X8 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=1.29
X9 VDD2.t6 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=1.29
X10 VDD1.t9 VP.t4 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=1.29
X11 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=1.29
X12 VTAIL.t14 VP.t5 VDD1.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X13 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X14 VDD2.t4 VN.t5 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=1.29
X15 VDD2.t3 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X16 VDD1.t4 VP.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X17 VDD1.t5 VP.t7 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=1.29
X18 VTAIL.t11 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X19 VDD1.t8 VP.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X20 VTAIL.t1 VN.t7 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X21 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=1.29
X23 VTAIL.t8 VN.t9 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=1.29
R0 VP.n33 VP.n7 174.089
R1 VP.n56 VP.n55 174.089
R2 VP.n32 VP.n31 174.089
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n12 161.3
R5 VP.n19 VP.n18 161.3
R6 VP.n20 VP.n11 161.3
R7 VP.n22 VP.n21 161.3
R8 VP.n23 VP.n10 161.3
R9 VP.n26 VP.n25 161.3
R10 VP.n27 VP.n9 161.3
R11 VP.n29 VP.n28 161.3
R12 VP.n30 VP.n8 161.3
R13 VP.n54 VP.n0 161.3
R14 VP.n53 VP.n52 161.3
R15 VP.n51 VP.n1 161.3
R16 VP.n50 VP.n49 161.3
R17 VP.n47 VP.n2 161.3
R18 VP.n46 VP.n45 161.3
R19 VP.n44 VP.n3 161.3
R20 VP.n43 VP.n42 161.3
R21 VP.n41 VP.n4 161.3
R22 VP.n40 VP.n39 161.3
R23 VP.n38 VP.n37 161.3
R24 VP.n36 VP.n6 161.3
R25 VP.n35 VP.n34 161.3
R26 VP.n14 VP.t1 80.1495
R27 VP.n14 VP.n13 59.2496
R28 VP.n42 VP.n41 56.5617
R29 VP.n47 VP.n46 56.5617
R30 VP.n23 VP.n22 56.5617
R31 VP.n18 VP.n17 56.5617
R32 VP.n3 VP.t6 51.1896
R33 VP.n7 VP.t7 51.1896
R34 VP.n5 VP.t2 51.1896
R35 VP.n48 VP.t8 51.1896
R36 VP.n55 VP.t3 51.1896
R37 VP.n11 VP.t9 51.1896
R38 VP.n31 VP.t4 51.1896
R39 VP.n24 VP.t0 51.1896
R40 VP.n13 VP.t5 51.1896
R41 VP.n37 VP.n36 47.3584
R42 VP.n53 VP.n1 47.3584
R43 VP.n29 VP.n9 47.3584
R44 VP.n33 VP.n32 38.8793
R45 VP.n36 VP.n35 33.7956
R46 VP.n54 VP.n53 33.7956
R47 VP.n30 VP.n29 33.7956
R48 VP.n15 VP.n14 27.2704
R49 VP.n41 VP.n40 24.5923
R50 VP.n42 VP.n3 24.5923
R51 VP.n46 VP.n3 24.5923
R52 VP.n49 VP.n47 24.5923
R53 VP.n25 VP.n23 24.5923
R54 VP.n18 VP.n11 24.5923
R55 VP.n22 VP.n11 24.5923
R56 VP.n17 VP.n16 24.5923
R57 VP.n37 VP.n5 18.6903
R58 VP.n48 VP.n1 18.6903
R59 VP.n24 VP.n9 18.6903
R60 VP.n35 VP.n7 11.8046
R61 VP.n55 VP.n54 11.8046
R62 VP.n31 VP.n30 11.8046
R63 VP.n40 VP.n5 5.90254
R64 VP.n49 VP.n48 5.90254
R65 VP.n25 VP.n24 5.90254
R66 VP.n16 VP.n13 5.90254
R67 VP.n15 VP.n12 0.189894
R68 VP.n19 VP.n12 0.189894
R69 VP.n20 VP.n19 0.189894
R70 VP.n21 VP.n20 0.189894
R71 VP.n21 VP.n10 0.189894
R72 VP.n26 VP.n10 0.189894
R73 VP.n27 VP.n26 0.189894
R74 VP.n28 VP.n27 0.189894
R75 VP.n28 VP.n8 0.189894
R76 VP.n32 VP.n8 0.189894
R77 VP.n34 VP.n33 0.189894
R78 VP.n34 VP.n6 0.189894
R79 VP.n38 VP.n6 0.189894
R80 VP.n39 VP.n38 0.189894
R81 VP.n39 VP.n4 0.189894
R82 VP.n43 VP.n4 0.189894
R83 VP.n44 VP.n43 0.189894
R84 VP.n45 VP.n44 0.189894
R85 VP.n45 VP.n2 0.189894
R86 VP.n50 VP.n2 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n0 0.189894
R90 VP.n56 VP.n0 0.189894
R91 VP VP.n56 0.0516364
R92 VDD1.n1 VDD1.t3 89.0635
R93 VDD1.n3 VDD1.t5 89.0633
R94 VDD1.n5 VDD1.n4 81.4325
R95 VDD1.n1 VDD1.n0 80.4407
R96 VDD1.n7 VDD1.n6 80.4406
R97 VDD1.n3 VDD1.n2 80.4405
R98 VDD1.n7 VDD1.n5 33.9923
R99 VDD1.n6 VDD1.t6 7.22678
R100 VDD1.n6 VDD1.t9 7.22678
R101 VDD1.n0 VDD1.t2 7.22678
R102 VDD1.n0 VDD1.t8 7.22678
R103 VDD1.n4 VDD1.t1 7.22678
R104 VDD1.n4 VDD1.t0 7.22678
R105 VDD1.n2 VDD1.t7 7.22678
R106 VDD1.n2 VDD1.t4 7.22678
R107 VDD1 VDD1.n7 0.989724
R108 VDD1 VDD1.n1 0.407828
R109 VDD1.n5 VDD1.n3 0.294292
R110 VTAIL.n11 VTAIL.t9 70.9882
R111 VTAIL.n17 VTAIL.t3 70.9879
R112 VTAIL.n2 VTAIL.t16 70.9879
R113 VTAIL.n16 VTAIL.t15 70.9879
R114 VTAIL.n15 VTAIL.n14 63.7619
R115 VTAIL.n13 VTAIL.n12 63.7619
R116 VTAIL.n10 VTAIL.n9 63.7619
R117 VTAIL.n8 VTAIL.n7 63.7619
R118 VTAIL.n19 VTAIL.n18 63.7617
R119 VTAIL.n1 VTAIL.n0 63.7617
R120 VTAIL.n4 VTAIL.n3 63.7617
R121 VTAIL.n6 VTAIL.n5 63.7617
R122 VTAIL.n8 VTAIL.n6 17.5221
R123 VTAIL.n17 VTAIL.n16 16.1255
R124 VTAIL.n18 VTAIL.t2 7.22678
R125 VTAIL.n18 VTAIL.t4 7.22678
R126 VTAIL.n0 VTAIL.t5 7.22678
R127 VTAIL.n0 VTAIL.t8 7.22678
R128 VTAIL.n3 VTAIL.t13 7.22678
R129 VTAIL.n3 VTAIL.t11 7.22678
R130 VTAIL.n5 VTAIL.t12 7.22678
R131 VTAIL.n5 VTAIL.t17 7.22678
R132 VTAIL.n14 VTAIL.t10 7.22678
R133 VTAIL.n14 VTAIL.t19 7.22678
R134 VTAIL.n12 VTAIL.t18 7.22678
R135 VTAIL.n12 VTAIL.t14 7.22678
R136 VTAIL.n9 VTAIL.t6 7.22678
R137 VTAIL.n9 VTAIL.t0 7.22678
R138 VTAIL.n7 VTAIL.t7 7.22678
R139 VTAIL.n7 VTAIL.t1 7.22678
R140 VTAIL.n10 VTAIL.n8 1.39705
R141 VTAIL.n11 VTAIL.n10 1.39705
R142 VTAIL.n15 VTAIL.n13 1.39705
R143 VTAIL.n16 VTAIL.n15 1.39705
R144 VTAIL.n6 VTAIL.n4 1.39705
R145 VTAIL.n4 VTAIL.n2 1.39705
R146 VTAIL.n19 VTAIL.n17 1.39705
R147 VTAIL.n13 VTAIL.n11 1.1686
R148 VTAIL.n2 VTAIL.n1 1.1686
R149 VTAIL VTAIL.n1 1.1061
R150 VTAIL VTAIL.n19 0.291448
R151 B.n493 B.n492 585
R152 B.n164 B.n87 585
R153 B.n163 B.n162 585
R154 B.n161 B.n160 585
R155 B.n159 B.n158 585
R156 B.n157 B.n156 585
R157 B.n155 B.n154 585
R158 B.n153 B.n152 585
R159 B.n151 B.n150 585
R160 B.n149 B.n148 585
R161 B.n147 B.n146 585
R162 B.n145 B.n144 585
R163 B.n143 B.n142 585
R164 B.n141 B.n140 585
R165 B.n139 B.n138 585
R166 B.n137 B.n136 585
R167 B.n135 B.n134 585
R168 B.n133 B.n132 585
R169 B.n131 B.n130 585
R170 B.n129 B.n128 585
R171 B.n127 B.n126 585
R172 B.n125 B.n124 585
R173 B.n123 B.n122 585
R174 B.n121 B.n120 585
R175 B.n119 B.n118 585
R176 B.n117 B.n116 585
R177 B.n115 B.n114 585
R178 B.n113 B.n112 585
R179 B.n111 B.n110 585
R180 B.n109 B.n108 585
R181 B.n107 B.n106 585
R182 B.n105 B.n104 585
R183 B.n103 B.n102 585
R184 B.n101 B.n100 585
R185 B.n99 B.n98 585
R186 B.n97 B.n96 585
R187 B.n95 B.n94 585
R188 B.n67 B.n66 585
R189 B.n491 B.n68 585
R190 B.n496 B.n68 585
R191 B.n490 B.n489 585
R192 B.n489 B.n64 585
R193 B.n488 B.n63 585
R194 B.n502 B.n63 585
R195 B.n487 B.n62 585
R196 B.n503 B.n62 585
R197 B.n486 B.n61 585
R198 B.n504 B.n61 585
R199 B.n485 B.n484 585
R200 B.n484 B.n60 585
R201 B.n483 B.n56 585
R202 B.n510 B.n56 585
R203 B.n482 B.n55 585
R204 B.n511 B.n55 585
R205 B.n481 B.n54 585
R206 B.n512 B.n54 585
R207 B.n480 B.n479 585
R208 B.n479 B.n50 585
R209 B.n478 B.n49 585
R210 B.n518 B.n49 585
R211 B.n477 B.n48 585
R212 B.n519 B.n48 585
R213 B.n476 B.n47 585
R214 B.n520 B.n47 585
R215 B.n475 B.n474 585
R216 B.n474 B.n46 585
R217 B.n473 B.n42 585
R218 B.n526 B.n42 585
R219 B.n472 B.n41 585
R220 B.n527 B.n41 585
R221 B.n471 B.n40 585
R222 B.n528 B.n40 585
R223 B.n470 B.n469 585
R224 B.n469 B.n36 585
R225 B.n468 B.n35 585
R226 B.n534 B.n35 585
R227 B.n467 B.n34 585
R228 B.n535 B.n34 585
R229 B.n466 B.n33 585
R230 B.n536 B.n33 585
R231 B.n465 B.n464 585
R232 B.n464 B.n29 585
R233 B.n463 B.n28 585
R234 B.n542 B.n28 585
R235 B.n462 B.n27 585
R236 B.n543 B.n27 585
R237 B.n461 B.n26 585
R238 B.n544 B.n26 585
R239 B.n460 B.n459 585
R240 B.n459 B.n22 585
R241 B.n458 B.n21 585
R242 B.n550 B.n21 585
R243 B.n457 B.n20 585
R244 B.n551 B.n20 585
R245 B.n456 B.n19 585
R246 B.n552 B.n19 585
R247 B.n455 B.n454 585
R248 B.n454 B.n15 585
R249 B.n453 B.n14 585
R250 B.n558 B.n14 585
R251 B.n452 B.n13 585
R252 B.n559 B.n13 585
R253 B.n451 B.n12 585
R254 B.n560 B.n12 585
R255 B.n450 B.n449 585
R256 B.n449 B.n448 585
R257 B.n447 B.n446 585
R258 B.n447 B.n8 585
R259 B.n445 B.n7 585
R260 B.n567 B.n7 585
R261 B.n444 B.n6 585
R262 B.n568 B.n6 585
R263 B.n443 B.n5 585
R264 B.n569 B.n5 585
R265 B.n442 B.n441 585
R266 B.n441 B.n4 585
R267 B.n440 B.n165 585
R268 B.n440 B.n439 585
R269 B.n430 B.n166 585
R270 B.n167 B.n166 585
R271 B.n432 B.n431 585
R272 B.n433 B.n432 585
R273 B.n429 B.n172 585
R274 B.n172 B.n171 585
R275 B.n428 B.n427 585
R276 B.n427 B.n426 585
R277 B.n174 B.n173 585
R278 B.n175 B.n174 585
R279 B.n419 B.n418 585
R280 B.n420 B.n419 585
R281 B.n417 B.n179 585
R282 B.n183 B.n179 585
R283 B.n416 B.n415 585
R284 B.n415 B.n414 585
R285 B.n181 B.n180 585
R286 B.n182 B.n181 585
R287 B.n407 B.n406 585
R288 B.n408 B.n407 585
R289 B.n405 B.n188 585
R290 B.n188 B.n187 585
R291 B.n404 B.n403 585
R292 B.n403 B.n402 585
R293 B.n190 B.n189 585
R294 B.n191 B.n190 585
R295 B.n395 B.n394 585
R296 B.n396 B.n395 585
R297 B.n393 B.n196 585
R298 B.n196 B.n195 585
R299 B.n392 B.n391 585
R300 B.n391 B.n390 585
R301 B.n198 B.n197 585
R302 B.n199 B.n198 585
R303 B.n383 B.n382 585
R304 B.n384 B.n383 585
R305 B.n381 B.n204 585
R306 B.n204 B.n203 585
R307 B.n380 B.n379 585
R308 B.n379 B.n378 585
R309 B.n206 B.n205 585
R310 B.n371 B.n206 585
R311 B.n370 B.n369 585
R312 B.n372 B.n370 585
R313 B.n368 B.n211 585
R314 B.n211 B.n210 585
R315 B.n367 B.n366 585
R316 B.n366 B.n365 585
R317 B.n213 B.n212 585
R318 B.n214 B.n213 585
R319 B.n358 B.n357 585
R320 B.n359 B.n358 585
R321 B.n356 B.n219 585
R322 B.n219 B.n218 585
R323 B.n355 B.n354 585
R324 B.n354 B.n353 585
R325 B.n221 B.n220 585
R326 B.n346 B.n221 585
R327 B.n345 B.n344 585
R328 B.n347 B.n345 585
R329 B.n343 B.n226 585
R330 B.n226 B.n225 585
R331 B.n342 B.n341 585
R332 B.n341 B.n340 585
R333 B.n228 B.n227 585
R334 B.n229 B.n228 585
R335 B.n333 B.n332 585
R336 B.n334 B.n333 585
R337 B.n232 B.n231 585
R338 B.n257 B.n255 585
R339 B.n258 B.n254 585
R340 B.n258 B.n233 585
R341 B.n261 B.n260 585
R342 B.n262 B.n253 585
R343 B.n264 B.n263 585
R344 B.n266 B.n252 585
R345 B.n269 B.n268 585
R346 B.n270 B.n251 585
R347 B.n272 B.n271 585
R348 B.n274 B.n250 585
R349 B.n277 B.n276 585
R350 B.n278 B.n249 585
R351 B.n283 B.n282 585
R352 B.n285 B.n248 585
R353 B.n288 B.n287 585
R354 B.n289 B.n247 585
R355 B.n291 B.n290 585
R356 B.n293 B.n246 585
R357 B.n296 B.n295 585
R358 B.n297 B.n245 585
R359 B.n299 B.n298 585
R360 B.n301 B.n244 585
R361 B.n304 B.n303 585
R362 B.n306 B.n241 585
R363 B.n308 B.n307 585
R364 B.n310 B.n240 585
R365 B.n313 B.n312 585
R366 B.n314 B.n239 585
R367 B.n316 B.n315 585
R368 B.n318 B.n238 585
R369 B.n321 B.n320 585
R370 B.n322 B.n237 585
R371 B.n324 B.n323 585
R372 B.n326 B.n236 585
R373 B.n327 B.n235 585
R374 B.n330 B.n329 585
R375 B.n331 B.n234 585
R376 B.n234 B.n233 585
R377 B.n336 B.n335 585
R378 B.n335 B.n334 585
R379 B.n337 B.n230 585
R380 B.n230 B.n229 585
R381 B.n339 B.n338 585
R382 B.n340 B.n339 585
R383 B.n224 B.n223 585
R384 B.n225 B.n224 585
R385 B.n349 B.n348 585
R386 B.n348 B.n347 585
R387 B.n350 B.n222 585
R388 B.n346 B.n222 585
R389 B.n352 B.n351 585
R390 B.n353 B.n352 585
R391 B.n217 B.n216 585
R392 B.n218 B.n217 585
R393 B.n361 B.n360 585
R394 B.n360 B.n359 585
R395 B.n362 B.n215 585
R396 B.n215 B.n214 585
R397 B.n364 B.n363 585
R398 B.n365 B.n364 585
R399 B.n209 B.n208 585
R400 B.n210 B.n209 585
R401 B.n374 B.n373 585
R402 B.n373 B.n372 585
R403 B.n375 B.n207 585
R404 B.n371 B.n207 585
R405 B.n377 B.n376 585
R406 B.n378 B.n377 585
R407 B.n202 B.n201 585
R408 B.n203 B.n202 585
R409 B.n386 B.n385 585
R410 B.n385 B.n384 585
R411 B.n387 B.n200 585
R412 B.n200 B.n199 585
R413 B.n389 B.n388 585
R414 B.n390 B.n389 585
R415 B.n194 B.n193 585
R416 B.n195 B.n194 585
R417 B.n398 B.n397 585
R418 B.n397 B.n396 585
R419 B.n399 B.n192 585
R420 B.n192 B.n191 585
R421 B.n401 B.n400 585
R422 B.n402 B.n401 585
R423 B.n186 B.n185 585
R424 B.n187 B.n186 585
R425 B.n410 B.n409 585
R426 B.n409 B.n408 585
R427 B.n411 B.n184 585
R428 B.n184 B.n182 585
R429 B.n413 B.n412 585
R430 B.n414 B.n413 585
R431 B.n178 B.n177 585
R432 B.n183 B.n178 585
R433 B.n422 B.n421 585
R434 B.n421 B.n420 585
R435 B.n423 B.n176 585
R436 B.n176 B.n175 585
R437 B.n425 B.n424 585
R438 B.n426 B.n425 585
R439 B.n170 B.n169 585
R440 B.n171 B.n170 585
R441 B.n435 B.n434 585
R442 B.n434 B.n433 585
R443 B.n436 B.n168 585
R444 B.n168 B.n167 585
R445 B.n438 B.n437 585
R446 B.n439 B.n438 585
R447 B.n3 B.n0 585
R448 B.n4 B.n3 585
R449 B.n566 B.n1 585
R450 B.n567 B.n566 585
R451 B.n565 B.n564 585
R452 B.n565 B.n8 585
R453 B.n563 B.n9 585
R454 B.n448 B.n9 585
R455 B.n562 B.n561 585
R456 B.n561 B.n560 585
R457 B.n11 B.n10 585
R458 B.n559 B.n11 585
R459 B.n557 B.n556 585
R460 B.n558 B.n557 585
R461 B.n555 B.n16 585
R462 B.n16 B.n15 585
R463 B.n554 B.n553 585
R464 B.n553 B.n552 585
R465 B.n18 B.n17 585
R466 B.n551 B.n18 585
R467 B.n549 B.n548 585
R468 B.n550 B.n549 585
R469 B.n547 B.n23 585
R470 B.n23 B.n22 585
R471 B.n546 B.n545 585
R472 B.n545 B.n544 585
R473 B.n25 B.n24 585
R474 B.n543 B.n25 585
R475 B.n541 B.n540 585
R476 B.n542 B.n541 585
R477 B.n539 B.n30 585
R478 B.n30 B.n29 585
R479 B.n538 B.n537 585
R480 B.n537 B.n536 585
R481 B.n32 B.n31 585
R482 B.n535 B.n32 585
R483 B.n533 B.n532 585
R484 B.n534 B.n533 585
R485 B.n531 B.n37 585
R486 B.n37 B.n36 585
R487 B.n530 B.n529 585
R488 B.n529 B.n528 585
R489 B.n39 B.n38 585
R490 B.n527 B.n39 585
R491 B.n525 B.n524 585
R492 B.n526 B.n525 585
R493 B.n523 B.n43 585
R494 B.n46 B.n43 585
R495 B.n522 B.n521 585
R496 B.n521 B.n520 585
R497 B.n45 B.n44 585
R498 B.n519 B.n45 585
R499 B.n517 B.n516 585
R500 B.n518 B.n517 585
R501 B.n515 B.n51 585
R502 B.n51 B.n50 585
R503 B.n514 B.n513 585
R504 B.n513 B.n512 585
R505 B.n53 B.n52 585
R506 B.n511 B.n53 585
R507 B.n509 B.n508 585
R508 B.n510 B.n509 585
R509 B.n507 B.n57 585
R510 B.n60 B.n57 585
R511 B.n506 B.n505 585
R512 B.n505 B.n504 585
R513 B.n59 B.n58 585
R514 B.n503 B.n59 585
R515 B.n501 B.n500 585
R516 B.n502 B.n501 585
R517 B.n499 B.n65 585
R518 B.n65 B.n64 585
R519 B.n498 B.n497 585
R520 B.n497 B.n496 585
R521 B.n570 B.n569 585
R522 B.n568 B.n2 585
R523 B.n497 B.n67 559.769
R524 B.n493 B.n68 559.769
R525 B.n333 B.n234 559.769
R526 B.n335 B.n232 559.769
R527 B.n495 B.n494 256.663
R528 B.n495 B.n86 256.663
R529 B.n495 B.n85 256.663
R530 B.n495 B.n84 256.663
R531 B.n495 B.n83 256.663
R532 B.n495 B.n82 256.663
R533 B.n495 B.n81 256.663
R534 B.n495 B.n80 256.663
R535 B.n495 B.n79 256.663
R536 B.n495 B.n78 256.663
R537 B.n495 B.n77 256.663
R538 B.n495 B.n76 256.663
R539 B.n495 B.n75 256.663
R540 B.n495 B.n74 256.663
R541 B.n495 B.n73 256.663
R542 B.n495 B.n72 256.663
R543 B.n495 B.n71 256.663
R544 B.n495 B.n70 256.663
R545 B.n495 B.n69 256.663
R546 B.n256 B.n233 256.663
R547 B.n259 B.n233 256.663
R548 B.n265 B.n233 256.663
R549 B.n267 B.n233 256.663
R550 B.n273 B.n233 256.663
R551 B.n275 B.n233 256.663
R552 B.n284 B.n233 256.663
R553 B.n286 B.n233 256.663
R554 B.n292 B.n233 256.663
R555 B.n294 B.n233 256.663
R556 B.n300 B.n233 256.663
R557 B.n302 B.n233 256.663
R558 B.n309 B.n233 256.663
R559 B.n311 B.n233 256.663
R560 B.n317 B.n233 256.663
R561 B.n319 B.n233 256.663
R562 B.n325 B.n233 256.663
R563 B.n328 B.n233 256.663
R564 B.n572 B.n571 256.663
R565 B.n91 B.t18 255.751
R566 B.n88 B.t14 255.751
R567 B.n242 B.t21 255.751
R568 B.n279 B.t10 255.751
R569 B.n334 B.n233 188.023
R570 B.n496 B.n495 188.023
R571 B.n96 B.n95 163.367
R572 B.n100 B.n99 163.367
R573 B.n104 B.n103 163.367
R574 B.n108 B.n107 163.367
R575 B.n112 B.n111 163.367
R576 B.n116 B.n115 163.367
R577 B.n120 B.n119 163.367
R578 B.n124 B.n123 163.367
R579 B.n128 B.n127 163.367
R580 B.n132 B.n131 163.367
R581 B.n136 B.n135 163.367
R582 B.n140 B.n139 163.367
R583 B.n144 B.n143 163.367
R584 B.n148 B.n147 163.367
R585 B.n152 B.n151 163.367
R586 B.n156 B.n155 163.367
R587 B.n160 B.n159 163.367
R588 B.n162 B.n87 163.367
R589 B.n333 B.n228 163.367
R590 B.n341 B.n228 163.367
R591 B.n341 B.n226 163.367
R592 B.n345 B.n226 163.367
R593 B.n345 B.n221 163.367
R594 B.n354 B.n221 163.367
R595 B.n354 B.n219 163.367
R596 B.n358 B.n219 163.367
R597 B.n358 B.n213 163.367
R598 B.n366 B.n213 163.367
R599 B.n366 B.n211 163.367
R600 B.n370 B.n211 163.367
R601 B.n370 B.n206 163.367
R602 B.n379 B.n206 163.367
R603 B.n379 B.n204 163.367
R604 B.n383 B.n204 163.367
R605 B.n383 B.n198 163.367
R606 B.n391 B.n198 163.367
R607 B.n391 B.n196 163.367
R608 B.n395 B.n196 163.367
R609 B.n395 B.n190 163.367
R610 B.n403 B.n190 163.367
R611 B.n403 B.n188 163.367
R612 B.n407 B.n188 163.367
R613 B.n407 B.n181 163.367
R614 B.n415 B.n181 163.367
R615 B.n415 B.n179 163.367
R616 B.n419 B.n179 163.367
R617 B.n419 B.n174 163.367
R618 B.n427 B.n174 163.367
R619 B.n427 B.n172 163.367
R620 B.n432 B.n172 163.367
R621 B.n432 B.n166 163.367
R622 B.n440 B.n166 163.367
R623 B.n441 B.n440 163.367
R624 B.n441 B.n5 163.367
R625 B.n6 B.n5 163.367
R626 B.n7 B.n6 163.367
R627 B.n447 B.n7 163.367
R628 B.n449 B.n447 163.367
R629 B.n449 B.n12 163.367
R630 B.n13 B.n12 163.367
R631 B.n14 B.n13 163.367
R632 B.n454 B.n14 163.367
R633 B.n454 B.n19 163.367
R634 B.n20 B.n19 163.367
R635 B.n21 B.n20 163.367
R636 B.n459 B.n21 163.367
R637 B.n459 B.n26 163.367
R638 B.n27 B.n26 163.367
R639 B.n28 B.n27 163.367
R640 B.n464 B.n28 163.367
R641 B.n464 B.n33 163.367
R642 B.n34 B.n33 163.367
R643 B.n35 B.n34 163.367
R644 B.n469 B.n35 163.367
R645 B.n469 B.n40 163.367
R646 B.n41 B.n40 163.367
R647 B.n42 B.n41 163.367
R648 B.n474 B.n42 163.367
R649 B.n474 B.n47 163.367
R650 B.n48 B.n47 163.367
R651 B.n49 B.n48 163.367
R652 B.n479 B.n49 163.367
R653 B.n479 B.n54 163.367
R654 B.n55 B.n54 163.367
R655 B.n56 B.n55 163.367
R656 B.n484 B.n56 163.367
R657 B.n484 B.n61 163.367
R658 B.n62 B.n61 163.367
R659 B.n63 B.n62 163.367
R660 B.n489 B.n63 163.367
R661 B.n489 B.n68 163.367
R662 B.n258 B.n257 163.367
R663 B.n260 B.n258 163.367
R664 B.n264 B.n253 163.367
R665 B.n268 B.n266 163.367
R666 B.n272 B.n251 163.367
R667 B.n276 B.n274 163.367
R668 B.n283 B.n249 163.367
R669 B.n287 B.n285 163.367
R670 B.n291 B.n247 163.367
R671 B.n295 B.n293 163.367
R672 B.n299 B.n245 163.367
R673 B.n303 B.n301 163.367
R674 B.n308 B.n241 163.367
R675 B.n312 B.n310 163.367
R676 B.n316 B.n239 163.367
R677 B.n320 B.n318 163.367
R678 B.n324 B.n237 163.367
R679 B.n327 B.n326 163.367
R680 B.n329 B.n234 163.367
R681 B.n335 B.n230 163.367
R682 B.n339 B.n230 163.367
R683 B.n339 B.n224 163.367
R684 B.n348 B.n224 163.367
R685 B.n348 B.n222 163.367
R686 B.n352 B.n222 163.367
R687 B.n352 B.n217 163.367
R688 B.n360 B.n217 163.367
R689 B.n360 B.n215 163.367
R690 B.n364 B.n215 163.367
R691 B.n364 B.n209 163.367
R692 B.n373 B.n209 163.367
R693 B.n373 B.n207 163.367
R694 B.n377 B.n207 163.367
R695 B.n377 B.n202 163.367
R696 B.n385 B.n202 163.367
R697 B.n385 B.n200 163.367
R698 B.n389 B.n200 163.367
R699 B.n389 B.n194 163.367
R700 B.n397 B.n194 163.367
R701 B.n397 B.n192 163.367
R702 B.n401 B.n192 163.367
R703 B.n401 B.n186 163.367
R704 B.n409 B.n186 163.367
R705 B.n409 B.n184 163.367
R706 B.n413 B.n184 163.367
R707 B.n413 B.n178 163.367
R708 B.n421 B.n178 163.367
R709 B.n421 B.n176 163.367
R710 B.n425 B.n176 163.367
R711 B.n425 B.n170 163.367
R712 B.n434 B.n170 163.367
R713 B.n434 B.n168 163.367
R714 B.n438 B.n168 163.367
R715 B.n438 B.n3 163.367
R716 B.n570 B.n3 163.367
R717 B.n566 B.n2 163.367
R718 B.n566 B.n565 163.367
R719 B.n565 B.n9 163.367
R720 B.n561 B.n9 163.367
R721 B.n561 B.n11 163.367
R722 B.n557 B.n11 163.367
R723 B.n557 B.n16 163.367
R724 B.n553 B.n16 163.367
R725 B.n553 B.n18 163.367
R726 B.n549 B.n18 163.367
R727 B.n549 B.n23 163.367
R728 B.n545 B.n23 163.367
R729 B.n545 B.n25 163.367
R730 B.n541 B.n25 163.367
R731 B.n541 B.n30 163.367
R732 B.n537 B.n30 163.367
R733 B.n537 B.n32 163.367
R734 B.n533 B.n32 163.367
R735 B.n533 B.n37 163.367
R736 B.n529 B.n37 163.367
R737 B.n529 B.n39 163.367
R738 B.n525 B.n39 163.367
R739 B.n525 B.n43 163.367
R740 B.n521 B.n43 163.367
R741 B.n521 B.n45 163.367
R742 B.n517 B.n45 163.367
R743 B.n517 B.n51 163.367
R744 B.n513 B.n51 163.367
R745 B.n513 B.n53 163.367
R746 B.n509 B.n53 163.367
R747 B.n509 B.n57 163.367
R748 B.n505 B.n57 163.367
R749 B.n505 B.n59 163.367
R750 B.n501 B.n59 163.367
R751 B.n501 B.n65 163.367
R752 B.n497 B.n65 163.367
R753 B.n88 B.t16 107.617
R754 B.n242 B.t23 107.617
R755 B.n91 B.t19 107.615
R756 B.n279 B.t13 107.615
R757 B.n334 B.n229 93.3255
R758 B.n340 B.n229 93.3255
R759 B.n340 B.n225 93.3255
R760 B.n347 B.n225 93.3255
R761 B.n347 B.n346 93.3255
R762 B.n353 B.n218 93.3255
R763 B.n359 B.n218 93.3255
R764 B.n359 B.n214 93.3255
R765 B.n365 B.n214 93.3255
R766 B.n365 B.n210 93.3255
R767 B.n372 B.n210 93.3255
R768 B.n372 B.n371 93.3255
R769 B.n378 B.n203 93.3255
R770 B.n384 B.n203 93.3255
R771 B.n384 B.n199 93.3255
R772 B.n390 B.n199 93.3255
R773 B.n396 B.n195 93.3255
R774 B.n396 B.n191 93.3255
R775 B.n402 B.n191 93.3255
R776 B.n408 B.n187 93.3255
R777 B.n408 B.n182 93.3255
R778 B.n414 B.n182 93.3255
R779 B.n414 B.n183 93.3255
R780 B.n420 B.n175 93.3255
R781 B.n426 B.n175 93.3255
R782 B.n426 B.n171 93.3255
R783 B.n433 B.n171 93.3255
R784 B.n439 B.n167 93.3255
R785 B.n439 B.n4 93.3255
R786 B.n569 B.n4 93.3255
R787 B.n569 B.n568 93.3255
R788 B.n568 B.n567 93.3255
R789 B.n567 B.n8 93.3255
R790 B.n448 B.n8 93.3255
R791 B.n560 B.n559 93.3255
R792 B.n559 B.n558 93.3255
R793 B.n558 B.n15 93.3255
R794 B.n552 B.n15 93.3255
R795 B.n551 B.n550 93.3255
R796 B.n550 B.n22 93.3255
R797 B.n544 B.n22 93.3255
R798 B.n544 B.n543 93.3255
R799 B.n542 B.n29 93.3255
R800 B.n536 B.n29 93.3255
R801 B.n536 B.n535 93.3255
R802 B.n534 B.n36 93.3255
R803 B.n528 B.n36 93.3255
R804 B.n528 B.n527 93.3255
R805 B.n527 B.n526 93.3255
R806 B.n520 B.n46 93.3255
R807 B.n520 B.n519 93.3255
R808 B.n519 B.n518 93.3255
R809 B.n518 B.n50 93.3255
R810 B.n512 B.n50 93.3255
R811 B.n512 B.n511 93.3255
R812 B.n511 B.n510 93.3255
R813 B.n504 B.n60 93.3255
R814 B.n504 B.n503 93.3255
R815 B.n503 B.n502 93.3255
R816 B.n502 B.n64 93.3255
R817 B.n496 B.n64 93.3255
R818 B.n402 B.t6 91.9531
R819 B.t2 B.n542 91.9531
R820 B.n89 B.t17 76.1987
R821 B.n243 B.t22 76.1987
R822 B.n92 B.t20 76.1968
R823 B.n280 B.t12 76.1968
R824 B.t1 B.n195 72.7391
R825 B.n535 B.t4 72.7391
R826 B.n69 B.n67 71.676
R827 B.n96 B.n70 71.676
R828 B.n100 B.n71 71.676
R829 B.n104 B.n72 71.676
R830 B.n108 B.n73 71.676
R831 B.n112 B.n74 71.676
R832 B.n116 B.n75 71.676
R833 B.n120 B.n76 71.676
R834 B.n124 B.n77 71.676
R835 B.n128 B.n78 71.676
R836 B.n132 B.n79 71.676
R837 B.n136 B.n80 71.676
R838 B.n140 B.n81 71.676
R839 B.n144 B.n82 71.676
R840 B.n148 B.n83 71.676
R841 B.n152 B.n84 71.676
R842 B.n156 B.n85 71.676
R843 B.n160 B.n86 71.676
R844 B.n494 B.n87 71.676
R845 B.n494 B.n493 71.676
R846 B.n162 B.n86 71.676
R847 B.n159 B.n85 71.676
R848 B.n155 B.n84 71.676
R849 B.n151 B.n83 71.676
R850 B.n147 B.n82 71.676
R851 B.n143 B.n81 71.676
R852 B.n139 B.n80 71.676
R853 B.n135 B.n79 71.676
R854 B.n131 B.n78 71.676
R855 B.n127 B.n77 71.676
R856 B.n123 B.n76 71.676
R857 B.n119 B.n75 71.676
R858 B.n115 B.n74 71.676
R859 B.n111 B.n73 71.676
R860 B.n107 B.n72 71.676
R861 B.n103 B.n71 71.676
R862 B.n99 B.n70 71.676
R863 B.n95 B.n69 71.676
R864 B.n256 B.n232 71.676
R865 B.n260 B.n259 71.676
R866 B.n265 B.n264 71.676
R867 B.n268 B.n267 71.676
R868 B.n273 B.n272 71.676
R869 B.n276 B.n275 71.676
R870 B.n284 B.n283 71.676
R871 B.n287 B.n286 71.676
R872 B.n292 B.n291 71.676
R873 B.n295 B.n294 71.676
R874 B.n300 B.n299 71.676
R875 B.n303 B.n302 71.676
R876 B.n309 B.n308 71.676
R877 B.n312 B.n311 71.676
R878 B.n317 B.n316 71.676
R879 B.n320 B.n319 71.676
R880 B.n325 B.n324 71.676
R881 B.n328 B.n327 71.676
R882 B.n257 B.n256 71.676
R883 B.n259 B.n253 71.676
R884 B.n266 B.n265 71.676
R885 B.n267 B.n251 71.676
R886 B.n274 B.n273 71.676
R887 B.n275 B.n249 71.676
R888 B.n285 B.n284 71.676
R889 B.n286 B.n247 71.676
R890 B.n293 B.n292 71.676
R891 B.n294 B.n245 71.676
R892 B.n301 B.n300 71.676
R893 B.n302 B.n241 71.676
R894 B.n310 B.n309 71.676
R895 B.n311 B.n239 71.676
R896 B.n318 B.n317 71.676
R897 B.n319 B.n237 71.676
R898 B.n326 B.n325 71.676
R899 B.n329 B.n328 71.676
R900 B.n571 B.n570 71.676
R901 B.n571 B.n2 71.676
R902 B.n183 B.t0 69.9943
R903 B.t8 B.n551 69.9943
R904 B.n93 B.n92 59.5399
R905 B.n90 B.n89 59.5399
R906 B.n305 B.n243 59.5399
R907 B.n281 B.n280 59.5399
R908 B.n378 B.t7 50.7803
R909 B.n526 B.t3 50.7803
R910 B.n353 B.t11 48.0354
R911 B.n433 B.t9 48.0354
R912 B.n560 B.t5 48.0354
R913 B.n510 B.t15 48.0354
R914 B.n346 B.t11 45.2906
R915 B.t9 B.n167 45.2906
R916 B.n448 B.t5 45.2906
R917 B.n60 B.t15 45.2906
R918 B.n371 B.t7 42.5457
R919 B.n46 B.t3 42.5457
R920 B.n336 B.n231 36.3712
R921 B.n332 B.n331 36.3712
R922 B.n492 B.n491 36.3712
R923 B.n498 B.n66 36.3712
R924 B.n92 B.n91 31.4187
R925 B.n89 B.n88 31.4187
R926 B.n243 B.n242 31.4187
R927 B.n280 B.n279 31.4187
R928 B.n420 B.t0 23.3318
R929 B.n552 B.t8 23.3318
R930 B.n390 B.t1 20.5869
R931 B.t4 B.n534 20.5869
R932 B B.n572 18.0485
R933 B.n337 B.n336 10.6151
R934 B.n338 B.n337 10.6151
R935 B.n338 B.n223 10.6151
R936 B.n349 B.n223 10.6151
R937 B.n350 B.n349 10.6151
R938 B.n351 B.n350 10.6151
R939 B.n351 B.n216 10.6151
R940 B.n361 B.n216 10.6151
R941 B.n362 B.n361 10.6151
R942 B.n363 B.n362 10.6151
R943 B.n363 B.n208 10.6151
R944 B.n374 B.n208 10.6151
R945 B.n375 B.n374 10.6151
R946 B.n376 B.n375 10.6151
R947 B.n376 B.n201 10.6151
R948 B.n386 B.n201 10.6151
R949 B.n387 B.n386 10.6151
R950 B.n388 B.n387 10.6151
R951 B.n388 B.n193 10.6151
R952 B.n398 B.n193 10.6151
R953 B.n399 B.n398 10.6151
R954 B.n400 B.n399 10.6151
R955 B.n400 B.n185 10.6151
R956 B.n410 B.n185 10.6151
R957 B.n411 B.n410 10.6151
R958 B.n412 B.n411 10.6151
R959 B.n412 B.n177 10.6151
R960 B.n422 B.n177 10.6151
R961 B.n423 B.n422 10.6151
R962 B.n424 B.n423 10.6151
R963 B.n424 B.n169 10.6151
R964 B.n435 B.n169 10.6151
R965 B.n436 B.n435 10.6151
R966 B.n437 B.n436 10.6151
R967 B.n437 B.n0 10.6151
R968 B.n255 B.n231 10.6151
R969 B.n255 B.n254 10.6151
R970 B.n261 B.n254 10.6151
R971 B.n262 B.n261 10.6151
R972 B.n263 B.n262 10.6151
R973 B.n263 B.n252 10.6151
R974 B.n269 B.n252 10.6151
R975 B.n270 B.n269 10.6151
R976 B.n271 B.n270 10.6151
R977 B.n271 B.n250 10.6151
R978 B.n277 B.n250 10.6151
R979 B.n278 B.n277 10.6151
R980 B.n282 B.n278 10.6151
R981 B.n288 B.n248 10.6151
R982 B.n289 B.n288 10.6151
R983 B.n290 B.n289 10.6151
R984 B.n290 B.n246 10.6151
R985 B.n296 B.n246 10.6151
R986 B.n297 B.n296 10.6151
R987 B.n298 B.n297 10.6151
R988 B.n298 B.n244 10.6151
R989 B.n304 B.n244 10.6151
R990 B.n307 B.n306 10.6151
R991 B.n307 B.n240 10.6151
R992 B.n313 B.n240 10.6151
R993 B.n314 B.n313 10.6151
R994 B.n315 B.n314 10.6151
R995 B.n315 B.n238 10.6151
R996 B.n321 B.n238 10.6151
R997 B.n322 B.n321 10.6151
R998 B.n323 B.n322 10.6151
R999 B.n323 B.n236 10.6151
R1000 B.n236 B.n235 10.6151
R1001 B.n330 B.n235 10.6151
R1002 B.n331 B.n330 10.6151
R1003 B.n332 B.n227 10.6151
R1004 B.n342 B.n227 10.6151
R1005 B.n343 B.n342 10.6151
R1006 B.n344 B.n343 10.6151
R1007 B.n344 B.n220 10.6151
R1008 B.n355 B.n220 10.6151
R1009 B.n356 B.n355 10.6151
R1010 B.n357 B.n356 10.6151
R1011 B.n357 B.n212 10.6151
R1012 B.n367 B.n212 10.6151
R1013 B.n368 B.n367 10.6151
R1014 B.n369 B.n368 10.6151
R1015 B.n369 B.n205 10.6151
R1016 B.n380 B.n205 10.6151
R1017 B.n381 B.n380 10.6151
R1018 B.n382 B.n381 10.6151
R1019 B.n382 B.n197 10.6151
R1020 B.n392 B.n197 10.6151
R1021 B.n393 B.n392 10.6151
R1022 B.n394 B.n393 10.6151
R1023 B.n394 B.n189 10.6151
R1024 B.n404 B.n189 10.6151
R1025 B.n405 B.n404 10.6151
R1026 B.n406 B.n405 10.6151
R1027 B.n406 B.n180 10.6151
R1028 B.n416 B.n180 10.6151
R1029 B.n417 B.n416 10.6151
R1030 B.n418 B.n417 10.6151
R1031 B.n418 B.n173 10.6151
R1032 B.n428 B.n173 10.6151
R1033 B.n429 B.n428 10.6151
R1034 B.n431 B.n429 10.6151
R1035 B.n431 B.n430 10.6151
R1036 B.n430 B.n165 10.6151
R1037 B.n442 B.n165 10.6151
R1038 B.n443 B.n442 10.6151
R1039 B.n444 B.n443 10.6151
R1040 B.n445 B.n444 10.6151
R1041 B.n446 B.n445 10.6151
R1042 B.n450 B.n446 10.6151
R1043 B.n451 B.n450 10.6151
R1044 B.n452 B.n451 10.6151
R1045 B.n453 B.n452 10.6151
R1046 B.n455 B.n453 10.6151
R1047 B.n456 B.n455 10.6151
R1048 B.n457 B.n456 10.6151
R1049 B.n458 B.n457 10.6151
R1050 B.n460 B.n458 10.6151
R1051 B.n461 B.n460 10.6151
R1052 B.n462 B.n461 10.6151
R1053 B.n463 B.n462 10.6151
R1054 B.n465 B.n463 10.6151
R1055 B.n466 B.n465 10.6151
R1056 B.n467 B.n466 10.6151
R1057 B.n468 B.n467 10.6151
R1058 B.n470 B.n468 10.6151
R1059 B.n471 B.n470 10.6151
R1060 B.n472 B.n471 10.6151
R1061 B.n473 B.n472 10.6151
R1062 B.n475 B.n473 10.6151
R1063 B.n476 B.n475 10.6151
R1064 B.n477 B.n476 10.6151
R1065 B.n478 B.n477 10.6151
R1066 B.n480 B.n478 10.6151
R1067 B.n481 B.n480 10.6151
R1068 B.n482 B.n481 10.6151
R1069 B.n483 B.n482 10.6151
R1070 B.n485 B.n483 10.6151
R1071 B.n486 B.n485 10.6151
R1072 B.n487 B.n486 10.6151
R1073 B.n488 B.n487 10.6151
R1074 B.n490 B.n488 10.6151
R1075 B.n491 B.n490 10.6151
R1076 B.n564 B.n1 10.6151
R1077 B.n564 B.n563 10.6151
R1078 B.n563 B.n562 10.6151
R1079 B.n562 B.n10 10.6151
R1080 B.n556 B.n10 10.6151
R1081 B.n556 B.n555 10.6151
R1082 B.n555 B.n554 10.6151
R1083 B.n554 B.n17 10.6151
R1084 B.n548 B.n17 10.6151
R1085 B.n548 B.n547 10.6151
R1086 B.n547 B.n546 10.6151
R1087 B.n546 B.n24 10.6151
R1088 B.n540 B.n24 10.6151
R1089 B.n540 B.n539 10.6151
R1090 B.n539 B.n538 10.6151
R1091 B.n538 B.n31 10.6151
R1092 B.n532 B.n31 10.6151
R1093 B.n532 B.n531 10.6151
R1094 B.n531 B.n530 10.6151
R1095 B.n530 B.n38 10.6151
R1096 B.n524 B.n38 10.6151
R1097 B.n524 B.n523 10.6151
R1098 B.n523 B.n522 10.6151
R1099 B.n522 B.n44 10.6151
R1100 B.n516 B.n44 10.6151
R1101 B.n516 B.n515 10.6151
R1102 B.n515 B.n514 10.6151
R1103 B.n514 B.n52 10.6151
R1104 B.n508 B.n52 10.6151
R1105 B.n508 B.n507 10.6151
R1106 B.n507 B.n506 10.6151
R1107 B.n506 B.n58 10.6151
R1108 B.n500 B.n58 10.6151
R1109 B.n500 B.n499 10.6151
R1110 B.n499 B.n498 10.6151
R1111 B.n94 B.n66 10.6151
R1112 B.n97 B.n94 10.6151
R1113 B.n98 B.n97 10.6151
R1114 B.n101 B.n98 10.6151
R1115 B.n102 B.n101 10.6151
R1116 B.n105 B.n102 10.6151
R1117 B.n106 B.n105 10.6151
R1118 B.n109 B.n106 10.6151
R1119 B.n110 B.n109 10.6151
R1120 B.n113 B.n110 10.6151
R1121 B.n114 B.n113 10.6151
R1122 B.n117 B.n114 10.6151
R1123 B.n118 B.n117 10.6151
R1124 B.n122 B.n121 10.6151
R1125 B.n125 B.n122 10.6151
R1126 B.n126 B.n125 10.6151
R1127 B.n129 B.n126 10.6151
R1128 B.n130 B.n129 10.6151
R1129 B.n133 B.n130 10.6151
R1130 B.n134 B.n133 10.6151
R1131 B.n137 B.n134 10.6151
R1132 B.n138 B.n137 10.6151
R1133 B.n142 B.n141 10.6151
R1134 B.n145 B.n142 10.6151
R1135 B.n146 B.n145 10.6151
R1136 B.n149 B.n146 10.6151
R1137 B.n150 B.n149 10.6151
R1138 B.n153 B.n150 10.6151
R1139 B.n154 B.n153 10.6151
R1140 B.n157 B.n154 10.6151
R1141 B.n158 B.n157 10.6151
R1142 B.n161 B.n158 10.6151
R1143 B.n163 B.n161 10.6151
R1144 B.n164 B.n163 10.6151
R1145 B.n492 B.n164 10.6151
R1146 B.n282 B.n281 9.36635
R1147 B.n306 B.n305 9.36635
R1148 B.n118 B.n93 9.36635
R1149 B.n141 B.n90 9.36635
R1150 B.n572 B.n0 8.11757
R1151 B.n572 B.n1 8.11757
R1152 B.t6 B.n187 1.37293
R1153 B.n543 B.t2 1.37293
R1154 B.n281 B.n248 1.24928
R1155 B.n305 B.n304 1.24928
R1156 B.n121 B.n93 1.24928
R1157 B.n138 B.n90 1.24928
R1158 VN.n24 VN.n23 174.089
R1159 VN.n49 VN.n48 174.089
R1160 VN.n47 VN.n25 161.3
R1161 VN.n46 VN.n45 161.3
R1162 VN.n44 VN.n26 161.3
R1163 VN.n43 VN.n42 161.3
R1164 VN.n41 VN.n27 161.3
R1165 VN.n40 VN.n39 161.3
R1166 VN.n38 VN.n29 161.3
R1167 VN.n37 VN.n36 161.3
R1168 VN.n35 VN.n30 161.3
R1169 VN.n34 VN.n33 161.3
R1170 VN.n22 VN.n0 161.3
R1171 VN.n21 VN.n20 161.3
R1172 VN.n19 VN.n1 161.3
R1173 VN.n18 VN.n17 161.3
R1174 VN.n15 VN.n2 161.3
R1175 VN.n14 VN.n13 161.3
R1176 VN.n12 VN.n3 161.3
R1177 VN.n11 VN.n10 161.3
R1178 VN.n9 VN.n4 161.3
R1179 VN.n8 VN.n7 161.3
R1180 VN.n6 VN.t3 80.1495
R1181 VN.n32 VN.t5 80.1495
R1182 VN.n6 VN.n5 59.2496
R1183 VN.n32 VN.n31 59.2496
R1184 VN.n10 VN.n9 56.5617
R1185 VN.n15 VN.n14 56.5617
R1186 VN.n36 VN.n35 56.5617
R1187 VN.n41 VN.n40 56.5617
R1188 VN.n3 VN.t6 51.1896
R1189 VN.n5 VN.t9 51.1896
R1190 VN.n16 VN.t4 51.1896
R1191 VN.n23 VN.t2 51.1896
R1192 VN.n29 VN.t1 51.1896
R1193 VN.n31 VN.t8 51.1896
R1194 VN.n28 VN.t7 51.1896
R1195 VN.n48 VN.t0 51.1896
R1196 VN.n21 VN.n1 47.3584
R1197 VN.n46 VN.n26 47.3584
R1198 VN VN.n49 39.26
R1199 VN.n22 VN.n21 33.7956
R1200 VN.n47 VN.n46 33.7956
R1201 VN.n33 VN.n32 27.2704
R1202 VN.n7 VN.n6 27.2704
R1203 VN.n9 VN.n8 24.5923
R1204 VN.n10 VN.n3 24.5923
R1205 VN.n14 VN.n3 24.5923
R1206 VN.n17 VN.n15 24.5923
R1207 VN.n35 VN.n34 24.5923
R1208 VN.n40 VN.n29 24.5923
R1209 VN.n36 VN.n29 24.5923
R1210 VN.n42 VN.n41 24.5923
R1211 VN.n16 VN.n1 18.6903
R1212 VN.n28 VN.n26 18.6903
R1213 VN.n23 VN.n22 11.8046
R1214 VN.n48 VN.n47 11.8046
R1215 VN.n8 VN.n5 5.90254
R1216 VN.n17 VN.n16 5.90254
R1217 VN.n34 VN.n31 5.90254
R1218 VN.n42 VN.n28 5.90254
R1219 VN.n49 VN.n25 0.189894
R1220 VN.n45 VN.n25 0.189894
R1221 VN.n45 VN.n44 0.189894
R1222 VN.n44 VN.n43 0.189894
R1223 VN.n43 VN.n27 0.189894
R1224 VN.n39 VN.n27 0.189894
R1225 VN.n39 VN.n38 0.189894
R1226 VN.n38 VN.n37 0.189894
R1227 VN.n37 VN.n30 0.189894
R1228 VN.n33 VN.n30 0.189894
R1229 VN.n7 VN.n4 0.189894
R1230 VN.n11 VN.n4 0.189894
R1231 VN.n12 VN.n11 0.189894
R1232 VN.n13 VN.n12 0.189894
R1233 VN.n13 VN.n2 0.189894
R1234 VN.n18 VN.n2 0.189894
R1235 VN.n19 VN.n18 0.189894
R1236 VN.n20 VN.n19 0.189894
R1237 VN.n20 VN.n0 0.189894
R1238 VN.n24 VN.n0 0.189894
R1239 VN VN.n24 0.0516364
R1240 VDD2.n1 VDD2.t6 89.0633
R1241 VDD2.n4 VDD2.t9 87.667
R1242 VDD2.n3 VDD2.n2 81.4325
R1243 VDD2 VDD2.n7 81.4298
R1244 VDD2.n6 VDD2.n5 80.4407
R1245 VDD2.n1 VDD2.n0 80.4405
R1246 VDD2.n4 VDD2.n3 32.711
R1247 VDD2.n7 VDD2.t1 7.22678
R1248 VDD2.n7 VDD2.t4 7.22678
R1249 VDD2.n5 VDD2.t2 7.22678
R1250 VDD2.n5 VDD2.t8 7.22678
R1251 VDD2.n2 VDD2.t5 7.22678
R1252 VDD2.n2 VDD2.t7 7.22678
R1253 VDD2.n0 VDD2.t0 7.22678
R1254 VDD2.n0 VDD2.t3 7.22678
R1255 VDD2.n6 VDD2.n4 1.39705
R1256 VDD2 VDD2.n6 0.407828
R1257 VDD2.n3 VDD2.n1 0.294292
C0 VTAIL VDD1 5.08158f
C1 VN VDD2 2.37089f
C2 VTAIL VP 3.0142f
C3 VP VDD1 2.63424f
C4 VTAIL VN 3.00001f
C5 VTAIL VDD2 5.12535f
C6 VN VDD1 0.156141f
C7 VP VN 4.75656f
C8 VDD2 VDD1 1.33562f
C9 VP VDD2 0.422008f
C10 VDD2 B 3.994851f
C11 VDD1 B 3.96555f
C12 VTAIL B 3.305573f
C13 VN B 11.05412f
C14 VP B 9.529514f
C15 VDD2.t6 B 0.476477f
C16 VDD2.t0 B 0.050769f
C17 VDD2.t3 B 0.050769f
C18 VDD2.n0 B 0.37071f
C19 VDD2.n1 B 0.621262f
C20 VDD2.t5 B 0.050769f
C21 VDD2.t7 B 0.050769f
C22 VDD2.n2 B 0.375126f
C23 VDD2.n3 B 1.54604f
C24 VDD2.t9 B 0.471386f
C25 VDD2.n4 B 1.71588f
C26 VDD2.t2 B 0.050769f
C27 VDD2.t8 B 0.050769f
C28 VDD2.n5 B 0.370711f
C29 VDD2.n6 B 0.308312f
C30 VDD2.t1 B 0.050769f
C31 VDD2.t4 B 0.050769f
C32 VDD2.n7 B 0.375104f
C33 VN.n0 B 0.037198f
C34 VN.t2 B 0.32364f
C35 VN.n1 B 0.061789f
C36 VN.n2 B 0.037198f
C37 VN.t6 B 0.32364f
C38 VN.n3 B 0.191801f
C39 VN.n4 B 0.037198f
C40 VN.t9 B 0.32364f
C41 VN.n5 B 0.208076f
C42 VN.t3 B 0.422359f
C43 VN.n6 B 0.225863f
C44 VN.n7 B 0.195538f
C45 VN.n8 B 0.043099f
C46 VN.n9 B 0.047898f
C47 VN.n10 B 0.060247f
C48 VN.n11 B 0.037198f
C49 VN.n12 B 0.037198f
C50 VN.n13 B 0.037198f
C51 VN.n14 B 0.060247f
C52 VN.n15 B 0.047898f
C53 VN.t4 B 0.32364f
C54 VN.n16 B 0.156875f
C55 VN.n17 B 0.043099f
C56 VN.n18 B 0.037198f
C57 VN.n19 B 0.037198f
C58 VN.n20 B 0.037198f
C59 VN.n21 B 0.032434f
C60 VN.n22 B 0.057021f
C61 VN.n23 B 0.222681f
C62 VN.n24 B 0.034044f
C63 VN.n25 B 0.037198f
C64 VN.t0 B 0.32364f
C65 VN.n26 B 0.061789f
C66 VN.n27 B 0.037198f
C67 VN.t7 B 0.32364f
C68 VN.n28 B 0.156875f
C69 VN.t1 B 0.32364f
C70 VN.n29 B 0.191801f
C71 VN.n30 B 0.037198f
C72 VN.t8 B 0.32364f
C73 VN.n31 B 0.208076f
C74 VN.t5 B 0.422359f
C75 VN.n32 B 0.225863f
C76 VN.n33 B 0.195538f
C77 VN.n34 B 0.043099f
C78 VN.n35 B 0.047898f
C79 VN.n36 B 0.060247f
C80 VN.n37 B 0.037198f
C81 VN.n38 B 0.037198f
C82 VN.n39 B 0.037198f
C83 VN.n40 B 0.060247f
C84 VN.n41 B 0.047898f
C85 VN.n42 B 0.043099f
C86 VN.n43 B 0.037198f
C87 VN.n44 B 0.037198f
C88 VN.n45 B 0.037198f
C89 VN.n46 B 0.032434f
C90 VN.n47 B 0.057021f
C91 VN.n48 B 0.222681f
C92 VN.n49 B 1.37489f
C93 VTAIL.t5 B 0.067643f
C94 VTAIL.t8 B 0.067643f
C95 VTAIL.n0 B 0.435527f
C96 VTAIL.n1 B 0.474023f
C97 VTAIL.t16 B 0.56378f
C98 VTAIL.n2 B 0.55954f
C99 VTAIL.t13 B 0.067643f
C100 VTAIL.t11 B 0.067643f
C101 VTAIL.n3 B 0.435527f
C102 VTAIL.n4 B 0.526308f
C103 VTAIL.t12 B 0.067643f
C104 VTAIL.t17 B 0.067643f
C105 VTAIL.n5 B 0.435527f
C106 VTAIL.n6 B 1.32904f
C107 VTAIL.t7 B 0.067643f
C108 VTAIL.t1 B 0.067643f
C109 VTAIL.n7 B 0.435529f
C110 VTAIL.n8 B 1.32903f
C111 VTAIL.t6 B 0.067643f
C112 VTAIL.t0 B 0.067643f
C113 VTAIL.n9 B 0.435529f
C114 VTAIL.n10 B 0.526306f
C115 VTAIL.t9 B 0.563782f
C116 VTAIL.n11 B 0.559538f
C117 VTAIL.t18 B 0.067643f
C118 VTAIL.t14 B 0.067643f
C119 VTAIL.n12 B 0.435529f
C120 VTAIL.n13 B 0.503309f
C121 VTAIL.t10 B 0.067643f
C122 VTAIL.t19 B 0.067643f
C123 VTAIL.n14 B 0.435529f
C124 VTAIL.n15 B 0.526306f
C125 VTAIL.t15 B 0.56378f
C126 VTAIL.n16 B 1.24468f
C127 VTAIL.t3 B 0.56378f
C128 VTAIL.n17 B 1.24468f
C129 VTAIL.t2 B 0.067643f
C130 VTAIL.t4 B 0.067643f
C131 VTAIL.n18 B 0.435527f
C132 VTAIL.n19 B 0.415013f
C133 VDD1.t3 B 0.4836f
C134 VDD1.t2 B 0.051528f
C135 VDD1.t8 B 0.051528f
C136 VDD1.n0 B 0.376252f
C137 VDD1.n1 B 0.637374f
C138 VDD1.t5 B 0.483599f
C139 VDD1.t7 B 0.051528f
C140 VDD1.t4 B 0.051528f
C141 VDD1.n2 B 0.376251f
C142 VDD1.n3 B 0.630548f
C143 VDD1.t1 B 0.051528f
C144 VDD1.t0 B 0.051528f
C145 VDD1.n4 B 0.380733f
C146 VDD1.n5 B 1.65023f
C147 VDD1.t6 B 0.051528f
C148 VDD1.t9 B 0.051528f
C149 VDD1.n6 B 0.376251f
C150 VDD1.n7 B 1.78585f
C151 VP.n0 B 0.038122f
C152 VP.t3 B 0.331686f
C153 VP.n1 B 0.063325f
C154 VP.n2 B 0.038122f
C155 VP.t6 B 0.331686f
C156 VP.n3 B 0.19657f
C157 VP.n4 B 0.038122f
C158 VP.t2 B 0.331686f
C159 VP.n5 B 0.160775f
C160 VP.n6 B 0.038122f
C161 VP.t7 B 0.331686f
C162 VP.n7 B 0.228217f
C163 VP.n8 B 0.038122f
C164 VP.t4 B 0.331686f
C165 VP.n9 B 0.063325f
C166 VP.n10 B 0.038122f
C167 VP.t9 B 0.331686f
C168 VP.n11 B 0.19657f
C169 VP.n12 B 0.038122f
C170 VP.t5 B 0.331686f
C171 VP.n13 B 0.213249f
C172 VP.t1 B 0.432859f
C173 VP.n14 B 0.231479f
C174 VP.n15 B 0.2004f
C175 VP.n16 B 0.044171f
C176 VP.n17 B 0.049088f
C177 VP.n18 B 0.061745f
C178 VP.n19 B 0.038122f
C179 VP.n20 B 0.038122f
C180 VP.n21 B 0.038122f
C181 VP.n22 B 0.061745f
C182 VP.n23 B 0.049088f
C183 VP.t0 B 0.331686f
C184 VP.n24 B 0.160775f
C185 VP.n25 B 0.044171f
C186 VP.n26 B 0.038122f
C187 VP.n27 B 0.038122f
C188 VP.n28 B 0.038122f
C189 VP.n29 B 0.03324f
C190 VP.n30 B 0.058439f
C191 VP.n31 B 0.228217f
C192 VP.n32 B 1.38392f
C193 VP.n33 B 1.41927f
C194 VP.n34 B 0.038122f
C195 VP.n35 B 0.058439f
C196 VP.n36 B 0.03324f
C197 VP.n37 B 0.063325f
C198 VP.n38 B 0.038122f
C199 VP.n39 B 0.038122f
C200 VP.n40 B 0.044171f
C201 VP.n41 B 0.049088f
C202 VP.n42 B 0.061745f
C203 VP.n43 B 0.038122f
C204 VP.n44 B 0.038122f
C205 VP.n45 B 0.038122f
C206 VP.n46 B 0.061745f
C207 VP.n47 B 0.049088f
C208 VP.t8 B 0.331686f
C209 VP.n48 B 0.160775f
C210 VP.n49 B 0.044171f
C211 VP.n50 B 0.038122f
C212 VP.n51 B 0.038122f
C213 VP.n52 B 0.038122f
C214 VP.n53 B 0.03324f
C215 VP.n54 B 0.058439f
C216 VP.n55 B 0.228217f
C217 VP.n56 B 0.03489f
.ends

