* NGSPICE file created from diff_pair_sample_0181.ext - technology: sky130A

.subckt diff_pair_sample_0181 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=4.1262 ps=21.94 w=10.58 l=1.03
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=4.1262 ps=21.94 w=10.58 l=1.03
X2 B.t11 B.t9 B.t10 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=0 ps=0 w=10.58 l=1.03
X3 B.t8 B.t6 B.t7 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=0 ps=0 w=10.58 l=1.03
X4 VDD1.t0 VP.t1 VTAIL.t3 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=4.1262 ps=21.94 w=10.58 l=1.03
X5 VDD2.t0 VN.t1 VTAIL.t2 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=4.1262 ps=21.94 w=10.58 l=1.03
X6 B.t5 B.t3 B.t4 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=0 ps=0 w=10.58 l=1.03
X7 B.t2 B.t0 B.t1 w_n1514_n3088# sky130_fd_pr__pfet_01v8 ad=4.1262 pd=21.94 as=0 ps=0 w=10.58 l=1.03
R0 VN VN.t1 486.803
R1 VN VN.t0 447.041
R2 VTAIL.n226 VTAIL.n174 756.745
R3 VTAIL.n52 VTAIL.n0 756.745
R4 VTAIL.n168 VTAIL.n116 756.745
R5 VTAIL.n110 VTAIL.n58 756.745
R6 VTAIL.n193 VTAIL.n192 585
R7 VTAIL.n190 VTAIL.n189 585
R8 VTAIL.n199 VTAIL.n198 585
R9 VTAIL.n201 VTAIL.n200 585
R10 VTAIL.n186 VTAIL.n185 585
R11 VTAIL.n207 VTAIL.n206 585
R12 VTAIL.n210 VTAIL.n209 585
R13 VTAIL.n208 VTAIL.n182 585
R14 VTAIL.n215 VTAIL.n181 585
R15 VTAIL.n217 VTAIL.n216 585
R16 VTAIL.n219 VTAIL.n218 585
R17 VTAIL.n178 VTAIL.n177 585
R18 VTAIL.n225 VTAIL.n224 585
R19 VTAIL.n227 VTAIL.n226 585
R20 VTAIL.n19 VTAIL.n18 585
R21 VTAIL.n16 VTAIL.n15 585
R22 VTAIL.n25 VTAIL.n24 585
R23 VTAIL.n27 VTAIL.n26 585
R24 VTAIL.n12 VTAIL.n11 585
R25 VTAIL.n33 VTAIL.n32 585
R26 VTAIL.n36 VTAIL.n35 585
R27 VTAIL.n34 VTAIL.n8 585
R28 VTAIL.n41 VTAIL.n7 585
R29 VTAIL.n43 VTAIL.n42 585
R30 VTAIL.n45 VTAIL.n44 585
R31 VTAIL.n4 VTAIL.n3 585
R32 VTAIL.n51 VTAIL.n50 585
R33 VTAIL.n53 VTAIL.n52 585
R34 VTAIL.n169 VTAIL.n168 585
R35 VTAIL.n167 VTAIL.n166 585
R36 VTAIL.n120 VTAIL.n119 585
R37 VTAIL.n161 VTAIL.n160 585
R38 VTAIL.n159 VTAIL.n158 585
R39 VTAIL.n157 VTAIL.n123 585
R40 VTAIL.n127 VTAIL.n124 585
R41 VTAIL.n152 VTAIL.n151 585
R42 VTAIL.n150 VTAIL.n149 585
R43 VTAIL.n129 VTAIL.n128 585
R44 VTAIL.n144 VTAIL.n143 585
R45 VTAIL.n142 VTAIL.n141 585
R46 VTAIL.n133 VTAIL.n132 585
R47 VTAIL.n136 VTAIL.n135 585
R48 VTAIL.n111 VTAIL.n110 585
R49 VTAIL.n109 VTAIL.n108 585
R50 VTAIL.n62 VTAIL.n61 585
R51 VTAIL.n103 VTAIL.n102 585
R52 VTAIL.n101 VTAIL.n100 585
R53 VTAIL.n99 VTAIL.n65 585
R54 VTAIL.n69 VTAIL.n66 585
R55 VTAIL.n94 VTAIL.n93 585
R56 VTAIL.n92 VTAIL.n91 585
R57 VTAIL.n71 VTAIL.n70 585
R58 VTAIL.n86 VTAIL.n85 585
R59 VTAIL.n84 VTAIL.n83 585
R60 VTAIL.n75 VTAIL.n74 585
R61 VTAIL.n78 VTAIL.n77 585
R62 VTAIL.t0 VTAIL.n134 329.038
R63 VTAIL.t2 VTAIL.n76 329.038
R64 VTAIL.t1 VTAIL.n191 329.038
R65 VTAIL.t3 VTAIL.n17 329.038
R66 VTAIL.n192 VTAIL.n189 171.744
R67 VTAIL.n199 VTAIL.n189 171.744
R68 VTAIL.n200 VTAIL.n199 171.744
R69 VTAIL.n200 VTAIL.n185 171.744
R70 VTAIL.n207 VTAIL.n185 171.744
R71 VTAIL.n209 VTAIL.n207 171.744
R72 VTAIL.n209 VTAIL.n208 171.744
R73 VTAIL.n208 VTAIL.n181 171.744
R74 VTAIL.n217 VTAIL.n181 171.744
R75 VTAIL.n218 VTAIL.n217 171.744
R76 VTAIL.n218 VTAIL.n177 171.744
R77 VTAIL.n225 VTAIL.n177 171.744
R78 VTAIL.n226 VTAIL.n225 171.744
R79 VTAIL.n18 VTAIL.n15 171.744
R80 VTAIL.n25 VTAIL.n15 171.744
R81 VTAIL.n26 VTAIL.n25 171.744
R82 VTAIL.n26 VTAIL.n11 171.744
R83 VTAIL.n33 VTAIL.n11 171.744
R84 VTAIL.n35 VTAIL.n33 171.744
R85 VTAIL.n35 VTAIL.n34 171.744
R86 VTAIL.n34 VTAIL.n7 171.744
R87 VTAIL.n43 VTAIL.n7 171.744
R88 VTAIL.n44 VTAIL.n43 171.744
R89 VTAIL.n44 VTAIL.n3 171.744
R90 VTAIL.n51 VTAIL.n3 171.744
R91 VTAIL.n52 VTAIL.n51 171.744
R92 VTAIL.n168 VTAIL.n167 171.744
R93 VTAIL.n167 VTAIL.n119 171.744
R94 VTAIL.n160 VTAIL.n119 171.744
R95 VTAIL.n160 VTAIL.n159 171.744
R96 VTAIL.n159 VTAIL.n123 171.744
R97 VTAIL.n127 VTAIL.n123 171.744
R98 VTAIL.n151 VTAIL.n127 171.744
R99 VTAIL.n151 VTAIL.n150 171.744
R100 VTAIL.n150 VTAIL.n128 171.744
R101 VTAIL.n143 VTAIL.n128 171.744
R102 VTAIL.n143 VTAIL.n142 171.744
R103 VTAIL.n142 VTAIL.n132 171.744
R104 VTAIL.n135 VTAIL.n132 171.744
R105 VTAIL.n110 VTAIL.n109 171.744
R106 VTAIL.n109 VTAIL.n61 171.744
R107 VTAIL.n102 VTAIL.n61 171.744
R108 VTAIL.n102 VTAIL.n101 171.744
R109 VTAIL.n101 VTAIL.n65 171.744
R110 VTAIL.n69 VTAIL.n65 171.744
R111 VTAIL.n93 VTAIL.n69 171.744
R112 VTAIL.n93 VTAIL.n92 171.744
R113 VTAIL.n92 VTAIL.n70 171.744
R114 VTAIL.n85 VTAIL.n70 171.744
R115 VTAIL.n85 VTAIL.n84 171.744
R116 VTAIL.n84 VTAIL.n74 171.744
R117 VTAIL.n77 VTAIL.n74 171.744
R118 VTAIL.n192 VTAIL.t1 85.8723
R119 VTAIL.n18 VTAIL.t3 85.8723
R120 VTAIL.n135 VTAIL.t0 85.8723
R121 VTAIL.n77 VTAIL.t2 85.8723
R122 VTAIL.n231 VTAIL.n230 30.246
R123 VTAIL.n57 VTAIL.n56 30.246
R124 VTAIL.n173 VTAIL.n172 30.246
R125 VTAIL.n115 VTAIL.n114 30.246
R126 VTAIL.n115 VTAIL.n57 23.8496
R127 VTAIL.n231 VTAIL.n173 22.6772
R128 VTAIL.n216 VTAIL.n215 13.1884
R129 VTAIL.n42 VTAIL.n41 13.1884
R130 VTAIL.n158 VTAIL.n157 13.1884
R131 VTAIL.n100 VTAIL.n99 13.1884
R132 VTAIL.n214 VTAIL.n182 12.8005
R133 VTAIL.n219 VTAIL.n180 12.8005
R134 VTAIL.n40 VTAIL.n8 12.8005
R135 VTAIL.n45 VTAIL.n6 12.8005
R136 VTAIL.n161 VTAIL.n122 12.8005
R137 VTAIL.n156 VTAIL.n124 12.8005
R138 VTAIL.n103 VTAIL.n64 12.8005
R139 VTAIL.n98 VTAIL.n66 12.8005
R140 VTAIL.n211 VTAIL.n210 12.0247
R141 VTAIL.n220 VTAIL.n178 12.0247
R142 VTAIL.n37 VTAIL.n36 12.0247
R143 VTAIL.n46 VTAIL.n4 12.0247
R144 VTAIL.n162 VTAIL.n120 12.0247
R145 VTAIL.n153 VTAIL.n152 12.0247
R146 VTAIL.n104 VTAIL.n62 12.0247
R147 VTAIL.n95 VTAIL.n94 12.0247
R148 VTAIL.n206 VTAIL.n184 11.249
R149 VTAIL.n224 VTAIL.n223 11.249
R150 VTAIL.n32 VTAIL.n10 11.249
R151 VTAIL.n50 VTAIL.n49 11.249
R152 VTAIL.n166 VTAIL.n165 11.249
R153 VTAIL.n149 VTAIL.n126 11.249
R154 VTAIL.n108 VTAIL.n107 11.249
R155 VTAIL.n91 VTAIL.n68 11.249
R156 VTAIL.n193 VTAIL.n191 10.7239
R157 VTAIL.n19 VTAIL.n17 10.7239
R158 VTAIL.n136 VTAIL.n134 10.7239
R159 VTAIL.n78 VTAIL.n76 10.7239
R160 VTAIL.n205 VTAIL.n186 10.4732
R161 VTAIL.n227 VTAIL.n176 10.4732
R162 VTAIL.n31 VTAIL.n12 10.4732
R163 VTAIL.n53 VTAIL.n2 10.4732
R164 VTAIL.n169 VTAIL.n118 10.4732
R165 VTAIL.n148 VTAIL.n129 10.4732
R166 VTAIL.n111 VTAIL.n60 10.4732
R167 VTAIL.n90 VTAIL.n71 10.4732
R168 VTAIL.n202 VTAIL.n201 9.69747
R169 VTAIL.n228 VTAIL.n174 9.69747
R170 VTAIL.n28 VTAIL.n27 9.69747
R171 VTAIL.n54 VTAIL.n0 9.69747
R172 VTAIL.n170 VTAIL.n116 9.69747
R173 VTAIL.n145 VTAIL.n144 9.69747
R174 VTAIL.n112 VTAIL.n58 9.69747
R175 VTAIL.n87 VTAIL.n86 9.69747
R176 VTAIL.n230 VTAIL.n229 9.45567
R177 VTAIL.n56 VTAIL.n55 9.45567
R178 VTAIL.n172 VTAIL.n171 9.45567
R179 VTAIL.n114 VTAIL.n113 9.45567
R180 VTAIL.n229 VTAIL.n228 9.3005
R181 VTAIL.n176 VTAIL.n175 9.3005
R182 VTAIL.n223 VTAIL.n222 9.3005
R183 VTAIL.n221 VTAIL.n220 9.3005
R184 VTAIL.n180 VTAIL.n179 9.3005
R185 VTAIL.n195 VTAIL.n194 9.3005
R186 VTAIL.n197 VTAIL.n196 9.3005
R187 VTAIL.n188 VTAIL.n187 9.3005
R188 VTAIL.n203 VTAIL.n202 9.3005
R189 VTAIL.n205 VTAIL.n204 9.3005
R190 VTAIL.n184 VTAIL.n183 9.3005
R191 VTAIL.n212 VTAIL.n211 9.3005
R192 VTAIL.n214 VTAIL.n213 9.3005
R193 VTAIL.n55 VTAIL.n54 9.3005
R194 VTAIL.n2 VTAIL.n1 9.3005
R195 VTAIL.n49 VTAIL.n48 9.3005
R196 VTAIL.n47 VTAIL.n46 9.3005
R197 VTAIL.n6 VTAIL.n5 9.3005
R198 VTAIL.n21 VTAIL.n20 9.3005
R199 VTAIL.n23 VTAIL.n22 9.3005
R200 VTAIL.n14 VTAIL.n13 9.3005
R201 VTAIL.n29 VTAIL.n28 9.3005
R202 VTAIL.n31 VTAIL.n30 9.3005
R203 VTAIL.n10 VTAIL.n9 9.3005
R204 VTAIL.n38 VTAIL.n37 9.3005
R205 VTAIL.n40 VTAIL.n39 9.3005
R206 VTAIL.n138 VTAIL.n137 9.3005
R207 VTAIL.n140 VTAIL.n139 9.3005
R208 VTAIL.n131 VTAIL.n130 9.3005
R209 VTAIL.n146 VTAIL.n145 9.3005
R210 VTAIL.n148 VTAIL.n147 9.3005
R211 VTAIL.n126 VTAIL.n125 9.3005
R212 VTAIL.n154 VTAIL.n153 9.3005
R213 VTAIL.n156 VTAIL.n155 9.3005
R214 VTAIL.n171 VTAIL.n170 9.3005
R215 VTAIL.n118 VTAIL.n117 9.3005
R216 VTAIL.n165 VTAIL.n164 9.3005
R217 VTAIL.n163 VTAIL.n162 9.3005
R218 VTAIL.n122 VTAIL.n121 9.3005
R219 VTAIL.n80 VTAIL.n79 9.3005
R220 VTAIL.n82 VTAIL.n81 9.3005
R221 VTAIL.n73 VTAIL.n72 9.3005
R222 VTAIL.n88 VTAIL.n87 9.3005
R223 VTAIL.n90 VTAIL.n89 9.3005
R224 VTAIL.n68 VTAIL.n67 9.3005
R225 VTAIL.n96 VTAIL.n95 9.3005
R226 VTAIL.n98 VTAIL.n97 9.3005
R227 VTAIL.n113 VTAIL.n112 9.3005
R228 VTAIL.n60 VTAIL.n59 9.3005
R229 VTAIL.n107 VTAIL.n106 9.3005
R230 VTAIL.n105 VTAIL.n104 9.3005
R231 VTAIL.n64 VTAIL.n63 9.3005
R232 VTAIL.n198 VTAIL.n188 8.92171
R233 VTAIL.n24 VTAIL.n14 8.92171
R234 VTAIL.n141 VTAIL.n131 8.92171
R235 VTAIL.n83 VTAIL.n73 8.92171
R236 VTAIL.n197 VTAIL.n190 8.14595
R237 VTAIL.n23 VTAIL.n16 8.14595
R238 VTAIL.n140 VTAIL.n133 8.14595
R239 VTAIL.n82 VTAIL.n75 8.14595
R240 VTAIL.n194 VTAIL.n193 7.3702
R241 VTAIL.n20 VTAIL.n19 7.3702
R242 VTAIL.n137 VTAIL.n136 7.3702
R243 VTAIL.n79 VTAIL.n78 7.3702
R244 VTAIL.n194 VTAIL.n190 5.81868
R245 VTAIL.n20 VTAIL.n16 5.81868
R246 VTAIL.n137 VTAIL.n133 5.81868
R247 VTAIL.n79 VTAIL.n75 5.81868
R248 VTAIL.n198 VTAIL.n197 5.04292
R249 VTAIL.n24 VTAIL.n23 5.04292
R250 VTAIL.n141 VTAIL.n140 5.04292
R251 VTAIL.n83 VTAIL.n82 5.04292
R252 VTAIL.n201 VTAIL.n188 4.26717
R253 VTAIL.n230 VTAIL.n174 4.26717
R254 VTAIL.n27 VTAIL.n14 4.26717
R255 VTAIL.n56 VTAIL.n0 4.26717
R256 VTAIL.n172 VTAIL.n116 4.26717
R257 VTAIL.n144 VTAIL.n131 4.26717
R258 VTAIL.n114 VTAIL.n58 4.26717
R259 VTAIL.n86 VTAIL.n73 4.26717
R260 VTAIL.n202 VTAIL.n186 3.49141
R261 VTAIL.n228 VTAIL.n227 3.49141
R262 VTAIL.n28 VTAIL.n12 3.49141
R263 VTAIL.n54 VTAIL.n53 3.49141
R264 VTAIL.n170 VTAIL.n169 3.49141
R265 VTAIL.n145 VTAIL.n129 3.49141
R266 VTAIL.n112 VTAIL.n111 3.49141
R267 VTAIL.n87 VTAIL.n71 3.49141
R268 VTAIL.n206 VTAIL.n205 2.71565
R269 VTAIL.n224 VTAIL.n176 2.71565
R270 VTAIL.n32 VTAIL.n31 2.71565
R271 VTAIL.n50 VTAIL.n2 2.71565
R272 VTAIL.n166 VTAIL.n118 2.71565
R273 VTAIL.n149 VTAIL.n148 2.71565
R274 VTAIL.n108 VTAIL.n60 2.71565
R275 VTAIL.n91 VTAIL.n90 2.71565
R276 VTAIL.n195 VTAIL.n191 2.41282
R277 VTAIL.n21 VTAIL.n17 2.41282
R278 VTAIL.n138 VTAIL.n134 2.41282
R279 VTAIL.n80 VTAIL.n76 2.41282
R280 VTAIL.n210 VTAIL.n184 1.93989
R281 VTAIL.n223 VTAIL.n178 1.93989
R282 VTAIL.n36 VTAIL.n10 1.93989
R283 VTAIL.n49 VTAIL.n4 1.93989
R284 VTAIL.n165 VTAIL.n120 1.93989
R285 VTAIL.n152 VTAIL.n126 1.93989
R286 VTAIL.n107 VTAIL.n62 1.93989
R287 VTAIL.n94 VTAIL.n68 1.93989
R288 VTAIL.n211 VTAIL.n182 1.16414
R289 VTAIL.n220 VTAIL.n219 1.16414
R290 VTAIL.n37 VTAIL.n8 1.16414
R291 VTAIL.n46 VTAIL.n45 1.16414
R292 VTAIL.n162 VTAIL.n161 1.16414
R293 VTAIL.n153 VTAIL.n124 1.16414
R294 VTAIL.n104 VTAIL.n103 1.16414
R295 VTAIL.n95 VTAIL.n66 1.16414
R296 VTAIL.n173 VTAIL.n115 1.05653
R297 VTAIL VTAIL.n57 0.821621
R298 VTAIL.n215 VTAIL.n214 0.388379
R299 VTAIL.n216 VTAIL.n180 0.388379
R300 VTAIL.n41 VTAIL.n40 0.388379
R301 VTAIL.n42 VTAIL.n6 0.388379
R302 VTAIL.n158 VTAIL.n122 0.388379
R303 VTAIL.n157 VTAIL.n156 0.388379
R304 VTAIL.n100 VTAIL.n64 0.388379
R305 VTAIL.n99 VTAIL.n98 0.388379
R306 VTAIL VTAIL.n231 0.235414
R307 VTAIL.n196 VTAIL.n195 0.155672
R308 VTAIL.n196 VTAIL.n187 0.155672
R309 VTAIL.n203 VTAIL.n187 0.155672
R310 VTAIL.n204 VTAIL.n203 0.155672
R311 VTAIL.n204 VTAIL.n183 0.155672
R312 VTAIL.n212 VTAIL.n183 0.155672
R313 VTAIL.n213 VTAIL.n212 0.155672
R314 VTAIL.n213 VTAIL.n179 0.155672
R315 VTAIL.n221 VTAIL.n179 0.155672
R316 VTAIL.n222 VTAIL.n221 0.155672
R317 VTAIL.n222 VTAIL.n175 0.155672
R318 VTAIL.n229 VTAIL.n175 0.155672
R319 VTAIL.n22 VTAIL.n21 0.155672
R320 VTAIL.n22 VTAIL.n13 0.155672
R321 VTAIL.n29 VTAIL.n13 0.155672
R322 VTAIL.n30 VTAIL.n29 0.155672
R323 VTAIL.n30 VTAIL.n9 0.155672
R324 VTAIL.n38 VTAIL.n9 0.155672
R325 VTAIL.n39 VTAIL.n38 0.155672
R326 VTAIL.n39 VTAIL.n5 0.155672
R327 VTAIL.n47 VTAIL.n5 0.155672
R328 VTAIL.n48 VTAIL.n47 0.155672
R329 VTAIL.n48 VTAIL.n1 0.155672
R330 VTAIL.n55 VTAIL.n1 0.155672
R331 VTAIL.n171 VTAIL.n117 0.155672
R332 VTAIL.n164 VTAIL.n117 0.155672
R333 VTAIL.n164 VTAIL.n163 0.155672
R334 VTAIL.n163 VTAIL.n121 0.155672
R335 VTAIL.n155 VTAIL.n121 0.155672
R336 VTAIL.n155 VTAIL.n154 0.155672
R337 VTAIL.n154 VTAIL.n125 0.155672
R338 VTAIL.n147 VTAIL.n125 0.155672
R339 VTAIL.n147 VTAIL.n146 0.155672
R340 VTAIL.n146 VTAIL.n130 0.155672
R341 VTAIL.n139 VTAIL.n130 0.155672
R342 VTAIL.n139 VTAIL.n138 0.155672
R343 VTAIL.n113 VTAIL.n59 0.155672
R344 VTAIL.n106 VTAIL.n59 0.155672
R345 VTAIL.n106 VTAIL.n105 0.155672
R346 VTAIL.n105 VTAIL.n63 0.155672
R347 VTAIL.n97 VTAIL.n63 0.155672
R348 VTAIL.n97 VTAIL.n96 0.155672
R349 VTAIL.n96 VTAIL.n67 0.155672
R350 VTAIL.n89 VTAIL.n67 0.155672
R351 VTAIL.n89 VTAIL.n88 0.155672
R352 VTAIL.n88 VTAIL.n72 0.155672
R353 VTAIL.n81 VTAIL.n72 0.155672
R354 VTAIL.n81 VTAIL.n80 0.155672
R355 VDD2.n109 VDD2.n57 756.745
R356 VDD2.n52 VDD2.n0 756.745
R357 VDD2.n110 VDD2.n109 585
R358 VDD2.n108 VDD2.n107 585
R359 VDD2.n61 VDD2.n60 585
R360 VDD2.n102 VDD2.n101 585
R361 VDD2.n100 VDD2.n99 585
R362 VDD2.n98 VDD2.n64 585
R363 VDD2.n68 VDD2.n65 585
R364 VDD2.n93 VDD2.n92 585
R365 VDD2.n91 VDD2.n90 585
R366 VDD2.n70 VDD2.n69 585
R367 VDD2.n85 VDD2.n84 585
R368 VDD2.n83 VDD2.n82 585
R369 VDD2.n74 VDD2.n73 585
R370 VDD2.n77 VDD2.n76 585
R371 VDD2.n19 VDD2.n18 585
R372 VDD2.n16 VDD2.n15 585
R373 VDD2.n25 VDD2.n24 585
R374 VDD2.n27 VDD2.n26 585
R375 VDD2.n12 VDD2.n11 585
R376 VDD2.n33 VDD2.n32 585
R377 VDD2.n36 VDD2.n35 585
R378 VDD2.n34 VDD2.n8 585
R379 VDD2.n41 VDD2.n7 585
R380 VDD2.n43 VDD2.n42 585
R381 VDD2.n45 VDD2.n44 585
R382 VDD2.n4 VDD2.n3 585
R383 VDD2.n51 VDD2.n50 585
R384 VDD2.n53 VDD2.n52 585
R385 VDD2.t0 VDD2.n75 329.038
R386 VDD2.t1 VDD2.n17 329.038
R387 VDD2.n109 VDD2.n108 171.744
R388 VDD2.n108 VDD2.n60 171.744
R389 VDD2.n101 VDD2.n60 171.744
R390 VDD2.n101 VDD2.n100 171.744
R391 VDD2.n100 VDD2.n64 171.744
R392 VDD2.n68 VDD2.n64 171.744
R393 VDD2.n92 VDD2.n68 171.744
R394 VDD2.n92 VDD2.n91 171.744
R395 VDD2.n91 VDD2.n69 171.744
R396 VDD2.n84 VDD2.n69 171.744
R397 VDD2.n84 VDD2.n83 171.744
R398 VDD2.n83 VDD2.n73 171.744
R399 VDD2.n76 VDD2.n73 171.744
R400 VDD2.n18 VDD2.n15 171.744
R401 VDD2.n25 VDD2.n15 171.744
R402 VDD2.n26 VDD2.n25 171.744
R403 VDD2.n26 VDD2.n11 171.744
R404 VDD2.n33 VDD2.n11 171.744
R405 VDD2.n35 VDD2.n33 171.744
R406 VDD2.n35 VDD2.n34 171.744
R407 VDD2.n34 VDD2.n7 171.744
R408 VDD2.n43 VDD2.n7 171.744
R409 VDD2.n44 VDD2.n43 171.744
R410 VDD2.n44 VDD2.n3 171.744
R411 VDD2.n51 VDD2.n3 171.744
R412 VDD2.n52 VDD2.n51 171.744
R413 VDD2.n76 VDD2.t0 85.8723
R414 VDD2.n18 VDD2.t1 85.8723
R415 VDD2.n114 VDD2.n56 82.0669
R416 VDD2.n114 VDD2.n113 46.9247
R417 VDD2.n99 VDD2.n98 13.1884
R418 VDD2.n42 VDD2.n41 13.1884
R419 VDD2.n102 VDD2.n63 12.8005
R420 VDD2.n97 VDD2.n65 12.8005
R421 VDD2.n40 VDD2.n8 12.8005
R422 VDD2.n45 VDD2.n6 12.8005
R423 VDD2.n103 VDD2.n61 12.0247
R424 VDD2.n94 VDD2.n93 12.0247
R425 VDD2.n37 VDD2.n36 12.0247
R426 VDD2.n46 VDD2.n4 12.0247
R427 VDD2.n107 VDD2.n106 11.249
R428 VDD2.n90 VDD2.n67 11.249
R429 VDD2.n32 VDD2.n10 11.249
R430 VDD2.n50 VDD2.n49 11.249
R431 VDD2.n77 VDD2.n75 10.7239
R432 VDD2.n19 VDD2.n17 10.7239
R433 VDD2.n110 VDD2.n59 10.4732
R434 VDD2.n89 VDD2.n70 10.4732
R435 VDD2.n31 VDD2.n12 10.4732
R436 VDD2.n53 VDD2.n2 10.4732
R437 VDD2.n111 VDD2.n57 9.69747
R438 VDD2.n86 VDD2.n85 9.69747
R439 VDD2.n28 VDD2.n27 9.69747
R440 VDD2.n54 VDD2.n0 9.69747
R441 VDD2.n113 VDD2.n112 9.45567
R442 VDD2.n56 VDD2.n55 9.45567
R443 VDD2.n79 VDD2.n78 9.3005
R444 VDD2.n81 VDD2.n80 9.3005
R445 VDD2.n72 VDD2.n71 9.3005
R446 VDD2.n87 VDD2.n86 9.3005
R447 VDD2.n89 VDD2.n88 9.3005
R448 VDD2.n67 VDD2.n66 9.3005
R449 VDD2.n95 VDD2.n94 9.3005
R450 VDD2.n97 VDD2.n96 9.3005
R451 VDD2.n112 VDD2.n111 9.3005
R452 VDD2.n59 VDD2.n58 9.3005
R453 VDD2.n106 VDD2.n105 9.3005
R454 VDD2.n104 VDD2.n103 9.3005
R455 VDD2.n63 VDD2.n62 9.3005
R456 VDD2.n55 VDD2.n54 9.3005
R457 VDD2.n2 VDD2.n1 9.3005
R458 VDD2.n49 VDD2.n48 9.3005
R459 VDD2.n47 VDD2.n46 9.3005
R460 VDD2.n6 VDD2.n5 9.3005
R461 VDD2.n21 VDD2.n20 9.3005
R462 VDD2.n23 VDD2.n22 9.3005
R463 VDD2.n14 VDD2.n13 9.3005
R464 VDD2.n29 VDD2.n28 9.3005
R465 VDD2.n31 VDD2.n30 9.3005
R466 VDD2.n10 VDD2.n9 9.3005
R467 VDD2.n38 VDD2.n37 9.3005
R468 VDD2.n40 VDD2.n39 9.3005
R469 VDD2.n82 VDD2.n72 8.92171
R470 VDD2.n24 VDD2.n14 8.92171
R471 VDD2.n81 VDD2.n74 8.14595
R472 VDD2.n23 VDD2.n16 8.14595
R473 VDD2.n78 VDD2.n77 7.3702
R474 VDD2.n20 VDD2.n19 7.3702
R475 VDD2.n78 VDD2.n74 5.81868
R476 VDD2.n20 VDD2.n16 5.81868
R477 VDD2.n82 VDD2.n81 5.04292
R478 VDD2.n24 VDD2.n23 5.04292
R479 VDD2.n113 VDD2.n57 4.26717
R480 VDD2.n85 VDD2.n72 4.26717
R481 VDD2.n27 VDD2.n14 4.26717
R482 VDD2.n56 VDD2.n0 4.26717
R483 VDD2.n111 VDD2.n110 3.49141
R484 VDD2.n86 VDD2.n70 3.49141
R485 VDD2.n28 VDD2.n12 3.49141
R486 VDD2.n54 VDD2.n53 3.49141
R487 VDD2.n107 VDD2.n59 2.71565
R488 VDD2.n90 VDD2.n89 2.71565
R489 VDD2.n32 VDD2.n31 2.71565
R490 VDD2.n50 VDD2.n2 2.71565
R491 VDD2.n79 VDD2.n75 2.41282
R492 VDD2.n21 VDD2.n17 2.41282
R493 VDD2.n106 VDD2.n61 1.93989
R494 VDD2.n93 VDD2.n67 1.93989
R495 VDD2.n36 VDD2.n10 1.93989
R496 VDD2.n49 VDD2.n4 1.93989
R497 VDD2.n103 VDD2.n102 1.16414
R498 VDD2.n94 VDD2.n65 1.16414
R499 VDD2.n37 VDD2.n8 1.16414
R500 VDD2.n46 VDD2.n45 1.16414
R501 VDD2.n99 VDD2.n63 0.388379
R502 VDD2.n98 VDD2.n97 0.388379
R503 VDD2.n41 VDD2.n40 0.388379
R504 VDD2.n42 VDD2.n6 0.388379
R505 VDD2 VDD2.n114 0.351793
R506 VDD2.n112 VDD2.n58 0.155672
R507 VDD2.n105 VDD2.n58 0.155672
R508 VDD2.n105 VDD2.n104 0.155672
R509 VDD2.n104 VDD2.n62 0.155672
R510 VDD2.n96 VDD2.n62 0.155672
R511 VDD2.n96 VDD2.n95 0.155672
R512 VDD2.n95 VDD2.n66 0.155672
R513 VDD2.n88 VDD2.n66 0.155672
R514 VDD2.n88 VDD2.n87 0.155672
R515 VDD2.n87 VDD2.n71 0.155672
R516 VDD2.n80 VDD2.n71 0.155672
R517 VDD2.n80 VDD2.n79 0.155672
R518 VDD2.n22 VDD2.n21 0.155672
R519 VDD2.n22 VDD2.n13 0.155672
R520 VDD2.n29 VDD2.n13 0.155672
R521 VDD2.n30 VDD2.n29 0.155672
R522 VDD2.n30 VDD2.n9 0.155672
R523 VDD2.n38 VDD2.n9 0.155672
R524 VDD2.n39 VDD2.n38 0.155672
R525 VDD2.n39 VDD2.n5 0.155672
R526 VDD2.n47 VDD2.n5 0.155672
R527 VDD2.n48 VDD2.n47 0.155672
R528 VDD2.n48 VDD2.n1 0.155672
R529 VDD2.n55 VDD2.n1 0.155672
R530 VP.n0 VP.t0 486.423
R531 VP.n0 VP.t1 446.99
R532 VP VP.n0 0.0516364
R533 VDD1.n52 VDD1.n0 756.745
R534 VDD1.n109 VDD1.n57 756.745
R535 VDD1.n53 VDD1.n52 585
R536 VDD1.n51 VDD1.n50 585
R537 VDD1.n4 VDD1.n3 585
R538 VDD1.n45 VDD1.n44 585
R539 VDD1.n43 VDD1.n42 585
R540 VDD1.n41 VDD1.n7 585
R541 VDD1.n11 VDD1.n8 585
R542 VDD1.n36 VDD1.n35 585
R543 VDD1.n34 VDD1.n33 585
R544 VDD1.n13 VDD1.n12 585
R545 VDD1.n28 VDD1.n27 585
R546 VDD1.n26 VDD1.n25 585
R547 VDD1.n17 VDD1.n16 585
R548 VDD1.n20 VDD1.n19 585
R549 VDD1.n76 VDD1.n75 585
R550 VDD1.n73 VDD1.n72 585
R551 VDD1.n82 VDD1.n81 585
R552 VDD1.n84 VDD1.n83 585
R553 VDD1.n69 VDD1.n68 585
R554 VDD1.n90 VDD1.n89 585
R555 VDD1.n93 VDD1.n92 585
R556 VDD1.n91 VDD1.n65 585
R557 VDD1.n98 VDD1.n64 585
R558 VDD1.n100 VDD1.n99 585
R559 VDD1.n102 VDD1.n101 585
R560 VDD1.n61 VDD1.n60 585
R561 VDD1.n108 VDD1.n107 585
R562 VDD1.n110 VDD1.n109 585
R563 VDD1.t1 VDD1.n18 329.038
R564 VDD1.t0 VDD1.n74 329.038
R565 VDD1.n52 VDD1.n51 171.744
R566 VDD1.n51 VDD1.n3 171.744
R567 VDD1.n44 VDD1.n3 171.744
R568 VDD1.n44 VDD1.n43 171.744
R569 VDD1.n43 VDD1.n7 171.744
R570 VDD1.n11 VDD1.n7 171.744
R571 VDD1.n35 VDD1.n11 171.744
R572 VDD1.n35 VDD1.n34 171.744
R573 VDD1.n34 VDD1.n12 171.744
R574 VDD1.n27 VDD1.n12 171.744
R575 VDD1.n27 VDD1.n26 171.744
R576 VDD1.n26 VDD1.n16 171.744
R577 VDD1.n19 VDD1.n16 171.744
R578 VDD1.n75 VDD1.n72 171.744
R579 VDD1.n82 VDD1.n72 171.744
R580 VDD1.n83 VDD1.n82 171.744
R581 VDD1.n83 VDD1.n68 171.744
R582 VDD1.n90 VDD1.n68 171.744
R583 VDD1.n92 VDD1.n90 171.744
R584 VDD1.n92 VDD1.n91 171.744
R585 VDD1.n91 VDD1.n64 171.744
R586 VDD1.n100 VDD1.n64 171.744
R587 VDD1.n101 VDD1.n100 171.744
R588 VDD1.n101 VDD1.n60 171.744
R589 VDD1.n108 VDD1.n60 171.744
R590 VDD1.n109 VDD1.n108 171.744
R591 VDD1.n19 VDD1.t1 85.8723
R592 VDD1.n75 VDD1.t0 85.8723
R593 VDD1 VDD1.n113 82.8849
R594 VDD1 VDD1.n56 47.276
R595 VDD1.n42 VDD1.n41 13.1884
R596 VDD1.n99 VDD1.n98 13.1884
R597 VDD1.n45 VDD1.n6 12.8005
R598 VDD1.n40 VDD1.n8 12.8005
R599 VDD1.n97 VDD1.n65 12.8005
R600 VDD1.n102 VDD1.n63 12.8005
R601 VDD1.n46 VDD1.n4 12.0247
R602 VDD1.n37 VDD1.n36 12.0247
R603 VDD1.n94 VDD1.n93 12.0247
R604 VDD1.n103 VDD1.n61 12.0247
R605 VDD1.n50 VDD1.n49 11.249
R606 VDD1.n33 VDD1.n10 11.249
R607 VDD1.n89 VDD1.n67 11.249
R608 VDD1.n107 VDD1.n106 11.249
R609 VDD1.n20 VDD1.n18 10.7239
R610 VDD1.n76 VDD1.n74 10.7239
R611 VDD1.n53 VDD1.n2 10.4732
R612 VDD1.n32 VDD1.n13 10.4732
R613 VDD1.n88 VDD1.n69 10.4732
R614 VDD1.n110 VDD1.n59 10.4732
R615 VDD1.n54 VDD1.n0 9.69747
R616 VDD1.n29 VDD1.n28 9.69747
R617 VDD1.n85 VDD1.n84 9.69747
R618 VDD1.n111 VDD1.n57 9.69747
R619 VDD1.n56 VDD1.n55 9.45567
R620 VDD1.n113 VDD1.n112 9.45567
R621 VDD1.n22 VDD1.n21 9.3005
R622 VDD1.n24 VDD1.n23 9.3005
R623 VDD1.n15 VDD1.n14 9.3005
R624 VDD1.n30 VDD1.n29 9.3005
R625 VDD1.n32 VDD1.n31 9.3005
R626 VDD1.n10 VDD1.n9 9.3005
R627 VDD1.n38 VDD1.n37 9.3005
R628 VDD1.n40 VDD1.n39 9.3005
R629 VDD1.n55 VDD1.n54 9.3005
R630 VDD1.n2 VDD1.n1 9.3005
R631 VDD1.n49 VDD1.n48 9.3005
R632 VDD1.n47 VDD1.n46 9.3005
R633 VDD1.n6 VDD1.n5 9.3005
R634 VDD1.n112 VDD1.n111 9.3005
R635 VDD1.n59 VDD1.n58 9.3005
R636 VDD1.n106 VDD1.n105 9.3005
R637 VDD1.n104 VDD1.n103 9.3005
R638 VDD1.n63 VDD1.n62 9.3005
R639 VDD1.n78 VDD1.n77 9.3005
R640 VDD1.n80 VDD1.n79 9.3005
R641 VDD1.n71 VDD1.n70 9.3005
R642 VDD1.n86 VDD1.n85 9.3005
R643 VDD1.n88 VDD1.n87 9.3005
R644 VDD1.n67 VDD1.n66 9.3005
R645 VDD1.n95 VDD1.n94 9.3005
R646 VDD1.n97 VDD1.n96 9.3005
R647 VDD1.n25 VDD1.n15 8.92171
R648 VDD1.n81 VDD1.n71 8.92171
R649 VDD1.n24 VDD1.n17 8.14595
R650 VDD1.n80 VDD1.n73 8.14595
R651 VDD1.n21 VDD1.n20 7.3702
R652 VDD1.n77 VDD1.n76 7.3702
R653 VDD1.n21 VDD1.n17 5.81868
R654 VDD1.n77 VDD1.n73 5.81868
R655 VDD1.n25 VDD1.n24 5.04292
R656 VDD1.n81 VDD1.n80 5.04292
R657 VDD1.n56 VDD1.n0 4.26717
R658 VDD1.n28 VDD1.n15 4.26717
R659 VDD1.n84 VDD1.n71 4.26717
R660 VDD1.n113 VDD1.n57 4.26717
R661 VDD1.n54 VDD1.n53 3.49141
R662 VDD1.n29 VDD1.n13 3.49141
R663 VDD1.n85 VDD1.n69 3.49141
R664 VDD1.n111 VDD1.n110 3.49141
R665 VDD1.n50 VDD1.n2 2.71565
R666 VDD1.n33 VDD1.n32 2.71565
R667 VDD1.n89 VDD1.n88 2.71565
R668 VDD1.n107 VDD1.n59 2.71565
R669 VDD1.n22 VDD1.n18 2.41282
R670 VDD1.n78 VDD1.n74 2.41282
R671 VDD1.n49 VDD1.n4 1.93989
R672 VDD1.n36 VDD1.n10 1.93989
R673 VDD1.n93 VDD1.n67 1.93989
R674 VDD1.n106 VDD1.n61 1.93989
R675 VDD1.n46 VDD1.n45 1.16414
R676 VDD1.n37 VDD1.n8 1.16414
R677 VDD1.n94 VDD1.n65 1.16414
R678 VDD1.n103 VDD1.n102 1.16414
R679 VDD1.n42 VDD1.n6 0.388379
R680 VDD1.n41 VDD1.n40 0.388379
R681 VDD1.n98 VDD1.n97 0.388379
R682 VDD1.n99 VDD1.n63 0.388379
R683 VDD1.n55 VDD1.n1 0.155672
R684 VDD1.n48 VDD1.n1 0.155672
R685 VDD1.n48 VDD1.n47 0.155672
R686 VDD1.n47 VDD1.n5 0.155672
R687 VDD1.n39 VDD1.n5 0.155672
R688 VDD1.n39 VDD1.n38 0.155672
R689 VDD1.n38 VDD1.n9 0.155672
R690 VDD1.n31 VDD1.n9 0.155672
R691 VDD1.n31 VDD1.n30 0.155672
R692 VDD1.n30 VDD1.n14 0.155672
R693 VDD1.n23 VDD1.n14 0.155672
R694 VDD1.n23 VDD1.n22 0.155672
R695 VDD1.n79 VDD1.n78 0.155672
R696 VDD1.n79 VDD1.n70 0.155672
R697 VDD1.n86 VDD1.n70 0.155672
R698 VDD1.n87 VDD1.n86 0.155672
R699 VDD1.n87 VDD1.n66 0.155672
R700 VDD1.n95 VDD1.n66 0.155672
R701 VDD1.n96 VDD1.n95 0.155672
R702 VDD1.n96 VDD1.n62 0.155672
R703 VDD1.n104 VDD1.n62 0.155672
R704 VDD1.n105 VDD1.n104 0.155672
R705 VDD1.n105 VDD1.n58 0.155672
R706 VDD1.n112 VDD1.n58 0.155672
R707 B.n329 B.n56 585
R708 B.n331 B.n330 585
R709 B.n332 B.n55 585
R710 B.n334 B.n333 585
R711 B.n335 B.n54 585
R712 B.n337 B.n336 585
R713 B.n338 B.n53 585
R714 B.n340 B.n339 585
R715 B.n341 B.n52 585
R716 B.n343 B.n342 585
R717 B.n344 B.n51 585
R718 B.n346 B.n345 585
R719 B.n347 B.n50 585
R720 B.n349 B.n348 585
R721 B.n350 B.n49 585
R722 B.n352 B.n351 585
R723 B.n353 B.n48 585
R724 B.n355 B.n354 585
R725 B.n356 B.n47 585
R726 B.n358 B.n357 585
R727 B.n359 B.n46 585
R728 B.n361 B.n360 585
R729 B.n362 B.n45 585
R730 B.n364 B.n363 585
R731 B.n365 B.n44 585
R732 B.n367 B.n366 585
R733 B.n368 B.n43 585
R734 B.n370 B.n369 585
R735 B.n371 B.n42 585
R736 B.n373 B.n372 585
R737 B.n374 B.n41 585
R738 B.n376 B.n375 585
R739 B.n377 B.n40 585
R740 B.n379 B.n378 585
R741 B.n380 B.n39 585
R742 B.n382 B.n381 585
R743 B.n383 B.n38 585
R744 B.n385 B.n384 585
R745 B.n387 B.n35 585
R746 B.n389 B.n388 585
R747 B.n390 B.n34 585
R748 B.n392 B.n391 585
R749 B.n393 B.n33 585
R750 B.n395 B.n394 585
R751 B.n396 B.n32 585
R752 B.n398 B.n397 585
R753 B.n399 B.n29 585
R754 B.n402 B.n401 585
R755 B.n403 B.n28 585
R756 B.n405 B.n404 585
R757 B.n406 B.n27 585
R758 B.n408 B.n407 585
R759 B.n409 B.n26 585
R760 B.n411 B.n410 585
R761 B.n412 B.n25 585
R762 B.n414 B.n413 585
R763 B.n415 B.n24 585
R764 B.n417 B.n416 585
R765 B.n418 B.n23 585
R766 B.n420 B.n419 585
R767 B.n421 B.n22 585
R768 B.n423 B.n422 585
R769 B.n424 B.n21 585
R770 B.n426 B.n425 585
R771 B.n427 B.n20 585
R772 B.n429 B.n428 585
R773 B.n430 B.n19 585
R774 B.n432 B.n431 585
R775 B.n433 B.n18 585
R776 B.n435 B.n434 585
R777 B.n436 B.n17 585
R778 B.n438 B.n437 585
R779 B.n439 B.n16 585
R780 B.n441 B.n440 585
R781 B.n442 B.n15 585
R782 B.n444 B.n443 585
R783 B.n445 B.n14 585
R784 B.n447 B.n446 585
R785 B.n448 B.n13 585
R786 B.n450 B.n449 585
R787 B.n451 B.n12 585
R788 B.n453 B.n452 585
R789 B.n454 B.n11 585
R790 B.n456 B.n455 585
R791 B.n457 B.n10 585
R792 B.n328 B.n327 585
R793 B.n326 B.n57 585
R794 B.n325 B.n324 585
R795 B.n323 B.n58 585
R796 B.n322 B.n321 585
R797 B.n320 B.n59 585
R798 B.n319 B.n318 585
R799 B.n317 B.n60 585
R800 B.n316 B.n315 585
R801 B.n314 B.n61 585
R802 B.n313 B.n312 585
R803 B.n311 B.n62 585
R804 B.n310 B.n309 585
R805 B.n308 B.n63 585
R806 B.n307 B.n306 585
R807 B.n305 B.n64 585
R808 B.n304 B.n303 585
R809 B.n302 B.n65 585
R810 B.n301 B.n300 585
R811 B.n299 B.n66 585
R812 B.n298 B.n297 585
R813 B.n296 B.n67 585
R814 B.n295 B.n294 585
R815 B.n293 B.n68 585
R816 B.n292 B.n291 585
R817 B.n290 B.n69 585
R818 B.n289 B.n288 585
R819 B.n287 B.n70 585
R820 B.n286 B.n285 585
R821 B.n284 B.n71 585
R822 B.n283 B.n282 585
R823 B.n281 B.n72 585
R824 B.n280 B.n279 585
R825 B.n151 B.n150 585
R826 B.n152 B.n119 585
R827 B.n154 B.n153 585
R828 B.n155 B.n118 585
R829 B.n157 B.n156 585
R830 B.n158 B.n117 585
R831 B.n160 B.n159 585
R832 B.n161 B.n116 585
R833 B.n163 B.n162 585
R834 B.n164 B.n115 585
R835 B.n166 B.n165 585
R836 B.n167 B.n114 585
R837 B.n169 B.n168 585
R838 B.n170 B.n113 585
R839 B.n172 B.n171 585
R840 B.n173 B.n112 585
R841 B.n175 B.n174 585
R842 B.n176 B.n111 585
R843 B.n178 B.n177 585
R844 B.n179 B.n110 585
R845 B.n181 B.n180 585
R846 B.n182 B.n109 585
R847 B.n184 B.n183 585
R848 B.n185 B.n108 585
R849 B.n187 B.n186 585
R850 B.n188 B.n107 585
R851 B.n190 B.n189 585
R852 B.n191 B.n106 585
R853 B.n193 B.n192 585
R854 B.n194 B.n105 585
R855 B.n196 B.n195 585
R856 B.n197 B.n104 585
R857 B.n199 B.n198 585
R858 B.n200 B.n103 585
R859 B.n202 B.n201 585
R860 B.n203 B.n102 585
R861 B.n205 B.n204 585
R862 B.n206 B.n99 585
R863 B.n209 B.n208 585
R864 B.n210 B.n98 585
R865 B.n212 B.n211 585
R866 B.n213 B.n97 585
R867 B.n215 B.n214 585
R868 B.n216 B.n96 585
R869 B.n218 B.n217 585
R870 B.n219 B.n95 585
R871 B.n221 B.n220 585
R872 B.n223 B.n222 585
R873 B.n224 B.n91 585
R874 B.n226 B.n225 585
R875 B.n227 B.n90 585
R876 B.n229 B.n228 585
R877 B.n230 B.n89 585
R878 B.n232 B.n231 585
R879 B.n233 B.n88 585
R880 B.n235 B.n234 585
R881 B.n236 B.n87 585
R882 B.n238 B.n237 585
R883 B.n239 B.n86 585
R884 B.n241 B.n240 585
R885 B.n242 B.n85 585
R886 B.n244 B.n243 585
R887 B.n245 B.n84 585
R888 B.n247 B.n246 585
R889 B.n248 B.n83 585
R890 B.n250 B.n249 585
R891 B.n251 B.n82 585
R892 B.n253 B.n252 585
R893 B.n254 B.n81 585
R894 B.n256 B.n255 585
R895 B.n257 B.n80 585
R896 B.n259 B.n258 585
R897 B.n260 B.n79 585
R898 B.n262 B.n261 585
R899 B.n263 B.n78 585
R900 B.n265 B.n264 585
R901 B.n266 B.n77 585
R902 B.n268 B.n267 585
R903 B.n269 B.n76 585
R904 B.n271 B.n270 585
R905 B.n272 B.n75 585
R906 B.n274 B.n273 585
R907 B.n275 B.n74 585
R908 B.n277 B.n276 585
R909 B.n278 B.n73 585
R910 B.n149 B.n120 585
R911 B.n148 B.n147 585
R912 B.n146 B.n121 585
R913 B.n145 B.n144 585
R914 B.n143 B.n122 585
R915 B.n142 B.n141 585
R916 B.n140 B.n123 585
R917 B.n139 B.n138 585
R918 B.n137 B.n124 585
R919 B.n136 B.n135 585
R920 B.n134 B.n125 585
R921 B.n133 B.n132 585
R922 B.n131 B.n126 585
R923 B.n130 B.n129 585
R924 B.n128 B.n127 585
R925 B.n2 B.n0 585
R926 B.n481 B.n1 585
R927 B.n480 B.n479 585
R928 B.n478 B.n3 585
R929 B.n477 B.n476 585
R930 B.n475 B.n4 585
R931 B.n474 B.n473 585
R932 B.n472 B.n5 585
R933 B.n471 B.n470 585
R934 B.n469 B.n6 585
R935 B.n468 B.n467 585
R936 B.n466 B.n7 585
R937 B.n465 B.n464 585
R938 B.n463 B.n8 585
R939 B.n462 B.n461 585
R940 B.n460 B.n9 585
R941 B.n459 B.n458 585
R942 B.n483 B.n482 585
R943 B.n150 B.n149 482.89
R944 B.n458 B.n457 482.89
R945 B.n280 B.n73 482.89
R946 B.n329 B.n328 482.89
R947 B.n92 B.t9 450.678
R948 B.n100 B.t6 450.678
R949 B.n30 B.t0 450.678
R950 B.n36 B.t3 450.678
R951 B.n92 B.t11 376.252
R952 B.n36 B.t4 376.252
R953 B.n100 B.t8 376.252
R954 B.n30 B.t1 376.252
R955 B.n93 B.t10 349.877
R956 B.n37 B.t5 349.877
R957 B.n101 B.t7 349.877
R958 B.n31 B.t2 349.877
R959 B.n149 B.n148 163.367
R960 B.n148 B.n121 163.367
R961 B.n144 B.n121 163.367
R962 B.n144 B.n143 163.367
R963 B.n143 B.n142 163.367
R964 B.n142 B.n123 163.367
R965 B.n138 B.n123 163.367
R966 B.n138 B.n137 163.367
R967 B.n137 B.n136 163.367
R968 B.n136 B.n125 163.367
R969 B.n132 B.n125 163.367
R970 B.n132 B.n131 163.367
R971 B.n131 B.n130 163.367
R972 B.n130 B.n127 163.367
R973 B.n127 B.n2 163.367
R974 B.n482 B.n2 163.367
R975 B.n482 B.n481 163.367
R976 B.n481 B.n480 163.367
R977 B.n480 B.n3 163.367
R978 B.n476 B.n3 163.367
R979 B.n476 B.n475 163.367
R980 B.n475 B.n474 163.367
R981 B.n474 B.n5 163.367
R982 B.n470 B.n5 163.367
R983 B.n470 B.n469 163.367
R984 B.n469 B.n468 163.367
R985 B.n468 B.n7 163.367
R986 B.n464 B.n7 163.367
R987 B.n464 B.n463 163.367
R988 B.n463 B.n462 163.367
R989 B.n462 B.n9 163.367
R990 B.n458 B.n9 163.367
R991 B.n150 B.n119 163.367
R992 B.n154 B.n119 163.367
R993 B.n155 B.n154 163.367
R994 B.n156 B.n155 163.367
R995 B.n156 B.n117 163.367
R996 B.n160 B.n117 163.367
R997 B.n161 B.n160 163.367
R998 B.n162 B.n161 163.367
R999 B.n162 B.n115 163.367
R1000 B.n166 B.n115 163.367
R1001 B.n167 B.n166 163.367
R1002 B.n168 B.n167 163.367
R1003 B.n168 B.n113 163.367
R1004 B.n172 B.n113 163.367
R1005 B.n173 B.n172 163.367
R1006 B.n174 B.n173 163.367
R1007 B.n174 B.n111 163.367
R1008 B.n178 B.n111 163.367
R1009 B.n179 B.n178 163.367
R1010 B.n180 B.n179 163.367
R1011 B.n180 B.n109 163.367
R1012 B.n184 B.n109 163.367
R1013 B.n185 B.n184 163.367
R1014 B.n186 B.n185 163.367
R1015 B.n186 B.n107 163.367
R1016 B.n190 B.n107 163.367
R1017 B.n191 B.n190 163.367
R1018 B.n192 B.n191 163.367
R1019 B.n192 B.n105 163.367
R1020 B.n196 B.n105 163.367
R1021 B.n197 B.n196 163.367
R1022 B.n198 B.n197 163.367
R1023 B.n198 B.n103 163.367
R1024 B.n202 B.n103 163.367
R1025 B.n203 B.n202 163.367
R1026 B.n204 B.n203 163.367
R1027 B.n204 B.n99 163.367
R1028 B.n209 B.n99 163.367
R1029 B.n210 B.n209 163.367
R1030 B.n211 B.n210 163.367
R1031 B.n211 B.n97 163.367
R1032 B.n215 B.n97 163.367
R1033 B.n216 B.n215 163.367
R1034 B.n217 B.n216 163.367
R1035 B.n217 B.n95 163.367
R1036 B.n221 B.n95 163.367
R1037 B.n222 B.n221 163.367
R1038 B.n222 B.n91 163.367
R1039 B.n226 B.n91 163.367
R1040 B.n227 B.n226 163.367
R1041 B.n228 B.n227 163.367
R1042 B.n228 B.n89 163.367
R1043 B.n232 B.n89 163.367
R1044 B.n233 B.n232 163.367
R1045 B.n234 B.n233 163.367
R1046 B.n234 B.n87 163.367
R1047 B.n238 B.n87 163.367
R1048 B.n239 B.n238 163.367
R1049 B.n240 B.n239 163.367
R1050 B.n240 B.n85 163.367
R1051 B.n244 B.n85 163.367
R1052 B.n245 B.n244 163.367
R1053 B.n246 B.n245 163.367
R1054 B.n246 B.n83 163.367
R1055 B.n250 B.n83 163.367
R1056 B.n251 B.n250 163.367
R1057 B.n252 B.n251 163.367
R1058 B.n252 B.n81 163.367
R1059 B.n256 B.n81 163.367
R1060 B.n257 B.n256 163.367
R1061 B.n258 B.n257 163.367
R1062 B.n258 B.n79 163.367
R1063 B.n262 B.n79 163.367
R1064 B.n263 B.n262 163.367
R1065 B.n264 B.n263 163.367
R1066 B.n264 B.n77 163.367
R1067 B.n268 B.n77 163.367
R1068 B.n269 B.n268 163.367
R1069 B.n270 B.n269 163.367
R1070 B.n270 B.n75 163.367
R1071 B.n274 B.n75 163.367
R1072 B.n275 B.n274 163.367
R1073 B.n276 B.n275 163.367
R1074 B.n276 B.n73 163.367
R1075 B.n281 B.n280 163.367
R1076 B.n282 B.n281 163.367
R1077 B.n282 B.n71 163.367
R1078 B.n286 B.n71 163.367
R1079 B.n287 B.n286 163.367
R1080 B.n288 B.n287 163.367
R1081 B.n288 B.n69 163.367
R1082 B.n292 B.n69 163.367
R1083 B.n293 B.n292 163.367
R1084 B.n294 B.n293 163.367
R1085 B.n294 B.n67 163.367
R1086 B.n298 B.n67 163.367
R1087 B.n299 B.n298 163.367
R1088 B.n300 B.n299 163.367
R1089 B.n300 B.n65 163.367
R1090 B.n304 B.n65 163.367
R1091 B.n305 B.n304 163.367
R1092 B.n306 B.n305 163.367
R1093 B.n306 B.n63 163.367
R1094 B.n310 B.n63 163.367
R1095 B.n311 B.n310 163.367
R1096 B.n312 B.n311 163.367
R1097 B.n312 B.n61 163.367
R1098 B.n316 B.n61 163.367
R1099 B.n317 B.n316 163.367
R1100 B.n318 B.n317 163.367
R1101 B.n318 B.n59 163.367
R1102 B.n322 B.n59 163.367
R1103 B.n323 B.n322 163.367
R1104 B.n324 B.n323 163.367
R1105 B.n324 B.n57 163.367
R1106 B.n328 B.n57 163.367
R1107 B.n457 B.n456 163.367
R1108 B.n456 B.n11 163.367
R1109 B.n452 B.n11 163.367
R1110 B.n452 B.n451 163.367
R1111 B.n451 B.n450 163.367
R1112 B.n450 B.n13 163.367
R1113 B.n446 B.n13 163.367
R1114 B.n446 B.n445 163.367
R1115 B.n445 B.n444 163.367
R1116 B.n444 B.n15 163.367
R1117 B.n440 B.n15 163.367
R1118 B.n440 B.n439 163.367
R1119 B.n439 B.n438 163.367
R1120 B.n438 B.n17 163.367
R1121 B.n434 B.n17 163.367
R1122 B.n434 B.n433 163.367
R1123 B.n433 B.n432 163.367
R1124 B.n432 B.n19 163.367
R1125 B.n428 B.n19 163.367
R1126 B.n428 B.n427 163.367
R1127 B.n427 B.n426 163.367
R1128 B.n426 B.n21 163.367
R1129 B.n422 B.n21 163.367
R1130 B.n422 B.n421 163.367
R1131 B.n421 B.n420 163.367
R1132 B.n420 B.n23 163.367
R1133 B.n416 B.n23 163.367
R1134 B.n416 B.n415 163.367
R1135 B.n415 B.n414 163.367
R1136 B.n414 B.n25 163.367
R1137 B.n410 B.n25 163.367
R1138 B.n410 B.n409 163.367
R1139 B.n409 B.n408 163.367
R1140 B.n408 B.n27 163.367
R1141 B.n404 B.n27 163.367
R1142 B.n404 B.n403 163.367
R1143 B.n403 B.n402 163.367
R1144 B.n402 B.n29 163.367
R1145 B.n397 B.n29 163.367
R1146 B.n397 B.n396 163.367
R1147 B.n396 B.n395 163.367
R1148 B.n395 B.n33 163.367
R1149 B.n391 B.n33 163.367
R1150 B.n391 B.n390 163.367
R1151 B.n390 B.n389 163.367
R1152 B.n389 B.n35 163.367
R1153 B.n384 B.n35 163.367
R1154 B.n384 B.n383 163.367
R1155 B.n383 B.n382 163.367
R1156 B.n382 B.n39 163.367
R1157 B.n378 B.n39 163.367
R1158 B.n378 B.n377 163.367
R1159 B.n377 B.n376 163.367
R1160 B.n376 B.n41 163.367
R1161 B.n372 B.n41 163.367
R1162 B.n372 B.n371 163.367
R1163 B.n371 B.n370 163.367
R1164 B.n370 B.n43 163.367
R1165 B.n366 B.n43 163.367
R1166 B.n366 B.n365 163.367
R1167 B.n365 B.n364 163.367
R1168 B.n364 B.n45 163.367
R1169 B.n360 B.n45 163.367
R1170 B.n360 B.n359 163.367
R1171 B.n359 B.n358 163.367
R1172 B.n358 B.n47 163.367
R1173 B.n354 B.n47 163.367
R1174 B.n354 B.n353 163.367
R1175 B.n353 B.n352 163.367
R1176 B.n352 B.n49 163.367
R1177 B.n348 B.n49 163.367
R1178 B.n348 B.n347 163.367
R1179 B.n347 B.n346 163.367
R1180 B.n346 B.n51 163.367
R1181 B.n342 B.n51 163.367
R1182 B.n342 B.n341 163.367
R1183 B.n341 B.n340 163.367
R1184 B.n340 B.n53 163.367
R1185 B.n336 B.n53 163.367
R1186 B.n336 B.n335 163.367
R1187 B.n335 B.n334 163.367
R1188 B.n334 B.n55 163.367
R1189 B.n330 B.n55 163.367
R1190 B.n330 B.n329 163.367
R1191 B.n94 B.n93 59.5399
R1192 B.n207 B.n101 59.5399
R1193 B.n400 B.n31 59.5399
R1194 B.n386 B.n37 59.5399
R1195 B.n459 B.n10 31.3761
R1196 B.n327 B.n56 31.3761
R1197 B.n279 B.n278 31.3761
R1198 B.n151 B.n120 31.3761
R1199 B.n93 B.n92 26.3763
R1200 B.n101 B.n100 26.3763
R1201 B.n31 B.n30 26.3763
R1202 B.n37 B.n36 26.3763
R1203 B B.n483 18.0485
R1204 B.n455 B.n10 10.6151
R1205 B.n455 B.n454 10.6151
R1206 B.n454 B.n453 10.6151
R1207 B.n453 B.n12 10.6151
R1208 B.n449 B.n12 10.6151
R1209 B.n449 B.n448 10.6151
R1210 B.n448 B.n447 10.6151
R1211 B.n447 B.n14 10.6151
R1212 B.n443 B.n14 10.6151
R1213 B.n443 B.n442 10.6151
R1214 B.n442 B.n441 10.6151
R1215 B.n441 B.n16 10.6151
R1216 B.n437 B.n16 10.6151
R1217 B.n437 B.n436 10.6151
R1218 B.n436 B.n435 10.6151
R1219 B.n435 B.n18 10.6151
R1220 B.n431 B.n18 10.6151
R1221 B.n431 B.n430 10.6151
R1222 B.n430 B.n429 10.6151
R1223 B.n429 B.n20 10.6151
R1224 B.n425 B.n20 10.6151
R1225 B.n425 B.n424 10.6151
R1226 B.n424 B.n423 10.6151
R1227 B.n423 B.n22 10.6151
R1228 B.n419 B.n22 10.6151
R1229 B.n419 B.n418 10.6151
R1230 B.n418 B.n417 10.6151
R1231 B.n417 B.n24 10.6151
R1232 B.n413 B.n24 10.6151
R1233 B.n413 B.n412 10.6151
R1234 B.n412 B.n411 10.6151
R1235 B.n411 B.n26 10.6151
R1236 B.n407 B.n26 10.6151
R1237 B.n407 B.n406 10.6151
R1238 B.n406 B.n405 10.6151
R1239 B.n405 B.n28 10.6151
R1240 B.n401 B.n28 10.6151
R1241 B.n399 B.n398 10.6151
R1242 B.n398 B.n32 10.6151
R1243 B.n394 B.n32 10.6151
R1244 B.n394 B.n393 10.6151
R1245 B.n393 B.n392 10.6151
R1246 B.n392 B.n34 10.6151
R1247 B.n388 B.n34 10.6151
R1248 B.n388 B.n387 10.6151
R1249 B.n385 B.n38 10.6151
R1250 B.n381 B.n38 10.6151
R1251 B.n381 B.n380 10.6151
R1252 B.n380 B.n379 10.6151
R1253 B.n379 B.n40 10.6151
R1254 B.n375 B.n40 10.6151
R1255 B.n375 B.n374 10.6151
R1256 B.n374 B.n373 10.6151
R1257 B.n373 B.n42 10.6151
R1258 B.n369 B.n42 10.6151
R1259 B.n369 B.n368 10.6151
R1260 B.n368 B.n367 10.6151
R1261 B.n367 B.n44 10.6151
R1262 B.n363 B.n44 10.6151
R1263 B.n363 B.n362 10.6151
R1264 B.n362 B.n361 10.6151
R1265 B.n361 B.n46 10.6151
R1266 B.n357 B.n46 10.6151
R1267 B.n357 B.n356 10.6151
R1268 B.n356 B.n355 10.6151
R1269 B.n355 B.n48 10.6151
R1270 B.n351 B.n48 10.6151
R1271 B.n351 B.n350 10.6151
R1272 B.n350 B.n349 10.6151
R1273 B.n349 B.n50 10.6151
R1274 B.n345 B.n50 10.6151
R1275 B.n345 B.n344 10.6151
R1276 B.n344 B.n343 10.6151
R1277 B.n343 B.n52 10.6151
R1278 B.n339 B.n52 10.6151
R1279 B.n339 B.n338 10.6151
R1280 B.n338 B.n337 10.6151
R1281 B.n337 B.n54 10.6151
R1282 B.n333 B.n54 10.6151
R1283 B.n333 B.n332 10.6151
R1284 B.n332 B.n331 10.6151
R1285 B.n331 B.n56 10.6151
R1286 B.n279 B.n72 10.6151
R1287 B.n283 B.n72 10.6151
R1288 B.n284 B.n283 10.6151
R1289 B.n285 B.n284 10.6151
R1290 B.n285 B.n70 10.6151
R1291 B.n289 B.n70 10.6151
R1292 B.n290 B.n289 10.6151
R1293 B.n291 B.n290 10.6151
R1294 B.n291 B.n68 10.6151
R1295 B.n295 B.n68 10.6151
R1296 B.n296 B.n295 10.6151
R1297 B.n297 B.n296 10.6151
R1298 B.n297 B.n66 10.6151
R1299 B.n301 B.n66 10.6151
R1300 B.n302 B.n301 10.6151
R1301 B.n303 B.n302 10.6151
R1302 B.n303 B.n64 10.6151
R1303 B.n307 B.n64 10.6151
R1304 B.n308 B.n307 10.6151
R1305 B.n309 B.n308 10.6151
R1306 B.n309 B.n62 10.6151
R1307 B.n313 B.n62 10.6151
R1308 B.n314 B.n313 10.6151
R1309 B.n315 B.n314 10.6151
R1310 B.n315 B.n60 10.6151
R1311 B.n319 B.n60 10.6151
R1312 B.n320 B.n319 10.6151
R1313 B.n321 B.n320 10.6151
R1314 B.n321 B.n58 10.6151
R1315 B.n325 B.n58 10.6151
R1316 B.n326 B.n325 10.6151
R1317 B.n327 B.n326 10.6151
R1318 B.n152 B.n151 10.6151
R1319 B.n153 B.n152 10.6151
R1320 B.n153 B.n118 10.6151
R1321 B.n157 B.n118 10.6151
R1322 B.n158 B.n157 10.6151
R1323 B.n159 B.n158 10.6151
R1324 B.n159 B.n116 10.6151
R1325 B.n163 B.n116 10.6151
R1326 B.n164 B.n163 10.6151
R1327 B.n165 B.n164 10.6151
R1328 B.n165 B.n114 10.6151
R1329 B.n169 B.n114 10.6151
R1330 B.n170 B.n169 10.6151
R1331 B.n171 B.n170 10.6151
R1332 B.n171 B.n112 10.6151
R1333 B.n175 B.n112 10.6151
R1334 B.n176 B.n175 10.6151
R1335 B.n177 B.n176 10.6151
R1336 B.n177 B.n110 10.6151
R1337 B.n181 B.n110 10.6151
R1338 B.n182 B.n181 10.6151
R1339 B.n183 B.n182 10.6151
R1340 B.n183 B.n108 10.6151
R1341 B.n187 B.n108 10.6151
R1342 B.n188 B.n187 10.6151
R1343 B.n189 B.n188 10.6151
R1344 B.n189 B.n106 10.6151
R1345 B.n193 B.n106 10.6151
R1346 B.n194 B.n193 10.6151
R1347 B.n195 B.n194 10.6151
R1348 B.n195 B.n104 10.6151
R1349 B.n199 B.n104 10.6151
R1350 B.n200 B.n199 10.6151
R1351 B.n201 B.n200 10.6151
R1352 B.n201 B.n102 10.6151
R1353 B.n205 B.n102 10.6151
R1354 B.n206 B.n205 10.6151
R1355 B.n208 B.n98 10.6151
R1356 B.n212 B.n98 10.6151
R1357 B.n213 B.n212 10.6151
R1358 B.n214 B.n213 10.6151
R1359 B.n214 B.n96 10.6151
R1360 B.n218 B.n96 10.6151
R1361 B.n219 B.n218 10.6151
R1362 B.n220 B.n219 10.6151
R1363 B.n224 B.n223 10.6151
R1364 B.n225 B.n224 10.6151
R1365 B.n225 B.n90 10.6151
R1366 B.n229 B.n90 10.6151
R1367 B.n230 B.n229 10.6151
R1368 B.n231 B.n230 10.6151
R1369 B.n231 B.n88 10.6151
R1370 B.n235 B.n88 10.6151
R1371 B.n236 B.n235 10.6151
R1372 B.n237 B.n236 10.6151
R1373 B.n237 B.n86 10.6151
R1374 B.n241 B.n86 10.6151
R1375 B.n242 B.n241 10.6151
R1376 B.n243 B.n242 10.6151
R1377 B.n243 B.n84 10.6151
R1378 B.n247 B.n84 10.6151
R1379 B.n248 B.n247 10.6151
R1380 B.n249 B.n248 10.6151
R1381 B.n249 B.n82 10.6151
R1382 B.n253 B.n82 10.6151
R1383 B.n254 B.n253 10.6151
R1384 B.n255 B.n254 10.6151
R1385 B.n255 B.n80 10.6151
R1386 B.n259 B.n80 10.6151
R1387 B.n260 B.n259 10.6151
R1388 B.n261 B.n260 10.6151
R1389 B.n261 B.n78 10.6151
R1390 B.n265 B.n78 10.6151
R1391 B.n266 B.n265 10.6151
R1392 B.n267 B.n266 10.6151
R1393 B.n267 B.n76 10.6151
R1394 B.n271 B.n76 10.6151
R1395 B.n272 B.n271 10.6151
R1396 B.n273 B.n272 10.6151
R1397 B.n273 B.n74 10.6151
R1398 B.n277 B.n74 10.6151
R1399 B.n278 B.n277 10.6151
R1400 B.n147 B.n120 10.6151
R1401 B.n147 B.n146 10.6151
R1402 B.n146 B.n145 10.6151
R1403 B.n145 B.n122 10.6151
R1404 B.n141 B.n122 10.6151
R1405 B.n141 B.n140 10.6151
R1406 B.n140 B.n139 10.6151
R1407 B.n139 B.n124 10.6151
R1408 B.n135 B.n124 10.6151
R1409 B.n135 B.n134 10.6151
R1410 B.n134 B.n133 10.6151
R1411 B.n133 B.n126 10.6151
R1412 B.n129 B.n126 10.6151
R1413 B.n129 B.n128 10.6151
R1414 B.n128 B.n0 10.6151
R1415 B.n479 B.n1 10.6151
R1416 B.n479 B.n478 10.6151
R1417 B.n478 B.n477 10.6151
R1418 B.n477 B.n4 10.6151
R1419 B.n473 B.n4 10.6151
R1420 B.n473 B.n472 10.6151
R1421 B.n472 B.n471 10.6151
R1422 B.n471 B.n6 10.6151
R1423 B.n467 B.n6 10.6151
R1424 B.n467 B.n466 10.6151
R1425 B.n466 B.n465 10.6151
R1426 B.n465 B.n8 10.6151
R1427 B.n461 B.n8 10.6151
R1428 B.n461 B.n460 10.6151
R1429 B.n460 B.n459 10.6151
R1430 B.n400 B.n399 7.18099
R1431 B.n387 B.n386 7.18099
R1432 B.n208 B.n207 7.18099
R1433 B.n220 B.n94 7.18099
R1434 B.n401 B.n400 3.43465
R1435 B.n386 B.n385 3.43465
R1436 B.n207 B.n206 3.43465
R1437 B.n223 B.n94 3.43465
R1438 B.n483 B.n0 2.81026
R1439 B.n483 B.n1 2.81026
C0 VP B 1.07514f
C1 VTAIL VP 1.63487f
C2 VN B 0.769941f
C3 VTAIL VN 1.6204f
C4 VP VDD2 0.268864f
C5 VTAIL B 2.63241f
C6 VN VDD2 2.01687f
C7 VDD1 VP 2.13324f
C8 B VDD2 1.38447f
C9 VTAIL VDD2 4.85101f
C10 VDD1 VN 0.149073f
C11 VDD1 B 1.3676f
C12 VDD1 VTAIL 4.81314f
C13 VP w_n1514_n3088# 2.10864f
C14 VN w_n1514_n3088# 1.91917f
C15 VDD1 VDD2 0.494896f
C16 w_n1514_n3088# B 6.7191f
C17 VTAIL w_n1514_n3088# 2.63988f
C18 w_n1514_n3088# VDD2 1.51214f
C19 VN VP 4.44558f
C20 VDD1 w_n1514_n3088# 1.50417f
C21 VDD2 VSUBS 0.724074f
C22 VDD1 VSUBS 3.03925f
C23 VTAIL VSUBS 0.744007f
C24 VN VSUBS 5.1964f
C25 VP VSUBS 1.153098f
C26 B VSUBS 2.618409f
C27 w_n1514_n3088# VSUBS 57.6834f
C28 B.n0 VSUBS 0.004591f
C29 B.n1 VSUBS 0.004591f
C30 B.n2 VSUBS 0.00726f
C31 B.n3 VSUBS 0.00726f
C32 B.n4 VSUBS 0.00726f
C33 B.n5 VSUBS 0.00726f
C34 B.n6 VSUBS 0.00726f
C35 B.n7 VSUBS 0.00726f
C36 B.n8 VSUBS 0.00726f
C37 B.n9 VSUBS 0.00726f
C38 B.n10 VSUBS 0.017213f
C39 B.n11 VSUBS 0.00726f
C40 B.n12 VSUBS 0.00726f
C41 B.n13 VSUBS 0.00726f
C42 B.n14 VSUBS 0.00726f
C43 B.n15 VSUBS 0.00726f
C44 B.n16 VSUBS 0.00726f
C45 B.n17 VSUBS 0.00726f
C46 B.n18 VSUBS 0.00726f
C47 B.n19 VSUBS 0.00726f
C48 B.n20 VSUBS 0.00726f
C49 B.n21 VSUBS 0.00726f
C50 B.n22 VSUBS 0.00726f
C51 B.n23 VSUBS 0.00726f
C52 B.n24 VSUBS 0.00726f
C53 B.n25 VSUBS 0.00726f
C54 B.n26 VSUBS 0.00726f
C55 B.n27 VSUBS 0.00726f
C56 B.n28 VSUBS 0.00726f
C57 B.n29 VSUBS 0.00726f
C58 B.t2 VSUBS 0.186388f
C59 B.t1 VSUBS 0.202043f
C60 B.t0 VSUBS 0.484089f
C61 B.n30 VSUBS 0.308495f
C62 B.n31 VSUBS 0.233681f
C63 B.n32 VSUBS 0.00726f
C64 B.n33 VSUBS 0.00726f
C65 B.n34 VSUBS 0.00726f
C66 B.n35 VSUBS 0.00726f
C67 B.t5 VSUBS 0.186391f
C68 B.t4 VSUBS 0.202046f
C69 B.t3 VSUBS 0.484089f
C70 B.n36 VSUBS 0.308493f
C71 B.n37 VSUBS 0.233678f
C72 B.n38 VSUBS 0.00726f
C73 B.n39 VSUBS 0.00726f
C74 B.n40 VSUBS 0.00726f
C75 B.n41 VSUBS 0.00726f
C76 B.n42 VSUBS 0.00726f
C77 B.n43 VSUBS 0.00726f
C78 B.n44 VSUBS 0.00726f
C79 B.n45 VSUBS 0.00726f
C80 B.n46 VSUBS 0.00726f
C81 B.n47 VSUBS 0.00726f
C82 B.n48 VSUBS 0.00726f
C83 B.n49 VSUBS 0.00726f
C84 B.n50 VSUBS 0.00726f
C85 B.n51 VSUBS 0.00726f
C86 B.n52 VSUBS 0.00726f
C87 B.n53 VSUBS 0.00726f
C88 B.n54 VSUBS 0.00726f
C89 B.n55 VSUBS 0.00726f
C90 B.n56 VSUBS 0.01632f
C91 B.n57 VSUBS 0.00726f
C92 B.n58 VSUBS 0.00726f
C93 B.n59 VSUBS 0.00726f
C94 B.n60 VSUBS 0.00726f
C95 B.n61 VSUBS 0.00726f
C96 B.n62 VSUBS 0.00726f
C97 B.n63 VSUBS 0.00726f
C98 B.n64 VSUBS 0.00726f
C99 B.n65 VSUBS 0.00726f
C100 B.n66 VSUBS 0.00726f
C101 B.n67 VSUBS 0.00726f
C102 B.n68 VSUBS 0.00726f
C103 B.n69 VSUBS 0.00726f
C104 B.n70 VSUBS 0.00726f
C105 B.n71 VSUBS 0.00726f
C106 B.n72 VSUBS 0.00726f
C107 B.n73 VSUBS 0.017213f
C108 B.n74 VSUBS 0.00726f
C109 B.n75 VSUBS 0.00726f
C110 B.n76 VSUBS 0.00726f
C111 B.n77 VSUBS 0.00726f
C112 B.n78 VSUBS 0.00726f
C113 B.n79 VSUBS 0.00726f
C114 B.n80 VSUBS 0.00726f
C115 B.n81 VSUBS 0.00726f
C116 B.n82 VSUBS 0.00726f
C117 B.n83 VSUBS 0.00726f
C118 B.n84 VSUBS 0.00726f
C119 B.n85 VSUBS 0.00726f
C120 B.n86 VSUBS 0.00726f
C121 B.n87 VSUBS 0.00726f
C122 B.n88 VSUBS 0.00726f
C123 B.n89 VSUBS 0.00726f
C124 B.n90 VSUBS 0.00726f
C125 B.n91 VSUBS 0.00726f
C126 B.t10 VSUBS 0.186391f
C127 B.t11 VSUBS 0.202046f
C128 B.t9 VSUBS 0.484089f
C129 B.n92 VSUBS 0.308493f
C130 B.n93 VSUBS 0.233678f
C131 B.n94 VSUBS 0.016821f
C132 B.n95 VSUBS 0.00726f
C133 B.n96 VSUBS 0.00726f
C134 B.n97 VSUBS 0.00726f
C135 B.n98 VSUBS 0.00726f
C136 B.n99 VSUBS 0.00726f
C137 B.t7 VSUBS 0.186388f
C138 B.t8 VSUBS 0.202043f
C139 B.t6 VSUBS 0.484089f
C140 B.n100 VSUBS 0.308495f
C141 B.n101 VSUBS 0.233681f
C142 B.n102 VSUBS 0.00726f
C143 B.n103 VSUBS 0.00726f
C144 B.n104 VSUBS 0.00726f
C145 B.n105 VSUBS 0.00726f
C146 B.n106 VSUBS 0.00726f
C147 B.n107 VSUBS 0.00726f
C148 B.n108 VSUBS 0.00726f
C149 B.n109 VSUBS 0.00726f
C150 B.n110 VSUBS 0.00726f
C151 B.n111 VSUBS 0.00726f
C152 B.n112 VSUBS 0.00726f
C153 B.n113 VSUBS 0.00726f
C154 B.n114 VSUBS 0.00726f
C155 B.n115 VSUBS 0.00726f
C156 B.n116 VSUBS 0.00726f
C157 B.n117 VSUBS 0.00726f
C158 B.n118 VSUBS 0.00726f
C159 B.n119 VSUBS 0.00726f
C160 B.n120 VSUBS 0.015885f
C161 B.n121 VSUBS 0.00726f
C162 B.n122 VSUBS 0.00726f
C163 B.n123 VSUBS 0.00726f
C164 B.n124 VSUBS 0.00726f
C165 B.n125 VSUBS 0.00726f
C166 B.n126 VSUBS 0.00726f
C167 B.n127 VSUBS 0.00726f
C168 B.n128 VSUBS 0.00726f
C169 B.n129 VSUBS 0.00726f
C170 B.n130 VSUBS 0.00726f
C171 B.n131 VSUBS 0.00726f
C172 B.n132 VSUBS 0.00726f
C173 B.n133 VSUBS 0.00726f
C174 B.n134 VSUBS 0.00726f
C175 B.n135 VSUBS 0.00726f
C176 B.n136 VSUBS 0.00726f
C177 B.n137 VSUBS 0.00726f
C178 B.n138 VSUBS 0.00726f
C179 B.n139 VSUBS 0.00726f
C180 B.n140 VSUBS 0.00726f
C181 B.n141 VSUBS 0.00726f
C182 B.n142 VSUBS 0.00726f
C183 B.n143 VSUBS 0.00726f
C184 B.n144 VSUBS 0.00726f
C185 B.n145 VSUBS 0.00726f
C186 B.n146 VSUBS 0.00726f
C187 B.n147 VSUBS 0.00726f
C188 B.n148 VSUBS 0.00726f
C189 B.n149 VSUBS 0.015885f
C190 B.n150 VSUBS 0.017213f
C191 B.n151 VSUBS 0.017213f
C192 B.n152 VSUBS 0.00726f
C193 B.n153 VSUBS 0.00726f
C194 B.n154 VSUBS 0.00726f
C195 B.n155 VSUBS 0.00726f
C196 B.n156 VSUBS 0.00726f
C197 B.n157 VSUBS 0.00726f
C198 B.n158 VSUBS 0.00726f
C199 B.n159 VSUBS 0.00726f
C200 B.n160 VSUBS 0.00726f
C201 B.n161 VSUBS 0.00726f
C202 B.n162 VSUBS 0.00726f
C203 B.n163 VSUBS 0.00726f
C204 B.n164 VSUBS 0.00726f
C205 B.n165 VSUBS 0.00726f
C206 B.n166 VSUBS 0.00726f
C207 B.n167 VSUBS 0.00726f
C208 B.n168 VSUBS 0.00726f
C209 B.n169 VSUBS 0.00726f
C210 B.n170 VSUBS 0.00726f
C211 B.n171 VSUBS 0.00726f
C212 B.n172 VSUBS 0.00726f
C213 B.n173 VSUBS 0.00726f
C214 B.n174 VSUBS 0.00726f
C215 B.n175 VSUBS 0.00726f
C216 B.n176 VSUBS 0.00726f
C217 B.n177 VSUBS 0.00726f
C218 B.n178 VSUBS 0.00726f
C219 B.n179 VSUBS 0.00726f
C220 B.n180 VSUBS 0.00726f
C221 B.n181 VSUBS 0.00726f
C222 B.n182 VSUBS 0.00726f
C223 B.n183 VSUBS 0.00726f
C224 B.n184 VSUBS 0.00726f
C225 B.n185 VSUBS 0.00726f
C226 B.n186 VSUBS 0.00726f
C227 B.n187 VSUBS 0.00726f
C228 B.n188 VSUBS 0.00726f
C229 B.n189 VSUBS 0.00726f
C230 B.n190 VSUBS 0.00726f
C231 B.n191 VSUBS 0.00726f
C232 B.n192 VSUBS 0.00726f
C233 B.n193 VSUBS 0.00726f
C234 B.n194 VSUBS 0.00726f
C235 B.n195 VSUBS 0.00726f
C236 B.n196 VSUBS 0.00726f
C237 B.n197 VSUBS 0.00726f
C238 B.n198 VSUBS 0.00726f
C239 B.n199 VSUBS 0.00726f
C240 B.n200 VSUBS 0.00726f
C241 B.n201 VSUBS 0.00726f
C242 B.n202 VSUBS 0.00726f
C243 B.n203 VSUBS 0.00726f
C244 B.n204 VSUBS 0.00726f
C245 B.n205 VSUBS 0.00726f
C246 B.n206 VSUBS 0.004805f
C247 B.n207 VSUBS 0.016821f
C248 B.n208 VSUBS 0.006086f
C249 B.n209 VSUBS 0.00726f
C250 B.n210 VSUBS 0.00726f
C251 B.n211 VSUBS 0.00726f
C252 B.n212 VSUBS 0.00726f
C253 B.n213 VSUBS 0.00726f
C254 B.n214 VSUBS 0.00726f
C255 B.n215 VSUBS 0.00726f
C256 B.n216 VSUBS 0.00726f
C257 B.n217 VSUBS 0.00726f
C258 B.n218 VSUBS 0.00726f
C259 B.n219 VSUBS 0.00726f
C260 B.n220 VSUBS 0.006086f
C261 B.n221 VSUBS 0.00726f
C262 B.n222 VSUBS 0.00726f
C263 B.n223 VSUBS 0.004805f
C264 B.n224 VSUBS 0.00726f
C265 B.n225 VSUBS 0.00726f
C266 B.n226 VSUBS 0.00726f
C267 B.n227 VSUBS 0.00726f
C268 B.n228 VSUBS 0.00726f
C269 B.n229 VSUBS 0.00726f
C270 B.n230 VSUBS 0.00726f
C271 B.n231 VSUBS 0.00726f
C272 B.n232 VSUBS 0.00726f
C273 B.n233 VSUBS 0.00726f
C274 B.n234 VSUBS 0.00726f
C275 B.n235 VSUBS 0.00726f
C276 B.n236 VSUBS 0.00726f
C277 B.n237 VSUBS 0.00726f
C278 B.n238 VSUBS 0.00726f
C279 B.n239 VSUBS 0.00726f
C280 B.n240 VSUBS 0.00726f
C281 B.n241 VSUBS 0.00726f
C282 B.n242 VSUBS 0.00726f
C283 B.n243 VSUBS 0.00726f
C284 B.n244 VSUBS 0.00726f
C285 B.n245 VSUBS 0.00726f
C286 B.n246 VSUBS 0.00726f
C287 B.n247 VSUBS 0.00726f
C288 B.n248 VSUBS 0.00726f
C289 B.n249 VSUBS 0.00726f
C290 B.n250 VSUBS 0.00726f
C291 B.n251 VSUBS 0.00726f
C292 B.n252 VSUBS 0.00726f
C293 B.n253 VSUBS 0.00726f
C294 B.n254 VSUBS 0.00726f
C295 B.n255 VSUBS 0.00726f
C296 B.n256 VSUBS 0.00726f
C297 B.n257 VSUBS 0.00726f
C298 B.n258 VSUBS 0.00726f
C299 B.n259 VSUBS 0.00726f
C300 B.n260 VSUBS 0.00726f
C301 B.n261 VSUBS 0.00726f
C302 B.n262 VSUBS 0.00726f
C303 B.n263 VSUBS 0.00726f
C304 B.n264 VSUBS 0.00726f
C305 B.n265 VSUBS 0.00726f
C306 B.n266 VSUBS 0.00726f
C307 B.n267 VSUBS 0.00726f
C308 B.n268 VSUBS 0.00726f
C309 B.n269 VSUBS 0.00726f
C310 B.n270 VSUBS 0.00726f
C311 B.n271 VSUBS 0.00726f
C312 B.n272 VSUBS 0.00726f
C313 B.n273 VSUBS 0.00726f
C314 B.n274 VSUBS 0.00726f
C315 B.n275 VSUBS 0.00726f
C316 B.n276 VSUBS 0.00726f
C317 B.n277 VSUBS 0.00726f
C318 B.n278 VSUBS 0.017213f
C319 B.n279 VSUBS 0.015885f
C320 B.n280 VSUBS 0.015885f
C321 B.n281 VSUBS 0.00726f
C322 B.n282 VSUBS 0.00726f
C323 B.n283 VSUBS 0.00726f
C324 B.n284 VSUBS 0.00726f
C325 B.n285 VSUBS 0.00726f
C326 B.n286 VSUBS 0.00726f
C327 B.n287 VSUBS 0.00726f
C328 B.n288 VSUBS 0.00726f
C329 B.n289 VSUBS 0.00726f
C330 B.n290 VSUBS 0.00726f
C331 B.n291 VSUBS 0.00726f
C332 B.n292 VSUBS 0.00726f
C333 B.n293 VSUBS 0.00726f
C334 B.n294 VSUBS 0.00726f
C335 B.n295 VSUBS 0.00726f
C336 B.n296 VSUBS 0.00726f
C337 B.n297 VSUBS 0.00726f
C338 B.n298 VSUBS 0.00726f
C339 B.n299 VSUBS 0.00726f
C340 B.n300 VSUBS 0.00726f
C341 B.n301 VSUBS 0.00726f
C342 B.n302 VSUBS 0.00726f
C343 B.n303 VSUBS 0.00726f
C344 B.n304 VSUBS 0.00726f
C345 B.n305 VSUBS 0.00726f
C346 B.n306 VSUBS 0.00726f
C347 B.n307 VSUBS 0.00726f
C348 B.n308 VSUBS 0.00726f
C349 B.n309 VSUBS 0.00726f
C350 B.n310 VSUBS 0.00726f
C351 B.n311 VSUBS 0.00726f
C352 B.n312 VSUBS 0.00726f
C353 B.n313 VSUBS 0.00726f
C354 B.n314 VSUBS 0.00726f
C355 B.n315 VSUBS 0.00726f
C356 B.n316 VSUBS 0.00726f
C357 B.n317 VSUBS 0.00726f
C358 B.n318 VSUBS 0.00726f
C359 B.n319 VSUBS 0.00726f
C360 B.n320 VSUBS 0.00726f
C361 B.n321 VSUBS 0.00726f
C362 B.n322 VSUBS 0.00726f
C363 B.n323 VSUBS 0.00726f
C364 B.n324 VSUBS 0.00726f
C365 B.n325 VSUBS 0.00726f
C366 B.n326 VSUBS 0.00726f
C367 B.n327 VSUBS 0.016778f
C368 B.n328 VSUBS 0.015885f
C369 B.n329 VSUBS 0.017213f
C370 B.n330 VSUBS 0.00726f
C371 B.n331 VSUBS 0.00726f
C372 B.n332 VSUBS 0.00726f
C373 B.n333 VSUBS 0.00726f
C374 B.n334 VSUBS 0.00726f
C375 B.n335 VSUBS 0.00726f
C376 B.n336 VSUBS 0.00726f
C377 B.n337 VSUBS 0.00726f
C378 B.n338 VSUBS 0.00726f
C379 B.n339 VSUBS 0.00726f
C380 B.n340 VSUBS 0.00726f
C381 B.n341 VSUBS 0.00726f
C382 B.n342 VSUBS 0.00726f
C383 B.n343 VSUBS 0.00726f
C384 B.n344 VSUBS 0.00726f
C385 B.n345 VSUBS 0.00726f
C386 B.n346 VSUBS 0.00726f
C387 B.n347 VSUBS 0.00726f
C388 B.n348 VSUBS 0.00726f
C389 B.n349 VSUBS 0.00726f
C390 B.n350 VSUBS 0.00726f
C391 B.n351 VSUBS 0.00726f
C392 B.n352 VSUBS 0.00726f
C393 B.n353 VSUBS 0.00726f
C394 B.n354 VSUBS 0.00726f
C395 B.n355 VSUBS 0.00726f
C396 B.n356 VSUBS 0.00726f
C397 B.n357 VSUBS 0.00726f
C398 B.n358 VSUBS 0.00726f
C399 B.n359 VSUBS 0.00726f
C400 B.n360 VSUBS 0.00726f
C401 B.n361 VSUBS 0.00726f
C402 B.n362 VSUBS 0.00726f
C403 B.n363 VSUBS 0.00726f
C404 B.n364 VSUBS 0.00726f
C405 B.n365 VSUBS 0.00726f
C406 B.n366 VSUBS 0.00726f
C407 B.n367 VSUBS 0.00726f
C408 B.n368 VSUBS 0.00726f
C409 B.n369 VSUBS 0.00726f
C410 B.n370 VSUBS 0.00726f
C411 B.n371 VSUBS 0.00726f
C412 B.n372 VSUBS 0.00726f
C413 B.n373 VSUBS 0.00726f
C414 B.n374 VSUBS 0.00726f
C415 B.n375 VSUBS 0.00726f
C416 B.n376 VSUBS 0.00726f
C417 B.n377 VSUBS 0.00726f
C418 B.n378 VSUBS 0.00726f
C419 B.n379 VSUBS 0.00726f
C420 B.n380 VSUBS 0.00726f
C421 B.n381 VSUBS 0.00726f
C422 B.n382 VSUBS 0.00726f
C423 B.n383 VSUBS 0.00726f
C424 B.n384 VSUBS 0.00726f
C425 B.n385 VSUBS 0.004805f
C426 B.n386 VSUBS 0.016821f
C427 B.n387 VSUBS 0.006086f
C428 B.n388 VSUBS 0.00726f
C429 B.n389 VSUBS 0.00726f
C430 B.n390 VSUBS 0.00726f
C431 B.n391 VSUBS 0.00726f
C432 B.n392 VSUBS 0.00726f
C433 B.n393 VSUBS 0.00726f
C434 B.n394 VSUBS 0.00726f
C435 B.n395 VSUBS 0.00726f
C436 B.n396 VSUBS 0.00726f
C437 B.n397 VSUBS 0.00726f
C438 B.n398 VSUBS 0.00726f
C439 B.n399 VSUBS 0.006086f
C440 B.n400 VSUBS 0.016821f
C441 B.n401 VSUBS 0.004805f
C442 B.n402 VSUBS 0.00726f
C443 B.n403 VSUBS 0.00726f
C444 B.n404 VSUBS 0.00726f
C445 B.n405 VSUBS 0.00726f
C446 B.n406 VSUBS 0.00726f
C447 B.n407 VSUBS 0.00726f
C448 B.n408 VSUBS 0.00726f
C449 B.n409 VSUBS 0.00726f
C450 B.n410 VSUBS 0.00726f
C451 B.n411 VSUBS 0.00726f
C452 B.n412 VSUBS 0.00726f
C453 B.n413 VSUBS 0.00726f
C454 B.n414 VSUBS 0.00726f
C455 B.n415 VSUBS 0.00726f
C456 B.n416 VSUBS 0.00726f
C457 B.n417 VSUBS 0.00726f
C458 B.n418 VSUBS 0.00726f
C459 B.n419 VSUBS 0.00726f
C460 B.n420 VSUBS 0.00726f
C461 B.n421 VSUBS 0.00726f
C462 B.n422 VSUBS 0.00726f
C463 B.n423 VSUBS 0.00726f
C464 B.n424 VSUBS 0.00726f
C465 B.n425 VSUBS 0.00726f
C466 B.n426 VSUBS 0.00726f
C467 B.n427 VSUBS 0.00726f
C468 B.n428 VSUBS 0.00726f
C469 B.n429 VSUBS 0.00726f
C470 B.n430 VSUBS 0.00726f
C471 B.n431 VSUBS 0.00726f
C472 B.n432 VSUBS 0.00726f
C473 B.n433 VSUBS 0.00726f
C474 B.n434 VSUBS 0.00726f
C475 B.n435 VSUBS 0.00726f
C476 B.n436 VSUBS 0.00726f
C477 B.n437 VSUBS 0.00726f
C478 B.n438 VSUBS 0.00726f
C479 B.n439 VSUBS 0.00726f
C480 B.n440 VSUBS 0.00726f
C481 B.n441 VSUBS 0.00726f
C482 B.n442 VSUBS 0.00726f
C483 B.n443 VSUBS 0.00726f
C484 B.n444 VSUBS 0.00726f
C485 B.n445 VSUBS 0.00726f
C486 B.n446 VSUBS 0.00726f
C487 B.n447 VSUBS 0.00726f
C488 B.n448 VSUBS 0.00726f
C489 B.n449 VSUBS 0.00726f
C490 B.n450 VSUBS 0.00726f
C491 B.n451 VSUBS 0.00726f
C492 B.n452 VSUBS 0.00726f
C493 B.n453 VSUBS 0.00726f
C494 B.n454 VSUBS 0.00726f
C495 B.n455 VSUBS 0.00726f
C496 B.n456 VSUBS 0.00726f
C497 B.n457 VSUBS 0.017213f
C498 B.n458 VSUBS 0.015885f
C499 B.n459 VSUBS 0.015885f
C500 B.n460 VSUBS 0.00726f
C501 B.n461 VSUBS 0.00726f
C502 B.n462 VSUBS 0.00726f
C503 B.n463 VSUBS 0.00726f
C504 B.n464 VSUBS 0.00726f
C505 B.n465 VSUBS 0.00726f
C506 B.n466 VSUBS 0.00726f
C507 B.n467 VSUBS 0.00726f
C508 B.n468 VSUBS 0.00726f
C509 B.n469 VSUBS 0.00726f
C510 B.n470 VSUBS 0.00726f
C511 B.n471 VSUBS 0.00726f
C512 B.n472 VSUBS 0.00726f
C513 B.n473 VSUBS 0.00726f
C514 B.n474 VSUBS 0.00726f
C515 B.n475 VSUBS 0.00726f
C516 B.n476 VSUBS 0.00726f
C517 B.n477 VSUBS 0.00726f
C518 B.n478 VSUBS 0.00726f
C519 B.n479 VSUBS 0.00726f
C520 B.n480 VSUBS 0.00726f
C521 B.n481 VSUBS 0.00726f
C522 B.n482 VSUBS 0.00726f
C523 B.n483 VSUBS 0.01644f
C524 VDD1.n0 VSUBS 0.020748f
C525 VDD1.n1 VSUBS 0.020375f
C526 VDD1.n2 VSUBS 0.010949f
C527 VDD1.n3 VSUBS 0.025879f
C528 VDD1.n4 VSUBS 0.011593f
C529 VDD1.n5 VSUBS 0.020375f
C530 VDD1.n6 VSUBS 0.010949f
C531 VDD1.n7 VSUBS 0.025879f
C532 VDD1.n8 VSUBS 0.011593f
C533 VDD1.n9 VSUBS 0.020375f
C534 VDD1.n10 VSUBS 0.010949f
C535 VDD1.n11 VSUBS 0.025879f
C536 VDD1.n12 VSUBS 0.025879f
C537 VDD1.n13 VSUBS 0.011593f
C538 VDD1.n14 VSUBS 0.020375f
C539 VDD1.n15 VSUBS 0.010949f
C540 VDD1.n16 VSUBS 0.025879f
C541 VDD1.n17 VSUBS 0.011593f
C542 VDD1.n18 VSUBS 0.147387f
C543 VDD1.t1 VSUBS 0.055672f
C544 VDD1.n19 VSUBS 0.019409f
C545 VDD1.n20 VSUBS 0.019467f
C546 VDD1.n21 VSUBS 0.010949f
C547 VDD1.n22 VSUBS 0.874314f
C548 VDD1.n23 VSUBS 0.020375f
C549 VDD1.n24 VSUBS 0.010949f
C550 VDD1.n25 VSUBS 0.011593f
C551 VDD1.n26 VSUBS 0.025879f
C552 VDD1.n27 VSUBS 0.025879f
C553 VDD1.n28 VSUBS 0.011593f
C554 VDD1.n29 VSUBS 0.010949f
C555 VDD1.n30 VSUBS 0.020375f
C556 VDD1.n31 VSUBS 0.020375f
C557 VDD1.n32 VSUBS 0.010949f
C558 VDD1.n33 VSUBS 0.011593f
C559 VDD1.n34 VSUBS 0.025879f
C560 VDD1.n35 VSUBS 0.025879f
C561 VDD1.n36 VSUBS 0.011593f
C562 VDD1.n37 VSUBS 0.010949f
C563 VDD1.n38 VSUBS 0.020375f
C564 VDD1.n39 VSUBS 0.020375f
C565 VDD1.n40 VSUBS 0.010949f
C566 VDD1.n41 VSUBS 0.011271f
C567 VDD1.n42 VSUBS 0.011271f
C568 VDD1.n43 VSUBS 0.025879f
C569 VDD1.n44 VSUBS 0.025879f
C570 VDD1.n45 VSUBS 0.011593f
C571 VDD1.n46 VSUBS 0.010949f
C572 VDD1.n47 VSUBS 0.020375f
C573 VDD1.n48 VSUBS 0.020375f
C574 VDD1.n49 VSUBS 0.010949f
C575 VDD1.n50 VSUBS 0.011593f
C576 VDD1.n51 VSUBS 0.025879f
C577 VDD1.n52 VSUBS 0.057064f
C578 VDD1.n53 VSUBS 0.011593f
C579 VDD1.n54 VSUBS 0.010949f
C580 VDD1.n55 VSUBS 0.044313f
C581 VDD1.n56 VSUBS 0.042904f
C582 VDD1.n57 VSUBS 0.020748f
C583 VDD1.n58 VSUBS 0.020375f
C584 VDD1.n59 VSUBS 0.010949f
C585 VDD1.n60 VSUBS 0.025879f
C586 VDD1.n61 VSUBS 0.011593f
C587 VDD1.n62 VSUBS 0.020375f
C588 VDD1.n63 VSUBS 0.010949f
C589 VDD1.n64 VSUBS 0.025879f
C590 VDD1.n65 VSUBS 0.011593f
C591 VDD1.n66 VSUBS 0.020375f
C592 VDD1.n67 VSUBS 0.010949f
C593 VDD1.n68 VSUBS 0.025879f
C594 VDD1.n69 VSUBS 0.011593f
C595 VDD1.n70 VSUBS 0.020375f
C596 VDD1.n71 VSUBS 0.010949f
C597 VDD1.n72 VSUBS 0.025879f
C598 VDD1.n73 VSUBS 0.011593f
C599 VDD1.n74 VSUBS 0.147387f
C600 VDD1.t0 VSUBS 0.055672f
C601 VDD1.n75 VSUBS 0.019409f
C602 VDD1.n76 VSUBS 0.019467f
C603 VDD1.n77 VSUBS 0.010949f
C604 VDD1.n78 VSUBS 0.874314f
C605 VDD1.n79 VSUBS 0.020375f
C606 VDD1.n80 VSUBS 0.010949f
C607 VDD1.n81 VSUBS 0.011593f
C608 VDD1.n82 VSUBS 0.025879f
C609 VDD1.n83 VSUBS 0.025879f
C610 VDD1.n84 VSUBS 0.011593f
C611 VDD1.n85 VSUBS 0.010949f
C612 VDD1.n86 VSUBS 0.020375f
C613 VDD1.n87 VSUBS 0.020375f
C614 VDD1.n88 VSUBS 0.010949f
C615 VDD1.n89 VSUBS 0.011593f
C616 VDD1.n90 VSUBS 0.025879f
C617 VDD1.n91 VSUBS 0.025879f
C618 VDD1.n92 VSUBS 0.025879f
C619 VDD1.n93 VSUBS 0.011593f
C620 VDD1.n94 VSUBS 0.010949f
C621 VDD1.n95 VSUBS 0.020375f
C622 VDD1.n96 VSUBS 0.020375f
C623 VDD1.n97 VSUBS 0.010949f
C624 VDD1.n98 VSUBS 0.011271f
C625 VDD1.n99 VSUBS 0.011271f
C626 VDD1.n100 VSUBS 0.025879f
C627 VDD1.n101 VSUBS 0.025879f
C628 VDD1.n102 VSUBS 0.011593f
C629 VDD1.n103 VSUBS 0.010949f
C630 VDD1.n104 VSUBS 0.020375f
C631 VDD1.n105 VSUBS 0.020375f
C632 VDD1.n106 VSUBS 0.010949f
C633 VDD1.n107 VSUBS 0.011593f
C634 VDD1.n108 VSUBS 0.025879f
C635 VDD1.n109 VSUBS 0.057064f
C636 VDD1.n110 VSUBS 0.011593f
C637 VDD1.n111 VSUBS 0.010949f
C638 VDD1.n112 VSUBS 0.044313f
C639 VDD1.n113 VSUBS 0.514725f
C640 VP.t0 VSUBS 2.07575f
C641 VP.t1 VSUBS 1.88169f
C642 VP.n0 VSUBS 4.61342f
C643 VDD2.n0 VSUBS 0.020977f
C644 VDD2.n1 VSUBS 0.0206f
C645 VDD2.n2 VSUBS 0.011069f
C646 VDD2.n3 VSUBS 0.026164f
C647 VDD2.n4 VSUBS 0.011721f
C648 VDD2.n5 VSUBS 0.0206f
C649 VDD2.n6 VSUBS 0.011069f
C650 VDD2.n7 VSUBS 0.026164f
C651 VDD2.n8 VSUBS 0.011721f
C652 VDD2.n9 VSUBS 0.0206f
C653 VDD2.n10 VSUBS 0.011069f
C654 VDD2.n11 VSUBS 0.026164f
C655 VDD2.n12 VSUBS 0.011721f
C656 VDD2.n13 VSUBS 0.0206f
C657 VDD2.n14 VSUBS 0.011069f
C658 VDD2.n15 VSUBS 0.026164f
C659 VDD2.n16 VSUBS 0.011721f
C660 VDD2.n17 VSUBS 0.149012f
C661 VDD2.t1 VSUBS 0.056286f
C662 VDD2.n18 VSUBS 0.019623f
C663 VDD2.n19 VSUBS 0.019682f
C664 VDD2.n20 VSUBS 0.011069f
C665 VDD2.n21 VSUBS 0.883955f
C666 VDD2.n22 VSUBS 0.0206f
C667 VDD2.n23 VSUBS 0.011069f
C668 VDD2.n24 VSUBS 0.011721f
C669 VDD2.n25 VSUBS 0.026164f
C670 VDD2.n26 VSUBS 0.026164f
C671 VDD2.n27 VSUBS 0.011721f
C672 VDD2.n28 VSUBS 0.011069f
C673 VDD2.n29 VSUBS 0.0206f
C674 VDD2.n30 VSUBS 0.0206f
C675 VDD2.n31 VSUBS 0.011069f
C676 VDD2.n32 VSUBS 0.011721f
C677 VDD2.n33 VSUBS 0.026164f
C678 VDD2.n34 VSUBS 0.026164f
C679 VDD2.n35 VSUBS 0.026164f
C680 VDD2.n36 VSUBS 0.011721f
C681 VDD2.n37 VSUBS 0.011069f
C682 VDD2.n38 VSUBS 0.0206f
C683 VDD2.n39 VSUBS 0.0206f
C684 VDD2.n40 VSUBS 0.011069f
C685 VDD2.n41 VSUBS 0.011395f
C686 VDD2.n42 VSUBS 0.011395f
C687 VDD2.n43 VSUBS 0.026164f
C688 VDD2.n44 VSUBS 0.026164f
C689 VDD2.n45 VSUBS 0.011721f
C690 VDD2.n46 VSUBS 0.011069f
C691 VDD2.n47 VSUBS 0.0206f
C692 VDD2.n48 VSUBS 0.0206f
C693 VDD2.n49 VSUBS 0.011069f
C694 VDD2.n50 VSUBS 0.011721f
C695 VDD2.n51 VSUBS 0.026164f
C696 VDD2.n52 VSUBS 0.057693f
C697 VDD2.n53 VSUBS 0.011721f
C698 VDD2.n54 VSUBS 0.011069f
C699 VDD2.n55 VSUBS 0.044801f
C700 VDD2.n56 VSUBS 0.490981f
C701 VDD2.n57 VSUBS 0.020977f
C702 VDD2.n58 VSUBS 0.0206f
C703 VDD2.n59 VSUBS 0.011069f
C704 VDD2.n60 VSUBS 0.026164f
C705 VDD2.n61 VSUBS 0.011721f
C706 VDD2.n62 VSUBS 0.0206f
C707 VDD2.n63 VSUBS 0.011069f
C708 VDD2.n64 VSUBS 0.026164f
C709 VDD2.n65 VSUBS 0.011721f
C710 VDD2.n66 VSUBS 0.0206f
C711 VDD2.n67 VSUBS 0.011069f
C712 VDD2.n68 VSUBS 0.026164f
C713 VDD2.n69 VSUBS 0.026164f
C714 VDD2.n70 VSUBS 0.011721f
C715 VDD2.n71 VSUBS 0.0206f
C716 VDD2.n72 VSUBS 0.011069f
C717 VDD2.n73 VSUBS 0.026164f
C718 VDD2.n74 VSUBS 0.011721f
C719 VDD2.n75 VSUBS 0.149012f
C720 VDD2.t0 VSUBS 0.056286f
C721 VDD2.n76 VSUBS 0.019623f
C722 VDD2.n77 VSUBS 0.019682f
C723 VDD2.n78 VSUBS 0.011069f
C724 VDD2.n79 VSUBS 0.883955f
C725 VDD2.n80 VSUBS 0.0206f
C726 VDD2.n81 VSUBS 0.011069f
C727 VDD2.n82 VSUBS 0.011721f
C728 VDD2.n83 VSUBS 0.026164f
C729 VDD2.n84 VSUBS 0.026164f
C730 VDD2.n85 VSUBS 0.011721f
C731 VDD2.n86 VSUBS 0.011069f
C732 VDD2.n87 VSUBS 0.0206f
C733 VDD2.n88 VSUBS 0.0206f
C734 VDD2.n89 VSUBS 0.011069f
C735 VDD2.n90 VSUBS 0.011721f
C736 VDD2.n91 VSUBS 0.026164f
C737 VDD2.n92 VSUBS 0.026164f
C738 VDD2.n93 VSUBS 0.011721f
C739 VDD2.n94 VSUBS 0.011069f
C740 VDD2.n95 VSUBS 0.0206f
C741 VDD2.n96 VSUBS 0.0206f
C742 VDD2.n97 VSUBS 0.011069f
C743 VDD2.n98 VSUBS 0.011395f
C744 VDD2.n99 VSUBS 0.011395f
C745 VDD2.n100 VSUBS 0.026164f
C746 VDD2.n101 VSUBS 0.026164f
C747 VDD2.n102 VSUBS 0.011721f
C748 VDD2.n103 VSUBS 0.011069f
C749 VDD2.n104 VSUBS 0.0206f
C750 VDD2.n105 VSUBS 0.0206f
C751 VDD2.n106 VSUBS 0.011069f
C752 VDD2.n107 VSUBS 0.011721f
C753 VDD2.n108 VSUBS 0.026164f
C754 VDD2.n109 VSUBS 0.057693f
C755 VDD2.n110 VSUBS 0.011721f
C756 VDD2.n111 VSUBS 0.011069f
C757 VDD2.n112 VSUBS 0.044801f
C758 VDD2.n113 VSUBS 0.042921f
C759 VDD2.n114 VSUBS 2.12687f
C760 VTAIL.n0 VSUBS 0.024372f
C761 VTAIL.n1 VSUBS 0.023934f
C762 VTAIL.n2 VSUBS 0.012861f
C763 VTAIL.n3 VSUBS 0.030399f
C764 VTAIL.n4 VSUBS 0.013618f
C765 VTAIL.n5 VSUBS 0.023934f
C766 VTAIL.n6 VSUBS 0.012861f
C767 VTAIL.n7 VSUBS 0.030399f
C768 VTAIL.n8 VSUBS 0.013618f
C769 VTAIL.n9 VSUBS 0.023934f
C770 VTAIL.n10 VSUBS 0.012861f
C771 VTAIL.n11 VSUBS 0.030399f
C772 VTAIL.n12 VSUBS 0.013618f
C773 VTAIL.n13 VSUBS 0.023934f
C774 VTAIL.n14 VSUBS 0.012861f
C775 VTAIL.n15 VSUBS 0.030399f
C776 VTAIL.n16 VSUBS 0.013618f
C777 VTAIL.n17 VSUBS 0.17313f
C778 VTAIL.t3 VSUBS 0.065396f
C779 VTAIL.n18 VSUBS 0.022799f
C780 VTAIL.n19 VSUBS 0.022868f
C781 VTAIL.n20 VSUBS 0.012861f
C782 VTAIL.n21 VSUBS 1.02702f
C783 VTAIL.n22 VSUBS 0.023934f
C784 VTAIL.n23 VSUBS 0.012861f
C785 VTAIL.n24 VSUBS 0.013618f
C786 VTAIL.n25 VSUBS 0.030399f
C787 VTAIL.n26 VSUBS 0.030399f
C788 VTAIL.n27 VSUBS 0.013618f
C789 VTAIL.n28 VSUBS 0.012861f
C790 VTAIL.n29 VSUBS 0.023934f
C791 VTAIL.n30 VSUBS 0.023934f
C792 VTAIL.n31 VSUBS 0.012861f
C793 VTAIL.n32 VSUBS 0.013618f
C794 VTAIL.n33 VSUBS 0.030399f
C795 VTAIL.n34 VSUBS 0.030399f
C796 VTAIL.n35 VSUBS 0.030399f
C797 VTAIL.n36 VSUBS 0.013618f
C798 VTAIL.n37 VSUBS 0.012861f
C799 VTAIL.n38 VSUBS 0.023934f
C800 VTAIL.n39 VSUBS 0.023934f
C801 VTAIL.n40 VSUBS 0.012861f
C802 VTAIL.n41 VSUBS 0.013239f
C803 VTAIL.n42 VSUBS 0.013239f
C804 VTAIL.n43 VSUBS 0.030399f
C805 VTAIL.n44 VSUBS 0.030399f
C806 VTAIL.n45 VSUBS 0.013618f
C807 VTAIL.n46 VSUBS 0.012861f
C808 VTAIL.n47 VSUBS 0.023934f
C809 VTAIL.n48 VSUBS 0.023934f
C810 VTAIL.n49 VSUBS 0.012861f
C811 VTAIL.n50 VSUBS 0.013618f
C812 VTAIL.n51 VSUBS 0.030399f
C813 VTAIL.n52 VSUBS 0.067031f
C814 VTAIL.n53 VSUBS 0.013618f
C815 VTAIL.n54 VSUBS 0.012861f
C816 VTAIL.n55 VSUBS 0.052052f
C817 VTAIL.n56 VSUBS 0.033314f
C818 VTAIL.n57 VSUBS 1.29259f
C819 VTAIL.n58 VSUBS 0.024372f
C820 VTAIL.n59 VSUBS 0.023934f
C821 VTAIL.n60 VSUBS 0.012861f
C822 VTAIL.n61 VSUBS 0.030399f
C823 VTAIL.n62 VSUBS 0.013618f
C824 VTAIL.n63 VSUBS 0.023934f
C825 VTAIL.n64 VSUBS 0.012861f
C826 VTAIL.n65 VSUBS 0.030399f
C827 VTAIL.n66 VSUBS 0.013618f
C828 VTAIL.n67 VSUBS 0.023934f
C829 VTAIL.n68 VSUBS 0.012861f
C830 VTAIL.n69 VSUBS 0.030399f
C831 VTAIL.n70 VSUBS 0.030399f
C832 VTAIL.n71 VSUBS 0.013618f
C833 VTAIL.n72 VSUBS 0.023934f
C834 VTAIL.n73 VSUBS 0.012861f
C835 VTAIL.n74 VSUBS 0.030399f
C836 VTAIL.n75 VSUBS 0.013618f
C837 VTAIL.n76 VSUBS 0.17313f
C838 VTAIL.t2 VSUBS 0.065396f
C839 VTAIL.n77 VSUBS 0.022799f
C840 VTAIL.n78 VSUBS 0.022868f
C841 VTAIL.n79 VSUBS 0.012861f
C842 VTAIL.n80 VSUBS 1.02702f
C843 VTAIL.n81 VSUBS 0.023934f
C844 VTAIL.n82 VSUBS 0.012861f
C845 VTAIL.n83 VSUBS 0.013618f
C846 VTAIL.n84 VSUBS 0.030399f
C847 VTAIL.n85 VSUBS 0.030399f
C848 VTAIL.n86 VSUBS 0.013618f
C849 VTAIL.n87 VSUBS 0.012861f
C850 VTAIL.n88 VSUBS 0.023934f
C851 VTAIL.n89 VSUBS 0.023934f
C852 VTAIL.n90 VSUBS 0.012861f
C853 VTAIL.n91 VSUBS 0.013618f
C854 VTAIL.n92 VSUBS 0.030399f
C855 VTAIL.n93 VSUBS 0.030399f
C856 VTAIL.n94 VSUBS 0.013618f
C857 VTAIL.n95 VSUBS 0.012861f
C858 VTAIL.n96 VSUBS 0.023934f
C859 VTAIL.n97 VSUBS 0.023934f
C860 VTAIL.n98 VSUBS 0.012861f
C861 VTAIL.n99 VSUBS 0.013239f
C862 VTAIL.n100 VSUBS 0.013239f
C863 VTAIL.n101 VSUBS 0.030399f
C864 VTAIL.n102 VSUBS 0.030399f
C865 VTAIL.n103 VSUBS 0.013618f
C866 VTAIL.n104 VSUBS 0.012861f
C867 VTAIL.n105 VSUBS 0.023934f
C868 VTAIL.n106 VSUBS 0.023934f
C869 VTAIL.n107 VSUBS 0.012861f
C870 VTAIL.n108 VSUBS 0.013618f
C871 VTAIL.n109 VSUBS 0.030399f
C872 VTAIL.n110 VSUBS 0.067031f
C873 VTAIL.n111 VSUBS 0.013618f
C874 VTAIL.n112 VSUBS 0.012861f
C875 VTAIL.n113 VSUBS 0.052052f
C876 VTAIL.n114 VSUBS 0.033314f
C877 VTAIL.n115 VSUBS 1.3107f
C878 VTAIL.n116 VSUBS 0.024372f
C879 VTAIL.n117 VSUBS 0.023934f
C880 VTAIL.n118 VSUBS 0.012861f
C881 VTAIL.n119 VSUBS 0.030399f
C882 VTAIL.n120 VSUBS 0.013618f
C883 VTAIL.n121 VSUBS 0.023934f
C884 VTAIL.n122 VSUBS 0.012861f
C885 VTAIL.n123 VSUBS 0.030399f
C886 VTAIL.n124 VSUBS 0.013618f
C887 VTAIL.n125 VSUBS 0.023934f
C888 VTAIL.n126 VSUBS 0.012861f
C889 VTAIL.n127 VSUBS 0.030399f
C890 VTAIL.n128 VSUBS 0.030399f
C891 VTAIL.n129 VSUBS 0.013618f
C892 VTAIL.n130 VSUBS 0.023934f
C893 VTAIL.n131 VSUBS 0.012861f
C894 VTAIL.n132 VSUBS 0.030399f
C895 VTAIL.n133 VSUBS 0.013618f
C896 VTAIL.n134 VSUBS 0.17313f
C897 VTAIL.t0 VSUBS 0.065396f
C898 VTAIL.n135 VSUBS 0.022799f
C899 VTAIL.n136 VSUBS 0.022868f
C900 VTAIL.n137 VSUBS 0.012861f
C901 VTAIL.n138 VSUBS 1.02702f
C902 VTAIL.n139 VSUBS 0.023934f
C903 VTAIL.n140 VSUBS 0.012861f
C904 VTAIL.n141 VSUBS 0.013618f
C905 VTAIL.n142 VSUBS 0.030399f
C906 VTAIL.n143 VSUBS 0.030399f
C907 VTAIL.n144 VSUBS 0.013618f
C908 VTAIL.n145 VSUBS 0.012861f
C909 VTAIL.n146 VSUBS 0.023934f
C910 VTAIL.n147 VSUBS 0.023934f
C911 VTAIL.n148 VSUBS 0.012861f
C912 VTAIL.n149 VSUBS 0.013618f
C913 VTAIL.n150 VSUBS 0.030399f
C914 VTAIL.n151 VSUBS 0.030399f
C915 VTAIL.n152 VSUBS 0.013618f
C916 VTAIL.n153 VSUBS 0.012861f
C917 VTAIL.n154 VSUBS 0.023934f
C918 VTAIL.n155 VSUBS 0.023934f
C919 VTAIL.n156 VSUBS 0.012861f
C920 VTAIL.n157 VSUBS 0.013239f
C921 VTAIL.n158 VSUBS 0.013239f
C922 VTAIL.n159 VSUBS 0.030399f
C923 VTAIL.n160 VSUBS 0.030399f
C924 VTAIL.n161 VSUBS 0.013618f
C925 VTAIL.n162 VSUBS 0.012861f
C926 VTAIL.n163 VSUBS 0.023934f
C927 VTAIL.n164 VSUBS 0.023934f
C928 VTAIL.n165 VSUBS 0.012861f
C929 VTAIL.n166 VSUBS 0.013618f
C930 VTAIL.n167 VSUBS 0.030399f
C931 VTAIL.n168 VSUBS 0.067031f
C932 VTAIL.n169 VSUBS 0.013618f
C933 VTAIL.n170 VSUBS 0.012861f
C934 VTAIL.n171 VSUBS 0.052052f
C935 VTAIL.n172 VSUBS 0.033314f
C936 VTAIL.n173 VSUBS 1.22029f
C937 VTAIL.n174 VSUBS 0.024372f
C938 VTAIL.n175 VSUBS 0.023934f
C939 VTAIL.n176 VSUBS 0.012861f
C940 VTAIL.n177 VSUBS 0.030399f
C941 VTAIL.n178 VSUBS 0.013618f
C942 VTAIL.n179 VSUBS 0.023934f
C943 VTAIL.n180 VSUBS 0.012861f
C944 VTAIL.n181 VSUBS 0.030399f
C945 VTAIL.n182 VSUBS 0.013618f
C946 VTAIL.n183 VSUBS 0.023934f
C947 VTAIL.n184 VSUBS 0.012861f
C948 VTAIL.n185 VSUBS 0.030399f
C949 VTAIL.n186 VSUBS 0.013618f
C950 VTAIL.n187 VSUBS 0.023934f
C951 VTAIL.n188 VSUBS 0.012861f
C952 VTAIL.n189 VSUBS 0.030399f
C953 VTAIL.n190 VSUBS 0.013618f
C954 VTAIL.n191 VSUBS 0.17313f
C955 VTAIL.t1 VSUBS 0.065396f
C956 VTAIL.n192 VSUBS 0.022799f
C957 VTAIL.n193 VSUBS 0.022868f
C958 VTAIL.n194 VSUBS 0.012861f
C959 VTAIL.n195 VSUBS 1.02702f
C960 VTAIL.n196 VSUBS 0.023934f
C961 VTAIL.n197 VSUBS 0.012861f
C962 VTAIL.n198 VSUBS 0.013618f
C963 VTAIL.n199 VSUBS 0.030399f
C964 VTAIL.n200 VSUBS 0.030399f
C965 VTAIL.n201 VSUBS 0.013618f
C966 VTAIL.n202 VSUBS 0.012861f
C967 VTAIL.n203 VSUBS 0.023934f
C968 VTAIL.n204 VSUBS 0.023934f
C969 VTAIL.n205 VSUBS 0.012861f
C970 VTAIL.n206 VSUBS 0.013618f
C971 VTAIL.n207 VSUBS 0.030399f
C972 VTAIL.n208 VSUBS 0.030399f
C973 VTAIL.n209 VSUBS 0.030399f
C974 VTAIL.n210 VSUBS 0.013618f
C975 VTAIL.n211 VSUBS 0.012861f
C976 VTAIL.n212 VSUBS 0.023934f
C977 VTAIL.n213 VSUBS 0.023934f
C978 VTAIL.n214 VSUBS 0.012861f
C979 VTAIL.n215 VSUBS 0.013239f
C980 VTAIL.n216 VSUBS 0.013239f
C981 VTAIL.n217 VSUBS 0.030399f
C982 VTAIL.n218 VSUBS 0.030399f
C983 VTAIL.n219 VSUBS 0.013618f
C984 VTAIL.n220 VSUBS 0.012861f
C985 VTAIL.n221 VSUBS 0.023934f
C986 VTAIL.n222 VSUBS 0.023934f
C987 VTAIL.n223 VSUBS 0.012861f
C988 VTAIL.n224 VSUBS 0.013618f
C989 VTAIL.n225 VSUBS 0.030399f
C990 VTAIL.n226 VSUBS 0.067031f
C991 VTAIL.n227 VSUBS 0.013618f
C992 VTAIL.n228 VSUBS 0.012861f
C993 VTAIL.n229 VSUBS 0.052052f
C994 VTAIL.n230 VSUBS 0.033314f
C995 VTAIL.n231 VSUBS 1.15696f
C996 VN.t0 VSUBS 1.38838f
C997 VN.t1 VSUBS 1.53489f
.ends

