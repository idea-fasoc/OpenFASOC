* NGSPICE file created from diff_pair_sample_0502.ext - technology: sky130A

.subckt diff_pair_sample_0502 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=0 ps=0 w=15.15 l=1.48
X1 VDD2.t5 VN.t0 VTAIL.t5 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=2.49975 ps=15.48 w=15.15 l=1.48
X2 B.t8 B.t6 B.t7 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=0 ps=0 w=15.15 l=1.48
X3 VDD1.t5 VP.t0 VTAIL.t3 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=2.49975 ps=15.48 w=15.15 l=1.48
X4 VDD2.t4 VN.t1 VTAIL.t6 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=5.9085 ps=31.08 w=15.15 l=1.48
X5 B.t5 B.t3 B.t4 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=0 ps=0 w=15.15 l=1.48
X6 B.t2 B.t0 B.t1 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=0 ps=0 w=15.15 l=1.48
X7 VDD2.t3 VN.t2 VTAIL.t9 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=2.49975 ps=15.48 w=15.15 l=1.48
X8 VDD2.t2 VN.t3 VTAIL.t7 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=5.9085 ps=31.08 w=15.15 l=1.48
X9 VTAIL.t8 VN.t4 VDD2.t1 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=2.49975 ps=15.48 w=15.15 l=1.48
X10 VTAIL.t0 VP.t1 VDD1.t4 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=2.49975 ps=15.48 w=15.15 l=1.48
X11 VDD1.t3 VP.t2 VTAIL.t4 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=5.9085 ps=31.08 w=15.15 l=1.48
X12 VDD1.t2 VP.t3 VTAIL.t1 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=5.9085 ps=31.08 w=15.15 l=1.48
X13 VTAIL.t11 VP.t4 VDD1.t1 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=2.49975 ps=15.48 w=15.15 l=1.48
X14 VDD1.t0 VP.t5 VTAIL.t2 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=5.9085 pd=31.08 as=2.49975 ps=15.48 w=15.15 l=1.48
X15 VTAIL.t10 VN.t5 VDD2.t0 w_n2418_n3998# sky130_fd_pr__pfet_01v8 ad=2.49975 pd=15.48 as=2.49975 ps=15.48 w=15.15 l=1.48
R0 B.n390 B.n389 585
R1 B.n388 B.n107 585
R2 B.n387 B.n386 585
R3 B.n385 B.n108 585
R4 B.n384 B.n383 585
R5 B.n382 B.n109 585
R6 B.n381 B.n380 585
R7 B.n379 B.n110 585
R8 B.n378 B.n377 585
R9 B.n376 B.n111 585
R10 B.n375 B.n374 585
R11 B.n373 B.n112 585
R12 B.n372 B.n371 585
R13 B.n370 B.n113 585
R14 B.n369 B.n368 585
R15 B.n367 B.n114 585
R16 B.n366 B.n365 585
R17 B.n364 B.n115 585
R18 B.n363 B.n362 585
R19 B.n361 B.n116 585
R20 B.n360 B.n359 585
R21 B.n358 B.n117 585
R22 B.n357 B.n356 585
R23 B.n355 B.n118 585
R24 B.n354 B.n353 585
R25 B.n352 B.n119 585
R26 B.n351 B.n350 585
R27 B.n349 B.n120 585
R28 B.n348 B.n347 585
R29 B.n346 B.n121 585
R30 B.n345 B.n344 585
R31 B.n343 B.n122 585
R32 B.n342 B.n341 585
R33 B.n340 B.n123 585
R34 B.n339 B.n338 585
R35 B.n337 B.n124 585
R36 B.n336 B.n335 585
R37 B.n334 B.n125 585
R38 B.n333 B.n332 585
R39 B.n331 B.n126 585
R40 B.n330 B.n329 585
R41 B.n328 B.n127 585
R42 B.n327 B.n326 585
R43 B.n325 B.n128 585
R44 B.n324 B.n323 585
R45 B.n322 B.n129 585
R46 B.n321 B.n320 585
R47 B.n319 B.n130 585
R48 B.n318 B.n317 585
R49 B.n316 B.n131 585
R50 B.n315 B.n314 585
R51 B.n313 B.n312 585
R52 B.n311 B.n135 585
R53 B.n310 B.n309 585
R54 B.n308 B.n136 585
R55 B.n307 B.n306 585
R56 B.n305 B.n137 585
R57 B.n304 B.n303 585
R58 B.n302 B.n138 585
R59 B.n301 B.n300 585
R60 B.n298 B.n139 585
R61 B.n297 B.n296 585
R62 B.n295 B.n142 585
R63 B.n294 B.n293 585
R64 B.n292 B.n143 585
R65 B.n291 B.n290 585
R66 B.n289 B.n144 585
R67 B.n288 B.n287 585
R68 B.n286 B.n145 585
R69 B.n285 B.n284 585
R70 B.n283 B.n146 585
R71 B.n282 B.n281 585
R72 B.n280 B.n147 585
R73 B.n279 B.n278 585
R74 B.n277 B.n148 585
R75 B.n276 B.n275 585
R76 B.n274 B.n149 585
R77 B.n273 B.n272 585
R78 B.n271 B.n150 585
R79 B.n270 B.n269 585
R80 B.n268 B.n151 585
R81 B.n267 B.n266 585
R82 B.n265 B.n152 585
R83 B.n264 B.n263 585
R84 B.n262 B.n153 585
R85 B.n261 B.n260 585
R86 B.n259 B.n154 585
R87 B.n258 B.n257 585
R88 B.n256 B.n155 585
R89 B.n255 B.n254 585
R90 B.n253 B.n156 585
R91 B.n252 B.n251 585
R92 B.n250 B.n157 585
R93 B.n249 B.n248 585
R94 B.n247 B.n158 585
R95 B.n246 B.n245 585
R96 B.n244 B.n159 585
R97 B.n243 B.n242 585
R98 B.n241 B.n160 585
R99 B.n240 B.n239 585
R100 B.n238 B.n161 585
R101 B.n237 B.n236 585
R102 B.n235 B.n162 585
R103 B.n234 B.n233 585
R104 B.n232 B.n163 585
R105 B.n231 B.n230 585
R106 B.n229 B.n164 585
R107 B.n228 B.n227 585
R108 B.n226 B.n165 585
R109 B.n225 B.n224 585
R110 B.n223 B.n166 585
R111 B.n391 B.n106 585
R112 B.n393 B.n392 585
R113 B.n394 B.n105 585
R114 B.n396 B.n395 585
R115 B.n397 B.n104 585
R116 B.n399 B.n398 585
R117 B.n400 B.n103 585
R118 B.n402 B.n401 585
R119 B.n403 B.n102 585
R120 B.n405 B.n404 585
R121 B.n406 B.n101 585
R122 B.n408 B.n407 585
R123 B.n409 B.n100 585
R124 B.n411 B.n410 585
R125 B.n412 B.n99 585
R126 B.n414 B.n413 585
R127 B.n415 B.n98 585
R128 B.n417 B.n416 585
R129 B.n418 B.n97 585
R130 B.n420 B.n419 585
R131 B.n421 B.n96 585
R132 B.n423 B.n422 585
R133 B.n424 B.n95 585
R134 B.n426 B.n425 585
R135 B.n427 B.n94 585
R136 B.n429 B.n428 585
R137 B.n430 B.n93 585
R138 B.n432 B.n431 585
R139 B.n433 B.n92 585
R140 B.n435 B.n434 585
R141 B.n436 B.n91 585
R142 B.n438 B.n437 585
R143 B.n439 B.n90 585
R144 B.n441 B.n440 585
R145 B.n442 B.n89 585
R146 B.n444 B.n443 585
R147 B.n445 B.n88 585
R148 B.n447 B.n446 585
R149 B.n448 B.n87 585
R150 B.n450 B.n449 585
R151 B.n451 B.n86 585
R152 B.n453 B.n452 585
R153 B.n454 B.n85 585
R154 B.n456 B.n455 585
R155 B.n457 B.n84 585
R156 B.n459 B.n458 585
R157 B.n460 B.n83 585
R158 B.n462 B.n461 585
R159 B.n463 B.n82 585
R160 B.n465 B.n464 585
R161 B.n466 B.n81 585
R162 B.n468 B.n467 585
R163 B.n469 B.n80 585
R164 B.n471 B.n470 585
R165 B.n472 B.n79 585
R166 B.n474 B.n473 585
R167 B.n475 B.n78 585
R168 B.n477 B.n476 585
R169 B.n478 B.n77 585
R170 B.n480 B.n479 585
R171 B.n648 B.n647 585
R172 B.n646 B.n17 585
R173 B.n645 B.n644 585
R174 B.n643 B.n18 585
R175 B.n642 B.n641 585
R176 B.n640 B.n19 585
R177 B.n639 B.n638 585
R178 B.n637 B.n20 585
R179 B.n636 B.n635 585
R180 B.n634 B.n21 585
R181 B.n633 B.n632 585
R182 B.n631 B.n22 585
R183 B.n630 B.n629 585
R184 B.n628 B.n23 585
R185 B.n627 B.n626 585
R186 B.n625 B.n24 585
R187 B.n624 B.n623 585
R188 B.n622 B.n25 585
R189 B.n621 B.n620 585
R190 B.n619 B.n26 585
R191 B.n618 B.n617 585
R192 B.n616 B.n27 585
R193 B.n615 B.n614 585
R194 B.n613 B.n28 585
R195 B.n612 B.n611 585
R196 B.n610 B.n29 585
R197 B.n609 B.n608 585
R198 B.n607 B.n30 585
R199 B.n606 B.n605 585
R200 B.n604 B.n31 585
R201 B.n603 B.n602 585
R202 B.n601 B.n32 585
R203 B.n600 B.n599 585
R204 B.n598 B.n33 585
R205 B.n597 B.n596 585
R206 B.n595 B.n34 585
R207 B.n594 B.n593 585
R208 B.n592 B.n35 585
R209 B.n591 B.n590 585
R210 B.n589 B.n36 585
R211 B.n588 B.n587 585
R212 B.n586 B.n37 585
R213 B.n585 B.n584 585
R214 B.n583 B.n38 585
R215 B.n582 B.n581 585
R216 B.n580 B.n39 585
R217 B.n579 B.n578 585
R218 B.n577 B.n40 585
R219 B.n576 B.n575 585
R220 B.n574 B.n41 585
R221 B.n573 B.n572 585
R222 B.n571 B.n570 585
R223 B.n569 B.n45 585
R224 B.n568 B.n567 585
R225 B.n566 B.n46 585
R226 B.n565 B.n564 585
R227 B.n563 B.n47 585
R228 B.n562 B.n561 585
R229 B.n560 B.n48 585
R230 B.n559 B.n558 585
R231 B.n556 B.n49 585
R232 B.n555 B.n554 585
R233 B.n553 B.n52 585
R234 B.n552 B.n551 585
R235 B.n550 B.n53 585
R236 B.n549 B.n548 585
R237 B.n547 B.n54 585
R238 B.n546 B.n545 585
R239 B.n544 B.n55 585
R240 B.n543 B.n542 585
R241 B.n541 B.n56 585
R242 B.n540 B.n539 585
R243 B.n538 B.n57 585
R244 B.n537 B.n536 585
R245 B.n535 B.n58 585
R246 B.n534 B.n533 585
R247 B.n532 B.n59 585
R248 B.n531 B.n530 585
R249 B.n529 B.n60 585
R250 B.n528 B.n527 585
R251 B.n526 B.n61 585
R252 B.n525 B.n524 585
R253 B.n523 B.n62 585
R254 B.n522 B.n521 585
R255 B.n520 B.n63 585
R256 B.n519 B.n518 585
R257 B.n517 B.n64 585
R258 B.n516 B.n515 585
R259 B.n514 B.n65 585
R260 B.n513 B.n512 585
R261 B.n511 B.n66 585
R262 B.n510 B.n509 585
R263 B.n508 B.n67 585
R264 B.n507 B.n506 585
R265 B.n505 B.n68 585
R266 B.n504 B.n503 585
R267 B.n502 B.n69 585
R268 B.n501 B.n500 585
R269 B.n499 B.n70 585
R270 B.n498 B.n497 585
R271 B.n496 B.n71 585
R272 B.n495 B.n494 585
R273 B.n493 B.n72 585
R274 B.n492 B.n491 585
R275 B.n490 B.n73 585
R276 B.n489 B.n488 585
R277 B.n487 B.n74 585
R278 B.n486 B.n485 585
R279 B.n484 B.n75 585
R280 B.n483 B.n482 585
R281 B.n481 B.n76 585
R282 B.n649 B.n16 585
R283 B.n651 B.n650 585
R284 B.n652 B.n15 585
R285 B.n654 B.n653 585
R286 B.n655 B.n14 585
R287 B.n657 B.n656 585
R288 B.n658 B.n13 585
R289 B.n660 B.n659 585
R290 B.n661 B.n12 585
R291 B.n663 B.n662 585
R292 B.n664 B.n11 585
R293 B.n666 B.n665 585
R294 B.n667 B.n10 585
R295 B.n669 B.n668 585
R296 B.n670 B.n9 585
R297 B.n672 B.n671 585
R298 B.n673 B.n8 585
R299 B.n675 B.n674 585
R300 B.n676 B.n7 585
R301 B.n678 B.n677 585
R302 B.n679 B.n6 585
R303 B.n681 B.n680 585
R304 B.n682 B.n5 585
R305 B.n684 B.n683 585
R306 B.n685 B.n4 585
R307 B.n687 B.n686 585
R308 B.n688 B.n3 585
R309 B.n690 B.n689 585
R310 B.n691 B.n0 585
R311 B.n2 B.n1 585
R312 B.n181 B.n180 585
R313 B.n183 B.n182 585
R314 B.n184 B.n179 585
R315 B.n186 B.n185 585
R316 B.n187 B.n178 585
R317 B.n189 B.n188 585
R318 B.n190 B.n177 585
R319 B.n192 B.n191 585
R320 B.n193 B.n176 585
R321 B.n195 B.n194 585
R322 B.n196 B.n175 585
R323 B.n198 B.n197 585
R324 B.n199 B.n174 585
R325 B.n201 B.n200 585
R326 B.n202 B.n173 585
R327 B.n204 B.n203 585
R328 B.n205 B.n172 585
R329 B.n207 B.n206 585
R330 B.n208 B.n171 585
R331 B.n210 B.n209 585
R332 B.n211 B.n170 585
R333 B.n213 B.n212 585
R334 B.n214 B.n169 585
R335 B.n216 B.n215 585
R336 B.n217 B.n168 585
R337 B.n219 B.n218 585
R338 B.n220 B.n167 585
R339 B.n222 B.n221 585
R340 B.n223 B.n222 511.721
R341 B.n391 B.n390 511.721
R342 B.n481 B.n480 511.721
R343 B.n649 B.n648 511.721
R344 B.n140 B.t3 452.063
R345 B.n132 B.t0 452.063
R346 B.n50 B.t9 452.063
R347 B.n42 B.t6 452.063
R348 B.n693 B.n692 256.663
R349 B.n692 B.n691 235.042
R350 B.n692 B.n2 235.042
R351 B.n224 B.n223 163.367
R352 B.n224 B.n165 163.367
R353 B.n228 B.n165 163.367
R354 B.n229 B.n228 163.367
R355 B.n230 B.n229 163.367
R356 B.n230 B.n163 163.367
R357 B.n234 B.n163 163.367
R358 B.n235 B.n234 163.367
R359 B.n236 B.n235 163.367
R360 B.n236 B.n161 163.367
R361 B.n240 B.n161 163.367
R362 B.n241 B.n240 163.367
R363 B.n242 B.n241 163.367
R364 B.n242 B.n159 163.367
R365 B.n246 B.n159 163.367
R366 B.n247 B.n246 163.367
R367 B.n248 B.n247 163.367
R368 B.n248 B.n157 163.367
R369 B.n252 B.n157 163.367
R370 B.n253 B.n252 163.367
R371 B.n254 B.n253 163.367
R372 B.n254 B.n155 163.367
R373 B.n258 B.n155 163.367
R374 B.n259 B.n258 163.367
R375 B.n260 B.n259 163.367
R376 B.n260 B.n153 163.367
R377 B.n264 B.n153 163.367
R378 B.n265 B.n264 163.367
R379 B.n266 B.n265 163.367
R380 B.n266 B.n151 163.367
R381 B.n270 B.n151 163.367
R382 B.n271 B.n270 163.367
R383 B.n272 B.n271 163.367
R384 B.n272 B.n149 163.367
R385 B.n276 B.n149 163.367
R386 B.n277 B.n276 163.367
R387 B.n278 B.n277 163.367
R388 B.n278 B.n147 163.367
R389 B.n282 B.n147 163.367
R390 B.n283 B.n282 163.367
R391 B.n284 B.n283 163.367
R392 B.n284 B.n145 163.367
R393 B.n288 B.n145 163.367
R394 B.n289 B.n288 163.367
R395 B.n290 B.n289 163.367
R396 B.n290 B.n143 163.367
R397 B.n294 B.n143 163.367
R398 B.n295 B.n294 163.367
R399 B.n296 B.n295 163.367
R400 B.n296 B.n139 163.367
R401 B.n301 B.n139 163.367
R402 B.n302 B.n301 163.367
R403 B.n303 B.n302 163.367
R404 B.n303 B.n137 163.367
R405 B.n307 B.n137 163.367
R406 B.n308 B.n307 163.367
R407 B.n309 B.n308 163.367
R408 B.n309 B.n135 163.367
R409 B.n313 B.n135 163.367
R410 B.n314 B.n313 163.367
R411 B.n314 B.n131 163.367
R412 B.n318 B.n131 163.367
R413 B.n319 B.n318 163.367
R414 B.n320 B.n319 163.367
R415 B.n320 B.n129 163.367
R416 B.n324 B.n129 163.367
R417 B.n325 B.n324 163.367
R418 B.n326 B.n325 163.367
R419 B.n326 B.n127 163.367
R420 B.n330 B.n127 163.367
R421 B.n331 B.n330 163.367
R422 B.n332 B.n331 163.367
R423 B.n332 B.n125 163.367
R424 B.n336 B.n125 163.367
R425 B.n337 B.n336 163.367
R426 B.n338 B.n337 163.367
R427 B.n338 B.n123 163.367
R428 B.n342 B.n123 163.367
R429 B.n343 B.n342 163.367
R430 B.n344 B.n343 163.367
R431 B.n344 B.n121 163.367
R432 B.n348 B.n121 163.367
R433 B.n349 B.n348 163.367
R434 B.n350 B.n349 163.367
R435 B.n350 B.n119 163.367
R436 B.n354 B.n119 163.367
R437 B.n355 B.n354 163.367
R438 B.n356 B.n355 163.367
R439 B.n356 B.n117 163.367
R440 B.n360 B.n117 163.367
R441 B.n361 B.n360 163.367
R442 B.n362 B.n361 163.367
R443 B.n362 B.n115 163.367
R444 B.n366 B.n115 163.367
R445 B.n367 B.n366 163.367
R446 B.n368 B.n367 163.367
R447 B.n368 B.n113 163.367
R448 B.n372 B.n113 163.367
R449 B.n373 B.n372 163.367
R450 B.n374 B.n373 163.367
R451 B.n374 B.n111 163.367
R452 B.n378 B.n111 163.367
R453 B.n379 B.n378 163.367
R454 B.n380 B.n379 163.367
R455 B.n380 B.n109 163.367
R456 B.n384 B.n109 163.367
R457 B.n385 B.n384 163.367
R458 B.n386 B.n385 163.367
R459 B.n386 B.n107 163.367
R460 B.n390 B.n107 163.367
R461 B.n480 B.n77 163.367
R462 B.n476 B.n77 163.367
R463 B.n476 B.n475 163.367
R464 B.n475 B.n474 163.367
R465 B.n474 B.n79 163.367
R466 B.n470 B.n79 163.367
R467 B.n470 B.n469 163.367
R468 B.n469 B.n468 163.367
R469 B.n468 B.n81 163.367
R470 B.n464 B.n81 163.367
R471 B.n464 B.n463 163.367
R472 B.n463 B.n462 163.367
R473 B.n462 B.n83 163.367
R474 B.n458 B.n83 163.367
R475 B.n458 B.n457 163.367
R476 B.n457 B.n456 163.367
R477 B.n456 B.n85 163.367
R478 B.n452 B.n85 163.367
R479 B.n452 B.n451 163.367
R480 B.n451 B.n450 163.367
R481 B.n450 B.n87 163.367
R482 B.n446 B.n87 163.367
R483 B.n446 B.n445 163.367
R484 B.n445 B.n444 163.367
R485 B.n444 B.n89 163.367
R486 B.n440 B.n89 163.367
R487 B.n440 B.n439 163.367
R488 B.n439 B.n438 163.367
R489 B.n438 B.n91 163.367
R490 B.n434 B.n91 163.367
R491 B.n434 B.n433 163.367
R492 B.n433 B.n432 163.367
R493 B.n432 B.n93 163.367
R494 B.n428 B.n93 163.367
R495 B.n428 B.n427 163.367
R496 B.n427 B.n426 163.367
R497 B.n426 B.n95 163.367
R498 B.n422 B.n95 163.367
R499 B.n422 B.n421 163.367
R500 B.n421 B.n420 163.367
R501 B.n420 B.n97 163.367
R502 B.n416 B.n97 163.367
R503 B.n416 B.n415 163.367
R504 B.n415 B.n414 163.367
R505 B.n414 B.n99 163.367
R506 B.n410 B.n99 163.367
R507 B.n410 B.n409 163.367
R508 B.n409 B.n408 163.367
R509 B.n408 B.n101 163.367
R510 B.n404 B.n101 163.367
R511 B.n404 B.n403 163.367
R512 B.n403 B.n402 163.367
R513 B.n402 B.n103 163.367
R514 B.n398 B.n103 163.367
R515 B.n398 B.n397 163.367
R516 B.n397 B.n396 163.367
R517 B.n396 B.n105 163.367
R518 B.n392 B.n105 163.367
R519 B.n392 B.n391 163.367
R520 B.n648 B.n17 163.367
R521 B.n644 B.n17 163.367
R522 B.n644 B.n643 163.367
R523 B.n643 B.n642 163.367
R524 B.n642 B.n19 163.367
R525 B.n638 B.n19 163.367
R526 B.n638 B.n637 163.367
R527 B.n637 B.n636 163.367
R528 B.n636 B.n21 163.367
R529 B.n632 B.n21 163.367
R530 B.n632 B.n631 163.367
R531 B.n631 B.n630 163.367
R532 B.n630 B.n23 163.367
R533 B.n626 B.n23 163.367
R534 B.n626 B.n625 163.367
R535 B.n625 B.n624 163.367
R536 B.n624 B.n25 163.367
R537 B.n620 B.n25 163.367
R538 B.n620 B.n619 163.367
R539 B.n619 B.n618 163.367
R540 B.n618 B.n27 163.367
R541 B.n614 B.n27 163.367
R542 B.n614 B.n613 163.367
R543 B.n613 B.n612 163.367
R544 B.n612 B.n29 163.367
R545 B.n608 B.n29 163.367
R546 B.n608 B.n607 163.367
R547 B.n607 B.n606 163.367
R548 B.n606 B.n31 163.367
R549 B.n602 B.n31 163.367
R550 B.n602 B.n601 163.367
R551 B.n601 B.n600 163.367
R552 B.n600 B.n33 163.367
R553 B.n596 B.n33 163.367
R554 B.n596 B.n595 163.367
R555 B.n595 B.n594 163.367
R556 B.n594 B.n35 163.367
R557 B.n590 B.n35 163.367
R558 B.n590 B.n589 163.367
R559 B.n589 B.n588 163.367
R560 B.n588 B.n37 163.367
R561 B.n584 B.n37 163.367
R562 B.n584 B.n583 163.367
R563 B.n583 B.n582 163.367
R564 B.n582 B.n39 163.367
R565 B.n578 B.n39 163.367
R566 B.n578 B.n577 163.367
R567 B.n577 B.n576 163.367
R568 B.n576 B.n41 163.367
R569 B.n572 B.n41 163.367
R570 B.n572 B.n571 163.367
R571 B.n571 B.n45 163.367
R572 B.n567 B.n45 163.367
R573 B.n567 B.n566 163.367
R574 B.n566 B.n565 163.367
R575 B.n565 B.n47 163.367
R576 B.n561 B.n47 163.367
R577 B.n561 B.n560 163.367
R578 B.n560 B.n559 163.367
R579 B.n559 B.n49 163.367
R580 B.n554 B.n49 163.367
R581 B.n554 B.n553 163.367
R582 B.n553 B.n552 163.367
R583 B.n552 B.n53 163.367
R584 B.n548 B.n53 163.367
R585 B.n548 B.n547 163.367
R586 B.n547 B.n546 163.367
R587 B.n546 B.n55 163.367
R588 B.n542 B.n55 163.367
R589 B.n542 B.n541 163.367
R590 B.n541 B.n540 163.367
R591 B.n540 B.n57 163.367
R592 B.n536 B.n57 163.367
R593 B.n536 B.n535 163.367
R594 B.n535 B.n534 163.367
R595 B.n534 B.n59 163.367
R596 B.n530 B.n59 163.367
R597 B.n530 B.n529 163.367
R598 B.n529 B.n528 163.367
R599 B.n528 B.n61 163.367
R600 B.n524 B.n61 163.367
R601 B.n524 B.n523 163.367
R602 B.n523 B.n522 163.367
R603 B.n522 B.n63 163.367
R604 B.n518 B.n63 163.367
R605 B.n518 B.n517 163.367
R606 B.n517 B.n516 163.367
R607 B.n516 B.n65 163.367
R608 B.n512 B.n65 163.367
R609 B.n512 B.n511 163.367
R610 B.n511 B.n510 163.367
R611 B.n510 B.n67 163.367
R612 B.n506 B.n67 163.367
R613 B.n506 B.n505 163.367
R614 B.n505 B.n504 163.367
R615 B.n504 B.n69 163.367
R616 B.n500 B.n69 163.367
R617 B.n500 B.n499 163.367
R618 B.n499 B.n498 163.367
R619 B.n498 B.n71 163.367
R620 B.n494 B.n71 163.367
R621 B.n494 B.n493 163.367
R622 B.n493 B.n492 163.367
R623 B.n492 B.n73 163.367
R624 B.n488 B.n73 163.367
R625 B.n488 B.n487 163.367
R626 B.n487 B.n486 163.367
R627 B.n486 B.n75 163.367
R628 B.n482 B.n75 163.367
R629 B.n482 B.n481 163.367
R630 B.n650 B.n649 163.367
R631 B.n650 B.n15 163.367
R632 B.n654 B.n15 163.367
R633 B.n655 B.n654 163.367
R634 B.n656 B.n655 163.367
R635 B.n656 B.n13 163.367
R636 B.n660 B.n13 163.367
R637 B.n661 B.n660 163.367
R638 B.n662 B.n661 163.367
R639 B.n662 B.n11 163.367
R640 B.n666 B.n11 163.367
R641 B.n667 B.n666 163.367
R642 B.n668 B.n667 163.367
R643 B.n668 B.n9 163.367
R644 B.n672 B.n9 163.367
R645 B.n673 B.n672 163.367
R646 B.n674 B.n673 163.367
R647 B.n674 B.n7 163.367
R648 B.n678 B.n7 163.367
R649 B.n679 B.n678 163.367
R650 B.n680 B.n679 163.367
R651 B.n680 B.n5 163.367
R652 B.n684 B.n5 163.367
R653 B.n685 B.n684 163.367
R654 B.n686 B.n685 163.367
R655 B.n686 B.n3 163.367
R656 B.n690 B.n3 163.367
R657 B.n691 B.n690 163.367
R658 B.n181 B.n2 163.367
R659 B.n182 B.n181 163.367
R660 B.n182 B.n179 163.367
R661 B.n186 B.n179 163.367
R662 B.n187 B.n186 163.367
R663 B.n188 B.n187 163.367
R664 B.n188 B.n177 163.367
R665 B.n192 B.n177 163.367
R666 B.n193 B.n192 163.367
R667 B.n194 B.n193 163.367
R668 B.n194 B.n175 163.367
R669 B.n198 B.n175 163.367
R670 B.n199 B.n198 163.367
R671 B.n200 B.n199 163.367
R672 B.n200 B.n173 163.367
R673 B.n204 B.n173 163.367
R674 B.n205 B.n204 163.367
R675 B.n206 B.n205 163.367
R676 B.n206 B.n171 163.367
R677 B.n210 B.n171 163.367
R678 B.n211 B.n210 163.367
R679 B.n212 B.n211 163.367
R680 B.n212 B.n169 163.367
R681 B.n216 B.n169 163.367
R682 B.n217 B.n216 163.367
R683 B.n218 B.n217 163.367
R684 B.n218 B.n167 163.367
R685 B.n222 B.n167 163.367
R686 B.n132 B.t1 145.327
R687 B.n50 B.t11 145.327
R688 B.n140 B.t4 145.309
R689 B.n42 B.t8 145.309
R690 B.n133 B.t2 110.225
R691 B.n51 B.t10 110.225
R692 B.n141 B.t5 110.206
R693 B.n43 B.t7 110.206
R694 B.n299 B.n141 59.5399
R695 B.n134 B.n133 59.5399
R696 B.n557 B.n51 59.5399
R697 B.n44 B.n43 59.5399
R698 B.n141 B.n140 35.1035
R699 B.n133 B.n132 35.1035
R700 B.n51 B.n50 35.1035
R701 B.n43 B.n42 35.1035
R702 B.n647 B.n16 33.2493
R703 B.n479 B.n76 33.2493
R704 B.n389 B.n106 33.2493
R705 B.n221 B.n166 33.2493
R706 B B.n693 18.0485
R707 B.n651 B.n16 10.6151
R708 B.n652 B.n651 10.6151
R709 B.n653 B.n652 10.6151
R710 B.n653 B.n14 10.6151
R711 B.n657 B.n14 10.6151
R712 B.n658 B.n657 10.6151
R713 B.n659 B.n658 10.6151
R714 B.n659 B.n12 10.6151
R715 B.n663 B.n12 10.6151
R716 B.n664 B.n663 10.6151
R717 B.n665 B.n664 10.6151
R718 B.n665 B.n10 10.6151
R719 B.n669 B.n10 10.6151
R720 B.n670 B.n669 10.6151
R721 B.n671 B.n670 10.6151
R722 B.n671 B.n8 10.6151
R723 B.n675 B.n8 10.6151
R724 B.n676 B.n675 10.6151
R725 B.n677 B.n676 10.6151
R726 B.n677 B.n6 10.6151
R727 B.n681 B.n6 10.6151
R728 B.n682 B.n681 10.6151
R729 B.n683 B.n682 10.6151
R730 B.n683 B.n4 10.6151
R731 B.n687 B.n4 10.6151
R732 B.n688 B.n687 10.6151
R733 B.n689 B.n688 10.6151
R734 B.n689 B.n0 10.6151
R735 B.n647 B.n646 10.6151
R736 B.n646 B.n645 10.6151
R737 B.n645 B.n18 10.6151
R738 B.n641 B.n18 10.6151
R739 B.n641 B.n640 10.6151
R740 B.n640 B.n639 10.6151
R741 B.n639 B.n20 10.6151
R742 B.n635 B.n20 10.6151
R743 B.n635 B.n634 10.6151
R744 B.n634 B.n633 10.6151
R745 B.n633 B.n22 10.6151
R746 B.n629 B.n22 10.6151
R747 B.n629 B.n628 10.6151
R748 B.n628 B.n627 10.6151
R749 B.n627 B.n24 10.6151
R750 B.n623 B.n24 10.6151
R751 B.n623 B.n622 10.6151
R752 B.n622 B.n621 10.6151
R753 B.n621 B.n26 10.6151
R754 B.n617 B.n26 10.6151
R755 B.n617 B.n616 10.6151
R756 B.n616 B.n615 10.6151
R757 B.n615 B.n28 10.6151
R758 B.n611 B.n28 10.6151
R759 B.n611 B.n610 10.6151
R760 B.n610 B.n609 10.6151
R761 B.n609 B.n30 10.6151
R762 B.n605 B.n30 10.6151
R763 B.n605 B.n604 10.6151
R764 B.n604 B.n603 10.6151
R765 B.n603 B.n32 10.6151
R766 B.n599 B.n32 10.6151
R767 B.n599 B.n598 10.6151
R768 B.n598 B.n597 10.6151
R769 B.n597 B.n34 10.6151
R770 B.n593 B.n34 10.6151
R771 B.n593 B.n592 10.6151
R772 B.n592 B.n591 10.6151
R773 B.n591 B.n36 10.6151
R774 B.n587 B.n36 10.6151
R775 B.n587 B.n586 10.6151
R776 B.n586 B.n585 10.6151
R777 B.n585 B.n38 10.6151
R778 B.n581 B.n38 10.6151
R779 B.n581 B.n580 10.6151
R780 B.n580 B.n579 10.6151
R781 B.n579 B.n40 10.6151
R782 B.n575 B.n40 10.6151
R783 B.n575 B.n574 10.6151
R784 B.n574 B.n573 10.6151
R785 B.n570 B.n569 10.6151
R786 B.n569 B.n568 10.6151
R787 B.n568 B.n46 10.6151
R788 B.n564 B.n46 10.6151
R789 B.n564 B.n563 10.6151
R790 B.n563 B.n562 10.6151
R791 B.n562 B.n48 10.6151
R792 B.n558 B.n48 10.6151
R793 B.n556 B.n555 10.6151
R794 B.n555 B.n52 10.6151
R795 B.n551 B.n52 10.6151
R796 B.n551 B.n550 10.6151
R797 B.n550 B.n549 10.6151
R798 B.n549 B.n54 10.6151
R799 B.n545 B.n54 10.6151
R800 B.n545 B.n544 10.6151
R801 B.n544 B.n543 10.6151
R802 B.n543 B.n56 10.6151
R803 B.n539 B.n56 10.6151
R804 B.n539 B.n538 10.6151
R805 B.n538 B.n537 10.6151
R806 B.n537 B.n58 10.6151
R807 B.n533 B.n58 10.6151
R808 B.n533 B.n532 10.6151
R809 B.n532 B.n531 10.6151
R810 B.n531 B.n60 10.6151
R811 B.n527 B.n60 10.6151
R812 B.n527 B.n526 10.6151
R813 B.n526 B.n525 10.6151
R814 B.n525 B.n62 10.6151
R815 B.n521 B.n62 10.6151
R816 B.n521 B.n520 10.6151
R817 B.n520 B.n519 10.6151
R818 B.n519 B.n64 10.6151
R819 B.n515 B.n64 10.6151
R820 B.n515 B.n514 10.6151
R821 B.n514 B.n513 10.6151
R822 B.n513 B.n66 10.6151
R823 B.n509 B.n66 10.6151
R824 B.n509 B.n508 10.6151
R825 B.n508 B.n507 10.6151
R826 B.n507 B.n68 10.6151
R827 B.n503 B.n68 10.6151
R828 B.n503 B.n502 10.6151
R829 B.n502 B.n501 10.6151
R830 B.n501 B.n70 10.6151
R831 B.n497 B.n70 10.6151
R832 B.n497 B.n496 10.6151
R833 B.n496 B.n495 10.6151
R834 B.n495 B.n72 10.6151
R835 B.n491 B.n72 10.6151
R836 B.n491 B.n490 10.6151
R837 B.n490 B.n489 10.6151
R838 B.n489 B.n74 10.6151
R839 B.n485 B.n74 10.6151
R840 B.n485 B.n484 10.6151
R841 B.n484 B.n483 10.6151
R842 B.n483 B.n76 10.6151
R843 B.n479 B.n478 10.6151
R844 B.n478 B.n477 10.6151
R845 B.n477 B.n78 10.6151
R846 B.n473 B.n78 10.6151
R847 B.n473 B.n472 10.6151
R848 B.n472 B.n471 10.6151
R849 B.n471 B.n80 10.6151
R850 B.n467 B.n80 10.6151
R851 B.n467 B.n466 10.6151
R852 B.n466 B.n465 10.6151
R853 B.n465 B.n82 10.6151
R854 B.n461 B.n82 10.6151
R855 B.n461 B.n460 10.6151
R856 B.n460 B.n459 10.6151
R857 B.n459 B.n84 10.6151
R858 B.n455 B.n84 10.6151
R859 B.n455 B.n454 10.6151
R860 B.n454 B.n453 10.6151
R861 B.n453 B.n86 10.6151
R862 B.n449 B.n86 10.6151
R863 B.n449 B.n448 10.6151
R864 B.n448 B.n447 10.6151
R865 B.n447 B.n88 10.6151
R866 B.n443 B.n88 10.6151
R867 B.n443 B.n442 10.6151
R868 B.n442 B.n441 10.6151
R869 B.n441 B.n90 10.6151
R870 B.n437 B.n90 10.6151
R871 B.n437 B.n436 10.6151
R872 B.n436 B.n435 10.6151
R873 B.n435 B.n92 10.6151
R874 B.n431 B.n92 10.6151
R875 B.n431 B.n430 10.6151
R876 B.n430 B.n429 10.6151
R877 B.n429 B.n94 10.6151
R878 B.n425 B.n94 10.6151
R879 B.n425 B.n424 10.6151
R880 B.n424 B.n423 10.6151
R881 B.n423 B.n96 10.6151
R882 B.n419 B.n96 10.6151
R883 B.n419 B.n418 10.6151
R884 B.n418 B.n417 10.6151
R885 B.n417 B.n98 10.6151
R886 B.n413 B.n98 10.6151
R887 B.n413 B.n412 10.6151
R888 B.n412 B.n411 10.6151
R889 B.n411 B.n100 10.6151
R890 B.n407 B.n100 10.6151
R891 B.n407 B.n406 10.6151
R892 B.n406 B.n405 10.6151
R893 B.n405 B.n102 10.6151
R894 B.n401 B.n102 10.6151
R895 B.n401 B.n400 10.6151
R896 B.n400 B.n399 10.6151
R897 B.n399 B.n104 10.6151
R898 B.n395 B.n104 10.6151
R899 B.n395 B.n394 10.6151
R900 B.n394 B.n393 10.6151
R901 B.n393 B.n106 10.6151
R902 B.n180 B.n1 10.6151
R903 B.n183 B.n180 10.6151
R904 B.n184 B.n183 10.6151
R905 B.n185 B.n184 10.6151
R906 B.n185 B.n178 10.6151
R907 B.n189 B.n178 10.6151
R908 B.n190 B.n189 10.6151
R909 B.n191 B.n190 10.6151
R910 B.n191 B.n176 10.6151
R911 B.n195 B.n176 10.6151
R912 B.n196 B.n195 10.6151
R913 B.n197 B.n196 10.6151
R914 B.n197 B.n174 10.6151
R915 B.n201 B.n174 10.6151
R916 B.n202 B.n201 10.6151
R917 B.n203 B.n202 10.6151
R918 B.n203 B.n172 10.6151
R919 B.n207 B.n172 10.6151
R920 B.n208 B.n207 10.6151
R921 B.n209 B.n208 10.6151
R922 B.n209 B.n170 10.6151
R923 B.n213 B.n170 10.6151
R924 B.n214 B.n213 10.6151
R925 B.n215 B.n214 10.6151
R926 B.n215 B.n168 10.6151
R927 B.n219 B.n168 10.6151
R928 B.n220 B.n219 10.6151
R929 B.n221 B.n220 10.6151
R930 B.n225 B.n166 10.6151
R931 B.n226 B.n225 10.6151
R932 B.n227 B.n226 10.6151
R933 B.n227 B.n164 10.6151
R934 B.n231 B.n164 10.6151
R935 B.n232 B.n231 10.6151
R936 B.n233 B.n232 10.6151
R937 B.n233 B.n162 10.6151
R938 B.n237 B.n162 10.6151
R939 B.n238 B.n237 10.6151
R940 B.n239 B.n238 10.6151
R941 B.n239 B.n160 10.6151
R942 B.n243 B.n160 10.6151
R943 B.n244 B.n243 10.6151
R944 B.n245 B.n244 10.6151
R945 B.n245 B.n158 10.6151
R946 B.n249 B.n158 10.6151
R947 B.n250 B.n249 10.6151
R948 B.n251 B.n250 10.6151
R949 B.n251 B.n156 10.6151
R950 B.n255 B.n156 10.6151
R951 B.n256 B.n255 10.6151
R952 B.n257 B.n256 10.6151
R953 B.n257 B.n154 10.6151
R954 B.n261 B.n154 10.6151
R955 B.n262 B.n261 10.6151
R956 B.n263 B.n262 10.6151
R957 B.n263 B.n152 10.6151
R958 B.n267 B.n152 10.6151
R959 B.n268 B.n267 10.6151
R960 B.n269 B.n268 10.6151
R961 B.n269 B.n150 10.6151
R962 B.n273 B.n150 10.6151
R963 B.n274 B.n273 10.6151
R964 B.n275 B.n274 10.6151
R965 B.n275 B.n148 10.6151
R966 B.n279 B.n148 10.6151
R967 B.n280 B.n279 10.6151
R968 B.n281 B.n280 10.6151
R969 B.n281 B.n146 10.6151
R970 B.n285 B.n146 10.6151
R971 B.n286 B.n285 10.6151
R972 B.n287 B.n286 10.6151
R973 B.n287 B.n144 10.6151
R974 B.n291 B.n144 10.6151
R975 B.n292 B.n291 10.6151
R976 B.n293 B.n292 10.6151
R977 B.n293 B.n142 10.6151
R978 B.n297 B.n142 10.6151
R979 B.n298 B.n297 10.6151
R980 B.n300 B.n138 10.6151
R981 B.n304 B.n138 10.6151
R982 B.n305 B.n304 10.6151
R983 B.n306 B.n305 10.6151
R984 B.n306 B.n136 10.6151
R985 B.n310 B.n136 10.6151
R986 B.n311 B.n310 10.6151
R987 B.n312 B.n311 10.6151
R988 B.n316 B.n315 10.6151
R989 B.n317 B.n316 10.6151
R990 B.n317 B.n130 10.6151
R991 B.n321 B.n130 10.6151
R992 B.n322 B.n321 10.6151
R993 B.n323 B.n322 10.6151
R994 B.n323 B.n128 10.6151
R995 B.n327 B.n128 10.6151
R996 B.n328 B.n327 10.6151
R997 B.n329 B.n328 10.6151
R998 B.n329 B.n126 10.6151
R999 B.n333 B.n126 10.6151
R1000 B.n334 B.n333 10.6151
R1001 B.n335 B.n334 10.6151
R1002 B.n335 B.n124 10.6151
R1003 B.n339 B.n124 10.6151
R1004 B.n340 B.n339 10.6151
R1005 B.n341 B.n340 10.6151
R1006 B.n341 B.n122 10.6151
R1007 B.n345 B.n122 10.6151
R1008 B.n346 B.n345 10.6151
R1009 B.n347 B.n346 10.6151
R1010 B.n347 B.n120 10.6151
R1011 B.n351 B.n120 10.6151
R1012 B.n352 B.n351 10.6151
R1013 B.n353 B.n352 10.6151
R1014 B.n353 B.n118 10.6151
R1015 B.n357 B.n118 10.6151
R1016 B.n358 B.n357 10.6151
R1017 B.n359 B.n358 10.6151
R1018 B.n359 B.n116 10.6151
R1019 B.n363 B.n116 10.6151
R1020 B.n364 B.n363 10.6151
R1021 B.n365 B.n364 10.6151
R1022 B.n365 B.n114 10.6151
R1023 B.n369 B.n114 10.6151
R1024 B.n370 B.n369 10.6151
R1025 B.n371 B.n370 10.6151
R1026 B.n371 B.n112 10.6151
R1027 B.n375 B.n112 10.6151
R1028 B.n376 B.n375 10.6151
R1029 B.n377 B.n376 10.6151
R1030 B.n377 B.n110 10.6151
R1031 B.n381 B.n110 10.6151
R1032 B.n382 B.n381 10.6151
R1033 B.n383 B.n382 10.6151
R1034 B.n383 B.n108 10.6151
R1035 B.n387 B.n108 10.6151
R1036 B.n388 B.n387 10.6151
R1037 B.n389 B.n388 10.6151
R1038 B.n693 B.n0 8.11757
R1039 B.n693 B.n1 8.11757
R1040 B.n570 B.n44 6.5566
R1041 B.n558 B.n557 6.5566
R1042 B.n300 B.n299 6.5566
R1043 B.n312 B.n134 6.5566
R1044 B.n573 B.n44 4.05904
R1045 B.n557 B.n556 4.05904
R1046 B.n299 B.n298 4.05904
R1047 B.n315 B.n134 4.05904
R1048 VN.n3 VN.t0 283.916
R1049 VN.n13 VN.t1 283.916
R1050 VN.n2 VN.t5 246.7
R1051 VN.n8 VN.t3 246.7
R1052 VN.n12 VN.t4 246.7
R1053 VN.n18 VN.t2 246.7
R1054 VN.n9 VN.n8 170.597
R1055 VN.n19 VN.n18 170.597
R1056 VN.n17 VN.n10 161.3
R1057 VN.n16 VN.n15 161.3
R1058 VN.n14 VN.n11 161.3
R1059 VN.n7 VN.n0 161.3
R1060 VN.n6 VN.n5 161.3
R1061 VN.n4 VN.n1 161.3
R1062 VN.n6 VN.n1 49.7204
R1063 VN.n16 VN.n11 49.7204
R1064 VN VN.n19 47.0516
R1065 VN.n3 VN.n2 41.8757
R1066 VN.n13 VN.n12 41.8757
R1067 VN.n7 VN.n6 31.2664
R1068 VN.n17 VN.n16 31.2664
R1069 VN.n2 VN.n1 24.4675
R1070 VN.n12 VN.n11 24.4675
R1071 VN.n14 VN.n13 17.226
R1072 VN.n4 VN.n3 17.226
R1073 VN.n8 VN.n7 15.17
R1074 VN.n18 VN.n17 15.17
R1075 VN.n19 VN.n10 0.189894
R1076 VN.n15 VN.n10 0.189894
R1077 VN.n15 VN.n14 0.189894
R1078 VN.n5 VN.n4 0.189894
R1079 VN.n5 VN.n0 0.189894
R1080 VN.n9 VN.n0 0.189894
R1081 VN VN.n9 0.0516364
R1082 VTAIL.n7 VTAIL.t6 58.881
R1083 VTAIL.n11 VTAIL.t7 58.8807
R1084 VTAIL.n2 VTAIL.t4 58.8807
R1085 VTAIL.n10 VTAIL.t1 58.8807
R1086 VTAIL.n9 VTAIL.n8 56.7355
R1087 VTAIL.n6 VTAIL.n5 56.7355
R1088 VTAIL.n1 VTAIL.n0 56.7352
R1089 VTAIL.n4 VTAIL.n3 56.7352
R1090 VTAIL.n6 VTAIL.n4 28.5479
R1091 VTAIL.n11 VTAIL.n10 26.9876
R1092 VTAIL.n0 VTAIL.t5 2.14604
R1093 VTAIL.n0 VTAIL.t10 2.14604
R1094 VTAIL.n3 VTAIL.t3 2.14604
R1095 VTAIL.n3 VTAIL.t11 2.14604
R1096 VTAIL.n8 VTAIL.t2 2.14604
R1097 VTAIL.n8 VTAIL.t0 2.14604
R1098 VTAIL.n5 VTAIL.t9 2.14604
R1099 VTAIL.n5 VTAIL.t8 2.14604
R1100 VTAIL.n7 VTAIL.n6 1.56084
R1101 VTAIL.n10 VTAIL.n9 1.56084
R1102 VTAIL.n4 VTAIL.n2 1.56084
R1103 VTAIL.n9 VTAIL.n7 1.2505
R1104 VTAIL.n2 VTAIL.n1 1.2505
R1105 VTAIL VTAIL.n11 1.11257
R1106 VTAIL VTAIL.n1 0.448776
R1107 VDD2.n1 VDD2.t5 76.6745
R1108 VDD2.n2 VDD2.t3 75.5598
R1109 VDD2.n1 VDD2.n0 73.7487
R1110 VDD2 VDD2.n3 73.746
R1111 VDD2.n2 VDD2.n1 41.8468
R1112 VDD2.n3 VDD2.t1 2.14604
R1113 VDD2.n3 VDD2.t4 2.14604
R1114 VDD2.n0 VDD2.t0 2.14604
R1115 VDD2.n0 VDD2.t2 2.14604
R1116 VDD2 VDD2.n2 1.22895
R1117 VP.n7 VP.t5 283.916
R1118 VP.n20 VP.t4 246.7
R1119 VP.n14 VP.t0 246.7
R1120 VP.n26 VP.t2 246.7
R1121 VP.n6 VP.t1 246.7
R1122 VP.n12 VP.t3 246.7
R1123 VP.n15 VP.n14 170.597
R1124 VP.n27 VP.n26 170.597
R1125 VP.n13 VP.n12 170.597
R1126 VP.n8 VP.n5 161.3
R1127 VP.n10 VP.n9 161.3
R1128 VP.n11 VP.n4 161.3
R1129 VP.n25 VP.n0 161.3
R1130 VP.n24 VP.n23 161.3
R1131 VP.n22 VP.n1 161.3
R1132 VP.n21 VP.n20 161.3
R1133 VP.n19 VP.n2 161.3
R1134 VP.n18 VP.n17 161.3
R1135 VP.n16 VP.n3 161.3
R1136 VP.n19 VP.n18 49.7204
R1137 VP.n24 VP.n1 49.7204
R1138 VP.n10 VP.n5 49.7204
R1139 VP.n15 VP.n13 46.671
R1140 VP.n7 VP.n6 41.8757
R1141 VP.n18 VP.n3 31.2664
R1142 VP.n25 VP.n24 31.2664
R1143 VP.n11 VP.n10 31.2664
R1144 VP.n20 VP.n19 24.4675
R1145 VP.n20 VP.n1 24.4675
R1146 VP.n6 VP.n5 24.4675
R1147 VP.n8 VP.n7 17.226
R1148 VP.n14 VP.n3 15.17
R1149 VP.n26 VP.n25 15.17
R1150 VP.n12 VP.n11 15.17
R1151 VP.n9 VP.n8 0.189894
R1152 VP.n9 VP.n4 0.189894
R1153 VP.n13 VP.n4 0.189894
R1154 VP.n16 VP.n15 0.189894
R1155 VP.n17 VP.n16 0.189894
R1156 VP.n17 VP.n2 0.189894
R1157 VP.n21 VP.n2 0.189894
R1158 VP.n22 VP.n21 0.189894
R1159 VP.n23 VP.n22 0.189894
R1160 VP.n23 VP.n0 0.189894
R1161 VP.n27 VP.n0 0.189894
R1162 VP VP.n27 0.0516364
R1163 VDD1 VDD1.t0 76.7883
R1164 VDD1.n1 VDD1.t5 76.6745
R1165 VDD1.n1 VDD1.n0 73.7487
R1166 VDD1.n3 VDD1.n2 73.4141
R1167 VDD1.n3 VDD1.n1 43.2099
R1168 VDD1.n2 VDD1.t4 2.14604
R1169 VDD1.n2 VDD1.t2 2.14604
R1170 VDD1.n0 VDD1.t1 2.14604
R1171 VDD1.n0 VDD1.t3 2.14604
R1172 VDD1 VDD1.n3 0.332397
C0 VN VDD1 0.149142f
C1 VTAIL VDD1 9.463861f
C2 VN VP 6.41818f
C3 VTAIL VP 7.08382f
C4 VDD2 VN 7.29712f
C5 VDD2 VTAIL 9.50429f
C6 B VN 0.967219f
C7 B VTAIL 3.80999f
C8 VDD1 w_n2418_n3998# 2.23936f
C9 VN VTAIL 7.06932f
C10 VP w_n2418_n3998# 4.67019f
C11 VDD2 w_n2418_n3998# 2.28836f
C12 B w_n2418_n3998# 9.01265f
C13 VN w_n2418_n3998# 4.3607f
C14 VTAIL w_n2418_n3998# 3.36649f
C15 VP VDD1 7.50725f
C16 VDD2 VDD1 0.999731f
C17 VDD2 VP 0.363784f
C18 B VDD1 2.02912f
C19 B VP 1.47831f
C20 VDD2 B 2.07648f
C21 VDD2 VSUBS 1.693967f
C22 VDD1 VSUBS 2.071727f
C23 VTAIL VSUBS 1.079337f
C24 VN VSUBS 5.04267f
C25 VP VSUBS 2.178005f
C26 B VSUBS 3.798458f
C27 w_n2418_n3998# VSUBS 0.11853p
C28 VDD1.t0 VSUBS 3.46932f
C29 VDD1.t5 VSUBS 3.46813f
C30 VDD1.t1 VSUBS 0.325971f
C31 VDD1.t3 VSUBS 0.325971f
C32 VDD1.n0 VSUBS 2.66343f
C33 VDD1.n1 VSUBS 3.54468f
C34 VDD1.t4 VSUBS 0.325971f
C35 VDD1.t2 VSUBS 0.325971f
C36 VDD1.n2 VSUBS 2.66029f
C37 VDD1.n3 VSUBS 3.24399f
C38 VP.n0 VSUBS 0.039877f
C39 VP.t2 VSUBS 2.45059f
C40 VP.n1 VSUBS 0.073574f
C41 VP.n2 VSUBS 0.039877f
C42 VP.t4 VSUBS 2.45059f
C43 VP.n3 VSUBS 0.066122f
C44 VP.n4 VSUBS 0.039877f
C45 VP.t3 VSUBS 2.45059f
C46 VP.n5 VSUBS 0.073574f
C47 VP.t5 VSUBS 2.58556f
C48 VP.t1 VSUBS 2.45059f
C49 VP.n6 VSUBS 0.965397f
C50 VP.n7 VSUBS 0.95285f
C51 VP.n8 VSUBS 0.254697f
C52 VP.n9 VSUBS 0.039877f
C53 VP.n10 VSUBS 0.037113f
C54 VP.n11 VSUBS 0.066122f
C55 VP.n12 VSUBS 0.962324f
C56 VP.n13 VSUBS 1.95607f
C57 VP.t0 VSUBS 2.45059f
C58 VP.n14 VSUBS 0.962324f
C59 VP.n15 VSUBS 1.98679f
C60 VP.n16 VSUBS 0.039877f
C61 VP.n17 VSUBS 0.039877f
C62 VP.n18 VSUBS 0.037113f
C63 VP.n19 VSUBS 0.073574f
C64 VP.n20 VSUBS 0.90956f
C65 VP.n21 VSUBS 0.039877f
C66 VP.n22 VSUBS 0.039877f
C67 VP.n23 VSUBS 0.039877f
C68 VP.n24 VSUBS 0.037113f
C69 VP.n25 VSUBS 0.066122f
C70 VP.n26 VSUBS 0.962324f
C71 VP.n27 VSUBS 0.036113f
C72 VDD2.t5 VSUBS 3.48466f
C73 VDD2.t0 VSUBS 0.327525f
C74 VDD2.t2 VSUBS 0.327525f
C75 VDD2.n0 VSUBS 2.67613f
C76 VDD2.n1 VSUBS 3.45509f
C77 VDD2.t3 VSUBS 3.47427f
C78 VDD2.n2 VSUBS 3.29833f
C79 VDD2.t1 VSUBS 0.327525f
C80 VDD2.t4 VSUBS 0.327525f
C81 VDD2.n3 VSUBS 2.67608f
C82 VTAIL.t5 VSUBS 0.332109f
C83 VTAIL.t10 VSUBS 0.332109f
C84 VTAIL.n0 VSUBS 2.559f
C85 VTAIL.n1 VSUBS 0.785752f
C86 VTAIL.t4 VSUBS 3.3506f
C87 VTAIL.n2 VSUBS 0.999306f
C88 VTAIL.t3 VSUBS 0.332109f
C89 VTAIL.t11 VSUBS 0.332109f
C90 VTAIL.n3 VSUBS 2.559f
C91 VTAIL.n4 VSUBS 2.59661f
C92 VTAIL.t9 VSUBS 0.332109f
C93 VTAIL.t8 VSUBS 0.332109f
C94 VTAIL.n5 VSUBS 2.55901f
C95 VTAIL.n6 VSUBS 2.5966f
C96 VTAIL.t6 VSUBS 3.35061f
C97 VTAIL.n7 VSUBS 0.999301f
C98 VTAIL.t2 VSUBS 0.332109f
C99 VTAIL.t0 VSUBS 0.332109f
C100 VTAIL.n8 VSUBS 2.55901f
C101 VTAIL.n9 VSUBS 0.885151f
C102 VTAIL.t1 VSUBS 3.3506f
C103 VTAIL.n10 VSUBS 2.57128f
C104 VTAIL.t7 VSUBS 3.3506f
C105 VTAIL.n11 VSUBS 2.53121f
C106 VN.n0 VSUBS 0.039016f
C107 VN.t3 VSUBS 2.39768f
C108 VN.n1 VSUBS 0.071986f
C109 VN.t0 VSUBS 2.52974f
C110 VN.t5 VSUBS 2.39768f
C111 VN.n2 VSUBS 0.944555f
C112 VN.n3 VSUBS 0.932279f
C113 VN.n4 VSUBS 0.249198f
C114 VN.n5 VSUBS 0.039016f
C115 VN.n6 VSUBS 0.036312f
C116 VN.n7 VSUBS 0.064694f
C117 VN.n8 VSUBS 0.941548f
C118 VN.n9 VSUBS 0.035333f
C119 VN.n10 VSUBS 0.039016f
C120 VN.t2 VSUBS 2.39768f
C121 VN.n11 VSUBS 0.071986f
C122 VN.t1 VSUBS 2.52974f
C123 VN.t4 VSUBS 2.39768f
C124 VN.n12 VSUBS 0.944555f
C125 VN.n13 VSUBS 0.932279f
C126 VN.n14 VSUBS 0.249198f
C127 VN.n15 VSUBS 0.039016f
C128 VN.n16 VSUBS 0.036312f
C129 VN.n17 VSUBS 0.064694f
C130 VN.n18 VSUBS 0.941548f
C131 VN.n19 VSUBS 1.9393f
C132 B.n0 VSUBS 0.007389f
C133 B.n1 VSUBS 0.007389f
C134 B.n2 VSUBS 0.010928f
C135 B.n3 VSUBS 0.008374f
C136 B.n4 VSUBS 0.008374f
C137 B.n5 VSUBS 0.008374f
C138 B.n6 VSUBS 0.008374f
C139 B.n7 VSUBS 0.008374f
C140 B.n8 VSUBS 0.008374f
C141 B.n9 VSUBS 0.008374f
C142 B.n10 VSUBS 0.008374f
C143 B.n11 VSUBS 0.008374f
C144 B.n12 VSUBS 0.008374f
C145 B.n13 VSUBS 0.008374f
C146 B.n14 VSUBS 0.008374f
C147 B.n15 VSUBS 0.008374f
C148 B.n16 VSUBS 0.019578f
C149 B.n17 VSUBS 0.008374f
C150 B.n18 VSUBS 0.008374f
C151 B.n19 VSUBS 0.008374f
C152 B.n20 VSUBS 0.008374f
C153 B.n21 VSUBS 0.008374f
C154 B.n22 VSUBS 0.008374f
C155 B.n23 VSUBS 0.008374f
C156 B.n24 VSUBS 0.008374f
C157 B.n25 VSUBS 0.008374f
C158 B.n26 VSUBS 0.008374f
C159 B.n27 VSUBS 0.008374f
C160 B.n28 VSUBS 0.008374f
C161 B.n29 VSUBS 0.008374f
C162 B.n30 VSUBS 0.008374f
C163 B.n31 VSUBS 0.008374f
C164 B.n32 VSUBS 0.008374f
C165 B.n33 VSUBS 0.008374f
C166 B.n34 VSUBS 0.008374f
C167 B.n35 VSUBS 0.008374f
C168 B.n36 VSUBS 0.008374f
C169 B.n37 VSUBS 0.008374f
C170 B.n38 VSUBS 0.008374f
C171 B.n39 VSUBS 0.008374f
C172 B.n40 VSUBS 0.008374f
C173 B.n41 VSUBS 0.008374f
C174 B.t7 VSUBS 0.603848f
C175 B.t8 VSUBS 0.620423f
C176 B.t6 VSUBS 1.15308f
C177 B.n42 VSUBS 0.270367f
C178 B.n43 VSUBS 0.080554f
C179 B.n44 VSUBS 0.019402f
C180 B.n45 VSUBS 0.008374f
C181 B.n46 VSUBS 0.008374f
C182 B.n47 VSUBS 0.008374f
C183 B.n48 VSUBS 0.008374f
C184 B.n49 VSUBS 0.008374f
C185 B.t10 VSUBS 0.603831f
C186 B.t11 VSUBS 0.620407f
C187 B.t9 VSUBS 1.15308f
C188 B.n50 VSUBS 0.270382f
C189 B.n51 VSUBS 0.080571f
C190 B.n52 VSUBS 0.008374f
C191 B.n53 VSUBS 0.008374f
C192 B.n54 VSUBS 0.008374f
C193 B.n55 VSUBS 0.008374f
C194 B.n56 VSUBS 0.008374f
C195 B.n57 VSUBS 0.008374f
C196 B.n58 VSUBS 0.008374f
C197 B.n59 VSUBS 0.008374f
C198 B.n60 VSUBS 0.008374f
C199 B.n61 VSUBS 0.008374f
C200 B.n62 VSUBS 0.008374f
C201 B.n63 VSUBS 0.008374f
C202 B.n64 VSUBS 0.008374f
C203 B.n65 VSUBS 0.008374f
C204 B.n66 VSUBS 0.008374f
C205 B.n67 VSUBS 0.008374f
C206 B.n68 VSUBS 0.008374f
C207 B.n69 VSUBS 0.008374f
C208 B.n70 VSUBS 0.008374f
C209 B.n71 VSUBS 0.008374f
C210 B.n72 VSUBS 0.008374f
C211 B.n73 VSUBS 0.008374f
C212 B.n74 VSUBS 0.008374f
C213 B.n75 VSUBS 0.008374f
C214 B.n76 VSUBS 0.020076f
C215 B.n77 VSUBS 0.008374f
C216 B.n78 VSUBS 0.008374f
C217 B.n79 VSUBS 0.008374f
C218 B.n80 VSUBS 0.008374f
C219 B.n81 VSUBS 0.008374f
C220 B.n82 VSUBS 0.008374f
C221 B.n83 VSUBS 0.008374f
C222 B.n84 VSUBS 0.008374f
C223 B.n85 VSUBS 0.008374f
C224 B.n86 VSUBS 0.008374f
C225 B.n87 VSUBS 0.008374f
C226 B.n88 VSUBS 0.008374f
C227 B.n89 VSUBS 0.008374f
C228 B.n90 VSUBS 0.008374f
C229 B.n91 VSUBS 0.008374f
C230 B.n92 VSUBS 0.008374f
C231 B.n93 VSUBS 0.008374f
C232 B.n94 VSUBS 0.008374f
C233 B.n95 VSUBS 0.008374f
C234 B.n96 VSUBS 0.008374f
C235 B.n97 VSUBS 0.008374f
C236 B.n98 VSUBS 0.008374f
C237 B.n99 VSUBS 0.008374f
C238 B.n100 VSUBS 0.008374f
C239 B.n101 VSUBS 0.008374f
C240 B.n102 VSUBS 0.008374f
C241 B.n103 VSUBS 0.008374f
C242 B.n104 VSUBS 0.008374f
C243 B.n105 VSUBS 0.008374f
C244 B.n106 VSUBS 0.02055f
C245 B.n107 VSUBS 0.008374f
C246 B.n108 VSUBS 0.008374f
C247 B.n109 VSUBS 0.008374f
C248 B.n110 VSUBS 0.008374f
C249 B.n111 VSUBS 0.008374f
C250 B.n112 VSUBS 0.008374f
C251 B.n113 VSUBS 0.008374f
C252 B.n114 VSUBS 0.008374f
C253 B.n115 VSUBS 0.008374f
C254 B.n116 VSUBS 0.008374f
C255 B.n117 VSUBS 0.008374f
C256 B.n118 VSUBS 0.008374f
C257 B.n119 VSUBS 0.008374f
C258 B.n120 VSUBS 0.008374f
C259 B.n121 VSUBS 0.008374f
C260 B.n122 VSUBS 0.008374f
C261 B.n123 VSUBS 0.008374f
C262 B.n124 VSUBS 0.008374f
C263 B.n125 VSUBS 0.008374f
C264 B.n126 VSUBS 0.008374f
C265 B.n127 VSUBS 0.008374f
C266 B.n128 VSUBS 0.008374f
C267 B.n129 VSUBS 0.008374f
C268 B.n130 VSUBS 0.008374f
C269 B.n131 VSUBS 0.008374f
C270 B.t2 VSUBS 0.603831f
C271 B.t1 VSUBS 0.620407f
C272 B.t0 VSUBS 1.15308f
C273 B.n132 VSUBS 0.270382f
C274 B.n133 VSUBS 0.080571f
C275 B.n134 VSUBS 0.019402f
C276 B.n135 VSUBS 0.008374f
C277 B.n136 VSUBS 0.008374f
C278 B.n137 VSUBS 0.008374f
C279 B.n138 VSUBS 0.008374f
C280 B.n139 VSUBS 0.008374f
C281 B.t5 VSUBS 0.603848f
C282 B.t4 VSUBS 0.620423f
C283 B.t3 VSUBS 1.15308f
C284 B.n140 VSUBS 0.270367f
C285 B.n141 VSUBS 0.080554f
C286 B.n142 VSUBS 0.008374f
C287 B.n143 VSUBS 0.008374f
C288 B.n144 VSUBS 0.008374f
C289 B.n145 VSUBS 0.008374f
C290 B.n146 VSUBS 0.008374f
C291 B.n147 VSUBS 0.008374f
C292 B.n148 VSUBS 0.008374f
C293 B.n149 VSUBS 0.008374f
C294 B.n150 VSUBS 0.008374f
C295 B.n151 VSUBS 0.008374f
C296 B.n152 VSUBS 0.008374f
C297 B.n153 VSUBS 0.008374f
C298 B.n154 VSUBS 0.008374f
C299 B.n155 VSUBS 0.008374f
C300 B.n156 VSUBS 0.008374f
C301 B.n157 VSUBS 0.008374f
C302 B.n158 VSUBS 0.008374f
C303 B.n159 VSUBS 0.008374f
C304 B.n160 VSUBS 0.008374f
C305 B.n161 VSUBS 0.008374f
C306 B.n162 VSUBS 0.008374f
C307 B.n163 VSUBS 0.008374f
C308 B.n164 VSUBS 0.008374f
C309 B.n165 VSUBS 0.008374f
C310 B.n166 VSUBS 0.020076f
C311 B.n167 VSUBS 0.008374f
C312 B.n168 VSUBS 0.008374f
C313 B.n169 VSUBS 0.008374f
C314 B.n170 VSUBS 0.008374f
C315 B.n171 VSUBS 0.008374f
C316 B.n172 VSUBS 0.008374f
C317 B.n173 VSUBS 0.008374f
C318 B.n174 VSUBS 0.008374f
C319 B.n175 VSUBS 0.008374f
C320 B.n176 VSUBS 0.008374f
C321 B.n177 VSUBS 0.008374f
C322 B.n178 VSUBS 0.008374f
C323 B.n179 VSUBS 0.008374f
C324 B.n180 VSUBS 0.008374f
C325 B.n181 VSUBS 0.008374f
C326 B.n182 VSUBS 0.008374f
C327 B.n183 VSUBS 0.008374f
C328 B.n184 VSUBS 0.008374f
C329 B.n185 VSUBS 0.008374f
C330 B.n186 VSUBS 0.008374f
C331 B.n187 VSUBS 0.008374f
C332 B.n188 VSUBS 0.008374f
C333 B.n189 VSUBS 0.008374f
C334 B.n190 VSUBS 0.008374f
C335 B.n191 VSUBS 0.008374f
C336 B.n192 VSUBS 0.008374f
C337 B.n193 VSUBS 0.008374f
C338 B.n194 VSUBS 0.008374f
C339 B.n195 VSUBS 0.008374f
C340 B.n196 VSUBS 0.008374f
C341 B.n197 VSUBS 0.008374f
C342 B.n198 VSUBS 0.008374f
C343 B.n199 VSUBS 0.008374f
C344 B.n200 VSUBS 0.008374f
C345 B.n201 VSUBS 0.008374f
C346 B.n202 VSUBS 0.008374f
C347 B.n203 VSUBS 0.008374f
C348 B.n204 VSUBS 0.008374f
C349 B.n205 VSUBS 0.008374f
C350 B.n206 VSUBS 0.008374f
C351 B.n207 VSUBS 0.008374f
C352 B.n208 VSUBS 0.008374f
C353 B.n209 VSUBS 0.008374f
C354 B.n210 VSUBS 0.008374f
C355 B.n211 VSUBS 0.008374f
C356 B.n212 VSUBS 0.008374f
C357 B.n213 VSUBS 0.008374f
C358 B.n214 VSUBS 0.008374f
C359 B.n215 VSUBS 0.008374f
C360 B.n216 VSUBS 0.008374f
C361 B.n217 VSUBS 0.008374f
C362 B.n218 VSUBS 0.008374f
C363 B.n219 VSUBS 0.008374f
C364 B.n220 VSUBS 0.008374f
C365 B.n221 VSUBS 0.019578f
C366 B.n222 VSUBS 0.019578f
C367 B.n223 VSUBS 0.020076f
C368 B.n224 VSUBS 0.008374f
C369 B.n225 VSUBS 0.008374f
C370 B.n226 VSUBS 0.008374f
C371 B.n227 VSUBS 0.008374f
C372 B.n228 VSUBS 0.008374f
C373 B.n229 VSUBS 0.008374f
C374 B.n230 VSUBS 0.008374f
C375 B.n231 VSUBS 0.008374f
C376 B.n232 VSUBS 0.008374f
C377 B.n233 VSUBS 0.008374f
C378 B.n234 VSUBS 0.008374f
C379 B.n235 VSUBS 0.008374f
C380 B.n236 VSUBS 0.008374f
C381 B.n237 VSUBS 0.008374f
C382 B.n238 VSUBS 0.008374f
C383 B.n239 VSUBS 0.008374f
C384 B.n240 VSUBS 0.008374f
C385 B.n241 VSUBS 0.008374f
C386 B.n242 VSUBS 0.008374f
C387 B.n243 VSUBS 0.008374f
C388 B.n244 VSUBS 0.008374f
C389 B.n245 VSUBS 0.008374f
C390 B.n246 VSUBS 0.008374f
C391 B.n247 VSUBS 0.008374f
C392 B.n248 VSUBS 0.008374f
C393 B.n249 VSUBS 0.008374f
C394 B.n250 VSUBS 0.008374f
C395 B.n251 VSUBS 0.008374f
C396 B.n252 VSUBS 0.008374f
C397 B.n253 VSUBS 0.008374f
C398 B.n254 VSUBS 0.008374f
C399 B.n255 VSUBS 0.008374f
C400 B.n256 VSUBS 0.008374f
C401 B.n257 VSUBS 0.008374f
C402 B.n258 VSUBS 0.008374f
C403 B.n259 VSUBS 0.008374f
C404 B.n260 VSUBS 0.008374f
C405 B.n261 VSUBS 0.008374f
C406 B.n262 VSUBS 0.008374f
C407 B.n263 VSUBS 0.008374f
C408 B.n264 VSUBS 0.008374f
C409 B.n265 VSUBS 0.008374f
C410 B.n266 VSUBS 0.008374f
C411 B.n267 VSUBS 0.008374f
C412 B.n268 VSUBS 0.008374f
C413 B.n269 VSUBS 0.008374f
C414 B.n270 VSUBS 0.008374f
C415 B.n271 VSUBS 0.008374f
C416 B.n272 VSUBS 0.008374f
C417 B.n273 VSUBS 0.008374f
C418 B.n274 VSUBS 0.008374f
C419 B.n275 VSUBS 0.008374f
C420 B.n276 VSUBS 0.008374f
C421 B.n277 VSUBS 0.008374f
C422 B.n278 VSUBS 0.008374f
C423 B.n279 VSUBS 0.008374f
C424 B.n280 VSUBS 0.008374f
C425 B.n281 VSUBS 0.008374f
C426 B.n282 VSUBS 0.008374f
C427 B.n283 VSUBS 0.008374f
C428 B.n284 VSUBS 0.008374f
C429 B.n285 VSUBS 0.008374f
C430 B.n286 VSUBS 0.008374f
C431 B.n287 VSUBS 0.008374f
C432 B.n288 VSUBS 0.008374f
C433 B.n289 VSUBS 0.008374f
C434 B.n290 VSUBS 0.008374f
C435 B.n291 VSUBS 0.008374f
C436 B.n292 VSUBS 0.008374f
C437 B.n293 VSUBS 0.008374f
C438 B.n294 VSUBS 0.008374f
C439 B.n295 VSUBS 0.008374f
C440 B.n296 VSUBS 0.008374f
C441 B.n297 VSUBS 0.008374f
C442 B.n298 VSUBS 0.005788f
C443 B.n299 VSUBS 0.019402f
C444 B.n300 VSUBS 0.006773f
C445 B.n301 VSUBS 0.008374f
C446 B.n302 VSUBS 0.008374f
C447 B.n303 VSUBS 0.008374f
C448 B.n304 VSUBS 0.008374f
C449 B.n305 VSUBS 0.008374f
C450 B.n306 VSUBS 0.008374f
C451 B.n307 VSUBS 0.008374f
C452 B.n308 VSUBS 0.008374f
C453 B.n309 VSUBS 0.008374f
C454 B.n310 VSUBS 0.008374f
C455 B.n311 VSUBS 0.008374f
C456 B.n312 VSUBS 0.006773f
C457 B.n313 VSUBS 0.008374f
C458 B.n314 VSUBS 0.008374f
C459 B.n315 VSUBS 0.005788f
C460 B.n316 VSUBS 0.008374f
C461 B.n317 VSUBS 0.008374f
C462 B.n318 VSUBS 0.008374f
C463 B.n319 VSUBS 0.008374f
C464 B.n320 VSUBS 0.008374f
C465 B.n321 VSUBS 0.008374f
C466 B.n322 VSUBS 0.008374f
C467 B.n323 VSUBS 0.008374f
C468 B.n324 VSUBS 0.008374f
C469 B.n325 VSUBS 0.008374f
C470 B.n326 VSUBS 0.008374f
C471 B.n327 VSUBS 0.008374f
C472 B.n328 VSUBS 0.008374f
C473 B.n329 VSUBS 0.008374f
C474 B.n330 VSUBS 0.008374f
C475 B.n331 VSUBS 0.008374f
C476 B.n332 VSUBS 0.008374f
C477 B.n333 VSUBS 0.008374f
C478 B.n334 VSUBS 0.008374f
C479 B.n335 VSUBS 0.008374f
C480 B.n336 VSUBS 0.008374f
C481 B.n337 VSUBS 0.008374f
C482 B.n338 VSUBS 0.008374f
C483 B.n339 VSUBS 0.008374f
C484 B.n340 VSUBS 0.008374f
C485 B.n341 VSUBS 0.008374f
C486 B.n342 VSUBS 0.008374f
C487 B.n343 VSUBS 0.008374f
C488 B.n344 VSUBS 0.008374f
C489 B.n345 VSUBS 0.008374f
C490 B.n346 VSUBS 0.008374f
C491 B.n347 VSUBS 0.008374f
C492 B.n348 VSUBS 0.008374f
C493 B.n349 VSUBS 0.008374f
C494 B.n350 VSUBS 0.008374f
C495 B.n351 VSUBS 0.008374f
C496 B.n352 VSUBS 0.008374f
C497 B.n353 VSUBS 0.008374f
C498 B.n354 VSUBS 0.008374f
C499 B.n355 VSUBS 0.008374f
C500 B.n356 VSUBS 0.008374f
C501 B.n357 VSUBS 0.008374f
C502 B.n358 VSUBS 0.008374f
C503 B.n359 VSUBS 0.008374f
C504 B.n360 VSUBS 0.008374f
C505 B.n361 VSUBS 0.008374f
C506 B.n362 VSUBS 0.008374f
C507 B.n363 VSUBS 0.008374f
C508 B.n364 VSUBS 0.008374f
C509 B.n365 VSUBS 0.008374f
C510 B.n366 VSUBS 0.008374f
C511 B.n367 VSUBS 0.008374f
C512 B.n368 VSUBS 0.008374f
C513 B.n369 VSUBS 0.008374f
C514 B.n370 VSUBS 0.008374f
C515 B.n371 VSUBS 0.008374f
C516 B.n372 VSUBS 0.008374f
C517 B.n373 VSUBS 0.008374f
C518 B.n374 VSUBS 0.008374f
C519 B.n375 VSUBS 0.008374f
C520 B.n376 VSUBS 0.008374f
C521 B.n377 VSUBS 0.008374f
C522 B.n378 VSUBS 0.008374f
C523 B.n379 VSUBS 0.008374f
C524 B.n380 VSUBS 0.008374f
C525 B.n381 VSUBS 0.008374f
C526 B.n382 VSUBS 0.008374f
C527 B.n383 VSUBS 0.008374f
C528 B.n384 VSUBS 0.008374f
C529 B.n385 VSUBS 0.008374f
C530 B.n386 VSUBS 0.008374f
C531 B.n387 VSUBS 0.008374f
C532 B.n388 VSUBS 0.008374f
C533 B.n389 VSUBS 0.019104f
C534 B.n390 VSUBS 0.020076f
C535 B.n391 VSUBS 0.019578f
C536 B.n392 VSUBS 0.008374f
C537 B.n393 VSUBS 0.008374f
C538 B.n394 VSUBS 0.008374f
C539 B.n395 VSUBS 0.008374f
C540 B.n396 VSUBS 0.008374f
C541 B.n397 VSUBS 0.008374f
C542 B.n398 VSUBS 0.008374f
C543 B.n399 VSUBS 0.008374f
C544 B.n400 VSUBS 0.008374f
C545 B.n401 VSUBS 0.008374f
C546 B.n402 VSUBS 0.008374f
C547 B.n403 VSUBS 0.008374f
C548 B.n404 VSUBS 0.008374f
C549 B.n405 VSUBS 0.008374f
C550 B.n406 VSUBS 0.008374f
C551 B.n407 VSUBS 0.008374f
C552 B.n408 VSUBS 0.008374f
C553 B.n409 VSUBS 0.008374f
C554 B.n410 VSUBS 0.008374f
C555 B.n411 VSUBS 0.008374f
C556 B.n412 VSUBS 0.008374f
C557 B.n413 VSUBS 0.008374f
C558 B.n414 VSUBS 0.008374f
C559 B.n415 VSUBS 0.008374f
C560 B.n416 VSUBS 0.008374f
C561 B.n417 VSUBS 0.008374f
C562 B.n418 VSUBS 0.008374f
C563 B.n419 VSUBS 0.008374f
C564 B.n420 VSUBS 0.008374f
C565 B.n421 VSUBS 0.008374f
C566 B.n422 VSUBS 0.008374f
C567 B.n423 VSUBS 0.008374f
C568 B.n424 VSUBS 0.008374f
C569 B.n425 VSUBS 0.008374f
C570 B.n426 VSUBS 0.008374f
C571 B.n427 VSUBS 0.008374f
C572 B.n428 VSUBS 0.008374f
C573 B.n429 VSUBS 0.008374f
C574 B.n430 VSUBS 0.008374f
C575 B.n431 VSUBS 0.008374f
C576 B.n432 VSUBS 0.008374f
C577 B.n433 VSUBS 0.008374f
C578 B.n434 VSUBS 0.008374f
C579 B.n435 VSUBS 0.008374f
C580 B.n436 VSUBS 0.008374f
C581 B.n437 VSUBS 0.008374f
C582 B.n438 VSUBS 0.008374f
C583 B.n439 VSUBS 0.008374f
C584 B.n440 VSUBS 0.008374f
C585 B.n441 VSUBS 0.008374f
C586 B.n442 VSUBS 0.008374f
C587 B.n443 VSUBS 0.008374f
C588 B.n444 VSUBS 0.008374f
C589 B.n445 VSUBS 0.008374f
C590 B.n446 VSUBS 0.008374f
C591 B.n447 VSUBS 0.008374f
C592 B.n448 VSUBS 0.008374f
C593 B.n449 VSUBS 0.008374f
C594 B.n450 VSUBS 0.008374f
C595 B.n451 VSUBS 0.008374f
C596 B.n452 VSUBS 0.008374f
C597 B.n453 VSUBS 0.008374f
C598 B.n454 VSUBS 0.008374f
C599 B.n455 VSUBS 0.008374f
C600 B.n456 VSUBS 0.008374f
C601 B.n457 VSUBS 0.008374f
C602 B.n458 VSUBS 0.008374f
C603 B.n459 VSUBS 0.008374f
C604 B.n460 VSUBS 0.008374f
C605 B.n461 VSUBS 0.008374f
C606 B.n462 VSUBS 0.008374f
C607 B.n463 VSUBS 0.008374f
C608 B.n464 VSUBS 0.008374f
C609 B.n465 VSUBS 0.008374f
C610 B.n466 VSUBS 0.008374f
C611 B.n467 VSUBS 0.008374f
C612 B.n468 VSUBS 0.008374f
C613 B.n469 VSUBS 0.008374f
C614 B.n470 VSUBS 0.008374f
C615 B.n471 VSUBS 0.008374f
C616 B.n472 VSUBS 0.008374f
C617 B.n473 VSUBS 0.008374f
C618 B.n474 VSUBS 0.008374f
C619 B.n475 VSUBS 0.008374f
C620 B.n476 VSUBS 0.008374f
C621 B.n477 VSUBS 0.008374f
C622 B.n478 VSUBS 0.008374f
C623 B.n479 VSUBS 0.019578f
C624 B.n480 VSUBS 0.019578f
C625 B.n481 VSUBS 0.020076f
C626 B.n482 VSUBS 0.008374f
C627 B.n483 VSUBS 0.008374f
C628 B.n484 VSUBS 0.008374f
C629 B.n485 VSUBS 0.008374f
C630 B.n486 VSUBS 0.008374f
C631 B.n487 VSUBS 0.008374f
C632 B.n488 VSUBS 0.008374f
C633 B.n489 VSUBS 0.008374f
C634 B.n490 VSUBS 0.008374f
C635 B.n491 VSUBS 0.008374f
C636 B.n492 VSUBS 0.008374f
C637 B.n493 VSUBS 0.008374f
C638 B.n494 VSUBS 0.008374f
C639 B.n495 VSUBS 0.008374f
C640 B.n496 VSUBS 0.008374f
C641 B.n497 VSUBS 0.008374f
C642 B.n498 VSUBS 0.008374f
C643 B.n499 VSUBS 0.008374f
C644 B.n500 VSUBS 0.008374f
C645 B.n501 VSUBS 0.008374f
C646 B.n502 VSUBS 0.008374f
C647 B.n503 VSUBS 0.008374f
C648 B.n504 VSUBS 0.008374f
C649 B.n505 VSUBS 0.008374f
C650 B.n506 VSUBS 0.008374f
C651 B.n507 VSUBS 0.008374f
C652 B.n508 VSUBS 0.008374f
C653 B.n509 VSUBS 0.008374f
C654 B.n510 VSUBS 0.008374f
C655 B.n511 VSUBS 0.008374f
C656 B.n512 VSUBS 0.008374f
C657 B.n513 VSUBS 0.008374f
C658 B.n514 VSUBS 0.008374f
C659 B.n515 VSUBS 0.008374f
C660 B.n516 VSUBS 0.008374f
C661 B.n517 VSUBS 0.008374f
C662 B.n518 VSUBS 0.008374f
C663 B.n519 VSUBS 0.008374f
C664 B.n520 VSUBS 0.008374f
C665 B.n521 VSUBS 0.008374f
C666 B.n522 VSUBS 0.008374f
C667 B.n523 VSUBS 0.008374f
C668 B.n524 VSUBS 0.008374f
C669 B.n525 VSUBS 0.008374f
C670 B.n526 VSUBS 0.008374f
C671 B.n527 VSUBS 0.008374f
C672 B.n528 VSUBS 0.008374f
C673 B.n529 VSUBS 0.008374f
C674 B.n530 VSUBS 0.008374f
C675 B.n531 VSUBS 0.008374f
C676 B.n532 VSUBS 0.008374f
C677 B.n533 VSUBS 0.008374f
C678 B.n534 VSUBS 0.008374f
C679 B.n535 VSUBS 0.008374f
C680 B.n536 VSUBS 0.008374f
C681 B.n537 VSUBS 0.008374f
C682 B.n538 VSUBS 0.008374f
C683 B.n539 VSUBS 0.008374f
C684 B.n540 VSUBS 0.008374f
C685 B.n541 VSUBS 0.008374f
C686 B.n542 VSUBS 0.008374f
C687 B.n543 VSUBS 0.008374f
C688 B.n544 VSUBS 0.008374f
C689 B.n545 VSUBS 0.008374f
C690 B.n546 VSUBS 0.008374f
C691 B.n547 VSUBS 0.008374f
C692 B.n548 VSUBS 0.008374f
C693 B.n549 VSUBS 0.008374f
C694 B.n550 VSUBS 0.008374f
C695 B.n551 VSUBS 0.008374f
C696 B.n552 VSUBS 0.008374f
C697 B.n553 VSUBS 0.008374f
C698 B.n554 VSUBS 0.008374f
C699 B.n555 VSUBS 0.008374f
C700 B.n556 VSUBS 0.005788f
C701 B.n557 VSUBS 0.019402f
C702 B.n558 VSUBS 0.006773f
C703 B.n559 VSUBS 0.008374f
C704 B.n560 VSUBS 0.008374f
C705 B.n561 VSUBS 0.008374f
C706 B.n562 VSUBS 0.008374f
C707 B.n563 VSUBS 0.008374f
C708 B.n564 VSUBS 0.008374f
C709 B.n565 VSUBS 0.008374f
C710 B.n566 VSUBS 0.008374f
C711 B.n567 VSUBS 0.008374f
C712 B.n568 VSUBS 0.008374f
C713 B.n569 VSUBS 0.008374f
C714 B.n570 VSUBS 0.006773f
C715 B.n571 VSUBS 0.008374f
C716 B.n572 VSUBS 0.008374f
C717 B.n573 VSUBS 0.005788f
C718 B.n574 VSUBS 0.008374f
C719 B.n575 VSUBS 0.008374f
C720 B.n576 VSUBS 0.008374f
C721 B.n577 VSUBS 0.008374f
C722 B.n578 VSUBS 0.008374f
C723 B.n579 VSUBS 0.008374f
C724 B.n580 VSUBS 0.008374f
C725 B.n581 VSUBS 0.008374f
C726 B.n582 VSUBS 0.008374f
C727 B.n583 VSUBS 0.008374f
C728 B.n584 VSUBS 0.008374f
C729 B.n585 VSUBS 0.008374f
C730 B.n586 VSUBS 0.008374f
C731 B.n587 VSUBS 0.008374f
C732 B.n588 VSUBS 0.008374f
C733 B.n589 VSUBS 0.008374f
C734 B.n590 VSUBS 0.008374f
C735 B.n591 VSUBS 0.008374f
C736 B.n592 VSUBS 0.008374f
C737 B.n593 VSUBS 0.008374f
C738 B.n594 VSUBS 0.008374f
C739 B.n595 VSUBS 0.008374f
C740 B.n596 VSUBS 0.008374f
C741 B.n597 VSUBS 0.008374f
C742 B.n598 VSUBS 0.008374f
C743 B.n599 VSUBS 0.008374f
C744 B.n600 VSUBS 0.008374f
C745 B.n601 VSUBS 0.008374f
C746 B.n602 VSUBS 0.008374f
C747 B.n603 VSUBS 0.008374f
C748 B.n604 VSUBS 0.008374f
C749 B.n605 VSUBS 0.008374f
C750 B.n606 VSUBS 0.008374f
C751 B.n607 VSUBS 0.008374f
C752 B.n608 VSUBS 0.008374f
C753 B.n609 VSUBS 0.008374f
C754 B.n610 VSUBS 0.008374f
C755 B.n611 VSUBS 0.008374f
C756 B.n612 VSUBS 0.008374f
C757 B.n613 VSUBS 0.008374f
C758 B.n614 VSUBS 0.008374f
C759 B.n615 VSUBS 0.008374f
C760 B.n616 VSUBS 0.008374f
C761 B.n617 VSUBS 0.008374f
C762 B.n618 VSUBS 0.008374f
C763 B.n619 VSUBS 0.008374f
C764 B.n620 VSUBS 0.008374f
C765 B.n621 VSUBS 0.008374f
C766 B.n622 VSUBS 0.008374f
C767 B.n623 VSUBS 0.008374f
C768 B.n624 VSUBS 0.008374f
C769 B.n625 VSUBS 0.008374f
C770 B.n626 VSUBS 0.008374f
C771 B.n627 VSUBS 0.008374f
C772 B.n628 VSUBS 0.008374f
C773 B.n629 VSUBS 0.008374f
C774 B.n630 VSUBS 0.008374f
C775 B.n631 VSUBS 0.008374f
C776 B.n632 VSUBS 0.008374f
C777 B.n633 VSUBS 0.008374f
C778 B.n634 VSUBS 0.008374f
C779 B.n635 VSUBS 0.008374f
C780 B.n636 VSUBS 0.008374f
C781 B.n637 VSUBS 0.008374f
C782 B.n638 VSUBS 0.008374f
C783 B.n639 VSUBS 0.008374f
C784 B.n640 VSUBS 0.008374f
C785 B.n641 VSUBS 0.008374f
C786 B.n642 VSUBS 0.008374f
C787 B.n643 VSUBS 0.008374f
C788 B.n644 VSUBS 0.008374f
C789 B.n645 VSUBS 0.008374f
C790 B.n646 VSUBS 0.008374f
C791 B.n647 VSUBS 0.020076f
C792 B.n648 VSUBS 0.020076f
C793 B.n649 VSUBS 0.019578f
C794 B.n650 VSUBS 0.008374f
C795 B.n651 VSUBS 0.008374f
C796 B.n652 VSUBS 0.008374f
C797 B.n653 VSUBS 0.008374f
C798 B.n654 VSUBS 0.008374f
C799 B.n655 VSUBS 0.008374f
C800 B.n656 VSUBS 0.008374f
C801 B.n657 VSUBS 0.008374f
C802 B.n658 VSUBS 0.008374f
C803 B.n659 VSUBS 0.008374f
C804 B.n660 VSUBS 0.008374f
C805 B.n661 VSUBS 0.008374f
C806 B.n662 VSUBS 0.008374f
C807 B.n663 VSUBS 0.008374f
C808 B.n664 VSUBS 0.008374f
C809 B.n665 VSUBS 0.008374f
C810 B.n666 VSUBS 0.008374f
C811 B.n667 VSUBS 0.008374f
C812 B.n668 VSUBS 0.008374f
C813 B.n669 VSUBS 0.008374f
C814 B.n670 VSUBS 0.008374f
C815 B.n671 VSUBS 0.008374f
C816 B.n672 VSUBS 0.008374f
C817 B.n673 VSUBS 0.008374f
C818 B.n674 VSUBS 0.008374f
C819 B.n675 VSUBS 0.008374f
C820 B.n676 VSUBS 0.008374f
C821 B.n677 VSUBS 0.008374f
C822 B.n678 VSUBS 0.008374f
C823 B.n679 VSUBS 0.008374f
C824 B.n680 VSUBS 0.008374f
C825 B.n681 VSUBS 0.008374f
C826 B.n682 VSUBS 0.008374f
C827 B.n683 VSUBS 0.008374f
C828 B.n684 VSUBS 0.008374f
C829 B.n685 VSUBS 0.008374f
C830 B.n686 VSUBS 0.008374f
C831 B.n687 VSUBS 0.008374f
C832 B.n688 VSUBS 0.008374f
C833 B.n689 VSUBS 0.008374f
C834 B.n690 VSUBS 0.008374f
C835 B.n691 VSUBS 0.010928f
C836 B.n692 VSUBS 0.011641f
C837 B.n693 VSUBS 0.023149f
.ends

