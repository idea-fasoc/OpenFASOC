* NGSPICE file created from diff_pair_sample_1030.ext - technology: sky130A

.subckt diff_pair_sample_1030 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X1 VTAIL.t8 VP.t0 VDD1.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X2 VDD2.t7 VN.t1 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=2.43375 ps=15.08 w=14.75 l=1.84
X3 VDD1.t8 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X4 VTAIL.t16 VN.t2 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X5 B.t22 B.t20 B.t21 B.t10 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=0 ps=0 w=14.75 l=1.84
X6 VDD2.t9 VN.t3 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X7 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=0 ps=0 w=14.75 l=1.84
X8 VTAIL.t3 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X9 VDD1.t6 VP.t3 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=2.43375 ps=15.08 w=14.75 l=1.84
X10 VTAIL.t14 VN.t4 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X11 VDD2.t1 VN.t5 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X12 VTAIL.t5 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X13 VTAIL.t12 VN.t6 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X14 VDD1.t4 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=5.7525 ps=30.28 w=14.75 l=1.84
X15 VDD1.t3 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=5.7525 ps=30.28 w=14.75 l=1.84
X16 VDD2.t4 VN.t7 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=5.7525 ps=30.28 w=14.75 l=1.84
X17 VDD2.t3 VN.t8 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=5.7525 ps=30.28 w=14.75 l=1.84
X18 VTAIL.t0 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X19 VDD1.t1 VP.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=2.43375 ps=15.08 w=14.75 l=1.84
X20 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=0 ps=0 w=14.75 l=1.84
X21 VDD2.t2 VN.t9 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=2.43375 ps=15.08 w=14.75 l=1.84
X22 VDD1.t0 VP.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.43375 pd=15.08 as=2.43375 ps=15.08 w=14.75 l=1.84
X23 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.7525 pd=30.28 as=0 ps=0 w=14.75 l=1.84
R0 VN.n7 VN.t1 228.012
R1 VN.n39 VN.t7 228.012
R2 VN.n8 VN.t6 193.194
R3 VN.n15 VN.t3 193.194
R4 VN.n22 VN.t0 193.194
R5 VN.n30 VN.t8 193.194
R6 VN.n40 VN.t4 193.194
R7 VN.n47 VN.t5 193.194
R8 VN.n54 VN.t2 193.194
R9 VN.n62 VN.t9 193.194
R10 VN.n31 VN.n30 181.363
R11 VN.n63 VN.n62 181.363
R12 VN.n61 VN.n32 161.3
R13 VN.n60 VN.n59 161.3
R14 VN.n58 VN.n33 161.3
R15 VN.n57 VN.n56 161.3
R16 VN.n55 VN.n34 161.3
R17 VN.n53 VN.n52 161.3
R18 VN.n51 VN.n35 161.3
R19 VN.n50 VN.n49 161.3
R20 VN.n48 VN.n36 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n37 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n41 VN.n38 161.3
R25 VN.n29 VN.n0 161.3
R26 VN.n28 VN.n27 161.3
R27 VN.n26 VN.n1 161.3
R28 VN.n25 VN.n24 161.3
R29 VN.n23 VN.n2 161.3
R30 VN.n21 VN.n20 161.3
R31 VN.n19 VN.n3 161.3
R32 VN.n18 VN.n17 161.3
R33 VN.n16 VN.n4 161.3
R34 VN.n14 VN.n13 161.3
R35 VN.n12 VN.n5 161.3
R36 VN.n11 VN.n10 161.3
R37 VN.n9 VN.n6 161.3
R38 VN.n10 VN.n5 56.5193
R39 VN.n17 VN.n3 56.5193
R40 VN.n42 VN.n37 56.5193
R41 VN.n49 VN.n35 56.5193
R42 VN VN.n63 51.3698
R43 VN.n8 VN.n7 48.825
R44 VN.n40 VN.n39 48.825
R45 VN.n28 VN.n1 40.979
R46 VN.n60 VN.n33 40.979
R47 VN.n24 VN.n1 40.0078
R48 VN.n56 VN.n33 40.0078
R49 VN.n10 VN.n9 24.4675
R50 VN.n14 VN.n5 24.4675
R51 VN.n17 VN.n16 24.4675
R52 VN.n21 VN.n3 24.4675
R53 VN.n24 VN.n23 24.4675
R54 VN.n29 VN.n28 24.4675
R55 VN.n42 VN.n41 24.4675
R56 VN.n49 VN.n48 24.4675
R57 VN.n46 VN.n37 24.4675
R58 VN.n56 VN.n55 24.4675
R59 VN.n53 VN.n35 24.4675
R60 VN.n61 VN.n60 24.4675
R61 VN.n9 VN.n8 20.5528
R62 VN.n22 VN.n21 20.5528
R63 VN.n41 VN.n40 20.5528
R64 VN.n54 VN.n53 20.5528
R65 VN.n39 VN.n38 12.2488
R66 VN.n7 VN.n6 12.2488
R67 VN.n15 VN.n14 12.234
R68 VN.n16 VN.n15 12.234
R69 VN.n48 VN.n47 12.234
R70 VN.n47 VN.n46 12.234
R71 VN.n30 VN.n29 4.40456
R72 VN.n62 VN.n61 4.40456
R73 VN.n23 VN.n22 3.91522
R74 VN.n55 VN.n54 3.91522
R75 VN.n63 VN.n32 0.189894
R76 VN.n59 VN.n32 0.189894
R77 VN.n59 VN.n58 0.189894
R78 VN.n58 VN.n57 0.189894
R79 VN.n57 VN.n34 0.189894
R80 VN.n52 VN.n34 0.189894
R81 VN.n52 VN.n51 0.189894
R82 VN.n51 VN.n50 0.189894
R83 VN.n50 VN.n36 0.189894
R84 VN.n45 VN.n36 0.189894
R85 VN.n45 VN.n44 0.189894
R86 VN.n44 VN.n43 0.189894
R87 VN.n43 VN.n38 0.189894
R88 VN.n11 VN.n6 0.189894
R89 VN.n12 VN.n11 0.189894
R90 VN.n13 VN.n12 0.189894
R91 VN.n13 VN.n4 0.189894
R92 VN.n18 VN.n4 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n20 VN.n19 0.189894
R95 VN.n20 VN.n2 0.189894
R96 VN.n25 VN.n2 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n27 VN.n26 0.189894
R99 VN.n27 VN.n0 0.189894
R100 VN.n31 VN.n0 0.189894
R101 VN VN.n31 0.0516364
R102 VDD2.n161 VDD2.n85 289.615
R103 VDD2.n76 VDD2.n0 289.615
R104 VDD2.n162 VDD2.n161 185
R105 VDD2.n160 VDD2.n159 185
R106 VDD2.n158 VDD2.n88 185
R107 VDD2.n92 VDD2.n89 185
R108 VDD2.n153 VDD2.n152 185
R109 VDD2.n151 VDD2.n150 185
R110 VDD2.n94 VDD2.n93 185
R111 VDD2.n145 VDD2.n144 185
R112 VDD2.n143 VDD2.n142 185
R113 VDD2.n98 VDD2.n97 185
R114 VDD2.n137 VDD2.n136 185
R115 VDD2.n135 VDD2.n134 185
R116 VDD2.n102 VDD2.n101 185
R117 VDD2.n129 VDD2.n128 185
R118 VDD2.n127 VDD2.n126 185
R119 VDD2.n106 VDD2.n105 185
R120 VDD2.n121 VDD2.n120 185
R121 VDD2.n119 VDD2.n118 185
R122 VDD2.n110 VDD2.n109 185
R123 VDD2.n113 VDD2.n112 185
R124 VDD2.n27 VDD2.n26 185
R125 VDD2.n24 VDD2.n23 185
R126 VDD2.n33 VDD2.n32 185
R127 VDD2.n35 VDD2.n34 185
R128 VDD2.n20 VDD2.n19 185
R129 VDD2.n41 VDD2.n40 185
R130 VDD2.n43 VDD2.n42 185
R131 VDD2.n16 VDD2.n15 185
R132 VDD2.n49 VDD2.n48 185
R133 VDD2.n51 VDD2.n50 185
R134 VDD2.n12 VDD2.n11 185
R135 VDD2.n57 VDD2.n56 185
R136 VDD2.n59 VDD2.n58 185
R137 VDD2.n8 VDD2.n7 185
R138 VDD2.n65 VDD2.n64 185
R139 VDD2.n68 VDD2.n67 185
R140 VDD2.n66 VDD2.n4 185
R141 VDD2.n73 VDD2.n3 185
R142 VDD2.n75 VDD2.n74 185
R143 VDD2.n77 VDD2.n76 185
R144 VDD2.t2 VDD2.n111 147.659
R145 VDD2.t7 VDD2.n25 147.659
R146 VDD2.n161 VDD2.n160 104.615
R147 VDD2.n160 VDD2.n88 104.615
R148 VDD2.n92 VDD2.n88 104.615
R149 VDD2.n152 VDD2.n92 104.615
R150 VDD2.n152 VDD2.n151 104.615
R151 VDD2.n151 VDD2.n93 104.615
R152 VDD2.n144 VDD2.n93 104.615
R153 VDD2.n144 VDD2.n143 104.615
R154 VDD2.n143 VDD2.n97 104.615
R155 VDD2.n136 VDD2.n97 104.615
R156 VDD2.n136 VDD2.n135 104.615
R157 VDD2.n135 VDD2.n101 104.615
R158 VDD2.n128 VDD2.n101 104.615
R159 VDD2.n128 VDD2.n127 104.615
R160 VDD2.n127 VDD2.n105 104.615
R161 VDD2.n120 VDD2.n105 104.615
R162 VDD2.n120 VDD2.n119 104.615
R163 VDD2.n119 VDD2.n109 104.615
R164 VDD2.n112 VDD2.n109 104.615
R165 VDD2.n26 VDD2.n23 104.615
R166 VDD2.n33 VDD2.n23 104.615
R167 VDD2.n34 VDD2.n33 104.615
R168 VDD2.n34 VDD2.n19 104.615
R169 VDD2.n41 VDD2.n19 104.615
R170 VDD2.n42 VDD2.n41 104.615
R171 VDD2.n42 VDD2.n15 104.615
R172 VDD2.n49 VDD2.n15 104.615
R173 VDD2.n50 VDD2.n49 104.615
R174 VDD2.n50 VDD2.n11 104.615
R175 VDD2.n57 VDD2.n11 104.615
R176 VDD2.n58 VDD2.n57 104.615
R177 VDD2.n58 VDD2.n7 104.615
R178 VDD2.n65 VDD2.n7 104.615
R179 VDD2.n67 VDD2.n65 104.615
R180 VDD2.n67 VDD2.n66 104.615
R181 VDD2.n66 VDD2.n3 104.615
R182 VDD2.n75 VDD2.n3 104.615
R183 VDD2.n76 VDD2.n75 104.615
R184 VDD2.n84 VDD2.n83 64.4019
R185 VDD2 VDD2.n169 64.3991
R186 VDD2.n168 VDD2.n167 63.0544
R187 VDD2.n82 VDD2.n81 63.0542
R188 VDD2.n82 VDD2.n80 52.8682
R189 VDD2.n112 VDD2.t2 52.3082
R190 VDD2.n26 VDD2.t7 52.3082
R191 VDD2.n166 VDD2.n165 50.9975
R192 VDD2.n166 VDD2.n84 45.3166
R193 VDD2.n113 VDD2.n111 15.6677
R194 VDD2.n27 VDD2.n25 15.6677
R195 VDD2.n159 VDD2.n158 13.1884
R196 VDD2.n74 VDD2.n73 13.1884
R197 VDD2.n162 VDD2.n87 12.8005
R198 VDD2.n157 VDD2.n89 12.8005
R199 VDD2.n114 VDD2.n110 12.8005
R200 VDD2.n28 VDD2.n24 12.8005
R201 VDD2.n72 VDD2.n4 12.8005
R202 VDD2.n77 VDD2.n2 12.8005
R203 VDD2.n163 VDD2.n85 12.0247
R204 VDD2.n154 VDD2.n153 12.0247
R205 VDD2.n118 VDD2.n117 12.0247
R206 VDD2.n32 VDD2.n31 12.0247
R207 VDD2.n69 VDD2.n68 12.0247
R208 VDD2.n78 VDD2.n0 12.0247
R209 VDD2.n150 VDD2.n91 11.249
R210 VDD2.n121 VDD2.n108 11.249
R211 VDD2.n35 VDD2.n22 11.249
R212 VDD2.n64 VDD2.n6 11.249
R213 VDD2.n149 VDD2.n94 10.4732
R214 VDD2.n122 VDD2.n106 10.4732
R215 VDD2.n36 VDD2.n20 10.4732
R216 VDD2.n63 VDD2.n8 10.4732
R217 VDD2.n146 VDD2.n145 9.69747
R218 VDD2.n126 VDD2.n125 9.69747
R219 VDD2.n40 VDD2.n39 9.69747
R220 VDD2.n60 VDD2.n59 9.69747
R221 VDD2.n165 VDD2.n164 9.45567
R222 VDD2.n80 VDD2.n79 9.45567
R223 VDD2.n139 VDD2.n138 9.3005
R224 VDD2.n141 VDD2.n140 9.3005
R225 VDD2.n96 VDD2.n95 9.3005
R226 VDD2.n147 VDD2.n146 9.3005
R227 VDD2.n149 VDD2.n148 9.3005
R228 VDD2.n91 VDD2.n90 9.3005
R229 VDD2.n155 VDD2.n154 9.3005
R230 VDD2.n157 VDD2.n156 9.3005
R231 VDD2.n164 VDD2.n163 9.3005
R232 VDD2.n87 VDD2.n86 9.3005
R233 VDD2.n100 VDD2.n99 9.3005
R234 VDD2.n133 VDD2.n132 9.3005
R235 VDD2.n131 VDD2.n130 9.3005
R236 VDD2.n104 VDD2.n103 9.3005
R237 VDD2.n125 VDD2.n124 9.3005
R238 VDD2.n123 VDD2.n122 9.3005
R239 VDD2.n108 VDD2.n107 9.3005
R240 VDD2.n117 VDD2.n116 9.3005
R241 VDD2.n115 VDD2.n114 9.3005
R242 VDD2.n79 VDD2.n78 9.3005
R243 VDD2.n2 VDD2.n1 9.3005
R244 VDD2.n47 VDD2.n46 9.3005
R245 VDD2.n45 VDD2.n44 9.3005
R246 VDD2.n18 VDD2.n17 9.3005
R247 VDD2.n39 VDD2.n38 9.3005
R248 VDD2.n37 VDD2.n36 9.3005
R249 VDD2.n22 VDD2.n21 9.3005
R250 VDD2.n31 VDD2.n30 9.3005
R251 VDD2.n29 VDD2.n28 9.3005
R252 VDD2.n14 VDD2.n13 9.3005
R253 VDD2.n53 VDD2.n52 9.3005
R254 VDD2.n55 VDD2.n54 9.3005
R255 VDD2.n10 VDD2.n9 9.3005
R256 VDD2.n61 VDD2.n60 9.3005
R257 VDD2.n63 VDD2.n62 9.3005
R258 VDD2.n6 VDD2.n5 9.3005
R259 VDD2.n70 VDD2.n69 9.3005
R260 VDD2.n72 VDD2.n71 9.3005
R261 VDD2.n142 VDD2.n96 8.92171
R262 VDD2.n129 VDD2.n104 8.92171
R263 VDD2.n43 VDD2.n18 8.92171
R264 VDD2.n56 VDD2.n10 8.92171
R265 VDD2.n141 VDD2.n98 8.14595
R266 VDD2.n130 VDD2.n102 8.14595
R267 VDD2.n44 VDD2.n16 8.14595
R268 VDD2.n55 VDD2.n12 8.14595
R269 VDD2.n138 VDD2.n137 7.3702
R270 VDD2.n134 VDD2.n133 7.3702
R271 VDD2.n48 VDD2.n47 7.3702
R272 VDD2.n52 VDD2.n51 7.3702
R273 VDD2.n137 VDD2.n100 6.59444
R274 VDD2.n134 VDD2.n100 6.59444
R275 VDD2.n48 VDD2.n14 6.59444
R276 VDD2.n51 VDD2.n14 6.59444
R277 VDD2.n138 VDD2.n98 5.81868
R278 VDD2.n133 VDD2.n102 5.81868
R279 VDD2.n47 VDD2.n16 5.81868
R280 VDD2.n52 VDD2.n12 5.81868
R281 VDD2.n142 VDD2.n141 5.04292
R282 VDD2.n130 VDD2.n129 5.04292
R283 VDD2.n44 VDD2.n43 5.04292
R284 VDD2.n56 VDD2.n55 5.04292
R285 VDD2.n115 VDD2.n111 4.38563
R286 VDD2.n29 VDD2.n25 4.38563
R287 VDD2.n145 VDD2.n96 4.26717
R288 VDD2.n126 VDD2.n104 4.26717
R289 VDD2.n40 VDD2.n18 4.26717
R290 VDD2.n59 VDD2.n10 4.26717
R291 VDD2.n146 VDD2.n94 3.49141
R292 VDD2.n125 VDD2.n106 3.49141
R293 VDD2.n39 VDD2.n20 3.49141
R294 VDD2.n60 VDD2.n8 3.49141
R295 VDD2.n150 VDD2.n149 2.71565
R296 VDD2.n122 VDD2.n121 2.71565
R297 VDD2.n36 VDD2.n35 2.71565
R298 VDD2.n64 VDD2.n63 2.71565
R299 VDD2.n165 VDD2.n85 1.93989
R300 VDD2.n153 VDD2.n91 1.93989
R301 VDD2.n118 VDD2.n108 1.93989
R302 VDD2.n32 VDD2.n22 1.93989
R303 VDD2.n68 VDD2.n6 1.93989
R304 VDD2.n80 VDD2.n0 1.93989
R305 VDD2.n168 VDD2.n166 1.87119
R306 VDD2.n169 VDD2.t8 1.34287
R307 VDD2.n169 VDD2.t4 1.34287
R308 VDD2.n167 VDD2.t6 1.34287
R309 VDD2.n167 VDD2.t1 1.34287
R310 VDD2.n83 VDD2.t5 1.34287
R311 VDD2.n83 VDD2.t3 1.34287
R312 VDD2.n81 VDD2.t0 1.34287
R313 VDD2.n81 VDD2.t9 1.34287
R314 VDD2.n163 VDD2.n162 1.16414
R315 VDD2.n154 VDD2.n89 1.16414
R316 VDD2.n117 VDD2.n110 1.16414
R317 VDD2.n31 VDD2.n24 1.16414
R318 VDD2.n69 VDD2.n4 1.16414
R319 VDD2.n78 VDD2.n77 1.16414
R320 VDD2 VDD2.n168 0.526362
R321 VDD2.n84 VDD2.n82 0.412826
R322 VDD2.n159 VDD2.n87 0.388379
R323 VDD2.n158 VDD2.n157 0.388379
R324 VDD2.n114 VDD2.n113 0.388379
R325 VDD2.n28 VDD2.n27 0.388379
R326 VDD2.n73 VDD2.n72 0.388379
R327 VDD2.n74 VDD2.n2 0.388379
R328 VDD2.n164 VDD2.n86 0.155672
R329 VDD2.n156 VDD2.n86 0.155672
R330 VDD2.n156 VDD2.n155 0.155672
R331 VDD2.n155 VDD2.n90 0.155672
R332 VDD2.n148 VDD2.n90 0.155672
R333 VDD2.n148 VDD2.n147 0.155672
R334 VDD2.n147 VDD2.n95 0.155672
R335 VDD2.n140 VDD2.n95 0.155672
R336 VDD2.n140 VDD2.n139 0.155672
R337 VDD2.n139 VDD2.n99 0.155672
R338 VDD2.n132 VDD2.n99 0.155672
R339 VDD2.n132 VDD2.n131 0.155672
R340 VDD2.n131 VDD2.n103 0.155672
R341 VDD2.n124 VDD2.n103 0.155672
R342 VDD2.n124 VDD2.n123 0.155672
R343 VDD2.n123 VDD2.n107 0.155672
R344 VDD2.n116 VDD2.n107 0.155672
R345 VDD2.n116 VDD2.n115 0.155672
R346 VDD2.n30 VDD2.n29 0.155672
R347 VDD2.n30 VDD2.n21 0.155672
R348 VDD2.n37 VDD2.n21 0.155672
R349 VDD2.n38 VDD2.n37 0.155672
R350 VDD2.n38 VDD2.n17 0.155672
R351 VDD2.n45 VDD2.n17 0.155672
R352 VDD2.n46 VDD2.n45 0.155672
R353 VDD2.n46 VDD2.n13 0.155672
R354 VDD2.n53 VDD2.n13 0.155672
R355 VDD2.n54 VDD2.n53 0.155672
R356 VDD2.n54 VDD2.n9 0.155672
R357 VDD2.n61 VDD2.n9 0.155672
R358 VDD2.n62 VDD2.n61 0.155672
R359 VDD2.n62 VDD2.n5 0.155672
R360 VDD2.n70 VDD2.n5 0.155672
R361 VDD2.n71 VDD2.n70 0.155672
R362 VDD2.n71 VDD2.n1 0.155672
R363 VDD2.n79 VDD2.n1 0.155672
R364 VTAIL.n336 VTAIL.n260 289.615
R365 VTAIL.n78 VTAIL.n2 289.615
R366 VTAIL.n254 VTAIL.n178 289.615
R367 VTAIL.n168 VTAIL.n92 289.615
R368 VTAIL.n287 VTAIL.n286 185
R369 VTAIL.n284 VTAIL.n283 185
R370 VTAIL.n293 VTAIL.n292 185
R371 VTAIL.n295 VTAIL.n294 185
R372 VTAIL.n280 VTAIL.n279 185
R373 VTAIL.n301 VTAIL.n300 185
R374 VTAIL.n303 VTAIL.n302 185
R375 VTAIL.n276 VTAIL.n275 185
R376 VTAIL.n309 VTAIL.n308 185
R377 VTAIL.n311 VTAIL.n310 185
R378 VTAIL.n272 VTAIL.n271 185
R379 VTAIL.n317 VTAIL.n316 185
R380 VTAIL.n319 VTAIL.n318 185
R381 VTAIL.n268 VTAIL.n267 185
R382 VTAIL.n325 VTAIL.n324 185
R383 VTAIL.n328 VTAIL.n327 185
R384 VTAIL.n326 VTAIL.n264 185
R385 VTAIL.n333 VTAIL.n263 185
R386 VTAIL.n335 VTAIL.n334 185
R387 VTAIL.n337 VTAIL.n336 185
R388 VTAIL.n29 VTAIL.n28 185
R389 VTAIL.n26 VTAIL.n25 185
R390 VTAIL.n35 VTAIL.n34 185
R391 VTAIL.n37 VTAIL.n36 185
R392 VTAIL.n22 VTAIL.n21 185
R393 VTAIL.n43 VTAIL.n42 185
R394 VTAIL.n45 VTAIL.n44 185
R395 VTAIL.n18 VTAIL.n17 185
R396 VTAIL.n51 VTAIL.n50 185
R397 VTAIL.n53 VTAIL.n52 185
R398 VTAIL.n14 VTAIL.n13 185
R399 VTAIL.n59 VTAIL.n58 185
R400 VTAIL.n61 VTAIL.n60 185
R401 VTAIL.n10 VTAIL.n9 185
R402 VTAIL.n67 VTAIL.n66 185
R403 VTAIL.n70 VTAIL.n69 185
R404 VTAIL.n68 VTAIL.n6 185
R405 VTAIL.n75 VTAIL.n5 185
R406 VTAIL.n77 VTAIL.n76 185
R407 VTAIL.n79 VTAIL.n78 185
R408 VTAIL.n255 VTAIL.n254 185
R409 VTAIL.n253 VTAIL.n252 185
R410 VTAIL.n251 VTAIL.n181 185
R411 VTAIL.n185 VTAIL.n182 185
R412 VTAIL.n246 VTAIL.n245 185
R413 VTAIL.n244 VTAIL.n243 185
R414 VTAIL.n187 VTAIL.n186 185
R415 VTAIL.n238 VTAIL.n237 185
R416 VTAIL.n236 VTAIL.n235 185
R417 VTAIL.n191 VTAIL.n190 185
R418 VTAIL.n230 VTAIL.n229 185
R419 VTAIL.n228 VTAIL.n227 185
R420 VTAIL.n195 VTAIL.n194 185
R421 VTAIL.n222 VTAIL.n221 185
R422 VTAIL.n220 VTAIL.n219 185
R423 VTAIL.n199 VTAIL.n198 185
R424 VTAIL.n214 VTAIL.n213 185
R425 VTAIL.n212 VTAIL.n211 185
R426 VTAIL.n203 VTAIL.n202 185
R427 VTAIL.n206 VTAIL.n205 185
R428 VTAIL.n169 VTAIL.n168 185
R429 VTAIL.n167 VTAIL.n166 185
R430 VTAIL.n165 VTAIL.n95 185
R431 VTAIL.n99 VTAIL.n96 185
R432 VTAIL.n160 VTAIL.n159 185
R433 VTAIL.n158 VTAIL.n157 185
R434 VTAIL.n101 VTAIL.n100 185
R435 VTAIL.n152 VTAIL.n151 185
R436 VTAIL.n150 VTAIL.n149 185
R437 VTAIL.n105 VTAIL.n104 185
R438 VTAIL.n144 VTAIL.n143 185
R439 VTAIL.n142 VTAIL.n141 185
R440 VTAIL.n109 VTAIL.n108 185
R441 VTAIL.n136 VTAIL.n135 185
R442 VTAIL.n134 VTAIL.n133 185
R443 VTAIL.n113 VTAIL.n112 185
R444 VTAIL.n128 VTAIL.n127 185
R445 VTAIL.n126 VTAIL.n125 185
R446 VTAIL.n117 VTAIL.n116 185
R447 VTAIL.n120 VTAIL.n119 185
R448 VTAIL.t6 VTAIL.n204 147.659
R449 VTAIL.t11 VTAIL.n118 147.659
R450 VTAIL.t10 VTAIL.n285 147.659
R451 VTAIL.t1 VTAIL.n27 147.659
R452 VTAIL.n286 VTAIL.n283 104.615
R453 VTAIL.n293 VTAIL.n283 104.615
R454 VTAIL.n294 VTAIL.n293 104.615
R455 VTAIL.n294 VTAIL.n279 104.615
R456 VTAIL.n301 VTAIL.n279 104.615
R457 VTAIL.n302 VTAIL.n301 104.615
R458 VTAIL.n302 VTAIL.n275 104.615
R459 VTAIL.n309 VTAIL.n275 104.615
R460 VTAIL.n310 VTAIL.n309 104.615
R461 VTAIL.n310 VTAIL.n271 104.615
R462 VTAIL.n317 VTAIL.n271 104.615
R463 VTAIL.n318 VTAIL.n317 104.615
R464 VTAIL.n318 VTAIL.n267 104.615
R465 VTAIL.n325 VTAIL.n267 104.615
R466 VTAIL.n327 VTAIL.n325 104.615
R467 VTAIL.n327 VTAIL.n326 104.615
R468 VTAIL.n326 VTAIL.n263 104.615
R469 VTAIL.n335 VTAIL.n263 104.615
R470 VTAIL.n336 VTAIL.n335 104.615
R471 VTAIL.n28 VTAIL.n25 104.615
R472 VTAIL.n35 VTAIL.n25 104.615
R473 VTAIL.n36 VTAIL.n35 104.615
R474 VTAIL.n36 VTAIL.n21 104.615
R475 VTAIL.n43 VTAIL.n21 104.615
R476 VTAIL.n44 VTAIL.n43 104.615
R477 VTAIL.n44 VTAIL.n17 104.615
R478 VTAIL.n51 VTAIL.n17 104.615
R479 VTAIL.n52 VTAIL.n51 104.615
R480 VTAIL.n52 VTAIL.n13 104.615
R481 VTAIL.n59 VTAIL.n13 104.615
R482 VTAIL.n60 VTAIL.n59 104.615
R483 VTAIL.n60 VTAIL.n9 104.615
R484 VTAIL.n67 VTAIL.n9 104.615
R485 VTAIL.n69 VTAIL.n67 104.615
R486 VTAIL.n69 VTAIL.n68 104.615
R487 VTAIL.n68 VTAIL.n5 104.615
R488 VTAIL.n77 VTAIL.n5 104.615
R489 VTAIL.n78 VTAIL.n77 104.615
R490 VTAIL.n254 VTAIL.n253 104.615
R491 VTAIL.n253 VTAIL.n181 104.615
R492 VTAIL.n185 VTAIL.n181 104.615
R493 VTAIL.n245 VTAIL.n185 104.615
R494 VTAIL.n245 VTAIL.n244 104.615
R495 VTAIL.n244 VTAIL.n186 104.615
R496 VTAIL.n237 VTAIL.n186 104.615
R497 VTAIL.n237 VTAIL.n236 104.615
R498 VTAIL.n236 VTAIL.n190 104.615
R499 VTAIL.n229 VTAIL.n190 104.615
R500 VTAIL.n229 VTAIL.n228 104.615
R501 VTAIL.n228 VTAIL.n194 104.615
R502 VTAIL.n221 VTAIL.n194 104.615
R503 VTAIL.n221 VTAIL.n220 104.615
R504 VTAIL.n220 VTAIL.n198 104.615
R505 VTAIL.n213 VTAIL.n198 104.615
R506 VTAIL.n213 VTAIL.n212 104.615
R507 VTAIL.n212 VTAIL.n202 104.615
R508 VTAIL.n205 VTAIL.n202 104.615
R509 VTAIL.n168 VTAIL.n167 104.615
R510 VTAIL.n167 VTAIL.n95 104.615
R511 VTAIL.n99 VTAIL.n95 104.615
R512 VTAIL.n159 VTAIL.n99 104.615
R513 VTAIL.n159 VTAIL.n158 104.615
R514 VTAIL.n158 VTAIL.n100 104.615
R515 VTAIL.n151 VTAIL.n100 104.615
R516 VTAIL.n151 VTAIL.n150 104.615
R517 VTAIL.n150 VTAIL.n104 104.615
R518 VTAIL.n143 VTAIL.n104 104.615
R519 VTAIL.n143 VTAIL.n142 104.615
R520 VTAIL.n142 VTAIL.n108 104.615
R521 VTAIL.n135 VTAIL.n108 104.615
R522 VTAIL.n135 VTAIL.n134 104.615
R523 VTAIL.n134 VTAIL.n112 104.615
R524 VTAIL.n127 VTAIL.n112 104.615
R525 VTAIL.n127 VTAIL.n126 104.615
R526 VTAIL.n126 VTAIL.n116 104.615
R527 VTAIL.n119 VTAIL.n116 104.615
R528 VTAIL.n286 VTAIL.t10 52.3082
R529 VTAIL.n28 VTAIL.t1 52.3082
R530 VTAIL.n205 VTAIL.t6 52.3082
R531 VTAIL.n119 VTAIL.t11 52.3082
R532 VTAIL.n177 VTAIL.n176 46.3756
R533 VTAIL.n175 VTAIL.n174 46.3756
R534 VTAIL.n91 VTAIL.n90 46.3756
R535 VTAIL.n89 VTAIL.n88 46.3756
R536 VTAIL.n343 VTAIL.n342 46.3755
R537 VTAIL.n1 VTAIL.n0 46.3755
R538 VTAIL.n85 VTAIL.n84 46.3755
R539 VTAIL.n87 VTAIL.n86 46.3755
R540 VTAIL.n341 VTAIL.n340 34.3187
R541 VTAIL.n83 VTAIL.n82 34.3187
R542 VTAIL.n259 VTAIL.n258 34.3187
R543 VTAIL.n173 VTAIL.n172 34.3187
R544 VTAIL.n89 VTAIL.n87 28.8238
R545 VTAIL.n341 VTAIL.n259 26.9531
R546 VTAIL.n287 VTAIL.n285 15.6677
R547 VTAIL.n29 VTAIL.n27 15.6677
R548 VTAIL.n206 VTAIL.n204 15.6677
R549 VTAIL.n120 VTAIL.n118 15.6677
R550 VTAIL.n334 VTAIL.n333 13.1884
R551 VTAIL.n76 VTAIL.n75 13.1884
R552 VTAIL.n252 VTAIL.n251 13.1884
R553 VTAIL.n166 VTAIL.n165 13.1884
R554 VTAIL.n288 VTAIL.n284 12.8005
R555 VTAIL.n332 VTAIL.n264 12.8005
R556 VTAIL.n337 VTAIL.n262 12.8005
R557 VTAIL.n30 VTAIL.n26 12.8005
R558 VTAIL.n74 VTAIL.n6 12.8005
R559 VTAIL.n79 VTAIL.n4 12.8005
R560 VTAIL.n255 VTAIL.n180 12.8005
R561 VTAIL.n250 VTAIL.n182 12.8005
R562 VTAIL.n207 VTAIL.n203 12.8005
R563 VTAIL.n169 VTAIL.n94 12.8005
R564 VTAIL.n164 VTAIL.n96 12.8005
R565 VTAIL.n121 VTAIL.n117 12.8005
R566 VTAIL.n292 VTAIL.n291 12.0247
R567 VTAIL.n329 VTAIL.n328 12.0247
R568 VTAIL.n338 VTAIL.n260 12.0247
R569 VTAIL.n34 VTAIL.n33 12.0247
R570 VTAIL.n71 VTAIL.n70 12.0247
R571 VTAIL.n80 VTAIL.n2 12.0247
R572 VTAIL.n256 VTAIL.n178 12.0247
R573 VTAIL.n247 VTAIL.n246 12.0247
R574 VTAIL.n211 VTAIL.n210 12.0247
R575 VTAIL.n170 VTAIL.n92 12.0247
R576 VTAIL.n161 VTAIL.n160 12.0247
R577 VTAIL.n125 VTAIL.n124 12.0247
R578 VTAIL.n295 VTAIL.n282 11.249
R579 VTAIL.n324 VTAIL.n266 11.249
R580 VTAIL.n37 VTAIL.n24 11.249
R581 VTAIL.n66 VTAIL.n8 11.249
R582 VTAIL.n243 VTAIL.n184 11.249
R583 VTAIL.n214 VTAIL.n201 11.249
R584 VTAIL.n157 VTAIL.n98 11.249
R585 VTAIL.n128 VTAIL.n115 11.249
R586 VTAIL.n296 VTAIL.n280 10.4732
R587 VTAIL.n323 VTAIL.n268 10.4732
R588 VTAIL.n38 VTAIL.n22 10.4732
R589 VTAIL.n65 VTAIL.n10 10.4732
R590 VTAIL.n242 VTAIL.n187 10.4732
R591 VTAIL.n215 VTAIL.n199 10.4732
R592 VTAIL.n156 VTAIL.n101 10.4732
R593 VTAIL.n129 VTAIL.n113 10.4732
R594 VTAIL.n300 VTAIL.n299 9.69747
R595 VTAIL.n320 VTAIL.n319 9.69747
R596 VTAIL.n42 VTAIL.n41 9.69747
R597 VTAIL.n62 VTAIL.n61 9.69747
R598 VTAIL.n239 VTAIL.n238 9.69747
R599 VTAIL.n219 VTAIL.n218 9.69747
R600 VTAIL.n153 VTAIL.n152 9.69747
R601 VTAIL.n133 VTAIL.n132 9.69747
R602 VTAIL.n340 VTAIL.n339 9.45567
R603 VTAIL.n82 VTAIL.n81 9.45567
R604 VTAIL.n258 VTAIL.n257 9.45567
R605 VTAIL.n172 VTAIL.n171 9.45567
R606 VTAIL.n339 VTAIL.n338 9.3005
R607 VTAIL.n262 VTAIL.n261 9.3005
R608 VTAIL.n307 VTAIL.n306 9.3005
R609 VTAIL.n305 VTAIL.n304 9.3005
R610 VTAIL.n278 VTAIL.n277 9.3005
R611 VTAIL.n299 VTAIL.n298 9.3005
R612 VTAIL.n297 VTAIL.n296 9.3005
R613 VTAIL.n282 VTAIL.n281 9.3005
R614 VTAIL.n291 VTAIL.n290 9.3005
R615 VTAIL.n289 VTAIL.n288 9.3005
R616 VTAIL.n274 VTAIL.n273 9.3005
R617 VTAIL.n313 VTAIL.n312 9.3005
R618 VTAIL.n315 VTAIL.n314 9.3005
R619 VTAIL.n270 VTAIL.n269 9.3005
R620 VTAIL.n321 VTAIL.n320 9.3005
R621 VTAIL.n323 VTAIL.n322 9.3005
R622 VTAIL.n266 VTAIL.n265 9.3005
R623 VTAIL.n330 VTAIL.n329 9.3005
R624 VTAIL.n332 VTAIL.n331 9.3005
R625 VTAIL.n81 VTAIL.n80 9.3005
R626 VTAIL.n4 VTAIL.n3 9.3005
R627 VTAIL.n49 VTAIL.n48 9.3005
R628 VTAIL.n47 VTAIL.n46 9.3005
R629 VTAIL.n20 VTAIL.n19 9.3005
R630 VTAIL.n41 VTAIL.n40 9.3005
R631 VTAIL.n39 VTAIL.n38 9.3005
R632 VTAIL.n24 VTAIL.n23 9.3005
R633 VTAIL.n33 VTAIL.n32 9.3005
R634 VTAIL.n31 VTAIL.n30 9.3005
R635 VTAIL.n16 VTAIL.n15 9.3005
R636 VTAIL.n55 VTAIL.n54 9.3005
R637 VTAIL.n57 VTAIL.n56 9.3005
R638 VTAIL.n12 VTAIL.n11 9.3005
R639 VTAIL.n63 VTAIL.n62 9.3005
R640 VTAIL.n65 VTAIL.n64 9.3005
R641 VTAIL.n8 VTAIL.n7 9.3005
R642 VTAIL.n72 VTAIL.n71 9.3005
R643 VTAIL.n74 VTAIL.n73 9.3005
R644 VTAIL.n232 VTAIL.n231 9.3005
R645 VTAIL.n234 VTAIL.n233 9.3005
R646 VTAIL.n189 VTAIL.n188 9.3005
R647 VTAIL.n240 VTAIL.n239 9.3005
R648 VTAIL.n242 VTAIL.n241 9.3005
R649 VTAIL.n184 VTAIL.n183 9.3005
R650 VTAIL.n248 VTAIL.n247 9.3005
R651 VTAIL.n250 VTAIL.n249 9.3005
R652 VTAIL.n257 VTAIL.n256 9.3005
R653 VTAIL.n180 VTAIL.n179 9.3005
R654 VTAIL.n193 VTAIL.n192 9.3005
R655 VTAIL.n226 VTAIL.n225 9.3005
R656 VTAIL.n224 VTAIL.n223 9.3005
R657 VTAIL.n197 VTAIL.n196 9.3005
R658 VTAIL.n218 VTAIL.n217 9.3005
R659 VTAIL.n216 VTAIL.n215 9.3005
R660 VTAIL.n201 VTAIL.n200 9.3005
R661 VTAIL.n210 VTAIL.n209 9.3005
R662 VTAIL.n208 VTAIL.n207 9.3005
R663 VTAIL.n146 VTAIL.n145 9.3005
R664 VTAIL.n148 VTAIL.n147 9.3005
R665 VTAIL.n103 VTAIL.n102 9.3005
R666 VTAIL.n154 VTAIL.n153 9.3005
R667 VTAIL.n156 VTAIL.n155 9.3005
R668 VTAIL.n98 VTAIL.n97 9.3005
R669 VTAIL.n162 VTAIL.n161 9.3005
R670 VTAIL.n164 VTAIL.n163 9.3005
R671 VTAIL.n171 VTAIL.n170 9.3005
R672 VTAIL.n94 VTAIL.n93 9.3005
R673 VTAIL.n107 VTAIL.n106 9.3005
R674 VTAIL.n140 VTAIL.n139 9.3005
R675 VTAIL.n138 VTAIL.n137 9.3005
R676 VTAIL.n111 VTAIL.n110 9.3005
R677 VTAIL.n132 VTAIL.n131 9.3005
R678 VTAIL.n130 VTAIL.n129 9.3005
R679 VTAIL.n115 VTAIL.n114 9.3005
R680 VTAIL.n124 VTAIL.n123 9.3005
R681 VTAIL.n122 VTAIL.n121 9.3005
R682 VTAIL.n303 VTAIL.n278 8.92171
R683 VTAIL.n316 VTAIL.n270 8.92171
R684 VTAIL.n45 VTAIL.n20 8.92171
R685 VTAIL.n58 VTAIL.n12 8.92171
R686 VTAIL.n235 VTAIL.n189 8.92171
R687 VTAIL.n222 VTAIL.n197 8.92171
R688 VTAIL.n149 VTAIL.n103 8.92171
R689 VTAIL.n136 VTAIL.n111 8.92171
R690 VTAIL.n304 VTAIL.n276 8.14595
R691 VTAIL.n315 VTAIL.n272 8.14595
R692 VTAIL.n46 VTAIL.n18 8.14595
R693 VTAIL.n57 VTAIL.n14 8.14595
R694 VTAIL.n234 VTAIL.n191 8.14595
R695 VTAIL.n223 VTAIL.n195 8.14595
R696 VTAIL.n148 VTAIL.n105 8.14595
R697 VTAIL.n137 VTAIL.n109 8.14595
R698 VTAIL.n308 VTAIL.n307 7.3702
R699 VTAIL.n312 VTAIL.n311 7.3702
R700 VTAIL.n50 VTAIL.n49 7.3702
R701 VTAIL.n54 VTAIL.n53 7.3702
R702 VTAIL.n231 VTAIL.n230 7.3702
R703 VTAIL.n227 VTAIL.n226 7.3702
R704 VTAIL.n145 VTAIL.n144 7.3702
R705 VTAIL.n141 VTAIL.n140 7.3702
R706 VTAIL.n308 VTAIL.n274 6.59444
R707 VTAIL.n311 VTAIL.n274 6.59444
R708 VTAIL.n50 VTAIL.n16 6.59444
R709 VTAIL.n53 VTAIL.n16 6.59444
R710 VTAIL.n230 VTAIL.n193 6.59444
R711 VTAIL.n227 VTAIL.n193 6.59444
R712 VTAIL.n144 VTAIL.n107 6.59444
R713 VTAIL.n141 VTAIL.n107 6.59444
R714 VTAIL.n307 VTAIL.n276 5.81868
R715 VTAIL.n312 VTAIL.n272 5.81868
R716 VTAIL.n49 VTAIL.n18 5.81868
R717 VTAIL.n54 VTAIL.n14 5.81868
R718 VTAIL.n231 VTAIL.n191 5.81868
R719 VTAIL.n226 VTAIL.n195 5.81868
R720 VTAIL.n145 VTAIL.n105 5.81868
R721 VTAIL.n140 VTAIL.n109 5.81868
R722 VTAIL.n304 VTAIL.n303 5.04292
R723 VTAIL.n316 VTAIL.n315 5.04292
R724 VTAIL.n46 VTAIL.n45 5.04292
R725 VTAIL.n58 VTAIL.n57 5.04292
R726 VTAIL.n235 VTAIL.n234 5.04292
R727 VTAIL.n223 VTAIL.n222 5.04292
R728 VTAIL.n149 VTAIL.n148 5.04292
R729 VTAIL.n137 VTAIL.n136 5.04292
R730 VTAIL.n208 VTAIL.n204 4.38563
R731 VTAIL.n122 VTAIL.n118 4.38563
R732 VTAIL.n289 VTAIL.n285 4.38563
R733 VTAIL.n31 VTAIL.n27 4.38563
R734 VTAIL.n300 VTAIL.n278 4.26717
R735 VTAIL.n319 VTAIL.n270 4.26717
R736 VTAIL.n42 VTAIL.n20 4.26717
R737 VTAIL.n61 VTAIL.n12 4.26717
R738 VTAIL.n238 VTAIL.n189 4.26717
R739 VTAIL.n219 VTAIL.n197 4.26717
R740 VTAIL.n152 VTAIL.n103 4.26717
R741 VTAIL.n133 VTAIL.n111 4.26717
R742 VTAIL.n299 VTAIL.n280 3.49141
R743 VTAIL.n320 VTAIL.n268 3.49141
R744 VTAIL.n41 VTAIL.n22 3.49141
R745 VTAIL.n62 VTAIL.n10 3.49141
R746 VTAIL.n239 VTAIL.n187 3.49141
R747 VTAIL.n218 VTAIL.n199 3.49141
R748 VTAIL.n153 VTAIL.n101 3.49141
R749 VTAIL.n132 VTAIL.n113 3.49141
R750 VTAIL.n296 VTAIL.n295 2.71565
R751 VTAIL.n324 VTAIL.n323 2.71565
R752 VTAIL.n38 VTAIL.n37 2.71565
R753 VTAIL.n66 VTAIL.n65 2.71565
R754 VTAIL.n243 VTAIL.n242 2.71565
R755 VTAIL.n215 VTAIL.n214 2.71565
R756 VTAIL.n157 VTAIL.n156 2.71565
R757 VTAIL.n129 VTAIL.n128 2.71565
R758 VTAIL.n292 VTAIL.n282 1.93989
R759 VTAIL.n328 VTAIL.n266 1.93989
R760 VTAIL.n340 VTAIL.n260 1.93989
R761 VTAIL.n34 VTAIL.n24 1.93989
R762 VTAIL.n70 VTAIL.n8 1.93989
R763 VTAIL.n82 VTAIL.n2 1.93989
R764 VTAIL.n258 VTAIL.n178 1.93989
R765 VTAIL.n246 VTAIL.n184 1.93989
R766 VTAIL.n211 VTAIL.n201 1.93989
R767 VTAIL.n172 VTAIL.n92 1.93989
R768 VTAIL.n160 VTAIL.n98 1.93989
R769 VTAIL.n125 VTAIL.n115 1.93989
R770 VTAIL.n91 VTAIL.n89 1.87119
R771 VTAIL.n173 VTAIL.n91 1.87119
R772 VTAIL.n177 VTAIL.n175 1.87119
R773 VTAIL.n259 VTAIL.n177 1.87119
R774 VTAIL.n87 VTAIL.n85 1.87119
R775 VTAIL.n85 VTAIL.n83 1.87119
R776 VTAIL.n343 VTAIL.n341 1.87119
R777 VTAIL VTAIL.n1 1.46171
R778 VTAIL.n175 VTAIL.n173 1.40567
R779 VTAIL.n83 VTAIL.n1 1.40567
R780 VTAIL.n342 VTAIL.t15 1.34287
R781 VTAIL.n342 VTAIL.t18 1.34287
R782 VTAIL.n0 VTAIL.t17 1.34287
R783 VTAIL.n0 VTAIL.t12 1.34287
R784 VTAIL.n84 VTAIL.t7 1.34287
R785 VTAIL.n84 VTAIL.t3 1.34287
R786 VTAIL.n86 VTAIL.t19 1.34287
R787 VTAIL.n86 VTAIL.t0 1.34287
R788 VTAIL.n176 VTAIL.t4 1.34287
R789 VTAIL.n176 VTAIL.t8 1.34287
R790 VTAIL.n174 VTAIL.t2 1.34287
R791 VTAIL.n174 VTAIL.t5 1.34287
R792 VTAIL.n90 VTAIL.t13 1.34287
R793 VTAIL.n90 VTAIL.t14 1.34287
R794 VTAIL.n88 VTAIL.t9 1.34287
R795 VTAIL.n88 VTAIL.t16 1.34287
R796 VTAIL.n291 VTAIL.n284 1.16414
R797 VTAIL.n329 VTAIL.n264 1.16414
R798 VTAIL.n338 VTAIL.n337 1.16414
R799 VTAIL.n33 VTAIL.n26 1.16414
R800 VTAIL.n71 VTAIL.n6 1.16414
R801 VTAIL.n80 VTAIL.n79 1.16414
R802 VTAIL.n256 VTAIL.n255 1.16414
R803 VTAIL.n247 VTAIL.n182 1.16414
R804 VTAIL.n210 VTAIL.n203 1.16414
R805 VTAIL.n170 VTAIL.n169 1.16414
R806 VTAIL.n161 VTAIL.n96 1.16414
R807 VTAIL.n124 VTAIL.n117 1.16414
R808 VTAIL VTAIL.n343 0.409983
R809 VTAIL.n288 VTAIL.n287 0.388379
R810 VTAIL.n333 VTAIL.n332 0.388379
R811 VTAIL.n334 VTAIL.n262 0.388379
R812 VTAIL.n30 VTAIL.n29 0.388379
R813 VTAIL.n75 VTAIL.n74 0.388379
R814 VTAIL.n76 VTAIL.n4 0.388379
R815 VTAIL.n252 VTAIL.n180 0.388379
R816 VTAIL.n251 VTAIL.n250 0.388379
R817 VTAIL.n207 VTAIL.n206 0.388379
R818 VTAIL.n166 VTAIL.n94 0.388379
R819 VTAIL.n165 VTAIL.n164 0.388379
R820 VTAIL.n121 VTAIL.n120 0.388379
R821 VTAIL.n290 VTAIL.n289 0.155672
R822 VTAIL.n290 VTAIL.n281 0.155672
R823 VTAIL.n297 VTAIL.n281 0.155672
R824 VTAIL.n298 VTAIL.n297 0.155672
R825 VTAIL.n298 VTAIL.n277 0.155672
R826 VTAIL.n305 VTAIL.n277 0.155672
R827 VTAIL.n306 VTAIL.n305 0.155672
R828 VTAIL.n306 VTAIL.n273 0.155672
R829 VTAIL.n313 VTAIL.n273 0.155672
R830 VTAIL.n314 VTAIL.n313 0.155672
R831 VTAIL.n314 VTAIL.n269 0.155672
R832 VTAIL.n321 VTAIL.n269 0.155672
R833 VTAIL.n322 VTAIL.n321 0.155672
R834 VTAIL.n322 VTAIL.n265 0.155672
R835 VTAIL.n330 VTAIL.n265 0.155672
R836 VTAIL.n331 VTAIL.n330 0.155672
R837 VTAIL.n331 VTAIL.n261 0.155672
R838 VTAIL.n339 VTAIL.n261 0.155672
R839 VTAIL.n32 VTAIL.n31 0.155672
R840 VTAIL.n32 VTAIL.n23 0.155672
R841 VTAIL.n39 VTAIL.n23 0.155672
R842 VTAIL.n40 VTAIL.n39 0.155672
R843 VTAIL.n40 VTAIL.n19 0.155672
R844 VTAIL.n47 VTAIL.n19 0.155672
R845 VTAIL.n48 VTAIL.n47 0.155672
R846 VTAIL.n48 VTAIL.n15 0.155672
R847 VTAIL.n55 VTAIL.n15 0.155672
R848 VTAIL.n56 VTAIL.n55 0.155672
R849 VTAIL.n56 VTAIL.n11 0.155672
R850 VTAIL.n63 VTAIL.n11 0.155672
R851 VTAIL.n64 VTAIL.n63 0.155672
R852 VTAIL.n64 VTAIL.n7 0.155672
R853 VTAIL.n72 VTAIL.n7 0.155672
R854 VTAIL.n73 VTAIL.n72 0.155672
R855 VTAIL.n73 VTAIL.n3 0.155672
R856 VTAIL.n81 VTAIL.n3 0.155672
R857 VTAIL.n257 VTAIL.n179 0.155672
R858 VTAIL.n249 VTAIL.n179 0.155672
R859 VTAIL.n249 VTAIL.n248 0.155672
R860 VTAIL.n248 VTAIL.n183 0.155672
R861 VTAIL.n241 VTAIL.n183 0.155672
R862 VTAIL.n241 VTAIL.n240 0.155672
R863 VTAIL.n240 VTAIL.n188 0.155672
R864 VTAIL.n233 VTAIL.n188 0.155672
R865 VTAIL.n233 VTAIL.n232 0.155672
R866 VTAIL.n232 VTAIL.n192 0.155672
R867 VTAIL.n225 VTAIL.n192 0.155672
R868 VTAIL.n225 VTAIL.n224 0.155672
R869 VTAIL.n224 VTAIL.n196 0.155672
R870 VTAIL.n217 VTAIL.n196 0.155672
R871 VTAIL.n217 VTAIL.n216 0.155672
R872 VTAIL.n216 VTAIL.n200 0.155672
R873 VTAIL.n209 VTAIL.n200 0.155672
R874 VTAIL.n209 VTAIL.n208 0.155672
R875 VTAIL.n171 VTAIL.n93 0.155672
R876 VTAIL.n163 VTAIL.n93 0.155672
R877 VTAIL.n163 VTAIL.n162 0.155672
R878 VTAIL.n162 VTAIL.n97 0.155672
R879 VTAIL.n155 VTAIL.n97 0.155672
R880 VTAIL.n155 VTAIL.n154 0.155672
R881 VTAIL.n154 VTAIL.n102 0.155672
R882 VTAIL.n147 VTAIL.n102 0.155672
R883 VTAIL.n147 VTAIL.n146 0.155672
R884 VTAIL.n146 VTAIL.n106 0.155672
R885 VTAIL.n139 VTAIL.n106 0.155672
R886 VTAIL.n139 VTAIL.n138 0.155672
R887 VTAIL.n138 VTAIL.n110 0.155672
R888 VTAIL.n131 VTAIL.n110 0.155672
R889 VTAIL.n131 VTAIL.n130 0.155672
R890 VTAIL.n130 VTAIL.n114 0.155672
R891 VTAIL.n123 VTAIL.n114 0.155672
R892 VTAIL.n123 VTAIL.n122 0.155672
R893 B.n713 B.n712 585
R894 B.n713 B.n86 585
R895 B.n716 B.n715 585
R896 B.n717 B.n145 585
R897 B.n719 B.n718 585
R898 B.n721 B.n144 585
R899 B.n724 B.n723 585
R900 B.n725 B.n143 585
R901 B.n727 B.n726 585
R902 B.n729 B.n142 585
R903 B.n732 B.n731 585
R904 B.n733 B.n141 585
R905 B.n735 B.n734 585
R906 B.n737 B.n140 585
R907 B.n740 B.n739 585
R908 B.n741 B.n139 585
R909 B.n743 B.n742 585
R910 B.n745 B.n138 585
R911 B.n748 B.n747 585
R912 B.n749 B.n137 585
R913 B.n751 B.n750 585
R914 B.n753 B.n136 585
R915 B.n756 B.n755 585
R916 B.n757 B.n135 585
R917 B.n759 B.n758 585
R918 B.n761 B.n134 585
R919 B.n764 B.n763 585
R920 B.n765 B.n133 585
R921 B.n767 B.n766 585
R922 B.n769 B.n132 585
R923 B.n772 B.n771 585
R924 B.n773 B.n131 585
R925 B.n775 B.n774 585
R926 B.n777 B.n130 585
R927 B.n780 B.n779 585
R928 B.n781 B.n129 585
R929 B.n783 B.n782 585
R930 B.n785 B.n128 585
R931 B.n788 B.n787 585
R932 B.n789 B.n127 585
R933 B.n791 B.n790 585
R934 B.n793 B.n126 585
R935 B.n796 B.n795 585
R936 B.n797 B.n125 585
R937 B.n799 B.n798 585
R938 B.n801 B.n124 585
R939 B.n804 B.n803 585
R940 B.n805 B.n123 585
R941 B.n807 B.n806 585
R942 B.n809 B.n122 585
R943 B.n812 B.n811 585
R944 B.n814 B.n119 585
R945 B.n816 B.n815 585
R946 B.n818 B.n118 585
R947 B.n821 B.n820 585
R948 B.n822 B.n117 585
R949 B.n824 B.n823 585
R950 B.n826 B.n116 585
R951 B.n828 B.n827 585
R952 B.n830 B.n829 585
R953 B.n833 B.n832 585
R954 B.n834 B.n111 585
R955 B.n836 B.n835 585
R956 B.n838 B.n110 585
R957 B.n841 B.n840 585
R958 B.n842 B.n109 585
R959 B.n844 B.n843 585
R960 B.n846 B.n108 585
R961 B.n849 B.n848 585
R962 B.n850 B.n107 585
R963 B.n852 B.n851 585
R964 B.n854 B.n106 585
R965 B.n857 B.n856 585
R966 B.n858 B.n105 585
R967 B.n860 B.n859 585
R968 B.n862 B.n104 585
R969 B.n865 B.n864 585
R970 B.n866 B.n103 585
R971 B.n868 B.n867 585
R972 B.n870 B.n102 585
R973 B.n873 B.n872 585
R974 B.n874 B.n101 585
R975 B.n876 B.n875 585
R976 B.n878 B.n100 585
R977 B.n881 B.n880 585
R978 B.n882 B.n99 585
R979 B.n884 B.n883 585
R980 B.n886 B.n98 585
R981 B.n889 B.n888 585
R982 B.n890 B.n97 585
R983 B.n892 B.n891 585
R984 B.n894 B.n96 585
R985 B.n897 B.n896 585
R986 B.n898 B.n95 585
R987 B.n900 B.n899 585
R988 B.n902 B.n94 585
R989 B.n905 B.n904 585
R990 B.n906 B.n93 585
R991 B.n908 B.n907 585
R992 B.n910 B.n92 585
R993 B.n913 B.n912 585
R994 B.n914 B.n91 585
R995 B.n916 B.n915 585
R996 B.n918 B.n90 585
R997 B.n921 B.n920 585
R998 B.n922 B.n89 585
R999 B.n924 B.n923 585
R1000 B.n926 B.n88 585
R1001 B.n929 B.n928 585
R1002 B.n930 B.n87 585
R1003 B.n711 B.n85 585
R1004 B.n933 B.n85 585
R1005 B.n710 B.n84 585
R1006 B.n934 B.n84 585
R1007 B.n709 B.n83 585
R1008 B.n935 B.n83 585
R1009 B.n708 B.n707 585
R1010 B.n707 B.n79 585
R1011 B.n706 B.n78 585
R1012 B.n941 B.n78 585
R1013 B.n705 B.n77 585
R1014 B.n942 B.n77 585
R1015 B.n704 B.n76 585
R1016 B.n943 B.n76 585
R1017 B.n703 B.n702 585
R1018 B.n702 B.n72 585
R1019 B.n701 B.n71 585
R1020 B.n949 B.n71 585
R1021 B.n700 B.n70 585
R1022 B.n950 B.n70 585
R1023 B.n699 B.n69 585
R1024 B.n951 B.n69 585
R1025 B.n698 B.n697 585
R1026 B.n697 B.n65 585
R1027 B.n696 B.n64 585
R1028 B.n957 B.n64 585
R1029 B.n695 B.n63 585
R1030 B.n958 B.n63 585
R1031 B.n694 B.n62 585
R1032 B.n959 B.n62 585
R1033 B.n693 B.n692 585
R1034 B.n692 B.n58 585
R1035 B.n691 B.n57 585
R1036 B.n965 B.n57 585
R1037 B.n690 B.n56 585
R1038 B.n966 B.n56 585
R1039 B.n689 B.n55 585
R1040 B.n967 B.n55 585
R1041 B.n688 B.n687 585
R1042 B.n687 B.n51 585
R1043 B.n686 B.n50 585
R1044 B.n973 B.n50 585
R1045 B.n685 B.n49 585
R1046 B.n974 B.n49 585
R1047 B.n684 B.n48 585
R1048 B.n975 B.n48 585
R1049 B.n683 B.n682 585
R1050 B.n682 B.n44 585
R1051 B.n681 B.n43 585
R1052 B.n981 B.n43 585
R1053 B.n680 B.n42 585
R1054 B.n982 B.n42 585
R1055 B.n679 B.n41 585
R1056 B.n983 B.n41 585
R1057 B.n678 B.n677 585
R1058 B.n677 B.n37 585
R1059 B.n676 B.n36 585
R1060 B.n989 B.n36 585
R1061 B.n675 B.n35 585
R1062 B.n990 B.n35 585
R1063 B.n674 B.n34 585
R1064 B.n991 B.n34 585
R1065 B.n673 B.n672 585
R1066 B.n672 B.n30 585
R1067 B.n671 B.n29 585
R1068 B.n997 B.n29 585
R1069 B.n670 B.n28 585
R1070 B.n998 B.n28 585
R1071 B.n669 B.n27 585
R1072 B.n999 B.n27 585
R1073 B.n668 B.n667 585
R1074 B.n667 B.n26 585
R1075 B.n666 B.n22 585
R1076 B.n1005 B.n22 585
R1077 B.n665 B.n21 585
R1078 B.n1006 B.n21 585
R1079 B.n664 B.n20 585
R1080 B.n1007 B.n20 585
R1081 B.n663 B.n662 585
R1082 B.n662 B.n16 585
R1083 B.n661 B.n15 585
R1084 B.n1013 B.n15 585
R1085 B.n660 B.n14 585
R1086 B.n1014 B.n14 585
R1087 B.n659 B.n13 585
R1088 B.n1015 B.n13 585
R1089 B.n658 B.n657 585
R1090 B.n657 B.n12 585
R1091 B.n656 B.n655 585
R1092 B.n656 B.n8 585
R1093 B.n654 B.n7 585
R1094 B.n1022 B.n7 585
R1095 B.n653 B.n6 585
R1096 B.n1023 B.n6 585
R1097 B.n652 B.n5 585
R1098 B.n1024 B.n5 585
R1099 B.n651 B.n650 585
R1100 B.n650 B.n4 585
R1101 B.n649 B.n146 585
R1102 B.n649 B.n648 585
R1103 B.n639 B.n147 585
R1104 B.n148 B.n147 585
R1105 B.n641 B.n640 585
R1106 B.n642 B.n641 585
R1107 B.n638 B.n152 585
R1108 B.n156 B.n152 585
R1109 B.n637 B.n636 585
R1110 B.n636 B.n635 585
R1111 B.n154 B.n153 585
R1112 B.n155 B.n154 585
R1113 B.n628 B.n627 585
R1114 B.n629 B.n628 585
R1115 B.n626 B.n161 585
R1116 B.n161 B.n160 585
R1117 B.n625 B.n624 585
R1118 B.n624 B.n623 585
R1119 B.n163 B.n162 585
R1120 B.n616 B.n163 585
R1121 B.n615 B.n614 585
R1122 B.n617 B.n615 585
R1123 B.n613 B.n168 585
R1124 B.n168 B.n167 585
R1125 B.n612 B.n611 585
R1126 B.n611 B.n610 585
R1127 B.n170 B.n169 585
R1128 B.n171 B.n170 585
R1129 B.n603 B.n602 585
R1130 B.n604 B.n603 585
R1131 B.n601 B.n176 585
R1132 B.n176 B.n175 585
R1133 B.n600 B.n599 585
R1134 B.n599 B.n598 585
R1135 B.n178 B.n177 585
R1136 B.n179 B.n178 585
R1137 B.n591 B.n590 585
R1138 B.n592 B.n591 585
R1139 B.n589 B.n184 585
R1140 B.n184 B.n183 585
R1141 B.n588 B.n587 585
R1142 B.n587 B.n586 585
R1143 B.n186 B.n185 585
R1144 B.n187 B.n186 585
R1145 B.n579 B.n578 585
R1146 B.n580 B.n579 585
R1147 B.n577 B.n192 585
R1148 B.n192 B.n191 585
R1149 B.n576 B.n575 585
R1150 B.n575 B.n574 585
R1151 B.n194 B.n193 585
R1152 B.n195 B.n194 585
R1153 B.n567 B.n566 585
R1154 B.n568 B.n567 585
R1155 B.n565 B.n200 585
R1156 B.n200 B.n199 585
R1157 B.n564 B.n563 585
R1158 B.n563 B.n562 585
R1159 B.n202 B.n201 585
R1160 B.n203 B.n202 585
R1161 B.n555 B.n554 585
R1162 B.n556 B.n555 585
R1163 B.n553 B.n208 585
R1164 B.n208 B.n207 585
R1165 B.n552 B.n551 585
R1166 B.n551 B.n550 585
R1167 B.n210 B.n209 585
R1168 B.n211 B.n210 585
R1169 B.n543 B.n542 585
R1170 B.n544 B.n543 585
R1171 B.n541 B.n216 585
R1172 B.n216 B.n215 585
R1173 B.n540 B.n539 585
R1174 B.n539 B.n538 585
R1175 B.n218 B.n217 585
R1176 B.n219 B.n218 585
R1177 B.n531 B.n530 585
R1178 B.n532 B.n531 585
R1179 B.n529 B.n224 585
R1180 B.n224 B.n223 585
R1181 B.n528 B.n527 585
R1182 B.n527 B.n526 585
R1183 B.n226 B.n225 585
R1184 B.n227 B.n226 585
R1185 B.n519 B.n518 585
R1186 B.n520 B.n519 585
R1187 B.n517 B.n232 585
R1188 B.n232 B.n231 585
R1189 B.n516 B.n515 585
R1190 B.n515 B.n514 585
R1191 B.n511 B.n236 585
R1192 B.n510 B.n509 585
R1193 B.n507 B.n237 585
R1194 B.n507 B.n235 585
R1195 B.n506 B.n505 585
R1196 B.n504 B.n503 585
R1197 B.n502 B.n239 585
R1198 B.n500 B.n499 585
R1199 B.n498 B.n240 585
R1200 B.n497 B.n496 585
R1201 B.n494 B.n241 585
R1202 B.n492 B.n491 585
R1203 B.n490 B.n242 585
R1204 B.n489 B.n488 585
R1205 B.n486 B.n243 585
R1206 B.n484 B.n483 585
R1207 B.n482 B.n244 585
R1208 B.n481 B.n480 585
R1209 B.n478 B.n245 585
R1210 B.n476 B.n475 585
R1211 B.n474 B.n246 585
R1212 B.n473 B.n472 585
R1213 B.n470 B.n247 585
R1214 B.n468 B.n467 585
R1215 B.n466 B.n248 585
R1216 B.n465 B.n464 585
R1217 B.n462 B.n249 585
R1218 B.n460 B.n459 585
R1219 B.n458 B.n250 585
R1220 B.n457 B.n456 585
R1221 B.n454 B.n251 585
R1222 B.n452 B.n451 585
R1223 B.n450 B.n252 585
R1224 B.n449 B.n448 585
R1225 B.n446 B.n253 585
R1226 B.n444 B.n443 585
R1227 B.n442 B.n254 585
R1228 B.n441 B.n440 585
R1229 B.n438 B.n255 585
R1230 B.n436 B.n435 585
R1231 B.n434 B.n256 585
R1232 B.n433 B.n432 585
R1233 B.n430 B.n257 585
R1234 B.n428 B.n427 585
R1235 B.n426 B.n258 585
R1236 B.n425 B.n424 585
R1237 B.n422 B.n259 585
R1238 B.n420 B.n419 585
R1239 B.n418 B.n260 585
R1240 B.n417 B.n416 585
R1241 B.n414 B.n261 585
R1242 B.n412 B.n411 585
R1243 B.n410 B.n262 585
R1244 B.n409 B.n408 585
R1245 B.n406 B.n266 585
R1246 B.n404 B.n403 585
R1247 B.n402 B.n267 585
R1248 B.n401 B.n400 585
R1249 B.n398 B.n268 585
R1250 B.n396 B.n395 585
R1251 B.n393 B.n269 585
R1252 B.n392 B.n391 585
R1253 B.n389 B.n272 585
R1254 B.n387 B.n386 585
R1255 B.n385 B.n273 585
R1256 B.n384 B.n383 585
R1257 B.n381 B.n274 585
R1258 B.n379 B.n378 585
R1259 B.n377 B.n275 585
R1260 B.n376 B.n375 585
R1261 B.n373 B.n276 585
R1262 B.n371 B.n370 585
R1263 B.n369 B.n277 585
R1264 B.n368 B.n367 585
R1265 B.n365 B.n278 585
R1266 B.n363 B.n362 585
R1267 B.n361 B.n279 585
R1268 B.n360 B.n359 585
R1269 B.n357 B.n280 585
R1270 B.n355 B.n354 585
R1271 B.n353 B.n281 585
R1272 B.n352 B.n351 585
R1273 B.n349 B.n282 585
R1274 B.n347 B.n346 585
R1275 B.n345 B.n283 585
R1276 B.n344 B.n343 585
R1277 B.n341 B.n284 585
R1278 B.n339 B.n338 585
R1279 B.n337 B.n285 585
R1280 B.n336 B.n335 585
R1281 B.n333 B.n286 585
R1282 B.n331 B.n330 585
R1283 B.n329 B.n287 585
R1284 B.n328 B.n327 585
R1285 B.n325 B.n288 585
R1286 B.n323 B.n322 585
R1287 B.n321 B.n289 585
R1288 B.n320 B.n319 585
R1289 B.n317 B.n290 585
R1290 B.n315 B.n314 585
R1291 B.n313 B.n291 585
R1292 B.n312 B.n311 585
R1293 B.n309 B.n292 585
R1294 B.n307 B.n306 585
R1295 B.n305 B.n293 585
R1296 B.n304 B.n303 585
R1297 B.n301 B.n294 585
R1298 B.n299 B.n298 585
R1299 B.n297 B.n296 585
R1300 B.n234 B.n233 585
R1301 B.n513 B.n512 585
R1302 B.n514 B.n513 585
R1303 B.n230 B.n229 585
R1304 B.n231 B.n230 585
R1305 B.n522 B.n521 585
R1306 B.n521 B.n520 585
R1307 B.n523 B.n228 585
R1308 B.n228 B.n227 585
R1309 B.n525 B.n524 585
R1310 B.n526 B.n525 585
R1311 B.n222 B.n221 585
R1312 B.n223 B.n222 585
R1313 B.n534 B.n533 585
R1314 B.n533 B.n532 585
R1315 B.n535 B.n220 585
R1316 B.n220 B.n219 585
R1317 B.n537 B.n536 585
R1318 B.n538 B.n537 585
R1319 B.n214 B.n213 585
R1320 B.n215 B.n214 585
R1321 B.n546 B.n545 585
R1322 B.n545 B.n544 585
R1323 B.n547 B.n212 585
R1324 B.n212 B.n211 585
R1325 B.n549 B.n548 585
R1326 B.n550 B.n549 585
R1327 B.n206 B.n205 585
R1328 B.n207 B.n206 585
R1329 B.n558 B.n557 585
R1330 B.n557 B.n556 585
R1331 B.n559 B.n204 585
R1332 B.n204 B.n203 585
R1333 B.n561 B.n560 585
R1334 B.n562 B.n561 585
R1335 B.n198 B.n197 585
R1336 B.n199 B.n198 585
R1337 B.n570 B.n569 585
R1338 B.n569 B.n568 585
R1339 B.n571 B.n196 585
R1340 B.n196 B.n195 585
R1341 B.n573 B.n572 585
R1342 B.n574 B.n573 585
R1343 B.n190 B.n189 585
R1344 B.n191 B.n190 585
R1345 B.n582 B.n581 585
R1346 B.n581 B.n580 585
R1347 B.n583 B.n188 585
R1348 B.n188 B.n187 585
R1349 B.n585 B.n584 585
R1350 B.n586 B.n585 585
R1351 B.n182 B.n181 585
R1352 B.n183 B.n182 585
R1353 B.n594 B.n593 585
R1354 B.n593 B.n592 585
R1355 B.n595 B.n180 585
R1356 B.n180 B.n179 585
R1357 B.n597 B.n596 585
R1358 B.n598 B.n597 585
R1359 B.n174 B.n173 585
R1360 B.n175 B.n174 585
R1361 B.n606 B.n605 585
R1362 B.n605 B.n604 585
R1363 B.n607 B.n172 585
R1364 B.n172 B.n171 585
R1365 B.n609 B.n608 585
R1366 B.n610 B.n609 585
R1367 B.n166 B.n165 585
R1368 B.n167 B.n166 585
R1369 B.n619 B.n618 585
R1370 B.n618 B.n617 585
R1371 B.n620 B.n164 585
R1372 B.n616 B.n164 585
R1373 B.n622 B.n621 585
R1374 B.n623 B.n622 585
R1375 B.n159 B.n158 585
R1376 B.n160 B.n159 585
R1377 B.n631 B.n630 585
R1378 B.n630 B.n629 585
R1379 B.n632 B.n157 585
R1380 B.n157 B.n155 585
R1381 B.n634 B.n633 585
R1382 B.n635 B.n634 585
R1383 B.n151 B.n150 585
R1384 B.n156 B.n151 585
R1385 B.n644 B.n643 585
R1386 B.n643 B.n642 585
R1387 B.n645 B.n149 585
R1388 B.n149 B.n148 585
R1389 B.n647 B.n646 585
R1390 B.n648 B.n647 585
R1391 B.n3 B.n0 585
R1392 B.n4 B.n3 585
R1393 B.n1021 B.n1 585
R1394 B.n1022 B.n1021 585
R1395 B.n1020 B.n1019 585
R1396 B.n1020 B.n8 585
R1397 B.n1018 B.n9 585
R1398 B.n12 B.n9 585
R1399 B.n1017 B.n1016 585
R1400 B.n1016 B.n1015 585
R1401 B.n11 B.n10 585
R1402 B.n1014 B.n11 585
R1403 B.n1012 B.n1011 585
R1404 B.n1013 B.n1012 585
R1405 B.n1010 B.n17 585
R1406 B.n17 B.n16 585
R1407 B.n1009 B.n1008 585
R1408 B.n1008 B.n1007 585
R1409 B.n19 B.n18 585
R1410 B.n1006 B.n19 585
R1411 B.n1004 B.n1003 585
R1412 B.n1005 B.n1004 585
R1413 B.n1002 B.n23 585
R1414 B.n26 B.n23 585
R1415 B.n1001 B.n1000 585
R1416 B.n1000 B.n999 585
R1417 B.n25 B.n24 585
R1418 B.n998 B.n25 585
R1419 B.n996 B.n995 585
R1420 B.n997 B.n996 585
R1421 B.n994 B.n31 585
R1422 B.n31 B.n30 585
R1423 B.n993 B.n992 585
R1424 B.n992 B.n991 585
R1425 B.n33 B.n32 585
R1426 B.n990 B.n33 585
R1427 B.n988 B.n987 585
R1428 B.n989 B.n988 585
R1429 B.n986 B.n38 585
R1430 B.n38 B.n37 585
R1431 B.n985 B.n984 585
R1432 B.n984 B.n983 585
R1433 B.n40 B.n39 585
R1434 B.n982 B.n40 585
R1435 B.n980 B.n979 585
R1436 B.n981 B.n980 585
R1437 B.n978 B.n45 585
R1438 B.n45 B.n44 585
R1439 B.n977 B.n976 585
R1440 B.n976 B.n975 585
R1441 B.n47 B.n46 585
R1442 B.n974 B.n47 585
R1443 B.n972 B.n971 585
R1444 B.n973 B.n972 585
R1445 B.n970 B.n52 585
R1446 B.n52 B.n51 585
R1447 B.n969 B.n968 585
R1448 B.n968 B.n967 585
R1449 B.n54 B.n53 585
R1450 B.n966 B.n54 585
R1451 B.n964 B.n963 585
R1452 B.n965 B.n964 585
R1453 B.n962 B.n59 585
R1454 B.n59 B.n58 585
R1455 B.n961 B.n960 585
R1456 B.n960 B.n959 585
R1457 B.n61 B.n60 585
R1458 B.n958 B.n61 585
R1459 B.n956 B.n955 585
R1460 B.n957 B.n956 585
R1461 B.n954 B.n66 585
R1462 B.n66 B.n65 585
R1463 B.n953 B.n952 585
R1464 B.n952 B.n951 585
R1465 B.n68 B.n67 585
R1466 B.n950 B.n68 585
R1467 B.n948 B.n947 585
R1468 B.n949 B.n948 585
R1469 B.n946 B.n73 585
R1470 B.n73 B.n72 585
R1471 B.n945 B.n944 585
R1472 B.n944 B.n943 585
R1473 B.n75 B.n74 585
R1474 B.n942 B.n75 585
R1475 B.n940 B.n939 585
R1476 B.n941 B.n940 585
R1477 B.n938 B.n80 585
R1478 B.n80 B.n79 585
R1479 B.n937 B.n936 585
R1480 B.n936 B.n935 585
R1481 B.n82 B.n81 585
R1482 B.n934 B.n82 585
R1483 B.n932 B.n931 585
R1484 B.n933 B.n932 585
R1485 B.n1025 B.n1024 585
R1486 B.n1023 B.n2 585
R1487 B.n932 B.n87 482.89
R1488 B.n713 B.n85 482.89
R1489 B.n515 B.n234 482.89
R1490 B.n513 B.n236 482.89
R1491 B.n112 B.t13 399.709
R1492 B.n120 B.t17 399.709
R1493 B.n270 B.t9 399.709
R1494 B.n263 B.t20 399.709
R1495 B.n112 B.t15 371.524
R1496 B.n120 B.t18 371.524
R1497 B.n270 B.t12 371.524
R1498 B.n263 B.t22 371.524
R1499 B.n121 B.t19 329.44
R1500 B.n271 B.t11 329.44
R1501 B.n113 B.t16 329.44
R1502 B.n264 B.t21 329.44
R1503 B.n714 B.n86 256.663
R1504 B.n720 B.n86 256.663
R1505 B.n722 B.n86 256.663
R1506 B.n728 B.n86 256.663
R1507 B.n730 B.n86 256.663
R1508 B.n736 B.n86 256.663
R1509 B.n738 B.n86 256.663
R1510 B.n744 B.n86 256.663
R1511 B.n746 B.n86 256.663
R1512 B.n752 B.n86 256.663
R1513 B.n754 B.n86 256.663
R1514 B.n760 B.n86 256.663
R1515 B.n762 B.n86 256.663
R1516 B.n768 B.n86 256.663
R1517 B.n770 B.n86 256.663
R1518 B.n776 B.n86 256.663
R1519 B.n778 B.n86 256.663
R1520 B.n784 B.n86 256.663
R1521 B.n786 B.n86 256.663
R1522 B.n792 B.n86 256.663
R1523 B.n794 B.n86 256.663
R1524 B.n800 B.n86 256.663
R1525 B.n802 B.n86 256.663
R1526 B.n808 B.n86 256.663
R1527 B.n810 B.n86 256.663
R1528 B.n817 B.n86 256.663
R1529 B.n819 B.n86 256.663
R1530 B.n825 B.n86 256.663
R1531 B.n115 B.n86 256.663
R1532 B.n831 B.n86 256.663
R1533 B.n837 B.n86 256.663
R1534 B.n839 B.n86 256.663
R1535 B.n845 B.n86 256.663
R1536 B.n847 B.n86 256.663
R1537 B.n853 B.n86 256.663
R1538 B.n855 B.n86 256.663
R1539 B.n861 B.n86 256.663
R1540 B.n863 B.n86 256.663
R1541 B.n869 B.n86 256.663
R1542 B.n871 B.n86 256.663
R1543 B.n877 B.n86 256.663
R1544 B.n879 B.n86 256.663
R1545 B.n885 B.n86 256.663
R1546 B.n887 B.n86 256.663
R1547 B.n893 B.n86 256.663
R1548 B.n895 B.n86 256.663
R1549 B.n901 B.n86 256.663
R1550 B.n903 B.n86 256.663
R1551 B.n909 B.n86 256.663
R1552 B.n911 B.n86 256.663
R1553 B.n917 B.n86 256.663
R1554 B.n919 B.n86 256.663
R1555 B.n925 B.n86 256.663
R1556 B.n927 B.n86 256.663
R1557 B.n508 B.n235 256.663
R1558 B.n238 B.n235 256.663
R1559 B.n501 B.n235 256.663
R1560 B.n495 B.n235 256.663
R1561 B.n493 B.n235 256.663
R1562 B.n487 B.n235 256.663
R1563 B.n485 B.n235 256.663
R1564 B.n479 B.n235 256.663
R1565 B.n477 B.n235 256.663
R1566 B.n471 B.n235 256.663
R1567 B.n469 B.n235 256.663
R1568 B.n463 B.n235 256.663
R1569 B.n461 B.n235 256.663
R1570 B.n455 B.n235 256.663
R1571 B.n453 B.n235 256.663
R1572 B.n447 B.n235 256.663
R1573 B.n445 B.n235 256.663
R1574 B.n439 B.n235 256.663
R1575 B.n437 B.n235 256.663
R1576 B.n431 B.n235 256.663
R1577 B.n429 B.n235 256.663
R1578 B.n423 B.n235 256.663
R1579 B.n421 B.n235 256.663
R1580 B.n415 B.n235 256.663
R1581 B.n413 B.n235 256.663
R1582 B.n407 B.n235 256.663
R1583 B.n405 B.n235 256.663
R1584 B.n399 B.n235 256.663
R1585 B.n397 B.n235 256.663
R1586 B.n390 B.n235 256.663
R1587 B.n388 B.n235 256.663
R1588 B.n382 B.n235 256.663
R1589 B.n380 B.n235 256.663
R1590 B.n374 B.n235 256.663
R1591 B.n372 B.n235 256.663
R1592 B.n366 B.n235 256.663
R1593 B.n364 B.n235 256.663
R1594 B.n358 B.n235 256.663
R1595 B.n356 B.n235 256.663
R1596 B.n350 B.n235 256.663
R1597 B.n348 B.n235 256.663
R1598 B.n342 B.n235 256.663
R1599 B.n340 B.n235 256.663
R1600 B.n334 B.n235 256.663
R1601 B.n332 B.n235 256.663
R1602 B.n326 B.n235 256.663
R1603 B.n324 B.n235 256.663
R1604 B.n318 B.n235 256.663
R1605 B.n316 B.n235 256.663
R1606 B.n310 B.n235 256.663
R1607 B.n308 B.n235 256.663
R1608 B.n302 B.n235 256.663
R1609 B.n300 B.n235 256.663
R1610 B.n295 B.n235 256.663
R1611 B.n1027 B.n1026 256.663
R1612 B.n928 B.n926 163.367
R1613 B.n924 B.n89 163.367
R1614 B.n920 B.n918 163.367
R1615 B.n916 B.n91 163.367
R1616 B.n912 B.n910 163.367
R1617 B.n908 B.n93 163.367
R1618 B.n904 B.n902 163.367
R1619 B.n900 B.n95 163.367
R1620 B.n896 B.n894 163.367
R1621 B.n892 B.n97 163.367
R1622 B.n888 B.n886 163.367
R1623 B.n884 B.n99 163.367
R1624 B.n880 B.n878 163.367
R1625 B.n876 B.n101 163.367
R1626 B.n872 B.n870 163.367
R1627 B.n868 B.n103 163.367
R1628 B.n864 B.n862 163.367
R1629 B.n860 B.n105 163.367
R1630 B.n856 B.n854 163.367
R1631 B.n852 B.n107 163.367
R1632 B.n848 B.n846 163.367
R1633 B.n844 B.n109 163.367
R1634 B.n840 B.n838 163.367
R1635 B.n836 B.n111 163.367
R1636 B.n832 B.n830 163.367
R1637 B.n827 B.n826 163.367
R1638 B.n824 B.n117 163.367
R1639 B.n820 B.n818 163.367
R1640 B.n816 B.n119 163.367
R1641 B.n811 B.n809 163.367
R1642 B.n807 B.n123 163.367
R1643 B.n803 B.n801 163.367
R1644 B.n799 B.n125 163.367
R1645 B.n795 B.n793 163.367
R1646 B.n791 B.n127 163.367
R1647 B.n787 B.n785 163.367
R1648 B.n783 B.n129 163.367
R1649 B.n779 B.n777 163.367
R1650 B.n775 B.n131 163.367
R1651 B.n771 B.n769 163.367
R1652 B.n767 B.n133 163.367
R1653 B.n763 B.n761 163.367
R1654 B.n759 B.n135 163.367
R1655 B.n755 B.n753 163.367
R1656 B.n751 B.n137 163.367
R1657 B.n747 B.n745 163.367
R1658 B.n743 B.n139 163.367
R1659 B.n739 B.n737 163.367
R1660 B.n735 B.n141 163.367
R1661 B.n731 B.n729 163.367
R1662 B.n727 B.n143 163.367
R1663 B.n723 B.n721 163.367
R1664 B.n719 B.n145 163.367
R1665 B.n715 B.n713 163.367
R1666 B.n515 B.n232 163.367
R1667 B.n519 B.n232 163.367
R1668 B.n519 B.n226 163.367
R1669 B.n527 B.n226 163.367
R1670 B.n527 B.n224 163.367
R1671 B.n531 B.n224 163.367
R1672 B.n531 B.n218 163.367
R1673 B.n539 B.n218 163.367
R1674 B.n539 B.n216 163.367
R1675 B.n543 B.n216 163.367
R1676 B.n543 B.n210 163.367
R1677 B.n551 B.n210 163.367
R1678 B.n551 B.n208 163.367
R1679 B.n555 B.n208 163.367
R1680 B.n555 B.n202 163.367
R1681 B.n563 B.n202 163.367
R1682 B.n563 B.n200 163.367
R1683 B.n567 B.n200 163.367
R1684 B.n567 B.n194 163.367
R1685 B.n575 B.n194 163.367
R1686 B.n575 B.n192 163.367
R1687 B.n579 B.n192 163.367
R1688 B.n579 B.n186 163.367
R1689 B.n587 B.n186 163.367
R1690 B.n587 B.n184 163.367
R1691 B.n591 B.n184 163.367
R1692 B.n591 B.n178 163.367
R1693 B.n599 B.n178 163.367
R1694 B.n599 B.n176 163.367
R1695 B.n603 B.n176 163.367
R1696 B.n603 B.n170 163.367
R1697 B.n611 B.n170 163.367
R1698 B.n611 B.n168 163.367
R1699 B.n615 B.n168 163.367
R1700 B.n615 B.n163 163.367
R1701 B.n624 B.n163 163.367
R1702 B.n624 B.n161 163.367
R1703 B.n628 B.n161 163.367
R1704 B.n628 B.n154 163.367
R1705 B.n636 B.n154 163.367
R1706 B.n636 B.n152 163.367
R1707 B.n641 B.n152 163.367
R1708 B.n641 B.n147 163.367
R1709 B.n649 B.n147 163.367
R1710 B.n650 B.n649 163.367
R1711 B.n650 B.n5 163.367
R1712 B.n6 B.n5 163.367
R1713 B.n7 B.n6 163.367
R1714 B.n656 B.n7 163.367
R1715 B.n657 B.n656 163.367
R1716 B.n657 B.n13 163.367
R1717 B.n14 B.n13 163.367
R1718 B.n15 B.n14 163.367
R1719 B.n662 B.n15 163.367
R1720 B.n662 B.n20 163.367
R1721 B.n21 B.n20 163.367
R1722 B.n22 B.n21 163.367
R1723 B.n667 B.n22 163.367
R1724 B.n667 B.n27 163.367
R1725 B.n28 B.n27 163.367
R1726 B.n29 B.n28 163.367
R1727 B.n672 B.n29 163.367
R1728 B.n672 B.n34 163.367
R1729 B.n35 B.n34 163.367
R1730 B.n36 B.n35 163.367
R1731 B.n677 B.n36 163.367
R1732 B.n677 B.n41 163.367
R1733 B.n42 B.n41 163.367
R1734 B.n43 B.n42 163.367
R1735 B.n682 B.n43 163.367
R1736 B.n682 B.n48 163.367
R1737 B.n49 B.n48 163.367
R1738 B.n50 B.n49 163.367
R1739 B.n687 B.n50 163.367
R1740 B.n687 B.n55 163.367
R1741 B.n56 B.n55 163.367
R1742 B.n57 B.n56 163.367
R1743 B.n692 B.n57 163.367
R1744 B.n692 B.n62 163.367
R1745 B.n63 B.n62 163.367
R1746 B.n64 B.n63 163.367
R1747 B.n697 B.n64 163.367
R1748 B.n697 B.n69 163.367
R1749 B.n70 B.n69 163.367
R1750 B.n71 B.n70 163.367
R1751 B.n702 B.n71 163.367
R1752 B.n702 B.n76 163.367
R1753 B.n77 B.n76 163.367
R1754 B.n78 B.n77 163.367
R1755 B.n707 B.n78 163.367
R1756 B.n707 B.n83 163.367
R1757 B.n84 B.n83 163.367
R1758 B.n85 B.n84 163.367
R1759 B.n509 B.n507 163.367
R1760 B.n507 B.n506 163.367
R1761 B.n503 B.n502 163.367
R1762 B.n500 B.n240 163.367
R1763 B.n496 B.n494 163.367
R1764 B.n492 B.n242 163.367
R1765 B.n488 B.n486 163.367
R1766 B.n484 B.n244 163.367
R1767 B.n480 B.n478 163.367
R1768 B.n476 B.n246 163.367
R1769 B.n472 B.n470 163.367
R1770 B.n468 B.n248 163.367
R1771 B.n464 B.n462 163.367
R1772 B.n460 B.n250 163.367
R1773 B.n456 B.n454 163.367
R1774 B.n452 B.n252 163.367
R1775 B.n448 B.n446 163.367
R1776 B.n444 B.n254 163.367
R1777 B.n440 B.n438 163.367
R1778 B.n436 B.n256 163.367
R1779 B.n432 B.n430 163.367
R1780 B.n428 B.n258 163.367
R1781 B.n424 B.n422 163.367
R1782 B.n420 B.n260 163.367
R1783 B.n416 B.n414 163.367
R1784 B.n412 B.n262 163.367
R1785 B.n408 B.n406 163.367
R1786 B.n404 B.n267 163.367
R1787 B.n400 B.n398 163.367
R1788 B.n396 B.n269 163.367
R1789 B.n391 B.n389 163.367
R1790 B.n387 B.n273 163.367
R1791 B.n383 B.n381 163.367
R1792 B.n379 B.n275 163.367
R1793 B.n375 B.n373 163.367
R1794 B.n371 B.n277 163.367
R1795 B.n367 B.n365 163.367
R1796 B.n363 B.n279 163.367
R1797 B.n359 B.n357 163.367
R1798 B.n355 B.n281 163.367
R1799 B.n351 B.n349 163.367
R1800 B.n347 B.n283 163.367
R1801 B.n343 B.n341 163.367
R1802 B.n339 B.n285 163.367
R1803 B.n335 B.n333 163.367
R1804 B.n331 B.n287 163.367
R1805 B.n327 B.n325 163.367
R1806 B.n323 B.n289 163.367
R1807 B.n319 B.n317 163.367
R1808 B.n315 B.n291 163.367
R1809 B.n311 B.n309 163.367
R1810 B.n307 B.n293 163.367
R1811 B.n303 B.n301 163.367
R1812 B.n299 B.n296 163.367
R1813 B.n513 B.n230 163.367
R1814 B.n521 B.n230 163.367
R1815 B.n521 B.n228 163.367
R1816 B.n525 B.n228 163.367
R1817 B.n525 B.n222 163.367
R1818 B.n533 B.n222 163.367
R1819 B.n533 B.n220 163.367
R1820 B.n537 B.n220 163.367
R1821 B.n537 B.n214 163.367
R1822 B.n545 B.n214 163.367
R1823 B.n545 B.n212 163.367
R1824 B.n549 B.n212 163.367
R1825 B.n549 B.n206 163.367
R1826 B.n557 B.n206 163.367
R1827 B.n557 B.n204 163.367
R1828 B.n561 B.n204 163.367
R1829 B.n561 B.n198 163.367
R1830 B.n569 B.n198 163.367
R1831 B.n569 B.n196 163.367
R1832 B.n573 B.n196 163.367
R1833 B.n573 B.n190 163.367
R1834 B.n581 B.n190 163.367
R1835 B.n581 B.n188 163.367
R1836 B.n585 B.n188 163.367
R1837 B.n585 B.n182 163.367
R1838 B.n593 B.n182 163.367
R1839 B.n593 B.n180 163.367
R1840 B.n597 B.n180 163.367
R1841 B.n597 B.n174 163.367
R1842 B.n605 B.n174 163.367
R1843 B.n605 B.n172 163.367
R1844 B.n609 B.n172 163.367
R1845 B.n609 B.n166 163.367
R1846 B.n618 B.n166 163.367
R1847 B.n618 B.n164 163.367
R1848 B.n622 B.n164 163.367
R1849 B.n622 B.n159 163.367
R1850 B.n630 B.n159 163.367
R1851 B.n630 B.n157 163.367
R1852 B.n634 B.n157 163.367
R1853 B.n634 B.n151 163.367
R1854 B.n643 B.n151 163.367
R1855 B.n643 B.n149 163.367
R1856 B.n647 B.n149 163.367
R1857 B.n647 B.n3 163.367
R1858 B.n1025 B.n3 163.367
R1859 B.n1021 B.n2 163.367
R1860 B.n1021 B.n1020 163.367
R1861 B.n1020 B.n9 163.367
R1862 B.n1016 B.n9 163.367
R1863 B.n1016 B.n11 163.367
R1864 B.n1012 B.n11 163.367
R1865 B.n1012 B.n17 163.367
R1866 B.n1008 B.n17 163.367
R1867 B.n1008 B.n19 163.367
R1868 B.n1004 B.n19 163.367
R1869 B.n1004 B.n23 163.367
R1870 B.n1000 B.n23 163.367
R1871 B.n1000 B.n25 163.367
R1872 B.n996 B.n25 163.367
R1873 B.n996 B.n31 163.367
R1874 B.n992 B.n31 163.367
R1875 B.n992 B.n33 163.367
R1876 B.n988 B.n33 163.367
R1877 B.n988 B.n38 163.367
R1878 B.n984 B.n38 163.367
R1879 B.n984 B.n40 163.367
R1880 B.n980 B.n40 163.367
R1881 B.n980 B.n45 163.367
R1882 B.n976 B.n45 163.367
R1883 B.n976 B.n47 163.367
R1884 B.n972 B.n47 163.367
R1885 B.n972 B.n52 163.367
R1886 B.n968 B.n52 163.367
R1887 B.n968 B.n54 163.367
R1888 B.n964 B.n54 163.367
R1889 B.n964 B.n59 163.367
R1890 B.n960 B.n59 163.367
R1891 B.n960 B.n61 163.367
R1892 B.n956 B.n61 163.367
R1893 B.n956 B.n66 163.367
R1894 B.n952 B.n66 163.367
R1895 B.n952 B.n68 163.367
R1896 B.n948 B.n68 163.367
R1897 B.n948 B.n73 163.367
R1898 B.n944 B.n73 163.367
R1899 B.n944 B.n75 163.367
R1900 B.n940 B.n75 163.367
R1901 B.n940 B.n80 163.367
R1902 B.n936 B.n80 163.367
R1903 B.n936 B.n82 163.367
R1904 B.n932 B.n82 163.367
R1905 B.n927 B.n87 71.676
R1906 B.n926 B.n925 71.676
R1907 B.n919 B.n89 71.676
R1908 B.n918 B.n917 71.676
R1909 B.n911 B.n91 71.676
R1910 B.n910 B.n909 71.676
R1911 B.n903 B.n93 71.676
R1912 B.n902 B.n901 71.676
R1913 B.n895 B.n95 71.676
R1914 B.n894 B.n893 71.676
R1915 B.n887 B.n97 71.676
R1916 B.n886 B.n885 71.676
R1917 B.n879 B.n99 71.676
R1918 B.n878 B.n877 71.676
R1919 B.n871 B.n101 71.676
R1920 B.n870 B.n869 71.676
R1921 B.n863 B.n103 71.676
R1922 B.n862 B.n861 71.676
R1923 B.n855 B.n105 71.676
R1924 B.n854 B.n853 71.676
R1925 B.n847 B.n107 71.676
R1926 B.n846 B.n845 71.676
R1927 B.n839 B.n109 71.676
R1928 B.n838 B.n837 71.676
R1929 B.n831 B.n111 71.676
R1930 B.n830 B.n115 71.676
R1931 B.n826 B.n825 71.676
R1932 B.n819 B.n117 71.676
R1933 B.n818 B.n817 71.676
R1934 B.n810 B.n119 71.676
R1935 B.n809 B.n808 71.676
R1936 B.n802 B.n123 71.676
R1937 B.n801 B.n800 71.676
R1938 B.n794 B.n125 71.676
R1939 B.n793 B.n792 71.676
R1940 B.n786 B.n127 71.676
R1941 B.n785 B.n784 71.676
R1942 B.n778 B.n129 71.676
R1943 B.n777 B.n776 71.676
R1944 B.n770 B.n131 71.676
R1945 B.n769 B.n768 71.676
R1946 B.n762 B.n133 71.676
R1947 B.n761 B.n760 71.676
R1948 B.n754 B.n135 71.676
R1949 B.n753 B.n752 71.676
R1950 B.n746 B.n137 71.676
R1951 B.n745 B.n744 71.676
R1952 B.n738 B.n139 71.676
R1953 B.n737 B.n736 71.676
R1954 B.n730 B.n141 71.676
R1955 B.n729 B.n728 71.676
R1956 B.n722 B.n143 71.676
R1957 B.n721 B.n720 71.676
R1958 B.n714 B.n145 71.676
R1959 B.n715 B.n714 71.676
R1960 B.n720 B.n719 71.676
R1961 B.n723 B.n722 71.676
R1962 B.n728 B.n727 71.676
R1963 B.n731 B.n730 71.676
R1964 B.n736 B.n735 71.676
R1965 B.n739 B.n738 71.676
R1966 B.n744 B.n743 71.676
R1967 B.n747 B.n746 71.676
R1968 B.n752 B.n751 71.676
R1969 B.n755 B.n754 71.676
R1970 B.n760 B.n759 71.676
R1971 B.n763 B.n762 71.676
R1972 B.n768 B.n767 71.676
R1973 B.n771 B.n770 71.676
R1974 B.n776 B.n775 71.676
R1975 B.n779 B.n778 71.676
R1976 B.n784 B.n783 71.676
R1977 B.n787 B.n786 71.676
R1978 B.n792 B.n791 71.676
R1979 B.n795 B.n794 71.676
R1980 B.n800 B.n799 71.676
R1981 B.n803 B.n802 71.676
R1982 B.n808 B.n807 71.676
R1983 B.n811 B.n810 71.676
R1984 B.n817 B.n816 71.676
R1985 B.n820 B.n819 71.676
R1986 B.n825 B.n824 71.676
R1987 B.n827 B.n115 71.676
R1988 B.n832 B.n831 71.676
R1989 B.n837 B.n836 71.676
R1990 B.n840 B.n839 71.676
R1991 B.n845 B.n844 71.676
R1992 B.n848 B.n847 71.676
R1993 B.n853 B.n852 71.676
R1994 B.n856 B.n855 71.676
R1995 B.n861 B.n860 71.676
R1996 B.n864 B.n863 71.676
R1997 B.n869 B.n868 71.676
R1998 B.n872 B.n871 71.676
R1999 B.n877 B.n876 71.676
R2000 B.n880 B.n879 71.676
R2001 B.n885 B.n884 71.676
R2002 B.n888 B.n887 71.676
R2003 B.n893 B.n892 71.676
R2004 B.n896 B.n895 71.676
R2005 B.n901 B.n900 71.676
R2006 B.n904 B.n903 71.676
R2007 B.n909 B.n908 71.676
R2008 B.n912 B.n911 71.676
R2009 B.n917 B.n916 71.676
R2010 B.n920 B.n919 71.676
R2011 B.n925 B.n924 71.676
R2012 B.n928 B.n927 71.676
R2013 B.n508 B.n236 71.676
R2014 B.n506 B.n238 71.676
R2015 B.n502 B.n501 71.676
R2016 B.n495 B.n240 71.676
R2017 B.n494 B.n493 71.676
R2018 B.n487 B.n242 71.676
R2019 B.n486 B.n485 71.676
R2020 B.n479 B.n244 71.676
R2021 B.n478 B.n477 71.676
R2022 B.n471 B.n246 71.676
R2023 B.n470 B.n469 71.676
R2024 B.n463 B.n248 71.676
R2025 B.n462 B.n461 71.676
R2026 B.n455 B.n250 71.676
R2027 B.n454 B.n453 71.676
R2028 B.n447 B.n252 71.676
R2029 B.n446 B.n445 71.676
R2030 B.n439 B.n254 71.676
R2031 B.n438 B.n437 71.676
R2032 B.n431 B.n256 71.676
R2033 B.n430 B.n429 71.676
R2034 B.n423 B.n258 71.676
R2035 B.n422 B.n421 71.676
R2036 B.n415 B.n260 71.676
R2037 B.n414 B.n413 71.676
R2038 B.n407 B.n262 71.676
R2039 B.n406 B.n405 71.676
R2040 B.n399 B.n267 71.676
R2041 B.n398 B.n397 71.676
R2042 B.n390 B.n269 71.676
R2043 B.n389 B.n388 71.676
R2044 B.n382 B.n273 71.676
R2045 B.n381 B.n380 71.676
R2046 B.n374 B.n275 71.676
R2047 B.n373 B.n372 71.676
R2048 B.n366 B.n277 71.676
R2049 B.n365 B.n364 71.676
R2050 B.n358 B.n279 71.676
R2051 B.n357 B.n356 71.676
R2052 B.n350 B.n281 71.676
R2053 B.n349 B.n348 71.676
R2054 B.n342 B.n283 71.676
R2055 B.n341 B.n340 71.676
R2056 B.n334 B.n285 71.676
R2057 B.n333 B.n332 71.676
R2058 B.n326 B.n287 71.676
R2059 B.n325 B.n324 71.676
R2060 B.n318 B.n289 71.676
R2061 B.n317 B.n316 71.676
R2062 B.n310 B.n291 71.676
R2063 B.n309 B.n308 71.676
R2064 B.n302 B.n293 71.676
R2065 B.n301 B.n300 71.676
R2066 B.n296 B.n295 71.676
R2067 B.n509 B.n508 71.676
R2068 B.n503 B.n238 71.676
R2069 B.n501 B.n500 71.676
R2070 B.n496 B.n495 71.676
R2071 B.n493 B.n492 71.676
R2072 B.n488 B.n487 71.676
R2073 B.n485 B.n484 71.676
R2074 B.n480 B.n479 71.676
R2075 B.n477 B.n476 71.676
R2076 B.n472 B.n471 71.676
R2077 B.n469 B.n468 71.676
R2078 B.n464 B.n463 71.676
R2079 B.n461 B.n460 71.676
R2080 B.n456 B.n455 71.676
R2081 B.n453 B.n452 71.676
R2082 B.n448 B.n447 71.676
R2083 B.n445 B.n444 71.676
R2084 B.n440 B.n439 71.676
R2085 B.n437 B.n436 71.676
R2086 B.n432 B.n431 71.676
R2087 B.n429 B.n428 71.676
R2088 B.n424 B.n423 71.676
R2089 B.n421 B.n420 71.676
R2090 B.n416 B.n415 71.676
R2091 B.n413 B.n412 71.676
R2092 B.n408 B.n407 71.676
R2093 B.n405 B.n404 71.676
R2094 B.n400 B.n399 71.676
R2095 B.n397 B.n396 71.676
R2096 B.n391 B.n390 71.676
R2097 B.n388 B.n387 71.676
R2098 B.n383 B.n382 71.676
R2099 B.n380 B.n379 71.676
R2100 B.n375 B.n374 71.676
R2101 B.n372 B.n371 71.676
R2102 B.n367 B.n366 71.676
R2103 B.n364 B.n363 71.676
R2104 B.n359 B.n358 71.676
R2105 B.n356 B.n355 71.676
R2106 B.n351 B.n350 71.676
R2107 B.n348 B.n347 71.676
R2108 B.n343 B.n342 71.676
R2109 B.n340 B.n339 71.676
R2110 B.n335 B.n334 71.676
R2111 B.n332 B.n331 71.676
R2112 B.n327 B.n326 71.676
R2113 B.n324 B.n323 71.676
R2114 B.n319 B.n318 71.676
R2115 B.n316 B.n315 71.676
R2116 B.n311 B.n310 71.676
R2117 B.n308 B.n307 71.676
R2118 B.n303 B.n302 71.676
R2119 B.n300 B.n299 71.676
R2120 B.n295 B.n234 71.676
R2121 B.n1026 B.n1025 71.676
R2122 B.n1026 B.n2 71.676
R2123 B.n514 B.n235 64.2702
R2124 B.n933 B.n86 64.2702
R2125 B.n114 B.n113 59.5399
R2126 B.n813 B.n121 59.5399
R2127 B.n394 B.n271 59.5399
R2128 B.n265 B.n264 59.5399
R2129 B.n113 B.n112 42.0853
R2130 B.n121 B.n120 42.0853
R2131 B.n271 B.n270 42.0853
R2132 B.n264 B.n263 42.0853
R2133 B.n514 B.n231 37.3538
R2134 B.n520 B.n231 37.3538
R2135 B.n520 B.n227 37.3538
R2136 B.n526 B.n227 37.3538
R2137 B.n526 B.n223 37.3538
R2138 B.n532 B.n223 37.3538
R2139 B.n538 B.n219 37.3538
R2140 B.n538 B.n215 37.3538
R2141 B.n544 B.n215 37.3538
R2142 B.n544 B.n211 37.3538
R2143 B.n550 B.n211 37.3538
R2144 B.n550 B.n207 37.3538
R2145 B.n556 B.n207 37.3538
R2146 B.n556 B.n203 37.3538
R2147 B.n562 B.n203 37.3538
R2148 B.n568 B.n199 37.3538
R2149 B.n568 B.n195 37.3538
R2150 B.n574 B.n195 37.3538
R2151 B.n574 B.n191 37.3538
R2152 B.n580 B.n191 37.3538
R2153 B.n586 B.n187 37.3538
R2154 B.n586 B.n183 37.3538
R2155 B.n592 B.n183 37.3538
R2156 B.n592 B.n179 37.3538
R2157 B.n598 B.n179 37.3538
R2158 B.n604 B.n175 37.3538
R2159 B.n604 B.n171 37.3538
R2160 B.n610 B.n171 37.3538
R2161 B.n610 B.n167 37.3538
R2162 B.n617 B.n167 37.3538
R2163 B.n617 B.n616 37.3538
R2164 B.n623 B.n160 37.3538
R2165 B.n629 B.n160 37.3538
R2166 B.n629 B.n155 37.3538
R2167 B.n635 B.n155 37.3538
R2168 B.n635 B.n156 37.3538
R2169 B.n642 B.n148 37.3538
R2170 B.n648 B.n148 37.3538
R2171 B.n648 B.n4 37.3538
R2172 B.n1024 B.n4 37.3538
R2173 B.n1024 B.n1023 37.3538
R2174 B.n1023 B.n1022 37.3538
R2175 B.n1022 B.n8 37.3538
R2176 B.n12 B.n8 37.3538
R2177 B.n1015 B.n12 37.3538
R2178 B.n1014 B.n1013 37.3538
R2179 B.n1013 B.n16 37.3538
R2180 B.n1007 B.n16 37.3538
R2181 B.n1007 B.n1006 37.3538
R2182 B.n1006 B.n1005 37.3538
R2183 B.n999 B.n26 37.3538
R2184 B.n999 B.n998 37.3538
R2185 B.n998 B.n997 37.3538
R2186 B.n997 B.n30 37.3538
R2187 B.n991 B.n30 37.3538
R2188 B.n991 B.n990 37.3538
R2189 B.n989 B.n37 37.3538
R2190 B.n983 B.n37 37.3538
R2191 B.n983 B.n982 37.3538
R2192 B.n982 B.n981 37.3538
R2193 B.n981 B.n44 37.3538
R2194 B.n975 B.n974 37.3538
R2195 B.n974 B.n973 37.3538
R2196 B.n973 B.n51 37.3538
R2197 B.n967 B.n51 37.3538
R2198 B.n967 B.n966 37.3538
R2199 B.n965 B.n58 37.3538
R2200 B.n959 B.n58 37.3538
R2201 B.n959 B.n958 37.3538
R2202 B.n958 B.n957 37.3538
R2203 B.n957 B.n65 37.3538
R2204 B.n951 B.n65 37.3538
R2205 B.n951 B.n950 37.3538
R2206 B.n950 B.n949 37.3538
R2207 B.n949 B.n72 37.3538
R2208 B.n943 B.n942 37.3538
R2209 B.n942 B.n941 37.3538
R2210 B.n941 B.n79 37.3538
R2211 B.n935 B.n79 37.3538
R2212 B.n935 B.n934 37.3538
R2213 B.n934 B.n933 37.3538
R2214 B.n598 B.t7 35.1566
R2215 B.t4 B.n989 35.1566
R2216 B.n512 B.n511 31.3761
R2217 B.n516 B.n233 31.3761
R2218 B.n712 B.n711 31.3761
R2219 B.n931 B.n930 31.3761
R2220 B.t23 B.n199 30.762
R2221 B.n966 B.t6 30.762
R2222 B.n156 B.t1 26.3675
R2223 B.t2 B.n1014 26.3675
R2224 B.n623 B.t3 25.2689
R2225 B.n1005 B.t5 25.2689
R2226 B.n532 B.t10 21.973
R2227 B.n943 B.t14 21.973
R2228 B.n580 B.t0 20.8744
R2229 B.n975 B.t8 20.8744
R2230 B B.n1027 18.0485
R2231 B.t0 B.n187 16.4799
R2232 B.t8 B.n44 16.4799
R2233 B.t10 B.n219 15.3813
R2234 B.t14 B.n72 15.3813
R2235 B.n616 B.t3 12.0854
R2236 B.n26 B.t5 12.0854
R2237 B.n642 B.t1 10.9868
R2238 B.n1015 B.t2 10.9868
R2239 B.n512 B.n229 10.6151
R2240 B.n522 B.n229 10.6151
R2241 B.n523 B.n522 10.6151
R2242 B.n524 B.n523 10.6151
R2243 B.n524 B.n221 10.6151
R2244 B.n534 B.n221 10.6151
R2245 B.n535 B.n534 10.6151
R2246 B.n536 B.n535 10.6151
R2247 B.n536 B.n213 10.6151
R2248 B.n546 B.n213 10.6151
R2249 B.n547 B.n546 10.6151
R2250 B.n548 B.n547 10.6151
R2251 B.n548 B.n205 10.6151
R2252 B.n558 B.n205 10.6151
R2253 B.n559 B.n558 10.6151
R2254 B.n560 B.n559 10.6151
R2255 B.n560 B.n197 10.6151
R2256 B.n570 B.n197 10.6151
R2257 B.n571 B.n570 10.6151
R2258 B.n572 B.n571 10.6151
R2259 B.n572 B.n189 10.6151
R2260 B.n582 B.n189 10.6151
R2261 B.n583 B.n582 10.6151
R2262 B.n584 B.n583 10.6151
R2263 B.n584 B.n181 10.6151
R2264 B.n594 B.n181 10.6151
R2265 B.n595 B.n594 10.6151
R2266 B.n596 B.n595 10.6151
R2267 B.n596 B.n173 10.6151
R2268 B.n606 B.n173 10.6151
R2269 B.n607 B.n606 10.6151
R2270 B.n608 B.n607 10.6151
R2271 B.n608 B.n165 10.6151
R2272 B.n619 B.n165 10.6151
R2273 B.n620 B.n619 10.6151
R2274 B.n621 B.n620 10.6151
R2275 B.n621 B.n158 10.6151
R2276 B.n631 B.n158 10.6151
R2277 B.n632 B.n631 10.6151
R2278 B.n633 B.n632 10.6151
R2279 B.n633 B.n150 10.6151
R2280 B.n644 B.n150 10.6151
R2281 B.n645 B.n644 10.6151
R2282 B.n646 B.n645 10.6151
R2283 B.n646 B.n0 10.6151
R2284 B.n511 B.n510 10.6151
R2285 B.n510 B.n237 10.6151
R2286 B.n505 B.n237 10.6151
R2287 B.n505 B.n504 10.6151
R2288 B.n504 B.n239 10.6151
R2289 B.n499 B.n239 10.6151
R2290 B.n499 B.n498 10.6151
R2291 B.n498 B.n497 10.6151
R2292 B.n497 B.n241 10.6151
R2293 B.n491 B.n241 10.6151
R2294 B.n491 B.n490 10.6151
R2295 B.n490 B.n489 10.6151
R2296 B.n489 B.n243 10.6151
R2297 B.n483 B.n243 10.6151
R2298 B.n483 B.n482 10.6151
R2299 B.n482 B.n481 10.6151
R2300 B.n481 B.n245 10.6151
R2301 B.n475 B.n245 10.6151
R2302 B.n475 B.n474 10.6151
R2303 B.n474 B.n473 10.6151
R2304 B.n473 B.n247 10.6151
R2305 B.n467 B.n247 10.6151
R2306 B.n467 B.n466 10.6151
R2307 B.n466 B.n465 10.6151
R2308 B.n465 B.n249 10.6151
R2309 B.n459 B.n249 10.6151
R2310 B.n459 B.n458 10.6151
R2311 B.n458 B.n457 10.6151
R2312 B.n457 B.n251 10.6151
R2313 B.n451 B.n251 10.6151
R2314 B.n451 B.n450 10.6151
R2315 B.n450 B.n449 10.6151
R2316 B.n449 B.n253 10.6151
R2317 B.n443 B.n253 10.6151
R2318 B.n443 B.n442 10.6151
R2319 B.n442 B.n441 10.6151
R2320 B.n441 B.n255 10.6151
R2321 B.n435 B.n255 10.6151
R2322 B.n435 B.n434 10.6151
R2323 B.n434 B.n433 10.6151
R2324 B.n433 B.n257 10.6151
R2325 B.n427 B.n257 10.6151
R2326 B.n427 B.n426 10.6151
R2327 B.n426 B.n425 10.6151
R2328 B.n425 B.n259 10.6151
R2329 B.n419 B.n259 10.6151
R2330 B.n419 B.n418 10.6151
R2331 B.n418 B.n417 10.6151
R2332 B.n417 B.n261 10.6151
R2333 B.n411 B.n410 10.6151
R2334 B.n410 B.n409 10.6151
R2335 B.n409 B.n266 10.6151
R2336 B.n403 B.n266 10.6151
R2337 B.n403 B.n402 10.6151
R2338 B.n402 B.n401 10.6151
R2339 B.n401 B.n268 10.6151
R2340 B.n395 B.n268 10.6151
R2341 B.n393 B.n392 10.6151
R2342 B.n392 B.n272 10.6151
R2343 B.n386 B.n272 10.6151
R2344 B.n386 B.n385 10.6151
R2345 B.n385 B.n384 10.6151
R2346 B.n384 B.n274 10.6151
R2347 B.n378 B.n274 10.6151
R2348 B.n378 B.n377 10.6151
R2349 B.n377 B.n376 10.6151
R2350 B.n376 B.n276 10.6151
R2351 B.n370 B.n276 10.6151
R2352 B.n370 B.n369 10.6151
R2353 B.n369 B.n368 10.6151
R2354 B.n368 B.n278 10.6151
R2355 B.n362 B.n278 10.6151
R2356 B.n362 B.n361 10.6151
R2357 B.n361 B.n360 10.6151
R2358 B.n360 B.n280 10.6151
R2359 B.n354 B.n280 10.6151
R2360 B.n354 B.n353 10.6151
R2361 B.n353 B.n352 10.6151
R2362 B.n352 B.n282 10.6151
R2363 B.n346 B.n282 10.6151
R2364 B.n346 B.n345 10.6151
R2365 B.n345 B.n344 10.6151
R2366 B.n344 B.n284 10.6151
R2367 B.n338 B.n284 10.6151
R2368 B.n338 B.n337 10.6151
R2369 B.n337 B.n336 10.6151
R2370 B.n336 B.n286 10.6151
R2371 B.n330 B.n286 10.6151
R2372 B.n330 B.n329 10.6151
R2373 B.n329 B.n328 10.6151
R2374 B.n328 B.n288 10.6151
R2375 B.n322 B.n288 10.6151
R2376 B.n322 B.n321 10.6151
R2377 B.n321 B.n320 10.6151
R2378 B.n320 B.n290 10.6151
R2379 B.n314 B.n290 10.6151
R2380 B.n314 B.n313 10.6151
R2381 B.n313 B.n312 10.6151
R2382 B.n312 B.n292 10.6151
R2383 B.n306 B.n292 10.6151
R2384 B.n306 B.n305 10.6151
R2385 B.n305 B.n304 10.6151
R2386 B.n304 B.n294 10.6151
R2387 B.n298 B.n294 10.6151
R2388 B.n298 B.n297 10.6151
R2389 B.n297 B.n233 10.6151
R2390 B.n517 B.n516 10.6151
R2391 B.n518 B.n517 10.6151
R2392 B.n518 B.n225 10.6151
R2393 B.n528 B.n225 10.6151
R2394 B.n529 B.n528 10.6151
R2395 B.n530 B.n529 10.6151
R2396 B.n530 B.n217 10.6151
R2397 B.n540 B.n217 10.6151
R2398 B.n541 B.n540 10.6151
R2399 B.n542 B.n541 10.6151
R2400 B.n542 B.n209 10.6151
R2401 B.n552 B.n209 10.6151
R2402 B.n553 B.n552 10.6151
R2403 B.n554 B.n553 10.6151
R2404 B.n554 B.n201 10.6151
R2405 B.n564 B.n201 10.6151
R2406 B.n565 B.n564 10.6151
R2407 B.n566 B.n565 10.6151
R2408 B.n566 B.n193 10.6151
R2409 B.n576 B.n193 10.6151
R2410 B.n577 B.n576 10.6151
R2411 B.n578 B.n577 10.6151
R2412 B.n578 B.n185 10.6151
R2413 B.n588 B.n185 10.6151
R2414 B.n589 B.n588 10.6151
R2415 B.n590 B.n589 10.6151
R2416 B.n590 B.n177 10.6151
R2417 B.n600 B.n177 10.6151
R2418 B.n601 B.n600 10.6151
R2419 B.n602 B.n601 10.6151
R2420 B.n602 B.n169 10.6151
R2421 B.n612 B.n169 10.6151
R2422 B.n613 B.n612 10.6151
R2423 B.n614 B.n613 10.6151
R2424 B.n614 B.n162 10.6151
R2425 B.n625 B.n162 10.6151
R2426 B.n626 B.n625 10.6151
R2427 B.n627 B.n626 10.6151
R2428 B.n627 B.n153 10.6151
R2429 B.n637 B.n153 10.6151
R2430 B.n638 B.n637 10.6151
R2431 B.n640 B.n638 10.6151
R2432 B.n640 B.n639 10.6151
R2433 B.n639 B.n146 10.6151
R2434 B.n651 B.n146 10.6151
R2435 B.n652 B.n651 10.6151
R2436 B.n653 B.n652 10.6151
R2437 B.n654 B.n653 10.6151
R2438 B.n655 B.n654 10.6151
R2439 B.n658 B.n655 10.6151
R2440 B.n659 B.n658 10.6151
R2441 B.n660 B.n659 10.6151
R2442 B.n661 B.n660 10.6151
R2443 B.n663 B.n661 10.6151
R2444 B.n664 B.n663 10.6151
R2445 B.n665 B.n664 10.6151
R2446 B.n666 B.n665 10.6151
R2447 B.n668 B.n666 10.6151
R2448 B.n669 B.n668 10.6151
R2449 B.n670 B.n669 10.6151
R2450 B.n671 B.n670 10.6151
R2451 B.n673 B.n671 10.6151
R2452 B.n674 B.n673 10.6151
R2453 B.n675 B.n674 10.6151
R2454 B.n676 B.n675 10.6151
R2455 B.n678 B.n676 10.6151
R2456 B.n679 B.n678 10.6151
R2457 B.n680 B.n679 10.6151
R2458 B.n681 B.n680 10.6151
R2459 B.n683 B.n681 10.6151
R2460 B.n684 B.n683 10.6151
R2461 B.n685 B.n684 10.6151
R2462 B.n686 B.n685 10.6151
R2463 B.n688 B.n686 10.6151
R2464 B.n689 B.n688 10.6151
R2465 B.n690 B.n689 10.6151
R2466 B.n691 B.n690 10.6151
R2467 B.n693 B.n691 10.6151
R2468 B.n694 B.n693 10.6151
R2469 B.n695 B.n694 10.6151
R2470 B.n696 B.n695 10.6151
R2471 B.n698 B.n696 10.6151
R2472 B.n699 B.n698 10.6151
R2473 B.n700 B.n699 10.6151
R2474 B.n701 B.n700 10.6151
R2475 B.n703 B.n701 10.6151
R2476 B.n704 B.n703 10.6151
R2477 B.n705 B.n704 10.6151
R2478 B.n706 B.n705 10.6151
R2479 B.n708 B.n706 10.6151
R2480 B.n709 B.n708 10.6151
R2481 B.n710 B.n709 10.6151
R2482 B.n711 B.n710 10.6151
R2483 B.n1019 B.n1 10.6151
R2484 B.n1019 B.n1018 10.6151
R2485 B.n1018 B.n1017 10.6151
R2486 B.n1017 B.n10 10.6151
R2487 B.n1011 B.n10 10.6151
R2488 B.n1011 B.n1010 10.6151
R2489 B.n1010 B.n1009 10.6151
R2490 B.n1009 B.n18 10.6151
R2491 B.n1003 B.n18 10.6151
R2492 B.n1003 B.n1002 10.6151
R2493 B.n1002 B.n1001 10.6151
R2494 B.n1001 B.n24 10.6151
R2495 B.n995 B.n24 10.6151
R2496 B.n995 B.n994 10.6151
R2497 B.n994 B.n993 10.6151
R2498 B.n993 B.n32 10.6151
R2499 B.n987 B.n32 10.6151
R2500 B.n987 B.n986 10.6151
R2501 B.n986 B.n985 10.6151
R2502 B.n985 B.n39 10.6151
R2503 B.n979 B.n39 10.6151
R2504 B.n979 B.n978 10.6151
R2505 B.n978 B.n977 10.6151
R2506 B.n977 B.n46 10.6151
R2507 B.n971 B.n46 10.6151
R2508 B.n971 B.n970 10.6151
R2509 B.n970 B.n969 10.6151
R2510 B.n969 B.n53 10.6151
R2511 B.n963 B.n53 10.6151
R2512 B.n963 B.n962 10.6151
R2513 B.n962 B.n961 10.6151
R2514 B.n961 B.n60 10.6151
R2515 B.n955 B.n60 10.6151
R2516 B.n955 B.n954 10.6151
R2517 B.n954 B.n953 10.6151
R2518 B.n953 B.n67 10.6151
R2519 B.n947 B.n67 10.6151
R2520 B.n947 B.n946 10.6151
R2521 B.n946 B.n945 10.6151
R2522 B.n945 B.n74 10.6151
R2523 B.n939 B.n74 10.6151
R2524 B.n939 B.n938 10.6151
R2525 B.n938 B.n937 10.6151
R2526 B.n937 B.n81 10.6151
R2527 B.n931 B.n81 10.6151
R2528 B.n930 B.n929 10.6151
R2529 B.n929 B.n88 10.6151
R2530 B.n923 B.n88 10.6151
R2531 B.n923 B.n922 10.6151
R2532 B.n922 B.n921 10.6151
R2533 B.n921 B.n90 10.6151
R2534 B.n915 B.n90 10.6151
R2535 B.n915 B.n914 10.6151
R2536 B.n914 B.n913 10.6151
R2537 B.n913 B.n92 10.6151
R2538 B.n907 B.n92 10.6151
R2539 B.n907 B.n906 10.6151
R2540 B.n906 B.n905 10.6151
R2541 B.n905 B.n94 10.6151
R2542 B.n899 B.n94 10.6151
R2543 B.n899 B.n898 10.6151
R2544 B.n898 B.n897 10.6151
R2545 B.n897 B.n96 10.6151
R2546 B.n891 B.n96 10.6151
R2547 B.n891 B.n890 10.6151
R2548 B.n890 B.n889 10.6151
R2549 B.n889 B.n98 10.6151
R2550 B.n883 B.n98 10.6151
R2551 B.n883 B.n882 10.6151
R2552 B.n882 B.n881 10.6151
R2553 B.n881 B.n100 10.6151
R2554 B.n875 B.n100 10.6151
R2555 B.n875 B.n874 10.6151
R2556 B.n874 B.n873 10.6151
R2557 B.n873 B.n102 10.6151
R2558 B.n867 B.n102 10.6151
R2559 B.n867 B.n866 10.6151
R2560 B.n866 B.n865 10.6151
R2561 B.n865 B.n104 10.6151
R2562 B.n859 B.n104 10.6151
R2563 B.n859 B.n858 10.6151
R2564 B.n858 B.n857 10.6151
R2565 B.n857 B.n106 10.6151
R2566 B.n851 B.n106 10.6151
R2567 B.n851 B.n850 10.6151
R2568 B.n850 B.n849 10.6151
R2569 B.n849 B.n108 10.6151
R2570 B.n843 B.n108 10.6151
R2571 B.n843 B.n842 10.6151
R2572 B.n842 B.n841 10.6151
R2573 B.n841 B.n110 10.6151
R2574 B.n835 B.n110 10.6151
R2575 B.n835 B.n834 10.6151
R2576 B.n834 B.n833 10.6151
R2577 B.n829 B.n828 10.6151
R2578 B.n828 B.n116 10.6151
R2579 B.n823 B.n116 10.6151
R2580 B.n823 B.n822 10.6151
R2581 B.n822 B.n821 10.6151
R2582 B.n821 B.n118 10.6151
R2583 B.n815 B.n118 10.6151
R2584 B.n815 B.n814 10.6151
R2585 B.n812 B.n122 10.6151
R2586 B.n806 B.n122 10.6151
R2587 B.n806 B.n805 10.6151
R2588 B.n805 B.n804 10.6151
R2589 B.n804 B.n124 10.6151
R2590 B.n798 B.n124 10.6151
R2591 B.n798 B.n797 10.6151
R2592 B.n797 B.n796 10.6151
R2593 B.n796 B.n126 10.6151
R2594 B.n790 B.n126 10.6151
R2595 B.n790 B.n789 10.6151
R2596 B.n789 B.n788 10.6151
R2597 B.n788 B.n128 10.6151
R2598 B.n782 B.n128 10.6151
R2599 B.n782 B.n781 10.6151
R2600 B.n781 B.n780 10.6151
R2601 B.n780 B.n130 10.6151
R2602 B.n774 B.n130 10.6151
R2603 B.n774 B.n773 10.6151
R2604 B.n773 B.n772 10.6151
R2605 B.n772 B.n132 10.6151
R2606 B.n766 B.n132 10.6151
R2607 B.n766 B.n765 10.6151
R2608 B.n765 B.n764 10.6151
R2609 B.n764 B.n134 10.6151
R2610 B.n758 B.n134 10.6151
R2611 B.n758 B.n757 10.6151
R2612 B.n757 B.n756 10.6151
R2613 B.n756 B.n136 10.6151
R2614 B.n750 B.n136 10.6151
R2615 B.n750 B.n749 10.6151
R2616 B.n749 B.n748 10.6151
R2617 B.n748 B.n138 10.6151
R2618 B.n742 B.n138 10.6151
R2619 B.n742 B.n741 10.6151
R2620 B.n741 B.n740 10.6151
R2621 B.n740 B.n140 10.6151
R2622 B.n734 B.n140 10.6151
R2623 B.n734 B.n733 10.6151
R2624 B.n733 B.n732 10.6151
R2625 B.n732 B.n142 10.6151
R2626 B.n726 B.n142 10.6151
R2627 B.n726 B.n725 10.6151
R2628 B.n725 B.n724 10.6151
R2629 B.n724 B.n144 10.6151
R2630 B.n718 B.n144 10.6151
R2631 B.n718 B.n717 10.6151
R2632 B.n717 B.n716 10.6151
R2633 B.n716 B.n712 10.6151
R2634 B.n1027 B.n0 8.11757
R2635 B.n1027 B.n1 8.11757
R2636 B.n562 B.t23 6.59226
R2637 B.t6 B.n965 6.59226
R2638 B.n411 B.n265 6.5566
R2639 B.n395 B.n394 6.5566
R2640 B.n829 B.n114 6.5566
R2641 B.n814 B.n813 6.5566
R2642 B.n265 B.n261 4.05904
R2643 B.n394 B.n393 4.05904
R2644 B.n833 B.n114 4.05904
R2645 B.n813 B.n812 4.05904
R2646 B.t7 B.n175 2.19775
R2647 B.n990 B.t4 2.19775
R2648 VP.n17 VP.t8 228.012
R2649 VP.n9 VP.t3 193.194
R2650 VP.n51 VP.t7 193.194
R2651 VP.n58 VP.t9 193.194
R2652 VP.n65 VP.t2 193.194
R2653 VP.n73 VP.t6 193.194
R2654 VP.n40 VP.t5 193.194
R2655 VP.n32 VP.t0 193.194
R2656 VP.n25 VP.t1 193.194
R2657 VP.n18 VP.t4 193.194
R2658 VP.n42 VP.n9 181.363
R2659 VP.n74 VP.n73 181.363
R2660 VP.n41 VP.n40 181.363
R2661 VP.n19 VP.n16 161.3
R2662 VP.n21 VP.n20 161.3
R2663 VP.n22 VP.n15 161.3
R2664 VP.n24 VP.n23 161.3
R2665 VP.n26 VP.n14 161.3
R2666 VP.n28 VP.n27 161.3
R2667 VP.n29 VP.n13 161.3
R2668 VP.n31 VP.n30 161.3
R2669 VP.n33 VP.n12 161.3
R2670 VP.n35 VP.n34 161.3
R2671 VP.n36 VP.n11 161.3
R2672 VP.n38 VP.n37 161.3
R2673 VP.n39 VP.n10 161.3
R2674 VP.n72 VP.n0 161.3
R2675 VP.n71 VP.n70 161.3
R2676 VP.n69 VP.n1 161.3
R2677 VP.n68 VP.n67 161.3
R2678 VP.n66 VP.n2 161.3
R2679 VP.n64 VP.n63 161.3
R2680 VP.n62 VP.n3 161.3
R2681 VP.n61 VP.n60 161.3
R2682 VP.n59 VP.n4 161.3
R2683 VP.n57 VP.n56 161.3
R2684 VP.n55 VP.n5 161.3
R2685 VP.n54 VP.n53 161.3
R2686 VP.n52 VP.n6 161.3
R2687 VP.n50 VP.n49 161.3
R2688 VP.n48 VP.n7 161.3
R2689 VP.n47 VP.n46 161.3
R2690 VP.n45 VP.n8 161.3
R2691 VP.n44 VP.n43 161.3
R2692 VP.n53 VP.n5 56.5193
R2693 VP.n60 VP.n3 56.5193
R2694 VP.n27 VP.n13 56.5193
R2695 VP.n20 VP.n15 56.5193
R2696 VP.n42 VP.n41 50.9891
R2697 VP.n18 VP.n17 48.825
R2698 VP.n46 VP.n45 40.979
R2699 VP.n71 VP.n1 40.979
R2700 VP.n38 VP.n11 40.979
R2701 VP.n46 VP.n7 40.0078
R2702 VP.n67 VP.n1 40.0078
R2703 VP.n34 VP.n11 40.0078
R2704 VP.n45 VP.n44 24.4675
R2705 VP.n50 VP.n7 24.4675
R2706 VP.n53 VP.n52 24.4675
R2707 VP.n57 VP.n5 24.4675
R2708 VP.n60 VP.n59 24.4675
R2709 VP.n64 VP.n3 24.4675
R2710 VP.n67 VP.n66 24.4675
R2711 VP.n72 VP.n71 24.4675
R2712 VP.n39 VP.n38 24.4675
R2713 VP.n31 VP.n13 24.4675
R2714 VP.n34 VP.n33 24.4675
R2715 VP.n24 VP.n15 24.4675
R2716 VP.n27 VP.n26 24.4675
R2717 VP.n20 VP.n19 24.4675
R2718 VP.n52 VP.n51 20.5528
R2719 VP.n65 VP.n64 20.5528
R2720 VP.n32 VP.n31 20.5528
R2721 VP.n19 VP.n18 20.5528
R2722 VP.n17 VP.n16 12.2488
R2723 VP.n58 VP.n57 12.234
R2724 VP.n59 VP.n58 12.234
R2725 VP.n25 VP.n24 12.234
R2726 VP.n26 VP.n25 12.234
R2727 VP.n44 VP.n9 4.40456
R2728 VP.n73 VP.n72 4.40456
R2729 VP.n40 VP.n39 4.40456
R2730 VP.n51 VP.n50 3.91522
R2731 VP.n66 VP.n65 3.91522
R2732 VP.n33 VP.n32 3.91522
R2733 VP.n21 VP.n16 0.189894
R2734 VP.n22 VP.n21 0.189894
R2735 VP.n23 VP.n22 0.189894
R2736 VP.n23 VP.n14 0.189894
R2737 VP.n28 VP.n14 0.189894
R2738 VP.n29 VP.n28 0.189894
R2739 VP.n30 VP.n29 0.189894
R2740 VP.n30 VP.n12 0.189894
R2741 VP.n35 VP.n12 0.189894
R2742 VP.n36 VP.n35 0.189894
R2743 VP.n37 VP.n36 0.189894
R2744 VP.n37 VP.n10 0.189894
R2745 VP.n41 VP.n10 0.189894
R2746 VP.n43 VP.n42 0.189894
R2747 VP.n43 VP.n8 0.189894
R2748 VP.n47 VP.n8 0.189894
R2749 VP.n48 VP.n47 0.189894
R2750 VP.n49 VP.n48 0.189894
R2751 VP.n49 VP.n6 0.189894
R2752 VP.n54 VP.n6 0.189894
R2753 VP.n55 VP.n54 0.189894
R2754 VP.n56 VP.n55 0.189894
R2755 VP.n56 VP.n4 0.189894
R2756 VP.n61 VP.n4 0.189894
R2757 VP.n62 VP.n61 0.189894
R2758 VP.n63 VP.n62 0.189894
R2759 VP.n63 VP.n2 0.189894
R2760 VP.n68 VP.n2 0.189894
R2761 VP.n69 VP.n68 0.189894
R2762 VP.n70 VP.n69 0.189894
R2763 VP.n70 VP.n0 0.189894
R2764 VP.n74 VP.n0 0.189894
R2765 VP VP.n74 0.0516364
R2766 VDD1.n76 VDD1.n0 289.615
R2767 VDD1.n159 VDD1.n83 289.615
R2768 VDD1.n77 VDD1.n76 185
R2769 VDD1.n75 VDD1.n74 185
R2770 VDD1.n73 VDD1.n3 185
R2771 VDD1.n7 VDD1.n4 185
R2772 VDD1.n68 VDD1.n67 185
R2773 VDD1.n66 VDD1.n65 185
R2774 VDD1.n9 VDD1.n8 185
R2775 VDD1.n60 VDD1.n59 185
R2776 VDD1.n58 VDD1.n57 185
R2777 VDD1.n13 VDD1.n12 185
R2778 VDD1.n52 VDD1.n51 185
R2779 VDD1.n50 VDD1.n49 185
R2780 VDD1.n17 VDD1.n16 185
R2781 VDD1.n44 VDD1.n43 185
R2782 VDD1.n42 VDD1.n41 185
R2783 VDD1.n21 VDD1.n20 185
R2784 VDD1.n36 VDD1.n35 185
R2785 VDD1.n34 VDD1.n33 185
R2786 VDD1.n25 VDD1.n24 185
R2787 VDD1.n28 VDD1.n27 185
R2788 VDD1.n110 VDD1.n109 185
R2789 VDD1.n107 VDD1.n106 185
R2790 VDD1.n116 VDD1.n115 185
R2791 VDD1.n118 VDD1.n117 185
R2792 VDD1.n103 VDD1.n102 185
R2793 VDD1.n124 VDD1.n123 185
R2794 VDD1.n126 VDD1.n125 185
R2795 VDD1.n99 VDD1.n98 185
R2796 VDD1.n132 VDD1.n131 185
R2797 VDD1.n134 VDD1.n133 185
R2798 VDD1.n95 VDD1.n94 185
R2799 VDD1.n140 VDD1.n139 185
R2800 VDD1.n142 VDD1.n141 185
R2801 VDD1.n91 VDD1.n90 185
R2802 VDD1.n148 VDD1.n147 185
R2803 VDD1.n151 VDD1.n150 185
R2804 VDD1.n149 VDD1.n87 185
R2805 VDD1.n156 VDD1.n86 185
R2806 VDD1.n158 VDD1.n157 185
R2807 VDD1.n160 VDD1.n159 185
R2808 VDD1.t1 VDD1.n26 147.659
R2809 VDD1.t6 VDD1.n108 147.659
R2810 VDD1.n76 VDD1.n75 104.615
R2811 VDD1.n75 VDD1.n3 104.615
R2812 VDD1.n7 VDD1.n3 104.615
R2813 VDD1.n67 VDD1.n7 104.615
R2814 VDD1.n67 VDD1.n66 104.615
R2815 VDD1.n66 VDD1.n8 104.615
R2816 VDD1.n59 VDD1.n8 104.615
R2817 VDD1.n59 VDD1.n58 104.615
R2818 VDD1.n58 VDD1.n12 104.615
R2819 VDD1.n51 VDD1.n12 104.615
R2820 VDD1.n51 VDD1.n50 104.615
R2821 VDD1.n50 VDD1.n16 104.615
R2822 VDD1.n43 VDD1.n16 104.615
R2823 VDD1.n43 VDD1.n42 104.615
R2824 VDD1.n42 VDD1.n20 104.615
R2825 VDD1.n35 VDD1.n20 104.615
R2826 VDD1.n35 VDD1.n34 104.615
R2827 VDD1.n34 VDD1.n24 104.615
R2828 VDD1.n27 VDD1.n24 104.615
R2829 VDD1.n109 VDD1.n106 104.615
R2830 VDD1.n116 VDD1.n106 104.615
R2831 VDD1.n117 VDD1.n116 104.615
R2832 VDD1.n117 VDD1.n102 104.615
R2833 VDD1.n124 VDD1.n102 104.615
R2834 VDD1.n125 VDD1.n124 104.615
R2835 VDD1.n125 VDD1.n98 104.615
R2836 VDD1.n132 VDD1.n98 104.615
R2837 VDD1.n133 VDD1.n132 104.615
R2838 VDD1.n133 VDD1.n94 104.615
R2839 VDD1.n140 VDD1.n94 104.615
R2840 VDD1.n141 VDD1.n140 104.615
R2841 VDD1.n141 VDD1.n90 104.615
R2842 VDD1.n148 VDD1.n90 104.615
R2843 VDD1.n150 VDD1.n148 104.615
R2844 VDD1.n150 VDD1.n149 104.615
R2845 VDD1.n149 VDD1.n86 104.615
R2846 VDD1.n158 VDD1.n86 104.615
R2847 VDD1.n159 VDD1.n158 104.615
R2848 VDD1.n167 VDD1.n166 64.4019
R2849 VDD1.n82 VDD1.n81 63.0544
R2850 VDD1.n169 VDD1.n168 63.0542
R2851 VDD1.n165 VDD1.n164 63.0542
R2852 VDD1.n82 VDD1.n80 52.8682
R2853 VDD1.n165 VDD1.n163 52.8682
R2854 VDD1.n27 VDD1.t1 52.3082
R2855 VDD1.n109 VDD1.t6 52.3082
R2856 VDD1.n169 VDD1.n167 46.8349
R2857 VDD1.n28 VDD1.n26 15.6677
R2858 VDD1.n110 VDD1.n108 15.6677
R2859 VDD1.n74 VDD1.n73 13.1884
R2860 VDD1.n157 VDD1.n156 13.1884
R2861 VDD1.n77 VDD1.n2 12.8005
R2862 VDD1.n72 VDD1.n4 12.8005
R2863 VDD1.n29 VDD1.n25 12.8005
R2864 VDD1.n111 VDD1.n107 12.8005
R2865 VDD1.n155 VDD1.n87 12.8005
R2866 VDD1.n160 VDD1.n85 12.8005
R2867 VDD1.n78 VDD1.n0 12.0247
R2868 VDD1.n69 VDD1.n68 12.0247
R2869 VDD1.n33 VDD1.n32 12.0247
R2870 VDD1.n115 VDD1.n114 12.0247
R2871 VDD1.n152 VDD1.n151 12.0247
R2872 VDD1.n161 VDD1.n83 12.0247
R2873 VDD1.n65 VDD1.n6 11.249
R2874 VDD1.n36 VDD1.n23 11.249
R2875 VDD1.n118 VDD1.n105 11.249
R2876 VDD1.n147 VDD1.n89 11.249
R2877 VDD1.n64 VDD1.n9 10.4732
R2878 VDD1.n37 VDD1.n21 10.4732
R2879 VDD1.n119 VDD1.n103 10.4732
R2880 VDD1.n146 VDD1.n91 10.4732
R2881 VDD1.n61 VDD1.n60 9.69747
R2882 VDD1.n41 VDD1.n40 9.69747
R2883 VDD1.n123 VDD1.n122 9.69747
R2884 VDD1.n143 VDD1.n142 9.69747
R2885 VDD1.n80 VDD1.n79 9.45567
R2886 VDD1.n163 VDD1.n162 9.45567
R2887 VDD1.n54 VDD1.n53 9.3005
R2888 VDD1.n56 VDD1.n55 9.3005
R2889 VDD1.n11 VDD1.n10 9.3005
R2890 VDD1.n62 VDD1.n61 9.3005
R2891 VDD1.n64 VDD1.n63 9.3005
R2892 VDD1.n6 VDD1.n5 9.3005
R2893 VDD1.n70 VDD1.n69 9.3005
R2894 VDD1.n72 VDD1.n71 9.3005
R2895 VDD1.n79 VDD1.n78 9.3005
R2896 VDD1.n2 VDD1.n1 9.3005
R2897 VDD1.n15 VDD1.n14 9.3005
R2898 VDD1.n48 VDD1.n47 9.3005
R2899 VDD1.n46 VDD1.n45 9.3005
R2900 VDD1.n19 VDD1.n18 9.3005
R2901 VDD1.n40 VDD1.n39 9.3005
R2902 VDD1.n38 VDD1.n37 9.3005
R2903 VDD1.n23 VDD1.n22 9.3005
R2904 VDD1.n32 VDD1.n31 9.3005
R2905 VDD1.n30 VDD1.n29 9.3005
R2906 VDD1.n162 VDD1.n161 9.3005
R2907 VDD1.n85 VDD1.n84 9.3005
R2908 VDD1.n130 VDD1.n129 9.3005
R2909 VDD1.n128 VDD1.n127 9.3005
R2910 VDD1.n101 VDD1.n100 9.3005
R2911 VDD1.n122 VDD1.n121 9.3005
R2912 VDD1.n120 VDD1.n119 9.3005
R2913 VDD1.n105 VDD1.n104 9.3005
R2914 VDD1.n114 VDD1.n113 9.3005
R2915 VDD1.n112 VDD1.n111 9.3005
R2916 VDD1.n97 VDD1.n96 9.3005
R2917 VDD1.n136 VDD1.n135 9.3005
R2918 VDD1.n138 VDD1.n137 9.3005
R2919 VDD1.n93 VDD1.n92 9.3005
R2920 VDD1.n144 VDD1.n143 9.3005
R2921 VDD1.n146 VDD1.n145 9.3005
R2922 VDD1.n89 VDD1.n88 9.3005
R2923 VDD1.n153 VDD1.n152 9.3005
R2924 VDD1.n155 VDD1.n154 9.3005
R2925 VDD1.n57 VDD1.n11 8.92171
R2926 VDD1.n44 VDD1.n19 8.92171
R2927 VDD1.n126 VDD1.n101 8.92171
R2928 VDD1.n139 VDD1.n93 8.92171
R2929 VDD1.n56 VDD1.n13 8.14595
R2930 VDD1.n45 VDD1.n17 8.14595
R2931 VDD1.n127 VDD1.n99 8.14595
R2932 VDD1.n138 VDD1.n95 8.14595
R2933 VDD1.n53 VDD1.n52 7.3702
R2934 VDD1.n49 VDD1.n48 7.3702
R2935 VDD1.n131 VDD1.n130 7.3702
R2936 VDD1.n135 VDD1.n134 7.3702
R2937 VDD1.n52 VDD1.n15 6.59444
R2938 VDD1.n49 VDD1.n15 6.59444
R2939 VDD1.n131 VDD1.n97 6.59444
R2940 VDD1.n134 VDD1.n97 6.59444
R2941 VDD1.n53 VDD1.n13 5.81868
R2942 VDD1.n48 VDD1.n17 5.81868
R2943 VDD1.n130 VDD1.n99 5.81868
R2944 VDD1.n135 VDD1.n95 5.81868
R2945 VDD1.n57 VDD1.n56 5.04292
R2946 VDD1.n45 VDD1.n44 5.04292
R2947 VDD1.n127 VDD1.n126 5.04292
R2948 VDD1.n139 VDD1.n138 5.04292
R2949 VDD1.n30 VDD1.n26 4.38563
R2950 VDD1.n112 VDD1.n108 4.38563
R2951 VDD1.n60 VDD1.n11 4.26717
R2952 VDD1.n41 VDD1.n19 4.26717
R2953 VDD1.n123 VDD1.n101 4.26717
R2954 VDD1.n142 VDD1.n93 4.26717
R2955 VDD1.n61 VDD1.n9 3.49141
R2956 VDD1.n40 VDD1.n21 3.49141
R2957 VDD1.n122 VDD1.n103 3.49141
R2958 VDD1.n143 VDD1.n91 3.49141
R2959 VDD1.n65 VDD1.n64 2.71565
R2960 VDD1.n37 VDD1.n36 2.71565
R2961 VDD1.n119 VDD1.n118 2.71565
R2962 VDD1.n147 VDD1.n146 2.71565
R2963 VDD1.n80 VDD1.n0 1.93989
R2964 VDD1.n68 VDD1.n6 1.93989
R2965 VDD1.n33 VDD1.n23 1.93989
R2966 VDD1.n115 VDD1.n105 1.93989
R2967 VDD1.n151 VDD1.n89 1.93989
R2968 VDD1.n163 VDD1.n83 1.93989
R2969 VDD1 VDD1.n169 1.34533
R2970 VDD1.n168 VDD1.t9 1.34287
R2971 VDD1.n168 VDD1.t4 1.34287
R2972 VDD1.n81 VDD1.t5 1.34287
R2973 VDD1.n81 VDD1.t8 1.34287
R2974 VDD1.n166 VDD1.t7 1.34287
R2975 VDD1.n166 VDD1.t3 1.34287
R2976 VDD1.n164 VDD1.t2 1.34287
R2977 VDD1.n164 VDD1.t0 1.34287
R2978 VDD1.n78 VDD1.n77 1.16414
R2979 VDD1.n69 VDD1.n4 1.16414
R2980 VDD1.n32 VDD1.n25 1.16414
R2981 VDD1.n114 VDD1.n107 1.16414
R2982 VDD1.n152 VDD1.n87 1.16414
R2983 VDD1.n161 VDD1.n160 1.16414
R2984 VDD1 VDD1.n82 0.526362
R2985 VDD1.n167 VDD1.n165 0.412826
R2986 VDD1.n74 VDD1.n2 0.388379
R2987 VDD1.n73 VDD1.n72 0.388379
R2988 VDD1.n29 VDD1.n28 0.388379
R2989 VDD1.n111 VDD1.n110 0.388379
R2990 VDD1.n156 VDD1.n155 0.388379
R2991 VDD1.n157 VDD1.n85 0.388379
R2992 VDD1.n79 VDD1.n1 0.155672
R2993 VDD1.n71 VDD1.n1 0.155672
R2994 VDD1.n71 VDD1.n70 0.155672
R2995 VDD1.n70 VDD1.n5 0.155672
R2996 VDD1.n63 VDD1.n5 0.155672
R2997 VDD1.n63 VDD1.n62 0.155672
R2998 VDD1.n62 VDD1.n10 0.155672
R2999 VDD1.n55 VDD1.n10 0.155672
R3000 VDD1.n55 VDD1.n54 0.155672
R3001 VDD1.n54 VDD1.n14 0.155672
R3002 VDD1.n47 VDD1.n14 0.155672
R3003 VDD1.n47 VDD1.n46 0.155672
R3004 VDD1.n46 VDD1.n18 0.155672
R3005 VDD1.n39 VDD1.n18 0.155672
R3006 VDD1.n39 VDD1.n38 0.155672
R3007 VDD1.n38 VDD1.n22 0.155672
R3008 VDD1.n31 VDD1.n22 0.155672
R3009 VDD1.n31 VDD1.n30 0.155672
R3010 VDD1.n113 VDD1.n112 0.155672
R3011 VDD1.n113 VDD1.n104 0.155672
R3012 VDD1.n120 VDD1.n104 0.155672
R3013 VDD1.n121 VDD1.n120 0.155672
R3014 VDD1.n121 VDD1.n100 0.155672
R3015 VDD1.n128 VDD1.n100 0.155672
R3016 VDD1.n129 VDD1.n128 0.155672
R3017 VDD1.n129 VDD1.n96 0.155672
R3018 VDD1.n136 VDD1.n96 0.155672
R3019 VDD1.n137 VDD1.n136 0.155672
R3020 VDD1.n137 VDD1.n92 0.155672
R3021 VDD1.n144 VDD1.n92 0.155672
R3022 VDD1.n145 VDD1.n144 0.155672
R3023 VDD1.n145 VDD1.n88 0.155672
R3024 VDD1.n153 VDD1.n88 0.155672
R3025 VDD1.n154 VDD1.n153 0.155672
R3026 VDD1.n154 VDD1.n84 0.155672
R3027 VDD1.n162 VDD1.n84 0.155672
C0 VTAIL VP 12.2094f
C1 VDD1 VP 12.3122f
C2 VN VTAIL 12.194901f
C3 VDD2 VP 0.486806f
C4 VDD1 VN 0.151468f
C5 VDD1 VTAIL 12.059099f
C6 VDD2 VN 11.9814f
C7 VDD2 VTAIL 12.1031f
C8 VDD1 VDD2 1.67941f
C9 VN VP 7.78541f
C10 VDD2 B 6.785696f
C11 VDD1 B 6.773514f
C12 VTAIL B 8.668303f
C13 VN B 14.81092f
C14 VP B 13.174145f
C15 VDD1.n0 B 0.030116f
C16 VDD1.n1 B 0.022394f
C17 VDD1.n2 B 0.012033f
C18 VDD1.n3 B 0.028443f
C19 VDD1.n4 B 0.012741f
C20 VDD1.n5 B 0.022394f
C21 VDD1.n6 B 0.012033f
C22 VDD1.n7 B 0.028443f
C23 VDD1.n8 B 0.028443f
C24 VDD1.n9 B 0.012741f
C25 VDD1.n10 B 0.022394f
C26 VDD1.n11 B 0.012033f
C27 VDD1.n12 B 0.028443f
C28 VDD1.n13 B 0.012741f
C29 VDD1.n14 B 0.022394f
C30 VDD1.n15 B 0.012033f
C31 VDD1.n16 B 0.028443f
C32 VDD1.n17 B 0.012741f
C33 VDD1.n18 B 0.022394f
C34 VDD1.n19 B 0.012033f
C35 VDD1.n20 B 0.028443f
C36 VDD1.n21 B 0.012741f
C37 VDD1.n22 B 0.022394f
C38 VDD1.n23 B 0.012033f
C39 VDD1.n24 B 0.028443f
C40 VDD1.n25 B 0.012741f
C41 VDD1.n26 B 0.144652f
C42 VDD1.t1 B 0.046879f
C43 VDD1.n27 B 0.021332f
C44 VDD1.n28 B 0.016802f
C45 VDD1.n29 B 0.012033f
C46 VDD1.n30 B 1.4313f
C47 VDD1.n31 B 0.022394f
C48 VDD1.n32 B 0.012033f
C49 VDD1.n33 B 0.012741f
C50 VDD1.n34 B 0.028443f
C51 VDD1.n35 B 0.028443f
C52 VDD1.n36 B 0.012741f
C53 VDD1.n37 B 0.012033f
C54 VDD1.n38 B 0.022394f
C55 VDD1.n39 B 0.022394f
C56 VDD1.n40 B 0.012033f
C57 VDD1.n41 B 0.012741f
C58 VDD1.n42 B 0.028443f
C59 VDD1.n43 B 0.028443f
C60 VDD1.n44 B 0.012741f
C61 VDD1.n45 B 0.012033f
C62 VDD1.n46 B 0.022394f
C63 VDD1.n47 B 0.022394f
C64 VDD1.n48 B 0.012033f
C65 VDD1.n49 B 0.012741f
C66 VDD1.n50 B 0.028443f
C67 VDD1.n51 B 0.028443f
C68 VDD1.n52 B 0.012741f
C69 VDD1.n53 B 0.012033f
C70 VDD1.n54 B 0.022394f
C71 VDD1.n55 B 0.022394f
C72 VDD1.n56 B 0.012033f
C73 VDD1.n57 B 0.012741f
C74 VDD1.n58 B 0.028443f
C75 VDD1.n59 B 0.028443f
C76 VDD1.n60 B 0.012741f
C77 VDD1.n61 B 0.012033f
C78 VDD1.n62 B 0.022394f
C79 VDD1.n63 B 0.022394f
C80 VDD1.n64 B 0.012033f
C81 VDD1.n65 B 0.012741f
C82 VDD1.n66 B 0.028443f
C83 VDD1.n67 B 0.028443f
C84 VDD1.n68 B 0.012741f
C85 VDD1.n69 B 0.012033f
C86 VDD1.n70 B 0.022394f
C87 VDD1.n71 B 0.022394f
C88 VDD1.n72 B 0.012033f
C89 VDD1.n73 B 0.012387f
C90 VDD1.n74 B 0.012387f
C91 VDD1.n75 B 0.028443f
C92 VDD1.n76 B 0.059168f
C93 VDD1.n77 B 0.012741f
C94 VDD1.n78 B 0.012033f
C95 VDD1.n79 B 0.055127f
C96 VDD1.n80 B 0.054768f
C97 VDD1.t5 B 0.261018f
C98 VDD1.t8 B 0.261018f
C99 VDD1.n81 B 2.35956f
C100 VDD1.n82 B 0.527635f
C101 VDD1.n83 B 0.030116f
C102 VDD1.n84 B 0.022394f
C103 VDD1.n85 B 0.012033f
C104 VDD1.n86 B 0.028443f
C105 VDD1.n87 B 0.012741f
C106 VDD1.n88 B 0.022394f
C107 VDD1.n89 B 0.012033f
C108 VDD1.n90 B 0.028443f
C109 VDD1.n91 B 0.012741f
C110 VDD1.n92 B 0.022394f
C111 VDD1.n93 B 0.012033f
C112 VDD1.n94 B 0.028443f
C113 VDD1.n95 B 0.012741f
C114 VDD1.n96 B 0.022394f
C115 VDD1.n97 B 0.012033f
C116 VDD1.n98 B 0.028443f
C117 VDD1.n99 B 0.012741f
C118 VDD1.n100 B 0.022394f
C119 VDD1.n101 B 0.012033f
C120 VDD1.n102 B 0.028443f
C121 VDD1.n103 B 0.012741f
C122 VDD1.n104 B 0.022394f
C123 VDD1.n105 B 0.012033f
C124 VDD1.n106 B 0.028443f
C125 VDD1.n107 B 0.012741f
C126 VDD1.n108 B 0.144652f
C127 VDD1.t6 B 0.046879f
C128 VDD1.n109 B 0.021332f
C129 VDD1.n110 B 0.016802f
C130 VDD1.n111 B 0.012033f
C131 VDD1.n112 B 1.4313f
C132 VDD1.n113 B 0.022394f
C133 VDD1.n114 B 0.012033f
C134 VDD1.n115 B 0.012741f
C135 VDD1.n116 B 0.028443f
C136 VDD1.n117 B 0.028443f
C137 VDD1.n118 B 0.012741f
C138 VDD1.n119 B 0.012033f
C139 VDD1.n120 B 0.022394f
C140 VDD1.n121 B 0.022394f
C141 VDD1.n122 B 0.012033f
C142 VDD1.n123 B 0.012741f
C143 VDD1.n124 B 0.028443f
C144 VDD1.n125 B 0.028443f
C145 VDD1.n126 B 0.012741f
C146 VDD1.n127 B 0.012033f
C147 VDD1.n128 B 0.022394f
C148 VDD1.n129 B 0.022394f
C149 VDD1.n130 B 0.012033f
C150 VDD1.n131 B 0.012741f
C151 VDD1.n132 B 0.028443f
C152 VDD1.n133 B 0.028443f
C153 VDD1.n134 B 0.012741f
C154 VDD1.n135 B 0.012033f
C155 VDD1.n136 B 0.022394f
C156 VDD1.n137 B 0.022394f
C157 VDD1.n138 B 0.012033f
C158 VDD1.n139 B 0.012741f
C159 VDD1.n140 B 0.028443f
C160 VDD1.n141 B 0.028443f
C161 VDD1.n142 B 0.012741f
C162 VDD1.n143 B 0.012033f
C163 VDD1.n144 B 0.022394f
C164 VDD1.n145 B 0.022394f
C165 VDD1.n146 B 0.012033f
C166 VDD1.n147 B 0.012741f
C167 VDD1.n148 B 0.028443f
C168 VDD1.n149 B 0.028443f
C169 VDD1.n150 B 0.028443f
C170 VDD1.n151 B 0.012741f
C171 VDD1.n152 B 0.012033f
C172 VDD1.n153 B 0.022394f
C173 VDD1.n154 B 0.022394f
C174 VDD1.n155 B 0.012033f
C175 VDD1.n156 B 0.012387f
C176 VDD1.n157 B 0.012387f
C177 VDD1.n158 B 0.028443f
C178 VDD1.n159 B 0.059168f
C179 VDD1.n160 B 0.012741f
C180 VDD1.n161 B 0.012033f
C181 VDD1.n162 B 0.055127f
C182 VDD1.n163 B 0.054768f
C183 VDD1.t2 B 0.261018f
C184 VDD1.t0 B 0.261018f
C185 VDD1.n164 B 2.35955f
C186 VDD1.n165 B 0.52071f
C187 VDD1.t7 B 0.261018f
C188 VDD1.t3 B 0.261018f
C189 VDD1.n166 B 2.36839f
C190 VDD1.n167 B 2.49051f
C191 VDD1.t9 B 0.261018f
C192 VDD1.t4 B 0.261018f
C193 VDD1.n168 B 2.35955f
C194 VDD1.n169 B 2.74535f
C195 VP.n0 B 0.026472f
C196 VP.t6 B 1.96793f
C197 VP.n1 B 0.02141f
C198 VP.n2 B 0.026472f
C199 VP.t2 B 1.96793f
C200 VP.n3 B 0.032377f
C201 VP.n4 B 0.026472f
C202 VP.t9 B 1.96793f
C203 VP.n5 B 0.044917f
C204 VP.n6 B 0.026472f
C205 VP.t7 B 1.96793f
C206 VP.n7 B 0.052743f
C207 VP.n8 B 0.026472f
C208 VP.t3 B 1.96793f
C209 VP.n9 B 0.75801f
C210 VP.n10 B 0.026472f
C211 VP.t5 B 1.96793f
C212 VP.n11 B 0.02141f
C213 VP.n12 B 0.026472f
C214 VP.t0 B 1.96793f
C215 VP.n13 B 0.032377f
C216 VP.n14 B 0.026472f
C217 VP.t1 B 1.96793f
C218 VP.n15 B 0.044917f
C219 VP.n16 B 0.196088f
C220 VP.t4 B 1.96793f
C221 VP.t8 B 2.09365f
C222 VP.n17 B 0.754632f
C223 VP.n18 B 0.763503f
C224 VP.n19 B 0.04544f
C225 VP.n20 B 0.032377f
C226 VP.n21 B 0.026472f
C227 VP.n22 B 0.026472f
C228 VP.n23 B 0.026472f
C229 VP.n24 B 0.037158f
C230 VP.n25 B 0.6955f
C231 VP.n26 B 0.037158f
C232 VP.n27 B 0.044917f
C233 VP.n28 B 0.026472f
C234 VP.n29 B 0.026472f
C235 VP.n30 B 0.026472f
C236 VP.n31 B 0.04544f
C237 VP.n32 B 0.6955f
C238 VP.n33 B 0.028876f
C239 VP.n34 B 0.052743f
C240 VP.n35 B 0.026472f
C241 VP.n36 B 0.026472f
C242 VP.n37 B 0.026472f
C243 VP.n38 B 0.052478f
C244 VP.n39 B 0.029364f
C245 VP.n40 B 0.75801f
C246 VP.n41 B 1.48977f
C247 VP.n42 B 1.50843f
C248 VP.n43 B 0.026472f
C249 VP.n44 B 0.029364f
C250 VP.n45 B 0.052478f
C251 VP.n46 B 0.02141f
C252 VP.n47 B 0.026472f
C253 VP.n48 B 0.026472f
C254 VP.n49 B 0.026472f
C255 VP.n50 B 0.028876f
C256 VP.n51 B 0.6955f
C257 VP.n52 B 0.04544f
C258 VP.n53 B 0.032377f
C259 VP.n54 B 0.026472f
C260 VP.n55 B 0.026472f
C261 VP.n56 B 0.026472f
C262 VP.n57 B 0.037158f
C263 VP.n58 B 0.6955f
C264 VP.n59 B 0.037158f
C265 VP.n60 B 0.044917f
C266 VP.n61 B 0.026472f
C267 VP.n62 B 0.026472f
C268 VP.n63 B 0.026472f
C269 VP.n64 B 0.04544f
C270 VP.n65 B 0.6955f
C271 VP.n66 B 0.028876f
C272 VP.n67 B 0.052743f
C273 VP.n68 B 0.026472f
C274 VP.n69 B 0.026472f
C275 VP.n70 B 0.026472f
C276 VP.n71 B 0.052478f
C277 VP.n72 B 0.029364f
C278 VP.n73 B 0.75801f
C279 VP.n74 B 0.02829f
C280 VTAIL.t17 B 0.279367f
C281 VTAIL.t12 B 0.279367f
C282 VTAIL.n0 B 2.45738f
C283 VTAIL.n1 B 0.450628f
C284 VTAIL.n2 B 0.032234f
C285 VTAIL.n3 B 0.023968f
C286 VTAIL.n4 B 0.012879f
C287 VTAIL.n5 B 0.030442f
C288 VTAIL.n6 B 0.013637f
C289 VTAIL.n7 B 0.023968f
C290 VTAIL.n8 B 0.012879f
C291 VTAIL.n9 B 0.030442f
C292 VTAIL.n10 B 0.013637f
C293 VTAIL.n11 B 0.023968f
C294 VTAIL.n12 B 0.012879f
C295 VTAIL.n13 B 0.030442f
C296 VTAIL.n14 B 0.013637f
C297 VTAIL.n15 B 0.023968f
C298 VTAIL.n16 B 0.012879f
C299 VTAIL.n17 B 0.030442f
C300 VTAIL.n18 B 0.013637f
C301 VTAIL.n19 B 0.023968f
C302 VTAIL.n20 B 0.012879f
C303 VTAIL.n21 B 0.030442f
C304 VTAIL.n22 B 0.013637f
C305 VTAIL.n23 B 0.023968f
C306 VTAIL.n24 B 0.012879f
C307 VTAIL.n25 B 0.030442f
C308 VTAIL.n26 B 0.013637f
C309 VTAIL.n27 B 0.154821f
C310 VTAIL.t1 B 0.050175f
C311 VTAIL.n28 B 0.022831f
C312 VTAIL.n29 B 0.017983f
C313 VTAIL.n30 B 0.012879f
C314 VTAIL.n31 B 1.53192f
C315 VTAIL.n32 B 0.023968f
C316 VTAIL.n33 B 0.012879f
C317 VTAIL.n34 B 0.013637f
C318 VTAIL.n35 B 0.030442f
C319 VTAIL.n36 B 0.030442f
C320 VTAIL.n37 B 0.013637f
C321 VTAIL.n38 B 0.012879f
C322 VTAIL.n39 B 0.023968f
C323 VTAIL.n40 B 0.023968f
C324 VTAIL.n41 B 0.012879f
C325 VTAIL.n42 B 0.013637f
C326 VTAIL.n43 B 0.030442f
C327 VTAIL.n44 B 0.030442f
C328 VTAIL.n45 B 0.013637f
C329 VTAIL.n46 B 0.012879f
C330 VTAIL.n47 B 0.023968f
C331 VTAIL.n48 B 0.023968f
C332 VTAIL.n49 B 0.012879f
C333 VTAIL.n50 B 0.013637f
C334 VTAIL.n51 B 0.030442f
C335 VTAIL.n52 B 0.030442f
C336 VTAIL.n53 B 0.013637f
C337 VTAIL.n54 B 0.012879f
C338 VTAIL.n55 B 0.023968f
C339 VTAIL.n56 B 0.023968f
C340 VTAIL.n57 B 0.012879f
C341 VTAIL.n58 B 0.013637f
C342 VTAIL.n59 B 0.030442f
C343 VTAIL.n60 B 0.030442f
C344 VTAIL.n61 B 0.013637f
C345 VTAIL.n62 B 0.012879f
C346 VTAIL.n63 B 0.023968f
C347 VTAIL.n64 B 0.023968f
C348 VTAIL.n65 B 0.012879f
C349 VTAIL.n66 B 0.013637f
C350 VTAIL.n67 B 0.030442f
C351 VTAIL.n68 B 0.030442f
C352 VTAIL.n69 B 0.030442f
C353 VTAIL.n70 B 0.013637f
C354 VTAIL.n71 B 0.012879f
C355 VTAIL.n72 B 0.023968f
C356 VTAIL.n73 B 0.023968f
C357 VTAIL.n74 B 0.012879f
C358 VTAIL.n75 B 0.013258f
C359 VTAIL.n76 B 0.013258f
C360 VTAIL.n77 B 0.030442f
C361 VTAIL.n78 B 0.063328f
C362 VTAIL.n79 B 0.013637f
C363 VTAIL.n80 B 0.012879f
C364 VTAIL.n81 B 0.059002f
C365 VTAIL.n82 B 0.035278f
C366 VTAIL.n83 B 0.275501f
C367 VTAIL.t7 B 0.279367f
C368 VTAIL.t3 B 0.279367f
C369 VTAIL.n84 B 2.45738f
C370 VTAIL.n85 B 0.518205f
C371 VTAIL.t19 B 0.279367f
C372 VTAIL.t0 B 0.279367f
C373 VTAIL.n86 B 2.45738f
C374 VTAIL.n87 B 1.97027f
C375 VTAIL.t9 B 0.279367f
C376 VTAIL.t16 B 0.279367f
C377 VTAIL.n88 B 2.45739f
C378 VTAIL.n89 B 1.97026f
C379 VTAIL.t13 B 0.279367f
C380 VTAIL.t14 B 0.279367f
C381 VTAIL.n90 B 2.45739f
C382 VTAIL.n91 B 0.518193f
C383 VTAIL.n92 B 0.032234f
C384 VTAIL.n93 B 0.023968f
C385 VTAIL.n94 B 0.012879f
C386 VTAIL.n95 B 0.030442f
C387 VTAIL.n96 B 0.013637f
C388 VTAIL.n97 B 0.023968f
C389 VTAIL.n98 B 0.012879f
C390 VTAIL.n99 B 0.030442f
C391 VTAIL.n100 B 0.030442f
C392 VTAIL.n101 B 0.013637f
C393 VTAIL.n102 B 0.023968f
C394 VTAIL.n103 B 0.012879f
C395 VTAIL.n104 B 0.030442f
C396 VTAIL.n105 B 0.013637f
C397 VTAIL.n106 B 0.023968f
C398 VTAIL.n107 B 0.012879f
C399 VTAIL.n108 B 0.030442f
C400 VTAIL.n109 B 0.013637f
C401 VTAIL.n110 B 0.023968f
C402 VTAIL.n111 B 0.012879f
C403 VTAIL.n112 B 0.030442f
C404 VTAIL.n113 B 0.013637f
C405 VTAIL.n114 B 0.023968f
C406 VTAIL.n115 B 0.012879f
C407 VTAIL.n116 B 0.030442f
C408 VTAIL.n117 B 0.013637f
C409 VTAIL.n118 B 0.154821f
C410 VTAIL.t11 B 0.050175f
C411 VTAIL.n119 B 0.022831f
C412 VTAIL.n120 B 0.017983f
C413 VTAIL.n121 B 0.012879f
C414 VTAIL.n122 B 1.53192f
C415 VTAIL.n123 B 0.023968f
C416 VTAIL.n124 B 0.012879f
C417 VTAIL.n125 B 0.013637f
C418 VTAIL.n126 B 0.030442f
C419 VTAIL.n127 B 0.030442f
C420 VTAIL.n128 B 0.013637f
C421 VTAIL.n129 B 0.012879f
C422 VTAIL.n130 B 0.023968f
C423 VTAIL.n131 B 0.023968f
C424 VTAIL.n132 B 0.012879f
C425 VTAIL.n133 B 0.013637f
C426 VTAIL.n134 B 0.030442f
C427 VTAIL.n135 B 0.030442f
C428 VTAIL.n136 B 0.013637f
C429 VTAIL.n137 B 0.012879f
C430 VTAIL.n138 B 0.023968f
C431 VTAIL.n139 B 0.023968f
C432 VTAIL.n140 B 0.012879f
C433 VTAIL.n141 B 0.013637f
C434 VTAIL.n142 B 0.030442f
C435 VTAIL.n143 B 0.030442f
C436 VTAIL.n144 B 0.013637f
C437 VTAIL.n145 B 0.012879f
C438 VTAIL.n146 B 0.023968f
C439 VTAIL.n147 B 0.023968f
C440 VTAIL.n148 B 0.012879f
C441 VTAIL.n149 B 0.013637f
C442 VTAIL.n150 B 0.030442f
C443 VTAIL.n151 B 0.030442f
C444 VTAIL.n152 B 0.013637f
C445 VTAIL.n153 B 0.012879f
C446 VTAIL.n154 B 0.023968f
C447 VTAIL.n155 B 0.023968f
C448 VTAIL.n156 B 0.012879f
C449 VTAIL.n157 B 0.013637f
C450 VTAIL.n158 B 0.030442f
C451 VTAIL.n159 B 0.030442f
C452 VTAIL.n160 B 0.013637f
C453 VTAIL.n161 B 0.012879f
C454 VTAIL.n162 B 0.023968f
C455 VTAIL.n163 B 0.023968f
C456 VTAIL.n164 B 0.012879f
C457 VTAIL.n165 B 0.013258f
C458 VTAIL.n166 B 0.013258f
C459 VTAIL.n167 B 0.030442f
C460 VTAIL.n168 B 0.063328f
C461 VTAIL.n169 B 0.013637f
C462 VTAIL.n170 B 0.012879f
C463 VTAIL.n171 B 0.059002f
C464 VTAIL.n172 B 0.035278f
C465 VTAIL.n173 B 0.275501f
C466 VTAIL.t2 B 0.279367f
C467 VTAIL.t5 B 0.279367f
C468 VTAIL.n174 B 2.45739f
C469 VTAIL.n175 B 0.482241f
C470 VTAIL.t4 B 0.279367f
C471 VTAIL.t8 B 0.279367f
C472 VTAIL.n176 B 2.45739f
C473 VTAIL.n177 B 0.518193f
C474 VTAIL.n178 B 0.032234f
C475 VTAIL.n179 B 0.023968f
C476 VTAIL.n180 B 0.012879f
C477 VTAIL.n181 B 0.030442f
C478 VTAIL.n182 B 0.013637f
C479 VTAIL.n183 B 0.023968f
C480 VTAIL.n184 B 0.012879f
C481 VTAIL.n185 B 0.030442f
C482 VTAIL.n186 B 0.030442f
C483 VTAIL.n187 B 0.013637f
C484 VTAIL.n188 B 0.023968f
C485 VTAIL.n189 B 0.012879f
C486 VTAIL.n190 B 0.030442f
C487 VTAIL.n191 B 0.013637f
C488 VTAIL.n192 B 0.023968f
C489 VTAIL.n193 B 0.012879f
C490 VTAIL.n194 B 0.030442f
C491 VTAIL.n195 B 0.013637f
C492 VTAIL.n196 B 0.023968f
C493 VTAIL.n197 B 0.012879f
C494 VTAIL.n198 B 0.030442f
C495 VTAIL.n199 B 0.013637f
C496 VTAIL.n200 B 0.023968f
C497 VTAIL.n201 B 0.012879f
C498 VTAIL.n202 B 0.030442f
C499 VTAIL.n203 B 0.013637f
C500 VTAIL.n204 B 0.154821f
C501 VTAIL.t6 B 0.050175f
C502 VTAIL.n205 B 0.022831f
C503 VTAIL.n206 B 0.017983f
C504 VTAIL.n207 B 0.012879f
C505 VTAIL.n208 B 1.53192f
C506 VTAIL.n209 B 0.023968f
C507 VTAIL.n210 B 0.012879f
C508 VTAIL.n211 B 0.013637f
C509 VTAIL.n212 B 0.030442f
C510 VTAIL.n213 B 0.030442f
C511 VTAIL.n214 B 0.013637f
C512 VTAIL.n215 B 0.012879f
C513 VTAIL.n216 B 0.023968f
C514 VTAIL.n217 B 0.023968f
C515 VTAIL.n218 B 0.012879f
C516 VTAIL.n219 B 0.013637f
C517 VTAIL.n220 B 0.030442f
C518 VTAIL.n221 B 0.030442f
C519 VTAIL.n222 B 0.013637f
C520 VTAIL.n223 B 0.012879f
C521 VTAIL.n224 B 0.023968f
C522 VTAIL.n225 B 0.023968f
C523 VTAIL.n226 B 0.012879f
C524 VTAIL.n227 B 0.013637f
C525 VTAIL.n228 B 0.030442f
C526 VTAIL.n229 B 0.030442f
C527 VTAIL.n230 B 0.013637f
C528 VTAIL.n231 B 0.012879f
C529 VTAIL.n232 B 0.023968f
C530 VTAIL.n233 B 0.023968f
C531 VTAIL.n234 B 0.012879f
C532 VTAIL.n235 B 0.013637f
C533 VTAIL.n236 B 0.030442f
C534 VTAIL.n237 B 0.030442f
C535 VTAIL.n238 B 0.013637f
C536 VTAIL.n239 B 0.012879f
C537 VTAIL.n240 B 0.023968f
C538 VTAIL.n241 B 0.023968f
C539 VTAIL.n242 B 0.012879f
C540 VTAIL.n243 B 0.013637f
C541 VTAIL.n244 B 0.030442f
C542 VTAIL.n245 B 0.030442f
C543 VTAIL.n246 B 0.013637f
C544 VTAIL.n247 B 0.012879f
C545 VTAIL.n248 B 0.023968f
C546 VTAIL.n249 B 0.023968f
C547 VTAIL.n250 B 0.012879f
C548 VTAIL.n251 B 0.013258f
C549 VTAIL.n252 B 0.013258f
C550 VTAIL.n253 B 0.030442f
C551 VTAIL.n254 B 0.063328f
C552 VTAIL.n255 B 0.013637f
C553 VTAIL.n256 B 0.012879f
C554 VTAIL.n257 B 0.059002f
C555 VTAIL.n258 B 0.035278f
C556 VTAIL.n259 B 1.61905f
C557 VTAIL.n260 B 0.032234f
C558 VTAIL.n261 B 0.023968f
C559 VTAIL.n262 B 0.012879f
C560 VTAIL.n263 B 0.030442f
C561 VTAIL.n264 B 0.013637f
C562 VTAIL.n265 B 0.023968f
C563 VTAIL.n266 B 0.012879f
C564 VTAIL.n267 B 0.030442f
C565 VTAIL.n268 B 0.013637f
C566 VTAIL.n269 B 0.023968f
C567 VTAIL.n270 B 0.012879f
C568 VTAIL.n271 B 0.030442f
C569 VTAIL.n272 B 0.013637f
C570 VTAIL.n273 B 0.023968f
C571 VTAIL.n274 B 0.012879f
C572 VTAIL.n275 B 0.030442f
C573 VTAIL.n276 B 0.013637f
C574 VTAIL.n277 B 0.023968f
C575 VTAIL.n278 B 0.012879f
C576 VTAIL.n279 B 0.030442f
C577 VTAIL.n280 B 0.013637f
C578 VTAIL.n281 B 0.023968f
C579 VTAIL.n282 B 0.012879f
C580 VTAIL.n283 B 0.030442f
C581 VTAIL.n284 B 0.013637f
C582 VTAIL.n285 B 0.154821f
C583 VTAIL.t10 B 0.050175f
C584 VTAIL.n286 B 0.022831f
C585 VTAIL.n287 B 0.017983f
C586 VTAIL.n288 B 0.012879f
C587 VTAIL.n289 B 1.53192f
C588 VTAIL.n290 B 0.023968f
C589 VTAIL.n291 B 0.012879f
C590 VTAIL.n292 B 0.013637f
C591 VTAIL.n293 B 0.030442f
C592 VTAIL.n294 B 0.030442f
C593 VTAIL.n295 B 0.013637f
C594 VTAIL.n296 B 0.012879f
C595 VTAIL.n297 B 0.023968f
C596 VTAIL.n298 B 0.023968f
C597 VTAIL.n299 B 0.012879f
C598 VTAIL.n300 B 0.013637f
C599 VTAIL.n301 B 0.030442f
C600 VTAIL.n302 B 0.030442f
C601 VTAIL.n303 B 0.013637f
C602 VTAIL.n304 B 0.012879f
C603 VTAIL.n305 B 0.023968f
C604 VTAIL.n306 B 0.023968f
C605 VTAIL.n307 B 0.012879f
C606 VTAIL.n308 B 0.013637f
C607 VTAIL.n309 B 0.030442f
C608 VTAIL.n310 B 0.030442f
C609 VTAIL.n311 B 0.013637f
C610 VTAIL.n312 B 0.012879f
C611 VTAIL.n313 B 0.023968f
C612 VTAIL.n314 B 0.023968f
C613 VTAIL.n315 B 0.012879f
C614 VTAIL.n316 B 0.013637f
C615 VTAIL.n317 B 0.030442f
C616 VTAIL.n318 B 0.030442f
C617 VTAIL.n319 B 0.013637f
C618 VTAIL.n320 B 0.012879f
C619 VTAIL.n321 B 0.023968f
C620 VTAIL.n322 B 0.023968f
C621 VTAIL.n323 B 0.012879f
C622 VTAIL.n324 B 0.013637f
C623 VTAIL.n325 B 0.030442f
C624 VTAIL.n326 B 0.030442f
C625 VTAIL.n327 B 0.030442f
C626 VTAIL.n328 B 0.013637f
C627 VTAIL.n329 B 0.012879f
C628 VTAIL.n330 B 0.023968f
C629 VTAIL.n331 B 0.023968f
C630 VTAIL.n332 B 0.012879f
C631 VTAIL.n333 B 0.013258f
C632 VTAIL.n334 B 0.013258f
C633 VTAIL.n335 B 0.030442f
C634 VTAIL.n336 B 0.063328f
C635 VTAIL.n337 B 0.013637f
C636 VTAIL.n338 B 0.012879f
C637 VTAIL.n339 B 0.059002f
C638 VTAIL.n340 B 0.035278f
C639 VTAIL.n341 B 1.61905f
C640 VTAIL.t15 B 0.279367f
C641 VTAIL.t18 B 0.279367f
C642 VTAIL.n342 B 2.45738f
C643 VTAIL.n343 B 0.405356f
C644 VDD2.n0 B 0.029847f
C645 VDD2.n1 B 0.022194f
C646 VDD2.n2 B 0.011926f
C647 VDD2.n3 B 0.028188f
C648 VDD2.n4 B 0.012627f
C649 VDD2.n5 B 0.022194f
C650 VDD2.n6 B 0.011926f
C651 VDD2.n7 B 0.028188f
C652 VDD2.n8 B 0.012627f
C653 VDD2.n9 B 0.022194f
C654 VDD2.n10 B 0.011926f
C655 VDD2.n11 B 0.028188f
C656 VDD2.n12 B 0.012627f
C657 VDD2.n13 B 0.022194f
C658 VDD2.n14 B 0.011926f
C659 VDD2.n15 B 0.028188f
C660 VDD2.n16 B 0.012627f
C661 VDD2.n17 B 0.022194f
C662 VDD2.n18 B 0.011926f
C663 VDD2.n19 B 0.028188f
C664 VDD2.n20 B 0.012627f
C665 VDD2.n21 B 0.022194f
C666 VDD2.n22 B 0.011926f
C667 VDD2.n23 B 0.028188f
C668 VDD2.n24 B 0.012627f
C669 VDD2.n25 B 0.14336f
C670 VDD2.t7 B 0.04646f
C671 VDD2.n26 B 0.021141f
C672 VDD2.n27 B 0.016652f
C673 VDD2.n28 B 0.011926f
C674 VDD2.n29 B 1.41851f
C675 VDD2.n30 B 0.022194f
C676 VDD2.n31 B 0.011926f
C677 VDD2.n32 B 0.012627f
C678 VDD2.n33 B 0.028188f
C679 VDD2.n34 B 0.028188f
C680 VDD2.n35 B 0.012627f
C681 VDD2.n36 B 0.011926f
C682 VDD2.n37 B 0.022194f
C683 VDD2.n38 B 0.022194f
C684 VDD2.n39 B 0.011926f
C685 VDD2.n40 B 0.012627f
C686 VDD2.n41 B 0.028188f
C687 VDD2.n42 B 0.028188f
C688 VDD2.n43 B 0.012627f
C689 VDD2.n44 B 0.011926f
C690 VDD2.n45 B 0.022194f
C691 VDD2.n46 B 0.022194f
C692 VDD2.n47 B 0.011926f
C693 VDD2.n48 B 0.012627f
C694 VDD2.n49 B 0.028188f
C695 VDD2.n50 B 0.028188f
C696 VDD2.n51 B 0.012627f
C697 VDD2.n52 B 0.011926f
C698 VDD2.n53 B 0.022194f
C699 VDD2.n54 B 0.022194f
C700 VDD2.n55 B 0.011926f
C701 VDD2.n56 B 0.012627f
C702 VDD2.n57 B 0.028188f
C703 VDD2.n58 B 0.028188f
C704 VDD2.n59 B 0.012627f
C705 VDD2.n60 B 0.011926f
C706 VDD2.n61 B 0.022194f
C707 VDD2.n62 B 0.022194f
C708 VDD2.n63 B 0.011926f
C709 VDD2.n64 B 0.012627f
C710 VDD2.n65 B 0.028188f
C711 VDD2.n66 B 0.028188f
C712 VDD2.n67 B 0.028188f
C713 VDD2.n68 B 0.012627f
C714 VDD2.n69 B 0.011926f
C715 VDD2.n70 B 0.022194f
C716 VDD2.n71 B 0.022194f
C717 VDD2.n72 B 0.011926f
C718 VDD2.n73 B 0.012277f
C719 VDD2.n74 B 0.012277f
C720 VDD2.n75 B 0.028188f
C721 VDD2.n76 B 0.05864f
C722 VDD2.n77 B 0.012627f
C723 VDD2.n78 B 0.011926f
C724 VDD2.n79 B 0.054634f
C725 VDD2.n80 B 0.054279f
C726 VDD2.t0 B 0.258685f
C727 VDD2.t9 B 0.258685f
C728 VDD2.n81 B 2.33846f
C729 VDD2.n82 B 0.516057f
C730 VDD2.t5 B 0.258685f
C731 VDD2.t3 B 0.258685f
C732 VDD2.n83 B 2.34723f
C733 VDD2.n84 B 2.37367f
C734 VDD2.n85 B 0.029847f
C735 VDD2.n86 B 0.022194f
C736 VDD2.n87 B 0.011926f
C737 VDD2.n88 B 0.028188f
C738 VDD2.n89 B 0.012627f
C739 VDD2.n90 B 0.022194f
C740 VDD2.n91 B 0.011926f
C741 VDD2.n92 B 0.028188f
C742 VDD2.n93 B 0.028188f
C743 VDD2.n94 B 0.012627f
C744 VDD2.n95 B 0.022194f
C745 VDD2.n96 B 0.011926f
C746 VDD2.n97 B 0.028188f
C747 VDD2.n98 B 0.012627f
C748 VDD2.n99 B 0.022194f
C749 VDD2.n100 B 0.011926f
C750 VDD2.n101 B 0.028188f
C751 VDD2.n102 B 0.012627f
C752 VDD2.n103 B 0.022194f
C753 VDD2.n104 B 0.011926f
C754 VDD2.n105 B 0.028188f
C755 VDD2.n106 B 0.012627f
C756 VDD2.n107 B 0.022194f
C757 VDD2.n108 B 0.011926f
C758 VDD2.n109 B 0.028188f
C759 VDD2.n110 B 0.012627f
C760 VDD2.n111 B 0.14336f
C761 VDD2.t2 B 0.04646f
C762 VDD2.n112 B 0.021141f
C763 VDD2.n113 B 0.016652f
C764 VDD2.n114 B 0.011926f
C765 VDD2.n115 B 1.41851f
C766 VDD2.n116 B 0.022194f
C767 VDD2.n117 B 0.011926f
C768 VDD2.n118 B 0.012627f
C769 VDD2.n119 B 0.028188f
C770 VDD2.n120 B 0.028188f
C771 VDD2.n121 B 0.012627f
C772 VDD2.n122 B 0.011926f
C773 VDD2.n123 B 0.022194f
C774 VDD2.n124 B 0.022194f
C775 VDD2.n125 B 0.011926f
C776 VDD2.n126 B 0.012627f
C777 VDD2.n127 B 0.028188f
C778 VDD2.n128 B 0.028188f
C779 VDD2.n129 B 0.012627f
C780 VDD2.n130 B 0.011926f
C781 VDD2.n131 B 0.022194f
C782 VDD2.n132 B 0.022194f
C783 VDD2.n133 B 0.011926f
C784 VDD2.n134 B 0.012627f
C785 VDD2.n135 B 0.028188f
C786 VDD2.n136 B 0.028188f
C787 VDD2.n137 B 0.012627f
C788 VDD2.n138 B 0.011926f
C789 VDD2.n139 B 0.022194f
C790 VDD2.n140 B 0.022194f
C791 VDD2.n141 B 0.011926f
C792 VDD2.n142 B 0.012627f
C793 VDD2.n143 B 0.028188f
C794 VDD2.n144 B 0.028188f
C795 VDD2.n145 B 0.012627f
C796 VDD2.n146 B 0.011926f
C797 VDD2.n147 B 0.022194f
C798 VDD2.n148 B 0.022194f
C799 VDD2.n149 B 0.011926f
C800 VDD2.n150 B 0.012627f
C801 VDD2.n151 B 0.028188f
C802 VDD2.n152 B 0.028188f
C803 VDD2.n153 B 0.012627f
C804 VDD2.n154 B 0.011926f
C805 VDD2.n155 B 0.022194f
C806 VDD2.n156 B 0.022194f
C807 VDD2.n157 B 0.011926f
C808 VDD2.n158 B 0.012277f
C809 VDD2.n159 B 0.012277f
C810 VDD2.n160 B 0.028188f
C811 VDD2.n161 B 0.05864f
C812 VDD2.n162 B 0.012627f
C813 VDD2.n163 B 0.011926f
C814 VDD2.n164 B 0.054634f
C815 VDD2.n165 B 0.047966f
C816 VDD2.n166 B 2.49353f
C817 VDD2.t6 B 0.258685f
C818 VDD2.t1 B 0.258685f
C819 VDD2.n167 B 2.33847f
C820 VDD2.n168 B 0.350811f
C821 VDD2.t8 B 0.258685f
C822 VDD2.t4 B 0.258685f
C823 VDD2.n169 B 2.3472f
C824 VN.n0 B 0.026196f
C825 VN.t8 B 1.9474f
C826 VN.n1 B 0.021186f
C827 VN.n2 B 0.026196f
C828 VN.t0 B 1.9474f
C829 VN.n3 B 0.032039f
C830 VN.n4 B 0.026196f
C831 VN.t3 B 1.9474f
C832 VN.n5 B 0.044448f
C833 VN.n6 B 0.194043f
C834 VN.t6 B 1.9474f
C835 VN.t1 B 2.07181f
C836 VN.n7 B 0.746763f
C837 VN.n8 B 0.755541f
C838 VN.n9 B 0.044966f
C839 VN.n10 B 0.032039f
C840 VN.n11 B 0.026196f
C841 VN.n12 B 0.026196f
C842 VN.n13 B 0.026196f
C843 VN.n14 B 0.036771f
C844 VN.n15 B 0.688247f
C845 VN.n16 B 0.036771f
C846 VN.n17 B 0.044448f
C847 VN.n18 B 0.026196f
C848 VN.n19 B 0.026196f
C849 VN.n20 B 0.026196f
C850 VN.n21 B 0.044966f
C851 VN.n22 B 0.688247f
C852 VN.n23 B 0.028575f
C853 VN.n24 B 0.052193f
C854 VN.n25 B 0.026196f
C855 VN.n26 B 0.026196f
C856 VN.n27 B 0.026196f
C857 VN.n28 B 0.05193f
C858 VN.n29 B 0.029057f
C859 VN.n30 B 0.750105f
C860 VN.n31 B 0.027995f
C861 VN.n32 B 0.026196f
C862 VN.t9 B 1.9474f
C863 VN.n33 B 0.021186f
C864 VN.n34 B 0.026196f
C865 VN.t2 B 1.9474f
C866 VN.n35 B 0.032039f
C867 VN.n36 B 0.026196f
C868 VN.t5 B 1.9474f
C869 VN.n37 B 0.044448f
C870 VN.n38 B 0.194043f
C871 VN.t4 B 1.9474f
C872 VN.t7 B 2.07181f
C873 VN.n39 B 0.746763f
C874 VN.n40 B 0.755541f
C875 VN.n41 B 0.044966f
C876 VN.n42 B 0.032039f
C877 VN.n43 B 0.026196f
C878 VN.n44 B 0.026196f
C879 VN.n45 B 0.026196f
C880 VN.n46 B 0.036771f
C881 VN.n47 B 0.688247f
C882 VN.n48 B 0.036771f
C883 VN.n49 B 0.044448f
C884 VN.n50 B 0.026196f
C885 VN.n51 B 0.026196f
C886 VN.n52 B 0.026196f
C887 VN.n53 B 0.044966f
C888 VN.n54 B 0.688247f
C889 VN.n55 B 0.028575f
C890 VN.n56 B 0.052193f
C891 VN.n57 B 0.026196f
C892 VN.n58 B 0.026196f
C893 VN.n59 B 0.026196f
C894 VN.n60 B 0.05193f
C895 VN.n61 B 0.029057f
C896 VN.n62 B 0.750105f
C897 VN.n63 B 1.49125f
.ends

