* NGSPICE file created from diff_pair_sample_1614.ext - technology: sky130A

.subckt diff_pair_sample_1614 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=5.7993 ps=30.52 w=14.87 l=0.59
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=0 ps=0 w=14.87 l=0.59
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=0 ps=0 w=14.87 l=0.59
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=0 ps=0 w=14.87 l=0.59
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=5.7993 ps=30.52 w=14.87 l=0.59
X5 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=5.7993 ps=30.52 w=14.87 l=0.59
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=0 ps=0 w=14.87 l=0.59
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7993 pd=30.52 as=5.7993 ps=30.52 w=14.87 l=0.59
R0 VN VN.t0 877.587
R1 VN VN.t1 835.744
R2 VTAIL.n322 VTAIL.n246 289.615
R3 VTAIL.n76 VTAIL.n0 289.615
R4 VTAIL.n240 VTAIL.n164 289.615
R5 VTAIL.n158 VTAIL.n82 289.615
R6 VTAIL.n273 VTAIL.n272 185
R7 VTAIL.n270 VTAIL.n269 185
R8 VTAIL.n279 VTAIL.n278 185
R9 VTAIL.n281 VTAIL.n280 185
R10 VTAIL.n266 VTAIL.n265 185
R11 VTAIL.n287 VTAIL.n286 185
R12 VTAIL.n289 VTAIL.n288 185
R13 VTAIL.n262 VTAIL.n261 185
R14 VTAIL.n295 VTAIL.n294 185
R15 VTAIL.n297 VTAIL.n296 185
R16 VTAIL.n258 VTAIL.n257 185
R17 VTAIL.n303 VTAIL.n302 185
R18 VTAIL.n305 VTAIL.n304 185
R19 VTAIL.n254 VTAIL.n253 185
R20 VTAIL.n311 VTAIL.n310 185
R21 VTAIL.n314 VTAIL.n313 185
R22 VTAIL.n312 VTAIL.n250 185
R23 VTAIL.n319 VTAIL.n249 185
R24 VTAIL.n321 VTAIL.n320 185
R25 VTAIL.n323 VTAIL.n322 185
R26 VTAIL.n27 VTAIL.n26 185
R27 VTAIL.n24 VTAIL.n23 185
R28 VTAIL.n33 VTAIL.n32 185
R29 VTAIL.n35 VTAIL.n34 185
R30 VTAIL.n20 VTAIL.n19 185
R31 VTAIL.n41 VTAIL.n40 185
R32 VTAIL.n43 VTAIL.n42 185
R33 VTAIL.n16 VTAIL.n15 185
R34 VTAIL.n49 VTAIL.n48 185
R35 VTAIL.n51 VTAIL.n50 185
R36 VTAIL.n12 VTAIL.n11 185
R37 VTAIL.n57 VTAIL.n56 185
R38 VTAIL.n59 VTAIL.n58 185
R39 VTAIL.n8 VTAIL.n7 185
R40 VTAIL.n65 VTAIL.n64 185
R41 VTAIL.n68 VTAIL.n67 185
R42 VTAIL.n66 VTAIL.n4 185
R43 VTAIL.n73 VTAIL.n3 185
R44 VTAIL.n75 VTAIL.n74 185
R45 VTAIL.n77 VTAIL.n76 185
R46 VTAIL.n241 VTAIL.n240 185
R47 VTAIL.n239 VTAIL.n238 185
R48 VTAIL.n237 VTAIL.n167 185
R49 VTAIL.n171 VTAIL.n168 185
R50 VTAIL.n232 VTAIL.n231 185
R51 VTAIL.n230 VTAIL.n229 185
R52 VTAIL.n173 VTAIL.n172 185
R53 VTAIL.n224 VTAIL.n223 185
R54 VTAIL.n222 VTAIL.n221 185
R55 VTAIL.n177 VTAIL.n176 185
R56 VTAIL.n216 VTAIL.n215 185
R57 VTAIL.n214 VTAIL.n213 185
R58 VTAIL.n181 VTAIL.n180 185
R59 VTAIL.n208 VTAIL.n207 185
R60 VTAIL.n206 VTAIL.n205 185
R61 VTAIL.n185 VTAIL.n184 185
R62 VTAIL.n200 VTAIL.n199 185
R63 VTAIL.n198 VTAIL.n197 185
R64 VTAIL.n189 VTAIL.n188 185
R65 VTAIL.n192 VTAIL.n191 185
R66 VTAIL.n159 VTAIL.n158 185
R67 VTAIL.n157 VTAIL.n156 185
R68 VTAIL.n155 VTAIL.n85 185
R69 VTAIL.n89 VTAIL.n86 185
R70 VTAIL.n150 VTAIL.n149 185
R71 VTAIL.n148 VTAIL.n147 185
R72 VTAIL.n91 VTAIL.n90 185
R73 VTAIL.n142 VTAIL.n141 185
R74 VTAIL.n140 VTAIL.n139 185
R75 VTAIL.n95 VTAIL.n94 185
R76 VTAIL.n134 VTAIL.n133 185
R77 VTAIL.n132 VTAIL.n131 185
R78 VTAIL.n99 VTAIL.n98 185
R79 VTAIL.n126 VTAIL.n125 185
R80 VTAIL.n124 VTAIL.n123 185
R81 VTAIL.n103 VTAIL.n102 185
R82 VTAIL.n118 VTAIL.n117 185
R83 VTAIL.n116 VTAIL.n115 185
R84 VTAIL.n107 VTAIL.n106 185
R85 VTAIL.n110 VTAIL.n109 185
R86 VTAIL.t0 VTAIL.n190 147.659
R87 VTAIL.t2 VTAIL.n108 147.659
R88 VTAIL.t3 VTAIL.n271 147.659
R89 VTAIL.t1 VTAIL.n25 147.659
R90 VTAIL.n272 VTAIL.n269 104.615
R91 VTAIL.n279 VTAIL.n269 104.615
R92 VTAIL.n280 VTAIL.n279 104.615
R93 VTAIL.n280 VTAIL.n265 104.615
R94 VTAIL.n287 VTAIL.n265 104.615
R95 VTAIL.n288 VTAIL.n287 104.615
R96 VTAIL.n288 VTAIL.n261 104.615
R97 VTAIL.n295 VTAIL.n261 104.615
R98 VTAIL.n296 VTAIL.n295 104.615
R99 VTAIL.n296 VTAIL.n257 104.615
R100 VTAIL.n303 VTAIL.n257 104.615
R101 VTAIL.n304 VTAIL.n303 104.615
R102 VTAIL.n304 VTAIL.n253 104.615
R103 VTAIL.n311 VTAIL.n253 104.615
R104 VTAIL.n313 VTAIL.n311 104.615
R105 VTAIL.n313 VTAIL.n312 104.615
R106 VTAIL.n312 VTAIL.n249 104.615
R107 VTAIL.n321 VTAIL.n249 104.615
R108 VTAIL.n322 VTAIL.n321 104.615
R109 VTAIL.n26 VTAIL.n23 104.615
R110 VTAIL.n33 VTAIL.n23 104.615
R111 VTAIL.n34 VTAIL.n33 104.615
R112 VTAIL.n34 VTAIL.n19 104.615
R113 VTAIL.n41 VTAIL.n19 104.615
R114 VTAIL.n42 VTAIL.n41 104.615
R115 VTAIL.n42 VTAIL.n15 104.615
R116 VTAIL.n49 VTAIL.n15 104.615
R117 VTAIL.n50 VTAIL.n49 104.615
R118 VTAIL.n50 VTAIL.n11 104.615
R119 VTAIL.n57 VTAIL.n11 104.615
R120 VTAIL.n58 VTAIL.n57 104.615
R121 VTAIL.n58 VTAIL.n7 104.615
R122 VTAIL.n65 VTAIL.n7 104.615
R123 VTAIL.n67 VTAIL.n65 104.615
R124 VTAIL.n67 VTAIL.n66 104.615
R125 VTAIL.n66 VTAIL.n3 104.615
R126 VTAIL.n75 VTAIL.n3 104.615
R127 VTAIL.n76 VTAIL.n75 104.615
R128 VTAIL.n240 VTAIL.n239 104.615
R129 VTAIL.n239 VTAIL.n167 104.615
R130 VTAIL.n171 VTAIL.n167 104.615
R131 VTAIL.n231 VTAIL.n171 104.615
R132 VTAIL.n231 VTAIL.n230 104.615
R133 VTAIL.n230 VTAIL.n172 104.615
R134 VTAIL.n223 VTAIL.n172 104.615
R135 VTAIL.n223 VTAIL.n222 104.615
R136 VTAIL.n222 VTAIL.n176 104.615
R137 VTAIL.n215 VTAIL.n176 104.615
R138 VTAIL.n215 VTAIL.n214 104.615
R139 VTAIL.n214 VTAIL.n180 104.615
R140 VTAIL.n207 VTAIL.n180 104.615
R141 VTAIL.n207 VTAIL.n206 104.615
R142 VTAIL.n206 VTAIL.n184 104.615
R143 VTAIL.n199 VTAIL.n184 104.615
R144 VTAIL.n199 VTAIL.n198 104.615
R145 VTAIL.n198 VTAIL.n188 104.615
R146 VTAIL.n191 VTAIL.n188 104.615
R147 VTAIL.n158 VTAIL.n157 104.615
R148 VTAIL.n157 VTAIL.n85 104.615
R149 VTAIL.n89 VTAIL.n85 104.615
R150 VTAIL.n149 VTAIL.n89 104.615
R151 VTAIL.n149 VTAIL.n148 104.615
R152 VTAIL.n148 VTAIL.n90 104.615
R153 VTAIL.n141 VTAIL.n90 104.615
R154 VTAIL.n141 VTAIL.n140 104.615
R155 VTAIL.n140 VTAIL.n94 104.615
R156 VTAIL.n133 VTAIL.n94 104.615
R157 VTAIL.n133 VTAIL.n132 104.615
R158 VTAIL.n132 VTAIL.n98 104.615
R159 VTAIL.n125 VTAIL.n98 104.615
R160 VTAIL.n125 VTAIL.n124 104.615
R161 VTAIL.n124 VTAIL.n102 104.615
R162 VTAIL.n117 VTAIL.n102 104.615
R163 VTAIL.n117 VTAIL.n116 104.615
R164 VTAIL.n116 VTAIL.n106 104.615
R165 VTAIL.n109 VTAIL.n106 104.615
R166 VTAIL.n272 VTAIL.t3 52.3082
R167 VTAIL.n26 VTAIL.t1 52.3082
R168 VTAIL.n191 VTAIL.t0 52.3082
R169 VTAIL.n109 VTAIL.t2 52.3082
R170 VTAIL.n327 VTAIL.n326 36.646
R171 VTAIL.n81 VTAIL.n80 36.646
R172 VTAIL.n245 VTAIL.n244 36.646
R173 VTAIL.n163 VTAIL.n162 36.646
R174 VTAIL.n163 VTAIL.n81 26.7893
R175 VTAIL.n327 VTAIL.n245 25.9962
R176 VTAIL.n273 VTAIL.n271 15.6677
R177 VTAIL.n27 VTAIL.n25 15.6677
R178 VTAIL.n192 VTAIL.n190 15.6677
R179 VTAIL.n110 VTAIL.n108 15.6677
R180 VTAIL.n320 VTAIL.n319 13.1884
R181 VTAIL.n74 VTAIL.n73 13.1884
R182 VTAIL.n238 VTAIL.n237 13.1884
R183 VTAIL.n156 VTAIL.n155 13.1884
R184 VTAIL.n274 VTAIL.n270 12.8005
R185 VTAIL.n318 VTAIL.n250 12.8005
R186 VTAIL.n323 VTAIL.n248 12.8005
R187 VTAIL.n28 VTAIL.n24 12.8005
R188 VTAIL.n72 VTAIL.n4 12.8005
R189 VTAIL.n77 VTAIL.n2 12.8005
R190 VTAIL.n241 VTAIL.n166 12.8005
R191 VTAIL.n236 VTAIL.n168 12.8005
R192 VTAIL.n193 VTAIL.n189 12.8005
R193 VTAIL.n159 VTAIL.n84 12.8005
R194 VTAIL.n154 VTAIL.n86 12.8005
R195 VTAIL.n111 VTAIL.n107 12.8005
R196 VTAIL.n278 VTAIL.n277 12.0247
R197 VTAIL.n315 VTAIL.n314 12.0247
R198 VTAIL.n324 VTAIL.n246 12.0247
R199 VTAIL.n32 VTAIL.n31 12.0247
R200 VTAIL.n69 VTAIL.n68 12.0247
R201 VTAIL.n78 VTAIL.n0 12.0247
R202 VTAIL.n242 VTAIL.n164 12.0247
R203 VTAIL.n233 VTAIL.n232 12.0247
R204 VTAIL.n197 VTAIL.n196 12.0247
R205 VTAIL.n160 VTAIL.n82 12.0247
R206 VTAIL.n151 VTAIL.n150 12.0247
R207 VTAIL.n115 VTAIL.n114 12.0247
R208 VTAIL.n281 VTAIL.n268 11.249
R209 VTAIL.n310 VTAIL.n252 11.249
R210 VTAIL.n35 VTAIL.n22 11.249
R211 VTAIL.n64 VTAIL.n6 11.249
R212 VTAIL.n229 VTAIL.n170 11.249
R213 VTAIL.n200 VTAIL.n187 11.249
R214 VTAIL.n147 VTAIL.n88 11.249
R215 VTAIL.n118 VTAIL.n105 11.249
R216 VTAIL.n282 VTAIL.n266 10.4732
R217 VTAIL.n309 VTAIL.n254 10.4732
R218 VTAIL.n36 VTAIL.n20 10.4732
R219 VTAIL.n63 VTAIL.n8 10.4732
R220 VTAIL.n228 VTAIL.n173 10.4732
R221 VTAIL.n201 VTAIL.n185 10.4732
R222 VTAIL.n146 VTAIL.n91 10.4732
R223 VTAIL.n119 VTAIL.n103 10.4732
R224 VTAIL.n286 VTAIL.n285 9.69747
R225 VTAIL.n306 VTAIL.n305 9.69747
R226 VTAIL.n40 VTAIL.n39 9.69747
R227 VTAIL.n60 VTAIL.n59 9.69747
R228 VTAIL.n225 VTAIL.n224 9.69747
R229 VTAIL.n205 VTAIL.n204 9.69747
R230 VTAIL.n143 VTAIL.n142 9.69747
R231 VTAIL.n123 VTAIL.n122 9.69747
R232 VTAIL.n326 VTAIL.n325 9.45567
R233 VTAIL.n80 VTAIL.n79 9.45567
R234 VTAIL.n244 VTAIL.n243 9.45567
R235 VTAIL.n162 VTAIL.n161 9.45567
R236 VTAIL.n325 VTAIL.n324 9.3005
R237 VTAIL.n248 VTAIL.n247 9.3005
R238 VTAIL.n293 VTAIL.n292 9.3005
R239 VTAIL.n291 VTAIL.n290 9.3005
R240 VTAIL.n264 VTAIL.n263 9.3005
R241 VTAIL.n285 VTAIL.n284 9.3005
R242 VTAIL.n283 VTAIL.n282 9.3005
R243 VTAIL.n268 VTAIL.n267 9.3005
R244 VTAIL.n277 VTAIL.n276 9.3005
R245 VTAIL.n275 VTAIL.n274 9.3005
R246 VTAIL.n260 VTAIL.n259 9.3005
R247 VTAIL.n299 VTAIL.n298 9.3005
R248 VTAIL.n301 VTAIL.n300 9.3005
R249 VTAIL.n256 VTAIL.n255 9.3005
R250 VTAIL.n307 VTAIL.n306 9.3005
R251 VTAIL.n309 VTAIL.n308 9.3005
R252 VTAIL.n252 VTAIL.n251 9.3005
R253 VTAIL.n316 VTAIL.n315 9.3005
R254 VTAIL.n318 VTAIL.n317 9.3005
R255 VTAIL.n79 VTAIL.n78 9.3005
R256 VTAIL.n2 VTAIL.n1 9.3005
R257 VTAIL.n47 VTAIL.n46 9.3005
R258 VTAIL.n45 VTAIL.n44 9.3005
R259 VTAIL.n18 VTAIL.n17 9.3005
R260 VTAIL.n39 VTAIL.n38 9.3005
R261 VTAIL.n37 VTAIL.n36 9.3005
R262 VTAIL.n22 VTAIL.n21 9.3005
R263 VTAIL.n31 VTAIL.n30 9.3005
R264 VTAIL.n29 VTAIL.n28 9.3005
R265 VTAIL.n14 VTAIL.n13 9.3005
R266 VTAIL.n53 VTAIL.n52 9.3005
R267 VTAIL.n55 VTAIL.n54 9.3005
R268 VTAIL.n10 VTAIL.n9 9.3005
R269 VTAIL.n61 VTAIL.n60 9.3005
R270 VTAIL.n63 VTAIL.n62 9.3005
R271 VTAIL.n6 VTAIL.n5 9.3005
R272 VTAIL.n70 VTAIL.n69 9.3005
R273 VTAIL.n72 VTAIL.n71 9.3005
R274 VTAIL.n218 VTAIL.n217 9.3005
R275 VTAIL.n220 VTAIL.n219 9.3005
R276 VTAIL.n175 VTAIL.n174 9.3005
R277 VTAIL.n226 VTAIL.n225 9.3005
R278 VTAIL.n228 VTAIL.n227 9.3005
R279 VTAIL.n170 VTAIL.n169 9.3005
R280 VTAIL.n234 VTAIL.n233 9.3005
R281 VTAIL.n236 VTAIL.n235 9.3005
R282 VTAIL.n243 VTAIL.n242 9.3005
R283 VTAIL.n166 VTAIL.n165 9.3005
R284 VTAIL.n179 VTAIL.n178 9.3005
R285 VTAIL.n212 VTAIL.n211 9.3005
R286 VTAIL.n210 VTAIL.n209 9.3005
R287 VTAIL.n183 VTAIL.n182 9.3005
R288 VTAIL.n204 VTAIL.n203 9.3005
R289 VTAIL.n202 VTAIL.n201 9.3005
R290 VTAIL.n187 VTAIL.n186 9.3005
R291 VTAIL.n196 VTAIL.n195 9.3005
R292 VTAIL.n194 VTAIL.n193 9.3005
R293 VTAIL.n136 VTAIL.n135 9.3005
R294 VTAIL.n138 VTAIL.n137 9.3005
R295 VTAIL.n93 VTAIL.n92 9.3005
R296 VTAIL.n144 VTAIL.n143 9.3005
R297 VTAIL.n146 VTAIL.n145 9.3005
R298 VTAIL.n88 VTAIL.n87 9.3005
R299 VTAIL.n152 VTAIL.n151 9.3005
R300 VTAIL.n154 VTAIL.n153 9.3005
R301 VTAIL.n161 VTAIL.n160 9.3005
R302 VTAIL.n84 VTAIL.n83 9.3005
R303 VTAIL.n97 VTAIL.n96 9.3005
R304 VTAIL.n130 VTAIL.n129 9.3005
R305 VTAIL.n128 VTAIL.n127 9.3005
R306 VTAIL.n101 VTAIL.n100 9.3005
R307 VTAIL.n122 VTAIL.n121 9.3005
R308 VTAIL.n120 VTAIL.n119 9.3005
R309 VTAIL.n105 VTAIL.n104 9.3005
R310 VTAIL.n114 VTAIL.n113 9.3005
R311 VTAIL.n112 VTAIL.n111 9.3005
R312 VTAIL.n289 VTAIL.n264 8.92171
R313 VTAIL.n302 VTAIL.n256 8.92171
R314 VTAIL.n43 VTAIL.n18 8.92171
R315 VTAIL.n56 VTAIL.n10 8.92171
R316 VTAIL.n221 VTAIL.n175 8.92171
R317 VTAIL.n208 VTAIL.n183 8.92171
R318 VTAIL.n139 VTAIL.n93 8.92171
R319 VTAIL.n126 VTAIL.n101 8.92171
R320 VTAIL.n290 VTAIL.n262 8.14595
R321 VTAIL.n301 VTAIL.n258 8.14595
R322 VTAIL.n44 VTAIL.n16 8.14595
R323 VTAIL.n55 VTAIL.n12 8.14595
R324 VTAIL.n220 VTAIL.n177 8.14595
R325 VTAIL.n209 VTAIL.n181 8.14595
R326 VTAIL.n138 VTAIL.n95 8.14595
R327 VTAIL.n127 VTAIL.n99 8.14595
R328 VTAIL.n294 VTAIL.n293 7.3702
R329 VTAIL.n298 VTAIL.n297 7.3702
R330 VTAIL.n48 VTAIL.n47 7.3702
R331 VTAIL.n52 VTAIL.n51 7.3702
R332 VTAIL.n217 VTAIL.n216 7.3702
R333 VTAIL.n213 VTAIL.n212 7.3702
R334 VTAIL.n135 VTAIL.n134 7.3702
R335 VTAIL.n131 VTAIL.n130 7.3702
R336 VTAIL.n294 VTAIL.n260 6.59444
R337 VTAIL.n297 VTAIL.n260 6.59444
R338 VTAIL.n48 VTAIL.n14 6.59444
R339 VTAIL.n51 VTAIL.n14 6.59444
R340 VTAIL.n216 VTAIL.n179 6.59444
R341 VTAIL.n213 VTAIL.n179 6.59444
R342 VTAIL.n134 VTAIL.n97 6.59444
R343 VTAIL.n131 VTAIL.n97 6.59444
R344 VTAIL.n293 VTAIL.n262 5.81868
R345 VTAIL.n298 VTAIL.n258 5.81868
R346 VTAIL.n47 VTAIL.n16 5.81868
R347 VTAIL.n52 VTAIL.n12 5.81868
R348 VTAIL.n217 VTAIL.n177 5.81868
R349 VTAIL.n212 VTAIL.n181 5.81868
R350 VTAIL.n135 VTAIL.n95 5.81868
R351 VTAIL.n130 VTAIL.n99 5.81868
R352 VTAIL.n290 VTAIL.n289 5.04292
R353 VTAIL.n302 VTAIL.n301 5.04292
R354 VTAIL.n44 VTAIL.n43 5.04292
R355 VTAIL.n56 VTAIL.n55 5.04292
R356 VTAIL.n221 VTAIL.n220 5.04292
R357 VTAIL.n209 VTAIL.n208 5.04292
R358 VTAIL.n139 VTAIL.n138 5.04292
R359 VTAIL.n127 VTAIL.n126 5.04292
R360 VTAIL.n194 VTAIL.n190 4.38563
R361 VTAIL.n112 VTAIL.n108 4.38563
R362 VTAIL.n275 VTAIL.n271 4.38563
R363 VTAIL.n29 VTAIL.n25 4.38563
R364 VTAIL.n286 VTAIL.n264 4.26717
R365 VTAIL.n305 VTAIL.n256 4.26717
R366 VTAIL.n40 VTAIL.n18 4.26717
R367 VTAIL.n59 VTAIL.n10 4.26717
R368 VTAIL.n224 VTAIL.n175 4.26717
R369 VTAIL.n205 VTAIL.n183 4.26717
R370 VTAIL.n142 VTAIL.n93 4.26717
R371 VTAIL.n123 VTAIL.n101 4.26717
R372 VTAIL.n285 VTAIL.n266 3.49141
R373 VTAIL.n306 VTAIL.n254 3.49141
R374 VTAIL.n39 VTAIL.n20 3.49141
R375 VTAIL.n60 VTAIL.n8 3.49141
R376 VTAIL.n225 VTAIL.n173 3.49141
R377 VTAIL.n204 VTAIL.n185 3.49141
R378 VTAIL.n143 VTAIL.n91 3.49141
R379 VTAIL.n122 VTAIL.n103 3.49141
R380 VTAIL.n282 VTAIL.n281 2.71565
R381 VTAIL.n310 VTAIL.n309 2.71565
R382 VTAIL.n36 VTAIL.n35 2.71565
R383 VTAIL.n64 VTAIL.n63 2.71565
R384 VTAIL.n229 VTAIL.n228 2.71565
R385 VTAIL.n201 VTAIL.n200 2.71565
R386 VTAIL.n147 VTAIL.n146 2.71565
R387 VTAIL.n119 VTAIL.n118 2.71565
R388 VTAIL.n278 VTAIL.n268 1.93989
R389 VTAIL.n314 VTAIL.n252 1.93989
R390 VTAIL.n326 VTAIL.n246 1.93989
R391 VTAIL.n32 VTAIL.n22 1.93989
R392 VTAIL.n68 VTAIL.n6 1.93989
R393 VTAIL.n80 VTAIL.n0 1.93989
R394 VTAIL.n244 VTAIL.n164 1.93989
R395 VTAIL.n232 VTAIL.n170 1.93989
R396 VTAIL.n197 VTAIL.n187 1.93989
R397 VTAIL.n162 VTAIL.n82 1.93989
R398 VTAIL.n150 VTAIL.n88 1.93989
R399 VTAIL.n115 VTAIL.n105 1.93989
R400 VTAIL.n277 VTAIL.n270 1.16414
R401 VTAIL.n315 VTAIL.n250 1.16414
R402 VTAIL.n324 VTAIL.n323 1.16414
R403 VTAIL.n31 VTAIL.n24 1.16414
R404 VTAIL.n69 VTAIL.n4 1.16414
R405 VTAIL.n78 VTAIL.n77 1.16414
R406 VTAIL.n242 VTAIL.n241 1.16414
R407 VTAIL.n233 VTAIL.n168 1.16414
R408 VTAIL.n196 VTAIL.n189 1.16414
R409 VTAIL.n160 VTAIL.n159 1.16414
R410 VTAIL.n151 VTAIL.n86 1.16414
R411 VTAIL.n114 VTAIL.n107 1.16414
R412 VTAIL.n245 VTAIL.n163 0.866879
R413 VTAIL VTAIL.n81 0.726793
R414 VTAIL.n274 VTAIL.n273 0.388379
R415 VTAIL.n319 VTAIL.n318 0.388379
R416 VTAIL.n320 VTAIL.n248 0.388379
R417 VTAIL.n28 VTAIL.n27 0.388379
R418 VTAIL.n73 VTAIL.n72 0.388379
R419 VTAIL.n74 VTAIL.n2 0.388379
R420 VTAIL.n238 VTAIL.n166 0.388379
R421 VTAIL.n237 VTAIL.n236 0.388379
R422 VTAIL.n193 VTAIL.n192 0.388379
R423 VTAIL.n156 VTAIL.n84 0.388379
R424 VTAIL.n155 VTAIL.n154 0.388379
R425 VTAIL.n111 VTAIL.n110 0.388379
R426 VTAIL.n276 VTAIL.n275 0.155672
R427 VTAIL.n276 VTAIL.n267 0.155672
R428 VTAIL.n283 VTAIL.n267 0.155672
R429 VTAIL.n284 VTAIL.n283 0.155672
R430 VTAIL.n284 VTAIL.n263 0.155672
R431 VTAIL.n291 VTAIL.n263 0.155672
R432 VTAIL.n292 VTAIL.n291 0.155672
R433 VTAIL.n292 VTAIL.n259 0.155672
R434 VTAIL.n299 VTAIL.n259 0.155672
R435 VTAIL.n300 VTAIL.n299 0.155672
R436 VTAIL.n300 VTAIL.n255 0.155672
R437 VTAIL.n307 VTAIL.n255 0.155672
R438 VTAIL.n308 VTAIL.n307 0.155672
R439 VTAIL.n308 VTAIL.n251 0.155672
R440 VTAIL.n316 VTAIL.n251 0.155672
R441 VTAIL.n317 VTAIL.n316 0.155672
R442 VTAIL.n317 VTAIL.n247 0.155672
R443 VTAIL.n325 VTAIL.n247 0.155672
R444 VTAIL.n30 VTAIL.n29 0.155672
R445 VTAIL.n30 VTAIL.n21 0.155672
R446 VTAIL.n37 VTAIL.n21 0.155672
R447 VTAIL.n38 VTAIL.n37 0.155672
R448 VTAIL.n38 VTAIL.n17 0.155672
R449 VTAIL.n45 VTAIL.n17 0.155672
R450 VTAIL.n46 VTAIL.n45 0.155672
R451 VTAIL.n46 VTAIL.n13 0.155672
R452 VTAIL.n53 VTAIL.n13 0.155672
R453 VTAIL.n54 VTAIL.n53 0.155672
R454 VTAIL.n54 VTAIL.n9 0.155672
R455 VTAIL.n61 VTAIL.n9 0.155672
R456 VTAIL.n62 VTAIL.n61 0.155672
R457 VTAIL.n62 VTAIL.n5 0.155672
R458 VTAIL.n70 VTAIL.n5 0.155672
R459 VTAIL.n71 VTAIL.n70 0.155672
R460 VTAIL.n71 VTAIL.n1 0.155672
R461 VTAIL.n79 VTAIL.n1 0.155672
R462 VTAIL.n243 VTAIL.n165 0.155672
R463 VTAIL.n235 VTAIL.n165 0.155672
R464 VTAIL.n235 VTAIL.n234 0.155672
R465 VTAIL.n234 VTAIL.n169 0.155672
R466 VTAIL.n227 VTAIL.n169 0.155672
R467 VTAIL.n227 VTAIL.n226 0.155672
R468 VTAIL.n226 VTAIL.n174 0.155672
R469 VTAIL.n219 VTAIL.n174 0.155672
R470 VTAIL.n219 VTAIL.n218 0.155672
R471 VTAIL.n218 VTAIL.n178 0.155672
R472 VTAIL.n211 VTAIL.n178 0.155672
R473 VTAIL.n211 VTAIL.n210 0.155672
R474 VTAIL.n210 VTAIL.n182 0.155672
R475 VTAIL.n203 VTAIL.n182 0.155672
R476 VTAIL.n203 VTAIL.n202 0.155672
R477 VTAIL.n202 VTAIL.n186 0.155672
R478 VTAIL.n195 VTAIL.n186 0.155672
R479 VTAIL.n195 VTAIL.n194 0.155672
R480 VTAIL.n161 VTAIL.n83 0.155672
R481 VTAIL.n153 VTAIL.n83 0.155672
R482 VTAIL.n153 VTAIL.n152 0.155672
R483 VTAIL.n152 VTAIL.n87 0.155672
R484 VTAIL.n145 VTAIL.n87 0.155672
R485 VTAIL.n145 VTAIL.n144 0.155672
R486 VTAIL.n144 VTAIL.n92 0.155672
R487 VTAIL.n137 VTAIL.n92 0.155672
R488 VTAIL.n137 VTAIL.n136 0.155672
R489 VTAIL.n136 VTAIL.n96 0.155672
R490 VTAIL.n129 VTAIL.n96 0.155672
R491 VTAIL.n129 VTAIL.n128 0.155672
R492 VTAIL.n128 VTAIL.n100 0.155672
R493 VTAIL.n121 VTAIL.n100 0.155672
R494 VTAIL.n121 VTAIL.n120 0.155672
R495 VTAIL.n120 VTAIL.n104 0.155672
R496 VTAIL.n113 VTAIL.n104 0.155672
R497 VTAIL.n113 VTAIL.n112 0.155672
R498 VTAIL VTAIL.n327 0.140586
R499 VDD2.n157 VDD2.n81 289.615
R500 VDD2.n76 VDD2.n0 289.615
R501 VDD2.n158 VDD2.n157 185
R502 VDD2.n156 VDD2.n155 185
R503 VDD2.n154 VDD2.n84 185
R504 VDD2.n88 VDD2.n85 185
R505 VDD2.n149 VDD2.n148 185
R506 VDD2.n147 VDD2.n146 185
R507 VDD2.n90 VDD2.n89 185
R508 VDD2.n141 VDD2.n140 185
R509 VDD2.n139 VDD2.n138 185
R510 VDD2.n94 VDD2.n93 185
R511 VDD2.n133 VDD2.n132 185
R512 VDD2.n131 VDD2.n130 185
R513 VDD2.n98 VDD2.n97 185
R514 VDD2.n125 VDD2.n124 185
R515 VDD2.n123 VDD2.n122 185
R516 VDD2.n102 VDD2.n101 185
R517 VDD2.n117 VDD2.n116 185
R518 VDD2.n115 VDD2.n114 185
R519 VDD2.n106 VDD2.n105 185
R520 VDD2.n109 VDD2.n108 185
R521 VDD2.n27 VDD2.n26 185
R522 VDD2.n24 VDD2.n23 185
R523 VDD2.n33 VDD2.n32 185
R524 VDD2.n35 VDD2.n34 185
R525 VDD2.n20 VDD2.n19 185
R526 VDD2.n41 VDD2.n40 185
R527 VDD2.n43 VDD2.n42 185
R528 VDD2.n16 VDD2.n15 185
R529 VDD2.n49 VDD2.n48 185
R530 VDD2.n51 VDD2.n50 185
R531 VDD2.n12 VDD2.n11 185
R532 VDD2.n57 VDD2.n56 185
R533 VDD2.n59 VDD2.n58 185
R534 VDD2.n8 VDD2.n7 185
R535 VDD2.n65 VDD2.n64 185
R536 VDD2.n68 VDD2.n67 185
R537 VDD2.n66 VDD2.n4 185
R538 VDD2.n73 VDD2.n3 185
R539 VDD2.n75 VDD2.n74 185
R540 VDD2.n77 VDD2.n76 185
R541 VDD2.t1 VDD2.n107 147.659
R542 VDD2.t0 VDD2.n25 147.659
R543 VDD2.n157 VDD2.n156 104.615
R544 VDD2.n156 VDD2.n84 104.615
R545 VDD2.n88 VDD2.n84 104.615
R546 VDD2.n148 VDD2.n88 104.615
R547 VDD2.n148 VDD2.n147 104.615
R548 VDD2.n147 VDD2.n89 104.615
R549 VDD2.n140 VDD2.n89 104.615
R550 VDD2.n140 VDD2.n139 104.615
R551 VDD2.n139 VDD2.n93 104.615
R552 VDD2.n132 VDD2.n93 104.615
R553 VDD2.n132 VDD2.n131 104.615
R554 VDD2.n131 VDD2.n97 104.615
R555 VDD2.n124 VDD2.n97 104.615
R556 VDD2.n124 VDD2.n123 104.615
R557 VDD2.n123 VDD2.n101 104.615
R558 VDD2.n116 VDD2.n101 104.615
R559 VDD2.n116 VDD2.n115 104.615
R560 VDD2.n115 VDD2.n105 104.615
R561 VDD2.n108 VDD2.n105 104.615
R562 VDD2.n26 VDD2.n23 104.615
R563 VDD2.n33 VDD2.n23 104.615
R564 VDD2.n34 VDD2.n33 104.615
R565 VDD2.n34 VDD2.n19 104.615
R566 VDD2.n41 VDD2.n19 104.615
R567 VDD2.n42 VDD2.n41 104.615
R568 VDD2.n42 VDD2.n15 104.615
R569 VDD2.n49 VDD2.n15 104.615
R570 VDD2.n50 VDD2.n49 104.615
R571 VDD2.n50 VDD2.n11 104.615
R572 VDD2.n57 VDD2.n11 104.615
R573 VDD2.n58 VDD2.n57 104.615
R574 VDD2.n58 VDD2.n7 104.615
R575 VDD2.n65 VDD2.n7 104.615
R576 VDD2.n67 VDD2.n65 104.615
R577 VDD2.n67 VDD2.n66 104.615
R578 VDD2.n66 VDD2.n3 104.615
R579 VDD2.n75 VDD2.n3 104.615
R580 VDD2.n76 VDD2.n75 104.615
R581 VDD2.n162 VDD2.n80 91.4066
R582 VDD2.n162 VDD2.n161 53.3247
R583 VDD2.n108 VDD2.t1 52.3082
R584 VDD2.n26 VDD2.t0 52.3082
R585 VDD2.n109 VDD2.n107 15.6677
R586 VDD2.n27 VDD2.n25 15.6677
R587 VDD2.n155 VDD2.n154 13.1884
R588 VDD2.n74 VDD2.n73 13.1884
R589 VDD2.n158 VDD2.n83 12.8005
R590 VDD2.n153 VDD2.n85 12.8005
R591 VDD2.n110 VDD2.n106 12.8005
R592 VDD2.n28 VDD2.n24 12.8005
R593 VDD2.n72 VDD2.n4 12.8005
R594 VDD2.n77 VDD2.n2 12.8005
R595 VDD2.n159 VDD2.n81 12.0247
R596 VDD2.n150 VDD2.n149 12.0247
R597 VDD2.n114 VDD2.n113 12.0247
R598 VDD2.n32 VDD2.n31 12.0247
R599 VDD2.n69 VDD2.n68 12.0247
R600 VDD2.n78 VDD2.n0 12.0247
R601 VDD2.n146 VDD2.n87 11.249
R602 VDD2.n117 VDD2.n104 11.249
R603 VDD2.n35 VDD2.n22 11.249
R604 VDD2.n64 VDD2.n6 11.249
R605 VDD2.n145 VDD2.n90 10.4732
R606 VDD2.n118 VDD2.n102 10.4732
R607 VDD2.n36 VDD2.n20 10.4732
R608 VDD2.n63 VDD2.n8 10.4732
R609 VDD2.n142 VDD2.n141 9.69747
R610 VDD2.n122 VDD2.n121 9.69747
R611 VDD2.n40 VDD2.n39 9.69747
R612 VDD2.n60 VDD2.n59 9.69747
R613 VDD2.n161 VDD2.n160 9.45567
R614 VDD2.n80 VDD2.n79 9.45567
R615 VDD2.n135 VDD2.n134 9.3005
R616 VDD2.n137 VDD2.n136 9.3005
R617 VDD2.n92 VDD2.n91 9.3005
R618 VDD2.n143 VDD2.n142 9.3005
R619 VDD2.n145 VDD2.n144 9.3005
R620 VDD2.n87 VDD2.n86 9.3005
R621 VDD2.n151 VDD2.n150 9.3005
R622 VDD2.n153 VDD2.n152 9.3005
R623 VDD2.n160 VDD2.n159 9.3005
R624 VDD2.n83 VDD2.n82 9.3005
R625 VDD2.n96 VDD2.n95 9.3005
R626 VDD2.n129 VDD2.n128 9.3005
R627 VDD2.n127 VDD2.n126 9.3005
R628 VDD2.n100 VDD2.n99 9.3005
R629 VDD2.n121 VDD2.n120 9.3005
R630 VDD2.n119 VDD2.n118 9.3005
R631 VDD2.n104 VDD2.n103 9.3005
R632 VDD2.n113 VDD2.n112 9.3005
R633 VDD2.n111 VDD2.n110 9.3005
R634 VDD2.n79 VDD2.n78 9.3005
R635 VDD2.n2 VDD2.n1 9.3005
R636 VDD2.n47 VDD2.n46 9.3005
R637 VDD2.n45 VDD2.n44 9.3005
R638 VDD2.n18 VDD2.n17 9.3005
R639 VDD2.n39 VDD2.n38 9.3005
R640 VDD2.n37 VDD2.n36 9.3005
R641 VDD2.n22 VDD2.n21 9.3005
R642 VDD2.n31 VDD2.n30 9.3005
R643 VDD2.n29 VDD2.n28 9.3005
R644 VDD2.n14 VDD2.n13 9.3005
R645 VDD2.n53 VDD2.n52 9.3005
R646 VDD2.n55 VDD2.n54 9.3005
R647 VDD2.n10 VDD2.n9 9.3005
R648 VDD2.n61 VDD2.n60 9.3005
R649 VDD2.n63 VDD2.n62 9.3005
R650 VDD2.n6 VDD2.n5 9.3005
R651 VDD2.n70 VDD2.n69 9.3005
R652 VDD2.n72 VDD2.n71 9.3005
R653 VDD2.n138 VDD2.n92 8.92171
R654 VDD2.n125 VDD2.n100 8.92171
R655 VDD2.n43 VDD2.n18 8.92171
R656 VDD2.n56 VDD2.n10 8.92171
R657 VDD2.n137 VDD2.n94 8.14595
R658 VDD2.n126 VDD2.n98 8.14595
R659 VDD2.n44 VDD2.n16 8.14595
R660 VDD2.n55 VDD2.n12 8.14595
R661 VDD2.n134 VDD2.n133 7.3702
R662 VDD2.n130 VDD2.n129 7.3702
R663 VDD2.n48 VDD2.n47 7.3702
R664 VDD2.n52 VDD2.n51 7.3702
R665 VDD2.n133 VDD2.n96 6.59444
R666 VDD2.n130 VDD2.n96 6.59444
R667 VDD2.n48 VDD2.n14 6.59444
R668 VDD2.n51 VDD2.n14 6.59444
R669 VDD2.n134 VDD2.n94 5.81868
R670 VDD2.n129 VDD2.n98 5.81868
R671 VDD2.n47 VDD2.n16 5.81868
R672 VDD2.n52 VDD2.n12 5.81868
R673 VDD2.n138 VDD2.n137 5.04292
R674 VDD2.n126 VDD2.n125 5.04292
R675 VDD2.n44 VDD2.n43 5.04292
R676 VDD2.n56 VDD2.n55 5.04292
R677 VDD2.n111 VDD2.n107 4.38563
R678 VDD2.n29 VDD2.n25 4.38563
R679 VDD2.n141 VDD2.n92 4.26717
R680 VDD2.n122 VDD2.n100 4.26717
R681 VDD2.n40 VDD2.n18 4.26717
R682 VDD2.n59 VDD2.n10 4.26717
R683 VDD2.n142 VDD2.n90 3.49141
R684 VDD2.n121 VDD2.n102 3.49141
R685 VDD2.n39 VDD2.n20 3.49141
R686 VDD2.n60 VDD2.n8 3.49141
R687 VDD2.n146 VDD2.n145 2.71565
R688 VDD2.n118 VDD2.n117 2.71565
R689 VDD2.n36 VDD2.n35 2.71565
R690 VDD2.n64 VDD2.n63 2.71565
R691 VDD2.n161 VDD2.n81 1.93989
R692 VDD2.n149 VDD2.n87 1.93989
R693 VDD2.n114 VDD2.n104 1.93989
R694 VDD2.n32 VDD2.n22 1.93989
R695 VDD2.n68 VDD2.n6 1.93989
R696 VDD2.n80 VDD2.n0 1.93989
R697 VDD2.n159 VDD2.n158 1.16414
R698 VDD2.n150 VDD2.n85 1.16414
R699 VDD2.n113 VDD2.n106 1.16414
R700 VDD2.n31 VDD2.n24 1.16414
R701 VDD2.n69 VDD2.n4 1.16414
R702 VDD2.n78 VDD2.n77 1.16414
R703 VDD2.n155 VDD2.n83 0.388379
R704 VDD2.n154 VDD2.n153 0.388379
R705 VDD2.n110 VDD2.n109 0.388379
R706 VDD2.n28 VDD2.n27 0.388379
R707 VDD2.n73 VDD2.n72 0.388379
R708 VDD2.n74 VDD2.n2 0.388379
R709 VDD2 VDD2.n162 0.256966
R710 VDD2.n160 VDD2.n82 0.155672
R711 VDD2.n152 VDD2.n82 0.155672
R712 VDD2.n152 VDD2.n151 0.155672
R713 VDD2.n151 VDD2.n86 0.155672
R714 VDD2.n144 VDD2.n86 0.155672
R715 VDD2.n144 VDD2.n143 0.155672
R716 VDD2.n143 VDD2.n91 0.155672
R717 VDD2.n136 VDD2.n91 0.155672
R718 VDD2.n136 VDD2.n135 0.155672
R719 VDD2.n135 VDD2.n95 0.155672
R720 VDD2.n128 VDD2.n95 0.155672
R721 VDD2.n128 VDD2.n127 0.155672
R722 VDD2.n127 VDD2.n99 0.155672
R723 VDD2.n120 VDD2.n99 0.155672
R724 VDD2.n120 VDD2.n119 0.155672
R725 VDD2.n119 VDD2.n103 0.155672
R726 VDD2.n112 VDD2.n103 0.155672
R727 VDD2.n112 VDD2.n111 0.155672
R728 VDD2.n30 VDD2.n29 0.155672
R729 VDD2.n30 VDD2.n21 0.155672
R730 VDD2.n37 VDD2.n21 0.155672
R731 VDD2.n38 VDD2.n37 0.155672
R732 VDD2.n38 VDD2.n17 0.155672
R733 VDD2.n45 VDD2.n17 0.155672
R734 VDD2.n46 VDD2.n45 0.155672
R735 VDD2.n46 VDD2.n13 0.155672
R736 VDD2.n53 VDD2.n13 0.155672
R737 VDD2.n54 VDD2.n53 0.155672
R738 VDD2.n54 VDD2.n9 0.155672
R739 VDD2.n61 VDD2.n9 0.155672
R740 VDD2.n62 VDD2.n61 0.155672
R741 VDD2.n62 VDD2.n5 0.155672
R742 VDD2.n70 VDD2.n5 0.155672
R743 VDD2.n71 VDD2.n70 0.155672
R744 VDD2.n71 VDD2.n1 0.155672
R745 VDD2.n79 VDD2.n1 0.155672
R746 B.n87 B.t2 811.971
R747 B.n84 B.t6 811.971
R748 B.n389 B.t13 811.971
R749 B.n387 B.t9 811.971
R750 B.n670 B.n669 585
R751 B.n306 B.n83 585
R752 B.n305 B.n304 585
R753 B.n303 B.n302 585
R754 B.n301 B.n300 585
R755 B.n299 B.n298 585
R756 B.n297 B.n296 585
R757 B.n295 B.n294 585
R758 B.n293 B.n292 585
R759 B.n291 B.n290 585
R760 B.n289 B.n288 585
R761 B.n287 B.n286 585
R762 B.n285 B.n284 585
R763 B.n283 B.n282 585
R764 B.n281 B.n280 585
R765 B.n279 B.n278 585
R766 B.n277 B.n276 585
R767 B.n275 B.n274 585
R768 B.n273 B.n272 585
R769 B.n271 B.n270 585
R770 B.n269 B.n268 585
R771 B.n267 B.n266 585
R772 B.n265 B.n264 585
R773 B.n263 B.n262 585
R774 B.n261 B.n260 585
R775 B.n259 B.n258 585
R776 B.n257 B.n256 585
R777 B.n255 B.n254 585
R778 B.n253 B.n252 585
R779 B.n251 B.n250 585
R780 B.n249 B.n248 585
R781 B.n247 B.n246 585
R782 B.n245 B.n244 585
R783 B.n243 B.n242 585
R784 B.n241 B.n240 585
R785 B.n239 B.n238 585
R786 B.n237 B.n236 585
R787 B.n235 B.n234 585
R788 B.n233 B.n232 585
R789 B.n231 B.n230 585
R790 B.n229 B.n228 585
R791 B.n227 B.n226 585
R792 B.n225 B.n224 585
R793 B.n223 B.n222 585
R794 B.n221 B.n220 585
R795 B.n219 B.n218 585
R796 B.n217 B.n216 585
R797 B.n215 B.n214 585
R798 B.n213 B.n212 585
R799 B.n211 B.n210 585
R800 B.n209 B.n208 585
R801 B.n207 B.n206 585
R802 B.n205 B.n204 585
R803 B.n203 B.n202 585
R804 B.n201 B.n200 585
R805 B.n199 B.n198 585
R806 B.n197 B.n196 585
R807 B.n195 B.n194 585
R808 B.n193 B.n192 585
R809 B.n191 B.n190 585
R810 B.n189 B.n188 585
R811 B.n187 B.n186 585
R812 B.n185 B.n184 585
R813 B.n183 B.n182 585
R814 B.n181 B.n180 585
R815 B.n179 B.n178 585
R816 B.n177 B.n176 585
R817 B.n175 B.n174 585
R818 B.n173 B.n172 585
R819 B.n171 B.n170 585
R820 B.n169 B.n168 585
R821 B.n167 B.n166 585
R822 B.n165 B.n164 585
R823 B.n163 B.n162 585
R824 B.n161 B.n160 585
R825 B.n159 B.n158 585
R826 B.n157 B.n156 585
R827 B.n155 B.n154 585
R828 B.n153 B.n152 585
R829 B.n151 B.n150 585
R830 B.n149 B.n148 585
R831 B.n147 B.n146 585
R832 B.n145 B.n144 585
R833 B.n143 B.n142 585
R834 B.n141 B.n140 585
R835 B.n139 B.n138 585
R836 B.n137 B.n136 585
R837 B.n135 B.n134 585
R838 B.n133 B.n132 585
R839 B.n131 B.n130 585
R840 B.n129 B.n128 585
R841 B.n127 B.n126 585
R842 B.n125 B.n124 585
R843 B.n123 B.n122 585
R844 B.n121 B.n120 585
R845 B.n119 B.n118 585
R846 B.n117 B.n116 585
R847 B.n115 B.n114 585
R848 B.n113 B.n112 585
R849 B.n111 B.n110 585
R850 B.n109 B.n108 585
R851 B.n107 B.n106 585
R852 B.n105 B.n104 585
R853 B.n103 B.n102 585
R854 B.n101 B.n100 585
R855 B.n99 B.n98 585
R856 B.n97 B.n96 585
R857 B.n95 B.n94 585
R858 B.n93 B.n92 585
R859 B.n91 B.n90 585
R860 B.n668 B.n28 585
R861 B.n673 B.n28 585
R862 B.n667 B.n27 585
R863 B.n674 B.n27 585
R864 B.n666 B.n665 585
R865 B.n665 B.n23 585
R866 B.n664 B.n22 585
R867 B.n680 B.n22 585
R868 B.n663 B.n21 585
R869 B.n681 B.n21 585
R870 B.n662 B.n20 585
R871 B.n682 B.n20 585
R872 B.n661 B.n660 585
R873 B.n660 B.n16 585
R874 B.n659 B.n15 585
R875 B.n688 B.n15 585
R876 B.n658 B.n14 585
R877 B.n689 B.n14 585
R878 B.n657 B.n13 585
R879 B.n690 B.n13 585
R880 B.n656 B.n655 585
R881 B.n655 B.n12 585
R882 B.n654 B.n653 585
R883 B.n654 B.n8 585
R884 B.n652 B.n7 585
R885 B.n697 B.n7 585
R886 B.n651 B.n6 585
R887 B.n698 B.n6 585
R888 B.n650 B.n5 585
R889 B.n699 B.n5 585
R890 B.n649 B.n648 585
R891 B.n648 B.n4 585
R892 B.n647 B.n307 585
R893 B.n647 B.n646 585
R894 B.n636 B.n308 585
R895 B.n639 B.n308 585
R896 B.n638 B.n637 585
R897 B.n640 B.n638 585
R898 B.n635 B.n313 585
R899 B.n313 B.n312 585
R900 B.n634 B.n633 585
R901 B.n633 B.n632 585
R902 B.n315 B.n314 585
R903 B.n316 B.n315 585
R904 B.n625 B.n624 585
R905 B.n626 B.n625 585
R906 B.n623 B.n320 585
R907 B.n324 B.n320 585
R908 B.n622 B.n621 585
R909 B.n621 B.n620 585
R910 B.n322 B.n321 585
R911 B.n323 B.n322 585
R912 B.n613 B.n612 585
R913 B.n614 B.n613 585
R914 B.n611 B.n329 585
R915 B.n329 B.n328 585
R916 B.n606 B.n605 585
R917 B.n604 B.n386 585
R918 B.n603 B.n385 585
R919 B.n608 B.n385 585
R920 B.n602 B.n601 585
R921 B.n600 B.n599 585
R922 B.n598 B.n597 585
R923 B.n596 B.n595 585
R924 B.n594 B.n593 585
R925 B.n592 B.n591 585
R926 B.n590 B.n589 585
R927 B.n588 B.n587 585
R928 B.n586 B.n585 585
R929 B.n584 B.n583 585
R930 B.n582 B.n581 585
R931 B.n580 B.n579 585
R932 B.n578 B.n577 585
R933 B.n576 B.n575 585
R934 B.n574 B.n573 585
R935 B.n572 B.n571 585
R936 B.n570 B.n569 585
R937 B.n568 B.n567 585
R938 B.n566 B.n565 585
R939 B.n564 B.n563 585
R940 B.n562 B.n561 585
R941 B.n560 B.n559 585
R942 B.n558 B.n557 585
R943 B.n556 B.n555 585
R944 B.n554 B.n553 585
R945 B.n552 B.n551 585
R946 B.n550 B.n549 585
R947 B.n548 B.n547 585
R948 B.n546 B.n545 585
R949 B.n544 B.n543 585
R950 B.n542 B.n541 585
R951 B.n540 B.n539 585
R952 B.n538 B.n537 585
R953 B.n536 B.n535 585
R954 B.n534 B.n533 585
R955 B.n532 B.n531 585
R956 B.n530 B.n529 585
R957 B.n528 B.n527 585
R958 B.n526 B.n525 585
R959 B.n524 B.n523 585
R960 B.n522 B.n521 585
R961 B.n520 B.n519 585
R962 B.n518 B.n517 585
R963 B.n516 B.n515 585
R964 B.n514 B.n513 585
R965 B.n512 B.n511 585
R966 B.n510 B.n509 585
R967 B.n507 B.n506 585
R968 B.n505 B.n504 585
R969 B.n503 B.n502 585
R970 B.n501 B.n500 585
R971 B.n499 B.n498 585
R972 B.n497 B.n496 585
R973 B.n495 B.n494 585
R974 B.n493 B.n492 585
R975 B.n491 B.n490 585
R976 B.n489 B.n488 585
R977 B.n486 B.n485 585
R978 B.n484 B.n483 585
R979 B.n482 B.n481 585
R980 B.n480 B.n479 585
R981 B.n478 B.n477 585
R982 B.n476 B.n475 585
R983 B.n474 B.n473 585
R984 B.n472 B.n471 585
R985 B.n470 B.n469 585
R986 B.n468 B.n467 585
R987 B.n466 B.n465 585
R988 B.n464 B.n463 585
R989 B.n462 B.n461 585
R990 B.n460 B.n459 585
R991 B.n458 B.n457 585
R992 B.n456 B.n455 585
R993 B.n454 B.n453 585
R994 B.n452 B.n451 585
R995 B.n450 B.n449 585
R996 B.n448 B.n447 585
R997 B.n446 B.n445 585
R998 B.n444 B.n443 585
R999 B.n442 B.n441 585
R1000 B.n440 B.n439 585
R1001 B.n438 B.n437 585
R1002 B.n436 B.n435 585
R1003 B.n434 B.n433 585
R1004 B.n432 B.n431 585
R1005 B.n430 B.n429 585
R1006 B.n428 B.n427 585
R1007 B.n426 B.n425 585
R1008 B.n424 B.n423 585
R1009 B.n422 B.n421 585
R1010 B.n420 B.n419 585
R1011 B.n418 B.n417 585
R1012 B.n416 B.n415 585
R1013 B.n414 B.n413 585
R1014 B.n412 B.n411 585
R1015 B.n410 B.n409 585
R1016 B.n408 B.n407 585
R1017 B.n406 B.n405 585
R1018 B.n404 B.n403 585
R1019 B.n402 B.n401 585
R1020 B.n400 B.n399 585
R1021 B.n398 B.n397 585
R1022 B.n396 B.n395 585
R1023 B.n394 B.n393 585
R1024 B.n392 B.n391 585
R1025 B.n331 B.n330 585
R1026 B.n610 B.n609 585
R1027 B.n609 B.n608 585
R1028 B.n327 B.n326 585
R1029 B.n328 B.n327 585
R1030 B.n616 B.n615 585
R1031 B.n615 B.n614 585
R1032 B.n617 B.n325 585
R1033 B.n325 B.n323 585
R1034 B.n619 B.n618 585
R1035 B.n620 B.n619 585
R1036 B.n319 B.n318 585
R1037 B.n324 B.n319 585
R1038 B.n628 B.n627 585
R1039 B.n627 B.n626 585
R1040 B.n629 B.n317 585
R1041 B.n317 B.n316 585
R1042 B.n631 B.n630 585
R1043 B.n632 B.n631 585
R1044 B.n311 B.n310 585
R1045 B.n312 B.n311 585
R1046 B.n642 B.n641 585
R1047 B.n641 B.n640 585
R1048 B.n643 B.n309 585
R1049 B.n639 B.n309 585
R1050 B.n645 B.n644 585
R1051 B.n646 B.n645 585
R1052 B.n3 B.n0 585
R1053 B.n4 B.n3 585
R1054 B.n696 B.n1 585
R1055 B.n697 B.n696 585
R1056 B.n695 B.n694 585
R1057 B.n695 B.n8 585
R1058 B.n693 B.n9 585
R1059 B.n12 B.n9 585
R1060 B.n692 B.n691 585
R1061 B.n691 B.n690 585
R1062 B.n11 B.n10 585
R1063 B.n689 B.n11 585
R1064 B.n687 B.n686 585
R1065 B.n688 B.n687 585
R1066 B.n685 B.n17 585
R1067 B.n17 B.n16 585
R1068 B.n684 B.n683 585
R1069 B.n683 B.n682 585
R1070 B.n19 B.n18 585
R1071 B.n681 B.n19 585
R1072 B.n679 B.n678 585
R1073 B.n680 B.n679 585
R1074 B.n677 B.n24 585
R1075 B.n24 B.n23 585
R1076 B.n676 B.n675 585
R1077 B.n675 B.n674 585
R1078 B.n26 B.n25 585
R1079 B.n673 B.n26 585
R1080 B.n700 B.n699 585
R1081 B.n698 B.n2 585
R1082 B.n90 B.n26 487.695
R1083 B.n670 B.n28 487.695
R1084 B.n609 B.n329 487.695
R1085 B.n606 B.n327 487.695
R1086 B.n84 B.t7 349.61
R1087 B.n389 B.t15 349.61
R1088 B.n87 B.t4 349.61
R1089 B.n387 B.t12 349.61
R1090 B.n85 B.t8 331.767
R1091 B.n390 B.t14 331.767
R1092 B.n88 B.t5 331.767
R1093 B.n388 B.t11 331.767
R1094 B.n672 B.n671 256.663
R1095 B.n672 B.n82 256.663
R1096 B.n672 B.n81 256.663
R1097 B.n672 B.n80 256.663
R1098 B.n672 B.n79 256.663
R1099 B.n672 B.n78 256.663
R1100 B.n672 B.n77 256.663
R1101 B.n672 B.n76 256.663
R1102 B.n672 B.n75 256.663
R1103 B.n672 B.n74 256.663
R1104 B.n672 B.n73 256.663
R1105 B.n672 B.n72 256.663
R1106 B.n672 B.n71 256.663
R1107 B.n672 B.n70 256.663
R1108 B.n672 B.n69 256.663
R1109 B.n672 B.n68 256.663
R1110 B.n672 B.n67 256.663
R1111 B.n672 B.n66 256.663
R1112 B.n672 B.n65 256.663
R1113 B.n672 B.n64 256.663
R1114 B.n672 B.n63 256.663
R1115 B.n672 B.n62 256.663
R1116 B.n672 B.n61 256.663
R1117 B.n672 B.n60 256.663
R1118 B.n672 B.n59 256.663
R1119 B.n672 B.n58 256.663
R1120 B.n672 B.n57 256.663
R1121 B.n672 B.n56 256.663
R1122 B.n672 B.n55 256.663
R1123 B.n672 B.n54 256.663
R1124 B.n672 B.n53 256.663
R1125 B.n672 B.n52 256.663
R1126 B.n672 B.n51 256.663
R1127 B.n672 B.n50 256.663
R1128 B.n672 B.n49 256.663
R1129 B.n672 B.n48 256.663
R1130 B.n672 B.n47 256.663
R1131 B.n672 B.n46 256.663
R1132 B.n672 B.n45 256.663
R1133 B.n672 B.n44 256.663
R1134 B.n672 B.n43 256.663
R1135 B.n672 B.n42 256.663
R1136 B.n672 B.n41 256.663
R1137 B.n672 B.n40 256.663
R1138 B.n672 B.n39 256.663
R1139 B.n672 B.n38 256.663
R1140 B.n672 B.n37 256.663
R1141 B.n672 B.n36 256.663
R1142 B.n672 B.n35 256.663
R1143 B.n672 B.n34 256.663
R1144 B.n672 B.n33 256.663
R1145 B.n672 B.n32 256.663
R1146 B.n672 B.n31 256.663
R1147 B.n672 B.n30 256.663
R1148 B.n672 B.n29 256.663
R1149 B.n608 B.n607 256.663
R1150 B.n608 B.n332 256.663
R1151 B.n608 B.n333 256.663
R1152 B.n608 B.n334 256.663
R1153 B.n608 B.n335 256.663
R1154 B.n608 B.n336 256.663
R1155 B.n608 B.n337 256.663
R1156 B.n608 B.n338 256.663
R1157 B.n608 B.n339 256.663
R1158 B.n608 B.n340 256.663
R1159 B.n608 B.n341 256.663
R1160 B.n608 B.n342 256.663
R1161 B.n608 B.n343 256.663
R1162 B.n608 B.n344 256.663
R1163 B.n608 B.n345 256.663
R1164 B.n608 B.n346 256.663
R1165 B.n608 B.n347 256.663
R1166 B.n608 B.n348 256.663
R1167 B.n608 B.n349 256.663
R1168 B.n608 B.n350 256.663
R1169 B.n608 B.n351 256.663
R1170 B.n608 B.n352 256.663
R1171 B.n608 B.n353 256.663
R1172 B.n608 B.n354 256.663
R1173 B.n608 B.n355 256.663
R1174 B.n608 B.n356 256.663
R1175 B.n608 B.n357 256.663
R1176 B.n608 B.n358 256.663
R1177 B.n608 B.n359 256.663
R1178 B.n608 B.n360 256.663
R1179 B.n608 B.n361 256.663
R1180 B.n608 B.n362 256.663
R1181 B.n608 B.n363 256.663
R1182 B.n608 B.n364 256.663
R1183 B.n608 B.n365 256.663
R1184 B.n608 B.n366 256.663
R1185 B.n608 B.n367 256.663
R1186 B.n608 B.n368 256.663
R1187 B.n608 B.n369 256.663
R1188 B.n608 B.n370 256.663
R1189 B.n608 B.n371 256.663
R1190 B.n608 B.n372 256.663
R1191 B.n608 B.n373 256.663
R1192 B.n608 B.n374 256.663
R1193 B.n608 B.n375 256.663
R1194 B.n608 B.n376 256.663
R1195 B.n608 B.n377 256.663
R1196 B.n608 B.n378 256.663
R1197 B.n608 B.n379 256.663
R1198 B.n608 B.n380 256.663
R1199 B.n608 B.n381 256.663
R1200 B.n608 B.n382 256.663
R1201 B.n608 B.n383 256.663
R1202 B.n608 B.n384 256.663
R1203 B.n702 B.n701 256.663
R1204 B.n94 B.n93 163.367
R1205 B.n98 B.n97 163.367
R1206 B.n102 B.n101 163.367
R1207 B.n106 B.n105 163.367
R1208 B.n110 B.n109 163.367
R1209 B.n114 B.n113 163.367
R1210 B.n118 B.n117 163.367
R1211 B.n122 B.n121 163.367
R1212 B.n126 B.n125 163.367
R1213 B.n130 B.n129 163.367
R1214 B.n134 B.n133 163.367
R1215 B.n138 B.n137 163.367
R1216 B.n142 B.n141 163.367
R1217 B.n146 B.n145 163.367
R1218 B.n150 B.n149 163.367
R1219 B.n154 B.n153 163.367
R1220 B.n158 B.n157 163.367
R1221 B.n162 B.n161 163.367
R1222 B.n166 B.n165 163.367
R1223 B.n170 B.n169 163.367
R1224 B.n174 B.n173 163.367
R1225 B.n178 B.n177 163.367
R1226 B.n182 B.n181 163.367
R1227 B.n186 B.n185 163.367
R1228 B.n190 B.n189 163.367
R1229 B.n194 B.n193 163.367
R1230 B.n198 B.n197 163.367
R1231 B.n202 B.n201 163.367
R1232 B.n206 B.n205 163.367
R1233 B.n210 B.n209 163.367
R1234 B.n214 B.n213 163.367
R1235 B.n218 B.n217 163.367
R1236 B.n222 B.n221 163.367
R1237 B.n226 B.n225 163.367
R1238 B.n230 B.n229 163.367
R1239 B.n234 B.n233 163.367
R1240 B.n238 B.n237 163.367
R1241 B.n242 B.n241 163.367
R1242 B.n246 B.n245 163.367
R1243 B.n250 B.n249 163.367
R1244 B.n254 B.n253 163.367
R1245 B.n258 B.n257 163.367
R1246 B.n262 B.n261 163.367
R1247 B.n266 B.n265 163.367
R1248 B.n270 B.n269 163.367
R1249 B.n274 B.n273 163.367
R1250 B.n278 B.n277 163.367
R1251 B.n282 B.n281 163.367
R1252 B.n286 B.n285 163.367
R1253 B.n290 B.n289 163.367
R1254 B.n294 B.n293 163.367
R1255 B.n298 B.n297 163.367
R1256 B.n302 B.n301 163.367
R1257 B.n304 B.n83 163.367
R1258 B.n613 B.n329 163.367
R1259 B.n613 B.n322 163.367
R1260 B.n621 B.n322 163.367
R1261 B.n621 B.n320 163.367
R1262 B.n625 B.n320 163.367
R1263 B.n625 B.n315 163.367
R1264 B.n633 B.n315 163.367
R1265 B.n633 B.n313 163.367
R1266 B.n638 B.n313 163.367
R1267 B.n638 B.n308 163.367
R1268 B.n647 B.n308 163.367
R1269 B.n648 B.n647 163.367
R1270 B.n648 B.n5 163.367
R1271 B.n6 B.n5 163.367
R1272 B.n7 B.n6 163.367
R1273 B.n654 B.n7 163.367
R1274 B.n655 B.n654 163.367
R1275 B.n655 B.n13 163.367
R1276 B.n14 B.n13 163.367
R1277 B.n15 B.n14 163.367
R1278 B.n660 B.n15 163.367
R1279 B.n660 B.n20 163.367
R1280 B.n21 B.n20 163.367
R1281 B.n22 B.n21 163.367
R1282 B.n665 B.n22 163.367
R1283 B.n665 B.n27 163.367
R1284 B.n28 B.n27 163.367
R1285 B.n386 B.n385 163.367
R1286 B.n601 B.n385 163.367
R1287 B.n599 B.n598 163.367
R1288 B.n595 B.n594 163.367
R1289 B.n591 B.n590 163.367
R1290 B.n587 B.n586 163.367
R1291 B.n583 B.n582 163.367
R1292 B.n579 B.n578 163.367
R1293 B.n575 B.n574 163.367
R1294 B.n571 B.n570 163.367
R1295 B.n567 B.n566 163.367
R1296 B.n563 B.n562 163.367
R1297 B.n559 B.n558 163.367
R1298 B.n555 B.n554 163.367
R1299 B.n551 B.n550 163.367
R1300 B.n547 B.n546 163.367
R1301 B.n543 B.n542 163.367
R1302 B.n539 B.n538 163.367
R1303 B.n535 B.n534 163.367
R1304 B.n531 B.n530 163.367
R1305 B.n527 B.n526 163.367
R1306 B.n523 B.n522 163.367
R1307 B.n519 B.n518 163.367
R1308 B.n515 B.n514 163.367
R1309 B.n511 B.n510 163.367
R1310 B.n506 B.n505 163.367
R1311 B.n502 B.n501 163.367
R1312 B.n498 B.n497 163.367
R1313 B.n494 B.n493 163.367
R1314 B.n490 B.n489 163.367
R1315 B.n485 B.n484 163.367
R1316 B.n481 B.n480 163.367
R1317 B.n477 B.n476 163.367
R1318 B.n473 B.n472 163.367
R1319 B.n469 B.n468 163.367
R1320 B.n465 B.n464 163.367
R1321 B.n461 B.n460 163.367
R1322 B.n457 B.n456 163.367
R1323 B.n453 B.n452 163.367
R1324 B.n449 B.n448 163.367
R1325 B.n445 B.n444 163.367
R1326 B.n441 B.n440 163.367
R1327 B.n437 B.n436 163.367
R1328 B.n433 B.n432 163.367
R1329 B.n429 B.n428 163.367
R1330 B.n425 B.n424 163.367
R1331 B.n421 B.n420 163.367
R1332 B.n417 B.n416 163.367
R1333 B.n413 B.n412 163.367
R1334 B.n409 B.n408 163.367
R1335 B.n405 B.n404 163.367
R1336 B.n401 B.n400 163.367
R1337 B.n397 B.n396 163.367
R1338 B.n393 B.n392 163.367
R1339 B.n609 B.n331 163.367
R1340 B.n615 B.n327 163.367
R1341 B.n615 B.n325 163.367
R1342 B.n619 B.n325 163.367
R1343 B.n619 B.n319 163.367
R1344 B.n627 B.n319 163.367
R1345 B.n627 B.n317 163.367
R1346 B.n631 B.n317 163.367
R1347 B.n631 B.n311 163.367
R1348 B.n641 B.n311 163.367
R1349 B.n641 B.n309 163.367
R1350 B.n645 B.n309 163.367
R1351 B.n645 B.n3 163.367
R1352 B.n700 B.n3 163.367
R1353 B.n696 B.n2 163.367
R1354 B.n696 B.n695 163.367
R1355 B.n695 B.n9 163.367
R1356 B.n691 B.n9 163.367
R1357 B.n691 B.n11 163.367
R1358 B.n687 B.n11 163.367
R1359 B.n687 B.n17 163.367
R1360 B.n683 B.n17 163.367
R1361 B.n683 B.n19 163.367
R1362 B.n679 B.n19 163.367
R1363 B.n679 B.n24 163.367
R1364 B.n675 B.n24 163.367
R1365 B.n675 B.n26 163.367
R1366 B.n90 B.n29 71.676
R1367 B.n94 B.n30 71.676
R1368 B.n98 B.n31 71.676
R1369 B.n102 B.n32 71.676
R1370 B.n106 B.n33 71.676
R1371 B.n110 B.n34 71.676
R1372 B.n114 B.n35 71.676
R1373 B.n118 B.n36 71.676
R1374 B.n122 B.n37 71.676
R1375 B.n126 B.n38 71.676
R1376 B.n130 B.n39 71.676
R1377 B.n134 B.n40 71.676
R1378 B.n138 B.n41 71.676
R1379 B.n142 B.n42 71.676
R1380 B.n146 B.n43 71.676
R1381 B.n150 B.n44 71.676
R1382 B.n154 B.n45 71.676
R1383 B.n158 B.n46 71.676
R1384 B.n162 B.n47 71.676
R1385 B.n166 B.n48 71.676
R1386 B.n170 B.n49 71.676
R1387 B.n174 B.n50 71.676
R1388 B.n178 B.n51 71.676
R1389 B.n182 B.n52 71.676
R1390 B.n186 B.n53 71.676
R1391 B.n190 B.n54 71.676
R1392 B.n194 B.n55 71.676
R1393 B.n198 B.n56 71.676
R1394 B.n202 B.n57 71.676
R1395 B.n206 B.n58 71.676
R1396 B.n210 B.n59 71.676
R1397 B.n214 B.n60 71.676
R1398 B.n218 B.n61 71.676
R1399 B.n222 B.n62 71.676
R1400 B.n226 B.n63 71.676
R1401 B.n230 B.n64 71.676
R1402 B.n234 B.n65 71.676
R1403 B.n238 B.n66 71.676
R1404 B.n242 B.n67 71.676
R1405 B.n246 B.n68 71.676
R1406 B.n250 B.n69 71.676
R1407 B.n254 B.n70 71.676
R1408 B.n258 B.n71 71.676
R1409 B.n262 B.n72 71.676
R1410 B.n266 B.n73 71.676
R1411 B.n270 B.n74 71.676
R1412 B.n274 B.n75 71.676
R1413 B.n278 B.n76 71.676
R1414 B.n282 B.n77 71.676
R1415 B.n286 B.n78 71.676
R1416 B.n290 B.n79 71.676
R1417 B.n294 B.n80 71.676
R1418 B.n298 B.n81 71.676
R1419 B.n302 B.n82 71.676
R1420 B.n671 B.n83 71.676
R1421 B.n671 B.n670 71.676
R1422 B.n304 B.n82 71.676
R1423 B.n301 B.n81 71.676
R1424 B.n297 B.n80 71.676
R1425 B.n293 B.n79 71.676
R1426 B.n289 B.n78 71.676
R1427 B.n285 B.n77 71.676
R1428 B.n281 B.n76 71.676
R1429 B.n277 B.n75 71.676
R1430 B.n273 B.n74 71.676
R1431 B.n269 B.n73 71.676
R1432 B.n265 B.n72 71.676
R1433 B.n261 B.n71 71.676
R1434 B.n257 B.n70 71.676
R1435 B.n253 B.n69 71.676
R1436 B.n249 B.n68 71.676
R1437 B.n245 B.n67 71.676
R1438 B.n241 B.n66 71.676
R1439 B.n237 B.n65 71.676
R1440 B.n233 B.n64 71.676
R1441 B.n229 B.n63 71.676
R1442 B.n225 B.n62 71.676
R1443 B.n221 B.n61 71.676
R1444 B.n217 B.n60 71.676
R1445 B.n213 B.n59 71.676
R1446 B.n209 B.n58 71.676
R1447 B.n205 B.n57 71.676
R1448 B.n201 B.n56 71.676
R1449 B.n197 B.n55 71.676
R1450 B.n193 B.n54 71.676
R1451 B.n189 B.n53 71.676
R1452 B.n185 B.n52 71.676
R1453 B.n181 B.n51 71.676
R1454 B.n177 B.n50 71.676
R1455 B.n173 B.n49 71.676
R1456 B.n169 B.n48 71.676
R1457 B.n165 B.n47 71.676
R1458 B.n161 B.n46 71.676
R1459 B.n157 B.n45 71.676
R1460 B.n153 B.n44 71.676
R1461 B.n149 B.n43 71.676
R1462 B.n145 B.n42 71.676
R1463 B.n141 B.n41 71.676
R1464 B.n137 B.n40 71.676
R1465 B.n133 B.n39 71.676
R1466 B.n129 B.n38 71.676
R1467 B.n125 B.n37 71.676
R1468 B.n121 B.n36 71.676
R1469 B.n117 B.n35 71.676
R1470 B.n113 B.n34 71.676
R1471 B.n109 B.n33 71.676
R1472 B.n105 B.n32 71.676
R1473 B.n101 B.n31 71.676
R1474 B.n97 B.n30 71.676
R1475 B.n93 B.n29 71.676
R1476 B.n607 B.n606 71.676
R1477 B.n601 B.n332 71.676
R1478 B.n598 B.n333 71.676
R1479 B.n594 B.n334 71.676
R1480 B.n590 B.n335 71.676
R1481 B.n586 B.n336 71.676
R1482 B.n582 B.n337 71.676
R1483 B.n578 B.n338 71.676
R1484 B.n574 B.n339 71.676
R1485 B.n570 B.n340 71.676
R1486 B.n566 B.n341 71.676
R1487 B.n562 B.n342 71.676
R1488 B.n558 B.n343 71.676
R1489 B.n554 B.n344 71.676
R1490 B.n550 B.n345 71.676
R1491 B.n546 B.n346 71.676
R1492 B.n542 B.n347 71.676
R1493 B.n538 B.n348 71.676
R1494 B.n534 B.n349 71.676
R1495 B.n530 B.n350 71.676
R1496 B.n526 B.n351 71.676
R1497 B.n522 B.n352 71.676
R1498 B.n518 B.n353 71.676
R1499 B.n514 B.n354 71.676
R1500 B.n510 B.n355 71.676
R1501 B.n505 B.n356 71.676
R1502 B.n501 B.n357 71.676
R1503 B.n497 B.n358 71.676
R1504 B.n493 B.n359 71.676
R1505 B.n489 B.n360 71.676
R1506 B.n484 B.n361 71.676
R1507 B.n480 B.n362 71.676
R1508 B.n476 B.n363 71.676
R1509 B.n472 B.n364 71.676
R1510 B.n468 B.n365 71.676
R1511 B.n464 B.n366 71.676
R1512 B.n460 B.n367 71.676
R1513 B.n456 B.n368 71.676
R1514 B.n452 B.n369 71.676
R1515 B.n448 B.n370 71.676
R1516 B.n444 B.n371 71.676
R1517 B.n440 B.n372 71.676
R1518 B.n436 B.n373 71.676
R1519 B.n432 B.n374 71.676
R1520 B.n428 B.n375 71.676
R1521 B.n424 B.n376 71.676
R1522 B.n420 B.n377 71.676
R1523 B.n416 B.n378 71.676
R1524 B.n412 B.n379 71.676
R1525 B.n408 B.n380 71.676
R1526 B.n404 B.n381 71.676
R1527 B.n400 B.n382 71.676
R1528 B.n396 B.n383 71.676
R1529 B.n392 B.n384 71.676
R1530 B.n607 B.n386 71.676
R1531 B.n599 B.n332 71.676
R1532 B.n595 B.n333 71.676
R1533 B.n591 B.n334 71.676
R1534 B.n587 B.n335 71.676
R1535 B.n583 B.n336 71.676
R1536 B.n579 B.n337 71.676
R1537 B.n575 B.n338 71.676
R1538 B.n571 B.n339 71.676
R1539 B.n567 B.n340 71.676
R1540 B.n563 B.n341 71.676
R1541 B.n559 B.n342 71.676
R1542 B.n555 B.n343 71.676
R1543 B.n551 B.n344 71.676
R1544 B.n547 B.n345 71.676
R1545 B.n543 B.n346 71.676
R1546 B.n539 B.n347 71.676
R1547 B.n535 B.n348 71.676
R1548 B.n531 B.n349 71.676
R1549 B.n527 B.n350 71.676
R1550 B.n523 B.n351 71.676
R1551 B.n519 B.n352 71.676
R1552 B.n515 B.n353 71.676
R1553 B.n511 B.n354 71.676
R1554 B.n506 B.n355 71.676
R1555 B.n502 B.n356 71.676
R1556 B.n498 B.n357 71.676
R1557 B.n494 B.n358 71.676
R1558 B.n490 B.n359 71.676
R1559 B.n485 B.n360 71.676
R1560 B.n481 B.n361 71.676
R1561 B.n477 B.n362 71.676
R1562 B.n473 B.n363 71.676
R1563 B.n469 B.n364 71.676
R1564 B.n465 B.n365 71.676
R1565 B.n461 B.n366 71.676
R1566 B.n457 B.n367 71.676
R1567 B.n453 B.n368 71.676
R1568 B.n449 B.n369 71.676
R1569 B.n445 B.n370 71.676
R1570 B.n441 B.n371 71.676
R1571 B.n437 B.n372 71.676
R1572 B.n433 B.n373 71.676
R1573 B.n429 B.n374 71.676
R1574 B.n425 B.n375 71.676
R1575 B.n421 B.n376 71.676
R1576 B.n417 B.n377 71.676
R1577 B.n413 B.n378 71.676
R1578 B.n409 B.n379 71.676
R1579 B.n405 B.n380 71.676
R1580 B.n401 B.n381 71.676
R1581 B.n397 B.n382 71.676
R1582 B.n393 B.n383 71.676
R1583 B.n384 B.n331 71.676
R1584 B.n701 B.n700 71.676
R1585 B.n701 B.n2 71.676
R1586 B.n608 B.n328 68.188
R1587 B.n673 B.n672 68.188
R1588 B.n89 B.n88 59.5399
R1589 B.n86 B.n85 59.5399
R1590 B.n487 B.n390 59.5399
R1591 B.n508 B.n388 59.5399
R1592 B.n614 B.n328 37.0945
R1593 B.n614 B.n323 37.0945
R1594 B.n620 B.n323 37.0945
R1595 B.n620 B.n324 37.0945
R1596 B.n626 B.n316 37.0945
R1597 B.n632 B.n316 37.0945
R1598 B.n632 B.n312 37.0945
R1599 B.n640 B.n312 37.0945
R1600 B.n640 B.n639 37.0945
R1601 B.n646 B.n4 37.0945
R1602 B.n699 B.n4 37.0945
R1603 B.n699 B.n698 37.0945
R1604 B.n698 B.n697 37.0945
R1605 B.n697 B.n8 37.0945
R1606 B.n690 B.n12 37.0945
R1607 B.n690 B.n689 37.0945
R1608 B.n689 B.n688 37.0945
R1609 B.n688 B.n16 37.0945
R1610 B.n682 B.n16 37.0945
R1611 B.n681 B.n680 37.0945
R1612 B.n680 B.n23 37.0945
R1613 B.n674 B.n23 37.0945
R1614 B.n674 B.n673 37.0945
R1615 B.n605 B.n326 31.6883
R1616 B.n611 B.n610 31.6883
R1617 B.n669 B.n668 31.6883
R1618 B.n91 B.n25 31.6883
R1619 B.n324 B.t10 23.457
R1620 B.t3 B.n681 23.457
R1621 B.n639 B.t1 20.184
R1622 B.n12 B.t0 20.184
R1623 B B.n702 18.0485
R1624 B.n88 B.n87 17.8429
R1625 B.n85 B.n84 17.8429
R1626 B.n390 B.n389 17.8429
R1627 B.n388 B.n387 17.8429
R1628 B.n646 B.t1 16.911
R1629 B.t0 B.n8 16.911
R1630 B.n626 B.t10 13.638
R1631 B.n682 B.t3 13.638
R1632 B.n616 B.n326 10.6151
R1633 B.n617 B.n616 10.6151
R1634 B.n618 B.n617 10.6151
R1635 B.n618 B.n318 10.6151
R1636 B.n628 B.n318 10.6151
R1637 B.n629 B.n628 10.6151
R1638 B.n630 B.n629 10.6151
R1639 B.n630 B.n310 10.6151
R1640 B.n642 B.n310 10.6151
R1641 B.n643 B.n642 10.6151
R1642 B.n644 B.n643 10.6151
R1643 B.n644 B.n0 10.6151
R1644 B.n605 B.n604 10.6151
R1645 B.n604 B.n603 10.6151
R1646 B.n603 B.n602 10.6151
R1647 B.n602 B.n600 10.6151
R1648 B.n600 B.n597 10.6151
R1649 B.n597 B.n596 10.6151
R1650 B.n596 B.n593 10.6151
R1651 B.n593 B.n592 10.6151
R1652 B.n592 B.n589 10.6151
R1653 B.n589 B.n588 10.6151
R1654 B.n588 B.n585 10.6151
R1655 B.n585 B.n584 10.6151
R1656 B.n584 B.n581 10.6151
R1657 B.n581 B.n580 10.6151
R1658 B.n580 B.n577 10.6151
R1659 B.n577 B.n576 10.6151
R1660 B.n576 B.n573 10.6151
R1661 B.n573 B.n572 10.6151
R1662 B.n572 B.n569 10.6151
R1663 B.n569 B.n568 10.6151
R1664 B.n568 B.n565 10.6151
R1665 B.n565 B.n564 10.6151
R1666 B.n564 B.n561 10.6151
R1667 B.n561 B.n560 10.6151
R1668 B.n560 B.n557 10.6151
R1669 B.n557 B.n556 10.6151
R1670 B.n556 B.n553 10.6151
R1671 B.n553 B.n552 10.6151
R1672 B.n552 B.n549 10.6151
R1673 B.n549 B.n548 10.6151
R1674 B.n548 B.n545 10.6151
R1675 B.n545 B.n544 10.6151
R1676 B.n544 B.n541 10.6151
R1677 B.n541 B.n540 10.6151
R1678 B.n540 B.n537 10.6151
R1679 B.n537 B.n536 10.6151
R1680 B.n536 B.n533 10.6151
R1681 B.n533 B.n532 10.6151
R1682 B.n532 B.n529 10.6151
R1683 B.n529 B.n528 10.6151
R1684 B.n528 B.n525 10.6151
R1685 B.n525 B.n524 10.6151
R1686 B.n524 B.n521 10.6151
R1687 B.n521 B.n520 10.6151
R1688 B.n520 B.n517 10.6151
R1689 B.n517 B.n516 10.6151
R1690 B.n516 B.n513 10.6151
R1691 B.n513 B.n512 10.6151
R1692 B.n512 B.n509 10.6151
R1693 B.n507 B.n504 10.6151
R1694 B.n504 B.n503 10.6151
R1695 B.n503 B.n500 10.6151
R1696 B.n500 B.n499 10.6151
R1697 B.n499 B.n496 10.6151
R1698 B.n496 B.n495 10.6151
R1699 B.n495 B.n492 10.6151
R1700 B.n492 B.n491 10.6151
R1701 B.n491 B.n488 10.6151
R1702 B.n486 B.n483 10.6151
R1703 B.n483 B.n482 10.6151
R1704 B.n482 B.n479 10.6151
R1705 B.n479 B.n478 10.6151
R1706 B.n478 B.n475 10.6151
R1707 B.n475 B.n474 10.6151
R1708 B.n474 B.n471 10.6151
R1709 B.n471 B.n470 10.6151
R1710 B.n470 B.n467 10.6151
R1711 B.n467 B.n466 10.6151
R1712 B.n466 B.n463 10.6151
R1713 B.n463 B.n462 10.6151
R1714 B.n462 B.n459 10.6151
R1715 B.n459 B.n458 10.6151
R1716 B.n458 B.n455 10.6151
R1717 B.n455 B.n454 10.6151
R1718 B.n454 B.n451 10.6151
R1719 B.n451 B.n450 10.6151
R1720 B.n450 B.n447 10.6151
R1721 B.n447 B.n446 10.6151
R1722 B.n446 B.n443 10.6151
R1723 B.n443 B.n442 10.6151
R1724 B.n442 B.n439 10.6151
R1725 B.n439 B.n438 10.6151
R1726 B.n438 B.n435 10.6151
R1727 B.n435 B.n434 10.6151
R1728 B.n434 B.n431 10.6151
R1729 B.n431 B.n430 10.6151
R1730 B.n430 B.n427 10.6151
R1731 B.n427 B.n426 10.6151
R1732 B.n426 B.n423 10.6151
R1733 B.n423 B.n422 10.6151
R1734 B.n422 B.n419 10.6151
R1735 B.n419 B.n418 10.6151
R1736 B.n418 B.n415 10.6151
R1737 B.n415 B.n414 10.6151
R1738 B.n414 B.n411 10.6151
R1739 B.n411 B.n410 10.6151
R1740 B.n410 B.n407 10.6151
R1741 B.n407 B.n406 10.6151
R1742 B.n406 B.n403 10.6151
R1743 B.n403 B.n402 10.6151
R1744 B.n402 B.n399 10.6151
R1745 B.n399 B.n398 10.6151
R1746 B.n398 B.n395 10.6151
R1747 B.n395 B.n394 10.6151
R1748 B.n394 B.n391 10.6151
R1749 B.n391 B.n330 10.6151
R1750 B.n610 B.n330 10.6151
R1751 B.n612 B.n611 10.6151
R1752 B.n612 B.n321 10.6151
R1753 B.n622 B.n321 10.6151
R1754 B.n623 B.n622 10.6151
R1755 B.n624 B.n623 10.6151
R1756 B.n624 B.n314 10.6151
R1757 B.n634 B.n314 10.6151
R1758 B.n635 B.n634 10.6151
R1759 B.n637 B.n635 10.6151
R1760 B.n637 B.n636 10.6151
R1761 B.n636 B.n307 10.6151
R1762 B.n649 B.n307 10.6151
R1763 B.n650 B.n649 10.6151
R1764 B.n651 B.n650 10.6151
R1765 B.n652 B.n651 10.6151
R1766 B.n653 B.n652 10.6151
R1767 B.n656 B.n653 10.6151
R1768 B.n657 B.n656 10.6151
R1769 B.n658 B.n657 10.6151
R1770 B.n659 B.n658 10.6151
R1771 B.n661 B.n659 10.6151
R1772 B.n662 B.n661 10.6151
R1773 B.n663 B.n662 10.6151
R1774 B.n664 B.n663 10.6151
R1775 B.n666 B.n664 10.6151
R1776 B.n667 B.n666 10.6151
R1777 B.n668 B.n667 10.6151
R1778 B.n694 B.n1 10.6151
R1779 B.n694 B.n693 10.6151
R1780 B.n693 B.n692 10.6151
R1781 B.n692 B.n10 10.6151
R1782 B.n686 B.n10 10.6151
R1783 B.n686 B.n685 10.6151
R1784 B.n685 B.n684 10.6151
R1785 B.n684 B.n18 10.6151
R1786 B.n678 B.n18 10.6151
R1787 B.n678 B.n677 10.6151
R1788 B.n677 B.n676 10.6151
R1789 B.n676 B.n25 10.6151
R1790 B.n92 B.n91 10.6151
R1791 B.n95 B.n92 10.6151
R1792 B.n96 B.n95 10.6151
R1793 B.n99 B.n96 10.6151
R1794 B.n100 B.n99 10.6151
R1795 B.n103 B.n100 10.6151
R1796 B.n104 B.n103 10.6151
R1797 B.n107 B.n104 10.6151
R1798 B.n108 B.n107 10.6151
R1799 B.n111 B.n108 10.6151
R1800 B.n112 B.n111 10.6151
R1801 B.n115 B.n112 10.6151
R1802 B.n116 B.n115 10.6151
R1803 B.n119 B.n116 10.6151
R1804 B.n120 B.n119 10.6151
R1805 B.n123 B.n120 10.6151
R1806 B.n124 B.n123 10.6151
R1807 B.n127 B.n124 10.6151
R1808 B.n128 B.n127 10.6151
R1809 B.n131 B.n128 10.6151
R1810 B.n132 B.n131 10.6151
R1811 B.n135 B.n132 10.6151
R1812 B.n136 B.n135 10.6151
R1813 B.n139 B.n136 10.6151
R1814 B.n140 B.n139 10.6151
R1815 B.n143 B.n140 10.6151
R1816 B.n144 B.n143 10.6151
R1817 B.n147 B.n144 10.6151
R1818 B.n148 B.n147 10.6151
R1819 B.n151 B.n148 10.6151
R1820 B.n152 B.n151 10.6151
R1821 B.n155 B.n152 10.6151
R1822 B.n156 B.n155 10.6151
R1823 B.n159 B.n156 10.6151
R1824 B.n160 B.n159 10.6151
R1825 B.n163 B.n160 10.6151
R1826 B.n164 B.n163 10.6151
R1827 B.n167 B.n164 10.6151
R1828 B.n168 B.n167 10.6151
R1829 B.n171 B.n168 10.6151
R1830 B.n172 B.n171 10.6151
R1831 B.n175 B.n172 10.6151
R1832 B.n176 B.n175 10.6151
R1833 B.n179 B.n176 10.6151
R1834 B.n180 B.n179 10.6151
R1835 B.n183 B.n180 10.6151
R1836 B.n184 B.n183 10.6151
R1837 B.n187 B.n184 10.6151
R1838 B.n188 B.n187 10.6151
R1839 B.n192 B.n191 10.6151
R1840 B.n195 B.n192 10.6151
R1841 B.n196 B.n195 10.6151
R1842 B.n199 B.n196 10.6151
R1843 B.n200 B.n199 10.6151
R1844 B.n203 B.n200 10.6151
R1845 B.n204 B.n203 10.6151
R1846 B.n207 B.n204 10.6151
R1847 B.n208 B.n207 10.6151
R1848 B.n212 B.n211 10.6151
R1849 B.n215 B.n212 10.6151
R1850 B.n216 B.n215 10.6151
R1851 B.n219 B.n216 10.6151
R1852 B.n220 B.n219 10.6151
R1853 B.n223 B.n220 10.6151
R1854 B.n224 B.n223 10.6151
R1855 B.n227 B.n224 10.6151
R1856 B.n228 B.n227 10.6151
R1857 B.n231 B.n228 10.6151
R1858 B.n232 B.n231 10.6151
R1859 B.n235 B.n232 10.6151
R1860 B.n236 B.n235 10.6151
R1861 B.n239 B.n236 10.6151
R1862 B.n240 B.n239 10.6151
R1863 B.n243 B.n240 10.6151
R1864 B.n244 B.n243 10.6151
R1865 B.n247 B.n244 10.6151
R1866 B.n248 B.n247 10.6151
R1867 B.n251 B.n248 10.6151
R1868 B.n252 B.n251 10.6151
R1869 B.n255 B.n252 10.6151
R1870 B.n256 B.n255 10.6151
R1871 B.n259 B.n256 10.6151
R1872 B.n260 B.n259 10.6151
R1873 B.n263 B.n260 10.6151
R1874 B.n264 B.n263 10.6151
R1875 B.n267 B.n264 10.6151
R1876 B.n268 B.n267 10.6151
R1877 B.n271 B.n268 10.6151
R1878 B.n272 B.n271 10.6151
R1879 B.n275 B.n272 10.6151
R1880 B.n276 B.n275 10.6151
R1881 B.n279 B.n276 10.6151
R1882 B.n280 B.n279 10.6151
R1883 B.n283 B.n280 10.6151
R1884 B.n284 B.n283 10.6151
R1885 B.n287 B.n284 10.6151
R1886 B.n288 B.n287 10.6151
R1887 B.n291 B.n288 10.6151
R1888 B.n292 B.n291 10.6151
R1889 B.n295 B.n292 10.6151
R1890 B.n296 B.n295 10.6151
R1891 B.n299 B.n296 10.6151
R1892 B.n300 B.n299 10.6151
R1893 B.n303 B.n300 10.6151
R1894 B.n305 B.n303 10.6151
R1895 B.n306 B.n305 10.6151
R1896 B.n669 B.n306 10.6151
R1897 B.n509 B.n508 8.74196
R1898 B.n487 B.n486 8.74196
R1899 B.n188 B.n89 8.74196
R1900 B.n211 B.n86 8.74196
R1901 B.n702 B.n0 8.11757
R1902 B.n702 B.n1 8.11757
R1903 B.n508 B.n507 1.87367
R1904 B.n488 B.n487 1.87367
R1905 B.n191 B.n89 1.87367
R1906 B.n208 B.n86 1.87367
R1907 VP.n0 VP.t0 877.207
R1908 VP.n0 VP.t1 835.692
R1909 VP VP.n0 0.0516364
R1910 VDD1.n76 VDD1.n0 289.615
R1911 VDD1.n157 VDD1.n81 289.615
R1912 VDD1.n77 VDD1.n76 185
R1913 VDD1.n75 VDD1.n74 185
R1914 VDD1.n73 VDD1.n3 185
R1915 VDD1.n7 VDD1.n4 185
R1916 VDD1.n68 VDD1.n67 185
R1917 VDD1.n66 VDD1.n65 185
R1918 VDD1.n9 VDD1.n8 185
R1919 VDD1.n60 VDD1.n59 185
R1920 VDD1.n58 VDD1.n57 185
R1921 VDD1.n13 VDD1.n12 185
R1922 VDD1.n52 VDD1.n51 185
R1923 VDD1.n50 VDD1.n49 185
R1924 VDD1.n17 VDD1.n16 185
R1925 VDD1.n44 VDD1.n43 185
R1926 VDD1.n42 VDD1.n41 185
R1927 VDD1.n21 VDD1.n20 185
R1928 VDD1.n36 VDD1.n35 185
R1929 VDD1.n34 VDD1.n33 185
R1930 VDD1.n25 VDD1.n24 185
R1931 VDD1.n28 VDD1.n27 185
R1932 VDD1.n108 VDD1.n107 185
R1933 VDD1.n105 VDD1.n104 185
R1934 VDD1.n114 VDD1.n113 185
R1935 VDD1.n116 VDD1.n115 185
R1936 VDD1.n101 VDD1.n100 185
R1937 VDD1.n122 VDD1.n121 185
R1938 VDD1.n124 VDD1.n123 185
R1939 VDD1.n97 VDD1.n96 185
R1940 VDD1.n130 VDD1.n129 185
R1941 VDD1.n132 VDD1.n131 185
R1942 VDD1.n93 VDD1.n92 185
R1943 VDD1.n138 VDD1.n137 185
R1944 VDD1.n140 VDD1.n139 185
R1945 VDD1.n89 VDD1.n88 185
R1946 VDD1.n146 VDD1.n145 185
R1947 VDD1.n149 VDD1.n148 185
R1948 VDD1.n147 VDD1.n85 185
R1949 VDD1.n154 VDD1.n84 185
R1950 VDD1.n156 VDD1.n155 185
R1951 VDD1.n158 VDD1.n157 185
R1952 VDD1.t1 VDD1.n26 147.659
R1953 VDD1.t0 VDD1.n106 147.659
R1954 VDD1.n76 VDD1.n75 104.615
R1955 VDD1.n75 VDD1.n3 104.615
R1956 VDD1.n7 VDD1.n3 104.615
R1957 VDD1.n67 VDD1.n7 104.615
R1958 VDD1.n67 VDD1.n66 104.615
R1959 VDD1.n66 VDD1.n8 104.615
R1960 VDD1.n59 VDD1.n8 104.615
R1961 VDD1.n59 VDD1.n58 104.615
R1962 VDD1.n58 VDD1.n12 104.615
R1963 VDD1.n51 VDD1.n12 104.615
R1964 VDD1.n51 VDD1.n50 104.615
R1965 VDD1.n50 VDD1.n16 104.615
R1966 VDD1.n43 VDD1.n16 104.615
R1967 VDD1.n43 VDD1.n42 104.615
R1968 VDD1.n42 VDD1.n20 104.615
R1969 VDD1.n35 VDD1.n20 104.615
R1970 VDD1.n35 VDD1.n34 104.615
R1971 VDD1.n34 VDD1.n24 104.615
R1972 VDD1.n27 VDD1.n24 104.615
R1973 VDD1.n107 VDD1.n104 104.615
R1974 VDD1.n114 VDD1.n104 104.615
R1975 VDD1.n115 VDD1.n114 104.615
R1976 VDD1.n115 VDD1.n100 104.615
R1977 VDD1.n122 VDD1.n100 104.615
R1978 VDD1.n123 VDD1.n122 104.615
R1979 VDD1.n123 VDD1.n96 104.615
R1980 VDD1.n130 VDD1.n96 104.615
R1981 VDD1.n131 VDD1.n130 104.615
R1982 VDD1.n131 VDD1.n92 104.615
R1983 VDD1.n138 VDD1.n92 104.615
R1984 VDD1.n139 VDD1.n138 104.615
R1985 VDD1.n139 VDD1.n88 104.615
R1986 VDD1.n146 VDD1.n88 104.615
R1987 VDD1.n148 VDD1.n146 104.615
R1988 VDD1.n148 VDD1.n147 104.615
R1989 VDD1.n147 VDD1.n84 104.615
R1990 VDD1.n156 VDD1.n84 104.615
R1991 VDD1.n157 VDD1.n156 104.615
R1992 VDD1 VDD1.n161 92.1297
R1993 VDD1 VDD1.n80 53.5812
R1994 VDD1.n27 VDD1.t1 52.3082
R1995 VDD1.n107 VDD1.t0 52.3082
R1996 VDD1.n28 VDD1.n26 15.6677
R1997 VDD1.n108 VDD1.n106 15.6677
R1998 VDD1.n74 VDD1.n73 13.1884
R1999 VDD1.n155 VDD1.n154 13.1884
R2000 VDD1.n77 VDD1.n2 12.8005
R2001 VDD1.n72 VDD1.n4 12.8005
R2002 VDD1.n29 VDD1.n25 12.8005
R2003 VDD1.n109 VDD1.n105 12.8005
R2004 VDD1.n153 VDD1.n85 12.8005
R2005 VDD1.n158 VDD1.n83 12.8005
R2006 VDD1.n78 VDD1.n0 12.0247
R2007 VDD1.n69 VDD1.n68 12.0247
R2008 VDD1.n33 VDD1.n32 12.0247
R2009 VDD1.n113 VDD1.n112 12.0247
R2010 VDD1.n150 VDD1.n149 12.0247
R2011 VDD1.n159 VDD1.n81 12.0247
R2012 VDD1.n65 VDD1.n6 11.249
R2013 VDD1.n36 VDD1.n23 11.249
R2014 VDD1.n116 VDD1.n103 11.249
R2015 VDD1.n145 VDD1.n87 11.249
R2016 VDD1.n64 VDD1.n9 10.4732
R2017 VDD1.n37 VDD1.n21 10.4732
R2018 VDD1.n117 VDD1.n101 10.4732
R2019 VDD1.n144 VDD1.n89 10.4732
R2020 VDD1.n61 VDD1.n60 9.69747
R2021 VDD1.n41 VDD1.n40 9.69747
R2022 VDD1.n121 VDD1.n120 9.69747
R2023 VDD1.n141 VDD1.n140 9.69747
R2024 VDD1.n80 VDD1.n79 9.45567
R2025 VDD1.n161 VDD1.n160 9.45567
R2026 VDD1.n54 VDD1.n53 9.3005
R2027 VDD1.n56 VDD1.n55 9.3005
R2028 VDD1.n11 VDD1.n10 9.3005
R2029 VDD1.n62 VDD1.n61 9.3005
R2030 VDD1.n64 VDD1.n63 9.3005
R2031 VDD1.n6 VDD1.n5 9.3005
R2032 VDD1.n70 VDD1.n69 9.3005
R2033 VDD1.n72 VDD1.n71 9.3005
R2034 VDD1.n79 VDD1.n78 9.3005
R2035 VDD1.n2 VDD1.n1 9.3005
R2036 VDD1.n15 VDD1.n14 9.3005
R2037 VDD1.n48 VDD1.n47 9.3005
R2038 VDD1.n46 VDD1.n45 9.3005
R2039 VDD1.n19 VDD1.n18 9.3005
R2040 VDD1.n40 VDD1.n39 9.3005
R2041 VDD1.n38 VDD1.n37 9.3005
R2042 VDD1.n23 VDD1.n22 9.3005
R2043 VDD1.n32 VDD1.n31 9.3005
R2044 VDD1.n30 VDD1.n29 9.3005
R2045 VDD1.n160 VDD1.n159 9.3005
R2046 VDD1.n83 VDD1.n82 9.3005
R2047 VDD1.n128 VDD1.n127 9.3005
R2048 VDD1.n126 VDD1.n125 9.3005
R2049 VDD1.n99 VDD1.n98 9.3005
R2050 VDD1.n120 VDD1.n119 9.3005
R2051 VDD1.n118 VDD1.n117 9.3005
R2052 VDD1.n103 VDD1.n102 9.3005
R2053 VDD1.n112 VDD1.n111 9.3005
R2054 VDD1.n110 VDD1.n109 9.3005
R2055 VDD1.n95 VDD1.n94 9.3005
R2056 VDD1.n134 VDD1.n133 9.3005
R2057 VDD1.n136 VDD1.n135 9.3005
R2058 VDD1.n91 VDD1.n90 9.3005
R2059 VDD1.n142 VDD1.n141 9.3005
R2060 VDD1.n144 VDD1.n143 9.3005
R2061 VDD1.n87 VDD1.n86 9.3005
R2062 VDD1.n151 VDD1.n150 9.3005
R2063 VDD1.n153 VDD1.n152 9.3005
R2064 VDD1.n57 VDD1.n11 8.92171
R2065 VDD1.n44 VDD1.n19 8.92171
R2066 VDD1.n124 VDD1.n99 8.92171
R2067 VDD1.n137 VDD1.n91 8.92171
R2068 VDD1.n56 VDD1.n13 8.14595
R2069 VDD1.n45 VDD1.n17 8.14595
R2070 VDD1.n125 VDD1.n97 8.14595
R2071 VDD1.n136 VDD1.n93 8.14595
R2072 VDD1.n53 VDD1.n52 7.3702
R2073 VDD1.n49 VDD1.n48 7.3702
R2074 VDD1.n129 VDD1.n128 7.3702
R2075 VDD1.n133 VDD1.n132 7.3702
R2076 VDD1.n52 VDD1.n15 6.59444
R2077 VDD1.n49 VDD1.n15 6.59444
R2078 VDD1.n129 VDD1.n95 6.59444
R2079 VDD1.n132 VDD1.n95 6.59444
R2080 VDD1.n53 VDD1.n13 5.81868
R2081 VDD1.n48 VDD1.n17 5.81868
R2082 VDD1.n128 VDD1.n97 5.81868
R2083 VDD1.n133 VDD1.n93 5.81868
R2084 VDD1.n57 VDD1.n56 5.04292
R2085 VDD1.n45 VDD1.n44 5.04292
R2086 VDD1.n125 VDD1.n124 5.04292
R2087 VDD1.n137 VDD1.n136 5.04292
R2088 VDD1.n30 VDD1.n26 4.38563
R2089 VDD1.n110 VDD1.n106 4.38563
R2090 VDD1.n60 VDD1.n11 4.26717
R2091 VDD1.n41 VDD1.n19 4.26717
R2092 VDD1.n121 VDD1.n99 4.26717
R2093 VDD1.n140 VDD1.n91 4.26717
R2094 VDD1.n61 VDD1.n9 3.49141
R2095 VDD1.n40 VDD1.n21 3.49141
R2096 VDD1.n120 VDD1.n101 3.49141
R2097 VDD1.n141 VDD1.n89 3.49141
R2098 VDD1.n65 VDD1.n64 2.71565
R2099 VDD1.n37 VDD1.n36 2.71565
R2100 VDD1.n117 VDD1.n116 2.71565
R2101 VDD1.n145 VDD1.n144 2.71565
R2102 VDD1.n80 VDD1.n0 1.93989
R2103 VDD1.n68 VDD1.n6 1.93989
R2104 VDD1.n33 VDD1.n23 1.93989
R2105 VDD1.n113 VDD1.n103 1.93989
R2106 VDD1.n149 VDD1.n87 1.93989
R2107 VDD1.n161 VDD1.n81 1.93989
R2108 VDD1.n78 VDD1.n77 1.16414
R2109 VDD1.n69 VDD1.n4 1.16414
R2110 VDD1.n32 VDD1.n25 1.16414
R2111 VDD1.n112 VDD1.n105 1.16414
R2112 VDD1.n150 VDD1.n85 1.16414
R2113 VDD1.n159 VDD1.n158 1.16414
R2114 VDD1.n74 VDD1.n2 0.388379
R2115 VDD1.n73 VDD1.n72 0.388379
R2116 VDD1.n29 VDD1.n28 0.388379
R2117 VDD1.n109 VDD1.n108 0.388379
R2118 VDD1.n154 VDD1.n153 0.388379
R2119 VDD1.n155 VDD1.n83 0.388379
R2120 VDD1.n79 VDD1.n1 0.155672
R2121 VDD1.n71 VDD1.n1 0.155672
R2122 VDD1.n71 VDD1.n70 0.155672
R2123 VDD1.n70 VDD1.n5 0.155672
R2124 VDD1.n63 VDD1.n5 0.155672
R2125 VDD1.n63 VDD1.n62 0.155672
R2126 VDD1.n62 VDD1.n10 0.155672
R2127 VDD1.n55 VDD1.n10 0.155672
R2128 VDD1.n55 VDD1.n54 0.155672
R2129 VDD1.n54 VDD1.n14 0.155672
R2130 VDD1.n47 VDD1.n14 0.155672
R2131 VDD1.n47 VDD1.n46 0.155672
R2132 VDD1.n46 VDD1.n18 0.155672
R2133 VDD1.n39 VDD1.n18 0.155672
R2134 VDD1.n39 VDD1.n38 0.155672
R2135 VDD1.n38 VDD1.n22 0.155672
R2136 VDD1.n31 VDD1.n22 0.155672
R2137 VDD1.n31 VDD1.n30 0.155672
R2138 VDD1.n111 VDD1.n110 0.155672
R2139 VDD1.n111 VDD1.n102 0.155672
R2140 VDD1.n118 VDD1.n102 0.155672
R2141 VDD1.n119 VDD1.n118 0.155672
R2142 VDD1.n119 VDD1.n98 0.155672
R2143 VDD1.n126 VDD1.n98 0.155672
R2144 VDD1.n127 VDD1.n126 0.155672
R2145 VDD1.n127 VDD1.n94 0.155672
R2146 VDD1.n134 VDD1.n94 0.155672
R2147 VDD1.n135 VDD1.n134 0.155672
R2148 VDD1.n135 VDD1.n90 0.155672
R2149 VDD1.n142 VDD1.n90 0.155672
R2150 VDD1.n143 VDD1.n142 0.155672
R2151 VDD1.n143 VDD1.n86 0.155672
R2152 VDD1.n151 VDD1.n86 0.155672
R2153 VDD1.n152 VDD1.n151 0.155672
R2154 VDD1.n152 VDD1.n82 0.155672
R2155 VDD1.n160 VDD1.n82 0.155672
C0 VDD2 VDD1 0.452653f
C1 VN VDD1 0.148539f
C2 VDD1 VP 2.35281f
C3 VDD1 VTAIL 6.98948f
C4 VDD2 VN 2.25603f
C5 VDD2 VP 0.250891f
C6 VDD2 VTAIL 7.02042f
C7 VN VP 5.0435f
C8 VN VTAIL 1.60042f
C9 VTAIL VP 1.61519f
C10 VDD2 B 4.232365f
C11 VDD1 B 6.973589f
C12 VTAIL B 7.42718f
C13 VN B 8.79451f
C14 VP B 4.092576f
C15 VDD1.n0 B 0.030462f
C16 VDD1.n1 B 0.021364f
C17 VDD1.n2 B 0.01148f
C18 VDD1.n3 B 0.027135f
C19 VDD1.n4 B 0.012156f
C20 VDD1.n5 B 0.021364f
C21 VDD1.n6 B 0.01148f
C22 VDD1.n7 B 0.027135f
C23 VDD1.n8 B 0.027135f
C24 VDD1.n9 B 0.012156f
C25 VDD1.n10 B 0.021364f
C26 VDD1.n11 B 0.01148f
C27 VDD1.n12 B 0.027135f
C28 VDD1.n13 B 0.012156f
C29 VDD1.n14 B 0.021364f
C30 VDD1.n15 B 0.01148f
C31 VDD1.n16 B 0.027135f
C32 VDD1.n17 B 0.012156f
C33 VDD1.n18 B 0.021364f
C34 VDD1.n19 B 0.01148f
C35 VDD1.n20 B 0.027135f
C36 VDD1.n21 B 0.012156f
C37 VDD1.n22 B 0.021364f
C38 VDD1.n23 B 0.01148f
C39 VDD1.n24 B 0.027135f
C40 VDD1.n25 B 0.012156f
C41 VDD1.n26 B 0.138646f
C42 VDD1.t1 B 0.044733f
C43 VDD1.n27 B 0.020351f
C44 VDD1.n28 B 0.016029f
C45 VDD1.n29 B 0.01148f
C46 VDD1.n30 B 1.37726f
C47 VDD1.n31 B 0.021364f
C48 VDD1.n32 B 0.01148f
C49 VDD1.n33 B 0.012156f
C50 VDD1.n34 B 0.027135f
C51 VDD1.n35 B 0.027135f
C52 VDD1.n36 B 0.012156f
C53 VDD1.n37 B 0.01148f
C54 VDD1.n38 B 0.021364f
C55 VDD1.n39 B 0.021364f
C56 VDD1.n40 B 0.01148f
C57 VDD1.n41 B 0.012156f
C58 VDD1.n42 B 0.027135f
C59 VDD1.n43 B 0.027135f
C60 VDD1.n44 B 0.012156f
C61 VDD1.n45 B 0.01148f
C62 VDD1.n46 B 0.021364f
C63 VDD1.n47 B 0.021364f
C64 VDD1.n48 B 0.01148f
C65 VDD1.n49 B 0.012156f
C66 VDD1.n50 B 0.027135f
C67 VDD1.n51 B 0.027135f
C68 VDD1.n52 B 0.012156f
C69 VDD1.n53 B 0.01148f
C70 VDD1.n54 B 0.021364f
C71 VDD1.n55 B 0.021364f
C72 VDD1.n56 B 0.01148f
C73 VDD1.n57 B 0.012156f
C74 VDD1.n58 B 0.027135f
C75 VDD1.n59 B 0.027135f
C76 VDD1.n60 B 0.012156f
C77 VDD1.n61 B 0.01148f
C78 VDD1.n62 B 0.021364f
C79 VDD1.n63 B 0.021364f
C80 VDD1.n64 B 0.01148f
C81 VDD1.n65 B 0.012156f
C82 VDD1.n66 B 0.027135f
C83 VDD1.n67 B 0.027135f
C84 VDD1.n68 B 0.012156f
C85 VDD1.n69 B 0.01148f
C86 VDD1.n70 B 0.021364f
C87 VDD1.n71 B 0.021364f
C88 VDD1.n72 B 0.01148f
C89 VDD1.n73 B 0.011818f
C90 VDD1.n74 B 0.011818f
C91 VDD1.n75 B 0.027135f
C92 VDD1.n76 B 0.059508f
C93 VDD1.n77 B 0.012156f
C94 VDD1.n78 B 0.01148f
C95 VDD1.n79 B 0.056095f
C96 VDD1.n80 B 0.048576f
C97 VDD1.n81 B 0.030462f
C98 VDD1.n82 B 0.021364f
C99 VDD1.n83 B 0.01148f
C100 VDD1.n84 B 0.027135f
C101 VDD1.n85 B 0.012156f
C102 VDD1.n86 B 0.021364f
C103 VDD1.n87 B 0.01148f
C104 VDD1.n88 B 0.027135f
C105 VDD1.n89 B 0.012156f
C106 VDD1.n90 B 0.021364f
C107 VDD1.n91 B 0.01148f
C108 VDD1.n92 B 0.027135f
C109 VDD1.n93 B 0.012156f
C110 VDD1.n94 B 0.021364f
C111 VDD1.n95 B 0.01148f
C112 VDD1.n96 B 0.027135f
C113 VDD1.n97 B 0.012156f
C114 VDD1.n98 B 0.021364f
C115 VDD1.n99 B 0.01148f
C116 VDD1.n100 B 0.027135f
C117 VDD1.n101 B 0.012156f
C118 VDD1.n102 B 0.021364f
C119 VDD1.n103 B 0.01148f
C120 VDD1.n104 B 0.027135f
C121 VDD1.n105 B 0.012156f
C122 VDD1.n106 B 0.138646f
C123 VDD1.t0 B 0.044733f
C124 VDD1.n107 B 0.020351f
C125 VDD1.n108 B 0.016029f
C126 VDD1.n109 B 0.01148f
C127 VDD1.n110 B 1.37726f
C128 VDD1.n111 B 0.021364f
C129 VDD1.n112 B 0.01148f
C130 VDD1.n113 B 0.012156f
C131 VDD1.n114 B 0.027135f
C132 VDD1.n115 B 0.027135f
C133 VDD1.n116 B 0.012156f
C134 VDD1.n117 B 0.01148f
C135 VDD1.n118 B 0.021364f
C136 VDD1.n119 B 0.021364f
C137 VDD1.n120 B 0.01148f
C138 VDD1.n121 B 0.012156f
C139 VDD1.n122 B 0.027135f
C140 VDD1.n123 B 0.027135f
C141 VDD1.n124 B 0.012156f
C142 VDD1.n125 B 0.01148f
C143 VDD1.n126 B 0.021364f
C144 VDD1.n127 B 0.021364f
C145 VDD1.n128 B 0.01148f
C146 VDD1.n129 B 0.012156f
C147 VDD1.n130 B 0.027135f
C148 VDD1.n131 B 0.027135f
C149 VDD1.n132 B 0.012156f
C150 VDD1.n133 B 0.01148f
C151 VDD1.n134 B 0.021364f
C152 VDD1.n135 B 0.021364f
C153 VDD1.n136 B 0.01148f
C154 VDD1.n137 B 0.012156f
C155 VDD1.n138 B 0.027135f
C156 VDD1.n139 B 0.027135f
C157 VDD1.n140 B 0.012156f
C158 VDD1.n141 B 0.01148f
C159 VDD1.n142 B 0.021364f
C160 VDD1.n143 B 0.021364f
C161 VDD1.n144 B 0.01148f
C162 VDD1.n145 B 0.012156f
C163 VDD1.n146 B 0.027135f
C164 VDD1.n147 B 0.027135f
C165 VDD1.n148 B 0.027135f
C166 VDD1.n149 B 0.012156f
C167 VDD1.n150 B 0.01148f
C168 VDD1.n151 B 0.021364f
C169 VDD1.n152 B 0.021364f
C170 VDD1.n153 B 0.01148f
C171 VDD1.n154 B 0.011818f
C172 VDD1.n155 B 0.011818f
C173 VDD1.n156 B 0.027135f
C174 VDD1.n157 B 0.059508f
C175 VDD1.n158 B 0.012156f
C176 VDD1.n159 B 0.01148f
C177 VDD1.n160 B 0.056095f
C178 VDD1.n161 B 0.606247f
C179 VP.t0 B 1.42563f
C180 VP.t1 B 1.31371f
C181 VP.n0 B 4.6469f
C182 VDD2.n0 B 0.030393f
C183 VDD2.n1 B 0.021316f
C184 VDD2.n2 B 0.011454f
C185 VDD2.n3 B 0.027074f
C186 VDD2.n4 B 0.012128f
C187 VDD2.n5 B 0.021316f
C188 VDD2.n6 B 0.011454f
C189 VDD2.n7 B 0.027074f
C190 VDD2.n8 B 0.012128f
C191 VDD2.n9 B 0.021316f
C192 VDD2.n10 B 0.011454f
C193 VDD2.n11 B 0.027074f
C194 VDD2.n12 B 0.012128f
C195 VDD2.n13 B 0.021316f
C196 VDD2.n14 B 0.011454f
C197 VDD2.n15 B 0.027074f
C198 VDD2.n16 B 0.012128f
C199 VDD2.n17 B 0.021316f
C200 VDD2.n18 B 0.011454f
C201 VDD2.n19 B 0.027074f
C202 VDD2.n20 B 0.012128f
C203 VDD2.n21 B 0.021316f
C204 VDD2.n22 B 0.011454f
C205 VDD2.n23 B 0.027074f
C206 VDD2.n24 B 0.012128f
C207 VDD2.n25 B 0.138332f
C208 VDD2.t0 B 0.044632f
C209 VDD2.n26 B 0.020305f
C210 VDD2.n27 B 0.015993f
C211 VDD2.n28 B 0.011454f
C212 VDD2.n29 B 1.37414f
C213 VDD2.n30 B 0.021316f
C214 VDD2.n31 B 0.011454f
C215 VDD2.n32 B 0.012128f
C216 VDD2.n33 B 0.027074f
C217 VDD2.n34 B 0.027074f
C218 VDD2.n35 B 0.012128f
C219 VDD2.n36 B 0.011454f
C220 VDD2.n37 B 0.021316f
C221 VDD2.n38 B 0.021316f
C222 VDD2.n39 B 0.011454f
C223 VDD2.n40 B 0.012128f
C224 VDD2.n41 B 0.027074f
C225 VDD2.n42 B 0.027074f
C226 VDD2.n43 B 0.012128f
C227 VDD2.n44 B 0.011454f
C228 VDD2.n45 B 0.021316f
C229 VDD2.n46 B 0.021316f
C230 VDD2.n47 B 0.011454f
C231 VDD2.n48 B 0.012128f
C232 VDD2.n49 B 0.027074f
C233 VDD2.n50 B 0.027074f
C234 VDD2.n51 B 0.012128f
C235 VDD2.n52 B 0.011454f
C236 VDD2.n53 B 0.021316f
C237 VDD2.n54 B 0.021316f
C238 VDD2.n55 B 0.011454f
C239 VDD2.n56 B 0.012128f
C240 VDD2.n57 B 0.027074f
C241 VDD2.n58 B 0.027074f
C242 VDD2.n59 B 0.012128f
C243 VDD2.n60 B 0.011454f
C244 VDD2.n61 B 0.021316f
C245 VDD2.n62 B 0.021316f
C246 VDD2.n63 B 0.011454f
C247 VDD2.n64 B 0.012128f
C248 VDD2.n65 B 0.027074f
C249 VDD2.n66 B 0.027074f
C250 VDD2.n67 B 0.027074f
C251 VDD2.n68 B 0.012128f
C252 VDD2.n69 B 0.011454f
C253 VDD2.n70 B 0.021316f
C254 VDD2.n71 B 0.021316f
C255 VDD2.n72 B 0.011454f
C256 VDD2.n73 B 0.011791f
C257 VDD2.n74 B 0.011791f
C258 VDD2.n75 B 0.027074f
C259 VDD2.n76 B 0.059373f
C260 VDD2.n77 B 0.012128f
C261 VDD2.n78 B 0.011454f
C262 VDD2.n79 B 0.055968f
C263 VDD2.n80 B 0.577046f
C264 VDD2.n81 B 0.030393f
C265 VDD2.n82 B 0.021316f
C266 VDD2.n83 B 0.011454f
C267 VDD2.n84 B 0.027074f
C268 VDD2.n85 B 0.012128f
C269 VDD2.n86 B 0.021316f
C270 VDD2.n87 B 0.011454f
C271 VDD2.n88 B 0.027074f
C272 VDD2.n89 B 0.027074f
C273 VDD2.n90 B 0.012128f
C274 VDD2.n91 B 0.021316f
C275 VDD2.n92 B 0.011454f
C276 VDD2.n93 B 0.027074f
C277 VDD2.n94 B 0.012128f
C278 VDD2.n95 B 0.021316f
C279 VDD2.n96 B 0.011454f
C280 VDD2.n97 B 0.027074f
C281 VDD2.n98 B 0.012128f
C282 VDD2.n99 B 0.021316f
C283 VDD2.n100 B 0.011454f
C284 VDD2.n101 B 0.027074f
C285 VDD2.n102 B 0.012128f
C286 VDD2.n103 B 0.021316f
C287 VDD2.n104 B 0.011454f
C288 VDD2.n105 B 0.027074f
C289 VDD2.n106 B 0.012128f
C290 VDD2.n107 B 0.138332f
C291 VDD2.t1 B 0.044632f
C292 VDD2.n108 B 0.020305f
C293 VDD2.n109 B 0.015993f
C294 VDD2.n110 B 0.011454f
C295 VDD2.n111 B 1.37414f
C296 VDD2.n112 B 0.021316f
C297 VDD2.n113 B 0.011454f
C298 VDD2.n114 B 0.012128f
C299 VDD2.n115 B 0.027074f
C300 VDD2.n116 B 0.027074f
C301 VDD2.n117 B 0.012128f
C302 VDD2.n118 B 0.011454f
C303 VDD2.n119 B 0.021316f
C304 VDD2.n120 B 0.021316f
C305 VDD2.n121 B 0.011454f
C306 VDD2.n122 B 0.012128f
C307 VDD2.n123 B 0.027074f
C308 VDD2.n124 B 0.027074f
C309 VDD2.n125 B 0.012128f
C310 VDD2.n126 B 0.011454f
C311 VDD2.n127 B 0.021316f
C312 VDD2.n128 B 0.021316f
C313 VDD2.n129 B 0.011454f
C314 VDD2.n130 B 0.012128f
C315 VDD2.n131 B 0.027074f
C316 VDD2.n132 B 0.027074f
C317 VDD2.n133 B 0.012128f
C318 VDD2.n134 B 0.011454f
C319 VDD2.n135 B 0.021316f
C320 VDD2.n136 B 0.021316f
C321 VDD2.n137 B 0.011454f
C322 VDD2.n138 B 0.012128f
C323 VDD2.n139 B 0.027074f
C324 VDD2.n140 B 0.027074f
C325 VDD2.n141 B 0.012128f
C326 VDD2.n142 B 0.011454f
C327 VDD2.n143 B 0.021316f
C328 VDD2.n144 B 0.021316f
C329 VDD2.n145 B 0.011454f
C330 VDD2.n146 B 0.012128f
C331 VDD2.n147 B 0.027074f
C332 VDD2.n148 B 0.027074f
C333 VDD2.n149 B 0.012128f
C334 VDD2.n150 B 0.011454f
C335 VDD2.n151 B 0.021316f
C336 VDD2.n152 B 0.021316f
C337 VDD2.n153 B 0.011454f
C338 VDD2.n154 B 0.011791f
C339 VDD2.n155 B 0.011791f
C340 VDD2.n156 B 0.027074f
C341 VDD2.n157 B 0.059373f
C342 VDD2.n158 B 0.012128f
C343 VDD2.n159 B 0.011454f
C344 VDD2.n160 B 0.055968f
C345 VDD2.n161 B 0.048167f
C346 VDD2.n162 B 2.5569f
C347 VTAIL.n0 B 0.024153f
C348 VTAIL.n1 B 0.01694f
C349 VTAIL.n2 B 0.009103f
C350 VTAIL.n3 B 0.021516f
C351 VTAIL.n4 B 0.009638f
C352 VTAIL.n5 B 0.01694f
C353 VTAIL.n6 B 0.009103f
C354 VTAIL.n7 B 0.021516f
C355 VTAIL.n8 B 0.009638f
C356 VTAIL.n9 B 0.01694f
C357 VTAIL.n10 B 0.009103f
C358 VTAIL.n11 B 0.021516f
C359 VTAIL.n12 B 0.009638f
C360 VTAIL.n13 B 0.01694f
C361 VTAIL.n14 B 0.009103f
C362 VTAIL.n15 B 0.021516f
C363 VTAIL.n16 B 0.009638f
C364 VTAIL.n17 B 0.01694f
C365 VTAIL.n18 B 0.009103f
C366 VTAIL.n19 B 0.021516f
C367 VTAIL.n20 B 0.009638f
C368 VTAIL.n21 B 0.01694f
C369 VTAIL.n22 B 0.009103f
C370 VTAIL.n23 B 0.021516f
C371 VTAIL.n24 B 0.009638f
C372 VTAIL.n25 B 0.109934f
C373 VTAIL.t1 B 0.035469f
C374 VTAIL.n26 B 0.016137f
C375 VTAIL.n27 B 0.01271f
C376 VTAIL.n28 B 0.009103f
C377 VTAIL.n29 B 1.09204f
C378 VTAIL.n30 B 0.01694f
C379 VTAIL.n31 B 0.009103f
C380 VTAIL.n32 B 0.009638f
C381 VTAIL.n33 B 0.021516f
C382 VTAIL.n34 B 0.021516f
C383 VTAIL.n35 B 0.009638f
C384 VTAIL.n36 B 0.009103f
C385 VTAIL.n37 B 0.01694f
C386 VTAIL.n38 B 0.01694f
C387 VTAIL.n39 B 0.009103f
C388 VTAIL.n40 B 0.009638f
C389 VTAIL.n41 B 0.021516f
C390 VTAIL.n42 B 0.021516f
C391 VTAIL.n43 B 0.009638f
C392 VTAIL.n44 B 0.009103f
C393 VTAIL.n45 B 0.01694f
C394 VTAIL.n46 B 0.01694f
C395 VTAIL.n47 B 0.009103f
C396 VTAIL.n48 B 0.009638f
C397 VTAIL.n49 B 0.021516f
C398 VTAIL.n50 B 0.021516f
C399 VTAIL.n51 B 0.009638f
C400 VTAIL.n52 B 0.009103f
C401 VTAIL.n53 B 0.01694f
C402 VTAIL.n54 B 0.01694f
C403 VTAIL.n55 B 0.009103f
C404 VTAIL.n56 B 0.009638f
C405 VTAIL.n57 B 0.021516f
C406 VTAIL.n58 B 0.021516f
C407 VTAIL.n59 B 0.009638f
C408 VTAIL.n60 B 0.009103f
C409 VTAIL.n61 B 0.01694f
C410 VTAIL.n62 B 0.01694f
C411 VTAIL.n63 B 0.009103f
C412 VTAIL.n64 B 0.009638f
C413 VTAIL.n65 B 0.021516f
C414 VTAIL.n66 B 0.021516f
C415 VTAIL.n67 B 0.021516f
C416 VTAIL.n68 B 0.009638f
C417 VTAIL.n69 B 0.009103f
C418 VTAIL.n70 B 0.01694f
C419 VTAIL.n71 B 0.01694f
C420 VTAIL.n72 B 0.009103f
C421 VTAIL.n73 B 0.00937f
C422 VTAIL.n74 B 0.00937f
C423 VTAIL.n75 B 0.021516f
C424 VTAIL.n76 B 0.047184f
C425 VTAIL.n77 B 0.009638f
C426 VTAIL.n78 B 0.009103f
C427 VTAIL.n79 B 0.044478f
C428 VTAIL.n80 B 0.026618f
C429 VTAIL.n81 B 1.07447f
C430 VTAIL.n82 B 0.024153f
C431 VTAIL.n83 B 0.01694f
C432 VTAIL.n84 B 0.009103f
C433 VTAIL.n85 B 0.021516f
C434 VTAIL.n86 B 0.009638f
C435 VTAIL.n87 B 0.01694f
C436 VTAIL.n88 B 0.009103f
C437 VTAIL.n89 B 0.021516f
C438 VTAIL.n90 B 0.021516f
C439 VTAIL.n91 B 0.009638f
C440 VTAIL.n92 B 0.01694f
C441 VTAIL.n93 B 0.009103f
C442 VTAIL.n94 B 0.021516f
C443 VTAIL.n95 B 0.009638f
C444 VTAIL.n96 B 0.01694f
C445 VTAIL.n97 B 0.009103f
C446 VTAIL.n98 B 0.021516f
C447 VTAIL.n99 B 0.009638f
C448 VTAIL.n100 B 0.01694f
C449 VTAIL.n101 B 0.009103f
C450 VTAIL.n102 B 0.021516f
C451 VTAIL.n103 B 0.009638f
C452 VTAIL.n104 B 0.01694f
C453 VTAIL.n105 B 0.009103f
C454 VTAIL.n106 B 0.021516f
C455 VTAIL.n107 B 0.009638f
C456 VTAIL.n108 B 0.109934f
C457 VTAIL.t2 B 0.035469f
C458 VTAIL.n109 B 0.016137f
C459 VTAIL.n110 B 0.01271f
C460 VTAIL.n111 B 0.009103f
C461 VTAIL.n112 B 1.09204f
C462 VTAIL.n113 B 0.01694f
C463 VTAIL.n114 B 0.009103f
C464 VTAIL.n115 B 0.009638f
C465 VTAIL.n116 B 0.021516f
C466 VTAIL.n117 B 0.021516f
C467 VTAIL.n118 B 0.009638f
C468 VTAIL.n119 B 0.009103f
C469 VTAIL.n120 B 0.01694f
C470 VTAIL.n121 B 0.01694f
C471 VTAIL.n122 B 0.009103f
C472 VTAIL.n123 B 0.009638f
C473 VTAIL.n124 B 0.021516f
C474 VTAIL.n125 B 0.021516f
C475 VTAIL.n126 B 0.009638f
C476 VTAIL.n127 B 0.009103f
C477 VTAIL.n128 B 0.01694f
C478 VTAIL.n129 B 0.01694f
C479 VTAIL.n130 B 0.009103f
C480 VTAIL.n131 B 0.009638f
C481 VTAIL.n132 B 0.021516f
C482 VTAIL.n133 B 0.021516f
C483 VTAIL.n134 B 0.009638f
C484 VTAIL.n135 B 0.009103f
C485 VTAIL.n136 B 0.01694f
C486 VTAIL.n137 B 0.01694f
C487 VTAIL.n138 B 0.009103f
C488 VTAIL.n139 B 0.009638f
C489 VTAIL.n140 B 0.021516f
C490 VTAIL.n141 B 0.021516f
C491 VTAIL.n142 B 0.009638f
C492 VTAIL.n143 B 0.009103f
C493 VTAIL.n144 B 0.01694f
C494 VTAIL.n145 B 0.01694f
C495 VTAIL.n146 B 0.009103f
C496 VTAIL.n147 B 0.009638f
C497 VTAIL.n148 B 0.021516f
C498 VTAIL.n149 B 0.021516f
C499 VTAIL.n150 B 0.009638f
C500 VTAIL.n151 B 0.009103f
C501 VTAIL.n152 B 0.01694f
C502 VTAIL.n153 B 0.01694f
C503 VTAIL.n154 B 0.009103f
C504 VTAIL.n155 B 0.00937f
C505 VTAIL.n156 B 0.00937f
C506 VTAIL.n157 B 0.021516f
C507 VTAIL.n158 B 0.047184f
C508 VTAIL.n159 B 0.009638f
C509 VTAIL.n160 B 0.009103f
C510 VTAIL.n161 B 0.044478f
C511 VTAIL.n162 B 0.026618f
C512 VTAIL.n163 B 1.08212f
C513 VTAIL.n164 B 0.024153f
C514 VTAIL.n165 B 0.01694f
C515 VTAIL.n166 B 0.009103f
C516 VTAIL.n167 B 0.021516f
C517 VTAIL.n168 B 0.009638f
C518 VTAIL.n169 B 0.01694f
C519 VTAIL.n170 B 0.009103f
C520 VTAIL.n171 B 0.021516f
C521 VTAIL.n172 B 0.021516f
C522 VTAIL.n173 B 0.009638f
C523 VTAIL.n174 B 0.01694f
C524 VTAIL.n175 B 0.009103f
C525 VTAIL.n176 B 0.021516f
C526 VTAIL.n177 B 0.009638f
C527 VTAIL.n178 B 0.01694f
C528 VTAIL.n179 B 0.009103f
C529 VTAIL.n180 B 0.021516f
C530 VTAIL.n181 B 0.009638f
C531 VTAIL.n182 B 0.01694f
C532 VTAIL.n183 B 0.009103f
C533 VTAIL.n184 B 0.021516f
C534 VTAIL.n185 B 0.009638f
C535 VTAIL.n186 B 0.01694f
C536 VTAIL.n187 B 0.009103f
C537 VTAIL.n188 B 0.021516f
C538 VTAIL.n189 B 0.009638f
C539 VTAIL.n190 B 0.109934f
C540 VTAIL.t0 B 0.035469f
C541 VTAIL.n191 B 0.016137f
C542 VTAIL.n192 B 0.01271f
C543 VTAIL.n193 B 0.009103f
C544 VTAIL.n194 B 1.09204f
C545 VTAIL.n195 B 0.01694f
C546 VTAIL.n196 B 0.009103f
C547 VTAIL.n197 B 0.009638f
C548 VTAIL.n198 B 0.021516f
C549 VTAIL.n199 B 0.021516f
C550 VTAIL.n200 B 0.009638f
C551 VTAIL.n201 B 0.009103f
C552 VTAIL.n202 B 0.01694f
C553 VTAIL.n203 B 0.01694f
C554 VTAIL.n204 B 0.009103f
C555 VTAIL.n205 B 0.009638f
C556 VTAIL.n206 B 0.021516f
C557 VTAIL.n207 B 0.021516f
C558 VTAIL.n208 B 0.009638f
C559 VTAIL.n209 B 0.009103f
C560 VTAIL.n210 B 0.01694f
C561 VTAIL.n211 B 0.01694f
C562 VTAIL.n212 B 0.009103f
C563 VTAIL.n213 B 0.009638f
C564 VTAIL.n214 B 0.021516f
C565 VTAIL.n215 B 0.021516f
C566 VTAIL.n216 B 0.009638f
C567 VTAIL.n217 B 0.009103f
C568 VTAIL.n218 B 0.01694f
C569 VTAIL.n219 B 0.01694f
C570 VTAIL.n220 B 0.009103f
C571 VTAIL.n221 B 0.009638f
C572 VTAIL.n222 B 0.021516f
C573 VTAIL.n223 B 0.021516f
C574 VTAIL.n224 B 0.009638f
C575 VTAIL.n225 B 0.009103f
C576 VTAIL.n226 B 0.01694f
C577 VTAIL.n227 B 0.01694f
C578 VTAIL.n228 B 0.009103f
C579 VTAIL.n229 B 0.009638f
C580 VTAIL.n230 B 0.021516f
C581 VTAIL.n231 B 0.021516f
C582 VTAIL.n232 B 0.009638f
C583 VTAIL.n233 B 0.009103f
C584 VTAIL.n234 B 0.01694f
C585 VTAIL.n235 B 0.01694f
C586 VTAIL.n236 B 0.009103f
C587 VTAIL.n237 B 0.00937f
C588 VTAIL.n238 B 0.00937f
C589 VTAIL.n239 B 0.021516f
C590 VTAIL.n240 B 0.047184f
C591 VTAIL.n241 B 0.009638f
C592 VTAIL.n242 B 0.009103f
C593 VTAIL.n243 B 0.044478f
C594 VTAIL.n244 B 0.026618f
C595 VTAIL.n245 B 1.03883f
C596 VTAIL.n246 B 0.024153f
C597 VTAIL.n247 B 0.01694f
C598 VTAIL.n248 B 0.009103f
C599 VTAIL.n249 B 0.021516f
C600 VTAIL.n250 B 0.009638f
C601 VTAIL.n251 B 0.01694f
C602 VTAIL.n252 B 0.009103f
C603 VTAIL.n253 B 0.021516f
C604 VTAIL.n254 B 0.009638f
C605 VTAIL.n255 B 0.01694f
C606 VTAIL.n256 B 0.009103f
C607 VTAIL.n257 B 0.021516f
C608 VTAIL.n258 B 0.009638f
C609 VTAIL.n259 B 0.01694f
C610 VTAIL.n260 B 0.009103f
C611 VTAIL.n261 B 0.021516f
C612 VTAIL.n262 B 0.009638f
C613 VTAIL.n263 B 0.01694f
C614 VTAIL.n264 B 0.009103f
C615 VTAIL.n265 B 0.021516f
C616 VTAIL.n266 B 0.009638f
C617 VTAIL.n267 B 0.01694f
C618 VTAIL.n268 B 0.009103f
C619 VTAIL.n269 B 0.021516f
C620 VTAIL.n270 B 0.009638f
C621 VTAIL.n271 B 0.109934f
C622 VTAIL.t3 B 0.035469f
C623 VTAIL.n272 B 0.016137f
C624 VTAIL.n273 B 0.01271f
C625 VTAIL.n274 B 0.009103f
C626 VTAIL.n275 B 1.09204f
C627 VTAIL.n276 B 0.01694f
C628 VTAIL.n277 B 0.009103f
C629 VTAIL.n278 B 0.009638f
C630 VTAIL.n279 B 0.021516f
C631 VTAIL.n280 B 0.021516f
C632 VTAIL.n281 B 0.009638f
C633 VTAIL.n282 B 0.009103f
C634 VTAIL.n283 B 0.01694f
C635 VTAIL.n284 B 0.01694f
C636 VTAIL.n285 B 0.009103f
C637 VTAIL.n286 B 0.009638f
C638 VTAIL.n287 B 0.021516f
C639 VTAIL.n288 B 0.021516f
C640 VTAIL.n289 B 0.009638f
C641 VTAIL.n290 B 0.009103f
C642 VTAIL.n291 B 0.01694f
C643 VTAIL.n292 B 0.01694f
C644 VTAIL.n293 B 0.009103f
C645 VTAIL.n294 B 0.009638f
C646 VTAIL.n295 B 0.021516f
C647 VTAIL.n296 B 0.021516f
C648 VTAIL.n297 B 0.009638f
C649 VTAIL.n298 B 0.009103f
C650 VTAIL.n299 B 0.01694f
C651 VTAIL.n300 B 0.01694f
C652 VTAIL.n301 B 0.009103f
C653 VTAIL.n302 B 0.009638f
C654 VTAIL.n303 B 0.021516f
C655 VTAIL.n304 B 0.021516f
C656 VTAIL.n305 B 0.009638f
C657 VTAIL.n306 B 0.009103f
C658 VTAIL.n307 B 0.01694f
C659 VTAIL.n308 B 0.01694f
C660 VTAIL.n309 B 0.009103f
C661 VTAIL.n310 B 0.009638f
C662 VTAIL.n311 B 0.021516f
C663 VTAIL.n312 B 0.021516f
C664 VTAIL.n313 B 0.021516f
C665 VTAIL.n314 B 0.009638f
C666 VTAIL.n315 B 0.009103f
C667 VTAIL.n316 B 0.01694f
C668 VTAIL.n317 B 0.01694f
C669 VTAIL.n318 B 0.009103f
C670 VTAIL.n319 B 0.00937f
C671 VTAIL.n320 B 0.00937f
C672 VTAIL.n321 B 0.021516f
C673 VTAIL.n322 B 0.047184f
C674 VTAIL.n323 B 0.009638f
C675 VTAIL.n324 B 0.009103f
C676 VTAIL.n325 B 0.044478f
C677 VTAIL.n326 B 0.026618f
C678 VTAIL.n327 B 0.999181f
C679 VN.t1 B 1.28401f
C680 VN.t0 B 1.39583f
.ends

