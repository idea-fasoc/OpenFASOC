* NGSPICE file created from diff_pair_sample_1690.ext - technology: sky130A

.subckt diff_pair_sample_1690 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0 ps=0 w=1.7 l=0.68
X2 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0 ps=0 w=1.7 l=0.68
X3 VTAIL.t13 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0.2805 ps=2.03 w=1.7 l=0.68
X4 VDD1.t7 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X5 VDD2.t5 VN.t2 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X6 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0 ps=0 w=1.7 l=0.68
X7 VTAIL.t12 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X8 VTAIL.t7 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0.2805 ps=2.03 w=1.7 l=0.68
X9 VDD2.t3 VN.t4 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.663 ps=4.18 w=1.7 l=0.68
X10 VTAIL.t9 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X11 VDD2.t1 VN.t6 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.663 ps=4.18 w=1.7 l=0.68
X12 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.663 ps=4.18 w=1.7 l=0.68
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0 ps=0 w=1.7 l=0.68
X14 VDD1.t4 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.663 ps=4.18 w=1.7 l=0.68
X15 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X16 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
X17 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0.2805 ps=2.03 w=1.7 l=0.68
X18 VTAIL.t14 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.663 pd=4.18 as=0.2805 ps=2.03 w=1.7 l=0.68
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2805 pd=2.03 as=0.2805 ps=2.03 w=1.7 l=0.68
R0 VN.n9 VN.n8 161.3
R1 VN.n19 VN.n18 161.3
R2 VN.n17 VN.n10 161.3
R3 VN.n16 VN.n15 161.3
R4 VN.n14 VN.n11 161.3
R5 VN.n7 VN.n0 161.3
R6 VN.n6 VN.n5 161.3
R7 VN.n4 VN.n1 161.3
R8 VN.n3 VN.t1 139.417
R9 VN.n13 VN.t6 139.417
R10 VN.n2 VN.t2 118.019
R11 VN.n6 VN.t5 118.019
R12 VN.n8 VN.t4 118.019
R13 VN.n12 VN.t3 118.019
R14 VN.n16 VN.t0 118.019
R15 VN.n18 VN.t7 118.019
R16 VN.n14 VN.n13 44.853
R17 VN.n4 VN.n3 44.853
R18 VN VN.n19 34.4494
R19 VN.n8 VN.n7 25.5611
R20 VN.n18 VN.n17 25.5611
R21 VN.n2 VN.n1 24.1005
R22 VN.n6 VN.n1 24.1005
R23 VN.n16 VN.n11 24.1005
R24 VN.n12 VN.n11 24.1005
R25 VN.n7 VN.n6 22.6399
R26 VN.n17 VN.n16 22.6399
R27 VN.n3 VN.n2 20.5405
R28 VN.n13 VN.n12 20.5405
R29 VN.n19 VN.n10 0.189894
R30 VN.n15 VN.n10 0.189894
R31 VN.n15 VN.n14 0.189894
R32 VN.n5 VN.n4 0.189894
R33 VN.n5 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VTAIL.n15 VTAIL.t8 112.109
R37 VTAIL.n2 VTAIL.t13 112.109
R38 VTAIL.n3 VTAIL.t5 112.109
R39 VTAIL.n6 VTAIL.t4 112.109
R40 VTAIL.n14 VTAIL.t6 112.109
R41 VTAIL.n11 VTAIL.t7 112.109
R42 VTAIL.n10 VTAIL.t10 112.109
R43 VTAIL.n7 VTAIL.t14 112.109
R44 VTAIL.n1 VTAIL.n0 100.462
R45 VTAIL.n5 VTAIL.n4 100.462
R46 VTAIL.n13 VTAIL.n12 100.462
R47 VTAIL.n9 VTAIL.n8 100.462
R48 VTAIL.n15 VTAIL.n14 14.7031
R49 VTAIL.n7 VTAIL.n6 14.7031
R50 VTAIL.n0 VTAIL.t15 11.6476
R51 VTAIL.n0 VTAIL.t9 11.6476
R52 VTAIL.n4 VTAIL.t3 11.6476
R53 VTAIL.n4 VTAIL.t1 11.6476
R54 VTAIL.n12 VTAIL.t2 11.6476
R55 VTAIL.n12 VTAIL.t0 11.6476
R56 VTAIL.n8 VTAIL.t11 11.6476
R57 VTAIL.n8 VTAIL.t12 11.6476
R58 VTAIL.n9 VTAIL.n7 0.87119
R59 VTAIL.n10 VTAIL.n9 0.87119
R60 VTAIL.n13 VTAIL.n11 0.87119
R61 VTAIL.n14 VTAIL.n13 0.87119
R62 VTAIL.n6 VTAIL.n5 0.87119
R63 VTAIL.n5 VTAIL.n3 0.87119
R64 VTAIL.n2 VTAIL.n1 0.87119
R65 VTAIL VTAIL.n15 0.813
R66 VTAIL.n11 VTAIL.n10 0.470328
R67 VTAIL.n3 VTAIL.n2 0.470328
R68 VTAIL VTAIL.n1 0.0586897
R69 VDD2.n2 VDD2.n1 117.519
R70 VDD2.n2 VDD2.n0 117.519
R71 VDD2 VDD2.n5 117.517
R72 VDD2.n4 VDD2.n3 117.139
R73 VDD2.n4 VDD2.n2 29.0989
R74 VDD2.n5 VDD2.t4 11.6476
R75 VDD2.n5 VDD2.t1 11.6476
R76 VDD2.n3 VDD2.t0 11.6476
R77 VDD2.n3 VDD2.t7 11.6476
R78 VDD2.n1 VDD2.t2 11.6476
R79 VDD2.n1 VDD2.t3 11.6476
R80 VDD2.n0 VDD2.t6 11.6476
R81 VDD2.n0 VDD2.t5 11.6476
R82 VDD2 VDD2.n4 0.494034
R83 B.n353 B.n352 585
R84 B.n125 B.n61 585
R85 B.n124 B.n123 585
R86 B.n122 B.n121 585
R87 B.n120 B.n119 585
R88 B.n118 B.n117 585
R89 B.n116 B.n115 585
R90 B.n114 B.n113 585
R91 B.n112 B.n111 585
R92 B.n110 B.n109 585
R93 B.n108 B.n107 585
R94 B.n105 B.n104 585
R95 B.n103 B.n102 585
R96 B.n101 B.n100 585
R97 B.n99 B.n98 585
R98 B.n97 B.n96 585
R99 B.n95 B.n94 585
R100 B.n93 B.n92 585
R101 B.n91 B.n90 585
R102 B.n89 B.n88 585
R103 B.n87 B.n86 585
R104 B.n84 B.n83 585
R105 B.n82 B.n81 585
R106 B.n80 B.n79 585
R107 B.n78 B.n77 585
R108 B.n76 B.n75 585
R109 B.n74 B.n73 585
R110 B.n72 B.n71 585
R111 B.n70 B.n69 585
R112 B.n68 B.n67 585
R113 B.n46 B.n45 585
R114 B.n358 B.n357 585
R115 B.n351 B.n62 585
R116 B.n62 B.n43 585
R117 B.n350 B.n42 585
R118 B.n362 B.n42 585
R119 B.n349 B.n41 585
R120 B.n363 B.n41 585
R121 B.n348 B.n40 585
R122 B.n364 B.n40 585
R123 B.n347 B.n346 585
R124 B.n346 B.n39 585
R125 B.n345 B.n35 585
R126 B.n370 B.n35 585
R127 B.n344 B.n34 585
R128 B.n371 B.n34 585
R129 B.n343 B.n33 585
R130 B.n372 B.n33 585
R131 B.n342 B.n341 585
R132 B.n341 B.n29 585
R133 B.n340 B.n28 585
R134 B.n378 B.n28 585
R135 B.n339 B.n27 585
R136 B.n379 B.n27 585
R137 B.n338 B.n26 585
R138 B.t6 B.n26 585
R139 B.n337 B.n336 585
R140 B.n336 B.n22 585
R141 B.n335 B.n21 585
R142 B.n385 B.n21 585
R143 B.n334 B.n20 585
R144 B.n386 B.n20 585
R145 B.n333 B.n19 585
R146 B.n387 B.n19 585
R147 B.n332 B.n331 585
R148 B.n331 B.n18 585
R149 B.n330 B.n14 585
R150 B.n393 B.n14 585
R151 B.n329 B.n13 585
R152 B.n394 B.n13 585
R153 B.n328 B.n12 585
R154 B.n395 B.n12 585
R155 B.n327 B.n326 585
R156 B.n326 B.n8 585
R157 B.n325 B.n7 585
R158 B.n401 B.n7 585
R159 B.n324 B.n6 585
R160 B.n402 B.n6 585
R161 B.n323 B.n5 585
R162 B.n403 B.n5 585
R163 B.n322 B.n321 585
R164 B.n321 B.n4 585
R165 B.n320 B.n126 585
R166 B.n320 B.n319 585
R167 B.n310 B.n127 585
R168 B.n128 B.n127 585
R169 B.n312 B.n311 585
R170 B.n313 B.n312 585
R171 B.n309 B.n133 585
R172 B.n133 B.n132 585
R173 B.n308 B.n307 585
R174 B.n307 B.n306 585
R175 B.n135 B.n134 585
R176 B.n299 B.n135 585
R177 B.n298 B.n297 585
R178 B.n300 B.n298 585
R179 B.n296 B.n140 585
R180 B.n140 B.n139 585
R181 B.n295 B.n294 585
R182 B.n294 B.n293 585
R183 B.n142 B.n141 585
R184 B.n143 B.n142 585
R185 B.n287 B.n286 585
R186 B.t4 B.n287 585
R187 B.n285 B.n148 585
R188 B.n148 B.n147 585
R189 B.n284 B.n283 585
R190 B.n283 B.n282 585
R191 B.n150 B.n149 585
R192 B.n151 B.n150 585
R193 B.n275 B.n274 585
R194 B.n276 B.n275 585
R195 B.n273 B.n156 585
R196 B.n156 B.n155 585
R197 B.n272 B.n271 585
R198 B.n271 B.n270 585
R199 B.n158 B.n157 585
R200 B.n263 B.n158 585
R201 B.n262 B.n261 585
R202 B.n264 B.n262 585
R203 B.n260 B.n163 585
R204 B.n163 B.n162 585
R205 B.n259 B.n258 585
R206 B.n258 B.n257 585
R207 B.n165 B.n164 585
R208 B.n166 B.n165 585
R209 B.n253 B.n252 585
R210 B.n169 B.n168 585
R211 B.n249 B.n248 585
R212 B.n250 B.n249 585
R213 B.n247 B.n185 585
R214 B.n246 B.n245 585
R215 B.n244 B.n243 585
R216 B.n242 B.n241 585
R217 B.n240 B.n239 585
R218 B.n238 B.n237 585
R219 B.n236 B.n235 585
R220 B.n234 B.n233 585
R221 B.n232 B.n231 585
R222 B.n230 B.n229 585
R223 B.n228 B.n227 585
R224 B.n226 B.n225 585
R225 B.n224 B.n223 585
R226 B.n222 B.n221 585
R227 B.n220 B.n219 585
R228 B.n218 B.n217 585
R229 B.n216 B.n215 585
R230 B.n214 B.n213 585
R231 B.n212 B.n211 585
R232 B.n210 B.n209 585
R233 B.n208 B.n207 585
R234 B.n206 B.n205 585
R235 B.n204 B.n203 585
R236 B.n202 B.n201 585
R237 B.n200 B.n199 585
R238 B.n198 B.n197 585
R239 B.n196 B.n195 585
R240 B.n194 B.n193 585
R241 B.n192 B.n184 585
R242 B.n250 B.n184 585
R243 B.n254 B.n167 585
R244 B.n167 B.n166 585
R245 B.n256 B.n255 585
R246 B.n257 B.n256 585
R247 B.n161 B.n160 585
R248 B.n162 B.n161 585
R249 B.n266 B.n265 585
R250 B.n265 B.n264 585
R251 B.n267 B.n159 585
R252 B.n263 B.n159 585
R253 B.n269 B.n268 585
R254 B.n270 B.n269 585
R255 B.n154 B.n153 585
R256 B.n155 B.n154 585
R257 B.n278 B.n277 585
R258 B.n277 B.n276 585
R259 B.n279 B.n152 585
R260 B.n152 B.n151 585
R261 B.n281 B.n280 585
R262 B.n282 B.n281 585
R263 B.n146 B.n145 585
R264 B.n147 B.n146 585
R265 B.n289 B.n288 585
R266 B.n288 B.t4 585
R267 B.n290 B.n144 585
R268 B.n144 B.n143 585
R269 B.n292 B.n291 585
R270 B.n293 B.n292 585
R271 B.n138 B.n137 585
R272 B.n139 B.n138 585
R273 B.n302 B.n301 585
R274 B.n301 B.n300 585
R275 B.n303 B.n136 585
R276 B.n299 B.n136 585
R277 B.n305 B.n304 585
R278 B.n306 B.n305 585
R279 B.n131 B.n130 585
R280 B.n132 B.n131 585
R281 B.n315 B.n314 585
R282 B.n314 B.n313 585
R283 B.n316 B.n129 585
R284 B.n129 B.n128 585
R285 B.n318 B.n317 585
R286 B.n319 B.n318 585
R287 B.n2 B.n0 585
R288 B.n4 B.n2 585
R289 B.n3 B.n1 585
R290 B.n402 B.n3 585
R291 B.n400 B.n399 585
R292 B.n401 B.n400 585
R293 B.n398 B.n9 585
R294 B.n9 B.n8 585
R295 B.n397 B.n396 585
R296 B.n396 B.n395 585
R297 B.n11 B.n10 585
R298 B.n394 B.n11 585
R299 B.n392 B.n391 585
R300 B.n393 B.n392 585
R301 B.n390 B.n15 585
R302 B.n18 B.n15 585
R303 B.n389 B.n388 585
R304 B.n388 B.n387 585
R305 B.n17 B.n16 585
R306 B.n386 B.n17 585
R307 B.n384 B.n383 585
R308 B.n385 B.n384 585
R309 B.n382 B.n23 585
R310 B.n23 B.n22 585
R311 B.n381 B.n380 585
R312 B.n380 B.t6 585
R313 B.n25 B.n24 585
R314 B.n379 B.n25 585
R315 B.n377 B.n376 585
R316 B.n378 B.n377 585
R317 B.n375 B.n30 585
R318 B.n30 B.n29 585
R319 B.n374 B.n373 585
R320 B.n373 B.n372 585
R321 B.n32 B.n31 585
R322 B.n371 B.n32 585
R323 B.n369 B.n368 585
R324 B.n370 B.n369 585
R325 B.n367 B.n36 585
R326 B.n39 B.n36 585
R327 B.n366 B.n365 585
R328 B.n365 B.n364 585
R329 B.n38 B.n37 585
R330 B.n363 B.n38 585
R331 B.n361 B.n360 585
R332 B.n362 B.n361 585
R333 B.n359 B.n44 585
R334 B.n44 B.n43 585
R335 B.n405 B.n404 585
R336 B.n404 B.n403 585
R337 B.n252 B.n167 511.721
R338 B.n357 B.n44 511.721
R339 B.n184 B.n165 511.721
R340 B.n353 B.n62 511.721
R341 B.n189 B.t19 263.469
R342 B.n186 B.t12 263.469
R343 B.n65 B.t16 263.469
R344 B.n63 B.t8 263.469
R345 B.n355 B.n354 256.663
R346 B.n355 B.n60 256.663
R347 B.n355 B.n59 256.663
R348 B.n355 B.n58 256.663
R349 B.n355 B.n57 256.663
R350 B.n355 B.n56 256.663
R351 B.n355 B.n55 256.663
R352 B.n355 B.n54 256.663
R353 B.n355 B.n53 256.663
R354 B.n355 B.n52 256.663
R355 B.n355 B.n51 256.663
R356 B.n355 B.n50 256.663
R357 B.n355 B.n49 256.663
R358 B.n355 B.n48 256.663
R359 B.n355 B.n47 256.663
R360 B.n356 B.n355 256.663
R361 B.n251 B.n250 256.663
R362 B.n250 B.n170 256.663
R363 B.n250 B.n171 256.663
R364 B.n250 B.n172 256.663
R365 B.n250 B.n173 256.663
R366 B.n250 B.n174 256.663
R367 B.n250 B.n175 256.663
R368 B.n250 B.n176 256.663
R369 B.n250 B.n177 256.663
R370 B.n250 B.n178 256.663
R371 B.n250 B.n179 256.663
R372 B.n250 B.n180 256.663
R373 B.n250 B.n181 256.663
R374 B.n250 B.n182 256.663
R375 B.n250 B.n183 256.663
R376 B.n250 B.n166 190.825
R377 B.n355 B.n43 190.825
R378 B.n256 B.n167 163.367
R379 B.n256 B.n161 163.367
R380 B.n265 B.n161 163.367
R381 B.n265 B.n159 163.367
R382 B.n269 B.n159 163.367
R383 B.n269 B.n154 163.367
R384 B.n277 B.n154 163.367
R385 B.n277 B.n152 163.367
R386 B.n281 B.n152 163.367
R387 B.n281 B.n146 163.367
R388 B.n288 B.n146 163.367
R389 B.n288 B.n144 163.367
R390 B.n292 B.n144 163.367
R391 B.n292 B.n138 163.367
R392 B.n301 B.n138 163.367
R393 B.n301 B.n136 163.367
R394 B.n305 B.n136 163.367
R395 B.n305 B.n131 163.367
R396 B.n314 B.n131 163.367
R397 B.n314 B.n129 163.367
R398 B.n318 B.n129 163.367
R399 B.n318 B.n2 163.367
R400 B.n404 B.n2 163.367
R401 B.n404 B.n3 163.367
R402 B.n400 B.n3 163.367
R403 B.n400 B.n9 163.367
R404 B.n396 B.n9 163.367
R405 B.n396 B.n11 163.367
R406 B.n392 B.n11 163.367
R407 B.n392 B.n15 163.367
R408 B.n388 B.n15 163.367
R409 B.n388 B.n17 163.367
R410 B.n384 B.n17 163.367
R411 B.n384 B.n23 163.367
R412 B.n380 B.n23 163.367
R413 B.n380 B.n25 163.367
R414 B.n377 B.n25 163.367
R415 B.n377 B.n30 163.367
R416 B.n373 B.n30 163.367
R417 B.n373 B.n32 163.367
R418 B.n369 B.n32 163.367
R419 B.n369 B.n36 163.367
R420 B.n365 B.n36 163.367
R421 B.n365 B.n38 163.367
R422 B.n361 B.n38 163.367
R423 B.n361 B.n44 163.367
R424 B.n249 B.n169 163.367
R425 B.n249 B.n185 163.367
R426 B.n245 B.n244 163.367
R427 B.n241 B.n240 163.367
R428 B.n237 B.n236 163.367
R429 B.n233 B.n232 163.367
R430 B.n229 B.n228 163.367
R431 B.n225 B.n224 163.367
R432 B.n221 B.n220 163.367
R433 B.n217 B.n216 163.367
R434 B.n213 B.n212 163.367
R435 B.n209 B.n208 163.367
R436 B.n205 B.n204 163.367
R437 B.n201 B.n200 163.367
R438 B.n197 B.n196 163.367
R439 B.n193 B.n184 163.367
R440 B.n258 B.n165 163.367
R441 B.n258 B.n163 163.367
R442 B.n262 B.n163 163.367
R443 B.n262 B.n158 163.367
R444 B.n271 B.n158 163.367
R445 B.n271 B.n156 163.367
R446 B.n275 B.n156 163.367
R447 B.n275 B.n150 163.367
R448 B.n283 B.n150 163.367
R449 B.n283 B.n148 163.367
R450 B.n287 B.n148 163.367
R451 B.n287 B.n142 163.367
R452 B.n294 B.n142 163.367
R453 B.n294 B.n140 163.367
R454 B.n298 B.n140 163.367
R455 B.n298 B.n135 163.367
R456 B.n307 B.n135 163.367
R457 B.n307 B.n133 163.367
R458 B.n312 B.n133 163.367
R459 B.n312 B.n127 163.367
R460 B.n320 B.n127 163.367
R461 B.n321 B.n320 163.367
R462 B.n321 B.n5 163.367
R463 B.n6 B.n5 163.367
R464 B.n7 B.n6 163.367
R465 B.n326 B.n7 163.367
R466 B.n326 B.n12 163.367
R467 B.n13 B.n12 163.367
R468 B.n14 B.n13 163.367
R469 B.n331 B.n14 163.367
R470 B.n331 B.n19 163.367
R471 B.n20 B.n19 163.367
R472 B.n21 B.n20 163.367
R473 B.n336 B.n21 163.367
R474 B.n336 B.n26 163.367
R475 B.n27 B.n26 163.367
R476 B.n28 B.n27 163.367
R477 B.n341 B.n28 163.367
R478 B.n341 B.n33 163.367
R479 B.n34 B.n33 163.367
R480 B.n35 B.n34 163.367
R481 B.n346 B.n35 163.367
R482 B.n346 B.n40 163.367
R483 B.n41 B.n40 163.367
R484 B.n42 B.n41 163.367
R485 B.n62 B.n42 163.367
R486 B.n67 B.n46 163.367
R487 B.n71 B.n70 163.367
R488 B.n75 B.n74 163.367
R489 B.n79 B.n78 163.367
R490 B.n83 B.n82 163.367
R491 B.n88 B.n87 163.367
R492 B.n92 B.n91 163.367
R493 B.n96 B.n95 163.367
R494 B.n100 B.n99 163.367
R495 B.n104 B.n103 163.367
R496 B.n109 B.n108 163.367
R497 B.n113 B.n112 163.367
R498 B.n117 B.n116 163.367
R499 B.n121 B.n120 163.367
R500 B.n123 B.n61 163.367
R501 B.n189 B.t21 129.254
R502 B.n63 B.t10 129.254
R503 B.n186 B.t15 129.252
R504 B.n65 B.t17 129.252
R505 B.n190 B.t20 109.665
R506 B.n64 B.t11 109.665
R507 B.n187 B.t14 109.665
R508 B.n66 B.t18 109.665
R509 B.n257 B.n166 107.24
R510 B.n257 B.n162 107.24
R511 B.n264 B.n162 107.24
R512 B.n264 B.n263 107.24
R513 B.n270 B.n155 107.24
R514 B.n276 B.n155 107.24
R515 B.n276 B.n151 107.24
R516 B.n282 B.n151 107.24
R517 B.n282 B.n147 107.24
R518 B.t4 B.n147 107.24
R519 B.t4 B.n143 107.24
R520 B.n293 B.n143 107.24
R521 B.n300 B.n139 107.24
R522 B.n300 B.n299 107.24
R523 B.n306 B.n132 107.24
R524 B.n313 B.n132 107.24
R525 B.n319 B.n128 107.24
R526 B.n319 B.n4 107.24
R527 B.n403 B.n4 107.24
R528 B.n403 B.n402 107.24
R529 B.n402 B.n401 107.24
R530 B.n401 B.n8 107.24
R531 B.n395 B.n394 107.24
R532 B.n394 B.n393 107.24
R533 B.n387 B.n18 107.24
R534 B.n387 B.n386 107.24
R535 B.n385 B.n22 107.24
R536 B.t6 B.n22 107.24
R537 B.t6 B.n379 107.24
R538 B.n379 B.n378 107.24
R539 B.n378 B.n29 107.24
R540 B.n372 B.n29 107.24
R541 B.n372 B.n371 107.24
R542 B.n371 B.n370 107.24
R543 B.n364 B.n39 107.24
R544 B.n364 B.n363 107.24
R545 B.n363 B.n362 107.24
R546 B.n362 B.n43 107.24
R547 B.n293 B.t3 104.087
R548 B.t0 B.n385 104.087
R549 B.n299 B.t1 100.933
R550 B.n18 B.t2 100.933
R551 B.n313 B.t5 97.7783
R552 B.n395 B.t7 97.7783
R553 B.n263 B.t13 88.3159
R554 B.n39 B.t9 88.3159
R555 B.n252 B.n251 71.676
R556 B.n185 B.n170 71.676
R557 B.n244 B.n171 71.676
R558 B.n240 B.n172 71.676
R559 B.n236 B.n173 71.676
R560 B.n232 B.n174 71.676
R561 B.n228 B.n175 71.676
R562 B.n224 B.n176 71.676
R563 B.n220 B.n177 71.676
R564 B.n216 B.n178 71.676
R565 B.n212 B.n179 71.676
R566 B.n208 B.n180 71.676
R567 B.n204 B.n181 71.676
R568 B.n200 B.n182 71.676
R569 B.n196 B.n183 71.676
R570 B.n357 B.n356 71.676
R571 B.n67 B.n47 71.676
R572 B.n71 B.n48 71.676
R573 B.n75 B.n49 71.676
R574 B.n79 B.n50 71.676
R575 B.n83 B.n51 71.676
R576 B.n88 B.n52 71.676
R577 B.n92 B.n53 71.676
R578 B.n96 B.n54 71.676
R579 B.n100 B.n55 71.676
R580 B.n104 B.n56 71.676
R581 B.n109 B.n57 71.676
R582 B.n113 B.n58 71.676
R583 B.n117 B.n59 71.676
R584 B.n121 B.n60 71.676
R585 B.n354 B.n61 71.676
R586 B.n354 B.n353 71.676
R587 B.n123 B.n60 71.676
R588 B.n120 B.n59 71.676
R589 B.n116 B.n58 71.676
R590 B.n112 B.n57 71.676
R591 B.n108 B.n56 71.676
R592 B.n103 B.n55 71.676
R593 B.n99 B.n54 71.676
R594 B.n95 B.n53 71.676
R595 B.n91 B.n52 71.676
R596 B.n87 B.n51 71.676
R597 B.n82 B.n50 71.676
R598 B.n78 B.n49 71.676
R599 B.n74 B.n48 71.676
R600 B.n70 B.n47 71.676
R601 B.n356 B.n46 71.676
R602 B.n251 B.n169 71.676
R603 B.n245 B.n170 71.676
R604 B.n241 B.n171 71.676
R605 B.n237 B.n172 71.676
R606 B.n233 B.n173 71.676
R607 B.n229 B.n174 71.676
R608 B.n225 B.n175 71.676
R609 B.n221 B.n176 71.676
R610 B.n217 B.n177 71.676
R611 B.n213 B.n178 71.676
R612 B.n209 B.n179 71.676
R613 B.n205 B.n180 71.676
R614 B.n201 B.n181 71.676
R615 B.n197 B.n182 71.676
R616 B.n193 B.n183 71.676
R617 B.n191 B.n190 59.5399
R618 B.n188 B.n187 59.5399
R619 B.n85 B.n66 59.5399
R620 B.n106 B.n64 59.5399
R621 B.n359 B.n358 33.2493
R622 B.n352 B.n351 33.2493
R623 B.n192 B.n164 33.2493
R624 B.n254 B.n253 33.2493
R625 B.n190 B.n189 19.5884
R626 B.n187 B.n186 19.5884
R627 B.n66 B.n65 19.5884
R628 B.n64 B.n63 19.5884
R629 B.n270 B.t13 18.9252
R630 B.n370 B.t9 18.9252
R631 B B.n405 18.0485
R632 B.n358 B.n45 10.6151
R633 B.n68 B.n45 10.6151
R634 B.n69 B.n68 10.6151
R635 B.n72 B.n69 10.6151
R636 B.n73 B.n72 10.6151
R637 B.n76 B.n73 10.6151
R638 B.n77 B.n76 10.6151
R639 B.n80 B.n77 10.6151
R640 B.n81 B.n80 10.6151
R641 B.n84 B.n81 10.6151
R642 B.n89 B.n86 10.6151
R643 B.n90 B.n89 10.6151
R644 B.n93 B.n90 10.6151
R645 B.n94 B.n93 10.6151
R646 B.n97 B.n94 10.6151
R647 B.n98 B.n97 10.6151
R648 B.n101 B.n98 10.6151
R649 B.n102 B.n101 10.6151
R650 B.n105 B.n102 10.6151
R651 B.n110 B.n107 10.6151
R652 B.n111 B.n110 10.6151
R653 B.n114 B.n111 10.6151
R654 B.n115 B.n114 10.6151
R655 B.n118 B.n115 10.6151
R656 B.n119 B.n118 10.6151
R657 B.n122 B.n119 10.6151
R658 B.n124 B.n122 10.6151
R659 B.n125 B.n124 10.6151
R660 B.n352 B.n125 10.6151
R661 B.n259 B.n164 10.6151
R662 B.n260 B.n259 10.6151
R663 B.n261 B.n260 10.6151
R664 B.n261 B.n157 10.6151
R665 B.n272 B.n157 10.6151
R666 B.n273 B.n272 10.6151
R667 B.n274 B.n273 10.6151
R668 B.n274 B.n149 10.6151
R669 B.n284 B.n149 10.6151
R670 B.n285 B.n284 10.6151
R671 B.n286 B.n285 10.6151
R672 B.n286 B.n141 10.6151
R673 B.n295 B.n141 10.6151
R674 B.n296 B.n295 10.6151
R675 B.n297 B.n296 10.6151
R676 B.n297 B.n134 10.6151
R677 B.n308 B.n134 10.6151
R678 B.n309 B.n308 10.6151
R679 B.n311 B.n309 10.6151
R680 B.n311 B.n310 10.6151
R681 B.n310 B.n126 10.6151
R682 B.n322 B.n126 10.6151
R683 B.n323 B.n322 10.6151
R684 B.n324 B.n323 10.6151
R685 B.n325 B.n324 10.6151
R686 B.n327 B.n325 10.6151
R687 B.n328 B.n327 10.6151
R688 B.n329 B.n328 10.6151
R689 B.n330 B.n329 10.6151
R690 B.n332 B.n330 10.6151
R691 B.n333 B.n332 10.6151
R692 B.n334 B.n333 10.6151
R693 B.n335 B.n334 10.6151
R694 B.n337 B.n335 10.6151
R695 B.n338 B.n337 10.6151
R696 B.n339 B.n338 10.6151
R697 B.n340 B.n339 10.6151
R698 B.n342 B.n340 10.6151
R699 B.n343 B.n342 10.6151
R700 B.n344 B.n343 10.6151
R701 B.n345 B.n344 10.6151
R702 B.n347 B.n345 10.6151
R703 B.n348 B.n347 10.6151
R704 B.n349 B.n348 10.6151
R705 B.n350 B.n349 10.6151
R706 B.n351 B.n350 10.6151
R707 B.n253 B.n168 10.6151
R708 B.n248 B.n168 10.6151
R709 B.n248 B.n247 10.6151
R710 B.n247 B.n246 10.6151
R711 B.n246 B.n243 10.6151
R712 B.n243 B.n242 10.6151
R713 B.n242 B.n239 10.6151
R714 B.n239 B.n238 10.6151
R715 B.n238 B.n235 10.6151
R716 B.n235 B.n234 10.6151
R717 B.n231 B.n230 10.6151
R718 B.n230 B.n227 10.6151
R719 B.n227 B.n226 10.6151
R720 B.n226 B.n223 10.6151
R721 B.n223 B.n222 10.6151
R722 B.n222 B.n219 10.6151
R723 B.n219 B.n218 10.6151
R724 B.n218 B.n215 10.6151
R725 B.n215 B.n214 10.6151
R726 B.n211 B.n210 10.6151
R727 B.n210 B.n207 10.6151
R728 B.n207 B.n206 10.6151
R729 B.n206 B.n203 10.6151
R730 B.n203 B.n202 10.6151
R731 B.n202 B.n199 10.6151
R732 B.n199 B.n198 10.6151
R733 B.n198 B.n195 10.6151
R734 B.n195 B.n194 10.6151
R735 B.n194 B.n192 10.6151
R736 B.n255 B.n254 10.6151
R737 B.n255 B.n160 10.6151
R738 B.n266 B.n160 10.6151
R739 B.n267 B.n266 10.6151
R740 B.n268 B.n267 10.6151
R741 B.n268 B.n153 10.6151
R742 B.n278 B.n153 10.6151
R743 B.n279 B.n278 10.6151
R744 B.n280 B.n279 10.6151
R745 B.n280 B.n145 10.6151
R746 B.n289 B.n145 10.6151
R747 B.n290 B.n289 10.6151
R748 B.n291 B.n290 10.6151
R749 B.n291 B.n137 10.6151
R750 B.n302 B.n137 10.6151
R751 B.n303 B.n302 10.6151
R752 B.n304 B.n303 10.6151
R753 B.n304 B.n130 10.6151
R754 B.n315 B.n130 10.6151
R755 B.n316 B.n315 10.6151
R756 B.n317 B.n316 10.6151
R757 B.n317 B.n0 10.6151
R758 B.n399 B.n1 10.6151
R759 B.n399 B.n398 10.6151
R760 B.n398 B.n397 10.6151
R761 B.n397 B.n10 10.6151
R762 B.n391 B.n10 10.6151
R763 B.n391 B.n390 10.6151
R764 B.n390 B.n389 10.6151
R765 B.n389 B.n16 10.6151
R766 B.n383 B.n16 10.6151
R767 B.n383 B.n382 10.6151
R768 B.n382 B.n381 10.6151
R769 B.n381 B.n24 10.6151
R770 B.n376 B.n24 10.6151
R771 B.n376 B.n375 10.6151
R772 B.n375 B.n374 10.6151
R773 B.n374 B.n31 10.6151
R774 B.n368 B.n31 10.6151
R775 B.n368 B.n367 10.6151
R776 B.n367 B.n366 10.6151
R777 B.n366 B.n37 10.6151
R778 B.n360 B.n37 10.6151
R779 B.n360 B.n359 10.6151
R780 B.t5 B.n128 9.46287
R781 B.t7 B.n8 9.46287
R782 B.n85 B.n84 9.36635
R783 B.n107 B.n106 9.36635
R784 B.n234 B.n188 9.36635
R785 B.n211 B.n191 9.36635
R786 B.n306 B.t1 6.30874
R787 B.n393 B.t2 6.30874
R788 B.t3 B.n139 3.15462
R789 B.n386 B.t0 3.15462
R790 B.n405 B.n0 2.81026
R791 B.n405 B.n1 2.81026
R792 B.n86 B.n85 1.24928
R793 B.n106 B.n105 1.24928
R794 B.n231 B.n188 1.24928
R795 B.n214 B.n191 1.24928
R796 VP.n23 VP.n22 161.3
R797 VP.n8 VP.n7 161.3
R798 VP.n9 VP.n4 161.3
R799 VP.n10 VP.n3 161.3
R800 VP.n12 VP.n11 161.3
R801 VP.n21 VP.n0 161.3
R802 VP.n20 VP.n19 161.3
R803 VP.n18 VP.n1 161.3
R804 VP.n17 VP.n16 161.3
R805 VP.n15 VP.n2 161.3
R806 VP.n14 VP.n13 161.3
R807 VP.n6 VP.t1 139.417
R808 VP.n14 VP.t6 118.019
R809 VP.n16 VP.t5 118.019
R810 VP.n20 VP.t4 118.019
R811 VP.n22 VP.t3 118.019
R812 VP.n11 VP.t2 118.019
R813 VP.n9 VP.t7 118.019
R814 VP.n5 VP.t0 118.019
R815 VP.n7 VP.n6 44.853
R816 VP.n13 VP.n12 34.0687
R817 VP.n15 VP.n14 25.5611
R818 VP.n22 VP.n21 25.5611
R819 VP.n11 VP.n10 25.5611
R820 VP.n16 VP.n1 24.1005
R821 VP.n20 VP.n1 24.1005
R822 VP.n8 VP.n5 24.1005
R823 VP.n9 VP.n8 24.1005
R824 VP.n16 VP.n15 22.6399
R825 VP.n21 VP.n20 22.6399
R826 VP.n10 VP.n9 22.6399
R827 VP.n6 VP.n5 20.5405
R828 VP.n7 VP.n4 0.189894
R829 VP.n4 VP.n3 0.189894
R830 VP.n12 VP.n3 0.189894
R831 VP.n13 VP.n2 0.189894
R832 VP.n17 VP.n2 0.189894
R833 VP.n18 VP.n17 0.189894
R834 VP.n19 VP.n18 0.189894
R835 VP.n19 VP.n0 0.189894
R836 VP.n23 VP.n0 0.189894
R837 VP VP.n23 0.0516364
R838 VDD1 VDD1.n0 117.633
R839 VDD1.n3 VDD1.n2 117.519
R840 VDD1.n3 VDD1.n1 117.519
R841 VDD1.n5 VDD1.n4 117.139
R842 VDD1.n5 VDD1.n3 29.6819
R843 VDD1.n4 VDD1.t0 11.6476
R844 VDD1.n4 VDD1.t5 11.6476
R845 VDD1.n0 VDD1.t6 11.6476
R846 VDD1.n0 VDD1.t7 11.6476
R847 VDD1.n2 VDD1.t3 11.6476
R848 VDD1.n2 VDD1.t4 11.6476
R849 VDD1.n1 VDD1.t1 11.6476
R850 VDD1.n1 VDD1.t2 11.6476
R851 VDD1 VDD1.n5 0.377655
C0 VDD2 VDD1 0.812674f
C1 VP VDD2 0.322172f
C2 VTAIL VN 1.38357f
C3 VN VDD1 0.15423f
C4 VTAIL VDD1 3.39257f
C5 VP VN 3.41438f
C6 VTAIL VP 1.39767f
C7 VP VDD1 1.27622f
C8 VDD2 VN 1.10959f
C9 VTAIL VDD2 3.43411f
C10 VDD2 B 2.519791f
C11 VDD1 B 2.743768f
C12 VTAIL B 2.86132f
C13 VN B 6.620648f
C14 VP B 5.689229f
C15 VDD1.t6 B 0.025522f
C16 VDD1.t7 B 0.025522f
C17 VDD1.n0 B 0.148201f
C18 VDD1.t1 B 0.025522f
C19 VDD1.t2 B 0.025522f
C20 VDD1.n1 B 0.147956f
C21 VDD1.t3 B 0.025522f
C22 VDD1.t4 B 0.025522f
C23 VDD1.n2 B 0.147956f
C24 VDD1.n3 B 1.2001f
C25 VDD1.t0 B 0.025522f
C26 VDD1.t5 B 0.025522f
C27 VDD1.n4 B 0.147215f
C28 VDD1.n5 B 1.11693f
C29 VP.n0 B 0.027865f
C30 VP.n1 B 0.006323f
C31 VP.n2 B 0.027865f
C32 VP.n3 B 0.027865f
C33 VP.t2 B 0.101426f
C34 VP.t7 B 0.101426f
C35 VP.n4 B 0.027865f
C36 VP.t0 B 0.101426f
C37 VP.n5 B 0.078949f
C38 VP.t1 B 0.113127f
C39 VP.n6 B 0.067292f
C40 VP.n7 B 0.114516f
C41 VP.n8 B 0.006323f
C42 VP.n9 B 0.076778f
C43 VP.n10 B 0.006323f
C44 VP.n11 B 0.074287f
C45 VP.n12 B 0.787651f
C46 VP.n13 B 0.817138f
C47 VP.t6 B 0.101426f
C48 VP.n14 B 0.074287f
C49 VP.n15 B 0.006323f
C50 VP.t5 B 0.101426f
C51 VP.n16 B 0.076778f
C52 VP.n17 B 0.027865f
C53 VP.n18 B 0.027865f
C54 VP.n19 B 0.027865f
C55 VP.t4 B 0.101426f
C56 VP.n20 B 0.076778f
C57 VP.n21 B 0.006323f
C58 VP.t3 B 0.101426f
C59 VP.n22 B 0.074287f
C60 VP.n23 B 0.021595f
C61 VDD2.t6 B 0.02606f
C62 VDD2.t5 B 0.02606f
C63 VDD2.n0 B 0.151074f
C64 VDD2.t2 B 0.02606f
C65 VDD2.t3 B 0.02606f
C66 VDD2.n1 B 0.151074f
C67 VDD2.n2 B 1.18382f
C68 VDD2.t0 B 0.02606f
C69 VDD2.t7 B 0.02606f
C70 VDD2.n3 B 0.150317f
C71 VDD2.n4 B 1.11766f
C72 VDD2.t4 B 0.02606f
C73 VDD2.t1 B 0.02606f
C74 VDD2.n5 B 0.151064f
C75 VTAIL.t15 B 0.026628f
C76 VTAIL.t9 B 0.026628f
C77 VTAIL.n0 B 0.129279f
C78 VTAIL.n1 B 0.206912f
C79 VTAIL.t13 B 0.183691f
C80 VTAIL.n2 B 0.251412f
C81 VTAIL.t5 B 0.183691f
C82 VTAIL.n3 B 0.251412f
C83 VTAIL.t3 B 0.026628f
C84 VTAIL.t1 B 0.026628f
C85 VTAIL.n4 B 0.129279f
C86 VTAIL.n5 B 0.258805f
C87 VTAIL.t4 B 0.183691f
C88 VTAIL.n6 B 0.639866f
C89 VTAIL.t14 B 0.183692f
C90 VTAIL.n7 B 0.639866f
C91 VTAIL.t11 B 0.026628f
C92 VTAIL.t12 B 0.026628f
C93 VTAIL.n8 B 0.129279f
C94 VTAIL.n9 B 0.258805f
C95 VTAIL.t10 B 0.183692f
C96 VTAIL.n10 B 0.251411f
C97 VTAIL.t7 B 0.183692f
C98 VTAIL.n11 B 0.251411f
C99 VTAIL.t2 B 0.026628f
C100 VTAIL.t0 B 0.026628f
C101 VTAIL.n12 B 0.129279f
C102 VTAIL.n13 B 0.258805f
C103 VTAIL.t6 B 0.183692f
C104 VTAIL.n14 B 0.639866f
C105 VTAIL.t8 B 0.183691f
C106 VTAIL.n15 B 0.63615f
C107 VN.n0 B 0.027548f
C108 VN.n1 B 0.006251f
C109 VN.t1 B 0.111839f
C110 VN.t2 B 0.100271f
C111 VN.n2 B 0.07805f
C112 VN.n3 B 0.066526f
C113 VN.n4 B 0.113211f
C114 VN.n5 B 0.027548f
C115 VN.t5 B 0.100271f
C116 VN.n6 B 0.075904f
C117 VN.n7 B 0.006251f
C118 VN.t4 B 0.100271f
C119 VN.n8 B 0.073441f
C120 VN.n9 B 0.021349f
C121 VN.n10 B 0.027548f
C122 VN.n11 B 0.006251f
C123 VN.t0 B 0.100271f
C124 VN.t6 B 0.111839f
C125 VN.t3 B 0.100271f
C126 VN.n12 B 0.07805f
C127 VN.n13 B 0.066526f
C128 VN.n14 B 0.113211f
C129 VN.n15 B 0.027548f
C130 VN.n16 B 0.075904f
C131 VN.n17 B 0.006251f
C132 VN.t7 B 0.100271f
C133 VN.n18 B 0.073441f
C134 VN.n19 B 0.797029f
.ends

