* NGSPICE file created from diff_pair_sample_0157.ext - technology: sky130A

.subckt diff_pair_sample_0157 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X1 VDD1.t7 VP.t1 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=1.85
X2 VDD1.t2 VP.t2 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=1.85
X3 VTAIL.t3 VN.t0 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X4 VDD2.t8 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X5 VTAIL.t16 VP.t3 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X6 VDD1.t1 VP.t4 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=1.85
X7 VDD1.t6 VP.t5 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X8 VDD1.t5 VP.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X9 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=1.85
X10 VTAIL.t12 VP.t7 VDD1.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X11 VTAIL.t0 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X12 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=1.85
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=1.85
X14 VDD2.t6 VN.t3 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=1.85
X15 VDD1.t4 VP.t8 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=1.85
X16 VTAIL.t10 VP.t9 VDD1.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X17 VDD2.t5 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=1.85
X18 VDD2.t4 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X19 VDD2.t3 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=1.85
X20 VTAIL.t8 VN.t7 VDD2.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X21 VTAIL.t1 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=1.85
X22 VDD2.t0 VN.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=1.85
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=1.85
R0 VP.n42 VP.n9 180.482
R1 VP.n74 VP.n73 180.482
R2 VP.n41 VP.n40 180.482
R3 VP.n19 VP.n16 161.3
R4 VP.n21 VP.n20 161.3
R5 VP.n22 VP.n15 161.3
R6 VP.n24 VP.n23 161.3
R7 VP.n26 VP.n14 161.3
R8 VP.n28 VP.n27 161.3
R9 VP.n29 VP.n13 161.3
R10 VP.n31 VP.n30 161.3
R11 VP.n33 VP.n12 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n36 VP.n11 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n39 VP.n10 161.3
R16 VP.n72 VP.n0 161.3
R17 VP.n71 VP.n70 161.3
R18 VP.n69 VP.n1 161.3
R19 VP.n68 VP.n67 161.3
R20 VP.n66 VP.n2 161.3
R21 VP.n64 VP.n63 161.3
R22 VP.n62 VP.n3 161.3
R23 VP.n61 VP.n60 161.3
R24 VP.n59 VP.n4 161.3
R25 VP.n57 VP.n56 161.3
R26 VP.n55 VP.n5 161.3
R27 VP.n54 VP.n53 161.3
R28 VP.n52 VP.n6 161.3
R29 VP.n50 VP.n49 161.3
R30 VP.n48 VP.n7 161.3
R31 VP.n47 VP.n46 161.3
R32 VP.n45 VP.n8 161.3
R33 VP.n44 VP.n43 161.3
R34 VP.n17 VP.t2 92.324
R35 VP.n9 VP.t4 56.7983
R36 VP.n51 VP.t0 56.7983
R37 VP.n58 VP.t6 56.7983
R38 VP.n65 VP.t3 56.7983
R39 VP.n73 VP.t1 56.7983
R40 VP.n40 VP.t8 56.7983
R41 VP.n32 VP.t9 56.7983
R42 VP.n25 VP.t5 56.7983
R43 VP.n18 VP.t7 56.7983
R44 VP.n53 VP.n5 56.0773
R45 VP.n60 VP.n3 56.0773
R46 VP.n27 VP.n13 56.0773
R47 VP.n20 VP.n15 56.0773
R48 VP.n18 VP.n17 48.3759
R49 VP.n42 VP.n41 43.1899
R50 VP.n46 VP.n45 42.5146
R51 VP.n71 VP.n1 42.5146
R52 VP.n38 VP.n11 42.5146
R53 VP.n46 VP.n7 38.6395
R54 VP.n67 VP.n1 38.6395
R55 VP.n34 VP.n11 38.6395
R56 VP.n53 VP.n52 25.0767
R57 VP.n64 VP.n3 25.0767
R58 VP.n31 VP.n13 25.0767
R59 VP.n20 VP.n19 25.0767
R60 VP.n45 VP.n44 24.5923
R61 VP.n50 VP.n7 24.5923
R62 VP.n57 VP.n5 24.5923
R63 VP.n60 VP.n59 24.5923
R64 VP.n67 VP.n66 24.5923
R65 VP.n72 VP.n71 24.5923
R66 VP.n39 VP.n38 24.5923
R67 VP.n34 VP.n33 24.5923
R68 VP.n24 VP.n15 24.5923
R69 VP.n27 VP.n26 24.5923
R70 VP.n52 VP.n51 21.1495
R71 VP.n65 VP.n64 21.1495
R72 VP.n32 VP.n31 21.1495
R73 VP.n19 VP.n18 21.1495
R74 VP.n58 VP.n57 12.2964
R75 VP.n59 VP.n58 12.2964
R76 VP.n25 VP.n24 12.2964
R77 VP.n26 VP.n25 12.2964
R78 VP.n17 VP.n16 12.155
R79 VP.n44 VP.n9 5.4107
R80 VP.n73 VP.n72 5.4107
R81 VP.n40 VP.n39 5.4107
R82 VP.n51 VP.n50 3.44336
R83 VP.n66 VP.n65 3.44336
R84 VP.n33 VP.n32 3.44336
R85 VP.n21 VP.n16 0.189894
R86 VP.n22 VP.n21 0.189894
R87 VP.n23 VP.n22 0.189894
R88 VP.n23 VP.n14 0.189894
R89 VP.n28 VP.n14 0.189894
R90 VP.n29 VP.n28 0.189894
R91 VP.n30 VP.n29 0.189894
R92 VP.n30 VP.n12 0.189894
R93 VP.n35 VP.n12 0.189894
R94 VP.n36 VP.n35 0.189894
R95 VP.n37 VP.n36 0.189894
R96 VP.n37 VP.n10 0.189894
R97 VP.n41 VP.n10 0.189894
R98 VP.n43 VP.n42 0.189894
R99 VP.n43 VP.n8 0.189894
R100 VP.n47 VP.n8 0.189894
R101 VP.n48 VP.n47 0.189894
R102 VP.n49 VP.n48 0.189894
R103 VP.n49 VP.n6 0.189894
R104 VP.n54 VP.n6 0.189894
R105 VP.n55 VP.n54 0.189894
R106 VP.n56 VP.n55 0.189894
R107 VP.n56 VP.n4 0.189894
R108 VP.n61 VP.n4 0.189894
R109 VP.n62 VP.n61 0.189894
R110 VP.n63 VP.n62 0.189894
R111 VP.n63 VP.n2 0.189894
R112 VP.n68 VP.n2 0.189894
R113 VP.n69 VP.n68 0.189894
R114 VP.n70 VP.n69 0.189894
R115 VP.n70 VP.n0 0.189894
R116 VP.n74 VP.n0 0.189894
R117 VP VP.n74 0.0516364
R118 VDD1.n1 VDD1.t2 81.4421
R119 VDD1.n3 VDD1.t1 81.4418
R120 VDD1.n5 VDD1.n4 76.3754
R121 VDD1.n1 VDD1.n0 75.0215
R122 VDD1.n7 VDD1.n6 75.0213
R123 VDD1.n3 VDD1.n2 75.0213
R124 VDD1.n7 VDD1.n5 37.9233
R125 VDD1.n6 VDD1.t8 4.54178
R126 VDD1.n6 VDD1.t4 4.54178
R127 VDD1.n0 VDD1.t9 4.54178
R128 VDD1.n0 VDD1.t6 4.54178
R129 VDD1.n4 VDD1.t3 4.54178
R130 VDD1.n4 VDD1.t7 4.54178
R131 VDD1.n2 VDD1.t0 4.54178
R132 VDD1.n2 VDD1.t5 4.54178
R133 VDD1 VDD1.n7 1.35179
R134 VDD1 VDD1.n1 0.528517
R135 VDD1.n5 VDD1.n3 0.414982
R136 VTAIL.n11 VTAIL.t5 62.884
R137 VTAIL.n16 VTAIL.t11 62.8837
R138 VTAIL.n17 VTAIL.t7 62.8837
R139 VTAIL.n2 VTAIL.t18 62.8837
R140 VTAIL.n15 VTAIL.n14 58.3427
R141 VTAIL.n13 VTAIL.n12 58.3427
R142 VTAIL.n10 VTAIL.n9 58.3427
R143 VTAIL.n8 VTAIL.n7 58.3427
R144 VTAIL.n19 VTAIL.n18 58.3425
R145 VTAIL.n1 VTAIL.n0 58.3425
R146 VTAIL.n4 VTAIL.n3 58.3425
R147 VTAIL.n6 VTAIL.n5 58.3425
R148 VTAIL.n8 VTAIL.n6 19.8841
R149 VTAIL.n17 VTAIL.n16 18.0048
R150 VTAIL.n18 VTAIL.t2 4.54178
R151 VTAIL.n18 VTAIL.t3 4.54178
R152 VTAIL.n0 VTAIL.t4 4.54178
R153 VTAIL.n0 VTAIL.t1 4.54178
R154 VTAIL.n3 VTAIL.t13 4.54178
R155 VTAIL.n3 VTAIL.t16 4.54178
R156 VTAIL.n5 VTAIL.t15 4.54178
R157 VTAIL.n5 VTAIL.t19 4.54178
R158 VTAIL.n14 VTAIL.t14 4.54178
R159 VTAIL.n14 VTAIL.t10 4.54178
R160 VTAIL.n12 VTAIL.t17 4.54178
R161 VTAIL.n12 VTAIL.t12 4.54178
R162 VTAIL.n9 VTAIL.t6 4.54178
R163 VTAIL.n9 VTAIL.t8 4.54178
R164 VTAIL.n7 VTAIL.t9 4.54178
R165 VTAIL.n7 VTAIL.t0 4.54178
R166 VTAIL.n10 VTAIL.n8 1.87981
R167 VTAIL.n11 VTAIL.n10 1.87981
R168 VTAIL.n15 VTAIL.n13 1.87981
R169 VTAIL.n16 VTAIL.n15 1.87981
R170 VTAIL.n6 VTAIL.n4 1.87981
R171 VTAIL.n4 VTAIL.n2 1.87981
R172 VTAIL.n19 VTAIL.n17 1.87981
R173 VTAIL VTAIL.n1 1.46817
R174 VTAIL.n13 VTAIL.n11 1.40998
R175 VTAIL.n2 VTAIL.n1 1.40998
R176 VTAIL VTAIL.n19 0.412138
R177 B.n530 B.n529 585
R178 B.n532 B.n115 585
R179 B.n535 B.n534 585
R180 B.n536 B.n114 585
R181 B.n538 B.n537 585
R182 B.n540 B.n113 585
R183 B.n543 B.n542 585
R184 B.n544 B.n112 585
R185 B.n546 B.n545 585
R186 B.n548 B.n111 585
R187 B.n551 B.n550 585
R188 B.n552 B.n110 585
R189 B.n554 B.n553 585
R190 B.n556 B.n109 585
R191 B.n559 B.n558 585
R192 B.n560 B.n108 585
R193 B.n562 B.n561 585
R194 B.n564 B.n107 585
R195 B.n567 B.n566 585
R196 B.n569 B.n104 585
R197 B.n571 B.n570 585
R198 B.n573 B.n103 585
R199 B.n576 B.n575 585
R200 B.n577 B.n102 585
R201 B.n579 B.n578 585
R202 B.n581 B.n101 585
R203 B.n584 B.n583 585
R204 B.n585 B.n97 585
R205 B.n587 B.n586 585
R206 B.n589 B.n96 585
R207 B.n592 B.n591 585
R208 B.n593 B.n95 585
R209 B.n595 B.n594 585
R210 B.n597 B.n94 585
R211 B.n600 B.n599 585
R212 B.n601 B.n93 585
R213 B.n603 B.n602 585
R214 B.n605 B.n92 585
R215 B.n608 B.n607 585
R216 B.n609 B.n91 585
R217 B.n611 B.n610 585
R218 B.n613 B.n90 585
R219 B.n616 B.n615 585
R220 B.n617 B.n89 585
R221 B.n619 B.n618 585
R222 B.n621 B.n88 585
R223 B.n624 B.n623 585
R224 B.n625 B.n87 585
R225 B.n528 B.n85 585
R226 B.n628 B.n85 585
R227 B.n527 B.n84 585
R228 B.n629 B.n84 585
R229 B.n526 B.n83 585
R230 B.n630 B.n83 585
R231 B.n525 B.n524 585
R232 B.n524 B.n79 585
R233 B.n523 B.n78 585
R234 B.n636 B.n78 585
R235 B.n522 B.n77 585
R236 B.n637 B.n77 585
R237 B.n521 B.n76 585
R238 B.n638 B.n76 585
R239 B.n520 B.n519 585
R240 B.n519 B.n72 585
R241 B.n518 B.n71 585
R242 B.n644 B.n71 585
R243 B.n517 B.n70 585
R244 B.n645 B.n70 585
R245 B.n516 B.n69 585
R246 B.n646 B.n69 585
R247 B.n515 B.n514 585
R248 B.n514 B.n65 585
R249 B.n513 B.n64 585
R250 B.n652 B.n64 585
R251 B.n512 B.n63 585
R252 B.n653 B.n63 585
R253 B.n511 B.n62 585
R254 B.n654 B.n62 585
R255 B.n510 B.n509 585
R256 B.n509 B.n58 585
R257 B.n508 B.n57 585
R258 B.n660 B.n57 585
R259 B.n507 B.n56 585
R260 B.n661 B.n56 585
R261 B.n506 B.n55 585
R262 B.n662 B.n55 585
R263 B.n505 B.n504 585
R264 B.n504 B.n51 585
R265 B.n503 B.n50 585
R266 B.n668 B.n50 585
R267 B.n502 B.n49 585
R268 B.n669 B.n49 585
R269 B.n501 B.n48 585
R270 B.n670 B.n48 585
R271 B.n500 B.n499 585
R272 B.n499 B.n44 585
R273 B.n498 B.n43 585
R274 B.n676 B.n43 585
R275 B.n497 B.n42 585
R276 B.n677 B.n42 585
R277 B.n496 B.n41 585
R278 B.n678 B.n41 585
R279 B.n495 B.n494 585
R280 B.n494 B.n37 585
R281 B.n493 B.n36 585
R282 B.n684 B.n36 585
R283 B.n492 B.n35 585
R284 B.n685 B.n35 585
R285 B.n491 B.n34 585
R286 B.n686 B.n34 585
R287 B.n490 B.n489 585
R288 B.n489 B.n30 585
R289 B.n488 B.n29 585
R290 B.n692 B.n29 585
R291 B.n487 B.n28 585
R292 B.n693 B.n28 585
R293 B.n486 B.n27 585
R294 B.n694 B.n27 585
R295 B.n485 B.n484 585
R296 B.n484 B.n26 585
R297 B.n483 B.n22 585
R298 B.n700 B.n22 585
R299 B.n482 B.n21 585
R300 B.n701 B.n21 585
R301 B.n481 B.n20 585
R302 B.n702 B.n20 585
R303 B.n480 B.n479 585
R304 B.n479 B.n16 585
R305 B.n478 B.n15 585
R306 B.n708 B.n15 585
R307 B.n477 B.n14 585
R308 B.n709 B.n14 585
R309 B.n476 B.n13 585
R310 B.n710 B.n13 585
R311 B.n475 B.n474 585
R312 B.n474 B.n12 585
R313 B.n473 B.n472 585
R314 B.n473 B.n8 585
R315 B.n471 B.n7 585
R316 B.n717 B.n7 585
R317 B.n470 B.n6 585
R318 B.n718 B.n6 585
R319 B.n469 B.n5 585
R320 B.n719 B.n5 585
R321 B.n468 B.n467 585
R322 B.n467 B.n4 585
R323 B.n466 B.n116 585
R324 B.n466 B.n465 585
R325 B.n456 B.n117 585
R326 B.n118 B.n117 585
R327 B.n458 B.n457 585
R328 B.n459 B.n458 585
R329 B.n455 B.n122 585
R330 B.n126 B.n122 585
R331 B.n454 B.n453 585
R332 B.n453 B.n452 585
R333 B.n124 B.n123 585
R334 B.n125 B.n124 585
R335 B.n445 B.n444 585
R336 B.n446 B.n445 585
R337 B.n443 B.n131 585
R338 B.n131 B.n130 585
R339 B.n442 B.n441 585
R340 B.n441 B.n440 585
R341 B.n133 B.n132 585
R342 B.n433 B.n133 585
R343 B.n432 B.n431 585
R344 B.n434 B.n432 585
R345 B.n430 B.n138 585
R346 B.n138 B.n137 585
R347 B.n429 B.n428 585
R348 B.n428 B.n427 585
R349 B.n140 B.n139 585
R350 B.n141 B.n140 585
R351 B.n420 B.n419 585
R352 B.n421 B.n420 585
R353 B.n418 B.n146 585
R354 B.n146 B.n145 585
R355 B.n417 B.n416 585
R356 B.n416 B.n415 585
R357 B.n148 B.n147 585
R358 B.n149 B.n148 585
R359 B.n408 B.n407 585
R360 B.n409 B.n408 585
R361 B.n406 B.n154 585
R362 B.n154 B.n153 585
R363 B.n405 B.n404 585
R364 B.n404 B.n403 585
R365 B.n156 B.n155 585
R366 B.n157 B.n156 585
R367 B.n396 B.n395 585
R368 B.n397 B.n396 585
R369 B.n394 B.n162 585
R370 B.n162 B.n161 585
R371 B.n393 B.n392 585
R372 B.n392 B.n391 585
R373 B.n164 B.n163 585
R374 B.n165 B.n164 585
R375 B.n384 B.n383 585
R376 B.n385 B.n384 585
R377 B.n382 B.n170 585
R378 B.n170 B.n169 585
R379 B.n381 B.n380 585
R380 B.n380 B.n379 585
R381 B.n172 B.n171 585
R382 B.n173 B.n172 585
R383 B.n372 B.n371 585
R384 B.n373 B.n372 585
R385 B.n370 B.n178 585
R386 B.n178 B.n177 585
R387 B.n369 B.n368 585
R388 B.n368 B.n367 585
R389 B.n180 B.n179 585
R390 B.n181 B.n180 585
R391 B.n360 B.n359 585
R392 B.n361 B.n360 585
R393 B.n358 B.n186 585
R394 B.n186 B.n185 585
R395 B.n357 B.n356 585
R396 B.n356 B.n355 585
R397 B.n188 B.n187 585
R398 B.n189 B.n188 585
R399 B.n348 B.n347 585
R400 B.n349 B.n348 585
R401 B.n346 B.n194 585
R402 B.n194 B.n193 585
R403 B.n345 B.n344 585
R404 B.n344 B.n343 585
R405 B.n196 B.n195 585
R406 B.n197 B.n196 585
R407 B.n336 B.n335 585
R408 B.n337 B.n336 585
R409 B.n334 B.n202 585
R410 B.n202 B.n201 585
R411 B.n333 B.n332 585
R412 B.n332 B.n331 585
R413 B.n328 B.n206 585
R414 B.n327 B.n326 585
R415 B.n324 B.n207 585
R416 B.n324 B.n205 585
R417 B.n323 B.n322 585
R418 B.n321 B.n320 585
R419 B.n319 B.n209 585
R420 B.n317 B.n316 585
R421 B.n315 B.n210 585
R422 B.n314 B.n313 585
R423 B.n311 B.n211 585
R424 B.n309 B.n308 585
R425 B.n307 B.n212 585
R426 B.n306 B.n305 585
R427 B.n303 B.n213 585
R428 B.n301 B.n300 585
R429 B.n299 B.n214 585
R430 B.n298 B.n297 585
R431 B.n295 B.n215 585
R432 B.n293 B.n292 585
R433 B.n290 B.n216 585
R434 B.n289 B.n288 585
R435 B.n286 B.n219 585
R436 B.n284 B.n283 585
R437 B.n282 B.n220 585
R438 B.n281 B.n280 585
R439 B.n278 B.n221 585
R440 B.n276 B.n275 585
R441 B.n274 B.n222 585
R442 B.n273 B.n272 585
R443 B.n270 B.n269 585
R444 B.n268 B.n267 585
R445 B.n266 B.n227 585
R446 B.n264 B.n263 585
R447 B.n262 B.n228 585
R448 B.n261 B.n260 585
R449 B.n258 B.n229 585
R450 B.n256 B.n255 585
R451 B.n254 B.n230 585
R452 B.n253 B.n252 585
R453 B.n250 B.n231 585
R454 B.n248 B.n247 585
R455 B.n246 B.n232 585
R456 B.n245 B.n244 585
R457 B.n242 B.n233 585
R458 B.n240 B.n239 585
R459 B.n238 B.n234 585
R460 B.n237 B.n236 585
R461 B.n204 B.n203 585
R462 B.n205 B.n204 585
R463 B.n330 B.n329 585
R464 B.n331 B.n330 585
R465 B.n200 B.n199 585
R466 B.n201 B.n200 585
R467 B.n339 B.n338 585
R468 B.n338 B.n337 585
R469 B.n340 B.n198 585
R470 B.n198 B.n197 585
R471 B.n342 B.n341 585
R472 B.n343 B.n342 585
R473 B.n192 B.n191 585
R474 B.n193 B.n192 585
R475 B.n351 B.n350 585
R476 B.n350 B.n349 585
R477 B.n352 B.n190 585
R478 B.n190 B.n189 585
R479 B.n354 B.n353 585
R480 B.n355 B.n354 585
R481 B.n184 B.n183 585
R482 B.n185 B.n184 585
R483 B.n363 B.n362 585
R484 B.n362 B.n361 585
R485 B.n364 B.n182 585
R486 B.n182 B.n181 585
R487 B.n366 B.n365 585
R488 B.n367 B.n366 585
R489 B.n176 B.n175 585
R490 B.n177 B.n176 585
R491 B.n375 B.n374 585
R492 B.n374 B.n373 585
R493 B.n376 B.n174 585
R494 B.n174 B.n173 585
R495 B.n378 B.n377 585
R496 B.n379 B.n378 585
R497 B.n168 B.n167 585
R498 B.n169 B.n168 585
R499 B.n387 B.n386 585
R500 B.n386 B.n385 585
R501 B.n388 B.n166 585
R502 B.n166 B.n165 585
R503 B.n390 B.n389 585
R504 B.n391 B.n390 585
R505 B.n160 B.n159 585
R506 B.n161 B.n160 585
R507 B.n399 B.n398 585
R508 B.n398 B.n397 585
R509 B.n400 B.n158 585
R510 B.n158 B.n157 585
R511 B.n402 B.n401 585
R512 B.n403 B.n402 585
R513 B.n152 B.n151 585
R514 B.n153 B.n152 585
R515 B.n411 B.n410 585
R516 B.n410 B.n409 585
R517 B.n412 B.n150 585
R518 B.n150 B.n149 585
R519 B.n414 B.n413 585
R520 B.n415 B.n414 585
R521 B.n144 B.n143 585
R522 B.n145 B.n144 585
R523 B.n423 B.n422 585
R524 B.n422 B.n421 585
R525 B.n424 B.n142 585
R526 B.n142 B.n141 585
R527 B.n426 B.n425 585
R528 B.n427 B.n426 585
R529 B.n136 B.n135 585
R530 B.n137 B.n136 585
R531 B.n436 B.n435 585
R532 B.n435 B.n434 585
R533 B.n437 B.n134 585
R534 B.n433 B.n134 585
R535 B.n439 B.n438 585
R536 B.n440 B.n439 585
R537 B.n129 B.n128 585
R538 B.n130 B.n129 585
R539 B.n448 B.n447 585
R540 B.n447 B.n446 585
R541 B.n449 B.n127 585
R542 B.n127 B.n125 585
R543 B.n451 B.n450 585
R544 B.n452 B.n451 585
R545 B.n121 B.n120 585
R546 B.n126 B.n121 585
R547 B.n461 B.n460 585
R548 B.n460 B.n459 585
R549 B.n462 B.n119 585
R550 B.n119 B.n118 585
R551 B.n464 B.n463 585
R552 B.n465 B.n464 585
R553 B.n3 B.n0 585
R554 B.n4 B.n3 585
R555 B.n716 B.n1 585
R556 B.n717 B.n716 585
R557 B.n715 B.n714 585
R558 B.n715 B.n8 585
R559 B.n713 B.n9 585
R560 B.n12 B.n9 585
R561 B.n712 B.n711 585
R562 B.n711 B.n710 585
R563 B.n11 B.n10 585
R564 B.n709 B.n11 585
R565 B.n707 B.n706 585
R566 B.n708 B.n707 585
R567 B.n705 B.n17 585
R568 B.n17 B.n16 585
R569 B.n704 B.n703 585
R570 B.n703 B.n702 585
R571 B.n19 B.n18 585
R572 B.n701 B.n19 585
R573 B.n699 B.n698 585
R574 B.n700 B.n699 585
R575 B.n697 B.n23 585
R576 B.n26 B.n23 585
R577 B.n696 B.n695 585
R578 B.n695 B.n694 585
R579 B.n25 B.n24 585
R580 B.n693 B.n25 585
R581 B.n691 B.n690 585
R582 B.n692 B.n691 585
R583 B.n689 B.n31 585
R584 B.n31 B.n30 585
R585 B.n688 B.n687 585
R586 B.n687 B.n686 585
R587 B.n33 B.n32 585
R588 B.n685 B.n33 585
R589 B.n683 B.n682 585
R590 B.n684 B.n683 585
R591 B.n681 B.n38 585
R592 B.n38 B.n37 585
R593 B.n680 B.n679 585
R594 B.n679 B.n678 585
R595 B.n40 B.n39 585
R596 B.n677 B.n40 585
R597 B.n675 B.n674 585
R598 B.n676 B.n675 585
R599 B.n673 B.n45 585
R600 B.n45 B.n44 585
R601 B.n672 B.n671 585
R602 B.n671 B.n670 585
R603 B.n47 B.n46 585
R604 B.n669 B.n47 585
R605 B.n667 B.n666 585
R606 B.n668 B.n667 585
R607 B.n665 B.n52 585
R608 B.n52 B.n51 585
R609 B.n664 B.n663 585
R610 B.n663 B.n662 585
R611 B.n54 B.n53 585
R612 B.n661 B.n54 585
R613 B.n659 B.n658 585
R614 B.n660 B.n659 585
R615 B.n657 B.n59 585
R616 B.n59 B.n58 585
R617 B.n656 B.n655 585
R618 B.n655 B.n654 585
R619 B.n61 B.n60 585
R620 B.n653 B.n61 585
R621 B.n651 B.n650 585
R622 B.n652 B.n651 585
R623 B.n649 B.n66 585
R624 B.n66 B.n65 585
R625 B.n648 B.n647 585
R626 B.n647 B.n646 585
R627 B.n68 B.n67 585
R628 B.n645 B.n68 585
R629 B.n643 B.n642 585
R630 B.n644 B.n643 585
R631 B.n641 B.n73 585
R632 B.n73 B.n72 585
R633 B.n640 B.n639 585
R634 B.n639 B.n638 585
R635 B.n75 B.n74 585
R636 B.n637 B.n75 585
R637 B.n635 B.n634 585
R638 B.n636 B.n635 585
R639 B.n633 B.n80 585
R640 B.n80 B.n79 585
R641 B.n632 B.n631 585
R642 B.n631 B.n630 585
R643 B.n82 B.n81 585
R644 B.n629 B.n82 585
R645 B.n627 B.n626 585
R646 B.n628 B.n627 585
R647 B.n720 B.n719 585
R648 B.n718 B.n2 585
R649 B.n627 B.n87 502.111
R650 B.n530 B.n85 502.111
R651 B.n332 B.n204 502.111
R652 B.n330 B.n206 502.111
R653 B.n98 B.t14 263.341
R654 B.n105 B.t18 263.341
R655 B.n223 B.t21 263.341
R656 B.n217 B.t10 263.341
R657 B.n531 B.n86 256.663
R658 B.n533 B.n86 256.663
R659 B.n539 B.n86 256.663
R660 B.n541 B.n86 256.663
R661 B.n547 B.n86 256.663
R662 B.n549 B.n86 256.663
R663 B.n555 B.n86 256.663
R664 B.n557 B.n86 256.663
R665 B.n563 B.n86 256.663
R666 B.n565 B.n86 256.663
R667 B.n572 B.n86 256.663
R668 B.n574 B.n86 256.663
R669 B.n580 B.n86 256.663
R670 B.n582 B.n86 256.663
R671 B.n588 B.n86 256.663
R672 B.n590 B.n86 256.663
R673 B.n596 B.n86 256.663
R674 B.n598 B.n86 256.663
R675 B.n604 B.n86 256.663
R676 B.n606 B.n86 256.663
R677 B.n612 B.n86 256.663
R678 B.n614 B.n86 256.663
R679 B.n620 B.n86 256.663
R680 B.n622 B.n86 256.663
R681 B.n325 B.n205 256.663
R682 B.n208 B.n205 256.663
R683 B.n318 B.n205 256.663
R684 B.n312 B.n205 256.663
R685 B.n310 B.n205 256.663
R686 B.n304 B.n205 256.663
R687 B.n302 B.n205 256.663
R688 B.n296 B.n205 256.663
R689 B.n294 B.n205 256.663
R690 B.n287 B.n205 256.663
R691 B.n285 B.n205 256.663
R692 B.n279 B.n205 256.663
R693 B.n277 B.n205 256.663
R694 B.n271 B.n205 256.663
R695 B.n226 B.n205 256.663
R696 B.n265 B.n205 256.663
R697 B.n259 B.n205 256.663
R698 B.n257 B.n205 256.663
R699 B.n251 B.n205 256.663
R700 B.n249 B.n205 256.663
R701 B.n243 B.n205 256.663
R702 B.n241 B.n205 256.663
R703 B.n235 B.n205 256.663
R704 B.n722 B.n721 256.663
R705 B.n623 B.n621 163.367
R706 B.n619 B.n89 163.367
R707 B.n615 B.n613 163.367
R708 B.n611 B.n91 163.367
R709 B.n607 B.n605 163.367
R710 B.n603 B.n93 163.367
R711 B.n599 B.n597 163.367
R712 B.n595 B.n95 163.367
R713 B.n591 B.n589 163.367
R714 B.n587 B.n97 163.367
R715 B.n583 B.n581 163.367
R716 B.n579 B.n102 163.367
R717 B.n575 B.n573 163.367
R718 B.n571 B.n104 163.367
R719 B.n566 B.n564 163.367
R720 B.n562 B.n108 163.367
R721 B.n558 B.n556 163.367
R722 B.n554 B.n110 163.367
R723 B.n550 B.n548 163.367
R724 B.n546 B.n112 163.367
R725 B.n542 B.n540 163.367
R726 B.n538 B.n114 163.367
R727 B.n534 B.n532 163.367
R728 B.n332 B.n202 163.367
R729 B.n336 B.n202 163.367
R730 B.n336 B.n196 163.367
R731 B.n344 B.n196 163.367
R732 B.n344 B.n194 163.367
R733 B.n348 B.n194 163.367
R734 B.n348 B.n188 163.367
R735 B.n356 B.n188 163.367
R736 B.n356 B.n186 163.367
R737 B.n360 B.n186 163.367
R738 B.n360 B.n180 163.367
R739 B.n368 B.n180 163.367
R740 B.n368 B.n178 163.367
R741 B.n372 B.n178 163.367
R742 B.n372 B.n172 163.367
R743 B.n380 B.n172 163.367
R744 B.n380 B.n170 163.367
R745 B.n384 B.n170 163.367
R746 B.n384 B.n164 163.367
R747 B.n392 B.n164 163.367
R748 B.n392 B.n162 163.367
R749 B.n396 B.n162 163.367
R750 B.n396 B.n156 163.367
R751 B.n404 B.n156 163.367
R752 B.n404 B.n154 163.367
R753 B.n408 B.n154 163.367
R754 B.n408 B.n148 163.367
R755 B.n416 B.n148 163.367
R756 B.n416 B.n146 163.367
R757 B.n420 B.n146 163.367
R758 B.n420 B.n140 163.367
R759 B.n428 B.n140 163.367
R760 B.n428 B.n138 163.367
R761 B.n432 B.n138 163.367
R762 B.n432 B.n133 163.367
R763 B.n441 B.n133 163.367
R764 B.n441 B.n131 163.367
R765 B.n445 B.n131 163.367
R766 B.n445 B.n124 163.367
R767 B.n453 B.n124 163.367
R768 B.n453 B.n122 163.367
R769 B.n458 B.n122 163.367
R770 B.n458 B.n117 163.367
R771 B.n466 B.n117 163.367
R772 B.n467 B.n466 163.367
R773 B.n467 B.n5 163.367
R774 B.n6 B.n5 163.367
R775 B.n7 B.n6 163.367
R776 B.n473 B.n7 163.367
R777 B.n474 B.n473 163.367
R778 B.n474 B.n13 163.367
R779 B.n14 B.n13 163.367
R780 B.n15 B.n14 163.367
R781 B.n479 B.n15 163.367
R782 B.n479 B.n20 163.367
R783 B.n21 B.n20 163.367
R784 B.n22 B.n21 163.367
R785 B.n484 B.n22 163.367
R786 B.n484 B.n27 163.367
R787 B.n28 B.n27 163.367
R788 B.n29 B.n28 163.367
R789 B.n489 B.n29 163.367
R790 B.n489 B.n34 163.367
R791 B.n35 B.n34 163.367
R792 B.n36 B.n35 163.367
R793 B.n494 B.n36 163.367
R794 B.n494 B.n41 163.367
R795 B.n42 B.n41 163.367
R796 B.n43 B.n42 163.367
R797 B.n499 B.n43 163.367
R798 B.n499 B.n48 163.367
R799 B.n49 B.n48 163.367
R800 B.n50 B.n49 163.367
R801 B.n504 B.n50 163.367
R802 B.n504 B.n55 163.367
R803 B.n56 B.n55 163.367
R804 B.n57 B.n56 163.367
R805 B.n509 B.n57 163.367
R806 B.n509 B.n62 163.367
R807 B.n63 B.n62 163.367
R808 B.n64 B.n63 163.367
R809 B.n514 B.n64 163.367
R810 B.n514 B.n69 163.367
R811 B.n70 B.n69 163.367
R812 B.n71 B.n70 163.367
R813 B.n519 B.n71 163.367
R814 B.n519 B.n76 163.367
R815 B.n77 B.n76 163.367
R816 B.n78 B.n77 163.367
R817 B.n524 B.n78 163.367
R818 B.n524 B.n83 163.367
R819 B.n84 B.n83 163.367
R820 B.n85 B.n84 163.367
R821 B.n326 B.n324 163.367
R822 B.n324 B.n323 163.367
R823 B.n320 B.n319 163.367
R824 B.n317 B.n210 163.367
R825 B.n313 B.n311 163.367
R826 B.n309 B.n212 163.367
R827 B.n305 B.n303 163.367
R828 B.n301 B.n214 163.367
R829 B.n297 B.n295 163.367
R830 B.n293 B.n216 163.367
R831 B.n288 B.n286 163.367
R832 B.n284 B.n220 163.367
R833 B.n280 B.n278 163.367
R834 B.n276 B.n222 163.367
R835 B.n272 B.n270 163.367
R836 B.n267 B.n266 163.367
R837 B.n264 B.n228 163.367
R838 B.n260 B.n258 163.367
R839 B.n256 B.n230 163.367
R840 B.n252 B.n250 163.367
R841 B.n248 B.n232 163.367
R842 B.n244 B.n242 163.367
R843 B.n240 B.n234 163.367
R844 B.n236 B.n204 163.367
R845 B.n330 B.n200 163.367
R846 B.n338 B.n200 163.367
R847 B.n338 B.n198 163.367
R848 B.n342 B.n198 163.367
R849 B.n342 B.n192 163.367
R850 B.n350 B.n192 163.367
R851 B.n350 B.n190 163.367
R852 B.n354 B.n190 163.367
R853 B.n354 B.n184 163.367
R854 B.n362 B.n184 163.367
R855 B.n362 B.n182 163.367
R856 B.n366 B.n182 163.367
R857 B.n366 B.n176 163.367
R858 B.n374 B.n176 163.367
R859 B.n374 B.n174 163.367
R860 B.n378 B.n174 163.367
R861 B.n378 B.n168 163.367
R862 B.n386 B.n168 163.367
R863 B.n386 B.n166 163.367
R864 B.n390 B.n166 163.367
R865 B.n390 B.n160 163.367
R866 B.n398 B.n160 163.367
R867 B.n398 B.n158 163.367
R868 B.n402 B.n158 163.367
R869 B.n402 B.n152 163.367
R870 B.n410 B.n152 163.367
R871 B.n410 B.n150 163.367
R872 B.n414 B.n150 163.367
R873 B.n414 B.n144 163.367
R874 B.n422 B.n144 163.367
R875 B.n422 B.n142 163.367
R876 B.n426 B.n142 163.367
R877 B.n426 B.n136 163.367
R878 B.n435 B.n136 163.367
R879 B.n435 B.n134 163.367
R880 B.n439 B.n134 163.367
R881 B.n439 B.n129 163.367
R882 B.n447 B.n129 163.367
R883 B.n447 B.n127 163.367
R884 B.n451 B.n127 163.367
R885 B.n451 B.n121 163.367
R886 B.n460 B.n121 163.367
R887 B.n460 B.n119 163.367
R888 B.n464 B.n119 163.367
R889 B.n464 B.n3 163.367
R890 B.n720 B.n3 163.367
R891 B.n716 B.n2 163.367
R892 B.n716 B.n715 163.367
R893 B.n715 B.n9 163.367
R894 B.n711 B.n9 163.367
R895 B.n711 B.n11 163.367
R896 B.n707 B.n11 163.367
R897 B.n707 B.n17 163.367
R898 B.n703 B.n17 163.367
R899 B.n703 B.n19 163.367
R900 B.n699 B.n19 163.367
R901 B.n699 B.n23 163.367
R902 B.n695 B.n23 163.367
R903 B.n695 B.n25 163.367
R904 B.n691 B.n25 163.367
R905 B.n691 B.n31 163.367
R906 B.n687 B.n31 163.367
R907 B.n687 B.n33 163.367
R908 B.n683 B.n33 163.367
R909 B.n683 B.n38 163.367
R910 B.n679 B.n38 163.367
R911 B.n679 B.n40 163.367
R912 B.n675 B.n40 163.367
R913 B.n675 B.n45 163.367
R914 B.n671 B.n45 163.367
R915 B.n671 B.n47 163.367
R916 B.n667 B.n47 163.367
R917 B.n667 B.n52 163.367
R918 B.n663 B.n52 163.367
R919 B.n663 B.n54 163.367
R920 B.n659 B.n54 163.367
R921 B.n659 B.n59 163.367
R922 B.n655 B.n59 163.367
R923 B.n655 B.n61 163.367
R924 B.n651 B.n61 163.367
R925 B.n651 B.n66 163.367
R926 B.n647 B.n66 163.367
R927 B.n647 B.n68 163.367
R928 B.n643 B.n68 163.367
R929 B.n643 B.n73 163.367
R930 B.n639 B.n73 163.367
R931 B.n639 B.n75 163.367
R932 B.n635 B.n75 163.367
R933 B.n635 B.n80 163.367
R934 B.n631 B.n80 163.367
R935 B.n631 B.n82 163.367
R936 B.n627 B.n82 163.367
R937 B.n331 B.n205 147.276
R938 B.n628 B.n86 147.276
R939 B.n105 B.t19 118.665
R940 B.n223 B.t23 118.665
R941 B.n98 B.t16 118.662
R942 B.n217 B.t13 118.662
R943 B.n331 B.n201 77.6341
R944 B.n337 B.n201 77.6341
R945 B.n337 B.n197 77.6341
R946 B.n343 B.n197 77.6341
R947 B.n343 B.n193 77.6341
R948 B.n349 B.n193 77.6341
R949 B.n355 B.n189 77.6341
R950 B.n355 B.n185 77.6341
R951 B.n361 B.n185 77.6341
R952 B.n361 B.n181 77.6341
R953 B.n367 B.n181 77.6341
R954 B.n367 B.n177 77.6341
R955 B.n373 B.n177 77.6341
R956 B.n373 B.n173 77.6341
R957 B.n379 B.n173 77.6341
R958 B.n385 B.n169 77.6341
R959 B.n385 B.n165 77.6341
R960 B.n391 B.n165 77.6341
R961 B.n391 B.n161 77.6341
R962 B.n397 B.n161 77.6341
R963 B.n403 B.n157 77.6341
R964 B.n403 B.n153 77.6341
R965 B.n409 B.n153 77.6341
R966 B.n409 B.n149 77.6341
R967 B.n415 B.n149 77.6341
R968 B.n421 B.n145 77.6341
R969 B.n421 B.n141 77.6341
R970 B.n427 B.n141 77.6341
R971 B.n427 B.n137 77.6341
R972 B.n434 B.n137 77.6341
R973 B.n434 B.n433 77.6341
R974 B.n440 B.n130 77.6341
R975 B.n446 B.n130 77.6341
R976 B.n446 B.n125 77.6341
R977 B.n452 B.n125 77.6341
R978 B.n452 B.n126 77.6341
R979 B.n459 B.n118 77.6341
R980 B.n465 B.n118 77.6341
R981 B.n465 B.n4 77.6341
R982 B.n719 B.n4 77.6341
R983 B.n719 B.n718 77.6341
R984 B.n718 B.n717 77.6341
R985 B.n717 B.n8 77.6341
R986 B.n12 B.n8 77.6341
R987 B.n710 B.n12 77.6341
R988 B.n709 B.n708 77.6341
R989 B.n708 B.n16 77.6341
R990 B.n702 B.n16 77.6341
R991 B.n702 B.n701 77.6341
R992 B.n701 B.n700 77.6341
R993 B.n694 B.n26 77.6341
R994 B.n694 B.n693 77.6341
R995 B.n693 B.n692 77.6341
R996 B.n692 B.n30 77.6341
R997 B.n686 B.n30 77.6341
R998 B.n686 B.n685 77.6341
R999 B.n684 B.n37 77.6341
R1000 B.n678 B.n37 77.6341
R1001 B.n678 B.n677 77.6341
R1002 B.n677 B.n676 77.6341
R1003 B.n676 B.n44 77.6341
R1004 B.n670 B.n669 77.6341
R1005 B.n669 B.n668 77.6341
R1006 B.n668 B.n51 77.6341
R1007 B.n662 B.n51 77.6341
R1008 B.n662 B.n661 77.6341
R1009 B.n660 B.n58 77.6341
R1010 B.n654 B.n58 77.6341
R1011 B.n654 B.n653 77.6341
R1012 B.n653 B.n652 77.6341
R1013 B.n652 B.n65 77.6341
R1014 B.n646 B.n65 77.6341
R1015 B.n646 B.n645 77.6341
R1016 B.n645 B.n644 77.6341
R1017 B.n644 B.n72 77.6341
R1018 B.n638 B.n637 77.6341
R1019 B.n637 B.n636 77.6341
R1020 B.n636 B.n79 77.6341
R1021 B.n630 B.n79 77.6341
R1022 B.n630 B.n629 77.6341
R1023 B.n629 B.n628 77.6341
R1024 B.n106 B.t20 76.3861
R1025 B.n224 B.t22 76.3861
R1026 B.n99 B.t17 76.3822
R1027 B.n218 B.t12 76.3822
R1028 B.t9 B.n169 74.2091
R1029 B.n661 B.t7 74.2091
R1030 B.n622 B.n87 71.676
R1031 B.n621 B.n620 71.676
R1032 B.n614 B.n89 71.676
R1033 B.n613 B.n612 71.676
R1034 B.n606 B.n91 71.676
R1035 B.n605 B.n604 71.676
R1036 B.n598 B.n93 71.676
R1037 B.n597 B.n596 71.676
R1038 B.n590 B.n95 71.676
R1039 B.n589 B.n588 71.676
R1040 B.n582 B.n97 71.676
R1041 B.n581 B.n580 71.676
R1042 B.n574 B.n102 71.676
R1043 B.n573 B.n572 71.676
R1044 B.n565 B.n104 71.676
R1045 B.n564 B.n563 71.676
R1046 B.n557 B.n108 71.676
R1047 B.n556 B.n555 71.676
R1048 B.n549 B.n110 71.676
R1049 B.n548 B.n547 71.676
R1050 B.n541 B.n112 71.676
R1051 B.n540 B.n539 71.676
R1052 B.n533 B.n114 71.676
R1053 B.n532 B.n531 71.676
R1054 B.n531 B.n530 71.676
R1055 B.n534 B.n533 71.676
R1056 B.n539 B.n538 71.676
R1057 B.n542 B.n541 71.676
R1058 B.n547 B.n546 71.676
R1059 B.n550 B.n549 71.676
R1060 B.n555 B.n554 71.676
R1061 B.n558 B.n557 71.676
R1062 B.n563 B.n562 71.676
R1063 B.n566 B.n565 71.676
R1064 B.n572 B.n571 71.676
R1065 B.n575 B.n574 71.676
R1066 B.n580 B.n579 71.676
R1067 B.n583 B.n582 71.676
R1068 B.n588 B.n587 71.676
R1069 B.n591 B.n590 71.676
R1070 B.n596 B.n595 71.676
R1071 B.n599 B.n598 71.676
R1072 B.n604 B.n603 71.676
R1073 B.n607 B.n606 71.676
R1074 B.n612 B.n611 71.676
R1075 B.n615 B.n614 71.676
R1076 B.n620 B.n619 71.676
R1077 B.n623 B.n622 71.676
R1078 B.n325 B.n206 71.676
R1079 B.n323 B.n208 71.676
R1080 B.n319 B.n318 71.676
R1081 B.n312 B.n210 71.676
R1082 B.n311 B.n310 71.676
R1083 B.n304 B.n212 71.676
R1084 B.n303 B.n302 71.676
R1085 B.n296 B.n214 71.676
R1086 B.n295 B.n294 71.676
R1087 B.n287 B.n216 71.676
R1088 B.n286 B.n285 71.676
R1089 B.n279 B.n220 71.676
R1090 B.n278 B.n277 71.676
R1091 B.n271 B.n222 71.676
R1092 B.n270 B.n226 71.676
R1093 B.n266 B.n265 71.676
R1094 B.n259 B.n228 71.676
R1095 B.n258 B.n257 71.676
R1096 B.n251 B.n230 71.676
R1097 B.n250 B.n249 71.676
R1098 B.n243 B.n232 71.676
R1099 B.n242 B.n241 71.676
R1100 B.n235 B.n234 71.676
R1101 B.n326 B.n325 71.676
R1102 B.n320 B.n208 71.676
R1103 B.n318 B.n317 71.676
R1104 B.n313 B.n312 71.676
R1105 B.n310 B.n309 71.676
R1106 B.n305 B.n304 71.676
R1107 B.n302 B.n301 71.676
R1108 B.n297 B.n296 71.676
R1109 B.n294 B.n293 71.676
R1110 B.n288 B.n287 71.676
R1111 B.n285 B.n284 71.676
R1112 B.n280 B.n279 71.676
R1113 B.n277 B.n276 71.676
R1114 B.n272 B.n271 71.676
R1115 B.n267 B.n226 71.676
R1116 B.n265 B.n264 71.676
R1117 B.n260 B.n259 71.676
R1118 B.n257 B.n256 71.676
R1119 B.n252 B.n251 71.676
R1120 B.n249 B.n248 71.676
R1121 B.n244 B.n243 71.676
R1122 B.n241 B.n240 71.676
R1123 B.n236 B.n235 71.676
R1124 B.n721 B.n720 71.676
R1125 B.n721 B.n2 71.676
R1126 B.n415 B.t6 67.3591
R1127 B.t2 B.n684 67.3591
R1128 B.n100 B.n99 59.5399
R1129 B.n568 B.n106 59.5399
R1130 B.n225 B.n224 59.5399
R1131 B.n291 B.n218 59.5399
R1132 B.n440 B.t8 55.9424
R1133 B.n700 B.t1 55.9424
R1134 B.n126 B.t5 53.659
R1135 B.t4 B.n709 53.659
R1136 B.t11 B.n189 44.5257
R1137 B.t15 B.n72 44.5257
R1138 B.n99 B.n98 42.2793
R1139 B.n106 B.n105 42.2793
R1140 B.n224 B.n223 42.2793
R1141 B.n218 B.n217 42.2793
R1142 B.t0 B.n157 42.2423
R1143 B.t3 B.n44 42.2423
R1144 B.n397 B.t0 35.3923
R1145 B.n670 B.t3 35.3923
R1146 B.n349 B.t11 33.109
R1147 B.n638 B.t15 33.109
R1148 B.n329 B.n328 32.6249
R1149 B.n333 B.n203 32.6249
R1150 B.n529 B.n528 32.6249
R1151 B.n626 B.n625 32.6249
R1152 B.n459 B.t5 23.9756
R1153 B.n710 B.t4 23.9756
R1154 B.n433 B.t8 21.6922
R1155 B.n26 B.t1 21.6922
R1156 B B.n722 18.0485
R1157 B.n329 B.n199 10.6151
R1158 B.n339 B.n199 10.6151
R1159 B.n340 B.n339 10.6151
R1160 B.n341 B.n340 10.6151
R1161 B.n341 B.n191 10.6151
R1162 B.n351 B.n191 10.6151
R1163 B.n352 B.n351 10.6151
R1164 B.n353 B.n352 10.6151
R1165 B.n353 B.n183 10.6151
R1166 B.n363 B.n183 10.6151
R1167 B.n364 B.n363 10.6151
R1168 B.n365 B.n364 10.6151
R1169 B.n365 B.n175 10.6151
R1170 B.n375 B.n175 10.6151
R1171 B.n376 B.n375 10.6151
R1172 B.n377 B.n376 10.6151
R1173 B.n377 B.n167 10.6151
R1174 B.n387 B.n167 10.6151
R1175 B.n388 B.n387 10.6151
R1176 B.n389 B.n388 10.6151
R1177 B.n389 B.n159 10.6151
R1178 B.n399 B.n159 10.6151
R1179 B.n400 B.n399 10.6151
R1180 B.n401 B.n400 10.6151
R1181 B.n401 B.n151 10.6151
R1182 B.n411 B.n151 10.6151
R1183 B.n412 B.n411 10.6151
R1184 B.n413 B.n412 10.6151
R1185 B.n413 B.n143 10.6151
R1186 B.n423 B.n143 10.6151
R1187 B.n424 B.n423 10.6151
R1188 B.n425 B.n424 10.6151
R1189 B.n425 B.n135 10.6151
R1190 B.n436 B.n135 10.6151
R1191 B.n437 B.n436 10.6151
R1192 B.n438 B.n437 10.6151
R1193 B.n438 B.n128 10.6151
R1194 B.n448 B.n128 10.6151
R1195 B.n449 B.n448 10.6151
R1196 B.n450 B.n449 10.6151
R1197 B.n450 B.n120 10.6151
R1198 B.n461 B.n120 10.6151
R1199 B.n462 B.n461 10.6151
R1200 B.n463 B.n462 10.6151
R1201 B.n463 B.n0 10.6151
R1202 B.n328 B.n327 10.6151
R1203 B.n327 B.n207 10.6151
R1204 B.n322 B.n207 10.6151
R1205 B.n322 B.n321 10.6151
R1206 B.n321 B.n209 10.6151
R1207 B.n316 B.n209 10.6151
R1208 B.n316 B.n315 10.6151
R1209 B.n315 B.n314 10.6151
R1210 B.n314 B.n211 10.6151
R1211 B.n308 B.n211 10.6151
R1212 B.n308 B.n307 10.6151
R1213 B.n307 B.n306 10.6151
R1214 B.n306 B.n213 10.6151
R1215 B.n300 B.n213 10.6151
R1216 B.n300 B.n299 10.6151
R1217 B.n299 B.n298 10.6151
R1218 B.n298 B.n215 10.6151
R1219 B.n292 B.n215 10.6151
R1220 B.n290 B.n289 10.6151
R1221 B.n289 B.n219 10.6151
R1222 B.n283 B.n219 10.6151
R1223 B.n283 B.n282 10.6151
R1224 B.n282 B.n281 10.6151
R1225 B.n281 B.n221 10.6151
R1226 B.n275 B.n221 10.6151
R1227 B.n275 B.n274 10.6151
R1228 B.n274 B.n273 10.6151
R1229 B.n269 B.n268 10.6151
R1230 B.n268 B.n227 10.6151
R1231 B.n263 B.n227 10.6151
R1232 B.n263 B.n262 10.6151
R1233 B.n262 B.n261 10.6151
R1234 B.n261 B.n229 10.6151
R1235 B.n255 B.n229 10.6151
R1236 B.n255 B.n254 10.6151
R1237 B.n254 B.n253 10.6151
R1238 B.n253 B.n231 10.6151
R1239 B.n247 B.n231 10.6151
R1240 B.n247 B.n246 10.6151
R1241 B.n246 B.n245 10.6151
R1242 B.n245 B.n233 10.6151
R1243 B.n239 B.n233 10.6151
R1244 B.n239 B.n238 10.6151
R1245 B.n238 B.n237 10.6151
R1246 B.n237 B.n203 10.6151
R1247 B.n334 B.n333 10.6151
R1248 B.n335 B.n334 10.6151
R1249 B.n335 B.n195 10.6151
R1250 B.n345 B.n195 10.6151
R1251 B.n346 B.n345 10.6151
R1252 B.n347 B.n346 10.6151
R1253 B.n347 B.n187 10.6151
R1254 B.n357 B.n187 10.6151
R1255 B.n358 B.n357 10.6151
R1256 B.n359 B.n358 10.6151
R1257 B.n359 B.n179 10.6151
R1258 B.n369 B.n179 10.6151
R1259 B.n370 B.n369 10.6151
R1260 B.n371 B.n370 10.6151
R1261 B.n371 B.n171 10.6151
R1262 B.n381 B.n171 10.6151
R1263 B.n382 B.n381 10.6151
R1264 B.n383 B.n382 10.6151
R1265 B.n383 B.n163 10.6151
R1266 B.n393 B.n163 10.6151
R1267 B.n394 B.n393 10.6151
R1268 B.n395 B.n394 10.6151
R1269 B.n395 B.n155 10.6151
R1270 B.n405 B.n155 10.6151
R1271 B.n406 B.n405 10.6151
R1272 B.n407 B.n406 10.6151
R1273 B.n407 B.n147 10.6151
R1274 B.n417 B.n147 10.6151
R1275 B.n418 B.n417 10.6151
R1276 B.n419 B.n418 10.6151
R1277 B.n419 B.n139 10.6151
R1278 B.n429 B.n139 10.6151
R1279 B.n430 B.n429 10.6151
R1280 B.n431 B.n430 10.6151
R1281 B.n431 B.n132 10.6151
R1282 B.n442 B.n132 10.6151
R1283 B.n443 B.n442 10.6151
R1284 B.n444 B.n443 10.6151
R1285 B.n444 B.n123 10.6151
R1286 B.n454 B.n123 10.6151
R1287 B.n455 B.n454 10.6151
R1288 B.n457 B.n455 10.6151
R1289 B.n457 B.n456 10.6151
R1290 B.n456 B.n116 10.6151
R1291 B.n468 B.n116 10.6151
R1292 B.n469 B.n468 10.6151
R1293 B.n470 B.n469 10.6151
R1294 B.n471 B.n470 10.6151
R1295 B.n472 B.n471 10.6151
R1296 B.n475 B.n472 10.6151
R1297 B.n476 B.n475 10.6151
R1298 B.n477 B.n476 10.6151
R1299 B.n478 B.n477 10.6151
R1300 B.n480 B.n478 10.6151
R1301 B.n481 B.n480 10.6151
R1302 B.n482 B.n481 10.6151
R1303 B.n483 B.n482 10.6151
R1304 B.n485 B.n483 10.6151
R1305 B.n486 B.n485 10.6151
R1306 B.n487 B.n486 10.6151
R1307 B.n488 B.n487 10.6151
R1308 B.n490 B.n488 10.6151
R1309 B.n491 B.n490 10.6151
R1310 B.n492 B.n491 10.6151
R1311 B.n493 B.n492 10.6151
R1312 B.n495 B.n493 10.6151
R1313 B.n496 B.n495 10.6151
R1314 B.n497 B.n496 10.6151
R1315 B.n498 B.n497 10.6151
R1316 B.n500 B.n498 10.6151
R1317 B.n501 B.n500 10.6151
R1318 B.n502 B.n501 10.6151
R1319 B.n503 B.n502 10.6151
R1320 B.n505 B.n503 10.6151
R1321 B.n506 B.n505 10.6151
R1322 B.n507 B.n506 10.6151
R1323 B.n508 B.n507 10.6151
R1324 B.n510 B.n508 10.6151
R1325 B.n511 B.n510 10.6151
R1326 B.n512 B.n511 10.6151
R1327 B.n513 B.n512 10.6151
R1328 B.n515 B.n513 10.6151
R1329 B.n516 B.n515 10.6151
R1330 B.n517 B.n516 10.6151
R1331 B.n518 B.n517 10.6151
R1332 B.n520 B.n518 10.6151
R1333 B.n521 B.n520 10.6151
R1334 B.n522 B.n521 10.6151
R1335 B.n523 B.n522 10.6151
R1336 B.n525 B.n523 10.6151
R1337 B.n526 B.n525 10.6151
R1338 B.n527 B.n526 10.6151
R1339 B.n528 B.n527 10.6151
R1340 B.n714 B.n1 10.6151
R1341 B.n714 B.n713 10.6151
R1342 B.n713 B.n712 10.6151
R1343 B.n712 B.n10 10.6151
R1344 B.n706 B.n10 10.6151
R1345 B.n706 B.n705 10.6151
R1346 B.n705 B.n704 10.6151
R1347 B.n704 B.n18 10.6151
R1348 B.n698 B.n18 10.6151
R1349 B.n698 B.n697 10.6151
R1350 B.n697 B.n696 10.6151
R1351 B.n696 B.n24 10.6151
R1352 B.n690 B.n24 10.6151
R1353 B.n690 B.n689 10.6151
R1354 B.n689 B.n688 10.6151
R1355 B.n688 B.n32 10.6151
R1356 B.n682 B.n32 10.6151
R1357 B.n682 B.n681 10.6151
R1358 B.n681 B.n680 10.6151
R1359 B.n680 B.n39 10.6151
R1360 B.n674 B.n39 10.6151
R1361 B.n674 B.n673 10.6151
R1362 B.n673 B.n672 10.6151
R1363 B.n672 B.n46 10.6151
R1364 B.n666 B.n46 10.6151
R1365 B.n666 B.n665 10.6151
R1366 B.n665 B.n664 10.6151
R1367 B.n664 B.n53 10.6151
R1368 B.n658 B.n53 10.6151
R1369 B.n658 B.n657 10.6151
R1370 B.n657 B.n656 10.6151
R1371 B.n656 B.n60 10.6151
R1372 B.n650 B.n60 10.6151
R1373 B.n650 B.n649 10.6151
R1374 B.n649 B.n648 10.6151
R1375 B.n648 B.n67 10.6151
R1376 B.n642 B.n67 10.6151
R1377 B.n642 B.n641 10.6151
R1378 B.n641 B.n640 10.6151
R1379 B.n640 B.n74 10.6151
R1380 B.n634 B.n74 10.6151
R1381 B.n634 B.n633 10.6151
R1382 B.n633 B.n632 10.6151
R1383 B.n632 B.n81 10.6151
R1384 B.n626 B.n81 10.6151
R1385 B.n625 B.n624 10.6151
R1386 B.n624 B.n88 10.6151
R1387 B.n618 B.n88 10.6151
R1388 B.n618 B.n617 10.6151
R1389 B.n617 B.n616 10.6151
R1390 B.n616 B.n90 10.6151
R1391 B.n610 B.n90 10.6151
R1392 B.n610 B.n609 10.6151
R1393 B.n609 B.n608 10.6151
R1394 B.n608 B.n92 10.6151
R1395 B.n602 B.n92 10.6151
R1396 B.n602 B.n601 10.6151
R1397 B.n601 B.n600 10.6151
R1398 B.n600 B.n94 10.6151
R1399 B.n594 B.n94 10.6151
R1400 B.n594 B.n593 10.6151
R1401 B.n593 B.n592 10.6151
R1402 B.n592 B.n96 10.6151
R1403 B.n586 B.n585 10.6151
R1404 B.n585 B.n584 10.6151
R1405 B.n584 B.n101 10.6151
R1406 B.n578 B.n101 10.6151
R1407 B.n578 B.n577 10.6151
R1408 B.n577 B.n576 10.6151
R1409 B.n576 B.n103 10.6151
R1410 B.n570 B.n103 10.6151
R1411 B.n570 B.n569 10.6151
R1412 B.n567 B.n107 10.6151
R1413 B.n561 B.n107 10.6151
R1414 B.n561 B.n560 10.6151
R1415 B.n560 B.n559 10.6151
R1416 B.n559 B.n109 10.6151
R1417 B.n553 B.n109 10.6151
R1418 B.n553 B.n552 10.6151
R1419 B.n552 B.n551 10.6151
R1420 B.n551 B.n111 10.6151
R1421 B.n545 B.n111 10.6151
R1422 B.n545 B.n544 10.6151
R1423 B.n544 B.n543 10.6151
R1424 B.n543 B.n113 10.6151
R1425 B.n537 B.n113 10.6151
R1426 B.n537 B.n536 10.6151
R1427 B.n536 B.n535 10.6151
R1428 B.n535 B.n115 10.6151
R1429 B.n529 B.n115 10.6151
R1430 B.t6 B.n145 10.2755
R1431 B.n685 B.t2 10.2755
R1432 B.n292 B.n291 9.36635
R1433 B.n269 B.n225 9.36635
R1434 B.n100 B.n96 9.36635
R1435 B.n568 B.n567 9.36635
R1436 B.n722 B.n0 8.11757
R1437 B.n722 B.n1 8.11757
R1438 B.n379 B.t9 3.42551
R1439 B.t7 B.n660 3.42551
R1440 B.n291 B.n290 1.24928
R1441 B.n273 B.n225 1.24928
R1442 B.n586 B.n100 1.24928
R1443 B.n569 B.n568 1.24928
R1444 VN.n31 VN.n30 180.482
R1445 VN.n63 VN.n62 180.482
R1446 VN.n61 VN.n32 161.3
R1447 VN.n60 VN.n59 161.3
R1448 VN.n58 VN.n33 161.3
R1449 VN.n57 VN.n56 161.3
R1450 VN.n55 VN.n34 161.3
R1451 VN.n53 VN.n52 161.3
R1452 VN.n51 VN.n35 161.3
R1453 VN.n50 VN.n49 161.3
R1454 VN.n48 VN.n36 161.3
R1455 VN.n46 VN.n45 161.3
R1456 VN.n44 VN.n37 161.3
R1457 VN.n43 VN.n42 161.3
R1458 VN.n41 VN.n38 161.3
R1459 VN.n29 VN.n0 161.3
R1460 VN.n28 VN.n27 161.3
R1461 VN.n26 VN.n1 161.3
R1462 VN.n25 VN.n24 161.3
R1463 VN.n23 VN.n2 161.3
R1464 VN.n21 VN.n20 161.3
R1465 VN.n19 VN.n3 161.3
R1466 VN.n18 VN.n17 161.3
R1467 VN.n16 VN.n4 161.3
R1468 VN.n14 VN.n13 161.3
R1469 VN.n12 VN.n5 161.3
R1470 VN.n11 VN.n10 161.3
R1471 VN.n9 VN.n6 161.3
R1472 VN.n7 VN.t6 92.324
R1473 VN.n39 VN.t4 92.324
R1474 VN.n8 VN.t8 56.7983
R1475 VN.n15 VN.t5 56.7983
R1476 VN.n22 VN.t0 56.7983
R1477 VN.n30 VN.t9 56.7983
R1478 VN.n40 VN.t7 56.7983
R1479 VN.n47 VN.t1 56.7983
R1480 VN.n54 VN.t2 56.7983
R1481 VN.n62 VN.t3 56.7983
R1482 VN.n10 VN.n5 56.0773
R1483 VN.n17 VN.n3 56.0773
R1484 VN.n42 VN.n37 56.0773
R1485 VN.n49 VN.n35 56.0773
R1486 VN.n8 VN.n7 48.3759
R1487 VN.n40 VN.n39 48.3759
R1488 VN VN.n63 43.5706
R1489 VN.n28 VN.n1 42.5146
R1490 VN.n60 VN.n33 42.5146
R1491 VN.n24 VN.n1 38.6395
R1492 VN.n56 VN.n33 38.6395
R1493 VN.n10 VN.n9 25.0767
R1494 VN.n21 VN.n3 25.0767
R1495 VN.n42 VN.n41 25.0767
R1496 VN.n53 VN.n35 25.0767
R1497 VN.n14 VN.n5 24.5923
R1498 VN.n17 VN.n16 24.5923
R1499 VN.n24 VN.n23 24.5923
R1500 VN.n29 VN.n28 24.5923
R1501 VN.n49 VN.n48 24.5923
R1502 VN.n46 VN.n37 24.5923
R1503 VN.n56 VN.n55 24.5923
R1504 VN.n61 VN.n60 24.5923
R1505 VN.n9 VN.n8 21.1495
R1506 VN.n22 VN.n21 21.1495
R1507 VN.n41 VN.n40 21.1495
R1508 VN.n54 VN.n53 21.1495
R1509 VN.n15 VN.n14 12.2964
R1510 VN.n16 VN.n15 12.2964
R1511 VN.n48 VN.n47 12.2964
R1512 VN.n47 VN.n46 12.2964
R1513 VN.n39 VN.n38 12.155
R1514 VN.n7 VN.n6 12.155
R1515 VN.n30 VN.n29 5.4107
R1516 VN.n62 VN.n61 5.4107
R1517 VN.n23 VN.n22 3.44336
R1518 VN.n55 VN.n54 3.44336
R1519 VN.n63 VN.n32 0.189894
R1520 VN.n59 VN.n32 0.189894
R1521 VN.n59 VN.n58 0.189894
R1522 VN.n58 VN.n57 0.189894
R1523 VN.n57 VN.n34 0.189894
R1524 VN.n52 VN.n34 0.189894
R1525 VN.n52 VN.n51 0.189894
R1526 VN.n51 VN.n50 0.189894
R1527 VN.n50 VN.n36 0.189894
R1528 VN.n45 VN.n36 0.189894
R1529 VN.n45 VN.n44 0.189894
R1530 VN.n44 VN.n43 0.189894
R1531 VN.n43 VN.n38 0.189894
R1532 VN.n11 VN.n6 0.189894
R1533 VN.n12 VN.n11 0.189894
R1534 VN.n13 VN.n12 0.189894
R1535 VN.n13 VN.n4 0.189894
R1536 VN.n18 VN.n4 0.189894
R1537 VN.n19 VN.n18 0.189894
R1538 VN.n20 VN.n19 0.189894
R1539 VN.n20 VN.n2 0.189894
R1540 VN.n25 VN.n2 0.189894
R1541 VN.n26 VN.n25 0.189894
R1542 VN.n27 VN.n26 0.189894
R1543 VN.n27 VN.n0 0.189894
R1544 VN.n31 VN.n0 0.189894
R1545 VN VN.n31 0.0516364
R1546 VDD2.n1 VDD2.t3 81.4418
R1547 VDD2.n4 VDD2.t6 79.5627
R1548 VDD2.n3 VDD2.n2 76.3754
R1549 VDD2 VDD2.n7 76.3726
R1550 VDD2.n6 VDD2.n5 75.0215
R1551 VDD2.n1 VDD2.n0 75.0213
R1552 VDD2.n4 VDD2.n3 36.4006
R1553 VDD2.n7 VDD2.t2 4.54178
R1554 VDD2.n7 VDD2.t5 4.54178
R1555 VDD2.n5 VDD2.t7 4.54178
R1556 VDD2.n5 VDD2.t8 4.54178
R1557 VDD2.n2 VDD2.t9 4.54178
R1558 VDD2.n2 VDD2.t0 4.54178
R1559 VDD2.n0 VDD2.t1 4.54178
R1560 VDD2.n0 VDD2.t4 4.54178
R1561 VDD2.n6 VDD2.n4 1.87981
R1562 VDD2 VDD2.n6 0.528517
R1563 VDD2.n3 VDD2.n1 0.414982
C0 VTAIL VDD1 6.32393f
C1 VDD1 VDD2 1.6844f
C2 VDD1 VP 4.230259f
C3 VTAIL VN 4.72027f
C4 VDD2 VN 3.89707f
C5 VN VP 5.87513f
C6 VDD1 VN 0.15596f
C7 VTAIL VDD2 6.37123f
C8 VTAIL VP 4.73447f
C9 VDD2 VP 0.491999f
C10 VDD2 B 4.952646f
C11 VDD1 B 4.931407f
C12 VTAIL B 4.281471f
C13 VN B 13.78623f
C14 VP B 12.301999f
C15 VDD2.t3 B 0.809403f
C16 VDD2.t1 B 0.078947f
C17 VDD2.t4 B 0.078947f
C18 VDD2.n0 B 0.629206f
C19 VDD2.n1 B 0.714332f
C20 VDD2.t9 B 0.078947f
C21 VDD2.t0 B 0.078947f
C22 VDD2.n2 B 0.636806f
C23 VDD2.n3 B 1.87559f
C24 VDD2.t6 B 0.800822f
C25 VDD2.n4 B 2.019f
C26 VDD2.t7 B 0.078947f
C27 VDD2.t8 B 0.078947f
C28 VDD2.n5 B 0.629208f
C29 VDD2.n6 B 0.358036f
C30 VDD2.t2 B 0.078947f
C31 VDD2.t5 B 0.078947f
C32 VDD2.n7 B 0.636779f
C33 VN.n0 B 0.029993f
C34 VN.t9 B 0.626151f
C35 VN.n1 B 0.024378f
C36 VN.n2 B 0.029993f
C37 VN.t0 B 0.626151f
C38 VN.n3 B 0.035685f
C39 VN.n4 B 0.029993f
C40 VN.t5 B 0.626151f
C41 VN.n5 B 0.050994f
C42 VN.n6 B 0.222804f
C43 VN.t8 B 0.626151f
C44 VN.t6 B 0.779476f
C45 VN.n7 B 0.310343f
C46 VN.n8 B 0.330833f
C47 VN.n9 B 0.052295f
C48 VN.n10 B 0.035685f
C49 VN.n11 B 0.029993f
C50 VN.n12 B 0.029993f
C51 VN.n13 B 0.029993f
C52 VN.n14 B 0.04189f
C53 VN.n15 B 0.253453f
C54 VN.n16 B 0.04189f
C55 VN.n17 B 0.050994f
C56 VN.n18 B 0.029993f
C57 VN.n19 B 0.029993f
C58 VN.n20 B 0.029993f
C59 VN.n21 B 0.052295f
C60 VN.n22 B 0.253453f
C61 VN.n23 B 0.032006f
C62 VN.n24 B 0.059812f
C63 VN.n25 B 0.029993f
C64 VN.n26 B 0.029993f
C65 VN.n27 B 0.029993f
C66 VN.n28 B 0.058629f
C67 VN.n29 B 0.034202f
C68 VN.n30 B 0.325737f
C69 VN.n31 B 0.03184f
C70 VN.n32 B 0.029993f
C71 VN.t3 B 0.626151f
C72 VN.n33 B 0.024378f
C73 VN.n34 B 0.029993f
C74 VN.t2 B 0.626151f
C75 VN.n35 B 0.035685f
C76 VN.n36 B 0.029993f
C77 VN.t1 B 0.626151f
C78 VN.n37 B 0.050994f
C79 VN.n38 B 0.222804f
C80 VN.t7 B 0.626151f
C81 VN.t4 B 0.779476f
C82 VN.n39 B 0.310343f
C83 VN.n40 B 0.330833f
C84 VN.n41 B 0.052295f
C85 VN.n42 B 0.035685f
C86 VN.n43 B 0.029993f
C87 VN.n44 B 0.029993f
C88 VN.n45 B 0.029993f
C89 VN.n46 B 0.04189f
C90 VN.n47 B 0.253453f
C91 VN.n48 B 0.04189f
C92 VN.n49 B 0.050994f
C93 VN.n50 B 0.029993f
C94 VN.n51 B 0.029993f
C95 VN.n52 B 0.029993f
C96 VN.n53 B 0.052295f
C97 VN.n54 B 0.253453f
C98 VN.n55 B 0.032006f
C99 VN.n56 B 0.059812f
C100 VN.n57 B 0.029993f
C101 VN.n58 B 0.029993f
C102 VN.n59 B 0.029993f
C103 VN.n60 B 0.058629f
C104 VN.n61 B 0.034202f
C105 VN.n62 B 0.325737f
C106 VN.n63 B 1.32468f
C107 VTAIL.t4 B 0.100918f
C108 VTAIL.t1 B 0.100918f
C109 VTAIL.n0 B 0.740017f
C110 VTAIL.n1 B 0.526501f
C111 VTAIL.t18 B 0.949217f
C112 VTAIL.n2 B 0.631383f
C113 VTAIL.t13 B 0.100918f
C114 VTAIL.t16 B 0.100918f
C115 VTAIL.n3 B 0.740017f
C116 VTAIL.n4 B 0.609695f
C117 VTAIL.t15 B 0.100918f
C118 VTAIL.t19 B 0.100918f
C119 VTAIL.n5 B 0.740017f
C120 VTAIL.n6 B 1.53969f
C121 VTAIL.t9 B 0.100918f
C122 VTAIL.t0 B 0.100918f
C123 VTAIL.n7 B 0.740021f
C124 VTAIL.n8 B 1.53968f
C125 VTAIL.t6 B 0.100918f
C126 VTAIL.t8 B 0.100918f
C127 VTAIL.n9 B 0.740021f
C128 VTAIL.n10 B 0.609691f
C129 VTAIL.t5 B 0.949221f
C130 VTAIL.n11 B 0.631379f
C131 VTAIL.t17 B 0.100918f
C132 VTAIL.t12 B 0.100918f
C133 VTAIL.n12 B 0.740021f
C134 VTAIL.n13 B 0.565348f
C135 VTAIL.t14 B 0.100918f
C136 VTAIL.t10 B 0.100918f
C137 VTAIL.n14 B 0.740021f
C138 VTAIL.n15 B 0.609691f
C139 VTAIL.t11 B 0.949217f
C140 VTAIL.n16 B 1.42835f
C141 VTAIL.t7 B 0.949217f
C142 VTAIL.n17 B 1.42835f
C143 VTAIL.t2 B 0.100918f
C144 VTAIL.t3 B 0.100918f
C145 VTAIL.n18 B 0.740017f
C146 VTAIL.n19 B 0.471174f
C147 VDD1.t2 B 0.818397f
C148 VDD1.t9 B 0.079825f
C149 VDD1.t6 B 0.079825f
C150 VDD1.n0 B 0.636198f
C151 VDD1.n1 B 0.729444f
C152 VDD1.t1 B 0.818396f
C153 VDD1.t0 B 0.079825f
C154 VDD1.t5 B 0.079825f
C155 VDD1.n2 B 0.636196f
C156 VDD1.n3 B 0.722268f
C157 VDD1.t3 B 0.079825f
C158 VDD1.t7 B 0.079825f
C159 VDD1.n4 B 0.643881f
C160 VDD1.n5 B 1.98885f
C161 VDD1.t8 B 0.079825f
C162 VDD1.t4 B 0.079825f
C163 VDD1.n6 B 0.636195f
C164 VDD1.n7 B 2.09128f
C165 VP.n0 B 0.030703f
C166 VP.t1 B 0.64097f
C167 VP.n1 B 0.024955f
C168 VP.n2 B 0.030703f
C169 VP.t3 B 0.64097f
C170 VP.n3 B 0.03653f
C171 VP.n4 B 0.030703f
C172 VP.t6 B 0.64097f
C173 VP.n5 B 0.052201f
C174 VP.n6 B 0.030703f
C175 VP.t0 B 0.64097f
C176 VP.n7 B 0.061228f
C177 VP.n8 B 0.030703f
C178 VP.t4 B 0.64097f
C179 VP.n9 B 0.333446f
C180 VP.n10 B 0.030703f
C181 VP.t8 B 0.64097f
C182 VP.n11 B 0.024955f
C183 VP.n12 B 0.030703f
C184 VP.t9 B 0.64097f
C185 VP.n13 B 0.03653f
C186 VP.n14 B 0.030703f
C187 VP.t5 B 0.64097f
C188 VP.n15 B 0.052201f
C189 VP.n16 B 0.228077f
C190 VP.t7 B 0.64097f
C191 VP.t2 B 0.797923f
C192 VP.n17 B 0.317688f
C193 VP.n18 B 0.338663f
C194 VP.n19 B 0.053533f
C195 VP.n20 B 0.03653f
C196 VP.n21 B 0.030703f
C197 VP.n22 B 0.030703f
C198 VP.n23 B 0.030703f
C199 VP.n24 B 0.042882f
C200 VP.n25 B 0.259451f
C201 VP.n26 B 0.042882f
C202 VP.n27 B 0.052201f
C203 VP.n28 B 0.030703f
C204 VP.n29 B 0.030703f
C205 VP.n30 B 0.030703f
C206 VP.n31 B 0.053533f
C207 VP.n32 B 0.259451f
C208 VP.n33 B 0.032763f
C209 VP.n34 B 0.061228f
C210 VP.n35 B 0.030703f
C211 VP.n36 B 0.030703f
C212 VP.n37 B 0.030703f
C213 VP.n38 B 0.060016f
C214 VP.n39 B 0.035012f
C215 VP.n40 B 0.333446f
C216 VP.n41 B 1.33591f
C217 VP.n42 B 1.36154f
C218 VP.n43 B 0.030703f
C219 VP.n44 B 0.035012f
C220 VP.n45 B 0.060016f
C221 VP.n46 B 0.024955f
C222 VP.n47 B 0.030703f
C223 VP.n48 B 0.030703f
C224 VP.n49 B 0.030703f
C225 VP.n50 B 0.032763f
C226 VP.n51 B 0.259451f
C227 VP.n52 B 0.053533f
C228 VP.n53 B 0.03653f
C229 VP.n54 B 0.030703f
C230 VP.n55 B 0.030703f
C231 VP.n56 B 0.030703f
C232 VP.n57 B 0.042882f
C233 VP.n58 B 0.259451f
C234 VP.n59 B 0.042882f
C235 VP.n60 B 0.052201f
C236 VP.n61 B 0.030703f
C237 VP.n62 B 0.030703f
C238 VP.n63 B 0.030703f
C239 VP.n64 B 0.053533f
C240 VP.n65 B 0.259451f
C241 VP.n66 B 0.032763f
C242 VP.n67 B 0.061228f
C243 VP.n68 B 0.030703f
C244 VP.n69 B 0.030703f
C245 VP.n70 B 0.030703f
C246 VP.n71 B 0.060016f
C247 VP.n72 B 0.035012f
C248 VP.n73 B 0.333446f
C249 VP.n74 B 0.032593f
.ends

