* NGSPICE file created from tg_sample_0007.ext - technology: sky130A

.subckt tg_sample_0007 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t4 VGN.t0 VIN.t4 VSS.t2 sky130_fd_pr__nfet_01v8 ad=1.5366 pd=8.66 as=0.6501 ps=4.27 w=3.94 l=1.82
X1 VCC.t9 VCC.t6 VCC.t8 VCC.t7 sky130_fd_pr__pfet_01v8 ad=1.1388 pd=6.62 as=0 ps=0 w=2.92 l=3.64
X2 VOUT.t1 VGP.t0 VIN.t1 VCC.t1 sky130_fd_pr__pfet_01v8 ad=0.4818 pd=3.25 as=1.1388 ps=6.62 w=2.92 l=3.64
X3 VCC.t5 VCC.t2 VCC.t4 VCC.t3 sky130_fd_pr__pfet_01v8 ad=1.1388 pd=6.62 as=0 ps=0 w=2.92 l=3.64
X4 VOUT.t0 VGP.t1 VIN.t0 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.1388 pd=6.62 as=0.4818 ps=3.25 w=2.92 l=3.64
X5 VSS.t10 VSS.t7 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=1.5366 pd=8.66 as=0 ps=0 w=3.94 l=1.82
X6 VOUT.t3 VGN.t1 VIN.t3 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.6501 pd=4.27 as=1.5366 ps=8.66 w=3.94 l=1.82
X7 VIN.t2 VGN.t2 VOUT.t2 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.6501 pd=4.27 as=0.6501 ps=4.27 w=3.94 l=1.82
X8 VIN.t5 VGP.t2 VOUT.t5 VCC.t10 sky130_fd_pr__pfet_01v8 ad=0.4818 pd=3.25 as=0.4818 ps=3.25 w=2.92 l=3.64
X9 VSS.t6 VSS.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=1.5366 pd=8.66 as=0 ps=0 w=3.94 l=1.82
R0 VGN.n9 VGN.n0 161.3
R1 VGN.n8 VGN.n7 161.3
R2 VGN.n6 VGN.n1 161.3
R3 VGN.n5 VGN.n4 161.3
R4 VGN.n11 VGN.n10 91.2348
R5 VGN.n2 VGN.t1 82.5204
R6 VGN.n3 VGN.n2 57.6647
R7 VGN.n8 VGN.n1 56.5617
R8 VGN.n3 VGN.t2 52.173
R9 VGN.n10 VGN.t0 52.173
R10 VGN.n4 VGN.n1 24.5923
R11 VGN.n9 VGN.n8 24.5923
R12 VGN.n10 VGN.n9 19.674
R13 VGN.n5 VGN.n2 13.3418
R14 VGN.n4 VGN.n3 12.2964
R15 VGN.n11 VGN.n0 0.278335
R16 VGN.n7 VGN.n0 0.189894
R17 VGN.n7 VGN.n6 0.189894
R18 VGN.n6 VGN.n5 0.189894
R19 VGN VGN.n11 0.168637
R20 VIN.n16 VIN.n2 289.615
R21 VIN.n17 VIN.n16 185
R22 VIN.n15 VIN.n14 185
R23 VIN.n6 VIN.n5 185
R24 VIN.n9 VIN.n8 185
R25 VIN.t3 VIN.n7 147.888
R26 VIN.n1 VIN.t1 139.048
R27 VIN.n1 VIN.n0 124.495
R28 VIN.n16 VIN.n15 104.615
R29 VIN.n15 VIN.n5 104.615
R30 VIN.n8 VIN.n5 104.615
R31 VIN.n22 VIN.n21 58.7247
R32 VIN.n8 VIN.t3 52.3082
R33 VIN.n22 VIN.n20 35.9782
R34 VIN.n9 VIN.n7 15.6496
R35 VIN VIN.n1 14.2548
R36 VIN.n10 VIN.n6 12.8005
R37 VIN.n14 VIN.n13 12.0247
R38 VIN.n17 VIN.n4 11.249
R39 VIN.n0 VIN.t0 11.1323
R40 VIN.n0 VIN.t5 11.1323
R41 VIN.n18 VIN.n2 10.4732
R42 VIN.n20 VIN.n19 9.45567
R43 VIN.n19 VIN.n18 9.3005
R44 VIN.n4 VIN.n3 9.3005
R45 VIN.n13 VIN.n12 9.3005
R46 VIN.n11 VIN.n10 9.3005
R47 VIN.n21 VIN.t4 5.02588
R48 VIN.n21 VIN.t2 5.02588
R49 VIN.n11 VIN.n7 4.40546
R50 VIN.n20 VIN.n2 3.49141
R51 VIN.n18 VIN.n17 2.71565
R52 VIN.n14 VIN.n4 1.93989
R53 VIN.n13 VIN.n6 1.16414
R54 VIN VIN.n22 0.931535
R55 VIN.n10 VIN.n9 0.388379
R56 VIN.n19 VIN.n3 0.155672
R57 VIN.n12 VIN.n3 0.155672
R58 VIN.n12 VIN.n11 0.155672
R59 VOUT.n16 VOUT.n2 289.615
R60 VOUT.n17 VOUT.n16 185
R61 VOUT.n15 VOUT.n14 185
R62 VOUT.n6 VOUT.n5 185
R63 VOUT.n9 VOUT.n8 185
R64 VOUT.n1 VOUT.t0 155.727
R65 VOUT.t4 VOUT.n7 147.888
R66 VOUT.n1 VOUT.n0 141.172
R67 VOUT.n16 VOUT.n15 104.615
R68 VOUT.n15 VOUT.n5 104.615
R69 VOUT.n8 VOUT.n5 104.615
R70 VOUT.n22 VOUT.n21 75.4035
R71 VOUT.n22 VOUT.n20 52.657
R72 VOUT.n8 VOUT.t4 52.3082
R73 VOUT.n9 VOUT.n7 15.6496
R74 VOUT VOUT.n22 12.8626
R75 VOUT.n10 VOUT.n6 12.8005
R76 VOUT.n14 VOUT.n13 12.0247
R77 VOUT.n17 VOUT.n4 11.249
R78 VOUT.n0 VOUT.t5 11.1323
R79 VOUT.n0 VOUT.t1 11.1323
R80 VOUT.n18 VOUT.n2 10.4732
R81 VOUT.n20 VOUT.n19 9.45567
R82 VOUT.n19 VOUT.n18 9.3005
R83 VOUT.n4 VOUT.n3 9.3005
R84 VOUT.n13 VOUT.n12 9.3005
R85 VOUT.n11 VOUT.n10 9.3005
R86 VOUT.n21 VOUT.t2 5.02588
R87 VOUT.n21 VOUT.t3 5.02588
R88 VOUT.n11 VOUT.n7 4.40546
R89 VOUT.n20 VOUT.n2 3.49141
R90 VOUT.n18 VOUT.n17 2.71565
R91 VOUT.n14 VOUT.n4 1.93989
R92 VOUT VOUT.n1 1.8324
R93 VOUT.n13 VOUT.n6 1.16414
R94 VOUT.n10 VOUT.n9 0.388379
R95 VOUT.n19 VOUT.n3 0.155672
R96 VOUT.n12 VOUT.n3 0.155672
R97 VOUT.n12 VOUT.n11 0.155672
R98 VSS.n137 VSS.n136 585
R99 VSS.n136 VSS.n135 585
R100 VSS.n80 VSS.n79 585
R101 VSS.n79 VSS.n78 585
R102 VSS.n142 VSS.n141 585
R103 VSS.n143 VSS.n142 585
R104 VSS.n71 VSS.n70 585
R105 VSS.n72 VSS.n71 585
R106 VSS.n153 VSS.n152 585
R107 VSS.n152 VSS.n151 585
R108 VSS.n68 VSS.n67 585
R109 VSS.n67 VSS.n66 585
R110 VSS.n158 VSS.n157 585
R111 VSS.n159 VSS.n158 585
R112 VSS.n59 VSS.n58 585
R113 VSS.n60 VSS.n59 585
R114 VSS.n170 VSS.n169 585
R115 VSS.n169 VSS.n168 585
R116 VSS.n55 VSS.n53 585
R117 VSS.n167 VSS.n53 585
R118 VSS.n176 VSS.n175 585
R119 VSS.n177 VSS.n176 585
R120 VSS.n56 VSS.n54 585
R121 VSS.n54 VSS.n52 585
R122 VSS.n45 VSS.n44 585
R123 VSS.n46 VSS.n45 585
R124 VSS.n188 VSS.n187 585
R125 VSS.n187 VSS.n186 585
R126 VSS.n42 VSS.n41 585
R127 VSS.n41 VSS.n40 585
R128 VSS.n193 VSS.n192 585
R129 VSS.n194 VSS.n193 585
R130 VSS.n39 VSS.n38 585
R131 VSS.n195 VSS.n39 585
R132 VSS.n199 VSS.n198 585
R133 VSS.n198 VSS.n197 585
R134 VSS.n36 VSS.n35 585
R135 VSS.n35 VSS.n34 585
R136 VSS.n204 VSS.n203 585
R137 VSS.n205 VSS.n204 585
R138 VSS.n33 VSS.n32 585
R139 VSS.n206 VSS.n33 585
R140 VSS.n210 VSS.n209 585
R141 VSS.n209 VSS.n208 585
R142 VSS.n30 VSS.n29 585
R143 VSS.n29 VSS.n28 585
R144 VSS.n215 VSS.n214 585
R145 VSS.n216 VSS.n215 585
R146 VSS.n27 VSS.n26 585
R147 VSS.n217 VSS.n27 585
R148 VSS.n221 VSS.n220 585
R149 VSS.n220 VSS.n219 585
R150 VSS.n24 VSS.n22 585
R151 VSS.n22 VSS.n20 585
R152 VSS.n274 VSS.n273 585
R153 VSS.n275 VSS.n274 585
R154 VSS.n277 VSS.n276 585
R155 VSS.n276 VSS.n275 585
R156 VSS.n278 VSS.n18 585
R157 VSS.n20 VSS.n18 585
R158 VSS.n218 VSS.n16 585
R159 VSS.n219 VSS.n218 585
R160 VSS.n282 VSS.n15 585
R161 VSS.n217 VSS.n15 585
R162 VSS.n283 VSS.n14 585
R163 VSS.n216 VSS.n14 585
R164 VSS.n284 VSS.n13 585
R165 VSS.n28 VSS.n13 585
R166 VSS.n207 VSS.n11 585
R167 VSS.n208 VSS.n207 585
R168 VSS.n288 VSS.n10 585
R169 VSS.n206 VSS.n10 585
R170 VSS.n289 VSS.n9 585
R171 VSS.n205 VSS.n9 585
R172 VSS.n290 VSS.n8 585
R173 VSS.n34 VSS.n8 585
R174 VSS.n196 VSS.n6 585
R175 VSS.n197 VSS.n196 585
R176 VSS.n294 VSS.n5 585
R177 VSS.n195 VSS.n5 585
R178 VSS.n295 VSS.n4 585
R179 VSS.n194 VSS.n4 585
R180 VSS.n296 VSS.n3 585
R181 VSS.n40 VSS.n3 585
R182 VSS.n185 VSS.n2 585
R183 VSS.n186 VSS.n185 585
R184 VSS.n184 VSS.n183 585
R185 VSS.n184 VSS.n46 585
R186 VSS.n48 VSS.n47 585
R187 VSS.n52 VSS.n47 585
R188 VSS.n179 VSS.n178 585
R189 VSS.n178 VSS.n177 585
R190 VSS.n51 VSS.n50 585
R191 VSS.n167 VSS.n51 585
R192 VSS.n166 VSS.n165 585
R193 VSS.n168 VSS.n166 585
R194 VSS.n62 VSS.n61 585
R195 VSS.n61 VSS.n60 585
R196 VSS.n161 VSS.n160 585
R197 VSS.n160 VSS.n159 585
R198 VSS.n65 VSS.n64 585
R199 VSS.n66 VSS.n65 585
R200 VSS.n150 VSS.n149 585
R201 VSS.n151 VSS.n150 585
R202 VSS.n74 VSS.n73 585
R203 VSS.n73 VSS.n72 585
R204 VSS.n145 VSS.n144 585
R205 VSS.n144 VSS.n143 585
R206 VSS.n77 VSS.n76 585
R207 VSS.n78 VSS.n77 585
R208 VSS.n134 VSS.n133 585
R209 VSS.n135 VSS.n134 585
R210 VSS.n240 VSS.n19 585
R211 VSS.n241 VSS.n236 585
R212 VSS.n243 VSS.n242 585
R213 VSS.n245 VSS.n233 585
R214 VSS.n247 VSS.n246 585
R215 VSS.n248 VSS.n232 585
R216 VSS.n250 VSS.n249 585
R217 VSS.n252 VSS.n230 585
R218 VSS.n254 VSS.n253 585
R219 VSS.n255 VSS.n229 585
R220 VSS.n257 VSS.n256 585
R221 VSS.n259 VSS.n227 585
R222 VSS.n261 VSS.n260 585
R223 VSS.n262 VSS.n226 585
R224 VSS.n264 VSS.n263 585
R225 VSS.n266 VSS.n225 585
R226 VSS.n267 VSS.n224 585
R227 VSS.n270 VSS.n269 585
R228 VSS.n271 VSS.n23 585
R229 VSS.n23 VSS.n21 585
R230 VSS.n82 VSS.n81 585
R231 VSS.n95 VSS.n94 585
R232 VSS.n96 VSS.n92 585
R233 VSS.n92 VSS.n83 585
R234 VSS.n98 VSS.n97 585
R235 VSS.n100 VSS.n91 585
R236 VSS.n103 VSS.n102 585
R237 VSS.n104 VSS.n90 585
R238 VSS.n106 VSS.n105 585
R239 VSS.n108 VSS.n89 585
R240 VSS.n111 VSS.n110 585
R241 VSS.n112 VSS.n88 585
R242 VSS.n114 VSS.n113 585
R243 VSS.n116 VSS.n87 585
R244 VSS.n119 VSS.n118 585
R245 VSS.n120 VSS.n86 585
R246 VSS.n125 VSS.n124 585
R247 VSS.n127 VSS.n85 585
R248 VSS.n130 VSS.n129 585
R249 VSS.n131 VSS.n84 585
R250 VSS.n136 VSS.n82 569.379
R251 VSS.n134 VSS.n84 569.379
R252 VSS.n274 VSS.n23 569.379
R253 VSS.n276 VSS.n19 569.379
R254 VSS.n135 VSS.n83 417.82
R255 VSS.n275 VSS.n21 417.82
R256 VSS.n237 VSS.t3 258.635
R257 VSS.n121 VSS.t7 258.635
R258 VSS.n135 VSS.n78 257.913
R259 VSS.n143 VSS.n78 257.913
R260 VSS.n151 VSS.n72 257.913
R261 VSS.n151 VSS.n66 257.913
R262 VSS.n159 VSS.n66 257.913
R263 VSS.n159 VSS.n60 257.913
R264 VSS.n168 VSS.n60 257.913
R265 VSS.n168 VSS.n167 257.913
R266 VSS.n177 VSS.n52 257.913
R267 VSS.n52 VSS.n46 257.913
R268 VSS.n186 VSS.n46 257.913
R269 VSS.n194 VSS.n40 257.913
R270 VSS.n195 VSS.n194 257.913
R271 VSS.n197 VSS.n195 257.913
R272 VSS.n205 VSS.n34 257.913
R273 VSS.n206 VSS.n205 257.913
R274 VSS.n208 VSS.n206 257.913
R275 VSS.n208 VSS.n28 257.913
R276 VSS.n216 VSS.n28 257.913
R277 VSS.n217 VSS.n216 257.913
R278 VSS.n219 VSS.n20 257.913
R279 VSS.n275 VSS.n20 257.913
R280 VSS.n235 VSS.n21 256.663
R281 VSS.n244 VSS.n21 256.663
R282 VSS.n234 VSS.n21 256.663
R283 VSS.n251 VSS.n21 256.663
R284 VSS.n231 VSS.n21 256.663
R285 VSS.n258 VSS.n21 256.663
R286 VSS.n228 VSS.n21 256.663
R287 VSS.n265 VSS.n21 256.663
R288 VSS.n268 VSS.n21 256.663
R289 VSS.n93 VSS.n83 256.663
R290 VSS.n99 VSS.n83 256.663
R291 VSS.n101 VSS.n83 256.663
R292 VSS.n107 VSS.n83 256.663
R293 VSS.n109 VSS.n83 256.663
R294 VSS.n115 VSS.n83 256.663
R295 VSS.n117 VSS.n83 256.663
R296 VSS.n126 VSS.n83 256.663
R297 VSS.n128 VSS.n83 256.663
R298 VSS.n136 VSS.n79 240.244
R299 VSS.n142 VSS.n79 240.244
R300 VSS.n142 VSS.n71 240.244
R301 VSS.n152 VSS.n71 240.244
R302 VSS.n152 VSS.n67 240.244
R303 VSS.n158 VSS.n67 240.244
R304 VSS.n158 VSS.n59 240.244
R305 VSS.n169 VSS.n59 240.244
R306 VSS.n169 VSS.n53 240.244
R307 VSS.n176 VSS.n53 240.244
R308 VSS.n176 VSS.n54 240.244
R309 VSS.n54 VSS.n45 240.244
R310 VSS.n187 VSS.n45 240.244
R311 VSS.n187 VSS.n41 240.244
R312 VSS.n193 VSS.n41 240.244
R313 VSS.n193 VSS.n39 240.244
R314 VSS.n198 VSS.n39 240.244
R315 VSS.n198 VSS.n35 240.244
R316 VSS.n204 VSS.n35 240.244
R317 VSS.n204 VSS.n33 240.244
R318 VSS.n209 VSS.n33 240.244
R319 VSS.n209 VSS.n29 240.244
R320 VSS.n215 VSS.n29 240.244
R321 VSS.n215 VSS.n27 240.244
R322 VSS.n220 VSS.n27 240.244
R323 VSS.n220 VSS.n22 240.244
R324 VSS.n274 VSS.n22 240.244
R325 VSS.n134 VSS.n77 240.244
R326 VSS.n144 VSS.n77 240.244
R327 VSS.n144 VSS.n73 240.244
R328 VSS.n150 VSS.n73 240.244
R329 VSS.n150 VSS.n65 240.244
R330 VSS.n160 VSS.n65 240.244
R331 VSS.n160 VSS.n61 240.244
R332 VSS.n166 VSS.n61 240.244
R333 VSS.n166 VSS.n51 240.244
R334 VSS.n178 VSS.n51 240.244
R335 VSS.n178 VSS.n47 240.244
R336 VSS.n184 VSS.n47 240.244
R337 VSS.n185 VSS.n184 240.244
R338 VSS.n185 VSS.n3 240.244
R339 VSS.n4 VSS.n3 240.244
R340 VSS.n5 VSS.n4 240.244
R341 VSS.n196 VSS.n5 240.244
R342 VSS.n196 VSS.n8 240.244
R343 VSS.n9 VSS.n8 240.244
R344 VSS.n10 VSS.n9 240.244
R345 VSS.n207 VSS.n10 240.244
R346 VSS.n207 VSS.n13 240.244
R347 VSS.n14 VSS.n13 240.244
R348 VSS.n15 VSS.n14 240.244
R349 VSS.n218 VSS.n15 240.244
R350 VSS.n218 VSS.n18 240.244
R351 VSS.n276 VSS.n18 240.244
R352 VSS.n177 VSS.t2 206.332
R353 VSS.n197 VSS.t1 206.332
R354 VSS.n237 VSS.t5 185.793
R355 VSS.n121 VSS.t10 185.793
R356 VSS.n143 VSS.t8 185.698
R357 VSS.n219 VSS.t4 185.698
R358 VSS.n94 VSS.n92 163.367
R359 VSS.n98 VSS.n92 163.367
R360 VSS.n102 VSS.n100 163.367
R361 VSS.n106 VSS.n90 163.367
R362 VSS.n110 VSS.n108 163.367
R363 VSS.n114 VSS.n88 163.367
R364 VSS.n118 VSS.n116 163.367
R365 VSS.n125 VSS.n86 163.367
R366 VSS.n129 VSS.n127 163.367
R367 VSS.n269 VSS.n23 163.367
R368 VSS.n267 VSS.n266 163.367
R369 VSS.n264 VSS.n226 163.367
R370 VSS.n260 VSS.n259 163.367
R371 VSS.n257 VSS.n229 163.367
R372 VSS.n253 VSS.n252 163.367
R373 VSS.n250 VSS.n232 163.367
R374 VSS.n246 VSS.n245 163.367
R375 VSS.n243 VSS.n236 163.367
R376 VSS.n238 VSS.t6 144.096
R377 VSS.n122 VSS.t9 144.096
R378 VSS.n186 VSS.t0 128.958
R379 VSS.t0 VSS.n40 128.958
R380 VSS.t8 VSS.n72 72.2162
R381 VSS.t4 VSS.n217 72.2162
R382 VSS.n93 VSS.n82 71.676
R383 VSS.n99 VSS.n98 71.676
R384 VSS.n102 VSS.n101 71.676
R385 VSS.n107 VSS.n106 71.676
R386 VSS.n110 VSS.n109 71.676
R387 VSS.n115 VSS.n114 71.676
R388 VSS.n118 VSS.n117 71.676
R389 VSS.n126 VSS.n125 71.676
R390 VSS.n129 VSS.n128 71.676
R391 VSS.n268 VSS.n267 71.676
R392 VSS.n265 VSS.n264 71.676
R393 VSS.n260 VSS.n228 71.676
R394 VSS.n258 VSS.n257 71.676
R395 VSS.n253 VSS.n231 71.676
R396 VSS.n251 VSS.n250 71.676
R397 VSS.n246 VSS.n234 71.676
R398 VSS.n244 VSS.n243 71.676
R399 VSS.n235 VSS.n19 71.676
R400 VSS.n236 VSS.n235 71.676
R401 VSS.n245 VSS.n244 71.676
R402 VSS.n234 VSS.n232 71.676
R403 VSS.n252 VSS.n251 71.676
R404 VSS.n231 VSS.n229 71.676
R405 VSS.n259 VSS.n258 71.676
R406 VSS.n228 VSS.n226 71.676
R407 VSS.n266 VSS.n265 71.676
R408 VSS.n269 VSS.n268 71.676
R409 VSS.n94 VSS.n93 71.676
R410 VSS.n100 VSS.n99 71.676
R411 VSS.n101 VSS.n90 71.676
R412 VSS.n108 VSS.n107 71.676
R413 VSS.n109 VSS.n88 71.676
R414 VSS.n116 VSS.n115 71.676
R415 VSS.n117 VSS.n86 71.676
R416 VSS.n127 VSS.n126 71.676
R417 VSS.n128 VSS.n84 71.676
R418 VSS.n167 VSS.t2 51.5831
R419 VSS.t1 VSS.n34 51.5831
R420 VSS.n238 VSS.n237 41.6975
R421 VSS.n122 VSS.n121 41.6975
R422 VSS.n239 VSS.n238 34.5217
R423 VSS.n123 VSS.n122 34.5217
R424 VSS.n272 VSS.n271 27.6548
R425 VSS.n240 VSS.n17 27.6548
R426 VSS.n138 VSS.n81 27.6548
R427 VSS.n132 VSS.n131 27.6548
R428 VSS.n137 VSS.n80 19.3944
R429 VSS.n141 VSS.n80 19.3944
R430 VSS.n141 VSS.n70 19.3944
R431 VSS.n153 VSS.n70 19.3944
R432 VSS.n153 VSS.n68 19.3944
R433 VSS.n157 VSS.n68 19.3944
R434 VSS.n157 VSS.n58 19.3944
R435 VSS.n170 VSS.n58 19.3944
R436 VSS.n170 VSS.n55 19.3944
R437 VSS.n175 VSS.n55 19.3944
R438 VSS.n175 VSS.n56 19.3944
R439 VSS.n56 VSS.n44 19.3944
R440 VSS.n188 VSS.n44 19.3944
R441 VSS.n188 VSS.n42 19.3944
R442 VSS.n192 VSS.n42 19.3944
R443 VSS.n192 VSS.n38 19.3944
R444 VSS.n199 VSS.n38 19.3944
R445 VSS.n199 VSS.n36 19.3944
R446 VSS.n203 VSS.n36 19.3944
R447 VSS.n203 VSS.n32 19.3944
R448 VSS.n210 VSS.n32 19.3944
R449 VSS.n210 VSS.n30 19.3944
R450 VSS.n214 VSS.n30 19.3944
R451 VSS.n214 VSS.n26 19.3944
R452 VSS.n221 VSS.n26 19.3944
R453 VSS.n221 VSS.n24 19.3944
R454 VSS.n273 VSS.n24 19.3944
R455 VSS.n133 VSS.n76 19.3944
R456 VSS.n145 VSS.n76 19.3944
R457 VSS.n145 VSS.n74 19.3944
R458 VSS.n149 VSS.n74 19.3944
R459 VSS.n149 VSS.n64 19.3944
R460 VSS.n161 VSS.n64 19.3944
R461 VSS.n161 VSS.n62 19.3944
R462 VSS.n165 VSS.n62 19.3944
R463 VSS.n165 VSS.n50 19.3944
R464 VSS.n179 VSS.n50 19.3944
R465 VSS.n179 VSS.n48 19.3944
R466 VSS.n183 VSS.n48 19.3944
R467 VSS.n183 VSS.n2 19.3944
R468 VSS.n296 VSS.n2 19.3944
R469 VSS.n296 VSS.n295 19.3944
R470 VSS.n295 VSS.n294 19.3944
R471 VSS.n294 VSS.n6 19.3944
R472 VSS.n290 VSS.n6 19.3944
R473 VSS.n290 VSS.n289 19.3944
R474 VSS.n289 VSS.n288 19.3944
R475 VSS.n288 VSS.n11 19.3944
R476 VSS.n284 VSS.n11 19.3944
R477 VSS.n284 VSS.n283 19.3944
R478 VSS.n283 VSS.n282 19.3944
R479 VSS.n282 VSS.n16 19.3944
R480 VSS.n278 VSS.n16 19.3944
R481 VSS.n278 VSS.n277 19.3944
R482 VSS.n271 VSS.n270 10.6151
R483 VSS.n270 VSS.n224 10.6151
R484 VSS.n225 VSS.n224 10.6151
R485 VSS.n263 VSS.n225 10.6151
R486 VSS.n263 VSS.n262 10.6151
R487 VSS.n262 VSS.n261 10.6151
R488 VSS.n261 VSS.n227 10.6151
R489 VSS.n256 VSS.n227 10.6151
R490 VSS.n256 VSS.n255 10.6151
R491 VSS.n255 VSS.n254 10.6151
R492 VSS.n254 VSS.n230 10.6151
R493 VSS.n249 VSS.n230 10.6151
R494 VSS.n249 VSS.n248 10.6151
R495 VSS.n248 VSS.n247 10.6151
R496 VSS.n247 VSS.n233 10.6151
R497 VSS.n242 VSS.n241 10.6151
R498 VSS.n241 VSS.n240 10.6151
R499 VSS.n95 VSS.n81 10.6151
R500 VSS.n96 VSS.n95 10.6151
R501 VSS.n97 VSS.n96 10.6151
R502 VSS.n97 VSS.n91 10.6151
R503 VSS.n103 VSS.n91 10.6151
R504 VSS.n104 VSS.n103 10.6151
R505 VSS.n105 VSS.n104 10.6151
R506 VSS.n105 VSS.n89 10.6151
R507 VSS.n111 VSS.n89 10.6151
R508 VSS.n112 VSS.n111 10.6151
R509 VSS.n113 VSS.n112 10.6151
R510 VSS.n113 VSS.n87 10.6151
R511 VSS.n119 VSS.n87 10.6151
R512 VSS.n120 VSS.n119 10.6151
R513 VSS.n124 VSS.n120 10.6151
R514 VSS.n130 VSS.n85 10.6151
R515 VSS.n131 VSS.n130 10.6151
R516 VSS.n295 VSS.n0 9.3005
R517 VSS.n294 VSS.n293 9.3005
R518 VSS.n292 VSS.n6 9.3005
R519 VSS.n291 VSS.n290 9.3005
R520 VSS.n289 VSS.n7 9.3005
R521 VSS.n288 VSS.n287 9.3005
R522 VSS.n286 VSS.n11 9.3005
R523 VSS.n285 VSS.n284 9.3005
R524 VSS.n283 VSS.n12 9.3005
R525 VSS.n282 VSS.n281 9.3005
R526 VSS.n280 VSS.n16 9.3005
R527 VSS.n279 VSS.n278 9.3005
R528 VSS.n277 VSS.n17 9.3005
R529 VSS.n138 VSS.n137 9.3005
R530 VSS.n139 VSS.n80 9.3005
R531 VSS.n141 VSS.n140 9.3005
R532 VSS.n70 VSS.n69 9.3005
R533 VSS.n154 VSS.n153 9.3005
R534 VSS.n155 VSS.n68 9.3005
R535 VSS.n157 VSS.n156 9.3005
R536 VSS.n58 VSS.n57 9.3005
R537 VSS.n171 VSS.n170 9.3005
R538 VSS.n172 VSS.n55 9.3005
R539 VSS.n175 VSS.n174 9.3005
R540 VSS.n173 VSS.n56 9.3005
R541 VSS.n44 VSS.n43 9.3005
R542 VSS.n189 VSS.n188 9.3005
R543 VSS.n190 VSS.n42 9.3005
R544 VSS.n192 VSS.n191 9.3005
R545 VSS.n38 VSS.n37 9.3005
R546 VSS.n200 VSS.n199 9.3005
R547 VSS.n201 VSS.n36 9.3005
R548 VSS.n203 VSS.n202 9.3005
R549 VSS.n32 VSS.n31 9.3005
R550 VSS.n211 VSS.n210 9.3005
R551 VSS.n212 VSS.n30 9.3005
R552 VSS.n214 VSS.n213 9.3005
R553 VSS.n26 VSS.n25 9.3005
R554 VSS.n222 VSS.n221 9.3005
R555 VSS.n223 VSS.n24 9.3005
R556 VSS.n273 VSS.n272 9.3005
R557 VSS.n76 VSS.n75 9.3005
R558 VSS.n146 VSS.n145 9.3005
R559 VSS.n147 VSS.n74 9.3005
R560 VSS.n149 VSS.n148 9.3005
R561 VSS.n64 VSS.n63 9.3005
R562 VSS.n162 VSS.n161 9.3005
R563 VSS.n163 VSS.n62 9.3005
R564 VSS.n165 VSS.n164 9.3005
R565 VSS.n50 VSS.n49 9.3005
R566 VSS.n180 VSS.n179 9.3005
R567 VSS.n181 VSS.n48 9.3005
R568 VSS.n183 VSS.n182 9.3005
R569 VSS.n2 VSS.n1 9.3005
R570 VSS.n133 VSS.n132 9.3005
R571 VSS VSS.n296 9.3005
R572 VSS.n239 VSS.n233 8.58587
R573 VSS.n124 VSS.n123 8.58587
R574 VSS.n242 VSS.n239 2.02977
R575 VSS.n123 VSS.n85 2.02977
R576 VSS VSS.n0 0.152939
R577 VSS.n293 VSS.n0 0.152939
R578 VSS.n293 VSS.n292 0.152939
R579 VSS.n292 VSS.n291 0.152939
R580 VSS.n291 VSS.n7 0.152939
R581 VSS.n287 VSS.n7 0.152939
R582 VSS.n287 VSS.n286 0.152939
R583 VSS.n286 VSS.n285 0.152939
R584 VSS.n285 VSS.n12 0.152939
R585 VSS.n281 VSS.n12 0.152939
R586 VSS.n281 VSS.n280 0.152939
R587 VSS.n280 VSS.n279 0.152939
R588 VSS.n279 VSS.n17 0.152939
R589 VSS.n139 VSS.n138 0.152939
R590 VSS.n140 VSS.n139 0.152939
R591 VSS.n140 VSS.n69 0.152939
R592 VSS.n154 VSS.n69 0.152939
R593 VSS.n155 VSS.n154 0.152939
R594 VSS.n156 VSS.n155 0.152939
R595 VSS.n156 VSS.n57 0.152939
R596 VSS.n171 VSS.n57 0.152939
R597 VSS.n172 VSS.n171 0.152939
R598 VSS.n174 VSS.n172 0.152939
R599 VSS.n174 VSS.n173 0.152939
R600 VSS.n173 VSS.n43 0.152939
R601 VSS.n189 VSS.n43 0.152939
R602 VSS.n190 VSS.n189 0.152939
R603 VSS.n191 VSS.n190 0.152939
R604 VSS.n191 VSS.n37 0.152939
R605 VSS.n200 VSS.n37 0.152939
R606 VSS.n201 VSS.n200 0.152939
R607 VSS.n202 VSS.n201 0.152939
R608 VSS.n202 VSS.n31 0.152939
R609 VSS.n211 VSS.n31 0.152939
R610 VSS.n212 VSS.n211 0.152939
R611 VSS.n213 VSS.n212 0.152939
R612 VSS.n213 VSS.n25 0.152939
R613 VSS.n222 VSS.n25 0.152939
R614 VSS.n223 VSS.n222 0.152939
R615 VSS.n272 VSS.n223 0.152939
R616 VSS.n132 VSS.n75 0.152939
R617 VSS.n146 VSS.n75 0.152939
R618 VSS.n147 VSS.n146 0.152939
R619 VSS.n148 VSS.n147 0.152939
R620 VSS.n148 VSS.n63 0.152939
R621 VSS.n162 VSS.n63 0.152939
R622 VSS.n163 VSS.n162 0.152939
R623 VSS.n164 VSS.n163 0.152939
R624 VSS.n164 VSS.n49 0.152939
R625 VSS.n180 VSS.n49 0.152939
R626 VSS.n181 VSS.n180 0.152939
R627 VSS.n182 VSS.n181 0.152939
R628 VSS.n182 VSS.n1 0.152939
R629 VSS VSS.n1 0.1255
R630 VCC.n359 VCC.n30 406.829
R631 VCC.n332 VCC.n331 406.829
R632 VCC.n182 VCC.n138 406.829
R633 VCC.n180 VCC.n140 406.829
R634 VCC.n41 VCC.t2 228.548
R635 VCC.n141 VCC.t6 228.548
R636 VCC.n41 VCC.t4 220.963
R637 VCC.n141 VCC.t9 220.963
R638 VCC.n331 VCC.n330 185
R639 VCC.n331 VCC.n33 185
R640 VCC.n329 VCC.n45 185
R641 VCC.n320 VCC.n45 185
R642 VCC.n50 VCC.n46 185
R643 VCC.n321 VCC.n50 185
R644 VCC.n325 VCC.n324 185
R645 VCC.n324 VCC.n323 185
R646 VCC.n49 VCC.n48 185
R647 VCC.n319 VCC.n49 185
R648 VCC.n317 VCC.n316 185
R649 VCC.n318 VCC.n317 185
R650 VCC.n53 VCC.n52 185
R651 VCC.n52 VCC.n51 185
R652 VCC.n312 VCC.n311 185
R653 VCC.n311 VCC.n310 185
R654 VCC.n56 VCC.n55 185
R655 VCC.n308 VCC.n56 185
R656 VCC.n306 VCC.n305 185
R657 VCC.n307 VCC.n306 185
R658 VCC.n59 VCC.n58 185
R659 VCC.n58 VCC.n57 185
R660 VCC.n301 VCC.n300 185
R661 VCC.n300 VCC.n299 185
R662 VCC.n62 VCC.n61 185
R663 VCC.n297 VCC.n62 185
R664 VCC.n295 VCC.n294 185
R665 VCC.n296 VCC.n295 185
R666 VCC.n65 VCC.n64 185
R667 VCC.n64 VCC.n63 185
R668 VCC.n290 VCC.n289 185
R669 VCC.n289 VCC.n288 185
R670 VCC.n68 VCC.n67 185
R671 VCC.n286 VCC.n68 185
R672 VCC.n284 VCC.n283 185
R673 VCC.n285 VCC.n284 185
R674 VCC.n71 VCC.n70 185
R675 VCC.n70 VCC.n69 185
R676 VCC.n279 VCC.n278 185
R677 VCC.n278 VCC.n277 185
R678 VCC.n74 VCC.n73 185
R679 VCC.n275 VCC.n74 185
R680 VCC.n273 VCC.n272 185
R681 VCC.n274 VCC.n273 185
R682 VCC.n76 VCC.n75 185
R683 VCC.n75 VCC.t10 185
R684 VCC.n268 VCC.n267 185
R685 VCC.n267 VCC.n266 185
R686 VCC.n79 VCC.n78 185
R687 VCC.n80 VCC.n79 185
R688 VCC.n255 VCC.n254 185
R689 VCC.n256 VCC.n255 185
R690 VCC.n88 VCC.n87 185
R691 VCC.n257 VCC.n87 185
R692 VCC.n250 VCC.n249 185
R693 VCC.n249 VCC.n86 185
R694 VCC.n248 VCC.n90 185
R695 VCC.n248 VCC.n247 185
R696 VCC.n101 VCC.n91 185
R697 VCC.n92 VCC.n91 185
R698 VCC.n238 VCC.n237 185
R699 VCC.n239 VCC.n238 185
R700 VCC.n100 VCC.n99 185
R701 VCC.n99 VCC.n98 185
R702 VCC.n232 VCC.n231 185
R703 VCC.n231 VCC.n230 185
R704 VCC.n104 VCC.n103 185
R705 VCC.n105 VCC.n104 185
R706 VCC.n221 VCC.n220 185
R707 VCC.n222 VCC.n221 185
R708 VCC.n113 VCC.n112 185
R709 VCC.n112 VCC.n111 185
R710 VCC.n216 VCC.n215 185
R711 VCC.n215 VCC.n214 185
R712 VCC.n116 VCC.n115 185
R713 VCC.n117 VCC.n116 185
R714 VCC.n205 VCC.n204 185
R715 VCC.n206 VCC.n205 185
R716 VCC.n125 VCC.n124 185
R717 VCC.n124 VCC.n123 185
R718 VCC.n200 VCC.n199 185
R719 VCC.n199 VCC.n198 185
R720 VCC.n128 VCC.n127 185
R721 VCC.n189 VCC.n128 185
R722 VCC.n188 VCC.n187 185
R723 VCC.n190 VCC.n188 185
R724 VCC.n136 VCC.n135 185
R725 VCC.n135 VCC.n134 185
R726 VCC.n183 VCC.n182 185
R727 VCC.n182 VCC.n181 185
R728 VCC.n180 VCC.n179 185
R729 VCC.n181 VCC.n180 185
R730 VCC.n133 VCC.n132 185
R731 VCC.n134 VCC.n133 185
R732 VCC.n192 VCC.n191 185
R733 VCC.n191 VCC.n190 185
R734 VCC.n130 VCC.n129 185
R735 VCC.n189 VCC.n129 185
R736 VCC.n197 VCC.n196 185
R737 VCC.n198 VCC.n197 185
R738 VCC.n122 VCC.n121 185
R739 VCC.n123 VCC.n122 185
R740 VCC.n208 VCC.n207 185
R741 VCC.n207 VCC.n206 185
R742 VCC.n119 VCC.n118 185
R743 VCC.n118 VCC.n117 185
R744 VCC.n213 VCC.n212 185
R745 VCC.n214 VCC.n213 185
R746 VCC.n110 VCC.n109 185
R747 VCC.n111 VCC.n110 185
R748 VCC.n224 VCC.n223 185
R749 VCC.n223 VCC.n222 185
R750 VCC.n107 VCC.n106 185
R751 VCC.n106 VCC.n105 185
R752 VCC.n229 VCC.n228 185
R753 VCC.n230 VCC.n229 185
R754 VCC.n97 VCC.n96 185
R755 VCC.n98 VCC.n97 185
R756 VCC.n241 VCC.n240 185
R757 VCC.n240 VCC.n239 185
R758 VCC.n94 VCC.n93 185
R759 VCC.n93 VCC.n92 185
R760 VCC.n246 VCC.n245 185
R761 VCC.n247 VCC.n246 185
R762 VCC.n85 VCC.n84 185
R763 VCC.n86 VCC.n85 185
R764 VCC.n259 VCC.n258 185
R765 VCC.n258 VCC.n257 185
R766 VCC.n82 VCC.n81 185
R767 VCC.n256 VCC.n81 185
R768 VCC.n264 VCC.n263 185
R769 VCC.n264 VCC.n80 185
R770 VCC.n265 VCC.n2 185
R771 VCC.n266 VCC.n265 185
R772 VCC.n394 VCC.n3 185
R773 VCC.t10 VCC.n3 185
R774 VCC.n393 VCC.n4 185
R775 VCC.n274 VCC.n4 185
R776 VCC.n392 VCC.n5 185
R777 VCC.n275 VCC.n5 185
R778 VCC.n276 VCC.n6 185
R779 VCC.n277 VCC.n276 185
R780 VCC.n388 VCC.n8 185
R781 VCC.n69 VCC.n8 185
R782 VCC.n387 VCC.n9 185
R783 VCC.n285 VCC.n9 185
R784 VCC.n386 VCC.n10 185
R785 VCC.n286 VCC.n10 185
R786 VCC.n287 VCC.n11 185
R787 VCC.n288 VCC.n287 185
R788 VCC.n382 VCC.n13 185
R789 VCC.n63 VCC.n13 185
R790 VCC.n381 VCC.n14 185
R791 VCC.n296 VCC.n14 185
R792 VCC.n380 VCC.n15 185
R793 VCC.n297 VCC.n15 185
R794 VCC.n298 VCC.n16 185
R795 VCC.n299 VCC.n298 185
R796 VCC.n376 VCC.n18 185
R797 VCC.n57 VCC.n18 185
R798 VCC.n375 VCC.n19 185
R799 VCC.n307 VCC.n19 185
R800 VCC.n374 VCC.n20 185
R801 VCC.n308 VCC.n20 185
R802 VCC.n309 VCC.n21 185
R803 VCC.n310 VCC.n309 185
R804 VCC.n370 VCC.n23 185
R805 VCC.n51 VCC.n23 185
R806 VCC.n369 VCC.n24 185
R807 VCC.n318 VCC.n24 185
R808 VCC.n368 VCC.n25 185
R809 VCC.n319 VCC.n25 185
R810 VCC.n322 VCC.n26 185
R811 VCC.n323 VCC.n322 185
R812 VCC.n364 VCC.n28 185
R813 VCC.n321 VCC.n28 185
R814 VCC.n363 VCC.n29 185
R815 VCC.n320 VCC.n29 185
R816 VCC.n362 VCC.n30 185
R817 VCC.n33 VCC.n30 185
R818 VCC.n333 VCC.n332 185
R819 VCC.n335 VCC.n334 185
R820 VCC.n337 VCC.n336 185
R821 VCC.n339 VCC.n338 185
R822 VCC.n341 VCC.n340 185
R823 VCC.n343 VCC.n342 185
R824 VCC.n345 VCC.n344 185
R825 VCC.n347 VCC.n346 185
R826 VCC.n349 VCC.n348 185
R827 VCC.n351 VCC.n350 185
R828 VCC.n353 VCC.n352 185
R829 VCC.n354 VCC.n40 185
R830 VCC.n356 VCC.n355 185
R831 VCC.n32 VCC.n31 185
R832 VCC.n360 VCC.n359 185
R833 VCC.n359 VCC.n358 185
R834 VCC.n177 VCC.n140 185
R835 VCC.n176 VCC.n175 185
R836 VCC.n173 VCC.n172 185
R837 VCC.n173 VCC.n139 185
R838 VCC.n171 VCC.n144 185
R839 VCC.n170 VCC.n169 185
R840 VCC.n167 VCC.n145 185
R841 VCC.n165 VCC.n164 185
R842 VCC.n163 VCC.n146 185
R843 VCC.n162 VCC.n161 185
R844 VCC.n159 VCC.n147 185
R845 VCC.n157 VCC.n156 185
R846 VCC.n155 VCC.n148 185
R847 VCC.n154 VCC.n153 185
R848 VCC.n151 VCC.n149 185
R849 VCC.n138 VCC.n137 185
R850 VCC.n182 VCC.n135 146.341
R851 VCC.n188 VCC.n135 146.341
R852 VCC.n188 VCC.n128 146.341
R853 VCC.n199 VCC.n128 146.341
R854 VCC.n199 VCC.n124 146.341
R855 VCC.n205 VCC.n124 146.341
R856 VCC.n205 VCC.n116 146.341
R857 VCC.n215 VCC.n116 146.341
R858 VCC.n215 VCC.n112 146.341
R859 VCC.n221 VCC.n112 146.341
R860 VCC.n221 VCC.n104 146.341
R861 VCC.n231 VCC.n104 146.341
R862 VCC.n231 VCC.n99 146.341
R863 VCC.n238 VCC.n99 146.341
R864 VCC.n238 VCC.n91 146.341
R865 VCC.n248 VCC.n91 146.341
R866 VCC.n249 VCC.n248 146.341
R867 VCC.n249 VCC.n87 146.341
R868 VCC.n255 VCC.n87 146.341
R869 VCC.n255 VCC.n79 146.341
R870 VCC.n267 VCC.n79 146.341
R871 VCC.n267 VCC.n75 146.341
R872 VCC.n273 VCC.n75 146.341
R873 VCC.n273 VCC.n74 146.341
R874 VCC.n278 VCC.n74 146.341
R875 VCC.n278 VCC.n70 146.341
R876 VCC.n284 VCC.n70 146.341
R877 VCC.n284 VCC.n68 146.341
R878 VCC.n289 VCC.n68 146.341
R879 VCC.n289 VCC.n64 146.341
R880 VCC.n295 VCC.n64 146.341
R881 VCC.n295 VCC.n62 146.341
R882 VCC.n300 VCC.n62 146.341
R883 VCC.n300 VCC.n58 146.341
R884 VCC.n306 VCC.n58 146.341
R885 VCC.n306 VCC.n56 146.341
R886 VCC.n311 VCC.n56 146.341
R887 VCC.n311 VCC.n52 146.341
R888 VCC.n317 VCC.n52 146.341
R889 VCC.n317 VCC.n49 146.341
R890 VCC.n324 VCC.n49 146.341
R891 VCC.n324 VCC.n50 146.341
R892 VCC.n50 VCC.n45 146.341
R893 VCC.n331 VCC.n45 146.341
R894 VCC.n180 VCC.n133 146.341
R895 VCC.n191 VCC.n133 146.341
R896 VCC.n191 VCC.n129 146.341
R897 VCC.n197 VCC.n129 146.341
R898 VCC.n197 VCC.n122 146.341
R899 VCC.n207 VCC.n122 146.341
R900 VCC.n207 VCC.n118 146.341
R901 VCC.n213 VCC.n118 146.341
R902 VCC.n213 VCC.n110 146.341
R903 VCC.n223 VCC.n110 146.341
R904 VCC.n223 VCC.n106 146.341
R905 VCC.n229 VCC.n106 146.341
R906 VCC.n229 VCC.n97 146.341
R907 VCC.n240 VCC.n97 146.341
R908 VCC.n240 VCC.n93 146.341
R909 VCC.n246 VCC.n93 146.341
R910 VCC.n246 VCC.n85 146.341
R911 VCC.n258 VCC.n85 146.341
R912 VCC.n258 VCC.n81 146.341
R913 VCC.n264 VCC.n81 146.341
R914 VCC.n265 VCC.n264 146.341
R915 VCC.n265 VCC.n3 146.341
R916 VCC.n4 VCC.n3 146.341
R917 VCC.n5 VCC.n4 146.341
R918 VCC.n276 VCC.n5 146.341
R919 VCC.n276 VCC.n8 146.341
R920 VCC.n9 VCC.n8 146.341
R921 VCC.n10 VCC.n9 146.341
R922 VCC.n287 VCC.n10 146.341
R923 VCC.n287 VCC.n13 146.341
R924 VCC.n14 VCC.n13 146.341
R925 VCC.n15 VCC.n14 146.341
R926 VCC.n298 VCC.n15 146.341
R927 VCC.n298 VCC.n18 146.341
R928 VCC.n19 VCC.n18 146.341
R929 VCC.n20 VCC.n19 146.341
R930 VCC.n309 VCC.n20 146.341
R931 VCC.n309 VCC.n23 146.341
R932 VCC.n24 VCC.n23 146.341
R933 VCC.n25 VCC.n24 146.341
R934 VCC.n322 VCC.n25 146.341
R935 VCC.n322 VCC.n28 146.341
R936 VCC.n29 VCC.n28 146.341
R937 VCC.n30 VCC.n29 146.341
R938 VCC.n42 VCC.t5 143.969
R939 VCC.n142 VCC.t8 143.969
R940 VCC.n181 VCC.n139 131.757
R941 VCC.n358 VCC.n33 131.757
R942 VCC.n359 VCC.n32 99.5127
R943 VCC.n356 VCC.n40 99.5127
R944 VCC.n352 VCC.n351 99.5127
R945 VCC.n348 VCC.n347 99.5127
R946 VCC.n344 VCC.n343 99.5127
R947 VCC.n340 VCC.n339 99.5127
R948 VCC.n336 VCC.n335 99.5127
R949 VCC.n175 VCC.n173 99.5127
R950 VCC.n173 VCC.n144 99.5127
R951 VCC.n169 VCC.n167 99.5127
R952 VCC.n165 VCC.n146 99.5127
R953 VCC.n161 VCC.n159 99.5127
R954 VCC.n157 VCC.n148 99.5127
R955 VCC.n153 VCC.n151 99.5127
R956 VCC.n42 VCC.n41 76.9944
R957 VCC.n142 VCC.n141 76.9944
R958 VCC.n358 VCC.n34 72.8958
R959 VCC.n358 VCC.n35 72.8958
R960 VCC.n358 VCC.n36 72.8958
R961 VCC.n358 VCC.n37 72.8958
R962 VCC.n358 VCC.n38 72.8958
R963 VCC.n358 VCC.n39 72.8958
R964 VCC.n358 VCC.n357 72.8958
R965 VCC.n174 VCC.n139 72.8958
R966 VCC.n168 VCC.n139 72.8958
R967 VCC.n166 VCC.n139 72.8958
R968 VCC.n160 VCC.n139 72.8958
R969 VCC.n158 VCC.n139 72.8958
R970 VCC.n152 VCC.n139 72.8958
R971 VCC.n150 VCC.n139 72.8958
R972 VCC.n181 VCC.n134 67.5681
R973 VCC.n190 VCC.n134 67.5681
R974 VCC.n190 VCC.n189 67.5681
R975 VCC.n198 VCC.n123 67.5681
R976 VCC.n206 VCC.n123 67.5681
R977 VCC.n206 VCC.n117 67.5681
R978 VCC.n214 VCC.n117 67.5681
R979 VCC.n214 VCC.n111 67.5681
R980 VCC.n222 VCC.n111 67.5681
R981 VCC.n222 VCC.n105 67.5681
R982 VCC.n230 VCC.n105 67.5681
R983 VCC.n230 VCC.n98 67.5681
R984 VCC.n239 VCC.n98 67.5681
R985 VCC.n247 VCC.n92 67.5681
R986 VCC.n247 VCC.n86 67.5681
R987 VCC.n257 VCC.n86 67.5681
R988 VCC.n257 VCC.n256 67.5681
R989 VCC.n256 VCC.n80 67.5681
R990 VCC.n266 VCC.n80 67.5681
R991 VCC.n266 VCC.t10 67.5681
R992 VCC.n274 VCC.t10 67.5681
R993 VCC.n275 VCC.n274 67.5681
R994 VCC.n277 VCC.n275 67.5681
R995 VCC.n277 VCC.n69 67.5681
R996 VCC.n285 VCC.n69 67.5681
R997 VCC.n286 VCC.n285 67.5681
R998 VCC.n288 VCC.n286 67.5681
R999 VCC.n296 VCC.n63 67.5681
R1000 VCC.n297 VCC.n296 67.5681
R1001 VCC.n299 VCC.n297 67.5681
R1002 VCC.n299 VCC.n57 67.5681
R1003 VCC.n307 VCC.n57 67.5681
R1004 VCC.n308 VCC.n307 67.5681
R1005 VCC.n310 VCC.n308 67.5681
R1006 VCC.n310 VCC.n51 67.5681
R1007 VCC.n318 VCC.n51 67.5681
R1008 VCC.n319 VCC.n318 67.5681
R1009 VCC.n323 VCC.n321 67.5681
R1010 VCC.n321 VCC.n320 67.5681
R1011 VCC.n320 VCC.n33 67.5681
R1012 VCC.n189 VCC.t7 63.514
R1013 VCC.t0 VCC.n92 63.514
R1014 VCC.n288 VCC.t1 63.514
R1015 VCC.n323 VCC.t3 63.514
R1016 VCC.n357 VCC.n356 39.2114
R1017 VCC.n352 VCC.n39 39.2114
R1018 VCC.n348 VCC.n38 39.2114
R1019 VCC.n344 VCC.n37 39.2114
R1020 VCC.n340 VCC.n36 39.2114
R1021 VCC.n336 VCC.n35 39.2114
R1022 VCC.n332 VCC.n34 39.2114
R1023 VCC.n174 VCC.n140 39.2114
R1024 VCC.n168 VCC.n144 39.2114
R1025 VCC.n167 VCC.n166 39.2114
R1026 VCC.n160 VCC.n146 39.2114
R1027 VCC.n159 VCC.n158 39.2114
R1028 VCC.n152 VCC.n148 39.2114
R1029 VCC.n151 VCC.n150 39.2114
R1030 VCC.n335 VCC.n34 39.2114
R1031 VCC.n339 VCC.n35 39.2114
R1032 VCC.n343 VCC.n36 39.2114
R1033 VCC.n347 VCC.n37 39.2114
R1034 VCC.n351 VCC.n38 39.2114
R1035 VCC.n40 VCC.n39 39.2114
R1036 VCC.n357 VCC.n32 39.2114
R1037 VCC.n175 VCC.n174 39.2114
R1038 VCC.n169 VCC.n168 39.2114
R1039 VCC.n166 VCC.n165 39.2114
R1040 VCC.n161 VCC.n160 39.2114
R1041 VCC.n158 VCC.n157 39.2114
R1042 VCC.n153 VCC.n152 39.2114
R1043 VCC.n150 VCC.n138 39.2114
R1044 VCC.n43 VCC.n42 29.2853
R1045 VCC.n143 VCC.n142 29.2853
R1046 VCC.n361 VCC.n360 28.9539
R1047 VCC.n333 VCC.n44 28.9539
R1048 VCC.n178 VCC.n177 28.9539
R1049 VCC.n184 VCC.n137 28.9539
R1050 VCC.n183 VCC.n136 19.3944
R1051 VCC.n187 VCC.n136 19.3944
R1052 VCC.n187 VCC.n127 19.3944
R1053 VCC.n200 VCC.n127 19.3944
R1054 VCC.n200 VCC.n125 19.3944
R1055 VCC.n204 VCC.n125 19.3944
R1056 VCC.n204 VCC.n115 19.3944
R1057 VCC.n216 VCC.n115 19.3944
R1058 VCC.n216 VCC.n113 19.3944
R1059 VCC.n220 VCC.n113 19.3944
R1060 VCC.n220 VCC.n103 19.3944
R1061 VCC.n232 VCC.n103 19.3944
R1062 VCC.n232 VCC.n100 19.3944
R1063 VCC.n237 VCC.n100 19.3944
R1064 VCC.n237 VCC.n101 19.3944
R1065 VCC.n101 VCC.n90 19.3944
R1066 VCC.n250 VCC.n90 19.3944
R1067 VCC.n250 VCC.n88 19.3944
R1068 VCC.n254 VCC.n88 19.3944
R1069 VCC.n254 VCC.n78 19.3944
R1070 VCC.n268 VCC.n78 19.3944
R1071 VCC.n268 VCC.n76 19.3944
R1072 VCC.n272 VCC.n76 19.3944
R1073 VCC.n272 VCC.n73 19.3944
R1074 VCC.n279 VCC.n73 19.3944
R1075 VCC.n279 VCC.n71 19.3944
R1076 VCC.n283 VCC.n71 19.3944
R1077 VCC.n283 VCC.n67 19.3944
R1078 VCC.n290 VCC.n67 19.3944
R1079 VCC.n290 VCC.n65 19.3944
R1080 VCC.n294 VCC.n65 19.3944
R1081 VCC.n294 VCC.n61 19.3944
R1082 VCC.n301 VCC.n61 19.3944
R1083 VCC.n301 VCC.n59 19.3944
R1084 VCC.n305 VCC.n59 19.3944
R1085 VCC.n305 VCC.n55 19.3944
R1086 VCC.n312 VCC.n55 19.3944
R1087 VCC.n312 VCC.n53 19.3944
R1088 VCC.n316 VCC.n53 19.3944
R1089 VCC.n316 VCC.n48 19.3944
R1090 VCC.n325 VCC.n48 19.3944
R1091 VCC.n325 VCC.n46 19.3944
R1092 VCC.n329 VCC.n46 19.3944
R1093 VCC.n330 VCC.n329 19.3944
R1094 VCC.n179 VCC.n132 19.3944
R1095 VCC.n192 VCC.n132 19.3944
R1096 VCC.n192 VCC.n130 19.3944
R1097 VCC.n196 VCC.n130 19.3944
R1098 VCC.n196 VCC.n121 19.3944
R1099 VCC.n208 VCC.n121 19.3944
R1100 VCC.n208 VCC.n119 19.3944
R1101 VCC.n212 VCC.n119 19.3944
R1102 VCC.n212 VCC.n109 19.3944
R1103 VCC.n224 VCC.n109 19.3944
R1104 VCC.n224 VCC.n107 19.3944
R1105 VCC.n228 VCC.n107 19.3944
R1106 VCC.n228 VCC.n96 19.3944
R1107 VCC.n241 VCC.n96 19.3944
R1108 VCC.n241 VCC.n94 19.3944
R1109 VCC.n245 VCC.n94 19.3944
R1110 VCC.n245 VCC.n84 19.3944
R1111 VCC.n259 VCC.n84 19.3944
R1112 VCC.n259 VCC.n82 19.3944
R1113 VCC.n263 VCC.n82 19.3944
R1114 VCC.n263 VCC.n2 19.3944
R1115 VCC.n394 VCC.n2 19.3944
R1116 VCC.n394 VCC.n393 19.3944
R1117 VCC.n393 VCC.n392 19.3944
R1118 VCC.n392 VCC.n6 19.3944
R1119 VCC.n388 VCC.n6 19.3944
R1120 VCC.n388 VCC.n387 19.3944
R1121 VCC.n387 VCC.n386 19.3944
R1122 VCC.n386 VCC.n11 19.3944
R1123 VCC.n382 VCC.n11 19.3944
R1124 VCC.n382 VCC.n381 19.3944
R1125 VCC.n381 VCC.n380 19.3944
R1126 VCC.n380 VCC.n16 19.3944
R1127 VCC.n376 VCC.n16 19.3944
R1128 VCC.n376 VCC.n375 19.3944
R1129 VCC.n375 VCC.n374 19.3944
R1130 VCC.n374 VCC.n21 19.3944
R1131 VCC.n370 VCC.n21 19.3944
R1132 VCC.n370 VCC.n369 19.3944
R1133 VCC.n369 VCC.n368 19.3944
R1134 VCC.n368 VCC.n26 19.3944
R1135 VCC.n364 VCC.n26 19.3944
R1136 VCC.n364 VCC.n363 19.3944
R1137 VCC.n363 VCC.n362 19.3944
R1138 VCC.n360 VCC.n31 10.6151
R1139 VCC.n355 VCC.n354 10.6151
R1140 VCC.n354 VCC.n353 10.6151
R1141 VCC.n353 VCC.n350 10.6151
R1142 VCC.n350 VCC.n349 10.6151
R1143 VCC.n349 VCC.n346 10.6151
R1144 VCC.n346 VCC.n345 10.6151
R1145 VCC.n345 VCC.n342 10.6151
R1146 VCC.n342 VCC.n341 10.6151
R1147 VCC.n341 VCC.n338 10.6151
R1148 VCC.n338 VCC.n337 10.6151
R1149 VCC.n337 VCC.n334 10.6151
R1150 VCC.n334 VCC.n333 10.6151
R1151 VCC.n177 VCC.n176 10.6151
R1152 VCC.n172 VCC.n171 10.6151
R1153 VCC.n171 VCC.n170 10.6151
R1154 VCC.n170 VCC.n145 10.6151
R1155 VCC.n164 VCC.n145 10.6151
R1156 VCC.n164 VCC.n163 10.6151
R1157 VCC.n163 VCC.n162 10.6151
R1158 VCC.n162 VCC.n147 10.6151
R1159 VCC.n156 VCC.n147 10.6151
R1160 VCC.n156 VCC.n155 10.6151
R1161 VCC.n155 VCC.n154 10.6151
R1162 VCC.n154 VCC.n149 10.6151
R1163 VCC.n149 VCC.n137 10.6151
R1164 VCC.n393 VCC.n0 9.3005
R1165 VCC.n392 VCC.n391 9.3005
R1166 VCC.n390 VCC.n6 9.3005
R1167 VCC.n389 VCC.n388 9.3005
R1168 VCC.n387 VCC.n7 9.3005
R1169 VCC.n386 VCC.n385 9.3005
R1170 VCC.n384 VCC.n11 9.3005
R1171 VCC.n383 VCC.n382 9.3005
R1172 VCC.n381 VCC.n12 9.3005
R1173 VCC.n380 VCC.n379 9.3005
R1174 VCC.n378 VCC.n16 9.3005
R1175 VCC.n377 VCC.n376 9.3005
R1176 VCC.n375 VCC.n17 9.3005
R1177 VCC.n374 VCC.n373 9.3005
R1178 VCC.n372 VCC.n21 9.3005
R1179 VCC.n371 VCC.n370 9.3005
R1180 VCC.n369 VCC.n22 9.3005
R1181 VCC.n368 VCC.n367 9.3005
R1182 VCC.n366 VCC.n26 9.3005
R1183 VCC.n365 VCC.n364 9.3005
R1184 VCC.n363 VCC.n27 9.3005
R1185 VCC.n362 VCC.n361 9.3005
R1186 VCC.n185 VCC.n136 9.3005
R1187 VCC.n187 VCC.n186 9.3005
R1188 VCC.n127 VCC.n126 9.3005
R1189 VCC.n201 VCC.n200 9.3005
R1190 VCC.n202 VCC.n125 9.3005
R1191 VCC.n204 VCC.n203 9.3005
R1192 VCC.n115 VCC.n114 9.3005
R1193 VCC.n217 VCC.n216 9.3005
R1194 VCC.n218 VCC.n113 9.3005
R1195 VCC.n220 VCC.n219 9.3005
R1196 VCC.n103 VCC.n102 9.3005
R1197 VCC.n233 VCC.n232 9.3005
R1198 VCC.n234 VCC.n100 9.3005
R1199 VCC.n237 VCC.n236 9.3005
R1200 VCC.n235 VCC.n101 9.3005
R1201 VCC.n90 VCC.n89 9.3005
R1202 VCC.n251 VCC.n250 9.3005
R1203 VCC.n252 VCC.n88 9.3005
R1204 VCC.n254 VCC.n253 9.3005
R1205 VCC.n78 VCC.n77 9.3005
R1206 VCC.n269 VCC.n268 9.3005
R1207 VCC.n270 VCC.n76 9.3005
R1208 VCC.n272 VCC.n271 9.3005
R1209 VCC.n73 VCC.n72 9.3005
R1210 VCC.n280 VCC.n279 9.3005
R1211 VCC.n281 VCC.n71 9.3005
R1212 VCC.n283 VCC.n282 9.3005
R1213 VCC.n67 VCC.n66 9.3005
R1214 VCC.n291 VCC.n290 9.3005
R1215 VCC.n292 VCC.n65 9.3005
R1216 VCC.n294 VCC.n293 9.3005
R1217 VCC.n61 VCC.n60 9.3005
R1218 VCC.n302 VCC.n301 9.3005
R1219 VCC.n303 VCC.n59 9.3005
R1220 VCC.n305 VCC.n304 9.3005
R1221 VCC.n55 VCC.n54 9.3005
R1222 VCC.n313 VCC.n312 9.3005
R1223 VCC.n314 VCC.n53 9.3005
R1224 VCC.n316 VCC.n315 9.3005
R1225 VCC.n48 VCC.n47 9.3005
R1226 VCC.n326 VCC.n325 9.3005
R1227 VCC.n327 VCC.n46 9.3005
R1228 VCC.n329 VCC.n328 9.3005
R1229 VCC.n330 VCC.n44 9.3005
R1230 VCC.n184 VCC.n183 9.3005
R1231 VCC.n179 VCC.n178 9.3005
R1232 VCC.n132 VCC.n131 9.3005
R1233 VCC.n193 VCC.n192 9.3005
R1234 VCC.n194 VCC.n130 9.3005
R1235 VCC.n196 VCC.n195 9.3005
R1236 VCC.n121 VCC.n120 9.3005
R1237 VCC.n209 VCC.n208 9.3005
R1238 VCC.n210 VCC.n119 9.3005
R1239 VCC.n212 VCC.n211 9.3005
R1240 VCC.n109 VCC.n108 9.3005
R1241 VCC.n225 VCC.n224 9.3005
R1242 VCC.n226 VCC.n107 9.3005
R1243 VCC.n228 VCC.n227 9.3005
R1244 VCC.n96 VCC.n95 9.3005
R1245 VCC.n242 VCC.n241 9.3005
R1246 VCC.n243 VCC.n94 9.3005
R1247 VCC.n245 VCC.n244 9.3005
R1248 VCC.n84 VCC.n83 9.3005
R1249 VCC.n260 VCC.n259 9.3005
R1250 VCC.n261 VCC.n82 9.3005
R1251 VCC.n263 VCC.n262 9.3005
R1252 VCC.n2 VCC.n1 9.3005
R1253 VCC.n395 VCC.n394 9.3005
R1254 VCC.n43 VCC.n31 7.33709
R1255 VCC.n176 VCC.n143 7.33709
R1256 VCC.n198 VCC.t7 4.05455
R1257 VCC.n239 VCC.t0 4.05455
R1258 VCC.t1 VCC.n63 4.05455
R1259 VCC.t3 VCC.n319 4.05455
R1260 VCC.n355 VCC.n43 3.27855
R1261 VCC.n172 VCC.n143 3.27855
R1262 VCC.n391 VCC.n0 0.152939
R1263 VCC.n391 VCC.n390 0.152939
R1264 VCC.n390 VCC.n389 0.152939
R1265 VCC.n389 VCC.n7 0.152939
R1266 VCC.n385 VCC.n7 0.152939
R1267 VCC.n385 VCC.n384 0.152939
R1268 VCC.n384 VCC.n383 0.152939
R1269 VCC.n383 VCC.n12 0.152939
R1270 VCC.n379 VCC.n12 0.152939
R1271 VCC.n379 VCC.n378 0.152939
R1272 VCC.n378 VCC.n377 0.152939
R1273 VCC.n377 VCC.n17 0.152939
R1274 VCC.n373 VCC.n17 0.152939
R1275 VCC.n373 VCC.n372 0.152939
R1276 VCC.n372 VCC.n371 0.152939
R1277 VCC.n371 VCC.n22 0.152939
R1278 VCC.n367 VCC.n22 0.152939
R1279 VCC.n367 VCC.n366 0.152939
R1280 VCC.n366 VCC.n365 0.152939
R1281 VCC.n365 VCC.n27 0.152939
R1282 VCC.n361 VCC.n27 0.152939
R1283 VCC.n185 VCC.n184 0.152939
R1284 VCC.n186 VCC.n185 0.152939
R1285 VCC.n186 VCC.n126 0.152939
R1286 VCC.n201 VCC.n126 0.152939
R1287 VCC.n202 VCC.n201 0.152939
R1288 VCC.n203 VCC.n202 0.152939
R1289 VCC.n203 VCC.n114 0.152939
R1290 VCC.n217 VCC.n114 0.152939
R1291 VCC.n218 VCC.n217 0.152939
R1292 VCC.n219 VCC.n218 0.152939
R1293 VCC.n219 VCC.n102 0.152939
R1294 VCC.n233 VCC.n102 0.152939
R1295 VCC.n234 VCC.n233 0.152939
R1296 VCC.n236 VCC.n234 0.152939
R1297 VCC.n236 VCC.n235 0.152939
R1298 VCC.n235 VCC.n89 0.152939
R1299 VCC.n251 VCC.n89 0.152939
R1300 VCC.n252 VCC.n251 0.152939
R1301 VCC.n253 VCC.n252 0.152939
R1302 VCC.n253 VCC.n77 0.152939
R1303 VCC.n269 VCC.n77 0.152939
R1304 VCC.n270 VCC.n269 0.152939
R1305 VCC.n271 VCC.n270 0.152939
R1306 VCC.n271 VCC.n72 0.152939
R1307 VCC.n280 VCC.n72 0.152939
R1308 VCC.n281 VCC.n280 0.152939
R1309 VCC.n282 VCC.n281 0.152939
R1310 VCC.n282 VCC.n66 0.152939
R1311 VCC.n291 VCC.n66 0.152939
R1312 VCC.n292 VCC.n291 0.152939
R1313 VCC.n293 VCC.n292 0.152939
R1314 VCC.n293 VCC.n60 0.152939
R1315 VCC.n302 VCC.n60 0.152939
R1316 VCC.n303 VCC.n302 0.152939
R1317 VCC.n304 VCC.n303 0.152939
R1318 VCC.n304 VCC.n54 0.152939
R1319 VCC.n313 VCC.n54 0.152939
R1320 VCC.n314 VCC.n313 0.152939
R1321 VCC.n315 VCC.n314 0.152939
R1322 VCC.n315 VCC.n47 0.152939
R1323 VCC.n326 VCC.n47 0.152939
R1324 VCC.n327 VCC.n326 0.152939
R1325 VCC.n328 VCC.n327 0.152939
R1326 VCC.n328 VCC.n44 0.152939
R1327 VCC.n178 VCC.n131 0.152939
R1328 VCC.n193 VCC.n131 0.152939
R1329 VCC.n194 VCC.n193 0.152939
R1330 VCC.n195 VCC.n194 0.152939
R1331 VCC.n195 VCC.n120 0.152939
R1332 VCC.n209 VCC.n120 0.152939
R1333 VCC.n210 VCC.n209 0.152939
R1334 VCC.n211 VCC.n210 0.152939
R1335 VCC.n211 VCC.n108 0.152939
R1336 VCC.n225 VCC.n108 0.152939
R1337 VCC.n226 VCC.n225 0.152939
R1338 VCC.n227 VCC.n226 0.152939
R1339 VCC.n227 VCC.n95 0.152939
R1340 VCC.n242 VCC.n95 0.152939
R1341 VCC.n243 VCC.n242 0.152939
R1342 VCC.n244 VCC.n243 0.152939
R1343 VCC.n244 VCC.n83 0.152939
R1344 VCC.n260 VCC.n83 0.152939
R1345 VCC.n261 VCC.n260 0.152939
R1346 VCC.n262 VCC.n261 0.152939
R1347 VCC.n262 VCC.n1 0.152939
R1348 VCC.n395 VCC.n1 0.13922
R1349 VCC VCC.n0 0.0767195
R1350 VCC VCC.n395 0.063
R1351 VGP.n18 VGP.n17 161.3
R1352 VGP.n16 VGP.n1 161.3
R1353 VGP.n15 VGP.n14 161.3
R1354 VGP.n13 VGP.n2 161.3
R1355 VGP.n12 VGP.n11 161.3
R1356 VGP.n10 VGP.n3 161.3
R1357 VGP.n9 VGP.n8 161.3
R1358 VGP.n7 VGP.n4 161.3
R1359 VGP.n19 VGP.n0 79.4252
R1360 VGP.n6 VGP.n5 62.5662
R1361 VGP.n11 VGP.n2 56.5617
R1362 VGP.n6 VGP.t0 52.9281
R1363 VGP.n11 VGP.n10 24.5923
R1364 VGP.n10 VGP.n9 24.5923
R1365 VGP.n9 VGP.n4 24.5923
R1366 VGP.n17 VGP.n16 24.5923
R1367 VGP.n16 VGP.n15 24.5923
R1368 VGP.n15 VGP.n2 24.5923
R1369 VGP.n5 VGP.t2 19.3335
R1370 VGP.n0 VGP.t1 19.3335
R1371 VGP.n5 VGP.n4 12.2964
R1372 VGP.n17 VGP.n0 10.8209
R1373 VGP.n7 VGP.n6 3.11924
R1374 VGP VGP.n19 0.369343
R1375 VGP.n19 VGP.n18 0.354861
R1376 VGP.n18 VGP.n1 0.189894
R1377 VGP.n14 VGP.n1 0.189894
R1378 VGP.n14 VGP.n13 0.189894
R1379 VGP.n13 VGP.n12 0.189894
R1380 VGP.n12 VGP.n3 0.189894
R1381 VGP.n8 VGP.n3 0.189894
R1382 VGP.n8 VGP.n7 0.189894
C0 VGN VOUT 0.940727f
C1 VIN VOUT 3.02959f
C2 VGN VCC 0.020914f
C3 VIN VCC 0.723793f
C4 VOUT VGP 0.842585f
C5 VGP VCC 4.3411f
C6 VIN VGN 1.22517f
C7 VGN VGP 0.02055f
C8 VIN VGP 1.42528f
C9 VOUT VCC 1.75974f
C10 VGN VSS 3.00185f
C11 VOUT VSS 2.010797f
C12 VIN VSS 1.570576f
C13 VGP VSS 1.507077f
C14 VCC VSS 24.475286f
C15 VGP.t1 VSS 0.655412f
C16 VGP.n0 VSS 0.369237f
C17 VGP.n1 VSS 0.024839f
C18 VGP.n2 VSS 0.037138f
C19 VGP.n3 VSS 0.024839f
C20 VGP.n4 VSS 0.034692f
C21 VGP.t0 VSS 0.946909f
C22 VGP.t2 VSS 0.655412f
C23 VGP.n5 VSS 0.355523f
C24 VGP.n6 VSS 0.367229f
C25 VGP.n7 VSS 0.310462f
C26 VGP.n8 VSS 0.024839f
C27 VGP.n9 VSS 0.046061f
C28 VGP.n10 VSS 0.046061f
C29 VGP.n11 VSS 0.035076f
C30 VGP.n12 VSS 0.024839f
C31 VGP.n13 VSS 0.024839f
C32 VGP.n14 VSS 0.024839f
C33 VGP.n15 VSS 0.046061f
C34 VGP.n16 VSS 0.046061f
C35 VGP.n17 VSS 0.033327f
C36 VGP.n18 VSS 0.040083f
C37 VGP.n19 VSS 0.080594f
C38 VCC.n0 VSS 0.002416f
C39 VCC.n1 VSS 0.003222f
C40 VCC.n2 VSS 0.002593f
C41 VCC.n3 VSS 0.003222f
C42 VCC.n4 VSS 0.003222f
C43 VCC.n5 VSS 0.003222f
C44 VCC.n6 VSS 0.002593f
C45 VCC.n7 VSS 0.003222f
C46 VCC.n8 VSS 0.003222f
C47 VCC.n9 VSS 0.003222f
C48 VCC.n10 VSS 0.003222f
C49 VCC.n11 VSS 0.002593f
C50 VCC.n12 VSS 0.003222f
C51 VCC.n13 VSS 0.003222f
C52 VCC.n14 VSS 0.003222f
C53 VCC.n15 VSS 0.003222f
C54 VCC.n16 VSS 0.002593f
C55 VCC.n17 VSS 0.003222f
C56 VCC.n18 VSS 0.003222f
C57 VCC.n19 VSS 0.003222f
C58 VCC.n20 VSS 0.003222f
C59 VCC.n21 VSS 0.002593f
C60 VCC.n22 VSS 0.003222f
C61 VCC.n23 VSS 0.003222f
C62 VCC.n24 VSS 0.003222f
C63 VCC.n25 VSS 0.003222f
C64 VCC.n26 VSS 0.002593f
C65 VCC.n27 VSS 0.003222f
C66 VCC.n28 VSS 0.003222f
C67 VCC.n29 VSS 0.003222f
C68 VCC.n30 VSS 0.006483f
C69 VCC.n31 VSS 0.001852f
C70 VCC.n32 VSS 0.002191f
C71 VCC.n33 VSS 0.081476f
C72 VCC.n40 VSS 0.002191f
C73 VCC.t5 VSS 0.021806f
C74 VCC.t4 VSS 0.028264f
C75 VCC.t2 VSS 0.163172f
C76 VCC.n41 VSS 0.027939f
C77 VCC.n42 VSS 0.019634f
C78 VCC.n43 VSS 0.003053f
C79 VCC.n44 VSS 0.011386f
C80 VCC.n45 VSS 0.003222f
C81 VCC.n46 VSS 0.002593f
C82 VCC.n47 VSS 0.003222f
C83 VCC.n48 VSS 0.002593f
C84 VCC.n49 VSS 0.003222f
C85 VCC.n50 VSS 0.003222f
C86 VCC.n51 VSS 0.055238f
C87 VCC.n52 VSS 0.003222f
C88 VCC.n53 VSS 0.002593f
C89 VCC.n54 VSS 0.003222f
C90 VCC.n55 VSS 0.002593f
C91 VCC.n56 VSS 0.003222f
C92 VCC.n57 VSS 0.055238f
C93 VCC.n58 VSS 0.003222f
C94 VCC.n59 VSS 0.002593f
C95 VCC.n60 VSS 0.003222f
C96 VCC.n61 VSS 0.002593f
C97 VCC.n62 VSS 0.003222f
C98 VCC.n63 VSS 0.029276f
C99 VCC.n64 VSS 0.003222f
C100 VCC.n65 VSS 0.002593f
C101 VCC.n66 VSS 0.003222f
C102 VCC.n67 VSS 0.002593f
C103 VCC.n68 VSS 0.003222f
C104 VCC.n69 VSS 0.055238f
C105 VCC.n70 VSS 0.003222f
C106 VCC.n71 VSS 0.002593f
C107 VCC.n72 VSS 0.003222f
C108 VCC.n73 VSS 0.002593f
C109 VCC.n74 VSS 0.003222f
C110 VCC.t10 VSS 0.055238f
C111 VCC.n75 VSS 0.003222f
C112 VCC.n76 VSS 0.002593f
C113 VCC.n77 VSS 0.003222f
C114 VCC.n78 VSS 0.002593f
C115 VCC.n79 VSS 0.003222f
C116 VCC.n80 VSS 0.055238f
C117 VCC.n81 VSS 0.003222f
C118 VCC.n82 VSS 0.002593f
C119 VCC.n83 VSS 0.003222f
C120 VCC.n84 VSS 0.002593f
C121 VCC.n85 VSS 0.003222f
C122 VCC.n86 VSS 0.055238f
C123 VCC.n87 VSS 0.003222f
C124 VCC.n88 VSS 0.002593f
C125 VCC.n89 VSS 0.003222f
C126 VCC.n90 VSS 0.002593f
C127 VCC.n91 VSS 0.003222f
C128 VCC.n92 VSS 0.053581f
C129 VCC.n93 VSS 0.003222f
C130 VCC.n94 VSS 0.002593f
C131 VCC.n95 VSS 0.003222f
C132 VCC.n96 VSS 0.002593f
C133 VCC.n97 VSS 0.003222f
C134 VCC.n98 VSS 0.055238f
C135 VCC.n99 VSS 0.003222f
C136 VCC.n100 VSS 0.002593f
C137 VCC.n101 VSS 0.002593f
C138 VCC.n102 VSS 0.003222f
C139 VCC.n103 VSS 0.002593f
C140 VCC.n104 VSS 0.003222f
C141 VCC.n105 VSS 0.055238f
C142 VCC.n106 VSS 0.003222f
C143 VCC.n107 VSS 0.002593f
C144 VCC.n108 VSS 0.003222f
C145 VCC.n109 VSS 0.002593f
C146 VCC.n110 VSS 0.003222f
C147 VCC.n111 VSS 0.055238f
C148 VCC.n112 VSS 0.003222f
C149 VCC.n113 VSS 0.002593f
C150 VCC.n114 VSS 0.003222f
C151 VCC.n115 VSS 0.002593f
C152 VCC.n116 VSS 0.003222f
C153 VCC.n117 VSS 0.055238f
C154 VCC.n118 VSS 0.003222f
C155 VCC.n119 VSS 0.002593f
C156 VCC.n120 VSS 0.003222f
C157 VCC.n121 VSS 0.002593f
C158 VCC.n122 VSS 0.003222f
C159 VCC.n123 VSS 0.055238f
C160 VCC.n124 VSS 0.003222f
C161 VCC.n125 VSS 0.002593f
C162 VCC.n126 VSS 0.003222f
C163 VCC.n127 VSS 0.002593f
C164 VCC.n128 VSS 0.003222f
C165 VCC.t7 VSS 0.027619f
C166 VCC.n129 VSS 0.003222f
C167 VCC.n130 VSS 0.002593f
C168 VCC.n131 VSS 0.003222f
C169 VCC.n132 VSS 0.002593f
C170 VCC.n133 VSS 0.003222f
C171 VCC.n134 VSS 0.055238f
C172 VCC.n135 VSS 0.003222f
C173 VCC.n136 VSS 0.002593f
C174 VCC.n137 VSS 0.004238f
C175 VCC.n138 VSS 0.0065f
C176 VCC.n139 VSS 0.110752f
C177 VCC.n140 VSS 0.0065f
C178 VCC.t8 VSS 0.021806f
C179 VCC.t9 VSS 0.028264f
C180 VCC.t6 VSS 0.163172f
C181 VCC.n141 VSS 0.027939f
C182 VCC.n142 VSS 0.019634f
C183 VCC.n143 VSS 0.003053f
C184 VCC.n144 VSS 0.002191f
C185 VCC.n145 VSS 0.002191f
C186 VCC.n146 VSS 0.002191f
C187 VCC.n147 VSS 0.002191f
C188 VCC.n148 VSS 0.002191f
C189 VCC.n149 VSS 0.002191f
C190 VCC.n151 VSS 0.002191f
C191 VCC.n153 VSS 0.002191f
C192 VCC.n154 VSS 0.002191f
C193 VCC.n155 VSS 0.002191f
C194 VCC.n156 VSS 0.002191f
C195 VCC.n157 VSS 0.002191f
C196 VCC.n159 VSS 0.002191f
C197 VCC.n161 VSS 0.002191f
C198 VCC.n162 VSS 0.002191f
C199 VCC.n163 VSS 0.002191f
C200 VCC.n164 VSS 0.002191f
C201 VCC.n165 VSS 0.002191f
C202 VCC.n167 VSS 0.002191f
C203 VCC.n169 VSS 0.002191f
C204 VCC.n170 VSS 0.002191f
C205 VCC.n171 VSS 0.002191f
C206 VCC.n172 VSS 0.001434f
C207 VCC.n173 VSS 0.002191f
C208 VCC.n175 VSS 0.002191f
C209 VCC.n176 VSS 0.001852f
C210 VCC.n177 VSS 0.004238f
C211 VCC.n178 VSS 0.011386f
C212 VCC.n179 VSS 0.002152f
C213 VCC.n180 VSS 0.006483f
C214 VCC.n181 VSS 0.081476f
C215 VCC.n182 VSS 0.006483f
C216 VCC.n183 VSS 0.002152f
C217 VCC.n184 VSS 0.011386f
C218 VCC.n185 VSS 0.003222f
C219 VCC.n186 VSS 0.003222f
C220 VCC.n187 VSS 0.002593f
C221 VCC.n188 VSS 0.003222f
C222 VCC.n189 VSS 0.053581f
C223 VCC.n190 VSS 0.055238f
C224 VCC.n191 VSS 0.003222f
C225 VCC.n192 VSS 0.002593f
C226 VCC.n193 VSS 0.003222f
C227 VCC.n194 VSS 0.003222f
C228 VCC.n195 VSS 0.003222f
C229 VCC.n196 VSS 0.002593f
C230 VCC.n197 VSS 0.003222f
C231 VCC.n198 VSS 0.029276f
C232 VCC.n199 VSS 0.003222f
C233 VCC.n200 VSS 0.002593f
C234 VCC.n201 VSS 0.003222f
C235 VCC.n202 VSS 0.003222f
C236 VCC.n203 VSS 0.003222f
C237 VCC.n204 VSS 0.002593f
C238 VCC.n205 VSS 0.003222f
C239 VCC.n206 VSS 0.055238f
C240 VCC.n207 VSS 0.003222f
C241 VCC.n208 VSS 0.002593f
C242 VCC.n209 VSS 0.003222f
C243 VCC.n210 VSS 0.003222f
C244 VCC.n211 VSS 0.003222f
C245 VCC.n212 VSS 0.002593f
C246 VCC.n213 VSS 0.003222f
C247 VCC.n214 VSS 0.055238f
C248 VCC.n215 VSS 0.003222f
C249 VCC.n216 VSS 0.002593f
C250 VCC.n217 VSS 0.003222f
C251 VCC.n218 VSS 0.003222f
C252 VCC.n219 VSS 0.003222f
C253 VCC.n220 VSS 0.002593f
C254 VCC.n221 VSS 0.003222f
C255 VCC.n222 VSS 0.055238f
C256 VCC.n223 VSS 0.003222f
C257 VCC.n224 VSS 0.002593f
C258 VCC.n225 VSS 0.003222f
C259 VCC.n226 VSS 0.003222f
C260 VCC.n227 VSS 0.003222f
C261 VCC.n228 VSS 0.002593f
C262 VCC.n229 VSS 0.003222f
C263 VCC.n230 VSS 0.055238f
C264 VCC.n231 VSS 0.003222f
C265 VCC.n232 VSS 0.002593f
C266 VCC.n233 VSS 0.003222f
C267 VCC.n234 VSS 0.003222f
C268 VCC.n235 VSS 0.003222f
C269 VCC.n236 VSS 0.003222f
C270 VCC.n237 VSS 0.002593f
C271 VCC.n238 VSS 0.003222f
C272 VCC.t0 VSS 0.027619f
C273 VCC.n239 VSS 0.029276f
C274 VCC.n240 VSS 0.003222f
C275 VCC.n241 VSS 0.002593f
C276 VCC.n242 VSS 0.003222f
C277 VCC.n243 VSS 0.003222f
C278 VCC.n244 VSS 0.003222f
C279 VCC.n245 VSS 0.002593f
C280 VCC.n246 VSS 0.003222f
C281 VCC.n247 VSS 0.055238f
C282 VCC.n248 VSS 0.003222f
C283 VCC.n249 VSS 0.003222f
C284 VCC.n250 VSS 0.002593f
C285 VCC.n251 VSS 0.003222f
C286 VCC.n252 VSS 0.003222f
C287 VCC.n253 VSS 0.003222f
C288 VCC.n254 VSS 0.002593f
C289 VCC.n255 VSS 0.003222f
C290 VCC.n256 VSS 0.055238f
C291 VCC.n257 VSS 0.055238f
C292 VCC.n258 VSS 0.003222f
C293 VCC.n259 VSS 0.002593f
C294 VCC.n260 VSS 0.003222f
C295 VCC.n261 VSS 0.003222f
C296 VCC.n262 VSS 0.003222f
C297 VCC.n263 VSS 0.002593f
C298 VCC.n264 VSS 0.003222f
C299 VCC.n265 VSS 0.003222f
C300 VCC.n266 VSS 0.055238f
C301 VCC.n267 VSS 0.003222f
C302 VCC.n268 VSS 0.002593f
C303 VCC.n269 VSS 0.003222f
C304 VCC.n270 VSS 0.003222f
C305 VCC.n271 VSS 0.003222f
C306 VCC.n272 VSS 0.002593f
C307 VCC.n273 VSS 0.003222f
C308 VCC.n274 VSS 0.055238f
C309 VCC.n275 VSS 0.055238f
C310 VCC.n276 VSS 0.003222f
C311 VCC.n277 VSS 0.055238f
C312 VCC.n278 VSS 0.003222f
C313 VCC.n279 VSS 0.002593f
C314 VCC.n280 VSS 0.003222f
C315 VCC.n281 VSS 0.003222f
C316 VCC.n282 VSS 0.003222f
C317 VCC.n283 VSS 0.002593f
C318 VCC.n284 VSS 0.003222f
C319 VCC.n285 VSS 0.055238f
C320 VCC.n286 VSS 0.055238f
C321 VCC.t1 VSS 0.027619f
C322 VCC.n287 VSS 0.003222f
C323 VCC.n288 VSS 0.053581f
C324 VCC.n289 VSS 0.003222f
C325 VCC.n290 VSS 0.002593f
C326 VCC.n291 VSS 0.003222f
C327 VCC.n292 VSS 0.003222f
C328 VCC.n293 VSS 0.003222f
C329 VCC.n294 VSS 0.002593f
C330 VCC.n295 VSS 0.003222f
C331 VCC.n296 VSS 0.055238f
C332 VCC.n297 VSS 0.055238f
C333 VCC.n298 VSS 0.003222f
C334 VCC.n299 VSS 0.055238f
C335 VCC.n300 VSS 0.003222f
C336 VCC.n301 VSS 0.002593f
C337 VCC.n302 VSS 0.003222f
C338 VCC.n303 VSS 0.003222f
C339 VCC.n304 VSS 0.003222f
C340 VCC.n305 VSS 0.002593f
C341 VCC.n306 VSS 0.003222f
C342 VCC.n307 VSS 0.055238f
C343 VCC.n308 VSS 0.055238f
C344 VCC.n309 VSS 0.003222f
C345 VCC.n310 VSS 0.055238f
C346 VCC.n311 VSS 0.003222f
C347 VCC.n312 VSS 0.002593f
C348 VCC.n313 VSS 0.003222f
C349 VCC.n314 VSS 0.003222f
C350 VCC.n315 VSS 0.003222f
C351 VCC.n316 VSS 0.002593f
C352 VCC.n317 VSS 0.003222f
C353 VCC.n318 VSS 0.055238f
C354 VCC.n319 VSS 0.029276f
C355 VCC.t3 VSS 0.027619f
C356 VCC.n320 VSS 0.055238f
C357 VCC.n321 VSS 0.055238f
C358 VCC.n322 VSS 0.003222f
C359 VCC.n323 VSS 0.053581f
C360 VCC.n324 VSS 0.003222f
C361 VCC.n325 VSS 0.002593f
C362 VCC.n326 VSS 0.003222f
C363 VCC.n327 VSS 0.003222f
C364 VCC.n328 VSS 0.003222f
C365 VCC.n329 VSS 0.002593f
C366 VCC.n330 VSS 0.002152f
C367 VCC.n331 VSS 0.006483f
C368 VCC.n332 VSS 0.0065f
C369 VCC.n333 VSS 0.004238f
C370 VCC.n334 VSS 0.002191f
C371 VCC.n335 VSS 0.002191f
C372 VCC.n336 VSS 0.002191f
C373 VCC.n337 VSS 0.002191f
C374 VCC.n338 VSS 0.002191f
C375 VCC.n339 VSS 0.002191f
C376 VCC.n340 VSS 0.002191f
C377 VCC.n341 VSS 0.002191f
C378 VCC.n342 VSS 0.002191f
C379 VCC.n343 VSS 0.002191f
C380 VCC.n344 VSS 0.002191f
C381 VCC.n345 VSS 0.002191f
C382 VCC.n346 VSS 0.002191f
C383 VCC.n347 VSS 0.002191f
C384 VCC.n348 VSS 0.002191f
C385 VCC.n349 VSS 0.002191f
C386 VCC.n350 VSS 0.002191f
C387 VCC.n351 VSS 0.002191f
C388 VCC.n352 VSS 0.002191f
C389 VCC.n353 VSS 0.002191f
C390 VCC.n354 VSS 0.002191f
C391 VCC.n355 VSS 0.001434f
C392 VCC.n356 VSS 0.002191f
C393 VCC.n358 VSS 0.110752f
C394 VCC.n359 VSS 0.0065f
C395 VCC.n360 VSS 0.004238f
C396 VCC.n361 VSS 0.011386f
C397 VCC.n362 VSS 0.002152f
C398 VCC.n363 VSS 0.002593f
C399 VCC.n364 VSS 0.002593f
C400 VCC.n365 VSS 0.003222f
C401 VCC.n366 VSS 0.003222f
C402 VCC.n367 VSS 0.003222f
C403 VCC.n368 VSS 0.002593f
C404 VCC.n369 VSS 0.002593f
C405 VCC.n370 VSS 0.002593f
C406 VCC.n371 VSS 0.003222f
C407 VCC.n372 VSS 0.003222f
C408 VCC.n373 VSS 0.003222f
C409 VCC.n374 VSS 0.002593f
C410 VCC.n375 VSS 0.002593f
C411 VCC.n376 VSS 0.002593f
C412 VCC.n377 VSS 0.003222f
C413 VCC.n378 VSS 0.003222f
C414 VCC.n379 VSS 0.003222f
C415 VCC.n380 VSS 0.002593f
C416 VCC.n381 VSS 0.002593f
C417 VCC.n382 VSS 0.002593f
C418 VCC.n383 VSS 0.003222f
C419 VCC.n384 VSS 0.003222f
C420 VCC.n385 VSS 0.003222f
C421 VCC.n386 VSS 0.002593f
C422 VCC.n387 VSS 0.002593f
C423 VCC.n388 VSS 0.002593f
C424 VCC.n389 VSS 0.003222f
C425 VCC.n390 VSS 0.003222f
C426 VCC.n391 VSS 0.003222f
C427 VCC.n392 VSS 0.002593f
C428 VCC.n393 VSS 0.002593f
C429 VCC.n394 VSS 0.002593f
C430 VCC.n395 VSS 0.002947f
C431 VOUT.t0 VSS 0.245184f
C432 VOUT.t5 VSS 0.032057f
C433 VOUT.t1 VSS 0.032057f
C434 VOUT.n0 VSS 0.166284f
C435 VOUT.n1 VSS 0.750729f
C436 VOUT.n2 VSS 0.01934f
C437 VOUT.n3 VSS 0.013893f
C438 VOUT.n4 VSS 0.007465f
C439 VOUT.n5 VSS 0.017645f
C440 VOUT.n6 VSS 0.007904f
C441 VOUT.n7 VSS 0.053367f
C442 VOUT.t4 VSS 0.029286f
C443 VOUT.n8 VSS 0.013234f
C444 VOUT.n9 VSS 0.010385f
C445 VOUT.n10 VSS 0.007465f
C446 VOUT.n11 VSS 0.197724f
C447 VOUT.n12 VSS 0.013893f
C448 VOUT.n13 VSS 0.007465f
C449 VOUT.n14 VSS 0.007904f
C450 VOUT.n15 VSS 0.017645f
C451 VOUT.n16 VSS 0.037868f
C452 VOUT.n17 VSS 0.007904f
C453 VOUT.n18 VSS 0.007465f
C454 VOUT.n19 VSS 0.03401f
C455 VOUT.n20 VSS 0.03469f
C456 VOUT.t2 VSS 0.043255f
C457 VOUT.t3 VSS 0.043255f
C458 VOUT.n21 VSS 0.33896f
C459 VOUT.n22 VSS 0.571847f
C460 VIN.t1 VSS 0.225501f
C461 VIN.t0 VSS 0.032398f
C462 VIN.t5 VSS 0.032398f
C463 VIN.n0 VSS 0.144837f
C464 VIN.n1 VSS 0.973234f
C465 VIN.n2 VSS 0.019545f
C466 VIN.n3 VSS 0.01404f
C467 VIN.n4 VSS 0.007545f
C468 VIN.n5 VSS 0.017833f
C469 VIN.n6 VSS 0.007988f
C470 VIN.n7 VSS 0.053934f
C471 VIN.t3 VSS 0.029597f
C472 VIN.n8 VSS 0.013375f
C473 VIN.n9 VSS 0.010496f
C474 VIN.n10 VSS 0.007545f
C475 VIN.n11 VSS 0.199824f
C476 VIN.n12 VSS 0.01404f
C477 VIN.n13 VSS 0.007545f
C478 VIN.n14 VSS 0.007988f
C479 VIN.n15 VSS 0.017833f
C480 VIN.n16 VSS 0.03827f
C481 VIN.n17 VSS 0.007988f
C482 VIN.n18 VSS 0.007545f
C483 VIN.n19 VSS 0.034371f
C484 VIN.n20 VSS 0.026721f
C485 VIN.t4 VSS 0.043715f
C486 VIN.t2 VSS 0.043715f
C487 VIN.n21 VSS 0.312329f
C488 VIN.n22 VSS 0.343535f
.ends

