* NGSPICE file created from diff_pair_sample_1154.ext - technology: sky130A

.subckt diff_pair_sample_1154 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=1.83
X1 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=1.83
X2 VTAIL.t6 VN.t1 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=1.83
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=1.83
X4 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=1.83
X5 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=1.83
X6 VDD2.t3 VN.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=1.83
X7 VDD2.t0 VN.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=1.83
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=1.83
X9 VDD1.t0 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=1.83
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=1.83
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=1.83
R0 VN.n0 VN.t1 83.4755
R1 VN.n1 VN.t3 83.4755
R2 VN.n0 VN.t2 83.0418
R3 VN.n1 VN.t0 83.0418
R4 VN VN.n1 47.0894
R5 VN VN.n0 9.24472
R6 VDD2.n2 VDD2.n0 108.674
R7 VDD2.n2 VDD2.n1 76.3302
R8 VDD2.n1 VDD2.t2 5.60957
R9 VDD2.n1 VDD2.t0 5.60957
R10 VDD2.n0 VDD2.t1 5.60957
R11 VDD2.n0 VDD2.t3 5.60957
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t0 65.2605
R14 VTAIL.n4 VTAIL.t4 65.2605
R15 VTAIL.n3 VTAIL.t7 65.2605
R16 VTAIL.n7 VTAIL.t5 65.2605
R17 VTAIL.n0 VTAIL.t6 65.2605
R18 VTAIL.n1 VTAIL.t3 65.2605
R19 VTAIL.n2 VTAIL.t1 65.2605
R20 VTAIL.n6 VTAIL.t2 65.2605
R21 VTAIL.n7 VTAIL.n6 17.2721
R22 VTAIL.n3 VTAIL.n2 17.2721
R23 VTAIL.n4 VTAIL.n3 1.86257
R24 VTAIL.n6 VTAIL.n5 1.86257
R25 VTAIL.n2 VTAIL.n1 1.86257
R26 VTAIL VTAIL.n0 0.989724
R27 VTAIL VTAIL.n7 0.873345
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n442 B.n441 585
R31 B.n443 B.n442 585
R32 B.n160 B.n74 585
R33 B.n159 B.n158 585
R34 B.n157 B.n156 585
R35 B.n155 B.n154 585
R36 B.n153 B.n152 585
R37 B.n151 B.n150 585
R38 B.n149 B.n148 585
R39 B.n147 B.n146 585
R40 B.n145 B.n144 585
R41 B.n143 B.n142 585
R42 B.n141 B.n140 585
R43 B.n139 B.n138 585
R44 B.n137 B.n136 585
R45 B.n135 B.n134 585
R46 B.n133 B.n132 585
R47 B.n131 B.n130 585
R48 B.n129 B.n128 585
R49 B.n127 B.n126 585
R50 B.n125 B.n124 585
R51 B.n123 B.n122 585
R52 B.n121 B.n120 585
R53 B.n119 B.n118 585
R54 B.n117 B.n116 585
R55 B.n115 B.n114 585
R56 B.n113 B.n112 585
R57 B.n110 B.n109 585
R58 B.n108 B.n107 585
R59 B.n106 B.n105 585
R60 B.n104 B.n103 585
R61 B.n102 B.n101 585
R62 B.n100 B.n99 585
R63 B.n98 B.n97 585
R64 B.n96 B.n95 585
R65 B.n94 B.n93 585
R66 B.n92 B.n91 585
R67 B.n90 B.n89 585
R68 B.n88 B.n87 585
R69 B.n86 B.n85 585
R70 B.n84 B.n83 585
R71 B.n82 B.n81 585
R72 B.n53 B.n52 585
R73 B.n446 B.n445 585
R74 B.n440 B.n75 585
R75 B.n75 B.n50 585
R76 B.n439 B.n49 585
R77 B.n450 B.n49 585
R78 B.n438 B.n48 585
R79 B.n451 B.n48 585
R80 B.n437 B.n47 585
R81 B.n452 B.n47 585
R82 B.n436 B.n435 585
R83 B.n435 B.n43 585
R84 B.n434 B.n42 585
R85 B.n458 B.n42 585
R86 B.n433 B.n41 585
R87 B.n459 B.n41 585
R88 B.n432 B.n40 585
R89 B.n460 B.n40 585
R90 B.n431 B.n430 585
R91 B.n430 B.n36 585
R92 B.n429 B.n35 585
R93 B.n466 B.n35 585
R94 B.n428 B.n34 585
R95 B.n467 B.n34 585
R96 B.n427 B.n33 585
R97 B.n468 B.n33 585
R98 B.n426 B.n425 585
R99 B.n425 B.n29 585
R100 B.n424 B.n28 585
R101 B.n474 B.n28 585
R102 B.n423 B.n27 585
R103 B.n475 B.n27 585
R104 B.n422 B.n26 585
R105 B.n476 B.n26 585
R106 B.n421 B.n420 585
R107 B.n420 B.n22 585
R108 B.n419 B.n21 585
R109 B.n482 B.n21 585
R110 B.n418 B.n20 585
R111 B.n483 B.n20 585
R112 B.n417 B.n19 585
R113 B.n484 B.n19 585
R114 B.n416 B.n415 585
R115 B.n415 B.n15 585
R116 B.n414 B.n14 585
R117 B.n490 B.n14 585
R118 B.n413 B.n13 585
R119 B.n491 B.n13 585
R120 B.n412 B.n12 585
R121 B.n492 B.n12 585
R122 B.n411 B.n410 585
R123 B.n410 B.n8 585
R124 B.n409 B.n7 585
R125 B.n498 B.n7 585
R126 B.n408 B.n6 585
R127 B.n499 B.n6 585
R128 B.n407 B.n5 585
R129 B.n500 B.n5 585
R130 B.n406 B.n405 585
R131 B.n405 B.n4 585
R132 B.n404 B.n161 585
R133 B.n404 B.n403 585
R134 B.n394 B.n162 585
R135 B.n163 B.n162 585
R136 B.n396 B.n395 585
R137 B.n397 B.n396 585
R138 B.n393 B.n167 585
R139 B.n171 B.n167 585
R140 B.n392 B.n391 585
R141 B.n391 B.n390 585
R142 B.n169 B.n168 585
R143 B.n170 B.n169 585
R144 B.n383 B.n382 585
R145 B.n384 B.n383 585
R146 B.n381 B.n176 585
R147 B.n176 B.n175 585
R148 B.n380 B.n379 585
R149 B.n379 B.n378 585
R150 B.n178 B.n177 585
R151 B.n179 B.n178 585
R152 B.n371 B.n370 585
R153 B.n372 B.n371 585
R154 B.n369 B.n184 585
R155 B.n184 B.n183 585
R156 B.n368 B.n367 585
R157 B.n367 B.n366 585
R158 B.n186 B.n185 585
R159 B.n187 B.n186 585
R160 B.n359 B.n358 585
R161 B.n360 B.n359 585
R162 B.n357 B.n192 585
R163 B.n192 B.n191 585
R164 B.n356 B.n355 585
R165 B.n355 B.n354 585
R166 B.n194 B.n193 585
R167 B.n195 B.n194 585
R168 B.n347 B.n346 585
R169 B.n348 B.n347 585
R170 B.n345 B.n199 585
R171 B.n203 B.n199 585
R172 B.n344 B.n343 585
R173 B.n343 B.n342 585
R174 B.n201 B.n200 585
R175 B.n202 B.n201 585
R176 B.n335 B.n334 585
R177 B.n336 B.n335 585
R178 B.n333 B.n208 585
R179 B.n208 B.n207 585
R180 B.n332 B.n331 585
R181 B.n331 B.n330 585
R182 B.n210 B.n209 585
R183 B.n211 B.n210 585
R184 B.n326 B.n325 585
R185 B.n214 B.n213 585
R186 B.n322 B.n321 585
R187 B.n323 B.n322 585
R188 B.n320 B.n235 585
R189 B.n319 B.n318 585
R190 B.n317 B.n316 585
R191 B.n315 B.n314 585
R192 B.n313 B.n312 585
R193 B.n311 B.n310 585
R194 B.n309 B.n308 585
R195 B.n307 B.n306 585
R196 B.n305 B.n304 585
R197 B.n303 B.n302 585
R198 B.n301 B.n300 585
R199 B.n299 B.n298 585
R200 B.n297 B.n296 585
R201 B.n295 B.n294 585
R202 B.n293 B.n292 585
R203 B.n291 B.n290 585
R204 B.n289 B.n288 585
R205 B.n287 B.n286 585
R206 B.n285 B.n284 585
R207 B.n283 B.n282 585
R208 B.n281 B.n280 585
R209 B.n279 B.n278 585
R210 B.n277 B.n276 585
R211 B.n274 B.n273 585
R212 B.n272 B.n271 585
R213 B.n270 B.n269 585
R214 B.n268 B.n267 585
R215 B.n266 B.n265 585
R216 B.n264 B.n263 585
R217 B.n262 B.n261 585
R218 B.n260 B.n259 585
R219 B.n258 B.n257 585
R220 B.n256 B.n255 585
R221 B.n254 B.n253 585
R222 B.n252 B.n251 585
R223 B.n250 B.n249 585
R224 B.n248 B.n247 585
R225 B.n246 B.n245 585
R226 B.n244 B.n243 585
R227 B.n242 B.n241 585
R228 B.n327 B.n212 585
R229 B.n212 B.n211 585
R230 B.n329 B.n328 585
R231 B.n330 B.n329 585
R232 B.n206 B.n205 585
R233 B.n207 B.n206 585
R234 B.n338 B.n337 585
R235 B.n337 B.n336 585
R236 B.n339 B.n204 585
R237 B.n204 B.n202 585
R238 B.n341 B.n340 585
R239 B.n342 B.n341 585
R240 B.n198 B.n197 585
R241 B.n203 B.n198 585
R242 B.n350 B.n349 585
R243 B.n349 B.n348 585
R244 B.n351 B.n196 585
R245 B.n196 B.n195 585
R246 B.n353 B.n352 585
R247 B.n354 B.n353 585
R248 B.n190 B.n189 585
R249 B.n191 B.n190 585
R250 B.n362 B.n361 585
R251 B.n361 B.n360 585
R252 B.n363 B.n188 585
R253 B.n188 B.n187 585
R254 B.n365 B.n364 585
R255 B.n366 B.n365 585
R256 B.n182 B.n181 585
R257 B.n183 B.n182 585
R258 B.n374 B.n373 585
R259 B.n373 B.n372 585
R260 B.n375 B.n180 585
R261 B.n180 B.n179 585
R262 B.n377 B.n376 585
R263 B.n378 B.n377 585
R264 B.n174 B.n173 585
R265 B.n175 B.n174 585
R266 B.n386 B.n385 585
R267 B.n385 B.n384 585
R268 B.n387 B.n172 585
R269 B.n172 B.n170 585
R270 B.n389 B.n388 585
R271 B.n390 B.n389 585
R272 B.n166 B.n165 585
R273 B.n171 B.n166 585
R274 B.n399 B.n398 585
R275 B.n398 B.n397 585
R276 B.n400 B.n164 585
R277 B.n164 B.n163 585
R278 B.n402 B.n401 585
R279 B.n403 B.n402 585
R280 B.n2 B.n0 585
R281 B.n4 B.n2 585
R282 B.n3 B.n1 585
R283 B.n499 B.n3 585
R284 B.n497 B.n496 585
R285 B.n498 B.n497 585
R286 B.n495 B.n9 585
R287 B.n9 B.n8 585
R288 B.n494 B.n493 585
R289 B.n493 B.n492 585
R290 B.n11 B.n10 585
R291 B.n491 B.n11 585
R292 B.n489 B.n488 585
R293 B.n490 B.n489 585
R294 B.n487 B.n16 585
R295 B.n16 B.n15 585
R296 B.n486 B.n485 585
R297 B.n485 B.n484 585
R298 B.n18 B.n17 585
R299 B.n483 B.n18 585
R300 B.n481 B.n480 585
R301 B.n482 B.n481 585
R302 B.n479 B.n23 585
R303 B.n23 B.n22 585
R304 B.n478 B.n477 585
R305 B.n477 B.n476 585
R306 B.n25 B.n24 585
R307 B.n475 B.n25 585
R308 B.n473 B.n472 585
R309 B.n474 B.n473 585
R310 B.n471 B.n30 585
R311 B.n30 B.n29 585
R312 B.n470 B.n469 585
R313 B.n469 B.n468 585
R314 B.n32 B.n31 585
R315 B.n467 B.n32 585
R316 B.n465 B.n464 585
R317 B.n466 B.n465 585
R318 B.n463 B.n37 585
R319 B.n37 B.n36 585
R320 B.n462 B.n461 585
R321 B.n461 B.n460 585
R322 B.n39 B.n38 585
R323 B.n459 B.n39 585
R324 B.n457 B.n456 585
R325 B.n458 B.n457 585
R326 B.n455 B.n44 585
R327 B.n44 B.n43 585
R328 B.n454 B.n453 585
R329 B.n453 B.n452 585
R330 B.n46 B.n45 585
R331 B.n451 B.n46 585
R332 B.n449 B.n448 585
R333 B.n450 B.n449 585
R334 B.n447 B.n51 585
R335 B.n51 B.n50 585
R336 B.n502 B.n501 585
R337 B.n501 B.n500 585
R338 B.n325 B.n212 526.135
R339 B.n445 B.n51 526.135
R340 B.n241 B.n210 526.135
R341 B.n442 B.n75 526.135
R342 B.n443 B.n73 256.663
R343 B.n443 B.n72 256.663
R344 B.n443 B.n71 256.663
R345 B.n443 B.n70 256.663
R346 B.n443 B.n69 256.663
R347 B.n443 B.n68 256.663
R348 B.n443 B.n67 256.663
R349 B.n443 B.n66 256.663
R350 B.n443 B.n65 256.663
R351 B.n443 B.n64 256.663
R352 B.n443 B.n63 256.663
R353 B.n443 B.n62 256.663
R354 B.n443 B.n61 256.663
R355 B.n443 B.n60 256.663
R356 B.n443 B.n59 256.663
R357 B.n443 B.n58 256.663
R358 B.n443 B.n57 256.663
R359 B.n443 B.n56 256.663
R360 B.n443 B.n55 256.663
R361 B.n443 B.n54 256.663
R362 B.n444 B.n443 256.663
R363 B.n324 B.n323 256.663
R364 B.n323 B.n215 256.663
R365 B.n323 B.n216 256.663
R366 B.n323 B.n217 256.663
R367 B.n323 B.n218 256.663
R368 B.n323 B.n219 256.663
R369 B.n323 B.n220 256.663
R370 B.n323 B.n221 256.663
R371 B.n323 B.n222 256.663
R372 B.n323 B.n223 256.663
R373 B.n323 B.n224 256.663
R374 B.n323 B.n225 256.663
R375 B.n323 B.n226 256.663
R376 B.n323 B.n227 256.663
R377 B.n323 B.n228 256.663
R378 B.n323 B.n229 256.663
R379 B.n323 B.n230 256.663
R380 B.n323 B.n231 256.663
R381 B.n323 B.n232 256.663
R382 B.n323 B.n233 256.663
R383 B.n323 B.n234 256.663
R384 B.n239 B.t4 252.976
R385 B.n236 B.t15 252.976
R386 B.n79 B.t12 252.976
R387 B.n76 B.t8 252.976
R388 B.n323 B.n211 168.655
R389 B.n443 B.n50 168.655
R390 B.n329 B.n212 163.367
R391 B.n329 B.n206 163.367
R392 B.n337 B.n206 163.367
R393 B.n337 B.n204 163.367
R394 B.n341 B.n204 163.367
R395 B.n341 B.n198 163.367
R396 B.n349 B.n198 163.367
R397 B.n349 B.n196 163.367
R398 B.n353 B.n196 163.367
R399 B.n353 B.n190 163.367
R400 B.n361 B.n190 163.367
R401 B.n361 B.n188 163.367
R402 B.n365 B.n188 163.367
R403 B.n365 B.n182 163.367
R404 B.n373 B.n182 163.367
R405 B.n373 B.n180 163.367
R406 B.n377 B.n180 163.367
R407 B.n377 B.n174 163.367
R408 B.n385 B.n174 163.367
R409 B.n385 B.n172 163.367
R410 B.n389 B.n172 163.367
R411 B.n389 B.n166 163.367
R412 B.n398 B.n166 163.367
R413 B.n398 B.n164 163.367
R414 B.n402 B.n164 163.367
R415 B.n402 B.n2 163.367
R416 B.n501 B.n2 163.367
R417 B.n501 B.n3 163.367
R418 B.n497 B.n3 163.367
R419 B.n497 B.n9 163.367
R420 B.n493 B.n9 163.367
R421 B.n493 B.n11 163.367
R422 B.n489 B.n11 163.367
R423 B.n489 B.n16 163.367
R424 B.n485 B.n16 163.367
R425 B.n485 B.n18 163.367
R426 B.n481 B.n18 163.367
R427 B.n481 B.n23 163.367
R428 B.n477 B.n23 163.367
R429 B.n477 B.n25 163.367
R430 B.n473 B.n25 163.367
R431 B.n473 B.n30 163.367
R432 B.n469 B.n30 163.367
R433 B.n469 B.n32 163.367
R434 B.n465 B.n32 163.367
R435 B.n465 B.n37 163.367
R436 B.n461 B.n37 163.367
R437 B.n461 B.n39 163.367
R438 B.n457 B.n39 163.367
R439 B.n457 B.n44 163.367
R440 B.n453 B.n44 163.367
R441 B.n453 B.n46 163.367
R442 B.n449 B.n46 163.367
R443 B.n449 B.n51 163.367
R444 B.n322 B.n214 163.367
R445 B.n322 B.n235 163.367
R446 B.n318 B.n317 163.367
R447 B.n314 B.n313 163.367
R448 B.n310 B.n309 163.367
R449 B.n306 B.n305 163.367
R450 B.n302 B.n301 163.367
R451 B.n298 B.n297 163.367
R452 B.n294 B.n293 163.367
R453 B.n290 B.n289 163.367
R454 B.n286 B.n285 163.367
R455 B.n282 B.n281 163.367
R456 B.n278 B.n277 163.367
R457 B.n273 B.n272 163.367
R458 B.n269 B.n268 163.367
R459 B.n265 B.n264 163.367
R460 B.n261 B.n260 163.367
R461 B.n257 B.n256 163.367
R462 B.n253 B.n252 163.367
R463 B.n249 B.n248 163.367
R464 B.n245 B.n244 163.367
R465 B.n331 B.n210 163.367
R466 B.n331 B.n208 163.367
R467 B.n335 B.n208 163.367
R468 B.n335 B.n201 163.367
R469 B.n343 B.n201 163.367
R470 B.n343 B.n199 163.367
R471 B.n347 B.n199 163.367
R472 B.n347 B.n194 163.367
R473 B.n355 B.n194 163.367
R474 B.n355 B.n192 163.367
R475 B.n359 B.n192 163.367
R476 B.n359 B.n186 163.367
R477 B.n367 B.n186 163.367
R478 B.n367 B.n184 163.367
R479 B.n371 B.n184 163.367
R480 B.n371 B.n178 163.367
R481 B.n379 B.n178 163.367
R482 B.n379 B.n176 163.367
R483 B.n383 B.n176 163.367
R484 B.n383 B.n169 163.367
R485 B.n391 B.n169 163.367
R486 B.n391 B.n167 163.367
R487 B.n396 B.n167 163.367
R488 B.n396 B.n162 163.367
R489 B.n404 B.n162 163.367
R490 B.n405 B.n404 163.367
R491 B.n405 B.n5 163.367
R492 B.n6 B.n5 163.367
R493 B.n7 B.n6 163.367
R494 B.n410 B.n7 163.367
R495 B.n410 B.n12 163.367
R496 B.n13 B.n12 163.367
R497 B.n14 B.n13 163.367
R498 B.n415 B.n14 163.367
R499 B.n415 B.n19 163.367
R500 B.n20 B.n19 163.367
R501 B.n21 B.n20 163.367
R502 B.n420 B.n21 163.367
R503 B.n420 B.n26 163.367
R504 B.n27 B.n26 163.367
R505 B.n28 B.n27 163.367
R506 B.n425 B.n28 163.367
R507 B.n425 B.n33 163.367
R508 B.n34 B.n33 163.367
R509 B.n35 B.n34 163.367
R510 B.n430 B.n35 163.367
R511 B.n430 B.n40 163.367
R512 B.n41 B.n40 163.367
R513 B.n42 B.n41 163.367
R514 B.n435 B.n42 163.367
R515 B.n435 B.n47 163.367
R516 B.n48 B.n47 163.367
R517 B.n49 B.n48 163.367
R518 B.n75 B.n49 163.367
R519 B.n81 B.n53 163.367
R520 B.n85 B.n84 163.367
R521 B.n89 B.n88 163.367
R522 B.n93 B.n92 163.367
R523 B.n97 B.n96 163.367
R524 B.n101 B.n100 163.367
R525 B.n105 B.n104 163.367
R526 B.n109 B.n108 163.367
R527 B.n114 B.n113 163.367
R528 B.n118 B.n117 163.367
R529 B.n122 B.n121 163.367
R530 B.n126 B.n125 163.367
R531 B.n130 B.n129 163.367
R532 B.n134 B.n133 163.367
R533 B.n138 B.n137 163.367
R534 B.n142 B.n141 163.367
R535 B.n146 B.n145 163.367
R536 B.n150 B.n149 163.367
R537 B.n154 B.n153 163.367
R538 B.n158 B.n157 163.367
R539 B.n442 B.n74 163.367
R540 B.n239 B.t7 116.983
R541 B.n76 B.t10 116.983
R542 B.n236 B.t17 116.98
R543 B.n79 B.t13 116.98
R544 B.n330 B.n211 84.9522
R545 B.n330 B.n207 84.9522
R546 B.n336 B.n207 84.9522
R547 B.n336 B.n202 84.9522
R548 B.n342 B.n202 84.9522
R549 B.n342 B.n203 84.9522
R550 B.n348 B.n195 84.9522
R551 B.n354 B.n195 84.9522
R552 B.n354 B.n191 84.9522
R553 B.n360 B.n191 84.9522
R554 B.n360 B.n187 84.9522
R555 B.n366 B.n187 84.9522
R556 B.n366 B.n183 84.9522
R557 B.n372 B.n183 84.9522
R558 B.n378 B.n179 84.9522
R559 B.n378 B.n175 84.9522
R560 B.n384 B.n175 84.9522
R561 B.n384 B.n170 84.9522
R562 B.n390 B.n170 84.9522
R563 B.n390 B.n171 84.9522
R564 B.n397 B.n163 84.9522
R565 B.n403 B.n163 84.9522
R566 B.n403 B.n4 84.9522
R567 B.n500 B.n4 84.9522
R568 B.n500 B.n499 84.9522
R569 B.n499 B.n498 84.9522
R570 B.n498 B.n8 84.9522
R571 B.n492 B.n8 84.9522
R572 B.n491 B.n490 84.9522
R573 B.n490 B.n15 84.9522
R574 B.n484 B.n15 84.9522
R575 B.n484 B.n483 84.9522
R576 B.n483 B.n482 84.9522
R577 B.n482 B.n22 84.9522
R578 B.n476 B.n475 84.9522
R579 B.n475 B.n474 84.9522
R580 B.n474 B.n29 84.9522
R581 B.n468 B.n29 84.9522
R582 B.n468 B.n467 84.9522
R583 B.n467 B.n466 84.9522
R584 B.n466 B.n36 84.9522
R585 B.n460 B.n36 84.9522
R586 B.n459 B.n458 84.9522
R587 B.n458 B.n43 84.9522
R588 B.n452 B.n43 84.9522
R589 B.n452 B.n451 84.9522
R590 B.n451 B.n450 84.9522
R591 B.n450 B.n50 84.9522
R592 B.n240 B.t6 75.0918
R593 B.n77 B.t11 75.0918
R594 B.n237 B.t16 75.0889
R595 B.n80 B.t14 75.0889
R596 B.n372 B.t1 73.7086
R597 B.n476 B.t2 73.7086
R598 B.n325 B.n324 71.676
R599 B.n235 B.n215 71.676
R600 B.n317 B.n216 71.676
R601 B.n313 B.n217 71.676
R602 B.n309 B.n218 71.676
R603 B.n305 B.n219 71.676
R604 B.n301 B.n220 71.676
R605 B.n297 B.n221 71.676
R606 B.n293 B.n222 71.676
R607 B.n289 B.n223 71.676
R608 B.n285 B.n224 71.676
R609 B.n281 B.n225 71.676
R610 B.n277 B.n226 71.676
R611 B.n272 B.n227 71.676
R612 B.n268 B.n228 71.676
R613 B.n264 B.n229 71.676
R614 B.n260 B.n230 71.676
R615 B.n256 B.n231 71.676
R616 B.n252 B.n232 71.676
R617 B.n248 B.n233 71.676
R618 B.n244 B.n234 71.676
R619 B.n445 B.n444 71.676
R620 B.n81 B.n54 71.676
R621 B.n85 B.n55 71.676
R622 B.n89 B.n56 71.676
R623 B.n93 B.n57 71.676
R624 B.n97 B.n58 71.676
R625 B.n101 B.n59 71.676
R626 B.n105 B.n60 71.676
R627 B.n109 B.n61 71.676
R628 B.n114 B.n62 71.676
R629 B.n118 B.n63 71.676
R630 B.n122 B.n64 71.676
R631 B.n126 B.n65 71.676
R632 B.n130 B.n66 71.676
R633 B.n134 B.n67 71.676
R634 B.n138 B.n68 71.676
R635 B.n142 B.n69 71.676
R636 B.n146 B.n70 71.676
R637 B.n150 B.n71 71.676
R638 B.n154 B.n72 71.676
R639 B.n158 B.n73 71.676
R640 B.n74 B.n73 71.676
R641 B.n157 B.n72 71.676
R642 B.n153 B.n71 71.676
R643 B.n149 B.n70 71.676
R644 B.n145 B.n69 71.676
R645 B.n141 B.n68 71.676
R646 B.n137 B.n67 71.676
R647 B.n133 B.n66 71.676
R648 B.n129 B.n65 71.676
R649 B.n125 B.n64 71.676
R650 B.n121 B.n63 71.676
R651 B.n117 B.n62 71.676
R652 B.n113 B.n61 71.676
R653 B.n108 B.n60 71.676
R654 B.n104 B.n59 71.676
R655 B.n100 B.n58 71.676
R656 B.n96 B.n57 71.676
R657 B.n92 B.n56 71.676
R658 B.n88 B.n55 71.676
R659 B.n84 B.n54 71.676
R660 B.n444 B.n53 71.676
R661 B.n324 B.n214 71.676
R662 B.n318 B.n215 71.676
R663 B.n314 B.n216 71.676
R664 B.n310 B.n217 71.676
R665 B.n306 B.n218 71.676
R666 B.n302 B.n219 71.676
R667 B.n298 B.n220 71.676
R668 B.n294 B.n221 71.676
R669 B.n290 B.n222 71.676
R670 B.n286 B.n223 71.676
R671 B.n282 B.n224 71.676
R672 B.n278 B.n225 71.676
R673 B.n273 B.n226 71.676
R674 B.n269 B.n227 71.676
R675 B.n265 B.n228 71.676
R676 B.n261 B.n229 71.676
R677 B.n257 B.n230 71.676
R678 B.n253 B.n231 71.676
R679 B.n249 B.n232 71.676
R680 B.n245 B.n233 71.676
R681 B.n241 B.n234 71.676
R682 B.n397 B.t3 66.2129
R683 B.n492 B.t0 66.2129
R684 B.n275 B.n240 59.5399
R685 B.n238 B.n237 59.5399
R686 B.n111 B.n80 59.5399
R687 B.n78 B.n77 59.5399
R688 B.n348 B.t5 58.7171
R689 B.n460 B.t9 58.7171
R690 B.n240 B.n239 41.8914
R691 B.n237 B.n236 41.8914
R692 B.n80 B.n79 41.8914
R693 B.n77 B.n76 41.8914
R694 B.n447 B.n446 34.1859
R695 B.n441 B.n440 34.1859
R696 B.n242 B.n209 34.1859
R697 B.n327 B.n326 34.1859
R698 B.n203 B.t5 26.2356
R699 B.t9 B.n459 26.2356
R700 B.n171 B.t3 18.7399
R701 B.t0 B.n491 18.7399
R702 B B.n502 18.0485
R703 B.t1 B.n179 11.2441
R704 B.t2 B.n22 11.2441
R705 B.n446 B.n52 10.6151
R706 B.n82 B.n52 10.6151
R707 B.n83 B.n82 10.6151
R708 B.n86 B.n83 10.6151
R709 B.n87 B.n86 10.6151
R710 B.n90 B.n87 10.6151
R711 B.n91 B.n90 10.6151
R712 B.n94 B.n91 10.6151
R713 B.n95 B.n94 10.6151
R714 B.n98 B.n95 10.6151
R715 B.n99 B.n98 10.6151
R716 B.n102 B.n99 10.6151
R717 B.n103 B.n102 10.6151
R718 B.n106 B.n103 10.6151
R719 B.n107 B.n106 10.6151
R720 B.n110 B.n107 10.6151
R721 B.n115 B.n112 10.6151
R722 B.n116 B.n115 10.6151
R723 B.n119 B.n116 10.6151
R724 B.n120 B.n119 10.6151
R725 B.n123 B.n120 10.6151
R726 B.n124 B.n123 10.6151
R727 B.n127 B.n124 10.6151
R728 B.n128 B.n127 10.6151
R729 B.n132 B.n131 10.6151
R730 B.n135 B.n132 10.6151
R731 B.n136 B.n135 10.6151
R732 B.n139 B.n136 10.6151
R733 B.n140 B.n139 10.6151
R734 B.n143 B.n140 10.6151
R735 B.n144 B.n143 10.6151
R736 B.n147 B.n144 10.6151
R737 B.n148 B.n147 10.6151
R738 B.n151 B.n148 10.6151
R739 B.n152 B.n151 10.6151
R740 B.n155 B.n152 10.6151
R741 B.n156 B.n155 10.6151
R742 B.n159 B.n156 10.6151
R743 B.n160 B.n159 10.6151
R744 B.n441 B.n160 10.6151
R745 B.n332 B.n209 10.6151
R746 B.n333 B.n332 10.6151
R747 B.n334 B.n333 10.6151
R748 B.n334 B.n200 10.6151
R749 B.n344 B.n200 10.6151
R750 B.n345 B.n344 10.6151
R751 B.n346 B.n345 10.6151
R752 B.n346 B.n193 10.6151
R753 B.n356 B.n193 10.6151
R754 B.n357 B.n356 10.6151
R755 B.n358 B.n357 10.6151
R756 B.n358 B.n185 10.6151
R757 B.n368 B.n185 10.6151
R758 B.n369 B.n368 10.6151
R759 B.n370 B.n369 10.6151
R760 B.n370 B.n177 10.6151
R761 B.n380 B.n177 10.6151
R762 B.n381 B.n380 10.6151
R763 B.n382 B.n381 10.6151
R764 B.n382 B.n168 10.6151
R765 B.n392 B.n168 10.6151
R766 B.n393 B.n392 10.6151
R767 B.n395 B.n393 10.6151
R768 B.n395 B.n394 10.6151
R769 B.n394 B.n161 10.6151
R770 B.n406 B.n161 10.6151
R771 B.n407 B.n406 10.6151
R772 B.n408 B.n407 10.6151
R773 B.n409 B.n408 10.6151
R774 B.n411 B.n409 10.6151
R775 B.n412 B.n411 10.6151
R776 B.n413 B.n412 10.6151
R777 B.n414 B.n413 10.6151
R778 B.n416 B.n414 10.6151
R779 B.n417 B.n416 10.6151
R780 B.n418 B.n417 10.6151
R781 B.n419 B.n418 10.6151
R782 B.n421 B.n419 10.6151
R783 B.n422 B.n421 10.6151
R784 B.n423 B.n422 10.6151
R785 B.n424 B.n423 10.6151
R786 B.n426 B.n424 10.6151
R787 B.n427 B.n426 10.6151
R788 B.n428 B.n427 10.6151
R789 B.n429 B.n428 10.6151
R790 B.n431 B.n429 10.6151
R791 B.n432 B.n431 10.6151
R792 B.n433 B.n432 10.6151
R793 B.n434 B.n433 10.6151
R794 B.n436 B.n434 10.6151
R795 B.n437 B.n436 10.6151
R796 B.n438 B.n437 10.6151
R797 B.n439 B.n438 10.6151
R798 B.n440 B.n439 10.6151
R799 B.n326 B.n213 10.6151
R800 B.n321 B.n213 10.6151
R801 B.n321 B.n320 10.6151
R802 B.n320 B.n319 10.6151
R803 B.n319 B.n316 10.6151
R804 B.n316 B.n315 10.6151
R805 B.n315 B.n312 10.6151
R806 B.n312 B.n311 10.6151
R807 B.n311 B.n308 10.6151
R808 B.n308 B.n307 10.6151
R809 B.n307 B.n304 10.6151
R810 B.n304 B.n303 10.6151
R811 B.n303 B.n300 10.6151
R812 B.n300 B.n299 10.6151
R813 B.n299 B.n296 10.6151
R814 B.n296 B.n295 10.6151
R815 B.n292 B.n291 10.6151
R816 B.n291 B.n288 10.6151
R817 B.n288 B.n287 10.6151
R818 B.n287 B.n284 10.6151
R819 B.n284 B.n283 10.6151
R820 B.n283 B.n280 10.6151
R821 B.n280 B.n279 10.6151
R822 B.n279 B.n276 10.6151
R823 B.n274 B.n271 10.6151
R824 B.n271 B.n270 10.6151
R825 B.n270 B.n267 10.6151
R826 B.n267 B.n266 10.6151
R827 B.n266 B.n263 10.6151
R828 B.n263 B.n262 10.6151
R829 B.n262 B.n259 10.6151
R830 B.n259 B.n258 10.6151
R831 B.n258 B.n255 10.6151
R832 B.n255 B.n254 10.6151
R833 B.n254 B.n251 10.6151
R834 B.n251 B.n250 10.6151
R835 B.n250 B.n247 10.6151
R836 B.n247 B.n246 10.6151
R837 B.n246 B.n243 10.6151
R838 B.n243 B.n242 10.6151
R839 B.n328 B.n327 10.6151
R840 B.n328 B.n205 10.6151
R841 B.n338 B.n205 10.6151
R842 B.n339 B.n338 10.6151
R843 B.n340 B.n339 10.6151
R844 B.n340 B.n197 10.6151
R845 B.n350 B.n197 10.6151
R846 B.n351 B.n350 10.6151
R847 B.n352 B.n351 10.6151
R848 B.n352 B.n189 10.6151
R849 B.n362 B.n189 10.6151
R850 B.n363 B.n362 10.6151
R851 B.n364 B.n363 10.6151
R852 B.n364 B.n181 10.6151
R853 B.n374 B.n181 10.6151
R854 B.n375 B.n374 10.6151
R855 B.n376 B.n375 10.6151
R856 B.n376 B.n173 10.6151
R857 B.n386 B.n173 10.6151
R858 B.n387 B.n386 10.6151
R859 B.n388 B.n387 10.6151
R860 B.n388 B.n165 10.6151
R861 B.n399 B.n165 10.6151
R862 B.n400 B.n399 10.6151
R863 B.n401 B.n400 10.6151
R864 B.n401 B.n0 10.6151
R865 B.n496 B.n1 10.6151
R866 B.n496 B.n495 10.6151
R867 B.n495 B.n494 10.6151
R868 B.n494 B.n10 10.6151
R869 B.n488 B.n10 10.6151
R870 B.n488 B.n487 10.6151
R871 B.n487 B.n486 10.6151
R872 B.n486 B.n17 10.6151
R873 B.n480 B.n17 10.6151
R874 B.n480 B.n479 10.6151
R875 B.n479 B.n478 10.6151
R876 B.n478 B.n24 10.6151
R877 B.n472 B.n24 10.6151
R878 B.n472 B.n471 10.6151
R879 B.n471 B.n470 10.6151
R880 B.n470 B.n31 10.6151
R881 B.n464 B.n31 10.6151
R882 B.n464 B.n463 10.6151
R883 B.n463 B.n462 10.6151
R884 B.n462 B.n38 10.6151
R885 B.n456 B.n38 10.6151
R886 B.n456 B.n455 10.6151
R887 B.n455 B.n454 10.6151
R888 B.n454 B.n45 10.6151
R889 B.n448 B.n45 10.6151
R890 B.n448 B.n447 10.6151
R891 B.n112 B.n111 6.5566
R892 B.n128 B.n78 6.5566
R893 B.n292 B.n238 6.5566
R894 B.n276 B.n275 6.5566
R895 B.n111 B.n110 4.05904
R896 B.n131 B.n78 4.05904
R897 B.n295 B.n238 4.05904
R898 B.n275 B.n274 4.05904
R899 B.n502 B.n0 2.81026
R900 B.n502 B.n1 2.81026
R901 VP.n5 VP.n4 181.852
R902 VP.n14 VP.n13 181.852
R903 VP.n12 VP.n0 161.3
R904 VP.n11 VP.n10 161.3
R905 VP.n9 VP.n1 161.3
R906 VP.n8 VP.n7 161.3
R907 VP.n6 VP.n2 161.3
R908 VP.n3 VP.t1 83.4755
R909 VP.n3 VP.t3 83.0418
R910 VP.n4 VP.n3 46.7087
R911 VP.n5 VP.t2 46.4885
R912 VP.n13 VP.t0 46.4885
R913 VP.n7 VP.n1 40.4934
R914 VP.n11 VP.n1 40.4934
R915 VP.n7 VP.n6 24.4675
R916 VP.n12 VP.n11 24.4675
R917 VP.n6 VP.n5 3.91522
R918 VP.n13 VP.n12 3.91522
R919 VP.n4 VP.n2 0.189894
R920 VP.n8 VP.n2 0.189894
R921 VP.n9 VP.n8 0.189894
R922 VP.n10 VP.n9 0.189894
R923 VP.n10 VP.n0 0.189894
R924 VP.n14 VP.n0 0.189894
R925 VP VP.n14 0.0516364
R926 VDD1 VDD1.n1 109.2
R927 VDD1 VDD1.n0 76.3884
R928 VDD1.n0 VDD1.t2 5.60957
R929 VDD1.n0 VDD1.t0 5.60957
R930 VDD1.n1 VDD1.t1 5.60957
R931 VDD1.n1 VDD1.t3 5.60957
C0 VTAIL VN 1.79257f
C1 VTAIL VP 1.80668f
C2 VTAIL VDD2 3.12772f
C3 VDD1 VTAIL 3.07868f
C4 VP VN 4.07204f
C5 VDD2 VN 1.52217f
C6 VDD1 VN 0.152675f
C7 VP VDD2 0.350142f
C8 VDD1 VDD2 0.839251f
C9 VDD1 VP 1.7186f
C10 VDD2 B 2.607548f
C11 VDD1 B 4.63037f
C12 VTAIL B 4.326764f
C13 VN B 7.70496f
C14 VP B 6.548549f
C15 VDD1.t2 B 0.05019f
C16 VDD1.t0 B 0.05019f
C17 VDD1.n0 B 0.385861f
C18 VDD1.t1 B 0.05019f
C19 VDD1.t3 B 0.05019f
C20 VDD1.n1 B 0.610334f
C21 VP.n0 B 0.020581f
C22 VP.t0 B 0.337406f
C23 VP.n1 B 0.016638f
C24 VP.n2 B 0.020581f
C25 VP.t2 B 0.337406f
C26 VP.t1 B 0.445902f
C27 VP.t3 B 0.444661f
C28 VP.n3 B 0.985057f
C29 VP.n4 B 0.88857f
C30 VP.n5 B 0.19093f
C31 VP.n6 B 0.02245f
C32 VP.n7 B 0.040904f
C33 VP.n8 B 0.020581f
C34 VP.n9 B 0.020581f
C35 VP.n10 B 0.020581f
C36 VP.n11 B 0.040904f
C37 VP.n12 B 0.02245f
C38 VP.n13 B 0.19093f
C39 VP.n14 B 0.022039f
C40 VTAIL.t6 B 0.339534f
C41 VTAIL.n0 B 0.206869f
C42 VTAIL.t3 B 0.339534f
C43 VTAIL.n1 B 0.245252f
C44 VTAIL.t1 B 0.339534f
C45 VTAIL.n2 B 0.62568f
C46 VTAIL.t7 B 0.339536f
C47 VTAIL.n3 B 0.625678f
C48 VTAIL.t4 B 0.339536f
C49 VTAIL.n4 B 0.24525f
C50 VTAIL.t0 B 0.339536f
C51 VTAIL.n5 B 0.24525f
C52 VTAIL.t2 B 0.339534f
C53 VTAIL.n6 B 0.62568f
C54 VTAIL.t5 B 0.339534f
C55 VTAIL.n7 B 0.582179f
C56 VDD2.t1 B 0.05129f
C57 VDD2.t3 B 0.05129f
C58 VDD2.n0 B 0.609975f
C59 VDD2.t2 B 0.05129f
C60 VDD2.t0 B 0.05129f
C61 VDD2.n1 B 0.394114f
C62 VDD2.n2 B 1.77647f
C63 VN.t1 B 0.442778f
C64 VN.t2 B 0.441546f
C65 VN.n0 B 0.312332f
C66 VN.t3 B 0.442778f
C67 VN.t0 B 0.441546f
C68 VN.n1 B 0.990353f
.ends

