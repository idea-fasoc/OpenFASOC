* NGSPICE file created from diff_pair_sample_1136.ext - technology: sky130A

.subckt diff_pair_sample_1136 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0.7062 ps=4.61 w=4.28 l=3.76
X1 VDD2.t9 VN.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0.7062 ps=4.61 w=4.28 l=3.76
X2 VDD1.t8 VP.t1 VTAIL.t19 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X3 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0 ps=0 w=4.28 l=3.76
X4 VDD2.t8 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X5 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0 ps=0 w=4.28 l=3.76
X6 VDD1.t7 VP.t2 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=1.6692 ps=9.34 w=4.28 l=3.76
X7 VTAIL.t9 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X8 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X9 VTAIL.t16 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X10 VTAIL.t11 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X11 VTAIL.t13 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X12 VDD2.t5 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0.7062 ps=4.61 w=4.28 l=3.76
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0 ps=0 w=4.28 l=3.76
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0 ps=0 w=4.28 l=3.76
X15 VDD1.t3 VP.t6 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6692 pd=9.34 as=0.7062 ps=4.61 w=4.28 l=3.76
X16 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=1.6692 ps=9.34 w=4.28 l=3.76
X17 VTAIL.t2 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X18 VTAIL.t5 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X19 VTAIL.t10 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X20 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
X21 VDD1.t1 VP.t8 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=1.6692 ps=9.34 w=4.28 l=3.76
X22 VDD2.t0 VN.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=1.6692 ps=9.34 w=4.28 l=3.76
X23 VDD1.t0 VP.t9 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=3.76
R0 VP.n31 VP.n30 161.3
R1 VP.n32 VP.n27 161.3
R2 VP.n34 VP.n33 161.3
R3 VP.n35 VP.n26 161.3
R4 VP.n37 VP.n36 161.3
R5 VP.n38 VP.n25 161.3
R6 VP.n40 VP.n39 161.3
R7 VP.n41 VP.n24 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n23 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n22 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n21 161.3
R14 VP.n53 VP.n52 161.3
R15 VP.n54 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n17 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n67 VP.n16 161.3
R24 VP.n122 VP.n0 161.3
R25 VP.n121 VP.n120 161.3
R26 VP.n119 VP.n1 161.3
R27 VP.n118 VP.n117 161.3
R28 VP.n116 VP.n2 161.3
R29 VP.n115 VP.n114 161.3
R30 VP.n113 VP.n3 161.3
R31 VP.n112 VP.n111 161.3
R32 VP.n109 VP.n4 161.3
R33 VP.n108 VP.n107 161.3
R34 VP.n106 VP.n5 161.3
R35 VP.n105 VP.n104 161.3
R36 VP.n103 VP.n6 161.3
R37 VP.n102 VP.n101 161.3
R38 VP.n100 VP.n7 161.3
R39 VP.n99 VP.n98 161.3
R40 VP.n96 VP.n8 161.3
R41 VP.n95 VP.n94 161.3
R42 VP.n93 VP.n9 161.3
R43 VP.n92 VP.n91 161.3
R44 VP.n90 VP.n10 161.3
R45 VP.n89 VP.n88 161.3
R46 VP.n87 VP.n11 161.3
R47 VP.n86 VP.n85 161.3
R48 VP.n83 VP.n12 161.3
R49 VP.n82 VP.n81 161.3
R50 VP.n80 VP.n13 161.3
R51 VP.n79 VP.n78 161.3
R52 VP.n77 VP.n14 161.3
R53 VP.n76 VP.n75 161.3
R54 VP.n74 VP.n15 161.3
R55 VP.n73 VP.n72 161.3
R56 VP.n71 VP.n70 61.2309
R57 VP.n124 VP.n123 61.2309
R58 VP.n69 VP.n68 61.2309
R59 VP.n28 VP.t6 59.7966
R60 VP.n29 VP.n28 58.5323
R61 VP.n91 VP.n90 56.5617
R62 VP.n104 VP.n103 56.5617
R63 VP.n49 VP.n48 56.5617
R64 VP.n36 VP.n35 56.5617
R65 VP.n70 VP.n69 53.7734
R66 VP.n78 VP.n77 51.7179
R67 VP.n117 VP.n116 51.7179
R68 VP.n62 VP.n61 51.7179
R69 VP.n77 VP.n76 29.4362
R70 VP.n117 VP.n1 29.4362
R71 VP.n62 VP.n17 29.4362
R72 VP.n71 VP.t0 27.4335
R73 VP.n84 VP.t4 27.4335
R74 VP.n97 VP.t1 27.4335
R75 VP.n110 VP.t7 27.4335
R76 VP.n123 VP.t2 27.4335
R77 VP.n68 VP.t8 27.4335
R78 VP.n55 VP.t5 27.4335
R79 VP.n42 VP.t9 27.4335
R80 VP.n29 VP.t3 27.4335
R81 VP.n72 VP.n15 24.5923
R82 VP.n76 VP.n15 24.5923
R83 VP.n78 VP.n13 24.5923
R84 VP.n82 VP.n13 24.5923
R85 VP.n83 VP.n82 24.5923
R86 VP.n85 VP.n11 24.5923
R87 VP.n89 VP.n11 24.5923
R88 VP.n90 VP.n89 24.5923
R89 VP.n91 VP.n9 24.5923
R90 VP.n95 VP.n9 24.5923
R91 VP.n96 VP.n95 24.5923
R92 VP.n98 VP.n7 24.5923
R93 VP.n102 VP.n7 24.5923
R94 VP.n103 VP.n102 24.5923
R95 VP.n104 VP.n5 24.5923
R96 VP.n108 VP.n5 24.5923
R97 VP.n109 VP.n108 24.5923
R98 VP.n111 VP.n3 24.5923
R99 VP.n115 VP.n3 24.5923
R100 VP.n116 VP.n115 24.5923
R101 VP.n121 VP.n1 24.5923
R102 VP.n122 VP.n121 24.5923
R103 VP.n66 VP.n17 24.5923
R104 VP.n67 VP.n66 24.5923
R105 VP.n49 VP.n21 24.5923
R106 VP.n53 VP.n21 24.5923
R107 VP.n54 VP.n53 24.5923
R108 VP.n56 VP.n19 24.5923
R109 VP.n60 VP.n19 24.5923
R110 VP.n61 VP.n60 24.5923
R111 VP.n36 VP.n25 24.5923
R112 VP.n40 VP.n25 24.5923
R113 VP.n41 VP.n40 24.5923
R114 VP.n43 VP.n23 24.5923
R115 VP.n47 VP.n23 24.5923
R116 VP.n48 VP.n47 24.5923
R117 VP.n30 VP.n27 24.5923
R118 VP.n34 VP.n27 24.5923
R119 VP.n35 VP.n34 24.5923
R120 VP.n72 VP.n71 21.1495
R121 VP.n123 VP.n122 21.1495
R122 VP.n68 VP.n67 21.1495
R123 VP.n85 VP.n84 16.7229
R124 VP.n110 VP.n109 16.7229
R125 VP.n55 VP.n54 16.7229
R126 VP.n30 VP.n29 16.7229
R127 VP.n97 VP.n96 12.2964
R128 VP.n98 VP.n97 12.2964
R129 VP.n42 VP.n41 12.2964
R130 VP.n43 VP.n42 12.2964
R131 VP.n84 VP.n83 7.86989
R132 VP.n111 VP.n110 7.86989
R133 VP.n56 VP.n55 7.86989
R134 VP.n31 VP.n28 2.63942
R135 VP.n69 VP.n16 0.417304
R136 VP.n73 VP.n70 0.417304
R137 VP.n124 VP.n0 0.417304
R138 VP VP.n124 0.394524
R139 VP.n32 VP.n31 0.189894
R140 VP.n33 VP.n32 0.189894
R141 VP.n33 VP.n26 0.189894
R142 VP.n37 VP.n26 0.189894
R143 VP.n38 VP.n37 0.189894
R144 VP.n39 VP.n38 0.189894
R145 VP.n39 VP.n24 0.189894
R146 VP.n44 VP.n24 0.189894
R147 VP.n45 VP.n44 0.189894
R148 VP.n46 VP.n45 0.189894
R149 VP.n46 VP.n22 0.189894
R150 VP.n50 VP.n22 0.189894
R151 VP.n51 VP.n50 0.189894
R152 VP.n52 VP.n51 0.189894
R153 VP.n52 VP.n20 0.189894
R154 VP.n57 VP.n20 0.189894
R155 VP.n58 VP.n57 0.189894
R156 VP.n59 VP.n58 0.189894
R157 VP.n59 VP.n18 0.189894
R158 VP.n63 VP.n18 0.189894
R159 VP.n64 VP.n63 0.189894
R160 VP.n65 VP.n64 0.189894
R161 VP.n65 VP.n16 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n75 VP.n74 0.189894
R164 VP.n75 VP.n14 0.189894
R165 VP.n79 VP.n14 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n81 VP.n80 0.189894
R168 VP.n81 VP.n12 0.189894
R169 VP.n86 VP.n12 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n88 VP.n87 0.189894
R172 VP.n88 VP.n10 0.189894
R173 VP.n92 VP.n10 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n94 VP.n93 0.189894
R176 VP.n94 VP.n8 0.189894
R177 VP.n99 VP.n8 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n101 VP.n100 0.189894
R180 VP.n101 VP.n6 0.189894
R181 VP.n105 VP.n6 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n107 VP.n106 0.189894
R184 VP.n107 VP.n4 0.189894
R185 VP.n112 VP.n4 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n114 VP.n113 0.189894
R188 VP.n114 VP.n2 0.189894
R189 VP.n118 VP.n2 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n120 VP.n119 0.189894
R192 VP.n120 VP.n0 0.189894
R193 VTAIL.n11 VTAIL.t1 61.4173
R194 VTAIL.n16 VTAIL.t17 61.4171
R195 VTAIL.n17 VTAIL.t8 61.4171
R196 VTAIL.n2 VTAIL.t12 61.4171
R197 VTAIL.n15 VTAIL.n14 56.7912
R198 VTAIL.n13 VTAIL.n12 56.7912
R199 VTAIL.n10 VTAIL.n9 56.7912
R200 VTAIL.n8 VTAIL.n7 56.7912
R201 VTAIL.n19 VTAIL.n18 56.7909
R202 VTAIL.n1 VTAIL.n0 56.7909
R203 VTAIL.n4 VTAIL.n3 56.7909
R204 VTAIL.n6 VTAIL.n5 56.7909
R205 VTAIL.n8 VTAIL.n6 23.1083
R206 VTAIL.n17 VTAIL.n16 19.5824
R207 VTAIL.n18 VTAIL.t6 4.62667
R208 VTAIL.n18 VTAIL.t2 4.62667
R209 VTAIL.n0 VTAIL.t7 4.62667
R210 VTAIL.n0 VTAIL.t0 4.62667
R211 VTAIL.n3 VTAIL.t19 4.62667
R212 VTAIL.n3 VTAIL.t10 4.62667
R213 VTAIL.n5 VTAIL.t18 4.62667
R214 VTAIL.n5 VTAIL.t11 4.62667
R215 VTAIL.n14 VTAIL.t14 4.62667
R216 VTAIL.n14 VTAIL.t13 4.62667
R217 VTAIL.n12 VTAIL.t15 4.62667
R218 VTAIL.n12 VTAIL.t16 4.62667
R219 VTAIL.n9 VTAIL.t4 4.62667
R220 VTAIL.n9 VTAIL.t9 4.62667
R221 VTAIL.n7 VTAIL.t3 4.62667
R222 VTAIL.n7 VTAIL.t5 4.62667
R223 VTAIL.n10 VTAIL.n8 3.52636
R224 VTAIL.n11 VTAIL.n10 3.52636
R225 VTAIL.n15 VTAIL.n13 3.52636
R226 VTAIL.n16 VTAIL.n15 3.52636
R227 VTAIL.n6 VTAIL.n4 3.52636
R228 VTAIL.n4 VTAIL.n2 3.52636
R229 VTAIL.n19 VTAIL.n17 3.52636
R230 VTAIL VTAIL.n1 2.70309
R231 VTAIL.n13 VTAIL.n11 2.23326
R232 VTAIL.n2 VTAIL.n1 2.23326
R233 VTAIL VTAIL.n19 0.823776
R234 VDD1.n1 VDD1.t3 81.622
R235 VDD1.n3 VDD1.t9 81.6218
R236 VDD1.n5 VDD1.n4 76.0588
R237 VDD1.n1 VDD1.n0 73.47
R238 VDD1.n7 VDD1.n6 73.4698
R239 VDD1.n3 VDD1.n2 73.4697
R240 VDD1.n7 VDD1.n5 46.4987
R241 VDD1.n6 VDD1.t4 4.62667
R242 VDD1.n6 VDD1.t1 4.62667
R243 VDD1.n0 VDD1.t6 4.62667
R244 VDD1.n0 VDD1.t0 4.62667
R245 VDD1.n4 VDD1.t2 4.62667
R246 VDD1.n4 VDD1.t7 4.62667
R247 VDD1.n2 VDD1.t5 4.62667
R248 VDD1.n2 VDD1.t8 4.62667
R249 VDD1 VDD1.n7 2.58671
R250 VDD1 VDD1.n1 0.940155
R251 VDD1.n5 VDD1.n3 0.826619
R252 B.n891 B.n890 585
R253 B.n892 B.n891 585
R254 B.n265 B.n170 585
R255 B.n264 B.n263 585
R256 B.n262 B.n261 585
R257 B.n260 B.n259 585
R258 B.n258 B.n257 585
R259 B.n256 B.n255 585
R260 B.n254 B.n253 585
R261 B.n252 B.n251 585
R262 B.n250 B.n249 585
R263 B.n248 B.n247 585
R264 B.n246 B.n245 585
R265 B.n244 B.n243 585
R266 B.n242 B.n241 585
R267 B.n240 B.n239 585
R268 B.n238 B.n237 585
R269 B.n236 B.n235 585
R270 B.n234 B.n233 585
R271 B.n232 B.n231 585
R272 B.n230 B.n229 585
R273 B.n228 B.n227 585
R274 B.n226 B.n225 585
R275 B.n224 B.n223 585
R276 B.n222 B.n221 585
R277 B.n220 B.n219 585
R278 B.n218 B.n217 585
R279 B.n216 B.n215 585
R280 B.n214 B.n213 585
R281 B.n211 B.n210 585
R282 B.n209 B.n208 585
R283 B.n207 B.n206 585
R284 B.n205 B.n204 585
R285 B.n203 B.n202 585
R286 B.n201 B.n200 585
R287 B.n199 B.n198 585
R288 B.n197 B.n196 585
R289 B.n195 B.n194 585
R290 B.n193 B.n192 585
R291 B.n191 B.n190 585
R292 B.n189 B.n188 585
R293 B.n187 B.n186 585
R294 B.n185 B.n184 585
R295 B.n183 B.n182 585
R296 B.n181 B.n180 585
R297 B.n179 B.n178 585
R298 B.n177 B.n176 585
R299 B.n145 B.n144 585
R300 B.n889 B.n146 585
R301 B.n893 B.n146 585
R302 B.n888 B.n887 585
R303 B.n887 B.n142 585
R304 B.n886 B.n141 585
R305 B.n899 B.n141 585
R306 B.n885 B.n140 585
R307 B.n900 B.n140 585
R308 B.n884 B.n139 585
R309 B.n901 B.n139 585
R310 B.n883 B.n882 585
R311 B.n882 B.n135 585
R312 B.n881 B.n134 585
R313 B.n907 B.n134 585
R314 B.n880 B.n133 585
R315 B.n908 B.n133 585
R316 B.n879 B.n132 585
R317 B.n909 B.n132 585
R318 B.n878 B.n877 585
R319 B.n877 B.n131 585
R320 B.n876 B.n127 585
R321 B.n915 B.n127 585
R322 B.n875 B.n126 585
R323 B.n916 B.n126 585
R324 B.n874 B.n125 585
R325 B.n917 B.n125 585
R326 B.n873 B.n872 585
R327 B.n872 B.n121 585
R328 B.n871 B.n120 585
R329 B.n923 B.n120 585
R330 B.n870 B.n119 585
R331 B.n924 B.n119 585
R332 B.n869 B.n118 585
R333 B.n925 B.n118 585
R334 B.n868 B.n867 585
R335 B.n867 B.n114 585
R336 B.n866 B.n113 585
R337 B.n931 B.n113 585
R338 B.n865 B.n112 585
R339 B.n932 B.n112 585
R340 B.n864 B.n111 585
R341 B.n933 B.n111 585
R342 B.n863 B.n862 585
R343 B.n862 B.n107 585
R344 B.n861 B.n106 585
R345 B.n939 B.n106 585
R346 B.n860 B.n105 585
R347 B.n940 B.n105 585
R348 B.n859 B.n104 585
R349 B.n941 B.n104 585
R350 B.n858 B.n857 585
R351 B.n857 B.n100 585
R352 B.n856 B.n99 585
R353 B.n947 B.n99 585
R354 B.n855 B.n98 585
R355 B.n948 B.n98 585
R356 B.n854 B.n97 585
R357 B.n949 B.n97 585
R358 B.n853 B.n852 585
R359 B.n852 B.n93 585
R360 B.n851 B.n92 585
R361 B.n955 B.n92 585
R362 B.n850 B.n91 585
R363 B.n956 B.n91 585
R364 B.n849 B.n90 585
R365 B.n957 B.n90 585
R366 B.n848 B.n847 585
R367 B.n847 B.n86 585
R368 B.n846 B.n85 585
R369 B.n963 B.n85 585
R370 B.n845 B.n84 585
R371 B.n964 B.n84 585
R372 B.n844 B.n83 585
R373 B.n965 B.n83 585
R374 B.n843 B.n842 585
R375 B.n842 B.n79 585
R376 B.n841 B.n78 585
R377 B.n971 B.n78 585
R378 B.n840 B.n77 585
R379 B.n972 B.n77 585
R380 B.n839 B.n76 585
R381 B.n973 B.n76 585
R382 B.n838 B.n837 585
R383 B.n837 B.n72 585
R384 B.n836 B.n71 585
R385 B.n979 B.n71 585
R386 B.n835 B.n70 585
R387 B.n980 B.n70 585
R388 B.n834 B.n69 585
R389 B.n981 B.n69 585
R390 B.n833 B.n832 585
R391 B.n832 B.n65 585
R392 B.n831 B.n64 585
R393 B.n987 B.n64 585
R394 B.n830 B.n63 585
R395 B.n988 B.n63 585
R396 B.n829 B.n62 585
R397 B.n989 B.n62 585
R398 B.n828 B.n827 585
R399 B.n827 B.n58 585
R400 B.n826 B.n57 585
R401 B.n995 B.n57 585
R402 B.n825 B.n56 585
R403 B.n996 B.n56 585
R404 B.n824 B.n55 585
R405 B.n997 B.n55 585
R406 B.n823 B.n822 585
R407 B.n822 B.n51 585
R408 B.n821 B.n50 585
R409 B.n1003 B.n50 585
R410 B.n820 B.n49 585
R411 B.n1004 B.n49 585
R412 B.n819 B.n48 585
R413 B.n1005 B.n48 585
R414 B.n818 B.n817 585
R415 B.n817 B.n44 585
R416 B.n816 B.n43 585
R417 B.n1011 B.n43 585
R418 B.n815 B.n42 585
R419 B.n1012 B.n42 585
R420 B.n814 B.n41 585
R421 B.n1013 B.n41 585
R422 B.n813 B.n812 585
R423 B.n812 B.n37 585
R424 B.n811 B.n36 585
R425 B.n1019 B.n36 585
R426 B.n810 B.n35 585
R427 B.n1020 B.n35 585
R428 B.n809 B.n34 585
R429 B.n1021 B.n34 585
R430 B.n808 B.n807 585
R431 B.n807 B.n30 585
R432 B.n806 B.n29 585
R433 B.n1027 B.n29 585
R434 B.n805 B.n28 585
R435 B.n1028 B.n28 585
R436 B.n804 B.n27 585
R437 B.n1029 B.n27 585
R438 B.n803 B.n802 585
R439 B.n802 B.n23 585
R440 B.n801 B.n22 585
R441 B.n1035 B.n22 585
R442 B.n800 B.n21 585
R443 B.n1036 B.n21 585
R444 B.n799 B.n20 585
R445 B.n1037 B.n20 585
R446 B.n798 B.n797 585
R447 B.n797 B.n16 585
R448 B.n796 B.n15 585
R449 B.n1043 B.n15 585
R450 B.n795 B.n14 585
R451 B.n1044 B.n14 585
R452 B.n794 B.n13 585
R453 B.n1045 B.n13 585
R454 B.n793 B.n792 585
R455 B.n792 B.n12 585
R456 B.n791 B.n790 585
R457 B.n791 B.n8 585
R458 B.n789 B.n7 585
R459 B.n1052 B.n7 585
R460 B.n788 B.n6 585
R461 B.n1053 B.n6 585
R462 B.n787 B.n5 585
R463 B.n1054 B.n5 585
R464 B.n786 B.n785 585
R465 B.n785 B.n4 585
R466 B.n784 B.n266 585
R467 B.n784 B.n783 585
R468 B.n774 B.n267 585
R469 B.n268 B.n267 585
R470 B.n776 B.n775 585
R471 B.n777 B.n776 585
R472 B.n773 B.n273 585
R473 B.n273 B.n272 585
R474 B.n772 B.n771 585
R475 B.n771 B.n770 585
R476 B.n275 B.n274 585
R477 B.n276 B.n275 585
R478 B.n763 B.n762 585
R479 B.n764 B.n763 585
R480 B.n761 B.n281 585
R481 B.n281 B.n280 585
R482 B.n760 B.n759 585
R483 B.n759 B.n758 585
R484 B.n283 B.n282 585
R485 B.n284 B.n283 585
R486 B.n751 B.n750 585
R487 B.n752 B.n751 585
R488 B.n749 B.n289 585
R489 B.n289 B.n288 585
R490 B.n748 B.n747 585
R491 B.n747 B.n746 585
R492 B.n291 B.n290 585
R493 B.n292 B.n291 585
R494 B.n739 B.n738 585
R495 B.n740 B.n739 585
R496 B.n737 B.n297 585
R497 B.n297 B.n296 585
R498 B.n736 B.n735 585
R499 B.n735 B.n734 585
R500 B.n299 B.n298 585
R501 B.n300 B.n299 585
R502 B.n727 B.n726 585
R503 B.n728 B.n727 585
R504 B.n725 B.n305 585
R505 B.n305 B.n304 585
R506 B.n724 B.n723 585
R507 B.n723 B.n722 585
R508 B.n307 B.n306 585
R509 B.n308 B.n307 585
R510 B.n715 B.n714 585
R511 B.n716 B.n715 585
R512 B.n713 B.n313 585
R513 B.n313 B.n312 585
R514 B.n712 B.n711 585
R515 B.n711 B.n710 585
R516 B.n315 B.n314 585
R517 B.n316 B.n315 585
R518 B.n703 B.n702 585
R519 B.n704 B.n703 585
R520 B.n701 B.n321 585
R521 B.n321 B.n320 585
R522 B.n700 B.n699 585
R523 B.n699 B.n698 585
R524 B.n323 B.n322 585
R525 B.n324 B.n323 585
R526 B.n691 B.n690 585
R527 B.n692 B.n691 585
R528 B.n689 B.n329 585
R529 B.n329 B.n328 585
R530 B.n688 B.n687 585
R531 B.n687 B.n686 585
R532 B.n331 B.n330 585
R533 B.n332 B.n331 585
R534 B.n679 B.n678 585
R535 B.n680 B.n679 585
R536 B.n677 B.n337 585
R537 B.n337 B.n336 585
R538 B.n676 B.n675 585
R539 B.n675 B.n674 585
R540 B.n339 B.n338 585
R541 B.n340 B.n339 585
R542 B.n667 B.n666 585
R543 B.n668 B.n667 585
R544 B.n665 B.n345 585
R545 B.n345 B.n344 585
R546 B.n664 B.n663 585
R547 B.n663 B.n662 585
R548 B.n347 B.n346 585
R549 B.n348 B.n347 585
R550 B.n655 B.n654 585
R551 B.n656 B.n655 585
R552 B.n653 B.n353 585
R553 B.n353 B.n352 585
R554 B.n652 B.n651 585
R555 B.n651 B.n650 585
R556 B.n355 B.n354 585
R557 B.n356 B.n355 585
R558 B.n643 B.n642 585
R559 B.n644 B.n643 585
R560 B.n641 B.n361 585
R561 B.n361 B.n360 585
R562 B.n640 B.n639 585
R563 B.n639 B.n638 585
R564 B.n363 B.n362 585
R565 B.n364 B.n363 585
R566 B.n631 B.n630 585
R567 B.n632 B.n631 585
R568 B.n629 B.n369 585
R569 B.n369 B.n368 585
R570 B.n628 B.n627 585
R571 B.n627 B.n626 585
R572 B.n371 B.n370 585
R573 B.n372 B.n371 585
R574 B.n619 B.n618 585
R575 B.n620 B.n619 585
R576 B.n617 B.n377 585
R577 B.n377 B.n376 585
R578 B.n616 B.n615 585
R579 B.n615 B.n614 585
R580 B.n379 B.n378 585
R581 B.n380 B.n379 585
R582 B.n607 B.n606 585
R583 B.n608 B.n607 585
R584 B.n605 B.n385 585
R585 B.n385 B.n384 585
R586 B.n604 B.n603 585
R587 B.n603 B.n602 585
R588 B.n387 B.n386 585
R589 B.n388 B.n387 585
R590 B.n595 B.n594 585
R591 B.n596 B.n595 585
R592 B.n593 B.n393 585
R593 B.n393 B.n392 585
R594 B.n592 B.n591 585
R595 B.n591 B.n590 585
R596 B.n395 B.n394 585
R597 B.n396 B.n395 585
R598 B.n583 B.n582 585
R599 B.n584 B.n583 585
R600 B.n581 B.n401 585
R601 B.n401 B.n400 585
R602 B.n580 B.n579 585
R603 B.n579 B.n578 585
R604 B.n403 B.n402 585
R605 B.n571 B.n403 585
R606 B.n570 B.n569 585
R607 B.n572 B.n570 585
R608 B.n568 B.n408 585
R609 B.n408 B.n407 585
R610 B.n567 B.n566 585
R611 B.n566 B.n565 585
R612 B.n410 B.n409 585
R613 B.n411 B.n410 585
R614 B.n558 B.n557 585
R615 B.n559 B.n558 585
R616 B.n556 B.n416 585
R617 B.n416 B.n415 585
R618 B.n555 B.n554 585
R619 B.n554 B.n553 585
R620 B.n418 B.n417 585
R621 B.n419 B.n418 585
R622 B.n546 B.n545 585
R623 B.n547 B.n546 585
R624 B.n422 B.n421 585
R625 B.n451 B.n450 585
R626 B.n452 B.n448 585
R627 B.n448 B.n423 585
R628 B.n454 B.n453 585
R629 B.n456 B.n447 585
R630 B.n459 B.n458 585
R631 B.n460 B.n446 585
R632 B.n462 B.n461 585
R633 B.n464 B.n445 585
R634 B.n467 B.n466 585
R635 B.n468 B.n444 585
R636 B.n470 B.n469 585
R637 B.n472 B.n443 585
R638 B.n475 B.n474 585
R639 B.n476 B.n442 585
R640 B.n478 B.n477 585
R641 B.n480 B.n441 585
R642 B.n483 B.n482 585
R643 B.n484 B.n438 585
R644 B.n487 B.n486 585
R645 B.n489 B.n437 585
R646 B.n492 B.n491 585
R647 B.n493 B.n436 585
R648 B.n495 B.n494 585
R649 B.n497 B.n435 585
R650 B.n500 B.n499 585
R651 B.n501 B.n434 585
R652 B.n506 B.n505 585
R653 B.n508 B.n433 585
R654 B.n511 B.n510 585
R655 B.n512 B.n432 585
R656 B.n514 B.n513 585
R657 B.n516 B.n431 585
R658 B.n519 B.n518 585
R659 B.n520 B.n430 585
R660 B.n522 B.n521 585
R661 B.n524 B.n429 585
R662 B.n527 B.n526 585
R663 B.n528 B.n428 585
R664 B.n530 B.n529 585
R665 B.n532 B.n427 585
R666 B.n535 B.n534 585
R667 B.n536 B.n426 585
R668 B.n538 B.n537 585
R669 B.n540 B.n425 585
R670 B.n543 B.n542 585
R671 B.n544 B.n424 585
R672 B.n549 B.n548 585
R673 B.n548 B.n547 585
R674 B.n550 B.n420 585
R675 B.n420 B.n419 585
R676 B.n552 B.n551 585
R677 B.n553 B.n552 585
R678 B.n414 B.n413 585
R679 B.n415 B.n414 585
R680 B.n561 B.n560 585
R681 B.n560 B.n559 585
R682 B.n562 B.n412 585
R683 B.n412 B.n411 585
R684 B.n564 B.n563 585
R685 B.n565 B.n564 585
R686 B.n406 B.n405 585
R687 B.n407 B.n406 585
R688 B.n574 B.n573 585
R689 B.n573 B.n572 585
R690 B.n575 B.n404 585
R691 B.n571 B.n404 585
R692 B.n577 B.n576 585
R693 B.n578 B.n577 585
R694 B.n399 B.n398 585
R695 B.n400 B.n399 585
R696 B.n586 B.n585 585
R697 B.n585 B.n584 585
R698 B.n587 B.n397 585
R699 B.n397 B.n396 585
R700 B.n589 B.n588 585
R701 B.n590 B.n589 585
R702 B.n391 B.n390 585
R703 B.n392 B.n391 585
R704 B.n598 B.n597 585
R705 B.n597 B.n596 585
R706 B.n599 B.n389 585
R707 B.n389 B.n388 585
R708 B.n601 B.n600 585
R709 B.n602 B.n601 585
R710 B.n383 B.n382 585
R711 B.n384 B.n383 585
R712 B.n610 B.n609 585
R713 B.n609 B.n608 585
R714 B.n611 B.n381 585
R715 B.n381 B.n380 585
R716 B.n613 B.n612 585
R717 B.n614 B.n613 585
R718 B.n375 B.n374 585
R719 B.n376 B.n375 585
R720 B.n622 B.n621 585
R721 B.n621 B.n620 585
R722 B.n623 B.n373 585
R723 B.n373 B.n372 585
R724 B.n625 B.n624 585
R725 B.n626 B.n625 585
R726 B.n367 B.n366 585
R727 B.n368 B.n367 585
R728 B.n634 B.n633 585
R729 B.n633 B.n632 585
R730 B.n635 B.n365 585
R731 B.n365 B.n364 585
R732 B.n637 B.n636 585
R733 B.n638 B.n637 585
R734 B.n359 B.n358 585
R735 B.n360 B.n359 585
R736 B.n646 B.n645 585
R737 B.n645 B.n644 585
R738 B.n647 B.n357 585
R739 B.n357 B.n356 585
R740 B.n649 B.n648 585
R741 B.n650 B.n649 585
R742 B.n351 B.n350 585
R743 B.n352 B.n351 585
R744 B.n658 B.n657 585
R745 B.n657 B.n656 585
R746 B.n659 B.n349 585
R747 B.n349 B.n348 585
R748 B.n661 B.n660 585
R749 B.n662 B.n661 585
R750 B.n343 B.n342 585
R751 B.n344 B.n343 585
R752 B.n670 B.n669 585
R753 B.n669 B.n668 585
R754 B.n671 B.n341 585
R755 B.n341 B.n340 585
R756 B.n673 B.n672 585
R757 B.n674 B.n673 585
R758 B.n335 B.n334 585
R759 B.n336 B.n335 585
R760 B.n682 B.n681 585
R761 B.n681 B.n680 585
R762 B.n683 B.n333 585
R763 B.n333 B.n332 585
R764 B.n685 B.n684 585
R765 B.n686 B.n685 585
R766 B.n327 B.n326 585
R767 B.n328 B.n327 585
R768 B.n694 B.n693 585
R769 B.n693 B.n692 585
R770 B.n695 B.n325 585
R771 B.n325 B.n324 585
R772 B.n697 B.n696 585
R773 B.n698 B.n697 585
R774 B.n319 B.n318 585
R775 B.n320 B.n319 585
R776 B.n706 B.n705 585
R777 B.n705 B.n704 585
R778 B.n707 B.n317 585
R779 B.n317 B.n316 585
R780 B.n709 B.n708 585
R781 B.n710 B.n709 585
R782 B.n311 B.n310 585
R783 B.n312 B.n311 585
R784 B.n718 B.n717 585
R785 B.n717 B.n716 585
R786 B.n719 B.n309 585
R787 B.n309 B.n308 585
R788 B.n721 B.n720 585
R789 B.n722 B.n721 585
R790 B.n303 B.n302 585
R791 B.n304 B.n303 585
R792 B.n730 B.n729 585
R793 B.n729 B.n728 585
R794 B.n731 B.n301 585
R795 B.n301 B.n300 585
R796 B.n733 B.n732 585
R797 B.n734 B.n733 585
R798 B.n295 B.n294 585
R799 B.n296 B.n295 585
R800 B.n742 B.n741 585
R801 B.n741 B.n740 585
R802 B.n743 B.n293 585
R803 B.n293 B.n292 585
R804 B.n745 B.n744 585
R805 B.n746 B.n745 585
R806 B.n287 B.n286 585
R807 B.n288 B.n287 585
R808 B.n754 B.n753 585
R809 B.n753 B.n752 585
R810 B.n755 B.n285 585
R811 B.n285 B.n284 585
R812 B.n757 B.n756 585
R813 B.n758 B.n757 585
R814 B.n279 B.n278 585
R815 B.n280 B.n279 585
R816 B.n766 B.n765 585
R817 B.n765 B.n764 585
R818 B.n767 B.n277 585
R819 B.n277 B.n276 585
R820 B.n769 B.n768 585
R821 B.n770 B.n769 585
R822 B.n271 B.n270 585
R823 B.n272 B.n271 585
R824 B.n779 B.n778 585
R825 B.n778 B.n777 585
R826 B.n780 B.n269 585
R827 B.n269 B.n268 585
R828 B.n782 B.n781 585
R829 B.n783 B.n782 585
R830 B.n3 B.n0 585
R831 B.n4 B.n3 585
R832 B.n1051 B.n1 585
R833 B.n1052 B.n1051 585
R834 B.n1050 B.n1049 585
R835 B.n1050 B.n8 585
R836 B.n1048 B.n9 585
R837 B.n12 B.n9 585
R838 B.n1047 B.n1046 585
R839 B.n1046 B.n1045 585
R840 B.n11 B.n10 585
R841 B.n1044 B.n11 585
R842 B.n1042 B.n1041 585
R843 B.n1043 B.n1042 585
R844 B.n1040 B.n17 585
R845 B.n17 B.n16 585
R846 B.n1039 B.n1038 585
R847 B.n1038 B.n1037 585
R848 B.n19 B.n18 585
R849 B.n1036 B.n19 585
R850 B.n1034 B.n1033 585
R851 B.n1035 B.n1034 585
R852 B.n1032 B.n24 585
R853 B.n24 B.n23 585
R854 B.n1031 B.n1030 585
R855 B.n1030 B.n1029 585
R856 B.n26 B.n25 585
R857 B.n1028 B.n26 585
R858 B.n1026 B.n1025 585
R859 B.n1027 B.n1026 585
R860 B.n1024 B.n31 585
R861 B.n31 B.n30 585
R862 B.n1023 B.n1022 585
R863 B.n1022 B.n1021 585
R864 B.n33 B.n32 585
R865 B.n1020 B.n33 585
R866 B.n1018 B.n1017 585
R867 B.n1019 B.n1018 585
R868 B.n1016 B.n38 585
R869 B.n38 B.n37 585
R870 B.n1015 B.n1014 585
R871 B.n1014 B.n1013 585
R872 B.n40 B.n39 585
R873 B.n1012 B.n40 585
R874 B.n1010 B.n1009 585
R875 B.n1011 B.n1010 585
R876 B.n1008 B.n45 585
R877 B.n45 B.n44 585
R878 B.n1007 B.n1006 585
R879 B.n1006 B.n1005 585
R880 B.n47 B.n46 585
R881 B.n1004 B.n47 585
R882 B.n1002 B.n1001 585
R883 B.n1003 B.n1002 585
R884 B.n1000 B.n52 585
R885 B.n52 B.n51 585
R886 B.n999 B.n998 585
R887 B.n998 B.n997 585
R888 B.n54 B.n53 585
R889 B.n996 B.n54 585
R890 B.n994 B.n993 585
R891 B.n995 B.n994 585
R892 B.n992 B.n59 585
R893 B.n59 B.n58 585
R894 B.n991 B.n990 585
R895 B.n990 B.n989 585
R896 B.n61 B.n60 585
R897 B.n988 B.n61 585
R898 B.n986 B.n985 585
R899 B.n987 B.n986 585
R900 B.n984 B.n66 585
R901 B.n66 B.n65 585
R902 B.n983 B.n982 585
R903 B.n982 B.n981 585
R904 B.n68 B.n67 585
R905 B.n980 B.n68 585
R906 B.n978 B.n977 585
R907 B.n979 B.n978 585
R908 B.n976 B.n73 585
R909 B.n73 B.n72 585
R910 B.n975 B.n974 585
R911 B.n974 B.n973 585
R912 B.n75 B.n74 585
R913 B.n972 B.n75 585
R914 B.n970 B.n969 585
R915 B.n971 B.n970 585
R916 B.n968 B.n80 585
R917 B.n80 B.n79 585
R918 B.n967 B.n966 585
R919 B.n966 B.n965 585
R920 B.n82 B.n81 585
R921 B.n964 B.n82 585
R922 B.n962 B.n961 585
R923 B.n963 B.n962 585
R924 B.n960 B.n87 585
R925 B.n87 B.n86 585
R926 B.n959 B.n958 585
R927 B.n958 B.n957 585
R928 B.n89 B.n88 585
R929 B.n956 B.n89 585
R930 B.n954 B.n953 585
R931 B.n955 B.n954 585
R932 B.n952 B.n94 585
R933 B.n94 B.n93 585
R934 B.n951 B.n950 585
R935 B.n950 B.n949 585
R936 B.n96 B.n95 585
R937 B.n948 B.n96 585
R938 B.n946 B.n945 585
R939 B.n947 B.n946 585
R940 B.n944 B.n101 585
R941 B.n101 B.n100 585
R942 B.n943 B.n942 585
R943 B.n942 B.n941 585
R944 B.n103 B.n102 585
R945 B.n940 B.n103 585
R946 B.n938 B.n937 585
R947 B.n939 B.n938 585
R948 B.n936 B.n108 585
R949 B.n108 B.n107 585
R950 B.n935 B.n934 585
R951 B.n934 B.n933 585
R952 B.n110 B.n109 585
R953 B.n932 B.n110 585
R954 B.n930 B.n929 585
R955 B.n931 B.n930 585
R956 B.n928 B.n115 585
R957 B.n115 B.n114 585
R958 B.n927 B.n926 585
R959 B.n926 B.n925 585
R960 B.n117 B.n116 585
R961 B.n924 B.n117 585
R962 B.n922 B.n921 585
R963 B.n923 B.n922 585
R964 B.n920 B.n122 585
R965 B.n122 B.n121 585
R966 B.n919 B.n918 585
R967 B.n918 B.n917 585
R968 B.n124 B.n123 585
R969 B.n916 B.n124 585
R970 B.n914 B.n913 585
R971 B.n915 B.n914 585
R972 B.n912 B.n128 585
R973 B.n131 B.n128 585
R974 B.n911 B.n910 585
R975 B.n910 B.n909 585
R976 B.n130 B.n129 585
R977 B.n908 B.n130 585
R978 B.n906 B.n905 585
R979 B.n907 B.n906 585
R980 B.n904 B.n136 585
R981 B.n136 B.n135 585
R982 B.n903 B.n902 585
R983 B.n902 B.n901 585
R984 B.n138 B.n137 585
R985 B.n900 B.n138 585
R986 B.n898 B.n897 585
R987 B.n899 B.n898 585
R988 B.n896 B.n143 585
R989 B.n143 B.n142 585
R990 B.n895 B.n894 585
R991 B.n894 B.n893 585
R992 B.n1055 B.n1054 585
R993 B.n1053 B.n2 585
R994 B.n894 B.n145 497.305
R995 B.n891 B.n146 497.305
R996 B.n546 B.n424 497.305
R997 B.n548 B.n422 497.305
R998 B.n892 B.n169 256.663
R999 B.n892 B.n168 256.663
R1000 B.n892 B.n167 256.663
R1001 B.n892 B.n166 256.663
R1002 B.n892 B.n165 256.663
R1003 B.n892 B.n164 256.663
R1004 B.n892 B.n163 256.663
R1005 B.n892 B.n162 256.663
R1006 B.n892 B.n161 256.663
R1007 B.n892 B.n160 256.663
R1008 B.n892 B.n159 256.663
R1009 B.n892 B.n158 256.663
R1010 B.n892 B.n157 256.663
R1011 B.n892 B.n156 256.663
R1012 B.n892 B.n155 256.663
R1013 B.n892 B.n154 256.663
R1014 B.n892 B.n153 256.663
R1015 B.n892 B.n152 256.663
R1016 B.n892 B.n151 256.663
R1017 B.n892 B.n150 256.663
R1018 B.n892 B.n149 256.663
R1019 B.n892 B.n148 256.663
R1020 B.n892 B.n147 256.663
R1021 B.n449 B.n423 256.663
R1022 B.n455 B.n423 256.663
R1023 B.n457 B.n423 256.663
R1024 B.n463 B.n423 256.663
R1025 B.n465 B.n423 256.663
R1026 B.n471 B.n423 256.663
R1027 B.n473 B.n423 256.663
R1028 B.n479 B.n423 256.663
R1029 B.n481 B.n423 256.663
R1030 B.n488 B.n423 256.663
R1031 B.n490 B.n423 256.663
R1032 B.n496 B.n423 256.663
R1033 B.n498 B.n423 256.663
R1034 B.n507 B.n423 256.663
R1035 B.n509 B.n423 256.663
R1036 B.n515 B.n423 256.663
R1037 B.n517 B.n423 256.663
R1038 B.n523 B.n423 256.663
R1039 B.n525 B.n423 256.663
R1040 B.n531 B.n423 256.663
R1041 B.n533 B.n423 256.663
R1042 B.n539 B.n423 256.663
R1043 B.n541 B.n423 256.663
R1044 B.n1057 B.n1056 256.663
R1045 B.n174 B.t21 236.745
R1046 B.n171 B.t14 236.745
R1047 B.n502 B.t18 236.745
R1048 B.n439 B.t10 236.745
R1049 B.n178 B.n177 163.367
R1050 B.n182 B.n181 163.367
R1051 B.n186 B.n185 163.367
R1052 B.n190 B.n189 163.367
R1053 B.n194 B.n193 163.367
R1054 B.n198 B.n197 163.367
R1055 B.n202 B.n201 163.367
R1056 B.n206 B.n205 163.367
R1057 B.n210 B.n209 163.367
R1058 B.n215 B.n214 163.367
R1059 B.n219 B.n218 163.367
R1060 B.n223 B.n222 163.367
R1061 B.n227 B.n226 163.367
R1062 B.n231 B.n230 163.367
R1063 B.n235 B.n234 163.367
R1064 B.n239 B.n238 163.367
R1065 B.n243 B.n242 163.367
R1066 B.n247 B.n246 163.367
R1067 B.n251 B.n250 163.367
R1068 B.n255 B.n254 163.367
R1069 B.n259 B.n258 163.367
R1070 B.n263 B.n262 163.367
R1071 B.n891 B.n170 163.367
R1072 B.n546 B.n418 163.367
R1073 B.n554 B.n418 163.367
R1074 B.n554 B.n416 163.367
R1075 B.n558 B.n416 163.367
R1076 B.n558 B.n410 163.367
R1077 B.n566 B.n410 163.367
R1078 B.n566 B.n408 163.367
R1079 B.n570 B.n408 163.367
R1080 B.n570 B.n403 163.367
R1081 B.n579 B.n403 163.367
R1082 B.n579 B.n401 163.367
R1083 B.n583 B.n401 163.367
R1084 B.n583 B.n395 163.367
R1085 B.n591 B.n395 163.367
R1086 B.n591 B.n393 163.367
R1087 B.n595 B.n393 163.367
R1088 B.n595 B.n387 163.367
R1089 B.n603 B.n387 163.367
R1090 B.n603 B.n385 163.367
R1091 B.n607 B.n385 163.367
R1092 B.n607 B.n379 163.367
R1093 B.n615 B.n379 163.367
R1094 B.n615 B.n377 163.367
R1095 B.n619 B.n377 163.367
R1096 B.n619 B.n371 163.367
R1097 B.n627 B.n371 163.367
R1098 B.n627 B.n369 163.367
R1099 B.n631 B.n369 163.367
R1100 B.n631 B.n363 163.367
R1101 B.n639 B.n363 163.367
R1102 B.n639 B.n361 163.367
R1103 B.n643 B.n361 163.367
R1104 B.n643 B.n355 163.367
R1105 B.n651 B.n355 163.367
R1106 B.n651 B.n353 163.367
R1107 B.n655 B.n353 163.367
R1108 B.n655 B.n347 163.367
R1109 B.n663 B.n347 163.367
R1110 B.n663 B.n345 163.367
R1111 B.n667 B.n345 163.367
R1112 B.n667 B.n339 163.367
R1113 B.n675 B.n339 163.367
R1114 B.n675 B.n337 163.367
R1115 B.n679 B.n337 163.367
R1116 B.n679 B.n331 163.367
R1117 B.n687 B.n331 163.367
R1118 B.n687 B.n329 163.367
R1119 B.n691 B.n329 163.367
R1120 B.n691 B.n323 163.367
R1121 B.n699 B.n323 163.367
R1122 B.n699 B.n321 163.367
R1123 B.n703 B.n321 163.367
R1124 B.n703 B.n315 163.367
R1125 B.n711 B.n315 163.367
R1126 B.n711 B.n313 163.367
R1127 B.n715 B.n313 163.367
R1128 B.n715 B.n307 163.367
R1129 B.n723 B.n307 163.367
R1130 B.n723 B.n305 163.367
R1131 B.n727 B.n305 163.367
R1132 B.n727 B.n299 163.367
R1133 B.n735 B.n299 163.367
R1134 B.n735 B.n297 163.367
R1135 B.n739 B.n297 163.367
R1136 B.n739 B.n291 163.367
R1137 B.n747 B.n291 163.367
R1138 B.n747 B.n289 163.367
R1139 B.n751 B.n289 163.367
R1140 B.n751 B.n283 163.367
R1141 B.n759 B.n283 163.367
R1142 B.n759 B.n281 163.367
R1143 B.n763 B.n281 163.367
R1144 B.n763 B.n275 163.367
R1145 B.n771 B.n275 163.367
R1146 B.n771 B.n273 163.367
R1147 B.n776 B.n273 163.367
R1148 B.n776 B.n267 163.367
R1149 B.n784 B.n267 163.367
R1150 B.n785 B.n784 163.367
R1151 B.n785 B.n5 163.367
R1152 B.n6 B.n5 163.367
R1153 B.n7 B.n6 163.367
R1154 B.n791 B.n7 163.367
R1155 B.n792 B.n791 163.367
R1156 B.n792 B.n13 163.367
R1157 B.n14 B.n13 163.367
R1158 B.n15 B.n14 163.367
R1159 B.n797 B.n15 163.367
R1160 B.n797 B.n20 163.367
R1161 B.n21 B.n20 163.367
R1162 B.n22 B.n21 163.367
R1163 B.n802 B.n22 163.367
R1164 B.n802 B.n27 163.367
R1165 B.n28 B.n27 163.367
R1166 B.n29 B.n28 163.367
R1167 B.n807 B.n29 163.367
R1168 B.n807 B.n34 163.367
R1169 B.n35 B.n34 163.367
R1170 B.n36 B.n35 163.367
R1171 B.n812 B.n36 163.367
R1172 B.n812 B.n41 163.367
R1173 B.n42 B.n41 163.367
R1174 B.n43 B.n42 163.367
R1175 B.n817 B.n43 163.367
R1176 B.n817 B.n48 163.367
R1177 B.n49 B.n48 163.367
R1178 B.n50 B.n49 163.367
R1179 B.n822 B.n50 163.367
R1180 B.n822 B.n55 163.367
R1181 B.n56 B.n55 163.367
R1182 B.n57 B.n56 163.367
R1183 B.n827 B.n57 163.367
R1184 B.n827 B.n62 163.367
R1185 B.n63 B.n62 163.367
R1186 B.n64 B.n63 163.367
R1187 B.n832 B.n64 163.367
R1188 B.n832 B.n69 163.367
R1189 B.n70 B.n69 163.367
R1190 B.n71 B.n70 163.367
R1191 B.n837 B.n71 163.367
R1192 B.n837 B.n76 163.367
R1193 B.n77 B.n76 163.367
R1194 B.n78 B.n77 163.367
R1195 B.n842 B.n78 163.367
R1196 B.n842 B.n83 163.367
R1197 B.n84 B.n83 163.367
R1198 B.n85 B.n84 163.367
R1199 B.n847 B.n85 163.367
R1200 B.n847 B.n90 163.367
R1201 B.n91 B.n90 163.367
R1202 B.n92 B.n91 163.367
R1203 B.n852 B.n92 163.367
R1204 B.n852 B.n97 163.367
R1205 B.n98 B.n97 163.367
R1206 B.n99 B.n98 163.367
R1207 B.n857 B.n99 163.367
R1208 B.n857 B.n104 163.367
R1209 B.n105 B.n104 163.367
R1210 B.n106 B.n105 163.367
R1211 B.n862 B.n106 163.367
R1212 B.n862 B.n111 163.367
R1213 B.n112 B.n111 163.367
R1214 B.n113 B.n112 163.367
R1215 B.n867 B.n113 163.367
R1216 B.n867 B.n118 163.367
R1217 B.n119 B.n118 163.367
R1218 B.n120 B.n119 163.367
R1219 B.n872 B.n120 163.367
R1220 B.n872 B.n125 163.367
R1221 B.n126 B.n125 163.367
R1222 B.n127 B.n126 163.367
R1223 B.n877 B.n127 163.367
R1224 B.n877 B.n132 163.367
R1225 B.n133 B.n132 163.367
R1226 B.n134 B.n133 163.367
R1227 B.n882 B.n134 163.367
R1228 B.n882 B.n139 163.367
R1229 B.n140 B.n139 163.367
R1230 B.n141 B.n140 163.367
R1231 B.n887 B.n141 163.367
R1232 B.n887 B.n146 163.367
R1233 B.n450 B.n448 163.367
R1234 B.n454 B.n448 163.367
R1235 B.n458 B.n456 163.367
R1236 B.n462 B.n446 163.367
R1237 B.n466 B.n464 163.367
R1238 B.n470 B.n444 163.367
R1239 B.n474 B.n472 163.367
R1240 B.n478 B.n442 163.367
R1241 B.n482 B.n480 163.367
R1242 B.n487 B.n438 163.367
R1243 B.n491 B.n489 163.367
R1244 B.n495 B.n436 163.367
R1245 B.n499 B.n497 163.367
R1246 B.n506 B.n434 163.367
R1247 B.n510 B.n508 163.367
R1248 B.n514 B.n432 163.367
R1249 B.n518 B.n516 163.367
R1250 B.n522 B.n430 163.367
R1251 B.n526 B.n524 163.367
R1252 B.n530 B.n428 163.367
R1253 B.n534 B.n532 163.367
R1254 B.n538 B.n426 163.367
R1255 B.n542 B.n540 163.367
R1256 B.n548 B.n420 163.367
R1257 B.n552 B.n420 163.367
R1258 B.n552 B.n414 163.367
R1259 B.n560 B.n414 163.367
R1260 B.n560 B.n412 163.367
R1261 B.n564 B.n412 163.367
R1262 B.n564 B.n406 163.367
R1263 B.n573 B.n406 163.367
R1264 B.n573 B.n404 163.367
R1265 B.n577 B.n404 163.367
R1266 B.n577 B.n399 163.367
R1267 B.n585 B.n399 163.367
R1268 B.n585 B.n397 163.367
R1269 B.n589 B.n397 163.367
R1270 B.n589 B.n391 163.367
R1271 B.n597 B.n391 163.367
R1272 B.n597 B.n389 163.367
R1273 B.n601 B.n389 163.367
R1274 B.n601 B.n383 163.367
R1275 B.n609 B.n383 163.367
R1276 B.n609 B.n381 163.367
R1277 B.n613 B.n381 163.367
R1278 B.n613 B.n375 163.367
R1279 B.n621 B.n375 163.367
R1280 B.n621 B.n373 163.367
R1281 B.n625 B.n373 163.367
R1282 B.n625 B.n367 163.367
R1283 B.n633 B.n367 163.367
R1284 B.n633 B.n365 163.367
R1285 B.n637 B.n365 163.367
R1286 B.n637 B.n359 163.367
R1287 B.n645 B.n359 163.367
R1288 B.n645 B.n357 163.367
R1289 B.n649 B.n357 163.367
R1290 B.n649 B.n351 163.367
R1291 B.n657 B.n351 163.367
R1292 B.n657 B.n349 163.367
R1293 B.n661 B.n349 163.367
R1294 B.n661 B.n343 163.367
R1295 B.n669 B.n343 163.367
R1296 B.n669 B.n341 163.367
R1297 B.n673 B.n341 163.367
R1298 B.n673 B.n335 163.367
R1299 B.n681 B.n335 163.367
R1300 B.n681 B.n333 163.367
R1301 B.n685 B.n333 163.367
R1302 B.n685 B.n327 163.367
R1303 B.n693 B.n327 163.367
R1304 B.n693 B.n325 163.367
R1305 B.n697 B.n325 163.367
R1306 B.n697 B.n319 163.367
R1307 B.n705 B.n319 163.367
R1308 B.n705 B.n317 163.367
R1309 B.n709 B.n317 163.367
R1310 B.n709 B.n311 163.367
R1311 B.n717 B.n311 163.367
R1312 B.n717 B.n309 163.367
R1313 B.n721 B.n309 163.367
R1314 B.n721 B.n303 163.367
R1315 B.n729 B.n303 163.367
R1316 B.n729 B.n301 163.367
R1317 B.n733 B.n301 163.367
R1318 B.n733 B.n295 163.367
R1319 B.n741 B.n295 163.367
R1320 B.n741 B.n293 163.367
R1321 B.n745 B.n293 163.367
R1322 B.n745 B.n287 163.367
R1323 B.n753 B.n287 163.367
R1324 B.n753 B.n285 163.367
R1325 B.n757 B.n285 163.367
R1326 B.n757 B.n279 163.367
R1327 B.n765 B.n279 163.367
R1328 B.n765 B.n277 163.367
R1329 B.n769 B.n277 163.367
R1330 B.n769 B.n271 163.367
R1331 B.n778 B.n271 163.367
R1332 B.n778 B.n269 163.367
R1333 B.n782 B.n269 163.367
R1334 B.n782 B.n3 163.367
R1335 B.n1055 B.n3 163.367
R1336 B.n1051 B.n2 163.367
R1337 B.n1051 B.n1050 163.367
R1338 B.n1050 B.n9 163.367
R1339 B.n1046 B.n9 163.367
R1340 B.n1046 B.n11 163.367
R1341 B.n1042 B.n11 163.367
R1342 B.n1042 B.n17 163.367
R1343 B.n1038 B.n17 163.367
R1344 B.n1038 B.n19 163.367
R1345 B.n1034 B.n19 163.367
R1346 B.n1034 B.n24 163.367
R1347 B.n1030 B.n24 163.367
R1348 B.n1030 B.n26 163.367
R1349 B.n1026 B.n26 163.367
R1350 B.n1026 B.n31 163.367
R1351 B.n1022 B.n31 163.367
R1352 B.n1022 B.n33 163.367
R1353 B.n1018 B.n33 163.367
R1354 B.n1018 B.n38 163.367
R1355 B.n1014 B.n38 163.367
R1356 B.n1014 B.n40 163.367
R1357 B.n1010 B.n40 163.367
R1358 B.n1010 B.n45 163.367
R1359 B.n1006 B.n45 163.367
R1360 B.n1006 B.n47 163.367
R1361 B.n1002 B.n47 163.367
R1362 B.n1002 B.n52 163.367
R1363 B.n998 B.n52 163.367
R1364 B.n998 B.n54 163.367
R1365 B.n994 B.n54 163.367
R1366 B.n994 B.n59 163.367
R1367 B.n990 B.n59 163.367
R1368 B.n990 B.n61 163.367
R1369 B.n986 B.n61 163.367
R1370 B.n986 B.n66 163.367
R1371 B.n982 B.n66 163.367
R1372 B.n982 B.n68 163.367
R1373 B.n978 B.n68 163.367
R1374 B.n978 B.n73 163.367
R1375 B.n974 B.n73 163.367
R1376 B.n974 B.n75 163.367
R1377 B.n970 B.n75 163.367
R1378 B.n970 B.n80 163.367
R1379 B.n966 B.n80 163.367
R1380 B.n966 B.n82 163.367
R1381 B.n962 B.n82 163.367
R1382 B.n962 B.n87 163.367
R1383 B.n958 B.n87 163.367
R1384 B.n958 B.n89 163.367
R1385 B.n954 B.n89 163.367
R1386 B.n954 B.n94 163.367
R1387 B.n950 B.n94 163.367
R1388 B.n950 B.n96 163.367
R1389 B.n946 B.n96 163.367
R1390 B.n946 B.n101 163.367
R1391 B.n942 B.n101 163.367
R1392 B.n942 B.n103 163.367
R1393 B.n938 B.n103 163.367
R1394 B.n938 B.n108 163.367
R1395 B.n934 B.n108 163.367
R1396 B.n934 B.n110 163.367
R1397 B.n930 B.n110 163.367
R1398 B.n930 B.n115 163.367
R1399 B.n926 B.n115 163.367
R1400 B.n926 B.n117 163.367
R1401 B.n922 B.n117 163.367
R1402 B.n922 B.n122 163.367
R1403 B.n918 B.n122 163.367
R1404 B.n918 B.n124 163.367
R1405 B.n914 B.n124 163.367
R1406 B.n914 B.n128 163.367
R1407 B.n910 B.n128 163.367
R1408 B.n910 B.n130 163.367
R1409 B.n906 B.n130 163.367
R1410 B.n906 B.n136 163.367
R1411 B.n902 B.n136 163.367
R1412 B.n902 B.n138 163.367
R1413 B.n898 B.n138 163.367
R1414 B.n898 B.n143 163.367
R1415 B.n894 B.n143 163.367
R1416 B.n171 B.t16 154.24
R1417 B.n502 B.t20 154.24
R1418 B.n174 B.t22 154.237
R1419 B.n439 B.t13 154.237
R1420 B.n547 B.n423 125.484
R1421 B.n893 B.n892 125.484
R1422 B.n175 B.n174 79.3217
R1423 B.n172 B.n171 79.3217
R1424 B.n503 B.n502 79.3217
R1425 B.n440 B.n439 79.3217
R1426 B.n547 B.n419 78.2841
R1427 B.n553 B.n419 78.2841
R1428 B.n553 B.n415 78.2841
R1429 B.n559 B.n415 78.2841
R1430 B.n559 B.n411 78.2841
R1431 B.n565 B.n411 78.2841
R1432 B.n565 B.n407 78.2841
R1433 B.n572 B.n407 78.2841
R1434 B.n572 B.n571 78.2841
R1435 B.n578 B.n400 78.2841
R1436 B.n584 B.n400 78.2841
R1437 B.n584 B.n396 78.2841
R1438 B.n590 B.n396 78.2841
R1439 B.n590 B.n392 78.2841
R1440 B.n596 B.n392 78.2841
R1441 B.n596 B.n388 78.2841
R1442 B.n602 B.n388 78.2841
R1443 B.n602 B.n384 78.2841
R1444 B.n608 B.n384 78.2841
R1445 B.n608 B.n380 78.2841
R1446 B.n614 B.n380 78.2841
R1447 B.n614 B.n376 78.2841
R1448 B.n620 B.n376 78.2841
R1449 B.n626 B.n372 78.2841
R1450 B.n626 B.n368 78.2841
R1451 B.n632 B.n368 78.2841
R1452 B.n632 B.n364 78.2841
R1453 B.n638 B.n364 78.2841
R1454 B.n638 B.n360 78.2841
R1455 B.n644 B.n360 78.2841
R1456 B.n644 B.n356 78.2841
R1457 B.n650 B.n356 78.2841
R1458 B.n650 B.n352 78.2841
R1459 B.n656 B.n352 78.2841
R1460 B.n662 B.n348 78.2841
R1461 B.n662 B.n344 78.2841
R1462 B.n668 B.n344 78.2841
R1463 B.n668 B.n340 78.2841
R1464 B.n674 B.n340 78.2841
R1465 B.n674 B.n336 78.2841
R1466 B.n680 B.n336 78.2841
R1467 B.n680 B.n332 78.2841
R1468 B.n686 B.n332 78.2841
R1469 B.n686 B.n328 78.2841
R1470 B.n692 B.n328 78.2841
R1471 B.n698 B.n324 78.2841
R1472 B.n698 B.n320 78.2841
R1473 B.n704 B.n320 78.2841
R1474 B.n704 B.n316 78.2841
R1475 B.n710 B.n316 78.2841
R1476 B.n710 B.n312 78.2841
R1477 B.n716 B.n312 78.2841
R1478 B.n716 B.n308 78.2841
R1479 B.n722 B.n308 78.2841
R1480 B.n722 B.n304 78.2841
R1481 B.n728 B.n304 78.2841
R1482 B.n734 B.n300 78.2841
R1483 B.n734 B.n296 78.2841
R1484 B.n740 B.n296 78.2841
R1485 B.n740 B.n292 78.2841
R1486 B.n746 B.n292 78.2841
R1487 B.n746 B.n288 78.2841
R1488 B.n752 B.n288 78.2841
R1489 B.n752 B.n284 78.2841
R1490 B.n758 B.n284 78.2841
R1491 B.n758 B.n280 78.2841
R1492 B.n764 B.n280 78.2841
R1493 B.n770 B.n276 78.2841
R1494 B.n770 B.n272 78.2841
R1495 B.n777 B.n272 78.2841
R1496 B.n777 B.n268 78.2841
R1497 B.n783 B.n268 78.2841
R1498 B.n783 B.n4 78.2841
R1499 B.n1054 B.n4 78.2841
R1500 B.n1054 B.n1053 78.2841
R1501 B.n1053 B.n1052 78.2841
R1502 B.n1052 B.n8 78.2841
R1503 B.n12 B.n8 78.2841
R1504 B.n1045 B.n12 78.2841
R1505 B.n1045 B.n1044 78.2841
R1506 B.n1044 B.n1043 78.2841
R1507 B.n1043 B.n16 78.2841
R1508 B.n1037 B.n1036 78.2841
R1509 B.n1036 B.n1035 78.2841
R1510 B.n1035 B.n23 78.2841
R1511 B.n1029 B.n23 78.2841
R1512 B.n1029 B.n1028 78.2841
R1513 B.n1028 B.n1027 78.2841
R1514 B.n1027 B.n30 78.2841
R1515 B.n1021 B.n30 78.2841
R1516 B.n1021 B.n1020 78.2841
R1517 B.n1020 B.n1019 78.2841
R1518 B.n1019 B.n37 78.2841
R1519 B.n1013 B.n1012 78.2841
R1520 B.n1012 B.n1011 78.2841
R1521 B.n1011 B.n44 78.2841
R1522 B.n1005 B.n44 78.2841
R1523 B.n1005 B.n1004 78.2841
R1524 B.n1004 B.n1003 78.2841
R1525 B.n1003 B.n51 78.2841
R1526 B.n997 B.n51 78.2841
R1527 B.n997 B.n996 78.2841
R1528 B.n996 B.n995 78.2841
R1529 B.n995 B.n58 78.2841
R1530 B.n989 B.n988 78.2841
R1531 B.n988 B.n987 78.2841
R1532 B.n987 B.n65 78.2841
R1533 B.n981 B.n65 78.2841
R1534 B.n981 B.n980 78.2841
R1535 B.n980 B.n979 78.2841
R1536 B.n979 B.n72 78.2841
R1537 B.n973 B.n72 78.2841
R1538 B.n973 B.n972 78.2841
R1539 B.n972 B.n971 78.2841
R1540 B.n971 B.n79 78.2841
R1541 B.n965 B.n964 78.2841
R1542 B.n964 B.n963 78.2841
R1543 B.n963 B.n86 78.2841
R1544 B.n957 B.n86 78.2841
R1545 B.n957 B.n956 78.2841
R1546 B.n956 B.n955 78.2841
R1547 B.n955 B.n93 78.2841
R1548 B.n949 B.n93 78.2841
R1549 B.n949 B.n948 78.2841
R1550 B.n948 B.n947 78.2841
R1551 B.n947 B.n100 78.2841
R1552 B.n941 B.n940 78.2841
R1553 B.n940 B.n939 78.2841
R1554 B.n939 B.n107 78.2841
R1555 B.n933 B.n107 78.2841
R1556 B.n933 B.n932 78.2841
R1557 B.n932 B.n931 78.2841
R1558 B.n931 B.n114 78.2841
R1559 B.n925 B.n114 78.2841
R1560 B.n925 B.n924 78.2841
R1561 B.n924 B.n923 78.2841
R1562 B.n923 B.n121 78.2841
R1563 B.n917 B.n121 78.2841
R1564 B.n917 B.n916 78.2841
R1565 B.n916 B.n915 78.2841
R1566 B.n909 B.n131 78.2841
R1567 B.n909 B.n908 78.2841
R1568 B.n908 B.n907 78.2841
R1569 B.n907 B.n135 78.2841
R1570 B.n901 B.n135 78.2841
R1571 B.n901 B.n900 78.2841
R1572 B.n900 B.n899 78.2841
R1573 B.n899 B.n142 78.2841
R1574 B.n893 B.n142 78.2841
R1575 B.n172 B.t17 74.9195
R1576 B.n503 B.t19 74.9195
R1577 B.n175 B.t23 74.9156
R1578 B.n440 B.t12 74.9156
R1579 B.n147 B.n145 71.676
R1580 B.n178 B.n148 71.676
R1581 B.n182 B.n149 71.676
R1582 B.n186 B.n150 71.676
R1583 B.n190 B.n151 71.676
R1584 B.n194 B.n152 71.676
R1585 B.n198 B.n153 71.676
R1586 B.n202 B.n154 71.676
R1587 B.n206 B.n155 71.676
R1588 B.n210 B.n156 71.676
R1589 B.n215 B.n157 71.676
R1590 B.n219 B.n158 71.676
R1591 B.n223 B.n159 71.676
R1592 B.n227 B.n160 71.676
R1593 B.n231 B.n161 71.676
R1594 B.n235 B.n162 71.676
R1595 B.n239 B.n163 71.676
R1596 B.n243 B.n164 71.676
R1597 B.n247 B.n165 71.676
R1598 B.n251 B.n166 71.676
R1599 B.n255 B.n167 71.676
R1600 B.n259 B.n168 71.676
R1601 B.n263 B.n169 71.676
R1602 B.n170 B.n169 71.676
R1603 B.n262 B.n168 71.676
R1604 B.n258 B.n167 71.676
R1605 B.n254 B.n166 71.676
R1606 B.n250 B.n165 71.676
R1607 B.n246 B.n164 71.676
R1608 B.n242 B.n163 71.676
R1609 B.n238 B.n162 71.676
R1610 B.n234 B.n161 71.676
R1611 B.n230 B.n160 71.676
R1612 B.n226 B.n159 71.676
R1613 B.n222 B.n158 71.676
R1614 B.n218 B.n157 71.676
R1615 B.n214 B.n156 71.676
R1616 B.n209 B.n155 71.676
R1617 B.n205 B.n154 71.676
R1618 B.n201 B.n153 71.676
R1619 B.n197 B.n152 71.676
R1620 B.n193 B.n151 71.676
R1621 B.n189 B.n150 71.676
R1622 B.n185 B.n149 71.676
R1623 B.n181 B.n148 71.676
R1624 B.n177 B.n147 71.676
R1625 B.n449 B.n422 71.676
R1626 B.n455 B.n454 71.676
R1627 B.n458 B.n457 71.676
R1628 B.n463 B.n462 71.676
R1629 B.n466 B.n465 71.676
R1630 B.n471 B.n470 71.676
R1631 B.n474 B.n473 71.676
R1632 B.n479 B.n478 71.676
R1633 B.n482 B.n481 71.676
R1634 B.n488 B.n487 71.676
R1635 B.n491 B.n490 71.676
R1636 B.n496 B.n495 71.676
R1637 B.n499 B.n498 71.676
R1638 B.n507 B.n506 71.676
R1639 B.n510 B.n509 71.676
R1640 B.n515 B.n514 71.676
R1641 B.n518 B.n517 71.676
R1642 B.n523 B.n522 71.676
R1643 B.n526 B.n525 71.676
R1644 B.n531 B.n530 71.676
R1645 B.n534 B.n533 71.676
R1646 B.n539 B.n538 71.676
R1647 B.n542 B.n541 71.676
R1648 B.n450 B.n449 71.676
R1649 B.n456 B.n455 71.676
R1650 B.n457 B.n446 71.676
R1651 B.n464 B.n463 71.676
R1652 B.n465 B.n444 71.676
R1653 B.n472 B.n471 71.676
R1654 B.n473 B.n442 71.676
R1655 B.n480 B.n479 71.676
R1656 B.n481 B.n438 71.676
R1657 B.n489 B.n488 71.676
R1658 B.n490 B.n436 71.676
R1659 B.n497 B.n496 71.676
R1660 B.n498 B.n434 71.676
R1661 B.n508 B.n507 71.676
R1662 B.n509 B.n432 71.676
R1663 B.n516 B.n515 71.676
R1664 B.n517 B.n430 71.676
R1665 B.n524 B.n523 71.676
R1666 B.n525 B.n428 71.676
R1667 B.n532 B.n531 71.676
R1668 B.n533 B.n426 71.676
R1669 B.n540 B.n539 71.676
R1670 B.n541 B.n424 71.676
R1671 B.n1056 B.n1055 71.676
R1672 B.n1056 B.n2 71.676
R1673 B.n764 B.t1 69.0743
R1674 B.n1037 B.t7 69.0743
R1675 B.n728 B.t9 66.7718
R1676 B.n1013 B.t0 66.7718
R1677 B.n692 B.t4 64.4694
R1678 B.n989 B.t6 64.4694
R1679 B.n656 B.t5 62.1669
R1680 B.n965 B.t2 62.1669
R1681 B.n620 B.t3 59.8644
R1682 B.n941 B.t8 59.8644
R1683 B.n212 B.n175 59.5399
R1684 B.n173 B.n172 59.5399
R1685 B.n504 B.n503 59.5399
R1686 B.n485 B.n440 59.5399
R1687 B.n571 B.t11 41.4448
R1688 B.n131 B.t15 41.4448
R1689 B.n578 B.t11 36.8399
R1690 B.n915 B.t15 36.8399
R1691 B.n549 B.n421 32.3127
R1692 B.n545 B.n544 32.3127
R1693 B.n890 B.n889 32.3127
R1694 B.n895 B.n144 32.3127
R1695 B.t3 B.n372 18.4202
R1696 B.t8 B.n100 18.4202
R1697 B B.n1057 18.0485
R1698 B.t5 B.n348 16.1177
R1699 B.t2 B.n79 16.1177
R1700 B.t4 B.n324 13.8153
R1701 B.t6 B.n58 13.8153
R1702 B.t9 B.n300 11.5128
R1703 B.t0 B.n37 11.5128
R1704 B.n550 B.n549 10.6151
R1705 B.n551 B.n550 10.6151
R1706 B.n551 B.n413 10.6151
R1707 B.n561 B.n413 10.6151
R1708 B.n562 B.n561 10.6151
R1709 B.n563 B.n562 10.6151
R1710 B.n563 B.n405 10.6151
R1711 B.n574 B.n405 10.6151
R1712 B.n575 B.n574 10.6151
R1713 B.n576 B.n575 10.6151
R1714 B.n576 B.n398 10.6151
R1715 B.n586 B.n398 10.6151
R1716 B.n587 B.n586 10.6151
R1717 B.n588 B.n587 10.6151
R1718 B.n588 B.n390 10.6151
R1719 B.n598 B.n390 10.6151
R1720 B.n599 B.n598 10.6151
R1721 B.n600 B.n599 10.6151
R1722 B.n600 B.n382 10.6151
R1723 B.n610 B.n382 10.6151
R1724 B.n611 B.n610 10.6151
R1725 B.n612 B.n611 10.6151
R1726 B.n612 B.n374 10.6151
R1727 B.n622 B.n374 10.6151
R1728 B.n623 B.n622 10.6151
R1729 B.n624 B.n623 10.6151
R1730 B.n624 B.n366 10.6151
R1731 B.n634 B.n366 10.6151
R1732 B.n635 B.n634 10.6151
R1733 B.n636 B.n635 10.6151
R1734 B.n636 B.n358 10.6151
R1735 B.n646 B.n358 10.6151
R1736 B.n647 B.n646 10.6151
R1737 B.n648 B.n647 10.6151
R1738 B.n648 B.n350 10.6151
R1739 B.n658 B.n350 10.6151
R1740 B.n659 B.n658 10.6151
R1741 B.n660 B.n659 10.6151
R1742 B.n660 B.n342 10.6151
R1743 B.n670 B.n342 10.6151
R1744 B.n671 B.n670 10.6151
R1745 B.n672 B.n671 10.6151
R1746 B.n672 B.n334 10.6151
R1747 B.n682 B.n334 10.6151
R1748 B.n683 B.n682 10.6151
R1749 B.n684 B.n683 10.6151
R1750 B.n684 B.n326 10.6151
R1751 B.n694 B.n326 10.6151
R1752 B.n695 B.n694 10.6151
R1753 B.n696 B.n695 10.6151
R1754 B.n696 B.n318 10.6151
R1755 B.n706 B.n318 10.6151
R1756 B.n707 B.n706 10.6151
R1757 B.n708 B.n707 10.6151
R1758 B.n708 B.n310 10.6151
R1759 B.n718 B.n310 10.6151
R1760 B.n719 B.n718 10.6151
R1761 B.n720 B.n719 10.6151
R1762 B.n720 B.n302 10.6151
R1763 B.n730 B.n302 10.6151
R1764 B.n731 B.n730 10.6151
R1765 B.n732 B.n731 10.6151
R1766 B.n732 B.n294 10.6151
R1767 B.n742 B.n294 10.6151
R1768 B.n743 B.n742 10.6151
R1769 B.n744 B.n743 10.6151
R1770 B.n744 B.n286 10.6151
R1771 B.n754 B.n286 10.6151
R1772 B.n755 B.n754 10.6151
R1773 B.n756 B.n755 10.6151
R1774 B.n756 B.n278 10.6151
R1775 B.n766 B.n278 10.6151
R1776 B.n767 B.n766 10.6151
R1777 B.n768 B.n767 10.6151
R1778 B.n768 B.n270 10.6151
R1779 B.n779 B.n270 10.6151
R1780 B.n780 B.n779 10.6151
R1781 B.n781 B.n780 10.6151
R1782 B.n781 B.n0 10.6151
R1783 B.n451 B.n421 10.6151
R1784 B.n452 B.n451 10.6151
R1785 B.n453 B.n452 10.6151
R1786 B.n453 B.n447 10.6151
R1787 B.n459 B.n447 10.6151
R1788 B.n460 B.n459 10.6151
R1789 B.n461 B.n460 10.6151
R1790 B.n461 B.n445 10.6151
R1791 B.n467 B.n445 10.6151
R1792 B.n468 B.n467 10.6151
R1793 B.n469 B.n468 10.6151
R1794 B.n469 B.n443 10.6151
R1795 B.n475 B.n443 10.6151
R1796 B.n476 B.n475 10.6151
R1797 B.n477 B.n476 10.6151
R1798 B.n477 B.n441 10.6151
R1799 B.n483 B.n441 10.6151
R1800 B.n484 B.n483 10.6151
R1801 B.n486 B.n437 10.6151
R1802 B.n492 B.n437 10.6151
R1803 B.n493 B.n492 10.6151
R1804 B.n494 B.n493 10.6151
R1805 B.n494 B.n435 10.6151
R1806 B.n500 B.n435 10.6151
R1807 B.n501 B.n500 10.6151
R1808 B.n505 B.n501 10.6151
R1809 B.n511 B.n433 10.6151
R1810 B.n512 B.n511 10.6151
R1811 B.n513 B.n512 10.6151
R1812 B.n513 B.n431 10.6151
R1813 B.n519 B.n431 10.6151
R1814 B.n520 B.n519 10.6151
R1815 B.n521 B.n520 10.6151
R1816 B.n521 B.n429 10.6151
R1817 B.n527 B.n429 10.6151
R1818 B.n528 B.n527 10.6151
R1819 B.n529 B.n528 10.6151
R1820 B.n529 B.n427 10.6151
R1821 B.n535 B.n427 10.6151
R1822 B.n536 B.n535 10.6151
R1823 B.n537 B.n536 10.6151
R1824 B.n537 B.n425 10.6151
R1825 B.n543 B.n425 10.6151
R1826 B.n544 B.n543 10.6151
R1827 B.n545 B.n417 10.6151
R1828 B.n555 B.n417 10.6151
R1829 B.n556 B.n555 10.6151
R1830 B.n557 B.n556 10.6151
R1831 B.n557 B.n409 10.6151
R1832 B.n567 B.n409 10.6151
R1833 B.n568 B.n567 10.6151
R1834 B.n569 B.n568 10.6151
R1835 B.n569 B.n402 10.6151
R1836 B.n580 B.n402 10.6151
R1837 B.n581 B.n580 10.6151
R1838 B.n582 B.n581 10.6151
R1839 B.n582 B.n394 10.6151
R1840 B.n592 B.n394 10.6151
R1841 B.n593 B.n592 10.6151
R1842 B.n594 B.n593 10.6151
R1843 B.n594 B.n386 10.6151
R1844 B.n604 B.n386 10.6151
R1845 B.n605 B.n604 10.6151
R1846 B.n606 B.n605 10.6151
R1847 B.n606 B.n378 10.6151
R1848 B.n616 B.n378 10.6151
R1849 B.n617 B.n616 10.6151
R1850 B.n618 B.n617 10.6151
R1851 B.n618 B.n370 10.6151
R1852 B.n628 B.n370 10.6151
R1853 B.n629 B.n628 10.6151
R1854 B.n630 B.n629 10.6151
R1855 B.n630 B.n362 10.6151
R1856 B.n640 B.n362 10.6151
R1857 B.n641 B.n640 10.6151
R1858 B.n642 B.n641 10.6151
R1859 B.n642 B.n354 10.6151
R1860 B.n652 B.n354 10.6151
R1861 B.n653 B.n652 10.6151
R1862 B.n654 B.n653 10.6151
R1863 B.n654 B.n346 10.6151
R1864 B.n664 B.n346 10.6151
R1865 B.n665 B.n664 10.6151
R1866 B.n666 B.n665 10.6151
R1867 B.n666 B.n338 10.6151
R1868 B.n676 B.n338 10.6151
R1869 B.n677 B.n676 10.6151
R1870 B.n678 B.n677 10.6151
R1871 B.n678 B.n330 10.6151
R1872 B.n688 B.n330 10.6151
R1873 B.n689 B.n688 10.6151
R1874 B.n690 B.n689 10.6151
R1875 B.n690 B.n322 10.6151
R1876 B.n700 B.n322 10.6151
R1877 B.n701 B.n700 10.6151
R1878 B.n702 B.n701 10.6151
R1879 B.n702 B.n314 10.6151
R1880 B.n712 B.n314 10.6151
R1881 B.n713 B.n712 10.6151
R1882 B.n714 B.n713 10.6151
R1883 B.n714 B.n306 10.6151
R1884 B.n724 B.n306 10.6151
R1885 B.n725 B.n724 10.6151
R1886 B.n726 B.n725 10.6151
R1887 B.n726 B.n298 10.6151
R1888 B.n736 B.n298 10.6151
R1889 B.n737 B.n736 10.6151
R1890 B.n738 B.n737 10.6151
R1891 B.n738 B.n290 10.6151
R1892 B.n748 B.n290 10.6151
R1893 B.n749 B.n748 10.6151
R1894 B.n750 B.n749 10.6151
R1895 B.n750 B.n282 10.6151
R1896 B.n760 B.n282 10.6151
R1897 B.n761 B.n760 10.6151
R1898 B.n762 B.n761 10.6151
R1899 B.n762 B.n274 10.6151
R1900 B.n772 B.n274 10.6151
R1901 B.n773 B.n772 10.6151
R1902 B.n775 B.n773 10.6151
R1903 B.n775 B.n774 10.6151
R1904 B.n774 B.n266 10.6151
R1905 B.n786 B.n266 10.6151
R1906 B.n787 B.n786 10.6151
R1907 B.n788 B.n787 10.6151
R1908 B.n789 B.n788 10.6151
R1909 B.n790 B.n789 10.6151
R1910 B.n793 B.n790 10.6151
R1911 B.n794 B.n793 10.6151
R1912 B.n795 B.n794 10.6151
R1913 B.n796 B.n795 10.6151
R1914 B.n798 B.n796 10.6151
R1915 B.n799 B.n798 10.6151
R1916 B.n800 B.n799 10.6151
R1917 B.n801 B.n800 10.6151
R1918 B.n803 B.n801 10.6151
R1919 B.n804 B.n803 10.6151
R1920 B.n805 B.n804 10.6151
R1921 B.n806 B.n805 10.6151
R1922 B.n808 B.n806 10.6151
R1923 B.n809 B.n808 10.6151
R1924 B.n810 B.n809 10.6151
R1925 B.n811 B.n810 10.6151
R1926 B.n813 B.n811 10.6151
R1927 B.n814 B.n813 10.6151
R1928 B.n815 B.n814 10.6151
R1929 B.n816 B.n815 10.6151
R1930 B.n818 B.n816 10.6151
R1931 B.n819 B.n818 10.6151
R1932 B.n820 B.n819 10.6151
R1933 B.n821 B.n820 10.6151
R1934 B.n823 B.n821 10.6151
R1935 B.n824 B.n823 10.6151
R1936 B.n825 B.n824 10.6151
R1937 B.n826 B.n825 10.6151
R1938 B.n828 B.n826 10.6151
R1939 B.n829 B.n828 10.6151
R1940 B.n830 B.n829 10.6151
R1941 B.n831 B.n830 10.6151
R1942 B.n833 B.n831 10.6151
R1943 B.n834 B.n833 10.6151
R1944 B.n835 B.n834 10.6151
R1945 B.n836 B.n835 10.6151
R1946 B.n838 B.n836 10.6151
R1947 B.n839 B.n838 10.6151
R1948 B.n840 B.n839 10.6151
R1949 B.n841 B.n840 10.6151
R1950 B.n843 B.n841 10.6151
R1951 B.n844 B.n843 10.6151
R1952 B.n845 B.n844 10.6151
R1953 B.n846 B.n845 10.6151
R1954 B.n848 B.n846 10.6151
R1955 B.n849 B.n848 10.6151
R1956 B.n850 B.n849 10.6151
R1957 B.n851 B.n850 10.6151
R1958 B.n853 B.n851 10.6151
R1959 B.n854 B.n853 10.6151
R1960 B.n855 B.n854 10.6151
R1961 B.n856 B.n855 10.6151
R1962 B.n858 B.n856 10.6151
R1963 B.n859 B.n858 10.6151
R1964 B.n860 B.n859 10.6151
R1965 B.n861 B.n860 10.6151
R1966 B.n863 B.n861 10.6151
R1967 B.n864 B.n863 10.6151
R1968 B.n865 B.n864 10.6151
R1969 B.n866 B.n865 10.6151
R1970 B.n868 B.n866 10.6151
R1971 B.n869 B.n868 10.6151
R1972 B.n870 B.n869 10.6151
R1973 B.n871 B.n870 10.6151
R1974 B.n873 B.n871 10.6151
R1975 B.n874 B.n873 10.6151
R1976 B.n875 B.n874 10.6151
R1977 B.n876 B.n875 10.6151
R1978 B.n878 B.n876 10.6151
R1979 B.n879 B.n878 10.6151
R1980 B.n880 B.n879 10.6151
R1981 B.n881 B.n880 10.6151
R1982 B.n883 B.n881 10.6151
R1983 B.n884 B.n883 10.6151
R1984 B.n885 B.n884 10.6151
R1985 B.n886 B.n885 10.6151
R1986 B.n888 B.n886 10.6151
R1987 B.n889 B.n888 10.6151
R1988 B.n1049 B.n1 10.6151
R1989 B.n1049 B.n1048 10.6151
R1990 B.n1048 B.n1047 10.6151
R1991 B.n1047 B.n10 10.6151
R1992 B.n1041 B.n10 10.6151
R1993 B.n1041 B.n1040 10.6151
R1994 B.n1040 B.n1039 10.6151
R1995 B.n1039 B.n18 10.6151
R1996 B.n1033 B.n18 10.6151
R1997 B.n1033 B.n1032 10.6151
R1998 B.n1032 B.n1031 10.6151
R1999 B.n1031 B.n25 10.6151
R2000 B.n1025 B.n25 10.6151
R2001 B.n1025 B.n1024 10.6151
R2002 B.n1024 B.n1023 10.6151
R2003 B.n1023 B.n32 10.6151
R2004 B.n1017 B.n32 10.6151
R2005 B.n1017 B.n1016 10.6151
R2006 B.n1016 B.n1015 10.6151
R2007 B.n1015 B.n39 10.6151
R2008 B.n1009 B.n39 10.6151
R2009 B.n1009 B.n1008 10.6151
R2010 B.n1008 B.n1007 10.6151
R2011 B.n1007 B.n46 10.6151
R2012 B.n1001 B.n46 10.6151
R2013 B.n1001 B.n1000 10.6151
R2014 B.n1000 B.n999 10.6151
R2015 B.n999 B.n53 10.6151
R2016 B.n993 B.n53 10.6151
R2017 B.n993 B.n992 10.6151
R2018 B.n992 B.n991 10.6151
R2019 B.n991 B.n60 10.6151
R2020 B.n985 B.n60 10.6151
R2021 B.n985 B.n984 10.6151
R2022 B.n984 B.n983 10.6151
R2023 B.n983 B.n67 10.6151
R2024 B.n977 B.n67 10.6151
R2025 B.n977 B.n976 10.6151
R2026 B.n976 B.n975 10.6151
R2027 B.n975 B.n74 10.6151
R2028 B.n969 B.n74 10.6151
R2029 B.n969 B.n968 10.6151
R2030 B.n968 B.n967 10.6151
R2031 B.n967 B.n81 10.6151
R2032 B.n961 B.n81 10.6151
R2033 B.n961 B.n960 10.6151
R2034 B.n960 B.n959 10.6151
R2035 B.n959 B.n88 10.6151
R2036 B.n953 B.n88 10.6151
R2037 B.n953 B.n952 10.6151
R2038 B.n952 B.n951 10.6151
R2039 B.n951 B.n95 10.6151
R2040 B.n945 B.n95 10.6151
R2041 B.n945 B.n944 10.6151
R2042 B.n944 B.n943 10.6151
R2043 B.n943 B.n102 10.6151
R2044 B.n937 B.n102 10.6151
R2045 B.n937 B.n936 10.6151
R2046 B.n936 B.n935 10.6151
R2047 B.n935 B.n109 10.6151
R2048 B.n929 B.n109 10.6151
R2049 B.n929 B.n928 10.6151
R2050 B.n928 B.n927 10.6151
R2051 B.n927 B.n116 10.6151
R2052 B.n921 B.n116 10.6151
R2053 B.n921 B.n920 10.6151
R2054 B.n920 B.n919 10.6151
R2055 B.n919 B.n123 10.6151
R2056 B.n913 B.n123 10.6151
R2057 B.n913 B.n912 10.6151
R2058 B.n912 B.n911 10.6151
R2059 B.n911 B.n129 10.6151
R2060 B.n905 B.n129 10.6151
R2061 B.n905 B.n904 10.6151
R2062 B.n904 B.n903 10.6151
R2063 B.n903 B.n137 10.6151
R2064 B.n897 B.n137 10.6151
R2065 B.n897 B.n896 10.6151
R2066 B.n896 B.n895 10.6151
R2067 B.n176 B.n144 10.6151
R2068 B.n179 B.n176 10.6151
R2069 B.n180 B.n179 10.6151
R2070 B.n183 B.n180 10.6151
R2071 B.n184 B.n183 10.6151
R2072 B.n187 B.n184 10.6151
R2073 B.n188 B.n187 10.6151
R2074 B.n191 B.n188 10.6151
R2075 B.n192 B.n191 10.6151
R2076 B.n195 B.n192 10.6151
R2077 B.n196 B.n195 10.6151
R2078 B.n199 B.n196 10.6151
R2079 B.n200 B.n199 10.6151
R2080 B.n203 B.n200 10.6151
R2081 B.n204 B.n203 10.6151
R2082 B.n207 B.n204 10.6151
R2083 B.n208 B.n207 10.6151
R2084 B.n211 B.n208 10.6151
R2085 B.n216 B.n213 10.6151
R2086 B.n217 B.n216 10.6151
R2087 B.n220 B.n217 10.6151
R2088 B.n221 B.n220 10.6151
R2089 B.n224 B.n221 10.6151
R2090 B.n225 B.n224 10.6151
R2091 B.n228 B.n225 10.6151
R2092 B.n229 B.n228 10.6151
R2093 B.n233 B.n232 10.6151
R2094 B.n236 B.n233 10.6151
R2095 B.n237 B.n236 10.6151
R2096 B.n240 B.n237 10.6151
R2097 B.n241 B.n240 10.6151
R2098 B.n244 B.n241 10.6151
R2099 B.n245 B.n244 10.6151
R2100 B.n248 B.n245 10.6151
R2101 B.n249 B.n248 10.6151
R2102 B.n252 B.n249 10.6151
R2103 B.n253 B.n252 10.6151
R2104 B.n256 B.n253 10.6151
R2105 B.n257 B.n256 10.6151
R2106 B.n260 B.n257 10.6151
R2107 B.n261 B.n260 10.6151
R2108 B.n264 B.n261 10.6151
R2109 B.n265 B.n264 10.6151
R2110 B.n890 B.n265 10.6151
R2111 B.t1 B.n276 9.21034
R2112 B.t7 B.n16 9.21034
R2113 B.n1057 B.n0 8.11757
R2114 B.n1057 B.n1 8.11757
R2115 B.n486 B.n485 6.5566
R2116 B.n505 B.n504 6.5566
R2117 B.n213 B.n212 6.5566
R2118 B.n229 B.n173 6.5566
R2119 B.n485 B.n484 4.05904
R2120 B.n504 B.n433 4.05904
R2121 B.n212 B.n211 4.05904
R2122 B.n232 B.n173 4.05904
R2123 VN.n105 VN.n54 161.3
R2124 VN.n104 VN.n103 161.3
R2125 VN.n102 VN.n55 161.3
R2126 VN.n101 VN.n100 161.3
R2127 VN.n99 VN.n56 161.3
R2128 VN.n98 VN.n97 161.3
R2129 VN.n96 VN.n57 161.3
R2130 VN.n95 VN.n94 161.3
R2131 VN.n92 VN.n58 161.3
R2132 VN.n91 VN.n90 161.3
R2133 VN.n89 VN.n59 161.3
R2134 VN.n88 VN.n87 161.3
R2135 VN.n86 VN.n60 161.3
R2136 VN.n85 VN.n84 161.3
R2137 VN.n83 VN.n61 161.3
R2138 VN.n82 VN.n81 161.3
R2139 VN.n79 VN.n62 161.3
R2140 VN.n78 VN.n77 161.3
R2141 VN.n76 VN.n63 161.3
R2142 VN.n75 VN.n74 161.3
R2143 VN.n73 VN.n64 161.3
R2144 VN.n72 VN.n71 161.3
R2145 VN.n70 VN.n65 161.3
R2146 VN.n69 VN.n68 161.3
R2147 VN.n51 VN.n0 161.3
R2148 VN.n50 VN.n49 161.3
R2149 VN.n48 VN.n1 161.3
R2150 VN.n47 VN.n46 161.3
R2151 VN.n45 VN.n2 161.3
R2152 VN.n44 VN.n43 161.3
R2153 VN.n42 VN.n3 161.3
R2154 VN.n41 VN.n40 161.3
R2155 VN.n38 VN.n4 161.3
R2156 VN.n37 VN.n36 161.3
R2157 VN.n35 VN.n5 161.3
R2158 VN.n34 VN.n33 161.3
R2159 VN.n32 VN.n6 161.3
R2160 VN.n31 VN.n30 161.3
R2161 VN.n29 VN.n7 161.3
R2162 VN.n28 VN.n27 161.3
R2163 VN.n25 VN.n8 161.3
R2164 VN.n24 VN.n23 161.3
R2165 VN.n22 VN.n9 161.3
R2166 VN.n21 VN.n20 161.3
R2167 VN.n19 VN.n10 161.3
R2168 VN.n18 VN.n17 161.3
R2169 VN.n16 VN.n11 161.3
R2170 VN.n15 VN.n14 161.3
R2171 VN.n53 VN.n52 61.2309
R2172 VN.n107 VN.n106 61.2309
R2173 VN.n12 VN.t0 59.797
R2174 VN.n66 VN.t5 59.797
R2175 VN.n13 VN.n12 58.5323
R2176 VN.n67 VN.n66 58.5323
R2177 VN.n20 VN.n19 56.5617
R2178 VN.n33 VN.n32 56.5617
R2179 VN.n74 VN.n73 56.5617
R2180 VN.n87 VN.n86 56.5617
R2181 VN VN.n107 53.8112
R2182 VN.n46 VN.n45 51.7179
R2183 VN.n100 VN.n99 51.7179
R2184 VN.n46 VN.n1 29.4362
R2185 VN.n100 VN.n55 29.4362
R2186 VN.n13 VN.t8 27.4335
R2187 VN.n26 VN.t3 27.4335
R2188 VN.n39 VN.t6 27.4335
R2189 VN.n52 VN.t9 27.4335
R2190 VN.n67 VN.t2 27.4335
R2191 VN.n80 VN.t1 27.4335
R2192 VN.n93 VN.t7 27.4335
R2193 VN.n106 VN.t4 27.4335
R2194 VN.n14 VN.n11 24.5923
R2195 VN.n18 VN.n11 24.5923
R2196 VN.n19 VN.n18 24.5923
R2197 VN.n20 VN.n9 24.5923
R2198 VN.n24 VN.n9 24.5923
R2199 VN.n25 VN.n24 24.5923
R2200 VN.n27 VN.n7 24.5923
R2201 VN.n31 VN.n7 24.5923
R2202 VN.n32 VN.n31 24.5923
R2203 VN.n33 VN.n5 24.5923
R2204 VN.n37 VN.n5 24.5923
R2205 VN.n38 VN.n37 24.5923
R2206 VN.n40 VN.n3 24.5923
R2207 VN.n44 VN.n3 24.5923
R2208 VN.n45 VN.n44 24.5923
R2209 VN.n50 VN.n1 24.5923
R2210 VN.n51 VN.n50 24.5923
R2211 VN.n73 VN.n72 24.5923
R2212 VN.n72 VN.n65 24.5923
R2213 VN.n68 VN.n65 24.5923
R2214 VN.n86 VN.n85 24.5923
R2215 VN.n85 VN.n61 24.5923
R2216 VN.n81 VN.n61 24.5923
R2217 VN.n79 VN.n78 24.5923
R2218 VN.n78 VN.n63 24.5923
R2219 VN.n74 VN.n63 24.5923
R2220 VN.n99 VN.n98 24.5923
R2221 VN.n98 VN.n57 24.5923
R2222 VN.n94 VN.n57 24.5923
R2223 VN.n92 VN.n91 24.5923
R2224 VN.n91 VN.n59 24.5923
R2225 VN.n87 VN.n59 24.5923
R2226 VN.n105 VN.n104 24.5923
R2227 VN.n104 VN.n55 24.5923
R2228 VN.n52 VN.n51 21.1495
R2229 VN.n106 VN.n105 21.1495
R2230 VN.n14 VN.n13 16.7229
R2231 VN.n39 VN.n38 16.7229
R2232 VN.n68 VN.n67 16.7229
R2233 VN.n93 VN.n92 16.7229
R2234 VN.n26 VN.n25 12.2964
R2235 VN.n27 VN.n26 12.2964
R2236 VN.n81 VN.n80 12.2964
R2237 VN.n80 VN.n79 12.2964
R2238 VN.n40 VN.n39 7.86989
R2239 VN.n94 VN.n93 7.86989
R2240 VN.n69 VN.n66 2.63944
R2241 VN.n15 VN.n12 2.63944
R2242 VN.n107 VN.n54 0.417304
R2243 VN.n53 VN.n0 0.417304
R2244 VN VN.n53 0.394524
R2245 VN.n103 VN.n54 0.189894
R2246 VN.n103 VN.n102 0.189894
R2247 VN.n102 VN.n101 0.189894
R2248 VN.n101 VN.n56 0.189894
R2249 VN.n97 VN.n56 0.189894
R2250 VN.n97 VN.n96 0.189894
R2251 VN.n96 VN.n95 0.189894
R2252 VN.n95 VN.n58 0.189894
R2253 VN.n90 VN.n58 0.189894
R2254 VN.n90 VN.n89 0.189894
R2255 VN.n89 VN.n88 0.189894
R2256 VN.n88 VN.n60 0.189894
R2257 VN.n84 VN.n60 0.189894
R2258 VN.n84 VN.n83 0.189894
R2259 VN.n83 VN.n82 0.189894
R2260 VN.n82 VN.n62 0.189894
R2261 VN.n77 VN.n62 0.189894
R2262 VN.n77 VN.n76 0.189894
R2263 VN.n76 VN.n75 0.189894
R2264 VN.n75 VN.n64 0.189894
R2265 VN.n71 VN.n64 0.189894
R2266 VN.n71 VN.n70 0.189894
R2267 VN.n70 VN.n69 0.189894
R2268 VN.n16 VN.n15 0.189894
R2269 VN.n17 VN.n16 0.189894
R2270 VN.n17 VN.n10 0.189894
R2271 VN.n21 VN.n10 0.189894
R2272 VN.n22 VN.n21 0.189894
R2273 VN.n23 VN.n22 0.189894
R2274 VN.n23 VN.n8 0.189894
R2275 VN.n28 VN.n8 0.189894
R2276 VN.n29 VN.n28 0.189894
R2277 VN.n30 VN.n29 0.189894
R2278 VN.n30 VN.n6 0.189894
R2279 VN.n34 VN.n6 0.189894
R2280 VN.n35 VN.n34 0.189894
R2281 VN.n36 VN.n35 0.189894
R2282 VN.n36 VN.n4 0.189894
R2283 VN.n41 VN.n4 0.189894
R2284 VN.n42 VN.n41 0.189894
R2285 VN.n43 VN.n42 0.189894
R2286 VN.n43 VN.n2 0.189894
R2287 VN.n47 VN.n2 0.189894
R2288 VN.n48 VN.n47 0.189894
R2289 VN.n49 VN.n48 0.189894
R2290 VN.n49 VN.n0 0.189894
R2291 VDD2.n1 VDD2.t9 81.6218
R2292 VDD2.n4 VDD2.t5 78.0961
R2293 VDD2.n3 VDD2.n2 76.0588
R2294 VDD2 VDD2.n7 76.056
R2295 VDD2.n6 VDD2.n5 73.47
R2296 VDD2.n1 VDD2.n0 73.4697
R2297 VDD2.n4 VDD2.n3 44.1528
R2298 VDD2.n7 VDD2.t7 4.62667
R2299 VDD2.n7 VDD2.t4 4.62667
R2300 VDD2.n5 VDD2.t2 4.62667
R2301 VDD2.n5 VDD2.t8 4.62667
R2302 VDD2.n2 VDD2.t3 4.62667
R2303 VDD2.n2 VDD2.t0 4.62667
R2304 VDD2.n0 VDD2.t1 4.62667
R2305 VDD2.n0 VDD2.t6 4.62667
R2306 VDD2.n6 VDD2.n4 3.52636
R2307 VDD2 VDD2.n6 0.940155
R2308 VDD2.n3 VDD2.n1 0.826619
C0 VN VDD2 4.40601f
C1 VDD1 VDD2 2.93014f
C2 VTAIL VDD2 8.03917f
C3 VN VP 8.68139f
C4 VDD1 VP 4.97789f
C5 VTAIL VP 6.25027f
C6 VP VDD2 0.736346f
C7 VN VDD1 0.160588f
C8 VN VTAIL 6.23597f
C9 VTAIL VDD1 7.9783f
C10 VDD2 B 7.29671f
C11 VDD1 B 7.195543f
C12 VTAIL B 5.323847f
C13 VN B 22.94935f
C14 VP B 21.418533f
C15 VDD2.t9 B 0.98001f
C16 VDD2.t1 B 0.094419f
C17 VDD2.t6 B 0.094419f
C18 VDD2.n0 B 0.750656f
C19 VDD2.n1 B 1.18639f
C20 VDD2.t3 B 0.094419f
C21 VDD2.t0 B 0.094419f
C22 VDD2.n2 B 0.777219f
C23 VDD2.n3 B 3.38298f
C24 VDD2.t5 B 0.954037f
C25 VDD2.n4 B 3.29459f
C26 VDD2.t2 B 0.094419f
C27 VDD2.t8 B 0.094419f
C28 VDD2.n5 B 0.750659f
C29 VDD2.n6 B 0.62047f
C30 VDD2.t7 B 0.094419f
C31 VDD2.t4 B 0.094419f
C32 VDD2.n7 B 0.777173f
C33 VN.n0 B 0.039966f
C34 VN.t9 B 0.883878f
C35 VN.n1 B 0.041974f
C36 VN.n2 B 0.021254f
C37 VN.n3 B 0.039413f
C38 VN.n4 B 0.021254f
C39 VN.t6 B 0.883878f
C40 VN.n5 B 0.039413f
C41 VN.n6 B 0.021254f
C42 VN.n7 B 0.039413f
C43 VN.n8 B 0.021254f
C44 VN.t3 B 0.883878f
C45 VN.n9 B 0.039413f
C46 VN.n10 B 0.021254f
C47 VN.n11 B 0.039413f
C48 VN.t0 B 1.15554f
C49 VN.n12 B 0.417457f
C50 VN.t8 B 0.883878f
C51 VN.n13 B 0.418034f
C52 VN.n14 B 0.033187f
C53 VN.n15 B 0.276547f
C54 VN.n16 B 0.021254f
C55 VN.n17 B 0.021254f
C56 VN.n18 B 0.039413f
C57 VN.n19 B 0.028249f
C58 VN.n20 B 0.033542f
C59 VN.n21 B 0.021254f
C60 VN.n22 B 0.021254f
C61 VN.n23 B 0.021254f
C62 VN.n24 B 0.039413f
C63 VN.n25 B 0.029684f
C64 VN.n26 B 0.338967f
C65 VN.n27 B 0.029684f
C66 VN.n28 B 0.021254f
C67 VN.n29 B 0.021254f
C68 VN.n30 B 0.021254f
C69 VN.n31 B 0.039413f
C70 VN.n32 B 0.033542f
C71 VN.n33 B 0.028249f
C72 VN.n34 B 0.021254f
C73 VN.n35 B 0.021254f
C74 VN.n36 B 0.021254f
C75 VN.n37 B 0.039413f
C76 VN.n38 B 0.033187f
C77 VN.n39 B 0.338967f
C78 VN.n40 B 0.026182f
C79 VN.n41 B 0.021254f
C80 VN.n42 B 0.021254f
C81 VN.n43 B 0.021254f
C82 VN.n44 B 0.039413f
C83 VN.n45 B 0.038188f
C84 VN.n46 B 0.021041f
C85 VN.n47 B 0.021254f
C86 VN.n48 B 0.021254f
C87 VN.n49 B 0.021254f
C88 VN.n50 B 0.039413f
C89 VN.n51 B 0.036689f
C90 VN.n52 B 0.428932f
C91 VN.n53 B 0.064691f
C92 VN.n54 B 0.039966f
C93 VN.t4 B 0.883878f
C94 VN.n55 B 0.041974f
C95 VN.n56 B 0.021254f
C96 VN.n57 B 0.039413f
C97 VN.n58 B 0.021254f
C98 VN.t7 B 0.883878f
C99 VN.n59 B 0.039413f
C100 VN.n60 B 0.021254f
C101 VN.n61 B 0.039413f
C102 VN.n62 B 0.021254f
C103 VN.t1 B 0.883878f
C104 VN.n63 B 0.039413f
C105 VN.n64 B 0.021254f
C106 VN.n65 B 0.039413f
C107 VN.t5 B 1.15554f
C108 VN.n66 B 0.417457f
C109 VN.t2 B 0.883878f
C110 VN.n67 B 0.418034f
C111 VN.n68 B 0.033187f
C112 VN.n69 B 0.276547f
C113 VN.n70 B 0.021254f
C114 VN.n71 B 0.021254f
C115 VN.n72 B 0.039413f
C116 VN.n73 B 0.028249f
C117 VN.n74 B 0.033542f
C118 VN.n75 B 0.021254f
C119 VN.n76 B 0.021254f
C120 VN.n77 B 0.021254f
C121 VN.n78 B 0.039413f
C122 VN.n79 B 0.029684f
C123 VN.n80 B 0.338967f
C124 VN.n81 B 0.029684f
C125 VN.n82 B 0.021254f
C126 VN.n83 B 0.021254f
C127 VN.n84 B 0.021254f
C128 VN.n85 B 0.039413f
C129 VN.n86 B 0.033542f
C130 VN.n87 B 0.028249f
C131 VN.n88 B 0.021254f
C132 VN.n89 B 0.021254f
C133 VN.n90 B 0.021254f
C134 VN.n91 B 0.039413f
C135 VN.n92 B 0.033187f
C136 VN.n93 B 0.338967f
C137 VN.n94 B 0.026182f
C138 VN.n95 B 0.021254f
C139 VN.n96 B 0.021254f
C140 VN.n97 B 0.021254f
C141 VN.n98 B 0.039413f
C142 VN.n99 B 0.038188f
C143 VN.n100 B 0.021041f
C144 VN.n101 B 0.021254f
C145 VN.n102 B 0.021254f
C146 VN.n103 B 0.021254f
C147 VN.n104 B 0.039413f
C148 VN.n105 B 0.036689f
C149 VN.n106 B 0.428932f
C150 VN.n107 B 1.36876f
C151 VDD1.t3 B 1.01163f
C152 VDD1.t6 B 0.097465f
C153 VDD1.t0 B 0.097465f
C154 VDD1.n0 B 0.774875f
C155 VDD1.n1 B 1.23439f
C156 VDD1.t9 B 1.01162f
C157 VDD1.t5 B 0.097465f
C158 VDD1.t8 B 0.097465f
C159 VDD1.n2 B 0.774872f
C160 VDD1.n3 B 1.22466f
C161 VDD1.t2 B 0.097465f
C162 VDD1.t7 B 0.097465f
C163 VDD1.n4 B 0.802292f
C164 VDD1.n5 B 3.66452f
C165 VDD1.t4 B 0.097465f
C166 VDD1.t1 B 0.097465f
C167 VDD1.n6 B 0.774871f
C168 VDD1.n7 B 3.51917f
C169 VTAIL.t7 B 0.110537f
C170 VTAIL.t0 B 0.110537f
C171 VTAIL.n0 B 0.805409f
C172 VTAIL.n1 B 0.80485f
C173 VTAIL.t12 B 1.03183f
C174 VTAIL.n2 B 0.966597f
C175 VTAIL.t19 B 0.110537f
C176 VTAIL.t10 B 0.110537f
C177 VTAIL.n3 B 0.805409f
C178 VTAIL.n4 B 1.02772f
C179 VTAIL.t18 B 0.110537f
C180 VTAIL.t11 B 0.110537f
C181 VTAIL.n5 B 0.805409f
C182 VTAIL.n6 B 2.23154f
C183 VTAIL.t3 B 0.110537f
C184 VTAIL.t5 B 0.110537f
C185 VTAIL.n7 B 0.805413f
C186 VTAIL.n8 B 2.23153f
C187 VTAIL.t4 B 0.110537f
C188 VTAIL.t9 B 0.110537f
C189 VTAIL.n9 B 0.805413f
C190 VTAIL.n10 B 1.02772f
C191 VTAIL.t1 B 1.03183f
C192 VTAIL.n11 B 0.966593f
C193 VTAIL.t15 B 0.110537f
C194 VTAIL.t16 B 0.110537f
C195 VTAIL.n12 B 0.805413f
C196 VTAIL.n13 B 0.891545f
C197 VTAIL.t14 B 0.110537f
C198 VTAIL.t13 B 0.110537f
C199 VTAIL.n14 B 0.805413f
C200 VTAIL.n15 B 1.02772f
C201 VTAIL.t17 B 1.03183f
C202 VTAIL.n16 B 1.93528f
C203 VTAIL.t8 B 1.03183f
C204 VTAIL.n17 B 1.93528f
C205 VTAIL.t6 B 0.110537f
C206 VTAIL.t2 B 0.110537f
C207 VTAIL.n18 B 0.805409f
C208 VTAIL.n19 B 0.743117f
C209 VP.n0 B 0.04148f
C210 VP.t2 B 0.917355f
C211 VP.n1 B 0.043564f
C212 VP.n2 B 0.022059f
C213 VP.n3 B 0.040906f
C214 VP.n4 B 0.022059f
C215 VP.t7 B 0.917355f
C216 VP.n5 B 0.040906f
C217 VP.n6 B 0.022059f
C218 VP.n7 B 0.040906f
C219 VP.n8 B 0.022059f
C220 VP.t1 B 0.917355f
C221 VP.n9 B 0.040906f
C222 VP.n10 B 0.022059f
C223 VP.n11 B 0.040906f
C224 VP.n12 B 0.022059f
C225 VP.t4 B 0.917355f
C226 VP.n13 B 0.040906f
C227 VP.n14 B 0.022059f
C228 VP.n15 B 0.040906f
C229 VP.n16 B 0.04148f
C230 VP.t8 B 0.917355f
C231 VP.n17 B 0.043564f
C232 VP.n18 B 0.022059f
C233 VP.n19 B 0.040906f
C234 VP.n20 B 0.022059f
C235 VP.t5 B 0.917355f
C236 VP.n21 B 0.040906f
C237 VP.n22 B 0.022059f
C238 VP.n23 B 0.040906f
C239 VP.n24 B 0.022059f
C240 VP.t9 B 0.917355f
C241 VP.n25 B 0.040906f
C242 VP.n26 B 0.022059f
C243 VP.n27 B 0.040906f
C244 VP.t6 B 1.19931f
C245 VP.n28 B 0.43327f
C246 VP.t3 B 0.917355f
C247 VP.n29 B 0.433868f
C248 VP.n30 B 0.034444f
C249 VP.n31 B 0.287022f
C250 VP.n32 B 0.022059f
C251 VP.n33 B 0.022059f
C252 VP.n34 B 0.040906f
C253 VP.n35 B 0.029319f
C254 VP.n36 B 0.034812f
C255 VP.n37 B 0.022059f
C256 VP.n38 B 0.022059f
C257 VP.n39 B 0.022059f
C258 VP.n40 B 0.040906f
C259 VP.n41 B 0.030809f
C260 VP.n42 B 0.351806f
C261 VP.n43 B 0.030809f
C262 VP.n44 B 0.022059f
C263 VP.n45 B 0.022059f
C264 VP.n46 B 0.022059f
C265 VP.n47 B 0.040906f
C266 VP.n48 B 0.034812f
C267 VP.n49 B 0.029319f
C268 VP.n50 B 0.022059f
C269 VP.n51 B 0.022059f
C270 VP.n52 B 0.022059f
C271 VP.n53 B 0.040906f
C272 VP.n54 B 0.034444f
C273 VP.n55 B 0.351806f
C274 VP.n56 B 0.027174f
C275 VP.n57 B 0.022059f
C276 VP.n58 B 0.022059f
C277 VP.n59 B 0.022059f
C278 VP.n60 B 0.040906f
C279 VP.n61 B 0.039635f
C280 VP.n62 B 0.021838f
C281 VP.n63 B 0.022059f
C282 VP.n64 B 0.022059f
C283 VP.n65 B 0.022059f
C284 VP.n66 B 0.040906f
C285 VP.n67 B 0.038078f
C286 VP.n68 B 0.445178f
C287 VP.n69 B 1.41513f
C288 VP.n70 B 1.42992f
C289 VP.t0 B 0.917355f
C290 VP.n71 B 0.445178f
C291 VP.n72 B 0.038078f
C292 VP.n73 B 0.04148f
C293 VP.n74 B 0.022059f
C294 VP.n75 B 0.022059f
C295 VP.n76 B 0.043564f
C296 VP.n77 B 0.021838f
C297 VP.n78 B 0.039635f
C298 VP.n79 B 0.022059f
C299 VP.n80 B 0.022059f
C300 VP.n81 B 0.022059f
C301 VP.n82 B 0.040906f
C302 VP.n83 B 0.027174f
C303 VP.n84 B 0.351806f
C304 VP.n85 B 0.034444f
C305 VP.n86 B 0.022059f
C306 VP.n87 B 0.022059f
C307 VP.n88 B 0.022059f
C308 VP.n89 B 0.040906f
C309 VP.n90 B 0.029319f
C310 VP.n91 B 0.034812f
C311 VP.n92 B 0.022059f
C312 VP.n93 B 0.022059f
C313 VP.n94 B 0.022059f
C314 VP.n95 B 0.040906f
C315 VP.n96 B 0.030809f
C316 VP.n97 B 0.351806f
C317 VP.n98 B 0.030809f
C318 VP.n99 B 0.022059f
C319 VP.n100 B 0.022059f
C320 VP.n101 B 0.022059f
C321 VP.n102 B 0.040906f
C322 VP.n103 B 0.034812f
C323 VP.n104 B 0.029319f
C324 VP.n105 B 0.022059f
C325 VP.n106 B 0.022059f
C326 VP.n107 B 0.022059f
C327 VP.n108 B 0.040906f
C328 VP.n109 B 0.034444f
C329 VP.n110 B 0.351806f
C330 VP.n111 B 0.027174f
C331 VP.n112 B 0.022059f
C332 VP.n113 B 0.022059f
C333 VP.n114 B 0.022059f
C334 VP.n115 B 0.040906f
C335 VP.n116 B 0.039635f
C336 VP.n117 B 0.021838f
C337 VP.n118 B 0.022059f
C338 VP.n119 B 0.022059f
C339 VP.n120 B 0.022059f
C340 VP.n121 B 0.040906f
C341 VP.n122 B 0.038078f
C342 VP.n123 B 0.445178f
C343 VP.n124 B 0.067141f
.ends

