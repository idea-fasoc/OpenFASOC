* NGSPICE file created from diff_pair_sample_0898.ext - technology: sky130A

.subckt diff_pair_sample_0898 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=1.17645 ps=7.46 w=7.13 l=0.96
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=0 ps=0 w=7.13 l=0.96
X2 VTAIL.t1 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=1.17645 ps=7.46 w=7.13 l=0.96
X3 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=1.17645 ps=7.46 w=7.13 l=0.96
X4 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=0 ps=0 w=7.13 l=0.96
X5 VTAIL.t2 VN.t2 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=1.17645 ps=7.46 w=7.13 l=0.96
X6 VDD1.t4 VP.t1 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=2.7807 ps=15.04 w=7.13 l=0.96
X7 VDD1.t5 VP.t2 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=1.17645 ps=7.46 w=7.13 l=0.96
X8 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=2.7807 ps=15.04 w=7.13 l=0.96
X9 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=2.7807 ps=15.04 w=7.13 l=0.96
X10 VTAIL.t7 VP.t3 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=1.17645 ps=7.46 w=7.13 l=0.96
X11 VDD1.t2 VP.t4 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.17645 pd=7.46 as=2.7807 ps=15.04 w=7.13 l=0.96
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=0 ps=0 w=7.13 l=0.96
X13 VDD1.t0 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=1.17645 ps=7.46 w=7.13 l=0.96
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=0 ps=0 w=7.13 l=0.96
X15 VDD2.t0 VN.t5 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7807 pd=15.04 as=1.17645 ps=7.46 w=7.13 l=0.96
R0 VP.n5 VP.t2 239.105
R1 VP.n12 VP.t5 220.165
R2 VP.n19 VP.t1 220.165
R3 VP.n9 VP.t4 220.165
R4 VP.n1 VP.t3 178.994
R5 VP.n4 VP.t0 178.994
R6 VP.n20 VP.n19 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n8 VP.n3 161.3
R9 VP.n10 VP.n9 161.3
R10 VP.n18 VP.n0 161.3
R11 VP.n17 VP.n16 161.3
R12 VP.n15 VP.n14 161.3
R13 VP.n13 VP.n2 161.3
R14 VP.n12 VP.n11 161.3
R15 VP.n14 VP.n13 50.6917
R16 VP.n18 VP.n17 50.6917
R17 VP.n8 VP.n7 50.6917
R18 VP.n6 VP.n5 43.2502
R19 VP.n5 VP.n4 42.2819
R20 VP.n11 VP.n10 38.6028
R21 VP.n14 VP.n1 12.234
R22 VP.n17 VP.n1 12.234
R23 VP.n7 VP.n4 12.234
R24 VP.n13 VP.n12 8.76414
R25 VP.n19 VP.n18 8.76414
R26 VP.n9 VP.n8 8.76414
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VDD1 VDD1.t5 70.2502
R36 VDD1.n1 VDD1.t0 70.1364
R37 VDD1.n1 VDD1.n0 66.8036
R38 VDD1.n3 VDD1.n2 66.5808
R39 VDD1.n3 VDD1.n1 34.6151
R40 VDD1.n2 VDD1.t1 2.7775
R41 VDD1.n2 VDD1.t2 2.7775
R42 VDD1.n0 VDD1.t3 2.7775
R43 VDD1.n0 VDD1.t4 2.7775
R44 VDD1 VDD1.n3 0.220328
R45 VTAIL.n7 VTAIL.t3 52.6791
R46 VTAIL.n10 VTAIL.t6 52.6789
R47 VTAIL.n11 VTAIL.t4 52.6789
R48 VTAIL.n2 VTAIL.t9 52.6789
R49 VTAIL.n9 VTAIL.n8 49.9021
R50 VTAIL.n6 VTAIL.n5 49.9021
R51 VTAIL.n1 VTAIL.n0 49.9021
R52 VTAIL.n4 VTAIL.n3 49.9021
R53 VTAIL.n6 VTAIL.n4 20.7376
R54 VTAIL.n11 VTAIL.n10 19.6255
R55 VTAIL.n0 VTAIL.t0 2.7775
R56 VTAIL.n0 VTAIL.t1 2.7775
R57 VTAIL.n3 VTAIL.t5 2.7775
R58 VTAIL.n3 VTAIL.t7 2.7775
R59 VTAIL.n8 VTAIL.t8 2.7775
R60 VTAIL.n8 VTAIL.t10 2.7775
R61 VTAIL.n5 VTAIL.t11 2.7775
R62 VTAIL.n5 VTAIL.t2 2.7775
R63 VTAIL.n7 VTAIL.n6 1.11257
R64 VTAIL.n10 VTAIL.n9 1.11257
R65 VTAIL.n4 VTAIL.n2 1.11257
R66 VTAIL.n9 VTAIL.n7 1.02636
R67 VTAIL.n2 VTAIL.n1 1.02636
R68 VTAIL VTAIL.n11 0.776362
R69 VTAIL VTAIL.n1 0.336707
R70 B.n515 B.n514 585
R71 B.n205 B.n77 585
R72 B.n204 B.n203 585
R73 B.n202 B.n201 585
R74 B.n200 B.n199 585
R75 B.n198 B.n197 585
R76 B.n196 B.n195 585
R77 B.n194 B.n193 585
R78 B.n192 B.n191 585
R79 B.n190 B.n189 585
R80 B.n188 B.n187 585
R81 B.n186 B.n185 585
R82 B.n184 B.n183 585
R83 B.n182 B.n181 585
R84 B.n180 B.n179 585
R85 B.n178 B.n177 585
R86 B.n176 B.n175 585
R87 B.n174 B.n173 585
R88 B.n172 B.n171 585
R89 B.n170 B.n169 585
R90 B.n168 B.n167 585
R91 B.n166 B.n165 585
R92 B.n164 B.n163 585
R93 B.n162 B.n161 585
R94 B.n160 B.n159 585
R95 B.n158 B.n157 585
R96 B.n156 B.n155 585
R97 B.n153 B.n152 585
R98 B.n151 B.n150 585
R99 B.n149 B.n148 585
R100 B.n147 B.n146 585
R101 B.n145 B.n144 585
R102 B.n143 B.n142 585
R103 B.n141 B.n140 585
R104 B.n139 B.n138 585
R105 B.n137 B.n136 585
R106 B.n135 B.n134 585
R107 B.n132 B.n131 585
R108 B.n130 B.n129 585
R109 B.n128 B.n127 585
R110 B.n126 B.n125 585
R111 B.n124 B.n123 585
R112 B.n122 B.n121 585
R113 B.n120 B.n119 585
R114 B.n118 B.n117 585
R115 B.n116 B.n115 585
R116 B.n114 B.n113 585
R117 B.n112 B.n111 585
R118 B.n110 B.n109 585
R119 B.n108 B.n107 585
R120 B.n106 B.n105 585
R121 B.n104 B.n103 585
R122 B.n102 B.n101 585
R123 B.n100 B.n99 585
R124 B.n98 B.n97 585
R125 B.n96 B.n95 585
R126 B.n94 B.n93 585
R127 B.n92 B.n91 585
R128 B.n90 B.n89 585
R129 B.n88 B.n87 585
R130 B.n86 B.n85 585
R131 B.n84 B.n83 585
R132 B.n46 B.n45 585
R133 B.n520 B.n519 585
R134 B.n513 B.n78 585
R135 B.n78 B.n43 585
R136 B.n512 B.n42 585
R137 B.n524 B.n42 585
R138 B.n511 B.n41 585
R139 B.n525 B.n41 585
R140 B.n510 B.n40 585
R141 B.n526 B.n40 585
R142 B.n509 B.n508 585
R143 B.n508 B.n36 585
R144 B.n507 B.n35 585
R145 B.n532 B.n35 585
R146 B.n506 B.n34 585
R147 B.n533 B.n34 585
R148 B.n505 B.n33 585
R149 B.n534 B.n33 585
R150 B.n504 B.n503 585
R151 B.n503 B.n29 585
R152 B.n502 B.n28 585
R153 B.n540 B.n28 585
R154 B.n501 B.n27 585
R155 B.n541 B.n27 585
R156 B.n500 B.n26 585
R157 B.n542 B.n26 585
R158 B.n499 B.n498 585
R159 B.n498 B.n25 585
R160 B.n497 B.n21 585
R161 B.n548 B.n21 585
R162 B.n496 B.n20 585
R163 B.n549 B.n20 585
R164 B.n495 B.n19 585
R165 B.n550 B.n19 585
R166 B.n494 B.n493 585
R167 B.n493 B.n18 585
R168 B.n492 B.n14 585
R169 B.n556 B.n14 585
R170 B.n491 B.n13 585
R171 B.n557 B.n13 585
R172 B.n490 B.n12 585
R173 B.n558 B.n12 585
R174 B.n489 B.n488 585
R175 B.n488 B.t0 585
R176 B.n487 B.n486 585
R177 B.n487 B.n8 585
R178 B.n485 B.n7 585
R179 B.n565 B.n7 585
R180 B.n484 B.n6 585
R181 B.n566 B.n6 585
R182 B.n483 B.n5 585
R183 B.n567 B.n5 585
R184 B.n482 B.n481 585
R185 B.n481 B.n4 585
R186 B.n480 B.n206 585
R187 B.n480 B.n479 585
R188 B.n470 B.n207 585
R189 B.t3 B.n207 585
R190 B.n472 B.n471 585
R191 B.n473 B.n472 585
R192 B.n469 B.n212 585
R193 B.n212 B.n211 585
R194 B.n468 B.n467 585
R195 B.n467 B.n466 585
R196 B.n214 B.n213 585
R197 B.n459 B.n214 585
R198 B.n458 B.n457 585
R199 B.n460 B.n458 585
R200 B.n456 B.n219 585
R201 B.n219 B.n218 585
R202 B.n455 B.n454 585
R203 B.n454 B.n453 585
R204 B.n221 B.n220 585
R205 B.n446 B.n221 585
R206 B.n445 B.n444 585
R207 B.n447 B.n445 585
R208 B.n443 B.n226 585
R209 B.n226 B.n225 585
R210 B.n442 B.n441 585
R211 B.n441 B.n440 585
R212 B.n228 B.n227 585
R213 B.n229 B.n228 585
R214 B.n433 B.n432 585
R215 B.n434 B.n433 585
R216 B.n431 B.n234 585
R217 B.n234 B.n233 585
R218 B.n430 B.n429 585
R219 B.n429 B.n428 585
R220 B.n236 B.n235 585
R221 B.n237 B.n236 585
R222 B.n421 B.n420 585
R223 B.n422 B.n421 585
R224 B.n419 B.n242 585
R225 B.n242 B.n241 585
R226 B.n418 B.n417 585
R227 B.n417 B.n416 585
R228 B.n244 B.n243 585
R229 B.n245 B.n244 585
R230 B.n412 B.n411 585
R231 B.n248 B.n247 585
R232 B.n408 B.n407 585
R233 B.n409 B.n408 585
R234 B.n406 B.n280 585
R235 B.n405 B.n404 585
R236 B.n403 B.n402 585
R237 B.n401 B.n400 585
R238 B.n399 B.n398 585
R239 B.n397 B.n396 585
R240 B.n395 B.n394 585
R241 B.n393 B.n392 585
R242 B.n391 B.n390 585
R243 B.n389 B.n388 585
R244 B.n387 B.n386 585
R245 B.n385 B.n384 585
R246 B.n383 B.n382 585
R247 B.n381 B.n380 585
R248 B.n379 B.n378 585
R249 B.n377 B.n376 585
R250 B.n375 B.n374 585
R251 B.n373 B.n372 585
R252 B.n371 B.n370 585
R253 B.n369 B.n368 585
R254 B.n367 B.n366 585
R255 B.n365 B.n364 585
R256 B.n363 B.n362 585
R257 B.n361 B.n360 585
R258 B.n359 B.n358 585
R259 B.n357 B.n356 585
R260 B.n355 B.n354 585
R261 B.n353 B.n352 585
R262 B.n351 B.n350 585
R263 B.n349 B.n348 585
R264 B.n347 B.n346 585
R265 B.n345 B.n344 585
R266 B.n343 B.n342 585
R267 B.n341 B.n340 585
R268 B.n339 B.n338 585
R269 B.n337 B.n336 585
R270 B.n335 B.n334 585
R271 B.n333 B.n332 585
R272 B.n331 B.n330 585
R273 B.n329 B.n328 585
R274 B.n327 B.n326 585
R275 B.n325 B.n324 585
R276 B.n323 B.n322 585
R277 B.n321 B.n320 585
R278 B.n319 B.n318 585
R279 B.n317 B.n316 585
R280 B.n315 B.n314 585
R281 B.n313 B.n312 585
R282 B.n311 B.n310 585
R283 B.n309 B.n308 585
R284 B.n307 B.n306 585
R285 B.n305 B.n304 585
R286 B.n303 B.n302 585
R287 B.n301 B.n300 585
R288 B.n299 B.n298 585
R289 B.n297 B.n296 585
R290 B.n295 B.n294 585
R291 B.n293 B.n292 585
R292 B.n291 B.n290 585
R293 B.n289 B.n288 585
R294 B.n287 B.n279 585
R295 B.n409 B.n279 585
R296 B.n413 B.n246 585
R297 B.n246 B.n245 585
R298 B.n415 B.n414 585
R299 B.n416 B.n415 585
R300 B.n240 B.n239 585
R301 B.n241 B.n240 585
R302 B.n424 B.n423 585
R303 B.n423 B.n422 585
R304 B.n425 B.n238 585
R305 B.n238 B.n237 585
R306 B.n427 B.n426 585
R307 B.n428 B.n427 585
R308 B.n232 B.n231 585
R309 B.n233 B.n232 585
R310 B.n436 B.n435 585
R311 B.n435 B.n434 585
R312 B.n437 B.n230 585
R313 B.n230 B.n229 585
R314 B.n439 B.n438 585
R315 B.n440 B.n439 585
R316 B.n224 B.n223 585
R317 B.n225 B.n224 585
R318 B.n449 B.n448 585
R319 B.n448 B.n447 585
R320 B.n450 B.n222 585
R321 B.n446 B.n222 585
R322 B.n452 B.n451 585
R323 B.n453 B.n452 585
R324 B.n217 B.n216 585
R325 B.n218 B.n217 585
R326 B.n462 B.n461 585
R327 B.n461 B.n460 585
R328 B.n463 B.n215 585
R329 B.n459 B.n215 585
R330 B.n465 B.n464 585
R331 B.n466 B.n465 585
R332 B.n210 B.n209 585
R333 B.n211 B.n210 585
R334 B.n475 B.n474 585
R335 B.n474 B.n473 585
R336 B.n476 B.n208 585
R337 B.n208 B.t3 585
R338 B.n478 B.n477 585
R339 B.n479 B.n478 585
R340 B.n3 B.n0 585
R341 B.n4 B.n3 585
R342 B.n564 B.n1 585
R343 B.n565 B.n564 585
R344 B.n563 B.n562 585
R345 B.n563 B.n8 585
R346 B.n561 B.n9 585
R347 B.t0 B.n9 585
R348 B.n560 B.n559 585
R349 B.n559 B.n558 585
R350 B.n11 B.n10 585
R351 B.n557 B.n11 585
R352 B.n555 B.n554 585
R353 B.n556 B.n555 585
R354 B.n553 B.n15 585
R355 B.n18 B.n15 585
R356 B.n552 B.n551 585
R357 B.n551 B.n550 585
R358 B.n17 B.n16 585
R359 B.n549 B.n17 585
R360 B.n547 B.n546 585
R361 B.n548 B.n547 585
R362 B.n545 B.n22 585
R363 B.n25 B.n22 585
R364 B.n544 B.n543 585
R365 B.n543 B.n542 585
R366 B.n24 B.n23 585
R367 B.n541 B.n24 585
R368 B.n539 B.n538 585
R369 B.n540 B.n539 585
R370 B.n537 B.n30 585
R371 B.n30 B.n29 585
R372 B.n536 B.n535 585
R373 B.n535 B.n534 585
R374 B.n32 B.n31 585
R375 B.n533 B.n32 585
R376 B.n531 B.n530 585
R377 B.n532 B.n531 585
R378 B.n529 B.n37 585
R379 B.n37 B.n36 585
R380 B.n528 B.n527 585
R381 B.n527 B.n526 585
R382 B.n39 B.n38 585
R383 B.n525 B.n39 585
R384 B.n523 B.n522 585
R385 B.n524 B.n523 585
R386 B.n521 B.n44 585
R387 B.n44 B.n43 585
R388 B.n568 B.n567 585
R389 B.n566 B.n2 585
R390 B.n519 B.n44 478.086
R391 B.n515 B.n78 478.086
R392 B.n279 B.n244 478.086
R393 B.n411 B.n246 478.086
R394 B.n81 B.t17 381.639
R395 B.n79 B.t10 381.639
R396 B.n284 B.t6 381.639
R397 B.n281 B.t14 381.639
R398 B.n517 B.n516 256.663
R399 B.n517 B.n76 256.663
R400 B.n517 B.n75 256.663
R401 B.n517 B.n74 256.663
R402 B.n517 B.n73 256.663
R403 B.n517 B.n72 256.663
R404 B.n517 B.n71 256.663
R405 B.n517 B.n70 256.663
R406 B.n517 B.n69 256.663
R407 B.n517 B.n68 256.663
R408 B.n517 B.n67 256.663
R409 B.n517 B.n66 256.663
R410 B.n517 B.n65 256.663
R411 B.n517 B.n64 256.663
R412 B.n517 B.n63 256.663
R413 B.n517 B.n62 256.663
R414 B.n517 B.n61 256.663
R415 B.n517 B.n60 256.663
R416 B.n517 B.n59 256.663
R417 B.n517 B.n58 256.663
R418 B.n517 B.n57 256.663
R419 B.n517 B.n56 256.663
R420 B.n517 B.n55 256.663
R421 B.n517 B.n54 256.663
R422 B.n517 B.n53 256.663
R423 B.n517 B.n52 256.663
R424 B.n517 B.n51 256.663
R425 B.n517 B.n50 256.663
R426 B.n517 B.n49 256.663
R427 B.n517 B.n48 256.663
R428 B.n517 B.n47 256.663
R429 B.n518 B.n517 256.663
R430 B.n410 B.n409 256.663
R431 B.n409 B.n249 256.663
R432 B.n409 B.n250 256.663
R433 B.n409 B.n251 256.663
R434 B.n409 B.n252 256.663
R435 B.n409 B.n253 256.663
R436 B.n409 B.n254 256.663
R437 B.n409 B.n255 256.663
R438 B.n409 B.n256 256.663
R439 B.n409 B.n257 256.663
R440 B.n409 B.n258 256.663
R441 B.n409 B.n259 256.663
R442 B.n409 B.n260 256.663
R443 B.n409 B.n261 256.663
R444 B.n409 B.n262 256.663
R445 B.n409 B.n263 256.663
R446 B.n409 B.n264 256.663
R447 B.n409 B.n265 256.663
R448 B.n409 B.n266 256.663
R449 B.n409 B.n267 256.663
R450 B.n409 B.n268 256.663
R451 B.n409 B.n269 256.663
R452 B.n409 B.n270 256.663
R453 B.n409 B.n271 256.663
R454 B.n409 B.n272 256.663
R455 B.n409 B.n273 256.663
R456 B.n409 B.n274 256.663
R457 B.n409 B.n275 256.663
R458 B.n409 B.n276 256.663
R459 B.n409 B.n277 256.663
R460 B.n409 B.n278 256.663
R461 B.n570 B.n569 256.663
R462 B.n83 B.n46 163.367
R463 B.n87 B.n86 163.367
R464 B.n91 B.n90 163.367
R465 B.n95 B.n94 163.367
R466 B.n99 B.n98 163.367
R467 B.n103 B.n102 163.367
R468 B.n107 B.n106 163.367
R469 B.n111 B.n110 163.367
R470 B.n115 B.n114 163.367
R471 B.n119 B.n118 163.367
R472 B.n123 B.n122 163.367
R473 B.n127 B.n126 163.367
R474 B.n131 B.n130 163.367
R475 B.n136 B.n135 163.367
R476 B.n140 B.n139 163.367
R477 B.n144 B.n143 163.367
R478 B.n148 B.n147 163.367
R479 B.n152 B.n151 163.367
R480 B.n157 B.n156 163.367
R481 B.n161 B.n160 163.367
R482 B.n165 B.n164 163.367
R483 B.n169 B.n168 163.367
R484 B.n173 B.n172 163.367
R485 B.n177 B.n176 163.367
R486 B.n181 B.n180 163.367
R487 B.n185 B.n184 163.367
R488 B.n189 B.n188 163.367
R489 B.n193 B.n192 163.367
R490 B.n197 B.n196 163.367
R491 B.n201 B.n200 163.367
R492 B.n203 B.n77 163.367
R493 B.n417 B.n244 163.367
R494 B.n417 B.n242 163.367
R495 B.n421 B.n242 163.367
R496 B.n421 B.n236 163.367
R497 B.n429 B.n236 163.367
R498 B.n429 B.n234 163.367
R499 B.n433 B.n234 163.367
R500 B.n433 B.n228 163.367
R501 B.n441 B.n228 163.367
R502 B.n441 B.n226 163.367
R503 B.n445 B.n226 163.367
R504 B.n445 B.n221 163.367
R505 B.n454 B.n221 163.367
R506 B.n454 B.n219 163.367
R507 B.n458 B.n219 163.367
R508 B.n458 B.n214 163.367
R509 B.n467 B.n214 163.367
R510 B.n467 B.n212 163.367
R511 B.n472 B.n212 163.367
R512 B.n472 B.n207 163.367
R513 B.n480 B.n207 163.367
R514 B.n481 B.n480 163.367
R515 B.n481 B.n5 163.367
R516 B.n6 B.n5 163.367
R517 B.n7 B.n6 163.367
R518 B.n487 B.n7 163.367
R519 B.n488 B.n487 163.367
R520 B.n488 B.n12 163.367
R521 B.n13 B.n12 163.367
R522 B.n14 B.n13 163.367
R523 B.n493 B.n14 163.367
R524 B.n493 B.n19 163.367
R525 B.n20 B.n19 163.367
R526 B.n21 B.n20 163.367
R527 B.n498 B.n21 163.367
R528 B.n498 B.n26 163.367
R529 B.n27 B.n26 163.367
R530 B.n28 B.n27 163.367
R531 B.n503 B.n28 163.367
R532 B.n503 B.n33 163.367
R533 B.n34 B.n33 163.367
R534 B.n35 B.n34 163.367
R535 B.n508 B.n35 163.367
R536 B.n508 B.n40 163.367
R537 B.n41 B.n40 163.367
R538 B.n42 B.n41 163.367
R539 B.n78 B.n42 163.367
R540 B.n408 B.n248 163.367
R541 B.n408 B.n280 163.367
R542 B.n404 B.n403 163.367
R543 B.n400 B.n399 163.367
R544 B.n396 B.n395 163.367
R545 B.n392 B.n391 163.367
R546 B.n388 B.n387 163.367
R547 B.n384 B.n383 163.367
R548 B.n380 B.n379 163.367
R549 B.n376 B.n375 163.367
R550 B.n372 B.n371 163.367
R551 B.n368 B.n367 163.367
R552 B.n364 B.n363 163.367
R553 B.n360 B.n359 163.367
R554 B.n356 B.n355 163.367
R555 B.n352 B.n351 163.367
R556 B.n348 B.n347 163.367
R557 B.n344 B.n343 163.367
R558 B.n340 B.n339 163.367
R559 B.n336 B.n335 163.367
R560 B.n332 B.n331 163.367
R561 B.n328 B.n327 163.367
R562 B.n324 B.n323 163.367
R563 B.n320 B.n319 163.367
R564 B.n316 B.n315 163.367
R565 B.n312 B.n311 163.367
R566 B.n308 B.n307 163.367
R567 B.n304 B.n303 163.367
R568 B.n300 B.n299 163.367
R569 B.n296 B.n295 163.367
R570 B.n292 B.n291 163.367
R571 B.n288 B.n279 163.367
R572 B.n415 B.n246 163.367
R573 B.n415 B.n240 163.367
R574 B.n423 B.n240 163.367
R575 B.n423 B.n238 163.367
R576 B.n427 B.n238 163.367
R577 B.n427 B.n232 163.367
R578 B.n435 B.n232 163.367
R579 B.n435 B.n230 163.367
R580 B.n439 B.n230 163.367
R581 B.n439 B.n224 163.367
R582 B.n448 B.n224 163.367
R583 B.n448 B.n222 163.367
R584 B.n452 B.n222 163.367
R585 B.n452 B.n217 163.367
R586 B.n461 B.n217 163.367
R587 B.n461 B.n215 163.367
R588 B.n465 B.n215 163.367
R589 B.n465 B.n210 163.367
R590 B.n474 B.n210 163.367
R591 B.n474 B.n208 163.367
R592 B.n478 B.n208 163.367
R593 B.n478 B.n3 163.367
R594 B.n568 B.n3 163.367
R595 B.n564 B.n2 163.367
R596 B.n564 B.n563 163.367
R597 B.n563 B.n9 163.367
R598 B.n559 B.n9 163.367
R599 B.n559 B.n11 163.367
R600 B.n555 B.n11 163.367
R601 B.n555 B.n15 163.367
R602 B.n551 B.n15 163.367
R603 B.n551 B.n17 163.367
R604 B.n547 B.n17 163.367
R605 B.n547 B.n22 163.367
R606 B.n543 B.n22 163.367
R607 B.n543 B.n24 163.367
R608 B.n539 B.n24 163.367
R609 B.n539 B.n30 163.367
R610 B.n535 B.n30 163.367
R611 B.n535 B.n32 163.367
R612 B.n531 B.n32 163.367
R613 B.n531 B.n37 163.367
R614 B.n527 B.n37 163.367
R615 B.n527 B.n39 163.367
R616 B.n523 B.n39 163.367
R617 B.n523 B.n44 163.367
R618 B.n79 B.t12 100.332
R619 B.n284 B.t9 100.332
R620 B.n81 B.t18 100.323
R621 B.n281 B.t16 100.323
R622 B.n409 B.n245 96.6551
R623 B.n517 B.n43 96.6551
R624 B.n80 B.t13 75.3134
R625 B.n285 B.t8 75.3134
R626 B.n82 B.t19 75.3057
R627 B.n282 B.t15 75.3057
R628 B.n519 B.n518 71.676
R629 B.n83 B.n47 71.676
R630 B.n87 B.n48 71.676
R631 B.n91 B.n49 71.676
R632 B.n95 B.n50 71.676
R633 B.n99 B.n51 71.676
R634 B.n103 B.n52 71.676
R635 B.n107 B.n53 71.676
R636 B.n111 B.n54 71.676
R637 B.n115 B.n55 71.676
R638 B.n119 B.n56 71.676
R639 B.n123 B.n57 71.676
R640 B.n127 B.n58 71.676
R641 B.n131 B.n59 71.676
R642 B.n136 B.n60 71.676
R643 B.n140 B.n61 71.676
R644 B.n144 B.n62 71.676
R645 B.n148 B.n63 71.676
R646 B.n152 B.n64 71.676
R647 B.n157 B.n65 71.676
R648 B.n161 B.n66 71.676
R649 B.n165 B.n67 71.676
R650 B.n169 B.n68 71.676
R651 B.n173 B.n69 71.676
R652 B.n177 B.n70 71.676
R653 B.n181 B.n71 71.676
R654 B.n185 B.n72 71.676
R655 B.n189 B.n73 71.676
R656 B.n193 B.n74 71.676
R657 B.n197 B.n75 71.676
R658 B.n201 B.n76 71.676
R659 B.n516 B.n77 71.676
R660 B.n516 B.n515 71.676
R661 B.n203 B.n76 71.676
R662 B.n200 B.n75 71.676
R663 B.n196 B.n74 71.676
R664 B.n192 B.n73 71.676
R665 B.n188 B.n72 71.676
R666 B.n184 B.n71 71.676
R667 B.n180 B.n70 71.676
R668 B.n176 B.n69 71.676
R669 B.n172 B.n68 71.676
R670 B.n168 B.n67 71.676
R671 B.n164 B.n66 71.676
R672 B.n160 B.n65 71.676
R673 B.n156 B.n64 71.676
R674 B.n151 B.n63 71.676
R675 B.n147 B.n62 71.676
R676 B.n143 B.n61 71.676
R677 B.n139 B.n60 71.676
R678 B.n135 B.n59 71.676
R679 B.n130 B.n58 71.676
R680 B.n126 B.n57 71.676
R681 B.n122 B.n56 71.676
R682 B.n118 B.n55 71.676
R683 B.n114 B.n54 71.676
R684 B.n110 B.n53 71.676
R685 B.n106 B.n52 71.676
R686 B.n102 B.n51 71.676
R687 B.n98 B.n50 71.676
R688 B.n94 B.n49 71.676
R689 B.n90 B.n48 71.676
R690 B.n86 B.n47 71.676
R691 B.n518 B.n46 71.676
R692 B.n411 B.n410 71.676
R693 B.n280 B.n249 71.676
R694 B.n403 B.n250 71.676
R695 B.n399 B.n251 71.676
R696 B.n395 B.n252 71.676
R697 B.n391 B.n253 71.676
R698 B.n387 B.n254 71.676
R699 B.n383 B.n255 71.676
R700 B.n379 B.n256 71.676
R701 B.n375 B.n257 71.676
R702 B.n371 B.n258 71.676
R703 B.n367 B.n259 71.676
R704 B.n363 B.n260 71.676
R705 B.n359 B.n261 71.676
R706 B.n355 B.n262 71.676
R707 B.n351 B.n263 71.676
R708 B.n347 B.n264 71.676
R709 B.n343 B.n265 71.676
R710 B.n339 B.n266 71.676
R711 B.n335 B.n267 71.676
R712 B.n331 B.n268 71.676
R713 B.n327 B.n269 71.676
R714 B.n323 B.n270 71.676
R715 B.n319 B.n271 71.676
R716 B.n315 B.n272 71.676
R717 B.n311 B.n273 71.676
R718 B.n307 B.n274 71.676
R719 B.n303 B.n275 71.676
R720 B.n299 B.n276 71.676
R721 B.n295 B.n277 71.676
R722 B.n291 B.n278 71.676
R723 B.n410 B.n248 71.676
R724 B.n404 B.n249 71.676
R725 B.n400 B.n250 71.676
R726 B.n396 B.n251 71.676
R727 B.n392 B.n252 71.676
R728 B.n388 B.n253 71.676
R729 B.n384 B.n254 71.676
R730 B.n380 B.n255 71.676
R731 B.n376 B.n256 71.676
R732 B.n372 B.n257 71.676
R733 B.n368 B.n258 71.676
R734 B.n364 B.n259 71.676
R735 B.n360 B.n260 71.676
R736 B.n356 B.n261 71.676
R737 B.n352 B.n262 71.676
R738 B.n348 B.n263 71.676
R739 B.n344 B.n264 71.676
R740 B.n340 B.n265 71.676
R741 B.n336 B.n266 71.676
R742 B.n332 B.n267 71.676
R743 B.n328 B.n268 71.676
R744 B.n324 B.n269 71.676
R745 B.n320 B.n270 71.676
R746 B.n316 B.n271 71.676
R747 B.n312 B.n272 71.676
R748 B.n308 B.n273 71.676
R749 B.n304 B.n274 71.676
R750 B.n300 B.n275 71.676
R751 B.n296 B.n276 71.676
R752 B.n292 B.n277 71.676
R753 B.n288 B.n278 71.676
R754 B.n569 B.n568 71.676
R755 B.n569 B.n2 71.676
R756 B.n416 B.n245 60.2988
R757 B.n416 B.n241 60.2988
R758 B.n422 B.n241 60.2988
R759 B.n422 B.n237 60.2988
R760 B.n428 B.n237 60.2988
R761 B.n434 B.n233 60.2988
R762 B.n434 B.n229 60.2988
R763 B.n440 B.n229 60.2988
R764 B.n440 B.n225 60.2988
R765 B.n447 B.n225 60.2988
R766 B.n447 B.n446 60.2988
R767 B.n453 B.n218 60.2988
R768 B.n460 B.n218 60.2988
R769 B.n460 B.n459 60.2988
R770 B.n466 B.n211 60.2988
R771 B.n473 B.n211 60.2988
R772 B.n473 B.t3 60.2988
R773 B.n479 B.t3 60.2988
R774 B.n479 B.n4 60.2988
R775 B.n567 B.n4 60.2988
R776 B.n567 B.n566 60.2988
R777 B.n566 B.n565 60.2988
R778 B.n565 B.n8 60.2988
R779 B.t0 B.n8 60.2988
R780 B.n558 B.t0 60.2988
R781 B.n558 B.n557 60.2988
R782 B.n557 B.n556 60.2988
R783 B.n550 B.n18 60.2988
R784 B.n550 B.n549 60.2988
R785 B.n549 B.n548 60.2988
R786 B.n542 B.n25 60.2988
R787 B.n542 B.n541 60.2988
R788 B.n541 B.n540 60.2988
R789 B.n540 B.n29 60.2988
R790 B.n534 B.n29 60.2988
R791 B.n534 B.n533 60.2988
R792 B.n532 B.n36 60.2988
R793 B.n526 B.n36 60.2988
R794 B.n526 B.n525 60.2988
R795 B.n525 B.n524 60.2988
R796 B.n524 B.n43 60.2988
R797 B.n133 B.n82 59.5399
R798 B.n154 B.n80 59.5399
R799 B.n286 B.n285 59.5399
R800 B.n283 B.n282 59.5399
R801 B.n466 B.t2 47.8844
R802 B.n556 B.t1 47.8844
R803 B.t7 B.n233 35.4701
R804 B.n453 B.t5 35.4701
R805 B.n548 B.t4 35.4701
R806 B.n533 B.t11 35.4701
R807 B.n413 B.n412 31.0639
R808 B.n287 B.n243 31.0639
R809 B.n514 B.n513 31.0639
R810 B.n521 B.n520 31.0639
R811 B.n82 B.n81 25.0187
R812 B.n80 B.n79 25.0187
R813 B.n285 B.n284 25.0187
R814 B.n282 B.n281 25.0187
R815 B.n428 B.t7 24.8292
R816 B.n446 B.t5 24.8292
R817 B.n25 B.t4 24.8292
R818 B.t11 B.n532 24.8292
R819 B B.n570 18.0485
R820 B.n459 B.t2 12.4148
R821 B.n18 B.t1 12.4148
R822 B.n414 B.n413 10.6151
R823 B.n414 B.n239 10.6151
R824 B.n424 B.n239 10.6151
R825 B.n425 B.n424 10.6151
R826 B.n426 B.n425 10.6151
R827 B.n426 B.n231 10.6151
R828 B.n436 B.n231 10.6151
R829 B.n437 B.n436 10.6151
R830 B.n438 B.n437 10.6151
R831 B.n438 B.n223 10.6151
R832 B.n449 B.n223 10.6151
R833 B.n450 B.n449 10.6151
R834 B.n451 B.n450 10.6151
R835 B.n451 B.n216 10.6151
R836 B.n462 B.n216 10.6151
R837 B.n463 B.n462 10.6151
R838 B.n464 B.n463 10.6151
R839 B.n464 B.n209 10.6151
R840 B.n475 B.n209 10.6151
R841 B.n476 B.n475 10.6151
R842 B.n477 B.n476 10.6151
R843 B.n477 B.n0 10.6151
R844 B.n412 B.n247 10.6151
R845 B.n407 B.n247 10.6151
R846 B.n407 B.n406 10.6151
R847 B.n406 B.n405 10.6151
R848 B.n405 B.n402 10.6151
R849 B.n402 B.n401 10.6151
R850 B.n401 B.n398 10.6151
R851 B.n398 B.n397 10.6151
R852 B.n397 B.n394 10.6151
R853 B.n394 B.n393 10.6151
R854 B.n393 B.n390 10.6151
R855 B.n390 B.n389 10.6151
R856 B.n389 B.n386 10.6151
R857 B.n386 B.n385 10.6151
R858 B.n385 B.n382 10.6151
R859 B.n382 B.n381 10.6151
R860 B.n381 B.n378 10.6151
R861 B.n378 B.n377 10.6151
R862 B.n377 B.n374 10.6151
R863 B.n374 B.n373 10.6151
R864 B.n373 B.n370 10.6151
R865 B.n370 B.n369 10.6151
R866 B.n369 B.n366 10.6151
R867 B.n366 B.n365 10.6151
R868 B.n365 B.n362 10.6151
R869 B.n362 B.n361 10.6151
R870 B.n358 B.n357 10.6151
R871 B.n357 B.n354 10.6151
R872 B.n354 B.n353 10.6151
R873 B.n353 B.n350 10.6151
R874 B.n350 B.n349 10.6151
R875 B.n349 B.n346 10.6151
R876 B.n346 B.n345 10.6151
R877 B.n345 B.n342 10.6151
R878 B.n342 B.n341 10.6151
R879 B.n338 B.n337 10.6151
R880 B.n337 B.n334 10.6151
R881 B.n334 B.n333 10.6151
R882 B.n333 B.n330 10.6151
R883 B.n330 B.n329 10.6151
R884 B.n329 B.n326 10.6151
R885 B.n326 B.n325 10.6151
R886 B.n325 B.n322 10.6151
R887 B.n322 B.n321 10.6151
R888 B.n321 B.n318 10.6151
R889 B.n318 B.n317 10.6151
R890 B.n317 B.n314 10.6151
R891 B.n314 B.n313 10.6151
R892 B.n313 B.n310 10.6151
R893 B.n310 B.n309 10.6151
R894 B.n309 B.n306 10.6151
R895 B.n306 B.n305 10.6151
R896 B.n305 B.n302 10.6151
R897 B.n302 B.n301 10.6151
R898 B.n301 B.n298 10.6151
R899 B.n298 B.n297 10.6151
R900 B.n297 B.n294 10.6151
R901 B.n294 B.n293 10.6151
R902 B.n293 B.n290 10.6151
R903 B.n290 B.n289 10.6151
R904 B.n289 B.n287 10.6151
R905 B.n418 B.n243 10.6151
R906 B.n419 B.n418 10.6151
R907 B.n420 B.n419 10.6151
R908 B.n420 B.n235 10.6151
R909 B.n430 B.n235 10.6151
R910 B.n431 B.n430 10.6151
R911 B.n432 B.n431 10.6151
R912 B.n432 B.n227 10.6151
R913 B.n442 B.n227 10.6151
R914 B.n443 B.n442 10.6151
R915 B.n444 B.n443 10.6151
R916 B.n444 B.n220 10.6151
R917 B.n455 B.n220 10.6151
R918 B.n456 B.n455 10.6151
R919 B.n457 B.n456 10.6151
R920 B.n457 B.n213 10.6151
R921 B.n468 B.n213 10.6151
R922 B.n469 B.n468 10.6151
R923 B.n471 B.n469 10.6151
R924 B.n471 B.n470 10.6151
R925 B.n470 B.n206 10.6151
R926 B.n482 B.n206 10.6151
R927 B.n483 B.n482 10.6151
R928 B.n484 B.n483 10.6151
R929 B.n485 B.n484 10.6151
R930 B.n486 B.n485 10.6151
R931 B.n489 B.n486 10.6151
R932 B.n490 B.n489 10.6151
R933 B.n491 B.n490 10.6151
R934 B.n492 B.n491 10.6151
R935 B.n494 B.n492 10.6151
R936 B.n495 B.n494 10.6151
R937 B.n496 B.n495 10.6151
R938 B.n497 B.n496 10.6151
R939 B.n499 B.n497 10.6151
R940 B.n500 B.n499 10.6151
R941 B.n501 B.n500 10.6151
R942 B.n502 B.n501 10.6151
R943 B.n504 B.n502 10.6151
R944 B.n505 B.n504 10.6151
R945 B.n506 B.n505 10.6151
R946 B.n507 B.n506 10.6151
R947 B.n509 B.n507 10.6151
R948 B.n510 B.n509 10.6151
R949 B.n511 B.n510 10.6151
R950 B.n512 B.n511 10.6151
R951 B.n513 B.n512 10.6151
R952 B.n562 B.n1 10.6151
R953 B.n562 B.n561 10.6151
R954 B.n561 B.n560 10.6151
R955 B.n560 B.n10 10.6151
R956 B.n554 B.n10 10.6151
R957 B.n554 B.n553 10.6151
R958 B.n553 B.n552 10.6151
R959 B.n552 B.n16 10.6151
R960 B.n546 B.n16 10.6151
R961 B.n546 B.n545 10.6151
R962 B.n545 B.n544 10.6151
R963 B.n544 B.n23 10.6151
R964 B.n538 B.n23 10.6151
R965 B.n538 B.n537 10.6151
R966 B.n537 B.n536 10.6151
R967 B.n536 B.n31 10.6151
R968 B.n530 B.n31 10.6151
R969 B.n530 B.n529 10.6151
R970 B.n529 B.n528 10.6151
R971 B.n528 B.n38 10.6151
R972 B.n522 B.n38 10.6151
R973 B.n522 B.n521 10.6151
R974 B.n520 B.n45 10.6151
R975 B.n84 B.n45 10.6151
R976 B.n85 B.n84 10.6151
R977 B.n88 B.n85 10.6151
R978 B.n89 B.n88 10.6151
R979 B.n92 B.n89 10.6151
R980 B.n93 B.n92 10.6151
R981 B.n96 B.n93 10.6151
R982 B.n97 B.n96 10.6151
R983 B.n100 B.n97 10.6151
R984 B.n101 B.n100 10.6151
R985 B.n104 B.n101 10.6151
R986 B.n105 B.n104 10.6151
R987 B.n108 B.n105 10.6151
R988 B.n109 B.n108 10.6151
R989 B.n112 B.n109 10.6151
R990 B.n113 B.n112 10.6151
R991 B.n116 B.n113 10.6151
R992 B.n117 B.n116 10.6151
R993 B.n120 B.n117 10.6151
R994 B.n121 B.n120 10.6151
R995 B.n124 B.n121 10.6151
R996 B.n125 B.n124 10.6151
R997 B.n128 B.n125 10.6151
R998 B.n129 B.n128 10.6151
R999 B.n132 B.n129 10.6151
R1000 B.n137 B.n134 10.6151
R1001 B.n138 B.n137 10.6151
R1002 B.n141 B.n138 10.6151
R1003 B.n142 B.n141 10.6151
R1004 B.n145 B.n142 10.6151
R1005 B.n146 B.n145 10.6151
R1006 B.n149 B.n146 10.6151
R1007 B.n150 B.n149 10.6151
R1008 B.n153 B.n150 10.6151
R1009 B.n158 B.n155 10.6151
R1010 B.n159 B.n158 10.6151
R1011 B.n162 B.n159 10.6151
R1012 B.n163 B.n162 10.6151
R1013 B.n166 B.n163 10.6151
R1014 B.n167 B.n166 10.6151
R1015 B.n170 B.n167 10.6151
R1016 B.n171 B.n170 10.6151
R1017 B.n174 B.n171 10.6151
R1018 B.n175 B.n174 10.6151
R1019 B.n178 B.n175 10.6151
R1020 B.n179 B.n178 10.6151
R1021 B.n182 B.n179 10.6151
R1022 B.n183 B.n182 10.6151
R1023 B.n186 B.n183 10.6151
R1024 B.n187 B.n186 10.6151
R1025 B.n190 B.n187 10.6151
R1026 B.n191 B.n190 10.6151
R1027 B.n194 B.n191 10.6151
R1028 B.n195 B.n194 10.6151
R1029 B.n198 B.n195 10.6151
R1030 B.n199 B.n198 10.6151
R1031 B.n202 B.n199 10.6151
R1032 B.n204 B.n202 10.6151
R1033 B.n205 B.n204 10.6151
R1034 B.n514 B.n205 10.6151
R1035 B.n361 B.n283 9.36635
R1036 B.n338 B.n286 9.36635
R1037 B.n133 B.n132 9.36635
R1038 B.n155 B.n154 9.36635
R1039 B.n570 B.n0 8.11757
R1040 B.n570 B.n1 8.11757
R1041 B.n358 B.n283 1.24928
R1042 B.n341 B.n286 1.24928
R1043 B.n134 B.n133 1.24928
R1044 B.n154 B.n153 1.24928
R1045 VN.n2 VN.t1 239.105
R1046 VN.n10 VN.t3 239.105
R1047 VN.n6 VN.t4 220.165
R1048 VN.n14 VN.t5 220.165
R1049 VN.n1 VN.t0 178.994
R1050 VN.n9 VN.t2 178.994
R1051 VN.n7 VN.n6 161.3
R1052 VN.n15 VN.n14 161.3
R1053 VN.n13 VN.n8 161.3
R1054 VN.n12 VN.n11 161.3
R1055 VN.n5 VN.n0 161.3
R1056 VN.n4 VN.n3 161.3
R1057 VN.n5 VN.n4 50.6917
R1058 VN.n13 VN.n12 50.6917
R1059 VN.n11 VN.n10 43.2502
R1060 VN.n3 VN.n2 43.2502
R1061 VN.n2 VN.n1 42.2819
R1062 VN.n10 VN.n9 42.2819
R1063 VN VN.n15 38.9835
R1064 VN.n4 VN.n1 12.234
R1065 VN.n12 VN.n9 12.234
R1066 VN.n6 VN.n5 8.76414
R1067 VN.n14 VN.n13 8.76414
R1068 VN.n15 VN.n8 0.189894
R1069 VN.n11 VN.n8 0.189894
R1070 VN.n3 VN.n0 0.189894
R1071 VN.n7 VN.n0 0.189894
R1072 VN VN.n7 0.0516364
R1073 VDD2.n1 VDD2.t4 70.1364
R1074 VDD2.n2 VDD2.t0 69.3579
R1075 VDD2.n1 VDD2.n0 66.8036
R1076 VDD2 VDD2.n3 66.8006
R1077 VDD2.n2 VDD2.n1 33.4761
R1078 VDD2.n3 VDD2.t3 2.7775
R1079 VDD2.n3 VDD2.t2 2.7775
R1080 VDD2.n0 VDD2.t5 2.7775
R1081 VDD2.n0 VDD2.t1 2.7775
R1082 VDD2 VDD2.n2 0.892741
C0 VN VDD2 3.11261f
C1 VN VTAIL 3.13104f
C2 VDD2 VTAIL 6.1783f
C3 VP VN 4.42835f
C4 VP VDD2 0.318835f
C5 VN VDD1 0.148442f
C6 VDD2 VDD1 0.804112f
C7 VP VTAIL 3.1454f
C8 VDD1 VTAIL 6.13921f
C9 VP VDD1 3.28031f
C10 VDD2 B 3.824251f
C11 VDD1 B 4.061924f
C12 VTAIL B 4.646599f
C13 VN B 7.74899f
C14 VP B 6.137735f
C15 VDD2.t4 B 1.38287f
C16 VDD2.t5 B 0.127438f
C17 VDD2.t1 B 0.127438f
C18 VDD2.n0 B 1.08514f
C19 VDD2.n1 B 1.71681f
C20 VDD2.t0 B 1.37949f
C21 VDD2.n2 B 1.76857f
C22 VDD2.t3 B 0.127438f
C23 VDD2.t2 B 0.127438f
C24 VDD2.n3 B 1.08512f
C25 VN.n0 B 0.04147f
C26 VN.t0 B 0.758293f
C27 VN.n1 B 0.344382f
C28 VN.t1 B 0.848121f
C29 VN.n2 B 0.355674f
C30 VN.n3 B 0.178783f
C31 VN.n4 B 0.056631f
C32 VN.n5 B 0.01484f
C33 VN.t4 B 0.819284f
C34 VN.n6 B 0.353203f
C35 VN.n7 B 0.032137f
C36 VN.n8 B 0.04147f
C37 VN.t2 B 0.758293f
C38 VN.n9 B 0.344382f
C39 VN.t3 B 0.848121f
C40 VN.n10 B 0.355674f
C41 VN.n11 B 0.178783f
C42 VN.n12 B 0.056631f
C43 VN.n13 B 0.01484f
C44 VN.t5 B 0.819284f
C45 VN.n14 B 0.353203f
C46 VN.n15 B 1.50824f
C47 VTAIL.t0 B 0.140505f
C48 VTAIL.t1 B 0.140505f
C49 VTAIL.n0 B 1.12838f
C50 VTAIL.n1 B 0.347554f
C51 VTAIL.t9 B 1.43929f
C52 VTAIL.n2 B 0.482178f
C53 VTAIL.t5 B 0.140505f
C54 VTAIL.t7 B 0.140505f
C55 VTAIL.n3 B 1.12838f
C56 VTAIL.n4 B 1.33882f
C57 VTAIL.t11 B 0.140505f
C58 VTAIL.t2 B 0.140505f
C59 VTAIL.n5 B 1.12838f
C60 VTAIL.n6 B 1.33882f
C61 VTAIL.t3 B 1.4393f
C62 VTAIL.n7 B 0.482172f
C63 VTAIL.t8 B 0.140505f
C64 VTAIL.t10 B 0.140505f
C65 VTAIL.n8 B 1.12838f
C66 VTAIL.n9 B 0.409895f
C67 VTAIL.t6 B 1.43929f
C68 VTAIL.n10 B 1.32174f
C69 VTAIL.t4 B 1.43929f
C70 VTAIL.n11 B 1.29473f
C71 VDD1.t5 B 1.38589f
C72 VDD1.t0 B 1.3853f
C73 VDD1.t3 B 0.127661f
C74 VDD1.t4 B 0.127661f
C75 VDD1.n0 B 1.08704f
C76 VDD1.n1 B 1.79308f
C77 VDD1.t1 B 0.127661f
C78 VDD1.t2 B 0.127661f
C79 VDD1.n2 B 1.08606f
C80 VDD1.n3 B 1.76189f
C81 VP.n0 B 0.042486f
C82 VP.t3 B 0.776873f
C83 VP.n1 B 0.310751f
C84 VP.n2 B 0.042486f
C85 VP.n3 B 0.042486f
C86 VP.t4 B 0.839358f
C87 VP.t0 B 0.776873f
C88 VP.n4 B 0.35282f
C89 VP.t2 B 0.868902f
C90 VP.n5 B 0.364389f
C91 VP.n6 B 0.183164f
C92 VP.n7 B 0.058018f
C93 VP.n8 B 0.015204f
C94 VP.n9 B 0.361858f
C95 VP.n10 B 1.51715f
C96 VP.n11 B 1.55671f
C97 VP.t5 B 0.839358f
C98 VP.n12 B 0.361858f
C99 VP.n13 B 0.015204f
C100 VP.n14 B 0.058018f
C101 VP.n15 B 0.042486f
C102 VP.n16 B 0.042486f
C103 VP.n17 B 0.058018f
C104 VP.n18 B 0.015204f
C105 VP.t1 B 0.839358f
C106 VP.n19 B 0.361858f
C107 VP.n20 B 0.032925f
.ends

