* NGSPICE file created from diff_pair_sample_0252.ext - technology: sky130A

.subckt diff_pair_sample_0252 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t13 VN.t0 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X1 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0 ps=0 w=3.11 l=2.24
X2 VTAIL.t15 VP.t0 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0.51315 ps=3.44 w=3.11 l=2.24
X3 VDD1.t6 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=1.2129 ps=7 w=3.11 l=2.24
X4 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X5 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0 ps=0 w=3.11 l=2.24
X6 VDD1.t4 VP.t3 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=1.2129 ps=7 w=3.11 l=2.24
X7 VTAIL.t12 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0.51315 ps=3.44 w=3.11 l=2.24
X8 VTAIL.t11 VN.t2 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X9 VDD2.t0 VN.t3 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X10 VDD2.t4 VN.t4 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=1.2129 ps=7 w=3.11 l=2.24
X11 VTAIL.t5 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0.51315 ps=3.44 w=3.11 l=2.24
X12 VDD2.t5 VN.t5 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=1.2129 ps=7 w=3.11 l=2.24
X13 VTAIL.t7 VN.t6 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0.51315 ps=3.44 w=3.11 l=2.24
X14 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X15 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0 ps=0 w=3.11 l=2.24
X16 VDD1.t1 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X17 VDD2.t3 VN.t7 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2129 pd=7 as=0 ps=0 w=3.11 l=2.24
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.51315 pd=3.44 as=0.51315 ps=3.44 w=3.11 l=2.24
R0 VN.n47 VN.n25 161.3
R1 VN.n46 VN.n45 161.3
R2 VN.n44 VN.n26 161.3
R3 VN.n43 VN.n42 161.3
R4 VN.n41 VN.n27 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n28 161.3
R7 VN.n36 VN.n35 161.3
R8 VN.n34 VN.n29 161.3
R9 VN.n33 VN.n32 161.3
R10 VN.n22 VN.n0 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n1 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n2 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n12 VN.n3 161.3
R17 VN.n11 VN.n10 161.3
R18 VN.n9 VN.n4 161.3
R19 VN.n8 VN.n7 161.3
R20 VN.n24 VN.n23 93.3849
R21 VN.n49 VN.n48 93.3849
R22 VN.n6 VN.t6 66.8891
R23 VN.n31 VN.t4 66.8891
R24 VN.n6 VN.n5 57.3618
R25 VN.n31 VN.n30 57.3618
R26 VN.n21 VN.n1 47.2923
R27 VN.n46 VN.n26 47.2923
R28 VN VN.n49 42.8012
R29 VN.n10 VN.n9 40.4934
R30 VN.n10 VN.n3 40.4934
R31 VN.n35 VN.n34 40.4934
R32 VN.n35 VN.n28 40.4934
R33 VN.n17 VN.n1 33.6945
R34 VN.n42 VN.n26 33.6945
R35 VN.n5 VN.t7 33.4608
R36 VN.n15 VN.t0 33.4608
R37 VN.n23 VN.t5 33.4608
R38 VN.n30 VN.t2 33.4608
R39 VN.n40 VN.t3 33.4608
R40 VN.n48 VN.t1 33.4608
R41 VN.n9 VN.n8 24.4675
R42 VN.n14 VN.n3 24.4675
R43 VN.n17 VN.n16 24.4675
R44 VN.n22 VN.n21 24.4675
R45 VN.n34 VN.n33 24.4675
R46 VN.n42 VN.n41 24.4675
R47 VN.n39 VN.n28 24.4675
R48 VN.n47 VN.n46 24.4675
R49 VN.n23 VN.n22 17.3721
R50 VN.n48 VN.n47 17.3721
R51 VN.n8 VN.n5 13.9467
R52 VN.n15 VN.n14 13.9467
R53 VN.n33 VN.n30 13.9467
R54 VN.n40 VN.n39 13.9467
R55 VN.n16 VN.n15 10.5213
R56 VN.n41 VN.n40 10.5213
R57 VN.n32 VN.n31 9.22138
R58 VN.n7 VN.n6 9.22138
R59 VN.n49 VN.n25 0.278367
R60 VN.n24 VN.n0 0.278367
R61 VN.n45 VN.n25 0.189894
R62 VN.n45 VN.n44 0.189894
R63 VN.n44 VN.n43 0.189894
R64 VN.n43 VN.n27 0.189894
R65 VN.n38 VN.n27 0.189894
R66 VN.n38 VN.n37 0.189894
R67 VN.n37 VN.n36 0.189894
R68 VN.n36 VN.n29 0.189894
R69 VN.n32 VN.n29 0.189894
R70 VN.n7 VN.n4 0.189894
R71 VN.n11 VN.n4 0.189894
R72 VN.n12 VN.n11 0.189894
R73 VN.n13 VN.n12 0.189894
R74 VN.n13 VN.n2 0.189894
R75 VN.n18 VN.n2 0.189894
R76 VN.n19 VN.n18 0.189894
R77 VN.n20 VN.n19 0.189894
R78 VN.n20 VN.n0 0.189894
R79 VN VN.n24 0.153454
R80 VDD2.n2 VDD2.n1 78.6075
R81 VDD2.n2 VDD2.n0 78.6075
R82 VDD2 VDD2.n5 78.6047
R83 VDD2.n4 VDD2.n3 77.5552
R84 VDD2.n4 VDD2.n2 36.3662
R85 VDD2.n5 VDD2.t7 6.36706
R86 VDD2.n5 VDD2.t4 6.36706
R87 VDD2.n3 VDD2.t6 6.36706
R88 VDD2.n3 VDD2.t0 6.36706
R89 VDD2.n1 VDD2.t1 6.36706
R90 VDD2.n1 VDD2.t5 6.36706
R91 VDD2.n0 VDD2.t2 6.36706
R92 VDD2.n0 VDD2.t3 6.36706
R93 VDD2 VDD2.n4 1.16645
R94 VTAIL.n130 VTAIL.n120 289.615
R95 VTAIL.n12 VTAIL.n2 289.615
R96 VTAIL.n28 VTAIL.n18 289.615
R97 VTAIL.n46 VTAIL.n36 289.615
R98 VTAIL.n114 VTAIL.n104 289.615
R99 VTAIL.n96 VTAIL.n86 289.615
R100 VTAIL.n80 VTAIL.n70 289.615
R101 VTAIL.n62 VTAIL.n52 289.615
R102 VTAIL.n124 VTAIL.n123 185
R103 VTAIL.n129 VTAIL.n128 185
R104 VTAIL.n131 VTAIL.n130 185
R105 VTAIL.n6 VTAIL.n5 185
R106 VTAIL.n11 VTAIL.n10 185
R107 VTAIL.n13 VTAIL.n12 185
R108 VTAIL.n22 VTAIL.n21 185
R109 VTAIL.n27 VTAIL.n26 185
R110 VTAIL.n29 VTAIL.n28 185
R111 VTAIL.n40 VTAIL.n39 185
R112 VTAIL.n45 VTAIL.n44 185
R113 VTAIL.n47 VTAIL.n46 185
R114 VTAIL.n115 VTAIL.n114 185
R115 VTAIL.n113 VTAIL.n112 185
R116 VTAIL.n108 VTAIL.n107 185
R117 VTAIL.n97 VTAIL.n96 185
R118 VTAIL.n95 VTAIL.n94 185
R119 VTAIL.n90 VTAIL.n89 185
R120 VTAIL.n81 VTAIL.n80 185
R121 VTAIL.n79 VTAIL.n78 185
R122 VTAIL.n74 VTAIL.n73 185
R123 VTAIL.n63 VTAIL.n62 185
R124 VTAIL.n61 VTAIL.n60 185
R125 VTAIL.n56 VTAIL.n55 185
R126 VTAIL.n125 VTAIL.t8 148.606
R127 VTAIL.n7 VTAIL.t7 148.606
R128 VTAIL.n23 VTAIL.t2 148.606
R129 VTAIL.n41 VTAIL.t15 148.606
R130 VTAIL.n109 VTAIL.t14 148.606
R131 VTAIL.n91 VTAIL.t5 148.606
R132 VTAIL.n75 VTAIL.t9 148.606
R133 VTAIL.n57 VTAIL.t12 148.606
R134 VTAIL.n129 VTAIL.n123 104.615
R135 VTAIL.n130 VTAIL.n129 104.615
R136 VTAIL.n11 VTAIL.n5 104.615
R137 VTAIL.n12 VTAIL.n11 104.615
R138 VTAIL.n27 VTAIL.n21 104.615
R139 VTAIL.n28 VTAIL.n27 104.615
R140 VTAIL.n45 VTAIL.n39 104.615
R141 VTAIL.n46 VTAIL.n45 104.615
R142 VTAIL.n114 VTAIL.n113 104.615
R143 VTAIL.n113 VTAIL.n107 104.615
R144 VTAIL.n96 VTAIL.n95 104.615
R145 VTAIL.n95 VTAIL.n89 104.615
R146 VTAIL.n80 VTAIL.n79 104.615
R147 VTAIL.n79 VTAIL.n73 104.615
R148 VTAIL.n62 VTAIL.n61 104.615
R149 VTAIL.n61 VTAIL.n55 104.615
R150 VTAIL.n103 VTAIL.n102 60.8765
R151 VTAIL.n69 VTAIL.n68 60.8765
R152 VTAIL.n1 VTAIL.n0 60.8763
R153 VTAIL.n35 VTAIL.n34 60.8763
R154 VTAIL.t8 VTAIL.n123 52.3082
R155 VTAIL.t7 VTAIL.n5 52.3082
R156 VTAIL.t2 VTAIL.n21 52.3082
R157 VTAIL.t15 VTAIL.n39 52.3082
R158 VTAIL.t14 VTAIL.n107 52.3082
R159 VTAIL.t5 VTAIL.n89 52.3082
R160 VTAIL.t9 VTAIL.n73 52.3082
R161 VTAIL.t12 VTAIL.n55 52.3082
R162 VTAIL.n135 VTAIL.n134 31.9914
R163 VTAIL.n17 VTAIL.n16 31.9914
R164 VTAIL.n33 VTAIL.n32 31.9914
R165 VTAIL.n51 VTAIL.n50 31.9914
R166 VTAIL.n119 VTAIL.n118 31.9914
R167 VTAIL.n101 VTAIL.n100 31.9914
R168 VTAIL.n85 VTAIL.n84 31.9914
R169 VTAIL.n67 VTAIL.n66 31.9914
R170 VTAIL.n135 VTAIL.n119 17.2634
R171 VTAIL.n67 VTAIL.n51 17.2634
R172 VTAIL.n125 VTAIL.n124 15.5966
R173 VTAIL.n7 VTAIL.n6 15.5966
R174 VTAIL.n23 VTAIL.n22 15.5966
R175 VTAIL.n41 VTAIL.n40 15.5966
R176 VTAIL.n109 VTAIL.n108 15.5966
R177 VTAIL.n91 VTAIL.n90 15.5966
R178 VTAIL.n75 VTAIL.n74 15.5966
R179 VTAIL.n57 VTAIL.n56 15.5966
R180 VTAIL.n128 VTAIL.n127 12.8005
R181 VTAIL.n10 VTAIL.n9 12.8005
R182 VTAIL.n26 VTAIL.n25 12.8005
R183 VTAIL.n44 VTAIL.n43 12.8005
R184 VTAIL.n112 VTAIL.n111 12.8005
R185 VTAIL.n94 VTAIL.n93 12.8005
R186 VTAIL.n78 VTAIL.n77 12.8005
R187 VTAIL.n60 VTAIL.n59 12.8005
R188 VTAIL.n131 VTAIL.n122 12.0247
R189 VTAIL.n13 VTAIL.n4 12.0247
R190 VTAIL.n29 VTAIL.n20 12.0247
R191 VTAIL.n47 VTAIL.n38 12.0247
R192 VTAIL.n115 VTAIL.n106 12.0247
R193 VTAIL.n97 VTAIL.n88 12.0247
R194 VTAIL.n81 VTAIL.n72 12.0247
R195 VTAIL.n63 VTAIL.n54 12.0247
R196 VTAIL.n132 VTAIL.n120 11.249
R197 VTAIL.n14 VTAIL.n2 11.249
R198 VTAIL.n30 VTAIL.n18 11.249
R199 VTAIL.n48 VTAIL.n36 11.249
R200 VTAIL.n116 VTAIL.n104 11.249
R201 VTAIL.n98 VTAIL.n86 11.249
R202 VTAIL.n82 VTAIL.n70 11.249
R203 VTAIL.n64 VTAIL.n52 11.249
R204 VTAIL.n134 VTAIL.n133 9.45567
R205 VTAIL.n16 VTAIL.n15 9.45567
R206 VTAIL.n32 VTAIL.n31 9.45567
R207 VTAIL.n50 VTAIL.n49 9.45567
R208 VTAIL.n118 VTAIL.n117 9.45567
R209 VTAIL.n100 VTAIL.n99 9.45567
R210 VTAIL.n84 VTAIL.n83 9.45567
R211 VTAIL.n66 VTAIL.n65 9.45567
R212 VTAIL.n133 VTAIL.n132 9.3005
R213 VTAIL.n122 VTAIL.n121 9.3005
R214 VTAIL.n127 VTAIL.n126 9.3005
R215 VTAIL.n15 VTAIL.n14 9.3005
R216 VTAIL.n4 VTAIL.n3 9.3005
R217 VTAIL.n9 VTAIL.n8 9.3005
R218 VTAIL.n31 VTAIL.n30 9.3005
R219 VTAIL.n20 VTAIL.n19 9.3005
R220 VTAIL.n25 VTAIL.n24 9.3005
R221 VTAIL.n49 VTAIL.n48 9.3005
R222 VTAIL.n38 VTAIL.n37 9.3005
R223 VTAIL.n43 VTAIL.n42 9.3005
R224 VTAIL.n117 VTAIL.n116 9.3005
R225 VTAIL.n106 VTAIL.n105 9.3005
R226 VTAIL.n111 VTAIL.n110 9.3005
R227 VTAIL.n99 VTAIL.n98 9.3005
R228 VTAIL.n88 VTAIL.n87 9.3005
R229 VTAIL.n93 VTAIL.n92 9.3005
R230 VTAIL.n83 VTAIL.n82 9.3005
R231 VTAIL.n72 VTAIL.n71 9.3005
R232 VTAIL.n77 VTAIL.n76 9.3005
R233 VTAIL.n65 VTAIL.n64 9.3005
R234 VTAIL.n54 VTAIL.n53 9.3005
R235 VTAIL.n59 VTAIL.n58 9.3005
R236 VTAIL.n0 VTAIL.t6 6.36706
R237 VTAIL.n0 VTAIL.t13 6.36706
R238 VTAIL.n34 VTAIL.t0 6.36706
R239 VTAIL.n34 VTAIL.t1 6.36706
R240 VTAIL.n102 VTAIL.t3 6.36706
R241 VTAIL.n102 VTAIL.t4 6.36706
R242 VTAIL.n68 VTAIL.t10 6.36706
R243 VTAIL.n68 VTAIL.t11 6.36706
R244 VTAIL.n126 VTAIL.n125 4.46457
R245 VTAIL.n8 VTAIL.n7 4.46457
R246 VTAIL.n24 VTAIL.n23 4.46457
R247 VTAIL.n42 VTAIL.n41 4.46457
R248 VTAIL.n110 VTAIL.n109 4.46457
R249 VTAIL.n92 VTAIL.n91 4.46457
R250 VTAIL.n76 VTAIL.n75 4.46457
R251 VTAIL.n58 VTAIL.n57 4.46457
R252 VTAIL.n134 VTAIL.n120 2.71565
R253 VTAIL.n16 VTAIL.n2 2.71565
R254 VTAIL.n32 VTAIL.n18 2.71565
R255 VTAIL.n50 VTAIL.n36 2.71565
R256 VTAIL.n118 VTAIL.n104 2.71565
R257 VTAIL.n100 VTAIL.n86 2.71565
R258 VTAIL.n84 VTAIL.n70 2.71565
R259 VTAIL.n66 VTAIL.n52 2.71565
R260 VTAIL.n69 VTAIL.n67 2.21602
R261 VTAIL.n85 VTAIL.n69 2.21602
R262 VTAIL.n103 VTAIL.n101 2.21602
R263 VTAIL.n119 VTAIL.n103 2.21602
R264 VTAIL.n51 VTAIL.n35 2.21602
R265 VTAIL.n35 VTAIL.n33 2.21602
R266 VTAIL.n17 VTAIL.n1 2.21602
R267 VTAIL VTAIL.n135 2.15783
R268 VTAIL.n132 VTAIL.n131 1.93989
R269 VTAIL.n14 VTAIL.n13 1.93989
R270 VTAIL.n30 VTAIL.n29 1.93989
R271 VTAIL.n48 VTAIL.n47 1.93989
R272 VTAIL.n116 VTAIL.n115 1.93989
R273 VTAIL.n98 VTAIL.n97 1.93989
R274 VTAIL.n82 VTAIL.n81 1.93989
R275 VTAIL.n64 VTAIL.n63 1.93989
R276 VTAIL.n128 VTAIL.n122 1.16414
R277 VTAIL.n10 VTAIL.n4 1.16414
R278 VTAIL.n26 VTAIL.n20 1.16414
R279 VTAIL.n44 VTAIL.n38 1.16414
R280 VTAIL.n112 VTAIL.n106 1.16414
R281 VTAIL.n94 VTAIL.n88 1.16414
R282 VTAIL.n78 VTAIL.n72 1.16414
R283 VTAIL.n60 VTAIL.n54 1.16414
R284 VTAIL.n101 VTAIL.n85 0.470328
R285 VTAIL.n33 VTAIL.n17 0.470328
R286 VTAIL.n127 VTAIL.n124 0.388379
R287 VTAIL.n9 VTAIL.n6 0.388379
R288 VTAIL.n25 VTAIL.n22 0.388379
R289 VTAIL.n43 VTAIL.n40 0.388379
R290 VTAIL.n111 VTAIL.n108 0.388379
R291 VTAIL.n93 VTAIL.n90 0.388379
R292 VTAIL.n77 VTAIL.n74 0.388379
R293 VTAIL.n59 VTAIL.n56 0.388379
R294 VTAIL.n126 VTAIL.n121 0.155672
R295 VTAIL.n133 VTAIL.n121 0.155672
R296 VTAIL.n8 VTAIL.n3 0.155672
R297 VTAIL.n15 VTAIL.n3 0.155672
R298 VTAIL.n24 VTAIL.n19 0.155672
R299 VTAIL.n31 VTAIL.n19 0.155672
R300 VTAIL.n42 VTAIL.n37 0.155672
R301 VTAIL.n49 VTAIL.n37 0.155672
R302 VTAIL.n117 VTAIL.n105 0.155672
R303 VTAIL.n110 VTAIL.n105 0.155672
R304 VTAIL.n99 VTAIL.n87 0.155672
R305 VTAIL.n92 VTAIL.n87 0.155672
R306 VTAIL.n83 VTAIL.n71 0.155672
R307 VTAIL.n76 VTAIL.n71 0.155672
R308 VTAIL.n65 VTAIL.n53 0.155672
R309 VTAIL.n58 VTAIL.n53 0.155672
R310 VTAIL VTAIL.n1 0.0586897
R311 B.n503 B.n502 585
R312 B.n505 B.n110 585
R313 B.n508 B.n507 585
R314 B.n509 B.n109 585
R315 B.n511 B.n510 585
R316 B.n513 B.n108 585
R317 B.n516 B.n515 585
R318 B.n517 B.n107 585
R319 B.n519 B.n518 585
R320 B.n521 B.n106 585
R321 B.n524 B.n523 585
R322 B.n525 B.n105 585
R323 B.n527 B.n526 585
R324 B.n529 B.n104 585
R325 B.n532 B.n531 585
R326 B.n534 B.n101 585
R327 B.n536 B.n535 585
R328 B.n538 B.n100 585
R329 B.n541 B.n540 585
R330 B.n542 B.n99 585
R331 B.n544 B.n543 585
R332 B.n546 B.n98 585
R333 B.n549 B.n548 585
R334 B.n550 B.n94 585
R335 B.n552 B.n551 585
R336 B.n554 B.n93 585
R337 B.n557 B.n556 585
R338 B.n558 B.n92 585
R339 B.n560 B.n559 585
R340 B.n562 B.n91 585
R341 B.n565 B.n564 585
R342 B.n566 B.n90 585
R343 B.n568 B.n567 585
R344 B.n570 B.n89 585
R345 B.n573 B.n572 585
R346 B.n574 B.n88 585
R347 B.n576 B.n575 585
R348 B.n578 B.n87 585
R349 B.n581 B.n580 585
R350 B.n582 B.n86 585
R351 B.n501 B.n84 585
R352 B.n585 B.n84 585
R353 B.n500 B.n83 585
R354 B.n586 B.n83 585
R355 B.n499 B.n82 585
R356 B.n587 B.n82 585
R357 B.n498 B.n497 585
R358 B.n497 B.n78 585
R359 B.n496 B.n77 585
R360 B.n593 B.n77 585
R361 B.n495 B.n76 585
R362 B.n594 B.n76 585
R363 B.n494 B.n75 585
R364 B.n595 B.n75 585
R365 B.n493 B.n492 585
R366 B.n492 B.n74 585
R367 B.n491 B.n70 585
R368 B.n601 B.n70 585
R369 B.n490 B.n69 585
R370 B.n602 B.n69 585
R371 B.n489 B.n68 585
R372 B.n603 B.n68 585
R373 B.n488 B.n487 585
R374 B.n487 B.n64 585
R375 B.n486 B.n63 585
R376 B.n609 B.n63 585
R377 B.n485 B.n62 585
R378 B.n610 B.n62 585
R379 B.n484 B.n61 585
R380 B.n611 B.n61 585
R381 B.n483 B.n482 585
R382 B.n482 B.n57 585
R383 B.n481 B.n56 585
R384 B.n617 B.n56 585
R385 B.n480 B.n55 585
R386 B.n618 B.n55 585
R387 B.n479 B.n54 585
R388 B.n619 B.n54 585
R389 B.n478 B.n477 585
R390 B.n477 B.n50 585
R391 B.n476 B.n49 585
R392 B.n625 B.n49 585
R393 B.n475 B.n48 585
R394 B.n626 B.n48 585
R395 B.n474 B.n47 585
R396 B.n627 B.n47 585
R397 B.n473 B.n472 585
R398 B.n472 B.n43 585
R399 B.n471 B.n42 585
R400 B.n633 B.n42 585
R401 B.n470 B.n41 585
R402 B.n634 B.n41 585
R403 B.n469 B.n40 585
R404 B.n635 B.n40 585
R405 B.n468 B.n467 585
R406 B.n467 B.n36 585
R407 B.n466 B.n35 585
R408 B.n641 B.n35 585
R409 B.n465 B.n34 585
R410 B.n642 B.n34 585
R411 B.n464 B.n33 585
R412 B.n643 B.n33 585
R413 B.n463 B.n462 585
R414 B.n462 B.n29 585
R415 B.n461 B.n28 585
R416 B.n649 B.n28 585
R417 B.n460 B.n27 585
R418 B.n650 B.n27 585
R419 B.n459 B.n26 585
R420 B.n651 B.n26 585
R421 B.n458 B.n457 585
R422 B.n457 B.n22 585
R423 B.n456 B.n21 585
R424 B.n657 B.n21 585
R425 B.n455 B.n20 585
R426 B.n658 B.n20 585
R427 B.n454 B.n19 585
R428 B.n659 B.n19 585
R429 B.n453 B.n452 585
R430 B.n452 B.n15 585
R431 B.n451 B.n14 585
R432 B.n665 B.n14 585
R433 B.n450 B.n13 585
R434 B.n666 B.n13 585
R435 B.n449 B.n12 585
R436 B.n667 B.n12 585
R437 B.n448 B.n447 585
R438 B.n447 B.n8 585
R439 B.n446 B.n7 585
R440 B.n673 B.n7 585
R441 B.n445 B.n6 585
R442 B.n674 B.n6 585
R443 B.n444 B.n5 585
R444 B.n675 B.n5 585
R445 B.n443 B.n442 585
R446 B.n442 B.n4 585
R447 B.n441 B.n111 585
R448 B.n441 B.n440 585
R449 B.n431 B.n112 585
R450 B.n113 B.n112 585
R451 B.n433 B.n432 585
R452 B.n434 B.n433 585
R453 B.n430 B.n118 585
R454 B.n118 B.n117 585
R455 B.n429 B.n428 585
R456 B.n428 B.n427 585
R457 B.n120 B.n119 585
R458 B.n121 B.n120 585
R459 B.n420 B.n419 585
R460 B.n421 B.n420 585
R461 B.n418 B.n126 585
R462 B.n126 B.n125 585
R463 B.n417 B.n416 585
R464 B.n416 B.n415 585
R465 B.n128 B.n127 585
R466 B.n129 B.n128 585
R467 B.n408 B.n407 585
R468 B.n409 B.n408 585
R469 B.n406 B.n133 585
R470 B.n137 B.n133 585
R471 B.n405 B.n404 585
R472 B.n404 B.n403 585
R473 B.n135 B.n134 585
R474 B.n136 B.n135 585
R475 B.n396 B.n395 585
R476 B.n397 B.n396 585
R477 B.n394 B.n142 585
R478 B.n142 B.n141 585
R479 B.n393 B.n392 585
R480 B.n392 B.n391 585
R481 B.n144 B.n143 585
R482 B.n145 B.n144 585
R483 B.n384 B.n383 585
R484 B.n385 B.n384 585
R485 B.n382 B.n149 585
R486 B.n153 B.n149 585
R487 B.n381 B.n380 585
R488 B.n380 B.n379 585
R489 B.n151 B.n150 585
R490 B.n152 B.n151 585
R491 B.n372 B.n371 585
R492 B.n373 B.n372 585
R493 B.n370 B.n158 585
R494 B.n158 B.n157 585
R495 B.n369 B.n368 585
R496 B.n368 B.n367 585
R497 B.n160 B.n159 585
R498 B.n161 B.n160 585
R499 B.n360 B.n359 585
R500 B.n361 B.n360 585
R501 B.n358 B.n165 585
R502 B.n169 B.n165 585
R503 B.n357 B.n356 585
R504 B.n356 B.n355 585
R505 B.n167 B.n166 585
R506 B.n168 B.n167 585
R507 B.n348 B.n347 585
R508 B.n349 B.n348 585
R509 B.n346 B.n174 585
R510 B.n174 B.n173 585
R511 B.n345 B.n344 585
R512 B.n344 B.n343 585
R513 B.n176 B.n175 585
R514 B.n177 B.n176 585
R515 B.n336 B.n335 585
R516 B.n337 B.n336 585
R517 B.n334 B.n182 585
R518 B.n182 B.n181 585
R519 B.n333 B.n332 585
R520 B.n332 B.n331 585
R521 B.n184 B.n183 585
R522 B.n324 B.n184 585
R523 B.n323 B.n322 585
R524 B.n325 B.n323 585
R525 B.n321 B.n189 585
R526 B.n189 B.n188 585
R527 B.n320 B.n319 585
R528 B.n319 B.n318 585
R529 B.n191 B.n190 585
R530 B.n192 B.n191 585
R531 B.n311 B.n310 585
R532 B.n312 B.n311 585
R533 B.n309 B.n197 585
R534 B.n197 B.n196 585
R535 B.n308 B.n307 585
R536 B.n307 B.n306 585
R537 B.n303 B.n201 585
R538 B.n302 B.n301 585
R539 B.n299 B.n202 585
R540 B.n299 B.n200 585
R541 B.n298 B.n297 585
R542 B.n296 B.n295 585
R543 B.n294 B.n204 585
R544 B.n292 B.n291 585
R545 B.n290 B.n205 585
R546 B.n289 B.n288 585
R547 B.n286 B.n206 585
R548 B.n284 B.n283 585
R549 B.n282 B.n207 585
R550 B.n281 B.n280 585
R551 B.n278 B.n208 585
R552 B.n276 B.n275 585
R553 B.n273 B.n209 585
R554 B.n272 B.n271 585
R555 B.n269 B.n212 585
R556 B.n267 B.n266 585
R557 B.n265 B.n213 585
R558 B.n264 B.n263 585
R559 B.n261 B.n214 585
R560 B.n259 B.n258 585
R561 B.n257 B.n215 585
R562 B.n256 B.n255 585
R563 B.n253 B.n252 585
R564 B.n251 B.n250 585
R565 B.n249 B.n220 585
R566 B.n247 B.n246 585
R567 B.n245 B.n221 585
R568 B.n244 B.n243 585
R569 B.n241 B.n222 585
R570 B.n239 B.n238 585
R571 B.n237 B.n223 585
R572 B.n236 B.n235 585
R573 B.n233 B.n224 585
R574 B.n231 B.n230 585
R575 B.n229 B.n225 585
R576 B.n228 B.n227 585
R577 B.n199 B.n198 585
R578 B.n200 B.n199 585
R579 B.n305 B.n304 585
R580 B.n306 B.n305 585
R581 B.n195 B.n194 585
R582 B.n196 B.n195 585
R583 B.n314 B.n313 585
R584 B.n313 B.n312 585
R585 B.n315 B.n193 585
R586 B.n193 B.n192 585
R587 B.n317 B.n316 585
R588 B.n318 B.n317 585
R589 B.n187 B.n186 585
R590 B.n188 B.n187 585
R591 B.n327 B.n326 585
R592 B.n326 B.n325 585
R593 B.n328 B.n185 585
R594 B.n324 B.n185 585
R595 B.n330 B.n329 585
R596 B.n331 B.n330 585
R597 B.n180 B.n179 585
R598 B.n181 B.n180 585
R599 B.n339 B.n338 585
R600 B.n338 B.n337 585
R601 B.n340 B.n178 585
R602 B.n178 B.n177 585
R603 B.n342 B.n341 585
R604 B.n343 B.n342 585
R605 B.n172 B.n171 585
R606 B.n173 B.n172 585
R607 B.n351 B.n350 585
R608 B.n350 B.n349 585
R609 B.n352 B.n170 585
R610 B.n170 B.n168 585
R611 B.n354 B.n353 585
R612 B.n355 B.n354 585
R613 B.n164 B.n163 585
R614 B.n169 B.n164 585
R615 B.n363 B.n362 585
R616 B.n362 B.n361 585
R617 B.n364 B.n162 585
R618 B.n162 B.n161 585
R619 B.n366 B.n365 585
R620 B.n367 B.n366 585
R621 B.n156 B.n155 585
R622 B.n157 B.n156 585
R623 B.n375 B.n374 585
R624 B.n374 B.n373 585
R625 B.n376 B.n154 585
R626 B.n154 B.n152 585
R627 B.n378 B.n377 585
R628 B.n379 B.n378 585
R629 B.n148 B.n147 585
R630 B.n153 B.n148 585
R631 B.n387 B.n386 585
R632 B.n386 B.n385 585
R633 B.n388 B.n146 585
R634 B.n146 B.n145 585
R635 B.n390 B.n389 585
R636 B.n391 B.n390 585
R637 B.n140 B.n139 585
R638 B.n141 B.n140 585
R639 B.n399 B.n398 585
R640 B.n398 B.n397 585
R641 B.n400 B.n138 585
R642 B.n138 B.n136 585
R643 B.n402 B.n401 585
R644 B.n403 B.n402 585
R645 B.n132 B.n131 585
R646 B.n137 B.n132 585
R647 B.n411 B.n410 585
R648 B.n410 B.n409 585
R649 B.n412 B.n130 585
R650 B.n130 B.n129 585
R651 B.n414 B.n413 585
R652 B.n415 B.n414 585
R653 B.n124 B.n123 585
R654 B.n125 B.n124 585
R655 B.n423 B.n422 585
R656 B.n422 B.n421 585
R657 B.n424 B.n122 585
R658 B.n122 B.n121 585
R659 B.n426 B.n425 585
R660 B.n427 B.n426 585
R661 B.n116 B.n115 585
R662 B.n117 B.n116 585
R663 B.n436 B.n435 585
R664 B.n435 B.n434 585
R665 B.n437 B.n114 585
R666 B.n114 B.n113 585
R667 B.n439 B.n438 585
R668 B.n440 B.n439 585
R669 B.n2 B.n0 585
R670 B.n4 B.n2 585
R671 B.n3 B.n1 585
R672 B.n674 B.n3 585
R673 B.n672 B.n671 585
R674 B.n673 B.n672 585
R675 B.n670 B.n9 585
R676 B.n9 B.n8 585
R677 B.n669 B.n668 585
R678 B.n668 B.n667 585
R679 B.n11 B.n10 585
R680 B.n666 B.n11 585
R681 B.n664 B.n663 585
R682 B.n665 B.n664 585
R683 B.n662 B.n16 585
R684 B.n16 B.n15 585
R685 B.n661 B.n660 585
R686 B.n660 B.n659 585
R687 B.n18 B.n17 585
R688 B.n658 B.n18 585
R689 B.n656 B.n655 585
R690 B.n657 B.n656 585
R691 B.n654 B.n23 585
R692 B.n23 B.n22 585
R693 B.n653 B.n652 585
R694 B.n652 B.n651 585
R695 B.n25 B.n24 585
R696 B.n650 B.n25 585
R697 B.n648 B.n647 585
R698 B.n649 B.n648 585
R699 B.n646 B.n30 585
R700 B.n30 B.n29 585
R701 B.n645 B.n644 585
R702 B.n644 B.n643 585
R703 B.n32 B.n31 585
R704 B.n642 B.n32 585
R705 B.n640 B.n639 585
R706 B.n641 B.n640 585
R707 B.n638 B.n37 585
R708 B.n37 B.n36 585
R709 B.n637 B.n636 585
R710 B.n636 B.n635 585
R711 B.n39 B.n38 585
R712 B.n634 B.n39 585
R713 B.n632 B.n631 585
R714 B.n633 B.n632 585
R715 B.n630 B.n44 585
R716 B.n44 B.n43 585
R717 B.n629 B.n628 585
R718 B.n628 B.n627 585
R719 B.n46 B.n45 585
R720 B.n626 B.n46 585
R721 B.n624 B.n623 585
R722 B.n625 B.n624 585
R723 B.n622 B.n51 585
R724 B.n51 B.n50 585
R725 B.n621 B.n620 585
R726 B.n620 B.n619 585
R727 B.n53 B.n52 585
R728 B.n618 B.n53 585
R729 B.n616 B.n615 585
R730 B.n617 B.n616 585
R731 B.n614 B.n58 585
R732 B.n58 B.n57 585
R733 B.n613 B.n612 585
R734 B.n612 B.n611 585
R735 B.n60 B.n59 585
R736 B.n610 B.n60 585
R737 B.n608 B.n607 585
R738 B.n609 B.n608 585
R739 B.n606 B.n65 585
R740 B.n65 B.n64 585
R741 B.n605 B.n604 585
R742 B.n604 B.n603 585
R743 B.n67 B.n66 585
R744 B.n602 B.n67 585
R745 B.n600 B.n599 585
R746 B.n601 B.n600 585
R747 B.n598 B.n71 585
R748 B.n74 B.n71 585
R749 B.n597 B.n596 585
R750 B.n596 B.n595 585
R751 B.n73 B.n72 585
R752 B.n594 B.n73 585
R753 B.n592 B.n591 585
R754 B.n593 B.n592 585
R755 B.n590 B.n79 585
R756 B.n79 B.n78 585
R757 B.n589 B.n588 585
R758 B.n588 B.n587 585
R759 B.n81 B.n80 585
R760 B.n586 B.n81 585
R761 B.n584 B.n583 585
R762 B.n585 B.n584 585
R763 B.n677 B.n676 585
R764 B.n676 B.n675 585
R765 B.n305 B.n201 526.135
R766 B.n584 B.n86 526.135
R767 B.n307 B.n199 526.135
R768 B.n503 B.n84 526.135
R769 B.n504 B.n85 256.663
R770 B.n506 B.n85 256.663
R771 B.n512 B.n85 256.663
R772 B.n514 B.n85 256.663
R773 B.n520 B.n85 256.663
R774 B.n522 B.n85 256.663
R775 B.n528 B.n85 256.663
R776 B.n530 B.n85 256.663
R777 B.n537 B.n85 256.663
R778 B.n539 B.n85 256.663
R779 B.n545 B.n85 256.663
R780 B.n547 B.n85 256.663
R781 B.n553 B.n85 256.663
R782 B.n555 B.n85 256.663
R783 B.n561 B.n85 256.663
R784 B.n563 B.n85 256.663
R785 B.n569 B.n85 256.663
R786 B.n571 B.n85 256.663
R787 B.n577 B.n85 256.663
R788 B.n579 B.n85 256.663
R789 B.n300 B.n200 256.663
R790 B.n203 B.n200 256.663
R791 B.n293 B.n200 256.663
R792 B.n287 B.n200 256.663
R793 B.n285 B.n200 256.663
R794 B.n279 B.n200 256.663
R795 B.n277 B.n200 256.663
R796 B.n270 B.n200 256.663
R797 B.n268 B.n200 256.663
R798 B.n262 B.n200 256.663
R799 B.n260 B.n200 256.663
R800 B.n254 B.n200 256.663
R801 B.n219 B.n200 256.663
R802 B.n248 B.n200 256.663
R803 B.n242 B.n200 256.663
R804 B.n240 B.n200 256.663
R805 B.n234 B.n200 256.663
R806 B.n232 B.n200 256.663
R807 B.n226 B.n200 256.663
R808 B.n216 B.t15 240.891
R809 B.n210 B.t19 240.891
R810 B.n95 B.t8 240.891
R811 B.n102 B.t12 240.891
R812 B.n216 B.t18 180.276
R813 B.n102 B.t13 180.276
R814 B.n210 B.t21 180.276
R815 B.n95 B.t10 180.276
R816 B.n305 B.n195 163.367
R817 B.n313 B.n195 163.367
R818 B.n313 B.n193 163.367
R819 B.n317 B.n193 163.367
R820 B.n317 B.n187 163.367
R821 B.n326 B.n187 163.367
R822 B.n326 B.n185 163.367
R823 B.n330 B.n185 163.367
R824 B.n330 B.n180 163.367
R825 B.n338 B.n180 163.367
R826 B.n338 B.n178 163.367
R827 B.n342 B.n178 163.367
R828 B.n342 B.n172 163.367
R829 B.n350 B.n172 163.367
R830 B.n350 B.n170 163.367
R831 B.n354 B.n170 163.367
R832 B.n354 B.n164 163.367
R833 B.n362 B.n164 163.367
R834 B.n362 B.n162 163.367
R835 B.n366 B.n162 163.367
R836 B.n366 B.n156 163.367
R837 B.n374 B.n156 163.367
R838 B.n374 B.n154 163.367
R839 B.n378 B.n154 163.367
R840 B.n378 B.n148 163.367
R841 B.n386 B.n148 163.367
R842 B.n386 B.n146 163.367
R843 B.n390 B.n146 163.367
R844 B.n390 B.n140 163.367
R845 B.n398 B.n140 163.367
R846 B.n398 B.n138 163.367
R847 B.n402 B.n138 163.367
R848 B.n402 B.n132 163.367
R849 B.n410 B.n132 163.367
R850 B.n410 B.n130 163.367
R851 B.n414 B.n130 163.367
R852 B.n414 B.n124 163.367
R853 B.n422 B.n124 163.367
R854 B.n422 B.n122 163.367
R855 B.n426 B.n122 163.367
R856 B.n426 B.n116 163.367
R857 B.n435 B.n116 163.367
R858 B.n435 B.n114 163.367
R859 B.n439 B.n114 163.367
R860 B.n439 B.n2 163.367
R861 B.n676 B.n2 163.367
R862 B.n676 B.n3 163.367
R863 B.n672 B.n3 163.367
R864 B.n672 B.n9 163.367
R865 B.n668 B.n9 163.367
R866 B.n668 B.n11 163.367
R867 B.n664 B.n11 163.367
R868 B.n664 B.n16 163.367
R869 B.n660 B.n16 163.367
R870 B.n660 B.n18 163.367
R871 B.n656 B.n18 163.367
R872 B.n656 B.n23 163.367
R873 B.n652 B.n23 163.367
R874 B.n652 B.n25 163.367
R875 B.n648 B.n25 163.367
R876 B.n648 B.n30 163.367
R877 B.n644 B.n30 163.367
R878 B.n644 B.n32 163.367
R879 B.n640 B.n32 163.367
R880 B.n640 B.n37 163.367
R881 B.n636 B.n37 163.367
R882 B.n636 B.n39 163.367
R883 B.n632 B.n39 163.367
R884 B.n632 B.n44 163.367
R885 B.n628 B.n44 163.367
R886 B.n628 B.n46 163.367
R887 B.n624 B.n46 163.367
R888 B.n624 B.n51 163.367
R889 B.n620 B.n51 163.367
R890 B.n620 B.n53 163.367
R891 B.n616 B.n53 163.367
R892 B.n616 B.n58 163.367
R893 B.n612 B.n58 163.367
R894 B.n612 B.n60 163.367
R895 B.n608 B.n60 163.367
R896 B.n608 B.n65 163.367
R897 B.n604 B.n65 163.367
R898 B.n604 B.n67 163.367
R899 B.n600 B.n67 163.367
R900 B.n600 B.n71 163.367
R901 B.n596 B.n71 163.367
R902 B.n596 B.n73 163.367
R903 B.n592 B.n73 163.367
R904 B.n592 B.n79 163.367
R905 B.n588 B.n79 163.367
R906 B.n588 B.n81 163.367
R907 B.n584 B.n81 163.367
R908 B.n301 B.n299 163.367
R909 B.n299 B.n298 163.367
R910 B.n295 B.n294 163.367
R911 B.n292 B.n205 163.367
R912 B.n288 B.n286 163.367
R913 B.n284 B.n207 163.367
R914 B.n280 B.n278 163.367
R915 B.n276 B.n209 163.367
R916 B.n271 B.n269 163.367
R917 B.n267 B.n213 163.367
R918 B.n263 B.n261 163.367
R919 B.n259 B.n215 163.367
R920 B.n255 B.n253 163.367
R921 B.n250 B.n249 163.367
R922 B.n247 B.n221 163.367
R923 B.n243 B.n241 163.367
R924 B.n239 B.n223 163.367
R925 B.n235 B.n233 163.367
R926 B.n231 B.n225 163.367
R927 B.n227 B.n199 163.367
R928 B.n307 B.n197 163.367
R929 B.n311 B.n197 163.367
R930 B.n311 B.n191 163.367
R931 B.n319 B.n191 163.367
R932 B.n319 B.n189 163.367
R933 B.n323 B.n189 163.367
R934 B.n323 B.n184 163.367
R935 B.n332 B.n184 163.367
R936 B.n332 B.n182 163.367
R937 B.n336 B.n182 163.367
R938 B.n336 B.n176 163.367
R939 B.n344 B.n176 163.367
R940 B.n344 B.n174 163.367
R941 B.n348 B.n174 163.367
R942 B.n348 B.n167 163.367
R943 B.n356 B.n167 163.367
R944 B.n356 B.n165 163.367
R945 B.n360 B.n165 163.367
R946 B.n360 B.n160 163.367
R947 B.n368 B.n160 163.367
R948 B.n368 B.n158 163.367
R949 B.n372 B.n158 163.367
R950 B.n372 B.n151 163.367
R951 B.n380 B.n151 163.367
R952 B.n380 B.n149 163.367
R953 B.n384 B.n149 163.367
R954 B.n384 B.n144 163.367
R955 B.n392 B.n144 163.367
R956 B.n392 B.n142 163.367
R957 B.n396 B.n142 163.367
R958 B.n396 B.n135 163.367
R959 B.n404 B.n135 163.367
R960 B.n404 B.n133 163.367
R961 B.n408 B.n133 163.367
R962 B.n408 B.n128 163.367
R963 B.n416 B.n128 163.367
R964 B.n416 B.n126 163.367
R965 B.n420 B.n126 163.367
R966 B.n420 B.n120 163.367
R967 B.n428 B.n120 163.367
R968 B.n428 B.n118 163.367
R969 B.n433 B.n118 163.367
R970 B.n433 B.n112 163.367
R971 B.n441 B.n112 163.367
R972 B.n442 B.n441 163.367
R973 B.n442 B.n5 163.367
R974 B.n6 B.n5 163.367
R975 B.n7 B.n6 163.367
R976 B.n447 B.n7 163.367
R977 B.n447 B.n12 163.367
R978 B.n13 B.n12 163.367
R979 B.n14 B.n13 163.367
R980 B.n452 B.n14 163.367
R981 B.n452 B.n19 163.367
R982 B.n20 B.n19 163.367
R983 B.n21 B.n20 163.367
R984 B.n457 B.n21 163.367
R985 B.n457 B.n26 163.367
R986 B.n27 B.n26 163.367
R987 B.n28 B.n27 163.367
R988 B.n462 B.n28 163.367
R989 B.n462 B.n33 163.367
R990 B.n34 B.n33 163.367
R991 B.n35 B.n34 163.367
R992 B.n467 B.n35 163.367
R993 B.n467 B.n40 163.367
R994 B.n41 B.n40 163.367
R995 B.n42 B.n41 163.367
R996 B.n472 B.n42 163.367
R997 B.n472 B.n47 163.367
R998 B.n48 B.n47 163.367
R999 B.n49 B.n48 163.367
R1000 B.n477 B.n49 163.367
R1001 B.n477 B.n54 163.367
R1002 B.n55 B.n54 163.367
R1003 B.n56 B.n55 163.367
R1004 B.n482 B.n56 163.367
R1005 B.n482 B.n61 163.367
R1006 B.n62 B.n61 163.367
R1007 B.n63 B.n62 163.367
R1008 B.n487 B.n63 163.367
R1009 B.n487 B.n68 163.367
R1010 B.n69 B.n68 163.367
R1011 B.n70 B.n69 163.367
R1012 B.n492 B.n70 163.367
R1013 B.n492 B.n75 163.367
R1014 B.n76 B.n75 163.367
R1015 B.n77 B.n76 163.367
R1016 B.n497 B.n77 163.367
R1017 B.n497 B.n82 163.367
R1018 B.n83 B.n82 163.367
R1019 B.n84 B.n83 163.367
R1020 B.n580 B.n578 163.367
R1021 B.n576 B.n88 163.367
R1022 B.n572 B.n570 163.367
R1023 B.n568 B.n90 163.367
R1024 B.n564 B.n562 163.367
R1025 B.n560 B.n92 163.367
R1026 B.n556 B.n554 163.367
R1027 B.n552 B.n94 163.367
R1028 B.n548 B.n546 163.367
R1029 B.n544 B.n99 163.367
R1030 B.n540 B.n538 163.367
R1031 B.n536 B.n101 163.367
R1032 B.n531 B.n529 163.367
R1033 B.n527 B.n105 163.367
R1034 B.n523 B.n521 163.367
R1035 B.n519 B.n107 163.367
R1036 B.n515 B.n513 163.367
R1037 B.n511 B.n109 163.367
R1038 B.n507 B.n505 163.367
R1039 B.n306 B.n200 153.488
R1040 B.n585 B.n85 153.488
R1041 B.n217 B.t17 130.434
R1042 B.n103 B.t14 130.434
R1043 B.n211 B.t20 130.434
R1044 B.n96 B.t11 130.434
R1045 B.n306 B.n196 89.2074
R1046 B.n312 B.n196 89.2074
R1047 B.n312 B.n192 89.2074
R1048 B.n318 B.n192 89.2074
R1049 B.n318 B.n188 89.2074
R1050 B.n325 B.n188 89.2074
R1051 B.n325 B.n324 89.2074
R1052 B.n331 B.n181 89.2074
R1053 B.n337 B.n181 89.2074
R1054 B.n337 B.n177 89.2074
R1055 B.n343 B.n177 89.2074
R1056 B.n343 B.n173 89.2074
R1057 B.n349 B.n173 89.2074
R1058 B.n349 B.n168 89.2074
R1059 B.n355 B.n168 89.2074
R1060 B.n355 B.n169 89.2074
R1061 B.n361 B.n161 89.2074
R1062 B.n367 B.n161 89.2074
R1063 B.n367 B.n157 89.2074
R1064 B.n373 B.n157 89.2074
R1065 B.n373 B.n152 89.2074
R1066 B.n379 B.n152 89.2074
R1067 B.n379 B.n153 89.2074
R1068 B.n385 B.n145 89.2074
R1069 B.n391 B.n145 89.2074
R1070 B.n391 B.n141 89.2074
R1071 B.n397 B.n141 89.2074
R1072 B.n397 B.n136 89.2074
R1073 B.n403 B.n136 89.2074
R1074 B.n403 B.n137 89.2074
R1075 B.n409 B.n129 89.2074
R1076 B.n415 B.n129 89.2074
R1077 B.n415 B.n125 89.2074
R1078 B.n421 B.n125 89.2074
R1079 B.n421 B.n121 89.2074
R1080 B.n427 B.n121 89.2074
R1081 B.n434 B.n117 89.2074
R1082 B.n434 B.n113 89.2074
R1083 B.n440 B.n113 89.2074
R1084 B.n440 B.n4 89.2074
R1085 B.n675 B.n4 89.2074
R1086 B.n675 B.n674 89.2074
R1087 B.n674 B.n673 89.2074
R1088 B.n673 B.n8 89.2074
R1089 B.n667 B.n8 89.2074
R1090 B.n667 B.n666 89.2074
R1091 B.n665 B.n15 89.2074
R1092 B.n659 B.n15 89.2074
R1093 B.n659 B.n658 89.2074
R1094 B.n658 B.n657 89.2074
R1095 B.n657 B.n22 89.2074
R1096 B.n651 B.n22 89.2074
R1097 B.n650 B.n649 89.2074
R1098 B.n649 B.n29 89.2074
R1099 B.n643 B.n29 89.2074
R1100 B.n643 B.n642 89.2074
R1101 B.n642 B.n641 89.2074
R1102 B.n641 B.n36 89.2074
R1103 B.n635 B.n36 89.2074
R1104 B.n634 B.n633 89.2074
R1105 B.n633 B.n43 89.2074
R1106 B.n627 B.n43 89.2074
R1107 B.n627 B.n626 89.2074
R1108 B.n626 B.n625 89.2074
R1109 B.n625 B.n50 89.2074
R1110 B.n619 B.n50 89.2074
R1111 B.n618 B.n617 89.2074
R1112 B.n617 B.n57 89.2074
R1113 B.n611 B.n57 89.2074
R1114 B.n611 B.n610 89.2074
R1115 B.n610 B.n609 89.2074
R1116 B.n609 B.n64 89.2074
R1117 B.n603 B.n64 89.2074
R1118 B.n603 B.n602 89.2074
R1119 B.n602 B.n601 89.2074
R1120 B.n595 B.n74 89.2074
R1121 B.n595 B.n594 89.2074
R1122 B.n594 B.n593 89.2074
R1123 B.n593 B.n78 89.2074
R1124 B.n587 B.n78 89.2074
R1125 B.n587 B.n586 89.2074
R1126 B.n586 B.n585 89.2074
R1127 B.n169 B.t7 83.9599
R1128 B.n409 B.t1 83.9599
R1129 B.n651 B.t3 83.9599
R1130 B.t6 B.n618 83.9599
R1131 B.n331 B.t16 73.465
R1132 B.n601 B.t9 73.465
R1133 B.n300 B.n201 71.676
R1134 B.n298 B.n203 71.676
R1135 B.n294 B.n293 71.676
R1136 B.n287 B.n205 71.676
R1137 B.n286 B.n285 71.676
R1138 B.n279 B.n207 71.676
R1139 B.n278 B.n277 71.676
R1140 B.n270 B.n209 71.676
R1141 B.n269 B.n268 71.676
R1142 B.n262 B.n213 71.676
R1143 B.n261 B.n260 71.676
R1144 B.n254 B.n215 71.676
R1145 B.n253 B.n219 71.676
R1146 B.n249 B.n248 71.676
R1147 B.n242 B.n221 71.676
R1148 B.n241 B.n240 71.676
R1149 B.n234 B.n223 71.676
R1150 B.n233 B.n232 71.676
R1151 B.n226 B.n225 71.676
R1152 B.n579 B.n86 71.676
R1153 B.n578 B.n577 71.676
R1154 B.n571 B.n88 71.676
R1155 B.n570 B.n569 71.676
R1156 B.n563 B.n90 71.676
R1157 B.n562 B.n561 71.676
R1158 B.n555 B.n92 71.676
R1159 B.n554 B.n553 71.676
R1160 B.n547 B.n94 71.676
R1161 B.n546 B.n545 71.676
R1162 B.n539 B.n99 71.676
R1163 B.n538 B.n537 71.676
R1164 B.n530 B.n101 71.676
R1165 B.n529 B.n528 71.676
R1166 B.n522 B.n105 71.676
R1167 B.n521 B.n520 71.676
R1168 B.n514 B.n107 71.676
R1169 B.n513 B.n512 71.676
R1170 B.n506 B.n109 71.676
R1171 B.n505 B.n504 71.676
R1172 B.n504 B.n503 71.676
R1173 B.n507 B.n506 71.676
R1174 B.n512 B.n511 71.676
R1175 B.n515 B.n514 71.676
R1176 B.n520 B.n519 71.676
R1177 B.n523 B.n522 71.676
R1178 B.n528 B.n527 71.676
R1179 B.n531 B.n530 71.676
R1180 B.n537 B.n536 71.676
R1181 B.n540 B.n539 71.676
R1182 B.n545 B.n544 71.676
R1183 B.n548 B.n547 71.676
R1184 B.n553 B.n552 71.676
R1185 B.n556 B.n555 71.676
R1186 B.n561 B.n560 71.676
R1187 B.n564 B.n563 71.676
R1188 B.n569 B.n568 71.676
R1189 B.n572 B.n571 71.676
R1190 B.n577 B.n576 71.676
R1191 B.n580 B.n579 71.676
R1192 B.n301 B.n300 71.676
R1193 B.n295 B.n203 71.676
R1194 B.n293 B.n292 71.676
R1195 B.n288 B.n287 71.676
R1196 B.n285 B.n284 71.676
R1197 B.n280 B.n279 71.676
R1198 B.n277 B.n276 71.676
R1199 B.n271 B.n270 71.676
R1200 B.n268 B.n267 71.676
R1201 B.n263 B.n262 71.676
R1202 B.n260 B.n259 71.676
R1203 B.n255 B.n254 71.676
R1204 B.n250 B.n219 71.676
R1205 B.n248 B.n247 71.676
R1206 B.n243 B.n242 71.676
R1207 B.n240 B.n239 71.676
R1208 B.n235 B.n234 71.676
R1209 B.n232 B.n231 71.676
R1210 B.n227 B.n226 71.676
R1211 B.n218 B.n217 59.5399
R1212 B.n274 B.n211 59.5399
R1213 B.n97 B.n96 59.5399
R1214 B.n533 B.n103 59.5399
R1215 B.n427 B.t2 55.0989
R1216 B.t5 B.n665 55.0989
R1217 B.n217 B.n216 49.8429
R1218 B.n211 B.n210 49.8429
R1219 B.n96 B.n95 49.8429
R1220 B.n103 B.n102 49.8429
R1221 B.n153 B.t0 44.604
R1222 B.n385 B.t0 44.604
R1223 B.n635 B.t4 44.604
R1224 B.t4 B.n634 44.604
R1225 B.n583 B.n582 34.1859
R1226 B.n502 B.n501 34.1859
R1227 B.n308 B.n198 34.1859
R1228 B.n304 B.n303 34.1859
R1229 B.t2 B.n117 34.109
R1230 B.n666 B.t5 34.109
R1231 B B.n677 18.0485
R1232 B.n324 B.t16 15.7429
R1233 B.n74 B.t9 15.7429
R1234 B.n582 B.n581 10.6151
R1235 B.n581 B.n87 10.6151
R1236 B.n575 B.n87 10.6151
R1237 B.n575 B.n574 10.6151
R1238 B.n574 B.n573 10.6151
R1239 B.n573 B.n89 10.6151
R1240 B.n567 B.n89 10.6151
R1241 B.n567 B.n566 10.6151
R1242 B.n566 B.n565 10.6151
R1243 B.n565 B.n91 10.6151
R1244 B.n559 B.n91 10.6151
R1245 B.n559 B.n558 10.6151
R1246 B.n558 B.n557 10.6151
R1247 B.n557 B.n93 10.6151
R1248 B.n551 B.n550 10.6151
R1249 B.n550 B.n549 10.6151
R1250 B.n549 B.n98 10.6151
R1251 B.n543 B.n98 10.6151
R1252 B.n543 B.n542 10.6151
R1253 B.n542 B.n541 10.6151
R1254 B.n541 B.n100 10.6151
R1255 B.n535 B.n100 10.6151
R1256 B.n535 B.n534 10.6151
R1257 B.n532 B.n104 10.6151
R1258 B.n526 B.n104 10.6151
R1259 B.n526 B.n525 10.6151
R1260 B.n525 B.n524 10.6151
R1261 B.n524 B.n106 10.6151
R1262 B.n518 B.n106 10.6151
R1263 B.n518 B.n517 10.6151
R1264 B.n517 B.n516 10.6151
R1265 B.n516 B.n108 10.6151
R1266 B.n510 B.n108 10.6151
R1267 B.n510 B.n509 10.6151
R1268 B.n509 B.n508 10.6151
R1269 B.n508 B.n110 10.6151
R1270 B.n502 B.n110 10.6151
R1271 B.n309 B.n308 10.6151
R1272 B.n310 B.n309 10.6151
R1273 B.n310 B.n190 10.6151
R1274 B.n320 B.n190 10.6151
R1275 B.n321 B.n320 10.6151
R1276 B.n322 B.n321 10.6151
R1277 B.n322 B.n183 10.6151
R1278 B.n333 B.n183 10.6151
R1279 B.n334 B.n333 10.6151
R1280 B.n335 B.n334 10.6151
R1281 B.n335 B.n175 10.6151
R1282 B.n345 B.n175 10.6151
R1283 B.n346 B.n345 10.6151
R1284 B.n347 B.n346 10.6151
R1285 B.n347 B.n166 10.6151
R1286 B.n357 B.n166 10.6151
R1287 B.n358 B.n357 10.6151
R1288 B.n359 B.n358 10.6151
R1289 B.n359 B.n159 10.6151
R1290 B.n369 B.n159 10.6151
R1291 B.n370 B.n369 10.6151
R1292 B.n371 B.n370 10.6151
R1293 B.n371 B.n150 10.6151
R1294 B.n381 B.n150 10.6151
R1295 B.n382 B.n381 10.6151
R1296 B.n383 B.n382 10.6151
R1297 B.n383 B.n143 10.6151
R1298 B.n393 B.n143 10.6151
R1299 B.n394 B.n393 10.6151
R1300 B.n395 B.n394 10.6151
R1301 B.n395 B.n134 10.6151
R1302 B.n405 B.n134 10.6151
R1303 B.n406 B.n405 10.6151
R1304 B.n407 B.n406 10.6151
R1305 B.n407 B.n127 10.6151
R1306 B.n417 B.n127 10.6151
R1307 B.n418 B.n417 10.6151
R1308 B.n419 B.n418 10.6151
R1309 B.n419 B.n119 10.6151
R1310 B.n429 B.n119 10.6151
R1311 B.n430 B.n429 10.6151
R1312 B.n432 B.n430 10.6151
R1313 B.n432 B.n431 10.6151
R1314 B.n431 B.n111 10.6151
R1315 B.n443 B.n111 10.6151
R1316 B.n444 B.n443 10.6151
R1317 B.n445 B.n444 10.6151
R1318 B.n446 B.n445 10.6151
R1319 B.n448 B.n446 10.6151
R1320 B.n449 B.n448 10.6151
R1321 B.n450 B.n449 10.6151
R1322 B.n451 B.n450 10.6151
R1323 B.n453 B.n451 10.6151
R1324 B.n454 B.n453 10.6151
R1325 B.n455 B.n454 10.6151
R1326 B.n456 B.n455 10.6151
R1327 B.n458 B.n456 10.6151
R1328 B.n459 B.n458 10.6151
R1329 B.n460 B.n459 10.6151
R1330 B.n461 B.n460 10.6151
R1331 B.n463 B.n461 10.6151
R1332 B.n464 B.n463 10.6151
R1333 B.n465 B.n464 10.6151
R1334 B.n466 B.n465 10.6151
R1335 B.n468 B.n466 10.6151
R1336 B.n469 B.n468 10.6151
R1337 B.n470 B.n469 10.6151
R1338 B.n471 B.n470 10.6151
R1339 B.n473 B.n471 10.6151
R1340 B.n474 B.n473 10.6151
R1341 B.n475 B.n474 10.6151
R1342 B.n476 B.n475 10.6151
R1343 B.n478 B.n476 10.6151
R1344 B.n479 B.n478 10.6151
R1345 B.n480 B.n479 10.6151
R1346 B.n481 B.n480 10.6151
R1347 B.n483 B.n481 10.6151
R1348 B.n484 B.n483 10.6151
R1349 B.n485 B.n484 10.6151
R1350 B.n486 B.n485 10.6151
R1351 B.n488 B.n486 10.6151
R1352 B.n489 B.n488 10.6151
R1353 B.n490 B.n489 10.6151
R1354 B.n491 B.n490 10.6151
R1355 B.n493 B.n491 10.6151
R1356 B.n494 B.n493 10.6151
R1357 B.n495 B.n494 10.6151
R1358 B.n496 B.n495 10.6151
R1359 B.n498 B.n496 10.6151
R1360 B.n499 B.n498 10.6151
R1361 B.n500 B.n499 10.6151
R1362 B.n501 B.n500 10.6151
R1363 B.n303 B.n302 10.6151
R1364 B.n302 B.n202 10.6151
R1365 B.n297 B.n202 10.6151
R1366 B.n297 B.n296 10.6151
R1367 B.n296 B.n204 10.6151
R1368 B.n291 B.n204 10.6151
R1369 B.n291 B.n290 10.6151
R1370 B.n290 B.n289 10.6151
R1371 B.n289 B.n206 10.6151
R1372 B.n283 B.n206 10.6151
R1373 B.n283 B.n282 10.6151
R1374 B.n282 B.n281 10.6151
R1375 B.n281 B.n208 10.6151
R1376 B.n275 B.n208 10.6151
R1377 B.n273 B.n272 10.6151
R1378 B.n272 B.n212 10.6151
R1379 B.n266 B.n212 10.6151
R1380 B.n266 B.n265 10.6151
R1381 B.n265 B.n264 10.6151
R1382 B.n264 B.n214 10.6151
R1383 B.n258 B.n214 10.6151
R1384 B.n258 B.n257 10.6151
R1385 B.n257 B.n256 10.6151
R1386 B.n252 B.n251 10.6151
R1387 B.n251 B.n220 10.6151
R1388 B.n246 B.n220 10.6151
R1389 B.n246 B.n245 10.6151
R1390 B.n245 B.n244 10.6151
R1391 B.n244 B.n222 10.6151
R1392 B.n238 B.n222 10.6151
R1393 B.n238 B.n237 10.6151
R1394 B.n237 B.n236 10.6151
R1395 B.n236 B.n224 10.6151
R1396 B.n230 B.n224 10.6151
R1397 B.n230 B.n229 10.6151
R1398 B.n229 B.n228 10.6151
R1399 B.n228 B.n198 10.6151
R1400 B.n304 B.n194 10.6151
R1401 B.n314 B.n194 10.6151
R1402 B.n315 B.n314 10.6151
R1403 B.n316 B.n315 10.6151
R1404 B.n316 B.n186 10.6151
R1405 B.n327 B.n186 10.6151
R1406 B.n328 B.n327 10.6151
R1407 B.n329 B.n328 10.6151
R1408 B.n329 B.n179 10.6151
R1409 B.n339 B.n179 10.6151
R1410 B.n340 B.n339 10.6151
R1411 B.n341 B.n340 10.6151
R1412 B.n341 B.n171 10.6151
R1413 B.n351 B.n171 10.6151
R1414 B.n352 B.n351 10.6151
R1415 B.n353 B.n352 10.6151
R1416 B.n353 B.n163 10.6151
R1417 B.n363 B.n163 10.6151
R1418 B.n364 B.n363 10.6151
R1419 B.n365 B.n364 10.6151
R1420 B.n365 B.n155 10.6151
R1421 B.n375 B.n155 10.6151
R1422 B.n376 B.n375 10.6151
R1423 B.n377 B.n376 10.6151
R1424 B.n377 B.n147 10.6151
R1425 B.n387 B.n147 10.6151
R1426 B.n388 B.n387 10.6151
R1427 B.n389 B.n388 10.6151
R1428 B.n389 B.n139 10.6151
R1429 B.n399 B.n139 10.6151
R1430 B.n400 B.n399 10.6151
R1431 B.n401 B.n400 10.6151
R1432 B.n401 B.n131 10.6151
R1433 B.n411 B.n131 10.6151
R1434 B.n412 B.n411 10.6151
R1435 B.n413 B.n412 10.6151
R1436 B.n413 B.n123 10.6151
R1437 B.n423 B.n123 10.6151
R1438 B.n424 B.n423 10.6151
R1439 B.n425 B.n424 10.6151
R1440 B.n425 B.n115 10.6151
R1441 B.n436 B.n115 10.6151
R1442 B.n437 B.n436 10.6151
R1443 B.n438 B.n437 10.6151
R1444 B.n438 B.n0 10.6151
R1445 B.n671 B.n1 10.6151
R1446 B.n671 B.n670 10.6151
R1447 B.n670 B.n669 10.6151
R1448 B.n669 B.n10 10.6151
R1449 B.n663 B.n10 10.6151
R1450 B.n663 B.n662 10.6151
R1451 B.n662 B.n661 10.6151
R1452 B.n661 B.n17 10.6151
R1453 B.n655 B.n17 10.6151
R1454 B.n655 B.n654 10.6151
R1455 B.n654 B.n653 10.6151
R1456 B.n653 B.n24 10.6151
R1457 B.n647 B.n24 10.6151
R1458 B.n647 B.n646 10.6151
R1459 B.n646 B.n645 10.6151
R1460 B.n645 B.n31 10.6151
R1461 B.n639 B.n31 10.6151
R1462 B.n639 B.n638 10.6151
R1463 B.n638 B.n637 10.6151
R1464 B.n637 B.n38 10.6151
R1465 B.n631 B.n38 10.6151
R1466 B.n631 B.n630 10.6151
R1467 B.n630 B.n629 10.6151
R1468 B.n629 B.n45 10.6151
R1469 B.n623 B.n45 10.6151
R1470 B.n623 B.n622 10.6151
R1471 B.n622 B.n621 10.6151
R1472 B.n621 B.n52 10.6151
R1473 B.n615 B.n52 10.6151
R1474 B.n615 B.n614 10.6151
R1475 B.n614 B.n613 10.6151
R1476 B.n613 B.n59 10.6151
R1477 B.n607 B.n59 10.6151
R1478 B.n607 B.n606 10.6151
R1479 B.n606 B.n605 10.6151
R1480 B.n605 B.n66 10.6151
R1481 B.n599 B.n66 10.6151
R1482 B.n599 B.n598 10.6151
R1483 B.n598 B.n597 10.6151
R1484 B.n597 B.n72 10.6151
R1485 B.n591 B.n72 10.6151
R1486 B.n591 B.n590 10.6151
R1487 B.n590 B.n589 10.6151
R1488 B.n589 B.n80 10.6151
R1489 B.n583 B.n80 10.6151
R1490 B.n97 B.n93 9.36635
R1491 B.n533 B.n532 9.36635
R1492 B.n275 B.n274 9.36635
R1493 B.n252 B.n218 9.36635
R1494 B.n361 B.t7 5.24797
R1495 B.n137 B.t1 5.24797
R1496 B.t3 B.n650 5.24797
R1497 B.n619 B.t6 5.24797
R1498 B.n677 B.n0 2.81026
R1499 B.n677 B.n1 2.81026
R1500 B.n551 B.n97 1.24928
R1501 B.n534 B.n533 1.24928
R1502 B.n274 B.n273 1.24928
R1503 B.n256 B.n218 1.24928
R1504 VP.n16 VP.n15 161.3
R1505 VP.n17 VP.n12 161.3
R1506 VP.n19 VP.n18 161.3
R1507 VP.n20 VP.n11 161.3
R1508 VP.n22 VP.n21 161.3
R1509 VP.n24 VP.n10 161.3
R1510 VP.n26 VP.n25 161.3
R1511 VP.n27 VP.n9 161.3
R1512 VP.n29 VP.n28 161.3
R1513 VP.n30 VP.n8 161.3
R1514 VP.n58 VP.n0 161.3
R1515 VP.n57 VP.n56 161.3
R1516 VP.n55 VP.n1 161.3
R1517 VP.n54 VP.n53 161.3
R1518 VP.n52 VP.n2 161.3
R1519 VP.n50 VP.n49 161.3
R1520 VP.n48 VP.n3 161.3
R1521 VP.n47 VP.n46 161.3
R1522 VP.n45 VP.n4 161.3
R1523 VP.n44 VP.n43 161.3
R1524 VP.n42 VP.n41 161.3
R1525 VP.n40 VP.n6 161.3
R1526 VP.n39 VP.n38 161.3
R1527 VP.n37 VP.n7 161.3
R1528 VP.n36 VP.n35 161.3
R1529 VP.n34 VP.n33 93.3849
R1530 VP.n60 VP.n59 93.3849
R1531 VP.n32 VP.n31 93.3849
R1532 VP.n14 VP.t4 66.8891
R1533 VP.n14 VP.n13 57.3618
R1534 VP.n39 VP.n7 47.2923
R1535 VP.n57 VP.n1 47.2923
R1536 VP.n29 VP.n9 47.2923
R1537 VP.n33 VP.n32 42.5223
R1538 VP.n46 VP.n45 40.4934
R1539 VP.n46 VP.n3 40.4934
R1540 VP.n18 VP.n11 40.4934
R1541 VP.n18 VP.n17 40.4934
R1542 VP.n40 VP.n39 33.6945
R1543 VP.n53 VP.n1 33.6945
R1544 VP.n25 VP.n9 33.6945
R1545 VP.n34 VP.t0 33.4608
R1546 VP.n5 VP.t7 33.4608
R1547 VP.n51 VP.t2 33.4608
R1548 VP.n59 VP.t1 33.4608
R1549 VP.n31 VP.t3 33.4608
R1550 VP.n23 VP.t5 33.4608
R1551 VP.n13 VP.t6 33.4608
R1552 VP.n35 VP.n7 24.4675
R1553 VP.n41 VP.n40 24.4675
R1554 VP.n45 VP.n44 24.4675
R1555 VP.n50 VP.n3 24.4675
R1556 VP.n53 VP.n52 24.4675
R1557 VP.n58 VP.n57 24.4675
R1558 VP.n30 VP.n29 24.4675
R1559 VP.n22 VP.n11 24.4675
R1560 VP.n25 VP.n24 24.4675
R1561 VP.n17 VP.n16 24.4675
R1562 VP.n35 VP.n34 17.3721
R1563 VP.n59 VP.n58 17.3721
R1564 VP.n31 VP.n30 17.3721
R1565 VP.n44 VP.n5 13.9467
R1566 VP.n51 VP.n50 13.9467
R1567 VP.n23 VP.n22 13.9467
R1568 VP.n16 VP.n13 13.9467
R1569 VP.n41 VP.n5 10.5213
R1570 VP.n52 VP.n51 10.5213
R1571 VP.n24 VP.n23 10.5213
R1572 VP.n15 VP.n14 9.22138
R1573 VP.n32 VP.n8 0.278367
R1574 VP.n36 VP.n33 0.278367
R1575 VP.n60 VP.n0 0.278367
R1576 VP.n15 VP.n12 0.189894
R1577 VP.n19 VP.n12 0.189894
R1578 VP.n20 VP.n19 0.189894
R1579 VP.n21 VP.n20 0.189894
R1580 VP.n21 VP.n10 0.189894
R1581 VP.n26 VP.n10 0.189894
R1582 VP.n27 VP.n26 0.189894
R1583 VP.n28 VP.n27 0.189894
R1584 VP.n28 VP.n8 0.189894
R1585 VP.n37 VP.n36 0.189894
R1586 VP.n38 VP.n37 0.189894
R1587 VP.n38 VP.n6 0.189894
R1588 VP.n42 VP.n6 0.189894
R1589 VP.n43 VP.n42 0.189894
R1590 VP.n43 VP.n4 0.189894
R1591 VP.n47 VP.n4 0.189894
R1592 VP.n48 VP.n47 0.189894
R1593 VP.n49 VP.n48 0.189894
R1594 VP.n49 VP.n2 0.189894
R1595 VP.n54 VP.n2 0.189894
R1596 VP.n55 VP.n54 0.189894
R1597 VP.n56 VP.n55 0.189894
R1598 VP.n56 VP.n0 0.189894
R1599 VP VP.n60 0.153454
R1600 VDD1 VDD1.n0 78.7212
R1601 VDD1.n3 VDD1.n2 78.6075
R1602 VDD1.n3 VDD1.n1 78.6075
R1603 VDD1.n5 VDD1.n4 77.5551
R1604 VDD1.n5 VDD1.n3 36.9492
R1605 VDD1.n4 VDD1.t2 6.36706
R1606 VDD1.n4 VDD1.t4 6.36706
R1607 VDD1.n0 VDD1.t3 6.36706
R1608 VDD1.n0 VDD1.t1 6.36706
R1609 VDD1.n2 VDD1.t5 6.36706
R1610 VDD1.n2 VDD1.t6 6.36706
R1611 VDD1.n1 VDD1.t7 6.36706
R1612 VDD1.n1 VDD1.t0 6.36706
R1613 VDD1 VDD1.n5 1.05007
C0 VN VTAIL 3.38487f
C1 VDD2 VTAIL 4.85936f
C2 VDD1 VTAIL 4.80735f
C3 VN VP 5.58194f
C4 VDD2 VP 0.48669f
C5 VP VDD1 2.84637f
C6 VN VDD2 2.51743f
C7 VP VTAIL 3.39897f
C8 VN VDD1 0.155688f
C9 VDD2 VDD1 1.58822f
C10 VDD2 B 4.281981f
C11 VDD1 B 4.682844f
C12 VTAIL B 4.567885f
C13 VN B 13.30595f
C14 VP B 11.859969f
C15 VDD1.t3 B 0.060751f
C16 VDD1.t1 B 0.060751f
C17 VDD1.n0 B 0.462655f
C18 VDD1.t7 B 0.060751f
C19 VDD1.t0 B 0.060751f
C20 VDD1.n1 B 0.461878f
C21 VDD1.t5 B 0.060751f
C22 VDD1.t6 B 0.060751f
C23 VDD1.n2 B 0.461878f
C24 VDD1.n3 B 2.51907f
C25 VDD1.t2 B 0.060751f
C26 VDD1.t4 B 0.060751f
C27 VDD1.n4 B 0.455773f
C28 VDD1.n5 B 2.11868f
C29 VP.n0 B 0.040747f
C30 VP.t1 B 0.538722f
C31 VP.n1 B 0.026987f
C32 VP.n2 B 0.030907f
C33 VP.t2 B 0.538722f
C34 VP.n3 B 0.061427f
C35 VP.n4 B 0.030907f
C36 VP.t7 B 0.538722f
C37 VP.n5 B 0.229567f
C38 VP.n6 B 0.030907f
C39 VP.n7 B 0.058423f
C40 VP.n8 B 0.040747f
C41 VP.t3 B 0.538722f
C42 VP.n9 B 0.026987f
C43 VP.n10 B 0.030907f
C44 VP.t5 B 0.538722f
C45 VP.n11 B 0.061427f
C46 VP.n12 B 0.030907f
C47 VP.t6 B 0.538722f
C48 VP.n13 B 0.311981f
C49 VP.t4 B 0.739295f
C50 VP.n14 B 0.297267f
C51 VP.n15 B 0.26433f
C52 VP.n16 B 0.045372f
C53 VP.n17 B 0.061427f
C54 VP.n18 B 0.024985f
C55 VP.n19 B 0.030907f
C56 VP.n20 B 0.030907f
C57 VP.n21 B 0.030907f
C58 VP.n22 B 0.045372f
C59 VP.n23 B 0.229567f
C60 VP.n24 B 0.041391f
C61 VP.n25 B 0.062429f
C62 VP.n26 B 0.030907f
C63 VP.n27 B 0.030907f
C64 VP.n28 B 0.030907f
C65 VP.n29 B 0.058423f
C66 VP.n30 B 0.049354f
C67 VP.n31 B 0.330884f
C68 VP.n32 B 1.33228f
C69 VP.n33 B 1.35841f
C70 VP.t0 B 0.538722f
C71 VP.n34 B 0.330884f
C72 VP.n35 B 0.049354f
C73 VP.n36 B 0.040747f
C74 VP.n37 B 0.030907f
C75 VP.n38 B 0.030907f
C76 VP.n39 B 0.026987f
C77 VP.n40 B 0.062429f
C78 VP.n41 B 0.041391f
C79 VP.n42 B 0.030907f
C80 VP.n43 B 0.030907f
C81 VP.n44 B 0.045372f
C82 VP.n45 B 0.061427f
C83 VP.n46 B 0.024985f
C84 VP.n47 B 0.030907f
C85 VP.n48 B 0.030907f
C86 VP.n49 B 0.030907f
C87 VP.n50 B 0.045372f
C88 VP.n51 B 0.229567f
C89 VP.n52 B 0.041391f
C90 VP.n53 B 0.062429f
C91 VP.n54 B 0.030907f
C92 VP.n55 B 0.030907f
C93 VP.n56 B 0.030907f
C94 VP.n57 B 0.058423f
C95 VP.n58 B 0.049354f
C96 VP.n59 B 0.330884f
C97 VP.n60 B 0.041068f
C98 VTAIL.t6 B 0.066932f
C99 VTAIL.t13 B 0.066932f
C100 VTAIL.n0 B 0.447671f
C101 VTAIL.n1 B 0.421016f
C102 VTAIL.n2 B 0.035157f
C103 VTAIL.n3 B 0.027235f
C104 VTAIL.n4 B 0.014635f
C105 VTAIL.n5 B 0.025943f
C106 VTAIL.n6 B 0.02017f
C107 VTAIL.t7 B 0.057762f
C108 VTAIL.n7 B 0.098998f
C109 VTAIL.n8 B 0.283725f
C110 VTAIL.n9 B 0.014635f
C111 VTAIL.n10 B 0.015496f
C112 VTAIL.n11 B 0.034591f
C113 VTAIL.n12 B 0.06936f
C114 VTAIL.n13 B 0.015496f
C115 VTAIL.n14 B 0.014635f
C116 VTAIL.n15 B 0.06258f
C117 VTAIL.n16 B 0.03823f
C118 VTAIL.n17 B 0.258706f
C119 VTAIL.n18 B 0.035157f
C120 VTAIL.n19 B 0.027235f
C121 VTAIL.n20 B 0.014635f
C122 VTAIL.n21 B 0.025943f
C123 VTAIL.n22 B 0.02017f
C124 VTAIL.t2 B 0.057762f
C125 VTAIL.n23 B 0.098998f
C126 VTAIL.n24 B 0.283725f
C127 VTAIL.n25 B 0.014635f
C128 VTAIL.n26 B 0.015496f
C129 VTAIL.n27 B 0.034591f
C130 VTAIL.n28 B 0.06936f
C131 VTAIL.n29 B 0.015496f
C132 VTAIL.n30 B 0.014635f
C133 VTAIL.n31 B 0.06258f
C134 VTAIL.n32 B 0.03823f
C135 VTAIL.n33 B 0.258706f
C136 VTAIL.t0 B 0.066932f
C137 VTAIL.t1 B 0.066932f
C138 VTAIL.n34 B 0.447671f
C139 VTAIL.n35 B 0.610335f
C140 VTAIL.n36 B 0.035157f
C141 VTAIL.n37 B 0.027235f
C142 VTAIL.n38 B 0.014635f
C143 VTAIL.n39 B 0.025943f
C144 VTAIL.n40 B 0.02017f
C145 VTAIL.t15 B 0.057762f
C146 VTAIL.n41 B 0.098998f
C147 VTAIL.n42 B 0.283725f
C148 VTAIL.n43 B 0.014635f
C149 VTAIL.n44 B 0.015496f
C150 VTAIL.n45 B 0.034591f
C151 VTAIL.n46 B 0.06936f
C152 VTAIL.n47 B 0.015496f
C153 VTAIL.n48 B 0.014635f
C154 VTAIL.n49 B 0.06258f
C155 VTAIL.n50 B 0.03823f
C156 VTAIL.n51 B 1.01713f
C157 VTAIL.n52 B 0.035157f
C158 VTAIL.n53 B 0.027235f
C159 VTAIL.n54 B 0.014635f
C160 VTAIL.n55 B 0.025943f
C161 VTAIL.n56 B 0.02017f
C162 VTAIL.t12 B 0.057762f
C163 VTAIL.n57 B 0.098998f
C164 VTAIL.n58 B 0.283725f
C165 VTAIL.n59 B 0.014635f
C166 VTAIL.n60 B 0.015496f
C167 VTAIL.n61 B 0.034591f
C168 VTAIL.n62 B 0.06936f
C169 VTAIL.n63 B 0.015496f
C170 VTAIL.n64 B 0.014635f
C171 VTAIL.n65 B 0.06258f
C172 VTAIL.n66 B 0.03823f
C173 VTAIL.n67 B 1.01713f
C174 VTAIL.t10 B 0.066932f
C175 VTAIL.t11 B 0.066932f
C176 VTAIL.n68 B 0.447674f
C177 VTAIL.n69 B 0.610331f
C178 VTAIL.n70 B 0.035157f
C179 VTAIL.n71 B 0.027235f
C180 VTAIL.n72 B 0.014635f
C181 VTAIL.n73 B 0.025943f
C182 VTAIL.n74 B 0.02017f
C183 VTAIL.t9 B 0.057762f
C184 VTAIL.n75 B 0.098998f
C185 VTAIL.n76 B 0.283725f
C186 VTAIL.n77 B 0.014635f
C187 VTAIL.n78 B 0.015496f
C188 VTAIL.n79 B 0.034591f
C189 VTAIL.n80 B 0.06936f
C190 VTAIL.n81 B 0.015496f
C191 VTAIL.n82 B 0.014635f
C192 VTAIL.n83 B 0.06258f
C193 VTAIL.n84 B 0.03823f
C194 VTAIL.n85 B 0.258706f
C195 VTAIL.n86 B 0.035157f
C196 VTAIL.n87 B 0.027235f
C197 VTAIL.n88 B 0.014635f
C198 VTAIL.n89 B 0.025943f
C199 VTAIL.n90 B 0.02017f
C200 VTAIL.t5 B 0.057762f
C201 VTAIL.n91 B 0.098998f
C202 VTAIL.n92 B 0.283725f
C203 VTAIL.n93 B 0.014635f
C204 VTAIL.n94 B 0.015496f
C205 VTAIL.n95 B 0.034591f
C206 VTAIL.n96 B 0.06936f
C207 VTAIL.n97 B 0.015496f
C208 VTAIL.n98 B 0.014635f
C209 VTAIL.n99 B 0.06258f
C210 VTAIL.n100 B 0.03823f
C211 VTAIL.n101 B 0.258706f
C212 VTAIL.t3 B 0.066932f
C213 VTAIL.t4 B 0.066932f
C214 VTAIL.n102 B 0.447674f
C215 VTAIL.n103 B 0.610331f
C216 VTAIL.n104 B 0.035157f
C217 VTAIL.n105 B 0.027235f
C218 VTAIL.n106 B 0.014635f
C219 VTAIL.n107 B 0.025943f
C220 VTAIL.n108 B 0.02017f
C221 VTAIL.t14 B 0.057762f
C222 VTAIL.n109 B 0.098998f
C223 VTAIL.n110 B 0.283725f
C224 VTAIL.n111 B 0.014635f
C225 VTAIL.n112 B 0.015496f
C226 VTAIL.n113 B 0.034591f
C227 VTAIL.n114 B 0.06936f
C228 VTAIL.n115 B 0.015496f
C229 VTAIL.n116 B 0.014635f
C230 VTAIL.n117 B 0.06258f
C231 VTAIL.n118 B 0.03823f
C232 VTAIL.n119 B 1.01713f
C233 VTAIL.n120 B 0.035157f
C234 VTAIL.n121 B 0.027235f
C235 VTAIL.n122 B 0.014635f
C236 VTAIL.n123 B 0.025943f
C237 VTAIL.n124 B 0.02017f
C238 VTAIL.t8 B 0.057762f
C239 VTAIL.n125 B 0.098998f
C240 VTAIL.n126 B 0.283725f
C241 VTAIL.n127 B 0.014635f
C242 VTAIL.n128 B 0.015496f
C243 VTAIL.n129 B 0.034591f
C244 VTAIL.n130 B 0.06936f
C245 VTAIL.n131 B 0.015496f
C246 VTAIL.n132 B 0.014635f
C247 VTAIL.n133 B 0.06258f
C248 VTAIL.n134 B 0.03823f
C249 VTAIL.n135 B 1.01202f
C250 VDD2.t2 B 0.059871f
C251 VDD2.t3 B 0.059871f
C252 VDD2.n0 B 0.455191f
C253 VDD2.t1 B 0.059871f
C254 VDD2.t5 B 0.059871f
C255 VDD2.n1 B 0.455191f
C256 VDD2.n2 B 2.43144f
C257 VDD2.t6 B 0.059871f
C258 VDD2.t0 B 0.059871f
C259 VDD2.n3 B 0.449177f
C260 VDD2.n4 B 2.05832f
C261 VDD2.t7 B 0.059871f
C262 VDD2.t4 B 0.059871f
C263 VDD2.n5 B 0.455165f
C264 VN.n0 B 0.039566f
C265 VN.t5 B 0.523099f
C266 VN.n1 B 0.026204f
C267 VN.n2 B 0.03001f
C268 VN.t0 B 0.523099f
C269 VN.n3 B 0.059645f
C270 VN.n4 B 0.03001f
C271 VN.t7 B 0.523099f
C272 VN.n5 B 0.302934f
C273 VN.t6 B 0.717856f
C274 VN.n6 B 0.288647f
C275 VN.n7 B 0.256665f
C276 VN.n8 B 0.044057f
C277 VN.n9 B 0.059645f
C278 VN.n10 B 0.024261f
C279 VN.n11 B 0.03001f
C280 VN.n12 B 0.03001f
C281 VN.n13 B 0.03001f
C282 VN.n14 B 0.044057f
C283 VN.n15 B 0.22291f
C284 VN.n16 B 0.04019f
C285 VN.n17 B 0.060618f
C286 VN.n18 B 0.03001f
C287 VN.n19 B 0.03001f
C288 VN.n20 B 0.03001f
C289 VN.n21 B 0.056729f
C290 VN.n22 B 0.047922f
C291 VN.n23 B 0.321289f
C292 VN.n24 B 0.039877f
C293 VN.n25 B 0.039566f
C294 VN.t1 B 0.523099f
C295 VN.n26 B 0.026204f
C296 VN.n27 B 0.03001f
C297 VN.t3 B 0.523099f
C298 VN.n28 B 0.059645f
C299 VN.n29 B 0.03001f
C300 VN.t2 B 0.523099f
C301 VN.n30 B 0.302934f
C302 VN.t4 B 0.717856f
C303 VN.n31 B 0.288647f
C304 VN.n32 B 0.256665f
C305 VN.n33 B 0.044057f
C306 VN.n34 B 0.059645f
C307 VN.n35 B 0.024261f
C308 VN.n36 B 0.03001f
C309 VN.n37 B 0.03001f
C310 VN.n38 B 0.03001f
C311 VN.n39 B 0.044057f
C312 VN.n40 B 0.22291f
C313 VN.n41 B 0.04019f
C314 VN.n42 B 0.060618f
C315 VN.n43 B 0.03001f
C316 VN.n44 B 0.03001f
C317 VN.n45 B 0.03001f
C318 VN.n46 B 0.056729f
C319 VN.n47 B 0.047922f
C320 VN.n48 B 0.321289f
C321 VN.n49 B 1.31022f
.ends

