* NGSPICE file created from diff_pair_sample_0303.ext - technology: sky130A

.subckt diff_pair_sample_0303 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t0 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=1.3365 ps=8.43 w=8.1 l=0.4
X1 VDD2.t1 VN.t1 VTAIL.t8 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.4
X2 VTAIL.t7 VN.t2 VDD2.t2 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=1.3365 ps=8.43 w=8.1 l=0.4
X3 VDD1.t5 VP.t0 VTAIL.t0 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.4
X4 VTAIL.t1 VP.t1 VDD1.t4 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=1.3365 ps=8.43 w=8.1 l=0.4
X5 VDD1.t3 VP.t2 VTAIL.t2 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.4
X6 VDD2.t3 VN.t3 VTAIL.t6 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.4
X7 VDD2.t4 VN.t4 VTAIL.t5 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.4
X8 B.t11 B.t9 B.t10 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.4
X9 B.t8 B.t6 B.t7 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.4
X10 VTAIL.t3 VP.t3 VDD1.t2 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=1.3365 pd=8.43 as=1.3365 ps=8.43 w=8.1 l=0.4
X11 B.t5 B.t3 B.t4 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.4
X12 VDD1.t1 VP.t4 VTAIL.t10 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.4
X13 VDD1.t0 VP.t5 VTAIL.t11 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.4
X14 B.t2 B.t0 B.t1 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.4
X15 VDD2.t5 VN.t5 VTAIL.t4 w_n1554_n2588# sky130_fd_pr__pfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.4
R0 VN.n0 VN.t5 609.918
R1 VN.n4 VN.t4 609.918
R2 VN.n2 VN.t3 590.615
R3 VN.n6 VN.t1 590.615
R4 VN.n1 VN.t0 586.232
R5 VN.n5 VN.t2 586.232
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 71.2425
R9 VN.n3 VN.n0 71.2425
R10 VN.n2 VN.n1 43.8187
R11 VN.n6 VN.n5 43.8187
R12 VN VN.n7 37.5289
R13 VN.n5 VN.n4 19.2801
R14 VN.n1 VN.n0 19.2801
R15 VN VN.n3 0.0516364
R16 VDD2.n83 VDD2.n45 756.745
R17 VDD2.n38 VDD2.n0 756.745
R18 VDD2.n84 VDD2.n83 585
R19 VDD2.n82 VDD2.n81 585
R20 VDD2.n49 VDD2.n48 585
R21 VDD2.n76 VDD2.n75 585
R22 VDD2.n74 VDD2.n73 585
R23 VDD2.n53 VDD2.n52 585
R24 VDD2.n68 VDD2.n67 585
R25 VDD2.n66 VDD2.n65 585
R26 VDD2.n57 VDD2.n56 585
R27 VDD2.n60 VDD2.n59 585
R28 VDD2.n15 VDD2.n14 585
R29 VDD2.n12 VDD2.n11 585
R30 VDD2.n21 VDD2.n20 585
R31 VDD2.n23 VDD2.n22 585
R32 VDD2.n8 VDD2.n7 585
R33 VDD2.n29 VDD2.n28 585
R34 VDD2.n31 VDD2.n30 585
R35 VDD2.n4 VDD2.n3 585
R36 VDD2.n37 VDD2.n36 585
R37 VDD2.n39 VDD2.n38 585
R38 VDD2.t1 VDD2.n58 327.473
R39 VDD2.t5 VDD2.n13 327.473
R40 VDD2.n83 VDD2.n82 171.744
R41 VDD2.n82 VDD2.n48 171.744
R42 VDD2.n75 VDD2.n48 171.744
R43 VDD2.n75 VDD2.n74 171.744
R44 VDD2.n74 VDD2.n52 171.744
R45 VDD2.n67 VDD2.n52 171.744
R46 VDD2.n67 VDD2.n66 171.744
R47 VDD2.n66 VDD2.n56 171.744
R48 VDD2.n59 VDD2.n56 171.744
R49 VDD2.n14 VDD2.n11 171.744
R50 VDD2.n21 VDD2.n11 171.744
R51 VDD2.n22 VDD2.n21 171.744
R52 VDD2.n22 VDD2.n7 171.744
R53 VDD2.n29 VDD2.n7 171.744
R54 VDD2.n30 VDD2.n29 171.744
R55 VDD2.n30 VDD2.n3 171.744
R56 VDD2.n37 VDD2.n3 171.744
R57 VDD2.n38 VDD2.n37 171.744
R58 VDD2.n59 VDD2.t1 85.8723
R59 VDD2.n14 VDD2.t5 85.8723
R60 VDD2.n44 VDD2.n43 81.7251
R61 VDD2 VDD2.n89 81.7225
R62 VDD2.n44 VDD2.n42 48.1171
R63 VDD2.n88 VDD2.n87 47.7005
R64 VDD2.n88 VDD2.n44 32.7433
R65 VDD2.n60 VDD2.n58 16.3894
R66 VDD2.n15 VDD2.n13 16.3894
R67 VDD2.n61 VDD2.n57 12.8005
R68 VDD2.n16 VDD2.n12 12.8005
R69 VDD2.n65 VDD2.n64 12.0247
R70 VDD2.n20 VDD2.n19 12.0247
R71 VDD2.n68 VDD2.n55 11.249
R72 VDD2.n23 VDD2.n10 11.249
R73 VDD2.n69 VDD2.n53 10.4732
R74 VDD2.n24 VDD2.n8 10.4732
R75 VDD2.n73 VDD2.n72 9.69747
R76 VDD2.n28 VDD2.n27 9.69747
R77 VDD2.n87 VDD2.n86 9.45567
R78 VDD2.n42 VDD2.n41 9.45567
R79 VDD2.n86 VDD2.n85 9.3005
R80 VDD2.n47 VDD2.n46 9.3005
R81 VDD2.n80 VDD2.n79 9.3005
R82 VDD2.n78 VDD2.n77 9.3005
R83 VDD2.n51 VDD2.n50 9.3005
R84 VDD2.n72 VDD2.n71 9.3005
R85 VDD2.n70 VDD2.n69 9.3005
R86 VDD2.n55 VDD2.n54 9.3005
R87 VDD2.n64 VDD2.n63 9.3005
R88 VDD2.n62 VDD2.n61 9.3005
R89 VDD2.n2 VDD2.n1 9.3005
R90 VDD2.n41 VDD2.n40 9.3005
R91 VDD2.n33 VDD2.n32 9.3005
R92 VDD2.n6 VDD2.n5 9.3005
R93 VDD2.n27 VDD2.n26 9.3005
R94 VDD2.n25 VDD2.n24 9.3005
R95 VDD2.n10 VDD2.n9 9.3005
R96 VDD2.n19 VDD2.n18 9.3005
R97 VDD2.n17 VDD2.n16 9.3005
R98 VDD2.n35 VDD2.n34 9.3005
R99 VDD2.n76 VDD2.n51 8.92171
R100 VDD2.n31 VDD2.n6 8.92171
R101 VDD2.n87 VDD2.n45 8.14595
R102 VDD2.n77 VDD2.n49 8.14595
R103 VDD2.n32 VDD2.n4 8.14595
R104 VDD2.n42 VDD2.n0 8.14595
R105 VDD2.n85 VDD2.n84 7.3702
R106 VDD2.n81 VDD2.n80 7.3702
R107 VDD2.n36 VDD2.n35 7.3702
R108 VDD2.n40 VDD2.n39 7.3702
R109 VDD2.n84 VDD2.n47 6.59444
R110 VDD2.n81 VDD2.n47 6.59444
R111 VDD2.n36 VDD2.n2 6.59444
R112 VDD2.n39 VDD2.n2 6.59444
R113 VDD2.n85 VDD2.n45 5.81868
R114 VDD2.n80 VDD2.n49 5.81868
R115 VDD2.n35 VDD2.n4 5.81868
R116 VDD2.n40 VDD2.n0 5.81868
R117 VDD2.n77 VDD2.n76 5.04292
R118 VDD2.n32 VDD2.n31 5.04292
R119 VDD2.n73 VDD2.n51 4.26717
R120 VDD2.n28 VDD2.n6 4.26717
R121 VDD2.n89 VDD2.t2 4.01346
R122 VDD2.n89 VDD2.t4 4.01346
R123 VDD2.n43 VDD2.t0 4.01346
R124 VDD2.n43 VDD2.t3 4.01346
R125 VDD2.n62 VDD2.n58 3.70995
R126 VDD2.n17 VDD2.n13 3.70995
R127 VDD2.n72 VDD2.n53 3.49141
R128 VDD2.n27 VDD2.n8 3.49141
R129 VDD2.n69 VDD2.n68 2.71565
R130 VDD2.n24 VDD2.n23 2.71565
R131 VDD2.n65 VDD2.n55 1.93989
R132 VDD2.n20 VDD2.n10 1.93989
R133 VDD2.n64 VDD2.n57 1.16414
R134 VDD2.n19 VDD2.n12 1.16414
R135 VDD2 VDD2.n88 0.530672
R136 VDD2.n61 VDD2.n60 0.388379
R137 VDD2.n16 VDD2.n15 0.388379
R138 VDD2.n86 VDD2.n46 0.155672
R139 VDD2.n79 VDD2.n46 0.155672
R140 VDD2.n79 VDD2.n78 0.155672
R141 VDD2.n78 VDD2.n50 0.155672
R142 VDD2.n71 VDD2.n50 0.155672
R143 VDD2.n71 VDD2.n70 0.155672
R144 VDD2.n70 VDD2.n54 0.155672
R145 VDD2.n63 VDD2.n54 0.155672
R146 VDD2.n63 VDD2.n62 0.155672
R147 VDD2.n18 VDD2.n17 0.155672
R148 VDD2.n18 VDD2.n9 0.155672
R149 VDD2.n25 VDD2.n9 0.155672
R150 VDD2.n26 VDD2.n25 0.155672
R151 VDD2.n26 VDD2.n5 0.155672
R152 VDD2.n33 VDD2.n5 0.155672
R153 VDD2.n34 VDD2.n33 0.155672
R154 VDD2.n34 VDD2.n1 0.155672
R155 VDD2.n41 VDD2.n1 0.155672
R156 VTAIL.n178 VTAIL.n140 756.745
R157 VTAIL.n40 VTAIL.n2 756.745
R158 VTAIL.n134 VTAIL.n96 756.745
R159 VTAIL.n88 VTAIL.n50 756.745
R160 VTAIL.n155 VTAIL.n154 585
R161 VTAIL.n152 VTAIL.n151 585
R162 VTAIL.n161 VTAIL.n160 585
R163 VTAIL.n163 VTAIL.n162 585
R164 VTAIL.n148 VTAIL.n147 585
R165 VTAIL.n169 VTAIL.n168 585
R166 VTAIL.n171 VTAIL.n170 585
R167 VTAIL.n144 VTAIL.n143 585
R168 VTAIL.n177 VTAIL.n176 585
R169 VTAIL.n179 VTAIL.n178 585
R170 VTAIL.n17 VTAIL.n16 585
R171 VTAIL.n14 VTAIL.n13 585
R172 VTAIL.n23 VTAIL.n22 585
R173 VTAIL.n25 VTAIL.n24 585
R174 VTAIL.n10 VTAIL.n9 585
R175 VTAIL.n31 VTAIL.n30 585
R176 VTAIL.n33 VTAIL.n32 585
R177 VTAIL.n6 VTAIL.n5 585
R178 VTAIL.n39 VTAIL.n38 585
R179 VTAIL.n41 VTAIL.n40 585
R180 VTAIL.n135 VTAIL.n134 585
R181 VTAIL.n133 VTAIL.n132 585
R182 VTAIL.n100 VTAIL.n99 585
R183 VTAIL.n127 VTAIL.n126 585
R184 VTAIL.n125 VTAIL.n124 585
R185 VTAIL.n104 VTAIL.n103 585
R186 VTAIL.n119 VTAIL.n118 585
R187 VTAIL.n117 VTAIL.n116 585
R188 VTAIL.n108 VTAIL.n107 585
R189 VTAIL.n111 VTAIL.n110 585
R190 VTAIL.n89 VTAIL.n88 585
R191 VTAIL.n87 VTAIL.n86 585
R192 VTAIL.n54 VTAIL.n53 585
R193 VTAIL.n81 VTAIL.n80 585
R194 VTAIL.n79 VTAIL.n78 585
R195 VTAIL.n58 VTAIL.n57 585
R196 VTAIL.n73 VTAIL.n72 585
R197 VTAIL.n71 VTAIL.n70 585
R198 VTAIL.n62 VTAIL.n61 585
R199 VTAIL.n65 VTAIL.n64 585
R200 VTAIL.t6 VTAIL.n153 327.473
R201 VTAIL.t2 VTAIL.n15 327.473
R202 VTAIL.t0 VTAIL.n109 327.473
R203 VTAIL.t5 VTAIL.n63 327.473
R204 VTAIL.n154 VTAIL.n151 171.744
R205 VTAIL.n161 VTAIL.n151 171.744
R206 VTAIL.n162 VTAIL.n161 171.744
R207 VTAIL.n162 VTAIL.n147 171.744
R208 VTAIL.n169 VTAIL.n147 171.744
R209 VTAIL.n170 VTAIL.n169 171.744
R210 VTAIL.n170 VTAIL.n143 171.744
R211 VTAIL.n177 VTAIL.n143 171.744
R212 VTAIL.n178 VTAIL.n177 171.744
R213 VTAIL.n16 VTAIL.n13 171.744
R214 VTAIL.n23 VTAIL.n13 171.744
R215 VTAIL.n24 VTAIL.n23 171.744
R216 VTAIL.n24 VTAIL.n9 171.744
R217 VTAIL.n31 VTAIL.n9 171.744
R218 VTAIL.n32 VTAIL.n31 171.744
R219 VTAIL.n32 VTAIL.n5 171.744
R220 VTAIL.n39 VTAIL.n5 171.744
R221 VTAIL.n40 VTAIL.n39 171.744
R222 VTAIL.n134 VTAIL.n133 171.744
R223 VTAIL.n133 VTAIL.n99 171.744
R224 VTAIL.n126 VTAIL.n99 171.744
R225 VTAIL.n126 VTAIL.n125 171.744
R226 VTAIL.n125 VTAIL.n103 171.744
R227 VTAIL.n118 VTAIL.n103 171.744
R228 VTAIL.n118 VTAIL.n117 171.744
R229 VTAIL.n117 VTAIL.n107 171.744
R230 VTAIL.n110 VTAIL.n107 171.744
R231 VTAIL.n88 VTAIL.n87 171.744
R232 VTAIL.n87 VTAIL.n53 171.744
R233 VTAIL.n80 VTAIL.n53 171.744
R234 VTAIL.n80 VTAIL.n79 171.744
R235 VTAIL.n79 VTAIL.n57 171.744
R236 VTAIL.n72 VTAIL.n57 171.744
R237 VTAIL.n72 VTAIL.n71 171.744
R238 VTAIL.n71 VTAIL.n61 171.744
R239 VTAIL.n64 VTAIL.n61 171.744
R240 VTAIL.n154 VTAIL.t6 85.8723
R241 VTAIL.n16 VTAIL.t2 85.8723
R242 VTAIL.n110 VTAIL.t0 85.8723
R243 VTAIL.n64 VTAIL.t5 85.8723
R244 VTAIL.n95 VTAIL.n94 64.9445
R245 VTAIL.n49 VTAIL.n48 64.9445
R246 VTAIL.n1 VTAIL.n0 64.9444
R247 VTAIL.n47 VTAIL.n46 64.9444
R248 VTAIL.n183 VTAIL.n182 31.0217
R249 VTAIL.n45 VTAIL.n44 31.0217
R250 VTAIL.n139 VTAIL.n138 31.0217
R251 VTAIL.n93 VTAIL.n92 31.0217
R252 VTAIL.n49 VTAIL.n47 20.6083
R253 VTAIL.n183 VTAIL.n139 19.9789
R254 VTAIL.n155 VTAIL.n153 16.3894
R255 VTAIL.n17 VTAIL.n15 16.3894
R256 VTAIL.n111 VTAIL.n109 16.3894
R257 VTAIL.n65 VTAIL.n63 16.3894
R258 VTAIL.n156 VTAIL.n152 12.8005
R259 VTAIL.n18 VTAIL.n14 12.8005
R260 VTAIL.n112 VTAIL.n108 12.8005
R261 VTAIL.n66 VTAIL.n62 12.8005
R262 VTAIL.n160 VTAIL.n159 12.0247
R263 VTAIL.n22 VTAIL.n21 12.0247
R264 VTAIL.n116 VTAIL.n115 12.0247
R265 VTAIL.n70 VTAIL.n69 12.0247
R266 VTAIL.n163 VTAIL.n150 11.249
R267 VTAIL.n25 VTAIL.n12 11.249
R268 VTAIL.n119 VTAIL.n106 11.249
R269 VTAIL.n73 VTAIL.n60 11.249
R270 VTAIL.n164 VTAIL.n148 10.4732
R271 VTAIL.n26 VTAIL.n10 10.4732
R272 VTAIL.n120 VTAIL.n104 10.4732
R273 VTAIL.n74 VTAIL.n58 10.4732
R274 VTAIL.n168 VTAIL.n167 9.69747
R275 VTAIL.n30 VTAIL.n29 9.69747
R276 VTAIL.n124 VTAIL.n123 9.69747
R277 VTAIL.n78 VTAIL.n77 9.69747
R278 VTAIL.n182 VTAIL.n181 9.45567
R279 VTAIL.n44 VTAIL.n43 9.45567
R280 VTAIL.n138 VTAIL.n137 9.45567
R281 VTAIL.n92 VTAIL.n91 9.45567
R282 VTAIL.n142 VTAIL.n141 9.3005
R283 VTAIL.n181 VTAIL.n180 9.3005
R284 VTAIL.n173 VTAIL.n172 9.3005
R285 VTAIL.n146 VTAIL.n145 9.3005
R286 VTAIL.n167 VTAIL.n166 9.3005
R287 VTAIL.n165 VTAIL.n164 9.3005
R288 VTAIL.n150 VTAIL.n149 9.3005
R289 VTAIL.n159 VTAIL.n158 9.3005
R290 VTAIL.n157 VTAIL.n156 9.3005
R291 VTAIL.n175 VTAIL.n174 9.3005
R292 VTAIL.n4 VTAIL.n3 9.3005
R293 VTAIL.n43 VTAIL.n42 9.3005
R294 VTAIL.n35 VTAIL.n34 9.3005
R295 VTAIL.n8 VTAIL.n7 9.3005
R296 VTAIL.n29 VTAIL.n28 9.3005
R297 VTAIL.n27 VTAIL.n26 9.3005
R298 VTAIL.n12 VTAIL.n11 9.3005
R299 VTAIL.n21 VTAIL.n20 9.3005
R300 VTAIL.n19 VTAIL.n18 9.3005
R301 VTAIL.n37 VTAIL.n36 9.3005
R302 VTAIL.n98 VTAIL.n97 9.3005
R303 VTAIL.n131 VTAIL.n130 9.3005
R304 VTAIL.n129 VTAIL.n128 9.3005
R305 VTAIL.n102 VTAIL.n101 9.3005
R306 VTAIL.n123 VTAIL.n122 9.3005
R307 VTAIL.n121 VTAIL.n120 9.3005
R308 VTAIL.n106 VTAIL.n105 9.3005
R309 VTAIL.n115 VTAIL.n114 9.3005
R310 VTAIL.n113 VTAIL.n112 9.3005
R311 VTAIL.n137 VTAIL.n136 9.3005
R312 VTAIL.n91 VTAIL.n90 9.3005
R313 VTAIL.n52 VTAIL.n51 9.3005
R314 VTAIL.n85 VTAIL.n84 9.3005
R315 VTAIL.n83 VTAIL.n82 9.3005
R316 VTAIL.n56 VTAIL.n55 9.3005
R317 VTAIL.n77 VTAIL.n76 9.3005
R318 VTAIL.n75 VTAIL.n74 9.3005
R319 VTAIL.n60 VTAIL.n59 9.3005
R320 VTAIL.n69 VTAIL.n68 9.3005
R321 VTAIL.n67 VTAIL.n66 9.3005
R322 VTAIL.n171 VTAIL.n146 8.92171
R323 VTAIL.n33 VTAIL.n8 8.92171
R324 VTAIL.n127 VTAIL.n102 8.92171
R325 VTAIL.n81 VTAIL.n56 8.92171
R326 VTAIL.n172 VTAIL.n144 8.14595
R327 VTAIL.n182 VTAIL.n140 8.14595
R328 VTAIL.n34 VTAIL.n6 8.14595
R329 VTAIL.n44 VTAIL.n2 8.14595
R330 VTAIL.n138 VTAIL.n96 8.14595
R331 VTAIL.n128 VTAIL.n100 8.14595
R332 VTAIL.n92 VTAIL.n50 8.14595
R333 VTAIL.n82 VTAIL.n54 8.14595
R334 VTAIL.n176 VTAIL.n175 7.3702
R335 VTAIL.n180 VTAIL.n179 7.3702
R336 VTAIL.n38 VTAIL.n37 7.3702
R337 VTAIL.n42 VTAIL.n41 7.3702
R338 VTAIL.n136 VTAIL.n135 7.3702
R339 VTAIL.n132 VTAIL.n131 7.3702
R340 VTAIL.n90 VTAIL.n89 7.3702
R341 VTAIL.n86 VTAIL.n85 7.3702
R342 VTAIL.n176 VTAIL.n142 6.59444
R343 VTAIL.n179 VTAIL.n142 6.59444
R344 VTAIL.n38 VTAIL.n4 6.59444
R345 VTAIL.n41 VTAIL.n4 6.59444
R346 VTAIL.n135 VTAIL.n98 6.59444
R347 VTAIL.n132 VTAIL.n98 6.59444
R348 VTAIL.n89 VTAIL.n52 6.59444
R349 VTAIL.n86 VTAIL.n52 6.59444
R350 VTAIL.n175 VTAIL.n144 5.81868
R351 VTAIL.n180 VTAIL.n140 5.81868
R352 VTAIL.n37 VTAIL.n6 5.81868
R353 VTAIL.n42 VTAIL.n2 5.81868
R354 VTAIL.n136 VTAIL.n96 5.81868
R355 VTAIL.n131 VTAIL.n100 5.81868
R356 VTAIL.n90 VTAIL.n50 5.81868
R357 VTAIL.n85 VTAIL.n54 5.81868
R358 VTAIL.n172 VTAIL.n171 5.04292
R359 VTAIL.n34 VTAIL.n33 5.04292
R360 VTAIL.n128 VTAIL.n127 5.04292
R361 VTAIL.n82 VTAIL.n81 5.04292
R362 VTAIL.n168 VTAIL.n146 4.26717
R363 VTAIL.n30 VTAIL.n8 4.26717
R364 VTAIL.n124 VTAIL.n102 4.26717
R365 VTAIL.n78 VTAIL.n56 4.26717
R366 VTAIL.n0 VTAIL.t4 4.01346
R367 VTAIL.n0 VTAIL.t9 4.01346
R368 VTAIL.n46 VTAIL.t11 4.01346
R369 VTAIL.n46 VTAIL.t3 4.01346
R370 VTAIL.n94 VTAIL.t10 4.01346
R371 VTAIL.n94 VTAIL.t1 4.01346
R372 VTAIL.n48 VTAIL.t8 4.01346
R373 VTAIL.n48 VTAIL.t7 4.01346
R374 VTAIL.n157 VTAIL.n153 3.70995
R375 VTAIL.n19 VTAIL.n15 3.70995
R376 VTAIL.n67 VTAIL.n63 3.70995
R377 VTAIL.n113 VTAIL.n109 3.70995
R378 VTAIL.n167 VTAIL.n148 3.49141
R379 VTAIL.n29 VTAIL.n10 3.49141
R380 VTAIL.n123 VTAIL.n104 3.49141
R381 VTAIL.n77 VTAIL.n58 3.49141
R382 VTAIL.n164 VTAIL.n163 2.71565
R383 VTAIL.n26 VTAIL.n25 2.71565
R384 VTAIL.n120 VTAIL.n119 2.71565
R385 VTAIL.n74 VTAIL.n73 2.71565
R386 VTAIL.n160 VTAIL.n150 1.93989
R387 VTAIL.n22 VTAIL.n12 1.93989
R388 VTAIL.n116 VTAIL.n106 1.93989
R389 VTAIL.n70 VTAIL.n60 1.93989
R390 VTAIL.n159 VTAIL.n152 1.16414
R391 VTAIL.n21 VTAIL.n14 1.16414
R392 VTAIL.n115 VTAIL.n108 1.16414
R393 VTAIL.n69 VTAIL.n62 1.16414
R394 VTAIL.n95 VTAIL.n93 0.784983
R395 VTAIL.n45 VTAIL.n1 0.784983
R396 VTAIL.n93 VTAIL.n49 0.62981
R397 VTAIL.n139 VTAIL.n95 0.62981
R398 VTAIL.n47 VTAIL.n45 0.62981
R399 VTAIL VTAIL.n183 0.414293
R400 VTAIL.n156 VTAIL.n155 0.388379
R401 VTAIL.n18 VTAIL.n17 0.388379
R402 VTAIL.n112 VTAIL.n111 0.388379
R403 VTAIL.n66 VTAIL.n65 0.388379
R404 VTAIL VTAIL.n1 0.216017
R405 VTAIL.n158 VTAIL.n157 0.155672
R406 VTAIL.n158 VTAIL.n149 0.155672
R407 VTAIL.n165 VTAIL.n149 0.155672
R408 VTAIL.n166 VTAIL.n165 0.155672
R409 VTAIL.n166 VTAIL.n145 0.155672
R410 VTAIL.n173 VTAIL.n145 0.155672
R411 VTAIL.n174 VTAIL.n173 0.155672
R412 VTAIL.n174 VTAIL.n141 0.155672
R413 VTAIL.n181 VTAIL.n141 0.155672
R414 VTAIL.n20 VTAIL.n19 0.155672
R415 VTAIL.n20 VTAIL.n11 0.155672
R416 VTAIL.n27 VTAIL.n11 0.155672
R417 VTAIL.n28 VTAIL.n27 0.155672
R418 VTAIL.n28 VTAIL.n7 0.155672
R419 VTAIL.n35 VTAIL.n7 0.155672
R420 VTAIL.n36 VTAIL.n35 0.155672
R421 VTAIL.n36 VTAIL.n3 0.155672
R422 VTAIL.n43 VTAIL.n3 0.155672
R423 VTAIL.n137 VTAIL.n97 0.155672
R424 VTAIL.n130 VTAIL.n97 0.155672
R425 VTAIL.n130 VTAIL.n129 0.155672
R426 VTAIL.n129 VTAIL.n101 0.155672
R427 VTAIL.n122 VTAIL.n101 0.155672
R428 VTAIL.n122 VTAIL.n121 0.155672
R429 VTAIL.n121 VTAIL.n105 0.155672
R430 VTAIL.n114 VTAIL.n105 0.155672
R431 VTAIL.n114 VTAIL.n113 0.155672
R432 VTAIL.n91 VTAIL.n51 0.155672
R433 VTAIL.n84 VTAIL.n51 0.155672
R434 VTAIL.n84 VTAIL.n83 0.155672
R435 VTAIL.n83 VTAIL.n55 0.155672
R436 VTAIL.n76 VTAIL.n55 0.155672
R437 VTAIL.n76 VTAIL.n75 0.155672
R438 VTAIL.n75 VTAIL.n59 0.155672
R439 VTAIL.n68 VTAIL.n59 0.155672
R440 VTAIL.n68 VTAIL.n67 0.155672
R441 VP.n1 VP.t4 609.918
R442 VP.n8 VP.t2 590.615
R443 VP.n6 VP.t5 590.615
R444 VP.n3 VP.t0 590.615
R445 VP.n7 VP.t3 586.232
R446 VP.n2 VP.t1 586.232
R447 VP.n9 VP.n8 161.3
R448 VP.n4 VP.n3 161.3
R449 VP.n7 VP.n0 161.3
R450 VP.n6 VP.n5 161.3
R451 VP.n4 VP.n1 71.2425
R452 VP.n7 VP.n6 43.8187
R453 VP.n8 VP.n7 43.8187
R454 VP.n3 VP.n2 43.8187
R455 VP.n5 VP.n4 37.1482
R456 VP.n2 VP.n1 19.2801
R457 VP.n5 VP.n0 0.189894
R458 VP.n9 VP.n0 0.189894
R459 VP VP.n9 0.0516364
R460 VDD1.n38 VDD1.n0 756.745
R461 VDD1.n81 VDD1.n43 756.745
R462 VDD1.n39 VDD1.n38 585
R463 VDD1.n37 VDD1.n36 585
R464 VDD1.n4 VDD1.n3 585
R465 VDD1.n31 VDD1.n30 585
R466 VDD1.n29 VDD1.n28 585
R467 VDD1.n8 VDD1.n7 585
R468 VDD1.n23 VDD1.n22 585
R469 VDD1.n21 VDD1.n20 585
R470 VDD1.n12 VDD1.n11 585
R471 VDD1.n15 VDD1.n14 585
R472 VDD1.n58 VDD1.n57 585
R473 VDD1.n55 VDD1.n54 585
R474 VDD1.n64 VDD1.n63 585
R475 VDD1.n66 VDD1.n65 585
R476 VDD1.n51 VDD1.n50 585
R477 VDD1.n72 VDD1.n71 585
R478 VDD1.n74 VDD1.n73 585
R479 VDD1.n47 VDD1.n46 585
R480 VDD1.n80 VDD1.n79 585
R481 VDD1.n82 VDD1.n81 585
R482 VDD1.t1 VDD1.n13 327.473
R483 VDD1.t0 VDD1.n56 327.473
R484 VDD1.n38 VDD1.n37 171.744
R485 VDD1.n37 VDD1.n3 171.744
R486 VDD1.n30 VDD1.n3 171.744
R487 VDD1.n30 VDD1.n29 171.744
R488 VDD1.n29 VDD1.n7 171.744
R489 VDD1.n22 VDD1.n7 171.744
R490 VDD1.n22 VDD1.n21 171.744
R491 VDD1.n21 VDD1.n11 171.744
R492 VDD1.n14 VDD1.n11 171.744
R493 VDD1.n57 VDD1.n54 171.744
R494 VDD1.n64 VDD1.n54 171.744
R495 VDD1.n65 VDD1.n64 171.744
R496 VDD1.n65 VDD1.n50 171.744
R497 VDD1.n72 VDD1.n50 171.744
R498 VDD1.n73 VDD1.n72 171.744
R499 VDD1.n73 VDD1.n46 171.744
R500 VDD1.n80 VDD1.n46 171.744
R501 VDD1.n81 VDD1.n80 171.744
R502 VDD1.n14 VDD1.t1 85.8723
R503 VDD1.n57 VDD1.t0 85.8723
R504 VDD1.n87 VDD1.n86 81.7251
R505 VDD1.n89 VDD1.n88 81.6233
R506 VDD1 VDD1.n42 48.2307
R507 VDD1.n87 VDD1.n85 48.1171
R508 VDD1.n89 VDD1.n87 33.641
R509 VDD1.n15 VDD1.n13 16.3894
R510 VDD1.n58 VDD1.n56 16.3894
R511 VDD1.n16 VDD1.n12 12.8005
R512 VDD1.n59 VDD1.n55 12.8005
R513 VDD1.n20 VDD1.n19 12.0247
R514 VDD1.n63 VDD1.n62 12.0247
R515 VDD1.n23 VDD1.n10 11.249
R516 VDD1.n66 VDD1.n53 11.249
R517 VDD1.n24 VDD1.n8 10.4732
R518 VDD1.n67 VDD1.n51 10.4732
R519 VDD1.n28 VDD1.n27 9.69747
R520 VDD1.n71 VDD1.n70 9.69747
R521 VDD1.n42 VDD1.n41 9.45567
R522 VDD1.n85 VDD1.n84 9.45567
R523 VDD1.n41 VDD1.n40 9.3005
R524 VDD1.n2 VDD1.n1 9.3005
R525 VDD1.n35 VDD1.n34 9.3005
R526 VDD1.n33 VDD1.n32 9.3005
R527 VDD1.n6 VDD1.n5 9.3005
R528 VDD1.n27 VDD1.n26 9.3005
R529 VDD1.n25 VDD1.n24 9.3005
R530 VDD1.n10 VDD1.n9 9.3005
R531 VDD1.n19 VDD1.n18 9.3005
R532 VDD1.n17 VDD1.n16 9.3005
R533 VDD1.n45 VDD1.n44 9.3005
R534 VDD1.n84 VDD1.n83 9.3005
R535 VDD1.n76 VDD1.n75 9.3005
R536 VDD1.n49 VDD1.n48 9.3005
R537 VDD1.n70 VDD1.n69 9.3005
R538 VDD1.n68 VDD1.n67 9.3005
R539 VDD1.n53 VDD1.n52 9.3005
R540 VDD1.n62 VDD1.n61 9.3005
R541 VDD1.n60 VDD1.n59 9.3005
R542 VDD1.n78 VDD1.n77 9.3005
R543 VDD1.n31 VDD1.n6 8.92171
R544 VDD1.n74 VDD1.n49 8.92171
R545 VDD1.n42 VDD1.n0 8.14595
R546 VDD1.n32 VDD1.n4 8.14595
R547 VDD1.n75 VDD1.n47 8.14595
R548 VDD1.n85 VDD1.n43 8.14595
R549 VDD1.n40 VDD1.n39 7.3702
R550 VDD1.n36 VDD1.n35 7.3702
R551 VDD1.n79 VDD1.n78 7.3702
R552 VDD1.n83 VDD1.n82 7.3702
R553 VDD1.n39 VDD1.n2 6.59444
R554 VDD1.n36 VDD1.n2 6.59444
R555 VDD1.n79 VDD1.n45 6.59444
R556 VDD1.n82 VDD1.n45 6.59444
R557 VDD1.n40 VDD1.n0 5.81868
R558 VDD1.n35 VDD1.n4 5.81868
R559 VDD1.n78 VDD1.n47 5.81868
R560 VDD1.n83 VDD1.n43 5.81868
R561 VDD1.n32 VDD1.n31 5.04292
R562 VDD1.n75 VDD1.n74 5.04292
R563 VDD1.n28 VDD1.n6 4.26717
R564 VDD1.n71 VDD1.n49 4.26717
R565 VDD1.n88 VDD1.t4 4.01346
R566 VDD1.n88 VDD1.t5 4.01346
R567 VDD1.n86 VDD1.t2 4.01346
R568 VDD1.n86 VDD1.t3 4.01346
R569 VDD1.n17 VDD1.n13 3.70995
R570 VDD1.n60 VDD1.n56 3.70995
R571 VDD1.n27 VDD1.n8 3.49141
R572 VDD1.n70 VDD1.n51 3.49141
R573 VDD1.n24 VDD1.n23 2.71565
R574 VDD1.n67 VDD1.n66 2.71565
R575 VDD1.n20 VDD1.n10 1.93989
R576 VDD1.n63 VDD1.n53 1.93989
R577 VDD1.n19 VDD1.n12 1.16414
R578 VDD1.n62 VDD1.n55 1.16414
R579 VDD1.n16 VDD1.n15 0.388379
R580 VDD1.n59 VDD1.n58 0.388379
R581 VDD1.n41 VDD1.n1 0.155672
R582 VDD1.n34 VDD1.n1 0.155672
R583 VDD1.n34 VDD1.n33 0.155672
R584 VDD1.n33 VDD1.n5 0.155672
R585 VDD1.n26 VDD1.n5 0.155672
R586 VDD1.n26 VDD1.n25 0.155672
R587 VDD1.n25 VDD1.n9 0.155672
R588 VDD1.n18 VDD1.n9 0.155672
R589 VDD1.n18 VDD1.n17 0.155672
R590 VDD1.n61 VDD1.n60 0.155672
R591 VDD1.n61 VDD1.n52 0.155672
R592 VDD1.n68 VDD1.n52 0.155672
R593 VDD1.n69 VDD1.n68 0.155672
R594 VDD1.n69 VDD1.n48 0.155672
R595 VDD1.n76 VDD1.n48 0.155672
R596 VDD1.n77 VDD1.n76 0.155672
R597 VDD1.n77 VDD1.n44 0.155672
R598 VDD1.n84 VDD1.n44 0.155672
R599 VDD1 VDD1.n89 0.0996379
R600 B.n177 B.t3 697.446
R601 B.n82 B.t6 697.446
R602 B.n32 B.t0 697.446
R603 B.n26 B.t9 697.446
R604 B.n242 B.n241 585
R605 B.n240 B.n67 585
R606 B.n239 B.n238 585
R607 B.n237 B.n68 585
R608 B.n236 B.n235 585
R609 B.n234 B.n69 585
R610 B.n233 B.n232 585
R611 B.n231 B.n70 585
R612 B.n230 B.n229 585
R613 B.n228 B.n71 585
R614 B.n227 B.n226 585
R615 B.n225 B.n72 585
R616 B.n224 B.n223 585
R617 B.n222 B.n73 585
R618 B.n221 B.n220 585
R619 B.n219 B.n74 585
R620 B.n218 B.n217 585
R621 B.n216 B.n75 585
R622 B.n215 B.n214 585
R623 B.n213 B.n76 585
R624 B.n212 B.n211 585
R625 B.n210 B.n77 585
R626 B.n209 B.n208 585
R627 B.n207 B.n78 585
R628 B.n206 B.n205 585
R629 B.n204 B.n79 585
R630 B.n203 B.n202 585
R631 B.n201 B.n80 585
R632 B.n200 B.n199 585
R633 B.n198 B.n81 585
R634 B.n196 B.n195 585
R635 B.n194 B.n84 585
R636 B.n193 B.n192 585
R637 B.n191 B.n85 585
R638 B.n190 B.n189 585
R639 B.n188 B.n86 585
R640 B.n187 B.n186 585
R641 B.n185 B.n87 585
R642 B.n184 B.n183 585
R643 B.n182 B.n88 585
R644 B.n181 B.n180 585
R645 B.n176 B.n89 585
R646 B.n175 B.n174 585
R647 B.n173 B.n90 585
R648 B.n172 B.n171 585
R649 B.n170 B.n91 585
R650 B.n169 B.n168 585
R651 B.n167 B.n92 585
R652 B.n166 B.n165 585
R653 B.n164 B.n93 585
R654 B.n163 B.n162 585
R655 B.n161 B.n94 585
R656 B.n160 B.n159 585
R657 B.n158 B.n95 585
R658 B.n157 B.n156 585
R659 B.n155 B.n96 585
R660 B.n154 B.n153 585
R661 B.n152 B.n97 585
R662 B.n151 B.n150 585
R663 B.n149 B.n98 585
R664 B.n148 B.n147 585
R665 B.n146 B.n99 585
R666 B.n145 B.n144 585
R667 B.n143 B.n100 585
R668 B.n142 B.n141 585
R669 B.n140 B.n101 585
R670 B.n139 B.n138 585
R671 B.n137 B.n102 585
R672 B.n136 B.n135 585
R673 B.n134 B.n103 585
R674 B.n243 B.n66 585
R675 B.n245 B.n244 585
R676 B.n246 B.n65 585
R677 B.n248 B.n247 585
R678 B.n249 B.n64 585
R679 B.n251 B.n250 585
R680 B.n252 B.n63 585
R681 B.n254 B.n253 585
R682 B.n255 B.n62 585
R683 B.n257 B.n256 585
R684 B.n258 B.n61 585
R685 B.n260 B.n259 585
R686 B.n261 B.n60 585
R687 B.n263 B.n262 585
R688 B.n264 B.n59 585
R689 B.n266 B.n265 585
R690 B.n267 B.n58 585
R691 B.n269 B.n268 585
R692 B.n270 B.n57 585
R693 B.n272 B.n271 585
R694 B.n273 B.n56 585
R695 B.n275 B.n274 585
R696 B.n276 B.n55 585
R697 B.n278 B.n277 585
R698 B.n279 B.n54 585
R699 B.n281 B.n280 585
R700 B.n282 B.n53 585
R701 B.n284 B.n283 585
R702 B.n285 B.n52 585
R703 B.n287 B.n286 585
R704 B.n288 B.n51 585
R705 B.n290 B.n289 585
R706 B.n291 B.n50 585
R707 B.n293 B.n292 585
R708 B.n399 B.n10 585
R709 B.n398 B.n397 585
R710 B.n396 B.n11 585
R711 B.n395 B.n394 585
R712 B.n393 B.n12 585
R713 B.n392 B.n391 585
R714 B.n390 B.n13 585
R715 B.n389 B.n388 585
R716 B.n387 B.n14 585
R717 B.n386 B.n385 585
R718 B.n384 B.n15 585
R719 B.n383 B.n382 585
R720 B.n381 B.n16 585
R721 B.n380 B.n379 585
R722 B.n378 B.n17 585
R723 B.n377 B.n376 585
R724 B.n375 B.n18 585
R725 B.n374 B.n373 585
R726 B.n372 B.n19 585
R727 B.n371 B.n370 585
R728 B.n369 B.n20 585
R729 B.n368 B.n367 585
R730 B.n366 B.n21 585
R731 B.n365 B.n364 585
R732 B.n363 B.n22 585
R733 B.n362 B.n361 585
R734 B.n360 B.n23 585
R735 B.n359 B.n358 585
R736 B.n357 B.n24 585
R737 B.n356 B.n355 585
R738 B.n353 B.n25 585
R739 B.n352 B.n351 585
R740 B.n350 B.n28 585
R741 B.n349 B.n348 585
R742 B.n347 B.n29 585
R743 B.n346 B.n345 585
R744 B.n344 B.n30 585
R745 B.n343 B.n342 585
R746 B.n341 B.n31 585
R747 B.n340 B.n339 585
R748 B.n338 B.n337 585
R749 B.n336 B.n35 585
R750 B.n335 B.n334 585
R751 B.n333 B.n36 585
R752 B.n332 B.n331 585
R753 B.n330 B.n37 585
R754 B.n329 B.n328 585
R755 B.n327 B.n38 585
R756 B.n326 B.n325 585
R757 B.n324 B.n39 585
R758 B.n323 B.n322 585
R759 B.n321 B.n40 585
R760 B.n320 B.n319 585
R761 B.n318 B.n41 585
R762 B.n317 B.n316 585
R763 B.n315 B.n42 585
R764 B.n314 B.n313 585
R765 B.n312 B.n43 585
R766 B.n311 B.n310 585
R767 B.n309 B.n44 585
R768 B.n308 B.n307 585
R769 B.n306 B.n45 585
R770 B.n305 B.n304 585
R771 B.n303 B.n46 585
R772 B.n302 B.n301 585
R773 B.n300 B.n47 585
R774 B.n299 B.n298 585
R775 B.n297 B.n48 585
R776 B.n296 B.n295 585
R777 B.n294 B.n49 585
R778 B.n401 B.n400 585
R779 B.n402 B.n9 585
R780 B.n404 B.n403 585
R781 B.n405 B.n8 585
R782 B.n407 B.n406 585
R783 B.n408 B.n7 585
R784 B.n410 B.n409 585
R785 B.n411 B.n6 585
R786 B.n413 B.n412 585
R787 B.n414 B.n5 585
R788 B.n416 B.n415 585
R789 B.n417 B.n4 585
R790 B.n419 B.n418 585
R791 B.n420 B.n3 585
R792 B.n422 B.n421 585
R793 B.n423 B.n0 585
R794 B.n2 B.n1 585
R795 B.n112 B.n111 585
R796 B.n113 B.n110 585
R797 B.n115 B.n114 585
R798 B.n116 B.n109 585
R799 B.n118 B.n117 585
R800 B.n119 B.n108 585
R801 B.n121 B.n120 585
R802 B.n122 B.n107 585
R803 B.n124 B.n123 585
R804 B.n125 B.n106 585
R805 B.n127 B.n126 585
R806 B.n128 B.n105 585
R807 B.n130 B.n129 585
R808 B.n131 B.n104 585
R809 B.n133 B.n132 585
R810 B.n132 B.n103 521.33
R811 B.n243 B.n242 521.33
R812 B.n292 B.n49 521.33
R813 B.n400 B.n399 521.33
R814 B.n82 B.t7 319.788
R815 B.n32 B.t2 319.788
R816 B.n177 B.t4 319.788
R817 B.n26 B.t11 319.788
R818 B.n83 B.t8 305.63
R819 B.n33 B.t1 305.63
R820 B.n178 B.t5 305.63
R821 B.n27 B.t10 305.63
R822 B.n425 B.n424 256.663
R823 B.n424 B.n423 235.042
R824 B.n424 B.n2 235.042
R825 B.n136 B.n103 163.367
R826 B.n137 B.n136 163.367
R827 B.n138 B.n137 163.367
R828 B.n138 B.n101 163.367
R829 B.n142 B.n101 163.367
R830 B.n143 B.n142 163.367
R831 B.n144 B.n143 163.367
R832 B.n144 B.n99 163.367
R833 B.n148 B.n99 163.367
R834 B.n149 B.n148 163.367
R835 B.n150 B.n149 163.367
R836 B.n150 B.n97 163.367
R837 B.n154 B.n97 163.367
R838 B.n155 B.n154 163.367
R839 B.n156 B.n155 163.367
R840 B.n156 B.n95 163.367
R841 B.n160 B.n95 163.367
R842 B.n161 B.n160 163.367
R843 B.n162 B.n161 163.367
R844 B.n162 B.n93 163.367
R845 B.n166 B.n93 163.367
R846 B.n167 B.n166 163.367
R847 B.n168 B.n167 163.367
R848 B.n168 B.n91 163.367
R849 B.n172 B.n91 163.367
R850 B.n173 B.n172 163.367
R851 B.n174 B.n173 163.367
R852 B.n174 B.n89 163.367
R853 B.n181 B.n89 163.367
R854 B.n182 B.n181 163.367
R855 B.n183 B.n182 163.367
R856 B.n183 B.n87 163.367
R857 B.n187 B.n87 163.367
R858 B.n188 B.n187 163.367
R859 B.n189 B.n188 163.367
R860 B.n189 B.n85 163.367
R861 B.n193 B.n85 163.367
R862 B.n194 B.n193 163.367
R863 B.n195 B.n194 163.367
R864 B.n195 B.n81 163.367
R865 B.n200 B.n81 163.367
R866 B.n201 B.n200 163.367
R867 B.n202 B.n201 163.367
R868 B.n202 B.n79 163.367
R869 B.n206 B.n79 163.367
R870 B.n207 B.n206 163.367
R871 B.n208 B.n207 163.367
R872 B.n208 B.n77 163.367
R873 B.n212 B.n77 163.367
R874 B.n213 B.n212 163.367
R875 B.n214 B.n213 163.367
R876 B.n214 B.n75 163.367
R877 B.n218 B.n75 163.367
R878 B.n219 B.n218 163.367
R879 B.n220 B.n219 163.367
R880 B.n220 B.n73 163.367
R881 B.n224 B.n73 163.367
R882 B.n225 B.n224 163.367
R883 B.n226 B.n225 163.367
R884 B.n226 B.n71 163.367
R885 B.n230 B.n71 163.367
R886 B.n231 B.n230 163.367
R887 B.n232 B.n231 163.367
R888 B.n232 B.n69 163.367
R889 B.n236 B.n69 163.367
R890 B.n237 B.n236 163.367
R891 B.n238 B.n237 163.367
R892 B.n238 B.n67 163.367
R893 B.n242 B.n67 163.367
R894 B.n292 B.n291 163.367
R895 B.n291 B.n290 163.367
R896 B.n290 B.n51 163.367
R897 B.n286 B.n51 163.367
R898 B.n286 B.n285 163.367
R899 B.n285 B.n284 163.367
R900 B.n284 B.n53 163.367
R901 B.n280 B.n53 163.367
R902 B.n280 B.n279 163.367
R903 B.n279 B.n278 163.367
R904 B.n278 B.n55 163.367
R905 B.n274 B.n55 163.367
R906 B.n274 B.n273 163.367
R907 B.n273 B.n272 163.367
R908 B.n272 B.n57 163.367
R909 B.n268 B.n57 163.367
R910 B.n268 B.n267 163.367
R911 B.n267 B.n266 163.367
R912 B.n266 B.n59 163.367
R913 B.n262 B.n59 163.367
R914 B.n262 B.n261 163.367
R915 B.n261 B.n260 163.367
R916 B.n260 B.n61 163.367
R917 B.n256 B.n61 163.367
R918 B.n256 B.n255 163.367
R919 B.n255 B.n254 163.367
R920 B.n254 B.n63 163.367
R921 B.n250 B.n63 163.367
R922 B.n250 B.n249 163.367
R923 B.n249 B.n248 163.367
R924 B.n248 B.n65 163.367
R925 B.n244 B.n65 163.367
R926 B.n244 B.n243 163.367
R927 B.n399 B.n398 163.367
R928 B.n398 B.n11 163.367
R929 B.n394 B.n11 163.367
R930 B.n394 B.n393 163.367
R931 B.n393 B.n392 163.367
R932 B.n392 B.n13 163.367
R933 B.n388 B.n13 163.367
R934 B.n388 B.n387 163.367
R935 B.n387 B.n386 163.367
R936 B.n386 B.n15 163.367
R937 B.n382 B.n15 163.367
R938 B.n382 B.n381 163.367
R939 B.n381 B.n380 163.367
R940 B.n380 B.n17 163.367
R941 B.n376 B.n17 163.367
R942 B.n376 B.n375 163.367
R943 B.n375 B.n374 163.367
R944 B.n374 B.n19 163.367
R945 B.n370 B.n19 163.367
R946 B.n370 B.n369 163.367
R947 B.n369 B.n368 163.367
R948 B.n368 B.n21 163.367
R949 B.n364 B.n21 163.367
R950 B.n364 B.n363 163.367
R951 B.n363 B.n362 163.367
R952 B.n362 B.n23 163.367
R953 B.n358 B.n23 163.367
R954 B.n358 B.n357 163.367
R955 B.n357 B.n356 163.367
R956 B.n356 B.n25 163.367
R957 B.n351 B.n25 163.367
R958 B.n351 B.n350 163.367
R959 B.n350 B.n349 163.367
R960 B.n349 B.n29 163.367
R961 B.n345 B.n29 163.367
R962 B.n345 B.n344 163.367
R963 B.n344 B.n343 163.367
R964 B.n343 B.n31 163.367
R965 B.n339 B.n31 163.367
R966 B.n339 B.n338 163.367
R967 B.n338 B.n35 163.367
R968 B.n334 B.n35 163.367
R969 B.n334 B.n333 163.367
R970 B.n333 B.n332 163.367
R971 B.n332 B.n37 163.367
R972 B.n328 B.n37 163.367
R973 B.n328 B.n327 163.367
R974 B.n327 B.n326 163.367
R975 B.n326 B.n39 163.367
R976 B.n322 B.n39 163.367
R977 B.n322 B.n321 163.367
R978 B.n321 B.n320 163.367
R979 B.n320 B.n41 163.367
R980 B.n316 B.n41 163.367
R981 B.n316 B.n315 163.367
R982 B.n315 B.n314 163.367
R983 B.n314 B.n43 163.367
R984 B.n310 B.n43 163.367
R985 B.n310 B.n309 163.367
R986 B.n309 B.n308 163.367
R987 B.n308 B.n45 163.367
R988 B.n304 B.n45 163.367
R989 B.n304 B.n303 163.367
R990 B.n303 B.n302 163.367
R991 B.n302 B.n47 163.367
R992 B.n298 B.n47 163.367
R993 B.n298 B.n297 163.367
R994 B.n297 B.n296 163.367
R995 B.n296 B.n49 163.367
R996 B.n400 B.n9 163.367
R997 B.n404 B.n9 163.367
R998 B.n405 B.n404 163.367
R999 B.n406 B.n405 163.367
R1000 B.n406 B.n7 163.367
R1001 B.n410 B.n7 163.367
R1002 B.n411 B.n410 163.367
R1003 B.n412 B.n411 163.367
R1004 B.n412 B.n5 163.367
R1005 B.n416 B.n5 163.367
R1006 B.n417 B.n416 163.367
R1007 B.n418 B.n417 163.367
R1008 B.n418 B.n3 163.367
R1009 B.n422 B.n3 163.367
R1010 B.n423 B.n422 163.367
R1011 B.n112 B.n2 163.367
R1012 B.n113 B.n112 163.367
R1013 B.n114 B.n113 163.367
R1014 B.n114 B.n109 163.367
R1015 B.n118 B.n109 163.367
R1016 B.n119 B.n118 163.367
R1017 B.n120 B.n119 163.367
R1018 B.n120 B.n107 163.367
R1019 B.n124 B.n107 163.367
R1020 B.n125 B.n124 163.367
R1021 B.n126 B.n125 163.367
R1022 B.n126 B.n105 163.367
R1023 B.n130 B.n105 163.367
R1024 B.n131 B.n130 163.367
R1025 B.n132 B.n131 163.367
R1026 B.n179 B.n178 59.5399
R1027 B.n197 B.n83 59.5399
R1028 B.n34 B.n33 59.5399
R1029 B.n354 B.n27 59.5399
R1030 B.n401 B.n10 33.8737
R1031 B.n294 B.n293 33.8737
R1032 B.n241 B.n66 33.8737
R1033 B.n134 B.n133 33.8737
R1034 B B.n425 18.0485
R1035 B.n178 B.n177 14.1581
R1036 B.n83 B.n82 14.1581
R1037 B.n33 B.n32 14.1581
R1038 B.n27 B.n26 14.1581
R1039 B.n402 B.n401 10.6151
R1040 B.n403 B.n402 10.6151
R1041 B.n403 B.n8 10.6151
R1042 B.n407 B.n8 10.6151
R1043 B.n408 B.n407 10.6151
R1044 B.n409 B.n408 10.6151
R1045 B.n409 B.n6 10.6151
R1046 B.n413 B.n6 10.6151
R1047 B.n414 B.n413 10.6151
R1048 B.n415 B.n414 10.6151
R1049 B.n415 B.n4 10.6151
R1050 B.n419 B.n4 10.6151
R1051 B.n420 B.n419 10.6151
R1052 B.n421 B.n420 10.6151
R1053 B.n421 B.n0 10.6151
R1054 B.n397 B.n10 10.6151
R1055 B.n397 B.n396 10.6151
R1056 B.n396 B.n395 10.6151
R1057 B.n395 B.n12 10.6151
R1058 B.n391 B.n12 10.6151
R1059 B.n391 B.n390 10.6151
R1060 B.n390 B.n389 10.6151
R1061 B.n389 B.n14 10.6151
R1062 B.n385 B.n14 10.6151
R1063 B.n385 B.n384 10.6151
R1064 B.n384 B.n383 10.6151
R1065 B.n383 B.n16 10.6151
R1066 B.n379 B.n16 10.6151
R1067 B.n379 B.n378 10.6151
R1068 B.n378 B.n377 10.6151
R1069 B.n377 B.n18 10.6151
R1070 B.n373 B.n18 10.6151
R1071 B.n373 B.n372 10.6151
R1072 B.n372 B.n371 10.6151
R1073 B.n371 B.n20 10.6151
R1074 B.n367 B.n20 10.6151
R1075 B.n367 B.n366 10.6151
R1076 B.n366 B.n365 10.6151
R1077 B.n365 B.n22 10.6151
R1078 B.n361 B.n22 10.6151
R1079 B.n361 B.n360 10.6151
R1080 B.n360 B.n359 10.6151
R1081 B.n359 B.n24 10.6151
R1082 B.n355 B.n24 10.6151
R1083 B.n353 B.n352 10.6151
R1084 B.n352 B.n28 10.6151
R1085 B.n348 B.n28 10.6151
R1086 B.n348 B.n347 10.6151
R1087 B.n347 B.n346 10.6151
R1088 B.n346 B.n30 10.6151
R1089 B.n342 B.n30 10.6151
R1090 B.n342 B.n341 10.6151
R1091 B.n341 B.n340 10.6151
R1092 B.n337 B.n336 10.6151
R1093 B.n336 B.n335 10.6151
R1094 B.n335 B.n36 10.6151
R1095 B.n331 B.n36 10.6151
R1096 B.n331 B.n330 10.6151
R1097 B.n330 B.n329 10.6151
R1098 B.n329 B.n38 10.6151
R1099 B.n325 B.n38 10.6151
R1100 B.n325 B.n324 10.6151
R1101 B.n324 B.n323 10.6151
R1102 B.n323 B.n40 10.6151
R1103 B.n319 B.n40 10.6151
R1104 B.n319 B.n318 10.6151
R1105 B.n318 B.n317 10.6151
R1106 B.n317 B.n42 10.6151
R1107 B.n313 B.n42 10.6151
R1108 B.n313 B.n312 10.6151
R1109 B.n312 B.n311 10.6151
R1110 B.n311 B.n44 10.6151
R1111 B.n307 B.n44 10.6151
R1112 B.n307 B.n306 10.6151
R1113 B.n306 B.n305 10.6151
R1114 B.n305 B.n46 10.6151
R1115 B.n301 B.n46 10.6151
R1116 B.n301 B.n300 10.6151
R1117 B.n300 B.n299 10.6151
R1118 B.n299 B.n48 10.6151
R1119 B.n295 B.n48 10.6151
R1120 B.n295 B.n294 10.6151
R1121 B.n293 B.n50 10.6151
R1122 B.n289 B.n50 10.6151
R1123 B.n289 B.n288 10.6151
R1124 B.n288 B.n287 10.6151
R1125 B.n287 B.n52 10.6151
R1126 B.n283 B.n52 10.6151
R1127 B.n283 B.n282 10.6151
R1128 B.n282 B.n281 10.6151
R1129 B.n281 B.n54 10.6151
R1130 B.n277 B.n54 10.6151
R1131 B.n277 B.n276 10.6151
R1132 B.n276 B.n275 10.6151
R1133 B.n275 B.n56 10.6151
R1134 B.n271 B.n56 10.6151
R1135 B.n271 B.n270 10.6151
R1136 B.n270 B.n269 10.6151
R1137 B.n269 B.n58 10.6151
R1138 B.n265 B.n58 10.6151
R1139 B.n265 B.n264 10.6151
R1140 B.n264 B.n263 10.6151
R1141 B.n263 B.n60 10.6151
R1142 B.n259 B.n60 10.6151
R1143 B.n259 B.n258 10.6151
R1144 B.n258 B.n257 10.6151
R1145 B.n257 B.n62 10.6151
R1146 B.n253 B.n62 10.6151
R1147 B.n253 B.n252 10.6151
R1148 B.n252 B.n251 10.6151
R1149 B.n251 B.n64 10.6151
R1150 B.n247 B.n64 10.6151
R1151 B.n247 B.n246 10.6151
R1152 B.n246 B.n245 10.6151
R1153 B.n245 B.n66 10.6151
R1154 B.n111 B.n1 10.6151
R1155 B.n111 B.n110 10.6151
R1156 B.n115 B.n110 10.6151
R1157 B.n116 B.n115 10.6151
R1158 B.n117 B.n116 10.6151
R1159 B.n117 B.n108 10.6151
R1160 B.n121 B.n108 10.6151
R1161 B.n122 B.n121 10.6151
R1162 B.n123 B.n122 10.6151
R1163 B.n123 B.n106 10.6151
R1164 B.n127 B.n106 10.6151
R1165 B.n128 B.n127 10.6151
R1166 B.n129 B.n128 10.6151
R1167 B.n129 B.n104 10.6151
R1168 B.n133 B.n104 10.6151
R1169 B.n135 B.n134 10.6151
R1170 B.n135 B.n102 10.6151
R1171 B.n139 B.n102 10.6151
R1172 B.n140 B.n139 10.6151
R1173 B.n141 B.n140 10.6151
R1174 B.n141 B.n100 10.6151
R1175 B.n145 B.n100 10.6151
R1176 B.n146 B.n145 10.6151
R1177 B.n147 B.n146 10.6151
R1178 B.n147 B.n98 10.6151
R1179 B.n151 B.n98 10.6151
R1180 B.n152 B.n151 10.6151
R1181 B.n153 B.n152 10.6151
R1182 B.n153 B.n96 10.6151
R1183 B.n157 B.n96 10.6151
R1184 B.n158 B.n157 10.6151
R1185 B.n159 B.n158 10.6151
R1186 B.n159 B.n94 10.6151
R1187 B.n163 B.n94 10.6151
R1188 B.n164 B.n163 10.6151
R1189 B.n165 B.n164 10.6151
R1190 B.n165 B.n92 10.6151
R1191 B.n169 B.n92 10.6151
R1192 B.n170 B.n169 10.6151
R1193 B.n171 B.n170 10.6151
R1194 B.n171 B.n90 10.6151
R1195 B.n175 B.n90 10.6151
R1196 B.n176 B.n175 10.6151
R1197 B.n180 B.n176 10.6151
R1198 B.n184 B.n88 10.6151
R1199 B.n185 B.n184 10.6151
R1200 B.n186 B.n185 10.6151
R1201 B.n186 B.n86 10.6151
R1202 B.n190 B.n86 10.6151
R1203 B.n191 B.n190 10.6151
R1204 B.n192 B.n191 10.6151
R1205 B.n192 B.n84 10.6151
R1206 B.n196 B.n84 10.6151
R1207 B.n199 B.n198 10.6151
R1208 B.n199 B.n80 10.6151
R1209 B.n203 B.n80 10.6151
R1210 B.n204 B.n203 10.6151
R1211 B.n205 B.n204 10.6151
R1212 B.n205 B.n78 10.6151
R1213 B.n209 B.n78 10.6151
R1214 B.n210 B.n209 10.6151
R1215 B.n211 B.n210 10.6151
R1216 B.n211 B.n76 10.6151
R1217 B.n215 B.n76 10.6151
R1218 B.n216 B.n215 10.6151
R1219 B.n217 B.n216 10.6151
R1220 B.n217 B.n74 10.6151
R1221 B.n221 B.n74 10.6151
R1222 B.n222 B.n221 10.6151
R1223 B.n223 B.n222 10.6151
R1224 B.n223 B.n72 10.6151
R1225 B.n227 B.n72 10.6151
R1226 B.n228 B.n227 10.6151
R1227 B.n229 B.n228 10.6151
R1228 B.n229 B.n70 10.6151
R1229 B.n233 B.n70 10.6151
R1230 B.n234 B.n233 10.6151
R1231 B.n235 B.n234 10.6151
R1232 B.n235 B.n68 10.6151
R1233 B.n239 B.n68 10.6151
R1234 B.n240 B.n239 10.6151
R1235 B.n241 B.n240 10.6151
R1236 B.n355 B.n354 9.36635
R1237 B.n337 B.n34 9.36635
R1238 B.n180 B.n179 9.36635
R1239 B.n198 B.n197 9.36635
R1240 B.n425 B.n0 8.11757
R1241 B.n425 B.n1 8.11757
R1242 B.n354 B.n353 1.24928
R1243 B.n340 B.n34 1.24928
R1244 B.n179 B.n88 1.24928
R1245 B.n197 B.n196 1.24928
C0 VDD2 VTAIL 8.94442f
C1 VDD2 VDD1 0.603387f
C2 VTAIL VDD1 8.9111f
C3 w_n1554_n2588# VN 2.33413f
C4 w_n1554_n2588# B 5.54799f
C5 VN VDD2 2.26463f
C6 VN VTAIL 2.00933f
C7 w_n1554_n2588# VP 2.52891f
C8 VN VDD1 0.148056f
C9 VDD2 B 1.21045f
C10 B VTAIL 1.84721f
C11 B VDD1 1.1882f
C12 VDD2 VP 0.272011f
C13 VP VTAIL 2.02384f
C14 VP VDD1 2.38515f
C15 VN B 0.654967f
C16 w_n1554_n2588# VDD2 1.44814f
C17 w_n1554_n2588# VTAIL 2.32829f
C18 VN VP 4.06399f
C19 w_n1554_n2588# VDD1 1.4332f
C20 VP B 0.969095f
C21 VDD2 VSUBS 1.159509f
C22 VDD1 VSUBS 0.918781f
C23 VTAIL VSUBS 0.531808f
C24 VN VSUBS 4.05547f
C25 VP VSUBS 1.102124f
C26 B VSUBS 2.115948f
C27 w_n1554_n2588# VSUBS 49.8834f
C28 B.n0 VSUBS 0.0054f
C29 B.n1 VSUBS 0.0054f
C30 B.n2 VSUBS 0.007986f
C31 B.n3 VSUBS 0.00612f
C32 B.n4 VSUBS 0.00612f
C33 B.n5 VSUBS 0.00612f
C34 B.n6 VSUBS 0.00612f
C35 B.n7 VSUBS 0.00612f
C36 B.n8 VSUBS 0.00612f
C37 B.n9 VSUBS 0.00612f
C38 B.n10 VSUBS 0.015155f
C39 B.n11 VSUBS 0.00612f
C40 B.n12 VSUBS 0.00612f
C41 B.n13 VSUBS 0.00612f
C42 B.n14 VSUBS 0.00612f
C43 B.n15 VSUBS 0.00612f
C44 B.n16 VSUBS 0.00612f
C45 B.n17 VSUBS 0.00612f
C46 B.n18 VSUBS 0.00612f
C47 B.n19 VSUBS 0.00612f
C48 B.n20 VSUBS 0.00612f
C49 B.n21 VSUBS 0.00612f
C50 B.n22 VSUBS 0.00612f
C51 B.n23 VSUBS 0.00612f
C52 B.n24 VSUBS 0.00612f
C53 B.n25 VSUBS 0.00612f
C54 B.t10 VSUBS 0.112604f
C55 B.t11 VSUBS 0.119338f
C56 B.t9 VSUBS 0.115279f
C57 B.n26 VSUBS 0.182398f
C58 B.n27 VSUBS 0.160826f
C59 B.n28 VSUBS 0.00612f
C60 B.n29 VSUBS 0.00612f
C61 B.n30 VSUBS 0.00612f
C62 B.n31 VSUBS 0.00612f
C63 B.t1 VSUBS 0.112606f
C64 B.t2 VSUBS 0.11934f
C65 B.t0 VSUBS 0.115279f
C66 B.n32 VSUBS 0.182396f
C67 B.n33 VSUBS 0.160824f
C68 B.n34 VSUBS 0.01418f
C69 B.n35 VSUBS 0.00612f
C70 B.n36 VSUBS 0.00612f
C71 B.n37 VSUBS 0.00612f
C72 B.n38 VSUBS 0.00612f
C73 B.n39 VSUBS 0.00612f
C74 B.n40 VSUBS 0.00612f
C75 B.n41 VSUBS 0.00612f
C76 B.n42 VSUBS 0.00612f
C77 B.n43 VSUBS 0.00612f
C78 B.n44 VSUBS 0.00612f
C79 B.n45 VSUBS 0.00612f
C80 B.n46 VSUBS 0.00612f
C81 B.n47 VSUBS 0.00612f
C82 B.n48 VSUBS 0.00612f
C83 B.n49 VSUBS 0.015155f
C84 B.n50 VSUBS 0.00612f
C85 B.n51 VSUBS 0.00612f
C86 B.n52 VSUBS 0.00612f
C87 B.n53 VSUBS 0.00612f
C88 B.n54 VSUBS 0.00612f
C89 B.n55 VSUBS 0.00612f
C90 B.n56 VSUBS 0.00612f
C91 B.n57 VSUBS 0.00612f
C92 B.n58 VSUBS 0.00612f
C93 B.n59 VSUBS 0.00612f
C94 B.n60 VSUBS 0.00612f
C95 B.n61 VSUBS 0.00612f
C96 B.n62 VSUBS 0.00612f
C97 B.n63 VSUBS 0.00612f
C98 B.n64 VSUBS 0.00612f
C99 B.n65 VSUBS 0.00612f
C100 B.n66 VSUBS 0.014883f
C101 B.n67 VSUBS 0.00612f
C102 B.n68 VSUBS 0.00612f
C103 B.n69 VSUBS 0.00612f
C104 B.n70 VSUBS 0.00612f
C105 B.n71 VSUBS 0.00612f
C106 B.n72 VSUBS 0.00612f
C107 B.n73 VSUBS 0.00612f
C108 B.n74 VSUBS 0.00612f
C109 B.n75 VSUBS 0.00612f
C110 B.n76 VSUBS 0.00612f
C111 B.n77 VSUBS 0.00612f
C112 B.n78 VSUBS 0.00612f
C113 B.n79 VSUBS 0.00612f
C114 B.n80 VSUBS 0.00612f
C115 B.n81 VSUBS 0.00612f
C116 B.t8 VSUBS 0.112606f
C117 B.t7 VSUBS 0.11934f
C118 B.t6 VSUBS 0.115279f
C119 B.n82 VSUBS 0.182396f
C120 B.n83 VSUBS 0.160824f
C121 B.n84 VSUBS 0.00612f
C122 B.n85 VSUBS 0.00612f
C123 B.n86 VSUBS 0.00612f
C124 B.n87 VSUBS 0.00612f
C125 B.n88 VSUBS 0.00342f
C126 B.n89 VSUBS 0.00612f
C127 B.n90 VSUBS 0.00612f
C128 B.n91 VSUBS 0.00612f
C129 B.n92 VSUBS 0.00612f
C130 B.n93 VSUBS 0.00612f
C131 B.n94 VSUBS 0.00612f
C132 B.n95 VSUBS 0.00612f
C133 B.n96 VSUBS 0.00612f
C134 B.n97 VSUBS 0.00612f
C135 B.n98 VSUBS 0.00612f
C136 B.n99 VSUBS 0.00612f
C137 B.n100 VSUBS 0.00612f
C138 B.n101 VSUBS 0.00612f
C139 B.n102 VSUBS 0.00612f
C140 B.n103 VSUBS 0.015155f
C141 B.n104 VSUBS 0.00612f
C142 B.n105 VSUBS 0.00612f
C143 B.n106 VSUBS 0.00612f
C144 B.n107 VSUBS 0.00612f
C145 B.n108 VSUBS 0.00612f
C146 B.n109 VSUBS 0.00612f
C147 B.n110 VSUBS 0.00612f
C148 B.n111 VSUBS 0.00612f
C149 B.n112 VSUBS 0.00612f
C150 B.n113 VSUBS 0.00612f
C151 B.n114 VSUBS 0.00612f
C152 B.n115 VSUBS 0.00612f
C153 B.n116 VSUBS 0.00612f
C154 B.n117 VSUBS 0.00612f
C155 B.n118 VSUBS 0.00612f
C156 B.n119 VSUBS 0.00612f
C157 B.n120 VSUBS 0.00612f
C158 B.n121 VSUBS 0.00612f
C159 B.n122 VSUBS 0.00612f
C160 B.n123 VSUBS 0.00612f
C161 B.n124 VSUBS 0.00612f
C162 B.n125 VSUBS 0.00612f
C163 B.n126 VSUBS 0.00612f
C164 B.n127 VSUBS 0.00612f
C165 B.n128 VSUBS 0.00612f
C166 B.n129 VSUBS 0.00612f
C167 B.n130 VSUBS 0.00612f
C168 B.n131 VSUBS 0.00612f
C169 B.n132 VSUBS 0.014186f
C170 B.n133 VSUBS 0.014186f
C171 B.n134 VSUBS 0.015155f
C172 B.n135 VSUBS 0.00612f
C173 B.n136 VSUBS 0.00612f
C174 B.n137 VSUBS 0.00612f
C175 B.n138 VSUBS 0.00612f
C176 B.n139 VSUBS 0.00612f
C177 B.n140 VSUBS 0.00612f
C178 B.n141 VSUBS 0.00612f
C179 B.n142 VSUBS 0.00612f
C180 B.n143 VSUBS 0.00612f
C181 B.n144 VSUBS 0.00612f
C182 B.n145 VSUBS 0.00612f
C183 B.n146 VSUBS 0.00612f
C184 B.n147 VSUBS 0.00612f
C185 B.n148 VSUBS 0.00612f
C186 B.n149 VSUBS 0.00612f
C187 B.n150 VSUBS 0.00612f
C188 B.n151 VSUBS 0.00612f
C189 B.n152 VSUBS 0.00612f
C190 B.n153 VSUBS 0.00612f
C191 B.n154 VSUBS 0.00612f
C192 B.n155 VSUBS 0.00612f
C193 B.n156 VSUBS 0.00612f
C194 B.n157 VSUBS 0.00612f
C195 B.n158 VSUBS 0.00612f
C196 B.n159 VSUBS 0.00612f
C197 B.n160 VSUBS 0.00612f
C198 B.n161 VSUBS 0.00612f
C199 B.n162 VSUBS 0.00612f
C200 B.n163 VSUBS 0.00612f
C201 B.n164 VSUBS 0.00612f
C202 B.n165 VSUBS 0.00612f
C203 B.n166 VSUBS 0.00612f
C204 B.n167 VSUBS 0.00612f
C205 B.n168 VSUBS 0.00612f
C206 B.n169 VSUBS 0.00612f
C207 B.n170 VSUBS 0.00612f
C208 B.n171 VSUBS 0.00612f
C209 B.n172 VSUBS 0.00612f
C210 B.n173 VSUBS 0.00612f
C211 B.n174 VSUBS 0.00612f
C212 B.n175 VSUBS 0.00612f
C213 B.n176 VSUBS 0.00612f
C214 B.t5 VSUBS 0.112604f
C215 B.t4 VSUBS 0.119338f
C216 B.t3 VSUBS 0.115279f
C217 B.n177 VSUBS 0.182398f
C218 B.n178 VSUBS 0.160826f
C219 B.n179 VSUBS 0.01418f
C220 B.n180 VSUBS 0.00576f
C221 B.n181 VSUBS 0.00612f
C222 B.n182 VSUBS 0.00612f
C223 B.n183 VSUBS 0.00612f
C224 B.n184 VSUBS 0.00612f
C225 B.n185 VSUBS 0.00612f
C226 B.n186 VSUBS 0.00612f
C227 B.n187 VSUBS 0.00612f
C228 B.n188 VSUBS 0.00612f
C229 B.n189 VSUBS 0.00612f
C230 B.n190 VSUBS 0.00612f
C231 B.n191 VSUBS 0.00612f
C232 B.n192 VSUBS 0.00612f
C233 B.n193 VSUBS 0.00612f
C234 B.n194 VSUBS 0.00612f
C235 B.n195 VSUBS 0.00612f
C236 B.n196 VSUBS 0.00342f
C237 B.n197 VSUBS 0.01418f
C238 B.n198 VSUBS 0.00576f
C239 B.n199 VSUBS 0.00612f
C240 B.n200 VSUBS 0.00612f
C241 B.n201 VSUBS 0.00612f
C242 B.n202 VSUBS 0.00612f
C243 B.n203 VSUBS 0.00612f
C244 B.n204 VSUBS 0.00612f
C245 B.n205 VSUBS 0.00612f
C246 B.n206 VSUBS 0.00612f
C247 B.n207 VSUBS 0.00612f
C248 B.n208 VSUBS 0.00612f
C249 B.n209 VSUBS 0.00612f
C250 B.n210 VSUBS 0.00612f
C251 B.n211 VSUBS 0.00612f
C252 B.n212 VSUBS 0.00612f
C253 B.n213 VSUBS 0.00612f
C254 B.n214 VSUBS 0.00612f
C255 B.n215 VSUBS 0.00612f
C256 B.n216 VSUBS 0.00612f
C257 B.n217 VSUBS 0.00612f
C258 B.n218 VSUBS 0.00612f
C259 B.n219 VSUBS 0.00612f
C260 B.n220 VSUBS 0.00612f
C261 B.n221 VSUBS 0.00612f
C262 B.n222 VSUBS 0.00612f
C263 B.n223 VSUBS 0.00612f
C264 B.n224 VSUBS 0.00612f
C265 B.n225 VSUBS 0.00612f
C266 B.n226 VSUBS 0.00612f
C267 B.n227 VSUBS 0.00612f
C268 B.n228 VSUBS 0.00612f
C269 B.n229 VSUBS 0.00612f
C270 B.n230 VSUBS 0.00612f
C271 B.n231 VSUBS 0.00612f
C272 B.n232 VSUBS 0.00612f
C273 B.n233 VSUBS 0.00612f
C274 B.n234 VSUBS 0.00612f
C275 B.n235 VSUBS 0.00612f
C276 B.n236 VSUBS 0.00612f
C277 B.n237 VSUBS 0.00612f
C278 B.n238 VSUBS 0.00612f
C279 B.n239 VSUBS 0.00612f
C280 B.n240 VSUBS 0.00612f
C281 B.n241 VSUBS 0.014458f
C282 B.n242 VSUBS 0.015155f
C283 B.n243 VSUBS 0.014186f
C284 B.n244 VSUBS 0.00612f
C285 B.n245 VSUBS 0.00612f
C286 B.n246 VSUBS 0.00612f
C287 B.n247 VSUBS 0.00612f
C288 B.n248 VSUBS 0.00612f
C289 B.n249 VSUBS 0.00612f
C290 B.n250 VSUBS 0.00612f
C291 B.n251 VSUBS 0.00612f
C292 B.n252 VSUBS 0.00612f
C293 B.n253 VSUBS 0.00612f
C294 B.n254 VSUBS 0.00612f
C295 B.n255 VSUBS 0.00612f
C296 B.n256 VSUBS 0.00612f
C297 B.n257 VSUBS 0.00612f
C298 B.n258 VSUBS 0.00612f
C299 B.n259 VSUBS 0.00612f
C300 B.n260 VSUBS 0.00612f
C301 B.n261 VSUBS 0.00612f
C302 B.n262 VSUBS 0.00612f
C303 B.n263 VSUBS 0.00612f
C304 B.n264 VSUBS 0.00612f
C305 B.n265 VSUBS 0.00612f
C306 B.n266 VSUBS 0.00612f
C307 B.n267 VSUBS 0.00612f
C308 B.n268 VSUBS 0.00612f
C309 B.n269 VSUBS 0.00612f
C310 B.n270 VSUBS 0.00612f
C311 B.n271 VSUBS 0.00612f
C312 B.n272 VSUBS 0.00612f
C313 B.n273 VSUBS 0.00612f
C314 B.n274 VSUBS 0.00612f
C315 B.n275 VSUBS 0.00612f
C316 B.n276 VSUBS 0.00612f
C317 B.n277 VSUBS 0.00612f
C318 B.n278 VSUBS 0.00612f
C319 B.n279 VSUBS 0.00612f
C320 B.n280 VSUBS 0.00612f
C321 B.n281 VSUBS 0.00612f
C322 B.n282 VSUBS 0.00612f
C323 B.n283 VSUBS 0.00612f
C324 B.n284 VSUBS 0.00612f
C325 B.n285 VSUBS 0.00612f
C326 B.n286 VSUBS 0.00612f
C327 B.n287 VSUBS 0.00612f
C328 B.n288 VSUBS 0.00612f
C329 B.n289 VSUBS 0.00612f
C330 B.n290 VSUBS 0.00612f
C331 B.n291 VSUBS 0.00612f
C332 B.n292 VSUBS 0.014186f
C333 B.n293 VSUBS 0.014186f
C334 B.n294 VSUBS 0.015155f
C335 B.n295 VSUBS 0.00612f
C336 B.n296 VSUBS 0.00612f
C337 B.n297 VSUBS 0.00612f
C338 B.n298 VSUBS 0.00612f
C339 B.n299 VSUBS 0.00612f
C340 B.n300 VSUBS 0.00612f
C341 B.n301 VSUBS 0.00612f
C342 B.n302 VSUBS 0.00612f
C343 B.n303 VSUBS 0.00612f
C344 B.n304 VSUBS 0.00612f
C345 B.n305 VSUBS 0.00612f
C346 B.n306 VSUBS 0.00612f
C347 B.n307 VSUBS 0.00612f
C348 B.n308 VSUBS 0.00612f
C349 B.n309 VSUBS 0.00612f
C350 B.n310 VSUBS 0.00612f
C351 B.n311 VSUBS 0.00612f
C352 B.n312 VSUBS 0.00612f
C353 B.n313 VSUBS 0.00612f
C354 B.n314 VSUBS 0.00612f
C355 B.n315 VSUBS 0.00612f
C356 B.n316 VSUBS 0.00612f
C357 B.n317 VSUBS 0.00612f
C358 B.n318 VSUBS 0.00612f
C359 B.n319 VSUBS 0.00612f
C360 B.n320 VSUBS 0.00612f
C361 B.n321 VSUBS 0.00612f
C362 B.n322 VSUBS 0.00612f
C363 B.n323 VSUBS 0.00612f
C364 B.n324 VSUBS 0.00612f
C365 B.n325 VSUBS 0.00612f
C366 B.n326 VSUBS 0.00612f
C367 B.n327 VSUBS 0.00612f
C368 B.n328 VSUBS 0.00612f
C369 B.n329 VSUBS 0.00612f
C370 B.n330 VSUBS 0.00612f
C371 B.n331 VSUBS 0.00612f
C372 B.n332 VSUBS 0.00612f
C373 B.n333 VSUBS 0.00612f
C374 B.n334 VSUBS 0.00612f
C375 B.n335 VSUBS 0.00612f
C376 B.n336 VSUBS 0.00612f
C377 B.n337 VSUBS 0.00576f
C378 B.n338 VSUBS 0.00612f
C379 B.n339 VSUBS 0.00612f
C380 B.n340 VSUBS 0.00342f
C381 B.n341 VSUBS 0.00612f
C382 B.n342 VSUBS 0.00612f
C383 B.n343 VSUBS 0.00612f
C384 B.n344 VSUBS 0.00612f
C385 B.n345 VSUBS 0.00612f
C386 B.n346 VSUBS 0.00612f
C387 B.n347 VSUBS 0.00612f
C388 B.n348 VSUBS 0.00612f
C389 B.n349 VSUBS 0.00612f
C390 B.n350 VSUBS 0.00612f
C391 B.n351 VSUBS 0.00612f
C392 B.n352 VSUBS 0.00612f
C393 B.n353 VSUBS 0.00342f
C394 B.n354 VSUBS 0.01418f
C395 B.n355 VSUBS 0.00576f
C396 B.n356 VSUBS 0.00612f
C397 B.n357 VSUBS 0.00612f
C398 B.n358 VSUBS 0.00612f
C399 B.n359 VSUBS 0.00612f
C400 B.n360 VSUBS 0.00612f
C401 B.n361 VSUBS 0.00612f
C402 B.n362 VSUBS 0.00612f
C403 B.n363 VSUBS 0.00612f
C404 B.n364 VSUBS 0.00612f
C405 B.n365 VSUBS 0.00612f
C406 B.n366 VSUBS 0.00612f
C407 B.n367 VSUBS 0.00612f
C408 B.n368 VSUBS 0.00612f
C409 B.n369 VSUBS 0.00612f
C410 B.n370 VSUBS 0.00612f
C411 B.n371 VSUBS 0.00612f
C412 B.n372 VSUBS 0.00612f
C413 B.n373 VSUBS 0.00612f
C414 B.n374 VSUBS 0.00612f
C415 B.n375 VSUBS 0.00612f
C416 B.n376 VSUBS 0.00612f
C417 B.n377 VSUBS 0.00612f
C418 B.n378 VSUBS 0.00612f
C419 B.n379 VSUBS 0.00612f
C420 B.n380 VSUBS 0.00612f
C421 B.n381 VSUBS 0.00612f
C422 B.n382 VSUBS 0.00612f
C423 B.n383 VSUBS 0.00612f
C424 B.n384 VSUBS 0.00612f
C425 B.n385 VSUBS 0.00612f
C426 B.n386 VSUBS 0.00612f
C427 B.n387 VSUBS 0.00612f
C428 B.n388 VSUBS 0.00612f
C429 B.n389 VSUBS 0.00612f
C430 B.n390 VSUBS 0.00612f
C431 B.n391 VSUBS 0.00612f
C432 B.n392 VSUBS 0.00612f
C433 B.n393 VSUBS 0.00612f
C434 B.n394 VSUBS 0.00612f
C435 B.n395 VSUBS 0.00612f
C436 B.n396 VSUBS 0.00612f
C437 B.n397 VSUBS 0.00612f
C438 B.n398 VSUBS 0.00612f
C439 B.n399 VSUBS 0.015155f
C440 B.n400 VSUBS 0.014186f
C441 B.n401 VSUBS 0.014186f
C442 B.n402 VSUBS 0.00612f
C443 B.n403 VSUBS 0.00612f
C444 B.n404 VSUBS 0.00612f
C445 B.n405 VSUBS 0.00612f
C446 B.n406 VSUBS 0.00612f
C447 B.n407 VSUBS 0.00612f
C448 B.n408 VSUBS 0.00612f
C449 B.n409 VSUBS 0.00612f
C450 B.n410 VSUBS 0.00612f
C451 B.n411 VSUBS 0.00612f
C452 B.n412 VSUBS 0.00612f
C453 B.n413 VSUBS 0.00612f
C454 B.n414 VSUBS 0.00612f
C455 B.n415 VSUBS 0.00612f
C456 B.n416 VSUBS 0.00612f
C457 B.n417 VSUBS 0.00612f
C458 B.n418 VSUBS 0.00612f
C459 B.n419 VSUBS 0.00612f
C460 B.n420 VSUBS 0.00612f
C461 B.n421 VSUBS 0.00612f
C462 B.n422 VSUBS 0.00612f
C463 B.n423 VSUBS 0.007986f
C464 B.n424 VSUBS 0.008508f
C465 B.n425 VSUBS 0.016918f
C466 VDD1.n0 VSUBS 0.028947f
C467 VDD1.n1 VSUBS 0.025844f
C468 VDD1.n2 VSUBS 0.013888f
C469 VDD1.n3 VSUBS 0.032825f
C470 VDD1.n4 VSUBS 0.014704f
C471 VDD1.n5 VSUBS 0.025844f
C472 VDD1.n6 VSUBS 0.013888f
C473 VDD1.n7 VSUBS 0.032825f
C474 VDD1.n8 VSUBS 0.014704f
C475 VDD1.n9 VSUBS 0.025844f
C476 VDD1.n10 VSUBS 0.013888f
C477 VDD1.n11 VSUBS 0.032825f
C478 VDD1.n12 VSUBS 0.014704f
C479 VDD1.n13 VSUBS 0.129751f
C480 VDD1.t1 VSUBS 0.07f
C481 VDD1.n14 VSUBS 0.024619f
C482 VDD1.n15 VSUBS 0.020881f
C483 VDD1.n16 VSUBS 0.013888f
C484 VDD1.n17 VSUBS 0.840315f
C485 VDD1.n18 VSUBS 0.025844f
C486 VDD1.n19 VSUBS 0.013888f
C487 VDD1.n20 VSUBS 0.014704f
C488 VDD1.n21 VSUBS 0.032825f
C489 VDD1.n22 VSUBS 0.032825f
C490 VDD1.n23 VSUBS 0.014704f
C491 VDD1.n24 VSUBS 0.013888f
C492 VDD1.n25 VSUBS 0.025844f
C493 VDD1.n26 VSUBS 0.025844f
C494 VDD1.n27 VSUBS 0.013888f
C495 VDD1.n28 VSUBS 0.014704f
C496 VDD1.n29 VSUBS 0.032825f
C497 VDD1.n30 VSUBS 0.032825f
C498 VDD1.n31 VSUBS 0.014704f
C499 VDD1.n32 VSUBS 0.013888f
C500 VDD1.n33 VSUBS 0.025844f
C501 VDD1.n34 VSUBS 0.025844f
C502 VDD1.n35 VSUBS 0.013888f
C503 VDD1.n36 VSUBS 0.014704f
C504 VDD1.n37 VSUBS 0.032825f
C505 VDD1.n38 VSUBS 0.081337f
C506 VDD1.n39 VSUBS 0.014704f
C507 VDD1.n40 VSUBS 0.013888f
C508 VDD1.n41 VSUBS 0.057619f
C509 VDD1.n42 VSUBS 0.059802f
C510 VDD1.n43 VSUBS 0.028947f
C511 VDD1.n44 VSUBS 0.025844f
C512 VDD1.n45 VSUBS 0.013888f
C513 VDD1.n46 VSUBS 0.032825f
C514 VDD1.n47 VSUBS 0.014704f
C515 VDD1.n48 VSUBS 0.025844f
C516 VDD1.n49 VSUBS 0.013888f
C517 VDD1.n50 VSUBS 0.032825f
C518 VDD1.n51 VSUBS 0.014704f
C519 VDD1.n52 VSUBS 0.025844f
C520 VDD1.n53 VSUBS 0.013888f
C521 VDD1.n54 VSUBS 0.032825f
C522 VDD1.n55 VSUBS 0.014704f
C523 VDD1.n56 VSUBS 0.129751f
C524 VDD1.t0 VSUBS 0.07f
C525 VDD1.n57 VSUBS 0.024619f
C526 VDD1.n58 VSUBS 0.020881f
C527 VDD1.n59 VSUBS 0.013888f
C528 VDD1.n60 VSUBS 0.840315f
C529 VDD1.n61 VSUBS 0.025844f
C530 VDD1.n62 VSUBS 0.013888f
C531 VDD1.n63 VSUBS 0.014704f
C532 VDD1.n64 VSUBS 0.032825f
C533 VDD1.n65 VSUBS 0.032825f
C534 VDD1.n66 VSUBS 0.014704f
C535 VDD1.n67 VSUBS 0.013888f
C536 VDD1.n68 VSUBS 0.025844f
C537 VDD1.n69 VSUBS 0.025844f
C538 VDD1.n70 VSUBS 0.013888f
C539 VDD1.n71 VSUBS 0.014704f
C540 VDD1.n72 VSUBS 0.032825f
C541 VDD1.n73 VSUBS 0.032825f
C542 VDD1.n74 VSUBS 0.014704f
C543 VDD1.n75 VSUBS 0.013888f
C544 VDD1.n76 VSUBS 0.025844f
C545 VDD1.n77 VSUBS 0.025844f
C546 VDD1.n78 VSUBS 0.013888f
C547 VDD1.n79 VSUBS 0.014704f
C548 VDD1.n80 VSUBS 0.032825f
C549 VDD1.n81 VSUBS 0.081337f
C550 VDD1.n82 VSUBS 0.014704f
C551 VDD1.n83 VSUBS 0.013888f
C552 VDD1.n84 VSUBS 0.057619f
C553 VDD1.n85 VSUBS 0.059516f
C554 VDD1.t2 VSUBS 0.165425f
C555 VDD1.t3 VSUBS 0.165425f
C556 VDD1.n86 VSUBS 1.18098f
C557 VDD1.n87 VSUBS 1.85531f
C558 VDD1.t4 VSUBS 0.165425f
C559 VDD1.t5 VSUBS 0.165425f
C560 VDD1.n88 VSUBS 1.18032f
C561 VDD1.n89 VSUBS 2.17021f
C562 VP.n0 VSUBS 0.071889f
C563 VP.t5 VSUBS 0.671753f
C564 VP.t4 VSUBS 0.681081f
C565 VP.n1 VSUBS 0.285858f
C566 VP.t1 VSUBS 0.669672f
C567 VP.n2 VSUBS 0.307377f
C568 VP.t0 VSUBS 0.671753f
C569 VP.n3 VSUBS 0.294659f
C570 VP.n4 VSUBS 2.55472f
C571 VP.n5 VSUBS 2.46528f
C572 VP.n6 VSUBS 0.294659f
C573 VP.t3 VSUBS 0.669672f
C574 VP.n7 VSUBS 0.307377f
C575 VP.t2 VSUBS 0.671753f
C576 VP.n8 VSUBS 0.294659f
C577 VP.n9 VSUBS 0.055711f
C578 VTAIL.t4 VSUBS 0.192683f
C579 VTAIL.t9 VSUBS 0.192683f
C580 VTAIL.n0 VSUBS 1.23882f
C581 VTAIL.n1 VSUBS 0.727265f
C582 VTAIL.n2 VSUBS 0.033716f
C583 VTAIL.n3 VSUBS 0.030103f
C584 VTAIL.n4 VSUBS 0.016176f
C585 VTAIL.n5 VSUBS 0.038234f
C586 VTAIL.n6 VSUBS 0.017127f
C587 VTAIL.n7 VSUBS 0.030103f
C588 VTAIL.n8 VSUBS 0.016176f
C589 VTAIL.n9 VSUBS 0.038234f
C590 VTAIL.n10 VSUBS 0.017127f
C591 VTAIL.n11 VSUBS 0.030103f
C592 VTAIL.n12 VSUBS 0.016176f
C593 VTAIL.n13 VSUBS 0.038234f
C594 VTAIL.n14 VSUBS 0.017127f
C595 VTAIL.n15 VSUBS 0.15113f
C596 VTAIL.t2 VSUBS 0.081535f
C597 VTAIL.n16 VSUBS 0.028675f
C598 VTAIL.n17 VSUBS 0.024322f
C599 VTAIL.n18 VSUBS 0.016176f
C600 VTAIL.n19 VSUBS 0.978779f
C601 VTAIL.n20 VSUBS 0.030103f
C602 VTAIL.n21 VSUBS 0.016176f
C603 VTAIL.n22 VSUBS 0.017127f
C604 VTAIL.n23 VSUBS 0.038234f
C605 VTAIL.n24 VSUBS 0.038234f
C606 VTAIL.n25 VSUBS 0.017127f
C607 VTAIL.n26 VSUBS 0.016176f
C608 VTAIL.n27 VSUBS 0.030103f
C609 VTAIL.n28 VSUBS 0.030103f
C610 VTAIL.n29 VSUBS 0.016176f
C611 VTAIL.n30 VSUBS 0.017127f
C612 VTAIL.n31 VSUBS 0.038234f
C613 VTAIL.n32 VSUBS 0.038234f
C614 VTAIL.n33 VSUBS 0.017127f
C615 VTAIL.n34 VSUBS 0.016176f
C616 VTAIL.n35 VSUBS 0.030103f
C617 VTAIL.n36 VSUBS 0.030103f
C618 VTAIL.n37 VSUBS 0.016176f
C619 VTAIL.n38 VSUBS 0.017127f
C620 VTAIL.n39 VSUBS 0.038234f
C621 VTAIL.n40 VSUBS 0.094739f
C622 VTAIL.n41 VSUBS 0.017127f
C623 VTAIL.n42 VSUBS 0.016176f
C624 VTAIL.n43 VSUBS 0.067113f
C625 VTAIL.n44 VSUBS 0.047663f
C626 VTAIL.n45 VSUBS 0.161453f
C627 VTAIL.t11 VSUBS 0.192683f
C628 VTAIL.t3 VSUBS 0.192683f
C629 VTAIL.n46 VSUBS 1.23882f
C630 VTAIL.n47 VSUBS 1.89961f
C631 VTAIL.t8 VSUBS 0.192683f
C632 VTAIL.t7 VSUBS 0.192683f
C633 VTAIL.n48 VSUBS 1.23883f
C634 VTAIL.n49 VSUBS 1.8996f
C635 VTAIL.n50 VSUBS 0.033716f
C636 VTAIL.n51 VSUBS 0.030103f
C637 VTAIL.n52 VSUBS 0.016176f
C638 VTAIL.n53 VSUBS 0.038234f
C639 VTAIL.n54 VSUBS 0.017127f
C640 VTAIL.n55 VSUBS 0.030103f
C641 VTAIL.n56 VSUBS 0.016176f
C642 VTAIL.n57 VSUBS 0.038234f
C643 VTAIL.n58 VSUBS 0.017127f
C644 VTAIL.n59 VSUBS 0.030103f
C645 VTAIL.n60 VSUBS 0.016176f
C646 VTAIL.n61 VSUBS 0.038234f
C647 VTAIL.n62 VSUBS 0.017127f
C648 VTAIL.n63 VSUBS 0.15113f
C649 VTAIL.t5 VSUBS 0.081535f
C650 VTAIL.n64 VSUBS 0.028675f
C651 VTAIL.n65 VSUBS 0.024322f
C652 VTAIL.n66 VSUBS 0.016176f
C653 VTAIL.n67 VSUBS 0.978779f
C654 VTAIL.n68 VSUBS 0.030103f
C655 VTAIL.n69 VSUBS 0.016176f
C656 VTAIL.n70 VSUBS 0.017127f
C657 VTAIL.n71 VSUBS 0.038234f
C658 VTAIL.n72 VSUBS 0.038234f
C659 VTAIL.n73 VSUBS 0.017127f
C660 VTAIL.n74 VSUBS 0.016176f
C661 VTAIL.n75 VSUBS 0.030103f
C662 VTAIL.n76 VSUBS 0.030103f
C663 VTAIL.n77 VSUBS 0.016176f
C664 VTAIL.n78 VSUBS 0.017127f
C665 VTAIL.n79 VSUBS 0.038234f
C666 VTAIL.n80 VSUBS 0.038234f
C667 VTAIL.n81 VSUBS 0.017127f
C668 VTAIL.n82 VSUBS 0.016176f
C669 VTAIL.n83 VSUBS 0.030103f
C670 VTAIL.n84 VSUBS 0.030103f
C671 VTAIL.n85 VSUBS 0.016176f
C672 VTAIL.n86 VSUBS 0.017127f
C673 VTAIL.n87 VSUBS 0.038234f
C674 VTAIL.n88 VSUBS 0.094739f
C675 VTAIL.n89 VSUBS 0.017127f
C676 VTAIL.n90 VSUBS 0.016176f
C677 VTAIL.n91 VSUBS 0.067113f
C678 VTAIL.n92 VSUBS 0.047663f
C679 VTAIL.n93 VSUBS 0.161453f
C680 VTAIL.t10 VSUBS 0.192683f
C681 VTAIL.t1 VSUBS 0.192683f
C682 VTAIL.n94 VSUBS 1.23883f
C683 VTAIL.n95 VSUBS 0.767392f
C684 VTAIL.n96 VSUBS 0.033716f
C685 VTAIL.n97 VSUBS 0.030103f
C686 VTAIL.n98 VSUBS 0.016176f
C687 VTAIL.n99 VSUBS 0.038234f
C688 VTAIL.n100 VSUBS 0.017127f
C689 VTAIL.n101 VSUBS 0.030103f
C690 VTAIL.n102 VSUBS 0.016176f
C691 VTAIL.n103 VSUBS 0.038234f
C692 VTAIL.n104 VSUBS 0.017127f
C693 VTAIL.n105 VSUBS 0.030103f
C694 VTAIL.n106 VSUBS 0.016176f
C695 VTAIL.n107 VSUBS 0.038234f
C696 VTAIL.n108 VSUBS 0.017127f
C697 VTAIL.n109 VSUBS 0.15113f
C698 VTAIL.t0 VSUBS 0.081535f
C699 VTAIL.n110 VSUBS 0.028675f
C700 VTAIL.n111 VSUBS 0.024322f
C701 VTAIL.n112 VSUBS 0.016176f
C702 VTAIL.n113 VSUBS 0.978779f
C703 VTAIL.n114 VSUBS 0.030103f
C704 VTAIL.n115 VSUBS 0.016176f
C705 VTAIL.n116 VSUBS 0.017127f
C706 VTAIL.n117 VSUBS 0.038234f
C707 VTAIL.n118 VSUBS 0.038234f
C708 VTAIL.n119 VSUBS 0.017127f
C709 VTAIL.n120 VSUBS 0.016176f
C710 VTAIL.n121 VSUBS 0.030103f
C711 VTAIL.n122 VSUBS 0.030103f
C712 VTAIL.n123 VSUBS 0.016176f
C713 VTAIL.n124 VSUBS 0.017127f
C714 VTAIL.n125 VSUBS 0.038234f
C715 VTAIL.n126 VSUBS 0.038234f
C716 VTAIL.n127 VSUBS 0.017127f
C717 VTAIL.n128 VSUBS 0.016176f
C718 VTAIL.n129 VSUBS 0.030103f
C719 VTAIL.n130 VSUBS 0.030103f
C720 VTAIL.n131 VSUBS 0.016176f
C721 VTAIL.n132 VSUBS 0.017127f
C722 VTAIL.n133 VSUBS 0.038234f
C723 VTAIL.n134 VSUBS 0.094739f
C724 VTAIL.n135 VSUBS 0.017127f
C725 VTAIL.n136 VSUBS 0.016176f
C726 VTAIL.n137 VSUBS 0.067113f
C727 VTAIL.n138 VSUBS 0.047663f
C728 VTAIL.n139 VSUBS 1.23262f
C729 VTAIL.n140 VSUBS 0.033716f
C730 VTAIL.n141 VSUBS 0.030103f
C731 VTAIL.n142 VSUBS 0.016176f
C732 VTAIL.n143 VSUBS 0.038234f
C733 VTAIL.n144 VSUBS 0.017127f
C734 VTAIL.n145 VSUBS 0.030103f
C735 VTAIL.n146 VSUBS 0.016176f
C736 VTAIL.n147 VSUBS 0.038234f
C737 VTAIL.n148 VSUBS 0.017127f
C738 VTAIL.n149 VSUBS 0.030103f
C739 VTAIL.n150 VSUBS 0.016176f
C740 VTAIL.n151 VSUBS 0.038234f
C741 VTAIL.n152 VSUBS 0.017127f
C742 VTAIL.n153 VSUBS 0.15113f
C743 VTAIL.t6 VSUBS 0.081535f
C744 VTAIL.n154 VSUBS 0.028675f
C745 VTAIL.n155 VSUBS 0.024322f
C746 VTAIL.n156 VSUBS 0.016176f
C747 VTAIL.n157 VSUBS 0.978779f
C748 VTAIL.n158 VSUBS 0.030103f
C749 VTAIL.n159 VSUBS 0.016176f
C750 VTAIL.n160 VSUBS 0.017127f
C751 VTAIL.n161 VSUBS 0.038234f
C752 VTAIL.n162 VSUBS 0.038234f
C753 VTAIL.n163 VSUBS 0.017127f
C754 VTAIL.n164 VSUBS 0.016176f
C755 VTAIL.n165 VSUBS 0.030103f
C756 VTAIL.n166 VSUBS 0.030103f
C757 VTAIL.n167 VSUBS 0.016176f
C758 VTAIL.n168 VSUBS 0.017127f
C759 VTAIL.n169 VSUBS 0.038234f
C760 VTAIL.n170 VSUBS 0.038234f
C761 VTAIL.n171 VSUBS 0.017127f
C762 VTAIL.n172 VSUBS 0.016176f
C763 VTAIL.n173 VSUBS 0.030103f
C764 VTAIL.n174 VSUBS 0.030103f
C765 VTAIL.n175 VSUBS 0.016176f
C766 VTAIL.n176 VSUBS 0.017127f
C767 VTAIL.n177 VSUBS 0.038234f
C768 VTAIL.n178 VSUBS 0.094739f
C769 VTAIL.n179 VSUBS 0.017127f
C770 VTAIL.n180 VSUBS 0.016176f
C771 VTAIL.n181 VSUBS 0.067113f
C772 VTAIL.n182 VSUBS 0.047663f
C773 VTAIL.n183 VSUBS 1.21172f
C774 VDD2.n0 VSUBS 0.028935f
C775 VDD2.n1 VSUBS 0.025834f
C776 VDD2.n2 VSUBS 0.013882f
C777 VDD2.n3 VSUBS 0.032812f
C778 VDD2.n4 VSUBS 0.014698f
C779 VDD2.n5 VSUBS 0.025834f
C780 VDD2.n6 VSUBS 0.013882f
C781 VDD2.n7 VSUBS 0.032812f
C782 VDD2.n8 VSUBS 0.014698f
C783 VDD2.n9 VSUBS 0.025834f
C784 VDD2.n10 VSUBS 0.013882f
C785 VDD2.n11 VSUBS 0.032812f
C786 VDD2.n12 VSUBS 0.014698f
C787 VDD2.n13 VSUBS 0.129698f
C788 VDD2.t5 VSUBS 0.069972f
C789 VDD2.n14 VSUBS 0.024609f
C790 VDD2.n15 VSUBS 0.020873f
C791 VDD2.n16 VSUBS 0.013882f
C792 VDD2.n17 VSUBS 0.839974f
C793 VDD2.n18 VSUBS 0.025834f
C794 VDD2.n19 VSUBS 0.013882f
C795 VDD2.n20 VSUBS 0.014698f
C796 VDD2.n21 VSUBS 0.032812f
C797 VDD2.n22 VSUBS 0.032812f
C798 VDD2.n23 VSUBS 0.014698f
C799 VDD2.n24 VSUBS 0.013882f
C800 VDD2.n25 VSUBS 0.025834f
C801 VDD2.n26 VSUBS 0.025834f
C802 VDD2.n27 VSUBS 0.013882f
C803 VDD2.n28 VSUBS 0.014698f
C804 VDD2.n29 VSUBS 0.032812f
C805 VDD2.n30 VSUBS 0.032812f
C806 VDD2.n31 VSUBS 0.014698f
C807 VDD2.n32 VSUBS 0.013882f
C808 VDD2.n33 VSUBS 0.025834f
C809 VDD2.n34 VSUBS 0.025834f
C810 VDD2.n35 VSUBS 0.013882f
C811 VDD2.n36 VSUBS 0.014698f
C812 VDD2.n37 VSUBS 0.032812f
C813 VDD2.n38 VSUBS 0.081304f
C814 VDD2.n39 VSUBS 0.014698f
C815 VDD2.n40 VSUBS 0.013882f
C816 VDD2.n41 VSUBS 0.057596f
C817 VDD2.n42 VSUBS 0.059492f
C818 VDD2.t0 VSUBS 0.165358f
C819 VDD2.t3 VSUBS 0.165358f
C820 VDD2.n43 VSUBS 1.1805f
C821 VDD2.n44 VSUBS 1.78307f
C822 VDD2.n45 VSUBS 0.028935f
C823 VDD2.n46 VSUBS 0.025834f
C824 VDD2.n47 VSUBS 0.013882f
C825 VDD2.n48 VSUBS 0.032812f
C826 VDD2.n49 VSUBS 0.014698f
C827 VDD2.n50 VSUBS 0.025834f
C828 VDD2.n51 VSUBS 0.013882f
C829 VDD2.n52 VSUBS 0.032812f
C830 VDD2.n53 VSUBS 0.014698f
C831 VDD2.n54 VSUBS 0.025834f
C832 VDD2.n55 VSUBS 0.013882f
C833 VDD2.n56 VSUBS 0.032812f
C834 VDD2.n57 VSUBS 0.014698f
C835 VDD2.n58 VSUBS 0.129698f
C836 VDD2.t1 VSUBS 0.069972f
C837 VDD2.n59 VSUBS 0.024609f
C838 VDD2.n60 VSUBS 0.020873f
C839 VDD2.n61 VSUBS 0.013882f
C840 VDD2.n62 VSUBS 0.839974f
C841 VDD2.n63 VSUBS 0.025834f
C842 VDD2.n64 VSUBS 0.013882f
C843 VDD2.n65 VSUBS 0.014698f
C844 VDD2.n66 VSUBS 0.032812f
C845 VDD2.n67 VSUBS 0.032812f
C846 VDD2.n68 VSUBS 0.014698f
C847 VDD2.n69 VSUBS 0.013882f
C848 VDD2.n70 VSUBS 0.025834f
C849 VDD2.n71 VSUBS 0.025834f
C850 VDD2.n72 VSUBS 0.013882f
C851 VDD2.n73 VSUBS 0.014698f
C852 VDD2.n74 VSUBS 0.032812f
C853 VDD2.n75 VSUBS 0.032812f
C854 VDD2.n76 VSUBS 0.014698f
C855 VDD2.n77 VSUBS 0.013882f
C856 VDD2.n78 VSUBS 0.025834f
C857 VDD2.n79 VSUBS 0.025834f
C858 VDD2.n80 VSUBS 0.013882f
C859 VDD2.n81 VSUBS 0.014698f
C860 VDD2.n82 VSUBS 0.032812f
C861 VDD2.n83 VSUBS 0.081304f
C862 VDD2.n84 VSUBS 0.014698f
C863 VDD2.n85 VSUBS 0.013882f
C864 VDD2.n86 VSUBS 0.057596f
C865 VDD2.n87 VSUBS 0.058759f
C866 VDD2.n88 VSUBS 1.70772f
C867 VDD2.t2 VSUBS 0.165358f
C868 VDD2.t4 VSUBS 0.165358f
C869 VDD2.n89 VSUBS 1.18048f
C870 VN.t5 VSUBS 0.656475f
C871 VN.n0 VSUBS 0.275531f
C872 VN.t0 VSUBS 0.645478f
C873 VN.n1 VSUBS 0.296272f
C874 VN.t3 VSUBS 0.647484f
C875 VN.n2 VSUBS 0.284014f
C876 VN.n3 VSUBS 0.207153f
C877 VN.t4 VSUBS 0.656475f
C878 VN.n4 VSUBS 0.275531f
C879 VN.t1 VSUBS 0.647484f
C880 VN.t2 VSUBS 0.645478f
C881 VN.n5 VSUBS 0.296272f
C882 VN.n6 VSUBS 0.284014f
C883 VN.n7 VSUBS 2.50828f
.ends

