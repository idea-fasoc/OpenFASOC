* NGSPICE file created from diff_pair_sample_0266.ext - technology: sky130A

.subckt diff_pair_sample_0266 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=1.29
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=1.29
X2 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=1.29
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=1.29
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=1.29
X5 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=1.29
X6 VDD1.t2 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=1.29
X7 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=1.29
X8 VDD1.t1 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=1.29
X9 VTAIL.t4 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=1.29
X10 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=1.29
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=1.29
R0 VP.n2 VP.t0 393.598
R1 VP.n2 VP.t1 393.372
R2 VP.n3 VP.t3 356.269
R3 VP.n9 VP.t2 356.269
R4 VP.n4 VP.n3 170.597
R5 VP.n10 VP.n9 170.597
R6 VP.n8 VP.n0 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n5 VP.n1 161.3
R9 VP.n4 VP.n2 65.6167
R10 VP.n7 VP.n1 40.4934
R11 VP.n8 VP.n7 40.4934
R12 VP.n3 VP.n1 15.17
R13 VP.n9 VP.n8 15.17
R14 VP.n5 VP.n4 0.189894
R15 VP.n6 VP.n5 0.189894
R16 VP.n6 VP.n0 0.189894
R17 VP.n10 VP.n0 0.189894
R18 VP VP.n10 0.0516364
R19 VDD1 VDD1.n1 107.201
R20 VDD1 VDD1.n0 62.3909
R21 VDD1.n0 VDD1.t3 1.03878
R22 VDD1.n0 VDD1.t2 1.03878
R23 VDD1.n1 VDD1.t0 1.03878
R24 VDD1.n1 VDD1.t1 1.03878
R25 VTAIL.n5 VTAIL.t7 46.6923
R26 VTAIL.n4 VTAIL.t1 46.6923
R27 VTAIL.n3 VTAIL.t2 46.6923
R28 VTAIL.n7 VTAIL.t0 46.6922
R29 VTAIL.n0 VTAIL.t3 46.6922
R30 VTAIL.n1 VTAIL.t5 46.6922
R31 VTAIL.n2 VTAIL.t4 46.6922
R32 VTAIL.n6 VTAIL.t6 46.6922
R33 VTAIL.n7 VTAIL.n6 30.2031
R34 VTAIL.n3 VTAIL.n2 30.2031
R35 VTAIL.n4 VTAIL.n3 1.39705
R36 VTAIL.n6 VTAIL.n5 1.39705
R37 VTAIL.n2 VTAIL.n1 1.39705
R38 VTAIL VTAIL.n0 0.756965
R39 VTAIL VTAIL.n7 0.640586
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 B.n598 B.n597 585
R43 B.n599 B.n116 585
R44 B.n601 B.n600 585
R45 B.n603 B.n115 585
R46 B.n606 B.n605 585
R47 B.n607 B.n114 585
R48 B.n609 B.n608 585
R49 B.n611 B.n113 585
R50 B.n614 B.n613 585
R51 B.n615 B.n112 585
R52 B.n617 B.n616 585
R53 B.n619 B.n111 585
R54 B.n622 B.n621 585
R55 B.n623 B.n110 585
R56 B.n625 B.n624 585
R57 B.n627 B.n109 585
R58 B.n630 B.n629 585
R59 B.n631 B.n108 585
R60 B.n633 B.n632 585
R61 B.n635 B.n107 585
R62 B.n638 B.n637 585
R63 B.n639 B.n106 585
R64 B.n641 B.n640 585
R65 B.n643 B.n105 585
R66 B.n646 B.n645 585
R67 B.n647 B.n104 585
R68 B.n649 B.n648 585
R69 B.n651 B.n103 585
R70 B.n654 B.n653 585
R71 B.n655 B.n102 585
R72 B.n657 B.n656 585
R73 B.n659 B.n101 585
R74 B.n662 B.n661 585
R75 B.n663 B.n100 585
R76 B.n665 B.n664 585
R77 B.n667 B.n99 585
R78 B.n670 B.n669 585
R79 B.n671 B.n98 585
R80 B.n673 B.n672 585
R81 B.n675 B.n97 585
R82 B.n678 B.n677 585
R83 B.n679 B.n96 585
R84 B.n681 B.n680 585
R85 B.n683 B.n95 585
R86 B.n686 B.n685 585
R87 B.n687 B.n94 585
R88 B.n689 B.n688 585
R89 B.n691 B.n93 585
R90 B.n694 B.n693 585
R91 B.n695 B.n92 585
R92 B.n697 B.n696 585
R93 B.n699 B.n91 585
R94 B.n702 B.n701 585
R95 B.n703 B.n90 585
R96 B.n705 B.n704 585
R97 B.n707 B.n89 585
R98 B.n710 B.n709 585
R99 B.n711 B.n88 585
R100 B.n713 B.n712 585
R101 B.n715 B.n87 585
R102 B.n717 B.n716 585
R103 B.n719 B.n718 585
R104 B.n722 B.n721 585
R105 B.n723 B.n82 585
R106 B.n725 B.n724 585
R107 B.n727 B.n81 585
R108 B.n730 B.n729 585
R109 B.n731 B.n80 585
R110 B.n733 B.n732 585
R111 B.n735 B.n79 585
R112 B.n737 B.n736 585
R113 B.n739 B.n738 585
R114 B.n742 B.n741 585
R115 B.n743 B.n74 585
R116 B.n745 B.n744 585
R117 B.n747 B.n73 585
R118 B.n750 B.n749 585
R119 B.n751 B.n72 585
R120 B.n753 B.n752 585
R121 B.n755 B.n71 585
R122 B.n758 B.n757 585
R123 B.n759 B.n70 585
R124 B.n761 B.n760 585
R125 B.n763 B.n69 585
R126 B.n766 B.n765 585
R127 B.n767 B.n68 585
R128 B.n769 B.n768 585
R129 B.n771 B.n67 585
R130 B.n774 B.n773 585
R131 B.n775 B.n66 585
R132 B.n777 B.n776 585
R133 B.n779 B.n65 585
R134 B.n782 B.n781 585
R135 B.n783 B.n64 585
R136 B.n785 B.n784 585
R137 B.n787 B.n63 585
R138 B.n790 B.n789 585
R139 B.n791 B.n62 585
R140 B.n793 B.n792 585
R141 B.n795 B.n61 585
R142 B.n798 B.n797 585
R143 B.n799 B.n60 585
R144 B.n801 B.n800 585
R145 B.n803 B.n59 585
R146 B.n806 B.n805 585
R147 B.n807 B.n58 585
R148 B.n809 B.n808 585
R149 B.n811 B.n57 585
R150 B.n814 B.n813 585
R151 B.n815 B.n56 585
R152 B.n817 B.n816 585
R153 B.n819 B.n55 585
R154 B.n822 B.n821 585
R155 B.n823 B.n54 585
R156 B.n825 B.n824 585
R157 B.n827 B.n53 585
R158 B.n830 B.n829 585
R159 B.n831 B.n52 585
R160 B.n833 B.n832 585
R161 B.n835 B.n51 585
R162 B.n838 B.n837 585
R163 B.n839 B.n50 585
R164 B.n841 B.n840 585
R165 B.n843 B.n49 585
R166 B.n846 B.n845 585
R167 B.n847 B.n48 585
R168 B.n849 B.n848 585
R169 B.n851 B.n47 585
R170 B.n854 B.n853 585
R171 B.n855 B.n46 585
R172 B.n857 B.n856 585
R173 B.n859 B.n45 585
R174 B.n862 B.n861 585
R175 B.n863 B.n44 585
R176 B.n595 B.n42 585
R177 B.n866 B.n42 585
R178 B.n594 B.n41 585
R179 B.n867 B.n41 585
R180 B.n593 B.n40 585
R181 B.n868 B.n40 585
R182 B.n592 B.n591 585
R183 B.n591 B.n36 585
R184 B.n590 B.n35 585
R185 B.n874 B.n35 585
R186 B.n589 B.n34 585
R187 B.n875 B.n34 585
R188 B.n588 B.n33 585
R189 B.n876 B.n33 585
R190 B.n587 B.n586 585
R191 B.n586 B.n29 585
R192 B.n585 B.n28 585
R193 B.n882 B.n28 585
R194 B.n584 B.n27 585
R195 B.n883 B.n27 585
R196 B.n583 B.n26 585
R197 B.n884 B.n26 585
R198 B.n582 B.n581 585
R199 B.n581 B.n22 585
R200 B.n580 B.n21 585
R201 B.n890 B.n21 585
R202 B.n579 B.n20 585
R203 B.n891 B.n20 585
R204 B.n578 B.n19 585
R205 B.n892 B.n19 585
R206 B.n577 B.n576 585
R207 B.n576 B.n15 585
R208 B.n575 B.n14 585
R209 B.n898 B.n14 585
R210 B.n574 B.n13 585
R211 B.n899 B.n13 585
R212 B.n573 B.n12 585
R213 B.n900 B.n12 585
R214 B.n572 B.n571 585
R215 B.n571 B.n570 585
R216 B.n569 B.n568 585
R217 B.n569 B.n8 585
R218 B.n567 B.n7 585
R219 B.n907 B.n7 585
R220 B.n566 B.n6 585
R221 B.n908 B.n6 585
R222 B.n565 B.n5 585
R223 B.n909 B.n5 585
R224 B.n564 B.n563 585
R225 B.n563 B.n4 585
R226 B.n562 B.n117 585
R227 B.n562 B.n561 585
R228 B.n552 B.n118 585
R229 B.n119 B.n118 585
R230 B.n554 B.n553 585
R231 B.n555 B.n554 585
R232 B.n551 B.n124 585
R233 B.n124 B.n123 585
R234 B.n550 B.n549 585
R235 B.n549 B.n548 585
R236 B.n126 B.n125 585
R237 B.n127 B.n126 585
R238 B.n541 B.n540 585
R239 B.n542 B.n541 585
R240 B.n539 B.n131 585
R241 B.n135 B.n131 585
R242 B.n538 B.n537 585
R243 B.n537 B.n536 585
R244 B.n133 B.n132 585
R245 B.n134 B.n133 585
R246 B.n529 B.n528 585
R247 B.n530 B.n529 585
R248 B.n527 B.n140 585
R249 B.n140 B.n139 585
R250 B.n526 B.n525 585
R251 B.n525 B.n524 585
R252 B.n142 B.n141 585
R253 B.n143 B.n142 585
R254 B.n517 B.n516 585
R255 B.n518 B.n517 585
R256 B.n515 B.n147 585
R257 B.n151 B.n147 585
R258 B.n514 B.n513 585
R259 B.n513 B.n512 585
R260 B.n149 B.n148 585
R261 B.n150 B.n149 585
R262 B.n505 B.n504 585
R263 B.n506 B.n505 585
R264 B.n503 B.n156 585
R265 B.n156 B.n155 585
R266 B.n502 B.n501 585
R267 B.n501 B.n500 585
R268 B.n497 B.n160 585
R269 B.n496 B.n495 585
R270 B.n493 B.n161 585
R271 B.n493 B.n159 585
R272 B.n492 B.n491 585
R273 B.n490 B.n489 585
R274 B.n488 B.n163 585
R275 B.n486 B.n485 585
R276 B.n484 B.n164 585
R277 B.n483 B.n482 585
R278 B.n480 B.n165 585
R279 B.n478 B.n477 585
R280 B.n476 B.n166 585
R281 B.n475 B.n474 585
R282 B.n472 B.n167 585
R283 B.n470 B.n469 585
R284 B.n468 B.n168 585
R285 B.n467 B.n466 585
R286 B.n464 B.n169 585
R287 B.n462 B.n461 585
R288 B.n460 B.n170 585
R289 B.n459 B.n458 585
R290 B.n456 B.n171 585
R291 B.n454 B.n453 585
R292 B.n452 B.n172 585
R293 B.n451 B.n450 585
R294 B.n448 B.n173 585
R295 B.n446 B.n445 585
R296 B.n444 B.n174 585
R297 B.n443 B.n442 585
R298 B.n440 B.n175 585
R299 B.n438 B.n437 585
R300 B.n436 B.n176 585
R301 B.n435 B.n434 585
R302 B.n432 B.n177 585
R303 B.n430 B.n429 585
R304 B.n428 B.n178 585
R305 B.n427 B.n426 585
R306 B.n424 B.n179 585
R307 B.n422 B.n421 585
R308 B.n420 B.n180 585
R309 B.n419 B.n418 585
R310 B.n416 B.n181 585
R311 B.n414 B.n413 585
R312 B.n412 B.n182 585
R313 B.n411 B.n410 585
R314 B.n408 B.n183 585
R315 B.n406 B.n405 585
R316 B.n404 B.n184 585
R317 B.n403 B.n402 585
R318 B.n400 B.n185 585
R319 B.n398 B.n397 585
R320 B.n396 B.n186 585
R321 B.n395 B.n394 585
R322 B.n392 B.n187 585
R323 B.n390 B.n389 585
R324 B.n388 B.n188 585
R325 B.n387 B.n386 585
R326 B.n384 B.n189 585
R327 B.n382 B.n381 585
R328 B.n380 B.n190 585
R329 B.n379 B.n378 585
R330 B.n376 B.n191 585
R331 B.n374 B.n373 585
R332 B.n372 B.n192 585
R333 B.n371 B.n370 585
R334 B.n368 B.n196 585
R335 B.n366 B.n365 585
R336 B.n364 B.n197 585
R337 B.n363 B.n362 585
R338 B.n360 B.n198 585
R339 B.n358 B.n357 585
R340 B.n356 B.n199 585
R341 B.n354 B.n353 585
R342 B.n351 B.n202 585
R343 B.n349 B.n348 585
R344 B.n347 B.n203 585
R345 B.n346 B.n345 585
R346 B.n343 B.n204 585
R347 B.n341 B.n340 585
R348 B.n339 B.n205 585
R349 B.n338 B.n337 585
R350 B.n335 B.n206 585
R351 B.n333 B.n332 585
R352 B.n331 B.n207 585
R353 B.n330 B.n329 585
R354 B.n327 B.n208 585
R355 B.n325 B.n324 585
R356 B.n323 B.n209 585
R357 B.n322 B.n321 585
R358 B.n319 B.n210 585
R359 B.n317 B.n316 585
R360 B.n315 B.n211 585
R361 B.n314 B.n313 585
R362 B.n311 B.n212 585
R363 B.n309 B.n308 585
R364 B.n307 B.n213 585
R365 B.n306 B.n305 585
R366 B.n303 B.n214 585
R367 B.n301 B.n300 585
R368 B.n299 B.n215 585
R369 B.n298 B.n297 585
R370 B.n295 B.n216 585
R371 B.n293 B.n292 585
R372 B.n291 B.n217 585
R373 B.n290 B.n289 585
R374 B.n287 B.n218 585
R375 B.n285 B.n284 585
R376 B.n283 B.n219 585
R377 B.n282 B.n281 585
R378 B.n279 B.n220 585
R379 B.n277 B.n276 585
R380 B.n275 B.n221 585
R381 B.n274 B.n273 585
R382 B.n271 B.n222 585
R383 B.n269 B.n268 585
R384 B.n267 B.n223 585
R385 B.n266 B.n265 585
R386 B.n263 B.n224 585
R387 B.n261 B.n260 585
R388 B.n259 B.n225 585
R389 B.n258 B.n257 585
R390 B.n255 B.n226 585
R391 B.n253 B.n252 585
R392 B.n251 B.n227 585
R393 B.n250 B.n249 585
R394 B.n247 B.n228 585
R395 B.n245 B.n244 585
R396 B.n243 B.n229 585
R397 B.n242 B.n241 585
R398 B.n239 B.n230 585
R399 B.n237 B.n236 585
R400 B.n235 B.n231 585
R401 B.n234 B.n233 585
R402 B.n158 B.n157 585
R403 B.n159 B.n158 585
R404 B.n499 B.n498 585
R405 B.n500 B.n499 585
R406 B.n154 B.n153 585
R407 B.n155 B.n154 585
R408 B.n508 B.n507 585
R409 B.n507 B.n506 585
R410 B.n509 B.n152 585
R411 B.n152 B.n150 585
R412 B.n511 B.n510 585
R413 B.n512 B.n511 585
R414 B.n146 B.n145 585
R415 B.n151 B.n146 585
R416 B.n520 B.n519 585
R417 B.n519 B.n518 585
R418 B.n521 B.n144 585
R419 B.n144 B.n143 585
R420 B.n523 B.n522 585
R421 B.n524 B.n523 585
R422 B.n138 B.n137 585
R423 B.n139 B.n138 585
R424 B.n532 B.n531 585
R425 B.n531 B.n530 585
R426 B.n533 B.n136 585
R427 B.n136 B.n134 585
R428 B.n535 B.n534 585
R429 B.n536 B.n535 585
R430 B.n130 B.n129 585
R431 B.n135 B.n130 585
R432 B.n544 B.n543 585
R433 B.n543 B.n542 585
R434 B.n545 B.n128 585
R435 B.n128 B.n127 585
R436 B.n547 B.n546 585
R437 B.n548 B.n547 585
R438 B.n122 B.n121 585
R439 B.n123 B.n122 585
R440 B.n557 B.n556 585
R441 B.n556 B.n555 585
R442 B.n558 B.n120 585
R443 B.n120 B.n119 585
R444 B.n560 B.n559 585
R445 B.n561 B.n560 585
R446 B.n3 B.n0 585
R447 B.n4 B.n3 585
R448 B.n906 B.n1 585
R449 B.n907 B.n906 585
R450 B.n905 B.n904 585
R451 B.n905 B.n8 585
R452 B.n903 B.n9 585
R453 B.n570 B.n9 585
R454 B.n902 B.n901 585
R455 B.n901 B.n900 585
R456 B.n11 B.n10 585
R457 B.n899 B.n11 585
R458 B.n897 B.n896 585
R459 B.n898 B.n897 585
R460 B.n895 B.n16 585
R461 B.n16 B.n15 585
R462 B.n894 B.n893 585
R463 B.n893 B.n892 585
R464 B.n18 B.n17 585
R465 B.n891 B.n18 585
R466 B.n889 B.n888 585
R467 B.n890 B.n889 585
R468 B.n887 B.n23 585
R469 B.n23 B.n22 585
R470 B.n886 B.n885 585
R471 B.n885 B.n884 585
R472 B.n25 B.n24 585
R473 B.n883 B.n25 585
R474 B.n881 B.n880 585
R475 B.n882 B.n881 585
R476 B.n879 B.n30 585
R477 B.n30 B.n29 585
R478 B.n878 B.n877 585
R479 B.n877 B.n876 585
R480 B.n32 B.n31 585
R481 B.n875 B.n32 585
R482 B.n873 B.n872 585
R483 B.n874 B.n873 585
R484 B.n871 B.n37 585
R485 B.n37 B.n36 585
R486 B.n870 B.n869 585
R487 B.n869 B.n868 585
R488 B.n39 B.n38 585
R489 B.n867 B.n39 585
R490 B.n865 B.n864 585
R491 B.n866 B.n865 585
R492 B.n910 B.n909 585
R493 B.n908 B.n2 585
R494 B.n75 B.t8 560.832
R495 B.n83 B.t12 560.832
R496 B.n200 B.t4 560.832
R497 B.n193 B.t15 560.832
R498 B.n865 B.n44 516.524
R499 B.n597 B.n42 516.524
R500 B.n501 B.n158 516.524
R501 B.n499 B.n160 516.524
R502 B.n596 B.n43 256.663
R503 B.n602 B.n43 256.663
R504 B.n604 B.n43 256.663
R505 B.n610 B.n43 256.663
R506 B.n612 B.n43 256.663
R507 B.n618 B.n43 256.663
R508 B.n620 B.n43 256.663
R509 B.n626 B.n43 256.663
R510 B.n628 B.n43 256.663
R511 B.n634 B.n43 256.663
R512 B.n636 B.n43 256.663
R513 B.n642 B.n43 256.663
R514 B.n644 B.n43 256.663
R515 B.n650 B.n43 256.663
R516 B.n652 B.n43 256.663
R517 B.n658 B.n43 256.663
R518 B.n660 B.n43 256.663
R519 B.n666 B.n43 256.663
R520 B.n668 B.n43 256.663
R521 B.n674 B.n43 256.663
R522 B.n676 B.n43 256.663
R523 B.n682 B.n43 256.663
R524 B.n684 B.n43 256.663
R525 B.n690 B.n43 256.663
R526 B.n692 B.n43 256.663
R527 B.n698 B.n43 256.663
R528 B.n700 B.n43 256.663
R529 B.n706 B.n43 256.663
R530 B.n708 B.n43 256.663
R531 B.n714 B.n43 256.663
R532 B.n86 B.n43 256.663
R533 B.n720 B.n43 256.663
R534 B.n726 B.n43 256.663
R535 B.n728 B.n43 256.663
R536 B.n734 B.n43 256.663
R537 B.n78 B.n43 256.663
R538 B.n740 B.n43 256.663
R539 B.n746 B.n43 256.663
R540 B.n748 B.n43 256.663
R541 B.n754 B.n43 256.663
R542 B.n756 B.n43 256.663
R543 B.n762 B.n43 256.663
R544 B.n764 B.n43 256.663
R545 B.n770 B.n43 256.663
R546 B.n772 B.n43 256.663
R547 B.n778 B.n43 256.663
R548 B.n780 B.n43 256.663
R549 B.n786 B.n43 256.663
R550 B.n788 B.n43 256.663
R551 B.n794 B.n43 256.663
R552 B.n796 B.n43 256.663
R553 B.n802 B.n43 256.663
R554 B.n804 B.n43 256.663
R555 B.n810 B.n43 256.663
R556 B.n812 B.n43 256.663
R557 B.n818 B.n43 256.663
R558 B.n820 B.n43 256.663
R559 B.n826 B.n43 256.663
R560 B.n828 B.n43 256.663
R561 B.n834 B.n43 256.663
R562 B.n836 B.n43 256.663
R563 B.n842 B.n43 256.663
R564 B.n844 B.n43 256.663
R565 B.n850 B.n43 256.663
R566 B.n852 B.n43 256.663
R567 B.n858 B.n43 256.663
R568 B.n860 B.n43 256.663
R569 B.n494 B.n159 256.663
R570 B.n162 B.n159 256.663
R571 B.n487 B.n159 256.663
R572 B.n481 B.n159 256.663
R573 B.n479 B.n159 256.663
R574 B.n473 B.n159 256.663
R575 B.n471 B.n159 256.663
R576 B.n465 B.n159 256.663
R577 B.n463 B.n159 256.663
R578 B.n457 B.n159 256.663
R579 B.n455 B.n159 256.663
R580 B.n449 B.n159 256.663
R581 B.n447 B.n159 256.663
R582 B.n441 B.n159 256.663
R583 B.n439 B.n159 256.663
R584 B.n433 B.n159 256.663
R585 B.n431 B.n159 256.663
R586 B.n425 B.n159 256.663
R587 B.n423 B.n159 256.663
R588 B.n417 B.n159 256.663
R589 B.n415 B.n159 256.663
R590 B.n409 B.n159 256.663
R591 B.n407 B.n159 256.663
R592 B.n401 B.n159 256.663
R593 B.n399 B.n159 256.663
R594 B.n393 B.n159 256.663
R595 B.n391 B.n159 256.663
R596 B.n385 B.n159 256.663
R597 B.n383 B.n159 256.663
R598 B.n377 B.n159 256.663
R599 B.n375 B.n159 256.663
R600 B.n369 B.n159 256.663
R601 B.n367 B.n159 256.663
R602 B.n361 B.n159 256.663
R603 B.n359 B.n159 256.663
R604 B.n352 B.n159 256.663
R605 B.n350 B.n159 256.663
R606 B.n344 B.n159 256.663
R607 B.n342 B.n159 256.663
R608 B.n336 B.n159 256.663
R609 B.n334 B.n159 256.663
R610 B.n328 B.n159 256.663
R611 B.n326 B.n159 256.663
R612 B.n320 B.n159 256.663
R613 B.n318 B.n159 256.663
R614 B.n312 B.n159 256.663
R615 B.n310 B.n159 256.663
R616 B.n304 B.n159 256.663
R617 B.n302 B.n159 256.663
R618 B.n296 B.n159 256.663
R619 B.n294 B.n159 256.663
R620 B.n288 B.n159 256.663
R621 B.n286 B.n159 256.663
R622 B.n280 B.n159 256.663
R623 B.n278 B.n159 256.663
R624 B.n272 B.n159 256.663
R625 B.n270 B.n159 256.663
R626 B.n264 B.n159 256.663
R627 B.n262 B.n159 256.663
R628 B.n256 B.n159 256.663
R629 B.n254 B.n159 256.663
R630 B.n248 B.n159 256.663
R631 B.n246 B.n159 256.663
R632 B.n240 B.n159 256.663
R633 B.n238 B.n159 256.663
R634 B.n232 B.n159 256.663
R635 B.n912 B.n911 256.663
R636 B.n861 B.n859 163.367
R637 B.n857 B.n46 163.367
R638 B.n853 B.n851 163.367
R639 B.n849 B.n48 163.367
R640 B.n845 B.n843 163.367
R641 B.n841 B.n50 163.367
R642 B.n837 B.n835 163.367
R643 B.n833 B.n52 163.367
R644 B.n829 B.n827 163.367
R645 B.n825 B.n54 163.367
R646 B.n821 B.n819 163.367
R647 B.n817 B.n56 163.367
R648 B.n813 B.n811 163.367
R649 B.n809 B.n58 163.367
R650 B.n805 B.n803 163.367
R651 B.n801 B.n60 163.367
R652 B.n797 B.n795 163.367
R653 B.n793 B.n62 163.367
R654 B.n789 B.n787 163.367
R655 B.n785 B.n64 163.367
R656 B.n781 B.n779 163.367
R657 B.n777 B.n66 163.367
R658 B.n773 B.n771 163.367
R659 B.n769 B.n68 163.367
R660 B.n765 B.n763 163.367
R661 B.n761 B.n70 163.367
R662 B.n757 B.n755 163.367
R663 B.n753 B.n72 163.367
R664 B.n749 B.n747 163.367
R665 B.n745 B.n74 163.367
R666 B.n741 B.n739 163.367
R667 B.n736 B.n735 163.367
R668 B.n733 B.n80 163.367
R669 B.n729 B.n727 163.367
R670 B.n725 B.n82 163.367
R671 B.n721 B.n719 163.367
R672 B.n716 B.n715 163.367
R673 B.n713 B.n88 163.367
R674 B.n709 B.n707 163.367
R675 B.n705 B.n90 163.367
R676 B.n701 B.n699 163.367
R677 B.n697 B.n92 163.367
R678 B.n693 B.n691 163.367
R679 B.n689 B.n94 163.367
R680 B.n685 B.n683 163.367
R681 B.n681 B.n96 163.367
R682 B.n677 B.n675 163.367
R683 B.n673 B.n98 163.367
R684 B.n669 B.n667 163.367
R685 B.n665 B.n100 163.367
R686 B.n661 B.n659 163.367
R687 B.n657 B.n102 163.367
R688 B.n653 B.n651 163.367
R689 B.n649 B.n104 163.367
R690 B.n645 B.n643 163.367
R691 B.n641 B.n106 163.367
R692 B.n637 B.n635 163.367
R693 B.n633 B.n108 163.367
R694 B.n629 B.n627 163.367
R695 B.n625 B.n110 163.367
R696 B.n621 B.n619 163.367
R697 B.n617 B.n112 163.367
R698 B.n613 B.n611 163.367
R699 B.n609 B.n114 163.367
R700 B.n605 B.n603 163.367
R701 B.n601 B.n116 163.367
R702 B.n501 B.n156 163.367
R703 B.n505 B.n156 163.367
R704 B.n505 B.n149 163.367
R705 B.n513 B.n149 163.367
R706 B.n513 B.n147 163.367
R707 B.n517 B.n147 163.367
R708 B.n517 B.n142 163.367
R709 B.n525 B.n142 163.367
R710 B.n525 B.n140 163.367
R711 B.n529 B.n140 163.367
R712 B.n529 B.n133 163.367
R713 B.n537 B.n133 163.367
R714 B.n537 B.n131 163.367
R715 B.n541 B.n131 163.367
R716 B.n541 B.n126 163.367
R717 B.n549 B.n126 163.367
R718 B.n549 B.n124 163.367
R719 B.n554 B.n124 163.367
R720 B.n554 B.n118 163.367
R721 B.n562 B.n118 163.367
R722 B.n563 B.n562 163.367
R723 B.n563 B.n5 163.367
R724 B.n6 B.n5 163.367
R725 B.n7 B.n6 163.367
R726 B.n569 B.n7 163.367
R727 B.n571 B.n569 163.367
R728 B.n571 B.n12 163.367
R729 B.n13 B.n12 163.367
R730 B.n14 B.n13 163.367
R731 B.n576 B.n14 163.367
R732 B.n576 B.n19 163.367
R733 B.n20 B.n19 163.367
R734 B.n21 B.n20 163.367
R735 B.n581 B.n21 163.367
R736 B.n581 B.n26 163.367
R737 B.n27 B.n26 163.367
R738 B.n28 B.n27 163.367
R739 B.n586 B.n28 163.367
R740 B.n586 B.n33 163.367
R741 B.n34 B.n33 163.367
R742 B.n35 B.n34 163.367
R743 B.n591 B.n35 163.367
R744 B.n591 B.n40 163.367
R745 B.n41 B.n40 163.367
R746 B.n42 B.n41 163.367
R747 B.n495 B.n493 163.367
R748 B.n493 B.n492 163.367
R749 B.n489 B.n488 163.367
R750 B.n486 B.n164 163.367
R751 B.n482 B.n480 163.367
R752 B.n478 B.n166 163.367
R753 B.n474 B.n472 163.367
R754 B.n470 B.n168 163.367
R755 B.n466 B.n464 163.367
R756 B.n462 B.n170 163.367
R757 B.n458 B.n456 163.367
R758 B.n454 B.n172 163.367
R759 B.n450 B.n448 163.367
R760 B.n446 B.n174 163.367
R761 B.n442 B.n440 163.367
R762 B.n438 B.n176 163.367
R763 B.n434 B.n432 163.367
R764 B.n430 B.n178 163.367
R765 B.n426 B.n424 163.367
R766 B.n422 B.n180 163.367
R767 B.n418 B.n416 163.367
R768 B.n414 B.n182 163.367
R769 B.n410 B.n408 163.367
R770 B.n406 B.n184 163.367
R771 B.n402 B.n400 163.367
R772 B.n398 B.n186 163.367
R773 B.n394 B.n392 163.367
R774 B.n390 B.n188 163.367
R775 B.n386 B.n384 163.367
R776 B.n382 B.n190 163.367
R777 B.n378 B.n376 163.367
R778 B.n374 B.n192 163.367
R779 B.n370 B.n368 163.367
R780 B.n366 B.n197 163.367
R781 B.n362 B.n360 163.367
R782 B.n358 B.n199 163.367
R783 B.n353 B.n351 163.367
R784 B.n349 B.n203 163.367
R785 B.n345 B.n343 163.367
R786 B.n341 B.n205 163.367
R787 B.n337 B.n335 163.367
R788 B.n333 B.n207 163.367
R789 B.n329 B.n327 163.367
R790 B.n325 B.n209 163.367
R791 B.n321 B.n319 163.367
R792 B.n317 B.n211 163.367
R793 B.n313 B.n311 163.367
R794 B.n309 B.n213 163.367
R795 B.n305 B.n303 163.367
R796 B.n301 B.n215 163.367
R797 B.n297 B.n295 163.367
R798 B.n293 B.n217 163.367
R799 B.n289 B.n287 163.367
R800 B.n285 B.n219 163.367
R801 B.n281 B.n279 163.367
R802 B.n277 B.n221 163.367
R803 B.n273 B.n271 163.367
R804 B.n269 B.n223 163.367
R805 B.n265 B.n263 163.367
R806 B.n261 B.n225 163.367
R807 B.n257 B.n255 163.367
R808 B.n253 B.n227 163.367
R809 B.n249 B.n247 163.367
R810 B.n245 B.n229 163.367
R811 B.n241 B.n239 163.367
R812 B.n237 B.n231 163.367
R813 B.n233 B.n158 163.367
R814 B.n499 B.n154 163.367
R815 B.n507 B.n154 163.367
R816 B.n507 B.n152 163.367
R817 B.n511 B.n152 163.367
R818 B.n511 B.n146 163.367
R819 B.n519 B.n146 163.367
R820 B.n519 B.n144 163.367
R821 B.n523 B.n144 163.367
R822 B.n523 B.n138 163.367
R823 B.n531 B.n138 163.367
R824 B.n531 B.n136 163.367
R825 B.n535 B.n136 163.367
R826 B.n535 B.n130 163.367
R827 B.n543 B.n130 163.367
R828 B.n543 B.n128 163.367
R829 B.n547 B.n128 163.367
R830 B.n547 B.n122 163.367
R831 B.n556 B.n122 163.367
R832 B.n556 B.n120 163.367
R833 B.n560 B.n120 163.367
R834 B.n560 B.n3 163.367
R835 B.n910 B.n3 163.367
R836 B.n906 B.n2 163.367
R837 B.n906 B.n905 163.367
R838 B.n905 B.n9 163.367
R839 B.n901 B.n9 163.367
R840 B.n901 B.n11 163.367
R841 B.n897 B.n11 163.367
R842 B.n897 B.n16 163.367
R843 B.n893 B.n16 163.367
R844 B.n893 B.n18 163.367
R845 B.n889 B.n18 163.367
R846 B.n889 B.n23 163.367
R847 B.n885 B.n23 163.367
R848 B.n885 B.n25 163.367
R849 B.n881 B.n25 163.367
R850 B.n881 B.n30 163.367
R851 B.n877 B.n30 163.367
R852 B.n877 B.n32 163.367
R853 B.n873 B.n32 163.367
R854 B.n873 B.n37 163.367
R855 B.n869 B.n37 163.367
R856 B.n869 B.n39 163.367
R857 B.n865 B.n39 163.367
R858 B.n83 B.t13 99.1887
R859 B.n200 B.t7 99.1887
R860 B.n75 B.t10 99.1629
R861 B.n193 B.t17 99.1629
R862 B.n860 B.n44 71.676
R863 B.n859 B.n858 71.676
R864 B.n852 B.n46 71.676
R865 B.n851 B.n850 71.676
R866 B.n844 B.n48 71.676
R867 B.n843 B.n842 71.676
R868 B.n836 B.n50 71.676
R869 B.n835 B.n834 71.676
R870 B.n828 B.n52 71.676
R871 B.n827 B.n826 71.676
R872 B.n820 B.n54 71.676
R873 B.n819 B.n818 71.676
R874 B.n812 B.n56 71.676
R875 B.n811 B.n810 71.676
R876 B.n804 B.n58 71.676
R877 B.n803 B.n802 71.676
R878 B.n796 B.n60 71.676
R879 B.n795 B.n794 71.676
R880 B.n788 B.n62 71.676
R881 B.n787 B.n786 71.676
R882 B.n780 B.n64 71.676
R883 B.n779 B.n778 71.676
R884 B.n772 B.n66 71.676
R885 B.n771 B.n770 71.676
R886 B.n764 B.n68 71.676
R887 B.n763 B.n762 71.676
R888 B.n756 B.n70 71.676
R889 B.n755 B.n754 71.676
R890 B.n748 B.n72 71.676
R891 B.n747 B.n746 71.676
R892 B.n740 B.n74 71.676
R893 B.n739 B.n78 71.676
R894 B.n735 B.n734 71.676
R895 B.n728 B.n80 71.676
R896 B.n727 B.n726 71.676
R897 B.n720 B.n82 71.676
R898 B.n719 B.n86 71.676
R899 B.n715 B.n714 71.676
R900 B.n708 B.n88 71.676
R901 B.n707 B.n706 71.676
R902 B.n700 B.n90 71.676
R903 B.n699 B.n698 71.676
R904 B.n692 B.n92 71.676
R905 B.n691 B.n690 71.676
R906 B.n684 B.n94 71.676
R907 B.n683 B.n682 71.676
R908 B.n676 B.n96 71.676
R909 B.n675 B.n674 71.676
R910 B.n668 B.n98 71.676
R911 B.n667 B.n666 71.676
R912 B.n660 B.n100 71.676
R913 B.n659 B.n658 71.676
R914 B.n652 B.n102 71.676
R915 B.n651 B.n650 71.676
R916 B.n644 B.n104 71.676
R917 B.n643 B.n642 71.676
R918 B.n636 B.n106 71.676
R919 B.n635 B.n634 71.676
R920 B.n628 B.n108 71.676
R921 B.n627 B.n626 71.676
R922 B.n620 B.n110 71.676
R923 B.n619 B.n618 71.676
R924 B.n612 B.n112 71.676
R925 B.n611 B.n610 71.676
R926 B.n604 B.n114 71.676
R927 B.n603 B.n602 71.676
R928 B.n596 B.n116 71.676
R929 B.n597 B.n596 71.676
R930 B.n602 B.n601 71.676
R931 B.n605 B.n604 71.676
R932 B.n610 B.n609 71.676
R933 B.n613 B.n612 71.676
R934 B.n618 B.n617 71.676
R935 B.n621 B.n620 71.676
R936 B.n626 B.n625 71.676
R937 B.n629 B.n628 71.676
R938 B.n634 B.n633 71.676
R939 B.n637 B.n636 71.676
R940 B.n642 B.n641 71.676
R941 B.n645 B.n644 71.676
R942 B.n650 B.n649 71.676
R943 B.n653 B.n652 71.676
R944 B.n658 B.n657 71.676
R945 B.n661 B.n660 71.676
R946 B.n666 B.n665 71.676
R947 B.n669 B.n668 71.676
R948 B.n674 B.n673 71.676
R949 B.n677 B.n676 71.676
R950 B.n682 B.n681 71.676
R951 B.n685 B.n684 71.676
R952 B.n690 B.n689 71.676
R953 B.n693 B.n692 71.676
R954 B.n698 B.n697 71.676
R955 B.n701 B.n700 71.676
R956 B.n706 B.n705 71.676
R957 B.n709 B.n708 71.676
R958 B.n714 B.n713 71.676
R959 B.n716 B.n86 71.676
R960 B.n721 B.n720 71.676
R961 B.n726 B.n725 71.676
R962 B.n729 B.n728 71.676
R963 B.n734 B.n733 71.676
R964 B.n736 B.n78 71.676
R965 B.n741 B.n740 71.676
R966 B.n746 B.n745 71.676
R967 B.n749 B.n748 71.676
R968 B.n754 B.n753 71.676
R969 B.n757 B.n756 71.676
R970 B.n762 B.n761 71.676
R971 B.n765 B.n764 71.676
R972 B.n770 B.n769 71.676
R973 B.n773 B.n772 71.676
R974 B.n778 B.n777 71.676
R975 B.n781 B.n780 71.676
R976 B.n786 B.n785 71.676
R977 B.n789 B.n788 71.676
R978 B.n794 B.n793 71.676
R979 B.n797 B.n796 71.676
R980 B.n802 B.n801 71.676
R981 B.n805 B.n804 71.676
R982 B.n810 B.n809 71.676
R983 B.n813 B.n812 71.676
R984 B.n818 B.n817 71.676
R985 B.n821 B.n820 71.676
R986 B.n826 B.n825 71.676
R987 B.n829 B.n828 71.676
R988 B.n834 B.n833 71.676
R989 B.n837 B.n836 71.676
R990 B.n842 B.n841 71.676
R991 B.n845 B.n844 71.676
R992 B.n850 B.n849 71.676
R993 B.n853 B.n852 71.676
R994 B.n858 B.n857 71.676
R995 B.n861 B.n860 71.676
R996 B.n494 B.n160 71.676
R997 B.n492 B.n162 71.676
R998 B.n488 B.n487 71.676
R999 B.n481 B.n164 71.676
R1000 B.n480 B.n479 71.676
R1001 B.n473 B.n166 71.676
R1002 B.n472 B.n471 71.676
R1003 B.n465 B.n168 71.676
R1004 B.n464 B.n463 71.676
R1005 B.n457 B.n170 71.676
R1006 B.n456 B.n455 71.676
R1007 B.n449 B.n172 71.676
R1008 B.n448 B.n447 71.676
R1009 B.n441 B.n174 71.676
R1010 B.n440 B.n439 71.676
R1011 B.n433 B.n176 71.676
R1012 B.n432 B.n431 71.676
R1013 B.n425 B.n178 71.676
R1014 B.n424 B.n423 71.676
R1015 B.n417 B.n180 71.676
R1016 B.n416 B.n415 71.676
R1017 B.n409 B.n182 71.676
R1018 B.n408 B.n407 71.676
R1019 B.n401 B.n184 71.676
R1020 B.n400 B.n399 71.676
R1021 B.n393 B.n186 71.676
R1022 B.n392 B.n391 71.676
R1023 B.n385 B.n188 71.676
R1024 B.n384 B.n383 71.676
R1025 B.n377 B.n190 71.676
R1026 B.n376 B.n375 71.676
R1027 B.n369 B.n192 71.676
R1028 B.n368 B.n367 71.676
R1029 B.n361 B.n197 71.676
R1030 B.n360 B.n359 71.676
R1031 B.n352 B.n199 71.676
R1032 B.n351 B.n350 71.676
R1033 B.n344 B.n203 71.676
R1034 B.n343 B.n342 71.676
R1035 B.n336 B.n205 71.676
R1036 B.n335 B.n334 71.676
R1037 B.n328 B.n207 71.676
R1038 B.n327 B.n326 71.676
R1039 B.n320 B.n209 71.676
R1040 B.n319 B.n318 71.676
R1041 B.n312 B.n211 71.676
R1042 B.n311 B.n310 71.676
R1043 B.n304 B.n213 71.676
R1044 B.n303 B.n302 71.676
R1045 B.n296 B.n215 71.676
R1046 B.n295 B.n294 71.676
R1047 B.n288 B.n217 71.676
R1048 B.n287 B.n286 71.676
R1049 B.n280 B.n219 71.676
R1050 B.n279 B.n278 71.676
R1051 B.n272 B.n221 71.676
R1052 B.n271 B.n270 71.676
R1053 B.n264 B.n223 71.676
R1054 B.n263 B.n262 71.676
R1055 B.n256 B.n225 71.676
R1056 B.n255 B.n254 71.676
R1057 B.n248 B.n227 71.676
R1058 B.n247 B.n246 71.676
R1059 B.n240 B.n229 71.676
R1060 B.n239 B.n238 71.676
R1061 B.n232 B.n231 71.676
R1062 B.n495 B.n494 71.676
R1063 B.n489 B.n162 71.676
R1064 B.n487 B.n486 71.676
R1065 B.n482 B.n481 71.676
R1066 B.n479 B.n478 71.676
R1067 B.n474 B.n473 71.676
R1068 B.n471 B.n470 71.676
R1069 B.n466 B.n465 71.676
R1070 B.n463 B.n462 71.676
R1071 B.n458 B.n457 71.676
R1072 B.n455 B.n454 71.676
R1073 B.n450 B.n449 71.676
R1074 B.n447 B.n446 71.676
R1075 B.n442 B.n441 71.676
R1076 B.n439 B.n438 71.676
R1077 B.n434 B.n433 71.676
R1078 B.n431 B.n430 71.676
R1079 B.n426 B.n425 71.676
R1080 B.n423 B.n422 71.676
R1081 B.n418 B.n417 71.676
R1082 B.n415 B.n414 71.676
R1083 B.n410 B.n409 71.676
R1084 B.n407 B.n406 71.676
R1085 B.n402 B.n401 71.676
R1086 B.n399 B.n398 71.676
R1087 B.n394 B.n393 71.676
R1088 B.n391 B.n390 71.676
R1089 B.n386 B.n385 71.676
R1090 B.n383 B.n382 71.676
R1091 B.n378 B.n377 71.676
R1092 B.n375 B.n374 71.676
R1093 B.n370 B.n369 71.676
R1094 B.n367 B.n366 71.676
R1095 B.n362 B.n361 71.676
R1096 B.n359 B.n358 71.676
R1097 B.n353 B.n352 71.676
R1098 B.n350 B.n349 71.676
R1099 B.n345 B.n344 71.676
R1100 B.n342 B.n341 71.676
R1101 B.n337 B.n336 71.676
R1102 B.n334 B.n333 71.676
R1103 B.n329 B.n328 71.676
R1104 B.n326 B.n325 71.676
R1105 B.n321 B.n320 71.676
R1106 B.n318 B.n317 71.676
R1107 B.n313 B.n312 71.676
R1108 B.n310 B.n309 71.676
R1109 B.n305 B.n304 71.676
R1110 B.n302 B.n301 71.676
R1111 B.n297 B.n296 71.676
R1112 B.n294 B.n293 71.676
R1113 B.n289 B.n288 71.676
R1114 B.n286 B.n285 71.676
R1115 B.n281 B.n280 71.676
R1116 B.n278 B.n277 71.676
R1117 B.n273 B.n272 71.676
R1118 B.n270 B.n269 71.676
R1119 B.n265 B.n264 71.676
R1120 B.n262 B.n261 71.676
R1121 B.n257 B.n256 71.676
R1122 B.n254 B.n253 71.676
R1123 B.n249 B.n248 71.676
R1124 B.n246 B.n245 71.676
R1125 B.n241 B.n240 71.676
R1126 B.n238 B.n237 71.676
R1127 B.n233 B.n232 71.676
R1128 B.n911 B.n910 71.676
R1129 B.n911 B.n2 71.676
R1130 B.n84 B.t14 67.7705
R1131 B.n201 B.t6 67.7705
R1132 B.n76 B.t11 67.7448
R1133 B.n194 B.t16 67.7448
R1134 B.n77 B.n76 59.5399
R1135 B.n85 B.n84 59.5399
R1136 B.n355 B.n201 59.5399
R1137 B.n195 B.n194 59.5399
R1138 B.n500 B.n159 52.8656
R1139 B.n866 B.n43 52.8656
R1140 B.n498 B.n497 33.5615
R1141 B.n502 B.n157 33.5615
R1142 B.n598 B.n595 33.5615
R1143 B.n864 B.n863 33.5615
R1144 B.n76 B.n75 31.4187
R1145 B.n84 B.n83 31.4187
R1146 B.n201 B.n200 31.4187
R1147 B.n194 B.n193 31.4187
R1148 B.n500 B.n155 30.7255
R1149 B.n506 B.n155 30.7255
R1150 B.n506 B.n150 30.7255
R1151 B.n512 B.n150 30.7255
R1152 B.n512 B.n151 30.7255
R1153 B.n518 B.n143 30.7255
R1154 B.n524 B.n143 30.7255
R1155 B.n524 B.n139 30.7255
R1156 B.n530 B.n139 30.7255
R1157 B.n530 B.n134 30.7255
R1158 B.n536 B.n134 30.7255
R1159 B.n536 B.n135 30.7255
R1160 B.n542 B.n127 30.7255
R1161 B.n548 B.n127 30.7255
R1162 B.n548 B.n123 30.7255
R1163 B.n555 B.n123 30.7255
R1164 B.n561 B.n119 30.7255
R1165 B.n561 B.n4 30.7255
R1166 B.n909 B.n4 30.7255
R1167 B.n909 B.n908 30.7255
R1168 B.n908 B.n907 30.7255
R1169 B.n907 B.n8 30.7255
R1170 B.n570 B.n8 30.7255
R1171 B.n900 B.n899 30.7255
R1172 B.n899 B.n898 30.7255
R1173 B.n898 B.n15 30.7255
R1174 B.n892 B.n15 30.7255
R1175 B.n891 B.n890 30.7255
R1176 B.n890 B.n22 30.7255
R1177 B.n884 B.n22 30.7255
R1178 B.n884 B.n883 30.7255
R1179 B.n883 B.n882 30.7255
R1180 B.n882 B.n29 30.7255
R1181 B.n876 B.n29 30.7255
R1182 B.n875 B.n874 30.7255
R1183 B.n874 B.n36 30.7255
R1184 B.n868 B.n36 30.7255
R1185 B.n868 B.n867 30.7255
R1186 B.n867 B.n866 30.7255
R1187 B.n151 B.t5 23.9479
R1188 B.t9 B.n875 23.9479
R1189 B.n135 B.t2 23.0442
R1190 B.t0 B.n891 23.0442
R1191 B B.n912 18.0485
R1192 B.n555 B.t1 15.8148
R1193 B.n900 B.t3 15.8148
R1194 B.t1 B.n119 14.9112
R1195 B.n570 B.t3 14.9112
R1196 B.n498 B.n153 10.6151
R1197 B.n508 B.n153 10.6151
R1198 B.n509 B.n508 10.6151
R1199 B.n510 B.n509 10.6151
R1200 B.n510 B.n145 10.6151
R1201 B.n520 B.n145 10.6151
R1202 B.n521 B.n520 10.6151
R1203 B.n522 B.n521 10.6151
R1204 B.n522 B.n137 10.6151
R1205 B.n532 B.n137 10.6151
R1206 B.n533 B.n532 10.6151
R1207 B.n534 B.n533 10.6151
R1208 B.n534 B.n129 10.6151
R1209 B.n544 B.n129 10.6151
R1210 B.n545 B.n544 10.6151
R1211 B.n546 B.n545 10.6151
R1212 B.n546 B.n121 10.6151
R1213 B.n557 B.n121 10.6151
R1214 B.n558 B.n557 10.6151
R1215 B.n559 B.n558 10.6151
R1216 B.n559 B.n0 10.6151
R1217 B.n497 B.n496 10.6151
R1218 B.n496 B.n161 10.6151
R1219 B.n491 B.n161 10.6151
R1220 B.n491 B.n490 10.6151
R1221 B.n490 B.n163 10.6151
R1222 B.n485 B.n163 10.6151
R1223 B.n485 B.n484 10.6151
R1224 B.n484 B.n483 10.6151
R1225 B.n483 B.n165 10.6151
R1226 B.n477 B.n165 10.6151
R1227 B.n477 B.n476 10.6151
R1228 B.n476 B.n475 10.6151
R1229 B.n475 B.n167 10.6151
R1230 B.n469 B.n167 10.6151
R1231 B.n469 B.n468 10.6151
R1232 B.n468 B.n467 10.6151
R1233 B.n467 B.n169 10.6151
R1234 B.n461 B.n169 10.6151
R1235 B.n461 B.n460 10.6151
R1236 B.n460 B.n459 10.6151
R1237 B.n459 B.n171 10.6151
R1238 B.n453 B.n171 10.6151
R1239 B.n453 B.n452 10.6151
R1240 B.n452 B.n451 10.6151
R1241 B.n451 B.n173 10.6151
R1242 B.n445 B.n173 10.6151
R1243 B.n445 B.n444 10.6151
R1244 B.n444 B.n443 10.6151
R1245 B.n443 B.n175 10.6151
R1246 B.n437 B.n175 10.6151
R1247 B.n437 B.n436 10.6151
R1248 B.n436 B.n435 10.6151
R1249 B.n435 B.n177 10.6151
R1250 B.n429 B.n177 10.6151
R1251 B.n429 B.n428 10.6151
R1252 B.n428 B.n427 10.6151
R1253 B.n427 B.n179 10.6151
R1254 B.n421 B.n179 10.6151
R1255 B.n421 B.n420 10.6151
R1256 B.n420 B.n419 10.6151
R1257 B.n419 B.n181 10.6151
R1258 B.n413 B.n181 10.6151
R1259 B.n413 B.n412 10.6151
R1260 B.n412 B.n411 10.6151
R1261 B.n411 B.n183 10.6151
R1262 B.n405 B.n183 10.6151
R1263 B.n405 B.n404 10.6151
R1264 B.n404 B.n403 10.6151
R1265 B.n403 B.n185 10.6151
R1266 B.n397 B.n185 10.6151
R1267 B.n397 B.n396 10.6151
R1268 B.n396 B.n395 10.6151
R1269 B.n395 B.n187 10.6151
R1270 B.n389 B.n187 10.6151
R1271 B.n389 B.n388 10.6151
R1272 B.n388 B.n387 10.6151
R1273 B.n387 B.n189 10.6151
R1274 B.n381 B.n189 10.6151
R1275 B.n381 B.n380 10.6151
R1276 B.n380 B.n379 10.6151
R1277 B.n379 B.n191 10.6151
R1278 B.n373 B.n372 10.6151
R1279 B.n372 B.n371 10.6151
R1280 B.n371 B.n196 10.6151
R1281 B.n365 B.n196 10.6151
R1282 B.n365 B.n364 10.6151
R1283 B.n364 B.n363 10.6151
R1284 B.n363 B.n198 10.6151
R1285 B.n357 B.n198 10.6151
R1286 B.n357 B.n356 10.6151
R1287 B.n354 B.n202 10.6151
R1288 B.n348 B.n202 10.6151
R1289 B.n348 B.n347 10.6151
R1290 B.n347 B.n346 10.6151
R1291 B.n346 B.n204 10.6151
R1292 B.n340 B.n204 10.6151
R1293 B.n340 B.n339 10.6151
R1294 B.n339 B.n338 10.6151
R1295 B.n338 B.n206 10.6151
R1296 B.n332 B.n206 10.6151
R1297 B.n332 B.n331 10.6151
R1298 B.n331 B.n330 10.6151
R1299 B.n330 B.n208 10.6151
R1300 B.n324 B.n208 10.6151
R1301 B.n324 B.n323 10.6151
R1302 B.n323 B.n322 10.6151
R1303 B.n322 B.n210 10.6151
R1304 B.n316 B.n210 10.6151
R1305 B.n316 B.n315 10.6151
R1306 B.n315 B.n314 10.6151
R1307 B.n314 B.n212 10.6151
R1308 B.n308 B.n212 10.6151
R1309 B.n308 B.n307 10.6151
R1310 B.n307 B.n306 10.6151
R1311 B.n306 B.n214 10.6151
R1312 B.n300 B.n214 10.6151
R1313 B.n300 B.n299 10.6151
R1314 B.n299 B.n298 10.6151
R1315 B.n298 B.n216 10.6151
R1316 B.n292 B.n216 10.6151
R1317 B.n292 B.n291 10.6151
R1318 B.n291 B.n290 10.6151
R1319 B.n290 B.n218 10.6151
R1320 B.n284 B.n218 10.6151
R1321 B.n284 B.n283 10.6151
R1322 B.n283 B.n282 10.6151
R1323 B.n282 B.n220 10.6151
R1324 B.n276 B.n220 10.6151
R1325 B.n276 B.n275 10.6151
R1326 B.n275 B.n274 10.6151
R1327 B.n274 B.n222 10.6151
R1328 B.n268 B.n222 10.6151
R1329 B.n268 B.n267 10.6151
R1330 B.n267 B.n266 10.6151
R1331 B.n266 B.n224 10.6151
R1332 B.n260 B.n224 10.6151
R1333 B.n260 B.n259 10.6151
R1334 B.n259 B.n258 10.6151
R1335 B.n258 B.n226 10.6151
R1336 B.n252 B.n226 10.6151
R1337 B.n252 B.n251 10.6151
R1338 B.n251 B.n250 10.6151
R1339 B.n250 B.n228 10.6151
R1340 B.n244 B.n228 10.6151
R1341 B.n244 B.n243 10.6151
R1342 B.n243 B.n242 10.6151
R1343 B.n242 B.n230 10.6151
R1344 B.n236 B.n230 10.6151
R1345 B.n236 B.n235 10.6151
R1346 B.n235 B.n234 10.6151
R1347 B.n234 B.n157 10.6151
R1348 B.n503 B.n502 10.6151
R1349 B.n504 B.n503 10.6151
R1350 B.n504 B.n148 10.6151
R1351 B.n514 B.n148 10.6151
R1352 B.n515 B.n514 10.6151
R1353 B.n516 B.n515 10.6151
R1354 B.n516 B.n141 10.6151
R1355 B.n526 B.n141 10.6151
R1356 B.n527 B.n526 10.6151
R1357 B.n528 B.n527 10.6151
R1358 B.n528 B.n132 10.6151
R1359 B.n538 B.n132 10.6151
R1360 B.n539 B.n538 10.6151
R1361 B.n540 B.n539 10.6151
R1362 B.n540 B.n125 10.6151
R1363 B.n550 B.n125 10.6151
R1364 B.n551 B.n550 10.6151
R1365 B.n553 B.n551 10.6151
R1366 B.n553 B.n552 10.6151
R1367 B.n552 B.n117 10.6151
R1368 B.n564 B.n117 10.6151
R1369 B.n565 B.n564 10.6151
R1370 B.n566 B.n565 10.6151
R1371 B.n567 B.n566 10.6151
R1372 B.n568 B.n567 10.6151
R1373 B.n572 B.n568 10.6151
R1374 B.n573 B.n572 10.6151
R1375 B.n574 B.n573 10.6151
R1376 B.n575 B.n574 10.6151
R1377 B.n577 B.n575 10.6151
R1378 B.n578 B.n577 10.6151
R1379 B.n579 B.n578 10.6151
R1380 B.n580 B.n579 10.6151
R1381 B.n582 B.n580 10.6151
R1382 B.n583 B.n582 10.6151
R1383 B.n584 B.n583 10.6151
R1384 B.n585 B.n584 10.6151
R1385 B.n587 B.n585 10.6151
R1386 B.n588 B.n587 10.6151
R1387 B.n589 B.n588 10.6151
R1388 B.n590 B.n589 10.6151
R1389 B.n592 B.n590 10.6151
R1390 B.n593 B.n592 10.6151
R1391 B.n594 B.n593 10.6151
R1392 B.n595 B.n594 10.6151
R1393 B.n904 B.n1 10.6151
R1394 B.n904 B.n903 10.6151
R1395 B.n903 B.n902 10.6151
R1396 B.n902 B.n10 10.6151
R1397 B.n896 B.n10 10.6151
R1398 B.n896 B.n895 10.6151
R1399 B.n895 B.n894 10.6151
R1400 B.n894 B.n17 10.6151
R1401 B.n888 B.n17 10.6151
R1402 B.n888 B.n887 10.6151
R1403 B.n887 B.n886 10.6151
R1404 B.n886 B.n24 10.6151
R1405 B.n880 B.n24 10.6151
R1406 B.n880 B.n879 10.6151
R1407 B.n879 B.n878 10.6151
R1408 B.n878 B.n31 10.6151
R1409 B.n872 B.n31 10.6151
R1410 B.n872 B.n871 10.6151
R1411 B.n871 B.n870 10.6151
R1412 B.n870 B.n38 10.6151
R1413 B.n864 B.n38 10.6151
R1414 B.n863 B.n862 10.6151
R1415 B.n862 B.n45 10.6151
R1416 B.n856 B.n45 10.6151
R1417 B.n856 B.n855 10.6151
R1418 B.n855 B.n854 10.6151
R1419 B.n854 B.n47 10.6151
R1420 B.n848 B.n47 10.6151
R1421 B.n848 B.n847 10.6151
R1422 B.n847 B.n846 10.6151
R1423 B.n846 B.n49 10.6151
R1424 B.n840 B.n49 10.6151
R1425 B.n840 B.n839 10.6151
R1426 B.n839 B.n838 10.6151
R1427 B.n838 B.n51 10.6151
R1428 B.n832 B.n51 10.6151
R1429 B.n832 B.n831 10.6151
R1430 B.n831 B.n830 10.6151
R1431 B.n830 B.n53 10.6151
R1432 B.n824 B.n53 10.6151
R1433 B.n824 B.n823 10.6151
R1434 B.n823 B.n822 10.6151
R1435 B.n822 B.n55 10.6151
R1436 B.n816 B.n55 10.6151
R1437 B.n816 B.n815 10.6151
R1438 B.n815 B.n814 10.6151
R1439 B.n814 B.n57 10.6151
R1440 B.n808 B.n57 10.6151
R1441 B.n808 B.n807 10.6151
R1442 B.n807 B.n806 10.6151
R1443 B.n806 B.n59 10.6151
R1444 B.n800 B.n59 10.6151
R1445 B.n800 B.n799 10.6151
R1446 B.n799 B.n798 10.6151
R1447 B.n798 B.n61 10.6151
R1448 B.n792 B.n61 10.6151
R1449 B.n792 B.n791 10.6151
R1450 B.n791 B.n790 10.6151
R1451 B.n790 B.n63 10.6151
R1452 B.n784 B.n63 10.6151
R1453 B.n784 B.n783 10.6151
R1454 B.n783 B.n782 10.6151
R1455 B.n782 B.n65 10.6151
R1456 B.n776 B.n65 10.6151
R1457 B.n776 B.n775 10.6151
R1458 B.n775 B.n774 10.6151
R1459 B.n774 B.n67 10.6151
R1460 B.n768 B.n67 10.6151
R1461 B.n768 B.n767 10.6151
R1462 B.n767 B.n766 10.6151
R1463 B.n766 B.n69 10.6151
R1464 B.n760 B.n69 10.6151
R1465 B.n760 B.n759 10.6151
R1466 B.n759 B.n758 10.6151
R1467 B.n758 B.n71 10.6151
R1468 B.n752 B.n71 10.6151
R1469 B.n752 B.n751 10.6151
R1470 B.n751 B.n750 10.6151
R1471 B.n750 B.n73 10.6151
R1472 B.n744 B.n73 10.6151
R1473 B.n744 B.n743 10.6151
R1474 B.n743 B.n742 10.6151
R1475 B.n738 B.n737 10.6151
R1476 B.n737 B.n79 10.6151
R1477 B.n732 B.n79 10.6151
R1478 B.n732 B.n731 10.6151
R1479 B.n731 B.n730 10.6151
R1480 B.n730 B.n81 10.6151
R1481 B.n724 B.n81 10.6151
R1482 B.n724 B.n723 10.6151
R1483 B.n723 B.n722 10.6151
R1484 B.n718 B.n717 10.6151
R1485 B.n717 B.n87 10.6151
R1486 B.n712 B.n87 10.6151
R1487 B.n712 B.n711 10.6151
R1488 B.n711 B.n710 10.6151
R1489 B.n710 B.n89 10.6151
R1490 B.n704 B.n89 10.6151
R1491 B.n704 B.n703 10.6151
R1492 B.n703 B.n702 10.6151
R1493 B.n702 B.n91 10.6151
R1494 B.n696 B.n91 10.6151
R1495 B.n696 B.n695 10.6151
R1496 B.n695 B.n694 10.6151
R1497 B.n694 B.n93 10.6151
R1498 B.n688 B.n93 10.6151
R1499 B.n688 B.n687 10.6151
R1500 B.n687 B.n686 10.6151
R1501 B.n686 B.n95 10.6151
R1502 B.n680 B.n95 10.6151
R1503 B.n680 B.n679 10.6151
R1504 B.n679 B.n678 10.6151
R1505 B.n678 B.n97 10.6151
R1506 B.n672 B.n97 10.6151
R1507 B.n672 B.n671 10.6151
R1508 B.n671 B.n670 10.6151
R1509 B.n670 B.n99 10.6151
R1510 B.n664 B.n99 10.6151
R1511 B.n664 B.n663 10.6151
R1512 B.n663 B.n662 10.6151
R1513 B.n662 B.n101 10.6151
R1514 B.n656 B.n101 10.6151
R1515 B.n656 B.n655 10.6151
R1516 B.n655 B.n654 10.6151
R1517 B.n654 B.n103 10.6151
R1518 B.n648 B.n103 10.6151
R1519 B.n648 B.n647 10.6151
R1520 B.n647 B.n646 10.6151
R1521 B.n646 B.n105 10.6151
R1522 B.n640 B.n105 10.6151
R1523 B.n640 B.n639 10.6151
R1524 B.n639 B.n638 10.6151
R1525 B.n638 B.n107 10.6151
R1526 B.n632 B.n107 10.6151
R1527 B.n632 B.n631 10.6151
R1528 B.n631 B.n630 10.6151
R1529 B.n630 B.n109 10.6151
R1530 B.n624 B.n109 10.6151
R1531 B.n624 B.n623 10.6151
R1532 B.n623 B.n622 10.6151
R1533 B.n622 B.n111 10.6151
R1534 B.n616 B.n111 10.6151
R1535 B.n616 B.n615 10.6151
R1536 B.n615 B.n614 10.6151
R1537 B.n614 B.n113 10.6151
R1538 B.n608 B.n113 10.6151
R1539 B.n608 B.n607 10.6151
R1540 B.n607 B.n606 10.6151
R1541 B.n606 B.n115 10.6151
R1542 B.n600 B.n115 10.6151
R1543 B.n600 B.n599 10.6151
R1544 B.n599 B.n598 10.6151
R1545 B.n195 B.n191 9.36635
R1546 B.n355 B.n354 9.36635
R1547 B.n742 B.n77 9.36635
R1548 B.n718 B.n85 9.36635
R1549 B.n912 B.n0 8.11757
R1550 B.n912 B.n1 8.11757
R1551 B.n542 B.t2 7.68175
R1552 B.n892 B.t0 7.68175
R1553 B.n518 B.t5 6.77807
R1554 B.n876 B.t9 6.77807
R1555 B.n373 B.n195 1.24928
R1556 B.n356 B.n355 1.24928
R1557 B.n738 B.n77 1.24928
R1558 B.n722 B.n85 1.24928
R1559 VN.n0 VN.t0 393.598
R1560 VN.n1 VN.t2 393.598
R1561 VN.n0 VN.t1 393.372
R1562 VN.n1 VN.t3 393.372
R1563 VN VN.n1 65.9973
R1564 VN VN.n0 18.0466
R1565 VDD2.n2 VDD2.n0 106.675
R1566 VDD2.n2 VDD2.n1 62.3327
R1567 VDD2.n1 VDD2.t0 1.03878
R1568 VDD2.n1 VDD2.t1 1.03878
R1569 VDD2.n0 VDD2.t3 1.03878
R1570 VDD2.n0 VDD2.t2 1.03878
R1571 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 5.59824f
C1 VTAIL VDD2 8.02008f
C2 VTAIL VP 5.61235f
C3 VDD2 VN 6.18597f
C4 VN VP 6.555779f
C5 VDD1 VTAIL 7.97466f
C6 VDD1 VN 0.14763f
C7 VDD2 VP 0.310762f
C8 VDD1 VDD2 0.706218f
C9 VDD1 VP 6.348701f
C10 VDD2 B 3.581594f
C11 VDD1 B 8.07815f
C12 VTAIL B 13.349462f
C13 VN B 9.380549f
C14 VP B 6.621935f
C15 VDD2.t3 B 0.403563f
C16 VDD2.t2 B 0.403563f
C17 VDD2.n0 B 4.54609f
C18 VDD2.t0 B 0.403563f
C19 VDD2.t1 B 0.403563f
C20 VDD2.n1 B 3.69271f
C21 VDD2.n2 B 4.22067f
C22 VN.t0 B 2.61676f
C23 VN.t1 B 2.61616f
C24 VN.n0 B 1.88471f
C25 VN.t2 B 2.61676f
C26 VN.t3 B 2.61616f
C27 VN.n1 B 3.38755f
C28 VTAIL.t3 B 2.59047f
C29 VTAIL.n0 B 0.256525f
C30 VTAIL.t5 B 2.59047f
C31 VTAIL.n1 B 0.28749f
C32 VTAIL.t4 B 2.59047f
C33 VTAIL.n2 B 1.33158f
C34 VTAIL.t2 B 2.59049f
C35 VTAIL.n3 B 1.33156f
C36 VTAIL.t1 B 2.59049f
C37 VTAIL.n4 B 0.287471f
C38 VTAIL.t7 B 2.59049f
C39 VTAIL.n5 B 0.287471f
C40 VTAIL.t6 B 2.59047f
C41 VTAIL.n6 B 1.33158f
C42 VTAIL.t0 B 2.59047f
C43 VTAIL.n7 B 1.29498f
C44 VDD1.t3 B 0.403594f
C45 VDD1.t2 B 0.403594f
C46 VDD1.n0 B 3.69331f
C47 VDD1.t0 B 0.403594f
C48 VDD1.t1 B 0.403594f
C49 VDD1.n1 B 4.57456f
C50 VP.n0 B 0.037516f
C51 VP.t2 B 2.5412f
C52 VP.n1 B 0.061445f
C53 VP.t0 B 2.63848f
C54 VP.t1 B 2.63788f
C55 VP.n2 B 3.39462f
C56 VP.t3 B 2.5412f
C57 VP.n3 B 0.969293f
C58 VP.n4 B 2.49108f
C59 VP.n5 B 0.037516f
C60 VP.n6 B 0.037516f
C61 VP.n7 B 0.030328f
C62 VP.n8 B 0.061445f
C63 VP.n9 B 0.969293f
C64 VP.n10 B 0.03326f
.ends

