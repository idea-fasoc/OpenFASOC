* NGSPICE file created from diff_pair_sample_0605.ext - technology: sky130A

.subckt diff_pair_sample_0605 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0 ps=0 w=5.37 l=3.12
X1 B.t8 B.t6 B.t7 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0 ps=0 w=5.37 l=3.12
X2 VDD1.t7 VP.t0 VTAIL.t9 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=2.0943 ps=11.52 w=5.37 l=3.12
X3 VDD1.t6 VP.t1 VTAIL.t12 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X4 VTAIL.t7 VN.t0 VDD2.t7 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0.88605 ps=5.7 w=5.37 l=3.12
X5 B.t5 B.t3 B.t4 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0 ps=0 w=5.37 l=3.12
X6 VTAIL.t4 VN.t1 VDD2.t6 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X7 B.t2 B.t0 B.t1 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0 ps=0 w=5.37 l=3.12
X8 VDD2.t5 VN.t2 VTAIL.t2 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=2.0943 ps=11.52 w=5.37 l=3.12
X9 VTAIL.t3 VN.t3 VDD2.t4 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X10 VTAIL.t10 VP.t2 VDD1.t5 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X11 VTAIL.t15 VP.t3 VDD1.t4 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0.88605 ps=5.7 w=5.37 l=3.12
X12 VTAIL.t13 VP.t4 VDD1.t3 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0.88605 ps=5.7 w=5.37 l=3.12
X13 VTAIL.t6 VN.t4 VDD2.t3 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=2.0943 pd=11.52 as=0.88605 ps=5.7 w=5.37 l=3.12
X14 VDD1.t2 VP.t5 VTAIL.t14 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X15 VTAIL.t8 VP.t6 VDD1.t1 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X16 VDD2.t2 VN.t5 VTAIL.t0 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X17 VDD2.t1 VN.t6 VTAIL.t5 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=0.88605 ps=5.7 w=5.37 l=3.12
X18 VDD1.t0 VP.t7 VTAIL.t11 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=2.0943 ps=11.52 w=5.37 l=3.12
X19 VDD2.t0 VN.t7 VTAIL.t1 w_n4420_n2042# sky130_fd_pr__pfet_01v8 ad=0.88605 pd=5.7 as=2.0943 ps=11.52 w=5.37 l=3.12
R0 B.n532 B.n63 585
R1 B.n534 B.n533 585
R2 B.n535 B.n62 585
R3 B.n537 B.n536 585
R4 B.n538 B.n61 585
R5 B.n540 B.n539 585
R6 B.n541 B.n60 585
R7 B.n543 B.n542 585
R8 B.n544 B.n59 585
R9 B.n546 B.n545 585
R10 B.n547 B.n58 585
R11 B.n549 B.n548 585
R12 B.n550 B.n57 585
R13 B.n552 B.n551 585
R14 B.n553 B.n56 585
R15 B.n555 B.n554 585
R16 B.n556 B.n55 585
R17 B.n558 B.n557 585
R18 B.n559 B.n54 585
R19 B.n561 B.n560 585
R20 B.n562 B.n53 585
R21 B.n564 B.n563 585
R22 B.n566 B.n50 585
R23 B.n568 B.n567 585
R24 B.n569 B.n49 585
R25 B.n571 B.n570 585
R26 B.n572 B.n48 585
R27 B.n574 B.n573 585
R28 B.n575 B.n47 585
R29 B.n577 B.n576 585
R30 B.n578 B.n43 585
R31 B.n580 B.n579 585
R32 B.n581 B.n42 585
R33 B.n583 B.n582 585
R34 B.n584 B.n41 585
R35 B.n586 B.n585 585
R36 B.n587 B.n40 585
R37 B.n589 B.n588 585
R38 B.n590 B.n39 585
R39 B.n592 B.n591 585
R40 B.n593 B.n38 585
R41 B.n595 B.n594 585
R42 B.n596 B.n37 585
R43 B.n598 B.n597 585
R44 B.n599 B.n36 585
R45 B.n601 B.n600 585
R46 B.n602 B.n35 585
R47 B.n604 B.n603 585
R48 B.n605 B.n34 585
R49 B.n607 B.n606 585
R50 B.n608 B.n33 585
R51 B.n610 B.n609 585
R52 B.n611 B.n32 585
R53 B.n613 B.n612 585
R54 B.n531 B.n530 585
R55 B.n529 B.n64 585
R56 B.n528 B.n527 585
R57 B.n526 B.n65 585
R58 B.n525 B.n524 585
R59 B.n523 B.n66 585
R60 B.n522 B.n521 585
R61 B.n520 B.n67 585
R62 B.n519 B.n518 585
R63 B.n517 B.n68 585
R64 B.n516 B.n515 585
R65 B.n514 B.n69 585
R66 B.n513 B.n512 585
R67 B.n511 B.n70 585
R68 B.n510 B.n509 585
R69 B.n508 B.n71 585
R70 B.n507 B.n506 585
R71 B.n505 B.n72 585
R72 B.n504 B.n503 585
R73 B.n502 B.n73 585
R74 B.n501 B.n500 585
R75 B.n499 B.n74 585
R76 B.n498 B.n497 585
R77 B.n496 B.n75 585
R78 B.n495 B.n494 585
R79 B.n493 B.n76 585
R80 B.n492 B.n491 585
R81 B.n490 B.n77 585
R82 B.n489 B.n488 585
R83 B.n487 B.n78 585
R84 B.n486 B.n485 585
R85 B.n484 B.n79 585
R86 B.n483 B.n482 585
R87 B.n481 B.n80 585
R88 B.n480 B.n479 585
R89 B.n478 B.n81 585
R90 B.n477 B.n476 585
R91 B.n475 B.n82 585
R92 B.n474 B.n473 585
R93 B.n472 B.n83 585
R94 B.n471 B.n470 585
R95 B.n469 B.n84 585
R96 B.n468 B.n467 585
R97 B.n466 B.n85 585
R98 B.n465 B.n464 585
R99 B.n463 B.n86 585
R100 B.n462 B.n461 585
R101 B.n460 B.n87 585
R102 B.n459 B.n458 585
R103 B.n457 B.n88 585
R104 B.n456 B.n455 585
R105 B.n454 B.n89 585
R106 B.n453 B.n452 585
R107 B.n451 B.n90 585
R108 B.n450 B.n449 585
R109 B.n448 B.n91 585
R110 B.n447 B.n446 585
R111 B.n445 B.n92 585
R112 B.n444 B.n443 585
R113 B.n442 B.n93 585
R114 B.n441 B.n440 585
R115 B.n439 B.n94 585
R116 B.n438 B.n437 585
R117 B.n436 B.n95 585
R118 B.n435 B.n434 585
R119 B.n433 B.n96 585
R120 B.n432 B.n431 585
R121 B.n430 B.n97 585
R122 B.n429 B.n428 585
R123 B.n427 B.n98 585
R124 B.n426 B.n425 585
R125 B.n424 B.n99 585
R126 B.n423 B.n422 585
R127 B.n421 B.n100 585
R128 B.n420 B.n419 585
R129 B.n418 B.n101 585
R130 B.n417 B.n416 585
R131 B.n415 B.n102 585
R132 B.n414 B.n413 585
R133 B.n412 B.n103 585
R134 B.n411 B.n410 585
R135 B.n409 B.n104 585
R136 B.n408 B.n407 585
R137 B.n406 B.n105 585
R138 B.n405 B.n404 585
R139 B.n403 B.n106 585
R140 B.n402 B.n401 585
R141 B.n400 B.n107 585
R142 B.n399 B.n398 585
R143 B.n397 B.n108 585
R144 B.n396 B.n395 585
R145 B.n394 B.n109 585
R146 B.n393 B.n392 585
R147 B.n391 B.n110 585
R148 B.n390 B.n389 585
R149 B.n388 B.n111 585
R150 B.n387 B.n386 585
R151 B.n385 B.n112 585
R152 B.n384 B.n383 585
R153 B.n382 B.n113 585
R154 B.n381 B.n380 585
R155 B.n379 B.n114 585
R156 B.n378 B.n377 585
R157 B.n376 B.n115 585
R158 B.n375 B.n374 585
R159 B.n373 B.n116 585
R160 B.n372 B.n371 585
R161 B.n370 B.n117 585
R162 B.n369 B.n368 585
R163 B.n367 B.n118 585
R164 B.n366 B.n365 585
R165 B.n364 B.n119 585
R166 B.n363 B.n362 585
R167 B.n361 B.n120 585
R168 B.n360 B.n359 585
R169 B.n358 B.n121 585
R170 B.n357 B.n356 585
R171 B.n355 B.n122 585
R172 B.n354 B.n353 585
R173 B.n271 B.n154 585
R174 B.n273 B.n272 585
R175 B.n274 B.n153 585
R176 B.n276 B.n275 585
R177 B.n277 B.n152 585
R178 B.n279 B.n278 585
R179 B.n280 B.n151 585
R180 B.n282 B.n281 585
R181 B.n283 B.n150 585
R182 B.n285 B.n284 585
R183 B.n286 B.n149 585
R184 B.n288 B.n287 585
R185 B.n289 B.n148 585
R186 B.n291 B.n290 585
R187 B.n292 B.n147 585
R188 B.n294 B.n293 585
R189 B.n295 B.n146 585
R190 B.n297 B.n296 585
R191 B.n298 B.n145 585
R192 B.n300 B.n299 585
R193 B.n301 B.n144 585
R194 B.n303 B.n302 585
R195 B.n305 B.n304 585
R196 B.n306 B.n140 585
R197 B.n308 B.n307 585
R198 B.n309 B.n139 585
R199 B.n311 B.n310 585
R200 B.n312 B.n138 585
R201 B.n314 B.n313 585
R202 B.n315 B.n137 585
R203 B.n317 B.n316 585
R204 B.n318 B.n134 585
R205 B.n321 B.n320 585
R206 B.n322 B.n133 585
R207 B.n324 B.n323 585
R208 B.n325 B.n132 585
R209 B.n327 B.n326 585
R210 B.n328 B.n131 585
R211 B.n330 B.n329 585
R212 B.n331 B.n130 585
R213 B.n333 B.n332 585
R214 B.n334 B.n129 585
R215 B.n336 B.n335 585
R216 B.n337 B.n128 585
R217 B.n339 B.n338 585
R218 B.n340 B.n127 585
R219 B.n342 B.n341 585
R220 B.n343 B.n126 585
R221 B.n345 B.n344 585
R222 B.n346 B.n125 585
R223 B.n348 B.n347 585
R224 B.n349 B.n124 585
R225 B.n351 B.n350 585
R226 B.n352 B.n123 585
R227 B.n270 B.n269 585
R228 B.n268 B.n155 585
R229 B.n267 B.n266 585
R230 B.n265 B.n156 585
R231 B.n264 B.n263 585
R232 B.n262 B.n157 585
R233 B.n261 B.n260 585
R234 B.n259 B.n158 585
R235 B.n258 B.n257 585
R236 B.n256 B.n159 585
R237 B.n255 B.n254 585
R238 B.n253 B.n160 585
R239 B.n252 B.n251 585
R240 B.n250 B.n161 585
R241 B.n249 B.n248 585
R242 B.n247 B.n162 585
R243 B.n246 B.n245 585
R244 B.n244 B.n163 585
R245 B.n243 B.n242 585
R246 B.n241 B.n164 585
R247 B.n240 B.n239 585
R248 B.n238 B.n165 585
R249 B.n237 B.n236 585
R250 B.n235 B.n166 585
R251 B.n234 B.n233 585
R252 B.n232 B.n167 585
R253 B.n231 B.n230 585
R254 B.n229 B.n168 585
R255 B.n228 B.n227 585
R256 B.n226 B.n169 585
R257 B.n225 B.n224 585
R258 B.n223 B.n170 585
R259 B.n222 B.n221 585
R260 B.n220 B.n171 585
R261 B.n219 B.n218 585
R262 B.n217 B.n172 585
R263 B.n216 B.n215 585
R264 B.n214 B.n173 585
R265 B.n213 B.n212 585
R266 B.n211 B.n174 585
R267 B.n210 B.n209 585
R268 B.n208 B.n175 585
R269 B.n207 B.n206 585
R270 B.n205 B.n176 585
R271 B.n204 B.n203 585
R272 B.n202 B.n177 585
R273 B.n201 B.n200 585
R274 B.n199 B.n178 585
R275 B.n198 B.n197 585
R276 B.n196 B.n179 585
R277 B.n195 B.n194 585
R278 B.n193 B.n180 585
R279 B.n192 B.n191 585
R280 B.n190 B.n181 585
R281 B.n189 B.n188 585
R282 B.n187 B.n182 585
R283 B.n186 B.n185 585
R284 B.n184 B.n183 585
R285 B.n2 B.n0 585
R286 B.n701 B.n1 585
R287 B.n700 B.n699 585
R288 B.n698 B.n3 585
R289 B.n697 B.n696 585
R290 B.n695 B.n4 585
R291 B.n694 B.n693 585
R292 B.n692 B.n5 585
R293 B.n691 B.n690 585
R294 B.n689 B.n6 585
R295 B.n688 B.n687 585
R296 B.n686 B.n7 585
R297 B.n685 B.n684 585
R298 B.n683 B.n8 585
R299 B.n682 B.n681 585
R300 B.n680 B.n9 585
R301 B.n679 B.n678 585
R302 B.n677 B.n10 585
R303 B.n676 B.n675 585
R304 B.n674 B.n11 585
R305 B.n673 B.n672 585
R306 B.n671 B.n12 585
R307 B.n670 B.n669 585
R308 B.n668 B.n13 585
R309 B.n667 B.n666 585
R310 B.n665 B.n14 585
R311 B.n664 B.n663 585
R312 B.n662 B.n15 585
R313 B.n661 B.n660 585
R314 B.n659 B.n16 585
R315 B.n658 B.n657 585
R316 B.n656 B.n17 585
R317 B.n655 B.n654 585
R318 B.n653 B.n18 585
R319 B.n652 B.n651 585
R320 B.n650 B.n19 585
R321 B.n649 B.n648 585
R322 B.n647 B.n20 585
R323 B.n646 B.n645 585
R324 B.n644 B.n21 585
R325 B.n643 B.n642 585
R326 B.n641 B.n22 585
R327 B.n640 B.n639 585
R328 B.n638 B.n23 585
R329 B.n637 B.n636 585
R330 B.n635 B.n24 585
R331 B.n634 B.n633 585
R332 B.n632 B.n25 585
R333 B.n631 B.n630 585
R334 B.n629 B.n26 585
R335 B.n628 B.n627 585
R336 B.n626 B.n27 585
R337 B.n625 B.n624 585
R338 B.n623 B.n28 585
R339 B.n622 B.n621 585
R340 B.n620 B.n29 585
R341 B.n619 B.n618 585
R342 B.n617 B.n30 585
R343 B.n616 B.n615 585
R344 B.n614 B.n31 585
R345 B.n703 B.n702 585
R346 B.n269 B.n154 458.866
R347 B.n612 B.n31 458.866
R348 B.n353 B.n352 458.866
R349 B.n532 B.n531 458.866
R350 B.n135 B.t11 324.303
R351 B.n51 B.t1 324.303
R352 B.n141 B.t8 324.303
R353 B.n44 B.t4 324.303
R354 B.n136 B.t10 257.394
R355 B.n52 B.t2 257.394
R356 B.n142 B.t7 257.394
R357 B.n45 B.t5 257.394
R358 B.n135 B.t9 250.196
R359 B.n141 B.t6 250.196
R360 B.n44 B.t3 250.196
R361 B.n51 B.t0 250.196
R362 B.n269 B.n268 163.367
R363 B.n268 B.n267 163.367
R364 B.n267 B.n156 163.367
R365 B.n263 B.n156 163.367
R366 B.n263 B.n262 163.367
R367 B.n262 B.n261 163.367
R368 B.n261 B.n158 163.367
R369 B.n257 B.n158 163.367
R370 B.n257 B.n256 163.367
R371 B.n256 B.n255 163.367
R372 B.n255 B.n160 163.367
R373 B.n251 B.n160 163.367
R374 B.n251 B.n250 163.367
R375 B.n250 B.n249 163.367
R376 B.n249 B.n162 163.367
R377 B.n245 B.n162 163.367
R378 B.n245 B.n244 163.367
R379 B.n244 B.n243 163.367
R380 B.n243 B.n164 163.367
R381 B.n239 B.n164 163.367
R382 B.n239 B.n238 163.367
R383 B.n238 B.n237 163.367
R384 B.n237 B.n166 163.367
R385 B.n233 B.n166 163.367
R386 B.n233 B.n232 163.367
R387 B.n232 B.n231 163.367
R388 B.n231 B.n168 163.367
R389 B.n227 B.n168 163.367
R390 B.n227 B.n226 163.367
R391 B.n226 B.n225 163.367
R392 B.n225 B.n170 163.367
R393 B.n221 B.n170 163.367
R394 B.n221 B.n220 163.367
R395 B.n220 B.n219 163.367
R396 B.n219 B.n172 163.367
R397 B.n215 B.n172 163.367
R398 B.n215 B.n214 163.367
R399 B.n214 B.n213 163.367
R400 B.n213 B.n174 163.367
R401 B.n209 B.n174 163.367
R402 B.n209 B.n208 163.367
R403 B.n208 B.n207 163.367
R404 B.n207 B.n176 163.367
R405 B.n203 B.n176 163.367
R406 B.n203 B.n202 163.367
R407 B.n202 B.n201 163.367
R408 B.n201 B.n178 163.367
R409 B.n197 B.n178 163.367
R410 B.n197 B.n196 163.367
R411 B.n196 B.n195 163.367
R412 B.n195 B.n180 163.367
R413 B.n191 B.n180 163.367
R414 B.n191 B.n190 163.367
R415 B.n190 B.n189 163.367
R416 B.n189 B.n182 163.367
R417 B.n185 B.n182 163.367
R418 B.n185 B.n184 163.367
R419 B.n184 B.n2 163.367
R420 B.n702 B.n2 163.367
R421 B.n702 B.n701 163.367
R422 B.n701 B.n700 163.367
R423 B.n700 B.n3 163.367
R424 B.n696 B.n3 163.367
R425 B.n696 B.n695 163.367
R426 B.n695 B.n694 163.367
R427 B.n694 B.n5 163.367
R428 B.n690 B.n5 163.367
R429 B.n690 B.n689 163.367
R430 B.n689 B.n688 163.367
R431 B.n688 B.n7 163.367
R432 B.n684 B.n7 163.367
R433 B.n684 B.n683 163.367
R434 B.n683 B.n682 163.367
R435 B.n682 B.n9 163.367
R436 B.n678 B.n9 163.367
R437 B.n678 B.n677 163.367
R438 B.n677 B.n676 163.367
R439 B.n676 B.n11 163.367
R440 B.n672 B.n11 163.367
R441 B.n672 B.n671 163.367
R442 B.n671 B.n670 163.367
R443 B.n670 B.n13 163.367
R444 B.n666 B.n13 163.367
R445 B.n666 B.n665 163.367
R446 B.n665 B.n664 163.367
R447 B.n664 B.n15 163.367
R448 B.n660 B.n15 163.367
R449 B.n660 B.n659 163.367
R450 B.n659 B.n658 163.367
R451 B.n658 B.n17 163.367
R452 B.n654 B.n17 163.367
R453 B.n654 B.n653 163.367
R454 B.n653 B.n652 163.367
R455 B.n652 B.n19 163.367
R456 B.n648 B.n19 163.367
R457 B.n648 B.n647 163.367
R458 B.n647 B.n646 163.367
R459 B.n646 B.n21 163.367
R460 B.n642 B.n21 163.367
R461 B.n642 B.n641 163.367
R462 B.n641 B.n640 163.367
R463 B.n640 B.n23 163.367
R464 B.n636 B.n23 163.367
R465 B.n636 B.n635 163.367
R466 B.n635 B.n634 163.367
R467 B.n634 B.n25 163.367
R468 B.n630 B.n25 163.367
R469 B.n630 B.n629 163.367
R470 B.n629 B.n628 163.367
R471 B.n628 B.n27 163.367
R472 B.n624 B.n27 163.367
R473 B.n624 B.n623 163.367
R474 B.n623 B.n622 163.367
R475 B.n622 B.n29 163.367
R476 B.n618 B.n29 163.367
R477 B.n618 B.n617 163.367
R478 B.n617 B.n616 163.367
R479 B.n616 B.n31 163.367
R480 B.n273 B.n154 163.367
R481 B.n274 B.n273 163.367
R482 B.n275 B.n274 163.367
R483 B.n275 B.n152 163.367
R484 B.n279 B.n152 163.367
R485 B.n280 B.n279 163.367
R486 B.n281 B.n280 163.367
R487 B.n281 B.n150 163.367
R488 B.n285 B.n150 163.367
R489 B.n286 B.n285 163.367
R490 B.n287 B.n286 163.367
R491 B.n287 B.n148 163.367
R492 B.n291 B.n148 163.367
R493 B.n292 B.n291 163.367
R494 B.n293 B.n292 163.367
R495 B.n293 B.n146 163.367
R496 B.n297 B.n146 163.367
R497 B.n298 B.n297 163.367
R498 B.n299 B.n298 163.367
R499 B.n299 B.n144 163.367
R500 B.n303 B.n144 163.367
R501 B.n304 B.n303 163.367
R502 B.n304 B.n140 163.367
R503 B.n308 B.n140 163.367
R504 B.n309 B.n308 163.367
R505 B.n310 B.n309 163.367
R506 B.n310 B.n138 163.367
R507 B.n314 B.n138 163.367
R508 B.n315 B.n314 163.367
R509 B.n316 B.n315 163.367
R510 B.n316 B.n134 163.367
R511 B.n321 B.n134 163.367
R512 B.n322 B.n321 163.367
R513 B.n323 B.n322 163.367
R514 B.n323 B.n132 163.367
R515 B.n327 B.n132 163.367
R516 B.n328 B.n327 163.367
R517 B.n329 B.n328 163.367
R518 B.n329 B.n130 163.367
R519 B.n333 B.n130 163.367
R520 B.n334 B.n333 163.367
R521 B.n335 B.n334 163.367
R522 B.n335 B.n128 163.367
R523 B.n339 B.n128 163.367
R524 B.n340 B.n339 163.367
R525 B.n341 B.n340 163.367
R526 B.n341 B.n126 163.367
R527 B.n345 B.n126 163.367
R528 B.n346 B.n345 163.367
R529 B.n347 B.n346 163.367
R530 B.n347 B.n124 163.367
R531 B.n351 B.n124 163.367
R532 B.n352 B.n351 163.367
R533 B.n353 B.n122 163.367
R534 B.n357 B.n122 163.367
R535 B.n358 B.n357 163.367
R536 B.n359 B.n358 163.367
R537 B.n359 B.n120 163.367
R538 B.n363 B.n120 163.367
R539 B.n364 B.n363 163.367
R540 B.n365 B.n364 163.367
R541 B.n365 B.n118 163.367
R542 B.n369 B.n118 163.367
R543 B.n370 B.n369 163.367
R544 B.n371 B.n370 163.367
R545 B.n371 B.n116 163.367
R546 B.n375 B.n116 163.367
R547 B.n376 B.n375 163.367
R548 B.n377 B.n376 163.367
R549 B.n377 B.n114 163.367
R550 B.n381 B.n114 163.367
R551 B.n382 B.n381 163.367
R552 B.n383 B.n382 163.367
R553 B.n383 B.n112 163.367
R554 B.n387 B.n112 163.367
R555 B.n388 B.n387 163.367
R556 B.n389 B.n388 163.367
R557 B.n389 B.n110 163.367
R558 B.n393 B.n110 163.367
R559 B.n394 B.n393 163.367
R560 B.n395 B.n394 163.367
R561 B.n395 B.n108 163.367
R562 B.n399 B.n108 163.367
R563 B.n400 B.n399 163.367
R564 B.n401 B.n400 163.367
R565 B.n401 B.n106 163.367
R566 B.n405 B.n106 163.367
R567 B.n406 B.n405 163.367
R568 B.n407 B.n406 163.367
R569 B.n407 B.n104 163.367
R570 B.n411 B.n104 163.367
R571 B.n412 B.n411 163.367
R572 B.n413 B.n412 163.367
R573 B.n413 B.n102 163.367
R574 B.n417 B.n102 163.367
R575 B.n418 B.n417 163.367
R576 B.n419 B.n418 163.367
R577 B.n419 B.n100 163.367
R578 B.n423 B.n100 163.367
R579 B.n424 B.n423 163.367
R580 B.n425 B.n424 163.367
R581 B.n425 B.n98 163.367
R582 B.n429 B.n98 163.367
R583 B.n430 B.n429 163.367
R584 B.n431 B.n430 163.367
R585 B.n431 B.n96 163.367
R586 B.n435 B.n96 163.367
R587 B.n436 B.n435 163.367
R588 B.n437 B.n436 163.367
R589 B.n437 B.n94 163.367
R590 B.n441 B.n94 163.367
R591 B.n442 B.n441 163.367
R592 B.n443 B.n442 163.367
R593 B.n443 B.n92 163.367
R594 B.n447 B.n92 163.367
R595 B.n448 B.n447 163.367
R596 B.n449 B.n448 163.367
R597 B.n449 B.n90 163.367
R598 B.n453 B.n90 163.367
R599 B.n454 B.n453 163.367
R600 B.n455 B.n454 163.367
R601 B.n455 B.n88 163.367
R602 B.n459 B.n88 163.367
R603 B.n460 B.n459 163.367
R604 B.n461 B.n460 163.367
R605 B.n461 B.n86 163.367
R606 B.n465 B.n86 163.367
R607 B.n466 B.n465 163.367
R608 B.n467 B.n466 163.367
R609 B.n467 B.n84 163.367
R610 B.n471 B.n84 163.367
R611 B.n472 B.n471 163.367
R612 B.n473 B.n472 163.367
R613 B.n473 B.n82 163.367
R614 B.n477 B.n82 163.367
R615 B.n478 B.n477 163.367
R616 B.n479 B.n478 163.367
R617 B.n479 B.n80 163.367
R618 B.n483 B.n80 163.367
R619 B.n484 B.n483 163.367
R620 B.n485 B.n484 163.367
R621 B.n485 B.n78 163.367
R622 B.n489 B.n78 163.367
R623 B.n490 B.n489 163.367
R624 B.n491 B.n490 163.367
R625 B.n491 B.n76 163.367
R626 B.n495 B.n76 163.367
R627 B.n496 B.n495 163.367
R628 B.n497 B.n496 163.367
R629 B.n497 B.n74 163.367
R630 B.n501 B.n74 163.367
R631 B.n502 B.n501 163.367
R632 B.n503 B.n502 163.367
R633 B.n503 B.n72 163.367
R634 B.n507 B.n72 163.367
R635 B.n508 B.n507 163.367
R636 B.n509 B.n508 163.367
R637 B.n509 B.n70 163.367
R638 B.n513 B.n70 163.367
R639 B.n514 B.n513 163.367
R640 B.n515 B.n514 163.367
R641 B.n515 B.n68 163.367
R642 B.n519 B.n68 163.367
R643 B.n520 B.n519 163.367
R644 B.n521 B.n520 163.367
R645 B.n521 B.n66 163.367
R646 B.n525 B.n66 163.367
R647 B.n526 B.n525 163.367
R648 B.n527 B.n526 163.367
R649 B.n527 B.n64 163.367
R650 B.n531 B.n64 163.367
R651 B.n612 B.n611 163.367
R652 B.n611 B.n610 163.367
R653 B.n610 B.n33 163.367
R654 B.n606 B.n33 163.367
R655 B.n606 B.n605 163.367
R656 B.n605 B.n604 163.367
R657 B.n604 B.n35 163.367
R658 B.n600 B.n35 163.367
R659 B.n600 B.n599 163.367
R660 B.n599 B.n598 163.367
R661 B.n598 B.n37 163.367
R662 B.n594 B.n37 163.367
R663 B.n594 B.n593 163.367
R664 B.n593 B.n592 163.367
R665 B.n592 B.n39 163.367
R666 B.n588 B.n39 163.367
R667 B.n588 B.n587 163.367
R668 B.n587 B.n586 163.367
R669 B.n586 B.n41 163.367
R670 B.n582 B.n41 163.367
R671 B.n582 B.n581 163.367
R672 B.n581 B.n580 163.367
R673 B.n580 B.n43 163.367
R674 B.n576 B.n43 163.367
R675 B.n576 B.n575 163.367
R676 B.n575 B.n574 163.367
R677 B.n574 B.n48 163.367
R678 B.n570 B.n48 163.367
R679 B.n570 B.n569 163.367
R680 B.n569 B.n568 163.367
R681 B.n568 B.n50 163.367
R682 B.n563 B.n50 163.367
R683 B.n563 B.n562 163.367
R684 B.n562 B.n561 163.367
R685 B.n561 B.n54 163.367
R686 B.n557 B.n54 163.367
R687 B.n557 B.n556 163.367
R688 B.n556 B.n555 163.367
R689 B.n555 B.n56 163.367
R690 B.n551 B.n56 163.367
R691 B.n551 B.n550 163.367
R692 B.n550 B.n549 163.367
R693 B.n549 B.n58 163.367
R694 B.n545 B.n58 163.367
R695 B.n545 B.n544 163.367
R696 B.n544 B.n543 163.367
R697 B.n543 B.n60 163.367
R698 B.n539 B.n60 163.367
R699 B.n539 B.n538 163.367
R700 B.n538 B.n537 163.367
R701 B.n537 B.n62 163.367
R702 B.n533 B.n62 163.367
R703 B.n533 B.n532 163.367
R704 B.n136 B.n135 66.9096
R705 B.n142 B.n141 66.9096
R706 B.n45 B.n44 66.9096
R707 B.n52 B.n51 66.9096
R708 B.n319 B.n136 59.5399
R709 B.n143 B.n142 59.5399
R710 B.n46 B.n45 59.5399
R711 B.n565 B.n52 59.5399
R712 B.n614 B.n613 29.8151
R713 B.n530 B.n63 29.8151
R714 B.n354 B.n123 29.8151
R715 B.n271 B.n270 29.8151
R716 B B.n703 18.0485
R717 B.n613 B.n32 10.6151
R718 B.n609 B.n32 10.6151
R719 B.n609 B.n608 10.6151
R720 B.n608 B.n607 10.6151
R721 B.n607 B.n34 10.6151
R722 B.n603 B.n34 10.6151
R723 B.n603 B.n602 10.6151
R724 B.n602 B.n601 10.6151
R725 B.n601 B.n36 10.6151
R726 B.n597 B.n36 10.6151
R727 B.n597 B.n596 10.6151
R728 B.n596 B.n595 10.6151
R729 B.n595 B.n38 10.6151
R730 B.n591 B.n38 10.6151
R731 B.n591 B.n590 10.6151
R732 B.n590 B.n589 10.6151
R733 B.n589 B.n40 10.6151
R734 B.n585 B.n40 10.6151
R735 B.n585 B.n584 10.6151
R736 B.n584 B.n583 10.6151
R737 B.n583 B.n42 10.6151
R738 B.n579 B.n578 10.6151
R739 B.n578 B.n577 10.6151
R740 B.n577 B.n47 10.6151
R741 B.n573 B.n47 10.6151
R742 B.n573 B.n572 10.6151
R743 B.n572 B.n571 10.6151
R744 B.n571 B.n49 10.6151
R745 B.n567 B.n49 10.6151
R746 B.n567 B.n566 10.6151
R747 B.n564 B.n53 10.6151
R748 B.n560 B.n53 10.6151
R749 B.n560 B.n559 10.6151
R750 B.n559 B.n558 10.6151
R751 B.n558 B.n55 10.6151
R752 B.n554 B.n55 10.6151
R753 B.n554 B.n553 10.6151
R754 B.n553 B.n552 10.6151
R755 B.n552 B.n57 10.6151
R756 B.n548 B.n57 10.6151
R757 B.n548 B.n547 10.6151
R758 B.n547 B.n546 10.6151
R759 B.n546 B.n59 10.6151
R760 B.n542 B.n59 10.6151
R761 B.n542 B.n541 10.6151
R762 B.n541 B.n540 10.6151
R763 B.n540 B.n61 10.6151
R764 B.n536 B.n61 10.6151
R765 B.n536 B.n535 10.6151
R766 B.n535 B.n534 10.6151
R767 B.n534 B.n63 10.6151
R768 B.n355 B.n354 10.6151
R769 B.n356 B.n355 10.6151
R770 B.n356 B.n121 10.6151
R771 B.n360 B.n121 10.6151
R772 B.n361 B.n360 10.6151
R773 B.n362 B.n361 10.6151
R774 B.n362 B.n119 10.6151
R775 B.n366 B.n119 10.6151
R776 B.n367 B.n366 10.6151
R777 B.n368 B.n367 10.6151
R778 B.n368 B.n117 10.6151
R779 B.n372 B.n117 10.6151
R780 B.n373 B.n372 10.6151
R781 B.n374 B.n373 10.6151
R782 B.n374 B.n115 10.6151
R783 B.n378 B.n115 10.6151
R784 B.n379 B.n378 10.6151
R785 B.n380 B.n379 10.6151
R786 B.n380 B.n113 10.6151
R787 B.n384 B.n113 10.6151
R788 B.n385 B.n384 10.6151
R789 B.n386 B.n385 10.6151
R790 B.n386 B.n111 10.6151
R791 B.n390 B.n111 10.6151
R792 B.n391 B.n390 10.6151
R793 B.n392 B.n391 10.6151
R794 B.n392 B.n109 10.6151
R795 B.n396 B.n109 10.6151
R796 B.n397 B.n396 10.6151
R797 B.n398 B.n397 10.6151
R798 B.n398 B.n107 10.6151
R799 B.n402 B.n107 10.6151
R800 B.n403 B.n402 10.6151
R801 B.n404 B.n403 10.6151
R802 B.n404 B.n105 10.6151
R803 B.n408 B.n105 10.6151
R804 B.n409 B.n408 10.6151
R805 B.n410 B.n409 10.6151
R806 B.n410 B.n103 10.6151
R807 B.n414 B.n103 10.6151
R808 B.n415 B.n414 10.6151
R809 B.n416 B.n415 10.6151
R810 B.n416 B.n101 10.6151
R811 B.n420 B.n101 10.6151
R812 B.n421 B.n420 10.6151
R813 B.n422 B.n421 10.6151
R814 B.n422 B.n99 10.6151
R815 B.n426 B.n99 10.6151
R816 B.n427 B.n426 10.6151
R817 B.n428 B.n427 10.6151
R818 B.n428 B.n97 10.6151
R819 B.n432 B.n97 10.6151
R820 B.n433 B.n432 10.6151
R821 B.n434 B.n433 10.6151
R822 B.n434 B.n95 10.6151
R823 B.n438 B.n95 10.6151
R824 B.n439 B.n438 10.6151
R825 B.n440 B.n439 10.6151
R826 B.n440 B.n93 10.6151
R827 B.n444 B.n93 10.6151
R828 B.n445 B.n444 10.6151
R829 B.n446 B.n445 10.6151
R830 B.n446 B.n91 10.6151
R831 B.n450 B.n91 10.6151
R832 B.n451 B.n450 10.6151
R833 B.n452 B.n451 10.6151
R834 B.n452 B.n89 10.6151
R835 B.n456 B.n89 10.6151
R836 B.n457 B.n456 10.6151
R837 B.n458 B.n457 10.6151
R838 B.n458 B.n87 10.6151
R839 B.n462 B.n87 10.6151
R840 B.n463 B.n462 10.6151
R841 B.n464 B.n463 10.6151
R842 B.n464 B.n85 10.6151
R843 B.n468 B.n85 10.6151
R844 B.n469 B.n468 10.6151
R845 B.n470 B.n469 10.6151
R846 B.n470 B.n83 10.6151
R847 B.n474 B.n83 10.6151
R848 B.n475 B.n474 10.6151
R849 B.n476 B.n475 10.6151
R850 B.n476 B.n81 10.6151
R851 B.n480 B.n81 10.6151
R852 B.n481 B.n480 10.6151
R853 B.n482 B.n481 10.6151
R854 B.n482 B.n79 10.6151
R855 B.n486 B.n79 10.6151
R856 B.n487 B.n486 10.6151
R857 B.n488 B.n487 10.6151
R858 B.n488 B.n77 10.6151
R859 B.n492 B.n77 10.6151
R860 B.n493 B.n492 10.6151
R861 B.n494 B.n493 10.6151
R862 B.n494 B.n75 10.6151
R863 B.n498 B.n75 10.6151
R864 B.n499 B.n498 10.6151
R865 B.n500 B.n499 10.6151
R866 B.n500 B.n73 10.6151
R867 B.n504 B.n73 10.6151
R868 B.n505 B.n504 10.6151
R869 B.n506 B.n505 10.6151
R870 B.n506 B.n71 10.6151
R871 B.n510 B.n71 10.6151
R872 B.n511 B.n510 10.6151
R873 B.n512 B.n511 10.6151
R874 B.n512 B.n69 10.6151
R875 B.n516 B.n69 10.6151
R876 B.n517 B.n516 10.6151
R877 B.n518 B.n517 10.6151
R878 B.n518 B.n67 10.6151
R879 B.n522 B.n67 10.6151
R880 B.n523 B.n522 10.6151
R881 B.n524 B.n523 10.6151
R882 B.n524 B.n65 10.6151
R883 B.n528 B.n65 10.6151
R884 B.n529 B.n528 10.6151
R885 B.n530 B.n529 10.6151
R886 B.n272 B.n271 10.6151
R887 B.n272 B.n153 10.6151
R888 B.n276 B.n153 10.6151
R889 B.n277 B.n276 10.6151
R890 B.n278 B.n277 10.6151
R891 B.n278 B.n151 10.6151
R892 B.n282 B.n151 10.6151
R893 B.n283 B.n282 10.6151
R894 B.n284 B.n283 10.6151
R895 B.n284 B.n149 10.6151
R896 B.n288 B.n149 10.6151
R897 B.n289 B.n288 10.6151
R898 B.n290 B.n289 10.6151
R899 B.n290 B.n147 10.6151
R900 B.n294 B.n147 10.6151
R901 B.n295 B.n294 10.6151
R902 B.n296 B.n295 10.6151
R903 B.n296 B.n145 10.6151
R904 B.n300 B.n145 10.6151
R905 B.n301 B.n300 10.6151
R906 B.n302 B.n301 10.6151
R907 B.n306 B.n305 10.6151
R908 B.n307 B.n306 10.6151
R909 B.n307 B.n139 10.6151
R910 B.n311 B.n139 10.6151
R911 B.n312 B.n311 10.6151
R912 B.n313 B.n312 10.6151
R913 B.n313 B.n137 10.6151
R914 B.n317 B.n137 10.6151
R915 B.n318 B.n317 10.6151
R916 B.n320 B.n133 10.6151
R917 B.n324 B.n133 10.6151
R918 B.n325 B.n324 10.6151
R919 B.n326 B.n325 10.6151
R920 B.n326 B.n131 10.6151
R921 B.n330 B.n131 10.6151
R922 B.n331 B.n330 10.6151
R923 B.n332 B.n331 10.6151
R924 B.n332 B.n129 10.6151
R925 B.n336 B.n129 10.6151
R926 B.n337 B.n336 10.6151
R927 B.n338 B.n337 10.6151
R928 B.n338 B.n127 10.6151
R929 B.n342 B.n127 10.6151
R930 B.n343 B.n342 10.6151
R931 B.n344 B.n343 10.6151
R932 B.n344 B.n125 10.6151
R933 B.n348 B.n125 10.6151
R934 B.n349 B.n348 10.6151
R935 B.n350 B.n349 10.6151
R936 B.n350 B.n123 10.6151
R937 B.n270 B.n155 10.6151
R938 B.n266 B.n155 10.6151
R939 B.n266 B.n265 10.6151
R940 B.n265 B.n264 10.6151
R941 B.n264 B.n157 10.6151
R942 B.n260 B.n157 10.6151
R943 B.n260 B.n259 10.6151
R944 B.n259 B.n258 10.6151
R945 B.n258 B.n159 10.6151
R946 B.n254 B.n159 10.6151
R947 B.n254 B.n253 10.6151
R948 B.n253 B.n252 10.6151
R949 B.n252 B.n161 10.6151
R950 B.n248 B.n161 10.6151
R951 B.n248 B.n247 10.6151
R952 B.n247 B.n246 10.6151
R953 B.n246 B.n163 10.6151
R954 B.n242 B.n163 10.6151
R955 B.n242 B.n241 10.6151
R956 B.n241 B.n240 10.6151
R957 B.n240 B.n165 10.6151
R958 B.n236 B.n165 10.6151
R959 B.n236 B.n235 10.6151
R960 B.n235 B.n234 10.6151
R961 B.n234 B.n167 10.6151
R962 B.n230 B.n167 10.6151
R963 B.n230 B.n229 10.6151
R964 B.n229 B.n228 10.6151
R965 B.n228 B.n169 10.6151
R966 B.n224 B.n169 10.6151
R967 B.n224 B.n223 10.6151
R968 B.n223 B.n222 10.6151
R969 B.n222 B.n171 10.6151
R970 B.n218 B.n171 10.6151
R971 B.n218 B.n217 10.6151
R972 B.n217 B.n216 10.6151
R973 B.n216 B.n173 10.6151
R974 B.n212 B.n173 10.6151
R975 B.n212 B.n211 10.6151
R976 B.n211 B.n210 10.6151
R977 B.n210 B.n175 10.6151
R978 B.n206 B.n175 10.6151
R979 B.n206 B.n205 10.6151
R980 B.n205 B.n204 10.6151
R981 B.n204 B.n177 10.6151
R982 B.n200 B.n177 10.6151
R983 B.n200 B.n199 10.6151
R984 B.n199 B.n198 10.6151
R985 B.n198 B.n179 10.6151
R986 B.n194 B.n179 10.6151
R987 B.n194 B.n193 10.6151
R988 B.n193 B.n192 10.6151
R989 B.n192 B.n181 10.6151
R990 B.n188 B.n181 10.6151
R991 B.n188 B.n187 10.6151
R992 B.n187 B.n186 10.6151
R993 B.n186 B.n183 10.6151
R994 B.n183 B.n0 10.6151
R995 B.n699 B.n1 10.6151
R996 B.n699 B.n698 10.6151
R997 B.n698 B.n697 10.6151
R998 B.n697 B.n4 10.6151
R999 B.n693 B.n4 10.6151
R1000 B.n693 B.n692 10.6151
R1001 B.n692 B.n691 10.6151
R1002 B.n691 B.n6 10.6151
R1003 B.n687 B.n6 10.6151
R1004 B.n687 B.n686 10.6151
R1005 B.n686 B.n685 10.6151
R1006 B.n685 B.n8 10.6151
R1007 B.n681 B.n8 10.6151
R1008 B.n681 B.n680 10.6151
R1009 B.n680 B.n679 10.6151
R1010 B.n679 B.n10 10.6151
R1011 B.n675 B.n10 10.6151
R1012 B.n675 B.n674 10.6151
R1013 B.n674 B.n673 10.6151
R1014 B.n673 B.n12 10.6151
R1015 B.n669 B.n12 10.6151
R1016 B.n669 B.n668 10.6151
R1017 B.n668 B.n667 10.6151
R1018 B.n667 B.n14 10.6151
R1019 B.n663 B.n14 10.6151
R1020 B.n663 B.n662 10.6151
R1021 B.n662 B.n661 10.6151
R1022 B.n661 B.n16 10.6151
R1023 B.n657 B.n16 10.6151
R1024 B.n657 B.n656 10.6151
R1025 B.n656 B.n655 10.6151
R1026 B.n655 B.n18 10.6151
R1027 B.n651 B.n18 10.6151
R1028 B.n651 B.n650 10.6151
R1029 B.n650 B.n649 10.6151
R1030 B.n649 B.n20 10.6151
R1031 B.n645 B.n20 10.6151
R1032 B.n645 B.n644 10.6151
R1033 B.n644 B.n643 10.6151
R1034 B.n643 B.n22 10.6151
R1035 B.n639 B.n22 10.6151
R1036 B.n639 B.n638 10.6151
R1037 B.n638 B.n637 10.6151
R1038 B.n637 B.n24 10.6151
R1039 B.n633 B.n24 10.6151
R1040 B.n633 B.n632 10.6151
R1041 B.n632 B.n631 10.6151
R1042 B.n631 B.n26 10.6151
R1043 B.n627 B.n26 10.6151
R1044 B.n627 B.n626 10.6151
R1045 B.n626 B.n625 10.6151
R1046 B.n625 B.n28 10.6151
R1047 B.n621 B.n28 10.6151
R1048 B.n621 B.n620 10.6151
R1049 B.n620 B.n619 10.6151
R1050 B.n619 B.n30 10.6151
R1051 B.n615 B.n30 10.6151
R1052 B.n615 B.n614 10.6151
R1053 B.n46 B.n42 9.36635
R1054 B.n565 B.n564 9.36635
R1055 B.n302 B.n143 9.36635
R1056 B.n320 B.n319 9.36635
R1057 B.n703 B.n0 2.81026
R1058 B.n703 B.n1 2.81026
R1059 B.n579 B.n46 1.24928
R1060 B.n566 B.n565 1.24928
R1061 B.n305 B.n143 1.24928
R1062 B.n319 B.n318 1.24928
R1063 VP.n21 VP.n18 161.3
R1064 VP.n23 VP.n22 161.3
R1065 VP.n24 VP.n17 161.3
R1066 VP.n26 VP.n25 161.3
R1067 VP.n27 VP.n16 161.3
R1068 VP.n29 VP.n28 161.3
R1069 VP.n31 VP.n30 161.3
R1070 VP.n32 VP.n14 161.3
R1071 VP.n34 VP.n33 161.3
R1072 VP.n35 VP.n13 161.3
R1073 VP.n37 VP.n36 161.3
R1074 VP.n38 VP.n12 161.3
R1075 VP.n40 VP.n39 161.3
R1076 VP.n75 VP.n74 161.3
R1077 VP.n73 VP.n1 161.3
R1078 VP.n72 VP.n71 161.3
R1079 VP.n70 VP.n2 161.3
R1080 VP.n69 VP.n68 161.3
R1081 VP.n67 VP.n3 161.3
R1082 VP.n66 VP.n65 161.3
R1083 VP.n64 VP.n63 161.3
R1084 VP.n62 VP.n5 161.3
R1085 VP.n61 VP.n60 161.3
R1086 VP.n59 VP.n6 161.3
R1087 VP.n58 VP.n57 161.3
R1088 VP.n56 VP.n7 161.3
R1089 VP.n54 VP.n53 161.3
R1090 VP.n52 VP.n8 161.3
R1091 VP.n51 VP.n50 161.3
R1092 VP.n49 VP.n9 161.3
R1093 VP.n48 VP.n47 161.3
R1094 VP.n46 VP.n10 161.3
R1095 VP.n45 VP.n44 161.3
R1096 VP.n19 VP.t3 74.8933
R1097 VP.n43 VP.n42 69.2705
R1098 VP.n76 VP.n0 69.2705
R1099 VP.n41 VP.n11 69.2705
R1100 VP.n49 VP.n48 56.5193
R1101 VP.n61 VP.n6 56.5193
R1102 VP.n72 VP.n2 56.5193
R1103 VP.n37 VP.n13 56.5193
R1104 VP.n26 VP.n17 56.5193
R1105 VP.n20 VP.n19 50.6608
R1106 VP.n42 VP.n41 48.469
R1107 VP.n43 VP.t4 41.4803
R1108 VP.n55 VP.t1 41.4803
R1109 VP.n4 VP.t6 41.4803
R1110 VP.n0 VP.t0 41.4803
R1111 VP.n11 VP.t7 41.4803
R1112 VP.n15 VP.t2 41.4803
R1113 VP.n20 VP.t5 41.4803
R1114 VP.n44 VP.n10 24.4675
R1115 VP.n48 VP.n10 24.4675
R1116 VP.n50 VP.n49 24.4675
R1117 VP.n50 VP.n8 24.4675
R1118 VP.n54 VP.n8 24.4675
R1119 VP.n57 VP.n56 24.4675
R1120 VP.n57 VP.n6 24.4675
R1121 VP.n62 VP.n61 24.4675
R1122 VP.n63 VP.n62 24.4675
R1123 VP.n67 VP.n66 24.4675
R1124 VP.n68 VP.n67 24.4675
R1125 VP.n68 VP.n2 24.4675
R1126 VP.n73 VP.n72 24.4675
R1127 VP.n74 VP.n73 24.4675
R1128 VP.n38 VP.n37 24.4675
R1129 VP.n39 VP.n38 24.4675
R1130 VP.n27 VP.n26 24.4675
R1131 VP.n28 VP.n27 24.4675
R1132 VP.n32 VP.n31 24.4675
R1133 VP.n33 VP.n32 24.4675
R1134 VP.n33 VP.n13 24.4675
R1135 VP.n22 VP.n21 24.4675
R1136 VP.n22 VP.n17 24.4675
R1137 VP.n56 VP.n55 23.2442
R1138 VP.n63 VP.n4 23.2442
R1139 VP.n28 VP.n15 23.2442
R1140 VP.n21 VP.n20 23.2442
R1141 VP.n44 VP.n43 20.7975
R1142 VP.n74 VP.n0 20.7975
R1143 VP.n39 VP.n11 20.7975
R1144 VP.n19 VP.n18 3.87631
R1145 VP.n55 VP.n54 1.22385
R1146 VP.n66 VP.n4 1.22385
R1147 VP.n31 VP.n15 1.22385
R1148 VP.n41 VP.n40 0.354971
R1149 VP.n45 VP.n42 0.354971
R1150 VP.n76 VP.n75 0.354971
R1151 VP VP.n76 0.26696
R1152 VP.n23 VP.n18 0.189894
R1153 VP.n24 VP.n23 0.189894
R1154 VP.n25 VP.n24 0.189894
R1155 VP.n25 VP.n16 0.189894
R1156 VP.n29 VP.n16 0.189894
R1157 VP.n30 VP.n29 0.189894
R1158 VP.n30 VP.n14 0.189894
R1159 VP.n34 VP.n14 0.189894
R1160 VP.n35 VP.n34 0.189894
R1161 VP.n36 VP.n35 0.189894
R1162 VP.n36 VP.n12 0.189894
R1163 VP.n40 VP.n12 0.189894
R1164 VP.n46 VP.n45 0.189894
R1165 VP.n47 VP.n46 0.189894
R1166 VP.n47 VP.n9 0.189894
R1167 VP.n51 VP.n9 0.189894
R1168 VP.n52 VP.n51 0.189894
R1169 VP.n53 VP.n52 0.189894
R1170 VP.n53 VP.n7 0.189894
R1171 VP.n58 VP.n7 0.189894
R1172 VP.n59 VP.n58 0.189894
R1173 VP.n60 VP.n59 0.189894
R1174 VP.n60 VP.n5 0.189894
R1175 VP.n64 VP.n5 0.189894
R1176 VP.n65 VP.n64 0.189894
R1177 VP.n65 VP.n3 0.189894
R1178 VP.n69 VP.n3 0.189894
R1179 VP.n70 VP.n69 0.189894
R1180 VP.n71 VP.n70 0.189894
R1181 VP.n71 VP.n1 0.189894
R1182 VP.n75 VP.n1 0.189894
R1183 VTAIL.n226 VTAIL.n204 756.745
R1184 VTAIL.n24 VTAIL.n2 756.745
R1185 VTAIL.n52 VTAIL.n30 756.745
R1186 VTAIL.n82 VTAIL.n60 756.745
R1187 VTAIL.n198 VTAIL.n176 756.745
R1188 VTAIL.n168 VTAIL.n146 756.745
R1189 VTAIL.n140 VTAIL.n118 756.745
R1190 VTAIL.n110 VTAIL.n88 756.745
R1191 VTAIL.n212 VTAIL.n211 585
R1192 VTAIL.n217 VTAIL.n216 585
R1193 VTAIL.n219 VTAIL.n218 585
R1194 VTAIL.n208 VTAIL.n207 585
R1195 VTAIL.n225 VTAIL.n224 585
R1196 VTAIL.n227 VTAIL.n226 585
R1197 VTAIL.n10 VTAIL.n9 585
R1198 VTAIL.n15 VTAIL.n14 585
R1199 VTAIL.n17 VTAIL.n16 585
R1200 VTAIL.n6 VTAIL.n5 585
R1201 VTAIL.n23 VTAIL.n22 585
R1202 VTAIL.n25 VTAIL.n24 585
R1203 VTAIL.n38 VTAIL.n37 585
R1204 VTAIL.n43 VTAIL.n42 585
R1205 VTAIL.n45 VTAIL.n44 585
R1206 VTAIL.n34 VTAIL.n33 585
R1207 VTAIL.n51 VTAIL.n50 585
R1208 VTAIL.n53 VTAIL.n52 585
R1209 VTAIL.n68 VTAIL.n67 585
R1210 VTAIL.n73 VTAIL.n72 585
R1211 VTAIL.n75 VTAIL.n74 585
R1212 VTAIL.n64 VTAIL.n63 585
R1213 VTAIL.n81 VTAIL.n80 585
R1214 VTAIL.n83 VTAIL.n82 585
R1215 VTAIL.n199 VTAIL.n198 585
R1216 VTAIL.n197 VTAIL.n196 585
R1217 VTAIL.n180 VTAIL.n179 585
R1218 VTAIL.n191 VTAIL.n190 585
R1219 VTAIL.n189 VTAIL.n188 585
R1220 VTAIL.n184 VTAIL.n183 585
R1221 VTAIL.n169 VTAIL.n168 585
R1222 VTAIL.n167 VTAIL.n166 585
R1223 VTAIL.n150 VTAIL.n149 585
R1224 VTAIL.n161 VTAIL.n160 585
R1225 VTAIL.n159 VTAIL.n158 585
R1226 VTAIL.n154 VTAIL.n153 585
R1227 VTAIL.n141 VTAIL.n140 585
R1228 VTAIL.n139 VTAIL.n138 585
R1229 VTAIL.n122 VTAIL.n121 585
R1230 VTAIL.n133 VTAIL.n132 585
R1231 VTAIL.n131 VTAIL.n130 585
R1232 VTAIL.n126 VTAIL.n125 585
R1233 VTAIL.n111 VTAIL.n110 585
R1234 VTAIL.n109 VTAIL.n108 585
R1235 VTAIL.n92 VTAIL.n91 585
R1236 VTAIL.n103 VTAIL.n102 585
R1237 VTAIL.n101 VTAIL.n100 585
R1238 VTAIL.n96 VTAIL.n95 585
R1239 VTAIL.n213 VTAIL.t1 327.856
R1240 VTAIL.n11 VTAIL.t7 327.856
R1241 VTAIL.n39 VTAIL.t9 327.856
R1242 VTAIL.n69 VTAIL.t13 327.856
R1243 VTAIL.n185 VTAIL.t11 327.856
R1244 VTAIL.n155 VTAIL.t15 327.856
R1245 VTAIL.n127 VTAIL.t2 327.856
R1246 VTAIL.n97 VTAIL.t6 327.856
R1247 VTAIL.n217 VTAIL.n211 171.744
R1248 VTAIL.n218 VTAIL.n217 171.744
R1249 VTAIL.n218 VTAIL.n207 171.744
R1250 VTAIL.n225 VTAIL.n207 171.744
R1251 VTAIL.n226 VTAIL.n225 171.744
R1252 VTAIL.n15 VTAIL.n9 171.744
R1253 VTAIL.n16 VTAIL.n15 171.744
R1254 VTAIL.n16 VTAIL.n5 171.744
R1255 VTAIL.n23 VTAIL.n5 171.744
R1256 VTAIL.n24 VTAIL.n23 171.744
R1257 VTAIL.n43 VTAIL.n37 171.744
R1258 VTAIL.n44 VTAIL.n43 171.744
R1259 VTAIL.n44 VTAIL.n33 171.744
R1260 VTAIL.n51 VTAIL.n33 171.744
R1261 VTAIL.n52 VTAIL.n51 171.744
R1262 VTAIL.n73 VTAIL.n67 171.744
R1263 VTAIL.n74 VTAIL.n73 171.744
R1264 VTAIL.n74 VTAIL.n63 171.744
R1265 VTAIL.n81 VTAIL.n63 171.744
R1266 VTAIL.n82 VTAIL.n81 171.744
R1267 VTAIL.n198 VTAIL.n197 171.744
R1268 VTAIL.n197 VTAIL.n179 171.744
R1269 VTAIL.n190 VTAIL.n179 171.744
R1270 VTAIL.n190 VTAIL.n189 171.744
R1271 VTAIL.n189 VTAIL.n183 171.744
R1272 VTAIL.n168 VTAIL.n167 171.744
R1273 VTAIL.n167 VTAIL.n149 171.744
R1274 VTAIL.n160 VTAIL.n149 171.744
R1275 VTAIL.n160 VTAIL.n159 171.744
R1276 VTAIL.n159 VTAIL.n153 171.744
R1277 VTAIL.n140 VTAIL.n139 171.744
R1278 VTAIL.n139 VTAIL.n121 171.744
R1279 VTAIL.n132 VTAIL.n121 171.744
R1280 VTAIL.n132 VTAIL.n131 171.744
R1281 VTAIL.n131 VTAIL.n125 171.744
R1282 VTAIL.n110 VTAIL.n109 171.744
R1283 VTAIL.n109 VTAIL.n91 171.744
R1284 VTAIL.n102 VTAIL.n91 171.744
R1285 VTAIL.n102 VTAIL.n101 171.744
R1286 VTAIL.n101 VTAIL.n95 171.744
R1287 VTAIL.t1 VTAIL.n211 85.8723
R1288 VTAIL.t7 VTAIL.n9 85.8723
R1289 VTAIL.t9 VTAIL.n37 85.8723
R1290 VTAIL.t13 VTAIL.n67 85.8723
R1291 VTAIL.t11 VTAIL.n183 85.8723
R1292 VTAIL.t15 VTAIL.n153 85.8723
R1293 VTAIL.t2 VTAIL.n125 85.8723
R1294 VTAIL.t6 VTAIL.n95 85.8723
R1295 VTAIL.n175 VTAIL.n174 82.3976
R1296 VTAIL.n117 VTAIL.n116 82.3976
R1297 VTAIL.n1 VTAIL.n0 82.3974
R1298 VTAIL.n59 VTAIL.n58 82.3974
R1299 VTAIL.n231 VTAIL.n230 33.9308
R1300 VTAIL.n29 VTAIL.n28 33.9308
R1301 VTAIL.n57 VTAIL.n56 33.9308
R1302 VTAIL.n87 VTAIL.n86 33.9308
R1303 VTAIL.n203 VTAIL.n202 33.9308
R1304 VTAIL.n173 VTAIL.n172 33.9308
R1305 VTAIL.n145 VTAIL.n144 33.9308
R1306 VTAIL.n115 VTAIL.n114 33.9308
R1307 VTAIL.n231 VTAIL.n203 19.9703
R1308 VTAIL.n115 VTAIL.n87 19.9703
R1309 VTAIL.n213 VTAIL.n212 16.381
R1310 VTAIL.n11 VTAIL.n10 16.381
R1311 VTAIL.n39 VTAIL.n38 16.381
R1312 VTAIL.n69 VTAIL.n68 16.381
R1313 VTAIL.n185 VTAIL.n184 16.381
R1314 VTAIL.n155 VTAIL.n154 16.381
R1315 VTAIL.n127 VTAIL.n126 16.381
R1316 VTAIL.n97 VTAIL.n96 16.381
R1317 VTAIL.n216 VTAIL.n215 12.8005
R1318 VTAIL.n14 VTAIL.n13 12.8005
R1319 VTAIL.n42 VTAIL.n41 12.8005
R1320 VTAIL.n72 VTAIL.n71 12.8005
R1321 VTAIL.n188 VTAIL.n187 12.8005
R1322 VTAIL.n158 VTAIL.n157 12.8005
R1323 VTAIL.n130 VTAIL.n129 12.8005
R1324 VTAIL.n100 VTAIL.n99 12.8005
R1325 VTAIL.n219 VTAIL.n210 12.0247
R1326 VTAIL.n17 VTAIL.n8 12.0247
R1327 VTAIL.n45 VTAIL.n36 12.0247
R1328 VTAIL.n75 VTAIL.n66 12.0247
R1329 VTAIL.n191 VTAIL.n182 12.0247
R1330 VTAIL.n161 VTAIL.n152 12.0247
R1331 VTAIL.n133 VTAIL.n124 12.0247
R1332 VTAIL.n103 VTAIL.n94 12.0247
R1333 VTAIL.n220 VTAIL.n208 11.249
R1334 VTAIL.n18 VTAIL.n6 11.249
R1335 VTAIL.n46 VTAIL.n34 11.249
R1336 VTAIL.n76 VTAIL.n64 11.249
R1337 VTAIL.n192 VTAIL.n180 11.249
R1338 VTAIL.n162 VTAIL.n150 11.249
R1339 VTAIL.n134 VTAIL.n122 11.249
R1340 VTAIL.n104 VTAIL.n92 11.249
R1341 VTAIL.n224 VTAIL.n223 10.4732
R1342 VTAIL.n22 VTAIL.n21 10.4732
R1343 VTAIL.n50 VTAIL.n49 10.4732
R1344 VTAIL.n80 VTAIL.n79 10.4732
R1345 VTAIL.n196 VTAIL.n195 10.4732
R1346 VTAIL.n166 VTAIL.n165 10.4732
R1347 VTAIL.n138 VTAIL.n137 10.4732
R1348 VTAIL.n108 VTAIL.n107 10.4732
R1349 VTAIL.n227 VTAIL.n206 9.69747
R1350 VTAIL.n25 VTAIL.n4 9.69747
R1351 VTAIL.n53 VTAIL.n32 9.69747
R1352 VTAIL.n83 VTAIL.n62 9.69747
R1353 VTAIL.n199 VTAIL.n178 9.69747
R1354 VTAIL.n169 VTAIL.n148 9.69747
R1355 VTAIL.n141 VTAIL.n120 9.69747
R1356 VTAIL.n111 VTAIL.n90 9.69747
R1357 VTAIL.n230 VTAIL.n229 9.45567
R1358 VTAIL.n28 VTAIL.n27 9.45567
R1359 VTAIL.n56 VTAIL.n55 9.45567
R1360 VTAIL.n86 VTAIL.n85 9.45567
R1361 VTAIL.n202 VTAIL.n201 9.45567
R1362 VTAIL.n172 VTAIL.n171 9.45567
R1363 VTAIL.n144 VTAIL.n143 9.45567
R1364 VTAIL.n114 VTAIL.n113 9.45567
R1365 VTAIL.n229 VTAIL.n228 9.3005
R1366 VTAIL.n206 VTAIL.n205 9.3005
R1367 VTAIL.n223 VTAIL.n222 9.3005
R1368 VTAIL.n221 VTAIL.n220 9.3005
R1369 VTAIL.n210 VTAIL.n209 9.3005
R1370 VTAIL.n215 VTAIL.n214 9.3005
R1371 VTAIL.n27 VTAIL.n26 9.3005
R1372 VTAIL.n4 VTAIL.n3 9.3005
R1373 VTAIL.n21 VTAIL.n20 9.3005
R1374 VTAIL.n19 VTAIL.n18 9.3005
R1375 VTAIL.n8 VTAIL.n7 9.3005
R1376 VTAIL.n13 VTAIL.n12 9.3005
R1377 VTAIL.n55 VTAIL.n54 9.3005
R1378 VTAIL.n32 VTAIL.n31 9.3005
R1379 VTAIL.n49 VTAIL.n48 9.3005
R1380 VTAIL.n47 VTAIL.n46 9.3005
R1381 VTAIL.n36 VTAIL.n35 9.3005
R1382 VTAIL.n41 VTAIL.n40 9.3005
R1383 VTAIL.n85 VTAIL.n84 9.3005
R1384 VTAIL.n62 VTAIL.n61 9.3005
R1385 VTAIL.n79 VTAIL.n78 9.3005
R1386 VTAIL.n77 VTAIL.n76 9.3005
R1387 VTAIL.n66 VTAIL.n65 9.3005
R1388 VTAIL.n71 VTAIL.n70 9.3005
R1389 VTAIL.n201 VTAIL.n200 9.3005
R1390 VTAIL.n178 VTAIL.n177 9.3005
R1391 VTAIL.n195 VTAIL.n194 9.3005
R1392 VTAIL.n193 VTAIL.n192 9.3005
R1393 VTAIL.n182 VTAIL.n181 9.3005
R1394 VTAIL.n187 VTAIL.n186 9.3005
R1395 VTAIL.n171 VTAIL.n170 9.3005
R1396 VTAIL.n148 VTAIL.n147 9.3005
R1397 VTAIL.n165 VTAIL.n164 9.3005
R1398 VTAIL.n163 VTAIL.n162 9.3005
R1399 VTAIL.n152 VTAIL.n151 9.3005
R1400 VTAIL.n157 VTAIL.n156 9.3005
R1401 VTAIL.n143 VTAIL.n142 9.3005
R1402 VTAIL.n120 VTAIL.n119 9.3005
R1403 VTAIL.n137 VTAIL.n136 9.3005
R1404 VTAIL.n135 VTAIL.n134 9.3005
R1405 VTAIL.n124 VTAIL.n123 9.3005
R1406 VTAIL.n129 VTAIL.n128 9.3005
R1407 VTAIL.n113 VTAIL.n112 9.3005
R1408 VTAIL.n90 VTAIL.n89 9.3005
R1409 VTAIL.n107 VTAIL.n106 9.3005
R1410 VTAIL.n105 VTAIL.n104 9.3005
R1411 VTAIL.n94 VTAIL.n93 9.3005
R1412 VTAIL.n99 VTAIL.n98 9.3005
R1413 VTAIL.n228 VTAIL.n204 8.92171
R1414 VTAIL.n26 VTAIL.n2 8.92171
R1415 VTAIL.n54 VTAIL.n30 8.92171
R1416 VTAIL.n84 VTAIL.n60 8.92171
R1417 VTAIL.n200 VTAIL.n176 8.92171
R1418 VTAIL.n170 VTAIL.n146 8.92171
R1419 VTAIL.n142 VTAIL.n118 8.92171
R1420 VTAIL.n112 VTAIL.n88 8.92171
R1421 VTAIL.n0 VTAIL.t5 6.05357
R1422 VTAIL.n0 VTAIL.t4 6.05357
R1423 VTAIL.n58 VTAIL.t12 6.05357
R1424 VTAIL.n58 VTAIL.t8 6.05357
R1425 VTAIL.n174 VTAIL.t14 6.05357
R1426 VTAIL.n174 VTAIL.t10 6.05357
R1427 VTAIL.n116 VTAIL.t0 6.05357
R1428 VTAIL.n116 VTAIL.t3 6.05357
R1429 VTAIL.n230 VTAIL.n204 5.04292
R1430 VTAIL.n28 VTAIL.n2 5.04292
R1431 VTAIL.n56 VTAIL.n30 5.04292
R1432 VTAIL.n86 VTAIL.n60 5.04292
R1433 VTAIL.n202 VTAIL.n176 5.04292
R1434 VTAIL.n172 VTAIL.n146 5.04292
R1435 VTAIL.n144 VTAIL.n118 5.04292
R1436 VTAIL.n114 VTAIL.n88 5.04292
R1437 VTAIL.n228 VTAIL.n227 4.26717
R1438 VTAIL.n26 VTAIL.n25 4.26717
R1439 VTAIL.n54 VTAIL.n53 4.26717
R1440 VTAIL.n84 VTAIL.n83 4.26717
R1441 VTAIL.n200 VTAIL.n199 4.26717
R1442 VTAIL.n170 VTAIL.n169 4.26717
R1443 VTAIL.n142 VTAIL.n141 4.26717
R1444 VTAIL.n112 VTAIL.n111 4.26717
R1445 VTAIL.n186 VTAIL.n185 3.71853
R1446 VTAIL.n156 VTAIL.n155 3.71853
R1447 VTAIL.n128 VTAIL.n127 3.71853
R1448 VTAIL.n98 VTAIL.n97 3.71853
R1449 VTAIL.n214 VTAIL.n213 3.71853
R1450 VTAIL.n12 VTAIL.n11 3.71853
R1451 VTAIL.n40 VTAIL.n39 3.71853
R1452 VTAIL.n70 VTAIL.n69 3.71853
R1453 VTAIL.n224 VTAIL.n206 3.49141
R1454 VTAIL.n22 VTAIL.n4 3.49141
R1455 VTAIL.n50 VTAIL.n32 3.49141
R1456 VTAIL.n80 VTAIL.n62 3.49141
R1457 VTAIL.n196 VTAIL.n178 3.49141
R1458 VTAIL.n166 VTAIL.n148 3.49141
R1459 VTAIL.n138 VTAIL.n120 3.49141
R1460 VTAIL.n108 VTAIL.n90 3.49141
R1461 VTAIL.n117 VTAIL.n115 2.97464
R1462 VTAIL.n145 VTAIL.n117 2.97464
R1463 VTAIL.n175 VTAIL.n173 2.97464
R1464 VTAIL.n203 VTAIL.n175 2.97464
R1465 VTAIL.n87 VTAIL.n59 2.97464
R1466 VTAIL.n59 VTAIL.n57 2.97464
R1467 VTAIL.n29 VTAIL.n1 2.97464
R1468 VTAIL VTAIL.n231 2.91645
R1469 VTAIL.n223 VTAIL.n208 2.71565
R1470 VTAIL.n21 VTAIL.n6 2.71565
R1471 VTAIL.n49 VTAIL.n34 2.71565
R1472 VTAIL.n79 VTAIL.n64 2.71565
R1473 VTAIL.n195 VTAIL.n180 2.71565
R1474 VTAIL.n165 VTAIL.n150 2.71565
R1475 VTAIL.n137 VTAIL.n122 2.71565
R1476 VTAIL.n107 VTAIL.n92 2.71565
R1477 VTAIL.n220 VTAIL.n219 1.93989
R1478 VTAIL.n18 VTAIL.n17 1.93989
R1479 VTAIL.n46 VTAIL.n45 1.93989
R1480 VTAIL.n76 VTAIL.n75 1.93989
R1481 VTAIL.n192 VTAIL.n191 1.93989
R1482 VTAIL.n162 VTAIL.n161 1.93989
R1483 VTAIL.n134 VTAIL.n133 1.93989
R1484 VTAIL.n104 VTAIL.n103 1.93989
R1485 VTAIL.n216 VTAIL.n210 1.16414
R1486 VTAIL.n14 VTAIL.n8 1.16414
R1487 VTAIL.n42 VTAIL.n36 1.16414
R1488 VTAIL.n72 VTAIL.n66 1.16414
R1489 VTAIL.n188 VTAIL.n182 1.16414
R1490 VTAIL.n158 VTAIL.n152 1.16414
R1491 VTAIL.n130 VTAIL.n124 1.16414
R1492 VTAIL.n100 VTAIL.n94 1.16414
R1493 VTAIL.n173 VTAIL.n145 0.470328
R1494 VTAIL.n57 VTAIL.n29 0.470328
R1495 VTAIL.n215 VTAIL.n212 0.388379
R1496 VTAIL.n13 VTAIL.n10 0.388379
R1497 VTAIL.n41 VTAIL.n38 0.388379
R1498 VTAIL.n71 VTAIL.n68 0.388379
R1499 VTAIL.n187 VTAIL.n184 0.388379
R1500 VTAIL.n157 VTAIL.n154 0.388379
R1501 VTAIL.n129 VTAIL.n126 0.388379
R1502 VTAIL.n99 VTAIL.n96 0.388379
R1503 VTAIL.n214 VTAIL.n209 0.155672
R1504 VTAIL.n221 VTAIL.n209 0.155672
R1505 VTAIL.n222 VTAIL.n221 0.155672
R1506 VTAIL.n222 VTAIL.n205 0.155672
R1507 VTAIL.n229 VTAIL.n205 0.155672
R1508 VTAIL.n12 VTAIL.n7 0.155672
R1509 VTAIL.n19 VTAIL.n7 0.155672
R1510 VTAIL.n20 VTAIL.n19 0.155672
R1511 VTAIL.n20 VTAIL.n3 0.155672
R1512 VTAIL.n27 VTAIL.n3 0.155672
R1513 VTAIL.n40 VTAIL.n35 0.155672
R1514 VTAIL.n47 VTAIL.n35 0.155672
R1515 VTAIL.n48 VTAIL.n47 0.155672
R1516 VTAIL.n48 VTAIL.n31 0.155672
R1517 VTAIL.n55 VTAIL.n31 0.155672
R1518 VTAIL.n70 VTAIL.n65 0.155672
R1519 VTAIL.n77 VTAIL.n65 0.155672
R1520 VTAIL.n78 VTAIL.n77 0.155672
R1521 VTAIL.n78 VTAIL.n61 0.155672
R1522 VTAIL.n85 VTAIL.n61 0.155672
R1523 VTAIL.n201 VTAIL.n177 0.155672
R1524 VTAIL.n194 VTAIL.n177 0.155672
R1525 VTAIL.n194 VTAIL.n193 0.155672
R1526 VTAIL.n193 VTAIL.n181 0.155672
R1527 VTAIL.n186 VTAIL.n181 0.155672
R1528 VTAIL.n171 VTAIL.n147 0.155672
R1529 VTAIL.n164 VTAIL.n147 0.155672
R1530 VTAIL.n164 VTAIL.n163 0.155672
R1531 VTAIL.n163 VTAIL.n151 0.155672
R1532 VTAIL.n156 VTAIL.n151 0.155672
R1533 VTAIL.n143 VTAIL.n119 0.155672
R1534 VTAIL.n136 VTAIL.n119 0.155672
R1535 VTAIL.n136 VTAIL.n135 0.155672
R1536 VTAIL.n135 VTAIL.n123 0.155672
R1537 VTAIL.n128 VTAIL.n123 0.155672
R1538 VTAIL.n113 VTAIL.n89 0.155672
R1539 VTAIL.n106 VTAIL.n89 0.155672
R1540 VTAIL.n106 VTAIL.n105 0.155672
R1541 VTAIL.n105 VTAIL.n93 0.155672
R1542 VTAIL.n98 VTAIL.n93 0.155672
R1543 VTAIL VTAIL.n1 0.0586897
R1544 VDD1 VDD1.n0 100.621
R1545 VDD1.n3 VDD1.n2 100.507
R1546 VDD1.n3 VDD1.n1 100.507
R1547 VDD1.n5 VDD1.n4 99.0762
R1548 VDD1.n5 VDD1.n3 42.3112
R1549 VDD1.n4 VDD1.t5 6.05357
R1550 VDD1.n4 VDD1.t0 6.05357
R1551 VDD1.n0 VDD1.t4 6.05357
R1552 VDD1.n0 VDD1.t2 6.05357
R1553 VDD1.n2 VDD1.t1 6.05357
R1554 VDD1.n2 VDD1.t7 6.05357
R1555 VDD1.n1 VDD1.t3 6.05357
R1556 VDD1.n1 VDD1.t6 6.05357
R1557 VDD1 VDD1.n5 1.42938
R1558 VN.n60 VN.n59 161.3
R1559 VN.n58 VN.n32 161.3
R1560 VN.n57 VN.n56 161.3
R1561 VN.n55 VN.n33 161.3
R1562 VN.n54 VN.n53 161.3
R1563 VN.n52 VN.n34 161.3
R1564 VN.n51 VN.n50 161.3
R1565 VN.n49 VN.n48 161.3
R1566 VN.n47 VN.n36 161.3
R1567 VN.n46 VN.n45 161.3
R1568 VN.n44 VN.n37 161.3
R1569 VN.n43 VN.n42 161.3
R1570 VN.n41 VN.n38 161.3
R1571 VN.n29 VN.n28 161.3
R1572 VN.n27 VN.n1 161.3
R1573 VN.n26 VN.n25 161.3
R1574 VN.n24 VN.n2 161.3
R1575 VN.n23 VN.n22 161.3
R1576 VN.n21 VN.n3 161.3
R1577 VN.n20 VN.n19 161.3
R1578 VN.n18 VN.n17 161.3
R1579 VN.n16 VN.n5 161.3
R1580 VN.n15 VN.n14 161.3
R1581 VN.n13 VN.n6 161.3
R1582 VN.n12 VN.n11 161.3
R1583 VN.n10 VN.n7 161.3
R1584 VN.n39 VN.t2 74.8935
R1585 VN.n8 VN.t0 74.8935
R1586 VN.n30 VN.n0 69.2705
R1587 VN.n61 VN.n31 69.2705
R1588 VN.n15 VN.n6 56.5193
R1589 VN.n26 VN.n2 56.5193
R1590 VN.n46 VN.n37 56.5193
R1591 VN.n57 VN.n33 56.5193
R1592 VN.n9 VN.n8 50.6608
R1593 VN.n40 VN.n39 50.6608
R1594 VN VN.n61 48.6344
R1595 VN.n9 VN.t6 41.4803
R1596 VN.n4 VN.t1 41.4803
R1597 VN.n0 VN.t7 41.4803
R1598 VN.n40 VN.t3 41.4803
R1599 VN.n35 VN.t5 41.4803
R1600 VN.n31 VN.t4 41.4803
R1601 VN.n11 VN.n10 24.4675
R1602 VN.n11 VN.n6 24.4675
R1603 VN.n16 VN.n15 24.4675
R1604 VN.n17 VN.n16 24.4675
R1605 VN.n21 VN.n20 24.4675
R1606 VN.n22 VN.n21 24.4675
R1607 VN.n22 VN.n2 24.4675
R1608 VN.n27 VN.n26 24.4675
R1609 VN.n28 VN.n27 24.4675
R1610 VN.n42 VN.n37 24.4675
R1611 VN.n42 VN.n41 24.4675
R1612 VN.n53 VN.n33 24.4675
R1613 VN.n53 VN.n52 24.4675
R1614 VN.n52 VN.n51 24.4675
R1615 VN.n48 VN.n47 24.4675
R1616 VN.n47 VN.n46 24.4675
R1617 VN.n59 VN.n58 24.4675
R1618 VN.n58 VN.n57 24.4675
R1619 VN.n10 VN.n9 23.2442
R1620 VN.n17 VN.n4 23.2442
R1621 VN.n41 VN.n40 23.2442
R1622 VN.n48 VN.n35 23.2442
R1623 VN.n28 VN.n0 20.7975
R1624 VN.n59 VN.n31 20.7975
R1625 VN.n39 VN.n38 3.87633
R1626 VN.n8 VN.n7 3.87633
R1627 VN.n20 VN.n4 1.22385
R1628 VN.n51 VN.n35 1.22385
R1629 VN.n61 VN.n60 0.354971
R1630 VN.n30 VN.n29 0.354971
R1631 VN VN.n30 0.26696
R1632 VN.n60 VN.n32 0.189894
R1633 VN.n56 VN.n32 0.189894
R1634 VN.n56 VN.n55 0.189894
R1635 VN.n55 VN.n54 0.189894
R1636 VN.n54 VN.n34 0.189894
R1637 VN.n50 VN.n34 0.189894
R1638 VN.n50 VN.n49 0.189894
R1639 VN.n49 VN.n36 0.189894
R1640 VN.n45 VN.n36 0.189894
R1641 VN.n45 VN.n44 0.189894
R1642 VN.n44 VN.n43 0.189894
R1643 VN.n43 VN.n38 0.189894
R1644 VN.n12 VN.n7 0.189894
R1645 VN.n13 VN.n12 0.189894
R1646 VN.n14 VN.n13 0.189894
R1647 VN.n14 VN.n5 0.189894
R1648 VN.n18 VN.n5 0.189894
R1649 VN.n19 VN.n18 0.189894
R1650 VN.n19 VN.n3 0.189894
R1651 VN.n23 VN.n3 0.189894
R1652 VN.n24 VN.n23 0.189894
R1653 VN.n25 VN.n24 0.189894
R1654 VN.n25 VN.n1 0.189894
R1655 VN.n29 VN.n1 0.189894
R1656 VDD2.n2 VDD2.n1 100.507
R1657 VDD2.n2 VDD2.n0 100.507
R1658 VDD2 VDD2.n5 100.505
R1659 VDD2.n4 VDD2.n3 99.0764
R1660 VDD2.n4 VDD2.n2 41.7282
R1661 VDD2.n5 VDD2.t4 6.05357
R1662 VDD2.n5 VDD2.t5 6.05357
R1663 VDD2.n3 VDD2.t3 6.05357
R1664 VDD2.n3 VDD2.t2 6.05357
R1665 VDD2.n1 VDD2.t6 6.05357
R1666 VDD2.n1 VDD2.t0 6.05357
R1667 VDD2.n0 VDD2.t7 6.05357
R1668 VDD2.n0 VDD2.t1 6.05357
R1669 VDD2 VDD2.n4 1.54576
C0 VDD2 w_n4420_n2042# 2.08325f
C1 VDD1 VN 0.152792f
C2 VDD2 VN 4.27387f
C3 B VTAIL 2.95312f
C4 VP B 2.22677f
C5 w_n4420_n2042# B 9.06845f
C6 VDD2 VDD1 2.04916f
C7 B VN 1.25953f
C8 VP VTAIL 5.37654f
C9 w_n4420_n2042# VTAIL 2.78392f
C10 VDD1 B 1.6291f
C11 w_n4420_n2042# VP 9.599191f
C12 VDD2 B 1.74168f
C13 VTAIL VN 5.36244f
C14 VP VN 7.07058f
C15 w_n4420_n2042# VN 9.0239f
C16 VDD1 VTAIL 6.2167f
C17 VDD1 VP 4.69446f
C18 VDD2 VTAIL 6.274601f
C19 VDD2 VP 0.579139f
C20 VDD1 w_n4420_n2042# 1.94696f
C21 VDD2 VSUBS 2.049717f
C22 VDD1 VSUBS 2.61484f
C23 VTAIL VSUBS 0.732869f
C24 VN VSUBS 7.238821f
C25 VP VSUBS 3.679238f
C26 B VSUBS 4.87009f
C27 w_n4420_n2042# VSUBS 0.112922p
C28 VDD2.t7 VSUBS 0.142523f
C29 VDD2.t1 VSUBS 0.142523f
C30 VDD2.n0 VSUBS 0.931099f
C31 VDD2.t6 VSUBS 0.142523f
C32 VDD2.t0 VSUBS 0.142523f
C33 VDD2.n1 VSUBS 0.931099f
C34 VDD2.n2 VSUBS 4.75895f
C35 VDD2.t3 VSUBS 0.142523f
C36 VDD2.t2 VSUBS 0.142523f
C37 VDD2.n3 VSUBS 0.916633f
C38 VDD2.n4 VSUBS 3.76856f
C39 VDD2.t4 VSUBS 0.142523f
C40 VDD2.t5 VSUBS 0.142523f
C41 VDD2.n5 VSUBS 0.931059f
C42 VN.t7 VSUBS 1.56051f
C43 VN.n0 VSUBS 0.734162f
C44 VN.n1 VSUBS 0.035435f
C45 VN.n2 VSUBS 0.046791f
C46 VN.n3 VSUBS 0.035435f
C47 VN.t1 VSUBS 1.56051f
C48 VN.n4 VSUBS 0.587198f
C49 VN.n5 VSUBS 0.035435f
C50 VN.n6 VSUBS 0.051728f
C51 VN.n7 VSUBS 0.404175f
C52 VN.t6 VSUBS 1.56051f
C53 VN.t0 VSUBS 1.93601f
C54 VN.n8 VSUBS 0.67502f
C55 VN.n9 VSUBS 0.718603f
C56 VN.n10 VSUBS 0.064409f
C57 VN.n11 VSUBS 0.066041f
C58 VN.n12 VSUBS 0.035435f
C59 VN.n13 VSUBS 0.035435f
C60 VN.n14 VSUBS 0.035435f
C61 VN.n15 VSUBS 0.051728f
C62 VN.n16 VSUBS 0.066041f
C63 VN.n17 VSUBS 0.064409f
C64 VN.n18 VSUBS 0.035435f
C65 VN.n19 VSUBS 0.035435f
C66 VN.n20 VSUBS 0.035065f
C67 VN.n21 VSUBS 0.066041f
C68 VN.n22 VSUBS 0.066041f
C69 VN.n23 VSUBS 0.035435f
C70 VN.n24 VSUBS 0.035435f
C71 VN.n25 VSUBS 0.035435f
C72 VN.n26 VSUBS 0.056665f
C73 VN.n27 VSUBS 0.066041f
C74 VN.n28 VSUBS 0.061149f
C75 VN.n29 VSUBS 0.057191f
C76 VN.n30 VSUBS 0.073781f
C77 VN.t4 VSUBS 1.56051f
C78 VN.n31 VSUBS 0.734162f
C79 VN.n32 VSUBS 0.035435f
C80 VN.n33 VSUBS 0.046791f
C81 VN.n34 VSUBS 0.035435f
C82 VN.t5 VSUBS 1.56051f
C83 VN.n35 VSUBS 0.587198f
C84 VN.n36 VSUBS 0.035435f
C85 VN.n37 VSUBS 0.051728f
C86 VN.n38 VSUBS 0.404175f
C87 VN.t3 VSUBS 1.56051f
C88 VN.t2 VSUBS 1.93601f
C89 VN.n39 VSUBS 0.67502f
C90 VN.n40 VSUBS 0.718603f
C91 VN.n41 VSUBS 0.064409f
C92 VN.n42 VSUBS 0.066041f
C93 VN.n43 VSUBS 0.035435f
C94 VN.n44 VSUBS 0.035435f
C95 VN.n45 VSUBS 0.035435f
C96 VN.n46 VSUBS 0.051728f
C97 VN.n47 VSUBS 0.066041f
C98 VN.n48 VSUBS 0.064409f
C99 VN.n49 VSUBS 0.035435f
C100 VN.n50 VSUBS 0.035435f
C101 VN.n51 VSUBS 0.035065f
C102 VN.n52 VSUBS 0.066041f
C103 VN.n53 VSUBS 0.066041f
C104 VN.n54 VSUBS 0.035435f
C105 VN.n55 VSUBS 0.035435f
C106 VN.n56 VSUBS 0.035435f
C107 VN.n57 VSUBS 0.056665f
C108 VN.n58 VSUBS 0.066041f
C109 VN.n59 VSUBS 0.061149f
C110 VN.n60 VSUBS 0.057191f
C111 VN.n61 VSUBS 1.93078f
C112 VDD1.t4 VSUBS 0.124024f
C113 VDD1.t2 VSUBS 0.124024f
C114 VDD1.n0 VSUBS 0.811393f
C115 VDD1.t3 VSUBS 0.124024f
C116 VDD1.t6 VSUBS 0.124024f
C117 VDD1.n1 VSUBS 0.810249f
C118 VDD1.t1 VSUBS 0.124024f
C119 VDD1.t7 VSUBS 0.124024f
C120 VDD1.n2 VSUBS 0.810249f
C121 VDD1.n3 VSUBS 4.20203f
C122 VDD1.t5 VSUBS 0.124024f
C123 VDD1.t0 VSUBS 0.124024f
C124 VDD1.n4 VSUBS 0.797657f
C125 VDD1.n5 VSUBS 3.31567f
C126 VTAIL.t5 VSUBS 0.131787f
C127 VTAIL.t4 VSUBS 0.131787f
C128 VTAIL.n0 VSUBS 0.750522f
C129 VTAIL.n1 VSUBS 0.843708f
C130 VTAIL.n2 VSUBS 0.034652f
C131 VTAIL.n3 VSUBS 0.031056f
C132 VTAIL.n4 VSUBS 0.016688f
C133 VTAIL.n5 VSUBS 0.039445f
C134 VTAIL.n6 VSUBS 0.01767f
C135 VTAIL.n7 VSUBS 0.031056f
C136 VTAIL.n8 VSUBS 0.016688f
C137 VTAIL.n9 VSUBS 0.029583f
C138 VTAIL.n10 VSUBS 0.025055f
C139 VTAIL.t7 VSUBS 0.085317f
C140 VTAIL.n11 VSUBS 0.132184f
C141 VTAIL.n12 VSUBS 0.622237f
C142 VTAIL.n13 VSUBS 0.016688f
C143 VTAIL.n14 VSUBS 0.01767f
C144 VTAIL.n15 VSUBS 0.039445f
C145 VTAIL.n16 VSUBS 0.039445f
C146 VTAIL.n17 VSUBS 0.01767f
C147 VTAIL.n18 VSUBS 0.016688f
C148 VTAIL.n19 VSUBS 0.031056f
C149 VTAIL.n20 VSUBS 0.031056f
C150 VTAIL.n21 VSUBS 0.016688f
C151 VTAIL.n22 VSUBS 0.01767f
C152 VTAIL.n23 VSUBS 0.039445f
C153 VTAIL.n24 VSUBS 0.097291f
C154 VTAIL.n25 VSUBS 0.01767f
C155 VTAIL.n26 VSUBS 0.016688f
C156 VTAIL.n27 VSUBS 0.075603f
C157 VTAIL.n28 VSUBS 0.049121f
C158 VTAIL.n29 VSUBS 0.373317f
C159 VTAIL.n30 VSUBS 0.034652f
C160 VTAIL.n31 VSUBS 0.031056f
C161 VTAIL.n32 VSUBS 0.016688f
C162 VTAIL.n33 VSUBS 0.039445f
C163 VTAIL.n34 VSUBS 0.01767f
C164 VTAIL.n35 VSUBS 0.031056f
C165 VTAIL.n36 VSUBS 0.016688f
C166 VTAIL.n37 VSUBS 0.029583f
C167 VTAIL.n38 VSUBS 0.025055f
C168 VTAIL.t9 VSUBS 0.085317f
C169 VTAIL.n39 VSUBS 0.132184f
C170 VTAIL.n40 VSUBS 0.622237f
C171 VTAIL.n41 VSUBS 0.016688f
C172 VTAIL.n42 VSUBS 0.01767f
C173 VTAIL.n43 VSUBS 0.039445f
C174 VTAIL.n44 VSUBS 0.039445f
C175 VTAIL.n45 VSUBS 0.01767f
C176 VTAIL.n46 VSUBS 0.016688f
C177 VTAIL.n47 VSUBS 0.031056f
C178 VTAIL.n48 VSUBS 0.031056f
C179 VTAIL.n49 VSUBS 0.016688f
C180 VTAIL.n50 VSUBS 0.01767f
C181 VTAIL.n51 VSUBS 0.039445f
C182 VTAIL.n52 VSUBS 0.097291f
C183 VTAIL.n53 VSUBS 0.01767f
C184 VTAIL.n54 VSUBS 0.016688f
C185 VTAIL.n55 VSUBS 0.075603f
C186 VTAIL.n56 VSUBS 0.049121f
C187 VTAIL.n57 VSUBS 0.373317f
C188 VTAIL.t12 VSUBS 0.131787f
C189 VTAIL.t8 VSUBS 0.131787f
C190 VTAIL.n58 VSUBS 0.750522f
C191 VTAIL.n59 VSUBS 1.13551f
C192 VTAIL.n60 VSUBS 0.034652f
C193 VTAIL.n61 VSUBS 0.031056f
C194 VTAIL.n62 VSUBS 0.016688f
C195 VTAIL.n63 VSUBS 0.039445f
C196 VTAIL.n64 VSUBS 0.01767f
C197 VTAIL.n65 VSUBS 0.031056f
C198 VTAIL.n66 VSUBS 0.016688f
C199 VTAIL.n67 VSUBS 0.029583f
C200 VTAIL.n68 VSUBS 0.025055f
C201 VTAIL.t13 VSUBS 0.085317f
C202 VTAIL.n69 VSUBS 0.132184f
C203 VTAIL.n70 VSUBS 0.622237f
C204 VTAIL.n71 VSUBS 0.016688f
C205 VTAIL.n72 VSUBS 0.01767f
C206 VTAIL.n73 VSUBS 0.039445f
C207 VTAIL.n74 VSUBS 0.039445f
C208 VTAIL.n75 VSUBS 0.01767f
C209 VTAIL.n76 VSUBS 0.016688f
C210 VTAIL.n77 VSUBS 0.031056f
C211 VTAIL.n78 VSUBS 0.031056f
C212 VTAIL.n79 VSUBS 0.016688f
C213 VTAIL.n80 VSUBS 0.01767f
C214 VTAIL.n81 VSUBS 0.039445f
C215 VTAIL.n82 VSUBS 0.097291f
C216 VTAIL.n83 VSUBS 0.01767f
C217 VTAIL.n84 VSUBS 0.016688f
C218 VTAIL.n85 VSUBS 0.075603f
C219 VTAIL.n86 VSUBS 0.049121f
C220 VTAIL.n87 VSUBS 1.50903f
C221 VTAIL.n88 VSUBS 0.034652f
C222 VTAIL.n89 VSUBS 0.031056f
C223 VTAIL.n90 VSUBS 0.016688f
C224 VTAIL.n91 VSUBS 0.039445f
C225 VTAIL.n92 VSUBS 0.01767f
C226 VTAIL.n93 VSUBS 0.031056f
C227 VTAIL.n94 VSUBS 0.016688f
C228 VTAIL.n95 VSUBS 0.029583f
C229 VTAIL.n96 VSUBS 0.025055f
C230 VTAIL.t6 VSUBS 0.085317f
C231 VTAIL.n97 VSUBS 0.132184f
C232 VTAIL.n98 VSUBS 0.622237f
C233 VTAIL.n99 VSUBS 0.016688f
C234 VTAIL.n100 VSUBS 0.01767f
C235 VTAIL.n101 VSUBS 0.039445f
C236 VTAIL.n102 VSUBS 0.039445f
C237 VTAIL.n103 VSUBS 0.01767f
C238 VTAIL.n104 VSUBS 0.016688f
C239 VTAIL.n105 VSUBS 0.031056f
C240 VTAIL.n106 VSUBS 0.031056f
C241 VTAIL.n107 VSUBS 0.016688f
C242 VTAIL.n108 VSUBS 0.01767f
C243 VTAIL.n109 VSUBS 0.039445f
C244 VTAIL.n110 VSUBS 0.097291f
C245 VTAIL.n111 VSUBS 0.01767f
C246 VTAIL.n112 VSUBS 0.016688f
C247 VTAIL.n113 VSUBS 0.075603f
C248 VTAIL.n114 VSUBS 0.049121f
C249 VTAIL.n115 VSUBS 1.50903f
C250 VTAIL.t0 VSUBS 0.131787f
C251 VTAIL.t3 VSUBS 0.131787f
C252 VTAIL.n116 VSUBS 0.750527f
C253 VTAIL.n117 VSUBS 1.1355f
C254 VTAIL.n118 VSUBS 0.034652f
C255 VTAIL.n119 VSUBS 0.031056f
C256 VTAIL.n120 VSUBS 0.016688f
C257 VTAIL.n121 VSUBS 0.039445f
C258 VTAIL.n122 VSUBS 0.01767f
C259 VTAIL.n123 VSUBS 0.031056f
C260 VTAIL.n124 VSUBS 0.016688f
C261 VTAIL.n125 VSUBS 0.029583f
C262 VTAIL.n126 VSUBS 0.025055f
C263 VTAIL.t2 VSUBS 0.085317f
C264 VTAIL.n127 VSUBS 0.132184f
C265 VTAIL.n128 VSUBS 0.622237f
C266 VTAIL.n129 VSUBS 0.016688f
C267 VTAIL.n130 VSUBS 0.01767f
C268 VTAIL.n131 VSUBS 0.039445f
C269 VTAIL.n132 VSUBS 0.039445f
C270 VTAIL.n133 VSUBS 0.01767f
C271 VTAIL.n134 VSUBS 0.016688f
C272 VTAIL.n135 VSUBS 0.031056f
C273 VTAIL.n136 VSUBS 0.031056f
C274 VTAIL.n137 VSUBS 0.016688f
C275 VTAIL.n138 VSUBS 0.01767f
C276 VTAIL.n139 VSUBS 0.039445f
C277 VTAIL.n140 VSUBS 0.097291f
C278 VTAIL.n141 VSUBS 0.01767f
C279 VTAIL.n142 VSUBS 0.016688f
C280 VTAIL.n143 VSUBS 0.075603f
C281 VTAIL.n144 VSUBS 0.049121f
C282 VTAIL.n145 VSUBS 0.373317f
C283 VTAIL.n146 VSUBS 0.034652f
C284 VTAIL.n147 VSUBS 0.031056f
C285 VTAIL.n148 VSUBS 0.016688f
C286 VTAIL.n149 VSUBS 0.039445f
C287 VTAIL.n150 VSUBS 0.01767f
C288 VTAIL.n151 VSUBS 0.031056f
C289 VTAIL.n152 VSUBS 0.016688f
C290 VTAIL.n153 VSUBS 0.029583f
C291 VTAIL.n154 VSUBS 0.025055f
C292 VTAIL.t15 VSUBS 0.085317f
C293 VTAIL.n155 VSUBS 0.132184f
C294 VTAIL.n156 VSUBS 0.622237f
C295 VTAIL.n157 VSUBS 0.016688f
C296 VTAIL.n158 VSUBS 0.01767f
C297 VTAIL.n159 VSUBS 0.039445f
C298 VTAIL.n160 VSUBS 0.039445f
C299 VTAIL.n161 VSUBS 0.01767f
C300 VTAIL.n162 VSUBS 0.016688f
C301 VTAIL.n163 VSUBS 0.031056f
C302 VTAIL.n164 VSUBS 0.031056f
C303 VTAIL.n165 VSUBS 0.016688f
C304 VTAIL.n166 VSUBS 0.01767f
C305 VTAIL.n167 VSUBS 0.039445f
C306 VTAIL.n168 VSUBS 0.097291f
C307 VTAIL.n169 VSUBS 0.01767f
C308 VTAIL.n170 VSUBS 0.016688f
C309 VTAIL.n171 VSUBS 0.075603f
C310 VTAIL.n172 VSUBS 0.049121f
C311 VTAIL.n173 VSUBS 0.373317f
C312 VTAIL.t14 VSUBS 0.131787f
C313 VTAIL.t10 VSUBS 0.131787f
C314 VTAIL.n174 VSUBS 0.750527f
C315 VTAIL.n175 VSUBS 1.1355f
C316 VTAIL.n176 VSUBS 0.034652f
C317 VTAIL.n177 VSUBS 0.031056f
C318 VTAIL.n178 VSUBS 0.016688f
C319 VTAIL.n179 VSUBS 0.039445f
C320 VTAIL.n180 VSUBS 0.01767f
C321 VTAIL.n181 VSUBS 0.031056f
C322 VTAIL.n182 VSUBS 0.016688f
C323 VTAIL.n183 VSUBS 0.029583f
C324 VTAIL.n184 VSUBS 0.025055f
C325 VTAIL.t11 VSUBS 0.085317f
C326 VTAIL.n185 VSUBS 0.132184f
C327 VTAIL.n186 VSUBS 0.622237f
C328 VTAIL.n187 VSUBS 0.016688f
C329 VTAIL.n188 VSUBS 0.01767f
C330 VTAIL.n189 VSUBS 0.039445f
C331 VTAIL.n190 VSUBS 0.039445f
C332 VTAIL.n191 VSUBS 0.01767f
C333 VTAIL.n192 VSUBS 0.016688f
C334 VTAIL.n193 VSUBS 0.031056f
C335 VTAIL.n194 VSUBS 0.031056f
C336 VTAIL.n195 VSUBS 0.016688f
C337 VTAIL.n196 VSUBS 0.01767f
C338 VTAIL.n197 VSUBS 0.039445f
C339 VTAIL.n198 VSUBS 0.097291f
C340 VTAIL.n199 VSUBS 0.01767f
C341 VTAIL.n200 VSUBS 0.016688f
C342 VTAIL.n201 VSUBS 0.075603f
C343 VTAIL.n202 VSUBS 0.049121f
C344 VTAIL.n203 VSUBS 1.50903f
C345 VTAIL.n204 VSUBS 0.034652f
C346 VTAIL.n205 VSUBS 0.031056f
C347 VTAIL.n206 VSUBS 0.016688f
C348 VTAIL.n207 VSUBS 0.039445f
C349 VTAIL.n208 VSUBS 0.01767f
C350 VTAIL.n209 VSUBS 0.031056f
C351 VTAIL.n210 VSUBS 0.016688f
C352 VTAIL.n211 VSUBS 0.029583f
C353 VTAIL.n212 VSUBS 0.025055f
C354 VTAIL.t1 VSUBS 0.085317f
C355 VTAIL.n213 VSUBS 0.132184f
C356 VTAIL.n214 VSUBS 0.622237f
C357 VTAIL.n215 VSUBS 0.016688f
C358 VTAIL.n216 VSUBS 0.01767f
C359 VTAIL.n217 VSUBS 0.039445f
C360 VTAIL.n218 VSUBS 0.039445f
C361 VTAIL.n219 VSUBS 0.01767f
C362 VTAIL.n220 VSUBS 0.016688f
C363 VTAIL.n221 VSUBS 0.031056f
C364 VTAIL.n222 VSUBS 0.031056f
C365 VTAIL.n223 VSUBS 0.016688f
C366 VTAIL.n224 VSUBS 0.01767f
C367 VTAIL.n225 VSUBS 0.039445f
C368 VTAIL.n226 VSUBS 0.097291f
C369 VTAIL.n227 VSUBS 0.01767f
C370 VTAIL.n228 VSUBS 0.016688f
C371 VTAIL.n229 VSUBS 0.075603f
C372 VTAIL.n230 VSUBS 0.049121f
C373 VTAIL.n231 VSUBS 1.50321f
C374 VP.t0 VSUBS 1.75746f
C375 VP.n0 VSUBS 0.826817f
C376 VP.n1 VSUBS 0.039907f
C377 VP.n2 VSUBS 0.052696f
C378 VP.n3 VSUBS 0.039907f
C379 VP.t6 VSUBS 1.75746f
C380 VP.n4 VSUBS 0.661305f
C381 VP.n5 VSUBS 0.039907f
C382 VP.n6 VSUBS 0.058257f
C383 VP.n7 VSUBS 0.039907f
C384 VP.t1 VSUBS 1.75746f
C385 VP.n8 VSUBS 0.074376f
C386 VP.n9 VSUBS 0.039907f
C387 VP.n10 VSUBS 0.074376f
C388 VP.t7 VSUBS 1.75746f
C389 VP.n11 VSUBS 0.826817f
C390 VP.n12 VSUBS 0.039907f
C391 VP.n13 VSUBS 0.052696f
C392 VP.n14 VSUBS 0.039907f
C393 VP.t2 VSUBS 1.75746f
C394 VP.n15 VSUBS 0.661305f
C395 VP.n16 VSUBS 0.039907f
C396 VP.n17 VSUBS 0.058257f
C397 VP.n18 VSUBS 0.455184f
C398 VP.t5 VSUBS 1.75746f
C399 VP.t3 VSUBS 2.18034f
C400 VP.n19 VSUBS 0.760213f
C401 VP.n20 VSUBS 0.809295f
C402 VP.n21 VSUBS 0.072538f
C403 VP.n22 VSUBS 0.074376f
C404 VP.n23 VSUBS 0.039907f
C405 VP.n24 VSUBS 0.039907f
C406 VP.n25 VSUBS 0.039907f
C407 VP.n26 VSUBS 0.058257f
C408 VP.n27 VSUBS 0.074376f
C409 VP.n28 VSUBS 0.072538f
C410 VP.n29 VSUBS 0.039907f
C411 VP.n30 VSUBS 0.039907f
C412 VP.n31 VSUBS 0.03949f
C413 VP.n32 VSUBS 0.074376f
C414 VP.n33 VSUBS 0.074376f
C415 VP.n34 VSUBS 0.039907f
C416 VP.n35 VSUBS 0.039907f
C417 VP.n36 VSUBS 0.039907f
C418 VP.n37 VSUBS 0.063817f
C419 VP.n38 VSUBS 0.074376f
C420 VP.n39 VSUBS 0.068866f
C421 VP.n40 VSUBS 0.064409f
C422 VP.n41 VSUBS 2.15796f
C423 VP.n42 VSUBS 2.18756f
C424 VP.t4 VSUBS 1.75746f
C425 VP.n43 VSUBS 0.826817f
C426 VP.n44 VSUBS 0.068866f
C427 VP.n45 VSUBS 0.064409f
C428 VP.n46 VSUBS 0.039907f
C429 VP.n47 VSUBS 0.039907f
C430 VP.n48 VSUBS 0.063817f
C431 VP.n49 VSUBS 0.052696f
C432 VP.n50 VSUBS 0.074376f
C433 VP.n51 VSUBS 0.039907f
C434 VP.n52 VSUBS 0.039907f
C435 VP.n53 VSUBS 0.039907f
C436 VP.n54 VSUBS 0.03949f
C437 VP.n55 VSUBS 0.661305f
C438 VP.n56 VSUBS 0.072538f
C439 VP.n57 VSUBS 0.074376f
C440 VP.n58 VSUBS 0.039907f
C441 VP.n59 VSUBS 0.039907f
C442 VP.n60 VSUBS 0.039907f
C443 VP.n61 VSUBS 0.058257f
C444 VP.n62 VSUBS 0.074376f
C445 VP.n63 VSUBS 0.072538f
C446 VP.n64 VSUBS 0.039907f
C447 VP.n65 VSUBS 0.039907f
C448 VP.n66 VSUBS 0.03949f
C449 VP.n67 VSUBS 0.074376f
C450 VP.n68 VSUBS 0.074376f
C451 VP.n69 VSUBS 0.039907f
C452 VP.n70 VSUBS 0.039907f
C453 VP.n71 VSUBS 0.039907f
C454 VP.n72 VSUBS 0.063817f
C455 VP.n73 VSUBS 0.074376f
C456 VP.n74 VSUBS 0.068866f
C457 VP.n75 VSUBS 0.064409f
C458 VP.n76 VSUBS 0.083093f
C459 B.n0 VSUBS 0.006142f
C460 B.n1 VSUBS 0.006142f
C461 B.n2 VSUBS 0.009712f
C462 B.n3 VSUBS 0.009712f
C463 B.n4 VSUBS 0.009712f
C464 B.n5 VSUBS 0.009712f
C465 B.n6 VSUBS 0.009712f
C466 B.n7 VSUBS 0.009712f
C467 B.n8 VSUBS 0.009712f
C468 B.n9 VSUBS 0.009712f
C469 B.n10 VSUBS 0.009712f
C470 B.n11 VSUBS 0.009712f
C471 B.n12 VSUBS 0.009712f
C472 B.n13 VSUBS 0.009712f
C473 B.n14 VSUBS 0.009712f
C474 B.n15 VSUBS 0.009712f
C475 B.n16 VSUBS 0.009712f
C476 B.n17 VSUBS 0.009712f
C477 B.n18 VSUBS 0.009712f
C478 B.n19 VSUBS 0.009712f
C479 B.n20 VSUBS 0.009712f
C480 B.n21 VSUBS 0.009712f
C481 B.n22 VSUBS 0.009712f
C482 B.n23 VSUBS 0.009712f
C483 B.n24 VSUBS 0.009712f
C484 B.n25 VSUBS 0.009712f
C485 B.n26 VSUBS 0.009712f
C486 B.n27 VSUBS 0.009712f
C487 B.n28 VSUBS 0.009712f
C488 B.n29 VSUBS 0.009712f
C489 B.n30 VSUBS 0.009712f
C490 B.n31 VSUBS 0.020888f
C491 B.n32 VSUBS 0.009712f
C492 B.n33 VSUBS 0.009712f
C493 B.n34 VSUBS 0.009712f
C494 B.n35 VSUBS 0.009712f
C495 B.n36 VSUBS 0.009712f
C496 B.n37 VSUBS 0.009712f
C497 B.n38 VSUBS 0.009712f
C498 B.n39 VSUBS 0.009712f
C499 B.n40 VSUBS 0.009712f
C500 B.n41 VSUBS 0.009712f
C501 B.n42 VSUBS 0.009141f
C502 B.n43 VSUBS 0.009712f
C503 B.t5 VSUBS 0.109529f
C504 B.t4 VSUBS 0.148569f
C505 B.t3 VSUBS 1.11367f
C506 B.n44 VSUBS 0.251081f
C507 B.n45 VSUBS 0.203076f
C508 B.n46 VSUBS 0.022502f
C509 B.n47 VSUBS 0.009712f
C510 B.n48 VSUBS 0.009712f
C511 B.n49 VSUBS 0.009712f
C512 B.n50 VSUBS 0.009712f
C513 B.t2 VSUBS 0.109532f
C514 B.t1 VSUBS 0.148571f
C515 B.t0 VSUBS 1.11367f
C516 B.n51 VSUBS 0.251079f
C517 B.n52 VSUBS 0.203074f
C518 B.n53 VSUBS 0.009712f
C519 B.n54 VSUBS 0.009712f
C520 B.n55 VSUBS 0.009712f
C521 B.n56 VSUBS 0.009712f
C522 B.n57 VSUBS 0.009712f
C523 B.n58 VSUBS 0.009712f
C524 B.n59 VSUBS 0.009712f
C525 B.n60 VSUBS 0.009712f
C526 B.n61 VSUBS 0.009712f
C527 B.n62 VSUBS 0.009712f
C528 B.n63 VSUBS 0.020704f
C529 B.n64 VSUBS 0.009712f
C530 B.n65 VSUBS 0.009712f
C531 B.n66 VSUBS 0.009712f
C532 B.n67 VSUBS 0.009712f
C533 B.n68 VSUBS 0.009712f
C534 B.n69 VSUBS 0.009712f
C535 B.n70 VSUBS 0.009712f
C536 B.n71 VSUBS 0.009712f
C537 B.n72 VSUBS 0.009712f
C538 B.n73 VSUBS 0.009712f
C539 B.n74 VSUBS 0.009712f
C540 B.n75 VSUBS 0.009712f
C541 B.n76 VSUBS 0.009712f
C542 B.n77 VSUBS 0.009712f
C543 B.n78 VSUBS 0.009712f
C544 B.n79 VSUBS 0.009712f
C545 B.n80 VSUBS 0.009712f
C546 B.n81 VSUBS 0.009712f
C547 B.n82 VSUBS 0.009712f
C548 B.n83 VSUBS 0.009712f
C549 B.n84 VSUBS 0.009712f
C550 B.n85 VSUBS 0.009712f
C551 B.n86 VSUBS 0.009712f
C552 B.n87 VSUBS 0.009712f
C553 B.n88 VSUBS 0.009712f
C554 B.n89 VSUBS 0.009712f
C555 B.n90 VSUBS 0.009712f
C556 B.n91 VSUBS 0.009712f
C557 B.n92 VSUBS 0.009712f
C558 B.n93 VSUBS 0.009712f
C559 B.n94 VSUBS 0.009712f
C560 B.n95 VSUBS 0.009712f
C561 B.n96 VSUBS 0.009712f
C562 B.n97 VSUBS 0.009712f
C563 B.n98 VSUBS 0.009712f
C564 B.n99 VSUBS 0.009712f
C565 B.n100 VSUBS 0.009712f
C566 B.n101 VSUBS 0.009712f
C567 B.n102 VSUBS 0.009712f
C568 B.n103 VSUBS 0.009712f
C569 B.n104 VSUBS 0.009712f
C570 B.n105 VSUBS 0.009712f
C571 B.n106 VSUBS 0.009712f
C572 B.n107 VSUBS 0.009712f
C573 B.n108 VSUBS 0.009712f
C574 B.n109 VSUBS 0.009712f
C575 B.n110 VSUBS 0.009712f
C576 B.n111 VSUBS 0.009712f
C577 B.n112 VSUBS 0.009712f
C578 B.n113 VSUBS 0.009712f
C579 B.n114 VSUBS 0.009712f
C580 B.n115 VSUBS 0.009712f
C581 B.n116 VSUBS 0.009712f
C582 B.n117 VSUBS 0.009712f
C583 B.n118 VSUBS 0.009712f
C584 B.n119 VSUBS 0.009712f
C585 B.n120 VSUBS 0.009712f
C586 B.n121 VSUBS 0.009712f
C587 B.n122 VSUBS 0.009712f
C588 B.n123 VSUBS 0.021961f
C589 B.n124 VSUBS 0.009712f
C590 B.n125 VSUBS 0.009712f
C591 B.n126 VSUBS 0.009712f
C592 B.n127 VSUBS 0.009712f
C593 B.n128 VSUBS 0.009712f
C594 B.n129 VSUBS 0.009712f
C595 B.n130 VSUBS 0.009712f
C596 B.n131 VSUBS 0.009712f
C597 B.n132 VSUBS 0.009712f
C598 B.n133 VSUBS 0.009712f
C599 B.n134 VSUBS 0.009712f
C600 B.t10 VSUBS 0.109532f
C601 B.t11 VSUBS 0.148571f
C602 B.t9 VSUBS 1.11367f
C603 B.n135 VSUBS 0.251079f
C604 B.n136 VSUBS 0.203074f
C605 B.n137 VSUBS 0.009712f
C606 B.n138 VSUBS 0.009712f
C607 B.n139 VSUBS 0.009712f
C608 B.n140 VSUBS 0.009712f
C609 B.t7 VSUBS 0.109529f
C610 B.t8 VSUBS 0.148569f
C611 B.t6 VSUBS 1.11367f
C612 B.n141 VSUBS 0.251081f
C613 B.n142 VSUBS 0.203076f
C614 B.n143 VSUBS 0.022502f
C615 B.n144 VSUBS 0.009712f
C616 B.n145 VSUBS 0.009712f
C617 B.n146 VSUBS 0.009712f
C618 B.n147 VSUBS 0.009712f
C619 B.n148 VSUBS 0.009712f
C620 B.n149 VSUBS 0.009712f
C621 B.n150 VSUBS 0.009712f
C622 B.n151 VSUBS 0.009712f
C623 B.n152 VSUBS 0.009712f
C624 B.n153 VSUBS 0.009712f
C625 B.n154 VSUBS 0.021961f
C626 B.n155 VSUBS 0.009712f
C627 B.n156 VSUBS 0.009712f
C628 B.n157 VSUBS 0.009712f
C629 B.n158 VSUBS 0.009712f
C630 B.n159 VSUBS 0.009712f
C631 B.n160 VSUBS 0.009712f
C632 B.n161 VSUBS 0.009712f
C633 B.n162 VSUBS 0.009712f
C634 B.n163 VSUBS 0.009712f
C635 B.n164 VSUBS 0.009712f
C636 B.n165 VSUBS 0.009712f
C637 B.n166 VSUBS 0.009712f
C638 B.n167 VSUBS 0.009712f
C639 B.n168 VSUBS 0.009712f
C640 B.n169 VSUBS 0.009712f
C641 B.n170 VSUBS 0.009712f
C642 B.n171 VSUBS 0.009712f
C643 B.n172 VSUBS 0.009712f
C644 B.n173 VSUBS 0.009712f
C645 B.n174 VSUBS 0.009712f
C646 B.n175 VSUBS 0.009712f
C647 B.n176 VSUBS 0.009712f
C648 B.n177 VSUBS 0.009712f
C649 B.n178 VSUBS 0.009712f
C650 B.n179 VSUBS 0.009712f
C651 B.n180 VSUBS 0.009712f
C652 B.n181 VSUBS 0.009712f
C653 B.n182 VSUBS 0.009712f
C654 B.n183 VSUBS 0.009712f
C655 B.n184 VSUBS 0.009712f
C656 B.n185 VSUBS 0.009712f
C657 B.n186 VSUBS 0.009712f
C658 B.n187 VSUBS 0.009712f
C659 B.n188 VSUBS 0.009712f
C660 B.n189 VSUBS 0.009712f
C661 B.n190 VSUBS 0.009712f
C662 B.n191 VSUBS 0.009712f
C663 B.n192 VSUBS 0.009712f
C664 B.n193 VSUBS 0.009712f
C665 B.n194 VSUBS 0.009712f
C666 B.n195 VSUBS 0.009712f
C667 B.n196 VSUBS 0.009712f
C668 B.n197 VSUBS 0.009712f
C669 B.n198 VSUBS 0.009712f
C670 B.n199 VSUBS 0.009712f
C671 B.n200 VSUBS 0.009712f
C672 B.n201 VSUBS 0.009712f
C673 B.n202 VSUBS 0.009712f
C674 B.n203 VSUBS 0.009712f
C675 B.n204 VSUBS 0.009712f
C676 B.n205 VSUBS 0.009712f
C677 B.n206 VSUBS 0.009712f
C678 B.n207 VSUBS 0.009712f
C679 B.n208 VSUBS 0.009712f
C680 B.n209 VSUBS 0.009712f
C681 B.n210 VSUBS 0.009712f
C682 B.n211 VSUBS 0.009712f
C683 B.n212 VSUBS 0.009712f
C684 B.n213 VSUBS 0.009712f
C685 B.n214 VSUBS 0.009712f
C686 B.n215 VSUBS 0.009712f
C687 B.n216 VSUBS 0.009712f
C688 B.n217 VSUBS 0.009712f
C689 B.n218 VSUBS 0.009712f
C690 B.n219 VSUBS 0.009712f
C691 B.n220 VSUBS 0.009712f
C692 B.n221 VSUBS 0.009712f
C693 B.n222 VSUBS 0.009712f
C694 B.n223 VSUBS 0.009712f
C695 B.n224 VSUBS 0.009712f
C696 B.n225 VSUBS 0.009712f
C697 B.n226 VSUBS 0.009712f
C698 B.n227 VSUBS 0.009712f
C699 B.n228 VSUBS 0.009712f
C700 B.n229 VSUBS 0.009712f
C701 B.n230 VSUBS 0.009712f
C702 B.n231 VSUBS 0.009712f
C703 B.n232 VSUBS 0.009712f
C704 B.n233 VSUBS 0.009712f
C705 B.n234 VSUBS 0.009712f
C706 B.n235 VSUBS 0.009712f
C707 B.n236 VSUBS 0.009712f
C708 B.n237 VSUBS 0.009712f
C709 B.n238 VSUBS 0.009712f
C710 B.n239 VSUBS 0.009712f
C711 B.n240 VSUBS 0.009712f
C712 B.n241 VSUBS 0.009712f
C713 B.n242 VSUBS 0.009712f
C714 B.n243 VSUBS 0.009712f
C715 B.n244 VSUBS 0.009712f
C716 B.n245 VSUBS 0.009712f
C717 B.n246 VSUBS 0.009712f
C718 B.n247 VSUBS 0.009712f
C719 B.n248 VSUBS 0.009712f
C720 B.n249 VSUBS 0.009712f
C721 B.n250 VSUBS 0.009712f
C722 B.n251 VSUBS 0.009712f
C723 B.n252 VSUBS 0.009712f
C724 B.n253 VSUBS 0.009712f
C725 B.n254 VSUBS 0.009712f
C726 B.n255 VSUBS 0.009712f
C727 B.n256 VSUBS 0.009712f
C728 B.n257 VSUBS 0.009712f
C729 B.n258 VSUBS 0.009712f
C730 B.n259 VSUBS 0.009712f
C731 B.n260 VSUBS 0.009712f
C732 B.n261 VSUBS 0.009712f
C733 B.n262 VSUBS 0.009712f
C734 B.n263 VSUBS 0.009712f
C735 B.n264 VSUBS 0.009712f
C736 B.n265 VSUBS 0.009712f
C737 B.n266 VSUBS 0.009712f
C738 B.n267 VSUBS 0.009712f
C739 B.n268 VSUBS 0.009712f
C740 B.n269 VSUBS 0.020888f
C741 B.n270 VSUBS 0.020888f
C742 B.n271 VSUBS 0.021961f
C743 B.n272 VSUBS 0.009712f
C744 B.n273 VSUBS 0.009712f
C745 B.n274 VSUBS 0.009712f
C746 B.n275 VSUBS 0.009712f
C747 B.n276 VSUBS 0.009712f
C748 B.n277 VSUBS 0.009712f
C749 B.n278 VSUBS 0.009712f
C750 B.n279 VSUBS 0.009712f
C751 B.n280 VSUBS 0.009712f
C752 B.n281 VSUBS 0.009712f
C753 B.n282 VSUBS 0.009712f
C754 B.n283 VSUBS 0.009712f
C755 B.n284 VSUBS 0.009712f
C756 B.n285 VSUBS 0.009712f
C757 B.n286 VSUBS 0.009712f
C758 B.n287 VSUBS 0.009712f
C759 B.n288 VSUBS 0.009712f
C760 B.n289 VSUBS 0.009712f
C761 B.n290 VSUBS 0.009712f
C762 B.n291 VSUBS 0.009712f
C763 B.n292 VSUBS 0.009712f
C764 B.n293 VSUBS 0.009712f
C765 B.n294 VSUBS 0.009712f
C766 B.n295 VSUBS 0.009712f
C767 B.n296 VSUBS 0.009712f
C768 B.n297 VSUBS 0.009712f
C769 B.n298 VSUBS 0.009712f
C770 B.n299 VSUBS 0.009712f
C771 B.n300 VSUBS 0.009712f
C772 B.n301 VSUBS 0.009712f
C773 B.n302 VSUBS 0.009141f
C774 B.n303 VSUBS 0.009712f
C775 B.n304 VSUBS 0.009712f
C776 B.n305 VSUBS 0.005427f
C777 B.n306 VSUBS 0.009712f
C778 B.n307 VSUBS 0.009712f
C779 B.n308 VSUBS 0.009712f
C780 B.n309 VSUBS 0.009712f
C781 B.n310 VSUBS 0.009712f
C782 B.n311 VSUBS 0.009712f
C783 B.n312 VSUBS 0.009712f
C784 B.n313 VSUBS 0.009712f
C785 B.n314 VSUBS 0.009712f
C786 B.n315 VSUBS 0.009712f
C787 B.n316 VSUBS 0.009712f
C788 B.n317 VSUBS 0.009712f
C789 B.n318 VSUBS 0.005427f
C790 B.n319 VSUBS 0.022502f
C791 B.n320 VSUBS 0.009141f
C792 B.n321 VSUBS 0.009712f
C793 B.n322 VSUBS 0.009712f
C794 B.n323 VSUBS 0.009712f
C795 B.n324 VSUBS 0.009712f
C796 B.n325 VSUBS 0.009712f
C797 B.n326 VSUBS 0.009712f
C798 B.n327 VSUBS 0.009712f
C799 B.n328 VSUBS 0.009712f
C800 B.n329 VSUBS 0.009712f
C801 B.n330 VSUBS 0.009712f
C802 B.n331 VSUBS 0.009712f
C803 B.n332 VSUBS 0.009712f
C804 B.n333 VSUBS 0.009712f
C805 B.n334 VSUBS 0.009712f
C806 B.n335 VSUBS 0.009712f
C807 B.n336 VSUBS 0.009712f
C808 B.n337 VSUBS 0.009712f
C809 B.n338 VSUBS 0.009712f
C810 B.n339 VSUBS 0.009712f
C811 B.n340 VSUBS 0.009712f
C812 B.n341 VSUBS 0.009712f
C813 B.n342 VSUBS 0.009712f
C814 B.n343 VSUBS 0.009712f
C815 B.n344 VSUBS 0.009712f
C816 B.n345 VSUBS 0.009712f
C817 B.n346 VSUBS 0.009712f
C818 B.n347 VSUBS 0.009712f
C819 B.n348 VSUBS 0.009712f
C820 B.n349 VSUBS 0.009712f
C821 B.n350 VSUBS 0.009712f
C822 B.n351 VSUBS 0.009712f
C823 B.n352 VSUBS 0.021961f
C824 B.n353 VSUBS 0.020888f
C825 B.n354 VSUBS 0.020888f
C826 B.n355 VSUBS 0.009712f
C827 B.n356 VSUBS 0.009712f
C828 B.n357 VSUBS 0.009712f
C829 B.n358 VSUBS 0.009712f
C830 B.n359 VSUBS 0.009712f
C831 B.n360 VSUBS 0.009712f
C832 B.n361 VSUBS 0.009712f
C833 B.n362 VSUBS 0.009712f
C834 B.n363 VSUBS 0.009712f
C835 B.n364 VSUBS 0.009712f
C836 B.n365 VSUBS 0.009712f
C837 B.n366 VSUBS 0.009712f
C838 B.n367 VSUBS 0.009712f
C839 B.n368 VSUBS 0.009712f
C840 B.n369 VSUBS 0.009712f
C841 B.n370 VSUBS 0.009712f
C842 B.n371 VSUBS 0.009712f
C843 B.n372 VSUBS 0.009712f
C844 B.n373 VSUBS 0.009712f
C845 B.n374 VSUBS 0.009712f
C846 B.n375 VSUBS 0.009712f
C847 B.n376 VSUBS 0.009712f
C848 B.n377 VSUBS 0.009712f
C849 B.n378 VSUBS 0.009712f
C850 B.n379 VSUBS 0.009712f
C851 B.n380 VSUBS 0.009712f
C852 B.n381 VSUBS 0.009712f
C853 B.n382 VSUBS 0.009712f
C854 B.n383 VSUBS 0.009712f
C855 B.n384 VSUBS 0.009712f
C856 B.n385 VSUBS 0.009712f
C857 B.n386 VSUBS 0.009712f
C858 B.n387 VSUBS 0.009712f
C859 B.n388 VSUBS 0.009712f
C860 B.n389 VSUBS 0.009712f
C861 B.n390 VSUBS 0.009712f
C862 B.n391 VSUBS 0.009712f
C863 B.n392 VSUBS 0.009712f
C864 B.n393 VSUBS 0.009712f
C865 B.n394 VSUBS 0.009712f
C866 B.n395 VSUBS 0.009712f
C867 B.n396 VSUBS 0.009712f
C868 B.n397 VSUBS 0.009712f
C869 B.n398 VSUBS 0.009712f
C870 B.n399 VSUBS 0.009712f
C871 B.n400 VSUBS 0.009712f
C872 B.n401 VSUBS 0.009712f
C873 B.n402 VSUBS 0.009712f
C874 B.n403 VSUBS 0.009712f
C875 B.n404 VSUBS 0.009712f
C876 B.n405 VSUBS 0.009712f
C877 B.n406 VSUBS 0.009712f
C878 B.n407 VSUBS 0.009712f
C879 B.n408 VSUBS 0.009712f
C880 B.n409 VSUBS 0.009712f
C881 B.n410 VSUBS 0.009712f
C882 B.n411 VSUBS 0.009712f
C883 B.n412 VSUBS 0.009712f
C884 B.n413 VSUBS 0.009712f
C885 B.n414 VSUBS 0.009712f
C886 B.n415 VSUBS 0.009712f
C887 B.n416 VSUBS 0.009712f
C888 B.n417 VSUBS 0.009712f
C889 B.n418 VSUBS 0.009712f
C890 B.n419 VSUBS 0.009712f
C891 B.n420 VSUBS 0.009712f
C892 B.n421 VSUBS 0.009712f
C893 B.n422 VSUBS 0.009712f
C894 B.n423 VSUBS 0.009712f
C895 B.n424 VSUBS 0.009712f
C896 B.n425 VSUBS 0.009712f
C897 B.n426 VSUBS 0.009712f
C898 B.n427 VSUBS 0.009712f
C899 B.n428 VSUBS 0.009712f
C900 B.n429 VSUBS 0.009712f
C901 B.n430 VSUBS 0.009712f
C902 B.n431 VSUBS 0.009712f
C903 B.n432 VSUBS 0.009712f
C904 B.n433 VSUBS 0.009712f
C905 B.n434 VSUBS 0.009712f
C906 B.n435 VSUBS 0.009712f
C907 B.n436 VSUBS 0.009712f
C908 B.n437 VSUBS 0.009712f
C909 B.n438 VSUBS 0.009712f
C910 B.n439 VSUBS 0.009712f
C911 B.n440 VSUBS 0.009712f
C912 B.n441 VSUBS 0.009712f
C913 B.n442 VSUBS 0.009712f
C914 B.n443 VSUBS 0.009712f
C915 B.n444 VSUBS 0.009712f
C916 B.n445 VSUBS 0.009712f
C917 B.n446 VSUBS 0.009712f
C918 B.n447 VSUBS 0.009712f
C919 B.n448 VSUBS 0.009712f
C920 B.n449 VSUBS 0.009712f
C921 B.n450 VSUBS 0.009712f
C922 B.n451 VSUBS 0.009712f
C923 B.n452 VSUBS 0.009712f
C924 B.n453 VSUBS 0.009712f
C925 B.n454 VSUBS 0.009712f
C926 B.n455 VSUBS 0.009712f
C927 B.n456 VSUBS 0.009712f
C928 B.n457 VSUBS 0.009712f
C929 B.n458 VSUBS 0.009712f
C930 B.n459 VSUBS 0.009712f
C931 B.n460 VSUBS 0.009712f
C932 B.n461 VSUBS 0.009712f
C933 B.n462 VSUBS 0.009712f
C934 B.n463 VSUBS 0.009712f
C935 B.n464 VSUBS 0.009712f
C936 B.n465 VSUBS 0.009712f
C937 B.n466 VSUBS 0.009712f
C938 B.n467 VSUBS 0.009712f
C939 B.n468 VSUBS 0.009712f
C940 B.n469 VSUBS 0.009712f
C941 B.n470 VSUBS 0.009712f
C942 B.n471 VSUBS 0.009712f
C943 B.n472 VSUBS 0.009712f
C944 B.n473 VSUBS 0.009712f
C945 B.n474 VSUBS 0.009712f
C946 B.n475 VSUBS 0.009712f
C947 B.n476 VSUBS 0.009712f
C948 B.n477 VSUBS 0.009712f
C949 B.n478 VSUBS 0.009712f
C950 B.n479 VSUBS 0.009712f
C951 B.n480 VSUBS 0.009712f
C952 B.n481 VSUBS 0.009712f
C953 B.n482 VSUBS 0.009712f
C954 B.n483 VSUBS 0.009712f
C955 B.n484 VSUBS 0.009712f
C956 B.n485 VSUBS 0.009712f
C957 B.n486 VSUBS 0.009712f
C958 B.n487 VSUBS 0.009712f
C959 B.n488 VSUBS 0.009712f
C960 B.n489 VSUBS 0.009712f
C961 B.n490 VSUBS 0.009712f
C962 B.n491 VSUBS 0.009712f
C963 B.n492 VSUBS 0.009712f
C964 B.n493 VSUBS 0.009712f
C965 B.n494 VSUBS 0.009712f
C966 B.n495 VSUBS 0.009712f
C967 B.n496 VSUBS 0.009712f
C968 B.n497 VSUBS 0.009712f
C969 B.n498 VSUBS 0.009712f
C970 B.n499 VSUBS 0.009712f
C971 B.n500 VSUBS 0.009712f
C972 B.n501 VSUBS 0.009712f
C973 B.n502 VSUBS 0.009712f
C974 B.n503 VSUBS 0.009712f
C975 B.n504 VSUBS 0.009712f
C976 B.n505 VSUBS 0.009712f
C977 B.n506 VSUBS 0.009712f
C978 B.n507 VSUBS 0.009712f
C979 B.n508 VSUBS 0.009712f
C980 B.n509 VSUBS 0.009712f
C981 B.n510 VSUBS 0.009712f
C982 B.n511 VSUBS 0.009712f
C983 B.n512 VSUBS 0.009712f
C984 B.n513 VSUBS 0.009712f
C985 B.n514 VSUBS 0.009712f
C986 B.n515 VSUBS 0.009712f
C987 B.n516 VSUBS 0.009712f
C988 B.n517 VSUBS 0.009712f
C989 B.n518 VSUBS 0.009712f
C990 B.n519 VSUBS 0.009712f
C991 B.n520 VSUBS 0.009712f
C992 B.n521 VSUBS 0.009712f
C993 B.n522 VSUBS 0.009712f
C994 B.n523 VSUBS 0.009712f
C995 B.n524 VSUBS 0.009712f
C996 B.n525 VSUBS 0.009712f
C997 B.n526 VSUBS 0.009712f
C998 B.n527 VSUBS 0.009712f
C999 B.n528 VSUBS 0.009712f
C1000 B.n529 VSUBS 0.009712f
C1001 B.n530 VSUBS 0.022145f
C1002 B.n531 VSUBS 0.020888f
C1003 B.n532 VSUBS 0.021961f
C1004 B.n533 VSUBS 0.009712f
C1005 B.n534 VSUBS 0.009712f
C1006 B.n535 VSUBS 0.009712f
C1007 B.n536 VSUBS 0.009712f
C1008 B.n537 VSUBS 0.009712f
C1009 B.n538 VSUBS 0.009712f
C1010 B.n539 VSUBS 0.009712f
C1011 B.n540 VSUBS 0.009712f
C1012 B.n541 VSUBS 0.009712f
C1013 B.n542 VSUBS 0.009712f
C1014 B.n543 VSUBS 0.009712f
C1015 B.n544 VSUBS 0.009712f
C1016 B.n545 VSUBS 0.009712f
C1017 B.n546 VSUBS 0.009712f
C1018 B.n547 VSUBS 0.009712f
C1019 B.n548 VSUBS 0.009712f
C1020 B.n549 VSUBS 0.009712f
C1021 B.n550 VSUBS 0.009712f
C1022 B.n551 VSUBS 0.009712f
C1023 B.n552 VSUBS 0.009712f
C1024 B.n553 VSUBS 0.009712f
C1025 B.n554 VSUBS 0.009712f
C1026 B.n555 VSUBS 0.009712f
C1027 B.n556 VSUBS 0.009712f
C1028 B.n557 VSUBS 0.009712f
C1029 B.n558 VSUBS 0.009712f
C1030 B.n559 VSUBS 0.009712f
C1031 B.n560 VSUBS 0.009712f
C1032 B.n561 VSUBS 0.009712f
C1033 B.n562 VSUBS 0.009712f
C1034 B.n563 VSUBS 0.009712f
C1035 B.n564 VSUBS 0.009141f
C1036 B.n565 VSUBS 0.022502f
C1037 B.n566 VSUBS 0.005427f
C1038 B.n567 VSUBS 0.009712f
C1039 B.n568 VSUBS 0.009712f
C1040 B.n569 VSUBS 0.009712f
C1041 B.n570 VSUBS 0.009712f
C1042 B.n571 VSUBS 0.009712f
C1043 B.n572 VSUBS 0.009712f
C1044 B.n573 VSUBS 0.009712f
C1045 B.n574 VSUBS 0.009712f
C1046 B.n575 VSUBS 0.009712f
C1047 B.n576 VSUBS 0.009712f
C1048 B.n577 VSUBS 0.009712f
C1049 B.n578 VSUBS 0.009712f
C1050 B.n579 VSUBS 0.005427f
C1051 B.n580 VSUBS 0.009712f
C1052 B.n581 VSUBS 0.009712f
C1053 B.n582 VSUBS 0.009712f
C1054 B.n583 VSUBS 0.009712f
C1055 B.n584 VSUBS 0.009712f
C1056 B.n585 VSUBS 0.009712f
C1057 B.n586 VSUBS 0.009712f
C1058 B.n587 VSUBS 0.009712f
C1059 B.n588 VSUBS 0.009712f
C1060 B.n589 VSUBS 0.009712f
C1061 B.n590 VSUBS 0.009712f
C1062 B.n591 VSUBS 0.009712f
C1063 B.n592 VSUBS 0.009712f
C1064 B.n593 VSUBS 0.009712f
C1065 B.n594 VSUBS 0.009712f
C1066 B.n595 VSUBS 0.009712f
C1067 B.n596 VSUBS 0.009712f
C1068 B.n597 VSUBS 0.009712f
C1069 B.n598 VSUBS 0.009712f
C1070 B.n599 VSUBS 0.009712f
C1071 B.n600 VSUBS 0.009712f
C1072 B.n601 VSUBS 0.009712f
C1073 B.n602 VSUBS 0.009712f
C1074 B.n603 VSUBS 0.009712f
C1075 B.n604 VSUBS 0.009712f
C1076 B.n605 VSUBS 0.009712f
C1077 B.n606 VSUBS 0.009712f
C1078 B.n607 VSUBS 0.009712f
C1079 B.n608 VSUBS 0.009712f
C1080 B.n609 VSUBS 0.009712f
C1081 B.n610 VSUBS 0.009712f
C1082 B.n611 VSUBS 0.009712f
C1083 B.n612 VSUBS 0.021961f
C1084 B.n613 VSUBS 0.021961f
C1085 B.n614 VSUBS 0.020888f
C1086 B.n615 VSUBS 0.009712f
C1087 B.n616 VSUBS 0.009712f
C1088 B.n617 VSUBS 0.009712f
C1089 B.n618 VSUBS 0.009712f
C1090 B.n619 VSUBS 0.009712f
C1091 B.n620 VSUBS 0.009712f
C1092 B.n621 VSUBS 0.009712f
C1093 B.n622 VSUBS 0.009712f
C1094 B.n623 VSUBS 0.009712f
C1095 B.n624 VSUBS 0.009712f
C1096 B.n625 VSUBS 0.009712f
C1097 B.n626 VSUBS 0.009712f
C1098 B.n627 VSUBS 0.009712f
C1099 B.n628 VSUBS 0.009712f
C1100 B.n629 VSUBS 0.009712f
C1101 B.n630 VSUBS 0.009712f
C1102 B.n631 VSUBS 0.009712f
C1103 B.n632 VSUBS 0.009712f
C1104 B.n633 VSUBS 0.009712f
C1105 B.n634 VSUBS 0.009712f
C1106 B.n635 VSUBS 0.009712f
C1107 B.n636 VSUBS 0.009712f
C1108 B.n637 VSUBS 0.009712f
C1109 B.n638 VSUBS 0.009712f
C1110 B.n639 VSUBS 0.009712f
C1111 B.n640 VSUBS 0.009712f
C1112 B.n641 VSUBS 0.009712f
C1113 B.n642 VSUBS 0.009712f
C1114 B.n643 VSUBS 0.009712f
C1115 B.n644 VSUBS 0.009712f
C1116 B.n645 VSUBS 0.009712f
C1117 B.n646 VSUBS 0.009712f
C1118 B.n647 VSUBS 0.009712f
C1119 B.n648 VSUBS 0.009712f
C1120 B.n649 VSUBS 0.009712f
C1121 B.n650 VSUBS 0.009712f
C1122 B.n651 VSUBS 0.009712f
C1123 B.n652 VSUBS 0.009712f
C1124 B.n653 VSUBS 0.009712f
C1125 B.n654 VSUBS 0.009712f
C1126 B.n655 VSUBS 0.009712f
C1127 B.n656 VSUBS 0.009712f
C1128 B.n657 VSUBS 0.009712f
C1129 B.n658 VSUBS 0.009712f
C1130 B.n659 VSUBS 0.009712f
C1131 B.n660 VSUBS 0.009712f
C1132 B.n661 VSUBS 0.009712f
C1133 B.n662 VSUBS 0.009712f
C1134 B.n663 VSUBS 0.009712f
C1135 B.n664 VSUBS 0.009712f
C1136 B.n665 VSUBS 0.009712f
C1137 B.n666 VSUBS 0.009712f
C1138 B.n667 VSUBS 0.009712f
C1139 B.n668 VSUBS 0.009712f
C1140 B.n669 VSUBS 0.009712f
C1141 B.n670 VSUBS 0.009712f
C1142 B.n671 VSUBS 0.009712f
C1143 B.n672 VSUBS 0.009712f
C1144 B.n673 VSUBS 0.009712f
C1145 B.n674 VSUBS 0.009712f
C1146 B.n675 VSUBS 0.009712f
C1147 B.n676 VSUBS 0.009712f
C1148 B.n677 VSUBS 0.009712f
C1149 B.n678 VSUBS 0.009712f
C1150 B.n679 VSUBS 0.009712f
C1151 B.n680 VSUBS 0.009712f
C1152 B.n681 VSUBS 0.009712f
C1153 B.n682 VSUBS 0.009712f
C1154 B.n683 VSUBS 0.009712f
C1155 B.n684 VSUBS 0.009712f
C1156 B.n685 VSUBS 0.009712f
C1157 B.n686 VSUBS 0.009712f
C1158 B.n687 VSUBS 0.009712f
C1159 B.n688 VSUBS 0.009712f
C1160 B.n689 VSUBS 0.009712f
C1161 B.n690 VSUBS 0.009712f
C1162 B.n691 VSUBS 0.009712f
C1163 B.n692 VSUBS 0.009712f
C1164 B.n693 VSUBS 0.009712f
C1165 B.n694 VSUBS 0.009712f
C1166 B.n695 VSUBS 0.009712f
C1167 B.n696 VSUBS 0.009712f
C1168 B.n697 VSUBS 0.009712f
C1169 B.n698 VSUBS 0.009712f
C1170 B.n699 VSUBS 0.009712f
C1171 B.n700 VSUBS 0.009712f
C1172 B.n701 VSUBS 0.009712f
C1173 B.n702 VSUBS 0.009712f
C1174 B.n703 VSUBS 0.021992f
.ends

