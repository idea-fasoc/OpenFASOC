* NGSPICE file created from diff_pair_sample_1510.ext - technology: sky130A

.subckt diff_pair_sample_1510 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=1.7292 ps=10.81 w=10.48 l=2.55
X1 VDD1.t9 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=4.0872 ps=21.74 w=10.48 l=2.55
X2 VTAIL.t9 VP.t1 VDD1.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X3 VDD2.t8 VN.t1 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=1.7292 ps=10.81 w=10.48 l=2.55
X4 VTAIL.t10 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X5 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=4.0872 ps=21.74 w=10.48 l=2.55
X6 VDD1.t6 VP.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X7 VTAIL.t12 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X8 VDD2.t5 VN.t4 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X9 VTAIL.t19 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X10 VDD2.t3 VN.t6 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X11 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=0 ps=0 w=10.48 l=2.55
X12 VTAIL.t8 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X13 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=0 ps=0 w=10.48 l=2.55
X14 VDD2.t2 VN.t7 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=4.0872 ps=21.74 w=10.48 l=2.55
X15 VDD2.t1 VN.t8 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=4.0872 ps=21.74 w=10.48 l=2.55
X16 VTAIL.t16 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X17 VDD1.t4 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X18 VTAIL.t3 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X19 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=1.7292 ps=10.81 w=10.48 l=2.55
X20 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=0 ps=0 w=10.48 l=2.55
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=0 ps=0 w=10.48 l=2.55
X22 VTAIL.t6 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7292 pd=10.81 as=1.7292 ps=10.81 w=10.48 l=2.55
X23 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.0872 pd=21.74 as=1.7292 ps=10.81 w=10.48 l=2.55
R0 VN.n75 VN.n39 161.3
R1 VN.n74 VN.n73 161.3
R2 VN.n72 VN.n40 161.3
R3 VN.n71 VN.n70 161.3
R4 VN.n69 VN.n41 161.3
R5 VN.n68 VN.n67 161.3
R6 VN.n66 VN.n65 161.3
R7 VN.n64 VN.n43 161.3
R8 VN.n63 VN.n62 161.3
R9 VN.n61 VN.n44 161.3
R10 VN.n60 VN.n59 161.3
R11 VN.n58 VN.n45 161.3
R12 VN.n57 VN.n56 161.3
R13 VN.n55 VN.n46 161.3
R14 VN.n54 VN.n53 161.3
R15 VN.n52 VN.n47 161.3
R16 VN.n51 VN.n50 161.3
R17 VN.n36 VN.n0 161.3
R18 VN.n35 VN.n34 161.3
R19 VN.n33 VN.n1 161.3
R20 VN.n32 VN.n31 161.3
R21 VN.n30 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n26 161.3
R24 VN.n25 VN.n4 161.3
R25 VN.n24 VN.n23 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n10 VN.t0 133.29
R35 VN.n49 VN.t8 133.29
R36 VN.n19 VN.t6 99.0468
R37 VN.n9 VN.t2 99.0468
R38 VN.n3 VN.t3 99.0468
R39 VN.n37 VN.t7 99.0468
R40 VN.n58 VN.t4 99.0468
R41 VN.n48 VN.t9 99.0468
R42 VN.n42 VN.t5 99.0468
R43 VN.n76 VN.t1 99.0468
R44 VN.n38 VN.n37 97.9476
R45 VN.n77 VN.n76 97.9476
R46 VN.n31 VN.n1 56.4773
R47 VN.n70 VN.n40 56.4773
R48 VN.n10 VN.n9 53.8957
R49 VN.n49 VN.n48 53.8957
R50 VN VN.n77 52.0208
R51 VN.n14 VN.n7 46.253
R52 VN.n24 VN.n5 46.253
R53 VN.n53 VN.n46 46.253
R54 VN.n63 VN.n44 46.253
R55 VN.n14 VN.n13 34.5682
R56 VN.n25 VN.n24 34.5682
R57 VN.n53 VN.n52 34.5682
R58 VN.n64 VN.n63 34.5682
R59 VN.n13 VN.n12 24.3439
R60 VN.n18 VN.n7 24.3439
R61 VN.n19 VN.n18 24.3439
R62 VN.n20 VN.n19 24.3439
R63 VN.n20 VN.n5 24.3439
R64 VN.n26 VN.n25 24.3439
R65 VN.n30 VN.n29 24.3439
R66 VN.n31 VN.n30 24.3439
R67 VN.n35 VN.n1 24.3439
R68 VN.n36 VN.n35 24.3439
R69 VN.n52 VN.n51 24.3439
R70 VN.n59 VN.n44 24.3439
R71 VN.n59 VN.n58 24.3439
R72 VN.n58 VN.n57 24.3439
R73 VN.n57 VN.n46 24.3439
R74 VN.n70 VN.n69 24.3439
R75 VN.n69 VN.n68 24.3439
R76 VN.n65 VN.n64 24.3439
R77 VN.n75 VN.n74 24.3439
R78 VN.n74 VN.n40 24.3439
R79 VN.n12 VN.n9 18.5015
R80 VN.n26 VN.n3 18.5015
R81 VN.n51 VN.n48 18.5015
R82 VN.n65 VN.n42 18.5015
R83 VN.n37 VN.n36 12.6591
R84 VN.n76 VN.n75 12.6591
R85 VN.n50 VN.n49 6.69845
R86 VN.n11 VN.n10 6.69845
R87 VN.n29 VN.n3 5.84292
R88 VN.n68 VN.n42 5.84292
R89 VN.n77 VN.n39 0.278398
R90 VN.n38 VN.n0 0.278398
R91 VN.n73 VN.n39 0.189894
R92 VN.n73 VN.n72 0.189894
R93 VN.n72 VN.n71 0.189894
R94 VN.n71 VN.n41 0.189894
R95 VN.n67 VN.n41 0.189894
R96 VN.n67 VN.n66 0.189894
R97 VN.n66 VN.n43 0.189894
R98 VN.n62 VN.n43 0.189894
R99 VN.n62 VN.n61 0.189894
R100 VN.n61 VN.n60 0.189894
R101 VN.n60 VN.n45 0.189894
R102 VN.n56 VN.n45 0.189894
R103 VN.n56 VN.n55 0.189894
R104 VN.n55 VN.n54 0.189894
R105 VN.n54 VN.n47 0.189894
R106 VN.n50 VN.n47 0.189894
R107 VN.n11 VN.n8 0.189894
R108 VN.n15 VN.n8 0.189894
R109 VN.n16 VN.n15 0.189894
R110 VN.n17 VN.n16 0.189894
R111 VN.n17 VN.n6 0.189894
R112 VN.n21 VN.n6 0.189894
R113 VN.n22 VN.n21 0.189894
R114 VN.n23 VN.n22 0.189894
R115 VN.n23 VN.n4 0.189894
R116 VN.n27 VN.n4 0.189894
R117 VN.n28 VN.n27 0.189894
R118 VN.n28 VN.n2 0.189894
R119 VN.n32 VN.n2 0.189894
R120 VN.n33 VN.n32 0.189894
R121 VN.n34 VN.n33 0.189894
R122 VN.n34 VN.n0 0.189894
R123 VN VN.n38 0.153422
R124 VTAIL.n11 VTAIL.t15 50.7966
R125 VTAIL.n17 VTAIL.t11 50.7963
R126 VTAIL.n2 VTAIL.t2 50.7963
R127 VTAIL.n16 VTAIL.t4 50.7963
R128 VTAIL.n15 VTAIL.n14 48.9072
R129 VTAIL.n13 VTAIL.n12 48.9072
R130 VTAIL.n10 VTAIL.n9 48.9072
R131 VTAIL.n8 VTAIL.n7 48.9072
R132 VTAIL.n19 VTAIL.n18 48.907
R133 VTAIL.n1 VTAIL.n0 48.907
R134 VTAIL.n4 VTAIL.n3 48.907
R135 VTAIL.n6 VTAIL.n5 48.907
R136 VTAIL.n8 VTAIL.n6 26.3669
R137 VTAIL.n17 VTAIL.n16 23.8841
R138 VTAIL.n10 VTAIL.n8 2.48326
R139 VTAIL.n11 VTAIL.n10 2.48326
R140 VTAIL.n15 VTAIL.n13 2.48326
R141 VTAIL.n16 VTAIL.n15 2.48326
R142 VTAIL.n6 VTAIL.n4 2.48326
R143 VTAIL.n4 VTAIL.n2 2.48326
R144 VTAIL.n19 VTAIL.n17 2.48326
R145 VTAIL VTAIL.n1 1.92076
R146 VTAIL.n18 VTAIL.t14 1.88981
R147 VTAIL.n18 VTAIL.t12 1.88981
R148 VTAIL.n0 VTAIL.t13 1.88981
R149 VTAIL.n0 VTAIL.t10 1.88981
R150 VTAIL.n3 VTAIL.t7 1.88981
R151 VTAIL.n3 VTAIL.t6 1.88981
R152 VTAIL.n5 VTAIL.t0 1.88981
R153 VTAIL.n5 VTAIL.t8 1.88981
R154 VTAIL.n14 VTAIL.t5 1.88981
R155 VTAIL.n14 VTAIL.t9 1.88981
R156 VTAIL.n12 VTAIL.t1 1.88981
R157 VTAIL.n12 VTAIL.t3 1.88981
R158 VTAIL.n9 VTAIL.t18 1.88981
R159 VTAIL.n9 VTAIL.t16 1.88981
R160 VTAIL.n7 VTAIL.t17 1.88981
R161 VTAIL.n7 VTAIL.t19 1.88981
R162 VTAIL.n13 VTAIL.n11 1.71171
R163 VTAIL.n2 VTAIL.n1 1.71171
R164 VTAIL VTAIL.n19 0.563
R165 VDD2.n1 VDD2.t9 69.9579
R166 VDD2.n4 VDD2.t8 67.4753
R167 VDD2.n3 VDD2.n2 67.3925
R168 VDD2 VDD2.n7 67.3897
R169 VDD2.n6 VDD2.n5 65.586
R170 VDD2.n1 VDD2.n0 65.5858
R171 VDD2.n4 VDD2.n3 44.5429
R172 VDD2.n6 VDD2.n4 2.48326
R173 VDD2.n7 VDD2.t0 1.88981
R174 VDD2.n7 VDD2.t1 1.88981
R175 VDD2.n5 VDD2.t4 1.88981
R176 VDD2.n5 VDD2.t5 1.88981
R177 VDD2.n2 VDD2.t6 1.88981
R178 VDD2.n2 VDD2.t2 1.88981
R179 VDD2.n0 VDD2.t7 1.88981
R180 VDD2.n0 VDD2.t3 1.88981
R181 VDD2 VDD2.n6 0.679379
R182 VDD2.n3 VDD2.n1 0.565844
R183 B.n902 B.n901 585
R184 B.n318 B.n150 585
R185 B.n317 B.n316 585
R186 B.n315 B.n314 585
R187 B.n313 B.n312 585
R188 B.n311 B.n310 585
R189 B.n309 B.n308 585
R190 B.n307 B.n306 585
R191 B.n305 B.n304 585
R192 B.n303 B.n302 585
R193 B.n301 B.n300 585
R194 B.n299 B.n298 585
R195 B.n297 B.n296 585
R196 B.n295 B.n294 585
R197 B.n293 B.n292 585
R198 B.n291 B.n290 585
R199 B.n289 B.n288 585
R200 B.n287 B.n286 585
R201 B.n285 B.n284 585
R202 B.n283 B.n282 585
R203 B.n281 B.n280 585
R204 B.n279 B.n278 585
R205 B.n277 B.n276 585
R206 B.n275 B.n274 585
R207 B.n273 B.n272 585
R208 B.n271 B.n270 585
R209 B.n269 B.n268 585
R210 B.n267 B.n266 585
R211 B.n265 B.n264 585
R212 B.n263 B.n262 585
R213 B.n261 B.n260 585
R214 B.n259 B.n258 585
R215 B.n257 B.n256 585
R216 B.n255 B.n254 585
R217 B.n253 B.n252 585
R218 B.n251 B.n250 585
R219 B.n249 B.n248 585
R220 B.n246 B.n245 585
R221 B.n244 B.n243 585
R222 B.n242 B.n241 585
R223 B.n240 B.n239 585
R224 B.n238 B.n237 585
R225 B.n236 B.n235 585
R226 B.n234 B.n233 585
R227 B.n232 B.n231 585
R228 B.n230 B.n229 585
R229 B.n228 B.n227 585
R230 B.n225 B.n224 585
R231 B.n223 B.n222 585
R232 B.n221 B.n220 585
R233 B.n219 B.n218 585
R234 B.n217 B.n216 585
R235 B.n215 B.n214 585
R236 B.n213 B.n212 585
R237 B.n211 B.n210 585
R238 B.n209 B.n208 585
R239 B.n207 B.n206 585
R240 B.n205 B.n204 585
R241 B.n203 B.n202 585
R242 B.n201 B.n200 585
R243 B.n199 B.n198 585
R244 B.n197 B.n196 585
R245 B.n195 B.n194 585
R246 B.n193 B.n192 585
R247 B.n191 B.n190 585
R248 B.n189 B.n188 585
R249 B.n187 B.n186 585
R250 B.n185 B.n184 585
R251 B.n183 B.n182 585
R252 B.n181 B.n180 585
R253 B.n179 B.n178 585
R254 B.n177 B.n176 585
R255 B.n175 B.n174 585
R256 B.n173 B.n172 585
R257 B.n171 B.n170 585
R258 B.n169 B.n168 585
R259 B.n167 B.n166 585
R260 B.n165 B.n164 585
R261 B.n163 B.n162 585
R262 B.n161 B.n160 585
R263 B.n159 B.n158 585
R264 B.n157 B.n156 585
R265 B.n109 B.n108 585
R266 B.n907 B.n906 585
R267 B.n900 B.n151 585
R268 B.n151 B.n106 585
R269 B.n899 B.n105 585
R270 B.n911 B.n105 585
R271 B.n898 B.n104 585
R272 B.n912 B.n104 585
R273 B.n897 B.n103 585
R274 B.n913 B.n103 585
R275 B.n896 B.n895 585
R276 B.n895 B.n99 585
R277 B.n894 B.n98 585
R278 B.n919 B.n98 585
R279 B.n893 B.n97 585
R280 B.n920 B.n97 585
R281 B.n892 B.n96 585
R282 B.n921 B.n96 585
R283 B.n891 B.n890 585
R284 B.n890 B.n92 585
R285 B.n889 B.n91 585
R286 B.n927 B.n91 585
R287 B.n888 B.n90 585
R288 B.n928 B.n90 585
R289 B.n887 B.n89 585
R290 B.n929 B.n89 585
R291 B.n886 B.n885 585
R292 B.n885 B.n85 585
R293 B.n884 B.n84 585
R294 B.n935 B.n84 585
R295 B.n883 B.n83 585
R296 B.n936 B.n83 585
R297 B.n882 B.n82 585
R298 B.n937 B.n82 585
R299 B.n881 B.n880 585
R300 B.n880 B.n78 585
R301 B.n879 B.n77 585
R302 B.n943 B.n77 585
R303 B.n878 B.n76 585
R304 B.n944 B.n76 585
R305 B.n877 B.n75 585
R306 B.n945 B.n75 585
R307 B.n876 B.n875 585
R308 B.n875 B.n71 585
R309 B.n874 B.n70 585
R310 B.n951 B.n70 585
R311 B.n873 B.n69 585
R312 B.n952 B.n69 585
R313 B.n872 B.n68 585
R314 B.n953 B.n68 585
R315 B.n871 B.n870 585
R316 B.n870 B.n64 585
R317 B.n869 B.n63 585
R318 B.n959 B.n63 585
R319 B.n868 B.n62 585
R320 B.n960 B.n62 585
R321 B.n867 B.n61 585
R322 B.n961 B.n61 585
R323 B.n866 B.n865 585
R324 B.n865 B.n57 585
R325 B.n864 B.n56 585
R326 B.n967 B.n56 585
R327 B.n863 B.n55 585
R328 B.n968 B.n55 585
R329 B.n862 B.n54 585
R330 B.n969 B.n54 585
R331 B.n861 B.n860 585
R332 B.n860 B.n50 585
R333 B.n859 B.n49 585
R334 B.n975 B.n49 585
R335 B.n858 B.n48 585
R336 B.n976 B.n48 585
R337 B.n857 B.n47 585
R338 B.n977 B.n47 585
R339 B.n856 B.n855 585
R340 B.n855 B.n46 585
R341 B.n854 B.n42 585
R342 B.n983 B.n42 585
R343 B.n853 B.n41 585
R344 B.n984 B.n41 585
R345 B.n852 B.n40 585
R346 B.n985 B.n40 585
R347 B.n851 B.n850 585
R348 B.n850 B.n36 585
R349 B.n849 B.n35 585
R350 B.n991 B.n35 585
R351 B.n848 B.n34 585
R352 B.n992 B.n34 585
R353 B.n847 B.n33 585
R354 B.n993 B.n33 585
R355 B.n846 B.n845 585
R356 B.n845 B.n32 585
R357 B.n844 B.n28 585
R358 B.n999 B.n28 585
R359 B.n843 B.n27 585
R360 B.n1000 B.n27 585
R361 B.n842 B.n26 585
R362 B.n1001 B.n26 585
R363 B.n841 B.n840 585
R364 B.n840 B.n22 585
R365 B.n839 B.n21 585
R366 B.n1007 B.n21 585
R367 B.n838 B.n20 585
R368 B.n1008 B.n20 585
R369 B.n837 B.n19 585
R370 B.n1009 B.n19 585
R371 B.n836 B.n835 585
R372 B.n835 B.n15 585
R373 B.n834 B.n14 585
R374 B.n1015 B.n14 585
R375 B.n833 B.n13 585
R376 B.n1016 B.n13 585
R377 B.n832 B.n12 585
R378 B.n1017 B.n12 585
R379 B.n831 B.n830 585
R380 B.n830 B.n8 585
R381 B.n829 B.n7 585
R382 B.n1023 B.n7 585
R383 B.n828 B.n6 585
R384 B.n1024 B.n6 585
R385 B.n827 B.n5 585
R386 B.n1025 B.n5 585
R387 B.n826 B.n825 585
R388 B.n825 B.n4 585
R389 B.n824 B.n319 585
R390 B.n824 B.n823 585
R391 B.n814 B.n320 585
R392 B.n321 B.n320 585
R393 B.n816 B.n815 585
R394 B.n817 B.n816 585
R395 B.n813 B.n326 585
R396 B.n326 B.n325 585
R397 B.n812 B.n811 585
R398 B.n811 B.n810 585
R399 B.n328 B.n327 585
R400 B.n329 B.n328 585
R401 B.n803 B.n802 585
R402 B.n804 B.n803 585
R403 B.n801 B.n334 585
R404 B.n334 B.n333 585
R405 B.n800 B.n799 585
R406 B.n799 B.n798 585
R407 B.n336 B.n335 585
R408 B.n337 B.n336 585
R409 B.n791 B.n790 585
R410 B.n792 B.n791 585
R411 B.n789 B.n342 585
R412 B.n342 B.n341 585
R413 B.n788 B.n787 585
R414 B.n787 B.n786 585
R415 B.n344 B.n343 585
R416 B.n779 B.n344 585
R417 B.n778 B.n777 585
R418 B.n780 B.n778 585
R419 B.n776 B.n349 585
R420 B.n349 B.n348 585
R421 B.n775 B.n774 585
R422 B.n774 B.n773 585
R423 B.n351 B.n350 585
R424 B.n352 B.n351 585
R425 B.n766 B.n765 585
R426 B.n767 B.n766 585
R427 B.n764 B.n357 585
R428 B.n357 B.n356 585
R429 B.n763 B.n762 585
R430 B.n762 B.n761 585
R431 B.n359 B.n358 585
R432 B.n754 B.n359 585
R433 B.n753 B.n752 585
R434 B.n755 B.n753 585
R435 B.n751 B.n364 585
R436 B.n364 B.n363 585
R437 B.n750 B.n749 585
R438 B.n749 B.n748 585
R439 B.n366 B.n365 585
R440 B.n367 B.n366 585
R441 B.n741 B.n740 585
R442 B.n742 B.n741 585
R443 B.n739 B.n372 585
R444 B.n372 B.n371 585
R445 B.n738 B.n737 585
R446 B.n737 B.n736 585
R447 B.n374 B.n373 585
R448 B.n375 B.n374 585
R449 B.n729 B.n728 585
R450 B.n730 B.n729 585
R451 B.n727 B.n380 585
R452 B.n380 B.n379 585
R453 B.n726 B.n725 585
R454 B.n725 B.n724 585
R455 B.n382 B.n381 585
R456 B.n383 B.n382 585
R457 B.n717 B.n716 585
R458 B.n718 B.n717 585
R459 B.n715 B.n388 585
R460 B.n388 B.n387 585
R461 B.n714 B.n713 585
R462 B.n713 B.n712 585
R463 B.n390 B.n389 585
R464 B.n391 B.n390 585
R465 B.n705 B.n704 585
R466 B.n706 B.n705 585
R467 B.n703 B.n396 585
R468 B.n396 B.n395 585
R469 B.n702 B.n701 585
R470 B.n701 B.n700 585
R471 B.n398 B.n397 585
R472 B.n399 B.n398 585
R473 B.n693 B.n692 585
R474 B.n694 B.n693 585
R475 B.n691 B.n404 585
R476 B.n404 B.n403 585
R477 B.n690 B.n689 585
R478 B.n689 B.n688 585
R479 B.n406 B.n405 585
R480 B.n407 B.n406 585
R481 B.n681 B.n680 585
R482 B.n682 B.n681 585
R483 B.n679 B.n412 585
R484 B.n412 B.n411 585
R485 B.n678 B.n677 585
R486 B.n677 B.n676 585
R487 B.n414 B.n413 585
R488 B.n415 B.n414 585
R489 B.n669 B.n668 585
R490 B.n670 B.n669 585
R491 B.n667 B.n420 585
R492 B.n420 B.n419 585
R493 B.n666 B.n665 585
R494 B.n665 B.n664 585
R495 B.n422 B.n421 585
R496 B.n423 B.n422 585
R497 B.n657 B.n656 585
R498 B.n658 B.n657 585
R499 B.n655 B.n428 585
R500 B.n428 B.n427 585
R501 B.n654 B.n653 585
R502 B.n653 B.n652 585
R503 B.n430 B.n429 585
R504 B.n431 B.n430 585
R505 B.n648 B.n647 585
R506 B.n434 B.n433 585
R507 B.n644 B.n643 585
R508 B.n645 B.n644 585
R509 B.n642 B.n476 585
R510 B.n641 B.n640 585
R511 B.n639 B.n638 585
R512 B.n637 B.n636 585
R513 B.n635 B.n634 585
R514 B.n633 B.n632 585
R515 B.n631 B.n630 585
R516 B.n629 B.n628 585
R517 B.n627 B.n626 585
R518 B.n625 B.n624 585
R519 B.n623 B.n622 585
R520 B.n621 B.n620 585
R521 B.n619 B.n618 585
R522 B.n617 B.n616 585
R523 B.n615 B.n614 585
R524 B.n613 B.n612 585
R525 B.n611 B.n610 585
R526 B.n609 B.n608 585
R527 B.n607 B.n606 585
R528 B.n605 B.n604 585
R529 B.n603 B.n602 585
R530 B.n601 B.n600 585
R531 B.n599 B.n598 585
R532 B.n597 B.n596 585
R533 B.n595 B.n594 585
R534 B.n593 B.n592 585
R535 B.n591 B.n590 585
R536 B.n589 B.n588 585
R537 B.n587 B.n586 585
R538 B.n585 B.n584 585
R539 B.n583 B.n582 585
R540 B.n581 B.n580 585
R541 B.n579 B.n578 585
R542 B.n577 B.n576 585
R543 B.n575 B.n574 585
R544 B.n573 B.n572 585
R545 B.n571 B.n570 585
R546 B.n569 B.n568 585
R547 B.n567 B.n566 585
R548 B.n565 B.n564 585
R549 B.n563 B.n562 585
R550 B.n561 B.n560 585
R551 B.n559 B.n558 585
R552 B.n557 B.n556 585
R553 B.n555 B.n554 585
R554 B.n553 B.n552 585
R555 B.n551 B.n550 585
R556 B.n549 B.n548 585
R557 B.n547 B.n546 585
R558 B.n545 B.n544 585
R559 B.n543 B.n542 585
R560 B.n541 B.n540 585
R561 B.n539 B.n538 585
R562 B.n537 B.n536 585
R563 B.n535 B.n534 585
R564 B.n533 B.n532 585
R565 B.n531 B.n530 585
R566 B.n529 B.n528 585
R567 B.n527 B.n526 585
R568 B.n525 B.n524 585
R569 B.n523 B.n522 585
R570 B.n521 B.n520 585
R571 B.n519 B.n518 585
R572 B.n517 B.n516 585
R573 B.n515 B.n514 585
R574 B.n513 B.n512 585
R575 B.n511 B.n510 585
R576 B.n509 B.n508 585
R577 B.n507 B.n506 585
R578 B.n505 B.n504 585
R579 B.n503 B.n502 585
R580 B.n501 B.n500 585
R581 B.n499 B.n498 585
R582 B.n497 B.n496 585
R583 B.n495 B.n494 585
R584 B.n493 B.n492 585
R585 B.n491 B.n490 585
R586 B.n489 B.n488 585
R587 B.n487 B.n486 585
R588 B.n485 B.n484 585
R589 B.n483 B.n475 585
R590 B.n645 B.n475 585
R591 B.n649 B.n432 585
R592 B.n432 B.n431 585
R593 B.n651 B.n650 585
R594 B.n652 B.n651 585
R595 B.n426 B.n425 585
R596 B.n427 B.n426 585
R597 B.n660 B.n659 585
R598 B.n659 B.n658 585
R599 B.n661 B.n424 585
R600 B.n424 B.n423 585
R601 B.n663 B.n662 585
R602 B.n664 B.n663 585
R603 B.n418 B.n417 585
R604 B.n419 B.n418 585
R605 B.n672 B.n671 585
R606 B.n671 B.n670 585
R607 B.n673 B.n416 585
R608 B.n416 B.n415 585
R609 B.n675 B.n674 585
R610 B.n676 B.n675 585
R611 B.n410 B.n409 585
R612 B.n411 B.n410 585
R613 B.n684 B.n683 585
R614 B.n683 B.n682 585
R615 B.n685 B.n408 585
R616 B.n408 B.n407 585
R617 B.n687 B.n686 585
R618 B.n688 B.n687 585
R619 B.n402 B.n401 585
R620 B.n403 B.n402 585
R621 B.n696 B.n695 585
R622 B.n695 B.n694 585
R623 B.n697 B.n400 585
R624 B.n400 B.n399 585
R625 B.n699 B.n698 585
R626 B.n700 B.n699 585
R627 B.n394 B.n393 585
R628 B.n395 B.n394 585
R629 B.n708 B.n707 585
R630 B.n707 B.n706 585
R631 B.n709 B.n392 585
R632 B.n392 B.n391 585
R633 B.n711 B.n710 585
R634 B.n712 B.n711 585
R635 B.n386 B.n385 585
R636 B.n387 B.n386 585
R637 B.n720 B.n719 585
R638 B.n719 B.n718 585
R639 B.n721 B.n384 585
R640 B.n384 B.n383 585
R641 B.n723 B.n722 585
R642 B.n724 B.n723 585
R643 B.n378 B.n377 585
R644 B.n379 B.n378 585
R645 B.n732 B.n731 585
R646 B.n731 B.n730 585
R647 B.n733 B.n376 585
R648 B.n376 B.n375 585
R649 B.n735 B.n734 585
R650 B.n736 B.n735 585
R651 B.n370 B.n369 585
R652 B.n371 B.n370 585
R653 B.n744 B.n743 585
R654 B.n743 B.n742 585
R655 B.n745 B.n368 585
R656 B.n368 B.n367 585
R657 B.n747 B.n746 585
R658 B.n748 B.n747 585
R659 B.n362 B.n361 585
R660 B.n363 B.n362 585
R661 B.n757 B.n756 585
R662 B.n756 B.n755 585
R663 B.n758 B.n360 585
R664 B.n754 B.n360 585
R665 B.n760 B.n759 585
R666 B.n761 B.n760 585
R667 B.n355 B.n354 585
R668 B.n356 B.n355 585
R669 B.n769 B.n768 585
R670 B.n768 B.n767 585
R671 B.n770 B.n353 585
R672 B.n353 B.n352 585
R673 B.n772 B.n771 585
R674 B.n773 B.n772 585
R675 B.n347 B.n346 585
R676 B.n348 B.n347 585
R677 B.n782 B.n781 585
R678 B.n781 B.n780 585
R679 B.n783 B.n345 585
R680 B.n779 B.n345 585
R681 B.n785 B.n784 585
R682 B.n786 B.n785 585
R683 B.n340 B.n339 585
R684 B.n341 B.n340 585
R685 B.n794 B.n793 585
R686 B.n793 B.n792 585
R687 B.n795 B.n338 585
R688 B.n338 B.n337 585
R689 B.n797 B.n796 585
R690 B.n798 B.n797 585
R691 B.n332 B.n331 585
R692 B.n333 B.n332 585
R693 B.n806 B.n805 585
R694 B.n805 B.n804 585
R695 B.n807 B.n330 585
R696 B.n330 B.n329 585
R697 B.n809 B.n808 585
R698 B.n810 B.n809 585
R699 B.n324 B.n323 585
R700 B.n325 B.n324 585
R701 B.n819 B.n818 585
R702 B.n818 B.n817 585
R703 B.n820 B.n322 585
R704 B.n322 B.n321 585
R705 B.n822 B.n821 585
R706 B.n823 B.n822 585
R707 B.n2 B.n0 585
R708 B.n4 B.n2 585
R709 B.n3 B.n1 585
R710 B.n1024 B.n3 585
R711 B.n1022 B.n1021 585
R712 B.n1023 B.n1022 585
R713 B.n1020 B.n9 585
R714 B.n9 B.n8 585
R715 B.n1019 B.n1018 585
R716 B.n1018 B.n1017 585
R717 B.n11 B.n10 585
R718 B.n1016 B.n11 585
R719 B.n1014 B.n1013 585
R720 B.n1015 B.n1014 585
R721 B.n1012 B.n16 585
R722 B.n16 B.n15 585
R723 B.n1011 B.n1010 585
R724 B.n1010 B.n1009 585
R725 B.n18 B.n17 585
R726 B.n1008 B.n18 585
R727 B.n1006 B.n1005 585
R728 B.n1007 B.n1006 585
R729 B.n1004 B.n23 585
R730 B.n23 B.n22 585
R731 B.n1003 B.n1002 585
R732 B.n1002 B.n1001 585
R733 B.n25 B.n24 585
R734 B.n1000 B.n25 585
R735 B.n998 B.n997 585
R736 B.n999 B.n998 585
R737 B.n996 B.n29 585
R738 B.n32 B.n29 585
R739 B.n995 B.n994 585
R740 B.n994 B.n993 585
R741 B.n31 B.n30 585
R742 B.n992 B.n31 585
R743 B.n990 B.n989 585
R744 B.n991 B.n990 585
R745 B.n988 B.n37 585
R746 B.n37 B.n36 585
R747 B.n987 B.n986 585
R748 B.n986 B.n985 585
R749 B.n39 B.n38 585
R750 B.n984 B.n39 585
R751 B.n982 B.n981 585
R752 B.n983 B.n982 585
R753 B.n980 B.n43 585
R754 B.n46 B.n43 585
R755 B.n979 B.n978 585
R756 B.n978 B.n977 585
R757 B.n45 B.n44 585
R758 B.n976 B.n45 585
R759 B.n974 B.n973 585
R760 B.n975 B.n974 585
R761 B.n972 B.n51 585
R762 B.n51 B.n50 585
R763 B.n971 B.n970 585
R764 B.n970 B.n969 585
R765 B.n53 B.n52 585
R766 B.n968 B.n53 585
R767 B.n966 B.n965 585
R768 B.n967 B.n966 585
R769 B.n964 B.n58 585
R770 B.n58 B.n57 585
R771 B.n963 B.n962 585
R772 B.n962 B.n961 585
R773 B.n60 B.n59 585
R774 B.n960 B.n60 585
R775 B.n958 B.n957 585
R776 B.n959 B.n958 585
R777 B.n956 B.n65 585
R778 B.n65 B.n64 585
R779 B.n955 B.n954 585
R780 B.n954 B.n953 585
R781 B.n67 B.n66 585
R782 B.n952 B.n67 585
R783 B.n950 B.n949 585
R784 B.n951 B.n950 585
R785 B.n948 B.n72 585
R786 B.n72 B.n71 585
R787 B.n947 B.n946 585
R788 B.n946 B.n945 585
R789 B.n74 B.n73 585
R790 B.n944 B.n74 585
R791 B.n942 B.n941 585
R792 B.n943 B.n942 585
R793 B.n940 B.n79 585
R794 B.n79 B.n78 585
R795 B.n939 B.n938 585
R796 B.n938 B.n937 585
R797 B.n81 B.n80 585
R798 B.n936 B.n81 585
R799 B.n934 B.n933 585
R800 B.n935 B.n934 585
R801 B.n932 B.n86 585
R802 B.n86 B.n85 585
R803 B.n931 B.n930 585
R804 B.n930 B.n929 585
R805 B.n88 B.n87 585
R806 B.n928 B.n88 585
R807 B.n926 B.n925 585
R808 B.n927 B.n926 585
R809 B.n924 B.n93 585
R810 B.n93 B.n92 585
R811 B.n923 B.n922 585
R812 B.n922 B.n921 585
R813 B.n95 B.n94 585
R814 B.n920 B.n95 585
R815 B.n918 B.n917 585
R816 B.n919 B.n918 585
R817 B.n916 B.n100 585
R818 B.n100 B.n99 585
R819 B.n915 B.n914 585
R820 B.n914 B.n913 585
R821 B.n102 B.n101 585
R822 B.n912 B.n102 585
R823 B.n910 B.n909 585
R824 B.n911 B.n910 585
R825 B.n908 B.n107 585
R826 B.n107 B.n106 585
R827 B.n1027 B.n1026 585
R828 B.n1026 B.n1025 585
R829 B.n647 B.n432 478.086
R830 B.n906 B.n107 478.086
R831 B.n475 B.n430 478.086
R832 B.n902 B.n151 478.086
R833 B.n480 B.t10 307.017
R834 B.n477 B.t21 307.017
R835 B.n154 B.t18 307.017
R836 B.n152 B.t14 307.017
R837 B.n904 B.n903 256.663
R838 B.n904 B.n149 256.663
R839 B.n904 B.n148 256.663
R840 B.n904 B.n147 256.663
R841 B.n904 B.n146 256.663
R842 B.n904 B.n145 256.663
R843 B.n904 B.n144 256.663
R844 B.n904 B.n143 256.663
R845 B.n904 B.n142 256.663
R846 B.n904 B.n141 256.663
R847 B.n904 B.n140 256.663
R848 B.n904 B.n139 256.663
R849 B.n904 B.n138 256.663
R850 B.n904 B.n137 256.663
R851 B.n904 B.n136 256.663
R852 B.n904 B.n135 256.663
R853 B.n904 B.n134 256.663
R854 B.n904 B.n133 256.663
R855 B.n904 B.n132 256.663
R856 B.n904 B.n131 256.663
R857 B.n904 B.n130 256.663
R858 B.n904 B.n129 256.663
R859 B.n904 B.n128 256.663
R860 B.n904 B.n127 256.663
R861 B.n904 B.n126 256.663
R862 B.n904 B.n125 256.663
R863 B.n904 B.n124 256.663
R864 B.n904 B.n123 256.663
R865 B.n904 B.n122 256.663
R866 B.n904 B.n121 256.663
R867 B.n904 B.n120 256.663
R868 B.n904 B.n119 256.663
R869 B.n904 B.n118 256.663
R870 B.n904 B.n117 256.663
R871 B.n904 B.n116 256.663
R872 B.n904 B.n115 256.663
R873 B.n904 B.n114 256.663
R874 B.n904 B.n113 256.663
R875 B.n904 B.n112 256.663
R876 B.n904 B.n111 256.663
R877 B.n904 B.n110 256.663
R878 B.n905 B.n904 256.663
R879 B.n646 B.n645 256.663
R880 B.n645 B.n435 256.663
R881 B.n645 B.n436 256.663
R882 B.n645 B.n437 256.663
R883 B.n645 B.n438 256.663
R884 B.n645 B.n439 256.663
R885 B.n645 B.n440 256.663
R886 B.n645 B.n441 256.663
R887 B.n645 B.n442 256.663
R888 B.n645 B.n443 256.663
R889 B.n645 B.n444 256.663
R890 B.n645 B.n445 256.663
R891 B.n645 B.n446 256.663
R892 B.n645 B.n447 256.663
R893 B.n645 B.n448 256.663
R894 B.n645 B.n449 256.663
R895 B.n645 B.n450 256.663
R896 B.n645 B.n451 256.663
R897 B.n645 B.n452 256.663
R898 B.n645 B.n453 256.663
R899 B.n645 B.n454 256.663
R900 B.n645 B.n455 256.663
R901 B.n645 B.n456 256.663
R902 B.n645 B.n457 256.663
R903 B.n645 B.n458 256.663
R904 B.n645 B.n459 256.663
R905 B.n645 B.n460 256.663
R906 B.n645 B.n461 256.663
R907 B.n645 B.n462 256.663
R908 B.n645 B.n463 256.663
R909 B.n645 B.n464 256.663
R910 B.n645 B.n465 256.663
R911 B.n645 B.n466 256.663
R912 B.n645 B.n467 256.663
R913 B.n645 B.n468 256.663
R914 B.n645 B.n469 256.663
R915 B.n645 B.n470 256.663
R916 B.n645 B.n471 256.663
R917 B.n645 B.n472 256.663
R918 B.n645 B.n473 256.663
R919 B.n645 B.n474 256.663
R920 B.n651 B.n432 163.367
R921 B.n651 B.n426 163.367
R922 B.n659 B.n426 163.367
R923 B.n659 B.n424 163.367
R924 B.n663 B.n424 163.367
R925 B.n663 B.n418 163.367
R926 B.n671 B.n418 163.367
R927 B.n671 B.n416 163.367
R928 B.n675 B.n416 163.367
R929 B.n675 B.n410 163.367
R930 B.n683 B.n410 163.367
R931 B.n683 B.n408 163.367
R932 B.n687 B.n408 163.367
R933 B.n687 B.n402 163.367
R934 B.n695 B.n402 163.367
R935 B.n695 B.n400 163.367
R936 B.n699 B.n400 163.367
R937 B.n699 B.n394 163.367
R938 B.n707 B.n394 163.367
R939 B.n707 B.n392 163.367
R940 B.n711 B.n392 163.367
R941 B.n711 B.n386 163.367
R942 B.n719 B.n386 163.367
R943 B.n719 B.n384 163.367
R944 B.n723 B.n384 163.367
R945 B.n723 B.n378 163.367
R946 B.n731 B.n378 163.367
R947 B.n731 B.n376 163.367
R948 B.n735 B.n376 163.367
R949 B.n735 B.n370 163.367
R950 B.n743 B.n370 163.367
R951 B.n743 B.n368 163.367
R952 B.n747 B.n368 163.367
R953 B.n747 B.n362 163.367
R954 B.n756 B.n362 163.367
R955 B.n756 B.n360 163.367
R956 B.n760 B.n360 163.367
R957 B.n760 B.n355 163.367
R958 B.n768 B.n355 163.367
R959 B.n768 B.n353 163.367
R960 B.n772 B.n353 163.367
R961 B.n772 B.n347 163.367
R962 B.n781 B.n347 163.367
R963 B.n781 B.n345 163.367
R964 B.n785 B.n345 163.367
R965 B.n785 B.n340 163.367
R966 B.n793 B.n340 163.367
R967 B.n793 B.n338 163.367
R968 B.n797 B.n338 163.367
R969 B.n797 B.n332 163.367
R970 B.n805 B.n332 163.367
R971 B.n805 B.n330 163.367
R972 B.n809 B.n330 163.367
R973 B.n809 B.n324 163.367
R974 B.n818 B.n324 163.367
R975 B.n818 B.n322 163.367
R976 B.n822 B.n322 163.367
R977 B.n822 B.n2 163.367
R978 B.n1026 B.n2 163.367
R979 B.n1026 B.n3 163.367
R980 B.n1022 B.n3 163.367
R981 B.n1022 B.n9 163.367
R982 B.n1018 B.n9 163.367
R983 B.n1018 B.n11 163.367
R984 B.n1014 B.n11 163.367
R985 B.n1014 B.n16 163.367
R986 B.n1010 B.n16 163.367
R987 B.n1010 B.n18 163.367
R988 B.n1006 B.n18 163.367
R989 B.n1006 B.n23 163.367
R990 B.n1002 B.n23 163.367
R991 B.n1002 B.n25 163.367
R992 B.n998 B.n25 163.367
R993 B.n998 B.n29 163.367
R994 B.n994 B.n29 163.367
R995 B.n994 B.n31 163.367
R996 B.n990 B.n31 163.367
R997 B.n990 B.n37 163.367
R998 B.n986 B.n37 163.367
R999 B.n986 B.n39 163.367
R1000 B.n982 B.n39 163.367
R1001 B.n982 B.n43 163.367
R1002 B.n978 B.n43 163.367
R1003 B.n978 B.n45 163.367
R1004 B.n974 B.n45 163.367
R1005 B.n974 B.n51 163.367
R1006 B.n970 B.n51 163.367
R1007 B.n970 B.n53 163.367
R1008 B.n966 B.n53 163.367
R1009 B.n966 B.n58 163.367
R1010 B.n962 B.n58 163.367
R1011 B.n962 B.n60 163.367
R1012 B.n958 B.n60 163.367
R1013 B.n958 B.n65 163.367
R1014 B.n954 B.n65 163.367
R1015 B.n954 B.n67 163.367
R1016 B.n950 B.n67 163.367
R1017 B.n950 B.n72 163.367
R1018 B.n946 B.n72 163.367
R1019 B.n946 B.n74 163.367
R1020 B.n942 B.n74 163.367
R1021 B.n942 B.n79 163.367
R1022 B.n938 B.n79 163.367
R1023 B.n938 B.n81 163.367
R1024 B.n934 B.n81 163.367
R1025 B.n934 B.n86 163.367
R1026 B.n930 B.n86 163.367
R1027 B.n930 B.n88 163.367
R1028 B.n926 B.n88 163.367
R1029 B.n926 B.n93 163.367
R1030 B.n922 B.n93 163.367
R1031 B.n922 B.n95 163.367
R1032 B.n918 B.n95 163.367
R1033 B.n918 B.n100 163.367
R1034 B.n914 B.n100 163.367
R1035 B.n914 B.n102 163.367
R1036 B.n910 B.n102 163.367
R1037 B.n910 B.n107 163.367
R1038 B.n644 B.n434 163.367
R1039 B.n644 B.n476 163.367
R1040 B.n640 B.n639 163.367
R1041 B.n636 B.n635 163.367
R1042 B.n632 B.n631 163.367
R1043 B.n628 B.n627 163.367
R1044 B.n624 B.n623 163.367
R1045 B.n620 B.n619 163.367
R1046 B.n616 B.n615 163.367
R1047 B.n612 B.n611 163.367
R1048 B.n608 B.n607 163.367
R1049 B.n604 B.n603 163.367
R1050 B.n600 B.n599 163.367
R1051 B.n596 B.n595 163.367
R1052 B.n592 B.n591 163.367
R1053 B.n588 B.n587 163.367
R1054 B.n584 B.n583 163.367
R1055 B.n580 B.n579 163.367
R1056 B.n576 B.n575 163.367
R1057 B.n572 B.n571 163.367
R1058 B.n568 B.n567 163.367
R1059 B.n564 B.n563 163.367
R1060 B.n560 B.n559 163.367
R1061 B.n556 B.n555 163.367
R1062 B.n552 B.n551 163.367
R1063 B.n548 B.n547 163.367
R1064 B.n544 B.n543 163.367
R1065 B.n540 B.n539 163.367
R1066 B.n536 B.n535 163.367
R1067 B.n532 B.n531 163.367
R1068 B.n528 B.n527 163.367
R1069 B.n524 B.n523 163.367
R1070 B.n520 B.n519 163.367
R1071 B.n516 B.n515 163.367
R1072 B.n512 B.n511 163.367
R1073 B.n508 B.n507 163.367
R1074 B.n504 B.n503 163.367
R1075 B.n500 B.n499 163.367
R1076 B.n496 B.n495 163.367
R1077 B.n492 B.n491 163.367
R1078 B.n488 B.n487 163.367
R1079 B.n484 B.n475 163.367
R1080 B.n653 B.n430 163.367
R1081 B.n653 B.n428 163.367
R1082 B.n657 B.n428 163.367
R1083 B.n657 B.n422 163.367
R1084 B.n665 B.n422 163.367
R1085 B.n665 B.n420 163.367
R1086 B.n669 B.n420 163.367
R1087 B.n669 B.n414 163.367
R1088 B.n677 B.n414 163.367
R1089 B.n677 B.n412 163.367
R1090 B.n681 B.n412 163.367
R1091 B.n681 B.n406 163.367
R1092 B.n689 B.n406 163.367
R1093 B.n689 B.n404 163.367
R1094 B.n693 B.n404 163.367
R1095 B.n693 B.n398 163.367
R1096 B.n701 B.n398 163.367
R1097 B.n701 B.n396 163.367
R1098 B.n705 B.n396 163.367
R1099 B.n705 B.n390 163.367
R1100 B.n713 B.n390 163.367
R1101 B.n713 B.n388 163.367
R1102 B.n717 B.n388 163.367
R1103 B.n717 B.n382 163.367
R1104 B.n725 B.n382 163.367
R1105 B.n725 B.n380 163.367
R1106 B.n729 B.n380 163.367
R1107 B.n729 B.n374 163.367
R1108 B.n737 B.n374 163.367
R1109 B.n737 B.n372 163.367
R1110 B.n741 B.n372 163.367
R1111 B.n741 B.n366 163.367
R1112 B.n749 B.n366 163.367
R1113 B.n749 B.n364 163.367
R1114 B.n753 B.n364 163.367
R1115 B.n753 B.n359 163.367
R1116 B.n762 B.n359 163.367
R1117 B.n762 B.n357 163.367
R1118 B.n766 B.n357 163.367
R1119 B.n766 B.n351 163.367
R1120 B.n774 B.n351 163.367
R1121 B.n774 B.n349 163.367
R1122 B.n778 B.n349 163.367
R1123 B.n778 B.n344 163.367
R1124 B.n787 B.n344 163.367
R1125 B.n787 B.n342 163.367
R1126 B.n791 B.n342 163.367
R1127 B.n791 B.n336 163.367
R1128 B.n799 B.n336 163.367
R1129 B.n799 B.n334 163.367
R1130 B.n803 B.n334 163.367
R1131 B.n803 B.n328 163.367
R1132 B.n811 B.n328 163.367
R1133 B.n811 B.n326 163.367
R1134 B.n816 B.n326 163.367
R1135 B.n816 B.n320 163.367
R1136 B.n824 B.n320 163.367
R1137 B.n825 B.n824 163.367
R1138 B.n825 B.n5 163.367
R1139 B.n6 B.n5 163.367
R1140 B.n7 B.n6 163.367
R1141 B.n830 B.n7 163.367
R1142 B.n830 B.n12 163.367
R1143 B.n13 B.n12 163.367
R1144 B.n14 B.n13 163.367
R1145 B.n835 B.n14 163.367
R1146 B.n835 B.n19 163.367
R1147 B.n20 B.n19 163.367
R1148 B.n21 B.n20 163.367
R1149 B.n840 B.n21 163.367
R1150 B.n840 B.n26 163.367
R1151 B.n27 B.n26 163.367
R1152 B.n28 B.n27 163.367
R1153 B.n845 B.n28 163.367
R1154 B.n845 B.n33 163.367
R1155 B.n34 B.n33 163.367
R1156 B.n35 B.n34 163.367
R1157 B.n850 B.n35 163.367
R1158 B.n850 B.n40 163.367
R1159 B.n41 B.n40 163.367
R1160 B.n42 B.n41 163.367
R1161 B.n855 B.n42 163.367
R1162 B.n855 B.n47 163.367
R1163 B.n48 B.n47 163.367
R1164 B.n49 B.n48 163.367
R1165 B.n860 B.n49 163.367
R1166 B.n860 B.n54 163.367
R1167 B.n55 B.n54 163.367
R1168 B.n56 B.n55 163.367
R1169 B.n865 B.n56 163.367
R1170 B.n865 B.n61 163.367
R1171 B.n62 B.n61 163.367
R1172 B.n63 B.n62 163.367
R1173 B.n870 B.n63 163.367
R1174 B.n870 B.n68 163.367
R1175 B.n69 B.n68 163.367
R1176 B.n70 B.n69 163.367
R1177 B.n875 B.n70 163.367
R1178 B.n875 B.n75 163.367
R1179 B.n76 B.n75 163.367
R1180 B.n77 B.n76 163.367
R1181 B.n880 B.n77 163.367
R1182 B.n880 B.n82 163.367
R1183 B.n83 B.n82 163.367
R1184 B.n84 B.n83 163.367
R1185 B.n885 B.n84 163.367
R1186 B.n885 B.n89 163.367
R1187 B.n90 B.n89 163.367
R1188 B.n91 B.n90 163.367
R1189 B.n890 B.n91 163.367
R1190 B.n890 B.n96 163.367
R1191 B.n97 B.n96 163.367
R1192 B.n98 B.n97 163.367
R1193 B.n895 B.n98 163.367
R1194 B.n895 B.n103 163.367
R1195 B.n104 B.n103 163.367
R1196 B.n105 B.n104 163.367
R1197 B.n151 B.n105 163.367
R1198 B.n156 B.n109 163.367
R1199 B.n160 B.n159 163.367
R1200 B.n164 B.n163 163.367
R1201 B.n168 B.n167 163.367
R1202 B.n172 B.n171 163.367
R1203 B.n176 B.n175 163.367
R1204 B.n180 B.n179 163.367
R1205 B.n184 B.n183 163.367
R1206 B.n188 B.n187 163.367
R1207 B.n192 B.n191 163.367
R1208 B.n196 B.n195 163.367
R1209 B.n200 B.n199 163.367
R1210 B.n204 B.n203 163.367
R1211 B.n208 B.n207 163.367
R1212 B.n212 B.n211 163.367
R1213 B.n216 B.n215 163.367
R1214 B.n220 B.n219 163.367
R1215 B.n224 B.n223 163.367
R1216 B.n229 B.n228 163.367
R1217 B.n233 B.n232 163.367
R1218 B.n237 B.n236 163.367
R1219 B.n241 B.n240 163.367
R1220 B.n245 B.n244 163.367
R1221 B.n250 B.n249 163.367
R1222 B.n254 B.n253 163.367
R1223 B.n258 B.n257 163.367
R1224 B.n262 B.n261 163.367
R1225 B.n266 B.n265 163.367
R1226 B.n270 B.n269 163.367
R1227 B.n274 B.n273 163.367
R1228 B.n278 B.n277 163.367
R1229 B.n282 B.n281 163.367
R1230 B.n286 B.n285 163.367
R1231 B.n290 B.n289 163.367
R1232 B.n294 B.n293 163.367
R1233 B.n298 B.n297 163.367
R1234 B.n302 B.n301 163.367
R1235 B.n306 B.n305 163.367
R1236 B.n310 B.n309 163.367
R1237 B.n314 B.n313 163.367
R1238 B.n316 B.n150 163.367
R1239 B.n480 B.t13 129.311
R1240 B.n152 B.t16 129.311
R1241 B.n477 B.t23 129.298
R1242 B.n154 B.t19 129.298
R1243 B.n645 B.n431 83.0852
R1244 B.n904 B.n106 83.0852
R1245 B.n481 B.t12 73.457
R1246 B.n153 B.t17 73.457
R1247 B.n478 B.t22 73.4443
R1248 B.n155 B.t20 73.4443
R1249 B.n647 B.n646 71.676
R1250 B.n476 B.n435 71.676
R1251 B.n639 B.n436 71.676
R1252 B.n635 B.n437 71.676
R1253 B.n631 B.n438 71.676
R1254 B.n627 B.n439 71.676
R1255 B.n623 B.n440 71.676
R1256 B.n619 B.n441 71.676
R1257 B.n615 B.n442 71.676
R1258 B.n611 B.n443 71.676
R1259 B.n607 B.n444 71.676
R1260 B.n603 B.n445 71.676
R1261 B.n599 B.n446 71.676
R1262 B.n595 B.n447 71.676
R1263 B.n591 B.n448 71.676
R1264 B.n587 B.n449 71.676
R1265 B.n583 B.n450 71.676
R1266 B.n579 B.n451 71.676
R1267 B.n575 B.n452 71.676
R1268 B.n571 B.n453 71.676
R1269 B.n567 B.n454 71.676
R1270 B.n563 B.n455 71.676
R1271 B.n559 B.n456 71.676
R1272 B.n555 B.n457 71.676
R1273 B.n551 B.n458 71.676
R1274 B.n547 B.n459 71.676
R1275 B.n543 B.n460 71.676
R1276 B.n539 B.n461 71.676
R1277 B.n535 B.n462 71.676
R1278 B.n531 B.n463 71.676
R1279 B.n527 B.n464 71.676
R1280 B.n523 B.n465 71.676
R1281 B.n519 B.n466 71.676
R1282 B.n515 B.n467 71.676
R1283 B.n511 B.n468 71.676
R1284 B.n507 B.n469 71.676
R1285 B.n503 B.n470 71.676
R1286 B.n499 B.n471 71.676
R1287 B.n495 B.n472 71.676
R1288 B.n491 B.n473 71.676
R1289 B.n487 B.n474 71.676
R1290 B.n906 B.n905 71.676
R1291 B.n156 B.n110 71.676
R1292 B.n160 B.n111 71.676
R1293 B.n164 B.n112 71.676
R1294 B.n168 B.n113 71.676
R1295 B.n172 B.n114 71.676
R1296 B.n176 B.n115 71.676
R1297 B.n180 B.n116 71.676
R1298 B.n184 B.n117 71.676
R1299 B.n188 B.n118 71.676
R1300 B.n192 B.n119 71.676
R1301 B.n196 B.n120 71.676
R1302 B.n200 B.n121 71.676
R1303 B.n204 B.n122 71.676
R1304 B.n208 B.n123 71.676
R1305 B.n212 B.n124 71.676
R1306 B.n216 B.n125 71.676
R1307 B.n220 B.n126 71.676
R1308 B.n224 B.n127 71.676
R1309 B.n229 B.n128 71.676
R1310 B.n233 B.n129 71.676
R1311 B.n237 B.n130 71.676
R1312 B.n241 B.n131 71.676
R1313 B.n245 B.n132 71.676
R1314 B.n250 B.n133 71.676
R1315 B.n254 B.n134 71.676
R1316 B.n258 B.n135 71.676
R1317 B.n262 B.n136 71.676
R1318 B.n266 B.n137 71.676
R1319 B.n270 B.n138 71.676
R1320 B.n274 B.n139 71.676
R1321 B.n278 B.n140 71.676
R1322 B.n282 B.n141 71.676
R1323 B.n286 B.n142 71.676
R1324 B.n290 B.n143 71.676
R1325 B.n294 B.n144 71.676
R1326 B.n298 B.n145 71.676
R1327 B.n302 B.n146 71.676
R1328 B.n306 B.n147 71.676
R1329 B.n310 B.n148 71.676
R1330 B.n314 B.n149 71.676
R1331 B.n903 B.n150 71.676
R1332 B.n903 B.n902 71.676
R1333 B.n316 B.n149 71.676
R1334 B.n313 B.n148 71.676
R1335 B.n309 B.n147 71.676
R1336 B.n305 B.n146 71.676
R1337 B.n301 B.n145 71.676
R1338 B.n297 B.n144 71.676
R1339 B.n293 B.n143 71.676
R1340 B.n289 B.n142 71.676
R1341 B.n285 B.n141 71.676
R1342 B.n281 B.n140 71.676
R1343 B.n277 B.n139 71.676
R1344 B.n273 B.n138 71.676
R1345 B.n269 B.n137 71.676
R1346 B.n265 B.n136 71.676
R1347 B.n261 B.n135 71.676
R1348 B.n257 B.n134 71.676
R1349 B.n253 B.n133 71.676
R1350 B.n249 B.n132 71.676
R1351 B.n244 B.n131 71.676
R1352 B.n240 B.n130 71.676
R1353 B.n236 B.n129 71.676
R1354 B.n232 B.n128 71.676
R1355 B.n228 B.n127 71.676
R1356 B.n223 B.n126 71.676
R1357 B.n219 B.n125 71.676
R1358 B.n215 B.n124 71.676
R1359 B.n211 B.n123 71.676
R1360 B.n207 B.n122 71.676
R1361 B.n203 B.n121 71.676
R1362 B.n199 B.n120 71.676
R1363 B.n195 B.n119 71.676
R1364 B.n191 B.n118 71.676
R1365 B.n187 B.n117 71.676
R1366 B.n183 B.n116 71.676
R1367 B.n179 B.n115 71.676
R1368 B.n175 B.n114 71.676
R1369 B.n171 B.n113 71.676
R1370 B.n167 B.n112 71.676
R1371 B.n163 B.n111 71.676
R1372 B.n159 B.n110 71.676
R1373 B.n905 B.n109 71.676
R1374 B.n646 B.n434 71.676
R1375 B.n640 B.n435 71.676
R1376 B.n636 B.n436 71.676
R1377 B.n632 B.n437 71.676
R1378 B.n628 B.n438 71.676
R1379 B.n624 B.n439 71.676
R1380 B.n620 B.n440 71.676
R1381 B.n616 B.n441 71.676
R1382 B.n612 B.n442 71.676
R1383 B.n608 B.n443 71.676
R1384 B.n604 B.n444 71.676
R1385 B.n600 B.n445 71.676
R1386 B.n596 B.n446 71.676
R1387 B.n592 B.n447 71.676
R1388 B.n588 B.n448 71.676
R1389 B.n584 B.n449 71.676
R1390 B.n580 B.n450 71.676
R1391 B.n576 B.n451 71.676
R1392 B.n572 B.n452 71.676
R1393 B.n568 B.n453 71.676
R1394 B.n564 B.n454 71.676
R1395 B.n560 B.n455 71.676
R1396 B.n556 B.n456 71.676
R1397 B.n552 B.n457 71.676
R1398 B.n548 B.n458 71.676
R1399 B.n544 B.n459 71.676
R1400 B.n540 B.n460 71.676
R1401 B.n536 B.n461 71.676
R1402 B.n532 B.n462 71.676
R1403 B.n528 B.n463 71.676
R1404 B.n524 B.n464 71.676
R1405 B.n520 B.n465 71.676
R1406 B.n516 B.n466 71.676
R1407 B.n512 B.n467 71.676
R1408 B.n508 B.n468 71.676
R1409 B.n504 B.n469 71.676
R1410 B.n500 B.n470 71.676
R1411 B.n496 B.n471 71.676
R1412 B.n492 B.n472 71.676
R1413 B.n488 B.n473 71.676
R1414 B.n484 B.n474 71.676
R1415 B.n482 B.n481 59.5399
R1416 B.n479 B.n478 59.5399
R1417 B.n226 B.n155 59.5399
R1418 B.n247 B.n153 59.5399
R1419 B.n481 B.n480 55.855
R1420 B.n478 B.n477 55.855
R1421 B.n155 B.n154 55.855
R1422 B.n153 B.n152 55.855
R1423 B.n652 B.n431 47.4775
R1424 B.n652 B.n427 47.4775
R1425 B.n658 B.n427 47.4775
R1426 B.n658 B.n423 47.4775
R1427 B.n664 B.n423 47.4775
R1428 B.n664 B.n419 47.4775
R1429 B.n670 B.n419 47.4775
R1430 B.n676 B.n415 47.4775
R1431 B.n676 B.n411 47.4775
R1432 B.n682 B.n411 47.4775
R1433 B.n682 B.n407 47.4775
R1434 B.n688 B.n407 47.4775
R1435 B.n688 B.n403 47.4775
R1436 B.n694 B.n403 47.4775
R1437 B.n694 B.n399 47.4775
R1438 B.n700 B.n399 47.4775
R1439 B.n700 B.n395 47.4775
R1440 B.n706 B.n395 47.4775
R1441 B.n712 B.n391 47.4775
R1442 B.n712 B.n387 47.4775
R1443 B.n718 B.n387 47.4775
R1444 B.n718 B.n383 47.4775
R1445 B.n724 B.n383 47.4775
R1446 B.n724 B.n379 47.4775
R1447 B.n730 B.n379 47.4775
R1448 B.n736 B.n375 47.4775
R1449 B.n736 B.n371 47.4775
R1450 B.n742 B.n371 47.4775
R1451 B.n742 B.n367 47.4775
R1452 B.n748 B.n367 47.4775
R1453 B.n748 B.n363 47.4775
R1454 B.n755 B.n363 47.4775
R1455 B.n755 B.n754 47.4775
R1456 B.n761 B.n356 47.4775
R1457 B.n767 B.n356 47.4775
R1458 B.n767 B.n352 47.4775
R1459 B.n773 B.n352 47.4775
R1460 B.n773 B.n348 47.4775
R1461 B.n780 B.n348 47.4775
R1462 B.n780 B.n779 47.4775
R1463 B.n786 B.n341 47.4775
R1464 B.n792 B.n341 47.4775
R1465 B.n792 B.n337 47.4775
R1466 B.n798 B.n337 47.4775
R1467 B.n798 B.n333 47.4775
R1468 B.n804 B.n333 47.4775
R1469 B.n804 B.n329 47.4775
R1470 B.n810 B.n329 47.4775
R1471 B.n817 B.n325 47.4775
R1472 B.n817 B.n321 47.4775
R1473 B.n823 B.n321 47.4775
R1474 B.n823 B.n4 47.4775
R1475 B.n1025 B.n4 47.4775
R1476 B.n1025 B.n1024 47.4775
R1477 B.n1024 B.n1023 47.4775
R1478 B.n1023 B.n8 47.4775
R1479 B.n1017 B.n8 47.4775
R1480 B.n1017 B.n1016 47.4775
R1481 B.n1015 B.n15 47.4775
R1482 B.n1009 B.n15 47.4775
R1483 B.n1009 B.n1008 47.4775
R1484 B.n1008 B.n1007 47.4775
R1485 B.n1007 B.n22 47.4775
R1486 B.n1001 B.n22 47.4775
R1487 B.n1001 B.n1000 47.4775
R1488 B.n1000 B.n999 47.4775
R1489 B.n993 B.n32 47.4775
R1490 B.n993 B.n992 47.4775
R1491 B.n992 B.n991 47.4775
R1492 B.n991 B.n36 47.4775
R1493 B.n985 B.n36 47.4775
R1494 B.n985 B.n984 47.4775
R1495 B.n984 B.n983 47.4775
R1496 B.n977 B.n46 47.4775
R1497 B.n977 B.n976 47.4775
R1498 B.n976 B.n975 47.4775
R1499 B.n975 B.n50 47.4775
R1500 B.n969 B.n50 47.4775
R1501 B.n969 B.n968 47.4775
R1502 B.n968 B.n967 47.4775
R1503 B.n967 B.n57 47.4775
R1504 B.n961 B.n960 47.4775
R1505 B.n960 B.n959 47.4775
R1506 B.n959 B.n64 47.4775
R1507 B.n953 B.n64 47.4775
R1508 B.n953 B.n952 47.4775
R1509 B.n952 B.n951 47.4775
R1510 B.n951 B.n71 47.4775
R1511 B.n945 B.n944 47.4775
R1512 B.n944 B.n943 47.4775
R1513 B.n943 B.n78 47.4775
R1514 B.n937 B.n78 47.4775
R1515 B.n937 B.n936 47.4775
R1516 B.n936 B.n935 47.4775
R1517 B.n935 B.n85 47.4775
R1518 B.n929 B.n85 47.4775
R1519 B.n929 B.n928 47.4775
R1520 B.n928 B.n927 47.4775
R1521 B.n927 B.n92 47.4775
R1522 B.n921 B.n920 47.4775
R1523 B.n920 B.n919 47.4775
R1524 B.n919 B.n99 47.4775
R1525 B.n913 B.n99 47.4775
R1526 B.n913 B.n912 47.4775
R1527 B.n912 B.n911 47.4775
R1528 B.n911 B.n106 47.4775
R1529 B.t2 B.n325 39.7974
R1530 B.n1016 B.t1 39.7974
R1531 B.n761 B.t7 37.0046
R1532 B.n983 B.t5 37.0046
R1533 B.n730 B.t8 35.6082
R1534 B.n961 B.t9 35.6082
R1535 B.t0 B.n391 34.2119
R1536 B.t4 B.n71 34.2119
R1537 B.n779 B.t6 32.8155
R1538 B.n32 B.t3 32.8155
R1539 B.n908 B.n907 31.0639
R1540 B.n901 B.n900 31.0639
R1541 B.n483 B.n429 31.0639
R1542 B.n649 B.n648 31.0639
R1543 B.n670 B.t11 28.6263
R1544 B.n921 B.t15 28.6263
R1545 B.t11 B.n415 18.8517
R1546 B.t15 B.n92 18.8517
R1547 B B.n1027 18.0485
R1548 B.n786 B.t6 14.6625
R1549 B.n999 B.t3 14.6625
R1550 B.n706 B.t0 13.2661
R1551 B.n945 B.t4 13.2661
R1552 B.t8 B.n375 11.8697
R1553 B.t9 B.n57 11.8697
R1554 B.n907 B.n108 10.6151
R1555 B.n157 B.n108 10.6151
R1556 B.n158 B.n157 10.6151
R1557 B.n161 B.n158 10.6151
R1558 B.n162 B.n161 10.6151
R1559 B.n165 B.n162 10.6151
R1560 B.n166 B.n165 10.6151
R1561 B.n169 B.n166 10.6151
R1562 B.n170 B.n169 10.6151
R1563 B.n173 B.n170 10.6151
R1564 B.n174 B.n173 10.6151
R1565 B.n177 B.n174 10.6151
R1566 B.n178 B.n177 10.6151
R1567 B.n181 B.n178 10.6151
R1568 B.n182 B.n181 10.6151
R1569 B.n185 B.n182 10.6151
R1570 B.n186 B.n185 10.6151
R1571 B.n189 B.n186 10.6151
R1572 B.n190 B.n189 10.6151
R1573 B.n193 B.n190 10.6151
R1574 B.n194 B.n193 10.6151
R1575 B.n197 B.n194 10.6151
R1576 B.n198 B.n197 10.6151
R1577 B.n201 B.n198 10.6151
R1578 B.n202 B.n201 10.6151
R1579 B.n205 B.n202 10.6151
R1580 B.n206 B.n205 10.6151
R1581 B.n209 B.n206 10.6151
R1582 B.n210 B.n209 10.6151
R1583 B.n213 B.n210 10.6151
R1584 B.n214 B.n213 10.6151
R1585 B.n217 B.n214 10.6151
R1586 B.n218 B.n217 10.6151
R1587 B.n221 B.n218 10.6151
R1588 B.n222 B.n221 10.6151
R1589 B.n225 B.n222 10.6151
R1590 B.n230 B.n227 10.6151
R1591 B.n231 B.n230 10.6151
R1592 B.n234 B.n231 10.6151
R1593 B.n235 B.n234 10.6151
R1594 B.n238 B.n235 10.6151
R1595 B.n239 B.n238 10.6151
R1596 B.n242 B.n239 10.6151
R1597 B.n243 B.n242 10.6151
R1598 B.n246 B.n243 10.6151
R1599 B.n251 B.n248 10.6151
R1600 B.n252 B.n251 10.6151
R1601 B.n255 B.n252 10.6151
R1602 B.n256 B.n255 10.6151
R1603 B.n259 B.n256 10.6151
R1604 B.n260 B.n259 10.6151
R1605 B.n263 B.n260 10.6151
R1606 B.n264 B.n263 10.6151
R1607 B.n267 B.n264 10.6151
R1608 B.n268 B.n267 10.6151
R1609 B.n271 B.n268 10.6151
R1610 B.n272 B.n271 10.6151
R1611 B.n275 B.n272 10.6151
R1612 B.n276 B.n275 10.6151
R1613 B.n279 B.n276 10.6151
R1614 B.n280 B.n279 10.6151
R1615 B.n283 B.n280 10.6151
R1616 B.n284 B.n283 10.6151
R1617 B.n287 B.n284 10.6151
R1618 B.n288 B.n287 10.6151
R1619 B.n291 B.n288 10.6151
R1620 B.n292 B.n291 10.6151
R1621 B.n295 B.n292 10.6151
R1622 B.n296 B.n295 10.6151
R1623 B.n299 B.n296 10.6151
R1624 B.n300 B.n299 10.6151
R1625 B.n303 B.n300 10.6151
R1626 B.n304 B.n303 10.6151
R1627 B.n307 B.n304 10.6151
R1628 B.n308 B.n307 10.6151
R1629 B.n311 B.n308 10.6151
R1630 B.n312 B.n311 10.6151
R1631 B.n315 B.n312 10.6151
R1632 B.n317 B.n315 10.6151
R1633 B.n318 B.n317 10.6151
R1634 B.n901 B.n318 10.6151
R1635 B.n654 B.n429 10.6151
R1636 B.n655 B.n654 10.6151
R1637 B.n656 B.n655 10.6151
R1638 B.n656 B.n421 10.6151
R1639 B.n666 B.n421 10.6151
R1640 B.n667 B.n666 10.6151
R1641 B.n668 B.n667 10.6151
R1642 B.n668 B.n413 10.6151
R1643 B.n678 B.n413 10.6151
R1644 B.n679 B.n678 10.6151
R1645 B.n680 B.n679 10.6151
R1646 B.n680 B.n405 10.6151
R1647 B.n690 B.n405 10.6151
R1648 B.n691 B.n690 10.6151
R1649 B.n692 B.n691 10.6151
R1650 B.n692 B.n397 10.6151
R1651 B.n702 B.n397 10.6151
R1652 B.n703 B.n702 10.6151
R1653 B.n704 B.n703 10.6151
R1654 B.n704 B.n389 10.6151
R1655 B.n714 B.n389 10.6151
R1656 B.n715 B.n714 10.6151
R1657 B.n716 B.n715 10.6151
R1658 B.n716 B.n381 10.6151
R1659 B.n726 B.n381 10.6151
R1660 B.n727 B.n726 10.6151
R1661 B.n728 B.n727 10.6151
R1662 B.n728 B.n373 10.6151
R1663 B.n738 B.n373 10.6151
R1664 B.n739 B.n738 10.6151
R1665 B.n740 B.n739 10.6151
R1666 B.n740 B.n365 10.6151
R1667 B.n750 B.n365 10.6151
R1668 B.n751 B.n750 10.6151
R1669 B.n752 B.n751 10.6151
R1670 B.n752 B.n358 10.6151
R1671 B.n763 B.n358 10.6151
R1672 B.n764 B.n763 10.6151
R1673 B.n765 B.n764 10.6151
R1674 B.n765 B.n350 10.6151
R1675 B.n775 B.n350 10.6151
R1676 B.n776 B.n775 10.6151
R1677 B.n777 B.n776 10.6151
R1678 B.n777 B.n343 10.6151
R1679 B.n788 B.n343 10.6151
R1680 B.n789 B.n788 10.6151
R1681 B.n790 B.n789 10.6151
R1682 B.n790 B.n335 10.6151
R1683 B.n800 B.n335 10.6151
R1684 B.n801 B.n800 10.6151
R1685 B.n802 B.n801 10.6151
R1686 B.n802 B.n327 10.6151
R1687 B.n812 B.n327 10.6151
R1688 B.n813 B.n812 10.6151
R1689 B.n815 B.n813 10.6151
R1690 B.n815 B.n814 10.6151
R1691 B.n814 B.n319 10.6151
R1692 B.n826 B.n319 10.6151
R1693 B.n827 B.n826 10.6151
R1694 B.n828 B.n827 10.6151
R1695 B.n829 B.n828 10.6151
R1696 B.n831 B.n829 10.6151
R1697 B.n832 B.n831 10.6151
R1698 B.n833 B.n832 10.6151
R1699 B.n834 B.n833 10.6151
R1700 B.n836 B.n834 10.6151
R1701 B.n837 B.n836 10.6151
R1702 B.n838 B.n837 10.6151
R1703 B.n839 B.n838 10.6151
R1704 B.n841 B.n839 10.6151
R1705 B.n842 B.n841 10.6151
R1706 B.n843 B.n842 10.6151
R1707 B.n844 B.n843 10.6151
R1708 B.n846 B.n844 10.6151
R1709 B.n847 B.n846 10.6151
R1710 B.n848 B.n847 10.6151
R1711 B.n849 B.n848 10.6151
R1712 B.n851 B.n849 10.6151
R1713 B.n852 B.n851 10.6151
R1714 B.n853 B.n852 10.6151
R1715 B.n854 B.n853 10.6151
R1716 B.n856 B.n854 10.6151
R1717 B.n857 B.n856 10.6151
R1718 B.n858 B.n857 10.6151
R1719 B.n859 B.n858 10.6151
R1720 B.n861 B.n859 10.6151
R1721 B.n862 B.n861 10.6151
R1722 B.n863 B.n862 10.6151
R1723 B.n864 B.n863 10.6151
R1724 B.n866 B.n864 10.6151
R1725 B.n867 B.n866 10.6151
R1726 B.n868 B.n867 10.6151
R1727 B.n869 B.n868 10.6151
R1728 B.n871 B.n869 10.6151
R1729 B.n872 B.n871 10.6151
R1730 B.n873 B.n872 10.6151
R1731 B.n874 B.n873 10.6151
R1732 B.n876 B.n874 10.6151
R1733 B.n877 B.n876 10.6151
R1734 B.n878 B.n877 10.6151
R1735 B.n879 B.n878 10.6151
R1736 B.n881 B.n879 10.6151
R1737 B.n882 B.n881 10.6151
R1738 B.n883 B.n882 10.6151
R1739 B.n884 B.n883 10.6151
R1740 B.n886 B.n884 10.6151
R1741 B.n887 B.n886 10.6151
R1742 B.n888 B.n887 10.6151
R1743 B.n889 B.n888 10.6151
R1744 B.n891 B.n889 10.6151
R1745 B.n892 B.n891 10.6151
R1746 B.n893 B.n892 10.6151
R1747 B.n894 B.n893 10.6151
R1748 B.n896 B.n894 10.6151
R1749 B.n897 B.n896 10.6151
R1750 B.n898 B.n897 10.6151
R1751 B.n899 B.n898 10.6151
R1752 B.n900 B.n899 10.6151
R1753 B.n648 B.n433 10.6151
R1754 B.n643 B.n433 10.6151
R1755 B.n643 B.n642 10.6151
R1756 B.n642 B.n641 10.6151
R1757 B.n641 B.n638 10.6151
R1758 B.n638 B.n637 10.6151
R1759 B.n637 B.n634 10.6151
R1760 B.n634 B.n633 10.6151
R1761 B.n633 B.n630 10.6151
R1762 B.n630 B.n629 10.6151
R1763 B.n629 B.n626 10.6151
R1764 B.n626 B.n625 10.6151
R1765 B.n625 B.n622 10.6151
R1766 B.n622 B.n621 10.6151
R1767 B.n621 B.n618 10.6151
R1768 B.n618 B.n617 10.6151
R1769 B.n617 B.n614 10.6151
R1770 B.n614 B.n613 10.6151
R1771 B.n613 B.n610 10.6151
R1772 B.n610 B.n609 10.6151
R1773 B.n609 B.n606 10.6151
R1774 B.n606 B.n605 10.6151
R1775 B.n605 B.n602 10.6151
R1776 B.n602 B.n601 10.6151
R1777 B.n601 B.n598 10.6151
R1778 B.n598 B.n597 10.6151
R1779 B.n597 B.n594 10.6151
R1780 B.n594 B.n593 10.6151
R1781 B.n593 B.n590 10.6151
R1782 B.n590 B.n589 10.6151
R1783 B.n589 B.n586 10.6151
R1784 B.n586 B.n585 10.6151
R1785 B.n585 B.n582 10.6151
R1786 B.n582 B.n581 10.6151
R1787 B.n581 B.n578 10.6151
R1788 B.n578 B.n577 10.6151
R1789 B.n574 B.n573 10.6151
R1790 B.n573 B.n570 10.6151
R1791 B.n570 B.n569 10.6151
R1792 B.n569 B.n566 10.6151
R1793 B.n566 B.n565 10.6151
R1794 B.n565 B.n562 10.6151
R1795 B.n562 B.n561 10.6151
R1796 B.n561 B.n558 10.6151
R1797 B.n558 B.n557 10.6151
R1798 B.n554 B.n553 10.6151
R1799 B.n553 B.n550 10.6151
R1800 B.n550 B.n549 10.6151
R1801 B.n549 B.n546 10.6151
R1802 B.n546 B.n545 10.6151
R1803 B.n545 B.n542 10.6151
R1804 B.n542 B.n541 10.6151
R1805 B.n541 B.n538 10.6151
R1806 B.n538 B.n537 10.6151
R1807 B.n537 B.n534 10.6151
R1808 B.n534 B.n533 10.6151
R1809 B.n533 B.n530 10.6151
R1810 B.n530 B.n529 10.6151
R1811 B.n529 B.n526 10.6151
R1812 B.n526 B.n525 10.6151
R1813 B.n525 B.n522 10.6151
R1814 B.n522 B.n521 10.6151
R1815 B.n521 B.n518 10.6151
R1816 B.n518 B.n517 10.6151
R1817 B.n517 B.n514 10.6151
R1818 B.n514 B.n513 10.6151
R1819 B.n513 B.n510 10.6151
R1820 B.n510 B.n509 10.6151
R1821 B.n509 B.n506 10.6151
R1822 B.n506 B.n505 10.6151
R1823 B.n505 B.n502 10.6151
R1824 B.n502 B.n501 10.6151
R1825 B.n501 B.n498 10.6151
R1826 B.n498 B.n497 10.6151
R1827 B.n497 B.n494 10.6151
R1828 B.n494 B.n493 10.6151
R1829 B.n493 B.n490 10.6151
R1830 B.n490 B.n489 10.6151
R1831 B.n489 B.n486 10.6151
R1832 B.n486 B.n485 10.6151
R1833 B.n485 B.n483 10.6151
R1834 B.n650 B.n649 10.6151
R1835 B.n650 B.n425 10.6151
R1836 B.n660 B.n425 10.6151
R1837 B.n661 B.n660 10.6151
R1838 B.n662 B.n661 10.6151
R1839 B.n662 B.n417 10.6151
R1840 B.n672 B.n417 10.6151
R1841 B.n673 B.n672 10.6151
R1842 B.n674 B.n673 10.6151
R1843 B.n674 B.n409 10.6151
R1844 B.n684 B.n409 10.6151
R1845 B.n685 B.n684 10.6151
R1846 B.n686 B.n685 10.6151
R1847 B.n686 B.n401 10.6151
R1848 B.n696 B.n401 10.6151
R1849 B.n697 B.n696 10.6151
R1850 B.n698 B.n697 10.6151
R1851 B.n698 B.n393 10.6151
R1852 B.n708 B.n393 10.6151
R1853 B.n709 B.n708 10.6151
R1854 B.n710 B.n709 10.6151
R1855 B.n710 B.n385 10.6151
R1856 B.n720 B.n385 10.6151
R1857 B.n721 B.n720 10.6151
R1858 B.n722 B.n721 10.6151
R1859 B.n722 B.n377 10.6151
R1860 B.n732 B.n377 10.6151
R1861 B.n733 B.n732 10.6151
R1862 B.n734 B.n733 10.6151
R1863 B.n734 B.n369 10.6151
R1864 B.n744 B.n369 10.6151
R1865 B.n745 B.n744 10.6151
R1866 B.n746 B.n745 10.6151
R1867 B.n746 B.n361 10.6151
R1868 B.n757 B.n361 10.6151
R1869 B.n758 B.n757 10.6151
R1870 B.n759 B.n758 10.6151
R1871 B.n759 B.n354 10.6151
R1872 B.n769 B.n354 10.6151
R1873 B.n770 B.n769 10.6151
R1874 B.n771 B.n770 10.6151
R1875 B.n771 B.n346 10.6151
R1876 B.n782 B.n346 10.6151
R1877 B.n783 B.n782 10.6151
R1878 B.n784 B.n783 10.6151
R1879 B.n784 B.n339 10.6151
R1880 B.n794 B.n339 10.6151
R1881 B.n795 B.n794 10.6151
R1882 B.n796 B.n795 10.6151
R1883 B.n796 B.n331 10.6151
R1884 B.n806 B.n331 10.6151
R1885 B.n807 B.n806 10.6151
R1886 B.n808 B.n807 10.6151
R1887 B.n808 B.n323 10.6151
R1888 B.n819 B.n323 10.6151
R1889 B.n820 B.n819 10.6151
R1890 B.n821 B.n820 10.6151
R1891 B.n821 B.n0 10.6151
R1892 B.n1021 B.n1 10.6151
R1893 B.n1021 B.n1020 10.6151
R1894 B.n1020 B.n1019 10.6151
R1895 B.n1019 B.n10 10.6151
R1896 B.n1013 B.n10 10.6151
R1897 B.n1013 B.n1012 10.6151
R1898 B.n1012 B.n1011 10.6151
R1899 B.n1011 B.n17 10.6151
R1900 B.n1005 B.n17 10.6151
R1901 B.n1005 B.n1004 10.6151
R1902 B.n1004 B.n1003 10.6151
R1903 B.n1003 B.n24 10.6151
R1904 B.n997 B.n24 10.6151
R1905 B.n997 B.n996 10.6151
R1906 B.n996 B.n995 10.6151
R1907 B.n995 B.n30 10.6151
R1908 B.n989 B.n30 10.6151
R1909 B.n989 B.n988 10.6151
R1910 B.n988 B.n987 10.6151
R1911 B.n987 B.n38 10.6151
R1912 B.n981 B.n38 10.6151
R1913 B.n981 B.n980 10.6151
R1914 B.n980 B.n979 10.6151
R1915 B.n979 B.n44 10.6151
R1916 B.n973 B.n44 10.6151
R1917 B.n973 B.n972 10.6151
R1918 B.n972 B.n971 10.6151
R1919 B.n971 B.n52 10.6151
R1920 B.n965 B.n52 10.6151
R1921 B.n965 B.n964 10.6151
R1922 B.n964 B.n963 10.6151
R1923 B.n963 B.n59 10.6151
R1924 B.n957 B.n59 10.6151
R1925 B.n957 B.n956 10.6151
R1926 B.n956 B.n955 10.6151
R1927 B.n955 B.n66 10.6151
R1928 B.n949 B.n66 10.6151
R1929 B.n949 B.n948 10.6151
R1930 B.n948 B.n947 10.6151
R1931 B.n947 B.n73 10.6151
R1932 B.n941 B.n73 10.6151
R1933 B.n941 B.n940 10.6151
R1934 B.n940 B.n939 10.6151
R1935 B.n939 B.n80 10.6151
R1936 B.n933 B.n80 10.6151
R1937 B.n933 B.n932 10.6151
R1938 B.n932 B.n931 10.6151
R1939 B.n931 B.n87 10.6151
R1940 B.n925 B.n87 10.6151
R1941 B.n925 B.n924 10.6151
R1942 B.n924 B.n923 10.6151
R1943 B.n923 B.n94 10.6151
R1944 B.n917 B.n94 10.6151
R1945 B.n917 B.n916 10.6151
R1946 B.n916 B.n915 10.6151
R1947 B.n915 B.n101 10.6151
R1948 B.n909 B.n101 10.6151
R1949 B.n909 B.n908 10.6151
R1950 B.n754 B.t7 10.4734
R1951 B.n46 B.t5 10.4734
R1952 B.n226 B.n225 9.36635
R1953 B.n248 B.n247 9.36635
R1954 B.n577 B.n479 9.36635
R1955 B.n554 B.n482 9.36635
R1956 B.n810 B.t2 7.6806
R1957 B.t1 B.n1015 7.6806
R1958 B.n1027 B.n0 2.81026
R1959 B.n1027 B.n1 2.81026
R1960 B.n227 B.n226 1.24928
R1961 B.n247 B.n246 1.24928
R1962 B.n574 B.n479 1.24928
R1963 B.n557 B.n482 1.24928
R1964 VP.n25 VP.n24 161.3
R1965 VP.n26 VP.n21 161.3
R1966 VP.n28 VP.n27 161.3
R1967 VP.n29 VP.n20 161.3
R1968 VP.n31 VP.n30 161.3
R1969 VP.n32 VP.n19 161.3
R1970 VP.n34 VP.n33 161.3
R1971 VP.n35 VP.n18 161.3
R1972 VP.n37 VP.n36 161.3
R1973 VP.n38 VP.n17 161.3
R1974 VP.n40 VP.n39 161.3
R1975 VP.n42 VP.n41 161.3
R1976 VP.n43 VP.n15 161.3
R1977 VP.n45 VP.n44 161.3
R1978 VP.n46 VP.n14 161.3
R1979 VP.n48 VP.n47 161.3
R1980 VP.n49 VP.n13 161.3
R1981 VP.n88 VP.n0 161.3
R1982 VP.n87 VP.n86 161.3
R1983 VP.n85 VP.n1 161.3
R1984 VP.n84 VP.n83 161.3
R1985 VP.n82 VP.n2 161.3
R1986 VP.n81 VP.n80 161.3
R1987 VP.n79 VP.n78 161.3
R1988 VP.n77 VP.n4 161.3
R1989 VP.n76 VP.n75 161.3
R1990 VP.n74 VP.n5 161.3
R1991 VP.n73 VP.n72 161.3
R1992 VP.n71 VP.n6 161.3
R1993 VP.n70 VP.n69 161.3
R1994 VP.n68 VP.n7 161.3
R1995 VP.n67 VP.n66 161.3
R1996 VP.n65 VP.n8 161.3
R1997 VP.n64 VP.n63 161.3
R1998 VP.n62 VP.n61 161.3
R1999 VP.n60 VP.n10 161.3
R2000 VP.n59 VP.n58 161.3
R2001 VP.n57 VP.n11 161.3
R2002 VP.n56 VP.n55 161.3
R2003 VP.n54 VP.n12 161.3
R2004 VP.n23 VP.t7 133.29
R2005 VP.n71 VP.t3 99.0468
R2006 VP.n53 VP.t9 99.0468
R2007 VP.n9 VP.t4 99.0468
R2008 VP.n3 VP.t8 99.0468
R2009 VP.n89 VP.t2 99.0468
R2010 VP.n32 VP.t5 99.0468
R2011 VP.n50 VP.t0 99.0468
R2012 VP.n16 VP.t1 99.0468
R2013 VP.n22 VP.t6 99.0468
R2014 VP.n53 VP.n52 97.9476
R2015 VP.n90 VP.n89 97.9476
R2016 VP.n51 VP.n50 97.9476
R2017 VP.n59 VP.n11 56.4773
R2018 VP.n83 VP.n1 56.4773
R2019 VP.n44 VP.n14 56.4773
R2020 VP.n23 VP.n22 53.8957
R2021 VP.n52 VP.n51 51.7419
R2022 VP.n66 VP.n7 46.253
R2023 VP.n76 VP.n5 46.253
R2024 VP.n37 VP.n18 46.253
R2025 VP.n27 VP.n20 46.253
R2026 VP.n66 VP.n65 34.5682
R2027 VP.n77 VP.n76 34.5682
R2028 VP.n38 VP.n37 34.5682
R2029 VP.n27 VP.n26 34.5682
R2030 VP.n55 VP.n54 24.3439
R2031 VP.n55 VP.n11 24.3439
R2032 VP.n60 VP.n59 24.3439
R2033 VP.n61 VP.n60 24.3439
R2034 VP.n65 VP.n64 24.3439
R2035 VP.n70 VP.n7 24.3439
R2036 VP.n71 VP.n70 24.3439
R2037 VP.n72 VP.n71 24.3439
R2038 VP.n72 VP.n5 24.3439
R2039 VP.n78 VP.n77 24.3439
R2040 VP.n82 VP.n81 24.3439
R2041 VP.n83 VP.n82 24.3439
R2042 VP.n87 VP.n1 24.3439
R2043 VP.n88 VP.n87 24.3439
R2044 VP.n48 VP.n14 24.3439
R2045 VP.n49 VP.n48 24.3439
R2046 VP.n39 VP.n38 24.3439
R2047 VP.n43 VP.n42 24.3439
R2048 VP.n44 VP.n43 24.3439
R2049 VP.n31 VP.n20 24.3439
R2050 VP.n32 VP.n31 24.3439
R2051 VP.n33 VP.n32 24.3439
R2052 VP.n33 VP.n18 24.3439
R2053 VP.n26 VP.n25 24.3439
R2054 VP.n64 VP.n9 18.5015
R2055 VP.n78 VP.n3 18.5015
R2056 VP.n39 VP.n16 18.5015
R2057 VP.n25 VP.n22 18.5015
R2058 VP.n54 VP.n53 12.6591
R2059 VP.n89 VP.n88 12.6591
R2060 VP.n50 VP.n49 12.6591
R2061 VP.n24 VP.n23 6.69844
R2062 VP.n61 VP.n9 5.84292
R2063 VP.n81 VP.n3 5.84292
R2064 VP.n42 VP.n16 5.84292
R2065 VP.n51 VP.n13 0.278398
R2066 VP.n52 VP.n12 0.278398
R2067 VP.n90 VP.n0 0.278398
R2068 VP.n24 VP.n21 0.189894
R2069 VP.n28 VP.n21 0.189894
R2070 VP.n29 VP.n28 0.189894
R2071 VP.n30 VP.n29 0.189894
R2072 VP.n30 VP.n19 0.189894
R2073 VP.n34 VP.n19 0.189894
R2074 VP.n35 VP.n34 0.189894
R2075 VP.n36 VP.n35 0.189894
R2076 VP.n36 VP.n17 0.189894
R2077 VP.n40 VP.n17 0.189894
R2078 VP.n41 VP.n40 0.189894
R2079 VP.n41 VP.n15 0.189894
R2080 VP.n45 VP.n15 0.189894
R2081 VP.n46 VP.n45 0.189894
R2082 VP.n47 VP.n46 0.189894
R2083 VP.n47 VP.n13 0.189894
R2084 VP.n56 VP.n12 0.189894
R2085 VP.n57 VP.n56 0.189894
R2086 VP.n58 VP.n57 0.189894
R2087 VP.n58 VP.n10 0.189894
R2088 VP.n62 VP.n10 0.189894
R2089 VP.n63 VP.n62 0.189894
R2090 VP.n63 VP.n8 0.189894
R2091 VP.n67 VP.n8 0.189894
R2092 VP.n68 VP.n67 0.189894
R2093 VP.n69 VP.n68 0.189894
R2094 VP.n69 VP.n6 0.189894
R2095 VP.n73 VP.n6 0.189894
R2096 VP.n74 VP.n73 0.189894
R2097 VP.n75 VP.n74 0.189894
R2098 VP.n75 VP.n4 0.189894
R2099 VP.n79 VP.n4 0.189894
R2100 VP.n80 VP.n79 0.189894
R2101 VP.n80 VP.n2 0.189894
R2102 VP.n84 VP.n2 0.189894
R2103 VP.n85 VP.n84 0.189894
R2104 VP.n86 VP.n85 0.189894
R2105 VP.n86 VP.n0 0.189894
R2106 VP VP.n90 0.153422
R2107 VDD1.n1 VDD1.t2 69.9581
R2108 VDD1.n3 VDD1.t0 69.9579
R2109 VDD1.n5 VDD1.n4 67.3925
R2110 VDD1.n1 VDD1.n0 65.586
R2111 VDD1.n7 VDD1.n6 65.5859
R2112 VDD1.n3 VDD1.n2 65.5858
R2113 VDD1.n7 VDD1.n5 46.3673
R2114 VDD1.n6 VDD1.t8 1.88981
R2115 VDD1.n6 VDD1.t9 1.88981
R2116 VDD1.n0 VDD1.t3 1.88981
R2117 VDD1.n0 VDD1.t4 1.88981
R2118 VDD1.n4 VDD1.t1 1.88981
R2119 VDD1.n4 VDD1.t7 1.88981
R2120 VDD1.n2 VDD1.t5 1.88981
R2121 VDD1.n2 VDD1.t6 1.88981
R2122 VDD1 VDD1.n7 1.80438
R2123 VDD1 VDD1.n1 0.679379
R2124 VDD1.n5 VDD1.n3 0.565844
C0 VTAIL VP 10.0458f
C1 VTAIL VDD1 9.67635f
C2 VDD2 VP 0.57671f
C3 VDD2 VDD1 2.14141f
C4 VN VP 8.04785f
C5 VN VDD1 0.152877f
C6 VTAIL VDD2 9.727269f
C7 VTAIL VN 10.031599f
C8 VDD1 VP 9.76454f
C9 VN VDD2 9.344291f
C10 VDD2 B 6.899719f
C11 VDD1 B 6.859751f
C12 VTAIL B 7.564786f
C13 VN B 17.776161f
C14 VP B 16.328098f
C15 VDD1.t2 B 2.34548f
C16 VDD1.t3 B 0.206492f
C17 VDD1.t4 B 0.206492f
C18 VDD1.n0 B 1.82669f
C19 VDD1.n1 B 0.91102f
C20 VDD1.t0 B 2.34548f
C21 VDD1.t5 B 0.206492f
C22 VDD1.t6 B 0.206492f
C23 VDD1.n2 B 1.82669f
C24 VDD1.n3 B 0.902928f
C25 VDD1.t1 B 0.206492f
C26 VDD1.t7 B 0.206492f
C27 VDD1.n4 B 1.84161f
C28 VDD1.n5 B 2.89769f
C29 VDD1.t8 B 0.206492f
C30 VDD1.t9 B 0.206492f
C31 VDD1.n6 B 1.82669f
C32 VDD1.n7 B 3.02432f
C33 VP.n0 B 0.029541f
C34 VP.t2 B 1.62464f
C35 VP.n1 B 0.028449f
C36 VP.n2 B 0.022405f
C37 VP.t8 B 1.62464f
C38 VP.n3 B 0.580058f
C39 VP.n4 B 0.022405f
C40 VP.n5 B 0.042949f
C41 VP.n6 B 0.022405f
C42 VP.t3 B 1.62464f
C43 VP.n7 B 0.042949f
C44 VP.n8 B 0.022405f
C45 VP.t4 B 1.62464f
C46 VP.n9 B 0.580058f
C47 VP.n10 B 0.022405f
C48 VP.n11 B 0.028449f
C49 VP.n12 B 0.029541f
C50 VP.t9 B 1.62464f
C51 VP.n13 B 0.029541f
C52 VP.t0 B 1.62464f
C53 VP.n14 B 0.028449f
C54 VP.n15 B 0.022405f
C55 VP.t1 B 1.62464f
C56 VP.n16 B 0.580058f
C57 VP.n17 B 0.022405f
C58 VP.n18 B 0.042949f
C59 VP.n19 B 0.022405f
C60 VP.t5 B 1.62464f
C61 VP.n20 B 0.042949f
C62 VP.n21 B 0.022405f
C63 VP.t6 B 1.62464f
C64 VP.n22 B 0.650296f
C65 VP.t7 B 1.80951f
C66 VP.n23 B 0.623684f
C67 VP.n24 B 0.215447f
C68 VP.n25 B 0.036994f
C69 VP.n26 B 0.045522f
C70 VP.n27 B 0.019197f
C71 VP.n28 B 0.022405f
C72 VP.n29 B 0.022405f
C73 VP.n30 B 0.022405f
C74 VP.n31 B 0.041967f
C75 VP.n32 B 0.601305f
C76 VP.n33 B 0.041967f
C77 VP.n34 B 0.022405f
C78 VP.n35 B 0.022405f
C79 VP.n36 B 0.022405f
C80 VP.n37 B 0.019197f
C81 VP.n38 B 0.045522f
C82 VP.n39 B 0.036994f
C83 VP.n40 B 0.022405f
C84 VP.n41 B 0.022405f
C85 VP.n42 B 0.02622f
C86 VP.n43 B 0.041967f
C87 VP.n44 B 0.037252f
C88 VP.n45 B 0.022405f
C89 VP.n46 B 0.022405f
C90 VP.n47 B 0.022405f
C91 VP.n48 B 0.041967f
C92 VP.n49 B 0.032021f
C93 VP.n50 B 0.65772f
C94 VP.n51 B 1.3089f
C95 VP.n52 B 1.32442f
C96 VP.n53 B 0.65772f
C97 VP.n54 B 0.032021f
C98 VP.n55 B 0.041967f
C99 VP.n56 B 0.022405f
C100 VP.n57 B 0.022405f
C101 VP.n58 B 0.022405f
C102 VP.n59 B 0.037252f
C103 VP.n60 B 0.041967f
C104 VP.n61 B 0.02622f
C105 VP.n62 B 0.022405f
C106 VP.n63 B 0.022405f
C107 VP.n64 B 0.036994f
C108 VP.n65 B 0.045522f
C109 VP.n66 B 0.019197f
C110 VP.n67 B 0.022405f
C111 VP.n68 B 0.022405f
C112 VP.n69 B 0.022405f
C113 VP.n70 B 0.041967f
C114 VP.n71 B 0.601305f
C115 VP.n72 B 0.041967f
C116 VP.n73 B 0.022405f
C117 VP.n74 B 0.022405f
C118 VP.n75 B 0.022405f
C119 VP.n76 B 0.019197f
C120 VP.n77 B 0.045522f
C121 VP.n78 B 0.036994f
C122 VP.n79 B 0.022405f
C123 VP.n80 B 0.022405f
C124 VP.n81 B 0.02622f
C125 VP.n82 B 0.041967f
C126 VP.n83 B 0.037252f
C127 VP.n84 B 0.022405f
C128 VP.n85 B 0.022405f
C129 VP.n86 B 0.022405f
C130 VP.n87 B 0.041967f
C131 VP.n88 B 0.032021f
C132 VP.n89 B 0.65772f
C133 VP.n90 B 0.034472f
C134 VDD2.t9 B 2.30099f
C135 VDD2.t7 B 0.202576f
C136 VDD2.t3 B 0.202576f
C137 VDD2.n0 B 1.79205f
C138 VDD2.n1 B 0.885803f
C139 VDD2.t6 B 0.202576f
C140 VDD2.t2 B 0.202576f
C141 VDD2.n2 B 1.80668f
C142 VDD2.n3 B 2.72273f
C143 VDD2.t8 B 2.28455f
C144 VDD2.n4 B 2.91441f
C145 VDD2.t4 B 0.202576f
C146 VDD2.t5 B 0.202576f
C147 VDD2.n5 B 1.79205f
C148 VDD2.n6 B 0.446932f
C149 VDD2.t0 B 0.202576f
C150 VDD2.t1 B 0.202576f
C151 VDD2.n7 B 1.80664f
C152 VTAIL.t13 B 0.210307f
C153 VTAIL.t10 B 0.210307f
C154 VTAIL.n0 B 1.79208f
C155 VTAIL.n1 B 0.53628f
C156 VTAIL.t2 B 2.28547f
C157 VTAIL.n2 B 0.662474f
C158 VTAIL.t7 B 0.210307f
C159 VTAIL.t6 B 0.210307f
C160 VTAIL.n3 B 1.79208f
C161 VTAIL.n4 B 0.645441f
C162 VTAIL.t0 B 0.210307f
C163 VTAIL.t8 B 0.210307f
C164 VTAIL.n5 B 1.79208f
C165 VTAIL.n6 B 1.93281f
C166 VTAIL.t17 B 0.210307f
C167 VTAIL.t19 B 0.210307f
C168 VTAIL.n7 B 1.79208f
C169 VTAIL.n8 B 1.93281f
C170 VTAIL.t18 B 0.210307f
C171 VTAIL.t16 B 0.210307f
C172 VTAIL.n9 B 1.79208f
C173 VTAIL.n10 B 0.645436f
C174 VTAIL.t15 B 2.28548f
C175 VTAIL.n11 B 0.662468f
C176 VTAIL.t1 B 0.210307f
C177 VTAIL.t3 B 0.210307f
C178 VTAIL.n12 B 1.79208f
C179 VTAIL.n13 B 0.582302f
C180 VTAIL.t5 B 0.210307f
C181 VTAIL.t9 B 0.210307f
C182 VTAIL.n14 B 1.79208f
C183 VTAIL.n15 B 0.645436f
C184 VTAIL.t4 B 2.28547f
C185 VTAIL.n16 B 1.80982f
C186 VTAIL.t11 B 2.28547f
C187 VTAIL.n17 B 1.80982f
C188 VTAIL.t14 B 0.210307f
C189 VTAIL.t12 B 0.210307f
C190 VTAIL.n18 B 1.79208f
C191 VTAIL.n19 B 0.488313f
C192 VN.n0 B 0.028977f
C193 VN.t7 B 1.59362f
C194 VN.n1 B 0.027905f
C195 VN.n2 B 0.021978f
C196 VN.t3 B 1.59362f
C197 VN.n3 B 0.568981f
C198 VN.n4 B 0.021978f
C199 VN.n5 B 0.042129f
C200 VN.n6 B 0.021978f
C201 VN.t6 B 1.59362f
C202 VN.n7 B 0.042129f
C203 VN.n8 B 0.021978f
C204 VN.t2 B 1.59362f
C205 VN.n9 B 0.637877f
C206 VN.t0 B 1.77496f
C207 VN.n10 B 0.611773f
C208 VN.n11 B 0.211332f
C209 VN.n12 B 0.036288f
C210 VN.n13 B 0.044653f
C211 VN.n14 B 0.01883f
C212 VN.n15 B 0.021978f
C213 VN.n16 B 0.021978f
C214 VN.n17 B 0.021978f
C215 VN.n18 B 0.041166f
C216 VN.n19 B 0.589822f
C217 VN.n20 B 0.041166f
C218 VN.n21 B 0.021978f
C219 VN.n22 B 0.021978f
C220 VN.n23 B 0.021978f
C221 VN.n24 B 0.01883f
C222 VN.n25 B 0.044653f
C223 VN.n26 B 0.036288f
C224 VN.n27 B 0.021978f
C225 VN.n28 B 0.021978f
C226 VN.n29 B 0.025719f
C227 VN.n30 B 0.041166f
C228 VN.n31 B 0.03654f
C229 VN.n32 B 0.021978f
C230 VN.n33 B 0.021978f
C231 VN.n34 B 0.021978f
C232 VN.n35 B 0.041166f
C233 VN.n36 B 0.03141f
C234 VN.n37 B 0.645159f
C235 VN.n38 B 0.033813f
C236 VN.n39 B 0.028977f
C237 VN.t1 B 1.59362f
C238 VN.n40 B 0.027905f
C239 VN.n41 B 0.021978f
C240 VN.t5 B 1.59362f
C241 VN.n42 B 0.568981f
C242 VN.n43 B 0.021978f
C243 VN.n44 B 0.042129f
C244 VN.n45 B 0.021978f
C245 VN.t4 B 1.59362f
C246 VN.n46 B 0.042129f
C247 VN.n47 B 0.021978f
C248 VN.t9 B 1.59362f
C249 VN.n48 B 0.637877f
C250 VN.t8 B 1.77496f
C251 VN.n49 B 0.611773f
C252 VN.n50 B 0.211332f
C253 VN.n51 B 0.036288f
C254 VN.n52 B 0.044653f
C255 VN.n53 B 0.01883f
C256 VN.n54 B 0.021978f
C257 VN.n55 B 0.021978f
C258 VN.n56 B 0.021978f
C259 VN.n57 B 0.041166f
C260 VN.n58 B 0.589822f
C261 VN.n59 B 0.041166f
C262 VN.n60 B 0.021978f
C263 VN.n61 B 0.021978f
C264 VN.n62 B 0.021978f
C265 VN.n63 B 0.01883f
C266 VN.n64 B 0.044653f
C267 VN.n65 B 0.036288f
C268 VN.n66 B 0.021978f
C269 VN.n67 B 0.021978f
C270 VN.n68 B 0.025719f
C271 VN.n69 B 0.041166f
C272 VN.n70 B 0.03654f
C273 VN.n71 B 0.021978f
C274 VN.n72 B 0.021978f
C275 VN.n73 B 0.021978f
C276 VN.n74 B 0.041166f
C277 VN.n75 B 0.03141f
C278 VN.n76 B 0.645159f
C279 VN.n77 B 1.29565f
.ends

