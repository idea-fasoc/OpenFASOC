* NGSPICE file created from diff_pair_sample_1791.ext - technology: sky130A

.subckt diff_pair_sample_1791 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=1.3662 ps=8.61 w=8.28 l=0.17
X1 VTAIL.t14 VN.t1 VDD2.t2 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X2 VTAIL.t6 VP.t0 VDD1.t7 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=1.3662 ps=8.61 w=8.28 l=0.17
X3 B.t11 B.t9 B.t10 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=0 ps=0 w=8.28 l=0.17
X4 VDD1.t6 VP.t1 VTAIL.t5 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=3.2292 ps=17.34 w=8.28 l=0.17
X5 VDD2.t3 VN.t2 VTAIL.t13 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=3.2292 ps=17.34 w=8.28 l=0.17
X6 VTAIL.t3 VP.t2 VDD1.t5 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=1.3662 ps=8.61 w=8.28 l=0.17
X7 VDD1.t4 VP.t3 VTAIL.t4 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X8 VTAIL.t12 VN.t3 VDD2.t4 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=1.3662 ps=8.61 w=8.28 l=0.17
X9 B.t8 B.t6 B.t7 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=0 ps=0 w=8.28 l=0.17
X10 VTAIL.t2 VP.t4 VDD1.t3 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X11 B.t5 B.t3 B.t4 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=0 ps=0 w=8.28 l=0.17
X12 VTAIL.t1 VP.t5 VDD1.t2 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X13 VDD1.t1 VP.t6 VTAIL.t7 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=3.2292 ps=17.34 w=8.28 l=0.17
X14 B.t2 B.t0 B.t1 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=3.2292 pd=17.34 as=0 ps=0 w=8.28 l=0.17
X15 VDD2.t5 VN.t4 VTAIL.t11 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=3.2292 ps=17.34 w=8.28 l=0.17
X16 VDD2.t6 VN.t5 VTAIL.t10 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X17 VTAIL.t9 VN.t6 VDD2.t7 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X18 VDD1.t0 VP.t7 VTAIL.t0 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
X19 VDD2.t1 VN.t7 VTAIL.t8 w_n1470_n2624# sky130_fd_pr__pfet_01v8 ad=1.3662 pd=8.61 as=1.3662 ps=8.61 w=8.28 l=0.17
R0 VN.n5 VN.t4 1394.62
R1 VN.n1 VN.t0 1394.62
R2 VN.n12 VN.t3 1394.62
R3 VN.n8 VN.t2 1394.62
R4 VN.n4 VN.t6 1358.11
R5 VN.n2 VN.t7 1358.11
R6 VN.n11 VN.t5 1358.11
R7 VN.n9 VN.t1 1358.11
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN VN.n13 37.1009
R15 VN.n2 VN.n1 36.5157
R16 VN.n3 VN.n2 36.5157
R17 VN.n4 VN.n3 36.5157
R18 VN.n5 VN.n4 36.5157
R19 VN.n12 VN.n11 36.5157
R20 VN.n11 VN.n10 36.5157
R21 VN.n10 VN.n9 36.5157
R22 VN.n9 VN.n8 36.5157
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VDD2.n2 VDD2.n1 83.772
R27 VDD2.n2 VDD2.n0 83.772
R28 VDD2 VDD2.n5 83.7693
R29 VDD2.n4 VDD2.n3 83.6121
R30 VDD2.n4 VDD2.n2 32.7929
R31 VDD2.n5 VDD2.t2 3.92622
R32 VDD2.n5 VDD2.t3 3.92622
R33 VDD2.n3 VDD2.t4 3.92622
R34 VDD2.n3 VDD2.t6 3.92622
R35 VDD2.n1 VDD2.t7 3.92622
R36 VDD2.n1 VDD2.t5 3.92622
R37 VDD2.n0 VDD2.t0 3.92622
R38 VDD2.n0 VDD2.t1 3.92622
R39 VDD2 VDD2.n4 0.274207
R40 VTAIL.n11 VTAIL.t6 70.859
R41 VTAIL.n10 VTAIL.t13 70.859
R42 VTAIL.n7 VTAIL.t12 70.859
R43 VTAIL.n14 VTAIL.t5 70.8589
R44 VTAIL.n15 VTAIL.t11 70.8589
R45 VTAIL.n2 VTAIL.t15 70.8589
R46 VTAIL.n3 VTAIL.t7 70.8589
R47 VTAIL.n6 VTAIL.t3 70.8589
R48 VTAIL.n13 VTAIL.n12 66.9333
R49 VTAIL.n9 VTAIL.n8 66.9333
R50 VTAIL.n1 VTAIL.n0 66.9331
R51 VTAIL.n5 VTAIL.n4 66.9331
R52 VTAIL.n15 VTAIL.n14 19.9358
R53 VTAIL.n7 VTAIL.n6 19.9358
R54 VTAIL.n0 VTAIL.t8 3.92622
R55 VTAIL.n0 VTAIL.t9 3.92622
R56 VTAIL.n4 VTAIL.t4 3.92622
R57 VTAIL.n4 VTAIL.t2 3.92622
R58 VTAIL.n12 VTAIL.t0 3.92622
R59 VTAIL.n12 VTAIL.t1 3.92622
R60 VTAIL.n8 VTAIL.t10 3.92622
R61 VTAIL.n8 VTAIL.t14 3.92622
R62 VTAIL.n11 VTAIL.n10 0.470328
R63 VTAIL.n3 VTAIL.n2 0.470328
R64 VTAIL.n9 VTAIL.n7 0.431534
R65 VTAIL.n10 VTAIL.n9 0.431534
R66 VTAIL.n13 VTAIL.n11 0.431534
R67 VTAIL.n14 VTAIL.n13 0.431534
R68 VTAIL.n6 VTAIL.n5 0.431534
R69 VTAIL.n5 VTAIL.n3 0.431534
R70 VTAIL.n2 VTAIL.n1 0.431534
R71 VTAIL VTAIL.n15 0.373345
R72 VTAIL VTAIL.n1 0.0586897
R73 VP.n13 VP.t6 1394.62
R74 VP.n9 VP.t2 1394.62
R75 VP.n2 VP.t0 1394.62
R76 VP.n6 VP.t1 1394.62
R77 VP.n12 VP.t4 1358.11
R78 VP.n10 VP.t3 1358.11
R79 VP.n3 VP.t7 1358.11
R80 VP.n5 VP.t5 1358.11
R81 VP.n2 VP.n1 161.489
R82 VP.n14 VP.n13 161.3
R83 VP.n4 VP.n1 161.3
R84 VP.n7 VP.n6 161.3
R85 VP.n11 VP.n0 161.3
R86 VP.n9 VP.n8 161.3
R87 VP.n8 VP.n7 36.7202
R88 VP.n10 VP.n9 36.5157
R89 VP.n11 VP.n10 36.5157
R90 VP.n12 VP.n11 36.5157
R91 VP.n13 VP.n12 36.5157
R92 VP.n3 VP.n2 36.5157
R93 VP.n4 VP.n3 36.5157
R94 VP.n5 VP.n4 36.5157
R95 VP.n6 VP.n5 36.5157
R96 VP.n7 VP.n1 0.189894
R97 VP.n8 VP.n0 0.189894
R98 VP.n14 VP.n0 0.189894
R99 VP VP.n14 0.0516364
R100 VDD1 VDD1.n0 83.8858
R101 VDD1.n3 VDD1.n2 83.772
R102 VDD1.n3 VDD1.n1 83.772
R103 VDD1.n5 VDD1.n4 83.612
R104 VDD1.n5 VDD1.n3 33.3759
R105 VDD1.n4 VDD1.t2 3.92622
R106 VDD1.n4 VDD1.t6 3.92622
R107 VDD1.n0 VDD1.t7 3.92622
R108 VDD1.n0 VDD1.t0 3.92622
R109 VDD1.n2 VDD1.t3 3.92622
R110 VDD1.n2 VDD1.t1 3.92622
R111 VDD1.n1 VDD1.t5 3.92622
R112 VDD1.n1 VDD1.t4 3.92622
R113 VDD1 VDD1.n5 0.157828
R114 B.n86 B.t6 1420.79
R115 B.n190 B.t3 1420.79
R116 B.n32 B.t9 1420.79
R117 B.n26 B.t0 1420.79
R118 B.n240 B.n65 585
R119 B.n239 B.n238 585
R120 B.n237 B.n66 585
R121 B.n236 B.n235 585
R122 B.n234 B.n67 585
R123 B.n233 B.n232 585
R124 B.n231 B.n68 585
R125 B.n230 B.n229 585
R126 B.n228 B.n69 585
R127 B.n227 B.n226 585
R128 B.n225 B.n70 585
R129 B.n224 B.n223 585
R130 B.n222 B.n71 585
R131 B.n221 B.n220 585
R132 B.n219 B.n72 585
R133 B.n218 B.n217 585
R134 B.n216 B.n73 585
R135 B.n215 B.n214 585
R136 B.n213 B.n74 585
R137 B.n212 B.n211 585
R138 B.n210 B.n75 585
R139 B.n209 B.n208 585
R140 B.n207 B.n76 585
R141 B.n206 B.n205 585
R142 B.n204 B.n77 585
R143 B.n203 B.n202 585
R144 B.n201 B.n78 585
R145 B.n200 B.n199 585
R146 B.n198 B.n79 585
R147 B.n197 B.n196 585
R148 B.n195 B.n80 585
R149 B.n194 B.n193 585
R150 B.n189 B.n81 585
R151 B.n188 B.n187 585
R152 B.n186 B.n82 585
R153 B.n185 B.n184 585
R154 B.n183 B.n83 585
R155 B.n182 B.n181 585
R156 B.n180 B.n84 585
R157 B.n179 B.n178 585
R158 B.n176 B.n85 585
R159 B.n175 B.n174 585
R160 B.n173 B.n88 585
R161 B.n172 B.n171 585
R162 B.n170 B.n89 585
R163 B.n169 B.n168 585
R164 B.n167 B.n90 585
R165 B.n166 B.n165 585
R166 B.n164 B.n91 585
R167 B.n163 B.n162 585
R168 B.n161 B.n92 585
R169 B.n160 B.n159 585
R170 B.n158 B.n93 585
R171 B.n157 B.n156 585
R172 B.n155 B.n94 585
R173 B.n154 B.n153 585
R174 B.n152 B.n95 585
R175 B.n151 B.n150 585
R176 B.n149 B.n96 585
R177 B.n148 B.n147 585
R178 B.n146 B.n97 585
R179 B.n145 B.n144 585
R180 B.n143 B.n98 585
R181 B.n142 B.n141 585
R182 B.n140 B.n99 585
R183 B.n139 B.n138 585
R184 B.n137 B.n100 585
R185 B.n136 B.n135 585
R186 B.n134 B.n101 585
R187 B.n133 B.n132 585
R188 B.n131 B.n102 585
R189 B.n242 B.n241 585
R190 B.n243 B.n64 585
R191 B.n245 B.n244 585
R192 B.n246 B.n63 585
R193 B.n248 B.n247 585
R194 B.n249 B.n62 585
R195 B.n251 B.n250 585
R196 B.n252 B.n61 585
R197 B.n254 B.n253 585
R198 B.n255 B.n60 585
R199 B.n257 B.n256 585
R200 B.n258 B.n59 585
R201 B.n260 B.n259 585
R202 B.n261 B.n58 585
R203 B.n263 B.n262 585
R204 B.n264 B.n57 585
R205 B.n266 B.n265 585
R206 B.n267 B.n56 585
R207 B.n269 B.n268 585
R208 B.n270 B.n55 585
R209 B.n272 B.n271 585
R210 B.n273 B.n54 585
R211 B.n275 B.n274 585
R212 B.n276 B.n53 585
R213 B.n278 B.n277 585
R214 B.n279 B.n52 585
R215 B.n281 B.n280 585
R216 B.n282 B.n51 585
R217 B.n284 B.n283 585
R218 B.n285 B.n50 585
R219 B.n287 B.n286 585
R220 B.n288 B.n49 585
R221 B.n397 B.n396 585
R222 B.n395 B.n10 585
R223 B.n394 B.n393 585
R224 B.n392 B.n11 585
R225 B.n391 B.n390 585
R226 B.n389 B.n12 585
R227 B.n388 B.n387 585
R228 B.n386 B.n13 585
R229 B.n385 B.n384 585
R230 B.n383 B.n14 585
R231 B.n382 B.n381 585
R232 B.n380 B.n15 585
R233 B.n379 B.n378 585
R234 B.n377 B.n16 585
R235 B.n376 B.n375 585
R236 B.n374 B.n17 585
R237 B.n373 B.n372 585
R238 B.n371 B.n18 585
R239 B.n370 B.n369 585
R240 B.n368 B.n19 585
R241 B.n367 B.n366 585
R242 B.n365 B.n20 585
R243 B.n364 B.n363 585
R244 B.n362 B.n21 585
R245 B.n361 B.n360 585
R246 B.n359 B.n22 585
R247 B.n358 B.n357 585
R248 B.n356 B.n23 585
R249 B.n355 B.n354 585
R250 B.n353 B.n24 585
R251 B.n352 B.n351 585
R252 B.n349 B.n25 585
R253 B.n348 B.n347 585
R254 B.n346 B.n28 585
R255 B.n345 B.n344 585
R256 B.n343 B.n29 585
R257 B.n342 B.n341 585
R258 B.n340 B.n30 585
R259 B.n339 B.n338 585
R260 B.n337 B.n31 585
R261 B.n335 B.n334 585
R262 B.n333 B.n34 585
R263 B.n332 B.n331 585
R264 B.n330 B.n35 585
R265 B.n329 B.n328 585
R266 B.n327 B.n36 585
R267 B.n326 B.n325 585
R268 B.n324 B.n37 585
R269 B.n323 B.n322 585
R270 B.n321 B.n38 585
R271 B.n320 B.n319 585
R272 B.n318 B.n39 585
R273 B.n317 B.n316 585
R274 B.n315 B.n40 585
R275 B.n314 B.n313 585
R276 B.n312 B.n41 585
R277 B.n311 B.n310 585
R278 B.n309 B.n42 585
R279 B.n308 B.n307 585
R280 B.n306 B.n43 585
R281 B.n305 B.n304 585
R282 B.n303 B.n44 585
R283 B.n302 B.n301 585
R284 B.n300 B.n45 585
R285 B.n299 B.n298 585
R286 B.n297 B.n46 585
R287 B.n296 B.n295 585
R288 B.n294 B.n47 585
R289 B.n293 B.n292 585
R290 B.n291 B.n48 585
R291 B.n290 B.n289 585
R292 B.n398 B.n9 585
R293 B.n400 B.n399 585
R294 B.n401 B.n8 585
R295 B.n403 B.n402 585
R296 B.n404 B.n7 585
R297 B.n406 B.n405 585
R298 B.n407 B.n6 585
R299 B.n409 B.n408 585
R300 B.n410 B.n5 585
R301 B.n412 B.n411 585
R302 B.n413 B.n4 585
R303 B.n415 B.n414 585
R304 B.n416 B.n3 585
R305 B.n418 B.n417 585
R306 B.n419 B.n0 585
R307 B.n2 B.n1 585
R308 B.n110 B.n109 585
R309 B.n112 B.n111 585
R310 B.n113 B.n108 585
R311 B.n115 B.n114 585
R312 B.n116 B.n107 585
R313 B.n118 B.n117 585
R314 B.n119 B.n106 585
R315 B.n121 B.n120 585
R316 B.n122 B.n105 585
R317 B.n124 B.n123 585
R318 B.n125 B.n104 585
R319 B.n127 B.n126 585
R320 B.n128 B.n103 585
R321 B.n130 B.n129 585
R322 B.n131 B.n130 487.695
R323 B.n242 B.n65 487.695
R324 B.n290 B.n49 487.695
R325 B.n396 B.n9 487.695
R326 B.n421 B.n420 256.663
R327 B.n420 B.n419 235.042
R328 B.n420 B.n2 235.042
R329 B.n132 B.n131 163.367
R330 B.n132 B.n101 163.367
R331 B.n136 B.n101 163.367
R332 B.n137 B.n136 163.367
R333 B.n138 B.n137 163.367
R334 B.n138 B.n99 163.367
R335 B.n142 B.n99 163.367
R336 B.n143 B.n142 163.367
R337 B.n144 B.n143 163.367
R338 B.n144 B.n97 163.367
R339 B.n148 B.n97 163.367
R340 B.n149 B.n148 163.367
R341 B.n150 B.n149 163.367
R342 B.n150 B.n95 163.367
R343 B.n154 B.n95 163.367
R344 B.n155 B.n154 163.367
R345 B.n156 B.n155 163.367
R346 B.n156 B.n93 163.367
R347 B.n160 B.n93 163.367
R348 B.n161 B.n160 163.367
R349 B.n162 B.n161 163.367
R350 B.n162 B.n91 163.367
R351 B.n166 B.n91 163.367
R352 B.n167 B.n166 163.367
R353 B.n168 B.n167 163.367
R354 B.n168 B.n89 163.367
R355 B.n172 B.n89 163.367
R356 B.n173 B.n172 163.367
R357 B.n174 B.n173 163.367
R358 B.n174 B.n85 163.367
R359 B.n179 B.n85 163.367
R360 B.n180 B.n179 163.367
R361 B.n181 B.n180 163.367
R362 B.n181 B.n83 163.367
R363 B.n185 B.n83 163.367
R364 B.n186 B.n185 163.367
R365 B.n187 B.n186 163.367
R366 B.n187 B.n81 163.367
R367 B.n194 B.n81 163.367
R368 B.n195 B.n194 163.367
R369 B.n196 B.n195 163.367
R370 B.n196 B.n79 163.367
R371 B.n200 B.n79 163.367
R372 B.n201 B.n200 163.367
R373 B.n202 B.n201 163.367
R374 B.n202 B.n77 163.367
R375 B.n206 B.n77 163.367
R376 B.n207 B.n206 163.367
R377 B.n208 B.n207 163.367
R378 B.n208 B.n75 163.367
R379 B.n212 B.n75 163.367
R380 B.n213 B.n212 163.367
R381 B.n214 B.n213 163.367
R382 B.n214 B.n73 163.367
R383 B.n218 B.n73 163.367
R384 B.n219 B.n218 163.367
R385 B.n220 B.n219 163.367
R386 B.n220 B.n71 163.367
R387 B.n224 B.n71 163.367
R388 B.n225 B.n224 163.367
R389 B.n226 B.n225 163.367
R390 B.n226 B.n69 163.367
R391 B.n230 B.n69 163.367
R392 B.n231 B.n230 163.367
R393 B.n232 B.n231 163.367
R394 B.n232 B.n67 163.367
R395 B.n236 B.n67 163.367
R396 B.n237 B.n236 163.367
R397 B.n238 B.n237 163.367
R398 B.n238 B.n65 163.367
R399 B.n286 B.n49 163.367
R400 B.n286 B.n285 163.367
R401 B.n285 B.n284 163.367
R402 B.n284 B.n51 163.367
R403 B.n280 B.n51 163.367
R404 B.n280 B.n279 163.367
R405 B.n279 B.n278 163.367
R406 B.n278 B.n53 163.367
R407 B.n274 B.n53 163.367
R408 B.n274 B.n273 163.367
R409 B.n273 B.n272 163.367
R410 B.n272 B.n55 163.367
R411 B.n268 B.n55 163.367
R412 B.n268 B.n267 163.367
R413 B.n267 B.n266 163.367
R414 B.n266 B.n57 163.367
R415 B.n262 B.n57 163.367
R416 B.n262 B.n261 163.367
R417 B.n261 B.n260 163.367
R418 B.n260 B.n59 163.367
R419 B.n256 B.n59 163.367
R420 B.n256 B.n255 163.367
R421 B.n255 B.n254 163.367
R422 B.n254 B.n61 163.367
R423 B.n250 B.n61 163.367
R424 B.n250 B.n249 163.367
R425 B.n249 B.n248 163.367
R426 B.n248 B.n63 163.367
R427 B.n244 B.n63 163.367
R428 B.n244 B.n243 163.367
R429 B.n243 B.n242 163.367
R430 B.n396 B.n395 163.367
R431 B.n395 B.n394 163.367
R432 B.n394 B.n11 163.367
R433 B.n390 B.n11 163.367
R434 B.n390 B.n389 163.367
R435 B.n389 B.n388 163.367
R436 B.n388 B.n13 163.367
R437 B.n384 B.n13 163.367
R438 B.n384 B.n383 163.367
R439 B.n383 B.n382 163.367
R440 B.n382 B.n15 163.367
R441 B.n378 B.n15 163.367
R442 B.n378 B.n377 163.367
R443 B.n377 B.n376 163.367
R444 B.n376 B.n17 163.367
R445 B.n372 B.n17 163.367
R446 B.n372 B.n371 163.367
R447 B.n371 B.n370 163.367
R448 B.n370 B.n19 163.367
R449 B.n366 B.n19 163.367
R450 B.n366 B.n365 163.367
R451 B.n365 B.n364 163.367
R452 B.n364 B.n21 163.367
R453 B.n360 B.n21 163.367
R454 B.n360 B.n359 163.367
R455 B.n359 B.n358 163.367
R456 B.n358 B.n23 163.367
R457 B.n354 B.n23 163.367
R458 B.n354 B.n353 163.367
R459 B.n353 B.n352 163.367
R460 B.n352 B.n25 163.367
R461 B.n347 B.n25 163.367
R462 B.n347 B.n346 163.367
R463 B.n346 B.n345 163.367
R464 B.n345 B.n29 163.367
R465 B.n341 B.n29 163.367
R466 B.n341 B.n340 163.367
R467 B.n340 B.n339 163.367
R468 B.n339 B.n31 163.367
R469 B.n334 B.n31 163.367
R470 B.n334 B.n333 163.367
R471 B.n333 B.n332 163.367
R472 B.n332 B.n35 163.367
R473 B.n328 B.n35 163.367
R474 B.n328 B.n327 163.367
R475 B.n327 B.n326 163.367
R476 B.n326 B.n37 163.367
R477 B.n322 B.n37 163.367
R478 B.n322 B.n321 163.367
R479 B.n321 B.n320 163.367
R480 B.n320 B.n39 163.367
R481 B.n316 B.n39 163.367
R482 B.n316 B.n315 163.367
R483 B.n315 B.n314 163.367
R484 B.n314 B.n41 163.367
R485 B.n310 B.n41 163.367
R486 B.n310 B.n309 163.367
R487 B.n309 B.n308 163.367
R488 B.n308 B.n43 163.367
R489 B.n304 B.n43 163.367
R490 B.n304 B.n303 163.367
R491 B.n303 B.n302 163.367
R492 B.n302 B.n45 163.367
R493 B.n298 B.n45 163.367
R494 B.n298 B.n297 163.367
R495 B.n297 B.n296 163.367
R496 B.n296 B.n47 163.367
R497 B.n292 B.n47 163.367
R498 B.n292 B.n291 163.367
R499 B.n291 B.n290 163.367
R500 B.n400 B.n9 163.367
R501 B.n401 B.n400 163.367
R502 B.n402 B.n401 163.367
R503 B.n402 B.n7 163.367
R504 B.n406 B.n7 163.367
R505 B.n407 B.n406 163.367
R506 B.n408 B.n407 163.367
R507 B.n408 B.n5 163.367
R508 B.n412 B.n5 163.367
R509 B.n413 B.n412 163.367
R510 B.n414 B.n413 163.367
R511 B.n414 B.n3 163.367
R512 B.n418 B.n3 163.367
R513 B.n419 B.n418 163.367
R514 B.n109 B.n2 163.367
R515 B.n112 B.n109 163.367
R516 B.n113 B.n112 163.367
R517 B.n114 B.n113 163.367
R518 B.n114 B.n107 163.367
R519 B.n118 B.n107 163.367
R520 B.n119 B.n118 163.367
R521 B.n120 B.n119 163.367
R522 B.n120 B.n105 163.367
R523 B.n124 B.n105 163.367
R524 B.n125 B.n124 163.367
R525 B.n126 B.n125 163.367
R526 B.n126 B.n103 163.367
R527 B.n130 B.n103 163.367
R528 B.n190 B.t4 120.511
R529 B.n32 B.t11 120.511
R530 B.n86 B.t7 120.502
R531 B.n26 B.t2 120.502
R532 B.n191 B.t5 110.814
R533 B.n33 B.t10 110.814
R534 B.n87 B.t8 110.805
R535 B.n27 B.t1 110.805
R536 B.n177 B.n87 59.5399
R537 B.n192 B.n191 59.5399
R538 B.n336 B.n33 59.5399
R539 B.n350 B.n27 59.5399
R540 B.n398 B.n397 31.6883
R541 B.n289 B.n288 31.6883
R542 B.n241 B.n240 31.6883
R543 B.n129 B.n102 31.6883
R544 B B.n421 18.0485
R545 B.n399 B.n398 10.6151
R546 B.n399 B.n8 10.6151
R547 B.n403 B.n8 10.6151
R548 B.n404 B.n403 10.6151
R549 B.n405 B.n404 10.6151
R550 B.n405 B.n6 10.6151
R551 B.n409 B.n6 10.6151
R552 B.n410 B.n409 10.6151
R553 B.n411 B.n410 10.6151
R554 B.n411 B.n4 10.6151
R555 B.n415 B.n4 10.6151
R556 B.n416 B.n415 10.6151
R557 B.n417 B.n416 10.6151
R558 B.n417 B.n0 10.6151
R559 B.n397 B.n10 10.6151
R560 B.n393 B.n10 10.6151
R561 B.n393 B.n392 10.6151
R562 B.n392 B.n391 10.6151
R563 B.n391 B.n12 10.6151
R564 B.n387 B.n12 10.6151
R565 B.n387 B.n386 10.6151
R566 B.n386 B.n385 10.6151
R567 B.n385 B.n14 10.6151
R568 B.n381 B.n14 10.6151
R569 B.n381 B.n380 10.6151
R570 B.n380 B.n379 10.6151
R571 B.n379 B.n16 10.6151
R572 B.n375 B.n16 10.6151
R573 B.n375 B.n374 10.6151
R574 B.n374 B.n373 10.6151
R575 B.n373 B.n18 10.6151
R576 B.n369 B.n18 10.6151
R577 B.n369 B.n368 10.6151
R578 B.n368 B.n367 10.6151
R579 B.n367 B.n20 10.6151
R580 B.n363 B.n20 10.6151
R581 B.n363 B.n362 10.6151
R582 B.n362 B.n361 10.6151
R583 B.n361 B.n22 10.6151
R584 B.n357 B.n22 10.6151
R585 B.n357 B.n356 10.6151
R586 B.n356 B.n355 10.6151
R587 B.n355 B.n24 10.6151
R588 B.n351 B.n24 10.6151
R589 B.n349 B.n348 10.6151
R590 B.n348 B.n28 10.6151
R591 B.n344 B.n28 10.6151
R592 B.n344 B.n343 10.6151
R593 B.n343 B.n342 10.6151
R594 B.n342 B.n30 10.6151
R595 B.n338 B.n30 10.6151
R596 B.n338 B.n337 10.6151
R597 B.n335 B.n34 10.6151
R598 B.n331 B.n34 10.6151
R599 B.n331 B.n330 10.6151
R600 B.n330 B.n329 10.6151
R601 B.n329 B.n36 10.6151
R602 B.n325 B.n36 10.6151
R603 B.n325 B.n324 10.6151
R604 B.n324 B.n323 10.6151
R605 B.n323 B.n38 10.6151
R606 B.n319 B.n38 10.6151
R607 B.n319 B.n318 10.6151
R608 B.n318 B.n317 10.6151
R609 B.n317 B.n40 10.6151
R610 B.n313 B.n40 10.6151
R611 B.n313 B.n312 10.6151
R612 B.n312 B.n311 10.6151
R613 B.n311 B.n42 10.6151
R614 B.n307 B.n42 10.6151
R615 B.n307 B.n306 10.6151
R616 B.n306 B.n305 10.6151
R617 B.n305 B.n44 10.6151
R618 B.n301 B.n44 10.6151
R619 B.n301 B.n300 10.6151
R620 B.n300 B.n299 10.6151
R621 B.n299 B.n46 10.6151
R622 B.n295 B.n46 10.6151
R623 B.n295 B.n294 10.6151
R624 B.n294 B.n293 10.6151
R625 B.n293 B.n48 10.6151
R626 B.n289 B.n48 10.6151
R627 B.n288 B.n287 10.6151
R628 B.n287 B.n50 10.6151
R629 B.n283 B.n50 10.6151
R630 B.n283 B.n282 10.6151
R631 B.n282 B.n281 10.6151
R632 B.n281 B.n52 10.6151
R633 B.n277 B.n52 10.6151
R634 B.n277 B.n276 10.6151
R635 B.n276 B.n275 10.6151
R636 B.n275 B.n54 10.6151
R637 B.n271 B.n54 10.6151
R638 B.n271 B.n270 10.6151
R639 B.n270 B.n269 10.6151
R640 B.n269 B.n56 10.6151
R641 B.n265 B.n56 10.6151
R642 B.n265 B.n264 10.6151
R643 B.n264 B.n263 10.6151
R644 B.n263 B.n58 10.6151
R645 B.n259 B.n58 10.6151
R646 B.n259 B.n258 10.6151
R647 B.n258 B.n257 10.6151
R648 B.n257 B.n60 10.6151
R649 B.n253 B.n60 10.6151
R650 B.n253 B.n252 10.6151
R651 B.n252 B.n251 10.6151
R652 B.n251 B.n62 10.6151
R653 B.n247 B.n62 10.6151
R654 B.n247 B.n246 10.6151
R655 B.n246 B.n245 10.6151
R656 B.n245 B.n64 10.6151
R657 B.n241 B.n64 10.6151
R658 B.n110 B.n1 10.6151
R659 B.n111 B.n110 10.6151
R660 B.n111 B.n108 10.6151
R661 B.n115 B.n108 10.6151
R662 B.n116 B.n115 10.6151
R663 B.n117 B.n116 10.6151
R664 B.n117 B.n106 10.6151
R665 B.n121 B.n106 10.6151
R666 B.n122 B.n121 10.6151
R667 B.n123 B.n122 10.6151
R668 B.n123 B.n104 10.6151
R669 B.n127 B.n104 10.6151
R670 B.n128 B.n127 10.6151
R671 B.n129 B.n128 10.6151
R672 B.n133 B.n102 10.6151
R673 B.n134 B.n133 10.6151
R674 B.n135 B.n134 10.6151
R675 B.n135 B.n100 10.6151
R676 B.n139 B.n100 10.6151
R677 B.n140 B.n139 10.6151
R678 B.n141 B.n140 10.6151
R679 B.n141 B.n98 10.6151
R680 B.n145 B.n98 10.6151
R681 B.n146 B.n145 10.6151
R682 B.n147 B.n146 10.6151
R683 B.n147 B.n96 10.6151
R684 B.n151 B.n96 10.6151
R685 B.n152 B.n151 10.6151
R686 B.n153 B.n152 10.6151
R687 B.n153 B.n94 10.6151
R688 B.n157 B.n94 10.6151
R689 B.n158 B.n157 10.6151
R690 B.n159 B.n158 10.6151
R691 B.n159 B.n92 10.6151
R692 B.n163 B.n92 10.6151
R693 B.n164 B.n163 10.6151
R694 B.n165 B.n164 10.6151
R695 B.n165 B.n90 10.6151
R696 B.n169 B.n90 10.6151
R697 B.n170 B.n169 10.6151
R698 B.n171 B.n170 10.6151
R699 B.n171 B.n88 10.6151
R700 B.n175 B.n88 10.6151
R701 B.n176 B.n175 10.6151
R702 B.n178 B.n84 10.6151
R703 B.n182 B.n84 10.6151
R704 B.n183 B.n182 10.6151
R705 B.n184 B.n183 10.6151
R706 B.n184 B.n82 10.6151
R707 B.n188 B.n82 10.6151
R708 B.n189 B.n188 10.6151
R709 B.n193 B.n189 10.6151
R710 B.n197 B.n80 10.6151
R711 B.n198 B.n197 10.6151
R712 B.n199 B.n198 10.6151
R713 B.n199 B.n78 10.6151
R714 B.n203 B.n78 10.6151
R715 B.n204 B.n203 10.6151
R716 B.n205 B.n204 10.6151
R717 B.n205 B.n76 10.6151
R718 B.n209 B.n76 10.6151
R719 B.n210 B.n209 10.6151
R720 B.n211 B.n210 10.6151
R721 B.n211 B.n74 10.6151
R722 B.n215 B.n74 10.6151
R723 B.n216 B.n215 10.6151
R724 B.n217 B.n216 10.6151
R725 B.n217 B.n72 10.6151
R726 B.n221 B.n72 10.6151
R727 B.n222 B.n221 10.6151
R728 B.n223 B.n222 10.6151
R729 B.n223 B.n70 10.6151
R730 B.n227 B.n70 10.6151
R731 B.n228 B.n227 10.6151
R732 B.n229 B.n228 10.6151
R733 B.n229 B.n68 10.6151
R734 B.n233 B.n68 10.6151
R735 B.n234 B.n233 10.6151
R736 B.n235 B.n234 10.6151
R737 B.n235 B.n66 10.6151
R738 B.n239 B.n66 10.6151
R739 B.n240 B.n239 10.6151
R740 B.n87 B.n86 9.69747
R741 B.n191 B.n190 9.69747
R742 B.n33 B.n32 9.69747
R743 B.n27 B.n26 9.69747
R744 B.n421 B.n0 8.11757
R745 B.n421 B.n1 8.11757
R746 B.n350 B.n349 6.5566
R747 B.n337 B.n336 6.5566
R748 B.n178 B.n177 6.5566
R749 B.n193 B.n192 6.5566
R750 B.n351 B.n350 4.05904
R751 B.n336 B.n335 4.05904
R752 B.n177 B.n176 4.05904
R753 B.n192 B.n80 4.05904
C0 VP VTAIL 1.4035f
C1 VP VDD1 1.85669f
C2 VP VN 4.00224f
C3 VDD2 B 0.828565f
C4 VDD2 w_n1470_n2624# 0.982738f
C5 VDD2 VTAIL 14.896599f
C6 VDD2 VDD1 0.568086f
C7 VDD2 VN 1.7431f
C8 w_n1470_n2624# B 5.42693f
C9 VTAIL B 2.46893f
C10 B VDD1 0.80767f
C11 VTAIL w_n1470_n2624# 3.32731f
C12 w_n1470_n2624# VDD1 0.969281f
C13 VTAIL VDD1 14.8585f
C14 VN B 0.612016f
C15 VP VDD2 0.260852f
C16 VN w_n1470_n2624# 2.25513f
C17 VN VTAIL 1.38939f
C18 VN VDD1 0.147094f
C19 VP B 0.906961f
C20 VP w_n1470_n2624# 2.4388f
C21 VDD2 VSUBS 1.212402f
C22 VDD1 VSUBS 1.405804f
C23 VTAIL VSUBS 0.520587f
C24 VN VSUBS 3.28143f
C25 VP VSUBS 0.961335f
C26 B VSUBS 1.967321f
C27 w_n1470_n2624# VSUBS 47.822f
C28 B.n0 VSUBS 0.008242f
C29 B.n1 VSUBS 0.008242f
C30 B.n2 VSUBS 0.01219f
C31 B.n3 VSUBS 0.009341f
C32 B.n4 VSUBS 0.009341f
C33 B.n5 VSUBS 0.009341f
C34 B.n6 VSUBS 0.009341f
C35 B.n7 VSUBS 0.009341f
C36 B.n8 VSUBS 0.009341f
C37 B.n9 VSUBS 0.020889f
C38 B.n10 VSUBS 0.009341f
C39 B.n11 VSUBS 0.009341f
C40 B.n12 VSUBS 0.009341f
C41 B.n13 VSUBS 0.009341f
C42 B.n14 VSUBS 0.009341f
C43 B.n15 VSUBS 0.009341f
C44 B.n16 VSUBS 0.009341f
C45 B.n17 VSUBS 0.009341f
C46 B.n18 VSUBS 0.009341f
C47 B.n19 VSUBS 0.009341f
C48 B.n20 VSUBS 0.009341f
C49 B.n21 VSUBS 0.009341f
C50 B.n22 VSUBS 0.009341f
C51 B.n23 VSUBS 0.009341f
C52 B.n24 VSUBS 0.009341f
C53 B.n25 VSUBS 0.009341f
C54 B.t1 VSUBS 0.34288f
C55 B.t2 VSUBS 0.348397f
C56 B.t0 VSUBS 0.07323f
C57 B.n26 VSUBS 0.096954f
C58 B.n27 VSUBS 0.081874f
C59 B.n28 VSUBS 0.009341f
C60 B.n29 VSUBS 0.009341f
C61 B.n30 VSUBS 0.009341f
C62 B.n31 VSUBS 0.009341f
C63 B.t10 VSUBS 0.342877f
C64 B.t11 VSUBS 0.348393f
C65 B.t9 VSUBS 0.07323f
C66 B.n32 VSUBS 0.096957f
C67 B.n33 VSUBS 0.081877f
C68 B.n34 VSUBS 0.009341f
C69 B.n35 VSUBS 0.009341f
C70 B.n36 VSUBS 0.009341f
C71 B.n37 VSUBS 0.009341f
C72 B.n38 VSUBS 0.009341f
C73 B.n39 VSUBS 0.009341f
C74 B.n40 VSUBS 0.009341f
C75 B.n41 VSUBS 0.009341f
C76 B.n42 VSUBS 0.009341f
C77 B.n43 VSUBS 0.009341f
C78 B.n44 VSUBS 0.009341f
C79 B.n45 VSUBS 0.009341f
C80 B.n46 VSUBS 0.009341f
C81 B.n47 VSUBS 0.009341f
C82 B.n48 VSUBS 0.009341f
C83 B.n49 VSUBS 0.020889f
C84 B.n50 VSUBS 0.009341f
C85 B.n51 VSUBS 0.009341f
C86 B.n52 VSUBS 0.009341f
C87 B.n53 VSUBS 0.009341f
C88 B.n54 VSUBS 0.009341f
C89 B.n55 VSUBS 0.009341f
C90 B.n56 VSUBS 0.009341f
C91 B.n57 VSUBS 0.009341f
C92 B.n58 VSUBS 0.009341f
C93 B.n59 VSUBS 0.009341f
C94 B.n60 VSUBS 0.009341f
C95 B.n61 VSUBS 0.009341f
C96 B.n62 VSUBS 0.009341f
C97 B.n63 VSUBS 0.009341f
C98 B.n64 VSUBS 0.009341f
C99 B.n65 VSUBS 0.021971f
C100 B.n66 VSUBS 0.009341f
C101 B.n67 VSUBS 0.009341f
C102 B.n68 VSUBS 0.009341f
C103 B.n69 VSUBS 0.009341f
C104 B.n70 VSUBS 0.009341f
C105 B.n71 VSUBS 0.009341f
C106 B.n72 VSUBS 0.009341f
C107 B.n73 VSUBS 0.009341f
C108 B.n74 VSUBS 0.009341f
C109 B.n75 VSUBS 0.009341f
C110 B.n76 VSUBS 0.009341f
C111 B.n77 VSUBS 0.009341f
C112 B.n78 VSUBS 0.009341f
C113 B.n79 VSUBS 0.009341f
C114 B.n80 VSUBS 0.006456f
C115 B.n81 VSUBS 0.009341f
C116 B.n82 VSUBS 0.009341f
C117 B.n83 VSUBS 0.009341f
C118 B.n84 VSUBS 0.009341f
C119 B.n85 VSUBS 0.009341f
C120 B.t8 VSUBS 0.34288f
C121 B.t7 VSUBS 0.348397f
C122 B.t6 VSUBS 0.07323f
C123 B.n86 VSUBS 0.096954f
C124 B.n87 VSUBS 0.081874f
C125 B.n88 VSUBS 0.009341f
C126 B.n89 VSUBS 0.009341f
C127 B.n90 VSUBS 0.009341f
C128 B.n91 VSUBS 0.009341f
C129 B.n92 VSUBS 0.009341f
C130 B.n93 VSUBS 0.009341f
C131 B.n94 VSUBS 0.009341f
C132 B.n95 VSUBS 0.009341f
C133 B.n96 VSUBS 0.009341f
C134 B.n97 VSUBS 0.009341f
C135 B.n98 VSUBS 0.009341f
C136 B.n99 VSUBS 0.009341f
C137 B.n100 VSUBS 0.009341f
C138 B.n101 VSUBS 0.009341f
C139 B.n102 VSUBS 0.021971f
C140 B.n103 VSUBS 0.009341f
C141 B.n104 VSUBS 0.009341f
C142 B.n105 VSUBS 0.009341f
C143 B.n106 VSUBS 0.009341f
C144 B.n107 VSUBS 0.009341f
C145 B.n108 VSUBS 0.009341f
C146 B.n109 VSUBS 0.009341f
C147 B.n110 VSUBS 0.009341f
C148 B.n111 VSUBS 0.009341f
C149 B.n112 VSUBS 0.009341f
C150 B.n113 VSUBS 0.009341f
C151 B.n114 VSUBS 0.009341f
C152 B.n115 VSUBS 0.009341f
C153 B.n116 VSUBS 0.009341f
C154 B.n117 VSUBS 0.009341f
C155 B.n118 VSUBS 0.009341f
C156 B.n119 VSUBS 0.009341f
C157 B.n120 VSUBS 0.009341f
C158 B.n121 VSUBS 0.009341f
C159 B.n122 VSUBS 0.009341f
C160 B.n123 VSUBS 0.009341f
C161 B.n124 VSUBS 0.009341f
C162 B.n125 VSUBS 0.009341f
C163 B.n126 VSUBS 0.009341f
C164 B.n127 VSUBS 0.009341f
C165 B.n128 VSUBS 0.009341f
C166 B.n129 VSUBS 0.020889f
C167 B.n130 VSUBS 0.020889f
C168 B.n131 VSUBS 0.021971f
C169 B.n132 VSUBS 0.009341f
C170 B.n133 VSUBS 0.009341f
C171 B.n134 VSUBS 0.009341f
C172 B.n135 VSUBS 0.009341f
C173 B.n136 VSUBS 0.009341f
C174 B.n137 VSUBS 0.009341f
C175 B.n138 VSUBS 0.009341f
C176 B.n139 VSUBS 0.009341f
C177 B.n140 VSUBS 0.009341f
C178 B.n141 VSUBS 0.009341f
C179 B.n142 VSUBS 0.009341f
C180 B.n143 VSUBS 0.009341f
C181 B.n144 VSUBS 0.009341f
C182 B.n145 VSUBS 0.009341f
C183 B.n146 VSUBS 0.009341f
C184 B.n147 VSUBS 0.009341f
C185 B.n148 VSUBS 0.009341f
C186 B.n149 VSUBS 0.009341f
C187 B.n150 VSUBS 0.009341f
C188 B.n151 VSUBS 0.009341f
C189 B.n152 VSUBS 0.009341f
C190 B.n153 VSUBS 0.009341f
C191 B.n154 VSUBS 0.009341f
C192 B.n155 VSUBS 0.009341f
C193 B.n156 VSUBS 0.009341f
C194 B.n157 VSUBS 0.009341f
C195 B.n158 VSUBS 0.009341f
C196 B.n159 VSUBS 0.009341f
C197 B.n160 VSUBS 0.009341f
C198 B.n161 VSUBS 0.009341f
C199 B.n162 VSUBS 0.009341f
C200 B.n163 VSUBS 0.009341f
C201 B.n164 VSUBS 0.009341f
C202 B.n165 VSUBS 0.009341f
C203 B.n166 VSUBS 0.009341f
C204 B.n167 VSUBS 0.009341f
C205 B.n168 VSUBS 0.009341f
C206 B.n169 VSUBS 0.009341f
C207 B.n170 VSUBS 0.009341f
C208 B.n171 VSUBS 0.009341f
C209 B.n172 VSUBS 0.009341f
C210 B.n173 VSUBS 0.009341f
C211 B.n174 VSUBS 0.009341f
C212 B.n175 VSUBS 0.009341f
C213 B.n176 VSUBS 0.006456f
C214 B.n177 VSUBS 0.021643f
C215 B.n178 VSUBS 0.007555f
C216 B.n179 VSUBS 0.009341f
C217 B.n180 VSUBS 0.009341f
C218 B.n181 VSUBS 0.009341f
C219 B.n182 VSUBS 0.009341f
C220 B.n183 VSUBS 0.009341f
C221 B.n184 VSUBS 0.009341f
C222 B.n185 VSUBS 0.009341f
C223 B.n186 VSUBS 0.009341f
C224 B.n187 VSUBS 0.009341f
C225 B.n188 VSUBS 0.009341f
C226 B.n189 VSUBS 0.009341f
C227 B.t5 VSUBS 0.342877f
C228 B.t4 VSUBS 0.348393f
C229 B.t3 VSUBS 0.07323f
C230 B.n190 VSUBS 0.096957f
C231 B.n191 VSUBS 0.081877f
C232 B.n192 VSUBS 0.021643f
C233 B.n193 VSUBS 0.007555f
C234 B.n194 VSUBS 0.009341f
C235 B.n195 VSUBS 0.009341f
C236 B.n196 VSUBS 0.009341f
C237 B.n197 VSUBS 0.009341f
C238 B.n198 VSUBS 0.009341f
C239 B.n199 VSUBS 0.009341f
C240 B.n200 VSUBS 0.009341f
C241 B.n201 VSUBS 0.009341f
C242 B.n202 VSUBS 0.009341f
C243 B.n203 VSUBS 0.009341f
C244 B.n204 VSUBS 0.009341f
C245 B.n205 VSUBS 0.009341f
C246 B.n206 VSUBS 0.009341f
C247 B.n207 VSUBS 0.009341f
C248 B.n208 VSUBS 0.009341f
C249 B.n209 VSUBS 0.009341f
C250 B.n210 VSUBS 0.009341f
C251 B.n211 VSUBS 0.009341f
C252 B.n212 VSUBS 0.009341f
C253 B.n213 VSUBS 0.009341f
C254 B.n214 VSUBS 0.009341f
C255 B.n215 VSUBS 0.009341f
C256 B.n216 VSUBS 0.009341f
C257 B.n217 VSUBS 0.009341f
C258 B.n218 VSUBS 0.009341f
C259 B.n219 VSUBS 0.009341f
C260 B.n220 VSUBS 0.009341f
C261 B.n221 VSUBS 0.009341f
C262 B.n222 VSUBS 0.009341f
C263 B.n223 VSUBS 0.009341f
C264 B.n224 VSUBS 0.009341f
C265 B.n225 VSUBS 0.009341f
C266 B.n226 VSUBS 0.009341f
C267 B.n227 VSUBS 0.009341f
C268 B.n228 VSUBS 0.009341f
C269 B.n229 VSUBS 0.009341f
C270 B.n230 VSUBS 0.009341f
C271 B.n231 VSUBS 0.009341f
C272 B.n232 VSUBS 0.009341f
C273 B.n233 VSUBS 0.009341f
C274 B.n234 VSUBS 0.009341f
C275 B.n235 VSUBS 0.009341f
C276 B.n236 VSUBS 0.009341f
C277 B.n237 VSUBS 0.009341f
C278 B.n238 VSUBS 0.009341f
C279 B.n239 VSUBS 0.009341f
C280 B.n240 VSUBS 0.020833f
C281 B.n241 VSUBS 0.022027f
C282 B.n242 VSUBS 0.020889f
C283 B.n243 VSUBS 0.009341f
C284 B.n244 VSUBS 0.009341f
C285 B.n245 VSUBS 0.009341f
C286 B.n246 VSUBS 0.009341f
C287 B.n247 VSUBS 0.009341f
C288 B.n248 VSUBS 0.009341f
C289 B.n249 VSUBS 0.009341f
C290 B.n250 VSUBS 0.009341f
C291 B.n251 VSUBS 0.009341f
C292 B.n252 VSUBS 0.009341f
C293 B.n253 VSUBS 0.009341f
C294 B.n254 VSUBS 0.009341f
C295 B.n255 VSUBS 0.009341f
C296 B.n256 VSUBS 0.009341f
C297 B.n257 VSUBS 0.009341f
C298 B.n258 VSUBS 0.009341f
C299 B.n259 VSUBS 0.009341f
C300 B.n260 VSUBS 0.009341f
C301 B.n261 VSUBS 0.009341f
C302 B.n262 VSUBS 0.009341f
C303 B.n263 VSUBS 0.009341f
C304 B.n264 VSUBS 0.009341f
C305 B.n265 VSUBS 0.009341f
C306 B.n266 VSUBS 0.009341f
C307 B.n267 VSUBS 0.009341f
C308 B.n268 VSUBS 0.009341f
C309 B.n269 VSUBS 0.009341f
C310 B.n270 VSUBS 0.009341f
C311 B.n271 VSUBS 0.009341f
C312 B.n272 VSUBS 0.009341f
C313 B.n273 VSUBS 0.009341f
C314 B.n274 VSUBS 0.009341f
C315 B.n275 VSUBS 0.009341f
C316 B.n276 VSUBS 0.009341f
C317 B.n277 VSUBS 0.009341f
C318 B.n278 VSUBS 0.009341f
C319 B.n279 VSUBS 0.009341f
C320 B.n280 VSUBS 0.009341f
C321 B.n281 VSUBS 0.009341f
C322 B.n282 VSUBS 0.009341f
C323 B.n283 VSUBS 0.009341f
C324 B.n284 VSUBS 0.009341f
C325 B.n285 VSUBS 0.009341f
C326 B.n286 VSUBS 0.009341f
C327 B.n287 VSUBS 0.009341f
C328 B.n288 VSUBS 0.020889f
C329 B.n289 VSUBS 0.021971f
C330 B.n290 VSUBS 0.021971f
C331 B.n291 VSUBS 0.009341f
C332 B.n292 VSUBS 0.009341f
C333 B.n293 VSUBS 0.009341f
C334 B.n294 VSUBS 0.009341f
C335 B.n295 VSUBS 0.009341f
C336 B.n296 VSUBS 0.009341f
C337 B.n297 VSUBS 0.009341f
C338 B.n298 VSUBS 0.009341f
C339 B.n299 VSUBS 0.009341f
C340 B.n300 VSUBS 0.009341f
C341 B.n301 VSUBS 0.009341f
C342 B.n302 VSUBS 0.009341f
C343 B.n303 VSUBS 0.009341f
C344 B.n304 VSUBS 0.009341f
C345 B.n305 VSUBS 0.009341f
C346 B.n306 VSUBS 0.009341f
C347 B.n307 VSUBS 0.009341f
C348 B.n308 VSUBS 0.009341f
C349 B.n309 VSUBS 0.009341f
C350 B.n310 VSUBS 0.009341f
C351 B.n311 VSUBS 0.009341f
C352 B.n312 VSUBS 0.009341f
C353 B.n313 VSUBS 0.009341f
C354 B.n314 VSUBS 0.009341f
C355 B.n315 VSUBS 0.009341f
C356 B.n316 VSUBS 0.009341f
C357 B.n317 VSUBS 0.009341f
C358 B.n318 VSUBS 0.009341f
C359 B.n319 VSUBS 0.009341f
C360 B.n320 VSUBS 0.009341f
C361 B.n321 VSUBS 0.009341f
C362 B.n322 VSUBS 0.009341f
C363 B.n323 VSUBS 0.009341f
C364 B.n324 VSUBS 0.009341f
C365 B.n325 VSUBS 0.009341f
C366 B.n326 VSUBS 0.009341f
C367 B.n327 VSUBS 0.009341f
C368 B.n328 VSUBS 0.009341f
C369 B.n329 VSUBS 0.009341f
C370 B.n330 VSUBS 0.009341f
C371 B.n331 VSUBS 0.009341f
C372 B.n332 VSUBS 0.009341f
C373 B.n333 VSUBS 0.009341f
C374 B.n334 VSUBS 0.009341f
C375 B.n335 VSUBS 0.006456f
C376 B.n336 VSUBS 0.021643f
C377 B.n337 VSUBS 0.007555f
C378 B.n338 VSUBS 0.009341f
C379 B.n339 VSUBS 0.009341f
C380 B.n340 VSUBS 0.009341f
C381 B.n341 VSUBS 0.009341f
C382 B.n342 VSUBS 0.009341f
C383 B.n343 VSUBS 0.009341f
C384 B.n344 VSUBS 0.009341f
C385 B.n345 VSUBS 0.009341f
C386 B.n346 VSUBS 0.009341f
C387 B.n347 VSUBS 0.009341f
C388 B.n348 VSUBS 0.009341f
C389 B.n349 VSUBS 0.007555f
C390 B.n350 VSUBS 0.021643f
C391 B.n351 VSUBS 0.006456f
C392 B.n352 VSUBS 0.009341f
C393 B.n353 VSUBS 0.009341f
C394 B.n354 VSUBS 0.009341f
C395 B.n355 VSUBS 0.009341f
C396 B.n356 VSUBS 0.009341f
C397 B.n357 VSUBS 0.009341f
C398 B.n358 VSUBS 0.009341f
C399 B.n359 VSUBS 0.009341f
C400 B.n360 VSUBS 0.009341f
C401 B.n361 VSUBS 0.009341f
C402 B.n362 VSUBS 0.009341f
C403 B.n363 VSUBS 0.009341f
C404 B.n364 VSUBS 0.009341f
C405 B.n365 VSUBS 0.009341f
C406 B.n366 VSUBS 0.009341f
C407 B.n367 VSUBS 0.009341f
C408 B.n368 VSUBS 0.009341f
C409 B.n369 VSUBS 0.009341f
C410 B.n370 VSUBS 0.009341f
C411 B.n371 VSUBS 0.009341f
C412 B.n372 VSUBS 0.009341f
C413 B.n373 VSUBS 0.009341f
C414 B.n374 VSUBS 0.009341f
C415 B.n375 VSUBS 0.009341f
C416 B.n376 VSUBS 0.009341f
C417 B.n377 VSUBS 0.009341f
C418 B.n378 VSUBS 0.009341f
C419 B.n379 VSUBS 0.009341f
C420 B.n380 VSUBS 0.009341f
C421 B.n381 VSUBS 0.009341f
C422 B.n382 VSUBS 0.009341f
C423 B.n383 VSUBS 0.009341f
C424 B.n384 VSUBS 0.009341f
C425 B.n385 VSUBS 0.009341f
C426 B.n386 VSUBS 0.009341f
C427 B.n387 VSUBS 0.009341f
C428 B.n388 VSUBS 0.009341f
C429 B.n389 VSUBS 0.009341f
C430 B.n390 VSUBS 0.009341f
C431 B.n391 VSUBS 0.009341f
C432 B.n392 VSUBS 0.009341f
C433 B.n393 VSUBS 0.009341f
C434 B.n394 VSUBS 0.009341f
C435 B.n395 VSUBS 0.009341f
C436 B.n396 VSUBS 0.021971f
C437 B.n397 VSUBS 0.021971f
C438 B.n398 VSUBS 0.020889f
C439 B.n399 VSUBS 0.009341f
C440 B.n400 VSUBS 0.009341f
C441 B.n401 VSUBS 0.009341f
C442 B.n402 VSUBS 0.009341f
C443 B.n403 VSUBS 0.009341f
C444 B.n404 VSUBS 0.009341f
C445 B.n405 VSUBS 0.009341f
C446 B.n406 VSUBS 0.009341f
C447 B.n407 VSUBS 0.009341f
C448 B.n408 VSUBS 0.009341f
C449 B.n409 VSUBS 0.009341f
C450 B.n410 VSUBS 0.009341f
C451 B.n411 VSUBS 0.009341f
C452 B.n412 VSUBS 0.009341f
C453 B.n413 VSUBS 0.009341f
C454 B.n414 VSUBS 0.009341f
C455 B.n415 VSUBS 0.009341f
C456 B.n416 VSUBS 0.009341f
C457 B.n417 VSUBS 0.009341f
C458 B.n418 VSUBS 0.009341f
C459 B.n419 VSUBS 0.01219f
C460 B.n420 VSUBS 0.012985f
C461 B.n421 VSUBS 0.025823f
C462 VDD1.t7 VSUBS 0.225493f
C463 VDD1.t0 VSUBS 0.225493f
C464 VDD1.n0 VSUBS 1.64803f
C465 VDD1.t5 VSUBS 0.225493f
C466 VDD1.t4 VSUBS 0.225493f
C467 VDD1.n1 VSUBS 1.64709f
C468 VDD1.t3 VSUBS 0.225493f
C469 VDD1.t1 VSUBS 0.225493f
C470 VDD1.n2 VSUBS 1.64709f
C471 VDD1.n3 VSUBS 2.94087f
C472 VDD1.t2 VSUBS 0.225493f
C473 VDD1.t6 VSUBS 0.225493f
C474 VDD1.n4 VSUBS 1.6458f
C475 VDD1.n5 VSUBS 2.84192f
C476 VP.n0 VSUBS 0.053871f
C477 VP.t4 VSUBS 0.215077f
C478 VP.t3 VSUBS 0.215077f
C479 VP.t2 VSUBS 0.217588f
C480 VP.n1 VSUBS 0.11332f
C481 VP.t5 VSUBS 0.215077f
C482 VP.t7 VSUBS 0.215077f
C483 VP.t0 VSUBS 0.217588f
C484 VP.n2 VSUBS 0.111338f
C485 VP.n3 VSUBS 0.098565f
C486 VP.n4 VSUBS 0.017871f
C487 VP.n5 VSUBS 0.098565f
C488 VP.t1 VSUBS 0.217588f
C489 VP.n6 VSUBS 0.111268f
C490 VP.n7 VSUBS 1.7573f
C491 VP.n8 VSUBS 1.81019f
C492 VP.n9 VSUBS 0.111268f
C493 VP.n10 VSUBS 0.098565f
C494 VP.n11 VSUBS 0.017871f
C495 VP.n12 VSUBS 0.098565f
C496 VP.t6 VSUBS 0.217588f
C497 VP.n13 VSUBS 0.111268f
C498 VP.n14 VSUBS 0.041748f
C499 VTAIL.t8 VSUBS 0.20494f
C500 VTAIL.t9 VSUBS 0.20494f
C501 VTAIL.n0 VSUBS 1.36423f
C502 VTAIL.n1 VSUBS 0.672302f
C503 VTAIL.t15 VSUBS 1.82796f
C504 VTAIL.n2 VSUBS 0.809045f
C505 VTAIL.t7 VSUBS 1.82796f
C506 VTAIL.n3 VSUBS 0.809045f
C507 VTAIL.t4 VSUBS 0.20494f
C508 VTAIL.t2 VSUBS 0.20494f
C509 VTAIL.n4 VSUBS 1.36423f
C510 VTAIL.n5 VSUBS 0.709932f
C511 VTAIL.t3 VSUBS 1.82796f
C512 VTAIL.n6 VSUBS 1.95099f
C513 VTAIL.t12 VSUBS 1.82797f
C514 VTAIL.n7 VSUBS 1.95098f
C515 VTAIL.t10 VSUBS 0.20494f
C516 VTAIL.t14 VSUBS 0.20494f
C517 VTAIL.n8 VSUBS 1.36424f
C518 VTAIL.n9 VSUBS 0.709927f
C519 VTAIL.t13 VSUBS 1.82797f
C520 VTAIL.n10 VSUBS 0.809032f
C521 VTAIL.t6 VSUBS 1.82797f
C522 VTAIL.n11 VSUBS 0.809032f
C523 VTAIL.t0 VSUBS 0.20494f
C524 VTAIL.t1 VSUBS 0.20494f
C525 VTAIL.n12 VSUBS 1.36424f
C526 VTAIL.n13 VSUBS 0.709927f
C527 VTAIL.t5 VSUBS 1.82796f
C528 VTAIL.n14 VSUBS 1.95099f
C529 VTAIL.t11 VSUBS 1.82796f
C530 VTAIL.n15 VSUBS 1.94512f
C531 VDD2.t0 VSUBS 0.227435f
C532 VDD2.t1 VSUBS 0.227435f
C533 VDD2.n0 VSUBS 1.66128f
C534 VDD2.t7 VSUBS 0.227435f
C535 VDD2.t5 VSUBS 0.227435f
C536 VDD2.n1 VSUBS 1.66128f
C537 VDD2.n2 VSUBS 2.89116f
C538 VDD2.t4 VSUBS 0.227435f
C539 VDD2.t6 VSUBS 0.227435f
C540 VDD2.n3 VSUBS 1.65999f
C541 VDD2.n4 VSUBS 2.8261f
C542 VDD2.t2 VSUBS 0.227435f
C543 VDD2.t3 VSUBS 0.227435f
C544 VDD2.n5 VSUBS 1.66124f
C545 VN.n0 VSUBS 0.110245f
C546 VN.t6 VSUBS 0.20924f
C547 VN.t7 VSUBS 0.20924f
C548 VN.t0 VSUBS 0.211683f
C549 VN.n1 VSUBS 0.108317f
C550 VN.n2 VSUBS 0.095891f
C551 VN.n3 VSUBS 0.017386f
C552 VN.n4 VSUBS 0.095891f
C553 VN.t4 VSUBS 0.211683f
C554 VN.n5 VSUBS 0.108249f
C555 VN.n6 VSUBS 0.040616f
C556 VN.n7 VSUBS 0.110245f
C557 VN.t3 VSUBS 0.211683f
C558 VN.t5 VSUBS 0.20924f
C559 VN.t1 VSUBS 0.20924f
C560 VN.t2 VSUBS 0.211683f
C561 VN.n8 VSUBS 0.108317f
C562 VN.n9 VSUBS 0.095891f
C563 VN.n10 VSUBS 0.017386f
C564 VN.n11 VSUBS 0.095891f
C565 VN.n12 VSUBS 0.108249f
C566 VN.n13 VSUBS 1.74433f
.ends

